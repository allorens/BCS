BZh91AY&SY�՝��o_�@q����� ����bL]�           {�RP�UR�R��*���Q�J�R��(�T"�*��H��J�*�H�UQ5���ITR��@*�h ���BQ
�%�T�@�Jh��UBUJJ��J������B�%v hT�%B�����fد7IP���0d0�+�f"�I�l�D"��m�h�(��$)U	$�$R�R�AJ�Q��Psu�@� T��� �u���2
h����-O� �И�ʱF�Z6�aZ�))�f�)��ݍ� )���T��%���Kϒ�� cy��)ERq��z{��S{D:��%Iw����)%g��=̨֥��ꪪE)w����*�*��=�J��
X��Ǥ���ך��J�/mU�z�@�
�m�QB�H�[�)@:���HQR���{�UT��<�AT��W��D�Q=�^q�WjjH{��:�*��Y��z��R ���GX�����UR�I]��y��]jK��P�EEP^�UI��T�{�p}E���u�w�����O�zU	!x��*�ԩ���*��A^{}�zj����ꤢRT�K�꒥J����z�T*E�+�=GY^���R ��T�)T���(� ޛ�)T*��y/{ʮ̅
��>�TD�@���J��l�D�J6
�G��JB�+ޕ�B�J���R���*�UIΞ��RJ��RD)�R��S���l��B��
+�>���y���U���:�**��s����\�۪��7*�UP피�v�RURU��+���Ug��@w$��J�
D�R�t>}T� >��
8�{�����P��=�=�7���V��� s�� �R竝T���(u�ˀr�JAD���*E��J( 7��PR�ÇB�ur�� ѝ��ܮ�[���{�@{�L��{�z��[`�������$��Ԫ���$��E  ;���#���m�àPs��(-�}�@�:
nV�k@0  �+ lq�� r��HR*H�P�y$�@ 7� � q�rTU�K� ���� ��x z�a�
��Y�< ���:P8; tP��N8����*�       L%)T  �b` D�щIRP      O&AIJ��L�0C  �O�RTɤd2d�hѡ�@��JR#*� d�   h �j3JIFFA4��CLLC	�`���?{��g��?t8J��T��ߛ�����ʬunϜ�s|7������*��J ��b ���eTW���b�@_�<��?@o��_?� U���$�O�PW��T�� E���?�������lb[��2�6��6Ķ�-�l[b[cl`�l`��6ĶSؖ���6��%�-��l`��6Ŷ-��`��6���m�l�hm��%�-�l`���b[Lb[�Ķ�m�l-�b[��6��%�-�lK`XĶ%�-�lKb[ؖ����:e�i�lK`[���%�-�c�Ķ%�-�l`[��Ķ%�-�lKb[�Ķ2ؖ���Ŷ�m�lKb[-��Ŷ�m�lKb[�lcؖĶ%�-�lK`�-�6���lb��6�L�%0-�l`[���%�-�al`��6��6Ķ%�-�2��Lb��6��%�-�lK�Ķ�-�lb[L�0m�l�6Ķ%�-�`��6Ķ-�-�lcLKb[Lb� �-�-���-�lm�l`[���6��LK`[���%�-�ldclK`[ؖĶ�-�lKaL#b[LKb[ؖ��%�-�������-�lKb[4��1-�lb�ؖ��cli�lKclb[b[����0�1�6Ķ6�ؖ����%��cl
clKb[���Fؠ�KbF 6�� �[bl@m����
���(�V�(�`�lB��[[b��(��Rؠ�`�l@cب�[`�lm����*��Fث�lm�-�Q���R�� `	lU-��[bl@t�R�*[ [`�lQm�1�6�Fب[Kbl-�%��
��0��T� 6���Kb#m��*6�� �`�lU-����`LPm���Q�"6��*[����A�6��l@m�����b�lU-��� 6�R�lP�Dm����*��� �b�lPm����T�(��"��T-�-��([� �(�-��lK`�l b+lEm��lQm���-��l�Fت�`+lb#l` i�l
`�[؂��*��-�������
�[ [b�lDKb([[`lEm������`l b+lQm���U�*���,` [؂�B� ��*��1Q�"���*6��"6��(������� ����ض��ؖ��`[��m�l`����-�l�6Ŷ-�-��b���6Ķ��`Sؖ���-�lKclc�ؖ���-�l`[ؖ�1�1-��m�lm�lb[��b[ؚ`[ؖ���-�0�%�4Ķ��%�-�l`[�%�m�lK`[e�#ؖ���m�l1�%�-�lK`�ؚal
b[�6��%�-�lKm��`[���%�-�l`�)�l`�lK`[�Ķ%��bS����b[clbi�lb�ض�1�lb[ؖ���-��l[b[ �!lB�S`�L`�ؖ��m��%�-�lb� �%�0-�lm�lKclc���%�-��[`[����Q���q����#�fX�����|�V]�y����ڣ!7�iE�����:�fD�8�d�-9/MKiӃZ�
�t�m�MSN��c+�^V�K�Eᱩڠ��Z'0V�j�٥*�Z-y�c,2�'�%�15ا�D�	L�����0��ö��i��f�op�Ȍ�Wgv�hi��,�J�Q�F��I�]Br�v����-UlZÓ��vb�d;(H��y�&�b#�7cǈ^�tMZɒ������(n���L^��(ٶ�6�[A��H�m��]y�n�eqh�2RW�m4�I
�J��e���E�:��!O3QfY�b��`�1Z2�9�x�Έ4\�������k���ʇm�2aag.���Շ������y�oZ���)�z��p,�[�rἽ�2�M٫wAOi�l���]j�N��^o-��K��F��Y��HZ8��U�U���{Cm�T0̔ǂ�0+D��ʭɣ%�,h�ʪۋWvl���f�K��2�+8��b	e�,T�����`;� �*f3�eDǥ�M�a�wwV��v	��e$©�14�e[��Sm1 6v�+F���V�����f�GE��!��4�主�G��η.i��U썲Ҁm�թ�i�Dӽ��R������a*Z��y3)��[�4M�
���z4)s"��nA�[���/5�n�"Շa��Ef��H�.ڢ^����&+�.;Y��O!����nX�(%�%s-�ޥ���"�m(B�4�ت�1[YG5�L�A͔e�*��Ǵ�t,�,h.�nX�V
��%�b��jY2^-���&�[��b(���M@a��4��*�գ����{uk2�:�S]�e�j�ʤ�Ree�v�LmJ�3L1Y9d�[��Fm�cL�aVjL�MX��m�m��J�S�)���dW��u�P-���x.�Y�����t�N�� ��YrL�Fd�n�m%nf�ӎ����;gV`�\ʓ2�8mY�&d��ݨ�����ZS�b3e]ѣh�R�Y%�94
�tޚPۧH��v�3K��{���6���,��*.Y�t,�X�����l�CoV01ۡ5	
(��i�H����A�#)L{[IM;���]EM6��P9��٧\��ռp�2��A���X#�f_t�۫ј������A�#M+� -���i���j(�*e��5]\�u��rkw0;�2�Z%�/5&�v�k��S	�B�V��R��B¿m^:I���b�z�t:��Օ��TV�5��bl���O5b��<���cG/e(̆��
w�K
`=c+N+���6��J�S��9��;_UإE̓i-j
��C��*x�(��v*�8Ԉ
QZ�X7C�CV&"Nb��2ͷ��1Tx���k*�eb�+(�tNE��zܨ��'75��R���v�!��]�%Y�\�J�FT�XF*�/x*��w�R����-,�j�\�6�s8eջ��6S�KE�+#"���]at㼰�ej��.���z��S.� f��R��i�3a������@�f��瞘�j�+:aI]dx�;u�0u��f���7qQ㦚n��3�V��1TU{�d��:<q�#�(;0wv��.�G�c�Zb�*?r�`�m�nȚQ*�f��"�t��r�"z����Ż�����(�
�7��T�YRm<ʂL)��-��I��{h���@�*��	ڂ�Rf11mbj=�2�UT�Ly(VK��^�\x���$3�m�&=(��ՋU�cr���b� и�ѻUDj"����Viݫx�w�Zr�w/p�'MO��M����S�8�Ѷ��Td˅emCx�&���a�];�J�V��2��e%��B0l]仍��·�NM;%�ʉ̼t���oE%�,�u�6�p�N�n^�9��ʤ�[E�z)̇+=O[tN\�tY�h͆�ܪAf�q��x�l�k`\�F�r�&%ַ���"C�Qh2�]�JP+@����PU2�����
�J:(n�"5m�q�����&���6�����0�ؙ��,+xt�$y�H�e�����w�U�+D�2](6��ъ�K��GX��jX�1R������^j9��$��D�6��v�Њ��ګ��u�sn�ؙ"�[�
�*��V�GM��%����M�eQ)�=~xB�z�v�9�'1V�	7e�q�fƪɠ�q��։�M����.�S�"Ĩ7f[Kq�0����FA`��xoi��,��+9�aN`�ۚu�֪�	�V	��q	e�Xǻ�w
+Z��$���3L��BCv*�ф�B�ʐ�J�ѻBȁ��$|��6�չ�����;u���l��#	������X���jۻ�ׯA�H]fE�MƎ6�I]*;m(T�)�f;X��~����!���5D5ۈ�Y1��^�S]�ۈW�2ፉO�L�Mҥ��� ��Җ7�2E�{��V���� ���G�ƪ��h���41.�<ڵakj�c�9���6+Y��d�P�Q��/����n�2��ތ�knÂ��126)8�����-��휆ȣ�?�{yd0`��3s*ʌfn�j�f2�h"���W����c'vˤ�EՉ�#��;�Ș�x���d�%j�{���$.Jy%*-��Ļ#[�pc.��4^M�2�b�i��3Q�J�2��{z�%2���j����6��E�ױ�&�` ^tY{8fT��5���S�x`�����ǘ���9X1lBB���wNm����')�ؚ)a7tS��S̪	�:�v �kj��x �[N���ʡ�ZH��ZiI&���O.���B�d�3c��֫*Z��Ob���j�8�ѐi�q�1@��v3%�T���r���ĻZ���Md�D�%J/�#�Cm�
�j�p͚�0�\�As�-�z��V�	-U�bVd�$��[Zsn�8�$!o�e�:nLԆ�g�5j�D�B��W��������צnU���!�Aʹ��h��K�KK�TJ�.hM^�%���Z�3t5ZM6�r�-�M[$`�f�f��N�8��5�n]�r��r��"6Tr
��ŧ�˧���
��Д]/$J!m�P�0,�s�Ai�H���+����.n�������dS&{nΫ��tD1���!eh�PX�R�Mu2ۅ4FXl�U�%8�����oJ���8�Mą���nDc�Su���0m[������x�/�X�1���a<-�B�U��n�J6�M��Eԏ(fS�ң�F
M5�.Σ�F���� �jP۽%Y�:N���Y�$���Uj��[^m��H��NΪW '��z�dȓB��l�Pw1ڊ��:�
�l��3���Y�i�ʎOγv���c��굪�]�+sQ���u�M@/f��V��I���	b��;֭3*7�BR8A8��\:&^%b�hH���a��HY�W��8lI��ac���L2�5jz*�/Hg[��I�+y�=�y����$ ��I�CNa^� �#�r��e'0�#��,����3b�Me��$V�h���FV�z݄�������m��(��+hS���*�fV��`$�NX�[��P�x�ݫ0;u�m[@Y��M�Qݽ+fE���v%U�l~A�3;.��u�j�5��$n��w�`�K�ɢ�dǎT���Ĺ+J���'U(��ǹ���bV��Nh����o7�U����",V��|�D1e��z�t�mIYJ]�G-���{�I�Z�() �U	�aҜڗ�v�q�5m�enѢtq��)��J�d�ie�d鼩�eäj P�G^�JY�n�m�n	�݉�c��z�uY�GX�5��J����4`6��̏5QZ��c[�&=x4,F���.��\9��ٔ�[ǵhyO�Qgd��,�&�.����V��[n�Gt�`��t�,�ո�n[����f�J�:�P Lge�5�d��+UL�۬(w�K͢j���ˑ�hk �0[����P�-'�����.��
U)�v�2�{kg}�Ֆ�a3-�"wqH`���c0�vK E�e�㗣���@q*��*�w���/*��h�+c�p���۫(ֳN��r'cS��Q�.Uơ/4{7q-����u6�[�f[�jPRյhI%6�u%�7Zk���rl-����ˢ�.D�Zj���̨P"=�(h�"�h���֧��T��2��ds��Z�xl���yc(&�Z,�6m��,w��YX�Kh��(��dG5\ǚ��Փ[��b.V�	���F�oAv�"�yjM�nIoE�E�5Oq���ת�.�0(P0�a7D2ab˫o^�tOj��ee���-T,��@0�r��[�QC-;!�yr��.�4^�ʎ�KU2e��T���{�)*�KM;�F�rӨ�Ӣ�\z�{`V�S���-�8��i˔a��7��5�)A��#�"H�Ӣ:��L����VRܥYvFcq�7M�ҥ����J6�1�*��7h�ˈ�,V��8j<��F��B��
�bњ�r���~��e���A(Pv��l����vZ5�)&�)�h�c��D\t3#m�8�h;�2�+�-n��X��� ��������uO]�D*�~�I�:�Nԓ$E�еa�P��.Y�i䈦7*��۱%.�vKWh�[6D-b
���v�4g��7�J�	5�0��m�N&E����p]���c�M9B��9�e���i�n���T��L�}��gek.e�,�5��$�@�"� �;I�;ze���y�t�ۡ[�j"�h��4���Bf���V��ɖ㼸�Z�3j�G6$jy 7KM�ҥkDeg��z%�dd��#�/R�*3n��6Mۧ%���a[�i0����ש�3/aR^��V�٤��T)��i��&�oM�A$³P���܊�vw$��(�wUmi)�:�Ź�dCf�AI��@�ݏq�x�txr�]�2�d�uVm�ue��
�Sam�A�sUݲ	X�����8�`��R�9+T��"��׫uZ����jB%�p�R-���%V�e]����ZoA&={A����["F��mĳK���+j\��*�ej�W�3=Գ�P���
�v���B�H�n(�-�e7W����v���&X�R��n�XB�$�y�l\������i<%�v����#[@Sj^�V��09��ð���)��x2������z�k��ǣS6��h����V���U�r��q��s3n�-�cNް�*w��b2����;ͨúm�
TT5)��k�B@�ق �5!Ӑf"[��yQ�� ��h޻t#W6��`vհ�+�t��M)fF����Z�B��VH������E�@�K1륨e0��Ec�z0 cҢ�8F�G.��|�{�{;�z�qf컑�M1w,����׳2!�0M����o]�Rܤ����#�5�
��2�Tj�m�h���
��s�d���V37-�U��Z� ���U<�o�T �2��KfC0�66�ц�����/"�oSYV]�p�eMo���%�b�ù/�����*�`�E�*^^��ˑ
٨?=���Ct�]���*{^���Q���k6
qn,���^J5`GS�0fnfA�Cv�j�J��ͧt;2x��v�B��nXu�H�m�=�ª?]����YYc[�@j�3EE���1n�R���iDͬ4T�4a(="1�xf�A����j����v���^ȭ���Wyj��mD��HvQ�*�[��)�P�bQS%bN��fP���U$u2c�����3[!���d���ދ�����Q�n�Dܴ�3h�T]�fʹ��u�����{���@�[N�(�T�I�&��v�gHE�5��H#�m
��T��8�y�4�uHn��r��w8Pf�KQ�X���[b�EV�"�d�Tf�(�n�v�7�Q�{mQ�'}v����6�9�v�%��ƴH�C�i��(�Q*I4�T��ȅ]��J�b�B/��Yi*���H�J�yQm�m!e�9gkKͺY�lZ3'Q����ą�jx�PJut���3�������aQ�w�F���y+B�V(vc���^̔}��r�]@.ʴ�-�.E����	n+��SY@-����t;J���
,`6�){p�ռ�D�RL�8�Q���j��5k�ԒI�j�*r��;��T�ɋZ���5�
!��$��BRv�#�B���[�B�ͳi��Tӳ��OV��J��������_%I�iPW��I\J��iL]k�ƍ���օӴ	m$�!o��C"x�{�ޥZ�%ZZ��ri0E�9`�R��e�-��7A���]����F2�d�؁ʧ֝�N����\ q/�����Ī7C�&u��n��I�͓��+�ZТ	%KgP%8�#3f�V�'E����ǫ�+���(�Z�.}��D"T�R|�ܻU��f�����}_<x�%J$.�U6)�*)���Geхd=[�Pݻ7\RM$���jk��G�]���/^�D��1�"�ꘅ-k���9���9��!�n]ǉb��cSP�a��76G-�L��q!g"KC�6AT��$2���tR�MT�N�J�E�,q�e!��Ň��W;m��ґ6� �簌�����JKʊ���W�i*���rs���bW'H������[��*X =��*D��;W0��o�r�S z���jIU����e1@a3��E���o\C4���q<U.a�oƍ�:Z՚�Z����k���Bj��!Eh2m(�຤�$F:�.TR%N����*fᎈ0���B�ZHqB-&�hq���^�b��Z��,5�4�J�-J���%ņi��ԡ�������~������_��`���7������'\����/��z��G%�o�`�Ӓ���~�ж�V�C�3��XT5�	[I��mvǝ����Nb��#��MG�@�
;|��kB��15��}c�V�|�5�i�Y�H�U�n7ݗ�֛������f��;Ʈ��@�-vq�G8>}��Z�j,�{@9��<�j�d���樎wG�n���-�t���v�׉��	��nA"�ը��S���%q�D��	�;�S��[�3���v@��%����u(s{�@��N�Tp\�ĸ��0�1Ҁ�]}�S��vTSA�'v8b����s*^M��XP�+Ŭ����ev�yH��eVV����eڙ���\��%˼��*��<V^�ι�"Vڃi��5��u�^�Cc�.���mTY�Ȋ��M�/�j[��iu�0T�,:y�u|Lo��ܠ�W�+��Q	t�1nvhշ���MK(�WT�I����fZ��mq�����P�]�yѝ����j�^�Մt�ջFim����M��
BAٛ+hQˉ^��8Ҁ@4a�_����-bZg�홨���do�v��I���t�u��7�/Aw�T�5��9�w�#s4e��<L�±�I�'ZZ��@S���qN]nf)�;�7ʐ�:�\GaU���tx9�v͵u�ӓ�
�ٷ��;x��˝�T�a�z
��k���*�n'/��׽��V�q6&-��j�c��hՌ�;^��.˝��e2�bCh�2�
��KG�5w5rD�]���`G��sm��������h���C��%����I�x}����K��dw0j��9������:��܎�T7�D�k��<t*	e_m�0�FÈ�݂s�ژ���T�0�K�+��v�:%�}��+pm�m�5���-���{���ze�ׁE*�5���˽�s�S��ՙK�����������Z�-4��dZ������c���Aj��|GR���|3�H�F����U%�9<�2m7q����Ō��J3/��\ھB��ܱ�9�`)3����f֨�����x�W@���P��p֭�m#�v�m��l2��"�=v��څ��z�Kbx�'��}ʢ1ҫ�T7�n7�v��˦޻y�<0(��sRd�Ӕ�U�y��|�B_7p��,�/(��u�f�#wۧ��om�/���|r�qCj�>�:�0��44_u����M
"�
عm��wt��ڻ���.���+#u9XWz��+2f�C���(��'v>��.�H^���'F6��[���x1Kw������ԺQ+�Ҳu���[1���h����{�4��V�pŇ2��-�"�{q�s�iDZ�N�x��56��w:��^ά]�ZF�i�,�Q2�]���;O@�6�_;�J��8���=j��T{N���:�,��W��e�Y[n��sq��+9��g��V��`����V;�؆���_bFs�?Q�]��[ݴ�nܪQ#�)N"��-K�����[��Q�rIYؼ����a���g+e/3�eM:�,��if�E+�iH_TCu�¼ȷ5�+*#0N�5ԩ����4
C���b5�6�q')�ż�:�^�}������2:�����E�� vm��x�6s`��g��Y:�ME#N��<�b��#�f�_eZ"��2��F��+�r���q�U�8`\.���o���/��N�!l���ك:��5M��	k���j kV�ܷ5��f�hR���{�/u�7���ɧ@�Jgr�7�]�L�6�]DNH���u U�' m��ೠ.���Fi�;��׬��W�9q���<���9سj��h��8�3�&	4nЦ��}	���:T7�ğ^y����3q!܃�czm����kGQ�j$�4k�>�cb6�lQj��(j踔�U엜D{Ԅ����=�	��|Q�ä���\�	�&��{�e7]}�r���&��-6%#�U*2u����Z�6��cE#N��DL��f�9�tj�zm]�m�J%��Л�����B���xHhQ�mf�^U�`\�c7��L��	�L��;G
�^y2B�W&V1��t9qV)G�*�~S���]#�ۘ���])o�=ga^ӯqfY�]�yo�j)Ȫ��%j�J���:Oko0j@�
�#�r�1T;�����ݬ=��s�YC{{���$AKɭ�(�ӗa��s'`��v�
��h-Y-��W�FS�^N��	�n�n���F'IBՅ*>�4PlE�,vf���y�0��6�Ayp��w��yJYQ�is5g��3}�9����{}w3F���Xq��tWX��y� q^̳qֺZ����U�*c�e9/gVx�3��8�e��ܑZW�Gu���g�tC��:ۡq�N��V���CPv�pΝ�������������᜼&��{8�o�IBEa;�
�c�7^�Gu%vd	���;�'W*�}�]�9`x���,�D�¢�c��꜉��9z^�ٴ�f���]e��P���<�[ʀ��v�\��0ÑU�|����9])�?v	�ta`�����x�l�r���fV�֛�hwYd�7�x-q�6����U���ݢ������3���o$ա�Ur��%p��,�yis�����Fd�kvi�9D�ָ�C�"�ݝ3�\]β���؅΢ �W]��ݗ��C2�ԩ4��S�j��%��w�{kfq���X\�8�]Wzm#��3{Z���	�Kq�p���u�wf��:3��U�5{�e;XL�]+:�飦H$�h��A'NWr�v�:6ŉ�M�%y��>�`���:�opn�dP�d���Ϋt��$�,�.�_tsX�l���rsiQ��+�8�n�[C1<���u�oC���j�����a�:�Af���P����S��Ы����b�|��^6�ԽB��vq��WVr��K�7'+�0�Wp�Y|�Y�vإ����o	�.v�<��b7*eS�ӣ��Սի���3�8����af������P�Y�^:p��C�m���ǌmءʇnG�儏�]���}�$�}k�gz-�rI�(^�*���R$2����H�@c�I`�m�b=Xh�{�+{���!1◌�����w�ZW,�����;Lu<va�g��)[Zw\ޣ�I�l�T鱛nN�i�W�I6��[YY����zd0y��b���V/�9�D֎��^R	�����C;+��^;������P���WE�`��=ˏb������ׇ"�-�ǅKm���VH4%�H�n"#��u�����;=��^�U'.�Dmb�@�%��/ML���n=/{��;Q�lqn���ٵE0d|)�ӗ��@���d9�%�}���(�������Uw��ʞ0���a'H�I�K�+	��+A�����΍�]b Y��mp�D�[ܴf�fn�̨�m�n�4BK5��.�h����'�H��+���Ĥ	�Bg%���k�	��N�%�Sn��;s{�d]�w`�:�*�C���s�L��T��&\�ٸ�<��ǝ��w���=�"���v��Vu8��D�H�4q��~u�'.�*�4a�H��'�������y*k�qfq:粣�
d�	ӝY��fn�\��^�)E�<�&w5�9ǐ�G�mZ��/t�,Qe�̶�(���tN��;]1�Jg���y�gWd{�gf+�.��T�8�h��Θ��w8�
���E��is)=���,��f���S(Rz�ޖLrWh�V���q��'�_l�80�����OE�5	��@g��DS��WJӓL��|G�SQ0l�p��+�Z0΍��;���g�Q���v���i�ά�m���۬�6�(���+^����u�`}-���"��J�V���W>!�.��_�$�v:�7ob�Z�A��Y��!˔�`��."u����]L�a��=��$Sk`�Q�Z*�n6e<Mu��I+M��T9�+��a�S�soȔ�"e���0�Xq�w	��=qJ[�I\{�W�@��"�G��0�ep��|�_:�r+��sܛtꆧ,ʀf�F�)���<z�����\UR︡S�W���z�*tZ���䃕�0�)��w,���W�+�e\컲�\��i XR۱�N�%N�]��앚D緉��H���<Yn�J�z
[�����ne�ۿ�q��u��o�G
|�5�2��ݎ�$$���R��s�p�,֣�gd�[�@��؁n��.{�ڗ}�ʮ����!��w����Hl�t�3�\�w���,k�Mfe	�^˛�r�&�^>�^�F�>ɚ��ԓ��-�S6_6mWn#6elCh,g�|kcZx�ێmݡY-8�}���uc낹\�W�]�ɷ�6���D�Ѓ�.��Y���)n"ũ���N���{j��q�c1�l%�q���<�x�nd�*��g)��>�,���rz$ܨ����(��؝�r�^T�sģ(up��RR�����jJTꊚ�Q�L���n�ҳV6U�&e�$�{��Ν��2;��WF	�ٹ�%���.�[�s��+��]�i��'7&�2�c��������Xd�U���<�1v0�5�
�a�����_u���oH�*�
���D��9nmv��������$JE���S��oclY�Ы��د�5Өgl��t�{��!�Bʏ�v�G@��E%�,�3�n.��k1�ڹc�5Z�pr�S&b��(r{Ԁ+�p��X+e'gbY.d�l�B��m�
ު�Qb���IY����G��jK��_W5]�d��`�o�11�Ոg=���p�U<W�<n����xZ}�6��o�4�$�C��� 7�0p0��˲:+�6�Yǘ-���˫q�Ѡ��f!1ޑ����]��6v��y3�&2�c�3w��<]�D�-��k��f8�����݃���TB�:u�d��OIl�=�,�Ю����U͗N����'��8�E��Mu���s��-�[0�5�V :��Z�y�+��洺���\o�O/r�8��f�3�^)�q���tEeܰ)���=; �37k�\).�ɹ�NFb=�YLF�h7u���P��u_�;����qC���7�q��6�G�10�苨b̐���Va/N�G ��åt�����x��Z1,n8Pr�����[.�D�:�R{3d��Q���ҶK�3#�:I��4�Z
	�t2�[^��2:n����[2�N����XVk������p��g�<�t\-`|��h�N��E��S[ٕ+o/�-eJxA[��4%wb��iVȴ\'Kz�%����F��֗e@f]s�_�����U[��B�:MV#��	����v�u�ynU^��`�]F�L�iC�^����ѥ̖�Z��<�A�3n���^�H�0�*�f���{-!�Zy�u��O��,�R���V9�8Px.��$KTD
Lsg3�����թ���LF���m�ς�
��Q���$�ΜU:��|��0��!�,2꧗q�n�A)�ػ�W�۔��Y��^u#��ݶepd���1��F�&��G�iY����Xl�����W�Ũ�֪r�&IS�B������N�R�r{&��uH2P}6�`������t��yʜK�˳}bon�s;��Sx��l���1fu�8.��t�Br���7��x_H	*�P���Vw[}ۜ�fd������[�Z�0���q��r��l��"��]b���Z��ǫ��f�٨�d��t$Y(^l,5zb�{R<܇qE��{�#,�I�-�7��ܹ)呶��̥ϥX��a��{�6��m��^�'�s�
<�T��sP�h��"��lf�W��Z::��.w�Nַj��&Z:"�+��W�Y��*	�3{.�xI�9pyӳ��oŢ��@�=�8-'"@t��ѥ����f��e\@�7�nuf��v�o;�鱀���R/yPz�ޝb]]�)Ӡ1���z��1g\�$�5zN�K�Ud���-�z����D�Ν�8�j�X�J�����̒�B26�O�{\9���2h�T3[�F���U�N�ƗQ�rDL��Q�t�QXei�	��H���i�(^�D���`�2	��&���U's!�(�yx��Y�v'�*~%�I
%��~n���<銋�[)	DUm:F�e��8q��2²%u0�4�6� ��aP�K]L�4�n�C&H*`�l����ۇ�F�%B��O#�(Z��߬��8joj8�
��6��F��|�K4�n�U�,P����v.���xZ��#K=NQ��.:�8�x*��k���E�-ۆ��3J�&tEASn�c�e��\Q�}*)Eju��UWR�"q�˳f�� ����mq�n�v]��D�t�#F)�@���D!-L2)4R9inU�Y�(�W��y��p��l"Pb�Q�  ��V@!�AV׮Yv�ՙ����d��D�,�!�S [7���ZR@�r�H�L��J�IKM-���^��KT��g���k�Q�.z5�pn]@�a0H��m��I��a�l6�O2ۭ�!�t��P6���#X�!*$$�I�I�J����h���b�@Ͱ���,P+U�@078�He
�a�i��q��K�f���R���Z�ДH����TY�0لe�Ih�r�W
֤�W􊠠���?��ڈ�(|�p�o��E?���PPG�����P��'���/�G�G�S��u��D���5�Z���RoV
�ڻ�������ݨ)�:y#��� $���Q���s/Ű�?u����FK\��t�싣�B���>�:9-����s�6wVC�هx��eJ��c�tnL��M��{��l��6�g9��r;xv>ap��v��b/���[�R� �3-@���	�W(��uGQN�אe����6�Ն�X�ƻ���F[2��N=6�M��1��Y[p��67�Y\��E�RWF#R�ө3"=4���vX��\U� 4�ayb���C]�K&���g0l�
�&��e)�;f���c��X��Ղ�w,*��z�P�L)t�X�/M`��{ّ�8Hҋ4:��n��8C*�}\7�Yƈ��]#��5%V�����\��%J�,�yJ�$jͦ{zZ."G@t���
�з�MyGn7R:���;�<V7���P�e���{��#�S	��LԼ�����g��d�yp3��g��h����v
Q��=�w���T��#,��"��
c+�VQ����|"�+���ٵ�+<u�&�Y3,�a(`��<����n���]��9�<͢�P<�!�)��o;q�q��t�8㏎8㍸�8ێ8㍾8�:|q�q���8�8���q�qǎ1�q�>8�8��q�q�x��8�8��q�t�q�}pqǎ8��8�n8�8��8ێ8㍸�8��8��q�\q���[�6`��Jx��fL��a��J��K2�v����|��5��M��1;Y<�oX�w��ԉsR�+7�+KF��:��C�m���&���/��T��z�"Ӥ�e1�ُ^�7]]0x�g��7��f�/��}[V)Vf+j���.��-����)H�c�E��Gn"k�:�D�W:�9�����V�g+$��-RW�ڡs�:�P��G����[�L3�}HnLXl�t��ዱ����Py\;6�M�x�o^�r��^Y�\9�ƪ�W��t���5����Ҍ���z��DF�z�ooKl�@�c���5�&���c�WJ�N\�%K��B�D%F�ԏ#���ܝST�]���Q�Oss2�WB�z�f�s�7���av���Zݱ�cS=���YR+�t�(���M��6@h�nݺ��lnš ��c�����d�b��e ��x�^�k��9��zө����m�˃(��Y��N�o�+���0��Q�(��=}aWb�g3��V�V�U0ͤEgV!���лJ618(����Z�r[v�]^�/��]2W.HU(�|R�����+&��VY}��iֺ�|�ZEwV/��!w_CS�;t�2�!��EU���7����������8�8�q�q�q�q�q�\q�N8�8��8ێ8�q�}q�c�8�8���8������㏎8㍸�8�8��q�8�8�q�q��q�c�8�8��q�q�v�88�8��8��q�q�q�q�M�ֵ�w�����g50%��m��.Z���aI�����xmwf�4�}��w/ �������+� ������HPg��71-�Y�.ع��.ږ2��p=Ъ1G��F���m���c&w��Ez
��XҼ���s3J������ɰ��`�ݴ7������*Y�1ٷgr��h'b�6x62AɍOgfb�,#ǐ0��s(>�h�/�+mf�+�J]��qw���f�<���V�VaJ�ĩ�u4V82�}E�h�y��:w\��hT�E�b�� ��`�e��%����F�������{Hd=�I�3��<c'8�=dbz��m�h��JFNb��]�,��e��.����d���s˺C��T���HA�ٺ\3D�;��v�)�X��r�^Xgqo,5�\��S_�K`���b���Ef [)��tv�ڲRYZ.4��[��e����Zƒ�{��r
����֥:M�L*�4:���l`Eۤ3��<���a��j�����AC�$�|/��>v���뜳�6lL[+MY��p3�L!~;~܎ٜ�9���A�����h�\ѻ%nD���#��ao��j��Ƅ���S7�����8��q�\q�q�q��q�qǎ1�q�qێ4�8�n8�>8�8ێ8㏎8�6㏣�����8��q�q�q�q�m�q��q�q��t�4�8�;pq�q�q�q�q�pq�q�\q�N8㏎>8�������'�
LS_;5[���_��Ø������s���W	�9����gb�T2�.��"2�+.H�me-W�K�&�D.]��K���_>�;*�G�\�j�k^�Z�(�[n�7��O�s8�Һ�K͘=�{̮]6&��n��V��7��0|�{��\�H�L|S���Xr"I�Vn�h�)�f^����0e�B�v�{ώ�7����Wn�N�ۛx��
U���z�XUoCr�]��2Q#�^u��Owf�T���M�F���fg��y�7���ɰS[t9�ei���߽4�&�m{a[���J�r�U����+;G.\�]��t�/r��-d��Ǐy+��q��y�Û	n$`t+C[�ء���:R���^� !ƀ��)vce��.�	�F]�����O �k.��V��4��Vc's,��b&���p��Χt���y���ugU����Z���8L��x���l0���0�2"�~�(9�-bh���'�huE��7��ofi(�\D�*����t�1L�o��Ỽ.�zԨS�t)T"]���ِ�{�F�@�)�:hn���\��F`�NF͡�ӣ5�xk$���D�+E).��W*=4�Q:
��B�͠��+����*jG���Y2��6L�*�{�Q���1+�����:GR	��Z��ڛu��]C6�7�����������{=��q��t�>8��qƜq�q�n8�8�8��8�8��q�q�\q�N8�8����___\q�88�8㏮8�q�|q�m�i�q�q�q�8�8��8ӎ8�8��i�q�v�q�q�q�w����{��G�R�F����y�����v���6�&�mZLQL+���\ihe-��c46}��-���]+i�I��u��%m]���C�T����T�8��Q�t���BV�^�s�Tl�s�e"졯A���g\٧*�,�\@{ն�RD7T;:V�ym֑�8�u��t:$z���m��Y��6]�T��uF���L�N�*P��ʑ�	,�J+��f�:1Y��te+B������=I���.��l�q0�n�Zޣ��4�5�#еl�l�����-i��t��=x�ΔÂ�BU4Zv ��8�+ٗ�"�2mr�Nɜ=u����Hi�Q�V��;���i��Lu�	E���VV .�=����Ces�����6���D+�U��6�kR���Q���!��S��(��7Ԋ�QZ���u���8�Ds���U�a��)��K�G��H2�6�>��d�J�M;�#��+jv��x��62�1S:�=�&ݺ�W�8�ږ�a$S��9��w�j易F���G���Оa��WQ�;�+.��qQ�RT�I%z�e�f���Y�b=u
W�]XV������&KF�sޘh[X�᫣�]=59u%m�Y�.n�/�N�RP�]T�n��fr�}i�V�A-%f��U!
 %:󮳱��fC�;��tt�����7o2�mQK9Ī�f��\Pi�dd��t9\ͩ^�N��%s�5���i������&5-g\���>G��*'�i(Ň��t�r,U۴4b
(A�>rGo��2�ф;.W�	��Yz�᚝��IJ�0�l#���TU�������>'�^���,��+�P���G�;�\����bemd��uxa��j.�޶��(����e���Dmje�D�ⷁC��O3�W��!Q�Q"	��&�+��Uݦηx������HU�\�tM�� ��|�`W�Z���<����4����oD|e��1GB����E�d����@N[2tS�(�����Ս��	d��0�ze�����x�58@�OfwR։�<l.�tT��N�{x%hT-��"�v��13u�GK�"�x"X�d B��8�_fl鵶�F�}Q ���"U������<d%h����%���#ׂu�����b�ݽP�ls����&�v/�V.R�F]oI�(�h��/+#{N[���^�Fqi�ϒ廙��N��W:�z��/�J,X�����IR�S7��}�T��wY��Nh�3�o�ᗃpQ�ۄ�Տ^.����<�����h>���;hn���t�q��G.뫋��C6��^qM�#�+O���,�n	*�3P�O����S�K�G��9/�VU7hw)	�y�
�e᱙�J�fCܹ �bA��er���VIë�n����^eѝ��;�T]�צ�e2^CJ�r��;���f���;{1�����J���f�G[1�t�r�_<y�wZW�]yq�[ee�L��Z��O��RLR���q�ldXU�-7^t':+�8�l�Z�Eк*�YZ{m�Wn��}��z-�����]�t��/v3�z�Q�=M`��}���Y�lQC�Z*zp��=z�L45I��:ۭ�K;Y9v��eT7��L��O���t�Dvv5g��WI�`�y۠m`
�{��ʥ���r���3��i��ݫA���l���ɡ�;-+�('�r<8��c"$�Ѕ���*-�Ut_gX�t��b;�Bw�j&�V��z�Џ.͝�%
WYrRdPRΚ~�e����u%Va�n2R��ѫS���k2�5&*S0Z�[S�*��Y��7�hxcnaT-��7}��r�����H��̼�gM���'HK7UI'bAӳ��������f*�%xQé���vL�t��v�:vz��xGvرw/�9X��r���J���YL�("�{�i�&�������r�5
N���m�[�էI�.a��3�ZcۖS;�9Gۧ�K�=W�E�1�Gh���c���7����.Y�ڣn��C��N{����܇�&K/'�Uթw�%�Ü{u�ɺ�ҭն�%�n����3��|6G��T����G��X��4�����u�]Q�;�l��cKX��u�J0�(E�K�s�֥���g:�muC:0�=�%;C&uU�����QӍ_��XB�s�4�y����ӎՈ���s.^un\�Fnrp�����/��۾8uzwN�wu<�����UWj�I���P�:�ۤ�dǹB�%���v%�=�� H�����(��#7�֑�aً��U�d�'�����$:{��6���PS
KB�Ԭ���v�V+a���=X�KYR�d�;V��̢n΍���}tg^k*���25͎�L�1I�{����y�ev={|�OE��P���(��-�9��ۧ�՛D[�����;])ja�U��2�����)s}/Jk�28�z,Y��'�vS��._8�i��]\D��vR+ᾩK�W��ս���pQY
+�t8�R��U�rlWy����A�+UU�I+q�4��-�w�*�.��z�aےЋ�٨��9��t���ݫӜ0g4���)���U��N����Ջ��r#n���{l۱f�"���N�ǽz�Sf��� ��Rq���g��H+"���^����Bn󺷒�Sy�M]ˠ��W6m�N����%����PJ��U
��F2�ټ���̬�3e�&wJ�T�.�A�k}������`�X�QZ�۝۹ǗY)�M�Gs�
�h`Ma������U�g�������ZNG����4T�n�.>�Ҟv�W��oS�HgS����Fo"�	P�q_C��k��;�o�Z�W�.������|t���O!F�ݕ����N˙g�9��]�&:�{�y�H�xN_�8QV��v)ѳ&n�W�:�m���$>�U�z�\�N�$r��G�u�8�f��NH����cUBx���|De�a�x�m�2㷂�V`d����sx���XI��������x%<on��������- �*	R�+��e�4qq�e��F��9���	��d�ٔ�����+��k`��ݲ�0��eX+$���)��{[�na�;��.����b���s�h��Z	��U�gS|o���X.�Jq�&_���B����|�;vۓ8t��.�ն�)A�h�=Wi��m"�R��˻BF7h%��SG��I�#!�s��WM�j��yJ��+��WG�-[.��!�v�����f�>Xp$k���ˮ��{�@���Y.��"R�6D�wG"��Yq>\ܐ㞩��T��][�8L����l=So�b�$�� ���/C�(&c�C������B�F�r˾��QV���.z��*�2j�3K�`��
Q�3kB���%u(y�A\�����/rU�V��P���}�:������\wn�GR�0\�a�J����.K��s[��T�w�A���ޮ�c���]�XQݢ_Y���\z���yɸ�!�T�<ۊ�e�p,���ԩ�oۦo`�rZqm	R5����t�wM���7}�������f�{L���>x��cm�tqˬG7�ۭ��1[ڻ��()RF^��h����u'����!�	��i�:f�G�S�>�uϲ��׃q�0,�S�X��vA�l���h�U���	�}c��V&���M�_i�G����9��Ɖzpe���oϊ[ip fT�����s!�rBQN[|�;H�u!`��[�A�x�2k]���6��6��=�Y�2v�x�h)�K�-8]ѼM!b�.�EDfӡV&�5dF:vD[(k�dk���q^�Mk�EM]�����,GxI�������3W�W������xBA����$�D"�e���?��}� ���/�_�����?�~���� H������+��!��{��?�aDArM�e&Z��$���"6�DZ�ŉ��ҷ^�=V�Ȕ�E�(Z	��C��5���p*Ԣ��j�:T�)S����b�u��x���`��W�`N��<2��Uْg!O�c����<���-��D�j���\�'܍�ͱ���/r�	yS����}+x���Zƅk���]]Lڌ�u����S�
j��T�*�ҋ�9�v�7�>s\S�v�뼛�7�,{��=����|�:����V���s���Vö&��t����B��=��Q�i��+y�,e�fk��gj���@�;��!����m�(�2
(��`
w��d̘��f�2z��y��3z N'u�	�`�(�j�ٹ�8�;wqkv�c�;�h�i�D,���J��h�)d�S�V��Rǆ�vh�e\�N{Z,�/^��A�|�
�yBƠ�X�~�AU�t�M�n7��nON��RT�i�/i^R�t1��-VT�y�%����z:�Y�3���Mӏ:ڭ��^���̮׺�6�Kyx��7�]�;�3:������;�nk�W׉W2���b�u����K��F�<�reb\��n\��2L/@�}�5�M���̼�e��I^�bA���0x3���Q�	�n�p���{�nu
ȩ��='��P�ZȲ��B�#l3(��D�a��p�^d ѧ�n#�a���(�"E������j� �O�J � �0&�XEKur�ֹI8ZUTp�3]˛M�C�㎟ϟ>>{�{��}���d�w#�䂃� �H�|ݸ����ȅ$rN>:||v��nݻv�xfB�J*�Yfd��8""w$	4�!�	QB*PB,�q�}q۷nݻy����ߟ��$�#������p�r _�����
B����A(d�1��q���v�۷��i�N��L�f�R�le�h�u.m�K{�����KZ6L���bƘrC���nmv�>����$;����;����u���U#N���z��۷nݻ}z��v?Y۵�wW�w�뷶����E�=�z��mqݖ\���#���],��g<c;�-m�aݝ��vure�#��Y�Z�wu��7af�'��8Bٳ+����L��16�5�{�쮽y�gi;�m��kfcZfλ/k��ZnT��y����{�~7����n��ݛn37RΝ���t���y�:�pw�k�ٷI/o{jk7�i�׺����q��e�h�K����DixF�I%۹gpVM��s�oi��u^�Zޕ�ye�w��gq�W�n��l����N��Ò�m�kC���mZ:Q8uy��%��޶o�|w�A���I~{{���Ȓ.8�i_�}��}��}���Z�I�n_έ>,�'�Ȋh-�5�۷�z�i�6u��p�x��N�^�Q��'Dlv$ΰ�n�\�F��Jsf��LEu��o�Me�>~8��*:)ϐ5(�@tL������Ќ�Q�ۗ���Wg%���Ms�f�����R�����b1݃��6m�W��ԍ2����p�U��� ʋj�[(�֕.D2���\��S�C�Uǭ�^4��Ҳ��������|�Z��I��,�1T�g�����b��ޑ��!W���������l�Lkj�T�R��/vVjRel�T�g�ն�^��TޖY�[��J[`��I�4�^�����y'Դ�Fײ�N�4,�)dǘg�qb�$C�h�^��L�4��S�i�}��8�~m�o�vj�������� ~�R���eL�(�,/�n�W��;l�5*k"ƙ�}]�}� �E|+.�}�=aDO�>XQ3�=fU�B�@�V�(����8 ��~�0��B��hY�Ϧ���t��K�K���#�1˜���f��PneC=�u�p��؎�닲dX��<>V������cV��Xm°����r?ڵ]s�wSF�m�./�t��p7�&z�C�{�y�2%!�ϳ
\1ں��d��Wg+�l�����s����y���A�B�G������y����"m�d�MWtq��B#L+�
�S�pN솶kk���/Im���^Ycc^"�c�X*��$�����wr>�Mn#��P	�qr���}T&弱��mS��Ag�ND�2<I�3�s]z�x�r��[��)7sh�Ǻ5���X�JUj�>�*gf�X�!HJ��}I-iݼgc)
��I�QD���!k,��6Y��
�U=D*FE-!M('�[�iY��)(l]���΍gƦb��(�D����#����j=B*�V��F9"�N�B�O�`1)6�e͔ިEz�*�i��Vĵ�}���xg���N����<�rc]a�OM�7�U�:�UA��n�N�;5.�Z��Ai�&�Zm�d�ɶ��J.��y)n��{{XDC�Xܝ֮�s�s�\�荄��6��h0~t��Y��Z�P\:�<��L����&v��ӷFڌY"�34,��ژ4��� �_�c�I��s��oe�}��:"M��p�>a�AQ�n�!R'V�bw��;2�g5Z/0r��0.o��ކ���EU����m�f�|�4��q�� cbjqc��`�QI���o*�Z�f�5?�d6��O�c&�L֭y�.�;��Ӝنa�Ҋ�9��}R��nzQڣb�C����33���[�l4����W[ ���H�sךۯ��1տd+��tg�6!�s����O�����x�[��ʙ��ݪW4P)"Vr�u�|w��;���s��X���gз<�;ǳ}D؍.^5&V��gS��uD�ՠ�-��@�6L��c��Pd��m������r��[C$����T�f�����p�Tc�PA�g��շNi>Ú�Yg1S�%��f���
h<*��J��Rb@�FBHG�&�l�����)qyv��z5��_���R���rj* L�ou�9t��Qbٶӻ�h���5� U�첽�S�^������0Խ��,S{������Z��vuf`N���%w�}�2���.|ᖷ�[���b^�~]��v������Yq�S��	�q��e�
�=q�C����,��b���a���ʾUl��0k�{���7�jCt%���:�����oBU��gy�kGnw��4oy\Kq����}��
�9�}K�m6�2��r�l4���@c�U^�FB�)�����ƭ��l��9t��8)�UKl����}�aQf*��n�ׄ����W븋˗M������a�SV���^ݐ�	6+j/JG)�U�&R��5
�j�(��6oN��Վa����s�w[b���
��Ze"��\f�k�H)��U��
��M�a�i�N���7f�b����HI��Ywe�a<+ݏ\/FQ�:aE%c�g�k��6yk�AR5F��	��6�JKIS��QHϩ�{0Y,�^I�ǾJt�l��&~}�;��ե�u^����i��+&�t,������o�r����ᥜ�ԯ�UO_���\0d�ET�Kt���i���΢�n/��V�&#/�Gv�O~Oub�+�|�/&�����,1X+)Ԡ�ʋ��Q�{���xu�ˏ�f����
���f�<��'�Xt�n\��'���Xw�w#}P����r�nҽ��+;��Q���V��q㋶�:ɝ��藎��f�ކ&UA$�t2�*�'E�y�ou;��U�%i��e�;=ָ+*����E�`�l����M��S�Z͊�fs��n� ��w�*��H��MK�m�T1�/xe$�<(Xf��p#�K4���Tm�(���IH���tp��ee�hk�Ņ2�4���!^��%o)Š����>��n!��45�I�	�*�f�db�����mh�a�>�ܯ��)��4�ӗ�O��(�ǹ��f�5r�:�{�Q2&./4*̿$VT��p�R��a��ʱZB��B����TF<�q*��̈́���g�"en=�a��uKR�/rƪ�M3���s	V�b��B$kͽ�f�]�g��W φg<��?��Ւ��^��+@;)$�ڽk|�o�^x��NG�EǑIJ��Ɩ|v2t֧���K)�;D�*��&|�vNٖ�.N�C��\b�L׋;Z�>Cf[<��S�<���|l��'��ߕ�z�Q�۲�T���0��Q5��1�UKw��'e���H�c�1xhI���qoYN�iё�	�Ի��s�
 ���}�_�n��=r�w,ֈ�c�PN�E'*v�T)݋��z��=e#>����"�ۋ�*S��g�K��C��y�l�!�-�V6-mW�o3T=P�A�
BU���f��=W���S�LW����xej�oz�$s��Gʛ��m����Lͻ����K(>��Jp�q�h�'�5Ӫ-���P��k�,10�����h|T��8�F͉{H�Q
*�߮�r��v����?~��&�>���,5�s�N����S�2�t���� k$���Co�j��������6���B��sz���7��f��u=�98q��{��:F���D_�S���K^.�r��)X�^x�&�r�jr$f�.Bp�ܨL����v�������Ͼ�r]�\�"�6���v؀,�U���+)+g�%�.�i�`!I�q��l�6���g���{�TL�e�*�(,�/����Y�c�Y��>����
�]�ܠ��t���육j���[u���`+Y�XI�Ӵ]���1���]�ܡ()t;p��q�	,��S7�_sճ$�v#�D�7C�i�^iI;�%+jC���MUѴ�3�EWs�l����cB���g��d�غ��_z������U4"�Ϋ_�a�;G]�۴�|*�˔^��N�.V�0̬���D�<��CT�
4�ؤsZm)G��>���x�4؎k�T
�>H��ˍ�u#HC�r�ٻ+z�I�ϳC�H8���+G�d��F�^rRݐ;���e3�]��>����3WG'�ڏ3�d4X#z����{�O�ioʾ����٩��:��p��A;�Y4ίRl�����ly�e)w-�5X���/�a���p�:�Q���LY�X+\�_q�;<K���_T�3�1�̑�*��W�����3s���2�͇<���ͪMNM]HOzs����E}B:��קL׹a������PU�f`:ђ�<N6��W(�I��D!mm��pl���s�c�d�4���n�?/���T?V��hV����!e>>`؝շ�{	)׬�S��{�Kܱ�ě��/{fD]�2�וd䂬��u�Xh����Q��H9���.��f�$Y��/�֝�c�\����T�H����r���&�N��5���z��)���^�f4�m��!���h����m��@��[cK86'd����,������"�%��d����o:Y�aMwM����o=��.���ξ��ж?�b�H���x��E�������?h,��eH��D�e�CIz4�̌�������ލ�>�a���!�R���nѫ��U�f�2	t#2�3AT���i ��D�����)��L�BL^i]��e��P�
����f"�[fA˹٧�k���hH�*���T�f�ҟL�[hX���tIl�-�J�N
���/35�*��қI
&p��\�Z���!D戬^AFƹKZ4�`�l]o5�i����~���߁ȶ��$
8~z�k?py���[Μ�
2ebg�5g*k�ͪζI���P����B�h[0�
/�V����#�	*�f�F�RX!��-T<Ӗ1�p�W|_<�q��4+uv��[�X���Wdx�n�$R���qfV,X�ge��_s�����0wA˨�]�kus��sy��xu�z4�"�=�j'����s�r���U�Z��!ɶ
TCD�7$�n: y7��n��v�z���QX�(�4
&B�����mϞ�3f
��!"�4��dн/�
�<jǽB���V�f�10y����x�2��D\6S���6T�*�G��9��n���!�L�N��Q5Jv<��ٲ�m���N*�FN,F�M���mÅ����K5�(錗�x�]L,�:䍃��9����5�_��W�U��d�ض0����@rj]S�35��{��EE�QgŶ���m2�f�^�,�©4��|�A����3�Tt�J	o:�ž�1�F�g�,�V�9h�!-I��;-U��(;��p�ޫ��ը��Y'�"D
�Rb�CP���`R�w"-��,O*W��jB�<P)ϔנAKY�?������䟦�cGN_Q�ޜum��ә���hN0-^��)���Р�V���}��}��n��l�M[!��c�:����dJ��AT��/w�E8Ny���o=������x�-ONV�z�6��}KD�[j�I0!�]��B�P	v�SU�����	Vڜ�9��m��V��!YV���eL����ʋ��+5}���*Ν��F�Z���˛r.�'��:6�E@r�"�O���2�F՘VLhѝO�]&�Yئ�g��P	e=sZIM�r!(�"(�IM��o4�}A���ŏb��H�l���t���{u>���c/0���ra��"^�f_�[E���(�%-y2j�F��k�ՁR�y��J�V�*�P�W��ة�M[�,�e?�$�%x�R�4�̬�u@����OVo���L3 ��<�Dm{/	�y����Яu2y���ݪ���h<�.���3�R�8`sg���y�6@�+(I��Nɛ���!��#U�О�,+)5�<Fߍ!~*��`͞�U�2�����U�<v�>����p�ɕ��C�!�6�y�����{"�}z��h��䎷Or=ھ�x�l����!�vr6�;��� ��?d,ȑ����굵��J�>���V63Zj�G�6���,�yk�
�:��ջ#&b�����h�&���_M���HDyO<�*�y�f�������ua��_%%)�ъ-}BN[���c:���ە��|H��EmF_��j${���۷)M�4+��v3o���ܫN�l���U�
�<�"�u١ƹ�ި[�a�d[Ÿ��W�;��#O8�MR���=�HA�Y
��'=�]�%�Y��+���enP7�f=;ѻY<��� ��^Լ<�n��f#gsV����e�gVA%�i>4��4���=��%����,�S���R�����}{�V?�}�ܕ�� �,a�	�w#jŠ�Ǖ���mN�o�\J��`}��v�Y��F^!u(�ۋ���]��JP-|�f0���9:K�ۙқ��d���t��J�4p�O�g�ٺ�%�<�!�F_+�R؜t�n�&r��!��qsћ�p�p���&y>ьN.��S�.��n�:�����U��7�%�G���kp���eڔ�5������4h�0Wn�6�Y	�:�M�B�XL������xqR�G���)���(��L�x��͝5�T�k.t�!�M�E�ؠ�t����0�7��_^�a�Y�7������ww�lф�M$�#�i"�}M�Н*�ع��G0\�2`�^T A�
�����ov3�a.�6����J,��Lޣ�ʣ���&�4�oE+�:���#ެ��A�ѽ�`׬q�X@qrK����-s�Kb���m�}Qr��vET����3�1��}3:�0c�*\�;&X�&/�>�au�]�xf̨�<�B����oX؉�g5t�,C"]����2�����f˘��e�e��[l1�5�9p')��#��F�-s�h<nv��լ:�>���W�xv7_�n/ gn�W���I����{�Gs��6r���t�#+����'�r���y9���=�Ȏj���2��qR
���{;���o*^oK�h=x�=���L��2��t�*�t�8��B�1slR��A}(AJ���sUWCw��W~�0F��ښ2s�+(�P��Vή�o�%l[{m��%5�t_v��4��'r&�T�2xa�CsJ�ZM��`�Ǡ�E�v:8QBcV��r'8���[���}W%�K1�)ݪ����7���Od��߮�Pܣ�J�eA��
vr���|p2]Y�ꡛ�-)���E��t�t�i5�7�Z���N�Z��"�oU#�]#����G��o�xS���;�>.�{%1Y��}3��$���N��cΑ��m��r,{�P�{[P�^Vb��q�Qu�SN�͡�����wh2��~�r�'I�{��	�9��Q[m�~��~7ň��k���FT�)��ׯ^;v��Ǐ�zǧd�P*MI
a I%WX�A�OkK��ސn��^|VE�v]dqrI#|m�v�۷nݻz��=N��g(���d'��&�l��c���]����I�\Ԑ���]�z�۷nݻv��~���GZ��V��� �~o=),��˃�$	�kTU2I!>�z���׏�v�۷�0��$d$r�XI)� );�O�����)�V@�Cn�^qe�%�n�M�Y�q�D�wf\���	�\[n���[�ךd�%���iE%�Qfrq|o#,�BGg��^6���~l��+H�:Z��S������MZ�vN�e�r�h�mĝ�G!gׯ�:|�\eey^^T�dGHwHVua�u	������2��V{�[�:u̳�lNp�t��������a�PX�z��(�)��E�뵥��2�Wp3)$W����)>��|��I�z�1�bq;Y�Ν�s:��qT�z\eՒ�6�O�Z�k�����HIT0����0��/��Q��U�HVa�e�fJ���<�xa�9�=xKոג<⮍xMn�a<�|�f�ǅ	ȴ��;��.�3gD���5p���$PI/�eXX@f}����:�[��/����1�.*� �C�n�&;[[��-��Uy:��p�M����t��E�(���F����,.�:y�&�1�����(O5���h0ɸ�
�����6����.����
H�ߜ_�c�=���4�)$��� 
��"����ge����g;+��
p5��Q5�`	e�k�i���U�~���}�>� .YJҿG�'��|�c/��j��7Y�d->�[[xE��£1�D_����DJ~��E0
�w+��sq��Ƹ~�w����3�b>,Y�b�m��-цD4�����5&@�f��ܾK�v�)�Ž�e�ɻ�_zr�ۺxxO�����x��zԇ�� �@�@���R+c���/`�CМ*��u�5��)�O,�l�y�aPܷ���y(h�]��Lp�x���Ô�a�ֺ5�$Vt��ڞ��*��*/:��j�عm# ��+�c�M��V;�u�-��n�C���Y����ڃ>aZ��֛�[����Wb�9F8i;�����Ȥ�p��E��F�kPy���I��ztٍǇ�dwD�D�Qr����5:�ܷC��z0#0+3/��j��^e%��|=޾|S���߄BiV�ؽ��kZ����<\�g=�ۨ�*&j{� ��oX�S.500[��iO�ө�]�m����V|4�M_6�n1g���7U�Wh@����Y("Rd�k}+�Xń����}��z�`i�㞯i��D���� "�Yы7IG�����=�sԻ'&Ԍ��\���BoG��QiN[�ɓPw�5�؂ de����w���x{H�^~6R��Û}�{A��?�\f�S�EC�iC��q�����N*>V8 5���ڨ���CP8/X�z`8y�H�.�c�WJ��͐;�,���'r��Y� ��³���yO�Y�Yʹ�O��%�DhT|�=�Ȧ=.M����N�1{d��҂��:���rnn�n�`�W Q��(�Z@��|��%fr���{�;�>���ls*�"Tʗ�;�WyK��6�G��<�cY��=v@�Sݲ?=��MC_b�~�b��w�<�z��T��K�;>��`60J˶�����#g��#��4cu�Sx�W�FX��B��E�H9���'��[�jÏ.H?U�C9�V��Ӥ�jk��2,j���N��>����@��M���$�H�44�/C�R9�q��,޽�{GR0��Cv9�v�j�׽�]t�w##jb�f,�m9F�.�:�2Υ�֧�����Sh(@2�)Ȕ��o��������(K$I���o8ɩ*S>,���> Y_��=w 
�!��^%|l�@q�1bO�w��:C����^A�U�o����xo;&��Q|o8
�}�r�:�]�XHN���Q�:Kq��7&�l���I�^ ape�f��7�>���Xw�p!���X�D��\
��s@Lx!�6���zʠ���r�0Z������`�i�)�:���}�Z@�6�3v��p�������_/��@L.�#�u���J�o,�:%���)�)?�r9�P��^
�s��B`�p�Xs;��[� ;��q����i�}]�>���6���WL�,a���I�(�M�����n�p�G*8cT�^A}�yc�޼ɺ�O��
>��
�a{>Z}R������qAԗQ�E�uؙ����.�M�>:���o$������^��x 1��ަX��|��`�@Xh��z|8ح�S�r��2j����-껆=c�P
� �1G�� �Ʃ}��PG�0.!�T"~��������6ZΧŹ��zż���w�<	x��޼�ߒ���[^f�V.���p%�;�@�����j9Q��Q���븎�WS����[BQJ��,to�;�ۼ��\fS��f}���o5����]�f����H���ѼE'k1*���{&�e�7: {�<�[�d�ޜzĜ+2�M�;
���C#��qN7�5��Ms�_Zy��k��+����{���������������up�	��[�G�2|~H|���}a���	9L����x=�o0�ƁB&�)��ݧ{�����S�G�}F�V���v��~��Ƭ����a��1
|t֎�<���!�y���+}���A��< �.:2����8*a����F6�C%w#RR�l��o��sՐ���F϶�2o�����ı��k�ch|x�h=Q�
1�p=~��������H��^�v37t�{�]}gj� =�n|8o;�4��2@���A�GexA���_��:����W*8�04���V��?L���>Q�8x"ꞛ��,9��˫��"��>����1J�~�/
,r�ׇr�Z�>�u�!M�l[�[D�S�C闖�����)�3G��e-����ފo_�P��x��~@���� �?
���� �F���)J�O�{��z�|�/R���Es�xOLqu�/�*� P5i�n/����@I ���"pN��GfokQ��
�?s���l���k���w�JL8=s�\�yk�}n��Qn�{���Q����O{��%��z=|v��|�h�ɇ�a����xU��Cо�`Z���X��E�]]yUMY�4~���5г;�~�����]��+��c���-���k駗-��ܕ�L��فE�����=���u53���G{j�wr����p��gl���,撧�W9�k�!o�U��J�����4�4�SM
B�H5y��9}�|���K�-��<>k�.��ySFO���[�6Qf�q�U�9S_�d�Ua��}�x^��u+�S��l^ $��c���>��O��]��8U�W:>ID��F?ߺ�m�xj1�=�1��ґ�Ǣ��һ�����;$ᘠc���#��&�F�7�<��d�/ve_k�������z����j�~Z�2c47 �ݡ2�#��@1�i�z>d4zlp�곷Tf��HH|<�
�C���5ʄ+?m��Gϖf�CNm�R{4 �(B����1�����K��8]�`;9<s	�~�xɟ�0�\||h5ǾS�@M)����NȌ���B�D�%ʬ�ƨ��gEl���$O�|5M�@�
]�N�$1ß�CN�}B���$��"kXѫ���f���7]9y?78{�_�������3H�j�XW����v�ޯP]�<���ܨ���=~�2An�3\�hޗИp aB5���@ ��~ׄ�{ Y��| &��H�p�*=4A�%�;�^��S�q���k��2x 1�L
�L�t��5<0ιD��<�T9�25Er�T��>gǮ�GGS���>���%۝�6�G��$�[ֆ�J�@��˘�묹-n��)C~�M��g�f�>�ό�HF��g(�+ʋ'+��Ek�S�]���O0��3!�sq����ڃ+f�����w۷:U�s������>�/ ����i��dRA �o���&���˧y�]0��<�*;A�q<����<�at�S*ʻY��x["���H�
�}at���VRj�<o<y��A�5�� 5`�K���cR���\B�
#�t��([yP�x�`[��d�ہ�F��c�n��}�7��K�@^]�o(�y��2�9�P��>k�,�@i�~u��yz��N��y�/������0�y��Ѽ�5�@6)�	@t�Ĭ�1C�#���p�
i�>�1�H����9����/q�Di�{��^:�|4�RߣuP���_Cq�����oHp���S>���5�YX�&��o
����K�w������@p�S���{��Dk�z��|2��(Z ��a��j#^j'1U)��'8�9�{��o:�%�����,cYc�a&3�S��%ǭQgfa0ƌ ��%���ރ�r�l��{��AQ�?7B:���?emw?����0���r���JsN��' [�zS��֙/ ho;��$g�,�����"#�}~�᧲@��,ڡZ`	OEC�b$v��}��{��*F��N����w�M���l�#g�;��������Hjs���/����t#���Sp�v��dO��o�@���֧�4ګ��t���=*�b�G32V�djѹ����=�k0U��.9thrFڮ��.�PP	���OBXٓyB��Yש\��yK�ǣ]�w�ᔝj\ĵ�/�	˲�J����5��m	V ��� �}�'Ӓ*��Ȣs� G4Д�@%4�%4�!  ��'� Tt>罫��K���H����b���#���9
)3�j���xL��~T��؜��ΧS�4q�:�µI;��]� Ct���/b����ɯ�&�W���4�M�7����S��X�l1Aw#���6�ʻ��c}�B[���Mp����nù�8�s�~���3��>�8�nb�ֿ�2�Ƈ&\0��Q}����� ����5��g�>����z�z�����Gh��"L��8�3[잍9V�t�5t��ˇ����*)�O�����WHhb_|�����{tމ��]�;��5�""�{�ږ{��o�y��}FZ���7}8}B����~��P΃�;������(7C��ٽ���ʒg iqMY��+^�EP8�U��uJ�v������sږ>��g��E��#�gk}�{�٧�6@�5(�O-����p�-#Vė�p���Q|�ԝ�j���1�E�i=_X����$J��h���d1d�=��~K���Yɤ�Z���(�N��9k{OCJ��Xkb�v�ߥ�:�OH3fJB���>9,��"9Q��x3�tdڢ�&�ѵ)[�صCp:a�\F�����n*��G�\��x�⬔��cmS�9��W�%���7��uǝw�V<�J&��eY{���݌���#<t
ǩ���}�Om����i�Jo�<���&��R+���cz���r��B�4ЩM4 �M
� H #�y{�>w�|����Iaa�/��@c�ǦÞ���"�y���̺"���I�`ϝp�²���JQ�-���I�U�y9�k�=C��O�8�#��զC9@h����8�w@ߍ{"m*��W���7L?E��A����8Ǘ��PM�@%0��0��[/�6R�<�J&�����r��p���������f3Ԣ�P��C�`�f���P���1�_��TDd��vs���!h��p��>�Ʈ*�/ �Pi(˴��-�k�<1��>��
�t�Wؾ599�V����z��C�{�����SSe\��{=w\�9*�M�S�P�(�˧`����;9[68���i-���<L���`�����9��p	�L��SX܂��,�����g͌=j���s�e����<����1Pꁊg����]6È/$|�F7E{��z4�4֌n��q�)-mr�+7��O=�f�]<m����v�ĦhJ���z��`�$�y�d%=>��+c��q��3~��,���ƻwx{���%?wG7�7z��ӳ���r^�+�+I�B���+j��T{��� ���"g�g��\{	fc,w��������]��X���eI�e�!�.{/��;��1�h�wtk"�S�c9ӛ���W�
=�f���؃���[����U͡���<��s�y�靧N����̈́A�c8WGv*�7��B-4ҠSM )M4���{��s$��>#�ч���6��W?&xnN���P�U�)�,�����k�	�ŧáu���vn��������x�,�;�ƚ�����w�eY�'�@�����@��|�:���P�[��Z�8c&�6=Є��m�`dO0�;��d��o�9�.�ʸʇ,V�*�*k��7�<�F����/�G@!i¤,(�\֑gEg}"�~���Ѭ���퓊񥽵[�j6Ǚ����q>����sl�S���,#}�ւ�[0᳢<!��d�+xɈnܫ]�,0�ep��5�ʭ}�aw������茌`�t\�!�K�R�n:36�C�הs��<1�F��1��t=�>�r����"K�gc#`3h.���͈���ؾ��=F�B�#�k|�7u������f�2�c�aAӒ4RQ�+���a�}y��G���b^1��r��[n�5�f��4��I��4>H�5�悭��E>�ؾ�m��y�<�G�Ƴ���@�|����w:����g��К��L$r����/ٕh��/p~Y����9C{�k;�Y��Tj)�!������t��|��AF�P�|V��θ��ȜO/H��@�>D/�_W�Cn`#�\�2\N7�;�>�R�	�hS�����N4X]���N�&v�����	�}�+���M%4ҁPE�4���BTI REIOkϝ�~I����=�����:�:��1j
c�ĉS��~�:�P����^�z�KO�k6���S��{S�k�6�5������Ǣ�=�%'�A
,P]��� s�>��۩S�c��\J��a��������{���$N5�2�&�xO��u�c1׬dZ�)P�d�����A��.��_oV��\�����
�5�b8'���(�\$sB��m񨽳�ȭ�d;L�#���G���O7���C�i�"�����5^�Jdb��~]Z��k���rCԴ�nِa]qN�M̝C�{c�,@Ʊ�$|�F�8�e;����G2��y���l|fꭵ���G❑��H近��t��!|�!��MB�����a������(��E�Z!uX�2�CS��@-�b-#il�\w���C;�Y��f�=L�͎d���Qo�e����۸Z;������I�D��5#~�G�*�hcb�4��G�|/ l������Q̠�=WwW���_��1�}���f�r����=�vY<�5�Q�	�rI�!=<<���������h+�Er~��ᖰ�V��&��u^p|�h��$�&�iӊ���\A�\o��x�e�Η�T�I�IW��`�e��W	�U{S���srMp��V^e���Dz䵠,�'��ʰ^��=NK�R���c��ջ�o�6���g���v��ؾx���� �C�-['���5��"�@�<���6s��[�w�������<j�T:!M�,R�ų����,����l+�U|�.���ը[�ev��MwЌ�i�b��������u�$ō�Z��:q^�Q�(E�.�M��.V�p�ޥ����� vf���&U�Z7��u�U�����x`]��� ��]��,��z��@�:D��sn���Uշ�+��76�J�+%��7e ;�_,ƚ3d�'�̡��,�op5Y��Z}��S;;�����"7C^ө�.�dB����W4����{ש�i:����6w��.��5U�>j����D�(�:�L�1��R���ZK4
:	R�>t�\ޗ�I�\���{t:)ݯ�˲��l㽜��K0��7�TyZhq��e1�Fc�L:9�]���{|���f�|��"NHA���@��fIyZɒ��O��.��9J�s�k�of�&WgbM�d���[��+%�1ʱ[��a�uƊ���-�$��A�S^�A�n5���3%��A��.�)��-�RLcd"iR\kB�-��"2���a��B3�S�3�g�>u�V��f���;Ĳ�%6�SQ�w)�)��𪭿������ti*,�VEa�Df�;�E���F+w���z�L^6u:�*.U.Bv�U����HW5Nu褦g$tI��{�-��-��`�ke��@]��ц�y|zPfr�C��(�Ŷ�bw����T�o'3��1��J��c ��'��q�*�<��ݍ�dd���9
M����p�1ףR�������EbT��m�GT��g����u�}l�Ul��c��5�H�r�'Y;��樊�6���eŵ����L����I���z�9r��Щ�	%tۍ�U��q��8l|H eΣMҳ��`���˄�K���a��,zi�u�M��;��Z�ݙk���7%��r�A���:�p�m�<�\�|����@gf�s�W	/ļ���]����Z#�Wǃ�K�+okn�v��kGv��hp��{e��Tc흐]���{c����a�=w�<��G%�T���ѭH��ަ�c##��t�Xc �9�9auԲ���ڌ�ɞ��y���G%tm��yu��g6�m�aީ��}���*�NѬ�O;Z8�)���:�Uɚ&�����P�ǌ�#�ף�+�;���#��|��F�ܲV��K^�$��L�x�Xn_^�'+��R`��A��fLjjK%���H-�(���bQ(Q5P
c�8�c��T� �]]�Z�[�^��$pzjhп{��i�Ϗ;���~�s�r$�.�����;��J��㔑!I$P� �ӧo^�x��ǎݻv�����I$aDI$�����Ipu$T"I!�qǯ^<x��ǎ޽����~w��qy�f�S�r[�x8Q��~w{PE�K��>GR1������o^<x��Ǐ��ߝ~N	�)N)��G8���G"�������SM��;z��Ǐ<z�{����nC��ƐGG�RQćY�y�N�#��0��yvGepe(8W��{�vGGqDY�m�m�Q_����r8���:9��!C�u��GAܑN�s㾕�W�w%��M7q��rtu������۳����v^Ϟ���zΈ�|՝|����H�:�����+U:2#D'J)�uۛ�/*%X3B���쨭�r�p��x���zխQ|'VPI�q���Y2%A�4L����+��:�`���T�x�1Ud�M"!����槐�ԩe����T
~4�Q�V A�B@$cM%EcM �@]���W>w�����p���_���^6e������=J-�	�u�������)��b�Cn^�8������[�^�|A�,=6c�q�5L;'ɵ#$v�~pl23L(��q)-ˏI����>3<�n�7�+=��A�l��v��L#�2ޞX���>�@m�b���9�>S=���*�5[]yʔ��,��h�v�TW@��v)阘\���η/����Cne�.w�	��qZ���^g��˲mj��'�x[��(< aqm��X�;	�d+՚�A�{ǅߦ�|Es����O�P�h�������CdY\�g̤��/^v9�5f�s�Uc�ԣ���v:��^�y��N��b����d	e]Ƶ�z
8���t���>���\r�CƸE|��1J���*��􎾑<�4�6z�T�Z}K�wj'o�?���l�Z�P�ܲCj"�� ��v�	TS�����G�O�>��)�iq�Y��.{;�j�1�w0ו�v�L���g���qd��/��ş1Qc�r����:������
�bJ�����Fw��i0��j��.��h�:�,�[���e�sc��^�s�n�s��y��c�1}{��hE,]ׂ��.u�A`�Unn�(F���k� ewL�ɷ��� �ekq�\�ƍӠ���~�i���F�Ji� �� (2 $��"����ڿ�|�/z�_~����^E'���
��Yz��d@�c���=�u���pe\i���W�eu���&��]j�$��~r{��C��`d��:���O�(�/��v�{p�'��r�/̧�dI�r��*�"����s�u�t�uC	����6$���~�������_�ڻ�&G1/b^K�(,�N.��L+��K)�� ������ˎ����1]�7�D�C��`��7�)�W1᭓jEu9��P(�k��I���d��ΡNn����;�Æ��j�{w��B<���lq���>~��,9��Yf%�W>,�p�r'c�Z�t`�́�z�v���ZB�	��=u>ٟ[�HР<
�yKhd���V��s���dN�]'k�V��zC����@��%�npg|t�ʋJ�a�W�'$;Ẫ��ǎ��[���p��;��m�8���oӿ8Xtp�}��^(�_l77�����<p�\Hp��^��[ϭ�ߋ�V�Oʠ!Ò�5�K�h��K;���`Jq�nj�Z�D]��Y�pP�tF�W�wW6Vi�{���b�_\
E�^�3@��4u�F�7�|w&D3���9{h��v����j�w�Ct�����Q۵���Z_9��ǚ�]��5{7�{�泓������UL���hA)���iP���2* �ͫ$�[Γ�����=�5�\���i=�qjE7o@��u�zPO7���mn�!Pή�3�]Y�޶�<��#�����J�!FhW�8�h=Q��e�U��@{�7�S3��v��3�P���vؿ��u�Q+��6YGE��$$܆ƿ������Wҩ�k~�=K��Z{Y�>7��<Ú��W��ER>����U$�!E��S�c�ҡ�R�^�]�͜��ʈa�\3�*=4F|E5;Q]�}�3��fO��wd���%UC�r�c����x����ݐ�0���3��o��Q��7S�\��2��@�4��WN��i;[�v��0�%%�C_��+���a�b�s��eI�LX�]Q.���7{�L�V؏���""�e��`a����O�Y���{�"xa����=#
��|*�]JRh�-����f���#f4�oA�5��a=��O��6�4b��o��c�:�9�>|=uYu��W1��iw�ث���~��O0�L@��Ddc>��-�CG�u�Y�N��*;�h� ��r���5��,j��Y�i�@♣'�K���}n�@�������SDА1��aG)��}���>����Z���'�Y�w��4`]�����4U*ޣ�1�M4�$ιhK��+L��C�5k/���(�^��}"�"�h)��
�i���A�3|�������K��{�㪎46��7�,,d��3W�\�LF�H�F���&vq�P��(,r��ՏݗW7���P����b�����@7b�>����W��M&�W���Lh;���N��f�g��W3�&�Oa�6�����9a@� �{��lw��sp���y�>�>��ܶ����B}3���V��	{���f�U|�0>~�3�j��%	�|��	�^]W���a��ܷ Ξ����Ik=I�;vzH�e��y���S�0>��[�_5�K%I��M���1���Q��v���|WW}K�a*�8�ݓ��7��R1QY�BT���y�ϱ�o!��񁭟P��kt�O��;�>}DO5ީ���;"S���f=zޭ�:���Uz�N�G�"����)�����؎/�a�1N6���jxn���=B;�<�ՙ�Er�H�I�����VGn�斣��~�8�Bi�8�r��#���Bǐ�9�{"S���E6&;������W�if]^�N���1���Q5�T#��/�ǩW������rR~�*L\�R�-$�ENc����𹳷�ӂAi-#{��f<+�_�~M�x	ːP�fl��I� ��G�f�K|�ޔ��q��q�ʇ%-m�%�G�W(����:&K����Q��%��dźK�<�������_k��iLw���1:���$�X5�h������ϡW�$~4���4�4ҫQcM	PE@�|<<	���0n���OvS���w�:!��d��NT|F�ϵ��|��<tC�1~0�È>:��v���K�ل_�e�a�xms�dQ�|Ъ��[!�6-?.f4ﯴ�ϱ��,�`�Q8O�0�t)ĳ�k��O����.����
���W�D���Z�̡�.�_��Ot�2���!�Vώx����f��'��ٺt�Y\�f̉/] @��ݞj��u�>�7���~���1hGk�PiV}�eh�Ȋ�"~[��a��:���#!�����ψ�p '2����w��uU��;�o�3짚`o#\%�A�A~�?��j���t%Y��pV�=������J���D��f݋�f��[�&~��	�+�(����K�{�R9���XPr�^���5���ZLb+z�[6��u�K�>�"yO*+�dI�f�-)�偩5��u�Ê�(9��{y+��H�����Bh=�]�84�2�砟9輜`�4��38З�W�����M���{�;�+����zf��[��/`���A����*��nN)������f^W0'���yOԧEX3���usz�>Y��y-����T�p2?K����tD������#Jc$�Y�s=����W��nX{ʸ>���i�7�K�v2F���ʞ��i�#�q)i��g�o�a�~re�9yg.Ϡ�(G�V�i
�H�ƚJi�J��� 5vv��O��}N�v�����Ͳ.��?u�YO�w�zP����څ�w3ѽdm�V��e����Hɞ��_�?�Xk��������;:�t�����*V�ܧ[�K
m��=�����&��|���r�O��%sfy�ǈ�%��t	��ceQ�b5��O{sdt��>�5Qq$@�t_O�,��=��$��xsB[�11�1�^�kX�C�$ֶ��M�Z���y0��z��L�lp՞�p����5��0�l����5僱�]��Xn{���I� ��ǳS��"u"c|�}���j�F�y8�Xa"q�p-�܆��_�o�=L$��a:,�/j���u�W��M*�9��7�F(B65_6y;�aq�=.�Xr[��?Je������A�	�Ɠ�����
��V�(	��YF��Fb���c��XC1���ƶH�'�}n�[��v;��.�^����hQ�g�ޛ��y8��Id��=y�h"<O	ZP7��F���Tib�l/�X�^P9�����4f�1j1�g&oC+��W��;hg5�5m\|6��0����u�8��,^�\,!}'��β���L�-�uM��K��Rqv`�W�����r���-V��R�by���Wu��/�&��P$ $��H�P#M"5�@)M4 5I@  9�i��go�|�X}@����-��S�^x}��;PР?Qg�(&����f�3�X������Mb�H���L3LJr��۔� �D��`[7�Db����&�57��M�ӗˣ>��k�<@|Bj��d�>8�.��̓�˾C��w�~�y��Y^{N*=_� �J����Ɲ����6ΈIĈ�Y�Տ!��\v���I��p�J��lSd���ڼ��6�<�EÃ�\�<*�����>!���B���P��6b���-�r>t��*ė��Χ18,���v �בdDT�kqAT>Q`P��y���^}ύ�^�񜳐e�z�u��|]H%�^���yYwgP�x��ۑoV��TQc�Ώ����^\��ժc���C�������J�D�����G}��A�9��J���J�r��;�ٴ�5���W]�Ã�޾���O�6g���@e�~ފeC�W0�6%��6������mڜ~�WgKUC�mzEИ,O��7[C��fJw��)g��a��W�u���P�4�O��%BpDa�n�4�#�8�&�4.d�_�>�?K¾̭�M����'q���y�;(\]W���WN�f�'��La�>��G;��C­�g �*����ѯB�K��S���9��}�3e^ø�[qir����NRu�g,�x�Ѿ���c��SM �4ТSM*�II {����s���j�]�?�HLs!����|8E�a;��D�k��l�0��*s��.��y��_^�y^�>�(W��\�C���KBد4h^����i�.�H�Y�@��_t��؛�O&b��S�B�>)+'~�W��o��n�lQ򔟶�O��`c����;W43>+�b��� �$]���x	ͤ>U��{���M��l�@�F׵�
a�[�ZM^�����+�Nr��=��7Sȣ�}��@�/�S��=8�T�Rۡ Ǣ�@z�ԎE�s��᫼�\ق�?h���̊�v�h���~aa����*�,ih�	�+Κ�na��q�N{��h��9RV�p��!�{L�ɜ=[휯�L����3��]�c��Ng�����.o����c�{W���>i�^B4p�-0���6�d�������Os�ȶ���S�	�P��0���#�Ra�Z�V5E&b�AifGØ4�����҇����k5�tNɊ� �TU��rh�ʑ��e]�lw,��3g9��]c`JLPB�|�����G�����v!�4�C+'J�\��\r��f.�E�\��!�ΣJE�̜�Ҝt��m_6�2O5�2���y�d��N�S��FU�Z��wNۜ����ww��|�gBC�U�N���
����ʌ�oe���mr���)�U�4�4<�5�9����[K�Z�R�K>�GO�B	M4"4�B4��TRAA�$|<����|����w�i+Ix{?�#6}Q�;�q�ϣ��֟�����,�qﭻO�"�'���Kʨ[ݦ�V��\0D�)T~�|Fu�o��+��"J��s�϶�|��U�	�κ��N�,��o��� H0 )�&��*���9��Z$
sk���������H�@Q����3WB���v�N4�c[:�2�5��_��
2��CZG��Ց�ƙ��w���۶�R�|[�y�$���i�h�<T��#�����l p�� ��w�M�U|
��@�]s2q\��^_tF�'��Q���	E���琚F�i�%����[xG�gd�s�&�T���o��4�3�����$L�Gjr+� q���������U>SH�cL��K"�����[(JaC�;�ם?L�N�`Kk��j��R�����@�C]%��F��l��^�ATc�go��(��6�"�^a`6GP_Z��/�L,9>�"���a���r��I�:�=�Үg��x�直��U��_���=+���T{�"�q_@��}����	��k��V�(DAڳY�T޵l�Ѣ���G��%�x]�i֛J���I�c0�0��hdx�����tj6���t/ OZ�!@����yJ̣[���(A��	k��pZ����7iz!0���W7�+�ټ!�&���k�����3��hh�ݛ�I>dK�[;��<��PJT����i������h j*��+"�H����s�s�����p�kָ�ʂA�e\`�(�`�o�|���v��AX�~��m��Nq�EƎ�o�k�~��~O`.�C�hsj}�����KM?�0�&'^��ٜ��Kտ�U�P��̎�Os��l|��W-.���+��`P%�o4��'"�sus�ɱ����9�f�x��K�*r�^���u�C�Hi��n.)��?h:�Y�e�b�l7�OT:=	`�;�T5T���"�-��(���Q�n>�����v����|�w��]����yˎي�L�
�~��𞚋��9]+.[�~�z�?M#yćl�,���z�@������g°&�/M�ޕE>��9��fr�CC���ēQ�C�WS'g����Y�ۏ~�y�K���#�>��
S�FR��;�g�H[�V���5�OU�6�vI��/�nxY�̃|+�@��̛�bn��Rz�*��q�z��L��}�|�ؖ\�������q =�}�����p�]���t��%=������sO�Nz(m�f��܁�ږ�w�՟/�u�v7s{��ߛ���M�۠��_s}P��"��5�w	b��4t�E�>��fk�|��t��˷!�/{$���nCzHzP�����ܪ�VqB���V�Z��X��s�5�{[��R�o�9v�1�{r@n*�:3E�T(S��Ü�W��9�Y�ٷ�e�2;��[i�J�NGw�k
�.�*FY��C6g>�������>�w�V_{��K�R"n�'����+}*ȮdK����x6Z�� ���XvN嫣+����y�x��׶��gi�/�v�|��FS1M �J��R+XV��t��ԩ���濆��k�:uUu��lK�yU��}Qz�wY�n��R;V�bW�q�0��
�b�\/�V�:���4��R�:>bJ}��J}0u,�V����[�vB��B���5#��+R��k�4����LޟFn���),vC�����+5�;б]U�G	�d�!Ա��Ln
s�qi7�����7Y�IH��I*���]��i,��g_��TJ:�eө;e\���Q��5�.�f=�8᫋y�}��B#A�u�ry��n�t�,޽��rr��i�|�5��JjqG��*�]:���ټ��Z��8n틭�/{��v	�L��u�g"mΗ4V'|�lF�*��Q_V�5l$�s9.ů'�<�o�X�^�P��kR��!@_��b���Z�o���h#�S�0Ȼ��T�����}[e��}R��6L��������<��h!��ȶ��ŵ��Be1��K�R�GНP��Wm��C}�g��3������Y�>�"�����u���6��X34�P�G^�A}�.�fc��b?S��Fkdkf����`I&^P���B�y���3$.�;9�7�e���n�m���J�k@���2�^��{�i�`�F�:��.�bkYx:��H=r��N��(���9% �͵+�^�3�d��XM�v�=B����]����t��:��D��ۇ��s����nX���oĎ#�޽�75��˘-�o��Kj�� ��K{v���6o0�OVn��Anc��a-wfdujn�fے�l8��,����
�"lBۦ×�lwnN�mӄ�=u %�qS�J�S��1��y�4A�"��퇝�X�͝�u��.��Pևwn�u�[� ��ov����)"�d���GFͮ�c�/"��>E�].���� �8�*����\܃zm�)��{ls�v�テ.Rg��]�4b���W* 6��bugX�՞�C���{$d��/��t;�\�ja1ժ�Lk��֪�8֓&mT%poh�3���	��e��l��x(0Ƣ�V�!z�dՑ�w[d����@x=Ko�_ߛ��:Ӵw���O7s
�P)��ǯ^�q�Ǐ<x���<�?�q�pq	�n��5��"rr�Ƕ���;w�}���o^<x��Ǐ^�:�M5(�F�o���m������N�5t�n8㷯<x��ǯG�����Jr��"�/�+H�!R�T	D�*Ni�M���;z��Ǐ<z��eB��	$u�r�)
3��B�<I|Z��h���)"A}o��/š'�u�t"˷����Pr�p�Dy�I��E��w$T�|v��{��ĂJ'��ו��W�׷nD�9ͬ���r	ϛ�|֒|vD�I��|��R��r��'��|u�>���w���������q�+�SR-����sL9ni����7k��R�[�'_0�v�ꕁ�RP��\�)�����ڳ��tܪ��U�)��Zi��i@�! F�E��"!�k��ϟoT_&����ƍts��rԉ4W0�̢��j��ˡ2�)�L�w��Ұ�yj����#=��t�><���&��~r�Z1��*�J׏5ߊ�L/�JeZVB��*��v�-!T('��.��SOG�Z�b�
�,!�>|v}�WX�_P{��z�9U
�Y�{��O�7��޼}�]/H없��kcX!{C�(|1�µ�p.Y=z��+���|��o�_�蝗i2l��s7��^�H��s V=��N�TH[2i��C3�
������r��>[�9�*{���R9�qQ��Nk�����Y��OI�#�:=#�(ߟ9�BG�������i�:v��|;��^���TT[{�^K0qW�y �Ԡ �
2�^��q�R�-��[���f�^��$oF&c�0J|A����˚����fZ��9z���'�!�kwUjx���[�1kv;��>��R��S*����?�Wn|��\����Ƥ[^b��qߪz���Rh��7r���k����s���@�����0�j�V{�x�72�o}�I./g��'�B�K�3N+W9��xBͫ���U�������S{Q�]e�I_XwWj[�=��6\�6g$����.�X�w̪��ӺPidk>�B��Yy�5���lm��������� ���e��r���-��׽�
 �* ����$i�R�i��*H$��
��<����>O����~��w� ���>j�B��3ٟCE5
6>VE�!c{�6R��e]�s�WG�G�7VF4�!%�i�Oˣ��~�<�.�H���U$�]�����6�n���Rx�5��|k�0��E�|`ا�4��t�b�xeη��w)�H�0��Nf�t]�
�=�ٝh�4OF+#���T7�Y�����:>����k�~a������S {Sm=D���8�NA��������C@���c�?0����m�Y�*l����*T;&��X9t��.�=���nL�y��k����~bLv��g�|�
͘zW˫��0�`���v�.�2Uv{oyx�ޮ>���	�H%�dɥ�
9�p�`g��`�ϥ��t�3aQU*裫T9���xL��YO���
����'�u�� uD�wd!�4k�]uE:��3��?	�GU$L�<�;J'\��0�}�[�f��?<]���}��9@Q�����ۙ�7AE�$�A��{����~/�ȏ�^
����~�]G����C�L��X�QCi�/j��c&t\��\�����;;��\�`�WSu%����DY�2��!y�6��Ǆھ�T%�;v��T����.ۛ�hВl5�P��P�|���S�=�s3A��d�g\X�R[�o[|:���̐��K��B��u[��\�Xʾ\V���suw�
�����r�jϧ"��G�J�ƚ@��h��F����  H H�=�u|����O�<ʱ
)$��f($gM���ZC�����Z�2Cdz�O�Ĳ��O=�+�s�y��ǰ�e�ł��cr�M�)�e�<P(ƙk�r�SJ~��B�-�ʱU�f1�a7�x�	L2K@� ���-.S5j
>b��>��|�*����
���'�l�0:�.���!������rF��w�!]d_(���6��(���|'���͜�N����'bȌ��X��W����<g�l�H�~ӄ?�>�P�ħ򕙏T�z�����}	�7y�N:H�ar"�;#<�C:KH1k�O��wM7G)�&G}*U�=α�Z��*+��(���H�	n�	�!��/�W#�8�K\��G[��J�\����r�%D^��Z��MMރ�%d\:�@P-�����.�{%�+��0�`7���:�U ,��h�!7G��еC���j�1�#k��"���ŵb8�`h9[� NxU>����_	�³�F+�k@�O-�,a��02~Ȓ�c۬-�$/p�W�pǼ>���>��w��0�,�r_9/�$��G"I>�����ngGxJǧjB��˿���Z���V�r����J�^���_tf���V0�{=n���p���7����j�ܩ���rIy�d�f����Kg�CDR���F���k�p�{�^�D�A���FD�	�4�M4M4�T 	 E7���s�_��0����'�LKm�:,�/+�~jG��WHX�4��E!t.)!"���[Y}��¸�t��'H�
b��x���_ߟR���Z���r�>4�Y��2:��� �g'q�����!�w�˾L����cH�c[��1��.����z2��3{��ֽ��
G<��L������k�
2.�pW	�4e۴FYkօ0�av���-)ͺj�a1Y��`zU(s7Զ�1Ǻw�vuc}U988���t�h��9�QZ
�aN����� *�0!.o��jɋ��΋�Ψ����Z���(��msV{՘��@�͔���pi<e�}����@�xS��HOn��9��!fѺ�G�{q�b�z��M��s.��ˌx2;I{ơѵƷ*�P�3��n����'��T�>a�]�|�5Pt��g�_�_O�ٽ����b��g�&��:��������Ј�&[>�(�1P(8�!��q�4i,�P��eZ�?��u	�W���n�:K{�,��������R�e61_^�����}	ł�Wl[��b�Te��Q��H��W��ۙyA���Kع��rB��$,�Ov�m^���^��|��F�^��ev���y��������׍w�6����b2G�Ji��$
i�! $i�
H��9�^s�g�'͙>COٛB�),%�nN1��{��|��p����t܌��|�����W3j.;N�����G���1jW>�}�#���?/1Qn���辑��@4dr�>Aq|�Pڗ�kbk3���5�{��k��*�,�>=�5@���o�%c�S䪓"�ݤ�*��3&���`��G��K�}�Y��m|���F=Y1�����g�1��^F�����1U�ݗι�:�d��k�VX����wT����=Õ�*�k/_s�f�����L�-��Ԫ�7K2EvR���|��%4��j�����1���S���g�H6`��+�7�M���{��Jw/�j�7�=MS²���8lj���
�+9,?x��օ��{�>"��9��]B�������J�7�P�[�د��R~�zDvTF ���[F"<̆�j��p[J�e;��;��d�i<.S�Ǥ<��{*���-��4��ll�	���&�� c	�[���M����X��d�1X�����i�OEC�����<2����01�Cܸ�g!�g��ҷ�7���&��x�7\\�מ��֩�TfMˇj'�n���y"���]���*}�|�M�a�_Q��u{�.7��w�y`�o��7���cO�:ғY���%�k-��I�k�ö��4�>�ߞp ?n읻V�Nݳ���.�#������җo|�����$_) G���q���foM����z��-�f��0�R7G&�V.$V֓�_�N0��%�gg%p�3�_�x�qФB�Rd{hp��P���f�۲���Y�쫪߷�)dY���8H��<{��P�t�{�=#�{��_z���Ip�T&y��m�(u��v��!�veK�k�c5�y.S�:���Cs��ӃE���BBv�f��N���.���a�����#q���͆�swZ�)�	�)�z�)��L�(�����q�w]�q��!��Rg�5'Ʊ����1<��9�3�R'��ڑ���2��_&>�93���M���ߴ8��r_(L�6`!j=c6es8O�o~ފe^�U�6���^#_b��$��r��s����[�a���O�����N�y����`�m?ne0��捛Wu�oP�����A>�GB@�a���KC�s�c��El����#�*<�$��4��~L���ϻ%�ٱ����&T8ʇ-��Y����k��a�| O���;;�-�1T����=�Ft񁵚�%:���3:�Z���	P��N�ܫX��R�D)£ό��������Z:�TT1��f��`��uʇ��=@\ێ덲�t=�^`=�}�ڧ�Dy�)�՚�S<P�k#5캏�����S��Zh�5��,�Ժ�
��e2)$i�i���F�V���H�I$���p������GZ�X���CaD	�.�B�3ӭ
�uC$�Ҷ�k�������l��twn������29C�z��d�dKl�ݮaCJ�ׯ���T*�P�] ��f,�@���z6.�6��ÆZ������Ͷ�+"�ToP�o1��£�o�����4��FML�ݯ���{�cS��Q�@��a>�Q���T#� S�:"r�9�t5?K#K@ܼޥu�!ΚE�U:��v��?�)/����C|tWʡY�߫f�e�N��)(����Κ]������,�pJ�nZٷ1��c�����sw=K�=+A��&5�*0��|�G����$Oz�Sg��@CE�0���=�QI���(=0W��@����w�^,n7�)�L堖������0�z���!jV,a��wM�MܲC�͜��ퟤ���9bL��Gޜ���j��2Z��W
<,-��Cc��vGt���^�#�j������ΰE�ߧ��?�FE=��'0}\�L��%1P(8"�6;T�>���mk؄����I��'������SBg`S�k����0�z��.��,�6�]P-mu��`NAK_�pa�5"�ߐ��Kk�@G��m�{Kv����嫡KFN�EΖ.�"���[�wl}UT�ն�>��S�b���Bc���Q�7q{�C�����})��)��)��*F�J�Ǌ6O[_m��?���>r�Ο-���a��
�||�c	Z������-��6!�Xp��0��9u�@��jn��xѧ�6�5��~C���0t�0��7�v�(���a�zz�x:�7���u��V��Yu��J���-H�'��C�Dp��|���S�2n���������;��ނ�{!�|~juE�A���3�Hհޗ	��b�vNe�QB������Z��Oi��L`�'�3��'"[hvb��x�jG2���K�c����P�m3,x�啧�:��ga�5���y�:}������:k���8^)�=�4r�X(�N%��7�:�w�S{^�¸K��J@����3���h�}�`BX��؏?)�li ��~��S��هy�y�4�����(٨C�����H���
��8�~UX�Իs�޼�4;��'��N��seq\Ǧ�PI���At��5���#]����ӣ����B��*1.�	�D�H<-����� ��^s�WlҢ@OEC�iC�������yQ�N�����a�����Bfd�\;�Z��Z��XB�*AXŗ��뚛e��O�o�}Y��la(J��1��#����y�f�K������w�q^�9�N08���[��ж�����ic:F����b��ɗ�4/ڹ8�둙	3$2{5e�cU:3Q������.����w��˵ݕ;v��v�vQ]�u�x�������#��~Cw�)jMb�����ɐ�w˹7��/���Qf��F\N��y�X8�c�|M;��ݣX���"�򣸜�;�����q�O�M]�9����7�DqЧ�x´_J����Q_-0�z��p,�A��$P�F�ʹq��Ƴ����Ⱥ�?j5�yҵ��éK�0�7��B*���`��H����>3
5G+<h���f>̢�k���k��l3��A�_5�.:��z��R�>̌3�MD�+�����K[��;�NZ$�n�tm*[{�D+�G1��}�ݦ2"'��t��yk���q�q�Ǧ��q��>�M�!~*܈��wkQ��� �}Q�C_8��Ṵx�F���ߣIX�e�G�Y�W����H~�Շn��=�i�a�虨�A��'6Q�ɍ�(=�����'�S�s����G�4S����l�v��Q��`��$;�@AƲm��K���Q;=�qD`�����7��ռ6�sci��ӧPU�kVb��8������w��㚧Т�!�O�̀�c~B��t��p�̺�v~"D�V��I@B� �J��"5��G��ћ�X�̧C\��NuY�ﾪ�e��[J�ݷ|�(H�Ĕ�j�#��@:g}���yZN|k^�&.�ʝ���c�NJi���wPVp�۠�t\���w8���gR�j�C�g��_��Mʯ����*,
hi��$i�*	 Ȓ!�s�����g�wϞH��U���OKx��B���|C� ��a�!id��Cz
�ϸTlGVk]�XOg��d�(�kחBOl�����Q��v��WY<O_<p})��������ӹ�9��6�11��z���u	�l�Ԭ�&�|T	�	P,��l	�3���0�'9�\L�ȭ�/���V�R��۠	R�&�>"-�'���<T;��8�@DD��=u����w=J�˺͝O8aX�J����(�Qʈ�̺���B�s�
*��U�19v��v�Z1l���R�c���P�������O��b�:��r�
iI��h�G	�Tx���Mc�'�{�K�wP>��}>1N�q����b���1�w!sD�]���BE����ه�p�j�.��P��N�a"ڷ ߙ�nH����B���j~�5�c�����m�-Ds\������9�ة���3B��$q��eK�U=��}�ҺSI��E](z���3i���C�D��}��0ݶ/���<�[�F��9}�X�DrO����.9�{�x��+u����4�ve�'�-R! ��"h�s{�l;��E�����)�k�9t�aZ�h�Yf�>������w�\7�f�җfa��^���n�\k4������;1e���w��˲��J��.�(�`��,,r��K#v��x4yPM�t�8�w���b���'8�J>��gs[ճD��SD��ILH�������񼏘=��<\�Z(餆<X�ɗ�Ib�Dg��wM��	l�3�{tFN�]�ޗg�� D]'�ݪtyw[��&�YAx/h:"�m�Iu�gK��7��6��gQ��F��(}��",[Y�(S�(Լ�k{����PL�]�Zo�:�Ȝ�=,c-��i2�F�Mw3� ��,Fr�
�3/�]��%gl�m�I�a�Cs�c��c�޼6R|��хnT��{�g;�uz��wշ��}�`u�tw���"��"x��4�je�w��7&��*��(�m	�5���������_.�E�n��u�9U�,�}Xm�R.:N>;}c��;)"����|�j�q8�Ed<X��Z��9y|�
�V���4fhP��5 ��vE�;��
=�T���Q��6�Л�X���+{�6
��D�f$̎a�۠�29����h���w�]��us�'��a&��+��WF:�u=�4�Y�rF���J�hŌlq��e�-�sE:��!kW
�c���Ս��L}��Z�^��iB��KLnIۘ��F��{:����Kcw�%��5BA0�Φdї�4r��$��f�9��%'��3�^$OR�7z�g;�H�Z�Vt�ӔU|�] ����+Q�KN�9]��+b\$��̺c��t���q�UÌi��bǤ=K[�}t�,�\.J�M��wI�*��ivCu�^/���y<���9-jN�˰{.Dk7��h�]�;d(���æD�O�JTK�n̣�*zF�X^�:�;��e�9ҁ�6�n��6�I648h��ٲ��� }ܮꩁ�&���3�ru\��=�{j=����jn�^���2���A��DړU��b��ۮO0dUh�ɨx���@���m����w���X�5$f#��x)u�ꫳi��_�_GYwN���/����">��Ou-<%436�ܩ�6����T�T4�3hᒭ�;��;�����Oe4B����ށr[����W:K��r���o�@��u�غ+2ɡq����Q��y���.�fcc�(�DU�yB�N�WY�J
�^b�[��B*z�LM��s�x�+nd+l%Q^G����ڇS٪�h�8L����I������c��^�J �R�Y�\wc��k-��M|��kb��2-��.h;<��N9���Y�e;}�1�`�ݍ�١nD�U �������Q)wR���E$��\��-�P�L؀���0��&�Ķ�"J�jX)��5L�˒!YUy궬R�i��n{v�cM�4�
���]�q����|�'*H���d		$ȕ$�}m���~�<x��ǯ^�؄���	!&�N;�k�gQ����v����x��Ǐ<x��d
�IE�$FIDdA)�q�x��Ǐ<x��r��BI53������Nì�rH�@�#�t�8��o^<x��ǯ^�5�%I����B)�EXwY�Tv�g�&V\۰�4��{qGҷ ��:���;�ۓ���=m�<�+-����ב��vqw���E�vV|��9#���w�y���󳓬�9�[�����㲎�,��N|U�l�\������Vu�ae?�����g������;�QDuٝu�_n΃��׻��{�"�%��;�r����\ݚ�v+��Ok�eh����}���ok-�Ϲ���{�,��2�G�V�M�����K�DB�N�t�iI�R	V�=�m��ߕ���]�ss�j�"@$�	�G�#&�|���\�7i�qg���=�ȗ2O�0;�l�B�z��3���L����~�j���=T����sWY�u�5U��^#�.�o��]�����鳔��J�O�>k8͔�[�;�f�:���b4yA�MN�ϯ�_c|a����r+`G��D��^
�U����N�i��8YS���/���t#����i��A�Y^/��DG<-�x_�Ğ�ŵ�q��������M^�WB�r��(z��5�W�P%�О���X�H� �I��/w2n�D��S�L@j��8|��T�9�"[�7hˊ��<^��_��\��N�P��"hzN�#,��i�z(X*I�<j�c|�q�2�1�� �$"gmX�r~��dd�1�s�zʀ�կaT���5M6�3�����㏣�s��,4
j��P5��>�}0�����ISq�,�L3�+w��蛼ղ�:%*�
�ڟf���.�z�8)"������
=���HY��������
tu�}~AB�}/ښH�6'�n%�Z"���%�~�O@0\{�:�]�)��}�T�_}[��_a)�����?�R1ij���!���Tmö�!��˞J��8Zwu٦wA�rBfi~OhrÛ4���mY�A���d��O�bc7����A�w�R1Vd��u��}�Y��%�@�|�FP�E]�bw���cѢ�vP����n�ڷj�nk�.::�=�`�C�<"�����U�К���	9ʤ|'^�1��..`Pz@��F�J�ȿ����O��O���Y�hLz9饻yH6b���}ӌPⶂ���g9H�EgK|�^��S]�\4!�qqq�(�	U���������_����͌�NM�6z#�g���?m.��j�Gdw�������2-���U~�}�� �V���v���^֛7{U��Q��{]��K�
���E���V3�f�"X|���/T�Dz�1��/�U'���<cFR�z�V��-p��|�;�S ;��S�$����8��[:�4�!�5hH�C����6Z�կNh8a��=��;�e;�O�Ү���9�X/"�t��F1=>G�^�W�t"���ڈ�@wd���*ّ����4¿c������EE�ހX�􍥳M,Kך}��9�_o�;�ב-2��+eE�a����!��<7�Q,h^�
�fQx��C�����s㿆�RK�����A������(���6>�.��|��!��2#<gWg���A5�zas��/9�K6���?4!���@��J]�(��������[���*R���������XN��L���0S�8nSH�1"^(S1l'K�}/�܎�,���o�}Պ�^���9�gw3��+k��e)�1�{�V`����勤�x����t
�"@���G�
h��Ti��,"]o��O��9��ڪGW�[�K�� �½����I|�T�Xn}zB��3�W/e�)m�교���E�>j�O�֔�X#�v"b ���@h|@��=�3�N���;�BɼZ:k����^����S@8��t�=p��O��FߢZ'9xh:�׬O�3V�^v�&J�(�/����x�Q]̒3\|���Mi@o����|��*��e���U��ؖ����2V��J$�8I��~��kf����~��
�4&�e'>��0���/�t���0%Sή��<]��R�OG(�"�3>�l����:=��������}�U�A��Tb��,a4y^�����wP�!>X_�8ہ��y@j�I��q��ю��n��S��3TP�c$�@��%�Fs^(8���.�}�Glڰ��B<���&���F���]�巕�u�v�����Y��_u�ꎝ"�J��+�/e�Q�;.7x�m�m�>�� e���F�YIvLWV��?s���˳f��uP���^���{��;P��r���辟�>����.۞��L鷫��Ǡ������:�`�'��(��\�_-��磕U�Si����'���t������G�OT�ɽX�y5ǫ	;��o�=��L�[�؂�i�Z���hق���d����f�n3�� �?�@>���&T�i��h(I ����;��sӿ'ת����hz������'����~L�w�)=gs��]�Gl�Gay��9uw���r/�ِO����` ^@��	n�f��ojO=��������S��f�y��{�Z;ޗ�����nuRH�L��"��A�M�?w�O���h�sw�(�3��3)R�GV]�N��O�o�S��u�,��p؍����H�.9�9��Nzc����H�duX����ׇv����;W0��%�خ�a r���I� �������ώ������4��,�ŦNp�-�c}ϝ��R�U�k�]	=�s��S�Z��k/h~'nė��^�w
��B�������z���Fk�`���b΀�	�����x�*u-�8I/O���-��a�&���!��ʉ5^���|��}*�=m��:�0{$������ݐ,�a��C_����Rө���a��;҈�^U��l~;�M��1��N�L�S� 7^�e�w[N�)��-��������O�H�4���#�c�4<�;�A$�n�o���9����?-�N^4]�ܡ�}@�u����M/��鷺ieU����r����rH�1���sbvn��:�Kٛ����@9��P���C��W8�e����������Z3!�}�*��w�hΆqN�๦Ӭ�N�Ws��)�SG9i�Q	���v�^'߽�^^>>K�� H���o~�u���*�����5�>��>�y��)�����זx�7��4��$���~|��ڳ�Q�{w�Ȩ���m�`o���2+v���G؂�Ȳ)���.|8g��Z0~��/���1�4��Aꁊ��7^�"Sw�G7WgP�x��ۯ/d^LI��KJǷ==���ō'�J�RGy��|yٵ��3\r�tq{�/�Ep�gF}�9�73Fo,���U�Y�O�]�|��
��ɔ\�/ɵ�M��^�n��Tl��\��عz����N(>=��ϵ�����a�0�he#��\B�O��Y�Zks�Klrj��\�ݘ,xkı��8����D�fJ~�<
�A�|r=9�ؔfX�qݺ:D:�ݘ��eW;���S�9b_�S��P峝�Y��}��,e��c+�]$-3:��9�gu�8�0�C<s��ZoWP�+�C��k(���/^�����!���w����hy��������}48D�"߈=�=�0�_Ddv�%�Ɨ\_�I�^y�uN����/;�����9JB��e��M��|i�v	޺|��2�%�+��:�OMN�e�����)��Ķ��\�.�pKZ���0�&u޷j	��@�o�Z�����2�,qܮ�`�J�4AfQ���V����[ڤ��uj���C��>5AM��4M�3>g;�>�����X���'h�t��t�#z��Y�o>w��uz��3�,�f��LͬKZ-J���5T�WtC4�����`���x��y�f�S�)r��0M1Y<�_+;a�2z��h0�xsK]���f��m�'L�����v��z���b�:.)�B������5ُq�m]�����g�E�4���|��B�
F��ңC^ġ�6��	�3�����Q�ȧ1 O*ɬ����*Z�
w�:up��"F���ɖA���q"�-=y����,���ܝM�ng�Drd��������=ޕ��{�B��R���6�7rݠ;�2�������ɨ��F�����~����%�BF�i�X��yHv�.�%B��x?(�v5O�Ȕ��qW��� ��5��o�/c���wjE)���b�0>�� 
Ȩ���c�WF7q9���s��+u�7{:{HQ(������sbOP���<�vt�\�U$��|��T�����S��\�埞�0�V����{�4��?o�H��⫚��o���5ӯ�1�Ws4�����$�~?0�훼�aJ̝�Q�[���]���{�-�º��ށz�9�ը&���8j�"����۩7{w_��^<����U����p�J���K0WXش��Y�5�S��V�Ջ+;�7���Y� |�Z���惄�?���%��>^H�/%�Au��}\;>��s�^?���� i��N�}�u��^E*�E�j�'�!����i�K͸��Ҕ����!���6���j�k�-��(�s��-��ސh#4�c�EK6��#TnVw�Lp�h�!؟}e��H1'�T|��_@���F���~j~纡��,��V��:������%���P��㲈c�c�!}�_�bb��4`��F���s�(ba���wT��&��^�D��	��1��HP��"
േ�i�fO����@��K͝���7��#�Z��B�ń�ls,{�F}U
c]�ܯFHh�#%,��q�-g�K�u�Di�ȕUw�]I�=�R����TK4o����ռ�������!�^0bѱ.c��w�U�P�a�u}�5�'�s�P*%= T;���x��J������@��=�]m=9��_N�����>0��$`���<��g� ����"+��dp/���*�G؜|}�s3�b�?M�9���<�^(��q�WDP{���M?L
rX�|��Ǡ�T}�J��M/�����wdj��z�̝s5���|7���r˜.��0[	<�ꤥ��x�Z��B>S���������-/���3Fm�Ul���u�������Y��,uʸ��(�Y����:�N*��%��s�UtT�#δ�WJ�N��Q1����}��>^H�/���1y���u%���:�Wv�y�/��P����͓av(U)2��!�ӓ����N�o����r�C��f�`�w[~��*G�mx@�r�؁+�19�>BOU�I�����~����Ɣ�$�GIG�/��]I����]"x�QaMAnN5Qp���|!7��۩�5a��<��'/�{&~ �������>|��˟܄�wA��:ދg�75
�ʠ��V��E�z@�.>e��0CZt��:�������<��^k��븪σ�sR�|f�}��RdF�$	p�f��i�>��g�se/#��6x��9=��*��L��w�\(W��39�mQܚ�)I�-�X堁ڙ�_@�@�s
2���y�%�������x�g*�P�_|��v�,����m�D����q����П���P�Ӯ��"�i�ճ��ߗu&/��uR��k
ѭ%�ܰ`ؘ3�F�9a��t�W�w������õ�	��0�l`�(׫��:o[SG>���S�@�z�+��o(Gwp;��8�.5��6��S�ߦq#g}��ˑZ~�7w�f��ob��wm��;���;s�+�o#nYEg���O�ˊ�#*�I/��]�8�|{���\�n��k�sd�K��R
��v�E��ܖ����pJ��u!���U8�n^t���47r*�T���+~�||||||D�-�����-(���ȱ���Q*�@h��zG��gt����M�����z���0Q��}��}{!���JS��W0&=���W�Zr��2{���xv{�Sn�W0��AP�q���p�/�F�W`�ó���#X��7�C\����Y棕�j)�]��4� �\^���ͻ�����V�x���Nr��$f{�<8T&~�[E������"���[s5r���5�י��=G���b�ׯ�HuH��}�,K��-W�AYd�WԆ}Dp::Ȕ3���ۊ)�=l���H���ێCq�̠R��sgH1P�^Y�T��fz_5V�񫓡n��Y�>�s�%Ahf��k����o@��:�_��5=�#��{�܊����t�u3]��
�����Q`X�G=?1&�����b� K����*���'��˧�ÛF7^N�P�f2�]�y�F�6	��p}j^��ԣ�R�!�[����c���t`! Z�Fl�']��3T�3�(�92_u&�~��Sr�<����U�
l��
��eB�~����߃]�ʚ���Fڷ`�s%l����:�8��j��?�k��֝���ΫZ�!�v�
�U��=�p� �\����V}o��@P>> �F�"�0�� �ܶ��^�Ǐs����K��О�Pk:O������ŝ]ܝ��s�e���r^��y��u�y��c�=�6��-e���G1|��T�&~��L����i|d�yҞ�>�>Z�˽�۳���sֳ1��-��$J�}~�(a��z<_9i]	�q�Z�<y��l��[knpЬR�խַ�ɡ�Κ僺`���P��[ �J��vS�)y�s��@���T/���ŕ-dԎ5r'�Y���q�XXFp"ߘAv.���bY��^oGb����u*g�5�����+~׫�Np�莎`���_���\c�t�N�?KΑ�Vr�r';�>̍۾{[Ì|��ù�yi`���9�XLp}�>���O�#��S���tVTl8w2���Q������U8w�Ĭ��c>,eO�gہA�@m��i pt�4?s��2��B��D*蝋ə���;0�m����V�Nl$�S@R4��
^���[i�_���p;w���ks�9��u�j�b�SJr�ǐJvD�d&*��y0��ȴ�� g�����6�V������a��rQF�֖-�L� � :�%��0K��|����Bˠ�{��&�Y!�x+}��(�0�4|Ɛ�q��X�8�ق�x��k$�#
��A�����j���.��ʝɵ;�W\��Uj���L�Uz�e_�5�Y�2��56SC)&����m�855���=�n������R(�ᷜ��s��*�^��+�!�D0a�5naC�n�
Sti;ڐ5���f�CZٚD�8��I�ڷ��ir�#�Bu�\�镳(��Z��;"���:��5�uѷ�T)�3��<��3�<��^f�&l�H�jeE@�T���E�8�U�H��w:�Z/1��U%�zuf�吶^�+I$n�L�Vh�e��Э32o�b�/V���4wb���s�]�V�OG$o���z��j�ڃ70��{t�k!���yߴ�ӽ[�q+/oF�ѻ��HH��$p�QL&��`岃vz̼9I����':l4�k/v�^��u=$�g�]��C��XD��{�����+�m"���)�u<o%��䇷�ʜ�JE�՝���8{��r3�;�-�G�K� �-��tY�::�g�y ���m��{ f>k��������@�s���[D���y_mM�E�1bm
�z�= X��B��W���δӜ��;��8$W���M�v5貞t[�s9���c2�u[VI�#��V�� �j2�1�L���t3�*.N��중��B��!�鵫��w-��3�^m�saf�(�C{����ޜ���#օ]��V�Z��';� �O���;��V�?�I��p��k�B�ay�Ur�A�}��\�Eˎ���М��\]C�����F��@R�z�ԧs�r�V[�6�t�F
�R�OW�A�9���4k��>������U*4��馦��4t������hɳ
�{�o��;��FP�n*}�z|��٫�Ќ54��.J����&(��r���udE�\�ww7���t-��a�H*x�$ݱsVq�v�:�iT�����֧ـǳZީ��B�L��4����Z9A��r�
�a�)�����K���j�Q���z���R���ma��Z/��8�_T�pane�Z�RĪZ�Umq��-�K�3V#���"7·Yʠ��]���ݍn�{O|�e�Ϙ�չ6�����:��G�oJ��L<���N	P�H�]\�ZoM�k;�,=H��,�w�w�f>֯l`��J�M��k�� �HJ���s�����-M�Q��|V�F����ҋj�0�V-ܘ�<�������ˑ3+�S�؄�>��2��`t�u�y�{���\� w9�%U|i�]�+	}xl�W���N�Y��i=ZhM|�3/�j���c��%��ǜ���nb�ң�����Ƀ�k�<��FEl��K�\:t����ǎ�x��Ǐ�}�;%@�'5������e~lU�|Yy֝����qǎݽx��Ǐ^�2!غ�P��u�y��^~mקǔ�:��O��8�ǎ޼x��ǯ\�26Vuq%G���<��e����@#O�>;q�ǎ޼x��ǯ\3�Dg�q4DȕSS˫�%CҐ&���5�|����� ����ȹ�m�8#�>,������;��;��+3�h䣱���F�&ݶ����Oz�Ug-d��b��Y^5���zXqw!�[������n�	w�j,�Ǵ�j������\���q�Dw�b�.Ԏ��zm"]��d[��[z��dx1�=���d���ї���t{m�e�%*w�9kKeٌ�a��E�Ns�����Z�>��� ���O9���{|e�����J0-����gʽ>��O'�C�.<��S�\stX<Ұ�M�ٓX/�V��N��z���a��]ڟRi>@M"P9��	"Z���>�c#�ц�3�͈���b����b��T;�$�z;�=��aZ�GU�=?y�Q"Xc��
�|Cr��D�i1UWۤ3���:�.�_��1�����P~�}��=/ȏ����a��P!�Mwm�y�ɦƆdw�,�J�[��&����>�|���x��nOOr�.^_v'xwN��~�#k˯d�c�V_],$�(����
=BuL ��c�󿹣���(�.�4��bՊ�]�R�3s�f����#����.�|��2�B<�=V�S19�#Elv�ޡ}"�M��{pw�e�^ǋ�;%p�ɰCa|�Aa@������A�;�ӯ�&�����&��/e84�K/:��>�_m!ޫ��ʣ�<�f�:K|c�="�Z�Y��wʄw��U��9�3�\W}�j��.�p��u>������(��m�h;���Ah �\t��X�s�J_)�l�#��~��{�rSV8�z.�Z[A3���M�(f��I�kx^4;7.���ڮ���k���;"=),#d���Ia��Mְ봷v7d0e�R�7��{\����p�PU����%*t硻�WI�L�I}���A{�#���}t4�+w�Vz��~��c����ϟ2��w�wW�Cs�aX�G�e�I�ss��L3�=�:c������^ �&TR��5=2�q�X;۴l������ҽ����O	��C�i*��(��ml樕8o< ��@Tӕy{{?(�x�m0;J}q�2�+�P��|�eW/�z�WF���O��~�VS����O�Z�>���=��Z�TR}�RV>AǸ:!�dXg�9^u.OR��&>�}qYZq��¤5�f\�Ԓ��=ɋ~��Κ]��>a�2�w6�a��;��Jg�c���8��Gc������yj�zs�*�bH�ټN�s�9����Ӭ��y��0E'�}�=�
��lv��64��z��ƍ���*�|W�Wt������(χ�qgaKT%QN>���К���}SuW�y�:H�}���ȁR�فm��U�n#�?��r��!*�}�}u�Z��=�{�}�g��=�S�?��rؼ�@��z�"�r�/"�0���g�W#�}�5�9[����&e2"���|��w/�� �@��F+&7��F!�ubUI�����P�[��b�>��}�	�0�w��!�T�'�fr�߸n��cj'�q�U-��z��Cf��>,nR����ʸ��.W8�+elY�1��rX�[���GrvsW��:*.z���Ųڠ��/w�]�����i�Uy[5W<�~T�:�1#1�	r���Lԣ1�7�>�-���敥�myl�vmgJ���pC�Q��f�<v���'�6�Z�r����Ʌ��/֮y��at&\T20_8H@�#b#Y"|x�68�{�o�����X�V�6��{}��iF���#�������HK�#�qF�R��3��ۚ��ۓ-hL���(J��Ã�^�k��HM)���-x�?��,%c��i���XH�������զ&�HQ�?n�g#7;%�W8X~�o��@�e����C�*��۔�s����{*�R'Y�"Jm���K�-�۽�A���fq�XX��V�OܷԀ��\
ޞ#~O�F�љ���f��˙�E���`N��P��m�w���0>mCP*"|�-���aQ��ءϵ�z����Hz��yW��<,��z�A��.����^%�d�	�i��.��R$N=V��:�BZQ'��&zTz��|��8����'��|`
w7�ƶ]�o�ˏXr��л�&
���Ǔ*E��㣌�{��R)�v�m�!���@�>��0�T9��gg��j�/*f���B����w.p�˩VGq&�'�5fa�U�YAv��Ի+�Y'e�Q���h}�v�w�����./��Ĝ^v����݈p��PG�%���B�ؘś�K�mv� ůk0�޷Ƴ]�ȏ:��%!�w������~�u=��-���~y�A��4[���T�v{�S��x���WgS5s��w�v^;�l�1�/+k���p���i8E��?Vo� �A+���1�Ђ٦&z;<z"�mD�x�Wu�{[f�����iH�h��{/l�D�GɈP���Kʖ;�^�~�I��TkN�õ?eۧ�̬�}�~�C9��}�������S� ��Ty�!�A���<7K���ug�W�=:����8����A�R~ag�y?iwM�ޜ�>�~��*��@�iIc��"�ۦm�`T�rķ^�P�u�u@�R/$I�<��ʓS�9bW8�n�
��4�����n�(D�L�WQ5�t�	�w�la��'�Xl�r�;\֑�s�NoF����YE.�K׻ �[l�;���ѻ�����Ի�#�<H�s�
�[P寨Wv<C��m�=�Ѥ�ᒎ� .�{�|�q��"E��[*5�^�<;Tפu[�2=LP�k�ߒ'h�� Q�eB7�m��F�x�4� �g��͟D�@]�%57!�>QA���`3hND����jk���).Y��%'���;F[��A�C�B�0[M177��/q����j��Й�o�U����X�*�m�I�n���^�m�x8����y@�f_eن:�g��ۣ���Z��jE�k=ǡ��N�^�8�]Bx-Xfn6�� �������뻈�<��v� ���=�B�Kh�.F�r<����3��b�M��`��mo�le�ɬ�ǉ�]T�Ɋ��	sV�Flr�E�S@R#P���[�v"��<2����.j�V����fJ�4p���gi�\�.[�X�'�WF��ħ��J��zOSE�u㷵��rj-���*
x1��T��!��#�FMv�H�=���]�l]e���]È���׽Kye��qς��׷�*�s&(!E���Lw��D}�Tyv�#�g.���(��dF�w�5����r��iUe���Z)�+�7�K�P��T�:���1z�}W����{	oF!�������OW���(s�Tlj��@�I81�r^5���Y�jU��������[�:�1��CL��1��t�>7ut�S�=C��	O���]���%]�#�"\
�q���w�6�S��tAe���)wI`X�����;[�g��;����(7��\c�����	�|�(���1�Z�|�����P8
�q���k�La�c�L���*��Z�.*0��bAv��ړ�R���3�'g*��*#U^�ۻhyܕ��.�|=D�>u�g
�9\xfW-�f^��q��w�k���n��Ү��E,��ݙ7T}9����ɛ�{�+�Og^_������o0f�o(�m���n�i�{�al�xQ�D���)��'h^�
�g�5�tْ`B��F"w�7��54��w������E'í��bG����f�����=_P dTg,�6�����k��R�^*+������e�w���ma!��̟��I�-�ٺ��r�6QgS�-�ԊV�%��:�c[�!��s���K�+"�b���D��%�XC�U��!u��3�[�<�vO�-H��W86�
h�ڜϮZ|xd�=�*�q�{�٤�ys�²��{�i�ֺ����mT�c5Q|��������W5O���>a�N�������
% (}�Z�\����Q�Y������o�553��6=IB�7���7�x{��_��J�bO¡S��*O�䪫�����z6��G����}0UĞ�kWw���/�9��W��@I�u;���dT�]��O�!�����Py��pen�̷��8R��iO��Tˆ1�W�s�1�[�q��7F2l��w�u�]������\�]'�"sK]˯`�<����ݫ}ź�����j_���.}h�i|����,�����C\�'��柷�����̜e�s)
�f*Ov; �//*9������Y�����U;�w��p�p�;�{%X"T����M�^��c� U����ݗ�߷�Қh}z�+W^��k���U>?O_H��:gǼ�v�dyO�ᯤ���A=1�����[�W��Z�W���)xh��Up�qֵ'˷�����JqC��tvf--Z���gO��[�~1m��_s�?Q!u�O��y���50��L=Bgn�k�Uo=�^��Q�iPJ
趱+��ZÝ�}�ZV)n�V�v�!n..�w��3�U�q��LS}˯S�O�0}�:����nLpBK�7�/�qE�Q����9٢�B�{r��U����j��Be��0�u������@^gm��3������y�UV{�5��Bz�H2,��`��vb�`gW���s������H94���G�P�������+�˻���C��!Y�c��Z��7WE������F{^��I�zٍi�z�1m�>]Yi�&�-���深��xb��
�P'�=1�yj�]@�bm��<	�y��q��lZ��{��F�a�M�Tg�2j�{!����������1}����TI�ݏ�e���n��9��p�Κ���*LR��>��{�o<��C��uH�qج�SܫY��"��.a�j�m�2�Y�PI�ܷ>��c�"P|9�I��y����J�B�[Ρ��w[n=���j�wH�]���Dc��gsǝc1hWe++7j�b����È��� �������>�d��۽�z��:N|��DSUΞF�I�0����>�yI^&�'���쩾�8����a�v7|�CvBO]�8;�H��I�br���7�8?|D���Б\j�*�|�2m��N��k��B��=5z��<.�׆*��}�#�j�6�w+��}�OH�\�S�PWSh1�u�OgU?h�È}N�%>.#g�"�<�H��r�S�r��{6q���54�V��E�����LQt>|a��@�G�Eǐ�� �g�����q��˾��w4^�B1(�Ծ,1Q��-馞Z���vc��QPDW�����Ұ��m��F1UN"�-hג}!�넱�8�}�H�wjF*+�J���!E��P���謘,�X��+�b�u�k�=�q�/S���:�t~�杻8�P�L��nc�{PLs�fk#>�~'�g���:�o
�
�z#��~ag�y?`/�8�%A�MN�y�Hw��v��
j�:�R�"D��@z���Dv������qeA��є�ˠN���r��ծ��|��R3B�6gM9�4��L�Bܾ�������{Y'q&)(�e	Ʈd�x�yؕ
�N����ƻB��t��m�}��;ˬc�^���\S����˖�Ky�]abw�&�MG�"tN��nΣ�� �	93�}�%�O����d*���5����Aa�硛ʆX[ԡ�fs�fQAu^V%e�Z*�t�#P�����$��L`xF��A�� �W�&%��dKݒ�OGc�Y�k��3���|ߧ��tx_�g|%�MCT������5��U�.0>���S���+�m�9�s3����m�a�P�c�,%>�z~zc�f50Q��(�� ��7���s!����=ga_M��-�U��?9��YG_�ǳK[���д��YM�8-"�N�Q�rw�o�ͽ�*����x=�����f�k����G'�b�<�A#PɈ������AS�+�F^�=N��g�!�s�\?7'�z��y>z�4&���U!
��T���Q��߹��l�|�To����2S�����
��|�z����vwMx�0�7h���Q��yQ��=�)�m����f�����C�0��aw�R�tG}L[N�8�]�L���+�;Z�6HnnǄ��c��ݨ��|�ԉC�1SA���I�}(��u����IY�;abOS����3$'�����u�93���}C3l��_E�6�Q��������A���m:�"�N�����ә��pV;%�WAk���PJ�9��f�d�C�L>9����cVj��ͽX�:=%'��K��yx��6{{����ٯ'�G8��%����/D���L�yjΙ+�ʤ�|���z�5m���L�jM�k��_L �Et&������\��aDO9�Ҽ��]ʹ��7$h;� ;�gH������T��l�($����������:��4�~��q�{%�i�=�@
#�u��)P�X5��]�p�f�m]g$�c�/�=�&Yu���p��9?5`�"r�N�v�-����pu�gm���*�9�^q��U�B+r$��#`=
ȯ�=0�׎�-3Ҟ�rs�B��Z�g��g�޵���m��i�䉸�Oܱ ��iY�����@-�����10�ܾ��f�H�[��~|�TR���Ww�5R��6ϾaC6<��}jV�S�л�YU���X�s�B�gg��y�1�XVQ6��y1�A������]�]��mb�iY
������?r.	aյ�����iLrR1��F�v�:t�%%�s�μ ���E3���?Qs���1�F��:@���xP��� \���8�Jv����e_7s���La������\���wW�x*E3�h*$+aV�7���}kl]:vj<��"�Z���N�.�K�yN�(E+�/lS6P���7�.vg]jK:>mn�:��l*��!k��t�.\la���������4"j��Ӗ��5��@���N���<��2��²o^�V7% ���j�r���]ɻ�4*�0���BR9ۺEWu�J�b4�ٮg)L�L]x�Y`�Uh�-9[�fS��+,,�sW6�)�`�j��p�yUU5�2��o�����ئ�t�+i �T���Բ>��͂�,���Y�F2Իc���=�w�y�Z�f��w�&ˠV��ӺbTU�Y{p�s�5�y���A��6�����v�a�i�Żz؜Ӆ����c�b4�Wd�l���7J	J3nw@i\�WL���������/6�8C���^��j�g!B��3]P��M\�'5](�Z]~L%s�̨��:�dj��Ӎ��eְ�& �r�>���s��j���/Mp�^���pn��\/�z�+u1H���� �d[�"sM�#l�]� �A��e"Y��|i�"�
�b$L�<-���hj��G�t�l�q��	1��_]��8����2���D������:Wo���p�Or\��������+v�@QU}���;R��^�Ҍ�Z��E^)K�#�veT����UI(�US�_��"�}�
�$v��Z{.��X8��]��{	e C�zM�1$��d^�X6C체Gj]����q�_Q�fޫRh��*��fv�	�M��V��leR���u�JՉ�QnFRv]��C(�K�pg���t56;����γE�o���.�{J��v���nJ=�8����N�.!��m���+9m6�t4�y�r�������j
*��7E��\���2��q�4«z��|֫�ٺ�G�k'�$Fbu�/sA�[���e9�*���t��"&�����9t\��]�t9Ibmq��=���->��0<��p7B�vVio�T�I6�W��r�F(��Me�S�#��.�R��ı�8���*O���ٴA���* z�dH���;W`���t�!*���JH�"��Uͮxi:��l=��ues�TZ��q��G�F��7����)���i�����v��44փ0:<�nC��aS���::0իӆĦ��\�����|�������㘵VD �z2PE�R���ܷ�鰖�Ofi��Ď��7�hL�]���>8����A[]�>�������g�S#6�d>S�:��&�YƚEu#t�Rw[]�a;�땋ֻj�nJ�۳o	��/�@;���S�OQ��]K���Z�e:M�us��*�l8�i7D{�����Ha�4�P�
�4�a8-@%0Z��t�f�V�3@��EѦ�!Ι7u��4��St)Mӌ�*��B��j��MCLP��Z�=����MD,�eu̅)L&�,���b� �4YY�i6��������n�Kk�����Yy�;ݧ��n<x����Ǐ=z�;T��6����Z�$�;��N	�
�\
iӏ�;q��o^<x�����g�;-�v�߾�3ml�����TJ�BFBD�$iӧq�<x��Ǐ=z�v��,�	*��g��slҨ:^֙�x!RD�����qǏ;z��Ǐ{��n��(��X�I~�=n���rq�ج���v]�u�g=���z�>/������z�eBq�d{j/�|/f����r���+���i5��L֋>3Ћ1,�˳����Y��؛Xqa���ڋ����n�ܙ&u��Y�rpM����Z[e�v�l�C�mն�;���5��`Gf�Y6�"m>n�¯����"��;Yq�ָ��2�̌����{�d�Õ�;����Π��˳��5]�#싙*��=gH짺#�p8�s���_0QE.�&�����iJd�@�Z/T�*Yt^���~1�SMSM@������`=��D�����`s�i�ސ6[}��sr2���X��굀x^Z����GH�b�
r��^�#Nǜ��hZ}J��5db"�� X}}��!�q���I3T��92pBww��H]҆yq\��w�H4�a8��a)��E�*��N�y��a�"��w��z�D�H�iE�D���ʰ��M�y���R�QkDȚ`ш;�Q��yM�����jS���j�Ʀ�LhuY `o���$�V�ý0��H�a:����xQ)T[�$��.J/+`�mv�|û��w|^�uk�I0�=`r1"=p
X�u�"���*2ze-��)�零�I�QRh��5�a�[v6���T�s��e����U5��a�&l&)7�[�20״�+[�f�%�g̼�U���qd��\10�j�̽��ֲ�M��{�Vx�,�w�v�-,��X׻vF㣣2y�8��nbhh���zuv�v��.�@ǒ�K|ne`�C�ډ����O�'u��r@tS�]�4Yv(�:_gYz#9�ӗ����fe�}oVG�N7k���Xi}���ڋ�tq/8sc�pb#7��޲^����� ���4����(���|�3}�y�9�+�ЈJc�S�x��]5zz���8e�-7����eY�Nf����Y��?P��"��%Hս����5Jx���ð�M^�~��+*<�'`���a�ty�O��D��n?��W����� �դiU^#b쾪���ܤ7{��s>�,�e��J����r��tb�6M�fT��������F-�6��k�Rz<����p��l��V9^8���	8ġ�J�U�ا23<^8(܈RhD�y���xq��0R�!�,ڝi�鞚��΁��m��"��;Nb�{~�VӺ.��=����X�F�X���������CB��2��_4],06�5i.w/���o�t����h��9���h��9��+�^tĿ)P�<T-���OU�R�m��[��&�|A��^u����u��^$��lq�/\�N��Y�W(�۵�s:�f��U�+���)����+.�H�_5��ik������E�����v���Y����P`entk�u��q�E��'�F	�n�G���d�\��s�[��y�$��f�����I?~x�}�+���y��Mo�\�7^����zT~wvs���.�[�^��������wΤ�qGc's����
� n��:��/Ӥ��Y[ޕt��BLG	�q������aj��'��Q�+y�Vk�=˦�kA�}�>h�&���k��n5��g/;y��ѝ�tLQٳG� �¥��޿.J}�9CI���V5�j5�!噁0��u���e��\@{����]o"����Y-OTv�mF�������;e�df�(	��e�?����{�0�OʦV��o6��j(	N�/ z{s��B���q�e����vzf騞� �"�w��%�g�Z()�6��[;���6�Ǵ��-��e�#uϪ�))��D'��:��u�F��L����:(�;o�&2��~��ǈ��FYh�̓�½�E�"ſ�h��5#��|�&�G�
��:q;v��M��E��tݻ���4�c/u�=�gQ�()��S�ǡu��{{�[��0ŪC]{���w��|&��%>oo.������%=�ilW��e��2;�,�K�����O��K�lx����4�M5M5D$r���3/�^V�?+}.���B� Cx|��E䪶ULz�w��V������.��CmQ݇���c���q`�8P��ԛ���ǧE�ܵ`�����e��ٰЉ�����#7}��݀g�9@{�����T]V�39w;�Ldq�7F^������PG0Oc�[�[5X�s5d''��nr;wq�o{�on��g���wO?|ﮏ�3itW���6yp�ʬ�X����b�JvX.��)ls�k^P+�Wrꭆ��n�g�v.v�2�2Y)�_΀�hGs�'O^�4�7qe�]�^Y�?WL�p���X�^������bP��M{�[!�pF���)�o4V��w_ ��q�#�\��3�s��O��.��<���`����	w�/�1�<n��߲K[e帄�yf��&���b����$qǂ������i�,y>K_Jh1sP�`�������2���Y����÷Ҏj��u`}����:��Q]��á1�P`ݼF����̻�l�OgO�|�Q�Y���df����n���I5:�P��@§F��mѼ�4�^ok7^�Zݚ|ERK���@ނnF� 8�"$Y��f��~//"B���Z����}zC)/"r.?��L�y�MV�����q��'�L��:l�;���r�s�tT�B���
6�w��Rw���)�7~�m��C��J��qM$37tD�wjۈY����~�j���6g��S���펢'���a�LZ���+XH�����B]�0cѥ���L�>��s8g���>�T�ӥweq�Ӕ{�>�V�MsEr���\�M�R���h#���[��JP�Z�{/�Ӭ���]�ipuL��x�j���u� ����9�^ۨ�
�{[���k�Ar[9�O�e���S�i��fy���eX��d����S7HiԚ���rȨ��̧�2�7p�9ُ6����u�礪�B����/S:ޙj�D���mѷ���66�4��'Ft���ݮ�$���)on֧�jesX�M8�i�nfe��ͻ6�3��*8�yh�6����0��؀�h�.�8v:���tj��z�H����nr�B·���(�'��S9]̹��ӄ�Wz���I0����<6D�.�༂vŎ�vF��R��q<��r����5M0#(�}�}�|�_�����5�;h��Q�+��������fGf���#�����Sm*�0A�5���R��8��⥲�CU:����n���n]�T���ٙ�N�����4z���V7�/�ɖ'��}L�oM�^�}���;��E0�N�Q��p������yq3�]{���^B\3�����1���*�L.����<�2uI�Ǫ��=�#�OBz�Ѹs7"�K�����ìj�0O���Αjz\��z�Mq�M��/3s�q$7ו�]k�oP���j>��y�!8��#څ߹{�=G�;��H��F �tXǱ�y��!ґ��Vkz.J} �%!���i��6�.{��i�6"�n�Dg\j�<}YP��VpA�V�}��贶��^��n�0���5=�+�PW��ѵ���&�Qh�Q�.g̱7{�ۚ���T�bm���NC�ӗEӼV�o]>&�l�vk�[��I�إo�cK�\��}�@���������(���w���3z]�NY�)�yA<�Y�з��+z��j�[�5 �v�^ɭk��=3gV��Nk%s��r����1���7y���i`�x����bnn�v⯌H�@G#l��b��.g�ǻM�Pk�O���0�7+��w*���g*�! ��=��5HܽdVޗӣL� n���.v�+s�`�-y�8S��.D���I��c3�՛����\*i�[Xǻ&�Δu��^������՝.�g�CS����O�cB�e�����`#}�lj��j���U�@YCyei�Y5�o�y|A�T��G���IX/�gI�%>+�W�D����{��RJ��1M�����G��D?[�冝�-��f�EYySy�ṵf�����5��	vJk�{�S�o3��v}^�Y���|�Ek��o.������+��H�ks��0���V��a+���M�W��WeE��)�{��Ii�m�k�z*�y%xT�i������w�u#���C쁪��9OtUM�aֵz&\�+�姍k�qCݣD���p�� ���iˮ[:�y}i�Q ���4��+ܖ"ԭ�o<�z�a�c�b鄱�����S��v���y
���M����*�X��n��}�Tv;�{�7����y���:pͺӛ~_a�=���U<��Wl����^�@�7�o�s�4u\�]�_E���=��+�>���tQ��`1�i��%��!�b!�%�}�Ns�fo4�ff�OI87b����]��^3�[nI�E82`43FGkX٫�XSS�,�����_W����\
�19��a��e�=ٜ@̌�Ybr�81O�a� ��L̹��2��Uyc�^_F�[��fm: �gm�Ik=I�0�@���W[3C[�r��˾�2��_;Z���v�=5��Iɴ6�)	W*��^WT�`}9����T\`��;dt{/p�j��cqW>�:�p�=���>+ۏ���oN��pU��/	1�Z��f�u��6���Y���C�OW����E��?<ޝ۔)�ͽ%��p�{��`H����E-�~F}�����˩؝})��s����eʣ9G�fdT�˫�p�n��{������}�!�Z�	ֺ�b�J}Msk6�F�q,��4K"^�au*��Nٮ=�qK;��z�u�
�R"�c}}����I�Q�P�u�v�D����Z��(�6�RA��F���K�P�w�������N�̟�ύ�A'{�2���Tv�:%��Z/My��w��ǲ^��jȒ�E����qKf<m��������į����ܐ�&��hH*���6�+���l���	���A��~Ak�jE��;da�o��u�J�S"�`v&�r�Ğ8�m�f���x1�����e��U8�A2#��9�3~�ٚ����xL����;Uf�NEη7{�zA���5C��r��t��Z��(��`,���#�a��*G[��'�M9��;�;����a�ѢdR����-S�9�^L��i���D�*.N�J��Ѱ|�G3�m�Z����3]7�U[^�8fz�S���k6�c` �(��}Q����+��T_��v������ ���[��[�tz�*qn�ң�9��#u)O]j-�>���,"�i0(�p���U�{�9̼�0X��)[�dӴv�,�&H���zD��Z�3�Э���QqY����wn�7=����ɡJ[�/C�â��6$ [��U5��j�D�m�Ӧ4�=o�x!Wݛ�2�9�4,���r�1������c��������[��BN=�>>>>>>?��U��>��Ep>�uim�:Gu!+��.;=��;�)h<�e�թȞ�UN`h8#Zm�8go=M{�b<�դ�-��
M�מ�9.p�g�XhV��|ݡ\������}
�
]j;�MD&��|����r�3Պ�"o��l���W1�|z�-�cĆ�a�9]	Lgb�sL���C����l�.8��v��w\�BZDj��5������Z����9'v������Z*]7�3���~�xME�f��ǩ�[q�u�ƍͤ�Q
"4;n���]s��k�+�\��׻�F��[&C>��~��eR��D�ӽ�U��dBB�sm��U@YEⓊ�й)����r#�)cl�v��wSpԚ�07ݯ�j��G7�
G����Ĩ�On�"���U�Kv�~�в[+��EK�5�rSzo�1+5on��	1OUB�5��*�2��[�SI�&�7af��;gV2��%K�,ǆ�5�����Y72��sy�v�\�s�\�W�sg�G��fܲ;C�fX��7�J��S�����$�y�!Hi|r������[4^̠i�ɺ�;ޏ���V����i��ݜIQ�
��m)�9���vRm�n�v�S���ʾ;��doS����aM}:sEQ�V�8;1܅�Y�R�)�c�Z�][�J%v%�FS���'F�s7���X�w��Av�c�k�ճ�a,ͪ��N�l��@���]pIZ�4����#{�od��>�߻T}r��
�30���2Jž]P%{N�;�'��r8W3��5펌w3��/�lk]��9˳��M��-��篸���.�zF\���G�����u."�&�֏�b��ǜ�nqnP��(�`���N������ �Xr��Rʐѝ���n��t�A��v�Q����ٓ�U`����-�V���ը���f(w��6A*b�g:b��i�}U��;�1���,S�6e�]�LD�W+-��t%��]�+=����s��um�"F��;gY'��Ůk��]h��1j�:b's�$��}�U����E�j�DR�w�ƻv7�8v�U�%��r��L��Bڼ�	+̓���o'������2���Qz�^��Gf-��z&�2[;�q�b�]��w���!�<rs@�j
������͞#�
�"��-*�6�#��q�b�#T:�M��k�u���n��[ӏjo�Hɜ��%h�\r��k��$�ش,H x��n�#�\o}X
���8oc"��h<r��譶xQ�=����e�q�R�pb��gb��Vc�Vo��P�ҙ�2h8;�.خJK�ͳ�k�[[�-w)���6J.��i�����W�.j�(vK�d���U�w��d��+4m�2����R�N��3�EN���yq� �>P�6�jN�
�^�6LZ�n� �PY�a`+�tSac����y����[��E�ߢ��v�f>P���=0��G�S�v��;V�RJ�XԜ=�gm4����+Z�,Z���nS�0뽹�`t�w7���&���[���턯�r��N����s��a�Up�7z9�ARb5������I��Y�vT��,���Ч�1��֎ne�a�"�;0���t��h��ũ!���eՙ�3�{S���r�[�R�jx���9��77��ʳ�QZ{"r�Y�y��Xr�S�J�%Y��R�t<�7e���㵁L�Or��vN��C�a,u������9cá�)i���a����$����J2H�ݓ����:U�B�_s��F(Cg���ov+s$��E᭹�'��R���+���*s9!��ռ���;`���l8b�Q -����Ԩ�����Z=�%-���fʹ�#�n���N��}m{fV^[���w�c��<x�Ǐ<z���dj��Sz��^�m�i�+�םm��۶ƙ�vE���޾��|t��<x�㷯<x���'j�֖do�o{ڀ��ZZna�m������]�2��*�UU*�0�)ӧ�8�<v�������{��R$(~�rK>{����`�8?w{ݭ��a�6�n��J�ӱ+:zێ8�Ǐ=x��ǯ^̢�ڢC�6���yG	ޗd�m�@��S�ٶr�l��}>�~x�Y�[c,����r�QvY�Ae�rgZf�,����:[6������^�5��GvѶ�Dڳ�E�dvu����][H��6�]{E�ͽ�J�,�Ď��qE��/N��;lE�bm��ޝ�K2�v}�8�-�)��d[Y&�"i B8jM�mfwZ�m�͑��[�)�-������>l��#�� ��!3�Chm �,�ưV�r��է����߯���� zdPc��o%{���k�^Jm�j��D���0ʙ7u���q�����{�����N{vxK��c���I5>����+�� �ߴ��7�¸f����U	��y���\�Y�ЇTz&6�h[n���mSu�b��Cg)��Dưe~y������
�Dōy��$b
��Y��_�Ě�*}S�n������zߧ�~��೵�M[+*'<��m���5:��W��v�0c��x�w�9BQhX(G��̆T[j�bu�]��oyw#Ck38rß�
!�u��B���Eob3~ ��]�1pz����D�Y��S��ǽJpL���󻞐�8��r��,�Q��U�A`�Y��:��E�f�i����~��p�z�:b穙;�g�@Z|]�m�o�V�vaU�h.��#��y;�a��S�r�ݻ���X/ g� \�UH�ĳ�����otL��;Ӫ1װr�}ӿ}ψ}�N,��O��7tI$�����Ӽ'��{p��USJ�V���4v� ��:�D�WXv����w4вI,B��jqHܩ���%F��W'n���7}�dWOV�0p~���]�̵H��J$b��7Y¯x�;���ʽr��@�(�����qP�5�޽��7������"GHM;i�&Ո�x�Td�N;ZUo�xy��o7�Ά^*�Ԛ��o{So+�h���u �4{L�6z�u��#�wxxYM9:^��M�s�����S���d��5�
|o�(�y�]����b�Uu�K��y�o��A�@�����q�C�8�� ñ���A;7��ʩ��f���lo6]
��
�ʦg�����R���¨Do[ҋ����K��:ڼ���]����)����;�@�S[i��P������V�%O����6�ò�^��V@E��Ba� �m�,Ia�(t�=1�̼�:�[v�W�ns\z�-�Jt��-�tQ��ȗ�mGĬ��I�p2�g��8?�K�Z���o[E���z�m�t�m��j�g2��T��δ��ا��gA�Qjb��n��ы�q�2m�]����$�D���:��b/uӱNdd��1i�u��|�B�/��TT�η3�r;C(<�&��MOm��ٹp�2��vxQP�"���A՜�ir�;��1��,���>��H>��-YxD��ښ;ja���H��R):�8����j��1���c.H�yw�Ew	�]������IR��Q�u�J�ijb��D Xd�[����P���v�EC��T��>��f�p�o·A�%\��6��\�^�/G�pђ0u�������Ź�]R�:����E�ÏX�a;�m�Ы2ni�er�Dnv1��ZumF(X�R #�[�c�k%ܡp�q��Q-�g����c�1�X'u��{�nL���]�\�]�@����k^Қ���t6u�:�S����ޮ����I����?�Ѿ#�c���D�]uvsX~{w���j4�|�&ob.�5;Ƃ8�6c���C�D�Y�X�͡cT�s4�jȃ��c��8�pF���=9\�l���Kn8c�peI׌m���7J���/E��Rɐ+V���r���~$tk瓵���m�a�)��#���ݍ�dM�m��n<������+�W\E]�9{L��+S�3R���=�����F���H���k��۬w�����l몕'82�{���������Vw��om�w���O%��qt�sS�U(�TH�V֊cѵ�A�ݼ9҂uo�Z^7u�r��"وbw&zt�!=C��I�:��g[[�g)4��㗌����3o+Ve>�c̝�̞��������K��O�ͻ��m�^�o?��C�9��
Ď��=;݀JZ��U��K��W7Og�w6:�=�W�������0��g�Wu{(8�����ܦt�p�AY6�`�SސS?�	3��C?,��ywMq*�ߚٙ�&+惄��{��uњ��r5k@���;,�ܶ��ȖS]xKb;���y��U=&�Y��";�<��6�z@&ߙ�n�˸�m��UK���|a꧚�MJ=^��4ݩ)b�
&�::,S�
��r��ca�3��� �8���8�OHw0:�/,c�U�!�V������:���کB5u
[���%|>׼D����GTrك��Q�|�����Vynpǅ~������;yt�ݸ�wT?�O����zH U�Y�h21ԀfF���wqyS�P��2�3�������r�%�N0��|'%�h+��E�Th�b]D>���6�^�)R�Ew.{��#�o��>=wz{��H��k�;8u��-��Z���uFN6n��ore'���;a�י&�2>+����Y{6��^���`w�������<���iP*����Ǎ���[%g�C���ܗ�S?�!r_gS
�7����+����ME���5�b�l��(��Ҏ�����.D��յJ�K܉s�
�#5����#��;��Gs�pZ5T4��%CKl�tEcUk��ZP�Y��Ϡ��B�x�F{��o��]�뒝�Z�R7�-�_����r�N7g!��3��N�]{#��6����t8�d����3���W���z�x�b�T\��q*��é��8��r�$��ꕕOh����ۙB4*�8�P�*�E1ĕ�[łȯu�`U�R��dfZ:+-�Xţv��ү����a榽�L��������=��l�6�Iy>||���y������Wl��G�1�5z�ㅃ�P{���"�eV�f3kv9��2�󌂨m1��~UQ􆵁�������|�pUSs ��W�B����n�e4J͓/<�X�P�;���@�]3��G���$>�>"��47�*�2��o��ʵ�9���B���6�qS�~oY��9"���o���|2�z��f�|��ʶ���t|y��	��1�c2K;�����w�}�m��f0�.�����t�)S���[���dQ�d�÷��Vh͌�'Ϙ.��yu{�����[w"��M[?}�i
hn�����{j�����N"����}���0��K��q�>^{6���>����3ך��?e�>��(��*=�JW�0�=K�WNyV�]O�wU���\�9��Wz�h�-���#B�Ǩ��of��=<��ʾ�83s&r�]\:���L6�j����aI�z+^�����m�����	V�;U�v�Ӽ��Z�(�L; b6��]PM�Ȼ���6]������J�'�K����9t��/Y�w������岸��-6��a�xVӎ���6;Ov�b��6&�L^Ono� ]_.�5
�k�D􉟐�� 1���t�'ͳ�9�N�IGV��K��j�\lb.�q�L}�[�/&��p�ݸz\�̓���خ]utL�f�$�>z��>�����7��7��;`��\�H��t��Gy�������9U�9tY�Z�6g�zC�ks���q���sfI�����U��Y�ۑ�;�V��P���fDdG䣧@�RK߼|||||}o/;����Bf�A�`-��1���:�R�=�g-�-�N��<qZ���+q��k(1f� ^�%�P��7O�X��19-�y�R�;2j����rw�N�X,�!��X���]�P;�F��*�P���M����y�''J`�Ģ^]}�O��Սo�=��q���ۮ��ۜ.������8���Fm�>�R�
x����ҙ��֚��%U��t��Ο
�t5p�낖�j9�.iћikq}7|%�d4l�gm�O`����[���N{�.��|��)wtq�q�x��r[��ȵ񶯩��t�?_���{����@�1��ּt)�[v�U�I��YZ��Y�Ķ��R��9ޞ�y*��?tz"�GU�tޖ�j���ʷ]���$*�f�ux��C^L�-�H��W�u��Xf�t8Ȅ4�,�a���~���pT�y޺�K(r��(�9�t�����i��L}�0:o������#���hx��8��F��P��՝��y�x�]��^�+K(L-Eڸ9V��Yv�'��ͬ�7%���;����WwrZ�Dp�{�F�V@��1�c�=��{.��s�_�"��E)�T���k[$��%��3<��fO����+8���
�ro%ݛe��M��(��\I�<'gm��-.{n��s�YU�&Pn��/��5^��K=���z���S��D��2;��A�\��ж���v���Q��z��HӸn���;]Q�;��j��exa��h6���8Ϝ�*��O�*�@��»���E;���?`=b�g��A�<�ʅ �e�Ӏ����F�ݘz4��鹖��0j��Gs�`��Ax��ܡ{5� S%�L��1�������>^��������a��A�"���^#H�F��{�C�me��u���%]: ��p1w>�7O�Q��r�=Ԅ�"*�[[&m$�<]w��}���ME�"������ɒ���\.�u�㰻=ۂ�m}\=�dvn[|���%&8���DL��g1}F���$qԁ�:�79�s������6�A}G������ήY��%��;�\I�pd�2q���5
�>ΐ���Wj�>������n��ڜy�����UB�xxT.��[��V��T��sZp,Bf=<���z/mC��-��Z�����g�|��Pw�m�����g���\��Qsj9�]6�Kh�Rq3���ץ�wK:⻺##��U+����6�wt�u�Д�To�K�7�P��t��uhwCB���N�`[ca��2Z� �*�a���,�pYB0 ���������9�1Oz����ߖɟl�̌�5Tdc���6Б
�\���l��q��QsJ��3"�g�+d���/cY߸g�ϢO�C�����z:�ק���9�Eڥ�*��W�31W{2�����1�j�}�����r��m�^^�[�����,�ܕe� cݳ�ʳ�O�&��K�s��4��y�,�H�B���:pj�laݣ�J�ʽ:hM��H���eK��x�w"^�SF��4>���Ŷ__Yjd7WX�vv%�6m�-n$���n '@���b�z����XD�BHR-����V��v~y^'��}�I��-��vX���]�"*J76 d�D��t"ޮM��Ģm��o��y��o0
rr���V)sťB��.��b&��%*�����&tCa!�X-��8�w$��q��<.���|İ�捑L%���L�98E�:'�E>D��ܫ䷱[��f�x
��ys9��G���W�B*���@�U H�Y�1��w2������Rj��=W:H$ǵJx�� ��{j�%wL<���&r�4v����k΅zz�nh�t�2����Q/[�����9C�U�1��G�a��^��aЧwg���9>[wQ.�U���pN����nWSkg]���M�t����c��]�˷�+0Sob�mWؿ+�7��E�|7�^�פǲ��'�v�%`�'�PΣ)j���Y��qOK)O�e�u:����d�ѡ@��袘��^{ɸ��ŋy��_�:U����V��{�ټeR��	��C8f�Pb;g�{f�t�o�8x��>���_���Ӈ��0~���/�ׅ�g0m	\��v����ڳb����U>&:�e��R���,q�T�S�Z�-�҄�ʄ�҂O/�r�<��vT]��7	GP.GI��u�3P�[3"���z]gG�����y�d�\'`�Kظ#���;�v�)7�yN�l�8�*\5ӷf�3Bo��2���ng:�d�k��#��K������V��M��畓"�]j�0��;)��I��ZM���q�5�l�Ojy��i)���s2�Tk���y ])�J�2�0�u��^"-t��gZOP�yͫڵ�4.ˆ�m:�������7�N�k�����!Lz���ol�f@�렼��k�����ҹ�R�,o껕�F D`;��t�{E�԰ս;��kz�z�xJ�cUu��k�w͌AR�3u>�0�]�c�kf�#o�v�N�Mu�9����5��]&�0-�7���L�zN���-U�\\ԂCzD��R�Q��t2����H�&i�Ք��ݶ����$�9�;Xv������+P�ƕ���ծ$�t��7���Zf6w�9�Y�Tn]c^��u�l�@V��wwT̠������2\3i�j֢�+�)fۙ���Bc��J��3N
�RP�(<v�O2�۵Ý�*{zdm�'5h�x�:�۾�����/AlU^f��Y*��\!Ԭ%�^)Ȧkc!�,4JAp��vT�=q��`�P��-�vq�0�N��H$::3xBٹ�6r26k�f���̥��"i�5��襋-�*w���9ٛhCB�d�a�\�uہkN�����Z���<Ț�$N�3z�q�˔�lԺ�B��/���Y\�CRX{7���gS��SL	s5���}��*��V���kT;Bc�J��y,�+�h��b\�[�-:y��e�p����\����Iu���\�@�����Xwo����>��#���p��V�ᑗw� ���=Z���_�0����m��!*"����y�h���v�l1���J4�;�1U�pͭ�ga��:��C��KH��޻�cY;�`�y�S��.T�����u�r{�����c˒�v�x'�ۜr�t���B�^��!l�
޾w��|�w+�����D���+/8MM=un5m<���A�B�6�q���|U.8���$9^k ST-;6�#5Q39ga°��-Ld><{5��LQ�ֈ���a�T���r�=`(,16]�&��-[=[{`*�\����nQ*G������m��TwCe�;3���ASafU�W��d��uq��fX��k��#��!�s�!�&�E6:�;.��*'/�Y{)���l������g/ի'�ӕw�y��ܷMaά��V��F��ۺ��ءI��&Q�JI����F�����5 �&�]2B�4���j��)�h&����JT�TZL�J�~uUD h��L� �D���n�PK�Mb�T^�mU�r�L4 $�?���%PH"O�Ev�nͶ���\d��L�%o�v�:8kwm4K0ʠ�T5CP����o��۷o��۷���ON�UL�ʪ��QR�Q*�-�k[[�}z���vg	�'"L��5d�*�����z�nݻ}z�ۏ^�ڃ�}oz�#���Y�md���ڊ[�P��Zr��s��%|wh��I	UT$�=z��n;v����n���~���ߵ�YI;�ps����4Vgg=��8�+4�t�(�Zݧi�UUB��!$#O^��ێݻv��۾�����ڿ\�ii-��F�l����;ksl#���{׎�����{�`n�v\Ne����I��͛hGmi��$�n�����lK�K+m�:�S�}��Μ{nC��M�:Ўe�����m�8f$e�;NlKk[js�j��[s۬�(:�p6�ZRt�����p[i)9׽X���h�DP�f)�n�����ڳ4�G)Bk$��Cm�����vۙ�mk�!����v��w���!9+����ڜ�s���ϑ�Y:k���w,���"f�M�����~~��������w�����Ń��w�0o�Wgt��n�R���8W12��ڏZ����D�H��s_��v�NV]h��"(�4�SJ*�'��������im0�ջ�ʴ6���[�o�yEwrKy1�Sn��Y�:X�f]Sa.!L���N�(\-=�·�R� �E�N�wGZ3����|i��`R���U���r�j7��dr�l�bk�#,=b�J��TGXS9]�����O�3��)��,����,�.\
�R�`����NP(ǖ�X��Z2�Xy7�U�M9��9�h�p�}� @��M�+{u��,��{Ke?��:;��ɘJ�^�KsA��+�Pg�g��0%>�֨FwH�n+h�\�ٹw��|u��a0;5T�,lDu�+ �:�^q��[��p�I9w�/�n���J�y�/��z��-AZ}[��R���e���P"Q[t���ς������H���椋���;�(���t�\��"�V��6�^pB��1;�ѻs����0�s>�#B��:h8V^!ݝ�����q�v��*��kIY�30�w&�j�P�_�d��ĳtVk!�ַMnљ/��.�hኘ�� ��f���25�}�鑊��\�Ԗ�����f��W�xjv��it�@���e7������sQ�Ȍd��qv�Dy�J�o߼<<<<<=ss[����4���m�j�~Vs�U�F�0��wOu;@�t����9�q�헋5K�" M�q�V���װ@_dr�^��%�w)�cL���6 �:fV�U{�.���T���s:������/+��������n#K�\nfy	Uy)o�Sf<lz�p��UN�uXjW�����C!Jڳ�F�\z�>���ÑĶ�׮��3ћh�ɠ|r������nڍ��y���#�q�'��=��\���t��0��s7q��0�i���Jbw�#:aI����Z{��@؃���VK�f�?"�n�=K���y�ށt���q�rm�)��@h9�҄�'JU��'����?g�+�<yWm\����k�=�J��������'k4�Vv��=@����yj0W�C>^x�Y�]{^)�G��+�]�x�VB�Z��cޝ�,��rr�'�ԯŭ�sr.f�N�<�M�]
��cwC}���]1;�	�W}Λ���Crv�{Spu�Q�dK�u�6�^ͭ��)*Q#/Rμ�(.tY6{��=��݇�&���/7����y��̳e!QW�M��Ԥa���h)�,vX��!�n
����W7uzD���}�6&���Y�|�tc7��!��Ƿ���QO׽L�F�@M��픾��m��aUnk#�Y;��yն��Ou!.��*9�B2���)�1�u�3/+�������C+�H`a���R:2���롸��<v\C�&�ij�㆝D��e�?���JۏSD�bk:��!0�_)��=76��Z"�^\Fr�cK2�#)z�R�aoUE���%_	 Ra��Ϫ<���N��P����BaY�
u@�㤳���誠�}�O��!�֭�6��4��6�cQ���@���0�\�����u�y]�hl��{�J�����(&\�/	z½�[�
�ѐC��ե��OP�<U�{9W�]�ɠs#fo����`O��S��(q��#i�y�vo��"�yڕw��hr�`������V��ڎ��6S�������e�Dv%fgj��W��}Β}UB3x
�����(^%C6o��1�f���K��+{;v3��:җ��zb��Ó;w������@c�bp�j�(�������L�n������˧�����p{�hD.������N�7/I��e��n��/v9ϣ�$W>��ۦ�B}�,!��`�y���m0B�1�����z{K
��ޢ�ޕ�-]bx�ƙ9�8�m� 5�������2Njs�,\�:�'�ޔi���KӉ t-�!Pe'�Rk���ǌ`���y�ЀTP�l1%a)��LrBG�L2��I�ғ����z���{bM���C?���^ rHN0��5?\V��_f�2�*1��ʃ�:
 p��S�&7�'}�3z�-��bKZL�͑�)�ޮ�� �-�����6�5�;���P�6�=Y	��,�"_t�:�2Qu�uz��uџ$o���jE�:��q�=q��6㹨o{���=\�����»�:8�8䅷u�%�=&��]$FŴ��
�ꛧ:��m�I�8l�s���9@J4����������]ۖ�X�^�'o��-V1j�x�ҙ5B�b��uvA�{5�5%�|z�r�z�Ꮰ�;4��H��S�F�O^��&�[�*�)�2�3��}4����,)
t�Pb��KL�c�1��5��<���;\�P��J~��.��]���3�P���G.��)�C�mCs�ѳ�o�ϓQ����P�/��%��F�v]�ݵ�*���,���d\���o�B���k��8 �z�al��9�,�Ff��f���m�%M�L��<�9�v���j���v=�y��)�Z&"bG�!g,΅:��t��4��$��c>�-�[a��(gfy�m��'�u4�f����̡[V(�R/���\�k��[����^��㊑���Pe��m�H�}��/�b��ل�]�#�s=�1{;�w�.�aH�<���$g�����y��qFSofy�:���?ng\`�C�{u���c(��I�훀f���&8t���C��X��Ⳬ�tZU�5^��������%��y�H�[} �:7tX�O��S�w`��ʼ�$_���Y�۷�	�Rt��]l�J��������R6���b�6o�3؅JZ^�u��jo��8�a�]94,u}vf�}��Qh�z��CѬ�-{o��^��X�MZ���!��,[���Ժ��obSI����*جq�GOky���~�����������_��⣨ꔙB,�؏Jǧ���`֗�C�udD�c3LC˳#4p��B�E^.�V��k�!��ve�䵂6�	�P��"�y���OU�^m�����^���;�߇'��{�0�{]I��u���#��J�r]�8����q�^�W��hu֮��
��$�}3x�"F��eѦE���&��hXdz��0���=�b�؍3�a���cs"�Cy�/��/7�SѪd���n�������+#�$R^�Z篞���2��g<Gs�U�.ʍ�}�R���O�n_�S����u9�G��\]B5y�0r�<z���J��Q.�@l�[ƭ0:��^�`d�E���B��Ý�j�T9�� ��ǫ8�*x�6u���}�s��0㶭u�gds�����(����^�u;jgռ�b���\A㏽��K$�1�L�2\��*�Єk(��*,C���|�.��:`�6L��vn��m;�]Q�LZlT+���ؖ�l��ra���pw��T���m�mL�ݨ�O�wr+
E|�}�Sڵ6����O�E�����ի/z��`]��?p���������W٧� �^u�c��H�ΘS����ȧ�+�LZ��D����df�՞�V�7|��S��cr=Jy�V�e|KE���3\rԬͣVzxB�''�K�63�>ac�y�r�@�η~�ٓ�F�#�ջƙ5♼rR0(C(�gg�?I0i�u�ð$�E�K����Y�2�C{";5vW�-_`�
t��)�,dfz��)մ���}5W۹+�>>ڱΏ<�uYz�19�H��5kA��]f����97������6��W@{�T"�dU?Z[z�!wQ�-�V7K�=֢�Z݁��Nx�8�%�:2}thŲ,S�ǩ�\�H'������2��f�Y�\�co��
�p�6&��b�(
o�We��є"��7�ѳ����;0��Vf���)��sK��i�pPg�U~���n�����vo�hIQ<ʕ��s��!�"�Gi���9<��o�#���,�7�j���ԘB�:�o+��C�y]@�z����X=w{����6��n���Ż�ԕv��CJ-��ҞF;�K ~����y���Һܴ*��&� ��Ig\Wu�s%��N��ף(�J�ӯ�.���f�i�����+g�K��q
=Ӛ�wZy=��>�3�`\��{1Tu�L�{a�-��n@~�FG(魯����_����Ñu�{q�80�0Ʀ�(u��B�gʄt�*�(�`��q�[j/�.�l�G*���%-/���q�l��m�9�a�NLn�0�fɲ�zv�֜�B�.��QS��i�^�il!��������Ҍ9������  N�z��W�&��<`o04bM�0�Xӵ��6��e��B����Qa��X�Pdf�hQrN�8���F��A�Wv�1'�X/�3���f��6��2��1�{��[�<u&�Z��WLU㡻F��oc�
����:�z*��zQ�>8�m׎����[�[���l�N��>)��hF�6�&�q���ԙ��0D.1�O%�Mu�U���Ybc��+{:�s�;�NJ>~)UR$ ^f'ͥal� l���4�F�� �vd��c���R�	�k�Ⱦ;2�}3:���5�X'n�rz�$lXSIUP�TJ)x�%q�*�����������P�����\��i�傠k˙��xLO	M=�R@��ff��3��!��oc6B
���?���l�E����<;=��X8oG��ɗk�̤ͫ+x���۽}
�t���{f��|���]	�ǥ�4�}����Hv�غ�O:j�b��a�kǽ��b�R�;���U�G$v��M:��/�󅫕D.7�ʗ0�4�Xuc.SwE�ϧa>��T�w_��S),���E��.�,_j�M4�K�}�t���|�ܪ;�O�ƶ[vFf�Ķi�M�T�)�v��=����~��7�+���QC��)���ZdL��{�5Y���ҥ�^W�^s���xt���qك�4��3�+ڋ͙�6~�ko��\��w����J��[3�fw{�5�1��xGnm�n���R��z7��]25"��s�+s�@,�7L��0�s(8�sY]����cf�#�����k�0�����4]��T5�f5V��إыC��5�΍���i��P] Q�s�x�:��u%'�����wEr[�:�N�7'CI�2\�nwdη��)5s#:4lĶ@����5�{Y��՞Yd��1�s3#���j�&w��Ρ��N֞�*��R�P�37)��,n�wTRF�����]�W�w0�V��)��m��Yҧ`]���ޞ�-�p��-�P}���{�^�
�:��>��^�`5u��Nn���ؽd�F�M���� h�Y4���1��?Z���t�8+^��H��/���2.�إ���M���n���!IC���yQ����Q���StR�g�]L^#�JП"^37�UE9�kT�/X?R~c*)^*�1L���!N�V�GA����[>C�+��cnm���ט��gٕ����Y��\e�E݅�{2�vZ��qC���>m� V��9�V��V%;-���Ὑ�2�̋8f]�9��;7�����zV�}r�5���)�:fV�ʯ)o�,���~���e�T��+4x�F��`ᦩ���e*��Ns;�WY8��f���1��i(�ٝ:��L5z�h�i]P��u�nZ1���Y��r _E�r�/�09;:/z�pÕ�G,��I�Nv�\�I5�n����}��U9��4���+H�����چ_X`X�vtd$�����Fp���,�e�ޣ:��w���A6T����J�H;9pV>f��jޤ�+5x�i*he��/�YR��evԒ��c�=6�]�[�����V�7��u�����ggfƐ,�!#���|P��^P���*��;P�	�b��:PZ봀|M�Vb���՛�돌���sw���G�o��-[�Z�m�`���ǵ�V���Gj#�q(�����J�7�DԳvb@ܦ�в��d��tæ�/q���_�a��Xm�M片�@a؜��m��B2�=�7V�a��Q��x��+F�}gz�f��z�wl�F�c�ט�˔�f�v�0)வن���^'���q�kvL}�kؚ�G��17P�$�o+FNx�!�A�\����FHoN��[4����C��ͺ��.�a��k�݇��N� �{[�؛�0:�M��^�I����s]���!Ԗ&�#�l���{�c���+��Q��{N�q��U(aL�0�Ÿ]�f�R���w����j�	�Q=Ym��j�9H�렭H��w{7�o2u^�m���Z�DU�5x�u^U魁G�������C5���Ѭ]!e� ���*9�Ia�ˎga����2[�˧ �VQ�{���z�a�R�ۀ��6��_Cft�J�p�'Kp�啳n�Z1��@��v�	E�S�>�9/v�v��fȦ����h�O+ې	nMY�f�i��un\�A�b��0�Q�}�4��h�X��I���C}���i�|�O����aÛ�l���b��Yܖ�����Rd�ƙZ��U�y��j�e.=�;;aۘp�v�Ӌw8s�[��R�I�6b7|�wG�џA�t�Ʀk"��!R��n��B̓Ę�x0fվ����j����s�'5�g�6ۭ�����x��p��A��K/(볕L���֧��n��[.��@&��&��z��9�2��XL�lnhT�m!A3��s�0.��sfҷˎ��R�u�%�yhj�F��/,lq�/����4��k+X5ⷸ8ٕ}!d�2�t4� �+�+쩪{�%�'ر�WMI�96��mp��TYMv]��ݸ��DB��\���ĩ����$��ȕ���ts]�������U�������:�NΊ��Y�5jiv5<�T���:�L��K��V�U��<��z����#��]ʞ[͖��~�ةY�����q�*�4n��qѕW(eq�9�p`�%�	��kB�򑧜�N��\8�q4̳���3wfN��=؛���f���g��;ݵMp��u��K3��.�R���l�]ݚ�z𕯼^]����<��m��8��9�k�]��r=8����Ɠ�
�S2���Y�i���$�A$�|A��8�
^�3�Af�A�X$�I�H�r��T�Ɲ6����nݻ~;v�׽��P!�Q(�T�6�d���� �l�'"��֗�B�EtUL�D!##`GO[z���nݻz�ۏ^w���a$dj�!"r)��$8�Ģ2�G '8�n�I��Q H�$$��޾8�nݻ}z��׹�!! 0�����J'fp��`t'$������RBI�!�i���_��۷n�^�q�ײG���\�QD�H��t�[d��#l���:Fͻlۿ�i���$�}m:p�Z�	s�E�� t���!�@�	[����̃�.E�ݜR�������qG����=��n���5�Ӆ!�ir���:GH9$�.8!�Br[]�E#f��N�8qs�6����Gs�3s�ޙe��b9'{V�'yYe���^v��mfس����^[��B����9{���ӠIB8mgQ�A�G.���Իx�3���w�k�&栝>�V�\隬J͉�c�km�����:��}�c����
�5~���y��o7���I�l�5q�g���Et�ܻ=w�܏��l@�ޏ?q�׽�mW�����S����4�wYz�~��)o�6;ﱮ+FS����h��h'��)�h!}�{f�"���8@<�N��Uq���l����j����_3�Ȯ�ZЦES:j�V(O�ك;}2+{^}�\.x��i?eȪ�15��<�ۨ$�%d�Y����^�ӿL<�h��ڿi�sFg�k+vx��"�U���!7�Q��L��f�����@���<��@��y���>[�Ӭ;����W� ��B�Y9>����0��pGY���
E�}�JL�X�EƝ������$r%0 o�<M�R
����u�@mm��b��5�K�7�����GBG�1�F�� imE5�a��	����0�m�U����<v�� 5��G���IU��]�Ի��Z�x��hb|v��YN]G�u�i�9�X���*������}��l���G��\��|a�mfU���N�^����
�!�n=�|v֭<�n$��ۂ,�����v1I��ɖ.gp�ik5��h�|]�˜齳�ji��]���������j�6�[��(�^�x��D{9�Zlμ���U?Z[W�O�MB��`4�Y���w�5�&�Vu.�lO�u�3!�qM���֌���0�TV�����A*2�3*�
U��	iF��� L��p ?�P�״���#~.��ܼ�c�y�O����^yOZ��G��c���� ��x��i�t�_�.����.�:tQ�Q3HI7^�tr ���x���U�U�2�s�=�;4�o���n�}���nDդ_�<s_��	�w_�ʞ�d���-���3e<?z��]#5���X��G0Sץ����6#i��nYk�����q��znӿ�rw�[��
�qf8��(٭�.�k=\(X�z����S*�f��u�X�$L�/��i�ݚ�kl1���5���F���b�++IN#T
G���J��ݞ���m���2<C�Ȯ���~��X���q�D�L����+]��{)wO>��k	��"��c+PTغ����pDj�.��0���L�]���4�Ji���+���'���8q�*�4GtL�b�ffW'�+��t0VR��	.�ΨA�]My��z>�S`��*�)��e
OD�\��1�F1�����\��ff茌Z�ٞ׬�%N��zo�WX�l�F �nn��\�}v����!U�``8�6�O{�S7�+��m�����n�7��)�t5 '|ϡ3�
�x,����W^&T���k{7���cL)k1V0Nw'z�{�;���>��ֲ*�`̫�հ�-���
�EZ#�J����G�
���߰��¾`s"�����pvv�U�}��v�gJ��3)zr{�T�Ij�Z��!�n��qK�[z��o��HødME[�y�"d����*�ϒ8�/-M�:�6ZV�ED��xf~|��Urt:/a�7�<��}X*��;��=Q�%m��2���DIY�(�q���7��g�md\z�b+�À��c��r�.眥��m�݊��Ӥ�Z�/��79-hM3���&D�9�����v�wl�Al"Qd�+{nK�����C��E�����F�
:�v�o�S�j�(�;�]�=�5����)eQ�� $�ϕ�oS����)ؑU�[�J���F:����Lh�MF�FoF]=lQ�Tn*�el��^Z39�{�ߴ�k��#�1I������3?�S��vg|�����<��ɍ�<��Z#f��:����[��-�����ˬ����h�&�\:Cٕ��QN��H�Ct�ν�]e��{^tϫ��˱/�RSG����7a�	1c�*�* �͇�4��Z_ͫ� ��.�ħJ���\�į����M�W<_^r�Up�^gzD@S!�oH�Θ�:0��݅qUȥCK)x�У)�F�R|�7<�����q���(���U�����(�eG�s|O٪�諲]~	~��d�m���6��8r��S�t�Ҽ����~�u��5͝��ޙ�ޝâL�A�k}�
#F'�Z��uK2�a����v,�7�u}�iL�6��dS��o�s؜�C�9���c����k���m�17��[|��MF�F�Uz3g��Ď�fW�$T[40�P)S�M9&ݍ���D����]Uh����S1B�D�m8zͅ��է]�~�G���xA>�Y�ms���
��;�P^�y�g8\畔�N��1� %�Z���>�;�[r��+�Н�yUo��1�/|�{��Uܩ�l޴lʞy�y�[�5�t�\���[��u娌���ɶ`�6�n��Oq�9�{m��P����_2g-)�qC��o�t�Q
�mN�L�������u��F���ޟ������
ߕ�깷;��a�=�
���`^�}=y
������W���η��[<̀��L��|Nd>R���5c
����#�uڻ�Wr��n<n��S���]�j�vf�WUPϤ�J��Q=�_�*��Q��G�2�le�E�ZQ*:-f+�^�YZ7��м#�+�m�_�y�V��
�=`s���lK��LU��[jT�ߖwOf��x>ᚗm;y+��b��f���ne��93�MF���ʃs%gs�C8�l��<}őDDoH�;!�M-~���1;o{�]�4�l�^�R�:�6Z�y���B8\�6ݻ�����}ȼ}���Y4jPlvm
pL��O���u9v���$?;ZA�]٩��6��F�!+8T:4u����7R�J���j�D�徺6����c���r;���#eFs�6w�g.q%�S=J�ūmK}k������ �o�V�K]��߀�κw�&�p��Cy�������ʙ����)�3wRE9����
7Z��c���l��J/Q�ʽ��@`_M��˻�ܮ~��H�O������Hq�$�wׇ<�qg/PJT��:SXX$��j��5/�6��'���a�h�Ja�t��u��Q�n��~A��33�hڕ��k[Z�.
#���������]��Kt> �9�Td��[�a�VU:7t!W*}�o�e�cg���Pn-������̋�uV��d"�3*r�W�R8ڍ�MDyO�s����=(�ǽ��'}������7��fr7;�Z���u*ꥹ���4�.����\�a���~�o7w[��<$}�M4��� r��x仹��Ow�|6��x^���G_cV��^��}"���r!�"M[�i��ǫf>}��uق�L�7m��C�GV"D�%);ܘ��Օ[s�Uc,M>W�)�]���'o9��cY!��1*�m�������C� ú�nT�x�� ��	[��,�t�f��+6(��rl�ա��)�7�vQUݺ�&��g�C�M쬣A9�QK��޳揞���|֟��s��=NUVg�WӀZ�&�ܕl2�0����7�s���/#z�t��μmܧ���:�a�*�ۏ-3�e��O#�Z��F�*��N7�5{���-'�
)<����HZ_��ykm��a��v���4a���f0��,�L4�(�_o:���Y��2�9�C5OqX��4�y��=(I�K�$�� ����3�+��]�#��v�ɣu�8��X�L>%������+�#�8Í�T��l�������n_=&�
�eY�LI����7@!��Svs��_��B���w��tT��pLc�n-��e��k�0Jާ�c��\`�޾��Sb�e�c�#]�����y�"�������]��yjE�	�ys6Y��߅��/3�g�=MI�X�B�s{����w���'uH�cDC@w�|Q��4��ֺ8%
�e�32�]%!�kr�F�\�t�j��-[�^]��՝�J%�v6l��aN�2�1c���.��]p��Q5�ŕky��c}�D����f8��H��川��E���S�W5'�x�s�,�2��=��Sv��rJL��C��+�>����������+��c��y�*�����D		i��^�)��tH�{�tM��,�E�	����i)��#�
�C���n��;�b堞�v䶶�4�4B��7�����+۱�4����X����l�,�q_Bɑ�w m1�&���W"9�9�=T�<Z���k�]�>�7n�]{��JL�����u+�b�#�k�k�0 �3�g)^�zs��c���r�����<��zS�vV�]��ÔP�\�W4���4��j�|oANȱk���
Y�x�z3W���owq��[d#0ϟfW
|�.�5ap�=�Q�5���`t\��	'��+S�ȫ\�Qݕ}��LC��j�����	��7a1^���G`xӺ{�i�h�`��^#z���`��8o\����|�����z7 
S�z��ٯx-�W6�i,Dg�B�v��ۺΝ���u��A^tbSZ��7�����Xue��F�c�l0���ǉ�V���x�_E�MU۽lR�<�29�C��qEr��u�C�+,��zx��yIG:v6yZ���=�;���zJ����s'�S<��x^p<� Y06Cdf���Ǚ��k'-5f�;95i���}�z�ͦ[:[kN�d5c��cۣ��T�ʻ�U�|���I�S*S��6@�w>��S��ؕ9[�h����)��1Ry��^������
��kƚ��_܈CU�t���8Oz �bp᩻�2���3�w�z�kˌ���W+��/�Ħ��>�\�lz8-&t�a��?M��hՆvv2M{c�%C�u�wl��W5��q4��\!�p�Y��F�Kl��T����o�-��*!���P=�T���	�����/UYz�(ڇ�|n����v���T���;In�t����k�R��[��]a9z7WtS	�f@O�ּ.��H�]M�`��Ɉ1云ǝ2"��[��Ɯ���G�m
�Vo.���X8�[G������֨����I��i,�7��\so0p]u+!-S�6>��KbT"��"�e��5]��+z��B�z��g�1	&ߚ��m"^	$Q�T�A�&�Y��*�I�c�I"�fY�	%fa���}s�����Z�}G�
�ֳlu���b�\�7���/���U�u0��l�`ܚv \�ޔ쌰��������r6=N�Nq���>�SǬ���]�;ZF:� ���o��v:c��O��q����+�=9؞F�:�nS�v�"'q(Κ�	BZ�<k��\}���(F{$�ƻ5/���ȩ4���%�ו�w��	��4��7uR� A��Ր6Y�y�C]�̺/�r����@X*�;�뺙+PGZ���t+҉�S���F�lmy�����v&�]b��u��a*:Ժ�,�I{�Aݩ���W>@ �[����o��Y����kwS��B�)�`m��G�b�y[��pϪ�Wo4��mc���}��������1���,V���(�U띇�x�a1c/;�F�H�S6T�Y���c^���O�(z�"+��>�#�
��@S��u�f�Яk�ީ	Q-0ѯ=�����x��;�W�^~���̿}R4" *��{��?քAA���4h�P@`yj��Q�$F,`���B$b	�$"0
FA���FD�\���9�8�wN�N]��$ (�d �`��$�X��F�d �b�A�$a8�wt���N8�]ҹt�	 �*A��@dB1��ӎ8�W8�u�9N�W.s��wK�NwWNr�\�9�t���9.N]�+�r�W8��W8�イda*����C�9�\�9WR��t�Ur���WN:��R����d �D )FA��
1� �D ��`� bFF dB ��h��1�d`�dB*�%B��0����0b��0���F�`����D ,�0��0�
�`"�`�(�����0�0+�1������b�*� �b(SU�`� �@`�( @b��"�@`("�@`((�@`�
�@b��@b���(�@` �@b�*�@`"�@`� �@`R�@b�
�@b��@b(�@` �@b(�րt�@`�A�$"�@`��$*��@`)T�B�(� �`	�(�
@b���� �րt�@`��$ ��@`)����FD 	TH$�bA���U���N��W+�td�@`�F?�y������t �P@�AQ#�p+���o����7�g����������Y���Q��o������W���o{�� U���������D_q� � ��G���̟�/�S��?r�A ��?X~_��/�H|�6��!�r������Q'��UF**B�`	 	�$�$"b	�� �(�H�X����H
@`)"D�$�$
D�$@�$B�`�`	* )b��H�AX
E�$ �P��F ��$
V(�X�E 	�$"	"`����@�� 	 b�(�b��D"�  �*@�$b"�")�F � �"�H#"���� � �� ��"�*��$�2
� �	A���� $� � )  *$ �����$����"�B(�b! 	 B �b!�$��X�b"@���B������O�dPI @$ �}� �������	?_����_B ������y��Ca{�x���~���q����}��A ~��!������' � �� �
�ʇ�A���QD]}�:� � ��
~�ڔ�k�ǣa4���a_��}�G���h�@Y�����}� ��I ���?8~'����s���"�����
��p�c�: �� �z�а�?���4~ J'�P~'����|�p"k�� U�=� �g��������A�;^�:�dEQ�`Pa���"��S�?��?��~!�?:��d�Md��<|�f�A@��̟\��{|��U'٪+ZT�*E��"�ڶ�ڈ J��U*���MB��*�R�D*kDT� [b4f$T$��IM���X�i5[Y�ժ��ՙ��2�64�-e[5�&�l[kl���jͥ�c靔�KK[���VV�f�)Ij�Zjڳem�R��+*�*���"��5M�e�����i�����֖�U���e
jɡ��m�P�-K5M��
��hm�5l����F�ZkMJ�٨[eQ#6�Vֱc+6�  [��_^��Z+7f���:���w:�ǦV��7g�{˭������v�a�Wl�&E�*�L&�Mi�{e��=��uv�͵��T%Gn5��UP�;n�m�P��J��  ��
2$(P���E
(P���㞽�B�(P��#��ܧl�۝m�{����]���ͳ��R�v���uݖ�n����'+��J頦����Z���D{fV�b��h͖���6̌� ;���kf���i����;cZ�er�M�4��%Ƶ�)S����m�]�K�;�\�T�]v�թm[[T&��]���[��wuJ��)�+f�a��bF"m�A>  ]z�Mݰ�)���lh�tu��T��5M�YR����tu,t:n���m�q�:���wj�GrvK�ִ�ʴlFm�lH�o  Z�cGe3#�u��\UV��ˉ:4:n��L����wA����Ѯ�*�V��:�S3�j�9j�k�v����6ʛF�ԩ
��k  &��v���r��k�h��h5nG+�u����sM�.��֭r�vՕwX}�w�8�s��^��W�	N��ݮ�Yf�mZf��/� 3� R����C8X� 7(�P���W  �` i8�Ӧ�:0  v�  �u�  6�@Ȫf��f�:�kV�  # �`  /v9� �'U� ��6�  gE�  m  [׋�@ v�t(��R�����ul�fZ٤���u%�am�  �  9��e�`:n� P l�n$  ��� ���  s���� -]p �b� }�{Z�յl͚�j�m�imEZ|    �X@�q�ր{γ� V�u������ �{=��  F = <�� ����Ȱ  ��O��*P)�IJT   E=�� ����*HF�Oz�ҕA��h�	H����@ j}�?��|E|����_	���N�mN�+
v�QvS�>(K�`�eg�����}_W�}�y�5DDW�  
��TDEܨ����
"+
  ��|�?��g79�������n���+6iP�z��8�Ӗ�Yc3Ps]�F���)�5��7iG��g/aP�h+U4K�pb+V�@�h[p������4I.�M��R!����b�p ��NV\O^�b�ҝ�۴�J�mce���M��'-��mLX���B��Z�
U��^Y$NH�̀��vo"�f���Y�l��2��)X(�*1���=��U�m��
r���*S��2�&r(��1͸S4�J��2"�Z��-#n����hP��o51-�[�0�Z,�P�0*�n�[�KT3$��Y�f���D�La�&Ѻ�͑����&'��f#�]���uoT�^L��u#w�ld��K"h;*�m�E�I,֨`�7y��n�I�͎i��^;MQ�tq��:wU�ˤ�wM��יj���t<���qU��:�b�ѵ������'w-�q�[u���æ�YV����Fڴ]��@�U{7V��;֚7��U��c:�!Q�f���&�dF/1͂��b[&���J3���4t[�1�e���(��wwZ)۰��f^���vN�ڷu�"��̦ek.!�-bVJȊ
��O�q��%��r�����~'R�����W4��#�r�W�8f:U�s+kv����Th$[j��cU�1f��x�L+���w����9��ge�$ͧW)�oZ��JQh�]EI�zl��5y��%�N*vN�l$7I�
hW��Eyܻ�c��{@l-8�',���d�5I)ub^
B]�l9A0���In�V�)\B�Xͅ����JQaQ�EV���"�4�`S���`-u�ej͟4���ų0PԪw���ޝAG�`��,cY��b��@�V7	]Xّ�m<r�̩*�U�a`٫Bq�[Nb�M��yk%,�0+C��2�j��gfج5���مP�����Sei`�-��e�6���j����Y�q]��1����y���m4�k*��&�{W`U�Ɖ.[�V�4^���l2��Y#+l �՘�M�5���0j�Gu\&��a����hZ3j�5Ƶ`r��-�r��M[mԏ�V`f�˷�Xwn7�]f��8Y6V��Jݼ�l�u��P��@Q��M]��/oEb
O"J�c��g��󀷯sZڗ�sN8]�vT
Pu�q�l��M �)�u��jƫ���/]0\�a]6Ḵ������ʺ�v��t��2j#�p�W����p��܍��f�`��oL[�����q�̧��6��Ѭ����"�ej����Z\�h�E,�hMqYV�QmͶs�Vx>�kz0P��W���q�.��Ԙn���.۹�n���a�VDR]�!M�wus.kU-�ȣu*�]� ��]hu�ށRK_+*;������j��h[ҵ�J�o�v����i[![�C�K�cdu����:��֋�Lk1�E�M%h9"9WL1�m�6]@�E'F9I5y���5��=F�݌�:��:lY����b̻8��%"i�xeB��V2%G%�;oL�����fѶ�\U�j�;��2lVIb����Z͛�[��:��KSl:o%)�O��WY7���,�.�Ft�7���ژv�m<x��s>ZB�\T�a�2���PX@��*++*;R���γX�
G����Ҫ	v���\����� ѱ �5utem雧q�/h��Yk&���J K.���8��tJ�ۚe����J�W��j3bKk��v(Y��{Ol�6�f���^�Ym��{^�[�ct� �t��.�s���*�i�,�q˃s
v6�K���n,
ʿ��jTݴF��=2ԢPY��-���mj�6=���^1�`�IV��n0�Z0�X�B��U�ef������0�:���$ٺ{f���Q�G��-���&�mV��ֺ!�â|d�ʂ ���6ͅ��Zw�yom�;+U��$k!��J�Y��,+�-:�(|���]A�����^^����i�%AKkn=K)Q׉lz����H%[A� ���pcl��kt��z[��m�yVv<o^- ���1l�e�r��P�(�*�v�v���+P��-�F����gi���=���]���n�\�kQ��bNJJ���иYܕ�e]XR�P�Ŵ�<�Ee&�vl�m��T��$JR4�fU�ܩ�f�6�@(Ay[7h�J7�K1H�T4��ų3KX�jl�JeJ��e60��e9qҫ6�,U���^�m�ÓF�p}*�A�<pi�1�l%x�F�TQO�Z�;+~���s��ͬ��T۽��@e�T�;�%l�EV|5����D���I���4��D�!�%B�n�7`�y�HX>K�|u:�&����շF�\٘���%#Xō��n�k�2�N�,Z֩W��{1غM�v^j���$鋥�T�+A�������ǥ���v��j�ۂ9��ne'@D�̏���D��c��&i2�0�kr�HQ���>��3q���9����QT��2�ZA���%HU*p^M5p,�-����L�
ڊ����%ص�"N���,� ��v�S�&�]� ��R����ɫ4�ˤI۩��M�ͩ�jT�X2�G(�r�b�Lݻ�ssɔ�S��M�2ڴi�)���A[�bc�@bȮ[ ��Z�4��/qmBf`�U�������l\�v��L8���6�ǈ	[²��6�Ev��%L����U<�V1�8���U �3mA����%��j�`�B�yN�V}*�`�Ze	�ʒ�D�S�T�	�nhe����n�� �]1�$Z�Ga'�&�&���nҩ,������%�+)[��Z���ɪO�Tm�X��m�U4�3`v���6�5ʸ۫�EZ��xԣ�U֚6R��}wY(�w�W ��R��&�L	]Y�sn�� �/)@Nڭ��������(��wK�W�P���*��$�ssEiXܰv*�y�M���6���z�V�ܻ%� �(���mJ`(Ykv��uk� V\͵���z���c ��QZu֌�����Rv���h5zǌ"�����q�ܭ.��Xr�fZw>;&tԢwK�+l�VX�&7V��U©��{����
kۧ��Ah�z�Dç!eY!Q�B<���Y`� @d�3p�tjT�V����x2�o,�3?ikJ]���z�]	u�KP�͟G>��<���eh�U�d$����uu���.�b�@D�d�#B�Տ�r��H�u��݁U�h���R�.�����#$S�ɡ�I�mRJ�l�.�f�5I��u�j^��bk��ela}z�̙�iؙ�C�ʺ@+Q	n޺{#M����X��{������L�+N��0'fU��y���ޑ/kS`l���3a� �v��5�0�� vШm�t6�lʩim�U������.V!��P�����ś0� C[��4���*b�����U�_٨TֳVS��i�A��e��賖�{o@ �X���L5�O��JB@�۳�D"P\�Ǎd�� 8���Q0��s/��K�xh�Y���i4�˽��iмf�;W�qV�C�&]�� �C#M{����G4����c�����K�$b�k
i���3Feʘ.�w2��\v�15ҙ�շ�%�mnT�7dО� ݔ���Uv-�[Pb�[ ���X�\�y=������� �T�(2�2��lLd![V��������R�:2�H'k(;,�fMy� �b�Y��+��jn�\��8v�Uy�挬 �j�*V�t�vA����t�
Y#�72]�C6��ف����.ޛ�bѱ���VL�w�N�ƠU���)�^�Ԋf��Q�6�Z_drk�Gc�nQ��)������Cl�V�!�l�B蛑U���GX�`��رLˎS�%�6�[#r�W*���xr՝�pQB�+}�n���oa�J�XYD`��+h���.!�T���j�Z�0 ζ��eA�XE�K�7�f^BF:{{�L�R�#[(��7 �Fl�- XB��|���%�ނ����@�Α�.��]˲��Sb�Q�In'YMY!Ib���Ȉ�wp,��0V�gH�&��Ɖ��R�`Gl�h��J�AV\�Nl���6Xʉ!�YbQe��+�����
�1�,� �p(�M`��M^LZd{��Q��74JۓrA7*�T����+�ج�%-l�.�q��(�(ܿ��S[��`|�iߵDwn3�"�WV�ŁQ
:����E��%�@t�,�QF�ϰ�c��b�krT��DR������8���grm+F���i�Fn0XۑH;�eau�j�sl\�V��U�Y�x��Z��r���a�9k#_%���Ma��we���i��K�S�F[���ʺh#��QɈ�]<�[�r�T��j��F;�%�6�Z���y��[ypm*��ļ�"�q+���&
�X��(�7 ܉��'XBa�j���A�V�X�d���	y,��h����wEb�����!��4���U��D[دJ��[���丷���
�&$qP2"��V��V�e��4Q8a�᪋LV����T�+]��y�d�݉I݇{�K(*�)��1f���ńb�f�7�&�L��2m�*��J�-i�#ˎ��7g�5�o>��6��wQX�%&n�ebύ[�p�۰��Kk�Ƕ��.Ω�T>Sm�+[���>���F�6h���NUӆݬWyPn�xH	���4"�V��<1o`B�a��ͳwF�6��������]�%lâ��r1Zi���Icv��n,9���R��	ge:B���]6�p�i�B5d�&�ڛI����ywW�.m
�t�y�l�����;V۶L�hdպr+���z�Gc�-	IPM+K#�;��2�
aW�*����6��P��M� ��F�6aK0^A���ieّHRuW�l:��Yze�"�-4r2	U�.�pm�{J���$��	+{J��NfV�EZŹ�Sn��vA�"�0R�l��B*��5$�s�gv�p{���1�
B�}53�W,곸��Ym!K�K���Z*"%1��<qO*Qʣh�Z�CV�l���#��3�Q�ͽ�Uժze���M�˵�������ނcr��8_�&�h��h�����]^�vF3�/: ]ј��gh�FN`b��1�*4�Գ1�׷j�M:Ŭ�Պ6t�7"�5O��B�`̦f���ji�I�I*6��f��,�A���:��{��ܲb����5��B��u6�V\��)�����;y2k�QW�%M��=̱-;j�"���RCx,��Is0&0�81	K�N�.n��ګv�ɘ1R��3j�0��X�J�-Sv��f�D�k)%u6�������W���qiwx-��]�Zd*Q1R��g�7+��4��>�#6�
̎ջAՅb�Q�Zb��m�uP��n*�����!P�2��5��b���T�*Ld�!%m���'.�ڸA��s:W:3\1�:QeV��Y�Dz
5����.��s�����c��&i���Zے��	����˧0>�l��Je��u}
�Z���Ddۖo]��"#U	̻�B���2����4+��r�A�������f��{��MX��g*)[�u��sQ.J�,��v"0�l�$c�Wc%:֣f��-&ҫ�K�tZ��y`�ҹ��i�v��%���Нa���yеE6 �
w)!6�Ć��(�Jҗ�J�[RQ���x�7��hg֦^n@S��������2һu�뷤+M����\�-U�YX�A p�Y����k�Y[OF�L�oM���䬡[w2��p�3h<���tE�g++[��6���j:�wm<��H���k�#����lѤ�`��b�I���!��U���y�t3r��v�ײ�d��l|��e#��m��Эe��H�Q��:_�'jaa���@�V�[Or_�V��I��@//�í�bM�����MV��fQ%�֥���$�'���P"��%ѬR��&�҈���HN�i^
�2٨�sC6%�гB�DnY�h�'kK��:u6(U,v,����p���Y��JnK�e��Rė��1��4h��*�'ml�7~wb0�#����p(�!���e:u���4�٫�[��b��!ڵ�e@g�!�H�;0E0�s[z�hm�Pd/5}��b7O7$-ZOcʻ�Dcu��[��VYi�f[��qfZ�yK���.-�gd����ă�9 �8�P´�.YִX��L�Tqm�Vp /fX8�rT��6bڐ���Ɠ�Cw�B��n�ڕ�/^P9�����=�	�qƥY8S���ѥ�5�
�ʙ6��,��`I)���]��(=Դ���N�[W���0*�Z�ܱ�7An�8�:�1B��rD7"�X��ɉ����O	{P]�l�fK���ݬ�y.iڒRre_֪^�!Ř�ʆæ�n���ZN��S0%Yw�A�[j( E��\�Y(�t�\��Ֆl�c]��vh���.b��ݧD�i���^l��̭r�0x�ق���3h�$�H��S��q��H��ݛ79FG'��)W-��y	i��@�w"�B#�����p���a͕b��+)^嬧E�<ˣ[��c�a����)�y�I�aͱzu=�Ͳ��8�6�I�M#(��GܭXc6hB�ۙGAOh��>%ި��� �.'d2T�b��ɣ�2��ٗE����Pv�DI�7,9e�CN���%a���aZ3hǶ�����K:�mÆ�e�Z�w��TeM	��V�I�6Xy1��Z�Gb���U��II �����D�8�@u)cjp�+s��=���=�j��ص���|�nt�r�|����j�;NM&gDT�2v�bĩ�]��\]\�9����XX\7peI@�-��I ��m�� e�{Cy\9͕�3$���+��۩�i�Q�k�rR4Aחwj����jhQ�^��c���b.^��r�kzE]vO%EW�v����:�*k���غN8����d��m�1�@�r�r��&[���|k�����#I��㌅��g��k���� ɽ���t�9b��-vkee��9��̮��%�Z� g}n�2��u )ݞ�KƏR�@<5�׏owr��̺��e�9��H��:�Bt�j���Q[Я�}��קP�e��;��u2�����<p�V��]�bJd-5��F��pj�=U>AC�CWh��o��il�喨^�a�C�G֨E��s6eg=�آ�+��ʾQ�ԥyk��<�!�ir�5������mI[f�ô��y�����j���b&��[�^��øZX)qS�̋�=��+Qi���SN��}�����z�-]tZ%a�R��P���+%1��WX��P�lS}�&�@��]���Cn��2�)�N�}�[F[����o;�	�b1��/uyod)��� \-|2��(om��l���:�m�C/���LN�=L�h�;��mmLr�ܷ�>@N�Qr�K)��Q�FsaX�;��IRIof�uI/ ����P<������m�.XL�o�i�0D��}݌���f�ֹeӢ�p$mr��v�(W@2�ԋ��3�p�]s"�ƗT���K-����j�͹X*X��h�qJu��$;�Os\��Jt-���o]���	��W- 8nY�(N��z^�]I��1gF�¶�3dp�69k�ڟ�v(�����>T��'�9�����襓	ǘ.;������]�zm�Yf��BQs����>��gvut���>6 m��r�KK����2�!@���n��Yx�o���9-q-�5ܹFU�g�׃l�o����s��|A�]\�)���桢&�i1��tp�%�$xi]I��&���0�)C&�:ح��成+�;uD읍>;�-#����Ya�;+Xjkx`B'�wXT-]q�h�T�+���{��&�l6�S��`B%X�J���bnݘw�O��/�V���+���M.;��1�߻�ނa��9��q�D����aS
��-:j��Z,v}��S�Gsk�n"�G �e:3��,��@ʾ�mE:n��b��\�>�D��v�Wq%���n�k>wzH�h���hñ
n�n�����|���va��K �۷�]��M����n�i-�k�آ	��u�rrsc�),ڋv^p{m��Q�]��R�'����}Rq2Ҏ���XomN���)��ժ�1��NV��')΃V��-Ӭ�E���+�X���&�"��@#3��M���4т���C:����`��m�[c�l�Y�����7.�`G�nͪ���7t�g�ԥ*�]�����9�C]V�F�L.������%�E�c,�����ֵ�j����m�yF?��}F֒�����59���x�ɏJ�����m����T�f.�����B��_^�@W��̙@j�3t��'�K�0�ͼ�
�
��dD���_�m�*K�M�Ss�������rյ�9:���u��A�o�U�Ɣg1B�W32/���	
Vv;+�U�J��n!y���w.cb�$*�4F��eΚ�]n��)���f�}��&5��r	���2nke:ӭ�8���:ᔊ�� �&��rXJU�:0��C��H��4�Z'z�4��@�>�1�����(SLJ!x����k'\�Fu�=�Z�9��Ep�:�l���?p�:�2ٙ��}��'�YX�@0�n�jh��q����ߋ���yloj����.�e����N���?e�Ɯ�KC#J�9m'�i�����
�QK��s�qp���ެ%^`V�(�ٿNV�f�n���K�\������|��ھǭ;y]{�C����'���r�.���ܮ��5�'+aM�۬aT�{!zr�Q�]i�w� T�ܩM�_gf�2�AgS���U(��qE0e��U�"�ubf�B�L�6���Cx5ư�]�{�O���"]��.���"��3�wQ���^��8�n;�A� 3�G��m��k]�D$�*M��f1P!�O+n��Bn��c*�5�T�������/�BY�mf>j��ۋi�R1Ř݈�ծm{��<��^<�#UaV�z:Ws�Ժ�
�aq�ê"�*be&{GܔO�r��P���J�c�-�睺�5�R�#_'Թ.��Q�)]��D�mju�,�J>�����s��"�;�Y�䍢��U���e�>%3��g۪���9r!�ݰd%u�twq�t���ԝo�x�$��e;��Sы,���s���U��� ��k8��f�P3�o:�.���_]���	��X^Eԫ/�L.%YX���8����@Қ��g4Z���vzc�Q�(��85`X��A�����ɷ��:�SE*���x��یsůtt�˹(&�x[�75��Vӡe��o�.����i�6wh:+��eY���kXj@�8�f��-�n�i�V�dJh�(�S�t��z���?[�撁��e�g,I��wRe,X�����,�>��kz�v��LեΟF�:l�x�U@n.�%�<� ��k�/�����&�W�Xd��.⯷H��YW�.)k����ͼEnCM��Ƭv�hMɄ�����em�DB|1�5"������D���5�%���Y��컢՚6X�k �`��v��{����,z��1 h☝Ŗڼ��3�eϡ-u�6��5 ?�0{�1�z�glxfr�{fA�v9�����AXp8�b���N����uuv7*+79����&�^َC/����tM��8��FY镪Qy*��p�G��n\}����s�]�!3r˨���Z=�]�	o]N�w��9�4�&>n�[V'_I�[��f�Xݜ jð�#���&Ԧ�}����07�cP�J;���(���a�A&��@�	ە�9&oK{8��.���3eG|�����:���;wt3��4$&���Q�9�@$[ǷtfУ�S�V��Ԓ���x�;:x��0d�1�5�;���3�p�z�UZ��m� �Y�D�x5R���Uy6��t{H�i�;�M՘vK&F�Օ�T�^qX�q�Apy����}A;kyN�RT�fޓ
�u٭�x�s�!��9w�H2�E��V�`�c�fb�ۭLx4]���[��#f;E҅�\U����C6�G�t�C2����lp�I
�5�6�LXht컏���̮���ܙ�
jW>�5�o'|�Zd�oKs/N�h��u����n'�*�>m���miz3��N�Xͽj�&�{Y�@�C��*e�P����+B�V���=fmA �҂��ܣb��"�n�U��lU.�qf.�մOd�g?�^=����M`[o��
��֫iU�6н�v����)�H[NA�Zxw��Z��@��:w�
O�6��7�m�2y��w�
�-v6$����6h��7ȃ�[op���Ŗ��:�^S�kz�Q��3ۢ�CPb�t2r�a�smp���ze�3�]#r�(�.�ɋ���DG���q��mņ�9i�֕�ף*m��b�-���N�fY�0��!Ԗ�1���P�#���=�kr�%EJ���9�X��vrs"�6,�N�t��@%֬Ds���)��3�ľq�b���,�n���.vL�V�3��^���d��2�T��Q�J���'��8��c�!�v�{�D�x ko��A���~.�?���/!�}�v�t�B�YǬ����;�v-�5FJEϸ�J�el�s�t��p�d�S��x�
�����];5ղ���
#D�$���ʻ֭����Z:Q�K��W6�$�T����n��&,�#��Ρ4E�V��N�^�43�K��X}����e8ͧ)Z�Uל8P&��j_fc�ٰ���[��b��^M2ы��u���:6�<���Q�
*�t�l�4j��j��u.�v����-��U�zʶ�wZ�4,�G�kp�(U�2!��h���-��Xc��J!����N�<3�h#��P����;ƒ��NI���B��~M(^��t������u3x�8�r�Pn�O�x��ɋw��tݷYς�|��]�R�oG�T·��bg��J�"��e��b���,�{���A[x�"
���2J�Ϋ"^2p�ʱ�4�z�_�Q�y�͊*�(�5�$�s[�1^n���L$9Rݿ^�;kV���V�Єr���^�-�8J����l��<�7]i-R�N`��y�^	��`I�.�*ubS7E���D4;��t��V�tƉ����|$��/�H�1f?*V���zs;[qi�9*-�ۺs+K����`�v�]�G�AXf�23�i�4�s���U�|-r�:U� �F�m�c���b\s8�e�i��/tpX2g&FÂ5��֨X�ObV����	l�{K��g�*:��!�Ԍ�y;+9v�L�T��B[�wI
��
F2�v���bg��!1����f�ޥ���7`�[}� f�����Sb�	Z�2�$�[��9�Z��'
7e�ODFB&�}ی���b���s��eN��r�]���6��,WS ���jڬ��E;;�s��2-�k�-ʽ��C��|%:�����^�u��u���(��9���l���+�X�4������m����e7���.�	��T�k�w(�Y<sF-�7�2�k��tn� �Q1�h3����B��pRe�w~��r^S��aPtLy��D4��a[�u ���j�Λ�n��(6���!�vU�o���0 p�k���=͸[��*l\�������
j����J��<���m�fsO�A�N�;>Bm`�].��{�j��i�*>�X���1WYfm>�-R��*[Г.s�in�@��ǌ���oN����W\�I��	z�=G���9s��o	�jở�^|��}Z��eӄr�a��j��lZĕ���s	h�3Y�;�&mH�L��;9�XU�E�!�/�:w���;���Vi�fs�V�զ�iP�%�����Y]�ӎ^�rr�q[&�J�JL��_-�S(wQ�c�^ͬ�	������(�XxH�Ġyaᥙ�r��e'�Ca֒��5�t��}3j͂i��}�+2��p�КC1�BM������e�cli�U!ye��ԻP�\�E�eg4{M91G���mA�\F�x��i�dD��l	�'��N*����S"hbv��n�s�ڏ9N�1S����Nm�vdyPq�@;�:�H�]r����&��i% �k�n��د�<�2����"r�'9}��1���ǹP�گ�.��:��L�>�Z|1�#�`.���	��P]��%R�N�m�S�rp��2���g;U�C�VD9v,pދ�N7���Ρcw�,�7kC�E�f�ޘ�Z��˝�_AI
Vc�#%*�jt}*%�NG�Cf܇�#0�c^�[��G÷qe���JF�s4*��ӋE]�ȡt3[�J{� �<!qqg`��y��rc�{:;���f�S{����t�Y�Ԕշ�ɺ62��A��&�1�M��2����N��ݝ�� �v���d##_*:�;�)�����%-�6�/���Wc��O��R`�T��wo�=	�W�d�)����#Y�a�Η�`�XF��C#z0��9����]�FD&�^Z�)e���ED��t{���i����Y`Q�[a�
���&��zrً�s�z��=�r�� �LQ�!��M�5w���2�8ڢ����7uGEK<\лt��n�F�`v��rÓ��u��0�t,t��:
�+�t/�_M)��e��H��a4��f�Rw�s��	s�&�ȧA��ɱ8v��.޽�MI���w�� 0�κ�d`�ru�0lA)�����s1)ܝM�O���2���p�-8s0ݞmB��9,�4�6"�<#<��_P�*Uܫ�=y[���b�����d�(�Au��p���w���܊���N���!��Wb���f��յ��?ػ��j'g�m΋X��[2c�e���nsخ���A��d������o*JP'[2�mp��
�Nr�t���;�����=��<]�Lm(4X��<`n�[�v�K(��%g*^˵}�{:�k�~#��Ϋ�u;/�0��x�X�}Z��fq�nraG��2�&OQ����z����w.��!��T�"��*�`�`�:��]ʱ���.;{�p�I�O�=u�����8�A*Ԥk�t]�ksN�{�m�2ȃ�z�vr�:s�9�,n)� Ӗ�Xr�1}l��7���9od�6��]�6Ѽ�̵Np��s�΢#B���7����E������L����щ�gd�n��%i�bUj�ƮA�}��%���I+�6]��w�r��$^j�Q��ظ�r�a�9�Vִ���g{��KV�x�t�;z]�)}L<BpB�Θ1�ñ�i�Uc���JDct���RP��2� ԝ�]^�Iti�mSPBu�|"#dޔڨA�Z�>��1��T=�
+����󎿊c�ؘ�RضT锳
�;o�2�h�G���9/iܻ����cL��+gR��1��:��.�L�i�qU�֪K�F_k,[Ҵ⏕�ޏ�P�G���c�̦+N�Ts�PṒȊ\ג�-�">rT/�^u���"��ì�dd͙7#���\ضW]쒚[6���w���]��u���߿�( ���""�O����Y���3&1���y%���{����P���G#h[��v:s��f��|� Q��X�f2!��'q∥�Tl-V�wfn�孛͢��{[.ާ�X�;/�����}d�&�)K 6^a傖��L�"ۨ��{��93&'*Nj]�󍨫�e�N�ml��U�|Ⱥ:|^%1�m9X2n��Z�E�V�_|vr%E���7&�w' �;һv���o����ጘ�[�V�0����f8J��S^�Sp����ؠ�T��|����f���G��UvJoP�6�(v�ۃ_1�v�kS�ЄS�~ɘ�W��e�4.��Ж���������]��y��I�H0�oZ�.IZ�mH;9C]��Xz�gn�#�:%r�J�OhnT�E�w��k2�:[���M���)|�oD�®�|"z��wW2�e��[�Ӥ�Q�pޅ��]l���1-�vAwL��wc]y��>��2�7�M�N�p��,��_}���B�;9�d��G�ʹY��B�+�;	nmr.Ϋ�.Rr;��U)��WB�qas#���3gV]-��7K����N�M�X�\�z�^�D�x7MZj
�ڦ$l�饭:�L��W�����K����^�g}�W/2.���"�6*Y��k�D�j�У�R��W��yO���Dp{�E�i��w�>�q��%�ꓺ��b�?�ǬQux��'\^ƭ�H]ַ2���:�;�pu�Pp��r�_wN�Cq!ʚ��΢ͨz��@&����G^��Z�$->,K���Z���އ��V vd�D�2�X|rB���^@��U�H�%݉}�(��J!P��k5�2��,^Vv6�t�I-�)ZT�:!������W������29 0��)�;،�-��^����C�GM.�|'9VAy��U�Ik�S���ͩ���hX��2_i�Rm�Ҷ��������c&�F�p�Q6��8�uK�!rt�T-lx�z,q��d8jⰩwmû�X^s�׫�w���(I��Gxow7yq C%.�귙�6F��[��T�`��c�uۃ+�-��qц�]����l� �ڴ�Vq��#�6or�ވ��1>���о2ې�n&]�Z��	 VNo�M���T�br�����ڗ�k}ֹW.���@>g"؁RmrG�b��A ǃ�]��T�M�X�^�\�Sb�wnL��R��3��Uv�#DU]�vd�^m�n_��7e
ˊ�6L�=	p�=�D^<�� rpIɝ��y�2��Rl�l��(�f���?��ݭ`�W�=�oue퀆S�X��2�J�1��S�H�BoM9]��K�hWo9�����}A�o_˃x��q��5� �3I��u>�î��s�Ck���]]=��jl��j�۹0D�
5ʻ���>�L�U�p�):�sTʨ�c{��Y�Φs��+����.����Sz��$�j[J�Mc�Z����yL95� �m��ʷ�M��u��B�t�-��P�P�h�q��sn�	i>:;��ڇ�
Ƅ��+�T*�ؙ"h�#z3ՄD!��DS�h��0rlۭ���vSH�R��u:g������2���NGkU+�P��_-p�I`b�칕�\�ǡ-\�q�U�=K�v����ƧUφ݊��S|�AI���ڦ�y�
�1�
=��(a�Vg 
H�ˣ�b�D����!A�Y1��b2�^��r��`�TА*�d�V��S�96a{���[��#�6�S�B,K�Pr����U��;���j��Z����1>��\&���k;R�ӱfr�N.R����%̆�S1���a�7�9XY�K�۽�Vڼ©�ťL��jK�����9J��nC�j�pl���Q
�9T��ث�"IZmof����
\�2ě0!��\���k�ƞY�t�U�(!;��ՔZ��(��kN�OfL�2��X��o\�c��:���]
!�����&D͹����Mc�г����^m�;J���7x���	�X7(7^�n��� �kX(r謥l!��2Q�GWo=咲'Z��j;Tj��+���_E�#k�c+���n�]�M�C]ɋ�q��D]�˵�PM6s���g�,c�Kw�n�]ݮ����@6��d��+I��>h�X�����B�ɖ�]r:�e�/���p(�<zg�LX�s����Vv;��Q��d���a6GK�9J�\�J��B�<�R�'L�3ŧo��iZ�N�0�͙[�z�lћp�5	7�躍t�c��1B��+&cwV�d��$ɮ�Ne���(�vW=1=�L�C3L�(I2�\�.��Z�`��8�ܾG�l+mGvs�����wg��z3���ڃ�I�E:�O;.��GC��Rj�ju����	5�1�ovȝC����>�+ȕ��[-�-,�E}N֣��vΫ����Z���R�1Z��
]����s��b�drMd�Џo*WS�4,�̺y������ �9\���[S��k&8zիqL]w�h̗�g5�Hn�.ʳ��W�Y��I�G-�w�b��'
Le�Wډ��Pen�#�Sa���ܖpMڅ��BrSSUӦ
���!)�Ư>��}�e.c������M�[�X�:�� 'z���h=��e0H��h������0�P�$�=���#����v�l�Qmvh[��Sf����b�NÜ7��a�r'N��:���wL�2�W,Zi�x�,�b�y˚�:.AY��X��3�M�v�5��%9�6Q11��K��+jf#d��R8�f+'��6�DI��7��k1��]��oۚ&u6wo�ثJ�]�/�`$�	5Y:ݫ��x�o�lo���Km}4��w3��׸�&C�Sh���!u�Ȏ����H�R�w�.�������lپ/�ՎD�������O�h�^S/�dB����5��[��.%��
Gnre�swc�aVP�e����CV��l�4�󣹜�r�A����C��<���r3(ܼ�0t�4���i+�q��Eǁ��ƻs�L8ɼ��YK%_V�Ġp`�� ���N��_n����.���ƪܻ+P�t�{�x�]G2v���+�6���s�i�R}���P�ɸƭ ��u��qws���oi�(�.�"�}�bc�#�+��R@*]�Sř[��J�Gw:ӂ)� Z�6��|V��g:Ej��Y'��W+)2gX�x
�{(�Y�B����p�vJ�[X��m�JC�l����S��4�0`kI�ZS6vi �o]tu�6��nB�;�ӤN���E(��ʀI�
��{�����d����w�9�n+��.e�VNU����f�u#�$��V����S��"�>��.��(:�l�Du'�Tݽ�`�^�1�A=�o�Z�U5�pָ��	@��y��or�ܾ�):^�7�&�g����e i+�n*��7�6�S���*J�0��ݍ3��y��q�N�ZCl֨umҦ�s�;V:�-��%+����
��A됔ņ�[�U�F�U�>4��)��job�}�@���vUX͉�M@�7m��u�l�R�T�-K�b�T��u̞��GR�����*�o͘�]���9+1�R}8qiБ�t�n0'�����O��7�:����g�2�:��VK�� ���1�yU2��&\�բj�i�l���"���(�9t�B�s����W(�1Xl��՛=z���*i��W\�8V=o�J����#�7��+2��:սIU�G�˻�<�%���Ӥ��������4/����0%�F\�I]��kҏWT"��A6�K[ńR�����i#\)�iB����Ֆ�����J�si8����ZX�z����3�0\�z��e>ӊ���5�
x]��kWP]��%�I�/��i�"�ą"�1�#��foʋ��Z��f9���c������f��@���*V�{>��X]����!J�R�Vp���Z���Jn�e��뫖D�9Z!�!ͻ���
E���f�����YF��գ�F-8�͓h�2Wor�x�]����sZS�B�
���4��q�A=0����j.��c��#�i�ev����(toP�Kr`2H2���%bnd˛���}.�F�J�[�����u�7��{H���7�&�$y��7WO;�M�u֦e��6���Ֆ
�Oq0zě]��S��N����oT�FU��#՛7�͏�K^]p��\5��x)7*�|��X���`ݞ=WeǇMj��`?*���)T���2�S����h��螥�/�
L���6���k�ru��j�P��U�Y�]��Syf�0��Χ�E��u:�
���0�P����m0�1�9����8t��z��8�VU�k��ew8YV�����Vt+�!dt��'}��S����w
��+nM*̼�0�)Je�o8�&q�*�T���ma��ɼ�����-�;t�R��3�*��,�)-t�v�>ҙ�G+Q���gV���cr���Ȝ�kl^��R0���Jmtj�I�t����8=�[�q�Ċ��wf�M��+7;W*wq�y��N���f�r]y&�2�ǮXv�j\`�u���8{�7�m�5֚:�n��ҕwV+��
�����Qn�~F�b����	'�C�����N��ŲV3�*�˘�NorcL����A�Xr����Tsw2sّV>���
���w��[g��2�;�t��N�˚^*iL8N�QHP��kT���w�o�+h�P�p�ԳA�7}0(m}��eh�w g+��O\�_��m�@���q`�gd�0+T*�sя@u��� �`=�����&_r�I��է�7ƅ�T��j��0k��s"�Y��_Z8����7]X�����	qj�R�4��{k+h�����Nn��-�pWE��}Z���
�7[ҕ%5����YP1���ڵ����u��Ӫ�u�
u���ݜ�8{�a� :���i�pb���c�*��f����Nު:�,�$�O�J�Z�:�j��c|/���L�̎:#Z�k8���w�4Ćq�"̙'|�\�I#I���LǙ��v[��=|�;R���G�"�%O���&���ȝ�`�[Pkh81%�Z����Y�Ү7-���Ge�q��=lV�ku�6�S�%$��ي:&��a��t��1�nɛgr�q��� "#��X�=`�9m��������D��׬���$۝�r�p��.��`�qg�>�P;���[���v:S�d��E.�z�[qǄ:PF)��y,���wu��g)8R[]�B���P]N\f���M�t��.�7xG?�싎���*�S��X���+���Kfi��	PW<�N+��Eu�A��K_n����j.h�Z�N�;��ϻ�i�nK�Ճ�9��u���j�Y[s�����B2�(86�9Qj�X�"�?��)3h��,��0��K��
�I�ۮ7x��i�#��pV�@a��ob�~�X4j#H�}�[�u�'�9�����L<�PcE�)(v}�혉�}�p^˭53r��pREӸ��1.�4�lo6�V	b�\(36��l]�&@�4ϥm�z΍WY���-�t��j	k���͒���h(�J,f吅�E��*o��NC2hڽ��v��W
ʂ��R��3dT������fe�%W϶�2j��ྋ��>���Ʉ�1���N'B.���eЍ�]l��-�L����B�jXw�^N����P����ܬgP����֣qū��;A�"�z�6�p�3@�d�Kmֱ�2�_@]c뵠�;-3�d[�j�堹u�KYL��%s��Jt��`_V۹L�A��ju�%�˕cE集e�81��U���+�p��T9�u!YJ��ؙB�m��pǒ=Nrĉ��{C���9�{�\]�۶Ͱ,��TD�m���qQ+â�$WA��`)��a���R���z.��*h�i��7�;��Ty��nk�U�䖪������u0�4����Z�6JW����\��C:u-/��$i��7[���36�� Zr��զ�T �v�8gsF�!8h��v��P1�Zwb4�[�
�.��VtJ�e1�=�ʺΗ8mr��S4�}ҹu�&��oR+n��(1��6�G��4���G��u�$ɰ�G��E�t�-�!{��Bu��� �+sC�cPZ��uYq�Ļ��:L7cz�Ag��c�뾜X�R�Ge;��q�(g�u�ھ���*�������u�$�ngI�`�ޓ
�7W����k�ĭ���i^OC*��$.kO���K�������U���+8J���D#��հ	�tr�\-�YU�Y�J�]YGs���`�{�Ccbl/�q5����ۅ"���P��7�tV����m��Öz�eS[��s0�jh��yְ��Ac-�Be��ۉ|�+%��n�ݑ"�M��m<V:<B4��6�Cp2�ھ�Vm,��CL��L7�(!w�jo.Qǒ+�����s9�g&5Ɋ46�[���# 7�>��i�[��t����m�Ώ̂���}2�wI�9��-qB�1ܨ�lxcL�J�Ć]�ri�ݪ�*��l��Ԟ��e��6�<��;�I_�j0�D4���pG�ZUdG�wv�Wz'X<��2��Ŕ�F$uK�cS;*�����ٻO�}�bY_+��tK
$]����q�mm�Ţ���orR����x�7�t|�V���o�yV����Z�5��𬗳jL�����\�����=5��:�Jb���#��b����C@�T��rvm�E-mIYB�>�+�5V�9�Nަ�rBޢi�G.\�B��1!Y|���\5�0����mW<���W��}_}��ᶞx��Kڐ���7�=/�݅	�x����"��05�`Ә��z�B�tN����]z�\H����w�����z���.|%=�is�;"�R���n����az�xT�	[Xj2����'AKw��LKnM��s�ﻫK�ʄ��؟��[��卢�T����]��`&��ͻt��]�p&o[�D9�&u��67�͸��l��r�)#'N+pW9`�uݜ7�p�5�>��rĭ"��+k�P�-eAZ��f�:��N�Z�_4ijR�$��y��ts��٨�!�'<=�r:T�G��>����hE�[sּ�y�裶Bn��Y�:�9x�3K$�c�]�s�aC҉z.R�}��O���ށ�*�&��$��m)���/w�����>|�H�ѝ;��-;r�|�KՏ��ĳcX��ү���^ϟ|f\����Q��	� ڒ�L��F��R��][����qs����Ic0�� ѺPJ��`�i[5ܩ\� Y;�E�������
/犂�8���qj�w�U�r��d�P�Kz���;�E=����螏i�N�{]EdE�F�O]�<���r���M=�X��1Xܾ�/��N+���x����ot�����X��=�nf������r�z��l+��\��7��f�%�=�rl�zs/v��Sf<�&�N�#$���ӌ��E�t�[�� >�P���z�P�)������Ѣ��@Š���UV��X˶
5UP��K4Plf�h�@P�mA��N�AK��QE1!�v�P@�QI6ɤ��tLV�)M%1@�e����@[U1	i�Q�@QKM	% UPhҔ��UQUTI@D�U%+Eh���"�����N�m�jb�Z)���)H�"h"hX�i����ulӥ�И��F����"����I�����j���"�����R��D�� ��i
�
B��hJti�$)
P��)
�
Z����h
����B�����Ώ�n���}� m��G*��Zx���7��r�j-������73��9�yK{���T��uq���:}���:TR�c�)[4ak��׌�S5'U��R�ve���2Y��"0��'j�ژ��,�Fi`>uJ��>�A�٭�Z9�h,R����u�m!�ۘ%.�ۺt�cD�}����X��uC-������YC�Oȹ�y����!��Ǣe�Ü�D��$W�-����酦/�N+�',O/��Cf(s��**�ڂ_Gpo˪ �|���l��%�XX�!36>�N���4�s���1G�
��WikH,�_�9�����d������U;Oӊa`Ob�_SO d:��{������gަ�]P����Yi�}̕�uƅ��⾰��`\]8��]~ S��B�yW75������2��gV�}�/�V���!�Ws;qU��>u����b�|9��;Z�ۧ��I��s����#�1��D.T����I�t�>�W�L�RX�m�flE��*Q&�z|S�ٲ��WH|©�~gG�g|��b�
�e����RA��ˁ�5�T"�����#2�c�������LTFq�1oY�U�	Ȧ֍8e!��{�-��m�A���-�^�wW��E����%�w�V�Jʹ���[HH2Cs2�M}�8v�v����Q�C(9:|+�ǈ`��m�7f�������
|�Ƅj�wE%Zw&L��<��X|��Gb9���<>��:�!�ܩf�9T�R�N�_F9Y�i�t�c@�5��M�..���xgBu�M�w��R��!oX�E\�4��������d@ި���PL`j�L-Ψ!�W�{\�g��Mȵ�L8�;5�bk+�f��
s&�J�ț��W�j	Bs4*�t>����;k��'��q���Zԃ|�5ktqք�c �n�L�k��q�h�y^'�`�.LlT}]�=o�a��G��������&Jn@�pxE1ά:��r�T
=��9N���KGh���wYd�5�yp����s�&�n\�����ќ >?�b���11��xv�Ӈ���1�Y�GE)�1q�����l!q�O�2:E}na��w��ۜ3,�F���P^\%9��^�y�ڰ��&;��0�A��ۨC�F��/T�sB�e�]׷Nw��_ux�]���&�Ӏf:��ؾUE�������X������
ɰ�, {'v��X��!�&f�{��4ӥ�Ɲ�7�-6�[5ou�O�ԭ���t���l�o�7�6$W�����w�_I�5�Y5-DN�n��g�9��'��15kZ�Eh�ϕ�%(�T��B�1/��m�$�#\��Jl󧽶�%�vj����S��tjr�o��
| �'�@�t���W�@�s��SKU�M�nl
�X��ֲ1U|�YL�����T��x�U���_�/r��Ȳ������[J}���8lc�yˣq�r�X�_�q=i+�;G��l��C��T�d��]��L�G�[�e\LT��o���C�3���������.2����B1�������9D�fp	��	&$����-T���Ĵb��gH����ml��~���:'��[S�^�K7��0f6 J@�.R2O�3���%J���VS���Z��ݥ���X�վT:�L@��k�  �G��GA��<y�U8������*s���졢�JE7��f��	��lM��hR�&\ќ��(�;ǅ4f��hO$�4��wt��{����+�Wzt��f8C��J��
��ّq.���"'X�ap��0m�2�s�.�D����F�}��C�S¤�D$��s�MVy�*����b�o����=[�;�WH��'0��:�أ�&���sq5��9�M��x��ͩ-Tk0�<�]`ja�sB[�)�sdM_�j{*u�Դx�݁����G2u^�wt���,�uuN�<�~�8hB���m\Q�2_`�0��(��Q�\��^#�k*f�:����CLoK[�*'<��1p���	��y�`p��񡛱ث�o��|gTU~�D`�Ug+���A��@��c�]r�	��Y�N���-mt+(^Y�|�>��� "���b���[B�o�'����;���~��
�R��Ǐ��K�zu�1<G%٫ċsT����b��T��G�٢��T.:���AJ�h4!�ΔKC��%; ����E77d��ՙ�u3�i� d	gY��یU��/hVM�%�~\��m�&*������4P�F��@vN��GK�f*v�[���u�jS�;��F�K�� �E[Vq/qź��X���Q��Gxd�}�U��y�#!ܦ{"�p|_	t�Zᶤ��1s�;��������(6�^��ɐ�F5Vk��2���p��t��s �Sy�}���CՈ�+
�� �Cy�2�� 9��D?��{=����̛��-)PV�^�c�H���C���Նќ@�#� x|���!t��<n���}ް%ТY5�M��]^M<`d3��ư*	�%ެ�m��,�VӜk%��OǹS�e��V��{#��M�	��6:���(nb�5'KhZT��冏>�.\��H)ni��苌g;�p�;f-���q`W|��W6X�<�s��K�;K�|1� k���F�6�۲1��+�ft�8ƐR* 7���j^�/)t��"����5�p'-�f0�Zq9�Vڡ���rH�}BM�޶������R}� ��ɋ��\2�9��?G	;AZ��&1�I��(�w�p�Jq���1t6���׬,ڢ�L��ā4)7V����GoY\�~m������1�s�'F��뙹�����o��S�/���=��j��X�B�s6�[]u�ߑ�S�N<���~�(����uU���4�Fhm�9`Ls�r8Տ���٭��c�%1J��*���7��J�vDs�_]�|�E�@
���c/�s8�� +��ڃ�b�5疩�ۜ(W{v;T7۳��:���G��ѫ����za��18�g5�1+f�nb�F��&0C��b���wهg5u{f(R���?{��_b�*y�ʃ>����3���?f�w?��1F�(b3a�ۻ�2ww
�& �P�a��깬7NX"�
~��|���@s1��w����̴M������@U�桴�+}��=�[��pr�y/Ww\`��T��o#�ٛ�.r���>� ��h��o�m�g�b�GI��eǰJ��R��m`��v��ʛ7"�DYMɗ��G��ޗEQ�9#e���ʻ�3gN�d&��Xl��]�5�33��y�D�����p��W� �]g�qt��l�o�cyW75��};.{㯪b��}e��W�NUpѹ��Ʋ�wE�$�h�A����{��(t.k~�Ϻ`�S��R�R�J�) ���w�&j���L�êt|�[<	<N�t=Υ�Hp�6V�z�uԃ�`�q�8�pZf��v����2�柘ڄ���Sl��jС��DA����9�z�q����w�I�X6���L�3p�W�JPc��]�w��=q�����s,�јp�R
w��������``	;)��@(D������tcN��z�'�� v�<w2�;� ��LTa�(zh@hFF&�zXU5���D@��=.>���k��ۂ4a�XK�!��wPgG%�X�u�)DA�{�$iFy�(N9��
��K����1[�)d�'�wE��`�'t#����U�U*qgW��~�k�u��@N�31:U{Z���Wܺ`��JS&M��yC�@)}�cϖ^Ƌ<�R��3��{��Rx4<g�Wc���>Q]'�rn�P��wW�&�+gH�#�M�ˁ�'�`s�Ngp]_�$�ќ��8�1�:�I�Ǳ<� ��V7c�ʓ8�k��M{����tXm)�w0(��Ohf`�|V%���#���ʠ�u�OLyn65�N�)�g��X~��Q�yp������ɦ��;m]h�.�}w�a4�����V����t*�11�k�
���1q���l!{��#:EE���w�����@3/bf�?-����f#��X�WڬH+�4����H1W�P���Q�o��O���&n�p�[U.[�y��l���y�B�\���*��_e|�V;�������|�(,NՌ����e92��@q�]y�2��[t��E���)�������U���>;��s�ȕX�)w2u�IͪP. j�Db�������ｱ�<�ƶ���PKD���x/`�]��c��5s���a�;`b�yˣi�eg�����B��r�K7]$���"�z*f��}/t]*mp�ͮ�9jhB�r���:C2�MT=
o�ٶ�	[����e֒'uX�j~dh��SJ�$�w������Wz�F/�r�l�8�?�j9�'->w7��e�m\vڔn }���	H�����[�]+�9u�OVg�ȫfN��r��v/����7ʶ�Eۢng�}�W#ŝkq*�D㜝��ryn^�t36���)b�Va1il̬{y4� NN����:�=�ۙn�����ޥD�M��t *�ݷ]R��5gR�t�qp9psd'���J��vj�%�Xų�{ǟ�'@o�0S�)䗖� V�dtSǞPU8�V\ �n
mP9�yN�^��s��d���y6M�p�D�BIB��J�$09��]�$�K(�p��^8Ⴃ^����Z�R�mr,�mv�~'�����d3i$-o�\!���l�oTls�L�Xs�H���+�-�ޒ)�Rb�I;,�9��wTd7&�
q��鞭����9�YT_�3�P;f*V�`,�4!�u�Wt!2�|ܰ�/��vPX�|{�fO��{*�R"0CVr�(2>Y�H��^f��Z���#��f�.�FϽ׾}�D��rA���Z�(V�zhS� O:Ǹ��\�Q{�
�R��#jS��\+1ۡ�9�ξL���@C�X��{�E��PF_����d��WYU�S���V�z�;�s;�c�� ���on;#�k����u_m�f�Z��fu���OS�hϭ����+sY�s�乞��=�Dj��:���41S��F3��
>�:'�L\G�<4��U����i�b͡57>]���W(P�z����J��l�>1���q1�ar�8�쳶D���r��T�)9t�92�H���9+��i9�-Q�8����s�*��R���oo�����қ.��r!%Cڅ���v:�&�5��u�s�Q�u�Fz�x[i�qB�"���g�e�싼X�w)�ϩ��\�����ZԀ�z�,�y�t�}f �.6g����━
��n�dk��0i��}9=�|.)�qr5ւO����S�@�QH�'��������Rixt9VP�f�6ޙz�a"*�G��d�=�w`�iz�zn1�!���v6rJD�z"O��xHnu����ն֙OyH��/&]L��㳶��=��L0�� FStEƟ���E9Dq� 7����=��S�5��
iF�@p&tD=;ʴ<��� ��Ӑ�ƈ���];�d\*��O]���3*h�M�P0 �	d�u�e�(u��v��E�"�-7T�_����ՔM�����z���%�:<��f�O�Py���D9��ۮ%�Ʒ������U���wUbFp~��X�p}
^g*��}�sU�)մn(�5�D���B�^�C�wd�"9����KR�]�p�P��4��f��,�Ϲ�9*��ƾ;6�un�����*�k��{Bo5��R�)7_W2�NU#R�����]K��M�F�}��mp�ML���N���ӽ���i���"�:���B�-�;Ȇ�Ar���5}�ѣ�_ή�l�8��(c!��j-ӃD���M���	��d�$�y�7ѻ�:�$ᵧ�H�2t���k���lGo*�<��� ���[�92O��wR�딇�{;�C2�A[Ź��Z�2wU�����4�x�~Ney�5X�W3�e��&��Q��r	���@�~�-֘���6��X6�����d�&��B
fl}��s9���R�]��:�4�#��j��[�9�t{�
��Z�����xT>ma�*��|�~O d:��z�,]���P���T�!����߻O�ە�mR*�����$���qt��t5�O᐀r�q�l;�%HM��i������\4n5��5�C��\I�D�_j5�.�JN{ev��+�x�ڼ\��L��wP�O���5~q�nU)���G���<	<��+ܡU�]Wv�y�a�I��G[�"�9(>68K3P��ӐԖ^���P��bʛeƜ�BRAn�:��\�b�A���) 1���-���L�2�OҊXq�]�w�r4�^�P�1u�m�YC/�Vw;*�h���?0vy��"��		R���g��']Ĉ�>dM�>�:�a�;7�a���tՒr���'����j6��fE,��y3I:�t�%����2��p�ף����E
�b�Q-D�`��j
�թlXԘ^�5��{C��F�97����f+�܌�]9��%� �h����]�
��n	�;�k�V�pmnb�l�D��a�`6�Y�y�`���L�Y�,��q��	Z8��
�( �|ؙ��z�,GR�Ah�Xk������
�0����7A��u���-��Ga�GP�g��x�$�J��@�}S�I#L�l5�
I�ʇ�,D{NR[��u�F&6��CE[�L���Z�� ���K:�NA:"��V�R�C��a��7mg|d4��OE����S�Q�Sd�IPq!��Mҧ��:I�wyq�z]��5�&�Y_]��4A�?���G�z0k�������2��� �ҭOn�6.�i��a�tި��Yd�E������y��KS�ͥl!Pu��i������g��+2H�M7'Ej�s��.�.����F4��S �3!���J���.�4��(ʨYƭN�-v�+�ۢ��������g#!U-N-�Re�����&T^dQ�WIT-�YV�Q�vrkW�Et\ʵh��s�L�z9j�&��kkJ�2�sC��-��f=�0��ʲ(;�$��Xg,�cݣp�����N��)�ASL�^gZӘ�
���Y��dU���j�`<������@v�;��c{n�s�V��H����e��;;���N�F���'~�����_�M�����{Ju���R&e�!�+�89�ʔ��ܖy,����u�H�qۨ�!��S�vl3�x%�t��G(����e/���X�v�������j�P{%��C[�Y}K�w%�'�/�n���n�T)�._pœd���u��z��G'y(6pI��9����Kr�Qg͗e�Ih�=��lQK����,���vf^Y���=���5F�e��R��q�W]XTS�%�%>[�>2��=4h��W	 �uR=QAݛCo�2��X�&]�\��2��S�M�Ep9�Fo(����C��}�ܗF��Rfar�fD�jd�et@ �u�̼'K a�f
�1�C��8��ׯ-cH���>q]h��էMƴ��<��ט?tlJ�^䚯�ɧZ�N`��_�c!�;tk"�҂��V1h���O�%�\�]��
���f���`��B�H�]�I�+�����!�󹀣"+��f�OC�[o�[�lNɉ����#��'�f�͙�/v>�AHsgRK��|�m19b�㜆��k$���=J�O�<TN�ث�D� ��m�]�H�9��ξ��7}5PsL�۽�nMI�G0�P��B��BKq���ji�(������?}������Ͽ��CEE-M4�A@DP����0R�ґ+@QI��	E����4�5EP$T�IB�R�14�.�(DV��CE-#C24P�J4�U	AB�д	T4�Z�IE-JLM$U)C4ZGE4&�EU4�@U	MP��RSLE4�4�,ED%N�JQQQ@�E+2�DT�4�KM����"SBPRP3N�E4UE%R�@Q��i��)H���JV��
hB�*� h���
�у�>��/%Y�ى�w{�d�r�8�͈��ĝ�-	=���
O��l�R���Q�j ��9���]�/־�7�]+�:%���xW��}Z)WY:���%Q�A����Ph�C��l����
9�K�:�sy���a�G�w�| �%�?����S�t����=�|�O��9�����]���{̽�����#�b$������/#�y�Bu?e�>�����	Oq�d��_�@F�h`��2���<����{�C�|��r>���ۨJ��uw��.>Qd,^^��s�ww�D���1򺏅�r^K���;���g�}ۨ���w6�y�C�z����M<���|{���wu	|��uK��r{�?��):9����a��>|�?w����������C�>��E�����G'������zM�U'���w ���s�0�#�R��y���M&�׵��>ƃO�?q��CC�������wr����s|��cu��|��
g!�����|G�}�}��pS���|�!s��u�7y�>��}��䝟�|��!)�O�y�G�>Oq�J������c�r{=��׹i���=�p#�G}�6>�?}""�!��3����Q��|�#���D ��LG���@K�?���?e���8c��nO�tw�c���*��NC��/z�|�i�]�?�w��~������/[) ���"������������\�]n&��F���8H�F��������>�����9�Q�9	T���ܾ��B^c�x��?K�(<�?e���>��pF�eݟ?�w܅�h������&�G����u���>e%Cs{�T��b>����yLP���K��s��Γ�N�B��}��>��:�}�����O ����8u	O�}�]����U=�c�C�gX9��r9~���i4�?��n��߿���{�/���+�3=��DCDG����hu�θ�{����:�y�O���~�G���>�s�]'��~��{�T�F����? �7׬�S�?nO|�S��S�z�c�:���������者ſi�jsz�|�h����+-:��=�t�/G��t�?���}<��UK�cy��9	}�����ʟ%�������\����#�%��T~�^C��������;󛿒���2�x &���{v�[��]�]�B�Wvb�Y휸����a�
�Z܆�i�
Q��c�\ק��������$4)�'w��	�ŀ�v�5Ɍ��;�CP�͌l���pƚϯoz}`��Ɣ�h1��̾U4�=�8��zs�&�S;:�ο�K��O�={�]e��:���x�/[.�F��}��!�����w	l�a��u��{'#�{�_<��u>G�r<����w	A�<㯲~����:��
��� G��k���2/���Bwk���M.���O$�[<�>���r_/���~�����p�|�� }�h������J%�~��V"8F���#�~]Q�Hj��Ur��'�r�w��9�h;�?a��^��3��i4��=�K�#GüuW�N޷Pu�w��O�y����F��|�}�?e�������|��#�`p7yu�ֹ��U�k�7���:\��o1���y˗��x'��	O����������PP~�'�n�/�������4h4�<�<����Q�%?eݝ{���F��WPȮ���񌎜�m
�io���M�?#��_�'�y��4k��ϞpNC������'q��i�{O=�w�^�c�#N�l��5�������y��-�����=�D!XN{3�>�q{�)�;wV7�N��|���~�����t?��%�ν�{���9/�޸���C^G��{�>�S�]�y�=��#O�{�N��hz����:��<�k�u/#��~����^N|@E�&=�i�9z����bGу������9�;��!����;>����r� �<��O��O#�y�:��`ѽ�s�>����~7�N�>ƓG����^@u��:����}dm���E�nX��h�b"D|oA����t<�	N���ݗ�߲��Or�'ې����A�0�|��y��Q�J��8y'��NO��=�@QA�=�3�%�-�|��ￂ�f�~t���t����_!UDQ����'�����>~�Q�%?��g��~A�K��:?���~=d�:�e�r{��2PF������|���~��?X��A(/���O�1B(G�i[>�4��Y��A�X���~��>���F�-.%�p����x�o���NG�>�#�J|��|�p���r�ޱ�=_d�$�w��`�ױ�'�u�i�?��_���]���VU��p�@�!��
�^���l��>s����v,J�He��P�]@R96�r.mA�!8v�y.1;(-x-��8��4Y���R�t��*T�8��u�����B;?
�\@N�8�6��V6	]�5��D�c���F��i��������¼���sK}�Y#�#�nb(A|����.{�Or��������uO�`��:�T���u�G �'f���������?����)�����>����y�I��1���<����?�S75y��:��:c�#��+����4�w]t��/����=���r��z��a�o���O��?e���>�d��?d����h���y]�rg��4}��p�|�;�����{���}���-�[�Ǿ!��G�D��=fG��䜟��|?��h����:?��	y�����{�א�F�]q}�O��y=���w	TGϾq;�������%�O����}�����?y|�ojgBCoˁ��}���}�"�0} G�HP��\�����&���y�����=����]���w��Е@~�����%���/���=�������} }�8F{���!#�f�nXY�c��������������?Aɥ������{̝@y~I��:�����5����{HS��|����s�����]�����p��u��q��$�MC�{&>�1"!���b��M_�������^|�i���:��?G!(���y��������'*M���3B^a�:yë���y~�:�o��N���^e����p���>,�ǽ_}�>���}�נ��jO�ߪ�>��߻�=J<%�:~ϯ�x�~��_����>T���r�u����i�����i9>G%��<��r9''��7P�KE6=��r�'gx��>^Q�˩�}��&~�O@�0�Do���fw[��DE�">� �C���"a��s�ʟ�|�@h��n^����{��5�~�{��*B�ߍ����/Q�27S��/���;���?j��Q� |Ԩ��Gm/,�F<b�Ew��A�a��G�j�����r>���C�!)�>s�:NG�~� >~�U>ï$�?����45�?�}�~@r4��{��y�^@y��p���"��������{4�#�[�����Bӷδ<��� ��ҙ�m��T̀O�.,Sr��ы��:��J�7ճ��`�Uh#eLB��·(f�13c�X6���+Rt��Yt��M��g��<%���J���\�H��X�x;�+~�g;�2@=�3m�Q�J���X��[9ӹ�}vOH��05��z�pPi7���⪾��ɐ�XWSg�8 GL�)lп�L1�
;O�a'h!�9j�8Lc'h�)�����^�����=$_+�:��+LN���Bs��K�{�]V+K��!��FiN���S"����>u~f�'�n���)�Pt�z�QW]Á����e�]�2Npm*�8`�nX^B3Cm��y�9*���;6�V�7���@�v��s�7����!J���'�����7� +_�͌�#i1�h�j�̭'tHkq�5��������a߼:����釦/��s�uLJͨ�1�X9V>]�rA���D�.OS3�+���N����>ep�ڞ�]|Iw�W'\�k�e(�z]�=[�s63T<]:�@�>�4c���P�����8�x`
�%�"����ܲ����"ZL^�eE��2��y�~��r�f���Y�f�Q_XGUs>��q�
�R�\X멫̂i<���YŵZ�k�-��?g�[���ڽ���Tr  �$��&� �lx"{(�*���kC$�<+[5y�v�*co�9��
�2JF�"a�+�OC�2w�h4[��W]�=�B2%֜�:��]�Z�s�W�Z�W-��Ѡq0�V�p�v�º�����K�3x��+�n}�49�������%��p�W�ﾈ'x�\k�0`o}�Uã���0B	�'p���Ҧ7>����\�������g@ռ�v�@=ݔ�J�Сn!7�n"�G#G#�	Fj�zr��ӣ�3�M\1pT�/ l�{4�LAUn�m.�fH!�6�:|򘸊��fժ�j����;�9z�'��W ڱ����X�z��fH����/�� ttW �� GW{��o��z�s�Up^�FJ
������>X&z�t��-�\O�T���(o�@�$@]Q5��©�Έ�kO�w����ԐYݲ+�.�����`cP���;���!�4� �fy�(N9��.���.f�.�̫�������wʡ�Pۮ�8#�uL�U[���D.4v~9�X]�K%�[�a��s��I�'Q�/K�܄������2d��p� 4R��cϒ�tg���2!�ʓ*N���׾��f���3�)i�=�}]ח!'wF.1�̚n\�T�u��S�x%Ud���k���? �L-����L8�<j��<LX���~��w���";]��Y~r�r�u��ɤY{���[��k;w��*����I|��N(���Kţc�u����#���]��1��?�7NZ�h��F#�����,r��o�u9:т⊋����gn���.Iv�k����̑s��Z��;����l�	�;]B7�o�#��۔���B=n+M�,ۜ<�'8d�� �Ra�І�(1����@Ѹ0[ ���-β��o9=���n������$rҘ�n�q�6�N�eչ9a��E��Թ����]pٙ��!�e�{\"��p���d�L�{�h�d��ڱ����_FۊkG0���o��u@,=ι��>�pw�6}�]{^}��TV)l���C�ի�_lH����_�^饱U���G&끊�TA�K.�e3ʚ����᳢؝�w'�ҟR��GoDN����@�P:K�m{�ˉ����>x���ޫ���W6�v���s�zm�*�W���<I��|��m*���w�������'�����ʾ�P��#;�8�!��N�Î�P��>����
��G�B��+�#�8�J�y;��|9Nn_D��u�VS��t��`�4�N�\�" L�2:�;s�����4x��y�*l�.��ԺH�9��&��M�n��'��h�^���Д��ˮz��P��C��yj�����V�[Al���]�R��&�U��@�m.�ѧq���4d��P���	���q���2��!	�p�+cXKs��/m��z
NV����[�K*�S��t��G�y�=�2+Ի/��R�L�7�^q�.��_W�ܝ᤯x;��4������0�.��1���.m���� ���fF5ϖjkw��4�z���8��D�ޱ�å@�A�k0��o2%�\4��zώQ��Zp�-�_��ڙ�Vo����k�9.�V�Q������4��X.�^���Pfw���]�G��[��x&)Y�����:6�)�@�_`o����mU:��?���^��\6�1;���������x\��L�B�|�U�&)�hEk�OP6;�
r^�lP�v8��ƴs��}e�y[\:�xn9:���1:�l7�e��F�0���8��Q�/�w�7�ِ�7� ͽ�Y�5ȁ�%�f۪�o�U��vP�q缪Fg�oVi]%���@,[~Dܜ�>��(	[\>�癁�y��ePLVe|�9�r��7��׬���5ꚴ/�b��QP[�i�x�E�řTW Tb�e�̑��7ny��n�����S��0��1�&����@r����'�u�I�'�n�}���ɭv
n��2� � �>rǍm�~��Q���
Fy�����oә�+&KAR�Do�R��:��ل�s�.8+\�"�7��N�DfM��m�>��%:�ͣnG[B6�ys��� �2BcI���YW����@���t̫s�+�����)egTҺl_�ﾯ������p3yIh��}��}�;����K|&���$�+�#�j?�R�&(_f�Q�Io�#$w|�6rIf6� ��c�C�%���l�j@��O vΊ�9We��z�Ј��qFt�qbۊ�2�a��L0��k�#j-�#.բ��gA��Q��4�m�N�v�'�6���9�9��!i��u��m��oeiϓ��V�A���xhm�o^��ۚ��7���m��D
��[4.)L1���~K䝠�|�,��1v���1���EuM��y��o;k9�ܑX@Q�ȿ��i:��v�/�Z�
���Oł��;�/���f.���T�y�3,yD`�1�D)�h=ht5�T{V Я\2�����Q�	�E����!�Ֆ�rUrn0���Ќ�ۇ#	�uJ����;6�ع�;���w[P6t�)�F�L`���갭r���(I���rf����B��2���h�3�2��U����\uH����7�|����5��w�o���^��0v���ďt5]��+�Q���Y":�`���9��lNb�f^�͇�9��W�poi��g�՗섑ɻ t�.�9{W/����;4s1��R�d㷒L�"��q��.�D�\��0�2�x��C�ʈ���_}_G�a����;>�L`��'t���0����]|Iw�}���9� �LX�̦�]*�Sˮ�N�j暱��a�������{�
�ß8��(	��|�+{�f��czK�u�erހ�Tk=�����Wkj�Qg	[e}`i�������+�T���{���� 1�@���\����b:��u�m��C��s;qQ� �_pT2o�v����n��`ڬ@����,C���v�0�>�
�`��N�3�c:V��ʺ�[<	=~\V�v�k�U��,=��7���B*"OF(έv��K/�?1�	��4ˬ�����z8����E$��W<+tN��A�~
x%1$�3��}4�0_=v��F��D^��{�|��«��&􏭽�#��K* :��P ���ryT���!u)u�t�Mt(�t�l*�v��5]���q<nR����5�"P@�e*@�~���s[~4�ӑ�t��n�cݍ�#C����y�A�M|���ռ�&C� ��#L�:�-����w0�p�&��$���rs|�6����;���ʞfF!�����r*s27f�V섻6�^��P�u�/��8�L�Qt�;�j��Cz�#f��X�Iomf@_�}7#]y�P�A��Rg}�Xס�a],��}��U��2]�҆8fU��|'��f�PɨM�� :��a�������.=���r۸M�t��w�|޽5� z�Ԟ�����EBR�2m7@s��
<"�9�X�f��x�N�A����
cE���?]R��u�i�v�I�٫��Kn\��}i�V�n�3�	y��<tp�\~�=�1�W��3���7�i��U뮐r5a��jB?6'#�!�ل�r��6�m��9�'jO���Rگqb1A�.-����*���:��������,�7S�<̈8z�ً���#7%i�3]����/}ơ@��*�ex�>�šY:��@�c�CUC�L1��"���+�����E������]K�͵�Ό*wϛ�3U�8%� V��x����i�M���u��}����a5+�M�<96��-0��.�L�ۊ�]1qJ@�G&��07�Ȗ]��2�)��lD�=|�\��$�E�cK�C0�<gIAᾠP��s���E�,o���^w��^���o�iAdCjN��c�#�=�]��=)�(�h�jr�mt�`�`��ͱ���&��57C�]1������Z��Q�L�.R=DTd������Hٛ6T��u�|z��e���^�[YA��*�]g�A��U�E�&��d��e���7��K��)���P�z���	��f�
|�V�f.g�K���{һ��՚��I��7�Y����MB�����i��]�RA�;8]���ǳR]��TH�u������q.��Z�WO����!���ׄ�A)]JMY�f*CE�W��|P%+�3���z��%��c`ji��ɲI(�uS�J9p�.�!��
S�>�&�^��F��L���.ّ	r�M�O�����Hی��mW[�>^���M�Z(P��uuJ�Yh)K]ӶF�ړ[�*��U�Kt�� ��:Fջ�e�7$9�ޠ��V�ďp��DU��m�b�����z����E�'���ثYN_�\71�5*�T|�-���q
���	g�͔���tQd�
w&�)���)m�WՙWG�6*4��b�	���nQ����꺰��A)f�'V�R�ǎ[�˯ic�0�����ղ���8����b��hԫ�8�EV��}
��Jb�eW]�K�Ru�o4�A����)K��˱\RRʆ�+j�!�O&efk�}pA�Q
QU�dP�=ڥ�y2�欴	��/!��Y�	=*X6�B5%���@����\��L�Q.�h��l����L�a��h�S� �J�q7Y[��Z�o{3-ŵr��A��v�TJ�f�b��b��.u����6P��F�bf�W��wg7$�B��5��DkiÙ���w���s�v��H��5�4���a�]��c�����S�$��ܗN[κN���QqF�n
[\�ƽ�{�WW��nE��g�y�w��\�o"4L�X�y�Z�@H!��2mq�.�u<�²D�n�<q�<M+P�o,�e�n��B��ӝ���ێ�HG�IM��Lus{δ����,5%X�ô�����.H�>VIXF�Gz!�[6�S���7�Zagtn�O����S���fc�ȃ��ؿP���C����b����vA�����CN9k͆���G� ��m��fK�������闪,/�+2s���jP�g��{����v:���>�ۋ��m��a���b7�X�u!��S�Ʌ�as��F�M��.�*�#�2t�YW0!���x�F�����ܝ!	W�K ��������������	wOtޒq�.���]%��Ů�-��V\���>'7u�s��f$8̺Ygd�-�s+	���;M�dw��Xû:i1cx�e"ڝn�[���ˣ;vQ�y��5��c�|u!�k�R�(�����cQ��s��Ӱ�=�[�ԝ+��M����hc��BtS�d�ʧ���5�:�ԀK��S;.ui\���M�5.��_WC0L�����_
__P�1	TP%@P�QR�UP���h�
J
(bj$(��������&���(�����J
J����JR�(*����iJ�����Jh�$"�i���" i���I��4�����(b�K�hMhĴQCE�!T4�Q�
���֊�(bZ)�N���� ��F������)�����DE4�U�&�P����dt�)K@�P4UP�M�P��9:1% �KACKR4�T�<�
QBD4U%�SA
P���s��)��|�	>��.]Ѱ�����op�)w�y[���Eۃ�=Kd���+4��Ce�]��������ꯪvV�J�Ͻ[.�g������?]|7@�$�Eh�}���Hxsش�D��k�"��R��h΂���C;pX�p�N��ö������%* 2�����}	�J�s;�o]��M�֚��5,�征��mۀ��1�1sͯ+�@>�֩���(�-'ҴOu<Ut����y]��ǳԑ�3�8^�i�#m�X��������M�ٹ�"��na̗�6xED���ρ|k�
�.��1��%t���X����O?��C�7D:�$.��`�H�:�XL������	���p=�/�&���E�����:��������͐�1���}΁�4��X-E�.���;��������fR��"��H����9`���>P*9�=��ug �Q�4:�؏��Y������e={�J����yU��Z�3VX��e3"7�Ԉ�A=��|o�P����Ef�1��!6�MYqF��3_^^���rt1c�bw>����eAk���W�-K���y��
94FD�@r9�n1�fV���)����f�9D1s��&�1[�I�ڽ�����g+.���4�/yTs�z���+��0l�'�j�[O`���Ⱦ��Kc�$�Y�4����5[YhB���Bz�1o菾���WQg��/ya��o�xޛ�d'M�W�u7�}BY�m����k:B��dmlLt(����������`0�N\_^��Q-	n�H}7�+k��\�09S�ʼ+s�<u��c�oR*�n8{z�\j����
����1N�B���`�t9_ֻ�5��t�U=k��w������U�i�S�m�Ϭ���8���m/qH�T�Nx�͉��7V�x{6��N�dk��2�����Mʺ��Q�G�=F~�[t"p��S��o������d��E�vt���Y�� <=�������j�e� ��/uM]�X�r%�g��3t�M}Fx�U���2�a�S.9�@����e���N��:�FC0���wکI�D7qd���j�T�����δ<�n�?
�Xz�����|.��s�[u{)c��yG=N]�B���e +�5|{SN*�ˠ`�{O��I���-Sɳ�-����3j�g05�J]^4���Р����]:<����������y��3���z�)����Aeb䶁�qmwΗ��.b+:W�9gW)�k�~��B�c���I�֒/���E�00��ݫ�<|�*+���8n�n�#��3i^��Cc��.,R��l�A���9�\��֎��(d���q����o'�����4�(�-��܍�>s�Bn���`k�"�P�1�3>g�'�F�]Js@U���R#��]�Nj(l��������"����M�r,���P����B�+�䎞��|��bc��T4l�u��eغ��� V*��sQ��١,V��ݗ��}��0�a���2~����V��2�o/��Zq:��TĪ�L�[�zs.�^6u_:��Ja���M�Q
����/����� �����)����7����8�i��~m�p��r~2mw�i�x�A@7�UA"&��ϩK`@,���Dv	�6�ZIص�����n�����H�����jQ~5)��1�e�x��7�dһ	��;��k.@X�W "�c Lo*���1r농kk�ƶ�v\�L	���"�҈���ȴ����"�lel��:�!�;�����So�ȵT���Bc��]�`���.P��u��)�CPV�v��K6�~C*9u��Ǒ�;��<�X/y�|�wmZ�[І�yު�=���.�ׇ$|:(��ݣ��si|�z����=(j�oc��.��Q#{÷����q8�ørL$�Cck)��n�6��ٺh-��wo'f����ʻo�#��L�RB��ɣ,�6O���G�} ���M��7(�i�(��JH!U�!ˁ`�EWM*��#������.3�OE#S&D��}C7�E=�>��P�;�,ڂ x�� ��Ϧ�!�pHۋ�� ��3��\�-�������wo]��J~��5�T@�4IJ��&05��ַ���wm�F�v�:YWqz�z��+�MZ^�3�MBn��V�*�bB`Ơ�`Psׁ̭�LD��m1����g�d�q�j�U�M���a[�`�ʪ�L1�M�F�z2j�MF4_OZ�c��?�C�^�ޙ��x?�t�	Jdɴ���
��i)�d���Ǵz��+@���cYF�
cE���|;��ʇ�-�t��6�:��E)��d��v�:�!� ��t6��Tp�����b���X#��{N,��.(U����;�:��g����+�,��"��0�ۆ�+M��m����v0��.�)0���%h��S��^���C�[u\q�p�O��s�t�f/��#7%i�3]����c�oO�����)(cNЧ����^-X�%]�jtn\tp� �ui����8q�`�����6�݄�v�^^n#�D�*�D�A%kW�6;/^��U�lXm�՘�ꕆ�܃miu��Z17k���s�{���&�UU}�}�3�7����zN�U�0c�cUUC���r��S�e����j� �ϔw 6�����oB�/v&��4�K���B��*��� &#y�21U|��L��u)��k�(�����+��N�l�`��>4ꉂ��DO�V����*��Ȩ�������zv@�Nt�M_n��-e������AK��":+Ø(T�.|.�^�뉊�7���m:b�^�/>�ހ��8k���m\>ϊ�F#l��&2���m*��K�y�;�v��l�v�]<��MvV	�R�J%��3�X�p�'n���F>�f6��
�������׮u3)�vZHz�3�z���R��pVS㺝�n#�̄%9�r� .�Z��ԫ#{$~����;i�l���v�GBB�v�Y�6�2n��SB'-L�Ν#/s���M�`͊v<gH�ih�~9�M����h�c�0�Ox-mS.�R7u��8B�3 ��zP����H��5�(�������<_o2$<5
���?Z��1�ƳV��
���͍�}k��nh:�J��}t�f�t�Ԝ�4�o葽4"�]�_f�Go,m�|(����X4�X�\���z:��`��i�ug8[oC�O@�v�<��}�[�Ђw qjrR�3�b�.*0�+׿���ﾏ�ySΤv���-Ç�s��
��4@���ڙ��m+f.�vy4+�<����1ھ
Sg�y��ݟ�-ک&C����3�
��*F�0F��B1�Q�PL5^/�m_:D�@g-WP����7�=i��tk��٫��AN��sB*R"�� ��l>#�����ǌҳ�0��2R��W`hT����٫��Crt1xꘝ�����T�ĥ{>��Ļ�w���dޕ��_?�Q,�� ��T(�c�����c���7U���ȼ��~^����Ϸw���pW_0s�}q}~?r%�-���u� ��>^}�B�ox�͚���=�36p�}CH����T�����M*�t���������X�2[�њ*^.@S�����u�#!ܦ{)��Ugu=6�(
�?N(�p_�/q�߻0 �'2)�����p��ٍ��5����a��� �>w=%T�\��@�b<nXI-�\�I�\�}�O4�El�L��ȑ�#�����K1��0W��ŞG�x�t'3�vŎ�A?*<����u�w��}<����
o�,����9�p}G¡}�o���w��o�u$l�r|l&��{	��^�_l�H��IC�^��vGku��q=���鼫H�v^�մ�ɡR��zc�308+��b]�[S�%�����"o\KW� T�N�G�G#QFx�qbۊ���\r5��H�����(��[+�>;Z#��]zAQ m�J�@�g�o����ZKvٌ�V����ߍd���@yz��g��W�����>��B�6�7(�\�P=�L[��2�9���� Qi*u��6îr���4,5<�['Sw�Qu�q��n�"$���q��[3M%X=�gx���e�ާw���W!�����ۮ%�X�Q�L7L}_)�tx_��h�}{�C��y��ҰM���S_eC����J�N#��`ip���b��o�x��zs���L�t�\�ą�����͌�u�n�����c�͈]�oN����`��61D�Q����5+E�Zv��N�!�e���󨗪ѭ�`0X�YG�y
=���������r��T��<P+���tU`�o���^�7�h���C�eOl��V��=w=��� ���ӝ�}����*��2��.�L�B ��0�ϊr�|����ε�Y�ګ+��pB��FΕuj����'�hE{����n���ƅe��������7���Y�]�'-&PrpHK4&q-��;Y7��n��n�^'��kI�5V's��bG^�׶7��/)�ޗ6L���˶�P�+x��o?}_W�U��Q2��'5��޽\u4�C��g�����<�Y�����23�x������#'�1��|M<����K����qi "�"��nkbS�����~^�v�9 q�����:� �Lܳ��h�B�WP�f��:�y��
�;N�3��LnD��]��cfBk{��{��3���t�9Զ��Dxr;	Fj!k��!�,�9��5��Ot�OU.ؤ�r]~�<<"��;���!�*�@�EH��"�Ƞ��O&�ur�;�E����,� ��[�O�9�!�ܩf�A�|g�� 4���+��9������N�	囙��W�-�:�%먜=�O͘�"T@�fFn3����N��	ίLk��3�b�j�'���cI��.[ȫ����Gq���؇e�z;�a�I�Y��FC㙰'�'��5
�J������\,�+)�]���d��;:	�گ|��ί��5�:��]wx?�NtC��(�T��ՄH}뭢�uL�YWg)����f�k�ʗ{�f�l�X�=!f��<�JF�|%�qj�G���V�_O���֦��p�5sj0�n��+��.Η����<�τ$*]1nK5�m�rX�'H���(�{�e��pUpp����J}�U휊H�a���_UW�j�ڞ��\�L����cv�ut�,F��v~<v�x�Lt�뎺Ww�C���Y-��9�jvw�s菾���v�6�ќ :�?�ኦ�U�:�^Á��Ʈ�����N��S�K�d>���=��{�OP-�@�u�CY�8s�r	���@�1η+�"��VC3v����c�s�^�5( ����e�S�9�hA��'��ޑ��N������5q�N��kLL�w���.'�&��1����p��Ӑ���s���Q�CLcvu�����[֐���@�t�,����jl�����Cl�cv�E�q�|����7}�P�T��z�z�X �L�%�]4�ʔ pӊ�:�dtD��v%��\)��"��m���yAK��� �9��@�.|>躮&*v����g�?����yX��pt�a`3���|�?t@�*�p
N���T���im�t�����q"/���4���p��8{Qo�'-��)}�`�_jb�8�*�B�:�E��*�!t/'���Z��}��<���̚�����M��[݇yuAW'��J����:���L������:��2�m�]7f��*5z�j��8\G#�)ʐ�u"�Xi-�&�����oѽ�;r;��3y�wmP�Ē��}�G���l�$��6��۩/6R��J�n'��ʇT����o ��h�j�R�R{�c��8�����ٺ����k��l`86����[7�{iv�X�����:��܄�B��r�S}���}�R\��o��q}��v���5w�ղ�3�:��S�,��눜�kFk���5�'=�^��V�������EgQGja�2�]�D�b�b9ۚ�����3s-Ob@f��P&�xk�m���.{S��X�%F�8f�q�x�dLs�y�5��4VJu��5�N,�sz��z�}��b���9΅��[�vӝ��j�}W�����coԳ4�y^��ma����3��V��/+�k�r�\~��7�[zU�A����T�0����=�1�M�T�Q�&ޭ�Qj^�{j�A�֭2�q΋�ܞ�fr���U���~�K:�R��^}�`}�;r�H�c���3���ym=���R�We�'�Ԉ/yTĩ^j��
u=JE��ݮ@�^��{t4�j;��<��72����o[��b��e��p��5ն3��{]�5���&{�8"�M,��,�23z�Zf�f�t*vL?*�{X�s�.����1��ka���,� �:v��&K��Z5�t�i����2Ǝx�z��rw��i��Nҫa���7�%W|@5`��\���ݤ��\�Z;60PS�	���R�$�!1�u�R�33�
9�1WAbɌ<b�鵵�u-4�U)�zJ3	pBE�ʘ-���x�
ސ �݋�΀����/L�Bǯw�����r��������Fx��f��Y���M�sV�a��&�5g�U@Ʉч��Y�#��+:�5�wo���#��EfK.qt�е��0�)݋�^/��L�[��	'{7������oEW�R,SG��-��ew&�7�����;w ��c-m���H�B���mf�f�vu��S��)QT-�L�l=�S_a�U�!F��˽�!4Ipd�D�v�R�f�+&ɷ��Vcx"��7�=若R���r������/㚨��Z���z�"rv�e%�{!]ۺ��q����N��kFb�"<&��Vp��ˮ9�j}:��;`=�Kgv��F�%��UϠ��g�|�ecŇdw��g�_>���XK�
��7ۦ�c��&�T�i������J����{z+�A���&I$Y�hx�r��x�2�T�M�G�^�#-;r�[4`Z�ISxOu�z2hCwP��2�]Si�]�����D�2�Ն3G|ի.`�*�0]U�mS��9
�갵"�g;K�ɳ�u����Gx:�h{\j��G��8�*-��N�ޖ.n�՛MZؔ8�*�`u���}�W4�=jd��d|!�`o9L��{��,�f;z��\�HLKxT�1y���&Xŷf¾WP��O�	ۗO(!M$nd�g�1����
��~��e A�0��8�G7V�/�7I�Y���#
+�+��o��WnKC�,7���z6�]���bZR�C�\���mdvH�Ļ�:Zư�����|�ij�P�DY}�j�r, UlWV+�u���}�U
p+;�G����R�7�p��Mޗq`��ύ�ُ�7Y�5Mv��Qj�dc�h�`"��Ƣ,�+�K�4�%�SX�"�m[��K�ّX3tD���Nc�ȓ`:�ʙ���wtܫ����dQnS�����,��73M�3�q�f��U���b��ٚJSh��n�����4��YS�܈;�tc���<t�:՝�d������r�]�]�N������$O\�����k�Rժ
�n�+��1_:��6R�q�&I,��G 蘪�q��գ��f��1'����jR�h#޼s�,pܜ��W���**�ZW�	Ԏl�2�΋�9C�U�Rmtc+P�_1�f.�/�;j��P�����4�P)%!J#CHGBR�7Y3%-MKM)Q4�@R5E14 Ҕ@P��M	�% R4��AH�HW- rWH4!IHPQ5PQ͆��Z�Z
�K`�P-PQM�5CEPJQE)T�t�-�˒��i�D�Ҧ����Xih"4��)�&��)��j��� �
�����󚀠yJF���M�.���(t�)j����)�����A�4s8yi��MkZR�
k���$/��v}맯�h\��1��Q�d� �wl�I_K3��GD$�4L����j�����;cy-�1c�ؐG��yՓ���������gc���r�ҵo�W�7�X��]X�te����ys�*q�y)�Hm���r&z�w:��X��|��Q���B��Ml��p1t�&�Y��qp��l�+/$�
���}]�������yx����28�5mޗrt��zl��t�;�Ww��Ng����/k�=��H�������ڷ�C��ev�g�J<�M��O��L3w��;G���I==�������iS5�%J�ɛ�W
�.y;�m�����������ϧ~f���q�t�!qs���E_=ܺ\����-1�.��/��2���盜�����^rA�p��6^�jwp�}��2�;��EDL�)�5�.���Z���jr&�Lr��q{��UB\����G"[�+�4��;�gY���X�nj��SQ=�5�u���U���mƻ�q�����:G�/t[�
�����RΗ�b�� � C�����WX���j�좴�
����*�(Xz7Q1�f��j���c��;�⭋L��M�u�N������^'/��ɵ�p���γ�"���]������f�Y���T�-�꯾���~���������cڶ`��d\���Ƥ����͵	];pa�s=�ά��:��s��~��ڽ5oڮNG���M��s<�.R����]&�
=<�؞=�z��ue^����Soj"R����z��C�H>�2qI>���>w�_vk짷�.������l�sW ���һ�׵��X���c�]�=G���w�����^�֛�~~_E�by�)�Z���$�WӰ��b���(���79��������T7�gko�/�o)�Ú��g {_��2�l-����P��M>������:�DHݭ���gfd��2�r���Q2�\R�k�����%���S�q��̀�y��v��ݷ�v7
��)���CKk���*��&�P�ц.����-���k�ڷ�):n��k�Zv�`o>�{�
��b����V��U�&�hsr��N��"M��F�Ocxeޚu� `��z��+�u��	�MK�0F;M��T*Q�{F}B�l�9��9�&��qZ��;p<�C� �h �ע��q}�&"2�;���^���;�M��҆�꼙�ɑ��ﾪ��C�=������=��q��'�3z��7!�/���;o;F�t���D�j6a�-f�[?_iI4��$�0TBo"�Ӑ�Z�	kq[t$~�2�Û�f�P�#�'�2ؾҒ�z|�l;�+���̃g���ۮc�WAÚɭ!�|6�
�5/�j1d�����vLR��4w!U���r%	ϭV���*����씽�6�ٖ��<����{䷻dNǼ�bU��jf�T�P���kF��uznv*�9UH�Obؼ�� [�\,�oy����*�{ҹk�4�$q�xo\�{�1j�5���v)0�-3)%��8�g=��W2�_ܟ=e��{�M���!<z�'�z�%1�\�g�/U��eDOp��;;S<�Խ}��u���xD�B�]/{�jt&e��~��Z�U��ʕ�tb����.������z���}���]@f���<��I�o[��q@�)6�d�1Xk����et��l��i8�-E��2�y�|�8����i�$���8kZ��-� �+�����Y�\�	y�����Ib6��k����$��W�v{�Yv��K=���¸����ꬿB����O];Ό�@�#�t�N�>�)���껡H\���Lҩ���.���n��OM^�|#�@�#���E�*�W��r.�17��V���hj��ƚ{|��T�0v��?}ӱ��ΛH�{��x�����om>������tr_�p��Ev��=)�1C+���
�3�d0֐�#i���+���ۉ�k��xc��ŕ�@%��Vz���>��+�B2C�������}�楐�:��rc���&�w4p-��䡼�#�{�F�{����.��*�.i���b�v��v�7��ݬþ
¸���F/v�h��uJv'���w9-�Cv���Y9�6BT�78k��L6bpD�b�yۚ�/� m����v%MGk<)��gTڪ���n�w�Q��ᚈmƻ����#�vD��϶��y<;ma�ƛ��>)��n��6V�S�s1:�اLg&F���V��]�!�K����SR(6�YB�؋�=�����tjE�m�
�÷��f��,�{ӡ��V>T��Z�%x�<<�T�p��OCV0��Ԟm����ϫ���狝%��h���-��3O�5i���p�[�u3��B�<�;Ut'u�9������^��nM��E��I�}ޭ����823OA�#���X���E/�k�m��Uȇ�7'$���N�_��i;��Y�qJۣmr��	��Y=��9��秓9���_g���,���j��W��|T��U����Ыs4?�^��->ϝ�W�����!�rh�V��zl�*!�1vm/�xfy�곑����3��������VuBkg���+�v��1��G~��I����=��sҪ߼o7��4��'�U򍲭F�qnM_t��F@�r����)ԗ�Q9���>�~^�=>�����+>2��_7�<u�<���}�o��H�MR�JWe�-k�;c����m�졎����޳�T����/�L�����l-��ӣ���0���rmG������C��ua�����:$.��fSerJ���5���"���2��ם@vh�Q7��߬Κ� q��7�>꘤��Rz��Z�2���­�UL��EGD:��̶\�m�qQ�{�r[���qGm�λ�}��E���n�eߡkq��V�ʉt�B�*���#OÞ�D�x��R,�e�V����q\�L-	A��ب.�D�ϸ��QЕ���W���	�q6�q���*�K��o��eƻ��&��!�@��ʜl�zA�2� �ɨ��j1f뵱�Q���4ۍw����ݽ������:�*\}W���7�m��Ȑ��t�G��Ok<�^ɂ��wEf����\�:�s���U���ھ�8z9G��7ƔO��}��ѕ�{��O8�uK����9�c�z��3�ue\k��E���U����V܁�s�0����֙=��7W�lr|�#\��{}��Ö�fTs�V����x�5�ov���;�Wюv>/�Z���<��}эl��X�Kde�*��X��y=�`��S�к1�E����ˤ���p��^���\v�O	��@�k-i�Բ��d���]Wn�v��:Te��TI���k+ξZ�PM]f
�NT����P�U���զ�ې5pˆV�x��d�x��Ч���L/���ͣ��ǒĭ���x��f��B-�okn��tb�;���}��Ga�Gw'�� ]p����G*�������I�&�Dь.��E�8�
��׏�yWiV��:[�.�����D���&_+�(�-o�j���t��t�,.���6��M�@�*� ���p�����7|l`�^�^К����3���S�.>KZ�q�V�e}	�v7_rӰhIW�^v����I�]Sj��AޯP�Q|����,}�	�x�W��M7!���q��hɜ����ű���Z�iZ�J��o��o"��9���6���,>����p[��ި��I[w�9�ҫ乚��l9�Y� �v��ev>1�Fa�<ٛP_Jx~�������aW.��M�$�/5�sv]\����-�ލVC�1q���K�rWf\A�B��N��.�\������y�{̷��n�S��\Lk��1lf-�^aj^Z,`��'0V�o�.�.�^���=W�SU�P��^�t��L[S�\��u;�9������'��"�Av��g��y>�=jؾ㐖%�aj��=�	�,�6��S������U�hU↭nҭ4,=��;�{m*t���!e~���x{�ܧ�?b0��1��>Z��E�Gn���޸0-����L+yqF���6�;'{J���71���e`��O��v��T7xr��� d��|�I��H����x�&�+�lv(����S<�Խ|���ԃL��Rӽu�qw9��77�a���gW���VS��46�g2�a�ۉ4r���s��I�J��窞�=U�ꂮ~�u��[^�Su��]3.��)^mC��sm��/���g&�\����<�Opp�]l�d����F��+dS�{�}븇�����ڈM=�*�F�[�Cb�����vW����&��n��;��Ҕ�5�#=����� n�����֔���}4���'��B��i��+���ې�fն2S<�i\��r"�c2�����iz���
�BJCg�]	��7d>���z�>��J�M�e3]g3�0eD�lfp˝�a@��c4�̽�aՙ�^�t�[�:­�݀GSy��E���IQ�F�������\�,AA\�>IH�L�C�9�i��-�5k_<�R�o�Nd�|d,:\�vH�[���b8�CǪt�.�vu%!;�M)���U}�stE������+�sPT�]!w�p9��Jח����5r�/oз4�I�qmb�q���:�n����_�D�CX��)غ��Sgu^P�״܉�Z�U�[�9�r�5	&�.5�Y���nj8����7s�pN�׸$=ql.��LۉO&��b;^;���i�-��ќ����vr�Ω��g��S<��Y�ʷ�Ǜ�&��o9�Z��[�u3�ˡ�S�~'/ ��;�ڱ�}�{*�j�����E�#�����<�'���h�Y<��4�8ӏ۹ܿ�ߪ�T?i�9WŘ��듪Q~�с�u�)���Q����kL�ZƱ�Ns���o���:���w���=w�.�N�]�it<��Q��E�i�C�ݶ�{���v�;�7�x�$^{hb�}KQ���q.7hd���b�sr�=_K�Vu&�zx��*�h+X���Aҭ���>��-���7v���-L�zjd^���k�r�4�i;�G(�H��R�P��ngw��JW.h�S2�K�uù�GG�[���+�:X�y�P�-�.���Ώ1��z�Wr˭TL֛{��Z���8^N��q����D%P��7�^�I�Q=�l��w���"�އ��g��t�P�G_mBb�7��Vm���~\�KbK�+�1�����5��K|��Q����z.�I���>��d�`ʃ�!����˘��N��cn�
���&yF&ZŽ�*��wAb{��vP�]�9��y��+:���Nm���w/\��3z�>O�U�2�%�5
dv�>��۞y�'�ZxB��=�p�-upU��W�^�M+������	��.�����'j�0Rus�z�׀w�5���R�&����).s�6�;�eƻ�,�n�{5:��{a���y�+�p�ޡ�%nMKy5�b7^+��Lmƺ�яIU���y.�~�)`�u�5{���ԇ��=�l�j�$9{���ػ����`��_K�q������{�v-�K#Ug����_\���Dz\S}諾`��3�%��Lz��]�*�å���s�f�Gv�l�]Zh5�vj��Ɔ�в�6*�@����R���
�]��K��U�]����̭�����'r�.C�ʈIu����rAvX�2�sLU�t��T��	��C2�HFb�jC�u��dZH�D�;,f�,=YZ�)z��66�d���Rv��;˼���[�2������.L�J�,�d&7Ux��s��)m�q��kB2���"�Ӯm��"�zF�("��Z��Z�WL��"�y�t,�(��:o�*�f,�5\�GP�u�IX+/�M�,e]L۽��6]s�S��u�ʶ��S_�I��IZ4�է6���ne�����G��������H6���t���JSN�>�u��u�*��4`��O���uz��1����uY�
����)0���-lݵV�fd��U�h-JvD��s0���n�e���\����.H�t[��]f0�x�@P��
��MDV��-�R����p�N����������Z̟oR߮>�c����Z)\����S8��hK�,�|Q��5��t��j�������t�Y��u��0k�����,��e��.�z�.Mګ�ɎjL8cQ�o@�k�ƴ�oTx�/<݆18l�&�}��_N�j�ôV�uga�.�r�L5����ڭ��[9��ܒV�cP�f!���:�<J}�f��ͥv�KK��c�2R�#��P些��`;�B�S�d _�]�wV3�Sη(���ĺ�w`���R����qj�qia��T8�Εj˺k";����	V���Ӯ�,<Y�����~Θ"����6��r��huyF&���.�K�ΠM�K�c7Q�xS㤹G��������h�dq)���u��x��dV�o�6�{�R���"��꺆,<�̑)SLL�	k^
���^U��p�,��]Ժ�]�0#���5 J�G $ʺ��
�h4�Yf��t�3��o	C8�6\ �[�9c|���ιP��W�E-�bD'��� x�2GU���V�PL�.�v�A���fF!TX4xl��<���{-���[��H���[�=�]luK�H��es�'2�Z�B��C�7�Yݩe���n}�,DgQ�]{�յ3�Y���2��Ԣ���u�L�x��'M��3,�۲NbEg���8ͧ8����]a=��D���ǀ�..׵ve�R��*zl}W���GUy]H�%�R	V�ʗ�ͩ$U��GQ����q�Ǯ�����*�>z��0�3�Ʌ������n�\nB̨&]�9;�b
=��2K'G��z����8ش��c�XJٶ��T�!�v�}��,�TE����\\�e�|�Ҟ�ިzAq���ŝ�����\�S�{�+-N�.�Z=�[��u��73������@�Ϯ8t�������/���ru5E-%4J�.�
S���AE#�u@Д�N�J
	�����iZt���M�h!O%�M4�P%:A�M��r)
)Z"���a(��t�h��N��(�J
���B��
6��Ck!�J�4�H�@4�˪���CI�5H�\�+AAT���HP�!IJ�ERR5�A�4����J퇒�&�hZ)�Z(��Z@���CV�@i(����SAHihh��h"M:M	m��#�>�+���`�x4eM�}˦]����EN���6�LD�����EE��o�&���!�+�f69�Ɋ��K�j��g�*���~]Kݧ�ӝ��){q��<e���3�ue^����Q6�`EJ2�T;9���{�}bݨ?M�뎙X9=jK��׸���B��̃�9��:u{�����L{Y���Qt��ũz���w��'j�t���4�C�:���BE����u=���@�P1D����ϝ���a�]�yp��KT�BO��,ܷ7e�W�WL@:�}���B�j��b�$�e�� �^��Hz��ު�њS�YҶ]�u�_�mV	 ��.<7W$�3k�䨶x<.Ƹ7���ɧ�U�cp��plWøO����K����+\o����v�-���Z�qy�o�Rt������)���Y�fo?y��z�=)��ܳ���p]�>��=�OʇT��nC.Ϊw3g�(�+z��o�e��%����5�l���P�J��o���}4_d^]��VE�Z8]�
�v�6�(ޒq	
٬i�},A����72�f�1��w�%�y&s��J�[RVi]�s�z��ё��v��-.Pݝ��v7�������u&d�����d��V;Hfm(�h�q��t��PD`�f/}�)֧A��u>*C�}��ʕ����Ҫ!.f�|#i˞���.�{T���;C�]*��q?'�9�k�7���g�3w�{-�$�ql!(_��V{�V�����Mƻ#\L\s�=�F�]���N&��ME[JA���o�bܚ�ʦ�8rہ����Q��O�*�9��K�w���������/mX~�O����VU���{p�Ú�H��7;M^��\�ռ�u�Úrf8�F�R��8�o�bV��9���t��p��q�Y�yr��Ζ�f�:"�{H0���ޮt�1��K�f�g�f*;��S�V�o��L��?C¯����-���$�9�Γ��g��r!��V3G���ڧV��RT�3�蝹t��+lL�.�ӫnSݶ�Sէ��v�s�:�}�*(�����E;\J����v��;�b/�nnO��^����T}���aQ�:��I��{�s���ݪĜ��*�Њ�4��M+=�B�.��Lq�*�c�����M�fP`��UeH)U:�e�h���y��?1��+���5�JL=.��3�7�rb��k�j[F���7n�U�
���uj��]�AS�^�7ه+�GZ�_V:]�<����z}2�_����5�������ڈM=����ª ��f�{��U;�,�f�u^Ԟ�qIaE;��n8y�o�Rt��j�ؼ�ם��w(g!�)��}m��iW�%f�s��wB�؜^V��[7��7Ml-���W�fm9���vP� %S酻���R��\�f�I�}]t�]�f��˥�>pTBLeC�sEHU!u@�#�IZ�`>9�)M<�dvEmF��N�[�6_p0���&!�e�b�u�Nt5��7��;C���~��e�����q{��}˨�I�Ì}�YK�����u���#����(�a�M�{�sݓX�c����Zp�6�ZܳZ��}�1s<.u��^��=�f�X^<�}�eZ���[k\9��H���R.#lC��f��K����պ��V��>=.*��vV���ͺ���C�o=��Btq,�:�x��+��+tE��5�(���aa�9�Z%�y��2��%eu�!����
�*�f�M�X�9n��O�՜M#�ke���=�i�������h�v�����A1�e��{�
w�@n|]�a�����.GQ �_F��}���J3[ɪ��D=�z��{�����.��Fb��ʞ��Q=*
B����Εy��������{+��x�f�ZW�^�0�'B�G�R��w�Yl�R���C�.��
Z}���m��ƶz��pU�w�@D��qҊ�-'=*�a��ъ+��.�ֽ��39�M]�:r�}��w+�r� �k��I}Q��B�J�kw��|�O,T���XI���s�ksx�����Tw�b�.D%�I|��������g���O�\��W�<����R�:o�nP��?�;��iW�'��k&ӛNgS�"Lv�g;�t�n8խ�k�׌ۙ\���}�F�_o=�6��41e�%�oz��ָ��v��q�9�q>���x|�8�~�?]d̶؆P�%��W}WgW(���7&�-�]}�$��/��q�M�W�]3Je��@�>$�W5(5�,Jۇ29MF��l�=@�H�c�%�4<����1<<؂�^4b4J���+���z��2�\F�7��F�%QlǱǍY!α;5ExJ�i짛#�7��F3�h���N��˦Q�%..^8���h�
Ѿo7�m��/�DD�1�:��~�F�鸕�5��wP�9m�k�\k��ȍ��oVOeKt8䕓��v+�x�Vݬ.�d*�y5�b��x�)=����&���f#���9��Pت�m��.��>�n�$9{����5o���{m�/�I̎H�ګJ�j�s��ϵ��k�f*�y����"��0�M�K�L��Q����=��u8��8�↩�r*��l��>��^vH���Y�3�OP����:e`�������yo*͸��0���c��z�%KV8��nr���W���ظTt�qp������;�E*�4CK�A�ȕ�<�,W �(�D�}Ctb��Kv�U�K6�w�T�P�wJW{�꯱-����
�u�!J���t3�i|���v�A���Y[�#�.����Vu-�q\��>U'���\�TrZ�s%�����t�Z:��8���4T�y�s�}��0�u�I�IR�+9��9¶�5�4DeJ�N���*��So�ezkb�|nsڶ���ʕ��9�~�*YQ��W�v�f��<6J���Rj��ȝ��C�N�ʙPԩ��Z�>]0���-����uq��~�T5���i�T��T.#�hw�yǵ��Y���/./�o�)��<(�{�=k�5�m[��7��}ʅp�՝a8�n�E�t��p3bC[�am�ӪWu����񜯝R���U]q��4j�ٝ(�ԍ�p��0#HJ&Ʈ��+~I�a��-#Մ��Sz����6w]��
��t�u}4��jV�XN~�Ғ�R���'Ta뷒�dԔݬپ
�"_����>"sћ��{�?�c@]g��w0p���.2:����uI�Л�vF����v�S�avZ����p�F	��}����t�Y�4���U4�Úmſp+��c�\�\�f*�۽{������s�
��ו�K7��p澷H��r��P>��ӵ0qt��Z�)�\�>�v�f��}��f'78��V�'���<��4�T/Z��׉�A���,���/i�l`r!:�wg��)��o+�o��7CT���[SUF^���z���Ph���&�G6Mx{DЉ��+�խ�ﴢ�ܓ��m��&0k�n��in5��7�3J=����\nw�IY�h<uf5_ �����w�x���x]�X�&�+��:�Gc簦y�W(nĶ�6J�Ek�Y����Hj�9��Vc�r*��Ռ�G��k����{A!T�`�U�p�<��SݸoU=Zx�/��}�`���V�J��W^�L��s
��ہ�&��4�D�{egWɭ�q\I|�S�-l1�7r2�&�8�7��;\��R����ކ�������m��vs�s~��d�3�W�́"���ȓ��+;
Sˎp֕��ߏ��<������o��D���te���rv�(�*������J�l�S��-����}9��=�1��2���}�F�Q�S酻ٺ�i�%{E>N&���#�<��l^�6���G�Nb���'���G���v��w.�u��$_.i2�;P�1�d#�\D��ף�ߖ���^��� +R�;�����ӛ�2�t��۔�Yv��l̎����0�5fH^b�})���X:�R`s��ʌ�0Rw������g+-��h� �i���k�WP[5j��U����z�tѢ�}f)N!�z�1,D]�9уYBC8��c��ܱ��	�so'����t��$ö\k������+��;��U[�='���̸��j1d��w�N��k�g2i�	,A0.�-�6�!+�y�5h��%��̾YH���n�ڠ]���9WO��)Gϧy&Vz�M�j����z\S|TY�DB�d1\�i�uӎ��1�=�e�l���r!�M�ȳ��<��<�zEoo��V�hOt8��W�<����یZ�����`Ua��kOp��Zx� %����c�Q���-=P��o�����rQ!xX�B��k��Z���R��B��d���&/�7.�����Y�'����_*�!��gw�yʁ��}R��-��[��p�cOuV��7&��k^�,�+��7��t��!�)W�{y� ��}���Cha��@�h�yg�l#Z�8ڦ��#Z��cxUk�ҺPj������un��<�Rc�bR��j�b���M��S�:���!�����u�71����kU���e�١tj�CIڸ^ӑ���R����;j佹T}yawr��k��M��)}�~;w	��;�X��W��/=g�v)��4�{��Ʒ^7��|꒸�p:�_r�BP�Dw->��r ״�Mq���o�����nZW��O�S�r��Lҙ*���`:�	�-=ln��=��-o~�ޚ���L_iT�J���loɽ���d�}w{��6��Z�ɖ�ޯ�5j��V��F'��l%�i���̸ք�)꽕;0��*�蜞�.�^��i\���:��X��<����2�P�W[d�M7[�Ϊ��ލW�S����<�{k��dTzx��);����	G*�8�bi�������z��[P6�����l%Y�5o�\���{nߢ��W������t�ֽ�{�Ƶ�9g����YW�fT؞k0M�4�C��Fv\N����+M�\J�������yo*��so,7F�ox8g��g8uoV׊������J��[����EX���$�WyKQt;�yd��vT�ظ�F�H�etH��ˊ��q1/Q���t��D��܍��B�1��v���E�z���FMu��X�ˀᎹŵ��	ѓgp}=Tn�l+X�{Ý.��Z���?Wg��x�hL?sb^�O�'��������W�l9��ɹ��1�TQ;˛�On:Ҹ��[E5r�w��I�S�n��g���|#9P;/��Qʢ�U�G=o7.6j[,�)�r�J�j�nv�|Zx�[�*������Q'��r���\�Y
�H��A\�Mv��ᬸ�i4�ʶ��U�Rw�Y]�AX�aUo�U�M-��N�k&����Z�q�V�br�@�-F��u�:e��J��g`��`j}6�=:�wXX�r���Є
L��n�L3�s.ԅ]�_m�BƬ-��)&���[Cw�2����=�!���]{��f!!9��'��x;��w[�Ldj:;�XWQ�=&�|�0��m�ad7,dL���ԕ�K�T(�0��[��~��ԫ�i�q�z��͉�M�ܷSd�Vl��	 R3#��
������e�8��mL�t�&l�R�뀼l9ΊC�n�mw��ע����JNПm+yM�3۵�F��e"ą0�5W=�R�:�%��)zC�4�w�e9�ۼԚ�e:����n<�W[Wץ�Me�t�	�*�Nur]@Æ���X`�:��Zfr�{6��ı;m�
)�2��P�(�&	O��;�3kt\t]���t����}�ЌI��.�3un�f�u2���M�Nk*_:��}�Ln2JC4KO`�֘s�ڲ�� ����)[mV��wC-��d(H�e��&�� c
�`\���O��Ϲ�6����vt� p_=�2���l%�.]���$��	s/����ɴBL���q%�'N��W��T�m�@�M�r��V��R-Ce���R-	ncO�Ȼ~�S�*��q!^�Y�V��o)�q��"�,4jytU�^C){�կ%�~��:����"�{��Q���B�=-+w�j̙F��J�.V���Te�#�G�^lZ��z=��Ƭ�t�t����.�=�n�J��J����eP��{M�Cxg+���!<}4�Toաv�v��C5���B�tt�|�OwS�,%<�ǅ��C����l⻰����Rm��CU�m�9J#s�,5Њ˫|�Ӂ�W$��vv�#�l�hCb>���}ȭg7/�U�]�Nc��"��L}&Ь9�5�/t�v���7ը�Aw�7�T�Y��B��r���EC�5�,�`�i淎�<�2˻r��)�=��h�mZu5q�X�F^j�V�r�N�:�P/�w1�
��]��3�e'oi��s�2�[����H���.�յ���:�l�u��H������!9݃��o��]���MA�gb]�ʺ�)*
�;��WJ��q��a�W9�WTs/o�[��g�f�:k֮��˘�7�[鍭x�b��c�áf3�L�9��*l�c,�ͺJiK��C{c�{E-�6�V��Y�R�`���(+���Z�A����s���N57X��n��j��9�wQ�����b��*�5�;�əݶ�̢r���V{��˗|L�D�w�v�����=�r�4Eꤻe%WX*S�9]�;�A֩�%PȨ��M��d�:��:WAΫ��]t�����YZU4��7w�kU��gEd���ͽ$�9E�D0Mqڗ� ����Zv����_l����S�{N5/q"��8��#ʧ8�	�J��.��l��Vg��<*(I�����T��:��L�=wf�.`���*�H%��G��-r��>�$7q�:iǘ���:����m �C"����k(�:��ܫ�W�����ӵ#! J��9uد㥔V���z�f"UZ\�ڝ;�+Rk+@wՙ���͜��GT��z�ht!�^q�OX�2�o\<�"��h�/nNH7��TJ��u�J_}�蹱��nv)��՗U�6Ɔ�R�"�]S��BQ@��h4i��
K`�])��it��К��ևJk@�KN�q4���+E%��E:e5�F ��9	��К9r9]	����R�P��9���4�:
6�Ph�C�HS�9Q%�յ:��P�2�A\��44�����E;`5��ZZV`(�:Z��T�֜��MAl�N��b����SA���*�� [6ʔ���"JV���4!�M:��5�"�k�Ɗ)tP��5@�mR�N��M%7|����6�;��F�И��`˚�w��\GP�8udu)�Y��MM�DTx����K][�ˢt�v�X�E�Ԫ��Z���u��q��"c\TLs�=b�F��L)�	��xRQ���Q&q�y5c��}�g�c�5�Ѽ|.�g���駊z��kwUSѧ}���^^}/�F���Y�/V�r�-�;7;4����T���t�t���_u@�J����K���*,���w{}���p����g�ݮ��Ov������b���`<U���O1أ;7xZCx|ġk66=�3�u�s�U]�!�six�g���@��s�C�0!�>=Tnd�v�)����6'��\���<��=�o=ZzhwiW?@:�Q�/m��X�w�j"mˍ�»`b�������c���Ml���P!L�K1v���k�$!f�׏�@󨓊�{�Ҕ�kwp�5��=���*�=�q��q�4Ok|k�aVm����0*�JU'��%��a��㇕[Zb��ב�\���lG����^��k!�\v�� ����6�(xD�-�s�.� p�YbV��-�w�Uu������o�[5�O�f���p��٩�0��\�}�|\�k*��QS�b��;.R�wfթO���<Y�Zܧ����w)8��y��7O�#�D���"fk���wg�-i�{A}�SJ+��\���Oh��:�q?��<��tTkjJcg�X���u'J�+o%D�i�9�z��v�kY�{���������!܄��w�[��X��W�\�^�1B*��ޛ�*�歗��@x¸�[�B,���.5�}P%Lut8͋�j��5/�k���]F�L;�\k��Ȗ�EA����}+�K�:৯�3��l����2?/_%F�ӆi�ȴ�9�o/%��t�<�\�[�ƫ^�W#�OLΑ�Y����6%��6�x7���)okF:���`��U��_U����ǥ�'���$�/kR���&�cJO|�<��Z�9g��{r�=�g.�fTt��U78,`�Ζ&޿�>�'.6|z�9 �S��ƽ�mr����WÊ\�U����O����[�mJ�����d{��N)���_����$Y�"&YU�oq�����Ik�ؽ�S���Ō��m��U�ʭ��+q�14w^G!T;��l��>�̏y��t^k��M_o[̓&m֞b�Y�G,H"�+���<T�f�5���N�mNy(�b�]/�"��5��Ψƶxկ*޿'��T�$~������v5˝R�9���1D�_.ns�i���{�FS̸����o�u<Ym���;J��D��*9-)p���7�n'a�c�o�����I?��v���+��U|��|�$�Q_+����M��u{О�M�(.Y͵����ڋ|��n6�_jPv��k�g��|��pJּ����47鞊v5�5�m|�s)k8������:���Nn��I(ه�ٸ{�r�b��|�h���K�j�S���.n��/Z���_.��턲\����b�J��W����b�{q��up���[��y�g���H�P�[7ɩ��z�L�s����pdf�&���hMc���Ďֺ�]����s��M�g�w�1n�%,����'�ىwu���ST�f̾C%=��|AѶ��컚�x�4�f��F��.�(�^�}�� |��ј��`�	%;�a�q�.Ȓ'4��n�k/,>�����[��+3{3P�P�""+��˓�x�c�ң{����tOOm)�*���7��)��nU�}P6���V9=4m�&9�w�`��׹�Ȼ��\�g�~�e[P6����5Q�O��TĲl�t7=���	}W�����p_���̯����q���,��9��ʽp3%��n>�^��e���Ϗ���-��V�z��\J����o��k�D��/725��kx�lo;o���*��T{ת�u�v���|�Խ|M��5�Nj���5ݞ����ܲJ�qh�V���7:�5z�U��.��V��o��Uv�Sս�_n�Z��=q\O�t��������}Qn��nX�KʽIevJ����I�i�Ĵ��Ψ����+��; >WTr؆4]�v7GZ�V��O�+���kyzᬸ�SO8�n��U�G�9Qú�S���R瑘p3�����J)�<}���žP�7GWl{��*��F��!�a��ߗ�1������y>�ݻ7f�=�z�B�⊎k�L�4�[G�c��Ҍ��36��r>�k�TA�ʎ��%^��|�G:^�A[����cN��������\t���Ƨsy+d�\�b+o�eɛ�8��T�-O�;)9�8�C?wӲ��~�ϭ�L�n��:J���y��MC�"�:�W)��6�WMoHu���%5t&��2OI�����ӑu�{'-o$��s*e��u��~N�B:�'?�i�ܝJ�ˀ�^a�K m�[0O%G�eJ�S��V�/��l���nX
Y�!u�7ʯ�Z���QHJ���x�����U����]F�L��k���&5�D�=p)�Q:'J݉fQ<�䏃͎��ª1���j���,p�p6����,ꛭ���� N-h[�a@�{jg��<��>Y�Os<�����`K��Od��v�˽w�i�|x�d�.�JK����������zOK3����������Nx��NB�5����-k˖[��T����Ƙ��RO���^=����V;�ۅ�0*�w�\��U�.��dyo�a����e��)H�Bcf��7�ʶ�/��cs��QLo'f���G��7,���b��^ѢǞ�B���H�;��^uyN�����S��\�}�N=z��R�)���Nm�V��pH���Q��5� �.d�[}N���Γc)yܱ>ҹl,��q;˜_�ym�{���OM킮�Y��f���'X��$r��K������i��/��|�d�6�U)[����E���3 k����*R��5�����އ�	���/��q����j��er����\��>D$GkQIa�R�[A��EL٫o; n8��+�Wm'��֋qΛ��T/�L�(�ү����i�1�D��/Jy��^�kq�^\�vI���� ���p��o
[rV[�3�Yw��|���]�g>��:����i1x���*c*S�*B��B��F��;!�wa���O%n\�ܰ�b�JK�L��<aC��n�����e�}쥴�ymg���g����iT{aU;�s����i$�a�>��.�N��G/���x>�\t穉6پh��,��>���#��Qi�#r�[��6M�gLiIh}[SvϜ���f���O<w��Y�4"ک�a�6H�~$R+9NN�r�a�)�K�-�To��+k��K��}��IM�vC1;�S��;�@�=�c�=t"	�܌d�8��s��;�ajG�>�x���f�(�&��7����zB:tM���xe/��:mc�Kٌ��<�j4���-5x�Ŋ�y����Kj�cp��:�͆����[��[��ʉX3�`�S������l��p��_L��I�;�,�����[8��~>��4�.=�����K_�z��=�뵞�θ��֫�Qp��l�n-x��u`�{%��*�Z�W�[��N����*zTc���t�qjZ}���n��]�9qM��7w��g�XL*���Q.z������b���ˮZQ�cM�o�rVK[{��v�]넖�O�W@�q%�Q�b�V5��Ea׹sX|���޷ru�!T��=:���hq�m��U8G~�KFF��y�RԲ�ॆ����w[����n�\�p�|�˶� j�wӳ�����:���)Qzq����C-��ۮXj���vF�ͨx�T:�����}8H���j��R9ˬ���j�t���S&�0ˢK{�'���U&����'zCsv��/o�
E�g��X��<�矏�֩���e��$x� mm�97��;k�Sr�E�����~�˻X��z���ws�Ȼ� �.X�Q&���8��#d��RF+�3bB[�aoc��ZL^�Op?�3��V�lU-]D��Į��_f�~	lԭyp_i[	4������^�E�s�,ޯW�B�Ô	ң�]P#V��[���iJ!.r��S,_m
Ź�ڤ��t�c���VCr�AT� �~AnNJy8�uQ���w�j�r��1M�nO8}�j�`�6�]�S����;r�>�n���D�X�dhx�L�!�睾��[�>�y�5��[k}jځ���|,�F�"��j���0r�l,'e�<����X�d��ޗ��kX垼r��N�JQ@��墹���jz�MT_b��qN�_��i=-���v�_r&�c�@tܷ��8�18X�S^(#��C�*�v��;�R�Kߦzz���M	H��@��6{���?)��d�����,9��Y���.&4��l�[�~�_"U�[��IP��F��Ō�TUd��F�wp���^�Rǧ��"=ī�r�L��=ɭ�z�^o:��ri�Y�w\�131v,�DN{*"���*�[ۅRR�KM�N ���j We�YS�i���0��(=
�\8���ϝ���v���{����9U���㚤�X�2��G�F5]��5ŨI�&�_���fg:�ڢ�;N�61
�����
;q��#����J5[�pը�SO;⭻�nSΤM���yY��˖#Oq�Y�!�#y��ZɨR�sƟS�'���wn�,��x9 ^{�|�OڢY=m	�>���uo���xg������s��D�����:�r��WU)��:_5"4��bƯ�o��J\Էҳ�	�l�勶��8��pUT������u\��B���Z��kz��Xp�Z۫��kn��.x�u˙���0�,���b��k�]_�zr*�5
�뵻�]>�3.y��<���9uI0k��k��ȝqQ<��pZW;����26S쾝�J��7�3�B�t;����X��Cn�58y��/.����+v5d��,[&偊N�"��]�y7LWM��\�S�8��	ԣ��YY˭F����
����H�wZ���EN�0�RSNu��+h;ȹ�˻Sn�[�rc.>�8;1�\�(�!t�C<� {J���D	�t����{+���U��dt�c�3۲է:�����M��N�F�t���=	!��xsy0�g���ߵ\��>����w�(�Z45��md��Ѽ�R��s�r�?��{ɇ6\��3~��,���^�{�x@�a(78��B�丝�뼵���֟��)T�V>6M���ok+�VN���������^��
ym�{��*����V;�e���&�.r�S˦U':����%��Q7�7)��%�g��HoW�9顭��߷�7�6�k�(��a��U1qS)���[�<����ȏp�3��#�ߴ��c�x�����m�zC����ږXD�l�n(�f�P^9m��ۧ~����ف�/�=��E(���jW����#m����:vK�����O0���أ(�$�\r3�7�=���������S�������a�F�������ul׽2�|��]L���ofY�si�ܒM��K�p��ޖ���u����l�V�PM���|����Z�eNr�q6*N����X�O;�@/�v�N/b��u�����'��VĞ�@�JU��%u)��\G7Yt.��5��;ed�韂업�;@C~�3���Z,��,����eit��}��ќ�6�/�te�ݵ��b
D6��-}�7��-:cm	��b��pVR�����xs
�;�2� 4��F3���p���b��J�Xq.�v���ۙ*+|���;^᭍��&��y��뿣3A͵��j> �+����e�H}/���
�@�1ٙ�Q�\���oV�o�^�b�8��hvF�b�K0�IP�`B�K��L5�gWY��b��E�'.ܠ4�t�t=/�cR��S2G\�W��j�V<���5#5���]
��e	e�{]� �{3�)�uuX�;�8�Q
�����0���DЉ�ړ9ͬDW9]L�2�Fv�a����i���ӽVmg����#��v
xu�>ϸU���l��|��Y-Ӻ3��}���45�j�v�V���w�a�Fy�ۖ�O?b�ak}���,�a#gE�VL��:������iv�?�Gu�)ag�c�̙>��Okm١X�oov쬇Z���K cr��Xu���n��d@{G�8�g6���I_��;�l5��쇦�U�N����5	��9O4��ವj}�F����݈m�,'i�-�#�ǘl*�w����jAQ��We��EMD��6�v,�x�*Z��]%������l��%(.�k����an�ˠ��1f��9M�N<5L[��G�%��W'*Cc�2V���#�M��(/�Cn��#�=������릻���05>���S��s���h�fL��e�Q��ʘ4���h�`_C����:�v�@����M.L^0��o���[�rGxKq@�v�wq�I5��Bd._��vJky��)�2�:����#JLo9Z>|N�p�}��N�fV�TqQefvX�6�ܠ.q�1Q����j�hM�;Sg>&^Mj� Mf���]�A���J�he�Q�4x�8��Z��r��X��aޗ�ln�X�����d��5d&_P���(�v;]�I[.;|���B(0�)�U�n�<�����gf�Ό��W��*�F��kѯ%ut-�o����H�:�N�<czSӌ�>��Ӏl/�+�W� Ր�
9k�.�9&��_q����59){ji��n�t�`����G�bu��կ��Y9�GJ����P�T�9�Ul��_[uo��F[:�]i]>Y)�N�v��e�G�Nu�J�u4hi�i<�\�j�c���"XX���ȃ��:�u�ÃN�go��suGO��!�	�Q�)����N歪�}�,���n�k���9K�L���V���o��w׋2�J�)+F�zqF'sy���+�>"����A�4�5�i]cd�ƚ4R�E!����ӣB�i�CAI
+ZJ���i4h�6)*$T�m�q�.�I����4&�i4V��B�֫KC�����4GN�4RĴiQA�)�	�	H֐�6��(#`�Қ�t�ví%��(j��h(�4�h�]M��i4��g��bM��N��gZlm�*����FjK�uEkE��l�5��j)M!ADIE	Z4kCA�Q4ҚIIZ�_�uS����>"�Y6�s��f@��ۛyjI�Ƕ�4��D�ہ:(�u��M�8��x[���8c;
|�z�ŵ�@9����{����<<�z�1��޿3�Oi7޸;u�̖uT�Ӧ��:��H<p��7����g�g��4.�<��@>
�\�m��c#��g�>>��.=1p7޿\L]���3U�طbu��T�C�#����/�Ѹ�-l���\��-5w"�m׉�G���v����0�w�ji��g��@{&�C����B��Mle��[)�y��w��17W%z�{`ܖ�W�㔖��UK�9���^346��m����2����6�s}^�q�/I�ib�F�hּ���{�i;���/w��>�H���LOg�t;�NL�����t>���4��צ[/��{1��w�d��x����ϕM{Lc~�^;�	�߫p�?~��8�H;:O�<�7��r��yK3���Q�S�N����p�B�O c�_x��|d꟏1F����t�4����I�?a�k�¹Q8�f3+�>���d֛�� y_�L	Z�-W��|��+}u���L<�W�τ�(����A��_���>�D �3�>�FY�C�g�]Y�]��O��ծ?�Bha�`�_�xmHF��QB+@�ݥժ��m�R��[nw\���n�f�;KK��V��u�.�;}njT�7%�z�S+�{��#���<����8�!�t�R7W-.�I�����q�Z��Y��%�˄م\yJ�,��stDfm�:E}����;'�h[�련�J$>(ʨwg��2�e�6�������{s����W�֟w�x�r7��r=n�8���Ӳ]��J���b�C�[�ˑ�G�� ��n�Z�>h��s\f�z��ȟ��x�����(�t�n�Z��e����.����ۘ�u9���Ӵ4d'޶��zF����߮�y;Gƪ���^q�=�ӕ�޸��2L�@��J��X微�W��������\MǷ��e���:�ޡh-�3��:��\�P��E��@p_���E�ۂa�]r�o���O������Y��\=5�Gu�A��}8�_�%�Ϫu%� �_W��Q|v�j�F�jy�J�3���=��)֮��ĥ�ؖ ���
�޻�7���L�?��������#��)�K�x�'��y��7��}��4�T��_��{ޠ;���*8B���9�s�t�����K�&�yW��j<d��?Rl�MB�ˏ%�0�}�Q�����FlyQ�6n;�	��?^�P����N7/B�����9���R�D޲���s����Z��1�H.'�5������Z�'z���[�����MhWrfֳ8,�_u Mu�,��O�w*�GVIe�Ε��콬3���5������F�d�E��7�n��y�cTҙ��1~���F�*}�D�����������ݑ��;Ӟ2����\W�ߗ��j�K���U��G�G��wl�%BwL;��q�t��`
�u0�]`/����6�iSU�HT��N��9X;Q�I����yuh�ٷ#qΓ�pf>UⲫM��_�WL ��#��������	��+[�<���)��xj^�'��zvE~TX'��-��e^O�(���yft�ݮW8�����L����my��D���g����O�F�y�1q�]%�RIU2¡3��=�.*�z���D��|k&=�zG�����@��>>���_����dZ���ƙ�H+N�u�BO����T��'u��#�'e����'9����������7}#�_�C�Y��ɵ#�g��o��s¯Ӈ��$�3�H-(�l�(/sǚ(9~��>G��þ��4"�Ƭ2X�οpUz����A���GzmO�}������Y�|k��n5�NW{�![~�ً�OXų��Eyz�q7}R6���v�{�'����k�$q���P+�������6��#(�ͭ��4���!L_U�ƺP��X�$�կ���N�U�!:�܁��{d2���s��|{vv�$�x�q�Pgʞ�>{rյ��7s>�V�' f	L6���Z�B��s�����216I��Y��T��,�q̽�i��ZF����#q��X�	p����S�~�~��������uh7޽�U~5r�b�U%��@��HW����͚3"� y����j#�m�����O���x�`u�T{�~$\��I�S$5�P��`�8f���=щ���}9<��+M\l�=ޒ&���o�d�~�@�g��lw�QghӺ�͝��B�ݻѓ�)�h����W�
��2�Uo��Ɵ�z��BU����({����������n��R�R�>��<>��T
��̕cݰ'tßN�آ����4U�屟r��x��N�ߏD�YK�:�O+��k��zq9��盒3";�	���n}�E��/�򌕃C�2��﫥-uNfw��uU{I�^��w��%o��w���ub	��?�5�������#�w���o����|��+��Wx�~ۄ���s���9�,dm0�m#�7�ǽ�\ט~��QB����7�����Tr�����W��7}��a��}r���_�k�������5�z���g���h�E9��4<�]@��_�c�?�^�=��:^�6�&�''/�FNA2/^)3� B2�����Xc�LW�!�YW��M��~r�;���hx�Q�[�#υص�Az�;���� ��ą\��; ���.��`V�\��m�.��Q�yYO�Ef����d�_#t�����V�����w\ӽ�kٺ�,q'������M)�����a��z�{��8�z�]Y7�5P�ڼ:�B�F��\s��R;&Y�D�Pf:��w�l�T�ƛʉ{�йuV�ʑ�2�O��'������jO�=���s�H�~������ '$h������k�gEF
�]�^��x��2k�_eE{�^��As�+��H�������f�=�|n�$���>d�=�+o<�W%.�:+���-�����0�;��G��=޸;q�̖{��Y�n��㓳W"����˂�yM�=����!�Cj��O��>��/�2�۫d�/��d՚��w��Q������z�TK�����^����b�5w!�>'�8��5nY?,��m�>=X������p)<�Q�d�#���պd?����鯗{oê�6g�ї<|�zV/\�G������d346���
���2� ��g��n��/O��"��7nf��^�+�ozO{�گ.rwh��P�y�'�ꑾrrf�z�(�>`l�{��ry�ѩ^�����,B���;�q�,�E T�|�ގ}6�n
h���ߍz[�L��@�)�S��ϖ.����i�i3�T�����
I�O�r� *A`j��s�`;ß;��[���$(���+�oVMs^n[�MP���N��7_��uC�T״�7���	Y������~��/�'/I���a0|%�I����|:tm�9GE�S�N��Y��cRyϫ|T{�^)w���d�g��3equޒ��Z}��٘�).�kMӐ<�i�?-v��/du^~��Þ�ɩ�ûo�Ǟ���mx\}���9g	J��<4g��^�F�� 52<c�=�Y�����\���4��ޯZ��з��AQD�zKE�EG^�W�P�	�g,���j��_��%W��d���J��>�#�۟o���޷^�/-��d��(Q<yL6�U-ar�zGY���C���w&?T��#�jk����#�O��#�W��p�#���`��,ۂ}l��-ݟP�;��MP����tĒ���-��7�hh�O�m�u}������v�>��D�x���u_r�6�z	�@� l��5����/_O�0�ӽlv��K������ÞجV~Z�1���./�`�K�Z������ p�+��o�/���U��C���}7���`:s.�]s���~i�Df�j��]�ǹlv����7�gqK�dYF 0Vы4��]�&�����ܬV�)jH!��}N;^� �E�N��3���F�}�NԮ���M�r%C,&���UЃº���������7��ڑGE��ٳhI/L��K+����ӡ7��.'�쉸uU�FIh�8���7_��6���.��_����<[��>����~��zP>� ���@�z��ܺ�L�>Sg��D����k���>��}]4��g���>�5�G����F)~&M�{ޠ;������Ճ��Q�P�����U�=X�J��+�<��[(Va�m/]���������k�ߚ�~� ,$�Wf�u����7J��gGx/sæF΅�T�:.��;l��ۼg*�df�P^���W�Y���b�Qz��?d���z?�����R ��a��a�Ee{�ӝn6�k=��*�z	���X�H���%�oUS�S��n�Y�Z�c�۪� ��]�Mv,��qE��� S�h�ǎG��=AV�o��s��:��~�Ab�����QYV��6�/atW:�O�p�WO~7_��u��6tb�^Z�d�х�􁜝/V��~+>�+����b��u)J�a^x���:�F�x_��%��}]!zo��^.;����>>����VEy�{���m��4���*}��N=�����t���wZ��D�]~�Vvo����csY�u�;��/D))����$��d��I��h:��N�)���I��H�z������ƥ3}EaTu��%��$��}��nm�R�\�)[�:g�:���!�էP�����o��zK�3u	�g�@���T������幠��}��ёޏS��=p��=�~������}Ϲ���Q���S�"�>�3�H)+��l�(/tCǚ([��н��z��}��_��h�����^�SM�����;j|X�3`�@+�W	�Ʊ{�&�<C�k}Bw^��K֖߰z��=�N�'�鑞�]�{�G�p��j	Cs�K��\e����a�-t���|}�jF��	��9������zǪ�Ʈ%�Z�$��z����ݍRm/q�҂}B��83��j#�m������'�#�9�}pzkć�$܆��ν��k�]��j�{+�V�mX�S�h\W�i�/o���Wta��2S��{ :�����S�"/�kO����n�x���Q^0��	�1_K[z2��M_�,j�l%���=3k�Fn�K��f{��� s�g�+JQs{�fJ���>��a�z�M�z}��S/j鋌�My׆�wv�Ź���8܆k���=��y�#2;�	ڈ����C���7����~Ӿ��y���R��Rnr)&rwu��s�gl@��Sl��]�3�s퓳������=Z����ߏ�r�|'y	9ǚ[κHSW�EZ�t��ͮѬ�k5_�-P��r����2�)��x��X@%�=��R��of�oRf���.ࣵ;v������ȝ�q�>��2U=%��������{�{+d�|�AӤ�#�#]�F8�}�C[��}o��}y�����U�u4�@�u�����	d*�5��S��ӷq퍗��t��i�.�v�N�{��2�]K���Hjtx�5�^��C�[�^������`�����eO���OOc�}g	~�,e<X���#qNC*�l��u tbc��X�O�]��`�;n�fo��9S�x��-_�=���b�}u�YD�Fc��T���Fd�'�� w�x3]��[:��gz��
����#Έ}q�[�K�A��f�Iu��|�і��T��D��܅>݉�Xͼ�W���J���"�����s�HΈ~���q�-�9q'���@�kznOmX�`����� ��|��qV��G ���a�F�������ul���@�ۂ{��*;U^�}��;�j�:��E�~��~�B�Ɩ�py�m����_����%��;��ߌ���1�;��:w٘7�͐�Z7��#{�@���п��x��#\�6����O��������ʊ?a��Ԇyg0M��ri;�7���$(��eXZ�e�)p4��0��>������7���F�%[ZU
���}#Sga��;sV,�3w���6�ԭ���'6�ʹq
�dol�s+��J������y�=�o�n�_u�ƽJ��S�f�����n$G���i�s�ͳ��j���\��UR*5�Q�ﺾ�ݺ���h�'���P���=�U��F�'���!���Ml-����;�G��h�������yV�O��������G�~���y��XfU�a�;8�wd,�y�w�}�=d�+���o��Y�°�4�5���ǳ�N�ސ=F�R��u#}�����P���Gx`�r�NO������z�1�R��7��5{}p��U5�1��)x�|'�����Ӟ3���mMڬ�7Xk�\+��;+�3��᳡�T�^�������vC
�<�����9�Mx�jw���{�T�;��w�f?G�6霈gI�=y|��d֛� y\m0�@��W��y�&%M�����U^����W9~WX;�}	�!{��H�Y�R�0�ў�w�z�����l��Y�䚆znu�^��Uo_��y�{�^�c��hxqyHs�련�J=Z5�P�#�֣w/��`Ô}���������L���{o�x�s��������yh<�;%ߔ��.W�ڳ����ֆ�m`ڼ�-d�ِD*m���)\�������\��)'����W������s�w6��7�E2ڠ��B<
������*v��/]�.��ǥ�#���\�7fZ�U�eOX����(��6K����8�ap5����lO-�e��s��FCc�Y��#��7"��m4�ǭ�L>�b���M�r\�jU�T,)��-�����l���B��=��rT�&uIԔ.f:���>�fK+h.䣆�7R�nbu�6�mp6k�6�!Q��C@���,�`�|��7W�6���v�$Xij6^J��7R������{ʔ�d�jb�����:���ѺY���/���U���y7���b/�B���˯9��Rո%�{ ���z��NÕ�g5�2����,��������oF�{uţ����m��F���*����E��)wBy��Kh�4�|IGt�:	;H����++�.I��-Sۓ� �&���� VPC��ȴ����s�L�Mj�K�pߕӇ��WZ	�� F��Ԝѯ:j��Mx�V�8�9�A��#t�D���b`�9u��(n�PP�4Vr�'�+�!:[⻖쨄�ܳZ���RD{��L�k����u�[�lԞ��MKl<��ll��b0M3�f�{Q�	ݕcxc�5;\��	��겤(qo�>��j�@uƸ�F�Ts^���i��*�wF�9o�uꦝ�n�a{6�H���b�ԕ�&����2��|N}��'eB��֨�h��(�R^�9n���܆�fb�#lsd���Н�k�U�q��zX�Ir�h�R���D7���w�>�;�����x^�}Y]ҥb�#b7;t���^3�%�kG6�ۙ��>��}vx��k�OU��eL����e��$�����n�Hq���(��b.�JX=;�B࣌��x����1M[�ƑoP�ǭ��8Cq��w}���j�
�xޭP=�q�}ϸuG�M�U��H2��}�Ő��ʹ)��������;j�2�7�V^r��U�m� ˻����ζ�jS>���h��]�ͼ����&ޘ�8k�śd�gqS�i�W1JhM
{ы?�����Q�����<����t�ʖ*S���%o>�I�|�{��l�`*d)mi I�b]���g�����*�(��)�1���T/��8�|�Μ/x�3�H�హvMʾ��yk��J�Mr6f�$ԝ7o�{���%�1�mγ��0��G��,�;�Ȟa��Xb�$�q	s�V� �lF��L�+L*��q+�C�Φ���(�^�[�w�V����|{��W)lĆ�U�r.x�PN����p�Wr�wY�oc��Y[N���vf�Y�;gw�;$��Q3�p�E*�{�u�,K�f���ؘ�Z�0ZBD2���3H��ػ�q[�6&�wo.��m`�O��������lF�"* �@h�*��M-	AIIi�+Im�F�5A�3U�������ZZ����K��"Z4�ҚX��:�&�&(���B�(���X���%CMQCU��4誠�)�V���*!���*
h��)(h��(�����C��&
�X����
ذkl�i���*f��H���LT�T��[`��tSDZ�j�����u�j�����*�FM ����"���b���bh����%�)f&��RX�����m�UDE����(��Qڎ�����y�Ħ�YY�eܭ���s�7�j[o���[hP�	枬�1�O����*���S4껛�Wk̻���Q׈M����L��=K�"��3>w�9�'����3����ߏ�����O"}E��IG�v3��g ����Nb�S��Z&�Ӵ4d'޶���؅~�h=�:�G���{�Z�p��8��mQ�3��	�\��=+�k>��������3ӽlq¸a�X��;di����"}�W��߮)əg~D@j���`�WQ���8L5Q��C���0aD��=·8���v���r��� ztx�~�h����7.��6��ѿ���`��Q���-ޝy�f'�}�{&_wu;��6}��j=m���J�Ƽ �`u�{�^e��f'�F��XݾU;}3۞��$��z�����5�n=���7�9~&O��|�:���G^��=W�2Dk�'�(w5|�ŷ��Ӄ�*}�D�g»헦�u��ϒ���}�Q�����롰e�3�.f�uo��V�.�FQ��A>�1�8=�DT�N���:N�������}ʽ��#�53՛F�"mN)J=���k3��u�qN�����pf<��{Y^�qNt�� ��u���>�<�$h�֤&u�o�f��H�:���o�nG�]�g6���0�u^'x�;R��p��InY�	�l"����M"��˜�"����D})rቶQ�<�7F�b��Qz��\":�ff9��T&��v��.��;�r�B� i\rJf�c�}ʚ��yM%;�{�G��f��Iݳ0��)�73�h��[6�XR22_A�U�^�� f�ﺝ&FC���)�~�Ab���u�U%ؙxA��1��
�	_�٫q]�9 揢��o���*�NW���P��W��vy�1{�t�2ԒV�N�d�Mv�����{�L�;��s�Ny�׋�ި��|}G������dAu��}�.���}�:���:;��Z}���<�E���HL�'=����������77�<x�,�/���S]�*�)Oye�Cѳh�zmK6�$��<�)+��l�T���ǚ(\:~�'Tv�����
=�9>H�/P���:@���ǰv���2 'Pf:��
=+�V@�|Qݛ��a�V�\M[C����%λC��y~�J���m��ث����� y�8�n�^ğ���WEn2qB!�=^��f�q���~��zgx��~>��n!�נ_��Ʈ%�Ū�Ի~�n}}�2/F��X�ԅ]O����5��;��~�p�>D����>_Z�5�D�S`��!k���e�ͭ�謽�y[�ذ��s��R� ���Ϧ]��kL6����@��J:,��}�7]�F,�ٳ{`Ճ��&Qs�ou�����-����#Q�D��Ӳۡ���&v�9:q���f�o��s3�a|��2����:���8�O�̑��V*%�3B|Vݗ���D6�U�߬�~>��p���)����~Gg�4�.�n��t�f�s��b�Z�є��j�e��]w���UCV��ƕ�KY������UK���=Ҁ=p�Ei��e@��Y���>�;�׫t�Qz}��S*�x��j��7�n_�Mr�ݟ`�2����5y��>���_�nH��;�	�<�̘}Y^F�ֽ\$��N�o�r���>��j���ȅU^�r!��^9ު𕑾��~�V��p9�2�T1o�rSHz��� ��*�2%��J�+�d��-S�x�~ۄ�z��NmOYx+Q�h��{υr���:�U�S��7������\�k�:����F��]mg���{p���
�zT9�?͊���|s�8JW�2����ϑ�C+�l�����
�Lz�+.��V&v�yY����L�E:ap��1�����,�J�1�k�*���H̟���a̦t�q��߮��j�)F�����r=�G������PjmK,"K�1�$�T9�u��u�j�#�e�x%�?�B=���Z��/ǥr�x�W���OO6�U�`�)��d���	����Pb4rY��l�:Բ�P��qP�¢��0��V٨ ���\Bٻ��C�;�>ɵ�m(��m�Q��ˑW+F���zU�v�F��ˁ��zBF��D��^�iȅ�s���=��<����d@��.܀�8�3�i��9;�
�ck�<2}� ��X��Ӵ�;��?H���Q�f��Ag�\Q�F�s��S�=�	9���_�҅d��Bޮϩ�9������q޸;�E���΁���#�;}�d�,�T��p$�54.������*�]r���c>��Y�ڕ{��s^p�yvt*�H��1p<���,Ϥ�H|�OY��}FCY4�e�.TCÆQꢏ�F���^��μO���/���*=�w���F�'��먩}[�>��v��.<���P�W_�w�����<۫�x�@z}��|����!��^�3*�����g9R�s�:rj����=:}E��9}�r�����h���.3�LOg�t:�Ύ������FXhzt^FL��x���7�(+��Cn��:oJ񨽾�x�k�a�D���UxJ�߯���C�~15i�?�ҟv�G�yH;:J~:=qS�t\R��XY��cRyW�翆��3�}f�f�ҿ��ǝ]��S��Y�$ym���N90���nH�3��3pփϡ(F�I�m��;lW�=��4� =�[�_��Fm�w!Ju��h3��A�4��I[��+����T:���C]�3A��]o��'�޽�yV9�ڦ>���PG��s��q-^c�k�Y����B�5���V�@��s]�K��/�j:znj��Zbg�o�yUyzV����s��B�7Ϯ�ȳ�����y^�F��>�s��J����\�9\�:��Pc|�*1z��5��c�}Hxj�����>�"�Q���k�2��,x��+�����v*�>�>��muW������}#�ۑ��9��ׇt��9%�(R�{<�mL�1��(�����3�U/�sL��^¼���;�<v��Y�g�������T\�3"��������8 'Fx	���ۘ��OӖ�h��Ӵ4g�����ޑ���,��sT�W��&��=���X����	��@����5����|<3��lJڰj`���W�:*߷r��.s�O�{��~���[��f���H'�+��n���\s�***F+��{ӻ����y/_�}��"}�=:<K�� >�\K�]W�n�Z 9�z�4�d�b������3�W����ԍC�m_������}p����ĺ�L��
d�L��'#{�yb�;[�.��Y!�˾fY���p�	��n��1��/~��Ȣp�h�r�Wo\E��()w=�&0��*��1u���S�ob�p��V��@���Q��So��C]��Nn�T����]��r��]�U��i�tz��]�;���z�ز�]�Lm�0H��~�g?�G(�xz;��wro��/���� o����d_��!��@����^�O��ڃ�r�.���B���}U��]N��iz�L(}�Q������v��x���:��fy��&���R	T2c��և'�plS�'t��ʫ(�^쁑ŷ�h@��/��<��xR�G�i�Y����~�m����9���q�s���0u�_wz����w=S<�37�{��zyח�<������V��f܍Ϝ�;��xG�Û��%����,��W_zS��{��� yo��*t�FGΫü�_��Y�h^��QY������y: �l�b�{�-֔iz��S7G�y�4�
���������?q^W�{l/�κJ�CgW�{�ձ�B�%�&XT&P늙jb✄���׋��_c��Q��~+"��=��1�zt�|�7��o/n�C��4�"A]�`�R���'9��������G���f���9Wལ���ε��>����՞1��R����:H�<[;S(/cǚ(;c��C�	�U��E]�[�)�f�?�3��]F��S[� �l+r@��lvn\��i�<:F�G/"��z��Mi��7j�b�I:�zڶ���]p}ة3Χv���@�,ԔKc����if�@M�j��2��7�l-��9)����k�I��Z�}Q��	��2������}=7��Χ�i��RK�z����S������0[��c�5�}��u���m�/��.��-Z��#��\8��o�F߮튿z��n y�8�z*\��az�O�=ZQ�����	�Ʊq�w߭��s��Y�V�o޽��W�W�b�Ċ�!��~�¯M�f��fx�H o���!WR��܀_�b�P�W�/�ȟl���k15r=d�
������GL�Վ�����Zj��z{�$>m]ыm�̑���Z���ۻ^�9�;��j`e�z�b�J��)<�QQF<��=�*Z�ёN}������1O^A��=zzzGW�{�������<�+M�ތ���2U��}t���n�O�Q/z|f-M83�۩IO�u屑��}�5y��=��y�#3��v���n�C�FY�>��o����T�$�z���NF��Q{}lb�����ׂ���UxJϷݚ.=쭓��Aӹ\6����v;=�=cc"�0��D��z��=U�3� )s�~ʎ�u�j>_"�Pp��j�y����pQDq��Ѭ+������ ��;˗��]�3�K����	YY��e5 o����W�Y�B%A՟��ɜ��w;8EKwb?!�(��팒�d�j�>��2�Jק�+@<r] ��\���
N�E�fܢuky[Hs
��ge�5Ӭ�~kr_������2�L�w.���#�o�,�/Wx�q�o�K��_�Y2��l{��JUz;}�����������fX���ē�v)�eX١�]��ڿ����{��j�:T����+�ԙY�C֣݅�[�X�:QU�TT~Ґ�ͯ�{^��ك5���YW�������uc��|��j�����PhvԳl�K:�*��v|��Z'=��h館{p��c�r-{n&�;���zG���@���I߮�=���� '*�Y�q���2��G�#�ú�G�� ����T;�t�"����;�޲6��ճ]�Ϸ2���5�ޮ��J}��p���`_����Y �8�x2�I�zs�����l}�|���y���Oo����9���OUQ2G����*u���L_m�W�J�`�/��^���7y$����,���%z :��^���n%�zM!��OY��}Gb�[5��z�t�Ue¼{|b���)S���{�]ȸM׉�G���Dq�T{���ר�2O�S��Nd{�G��^?Z �U��W0��p���L�&E9�wN�G��s��$�z��M�g�ƪa��s�A�J�ԭ�tӮU�ۻ3�7kv���A)ڣep���j�V�a�a����L���^����̬�/�qK4�Zͣ|��]�8�ı�F�&�Bʫ��w<釳�"o��<���椨���~��>�f�ߐہKՆeX6�3Y�J|��i����z�{�KL��i�������+�ޠ=F�=k�w��o?x�JE��z�a9Y���	�p�
�twVRT�'M�i^5{}pԙ���R���UxJ���9�.�w�Ev��ޡ^���Fzs�9�;;s?���·T��)�N��b�ݐN��Gӥ�}4!37�(�x~����weW;Zb�7ٷ\X�s6 �<���.+&��S�<�i�����uv��@����.C���=���@�u^~������AF���.�����6[��ٔrR�5\���s�n�_�y�T쁾�19^�ӈ�SY^�<;>�{h\?>�.Q%��v��ye�<2W�z=��U�3�F[7G�&o��L8�O���n����ǭׇd�����r��1�㳱Yط�{)@���g���Tu�S/��O�3�ni���;��"|^��=�UhC��$ɵ�z��W��=�W�N�����j�sJ~���D�:v��O�m2=~�K�wHU2�wz�c�]8�tB��'W| �!��<�{�Rvò���w����l�uy(���	mZto�2�y�ҹ��>V6m_D^Ä�1R�(�27y�f3��h}j�K���M�@C1P�ܷ��}��]�v �eR{�����O_�޸;q�a�mO�� &`�@�=+�kc�#���eZ���\�u^�R)�Ko��Ho��\MǷ���w늿�MK7�T	��W���Q|}������f�ưOr�Բ��}�ԲC	����D� ztx�~�h>�dIs>��d�E0>��&-q�S�e_zI�0t��s�j�����}��vڿQ~��|�k��9�7�z���:��L3{�(փ>�ko���U8��[^3�0��J�h�>g(��^����<M�ɿ���2n=�P��n��W�:ǫչ50�ЭW&x�G��m9P\:pzJӃ~�{^q���˯.%�1��� ��T�����&NN]���)(=���m�l�w��d�Q����>Ӣ��;q(z�n�0��0#�s����s��*�uW���Azw�|gTo�*��gU?e���e~���x����cg�g�ɻ�^��w��Oy <����UN������d{�w�8{�nF�9�wA�g"�C���iA�H��^W+6����FF�+�^ O�|���^��1�xw��d������u�VE����s�ͅ��ь3���ae>�5z,J��Ub�L�c��%6�Lj�WJ+�1,wsI��I0�X���ZJ�p������:�c
}#������zؓH�*^�
�L�&�74=K�O-c�P��+[R�L|�^*v9�5���h�31t��u������Ԡ�@�|d)�XA��´��M�@�Z���P��B��Y/O=��+K�����p��g^!C;��-�L�6�	�b�2�i���9,p
�������E���Ey�V��\m�A/�S�Es�m)��-c����V�GP���R�؞(;�^���Z�Wy��Ք�i��g�b�F�u;�V���:�qIy7P36r�"CUJh��9�w���v�yo,��olT���7� ������:����,��x([�)Iq�ފ�<�GjTI.�-R6o9�RCl����Q�D��dҖ��j��U�[b�Zr�)ޠ���fs��pb�S-�5:����]��o�u"i�}�����z�A;���j��J�VNԝ"[ P��q�ذX[�>�Y�J�H��%��.�˿�C���M��bl3��`h��ul�2urwa4P]k1�x7���`^l�y5�F������z�%�:��L�>�P�]-N�����o7ǰv�v(#�u��I����ɺ�A�tJ\5}+0l .�k�!�l	Z�$p�ǈ�}s[�l��U���
�R�
�FA˄�Z�ӵ9���]/q�*�枳j����.Ӳ����wt^ö�]m��h7�m�1�p7>�1�+ȫ���ft{@V,�SY`�\��2�L���gI�����f�J���V���#����Y���3-��۔�%s�K�ʲ�m�O�[b�u]�.f�Pp����BU�w��Ԝ��ܒ��Le�t��Π���f��)nN�R��#� �Sض�-���\���n�d;ߡ���s%��C:�ͱ&���Խ���:%v�\dh���"�|A�����,k�����r�u���:rӺ<���n�֪2b�9��sQ�J���GcS�@㏛</��<����[	�B�pۧt{$��Ku�u��w���J�V��q�v�� EQ�`�=6^��HW��Ok�ia�5�l�T2^�U-��3ܾ��
[#72�0��ө��l�XK�A&���-�>��kh�P��w�}**o9�k��*4t[�+���h�&�089�+1����;bN�̮�����8�Z��Sɛ�ge���=�T�N���*�Zb67W�M����&p��Wm��$�C]j�[h<&K����NR_A�7펬���i��ぞw��t��R� .P��k�L�уX9�:���Kn�����2�dI�FY&�T�����J.��y@����l��j�2�R�%��+��R��9L(�i���+�#(�N��� �! :��+��ө�x��ޮ�>�y���1SM$�DU��V�m�h�*�(�)(h��"(ыcN�vV�DV�MRQ-�"`���PU��m�U%E5K,��4$QKE�SD�,EDDUE5DAEQDAm���bj�'lTU�kDl�4��i)�EEE;cMh�5�J�"&6q�i5AS�A�DQ��h��j�
"��DUCUQS5��Di�Ql`�mQM�D51[h�4�m6խ&��"�֌S�E�k4h�AQUF�EDTl`�#j�TL�Ui�;[m��j*����(�(֢)�2Qږ���#j5���������*h����Vڦ��������룿��u�i�}0]�<�k6�c��\{�m��򔢾y/i�u�>�������'Պ��0B�yG��!Ĺ���ie)��?��.�.�W
G��������x���p�VW��vG�cW��� �z��{}[;풇��'İ�L�wS>S�'6�k���T
�����C�����pR����L�MWc����'���k|m��5�H�W}x	ȱu*��>N{�4��g��E=#�HL��n}�*�!y��{�u���a�mK7�(���<�� x�v*e��E%��Ы�5W��=���u���W�[�z�ԁ�o��GdϏ2 'Pf:��
RP�Ky�6[��«�	����y�X�|^ב��Ѥ����m��ث�z��X y�+S=��K��[r;���ɾ���3f�)�Ya��ơ�~�ω�>���}޽��U��7�HEN��4v�ݩa8=�z��$��HU�R�����.5����M�O�>9���CF@	7�7�-n��o(��SXH�O])7�)���.{ƅ�zV����w��pڻ�4!)ؐ��<�y�j��'��P9Ø���d
��QX.c���b����9������S�ww�gM3 �n�ʆU�I�v\�B��ĬY"H������e���������3���#��E�ʡ��%�v ����=�N���v���z���cM��w���e^fR�ަS����ID��](��>�����W��kfZ�\�1<���W�U%{��{���^{�=3� w��"����ʁQ��2U�.a��'tú�n�*ή�lW |������~�+=��*/o-��W���P��3�a�O�do�G,�~��XW���D�]?0�m���w�^�T���^���O�ok��3/	J|9�Gz��V�o{�['a������מ\+������P}:�Ui���J5������{M/3�^��[�p��?*~bcN�/z��3��NmO�C�:t�/ L�WS�:.)����U]��^��W$�{z	�Uك�3�;�zw��}ח�׬��]#�g	J̱�$�#�NC*�l���l���M��bs"���æ�j�y����=~��?�^�=��#���Ƃ$���y�*���H�yF���]h�AQ�W�l�HO���A����f�'��o�u����9/)����%����F��@ǹ��V!6��g�7S<�}m���:w�+�yο���甑��~�Ӳ_��������p�_dN+n� ��0@~���~7e�{n*�;H�s�iO�4�����������K��<�Hs�@��ߘ~=W���4^֧".���>+$�C4�p0�w+#�ǎd
�u���7�u"��W�����H��i��ՙ�R
�zJ#�p����`����o�L��[�+���N�o���ʸ����m�Yɘ[�_�mq/�f䩎��ӱ���w������7P s��\㋧�_K��c���-��t#b���X���D�<��+�.�����@�:`�4.)�x���]r�𭩏R�{ ��S�勷�0#΋>�>��/ z� W�~�WK��F�Dz_�u�t���6Ϧ�0�L��޿f��s�S��0���6��t6���#�|zF�
�
��F�'������m�5u�/<�*�D�V}_����һ�^	��/�Mǽ~������	�YK�{�$�8qn~���K3����LV���[G�?@��YF�/Ui{�����'�޺��7���fR�C����'k<ze{�@�p>����zN�ǯo��>��)x���v$�������%Y�&����'9�Μ�����@���(�S����ج�d1>��*�^��tPש%&�v�*��?Mx���Zb�}�u�!�'v����=o�
��x�������?���~�������E������+�67OG����]#B�K�3Dꆴ��ǻ�iAt��^]J3+dd,b��Oۛ٦�C7R]T}w�7}�M�(z�
C�z}����#ݔ\�g���Z��j�8WWzp+�Jr�*my�o��s쎄���Z�J���uN<%v��\J��p�l�lt�cb�ԕ��u�wQms?�B�S÷�ih������tkKlr�\{ ?M�d��j�
5������=�ǔ�������-���Y(��e����7�eE��pN.y��2����P/��L<�ޯa��no���z�xqwH?u璱z��ۼ]u��d�G�%��{��C��nb�}I�fY������/����)z�t:�_�Y�k!�>�ws����z���@��,��	ўb�|���S��[u�mӴ4[���n}O���#������[�~4�]�0�{j|m�:� t���=+�jz��ӎ�n�6E_ ���p��z�2=;��?Oi*=���>��EoΦ���D@j�H&
�u��P�Y&�f���O�H�C>vz��^�]�<.�3�O�����m�ՠ\���7.��7�2KG389z�G��ǣP�G�Ͼ7���Q�����Gڑ�w����R�5�� :�*#޻�3k ��Eס؂%{;Hy�/eT�$�O�M��}Z*�*}�t<;�w���ɻ�7�9~&Mǽ���w�g(���]<WD��hW���)*����p:pz�V�Ok¯e鯗^\<K�|ag��[�bC��ti����lĐ��,U�Nf���3�]�T��;�T�rP�&���)�NY�� өw��u� �4(VK���ǔ����1��t�m�(�U�˂�
��$U�u2�bUmv���t{04M'f��"p��wK�P2��9��ip�p.Dˡ�vO_:�[:�\s�iG�}� ��t6�<��7�zA*�L5p6�;��i�qNt���=��Q1�W9�{*�n롣Ѯ������"7�_�ET���ɜAUO�`6~_��b��o�!0S��]g
E��#���/Ksǽ��)�&+=ֆ|���9	ח�<������m�H��Iݳ0���G��X���f�f�!���Kн���h��L+Z�.z���u^�;�?m �{m�|먫�����?b�����L�A��wJ��.����
��
��x���e��Y�y\wj�@�xg�����Tg/GU<���c��>���e�Bg����r���^/ w�Dc��Q��qpO�����7����������}+�3�����ȱ%JS��"��s_��>8�x�uo�r��y���Ȉ�P���Q�o��vԳl�K��R$TKgv���9��'c}�q_���%K��:��F|���V��i��RM�_�=�@��`@L��I�)�X='�/Av�6����ǫ L{�b}q7��0��#��\8�����]��L�N�k�`X���������ZX���_SX���|�x%�w
���I�F�f=T`�5'"U�q�z^�69Y��U���Xp��fm��Tw�V����)�Yk/��o�\0�}�I
���Ί��^�H��D��Y{�.�c�ܥ��ulT_f�q曅�w�(���\}7�k�Ąd���K���0��ظ�;���m��}����A��^����OC�a���AK/�c���Y�K�'��T���$���HUԾ:7 �Q��;m_������l:���~˫�7o��e��D߾����H�w^�q
d����K��q^����;ޢ��0.�Gލ�wf[��]��s��6�>����b������EQ�.�`���~�>�[�7��}n��k��������{C��yUP�F?P��ǽ> ���V��FT
�e�*(���a惓�\��NV��W����o���E^�[���z��_ў�zr=��w����9�0�{۝[��^������1ފ�H�����{���cU='"��w��'��x6�&l�	�[��W�����ş����t��]�ыG�yU���(�Fb��{M/2z���l��w/z\����=���{�|n7�5�U�GN�%ᎂ\%���O�~��KW�]�����O�/s6r���!3��0=
�k�z��w���Y����r����2��,I>FY���3��ӳ/|9v��à��ee�[�H����M�:m��85`��ٷ���R�|��*r�H�����:�v& �c�Ϯ�,�;xE�&j �eY� ���wU^�{:��2�5س�e��N���S�l_KrB��f��7����*��Y�,�gj�J���{�W Wؼ=~���VDW�vZ�[����*�3F�ʦ)x�} �s���c����|<��WC���z�f�'��o�u����9���|;jYa]��Y����n;Ԯv���E@��g�n�P^9o*B�~��^��=���n3ʈۇ�l,����>Scn��˷����N�� �����x�v�����m�[�i.w�q~#�'~0
����T�+w;�Nm23޺�j�U�nE�L���?J��5��<�_��U�|<�ś�Bo���M��A���p߮Ϫ�dlK�,�*��O�
�N{�s�|���h�L���H�~����yN�zG{�r�*>,�wļ����~���5�6�Hj�M�}^��y�c��]�Q��΃�����<B�dx6��6�Ŀxπ�dq�W�.�R�_��#$������
Y|}p��5^�D�RӔR;WP���m�d&���c��z�c3Cn<��
���Ҽ��޶G0�fg� �\l��WJ�L�i�����Q{yp��^�������]1<�j����?
i�r�SU˚�5�2�n�H�������aDs�̽΄'<�M̎�q��ޝ~�|-3MQ�J[��.ss
��ę��96.�T,$��	���VQ��Dt| ��5+�m��<��s��
��{:�U���ew�3ح�;��e!%f~cg�u+��0,���գ���m{I�zW��uC�S^�����qbz��lf���G��(Oz?z�~�k�|z�gI�a��*r��G�9����� �� ����Vu.���3}lλ���z��#ޚ�K{ǘ��&v^�P��ڼ���~՚��A�lxQ�T����qmx��@L-��B��pΫ�ҷ�]`�9�m!{��H�Y�R�桧F��e�ٓ���)z�U3u���ڡ�k�*#��Mo���R�%�oϮ��W*��٘�g$�U��K�Q%�DIh��ȣ>F�(�	�}T�χz�c!����9�u��^����6W���&Iy���xt얊��3�L@j��L�1u>��E��e�a]�/����r�{�����2'������=��+��}Y��ӢY�p@N��0�k�|�Ē�������q�kK����}��;�z�=냷���y�S�� � o|d�yM61�X�\E�w�뵷��J�x9��z��~�����\N��߮*��Գ" 5P$�E����03���[g+�]�%Z-O�bm�)�7��3�`?	�8h��{�g�O�Rp!�G��]�V=劲"�)WQ]spk{jݞu�wr���
+�v���},B7-�'�NT�fs��c���������Y�/m25�JJ�� EÓ�	���]�oΘ�sĿN�p���."}~ț�u^�=�-����:�lO�,zNa i����5�ŤfD6��}�J�Ƽ �`u�z�dĵZ��C=W�;�Y�ު�����-H�C>�բ�������w{n%T�2�L���{�j�7�6{����1�w�꡷ʎKՃ��ς�6=�+N��{^{/J꺇�edS�WsFs݂{,���6��f=��W����p\?]��*8l_zA*8�Z6�9>Ӄb��;m,�J��r���d�y�������1�}ʟdd>��=4��{�����np���j�*�7����tMN��NC6u��y���p�s�Q�X��S.�S�sＦ����kǽ�r7�;��-�ꮷ�&��g/3UR�C��;1�uXd$OtF׀��+�}+�9�}>~�A/e!�2[�w�_��%�Q>�w�/ԗ��QD��(x;2���g0oz�9��f��*,�W�F��rwm%w��{���|뤡�B*��aA<EL�LK!�[5�\��;3�m�x#��/��<�2�]t3�i�]=����x�eӼR���%%c���΍��x��N=+.��)�v���)��V;���"��:]qCq�0� Έ!��G,8�s�;7k�Ю��؅���L�tML�εw]nAŌ�<����k�|�*��Ǌ����L���Q���kҸ�9�� �c�y:*U!qU>Nq�`~�s��d;�g�ɮ���ŏk�S��=o��݅�w7*Q�x���������fi�y�	;㦛����cݖ��$_Ο�B��:��<z��RK�z�� vԊD@�{��g
�w���/c�����@Q��7a���'��X�y>GT?To�����]�}@��rs}+������J}��� @k��@����`�|qt���m��[,��A�B6=�bw��O����������M\OU�p�O� �?O	��V����.5�~cB��2.@��qw�~R�r��='���"\9�=�e�zM���}�s�����#Z�zI�j�M ������EGJ���^�+�0�����;��2=�4@K�^�p�yW�z�W��o@wf��S�#<=�칵u��^Ɍ��x<3������z|y�N��e@��%X���{����ɨ+�<Ge�%^�螥��(�=��W��������J���x��Þ����\y�}�Bi��i	�1�wz;��p(��])���֯���֮�6Z=E�3�.</��`���da�V�bǿm�Y}�v}m�u{10/z��t�Q�͏��[!�������}@����&u��z���/v����(vː՚2%Ǜad���9��M������3�t2��m�h����Ӳ*BrD,����4�L�k:[�d�9@ŕ�k�K�-����KJ�)ȣ��xn�;n�b49�Qd��=�h҇��J� �B������"]��77��T�[
fw�N��d�}u��<���	�J�SʖH�JC!�ϵ��St;]/jo,Wu�WO6�:z��:ލ�V�f���4r�#�z�PV�����������Y+xnN�W8�8kDnb��8�o�!�&��Y,�����<m	Ym��Et*�npҡ�,�i͇a���u_�m���Ce�#T�:CCUţ�Y�V#D��J<�z�}���PUk���5�)��$B���)a6��t�f����4��=x�ܨuK�76ud&�:���&�Gq�Ȉ��gi���nc�]�5�[C�G��G�>G�e�YWޕ�렗��� �f?V�-T;\-Ll`��3U�=����:��*�JZM��"v�-��}i]���%>���I� �]��
�\����q-X�\��"��G�*�A��[hP'Fr+S��i��%�d�R���r*R��&���6�ܩ:�j�FeЮ6�	�Vei���xC��"g2d�Kj���sC[��Dך{Dy����Yz
���"��$,���x��,���*��b�C���y-,�q$��Jµ�ϴ���2���<zl�t�QNޞ9ie�6�Ť8X샘!�|�g�Nf�����b�t��-Nʼܽ=+�L���]�Ŀ�x/j���^g�q���0̻T2hY�2�:c���Ff�#�l��.U���РaӴ.�k��ګ��,U���m��~J��i���ꎅ�M����2�+�r�S��kq����c�ݒ��0�2sZ�Wz�BEǰ,��b��P����뵒��Z�E���YiV�Dr�=3R6u�3�ֈ�eu7�+!�n��C�λ-#!L��jTM�}�A��\skQ P�0��Gvk:���Ѽ!
��{Ky���K��h�᠐[��&]^��Ne��/����\zZ��C&:G�[7��<�lw��KV	m�P�Y�]���nl͒�e��8���5��ԝK.��,���$��]�u��B|�P�ٙ@ν�V�3u+0✪�ʘ�sG�W|������_\��E��k�k[��o`\!��/^\����T�о����u�A�)Ae�S��ͣs��]�4CWLsϻݶ��9a:N�S{/���u�ERW%4	\��5�[7�V�kW1o�a�$��L7���X���P���EAQ6�X��ƒ�����'cZ�I�Th1V��i53�*�KUT�6�Q�IDED���bو�R�QDU0U)N�QV�(���EKZ���m�*&(�B)�#g4���Ui(50P[)�5@DkQē���M�����K�5���Ĵm�X(��֦" ���i���J	����E�El�m�AQD�,�T1LEUE��)�J64�Ej�Ѧ$�"KmLKDA5A���kQ1���[&��*����Z*��������
)�v��*�m&�CT$T�ER4�N�HD�-1��t�*i*#Z+TZ"�+u������~�>]�}����2�l:�:�t��p���߯��sAY7�rE����N.dV�fV�����ASt��}i������n�G_Ք�D�a8o
񨽾���'>�#}U�<�"�y��;��r�W����}�R�k��z7�['qL9G�f�ⲫ��^$Tap;=��U4��9�HD�;&�i1��5��Y�����3�sת���}9�<�6f.G�����Q�qNG�ޖt�.����F/C��B�[���������Vǯ.;�޽�YUǬ�=��x�O��fy��}�Q^������W^ߠd�]�}pb~�	ϟ����R���~}t."�z����1��K�ϋ�=�;�U�Ǫe�qG�w������^�3���G��~�=�"^RmK#���Emǽ�[�^�>�O���<�7(�f����[���~�ϗ�y�f�����ٕٲ+�wN_�ک���w�~��:vO������S<R9g���Y��NиNw�q�3ޞ���ͭ b+'c$0����Fں�n#ޝ��pB.�d���x�V����pw�`̺���o�D�+Տ0ǜ筌�z{I��\���~2.UK6�W�$��W�hK=��NUMc�nB�C�M��L~�wJwi�[h�`�uGAF��Dh-���#$g���tV�k���&c��	��A9*���ݨ}�3��cG;��P�s紮Zw�
�1I�1Ru*�:�iat�F�(��46>������a������T�K��|�^?O���'��2}�_�&�\פ�ЦHj����/��ljq�J��-t�裞٫��TB�dEB]�q��>����@�z��W�����tp��ޮ�]�-��:|v�*%z�\D�3�yP��w{m��7W'����z�0de[�N�G��/Z����ܞ�#�����ӭ�Qz|/�/B�ˇ��w���Q74���v	>س[=u���<��}��7�6�������c	t�?�m�i:o�+���Di4[��?RݠOor<UR^�1�I�/�τ�����k�|s��A�ۉ��T@��Q&�J����[��i�g�z�7�<��w�!�2�}	���=����a}�ͺ�8Ne�fT	�/#���.��E�(f�S{�{��}PN����ZZ�/d3�OՃ�罴�����9��%!��ϗ��{�'յ��*{�z2�������#R��Q�\��rt�魈�SY�B6��m
٩�~���d���ÏR���!�D�}Z4fa�I�q�*#q��鎌r~���7����J2�rfh�+��������"oи+�y���ķ��Ϻ���k�-����f�������G�G�֫N�=<�9dG���a��D�mqt��s��w9N��`I�p��SQ�u�ă'
�8�M2�<�ze�A�l���S\��j�(�G&l��Yű����Ӳ}nP$���$yT9%ɟW#H�2���>�׶=�wW�9n�mt�*WY����#��a�g���	g�0x
P4��������&<�z�b�y�Nos�'κ�47����zF����)��x=�>6���1� �@Wf�(�U~@9��s���H�^t��^�p�Cפֿ�~��߷���S�fYH�>q�1b���VN���)``�ި�'�y��ֶ�0��3�=���&�~�h>�dO��z������������} 1��G�)�!�K���Z�[�5~�~���	��豗:���Z��VM�Ȋ��`~��ރu��j��,�aқ^%���/Mwz��j�N_�|�dݩ��ܯG�9�W�&O��*�@u^Tl�^��9��\�vK��W�����g����ו��Ƚ��4��������z+�oޗ ��H�)6a}ސJ�0��ևu>Ӣp!��o��vh�����wz�h�%�Q{w��^�}�7��fw=��G��s��A9�W^��sH��R;�;J2ԣ��zr���7���B�Xg�7��;�,cn?���6��/[V�3v�j�X��������!7�����g.;��0h��4	����Hc&�s�L�ǘ�v_u���.�L0lҊ�=����2�]�͒�Nۆ,�B�4�9�t	���>G��+�E*|n��;mCY�2S�9�z_��������nF�g�C�&X��Ը�{�s�q��f�&������@	�o����ԼF:��~�AE�!h�_�[��z��n6=흓�s����9z�_��C��;\������/?�>�o����~�γ�	�覮;���_{�t�2,�Q,,�3��>S�e-��[��X��>�o�Z��p=�v|}G>�����]G�)�:�+�3�jH*��t��X��
w{]��s�q�2��K��>�DzR��#|���7��cs���~w����6�Q�x���1�Ex{�����|=Vc�9>�དm���FB���Ϸ�<z�ԁ�o��dڑ�/}�3�PB��5��_��@���~7F����%�V�����?Lf�����}T���F������x�ߨW��7��F���@���}Y�|j1uC��m����l���-'��3/#�Ў��>��뭉?ş$O��EtH�~\����r ㋌ç�p��;9�,��j����ߣ 9|�_n�A����>�����ȯxOH�W,u��{UBH����&"��~�7����=K/�*'WF��|������}���7f��o����`���wZ7jҫ�h������݈��r��-�8vۙ�m˩Kb�b���k��|p�sĸ���U��t�#�"=.�;yw��e~�"�伜ؘ���z�_y3�\�ڪ��Q����@u��F��^�hǕ|'������f��G����֔I�h�9����������K�t/���f�ޟ����i�E�^�2Q�kr��Bc�:g3��_�v�D�����wJ+*�;��W���P�������^��s���jJ?�maɼ��!{�@�T�"7f��)/	�xW�^�Z���S>�~h�:{���T�5t�<�pIV4&����E��V��S�x�}�\n(�*0����K�k�t�s�2op$��ָ��N���;��w���?��ϻ���i��v����2�R�)�}~̺�S��"n�kSK�n����v�����{�u���DVym��,7i�Ol挌�������;�v��Շ�^�Ǯ�,�k��?_���?��C��1�?>�G�=:�O|��&�ȉ�J�g�eW��S:��A;}ty������{�s�1�*^Rt�S�+����19Uo��N��
�e:����O�c����:��}í�����U즎��Ȯhn<�0�up���X�9���{�7*5Ƀy]�	�7E�%5����gײ�-<@����*]dɦ�,!8�w��s4f���iWT���i�{[|���ۛԞ��"wU���=n�c<�WT+�2���e�����_�s��s������\��>n<��P�6V�s��>���-���d��r Nj$�����#tg��Şۊ�N�>�a��D���[ۅP����)D/H���?Y�g}��|m��@��@�{Ǆ��� ۀ6|���nP��	N�<��xǍ�0��{I~�AΊ�ߌ��UR� 5�$���B�˲h�&�_����1G���~�S��܇p��<|�����p�Q�*=���ܹ�ID���T�]�X�.b���0��B�_#﮶UEv�\l�z�+"�U����`k�wG�wE�yR���M��|�O��:�6xw�֨�X?#����zk��m��	��7�|=7�{��8��>�T�#�f_���%���ьm�JnJ�����g���n����hvv!m���^���s��鍕��w�w+�� �<���&�kc�@h��T�
��W��zNҼu�u	ڵ�=��W���1�c���w��{Ld/z)x����V~�q?�Mxώ|�H;;L�
�Ώ\EN~<�V�^$~6�cg�Hz��0s�N
�I���E+c�P����^h�b�����mk5�Z���h>�֐Urֆ��d��ާ�Np���q��q��P*[8%�*-{2�3�J� �F���j�,6�c�॑/��6V���i-����&]�l���J�;y��>���_�z�7=�gʩ�A��k�";�^)lw�i��f�i�gIݿ����iW��.ʊ�ֆN����V�S�e�E)�7NP*��] F���@�u^�J��Б^�Ao�]#���0#��O:�/�tNw��{=0��T�Ӑ<�g��@�@rr������ϫև�l�Gd��kc�����`����{.Q%�-��T;������&m�W��ޠ+�_�;�r�yh�!jS{�m�R��}����WQy���Op<��L�13�L�E��g®6f6~���nzK9����s���9������ݐ]g�� t�m� ��<��h71&=�u�t���l����V�ϥ)�E�Z&�z�4/o��q�z�<��Uxǐ����D�@{�j�t��}DA���k���-R	�������q�����۸��3�n׻면�3sDz��2�y�6�$& �����	���$1m�����l@���n�Z+�9N� 8>�]�R�N'�K�>��h����#ޕFC���\j���o�� }�s��A�L�l���n���VM�m�vJ�֎�W;r�6��bX�Mp#v_cH|��;6�"K�"��
����"�8��v���,������/x���gw���g13.��7�kd�+�b�y���T�ǖA��Ϙ	N}Z.��S0�6��w��l| ]���b�5�SYl�U~��S%���M��_W�\T��iz{�&�����{�>P��T7�V�r}��&K����
�*6E/VR�7>
�N
�+N�~����]3ҏ����W<��B�˅�����I^����~Tp�QސJ���mho�v{�^a�����Q�G�ϑ�>��x��^쌇ޡ��M�=�TN�;ʛ/� ��~�_�G�P����{�+�+�+)#t�Aݖ<:����UN��N��9�yMWN}���]���� �v�+�����*.�{籁�D6�,,����p�$^��`��W��x�u^�5��9P{���d����_�������ݷ�^�����'F���A��W_�����ipk���^�v���}rVF.���_y�:f5�?\w{�l/s���E�Q,^	��g�b✆��}uv�'��M���S;��@�^���9��W�T{W��#p�/�x� ��>
E�s��ˌ�@�.�(�����P�`�T��r-M<�������cs����q�ϋ�F@�e�Ir~g[�Z?�t/8~F�b����ޡ�� Y�@�]��DԘ뽶o����E�[Y�տ����Jw���|�"M{,vl�������R����^�Z�L�$JL�m蕽ѵ����:4u��f�TU$d���]>�ү��q�;�=�9��\���Z�<Gq�8�詟q������#�?^���3پ����@�~�Ty�ny_��|��/;�_r³Ӈ�2 'Pf: ��>�̓N�w�q6�C ��#���{��<��뽊�]�g6�F{�v�ZUS�@	�D��~-�
���Ud	�ƾ��p��^�Ƚ���nߛ�f~�*m=��Ow=�^�uh7�~�6�����˪%��T����:`/RqR��n|�'z6+f<T�Tǽ��s�����W����'�x߉q���_���U�7�!��V+�s�4.�wѬW��ex�\n%��b5gx��\��\6����6�g�>�L�{ :���z�����0��1�ބ�������?�F�VE)Zj��6��^�ۻ���ʈ���w�;��qތ�;�}3U�253��Ũ�~2v(�o��WJ�M���vu1�����3�����q��iy�����|K^���_������L�R�[�+�2[����)��1פ�������k߅_s�^y�'k�����~>�U1=���E��el��^����f�ߍV���;�;�\�����g�	���3�?��"�yd7WYkg� ���K;h�H͏�vV[��Pu�q�&WVm�NB��5�vJxY j���\�O�Xӿ6��9,74lU��Ǒ�2�.'���z�h�mM��6�u�L�=�oL��Aض�&/*l�*�:D��=��J�����5��>u������"5�x��O��t�,^J���:=��X��Vo�<�1ex=�Da@-�;�k�D:���������Q��|���8JW�26S��h�ӷ\s�6�N��=Ji���*��,� �M{<+}��VEz��8�t?>�G/N�*���4A�Fϧw�g�Y�_�3}<2�|�Ӑ�}tx;޼�x��X�8�����D�d��^ �V�er�h^����% >�n��Q.|9[��P�_�r;�<痈�������tS�J0F�R��d��� '='����Kf��(�o*+{״Ƀ^�[��w^�~�>�S��w��=g�dm���~��"��7P(^�*o�D�O����Ϧ.�9�{~�>�J�x�Sfzs��~=������W��d[��e@��P[��q��Skz�P����V��
�\�m��c#��g�>>��7޸����^E~�U[)�Ѿ����j���z�ہ A��]F�횽�s�d!p����Z�e��
� �}�D}�G��>�AT�*""��U_�*""�㊈�������
"+�Q�
�����Q_�*""��DE��Qʈ���Q�@DW� �"������
"+� Q_�TDE~��"��1AY&SYvPSqL�߀rY��=�ݐ?���aK���H�(
��
�($����H))�*�P
��
T"BT
J�UT���UJ�
�  A�bsrUR�$$�� �T)$��T�U)QU)"@*�"� �6*��7 ;v�%4j#�S@`�ʥF�mldSb�#cC��
��T� �IG`�*C�   �\  �  ��� 2�$�mm3T�iT�R�*���RIQ��A�P��*��(� 5Y�h�i���%2�$DUD��p ��!�6�m�$A�T�jج�2���a�(��	i�PU���JU��%��uB��RQckJ
�Tڊ�H�d��)�j�P���։1V���U*��. w5RiH�kCU,QR�&�U�&�)X�MR��V�
m���@���J`�#l�(�\ u��((eJc`i�֒���J�&����RH6���BY�)@P��� 8#�T[Pa�h�V�[55���T
�63l�ajh�QR� uH�h�V"B(�mA�mU)�H&�
��Rƕ$DI �p ������F���THBZm�T$B��Q�Q���ʑ@H  �&�1R�T1�M2d�L�� E<0R���@1�� `�"�ڌ�H�P�G��4��d�T� JT���0� �昙2h�`��` ���M$��R�i�!��&A�8�WS�]V��^y�9e�u�Z����V�4�I A���"�q ���,�D��鄐Ar0�)�U�rHb�Xl���t�e~/���T?z6�R����  ����5Y$Aʈ�T%U$� ʑ�ϗl��O׿��]�="@A���\��W��д�:5��y�l��+�-����,.��s��������s�í�˷Oozk���TpR;L��gŋ���R%_]cY���Q�n���M>G�f���������)�X�2֘ad��)�/r5��o�����`�Y�M�LG8
V�]�b�46��oKj^J[W�8޾|V���xX�3��#k�����̙��Tҍ���<��#"!T.%eԘL5t uy�*�����K�u!���F����[�A���іim�Hv�1��}n���gn�[C]���V����a�9@�_76�8vj��يeR_a 楘OnS�������g���Ǎ&�݋%:O����J�V�2��V��NaN�V3�SHH��af-	�b�q�
Z��.f��3��h��nV	��%v���z)4N�n�tᗗ��m�0�y������ڹh��A53p0l����gU4���|x����G�G>���u����w�ZR��n��;C!ߎ��[�^�R���4��we֭7�.�M�t�N���"��V��L��t`fu,Ú��/i�`�[D��B��r�öBݪȚ�m��towB�D6��Om�r�\�i�"sE^mޠ��FۋU��"nf�^U!����X�������"�gJ;L�@}{s\	�,�B�#Z��Z�Ñڲ��R�����gY�aٹf$Z������,�LeY[s3$�Ǯ�1���1KEm��Yǈ@�F8��m]Q���&�r�ɻvR����Kf��ȥ'�W�e�Emģ7"Ճ8;L���c�1��ѕj�oUB��J�A�s)`�q,&�V��d<ľ���y�r�.�U��L���Ё��[�	ʰ{4Wv�V���IY��֣�;0Pٽ���w��w�'b��CxѶ7([�Oj�MX��r͓[k3)�2-8���T�5e�6/.]�L

֓�s�VV�zJ�2�:�s�Z�"�ʸ"�%�i�Qmh�ϲ���|��+O
�}�D�J�(��S�`n��Z@݃raM��a͍���3����
��O��4���}[�.�j��8�+�F�ea��:���V�Z�b���н��Ӂ��z��(m��]Ǜ3�I��n��z�V%$F�x�IV��eۤM}����3Z*�F�f���f�ڨn�6H��D7[�1gRt���Phr�<��`㪬;ɲ
���nl��]f㩶��U�h�ǻX�%%�.`��fP��ywz�J����,tv $���PG��Q�A;�\�0�KDl�͈�Wy��܎�84:�A/��u���� Uޮ�v���tQE����Ϗ^��d�)�@�c{hn&{��i�;{MfD6�9��c"�۶R4U,:γJ���*��M�x��{hҬ� {��,��B՛�ˊ�a��Z^��e�i��h�:��Jynj�doU�q��LVb��ʍ�x���l��v�,%���nCP�㽼��g
Wgu�VeY6���vغ��!c�n�kC{.�����ET%X��n�*Z�Y8�ݪ�-��9��*�9f�J�e
c9�T��1�!�e��ly�ރV��� ��WQ��85X�&�˵�f�yե����2n\�S)n�C:��t-���h�5D�W,�:r��E�t�Xê��d�oYv�!���]=oV�勻��XY++q�;Ff3��@�q�PVؿ�f�I _g|��:��XyVX�}`��UYy�Z�¥���.*�� 5�n���.9�8�6�����fv���Yw���e��
U��坦Vp��M56�q��LZ��ݻ0a�C��ǆΚ+Z������M�6�Z;��PX�`=ڪ4)�/�R�R�f,�iF�$+U�]�a�����nn*lf۷dc������9�l�j�b�3^[I����Xw3b�H����SJ�2}2bt�䛥�2��	P[M$B�.��U��j}�>�9e�;���͡��l^��3�vtM�kw-�j8����f��mi����
(���Uf*K@��,<�O���h���^�� �k�wgZy��nP�/��
�"������c�A�e�ƃ�f���uMR�~��S#�SB[4�U���a.3z���Q�U��D�c:�
7�v�u��彶x2��뮞��0v�������A&�8��Ţ �]��3C�E�ˎu��}՘�</�V�E5��0�����o%d�x�匼H��� ǵ�16�V�����X�UaKjEJ� �Pҁ�y[R��Aܵ����h:w�ճuB��iC�l�cXUI�RQX�a���9n�{�H�n��vh�n�0 hF4���Q�D�(dǑj�9W�3	��I�APu7(m�e���ŵ��2���j��z����*��E.�[I��ky�4��re�G'eQ�,a��=�ۼ�4)u4СOnM��oé��eib���*奒�0�f뙲ڪ��"�JUXq"(��q�:�:�6�4Ԫ��U��m^��ɕ.�VGO�uJvr�v�PPo�㴖i6���;�{`)�"Z˹uu�c��%^��`5gsX �"��2�f�6K�j��+Q��d1�:t�Dތύ�mU�]2���`�j���	�#2#�*/-�1Zٟn�	`r&L���uB��,��w�e�Z���Z�#yF�������g�ΰ���O8
TC[���Z}��Jc
Z��j��Y��I���1)�p��l9��PY{�����6j�N�M+��wX�]��ٜ�S<lG�ʹ�����7C{�r��Y�
�m��
#TV�����E��9�9���Z�V ]�J�ZŁ����������q�o���KI+Ss",*�bX���vE)�e�Enl��B�h@�hخɨ�ĥ�6N��5B&%i�����=Y��!��rEnK?�r�6�e;2(d1�YN��&MӃ~']^���o2��Sj��nٱW��1�E�4�2_[�V(��[v�����l�^�Z��0���Ƹ�,�Վ�2�Q�蠅n��*�]�\�m�a56����+X.����,N����Skϭf��tR�x�ѕnn��X"���zc�R�4�۲�Mx^�%��a��j(�r��
�^���/m����V�&�,<_h���v��)+L֓�#��Nm�^�[.n<�������t�	=?^���{�^��ڑI�/C���5\T��X�feB�jZa�����N��f$��XFl�2K�ȼ �MU�e�"F*E}md�/P�UB��j�!5�0���3-��l�K�r�qokŚ��u�������ybz@�kxc�����khG���-
���Y�>˫�l���ѷ�/�nR�4cL,h����w h>ᦐw�ż��wo1(�֎L��港'���42����6�PԷ�+�7�m�)V.���U⭻`x2+r�=��lL�f4��F<z�oq��0���]���\�6����8��jY�L�mR)����3$/ub���M��s���|�����X�0Ib��t %bF$�ڻș&��N)�uQ��nc�K�b��N�U�D��B��]�ȕ]험ӃnZ�{����K��N�cr��sVm�ڲT&�9��QJӴ�7F�.��M=�:�n ���^K:(�#����ݡefcJ�
��Ȳ-;)A���.ʀ�����������h�Ju)�gՅUS����tf.c�h��N��K�`%v�K9r���+/�ڹ\X���`xC3.];��b��ԍU�����U�kF�z�5I��a��T��X0��cC�|�&�7���� �.Σ�v~j8��Ry�2ΐ�열��'��t	?3R�(MJ�hJ^��o(���z�+Q�T�	�#(=��������ִٝ�Nf+��^Y�RT��{v��n��1/���DF���#�W�z�{�y6����r����͜��t�Q=�	�`]تʃ6�\�:�Q���ƦҪ���L��
��R砅F�n�sr�
T:Zy��a�f`�&�LmuR��9	�]|�̮�s�����m��E��Lo��(9�u�K����sN�X�4�r��5��F�	.H� �O�fL|-�Is-q��FxME���B�	U�����*��v|2l(u����h�@��<!�>�>��5�F������y�#<��A�{���C�r~��WMk,ٖ%1���Y�elǻ�y�hjn�Sǲogݖ�9�e�+ي�ROv>V��w�x��V�f52���#N�fK�c�:̛0�;d4D�\lŬQ��+T�����O��̧���j9�
��;!L���҆�QcP����G�8�e8�zƷe��ɀng��\�9s����}9ܕuט.:����R7\�#�����.E�d��O,Zֻq�M��Q�bd"��qZ��Չg[�+K��ӊS5�!�k��-���6���拄�Ѵ��K'�J��9[fX�q�)�a��J�r��KLSTr�̣$vq�	y]���2�U�gV��ɬ٦5q}3�}��=�m\�o�"�>ͬ�55�r���ǎ��
�{q�N����(�m�������~N¦��`�Q�YF���\�x�SwT��ɒ�=V��sF=����[�rf��<ث���b����'���`Ze݌SF���1��V�L����x�8F!�6/��n������r���i�0e-B���;gX��}0@��u�>	S����C&s���\��Uޙx�.0�@m����{�X�2(C5�&Fi�� �qi��X�w����3Ni�sh`�"�r�5�`��,ُ��	��.#[\2�;<21�-~Lp����Z}��cfI�NL�9|3�a`��mE��Pɼ�n�z���Rn����B�(t�k^�x�f<���{�V!��8ce�N_5y�䍚6��bb{ku��MD_$t�[��z�A�޴��`��!&�P�5+a]{��:Z����H_J2m6�D�k�͘��s�6�$��EJk��R4+_f���ǟ�ѐfcr��v36_F,�E�&dΙ�{b=��:����b��z��*��K�q�7gEqwVZҌ�d�!�����S�W.��79�E�F���zgYj� he�4
��bܽ�iG%�̘(�;Ў�$�M.|�̼���6�t"��5�MŇ�R9w�]%+0��U���Jqu�(=� �X���8&ɼ�.��ĢC��ɛ��w�(� V�e^��c.��Mq��e�{�^�)���.�9��\�]�,���W[ �X4�PqB�M��l@�A�Q��m#B�uU�O���Nbaڢ2����wk�K|��f]WR�ј�KK�����!�/�K؁}�1�+������h�����ܚ��;Nd�;`*>UB�v�1�U�p�t��#z��x�,�Y:n^P�H�Z�0����q��u��fv"��_ln�Zц�F�PB�Td�ʹyd,>��V�����4:��WU投�a��(��T"i�u���2�����w�Q6��]�$���QO���?<��)X=��p'ie�Z�A��Sq<NM�Z.Ԁ��c�@��/��,"wBg��e�^�<mSW�.7٫l��|�v���f4O.N�gOWf�n�/����k�G|Hb���p�wP�R+9픋�{�8��lW�#��::(und�׹d1�c�R�e��\�6l�٥���=u�~P�w4o�����eB���5�-ӑE��!.�^�A��?�di͚ʗ��ѽ�(	!Y�w7��U��5+WV�ۛ��� <��U��^�v1�B��&qV�ELe#�ܤz��]��)P���!x���Pś��b�!E�gR������ۂc��	��B1PGu�fn�Џ7h7}5i�,nZ�t��3Ә�����sЈ��6�̺%#<�&�×p�4��������T�˟�/��P����셝��pj;.aqc[�|�����%�m5�S�MS��T�D�^���\8�'NLe
Pc�e�2����E��"��-A��Z�;l>���4Z�J�ܷ*�{�љ[3u%7�%#�ٯ�D�q��vg+��K��ſXb�%n�2�hܪhC[�V��ʙ�0=��6f���޽kqꔊ���vnlG6n=v
p;�&��s�;���T�.�ʼ�|̡`�˝!�\]��2jn�n,��f��1��t�섍�b�-�0u6�t}}3��z.�m�dW��r�Is���\tcyh+o�Z���J� \�۲����l��e˙u�#��ۛ��t�]Nr�U��9$�s*އ/�c��ƹ�xn�0�Z��R�C�^��9����{0l�iF�۩:p���V����k�Qhs��P��p�+�SJ=�mt�6�B��2o
])�������R��ݳ��I�*Z��v�쮛�����&� �=��rDV+ܲE��J}�m��&p_8ō�lhUԷtJ�����
��$�v<�w-��k6)^�	n�}M�q�T"�KN�ыS	�N��IG��Z��@ml�ͷ��^���}L�W�4�fet�����Х�T�*�Rld�}x��R��f��Z�וpp�q7y.�t�+�/6�R�t��6)�%�GV��Trm�sb��f,�H�c�5�ڗ������Sҽٝ(�	.�:���&$^�ۇF��a����ٽ�G�o7�ͅ6c����ž�3aK)!aT)�o8�kw"�r[�]�b'�/��U�m���*g�A�jahR�y��1*K
�Y5��g���]�u�ZT5�Q���n����c���"F�QК�M��U�Gم�m� m�6e{���`l���Y�-T�w��`f�JI��Щ
��נjsj��L�G��&Ӛ�p�&L��K�8�b�}�f�r��{�Ձ�_7LXUj��/i^�I��I^�'9\q�d�7����'t�I�i�b�@�ԥ"#���I�,��6S�'����G�սGZ2��:]���М6�Q��L��Z�-��2�5���f�� TU�!�ʹ��]$�;��}w	�rƘ��]])gpկ^J@�/	Û:h�2=�e����CL�P	�}}ٌݡ��̙`!�2�0>/:�[&^Q���1�������tDT���̋x��9 )�U(Η��8EY��\�Z���:�9���}F��)28!cks��{[զ���(VG��8!k�O��i���S.�N��f7Γ̈c�b�'f\e��X�q6t��������h9נ�r�[�l�sn)9�fWR��C�RjY)�fQ����ή���C��ɑ�kFw��ź;���mr r�Q)�� +�.V-�!ȑg"�ѫc��X{]L{Kg�4�q\��٢P�W���\#iŸ�"�V�Flp)$i�$�I$�I$�H�I% +A"�v�QEL�I)oH(1��d��B��#r��brYD���f�w&�fu��rΩ;��c��ڻH�C�kd鶡�-e�ڶ��턝�Z#�:�R��K`ܺ�"��b�-�}��YV�k���bGf�w3�i���i�k��W�W�]{�t��
"=�Ɣ��io3�o��yF����jB⛛,��ы7�_Nl9�6����r9O���XԱd<�2�'[���8`�{k֪��5�Ȕnp�����*9��\������_s�ر�,kx8)gZ=r�Ś�F�*=��W�VAaY�lJ�|	���@�&�;ў�1��+�5�r�-�N=S��:�O@�U���-(��꒒?��w��?��/�?*{Yo�}M��D/�)�7ՊH��~Z�'Z6j�UV���$ A��T�ߞ�������kا�{I�>�y������Z�1d�X����Kv�'7�r��4��6e@\3~
VD�W��m�j���s�~�h�]}�r�*�Ս����2t�y��BKLa�:���t��C*��
ɖ9��!�Ek����wga�b�n6u_Wg1, j:���o.����mwe�7��2UK��D�MtsL���Y��a�x�Թ��U�7:��.��ԩH^4�}57ۣ^�������ufX�ˀB�ֈ��ȁDK#s���JÙ��[�ʷ�V�÷,=�߀�a9˂i����l�6�����]��w�.*�՘�?�Z�SGis`�ҳ����R��i���{����
���.�%;3/>v�mk�WR0HZ�{�_)Q�x�ܩ|�#p�9����,c��I�,���Ż+"����]kF8�?����a��b�K��nAC��Q�(mb�et�R����#!޽��B�:���B=q^,�l�$����t��@˚@��L�2�tl�D;���
q����o*�gu�̕���Vv����8�قq�mjV��ma�����+��7�q_�#�>k�W��H~]�n��`lfag�-����:�o]ƕqj[�����,<��ŧ��g������F�e`��!U�Pj��Y�1��S=i9[�&3;f�P�<�s��f�M�ݾ3M�a�;aZwt�M�=�Pɔ�{6��0��)�Xa�L��jܮ�HS�;p��yv�%�a���7@囊�&�Er�k�+���"�f�f����ז�)���b�!�]��H&��*l�!�p�b�/˾4F5OppΆ4&��-E3m��.�kv㋶��k4<�r�\���RCi�n���ZCX7%����;���]�Y�^�p9�cn䙙,^� _��7��ը�1]H�4M�b����]�{�YԻo�byDRƆ�^�򞧩<�}Jb�6�'�	`�YGPޫ�b}WS�슍e�z�t�aX/����s0�Pç6A�2��ٽ�c�o�؜*hG��n�f��Z�|�.b���qz��v�ӻ���c��W�ഭ1���k�9w;��N���3
�*u�筶���V�3��c������w-YI����|�d��HK��6����/��XF(�d}���H��A�j�.V�w�-�1�wOs6ݩ�wtʊ�i�<w^�R��o�ҙ�¶��6ẹ\�T��vSU��^DPV�V0ֲh�x9�sJ�1r�+Tq�Uu։��y3Vr�]����ht*gh+��ջ�,
$��Y�t1Խ����`�c&�L��؁��,�.�GU�Sm�(�3UP��2XD�&+�n��u�{k]�%�t���p@���ͮ�U���"}�V%Qv�p�@��֓����WW��l�wJriV�á��N�r�`C�.�>Ud���C*l�Y�رy%��䋇h��*>�����S����kr�Ⰱ	#����		1ަlJ��F�Y	ݺ�%��d�`�}�LܫŰ�n�=uC���5�Z��wi�j���R��Uy(G�f�t-��bnyB�\C�ݼ���@�W�06k��v��)���k�<��%�4���ݹY{��!�h��<�c�v.U��Bz��Y�6�'�a޻�i�,f�:�b����f��e>�G.�⚰\�wAb��׀k�|�2y�7Q��6f^��kQ5J��|��!�2�Wk
��M�<��y�aՂԮ�"���GZ�^LV2�)n���\5�u��Q:��#�_gh�#+]q��t��CU�+�3!:=6wm������g��Ιx�����*I֙�0�\#R:U����w&�NX��F���-ٽI7!֣���3ev�4��ۚ.���Q�}l� XK��Tثo�������(���MDeW"�WJ��k-�8��-����X{o+vAV��U�� �4�ǹ9&�-��/FulAj+r��^�MUΫ�8�D����@A�)�v\�/�����ٴ���� ��̪�pM/�Kp!�5�{��j<��@"
�ݧ�����|vi�o��Zx.��ݻ�Vo�>�ӐX�M�q �5)�2a�u�Y��閎�ʻW[�S����v��alٯ3Xק�o��9Ҳ�y@�tɊԧ�-��膔*����Aa�&�N��jtj�b�޵�ڢ2&ٽ����i��P�͗J%�U�%���r����V9�Q�[:���jQ�+�,B��3�i�jgj!X��p�Y5��A�ʃe�t|�jub���G;�Ք#kA �ث%��t�mΜIl�R5�,W��4�3\R=�"�ڭ��t���[��䚏�,5w�9��:���m*w�8fБٛ5��\wn��ݪ��7Vl\K�������j)�q�����}�/�m��T���H�WQr����ܠkӚlu"�iδ��6�4����4��֥]��C�\Sھ.��f"�(��n����)��d�z
`M�Wn�h P�wm����V�����<yT�/�89f��ev��7T��E�� 6m��ϣ��|d떛lɽ}�4��Y����L1|6WCy����1Z�x\ʷ�:A���á�ve�>��ȳ>6M-�9^&k����[0'k�ѝ����Ѝ��X�a� �����Ͷk4����l�鏰���-�v;�^s���ƂeJ��q�Q:69�{�ݼ�T%�-gT�ʂ<t����^���j�ᡝi0�J���Y��Ν������fEc�0�GVqJ���H��b�v���W�F����vw1�q�/��7un�F�_L��n�3���SM�Kd�����,"�=��|�p��K��ͻ�T�S�I���@�����l�N���ƨ���,�N��t��_L`���ŗC#��E:��Z�L�e=��������I�K��ܲ3r�4]��g�T�\�*�l(3�_R�ʽ*�*��v���g֍hS���i�ٜ��C�[���Ѯ7#�tr���淧3����1>��Wt��#���U\��q2.]x�wB[��t*�Ō�|a�79AJ�ِ�ٮ���g�!��p�L��� d�}c:-���ؙ��z�MtF1�mZ�L�w�g*��+Wl��s\�ƪ1R�D�놼�%�u	dS�|%�4���-*� emf���G�_bG�����3�z~c�A�_1;L���U��zi�߷�A#5#�����]�9@��+���j���ط{m&�Rdq�%�����!Z���0������OwI1zm����U�v$Uf��Z�}wef�r��y�>}osyYj�E:���q���F�Ѧ#��|&�6���
�eUf�c�e�4�+�u��M����{yk�v�\�'WV#®K˴�yF����QT�i����oTu̩�۽����I���ދ a��>|.��)�s��r�u��&?�/k|�Z�Jʶ���C���8U�]p�Ȏm,��@.5�Zdv�7���ܚ���]�t݁ٲ�Z֌�uܱ�����

3�)�᪸��[|�ᳱ�9�c�F�H�p���\1C:"�g1��Wg\@��j�d�B��R�����WxW.�m��j;��ēu�������+@&*(pW�ϻ��Q��0��d]�[�e
�\�2�ww9㰟GX'2�kp\͘��}�/�B��E���囼|J9i�����
�q4mȦ��^с��y��S�����b8a4��[x�kzܘ̩���]��q�n�R�$33Sq,����� ]��Wl�>-�JWU�sr�J�;!
��]�U&I�0Y��B�(H�g^ֻ֓]G���੻��0w$@2�+�t�z��7�y����|�����O�~�� � ��끠�@F��@���0�g��/���h$���S(mw �˩�5����`��<����O0о��#(5C�n_r|���3�r��y��tNf���c�g/Z�p��$�'n�K�*�c��
9bQ�quL�1Ր��-�0��ևX�=Y@ Wr{;Aq��������CL�����%l���gNb���Mi�K��٢���7f��atnl��6���wR�Mz��>W��s�F�qE�}��*�s,�yb"�c�-t�zi	��(�����#���r���}�l���Q��p���@����7���I�s�L��'���n����`�;yPZ^�����`��ɶ���C!�]<M�t
���WF��e[5ꑎ}|L)�p3#q)*eҢ�C�3Wv��	�v����º�WJƆ�%��O݄BH�1��(,��(�Ũ�AP�)s3Vc(��G�	QA@PY��L1QAP�*��R��t�� �"���T-),�@��:ABt��Db ,�"�"2*�"��"�J���Ő1%IU� �
F�VL���±b�f0b�֠�
E�$QQ�1�T�=�Gh�a�����A�w=�!'�TW��Z�N֧�SF]���o�Eʯ��I�.?�}_�U�
ܒ
�#ۂc������1!�&��*��-%��oF[r��d��i�X3tR܄z\V��̮��ź���'��,�+!�!�t�dKJDw�q{.�T�m�k���m�3#�ַ�!�Ng��u]�k@qK�������>��ZW>v�Ͻ��<t��3je�Yix�K�&�/uX��c�w�y����򃶯���CQ��k������bى�����b/;���������c;I��:T������κ�\{�Y���b{���-����N����B�ag.c���M��K�iR�Xz2�K��#K);^P����}��Uk�cI\�S|o��[�e�|97S3��������B���Ѵ�m_Y��U7U;-���=fˠb~26'ms[�z���-b�pv�h2u��+ ��NՐ�8���=Y}����k+8�]���L Ȋ�Q.��5{��
2zN)��^�9SΌ�ec�ؖ�fV:�y��cҪn;�rD@ܤͩ݌tb��n��
&#<7ׂ��]n���>�o3KH��K�D�����ގW����ޖ���y�`P��� m�Ym����9Ԋ��^\���#@�c�;�^�v�B��%%��"eí�0�:�j�}:�Πxbw���[�� �O�ǲ�}c��X��)���%�ƭՅ�m���׵�W�((�<J�j��NPY��\b��gp���jOw�e�Rj݋�׽y �F{_H����ͣ�3���]>���Û���;�}m������;��_.5q3<�>��$��)��Mv�8VvBl�c&8��<�W/}����=�Kz���B��<�^ɼ�}a�̫~e�7�Ɖ�@�z�;AM�3D������d�)s��5����-Z1����2���.���:�ա�?R�P�Ms����{J��v%&�ot��:k��^Q���Ƿ�%pf��D�V�MTd#N&y�����]o�OF�l�c�3sO��yͽ�t�cP�8��ѤE��,G�g�r)��lk~,���宷X-�Ca�ͿH��J����m9:ҧ�b���P1᣹k����Wn�tQ/�-
*f�|�Uv��j�@][uWm����r��M���X�ͣ"��� g�h-�c�b���|�C�Z5g:i�_*�p)vc�%o5PF�k�}�~90U�Ռ���N��.0�ׂ����̿WD�M/\��s+>*�_b��I��83�X�'Ƕ��9�{3�A�^�1�W���"�j3X�s�<��[�{	�N�cR1�6���a�V�J�~��� 	!{]��y��0��}�4מ |�Y������#���}ކ����=��Ioa�x�i��_��m�@�#��Y����x�p��W�~(����6)_�yWR����͘�p���ˁ���$���!���S���u�b�Ne8m�ې������h<������ʸgI��\�Y<�(8�8:�8w���UyV����ڊ�/��P�o��`s��Z;س�eg��o;+Z|�j��j�I��̬E̅����1�F&�;��2;��ƪ�m=3�t�Gc�D��4awv�V��w1)��G��Z�.kZ�M9��X}^�I�4�����8�g�//�g�u��WQ�9��-qU0�F��bk�oc��Γ��C��3<�^-}�h�dp�G.��^��#N�(�ȓ=ؼ&� �f\�,�S���7�\��,!�F}������L=5wkUԍ��/|^��6�;�n;�mm��f�>�|OY)���M��-�׊��f*]��ܩ��\���^�%�{Ql+θ�^����E���,烻���VC0pku/+��x%�����~�x�,�9���7I!xܼ�xZ?<�ռS�����F�VG��1>�ӜV��nH9�-��B1ʀ(̑��&��g��TW^�W���;�,�d_�N���<�y���N�,"��zY6{V}��~��s��8��A���m���ٽ�����W����`�C7^�3+��e�;�!E�v�L��`GA4�NB�#&o�g�,��K3wހ�t�Cإ�n"�^Nog^C�5c�W���SD�N���hn[���\�D�ˬ�`�Ef�G�+�8�~��i>���{-S[��!Ш����?2Z�D���=�Ѭ�;0��n#f�v�1S~�Œd̠�����}^���yf����&�pN����PX�'>�Ṗ-��'	:�,@j�n�Ӗk���՝�Nm�`f�6�yYW�6y�t��i�&j��-��l�v�Ἰ|voi>��H��qLϮg�}Bf�]�Y�C�s�Ϡ�ߣ�M�k�=�Y6�i��}�i�''��)imǉ���c��4��QyN�o����D��x�t��6 Z�u+�i��n�Q�jFzD�V�{P7��v�Hm�b� �"��F�9uh�$�Z�I��S��>�h^x� l��wjN��ܕA�춛��vYK"}T��v�=6V�Z#xz���K�8����[6:��y�ؚ�Foi滧�*5ՌH��2v��ɗ7��C�PI���o���E����؃�%�=�}��/���c�c��V�@��Ϧ��.���<��]e��Ul-D�����X�Z���,�p�ANɋב��F�r���ЌS�|�2 �)kkz*�]��v��J��(�Ķ�Τ|tf��	���˻�鼡m��< T��|�Yvz��������X�jz�+�[���6.T�h���t��T��4�g�'�R�`�ĕ�(�^�b6e�Yc�K�`!�Z�^�4q�m�"њ����_*ł�:w)���(�f�� �r�e��4Zw��u�54/d=n��^B�c�e��!݆l��cFs[.g�V!��bL�2�!aW���]�Jd��'�������e�;O��T��JM��-T"�$��RUU���/Ms�$���B�>j��e''+G{�u�z8��g
˪��fF&\qbp�m�������Ѓ��YT���� ���t�[�_F-��q��Y����t��ɢ�Y��^�u5
G.�n��j,�p�b�4�յ�{s6���z�\�����*����ֿv�n��#�D���f���X+���ٽ���)���%zߴ��'j����;G\�j�1	߯q2l٪��x�[����]�%�-gw��3c���/e�]�������;�n=���b�m+8M�QaVx�J[#��Ԗ��_;��!��c#��#��9�ҥs=6�FTv��Z�WnfAv�Uug��s-��vWJ�
Ѵ@	�<��!�}Z��*��7N����1��7�ltEJ�1:�_FVw �X]� �Z��B�(��:v0�7ƌjڂ�>�Y�mbX+N��/W:jM�fr�����x�1B��
Y˽)�de��̝v���9V�Fe�8�X���]d����(��	fn�q(�7w�;N�崆�k�ӡw1]]�;$���B��؋T�6ݍ��R���fYa���\��t�N��f��ы��ְ�ԳT����/I��/'!�����I3�	v��/��y{��T���?}�	���u�)?������M���7���]�+�,�\�h�m��{�+#Wh�%@,�GnI�Nm��Ot٣D�����[�SC��ELW. �R�f���V,��Z���Pg7Zs��·�N��Vt��:��؆Y��k#;y6#E�$�F��y�yi����Ȯ��̡r�TX_U��f�a�nx�����F��:Vۄ�v�L/�;1Ź�n��_d=��	�$s*�6pL�D3;��U�dvs	�c9q�<�2��{{�/���;ca�Y��k4�⻅#�T��
�S�fIe��]<X�;mɔ�&��wj��q݊8G�3[�rX7��Or�1IC9`,1�$y�r0�e�̍Ĝ�3�4VX������YF�B�1��@t�K�t���L|>��Θ%Bi�J�Q՘�	�$XT��"��*LaPI�J!X"#!U�%Ak�ȑHbVAdP4ʁ�X�Q�P]2��֒�
 �E)%�� ���"�ńY�Af0�H�U�)��E�����0�/�}aM_�3���r�u%'*��614s2�c�Z{^f�MN��6ё���'u��9-�����t�׽+g3y��Y�$�@d�|�/��[���������H�Ea��_��~�moL���ǿ��J��Q^�B�[u�<��Ջ����>f��d�lGF�G1#-�mnu������ۓ��p����ewd"�r�r�*�y���XG��
��_v��q������h׌!�C���N���o�m �j�Z��F&c���pyxZ�4�7!�,����PV��c��t��'�o*�㾺����v$��G[oB5s�x���e@��]����Ɛ�W�����صJ��ڄLI�eE���)��-�^��#��J��\6��f��\'S������A-�^��/�=}�Y*7eE;I��o�'�w���ثް�K]P�KD��N-Eb�z#Y�3�yg-�7����֡ͪ��P4�Yuo*�³������*dJ�cӦ�`���|���p�>��#���x��ǜ�!@�����P�\��i�O�c�;�OU�q���r�YI3'�|ՊN�O�{�?{�e��.!ם^H���&����I�Wx�e�h�I���|��Y��ƞwF������[<2OZ}Gڍ�o��+�Ho�ԃgZO�mon:4���������6�Sf�F�0��G�	��?�_Tt�7�n���4���ؤ��hC�O�/�ÿ4"00�~΃e�̿���Ǌ��6��o�q���ے��d�\?������g����G|�q>��q�g�B���g�P��R�<כd�~�[^�2�9���R���l����xs�EU�稓�o[� ���d�)f��Y�L06�^���.�L�F�.Ҩs�#��5���W��S�s�>���W��G}֞y���}�P�'VI4������9��!�& �t��ݲO�u�Hv里���C�'�뛾������CFR/A��ݼ̡�;��:��f7vx˶�k��g�>�)X���h6�5ٶU�'��)JR�$p��A2o ���UT��q��Hi�?��B��v��xwv�>d�t!�3�`M�VC����2Ї���Ld�<����:�o}���P��hC��@�j��M�x����I��i�MwI� ì��<d;a�I���s���ws����IXz�RCz��C�C�O>a�݁��8�;B��'�����I�@�{d=BuΎs�}���7'���|�lB3�,I���\�I��L�6�q�!>@�&�J�z�ޱ��O~���sଓ�;���$���m�퀰�@�;݂�.P�%zd8�Y'v�>Z|���q��s:���}��C��6�̤�=�I�� ��m��kv�a�	�uCԕ�!���a枹�w�V�=�~s8l�IP�;�P���4r�|ɇ)��li$���Rm��N%Bz��4���9���z޻��9��>d8ux�+*a5�>d=`|��	ٺAI�'��@��}�d�wa<I��s��}9���]����C�C��q	�O�LBu� qq�T�q�8�I�Ch���E}�=d����Z�==�<�|�M���æI�>���3�'�<d+!�}RN��r��6�P�f$��}C�Q��?}���ƣ����l��ʗw����Ȩ��:��o"���p��fbu1�?r	ը�'�K����XV�3�J��@ �I�elL�O:k1�?�}�Q������ͤ���N�M��6����H���!�'f�1 ~2t�̇�����Xc$�;O�C�s]{�����@�i:`i��OwI:`z���Iē�ͲM2�!wC���7���HN��Foݬ4������菦=��A��l&������d�I�~w���42x��t����C��hd��$:מ�������I�N0�� m�����M���ĝ>2zɶI�oܒ�l�	� X��$�'�}���s�o��|�T8�X�'z�h��x��rϙ'�m��]o |���O���g9��$4�Py���k��oߠ(V��%d��ơ� svC�OP��&�i8�z��|����P2gV2Nٿ^��w������^3�t�v�I'l
ZI�M���b ����V��<d5� z�秴�l���	�s~q�ӧ������M2C�0���hm ���m��P���!�:5a�'���|�Щ��zu���r�f��u�7�>6���v�ۈd�>d�!��m��xy@�N�-��'��E�V�i��z��Y����o�w�����?0�!��a>@ז$�2C�J����l�x���)'l�+	�'l��{ǖ�������x{��j�c�Pfe�X:ڭ�XQ���M����d��t��:#�EB�Ħ�I��aB3�]a�ۂ���)�S�� N��{�{��x�m�wa���d;Ha�vOY'z1m�������M�`H�`(C�P>���z5�o�>���d��BfُI'�t��!�W�IR��$:g�R{`��I���ԝr�B�^gG�w�{/o����!����OP3t�ĝ=�!=d;�$9`i�d:~`z�*o�|�8�����9����g�}���p���}�$Y.��=d�d���t�1�:O�M���2j�i0�O�;��}��}���ߧ���a���P�a�d��d�ɴ���i��hC��!�Lā��N��!��G���s���=���4����d3������M�w�Hz�OI'�L�d�%N�!ϸm��~������o��C��;C�'�OmM�b@���a�������M<�t�<@73��������mֵ���N��u@�I��Cԁ����3T'i=C���O�=a5��{�<��3�1잂���=���)�������q$�hh|��q$��F�<a�&��P��>d�a�}�1�b�s��ky_X?%������}�<d4���I�큅���Ĭ!ی<`,2�z��Y�l�(��=�;ǸA����R�>�����4mX'�۔3Y��h`٘Y��әR��6���rv��P&��B���|��d�����K�&�s��}�}�G:�=�|=I�ē�(����|�<M��!�&��M����'i<OY*Դ=H��x��]^���>�N�w���a�����z����XN��M{a� γ$6�=Ch~XOK$�'��!�:9�n���|�|�|�4�P��x�'V�a�_���ɴ�	�d�@��d6��6�Y/����㿷���k���7�B�;�Y'��P���C���;B�Cg����)<f�Me	�=d�z�o�$/<�_o��w�y��I<`,��� T�,'l��̐�q%t��� �y@��x%ar��!�4n���.�7�y��^o�r��_��<@5�'��bk(C��1�$�2�4�|�>d�%d6��Ƶ�y���w�(i��� ��iY't�$9����I<d�;�!���~H�X'�>�n�y�}u�>�rS�CI��>`)���߾ם��溹�\�������v���N܈ײzF���6����ӭ��z���xj|��3�J�(�*r�Y9��茥�y؀UȗJ��׽�2��oe��c;��+��G�^�����vz�w(p�<9qû#�6�Hԉ�������Q5>�T&n~�F�Z�>���ˆݛ�n^)0 �(�3�V�<8�xo��_g,��A����؊b���淂�$�>+���أ��hέ��ы١�-�z�7�F@H�XϐʲNB�ϪC��#�E��8д��/!:��n.dLfP�(����а������(ㇵ�9��$�Y��
����d�Kt_O˸|���G�hmR��}�Qz�7^o:�^��� #�� \���my�l�O��������Й��=؇W4w�|jV�x������םu�����n�9��ɘ��u|�^����,�<D�,t!9�}_W�_Q��R}�����~�I��Q��v�S�}�"k�<iŮ��A��8ՓX�d��HR���W��y�y�G��^?a�*���I���[;=T���7�{��'�\�:���!j�<Pܝ��{6���\zrku�&{�J�8��{=�鱍���E��L���t�e_�q��`m�yE^	���W��]'���
�{��.<&:��[��($KޗU���k*���2]�f���h���Պ��!��7:z.����yV��ѵ��ꪉ��cMUʼ�9U���Z�g��r��᫫����Vx�ƻYd��4rAJ�:�ѐ�R^�qF�򾪪��ms-���S;qz����ڲ�Cf-�'[:�|���Kֵ���מ�S8���y������]*(tLoeO0����6��6w^ß\����:H�b����`-�G��Y��M���yS����[��m��U��B"�˴v!�sDk�I֓�qb5����0ͨ�8����[�tO.{P��K.;)����v��"烌��g�5}]�J��7�k�*^p������T����eƐ�b����f�e��~U���c�b1㒢�f��bo�l����՛XA		�vb��he�u����[�ZN��)�L����\(s��ɔ����V�R|���uӼ��^6k�>�pf�֭�F��]�ekA􇶊�N[ێ�gM�L���"V������pc���.m#8��5=O\�gv��V�&�;���oNo�\w�rΌ6�Vw;��l�ֻU�KtF2�_:ԟlZ���V6��	%Ck�J�+'	�f�;�ݖ��h��`c�W�4)}��밡�ϥ8�D��1b+Y��OyU�4���t�ǥ���J�Y!���b�R�*���O��ݏ^)u�s-�2���ᕺ�\�����5u�4�]��Ga��z�L���Q�{�dη��Gu�l�k�V0�#�uu_q]���"�|�ۻ�c	��1]9Wr��[N��/�6,�통Z��Ζ�ٵ}�v_����V���=����m��/M�QCl����<�9H�
+�/M�gV�}�z"�s����7yz5K"�~G��3c�*u�9��U:}����3�In�M��rK̩M�[]�p�˽�4b{�����0¨$���;�)��0��O�g:=����N��dG���C��qfm[f��ӗ��m�Պ�
�x93���6���s��;/��V��5-�W�F��\�T��kiV	��W���Sي���G�c�2�]K9j�̤�)U���*�5�%��@�i9gWt�v��2�la˽h[��W;�x��i{�o9�(�͔麽d�9��vm���D����b���"L�i�ۉ����*��ga۠�����y��Lƫ���]V��������ɿ���a���P�#�V�Hi��2�i	�IP��f$�hCB���J��2k)42AdQJ��Zæ���V�dX�Y4��T��D�m�Lb!�N����!��P�
�����%`b-e@�ɤ�B.1J���JɊ���*U@,:ez�E�jV�)Ӊ�醐1#���Y�#l�5NR�]����&59U���h��!@�,v��p5�n�\���'������V��+�?�c�߫���9���_�f��������r�YT�����{^g~j}3Ju�'��~K9�E֚���MGMI���D�s�'�z��+`"j���G[dS��Ma�T=�=��rL���)���|����qDy�s��ncM�e6�+��H��S0r�x�Y㈤ڠ�y6�L$������hZ炳��jxɉty��<_ ��&��5����zJRM�i�Ɋ�h�#6�{�m>j��_��o�j������tk��
����3q��N�D�{��p����v]f�Q�Vs��;4Xj�s�9��m����]�n������(�%W��t�GnW��wN��R��4�u:���t��z�9�w�ڈ�Z��Ԍ>ܕ]�|��J4�)xo����ʓX��V��(��ⲫ5U�uq���֕�8 n�3z�Lѫb���Y�F�<�c���"	z�N����ʗ�8o���[X��܋�Z��q�[*Ο(���7٥T:1U����l��4:hG�}v��L  ��Eߒ���׫��=0�x'�g����<�닐��_L���Վ������\�W��T}II�b֊7�T�X;[r���q�^�����÷G�ߙ��1/��z"��!)`�Z��7�n"w1�-#5�%Ӯ�E#��UUU_T��Y�Wt�����h9�y,u�UWK��-��-�Ӿf8Y��~�2v�%�d��rhm*����Z�¾9��F�����D1]�;D�W�;K�����R�	�2W�r˶#�����zٵ�jzw);B����oAs\R��%��5��*�>T)v��p���[{�V�RN*W�N��Ow�Ÿ�doo�[X�-n�ݳQ8��(l�vr쁹[e���!��v5O�ݓ���e��A���'�w�xf��McxҘ�!vU� 5�:�+��+.��@~�6��&����ڎ*r&��Cie�%�Ą�s-^�Rᚖ9F��ϫꪯ��bG�'��4��h�]{�bqco��n�8������t��#�lp�j��Yc�e˗�ݷ��Fq�2�)�D��g{�p�0�̨�����F�*����x�.5z��@�v���Z<�z�3��o�5��Cg�Zh�`�Ea�<�.I="�b/]��7I�TP�����M�c�m�Щ�Ea��R��7��1���c<��ɢ%�u��-N�b�&��������4�;Y�U�5:���<��Ѻ���^�����X��EӃ"����/H�Q�D�^\��K��n����:�=ޓ�ʼa�Y$�'��k�G74���Z[�*裼����z=���Kb~�;~���x;"�T�Fi�|#d1Y��r��[��U����>��f�T�]���^!�:u���ޯqw(`����d����:��Ms���%FM���'.m���ި��<��k�w�__&��U�����y��j�qbƩ4Q�C�"j.W��Uaz�'_b�`(�g����1a�S�i���.�ހ��y����/sۈ!�`�Ͳ�{Y\�T=�k��Y�^�]�Z$����݄u���aj��ر;��V�#94Ya:��V�I�9�IkS���b�u��m��S��n��v$gB$����_q���{����p�Ԏ�i���do'��^��1<��, �aU�[����+4�Z�Í9	C���J�����堦�x�$э���T���=N��������������*id&��}�{�(q�s�+t�Z�-�bm�c:|R��z�y��{�S��x�|��]�����yS��B���<�hd��k�Z7D[�7݅Rkͫ��M���C�^�囇|&��sv��U}�����z�Y��ͳ�A��Ubb �}BFh�P3�#�L|r�ۦ{gZ�|���+,�e�}.Ʊ]sc:
�.�LG]14�J$��1�W���:�]�E}��{�
��}Zj;8߾/,�4"��u�|)�WS&�Ԋ9��ϭ��/����(��.;Zk[����mvah��~��u�^��v.�c��r+�(�.� 2ھ�έZ��Jf(m�&��q��2	��ׅsޖ��3{+5��N�{�{|� �
���T�ʲ�ZMy,��Y��hlt7����Y�|�iXD�<a����Ji��bI����hR��b�x��'
���-z�f�'�U��fp9��X7Ƿ2�����/.���m��;wU�j�Y��]�7���T���S��y��վnv�ڛ��+��5�ePɹ
���$������؎.LV^`���}��ޙ�������>;�6�C�#*�%:s�hގ��N�}�����vo�r�D�lM+ogy����r����7T��Xɏ�O��|q�/�O[	X ��3�g�~	'�p=�ga:D>Gэ�響�b�r�^�Y.4����L��Om������Q��z�jy�-s1�$��$W%���	qw	�6��3��B
��1��bCx��2���n���Pf(��?5�D���5W���k<ݥ�3�ڍ�J���v?���i�Muko���TP��#��*�ή:ՙW
��}�wz�$i�F�I�˟�磌��H�=Q�gY�]��]�'�WU�����m��X����~�Ts
vө��{����[�}�I�޲<x������ ��U�'�;��=��5���]��b��'�J���Z{k2+� ��)R�i�������s2���E3De��n+CC�����ux�ބ�.S�v�����j��8�����	��L��=��5[~56�}���0EE{UDf�<t�}QNX��{�2>MpX,[�s����D_!n�j�⌽j���d�B���L�h�w,�u��E����c���@@pn�ُ$	�!{��x�<9$�]��*�\q�WHh1ʜ#e����憎q9 չ����͏���uf$7���9����#�F��wg�l�Bj�o��#M$!���B�=v���>�k�g�u[�tn����-���
:l�8=�ӷ����x���9�Ə����5w۬RXkQ�ߴ���r��D����1��!�@F����<�%�5"z��nJ���w/q���:���#���v��1�D}�	>�پ�(��<��b'��?�@�ڇ��^�O*��߷oH��_��͍-pbȣ���4��p�ϯ-���^�I{y>��q&z`�'�g�kbj5�n9g�.W���U����X�/���Di(c'KC5q��i`�}u �����ݐ�^e���S�=M��O�<V:�s<�Z�Ed[f��h���Y�X^�'��6U�n��ٽ2�u�F�<),:c�;Vm�˪��V$���5����f�9����(8�{hV�DS*�z7Xܰ�/�B�$P
.�TC�Tf�ʎf���>�]�h�d�p�]��Wt@�ԾZ��T�F݇jҁvB5U��R�﷥Y�f���U���H��V���)���u�s���n[�����Y|�JH��q�+u��ce��w�EJ�P���0�5�5kaU>�x�V�wp�{��Ky����
����aY�^�.�J.�^ǅE�V�{R�^�5Pg98�mu��N�q蝈L�eQ�Z���=����{|g2tX��']*w1�8e�C��u��ݚ;��:9.a��7w��[FQ�1}k���@�2S6��n��^���÷mP�w�+��s����߈�S��[6U��i�[-�rV�}-ܼ#{O�,޴�3+`{����A�tn�#�dM�I�s5f�z=s�7�������������\c^X��7u(��X9E�N����U�$gK˼l�ލEJ���OMF����d�Q�Ff>k��k�R,�����U����vno�	z�D	�5y&��EP� �x Hw�}ݩ�T�XL�é΍
E2���9��V-��T�`% �q�NN�Ttg[��I��!)�#WK:\�z{&��0��Z�%JFm�\��{3�%����/,	�O�	*��11��G9w�M�O,��R ���`�k����J��s�j�o�Xsj4�n�+�jU���}�f��s��{�	��s��	[��~� ��|��55�A@Ӊ"�ń�YP��"���+"�IYt��4ш��ĊVV��� �.uE+Q"0��TP�ҥQ�F�G2�'Y���E�TYRT��++Pֵ.P�Y�R�$����*+1̢�I���`)Rc/T�&��m���Ƞ�\�(T1E�R�!U��AQP�Re�Vc+YXJ�=fH`����"�$��&%j-E��J�Vc�����xj����m&����+<m\�B��na?wmՑ�׬6�jj���軑�>��{�Wel�x�BE��a�0��"~㜑&)x�:��'�Zൌ��t��CN҇�B`Ǡ��7(v�|jf�l�p6B�)a����$��f�Z��C^6g��Yc��ٞ��-{P�삌���⵬-���31/v4�6�E��^�6��߈'��+�F�D�#�61�/�[�ۄp��B���L�b�ʫ%���L��Q8�U���{WY��1��3v��w�V��";cU��c*J�h���Q�H�<���`{W�Y��2�g1�[�a̝�rU�7P�}���6H6}0�kҦH��U���c�8�;1����
��ަ4�19j�k�N�hW/�x��Ox���Q��w]�B쨚J����zm��n�4�+��ڙӋ϶w7��|mf�*̊�ZT��(J��`ٲ�:;���M)$�UU�#��欿�v3�ŔGO><w���ᣩ��*��YU���)M��S��֬�k�`���G�4�_f�hb��k��8;�e{}pUs�~������.��N �:E�$��lԙ3�@977"�"jIi�/ˈx�����wW��i�9i�F0��z�0Rc�ž0�5��1E4V�dNI��"t)����9�� "yi���P��y1,/�=۞��Md�������ll[X��zCHn�d.�F�5��2������Vz�U=e��BͿl�������*2�)���~�'m��y�ǧH
���Y��5�m<�)l�p:�ٴ��x�Oօ\��ź��"r�k�G�^շf��S�LFɣ.8̓'.��/����r�N�~$�C������s�j{!��#Q��\uR�ٮ��e��qj�v�.���ޏye����*~�!S��
��$������t�����-sK	d�W,��IR��>x,*� N�B5�*�־�]��� ˌ��f�����Bȣz�V��Y������|}H���N�� z��XYq����\�R/�S˽���zi�i�I����|�����G	��wL���>���!��T�t}B:�Ӟ�9�
Nk��d�6gf� ���OU1<�l���4�x��bΝS����#"E</^��*-4G�Z)�0U��^oni���e�D���ϱ�ӆ]�4��W�Orقs��٤������kY#H%�y��N��9��].��laR�g�afF\6o������4�R)X�O][���-���_D3J�t�c�esu��]JV�����^��r�h��}U�T`(�d�_�L�����%�G�㼑шs%5y_Y�+���C=�Ze6<h��q���J��O�O}a�w���.�R�EJa5�y��pjb�
�������a�X��ޤr����q0��fʘ�鞋����#7�$�b2T�'�U�ٮ���ON!�d��{\-�����v��_����ib�!#�X�$e�w^��'Ԭ���9H+BR����ޜ3цt��~�or��t�yP'X�SC��=y�f���b�IaL����ܼ;�A�'�CXCܪ ���)�p$��ة�p��:��=�;����冒|�ج�OKh����d^p���*'���auc�u�v����gWʉ���e>�kR���mf��FxkosK���\��j�2�I��&na��Pn~����z��z�R�kHkX�������a�;p�M�f����ON�ɧ"�2L�>#	ЅF�>li~�4��nU��M���y؉=J}2gT=0q�I��B�'

Qݼ��ECn��uu��m]����I�Nx���O{{�a�͑��n(ЪTC��|�yND�8���*{5]ww�"<9�4ט��Zf�v��s��6���zI�����@���0�^6G���0��~6F袯���z�s����A�%��M��q~��$D߄D���u:E�[)�9����'�|`��:t���_i��Ha���u��nG�����2��ǹ陬1K�X���3"����+��uO�����ۦf�*ȼ�wiF.��I��#�,ŭ�ۓ�0k��7%�����齋	)�B�H�ͼ��o��UWH�r0�����#�,�!��چg;�z��B�1�Í����3�:l�6���=���0��F�v)��WN���iδ"C�qY���O0�'V����>��z�Vg�b��c �qx��Li��&&	&M�C�o��w���X���tÅ���Ϗ���5Y$m�$h��6���&&׫G��&�����ϊ˳Or8'lh&�}}��P�-tA�\����˦���q��B�G��(t9�SvfL�y�.cl����.T���F��t��ݐ]W�x��~O\p�&a��J�]/zf�o�i��y��"˥Ac���L[vD�{q��B7��j����A�B:W|}�n��M��������\�m�r.Ժ������j�s���EYZk@�C�7�q�~���4@��w�kn��o��ηޝ����N$/��D}����J�{3��� Ej��1�͘o�X�Ǡ�GLTz��F���! 겹���2az��K�1F�O�a�t�'V�}�:5��$���`M~2���xkˍb���T���y����;�I�g�#�&c�Ųm�����,��3kuV���0H�ԏ!��6c�<x��Jl^�e�Q�B�e\xæ���E$*������z�^���d�q�g�r���dt߈�Lt�!B]ɓ/4�|�ei?`�|���s�><AU^۾��Y:��Q��a������Df��&X�7���#�>�Q�R��y�����i�Q�߅��h�+��h^����� m��c�p�m��x8�	�*#z"�
fl�ͽ�OFB���5��{��a%��تg�39 ��p�C(x���A!�by���{]��HG�iz���H���Y����Ŧ��S9������p3FX\|I�L=��A��Ն��!�6�7��^^^��A�ׅ���53 �����&zv�2Iv�>�m"}v�KB��)�s�ꙨwJo�"��/�a������f<��{W*A>�dd�����:I��N�e7�v�����q_�B�Z�L3�+��k�B��������Z�S�Y�B�k/گ�K�1��i���=ң=梔���˱@FTί�T4Q$o��5�l�s��	�G�)��৥��!�R�"0ľ����|eU��Xe�-�/2ߏ=O)�.2��
�<�{���ٽ�9�s�o���]F�ܜ\'N�;��M_G�܎�\���'��.�Ȣcq���)wFL�"�.p����7ҡ̓��m�u�2W�|I��r\�ͳ9��F H�D�Y�x����yY�0�p��4��A!t���_�G<��Yo���u��H�;ۓLI+5�${�:�����3p`og����̰ⶂ<A�=���D�+),7��h����8�L��3� �!�Q:{���fT��=������@wjg��{��|�<��N�B��c͝$��H��u���N�h������b3�\��J�N��<ī���g�C|��\v��A?1��BE{X�B���L�x/�.��{8�Jh���<��a�-��9^��E���d�$�[�������4�o��TI�D3)N���Xz���*W$�����5��er��ZS��t�Z\��қ��η[!����U(D���W_���^��t�l��Qw�r'e`s��N�*ySٺ��i�`z�j�7}�Q�}>�GP8y@q�����;&e�WI���J^�&zU�ߑs`NN '���91lC�S�Yc)ߦ+i�m�B�tk�]���J/K}��cfX�y���b�tg���U�4���'6��Z9�7"v�t촆>l�@{Wr�����}��{�ǆ/yA~b��ب�6Vw�G�Z�W�hFZ��L�y���+�Cc��CH�,Z�P ��d��N����(C�'�Ǐ�45��㼅��t�P�V��(��
:
T0[u���te�=hi�c5�>��Z\�+|W���Idv9i����+��c�~�La��y"Ї���	���;��ڨ��R�U����߫a�x)O�5�c3u�[�9
�S~�:������TŲ`b���Gc-^�E�U�wuj/fY�J�(�6��]ib����T$��pt\/k0� ��{�e6(��w��=kuMF^�ldv����`�u6'�$�; ��f�ZA�kyCu�[S��`��ah���Gs�Ѽ�v)`toچ3�ʸ����!�Vbh�y�Ć�a�w�c�f��|��&��pi��q����ζ��̣f�SU�܃.7��u�ґ=�O$J"����)�ar��#h$����B�&�x�
X��4vcMC�=�7wţt\sCb�{yəe,/�-���ؐ�s�&���zK
�8#�Y�:
qk��73^�*rF��x���U��ekڋ����g{�p���0Ouw3���l���n˛��#X�T���:�e�ų��H�["@Hu�xo�$n�fR�f ��g�u��ǋr���x�ZjKYOz���V������ڻ2�8��ۜ$���yehT�ے��E/����X�ϰ����f˵���?��^�ll����#a��>�7X�g`�+�� ��H��;�GoU��[����xxрס�"!��t���[���:ы���k[b[w��ݷ�1��`֯p�|�e��x��r��M����:��Le�,��e�Ӗ��"���<mۼ��+���oD�\�6R@*�C}ܡ���q���=0n�Wz�Ųr��H�w8<X��2�S|��1��@�REm7��Ad�J�UJ�m�9�kYRc*(��Ր�&�gl0@�m+n���8�Y����TQ���b[	�.Z��B��5Y�,��s.Z���U�1d�e�b��.9���+1�h��m���s&c��8�]`i�!U!oX��R[�QK��S2�YY�C9b�B�\�B��ڗ
ʘ�Tą�"�"T��i���P�m�Qco�Bl �	�OW��{���N�3���}��V�&�Б[S{	�6�lG"�ګ�jM?e�;��r��?˝�|��Ť&�˵9�F_U�ogQ��.a��<l���=WB����%�La��n^o��}�괇�>8Eb��0�㇢giVo^*��C��Vo���Ma��<A��m�J|���I�`�a�LN�|֗)�d��^�f�c�ڇgt�山mc$_����f�~�֎9�ő�!0&��UEG(��:��`����sݗ��t%�҂�_>c�O���SخZl{� $}x��5��w]�j���F�$����q�XtK�>��E�=پ�Ϣ�cH��*@��t OL������g���3R���0$Aں���o��A#�?�j�l�^A�·~����>D���Fc�������l�eC*2�|$:6tl�b�S#�ub�]WuP΋7:��Z}�XHѼy\� (�_���P���ha��Lx� Y�7�}�Y�%��&).�۽���>X|=2�)�gN�<0��3V�Ww�ѥ�G�n�%�,�0�ݣP9u4�)�oud���}���I��?2,� j�x���ֆ/�[g����ib?@|#�L�鏸l�:v}�u���;�Z�좚d����*%��֛Ն�_qQi�<lod��z�]li���$����鏿�㦱Ҙù�=�߾9�b��ɉ���#35���y�Y�A��{۝۾2��|��i�L���E�'�q�q�H�\=��37���))�0�ּe6<h��Lx�!	��Ф�s�p��Ϻd=Q�;졜m�U���Bą�v���u��usrr�r0�"��U����r<l�� {���U*1[�����L	3K�U,S�=�q=�z=�����1�{7�g� �qdB����L&�����XwJ��gz�6�fA����Zk�菓V����s���̚4m�ȉ����O����Ƴ��\�=�\�H�p�Los�޼H��7��!�y�陬1Z������Si�c�Ud�\���E�D�:��iӴ���=�m�8s��Gү�W{�
0�0�H��<v֚<w�W4��!\��b�<�n�gs*0�鎙��0O�4�B�JXzg�
�s{��2,=/P�s�`�%f�$��N�v~���*�s�nm_��;B���D�P�_nc'��Nj��Y��yQ,]��!NЩ�.VGV�Hi<�B�Z}��p�fUeN�3�K����n=�ݺ���v`{��;k+����1�Hb:���8+�ٛ�B�1_O�s�0R�9���{/I_{�,�In���^�F�\ķJc`��A�ny�������Y��-s����r�x���	J��s�@�>?i8�3�)�h�I�.y����ͭ�LA��=�m��;��^z��O��cF�����y�b[�������<��^��ݽ0W��!��<^!�,j���@����6}�k�+7�'Zƶd�Z��#t{ �:�	�GP!�����֓f!]�reL��g���ɞ�jW�C��{v��m"E�l3�&����Tg������ٌ��u*�=�Y!��i�Ek�����Wjv��ɥe�)�^���(VUJQ�Vo,�f-!�H�6�w 1|+ݕ-����έJĥΛ�BW��Zn���]C 7]�ۃ��T�͎��I�>���®ù��C��7��.� 0�s�8D�D�?�W�-���C2�����d���zDT��F��|�_�FΙK�Ϙ��ڱ�m!�ar�n�ߒ�����z�\�u|3 R�*T�q��Ϗ7�����s˞����!�BĢ��;_S<����i�o��7�V<����D��Ǎ��L]�ծ�<�D=�H2'N6�lU���Z K�T�4l�6h%��.|CԒ�@�1լ��wkD�K�0fxc��+GL,_8�k��p����Vgn1�O�x���������;R���A�l�{M����h�ZA;�����־���o��o��{Mu@�|6H�6]z��&.�c�f�0��P��*&ǽ��.���D�����[����0�X��Z�wY�;5|-붰�3L���[����s���-e^��Ҽ���x.@v<uӡ�)?��	���1�j:ns�f�Eb�/��K7�7�{���p�MQe�=妦�8tx�W�v4����n�4g/k~��B	��4�M���ݮ�g��_{׻�C�~����ŵψ����$@}I�t�wl�&�^�<��*�C���|6��WR��}nǷ~3(�zA����yK8Td^4�ᔀ����ӾX]��<�K����q��q�R��^2��<~ϭ_-��5�y�2�!&֟�hAyi����|�r��*���^Q�3W����Ӥa���X��茨��Z�ۨ��0ө�l�3"�>C:�t���O�)�=[}3n�/[11�!`bY�%��;�ʵq��_
�c��(�ػe��O�\�qA��5r�r�E�,y�L��9�B�
�D���JL\�BN�8����Eb�3���Ox�{�����/=���@j�[ݝ�z��S�<A�o�+�?c�׷t����U�j�Ly�0��'�=;��C�G�W��5������=�77ؑ�C�N$8��R����C��!�KY{:�;ꞽ�vp�Zp�^"��
�[\rs���:����wO�qxA^kn��j����u�j�/^��슿f��e�wUx�
~!�k�����:}y��(�7ԟzH�L�"�:��Tg&zw�4��H��iSaT��]L�Y�IY(�~d��aô���;�Zp�Ӭ��9�f�U0��tP���u
��Zl��W4�_rց�9�x�Sy5��FP��u�����B�R]�[B!mG��r:P�]c$�͗�Զ'�vciα���.^�狞�Zr��r~�vv�ov趥���jӄa��!��˺=�b��.�}�T^X�e��������8�$�$��Np��)n7�b�^λ>����C�cC���<�NN��`za^V��|�?TĠɨ��L�=�OkcI���H��fQ�/�ݥ��4����@�>"�GKи���,��_�G���:ct	2����^R��t�t��z{�uv���t%G�c��ZP��n�A��)Q���\�~���s����JD�F�4]��ɦ�Ӟi��<w ��z�VN,�/����SE�3��L���0ꑭO0K��{v��խ4FZE�U�����5^]B���V��C^�S�O��x�u8��&(�E��h�i�ˬF�W7c�C�o@y���U���;��T��ժ�"�Ή[4}��v��g>O��?}�R1�wU���ݪ�,�̖�u۷s�4>D{�����]X��[M!d1�?�B7���:Tq����B�����O\Ƒ�����`�P�\X�B5Kڇ��Q�<ݼ���^�!OޘA7Aa�HO2�ݪ��1n���S�Zv���=�^[�/�:l3�Va��AY�Az�K�j���ܰ���2lf� 㭱�r��ar�g����3��^��Etd�bk��Q</�ǌ8Ymy��7�VR��w��n�ج���S��R�s���G���R��n(���m��S5�<#��t#�v�S
�DK��@�ZL�Z_�8�!����ֿ�飆�	a�K��ZJzs5S���	��S1W��Gd��Q˞��͋C���Lw��k���16����ٴ�'�!���F�����l����˝�ʛ��A$�|�s��@�1����6:x��+�F2��j�T��"�Y*	},]G��c���:t��|C�(���u�h��]g�)�="~��Y.��q&��E��W�o���_�4�6H�᳈q�'-�g�^�3kid��E���`�����둮���ħ܃�0���Z��lW-4��%t���R�>��)�_4�ZC���ݖ-[����fv�BO/��<�۾Ń���F�C
(,vy�A�$�_�ӎ+ݶJ�~���Uc�E_S�Z���L��^	B8&�D˞�o����:I맧i9��MOI�ePr�;���#��h���,t���ӳ�<2���b��X_�B��%dx^M_���;�gS�À<=/���&���;����$w>ujD��m�����D�ݿ����e,7Sfp��0�f�r4���ӧ��s �;�w�HR%*[�ZP�;����3�3d���Ŵ5^�eCmu9Ûcv�*�<G#�I,[h����Ӈ��Z�eǸ@[����$�\��F���7�3��]�3:�Y���BuK@J�ó j�
%�9s�w�b`��K��e]��A���a� l;�-�\q�9�����a�9+�����F�������u��n����S�X�XE�M��.L{G�tRgS�7�(�>�B�	�NNU1�V���i�.��Z��ҫ� �y1o��K�{�������}�un��m��J�	WK�UE�&u��g�"C{��g;Ⱦ��*��Zm�I�[b�N��
�5�U]�ɴ;R;*�k9����v����ņjz�&�ֵf�+z;t���}�3=�j#ܽ*J�8h7�j*���^����d��oo��}u��e�Pv��dC*F�ڢ,4q�Ņ-;u١"���Z��/��w��r @/s+6�5�A�O}�:k�j$���pc`�]�2���WO����sΰ�]�f�L���jh+]L8��p����)��f��K��"�;:d���a��"���t�5rzfmof^`g:01�՘��yI�fK��LUۧ.������)�7�n�x��%�˷hM�v�N}��;_Mĕٕ!�+"��dG!M���ݶz�h�b����r��)(�3
'�pȨ��f��ӈ5��5�330�|�H���(�Kh(2��\ʘ�\E���T�m�lL>��bQl�`�s2UE1(�Y�9i[j4�b�(�%AE���2���хT����R���ma�\n7����3�[
&5L�U�X&TkYX�����2cU�E*��R���[��juJ�n���iif\E�6��f5h�][1Tm�B�YJ�%E-�Kik�G&\+�Z6�
��l�*�e�rٖj�`�m��I���rѢT���?o��o���?.��;��02AZ�O8hĭ4L�2j�S6��}��;��i���ß�r��4���ZG��k�yky*ͼ����\|p���x~dt�.�`��u�#��(��u��ֿofFaF��KP��d��Hx����{�QPK����.���,�/FI�"��p��0j$KZoVH~묻�&I<�>���k@��<L�
h���AC�B��{x�u=�.��ϭ�"��F�
��I�H�	80"R5u���N���.9[n|��M�e�'�<B�d�r]�{�6�mTn��f\9Ok���g���2S/�Gvp�����$�(h���� �qik厊��<s�_��v��e �[ ���/+Ԗ����Zk��� ���>�u�r5�yf�jvo�[8��T�@�ō�fl�lS�����W�wG�u�Jӷ'bF�u�����s��(5c�Y�NvM=��Fё���G�.�P�w�n��Ј��������Eɑ+�ojwK�.�s�9̖&=0
C��t桵������45���ݾ�px?x���_���ӧ)"R�!�t�
ಽ~��O�4<t��tP�������V��p<�COO�O�!I�������h�W�ic��XC��Ʉ����d���o0O<K Ka�H�0�V�����]6��D��mJ�Τ��a���C܇�cA ���NⲢ�X�|��}��Þ��q{��!�l�C���c��4�0��]_{z�G-4��t��������v�兔���:w��K���ع��;��H�����*�@��
ӎ�����Ǵ��H̭ழ^"{L/)�O���M��vٿV)���v��ew]n������Aؙݣ6n�H��Ea���.T�T�ϩ��R۽˷`�j���9)�?�7hU*#���g�H��Y�[70�Ds�;>���;U�z*hU�{�RoYɅ&�����b0��r��1��8wǏk-���>3m񖇟�ٓ�`.�ڴ������/��60	"%���U�����ݪ���3dX�v�Nu����X����1Z��b��ʃ5Q�"8�:�Kg���?r��Zo,E|���B���0f*wD��skKl���z�������,6XHc��%��G�e����a]��:�g1�[�~B鿽�̓d�gcͪ0i8��x��k��9S~Jr\�����򶰍�a1�/��Ǟ��0Ō>�}+2K��
���BL�|,�^y�c��!cN���δ����:x�y	K�Ҝ�s�����+�Z��&�5�v�ٷ�7͘��P�ґ��� ��D�v����Xx��-��Ϗ+1��}��wب6i!��%J���Z=���b�ͪ��Uu$R&�^�D���8m�D�1�OW��|�_��ǵ�����izsA8N���0�&��UД�C��ս�ﰛ��ۚ�]HB�`�t��I�*�Lt�X����ZIz����N"�����?G��\X���(b������v�������͔v(W:����u횒�x�wYD�O#;Ќ�����<C��D岘���0_0�)�Ÿ�>��Nd�����B�����k�V&z�Ù\�<@GIyI�e�������l�TYiz��^6)a�OܽU�5q��s4�S<#�4I�������k���szƖ]N��n�{t(����7��q�o���7e#���^����C�7����񚃎,v�˜`��kn��|�5��D�����\aֳs}�ZI�c�Ň ��`���b�1�Ҙ��/rm�Z��$���m�0>a�i�-;�Ɩ3�(,�o��˕f���{ۘӅ�l�d5��(zT�Qi�<�������}�����XX#�|G�Ce�6�ei���bi�5�����I
\��L���#�3T��O_��R3J��[��B���L��yX|��d��+���q}׺j[ =��B�\N�$���`rHӇN���Hv��ׇ,R��5{����Di��^B:t8I�3G�:�[x��6�˷1V<!
B�ս(��<t��Hc�kt��)4�����2����y'h%c���6�h����vV�0[��b��2���+z�rO��x�(�p��dx�v�J�����'^D͛����(��m_�]2'�E�r���d-����G��Ѣ4�ۭ�x�I-a��#0GT9z�J��g0�*�c3;&z]��F���(�P����sy�˾���{���|h��&/�W�U�8t�[����kX�.NR�7	�]�f�M׮����<w0�gO�T8>��2�sv�${i�k%�z`�5�1��0�l��I�ޣ����B>��?YQr�>:v���DY,���{�6�g��G������#g�	�E0t�Ц[�w�y��ק�/�!Z���Mᚴ�h ���(5�	0ó�x�����,���5�L�����J�xI��>�;�K�(�r��)w쾝�u�O[r#�z/f�n)(�N-���Ī(��j;�;Z[J�v`�c"ԠkM��Zs����u�m�d���D��Fn�s�_�[�b��tǑt�Xy���v&�����e{�����ky�8�2�ŧ�����*_!�y���0���O͍>v����@�Ϗ���x�\FT���[ѳ���W���]��ҫ�Q�W\�:As���<�r6:�лǷj�u��1ڹo����e1���JM<��U�Q?4��W1��}�<���+9��|F��s�FT��-��Gsg&���nFW��L���JZ@�un�oz���9�Q�԰���H�L�}����������+3��o��i��r����Jm���A�;)�H��<��1MF�G�>!5x��4�禧پ����p�XL��o�~Y0zk3��N��(�D�^�!pu�Q�\�I+1��u��M=��xo�C��Va�w@P�<
��I<W��"�4�H��k&?L��ua�F-ǀ�4��Y�y[��sW|/�1���>�+���(��FMl��U�t�Ug�������Y|��\�Hx��񳮼"�u�{�1�a�>'���
�|�1�V�NT�����+[�%�B�S&\�<~TV�����F���]ӷs�5�w���Ya!����{��-}O��} ~ o����ۣjV��yv��Nи�����ƈ�6�Q�˗IR�z���C���,6XK	w�u��kR:�,�LK��3H9�'U���ǭa�!V�]�Pn�fvv0��ؙ�=��Z�k��\X�
���g%zKҌU�D�Mű�{u�	Tf��Q�����&�s�u�]�@��Ho5���FރRØ�#7dsenE�)���T��s�����M�r({����}E�KlKx������Ha�o�!~Ǥ4�|�E1�͘e���~��U{�f�xS��r��UϬ�XbS�'�a��@�Zȼ�_ޓվ��	�����@;��(�;V羴�>��8��Q�uDW����EMĉ�/[F�gB̻���1KĖ3���Vz{�de��>�w�k�ޞ ��W6R̮��)r�y$p��W�]����iB�T��|5�����>7��n�_q�I1�,>Z��@.�0��i� ����↾���TY�v�ϱadaψ�<��sI<]�zE�V��컻��������>0!%[��a�40�UI���鸬�u����,IBa��ZA�3ϑYQz��ǳ�jo�"�=�~�>I�٠���Lۅ��3����[2_�z@��c�	����\�������7���bg�V��7�5�� �����י�.�8�a�\ya����F�:x�ì��i:�-/w����|��ӋM0����<tр���NDd���3�F��!�lpGN[|E���~C�6����x�6�[JJ�HƝ��]]ϑ}�8k2Z����SL���E���'[����'�\tg!��y��ad�6p���Deg[�w�w�r=HCD�:v+;��H��:"�*''�i�.(�)�t���<EEz��"�i���:#����n�C�;�v�<)��1�t���T��-�>#%e��W��K.�6�\��31�Ә�53S#�?0f�Z�c�}/�X9�"��EM��\Q��U�p�Ў!D�B�Ke�|3�;��3[�Y]�=3�d������lWU��2Ρ�[�`��WϘ�S��VC����еZ��-`WYϭ�FS]hic��v�\�2,�B��g �\���-K���B`�-i�,n��.l���M�l�ld��{w���>�\.�1��:����a��鴓8���ʫ?�T1� ��{�:c�1dhhg.J���^`�be���MQ�;����$剺���u,VF�+g�]�b�$��b2u���tusJ��K����I��W�I��Uf����9uH�oA\"u=Xk�zP*��Z�R��燓��}e�0ݱB6 ���n�NU�R+��zP�]ZN�|o���Hi��ґ�&ð���bkj�^�8����L2+��Je�p�Ve΀Й��"���K�3w]H��W�I�=��^����"��fp��R�B�PzZ�ns�=����܀�H�س���VC|�t�ҿ�T=�u0�G޵B��;�?�#C�=b�$�#��l
�yWU6��i?�ܧ�7w�#��(��K����ՊB���l2�]���ʽ �v�ziWy;A4AB���2�w(C3`rc��j��%�GD��fE�mWp��.��ڕ�*��_�tJ�-��G�D��*�<4b�:}#��wb=��5���W�{O���j�g4��U�mv�J���m�f�ce��n�b.��-�ݹmT͔(��IΏ6"ї4[�4S��,�R��k#�I��ȸ���1�NI#rwV.�ز�I����rh�����L�����a�{��)���ʸ�d-KZR��j�k�[V�pp��V�E��;�
��V5������J�c�R�1j�Z�[�+�P��V�ee�7.K,�]Z��p�j[]6G.�Fdn\S-kQk%-T�����ĳ�\0���%(���	R�t㙆`uk���QR�l����)���k��l5Kq�)h6-�+UZ�j�[��-q�J��ɔ3Ɉ̅� ���GIM5�j
(1+W��q]3X[l[�M]e�0+mKJB�EOĂV;�Zr�ڵ�z�R���}|忋��{ �Ja��T�/f��+��<p�y�1s������D�V�˗i��n��W���v4_��s�mN;-_��M4�d��Xym�.�k�xe-����K�l�E�#$F�WM�f�GLի�];�92�Qsi��˺ �jgP�o��D��9�N#I9�ɭ����<%�2�]�>2k(L6 ������ץp�;����f�L�ON��}a�b���q�)����ǧ��׊�ս��!����Q�M!�~�4���{>v��&yf����x�{r�b��%����XE�G��g��	A�s�>7������Fį2x� �k��N9)����R�Y~��}��ahz��ȟ���h�A�F���xJ�lD=��M�yr��"���T�4���V��Ȧo2Z��R�[QS��>L�޲6��eD�#_6���������f�t���n�\������S�1wk��.�8F�����#y
�1"�JZSX{Q��*�� ���ɦ|B:��2�o�mT9;�R�; jqx�]����	�ޚk�It���Wϊ��H��'���ᣇg�}�2�����x���0Ss	���{��ʖj��/�OK#�i�L�(�Xz�b��b���,v0�.��V��5��l�H����:�T8�s3��]TA�P؉�'Pd���<wʼ�Sa�b�GzUc�zM%��������6\`2�4x!��؆���={~�G�
�� ��d�b[?*���ǈ-��$��~�XMi���Q5�6f`�11��`h{'׉K��+�vΙ����>��,wM�ıS��w����Xr�y,⇠׳z�0Q����sXl���͂�Z�#�;��Y;g<'D̍[��ۨ�F��}��T0H�lm���r��û�'�j����\f-��:��i�Q��tIr�ġ�C�'-Q�G�p��Q_�֢s�/{ت�\C��^ �lyqb:���O8Gken��nv��Ҏ>��F����k����b�r��UB!t�s��M�i������K���䬽�n�ד�4�H�[�66�؆/n�Z���O��sU=OE��`�����8b\E�a��ekY�����並���z`��pѳL*,���קbb14��mq�ʉ�3�����H��<=8E�ȑ�)k)"@����|����� �A��缆�zx�z9�8�b����,�ᳲs�IUe�yuԆ)�y�l˧��4�ٚ��@�"��n�73��(=)�F�YկkS����o0���Q���{mENO���ꎁ�l����N�1��^P�8����<iU�-є���F�NH3U	���̑Ӹ"�t֑]�9�{}�����7h��6Fd!��r��,�-�Du���U��ܽ˨F�.#��p��GI�1Q���)�x��c''s������7���D֭#�}�Iǯ�T����7��5������q�[Q#Kť��1�d�}��]��g�|�����^�V0�.:t7��ޕ�}��CH�s�{Uy\*SDt��٘���L\��FD���n���E�72��$+@�w1@ݢp�����ߦ�(���{/�i:K���/n���%�'�*)�����^���y=F׾C5frN����(��W),�1u��n�т�RӶJ����}0tj��,Y�͈.�,���F������Fp���C�ΒZ����<�8��'��;[$��(�(�\�\2L�.Ȩ�"/A��gVO�'N�ΪLR����6�fj�.���_y�څ�-�������������џI��C�NL|fU�NL���*=�x����%����/�Kd��ii�2�K�1�5��B��Pn6��ں��;&lg1"�6�K�}]��k�Z\��j/���[�]7�N�"� ����l����mp��2(8.09V��]Ü���P�8�$����`�@�����C䇱�Y���4F��v,h[ZCZ���r�}�=�S��(��ޯ����ǢlC���>�����Ő����Wr)�7
�r7�c��pu��S�������,�n�d̬��0 h���Ӓ���
�J��f9������rnF����;�5��(��68��K�j�����E+.��ʕ�}��Ϩ*:FW�:b_k
�ai&��,��{�,�,�*&rb\v�O��D�����Zp��m��K�S��ݤ7��BR�=�P�1����h�A|~M(V�9w����
��.[�CJt{�LZ�C���q��Ǭ�����<~{�(ٿ[�7/0:�j���zR{}����>��!�My��c������s������e_�MWÖ��ܯ��!�@��;�"ڼG.��N��[�^�X�J".|/z�a�g�OD�H�5���6����8�dlO�`N�����w������L ������ȯ.�߽�x�Z�����`��G���N�-��*#g.�"���v}������M����NmL��c�2.�N��(Z�ji)�w����B�H��s����-�������)~a�5N���~�x�Ӆ ��a�'Vt�Z#�������;Is1�6�f+�D���S&oDc��ӌ)S��L��+�ݬ�Xt��y�<�$���|�*�\��Z^�^��Ӳ%L)@y��;B�c��PQ�E�<�
�bx;��#��kX(�ak���9����]߭
���z�^ ���5i4O���&�[}�����P��Nye\��ޣ"��à�p� ��K{���z��t� �-E���Zl��N�O?�Q3+�G������R��d���L��ܚC��D��Lf`ΓH�c��fIt^����[[R^��H�� UՏ^�zxֳ����7ĺ`#h�Uo��C�\�t����a�d˛}��_{�)$��s������.L�W�^�{�wj�0���{J�\1z����6+���=3P��,�
6���z��2�99�K�.&�9��������'�`}�гɗ.U��vz���a�HF��+KKSRC�[���l�Q��0Z�k�߹a`��v4���r�kD|.���[t��z[	�><�X�rC=�k���Ӂ�o�C,$秏���YD�չ$Ne*(u���;ٖ�$��d��dܚs(��cN��	��0�=��R<�����cj��M��
^��`�՛�XШI���,��}ʅ6�:3c:ފ������S:3��;.s@cfn*���B����<�!2���Iq}�@+1rb>����,̺�F� X���-��=�Q@v���ˮ�!S��fh��-E����8*v�L<�b�6O/n���.P��c�Q˔�ݫ�y��R��a������5�}P�Y���MA��q"s��I��P+Vg��S�n��e�½��s��g��F���3�t���n�id߹�"+���KlA7�D�I$J�˂z>�f1����4�o~&�s���c�p�}{�e�W��dTL�S�O��~��Q�e��PR�r��	������V�)�	�Wx��bC��X�\��+`y4�ug;�G�����6Jl�d�U�8$R�\��7���g����D�5F ���I�t]N�E�z�sWC����n�Nľ�P�c.�u�[�<u�+DҶ�n�6\>����!M��V��d�x(/zS�1���8C��b�0�.^�ԝc�u	���ܞ=v�z�7t��yZ�&�f2:s�+���ו�s�s8�|�7WK!�l(�}�F᛼�C",�2���ѡ�ث݅R}��%��jjA��*2�����7�!�&#�Y��Ɗ�Ｒ�R̉6"��`еB�n��n����=��JU-��!R�V� u<*n6�v�����y8���8�n���Õyi��o}�X<v��$f]Z<�7̎�[��`U�5.���TMs���;@N�Ε�Gpa�:��U�QO��G�n�9��o��3�BIĴ]�g��A���M��\;fM�U�`1�B�%W�Es¥�j�͙�[Ý�8l��N��UM(�X�Y���)�X��t?���X���q�A��"Wu��3`�F�ݜ��K�7r���D�Δ����T[�:��x�4�K�@��qi�+���B%j�_\շ���͘�A�b\��v�}Y�a���v���vÍ�Iٖ����d4����A�V�l��/��1���u�S�i�Ǻ����N
w�D�抻��`dR�H�ƺ��o��fd�йO�w�:��Ӗ^SӃ��K��\��n���f��+D=}V��5�]k�ڦ��s�V~r`� ���d��.��2��rPKu�L��f�1mc��E��7T'Q��[6Ὕ��yOjf�}V6� In�u���9��|�6d3.�x�"r�2�	ۤ%��"Fn`�Tqe�磨�
��f���i���驓��#jfL����j��'����c��j�`��*�wn'������XIٱ1X��jk�^����ث0�R��� �u��aBۢ���`�& +��h���;ġ�[KxJ:%n�Ŭ��B-�ty�'w_9@1�P�!�,s�7���Drq��$nl�W��3���Τv�VM���ڪE��\,|�f��� ����Y�
�KT���������cS֌W�,�L�3ѢZ�kj��(�K+*X��un�MZ�*,M!T���X1n\X,V8��FնUeh�����ʋ�Uc��i)��(���"%�DZ��E@Qcm1��F8ذ�0���bֳIX�1R�KejV�0Pb��i�E�*�Ad��.�QDR((�%B�(��aE�2��+Z�H�
E�A
���Dji%Uն��/IrʄoW2�(��AV(#*�Y�����"���w�o�5������W��&I�v�G2�_P�b�8��-�ܨa���¿�����r�VW���:�0�2���L~X��7Ԏ|�72̋<���w^�d%%�ޮ*����֋�ד���8��+uw���1���#�"k$��8�u:�0[W�Y٫U�x�D��^�9M�"Xp�2�c8�1�ZU��E����r^N��u�mD�1��*ˁ�N�T{���i��!K�[��f���s)&K��}�����N���Yo�{�
y�^�����b�x��:/̞���7��OhGwB�����9�� �ftz;�[OL�e1�&{1�NS��,�jg�NH�ѭ콳�)�o"o�j2Nn��]����tfG�,�]Ȅ�S�%�X�Y;�w\)�v�i��:1��q�Lh��mZN��G:>8�}����t��0���_7�v�-f����o6�*P�����P�j���(��!���\	*>^�P������{>��=%���Oy�w�S���W��Zt1��_.;jf^�c`=w�a����c=ue�So}�g��.#�ME�{u��2^whr�p�oѴ|ft��">`�����T�i^���n�8�5���e�-�_l=��6�~��wU�̳bB�t�;mٲ�`[M��V�v���9i��:���s&����O��G��w�4Q�����Kg���>��'�/��8)U�#�΍%VN�$dʣX��8��kf���1/�Wc���Z�g2�Nr��&�	�\���n�ޒ�9P7ql6(�Qfeբ�SS=ڞ�+�42��{k2�R
�Z�������O����/�Z/6}t�˝L�^����ym%��vfÅO�r��F��Ky}��-_>���݇�t0Ƣk�����A��S~���p�"��x� k��-l��]g�t����������}Vh�g��֓\�)Z��ỿ4�j���Ts�E	�k)�-4�f�K\ֳ�6��6�H������J��{�p��ݲwTg�R��X�o)�e��5��Vs��\k����ͼwՖ��.5P��[��Ժ�ĖU_?�yo�f��;.v��R{&5{��<��<���y� �T�vc r7����y��{�u��bmr�׏�=%��I(5�tq<s�4�,�L��@g��ޮЃ��sb1V��n[n�[�L:ݵētu���#7w�> {�D��NP�Y�e++��K�8����:��_���>�[=��XU`��[d�ȳ��N���؄��,l⭾�p5p��I�݉t]���]��U�S��;���Gx��Q@�Cm��W��t^���' �J<��G�(��׻w����E5V�f����f��W�a�oz7���ɉ�����^��]e@_���?T�952\ůx!$��,�N��v�%�/.��x|<�N?"�<��˨��xi�S�<�LU臣4C5���v���|q���[��0�&��XM��jAݗ���!���6or)v�\��2�K(��fF5������x�E�Q�`��c�7:p~�^t\tĝ��y��6x�m���on�Ov���Q�K��Ӳ���1Bp���Y� �@E����oW��j�ֵ�A=Ut��GEY�W+t��Urg<��]q���@t��cw~�[�3�H��e�x�B��-	�PGBkQܷnԪ�#�:	�;w~��5^o_��=�qyɵ��P��5����z��0m�����=w��F̯l�}=���Ǆl��p��B_:�o�@�����Is�f���U���Vl��(Р�2��EƔ1dk5�����h�������Qx�AW�=�cY��U2���0���^swZ˥o��I�z��x�X���}Å-��5ۧ�N��=�U�r[�M�F��ѫA�T�Gs�!�N�l��#A����b�wz���Y���C���.j���|�U)����ӶR�Uf82�I�s�i5sΆQD��b��Z޲E;}�؆�pE�M�G=Z�*�[ךN�w�� r*4z��B�B׻ b�2♩9V�B7Q����� ݠ�pFv�*�':{,�o�0����:�IqC)�7��oD�.m��HN&�~�e��m�g!C�^�@�EÁ�.&��r3ٟ&��E������w���Xo�;����Ѣ)/V��U]�v�nd�k�Z��BZ0N���tk��h�Rj]݌|-d�w�^	d��D�<��*��u�G�_Ȯ�]V5��h't�pܪ��Dj�r��͵�v�-�p�_�������١Q|�i��=�=�K4���4n�=x���@�#3�JU�=�.-]GMX�O�}XTӵ�����������{]�>�MB���j6ҴΕ���=H^�Kh^���ګ��ޞ>(ViP.6 ��`�z�+v���u� �!�x��ix��b����o*�1��1j�z�4�<
�����3���T|I��ڤ�W�_�:����k[��1uuω����J��^��>�l����b���z2%�ٮ(�K$���X��:�ڬ�h���rl3Ⱦ�a$5��'q�7P�b��u��h/N�<���"3E9t�z`�]�ΕTwW���)�3%{(��ih�l��4�Y�ݠ�z-u�":����)���N�ZhQ�q[��eLھ��8^�a�6�>�O?�q�;��X�6A�O^w��/���X'U���s�h�{���;���5t���B�}b6]Gr�f���u�eO����5\����꺙�'ۢ��6��G�e]������%�p�3Ŏ�c��Q�Ir�K��i����	E�,�ˁY9wf6̮�0t��4x��u�/�20y����{�x�1�Cϐ�4^�wX=��V��
��9=`�a��&<�F������->������u%]V_K�ne��rLvQ"LW]��K��,.�e6<� �*푈n/�;>M���3��t�),��GD�Ƒ	]b��/�z)�{c0I*ox�	����sm�V�\�*�YjMF!�`�Mq��$"��U��J��WL�g��vM�h��.�k͘ܫ��B�Vƙ^�#8�}�ـ�;�Y4�k�1IRN;�P	�����5�p�^n�_em��ۨܜ$F��8�v;�p�BwF�D\����L�P��FC���\a�������=��b���T`q��mc�HRy�P������I �{׵�,���J#�)6��e;!�7�X�A[�d��l�����q|yLUQ�{�E�B�К5:��T#�:��Ue���(�(hS��ҋ���2�7�q�}������x-e����<=�˥&�Ke�=P��^2e���}�*=��D�J�1�7.,��t���`h�Q<o*����%�X�t�,��Y:�j�Ws��o���5��;����ޠ&��zʫ�ar0��7.�w>����b�|N9���빋i��x����tF���PL�δq��x�Z�ǹ�w����5�:����J�P^v�kyf���k�o��� �����3n�ێ�4#gy��b|�c��F�M�f���

�N�J��d&���Ճ)�D�5����&|�:�V��� ��8�c�6���U7�y=�C�7��Y�8^$��zj��ѻ�F�\v�ѫ�"�m����7>����:�י��-�ڛ̠���4�!D��ؠs�n�*�>�G*��Ru7x���e���: �ۆ}�����9>�uKނ�X�/9.��X�˾��\��qu�z�lb��F�|'86�[���oZH)
�lɛ2��&�nX�2]E�88��x� �EiJULpX	Ȟ۹�Z�F�֤�Ƹ� ��J������큐�$�$b�R�Ij��Q��J]`,
�ӈ�#���*+iTA`�%q�SL��ZYF
,-���he��1+
�Q4�dX���cY�Z �b���4�XEDU��(�6E�UEAE�c(Ȣ5�AAD�	�5�!�
�B�
���,�Z�D+TUA�Ę�TDX�����(,�@bŬ�)��F��!�:j��QeH���"E������2�߃�\����T��Nbu�Ǜ�v�A���L��'�=p�cyTn	�]"�l�6�|Q~�h�W�*�
kA��B���,�W�gk�ǵ\Ȫ����W��˗�癮�g��[��/n���[�3W��ek��ס���ɸ�)�v�u�X�zrȆ��(�"I�̲Z�&��(�Op����m]��;yp؋�B7.��\�.���k��v��w�C��Zh�{=��ͅ7�KV/Q�2 �\��6�e=����Z�:F_@�u��r��'��l͝�Xc}n��	y��|Uۮ������w��HEw�|Q'����չ����j�렑H��Ǵ���1��E�.�@�j��o��(��3ϋ�h>�Ⱖ�9�����v��,I��ܩ�/���|oH�oQ�My=�xT���7��-g�?daH��C16�F�o�������]�i'�V�A�W��~t�9R#s�n냈�PD�C_���Ql�q�^R�-d=����,D���
׽u��x@�Q�|G��C2��'�z��Pޣ[�{��hkk��� �{K_�~�?dߏ��<��/�7�o4�C��cN3u7�L����{��\)m�瘲ņ���Rm�Kg�v{.�~�8xt�
�׽٥��ol�u�`�,@�p����;�b�b�O:�{q�J~�ҫ%?Y�0�t�XV}���8uD���D�����.&�%�gcgi�x��ݱR�M��q$(w�s�I�u��p,^�\�c��$��L�ol;1Չ��|����q4�q�^�<J��2�ژ?L��NPyg+�ڜ�N���k��˺l�4T�:�Wޘ3<+=���gX=y��#.���(�EY�HGA��ش�Yj7j�*C�wU�8�ц �^lYʣ�C�doXw>����r%�V�A�)cu%?w(� �]����ez�r��A�Zi�c���ɨ�"���q=��l���QN��]1b�54{]<s{@r���yDk=}pc�![��;�=��ܸ��Y�ѯw5WltV�VV�N�=�L�'�YG�{��O2ʗ4fy�<KlN�}HEf��=�d_g3�ᴙ�Em�z��wXj�����n-�k�یS�2kv�d2����;ֻ���Nv:�vٴw���b��ҁJ�7��J�Դ�'��:~~#���o������47\��AB:6�g^͖���Bт���#�L�4���32ƹqb �-7���lڋ�)*Wq#w+-Wmpb�|S��6	TegN���P�-;�r��-���N덀n���ȉe����8F뛦"������N��=� �M�������Ɣ�ی[�]E��sg���]ے�Ym�TvK��F���wm���-C�f�U�P����5��ʸ[��d;$�N.��tN��q�z�%���&�4��km����b�Db�A��s�WB�Xo��{3�C�Ew�r��ZU��߷�N�KO��ST��V�\��(��\�&q��ܳ��C����u��*s`-6e���s�/W'��;I����5M�dU��V�����ϯE�|�����5��D��%��o��_Upz+�N�sX��=ԙm�W��b!�f��D򜸢:w�tCf�W>z�M�����nQ���U�����:��l�4z�z�����֦G��\�^U�{��;q6%��6�52}�d�]N$Ye[�	֫DX���g�)����G�w����!�W�ݵ'�o������R�ˇ�_c⼵��><=H�`q5�v�xqme�DcW�����\�F�W�� 4>G�i��ۑq���xg�(����ۮ���g�w�qZ/,���'T��7�����ۜxm�p�i�f��\/p_,u���+�-�v@�75��gM����M�1$ǦΙ`]N����=o<�gF��'U��y�A�e_fO�����F�wYv`��˗�~;���U-{��\��)�Q(Z3�Ũ9L{YV}�yg8�.����5��C}Q�dg3���K��:�^�ٰaC���xo1��Ջu��f�B9�rU��"�P���Y٩S�b��쳎�mos7)ve��:A��u|������ �m�Ph�GO����ą�u�y� M� �[��'�QdEϻ�}}Y�o/}��^kzھy��iR#&��
x����l,;S����ɲo�k�G0�����x����s����I�����s�߈(&���1�2��z5�ךN嫢n�GA޶6�z3�Jv�I�{hiP��uhz(���t�8m�N�r��w�;�L�'�a�w$�n!ї"1c�km۝��W�
v6b�6 ��țy�C��ҫ��m��2,�wY��׶g��"�O'�̻��z�g��\ksE�'i�q�ɋ� ϶f�\ǈ=�D�w�Y]�1uQd���;�Z�	9­�̃�p�q �7��vHmZ�wYR�Y(p
�Y��+Y�7B��7��-�=�sUkO�8SjV�WVsT����c�8Fd(Kl����mw���f���٫��'�o�P��m�LNuK�9WI�^X��x��q,�BvjDn��Mo;=o�Y�FBpMd����m*(tl��l�@��H�4�.�)��h��8�;��[hB�Y67*6�mڳ t7��XwAR���������=���þ�0�no��$�ų�����h3� �0�c{�:N��ãz�����q��ǜH/0O<��&�QK)����ǑgF�Ŗ�+w�.Y�y��0݇�;�iw%١���;f�*Z|=��ت�S���t,�w�W0K4J��޻�%I��'��ȶ��3{w������[^�wY7���D2���W�^a����8I�ެ��{:���W;���KZ�vj2�镯Yi�S�t���������i���.�gJ����ʽ)��n9�<��Z9Z&���0ϱ!�!��u)I#;r�)�{�U�_��x�ȱ���we��ƻ�m�MT�U�y�0�i�XK��Ue��:]�z{���-��}�f�{W:P#���;�Lֲ�>��uT��(�ϐY��6�u�]�d��gpH;[��u�m�FoJ�,�����N>4��l�>�+)q�o��m�e��	�dz8� �x�9������y��'�w�k���T���|�S�խ�NؔzFl�;q��g���ޗ}��
�O^���i�}�ag۬TY�WL?*4-��u���5��"%����6/Nf������<�sC�A�|�U:�xM�z��L�߲��\";܁˫� ����۔u*�E9���];��n��!ۉ+¦�l�S>#�G��R����1<=����6ag; �9Mզv+k9���-l��WmgtU}͸or�#Dê�f���8��z]d�d�k ��e������s��b�u�bȴh�7�Hq��W@b:Sͤr��*o�6���'����j���v�Rw��$��ɻQYZ�����l	��3�19a��N���z�V���|o�Bp��hT��7ɍ�d�CY�o99y	Gi5�b�7Y�n�_D�Z��{�ְdt�tYA[�\��|7dsw��f̳;�%��R*7Ϝ�P��z�3''ٝ�pD�n���i �|��6frk�escF�у2;M�N�x��u�	��y[|�a���)�z�G��o�='���^��/3h<�H.�V33�=�o�7b#��r��Ӝ��
�����ʙz��\%�$F<���B*Х��J)3z�tsy�ܴ�Z-k'wVmnS��v�+;_Q�<�o3`�N����?�+�zs��.��]Ǭ�dR`jF�NTˤ�D6�R�+ 5r���qC@�;h����N{�<���D�
"��Db��V
,��*���Eq�,�qUb�D;K�VAE$F-aX媪=%V�A�V�*EV���t����1p�M$1��D��FI�u��S�T/WadY+
fd�`	i�& ��QE����� ,��"ȌP,'IPU^��t�%AV
(,QAc*[La��0R�nf�(����c
b���ٚ���	^�!-F��Ȣ�:���:f�;)K�H�I�u6���H��ͺ���`e�gV�J�����&����9`4��.z����ޮ�i�j"T,��탽YJ�>��<��)Sb��z��Ңs�	]�uQvY�L(巚�m��Ҽ�j�[]�YU���C���B�����>툅��U�e�Px,C��7�t��<�B2�o�ځ�9WШk���ݙ���;eb=9Y+/�xxР']A�q��"n�&��5g=��r*1Q�hD�}z}�o��&38/�zWf�ݡ����s/�_Z7�ߗt�Yx�Ȓ�F�lg4C�������+�]w��^���t��_l
���Zp�_	PqLl]��5�$���NfV����<6���/�&ޭ�d^�˧D��E��_J�Х�����i�W�!��ͅe�맕N����e�şO��+�m�#���C-!w���x��=q#�)���9i���ޚ���f�K{�ԛ�h��=R�r]˚aR�`'Wyl���=mu�]cu��{Ү}��O!H�v�h{��\�"= ��4M���&#�Ji�N�a��=��E���Y^�u�$��u�/+��}�o.a�{�֯��[�F�%|�/$�l���ُ͛W_�Y�L�'�w'Hmk���d�m�v�Vz�CO09Q�dwOQ�g��4x�z��ś�v�Sw��\�˛���e���/3�k�M# rܝZ�Q{�e��t5z$�//vYZ&���l�;x���T�]��E���9ȳޛs����X�7˯����;�	FR�{��b:.�v׽����*����:��<w��s�	�[m���4\p���	M"���x5D���1���e�/��r7������:yM}�.�&m���Y�����1�F��O8�ѩåԭц�M�X�sh�[Y��ü��t�q����;��R�1�oB�1bˀa�=���r�
�)�f�<�[�""Huf�Y��[�9c��e\�8��#��vE;�s�s��S�M�8�N�O�R�^���?��_�I�����r�oģZ��`����hE�&W�:1�|�c�y�ܼ�r �=�9ׄ+A�@gxk�Þ��������W�(�Vh|tf9O)�t�6w��9o��tȮ�,ll.��	}����R�ɳ�'�R�|j������p�����W�&z��)}5�cB�������{-^�k������S��{�i�� k����e��d8> �:ӕ��u��u�d	 �k;�nH����6J�d���y���/M�W�tC�D�%����
�����Q������H�;�sa��H�}��&7���X駝�������]��{���ʾ8�adt�w�{�aXa~
6�M������-���16o><<ԍiA��9��L,�=rMi��1Ū]�x����k�а��F��T���
�وV(ͅՙA���D]�sS
0׻tpk�R�${&0T'��ec�n��*�@9FөC�.�G��[7�Un=�#q���rd��KӶ)E`�����v�x^̶DAkΤ�\[ӌ޼lN��G��-�Gw�$t��BZ�v�ɽϋ�<4��f��27᪪�Y����������xG�	��x@�f��<L�׎���Ykz7����d�j���e��r�	�'|��}�-Gl�r��~S�X�2�L;�+�N��'�xgB��@~m����,-�Ɍ�0	��Ocic�M���ݥ;<�sz�=t�(�o��5�i�wT�iT	��Bz�6���]c��O^~�)9��o]].��KuQ�P0y�*��!�{���3�2򮧒Kjg���V���+=�3�!c(F��V�S3���4����8����:A=�\ݲG$���Y7�����#����S��f��r7�6��\�K(�;��+����<�UE[W�OZ������O��}P��؛�*�hX�njz�sò��և�7��{����[~��~����AH=\h{�˨=����K��=����z��I.��͟,� �^ޝ��j�q�$MޮKԷK��V�c�gGYFo(Oy�û5����c��Pإ��O��KI���y���>�UfnNk�V��]5���P�����^��&tDu�wɽ�9�JƑu(ͽ�Г��n�ɜ`��`C���vc#����T�5g��)!��j���hR�͐��q�q����g	��k����[Ì�k=~{���N0�ӽkZ��/D<�O7�u�����n�}@4���<ŧx���ۑ��&]2��쵳�r��++�[m����eE�]�ޏ��=� SV��/�ZJ7խ)����>��z��e���_�[���&8�=�c���}�����8W��~�M�)�����r�䋫��.��*�CB7��|�L���U������������V��A��E���l��Z��'*�!�ԜV�7fi�4���~�z���� �|c�-h\���w����ѡۯ�o��Zb���rmf�zU���㽓�YGwƅ�����yr �iķ�m������,�j����*kU�+8��E�<���O�@�5�jIuiU�,�~��o�yTaYإ�Q��	���
P=䷬>��3�f��~J8oy�{�ʖ�x��󮈇��i�M�P�n��u�SU�|���;��.��ɫ�@��tom�1���PJ�|ޕJ+�����4�u���n��A\Q�A�� ��÷��'7:�|F[�6�n����A�/���&�=ߺ�\���1&{�*���.Gu�Xp�gf����{9uξ@���P��0#s�-�u��C���eN�fk�d��c�55��ݷ�a{X��N�+���C���;At��ϓ�g�Չ{�]�dj�ܐ�����b^'��W�E�y-���ۮh�ѕ����q}nky���;���]j�49�Mm��Ȳ����gc4zz*v��p�-�ʍז˽m�9��}�{W=||"*�߉͚U
瞈�y��)�=qoٓ�:�I�3My����۾����eg�mݑ�w<)_?M7P���+�w9�j���[��z�&�����?�������b��R�Z�QT����D���g?dH=^�Y5D��a���*)S#�,��P�;ɞ_�P,4��?I���N�5�	���@aD� ��"AXZD� �!$���hf���']D褳Ľа?$O���?#5ܯ�1�ZKk�{Ӣ�$
J�՝Uo�c���܍��\��k>�)K̤ŉ���E�Xт3?v��e��//����x��<�XP09�::�h<�~��;����&�}���0��RfI��*��]���a�V9쟞D�#���m�?�����9��n;�*��LH4>�=��\�;T���ȹ��T���]�50R3�%�~��k#V�{Vb�$[�kw/���z8����TUL���s͑L��+�I�谐 �&���g�'^�ä����D�H @5�s�XjI=�R���)��fu\��7�L�#�(n؟�מ$�ș)UU%�Y��Lx���M���bץJ�{�5&&��Q�n����<C���7�,�|���&_���R�������xq<�nd�G��p���&�u7�p���c2=��y�����;%V)�LI�;M�Q���'9����{L��@A�u�J+N^����I�m�4hbh]J{ņ�Aע,�kH�rH�
)s���'��j+�D�J�#��ObXۂM<�h�,H��<��u�	!�T�@����QE&�yup�J>mI�Uf-&+I�f)#���LF�MxW�w��(��'݄Hd�����%��S1�,K�_M0>�I  �.w���-��t�
��k̓��Q�s�R���mO������8��7�\���q�k%|]T����'Vök�Q�b%�c�F;cH���,H:\�z+�J�J-e�w�{ѤW��ZO^&]�i.�Ϭ>�Q��{�~�i�g.܏G�zўCE�R�OW;0T�%��{r�>>��᩶����kQ��:j����^3MMg;��7dH/�֎H�0��r���ݙb��OFe��j7p&��Q�QeVgו���Ac֘�wl��%!��$�B�Ǌ5Q#����������;d�w'��06�Gge�#edY&���w�^{�R7ET�GlS�G=���8L��H�
�f�