BZh91AY&SY�L{���߀@q���"� ����bGw�          ��*��ERTH�B�(!J�A(J�I*(�$�R��	IP��%P%$	(.�F�U((�3g��*�ҴЦ�j����
h
[-dՆ� F�Ҁ &e ����)�!J ���`��l�J� �:�h��*��k�@I!X���[3-h��e"�l�+l4H4i�h
[V�@P������ *�  |��	 6�� ^  �gХΘ ��� n��� !��� �2
%'�i�{�'] �ݞ4X��h�WϩJ���/�� ����Zil�6׃�8*���Q�yޞ��j�R��z��ҊR�x�����_��w˽
hQ�{��_>����z���ۺ��T�PkC�|����3`ٛ歹(y6��5�henU�:Mg�{�j�w]�@������y罥@Ul�k�_�j[o���V�k��8�}��Ҁ��¼�y�JO�KMIL�� i���R�s����Sk*���xh*���/'{MJ/o}�}zh(�+���mA����+�h/m���z�5P����Eҧ��4{`+xwR��Jm�k 4R�c*��@[��)� |�>��K8�ހPzhޓt�����j��݅()�^{{j��X�\m)Sp�R�퓤�;`Zʥ�{r�I�kk�.������Mf�v5@@���R c�ҀG���89Qٕ[v�۞z�5[j\{���j�UoN�4Р8�t�E��q��ڕE����k4�G��6��j\S�{m��t
�Z��T�Kl
F��T� <����N\�TSls]p�R��r��֩�ɫ��N�)�i���y�P�y5
QvpluB�8�G@����Pҁ��>�� �w�U�㧻���=�᣶(v���At��UEY�����Т�,�R���;r��;i�UK�) ֲ)���_>����!>��\ѴP
v�����U��:��T�GwJ���̂���.�T��U��TR����H�W��5FThѣZ�Dd��J( ���T��Q*-�N5@�hhq�4�RwvJ�UU���T]p�T>���IT�6éry�  URUP�A!( ��2�*@#L  2i�S�ĕJ�j      ��"���     S�	5ETh�!��@� ��H�� � &�h "I��)%6��L�Q����4�O~o����ѝ���N��azcC��3�MQ�g]s���~r�~�=�W��P@`���TT�*
���c�J@Xx	�����O���8_� 
�?�RI$֑^�8S��������?��L���0)�lb��6Ķ��`��6Ķ-�m�lKc��)�lb[ض���%�m�l[`���[����%�-�l�-�lKe��b[����-�ldb[�Ķ%�-�lb[���m%1-�l`[���%�-�clKb[�Ķ%�m�lK`[4��4��%�-�lKb[����%�-�l`�ؖĶ�m��ؖ���6��%�-�l`�a����-�l`F[�60m�lb[�6Ķ%�-��lb[ؖ��%�-�c���%�-�l[b[�F6��%�-�l`�ؖ��4�b[Lb[�6Ķ%�m�������%�m�laLm�lM0m�l`��6Ķ�Ŷ%�m�l�[`Ŷ!lR�6�٦6Ħ���%���-�lK`[�ؖĶ%�-�lK`[���i�l
b[�6��%�-�lKcl�m�lb[�6���-�la�6��%�-�lK`[ؖĶ��-�lcl`[b[clK`[`F�cl`[�������%�-��ؖ�Lb[�Ķ��K`b�l-���"��R� �bl-�LT-���Kb�lDm�lm�%��"��R؈銥�T�*��F��b�K`#lDt�؀�blm�-�R��lEm��� �K`lPm����(6�� bLm����"6��(�`l[`	*[b�l@m����(6��lc b�lm��Q����%���`lm�-�A� ��2؂�b+lm��� 6��`�lDm�-�T�(��Fؠ� `�lE-���LD�����`	l-���E���� [`�lm��� ��V؀�# B�"�[` [[`([`b�li�-�E���F��Ŷ��F��`#lQm���E��"�[b�lm���-��lt�b�Lm���� ��V��[`�b�li���� 6�F��bl� [`Lm���Q�����J`6�V؂�-��(�� ��F؊��`�LEm��lDb�[[b��A�*6��(� [` [bl �m�lb[ؖ��%�-�`�ضŶ�m�L��tĶ�-�l`[�6���l`�ؖĶ�-�lcl�bS��ؖĶ�-�lcL�i��-��6���-��-�lal#����-�lKb[`[�lbi�lb[ؖ���m��0-�lm�lKb[ضĶ�l[`[ؖ��%�4�ILb[ؖĶ�-�l-�`[ؖ��%�m�lb[�b[�6���-�lK`[�l[bi�l[`��6��4����ؖĶ�m�li��-���-�l��m��Sb[LKb[�Ķ%������Ķ-�-�l`[0�%1-�lb[ؖ���-�clKclb[ؖ���-�2ؖ��b[ضĶ%5�������ۭ�WjS�/?�ؙO�����4PJnܒі%RZ�]]b��7f�0�fmˎ�j�����lN��jK��w[E����bz��4ٌ�iMۂ����#���<%��56�]Y�	I�ד1z�qT��q�7�#ht�N<��i�ֹ��3!Z6��iՈ
��9M��B�k�NG�噌�li^f�q�EMR�-���.�y6�Yp���;wI��6�F���Lۤ���i�/s��ښi�X���@�`�w��&� .Ű��r�f�J��C�j+WnX�8�ԛ(x��]2��6�N먐Z%Z�	24�&3)i0�n�I��"���F��	*��3�6��٭�k%d�Q<b&�͏)�����s`xUײe���5 XWZV)�#ZU���n���.���%�J��L�,+v� �KV� �"�r�4TI�n ��L��`���nP�v��뻂�H*�â����U/:�3�Gn���c�� �fY�AT��"\u�m��o3^=a��DK�f��q�.��eiPRH�OCܤFE�1mZ��z�S�<���t��;��FL^�ɦd�Ъ�k^�{@��ṵ̈̄�H���1:1(�:e��X�����3)1ɦ�bLu� Y�VC�u�����)��b�Z ��o,#��*�ު��EedX�U�Cu�T^ɘصF�v h�NK[�v�&�-��HhKr�CoE�-\�*���T.^
���`M�)k�2+=ۙˉ��%ݛ��a�r�d�+L;;2���0^%An�)�F��J��zf�f��$���Lwe(��@PʼT� +Hڒ�r2͌�n��ݴ�іl��$�vV�)���&Ɓ�[�*+v��h�� �f%��Z����D�a����Z놖��d뵺h㫺LL��,j��Y$%b�y�n�����kj-ݐ�*m��C*[M���×�	ol;�+C٫�*��&��ц�4"):��-إ�X1�n��8(��e�67e �2�,�2��+h%r��1aÌjr̫�7���O�g/ne�b᳈W� H�ȳlE�!U�lօ�d�N؅ф�[�J:uch�v�����ZQ!{3EETX�+uPL&dJM�WY��J�+V�թ�j�iށ�f�\x���gٹ�P$v$0,"��+w@yy�ҽ��5h�ɨT�hB���y��^ҼШ1�̔��֘�n��F֪��7tT!��gt�[��^���V5l�Z��.x�� �q��6+e&�lj���jR�Qm��f������qd�Y�JiJ̡��\:��YP-Q��h]�G���ɲ��'-Iw���(i5�y�=�R�<��`�.�������r]6b��`lm��
��؍�����#b�r�lZ��Y�Ӷ�����5��J�-X��`m��=�[uR��A7xV�+o2P�J	zflw�u�����n���/	�e�Gj���ar=��#�w6��J٦��a����6^��pu4�v'�X��;{cVڬ�4b�jGjC�T/6�v@��,���9�ͽ�f��IyN���:Q��Լ4f��Q`��=p�֍�72�G�Rd�J��N9��Q��n��WY)�&�Qȣ�.�гF4��nC�օ���t��&��T��݄��qL�71n��m"!
��+�f�Bk!��0�U9�0�MR8�Y6�T�^�8h�h�Rf����&�d�kM�ؓ�-/0n`<�%��{P�`�ہm�6i�a��R��_(r�c��.u<Y����)�Q�6�+A)$ȷNؠ�i���<\x�Mڲ����z�ڋ1��$�m��ŗ$���/t1���̈́f��%�?-ǒȼ)
a�4F"�!�l�^m�f�;�;{n��	ٳU��5�4��a;����P�:�r퍲�Q̽L�HU�-�P��*ݖQ�!Y᱙6�z5�Z6�!�6FR�\��(�;B�rJ��D �Z�+Rx�����)�qI�c�7��BV�a��v.7����5�J��l-�ʼJ=j��/MQaf*ӲF�).�7Ct�5�"��J�<��N=v'��v�q�Z�ghmds,�Ճv�4�*9����40�h���-l7��CB�m^�YhJ�{P���J�e��v�{)L��;;�;�^d�Y):��%V�8�m��Z�J��Z*d)�3Y����@j��2�����e!x$Ͱ�˛X��jJ�lѶff5�c�/!N�\�5P�SFۣ��ЎU��f嘓���{u����6a���рiN�i�è����r����;j��k)�:�l����!�ԕ��PC�nkrR	�1<�o@�-�DK5�N��j��[1f�h7%�+B�a�rbEŋu\��lA�5�"X�fXD)t��2�jJf�D
����*EN�[c/8���9����턹�m��i��K��`�7v����S�H]e6������i���uQ|����O0�.�)W��h�l.�ޔ�9��7h�;���,CNz_5`�6;�3LT�hS͊�2�3vK̼*�6J	��5fڬo6�*[��e�;�TM�9R�6��������U,�i��[��D�{\�J
e",b�s��ҕ�%�Ŭ%	]אʘ5R�iJ�F^���A���4^�Rb�e�H���]�����R��#2Zb�4ޱgAg ��Kxo�h��.��[Rjhk�BKw6�Z�D�-͋Y���+zV75U�V&ܴ�-
����db����S��p�w�Y���" t�iK=��K��5�G%��1���!tS���6�$�ݧ����a�j��0�Y��CR�U@�w�V��2�+�j���n�y����=�gm"Mmdo`ww�^n��C��A��d���e�{��N��Z��K�Y9��e���U��������nk�t/4�V9�V[��,��q"��^�m�b�cv��Bˣ%�KsX��M-���M�����]­M�J�֝v�j�4
#fAB�cf=Wm�������db��C	Ŭ� �5�8����n�ǲ�SM��[ŭ�5��I&��]D��d3]�g+vM�1f�n���5�[��l�dX�ɷ��ؒ���ְ��(ҵ3I;����v��u��k�n)E����GzF�hnS&h�E5��K[{e+y�2�qlo[��]IW
�φ���.����2��K\/���hЧXI�)2e�4%�vL�B�i�h�{o/�&,�[�D�/���\����Y.:	ӕ��Ų�D�!��Hm`�(��];݄��D�È�ow0���0��Kg),�G� ��!]^���2�U`�Ā�;j�H�tY����$��+��롛 ����Tp-;wJ�ڷ�Y��Y��;��]�Up�q^^��A�Y�\��_��-���6Ề�s&�lu��H���@ɗ��"�0p��s�їGV�.�ư��Cm䙥(Eї�Por�]���������FZ7��a�qK�m^Zz�[�^�z`���:�����8� �6V�L�ˊ�+Ve�Q裌[����ܐmf��@�,��\PL���5����KusEj�\��2K8]�Yq��ؤ�/]ѥl�mm�2���tf�,�R쩧b
��ꅇ#�����m�H��F�$�8�K�����Dm^�s������ܩ*�i�h=Q+�;NܻfM�9�)����KvA-���o!ѩ'.K���������/�&��1`8���Q��q����i�P�F�쬼ږ�f�v��6A÷!��u!����-0D�z����ǂd�����"bC^�6�Z���U�oY�婤�L�M�8�؞�����Vs^%e�u���02��h��)У�m��T�7�r�H�T�x�IL�s#��*�W���6��m�0�˙sn��`[��QV9��)�ӛ�R�7�e]](���3����"�xCܴ��*o^�]���܊z�F]6/3�p��շ�¥f�(iMm�)e��Hkq�K1KŅVa9V%F�������t���y�'��=�8�<[۩+2��E1�ʔn���n���:��X�٧XS)�	�;6�mD��<��ʽW�oY�0X��v�"̫!�v��g"�r��S&�4Л��j��2VY��Y�c��ޅS	4^�H$ Aj2�5�e��yyV�M�U��u��.���P�;�Vi0��u����fT��P�l:��U7]`�Y��6�7��G{��N,kj�jI��ȶ��o!�r���b�&ջ��o*�k�S.�D�R�٫[�l������m�M9�e�,�؆嗝Î����!�HV���`��{���L��$lKw�rWo,^�ٵ%�aƥ{��Ʀ����eʢc�C�K���2z�0&(��V�[�/�S���V�Yx�a�5��Sf�^9ErTA+)S���ҞH�-+�b�݌��A�j҆Դ3w]�4oj�m��^�OU�IKK^��-X�e�J�"��d��W[z��b�Z������/^Vԉc�5��<wzF����e�crL��vf� �X&m�.e�(��T�[0#��;�U��ְe���K,�4 �o.*d:��p%5���6�������˽$�>�lP�/E4f�e�Z��wBU�su%5-[.�7q��J*��'r�t$)4C��K�ۼX^9u��CVD�u(vk�ZT�1e�4V"����azW[%��\G��Ӣ6���<a���զ�u�hFm]�.]�e�Cv��9���w�tTk/C��CDU]_	ӡ��L�gZ�"�-	屳�݆�$��"�:��d*٣n�n
�i���+w�Pg"�P�^�DCy��ujM�Gy`�7cd�2ˢ��hͫG$�nK�d'��%^�͎�5�Yw��Jخ^ZV"�ĵ��j���Ŵ���jH�<7�Vj�6��6�!��6��yl6I�l�Q��$�dC/����6un1ke]c,m�aE���[N����2�-P�I��ZY>�2m۸ZR���e�E������<O��i��[��]�,�l0%�o��a�l^��	�sdo2����kb����l�����U^IF�E�(%e�ln��m=���j��I�Z,И7�CѲ�"ƥ���(�X�f�J��^	vj#��4[� �B�*B��%�ҳ����Z��/|b7���4d�Y���A��i�3]#[ڐ��(ݏX�A!PE�SHS�L
�d���^�B��bҍ���љbr�ix�j��T�u���b�6���Bu=��R2�F�Ƒ�[�n��̰�iؑ�`9%'bd��l�*;[�3�&�EM�������a	��F�8XͶ1��!6��tM"4㗋x2I��F���/eX.E�b��[�+U�)ť���4�ib��J�Y�r�Vfab����#َ�7C2]EOm���q'��J��#2�
Wj�v��f��=��Ȅ��z���ނ�V����fQȋ,T�7j�����ݴ�%s&�]6f9G4tCfE��v�Zxv�9�ܵ10DLb�w\����om�kbmٚ&���L�A{[��9��B��B�
B�k(d����L��N��;wj+���A�)HD��+lPu\{X���]�j��`�ׂ̙�������[�t��K�[��5͙��ٔ�ȱ��vD��f`���QOX�IA(�Ā�,�2 ��c۹�����6Ζ���{�n����
UD�fӚ0���0�Y�Y��`Zoq��ԁd������jf�@kVwf^hB����ZEZz��VE!�wNݪ�� �Q����7W�+�U���aܕ���њ�4�ĝL&T���9�9`�:�n��Ʋݺ�Q�����S`���2ya6q�Y�MWY�mY���)�Ñ�rB��jYn�	j��*��5���^�Ӵ}�i��\�;�aj�a}�}Ր�t�����]���vv�QuJR�iV)�"�LU�-ZP�Em�l�3p�}��M�O!��p�ε7Z��y��w2�S)����ݫ�˱_U���U�t����������4+'D������n%�d��op�z�X�ȱ(�rLP;�)�vM�i&���M&��5KR$�Iuj�Si=I�At�����3F_Ri%5m�
�iv���}�fg�_^l�VԜ����\R-i�V�ٹ0�L��+ͬ��b�P5ݛPgj[F� �ĳR�����-0N*J�a�{��uk\:�(�[�-e���gnc�"��v�����w�� �^�}%�-�z��c����/:��˚�)C�Z�ܷ��X^�Z�T��~��˱�"��W�G6�ak�Qv����r��&�R��k�WjZMh.-�[{���l�۫d����F.��,�ݼ�u-R�ԚM&�FՃ��V��:KڼGh�:�SuJ[&i+YՃ6�ή�Bm�������]���+B�8:�n��p��P�
��Kjl�i��v"GR8�&�J��̃�/��w�Լ��;�-m�bx��n֧�jН��Һ�b#��6�gC�a�k"�[�)ZTE%�GRz5�1���/V%B��7�w�!�q��$��">΃[}�1���[a4�ܧ7��;Z�ZF%iE��E�f�^�[xM�;v��������o
��O����\x���I���U�Xf�����>�^I'սF�iڸ&K^���X�U^C3�3u���N�[�uo4�Z��aX�($i����d�������S�НJ���⤨g{/fv����4q.����}��1M)�qe*K��A�6�E%X���l��X"˕rvgeZ9H�;3�6�wJ����5.����N�4��M�tB�-լӹjJ�34�ⵢ����S�&h��rw�%X���`�Z�v�i��Փoa���AT���{a=���V�����)5ڔ�.��½Vt�h.���P�qB;9��<#S�"�n☻��Yf]��[��u�R�*Nӭ�^���I'����DD��[iRt�,"�*J*�����-\W��|�/���#���.��{?@��,>������	����o�P�!�
���ѷ�M�}�-A*M��I$3)�Bt����39D��*ok���EKyU0��	�*�m���Y�@�-kE���K��<5�.T,���~bl7�Nk��Wgd���]V%,42**�ݣ&�F�
���ڧN�l*�EF[�F�]���{w!E"�!H�&�˷	L^ȥpC�&���,YOR���k��6����;Y[���z��՗�1�k�b��яP�T�oIU0�k}vs$N����CuJ�k���'�xv��{E��{�od�m� ��BQը�Zj�j�:;4`�ս��(�$�Z ���[��}{Z�q6�[��v�T��B�{�Qf����n�bX��.�;��We��X�_^=ĕ#��n���/B�aT��.�$K)�b�X3��P}�Iu�Z^s�*۬�wDq��$F�ƽ}������)�F$�񸑦)�6FQ�q�[��H�JK:�;���E͔�,�괶�}17���[h5Kz�}�4.'S���}���}�_c㨬�T��b�����uTǶD����R�����cN��0e)4,������tv�9�s��mC��HMju조�'���o[�'r��W���a�e��;R�K���uoz-T*��fa���Ӕux9�+rn�w.w5��FV�X�٠w5M�FádJqYQ��'	����o��\�,���͆���ǥ��0����ma�4e��fbwa�!E��'�AS[Z��q��';T��k��Q`Һ��liu�oI��^���Ԝ*].WIX�k-��z��]�
ur�yԎ�3�M���!WۃY�w�_iY׶wN��791��j��K;%��c�Y0B�5p�m��q��Q�:�0en��R�w[�T�8����2�-��V�	���ЉHи���m[9��F��[\:���VS�@�|ins�ntc�l�C�nս}{���k��N�t�[*���j�D�{15����.cZUb�,"��16Ĕ�n�.zh'{|b:7�����Tgh��
���]���1¡�}�tШ��6����gj]:���*�n�,-��K���t��u�]��g)à���K��F�X���a�*Q��KHͅޥ"4��:�Ld[e�b�a�u�4'��o,�.��74���@����Dw6��`��<����x�ҳ
's72�
^K(f��.�����2r�fY���PL�6V�i]��;��X��ASdQ�d��Q�ۙju�u!��˅ �Qv�L�o�%H�L�';o��{��\�ɍ���r0e���7뜻�L����.8.1꾷�J�c,N����%�/}`髋�r�L�M*_U��B89g:�e�f�=ߨ�W�0.�mD(�Ul�⃻�� �yo�y�aR���z��9���6o/^ 8soe�,�o`��P����L���s�Mԙ%������D��Z&��1վ��ѦA�;�+��HStc��������r	�Z����w���j�G��[�u{I�C=�s+^���v��55����x^ev��>ÒN�f��2�}��qSx�2[�4*w�oj�*2�����]xC�q�u����͂�p*��<\��0uG�[|�A�P�	��H]�9F�3��ڻ��o�JFH�˓5����՗&,��`���*�%�3/ I�3d:��i�2��Pm��ȸ�����.�B*�+}�h:��~��.oM��ח7/ ��ƪrD��5�pN�l�rv|�F1�v� �Vx�U1�5of!�J�y����ׅ������mhkk�\	��-V���Zkl�m� ��4 �y�z�-Nj'��cG��Ŕ�}�q�5wl��7V�阯r���|�l�ѕ���f�yM`N�{�9!�̗A�yb�������hY�;�S��$�<
�F ĈL26*7&�j�`�����j�2��gVN�����jo]��_w��Ƭ���Y�5r���e�z
Ő���aL:ڶ�b�wR�`�1�>��K�"�'U����4��ݛ��r�}�{��;-jN��s�N<{3�8p�Jû��8��]�C˔���3��s��X)�ǖ!�GJڂe���<1��%X�q�j��ɨ�9�������!�6fP�;��ݞ������J]{RLckjVq7�[��w���!��[��N���4��LYYgwS�n������Op�o�/���V�8؛P�p���쭆�oC8��Ki��7vv�X��=:����+���s-��sN�:��^!�5,|����]em�Ó��V2�f�V��:�3_t:�Mt�W%؜Ge�e�����n�	o�ͭn���ވتq�UՈm����̅�	1�f؂��k�G6�D�z��ctj�2�)#N�'�WI��T�E�Y�/�t�җ��L�8�f��a���8�B��r�w^��<���Nt�<c����������[������y}��L��Г���Y�V����B�1�n��ћŤKA����IXf.l-��T�tJM�}��F�g�f�z;}��F�y�9��䬋ܤ�K�7Ӕ���'m�g�%U����5�	���z����YO���s��"��4��E!��/2t��i�i7�v-��D!��$Mi�V�U}�t���BСy5�+7w�u��ܻ+0Iv�,Tm^F��s�sjo���ne�r�ч��y�nv���Y�z 15rW�|�oR�2n�䳝>�36���F1S
#A��ӯL��8��� +�ަ�PQ(��2kOn$� �Wۀ�P�F펮V��!B^�۽լ&�͠=x^o�2��zQ��̳�:�5۠V�T0V��YJ�S4�m6K%��t�f���A[[y�t��������\�e,A��"+�������m8[��"��']����7���	W7�g��r�=�����A��t2d���c���!�zM�G��Ԗ�K�o*��y%@sI:����vV̖D84ݣ6r�ﲍ��&Vs`��V&���[O-Z��:���˘V��zuwF[h`!�A<��Xz���-BeM�E��M"�D�«v,ֲыN?Y����[�An�C�36�0�#��m��ܻz�p���Z�����P�7W2[�R˷y������%���_gN�������셊�%�Xq%]�۰m��WNi��9����۸c9ܲ��{����NdI�gNȂ�$�Y�;T��cY��肚�̀]�r��H�7sX |�[�aQM2�,疇���9t���ज़5���oIK:�%�QX��N	mXz��L�ąs��YM�;٤��vk������t�4,�Zq;��T얯�5��I8�8W3S�mγ��W��zE]�rÚ�r�nv��H�j�M�^��:�#v+Nj
j!�Vx�+�*�ϸI�7}e�u�h�ssU�=�7fT��QMڠ�#2�v��Le����:5��;2�b��Ӆ��5����ݾ�����5
{��b�ۗ%`��.�jw�����X���m'�_y�g�U��&r��2$�ʷ�j���,ֈ�H�ZҒYK�U/U�d�Z\*=z�RY�1�:����a���l]jɗ�����rLKs�[����_;y�������J��^�J�m��Q֚1��s:��8�k�������ۮ��uLn�P\��F��W�H�6��/N�|,������^�����Ń����\a.�L���ƧnֽI�����z�Rcg٣gů���d�� ���X{�\[�����-m:pN.`WO�:[��+W,�L<�e�u)-���-	��)�&��-��Cjם��Q�ǯA���A��&ظ[B��]���;y4��(PүjP��^�X���Ѩv,���#��hC�]�����A�,0����h���η9�}z�p�e�g*�NX��6���9v�n\��֮.�D��i�����n-:��� �T펞'/�����<!
��'{�}�0X�	Å�\�_a��N�d��Xc*���nҮ��z�&0�#�N��cjV�u�E��e��ױЬ���Y�3{ Z���j�QV5᪫�ue�TV�%�H}5u�˛�SQ��+Q�x@H�-�aڈ�I(Ma ӹnccF��s�X��E���e�Ӣl�A�]F��-�Z�����yR�@`�M�Q�;b���;u bξ�,v��ѷ��6\\�ģ��Awzc�u��sh�I�J�ZFְ��]���*tf���Eu��8�'��ފ��x�k�n���8̚�V�Q^���"�=J�0�$s*
֎�TB����үiX��{OJ�P���;IR���QÝ՞w���n��l���q��\$��R�=�u���'`���;o:Eՙ�yhin1;`9��7^R�s����k��h�E��J���JX9�4ά����rz��8�4�خ�����=|��q�D�LYs�QB)��|���z^�#�]���b�۷awVA.� �J�͂���I���3�gz�m_AK��qtl5�U��7x3��UFkC���]J���.��(@�Ǹ��j���r�[��++��/�A&���f��q9��Zb��7f�̶��,����:��V�/���T��V�BW%�����]��҃\T�}��\5ט���Gu�\:��w%\�V��r��^7'N�pQ+�Y79ݵ�z;D4�o;�v����BnP��Fm�Z�4sap<����B/��G���}���t��������9
�DP�X��!��6�{\M�v�n�<V�g����ֽbt7t�!�w[��+a6fI����A����1e�')K��8��U����J�bŽht��"���h��:�sz�)0���r��eQ���[�6���i�qkr�����:]�fۗ����ܩ^.6�Њ��!tP��b�k$2�-��q�'9ntD��[R�8/T���u�b��U�<3�U��H���,��@lp���*��k�&�(��%��a��[�V1�-	5����n�VH|"9�:�nA&�=�S�,���V��ζn��YW�U�Y�5�җnS��y"��Su���k�-��q�9��wj{V�����5�^�o��޽�/st��Eu�0wQ.��G�1+��2���`y���;��*R7#tFT�a�T9�T@C��dN�˦�/�q���J,ъ��cNUs��)8{���w)*'	7�.8�+@�nD��cͭ���ol:w-�SS��R��L�S٬[�l�^�/1�R� Z �V��N��꾖�^Ǜ�;p&���ʔ��:�"ekU��	j���9%��ЂV**�]�b
�;X8�BY��8��d�j;mέ�Qv9��Z�ee�}�VI��$V�2���#���o�����,f(����䄭&�f�@�����9�b#�,�����*��f�Q��Y�KtYV^�ջ9�Ō]����W�N!&���_j�' �3�ޫ�4k����k)%Pa�qWߜV3�໇�R[!]ݚ�d (G[��_�/�N}ē?Xv��鵵G4Pvq�VLw4\�O���9�����:���*�-7'.�܇n�:��e���-��*��� [���vv��Ox<�wq��)Q�o��2/n[jK�*r oK��Cl��hA�i��ȫ�����5����k�+�b�$d���Y��b����٠�oqi&����82�in$ê�u�e����W^�$�pϺ���<w�G�ݡN�owo�h��o�zK����=C����ŝם���w��u���HL)�|7�{p����s8�2u����ll�b^ݭh�&��LP����L�cQ�:�6�Y;P$JT�6v�C��U˲���)ދWW�T�90m��g#E�-D��M,-0��Q��L*ZDMY�=�	�$��owGA,�󷐲���z��&�f�mniM��m��m��m�����l�L��b*��3F�ً�-fth��up#m�xG(�6�ѮpC�@�UP��"M�#9�	 �ac��+K���	EK��:FPC������)���][�K�u<{(pQ�4_ucP������@�c<�d�ݠk�#�#U��Ҵ�F�F�*�(�����[��-t��.ʋ���<��T4�ȊM�嘐��whpy;����=�H��c�i*�@e]hL�'�Ytv%L�4��*yF�����ؕ���Ҟ�[� ����H��>J���9P����H6#��1���~0Wǡ��혥H���s�(�am�O[�89�
�*�mq�:�a��]�9ʤY�Puܥ��,p�ST:�����R�쬳�G9����'�Z��!���澥-�ظ��+	��$wP�%�z�L @Q�$ :Ww�P.Т9��A�5�B=�9�8xF��i�9@j<�E�b�(#����mAE>�������~���� ?��@w������#�?���?�e��ۢ��ު��5ٕw[��
 �!I���
� �uҗTF����\���F@�F,נý�����U(�ZW��V�R�2�,��;x𹟘�wih��:�%e2�DAmc��W`<0V�2F^�/ ��u�Ww7%�ɦ�Qf�5�IE��՚G`��u&�[X��Z\2c��g���;��)% �t�:1��ն�H��擡�l�ik�FZ�x�����C+G`Ζ�*B#4k�0]�7%�B֎���W`��w���aww)�XaFx[,@mh�6�o)�B�Z٫ц���,�]oW\�`y(8�׎*�����͙%]�ie/I�[vI�1�F%����f+��\�x�QQ�:7[���}/(�or�Y��^�B]
}�����tD���7�WT9�c�팤$ö�wQ@�$]`�� �5�.��&�Z�MV���{����r�d9��Kk�m=PḼ�YW�9|���6l�cȯ�ik��*��6��r;�SkޖGc�#��W��[�u\WR�֯T�pl�]�a�QF�F�S;bN��ۨv�z�H�{v��W�љ2���[΁ScW2܌+p�c�����>U�*ȄQ�u�����ǎ>��㎜q�m�q��q�q�q��i�q�v�q�q�N8���\q�q�q�q���������q��q�8�8��1�q�qノ8�8��:q�q�q�qƜq��q�8�㎜q�q���8�8���q�qǎ1���K��� GB�n�܁��2]m,�Gn�.7e��Z�����U�Z�OiNG/"����!k��q�R�c�ޮٷ!Ӯ����&��ѣ{��˨�.����e��H�-�Zgwv�z��BѼZ\.��rJ�U�M����5Ύ����^�j���ӽ���3z�uo��iMK�gK[����%*���r�c<��j�=�d�<9fDZ.�
Ԡm��01X��P�%��. H��aC�V8A�l�*N����쥎�3w�bwCr�6UH�F�0˳��w�S�f؋[���.��W��Y�	&��v�#�v컕+z����^���UFDüS�*�j�D� �����B�i��ᇦ��="3�֟��J���]yyk3K�Vt���'M�A�u�U$:��I;R��4վ�`D���gS��j\��u$�ue�6�\���J#V�H��wf��QL3EX;���J�W�����̄�"{-i jz��'�W%����r�`�N,��hJ�b\{"p�Y#�"�b��%XHn�9��cj�v/z���^��#c�o-�An�(R�]�:��0uk�aJ`�Z�f�P�3����u��6��o�qێ4�8�8��q�q�\q�N8�8��8ێ8�q�}q�8�8�<q�q�q۱������v�8�8��8�n8�6�8��1�q�q��8㏎8㍸�8��8�n8�6�8��8�q�}q�8�8�v0o*R��P�KOl �`�b*;z��j����Ȯ"ul�W��!l�Gw�ќ�R�n��3�]+2��E:�9�x[zmd;�%�;q�M���ۣ�i�+�W��E�eӱ�� �3�^��jq`�Բ+ۨ�2uӮ�K�����F[�{���{�S�#��9�W���^���M���X����[n�5ғnm�x���wou#-��Vբ����J ۃ8��-�l�g�m[]�3)���]5��.�b���x8<�+UY�6�2�!l�.;�]���ݦ�*x��Vc���ٵK���Z��{��f��1`��hs�{ީ����3.o$� �X�GJ/�V�V6�c�1�8�ʅ��]�`"�D��,��֫�W"zn와W�4������̠��J��s�`a�X�������s�g)݊%���
/it!`sjW�N��M�h����\3;�_%��A/�Bu
�}�(^2���/.�ǫ�'!U�Fa�/{�X�B�nێn���W���Y������rK���lA�ڻ�łM�X3b�(nН�U�f��x*Z�r�C��8����Ϫ��j�#*�M4u�҇xp��q^�RÏL�rb�Hn��ʶ(�iKA�enѣ�L��u_V�*��F�*6�^&z�Ԩ���L$׮:i��^8㶜q�qێ8��8�8���8�8��q�q��q��q�8�8��8�>8�n�����8��q�q�n8ӎ8�>8�6�4�8�;pq�q�v�8�8�;qƜq�q��qӎ8�>8�6�8��q�C~B�^���=ti�Ht�dr�����l�w�����I�)�Vj��k��b�� �du��Ge�!��ӰC�VC�u&]>��ҕ�ԟiR��yu�1vhT�Z��ٍn�bar�qXY���@.��Y���lˬ�%I��(V��V{V�ӕ��,��3I�����eTB�ل�V�V�+��򾵕��&7��Fi���k���l�f�����E���hP�v"Z�8S���l��,e�鹸]eR�(����u��' ��x6n�]��&�ޛE�4�㓯���+��"/�[M�ah�/�e	�cPh���R���yj��P��M��0]��pܭ��;��r�1cf�Fi�K��|��D4�]}]r��N��F#��T:��$���/3�n�	׏��ؠ��%Q$M{��<�r��YK_Jø�W�y��9je�[i�,d�R����r͕\=p�[g-�*\:���[���ͳ���fb뱡J����Y�U�æ�Y���0���{5q���)�]��M��f-�w2J#����������-�K�C� Ѻ���{U5���t�IfG�s&X�:zP��gTSX�m�$ЗA]@���w<nU�]��`.���\�����ӱ;[��KF�kꌍ=���n�z�{��Vh�����(-��W�2��a�A�ޚ��B=Q��)��Y��-G�	d��.#V��ѡV�Ԫg�y����Dt�۶�8��qƜq�q�n8�q�q�Oq�\q�pq�q�\q�N8�8��8��q�q۷nݻt�ێ8��1�q�qノ8�8�i�q��q�|q�q�q��8�8�8ノ8�8�c�8�8�i�q�}q�qsu+[�C�
�L����h���;F�������
����}ؙV��]q�I�Օ1��1�k�ޔ�(\��c��a3�����:3�Q�V�v�S{[��2�`���Ӄ3V{��;|�ꔔ&��\�Ʌz����lt�4�,*b��!�ܔ�,b]���:.��ҩ"RIK��:C�f��!v�!J���E�����}�{[[@���k����=F�f���*+GoK�>wi�����;����VR5`Ci�V� q�E�������� ȹP-�ff�i����"���g�_PO�C��Arӫt��USHJ�t������i��V�
�!�F���b'�����Gřk�\���V�f�vX�d���Wq��#�[�W���9m��X����ڷ�l�)���r��k���^9|n�L{ӷC��:K�oZ�+��n�o��MXi*KE���o�xa�9kB�� ·��8���%�p�cپL��)\���t,,湹�u�[ܥ�2Q]���f��Gq!�����1���J��^�X�Vn�ԻX��)��#j��Ӻ��؆uLm�uV�z��Xl.���%��v�)/�(vGZ��t\@y�л۾�yd�S)7SP.�^7/�@�ia<*!��E�b ��ٯ�k{�;��NX����Y���R�h��r���i�6���V��m{q���mՋNΧW]�:��村f��UUn�)�'�Գ6���3a��qX4�R)�Db^����b�!-u#L1`�3 �3���Cb���2���[c-�Vu�bZT��N�V�mX�PU]Ց,i�vӏ��=�_��Pzm��z�󂢞�vE[yZ<�w��T[����a���7�W`�k0w��ǝb�kޏ�;�7z�5)*�Ӕ��� �o�x6��{&�x3w���L;�kWׅ��VU87�0�VČ����( zB��I�z��խ��OJ���_^���:���;����v�ڣ�zW[�:���cU�tʨ0XR�;l_DM���Q�欕S�t����;���xK=X�V�l��@D�
f͹�/au��c�ʲC!�x�=ݭ⫳7p�ڒ)3��:,J����Hz��弽S�y}���2������Bʓ��r�l�#�8=���iCu�t9�W���JYF���fHDLͪ�̬��_Ұ��b��y7�f����]1O-��ci��.KDܶsa����H4�F����4oX��1��Z�a �͢B�u�a:��yy���	M�q$M�aN1�l�Ս�^�wg�zݝ�t�w�����;�X�3EE���(��nm�A�x�b���YƦv�����8Ж4
�P��;�W@��=t��K!^y>����Je���qbu�|�tXT7Ҳ�%�-��p�Y��I]n�Y7m����EC��D��Fp�0�J�F�* {�T�s �tG���\���j���5��{y�y�t",��c��介{��*%F�ԋ��Z,W�%핪n+�@$O��f�Q�Y9���+��b{�"/8��7I,�ww.C�A�w�l������3��!λv��m��:�>�D�W#R��, �n�}��7�ov�goL��LgI���4e�N�����+�	m��+�.Э���j,9���3�)��Cr�P˗Jliɂ�U���Nڔ�Ѷ�.��q���U��J���'B��f�����Q|v�_KKjJa�J5���I�(�C8��8����8oM	�k�ᯖ�8���]��d��-����%�a�$.46�;������,���b��GK�R,٩��g�;�ȖbSj�d��N�C����Od�n�|zɉ_5�Vz� �Uً
Y�͙�57C��wٙ|�۽�Wٗ��ӆsر3��sc��6Ni�j�F�%f��0Х��ɚfV�&��Cvk� *q�5�zy�v��ɳx�����t��w�%��ZSo��To���e]CZ^�U8-�P�T�[da���� c/kT� �hU�mѡ����y���Uvi�H}t3!�M��uq3i[�rd����`�S8\���W��1�{#]:���!n��m���GL�息�о��{��i��R�B�hf!p7�mL��9�����9ו��4�o8hVn��|�W���.|�s���U:��"��v`ɒa�KsM�Gr�G�b#z#Y�r)�Hz9ζ��� r��<Ó�t���ޡ�}�f%A^^#���I���oZy��k��Ί�G��j�sj1]F�8Mڛ�IRG��}:�=;��Am �2�T+�]v�@��j�5��1P�aup�h�7���v�r�ֈ����h�Aw�
װFJ�$੽h���E�9*v`���jg+�h�*X���}r�[�r�Mʎev��9]p�16Fqҩ݇G�lSYa�Z��`�[��P�}-���td�XI�c`�Fu�wbM4����-G69���g�U�9Bū'1n���ڣ��8z$ݺ]$ޛ����ƌLcn�2����h�޶���-�,�Q�����ct2	�Hn�~}���Ҷ�M=���*�x�ZT܌Q`�{ݔO�§)�gA�%z�v2����wV�(�k1���&�)Q!�k�c�$Jx��+z��ݬ�����*t���c����Y5�Ѡt}� ����z.Z}�6W>�FR�E-�d��M��:�T\1���4���בK{D�����g�-���zxNr�HC{i^�"�� k���t��1O��Ch�u�����$�0"m2��e�'�����Y��Q4n���Yy/_�.�0�h]�rB1E:��퇽���m�a�]2��t�z��K"t$��ܐ�j�L��k�hRp��r�y�7&F�Yl��^	x֠kIѹL3 �ںZ,D�O)8.�����G0Z܀�v'��.�ք]Υ��@4�������x�I]�v��t��%�dTp;�%,�gn3��f�X�3�"�Pz��^�+U�͌]��Ph��MwH�p��&;5��5e�u�|k*�/���`�U�����Y��Y�F�uSoN����A�OtSd����7�`�4�D��k2����ؼ��������M[Քv]�\�779ظۮ�cW�=��q���I�e�S�e^e��P�L���n���ޣP��H��p�݉.�<x�J�ɗ6��,�ř�Ʊ8�A�}��N�1�ý˥�Z'v�\6+�;��7���Al�u��d�{@�ZZ�(�f[z�m=ݰ6�ULi��wV�QK�vf,�
�I�T��-����Z�4�#�[�8�+��F:eQ}}�UεZ�r;Yl[��xwi`*n��YWR�Qb��MW��s���io.���/pBR��ڋ�����i�]�T#��Y\ޅ@�w�,׊�g�`�\���8��ns=�Ӏ�ԕ_����ͬ��-9,��W�]�	��*s��3w���H1�*f����fY�[�_'h^��-!(Ȼ�
WoDi�n��jn^��0l���b��q�Çz���}������2�K�N�>��z�q�v����0DT����O{���������%^��k�����B��L���E\\��BrF���a<hT5�]�wt_e��x'����t��e�\�3���e�j�cgf-{J�G�I�d�Ů��p,uX,!��;}�X9�qv�f�7����-������|���Ή�oK#ר��y�S9]�����vW	ޜ����ݡ�{���S��X�W�+.ش']����5�ԥMRQ�Y�w�2�=��5�
�<a�WXJ��u�xC����mS��sD��N>�Ć�p��5yF�㕚@ٻ-�|4��R��gU����{d��@�֓[t��Q}�Y��H)<z��b�oc7 ��M�4f�+pZ(�*�P��J�J�6�;��Le�����	���p��j���� ���+��~?������������~�X�����Q�jFۍ�KaP�����P��H!i�dn�AD�q��T��)@�*E,��%*�hB�@�p7'���@�G���13�)¸�
�U8�&��$|��#��E�fX(¡�!�� B)��:9uI\�	�lR@cm�H)8��%l�ڄ$�f7�]58�eB`��$F�ađD��0�F��8Z�����^��Ӳ��x�����yz��>���>�*���-�%�;]bX�^���uD=s�����.�`��"��h+��$�v����bĝgOIr��dK�6�|�"��.l$kV��V�ι���
��ʱ`.pճf�u��[p�u���*��Ʋ�U^�0�H5����&�6��m���{rm�Ȧ�}����H�E�Fa�+$�m�����������X����^���V�n)�%�mjp-�rHk%��!�����	7�'7�)����Vfr�����ɛ׹�ng_/g��t���%iW[�k�^H&�U���y���6;���Gk��
�k0l|ʃ/�5FL�{�Ԣ�r�@ӝ�sV}or��ozX���^�w�jk��qޫ떨�8���e�؊i�a��Rs0��;���9��F( ����ӂ�ooed{%-,36�Ut�jf%��{(@�-J�Y�7:^����	3���V+{7�tf��oH�
�^�<088����zp�PS�A�9avTJ�l�R����(=�nظ�Đ\'S�0E�%g{�k(���R+�b��6"��쏝\��hP��v��7ݽח}yg�����YW�Gg��}�;j�Sg'���)�;�/5fV#�b�E4�O�L�6�Aq"pꦔd�BVH ��"Ce��M�hƠqē2p�BjH�m- �H����ƘDP4�@�Ը�*N9
7�$r�1�)6�㉲��IFNZp8���$��'(�P�J0�QHIM� ��<(J\q�L�eDۈ�d��M��%0���cE�\pERR$T��S���.((�-$H�x�N��T�d��4�4QG�n"[!4Ck�!*B�-� ��2
0�"���yE�ĒH�qqF�&`m0�(�p2�tjPa�P�B�@��l�ȡ$�S�B�mBCL"	�4���d� �H�AגTVq$̜'P�8�$6Yu�h�%(�@�ds��d��a���J(ɶ��i�
�A�9E��&gA�A �S��O}��u�!bf"����Ҙ���
m��o�;v�۷o�8� �nАł�#_n���)(�i#M�q�nݻv�۷�1��B#!%�u�хLe�݁`��N����D��@�ׯ^�v�۷nݻq�rU^��W��E<gp���\����ۜD�ܱw��T���wwl�s��$��:Y������v�Eκ뻹t��DJ�P	T�޾=z��nݻv�Ǭq�22H�IP�#Ci+��[T����u�ȱ�v�E�p����78���y��6�ή\�ǋ�w[x�Σ���];g�V��א���K�m�2�qܜj��K�"Ի��W<뢏�y�q.j��s�w�ߝi�������:��+��l���r���bW];w��'%n�uw>�O�0��m	�6��r�$Q�M*�ED%RP�!�5�7��ڢj����y��ܚwtD|��Q�wk���nT�M�/�}|�ވE��B"�\#חk���n�#Pz}/`Ɠ^-������&��qG�^�K��h(�$y�3�(TQ"APlN�H���X)��)4l��tY<�����!�%\�*�E;wJ��=��St
+n�������*������΍��Y�9���/n,�%�_e]�X��`2�5!e��T�M���,"� �F6ю!���C-��&q6���'P��D�Ah��a�J&�#���&�(�k�8�0m��9���W�]��tt��!\rI	!ڨ.��_�wyN�nk��kewl&�/�`�ɓ�9!��E�a�%�1�?����vg.���/�����^MۊZ�Ɩo>��\��'�ss�+��b�F���
��Ϙ�|0�eGv�Y)��f������$P��d�,<zg�hC��ɃFR$u;z���'�&!�[Ͼ�+]�ܝ3�q�;�8}©ꓹ-L��T�q�4��J���1M-Xk]�b��t�7\^Nėu.�\X���R�Mvm'l����7�yϻ~m��vi��NB09�/�eY�]�}�63�Z��=؟9`g6�#�t�ucs0�ϙ�R�T]�E�Eo��6*��^}$���w7����[g�­�p���]�,��h-�^|$n\��� \#ۍֹk,s����29����a�qɸ��3����}��p�}W�N�.�$E\L��UHqM;7Lr��R�Pذ�/vl��X���^�ՒE� e��� �M��e�r���#D�L��NqWN$VԽ��е
��^��Z#讚�0Zw�B�i�G: W���|6���vP�h�Pc��t;V�9�rM)C���67=�v�w���
�%XT�C��a��v��>�K�;�C�-���v��B��&��d��.���n��e,��O	�+Z嵗%�Y��v>��ݪ|`^[�^�m�}L��΂��؝���x
�Q�m��w����C�i��2�8z}���]��4�Y�`�;0��c���Ƕ�{���O}�f�侁���1��}�cz���z(ݻ�Ԝ,t�����꺉}�|@��Mq���,86�{#�qnd���9��6�=}���q��͞��bE<~��פUmI7q�I�N/�h�A͒cI$�mXt�F��b_��;-�N�iTq���d:�ﷴC��۱���ֱ�����Q٠������p��7����9<ꕆfq��B��uq݇���f9��u���b��'��B��\I�Eޮ������]� H�B�ssF��7O��Ӫ�O�
G��Oq��ŵ�����h{�V_��:�'���f�m髩�ݍ�Y?�� |ѝ7��/F�����2� ���鿋�]З&ټ۞�ؙ%�:]�_J�B���&xإla��3W9��ua�Qr�vTd�U��O8��ȋ��ڃ��䊷�Tz���5�3�Ԥw^&�t�z��rۮ\v�ۮ�䫲`ddN�'�d���qE��UCS1E�v]٧��p��F�wК�����g~�I���r�'y�U	m��l��S�i!��`Cﷺ���p*�'�j�X�D�SC��R*����>���{�6qgYTӄ[_B�-���Ű�8�zf��݋6KC���a3¯�����0'7Y]ϸ��G�]�q�(.6�\1�{Fƅ'� #T��D���t{K�"V�x�}_G3���ɼ�f��F�����Ly�.���2��/M�ok0�.)"_:���cS	pm��1�j#Fd*�ٛP�U�#�A�Z;�Jl6�jwա]ݱ�>0R��V�.Xi��-oB���E��Lng�\�a_t�kfW�e��2:�:�C�n�����Ӫ�A�n�/|Ry���l�[YW.�" ��X)��ݦ�%�K����Y��e��[�ǭO:0��Y_T\oc������:[1J��1)vh�ݎEU������"NP;��F��G;7��p���E�!w�:{��j�@b9��U�p���Sn�������!EP���`�qF�tnM��B�0�d�^��`N���}��'��4L&g{1�F��f/�ne��>���G�]y�ć��EX�D�.)[��j�D���~᛫��u��3]1!lh����Bx��|�lm�j�G�T�&�����9.�ƻ+�?@cM�T�N�v���l���K�����Q�������"^GR,櫄��Gb.�+3`5���$ߎcϾnxq�OVJ�Nq��E�WG�
��6Ӂj���VjҸ��W�)��U��/��l��j������bt.�B��7A��L[t��b����\�!����P����ǟ"Q#�c;}�6�D|n�RN꺛�`{8��we\]�yхʖ��^�o^W$�d}�(*Q�E7Wj�o9�(tbQ��a�Yfͣ�H�M�ǂwzɻ���g���D��@N��5e��s���-��i�?MC��/�-�]�
�D��k�[���:O`џd\��o�K��M1O-2o�X��`�3s,�G5�6�;��//!��l�Xӥ���mn��7dm���@��#b�2�pA9��+�`��{EE���7�^��c�ݏ{��N4�p�#�	��;5��蔦q�u�'��D�be��eF�;�v��}\�Y��0NյrM �8�%_PS��[ac��|����ۍaZ5ݏ�qF��}Yh����W�I�G���;��v���1K�5��譸սyR��ut9r�fxn���[�����P����ԑ�ˤ��{�3f��z�{�����T��6��歬w �\����u���C���՛���!��cE)��9w�q��Q��}�t�����m�:7�i�5<�+����ng�>ڑ�����#��U���%�������z�>��P�w���v�XKt�r�f�����,�^�Enc6���V1�����؞�>m�NU�:�~S4"�A�x�[޲ur���\'GT�;���n�O���ߋ�|ݭT��y����}+�X�vd���+>�s=�R6
�8;���}m�M�m�ꕘ7C(^N��ྎ
G���T�)j��z/<���#�' +���U;{+���X�B� ��KW����b-�P�8lv^$��5�����$E,�`�ن����7f�a���8]�y�S�; �%�p�ɸ��Ʀ��"~��c
o��fknI`�[�K�b�-f���W��������f��j,���%��vTGj�7�n�0л�+������]�=�W��	;'c_�7��k�vq>̆�/N|�8v6~�<�f�v�'8�EC�;qڶ�����S8a\��m��n}�*��h).hφ����3�p� j/*in� ;`]�� ����z���q�U���Ԥ�f2�5���7nN�-m�%��Kz.��֕�	΅�м�u��I(�;"��������t���E�_G*��B�W����q������d5���{���a��)fg�'�ab��a��aL��u�2��Stzj$Pg�����@u�j0̈�7�y����~oH��Tc� t��j�=��.o@�!��0
��ks��������#�[�ݣ����X�.>�ֻ��x�S������3V&i|�a����)�_�V\V�uf� ��+��ƍt����}����5*}j6�$�OBg�ң���:�s��t�8�B3-ܦmL��`T��bB&�r���U��@+5Y�V�ȅ�����m�����vO���s�ȑ�0i��C�ttGE�ډ�N붭�J#��5t��,�}.%�ۓ�=�B��!�k�c=٤Ov�t��NN����ma�*)�-��;x"e�O�����gF'[����27��3f�G�p!��O�-P�����c��5X�����Cs���z�e���h�S�лN��^(Rcbo�dl
��虩j��C�1⛩h�y���\FP��x[�e�Y�{oX�$��_`j���FYx��lTq
DK��v��m[eS��M����`�׀�|R�(�Ӱz�$�&��WW}M�<o-V����#�E��p^(�jGv.��q57�"ig|鑱O�00�fd�p�G**%���MY�.�2��'���Xv��Wg�Q$@ӆ�YC��;F�}9���L��ݙc�j�+t����w�_-�ʹhtD����z&n'u]p��s�ŧ
��?n؉�(G�c�-@-��&�2�}�9J�q�4V�'�픮���3���s�A�	�I2533m��{�|�����9���s�q�ߨns�e¨���>�6��gI�6�U��]��bِ��꟣.p�������a��h�ݬ�VHGIy�&�qRB�v��݅��T�f�@;<6x�S�qҚ�����>��4�k�Z��p��Cz8T�`ؘ��[�)Zg]�u�9b��8VF���D;���e)�g�x����\��v�+n����'���ʴb�b��e�q�j�@xq��;��N9�ʱ�cֶ������e+�y2������>�H=3Zڝ�;z�v���j��A*I�6跸�l���Gi͌�M�ϛ�u9�",-�� ȁƄ�\�sʔT��]-m>�����ŝ�|�9��]ޟD;� ���7l(����\�TC�Ǳ�\J�Z_	��x@����Z߳L�>33Һ�S���Y���k!o;�Gc��V���+�@[VHyB�}�5_,��S�?-�
�h9��yWf6�:un�H��h!��RX��{��/m����ɣ�N;�t�~}����	����1���MvX��u� ��s;Qq�1��|��7��[�`<�}�G���s��»O�G��"*��{0�.ͺ�lԣwi��|;���b�o�*ɣQ`A`�nn26�7?D!t�����3QT�M������T���1�4e\��p�N��Z]�/#�1B��t;�D඼�j�i2l�s��&I����Ƭ����0nuZЫr�*�������)���}��R̔���஛�ѓz�B�Q�o�\��M[sn)�t=�*�1�*}�D���wI��SS�{	a
���5�2}��y�,k��5u��HK�%��/h]��K�[�R��=�wsQ��t�Kt;>b��z��t����!l�<iju������Z_l��d��4�/�;�2��Y�8#����Y��Ȭ=ܡ�[ȩ�m>�q��V;$�`6�Z��z@�[��S���4.[�f�LD�9yfV�+�z�,p��o���ݍ暶D-�c����n���	�O:���&�_�Epݥx�+Sa<��w�ʾ�`��{@��ü+%��W�@{S�0�L��MPĞb|��_mrϲ�����o��Ǐ��ԧ��p�DO������ݪ�IXw��e��7'ȹ6ywF}!.�uu���g�F���=�w�K���ٯ��lу�A��=��y�m3Ým��_5��B"�!D�9��uء��#)l8�ٿ'���C=�;�QPr�R������I�Vϝ� �}N������s�r����B�u�&-V��s뎡u;f��aE��T��S��\	QPv��A���F˳o*6�75S&�n(b�ˢ+�_L�cH�[�wd�=��b�4*�ٔ�3ز
4@4�Λ;e�G`gg!�,ٺ�xK�1̝������ԖtR�P/Wa$����2E�{N{�1��0I��{�z�W i�E-st���twir'5��|�Q�8���Zb�`](n���ث)������\�TN�9a�^����ݠ�l�񋩂ծ�[�"�7*[	rm�F*Ŭ�h�[�۹�rIݵ1j'��"�����m#·G���T�7�3k)U���BY#U ӢBL���K�V{!f`�<����]��ܖ��6��O���M���$ѹw٥w2p^&�{ Ot�t��OK{��p��#2mʡ�&訋L���l����E�y�nӻrdH����eإ&�v����]h�EX}|9�7���q��o,tyuN@��n��b�w�b�ν;@;�K�hD�=���ٶ���7-q�9e"�+N5102�i�+�.���KUض������].�-m�}��̼S�{y;�Y�;��� ���z����["��C��z����?���u���+pѵtl@W/u��cs�J����3c�1:`F��P�k(��w��mc^����Nr�f�X��;n�P�6��O��%WT7�]j�l���]
B��=h����0��/�H�'F�E����_q��}���?a��,��{�g����\���}M]Dzm�wp䗁�'sm:s���5���׈_�C�Ɉ�,��{�b3���_se��{�d�!F�ѭ˽��N�v^�;�u ��\��W�A:�Ӕ��`H9.1�ْ��av����'����!�+a1��F�b���"fK:��H�pnaa3/��ˢPǰ�ֆ��_Em�ÑqH�c9*8ydZ5���X쌋;|.�[j�uWc9�kY�nj\�������.�v�X7;h��q!��V`ή3j�c�he�����QBye�`��r��oh�}[DY��f38��7m�ߪ�t��^�Vu�tp�uG��՗2�ei��)ܷ\�#��ܓ.�ܡ����i=�.���.6x$bͅW0��˽��m�8�c��V;Q5v�����:�Q�?k�H�:�����poJÊ������eLc�Hm��@�R�p�^A���pΤ\�s�$�c��e��y5�Ͱ�o,���Y2T�U��	���Qb�I�r]��N��ن���N�;.�:f����2�TG:�*�pֻ��l��m��zK%)����V�ͺj��z���oV���p��_~߻��]+�a$Ţ<U����t�������Sz�;Ǐ^�v�۷n�x���:FE�I	���/�q<n?hߝ�.���uP���!G�O�^��۷nݻv�X�;$�RvT�#9�x����A����s"��B�v�<�$�P#�o��޽x�۷nݻz�qp��@�*� Ο~w���=j��B�zk�l�5UL����F�=z��׏<v�۷���u��ں���d��`(ސ\ۺ��Wl)
 �׎b""�=����b��1����W8j#b�k h�+��ӷ����IF��]݊79��Psnk��ܻ�p����n�F�r�u���Ք���nU�p1�k�U�_x��UWb�b�c�Ѩڑ ��e�����!tx�w!;*�I�gZ��Rv�ُ)C��$ j1S�ai0L͊���}`�����w����ÙV�ruj��vt��E���e���p ��;!?N�T9��'<�j�r���.���� =��0h�#�|~���z�G�*�g���{냂�̌�Ν�Xr�MJ��G�>}�;g38@ X	��eo,�-���ń����1�Q��TSKAjT;�M��sN�����]V�/{�s$:��l+>'��ഘ���,/|��۲*���h\�c@�"SZ��Ƈ;��fRʫ��y�{�9>��{CS*Ȓ�I�o
�:g��1U��@����,0!��U����c4+F����)�B {5ϭ�q���@e���W(ׅ'�{l�t�M=���`&r���������=  ��ݰ87�S����2/��=4\�JE2ԥ57GG��fz.]h�qWuyen��xZkJ��ÜA�S!�>k�p`\S�3�� ��t�kRT[Ø��{0�lB=|4b�������0a=�<��c�1�о;q�6a��+}���>z�bp/y�AfL�,��n�Y���B��co cr�~�c����6x(xy�G���m3�O�t���)�!�P����$^+�d�g[�jW��,��&Z2�(R�T\�`�Rr�ħ�L�ݵ���3��8���L|6>
�	��wwB���QF$�N]]G����x�m�S:U0��V��O)�L�����r��fa^��V����n�ݺ�۷aWf��T����.�����/��`��|w��`j��c˘F���o�ǿ]Q+P
����9+���<0���9nts^1�'�X;�-&��:�|2����&@� Ha}JrELl��Z��G6�Vխ��~��G;��b�H��
S�����7߻9U��@�喅�֮X(�;��Hdgm�/����C���s� �ͤR�\�22}U{|���`LO��#�F8���fz:0L�0ޭ;9ܬ��6ogp/���Z��ȉ��$���	��d� ��Nu
`	/\aۘ� 7����T���+���/�h���C�X�A������GG�q9����eexN������ۧ궧u�&��pC���p��A��@K��ր�qg����6p����՞;>�bS� ��睳+�X	m�����_m��ԑ�忠:E���Y����N��0|�����`��I��0v����޵����[6ѝ=����0�z���4xbs���mM��W�aP6��=�f3�I^�ޏpp}+z�]�?��$^�4�C i�ݰ���^�P��� ��w�a�����������i����9�y!$�X���Y$Y�ɮ�ع�����ܱ���A���`�a�u��2��Be��e}W��7�"OT6g�+�j�_<��k��e޼o�����d�i�.���8�Yk�p�^�#�@(ۍ��[˞_OZcL��5AL��@<�^����;��[��Rr�����r�[�| 촉`|g�����&AT#�PC��f7�ޫ�x�Ť�|�,S7���Ǵl���ƨ�]O=�����^��h46q��c�)�8C�e5�pi�^�
��O�&X�1o!�;z��r�(oK	��]�s��  ��k��ׅ�zw�p!������y� t��yv�GT����ސ������ڇ�Ϫ�fq;���ڃγ�
nN��C��oT�m��}T� u>%E�./�<��pr���Ն�uQ7�nނ�j�vc"�l�xJ��xj�r.S�=��z���������$< <wyuم��I�olϗ�s��P^ Ch.���ܰ3��� Zqw�*�
�>��VW��
���Q�T��	��;^/��Nm^����8��� ��!�Gh
�0��@���x��=�*	p-�Ts_��U�x#�(��}�U��L��hp+"��|H����ᜩ���D���O�e�T:��X�8����"�X뚺8��/�,�
Bj��?N�%h\��мx
[j�FOǞ2�6��E�͈ݬ��n��8��	s.����^��M�����]����L<��.�=f�+o�ޫ�.ߜ��me�1���kЛ��TT�sCML��,$���E�e��k
*��	�+p
׸��������F� ����&�+(��3�2s��vL�+��D^���m���Π�f>�r�v��ٕ��+�+���v$#������B�iI$E�g����{>{��C��Ű#2F&
?����r���O0㖡�P$���<����q�U$����W��C{�Խ��p-��u����\�mD^k|�LC�:
n ��ͼ~)ߗ3k�m��c�xp�
��P[�����"�}��(�~|�1�NG����"p�1�঺&��-����>�� Z�W�:(��!e��~ F��@Y��c���{��Se���U�B����:�P�zw`ݯ��,��=����.��sf��v��;3���t�����>Z玓�-!K��0�pF_sr�@xYr�-Y��>>~���v���M!�~@U�J,�@'E��I�[���0V�1h��U�K>��g��8X�E ���I4�	��n�b��@�%)����O��> @���Bŏ"�̞��}���{�y]`��
`(1J=lُIoCo<�L9uJo\�,mO��7�m�������Hw���KL�e}5���p$u�b��;���sd�߅+8\Z�0�-�b���p* �pa��8��K�ꮗv����9J�i��%�|!��C҈�돤i��
⧡е kG�׊�`�rkT��8��cޗ��V�W��Q;�w,�*�ު��2l]1����1ؙf\+
�E6��R�ї�����z7�nznkUv"�m�J����24�xfv,r��Q�P�us��8��0_	�V7Cd�7�ޮʻ�,���1��I������B�BX�>w���|���d�T���i��:�A�P�p���)��9���Q�cO<�w���pp��UHV��R�5���;]`���;��Hq��o��Fj���.�+��su�<q���1�#_�����K�{i��S=y�@��nY���Ƽ s���q�v�����ц�� [�މ��{��X^��`��0�����!���6뽮wB�+�X`"�4�7�J\3n&Guk$8�>����q���[��[c{P��}V�ӻ�ţ��}� ��A��8���3���}��3�)7}�i���g@F�-���5��mN4��ܘ�x+�hVoH	��V��󰼺���F�VXx�MȎ9(x�<�Qt���%z�����|V��돀>������v9�Y��8 ���Q��� 7^XS 7U�o�,N����t�jp@�,��C�ʞ1���.U�Y���۳Mβx}��?wq��4�o��]���Zp �]���/�x\%��@"��
����@b�>���NZˉG���O�ӎ\dߜ
��8��C.~(�2�F�|���>6���[���ѕz��ft����|��)M0Y�ggq��="����Ы*�"L	U�5d{g6=#;��o;gR
i�U�N&��w�'Dd����Q��鋫�rm����ש�!�U���M�$�9��VY���%��������%���֒BE��Y�j�]�tV-cTU�jך�^����������~������b LK�<M��[�2X
e���y�vF7��ұ�V�\�]���� ����i�dH��)���#r:H�I8�|�)��),9���mn�a�aw>���Α�{)� ���G��A+��|'�Z�;� O�[ŨN�voc�C�p)?+�;1Y�����#{��x :��[0��^�#k��.�]�<<���è[L��M	�꾟&&z����^hQ�������}���W�%��I ��k��iǱ������G�k�;�0z�X��p^��`
����M�­t�xy~�Ϫ>�v��A_���w���!s.�ό(Ei��_}��D��7��r�X�c;%�!Ҏ2}5��W�q�#�bf =�Yr"Ix:�ޭ.�6���W����L�	�,u׮�����"�R-��Y�6�&�������nI�ʫx��ouR�c�����C�\p�� o��5�>C�_dc�=�6>{{[�-�~.�0�d[�D���V�9�:��"��{g���C`�渘)�C�Zs���5+�<����􀏨�g<@N�~�w��uֈ�]y��42U���$�y+�=u�O�Ϧi�7Q��X�S��8>L���9+�o�XI��U�x
r�Kw�>��t/��X���;c��k�W�t>�Cr�cv��oQ�?P���hN�k �΍k_@�O�SM(SM! 4�HH
"Ȅ��'y5�o�M�\�A�SKJ�yt��j!pP��*�"�cW����A�o|��}�˴�ƴ�:����|Q��O�^ac�+������4F���C8`�� �{Yڭ�\eנ�,���ԑ��/&�W���K�X0"ä�Ց��J,�s)����k�7�΃�?���i�:Om��ɩd	b���zU|��K�����N%4z�v��G�����G$<��hy�#�����|ki���}��v�b�	�Ҩ���trV���h`5��3^�͸:���>�Nz��x���A9k�p�޾�"�ָ-ט��Ķ4��M���	�FA�mRv<�]Օ��[���ˌQ�l'�-��N7�G���`���!�\A��0e1�5�Y�X.�����>fD|f����8׉p���~~�f<��1ơ���.��	�G<�q��6�y�n=<��h(&���k�'�l��3�ܷ�F��筍�I��'�D�Y��}khן�գ���u���Q���˸j��:U>hZ�
�/�s�W�ܢ�9bW�ø��|�C���鈍̚�Y�$�>!������^S���>�..��QaV�	�Sb�����Ι�I,��N��<�
���Y{ʚ����B9�ɾW�dZ���N�:[$^ʇg̋e�Ԙ�l��	݂�-��a;	�^���0Ko�aef�l�6�umi{:`�zr�l�VQ�v4Gh#�����e�!�Zke�ݻ�{�s~��k&$���D>4�$��֣hݻvֻv�ck`ՉE�^�����s���HK�ޖ[>`���|e��E��?N��,~*	{k��moqJa����q�Txq_]�K'X!x>�ᯥ�V3�]s�x��K?Mc�v��M��OS���(xl�|c����'��C��c�ߕ��A�x�c�JмE�Z���n�u���P��kc��n����&�1q� �yn��l����L=�P#C��E	zO�.[
i���Pg�TW?a�B�������0qW�#2F�0m�.ӇD�K<�7^��@���6�4��:7����l���C��ێ��	z�������}����HA>m�)�t=x�<�AW4��fk�=������C�w+���7}��|�2�V�8w��U��mmf_�|rd|=�w,>�	����x�l����z�����5�^ϟ{D��=!2y�/��:��bc�ϮW��.өÔ+���ޭᩭ��b�S�k��L�^�7�y���0�U��2;*�Y��� �"�zsf���^�`���M�ј��l���{I���>^�eF=�e�#}�uɪ;X+��
�������R^ԋR��\�]v�k:��Y@u `��-^�0�U��^�p_P�(�=(�>�]��f�l;�������)N��!��N���sln�b�TB��)Y���q:�`yXo����5�jy��yG�D�q��hv�ڋZ�۵�U*�j�,�)"����s�>|���3���,�Z�ϸ�w?|^%�=�t[�$i0��p�������֜u�_�Vqx^���� I��/� ��0\�B5):�o<��F�4噃c�̹�ƍ�8��,B��>��!2�09�E�5��N�o��_����ތ��L�:L8ݖ�����u��6���s�v������8��W���w�s;�^�\=Z�c����1D��Ku�y�O��d9�߱��"5�{��g�;�zb[L�K'ݞa���ǫ-5a��UK�����_���p�@U6�E���8��n ;�k���6��kq�]І���K��|�L?RXr�:�u�f{���[L�����k�4u�����:��&�;l�q���kk�B]��n5ǘ��g��u���`ֵܽ�W���F�wΦ�i�h�;+7:33� =1"�&�/h|��&�^�!����k݂gE��vLGJ?&/��H�J���z{psbַ��O�e�-�����UZ�c'�u�'6�7 ���t��]�|�j���:׈H�;��!�8q��Cj�G���v�v�L��V\���y_���G镁�E�|8���bm��5]��qp�W7��uD�D�n�����[[�ŋ�%k{�����$-So��j32,B�=��J����/���iEZi�Y)�֢�-lmXլV�ڏ��kfg^��;���/@��vg1
b���&}�0ջ����"|���˱H[�ټ)���򫴼��>���dt�{�/s6g�VW��\n�Ӳw��PQl	�3xj��l��5r���E;��x���Ƽ��Ő�������9�Fzp�A@�p6������]W[�ȹ����0�t@2,��5�A8��ܟ�Q�eȝQ���sft���0}��̐_x��z�'��)�W:���Y��v<��Ľ�D�V��cI*Ml�pm�Fxu�WM��Nnlgs�@{�����zqmPT��a�ka�P̞�f��T��t�!�"�.��=4SIٹ��ݾio>��X����}{"�_'#�?�A�lNO�	���z�Sz��Kc��s	͠�
�^����t_'6g,�t$��Q��c��އ�\�&},�2��;�	V��`��Qy	�_��?��;��a��`!��06��2/���vs�e)Jv�D^MQ<�g-�P�v1ײM��I���������}�秚���{�N���Z� 8B�-�1J�yw��gr�+wa�7��bS�_�ʮ�i���]ctP�B,֎��;��D ��Ѣ�u�٣6 \�� f%[�v��6�+��lX��]%��]��^[����Gf%��A��q��U)6��.^�֒�VyQ�i�;g]дpyp�:��k=0�)u'�d-�C4��׷xEV�Ƥͥ5]���t���w�K6[�tV�^�S�A2�m�˧r�u�d!;p�Z&.���U�ǄlF�c�n��b�M�ɛ@���%b�n^\��r�T�hN�yԻ���).�&xY5��-n:Gz��;�A���/S�ʕ�g	w����SX	3[n�z�U����jw�1ɹ"C'�X\X]����}B^"_m��m�į<�"�����)M�z��X�w�F�U*uus.��
�3�L�XzL@p}1��z�N�D�I�V�,���ѝeh��c�gw�eΤJo�w6↙LoV�U��h��YYj��t�SݽT�G0&0��ݥR�bg��d�B��c���{�[�FJ���5�jgu�*S��)c�?�������-'|�W&��#���,ԡ[��3��l����fY<N�ᔖ��@X�({��G��`��38uD�9kpF�mqF�i�r-��ԕ��Eؽt"�1�������,J�H�*�>B*��׀�؁����!��r�8*�e�-D�B	�"-��q��$z��J�ءO,�km�k��}s�Cm��\��'x�Tfh��Wq(���ӯ�Z$��Sk���R$vA��=���4d��o�FH���m�sAj���[ݠ*O#�a��u���n��;�Nי���q:�z�G4��}{zl?H�$7�w�S��ĦmCEL�{
��'TC�G��(L�����l�u���bG
�t���1�ˍ������
�$z.�}N��%�wW\�3(���3��4���}�흹k>�5����0�����c���*J�P�̫�ݗL���c���N1�5�׼o2�D�#�cR�l��X6uf���W�����:VA�pҵr���xff*��t-×6��*ɷC�����sa=(R���I"�&ñ��Nv�ڴ�ˉ�1��v��0SU�=d1k��t�nb�]zv��Xtw;؇x��Bs�B��ZI��
U�TC
<3��+{֒��V0���oP��c>�W�}�[hc��-=����#���"��/Pa�����k����J����Jܼr�\\l��om��:�K5N^�]��/���f=]D���H^Ц���3�V��A��o�y����M����_o^�{�#H�y�<re�'{�gt䓦��1���J����m$���'�:����}~�H)(-���8G�Em�ǯ^=z��Ǐ;v���F�V4m}�з��bɑj	%�)��q��x��Ǐ���-�����(�m��h#s!PME*j�ȱ�q�o^<x��Ǐ^�C"�9��,�&��m�5�wq��3z�lq��x��Ǐ=z=W# �b�5�ƨ�}�����k�v�5t�׍�b�-�Hy��59�SP"����Pi����܌TTx��\���9�����[�xܮW.m�-^w^9�mx�*�;��W�wv�y�sn�-�Q|��^�͍g�[���)ݻ����EE}��^g׫ש�~���BZ$�'"h��Y�	F)�
(��H�0�8�.H@�o��Wj!8m����$�j��'3&��ج�Ջm�]��j��ݮ^�[�*��.��n<�/f�z�1% �h$�Ji���$!�A&4�4��J�
�*5J$�U\D�Z�F��2�l�Pd�DD�HF��C) �)���Hʑ�+U/_a ��i�B�iU)��R�hP"�^w�׷檻�Ƌ6��e���&�g,�N`*�l���e]���H�����y�����/�̻pt�ߟ;�:�֡t�?[��M^�^�w����=��28��D���==�؏�@/�2�����>����z8������G+p���l��V�~�2DȠ�@��^�%����~���*��}��C}�&ߟ�[�u�J�vX���D錏� 1����V�`�1��,��'�P���G��j�ّF2R��r$���/2#�š�7�S��4�2�%�8ў���!��(E���Ⱥ�����5���mJ������E4]�Q�7#�&��N����בL�tgO>s�::E8x�Eu*���W�i����C�zaQp9P�4޶���I���r�Ƽ�V�׌v8���sc��%��Z�m����`��:�7��4�������`����+������t��X���w�����ir��~��O�e������/1w���c�rߎ�5��X]�N��]�p�Ƣ�f�5�v����x�T�j�"pM����f1�Ǘ��k��P�bt2}�T���M�L#q0�*�/sg�J��Wѧ�A�@�7)^�[a��Vb.��i�h�}n�3���wiİx`�Q6//�C�O)]�J��)��x�����8t�4�p^f��Ԅ� �jNƑ�;�m�&+�cT�y��Z��ֳ�y*��O� �4ЈSM
22(SM#"����"�+u]�y\�����X����(�$M
���+�ș�?�ɦ�"|�y���/�OT����W���%�m�v�����H��sy�m vk���)�ȱ�#c���7��e9�)��?x��u/Lf�|'���*�<7z��/`�,]q��8�'�q����U�q�b]��E/0r�529����:�;#�#���*�]�eN0� ��[�*z�:���4E�wR�8����`]7X4�h3*�U���pOB�⠗�a��meEU��u��6�7�/r�MH�~���7��'ë��^Q�v��q���v�wt�T��Zqs5����=�2���'�N�,4�3��0���e�u�I�~�2��[��Y�;_���yrXf�A��y����1���m��-���˺�^�5Oרn�D�E�:����W����|���8��`"w$izF#��c��k�<7W�@fQD�Эm>�f-.���p�.ܧ�/V��=om���B�	zJ�!C��g��u\�[Um
�F	���1˱0�%	ʺ���m�Ṻ*��76gI�@��%��S�nV<��Pr�e�	�u�m�@��[w�{b��kQ����)Vq��6�U��y@6m��=�U��S����s��6B��e��ys���� �M��4�B"SM��%4Ҡ�
�"�����!,&6_�'�z���������"���2<�C#Q�#�q8 թ�r���z�[�ѧۈ��vG�q�[�`�řc���+��ʀ��ވM^)�\vS:���y��֒/dO;T�r�s��AJ�,EE�u���m!���Y
z�R�ŋ��.�Sq��d�#�A1:���S��q�~�z�Ξi���ɑ|}f�X8�뫷a�s6;���
|�^��Uǐ͞�'s��%��z'�)�j�$i7y�DE�o]<�G^�_bIɽ�F7���W��p6,T�~v�e}��Qt��>�I�:��+�47�~2q�b�2�wO+�u��]�z��6�����M�/�I��N�o���P|�@jr�1Bb�Xn#SG���s��Rb�������u���|�_0���x.����^�B��Uu*�=��y��k&�Q�Æ�T�
��OK sH/N����!�=k���آ2$ټ��x�Z&��N�,�`^�-�e�*W>��z�4�*�~ض#@����~.�
}w��ؚj,���QF0V�ϫ�Ql��.���Rs4Vi�i}��/5%����f��(t��<�=��gƵ���#]M�"yw$l�u�A�oF	t"�-���!`7\o�q��2�B���B�4f�팾�c:fB^D�L����/y��B#��E��Q�E#M-4�"�$Y $���%b�]CS4��S'�#u�4�Y3��ϻ��<��0�
�D�	��<�3��b�������ס�rz�����feL�׬q�����^=�PહѰv2�WUT���,33,wD>��S�*l�62W��i�!�۰@/^��~c\M;3��.f�R;������`/�(�f���\+��o��B/����w��� �׍	�f�0N"���gL5�ͭ���� �̞HK�*R�3)�a��9�� =ŧ0�~|�SM��ă���dFF�um.� 'e��e���sȪ�P�vs�����}�A�X�[XЀ�W-��aM�5��/a��gqK�C��Mvzg�:k�S׊3�(�^=[ռ�v`��v��Ҹ�ɴo���s	B W<���S�!�.(i�d�{)�ez��Q�I��ۚ���֫�^E5����uP����\n�k
�.��ɈLKߟ�K�H	ƂJ�[q�uo�]f��̚!
��s���μ��%T�n��Z�Pٞ�;��O��&(ӎ{��a�?]`Y�nG�g"1u�_ay��dBPlܗH�_<�
m�!���l0�4��7�a�eв(�HKfv5l�٠p�&���j{�Ջ;�EY>��X�8�2���֜�<ܓ�8��a��e����`�`I2�e�1^�m+���O�E��B�M4(��BT �E#M*�E"�BE |r�ܶ"a�X��<��w��⦋�� eڕ���-Lb��qǜ��1����,1�{N��}���Cǘ9�a�5�������գ���ؖq��7��C��t���niy��h��	���
(�v#���]�fr�ڙ�>)�<��yK��B�2y��	��G�K��]�gw涯C���݆q�l�n���"�d���U�ֶ���(LxKt��s]��J{�2���UϣƪFVŻ��`��.�)隘����nw�3�`�>Z�h���Qi�,�P�X]�#�ïO���~���I�&a �y��ϯb�Y�=��D
��zke�sB�Cq��?��i�C���>L�.��y푻�)8�/�L(>�^UFb��^��e�yIq��@o��^��Ծ5�a �2�����/Z�d8L��P{yVi�Ў>>�tc7hޡ�5� �uL�F���`{�V�ʷ����q�ߙ��}��wNR������#|�^U��&���8A����5�؞�<���l���f"��D�豗/D��P�W�]��o��)��.qCr81d�mJ|h5^N2��l��K��h7=�5�3�Q�*��LT��#F�@�y�吙���V	':���ڣ���ν�-#�>iΆ��$ p�N�8ŤҼL��n�qm?��"���zВ��Ԛw:�+u��Y�E�;R��_T*�h4ov��GVJMM���/�5������E��ЉP#M �M4"��H�TU$FO{� � �ܹ$�e���p|ט{��m�5�t�ݮ�r��oR]:�F���m�g�nݒ���q6<�ΧzDC����}õ��!)�+:e�,f�?Z�rĬT)6�1�Ps�N�2o2ow�H7���r��ȩ�r���Ǟ_1w$���:����B7�ަ��3 ��/(~�y�0�o�K�t&��ۏMN�
����0���-��1
���5ᔐT�wZ�4��A
����c1V�Qt�������o1��-�p&'�ǫqf:L1�o1Uٵ>j�N!���S������˜�8�Ky�m�\��^�1��Y�t�]Y��]��Ŵ5�l+�n��D�2�N��<�~{nQ{*��P���gZ�p6�
%�D�a������c!|q!�s�=�^^� �}\V�Tg�-ts4��6�^`e
���w�Q�=���a�ک'�W�����\�SH�>��������f)T��bէڜ��cZ��[��Yj�:DƯ�|�:	\�[�,�4O��H�Zn�V���.��!�%���-���	 �Ԩ�s�K�3�c�(��bo>թG�+s���S�u'���I��?<��_P��@����೭��B�§�u�A�����FPȰ֓:*;9�;��vX��e��v)  ����TZi�A��v�Vۚ���m%k�""�����ߜ�|+_;b����<M���'��q�8��m= �����d3h7�����.��� ~80�<��
ڷ]�L�ν��z��މ/\a��Y�C���_F����Q��&��by�+�SqЇ�t¢������M����Hǁ>E8UKDcHsY5#�/�73B������r�H��h�%���o�2�7j�o�|dн�^��P�k�W�[m��[JW���<~]4�5��
v�1�Hy
\�{\G?�����Aڷ#��L��v�f!��~�{Пd!U��:��b� ��iR��R�-�^Y�c��5�3��&<M}m��P1�<�,���k�~�s*��B�߂��(�K�׭��i흐.���qM�Bd��<9�ɑs�k�On/pe�9��;�)5��HO�A`���ޮ��<�����o�+�R��"�M����v��"rX?�c�b�<��o�٠D��tE1���x�g�܃�؛)psR���(�˝�/��D&�!�2]e��y��Qt��]����c�Ԩr�d0�8��6��Hd�W6�,֜וStdbS�3��(yWq�60�o��ee��E�wW����u����ԍ���Q�pIq��Y�l}�}*@���\�|���a¯�Q�j!�}���ݱ��Y��8�;�w�v �;>����^�-���I*&�8:�oK}�lQ�3��3=�ѭV��Z�+��Z�i� �"�i�@�#h@j �H���|���s���o��\�*�ow���"+��\&��$�Jw/�|�uߞyt�O4�����}g>��C�S� W�B���ΰ^8WB��fr�f9���2*����=s��kDӑ��eN`��ߟ��	N�;����s>2�*K���<A�Gy��/umG{<��f�r�\&�OfkN�m�y<�=�K��?�WJy�EÔ5��k�0C�|�����/r�-Wa����vb���C�^��ga��|���>�򆆼]9q�'ʶ|�2a?���)��p_�	�z��$����Yȏ���Z�ֿt��_\XN(-n��҅d8����^��bIWמ���5�P*��x�-D�4/"T�xld�v�nt�l�K��opd����BN6��9ޡ����Z�g$���hp��a��o�⨼}�͙�Nnv�,�3Z���G��{-�"/iq����ԏ���]&lP�9b9��N,���y��H:�K�fDfO���-S+���2�I�k�K�=�Ϊ�++ӰRV�V�V�{�zꂣ_��� ����}u�:{�$CMv�n-�Y|�v�6'PP��xdg�"�[�wc��ԁZ����W_d�ӭm��]����ǅ(n0c���A֝[�7o�'a���&��\'*�R,��v1�w4����p���V�ݺ�W,Tݺ���ݺ�ͱ[cE��U��� ȁ���ޛ��z���/�sxrj�k�Z�T��2Ҳ7ܟ/���|2|���ˤ�Mi�>���
=�@l��t��%5�-<�����{q���5!j�K��R�{���ju��.+J��:r�K#(�k���f䎏��~�U��{[��7�Us_��b
a���qu�±Ƌ�8�Z09�*�ZR)�����fv�4ʷ'7c�Բ�p� ��h����!*�?P�a��@����5^p�fzwI��Te�0����=���ttCL�x�o��rבJ�W0�z0�y�<��Q�oɷ��0m�\.��g >A��9ې�S9����6��1i�&���o<��vi�s����+�\O��\�p�Lϖ��q�M�y�6v)��%�U��T*ӊ\�`��^�}<�,H|RS����1�����_�7���GH��fny�>�ʙ�T�������I���<�-\�T�n"��Tұ5�{�Q�o4j��	���X{Ǒ��z��6dR�����n�e�~�Ӿavjz���'�K];�s�3�O����b����%��<7��{�v���(�����'�?J/�1�]��yj��Xni�0j]��ϳ��TV纘j��	otαx����f�n�}9���7�Aurv1�ا-�����n����T5�Ǚ��:��Jj��p;Cl�V��y�E�b�U{�Ma��i�̩�9�s���k9~�+��#�hT�2i�� ��
�$i�R���{��Ov.��*k���fW4���j�;��L�����g'kػ�7����@n]����ǈ�*�^�{m$劶K�S]-�Æ� {��r���W'b��D@�Ϭ\sLL�ZF��A���<�Nv8��cW=�����	킝#�OC�5�C�m��ُ3�0�iG�j^�+5����!2�M��3H���pK����%`Kx2]��l���ӥM�Ң���o�w�_$������P�v������I��B�Z���q�k�����0����6o\!SնY�P�C�nsC�B �TV|e�8���+��h��rc�޶�7&>���Z���{'���y��&D�EИI�8X�M�����ɇ�hSf��n[��^:��N����q[6�Gs�iY�5��П����{��mRq5��r��^�1�j�'d�́p����^���A��_;5��́�FW��--]~���e��1�cdT+�옽Y|�1c�7��u��i[�#h��=;���z}�x7�eQs0ڞv�e���m�����m��^w8�2dIYu�Ү"A�6E��سC�S�V�l�&ǲ�9��	ǫm.�)�xrr��z.�v���Ns��*�����JU�m�8�f��N=�-ۗ��S��[�v�\Y�=��'�3����CX�;إw0����d���7�2oaj��!�G\���n�V(j!���lLm��-01�I�%l�2��<M%r���By x޶����q��r�
fk�&9����b�f4�e�[�ʳSMK۫�(Z.*�d��.��^]
���2k,	�þ7��l�h�ʼqp�]+��.˸����/��\듶\V�]�J�%̖�tH6�U��B�	s��ȫ�$�%lfE;����N�hT��Vo�p�7�Q31Z���obB����3'^ۥG�=��ʒan�Y�4VH�5V��ޓ��ح�}a.9M���&t����F��rid����F]��K�x�@cU�΂���׸+[�2�8��I�V�"J�R�W�X����5����sf��D;D��p#J�L��;%�qBub��(�WPa���*�C�Σ	���C7��2�hS��j�:
� v@��C�	 �uݫͷǳ	�7#�#en�D��>&�3��ɔ�"��(��H;}��ډ�^5Z"D�;}�nU�"�`��2�op�|V�T��lh�<����s;0�*h�to����%#�E�e�ѻܵ��gSWW;w�p� ��r4��E����"����ML�@��hE0��p�=�
��p�F�Ev_O�ŭ�'/e�E�z֡����[�e��_�M}N��vlw����u��a�̳;�kM���&�9��̓�Nĭ;wpR���֤.c��݊(d�/3�S�&�wk!�Ņ�m�	�H�H��+��MZ��+�eB�u��5�Yz'1���N�]��2%]g�_vV����T��*=6t�w����;&����uF�MWwuZ]ٙ�^��˕���lcCG�x�~ٮL�����E��m1��T��t�9�ds#�q}���]��%���m��Yw�ޒ����X٫7Ki�S��7&
4z)]�.nd=S�D�Q�1,��bn���q��`d�k��#�u9����ee�8巌�r�����m�n��]�k%:���٩s�Y/�����so}ki�9^tۖ�B
Twм
'd�e�J���r��y����,����M�-�{�e�89βr�s���LD_m�d�L�DM�p97ioXV:� λ��ɾ��qy�n�
Bg>�U��sh˔���~g��܂`�1cMZ�ȸND�*H��&��;Ҧ%��눥�MC;�LX�������F�mF,�E��Ҙ�b��A[�8�yJ���{4ҥ�.m���d쒧.��^��ŷ�[|�|v�V�n	А�I V��@�=x���n<x��Ǐ���*5�pX���Sx�����Q����[�骃"SM��8��Ǐ<x��׬}��nm����<�E宍@�P5���FBDtӦ�q�=x��Ǐ=z���PJ��G"�|�kƯnzk��b�����5ӧ\q��o^<x��ǯ^�`! \A��@�zg�����z��Ƈ��X��&�/:�a붮F7���kż^5���<r���x�x�yl*�*6��n[�������V-�Ѩ��g���׵��x�^9�x������oJ�m�y-��;��\����\��sT4\+}wQo�p�	�G�QE�':�gmt��v�u�{Ifu�]�hE�<ٮ��n@����r��j.�!�i��ۻ)LO��%�����~���iQ��r֛�nU��F�ZѶ�ڧ9d��?"߃�h	�d��`�"z��0����xjnQ{�PX��R���q�uUl�#o���S���;����F��	�����U&A��.+}�QaV�y��33̙�2{�n��K?:d�����A^d��h����<�{\�>��)P~�.*�!-�-e죝��=�ڏ:���*9���:W=����G��R�	>�T�N�s�{�=[���֪�ȶ�vcl9�t��t�=�p��zi �s#d3>��D&���w�h��$�6ԮJW��Gt�و�}���/��;z&�+���`c=<�˿r]�mBb�ǽz���Q���f�B·� �S���h�H�T]fK��U��cD[�+b�أ��MHѾ�7w�W����ML﭂tuW�>AZ��EV�ո�븳�-~˂o�id�!=|{��
�S�8j�ֳ��G[�<3b�!q�P3�K*�?�|�/y��_5ȃ��+Tf���xr�Yĵ��j�oJ3(���\
�f9q�_V�9��r�&Ag`��=��%A��Ю�r��T�٭���1=�L�9-��r�N�Y4m���Xr����w�x	,^� ��w ��B?!�W&�}�cƫ���&ɪ�h�$D��.������/��;v�;��e��2ҧJ&�6�ʹ����S;�'�dt�h��i����(�h��H���i�����o�a�{e<�N�IP-{�M��W6gs�5�S�R{U�;b�Lf����X��v���)�,!�okx���0*.�
���BJm�7��!�	��X�.���3�2)[�{U��)Z[r�||*�S�V�k���W�^�8�SS�8C=kʽ9����{�%�{���e/89�k���r�>�͜�[,q��j-�p��s��D>��]!H�]�z(�aa뤞ps�1v�1Mb��e-�kg�$��C��ֺIU�*/���~;Q���'�;��ā|g��Ƭǖ6�Ҹ҃�<5��gٯ���Ϛ�!ڂ��/1��<�x.����X�n�/dͺ����Oz�ڛXDHg���B��T��>������ sIzw���4 �����8u�x`n6!�*����m��nBx�a��k�	A/q�B�3}��g`0�w�|D@�.ε?G��栞~���u�0Z������|R3��K�gӎK�i{bÜ0�u'/���l���F|�<�I�W��gʡK@-�n����#�a�iC+���W�N?~������+�&���m0G$j���vEoK�Z�U]F\�nۣd�������JUwr���w�A��Oc��hY��I���v�1S��dν�a\9)\-�-���N�T�#��9�w��S�w�u9��ٺ7|�(�@T�4�4�4�Q�4PdQ>Y�����j|��/m~T�-����`��Ԟ!���S�в`�
��Eƶ������.邊��\���>M'�Cн� k��e᱒�����/[PK�����:qT}|�N�?l�Xν�~�%���d-��Fz$�Տ7�'�L޾ӕ��)v����۔��fu��r��y�H��K�Xꘀfb�0,>�g��>+v�C�Z�g%��)ڍ�ĺ׍����*�vA�)��^[A�oM{r,K�:��)�,8�Ȧf�Z_)ŷɮ�2}u��aʼc���P�k�҃&�𜮋o׫zi��|�,kTv��ݶ�\���t3D���<�����`}��/ɂ��	F��u�)�U+;��0�=�����i>P���|���z�E>�v�j�!�$�Z�d���U�<�M�μy㺼c{0�52��e?��c!��'���0:���)��ru��E��2�C����w��|כ�.�������e�$R���Ơ��K���=�l!�G�|D��a$7q'i�"���*;Ǣ㐞u�e�}��_��K=���y�M�<�;�;�?L[(ֿxʝ�5���3`}ĦG`��yT��:��u9�3_��9���G�pƞ͉#��,����vNXq�k�����L���[LW����h�s�i����]YP+C�E㨨r�Mf�&+�_�9�f\�9�]�d�=��t�~�&����ߴJ�O�$H�4-4�=��3v�騪[,m��]A1�ꅸ����Km^�W�y�HLe��zO��xw��l[;&�p:/Pv�!S�q���l!hhq���.��o�"u�T&�O�v�����'qk�<J�@VO�L����\��vf���Z��Z�C@�Hb������9����I�9��|eo������
n�6� )_l�3����o��s�`���}�y�f��f���4= ��`d["�`�6+鈜Sel]_a�:k7�v�4���qz_b�_w�lA��:ȃ�Y�8Bx�!�s(�Ws�R��WP���cB�n� ���d/q�=q�k�z�&��\<���c:��%�,8��`[s$^���J�涖��jz�͛$�hڇ�;8][
^Z�Ռ�O�et���<�8A���i�X��˥��̀�~�VNQ��Kջ���P��1�=ŷ(�_��'�.���υ��G-Id�ԑ����/�cpxbf�m��b����~tӽ�‰�$n�"���rϺ��x�;��ʹ�b�cy��fk+l'��ڱ�tq71P�ZC����	�����������\O�P�|�}��$)��Ao ikfY��y�����2��69�a�7�yK#�U��.<}D���r�]�R�m}�_I멪����
��� _)4M蹲`p�q�[�9)��d��$'���W	]7�s.�[�ȇ`mi��G����99��b�\!)<:O�e^+�Qx�6a�*��R?M@�M4�@�cM@dFI	$�g>N�3���K���w���U&���P�.i��D��yA��0�ϭ�
ǻ�T�����S�&�62z�l׿?D�V
42�zd��	�-�����$<z�S��w�j�O���;:����`�$cX��/b�eQc�.dC%m�(�y"hW����������d��f=�Eɝk�5�ڡ�;⌑0��<l��X�Lj�~��q�<�C�*hr�n��Τ�u�Эu�nc��2��t���kJ~y�W�1�S�&�ְ�W�g�4ܢ��:�ho5@��'/P�Zw���;�ޥ��p��6>;�BN3�U >��..��,B�^��a^ ;�j��5�϶2��=�b�R~rͨ�$k���!Y��^q�}�r���r�C�`��0�xzn)�үQ.+�n:�y>J��>�}��餻��p�������>*��x䖺�ڙ��I��5{gS`�OMc���p̍c�K	�^�9��������L�n���.`� �V�Ľu�|��Xo8�/f���vqȈ�Tg/v�;���������͹��&`�	̉	A�Q"�JM�P�j6"g���od��4u܌�����;Y�QڗKݷ�u���Cw!V��:!͵�mjM�RUn`��B�����+�}4��TvA�vd��z�+{�=߅��O�?f��i������;3{������w��ic��+aOG`����b_g6[��r�`��˶��3P��S�z�ߐ�VY;���<��L�P&�������'�"��'��m�mT�K����qx���Tt��t��u݃Jo5�>d.6�5x�[S�|t@r��/y}��Rȃ�1mRix4��k8�?�:����b���:��|⺵�{�V<(��Jj/�+��R�)>���Ծ��4�7s��vM����G��c�2k��+FD��G(P=�^���D�_z'������:x޴�DB�ӹ]��?�����3��_�j�)Օ%�j��w���}jgK2�mu����_K`��>1xt8��t\��S��&��3fQs��%�{��ll$i0���S43;T�3ک�7�v+�%d�j��u�����k�Ot�}�oEL,#R���<�9n\�r�Λ���-�fF�ܵ;�6�O�����t?hx��3>�O �LJ��1'���{��Q�%���_����8<�P�gA���'�\>��y�[h���p4�^�.2\`�5#r߭}l(1���΀�o�!� �a�e
�
E��%���I"���XdY����W";+�W4�b�c�c�)�F�~{B�F%V^j]��/ו-u�6>�2�s��%S����&1Z���6�k�_i�UC󏟜#�" .!R4�SL�IA$�r��j���k�k�y��G�7:�)$Hҋ4R*]�`�Te�\U�l�`��XcE�
���K#X�%C��u��ZŽ;����#Xa�;���H�OA����;}(����;ݯ[�Oj�3ޞ��Jd��9��`+
��?Lj�f�%���O�����<<���4z���B;��v��\��
���9>�J}8��y���Hm��n����
�`�z��*�1�e��0��?yNl"�*��d��体�>����cmq/������a��'��K�s���p���+���C&��q������Ր��!�b��˱�3�y���Q��[.�s@RI�i�[�F�Mv��s��o�q�yP��W^:����N:ѣ��<����ޔ�}���zL8���增�� ��	�E6n"��FM]'$q��e��3��>p��/�j���磃%�lhIyu�|���C��������6���!��x;6�w��%��Ǭj"SY�A�Q)��
5L(�^<Vj�x�x��G��N�fi�!�ň�1s�p��j���/���'�i�nz�ʺ�93vy	�WQ{��:rMCzb��G�(TY�hQ�5�4�k�!����3�a�,5I�C:�����Rv���{G���tk��^�?L��`��6��gW!�#�x����4�W��S�d�U��N�
��I��!�M4�SMQBBr{�����������:����Ξi��G8��&)���ap4H�8����t�󊎤tb\F��a��#�hnȦ RF�[X��;"����fF5BR&�˸�
��(��z� w��5ĳUݒ<�5' ���ay�5�VÚ�F��xض'��Jh<�4>��J��]�T�(^h�,�k1le�q�O�yҵ�$+�`dЗu�2Ԭ��8XC٭�Ugg�;!��C�"�(�ڽ4*�O�M�M�� s׋�,�1��Xe.�N�=׺��X�l�P2X:/�&��:ꄰ��-���\�;ҏ�x^OO'�Q�~F�;kE�՜� 	�3B�Ż��`Ά`��)4��n���}�;*E&����\zsZ˗⽳Xo���Mt/J��t�+ �W(vd��/�J8}�}�wO�fFwYo�,T�M�~
�<����f�P�\<盞�5�[����4k��.�p.y�
?Y��41>������1����ܽ����f�y5]ش�����U�ٰD�"ȭ�����/Er�z� f�ʝ;H��t�jUTऊ�t!S��c�s��j�Z�BN�̛c��!K��eم EjY�m�r�}&mv�u8��*Ѽ�J���-��2�#ؕs� ��tɚ8�+��[�̇�IR��Iʶ���X��~p����v���Z	������������Z�z%㓻Ty����㈳b��1	@A�}��}lNZ)�,�&�-T���ߩ����^��> ڳާK�i�@W�V�pbԖII�����좫{���I:��l���x��)�����z�m�˧ғ�`���ee��Xfh�����3] ��N��c(
���K���|�6n*�%��Ml�-�=R��z�IMx#{�ٯ]�!�߹���T)\���F7K�>�{gA�z��Ⱥ	?�0��s:,k?]-�f���_����˟|��XH�[c]]�S�S�L$�h���!�I{��_L���{ !��Kz����Ξ��t�[t�/@]��Nx4 �b6��Bk�v�ۺV�8��ǵ��4�t�T�C�}n!��ާi�<�=|de���!2��!�#�!�8�f�}:l{����c�8[�7%�H�g�	Qz[@�!�<1n�2'���
���޳r�����:�gS���過���������䨅��T	 ~\!i��ǎ�Լ�U&GO����?�;y��@8�n��0[�Zu�k3{��g,UU4�F��V3�fY�wȩ[���3��a�-�rU�~rJ�b�a_�Z$fr{��8��qE*��*鈱�Uo\������0���s�+:Y�(�g{.�t�se���t�����3A@�~� '�q?��0�޽ⷓGN��X��}�̦T��gL���(A�ü:W>l'蘦Ɣ��4���q�ev`�+e&��|�.0q�Z�T��%GK������~�����
(|5��~�uǹW�{�Tȉ�g�7��-���u����Ot��d��pzb�H��;�v��Z9yy����X�zÀOb���|�-%;X�ݳ9�������H���Nw�/سͣ/O��S��ɛB=S�R�|��ʈ����Ր���˂���{� ��:���ޅ�����&�}CX%��<��;~�5Z�f�ݿ������9	���jgz��7D�g<OO�����}B�����D�U�N���t�m�<�>�\<f,�լ^'�=��;�=�-
e9�-�+�C �n����;���6O$u#�օ�Y����������U��˙�^.X��K�m�$�ߏHL����9�jQ��7��E����&�FN��{��ww{��B������ �B�c}9��b��� Y�5�ĨEA`�aB�Cd�L <��{�x�������{F�����4UT�f����	�Í�혫Ybq*��G�����yY��
��ز�f��+%#�	n]����"ǙU�d�2�rtg,�K�k�B���^��*��R5v,�� p��6�^dx��F��pc�h�3�ֲ�W�%��ŵ�UqGȤ1��u��E�AX�u*�f�͛�r	�CeE;��w�"�#ւ�&_ ��LԚ8n�WOi"}���
�w�R�;:j��R�6�t�9��m���xh�Ee�p�ʖ��|&�s���c���Ƕ�C����]�\�/q�˃#�M<��g %Xr�j�c�� Ww�n�-K/fW.�DLx���Q�n�7�H6_,����v�ur�:Os�(�&��z��8�V��=*�P�x.�|'4�%����5���F����d�t{p��6�����'���)i�N�X2rbpMI��A�zɌs�k��h�=����	faՋ���J ���I�RL�.���,�B�dHU�/_�Nݑ��d;'P�媓t������\�Kk>[!wo1)CM���H�����8m��w�x)�%9YP��-un������%�X�љ5U�v���;�UV��QP����n]"�o7�����S��_��X8�J���^�vg]!��:LlP�.��P�ԐѮ�&]�-kye��q��U��Qc~����ƹ�g=N��b��d#��M�r%��dPV������we��_[9�:�[��q6��+}Y1&�؝��wQ_I�mK���;j�1-S���r�j'\؜�(l�o>��$Qu�&��*�mY��C�Ve�u��}�­23>2"�	y�D��ox����\�E%���L�5ܻn��]��wx6s=�S��7r�W�T�ۧ����%�)�s��^�x��ykWX�ս�r�_fh�D\IwF`\cB#�4��'Yc9%�3k��,�W��o���	�
���mI��:�e�a`E�V�&��n"e��{w�⼮�.S�!s+PP�"Z��oG6.,�ݮ{�썈��gJ+�'C��7qf;��|���=�Z�$�*�M@`�'�t)))��]�
%�C��J(ٝ����	�Yoqk�;AZOpb�zp5��<�����5 ��Ce��#�"�֛�V��KG
�u�׊뺫i՜؆�-�-��J���3)c��^੻�l'g��r��J�������_!gWj�q�"��C�J����a����J�����T�Չr}b��=vC솺�V�1�L�_>���H���T��Z����)]�{����M�Д�[���r�<�( {j���s��^�N���4(�]
���j�]tI��p�wi��[ju]ZM���C
�g`�5���<Y[P$�V�&ü�b���z��^1h��n���宍A$E�j	M6��x��x��Ǐ�z�`Ȕ��hE�#!! \��2 H�M6�8��o^<x��ǯ^��a"kT��^4�Q]AI*	M6�8�㷯<x��ׯC�	$D��D�R�p�jǊ�[םEr�㼄5U	��F�|q�n<x��Ǐ<x��Ӑ^��$e��&�B�F���֍�Ź{�j�b��ݸmͣQnj/^�x�[�EnTx���4jwWJ/%c��Q�Ur�\�禷�EzZ��k�ȩ*ח��/E�<V��ܯKzUڽ#K�CT{���昵{w��Z�^1F����<E�;������*�\�.#�#ދ��:%��>G!*�䁢D�rq2T!7IH�་�_h8��hgo<�R��8&j�+�J�E\���;��n�O ҝ!��{�qk��;D���EY��uf�C
��C�C"0�e�
��Dg!(ȓH����"�j���(�$�(RA��m��F4R��j81Dc����Ā\(�p�A3���p�G���k�o��OiQ`�bң.��$m��WW�<V4�qm��q�O7�E���̢��r�E_�ʛsU�:^9T�H���7�����(,�eO���A�W�#M�O��`�̧yz(�ab��l�ǉ��;���1�[�R��:ܵ;�؂����]�Z��ϋ���둆�mؓ��
g9����zv�'Ӊ�`W>�.WA���t�a؟t���G����ܡ��u�ٔ�n�KQr�N���5Q��L�0��j<K��*�=��f�U�����rf�F���9ĩ�Y���<1y8{Ou1,z�XH�T#v�\S�s�ck�#�r���*����w��_Ͻjm^5^���A��p&������cdgh���N�����K�%1ީ�&��T��VO\j��PM�	��

�%՟&O�RՁY=��=|�}!g�#>X���x��u�_��d8�O�t詋���,jM�����q>�Se����W�CfV��mi3[�SD��[��O@�x8�v��-�5�k������[鉐����t��J��o�ԷA���^����*ߝ�y�;{�9�L�V�.���Z:�B�Xϻ��-
���r�^����s�#�fi	޻y�38�ɦ�E�:��-Y}���sih	ݔ7l��g4�����	�_I�|~�)�j�)�H�a1�J���`��Ӛ�)���М��/ﲇ����!/�WT��<�
n�2s��ީ�l����<�-�
Tt��=S�@[I�vA�)��#��l�z�{xG�E�h��tv6�S���	����4�z�VO�B�hd`��DJ{�Y���N�$g4ֶtQR��ӣWq���_��m���x�n�������B%��@<�<�Z�cꎙ��Ĳ�h����jD]l��S.c[JZ��SS��şqX�J�ZN�~O�-�u��8�8�lv��ɪ"ﲔ�$s��E�>�뤠KIRkk�"@�ȹu^���0-��j���b�S���o˜�p˓���r�1�d��π�w)��"�RXs{� ?���4	�'�\�����M�i����� \��5���Q�����^����<�i�6���lxy��:L�Q��i�n^�ˀa�z`d/ �L�Uru÷�N	����@�Ni��%�����F#^�;��R�~j&�5xo��}��P�=C?�r F��0%�}���w�0�]�j:�G�]T��%�M��V\���	r1��:���`��앝8ΰm�7�=��"*�r,]M�H"�$� �Zp�fh���媵7B�&��sx�Q�j�9����Ԇa3�,Q#��ΊV�O��Ci��t�@��x!��;y��7��0k�K9FY���^�:�'<����.)�C@����bƈ��ʄZ�"�ƅ�̙qݘ�y�7�7Nĩ9�䋮y���)�i��NЇm�lky�(%��z`ea��D|��@�,�>T�^��ޤ����;f5@�/�L(qh��_�/g��ˉp&"PDب�=Cc-�L4W��f��r�Ӻ��b�$6<w�'5҃�������`S�.Ո�ѿu;V{�+���˧H>�Ã��g���@vox
����%�������5���ё{:��ެ�}�����KGX�
�����ķ�)�a\�q�1n	czd����;�5L�*��]Tvu���L[ ��r�]���ï(�ڢ)�g�۲y�yX1^%oZ�i=��]{�]�ˏ8Ϡ�c��ʏ�"��#�]@�����V|g�{�:��v�y����C ""�m����]��!��n�����s�ɀ�|]�臶����Z���gӓ4����~a�Toy����^5�0(������k���=-|�n#O3�_@�O:$;6�0݅�c-k�;�pk��i�'�y�:����^� @s�#�K�iʬ��.a��!�(�n�l�9R����ɺ4����Ms���r���'G��K�L�b�-{2�]��lL���e�WV����縗5M5I"Ho�%|��̾��>�V|��[peB�H�#6M&8���7H�1+�?_f�7
#��Wk�.�̃�-L�Q����]��uAh3��Θjَ(#LE�.��7Ϻ�4���ohő����̇/j��q�����0�-�sȖv��O�fa�����\3m�hi�=�HL��ޜ��޵X�������S"y4��&�6W��67�]��K�u9�~x��e�֣gYȓz�t��E�v'�Dʝa�'�֞g�OP� ��i�BW�a�����[��)z�.0�ڄ1Z����'8�Jׁd)%�>�;ju����}�?�G���!m�d�j�a�@{�vw7%�'n#C��Mk�0'����W���Ť3�X~w�~���{�3��7[7�: �)>�����	��~��{>���zO���pu6%U��y���1���W�я��'��<��/l�����Ёc��r����޽��������gѝ�����:�����$\^
�|^+�7Z�ZX��9�������ʪ��K����)�B'*aTZ!`�!��.f�Z��2�i]�/��U��^v2�n��o���v4�R.��Eh'k�c~4����]DJ�:�9Z����Hٕk�q}쫫<�9�J����^ޯ�/�i�^�L�� ���&��Ε�w�>�U����Z�7�	��UH��D'�?�c�/z�������c�Xhv;��N���7�(軚.i������������1K@ѥ��|��##�#� �2u��gM���v%���gn��f��Z�6��*-�X>|�$�ߏHL�ѡI��Q��sE�E�\z�U���ӖtFF%���&et�l�a ���R��p����\
��5EU5�=�}��)�m�Wym�A�g2Q�����)J�|"�m���XЯ�@ad;�|U�d���Y�n�K�������t�ﯸ�������a=xk�����Fk+����/���U�֣->�b[�� V_�!�S�o^"_�􅀾�x�6�=@0��y<.B]��2|v���U�T����sr�L\wGnR�-�nz^8Ů�3����Rq-`>Ϛ�&C�ȭa���
�g�~���Vi$�Z�z%�5���@I�_�̰����3A=sF�>P=���
��}j����`�ͻ�D=
XZz<���TĶJ�ʷg�����O)�T�ċ�y�SuE�UP�p�+=�U��^oM�J挙ʷ����"�L�Kk�w4X�(��P��O4����-&�
��/ W�3�p=�摋���hoI꫁1t�8�����Jy�v8m��u�U�����]�����32�v����<<<<<�������M�msW�=�z�0wm�A!�<ﮛaٻ����DJ���ti|�L�N;��K"�U��������dUȚ�ޭ�is4K�?|��zs�q_�0N?^�/��f
fB��Ş��ެ~�ŧ�zc>����7C���	��c�t��{�&%M��/���L���MvC�\����lY��!�v7�E�4��8C�o�J5��.��a�� �r��
�}��u����ݚ�s}�� f�8��U�3�A�º��Zkzq���i�7A8^��[�4�_�c<�Ǿ*&���4ϩǟ�Z[�.��"|�(��9!׳g
�L;�;����^���[`�����:���,:ב�P����V�%5ߏJ�����,�X�29��?b�y�Q�3��|H�<�Ɲ����|h�|<��@6bα¥��I��l-@����L�ȱ��1,`�/���s�:z���������C�l�{�tW�߮� �<�����.�)�@�T����q�^��&>|g�Y�����S�.���(f��ϧ�J�r����N��P�5u�PR`�^B�ew'_V��`��_u[-'�_ �ԏ˨Z<�c�T�H��p�勂jT��p�,�vF�@�+5�i>�r]>�N�<�̙Z�k)� <4�R��P�ռ���<<<<?�����s�I���0�Ӆ�ώI�/�ūX����ʱ�"�%E�1����x�����ߙ6�ݢ禑��'��"c�p��զ]�r9��q�O�y�o������٦
Zی���3ԕ��j6��0S�y�-6]�WL�Uru�E���Waw����ng�Y؁/ �<��4�˛e}�{�>���$,��8��<=�\ޤŸ�H�uޘ�>���{}�I�ͶVǽ�T����x����%�ll_��L�)q�B���'�ޤO�ی�����Y�pY�7D�-��ɚM�,%x-�����W>���JYk�m��d���WM�팬��4�� �U�4w&ލ�ɝ��`�,�F����i�-^~�&��6��^ø������k	�q
\Ĕ��n�� ��(��y��#��A�T+��Ixa��I1�8c�S�-[>�"3ӷ�!�l���Y�{�!������Q�/���`�����H��s��|��0}\3�#u�X��ݡ�P5���@�rMW�i5��O�g&6DT��<W�Cmt��Q�Hd[m����
^�����,��t�0��o XK�]���&G��o#�6�w֭�a���]ks���(� �h3Ξ�G��%%���N�;����P�B�#�j�n�ej���C�k.m����{�@�h������IG]rcQ^��r��w�9�����D3��S�^U��U��0��^�z���T�>a�+�O�]�"��>�4�丘�$��!�{�� �oG���X�WZ�e�Ok�ɋ�5�� �R!V����Zy�O+q�-_���)�մ�R2O2ϾTz��W����Ƕ��	�;�X�Ou C����!�]��B��W�+-u��I5K����
��A�<Bi���������_�R�b&�w�խ����oU3\���vo0CC�s"�ۃ-�pk�l�Lq�Ht	/iBq�,�bf*�Lo2N�&�2=���1�ϼ���uQ���ҍWO��n<�*�w��|��P8yL����W{+��uX�����X]�U7M��=7ԘRnt��O��$�O4l��yᐾ��P�*�%�F��%<;��|{Hk/�lx�Q�>^g���o*�ͮQo Vܔ��rWe�.�c2���L,�:�- ��Hx{D(W
��Jr�Jݭ��~f8��.�0ccy��q@���eA��%G7�����w=�}@���y�x�A��/W���E,��lͭ
�c1��=˚����
n>�Je�}���?0�}@�܊��yQT<.�P�j_�|�Vֈ3���temoVn=a���a◦��ܒ�=�t9��5؛B�r��[aI��k/�*���M5M2��TI�	�������mߺ'w���c�2*���r ��C����f�C����n%C�1�{�dV�3�-��4��}b&�}�^����a����	Z=�@�<!��[���b�m����w��E�oD��q�`;�G[>�w�גt;��iL��(��85D�>�G��Ч�E+�h��Y�א�z���Z���ޫ˭\���6^����jZ���1�� 3:�e���T=	z��]�����դөjу�t��G���5�~Lн`o�{�\3�qY���5B����I��4�&�3;I�˾*�B\F�	j��yQ̦��92u��l*aɛ���y_TQ�
��Ȉ�ǃ�l�G��K�O��Y#�7xJk��A2�F�'���L�=�����UDڙ���jΎ��������m%ĵ�@F|�|CO�F3a������
$�M.j����]��K̾��m,i��xZ�x�>VWT���0���P��I����3�͙E����Tl1��wХ�.�y$���w�=���P��ܞT5����� #� HGy��'k&�睨����Y�Nw(,�{L��W;�`K��:ʐ�.�;Ν�jj�|0d�g8�lĪ�]=X��4��9T��q{��y3Z���l��6����9���5>�5�7�y������q9���ҽї�ڬ�%���'A��縐 �qqy���� ;0���.�J�E��1\�|����0��X��hux�[�jp����Q�� M��羙���r[g��B��r$�b��;OC�����T����aQ�!ڂ��|�����=���� �}����u�2v��!3����	����h]�*�L:�����w=,�� �;��Ɠ�{�:�a��(:Baràg�	˨xl8&D�}�'���J�%	=��q֎����D�hjSZ2�iǝBP���`���U`]�"z�Q')`����9�=��r��[���A�k�ϽƷ>nK2Y*g(��r�5��VNE�#喁5n���~�E���.���q2�E?}��!��c���gt:=4;p�0�!��������Se߯�A}J�Q��lV\�w���t�0-G��Kn�O�~,}~���-��Mv�0!L~ ��p���(ܗ���}����:��|zl}9����\vQ�9���*r�TCU����i}�z���yz}���V����3��~��z9驳�*; �IE�-��q����P�q�6�ZWP�i�x��I�I�쬌t�lQF[��F��o%I�c
|��,��C,��%��7��Ճ6)����3�tڢH��q�D�����=Ǜ��-�&�X�^�zՑ~�
U�RFڻu]�Bl�9J��[[��f����9t��=D�S���q[[]b�t���DgK��r��AwLLA}���S�;�DE���;
�u����s��&�}J�E� އV�*���ǆ�Iw�(�y�^M����(��Hp�F��V���p���@�odڳ�3�7Bb�]��nPKu謱a�x�ۨʀC=�:�'I���[	��`����RP����$ja�\���k%����n2Se����ُ,�����so6L#GL��Ko#}%�ɰ��r�%f���Hup9��n�/]#K�r�^m�8��-j�`��7��uv̙R���mۅ�o{�Ơ�}*>'s��/5�A7G�.��NɅ��1�ݻ4�bI�&�8+�Q����O��3�ѣS������OT���7���N���T5�Օ��]�����'*�d˝��i��-�a��u���S��,d\B{V�T������8���-�� oYǤ�J�Mgk]j�0��e�3��"��)�O|���53o6)�MU����-N���õ գ��*Ww���+�r�;0�H�wqh�
��.����I��|���g_���w�ρ*J����=�`��Jc�M}v��`~��%������#|�˩���B�+q�U�,y�y�v��5|Yf^z]��X��8xwa�׺X�F�͹�0)T{"D�lJ��֕���Fw�P[��)�̎j�'fGڥ��gp�6.�~wO!���(6%y"JLe��һk�["�̈́�\�]�[q���E�uUA����0ogt�<
�;K	��b:���7h^�V,��Yەnd�<U�8���C�Ѝ]�f�:�s Q���ꂕ�m�4h��+FQ��c��L�7b���[S�*e���{>��sNb�zqh}�E�㈜��!�X����YF��Ѥ\#�ڟ^�t���gwS��,=�
��ʀ7�x�o)�]��μר�[��;��Њ�uu�,sVl�
	N/5���<�4��k}�1P!-���_M��֊�V$��R��9u����`�a��%�@Vy.b#��qˮ��틦��FD�F����t)ۋ���$ՙ�&d,yM��L(�����Q�Q��V��r_��n���A�q��0�F�X�Hi����@�T`-�LF���P74���E��&����~�M�#�gN.Iȗ��z�}]]�EoC0!!����=�̰d�b�����ڼ{����}O7��\��ϱf�����s
Uk��t���њ.h^@�F�e"E�I����UH{�+�Pص���u�˛x�+�*�W��m��x�ۏ<x��קb5]���c��nE�T�$�F�,i�8�;z��Ǐ7��ߗ㻶�h�cr�����*�RDjyT-®��Zi�n8�Ǐ�x��Ǐ^�|��Y$���s�����k�Z+�-�����.�"Ȕ��o��8��ǯ<x��פ�$�"j��Q�6y�񢷍\���>z��ס��sW+�}�����5��6�$��܋|-sG�n��mr������rޕ�淥�H`�[��ܱX�X�nk����rۆ�k��Ʒ�7�rŮ�r��m˕�nr�-QWwTmx��>��ܪ(�U�rŕ_>|�^�\iֵr�u���u6�����螸��#c����*Gϩr;7)p��؞T
�p36���}����_������A����fr�1NR������
�H�x���,91�&��!E�F�g��j�I��[.�p�5ZyQ<�iމ��/��(���]�1Y����D�xy��Ä\m ��)����lh���Vcw'����?�bYX�hM2��lkX�¼�)ZO�c����~ ������V��J��Oe���3�[��Y[㘔�b�+� +���� uȞȸuC�<�= ��T�uT�W6�N����`������C�i�änOL��/�\�b���)RTXsP��|�8��c�[l���҃\ɴ�:�T��n&V�v��E��Z~X����[�#H��n=���ׅ5��,� ��t���ߡp�o5�Lͽ�
���S��w��5�n��S�_L�O�з7�|�{W�`�i>j��c���B�k��^=��ᘽ�3�A�v���y�4\d���x}��)�_{��1��zW�xA��+�i�Dσ��%���c��霹PU��:��^��a��*��9�3������Xs�����>���h���	��(�4�������F%�S1RX:%j�X���vWl�b�jtMfv�%vu���֩����d���yW[�A� F�M����ޞ؉�8��b����ŉNW:��<�G�K]G8,̐T��py=z2*�*�钊�>W�^^o�������Ȥ�gV����ؿH�^`���k6Qz\�[ v�<�_����cY�Iɡ�k����R�)ge�x<B��s�9��6Ck��ڦa�^����^�a ����E�naۙ~��p���@�{M.W������,��)�����žS�*��u����Dݶ��
�4�����+�0��0�kW��ܬrk��~b?d0�l�؛�MTS:�%�vj�[�.3�,�g�hijˎ�2'�kɶ\����x��8!Cϡ�ޘT\?��i�7��l�f�4�Ne}����*LjU���&.:��֕��MF��5�W���aϐʻź�-�/P�y~��;����M�b�-||b�Z��2��v*X�R�*�
jrq��.
k`��,GG���[�f�w��ֱ�<?�?�Z�^�84S*�]�ɶ;�z[��]l+��燦�1�����G�}����3_��i���[t�/X�J�Su��t\�{�,2�� K�RL��@�5�F/�.yΚc�� ����#�9�&�o�P]O�]fL�+��r��LL���6�}%��q�=Qʣ��uޣ)oD8.U����H<����w�y4��}���ś��ݧ$��A�V��1dܷ77�FP��5;n��NJ0-Ul�x61Uښ�7�N_��\�>��`F1�i�2B��9f�]��[8��w�v��P 5�L�F���o4$Y����1�w��}�y}vq�� K/sZ:7���.��YD���w�Q����r�]p����d�D���_J�ż��0�L#*`52�L�1}
ꇡ9�}ꞬP�>(�4-�.�*rB��\V�*�Q�����^�#�Μ���2��a�UV�'ɔ����9H���zFנ���z�_���.+�J��PK�X��lƶsۿ-ǡ�yj�2���#;k�h���2�v��]����ʹ�q�^���q�qA49���C+g��u������T
�b�\����?�a7��� }��-ٮj��y�(�4$;IB�:S�j*������x�		��:鿔ܿ����ϝr*���v}��~�Z�f1��Vsqi����x܌O@���P��0}��\�u�L���	��y<�n���|��!�c>�fJ����o4y<�2�ƁW=S�?'���A�u���M]1p���a��=x�L�6�rk9�̽:���K�R*E4�E�nG5�C�'\=��sg
v�T�����p��nɼ����ǵ�5MTKA�#!M�n�Vm`���������Ju��Ay�r]%s��ZQO3+��D��e��t��5���9�*v�G��MhU��>w%Y��I9+������g\醗`\�a���L�0�ϝ��7�ʕ��^���ؗ�B|d���@�a���U����T��I�G(BU���n �~�X��̥��z����v��E���1 �	�>!�R�f�#��zf�.�{!��d�
�C�z�a"" X����٘�uYyR⶘"���+�#���/�{~�;u0���ϥ�8Ε�v{2����[�C��c^IRaA�/�z�3�\��A�q��&����q}�U�H�>�nƥ�FO0�;&9ϡx����ѩE�3��#I�oc�p���]�AH����8z�W����1���du�v'�_Rw|g��Z~b��X��L?5'SP��ԺY����)�k��o��=
�<�L���x�Q��a͹�(]�Ta�d�e.�&r�r1��Uxg��������"�J��:&)`c�"-~��ų-�S���M��s�PK�=��MI�m���]YǬR�P�3 ���q�t�<~P4q{G:��h_������ѱ8`l�#��$�Y������5g�D<�S˦�ݵ�:P(�q�W4u���^����K�|2���5�7*�(E=��W�R�]j�ڥ�94hܐPC���FlM2�:�Z��ݍ˴4h����E��t�5��#>ኃ��.Y�s�*b��2���&�'��3����{A넦kcKFZ��v��+g�;�yU/[���<_��y��o7��;*��0�|�s�#��v_��=|��cn�{\}���qW:�G
J����u�QX�UI�{��]�ۇu����VǤ>͚�ӻ qz��dq4�%�[�v"����k��U�5b�����Xz����&9��}Ox�og�WF��l�j�y�O�"��z2�*�r������7K�N.%�\�ǣ�����Q��Yؐ�(���qCD�]��]�h:������`�����a{���<��ל�����pSS�]�UJ|�x4����id/3�I��nq�x�f=[ռ�vg("�Kw�nR��S�OV�K"�o�K�����L����+�N��Qj�_++�R�� ���2ʪ7������zE��X/v@�4���N�~}�.�%"���57�^싇\��j�}���< ٙ��D���D?��P�PT����q����[.+��&�lu���"���XsY����1:j�e/_Q��^u���!7W�,6����+T�M[�E�Q�O�<�G3>�&[9�"�?`Q��q����f�$]n{kK�,]�M�r�Q��Y<{znr��z@�t`bWu7#�*��i�qR�-X�l���
A�ڗZD՜�]�l���˱���#�u��k�3�M�)��3�l�GfXN��t���AQL���p�� ����{������9��D�]
��w���Kn�?��V|�hDj��\d�9�~���A��vt�5�����o��4ׯ_��p���E�q,(��k�Q��R	��&-��P�3/����"C�=ݯ�ff:-�rQqk���ӊ��]Pۨ�q�8!��x�wvi���˲�����7p��W=٩���E*�Ҙm��?j�gݜ��M3�.��Cl4wi�Xx�ӯ�qj��@�й��9mO���7�S��1��-��5�%�ܱjzM��]OOFZ��v���G@�ˁ�Nmm�>?Z��l�A����jTO�~�o����ma�;�{N��{�0�>x �-���Jq��@��CN���9��ꅌVk���:ײ�/O�z&A=s
c��\Ո�9�O��-�=Ų/bn=3�lV��V��9����'{n�.'�&�+$�oPH�i��e@##��sӼ3�8'�RL��yW��39�g8+W�M�H[6ѝ	>5���=x�ʅ��g��qp��:�@A@��v�m�iRg��.cY�	:;:�4�����ôV���Z�t2L��Qk�k*AىoM�<6�%Gj.[`bi��ATa���K/��9VudL#
e��4�!0��nqa�9�|wud�*�ι/FD���ʗTO=�� � �@����}]������(�z��9,2ӥ"C([)��k����Z�t�f���>��nYI��R�����8�j.���k	Ɉn��J6���W'gC�&�?@����z��"�ߟZ��&<�����qS�*��+ fڻ����
�Z�h;��H{`��9��@n"�l)LC����TkZ�>��D����>d�0,@�|F�2&c����ڌ|:���w���*�[�><��VL;�yHӡ�{���c�������$V��E�	�0^��M���Gt(���M��!.v�J�'��ܢ�T4���w�H�!{x���P��}S�d�U�!��m��^Z✑�}<�<ٞ��P�vt�'���Vt��I>j��lR5Bc���R�	w���X0>�-�05���-sF�P�ҵ��A/mf��,*6�k�`�>��uv��y��3.�Lj���	���A��S�{�+�:G���ߘ�ֽ�LO���kX�9Qy�L�F�c�5��BY��Qa�3d3X.tBa�2߯���ٚ�Q`œ=��)!_��k|�&�hǽ�6�h�y+�cT�T�jTDn3:�j9��2��tƜ��1T	��M��I͊�؝��7]=����t�3���H����mѺ����1Y��̞{Ϡ�.�\�&��><�nd�������s}�M�������y��w²��F���%����C������]1�1���JyY
+>�ٽy���VU��o�0W�m���	މ�C.����9�(zTL��'������X�p�������7|r|.w�"ښi�ئp7��ג���y��%�Q�����TM���+��Q捭���=��Y�8^c�&x�AE���hn>��8�?D��wf��f�m���G�ՑSR��s.�������,-0�9���������@L�t�.�0M�^�z���t��n�xxf;�@Z��8i�(�
-�'�4��G�3�>!�>5����kY�6�z���>�z��w�����4��Z�v�@|v_�r���B�t_(MzW���8"n���~۲�SI�^S�;�����zm��R����\_�������kK�F�U�k���A�$�%�}��0��J.��)�������Ƃ�]S�Y���Fy��(ȥ����,C��0����{Y�I�Mជ�q�O�`�,h.�5'̈��/2�A�mɦS�;������$��m[GOo-�&j��f95����V�|�"�X�#�N���yo(��.���WܥLiW.���(�A���Ķ1*E�k�A��o-��X�BjB`+JU)5\u���;E�M�������T<1#E��������2����SO�`t��#ZD<s���5�5g�z�X�Ił]�8lb��q����M�f%V����#���v�9�C�V��O��3{c��/R�����F\�� �썀mr�GX|�]��Ј�x�4M�[����.�n>뛞�M���Q^��t|�L�q��	��o��s�Q��,u	B}�0�zMP<����W���l$xy������m��9���w/g
��8>�lk��k�_
<�ocU��f=!��B}�
+���K�.��ƀכ��J���$s�sQԆ��f�_s���)Fʾ��zik: C`.��:d�[��n=5="w6Kw� ��%�9�w�WA�ʚ���fBd/!/wO���3���A�o����<�ֹ�YIr��ԨW�!yx�.���⃍�&�1�k�d#�������C��gM��0:ב�*-�5s�T�fA�B
��!��୹��ɪ�z%=y#;�,}׺�Z)h����2.�jO�ǳ�~*��?�� 7X7l�x�K�=i[*��e�rK AmҔ*�j(^��$�&ՓH��û/r���<��O ��ю�U�r̬fIBKˮ�Y���p�^�ߠ��9��Z��y���<��c�����)�U����䕰��M1��)7�s�o��r�r���7����!8�1,��bYB��n>5{gO"���a��}�zΙg]o^jB�X@���EB�� a�}~$���S)Rkk�<��C����z�7-l}��*�]r�G@ƑȘ|��Ѭ��q#��$��b�sȥA�qE�4J�/�E�q���~) ߥ+��|%W�A;#�����t񞃸-�򕾈��|޽�-=;	�yl�]����ֶ��O$���Q�#�Fs���ЧQ[�z��P5���3�U:���A3gޠ�v��xB����^��sg�ŕ�lw�<5�YD?��� =�ǿT���h*pٰ�3�)�׋���`��\l�R�}#��TW����'��U	ѵ�;�]���=���\�b���%�X�/��֨p�τ*	@߹i#�Y�؁x%;ӈJ���K"u���u��d���#�\�v��C@�6�6��L��u�n�d�������┌>m�r�9�xo78[��Kɝub3M]}����QpLN�r��Vޒ�i�s���\ڌ�v��i���)176ae
7X�@��� ����R��p�+CX��Z���rӗ{ts')�GhH�6jԽ�Q3%���w�{"�OF��샀�˺��p��P�E^���zZV�hH,�����f{IX'�j�]�[2���*�/b��ҹ~t*]v�,���uն@�/�[�3��:P�a.�����*55���v͗���.���Bn&C����a"�J.Ի�iť���&%���9Z�ZouNnl�7V��N�5,��W3X�|������m�n��x��93ꂱ���q��{tGT�OG�Ȥ�$,��f�����l���%�%HE�<�7wP�Y�!F��h��IW]�i�ǣ;��X��T1U�剹LCґ��l ���Ze���_d7��}�gt���"(�fTf��C�qu	ܺ�t�nι�)
j�d��8��R���w1f����$�xN��^.�%�5��y.ɻWيނ��Ś:�z<�����s��j��}O�Xh٧�M�+��1y���a>��pҪ�KK�5�]©)Q.nŌ�L���d�D��y��B��2���O�QPh1}l���%���Wne�"����2�Z�٪W\�����[��Ƚ���r����B[�d=x��4�E��*cm+��w�9��ܥZE�V;�T
�'4�[(V�[��al������bH���v�4�;�P�6L �r5��0���U�k00�2�,��?�-M�v�����)5-�-�O��Ո�v�]�BUf�l�`�{�r�I�������\{%�Wg8�5t��\��3J�x��l�Iֹ��[�t�̶͋��R�2D	��h�0v��fs�QS##��<P�xv�e=�f�r���p��vr�Y�j��@ξګLe]�bТr�32�C4���u&�|�SU���fҺ�o�SË[��GO��z��5p\]i=�Wܫ4�Ĉ����¸�t�,z�˛�
5�� ��I^͔�e�زk��5�K���#t��1�	(�Ǖ�4�pD����5S�(jOq���.�U�Wj�
Y�1+��X����lN���u#d�%>^�֑�-���Zb�h��N@�,hO-��n˦�B/��w\Ng�tC4[�v��������N�7ۘ9�w���Ҹ,�K-t5c}״��\�����vż.���:0���p͠���X�����IJ72�W�w������A}F�:�����$m�.��;:�vt~�6�ډ���С�T9��Y�h��anSMU�\/Wk�3&BwF��,������TC0%&k)K���F9�X`m�4�-4;�$�^R{��'��Z�I"SD�1+�8)����4��7���W����mx�$��ڝ��[�ˍ�		$Jm�o�;x�����Ǐ=z�0�:! ��Fr6�[�����nZF=tێ8�Ǐ�x��ǯ^�,�To�5��عr�B���E��
�=tێ8�Ǐ�x��ǯ^��Ed$�UE4b����y6����[����M��8��Ǐ^<x��תHI'ںF�����G:Q�s|���7�q���e�]�x�QIF�݊�͌`�Qd�]�$iwp����9|w��&����t�X�jTEE�M�x���X5�AI���꙽�R�t���h؊M�q��"���4��,�$��gu�69WI�2X��,��6���j��W7���I4Iy�����ݼ�ӻԁ�B
8AH�#�mB��L��(�� �bj�y�b�yt��g#g�L�Vd']���5��:ɴ�N�/j=��wXD�j�rl�kJUU�^oP�l��(%5�F��1��m`dGl��b!�t�[�E�mDJNLe�Q�@f�<�A�M&
(Ap�#H \NF�p}�������\U{��T�DΩ��7��%'��;+M�7��N91P�ڙu��_w7��&��cC��t�Ǆ�Q2����룒A��4�ͫ�h��8t������'�dwsa[�]�F���Qk�r*�	�Sr&���GX�$�ޭ�U��@����N�e�X.(%��͹r�����r4FJQ��ty*���RR�L�TK��\�[w���� �cqК?T	�
��r�^8�:��\񥗞��*�u�ngҦ�R�ɘ���>⯗ѓ��H`��FS�x�%\5���w�(�z*V�2��ý�'�����m_w�r ��!��E�a	q�;��vT9���i�zGe݆Έ�1��c���HЎ�. �����j�{"�˝i�v.j>�X��5|�G����r��A��9�(]�{�I�l��j���K��y{�P�\��F��W�u�̧ԘKǺ[ 6辊�荃�Z�b*�*y��v�V����lZ`̔�c�&VavX:��̡��Y��U�br���>��4���S]�8�rB�X����a�a�ԶhsBF7S��C��ҩm8{z�H����e;ŭ0~�;(�:���E�(�y#UwB��}z,����%�ĸ�xxQ�gw���+�o���+��.�]��yr�-w�[��c��K)�[�Na��<�p1�L;Ŋ�7�E�R��ht��{�\�b�D� {c���-�y�����Dp���
a�0��H�{��]�zq;q-N��zqe��Z�O�%P��6z�2;<�t3V���	P�{����K%�?r=�DA��U��(ݒ�`������d����,ϞU����li��ռ�
o���ܒSߏwX��8���ܹ��@���
����+8osc3��zbjU�m�ם�Q�0<�E^b�g��T�'�����~��G���<$c�&��軟v��>�}�c[5�<:�=]��9ew�
�s=,��O������t�{���)P[[n�����r�r��Q'�={�ں�s�׌�vG�q�]9+�b���j﬘C��3�5X�HoJ,�YM]�X͑^vPy��!���nv2.�Һq�@�g�R�n��Jd..�/Y���W�x�_M9�W���A��^u��y1��]kfc���P���"�֙U�#���	��?�����o~?����k��ψ���5����gy��߀^����EU(a����Q�p�x�(x\یS=G�GCy���j{m{�f�m�
��Ē�\0^:lB3���(vآ��~}���U/9A�wK��ћ<��6��KL�����[np-����n�O�er(9A��8wO�:�g&��:�KQDϖ�״9l���L�yj1x�ٽo��	U�P��|���u3�&�x[�����s������uJ�8�'�9<�J�����F8&`'�Y�y�
��2��Ӌ%e�z'M�*���'���}~�ؘ2g�Qwᔲv<����0�WH;�{���fѶZU�
�wӄ؄��u=��V�&3i��hg3�G1�țO��0��Y�/����2;wO�5���|�����{���q�#~�P/C�xڎ������%���E�b�V�D�7<�&u��Q�$�2:����W�a��`�-����Ð����KRv+���S�h���ܾ9��_�*��ͮ]�뎾�vvm�	{�j`�y�x>Ha$���z�P_h�GD'���u:0R��V����0~�1���fzB��(� �p���Z�U�g�uVUx�}��y��o ����h�,ey�.ߘ�
���R�rk�ޚ�����ǅ���\ED��@�M��6�8wG؛ë�g:Be�tt��Rԯ.^b���]v�]�1��FdME"u7���3mO��l4�7���o`F���ڥ�V�\�gO���)�=���7�n �"�'� z�.i�ƅ��
�P��f6����W��*޶.�!#'�y��x�E.��.��Z���K,8�e0hY��O��}�ljќ�Wnzv4�W�Th�ߒ�Uߚ'�$�{�%5w�>�� �;�*�Uz@� ��;��7�O��~|��u���J�[�GE�O��<\���6܃p��^�-��k���ՕS��߶������v2���߯���]�Do;����c+d�Su>�ʌ����I���l�y���+�Wc���e�_��=��Kݮ|��n��)�u�C��e�����)_��W�u�y�[�}Ƙ��r�NA+1��M�����B�����NVd�g*��;�,��g#��}r�D<yՊ&@U��뚁���Un��
u<Lۖ&.�J���wr��*<R�U���yZ��$]��t@);�xxx|<<)t��|l�L=7�;�6f�Вe���mc����?M��꡿{ҽ��R���w�1�}���7�������{�2�?v�s����M��?G��H��=�M2��[H�w|t�`�F�D�dQ��j[M�_�vI9-��MJG�t�yܬ����-����}�` ��.x�ƥ٣)<�Gï`Q���7GR�}�r5����X/��4G��~��y�ȸ�/e��
$��䖯O^A(��8�����B�^�Z������0�/zң3f�;� ����w��~�+Byp�WJ}�u��`���r���1�N_s8�z�Д^+����޷��G<�ɹ�yb���no��7:�|�{A00A����֧�k�;I�fK�S�!����K/
�2���M<M3���r!(��*ᯗu��Jxgm؏{��P ;��v0��m�'u����;�/C�j�1SO]>�����X��������(�˺���lNgp�v���EB�K�E�-�+19s(b}��� �ǯ�社c�j��y��g�J&�,I��ݐ��v���y�oMݓ�g��l�R�=T<�Y�Npvd�IV�
��g�*� �K�����=����ع+�Ro����s9���*�X'}�V��>���5N��內�++��\q�����a���@�!��h���������#��q��W=[�֕U���4iwI�t��z�5��e5�"����v�.�:���讠6XI5�+�����q�%jf:����W��n�zęYx�x^s	��49���lʗ�24�j�+&�[dE�q��'wLaWڔ��� ��T����G�t$P���q�A�y��x/17k��]���چ �}#��Ǆ���ƅ,�|��sw���9ӧi�7�w,��Z8��ʂ��ztۙ,K:	�X2��V����nZQG�`��]<z3wPD�oO��N ���ڣ�������JƂ��ˋ���i�z�y��V��Q8��Q���
�;\xs��B��6�N����"â1.��;:��Ϛ���[����m���N)0~Ҳ��4Ȳ%N�\�V�.bk׊����pVk�H�#��߼<<<<<<0�7~-�᝙�Ѽ���M?�U�ff�e�qַ�Z�;�-��ye+���a����0�s�B|���Ѹ~��Z��s���|�
�ƾ��^���f��0λ�;m*�}[,�(�y�:B��]�Q*Zf�/�&Cߥ���N�v���v.�3L�RnN��M9�[�
��'%Ɂ��p�N��'}V�Sճ����l��d7_~��KaU���̟u5��@�H�{y�3��legf��-m�� B�����$�O�����	nEP�+�Q���9^6)}I����y�s�hw\�A��2�t��#�>��X��/B���p����E�ɫ���KQF�XҵFք�]��y��tt�ȶ����X=`ц!�k1U�d^�~��qP�%�+���|�1�r�S��e�>6�@4�/V��	��f����~г��y6��D�{lh�9AQʱ�����Ԯ��U�V�{��}
�Z���T��f������6��:�J3[X����"����)�+~�8:G.������$F�=�b��KnJA���_��\Gb��K~���בֶ�a�ǟ��Q�k=��^zɤ>��c���w������=gv>H���f@`��@M-�`��^�'�d8Ւ�.�m�Vnî��pɿ���^��Ž���b�E(�l�8���B��3i<��Us�.�NoM�*�����y���8Xq�	�?e�z"k|�	2� eF+����(�p`������e%Y0��H��3^�'�q\(���#V&���z�?xed�;�]ޘr����~ƚ�/{ɔ�,����k�W��UU�\����/+�����~腬�D�ڻ��j��LJ�ņ�c���ُ�d�>7c�5�J��BJh�$��5P�>�K˛
>�c�5w.%�g�V���oZ��&0�(�+�	�����=�"��3΂�h���q�0�y�[���P�9�U�z���q#�t�˹����ˀ�7];�I�c���O��Sh�Wd'�#�_�� ,ߊYE���^4�
�[�&�j 8ˮ�i��ON˫��������D(��N�*x�UQ
�'-8S��sDڴ %�V����Ɋʕ����n���x �n�ad95�[�:	}0d[�F݋i�_"{�*��$&q̷��C��E%��������>�� ��)�$ҫf�v��ō�f�ʂ��{$Ĉ_n���}ޕc��	C��&�������ѽ).bx�MH�~��sx�+�^���<�3�! &~��>��e�F}txS���Ҧ٪���w��_1�,���Cz�"گ}|:%"X�l���ޘ������;BA/7VI�}���>�^=fт��v<g��ZͰ�;����2��>��r�b6Us�S��UW���Rݿ��T�z�[`G��������p:X
�7$�{*�6���^8�)��ה���2bz��yڸ�����_�n�X�#�n<+R>�zgx�bv���F�k�#�2�k���Ot���ew�8�Ϋ��]�:�׭DL+��L��Ԓ��]�!_R���	�#�ϞW`�W������E+%���e[�2����B��$n��#4�@������4(X.��7!��K��&�(]��$��-0:!�OI{���	r�wm�#x-"����z�A%С�·��7˕�>�U�U.�z�$��/����Ql$��긲[ �hgL��6y\�i֒�򥩷vrb���N�V��ňu�(.�}�uf'Z`}�������h�=|e��_�U]�[�f��)Y�jJ��u|�\l��n<�����N�n1���\��R�-l�:�Ydt�xƒyE�ں��/���ut�Y़��Pp�N�^@<;T�R5v���I�fz�.4C�]��8|�*yH�/g����Oi�]JȄ��*��
&<�qM�x=�B
/���n��0MP{�#r�H�"�$���+���벽�eV��.�{ZN�cx5�s�%a����o���JG����.WՑ*��:��Pq���VY�l"�P�J�֊�F��+���X>�*�+u��\k�8]*�０7�	�+�M���D
�����0�%�>;�^T�gR#y�yW�r�l���; :�4bYD�=�MP�\��q�[��nV�؜�{����[�2�`�gC� uB�fc�BL��t� H趩9o{k�eK1�wi�!C��Z8��4��M�s������;�:���+^E�e[UՃ�3s�Bm֐���1��ȌI�pl���Eޅv3s,�-jh��8�>��Jvr�����R���K��r�eى�3ü��&��k���e��/�n�ݹhޒ����n�nu������3y:)�:LT�n�6��'Z��2���ug
WpK ��o��ɔ�H0�y����J��L6ҭ�d�w�N��Ǖ��{�)�Q!��ņĖ���F�BW��*頦�4;b*n�fwW#����qkj�;��e����%e����P�FwZ{��ؼ����.>��uq�M�	;�N�=C1f���zJ�$JU�kv�m��/E�]}4]��O��3���f^�WI���2������b_u�;�|XC�kDI}Z��>���M�Hx���͓��#e�K�h�^�[Ua�#5�n���p��	�d˶l!aε�+Z��;z�;�����諥�฻���h��B��2�䳶f�W�~�Vd���������=���a˧}!�d.��,��&�}�4�ő�ᔬ�5bdT�����	�5��7;v�����dՂY�B��Cd"�CbR�\'�1"��9N&�2+p���
á�'Q�"�p7R�y���ܠr:a��A��4���sL5�*n�ݗ��>ք���҅�!�-SF�7W3�>S��Q�e���G]���\��� ]�9RY��oz:�FA������`���7|���"�^��lZ�j$i�l���f�]�����݇�2n^���%�.��t5�0�ە	����e�C�v2�1��K�2���Ux,�O�i�A��Ø�vcCf!ݪ��modX�n�8��&IUl�eA�~� �}x/�w�L�g��=w�9�5��ۮ��*���q_I���nC�N�\Su�ƌ�_i��s�m[��^���5��^9��
��sX��԰�A
�K���
[���m �b�i�+x��sغ�vu�3{�.P&�b���T�{pq��;�β.>��.��� ~f�k�]7;BxDz�]��E��NP�*ke��ƙHe�}Ҏ*�U�m��ɉ�ؐ��]�d�f�B�(uBk����T���f;��&!�R��׽:�[Ѯ��2����Cwnr�ӠKm��J�w��i�s_;j�{WDCo�|R84u��ӦJ ۦk��N������m�C�(3#I�N��d�ΝwYI�jy�>u.˓.��;���j��ʼZ��n��ML%�*��q!s��o{���=\�f� �$S��gsp]�4ZQ��Ӡ��������ډ}���Xr�}r�C���t,�n߆���	�3f��0�x��,څJb�N�L�o2m��Ku0�M�S(��b�Ð#�+�Um�9�or���������.�F4�D$h�I}Y���0�|v�bl�T[�]������R�z�����<x�Ǐ<z��`T�	����2�:.�ɮ���ܸ���^:�@���qǏ<z��Ǐ^���w|�xed���~+�7=y�ch��X�lL�E�)���_\q�Ǐ�x��ש�����D�&0Zer�.��_�nd4� �j5�=m�8��ǎ޼x��ߕ�i4a�����E��ڼ�s���E��_+�F�7B��H��Q��1D&��E�˻�ܡK�Y* ьr����h�}��I^�v"�n�,B��ſ}t� �UȲ�=�;�JH-�׿9�����%C2HL�s����3xŹ�}+�K���Q$`{p'.0�u%��NF����RaI��DI$B��)݀����TQ��u�n�{��ݧ2�f�1l�E��*ڍ��mc�:yK�euⅼ&e�W����ײ�7�7�W7d���1�c ��{������4C�y�?�{�x�ٮ�o�������{��!;�J��&`��w:��oN!�,��$�`ha���<�Msf��~SU�%{�J���K��t�j��'����>'�GsS���:CX��yP�C/��;�I�+7�df��'�"H�%�	���tJ�
k+{H�W�
$�?;��{-W�@�NԲ-�u�vV�"���^�9q��7*j����l����qʂ5�����v�;0�09,5�7�L�.K��dI0�i��74�v�O{��r�����#r��`�}��a��o
���ұ\��rհ��T��g@�ȫ`�`��㵹'T����{^��3�pF�y��yP�d�IK]VK.i�u������^7u���ϵ1�׳�PJHs��j����=9��WR?~��rY_�jtFF^oC���s�n`Q!�V�9]��S�����k�{�Xs,�Ҭ�}��l�eD>��Թ���T�-��Se���V)Y؞9�qهe$,�,�P�U)�X\f�ގ�{{�r�t�eٍ�����5	���c^^��w�r��{��-��Сv�r���䑔R�d,iF�o	�O�%���t$iW�m�����#V�O�|���� -Y
�3���u�+�u��2��M�T����r߫Gkl���~x�Qݷ�̶�7��+ݚ+�uRi#<��w%�����~F'�'P�N�Q�l9���=�u�匠�+�^i� L 7u�~��֛�_/��qFP�N"[��7չ޻@8�T��:r<��O�Ws�X�d����mB&%�FX���`�+ν�&Y�ގ�3���F���t�쟩8[a�_41�d��/
wk�߷h1�kR��Y���]��D�#� b�4SZ�h��,�x��J痏m��~EtP�)P��4��S�cu"�.�N^d�\���,ƤV�?;BY�A<�WJF�?NM���A
��H莼��-u2<���f�Ab��j��<*D�dzR�C����)\jMwm��W�L��o(�xh�_��W��k��a�WLv^�I�B�AڻU��!�KK��FC6؛����B�;�U�N�>���>�7g�Jպ_�<<<<<=�)�/F`���e�yV�7�f�����P�Œ��ܽ{�˔R��hM�n�Hwxfx��ݥ��9*GBM�#6�����n�aBۧ�(��θ5Y9���\�)^'�X������yI��]r|{2E�9���)cq9�i�fv0�3�������	���z���FU]2]�MvUUv�s�qk�N�}^8Й�R�B��!�.o|2�Btxk?-%Q/:�L�|�a}׹F��"9�"�M�r��e1�K��c���iDA��{S���޸�c1��l�0�^��[����F�&����f<mݠ�rF`����ЦC�n�Q���5����=4<�V��|�d�����ۡ���st����s��n�z�6������)X�(�x��O�6�m����옉�tW=\��Hp0��g:^��q��(ȥ����U9;M������^fh�2;������F����Ք'���<&q�]�_�������fj���qcsݭB����x��Ssז���uc�#gm�^����ܵc�c���n�=�i�G0AJ��7���-g��F�F��}��d�zt�%�;2��dE�`{��j�y����P�Jj���j��Q��c�v������o�_;��\�ŗ����[�YȮ]��{�vc
�<W^���f��M���@��!��- m�g7�q���eu`�J��`z�^S�Ӗ*�j�Y7Y�DM]9�u�
������8����v���L��wf�ް"�K2X,��uݩ�oe.�Pwի_,f)/H�Rh
������p�/�s��-��ĈÙc{�$��W5 �9���d`�P�R/%vm��s�zue��k���,q{=�O�H�̵_e�w����`Xoz��j:opr�冣6N�*�yf*�g>��vW�_Pc� EeL�g��5�Hv�5#�=8�s�����{s_��TI|��C�ە]6�&���(6�n�W��.����e�q��'o��g¼QS���R7-��0>m�C �@V���&���'/➬�]]\x,;�˱�╷I(��l솪s>�@�&��Ɖw�R��Jv���Ц[���P�����%�D�h26�nח�*5n���oA*ͺiRT#��ŝ�jE�	8.j�lΕ�����b����hv�����jα��$>�kE��z�;57�892U~�������ٿw�jX7�Z��6�6V�Q\�
㌹yo>���w�m����х��m9���� �g��z�l�j3WǞh�)wp��t���8Lx��t�l����/�ǚhU{����g8�Uk��n�'���O�6p����t�E��l��p�{6Cv	8����|+-N�Ǚ���_gco38�r}����/�Ο̉_k��1d���_D+p�2����ʪ�͵�a��Yں����[m��~�P���!�v y�A�����	p��V��q�ٚ㗊.���w�>}{�2-��S�^���Us����'���ק�X����t�>�I4��"������L��f�Wwa�6���ӑ��B���*:��ټ��ޡ�C���B3t�-LuW����yu�]�z�c!+��ɯC�N��j�Vh(���2U(��ԫ�:�[QU�A�αp�4v^�(���Ym�:�Aޑ��
ÏnZ%��!���n�n6񝍒��︩���N��kB�²@F�ZQL�l�uf��A�Әn�/r�8rͩ�N`�xN��U^�L�=�C�9߅���
��:�=�/gw/]�Hݍ"���ә�g���&	G���x�+��l�Ձ׻~�Y��-T��٩���*��7d�>^��������t(��wLyU��h@�h�ǒ�IU˹��Yf�;N��{�w��|yכ�b�x����U-��J����2�MroW6vǺ�8����_�G@\��f�$����R�?t�V�aM^����)g�|����^������=9���hN����l���C.H#��%:��e6����z�=j{��1|Xs� 0[��dhS`&�v8��@YY�,_�6��=�h� ��8�L���n�������u�qM��f���w�}ԇr]EO�Ůny�pw�_����Kk��zF�f$8,$��R _�H��/�$7cy^F��]�(;����x/��R|��Y��Bw���t��{V#ms�[�[��,A��$�h},n����YP�[7�Y�N��^��Wv����HL���N�%%�hͰdZs��S�a]��33uY(\ٯ0��Es���4ɋ1�7FѮ�\���$펳��~��������2�����l��Ӎ���uv,�m*6ו��G���~�>��#�k�G87;Y@�s���!~2SQy�m��<�����j���c�v�K:��.��3I^��&���jb752���<��!Y�������*
X^R�{����S8�^��6;v���$z�f�h�]��vn'C�~�^��꧳�[�I�9ϩ�3�0EЩ�`Һ�E+F��֟fڛ�Q����Kk���5�һU��/҅^�Y�AP��R�G�*�ܹx�k�_x� ���l7���u��M�H�p��z��$�ap��7�<x�=��\���2N[�V歬@�.�D#@aB�q�{�R���*����"Wf�'�����#�=-��:���x�!� ]1�½`kq���_DV�䔱'�iƳ�݁K�"���s=b	�Rb$��"� ���0�r���mw�s!�@A�����MXz�pð�3^�nteְ��rt"1���5m��A	�:i�с2�Ew!z�{g�3N�nhB�}��K{v��fV5���ebk-�T�݄-]��2����/�����y��|n�'x�Ǝy�[�:�=�Ρ�~��:���y��:��u�u1Yd�<�J#���٭S5�\��f� ���VJ�N�s{o=�`K´�n���}<�1Q��Y�ɰ�1���t�LAJbޱ���:wJqײw8�uY�c|�v�����8<g����ۧw�x����n�?C��r�j=I�J˿xu���@~�j>��-���U8�ff{3����Hje���Hc��\3V�nkУ;�y�V"�S����a�g��a3j�M�g����ǒ�Du���t`� [��`��u�^��)g�7X-��`��v�Q�ָ�ӿO(x������j<���E\�S�h�{s��%u�
�p�f��_i���C_UwY�;܀�亞ae=T���~�?cHoz�V����Jo��.6��NkJۤ��K����XИ��M��P�h�0MS��1�ꋺ�t�{\�ZϾ�c�&���K\^����q����w��8;}�Q�^\��ZO-�%q%Ν/r=��.����;I$��	U����������R�}󃵩uWmӋ �G��`^���]��t�C��`z����;4I�<�K�C2F6���wM@���t(70�W
f�/79�Ncr��T�8��+/��
??�nɯ���H�	X�g��K�����o�Q-�����^��΄��A�ID�l�s~�*]��juԏ3v$<\�`j�5��y�U�+��teo>�;<STW�Y�Y�&�����z���T��7Y~�Y5�\Ѥh/7�x��Q���59���Q���'��,+���}[�肤A��j���F����=��vs���*N{6}��������×H��>�`iKt��y��B��2�;�/�P$B�"b'>{�f����m����F:_B'�G΄������77��mZ�:b;�7�)�g���`=93��`����1�b���(��L�GO*�j;S��n.�f1���T"ԣT�e�'�ۋ�8�̘�r��;�F!�*���������
rl��gDݨ��"�U�(�s2|h�`�$=՛t��g\�sM!r�匸'U�l�\������¼<<<1(ݬA�f~*(ڨhUNr4��a��2)�]�ޜs=i����-� �q�a�f��J&�M��u#�9�Ҏ�#�i��!UÃn��{���4��k��Bi�]��þ!xy���c������W��7C����8i;�K)�`"��mǲ�x������*X33O��]���w�"�etr���t��^:���I�i���әe��Uk��9l{��z=*��<֕��5��/�Ɨ�IeT��Q�ʉ{�*����j��֮���xJ�죷�*��2�Aɏ]��Y���*�J�	%�}�Φ�j�|�#<w]��W3�̏_��t��,w -�H�)di��s=��\01]6`���1�׾��v_X���1����>hΞ@$e�����j�WW�fN_c�vvG]�@6�S���Y�pZ��l¢[�0���1�k��AG5)��6�T���Y��&`��;=�o	�yӦ�y��;�����9�%:Ř���7�4F��"�J���Y4'n��[���1/5+���4mCs���`�v�Zf;�Ji!}���8�dk�e.@v�<�l-�};��M�-Բ2a��M�+�Ui������f1q�7v�CSf�^�1;oe�i��xu���r�K�VG!�%�w_7�k��j�>�50�\L&ulڳ�LHY�Q<y0����]�ǸCw�!w>��qEEt�5)w���Ry�/d�8����LZ�3�W)fc\Xvc������f'��1^:�t���Kڎ7����U��Cj������o��������=]T����{�v�N��35�ZC͎T�$y	���-j7VaX}�i�}G��8+.��}3��ŋ��阘�\�sҺƄ��Ε����"�$'	m)�d=�1�)�97��֛�v���l�2R��1׺�L�����ff��i��6�囙�r4�\b�KgF8�G��5|2�<X.+�!����]��X�2��gW�w�*�aL]�v�ѥ�j<�V6���H�s���aA��vӇ�o��ʷWkLس���@����rL>�͑^���;G3o^�h5���b���N�����#dN�%�kIf��n�0g,8.գ�����3�/�t ��B�.�:I'v1�IFYzI�P-���]��7~`<z���`g^KSj��O�&�ә��;���8���s��*�-��5x�e^����㽨z�;�t.����zm�u�ٽ���Gj�t�;�W{n�$���q�iwg����ݵO(��Yb]�e�/Q�̇�˽�ˋV��UݝX@OU�}]R��2�fh�i5�Y6��ݰ34�n麔c���8txr�j��R��ܸn�	N1̈WEzб]r��_q3wM���Q2E]�.h�Z��Cm@�Q�v����>����m$Ճ\z¥����5V�Z%А�Ɗ��i�E��q�H�����s�չG��4)g��k���D�=�k��G!Fc�n�^\�b�WKСE��:oZJ����1�ռ(i5��6�R7��D�����z��wU��x���wU�D^�{��}lh ,U͜�F��{�&RQTգ\�ܬ�1{��X:���t�a��:��ue�h�_kB��r(]&�v(*�T:�*���kfC�w���״t�&���r�Э�W%]�^�9W{�]�Lf�]�)^gtL����w���2� i�%>����fdk�Z@�M�[��_ms��Օ�+uSE>��zXH>�s�vH|D��e�ʻ�UPQ9I����jݑx�������ӆ�tM��xC��5`w��׏���
L�#J�,c�r���]1%{sh����ˌ�PӶ�|v�۷nݿgnߏ^��.W�rQ!0���xH`�XD��Dfz�'頌�!!$*:i���׮ݻv���|����7�]�h�\�� �~wXـQ%�Fȕ%Q>V�	I*:m�����nݻ߻�|����7�(!A_W]�۴̆=wh��;ל($]�RJ^uW"F&�^n��������v�۷�ݽz���HFHB>.2����B�{�����݂��߿^HKu���R$���]TPJBȇ;����I;��bM�F���u�.�qE�o����|��d�E ����˾x���s��2G�����$����>�ߝH.�̲���
��������1��Mp��v ��w����C߮��WcK0^9�JPL]���W���n�^��{x�[��z��� ��� E�xA<���Ei�HI�5Ċ&�?����J(� �Be����#��kTڣvҴ�S�%WL�]�q�v�NZ�(�M��Q+�����yֹGsd7���S$��*^Zl��$jF�U��i�������d5 �(�b�(�D�"$�0�SA�F1D�[H{!�	P%2�A�*��.��)����s��xo�Ni3:'��{��L�WC ����=��o5����9���S�"I��f0��c�]C���V��[y��gVt���m�Wi��"��l��t�_u��m�n����ㆫ]�T=Lug_I6���0���ʳQ
�L\���7��蜥7�L�t#ĉ6"�����R�/�'ͱ�V}��8�v2~?Z��j@�D;U�����~�Vy��M!4�	C���@U��X��wL��ۧ���]�JcS��n�T(�T���4+��p�<+5���3��q&J��u�����O�ǚ�P/�qtؗ��f�X�g;������Ed����QV^!M��8������%�s<EwKO�
�^]��-������l�\VQZ�+L���h�Q�W�������R�k�J�pð��B�ɫk�	��������P��䁯^x�'Imfq�J"��~�s(�Ķ~�,ȝ˫x�["�n��f뒖;h�b�/������ғ��Q�-i� �[�i$&�;��`[�+��3����[���w;U�tfU��L�מ
���o������ݣ��&w���;�z�6�;%��~�������M�Y�Ǽ����Aպ�X���-�K��{���M���Mf>fД���ʕnf���!?���`��j:���A��q4[5���ŋ���f竕<��	���@E�q��p(~
=8��z��7¥i�f8Ƣ޷���OD�*��;�����f<{m�[�=:���������4���sn%�ǽK�y;{Vk��S����֝l�x�c�㵙��Q,��a`��(٭3Z�����Wr�|.�x�d�ca��&���v��Y�\o݈Pн���y�d���T7��Z��lR��f���Q6��m>svEl���b���y�Fa�ތ�}ӵμ_EV��3*���������՗!�w�7ӄ�����J�Y`g_GM*�7��<ޥ�Mƪ�-�$�A�t�/X:wH>�W��qH��p�{Z�f�W��ͣ9��NѲz*b�T��A��n��ʇ�J�u��NfKNv]m���ub�G�U����d�����2U�� P�s?S,����'H����y\�O30��(�R��$�0�����+R��c���p�s����k�C��+�ޑ�T��~$�:'�m0!�R;A��;�a��[�91�|�z�ﲪ���2�y�r�U�nji�����P�;�t�s54L`*��d�Ů�h���q�T.��L�S̱l��÷2��go��zV��O�-�T=n��o{�쳼-o��rg-fGD�Tݵ��|E�y#1������3{lTK��pWa�yߠ*FE�;o4�g|���a��sZ�.iu��������Q6:i暀@�(6�k冗��8�g9f��P����ly�fyv;äU��s&��m�ù@�,l�E�A�2�+��ݦwυ�;iz8�I���II7_���S߂���d����QK��玪�Js��3�>��<�2
�"��=[=Tz��JV�ל{ۼPz��<_s#������U��;yu�1���j��z2��Y.�}�8 �1�� 8���TA�u��S�0
b^�2y���Y������=�rn�CUۼDM��Ȃ���	��B»ճ�hI�5��ۚ��Jq���=�ݚ^����X��y԰����5{�a�d>O!-]i$g��3�y��o7���ٚq#y�d_��|�s���h������D:�b�I�A��e_��Dt�ws��C	5){�Z��q -�<
�
D��Ǭ'�w~<�#����"����4CC��ߴ���k�qw�������|�ɋ�$pN� ���g6���D��:��ٜ]7��1�"�,x��Cn]�c�fm38���E���`5�1+.���o��q��C��ȶ)�[��ՇK�wj�jaL������V-�e��=yo��I>��iɨ�{�f��t�c�s�\��������Ko��e�1�Y�V�QO��,=띪�:�b{p���Ovϓ��{�*�YB���χ�r�[]��
�1��o��#���+1e{p�&��l�>Ƃ�/��W�$[Ǽ����S�+��2Ĳ�D�7����!V��
[������s"��k�DKf�\[جi�
Yצ�B�ֶ���Z�ܣbW�1�ٙ�5׷s4R'C��_kNd�\��R�8�1P��5^jS������fv�t�w�:���dؔ�s�� {��\�\�f&e�<��H����������ϲ�Ү��?Rn�?�Wݬ__zM-R��F�m'HI��S{]B�o6��#�k�GI�R�UN_�a[@�x����b��9���b���<[����븘&O��ɽ��$g\{% ��!���8��:|}W(�-��]�lf<~J���-�܍���:j��p�`k�|�����.���9z]sS ��p�y����ćv�,����]�)�I]1�`�f�t0Y����vϖ��w=:ݞy\�U�W��tϭv�l�xз�YUM���m1�	����-sy�o�7�t�EQR���9;K��#\BM�B7��i��g�}b2�qԦ]t^��p'�{��hӉ}Uf�n���잗1n�O�W�>�S?�,�q��2#v""};�N/y`��K{#g���N��su�zk��]��ߴY�u�}vL{5�#/+�S��\9���K����5�;d�����D�xh���P�Ui�!��l
<xU�z'���'��c�9vvJ�����k��jù�i��K{�M�!��ZVR��ݡA^�K/A����)z�~Z�<��3Gw��o"n�s�Dyy��o7��gi���D��0�v)�,`h'�T�S��2E{|��R�S�s��U~�Te�5r���/��ҽݜ\�~��U���H{!S�e�!9��.y�-�ݙ�m7�
���{�v![��ؕ���ͥ�L�3��f�xê���q�f8pF�{���nu���(2OZ���<҇(l���᮫F^�7뎰A��
��s��׏�G���z�(���D[y���n;U�wa�v�O�$߲�x�~���� Q�7]UuW���gU���D�%%<�Q�u����%/_*�O��7�3z���+�0�fR�ܸ׵礞]@�c���Q�����=��ת����B�A��k�iII�k��J���xm�Ѝ�\4Nե��v��	_�Ϯzv�D����W��]����IsP�"ⱺ&6.�S�KY|ń�#}�ԫ��y
.��Q�u�9��5�S+��X�v�G�Jys^�]�|�
,����(��)�Ӂy�_+Vow�r�T��Ï:��%�vq�u�l�nf��F��s=�)HFG��m�l��s�<<<<< ��3�9[f�8��>�}��a�@u��B�z�n�I���X亵��h��5��/cwv��%�T����f�\�"GOe�o,�n[{C����U��G�]�������#��_%��X~��I{�5&�|W��T�?���r�������j����9Xιs������L�h�N�离�sN�a��a�9�9���m���� ����s��Ͳ��M���.x,Z'Xs��JTf������ƿ��L�W�񷆝"Q�;W�d�����X�*���S�OI5�|C%\"����]к������Tz����s�����<X+�0:�L]�>�t�r��J^��TU�����&=��lDZ�\{X�KÜx���L^��w�IqYd�Tcz�nb���4�kҥ�m�iR�ɨ<���t��5 zk�̺9^�L*�\ʎ�_�n�W]�;�h�A�v�[)�]�w�{u�A��0Cɪ[J]+��j�����l�G:��38�1����YM�����L�^42���������y2;<�X-�OM5��Gx�f�Lj��NʶO��<<<<< �'w����.����iwr��
*|�*�����\*�5����3���G�}�Tƈ�Z���+�ͤ�m�R'|�[$�6RRp�������H����L�C���	�>��[<���Y������5���L�t|���Z� b�"n��Q��Fk��2c���Y'&��L���<_ި���_B�5+��«�<��v>���!]'��}���������%~�A�gԦ�+�b]�w�ݢ��^��;�r���gT?��JC���7�ex��V%t.����`g��)�h��F�cF��}����ͮD�R/J�c��{ǳ��ݻ�ɠ�]�w�= TFOg k1y��C��}׸ #)�u��{�c�u�$Ⱦ�3�w5}��hpn�*��G���Ƀ-o�
�ͣ�8ujq��ް�{Ӿb�(��Ħ@����#��ge�'���/�R��(��F���}�e��c�Ӻ�%�]1>��z�}��`
�z;*�B-�N�b�r�^�,Z������!Jjz$2��|u-�V�2��isɖ���-ӎ3�=������«ZO/���*\���G��Jے(����,X�r���#�TNG�x���{+��
cTF�����zI⣬^{R53Ë����~�h�p�i�b�kѧ9��U07C�V�p^��{�)���GoQ=k�6P�o E��ۮ���̀Oa����<1���UC����;gM�4���e_+�X���o��ck���K�vL�jw$�r���Ch��<@w�8;�b�b������GH�JW�<���f��,����Yܭ��M��St	�@W%7�C�����=�������j�zf�J�`o�~���k�Z���D|����M�5�#P�x�s�^�k��2����ǋV�qͰS��p�>��2�#�r��.�/���FYO�+Sa<>���y���u�ܡl[P�U
�q���{\�uc8L�Lb�����7�7�wd] ǩ㱹q����/[���ـ���u��ѣ�狴�W1��:#a��EM�y�i�g��:�Z�L�Q�ѭ8J+�T6ւD���k����R�}G��M�jS�VD��R6�#B�u$%v"PJV�F�j�U:�KJ8(N�K����t��˹�I���1��sھg9ޕʿ��w]�o�>w`�K��Q	����m9a�,g3�SW� ��Փ��6&�]02���m�d���s0���o6m��ə���g�>�0��Dp]��%�!��B[��ɯ'��7웺-���Ɲ�~�����{�D41���E1#�C��zy��ݲwr����j�A0��צ}V3R��pi�&��<��@"���W���'-��d���Wv������v�hnuDi��Uѝ�~���ޗ���X��^��:jdD�?paG�5�pW��g���owg�{ܢ�������T�rZ���,������ �ȫ�B�� ���>�k&.n�G 0���py��;�>�a�Qݟ\��
��P� ��b���a<�WY�;kr�m��]��r�F�u�*��G�'7>���=��>d$-b�kWYT���b;ј�HE�.�rŌn��c^cx"p!*Ȗfp�G-f����(^�+��X�khZT�������e�#@4����l�2T�olei�(��9�-`ʛ���SɃ؊[�Eϭr�27�zo$��4f�xt�f��ͨ����7��i�7�+���C�>��9W%Z�1Fi�N}��-S�26���"�G����z�J1�NZ.V�'���]��|��t��x����:���[2���zV�+(��ʂ�d���&i,f��.��.�-����w(��PZO3���\vZE�3U��J}��+PB���hP�h<X�'�;w�j��9�>/8��U�Ή�7:��,Zv�v����xVVVeG��xu��;ܼ��pɪ�/;U�E�!��{bm�fg�&ֻjY�;:r$]��\�V��3��Joh�dֵ7R�Y6PY���;d]�����귣E<�$7c�2Dּ��X�Fk�N����
��F�;2�X��e̤
�o9R���z�V�]q-l��L3�*q��|��۵����G���^����m^���:��/�R��K�.�a`[��w����ꡔE��#�-��k�:u�S�FX�w6���Y��'d�B- U���f�y��܂�L50�UN���V�Bs��Ye�wV-(; 2���]�!��^U�B�e���G˺��4.�ys]�5j��8=.!�Nk#G��[��y[��*Q;�A�h����^�uϮ�MC3��JU�>���� *p!q�sAS�ki��<KM�ۥ�uJѲ���4�n0��Ƌd����y�jft�he+Ạzt]RiK�aX�F���u4�fq�]�i����n��ųl�}�51*�)k���.��霭�����sj!�mlm�v�4���u�Ұ�VpĄ(i�\���a�X�Hr�wd�ݳ���yYm���i����73�i��U�w��&�)ѽ�W�ݖ�~̊Du�t3���"����w�t�H[@%ߖ�Ghc�pm�E�sZ[�yow)���p��9-
�nU���'��y�����A��%)��[R!t�޼K�Jb[��;e�]���:�Xҋs�kqv���_Z����r֗�kB�b�qjw.U�sT�ݗ��,
������JX����F�OZOF��{�"����1�5�nηyZ�S}�<��q��۫*�[�օ��P�[�%��L,ǖ��SqJ3�&ʀ�Ӕ�QPkn�J/o��,����/�� �[�]�����[���RMʄRە2��<��oRu�c%�h�g�᠖t����ww
�o�6����ݴX6���=Pq�}p��R\�I��h���{y�Flғ:�Ke:��ź�hbd3N�ԓ{Z&����7�nv�� �$�N ����#㮑1"1�Oh�Ԅ!!UT*}��i���׮ݻv���v���:$dʨLIB���vκ����/I!�j:t���}z�۷nݿ����%��`�� LC��|�r�y}����=:�$�N`�Q	!!R�!#�o�����n����;�~���w��$4b����"��nDf"E��ƹ�������o{�|}z�۷nݾ���H�	Gʹ
 �#�	*O��%����dtO��^.�np��FfQ`�R ���s�k�"�u��n�;�z��
'��P|�R$RĈ�dn�]|wG���p�f���^'t��s|������K�/A�ҹ���hO}n�.p�.����뜏:���a�{���Fn�����%�4X��s |uؔ��"�0�����=����eL�h�sY��&v���j��)�/N����-AN�*2� ��yml��Sxu������Ǉ������LN�~��l��|���㤸T���Wo5��i���v�%������\���#���ؓGԯ�ˍp'���o��G#-޽��i�n��Djkף=�M���g��S��"m:�K�H�T�v���[-dE��_�/mW�\���L֭z��������V�9n���v�%��S�i��yt3�{��v��h9��}=I*O3���N�;�
�t��\8�.j`���{L�<���󂌈ہFQEc��سS��."ާ�	���o#�{ ϱ�v�n�w�93�y�_��F�4FV����My�!�����ka���g�9�.�b:�/�B���T�w�֨#�X6�~����ey�}�poA�o7'ć{E�b�Y�/�a_7��p���.*��B�X��J��W�W]7`�H��'�=��̉<%�fj�cq�"&��_�
���a����nzi�9R�]"t��8����ќ���5�k�]jZp�YG���hg���etD*�mn�AE]\��m����}��7�3������˭΢���G��.m`�&m�O�����y��dV�q���N�W� c�>�y|�us5N�,0b{����S.�W\��Sy����n���X/�Z�k�8fu�zvJg�ֲ�{��8�t��^��M�j'����D��,�+��!��#eyz���O���� T�e�e{��VdЃʀ���:o�maԒ}Ε�pz2�3����M���'<hA>mĄ���9�U�S�n��a眽�[һ���%»��鹿P+x@�{Ȧ`�.��JW���g􄉥[�������6ݭG,%j�I>���F��ܮXT=���;�y�v����j���1U�,�;ݪ[��Al�0�i@� �.�]cdb�e�u�b�T��Ez���4���s﷫�L�o<�yPޖp:�!��,�V�P-��l�ͷ���:d����nq��oT��+vA���϶���m�ǲ� [xcw��	�C$$�aLV��^�Z(p)�rkέǆ�m2�'!n;Z�=��F�Zz�fH1We���#*n!�\�M�7�%2�W��P�p��dS�Z�^*�v�ǫ��h�ֺ��l��:��K��,��3-���fd�VKX+/��@���c,tl��Ww���[��}tF	�}����M��Et����������-�D⅕���ΝY^'��]�S}[�����V_:0�y��I�a2AL�c�ܣ�ת<������U�}�\��)ś�{��o����(���?��/�Q^�q[�f��P�M�(��&Rm�)w{e�ʢ~��Cz�xTj*����.*��<"������P�U���^�}T;����C�~�!>3(eC�SSՂ,�k��� G�"��'{�ɒ3�u4�Z��,�6}l������� ��ZC�FU�C����60+,v�R�2	�i�@��s;-��U>�n��T,��;�تd���6�s���*��poֱQ�խ�ˑ{-��n�ma��`��y[?�ۏ�._���"mH�:��	W!����"�.6�n�N9�n�I�}���[�ճ�Wv:�N��	>�+�������pƕ]7KV<-���n� �^���APW���n�ѱ��fTl�'� �9�4W�ʾLQ�D�uzp�ֻk���Q��x���/��L�x���	��ݧ��pN�W�̆>��RP��ܳ�Pt!0oX�5*	��ʹp��uZ��-�ݿ��_��������
���b���f�7�I*�����H��P���W'��EK)ɼc͗�{$�Q�}�i4��y2v�m�-���L1�%m�G��.m��<�UB���5����oR�e���B9���xj�tN�T��<[{[�n�q�˽�/I���
�G��Y]&�<�x���E���-�'�9G�S��NшY�d�丣>5=�S�c��3u�Q]c��8�w=k���:�0j2 m���gz�����F��NR�
j��M&�L�}��;���(J��2�t߁�Y�*��q�<�J{�1�{_DG@��<��i�-�E�1��#�S^�h31.�$A`�*��s]|k]���z5�H͟ŏM��ȧϳ������=,kg_����p�����F�-<�s�xzB6D��*��ا�mX̣��V�_�[ͷO
&&��ܧ��!I\�]Ar�\�N�z���}o�^j{�t��:���A��j�hU �{�.K�Jv��F�E���j��SV�N��g9�Nppt+Wf2�^���oꮒ1�Od}��C߼<+��¨z�ogsv��`�����z�욋����Xd"{֟R:�2"��(qx-���1�;��]�-�t��W�{�VN��.!f}���[�)���l���d��'�[v|��o2( �E��3k��d�VU�K��D�|)5��E %[��ӷs�{4���-�?n_�u' ݴ�|�p���eh�ӯ��6�ו�)*c6n��������rЖU����Zch���:�}z�z�,�yʕD���"��(6c��3�L�хw���NL��+�Ź�M��~���y�}*��Se��蚍۝x]�H�������6@k}���L�-w+qz�lyN>�Th2V=t�R��S"��O�Ľ��*��O�X�1��zժO-5�q�aUQ訣��
t�/vV�b׵��g�fԇ����/3qU��}/wI�� |�8t�IS�z���Z�G�q\YȾ碲�<^AEG��5M�����0r��z�e�/�sA�'�0)ʖ5���8t���7���l���	ƺF;�3ٕ]�.8�4���S�_"�ԳB׿�
���y��k��kf����n�	�W:�E|�}}�=�ފ���+>G���o�{t��:����j�>�o�>w�jv�_%d*�ɮ�a~�t���R*a�D�c	�>V:En^l��27��p��p�"�TUW��o��F^����5�)�Fq��8�<�{�/��1��R#�C�v�1���AJ���d��a��eϷ|�����F�Ů�VN�6���XG����=zÚ
ϖ���/�պ�����:��<בj�%3;��$]�v�gKՓkp�!Y��{ZOmV@����D�b�����>�֩��Y��wR�����d+2hA�TU�K�c6o"��6�v�y�8�����R�j�*M��ݣ��kʠ�����=��=�vi| &m���O$��|F���"�cc̫H��V9Z7��MZ�3T<��=[�V5W��e�Iњ�);Z�$�C�9����tkt �����w��5W�g��+T�S���}X�V���"W�qw;�k:�"^]��MýD���p,������zݻ�Ջ��-��Ju)���]o�xxxxxxy���~�u�7-yu�N�M8��*�L��v�d�5�SwF8g�qv�o/1�*]X\�X,e��2<�)��sϫg�U�ó�\�4-z�˽��e��?q�����^��,�M�#��y���673��Is[ܵY<��4����P���k�V���G�>��9��O����C8��%�*�4���*�:Y��?��q��, �3�u<xl7Pm`���y�)��FqXJ�5R�����*�n!�]j9�a��xX[R�?�(h���5�<�[Uxn��yE���V<<ֽ����Dx8rC����M����Eda�
t5���U��\7HSϗ�LG�(�0�U,��6-�����;�Z�/F��M��cjx�G��%��EsC��`;�U���X�sQ����::	=������S����]__�H�nU��jB53�{p�p=2]�W<k�N_ɬ���������r��{:俣"�@6�란��J��(̷�)�$�.���vJkmm�
�J���y�����(h��K�+ͮ���Duof������;)�.���N�Zk��xxxxxx{��枞-n�- �N�9�����|�o�{o,Ϯ��i*�m��暽Ŵ��3�Y����ظ*��R�j�mX�l՝�p�m�=�h�Љ)�{�qA�ڀ{VPt`>̵#�Б�}Ռ*m��j��_��z�|s4-����<u~G*��Q��|��7�)�Y�3;,�F&zA$�X��\��u>�
���}KeZ�v��رoa#*Gf������"�\u��Kv}�}!����&��6B��Q<S�y=��\y�X�"��V��U��^��t<���t�-���@J�F������A�����L	�f�rm+wA�êt��K:�u2������0Y�{�!��t{z��4�!k�8x�`Wr�~��Y�2N�dVt��L<=j�㧎�=5OØ!���>A�jQ�k�~�M|��e�FL�"�pڕN�޼��>��ڙ�w�j��`ШkF�P�Hn�]�p�HwT̖�JZy��H�!�CZ
��j}в_ČI��U���s;��v.��[g���C�7{un���γh�T���3!l!V�&2G}?G�E9K���xdE�<ޅ8�R��+`6Vko�p]�Ȁ��Ղ}s{9���Iܖ]���}�g��-=�m�Mc��D������;k=��oY:
��-�ڄI��Y�{�	�H��H��&r�`d6�y�SU����}�{z^	��I\LvK�҉�j�9�+j�T���
�,�K�3�`�@@ߠ=�h���ϡa;������c�;wqR�{kz������U���v�$'���QJ�U�\�0o����S�{;v�w�|�@��#{o|��9V���0l����󜀭\L�x�b+�j�}
���
H�<�|���;.��ĵ�]9�B�c`��݇�m�J`E���k��w�u��R8����tdC*��(�ܭ�2��8����)\q�W�J�h�� 3���^����U�[�|R�2�ʜ��y�N;���#��j1�{�"u�ÃȻXz�6�wn>Ü"�h��&��b�V*�����
�-�ի��ф��;�t��ju�7�-���h�ٓc��Ρ��[OD���[�xY�.����m�n�6E9�Mco�S2�X�R̫r�����WՌ'�����S#��`h�Cܪ[����?81	$R�����}�e��QJ�y�?���*�`��� �t�	γ�E�^�x-۝�E��wLAJO�}������o��y�0�([]��w���,J�f���L���9y6���:'a�YP�W�9^ذwףG�;��H�ט�	;������ǎ���:_��u�^���y�b�d�~�A����|-���w���1��~4	�	Bv���^l���ƪ5LX��5���\�{��ZvRn�B3ꕒ�3�]�]zde��|v���݄p�*ڑx�����Ks8��]�iP�ۛ����$��Dԙl;g�m�@z�������?ҿ��Ҡ�*��E���� ��#�QE?��J#��_�*ܬ�Ҳ�+5���Jʬ�֥em1�V���iY��ljmic53U�1��VmYbʬɌe����S,ڳQ�[,c-YXƦ��I������śm5&kY�Kk5�ٌ���Y32�L��ki�,f���e����5�����K&V��U��1f��5-Y�c5�c2ͭ+&1����S6��1��Y,�l�Y�*�Re�5�RɌ���6�d�����1�kfL�ͭ1�Z��1f���VX�Uf1�fՕ������&[eejV5mҫ�-ef�5,��Y������T�e����Ե�f�,Y������5m������b�l���e��VU��������Vkee�����YY�����������VZ�Fj�ͬ����`���PȨ�(�P1@ 0T�Y�U+-�R�[U+5�)�@ 1@ *کY�����R�U�C@ 1@5� �D�YV�VV�J�Z�Y�M1 (�@b( �@`
�j�ij�eZ�Y�����R�kU+*�J�mT��U4H�5� �P���Ҳ�+6�VU�e���$ 5H4�@b����ҳkJͭ+5iY�Jb��&�� ��@b��Ҳ�+-iY�J��VjҳV��ݭ�f�����f�,�-��em+6���Ҳ�MJf�K��^�QG���T 	#E$`�~�Ͽ��V~��>�����������R?d�������P�ҫ��G�^��_�����������P*���1 U��?�l����ba����������Ch����>���4�
���8�����2į����yD��EU� )�F(��ԥZe�T��ʬZ��m��il�i�V�-id��R�*�@H�4�iZU��ZU6�ҫ5eZT�R�V�f֕-��5��V��kM��*mi����ZҪj�eZjU���MJ��-YU6��H1��D�AR,T ,"�,"$#�Y��i�֛+ef��l�d��6�6�TՍ�Zʚحc[3Vi[&���k)Z�m�mcV6���idQ�PBAAO� 
�T$QYb�Z*�V�kF��i�RD #H��BP�_��?�1PFE�@	@g�p
���������������?3?wࠀ*�~���_�~��?���g�a�0����a��,�_�� ���(~������� ��  
����!�UUk�?X���F�]� ���)A�v��z6�f�v��/S�G���, �A U����~��� ��Ci �^����}�����@�?����( 
�����]  
�������'�^��ad��(8�ƃ��������&�� 
�'�H���֔��������6�~&u~���/I�O�*�"�������?���!����(+$�k#�  ���0
 ��d��G�|w��*AT
��*��	Q 
R�RTU(�E%TU*�)D�UQ�	(�ARJ�RB%	!@U T*��"�{5ER"�B�
D
U)�BAI BRBH�P@��TR�P��"�$��ى@-�j����UUB)$�*��$R�J�*��
TD�AT�J�$�B�T�T�(�UE@@�U*��ϬU*UBJ� ԽB���L4�SMkb���Kj4�L��MSR��R�%�5H�h�em�wh:6�eiZ+VDæ�iJe2��vԥv�P�!*U	%J)B� n�CС��t4-�z=
-� л��(P�B����VM�ֆ��Q�Ɣ3�*W`(#;��-����wuJ��Zwt҂�a��WJhV�JEUJ
%UT��ER�  � �m���ڔ*���l�Ҧ�jb��l26ţ���f�)[jR�Ri�L�V�Am@zܫH��Jk4`�h)	Vت�IJ+� � CY!*��C  ��^�����mP��T��� �J	��5�J�&hdRII%U�)"Tt�� 7�(Ҩ�`5�Ѓ`PT �-j�`=:�P*�N�bZ5F���أ[(�
4�UUIDQT��"���  ��U ٤�(���� 5���v:���(�h4[��i�vj��b�V55�rT㒥��BD��U@Wx  ^UE^�;��(��IRTL:������:�$�ZwU[���B�lp4R�qp�HT��4�R�s��B�.�1R*
�$R�  3=�Q
$��㊔�p�r�T��NwER�B7JgQD%S���u��E(�:-�RHT�v��%-j�ΫJ�L�9�H��
"��T<  =�*(P�r΂֔HܫqR6ĕi��UJn�w ���7�U�Ηt��@0ᡄ��[��A��!GuU:a*U%UQRU�� zPI�K�#[��蒪�V��m$��r�
��q��)@�Φ�%J��)����@E�ԡ)Jx)���P��S�0���4  *~2����O��E ��{M&�T� ��F�	=T�LUI��16���Ř���f�#5�AB��w�2�J[��ί޺�z���s��߮uu�;kZ�ۿ<����kZ��޵UV��-��km����km��kZ��mUU���{�����R���ʼ�y��+���Q۷*4.����5��r��4��SDeR@	��nZ��:���$��E�A��e���0�u36�e��A&$
�r�au#��X���j�i5�n�����w3w$46�<�8����2����
�{7�Fs�2�)D���)̒���
����f�R�2�ն�ZЙ�p(�1;ҥ�B��rM��P�pk��,���ռ&�b���J�5�A���~©����!�Q~U�N�EN��N�����0�o�j(t�Z~R� CM��iǁ��(��l�Y�n�:����-6b�L�k��V��%���wL"�ld�����+^"�T8�&K��`���T��jٺܷ�F2Q�]�/E�ì�aw�6��kbh�V������r:��e�yI�ni���� !^6�[zh�GoZ�i�c������q2%bi3u�[�r���$����6��eJ�"�t>�S-H��X/*pX�g2�]�usT֛R�(aMʹk5�U+�����6|��sn�ࣖⲘ���'q��(�p62��Т��)Ů��ze�kn��S*�YXi��鍾���R���(���M��]E2h�,P!8 V�I���Tx����F����~1��h0�T�*�g) L���I0ϯ Cvq&a��P��[q����Z�I��b��r�ӑ���V+2
��f]�*����C[@�&؎
����w���'��mT-�[�5���R̼�61�O�)ōѦ㫲�Y���a*�Ւm;��2�ڂCz�U���ո��*ڽgf�-����ӳa����p%�+E�i��-M���m�7����Z;����!�����Zpkذ�v�fՅ&*�Uὰ�̔� /J�]m�b�t�-gu�4���{�weJav�f���7z�:�+�5Zb|:�[wz�B�d�Z/1V�+��3F+��r�����Dp�/Ũ|fؔ%�bT��X,���q%�{����/M��i�5�L�g]*�aȁLV8��ڧ�Ɇ%k�y��o�mG��v2�ݖ��,j2�XF�1z�Ō/��(S��
���5Ù�uj�'�j�5{�+��,�!�v��P��%M:/T�(�0�hd3u][ٵ�G��Z!:M%��w�)��6��P���c*����L�R�da�lN�u�m�.n`�Zӧ�X�`
����@4���-��Kp������9.%��91cyF[�.�LU��;�&d˱�Gj����92S���1G&� �*�ǔ�J��v(2��3GF�4�f���i[r�쥦ږ�#0!��d��u���󥶄���Q7Z���"�[X]�4Ӳ�e�e�ɒu��8�u�&ԁ�c�"M��lg�]��3,�e^�z#x�#��0혲�b��iLH:U71�ef�L�%mf=���PJu�������*̌@koAU�CM��qm�Ӊ���Yc^7��s��`J��&�^��Z�xkB��J� r ��@i��VbZ(y1��&`��7�E'Gue��xe�x�ͽ+sH��ҏ*i7�j�d�A�i���- ��ҡ�O���5M��QD�y�l��y0�p�w�t''K"�$NK�%�'w&e�`��m��,�6�&�,� �m�_���9���B�ߍ虻�HLɱ�a��n
�~R7�,�y�D��[����jPS;F��N�ZUaג��`�w�E���c�^'���ٹqV�m၌waHf���S�v�m�� �Q��tuJ@�D�����{����gDq��r�۰m*�����h�y��b�a	:˔7,�\�P�M�q:�+��)ҡ[*��5 ������xi�[f�DE�A�r�Z�nJu��R��V-(Q�Vi�[��">�*M�]�XE���)Sg\{�a��s4Ĳ�n�6��^�ڡ4�G���7CnӳE42�<z�nI5:05d
��i�M�dʻeՕZ�U�e�V���ƞd�H���XwY.�иv�VX��i\�vF"�Y�"���KVa���T�]��qQZ^d��E)�n}n7��廒VE�e��`ۭ���ٮ�u1�b�Z�6A�Yz��6H��Fm�7��K��.�$Z������Ka�����ؙ�EM��p4v���IYce�%�Li��3$+76<�	�B�E��%��+�W��-����C\���f$�X�CMni���i`Ê��W�7$7.Zc�`jOi}l��AMe�qIj�b�2*ko$��0݂��ܦ~6wjQ��٦L4�O�ܓ[u��	JIW7B����-Oh޻�W�����ٛL\Ö+E�z����r}���dFi�T��b`n��ɔ�ށ.�z	�Vn�[)2�hѳHeYR
�uK�X�zu��{�i,�(;�V�Iz��06mۄm�{�J�cm%2�X��F]���jG��r�*7VܼyH�zTW�=��$L1�`X���؝�n����r��,A�i�F�a^�gn^�2ΖP�׆5t�R��VLUO&���t6�T�t��ҺW�V��j��-kb;�!T�i+�F�eM4�E��1�H�i5�V8&5r��=P޽E�o.���y7v��E^�i�q��&�̲��^�)#N\+&�$�Z9��T�7��!f���!P^�D����F3�A��L�ɖ�q�مK�֑�sZw��
�K,lK1#J��.:5cAn�(^�1]ܖ��
��t�J� 2D��H\q\,��v�дD���D;)1��W�	����[��Ȗ�Q˻�6�aZRhN
u����qAR'�dʕ��B:H+�������ND�MKvK�h蛠0ji�[A�b�]=�1�r�b���̬x^�&�Z�i�.¨�)��i�)�5���^|�M��w���l�X.�T�e��������1)����LV�ܶ��"ZE���%2�D�Z����Y�tCNU���)�MY����:K%k�d�e%�1R�e�N�Y7v��x��u�ta%�4�����̸X�fJ���Yn��('2����u�>�/Z�%��4[�F@�Yh�tܷ������̍j�V0�Of �m��$+N�X�j���V�5q�G!�2W�$�b��و}`4>��͇4쫬��	��Ub(�6c���ҽ35M��U�����:\D���+-�ַ4�)�� ,Q�Z 64j�u��ذ"*�x��N��Y�إ+%;Π1��)X�n�G*�K�����sT݅f�ˢ��.ق�<
�[�ñ�i���ƅ�{��^<�	]r'�V^���)�4��dJ�x�)�${�i�^�T��l�iTrV̐h�d���ov��$J�ּ'_�.��`'�m7R��4T��:��p��H�k`�R�����Z���,\�Q��j���$�X��[,�Y�ٳO;}S����i�[\+$�1�j��Z�ԋ�CFG����[��JS��Ø΀,�������e�o 0F��yB��11zj8+#�&�=�us]�b��L�
�c�E��q](8�6�\_e�z�$m�rmG���U��~Z���!�q�fea�Skt��o,h�p,vR��ݗ�n���l�i�uj�n�CwN&(��;�~Ɏ$4��Z��VR�)��j�ɫ)%��� N��4ܙ��ڇ0;
��Sh�N�>n����Z��Q�x��rиK�v�e�o����'jA@�MIx�Z�c.��2�%�4�7+Zt�ˑ��\�+`A��8$;Xp�գX�Яnb9r�;���l60��̢h��&J�xV丆J��]�U��"Ao&QT���:��kF4)Ex��4�QN��9�b1�Z��aj�%���2�qSg2�P`�Z�u�pn_ʱ�u���tA*��t�*�ͺC�5Lej��-�uͤ%;��&�3 ��f�M!�,��j''�DU�J��dq���Jq�[��S���P���F��La0� �suaZ��M��jHSi�`;�P��y@3�B.��X[p2f-��o[��[�-�`
��iDԃ/4�5Y{6�=CWI[
����{�\�3S�!"2D��F�d�YZ�;�4�M2�a�T+Y�Ĭ�WDk����.�#$�ecE"�wu�:�YX��u��$��g����f�ԙ=p���H͕v�#�m}n^�m*�BM�2�f�oi�"@C��Q� J�*���x��cf�3D�.M�3F�,�D+BB<7Z�J�}�3i���0P�X��8L��b��A�F�A�~�X@��"ˍ�ull�ǬһYY�������J'��5*`[�mÄV���f��C��l�к�Mޫ�E?�r^�c	�#&�ݺ3-�\�N��4ĕ�^ ��cu�������A�$�����V�Q��խ�v�lU� 4e���n�4&U��z����! �A���:PKS�Mjt��*��K\Z���s�S�H��[U�`ժl�ˋ+]�r�w��f�f$u9�`N���l�6��y���&�dj6+>[��ѽj)�KOu�4�J�9<9�I��z�qP.��)鹁 [[�^�Q=6�'����r�&#J��-R�\9A�Ujo.dr��0���ݘm����5,с�]
ڇ� �4۶)�M=XيSIz0Y��Z�Ocоkr�׋	W$rS��fQ�꭬i��/�i��*�*%2Tj���m淒��Q���YnQ7���:�ʙ�����tё;��4s
&�r�H�k��nI�8 �h���z���'z5�R*�r�Le�Fɧ��X�xY@f��dK���V�sm�ۄb�L"9P1fT�J���{�d�FeѤ�VX�g�/��tm�۴u]���ZSU�b��5%=�Ǐs2�F�-����j�⫹�E�)�	�d��jyAS܍�V����X��lFK�ff��3,F�	Xf]a� ���r��b��pJ��d�q����1j � Zf�:��Yz4���N��O�����A����62�<ch��Lmb���&4!�Ǧ�k,��Y6�]�sT+IUQK9�ǲ��1�_��3^@H)�92�؍�%�u�� }j�(��7��66�M4I�����ĉ���+!N4�0�!��'N��Sw��bʽK��YAKl�)i�:u<nL�t����K�6\�o\�sY���][Z���w� ��nS��ц�3��0NC`	@V6��uF��x��ӹfͽ%���܇L�d���E-��^&�h�3V�G&���[2�ke���a"�gt��ZȔV�D#u���7Ih��j{���X���iw�MJ�vL�[���	�Hf�$N��L�X���zn�ӓ7j{��Z7�͒�*�3�������M�J�m�oe��S+6R��mQy5����An�m�b�� `�����[���lXq^J��!�4�7PQv�@h���#r��T�L�������\)�.X��w�V��\I=TM�c�u���-*�'t�+��,��l��* �uwq�(�3Y�!RmR�W�Ƚ��#kY$�ܳ2*8E� {���w)1�]LWzm�o�],�&�����K+-��.zi��6 n������dXQ�32XUV���y����H�������hjm�v��5CG!�p�-u��5f��;!�ݰ�毝6�ڦ�������(�aʒ��X�٠)��,?@����ͽ�F�
V��K��D]f���%sk(dQ���k����\
�m,d�y7J͎�mX��cjE\hV�}S#R��a0�'+u��A���7.ZQ�g��Yk0���٦[ց׵�w2`hED	��r'oFem��Ռ��E<����8���Z�t��r�p�6����Lh�gN#kjR!�aAY
���r�5!6�Y��f�.��YB�٘)T�D��2@�G(��hL��t��KhE�k �2�ٹM�"!�;K�����"�r:o\V�2���� �*��y�+pP��جT��gg�h-���!�72Q6����B� �Pܲ����ו1a�wZ���q3������e�q�l��[P(�cG[�q��om+��ԃ�M����'�ց !���@Ǹ �9xw2���{���
���wss)i6.�q��e���ū���fiH)I�Uf�u���$�5$��lR6�T"����/j�k(���4�Ys#Y���\�)�ҵ�L݇q=�zX��j�LR��E�ʲ[���Q{�v�H�)|�+�N�P�k��(������i��O $�ք�R�aK7�H�K�_d5gh"�(M�ʎͼ�k��@eM3Q��ax��Z��*�=V�Q[�9�#*���Ҡ+m���$Z2��`�+dk]�v�4�5��I�X��a��%�]���7yCv7n@Ag"��9�7Lw� ƕ\�����@2�f��Y�0S�c)!�6�lU��]C19�+�VN^FHTb�)����M���V��)i����P\�+
��ņ���Xd��de�����{P���:V�	��-��pm�CY3��X��\rSj�;c�1KwoF���E�*�6���VS��^�����Ad�ZyIS:f4J��ڶ2��*:A�v��j�C�)���e��Z�"S[��Х�i��3�����t#a�E�$Ӛc��*<�^	�/�Y-�!�{.;�u�RCQ��h���J���g) q�ʒR�U��9(�d䈑�=����2R�Zb�'���G��ۀf�EK���,Y�l�ef�s2����!��ڲݔ����$R��r�#{R�.��F�`-�J�v�EjU=鸷�[� r��jzu�@i���,<i'���\u���iR��zwg^�&��U�-�u�ү���`�\kx��D�A�k����)\�`�s�(i�(�ɵn���sl��Ɓ���ٴֹ���⮻�K0�����j�r���]P=]٦�?��:t
C�����p��O�v�K�i��ZU��ᰟa�N�hv���	�C7��ܓ��Wjl��	+�0�G��W_r�����m:���=-�u�(qMP߮�`�|跻9�����b�e	���J�v���xn�lg#�K�0.�	�e��uN�[j;X�CG�h��*�I��&�3p���frtr�h\����Q�R�����Wk�/%sG�%5z�՟���|�<a�הæo�p�@�A&Z�e��[��
Yc�� h�>$�Ŝ^c+��k�ӥ1���]�Z� 7Doa9�s1'�R�+/C͵N�+�CIL�Nb��X�f�|�u�1���p�Yx0l,͵���t�oi�i]��4u��֕�q_<I��ݯ=s5]� q�)��2�`��3�C�8�x���jmυ�U݅4��	1�	\����)*�f��uK��]���G���f:U0a��#�x��*u��1n^�ހ~o���f@Uf���)���n�t��{�6�A��Q"�1����^�Χz�΀f�%�R9�Ru�/���C�׃Ec���X����9i�ɭԩ@�gt��˩��ܑ����dTZ��HڳK�Uz�ij]�yH7��eҦȰ��h*���LoY��r�4������=+�t
�Q����2
�뱽]U{�k���ll[V��`��D�a��7]�D��pP�Y���ȸaHe�f��!ʅ�:� �6*_|�ɩ�����_R����U���h��%�t!�hc���]�~0�����4��ܛ\�E�8�^M���BD��MJ�h>ë���@�n�����;u�'L�T�+���e�éZ�
 ,�UHo	�&�R㙷����>zR�o�� ���#̀�4���Z��%ӡS��]�s'Jv�z��,M1�����} �+n�Y�	Nb�y�^l��V��+j���}��:��}f�E5"Q�;R���;��|�c"ɞsk��s��g^�T�����L�&��k	T\{�ǝ(�e�>�U�#�G'��Z����m����������k%Xy��@}}���t�Q��-Kpm�
`�i�;�c��F�JI.��1fJf��n�7lu��V��1�Uֺ�j����ːtj[��1��s�f�2��wC	���Y[&N�+{5��N]�
]l��5��~���X��GqcC�'�e	�]t�p��� �m"�t�Gi�w�=�ԖD/-ˎ���Ỡ}q �`P2m�[]B]<�k�@;L1w@G��f4�um奁�;+,�JE,k��s6i�f��ΗA�����g�J�cQ�%�8ttV_F����^��%�=-��*�9�5�}|��4-������	]ǨWN��Yҗ���t�1�S�z��U3@��'���R��hՔڦ2َ����0������(�S,0���Y�bP�;���+���e]�e�]��re��j���3��kV�\�D
�<�z��oX�]���Oq�2��+���>�W�f:Z3,c�s趭��郵9���攬��}k�J�0Ǯ�l���%A��cT�(�St_G��s	�=�&S��Rm+�>]O�X�Ľ�G��BL��vs��К|�WU�S�EAk��c�Z�5g��!��oj�5�>�'I���A�؜�q�����U����\�|��_jˈM(h���5����{^F�wq;*U�w��ڮ� �6��ٽ �Z��ݼV�n�f��_�QQglO#G���X�]l���`�C(7Q�}{��f;����<�f���D�uc=�X���s����*��=��e��.A�S8��G�l�ɳv
o��Ț�ӧV�K:�M�J�$w)�����Xޅ���jV�y��t�3w�m��O�%������ښEF�j}.��ʴƺ���Sc���J^	�
,���䲹dZ+��&�j��WV<�W��.�=b ���KH֚�y���ֺ�U�� ��lX:�ڏ]��9d7�N�z����)���m�o��M��p�x}�pF�{&�p����c�s:%��š�]A��e
W.�f��IZ���X�}*��o;�b��R������ "�ٽvU�����&;��=��Q����6�44m�-[K�Ag`��%�����÷��Vc����Ѣ����03�}u���e�&=S��L����CZ��\��*K����ĺ!3ٹ�z��O��v<JYt6��^;��J���T<������2�#��ۇ�VQ.�PV�c��S�yt���S���wC�9���e��O��k���!7J��0,՘�(M�}PEC����ue�q�6�4_l��sK��&�[j�.��J��Ŧ����V�����]I�F��z&��֢XJ�ضe�y�0�������e�Mkޛ���)�[���:�=t��e+e�u��"��,��ٖ�V�5dW�����) �����!�獼}�E_Z���B=i�R;�U�N�ea��*�M�C�bU:�H��WLYv8S�CՖ�T��e,A�g�_j�i$���]�����+9���֦`�ڿ�q�V������rw��<�ٕ��<o�*��l�޻�z�	�����Or4�^E�uۅ��h�ԫI@up-�xkJpďm��2�YS�"벀6.��3+m0dԤ(�����9���%�˺��wn�0�4�S���e��p�y�C%/rR[ʧl���|kGm[y\�J�7����6���
ʆ�.וֹuqWv����q%&ୱk�s�|9EUn)ȺVr�+!AI���2��,4y���ʩ�-��/25YJ��Ҥ':{FD��N��'4wZ5)|0%M��4t{yI�m9�76��դ�X�������7B�+q��Z崷NR
��_7*V˦���@��ͥ-+��y�lt��Q��Ӧ5�&Jtc9i7��&�ʹ���"yó��i��nTC����7��/T_S�۩��opfT\&cr��3��ڏ9�i[]��<�A�3K��$.�Eu�g�ֆ��z��sM*����j=˩�A{��i"��׈Ԝ0ur�$�
ۣ�"�\�+�n` m;�\x�|��D����Օ;:�e*vh�T:���uM6�9�U3�+�(��󑑓�Z1(�Y����[e�=��_FP'�L(d��W"N"]sr�(]�+PP����hN5�oMy��ɕ�pd��\�^olםVI�Ӽk�7ju��F����}������)�[�6�a̼��`�8j�5��X��I)��9�u<8�b�s��dN��K3���E'ܕ(��p�O��e$�A���s�q�*�74�-7�@;f*�OU����Y�F5�T�$g�i�3-fG�=�(�X���� ]�є@¶Rm�TY�fY��.e���]i��z�[gz8TУ�t����즯B;a�*��Ŭ�;���6�(��⍍���V\7ҥo�u��\غ�,����`̗Գ4�bt�&_�1<<g����wv�e$�����]������N�ҕ����if��o����7\�g.�s�U�	�o�e���-���ج�mm{�z��@J@nCa���[���75=9@a뺝2��*�ĝwu���W#���@�g�ѝ�7D){�M)b���s�m��;�k��!s|�R��W¹�4��\�ΣVG3�Rz�[;�Q���͎A�[�#��}\�^�ohA@�u�bWNGX�B���+�;��ɯ �$}u96��X�	����d��k����N�>ݭ�U&.[*�+��3�uI��b_F�//P���ք�n�O8�.v�G	t�Z���F��v8u%��z�����|)reζWf4�+�AՖޮÎi+��(U�%:��E'M*5��,@Fc��� 	�ל��}�>�h��k������y��813����6e���ҮU�Eb:�^MՇ{I�&G�0I��eDwl(��W&5wҴnKD���폩3i�T�&)0��l�K�geM����h�e]��}�nvr�mʅA\�{�������s]֯���au^��:F���o�b�*��-0�U��:.ޏ�;+�^�A�"�y��--I.������j@�l �V�l�nNkEro�{aACr.5�{Ő��/U-�l.����M�l"����������"V�2��%� <�Q�vo����+T���kk��oJv�"LR�uÑ�E0���
�{-��
���bl!�;}��ṹkw\�_9���nŁ�례��H��nZSnC����ϲ���Ǽ�Ұ;8;c��T�\Z��'6��������ל'M�ol�G�G)�kG.����\Ԅ z�����`�s/e`��=��wv�nv�".�+�%Zky�� cP�����J<��Ou��I��1>�e,�>ݾ��ح�4/��\����X���tk�;��R	�	g�A"��-Q�!>�k���	��
5ʠsW2t}�ڂ�KJ��{����+Gi������vHX�]�2iU X��%��6�	�jή�3����v0`�ĵ/��o/i�n�q�	�����ճ �˕��h�������X�ޞ��ne�2K�DD��q�~Że@r��c�Nu*o6mvAJ"��b�G�g]��n�۴M�o�*�Q�0tcP]i��W�M�s���^bhJ�V�A��
���{@�ӛHJj�����v���ۭ��
;�W�.�Kb�
Dv�1�a+Ds�o'W��꺚z6��;v�/u�F��]��=2�e�܂��������t+)n-�]�����K�Qvg�G_��4�=���G:��\�f�8�5�]��W�;�����x s9h��5�4���D��I�d�ԑ�;�b����'[�����V�`�%h������:�܃.Yqu����hj��8
E)U�t�o��A����S
_5S�1��g-�S��H�Vf�p�S�ـ�����֪�6�p�}��70�!)i;��g^�r�8Mv��*E��ح�1�ă��.��v3G"��n����LNer��sa��w�k';��~2���Y������3j�����%F�R�+&;���-�EwJ!3��{P+���S�8��q����Ǩ�ֶ��x��k��I�an�g�e�i�lzd<(.��^:��Dx�]3z���>l�7B��i]�Wr����b_N�T�T��p�	�>B���ksk"�xm���}��*� �bmC���Suf���:I�W�)z6V`�� 6F��Ց�B�.��yNr�B4�&��1KW>=:�Q�>�n�n{_���`b�>����$���є�rI
�mѝ�.O��q෭q�5��Y|Eu���@����|n�plb�.���o3':��*q��M� �&'vٙeh�л.��&
�Q.h�iw<�b�U��]��� �x�vZ�ˇ
�f8����c2]�xyޭZ�Vִ�`[t��q.a.����F��eM"�YBf
��T��[�p}�̈�԰��g�;)m�c3�8�OKPe��D5dA{1f_�ɬ�>��܋����}����2ARY=xn^�}�ȴ�i:8�����8ܚ:��e���U��pu��mhCe�6:��k6���n@�qϱ^
�{!A�:2�rĻ3�ys��-�fB���G�6�[I>�x����K�-4
��Ϲ'F� �Zr&F;ۧ#���A�ǯ���ԁL�Nne_e�끷��Y��r1���sH����8��)��w����_
�)�'/Yһ���5���� �7����]�[�Ew
��7��̂We�!�$8 �N|�X�����5+�egRO(Bn�Z'���FP �7�-����,�ѹMo=\2u��9�գ��E���:�f���:r-�0���ҡ!�u!w@�ueN�:V2g��w�+������op���}k�W�T��i���pf�\N�S�����hu*@�
�W�X�}W�����Y���rZ/n�{���jUO�uy�p�u���ԯV�1{��J��v9���SWi�H��4`�|�I���l�Y&g��H�/X�$lb-F��e�����%u�w�,���z:�-���:ձ��2V!5�̐���$s�����%���ˉ�A��)�Hm�ڒm+���e�Kr�+����A�ЊY3�=�h��Po��D렿�ˋ%�� KhM�
3:�jk�i��$��n��s��ߘ���&Bg� J�2�e�|�m��u%�n��u� �+�Q�#�
ㆵ�˝�R�7���e3��,c/�E7;o���ӀCu`�02R6!����J����il빨Ù�ۖ�ms0!2kX��H���Ө+�F�����`r�7;��&��g�7��jT��S@�����6c��'�n9���O�"�"�kA3���N�ʹ-DU�rJ�yW�o���w7��W{��J�+��M��6�C��0\̛�V��vV�&>xk�	�k	�Ն:��M��Ki��.�マ��P�[�ɾKt��][�g�%�&��3@�(\U��d]�na9{x�6������{�\��t7wJ\v�Etawo}f=��ov��[�d[�7{�_D�f�
ۦ��J�A�R��%�e.Y]�J㫸�YJ�BJ��0d�q�ň�*�L��I�j�������B�7�o��lȪ�����؇=��nm�ɮ�\f�޷K�����Vul`a�}p*w�i��қ��Ǚ��L�`�[��WB�Zɧ_Z�60g޳Ӗ'�g*X�.��`e���\��wwI�:��W���T�-�p-�Õ�3z����̬Qt��O��شg':���٭v��9;&�}�&�p	I��3�ʾ�����ﾯ�����������A���sg�z��U+w"���&��&cU�A8fwi��h9���M�Ɓv6�N�\�Y�+i�i�E:����+�E�Λᗁ�Ϯ�B�)�3��l�NL-2��#sMU���TnVM�[��r�)����b�Y*���wdK%�0*��GR}���+ܴh6�l�,���v���h2�lwf�}�u�Xw۷|��\��*�C�I��"��K�aKX��2�ޖ���o�i
>}�N�7�]��`	���<=�:��V\ޤ��s�g��.��Dl��?�)gQ}�PŻ��A���W-A:n�-r��U���.�� �w.
ƺ[��v�kR����t�����ף���U��^���w܄ G���b[��z�h3��r�A[�ti��}6$�0�fʄw oD���/��8�lҵf�J�?���H�]9a��c���	���K�3i��b�tU,��1�9����H�]ccW�GՃ^�	�ph��lP��P��������~�b ��EԢ(���jt���}����X7��ux��<�p
f
;:���Es�z�@n�YSil�/f�Ѧ~�������F ��2���0�+&I9#PU�]�E���}�H*�Z-�B�۷��Vu3�a��ũ���Q[ъ�r��J��O0_KK)�\�ڜ�'�mtƶ�e�7O�C�j�7�ɚɩN��ûW�#b�'i��Zn�+��ǆ��r��.�o�n���V�V��s����=�Y�dl�3�����N��=ޫ�X�t��%2��k^���Յ�e��G���ް�Z'!0d�k�.?!�ekN��$��b;���I1',�4Ta��׉�b6υe�G�;{�w�+;v:��ք�S�r=\�������k��u���qEXD@.\�n�]^�yȴ�ٗ�vu��z��h��؀l��#�W �m�N�wĻQ[t^�@ǲ����k��H�53��'�٘���T��:Ո-}��#�cu]Ft�;X�L�{QS�B��,p�x����>��F��pݻ!�@���� T�Ǫ�{z{1�J���b�6�e,���n�wu{θ���r�-�o���^K��YR{ِxk~��Mm7�o[����2��ʶ���e2����v�f���(:.Ъ]��K��7o49�ҟW��y���"N�s��1�)���_P��VvȎ�n�8@���/#�Ѧ�=YB�(��r�x�ul��Z�e�������nʽ�7�xk�B�1�f���s^:�����B�XxG,��%�y[v����Fо]��j���4S;-j�ԃ�h8ƅ�z]��D��񼫝�j��M(M���O]�u1_=5�:��f�V>���f��q�����*���6�=��=W��6�-/���݂K�.Cδ_J������p:��ov�Ğʰ3i�h��]��GfS .��:�6�k�v;��H��y� ae�C����T���	�2:��;)�@L��[�}ǹ�Fej�Gx)Z��Ae���j��ei�s]�˰��%J^��r6@��v�*��:�|k�WQ}G'9k&�3op-eP�:k�W��%�mC[%e�C�9���qu:s�o�v4�m𷗄l��}|��rJ&N<���ҖQ�`�;����3�
�o�K��P$�͢RV�V�8��(\�ֲ��im>8��5���c\]�S�\+�N����GfY�+
u�o_3J�-#oq<��ڨR���BG��U��o�Z�%��Mj��#D�ʹV"��$�pj���ÊH
(�N�Ց}�P�ZYWU����J}��̨�J�jԻ/Fh�;>K����ˊ��
K���4�Y��e�i96���9[�09�=f����v�Q�8�������ة�q���m���.������+4�yfSKyD2��AGf]��o�����\�GuM���k -`��r�G6�'!���l��r��$/4� [�L�Ǳ;ۄ=�Dp8XUtɶؼ�99q��d�T�^���,�2q_-�P7(����t߱D7��o���eZ�9��Ճ���ޢw�ק��Tѳ��0ER�����@��&�F�դ�8�v҇B�y]�:�\V}����(��l�ҩ�.\e���H�\�ly\�v���a1�h��3>J;ٶB �b�A���V�X�~1�J'Ո�j���BeJ��D�[�`�QQ���7ق�8+N���[8#�Ss�͝�<i��N�^l�{:����s5ۂB^	�HYqK.���R�WKK�ph��».D�wg!5붻��U��D�q��KK�|.�-�C�[�(9ս�8���F�<s���{��"Ug!�qZ�rȦ��8���v��ٴ���2��f���v!� ����;�b���݅�ᮗ@�bub�ӪY�Պ떣��t{�i���_p�AH+���`6A��;I!a��J�s���p�9�Bnd��5F�$VR[��-���)c@���A�L��;wD>Ď�c�5_
W�V#�����OH1���	V���J��t*�E�&J �y��v�+�g�e���t�=���w���v����Mc��w5=wyL�O���A���U���\��: WS�@�4u�p *�6`wObcs��wW�-;��ڛ��6�:�Zw��bO����B�Z��	T�L��_^=R_tlln�cXxn�m�kG
����Y�&4�+�j��;&u�������Lw�^Q�m�닠����`�^�6<���^s���Mr5�:��u��*�Ax+[�؃D{�ַ����F�;{$�kQ�69�!�" ������7��i�4�X��m��ĳ�u���nL�v��vƲ
�ݫ�2S+%�-�����Lb�sv�&��:���&4/ftz�q�{,C:Ýz��2L�{VwEi��G]Jt����k=K^��`����t��xY�l8�m��xC�
�]�b��0-�	Z�t��rU̫������E3�ju\(���
����b��T�eV���v����7�GZ��I��닽��*�=Jp��h�ɧB��#O5��%������t��dޟ@�|p\Kպ+����a�`X�{���K6NE���eeBV�ػy.�����&m;2�#��j��n��_f ����q���-[vmɭl{Ձ�[\��A��Y�#�(3��|��m���X��
ز'P����JzC\�>�wh�P�1"�!�X����LP�`B�o%���rU��!��;<}����j\�nɸ�2ښ�j�,��wV�:[Ő򍩩���ʔ�Z�Ve�9���#��X�	�Kt���nw3�12��JӜ2���uN�3�u1״L#�iœ`ڴ���Z55S$�-iU�6�s��$��C,*I�p��rnt�E�^�h������\���ǲ>��n&J-6��>XX�z�c}�|E�n��YZ�%|o�=��,y9Lڎ�w]�ty+ۓ{pG�WuoJ��x���s9Xo �\��6�]��1��J���4j������ d��&�n���20��^>��a�t���r�V�%�m����L9.��iR�� ��rg����l^��e,tK�4C�]��
Ƥ�b�5ۙ� �-��A�fq��2+�XZ�]k5ٌ��+I��M�\ěAmr�u!�[�*wjK�49,���ǪS�@+:��W.���)ûF�g�m�>���^��5�2��/��mjXNh � ��J�<��r�$\�ㇻ�z�T��lQ̷�fk;ږm�=�Cu�]tk1�6��דS�O��kEJw�m���L�z֍o�l�)� ��d�1�!R��������_[����
�@_Ѥ���a{�`��,�i.�c	�ZX��G��\��o/���#2�\ژn���]OozWcAe��:݅�+��H4���n�����]X�`C0�Y��z��bV$ww7c�Պ���K��{Bi�.n���Lћ̺r��mғo��S���8�c�
�Y������/p�����J���ucʗO-1���b��V�w�]��n���QfҢj��w��N�pK�����{W�@fy�A�!���P�}5��:���p��])Z���REJ���Ql���g/:��9�$�5�cާ7��wf>�U�u��YI��K�4��+N������O���s2������C-VlH,�$h4kAq�P+J9���:��w��n��Y�fJ	h�+j�-�N��1�Wh��\n���W�\P2�!�v�U�W�Mr�⤁�������e
��(*�2��m����KLU�n��,�<��*���ؗ�D�y��Z݌� "ϸŽH�3/���+��FFI��F��Q�t�f��ZU�V�mhG^;틛�X�kE������Wm��/2\�G��uǪM�.rz�P��B@(�M���i�qg�d��C�0�Y��,s���x6��4Z�8�nf&�}g�������K�ݥw�jA�8#.�wcF%W�f7������H>�y.�jt��ϰ�>&�f������»-�C�]N�8��ԶRK�v��wMI�p�+3�,ٱDqV�o��+���{�Dh���5e�J�ܡ�Y���_��������l�HK\3���Q�l�-�GXS-i�#guVh� u�MGɃg&�չ��N���u�x��`&�I�tإ�߹S6N�H-���3E��Ͱ��'��(�U��KA��h͇�_N���8!4��[�]RLQY�ze�`ؗ3.0���{��Xn4WA��'����Oq�LtA�JKH��"^�H�_@���2t*6j}:��ߘ؂�f�_g6F��N�Q�J�pgti�l�2S!J���7�`YxMF�1v-�f:����c�r1)Oy�'xqηz���#���u��Ⱥ�F)R��չ��_Q��۬��z�g*H@Z����N�͊�}F��Bf�!h��ĭ
Y:mc�6�v-2�W������-S��B��%E�%$F�[X����Y�SZ3����9�x$����`���v�؇*�KUE�a T��pM�/���Oi�T��g<�B�k�(��0�'4ϲ�Ǵ��EY�!LJ��O.���ܫ���ԗ�PnW'o�e�;���aHs���|�Xs�+{ ��n�Ny']f��Dwj���m�Fsy}1ᏯWו7uX�Y%��Ey}z�QF�N�r����<�X�r� ����gm�l+X��n��������FRZ�Sg�;6���j3D��fap�Nf�kk`(k�h\���,!s-Ksm�'��b`X�U����1P]]\y�$>敁��s�ۅ]�8�T�/�)����gvJ���&�x.ϐGyu�;~�:�x�R����Œ���iRr�h	f]�n�n!H%5�_e�Xd��*��v��т�����4�Y��Z��-Ö�1)���poI/F��c<�k���qN�)J���.�����S�r��h ������{ۏ��f��$-�3�Ӷ��oe�|��WY|:��XH�ژӴ�!t�t{ǻ坡�*�ᅜ�`���	eqK�8���z�AV� ���6�����!t��wד�u����<�+��]Z��Z!�j��P�e���Y�E�c�ڱ�1�Tv%YS��p��w{���65v1��Զ��{A��HT�����l琹��b��l���I��̂����:����CG�ݜf����2���yTp�s4+{�E^�ӹ�:�z��]c�dõ�(x9�i��̇�����_�Z
mc쮠�@_]��vG�ɝb�
L5:�VΔ,����b���3V�W8���[#R�q�Z���m��J�C�m�Ţ���-���3;���>\^���K�qux-�t�:)�X~Mms�{N�a�kOQQ�-q�t�'_vhC�@K�A6�7�-5���-�v�4��O�j���V�Z�-�X9)��.�\�]���sT�ю����b����=�y��SN���Y�r Vv�]ҧD�8��vΡ`Ц�����R;��}y�v*�!��ā&pQT*�R�
V��{0P�Y��]��Ɉ��.���6-Y�ubCHmv!��2�Mk87ugn�B���=��b�5�@Ú지.vfg��'zk��� 
ř}V���:�����:���do��%�a�����sHNf�`u���u�9k�ݖ��-ˡ�����}�Mu���`�����U1n��,�F�\6�֜�J�/%ʛJ�v�w&ł�Z�J>"L+Wu��G,Dq�a��O��wV�r�	[`؈�F�o�"��1�T�kc뾱OM�K�����|��#�bj���+�%�%��u�p=��M
��wJW*�\wm��J`�%�mkم�{hҢ��Ro,��4�=`� ��:s�z�0�k���%����A$ƷC�]N�k�����yU���ԫ��&�B����So")�������H��������<֎oM�5����r�7s9Z�8Vr[�B,wocR���W��
N�7OV�p�dV�i���ܭXU��	#Q�t�Q�Ӭ����f!Z8^8�Ѕ^�|K��]��5ӭ�b]��gF3%���{+��N�EVM7V�-��%,k�"�#.����n3������{uvGcY�2�W����[NMal��ŕք4,C�G�F�f�RѦ�c$ɴ��n2\˱jV��.w
Ջ{&�@��N/	�<z��;�GGIn��%�ْ�[�jL�w\q�Н�=�#;��Ҭmf���k�t��b�q������lJn�n���"�������.�+��v����Ğtj�a��μ�B�m7��D���ɗ�m���*�8ƅ�lC����/+<%P��!o|�=��Y����6~Aga��s3M�-uEC��O.�=|�j>�����ֵ��n��~��}{���}�뿝�XDD�2����>�8C��깘j]����V��V�΀$�KU��5\ ��F��̮��HՍm3�EiQ�PB@*	c`J���Y�jՑV�.VQ깈q���'wV)��+�E�擽�w�u�qv�SK\�e!�DSշ�� ��{�;�Y�<�2�%A��Pd�
�2lqu�%�w�hwf!�E�÷S���I%Z]�-�V����3[X��A*�n�/�o
��;���k�ɚJ�ն��z�ʙWU!Zu�v�X�oP�l����.ȳ^�r���B ��;KFӕ��X�m��N�u��`�c��ؕvt�kYmY{ΰ�޼�}ZUh�h`���������%����t/&���B�ɋ��P}DKF����ޮe(sJ���4c�)�hӣOu%ύցw���U�x�^��)��j��+6����fPY��&k�v��#��m7����v#NufN����pn���]{{9ѷ��u�%f`���uD��<��Pw\�cïׯ���W[���� -��#OO;��|�"�U)�&����Wï2�	��y��'���Zʸ�W%>�2����-�}��@�֞��k�H��������R�u(�'e�ࣆ�ډH�7�ər �#ϔw+���%��Ç�}b�J��Թ���o^7��o��"$S�6U�^�vk3y��&l��  UP }��\�9Řh��؂����6⢊+���d]71E��nLXK+	��[��h��	�\�j6���s�D����E�4V��b�QX�Mb�IE��H㘀�\U�X�
5�\�Z4V,��m�b4��b�srY1��llb�k$PTj-`��n

*61bň�lb��C�\W%���Rj6LX�j��E��t��F�U�ۍ��1ch�-��H�[q����G���V�,P���T�ά��(��Ω
�����C�<m��
��6F�{ST�0�T�z��j�7;��m�ݵG���e�sX��������F�q�1��i�n�R��+wZM<���{�+:),=�'���S�\2�*,����9*ψ�A��a袴�7��W�a��/��vkiɹgSW|�cu�'��q�����P�����GE�Oʢ%����锷x���Nl�͗���t�.O*���t���'��k�)dN�	�X�m��c(�03�G��A�A�e���3x��>�@$X]����N���Y�Q��Lh�*�{�.�����e�HxS���W5��+e�*0�'�_4���F3{~����]çc�5-(9s�z�cǯ��s%�����it��i�"�ܩ75�<�!k���ȥ���+�r1Q8,s�����K.�Q�O�JF��}Ra�
�,(� epv�o>�DۘG�����"k�BFΕxe�[��y�5>gA']%�W�W]4��������{5]��Z&����x2�V�mIe�ϴ���j�S6��3��u܈!�!�A�~�w��67T"AfЍA:;�4m':�4{溼�)	˕����b/d��>p���_h�}�ﾭPl��$2�_�[z�Gm��r��9�f
��srY�:�c�5}u�pΈ��4��=��z���m#1LX�Q����6�1�5}�Ħ(�p�BU�Ê���yO�����:ԝ=q���N��z.K;�+�kv<����(Y�;Ԇu$ 4�)� �|�D��T�������븛����P�̷��J�o�9eЇ ������`k���ڀ�I�A��f�ƌ'����&�Q�~p�vu�
]�~(!�E�NQ#
�=��2��9����V�"ea2}�g�y�u�3@�'�c �N�p����-9�_/��?+潧�a�/��E]ݱ6齺�մ��;�!��4y7@s��=_0{�Z��^�`�.[g�w�u 8����M#=b��V�꺇��I����n\��Fo��i��HɄ�ǧ�ܐ�ލQ�_��W�XW�V�q��,fϻ��Fjt�a�ۄ�+M�=۬)a���o��,	o��ĳA9���ٯJj�K�p�n�mW}�󖌈�)D�i�J����$;����N(���l�2����ʰ�`#�=�L �}lgʪ��.��V�.C� �#����u��Y��r����i�v�cvt	�:i�]��/ b�����8�h�h�S���]6$�YʏD�w7a�tѬ�m2� �\��]��LX�� ��C.�1��F���@���ė}oy��f6GG����P�ʻ'+��9ݫ2uuum+�rr�u��e��Eh�g"��ArVi;
������t���B�Ɯ^<wߌ{<-v��p���w�pw�v΋������ѥ�U0<�qIFd�Ӱ�9ŉ�F,c���X,�6��VE5hB��7(Af�H=Pe������9����voWP�鞭'S��4!\it�����s�M\>ϊ�G돆���b��M�k�U7˫v�9���U��%�}u;��R��ы�{%�,p8v�,iĬ��B�-k������������R`:���e4����)ϗt��~ӘpJ*��{J��}'H���곗d�w���h15�7T\�  ��>�`�P(l�{Wו�s�~�\}��t{��e�\��/��pT�G��StFtS�iLI(TuI]7�3�*J��J�|N����^ފ�uVb��&G>��As!����+��x�>�n�z���8	܌��X�x��;+�C�D���a�L�FwT�jxT��I�g��p�*�D�^f���v��g-2Y���29�(�p]����f�삇\!VT�@��ڬ*[u���q�t삀�J���I�3������#�)ɕ�� 2}���|�=���Wָ<�x�ge�V8��_u�o�m�#CVjl��Z��i�c2Ds-���Q��2�.�to�SG�pي�}Q��vhB����/�J�E�,3M� 4�(�Ip�c��[�nd�n���U�D`���zƇ�.s�B�clՔ/�Ո�N�3CO{��p��vu*�!�A*_����
y�	��c��߰�V*��Iz�a�
���!��zy1����t1oj��~����Q#-O���f���S;��)R��q7�y��������D6�n}=5ȁ�E9���*�n�4\,��.&P�~]Kg���m���K��~ז�;��]����u��ϥ;l����p���s�x�@�u%��:�4R����>w�-U��2!Ĺ��2h>�U r��X���)��;�d�� ��z��T�d�s����K�jnϡ�+���U��i{L|��Q�� �Kw�#\L!�e��w*���lҫy�H�rK���8�m�0.��'A�������3旆�C�_M��WH����Y�S:ٹھB2Ę����=��o�'ޘT'�W �t�����Ų���[i���	%�Wu7��[���u����	l�ͣIp5��Ah�N3��v���=�2���:^��˙J�ZIe>߀K�d1�M(��;�)⹛\����#+F=S�`|��QY}+I�*_	��GS�HA-�P��.�C��+��ra�}�;iy,�����ڋn����Z+!��DTB�8��fUR�=-wlv
{�N�rf�F�Ӂ)T��NiZS1b�{΍���ŉK�<gQ���Ը��#V�� �����x����i�$�mYf �N�n��e�V����۬�df�b�iQl���8�Rd-16P{�D ��~��uļX�ch�����m�}`?��W�7J�� ��htǡ�Zͪ[]u���;����=�^��yݕ�9�,��z����SCC�02!��J��Ǝ͇u�[�Ǵ)_��j�}2eT4;9*�O��\�F��c F�2/!���,'�r�F�sb�|�-�}�^z�^�4�騀G�:,��+���bqZ�>�b�N��ŉF���cxk.l�M]Y~��kv�m��������9y(��t��\G'Z�>�e-��M�R��*ʦ�}��&��13w݂���*�!]�C��/�m��D�i�uQ��s��U��t�5�#;��	���Ś�$����s�r��>*U�ǯt>��k�+�u�E5����
�]��o�_"�	�Z��]�i���~�l��h�=��V����U�]����d�L޷\�rv�/X�z6�<ASά�Tܧj�O����z���/,{=�!=yE}'k�ഷ�l�/�
vx �w�{ɯIF��C�۹�u<#�cF�[V5�C�-$�h�V��5�,WP�.�����Wd����|�T=��eX��jӸLח/��sD��y�5*��I֖^�]t�+���(��\�Yt�g����	�5�ޖ�e�i�MT1�)�e�i�JH"~'@ݍ�܄T�]�JƼhO��L]L�f����Q
Pc�=v�{�1�k���ah��>s��r3,�j6(
�f�� i��[ ��tH�K�������'�:]���S����8�J������ h��PL`j-߻n B�I�C>s����]wYL�]�����^nE%���+��Ӆ8:�@v�THy�3�W܁?11�*S݀#u�gz+�F�=�f�d�N�)���b�`�*�u?������*K�z;��M9D� ���]�'�,�{�߷�m�9�E5 j�8���	j�9��7,E@��A���?u�~�;6	���܂�8�㷀n8����_�p/i�V��̝�z�}o1�6'i�B�G�=�Ӛ!d��e�e*n�)b��@��>T �;�؋�ѳ�6	��j0�;�iN�������\Q���N�u�7�<�b�2��X�����h������1��F��x�k�>�^�z�3[��M�@u��5߯�"7$ޭ̘����&4:��Â��8�hB�2hXB㺟ddjt�a��NⴸԪL�輓.ۉ�:\`�N���e���Y��HW�������`۷����넭+��+y���M��,we����6�k�D�m�}U�.1w�	���_g�*����Wc�=��]�jQ)�o�"���M�@=\�Fn��c�[�OEl�q�l\�K|Q�C(�Y����W".�/{�Э��95������FB��	�����pw�x΋���uD���%����C#J��-�qT�s�6�)S+$&��07�ˢ�L򈦯�(g��,�t�x����G	��ǰ��mA�1�"4��"�_9�SB���=P�`#����Ub?U�jMqrC���z� R�@�û5c�u�̄*fxsȴ�D��7�q-�{%�%sŴ�zv���q�<�X �p����v�6>�S��) 2�詟�V�zS���h��A]����)bGíY7(	���gj9�a޼���&h�㺩Q�7w*f�3�ܱ�jE�b���s��%�:�ynŵ,�� ���D�k6�1N�ۓ,,�̤]=�.��1�y^Aݒ��ݰx��@�^�̅j�����Z�.>��l\D�ᩫ�S��r��D����t���̄%���� L��@�L�d	�qou�"�6��#�7�?pX��c����ݑ���1$�]RWM� }�����[S*��$Wl^>7�VY��=Ƣ0�0�9u�p��Ź�D�x�9���n�u��<���{��3:N�1��ZcF٫���ht�Z*LTrN�9\�c�1Q�� �:*�/��u�1G�_=SG�ٟ=��ȭ���\�xj��=��b���\"�s5�r�n���G"gf39���Y��T
�!�9](2>U�Ć_]y,�7�8\w:���lC\R�x�%�u�̸sLj��P���F�<���=�Q�u���zdF�c��Wi��*�m�s��BV�q&Gi��t1oj�������2��1C�d��WYU��%;����;d~0�hs6��h�}^5F=�[.��@�,�7�u_m�*�l1xcE��� �/�Vo}&R���D=���O���w[!���X��}].��:l��W�\���
?m�YN��ú�����+Z㲈Ʋ��]��K���O�p�&�T���٤k��1N�.Ro�y�xѱO���ⱚ�W&���O��Z�F��=����a���i����#�nH�`�ګ�Tս֭]S&-s
�L[|@�KK�#;f�ﻻ�����D���(�w�=�3�P�y�#!ܦVC�����8C10��l��VN�����q� GlA��3ԅ�L�7�U�� �7Vk��0� �}�'man,_h�U_n
��,�n��$� ����#PFwL�њT� �Y����NL��q�d���ZB1��Kޔ5:����f�V��k�<�t|��8���M�9��3��X�ؗ`�<df�����^��U?e�=�-�;�Ed3:��AUL�����%�o'J� �8�u��3�6tD-;|�C�t� ^���NcDT[u.ݳ@�G�W�k���ٍ�b�3;�VS�L�f��Na��=��I;A������M&�蹳1|S�ç\۳�J]�:~�3+R#�( (֜E�J�Pu��Bs?rn��w��N�V�6��u�:���VLW���C�St�ϫJ'�a��׌�f�-Z�u����|�ؗ\7��ԣh�ܗ9�������ۂ��	��*��ƾ;6Lh?�G1��x�X��o0n3i�V�i�X�^'�;%��<���E���h��@����&nAp���˔��U��N�$�{�+Nr���0ӽ���CS��
}��f��q� �Y����N�6M}@0�YyQ%���e��p<9�j#�4���=��9sǇ*JRfc:��b���S�Ӊ���â�c F�'T2�Qɛ4ܡ�3�L>�a�j�;�s���xNykո�bp��?�+�Q]����w׼��	�X�m��c:/b�뜇�jkWCp�'�`�7��|�Y7>��\��p������u��2�v��1@�ϬYy[�(���p�����l���{O�ُ����s�<����=���2	<T��y�θ��}XX���/�)iQD��_@��pV�ഺ��l�/�
�����BC2�Ew3��ԜKf�fM?�?
���`˭�O�_��Βt�=ŕ���|!@�e�΢��_N���P�VgN��] <?!�ӸLźTƩ��˕k4��N�%�*�\Vc*l�O��uכ�نԔ�'�p8K3�����2��i���W\)�e��Q����X�`�5��5�����p.��j�M*����Q
Pc��]�Z'��~�N����L���,�3|�i.���4{�B�u�Z�k�G�S�xT�,g��g�c���>�����B7�8&���d�+��Mf�
"���ַ��@.�=�u�Z��]vë(w6^X�7nZ�V-�����a���Y�� ӣB+6�d��{v��\���H㕴��TzH�jc�]9L6�[,���`-��-A]�p5���wv�����))�[n�����>�7P�ھ[V���{���W��]bM�y���l���*%vj���"��ɕuϻ*�g.��Y�0'MŖ�!����e�}���۰�[3`�X�<��i��˫����]x٭�<���X���ј��u6EX�J*teG���I��-���4P�Z�j���Ҿ�Z�|�����n����Ӏ�Up1�XH+�{��`	\}���75J�˄&�	�k�(��7�V��'�8�@��t�b���V^�K/^$j^��	r*����!MG�=����	��^��F�w;����X4�/8B@)9�:�cS7{����f��=�xgֲ��Y!�/�u]��g�6v*��=�U�p�P��Se��|�@]*�׎+ǑpܛB��7�].�J`�Ӗ��5�jn�^KٜY�@|j���S )�#v� !oW��ꃸWnySڊ�9%)9w�E�[}9]��$=˸��ed�/��|zJ�Q��S�+/�ڢ�L�`�if���I���'��7)�s�K�9��e�AS��L�.CdW�ئ*�Y>���U���ĸ�u����"S^a
�a89��w�Kl�5o�m�ъ ��i�鐦Qݘ�kJ���z0��wY���&�t]�w:�� ��Zn�S��&�Y����;`�tP;�u����V��̺�nE�qlXjX�F��yMP�E	�����ݪ޵.W�iʙHl����C��b�j!��v��T[FmnnS����0��:
�f-w٤[���@�ިg�$]���m�GKX�>��Gnj�9�zʊ�h�yS��1o5mӺ
�3�.�����Np֥���j+��V�+8���q�[2Z�;����g����X`�+�o\�ԫ5���5`��\7e<�`9c>�l}1_RVV�Ǥ]���u�P�NE]�r�*��ǽBM�e>f��[ѷ�˙�וju�����,s{̩������r���R�`o#�+�k�r��]�i�c"'qJ� �N���\�"ژkOJ��
 *���[8A���Bf��G]�h�}[��-��[��
�Θ�,i�bȳn��xX�V�1Z��qqږW1��!�޾]�������w:����R�O_b��n�LN�t���t�"�I�.���nu,n�q.�r��Rq��@��{Xܔw&��������i�������s���9���[������um��D�t[f��w+��Պ�5ٷ�������_�k������l�ns_���^.��G5٩*+H��\]�<
�0nk�0��n����fm!U@U%F�"-%�4lFJ ��I(��E*"�[�q�m"�(ьc
JJ⸓FѢ�s����E��!E��X����b���q��\j��n8�Z�j��űlIUQ��+�U�F-�Z����Th�5\[�ƺ[t��k9�\j�*��qnM���Ӝ�\d���ι]5u4Rm��"�Q�n9-��ۍ�\\j5���-Ɗ�\Uj�b��j��F��h�q�n5��\Z�"����n(_�Uw_}`W�.��4�Iu���nz(�}�%����)�a�e%S�8�B�[��S�u����{��1s.�U�o�n�7�]w��F���=�����o�F������k���Z���Z���]-�\�67�꿷9v����������6�W��-н���[�r�Z}����������U�qy�����|DDԢ�9� z�\�E�n���_���鷵з��u�+�m�]y���-x�͹�o��~^������s�m���^o��qž��t�W9�_Λ�_z�5������y�龯�t���{��DG��-�]d�������+a��I_��_�������Zy��~��v>.�t��ߺ��o���7�s����ߛs�p�ʸ��qq����zz��\n���o��<v�����~r鸿��j5�}Y��D���R��ytw���T�Ӿ�j��+Ҽ]?o���}W�t�o�{�KŠן>��[�q�ϟz��-�].�6������k�q|~{�����q���Xy�\[���;W�s�;m�v�����UW�F�՜��o�л#�oJ�3��{�����7��m��u�6��O�}[�|x��s�om�o�{t׿�u�/����>���צ�t�z���{_Wj鼿~�n�scq�/[��ү,^�?}""�#u�Jkk�(�=����������~���Zr�׫���n*���\�6�齶��o˧�ߗB�������=���~ws�-q������6��������{y�m�K�y��U�  ���aub��7W�g��{��2��������_���KŽ������v�]5��W���v��^s�=��]->��y˵���n��s��q���\�����_W�ny��מ5��/_:���>�>�����~�|��ٞmL����x��N�~�������r��޵�ƣ}�����J�n{��9]��n����[��֍�^ۧ濗kA��|�+����y�+����t�|[��"�>�>�"�Vk�eMf�:yJ�;1��2�>� � ���!��0>1�q_��}m���o���ͼU�r^���׶�6�^���{^so����˥��N���{��5v�V���r��FC��>�p�DbQ�H�F��S��ϝ��}�z��؊��+�֮z���{~���v�Ww|����|�ͺUǺ��^-��>r�u������ܿ����W����o=����6��|m�9W�Ӧ�B��t��q�\����y����u��.�'��.d���:E]�[u֭V*�O�%?�1�VO��?R��S$�\���3��������\�m�RZ���fp����#�HB7Z�5>_`��,%9,D�ʶ�ӳ6+L�6�5in�СH�>�Kvq�2nȵ���]rN;�!��B���J_���NI}㯸���/�ܵ���9w�6�|]��9|m�9�˯}m�W���=��Zs�������/�t�-���}�֮����K�������W�z�}�q�����]�����L��#�=�ś�~@�Y�׿��k��ݮ6�kſnst���.6��ku�5|[��o�|��o�{��������q}[�ޛ��Z+�ok��ޯ��b#�;�\���Y ttg��,�X�F��KD������W�nr�+���u�گ�Ƹ�z�]_�t�������ݾ�q�5�;Wj��>s�o{�߽����v�뿽w���{m��|�֋�����(�t�%1O�LtՖ@�c�-�~��W>�����y��U�/KF��|��^5�}]-뜢�+���t�������_V�W���7߼ۦ��s��ѽ�������zZy�ϖ{�sN�ɜ�d�Y9��t}��ޗ��o����￺�U���o������W����׋�yk��~���m���W���ns�q�q��5��W]r����Ӝ���7����żrv��?|���]9�U�D} }�0}#��T|�`�W޿un�Z���}��[��W?/������oM��/���_�zU��/U���Z��/>��vۧ_yk�7�^6�t��B��'�|G��V�_M�_e��瞍ʊ����c�D��G���?��\U��=��s��o���+�}w].���^|���5�t����]��\[�o��W~�o��t����Z�W��\^}���z~mү?w�v�nڸ�������Ͽ�]���/ۂ��@�&��@�@��ۊ��˩���vۃo˟9���{��-��:[�>w^w�\o�z���wƼn�KGϼ���x�M�t��_��j��k��>��Zz����뷟�z������^������>�n=�Ү./�߽k�x�|��5��v�Z7�y�n��oJ�i������������ޝ7���h����n����ޖ�~W>��o����޿w�'�(E��8v�o��#�(�T�Z��=~���9͸�}�:Z5zq������W�Nr��~�^ޛ��]/�z��K��}_�\��ok�����{kںkל�_y\X����r�W���ۗ���}""�>�[�:��u��8vN��*n�6�.yCg:�I��>�bCA(i���)֗��pL4]��t�uťR0ksA�5�
��3��H`�Zg�n�jB �F3%5R�
u���@Q�<�9���{J�{fԂ��	۠���}��Me���>�m��8�[�/�>�^.6��U��}F��;z���Wm�n���T��ƻk�^~�[��Ҿ5��u떸ߕ�^��/�/���{n��^�M�т ��A��}��3f�}t�ֺ��]/߿z����_W�������ۥ^�߿��W�������v�^+����������qo��z]ͻn7����گ˝som��]j�o��Ҽ���]�1��u�9�]a{L]OE�[�Z�c�׍�t���t���]5�.����t6"������zZ~����w��>�Ү.]so��z�ͺ_+����h/�����y����?r眽6�o�����^�k���7�����޼�����z�~~�~�Ү�5��/K�����v���׾Z�ל�6�����_�q���9�����\Z
�����[��WKNr��޶��ߗ�_[�󾷥ţ{_����oK�o���̰i$Af�m[;q�v����|aG��o��6z�qc�����U�q�5��]w��ۥ_�����~s�F���\m���[�羫����z�h�m�Ͽ����ܺk�\��][���˥t|�
�(R��Q7g=�{Q��������x�k���}���7�񯋦�޹����-��u�Z}�+�뮮�x���z���]�ύ�k��7�ڸ����z�[�q_V��{��~�g��������H`+��cB�dK�w6��7���U�˟�������E�7������Z�}|��Z��]7��o/��7ƺ]5�|q��lD_��t���y˦��үW��v�x|Gɟ����ɱ��bl��ZKǛߪ�qh/���}���[�[����w�_�t7�^�ux����������o}\|ou�Ϋ�z�~��Ϋ���.��W���ۜ��Wk�\o���W�st� �� >��S����%w��C����+��םwޯn���k��z���/KF�z�����J�}��ߖ��_�����ݮ������z����*�q�������\�[t��~�Wm�۝s��_n>s�:��T�G�BZ��-Ώ,ѳQ�|�W����\zf/�hy��`Ұ�s*ۨ9;�f��<�k�������Zmfv�t��Z�.�raʞLx�o��=;��hru��ڕ$���;�a����6���ƮX���Q�9|ñ|i�>��4�=��I��uA�i�S���}Y:�tf�S��3u�z�����oqV�X_;eF�ͦ;?����#�m���9�Ç��@���S١(������?*�I�amYg l�+ �@�67է��n�^��w)�֟����kN"�g��v�y�l#����ipy�|��Ot�>y��>���9@j������)�to����먩\��xZ�\*ǌ����N�gdܙ�]^�\����6X_448��d��Ơ��w�un��v�W[J�ֹ����?�s�G�
W���s�����P��dڄ�\C�93wX8#�V�۪�S�;��h�n�~Q�˩zN�������a�N'Q����:$Js%;��V�D�k�X3u�Ť��1����8�R�	�(��/�Uh�㓭g>}4�Wˬ:�ڞ�a<���z� j�U�V+�n�^8e��Q|����O 	t��]�2���z���*���ߤ�K^�v�l��~bU�������0� )m��أ�ե���*Wr v����yLB��]o�|��q������H�Ek��5� �"�W�~��b��k��CY�Ȇ�9��Ǻ���H�B��1��Ҕ��
�	x�{�<�B.�nWG�SZwès��]M�yjl�0��9���+���o�gt�GR��n�n��'������]f�e� ���^���M��[(3q�zYD+|�C]_�}�W���d���Q�h��V�χ*���ӨL�t��S��V�!����X 
����xז��-S��dh��:7	Fj1;zr#��^�!���b�L�/>�8
8�rջ۹��[oyGU�C&��,�ē��Z���J`��봎�'O\��t�wr�-ho�]��#�<\( o:+@@� [�N��xR�o�'oC�^�o.�[�qٕ�öy7:񳂬�	���p*��ـ��$�J�05tv� ��(��I���g/�t_N �i��h�i7Z�w�D����0���v��9��W†4��#M����s�P��UM|ۮ�3Z"�`�wl�U��.��?bv���Xh?=���;���{�3+�Q��}Q˨��R�4m7@s��?HM; 3نj��UT�yGa����t�vG�(?�����:�XV�z��gܝܘ���Pܸn9��Pބ�����%vqW�,�����`��a��T��^�а��u>���:u�{���n�Pn����me@LUQff��!me�$h��i'�3u�I�^M�`�Sqgӟ�B&�DM��E������s�[�Z�Ӣ݉Mf����B���ǻ˘J�y�@���{�S[]Xj#�w��1��V��2�	���T����}�;}ڧ���D\N��5�͝BxX
ZϦ�HWܯA�ցʌ��ۨB�C� ��bXww����.U�-���t��CSB'M�=����	L`7b��<��Ê��O=Z�3v^��Q|9�5G� ��hduUB�L1�b���tg��^8�S�� ���hǵ!�ߜ�W�r躼�KϷx{�I��=��%&;�s#!U|�YL��p�F>עZ��A^*�},ar�����H���"��KEϩ���x��C^���uZ�]NS+"���!|ui��q��z�v��m�.i�K��
���Q Ȅ*g���K�9���C�>�z!��:f"��u-�0��zL�g7��7
�P:�/�L!�L�t���ҥ�8&��hm��2��6a�%��,p8i;w#��F�}��l	=�G˸Ϛ_X^���^�U{��^�}ض)ĭ�B��>;���3 ^ÚMD7T\�" L���ʘ�-���
Ź�X��Ô�������H�:!�����&썺ubB��P�%t��YD;�]�e�E�BI�Lݻ�̀F7��&Hq8pM��ݵ��"�"�y��(/u�zP��f��N��g�AO�<�Z���-�A�sך%���*�A��%k�;��Yi.=�.���j>(_J���.�k*M��3�A��*ND٭��|�� >���~\/��L���'t���+�&�.��As�s6�P� ��٠x���$���7�S��Q!��lmX��$PC��aL�guHAq�1��;,�s��@�����&U�N��˪��вDwe:6�~�F.V�`��/B�;]���%w#Q�]6�ݭڛ��[w������+�=V�:�\(�vς�?5�ve2�=��0O��yk.��.�Z��V�'V"�:�1!�JfD.qu"*5�'X0{L9��;~�c���wWnQ�ǋ�1�f������~�|�w�a=�b��X�O*$g��%�P<���
[�qv�o�=m��vޘϑ:tDg�OnOMr `�q���qM�^�"��-��r�p���p�}��ٳޤ�]q�m(͉���0�
�����s03�N�+jlFm�̠�$��e�4��]����i��������������!�@�p|�y�#{3�}�V֯W��l7�p��Bi��{�=7�C@h���+_	M/i�����ý{�lד2���#���B4]	˅m8��;�h�����B-	�:� ���>%d�����P�B�^f��ڀZ']<��X�-�W����*���"�;ʰ��5SJ�溁�g�wr\�9>�֧j���^d:��E�x�yh������
o��t{�:�ʍ�F�������zT��] �(�<I�3��5��Wq����1V����h]��Y���:l�ƽ��{ԇdC�����{�9�k�����N�����t��X����PH����֖�M�����0���ڶ쌸wV�ϙ�D�{)�/��S����H�_:�a#�. B�7δ7.�0��<�`qm���xGB�j8��\
�妃�TY�P@���<�hJ0���Q�?*�'h!��e��1$����*_:��{'����9��ejDwJ
?V�E��a��p��8w�A�%�\�}#Wh����\��k�J�X�W���>�י�҉��v:t�^3)��Ύ�BQ�*�SMV���塑	*�7`��nX^46ˋ0'�*���a���j�gf���n���H��:	��J�ܯ'<L
�{n����#�������p��p�^:ڕ�z�ת�}��&�X9����n��0�����q�S�'D�s�� 8�F�=	\n=q�l\�{F�T�-�ʺ���5;���,-�D��V�6���!��A,T�����XE ���j���"l�;W�X�s�3������ZfS8I��
t15j���)lm���1��7b���� �{���g��LP�)L_�p�8�N3�D��r�%����U��N����%[�P�����f�neƝ����,�2��`�	B���q;1��"�w���zLJ_)��e�A.���U������ 5<�Y~�w���3C>7�������^�vj�y�R�1&�fk{�@�e '���75�)�E����U��1��t�G�����)��{;��yӎŧ�%# =9�,.��
���;��\:T��B����3Q���g��A���fw���U$�C�J3_F'oO2x\i�MT1�f�cl�A�����l���p�� ��'@�x	)����eR���㞻H�5'O	 ̠��ܭ��^i�hV����!_�r�6��ʾ3�P� ?�-��t
_m��bs�3̯m��͉�Ũ�ꎚ��N�����J~����" 5*�&05��eM��3ڲ3�ν�T�\A�{ֆC��f2�M&�@�V�*�2$!Zh��$aG����y7<�Q�V��&�^*L��"�OmX��3���\����w }�Zn�5b�`�X���yl^�χ�+̇t��{�*��Y��U��j� �\�{�����u�v,�Jڎ���Ķ{�3��:m9-S���6ܫ��A�~���ﾏ���윭N�[��f���	�D��P��C�I��^C5��,!�Jwl3n�7�D.3N��}E�bf��WU����VV ���5��������a��%��<�:�+���{j�k싮5}�������b��%-[g���;Z�5�yp��N�L_�g�&�� ��.���f.�jx��y�q�`��t4�Q��:`Z��X��Y��+�Xx[�LA�n�����Uv5�F�Z9�ڔ��X?�ʗ���kX3͝AT�X~��M�	
�0��C��A����2�l7����y*84e���9M�7�=���Q�Jc��*{�!Y"��p��:R˾�C��O��]hgʪ��c�'��.9�p�s�c~G	��2�䶪�<�<�qgvZ�Y���ze3U�/�.Q(�;ι����CBf36�B����p߅^��p#$�:��KdI��l\�g�2�b━�a�;F*��ˢ��y�W��=a��8�1I�ꭝ<�Fa��p��S�A�W���B�:K^�M�r��4!_�]1���:C}�lMſ��F+Sw�h���M&PF�^��}�Q�N��#���^�2�h���b&Tz�u�o)g����̰V7mAE.S�� 
���ѠTrˡ��q�w]/��6zf#��Jf�I���%ֹ^ޮU.�	����ե�yo��]P�FF�H��a0	:@٠q��)C�����N��t���yǻT�m�V�g&��wԖ�6��uGbU�Ts�N���!������ :�pݑ��Ì����2�J�ѕ-}�=@Ss��wY�+29�4+Ǳ�V��C.��
��`c��� o�ۮS.�4ls�6��̬��o��Jjr�T�uh5em�}�QoS2n��o�uH4��{�q�B�[P�7��w�x��{W�� �헇u�і&�ϱVP��s�n-I�Э.��i��bYJWo�K���3Xd�C�OE����0YΡ"X�:�@O+�I׊�Y�͎�K(�-�hUÕ���!�'��;�%�S^��(��͙����wР㮣�ۆVj<X�l��6`<�L��`䌫YC`F��gQ�ʋn�w
�Á�0�T/�\��t�L\�����v��Xm�z���b����K1�ZQ�Q��]��Z�N�`�;h��:N���7%.Sl����9�rƦ7���o�4k�mǔ������m;�.���
��X|+˶�v���� ǀ� y�V�ZT���܆���"���פs��Wח%�c���� ����gm�#���܌Ӭ�U�
��in�X��6�ͺ"t�8z�.���G�,�	L̗��{�R����	��ۉZ+e{�)aޏ�p���[u��K[�2�M��Ю��p��Ik���8�`qa\r�{�%�}btԴ_+��h�ws����Uʵ�n��,z�d�We�uw`!�h�E4MKu�����F�eN4(���g%5Qz���:Я4ms�CGHL1lz;����WD��=�3:��ܕ{��d��l]������b������ӴT�q�cC;;��ڭ��������Mt79)��:�}����#:�s�v���TP��B�U��2�3���NNX\�g
v���[���}]1p�e�;{Cv�W��\�� }�����40�wQ�5؊|�Fe�����z�w8i�u#.%�g��X;(K���7՟�e�j� N�����I�:�R{�@x��6���v|���1C���z]�ܽ���A)��v�:��Ju}[Y�d��a���Tg h��@���9�4c�>"O�:k~�t�TV�/x037&�
�T�fyC��<��ٳrQ�@p�C�#���V5%����n�N��w�t�t�}�W{(�W,�ɾ�#��gjt��u�c��/N��c�I���5s�z�*-�tGC�ݱ[���̛�W�]�a����j�P���%N��3ۈ�o'}����ĥ�\T�H�#�"��U���'������\�ߝW�ؠ�n5F�6�U��\Z-���ƨ�\j��Q����Tckq�mŋ��8�k���8������Y5Q�E�՜��j�b��W��9�ӊѱq\Zs�Ʈ7�\mq\m��+js�ɨ㊸��F��*�����\�6��F�֍b��q������D�6�KF��j��Ʈ1�6�k���j.s���r�9��qmqq[��4WEq9�n.+���Ů1�(��m��~�������b�h��4����b��Ny|���Ehu�ob��*����G`�>΍}�ԁp�VNV�:�?�UW���V�9��
q�`I�ϝ�vDX��p�q%�h/�S0�L�yif�\�d�l[Z�|��]
�-zJ9Ŏ|����v�7��&c`IJ��.R=��m)�QP�U«&�/hˮS����kv�y�p�����S�3M� [�4��ꋔ �����XqR�y0up��ʒ���ΣՂaq�]��I.tBG ���7dm�:��LI(;3Twa�}oQ�Yi��'�\A AǄT���������]m.c�1nf�*�y�=^�J��%��L�}O�,�ǹ�H=H�mbb�*�A�f�w�U�:Q\jLW��;,��W�\����Wy��3��5���:���� =�~fW%���j.�V%.^��p�[��xX�5��3�.��U�Sʕ���9[!�� �i�`#?X�TT/}p��E]���?:^Wf}L�2RʹXѮ<ggv�����^GZ�4"Ӑ��s��'4"��]H�� �`��#1Wv�r޿��&�f�;�B����Y�̽�2 ��N��-�S������
|�FQ���rU���*���d�6��%�	L����)�'5�շRXd�&�C�W(�5�DV)�i�o�s�y�F%KS"\���ͦ��!SpC�
���[���V�ϝ�D]�ge3l�6lTh�n)�@�S/9��}��UU_qf���b��ţ�;og|NXj�on�<�Y�.��n�2z3 �b�E�>v)�8-�������?f;[�����ط�{T���*�z>u��|hZN�+��d���]Wk��(��p��53��(T���+	OɊ.C�\����4�X�j6t�U
�容6��+6!��[+>w\dȾ1I����[�~�(�|#K�gϐ�L�~3[9��W�}^fuС��y^�q0�c�����J����QC�=��|aAҨb1���-%O��f2���T·�"̏����9�C1�h����R����¡=+�y:�z�^�J}��pa ���MQ�S9im���(v�Sv��<��u=�E�G8��>���ͷ1�Y�jA�ӵ��0� �3�!i߯�hy��c �Ҵ���h���'$��ǹ�:��{%�X��8?��1 �١(����ӣ�P��8?mvJ����{��uN�4�x�	ԫ�FUE8U4��$%�@��C�TV�N�p���t�
��nS���p�/�ó�k�[�Lp��8��iW��)����"j�	 ��Vc੊��霮�rÈLN�<�s�k���K���tl%����3�C ���9N�Ř�T*ȵQZ���V-W�������q��}H��� M�庋#�xh�ٰntT?Ͼ���ﾊ�m�uvbx��?G��|��%�k�g�?���>|��:	>ӿ���hSU��n��A�g�f�k�Z�EflllG%W&�"�ܰ4�
hm�\Y�1T2U�����g�9�Y�c�tc]��Q��Evg��έR
��Z�����3\ �{͇��.k���y{p�Ck�m�Ib�`p\Y�?�����;y�,���L�1Ew�_��g�e#~\�l�-�gKyr$?�9��qňczN'��d�d�2�\!Ҫ�}����8E��o�&���Yԋ�'�OO�
�*��!�B��kҖ��h�E��V�����NK��܆���*�^ݥ�w��ĩ��?t;���F|o(���-*NW���`r���x�}]
�Z ��< ��I��r�r�u�F���~^�rQ� �pwJ����s�{����Lf���9��UL(� v��Bf:T�⬾��=���;�-�^�t#��:Q��uc�Id�=C<�g�H�P�l!(�Dbv��!�
0��+�ep�B��u	r#2��o:�:C4K�[LA�[ޯg}��҉X�yr8��R��8���Kp3��h|[�yu1Y�36�^{����P���I�E��(���4�fv��k������BU�m�9���2�_*��&���{i�uf�~�',�j��㞟�}_}���gpq�F�)�Ӽs�����JH"I�#�`��.�c�T��E,?�봉�(y4o:*�Ō��x�^$ �{��jv��4�n9TA�A� ���>�ρB'�֊��u5=����eu���xn7]��7pxتS�D70@@k~���_{"���	������Z�e8�p�V�9<�&cFP��R��ҟ��M�@}t�TѐocҬa��{��і`K�y��"w�Ӳ����p/>f�0E�0	���6����r6����Q;R^���NhFi~e*�WR���+Mo3_W.�"�JdѶ�� :�&bS{��I7U��u�`wMx�b�N�`���?].��U�Ú���H�J�/��.c�N�N�����t.���T�p� p��0��L`BJq���(e}�B��]4y:Ǹ2�:ꦝ[i)Gmt?�t&�����gPS�`=��}6�B�z
� �=eHk��hA�3s���L!��h�GG��O��dD���}I�]��
�A{_*ȹ߀9�b'elYR�w\��Ƣ{�xȟ���]B��ua������h�u�:吆j���>w^�Y���fy��{����d��-Jz�w�ޕ��Fhv��z|�\�k��b��\���v��\Fy�7�Q��f�;��r��諭���i��ǪaD��U� ����*�� A�[=�{\"��p�y[F�lYӭ�:4�H��2�;�=WѴ�AF�;0�mV��1���
 N�dgЪ�CBb�W�k�`�>W�#~���z�Ӂ�l׉���X9�T���hگ��@��P,�7�r�U]���TH飋K"ج߹�c4�)B7]$�2�T"�4��6����Ɋ�^�vf���b�x��2�n`3���|�?p�0�|�U� >(g�3W�3Û�bj�2�k\�T��+oU!!˞.9Ĵb�{%�,p8i;w#��F>�f6�J��P&H�1�����w�����fI��T��_ҕ�������x� �sA	�n���@�������5	j�!�z�a�.���Q���.�!��P^Vp��6�)Ո1��ml\���l�ܧa_8wQ��mI�$?�������:L*�.��1��8|[�E57Ȟ�c�Iս�z�߽�0�9�H=H�l����^W���=�{��=��Xי|����Tx�6zQԪXC|�P�ۻ����K}*6���ٲ�+|N�+�Gvm���}��s�e���,��T���,][�ww�
WXT�*���mPT R����LLڠ�m.�OtF0 W3݊/�>� ��=©�Vw^��
�}��D)����՚ƚ�.b1\Q)������gܗ���h�*��/Yr�!��xE����/��Kk>��wr-����� w��*5�T
�yfOE]��)y]���k�G�������"*>Z �иxM�pU���]�Lyb���s������6���ı�s��S��A�V(���dF��[5�e����t1p�����oD?mD�-�h�L.��G+o��۠�|NYfՌV�N��N��1Oj�:�
���u_hf+����,�ڸ����q���5�}֍����n����(͈�j�x	�U���u��F���[=J'�%GR�tA�p�';T��A��H�u���xG��:\���ݗ�*f��GGٽ�s����㨡!ܦVC����\k������UG�Ҿ+_����_�=x�}ʴړ���0�j��НXQ�&ˌt��w��j��,�F�$�?EQ��M����cn�u�OT�tg��:=��OݝM��r���C�p����y���
���'3� �c�S���*��TTD]�dFN��*﫻[�ܚ�w
��Vc8�3�b��\~�Ύ��|�Z�yŤY���o�&�G��X�l�論"CZ��w1��ך����vh�ouLNs��N[�Ż1��zb�R��z�V��'jz֓ߢ#ﾈ�y�ƩW&�y>�6>���Qg�g"�ۉ%���\s\�Vݑ�L�C]��3�����[3���qD�����Έ�¯�hx��f0�Ҵ���C�-e]̭����^�
���tnUl�Ń�9]D
� m@<�h])�2���Y����K��ȣ�#-���{���������9��f�Gu+F#��^��k44u���,����w�ՔB5�)�S�X�~�3�鏫�7N�K�ǎ���Q�"�;� �'y�������Pd����-��J�M�E�)�`iyM����+!�
�Q�r�"s�V����a�ާ�0�w��j«�t����s���Ίo�o+��[�9-�<�DI� U��l����b�ۜ�`�<6�(�d���Ջ�z���T�f�]����������Vyj���BՎ�_�Η+&�Z��m�Ī*x�PWSe��e����	��q��)o���L\F��8m2��0��zx:q;+���/{t�4���u���Z�3��7L��hK���Ώ��]O�;~�ۮ�����6��<ݾgz
�߹ 7ZWnT�*]c��˲�ڝˤ��/j�%���\�=q���{�:�
!�locE��n�P�Ձ�3F ��:�ΔW�m~����>�%c{�8�� y��_��<��������-�~~�w���;mݻ���U��8�׉��P�s!<_Ւm���+�(=ʓs[)�W.�h܎}_�65�$���x@�c������e����Ln��8�}����tF��p��f-Ҧ7e�Bs���F�gJ._mQ�	<N ��u28E}%�F����5��Ӝ�2������t��;ojKB��pD�=��(���& �Z�ʧ�ҭ�t��|�xX�����X�%�v�x��\����w�1FO��N��z.K:��ʠ�1 � `y=3U�����&T�s�����x���(?�V����<5��'�1����R�����Z$)�7�Y�6`�}��}�(W11���6!&��s���30���hӸ��"B �b�q�zTt�<��7jT���t{���߻4T.SOBn��3X"�uLR�W-t�lŐ�25[y�)��p����A�[
Oa�6���8��ٸ���)�F�t;�E�s�]uRF�4�SI�tN��j���s}�Y�N-����D,��ѕԩ�u�A��qA��Ϟ��n�"��r��a���}�g<������떨�K�\�1s,��e�R���攝�c�/��z��r�o���U7-g4Y�3��������Չ;��.� ��	�v�:��7(E@�c3�!��j�+9�p�\�x�����G8���tMM��{���{%Xfq�g��i��v�[0!͉Fه�9UX�YY�saMWv���p�i
88n��25: �������i�{�Xs�r	{V��V���^c�3}]���1�;+z0�~�=L��M+��7����Ɋ�
�߶����0�\FK�jal����n|�ncEDI|O\L �}ld��`����p��y\/�Ǖ�~*����[\��]nr]\I���+uqJ�Mш|k
�� ��dt��	���!�-���S͠�K���x΋�h�O�a,^�R� 43j�6�B�:P,�1o�q����S��t�7��Ğ��)��B�a�B7�A�,k�P�-z#k�������\�=�u��})[�5�u4>��o�0��C�*��nA$��:�/��2��=R�zE�M��sˊX��������v����):n��T��0v>�fk]�����ORɏr����q�^�a�?�-��H���r� mS�����ņ	�h��익����(wa�ɭ>����ǲUߛ���>Z*���5�a����b���v�Nȟ�oR�M���_=�*��ܛ|�p��.��k:��*7P��&��BM�>���>���E�r���
j���Q�Ԅ�� +}��f���uJj��Gq�=mN�9[���o�`b��M��}��iC��a�
�M���NB�r/0m�y�.qd���T�>��G>�����}�%�CZv�R��5�oS�����s����찜@y��B�s_q�f��5+�k��(4�J��s�nz�-jZd]��ž�����nj8��s�[�S�];wR���V&��T��ά�p���Þ��k�g+\dO;�-��34��շ�ε�^]���m�qf�>?I�|�^���Nu3��8�Z�tK�Uuh�沞�k��V?��YQ+g=�˭W��$�]��s��n{���q:����x���U陷޴�I�Z\J�z�����>"d����]*���=���=*�4j�z>\N>6L+��J+.�k������ǐ��J�'n�&R�F;ۯ[�%u�����,z�,��뜳!Zlk�)��7rњ���ٻ�Y8[͌��W��[�7iEI�Ӎ<�il�'䮊��M��/*P�[���ԠHG��4l�Ji��T3U]���]ޜt!�\�#�|!P���킎9��4�v�d���ΝfwZ�}���b㘘Ÿ�N=���Q�h�8�x]�	���WR}ъ���G�3!��:�㺨���:��ѥ��}��ѓ0е.��1:v�yӴ *���،9��A%�C�I-Z��y���"�ޜ�j�%דD��h<mos����Y.�v���C��Wcc��e�F�}����Պ�-vCFiZ�uj�Ҷ殸�gg�|�Mɞ@�M�/�?���!B<�'��r!Z�/G<�*L�@�s8'b�=#��,�[��BX���s���Fj^�xT��*-,���|t��$@�ցݹ��&���#���	�h������B�+���G+���ت���Nj�E�Fd��<�G�ݸqӤ �E�3p̎��ܢ-�T	Jzeڙ�8ԂZ��Meӻe�&����t�UG�;�K��yV�	�7�b�>r�rt�ʅ˱g�v@�l�h�K������L����^^�X{��p;jQҥ�)'׻ö<�pC�D^S�R���Mk�
�I��LR���5r�YK��������1}��/D��V<���/ywN�u�ފv���^w1e��t%�o��	�}KQ]ut�=�:�T�[�z�6��5������PP%nf�w&X6魂�ԅ��Ɏ���F����x��Rɼ�:�M�{n��#X[s��u�}*\ފT�|����kM���ث�N�h��5]��7�Xs,>�=ώ�푔�mI��v���=�inh`�+"�Å뼡m�+CD=����t�붅ҍ�­�ڸ�V&yʣ?1�����{���_��s-�p��LW*G��^�e��u�GUn|��ZG�̵Ȫ��f�F��Qu�r9�]'K����Uwa��G����g��ʗĕ�k)�t�aSi�����,��/�p�T�:[=�MMN�Z��ԓз�*p;�q�7���p�X.*��������v��w`xiΙYf�c����R"���=O{��"6�5ḍ��^��\M�ӧ����3ksx:Mi82�ꔐ�hf�Xz]ai���h����]�e%�F�&3��EXt�˩�{�:�[�:�,���>�W����+^Ҍ����#���v]en�v�Iw&�sf���N�]9Ƌv�~ɋ89Mu���u�t�ȶ�_("U�kxu�bò4����:�X=�I�Lubf�Fq4OE8J4r���Ƥ{(����֔
��u�{N�}K���6X/�,؂������0��b>�o��(@�-<�7$iޜӈ��mf���z�y�;��\[t��cq����Ɗ���n#�k�Q�l\mq�Nu�ū�q��9�s���q�⣊�[��m�ێ7�V4X��r��m�E�4j5�Eƨэq�qY5q��&�9�k&�\h��I��Tm\X���F�ms�����m�-�\lZ1G���9͓�c��9�Ů6���ns�����q�\[����J�Eq�ЛI��rF�Q�s��hs�-E\Z�V�
:�7�n#���1k�Epn-��q&�ۍq�MX��-Ƹ��p}D}�g�Xʴ�])���D]���_^�s�v^o�VWk	�d�F�%-pp܂
�)v��V��sv�v��z��uT��DG�9��V&oU��+[���a��k'�*�uAW0��=Q*m8ٟ��h�R[�z�M^uO8��Lv>nr��s�S}_&�zxz�d�\������I�W�8�Z�)�C��:Z��-������_����Nr��U.�{�}L��6fۃ�%mD����#�����i�-f�Ȼ�Rj�<�v�FW����#�ؤ����c��~���ڇ�}7_�L"u3�;2Gf���I�0����an�=w�^��;��M*��
��f����N��AR}����f�%k���6��C\a	g���%�)������1�	��e�)�5�.��@ծVs��U�Z^�����y9-��o\������q)�
m�G�7����v8s�m���t:�\���y��%F�&%�� )ʈ���
D�����"�������r�H-;j)Hhś�!tD�|��*t6��S�\�tNV�R���%Ͻ�|�R�̰���An�礇�^��PxL�I�{؛���ڦ9>Mr�t�8��0��w
��	v���������]B�5h�9g�m���W�_)���t�3K8�
[_�{/"^9�ř�K7�u��m��b+JRg�[�{Wu���q+B^���ڒ�e��ip�+��iO:է��粠�������䟧-{�V�9�녳)�ʽp3* ��œojV�_-�����dl��i��JgS=+G7�>�ݚ�1���,�T>]79uRK��C���%JB���A��p��.��<�*�)�<���<��7�>�Ts6�Oע^�:\�Y���߱צ�Q�D�$��6��/�o���Ʋ{!Q���x�����o����9Uc�����Tr��-F�߭B�z�,̻����w��UE��[�n��,���w0:�ݑ2�\E)Gw�_n]ڧ֤��G���XȚo�j4�F�
� ����w4w}>�֨;����aA�{��kΜ�p�Z��6���):n�N_/���:�Ynzb�,�Kl�b�ܠ��q����q :����N�C;���� �Q�5�R��刉]1T���Tp����\���h<^�嬢|��fgP��As���wCMC�	`fp�*���R릃qn'ǯ�d�v������Y�n֔uиk��c���B�}�}�׮��\���6��vj:_u����m��T�����o�5����`�<#3�JS�����;g�B��Vky��F�L�)��vc�q5:)��*��+�v��%�R�2�'1�UG.r���6ÿ�,�Jk&6�R��V͸�ך)���Pڟ��5/�q]�)}˨�rLL��lM92q
�W)Wp��q�L.��t��O�ܕٗ)��س:ic�Öe9�h(S[�ћ9F�aJJ8�8�F���s-s�K�<��/;~NEa����2H<�Ş���RgC�˽^U��k��g��i��e�M����8�J�6㵥�~�	�{
����V�@8۝����{�涻�b?Ei_v�q�zc�[�Q3&�µW�s�:�Tc�|��AS�,�����睛f�Γ��OC�9��)^A ��9��n�W���j��ԫ5�̏��J`N�B���e�53�{�E)���䗃]�腪:TU�v�y�*�Wc�g�Z�AT���1�z-�=3b��Z�`wZC`��u��uA�Ի��ʴ���u�]���kG��ڋ{:�R!,��`�s��6=3{ᘶ��>��c�e�������W݋e87G8sG��uv���l����<�a{֙m{�����{}��Φ֗<l�*��K嚺he��n��j��Fj�{y7OUx>&������[_&�ڛ�ql��\���>F>ܿ]�=;h���d���k�m	������KE�*KE����*�ַ`Қ�W�}��HT��uD�յ��͔�%�Oq���uJ{��A3uQ���mm)�["���cHN'���[1ۊ���W�/��P�}q�r�������u��:�����=�#L}5+^\�}�T%����y,v��n�Z�ꋵ�z���e�~Ȕ��B�s\B�S��j"Wd�'�C��&	��&໶enbwJ�=}F�L;��;�+��8���nk�����[���F:Y%^B�M�R��ݷ����J�|�Ú���7��"c���+L*�M-��n�)ɳ�>�^>wX�q� l�L�g���t ��j�8V|V\�N����q3�*��(5p����yG }��o�2����1b͟h++�ts+`�8
�Yc_d�Fl�
}�
�^-��j�����[.��޹h�LZ:T|���_W��y;�<�<�o�)v�z�%gZv�J���]��'�~Y��qf��c��^��k��VP�u6����~˭W���]��s�R�M7�5ܜoj�[�|��q�z}���U���}=ᕊ]=W��%��wծ�r����+��>������+2��ۣ�|=��En�W��Vpe�/�3շ}i�Z�����y�����]�����s�tܛC�U��Y왮��muo�v0zV<��MB7�gD�>nq�j��6j�߻ܲ�w2�tJ�c��
�n�L��:\Iݩ�N��)\n��V������Nr�eرNrN�e��|ڍ�%��#^�Ij��W�vs}᭼p���-�:��Z��U���^��d�
��W�؅o�Rv�1�Q'���KB��q�Z���*�
��Τ�p\U?��Tճ����B6�Q#y��[7�\��/�;˚R9@d`�Xp����'N����{��H���؝��~]������Y�.n�<,h�z�W��y�3���|m֊�F�eX�-e3D��bŬvR�ɾ����[����e��h̳H��w�1S�n�
ɥQ��Y�ǽ��[������ûÛ�ɮ����q=�Qm��T栩
���4�{5+^!�њ��3��[�r�ƭ
�&�7��fد�{��)�<�or�����I�.�-�NnMb}��.f�M�w�p�3��Snt\���{����{����w>nNY��S~\jr�KM��p��������Uo\�}]��7�6��mdKs��ir]4�7�u��k�9#r�<�.�J�HSW>s��,�F�"�Fb�y�`���?VU���إ��}�IyW7�ˊ;i���˞�{3�ܫ�2���~���{Q�e�PǢ�]�hw>�R�Co'3�����U鞑?5��b<�-kӌ�1�꼮��5�8ۉy�w����:]�OW��RO+��yi���W>[{R�̚];�q>����g��aqՅF�M̴��������GR�%�t�X$�Y���ռ�£.=NjgX(QȦ�Twf��Si�֌���E�t���������ZquұA�F��-rgB�o�n�YW�
琁Ϡ����ӕ�]��/QQQt:]uu6��kL�aR�V���{\6.�}���[��n�u�h8U��9���_L����Qʣ�qj>M>��;SX��Wax>��8��:_�sqtz��`>DwdD��t���'���p�0r�]����ɳ��3\�c���i��aR�د�p�ү��67m�~d<�{E�.�R��g<k^���eD'Mޜ�ܦ�	FX��r�Z�Ƣ��r�l�ųQ
Wt+}��{�����MCr|�j��q�*o �\'x)�c�$v>�g��
�&����cS{�=7����eS�M�Wzm����Ϧ�V�XNo����j!7��3l3&1Ƿ%gŹ�sc'�j�X*6mMG��m�r_d�bɈ�er�97[Ț�|CM���pؖ�F��+��qQ1����)��+�
w;�&��Pi�6�ȞJ;��Jv��:4��߹�k����bګK���U33+ ��X"�3�15!�o����r˲��fVl\��568=��"�{��R^��d�ܶ���C�D��МL��v8���_Lv[�L��uB��U��	���)j�A������֯'L�:4I{[�1^�:S6�
r�[�b���(���]y=���������y�����+z18fܳ�	��s̛��[���B���Vz����3��u~���Ε�u���o���{�	�N ꫣ������mw�����Ss�<�V(?_>wO8�)��O7���P�v��֊w{���`�
�ޯ�\�J�أ�0���|��x���q��=� z�!N�^��i�6���_����HzO9�����=t��[�*����7�i�|�Ψmiw�p}ʤ�r�ŝ�!�Zè]~o�#Y��VΫ��v�5��-����)�Cλ@���>޵X��z[��ֳ�%������:��%����5�c���N��8�������̦��ܴ�w�nA�b�����+*6��)w\o�!8�x͘��̕���n�3�Z�o�%�-�Ɛ�H��n���Х��ݰ�4��3|1�`�g>0]D�bЦ+�[xwO��1�ifq|K=Oݵ	����\ˮ\r���F�Ϋuy���}�i�n���f#[�G�=k�R]�+A�_t�9i$8�^�d�7/x�����zg�bҰ�y�U`.�0[�S,�h�'3���O����oV��b~���ܑ��������>]��=��V�R_EA��{cL�%�W)���6¸"a:sJe�q�mL�k�]���@٨��S����w;ΧiU�]F���w��q-��t�8���ܔdt���[<����⦊ۗ�'�c����i���qq��K���۩ѭ�
�TӅ���[���"�|p���8��s_<�;p��Ŋ�5�_s]�:-�|�^��b�Δ��]b�^���^$�k�ʪ��M���fp��C�;)���Q�=8��`�� f#g3����A���ȼH����0�p辎M:��"_��l�~ڥ䱚�im9~�J����v��o���C�	o�!�}��W(��m�D�Ϳ�ޯ�����\��v/^�n&�Wn5�sz|� 4W��.�����78�n����O_��u�z��u�8��ʛ��ܐ]��5�ѿ���k�����o���\"�
:{f]d�#�Υ�ZB���0PU$[���U+�9n����+	 �IӮ�cc��<�S��e򶖸	���k��]� �I}6��r&�ƒ�Y�Ӻ.��{�&"��g�R�7�����K�u�R��kwxᬼi�Ĵ���%¶����)�ˎ�'-��D��|����޸ko=����ٓ�Y�u�#��;���ï�}�N���Y��N������V!$��_v��Xi.�8��r�ҋ���2��T��8=��N�u�J������e*��øc��;�&'���}o{�s��<չ�{�����ߓ��s߻P�47خ<-bק�R�_d],��x1]��a�I4�|�lRob�ӚS.x���@f75�VF��S�qN�jwrj1��૗3P��ḷ�q)�mFXr4���7�s�SJt����ےS��œ��_%F�&&�q��C��Ea8�n9�ܗyU����5����W�����o՜���SO=��|q���tI�ގ�x��ܜ�׻�o��F�U�g�%�<��+[���>;�p�z�f�P}C{;��5֦R'���a�[agJ$p@4-�{�yD�&�-o�e��B�ZR`HRG*n�ۭ��g,3f�-��u+9���)t�`�j�cz2�Y����-�7^���-��˸{���eH4��G��I��|����0�Μ�70W��)ܕ����6m��k}��6xh���0U��U˕�9r�2�)
6jV����y�ڃq�Ê�����J� M�9&Ɋ>��-s�W{P���u�g=]w�{��)gN��Mt�L�����F1R�Y%�MR��֌����*���w�=�1�
��Z˫a�j����Xx��4k�6t�Ѻo�6�A�����N�{��S7�]�'��ט��������T�&�q�R}{V)G��O���;u�X�Z)��4�q��P꫷�/w5����
ʽ��[ɺE�i��*ՈuebX�M��v����c�Z��wkB�T�r���̇u�T(V��]�s��Xﻳg.��~|��+;�H�e�\ME�����M�)Wr�j���<���7d�)�:4-��ՁF�ꌌVC�7��<'�n^v^�1���(^v���1V�v�u�"�J�6�؆�Wl�{S�oL5����EO�H��8b;�Bn�UҏK�z]�;yOZ�;�9ȹ�t�Ae�~�1NI�Bۦ�����
2�<+3eJ�h�&�L��&P��!t��g�KIb1�x���d�kV��[`3�{�<��F%)JC���ɜ��Se_k�i�[��N����w��Y!��n��A��a�\�R�Z�rQ����#5AJ4�X�6��E*�\��(�Vqhf���<O�B�Q;J��Ȳ�>y���mgWs�����*<U��
�ʶ�c��C����iݠ\����&tڛ2ŝ.\���LM��u���5p�0θ���`lկ���Yƭp�x�F���D��:+�M��ʁ��Ww<2�5֔�̾�5��ыꕘ�nݪ�9߬G�SvWL�Y��n��L_�r�J=����/��9iD-۽̙Ԩb��-�n��<(��Q���z:�tIT��f�Ś7�oam�ț��]*g2-=����5��p�D�w��hF�h�,��-(^�X��\ӫ��n����-�8�<.�A�o:sT����p[�h�b���7�aKf�I[�����M��S�F�۷7@�Ѯ��V8C�]/��v1�^g1L�����4//6�^��^�]�a�xQ�G�b��Mdd��+��3Z��t���hֲFM�ݾ���7�V�Л��[C���f�88#ُ��0u��}݀�كYj4���If��¶�]%�Vͫ��\��P���S��˹w��D$���BN�����<mm��W��ڌ&�6v�����!��kO28�m�')�8'�W��˟Z�1���ˮ�|�����xt�{�q36بc��n�v
LY�[�Bd��yn��&佉W1��
�/F=��1<��ed���<w�����;��=y�#�\m�*��6+qE�I�5"�+�*��(�Dj�5���X��Ź�X�����n��-,TF1�qE���m�%cbL\mŸ���)ҷ3Wq�E�\\P\k��5�n'ms�QE�7�'.m\Z�\��-�\h�5kq����c���J,TFM���\nDۥ\U\n�Zu�qh�[�����cF���.��D���\����lV�rlln*���6��%qWW���\jK�q���n-�7.\����\lhJ1�%�n6#F6�"��"9�e�\j��nJ�QTG�}@W�|�h�`�p��G-�t�aF�e�y��݌�/���A�:J�$�Ë��cӭe�?d�tL�d�޼2&�ԱU�d�Sl��r�{�=��1~{.y����k�v��U6��*�VwW6W�ߕά�l>��74i�2�=v�_vF��usy�,��W"�RKX���2룖����ډ|:����p�Ϝ\)x�!<�y���8��.�]N.�"[�_I6^ok��Gb��-/W�՗XTLF�M�So�_f�cg�.j��C����k'���:K�u�"Tr��-X��s u�O+(y��:��m!�ׇ)�s�8컙A�����g���t]*��q�����eU8{��8Z�x�4�M�K�Rv�0W[W�+kip{����~�ظ%�e�ߦ{��z�d>��br�Di��ܤ��w���i|2���JC��^��<5q�^y�vt��>܆�E[cjR�nC˭6E�E����ÓN_$w�"���ġf��&����C9�7�(�φ���%Q�gpEa@_�o��X9]W���Ut#W��5*��#�Ѣ�T[��R�	&4�����U�]h\�������K����ၭ��o6��"�F�k����%�����H��J; ����NO��D*�K�w�ǵ`^3}��!x� �AyKO�L�Q���	���p�}}�r�=���^�v�mp��ʔ�ͭ��ȗ��|�������Z�_d⼌�V3C\V'�.��J6M�}���MƸU�y۞�}�l.�ϢS�fy�����)-�Ҿ�]5�*4���j#��k�����jb�;�#o=�r3�����>�m�q#�ʤ�B��m�9���s̛��Ʃ�鋞0��7����"nxM�S���w��v�ժV������{��5_+�ט)eޝJ��O
W�I�_:Q[[���57��T�)��9TaEP�)Ky�U��S����X��*�qϪÛ�{��t���Q�zx��eY�v�L�6v�Â��t�n�Q��]X�*��uW�_Wҡrrg��
��ڡ�(���j�:g�(p����O��|�+�miw�t��(OL5�i`��%eM��	|�����M>y�����Ʋ�@��Ksa�W�)͌,��ؘ��t-�]t�6�G^:4�7�wj�A�S2׎��t�3��Vf�.�Z��J[��W�2��6���\���+��kM37攟l=y�=�3��۱n��}3�o��j����=e�ж�M=�S|��eWиg�s%p�J�b�T���Vԕ�%󸤰�I�8k=j-���:nj�ae�͓����\d��f��`'�RVTF�sPR�O��N3vw:^OU��ES˄�*��u:�5�!R����J(j}7��l���R�oF��' s��u��ba�
��WΩ�)��#�.��ϰs���J�ܧ�a\O�ψ�O9� 7��6°�&�5
e�q�ԕ�7} R�D�CovyꝧNs^� ���5��}\L6*9Ӝ���b�ܗN�����We���D�ɨǝ��.���JJ14g*5�EPάD�����q����t�Q9le��y��͍Y1�V���\-p�yNvw�B�.��C�/W�Dn�W3�>�V�ma���=�֡��R®��s`)wƣ{h�����v��g��(�{�3xW-K��X���[�]�-/]�û���7�+H����`�c�u����i�Jg6����R�(Z�[��j�U����h�n�pZ�U���8L����j�'(i;�:��%�+j=��˚�ڪ9QW��n!�~�9p�0{�f*�����2�1@Km�x��;�������&m?�Kqj|���cg�oڼ�3��߇�N߰�-cdd���{ٞ�n�D�"��^k����'�\K�ۏ��Ʋ{��wW�XUG��4pm7t�Ν����D�>�����¢c�ss��W��B���5��@r)��[�\�+x�7�P����*9lb��kwxᬸƟ�lT�����.\��æJnk7vz�\I�!�!,��J#>��n��[�bA���y��g��HPȚp�v�B�n��K�[~��iT�NR���#����$�%A�-�ڦ�Z����{�3������0����V�v�K,LoG&o�S>�m������[��语��e�!Tw˧�*/0�94�8��]nR��k-�LGf�_BM(o�PͱI��e�%�}�*����a���� �n�E�Ǽ����3��w�œ��_��|">�/9W��q͡ �e�v*�/�B4�l�40�j�{ՠ�+����g$��TyY�*�ҟoXƶ�)[�*;)��ϵu*1�e1����:�b�yl�,Mޅ�؆LZ�V���J�v7| b]5���&��緂����o��e�;��w�Ut.�H�(X׏�uX]w���Pڒ�&�%<�ś���%F�bb`΍�)X��|��+7�����9Z��]6�_FS�̩X�1d�U���L��6�.��\����."ہ�	�V�#_����M���s�mg+]�۝^AEP�<�ƲznG����a�ѝK�<����D]VJ���\��YM�3�'JD振�M�ZzV���/w�׹Q�Z��H:b8��m�v�|,cf�����|�nr��c�#_.y�/'{�����C��(&$v�^�ǯq���ʂ�`U���P����
3y&�")�5&��X�mW\��ڌxZ��3�{�bW=��t���d��P�UT��lv�,��c�	NY��W{ކ���~����U��`�*�=ľY<r3u��}S:۵�����"�0Z��áp?�EY�h��K4#�����wl����b���"�[�:�m�TD`�W�r��_[:��jS�`�Y���lɲ�b��5-����2:}�����vA����P�߯h�B�q���,�(�JstY��Ko{/\5��g&��M��
�po���ĸ�S�����x�^���IŽJ�`����\�^u�����K�T7^�U��=��J[�2a�_r�;l�v=�R��}���lf��;l�x`�$�hnc�\�w��4��BƯ�b;4*��W�y��v-��Y��{�T�+���c=��E��'L<�a{��ne���ҫ�\��ZK��ң[Դ%��p'�3hu��?'LT)�;P_M���~ͬ�Y����R�v��ܝֺcT�KU�VR�Z�K����6�\*�Oյ=���}6���m��wOj���be�5R�vf�,��F�X�M6�ms����t�[m�4�;�l{�T�s:�j>�/2�������Wz�6�����cߧ�K~-�\�U�5�p���{�Z��t���3���]�կ�L���֟K�\E�lsj��Z�qVT��Bb�af�E��6��W�B12�ʺ
�#@t�2e�μv�?�e���SnR��T�\�,Τ�Z�2�oɪp�:�쏖Vrĉ}]�CTÄ�o%�G) v.�)�qX��׻��F���icWY�R��;�OZ��ى���-zrX�r���x�.U����5u��;'�����A�>jh���6p�w��r�T�V3�+J�MXr��TJ�Պ8��H/��T�^��^;WS;7��)w��U�l�Վꂮ������t�h�ˀM�8h�{	ň��o"�݌�6�|_<ⳛX_W�����6��=�q���)9��nc�qJR�-��է�mBi����\��J��Qzb)y����Ψn׾B��n��;���I��8km�[Qo�<�� 5f{T��U��s������!�%
 4�$����K�=��jFw���m<�O`��m�Ιs��u������������ŁJ���u4sm&��q��Ԝ��>0TBle:�!���#E�L�P��=~YCXH��Y~�ۊ��imsJ|��"a:sJe�G��V��{��՝2OrXVJ.��w��E�Ӹ9p3��j���ָ7VK܋��+6Q�ұ���7���T�
�Q�KJ���:J�H �ð!Z"�s���<�1L�ݥG|pV}9ޛ�K��Q.�����\ݝL,��ה	y�&CҬ�o�2�;�f9�ɬNs����Q�h7���������T��9������ӧ4q���/"yd�,�v���K9m�4�Z�e���+�q%2���stj=��{�mny!��q�H��R{a���M��*�kݜ�"���unC�;)�s���TF�����wΔ���.��N�uh>��ê9U��mum&�t���sq�����~�9k�3(��b�����k��˾G�\Ǝ���BT���C�(E�$s�_���땥��U�r���i٠b}�3�F�����}����M>ȗy����Y%i�9��#fR8r.+�S�u�NԸ]C%��Q1ع�t�/�sۈS|_J5f)G<���J�Y{S��0_@�q_TJ�U�)J5���e�4�# ������uy�Ez�%��+̓!�P���C�Q%*��_ԤOg7:���f�]b��fQ	�>7�z�.v>x��y����L=�����(�Z���kŜ�+u֪u}Z\5�	עg&�7 t���u�t Ve�+�%G�h��7(�V�˱B���V��mD^!\�A>g'f�}��;N���(p����t��xVr8��.�C����m�\�B�l񶷫����ޯc���n�z(-��)���p��D�O�����4rс�������>�A�V�ʇT��R�~	Ge��ZJc��k-R�Ae���k[-(w���m��uNh��\��voM���tw_1.^�Ok�}��BM+���1���e�_\U'2��92fq�]���R�TF����nMbs��W.f��7��̸Ʋ𮋨�{uUb	����C�ʸm�7�}��{���s��j�,����N�E �b\� =Ntʸ�sM�0/}���aNk����eD����ٕ��s��q��t�z�ˋ����rY[N!']p�Ú��mBs��,�k���T�R����n�P;�ߕ^�ut[��ݎ���]��'ޗ:��k��E��O2\��&�c��T9�ʭ�7�_K���&ޫ=+�z�K��{���һ(�ש-�n ����5�t&�]j�O��[�i�k3�;w�\� Ο��t1dK�i�̯zb�k�ϥ����&��ie���v�r�}�A�fɶ�O���wr�L��3�ܒ$d'����p�Zi�̱�1nDWv����X�/���ǲ�s�':;�<��U��z���3����wݞ];Ŷ�{~cpl����%ltGN%R�yV��~j�9�Y�騸�£y&�$���Av^(vӞ��U�OV9o5,]�O\W�u��������ڡve�EENv����YP��	���w��r��8��.�|ޜj�I
�h󊨕k���lGjp�y��놲�-�M=��M�zl*��!�V�1��G1y�Ր�$81K�N�j�MAI�;k^���e|�7q�
��Ñ/,�ީ�ό�8��E�]�!���Ϣ���7�-c"�N�Z�s�{H��/��h%5al�hU	4�<���1cp!Ȭ�8��m+ǻ����K9�<��;_°��jt�.��/����N�w8�G[��̸z�VͰ�,�N�F��q��Sk��}��&nYq-��C��!'��N����l.[V��O��^ɍV�������;Y��\R�5q��E�_rf��I$��Z'h��N$�}{O���L<��*ƻl�K-��>�h�I!y�Ԙ��O��ҎT��En.̭�SD ��汚�ݩ7�Qo�[R�ƖQ�`�X�u��{ڈ��.ıhg�ޘ����MKwl��^�ȥ�=�����h��Ӻ�7up�IC�+�>�(P��,ͪ����o/
�wJj�A1�Z�ve��]Kn.�m��yX��9J��ո���5���6\�f��O[�Z�W,��=��	E|��q���'���Y�ĎI�r�_S+,�[�qV%i���I�|:��Z@�V��v�*���
�WY\��Ń���[ܕ�1�"��f�Z�lir޳�m*��^����@��I=`�����4.�v��7��Z�R(�Ck/$����/��fJ�*>Z�o�-7 ٽ���|L��C]�+�MZǘ+����5�(�N�n��p�;��'�s��hu��v2�ζ�̣9��˕s�}�%���:���7�Y���C��7��%���aw+{t3û�J�nwS����|m��Z���iLuY�Yi�7q�G�ڼ�}w��C&��n]�v��ǘ���R�Բ�$:x�nM_<�,fm"�oyV73���
�ň�-<�^����=l�c�Wx\�t�����Ε���a�,�Hn���G67��һ%����n]p<����hj����G���
{��]l���k�6`=�vo �-�b��.��Mƺ����˦~ˊ��)��̻����u�� 6��Y�c#�j,��J�c�lL�x��\U�z��p�/�,N�w:��*����i�\��5i��}p!�]�ë�&c���=I��1��^.E����U�:�rn^1ݸ��.����41�Q�_P
�R��x���T��>�XC��e�����g���9R�#�
�� &g�� ;Ұ�q�ڹ�����MV�mR�¬���k�5���4w.Z�11�6�S:֮��P��0����9:��m`�k�#J��bau;{(r�bx�Y[��/��%��J��:
�	}pҌ3(��7OU��uc�\L�{�ӻ��Y�uoZ�(sl����]�m�����!R��jLͷ�f�PY�S�N칏or��b�P�]:wk�ڹ�x���<E]a�x��V�B��Մ,(�삚�VXطY�R��L:��b;����m�iXK�N��һ��/8����Z�3�������!Z9�t0�υNG��{)^+�y��O��{ӧ%����W8z���]�d�YuN�do7kx\Y:2g=�7�v,���^7��{&��5��2�i<nS��}�N2�ԝ��tח�p�L��V�
,��
¶^i2s�)��}ӷ��A[��hYխ^��q>���X~��$�CEƪ`\e-D9_�׾�y���j(��s���1��7"����(�6�$j4VH�ѵ��n)0��1�F�!DQ��s�����E#cHV5�r�.s���h
(��W�UB��r5A�.s��4D�,���P�Q��rC`H�DHE4m6�ےM#cF���\�B��hZ,j4d4Y"\�,Q %.M����l�Y�qs��\HQ�J�9Eq��6S
,QƌTQb���K���1!�#LdHP�(�E�*H,�=w����z��z�wϞ����;Rqr"/oz�d��O.��8.��uj����"N��&�\��FR?-�!}���#k��bU�E�D/���{�ҫ�K��G$��͸�q1�*&9۞����آ��F�P{�+�lp�)��&��{j���\�5��k����dc���i^�[9;�Ĭʕ�n5d�]Z���}q��5n��Nv:b�n�`���Z1�{54ځ���f:��}R�ebsYZ�:e`�O�d�z�9�e��ֳ��a'����p�������Q79Q<�Tb�|�����a;����g���g�;|k�C�H���?O(����U��Q.r�T>��%��YQya�JEo��D���E��ڧ�m�kg�*�us�:��-���Mt'��6�J7�d��Q�؋s&�\K�gWͭ.x������:��X���p
�3s��┥c[��p�=�M�]�:g���ust��N?���`�ʤ�Q{��Xk��p�<��5��Ko��2n�Ԏq|��,����5����|�i
��uU��A-��}O';4�gZ"�f�i�;�/���J���[�n��̕I^.��\�>\fӭ��4���=17M\��"�@ܘ.�w��G���S&�}�лCz��VD�ӲDsN����u�RvJ$4�$���l�K�ba:��c��f�Q<�/���g��'���9�8܇P��0ca(�����]��!N����S���qq���7���_�	�z��Rt��4����B�v��Q��ͻ�ά�������K���|�6¿�ȟ��5
e�q��7��Xj:<g,y%��w�w��f�H�W���M�0ḷ
�Cb��@J����=�g��җ�+hm��̿�<�W�v�w�Q�X��6�]��%R�����J���p�eeHlM��t��y-���_$syI��D��02r��,{[���ٌ�v=��7_��J'�-����S�Y[w�c�u(}�\������ۈ~�~���~�K~�U�ۇ.��Y�np�W���P���o_ǧ�\)x���v��wk:	6�Ғ�<��Y��w/
�Y��A� �8l��r�nY�׻�#kN��u߅z���꽫sض;��n��4��������T:�5A�Ńt�'Z�-w4ļU+$�Zi���N�:�/u����5�M����[�ԩo;�3�:I��sT�r1�z�a�c���>�|��i�C�͸o:���u�t��JчZ���.���9c��ɹԺ�d��¢~�\��;m9�k���T��^y	r���f���Yl��=2������1JQ��F8k.����TEE��;�u��X��q-��|� m�_.��ϑ	o�_)D;�vހ ��n9���7��㇝��[nm��6|��'`����}M���-T���W
w�)�V:��P��\rֻ>��6���&,=_r��n�P���)󮋜�y/��a�of�l�|���_��!=�V��2�"�0�f62�����l��n EF=��z����Ъ!&���6-����KY��j��a{
�J��;e��vk�}B5k��%nMbs�.g�|7�dmvG4�)�ܪ�[7��<�҆|�����>�RV��Jy5�b��x�U�ʖ���B�Z��(�|� uAX��L��1�Hr�s�ś�N�'V_�ڈ_N�|�R�sV*PU�R�!SF�һ6�9ݱ��'.��e`�jj�Y�:r�(�I3��fb�e�M�-���� ru�co9<$�j_T�B:v��n���Q�j��;�M���F������ꭟo�ڬ��+��������vEY��+��Z\�z�sV������n�z]�=�ލ����rAZ����K<������j���}���8�p�\��K�"鞡wA'Q��5��]�)K��[S�2���z�J�|�����������f��B��⽜5�����|�&�*S�+������[�{|-J��,畊�wu�䪱�{��m�R�����K�_Ժ������}���J'5Z1�c4f�l��3����&��_f�=U�O]p0WH:�}���������E��eTi}�����p���s��O�%��_j��S�p�����{��w��í}��-R��g�t�X���5�Yq��Bi�oE��\	��B��:�]��L�B��3��|�Zɯ�O/�5υ�G��e'M�w<�z�$�@ɱPԎ��uh�1e�����].��Y7&Εҋn⼲��͝�*�B �(��nA��S�{��J[ԯ�_7D��np��j�p�(%{Ҙy��:$�b�X�<4L���]F$ڶe6e��(wu��Bx�ã'Q�8f���s��"}f�����ϧb��{5��q����Dn�(n'��ǅ�7Ck�7T���*��S4��`,j���Щ&��{��!�9x;%�w�tզ�`���*�k�S%q�F�}7+s!6��г���OU�p���o��f�vD�t�)�5�.��+\ȃ�����r4v�onZ�U.!�Noˤ�$��n5�W�u�~[��@TT�Mk^X���o�����r���5�&;j���_,p�p6���~�F�U����N�4g�x��UƷ�K�U�Ks����g���U&z]��ߏ����u�9�u�Q����U%Z�>�V�oՇ�r�{�qwL�V��[AҜ֣��uӳ\�ʡ�V�9��[�U�K�Ҿ���p!,������`u*s���̕��v�l��gz����)ʞSW��k����Xss؅T��h�����=�ED$���h�;�|������uٮj�X����y�+�W@mb3�e\-�֘I�1�ҥ�p�qȸ93M�+�+�`��~�ƾX�o���}��v�����s�.��fW8�7	۱��;t�.�]-���pBn9]\�#�*yHug�.q�ڧ�ݮ�kg���uQ�:7��X��|u�<�Y�	�Վ�6�g��҉��[�M>�|��+9�������:'9FL�������4{Z]�*�.�5��p�[���&���f���4L��'$sSy���R�ߟ-�JU{��%������Z&�i<����sr��sH�]���'�¨_r���	|�Ϥ�:�1�0e,��)��=]��^M$3~�ٛç�!HU�YV�L٢�!����yQj�ʷY���ZJ�K <�_&�T:�4T��.���VZ6��A�����r�̿����V�\��o��m��0�9D�+9�T���<q��z���p2�]9�&���l��0���c�
�ٺ��.���5T�XU��}<FPYw�Jy5�'�׎��J�B�W�v�b�7bm���ѩ��,JL����i�L8��y�m�խ���A��W�}���63���3��q�c����c���x�csT���k#��J�;�1�d���h^V�iŻO���+=��Z�ξe.T⤄:�/�{��T:����Ga-���B2M��[����9���xb}F�T�+9��uY�9y��˫Yf��#�.�[�����9y.q3�9Ś�p:E���f*�m�D�ӽ��5��@�s�y"��Qp�j�=+/��v�\�nT?c����}���^n;kr�7_!��5�:���N&�eDc���kyGD)x��ݸ����y���ۦ�Q��������+�޿�V׫u�Q����)���6��t�o
Æ�s��^j��94-8��`u��P��d��*'�ss��Ù���g��f�k���o?���K'���U%�DJ�U�)JƷ{ј�B�ڜp�X��ބx��LLӈM�����|��U��:N��N��ݿVNҚ%Mǵ�/N8�y-�!���᭿��ڋ|��o�M�K�Cb�w����e��n�w�ӓ�n),5�����mE�1̥����C�Er#�D�OV�DxI��:�V���*�(̹ic��/��N��������MJ-�;�0�x{�����}���y.f���� N��S\C[JiU}K�.ђ�X㷊%��EN�_wj�O�a8O[���4bg��-��X�?�Vr�Z7��գ�5N븟D_r�:�_=w�;՜����D�f4,s�uEC�4;q��M�;��w��#HOd�wv�%�M+e�l[���+�Ջ�<���Rw=P�^�jͩ��>��\ܭ���;x*�\��a����\���u=Njg�P�A!�z��NXF��G����V�ԧ�Q�9p�3/;�𸹴�7��m*4�1-���NV�5�^��՞���"N�OC^�!�z|�fS��R�z}j��9f�:+�E��>��C�:-uM�i�����]e9�ʉx2�˚Y���k���0�ܬ|7����w����H����թq1���ڕ�*1A�z�J�|���}/�V^���ۧۏE�
l\�ji�����\ʾ�����b��\(����7����*9��<o��������ݳ�C�*߁ީs�*`qҎ� x<�.����L��ѭ���H�j8��[W;#�P�}��H5�v����a��1u2�a��י�QH�s�ɲ�m�X�V��z*�fq�BSfV�2]�l�>NVr���Χ��e���o�͈���t4�6(]m^�/U��oh���+���y��ި�ٷ�=U�d��p?�5_�_Ӵ����b�=*CQb6��Ά�.v�}q-=���onq��s(:����zV���s���DΧqJQ��7��ˈ�i4�ʶ�l�peㅜ�5�MVb�@c5�1P5�����Q'��O�mG��f��� f6��ŋ\�ʩ嗬o^8g�_r�;B��-�L7�/<�����oKe�bx�;;S���V9h��Ni��_5���(���[ׁYŸ��I�Gk9�������c9��M�T|]3Jd�!v����g4��tw�󽻌N�^�}����9��pͰ�ȘN��6��P�g�L�����	kβ�$:eľɨǓ����v#�b[q��+����6�
�+On�E���0�w�ܕ�<�j1d��V���Ec�<ہ���SE�X%'u6�Q о�(����{�۵���yَC���v^Դ^�oļ�`��[�c+�Ju�,	�|�Ω{�WT��v���ku�V4�R��8�ZW�:S���0�B���5�c��o]�-R��Q��ʙ�v��v��9ϨgE[^�V�-�����R��]����]��y�=�n��}���z�%��U��Ok|����-�yS��~�^���*Mt�m֐�Pq��}.u�^��d�X�uG���梶��P��˽�J~j�Co5_ǧ�YO'y��;\���r��)FN�ķy{��Jq��X�(��|��)-R�5�U�c[=tnCާ�W'�-�<sO����Y�z-!���K끊'��E��������o��*�
�+�s��*ޓ��\@=�X�3�fK�����tw�cu��%����q'����+�pl�(�,5呾�3�,�2�.��t�0�(�f����7��-ߴ�n�� ���SX�g��Lk��xhy�1t�S��0ω�1�*$����أ!��;�=a�{0wqڴ׶��ı=u�|�3�o�Ŝ����ӥ\U6�k��<��FH��#�|ߢ����_��K/�W�.]��貸I�m��]r}���kj��[�L:3%iZ�����H"�c�dAZ���}�K���Z�{A|n<�9X`Y�̪u>]����Q�7�L��4�̮W���4�\�FIՄ�y�mo.��:�����Z�t,VJ�+��[qipu������կM}�t(�n��i�w*o�^������e<S{ЙSqYR���h@B�P	���-E`傱��e��hq��]�^�q];��穼�Pb����S8�˗i����R����bɑc��;BpgpW;.]��!��oog6c2��IQ��rE��Y�(�$N�y:7u�ʚ�T��k]D��å��↡���v�
�6�B�]�Xb��C�!���֗s�Y�;h��6�z=Csi!�@�Q�/z0�]rz�F��{���W-�{N6.�`�/ Fsa�Ң)N�9V[�@]_X��ȰX��i�;���j��l��YS�ײ�&h	W�+T�{R���+�7A���u��e�]�E�`뮅��֎�s[B�����1��K�9��.oN�[dNξ��Fڵ����u�@�j�_a�zEvji>D,A�"�SsZ]{���%Q6�)�� �:[����>�J�t'5Z6�=V��T���:؏tU��C �eg57X���ї�ڱ�oV����u�:��S]kT_��R�}^7�^�2����&]b�(���goZJ�S���;�3%ɷ';��
�;y
9���h�f��/h&�;���JܟwQ�e�n�zI����Hk�Q�U(e��m�&t�����'j���[�gA��9t�@n�9�۸!�h���K�����q,oG�2I��rC7��+sr�}ۅ�W�r��'�$�ݶ��Z�"�÷u���N�;�DH�K=��@�Z���v�����N��8Z�}�,=[7�d��3-�ac�ڳ��)<]X��րnA6��x���zZ)e�����0�X��{�p+�[�t��0c�D��%�_��י�P�q���\�mkF��M�6Y�V�b�WbչC傲�'��q�x�Fc�B��"�8Q
��E���(�Zr�u5U�`�SM�@!��]ip�V(��Ϯ���� �h��u���*wR�M���x���R�ٴ�B%���l$�9�ޤ~W�.�U�M���ct�:L�Xn��T��驺������L\�3�.u�v"�:�$�rU��:s��f�70���j�vxW�Y�*3YcNK41��
u�����s�Z;y����ۥ���#%��.@�;67g
�oB�	�t{� ]]����S� 3)�V�L.WRN�6
�MR@�g2rp��*�m's���g>=z]�M/��¿�uwb�y��K�zfWkP���>\io
)��Cr\�����(��#��:�a٬�=)A�ʵj��"�7T
Z�.�+���E�,lY˾� �   CE���5�P�����eJL���QQfVB5��K%&%�!d�R�2`��9�d�(��0QEMh4�1�8�X�L�I�m���bF6�$i1EcF$� �EaLM�&��"Ĕ�$�!��E"�b �m"	EE1(�d�D�&TY�BEh%#%���"Y1S(��0��h�(�2%`S(I�A�$X��!���FL�L�"en9 �/�=���u��_�wy
̤#���D�����D�%��Nʠ�._t5�ñ$�H�s��(sI�=��E�]��(KS0@~�bU�YBj�C�̜�\j#=�����ف��l�x���7N��QS�5��1�oد�5��)gї僺������s�*+哌ߠ��uH|ڿ0��ώzg<K�ꍁO��/uǏ!	:>���M�k>|�ɓ�'��J�tn(��W,{R�rj�E��%�C�oӽ\c�Lx�5Y�ƞ�o{]Rc��UC3���1�b�FOb�>G��@Zgq�8��U&�d����dӮ�㞳����/Z�ϙ��2�/M��ߠ�v��Ԛ�3e������x3@[��+;�P�䪵���]������+|�FP֣�5X�Aҁ���f�����Q�����B���v\��f��E��Pu�7�N��#�y���<I�� �Wi���wƴ�� ��?��}���]v`~򭚜��I�cS�r(':M��Dz�P�;9�#�:�>nTfz���V�t������Ƣ���O���{�Ņ�Vi9�j�i�0��Z�/d�u��[��H�u��E������aN����0-�R��G	H��za�W����rV6�x,��Bo��){�����&�DX��&w�=���JaU7�Boͤ#u	�T	Y��nZ��X"��j�W]��J�R�*����<�m���|;�}u��4�Q�$]��Ci<{;�eq��=Z�ʺ{t�Sz4��j�z�첆��3d[Γ��u<ջ�gu�k�#��9�P>C7��9����۠��J=%���H��H���}3���W'��V�Ŕ�a��=����Ɇ]�[��f_K�ߺ��q�侇(UD�S>���%@�����Ҡ��c�i��%ACm�e�,����=C�C��_�g�x��`&��"/�w�����<���.��L���[u�n;CF'޶��8ug�@�U\G8��iùlD�ʽ��ˢ�p���� \���_���;�1z�xz_.��WF_��a4<�gﱘ��ǯ����--�%��<v C܉�Ȑu�F����pL4���9�;c=>�O� =ѥ˟W�S�����<K�Ȋ�O�P�S_i�{M|LAؚ4�a�V�2�����w��o�5}7Q��
���p{�2�D[��W�:��i�Iy:rj��p�O3h���k}�s�*�W��j��X��w���M��J5�mDc3�1F�C��j\m>�Ի1�*e��t߮��o��i��T��B��A�5�i�KG��9�Lz��4�'~��w*"���}�[�4���MLa���.��;Qݧ��Ҟ3�u3;53��G�ھˮo�Z�E��fH,vG$��(��+NIewɗ�Osq���,o����=qu��ᖍ���P���F��\�i���3Fb�PE]Ix�������FF�t�����!��*^��zt�҇��˼d%^Y��Q�}��L��yAB*��O����XV�n���;^�����Fc7d:��n)΃�,���c"U;�S�o��0��#j�t�<��0C�9��K��W����_�M�w@��^����Vid�Z�b15d,G���+�ѾvG�WJ_�xw{+��:�+"�	Cne��Ey-3!�t��`�g�����r#Xg�B�u�e��6w�=�y�y�}9EjI*�XU���_������4�5��]"|c�X���{�Ƅ :���<�?���ݐ]j6�Wg"ԐUZ���^��sz���B�A�Q�''D�|��[�7Μz4ct_��r���<��{=�j��A޷9�k7�<=�\�zp��g��|��f����-��"���z<����:r)�}��Gٗ!߆�)� ��~�p�8�n�1�&t����Q}�:k*������v��w{�tgj%eh�zs�?RM�����6�sC�D>�	�2r#��ȑ�o�v� �Z�hZT]����f.$��G��UfA�^�W���h[�d�f��ހ���4��0�/�a6�5����ط�1u<���#'A��tr����&�GW���ښ6��KcC��U�[ ��n���muBhv�ے�����6���U{��pM���V���˛��g��89�Ȋ�349$���h����5|=��y�A�$O�j�m�f��G��A�+�
[�M�/Ig�9�2_�r���5L��^M�fLv�{$fI��os�=�Nj��u���';eU˲��jc�{j����EnX�~�C�g�Y�S�G�����ebH-�*.(��G�{��lE9����j�dr�܊�j�ˈ7�;#:(��	������&.���hB��;@EH쨛�:\ߍ�E��gS+r��Ī���v:���p�;�v���sn�0ϟ��nhr�eн��mA�=5�C�/'���&�g�9���ʼ<��O��yB��=������ٗ
�<�\P�jѿl�7Bg�P.n:����#�ؼ���Sn#Wy���'9���旈�q�Q�q�!Vq��>ڞ	Ä�y�Q�xm�[w�{>[��1�>G"p���.#P��!f��Dzy�gZ�=x��*�e->��{~=6![�^��l����3� xeL�n��U��|"��B|]8\������4��ȃ1um�i��U>��Y�R�	jٝ=��즌t�L�����[2�g��´�ի"Re�ٌ�;�1s-l\�t7�u$W7���ry�D�X*���1�$���s�;�i�M�4KR�qW���)!�R�Uf�sl��⽽�;ԈԪ��c�O�Y�(��Ǒ�2��%#�S��}n�0�{׃}�����W��Y�n�{EQf7��p��R vT�l�K�3`�T9�$���]�Bo�����j�Wc�}9N����<#����b�I��3�{�DoI��7P#ŲV�#�D׏�.�sS����=e�̺@O:�>����,�}��ŵ+��҂�}�ƞ_	��US8�ʒ�[�Ԙ��'wK��WӐ�p�n,��k��.��\ݓ͠}�:�eEO*,�Z���%�:�Y��a�����H �SB�+��;�v.��W��|}�e�|�|��CB�v�YM��#unɛ��8'o�|�b46d��q�'�4k�Z٫��=Q�\�/��܋�7^'�H�{�U�5�vteg��{}~����]�wz�G`����A}=���s>^��;��'Br���dZ�y���x�S�Y_��3yD5@7N#��*.�غ�h���;8�w���}}�3���z�������n�;E��P��K�5�v�¼�J3\�L�Ƣ����f���{�R~^�A�SE�h��[=�PP5 ��i�=׹4�P��X�'	�s7���MV��TG�6�-a���.���>{��T��Y.{�	�_�#�R�)LГ�Euh����P{�뻫���]n��k�ϗg0dKz�*oE��]��LwT�P�w;��q�����}d٫8ʫ���������|ʯ
����7��N�֜��A������{�r���H�@���(踮���ˈ��y���ս��_|ܦwon�����������R�Q�Zxa9��߾�X�ɭ7N@��v�������ΐ�����a��w��\�����ӊ�)i��|N��$w�ii��@j6dx.�.��Q^�Ui
����N'r�{Ҙ�'��gM-���F���9'��:�P��H����B�~�Pמ�.SP�VgO�({*Ϸ�<^����Nz�xv:�A���.ܠID�ʡ�W��E�7�5#��/�8{�;��Sk����f���Y��,�f8�<Co�r����>�͸ 'Zyr�}�e,��4����R������Tϟ�-��.]!�=�.>��M��7@�U\G5�����rͪ���qe�_���@�FHy���ײ������Z}]����6�	��};Q���|�N�k6Zut&���t֘�,�WQ���>�0�-�!�o��?}�`������+㱞�tD�g�י/��Xs;)�^R�����8.�Q�`�q�X5�b�MAh����0���G?}�rQ0m�-R�{�m��5��ڳ����	�5!BٔR�|5՞Zc�T��*����G�.�A+��a�a\8M�]�\�t�fK�����Ǜ�����'[��r��I544�=���2bh�=��Z�)�ױ�uJQ�_R�i���w����F�6��̧�O�/�S��4ԍ$��95��W	aF3�{�w����Nh�,q�(^�C7j����%m��~�9(���_>^�.s�s���=\��{%f۱~��4�{]
�z�����U�{��ѯ9pr�ҋ��G����"��I!��s�-d�q�2��Ò�}�n�v�GG���j1��,��ɘ��˹�u����
��wK��n�w=���:}/DS�o� ��u�T��O�{5F�^���9m	]�g�=����.5NuuA&�~3�
rgN�;
 $�،���mG���W���y�Jf��Ǉ%�N���>^�B��:�+".p�6�eგ6\Ν��I���^]'�$�8m9�'�o�:���������=y�<���"�Z�J���U�.6A9Qg�'�m�;���Adƹ���3��ηR�#��9�:�<y{M��+��V�˖�<$��*�W�z�.8).w�\��n�ڷMJj�#��M��gf�S��q�7-�%�}���ӸdM$�R�b����>��D���v3�\���5<��z9��ҺRԴk�{$3i�Iad�����_r=ܗb���.tAi�.�<8�����`��vv�Y�6v'+��� ׌�3Ǆ�(uT�晐��<4gz=Ln�C:��ǻ�t��ڊ��l������|�l<���Q%ў~"E|}-���P^�o4H-��w���Vg��PfW�0߮��j-�o�A�i߮=�v���Ȁ����,��PGaͷ��W?X�z�|��-{�^����4�{M���^mƒ�VH��1�@l�P*K����%�������%��T�.v^��GYŢa$�#���>����y�q�j���rJOER{f"#/OuP��9u��=qW�=;�MB`)���en;{SG~�/Ie�L��9\B橓5-t�2"��GD<��6/ܺS1y�b�\�hK+ll�5���C�M]ɋ��M���G!�_h��m�ț�^K���.� {��a��b�%��N}���6�u�29z�C�H�Ot�$�,D�L�Ly>~�:�����,~�'hEH�"n���5vi���b�W��ts�n>�ڝ��ǫ��[�P���j��O31y���=�A6�}Mv�W���zɳ�k��^�T x�^.��jX�p,3jt�b���Y��=w�
��\�Bk/A����}`��e��U+����E������f�p��U�%�|ef���ݜ)��� ^N�ܡ]Q�b����|̩i�j�����"��Q�ǟ_Fj���HQ�nKqԗ��Y]��'�y8�|��c˯Fs�h߾ٸ6n�{� \�p�~�SZ�9���^O�oZ�1^'K��'��A�zV��<����t3}��a@{�ڞd��4=ݕ���3��4�(>!n1��Ѹ�����z#Pz�,�Zȃ�6s�z�盫�=Y��܎~D��c�*;x7aZ�j����@ˏ(3����zh.�����/�D!��Ӆ��s:�֯�K8]��Sg٧LSE�f�װ�oj�U�IU��4eSJGj��<�j:;эנ壻�z�lC��Hia�c���C��^[2�x�㤞FF���P�����f��;qSK*�5��_�׋X�ֳ�8�l���1�|�L{u~ϸ��>r NjO?�N��W��שꪵ����3���on&�[���3�ls�������t����PY�4�ǋG\	�R��=>�T
{����n,��ܝw��+����4>���꩕�3�7��Z�l�KTU�Ч7��#��	�?)��N{�p��c�wm8��y���ݳ�~�`��*̈��c��&L`��XOT�=@t��L���}h�ʇ(�,)hՀ�G��V�|�J���{���jp��\�[/�=j�]a�ɚ�]wF��p�y�I�%�[Gj�����]e�����]d�lyIWU$���{z��2��ۧ�&���������l�꣣'4]1�ut�SGI0�D`��Ѡ�mʡs���S7��a�pO�Q8f�w$U��<��D^�GP�B����SF��$�5��A}=���f�Zfg<���8�/^_��nڮ�xڤh;j!�n�F�f=a�]CZ�ڃQ�b�GZj������9��,���6��ѻ>���/.}��Z|;�hӺN{�(�֣�5X�AҾ>�P���(�TMN�su:3a�'qL/,����6j�e
��t�����}�Ĝ-�²�|�M���l�/��x�2�=�ϖ���6�Ύ������>'t�62��gҩ<��Ռ����R�J�p�rp�?J�����ˌ~���uŌ'3`�~��X��&��S�<�#i���l�/`��~����jf�EU���`�������S�Ao�]#�Y�R�0��A��w^�F✀�l��]�~�ܣի�vq�ź��e��N!�b��_���� �g�,��U�.Q%�ѣ*���gȹm��
��3�%Ώ`z)�E��,�����|��z�n�=� 듌�ܽ[�>���(UL�
>ܱ���=�Lw+麽�mN�v��&��=��p����{b�w����ȶ�]C��+gȫh,�s�	�4D�O��ЛX"�ñ��L�Y�pZ�б��1sv��A�C�)KH�L�c+��*��T��,[dQ�wq�M��;-,�̭��u�ōLG�ݧR�����R,�x!R����m�ջ��ބz�:�fTV�`�M���a��y�"���۹&�v�5�}ƅwE����]�n�p)U���6E�&|���[��䶉�i�p��lI�&���ˮWFbO,��dy,��ʄ�����3oWd��pP�5����ܔaV}Ɍ�1�cZ�=H����ͨ[�q��(:�x����.��r�/��Y�����qָ�ƲP�����D3�����V&i�
�_2��k�	w�M�%����f`��W]p^�'l�,t�B }՝��ڢ��>U��"V^��5pLޜdh�Lf���ё�ۀ}�Ui-�0L�І9r��W���Avi���:�A�K�s�a�R�B�6,����ﬦI�757:gu��Q�}��i�9WR�%�5�H��.�8��;�wC5�҂%�ܣƚ�[�s�V�T�Y�E�m��!��(gCӞ�E����%�U^$Ȼ���q�j��	���hb��d[��On�-��vq�K)7P�-�e��7��v���[�ء�����V(�x6�)h=���C��RY^���Wo���F�.ƪ�:흆��$�"*�Vge%V�6�����
S�z�*��,2�}�ɾt��;K�uš�YɊ��Cvwܩu�wD�‥�vw]�Ɇ��K�t�a�T4��ԫZ�{���L�ݔ��.�ڕ�q�Է��@�Pc�w%�V��`S]
��9gq%-Y��6�]nR��2��ٜ2�*�YI��Iv�4�E45Qg+k����f\�R$.��nnh�����#N�$dl����*%�L�ѥ\�SK Kq����g�o;`0#/��ІL�V�M���,C��;�R.�fE�U�ꋣ����/��Ҙ4W�^�Zh ��ݥ�����#lb��v���_r޼r��'u���K�W����G�l*'�a�q'w�;�s�<m�|�zu(����	�p����G4f�j�H��qcas�����,��}��d�tD	ٷ�)�5�I]�%u�m�m��	hkQ��ҭڷp)�:J����mvж+n��\�������S��u��ϗV�2�L���D�h[�u�٭JR�=��ٗI�vU�TJR�]�� ����Ռ��U�V��-��6�1Վ��"�A�����z�!OU�>1J�s�2���@��/{i�r�R{J0l��oPJe��B�˽��a��u��y{88$�%�8Kԝ�ݺ�c�.�1���z7;c��3�r[�ԕ���빽q�Y��g��G#ű�aH��n��8�j�2�k�zfhG�y�|��y箴4S2E��E,j	5���#4���M�&!	���	BF�(24�6J4�d4h�L�h��2g9�����dP1bLDh,L&ȚH`�	a5�hBCX��2�9pb#��B��QE
S!�D��RH�3�(Y&I1Ȉ��`&F1�4�$L��@d$M�q�1"P�	(dD�%�HD&L��*�eD.r�����c(%0L�A$i)���"�i))��|��P�{�0!�Y<-���]XV+n�_Sd��ՙ��
>�������XZK+��8M���U�A�.K΅vt�л�I*Nnu'9�O���̝�~S���t�3B���zK=g��1�+�h>�Mg����,��}�1��y�Nb���]��W����.
q��S;�|+�\K�H`��[GȜ;~�A̸�# �\�M��w�[Xc};E�p@L:d9:�W��ы��!×ˣ�.�2EӹCY���{S�s��}��<o�V�&��n!�� p���u�����R��\���I�y8�ߟE���}��ļ���d�sqS��rI���I�4	�2bh�G������Z�cn��Q`k�A���h��`�e8����!uNK�H�Kً*�'��纼�rt�K�Q^�R_������n=�&���=�d�A��1���]cQ�����ӹ����)IN_�+Z�m�c�O�Ҟ�qAm�
�z��:��uZG�M� �|�t7��|��{<J�.�������I=a�����S�:/�s��=ѹw������,��Y��MP��E�1���\��Xkz3������:����S�vX~��[s��|��q��_�9���?S�LNQ.��d?V��������#�^���FP>QW]�]:C��A�^�:.� ߜ��1��8�����¨�oi5b�̋Y]�����zE��ms4�t��z>
����eYܧ��3�V�4�X��Td�M^�N���^��Ͼ{*��<W��](��&�+������_#̝�(�|��٩k�e�Ȭ�܎c0���#��d(u^�����н󮢳�%�����B��S���������nc��FF@�>��p� o'O�շ�3�	��k�tU�V�Ǿ��N�͵u�;��5y���z'�g�<2I�؊�怾��{�-]n��G�l�Z�[�����!���3�H�K�,��OQX]d�.���b�U!qU>Ni�{�~��5�~���W��zg�D@�ESrN����k̎�e�g�I=�r"`���o�A{-��"�[���w!VruمsIwQW�훋jϛj,���:I��d@N��t	�� 8�\&ܲl-�	5T:j��3����V�Oa�5����1��\�E�q��҉�1�"3.-�#ӽ�9�`s��|�H�+�y:�u�|sx[6ڸ49�Ȋ����II�R{e�b�Y��U��3����B�9����Cۅ���Ѯr��|�|�~�G+�C��LyqY��O��C�Z���K�Z؈��4l��]V��H�顬���CHF��ko�لں;Z�+�h4�0�9��;���c���ݓ3����|6��O�z�
�K�-�p-��X�d*m�)�6���A�Y�/�^��M��K{M�}����ҡ۾�N�+����vN�W3���_�2�ٓ(F*�����Nvʳ�7x��W��U$V�:(�r�c�i�䭿X�F����{���Ԙ�`6��FeKGs�������N}��e�]Ua���|���`�!�Yͦ�W;����xy�'ŌbЌt���#��n���5vk�/O�:�ю3�8ME���"{����U������2��C��r�+]ߔ{��j��n��^OMP�Dm��m޼�*o��{,�>�Ƣ/o�UT�o'Ϟ��c˯Fv��ٸ6n�/�
���h/��+:j���U��*��E�:k�<#���I�f#g����,�^�F�}9�<>�^w
73�n���c���_	�:�U�<���z�!��Y�<鳶��/5�b�r��W�ml/`��j��_vR��>'v���x�u3�n��U��Y]���_���_8=��~�]]��ʨ��6åѹ�/iϲ�*4��������S;��JXO"��a��n5�ꍺ�|q�l��H-�����[8�H{�~�=�!�ReK6�$�c�\*�te���i߸ˡG7�������=�����p5-,-��F�m�9��䇓���Wt�0���6��Eb���?*��
��'y�dIVW���j�j\;�騔�NKi�vU՞:�EɃ�n�X�s2��1�f_+�g�j�3w-3�&9h{][f��J͍����������Nϵ�>�y$=+<���z������9#�C��r�u�ǳ+�K�T�4�;�ծ�M	���z|���c���7F.��\Ss0Y�����$u���gtXqG�L�P�0/�{�P������u�l�o[gO��m����s(���7o ���*
�(�ԑ�	�/)�,��(�|F.���ݴ�Ž��z�rdN,���(sy����<�bm:
��)�_lɎ�9f��d��6X�jW!�zB���t�}Y�܎ɚNa���'�\E�GP�B�*�-~��2K��xOb�>G�v��u��d��f�דsM^�6�=�C�ܩ�16�"�>2���]Z׌�Ѐl>6vp?tnW_��滮�#T<^�,#�s��/��ۮ�O��hӺNsS�kQ隠1���OU�5��;�xn{�E���@/-�����7�
����N��s��p���e��;��_�g���S��H���u{�V}������᳡�ENQ�t����,	��d1��<���z�^��ܩ�,f�uD�,<��תW����ƫ�CyT̊��/����-1jw����;X2���K5� %�u�̭�ZވYY���5�l�F�^Fņt�h�.���n��+�gc��J[���X���T�;��lZ���p{X�ERq;�D��_n��	���y�/ɝ�!�'twȰ��kM�N@��`J�h��}�w�]g�[�ˬj��.��[SQ�-�r8[쥧�Q�;�dw�3�u|�T�Ӑ�К�b���$޵ʦ�yء�3�!���V��>�u[3ܽ[9�ҍ�N�t�$��gP��k�6=���Vw��,#bٗ��?[�g���C�S�_:�A���.ܠI]0�p�^��b�+��Y��D8\�PS=�)KZϾ���h_u;>��Y�>�1�+�hvx9^e�i�9�^�е9έ:<��8 ���ۘ����9��Z&�Ӵ4b}�h��Rt�OGGKw�{�۩���r�e�A^�]�0����	ѐ:`��yM`,uF/_�W���V�Y��'·����F�!��ǟ5�Ms�p�N�	��G�0#������X�{��T�i�f4o����j����9��G�mi/�ϡ�@sk")�~
��W�m%� ��z�\ϰ�Ħ��wt����m��]�Mm���K��{�!s�pk��R(l�{=����!ӟ�ö���f9���|��K�oa�z^���+�$����D��U���IBv!W;��I$���z����ה��+�0���ޛ�;V�=�1�N��c�Y���if)bZ@�{Jph�zT�����υڙ�� �J�#�#o;�|s�?�����zks�F���x�xouT�s��i��1�����P�6W7MTh~�3��wjm�qZ�6z_Ƨ�(��:S�n%ܸX.z����C��괎�%��r���E�ِ�J�����s���Ȼ�m��5�͒N���X����t]9�v�P�}�w��J��E��ʘ�p���{�7��tW��obg;�^8��`2�vG_����Aݖ ������|r_/F��|�R��X֞9zfd�Ǌ��y(��a��0�GZ�Vq��Ǘ>��T�_L7����v����G�����Z�{�q��|��Y�����u�U%ٗ��S��וo�^?U,�~�c��a��zh\��13ys-X�6w�'�/<5�-���I.)l�J����gm��&���=_)�����L�C���Y�|9�g|u��g;��z�,Gfnl�{���|i��$Fx	�ȱu*��R���WJ���_?8��0�E���F����Vy_���(��롹�/2�e���X:� x�v�P^�o4H��{�Y�C[�t�:� )h߶:#B���V�q<P��s�C+f�Bd�lC訝�Z�'�&�g2\�f�	����S٢2F^]���ެ�������vZY�+�˼�݉�Z�T.��t��p�_U�q��]�K��cu�l���+.'���׏�M�J����������N��v��1�����~mk�0#y#OǹD#���W����J�f�Q���1�,[̠�O}����ގkc	��ыi.���sÌD>�	�:6�k�7�:��Wz��S�:�T\Vh�m�[g�x�l9�pk����-S3_rJOG�;�0�~qX��Z^S;��&"��[
��7#��n:���49��Yd�%�r��>D�^k/��7�qM�����G��WQ�S&���ON2��s�U\��x��P�ک"���E�[���Z��"����TcB7\4,'�(�/��4t"���R�ތ�>�W�Ʈ��§׼"�y�c�,T�vwG��1{��ˈ9�������d���ݑؚ�5�=e�d��:��e��5+g7�}�=�^_�*�����f��C��fb��Ԣ��mA�=1w#�Vu�ݠ�*��[�s\�#�&�}gYUu���R]d����Y��Rp��3��r�#��̦yϬی��'e޾���F�f�|XG:hYb'���0q���>;s���W���O��P�������x���ST�m�����������펟�ѱ�5�Ǯ�9Ӱ�d�Q�Z�������,{Z�gE���WR5�����]��q�r��{�(�Z1�yݩ\}S�U�����&p�ؑ��e���������Jڼ������6�~��p��/��KG��7�N�g�5=Bk�dG�����݇2X��JS�
5�1z�������8J@�x�b�|��9���C����1�� ����j��f�J)�'����|�l<�<��P��I�
;�J�ή�S;��J\ogP�i�1�$��V�=w�jk��l���yC���8�)s,�2�.��t	>UY�s�T?jaz��W��{N���S7��V�Гܟ�k�}9�#��dǛI��q�%ېsLK'uEZ���B�@z��P:_�>/�_��ܷi��<w��b�W��N�qC�hË�e7��[���n`�c�8LFTsB�;�ƣW�:��c����}:��[�h̳���Փ�:2w��4L�đ����d\��n}�!%��	�l��щ�W�������gޙ�Jχ���AX�)�[2c���� �KFc��J#e�xfe�gf�Sϧ)fy�+�cک��2_�9q�!Q�UC_��Zd���R��Wg�칳���Ŏ۳QoJ�"��a�m�x�[t�|Yw���;�P�Dr�r��OMsU�M�k A�*��܍�ț}"�mW(W�1y��v��'�R���� ��U�k���{�y|h'Աt�|�-��n��ws�l��.J0��r�Y�0��z������w3��1�Cl��6�ǻ�R5��CT�8�/�Ң��e��^�3*�;�ej��W,��������/�.ns��iа�r���%�>�j!�A�'<:Q��G�j���|��0�
�:<qZy�x�qC=gC���.�S�M��g]e:e�������<I���8�fD�u��K��~�?��Ӭ֕�NNtL�
�·'$��S����X~�;�T�@�@oO����>zON��;ۢ4z���iݰ3�l�u����;�a�	�,\VMi�� y_�L
�vO�}K�1��N.�o�.SS�zW/xG���=n�����[o���G������^�?�����#�'���kSE�*l����s�������VǇgβи��Ad\�J5%��}�fDj�ji���VpS�Z8#���;�1���/s��������u��χNIw*��ϛ��yMV�k��	(��$��-oWJ�7ܟ���Y�6�q��}�7�>>1�S8p�$�r�|��l>����!J���\EL���n�M�v��O�m��m^}U�%��+L�Ň��n�i�0�t� %ʄ���*P�[��թ�{f�bnۺNZ���1��w[�����6��uu�|��Y��F�U��Lz��3�8��|-"�|9`���"�����N�R�Z9�)1�s���=ЛwԷU��"y�gb��2qZBs6oͫ��
��a�d�p@N���d
���)��X�^�P� �]���*�vVqY�����Ʋ-��	���4�:@OJ<kL�@H&
�u����Ŋ]�x�3ϸ�����.��F6�}]-�%���2k�mdE|�?�2�ޙ'��1�=�͚ ˎBk2w{��uG�q��~<�
�m�4i��q."-�r��Ω���/5!T��-'�4d����~6�t����q�hY�*�����5�:�F�mDc�rQjS�K�*��W�
���N<a��v9r��A����a�>~��9X��9�:���H�c	�Y���qq*�{�^`=�j�Q�ҟ�z�E���<f��I�L5ckC��i�qNt���=Q�w��b�S����ʴ�������r��5�Л/��/c�&�&쎠���t�;�+�xny�V�(m�|-��r��c��txN����.��{*��<W�ʆ3��t��yL;~Χ���nI���7���S>��K�`�MY�ԼF:�jv!�i����󮢲�	Cj"1���-�Έ���B�(��^��ڭD;"�=7��쫗��2\՚���,St J�đ�#q\�q[Ý��L^�z+���x�2�>��F�F��X��u`���hK��\Sd��[��8��
��IH�n��A2�7�R���z���Y�u�����F��GU=-�:Aq�D���t�Q��R�z�èV����zu��L{W����m����83ʧe�?�e��zj��ͫXr��)jdeP�=�&6�����15�f�<�����u��v��l�S*�ةuي�����Ov��{J���.�ʋ1*���":����s�r#5�w:uC�vNJ%;$�v1�D�r��'GK���|��$S.�]:�N�@F�ˎ�z�n��P��;��MÖ���.�u@��Km@�ݲ(��D��,�	hN&
�2�9��t� ��ow;��qGo]�䬩.MZR�{�V��{�I
-�j"4M���z��:�,w 9HԻ){ԛ<����곒�9w1���F�]q�r�v4�`�4֪��^���Isb�΀���a[f'[�6�8/�;���u�cQ����,CDk����[h�÷��{��vS������0��Z6|��:�LU��Z�6�1�ŕ��1�L��v_OQ~�y�maW��ڋ�di���e�øق�*���B�]�`{\8cx/H�n�q6w��zHJ��A\�
z�1���w���bs]�h��E4x�T)��cnz���PmZ�:�%�дV3x壡$��g{��ZB�J�u+q+� =Wpޠ�p}f���x#��g}�(�}YH��M���B
��1�)u<SjR���g fT�����k��ZZ�]�0�/
r�@0Wa�������!�1�â��gq���QR��1U���N�!��ǲ����F+/d���]oa�Ҹk���%�P�E�-�wWչ�{���P*�v�Y0NΘ���M儘�]�6v5��m�7]j�"h�{WX����ݳE��aK3P�c��R�#t�Ic�ƭU�bnG+Kn�L��0UΜ�/������*��1��>��)�7FN�xe\�C��v�Tm3%l�Q�ܰ)��-sc�%�Yy��3u��2�#p
��)��g%�6��+���H�V=���zY��\�s��!��6n�jow��ݺ{)�+k;��
őe�iv�8ӛ�Yz�e�d�m	�S�%�X�mo�;U��Qd�$ҫ&n�V��`�4]�S���֭I�ƌ��X���Ε��+�jl*��s�7�r�f��>����*�Ǯ��a�F$���9׹"�nV��S8�S�$�J��`���d��$+���OB�\��SCΊmnWx�I�Lc�ʖ����f�L�v{!�4qQM܊;�\^.�Et��1IJs�#�(������U|2�l}|h�3)���+D�%I��5�U��=@i��:SD��Q�W�E���Om�k���`� 1��̈2���"�3"E1A� ��F�2�b�0Ri��8��"��0��$��c6'9�FE��P4�B�eA �)B���\�C!E(��n30�2�9q��&IBH�@��H��SH�����2BP�!4f���H�d���HDDi�b!P�,�M	D̓��$I("HF$&"@�	������&d�ј$�D�Q���Ҁ	!@U
 ,G��\i�.ɩ�����|�Bޥak�&����u3�p<�X��ۀ�E7G�Р�m7��긯�Zݨ^�:���G�����^X��d��yD-�\�WN�g�����^�a�H���z^��;���(���yL��NGx)��+���B�S=ﰴ!u��y}�[;�)�Y��n�3�fLǬrH��ˎ^���+��L�RA@��b�U!2|���nh9�~��ꆬu`����>XI��!	j)��g+�}q���<c���e�I`� �H�>��)��tU=RiR3��aT��;����&�ڸ��O���l�}����:���}�o d`��D{�EN��=�ŭ�o+3T_ ��r��	�ƞ���t�!�m=9c���kͣ_:��T�E�1�e���%��s2Ľ.�,�����!��w.of�sj����dE	j��}���D��#�����5W��{���T�� ;�!R_���Ƈojh����,�����VdO�G����p��i�!�ګ&(j�h�&�ъ�ON2�����\��/����j�my���uɹ�ܺ�MmeYۦ|S(�����dw�Q��Ed���c>���e9vU}s�y����u��3~�T��������Ԥ��3V+����J��䚬�mܹ��i< ͦU_s��6�1ӵ���8`ΟV���y�R�hظ��1N�a5Y��G!��&�}cIN�_o)���dܒ�wQ��y2����`�;{�$U^�vO�v3'7v^EC�uS󶡩��r���c�"�������ݑ���,�#�*:�E0����yx���ަ4U�塉%�|�P�ӵP�O�ʌ����=�j	��C�u�ޜ'S�S�2%|)���"�5��_U�WG�ԗY>�N5�=I��<�\W��Z77��2d���.`~���`������zn2��VhF�t���&1y�{"\��z����p�W���fcg?oSƲyo����ܖ��a������
�}GEӑ�:��.�W/Z��Z��v����Q(*�л�I>y����^{]�1{��H�% X���L�d2��/���<��m�ž-Uנk��p��k��:[|��"���I�}GI:��yT��2����ê��}'?6ǣ�
�_]{���A�8�=�G��~�=�e �eK7�(��>3��_��a`*�ۋ�{9�L��
g#��w]	�=���0�mܘ�,y�1m����g���EnI�S6�Q볂��ZJ;���I�&��_��є_���n�8\��?H���Qڽ78l{F�W
���`�*�^��EϭN} ڛ5���k����f��
�ďx/�b�hF9�}2�$�Z�;�r�|0٥6���M7.������ɭbU�9�|[�;�ESɧ�:���u�Ꝓ���\��B6r�zs��9�]�2p����Q����]L���9�P����W�Gt��D?Z�7r�7�.n��|�z�μK��P7Cj��'�<kT��#=^ʊ]8͈q���*c�V����jv�����Y�[]��ǎ�e���x�b9���R�5�&;A�G��4h"��r�e�����1������w�C=��\�-�w"�7^'�=>}��`�����5�Izh�&��>廊�M�󮹌�8w�/M���7:�Ǉw*F��j!�ӈ��GJ�{�Xּf{��� �z���a�-��~y����ᓃ�N�M�Z}ǃ�ۗ�!/]���@4i�'<9Ҍ����8��8z5�Z�����5[�2�r�8Q��h�p�/'JzɳBβ��(w�����&�Ɋ^Z�ȳ>\-����M~����a���N����·u9GD�����`N_�!�>�ʱ��0�/�,��1:����3�cm�B߮�6M�#���zz)zU���[��d��N:�{c�Ww�~��E��O{�<�9��5�>��[o���Q�;�fza��$���G`c���vI�CZ%�މ8
�8},vj�Md���}�)��ن�"`q�z2�:��R��5�5}3V�#�%��Q�	)��YǼq�`����Wȱ��=��Øƾ䜑�r�g�y���ћ�hG�YH�./�ݭ���9
�!�Anլ_��[ o\i�,��
�k��Mz���Ǯ���7Hs�۠��Qg0l��P�B�5He����g��g��FsX�f��]����0�_����]^��-�x_�.g���9������s'|�%��<�*�u2�����9晝n��}�'��Ϸ���Z޼�|F�1�)3Xr��{�3�,�������J��ߪe?N}m։�N�Ѽ��M�v}�I�R����'�t/�����9C��;q�f�I��� t�d
���l�S�^��[4��=�Uշ�}��mtC�.����&����N�	�=(�� 5�$�^��[8q:�}2�ϔK=���r~�`D���8����<�%�37���DPj���I54�'�������2�0��gg���h#�mU��_nl!��v�F�m����q�t�#�NF<�kg�ɍ�YY�}.�HcfN��ɨ;�p�<ͣq�7x�x�u����Q�# �w��������>�õ�N��j<a��z}�q�#���i�/g°�*5^\<��b�����~�Չ�[�?���:��.!˔��A�p���bWV��p�:B4y<�ج�V>v��J�4=��� ������.��az�ؾ�2:Aѡ5Ѵ��$�%]��WzS^�3Q�ְ�Z"��&�%��m�v� ۙ������������Y͝ٸ��S9����{Y�>:�nmM���tA��z�]j,͛�J��\�O��ߩΓ�(y�^s.�eb�,fy�Cq�'���Ide�Q�|�S+^!6s��/s���C�n��^O�@�&�^�~�T��I�a���^ܭ�K���o'�|ʇ�61⸫~�Q~6M��U>8a�������ՙic��Xh"���qbjȵ^��φ���H,^�B�κ��
��*U�rϖ%�[^}��&����e���-4,C�d������y1N�g�����G�v�'.'�!f�<�-�v<+d��eƯ�g#���,.�ޚ���{ᅡ�Գ�����*Q��'w;�_U��þ����]b6�Wf� ��� �$�C~��'9nh9�����)���|<��ڥ�<8� �9_}A�/2�e��C��y g"$;����[8e{���3�&Eɵbk8yN'#u�g�&������g(5�l��N���h�_q��"�+ޛ�]̸bV
��X�un�q�i��F�Cm�B{������s�d��h�Ӫ��M�\��Dv����b���,�m>KY�@}j��Sc�Wg*ޤ�#�x,���NY�+��n��=ԎIJ%Uހv8^���7�-/�Pֻ(����R����x��5��z=U���{��oiX]��.��GcS��u�}��r�;E3㏩5�i��O)L�����u�7'��#\��>��>�-��P�u�|��ه������9��{����-͏�|�a��$��P�%�� t�~�*�_���ơ�ɫ����a�>���>䳗������'��1@r�h�&;s����eE�l�=e}x��[�s]wM�H�W������H�7��r�c"�9�b4k�h�D=Ϣs�!=�W��[tp����d��s�����B��XC�4��[�P�Mǜ����f�1hB�FN��R;+蛲95�sP���a�����>8:��=�3ض.*�.��I�s�;Ud����^���w���_�X)�`5oկ4o���+�+$syv���l�y�W}lgʪ���ׂ��*�
Y��ѻ4��P.2g�|���kUYi1�pl�	��E��P^J�F�t�#������f#ܚ�;jޚ���z�};�XǱ�f�?+ƴ_�9)/t�Қ�����Z�K��B=U쎸�b�#z�{)���^|��([쥧�ݣ=@�$�#�S��j��e����,���׬z�T(L9�����/]�[Ր]:C����T
n�|qE����{�m��5��^𲞿4�ʊ�"U�^&ڻv9`��(��'�n
wi�Z�^��A��F�5�u�����@��M�����9���e��p}���˙�+&$�{sRU�j�!���Zp�����Y�#����"�$�3D,zs�0h6�Hu��[QZ��-)�y��P㽅��x[���1ף�t<>��8eL�̢K��Er&�f����[����q��=�Iq���'�?�N{���5���b���?LP�)�U��Nr�c���b"�X��Ѕ�9�5�2�㖽�[��f�{O��F��F�KY1�Z��Um������+Jy�A�C��]DL����P?J��5�.�#���/���.��{JR1v���.W_svM}���UL��<��CT��#<
��x��0�f�
q��_m_�n�LS��V�G�oh��3�OxCB�/�:tr�ѡ�&;hD�����\A�Nc��L���K��׳��������0�7��b����~��~:����P�t�64�/K����θ�Ʋ�2�oԘs�Yg���A�Cq�8�w*G��CZ�8�/�Ң�=�P���j�	��MnХj��9�vfxB��`�GRj��;.�a�*�^����O�cQwI��v�P|İJ��j��w':%$LKǶV;�2�/������FM� r��s�r�������4�Q\��t�췗yɗ�'<Β�&w,�B�s��z�Z�� &�'�_��r�,������.g#�«�!�G]$!2�,JYE)�q���f^��{���;~�Y��$����Q�C���ۊ���+Ưo�J���
��\	
|0+�W�崕��G������V��~��9�~�������᳡�T���sce��'y���z���U�h�ܙ�N��#Ó����3�x�l��륇�l�� ����_�Ҭ�~p����G����GGQq�5q����0w�Ѝ�9�sQvp7�b���ZTQҨeyg�&}���H�=�Џ���b���a��b�LÍ�,�_m���X~N4�^��lP��J7Z��i���Uý�ڧ��.O�Q���F{M#�7�}|�Gz1���na��[��g�\�fDW����{N�L�������NIW�	(�<�T�sS�L�[�fn5�����O��Yۨ���޳���HX�
7�����f�|��86���<"��|�E3��wO�^F��8W���!�n��dۨ��[���l���tUq�v��� 'F@��.J��Q�����Wb<����s�M�{�zu�cy�������&��t:t$��Ƙ��	�}�U1�ص�@���s���B��pm����=?,��.���	�t��]6�I��k_���Ԫ�*�_c�ߥ6"�L,//�RY�F�h��v�z�����v��w�aӒ���w$�W��?l��\��mu�I�١���z������e�����H�r��m���ǥ`���:�$���?��nG�a*[�C���<���37��ȊS�T9$���oG5��1U�6��<w��,d��ȸ���9�3����h�m����q��G+�����w<���V�Wb��_%�R4��8MBخ�g�ز��{*�\=��h�ħ��,l:���^�S�)�n�3{�<a|�z��R�j2}�훊�8Us�U�z�8�o��U��x�2�y�\��hǹ��Q�@7�ҋ�1�(��$��=#�\�v.��':N���S�*:r�$eNd�2�_{Ey��FǾ�]��F9�y)�������f#��d=Q>�8S�1scwq�s��K^��t-8�^�N0j]W���=�vo+�u��:l����"�j��f��D�bh��C�༕�G;B�D	�Ց*�/��Ú�~�Ag��h{��P�<^s+Ѳ.�?��g�N�����U����T08aH�y�Ԏ����,�~�5蕢���=����B�[���E����aW�g���򘿩�f�׊��f[�{j-��ի�6�3���K .�_MAg,׭��׋P���9��=���Vko�I�n�	�z�J]������euG�}{|��6�V�륲1j��Ν6,R����W]��w�3:� X��AbT�TrIO7���<�.�8�ۘ��v�*h$���*+u�R�Ѥ}�[:ԇ�:��J�L�֤������,IR��U>Nf���̐�E��X<�w�0�����G���o�K:��ǻ���J7�<I@��46;G�W.��޳��fE^ƿQ`T·����$\K~���{=�Y���p������h���xA��72(?tm��C7�c= *����F����mb��'�/�h^��hŴ�B��v�RZ����m�i֩u�Ó�  5��\�-;m�]λ������.���s���^�pV�k���㯽���^�S3%�T��n	���7R��n|�\jj�:dv���8���t<��m͓Ź�i;�\�2+�&��c�>�U	��TW�猯N���ZG�OwY/rwW����)��j��:1M�o�G!��a�k�h֐�����uq����w�Mĩ�c�R���yLd�����N�b�[P��r�2��Vh}�Z�����#����_W!&��O���:��ҿ�g�1t\!W^�Y�<7�a��j���s�6w�M���J�o�~ux��*�yr��^7����.���L��鄀@��F�t�!s��|�S�i",�z*	���Ӯ8���n����2P�J˖���hkj��ms�ljY8=��".l�Ӽ��
�5vM2�-�f��΃w�P���	=�V9�Vc[r����s�dԶ�QP�.h�.��� �����I�V�7i`�;��2��9���U�r���]�^%u%��Zl�T4ñy��5�ݐf1��e%�qL�c��b
�^�@c;���O�il�B��U���J�R��_r=���y�����󛮢�RwC���NuI�����q3��՛������"�P����A�Z2ҽ�8�tzP#��p��TX��Á��a�/��,S�p�o�د�2�]�(��k�i]8h���|MT�h��M�]�2��\�NѾC���e�Hfb�<皺�+PB5���[k)�j��I���Iv�,�6�8M77k8�����K+*Jf*��g��Httj�Rk�X���x�V��j�upL�B�X�����d�
����J�ܨnB��t6���2՗Yj}�*s'e;b��Eۘl�&[���gW^u��Ct��-�YL:O�(QAQv�txh��/��X�t�H���*�q�H�k$��g���ԛ��g���R���}c�lm�|r�o ���*���:�8����}��qn�ݬ��N���&�
���k�)�b�^˝���.�enf-c�
9H��G����>F�}���-���{S�WC7��M+�SM�B�3r�<����Gl�J�����5�iv-;��N�e��9�,��8���z�X�۶�j��ۤ-� K����yN��9#�yf���r�(s+`��<��pٓv��շ	��G^�wv�ڭư���2#�F�!{�kV9X�*��.r�*�I���Yջ�m�s���.))�t��o�qL��K	kT!��c�}���q�!�����3+k���9:��n��#3��i+F���z���Z�2B�T�
q��Xn���# ŋ!�-��d�J�]ՙ�	:�r�Es]D�ʎ�sU�Gݱc�+�۶�<�n����9kV	cC�,���t�>ʕ0� t^ݷ0H$�˯yP���qY���Ћ�	�}iÚ:u:*\��\��}[I7�:�ݠN躲�5I�"�̃�w˲:Mj��w��)K.!+�*�T�:�wR�	�3��� :�':U�/�;�2�.K�{y������n�f����Y4��eЉ��g;moG[���`@�!���lfs����XZ-�i���U�j	C�X���FmmJ�����b���s�M̡�õG.N�ƱU�R�r;[�FGN��;#�,tWej�IRW\9[$�>;���8®=J�s�����luNa�����P��w�"���b�Y��s$MQ�����Cg�L����
n��ʶ;Ǯw�A�I$cI�4���D�BC)��P�	�D0�EX���Id$�E�0)��1��1b��(��H�$!h���d&�H�b�#�8i�1R�%&JB4�i4��SI��M��&DRS6dQA�,���6#BHC4����lfQ�c	E�AQIc`�i0a!(���
�ƌd�%�#F��� �b ��h���63�#qF�Cch��~�u����_�kﯾ�{�\�e�̵o�q�&i�����|��^�u�̀wGԀ�05��&��"�� oZ0����\������w��A��Ƶo^���!߆�f�	ԝ��q���8[����P��g{7����y=�����c�C8���!2bǏ��P�	�[�#��jZlO�έA���G���Fe_W�з>�9�|sfb�����}GEӑ�7����ҌH9���읽JX��V�#�Λ;i���u��ۥ��Q�9�gc�A�!|%�ӎ]99L�i�A����E�B#�t�|��{�:[}�<��P��J(#��@��73D���*�*6[�D�JS�6�gz���}G�����Q�޼���;�z�H>>u�����}�מ.�U����\�O�ZA|d��
�?{v�:�>����4��yv=�n e�K}5{ʳ���l���� '5'��
`LJF���Z��M�-�	��Zg͜�c���]cK����_������uL���g�F��3��B�3�4 ��k#���:8(��z�����ˊ��!�v�ls>�89���S*(	��ھ����Tyt�7I�_?3)tbӈ�Sz�r�y|���6�����4��Ք����y�X:�T�d!lzz�1zk[<��<h˗��f�R��5���3��|�E/����;�8�q㵎��_A���j��t�3t�C�dC��A%�5�����^e����͕W��W�'�u1����G�{E�|ϙ5�4,B�N���SF�ٓ��ֈ=��]tA�#�������Ŵ��˕g���0/-��ݖO8r�-�GP�B� 5��*o��cDu�ER�p�[;.��,��B^����|�#�lf;��wr�zˆ��~�� 9��(�v�s<��D��6�)�c�zNW�Tv�P�&��#�\Tixj#��Ľv��H�S[���}�o�ӘV��!�{�u#<����P}#z}I�_)�&�:ʫ�8���Y�+H�nG�U˿ga�o8��|_�p��?�BC�4�g�~�&���<}&�J�⯬׫�nt�#�3R�R���P�s��E�����L���l��߮�\C8Ne��yB}�)	׹�0�*^ޑ}ًW��3}��ao�.%y{t�g46������e-*(�K�=b����+�:����|`�j��A9���pY�����ʷ����u[����4�p�qz�|�~{�����?�g谓�	/J�̎BL�5�:#4��N;э2^_?\?)]^���L�u��	����ϝ��R��={L��@fʴ.s�Z��KE�U΃�E�*�6�g����:	�=��M���uui�ɣ�	/�<�)E-Ay��rsz�d=Y]/�%���v]���M!|�lɕ`���ڼ�����u�wnR]\���a�VEnO��t�uL�@{#�ΐ�]r9ji�^�iu�)����߽��:�*8�P�9�n���+̿}�}�1�ȁ�`Ђ��W�gY���x���*�����}�]l\{^:�7��6r���~�fG���:��[ ��������g�iu��Fr�y5�C�{������ǭ�FXmf@y�|� S�G����:�t�~w�2n�+�S�(x���V�,�[�C��!��/���&���DPj����;.�U���B�jO��+�N�:7��o�̭��:���E�;�e����M�ڼ��S��-���{޻�o��Ԋ�fNʅ�Ф�>FŞ���C�!5w&�y���پ�Ҟ���zp�,k����EO���ρ�q�>�'<}�֜*笗��^�/Q}^#3��ئ;�T
l.F�� ��E�5B{$�_E�쨵q��7�+��,�&�.�w�M��KQ�w���~��|�S+<9�Xhs����s��{W��v���z��99_�c/:�;��8#[�'DyI��� Zgm�5}�4�
I����B�)��� ��19�h�AT��3ʶ���*�����x�Š�]�A����[nғ��V�sU٢�knB����ճ0�3��=�T7��y��'�p�9S"�,ᮔ��&;x��ѾN��k�0��������^x�3R�9	ח�<����ls�m��'A��I�,z����d����G�b�KƀGY9s�`{^С�ֳ����kcv���uf`f�l��7Ap�w[��N��S���Izˢ��/�G�?i�g�5�`1�ֳ/v��N��k=׹>�Y�L6��u�m��󭢅 ��|&x;��{"�]1��L�C4TC��̼����=�I�v򥖏2�����U���\e��$Fc� "��R�b��ˊ^��Ţ���8�=s�����`Ϸ��E�<G�P��x����)�CNu9>�~��
Z�p�ݬ�jwM|���D���z1z|�{�����p����y�3^1��]܊YS��1���dP�7�! rw�GYC<�Sݾ��O�ӗ�4/My�b�ӛ�+�o��e���<��`��%O��3�#L�J�T��עGa�����eϰ�$l�r���������-ݼ�����U~3n���B�-M� t�O	��Z|7~5��=�|v;�3}PvpvH�>�oz�@��_Vu��=�"�b{�ui�ʍ�]H��8[��RX�f�]��:��|�|��ď���sk�.f�U�]zө귀�P@ItA�l�=�}; U�����hL�w�ymc�ʆyU�7	�k����`}2X{l��TJp�o*�uE5��N�ϸ�}|�28Դt��#A㌨����)��6��	Ǟ7Y�s6��E��1�7��C{�l�{��9�b5ԴwHz�NQ� �>����Ǟo��C��X�{{f2{Uz{5�Lu�������Vq�H��FN���ֳ^�>N�eu���ϘX�O�4�����w��.]z�f4����fk�j���fb������CeV��4���NEy��} �H�ݨ��ex�9�⾫���|'Rv{��fo(d�W%Tb���q�>�M=��=�����/�������GY0�xD�X�7��URc���3nn'­�)ˋ}f!�\�O2.�ʙ�ϭNG�ܛ6HA���-�	��X#,�O��E�����������"4��	���j�`�ۥ����fP�x�7�g��������+s4��W{Z�>1�n.Tv��"0�t�}�ms=��l=���"���J(#���E��G9��*�Cř�AL��"�]����C�%�<C���C���-��pލ�7�o�)g(�&Ϋ<�0H�/�4e�YX\kx�C���ϔ���N|�K}�����g�3���T����`5���#BĮ�WA��
��7��X�l��xh�8L��f��2�6�K9@_!f�<�o5e�E�7r�s;ȥ�b�m��><���b��\��<I����=�>�)����}n`N%~�ϗ�y�g��|zE����sq�!!8\/G�����>�r Nk�< i�6�:ϫ]Гܶ9{xx�>ix�����P�Tsŷ1g(7F.�t����|y������@��{Ǆ���J��4M���z�)�{�<�k+x�|]�ts>�<���꩕�G�1�&#$�r�T��8���Lu�ޔ�b��x��)�Lv�'{E�9�2y���i�����}�&;`i�=]>�Ǻ�Z��O�Q�w.U\�hnm7Lot�_C�o��=��su��ڿ�;�Uϖ_lm'Ȱ̓�h� ��+��+C��?.����#]r�ӈ��Wn������*�����N��͏P���'k�*;Y��M]�G���,�����n��3y�w2�ʬ����y����q���؜��F2~�m)����U���)��F����J�6��a�5�{yB>��y��#����p��?�%��e3�t�s�3�*�:��@���t׼���Pwf� �|��ӫ�R���@���R�]��G��f]�}�2��.��@r���47%u��7��sƇ5}��N��1=Ψ��S�5�ݳ:f�X/+�;ṓ�\�lEZ�V���R��Rw)�ǃt����pFg �wÅ^��QJ��7�N�?e��C%W��~�g��gv���-��Eq�>�|���J�y��^ۦ��0�+�C��D��l�ׯ�=�6wͯFa���ث}����~�YS�������q'��(�!t�,4LGmć�yD-�\ܫ�ǞG�Ѝ�%@�������b��,��kC��J5$�Ϥ�+�8�PF^�G�o���D!�� ?0ִ�ᙹ�q!b�u�s�T�p�ϕm�r�%TL�D�z�I;�/��>Ҹ̊���;����N����eٶc���:��Y���87�RAtg�����OW[�7�pjs8���lr�^���}}բT�q���v�d��=@�9�2�E�p@LGdQ��v����9��nLC���#c+Z���]���-��%��:����E�iz�'+��^l���rG| vA�����}��0�f�?�>��|��2�Ȳk�mdE���EK�.٫9����^v��32���>F�d�Z�#�n��H�W�yu}��ѯ�k`�r
�������?�a�&َ�V�ژ�n�$�.���6�r��~�~���q|q�z���xgdu9Y+$��ԡ�y�t�!nK�YWG4JQq3�Z�����P���f��lp��>̦��+A]H� �ll�’���F�f�뵕)Z��p�W�z�
�mS��4ԋٓ�4MA�
�R��5g��x�|3�ML�ȟxWq���&�I{��(��"ވ�q��>^�;>�ƌ5Ӷn=����#*
ޞ�'$���H��W�w���"�[���9@k�X�Y�zI;b.GeE��P�7��ݠ�+S�=����3��U��ݗ�6��s.�e^s��ֻ�^>�	��+�]��r���=R��Va����΃��ǅ}{}lb�w��u����eCY>�\wz��\PP�zc<�ne[ZU�j1��7tdg��hu|����d��� ��^����U��L�7��Ys�z�3ٟ��{[�}U��w����V��s��ۉ���3�
��Zn���t8�+_�*��*Bs�js��7�zT{�dW�qݏ݌\F���C>�����X�'��^�����nE�����;���Uv�:��#��e��峾�����[=�|TZ�
���*Qc^l���y=���u_m��W-���So'ղ��CN*6�t����,����6�5����Q%�P����ٴ���~X]��}�6��^�+%�����9��6�yњ���Z\�{�L|�ѽ��2���1�)֗8-f�D�Y���1��2r1�}�u&;N��-]�sZ�=�k8�}No^KJ剥���o�|���)�G��3�����s��[����<."�_���n�H�oף>^�|s�<G�W��6k�t�9�6��D��s9��
�,�ȁ����b(��4�GY���B{����zr��/M��s������^��J��do�wlW)�� '$7��C����0����_����T��ʗ��q5lǲ�7*���|_�ڸ47��r�����CT�ٯ��ɍkaP
{�����.��14�y�鬿V-���?�eo/Ig�9�q=�\B�2��e����*4ON2�_k�b�bVE�{���˚�T��0�p��S�v�"(os��2�y�C�sQF!k�h�̇��*�����w^2)�V^T����9V�';eYq���xouT��������h+5�Z�0��܆�������2y�Hˡ~#�5vh"��غ.*�.��j��_5�;Ud�_��q�,>����Qo�Ǫb�uA*�F��C���i���8����c N���nA��-�J��Խ)�W���[�u��v��.��� ��u/%��:ɳq�3�;.n<���QF��^b���h��[�e`Ї��āt��6E� �jC��,��OenN�rSكT�$�g��㱙G�Rlj�-T�m�`[xw%��S���(u���8�.�μ;�9�sR���aVǴ����]���mV�ܦ�:�g,��^g��S���F���NmO��͙c(zPrrN��Y�����X����:�Ç�љ/�n#��@���Dp�t��	���w�����H�Y�R��p�V�x$��S����pץa�0��\�{��"6�]8]�5���-������)i���ʕK��Boۜ��q&�c0�A�R�{M��B��tw����lK�~x�=it<2��T���Ó���72m��<�b��:I��$�C��Bz\o
�^ݦϾ�N/:�M�V�w�g]�oO��:���:���q�%ېsQ'��	T���qFQ~9m���@95v��gK7���,=�g���1g+=�#o�V��8�|��]}2Cs���B��6���*x�q�u�\�a[������!�Y�n�`y��:�eA�ʀ�$��7<����QRP)���+�*hN�<��]r�~�Ϗ����9�2hst0C��W�S� #��Ċ���z����o�bS�s�/�kL=�޲�N���q/��*���}G��}���ֵ����mk[o�m�k[nm�k[o��kZ���ֵ����ֵ��m��km�궵����kZ����kZ���vֵ��ݵ�km͵�km��[kk_��V�U��kZ����ֵ���m�k[o��Zֶ���m�ʭ�km�Vֵ����
�2��0�x�b�������>�������|z$�J�H�J��BJP*H�B�RR�)owAR$V�*B���
ADR�ERJ�����)DT
��!U@PT��)*��*A�*#ͪD����CL6�L�`��Ƥ��l�cT[e�;��F�\ ���%�P�l  s   ]�  ;71NBCMR�TP��TF�lRWfJ%JUR�Bf�Tkj�Xա3YCJ2UJ����'J&��Bݸڹ ֻh+���6a�����A��@5$H�Znr�+��F �	.V
ћtZ��#@P�A�l�*M X)�5@@P.�@.[L��v ik
�nE��P�"�⨊�;���BY��$T�T����4�P�QCX���2��֠�n�A*�-6[m6����Z�D!��Vش(٢HU	Hn 6.F��kL��f�	��6i A,ƥ�i5��JM�0N�!�QJ���	B�3(*iI6�j��Q $   D��*RJ��� `�  )�IJ��& LL0&�4�ɓF�� �0F`��T�� 1 @142 $A �I�S�2#5�&������)�4f��2d�ɠ 0#r��n\0�W.Y_��,�1��ʱ��7Ȑg�#�aw�'S� ��H�$�~t��Լ$��V1~�*~3�~��L?z5�UJ��F0�IQe$i���&���T%UI&T��N\m�F?NV����Ј�8��%�K�u��f��;�>�%�ڣi���Z�]�rT/?��/�J���2ꙹ����Uh@�Vc�[[��Q�1Ϡ��im]9���#"!��ۥ��1-����9��L�k�zn�
���t@��w

`6��J�X�.�:ů�7ot�91�A������6�`���6Y܈���YRkܺ�6��>� �=��$i��T�/��v[ro�u�8���ҫ�a��m�#:��e0[�Z��&�U�Ud��=����
�m�Y5�z����[n�t����O)�u��ل*�1��4�Jf��(n��]!cr�n�*E,��� �*b�"���U��O@
*�9���W�F�P�7fG�sv��Qc�[�k�u�SuJh�
�U�5(`Ӡ�[�/���W��k��n�RU:.nCVI0�x��Z��Wb� ua���6�i
��T�����]`�J�j)٢�J�!P@R7�Y:"�W�{YW�Zj|���STTz+m�cnѼ��R�S̻I����P<n�U^�
0�9�Z��s6����k,��߫H�77]���1u�5ܠK0anKY2��@�j�oiQ5X�è�hKKn��5P��Q���M%y�t�
Kں���7w)"��QE�QV@jk�6���5�^��F:�(PB%�e�0�9���a�y35/4渂Z���JO^�Ӗ�������8�U��ޱWh\�۠�c��#X��B5�`e����>�����h��Dԣ�E�A��v~Xa�R|�R�M�ŌI�N�2a��y��:s��7fdih������@���S�B�Z�[�CR��+P�2���	��:Y�o�"R�H�J�`�ňirf�BA���2c�g��l���+}�����}q��c
�E�J�xHZ�4wN��]Z-@�v��P��,c'qҊO(nHZ�)�r�������c��̻�1��!�ޣ���{��f0�Ԍ������d�X��wMU$�d�^C�a���z�1ԌM�łh� ���XaFK�a9ta�HIQ��v>6�5�YqӋ�[��{��I�9��6���e�{D�����V��*$,捼��^-��T�|]R�k�X��CS�va�X���TA1V��o-�Zðƚ:�H�$B�$Ռ��w��%�����
z�YW���W�rZ�w$5��RK�Z[g	6A�dJ7����Me0�-����D�)gc"Ĕ�9kf@��7_hQ�W��ɶ#��匦�@)���a8�*H��5�`���AnA��76B^Ғ�R���T6��ȧ�b%�C��ո�����ȩ�H�s]����
�v0�;�Ԁ����E@��N�t.��oR�w%UҤ��bN
�ێ�Yi�[�&=q - ��͵l�����+2m)R��ܩ�e7f�(�����K#�>��5pŤ̥[�[�A'P�kf�5����#N[��`�f����nj��Y�ȳ�;��7`�^A�zݝWM�j(������75yf	�F�e��IDT�V�ı���M��i�K7�fM����mυ��&ޱ�A�7eՠ��kYb��H*��vh�,ח$��!V �h�IaI��ͣa��&�vb�W`^�0�ک2't��FLvkvȥ9z�Gt���+	·5IF��I�Wm�rjX�4�p��"�0���e�%� V�mL��oLW�e-�mn�1�ܦĒ�X�h�b.�QM�=)�t�`�/���[A�x��0Ê���R��%(�Y�Qͬ����G���u�Mx��+D� �e�Z�[U�ಶB3/�n�=�l«he�w2F-�<�t��Pn!�kY�_[/��-�E���h����J��\N��cfish^k�*�(Vm���

##4ȌQ�ub�E���R9���W�:���V�
Ih���&D��MƩ����	���j����J�����7V{W�q���i"��|)⬭���V��S��q�qaү-̛w�\���.���m嵓-f-v7P���s3jJ�b�13 7i��3�ĕtͰ����gr�6��V<��T�ܣ�ha;�V��s#%-��)���Jۙa��ai��#�K[aB-g�dg׻�`.@2�/��̢(n͂V�]����
�9z6�kf��8�J���n�ţF�۟r+ЛE�l�m���&=�����[��F�:{#pĂ����yr�Ͱ�$�r�í*!�+Cb3ۦ
��dٗ�����j��N۳c���%�K
}��#�L��j9(%�G��}�;4Z��VȚ]S�J�˱i�Bi�wH,TԀ&�2�
���C�!p��+Hkh0�7�������U73KlW����$A��em�і�7t�N�<2���p蔫6���[�q�F�;[�NmȈ�J��r�&��R��-Y�fSY2�GK���e�^}�Fm�[��tP�T5p��ND)� �I ZXݬ�ah94�L�;@*�M�OQB�n2o7�	�Q�#%�]nI��*�&�#*0�Y���B#LeD���d�nåj���J�A5�>L�:v���.۳H�
�^\�V~�[y7~N;���S~34B���Z��9�����shf챫5`כ�&��s֩�y�7
�0'�v��;(�� //.!��Kl��F[(R���ݿ�BTB���&a�dR\�{�c�T�f��f��n�\s���h	��Ґ�5]!��^r�;��)�@�x�*�ܤ[�N+{2��6[�;��if�����S�VZ�W�D�0t�	8�RY���/�~�����@ḐBb.�,�r�M%�Z��
�1�tڟ!JX!R���j����^U�Õ�m��PE�\���J�E^�B�f�(�/%$�(�ܼ���!+�L��HM؂��@F[���DF��7F5�x4�&i[@Pi..^���B�kZ�����4K�ia��{��ysjk�e���K�*��d74��;u[��iἽ��Ec� x�Y�xo0�&��o`��Y�`֞
�(�jQ�+/6�7�f�+��]��Ӣ�o7h��JX��m�'"w��]� MR�x)��t�c�vj������hf�wM���zE�׊�Mv���z��6Qn�mձ��E� ��~��G������Q�?��\�pH˟�������@M�C�����#G[�����Rf��%"�GuM��n]�~=L��!D��r��V�����n[�`us���̏��ݵ�J\iZJ0d��:���������}���[{w̠�T��8�5���%-��Mr�u�i�3��r�Q���e��zL�z�m��.�
�B�%WmfTp�+�̾X��!��� s�M�7�Q��T�';J�Y�����}QTP�Ţ{{I�ӝ����d?��J�f[���9Vnm�mr�[�T�J턬k�9%���7a[���B*�p6���8,ٗ*�f�r��^����=��#�o��v���J���508	6���}�}q�7h�T��L��(SL":��w�+�X���uv�7�c���'<$Y��w�L�t�PAb�u���,܈��G'&:`2m�c��Yٛ��n�׺�c]؎�L-��ww�2vVS�Ϗ\�ȸ-1]W�*e�'�1k3\w� rO$��9�KA\���v�v�Vo8�����'��B�z��À��h�0¹�<h���+8զ�oM�F,#��U��/*�o�oej�"U��1^j�����Ժ���Wr�|nV-�J������c2������+�k/��U�Y��K�B�۝w2��O�ٰ�]��ufr
��8�b��Z���*��$�uC,Y��M���G{]���ިH
;Z]X�鑜�׼�Z�V&���b4�jp�ڭ�r_m�*�����|;3ot���y6�4�/�Qk��xn-X��},Y�'Q���M��ٶ��#���1��G�1�����,�v�ȴ\�i��h��v�Rc���]��Fe1H�rR5��`�L�)˦�桀�u1��I��y�B�a�EY��5\��h����7-Ҿ����6��F�d$�pJӹZ]@;�>�H�-&��q��C3�Y�YEq���E+&\������j!c��X��Ǵ#����-�Iւ��鬀�9�C�\�b�������(�����쳉��w��>v��Ov,r��@C���ôq���m*%
/���+�����\��O�d)ȍ#N�����&:4���8˖����*����i#����r���imf[:3�
�T87�<vV�)�u��x��s.�vD��d��,�s�;�m��;�y�z�3�񠸮������坍n�n��N��ԥ�Xg���-�B��}Sr��T�_pR�t�	�՞�wR�mG���g銑���]A%��1�����eF�,��n���'3�����^h0B(n��"��I>y�t<�Mwi�g0c��t�͇5�\���3rL�8Dx�r�7U�̩5VG�7Y��zM�48���]�9�OiqQ�Iv���йw��am3W�5iz�@��ШY7��]
����-�;�P�/A����\z���z����hv��EN�l镇B�>���u&��;ttN�Ѹ�úk[�BƲ/��Q5ڳ	Ț&�'P�XZ0��*�B��N!�m�w�/DJ�S�؟]V<�w�X�����NhWqw͝��˒_@:w�t�ynH�`s#T�F��ܧ���v��J���͠�w-����ălE���cݟBx�f�=��浄��wV����d�.�J�Kt���3�?�ӻ�b�c6�gbvUU|U�aJ�y��T!uE!��ei[������su�[6�����6]�h��iKD�2������x���{;UV�Y�����nt�[[��d�A{�2�"�1Õz+��ԴY.dR�v;�mB�VU4GF(�g>Vb��|+���(rڳ9��\V�N��C����xwA�1R��6��r4�%ά�NP�틷O�Ho.��؋w+׍W*�vѶv�+�K��w�7[kz@�v��Ld�P5i:�-b��6���:t��wP��ke��#)p�=U��IU���u���;K��O��U����{h�;����n�\눙-�*k�V�Ɇ!F��l��ɕ�PEc�f�w�LR��P�>�oX-]��X�dĮ���s�{�;$�1�.�m�dq�uV2���+��;��tYE�	7N�;2A['��,qn�f<@�����kH�j��n�eK{��c��[V����V��{�:�-.�q����+iӻ�Ӆ7�qf�
�,X�yN���睲a=38N%��w�r�O���(�Rl���\��4w �ɖo嫻kp�u�]����+Wr��ۆ��P�Q����[1���nnl�����P�P��t�-���ȣ[�������9�Wۮ��<9�:�Y���P�֪�R�	`�-��uV�pX�Q�����K��� ��y(�f�vwe�Z�����9W`&����U��F*,���ң�x�Wk�u��י�;���%Խ��EUDo"��Z��4Ȱ��Z�� ���$���2�7N+��T���=���J�[�A}��<���{��gk��/�kwO#U�Gݗ�i_l[������s�w�KRc��U��{�D���jƛ�W�Y[���uN;n��=�3>��ڏ.��'&ID�JzM�k��)"��X�U�TQ�H�giޝ����&�5���Q�]R<��ȇ'1s�F��6����P�W�'R��@��񘰣QN����nS"�ɉ�����K��șư
�,u��]Z�U��)I1��r�K���^gN�����̅kC����T�}�d&�y@�w@��� 0��>�(�F���w��TMu-y=�xҩWԁ���L�!R��yFIQ�/9�����f����+��n����膁<���͝�tc���
����β�2���y-p��ֱ�iu\�;�l�ɬ�&2��;�h��_k/(c*��K�o9R)�;vL�X�17�/�3b����Y�2�����/�ǯ�1�)n�dnq���$6u����O3�"�˶�T�(_hӗ�j���ӈn	�"ro�,C@�N +���I@�On�h�$�e�fĖ�N�+X\��AI$�I$�I$�\�q��l�E-�'�vJ�]�gb��h���6�ijZ�2�v��E���j�
]��Q�ôBK2���M��I$))hJ�4PA#��'�e,���rI$A%.�����q*�6'KN�m�C��i.Y��%
������$�I$�I$�I$�I$�I$�I$�$�I.I$�I$�I$�I$�I$�I)K������S^���}�Ym�mK{�G�D	$�dS,���vZ��'j6i�UV��F''����l�}xv^�o5���/�Uf�������j�%՘q��8�]�P{v�f7X5���shh/(�4~[�(��%p�M9X�*5�,G��X+���'3����u��Uj 1aq����ݻmt㷽m�0�@�A��۬ދ����̅�v�r�:��#��;)$�ZO�,υ��a�[��-<ll�8e=[ӳ�.m�n��YJ��k�2�v�/��6�|Pr��*芻3�7	��p�t�8p��Ӹj�n�D�|z:���Y=�����9�omRK��#1����e��Kp2�SZ狠�����X��,**��թy4�g�����:��9��I�+]EZ��ug�VcS�`;�:㬑C����-��2K��&=����'��[�BG\��QR.o�;խ�0־D�b��\��v������	���Z�(��^�mE�e_@ٓ%w�wV\�sd��L{�X:;rP��HNk�̺�b
���8g����w2N�}����"���<��F\=�0R�Fw��NI�g;	Ε�����_l=/�dxͳ�'��Қ&���ئ'[������8�w!�ǝ�� p.���}�����X�u]���:Y�wOZՋq}o���%c\G	Wî){�uqf�y���l��������x�+6D.I���jה�֙a���Y��G��n�Nu��0�e��ٛ:��FZW*��xx��(+4� ����5�P�=�v��$"����ʳ�<��(�S[�bU��6sgUB�R�̣a�3�l_�,WqQ�L%OU���i�௱Ѻn��p�=���`���G��Wv�����h�P$s5��Vd�V��m�񕦄�p�f�f��ԋ;����#4�"W ���������1Ƒ)�T%�;K)2r]�����q�N`�N�&���]��	h��am��R3����,�ɥ�s�R^u<g,ڳ62�AMc0b�8/6̹%[�x���"�-��ͶP7u.Z6\ŉ��wx�:�������3�(m�w���A�j���e��*J`��b�B�t�5}Ge�p��
��)�Q��P�\C�l�˭�����%�C$ݪ����R���A��2Q��gXo�'7�&6<솺�V�py�*�+�NĪ�"�ăm�I���w�h�puK����SÙZW3OU�Um$q�q��xv�P���V�f��J/�h��o�`����sXubz��6����/��FVh���#��}!�Wq԰�WF+�Yj_h��X�LY��;t	#1��j�J����k宅�vh�zaY+hf]q��3Z<s6�jdK!��|�7Q\jJ�N�ޚnR<�E�%�U���0N�:w"0J�W����$�gf��1��3,�8���Y[%���9Vjv�wY��+g<� �:#[f1�΁R�!��s��-��#0ֽ�X�O��:��\ y�㵋e@ٵ�����@�PaAt�9�]F�
o����/�f>��L�|j�4��3�`wD���v��l�{������������U��m0����@K���*�+�����9�L��ʻ�����X����C���{�d�WF��I �ha���%\\��{���I�VSB yy�8�_��LkZ�v����ٻ�oq�t"}�H=Ь��ok�[�U
�Ƀ�,l�\�;�JM�/���sV�$��W�i�-��u�����k�<��e˃���_+��A>�wz\����&���r�A�#��a��& �Z���le�������볱��,}�Y	��t�s��e�K�0KJU��R"��K�����ղ��d��Y�v�k��#�C��ˉ]�]�ŕ�����3&������������( 9�id�Tkj�uv�����5��|���� v�ûړ#���4����0;���P��zݾێ�S�"Ʈ���ͺ��Y�G b�N�A�OG�༮�/��VV��P��H<!�����r�Ћq	��x��i��e����T�hh��Ў\�Ⱦ��S�5i��ClC���������ZPWØ.D�V��n�ޑ�:u������,���T�T�g�J��p��wg JѶ���	ic^��a����_N�Uw]�k8�!��sCSh��T]I�k��7��U�����ś�e���Q�R�r]��k�-�ԙ������uz��T�hD\}X�V���yk�C�V���;Q�);m��z9�M�բ�{���G�8�wW*��lN/����8zV��Nm����l�Ü��,��ҭÍ}�S�(X)M1b���F�4t��"îG�<�G�n��S��T���s冪�3��Ho�vܼ�K�����T��c7�\�$=�JG=B�ems���O�+�y;mT�Ӿ��!����Qa6�s��5���%i�à���b���wD]dÝ��9|�EYUo1v<�>��eU�0�&�Ʋ0;UzgZ�GF�$�o*����CɈ�F�u����vcn�v��Vk�E`�7a쭷](�By	G�t�먌:;Mh�����+iΠR���L��]��
�m'�(�%�t�.���B�i͆ib�G.���z��.�|��33/r��4VS�w)�cYM,�{d�T+�S�����k�\���f:=��ͷ��E�%=8���6*�9�[ޤ 6�8�FY�/$=�g6
g��<�衤�S=�g��Y�S�)}Qn�����H֊������4��/��gf��˞,��뾩͍�1juO���:��܊�:��[r���%CE�w{h.yX��WC�2�y��Gy���Q��wY�!L=ʙ�*���Ub��s��'�:�U��s�n.�\;C� �	Ř���*�1D�����KnՔ��.چ��8iɂ�l��-dy��7��ԁ0V��-z���*n�*Z��vXz���e�F�A���u��I�]\ˀ�zT����P�n�0��ܳQ�H�Z�g�x�X��Z�sYu�;��7���=1LV��ʲ\m�µ845��77U�իy�ܯsJ��$\��������r��V"s%CĶŕ�:cNLt�d
\����:Y��>��[�jiwZ�c�O��θ�p����!�з{�Z?e�B����rӲ������浬c�  ���2 #iP=����A�q������k�C��K��ђ*���8]���J��>μ(bLQ����\G�%n�͗yʸS�̅�W�:�[��Zr���n����� ;�_;��ָ�Y�qKG%m;yo�ڨl,Kif��,VnV�#����K��ɰn�Wd:F�u������dB�qC�9ZŚ5�Y��ܙh�=]���mYn�o�RG
vwMpǝ	��Nrs�Ǉ]�5�UJVu�^�P�T���F��z��t���5�5!:ˋ�oN��'mq��h���XO{mvF��̽D�n�G�uڶYV�-4)��F.�����+�����$���U��/���
#�H�AfRRy
AATVE21C����d��q�j�'0S,��
���1a��"���H�"DCJH,�e
�M��Ab���P��,)�sE(�YAM�t�n��i�*�)Ze$R(����ImU% �%:I|��"�#B*���K4��ZIIB!LR�J���d�ҝ��j0X��UW�_os����uE��{�ěn�-���MpՏ�������q/��?�����ٲ@�=x{q����{�)|�Tb��H��$`�(�p�
ʿK������C�ۂT~��x�1�Ku����RY�F��Q>���E-	�0�"���Ū������mW��1k-���6�o)��<�8*U�B�/7	�������t��d�n1��RD�`�>���G�B���|Q%r����U�)ʫSW�NO�_��!�Fu�b��ۗ�������J�߼ι}� �;����@�GĎ�{��|�ܧk3ymC�E���u���iC0�}����z�^�*���}z�����-�yhj8�<�c7*�g���,���v�e�:"n/pZl27l�O��Q����_d�ס��X�Vg�5w��),9N����ݕ�"'�d37 i���kw����B���:�s���_@����)��f�P@�``�o��	u�Ʈ�Y�S�jz7���^ưح���ݜO�pu=x�P�/u���
B/^2[\]�v�y��1А�f
;�V�r�:�ui��sA}����p�J����sa!Δ����Fu��]`RR�χ�RRsn0{_g�n�$I���t�P�U|���2��,���?Z������V�����&E���� ���4��.�P���Gc�1"�Q�{XMv���F�ٻ�v�-R:�x(����Hکtqc�S�N��a�&�{����8Gga-e��p�s�ت�U�4�[z���P�j6gU����"��2��.ņ;�se)l��K�ed�c9��R�X��%
�qC�	��ѕg�w�_f>�=�*n<8f؆�W���-ó��E����:{X]-�WS���\��ze����jF���t����W���`u(�͇z��ү9b�����+������'#Ըۋv����1���*�Z�G��^0 e�dښй>wk-E�M��E�c)��{c]!v\'Ɔ5��f2�o9=�x��X����wP�����)��n0=�!�'�A�����U�3��9�v��(���r�MΤ
�;E��ށ5fբ�	hۖt��o���9��=S,����NlЙ��nG�j�)��+���jh���j�BA��o������U�%�8�56��SX��)���B`Д�.;]i\*k	{p�߳�xf�k��T�$ްf(�����ӂ�Ll�39��e!���o��v`���ol�W�f��CF4��.�9u�囝aXm�kz)��k֤³����:�,m�g-=/'�7��Rʶ͒r�J5������D���5�=�[{��(S䡎mm���M=Y����T�ĚQ�����׃^�\&zl���F��N�']��j=NtZ��k�d�u��vJ�%a�(����ڽ�O��~�k�\/���x����A�5H��]^���4p \�h�פp���0xW�����BV��V-�UrS����[�'�Y���Wv�a��K1�#�U���2s3k:�U�|8�#5�>�]�C���	W�0h���WTC��3�s}d�����؞�4��DXۜ4�7D��䪳f�{Gn>�~7����ugf ��1���y}I͟>��W��
�y��+t-X�t b��n�̐`O�[U�\W&��5�T���a.i�z����y��A'���m�>��yΞ��ǃ��3dO� �Dg\#��%����>bbݖ��d2�@�Ԅ}�ٽ|u��7�nr�(x�FLy�ɂ�o0��������~� G �q����ᔰ���%�-��Cgq�����HQ9,�0n扱g״
���&׋\d�B}�lfǣ`yo4sŜ�I�Ԭ�<dڽ\�.��4#���-ݘ�Z�,h��G������*֞>�{rs�S�bSL��^7g��u'ڔH���W<�&p�%u�"��m��n�+�m1��:�KΧ�<��@/�`���I���6Z�i5[�r�fz�h���Le�ΩX��QY<{t�i<��C7>���h��q��spc�\�l�MqF�f�ym�1�ʄ7��Gs�x��U�{k/�u���A&���ۜ�"8��Q�LՋ�ڤ��l��r�AsZ��^8��K�;7l�u����t�L;���aY`����|*ϻw,;���eԧ�M�	�؅��rE�5y�Lէ�뮈��6w�� <�W�2{[�\y=<{Ў��&i��U1Z.S�ַ{0�}Y$+��P�����wV
 �4����e-ٿ:����l����Ԙ�p���Rf��AE.L�X�.<�̧��J��������/A���o+��in�:�a��3%2ά�f���&�����^/^�XY�8�����Uo���-�i1�cm�βa	��:z{���h�W�5�D���kL�����n�g=��r�/7�v=��)���������:�=�����)Gs��/s���%���Ut2��k�.�혞��;
�v�3t8O�\�XfN���o�`��vE��ӿL��x��Н���!�F����-��lO]D\�����ʔ�V�-�,�Ml<2���c��ʮ,.|6Ȼ�=z:`� W�Z�`g~��q���wǙ9���$*�z�Y������c�J�+�����k>r�Vpt��z��uѸ��ĭ�r�j��Y��̈́]Իt"&�Ga[�1h$TQ�/��v��?c�ưe�=�������򈽀>���V4qn*@���byS��!���x��G%�(鮮5�EqWI�`)8^��������<�C1k����ƶA��gtHp�T�j�`��lWZ��R-4��b �Li�$�=uX�����:�P�s(����Z��7bN�F����jRf+�n���c�k)�,�5g;�e5Wve\���}�=�IyF����]�;p+������'�(D��o�E�i9Z�·��~D��Q_r��DM�k*��hNa�Q=��3��U�6n���Y���,᫂B�	�(��7GR�>�A*�,;{`��G}z��᰾P�2�讵St���V8ܭzz��<�hM�w����|/��2	�����ˊ^�T�T�ۗ�+�m���jv+��v)���|:B��׻Ќ̈L�V�S���՛��f4�F���g��T�#�����ۯrC�.����َc�+�}�ev��4���n�n��K�5+��2[���aJ����ZNv���zr�=OeA�S��j�h٘��çi��;�Di�n:R�����q�ӽ�{����{^>�Z��t$F,��B�AV�iZT��*�-�T�lR��fY6�T)��B��*ƩJEY�(�E�2�e#TJT�(���AU)>l�(QX�%5t+m�i�
C)K��U,�e2(j�-hhB��dU�V��)�*��Jm��e
i--��4��Q*)uB
E�U2�awB�#t�"����J0�l�-�P�T�4Ȱ�Z��2�H�1p�$0ȴʺ)�FVa�U0-��I������KIh�TNJ��O=}���P���T���8k�Z��6w��В����z!����!Q��">�Eb�]�t�U�U����Z�����{�	���^��ꪱ��+1�T�go�=�y�=�Ӫ��3ww���>ؒ�}DOYp!�������W`��V0o�4�Ԃkz/����s �e���}�Q�y/���c5{E;�G��t^�}��T#ӏ��<{�aǨ���롷%"c0 �>�9���n0�׵}�MRg]���Rz��2��+Nu�,Oe.TW-F;��lY�I�5��;i�v9��N�S��5WmN	� ��25g��!����wӂv��6�����>(��ǛK!�N���Ų�'c�����@6zk�؆��%ᩋ�-�x밦z:�jbT�G��J��<t
�
Ӹ��:�׊�=��*���ʋ�f�y֔�ޠ����条.�\}4�.�zo���Yl���[[���`�����-|T�j9i�H���kwi-w����:�"r6��!�{�LBr��M;�wڷY�u�U3��J��P�6���8��6�З�.T�,(�����DGp�F����=0�H򸪸�N0S�W��b:��nƎ;������4�����B�ԝ�/cV�L�/��`�Gv���y|㞦�ނ�;%8]_�l�
��^�!/s�IӛK'q�A�24�R�\>:��l��m�VF���hU�}���'��N���ޢ�{��5���]}T��{U����^׵�C$��Ri ��r��I0���I�>Kd��m��/�!�Cu���|�w�1�o���U̠kj���jZ���4�K�Gg�E{�b ?Գ�}���x��7�̬��II48�Sf��<���ވ�����@����!��B�$6�8�w�l�RBm��L�Jd�]�OϾ�u��i�*C(!���4b�6ɤ�M2O2N�p���P'P�!�M01��g1�k7���s�O0�2�]C,�d>d�Y����2�U@���	�ZN2B�RBj�s�b�ƻ��l���`YT�<�>L⡤�}��a"��	��!�I��I���ٽ�s>���&��~�!l�`(CM |�`�
C䁟T��Hm�Q�'/w��~�۾@�I�4�q��C��Y&�m��@�Ha:�4���JB|�<ç�_{����5�0�0��;ʂ��3��<�8Õے2i��q�La��a�*��}�k����!��$�R��N�`g�C��D�d�)s�$;���	2��ލ�η����[��Ba q$�$��y�<��C�r�:��H�q�����#���s�vK@8É�C��q	ę��Ba$�>C?T��Q������&���N*�Fg���c�� d�)���jd�Q�Y;gjW�����W���e	^�'7�\AuW�J�Z����|^,��u�g?�wY��}����)-$�g�CHJ�����6��!�I�|�-�5G�!����Y�}��=��M$��Y8ɎԐ�L I0��m�i���
C�CL�By�њ	��a��{��*�����_Rl!��'M2O$���&X2m��L�00��Ql��v$k��^/Y�	�L��� ����a>;P>I.v��$�$0!�m	� �&P�,�\z�����`,�D�O2�6Ì��4͡�w�2���H{�	� ��?j��}�{�q`Za�>O]8C���T�Y:�3Rd��CIԘI6z�:Ɇd�es�}��{X��߾��d2��$��L��q����q�L��D��VY'0]@�	����<=����zI��'�T���d�C�$�EPC���3���8�b�C���q���;��޾I]l�	��
d� u��	6�Y&�a��M�X��k���U��5�w��4��M��Q!]��'P4������'�� s�$2�I�M�M�e��+:�g��?)݋��X�o�cwU�xD��oi��f�T�Hۗ
H�B��o�࠙�F��5w�6.�;��n�s������6�����ׯ���I��JB~���I�I�5-y��C��(�<�8��@RM$��kί�Ͼ�%����*a�q�<�m S�<��O$:��j
I,� u'̤!���j���w������6�a�I�j�̇��l ��G�C���w�W�Y�}�Ru�i!�Pd�6�:��KHL}A�	���H[!������:�>�\�u����{��hC٠��Lz�8���$�L2i%������	i�Z@�ʐ�����x�ڽ}�}��>1R��y��08�g��d�Hq%�N&�L�) i<����~��w[�B�@�'�i	�Q�63G�BϫHd�L���|�[�f�����q��^�=6�xI
|�̇����O!��HV��XO�a8ɦRa��HW����ߵ���a)�$���Cl��J���	4��L$!�u�m�wGC,��K�f��{�w��j�a�m��L0:�d���a���!�%�d��Q!_ou[���2Mߍ�X��kg���#���=����÷r�lcu/. �����;*M���;�;W�#���"��ђM�L�8���u>�I�q!���6�H���E(|t�	���q�0�g<�"YhB��|�>������5��C�_p1mH����A�n�3�������U����Qs���/���˪�m���77�֋��p7K{�܂t����Y+5�}��k|�[9�s��;��t�%�f��=M%lrZ�x��3�/rj5��f�e�;�%Rd>����Ç��x�^J(M�k	�d'�b��z�ɱ�y�w�{���*v�tgf��0�kC;d��Q�m+��z""<h���S]��Wx��$h7~�r��ȝ:���owE^[_����)}0(Onӫ͌[ܧ�@����#�7��x-��Foq/#Sq������c+~3�ɳ����wM�ܟZ���#���������Y�qOw0��v;����\���q�g�����Z�i���"������c�ۍ����/w&��"9Cʕ01�0�d��V���1�m��
����mp�������,�������[V^V8�Ɖ�Wv�H��Zm�[%$3Q�G�۹��?�� �OƜ��Gҽ��r��Z1���X���\�:����f�y�'`��8�el�	�vչ=�႒�6b�����es��o>T-���kut.���e,}q����l�^�˅��ɠ>x��bK{U�{}iD�M
�8����D�P@��;�(��yC˳gM+����~ց��8N��l�;�����Y�k3(���yE�(O��FZ�tȻ3��*x���rU���s2�$֞+Ӳ�R�����-��>�������>/�^�fm��\E��!V'8��-s�%����-�\��G8���Z�T���2������XZ�B˅�^�3�i�xd�S�6��V����*tle�zZ@��F��o���詘��Pv譕Nي��l�D�ܖ�\hC�e$��U�1����kE�N����6b��ni��R�=W��P�߿T�{�?��%]7�z᢬����,�oB)7t��t�ʩׯ�~���Ģ;{�
����2�2��%�I��D5R�;HT����̫�}C����Sv3KVn8�l���i���u�2ͻ�����l_�<7��*�	I���%mS��n�|�]��"ǳ�ܸ̚�R���̦Lﲰλ��Ӵo)�Pg6	�]8��:g	3l���ׯ1��5�V�'M�Hɢ����1�Leocy��/ h�mW��R:���0uu�jP=�Iv�
�f��\pDj�F9�NM��Ci��f�H��^�7��c9G7�w�w��n�L$o1e�RR2HT"v���ղ/@G�V�L,3���K��c>�w�_L�MoԮ\2�}��m`=�ل��b�U�i]�[%�,�Q�	�N�A��F��;y<s�*����:Z�nϷQ��}e֓��i^]�*�wJ����[��'6>L�klcq�s��)�VOqѺ%��aӃ{�f�<���`ꙧB[o'@i5 ��"p�e��N�C�zJD�/�<֜��N�uªtlnR��� �����c̦��!��`���q�۷�w��
Sq�,&ء�5��E�vRt �F��}hWE�q�C�,�[ֻc��t����W�!^=s�ˆ��/n�$4�y�w������yA��rĂ��)$�~z�?�=�> |�1R[-�1L8am���BИaiH�`RC>L�,��ZT{�AH~%$2���,6�����0Ȥ�&6�0��,
a1�h��5���O|_q�~W��A��iv�!�Q�;�m�6�q$�C�Ғ7��D{ވUۣ��.4+ޯ
�ű�P��NV*׷��5�.��ߞ�04�MO<U�E���Q4�^��P�y��Bg����s
�b[*!x6���9=Eb���㤎����Ʃp�Qi���UE���=d�Q���.�_��k��zMUq�x'�{1�T�J�
b��`��8e��N���l�{��̶�בrsԆ'R�j��f�B�xn�s��y��Xk�O��-�RP�pU������z�3�����B��K;��-��o'��ǎ���Z$��58I�xg���B�,��p�K��&��ۜ-���#�����&׹��s��>b��������3���7Z$���GC!��#v��_[[m�p�mDs+]�ux���ж]�8�>�}��='�jp�ؚ�=�����T����L�'�|�'t헏�ξ���Nt]�8N�v�e��l: ���f�"$f �N��K���]g8�ڛ�V`�Vi���}3����V��'[/�E)�<���j� KY�g�L&��7WJ��tw\��{�fo=��� WM��vTO���s-�;!��Xu�i�j�:�|���Op�� E1��s��ݵ�R*A�����c�[�13�,�.�u�\�S�N6���7Gث�d�!�1�l�+y���5ު�H�6�3Z�F��y�m�|8d�&cDY�qq�7�mb�>"m�k��4�ѻ��c�IK�
�ر�q�ii5;�w;�vs�'
�/-�NY����U�(����BŪG>f.�)BNW_LV��(�*�*Ճ��Y%$0_�"=�|#�1�:�4�w��$�F-]���{�"�!���j�/u�E�*�+pv��8�k��XEm_W�vy�8�\��{U�j��~V���>�q�Y�n&�>F�%�-��5�ԅ��m�\���S���*1�R������)�\���`�w	���a�ԙ(a16��S=��l ��v�z�=�>���<,�y�,�$�Ѳ���8���G�fXV��*%��S�jF�7���d��7Vx��k�z����{ l~D{��D%��$��@;bcf:�1���̳��۾���=�Nݦ,Tɿ6�l͂�����>�VG�ԕ����tK�~�.�`���J[�<�+�O���v�y;cO����(N�Պ�|�.�wn��=sO!Gď=�E�{�'l�E�+��d9���8�N6�5����̈E�u%GN��0μ��� �^�y�c22��}7�� ��'բb%�B��j�I�z�{��R�	�|��~�Ec�K:��ĸ �ʢ��R����(�����D{��	(�5��v��_lqR	���`�e3}V�:�N�f���-�vTM>�����-�)s���5���\�3��F�Ͳ�X��۵1�c.Y�P�H�:s&4�雜�y{��["����9ݬ�{��)'�>�ͅ@}�)�[&˓����~nelY��N�!������yty�G͜���W�o.=��b�LsѶj����ҷԆb��R�9���%��>�RU�d�
�����j�D-ގ�pRB%N��RZ���+��c���ﾯ���w&���H_X'�4�k�Te��恘�ȥ��e3�&3�cE�^:��9C�0����_h�0u�H�IH�q]G��U���]g� �;�y1�w�W	#9X��7��QC�և�ۮ lu�W��N��W������=债�`��ŷG2{+pC�$RTY��^�� ���S�Ѩ�2��Sf{6�rPhvx��͙;�^U�X�
���=Ĉ^W����GV9oC�4�n��%��u�/��<�tJtq�%�љ3j��l��!�l��nJ�z"=�4F����>�o2uס�'w����S�Ӟa�ںJ�e�>7Qt�q��è[ܪ���6BwU��-���p������MӘ�J�n���E�jƌW�m�0�r�c��Ou�z6�c����uF@�~�K�e�̒b(ؾ�����Z]�M�}W�y��b��殔���\s�72]WB�+Ӳ��yQ�Py{�d@v�e�ʋG�k��������ɖ�"Ĩ�o��+��9�lǹ��c���\6_k�`�z$�p}�G�'Z'4}9a_y��U��*�Onv�43<��w=�Ƹ��6ҫ�Jɼ�޺R�a1/��N\��kb���q�N�t'�t���ϊa��F����ѽ)��9е�ݰb��v��;m���#`������M�6�/�o:�bx����Ź6_<��>Ս)���&�:����]9qn�w�fʽ��<Րy��ya.;!��(�fQ�J/]������Y�Ǥa�Ug&�+m(�DV�7)K�d�;;��{z�]p��i���v���HDG���Ē��1�3��jbd]&��+�dT��}��mZ�++(��j�u!���(�%BG�=Мy���}j��Y��6S{��t��t����]����矮��e+�K!/4Kʤ��u�z����>U�����<E�$QfϽLbZt�F�!�����z���>�f˙8��!��m�h.��J9�U�eoުa�?�"fy|n�e����ξw�0�s.JV��߫x0�}����㥑H�w�����KS�4�<�-ԎK�b�^�9:�Y9����&\�㾟)2e:�:�����\�ޤ�h���U������|L��1�.q���u.�;��(�r��[y��x�3m�{;H��
��J a��NG�Ve�uK�j3���J����ćz�\.n�5���gؒW��Pa��f�R��G�kHv9Y��y��_4YǙI
l���Q�����E8gjh�9������!�H�}���80ܫRH���I��
�{ X�����I8�y.�N�'k{ن�u���CQ�՛���9��8���P�{����U�y\�����\��-���}>A=�X@ι�SdA�zk�IQĖX��tĶ�No#�a}��1E�X?>����Cm��`��pP��_f`碪^*>S9ÐC��W
�V7�vߨ��t�m��+:kGVڷҸ��������y!�����:2��e["���o���.�{��|%ϛ��fݞ��[��#��d\�1��¥��h�e�aG��r�.w��<4Ӈ
�iv�kj둶�`����ʍ&6��2�c�h���	��H��w��#��g�T(e �u�9V.�X{��-�H:���л%�*t��������w�Qr��wr�ǅ�k�[��;�l�_hw$31����9��m�J�l&�v�	ܺ�όro1��V�v����XD��e1��*�;��������޳]�H�H.I.�J\~�D:��4�)���
Jd���0�I��y%�ILR�P���O̦a�`[&نdYEa��X,��!N*�X[%002Ē�*�b�MHJVi5tAb3Hm�E6���@-�2�%2C@�3���6V�捷ϵ�Wk�p��ޅ�a*�ït�aTV����z"ZN�r����ʌ��5��Tό��X��JnW����)�
��)9J�ab�F��\����w��ǈ�8��0쯚d>��)|ٞߨ�[������>O�0Z���Y��B�I/����C9����C�?�mcL(�u�xЏy���DY/֬�O�ٟ<7]�V�,Dyz��J��m`?x�f/v�������xK��ɆJ��E�~3�-U�AT�e""�l�{h�*vp���TEgڄkǉՆ�!���
o��2�5D3i�S�B�Y��$fk\�<~A�;�ܫ��C�-�Y�9�w ���{MNy�����n֚�u�����v��l�{�T]y����鸙6#B����X�"=�Y���O�Fb�ʚ#�9���`0�|���痫�fP�No+�:��\��Ux�"�S�!5�gc�����5^a�����C��0�_f�x�:_�VK䎟Z��цt��i]i�<:������YȲ5���_���ÄN��RťZ���-r_u84}�1��X�D_+4Q���[��|,�v�z['�H�ޟ;CXY#ʂ��*=�M*a����+� ���<F0�6��+z(��W_"�ť��դ+�z�� ,�Y�xy����ρt�Za��Y��^#7ީtV��]���B�J�R�n��a���(��8�Y[�vh�ˬ<��8�]����X����W8OL-C7�yg:|�U�Iǉ��+j�~�S���[�_N8HT�,Ջ���p�~��ˏAON���o�u��lM5g���Q�*�FA�%痢��_��5�t�r�� ^�:p�V
e����W��P�ޜI�ψ�AR�Z�F���?Y<�����:�Q�v<�.��R���q�L��7��$��}��y��0�4l��%�<�X��!l?/���җ���W�j���ԽQ�(y�N��j��z�)�8�\�	h��ؕ=1���*�4�6t�C����3\����s�x�8�>���v$�̿TA�-���Vi�R�
���U��T��wtf�pvL�q�{���J�z��|#FwZOe�w��R�t�LV��\u��'��v�:��X�O�0��c��X�7�8~��c�8��7f�>,�lN_c�/��a%Z�1�>#��7}�(���6CK�9i�6�\��ZH:窳����Y�d!��d�����3�/o]���-G=@\�Ze�����d/!g�9<>ͯda�Ǐyy�?aq!��#Ŵ'5�l����MYӧ�����i����-6�YQʾ?^��I���^4x��E����[�D���=Uv뻤��|��b'�l�k��3ɜ�sT)���S�8F�0��NA��֚A{�nI���r�Ou,��r�&��N��2��e���X���ܖ��gR��}�����G�-�.��̖�a#��'��=9�]�ڏ�u�=qp��g,�k���%~cI��n�]|��F%WJ^�Lr��>9Fc�ɘջ�y�Fߵ����:M��Ӻ���[�<'��{/�L�T�� N�g�qC:m�Q�R�㕔07ɻ�UW�TkW�Q����b���#5����Y�uz���_x� ��t��R��y��A�p�b��ߺ^R��<F�> �~VcL���t�<]�ӓ��0� 4z�>L0h�h�*�,�����̷�Լ{���b�zaX�#QwF��EV�����!�bl���<~X��i�;I�͝�M_�r
���_E���'026і-n������/l�M蛼7!#Il���ZJG
�6���=3�SN�}�-��M�����7�,�.^��2".�*;�OD���^�́d
��m��=�-�g��ܧ�5Hx�+0�F�?0�4��:�%���w=���!z5�\ED0�"�Hɬa�����G���AVX���:Qˏ�h0����ǳ-3S��pp�Cm��`zx��K�]�H��ozV�zeM�הfEû��K��ʄ\P<͢9*�&I~V_�r�>"�I��!��qU]^���>\5���<l�~IQB/�x�=c��Y��^�UB!�>������haH�+4Q���/�UE3LAL�ƃ�1V��ƹ�=2�v���,��|IRb�f��qN��x/�X�Z�6�F�H��#�֢f���o�~����&85��Q�n��Lv�ӻ�7��P�y�]��<{�:|F��/G���;�{�ͥ�
C��
�i	�u+6@[�)��9�ڢ,��R
����YӀ�U��ws�Ue�e�#��P�� RWw���Ϙ��5�oNU�SNq�Zh��Ҙ�6ř�+ˏS�����ն^��o��f�sYQ��S#"����We��F<՞k��OZ��5adY�n����Ce�$��ZC�(�-h#�av�Y��[��D���G��B�+=J�ˍZg�o-���\��:�Y޾�9�u�a�O��Ya��ӫ�svnЧ׭�ܴd_Oq�Զ�j�KI��ވ����F�C6G�Ǝ5����!���a�[	����Owx��N���L��Ylg[t�<�_V�=��eІ���H�(f�����#����u������yX�Ɯ&�˺
No�ͻZݢ�������Ȅ�4��a�>8G�h��W��K�"��?]�8��l�#�yv��W�!�:u������Dm�6����`��^vPv��/T/�Ed�
��ӄ�G�ϳ������ز�æȳ�.}eK_����{��=�;Ob���3Xb���(�u! ?Y>w�����6�Cm���9��*sڅw�C�T�b����
�p��a��*�K0.+;�CY6�w�Ey�-��﯌��~�K��8oP�!����cO�
:o���f�v���A"!g�i����<F��+;���ݱ��I�{P@��uQ�yBO����<f�ew\�P�9�!V~��q�"�#Z$~�7�z���C~��S1��^�s{�˖�9�ەt*nyZ9��?X>#N��O���"��!����~��fȲ�ӏČM����H�>�!{\�a4y��!��	���~�C:|Bs�ywv�mi�����y��u��^�+�W�꙱�E���N���^���P�.+m��)9Y+��]g���r̍��B6$I{��¢s�eV�W�{D`Bu^kU���nds׷��s[���͌>qB+ '���E��j�c�߮�V��i�_��_4��^8켕�{�Z&���yf�#9v!�*�'���w}ɮ�f�6}k�_>0zޝ#���!�7�7J�4��,����1S��*�Fl�?,P�j��G���s�������?x�oW��bj�_�fW��7��Y��G�l�l�u@~�زf��W+�u-���c�}�TE6}�F��:��}���X���#g�h{�}��(�Q3<���mιHn/�*ώ��Do��9��2|=N�z��B�X#]1ڃ?`����q/�� ɃRˬyv��<�ա�0�[�6oelL�pܡ��{1hUݚ�Wo�|A*�k���,ҫT�Vt�p�jR��w�a��I��OS���0w]l�˲L֦�l�#;e�o2w#ҍ�&��}[�rg�`�2au.���J�u�ؖx�G�B/��AR�Q�O钕��vՇ�L����c�� �E�I���g>ҫ;ls�Y,ҌĈgkQ]4I9��.�iUs�72Gk�l$;��[i���8<U�<d�tK.�ޜ�t���E8^m�L��h�)�mY��f�t7:��4�Y�Ա�ڦN;<��.�	�ԫ>��[�-�,�2�p�У6��^X��|`���-�噽o��"�.�=�:xL_��X�w35��A�f��'�����^���p�2�ogU�3n���%�P9�<Th+�݋)R7:ܾY!�\�|u]�o��]�����y��s-�X8e�z�}ɶ��\��q�w{ؠ���=G;�j�¢êGr�N7��v)�B�>$Y���븍���k�[��NRt�ѦS�&������4�œHsn��3�c�F�fr��ٜv�}��,Xk��$Xtxb��]�b��ӸgL�Fƍ�[�w�$��l����dT�p/6���R�<���Z9e��Wݬ���ެ"�ޣ�0��m��*	��V�I$��I)�@��z��2�SUH,"�-�4�4�(H�(r��%�"�Z��- ����L4�d�$�-�r�BI
BS �T%"�e�B�� ����$X(�E0��H��Ѐ�a�ҊAb��P�L$3�>=}���<��&���/f���h���_wsv�z����jݫ�/���D�1�%�~�?6�˵.�qt;���(�X��b����+o�I����[)�EC׈� ��Ր��./�x�!�i$w�z�j)�#ڴ�ǈ:��#�������������P����'Z��~�����=)���+���IZ���A��x�p����nz�:||�ď:@���V1�Xp��pB}��G��G��/���?UkÞ��B������A�P�a�� ��^�����B�ެ�Lx�!甼E�צ�C�\���;�²��~��ҠLS"����F<V��kEwי��"�[�O��f2ޠ�r�- ����tE�]+wo;1 9N�)!�}�
�j9='�'��W�#K6s�!�JX��T��db�3V�@���ic�O@�!��5a��<�wP�6a�-0�"�w�M����)���?Q>
�Ȍ��jM�v�a�S®A[s9�����7ꯪ>\9��IdO�z�>�#h��'N��#�R��|!��q�5(�0��ś?x����>���L�8j������Lo/��>,�G���ҽ��SC�@͚�
�ɩ��U�z�dH,*�	�M��m��12�By@p�� �|f!��4~�܉w{w�4�P>.�r�،i��M�?m������R:�;0�=lֺ��N¡	a���[Cm"0�6�M���<�������X�G��}.���'��+��^�}������ś��K�'=>2��(G�^1wu_{i0,8p�yB"�	*~#N�����n4�dY���X~����i�O����y�Ua�}ye�J��C�qӚ�<��H��|7ձ�ߢ�zX��
r�><j,8g!dC;�Lic����z��n�/��k�Iy9�M,�7�o)��v��������bՖE��b$Qf�g��
���y�f-����:F���a��v�q� j\}��\��Ƀ���_D#_n�3_�1��f���>[�;�cO�:E���Zy/��~��<-"l������.�z���[
��5���x�\N���f�)٘1s��J�o|Q�#�!�}�a3'JG����r|٣�ל'����)���Tn�]�pUG��曩���|�㾌z./��:A��:L���MP�G�]%���Uz���!���W��{w��Oe�;)(��,�&���#, U>0RrS����:+�oc!]�����/�?�a�Fz���^�ݿZx|-zْ�}�� �D4Ѳ�n��N���^vh��,;1�~]:���³~&���c��c�˯FO�b���×&A�s��M����qJX~����`?i���B�s����OĻ�xR���Da���#W�`/-� ��-n��}˄��ho*Y�|���R�Ϡ��[�;�ג���.���v&1��U�mq.CӋ���,�͏Q��Q�R��U�+f6L��TT�S���x��vi�O[�������h�b���+�h���Y�0�ZIO��c��y�? |kW�gO���ǎ��HVE6�}L��^���3�\_c>z|Q�0�o��c�}	�_~V�Tv�C����uh�|J��8�PZ��g�r�W�$�)�$֦���m���W��}.�
����^!�~!J!.��Ͻ��B�����;ԥLOR���\�q�����ԙ�E5gg����K��v�����F�j�L��)��(����)����05Ǡ�GO��T0�a��{-�]D�Rq�:�� S��Vv꛷|E�T�n}�Bll6(��L���)�,d
)!o2r������d���*cf���ZB�{o�w�n��"FO�������c3\seˮ�~ޮ���hQ��3∣�	Y%��]�zXo�iC��a���Q��rBȔO��a��캱�Tv
~>��_�҃VrzO�"��%�ƖO_��nz�!�a�� WG�4<��=x_z�;��Mؙ��!�9��'�8G���j����tt��)i�93�g)W�r�;����οsp�
B�-C�8F�G�g�u!<�T����'�u�Pͷe����^l�9Ji37YB��:�4��>DS��⠬�45i���Cv����lZ�3��ơB�2�q����cnؖdWݧ��9��+��C�?W�o'�/.����w/jP�ˮ?���b�ٕ�xT��i!��'� ��!��$`��^l�y��u�k<tȾ�v�8Qd?!�e��G�}�q�Jsl�ܿ]��<5i�Fe��x�w�ǐ�,$�M:��Ѳ:G�j�x�a���9����ޫ����`V�7����9�b
����A��_{2�	�~#���C9adY�.|�2�O��g^��u���`��jv`��=8u�K���H��	yk��wNܳ�#���4l�fϼ��>�6� �u}�.g~���<�<n��H���圴��Ν�$���uSЏ`�:���@��-8�j����e�i���W�ݜ��Ռ�MY�&�U����������T��o�ix+@��pw�
�� F�$Qf�n6w��w��N=���ws�gHZ���k'"�/w� k�߅H)����Z�Y�e�h#������739"w㐙$�o�bd�G:񞘴��-=����пo�T].�9:dC=:i�����Ǜ8M[���Wnpk�|l��"��@��y�GAB�~k7w�>6Fb���K�<��F�?{4�]��i���/Q>aCȕK�J�9�U?#���N�3�0�#�/W��,�E��=�oVn^�}�Y�Fם�#�y�)�ڬ���!ci�G|r�zM��e6X�=��/���Z���87�*�n��ḁ�MuB��X/�l罓"�3�z���#WhDTO���/���v����|`��0j&O����j���[L���!�Ԥi:lա�y|��j�W2v�,"Zl�"��>�
Xiު�노�R�'
 p�
4_��9�30f�5�q���#�}U���w����<}hq�1��ج�"���T,G���&�GyC��g��x�#���V!
�gF�*ێ��w4f�9�J4���ǎ���z�g��!�.��~a��a��Z|Q�F���5;�x�1×�)2&�mrZG�y!�[G'z�Y��cO�'W��VY�@���^ >�a�@�.�-��
�X}@�|3�ܸ�6��6Z9��ܨ���;�wNIǣno���3�%��^�u� .4�\������I�P����é���Α�ȇ�h��Ew���x�r��P�����rk�,�!^�Q�cF�q�����+�O�����O����5W�{N֑�i	�⸇�y�]����r�Ou�c˿1��0�p�_4�Y��
,Wj��m+���t��!U�ah٢�Ӆ���R:O�+��u���5ԣ-a{b�GqB	����%�&V��=�3�Z� B�谌��0B;I�C�}�W�����G��x��Ӳ���`i����B�/��M󩷨���CX�r�j�5��-=����>�v�l����ĆK�(q��vҮ9�;H8�OeL]W�=�pv&�3{cհ堥s�|�T�pg�������l�r"dh�QT3]ͳ)�2�n����$��ma���ڷs�T�c�>]q�^�ǳ��ce�S��{R�XT���33�U�U��"�e�ꚁa��k�P��_07Z)k�S׎[C7�w�Q����iЭN�yE�0�qU#㋲eh�q��q��:[��S�j#�r����/��K�N���S&����C����E��+��V��C6�K���Hd���
�7�}L-P���5at�^麵�9y�z�����\sv��\�7��rm7���Ҳ��EVK/�D�:w�+�����X���ǽf�4|	���YQ&�s�wM���4tU�ה#�HC.��(�uZ�u�һXU40�.�\�eXiD}��H������|�v�0WQ\"�m�Z���W����p�%J��Q�m��1:��xl[���\�ڷ�c��<.�d3������F�.���Á�5v����Ϸ���S3�JH��`]��R��,�nھ��������t�7�Α��q+����]����+roP�^ԝad:�x�ūmv�ױ�c��X�����F����f�4�$S�Aw�}�E�\z;w�؊|�Y@���F�Jӕ{:����wI���9�������!�JH�"�Q�LU-���")�PE��I�"���X�e(���)�'�"���"�i(U�UG���X�QW��iiRꮨIx��EEb���E�e��m)�8JdF(����#2�j"��LEAQED�R3�V�H �8�9��O��wV�R��� ���j��85V��;~�t��^�zp~-,�@���<���"�<D�����4�_�߲X�G���#d�?2:��_���H�x�����ݎx��t�r\�o0�i8�k�u!���]{��vQ��Cܾ�x��AwJ����+q�y��}>�r�����b������������y7)W^�t"�Ҽ���&j�	�Hs�U�Q��|<%ʑ��tdMI���Y$��z><6�<�����I�⍔�A ���8�!&P������,�՞@3�E"%�s��*����b�7�o�`�Ŧb�Ő!ȝ�H��m����L��/V���u��,�o,)�뜁��Kw{+�j�2d�w���+z���g/g<���/�  �}�h���)H+x;�\ş$2�ŚM~��|��CEt��)���Xb�E��"��I��Vy!��9(��X�Ç�
Ї؆�}I�;�fA���6l���-"�8�-4x��'�h�U���dv��=M�4E����B���Ut|_
�Zx��X��t���,�Y8�/A�+�wd����k����3Wو�	N�}�����Ct���؁\G��zz7��Ag�"�כ;
���Y�Za>~�~$<K�3�{���2a��Z�dQ����N�ezi����[�q���{�s/��/:ȷᇨz9�*�wfc�&���uE�,u��������L�����ۀ������(��=BI��1b���ҁ����~���w���Ɨ����&��h�D
��p^V�e��x��s7�a|������_���Zʼ��<52�ƈ�H��]�b�؃�浫=���)|U��Ӧ>я�|���zt�kq���w��_z�l.i���B2��]���yASu<�ɓ���������`�C7�z��]�]��JA��܇�t�	a��[6��9I�j�>���ht�К��B��݊͛"ϖ�ѵ=7�;�8l�Xa��Z�ykW�B0�-
��B�;��6�v�'L7Ief�C���a�u���%C��������`�}��H��Wwʻ��v�MGC��~ NsY�wwt�7F����X���ӧ�ho���{��n��pxB�#�=>Bk/�yi���\�r���_f�p��JL�b�x��]k��Ϻ&�mCڗKÛ��5]~���s�E�/��//��'�P�#��d��7�����4w'���T�VNDm�F���ҝ�!������\F���-���R�v���j(z}��x�}�F���%ʲ��cƚ��� ȿ+�:��.��=��3ml��b>6Gta�aG��`������$0{��/����ޥ
��^p�	�#�����
��];�����Ȱ�Cd��(�f�����qd���k)V�|0�K��eG�4�����R�GI�}+&qΝ�{��!f�NMO��]�t�Ԧ/����q��H��C�|�k޻��2�̏v��,ЬY,WA,ؿ�i��-^єس)=�����1@�)�9���i���PD#�����k�>׆Rtxe�S�<���ƌE��b��DÞ�6��ʛ�0�G-���I�W��QRdʝ!|l���XB5򳔝�2�{�)ᚙ��o��B�i�ư��}�
����gB�l�$=��8t��ώ�E�1QX�װW����?�(t�~�'�0�/0h\t������Jk=�g�8i�y/�|���f;e���7j?�{�Ug�x"kA��&,Q������f�N��fzvc���Q��5s  ����yD�+�/]���r�����w;�z"�A����	��l_�+3��rC�Eߘw�R�.�z���C�1}i}�Y�퇫�v���ٚ��Z�	+V��;3�A�(��G����k5�{e;Hk�í`W-7�K��Y�.{��a[�ZF���(�-Q�*]�O,,gd>���$�O�Ҭ�f��TBv�S�)c�a�B���g��޹��D6~E�D�P��8|E��o����|!sW�h٣��G/0����<Y���Z�v��"Z���P;ˣ`u�U�i�m�]K����Op��t����#�+�����4Qy2��os��r�8�YL9ӈ�-<.��}��'�˷�}9�`�W��Vn֬+�b�s;���d�̳JbU�()���E�����b�K��!^�n�|�?�,_�g���ly���Or�����`�_z��C�,� ��H҈�t�W��[��=i$�)|ύc�<h{X'H9����^�p�x��y��V�O�W�� �r����\pӷ��=YP1/<F�$����Z�C#}�7L�o���B�h#y
�!�V��������h]�4�{o�
C�ٔ��˵LC<�?i��ݝ�}�0�~5�G"S7�N���R��5�P��5^�K���j���a�����;+�p��
T���F��Λ��v�3���6��KK�Խ�Wיۓ�����q�M-Vf� =�~���g�~Y����g/)�y�-��O�V�u����+=�޽}�O!��k��1�xl�0р����zx6�Y��6�#���
zl�*�p���A��m.ړ�
�e̵��j���y�Pb
!�9�#Y}]6���+�ǋ���a~_ p�Df�]�~����y�@t���O�\.����wҪ�x���d�H��f�D�%/��mb^#�˖���mF��,�8����6h�#W���d�3=^w�h�i,"R^�#	�^o�#M�g��w޹��OE���7��߈~\���W6mPm�.meG��QI�ﻊ�4~|��wR�u���Y�ή���b�-ؼ9�i����d����珲�7�	�}��׫��gU�?b���L�ݭ�. Tw!�
��k@ׄ���x*wqs��ۅn�$:��f�m���^�3�؄�I�HQ`j�Z�龾�1m�8@U�(���YN߈F�+�V<�i�_>#-
?e�x��K�)Ari��%��j�^T/"�0&)��U� �k�
!+Y�_{ں���B7�.sx��Ӳ���� F�՜��x����O�D"D�h��{U�@���+Qq���oR�����h���c礞:"�+��z�F�^��>:F���V~De��϶Y�}���N����uwKcס�e��ts`�w��1>��!{�]�a��U����Y9�r[�(��o��r�慺;�S��mTr�|��t��5��/�l�]M��R�W�8��8t��Y"ȝ���Z~�����,��"wP��3B�	�C]����X7�}}0'==1B����A��Q3n�ș{��ʽ(�3|�vl�t܏�ya!�Y���������!���0��������N�W׻eu?:����J�<����.Mצ'eLT==KR�Bn�Om9���y9i�Z_�,��\�xz��s.��Ez��|���'�/yG�<O1��ht�nn�H�~�TF�0�4F���L��7�:�wg\M��jO��t���L�5�V��m�>_K������,���C�,쳐�7�Y���)%z�U�`#�L����UUi9FPͲ�Gs�wE��D�,����?E�|O�Iu�>3�s���TWR�� �Qr��Ȩ��&��ٔ�Fv6��֨j�Z�Y+x�2��-6�ȉ `zV�[@��X0".�2��먙p����^�f\��k7�u��Y���tX�1�{��0�Ӓ���̩[V;�&~+E���fR���툭�>��ISqX��Q�޹�xH��;��hֈ5<�i𛃌��q1�D���T���)ט�'�vC�NHx����:ik`�#mU��|��/2�8�:��prć���.�4t�fk��0�2��L[��,Ӱ��J�o�����q�����
�u��ЏU�N���a�+��!�t�N��ܩ�L�e<}܌�o-YN����'iA�H�=���wf8�7Re1�����zfR�O���Wx�7]�h&iܐ~��|�%���7�,>�B(�Jy��[i����ox��we^�X	�6��6��^蜶|s֌���o3��' �\�8F�j�Z)��O�1J'��x��m.v�L�U%ٳdyvrs����u����1�Ӭ8H[�Z��gQ]�XW$�G�IH����ک������)�F(��H�R��DD"��L�J��" �"1�J��"$EL�"�ۺF�cR�YU)c���(�)BEi�m��n������B�P�4ұ�X����UCIWE(����)JE	U�
r�p�TZiS7v�EF��RU�V�(U���ZhR�U��EhX��"�14"SI��*
�
�$A�hDDV�Q����q��]_�N�rgsV3��d�T��j��2���uu_��Ѳ!x���4В���'(ɜ�����{��9�2�ͮ�;G��_�h��Y^��sQ�%L+���"j�u��X~�TC���އ����b��	�.S��5&c�X�ih����W���d���'y���� k����3_���Ђ���KI�3�"xvK�Wn�x�繙X8CR�q_�7�����W� �œ�!X�cحS1݊��:�K@�q�NŽ����Ԛ��W�g�^�V枡3�tJ,QCb�B瞘&$���w��d���q�
$��f�y�ir�n*m�9!1V	�f�9ϝ,�h��U������~���c@�������R��4Ө3U����T�Y#��1l�o����L`v&7����t7����)t~�4kP��������%��|�eq�h�Z��c��K��1��i-7�g�^�J��+P�x�:�N�n���:�%4�P�۸!�D��tr��3̊�>����=��B��y�n�r��ׄ�	��Ao�ֲ5D��]�Ty�8�{˳@�Q��fbY� �f��d�R]����.��I�\fL����xg�DZ��{o��H0@�ܸB̂�\
��=���e@@�qpQ����2��J,��߽[��]O[�� �j�Ɵ�����I��JNJ�v�����{�Ty�\��D���
�
��4��Թe"qw],}}�nz�"����tlg�\�U���4����☘�ӈ��ݧ�>�c=�i�k)K�\�(^S���k��anr��V;0��-�T�Y����n���Ӭ���ԚBt�.� Bޭ�C6��Iq�|l�t���PR�W��"+�g}V�y��ЅV����m���d�#�w��M��F�w�!��<�%snڸ��l*��ܹ.-
ӵx��oJ����*?EKUz�5�������@�oS�Ύ�2�u�^}X��>�=L�C�Z�	-~W��;f������CW��m���R��]4�FUPy��C��YZr�&.T]�~���N_
�P0�R6ύ��,���G�����aޥ\�t"�g>qmfj��DYT����ʧG�e�t�_0,���Vk���^���!����/#��k��z4>��@�Y�d����aj�����\�ɲb饳6z'�XØ��d����s2��;u�����Fi=����(L�9z�u��Q�$�d�׌���8�g���E9�ˣ��|ʷ��x����+&'����g��$վ�ډ�� ݾ70bǥ����ߺ~��fk%���o�Y���L���]�",-�0F���{u8fK{�� Ƣ� ��k�f�=y����Y: �gձ�ҝ=3&;��é9�:Q��!sy��UTk����>م���Q����&�s۸�v��Ɏ���"��)m����3vBF;��פ	���][aF�+��7=�w�N�� ��w.1����¹��'A|�q:����9�ėEn)}�ۭsJ�ec��׼�V��i&���Q��&%j��o�M_e�)fg���l�W#\�«Ԑە�ۨ���D��1�N,yG�oy�6�(��;zj��a�Ԧ/����r?X�z@��u g#�k|��Ά�2v�9��E�&����V��ϫ)5x,ob����rt%�}6Ds=��_Cmf�ݫ��V�|ϣy�{6]!z�����xL�5��TOv��2�
���yދ��sGB�ҭ�ŧ df�L1�e!-JjH5�\y�8F7u����1w{�fm��ASp{��[(��S2T%#�3��Ek4k�-n�
x����a74��(=�vv���!%���"��3\�d�����G+p����r��G�
�;��h�|/o���=�_E��ؒ�*Ke`*]���x)RJ�\�ޓw�T�.O=��w�Y��qcf�^���%w[H+]ҵW�X�{���Y�:Q�M�+�A��tZZ��n�a��*E�?B����e����8jg'dOI�:�7.���{���"� mFNk�8���ur�j���g^Lki�k¹g?k�� ��kҦ���F+�R�m@9������Ovܛ��˚�m����d����Z�^WH�����;�_!�񀗶 �A��&x����|��flY��mCcc�)��7A���b����pI�R��w臈�|����+���/6�o���&tĵ�:��޶;����{NRz�U��$9�Zv��*F�;��J�6i�u�	{�5�PS���̾���))����m����KC$�ί��`^����o�\���D��	��{^��!9"���<�׆��FXy7u���;\�5�H�����ў#�E6�FһSp�h��܋�m�xr]K�h�̖{���0FB�M�" R�f�J��v�^���n��6�)~�O���6�5�`����}q����wlqS����hkz���k���}�[W\�[��Z����.q�i��9�o��}�6��#v!���ȝ�lcʨ0)��P��dƗ�� ���^FŒy�g�9'�V �יw������tE(�}��;=1�G2�-��t��K"C.��W�"F��٨xfoJ�ϲyZ9~*jG癇>Ptv���#;3c�͚(l|��T2��L��+V:�:}ډ��k�����C�Ube�NӼ{&:�I^��H/M3/`�-Z'�G}�$9�lq��dۡ˨�A��	7A�[S�Q�(m���K�f�O,��S���C{6��Wb���gR��ZcfGNJ���gZ��k=U9��jJ�ƞ���L�zG+t<{�;�3�V�2���x�9��ĳ,uc��F��P�Q���Ƶh�,��7(��u�]Y�q�1�4u��wSv�"�ٰ�\�8�N�����X]��7g�s�/��w�\{��b̓vH-7���]C�᷄`-w]��2�)����w����B17����N�W�w�y��m����tlg9 �ձ��]��;ν�IЛ�g�ъ
cc�A#�WM��̸�}��1$�6�9{����]�v6����/��w��o����&�Z՛
�G%�d�B��������4m��X�/,U�w���eT��\Z�u��L��C( �1�:�k6U��l���h�薣.�^mmu���\z�Y�e��yu����u!Y��|5
���۶�1�bW�$�<ޤͭ2�-�پ�*��ԁ9���.���4$��,v�c��C��e��Y�ͤ-���7h���z�m�GYu*o�ru�zNk�w{���{�t�(���)b�*�Q�K(ȰQ^�*���V
1U�R
�*ƨ����(")1Xm�FH����Qb5YK*
�Mc.��iTMUT�"+�F,��b*�%[Q�-P�����Eb6���UQTХR҆Ɗ��+���"��T�(���B
",AU�T*E�AdU-Y��(�G��w�J���{��)��sDӀΈ�ݶt�g�6��U< ��o�룙{��J�C�>M��60��H��w����*D
���j,k�jon�7�`Í�@�1������⟇z�`�L@��r��VE�)��_R� g,��Uv��5͢�������+5��V`�`�Rj����1VЗ��d��GИX����,�$4�ٷYf�zg��'�Ӆo�u#����k�ɳЭ�����uq�z)�*��Lԇp�E{�횲}���V)���õ�{�k�e��'�o�\����k�3�Zc��7{j��%`YU�1�)�d�kw�}ۜ�r)�IwŊ���0v����w�&�L��[)�����s�2�fE՞u}t}�My�S1�����{�������`ڼ�yd:ݞ�̆�f{Zǵ��G�D��/7v/`�Wsf��tP�4V�h+�Ev�۔�g3�C����x.t�b�b���%�y�9zc���t��`�&8qE׭.�B{�\SW%������2/�}�&���n]�Wt�A{Q�����0�:9���-�����E٘�.	�Y�Ȝ��>���F!^�����9���#1vՌ�������������|c��E%���f2��X��v�,��n�j.�/#c���/z��e�Njޕl��%�l$DtX�#�p=�+��mg�6cQxF���.�P*hNӲy>�w��k���o]i�h=6O�)[��8X@o�?+X+4��U�
���T�ˣgx.@����<�U�f��s�'�v �S��t����R{��:s#evՓ+P�����E�࿄^��nlgO<1���ۧ��&�Q\�7omMg�.����"��ej[[�����k�l����]����j>-�ax��1����s���of�}W� J��g����i4~圤q�d�4׵�}핬b������;{pHEE���N9�����ƓrEFφm�f�7���w�d2^uD��=/K��w����3����Ξ��Gd�ԁ�����\y@l����+�E|d�5���Dh讣n��m�)v�~CC[o��^"ю>s��a0��ޝ��J]�u:��grP�%hyD�7���I�s�Z�)��<���mMB׃UX��euqEev.��w]�{�p�V�}�m�n�� 4Ċ�T�I�k�kO�`OF��Z���q�c�o �m�9�r+�X�PR�X�c�@s����d<9a�}:�c{��s|�NfgF�4�"H��=�)���=.z�(�ӎn�]tJ8v�7zX�b����3�K�t��N���+{�.c 4��/y�
�X��~�fLoR4�!���Y�-�}�d�R�;��1{�\N4��eڂ�X=@��t9uM�{	���ɤ���ǵ����}��){g��V�����F:�5����� ����T��f���y=��a�t��W���Ɓٯ���T(ٴ���O&M&��.oC���a}T�� �zz�zy���`�/)G������A�YU}v����C�|m����^e�%\(�u�*��Z07�7o�l�IS��D�P�
m+�����Rh��}��o�p��6[ͻ�&61���ƌՒ�ZN����rN\Q[Qn���	{7�u��~�G��V��3�&n��y�khu,s|z����Jj6�����OOJ��5�/��U+8+j/
O�r���k�s��O3��6w��k7�:�m�'bi�MD�;��<
:7u�����4��������1���y֛�p�޵�9wؙCt�N8�|m���7�t��'yX@b�-�O��▎�Kt	�9��eg���w=?�1�U�+�ο|���z~�xF<�D,20{i�ʑ\T��SXDa�V�Y\ȌJ����6"DUM�r�Z���5TK�A�ib9��n�<V�N&'����8b���O��gM�"�'U�ӫ�]z5|��D���NSm��b����9�eo��#ECl77C��t]E��.�5��YX�b[�2�Hr�`������?=��G.�%�W61��}68އ�.�yj�\B>�i�n�#�u/�q�j�}�a;{3���uL���-���̯C���t�a�6�����ޜ|��o��Eˈ������7P�q�So=;Ӕ(�/�lR@��60t�*Q�@�&���J/�D�tLOc�<Fow�:9eJ�D�#0mo���	Nv��LM�ҝ{�)O���2ֹ�b�*���x.�s/���Z�T<}�.����(I���}�;�z���$���+Z��z�	�T���Hạw�/���ނV�Brh�2�8��{5o9f_�!��;�5]��P��QX���W�)O՟���5�P��?su%D_���'*��w���O�&���<�=w��s}&���b͡�/�y��OWȝ���&[[=���=�&s>q�����!��uG�)ڷ�o�Zz�I;�,� �2��P��˄X��ʃ�YN�%�pGK=��6z��ͭ~�R9��.�Kr������UOcD�y�c6�C9X��hPѮ�[2����B����\���^�N�D�F5��A:����v�);�pjU���?��'�kk�č&�WI��]T�H�ǣޜ�A[��M��-�vf�CB�r�I�"�F��"dC;+Q+z�̄eKT�t�E$�`�C{JE��ɺ�(�*G������y[�S}�:glU��Wg(w;v�giD�v�\�Mi
."Y6�r�U�ݧ+��]\���1n��Cj+�sRCPB�/���op0$��70ƥ=Иq�t�]y�8�gu�r4,^6iQ[`�d�i��*s��MAR6��s��]�,��Xvj�1d+�s\�^qZìh���s�G7��ܪ��e��*fQ���j�G�S��_T���gL]C8�A���y�>�������;�"�D��++�a.�.mB��j�m��b��zW8��a���0q�U(����6���4��y��)rY]/X8�a��_a�Xh��y�$��R����:�+JAG���t�u�4�7{^��|���c�+2�7���z��dΕ�v��w4�mG�_�����|��&h��۶���ЙQ�pvՌ��y�7��7u��/lv�;����ht͕�M��fG�b�J�LE��Pkz��BoV���Rw;"������Q��嫚�K(ּ?Ē�w�a�4�b��,�r�yZ�s��3��+۸�nG���6WJ��ȥȅ�$�I$�*"fb&&U2,b
((���
�EFm���YLb
����cX,*�UX�i`�FF"�
�JU�Q�H*�AQ��V

"1R=��b*�Q���Y2�ER)5E �R"�QTPQb����Z"�� ��1UEb)FEu+-,�J*�PG)�Q@EB
*1\�E}�t���ޣ޽[���on�!�F�>��8I=�p<7�k�^��}�}{l ��l�}YN�s�
2K��с­�j���;��Xj�z�.�:���&M���ܘ�l�������Q�7�CC��>�A�ֽ���/I�7�p�U�j��:������M��+,�2r������9(�2W�+��i\TB���Ki-��b�s5����+��0�<5z�g���5(��LoR�;�bm} ��e��x���KƈhJ�ޣSr�ji�ʮ�I�Ty���J	&�.�e=�wo�vT�*���x;�W��b��,ɔ�g�ݙ�8<Z�[zƫ�)�#�Y}���7��fr�Q�:/F=�Y��7:�K7ޔ�xW!PQ�gue�������i�=b`��<! W[75GONՔT��u��k)H����]j�.Ņ1~ڙ�s�ސ\<�����s��a��q��,5�{�l c���)�m���}�ӿl�c$��p�~��m�u�n�Ԭ�o	Hd�V<�]Aˁ�e^� n��a.g&.�Tb�:�0�!u���՝� j�h�����v��5�c��h�����{#�s�P6���F�C��N��;�6*�ݮ�z�9&�2�Bߧ;�)�����,���Z���U�{O��y,�V������՞�70Hjq����"s�4�KE�.Rz3`f�vUɘ�g��»�@)�	��z٧u�y��q̶�%*1��#]���>�1�Qom���k]C���oz�!z*c�_G���贾�a`o�A���h4�k!���w��glE�l�]s6�]�iI�;1�*;��Е�?���qk�B��6w�m��n�c�8�vS%��*�+�Gu�����f��Z��Ryx��o&4?%��2qn��%�N+� r���Qq�����Z­���1��X�|�n��қ����ޝ48WI�Ⱅ�Nz,Z��GI�R�� nb����o&����l�I�bd�`�w���.�_g)/��
��7!5�ق�6l����
3|�~���v�v5��'M����{}�]Z��C/�8�����d+'J����4���r�2����gI%��Xc'�m�Bu�4��v�U�ɝ������q�o4I��/ t�O��'/�ۑ!F���� �c��&�1���p{j������h/v�Y�c���.��Ȝ��U�5�XR��סu�ay׎�d�n�S���'���L���D����҂괹a�V�� �}����G[LF�WW�v����ue��.�o��\�4����g���EL�Y�b�8��b��3L���N@5�-7�h��7��st�x�.3j-��]�"d�x9�p����i��L�~[�bC��=����:潊g���J�TEv��ʗ*�Ց"�ya�S��-섖�O��D���C]�c��7~�^��#X*�=?1���h�|�g9<�ר��Oط^�C*�E����#�Ow� e˹ε���]�E(δ`A���,�LUE۶jt�
*egD�E\�Cs�A���f:��E���f�Uup9m·Gw��x,ɳ�f�2�}D����]�$��tJ�K�貕N�=3Y����^eNYگL~�RY��hI��k�����aN���D��`�a���U6�ʴ��/�1��8��6�%HP<�s�L�LK��ŰѰk:���8�ԍx잝�輆�w�ѯY��ի�m����j�W�>��3��7"��Q�����K��~ж�x-哫�kۍ�I�陔�a�L��b�V�±�_l��u�w�k�Of�.�k�C���y>̲7Қ��[r]�xΣZ�r������Z��em�ά�=ү��,�������p�9.Œh�|����&�*\��c��<uF:�r2M%9���f�]딩��#bq���v���[�g�E�����aT��	l�^��ɭ����F��xI\U�^&��-�6�'9"B��A���o�&��5t�Z�ҩ/=0V�����Nf%b)���"i@:���,݋C�h��vÖ��;�ͽ$zD'C�t_w�N���[Z<���I���2LtU7�7x9ki��^U:��QLn���vh� �����S�D����2�g6�g�\s�C�-i����I���7Z���٣{�b���q��vK`28!�Ǫ�N�6�0d���΋�H6�&�������{�y۰��<�(�P��6��������+��ńQ�n��1�!C�A�eݼ�{FB��-������(�o6{���º��ȕ�L8�~��K[��+=��y��S�B:v/1��މ��v>�D0S v]�{gg6�����t��d�s5C2��;��jw9;�ՃY���U��lv��@L]�c��9G�>Y��1��y��]��]���Mmenֹvk��p��L�,� �=��AV�e���0E�lpY0��|-��ïC5��[��6-�����
��yUv�u[>������э�N�g��wGN����+GQ��Y����<N�
�d���к�x�f�y��;ڍI�����9n�s�I�z�Y�mi�73�7�Y:$�<s�k��}���ϋ�(}Mz���ǰ,�щ�>e�ߌQͭ��}+
�r㞯Z-U�g���|���)g�A�aҤ���٥�HՊ����k8�ݡ
��[PÑd]f�����໪ w����r�i�3^���F�ۛN�1�u��I˟M�萨}01iu��#b�c΍X�m9�1ug��?q(��zj�{��b��j��pv1ȯo���%��٣��6���s4wN�loظ�s�����Zޜ�ْr�^ot7�t���]vvt4�r�z��vÛ�ٮ�S��\�:��!b�i�T�|o�Q}d2n�<ɗ˯٣�tW+�SS3��3{	,S-V��ݍ���G)��t���"��,F�h}z#
O�M:`��Ⲝ��Ǒ�V�Y����V�|��O�ve\����"�poL.`J�2F���&\��k��E�<��l��xy��v&���5��Yņe곗U��ς'�7�����n�+U<$�#ΦM��±u����,-�W���u�pS�V+��_>������,l��+�:owEN�鶦,�`c�9O�L��#\��W[r���$d���{�kx����=5z:���E��I��6�i%B�2�N���IVN�ǝs��ël��Eŝ9r�Cȭ;�tϕ<����1`���(��.�r) ��\RI/���A�5u��Qb;���*���Rŀ��X���R�R�JU�iF
��"�2#dFE&(�1U����ADa�)rТ�DV�QU� *f�-�A�Fi�)V1��:m����ȟ��ت1�@�X��T�R�e0X��P�RP(
��R�+��&),UU`���)��
������35z��s]Ir�v��Zy�j��O���:a���9�ņٓ��V����Z�<��^&��R����x8>�u"����`.1J�ž���A�|y'�D�(�GU
��Y����VH[�^��E�^1���w5&�	Yz��o�Ǿ�N��� `h'��â6$1ה��Ç�Z��:�A�4�Y���;���Ұ�E{��E.404��/	��8+�]����ɹ�ˋ��1R�݂�;��hbb�P�� a<7����G���V���I弋���pV]��Wzuض����-4qc���D�ݽ'Bz�*��ٝN�qMX.���j�uɑ�#{QQ��.�,���L�L��ݓ��+V����*.�QT�"zu�(|׼6m�<i���&:�ª1�{]�T��I��K*�38cj�Zԣu�&چ�ws9$c��x��-ko��Z./z����]|\��p��uХ������d��5��$��\�Vq.�6�nm�0��6�'E$G�񎮐u���j��8�+�C��^�oL�az��ƺ��}g$m����k���Og'zH�\���qeq)�o$NBn�Y�DS5ݿu�����|al�"$Gg�En��d��d�0m�2pxt��d\\z0FO����e��X��� #2�Xn�5\"����v1�KT���C�+��ȅ�p�Dm�B��x�P<�����5/����j+z�q�4�wD����m�����~���z;�j֢�>}�&����A����.�;o3�}{��!}�.��M�e�lQ"��]���,O�f�$�7����"%d����x\t��U91B�~9>Oފ�zϷ�
u%bs>L�V�2���R�x̒m���{9��#���qA�F��>�P�z0.�"���A��Ǭƞ�m����7fgA�L5�"�Ơr�*Ѝ�v#oz��y����7�
.4��B�x���悓�[�9ȴ�A�p���뙯���[�C��3ز��a�pr���N���f����e���}���.�!&`���%�t�w}Q:霶,��G	��ޗO_)�}������	'g�ѯ�3����}r*�-�\O^�z5� �ĝV`^�=��,)+����5�1��ח٨f%�u�iu����E�̙��O9֥�֗�;�}�ɝ$�m8U�OT:1�;�-U�h��9�ʋ�aA����Pc��n��}˻�!w�X��z�@n�f�$p�å{�h��B��V9�@K�%&���~���x+ �/@���{���j濙�A��c)9#}����G�Iw�0���$ދ�s44bs�����+&�
$�;��f���S���aw�9�p��uS��ۅv�i���J��-��ŵ2;a߱���Ë�W}�.��њLl�O�b�w�{=�/��
��/�|��a��9ږΞ�9����%Ѧ�۬�m��X�ӫX�GMY�BJk������;}��ɍ������u)��]�.��e�[S�.C�+��BW/�!����f�"a�>B*OF�q��
��_����`��Pr�/���r��郢�S*rQ������#o����ʐ۬�$�Nעh�dy���j?��gse�3�T�`�B�̷@̘�foq��IY�Rܸ�,w3�^�+��s��qx�9�ɓb��k�8�u��;L��t>K��J�y�[3��e�\����ֶj�-��͈�<��[�0KH�"s{��z���8l�ۥF���0���G#����楻\�@�"8;=&F�Wuikͼ�q��tvQU�L�E�Zt�* �AjৄGt�E:ӫE�����]-��ӻwu��T��� �w*b�o[f��x�u����sC{��\૜�b���t������).E�*��f���d���owH0���e�f���>%�3O��Zޒ�|�O���D�"�M���s����3Y��n��s&g��>g2����VQ��=�<p���ݻ�_(F9H'NR�Zc_^ �(��p��#
��_X�h��q�b]۸}@äP*xt��]�sOn���E�N�oE���=���2X��c�	������$}FR���$b��n�#��ژ5������p�9ٹ�J}��6]�=��Gmd��ţ�ٛ���]�IȏD�����v���yQ�Fλlͭ��O�o:����1!؅r X�\�B(��s?&+\��_s���u��k/!�`Y��x{[��GJ�����Yh�7�k�W�}L��8���Fа*6l�G�)'�e�#1w�Z^oέ�-�G��WI�쒸��iLZ�i�XN�)��[����W8<��D�h�b��WmY�wmd�T]:뎄{<���o��ތ�~Yt�u�������Z�7ҍ�o&B��|���-`��gX��(nb�Vf��D]��9R9U��N�yTQ�c>��-�E����,��m�q���Jٹ���gt�H�@Fb9 A�uZ�1ݐ�r�θWd}lq�.!�n�>����+��Ux\V�po@n1��B�&i0�1�e��H0Ug��O L��,���+z/qٽ%��|,�a@�}W �	C��8�����:|��萢�\:u�5����{û��l6�����g쟼���?j�iUUU*���d@$�Y��DOb,�a �Y���TR�G�Y�qAvj��@�ê������L�Ǆ�uau�$��H�R�"AXZD� �!$g�n�3�e�e��
��Cd�Αm�F�"�%L2�����1�Imv��7�ЀI�RUm��kw�n:rݖ�܍p�\��i<�R��I�����A�6�sI�oAr�,�QD���[�߅ �a����w0�$ I�F�{�b���i��II3Ԑ	?2��O�QQi.�_��ѱ���|�'�x���\����O�w�NFӡ%Y����ď+X�rRR�4�"�G��]$b�s�
Fr�/�m5�+J=�1^�-��Zݫ�$��ފ7�+:��c���/U�I��Z���2T�I��XS��"& @ ���\I�p�@�IR���F�r�=�=�F�Pۭ?F�4@$�&D�J��,���C�1���a7=/yůJ���i�17Uf��M��~ƶ/�=ϰ-�����e�ٷ�T�H��KIMKÉ푵��>H�����0,��˅�MP�����[�˽�_q�*�NbO��ݠx�K�w̽�?�f����%IEh���J(�<[1M&��S��G-���#�"�R�	>ԟa�S�D�V�VG�^Icf	4{Jhc$mb�d�xH	22�J*��MB���d�|�l��$@��Rb���b�8��Rd~�Oa��i% ����	�H\�Z�?T#d;6r`�_��������C���kH����^�rOؤ����씞o�b}�Ʈ�����?��8"��A�M�,��vR�������sW}G�B%���F-��0�~� ���8c�¸��E�����"�0�Ii01�Vr����o5㧎�ڍ�x�mG�՞�f�hQ�/���J.K�+��}~�����FFn�5(��u[=~���i����n�ܡ ���#�F�>����mۖ*�
z�,��I��7k����(س>Y[��(�)�Gv��D��	?�T��^y�gi�G]yO[��i�s��'9:���)2L�Q��d��YI�T1�����{��Fت�������߭�_	����H�
!H}@