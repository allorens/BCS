BZh91AY&SYH{O=ڰ_�@qg���c� ����bO�         |���P�44k *I�D�R�Z�� VCDт��ĥ(�$�(5�@HMi)��
�[b�S@d��e*����j�/lJ�(�m�UM�SlֵH��R�զ�,ՄI�Z��"�Cfц���i�m("���QF�j���d4�U�Wl���y-�lUik�gk+R���U�ά�-V�k�Wc&��[�\�lҶ�i.�	*V��A�V����q��ކ�h�fm��������*���ծ��Fա*J8    ��_j'G[j����V���ڛ���e��f�]�.�!���A��� i��$R��Xm��M�ԍPUkjڭjG�  >����������l
w�yǪ�P)n�^��'����}(t:S�z� ==t�^�� [ާ�>�i�=�[����}7ڀT�wz{Uu�}��P�j����-��π  \��}R��
n:���cAZ5�����h>����������j�[�s��π�Ҽ����G׭�p����t�����������4��}|�򾞝��)*�mjZҨkR���� by�����L:�w���֔c��� zd/)�zS��r�}�πo�_g��y����ݨ[N�[燢}���� >����|�� S_>��|�_mJ�v}+Yh��imR��M5��   .�s��A[M^����Ҥ�g��w�>�hr�}��W�i����w�zol�D�^x��tQ����kA�z�7= ��[���=��@Җ�Ծ�����8۔iF����mj[Rm�o�  ���]��U�;烥|�t�x��}SM[m�3�O�}��@hW�����֒�7�m�Ͻ�7f��n�����>�iM�+�: yP��M�zһi�,q�@�]mo�-����TU4�����   ,�K��m�[h�=p{g]v��S���@һ�W ������A޼pMpZ��@N��={p ���$6�V�T��Ȫ�   ^ 4�9��9�� ��� [�u@s�0 :�zz�x� ���� u��p �]�t
�v��-�[L0�m[h6ś>   �����������(����nW�  .�p�n\С@�Lh�ӗ�x��o8p=t<�[k�:�E�Z�T5F��  ��F������ޗ�( -�=wU���c�u��z����[�q���/\z ���    �   a��2�)Bb��L�M2dS�R��CF�1A��ɠd��B��@4  �  T�U*� �    ������=�z��FL�	4�i�J@4�4��F�OHڙ>?7������tJ���k��`Tԩƚǳ9k2ϑw�������{�� I'���0	!�I$ �O�?� $���A�~����I�����A�$?�� 	$C������D $��3��>$?ń	$�����W�xX���!�������$=����"����r$9""C���Br0��D�"�'##9�7��ȁ�����d�@�@�e�999r$9D��NFIȐ�I�9��FNF���������`r2r<� r099�DF""C���؁���`r$9��#ؐ�`r r0ȇ#��Ȑ�Hr2n r09���G����ȁȁ���d�Hr09�DDD�@b#'#�����d�`r r r2r!b�F"NDDFOc��Ȑ�C"���DFNFMć#������c<��@�`r2��F"#�����Ñ$9D�""C�����d9��!Ȑ�Hr09�F"C�!����d9��"�d9=��D�DDDDF#'��'""C����999FNDDF#���'�D�ND�"C����ȁȇ#��d9����D�"C�FF$9���#$�d9'#�!Ȓp��#'#��Ȑ�`r r099q'"dIȁ���d�@�`r0=���DF�@�`r$9��#	ȁȐ�`j<��"C��Ȅ�2��#!��r&�I��r09D��!��r!9Ȑ�a9ND�� r!7�dc!��r$9�ND�"C�!�NF�!Ȅ��ND!FC���� 9 �0r Br0�9@���'"I����a=���# ���		���Ir$�r2B�!�`� B� ���FB�$!��I9�� "H�`F0r$�9H�!D �H�$FB#$�	�C�C�	�C��C�C�!!�� r$r$�99ȐD ��ID��"Cq��Ȓ@�d�r$�9r2CȄ���Hr$�9B��!D�B�	F�#n!$�Ir! dd$9B�ID�D��# C���I r0$9$20r0!9!'"�����d	�I!����@	���d����!	����I$5��!'#$��`9H����I r @�I r0Q�'"FH#$!Ȓ�!r2@�`r2���Br2�F��Ȑ�@�`r$�g"C�!��r0<����"C���a5F#'#���d�d�@�@�`r3��99r#���FC����������d�@��a999r2r {r r$99j'#���ȁ�Hr2�FC�!Ȅ�f�'#�!��Ȑ�d9�FC�!���K�FC�!���Hr2n!Ȅ�d209�NFC��Ȑ�d9�d�@�!��r$9<�!��+=����?{�9���P��ꄩȖ�:]�F�(�*d�+VP)��{����=��X��hU9tݷYPh�D+v������t�wyF9���@�؁�6���C�4XB9+p��wA�.�m٦���Uz�Q��\�t#��2��� 5]����e)"�����aQ��X���m-/,�ze՜0k���d��Vջ�IiV�3r,e�W65
� ���.�빷x�XCC.��N����o]ˣ[�,�mi ȷ!<A�j�|�c~}�u'X���=�;�k�5�����b���Y�2��8�c��y��Z�0�6wW���Q��飌.�0 ��r��.�����Z�&dy���Vn`@Z�aqn�%=�F@4�L�;��f��Cn	X%:��͐���M�]�w�i�EЏrLti�x��F�(1�ʂ���p�0JJ�a�D�ޛ��f�D����أ��Y�Hb<�驩V�%�q-uwc+u�g#o��5����*�ڭW�j�ʆ#�7����D�{���X0�S��cg&�3B���=���<m݋�l�i3K�PYz�
=�,i���a��@�0*b�P;v-�iMM�vJ��������[C6�E���̙V!��<�5��1x�Mf�ͱc wE�[��� �e9�p���Zf���a��7DR7L�Do1���FSU=�X��[��\z�lm]�{y�N��sUfnTR���*�y�X�hKa�x� ��#�!���)��ja��kPX5ZonB/��z��B��˽�
�B���!8�\P�d�Cs^V3��)(S7�]��q]�J!��B����Zy��*+����]C����
�Pm�.Z���UY��ٱ
� ���X�g0�S��/��f�;%O:��e��+��1{��ĝC��DܳOVCxT!�ypf-��,b�s��l8ʎ�Ʌ�9���J�U٤��3st��OD�+Y�6����V�{���Z!��l�`ɢ�^2���������%"MMG7��5�9�f�Z�\��`m����g_�V�C{zp�y�{�ؖMs7� '-����[ڹ��(�&;Ьb��̱�a<�S����Ԛ��ܱ�F[ӅK���)��J�s�h`%�?-���{a*�kM����YE�E`: 8(=��Yf�ȼge�f�f��XY7m���,�&9�p����'fP�Э[cjh�(�5Ȉ�w	��7V]n�t���tj܂�7c�.�-�o(]l'*�5�AOa��p�Wh��?��U&�M9�\�{Q��c2;������	Yfͧ�p������RH"���ё��N$֜�L��y,ݨ�@��V���5(�۴"eJp�LSx�L�H�VS����5�boMn���shd���c
����3�u�9څy0I�K���44V�j�U��6������W�lj�^�J�Xn�8e,[L[������A��V�jGGʵ�I�ń]�9�'WC^���)#*�M�ٽ1܈�c(�[�˲V�h���&��b��� ��j]m���,�c�L�t!!���74�^;~�'��09�Tjn��z7%Ժ�`�e�נ��"�.��j����C1�WVؚ"�7CW�����ma�����2��3���ҩʕ(�r�-�j��jܵ��ܐ�@؎��8u����N�df�6 \��3CDQ\j�2^�.k��kU�Iz�6>�ݰ��AA���Z��i�M#�9k�ʁ���Z��L��d���{F\��mn�R���ZqȂǐ�O+i).\˙��Nc��ܨC�24�U�`�
9h��!�� ��MlݠL4X�&�����F���,-�)ǻEB�&�j��2���*X\̻7�����U���A[*��I��N�w�X!�^�&��u�/�p�t*��S@�u� p��ї�C{%�{p�7�m��`ER�*d4q�.�ne��\��a�2K9z4dU��:6��TP��׉`���h�{4�ei@���<�1��1ȶA�[���IM�/wU�U!,�/U�n\��ãe6���MP�W�옜)6(�Z�[W�45����M�����+D���-鱆����,桮$�Spi�a���ݳ�ȤTl���S
�)0�@�;�rXݍ�((�G�a	ګ���K��m[�Jɔr���%Ce��Z�U�7;U�.�30���WBӬ��2�K=-V�ʶ�)+[�\��� �����{����2��S�N��$cL�WRhk5Ie�fx���m+"����52�JE�MVn-ڍIVe��:"�uAf�(��y���.���pRu�,�����[T���4��f��YL�v��E=���7��wtcn��F�3s-m�ވ[T3�u����8�a�b/^�ЃBs�W����w���΍��-��@�V��c%#��2� ����=���il�
,l�($�B�vfcoAoU�4j'*�	t1R׏�b�U;��� �^<��q�&�O2��b0Y�e�"���ڱ�95��bm���̲��G+p�6boa�a��޹ *ڇ�-�0�bسs�Wt�x��+cuf��oDc��؀���va���(:ʖ�j����6�*�Q�:[��-Z��dW��D�Kҥ���$,�����LX���V�eʷ��/r��l�m����JPm��X՝�����ZW�|����݄и�9n�+�jS�YZ��-���#��k7m㷌#��L��ia����r��+4�maZ�M�2Q���@W��΅Xֽ|�;����y�sIm�VP�9�E���wq]go�s�a�Væ��T�u7����<�)��{�Mڑ�VQ7�#��f顤�+(T����;wztU��7M$z�i�"�f�{��ejk#��W������4�7Rq���Z��e9ʦThGx�ǲ�M"�c�b�a��H��6�oa��l<�UI����@Y~��ܽ+6+���*�j�e k\(��!P��0��Q�� ?���3L�(������YB+f�U%���$�kRk�$y���ޠ���CNf�tq$S��X[(V�ཤ[�
��+3nK$%�3W���ףC{��əy6��7�51��j�Cf5T	!e�eU�M\�j^Э���՗�K���l�-���[h��jX�=Y$ةW�"LK3�B�����7��q\���U�l9N�ʔM�xI�E�l��ڵ�w)��٘�m�xt�q�]���.�� �q:E3xՌ�%��$t�2��Y�]f��wJ
Q��)D+L�tt��I���
d����sr�7-�(��ZZ༺ܚ��7ob�ѫN�@〈$Â���m��2���%g�ټ�L��Y.֠��صe�%eaG-Tqh��R�K^�n\�4�-c���<-�����Q����c��;�Q�V:[u2˒�ˍ��Z�а�����R�tCl^ӆ��"H�w���12їu���e�(��t^���6�V�W��^���+P���q��x�y�Vi[T�@8o-̞��sM�YrJ��X�dv�y	Y�x���4lk�Zѭ��[���cHݧy-ksH�˔��XE��7h�PI�+35{���a
Z�0�W������e	V�"�&�q3u���oPг�z�D�Թ�M�Z��[�/3MY8$Hv4�æ��M�o2�!��3M1NM;��փ�fYS0�jVԹV�7�(�n*rV��%JP�W����ʈ��U�s�ز�̳�M�0�U��D�e���MnH6��d8
����LG�5SQPf��,j�sk6�;2�m�R�dz�S�	�G ����a����Ӑe韓Q$�z�S5W�����ʼo:k�cO(ߖu-9�em����u��̭wy3��BBjX�YYteәj Õ�����'����T_�E�́�{o0��]�۴v���Bd���h��m�+*`��M���K��"6��[:�h�*ʺm<+$�9� ]����*�.,;6������� ���-�̦�B�Wa���Ye�X�f�&7i�BSGP��[�2;����ͽ��/%Y��[f���SQ#�Q��F���+4�mXv�Z�j��^#CgB�1�"����Ò���ڦ�$��%��(m�x��U��Ri�X0����lJ�G���y�To�cbBj����l�,%Y�̢��.�7V�,�y�N�	�8%(�%)��҃ܳ��Vn:���y5����ҿ&��m��U�u}��I��Y�b�� ;٫* 0J�9aZ1�Ʊ�\�CqU�Ka֘�œ�4�%������R���j#���uz�K%�f�ٛ�/7^R����/@��8�2�Xf,f����D���)�eYj��Q���B�NX;5��jL��s3]ژ�^����Cd*�lKPܨ$�F^Zz��  Ǐ4��u(�Q��ڧhff�.�-a���D����ѩ��i|)�C�N #��#j-V⫁YZ�Æ�+�)x7l��pXW�r�q�	c�gۭ܀�X�u{Xf�9hL�G�n���V��л��VZ��c��m�a��[�r�7Y��q�s/�!V"sfn��!�&_91��(�y@ݥ;2KI�-����m���EE�h8����Ց�,�T��bm▜��f-^:�u����q��V��ц�O`�C*�BE�8���޷�d�����̰ι.]��3�&-Jt7u#�E[���m�<�p4�vl0,;YEg��ne�*�F�xk�2�����n����T"n,�V%�Aұ6�����Y{fBԼ��Q-�)����Х@邘(�KUD!00��\]�o�il^I�h�t�ݹ	V�qn���d�������	Gle�#��n8�eV���E&ѧ4��͊B���ѡ���eh`��XkjΛ:yʢF�e����ƅ�`�]�P�����J#Oq�q����%�V���u����N�z�jՊ��������7F����%�r�
�e;��1I.�C� f��QjDm�Z�(�3**���;c��m-�j8������#DL�v0��$���=kB1RU����Em堷]+�&�������b!^ꗏ/��3R��O�������3Z��m���!b-�ŻCe��	��ںN6�,�<�E&�˦�k2a"n��f�;ǖ.xT��y���n)[an�!��0N�r��A:��Z�����;ZEfDn�܌̒,��w���t�ܦu��US)�� ��j�)a��[2�Z�(5e��n�7&�لSL�nġ�<u��L.nK�-i�4^�J�6HR�v�Yzsf�s^���k��.�h�C�����RR{���*A*
Y� �A�ZnÚ��IH�M[�P�$������-s0�zlZҤ����w�νb��LPW�S.6ẽ�!��u��Q[�N�+6Ƙ�J.��8�P��Ժ�e`:�Lt&��f^懢QG.Qe'��fc��������KPX�l���S�iY`͘���~j�.X/PT!��Hm�fGr]�e���hɕ{2l�iYl9XЃ´��x�m����K-���V��T	zq�V^^�@�Rۘ�m������Թ,,���o��_�n�¯55z����(e�t�Z[#$j�qTaaX�!�B��Ͳ'�-
�t�+�2��h��2�,���njOC2�#˹�(Z�łf��V��e�g2�񣉋�:Ւ�Vf#/sM@�{g^#����ǯ5c�X����&]�J�yS���/S�)�fn�؆�^5��⌊Cf��U֬���Ô�&a6���[܎�×smS��Ue�ά��
w��Nܹ*�7`��t�{L��J���wf���\�VU�Qb�B*'}��3N��N���m�ǻl��[�\�.�)[a���5B4��0Q[��"��ܻX��-��rb5 v��q��(��&av��T0,H�|��@ �rwK7����s{E���v�#][���
ýM�Ot*N<S�/lT0�x�
1U����z�A#5��cB�3v��r�E��2oKD
��z�ce$��8sb©466p�*�	��V�փ�mMq�1�R�����z�,Ǳ�. ��V�Zե���ܳ/b�M�U�,J
�Q� ���(0�r�M�j��ol�.fL�M	4cЛs-0U^+Gm>�K�o��K�)�v����(dZ*E�=]�"Mp=��,���n38T����"�*\�*�3c�*rq����~��$fV�.$V�K�l�	�#��-E}�5e J�$߷:��p0Y���,�.*#*�O���z��B97O)DH"�&�|�����4N���G���qPn�ޫ�	t��x�5�H%�]��ۀ�����hŸE��>�}7���O$���z��"�D]v�kV�[����q�2�:�Jl=�N��Nq,����2��hnD��h��)[���^��`�-���|p�*�g��(��}�o���N�ӑE�.�.�K�sF�xHJ�+.��x!�:d�g��Y�&5�Ӎ��V'v��cM��Jz�K.���t]!O�2�tҾ�"`|����]e�l��I�;��.��B$�t��t뗠�1� Ad��x�L� �	�ٹ�!9�ȴ ŕh�ء�'�^��+��x����o2D��C05��@f�JӮrh܁Q�	�{%V�mIR��3�ys���n$e�Ű]]�hy{F0�Xꋪei�=���2Y*Y&P��,�T�3�	wQ=���)�G��Ip��U _0�l�#*��8&�<+U
�"�:�L�2.���RC��ew@��F�ws9�_%_MG֣�R�yig��3�> ?]��`:�}����'��TM��B�Xq�E
�g�i�bǂ��"i�I6k[]�T��s9Y��{�2??�������?��P}~�|�GO_*��s�d�)�A7�}���s�)���o�t����^E#PS&)n���;�D�'�Ld�]���x��)y����]n�,�|�ߴ��Y$l�#���J���Ņb����t�3����6ewB�xb��%9��lj \��ɻ�HJs=�j��**���S��iCGk'�1L���$���2:�+��J7�V0K3^,�ޕ�N�o.�[ z��s���q���ˢ�|C٘�4��zm��Ε)m�#�ݪ	��m)֯S�����m��l�Uz�s�V�SxI�n�}M����2��{��F�X�f*���&ч�>TQXB��8��H4����¹��1^u��ͷ�[0H��%����jj�/(���}�/����IӗfI�n����á�z����7��7ia�j�t�h"F�u��uY��8n%]����[Ç'U�2��ͨ��i�1��Xu���:�wF��Ͱ��e�؛M���h���xh<�-`㹕.�]NN�dA~�V��[]1�]YPC[SK�`�����7ݹ�#j�a&�V���U�`KV�if ��w�wO�f��w[t�[wt�l�O��#�d��Z�&[ѝ�݌GDwu�n�]������m�9�I�T8���67�ɯCm$�ե�hyz�g��p�%��\&6�r���eI�I��5M�dM�Ac��ܢMS0R'�3k!T�a]`��}��5��O���h
:S�]q'V��(3��2��2��C(��?`k�S,�m�7�!z���=A�ֆ�Mp��Rv\�]À�jv��N2�j�lJ���ᮘ�^�XU\�y$�c"��"��i2t(.Baރ3k(�?l$R:.ͩ�PK7u�ُ�:�S���F95���HJ3*u/�7:-��cf����:|�E�.�G� �b5i��uP]8�)��,�.�������f��׼#˹4�5�	�5��z��q��
�:��V���ndY��������$Xʗ��v/���C����\�Fp�H!{�<7p*�.T�q�3t�k�*�՝���u�N9��kx`g)�oOi�S`��
I���<�z5*��2ٷ]��9�[wZ�w��⻅k���A��:��Z��$2G����-#Of3B��b�wt´�R��n� ��̶��a
�/"8ؖVΩ�=��]�o��Ol<�9��d��{G�u�x"�
Χ3��աΞ���-D����/�FEmu���oN��(؏���)C�4���,�3��Fh%�{�ٝA�ţ]��S��׷!�T�vr��`�@�m�N���/j֨�;�E�w ��~Vqk�%tV��h��q��cqs5q$ٝ{������S|��f���齨�g(��(GҞ4v��[�]�'8j2͚<������ͬ�����R.�ީxC�M�4﯆�F�X�ڧ(�%<O(kЗuB�nWL�ǧo�;{7
x���ٔ��Qs���oNgU�h�����IUjͽ�4[K����o5=�ZIx�"�v\6ʙ4{�����O�����l����tM]�lآ�k]7[MD8K]+������rvӧtPXM�uG�;c3w�Ȟ�N����x�hP��չ���[�G��ɴ��}v+s�#�S��;�:L�d`,#��]���H5�rZ�GSVP�u81�q�����7�ڒ�'��"c�hH-$��Lu��#c;Fb�e�G�0�0��9҇�����[�{V�۪��:V�9�uk��i�(Kje�^5���(�-�}���V�*eڴ7��Gc��&���!���0;Q� ��L�n+4Շ�f3Nn�/��J��-Y͉�������9�v͒�:Q3-Z����ݰ��ej��l�Kޤ;AV�3��T�m��V9�ca|)e'_Q��`0(�"�X����U貓5��
���͛MCH$�]:���д��8Fh�S&'Jk�ڏ:Z3�s��yp�WS�禱詛W{w[��p��%���iq�R��_l�[[�Ԓ�z����&��GQ��V3e
���B%���4��^7��I�4���e�m)�\��'x��6Kd�fpv!����s�p�\w{����U���р�K��K2&�=v�F�HUe-Z����2���S��2���*��N$���]xU�fe�K8��q��ju�0��]�d�j�K]fN�:���y�TYEц��<U���8g����M��P;
���m���u�$�f�[��+��Cj%L��M+�b��n�����`�v����zFi���[�oOR�(�'�&o����ʰnT�Y�5�C#��,��W2��.�I̶���{km5��M
��	.��KfEM]���˹�r�햞)nR�ۗu^��Ȉ�����[��϶+K��p��
��'\�����LWI��ݡu�c��U�È�S�[���OgtB�7}kA7n>���e�촭�����iBkN����f�/���#�˴w+��V��#.#I��Ƀ�����uMæ��R:"V*4� ɛG@�ڬ�Lnj�\2����Uڄ��=9�,�}j��XG>0ʾՌ��I�m��c+t���a�y��nH���c]!A�ݤ���� ҹ4zD]5���q]��u��z��_�\y�W���E�p���\?V���n<\�5vIy�(�W\9o*�x����D]\b����t�o�:����Y��js@���W6�rzQ�����}9�N*U��f�ue	
{\w9piZ`����f�`L��:$?��]�94�%:�1^���q��y�7�xUp�μjo1���8�Z���ys���Hh �e�k4���%�4�"�Cv��s�z�R��ղ,���t�Ǘ;�.4 �R�{�&t'V��%p�^v
x���u�X5[ǌ�-Mo4U��E�>�+�i��Ε-ECA�Y�z�i�IbQ+�Cp�H8E��r�W�6�'GeW��]�U�9\պ�ծ�Ƥ�h��l��lDYւ�eQܩ4��&�szGx�<�b�m	m�[S���wUb�Q�kf�c��]S�n��QGVJ�+xc��{J�+��2�=��fh��L�δel=o��}�GL�˷�(�5S#C'8�s����5�^B$>�6�0���b�G����S���xي���]:Ꝕ��ܻt)�-Z�{Z��TR��f�$k�\�P"��vHV��h��gJ�Jxڸ]iʆ_^ ��Dv��W�HE�X�/&�k�՚��i_J�V����Ln<c�K9E	9p�p�wYZ��4�-�E�C9������L�{G%hV�J�N�W�v��[vY��@M�ws&8I��8	�ShS�48�h��4z�`=r�:3MV�،��uZ�f]`8jA�U)��`�kkDA1i��,��XV�q�Ys����u�P׼��a��o0�޳���z���z�B�1��X��Vu�#G�|��Z�xMgio����qn�n1�#Pk\�"���
̪����ڼ�$���-a��kv/Ӗ�Wn؃W���[yeFg$49˭8櫴{��2��Vj�3�ˡ�֙�g�� ��~��8+,ҭ.�4=X}���U�ʁ�J�4I+T�ڈ��ݫ�cg.��"+�*��"�&�Rwi�bM����'U��9��&`�XT�[�,�N�]���Ca#��������[B��ZQw��s:SM����a�}��pC�F��bAR��^��ŽaVq�6B�]�3���h�J�oAy�f�wcI�ev8�H	\�# X�.AQ�B(�J{�ʸ�ږ�'k��aI{��`�V��]�t#89@������L;2렙9}�i��R��ˤ�ZDP�#7�w_�Am\ۅP}cvT��lU�g�w<�OA�K.��!�\�&ni��i|^�]"�u.�ĄsQ���d7O{�4e�0�9B^��9I��䜹n���%��퓚wM8+维�M����W�A�y�kk^*Z�}a��U��sT���vj�L��
&�SED`�e��:X�6p��j�7\��ep��UVfn�屩�k]�Iv���&�A�>�x��P	�ٻ�n��|pbҝ:y�@5�v�Sn��:�S�M_cS-��@k7��.�e��=�Q���	)�0os\�4�gԪ�FO�W�9�Zn7���1^�fB�WYb�,��4���J�tY����J7�Nk��1����r�V����r�r=�v�"�f��՝������QR۰����.���tĳ͂S��IkF�:܅�Nem� S2�X���SK����v]ܽ U�w���l�ӣ�G�B9	��K4��,�|��j�^j�SXo;���L�Der�����r��Km�6ix�.�lV��'N�1e!4�E�{pn�M�N�s�1p�趔����]��Cvq��+����F�zĺVt.�{d���Nm���~|��uPVԴ3��:��*����q�j����B�qf�-��8K��`�4Zb�˹�1�n�I��zV��ޅ2���f��f����y�!�Z���&{�i��Ӻ��[4�]�#���)��s52����μ��t�}-s�1��^b�.I�j�+F	���JSk)��M�`�����}�e��;7�9�B�D�7M�Vʁ����l�tv�k��7��h�:V����-���r�'p��jT�� 4�r��,�����7qs��3�Uջ`��̮��jIF����$ڡ�*��Xak��e5�U��v�oh&�kh��}\)f>��5V�6�j�t�݊�n�em��3��� o*I*l���V$W.�'Y
�7���:T0L�TL���{��f�Nm>sU���vl��Q���c[ڑ�/a3�������.G3����;���:oL�[{��ǁ��n�M��릆�-
Q[�����rs�Wj�g:t�e����s dmThW�2���D��^��ۘ��coC����Ì�N��+_���g�u����\����)W<+^#�K�݊����	���0up;{Ԕ�a�����9�n`S�edgxt���c�0<H1��2ޤ���T�x�5;<���5c�=ޥ�2P`�GJ�-&x�͘��][yi���e+��g1��a��AY5�%�8N;GuW�%hܸ�h�gT�̥Af��ʤn�4���;Il	�����^�e�M�.����n�{}�R�������ފ��ktT�rk���G�4lR�a��#�Gh�n�YΑ��f�v
����U3E]��wY���z �k�S'\]�Z��<*ol��1)��VJ���k���EH8�D��.�5n�%�P˦��*|�iY4��uG����Ԍf��Y�Un�k�w4D*!X4��	C��0����B��\w�%7��d�u����眤�!x�^G"�yt�`KU"@��[D跽�Z6�ѽ�eR��<T��7qE�u�n�s��[������V%�;��wT�,���pn�KF��6��cAc�x�(�mm_r�g_%�����"ԻtQ��˧w���ݼ�HLr����a�����6a�{y
�7τg���������ry���:��s^fp�� ^��vHho!��/=�@�b���l��=ݻ�ۅ3���Y�ܮ��P�T�2	�t)��X��`�5�[xA[���Dc{�7��=fe��$����5��VfP[\�pT��͓����7\�-h�T|���������	L�#���I]A��<D�;|u�h�Esc}���~����W_k�~�d��ّS��g*z"��g�C�Oa�V��I"�X.�c�k��O�����؏K�)��Ŕ�D�<eGv�n��HQ�:sTW��N���fz0���R9��̛�6^�<�g��n����P��4vK��͠��m���y0�;QEu{+l�{�N�-�^`���a6�HY]E��sqm�/���꓾�w�-J��;�z�o7���A�vi��G�k��$�Z{kY*壁�Ӊùˤ`ݥ��n�p˜	ɺ�.����׷����s��x:CV#�L��UU.�+�%:��w{����}:w��[� &���ɷ���*���??gz����s�r�]��.0����-�{t}ݡ�=|y�ԧ^E�o61���iX� �h�-Ή-��K�*�Si���k��N\��w��̊�&nu�V���B�3N%����yK���kW7n>��c��Rif���Om[M��9͈ �$m=�Dͭ0F�m�-�l;G^͎���bf(M���pKr岤GY��̴�Jx����M�9*°kc��޹R.�$VG涤!Dh3d�C!D$l���"q:���e�Հ�Sf�c_�c��}f��{�a��!�S˽kq(�l0	)"�J~�ی�a�\�C��<qLCNٖ��|�yi{���4s
�0\�0�%�/�浀&$�p(t�N?��~n�me�C)�0�T<�d���}]]�~>>=��z��h��(��DQ�̊�MQ�&b�[{f���g�+�k(Tt�����V���x̶.�p�f��q���/�u�H��e���n��Q���k����mY�����մ���:��e��e�i%��:z`����q~9I� v'vŹ6�f44Q�GL�>\Rj�������-��ޯ�1۵f�d��k��x�|ˎj�W,4�k����1��V<���ٻ�;dZ��;�λι�kn8�4��M���|o��9�&�+�.���HI	�?O�����	 @��~�?_��!�o�߳���~�$��������}#�(�����;��}1@� �C%s/[��Ԣu��ٮ�j��Я&qQ��jwu`�.�e¡��H���v1���c-�,�����r[�G��9��哮��vU�!l�ݕ�����0�z�Է��ז�M2:����ጋ"�����t��Hd8�;�{R[���sW)�H����G��Ķ�^����t�ԍ؃g�ruSǪ<���e c��F��w�r�K�yB��Kk���p-E�Z�!K��,{��R�h.�}r�:]k�p/X�u��8��	��ͫ�ڹt�g$�|�5��&)�;2�E!ҷp�Eyؒ;r"�T7�ⶪ�������ClT�铡x�P:��a��A^���q�9u�VG�����ӽ#��"���AjI�&��N�$�{��l�%��*�$���]��	�х�H�sx��p�r��|ֺ̇-٫7��b7ނ���uf��Ǝ��%�y>`�`%�&({��	_����-��ί�-X�t)�Y5��0<�Ń����\�Q���j�3f�^�SR� T\���):��Uv�w�$F�(�����2|�ۿ5H�IA憊��v5u��_J�f�]�՘9����@JZ*a�@��q��Z���3E�#��Q%������ �j�4B�C�y�����q%9��=-*Ѥp�&;�V5Z�}O+�k�{�fO&NNOg�������������������������vvY���e�vvv3�������������������w�����ʒ��p���3n�}G�9^�i�qԮ!�P��O%�.-�m�ΰ�����NV���koG$�u#J��C�DQ=���&�]�oB�uc��8x���6���ћ[B�sc�.���v�B/�9�x:��ղ��LD����`ۼ��ٮ���j��у������8*��Qj�0ʦHu,��o,�,b���Q�H̆�>��٥�5������Ψ� web�C�U�WZOv�s���l�za�>���W�*�uI�]�V�>ΈQ�٣H�G���^�z<�U�����Q�v�é12�V���]3
;HF�͆�u�YZ̺
�c=�Kg��#�7Sn]l�[j�7n�$��	�z"˹o�ݼ��:�_v���;,�9��ا)J�qm���*��sVSc�޵�	��9�YF��h��Y,�v�	����|3yV��x��an�=�}�ld+�pi4����f��	�/kN��V����z*<{�m��x�Nt�\*ԙ�r��n���MQ˗}�zd=3o@�em���}5_s0��[�1��e,�ZNL�uk3/s:��Q�7
�j����dJgz�I������kyB�lKM0�5!��Y;��u��}Yv5ۉ����3xsR<��Ë/4�%�L:�B���a1�!�5{��9\�sy�7.�<�V�ǗӸ�O���������}���{����������vvvvvvvvvrv3����,���쳳��������vvvvvvvvw��^;�Z�泤LԺ���j��P�/�<����w�k�|�+ZXj^��2�C.��;܋Se&��E�eF7Ks��X�<���y�W�^���3�7o.�ފY�u`(� ��8�=��$w�{�0�*k"+y!��͘��-��4�M?��u#��G*��td7VЏ�g���mčb&��Vj�!�ʗ� B��z�VzdMW&o/9>3C�.ʤ���#�nd�4h�
ң_6�׶�n�t';K.�c7��J9Z�]�ͫoӇY9uݳzT�r�F�����!���1t�[9��ZK���0֏u�w{�X<٧.���צP%�#��X�trV.U��;��P��A�o��&����HY�XPָ�z	�9z$R��^j;�þR�l�bf��4�w�V��������$U=�A3�9��Z��GK��鹩p�e[˥I�@��*5���ɷn�[�I�3�Y��f�;̚���W3����w��!���k�V�H��7�0�5d�n�LSQV���p��6^��+��7;4���t,f0��=�ʾ�q�I��&�M�5���wO^m��tWx#��,֘+���v�"&g'4I�6>˧Q<�{W��������#E+6�jNan��ui5��H�t��KZV��ͩ&]!�Ts���+*�������{}��u{���w��S����������������;;;,������̝�������������������L�f�����y	�1��څ�������gY�����8V𕳥�NK��xn��i��-7,�\�@i��}ojM�\1U���ښz�/��q�C��㼆�6݄;a��qd����r��p�-=�su��d�l�	X�kyj�!K�×9V�4^��V���gvO'7��5Ɖ<u�[깪�b.�[���;E����6�P��]3�_d�;���C��:���&-�rF-tX(]�5�Ia���=�;���59(�����¤�dv��Ȇ@�(�W���� ��3��p��y����t�1�C(O�t/4�W6���X��K���zd�X�eC�Lتn���>���b�w�4AW�u��r+���N�؛�ǧ"ܿS7,�|��Ä<��y6�V��(\����ܥX�].@�ԣ�X�*4^H�a�7/u���q�P�ؖ]�,��c4�4Noup�v�Q������B��)3OI�ނ�.���,�Pv�_0.,M�4w^w?Y�u��i{����RO^pSg����c�C��[r�b��$t�⛷f�rpi~Lq3��{
7G!q�l�2�,s��S�v�`�ﷂ����%�ɥ:�m����қ�1r�\�etz�Fzp�Z���d�Oe�cw!��������{}��g����{�gggggg'gc;;;;;;,����;;;,��gggggf�ggggg�����������{=��w�X�].�f�+�U��q	$����\iq5�0T�Ϸf�'1C�
ݮ���+���ݕ��'T#hg]R�q$�uV�j�힜�E��KV���ً��t*�q��[�	X���},^Ɓ�v���y[v���8��I��q9�V`ޚz*Vb:�d��Kgov�o�j��eT�#�l�0�4{ewI�̼�!X�Xj6A��4JF`�#tQ.�g#u��e� ^�gkr�1���2 �tk�{����e����P��M@��S�y�ꭃ4���� Lb�F�ŔI]�t�K(��FzP���G�Bv��M+_K�vqm��{\0ժ,�XL���aE�a�� �jb�ZW)�ԡ�
]9�͋:��.XK��T��,Lf��ͪ�j� e�?��3e_G:;A�9n�9A�˽�=�^�P�۵�E��l{�0�"v�T$�����y�72�b�g���G�]�1/��g�b�io2������ɩ=���v�F%�����w�R]@Q�	u���9ǭ����MaC���6X�:p�pm�F��b�X哝o��g��-E�]X'M��I�t��4�-k���]y3�TJ�Ɋ
�y�*�,�z�����K��Q�Y�3wEf9V�M��D(�Sy���y�}��o�{;;;;2vvvvvvnvvvY����������gggf�L�;;;;;;<���������{����w�������*s�J���4w��K���aa�ʕ4�v��T��7�Z�w�a^�T�7���cb8�-���a�q)�T��5�l�qq6�4��#���EYuیJ��k���k�)α��>܃�a��oq�P��Go�lif�`f[]S2u�k4�vի���{����]��a7����6�"����;O���Jp�b��ͭ&\Y�{}�WJ�fb��E�6ko�q�����x&�x�`�ʕm K7�׹vKҤ͗-��4V��[ݗwt/�۽.����x��^d$�̩X�1v�צ�]�4�Q��h�j��5����c;�7gw���Ê!���K޵�Z{��g5��t7*N�D3v�Qq���
F]�ͺ�Df@��v3�fAVУ���yܘx�k�Nt��W �BSvl�)U�3+-���U����Oڰ���X�Lø�y+�En��R�Qh	M���wc�1����m���s-�>�f�t+�J��(��o�.����*��ٗ��Q1��1�|_[�j�9�k��\��+d����Wλ�]R�ip�Sܒ�p^�c�ޱ3�hT�2��#@�F���Y��L�F�cT(R�tAY,��[.�{Wyˑ4&!��,����Y�Fj<�2%ø[�M����h����y�{=��w�����{��^����������������ٹ����̝�2Y������ٹ��ٓ�����������/b��*��Q{K�,���'�%�W:���Ж�2�@m�3+ c
��}�]�q���}��k��X=m`X�S�e)�zK�]ֳ��9��~V�HzWgC���n�^�lN���j��X<|��=yfȾ�����F��̖��b�cp�T���+�TO�D�ҧj��pF�˒e��`�nu�Y��w�.�K�I���iV��c�Ķ�:�Yy}2�Ǜ�O(m���]�]@>ޫU+����v�����1K�O�m��ctZ�Sh+4huiZ��k����Q0�R9Vm�36﷓yUEZ�z76h���4�+DUيKB����C!/�!�q3z-us�\'H�*�{ !����3]8qɹH�0Y����[mN�jr�kr�� 2#�,�q��]ḟh�}%�wV��u�2<���B<niW��w=$`Q\�M��p�ײ���H�Ϋr���pY����_H�̜mL�?u�l��;�NI�w��#��ˣ�ܺ�z�܃��+���9���]�2L�`�#�t��s1�d���2C☏�q<�q}��G��+��٠��j���i�P���3��#��-��^�ņ�a2ԼG!��9%N81u��m3��=2)�\��4�W]Pk�#v9M�k���d����MaR��%���;B��H�\����%��|�K�K��G�E�Y��*��n��&�'g�s��٩������������������������vvvYٓ'fFvvvvvvvv{;;,�������������w|��9a���[�P�yݓC+�$e���bU��6��a`D�0��#j�v�H	(�e�S6U��a+(��=)�����$��{:���"Me�<����-�fW z_;��</���9�7����.�S�HR_I� o=/0�dWmi���&f��,�f�s(��tm�>��G���@�4��=���{ju��z�ri�}B�&NG��6��)k�[�8�:= ����h4�c̆�4�O�l��a@8�0��w��Ji����K�|������gxn�+A�I�d�wQ��k2�8����[���]�5�R�����ʗQ����gP��jU2V'A f��of�YTW.�5GƠʕ�s*2'o�i�̹����`�HmSw�������[���	�bf3�Q�ݜ&��-����UЇW�)��<p���x�aJ���[�Wy�a���2��.�_>���	��Y����|�<�l�mOQ�|^قj��ٱ�Ӆn�ֳ�GS��3X�!O���v�O;J��3Z����lm��k�	�=5'Ln��@R�(��5�Ӛwn��W��
0��e]��c��+����[q�^�ˢp�v�K�S�&ĝ����c{5
<�/��o�E��e�q��6�yK�Y�H��#V�	�}�ڰ:nt����Y�\	��uܕ���3-���l��2���+M2�����k��s��&��zӖc��&aO�vv�z
����T�����wI�����z{}���w�����ggggf�ggfN������'gggf�gggfL�2t����������������������xxm/Q窸nv���ؠ �G�����[�A2	��N�������=}���_4��nrՙ]��|�S�{)����mݍ
��[[AH-D�>Qu�R�-S
�.;�7֙��*-�ʲ֓����U��<�#�ժ��֖�I������u�XF�m�TѲ�|+ �
#x����Vrӎ������mk���%�_r}M�zg��G>���L�1B+�EC	�7v���C����������Ud`c-��a�?KÙF��qr"���B`�'��Z���63"S�/���&�o`w�k�6�)��#�7.�.�s�l*<�ƘѴ���g7J,���Y8:Ҳ:�Pf.�gi�*b����h��F���1ˈ��@�t(n�OK[\�r�	+P�ŹĻ��-��<ԼzO�b��h8(0/���$�)�4�7]�u����b��u:ۙg�͑/��wd�\�v��7�����ZE�ŭ�^��ih�����������F]��u�-�V]ܛ3*䣨H膴Yd�:V;煸����!�R�a쭩�ʹ��N�祱x�PeZ����׌�yKɲ��Qa9|��mv5wkvU�7�`���ݭd7p`�W]�R�m��V�(�S0Qɍ,�G/ ޓ�5]P�=���<'��UܬFHU�T�Pr�/�m�MM�lm��T��rm)��]��7�b���(��KZ��\Ĺ,��Xٗr�qr��l�x2��4�.z�d[�O2����5P��Wۙ���f����ƛa�]Fvn�,0���[u.\�7q�9�Z*o-w�/A˸ ��Ult{�Ү���k��+�s��j���)�(e�	��W��4�i�K���d���"�kr!a�ѹJϟ�A������a��\��B0ة	T��͜��N�Y@���6��n�g��kU�%�K)�;]�;�:\b��ǜt�H����W'�vT�Zw:͝8WT�����%�=���\���uN��n�U֬!�0�����/��Þov�JU���U Sܪ���4ڏ+��͑J�m��lmB��t3�A�;�j�H��м���g G���n�!˸P�<'h���;:�˒��&M����SX���r�Εz���E,�F���U�G2�i;�xk�[��K�<�������<637�.De���`����7e���w:�1�&��]F"�VMŪ\�{�4��r��;9�hn�yI���8p]e�d�ӣr���&0:�`�ns�&�K]am��:�{�S��� ��]���x��܎(�
����޸�4�i�Z�Y��u%�Gקl�mIF\�w�_U��T�
4�X�Ɋ�=SD㒧�;��B� lG��!�w�+yS���L�h�@����>� }�������������������/����=.��VܰFD���C ��`�ȄH�?�X�玌tQ֬t#L�n�8eӖђ0`�0Yo�%�0I���)G���"�@�V�Hx�h+4,�b��b"R1��_�B����A�v�j���τ[��-W������L�P�l�/�Rs-A}fQ���ڷ��ڎ洯��u֥+��Q��	���m�Z��O�yM�R�ff��Dz�T����]8���,��vJ��XH���h�<��pc5�v��<l��O��%^����ni��Cl��z���t���f��E��{{�_q�<�O�-NSu�݂�e��^i�]�*��5��h���N��d$��f�,�t�4K�5Ҙqnʬߋ����I��N�?#í�uvX�d���c"L��FSͿ(�KB��ݳ�ZJ
ݖa�ю�<�7�fz�M1�]5�u��ս�(A,���1��8�c)=�4}`��T�Z��jગ�J1^���_Kg,�x��.�9�)��u�%`F�(�$'iZ�)wϘ����܍�-��A}Bg����%JXuM=��	<s�����B��dk���2
v$���������qR��&T8N����k���-�绦��Ύ>�o�t#�,�6�qn�r�+��w]�x�l����%w*���5�n��v�NZR䂄t�^h{���m���c�-�A3;�s��P��8���]��S1|�a���iMb��ηo#��t��*�NH�GbN>��.�ԝ� �Ճ2�6.)
m~I�b"�FSPA�Z,�b@ے8cP����TȂ8�m�C�(8TF("�ѨCI0h�R0��(��m6!"0B0@R8�D�,B�m�፯�(���ܖ�(B�����ȎQ&&a��h�U"�T�MxS��B����Z�El8&&�a0�lH�	��&!�B\�r �&��bi�2 �"L���J��&U~!Q�J,�Z֜tZ4�����\˃=1=�H�;�e`�Z"����eQ�U-Ab�[��6�ǩT�)mDA�m��Ԩ�[,ɩٹ��b��"��cn2����TcF(T������-m���e��g�ss�jo�`��A�BbVAb73'��Շ���b"���[�X��&&X�2{=����b�ʓ��U�u����Z �@�R�ҶЩS�b���(�k+�6hɖ�Y���nl�m-H�E-n8ņ_fB��j2���aXx��*VQW�sWUq�bbX������rr{6DkF)P�bcm�-!U���j9s!�ח�Lj
����x��X�れL�k��Ƌ�2UM+��M�Of�(,��s����V¢3,��k[m����.�V凗F���G�&&�ⵑR�e�mF���\lТ��e���m*�UV�u�b��F�'g����)�
ͳ/�]h,��],��QƗXb V�r�Df�8E���fd锉�ے{C1�mGBX#6aY��I��$1
_3"cf��1^�u��ˢһ��Wlɹ�s����
��(�6�Z´��K#X�2#[�h�JYhT,���T�[*ZS����IQ��T�+��X����fZ���kX�0̵(�mpW�Z�cZK���(������������D]2W-ƈ��W�*��*�M�ҥ�y�.�kY��0J�V�e�:�ʹk1�fh���m3&W���}N�;�Ή��~�v��|5�\}_��	�%r<�S�/:X�0���r�syo-j�i9k��&�LꜨ�X�������Y�U���--rwH�+x�3&��6ײ^t��{��e2�Aׄ�Y<-Z���^��!r��D?��X�m>x��,�������}bwc�#�O��+��\�����'�;���x^�~��@��l��Cx���Ȇn��3[Tz�|.i�,7������Ѻ����p��s�߅�}z�Hw�ׂw�t�1ƙ��31{��������Zg�hpō��u����r�w�{�7���<=�>w2tt�c�>������+����bu�}������QY�UyeD<ټ�޸2�~y<u���l��Ѧ���Ѿ=����
0##~~��m�d}<#�f{��7�g����]+�[��:������h^�=������H�OK����8o��5f|��Z�})V罇�����=�9Th_xP�C�����x�o�NA���mߚ�O�s�g��Zd���WQ�B�|B�ί��Ŀz;�����u��F���
޼��B��&$�ښ�B�l�N�zĥ�]p_���9��x_Q	7[V4(���ǲC�v�[yvl�Q.|j�gąqa��y�E$�jS-�Ǯ��)Iz��S*��yM��N��ۥ�{J�Q�
��ٹ��ogj�7 ��7U<�<�{E;�
{��,]�]�>����_1��3�o��Կe[՞u9��0�4> �\`�ޑl�Va��/y�vjEw�#�i	�W���*3��:����������|�<� ��O������d�ap.�\~$�P�����ʪ!}IV��B]���zT��Å�=ܚ�=�n.@�4.��GI��'���xd�==��g�P�ѝu�7D���dȋ����!̌�h�OGW`������Lz���xpᴀ6Uz�<�*�<!��K�ue�=ܾ�V��W�EW����U�ݗދ�÷Z^�=�x�>���\ߪ��K0�c�@�`W9�޲{^K���5���fh�rtc��zz{)b��:�6����xQ�m�Cz=X�'6j\�h���u���zx3����$�&WR��e��6+�;�bޓ�.�k��ks^
�f�E���lf}z�kB�.���Dt�#��UVH��#7'F	Y[B�+���iap���	]?�~�Aw��}�g3�S�0t�t�^�`�t^%�w�Q��(����aA��ۼwm�}���yܛ�V	��_�WEG+>^_?Q�ϼ@��籩)������Е5;Ԯ�s�26�3*��WmЊ�>��B��伇�{�/KϷ��O7����β��(ǝT�>۠�,)b�w�s��}�u���n���x���G �?'%��Զ��/�ض�԰_�}~_�?{,>���<���[���[���OJ]��A���5<*{��x���q`��wş�FK[�Bצ�XF�zu��P�;�ٳ�1�B�����^�c��}$�A��E0�1*�������m}f������|mOo��`�J�]������l��(lm[�����\/��iwl���e������޼�	��N@��=!�t�;��f�;�}����/}	V++b�Tz�Tn]Q$u��Xfc�@��q��jz��h�O�9k��������e}���x>�[������,���G7�q��0�/��4�V�\iG�\!:&�Ry����yZ]�:b���3�+6�/�$]/��A��q����ʇ�7O,�*96��v�A�32�oUԺ��g'0�niFQ�c���k��U=r�~7�_[��w\�{����b{������J2*'k���M�}<Ar� �wO����$г�I�k���;�9�<�i���V�f����F�[܃�dW�]��x��������i&�<Om<f�j6����+ճ�e_4�Axp޲ذX�&1:J���}<������ɺ�n��S͵;ҼYب!��=��r{'�����s9�~˗����y��VY�-*����w��'J��dXç´�<��d���y��W�9��on�i���(��q��~�8䙶m�y��K�Ѽ�I�8`T��&*s��\ɖ��!��Uxz�q�p�f���3M�ym&��a��	�!����xߥ����������߸zM߯��b-O>��z���o�/}{�;}��Q��烾�5x��۽���b�o4\�lǬ�W:%�>���WH;,w�a���f�ڴY^̜Qߝ�� #�b��k�n�5�G���kʧX��ȫ5}����o��B�fj^65d�7��n�WH+����M�j��L;PI��,�D��KÍ� E7��D�;�|�;oY��Di�D�\.V��Y����ӹ����G�]%��V��=�Hw� ML#�_f����6� J�.��w>��3���S����g#�<0_G���M����v^�ٌ��Tڝ6\����J{(����?h����ZX�U�uFW%�N"O�^~B!��O^��ʕo��1#c�TȺF|5x{ &Ȑ{�
�:����X�	n>�w����"v�~��}B��Ͻ�_m���&���z�	�i�m�a�[�����7����o.#���J����<n�ǻ\�����o�Eݏ����'4=�*�h�%D �hz�\���xj�o�R��D7�/�z��k��?$}��.�OВ������8��=��=��|�Cc�����q�c ��j{�8C�̲�L���a���6޼:�9:�6�[vHx�8['+�x����� Q���'��ɑgi�s�B������9A��[� >�HR.c{��M�����F��)�3�G�<����j<������'e�Y�Wl�KH�9�\Y��X��j�U�t�����ê�^��!ˮ���7��쾋�T��҆�Aئ̝�; ��2GK�D779�.[������������پp���H}1ׅ.�R-7n�Iݑ�m�����v|��N��	=/��w�߹�M�)OJw��Ga�볬_�`}#�;��=F=B;�{��:�<��͝mp�f��������������ͪa�!m���?zJ�ΎG]�{�NMnCgwo%U��	0T��C�t+�����]Ó�wUN��t��zJ{�_O
w3�)��t@�o�OôgPO��kJ�+z�W�����x��oࠖ꿂�9PW�GdD7G 4i�]�U{�K���pO3�\b�b�S�^n-IXK��/�B�7��,VVMt��^:V5�u��>ֽ�&W�����/~���/xjxL����W�ѵ����.M�����{҆��#�Vv�{���G8=������_^f���j�ưW�ք�cg���M^��G��ܸ�C�m�8�=P���Ei�H+�#\��@~ň�t�t�	͚6�;��KiEW�h�h� NZe�Q3�ݢ�}�R��m�c�t1�f��X2��Fp�G:�6���;�6�U|E�ʽ�y��*8�;���0�,�w��{n�	��D��Ȳ.�s��b^ Oh�w}:tN�I�n�P}��6���g:��:��{��ܸ�Pvcm+>�`Z�e��`�]��!�Y�&�kg�t�u����{=��N�2mǮaj�z��N���i�����SɞO~z�N8��t2�3o;���R4�;�}���`�
���ٯ՟gϣ�����&/Jg��5-w�����{�2R�����u��'�Ǎ��[���O����$���e@g����r�p�7ᮝ���>	�ހG�˾�{E�:oWۛ�.U��¦��pL�Z���soFx�/�P\��(/F,.�<�1�us�P{�e]{�k�\�*��驫�ע��<�����:"u�8���L��`v����e^��Ǧw�nGv����Plf�<4n `��9��=��d�g�Q��GF�2k�Ş���vw�h��J�o7*�ԫ�u�Y��Py��om���12k����չ�I�-T2��N�������1c��DBeMp<#t^V��OG�v��R��"q���7l�7۪��o�׌���As�4������g3����<<�{%�n�@� �Y��m�dԏv���2{�)9�߶������o`Zj��.�n���{�6�_�h��C���;����"&\��{�b.��7�/tM��W����DN�s ��a]���zg�Z��z䥙j�S<'@�~�	�o�	紣��٦h������[���^>�WǼ���o�9gR���A=g���6o=�Fj�%�շ4`�|�����W���T*����c�xX}�-��ƽ��=F����Fm���l����,������}c@>�#>��bL��C�������{}8�U�����xG׎�/Wi����n�����bu˱�5���fM�KC������+��C�rvM�֝��j�A���ú7���Y��o�9j^݂��e��d�J�]�,��t&(Ⱥ�PJ�k~4�
0<m�嗬�՜[�q㆝n�P"�G��������j�z6����H젊T�����'[����*9\��܊5�wH��A��ʹˎ:��op����h߀)�L�:r�Dl����n3�WIwM��	�[�f�*�?K��3��E��:�������`��]=]^O/�D��?z�ַ�ůL�u�L|ܽ�+�����.��A?�hW��	�=O���ǽ<���Y��lX.u��}�D�
��D��|����g�E8:B���d�1#��O��Tٟ@7 e�zOpb�ʾ�#UX}i�S���{W�f���A�{a�p-��g�ڀI�����h��uqy~�P��|�ʡ�Ey�-������3�^W�)Gݤ���=�X�^E?��U�ٮ����3r�[���I��C=�;�0!\%���g��~�ؽ|)t�L�3�O�d��ws�O��'��= �����uÄ��{Ύw��W}�����{a��ʪ	�X�!{��=�"����GX�i�dXto����,���~�cC�`��s�&}����ȯt�zm�%���Y�M�B�y���":6B�v�J;���-Z	.�%��D3wW8I]�#gϑ��$�Aj]�c��@�F��M��{�(7���Jv��!�
&��]�6 �b;v�-�,�/)^,sx�e�4ǽ)�/;��gTq�ޕL$w|;4����m���g�����}�S_	4o�-ٵ"��Lo+��/aK+s{���#$�X������x�b�޹9�_�^B�xx���<x�l�����c�Y�s^��tY�T��7���O{&��ʻ/O�\�o��<O�b���j��=,1�K��/��\̜�/G|�L-����v�k�f����bzL���DEH�M����6��S�S����g׾5PGfc�<�9ź$������6��Lk�,r���ܓU��(�
$�W�ߦ��h�dyr ���̃�ni��F���=���%��gxT��/���4�g���6�o���E-�2�~�D��@k���Cn��f�D�3jޤ���`v?w�z'`���(?�����mt�����e-}�-yn��9�5�I�N��]��Lz*[�9�� �/������=\�L�a����h��>�ot(�L�����ɘ꺕nhSZ�7�2&O>ڨC���i�oL�����Iq�Y!-���]��5�b�\{ԼΎM��DLd��͗z�U,U�^�Ucr$�\n�E|�=NH�j,��3���w�#pg �.����R��٦+��m�z����m��M�N\Դ6mÝ;TO,����+]�Uo���sD��ױ�W�u�4�]Sw�r?u�e70.V�5,U9{���7]1����ԣ�POo[@;��ݜTc{]We�\�Z�1��K�F��ɲl��걌wLa+Q���}8*��c��o����{�)Gr��mբ��{���.<A��:`�봞�����t:�'p���[�pP@�G��Tt#Y@���,�{������\��Y\jt2������⣉9Hު=���FTˮ�H����	�n�ʠd�V~����#%�v���f�E�(��HaK!*�����O�d!��7��f�ط����Y�GH�V����E����\\F`�U�K;Ε'���ۮB�K�$�^<�3mMY;����SA�b7}R_F._��ԫ�j�f��Mw��[������U��L�J�:��!�]��֩���+S).��t�ƚ�tԷ���w���&�8j_D�[���&Il��B�;�5]<ЕȰ�57c��*�*k;85Qv��6��o�f��,}�,p���fh�,�N�a��&X=j���-�ۛ��M�7\��纾\d���쭤_��E��|1dGۥJ�?	r7$r��?��~��G.�����f�����ސ�h)68ngud�.�52��-
�3k�V���M�2�@�U&��4�Yrd6�Z�r�׼��S%QG/*�k8d��M�g=+��*�GJmՆ��=�[P�r[��"�"�ؽ��i���|���W���8�g�T;f�0E*74f���z�>���hS��sʲ'��t���}��-�m1���B%7-kb�]Up�T��wź��5�\j�΃&朢�L;,�Ƕ0i�}�F�B-��luY��Q[�[�P�a��JX�q�w@���Γ��X]��4�۴��7����m�E�ŝ7�A¯i��v�d˦��R˷��Nv���j-/J9V64s��J����VMx&.�R�LO$��u��{��o8�v=u(�j9N��ֺ�5:�sɗJ�MG�����ouի��X�rv�A�X(�f���U�|I�q�6Λ�jcv3lԚ��������ѷi<���g�W;s+�H8��2̚�UT{�H$���]��_Rޔy�����"���LI77�����n^�ی�3��.���0iSK
�e��m�ݗ:��:�޾�8�r5n�&d��z����R���[�e�n1/u�Z�s�q�JsN=���\�y������f�g!�����Uj��ə�m)�#�%˙E��1��[㉈T���L��7n��`��f�j�SW-���q�3'��sss�sJ��Qb�ZQ,D�ƍo�M@�Y�T֭�ӿ3���%R����s<t
�4e�a�52d�rnnx���m���R��*��X��<@�c<��x���b�.�f/)T|M�y599776�wX�m���D�0*QEˬ���F#�B����1�֙jT<r.[�2v{;<��mU�]Z����
ֶڢ
Z�+
²�����7B��2d����/�\��-�5TTAOT��ժU��U+Aģ�,�s!�L�pS�m��>5q-fNNM�&��m�K�����\�G)U�fMd��`�h*�Mr�񢕖ҤTm�GY���9=���������v�EST�J�X*��E����2���M:�w�0�._CzʅJ�L|�0,������nU�d�����Z0��8��(�YY�3�2i2�D��{����TV:ˊ�+-lMRV""*���H劊�fŃ�.`(�����z��9��(��n���M�z�LA����rc
��v�3�u�J�l�4���Ihѡ�G���k��f|*�����������?�a�~�D�����3���'�G��~o@kbs��ph9S>Y]kz��౥�[� !�p*^�������n�P�2}���K(!^FK �M<��"nY�$@8���:��-�-�Y�h�id�� fz�g�G����#���m�z@A�xnN'	��9��*�Ֆ{*��4�qI4f�'��V� c�I�$��-ԥ6O=�Mz�%6)ڮ���jsZ�3��t4�/t�l������J�}^�D~�t��*�վ;�
/͕�%��G�/+ ���X�RW[rh�p���P�8�bY7�XH�2�U�i�=����{`��E=�Ǥ*$��8źa�T�q�=kxD`��,0p�|��w-H�l�j�=e��e�i�m�e]��e�0i+���/��Bz��=�?���y!�=*���b-9@����sxs�_N�N�.O]�Y����b�A���A��D�ٸ��x��.ݎ[��g�okl��|@w��$�jƳa
�'���f�wCpʦ<�έy!��`�yҒ9��_̈��vvZ�6�i�9N���/}�ѡ�9X|~)T)�t��;;6e�헕vm�u�T�dg��$t	"����ɦbv�gg5>U�]*ح�@��i⽄��u]&����S9�l�W��Z��H��f��S�3�˿�;m�(󫐾Az�	���AN�XzI����ƙl��x����6�Y���շ�kT>����P%�s��,(!��~n�vd�zdN�
��Sw�#Z�)�n�.��y���|�Q�ʠ=�d'4o���H2�F?��<���������s�4�5+�z�Y�`�`�MO�mP���q�:�d.��<�����\�p�G$[@^���t�/�_Y����GVKVo
�kn/��ޡ��y��a��aşïI�i/�ܵø}F�^�P!,�kyg��߬���Ec�����7ꁌ�J�m����"4q�(�v-�c�� o���]�K6n�V�R~�&{��M��A��m��$�������]�W��f�y�=��}��oal��� �^;�fq�n���`1�2�1�=Ų9*����ˠ1�/��܆ᒪ�f����� �ɫ�d��5g�6m�{ [:y�S�z���m�ȇ���0~O� ��)v[�=':hs��x�\�0Bp1��a	0��K+�����_�)�ڀ�����#�C�u*�96�/w�pmb�;>'�Di�NJ�?F8�^S��ׅ+UE�5*�i�m�e�B�Q�;bb���Z��P#{�)�)u�aǛw��XP�ޡ���+�l�
L@��ݏ�Gq������,!]����MHv�Nu�j�w1�:!Y���k�3�����|5�S�/VDqm�|�/���vA���zw�������xS����HDx��ݢ�2���>�6��35"|K����ΛB4r9�����l��ҙ7�xN�F��UE?���BYN�P��꽲;��`��[B��oHN5�r���!�>��K���T�g�`��{���&���@F����+��w�㠴�
�6^��m'+v�Y��Q�<�4;��v|"�QK�1�E��<�p��tk�]6�:��i�ǣ��1`J���)-�í;-1C�O�frk�\~��]Q�=��
;I�PY'�Z�f��)� 4��G�&�q[�� �* [�B�"q;�
GL�1��1����)ͪ4,�s=�.�D�y����E�����( ����P�D�G�-__��&L�`9��ͳ�~V3����t����<��B�s	�{�툕Ch&"��g�}d��yXwe��<�A~j���0�P̲}�~��Z����_�@�}�ӭWъ_4ow[��������.1~c������0sް�|&k���`u@n�6�wz��XZ�ʯi.֭ޮ�����]ۭ��ު� �{k��l�8��7�!ެ=�O��N��`�j-�R�B��7���전t��Lgk������=�Ҍڥ{�b�S��J���/�2��Y���Q�5쬳�Of��Î`��*�Y1�3�Kh��s���e�2�ow�W1�m4#�S�H����N�,��틵��s�O�S
��x������iD[*�Dہhlg	��Yv� u:����f9+/��Y�%V�����c�"�3!'� �� ����M4���MC�.�E3���d��a�y�����0C�p�q)�_	T&������b��I�RN'�y��F7�������yş;N��:)��3�|���>��g[�	>O�T�e@Z4��?eP�r�ORS��w��S��8�s�y��	l��v�6-�'\�0s�mF��$�m�V�U�>Teڳ�?�]��.��2��"�7��(��r�IPp�$��w*��O>��Czp��YQ5��74H���ޘ���-���px�E���L��^�KνL+���@ipy���Gܞo7�氳�9�]�r����s��Ȥ�&ʥY�ʖ�C��NZ�}DD��=�D̝�QW�;��;��K0�E�La�n�;�� ��v�~�Z~`/�AcAt�|�=�8�t�g��a���l��П������CM�"��XИ�꺤�-�Ǳ�h%Q��Z��3*|;���f�$l�\�g�eX��ߖ�Z�#�o�{,I;�A��Y~�^��t��w(ڗ���#�vݼTz��C[i�����1��sdY��l���x�8]����z�HFA������Q"i�&�w�*�}���ǲ��S��y������of���Pnݡ����h~.���<�O�N�G�(w`��4ت�[+�X��= .v�݋}_���ڛ�gw|��?�۩��2L��Bn�����	�SS�Һ��Ze�����˚�q�X�r���O�*��>3��������,��<<���p� D�~�lP�ˉ$�7�qys���f�f���-��lc�\,�F���?S�����?5��I����|������2.�����C��p�zKy5�^�����v���z	z��� ��яꘊ�L=�	Rȉ�lʛJ'(>f޺:+�PνBKhN[>��?�|�>0I�>�#�W��9A
�2aÞ8��:ٻ)]R̈́:�]Yu�p&�@��SČZZP4O�'-Չ�G<�� [O�%L�gd�n�K�T��%�tV+oe���S�6��>oN���n����Z��@)^l�|`�	ȯrRu���&1�)iޖ��й����C&�iM'���Qs^=zޭਕIp�(�h'"\3ա>]3�=�6.�3�å
	�S�!8���? ��`�F�]�u�5��t�[c���נ�ߏ~��w˜٣����N���p,�z?�ܓ�u�����֔���y�k��:�q>���a?"�rڟ�!����F�Y��q, �Õ�.�-7�F��MI�亝�1�{Q�pn�碒3 � ��Ww;�7�K�x���g���$��\J 6dp��\��}4�ɰ�Jr���Q�����nm�.D5f�2ۂ�oy��C�X�.�c�|�ߘ*�.��4��"����(���	���=uv�׫�z�qן#����f5��~�hLpn�q�%������;#�\�ٳ���Y��_;S�J�l�v�K�pϝ��M0���5zm���;���?O@�B�QkZ���ב�7+O<fVc�����렕$3S%�����'�my�=�>}�n������J(�r܄a�k�	����<�)O�T�y��Ļ�l�X�~C���e���:u<�/�v48N�2#"�Зf�c+6�K��5�"OL�_g�V}��*��~�57�t*Qy��wt�^f.�����M"3�mO����T#k�ԓ�~e�4���a�nm��_KLE�$���c��C��v{��@�	���-�c1��ڟ4k�q�5�r@��]ش`ïo8����5>_��H|�w�K?��͂%�!�E�.��̠ӭ�o]T���i)�CMb���|�i���B���Y��U�&�`��O{�>�t���D'm�o�Qk;��B}��/����PUW�X�c;\L_M.k���t]
�M���/SF�\���|e�6���ا�\"rs���.���AF���]�6v��<R��i���V`^�6����U�3�!H7�
������N]��2֙�>hI����P���2��ک�==��"D�;+�[�Wso�Ѽ�ƙY���x� C�VJE�z͛e��L����@�`d�	|��ŵC��vQ!�N����f��/F��7@[I�A���\-@�%t�8u�5{* �sW���ٹ]�^Եed�;���/X�os�(�3U�g��9��2-����1���F�7�� ��[Qm�����l���a˥��:��4 ����� $�^��BA�M�^~��$��2�i<X	���~��#j�]�$��;�ply!��v_��r�����#^?����/z]���J�)�OEGp��7}�СT�xcez�H�u��x��/@:�n<����
1�C���`��[�e��&*I�輫У�28�+U+^���X�74_Aqm���8���O䤰z���Y�c��{Aqs�N�ĥ� ����u�zz|'*�>k�$��W�ܢ�`� ����0��1D� �����d�.�=<����oS�R�qL� 	h/��P�~s'_<ٜUl(NU������N�0�*@��V��V�r���i h=ݝ�gu��R|{sljU�9:���a92���;�p���]�;,�W���A��?pU�ǖ�S*�_e<͚�%sk��)�X���8���������3�#$J�|U�Tm�%������>��#Ōb��������׾}�u�-��1i����T�����ذR��#'^�*	{k��'8�'42^y�UN������^ǰ�lx0�(|@@���?d��4�wߟ�{����`m����5���3w�#�|]��i�n`$�֘��h�dx<o�&��~��7�,�fǷ���ۨS�Μ�x���j�	tIp+�a۱�# O����y~W�~�c��$����yO�7!�v�;�l��a�����q�����!h��#�t�!��Z&;�T��WsՔ=�H)�:g�b�.}���gpq�V�^��<�.��V�cĤ^�d\
+$!^�\�c�:k��t޵�
z�klĆv^�v=�_��!b5�h�A�S\��cGEH�A�!c��A�,��~J�8}�p�TE�t��b�V��|?#���t�C� S<|#�pL|�#�G|�1�T�K���^�����o�^V���»��#�ن}~��ῇ�ݨ�S�tj�#�}U��Ŀ�h�S�Y��*�����2�=��ZO\~��g��L��i�B�F���>��3�V��'��C)��3�^&����ǅWy\T�^*FG�Ut��	�4�\C$}����M�cY�Z(���b�0��̾�o��s%�V$��R�����3|�U���,H^�C�ǭA����gF:��{uw�]nd�,�*�T�nD�p�ʎ�j}�i>�N�П�#1�b1�C����(t:[��Ё��4=<fJu��K"� n�e^(�o
��W8���O����͗u�[F"4�#[��լ%�L�!�����'y�(�o�R���0ʼ����:���^$�~
��`�Х+'���E�2y�����z`&��O_Jw��]O�Z�5�,it��75�C�l���j�p�|%.}`��a�`C��~�������˪X�7��!�y1�$wT�ozf_J�l��M]򝝿ywha�
d�gS��>a7K���ß�x��y���.A��� ����e�+��A(��/t�Ү�o=0~Ο�~� �z���** @�;j;_8ؼ���yڻR������I��(��xϧ�^�Ժ��z싆m���D"뛙�slS̍���=S�78�d�l�{)?[���q�<��e�q����Ű��3���wC�e���ڨ]�)W,ӯ�8"�C�?��4�)��wPn����v��%�qhHb\uK^/�͌��g����l��k1��]��Y�>�@���ʿE�׎�����H�{�h�)d�0�t��ύ�XFR�f�w��Z��NnP��Z��74�L2�f<A��:���#�t�A��ڊ�;�g/vR����{�{�4f���Ĥ1�,���"�6b{a���ɝ��ܠ��օrB���t^���[�jۗ7�]c��{Û�y��?"�� �o0�w�*�C.�Á�h��8��yˇ01AT�����w��S��lJ��\��͜р�Ax���#xLܮu媵�j�Õ���8�i�g�H�x��f-��Xt^|##���8��O9�#�5v��Cw3cs�x�#�&Pd֔O.{i>�)��*e6��i?�s
>�9� ��ᰭ�au��ezx��{@k6�	��d��Fi��P�]�sz��=���On�s�!�敄I��޼l������BW��4'��y�?D�@'.�BrB�ȣ)��G\�O$��6-���<�ه[�Ԇǟe�)� �f�re�7���-�a�&R~"����E����P��|�Y���,9��������c�L>��~��<5z<�o���0v??�|������V�w���UR�|�^BOZ���r1-�|���h��|��ב��\����_/5�Z�MgcV����*�xkt=��~���W�I�ҏ��ǿ�a���}\�hh�/6��>վ�.h��.����SuzU�n>�f{!?G8��at%����\{a�9���H��<=���ƛ%ޱc��X�� �ˌ����#���1���;��m#�0���ƫ8����yr ی��T<�F��P������	bi����X����z\a�z�U-�4�uRǏQKbV�}�(XUs&Π�UeL��(����;Gi*���X���c���B��KEf����oh���c{��.ʧ�Yy�7B\�3�S�:�mM�sq��3����V���8q{C��*�#o$��d��W�0V_>mw�Շ�|����Ϙ�{A��׎�X�9d���QKV�sۈu��;�GJ���q6`U�.��;��R���onu�*���W!ɔ<i��q@���۝�����2Ŵ���םT�n����v���ե�8p�`�J����',��7��չ@���JN��cA+v��ۡ��^�k{M&�A��pq�VF�r�v&�Xk;j���c�$�dJ�m-jr�x���w�rS^���U3m�WO�P��}��̝���ʱ���<bW]��3(��ꨝo��y��ͱ��D�-vI/�<��N㏫++Q�¬NE�ے�mM0V�mc�yc��5;2�`�S*�B�ai.��X�P����Ey�]�7P�;f��e���Z�br�k}���DR���7u�tq��4����©�CMM�P��\���(�壳ݶ.u����K�Kw|�o ����ɽ����6��.D�*�����T�й��MZrd����uڒ��*M<)��S&Y��j�Xe���q�Z�Q��E�ڏ��)�9���C�m�޽��[���z��ԟ(z�m$�z�����;D�c�����A:�>1͝��o[ӝ}��0��uzK�X�/f��s�|S;���*�!��P�%Kp� #읫��p�ܱ6������������
˙��G�1g�Gi��9s�$�^�54&��\�f��Y�I��V�~1;b��\+�
��;0MC�x0�z��}bV�7/����=h�;��*����W[G#�j	hd��׵b5;oM���9=He��ذ�������"h�`�xoo���rA�杻��tn"8�Â�\��5!|��Ƌ����v�v_�5�H�϶��boi{� �Zļ
�����m�D����Э.�M�Tٗ+�gm;�3X}���eN��mZb�n썹ð2)��QJ(h���.���
O6oT���
s�8�e�,+�y�v���m�B?�K�����>�w.������;�������(l����"��g��ت�N��7 �0����}]v,Z��\t�ɻw��\�wC/����҂JGƟ���Α�<�f�تs��:���ٮ=k2Rb�A}��ێem뒞�ۼng-)��a��� ��d��I���9.󩭲����%9:����� \��a��1�R���SZ�ȨY%�
m"����D�Y(��XL�R殾�]��2̥DX�a�E^�QX:�	1�_cb�R��CL��a`*��s��s`mXTyLE��jj����+E��e��KK�`kE3%u
�Fjy9977;b�.�U��̸�,Ę�jX	sM3�"j��i�6�����ٸ|���+rۘ�j,EDC�\�
�Lʶ��L��Т���B�f�''�slM��>K��]fR��1��\Io��<M5<������fb�\pr�������jm-����Y�GT��5���qAĨ�8��s[�Q�_�lh�R�N,ɹ�ɹ�;�ˑ
���*�X���2��L��[C�������͇7��Qrҳ2ܳMq��AJ��nR���sYd�:t��B�'����6��]ۖ�W2�epL���m�Ql+�+̎9J��1%�it�.R�q�eT���iDX�����ꈕ�Į$m��r�9,�3�P�jc0�4��t��10�e(��nL���Z2عJ��4��y^+[ �7�M�a�دo:'�>!�U�M��v!����v25��R�br#`�ٹ���2��nS}Q��_r=Y$ӇXS��$J���b�2�	V�f�5fycM��א�{�|3ƹ���g7��?T>�b1��F$�db�W�������|��g�{9�.7j��no*Ρ_�&�����X�o�1��K�1�e�ǣӝ&�|������'b�`�����é�\2����fYa�@tyS������>;^=�l*�.� �ٮm�˞���
���>˔mFEV�X�3�J�z����S�m(ճ�*{Y_�0�ٴ_���3E�ka�Q����|�U����Rv�B��L%���Q�O)�1�.#bVgn�b�����ϲ�e��g�c�B�̽�}���"��S�ڜd
0��Xg��zMV��@���o��uMG�0L!���M]>��[s��^�R��`���A�QY=��g�6m�cW�T��a~��)5lO�)����!�g;�y���
p1P5�0]'Ƴ�B�֠Kuc=�|jʀ.���^��M	��V���PfV8"q�C�{�|d�^������:�dJ *��Ji��П"3:�E�D�͌���)܏�o
p=?����|���i�C�SsP~��=��N�Z}��3+7c_�\��*�\]�Ͱ��"��>g�Q�K.���g� \M�����z��#�;���V\ypHM�Ѥ^��s��A��Kj%���/n�TV�����c���w��}ً��卢�q���kn����pG��H�fc��
��Ѽ�T��В묢%G�;�:���սw��������}����	�F$b1�c��� i^�a	���͍�@,��Ȥ�\h��.͔�������r�L�Rҗ�uM���n�?O!lW�M;H9S����E���#4�;Ͼw±:R|���Z���܊�mSW;�]7lSH�A�_E<��Fg_O��;'�C~��y*9�v����q��}������0�lQ���7Bv���D@,y�^u�I�E�q]��N�Z��3*u�j�Ʈ� ��P�ff6{y'hԨ�(S��r2;��E@���������J�)�zl��e��E�ު\d�e
`����G6s�P�A	�4{GAi
Dv���k��,5�9*wj�j"q����u-*�Æ��(v����>=��{�yå�PQa��	��c"�]1�9;1'�v�f�;l�nAR�¼�Iza��������G�9�W��m+���<�Ź��Ʃ����
+3^0MoL���Xݦa���7�.����L4�l�����6�M�����������,*��<����T�A����L�ɌvAʸhDך�e�o�S���_��t�����s���&أ�ӑ>S�#�Eʺ�ڼYкvw\�ܙcV�#!F�Jr=��j��;-%��_gn��9�/�J���s�Rl��Y��Fʭ!❙{W.a�����"y�e9��z����<�������C�0�H1��B1��# u��;���g���{	4ƻ��E>��{�[���qa�@Mж��HX��A���'��Y�9��.3�Ռ��yAM4��k���ϤJ��[9�L� ���:�ի�LZÔ$��0�::'q���8<T��d���n
�v�Z�����/Ý��',� ��s5;�F� r�x3Z:y[/9���Ύ2��&���w�ɼz��	���0�L����h���i��i=��D0�$s�8���g��h���,�u���uc,�]I�?C����/Z����8k+�7wKz����^�L;].Cu�Y}E�GdQt��뤞s��L��P�^1��OM�Oj�W��i�3:���_}�7��� 1���ǯ�>��N���5ʣ�?3��9��r+��W��hwpd:�L?5���Ba33��=P9niDkx.�uI`Z���vJ�/��w�=B��1UٸL3�]�Z�r���ܣ��.�RpTx���y�Ok#�بL��L8�ʴI�Jj����Z��N�NKԹ��ԍ��`�>����|�"qy�i��da��ۘ���6+���{���]�;�=؝Y�|�9P��f>�3�nk��D��jZ�Bq��e��Jv+�yaq�F/-�dJ��ͨ�3�n(xV��W�ڄv���_3C:����-WBQRq��טn&ͧFŵ,��,7]�H�qχ�~��2� � 1$�BA�Ox���%��&j��5M��ҔĲ��˾���ZW�~0f�'��`��0J<��?����USUweoaס�Or�dv�m��%9	��qh�8�x�yb���MT,��64��Տ���L�#ԗXTCX]�&�T��4���/k;H��H޸�'��CT�!�$���e�ӥn����_��5�6~��C���Z��{m�Q`��G>v�P֑���P������ɶ�]�S?fTzP����P^K���f�j�1a��H���DC��><�/Oa����sv5����i����h.����8�7
�#����z�=[��6*���IsZW@��ۻ�����XBLW���/��ɨZSI�*��E��M<���
MÛ�e��uUCݽ�9��ԅ$;]n@�>�U�A�.8�2N�D�3�Z�G[�P�t�՘`�a�g��Ŏ�@�؞q��`ew��2��s��G��%��S*(�ki�ݺ�r�,�3v�*e��u�뀠[9P͸&82��`��K��oQ��L�r�';�F�K�+
N����`�B�n��پ��+��=Su:"[�X��C�i���d�k}"��h��EO&�t"0�#�
n�Pu�R��.��vS���:���N?j�=��V�Z�\������U�"�M�f�&����W����t�:���������=׸i�.Y������c!$#@c$� A� =3d=�z��Bj*�$0i���m|;h�M^�\
|�>������r!1�`�3��Qɫ9��|XRW�CN��MR�&gV�˥�e���	}E�w.�a ��?BD�>�F=3�^���O!E��Em�S/�'�q��*���y�^���������8���>���=��F����E�4�V<�������
���T�n��k��I��b2m�T{<�de��cD�
d��{�߫�ni�GPS��ǖ@�j�]t	�ڄk�1L���z}[~�\�6R�!�2������ĥ���!�(PVWզ�+m/^�d�"��G{�b�pl23L(qh�����U/d��~̃�8�ޯ�����+	����$q���َ?�z�c�'���^ї��J����D��S*����.�L1j�\OC�<#�כx46D��2�y�����< �˥�_����z&��Xv����}���n^VNP��K�9~t�&a������S�<]�N�0#�F0P��#��͔��t�6���a�l�J��t&�ӕ�X؝ �G ��,�A�v���*o�E0�����-�͌%��Ϯ�1e�ě����|t:�	DyfX���,�_o	F��z��V������wu�d#�t0�h��m�i���my0U�ө�_�c�S�['����[]at�:�m�ɰ.r��k4��*��ʚo�8"Q*���[�9מ�?BI?H��$�@���@bF2I� >�}�߹��^��P���0��c����	���zO�`�ըƼWV3�1��݊踂\SV5'�C1��[W�3�.a��P����m��ǐ_4�.�>�q�1I��4)m�����V7M�O���n0֍���z�(�g�H����&FP�I�n9��; Qnk�L���9��[�w�9t�n5&�͋�N.��~�-�Ʒ�H���C$`�!��s�-�4�u�y�K{A�1��ڌ�����c�E'+��}~��;�<0���cH�!?E�\;Y*�:�M�v�B�t��K�W�᫶����q�d]axX�J���A����F���ԩ?�S�m��g����`S��C�d^�;�ؕ"M4�Ux�yj�r�͂���v���L��QM;��n����'\��>d�q7'�y�U�k�͹��,�%����f�V�};��H�?\5W��B�š�v�Rs��ԁ
�9
��n;�[7�Z�sŝ��a�J׊��v��~�y��UU��g�H�����a.�������1��/4Oٷ>#����2�X���%\�h;��v�7�m&wEv>;;x'���W'��$�na�Ŷ�mܭ!\�մ�i��i������ñ�vEa�N-3����W�J,��\����p|�=dRz�Q��xo$nc�U�nt)��尕͐C�ל�w�g�c  c!#@�����I t�|�>}�Jl��ͷ���6��r��/x��<�K�k�:X5��D&l��' �V���h�W͊s����f��#Qa\bK��ݏ@q�tE1>��/>��@�#Z۬��c$��9�Q{�8)�榯N���ݢCy�K7�^mhT(4��ꖠdE���<7lS����ݭ��8�#�V���}o�p�5fF4��\��;:K���d-%^kØqM���}�|:�h�A#�׏߲;jj�0Hny2Ϫ�������g8�^g��K�ߴ|e�����<;����V�Gz��B��S$���@d��J��K��[��no-oKLGS;3h<ؑ���ѡI�J�^=�~��V����xk�#0����O:�T��S��n��܈Z�C/U�\�lBmbS�*Kc�z��M�B�r�R� ��$ۼ�BF�n���Mή�ղ���0X�*}���u��K"�E2�i0�����7�,>d�vW�!i}@�T�j�n�@Azİ����A��9���O�ƍ\F)�])�D�w�����k��&�eS��)�X����~Ԇ��tzM�`���`o�,�a��7׆��Mљ����T�]����q��dS��o)��!��ʖ(W%/��'�H�f�������C!W��,uވ�4$���lX��NGf��ne��z�Of��Q�����H`bI#I b! 1 @��Ͽ=���~�[������O�T_�̐�.�#��O_O�a��㾋OhZ�2��]|��v�>�"?��fj4����pZm���wZH�Y�m�����_Z�g��-f2�3�	�ff,\8^]
FK(��n�i��	e ����#̂�Y�إ�!L�2�UD�����=�b�r�`���S�=K�JyTφk��]A�@@�����׼�6үg��L�
��~*9��C�}��n��uc���|d��j��g�/ldؾv
=T�;�>��k���uy��g1����y;.5�T�K�������9{�F/jR���gB1E�\��Z��N����x�)���/l�n�m���ӽ�- �jɇ�L�$���n��
"%k�!�P����Vѣg�T=j������7hz=�}M���s�\[j��ݮ�02\.ak˶�`÷�}y��<��Hǖx#�Z|�
>���&=���y�>��++7����f�L�ô�G �4T��ݵU��)I\��o	I�{R�|	1{�D����U�e!Dv�a>�:r<~���B�E�b�GoQИK]��2:��Ƒ��]��L��>�V��N�k��0�PXC/C�'Gm�Lj�я��-ڼ��FBm���h���CA��QH+��!���4�b��d�$��P&X5wf�����#� �@��$���b#�[�~}�߿{���q��4@��l�7���	M�8���D���N01�zǂ��Ƅ�l��֩
>�̓�L�CU��^kۧ�洇SOE�X�pH_o �W.�g=��y� �����D˷Pj�54��t>���k�Rps�s�������y�?Bd����YN��z4��1�U���n}G���;��/�ǟ5)K4Ð_j�):K��4i'��N��;�CS�8Xه�:�j�Q`Z��.Լ�AÃx�\m�v%�jŦ)�&�A��
c#K��	�^��-?,<�i��7��,3���69�O��pQ�"Aqp�V�&�D�bf'������S�-u}�(�.y�2z*;�����:XEC�c;C`v�;.�ݙ�tT��Iul��2%?WT�n~�[�oIN*�O��)���B��R%L��¥���oqV���A�!i����GT�Y��д�g��1̵�>��Y�*�;
w���̇j��.�`�:�Oz\6z}"8"S;c"���;�H��׳�'�t����X��&]7�2"�]\�cu7>9s+n��x�<]͋1��fSW(�#k��)y�䲸��
�@D����v�5EU�RҾ���w#ΰ��h1�j�t�#�LL�H�����&3���;l�{�r�Ct��{���#k<���>o4r���D�01�@bHA��$���b���>M��3*3 8-�=ywV�sZ�$Z>d��
-���7J�C�vU�V�h�t�M�G0˻��͵;[d/.�M�j����pt/E��o��:��.�;H�q���ܵ3���I�<LR��X�FѝUӳ�1{�oA.qRi�T6��sbzR���	C��E�o��6�nW�xpT���8�7�˛ic�q��1b�d
2of�W@�t�FTC5��[k�0�gs��`{	��X��� g�{���a����OBO�ga��C+����*fi���-�1P�\3!�+E�~A�6'��p��jC`=J}��z����M1Q������m,FN����7Z���}nb��:��r�-震-�Pf<�U	;c�P�_��6��bs�q��f^'�7[��$��h%S��40ɶ7#U�µ�"��&H8��t4rT2��W��aC~N����>*M|� )����c����4j���b©���r�l��[��v^��#�}n!�n��n�YS��S"�=�4�����=4^��s瀑�<=}��ѹ��j��8!C��*۩�1�W�&m-��e���D��2�z�s9ddy���;�x��֕�[�5t�&4�-�)�b掏�����*i�T�Q6����b�찍U�+D��5f��B�T�sW7�]*����ӆ�<�sd�#0�����X��۳.�yݴ�b&VAȬD�8���9W��Cy_J�M�9��iB*�ʝ
��ܶ��S��ل�\��P�hf���/p�ێ���R�3�7�*U�,��L����HS\�;���j�!�����YT:�h��2�Txc���Zs�?�I����Ӫ&u����D�}�8�#na�y�n�1�{(����ï9�(J0��)Sګ�S�q�[�L �A��Z@1��<@��x�V�1��=�O���� n�l^���k2b��O��^a޷G�[�*VU�@��Td>�����>t��jR�[}���8c���Ol���Ϊ�oUa=B��(���[eE}�.���
���ji�쫛�}�՚T��5��"��J���V�8K�����f�p6A��S�7?We���#�q��e�������y9��{���h�����ԛ�(M�����>�r���V�D<f��7���v��x��
�@�{�;�� )�!�p�Ya�3�ͽ��nJ�}XV��q!��d�:��*�=H�i��Xp�M��΄TM�5G���95!aWn���j����<h�!�K����/LJV~?=\:g���+��Z�&T�%&2�q+��Σ�b���zqJ�肭���_$m�0%�w��Jf!1���ܔ��Ļ�\<;gA;Q�a���+(g$�{˳x%+u<WA�G�]��5����N͍��_�l�j7ã<3LN�
fo*Tg{q��V���L��X�qM�Y��T�η2�,�{N U��j*�tU�S�L�~���U�`�[��nfź�2���縎�ñ��YG�f��8�Y�;U����ݹ��a���Cu�2�ər�2&Z�2Y;��6[�EL�9K(��[���CS}�R����+(Z�Su�6����Ǔ;#�v���<n,�ɫ1Brrt�!0�K�a���B6��E���L����F��4�ީt��۵I"��>�7��."�*l9+��%$�n��p�6D��m��ݒ�f,YJ�Z	qִ�-U������u
U��c�d9`�Wi��\�ǋ��0����;�y�OiW�&��	9��ٹU����U�C�Ll��1%�A�Y�x��὇�(*����lPs'*���l�YM���u�(�^]�I΃yJiꭗN'��|��r��:&*�s��7 �י�p�&�$%���9�d+C�r�1�%�H^o��vȲ@����w1+����(,r�:�cV��-�M?)��L���r�k_�x���w�֣5>N�&�Ǝ�e�㉈���ap��ۅ�m�e133�2Ĵ���{rj�����̞�f��d��:�T���0����)�jێ8��4�1Kej-I���e��1YQ�ԳSs�S��y���A�+|(^�A�Z�S��>�",�b��JB�2IB����̸�W�[�SS�S�s���_h��mʶ>Z��me|CBj�	Z.��Q�l\,�r����T��`�j<��Of���zѨ�aB�r��j��*WV�ˤX�,T��0�D�1��U�q�g��S�r���Ҷͳ+fZ���Q�շ�������Q�kF�Kjʕ�l�]dg�٩��6�+*Qm��TP�mx��cR��[n]6e����Է32k0D��m�5=���ʞ;�F�Fݡ�h��i�p�W%����L�1��75h�����9�s$�V���cD�S�<˩Z�Tr�r�R����z�1b�h�������^��*���G�S���C;��'%���,�C}�mb�bG��\�/:ڿvG�"���\���3��@'�I$�$�b#	�I� �$!�}~|��������X"ߚM����N�.[�̉�ԘUvI疳P���ܗ�sf��KwT�P��!ϥ��A��i7��Ju@GQ�l2v��RX-t�4�E1�%�g�6H�
!o��#��L)��!Q�!Y C���z�ҡf������u^ i�+󤣋˞������m�� �]<�B����Ǿ�x�s�lx�~����yy�ߦ�� ��5�Ҩ+�k��r����E�Pg9�����o[���ލʸ�f,��&�y�͗�K/�q�n��3�DSqL�󏢡���[z)_F�w ��s���P{���P��,ҋ%�o�"���6Gwy��(�!�i&���E��=��H:��N�&n��<�܅�fq�ğ�����*��Q�ǀ3�3C�	r��{�su�(f��+#t�N�p�2�w�	k��;K'��0��F�܃�D��.#�V���c#0����qJw��NԚ���3t�5��(��Y��&㦽C]���,X��o�}?;�a_T���q���#�]�nZ�_!�y�3�� �/բ���N�aM�����Ba�a��N����C�3����S5��G��ow�{҇��ʸ���^�H�uj��XI��y�/��C�6�j_k̑��؉����2�Oq�xV$�������v��9���s��� �	01� ��� � ��xb��;�Ȱ6Dc_�+��ZP#���C.D�u��zTJb�hi(�j.\KY��~L,��41�<�^���x!�|��A��f�!6�N��-�d���&Z�iF)+�*Yv�����WDOR˽�p����X��_,�;��8<�H�):��,���U�&��yu�j	�[����~̳�p���õ�ҽ��+�R�|�E��R���)��5���L�����GVBoִ�W�vX�|��^Ќ|v��}i���+_eݲh�ວ��ξ,�!G>2��P]&���h;�XG�̛���Ɵ�յ8�-x(�=H�i���6δ��l��^Ԩ�ը�1EP�zY���������r'��ΰ.���&�}�Ks�:0�W 'hSu=V·��{*	{����$J����\[���qPj���x���ʕ�x,s�D���dNʩئ[4:��5>�E��i;R�<�ۧNOv�1��{���3 (L����7��O���v�f��^*	�}MŜug���������')'�opr7��yzǂ� ����zWb�����#9�f�ve�W��:����Ǧ�ZB�F�
��D�'M�d�V����x9�T����f�7�}�9�r�Q3�k��`�X��\1�
�h���h��~�%�ʗ��c�۸8�%%��!��~ ~FH$�I c$� �����~���Nk����r�K��-)pAl*�Տ����h�M&8Ba#C��G�nl�62]������z	z����f���r�ou;ve2�gS0r�k��5�c�1��-�A����dh��f������܌�d&T�������v9�@���dÉ��zn_=dPfif�k�<P�ii(oi�rݝy"��OFm��K��u�1m#�T�1�C����Pz͜OX�κ���0�m�[�	��m�2��m����>B^=3�m�6��EzA�%6q�1�K��l4�ǡk�x�IF���jv�L����K�T��s�ㅂ-V���l�\P��=���+
�
y���E��W[x+�T�0V��)3�`|�ͨL`�&�<¯zA���zЙ'�)��y��͠0��Y���ſ��Ĵ�kk��'"��_�" ǘ��Bc\�S�>��rA�J��y�����;=�;��>� �;�vh���DJ��"���s�]������Ȅ�Se��i���t���v��y.�cŝ��#�K�����9�s@���[
��-�	���qG�v~�g�:ְ�"Z���=�����֕���d,s�U�W1ʷ���l$.�|)vn�y��)hA���s�ȅ�����7Q�lv��,�áN$CTr.}��9��s�N�
��n�ޜ��*K��8��uӤ�H՟�@�� �B �F$�1!�	�"�1�H��~����t��h�xc�^��m�R'���fB:�7�f&�I�&�%Ɏ��-�x������N!�ݹ�`����E7?t�V�I�k��͊S�U237��w�|�M�3��;T�!z�҈+�t�}֡��G6��4-Xu<é�k,{k��.�l�sr:l��-��u_q�.��N��a�d�B
�?+?!�z�]�`I<����|��=?K�W��_��Xuv��V���	�aaF(s	��d��q�,5�5U�+�V:Ζ�B�Q%��aۚ|Ls����DaH{���oo����hP��]7���E=�?�ϼN�usi���Ԏ��7g�J����EHA��-�I���	��fẩ��9ޛ��*{��E�V���=���[ǥߜ��Gf�Hb�%d���}+��]%����纮�}wy�[W
P�BA���UJ���'��{m��@�Z�,x������:8p�C���Ǹ�~4.������_�7��b~Rx�]j�������tH��{0�Wv����<O&��w��h���W����X��W��NV���[,#|�S���Ik&��9��G��x�;�V�E�5��1\�lj�v+��ˬ*ʧ#�7>M)\vO�k�y��1�����`�B1!#$�F!$bd!3�8s>��߅BF� �S�˚ �~��SP=s�]Qp�)���Ns�2O��C��(�^�ə�-��=õ�Cj-l�����"S�(�T�Jqo�L3ۑm���l� ���-�ҷ��N-���6���֠�g�wB����		��Fy�]��خzw�xa��{���}4J��5�2�_�c<�s�@�UeS���\��)�u��l�*��f%�P���]��X�*��jsb,,7�(D��m�x�ǎd���aU�'�Z�ܢ�
�Ǜ�)���J�i���nb8	L�aXʓ�;�Ј	���/%�u��'_<ـ��J1�k<���I�s�Y(h�2GY������Θ9RH �;�����ǨLe"|ۆ�͈�E��tjF�j�D�[��.�tf:*	{k��H[S�\�����+�`�×�f߾������M�K=U������W^Ia̱%@�e�X��0'+�hsI�^�{�GHfq��//���3���}����B
W��3t3!�&��>qiK���T;z�S"|�E1��l��3�g�b��>c63;]��Qv�,en1qL�3m\���\M9����٢T����4U��Eݘ����{aqd�iT`�/7�]	q\S*�����z��g����l�U��J�y� ᷕɓ�q5"PE��3J�}����]<<�{��s�� �HH�BF2 1�A�!�$c$#I��/�v�w�.?=a�<��{aAK�h<��J��|�	��ǅ`��]4�r�=j<��H�A�x���澽&�Ôk����\��ڹ��4���Y�W���6�85�����[����J��߆�}Zr.?���ʫ�~;�^W}�l�Q]1�U�>$���	������!�!�ne^JN�|ض똨s�,�8�G��ȸP�.�ל�Zs߭�P+��)c�MK	�%6X�!2�J�'�]�({�b�j�3++;������=�&G<����F�c�����+��q�N���1
J�w7�Z�Ξ�C��N�Pڍ���)u2�A�'�e�����/��lE�k��fW:��,�ŬP\�M�*�0UU�̫��&�s�A���7.@��.�8q@��,�	rM�7�]�(�C0�U(��vT��ck�;a�3��ud��R�bK��%x���v�F>;��}_$7V��g�Lխ�"fw˥�e�����0��>B=�-����!|p����5���&�}�=,{븶�Z��ܼ����e�F�VkG�f�zC�HX~*�+\�8�w0����j�W�|�����O�F�}|0N��	4�g:�cі�v:8sT�Dq���aL�a�j�E#vv'y�h�+����qI;O�����̺�w� ��a$b@�H Đ�I�	�!'77w_�Uu}���3�T�""�Er,-� Em�Uz��s6U_S�[��0�0��h�`Ha��3Q#o�neC�;���,�*bYU�ŷ?t��x�%�^RF��h�;n���R짅�����v�Az��y�]4�vl�dV�d�woF��gӏW�@�T�i,a�CF�ʺG�_��z����f��~h��O0���� ����� �w�u��?M4�_-ڿn���߿V�����$��A�?<��t]�6�.1������5XR9d�>R�~<�
(�4��-�#b*�d�<#����K����/V�VE6�a}qy��!���	�B�KIe�4^E��y���yd�>0����{�=�����t�|����UO��{u��z�	>[a"�vcW�Di�ݵU��JJ�`�7vV��&\Nm�=��8!��>s�\zd��	��O�)���2j�Iz+�Q�sE��΢����xKFj�x.���;@
�,.b< ���8��O�AqC�K$���+�;��*$���k>ch���by�DN���gWG,.V*F%Zm�&[�Xd��A,��DD]���;xƧ؂��ɔ~[��(���k�4�����2Z���+aCֺ�ݙS�,���#h�G9��y���j���Ǽ߻�翁	�$�(cF2H1 F$�bI#���{���|>�[[1����=���hO-k�(L	ฺ��`�`p�}+�<�	�y�')���%ۡ�]��}�X�
4���D�͜�V*<�gJ�C�gJ�C�Bh8��[M1�ܰlA�t]��3���&*ۥ5�S�9�=���Ƕ-� ���!6���ln��3��GF�W�������Le�q�NNy<�l\�7A٦;�?L[�\�	8k�TU��Y�:B�q"kВ}4�b��e���X�^�!1��7�1G�RA��J�F�p�ى֙��Dg`�!��wd�rdN���"����X�{ғ�P�����J|�pT��Un�A�l�Z�5)H���
Ь��"yq~�l�n�3�8�V�6�Q3�Tأ	��UV�J2q�ڽa�C�C�s�7���Spn:\2�v���Sz��s]C�W^�ۛ�p{\��
Z��&������	�Ι�<��G0`��L�'�+������>i�'�b�ʛ���>Ö����\�kc����_++�`�?���:�"Q���U��=�-7�`�ZO8;�^m��a�̟7ghw2~z����:���K�`��V��wSѢb���򼫂^]��{�� ��D��]��S.�r5�pI�=��E����G�g#Xc����3u��[��w���$$��@��	�0$c!#1�Ho[~����մ�~�d<��w�IQ�~�MQ�]~ݟ@̳B+z{ŝ���#�K�Zz�<��[p�I|��U��w�Ow̤l	��5��ɸ�ϲ��E�D8��1j+%�Q��6�ęK7T!�ٞ��V��t�](E��L�T��y�/���|c��v�;�����#\��C[v(�m|���˧���ØK���+jd�N��Iލ6��`������#�C�L����.��B\ЙP��WXUE�5�8�:���
{g� �����M"�0�kw��Gi!}%���d_�D�W��d���goXX]ѕ�8ށ!���+�%n�UL�W'`��/�d8@C��"���/��g)�5 MU&Y��?��z�6'���V���w��R�i�*Y�l�Y�d;y��e�� _|/=Y淩�rc�������mt�y�?Ia�!VRW"}��=3XuZ�!��rA��>�����>�!�z�M�jSQ�5l*�����,ܢ�[F���q��g�˿���RCm�n��!������B^K�F��a��-'jɆ���n~M�0&~��錢��V����'�q;�\�B�/�O7S��a�;wz7�Y�]ݬ�P/	תdn�94f�p�:Ȋh<-�@�1�*�ܻ0��3�i�����L���`�Oy�s�3��$>�!�@c$2 ��#@<�}���ߜ>��5����6y�ʲ������zp�1�����t8�CzY�4�*Qr�7�ܝ�0��l������*9�����<͘�x�tbr�܎�a�O*TE��~m�"WS.�"cl����P%��粠NQ49���(���g�y��+M�9<�
�{2;.����B0<��G�ԭdM�U�C�Ƒ��5awn��35棢-���7L�hhZ�G3��Bt�X��W$Yi$O��I�]�a̋ǵ�Y�p@A�!�۹xD������o�~�ٚ�&{&�0��
r��%A�U5M��b��}��)}�6������VH#���g��\s���NS	�0໐o8qf�kU	qW������^�(n,܅28dn=���e�:���gH���5�g�Ia#�O\�E��<D���33W�����;Br���)���L�ZT)<.����pLK���n߆��L�����3�k ��O��. n	S�=֧Y��-�bS�*K��B�FM�X�=uK��sH�+�kmP��y�E�+����3p\Fb���ő����iS�yˏ]\,�1e<��`�(0{�*-SRU�R�hv�G;��[Ld���m�=YeQ冯Fh�z=�c�pp���ݍի�7���bHf���+b���w��
죣�!��x�Gv��� <:�tW�s!y&캒�]�]\�Ƴ�˝��X�\�\�&���e�6!����waY���T�&��7��ɘ�m�Zi̙�V��V�:�JgR؍muې��'���֞=@����V�w�P-���A�����Fk#����|3�Z`�%����9�U��[j��FH�E�f���;�&��J�͵�i�oa41�
��y١������\.!�V�v�	���KQ[J����U�2�̶y>lH�=�v�3���
��ԷA$T�J�]��BL�rU�Ov���EKlͷu6\%l�����]�e�k����زɫWwx�)�SK��<�N�f\[|h�n�.]�����#�i&Ɯ��׏r>�G�s/\ֶ{J<��[1֚���'Q/Y�3���1��i�k;$�w�q��q�%S���P�}6
�p��X��-
u۔mK�ƅ�}4R�+��鸴K�Q�4�Jq��'w5W� �c��v7X귺L���8�X��x�����,���Vos���M�ܵzo�1p�I��4�4�~�uy��u�%��`��u݃P�Ԕ��5�wWZ}i^��t�\R"T;z�����u;;�����/����	i��[ ��	(��pf�p[X��/9��J�m�~�xa�[Y��?;xo#��s0TR��έ���j�k���3h�E�ew9)×2:،��h�I3|F��|�ruQf�lʗ ��[�#��m��1�ȫ$eʫ�h�{-hY�6C��P��B�W7�c�9�6����K�/����dp�|�`�����xx��]��[�����V�E�hd�r��6��g_i�Q���X	������)�(��.TTi.�Ss
P�eV����J�S�;���d���=�5m�i����.�W���q��'`r��L�-�Oo�[���6�:��^
��Z5���5�^.�OV4�s��xz:{.<���4���fc��[]r���CnEZ`�j�%�s636�Nhp7���vt�����QJ��`u���t�L��: �Ю�O�Ԫ�2�9�iӸ��[�X�1��p�K�Ѹ�2mn)5�&t ��	Z����K::��kv��R\%DH��c�q��Y�����͓J�Yw'9�ju/;'I��\W��I�i�ݐ��&ٲ2.K�E��5N���h�a���Kn�z
C�v�u�5�*!/>]���r�b���P=eG%�
*[](���"��\�U(O�RӣqB�h~��c6}櫪i�jb��9Z�i������Z�Q���L�����E�����,mr�5���e�<��Oɰ�ݵ�*ysv�U�[�I��&��ckV��X�-��je.��S&���7��qJ���φTq���\)��ޛS
X���R���1Og�����ܞ-�+�J����E����\+���Ҷ�q2�<��*��C�&���ɹ�-�R�X�-J�+m)eQF�2�SF6Z
���S�KKAK�<�M�����L�h����љ�f%J"WI��T�C㦘�QkX{2j{=���kEYUQR���"�Z��-�c���X6�x�n�L.��J�Vc�����N���w�4kX+E1�-ڹpqR����.)l���Z�4�O0�
�T��g�SSsٹ�6���Uq����������E�Z�����#l���ih���8U�T˝�F��+[�
�CQ��.4Fx���4�����<ш��*e��ի�yY6*/��"�&��c2��L�ތ�vkGj ���	O\[1.�ș��ҫ:5q#�/�QQٽ��Y�^�F̘N+2%��-e���j����靼7s|�ċ'\�ygR٩,+�.m̷�n��J�ژ��X��Gaq�r�j�� 'ؐ2 �@��c$ y���M����|��Be��r�te�b��8BKb�wDT�)�_@"@�5�脝����"�� ��j၄ԯ]uݮG.[���ƋB��'�M�A���`��2��
E��y�tQt�d*�~�y�U]�[��'�d��y�/��-^w�ޚ�f.�����ƽF:�����}�_I�<��;/@����
�Ƽ�L?5�O��C�̅�����^��~D�W��gFv�4ta�~�/m԰�'h]�qY���9�
���@����ǐ�a�q��le�wѹ�D0j��&%���v2��aCx��)�z�4�||��5#kzq��I�=s�5�r!�;[�u)�8e��P4|���_嘝s��}��|�>X�>��nc��s�vf=��y�
FZ�t�Ҥy����̼K�����&����.�|�B���O��爺��TP5h3��DFbp�h�"N����a��g�Rc%^ݩ�>�ۻ�q+qj}��\��-������CO�j�K�3C,�>�I"�Z+�����'���6OE)�~n�����_0`9��!7�t��Buj}��rc\x����F�{Ut:{�%ogBM=����_o1Zln�0��A*Я����-7�0���f��{/;���vY�J=�t\f�Vv�����!��ȣ�.�Å7��䓻�����1$$�cH��������s���<9m�ϹW�/�FoI`k�e(#&]lZ~h������D�S,ᳵm8�w��u�^~�/��By��[J���`� Ĩ����U��RWU��$^�����x{���.����`Y{C��D;�(ŰF��!q�/�����1D�Y�l�P��U�+HJ�t��J�Ϫa��	��f��d��[<��%�x9%�2ۄ��Z�
���Ց�="el)�iI\�B���5�8�BYqbm��غ&��V�^̻���2�6�i��������9�JW���J|��=�;^��G�80-�(fv��}�;"F��*�ov7M3�f}�*`�Ւ]ďF�|!1^N���sW��/A�<�l!#յ�F�$�Vd-��-��4��l��~�Df���~�;O����P7@;4�{�|���je溳U8�����X.5��^�����x����{#)�ΰ㬳y�r���x��g�����}xX���n��3��p��y���9n5uB�Վ��B;��zRq_���0}f����:��6��.��%��'A=+Y��;
P-凩�W�Ri?��ڭT�N�O]U蕦r�`����E�E_�g�Fl��}Kf]E�KW��^�ͮ�-���q���So��I2UX��s
�m�o�R(%��y���=?B@���bH1�0#��@b �O|��_�;���ޯ��g�n�>��s�z�;H��x-!�[�3���ڼp���B��ܖ�l�gX���h�Z�΀K��B�H�a~���c;B��C	�� q�a�ʽ.��;�(�M,��v힍wC���`�ɠ�%��P.q��Ƴ�Έ�v�
����P����Lً'���,Uf�}|�27�I�E�ii&9�I�Ӫ=�J�`�=
:��Ra�͡Bn����|,�
?��yPj���/0ݽ��׏CXO���$fB~kO�x�Ob_m�tYL�[��Ư\ߙ�4l	!񅇸�:�'=�꩹��PHq^��W2�� ����gj�Ɏof �z���xc	+��a-��z����\�&��B�I�8���VL�MF�j�t�c�P%�q��z1��sTܹ�p�N.��_�@��y�{d�u>��8���s�����m�u6�߉���FD�3�%�j.|�W���R���hAo@Y�42��p��Z��*:kt�x�S��l ��w=�Bd��ue
�R�IύC�]l����3��o���Ci�s�B�^��,��a�wB{��f�A��X캔�9ڰ�u3קI��^�E�V�����V�TpU��n�5F�${����1/4L���s�����q(f��T�]��t@v�)���՜��
�u�X���V]��^s~���a$�A� �B1�o0���ox{�,�Lb��S}od8v!��F�A��q�$��e���1\�%>�Ň�rlƍ��8�^m-��g�Y�����[!�sS�n!��V�;nLv��)�u��>O6�Σx]����Z3�kƨ	�	Aa�Ha֑`{9�� 	��"S�'/�Q-p�'��s���t;�S��FX��aq�a)�!��)��ڈ,��8�*t��n���{o{�ԝ�۫�2�gev��-J�
����}4�򳧌AV�A_���ZA�v�4T}�e�+�և01
nB�P�~u+\W�Ϻ��^�ʂ�Bڝj�=��8a\#�ںPٍ14��a���^D;1���	�8��.����/}Ƈ4��(�x��rKVlE)�A���U��o�	��&�)l��b{SU ��U�k
�K�v���Ulsľ5
-�F�;5���4!�-�F�EC�^��5)Y���۰��Fc��l�U5Kl���r�}��q����M	�E0'F��84�黔QJ^<4 ��{Z��a?&����j��B�z)�go)3�Geo��/V�+g����(��CY��7��P�j��ra햸���}�Vwgq䁩���1.XѝCz�)�7n�=�T�ɦ���^�Wl6��ȹ�͗Ҫ�&��`mt������g��}�g]輸\$!����Ā1	��`F2�gr�{];���I�.N�N�w�L�,/���"gͷN��b��^Y��s:N;�9����{K�vMn<	ʼYe�j���4-��
���|e��[k��E]:>?���|�KW�o���O�n�ny��㡏w��;0�78Il�2*��?޸_�?����o좺Yfֵ]�[�7W�]���۰�,�ĵ�@�$)���[H���1)�PX&Q�E��~g�㽬�wt�����XQb*I��B.� �c�:8�,k��w~���f��#B~����������&� ��yNC���O�ly������T\���K���ӷw�g~�>�;�o37����	uOx�ߵ�Xׁ͠�aa=�Zày4���2C\�j1��;k�+/MR�Ψu=�a���=/\b��YPXחI���- ��f�2mg�VZ;����[�b��{��H���?+�~#��-�vJ�/B�k*|;�[�b^��v@qi�t��ߺo�:�eН�&�8~/�&%�P��jcc�q����π��)��H3��C�W�5m�NJmBl�)�C^x�v<>1Y�q�uQ~�zm��H����f�ɺ�.��R�zi��+���	�]�`�/#p�뵌=�F��{��AGnV6�
����"�sr�Ƌ��,Ah��*�K;p�)x��Q�=���ݽ�{���H���BF$�E ,2) CY�|�ݒ���+a�q>!�y�;W�;3\��홶E���lcS��L�q�S�:�ـ�Ji�]]�P�ػE��K4�z�1��h]�YY�P���[v��nZݧ7#+�v�Fӂ=���t4�zr�A�!���~�{P�C ���[%g�3�
v���f>��;aV*���5#�x�@2OT4�1�M���.׺$�"�%��5��ЬKE��������/I�-����F�&��R2a�ޙ�g�r�x����zL�>�?J�M��n౩���,����O#n-�ǒ�c���S�(�������t7z٬5`VMʨ��;�c3�}n5��J;�yC�h��]��b���\D����Pd�eD�rw�_�2f�4.��	��F�n�&�J�*%5�$��"Ćr%�;	�ylp.Uj��t �^_m�B�h[L�ʥ��Ⱥ�ͣ_�&zD�(�Tc���JM��� ګƤCq�F�%ej�T�	y�Xspn��F݋��u&\M'9�S*՞6�=��7"{"��?��V�)K2ӑ��l7�-�Pb��?P2��ģ�E6vV����Y,�2��H��$@#9���r�`c�9ݹޯ��1����-I��U^5`�[\�[ l<@�=�Mf,��V�0\���\mfvE�*;��L7s�I�ٕ�5�dn.����>���F0��Bd2HĒ)>U��V�n���#����Xj�c��.�@x]ZN]�r�A*,W��OA�<��a�7u�c��U����X '�X����ٸ�|+L�_���K�zO�'��9�|7�M0w��D����c.���|<����c�J?B��C����z%��H���/6`&0�
��ݎ�W;i}��W�c0�|���I��e߸c���Pk�ޠ$��ꂏ.�f���HWn�a�F�s�su٪!놆1�!v<�]��H�F��z�٣'��m"=�^'duw&6j�!u�+�]ن�.�SȽ�]ڛ.xu��W�a1oc_����G����b3�8����⎟�̠ۯ�ag�'sy��KS��T���a�M0�ɠ�k��S����5��tG3���Gm�������:]C�m=�����F�K�8÷4���q'DYz�=���ºVn������Oj�1j�\3�b���۶��NG�_A.�
��y��n��̄����7�����ڡ���<�祫d3>�$e����	~�m����z��sm6��q]�C�;��j�Q9U[�D�з�&f���H��gz�U0�n\����zWw�E������}(�[�uZI�nC�g3&񗣪���f��oq��oC��P��}X�$�#��մ{tY����k;w=n����q��X���C��%8ӳ�N{��4{S��X�HF2$�@�11 ������ϿK��z�`�����Uq�_ʼ�'��/�wk�� �zn���f^,�(d�+c��Uyw>2�1�=Z�,J�}1����ȶ��d&�%�b�ᓛ���5֎~�n��^��%�� C-}=�L��
WહyŲ�c/P�Ol�zzf�!�\żE=\�J=/�b����F�&�} Ab^�D�VQ��L���FM���"���D��&��u]��;7�5���p��1�Tkpi�"Gt�L���X�I��"N�g�6{u�u�����W.͔��nFA>�C��1�d���3S�oR3r�w��/�j��"�,|�;�;��ë��Ճ�y�ÿ�JhC�#��*u�QD��~-���;�ܮ!Ѓ�3Q%nY%�fun��ڎ+��Nǻ6��&He%JT�[���ݠ&�z�����d�� u������r��@d
TXZ��3!0�`��kH�A��a�ZB���{�E�WH*�݇���X����R(�:���б���R[����G)Kc"J��:�!S��3~���n��Rp�"��C��C0�LO[���U�"�kWs��/�9�vv��*,g^H}�-�hL���\�l��=�N��kDs-N�Q�SU��9YM�)��:�eQ-�v���}X�n��n���u��k,V3^R�u��{�g���w�]f�c c ��!�1��I;�}��>o�Ͼ���X2�7�ѐ�DZ��ח)�m�P6t�=���Ceq��>`Qw�}��es�qzqZΐS���B�&��Cy3T�����c'/~�#{�yWy�ؖ�T��Y%���3"R�S�-��@�}y��7`�­H�)"ZOl��"�IUs���z������,�HuZ��\b�Q�pzg��-C�5�W��H~Bo�2�=}�y���7�s+�g|O}]�Yu�9.U� �O�\m:j鋇�yg��!I��<�34��5Twm�S�6D��^��:����f��9��(	I��|ضshlS8L�wV.l]��;#w��+�3+��q�^�-�qR�6xJl�q�	�%"S�(�
]��Y8Ϧy���5|Z���e�Քlb�<��Ȉ�R9�i�b�j~BS?���tT	�-���%�]�������B;�dz槚P1I\�B��8Ci8eک��|��D��锝\�E�kMл����}�]�C���v�"�6����ʁF��ƌB˷+"Xk	K��O�e��a�~SH7�=�)*DV�/]�gh����W!�ײ��v��;/��d��[��lf�;B���jD�Kz�C)�8:���2ag1󼢘�����e��4��(9^�5��<�l�zp��x.�s_<��Đ/{;	N��1�Q�R���s7�2?�|?�W�����1�V2`)�b,��|�.!Gl8L�E�0���瑅��VoP�}����/�kx\2C�����[g��[sxxGF�,Pܜj60ջ��>���8�'ְT4�L?2a~;�XG�����������z4(b��bH�v`��9"��Te��k���1u!���	=�3�يֲes��VC �!��@p�]PبNЦU�$^su-嘥��vY���+��k�!�v��+��ԍ������;#k��$n�z�@<��f�|�Lf-�~�'b��~o�����y|?v������@����J��'����ZsʿD~Y��9��妡}�j�ϯ{�n �ؽ�_�`�,m�)��(x�Xh��Bi?��"T�yz���Kh5��n�������{�c_�A�|�����oA/Ŝ'�A}����~�dK?��Ǟ���c���>�C��e�q�^����^���[�Xo��Uv�p΋O^L���K�y�6$��z8L�w*gT#Z@��@{��7��O���� %f���*q�j(�z������N�O��6�Py�^���@�xpV�I�R4II��}f��|�ýZʤ���xi�G�h樮؂����YSg8�a7j�U���n�\o+x�n��J^Awt�豖��\�Y��L�`����>�x��,��F-��-آݻ冘�%�<�n��צdc����]>���dw��Wf]�O���wx�Ф m�<1��u��++#���������*�����:0mord�%v�@�oN�{�.H	�������* e	[aL��lqR̹�Ѽ!�2�wI����ZV�fHi�
��(�a�ܑQyԯ7[N3��9O��oJ�#ET�ki.6�t�n�ͽ2�j������	�#��~�پ��f��&�!wS0����o��i��֑Y��;fVw����Y�x�s�O�3j�!��.���r���X�Q�٠��JmO��_$���ݝ�unf*BB5WR�N����@ѐ3��Z��f�8q�wQ����vn,�#DH�Dv
��=�Q8I�E[�	��.�f��o7\�70_u*�8l��f�Q޳.l��l�b�p���Q�=�v\�w���e�2mn�_aJ��5R�Y�e�;_oM�4)���O@t3����lbaC�i�K�@�"��f���>��1ZV�v����d���7N�
ʈU�t�o4�o��A����I�Pb=��K�r�usH0���,K[���/��V�/e6��3w��K�7ݘυ�	g�{�;�m��X�[�'�����%���������~^��Ӽ��m�����֮95�f�]6�I�]�4֤%����6uU�(�P��f1o1WF���7��fm0�r�Һ*y�������δwx�cz'wt]ba�����B�`�f������܎��e�&�Y���[��*
s`���]{yb�퀝η�٨�I��5��U�<G��J[LC�. ^��캥ۇ|`�W��_V��k�)���G���jP'��	˅�Q�r���f/p�xn�h>4�n�r�S\hN�s�<E��	4�DՎ��J>�Z�v�v�3��9.��R�S�31q�{lpF���3���.:����)a��'�Y�کer{�eM�e�-K��b�v����:ط�Y��RJ�pw�־���,���Gi[��":ۼ���Mǲ�Қ�G�ӛ�7p���ݳ�s�]ά�kL�1�9]� �4��v������Ӊ���4ki�]Ɲ��EǝL���x�Gy�h��ic�i�(��ݪ����U��aqg�x����"��u�˛2-3F��#q�vNDV�7�u�{����[��P���|�����fʆ���r'���M��zSWn���G���^s�KQ3[�����.a�j�f>W$h9�ݼ�/4��s��U�Ԓ��f���﫹�'�׼��b����_�E��`��]V�i�Ic�m�h�q��ڵ[f6�f3+�]�Z[f����s[�6ִ*��n
"�J�W5�6�4ʹ�[l����&#r��Vf�5��1�[3r�=�d�{75�
�lR��an5K�1�`�t9m-�F���Q�b�*'�ea��B����ԹL���S�Y�����y��o�V" �%�p���[kiE2ت�Y�3&L�KapR�h�/�
��m���=���f盥K��<q�|�.4|�娷W˙q�*���I�a��ST�iE�S׺4����"";5=���l��[g�i���Q2Ъ�Fŋ1�̱r�U�����\h�X�eYKAVY������4X��T���P��ur+��|lŷ31���fKVҊcDV��mE�EeW-F,�=��Of��/�T;Ou�����E*6��cR̵F�	m��cAuh�e�.&��Tǌ������<f�j*��[j�D�2��h�[k�j,[jyCu����B��X֎�S.�ֵ[j9�>h3��5�Ƹ�Z4T)Z����ZU�ES �ʑ�Q�P�S����:Jmc:���c��k�v���^���F�C18.���;�c�g,S�r�;���yݟ��Ba1��F0�d�a�7�^�_;��O|���g�~_�ԕO�!&��B�N��~RF�B_a�/��ɝ�ʹLn�Ì]�[����z/�o[�H���₁f�	�" $��6@�U����Ɔ�uH�x�\9��ؖ)�#4��J:�%�s�\���q�rm^ˈ��B훺vy�0�뾈�b���n~b\b%:�J�����kk���P�:<��mq�4R�k��c#/����fv!���Q�L:���w�F�|!1W��5�J��s�&(�������E����v��#̃�P����z���]���I��J���bӌ.vֳWn��xۙ�8�k���y���!������(����j�P�����La�e���<��]쥍�0��$�3�c%�C�T�ض)�6���9������0GD)7��e-�	�O5��z̍�Ic��ycG��&t�����{���]^F�(nw�P}���c~�`}���S���P_��h����� [�76�ș���\�Ĳ�/�Epk�����;�>=f\�y�*Y�S��k��[�Y뜮�(��+$d�x�k�����.��,ؤ(��^�;r����n�s2AuPn�u���oF�<��b��kT�_H�-�3i]hS#�χ�N�������{����!?"F"��#B1#E$���ݿy�_T�+i���%��"$��c�7�oi'
� 8հ)�,���'�rŨ;�׆y��v�f��/��y��[���fv�N� ۛ���͠�󝆅q�/^���d�{�x��ǫ\��5j��\/��i�Ē�^�*�Ѓ,x[���>�PY5]�z�:t�3,Њ�$�P*B���d��\�He\(d-�?4S�x����v�|�?�a���7�0����t��Y�f,�U�#ZD�����j�!�ٺปx=�J�ҁ#Xeܫ̪�����E!IᲶ�U[�s�䬥m�^��P%�]K^,(8���_@�#�?X��P����Jꞥo�ܺ=��@s�M".;��c�,~.�+�L�"�v~��s"�XU���;=a�r���i�����B����S�2��;��a1.]�:�Q���d�q�l'L���<�T\�[�w�Z��􆶠���D9���E�H�)��~�)9M-+���w��b;n%���t��-�pƢ컖G���O�A�E�B�9E�~+����Y��o¶졛w%94�`�bP+$=uPyb�ƍh/��S������$�FpjZ*�!�#Ki�EPB�)�[9z������G����q�r�}d����FS\VTz�#|����ʌ�'�]��.��'�K��{�3V�}�Y�e[p��'�H�d�b�đ�c$�ʬ��n-���s4`za�F�nh��x���\�-�_�(�I����s�t�(<�R`=��8�Ӯ/b�5�c�>���ţ�r0�0u嫪:6���c�c�d�G����.8�f�]\s�`���5U-�����nhu2u��%Qa^���fT��{mi���O� h0��;ӯ׿Y�Hoe�^=�4�8BAm��m	ΡjÙ:���`�%�Ts	[K��5���M�`*N;�}a�8ތ�8^$��(�̙��]s՝^J��\�=��H���7�ר�M��]�c&���M��ώ	C�����X���S1���O��I�FͶ�ld���ý�ݰ�T���G�����0��ad�p�/�|�2�VE:v~���"Qk�ytb�~���[S:���zF�t$�!����I���/���8!\O��'YJ�����f�3�5=꫸]r
@���h���l��; ���B��5�˦�z��k�<X�a���N�VFTnd��(!��p�����@�Bn���29�A��<��`z	J�f�"ڍ}U<>�CVrY�����|�c���#Q��%�4�a�y�ʺ ��@�J��}��C}f�B���PF_m
�he��eӾ�F���*,����̐��\����at�˚�Ǡ��3/R}�κ[9�4;`��R��ͥ�^g�Ʌ��=�����y��9��C�I#�d dcX�X�_�~%Ħ~�`���@��!�'-l��T�|ќ;C��u0Dȗ,!:����X�=r�5��h������-�]�@(�̮�
EL0�Þ��f�p�O�o筏�IjbS��5f�1W����/��*_��=�|�mo4�	RV'�'I��T�I���/�x�Z�P�Zb�s0��η�<7K��P(Ґ}���;M��A1�~#�L�?L��gJR�&��3�%�x�L9L"�{��ʂޡ�r�}�w>�l�;0��n��>�隅��_p)jR#��H��=Wԝ���z����,J�0����Z�}2��7��qUr���нI��cH�"��Kκ��8Ú��л�(�ը�1EP�zY������k��_�R���#�̂�Y��t�z��t��~*�\��;�;g(�\�H!{2;��9�l����C��i�;6[��S-�U�ՒVr�9�\���4Ѵ�_�J}8��9��3sH�<��	X%�a��R6kUy��U\a_[f��&l�	�bj#0�`y��j��[	�_`A��;�~'��'o40|(S�1D%�+t���/n�L�42ͼ��3v�i�ֲ�ά]n� �Sf�N�˥fTm
]�ج#N�L��b�=t��!���;#���0-�\��޿$?#D��Q��I�Q%~j��ߜ|��}�i���=-#y�lǅ�G�,4J2C#e%���
Q�.v�ⲙ�)U:务�A�Fu7��4�A/^Z'�蹏7�"���l�<e1�]PF[��Sҷ:�wP����-퐇�)�^��^�O��2:Dg���5Ⲃ�&�-:��/s���M�\��'�{�i��B�����5n��q�|�n-�rT�G!4
�`Z���O0ԓ��n.�R@��]x��)IZ���zB��"��>Ql	�M�yq���/���5��Y��t4�-�e�z����n׫P^b�%�y����D�f���Þ^x��Ӂ��4�4l[b��u�����%��M~H�2XTl[�����}ތ�erqJ�g����$5?8��iؗJ�L-�N���,;.��t�	�r�	��S"�������L"�X���%��S��{�t��P��F)fu�`�u�����7���>��[t�5�	8>���&7�v)���i�wy���gν��#���^��� \/>�R�"ߙ��֠�	�s7�B�`������]W<;d�.v��e�G}t���KẎc���6��.���'+�Qrq�3(M�Uej����B�Y|�Ŝ��ܗa4�wrx��wv��'1�{�����xm8�dʉNZ7��!�s�X�W;}��u���}�z{�~��$�(ă#�+�_7�Ͽ~�C��������h�Q�0�0f�Z�'�[j�P����X4��{�l=�MW�|�DGP̺���<9P	)(5YD1��6�忪?��a����W�7��F�W?p'��~l��~L�UU���mKgqB����ҟ@U22�-ݛ�H!��x��y�b�-b#��v������X���4,�u)�W�ƲǾ= �5O�L���A���5�~�_�=�r�Ӥ]+�5rٗ���c̨�(�嗽#{ ��.�l�X��՚��nZ�/a���h���J;8w���G������
^��U��w�ނ~�s���v�_�u�Om��-k�nd����)IT�w�>'��yՋZS.Ձ�N�۳����ҋ���7L�t�ݛ�Ui�1p���~�2��uо9��hx*��:�j��D�
V~��-��e�;&e�{z��=�b&bu���,M��3��~���1��K� H�!w'�T�a���*n%A�c�\� u	5m��{m;5'	�[6�|c����*��f!�R3��g�B/kp��L��^Jo;�٘��w�q�#g�wT�#{jh�2奺��l�0Wo�w+|dvVi�� =����ě��OV�.S�
����;s�YM�1�f�Ȕ�3���Ÿ�εss��VV��eT��][�'=v��ۓJ�[PC_������ 1 1�$x��^-��s�7�Q�R!��C�@�c����ƽc��������eAa�J�W0���8�!��f�7�r�u&��ڱ�[����fTiv����y����&~r���!(�.(`*f���S8��;��"ͽ�%c�к1��q�)z�C�� �>����{�'�U&X�LT�g�\�u:�Ԟ�n~R�㠴��=��v��1ł�hî匆�T�Ǟ/!��<�a�n����1:�5���ߔ-�'��Qi��$��%Ƅ:ӆT7���Ǫ(a�-v��^�.���P�=�a�i,%��%���^�T+��[�q#�]������OiP�hsB��7��mCK�A~J��8�T�k��͊U�'��4�ʐOP �י�����o�6�g��.ԃ�tں����P��8�~�Z��<$��'��JڝcC]�$���2��J3�?2��%_c-aG�k0c������ver2��3��m�Mc�`N)��jLj����uRqY�Q�L�*����85aq�+%�?|�c'/~�'���oT���W3��B��^�9�辍�]Gdn�VU=�G��n����o�����-
��W�-u����Ǔ}�lw�|�ʱ�zxE���g��M;:ju�WT���v
���v�K���X�"�`����k��JoK�D݌���
$��f�ƫ����Q$bHĀ�D�Ay��ߟ;��h�=O��v8��dH:"��`�s˼���]�����z|���8sz�27�C��;��1L��dw��y�~t~1����g�1�xy>��2£f^L��k	f�aJ�Խ��y��d�OC�t���4���M]1p���}O�e*�������0C�p�q)�K�S���
�N�h�@�Ru������5��w�`�Ź�l9[�8@Ə`0�} ���*���W����`��ZT)<q�;L1ƽ_*��ڹ��{�H�F�� �c1��ޭ�����y@�4��C�[����Z�1f��sc���c�%�Le��(����g��ф̋�JS��F�_�Ϛ��E@�����I�hR�U÷�k�@��bk4jh����ek�g�Eּ������˷(�a�%�1�!֯r�^c^���5z��9Pb�d;�\�<�0�ީE�k���[�.�`㖧p���zi�E�lv�f�aUZ!3� �P��lȕ})�oe���19nNX��������I��\��oPE�Y��о\��Ǝj+��j��'}K-���g=Tj*5�޹c�C,�Ƿp������S�}�H�A�lQ���ƸpǸz����M𷶫g��@��ޒ��zY�q�]84L�)0 �G	�o%��|s�_Sp��� �l^�Fǟ���I�����M��>���9S�%�l9�(�Uzi��*A.�B�ح�Gs7�B[Ӽ� ��Xt��z��s�C��VEo}>��Y��c����DG]�uދ`�!�U�!]pA� � �.򁣫�?td�*s%��TΓ!c:t��j�Ke�֪�����E��>�ʇ��0r�Q��Ð^�#�zs�l�����������Eăuܛ���fR��~c�y��@ܡ��n�G�u���L|�z?}+�%��������U9���MT-�oB/\Z�z��������Lܼ��'OI��R��~��
����>|`e��%�޶�k�3/�F��@e(#&v���
�SI��ս�ë�=ޕ��n����9L$6�<9o��<��ڟ&-�����-z\k�#����z�'t��:H���'�9���*)+�BM!ŴXt^}���z����^�-)�����"66M��Z5��C&��_J��#ۍ4��TJmQ�D��d&"e�n%���oya�{�IYq]2)���xuv)����u.�6�܍j����Dl�gn��z2��䖸��Ǵ���F���T*���J�XWv����݃�rcN6�S8�2��K��aE��M��q�W�A͹�e�[��v| ������`���-N`���$�?>�«o�}J�P��5��y��xcD|1����N�)����\b��a�fG	�����Jd�Mf"S��)ʀ(�kk�[5��+�2:i�/ݑ�|-,<��~w
/�!�*�jeU}��MF�2/g����I����H��%E�c[o}z�.��_k'��W.��u�`��!�n�pm�.�P�ߙ��-?,�,�3T-���*zn��o;����?�B�i�9ó���=^�l�:�U���Lx=Un�L�3�w^��ƞe�ڀ|J9RA�2M�RQ8Txl��zwd�o�D���!�.��kM�����sr�i�k��N*�O��0��R%�W�+!��x��!B���Q<6�T�-o%Ժc+,`��>z~�}����/�6�G`�A[W��(��gr�kvkC��"ز��ġ��O7�.2߹G�܌�2s�p��/��C�?\*��q+����<�p���銠��5�&l����qǺ&�,�4l�jb��v-��P�e�l�[�L:�-ff?�N&���
�S�\��Ιt�=��\�fee^��`\Ո�j#����TJNG-z7x/sk���o�l�mq�]乤�L�����!W-�O�����+��a�7��]وRX�5N�ɘ��eD2͒7!���M�k�;��Vi��r��ȬM�U��&��4��m��<�f�:"Ct�H�>!�g�c����=�Q�euF!c7v����C���;�)WY�y>q�e��7م*�F�âk��A�ƛ�b�F�|t�G���Ռ�g��Z�-� *<�Ӷ�R7Մ�!�_0d�W5��[��TC!����]ӶY-��2���O&��*�҆��oal'�p<������rЗo#�S����v��:�;.�����έq�`�I1:�qcݼ�Ѯ�"-�'r�x*���aͭ��ά�;����q����p6:�J(��M�-��;����	��c	yw��Vw�A��$�F_T�p�m���o��2B�.���F�'-�����͝Z�0� L
�;��aGYB��,����;�x�8���
ԅc&P���������>�כgn|Z�A�I����-։Z������8�pB����Zo���ǵ�<V:�[�H�c|G+���^jZ��3R���1$ܚ��:���㤲�˲i�
�WO�ې͌vU0�b���ع,5�/�Z2�.�5�m���l��#�M�
�`�ɘh�Xl��io�uue�aI�&�L��Έ3����I�<N�_�ة��2-xf9�1�SU׹nT�)u�ٴ�]����9;z�nQ�Ӹe�n�;E;�5LGN:�E��y]cR�h��MS��+)�9�J�2��Jߢ�gHF��K2>Ʀ�1�*k�K��qv�v*�N䷉�F&_GMuJ
��i��8�fV���8��2���W�Uc2�Yl��(���;FK�yj̩�F��I�˰�вn�ʆ�p��*LP.t�(�@�3+)�Ebb��G{1���}B�d~���x/�IxRց���k�����	�k�D�)�$��AzR��O��bؾ|�e�Ѡa�Y�1�RY]C��F��l�x@�No�18��m�����*�Y�^檾�n�cA�)َ�,��3P9�����=\�b�Ww3֕[����5C�]����tǱU���ʱt�d!�&p�����<:��0!�m�-��6ꂣx�S'��kyWl�eq�"�m'0%JP!���.�t	U�i��`WުY�r�Z�r,\�e�{M�sk9Yd<��q�^��:�+���"Y�|�Zb�ht�X�h%��Z�U���9ĕw%�"��*��V�J���q5!u|�Z�A9�b*9�m[�Pe������:l&�&�3�'\{�hgc�X4��^5W3-,�1��r��or8QMcr	��R�v��C6�"bI����^�"�#��V�D�g�"-6\�l*{���Dj�R�fS9sEU�Yp�&:գ.7 �FV�KQEZ�%�~MO'f�(�1�|BȘ���y��:�GTm*�LEb�3
[im���X.e�K�UY������n+��[h���)g�2�[V��Z��U����k-F�V��;��Si�.[R����1�Of��s�kD�QFT��ٍA��E���,���V�T�{��J��-�؊�V��������Wv�-+hm��jQkEY�PA2�ch-X���̹�

��f��Dd�����l7�m�Z:k~Y�e���ˈ�aJR�O媶�Tį�Mˆ:pL�Z��5�b�E�59<���|�F�ݭ��҇�Y��T�1�����L�.8�
��lm���PX�.Sar�%�iiEW2�4fL��g�a�E]�ۙab6��ũkF�K�U���`����mM#QQ�j���`�ڣ��j���3'����ٻPKR��z��v6�+h��AX�<n���!�^�Ǝj��Mf0O-r��bi�Gn��e�m*em#�QkJ�ʅEƂ!���pb[W(�b�L2�lt�#��J����,�[-� �Q/<õl��O-�փx��aM�~{۱竽c�{��6�0۫�Kk镦��ΡK2s�[9�H�Zk!L�j�d�в�����u|^�[·�՜q��:�&;�3؇<�]ʯ|�+E�U���*�j�$�ڪz�U��в�������f]���w�j�y(�W@�7��7�t�ｶG�d�PVW��$ǼHb4c���o�T�5�;��̾�.�n��w�&�ga�<�
M��|��솩4�=0�y/�i���=�(}���UA�՟��[�+���D�f�l��4.f�L�f��-�dJ���p&�bP�$�F�oH�7rJo��n����Xץ��4���Lz�,��qq��� ^�@�%W���K�l\U?G��*���������u}�,k"�¨&t82kO�Rx�]j����ּL��|$�*�aLv��;s�Ȑ�W4�+m��ul:�>�ǶY��zT]R��8�s����~"S��F�-���o5��R�*koWwHl��$v�[B���>m	��e`Tkpi��t�L�k��B��9b:��C,�	�ٹ� +h�)��?��p�FYw,�a��A��K7?gt��O[������8�r�R�W=�ĺ�p̛�.i@��)��^JKpC�;+�5��Y�>��=]����R�nH��5�*��+�Z��.Q{Ac@�0�
��;��\8\w�Ř�����*qfSVw]*��s&9Gշ&<�~ׯ�9	����;6��O�����h�h�Ǩ/e�t�[��!R�I����Z-�[&U�'���L9t��	�{VԵ�a\e��d=v�&�5B����~�Az��֋nb�3�7K=7n�n߾� �w.t��X�"�שyO�*AцN��T��5�U*�^�Zy�ô`i�=Pȷ=:�K�A�*k�n����Hpb�P=���R�8�Q��`�%�Ts���6�9	�[ g~��|���u�z�%�C�K�1��Q��?���˜G���M#�.��O�n���٫=�uDI^��;�Yz���z5{�����G���8a�ߎ���f����%"m��^��^9�v�z��:X�@�Z����XU��r�5�G�u��w%>�䠴���b�6��0�{�<f��]�1��=��`v`�&{'�����J�M���YY��	Du`pin��ޚ�#1��6�B/Id�("k�}��t�f0�c8Iao��*��/u�wg^���3Ću	����g�]�n��w�}kC;(1��(	I�l�<���)�d�������ul>3������9�k��a�l�	ʖ�5{zD���2,���aJ���MN�}t1�\��n:6r��t�)Jb��5����Cvy����M'�Df�~�
�'�P�4�;���E�oK���so#��f;G��R�/t��A�f�q��r��U��bo��3�_�HTY�3ξ"�Ȕ%|�Y��ݏ���i�?ǟs�r�y�i����f^�獧-��W�WF��[xƗN&E��Af��r��|?� }��WtK�mfy�q�����Mc��TXq�s�@��敘+�R�y�[�j�p��sj��o=�e;F]�����t���fJu��K"�YqS�Ʌ�qOw-�Ȗ�C^*YH3/�Q|���xK��7M�>��~���]0�RK�nx�P��8噃k��f�Um���Sw��;Qe���o9e`Tm���_Rw���g���?7	�.��գ�ҹ(T4��MY�)��@�6a0��c�����`�֘xN�jH9�9mx]���׭A�{��<���CI]3tTr�ΒY�m�B�4�zw�H��D�ä0����x�WX�V ��y�Zi��x��w2��[΂Q��ħ
b�u�=�#�� q��jY�����WFε�ߣ��˨b�*L�UԢ)z��?c����>4��Y�pB3�bF*��S*�;eW�MP��Q�ݽFp��i���\�4QF��UP����z�)�}�<�!c.��FF`��ѼN������>���ɳ�i�c�Um�>��ѱZzh�h S�n�#:9śj�qٲ��������*B�M˥l&��"���y�|�?]@�B�-q�5�����A2	j�ʖ:G��eϳj�z����5ÝTZ��3u��0Em�E���t�Q��������l���z��q��Nĥ�U�9���Ϳ"l�R����Wzs49�#7�TW��"����u8��
#���T������IW�mlLVi�rD�
��h��V�K/�Y��e2������x5P+g��&U��-9\?{����+esن���x��@�}J�v��sb��zj�a'/������r���F�3y�0a���ג2�)铵s�V�@�e�ǃ�}��\�{Mv2�楆-�C;KjF�<A$�VQUA���0��-昩�W�t�?nc��\���y`�-�}�'.���*j��]�e����p��\��>+��Hp�e��������[��Ng?5|
@��UK��G�єQ�;�������^��m �Ѧb�tl!��-�,��3��l�����|��u��,C8�joB�����^�'}��*�K7�"�5*6CɃZٖƔw�̜���/�b*���
�g����Vm��r���^��'V�+Њ�9�#j�wE4=W؊�Z�9w�Wa�x@a�-���M��ԝu���q=�ė�j�W.��г-wv�\�1t�6�O���ݴ�L��w��/�ml4�ʢ�����}9U�����)7�2��g�̈́�庝�p��?ϥ�P1g��:<��>z;.�u{Ww������������d�Gu��R	��ë�|�H9�z���+NOb]@1��+�&9>%�6A͈�A���E�.�Gs�]S�!�p,�e\���l�_Y�����;�Z�ܦz^p������)/x�s�@@_���C:��]��l
��|dmhk���V��v��I��;�j�VM����ޒ,��%S/׽�oi�ވμ}��s��]]��p��R4+u=,���g�E�C���[p�7�,��'���@\U�b>��׊�c�b�\�c�j��nmv��=�˃���X*4F@wP"��sͼ�((�6g��"��&m��jn�a,�ܼ8n>z쌫x�gj��\���Ș�xW�
���.�7�W���V.U8�7gYҬ�go�4�TS�;XJ�>6�u�����h�v�̱-3�bU\���`'�*$C��ձ�£.g��x��ݪ�ԥ����C���<]�QR���-SJ�ۀ�r5p�hY�+������~,F\�s�*{�L�H�ȑo�ȂG�o��0*њׂ۟��r�v��]�� �)_9������M�c9�1��H�!Ӈ�n�zI*���]���g�&(v���Taot�ع�J�>�H0j��g�Z�;#N�e�4/Q�����/� �g�=�5���N�=e+�N��]���3jt�v|��{��tO�z��z�9H�&�\��\��q��d��:�W8�73��S��S	�4@x�.��[�V�9:ueq�Ud@"m����RSa��T%,�4O��~��>�Pc��>�oCP*�]q�Ze=��E=�3�k�9����>%��N�b�F����Y �xK�����:>?������[�96�i8yPJT��uϸ��=>�ng�������5[��P��]�\(�͙R�R*��6e�f׏hi<�
��C?yg�}�����Uڣ��Ⱦl��}��j�(����_
Jх��m�[�HQ���κx	�v�L7p�L�}%uf���ftwZ5��s
�r��;�M����vw@F;�o;����^�ؼz�{g\�&D�N�liY��\�Ǘ�գ�޳���Ǔ+���s�vw"��A!~x��4��O�	j�Rb���/&ё�ȟ�M�W�WD^�V���Z���B�`��!�����ʨZ�è���mZ[:e�\a�ɂ8ma��)O��>��gB��	�	���=>��oa�^��ص��0�t�.�c�׫z�s>�d�Y7!�VGD�3�?B�Z�{�sGF�����c�a�M�V*7�����gM�z{n@(�;R��Rf��N�7�LGN�e���R;�%`�#^[&G}��A��^1���P#�E-wCT��ᜦ-�D����gx�di:d��M��m���b������ΎQ���?ް���6���I���^��R�`�V�W��9������}"���!�G���t~S��՜����Q�އ�Tܶ�34��g���;��k]��q�7�0އ	�����
����.z)�4?Q����Zr�*,���{^�E(�Ӥp:N��ihG�K�7y	�kx�i���mLZw�v鵱�p�h,�)�[ҷ)��s2��ܾ�c�y������b�k��'l����r8֝�g1��m�\ث��r`���|3��'��v��.Gh�j!Y��I�}�b9�G/3�K���A��ze�w[_A���~�A���ڜ��g���d�R�{LJ�2�v3��R�pwxh�/|d@6xe���u1��m�۾��*zCD�'�R�?5w_�}��4%@��2,�X"��m�F3W.,`��FE6���+�LK6�@���=�C8��W7�E\�q�w\��[�'����g.�����99��
7����f1������j�k�.`}���#��
�?~[����m�w���1iQG}�J��b�27�3)�d�1R�Y�P`����q!]xq@�(�v�&�$\Ӛ��h���t*�;]�ݝ�-��1��	'���d��JʟS*	T��AڽT�)O%������L5gs�8��@�_��40�T/x@�t_ͩ�IR��S=YWK,ʭ��V����Ex�9䓝y}ž͟%�������P�nLu�m�l�V;.1:�@I��.�ҵq�Ge&�AO�	]ӏ2N+͝�_U�"�5&#����yd�������y��uf
 ԧ��on������A�s5�7�Q���E�'��}�ckl(ߗ �7LS�3��"u�B͟\�'���!�19�E�6�$��q��r��n�&���"f����������\�6�)��je���ɾ��&��[���)Z}����+N%,���qC9�o\B]ϱ0bc=V�Fgr�3=��W���f�B����핸��w�Ȼ;�ʞw�
vӖq��bYx���fTG�;�:�"��T��`��+3�g7-���N�˾5�t2�5�㌨ۀ2�*~���V/X)ɸ@Y9q6T�\Iۨ�[����A�<���l��4eV��;�v@UɎh-4�}p�.��r����}9�h6�C8��`.�uG$�[t�&��\�f��5SF�uh��0&�[��q烢�7�͌�@���y����b����0/0��3�o�ifԅ�� �"|Qk�嶨t[��Jyp&�S�G�b������*v�R(�oi;���5�K�B��c��ؐ:�5ű,�f=�/�a�"��]���G+��"����	�Y��;&����{]�!�stM�#m�{s#ݷ'ek��J�]�xQ.=�Λ��]ݽ� �	�$���8�j�E�����u�My��
#6J��vB�e�̷%P��"��^]-�����]�F(z��J�۞=�C��T��[�cO�S�T0R7_ 4���gp;��v�G	��b�GH6����m஽� d�3�Q��2_bn�'�7-�Vvl��x�g.��ۯ_��6�ɘ���*;GG���EUggf�1��w��ة&�h-�􋭏r�B���A�r�)���A����(�Ϳt���+����T�#1��UOb��c4��x�X�w9���n���4u��r��\H�JF.m�v{�!��!uԾ������S�A^{�?�H�5��=m�H�wI�u*���=d5F;���Xt�e�J��kN\�U�@ɳ�U��ʭw�J���&����&+Cp�w"��,�6�8�!����a��;WY���P��@H�=yn	���6�l�4����k���#�͒b�8Jѩ�������-�i����z�,֙���+<'1@�qZb8�R{q�����K�M�cQ�(鬨t����x�]w�u$nI��;����J��܊ɂР�W�'�8�85O�-K�k3pp����oe�0XG:e����k�=V��;�qR��e�83�Ob�nR��T�
u����;�^�l]�h��PT
H�g��K��E��Cܑ�O8&0�v%�U�lՙ�e�s�����5.��"�6Y�n��Uző��{`ųvbE��/�����R(5�kܙ���c�O�]|��9���a�N�}U�Z|��O�*�gv�0�"�-7Q�G�^5�])ں���{���NvEB�v�ئ`�v�,gE����M��|�#u�&%=�_XQ��V��a���;Y"�&vAl+�����͂�+�ۉ
IP=��A�N\˱wJ�]`�S	N�Փ@�*&w�+T�{����T��ƕ�Ik���pq��%3�tWs+��N_e��P�\[%u&��UQ)-�,tN>y�a�e�b����/�Zx2�
ic�˽�� :Jh
)!!כ�fc�v ��|bju�η/@�@^�(���T}���6��YZ6*�'�(=�ze��@r˼vczmhT��zN��q�����r��[[7U��҉�;.)�R��	�b�ي���+#����E-ImݴK5+^jk�V�W��X���
7����är[�V��g���2[\��e`V���:[�ٽ)Mhmu�E�hñlP��o��v�ŷ,�&�7��.����8�P�2�T�a�ڱ2:�f��=��G6k�|�Q���>�jq${+$�O�M�#	p���	�W:hZ�/���f�d6{w����b��2�t�'|s�A���)Y�x�`�!{RYG&U�#��F"/�aїE����Z͢4v�Q\Lأ��ҙ�U�[,)�>�6_Y5tk�[N��]E��S3��QV��XLK�=z�L0�;��Bd�ۇi�5\����$u��26Z�H�B-�\���q`�@\�Ø���/�>Äbݐ`���7�,21w��\�B��4�z1�n����e#V���n]��J��f9s�°=�\*,q��o��E��Nļ�e�훳��0K:8b}��\f�;�2{��ݓ�����k5c�]=n��u�	�~v�{�h��0�������vY��}҇M&(t�|R�}]1�����?p�7��ʘ�oDhS뚳u�L�v3Y�2r�xj���§�cu ���ǜ+�ם/L��u ��m���٤�Lj뚃Ե;�dMB��ƺ����<Q\Yeckz�^p]QS����e�,��Loe88�n������';��;�繫���k�߼�CuK)j�TGm��֍ˈ��4���5[lR�#:ʩ�X�Vis�Z�S2nnvnm�.ؖ�(���ܥU`ۥq�z�:lM1.R�����Lʮ9nŶ��c��f8Vd���{7<f�[pb�d(�i4&�����o3�|sklQVң����W0�-̩�ֹ��Ɔ&9T��99976��J�lWl�=Lwf�.n�R��ˁO2�&4T�q��em�M�S�N4O0�ۋ�Բ���<������Q��WE3*�����
��-T-�����T��Kk13%D���Df��S'''�s�����U][�mK�\h墈��+>���X�-eNc|�K��Qg�k
��O'�sa�m��
��m̢%����m���d�L��)�UE�Z�"�6�UFY�����ڼj*��)rܴv��:J*��(����2ҬYe
���E������Q�ᒱC(�FY���nny�m*z�V9q�bQWY�+�asĥTD���UR���چfct�t�4�*5�B��ˁ���kC3�YKj�����pU8�t��cm�U��m��t�M	䯥����ߣ㴪�\�m���뒘�J�X+5g3�M9�.�J��'
uP�*=�Ǒ�x�8�d��#n���b�d3�>��ӽޓ��i�{�ko;�U0���w.�S�M8Uv#}��s���6����\�ob���c8���-�Ů5�^dQg��e��O�'W�7��wr�}�߯��`�����C |{vi�����+.���%�w�g'���ѹ�X�=!D�� ����[C����W;q	��k�
#B0��y�9���ϣB�Fȓܘ��mm��~�05c]�0GWk��w���,r��&���!�2��VY�@�k����|���t����5T���j�	���T�������.-�p:ڝ�fgL.YQ�I���գl�˕U�
��I��ͫ�P歭pɶ%�/Y�l
B��Q}�ĳ����d�bB��췉�N*��W>�eL-�Gf���l�+ʕ<���Y�خ��*Gt��:<�L�Ǐ+�'���N�C�*��3�{j'6��l�fhG_��P$9�"m�'�0^.��W���+����W��!��ׇ��G7���Fc5�bk���U��%�; �ٱ=�*�ݔf1���UϪm;C��Y��]��G蘀Y���b<)�������w@LAz�ň��
��dj�[�[��>wM)V9Z �c= ,�K�j��W��ܛY{��V�~ |q�4�@��d���/^������:ij�ޠ��ܶ^�9�Y�`����,�Gb���s#�ap��4���wug}��B�X��o DŊ�� ���t��4�:Y��oG�-��/�0��j��ܝ;=�Ϻ^��V�C3ư*�{ҟ�f.}��z����^������s�;�t|0T%��ٮ���^�o����3Z���F�+���nokwj�͙�o��-?�0^��ncƫ�o�۱�y��N��<�Fok2��a��* �x6^��]��f�D�<X�U(�|4ӻ�����r��R��~���ߜ!>�/��#RU�i�=��.a;DN�7gl�V�ޖ|�T�aK�]-�E9��{B�R0#����vҜ.�_��`�d�B�+O���Zq9p沭QA�IC8����$=�i5j��S{FI�������u�^h��V��6����Ҷ]2o�G6Z��a���v��v0���jw/���Y}�}�SD�1Z�>�����{6N���.�҃,"J%�߀��^p�%��+EZZ���v�|��;dt�6�3iH�n��+�����t#'�4]�j�b�F�v���oʗe=q�[�y�sM�󪽱
7.�[��ӌ1X�kGq�ү7ϤA��RH߳Ըw7�A�o�_j��>��#�c�h�X�v�a�vg�����m$k�h{���mH�9:J���ek��`!�5��t3��ͶJ�ۧ3�PӤ ?��^�F���Pmv&�ԝ��U]�����&���/ }�[!l��s*�lN��۫�
:c#Y�<�J�4���mkf{�ħ��\��<�lsKjmq��iՕj�wo�ʞ>���Wl�gbk�1EwH]�O�������5򌥏������}�׭k���"����X�jig���2V*�����U!;3����<�^ H���Rm��4���SY^��Nv����E�3�S)fef��7�ĉ��g&3C�g����KΈ����D�u%L�Wτ0�Pܚ�v��9:ղ�.��������a٪�N���x�]B9[�	ξ����KR�bwwS�p���j��@�a����6qzu013y�cn��<qf#��Ԇ3�G�A�~�j̟��bK���Uo�9�����yԉ臻��9�v�}�l������꺣��*�>tr�E(�{Vp��m��S�����x�o���}�΁o�N(�@'��T���};g�K�'W�r��S�H�����A�P��g�,4;�	H��H�=���}�ͳ��'ԀO�r��r���z�aAVC����\3a`�n���:��7�x7vϥ�P
�cUB�E�H����K$펑EI�WcK2U;F���M�"#s�G��>���:�:d��ke����ax"�vs.e��;����.{ӸA���������@Pm�\e,ئ}��պ���wWa3/˺�?
0������r�H��he�j�M�_���m���(}N�� Uz��?е@n�%q�6��j���3��r@�y�K�2�<Y~4�hc0��h��sU���m�w{�\��F���3��V������MJSq�*	{TG� ҩK!�b�xc�y��Uܩ�N�jf�m\�v��ܽ����g*ޝ�n.J�P�O�i����C#�w
?��)�s�5��NP�je�sҎ�[�nx״��z�H��^��|�v����"aw�ݎ{�����
�=E���Q�;�F�+���u®�A��+mssۍaNc�ϲ�ǲ@�`����BR�)��]˻Ʌ����-�N����d�l�"�wCO��z��_PAv,��^Z;=!wT�g{]2ҭ�*+�hq�����BW)��7F���b7����ߌ
�Ζ�'g�����s�L�n��[���F�k���hS��ͮ�Q]3�o`�Sx6��3^7�d��v.+ ��d�~���:�ۙ�+��Q	*�����|�ú�;�+P�@��F��:�xg�I	�8&Z����$�̊8'��n��a,�)����-H{JDMOP����18���#'A1/x���gnԜ6���/�g�s�Ʋ��� !&��9�s�4iX+��1Ъ�}yZڭP�پC�@yu+ތ�"���r��SȎ�q�(U`��dp��/f�e���e	۱��[ױ�D� {�vUn����(-qGY�^�^ys��EYZV�� �њ��CtzmA�+�C=dH�/�w8����$�ne�C ��f//xxfgW�l[螺W-U�Xi�<!v,��iy�l�̋������5q�˙����ˡܒ��w���ڼ��2*��q�g�1�95w�gad�=�oXw�<�a��:a7�>m^�@q��$yR���}��:��c��n���k[�Mfh���u��$_I����#�O��d��a�hF��8�?d{2(�g��v8)��ţ�6y.R�M�q��6>��\�S��g����Ӳ� ��a���|������(F�Ⱦ�5ɣ��W�Vj&)�s#�O���g`Ѷ���q~�d�y�\���Ӱ�*�{�4o0Ī�(l�̼-2�cs��"�sϸ�wPY] go7�G�!�|7�!�D>ޏ��J7���vi<��FN��ҡ����+��pf.FR}��#�QQ�Tud���a��9��7��1�_9����c@�/���[GX����T`H눻bR�hXJ,̥�Y�t�酩Ul�Ƽ���RZ�Z��CҶR�z��n,kԽB��S�!�N��3n?Wa�k�{����o�{��!;��^��%��n�Q����Sن�rmrJ����M"^���-�EQ�U_� P���q����:~1�6�c*H2O��4�	�&)�,�c���,ܴ�}'A��l�7� 3L�Q==*�]
�9R���`&³U,-*�klz��$.jC;V�3C_Tu�Vv#�P@}��t�[B�F4.�wqο �ܳS��K�?rt�ɭ7��ن��J��A�/��S�s>�g:M���Q5��Y����v�Σ�J�H����&Ң�4�ҟ�Q��ޠl�k}�+%tp�z�CUSo����<a��Q�ǭP�$�r����\��9]�iv��18��
<.7dt��d���5�2�$bS꧑��p���������T�ʫg����S����6�hx$�;�v�N�3]�y�����.�M�~�z�>�P�@�:������3��^�9o���h�Qu����S���<K������=�Cf>� ��Z��@'�%a�M��y�JZp�����}���E��$Mh+o7�^�'�wVc���֭��׃��kh�a�����rõF�4+�����+��joGD�P����R�	�ٛ]Mg�&J�Ų��q)ٚ8p��t�N)%���k��T9�����:e ei��~ӓ�@;�?��mK�����I��u���B�����?���X�~�b��]�����kǙ129�f=G(�c�8�i۫��ok�[^ߝs����ZR�[�w�B��ބ��"v��^a�̵yy��1���G�X�#
3q�iP�xW�va6�����<la��%�g�d�oHu����B���#�����Ԥ���>�f�9I�~����y��#�v����8��޸4�-��j�PJA��V��b=d������/��n���b��ļ�c���4<6� �.�^�Ɠ�1���3e��o�����/#No�@�A�v�ظ9Ƃ�_�����r6����� ���*�����q|OvH2�$�Y(tlM��l}s֜y���������Ca#檧Pu���eg0w0����v+OG�p;[
N����.����-|�\�=�eO���vhi��y�l�]��þ5RsuE�v�fEP��*��h��%�wr�na<�N�4q�3.��;OM2��U'Ʒ��T�x��,Ț"0c�Vє;,�إk[��G��7�mQ�r��7��4Fkz闷�*%�F/7����{oX���h"�koͼ��8x��j.�pr&�,�؛�R���OG����Р��&\&1��;^�*�u��oQb���^�QRq�{�>ܷ]��.�ޔ�{_I睈�ܜ�f��;9���q��v�'Y(�S⻼i��Z��^|�DC��w'����6p��V���m'7[�sʫM.89�b�� ��-C;K�4D�m�~�6�L��
��F4V�E���Q�t��mZo�iӕ���ِꝖh��	�vG�V�4A]|w�N�H�yu2c���ph�ۚa���*"�����g_�Y���������S��H�Rn�̾<N��븜�a<{+��R�+�l��7o�sY�b�͔�k*�mЉ<���t���Ia�#^e�u�.=�{{���87����0�EC�Ty��'to�r�B�U&�q�i��ZF��;���
$[[sF������D��9�CG��X��π��;�J~H�~]�0�Gk~�Q�y��v�k��_��˺�E��[[n�ǒ7����5֓nP�U�}�۷̇�6{	���4M3��P���>��ƽ�u�L��wcx���=>�nkIf�љ��s|p��Cwm��.�*��k۾�ٽ�0�p�r7���e�����r��w���L'�"�����$bd�E�ILMOW�2 �<�u�x�&00�$퓼Ϲ�n��ɤ�2:)��~�,w@�������|ʜ �˨Q6�18{zgkWZq
B�2�cO�-M�9�6YЧ�[��VO%����/���j{���c�n���b�FU)�ߨ{� �J�(e��S��	^����������嘃����=��i ��'����v<�����ִ=CFpq�u��Ge��X���@��!"����\��#Kd��W>6@��yª�oBMϱP[i̍���Է�ԧ��nO�|�H��2]�=83M�먞�f�ȳ�� ��M�RO����]��OD�������g�e;,��|,"�qVԳVH�A�U,£<��Xr�u����M�v����{j���qQwi֗2:��D�����8{�����U���պA��]aPS�j�2�Y�y����� �����N���!����=Ul�5h.�R��{�dݟ�^�;iK+;)$�9������nPX�%�0���K �5�m�Ջ�{�w�.���WT9{�	r;�_f�V�)������V�n�vb7��G��4��<w���� �{�Q�5u �eз	��M���5�ހ�ȕ�ok{uoe��:1ޟhW������g���e����n�)��ʲ{�4Q�0�U�wn�^r�U�c�7o��,��jm���Vl��a����^��L�FD;b�(�᠃:���P*��E�9T�Tz�;/.�b�骈]8�����<�\���Iv�>��Dv��y!,�p��Ӽ�(�:XɁ��Z��Vn�v��b��O��En�#�UL�u4�58�L�_Jr�e���,ٽ��܅e�Z_u�:6\�ƫtU������pcrc�5\�x�}��"��v���0q]3�(t��,j��i�e�����&g^s�P�Ib�=Ŋ浪��H�žC�a��W��i5�)�������z����ҳ����D�*�SM!3Wm�� 4��M�f��4����M:�m��8�v�(�6f�y�
����]�����U�e�<�]I�&�mx0���G��]�e{�B8����3��[��]��6�y����>���ӼU)����t��3{c��<Uמ�l�1��e+Cն�K.��+���%<��
�ঠ���Fۂ��ȫ��X�ًi��[�.��L��]6��u�Dcv�)+��]�ow�ź�p/�:���8�q�i��79i�&]�et��	�Nnw9��\E��E#��si~MM����ә��C.�����lT��\�u4ۈa�L�������
e����U�+��V���Q�"���L-ɽ�w�� ���3�%��q�qh�x�i��<Զ�ܣd�_Bz)��=ƶ��Jn��X�: X�&7N+O<�٩H&K�eJ�5M�5;'%�v��h�"���y�OR���(8 k�A���,����b�n�r��w��LrQ�h�++�����uz':���0��)��LR���1����R���r���Q*�+hw,ܜ��
Lڤ�ܮ�Lq#F�����;`}9��/��V�/L����<�������׶�!�nR�i�C�"���d�J Tn��5����w�)uH�-U;�u,E�I�C9����_J|,�[���^�	�/�J4����v������jN�;0�#(F��=p�����n^��M�w�q��p��7S�Ϻ�}sI���3qeǭd�]*�Y�rո�jq����;{����z�!��B��"�Y.�i&St(�D�RB�P]/Ċ}�����(��j��XT�R�Z�[DZ��j;�kL����p�(�Mm��ʋPKEYZ���b�SsS���͋�%TC���U��-��r�j�� ��-�
�jUQ�����֎V�AƵ�T�1gYtш*�s��ss�<O\�E"�J�AT�eKm咪2���c,���)im<�P`��(�Pg&�'�s�9B�)DU�Z���)�
�X�͗�UZ)m���S�Q���Zf��^[<�f����ssbWܳ�-hi�Q���C�e��o�,QOYZ����噕E+�Z����'�sa�*��DU����T���U��L�o�Qŵ�m�(��9d*�#2{=���h>�R���q���*�W���QҺCU��U,X�*�AEU<eq-������Ej{<�����e,�,Ȩ��2�2m���*)VYXUEF"�V�,UkJ�,��nnnQ6��dLj*��h����/�8���b֏�ĉ�Qy�NMR��0�V"Rʴ��|,�U#��%v،Xɪq0`�U��ܴX�����b%j�PC���ѥ7��I��K�1lߣ���~�ͨ1�}���]N�N�8,�e����*8�²��*8n̮+��^�;V�Ril�t��1�S�LV��#�wy���W�8v�;��N���U��.�7��0!)�Mng/����C{����o�V�1�'';X;�M�ʻ���^Vi��j3�H��/ ?f����MB�g#��g{v�̿r^�e�o�`�`�z��[�mq��loC�oE��Z�>�\���A�gdݩL7���D�P��c�m?O�F�W3�kt�up��6(Á^n*�nm���l�o�e�ԧ+�s� �w�y�(
'Kb�S[����A�[ҙ��Y�&<l���,�M�3Ezf|�>ǝ��}��*�5�~̃�\�7	���ѣ����¹���6^�D}��OQ��T�2}}��B��z{P]��=x)H^�~��j`Ѿ���E(Uru�ڷ�j�{��u������>��j�V!!Ք���Pg����
�:^���Vk�b�oN0�7��O�u�I	ht�����8�3�H�ee�y�";�%�.��w�w?pV��{�6��\,��v8�4��[j�^[6k�ӈ&2�(�J�y+�P[Tj�����x���e�\v�^����GwoK�y^5;�c����(l�U*ʥF�n�����c�t��=��4�P,��u�ֶ	[��TCy;4�����O�őd�H�X����w�,s�p����N��Nz�6�B��!\�\qXK$6ǉ����4���J�bX��|ڹ�K6��VMV�k�����'|6���^�A�a�b���M9���E�Ӎ�!�H�������Шt���y�PÂ����6���#H�����>7'6�9����=�Cf<�A\y�[2�1�j����j9��N��a#����6ZFw�ir�'ص��+���Xg�8�iԑ�p�>S��\u��q�8���!O���ϯL��[���\�ݫ���a�R�K�1�)�z"��wp��e0�D% ��	S�=&�?vUo%�[���J���@��1�n��C���z��y����u��J�yfV?q�c�!�*�C'�YEN�je��T޺p)��.���3��y���s�:�,��jY���e�zZ���͗3�|1xˠ8���=;Fz��m��/@\;k7�'�9���5Q���L�i��F�����c2�UW�Q�5JL���dc�bpͻ��g�p��X�A���_t���٩�����_!C�3r�$�绦�����Q�5
�t錃b��e']Z�9��|/�9~}�.b�����s�W7@�}#Lt���g�y����kǷ��^3��LgT��aA����6��-xS 9��%�-.ܞ,
#>�-���q��̻�.я���{�/@����>f��SE��D�?���%\ �p�ͬ����Gk���:��������@=T�Sg�&�/���ڸsY+���`@g����ZI������Y!@w5��_y4������G/sFTV�v���d�4���v��=���IͺCS_����U�<������E�t�"����E��k��r�O6c��0�)�Rіg&��K�B~=�V���o�"�BҸ�m���Na���h�������#����w��_��6)B�V�@sʴ�����KQn��:��=0����L__b����N���s��(�ȭEz��0��}�ܘ�a��4)������3�]^vX7�-�9�NYa,�{���(�P�r���hT:=�����K�1^�Z�M�c��������X�׼-bΒ�s��^m����'L���o�5�T�*T���!���.Y����3=}��e�sw���]���l09ޘ�z�-H$Ϭ�Wv�F�2�MǢ*����bs1rK�EJ}�7��϶����
���s�>���51&�UQ���GN��w��m�M]�W_�mOM~\���$r��;�4������276qj�e�z^�y�{x�w@�c���J��nw�s	�h������P�l�Pؾ�0w��������<��^ ���nǫW�0n��W�Y+�O7�/6��u���䗣��A���빫s]S��n�ɸsV���"�8ABl=%"�\ZڱXc��1'Ti��y���l���"c'h���ɦ��tSǶ�r	h{�5�~vk��6�ugU�}-O�(��˷t�U٤�v6��SsNz=>g6�{]�σ*�19������;".7��+>�0�ZR�u`;WQ.l
��ü<v�O@��F�5W���ot\/C�W�*j¼�����N@��ޗ�]�&u�	��RU���^�~n��(�vz�]exv���aYs�a{����$j��ͷ��Ζ�َ���3�a����5���t��[��������E?�$�+"�y��{L��k�������b�ܬ�j4i/^G@$��&<6շ��Ԥ��S�+*��o}�i�c^.|�\FV�=r��F��"���M>��'9��v�Rղ�N��M�5��mZ��ћ<��oP��,nv����T�t���K�wgC�jp�������/
	�u�b�O"Z:g#Z{�7g� Q2��3:�+������V�bV��У*t�S�]~�z�iF$R�y���I��B/�7�nUB�!��G^V�����	�B ��R��~��u-&��9���O���y��9��-s�[Kux���qڧ�2�e�������:���9@��T�
q;�ǯ��Vrv#�l`9�ϥ3���Fl�yf����=4-�	�TٌN�՚��>]4�t���L�c�����<+5��6m�~�jW�1l�v�wc��\|9'�����7��{՗����9W�����	7pԓ�7�&r���2��Ѫ���]�;-wUɓR���a� ��	���'/i��jS˹:9����L��LΦ)I$�`�:�P�����{�ߏ����cW �<�
3�OӐ�4 �ty�$jt2��y���8��O�s�s���W��4h�	�%�%k˝,�:ge`�O�3F�SR��.��.�vd@.�v���	\#��+�'�����|��sMBf��=�]�%-p�p'������|P=�J:x�M�a���=�;;�;�=Q��?N[p��P��s�\�7�=�Cn1�R�L���E����n}��}��ƀ@�W��
Ԏp_�~���}���DN7��a������6�x��0
*�5 �:�j�n����`o�0HX-��}��ϙ鮌G�� MR�ǉ�<��]G��lǁ��+듰̜��"���/�����&�����w��w�.Vv��k['��J�,LX��5N;Mf\����E�p1��߶�!�/�{g=Qڪ$Q(��>]��|�������72�v��x�U��,N�m�i�+:�7p�C}���?w���
_��\T�Ȯ����O��s4Z�����V)�_ASʎ���9V��`��{�Ϊ�:�j��&�a�b�����$�;ɺ]��T�[v�
`���c����ON�3��z�<�O�w���.����&���sy*Z��a���'<^X�R����\�����3g�7��F}p2�g��'�Qz�3�)�qY���4nۈ��ĸ���[ ��s
|��0�5�������l3�Q'�7�vz5�Ev�;*�&8Oa�3��wG��W�P��Xĕ�+{�dy�{QN�����mk�i��!YT3[c�lƘ���.	�:$�S�l�6�SabwVTA�'���)C]�x�z�����̾q��XiVA�{嶴D/^�ds�黪�M�z�:�����P9�w�w���`\���u��h9��^�@�ݽɍo���Ϋ~�Z	5Tu�,���c�%�n,3mY�}gU��$4M�{_(�	�i�*%�0V�B�@�~�#�o7�9>yR���K6��Č��q2��Q����藉jР���Z���ه������Y�L��W��i��z������o�g[�ȝ�&շ��=�f!��^{|�y+1�b~�0��}R��u<�J^������L\�`�G����W��(�U.��˂���&�ix���#qwﾞ��q$Cΰ�N����y��lI/	W�*Lq�qsꕳn�vdX��%4���,����j�O���Z�on�\G:Xg�������k���'��*t;������s}a�	b~��#h��V�G���c+��]"�Ce���WJ�a��òᴁ};!�g��vÐ��� V�]�X�_�^��/��H�uwo�G�|��4:���N���}]�WA4����[p�cW��\��nO��	�^{N;��*�3���6X9�G��s+y����&�#&ZOg4?V0U�o*��O���%��X�����^�G1T"{c�-i\�4C��� q��ĳ�%��n�^���wG���s�VғS��p��YX�ͬ�yH���b�C���=@ӹW�}Ժ��vo&k�D'�,�=*�:��+Y7L�h��h��U�{y�A�3҄��#�ձ �ޮ�	{p����1%��0�����S9�~��>?�c�ڼ����sD*��-x�_�xӞ��s�l~Ƕ�hk����!�����n�I�
���Ũ�;�T��|���|�j��KsQmx�t�ci�ٓ�=�"�;�7:���֢���M0H 4�w9q��7�Re�4�	��Y����x��}"�^|�,��)�����ש"�S�.�:�w>L����3ƽd��r��������C�|�5DF�����;��̕���Z�4/�w�,��� �WpY.Ƒyjni�쳡W��OW�K&s�����n�:��2�H���	�Y�h�:��ں�s�E�C�̗8&&����lE�=�S�˧,��]-�.��y*
J�UOE���'C[�Fweލ�ݏTE��p���!(�CV�wJJ�/�vv7n��s��qg����^~���s"5��1 \"���Q\���[_]��e�F�M��"ci�R]E+�����u�-��zq�7�#Tn��]�{~�E�Munn�M�[�m���}U�:;�5~��8g�~t�j�`��� ���J܇�t��B�	����^�y��q?�����l� k$+&g�J��kV�^$��!}��y��Z��F<ub�q*Ap��D�+�w�ޮ̛S���K5ga]z~�j�[���j�yd�����r�n�+��w���2v��s�~�o��ml젹��"�Q���F�1������(�;��ig�R;O���9{���l4����w�q�[vo�o-�뒒���i��b�,E���Zn�2�K��RQO��`.�p،qy�9�j���n�X���T�<hi7�A����0E�ێ9�#�5���I��Y�['ר�r�Ԟ��a3w��v}���Z<n��;�l��A�{���������9��툻���l��m���.,`׎�FF�?NC!���k�^lof�SWeأ�y�U*إ	^�<��M�J%ⲑ�wz�*�Z�����=9�K�����U�-Tr��n�JBY���m*.*���TI)���e����ֆ��ի�,����<�s=tL^g����4��'�3^f<8ٍ������4�qI{ٷ��}�vp��#��_�:o=,��G0q4�;'M�� �&��ka��k�zd��V�E[8�9�Ee��� fж�C0���(�N��nf^Z��3�TJ�Z�ԭ�웬��J=,������f����9���J�d���n�V�->�Y-�NK�w��{Է��Z��k7�Ƹ����CGYm�Q�Hy�Q���͏u^Py���ێr�;��g�)�V�=J雿j�I=&��۬Oj�����^DS	��D�w�-��ǫ���.ƈ�6v었����'3�vSڤk(�U�`���V�5�g���Ѡ�a��x���f=�S��y������N������̣�\��^�R��#���PV��:��l�s���=�D���7�ga����֩3t��C�����P��+m^˶w����E�c��:S@<�Iz%ɑV*<c�2�#��[�%k`���C.��*ۣ�R��,�a�Zp �fB
̔ �$�E���ȬrH_u��Ewe�R�
�+���)1�l����u[�7�g4�0�*چ�\w%S.i�����}�����i��Rj���=\�T�_t�Ppy���YB�2��o0a����5֔�e�|�=��ݳ9S˱��ΥT������$�7&\}�_:�v6\���_�:�Kj��)ԩ8���j�U�
�ip�k|_+.bĊ'��kM�b#5�Ң�tn���lm��i���P�Uϖ�c���m�eC4ӣr�B��/QڏN�Sv�4�bu�\��p[Im>k��tΉ���<��L�H�Wv��3�A�v���	�1�-[���^\s�Gf�L�zH����vA�t2.�n�}�?k���'q��:��%����UN�&���.�m�;���'�<��Fj�zR�[C���V�ܚ�oSr��'j�}��\S���^Wz�b�.�����l�h���ZӺ��^g�7r�V�hn[�]\y�����[U�R�:��,��h���7�EYi_S�����ӡ���W:��}�^���O5ݭ(����#+(]I�+�tb�j���\�*q؃����;�p���lJ[q��z�p�[A�0KY�Vش�:��ڽ�8���ܛ���
;��x(BU��P�6s��sܬ�w�q�JZz�N^���(ŽwW9�91�9�ub�1UkBଷ�]j��I,op�KwNm��l�7@���S�<8�1�2c���'�2N��k�bU����yC�M'j��EP�ˡ���M}Wp�'5�K��us����A��lВ:�i���9�uE,�F��R�ef����\\�U�R�ˆ�����{�{'Ӷ�jcv+�(U#܅d�O��j�-�6cS�e��0䧎Åd�����{�d8�PK�SpS΅�����NK��]���*|B$�X����_tS(t���r�ܸ���u��"e��}��ƪ)�!#��M\U�É�'-���n��IR��J�)��k�X,YmTX���+�qߖx���Kh��UT�e���z4}�Y����{76��UZQ�*����L�̲��""���4[|eC)iXq1�!g&�'�d�����b����W�AMXQdY��*Q��+����[iY*�����{6UT�QE]�*�F��D�5�fB�)Dq��b5*���fNOg'&�٬�M��Uam���r�=�՝C<���l�U�eE��P���[,�����mU=�*�g�V�hU���B�QE��Q�P*�kYR��f��ٸm�7-%j�N�K��R/Z�Օ���ƫ���QkE�)���Y�R��\A��NM��cPU�Q�[Kj�Ŋ,Z�P`�v�6�-lX��QK[+R�R��i��̚�������*�Ȫ�,PUm�C2ʊ�h��X �j\�Qe�V�,F�*Z�VQ�
��R"-��.�
8"Z����F>Y[hi��Y�M]�5�d�{V�_���mS!o����3��%�I���Ӌ3��S�1rR7v�R����x�W﾿\1g�����"y����|tI7�*�UB�d��@S�v�.�ɝ[���ۙY5x�Dux��E��wBKG:�<	��G��)#a�.d�,~���Ħty�4�'�z��N��8༉��S|iI)��^�ͷ��ɷ�kcW�X��f�
��j�D-~}��2�ؚ���������ҙl�ں���/��J/�e�(kf�i�.��d��?7�po$���q�u+У�{ޗgwW�e�_�Mŏh��޾�R�A޵<�qV��3s4���ۍ�"�됵�Q�Z�2��lo�o�Ã�0c����!6�囘��Q�%ׇ즭3����;*�1�{}���4�a�h��A
�m^��n;t�|���r�]D��:B���QE�p�#����V\L��V���h	�����"m������H�Qk�I�����ʒT��fOVK�#��ޖ��k Q��f�C��(�]��j�u1��kmĝ9��Ю��J[jB����R����U��˴^�o�p��C
�C���]P�UqQ"��l�҄%q�+W�GWl^N����dq3Y�ѓ:;zB�?vK���b��ȷͦoX耭�Yl�tE>�D]�oq��a\��\[�)OVC�M�74G�}��5[���`�	�f:����"Z��ؖ��Ɏ=[�@;�ύ�5�ZO\
�[��.�Ɂ�URǝ��Zg+���r~�LHW�(�̓^3����tSذ*���{zN����Z���}�j}�)� Ԁ؉6x[�R�W�T�J@ܷI�w�ֽ|�qV0���#�ՋC;�����݄�����cY?����AQ�眕~s�z;�(� �<+ϖ�]^����@��d�އm�+eq�ŷ����Sg]'`�UҤ��G����.AY!�.�B��l֣Bl����}=���fﳗ;L��@�q;ǎ{���.��^�:��3!�oTAL�wz��ݚ�W=2�Ĝ95�����W�nɽ��}�͏0����"���Y�y��ƞ?_���P�{൏gIs��x�j�VK�^sD#���{��{#<�x����3���c��4I��dG�%���iYv+��0v�M_�)UYC6��c���=��gsbswTMvD�V��Ё���
�F�S E������t_&I�w��*ѱfwR����-�r��8�)V�xj΀2�ze��ue{�p��3����n���Y�)�ݡ�n^i��	��P6��+�]7Zb�{`v,5�\'���d`Y��VqZl"~� Qѝ	�rwL��"�48ɞ-�(-P�x�=׋b��sV"ϱ[��� w��<*5h�Ǜw3.�Ԣl�a���ϕ�|u G|j��-`�!d��D��<�J.i>Kf�Um�O���xWv<�_udI�M7����l3��%>����9VT��V��8a�6�<t�X�P2��K�����ӝ�WR��Z�g5S�o#���Q����Q��(x� ^�Y^�)P��p�Z��$�]�s`H��郃4��{�p���Kñ�p7Y7/FB�#mlzC�tϥi=>H�uC�x���(�f�ۙdڹ�c�g��d�Y"�e�����a���,�&�W6���^=����*x1z��TN��^.�sp�c	&�&� ��ɭ,a�
T��XV����[%��W�Q�_�E�}OCX�k���v�'OE1��v���,���'y� 3=��wng����c���~5��}�T�\�j����ɞ<[��*]c�Ί��Er��.��*��<A����&��%�"�7I������&����'��r���Ig�ō�.[�~��5~���/�0Þ��V��:�m\��634�P��z4?4�!����a[U�Q�����uͮ�i��'�T�Y��Olng�.�������>�ϖ��-���7���5Q�;���g�������!�v���N�|�#�8�\e߆_E'~Z���qȾ���]�5�)���`xx��YFp����G< ���ǲ˾+�F���/usm���&��y�����'EwHj�2Ձ�³�"4B�9��V>��']+1����7��,`��z{E�'��������z��Fq� q�4i�#u�**�kۗu�c4�Ebpȗ�yJv)�gu��xDUd��^�.��I���;1(�U��m�Z��UM�Y��H��=ȍAڢ��X‎	�e��pZ���*(9C*�r���QmH�㑰�<�|�]L�^Jw?�ek��Yc�����N��5gsk�gX�Vg4��cd��|2,����'���چ>���!Gm��H���_�q��Q� �LK�=�`��լ������l��
�XnO�oL�%�-q
��ZeŎ��u���Ynr3�mc\�F�.i��d@�>���SJ��/�T�oO�m���7݄ļOhԂ�*�FW)3���U:�l���:*��c3B����3/�B���a��1$�fI*Oe�v������Xa�@͍�꾌�F_r~�d^���)X�\k�v/Z���W�a����ʾbŚ,_97���f��#�`��1�`
u8���ܧ��G�v;�Wa\����Y:���*]����DS ��-��}p���|���=m^�)BnP��:��7 ��v�is�6�������b�iwf5���L���9���k�����efϚf}%B�����6���6�d�)T�]���&���#r�zv%4�U|{uWl"hmAO2S���R�%2�%�o����7{	G�����7��Aʆ<ׄma��P=cb�u���%n�m.%�������v\���/zPwr�n�N��FC����JT<���E$�����z�ц����?2����s��}���6�x�x�E�����D̛7�{��-�r���d�ĺ��-���v����6�6j�=ʈ� �4]WVe�+
)m�]�	3�5�ѱ}ft�o6�y���{��1Tذ�ܼn�j�j�X��E�~T�H׳'ݙ��/�Q�C�Qys�;d��]�p򮎽?-aD(���E�#6��<S]t������&.tQ�|'y�²M�W~�]L��$�O�����1x��J�uKy��zxu�]väړ^K�����ӓ��`�6�	��f�3�FN�3*.�V�@i"�3n[PWC�3�}&��o$�y��;u�7S3u�kFooO0���Pq��e7�L>r$���Q�*j��"7��/Hx��Q�}�w0žb�j�X��*8�+�V��7`�`s�U��MJ]]t����[WC�-H���7�Q��c��}^]�&�b'J�$Х8{��[5xׇ%��^����F{9�B���@�ΨU��J����`NE۹;mw�x�i\��q�mޢ9T��tyt�2Kd�����UL��P�&�W�T�$��^��/��@���������Z��5!Zn�3���Wn�n��,L�K��|6(V�@۞W*j�1�`�]�����ˣΎm�v{�N5��	�R�1���LyMռ)c�^f�i�h霍X�%�4iwI�y��,�M�k�������0�j/Q�4�|�A�7R�'�Ј�]	=?o~���{���E�3q>�To�3*V^��0h�����D99�qc��r�loKu���}V�c�3����kw7W����Al�*���^�J�o̺���o?Ǳ��ea�yW3��1;]^���87�L᱃#!�/�%��\z�C�����I��ʫ=p���N�F��������:,��=k`�̉�2݊d�(�����\;pa\���N��(��X*=�/���p��B���"2�M�%��L'3��;i�\�@i����C�|M)�AwW�)��\���ڇS�RJL���B"�U-������:̷�]^��iv���\0�4�u����� ���$�*�5����pq���u��7w�U_�=Y��������ynu�wڌ6֞�����y!|o*�:��go�eڎF�)�=25��v�d�ʣ����C�Y^��k�YsNnH�ط��9ظ�?k���s]���nE�^�W[�?�JR��������39���9XC���
�ؘXG�. �A� m����0��U!�fq�z���
�nשF�N�t	�@ۄ�O��4W_���(_2f����M&�f�	��݈c�;&x�M�|u��H�p�
��y��!G3Ya���y����� wO~&�V��7Q6u�t5>4�,�A���f�NtwOt��n�*]V`υ��v$oR�`�eq~F�c2��Ր�sM��Pɉ{��/��L�c ��S�ug�%w����
ݕg�t�g&B�T�ﵹ��g��`����;2��o���m Q5��q�U�$�6MY>�`���y�@�!�:���)��V�f1*n���-�=ߏ9{�=	�lҙ퉵��k�ʨ[Ԅ!\�������E�>��sҩ�ǍY�R�6�\�1�2_�1N��4���й�%u�ӷٳ��Ms���Lnd�1��^�HE��_dR����e��r'������#���w<ƚ$kfky�9v�� t���g��݁�}�0�㭍y�3tfn}�I۾n��K�e�>�m��`�!��3�A7��@�6;�ǜ�p�_&;Z32��f\�����y�7-<�����qc�ׁ�(�ا�F��s�����������]î*�Uʠ7]�<�4�,V!(���[L�9�;����_N�<���|�ӎ���iѱ'T�Ƀ��#݉	ht�6�4���Ǎ�CD�w)�8m�e�6́t���P.�X&�ʲtEZ�Tk���G���<&.�7�9�;�j����v�9���
�7"YqĢR����z|�͜�~K6�nČT	�RWI,��*ٓ�r:���}��yjf�h��y9ۨ<l&�!�Dx�pԏ3� �J�EU\u���T*�-��	O�f��Vd�N`��� y�؝[7��;�%̸�y2	�Ǭ����L��&x&�W��h̺����Fk�_u����|Ecx�y����5h�;��Ӈԟ,�E�9�׊A�	�X��k_���=��>�g�>�.�SA:疫pw�����9H��\j�KVj��a�Y���^��e�1�G�^��{���T0����Gk�ۧ18�2�����.W����#�?g���u;���$e�L�����0\�u��)>�5�;kb5^ɉ����f�^r��;��G����E��W�L�;.�@*�m|g��vA�nT�.�3��ۇO(��bī򐮶E��C5����F�Ec���F��hs��x�ڮ�%p:�G�NFl���{w�IE�L�qݴr�	�%�u�P|�dòq��$V2�	t�},���`1{�h�!ꎾ��r�D4�^gڍ�E*�o��}���s�Os���xh��]��7�m,�ke���0���T�zi�����<��E��Y��Gg�цsp��9@��v�[}C��M�;�t΂���w����˴<M���h��]fl���"p2	�+�v�</(���ߚ|>]>e��s��?�����O��	�� $��		!$'�S�'��I	!$#��0���D,���Ic$c#b�b1�)@�V�($!�$ � �� �$�#	���d C{�44�dHI@�Q�!(T@� 2@0�d � #$ #$ 2�%  D� @� �@X� #  FH  D���JE $�B � .`� a H�@2@$ $X�c  F `,�$ $a "�H� �%H�"� "�b@ H��  ��H�d ,P�D� d�E�� �F,H 1H�D�@"��0�f0Hċ��X����D��E�b�#�H�F�F$`��X�1"ĉ2@c1"1c�A"1�c0��$F,X�HB�Ĉ�,X�@$ 3 � Z�	!���C�P�����	$Y!1 �  ���[������'���?�������>����)���D-�����������\ I'O�`d���G�BI	?��0$������?A�<>��2���~�� 	$���~����K�7�G�Á�S�R���H�m�D$$ H�$��
@� ,�I!�	 	 R@�2�� ,� D� X@�  � � � H 0d 0�   ��   �d�$ d� a � � �@d� � �2H� 0@ 	�!�� d@�	�I� �a�$�2 ȐD� 2H�H"@� �  � ,�H0XF��w����!$$�P �@ ��~�|?��_����P���4�a�3�����P�t?���k���鞐��aO��7g��}���2 $�G���?������� �O� $����=��RHI��?y3�I $�������z��`!C��_�y��Y�h0� �G������?���?�B I�{�Z���g?Y���?� �~������� ��B I��:'��D I'����������(r��g����5�>~w�ß�p $�C�������@|��{'ɳ����O�BI	?q5<(`~�~!$����������B�/�����)������G�l�8(���1#�{�|�U�4h(EBa
����*J�:j)�TT]2��6�AJ:i)v@k!���U�Ɲ��$֦�֭j�%V��2�fԪ�5��f-��kl��+m-Z�[kkY����UZ�m��+6�,E�J�l-�[&�-
j�j�6�����k]��N��d��f����r��[$���Zk[Y��j��(�ي��J��d���,��[�q��e��D�jm�S#n�V�ff�m��iR��R�h��R��R��˕�m|   U�[U����u]��u*s:�u�hwkvM�i��u:T�5���AM3��SF[��8U4(]��qӛ(9�7
�`v�[YQbF�j��8��J�   l�<�a�C�СB��:(P�B�
9��xQ*�"E�d(P�{�âhKֵW�o���R�ָ�.����;pn5�n�n��l� Gt�k.��[��J�׭uH�����{�\�MTM���   �{�B��iӶ�jj�;e��v�;�tS7-8�4��uۣu6ʻj�[�ҝ}ۦ�m�]9L��׳y��3luZVۙ��ܮ��=S��uBU�h�v�V��w)-T���5��   6{Tף�wZ���NN٭�m7]�)N�SU��d)is�uMPuݶ`*������B���wN�5@Z鴾�N�fֶ��u��*͘��   ���V������h��v���������T[uW(M���WF���h�Җ���6�7G\���kF��6���\����=cn��jU�i�mf�   ;�+�����UB���f� D�T�ұU�GD�;�PKZw]N�E��7u� �;�p(Q]����:6�mi��:�m���nͪƆR5[|  ���7Z�������% ��  �  ��  ����ӥ��  �[���7oy�*��f{V�V�ݽf�m�v�]+��  �� ��ٴ� ��  
�� P9��  �ͺ� ��  �0 
ݴ�  ���}:z��kf6`jӣ���kiJ��|  �>  >�p 0�� 	�� Ml  s^�  ��� �uÞ�� t�  =gU�  ���=��Z�f��Y���-"��   w��: o��)� � (z�ҝ ��q��<��  �� ��X������n  �O��*P)�)IT� ��F�O`��SS@ ��%*SM 4?�@QI� e*
�  f�����~>��h��Q�#�q��{�����w�Ob�b��g-���0T��j�����_W���=������1�co{`�m���c`�6�����m���1�v���?��ϟ��I}FfBɨ���Q�D�]Оm�1��peT7�
�n=I��uQZ�4�xZ�N^�w�G{+r�܀o1�,D�YFU��"��V��J��Ȩ �nϘF�͆�L��C- L�k��4���WL6@�� �mb�X�8��MAn�]�"��ar7���с�#�#p]<[�,+;��	bXP#�B����b�wbg�^
ʟA9��E����fm6��`�U�d�w~�k](�7���-te����`�eVj��P�m.#�< �J�½)i�6"Q��
^�$�]���V6�u�۰~:�k��������Lc���Q؋�9���D�P�D6dq�S3.c�2�V	`�m4�iaܨoQ��W�+Q�mb�R�jVҒٸHZ�pk��V�Ս�fM��O�˻Wl�� U�#������*m�j��TsM&ؖ���|����	�"�5��������#R�T�(e��ԊP�EZ�M�b�V�	�؊��9;��,R��3�h�9���iX�U�p0�.��St���q˒�m;��k�.�j��N��	*[YU�[`�V�9�V@�n����(�S�4�
�N�GV0��[�Y�`��CV��a�ɋd���ՑA�`��,|��V�b�(q�]�	D�(�o�u#|�rS��2d1�5&la��m�JY�j�h��%����ֽ���7yx�,��cd3!�!�"����
���.n�@���U���f7��c;�����E�C���`�6�޼(@1��5v�$♧#"��6um%ZR�B&V,�2�8,dt�G������9Rr�z��5pR���j�X`9sY-�:���I&^RZ0� 0e���Y�����!u��[��I�iH��u�3�f�����*һu�h��1��)6]��N��m�7)��N���e)e]JQЦ�;Y����3%��T�v�eM����#3ؚ͡	���J��.Q��7n�ƨj���Xlm���G^B	���ܢ ��8M�P�l-��ַ�D�;p�bŐ�����Їrn�h����Ct����p`��xx~w>�� ELun6�]L5��J5�4�*��F=��̓E��z����X��ˏwd�Ĉ�pV�9Oj
��Xs/%/�ە�[�RpC��4��
B1�x���7Tח �YZ�l�K�h�ba
ӡ@b��ݒ�����f��.a��T���K5`I���F��)�����M���~A�{/�����VZbɶ��\���ӛ�v���c1�'J���`y6��y��1Cc�֗�!�E%��3�(ì;Z�i� MQ�K^���*�� �`�Q�b�1췓Fi�7�Q��&m�t�yE(��/,���,�tb�kh��I�Rѻ JR�t�י�HƷ�]�ʴ�٭���YZN�}�����݉M�im��-�v9�"�4���y. 5*�͵��&*�eQT�
-Y7r^�D�{M�lP���
�J�7�����L��2��+r]̆`.�$8�mЎ�{��V�q�=ڧ�K֎���̺q� �Ͱ�MF���ي*�*�2�*ݵL�6¤H6�ahM�X�6J����3KGp$���;�`����z��Z�0b���雛��`Վ�x,���e1*,��bQl�5��BK���T-+3V�PVࡨ�k]-���1h��=��,��S޾��ͥ�vpi�Էu=j�Y�6niͫQ�`:ɦ�L��]a���[����I�� ���o>A�YQ="�t◄�Dn]��.fKZ��i�n֌H��1U�j���]�GNҐm�j�y��Ԭ�4�׊J&�	"��eb�F��$\�[�:,`6�#ЯVť���f���q��MH�NlT��6W�[*K�CԷ))�u�����S�̪aZ�Q�	5-&GhT�%Sb܂��5l�F�bΥ�n4�F����q�O/Z�i�%���� ��k��Q@��v���:��^��!�a�
�H���]*[K^iS0�<Y��i`5�P���f$�â�[şaŴl�(�ІPKU�U	�)V���2��c��W(:��*��u.+�ų��lg㒃���j˖�n�EeF�ꬓP��/�+$��K��AF�^e�32���QXdՂ�0u�J�jp��䗬-еMiD*8Ɔ�0��i��T��j%�<�7e�'[��c��(I�Z>=w��.S�����v�������Vԓ*�:�0���E�C]n`����
�P�)���v0TL:W�J�CS#`+�v��1un-됾��Q ��%wRN��cmU�fV%��[�%�bƧo%��Y#v'X�ѦN�e��v*^#�nAG.��uD��2��l�-G����E�֙�B�S$Wm�ؾ�]�M���meF���ʠl��sU�ksD�غP�����^��A&�1޳�#~��b��_<�m]`A��8&@-�Qh3kų�6�8�ٻD���q3��]A��L�0Rf�����*�0� �Z����HX�܋w����D�Un�+��m�Xy���:X�3����Z:q�fIgE0�oiS5�-�����E	W��, ��d�kR�KaˬI�K^��z7m7 6.�����,b;�ö-�DdShPeXn]+s#źI�
m�J:�[L�ؖU�Eq-���ͬ�䄧a�6n�/l�5d�N�o`ś���et�z"�1�˧�K�Zӑ乴�*b!�b����M����Wc1Ք����nl+i[Բ4�zL�&e�v�d��,dq�e��,h\��&�n��I�Y�Ɓ˖C
�Dq�l=H�����Ib�n�ې���i�RbOb

��ba��/!��]@�e=��zi��A��9Y���,�Mɸ�n�]h��Ì��C]c�&ǘ�;��B��{y*ӭ�R�P�t���׹���l� �ʴ�B�4�d��) !�s4�%	�,����{��6,��V�J��q&T�󡎪�� hm����
-�5j�GH��P�\%ɮ����\e��8�w*�gP��hטA��VR-+�n��eh b�@,}��`d�m<�wu(��t�PmLZ֨aN�V�u�6�6ոt�nMͅku���Y̤t/��|.E�lEn�LA2ʨ�ۼ[Z7t�\�*#�w`:��>Ue:n�݃�w*�����7�q��I����d������9�d�z/6��W{[a���+5�7�2h�)�W�͑���C�b���d�.�D�z�=�-����u60�y��g\���%m��v��Y�v�#$�o%G��n�H=h�/#��m^U�D"#Td	���ѺR�I�oS��h�^�@�ٚZ�`̡����b�Lh�+"Sh���9c�5En�Yw�S�LLn"�YXY�&�Dn�f`��@p]a�P=���*�Cŷn���i�����juk�k�ԯ+;�l�Z��ն�|.�`8Mʛr�އ�*�*��|�f��p�C6�Z����U��mY��7/u��ʤė�X3]:໭�v�@!�g�R_Z`4�%V��X-��q�Q��Ma�b�F0�l�*b�jΩIH^�Ц�^'�闖%bQ�6-7��G5Շ�Y&,�&n̬�VU���D � z�Û𤩪�X�YA(���ܢ���Wߠ�#c��(�&��(�
�#@K�PD�˷{J�w�fX�h�!g��"��lPT�,;q�(�K5�k�*�#X.1������m&�y�*�򶥧��� ����U]`�6�@{�L3�cx�Sٔ٭�ti�Q����!F����B=}O����f��V��M������h�F�QBCb�ː�2�/��qӓ)S�.�N1��MgE�#�K�x�S�@��Z�Jm��q�']Jb��j�^��*�Yt�fIQ(C�(��0�x��0͚�і���;�T�e���X��ÎT��]3 �sr�P�"9M�٬�Ŏ�d^T[B�|5L0�5�mhۙ��nBk�����T5�rP��k��.���BQ%�L�� �oi8� E=�㼂��k7H����aВ8�hӄ�k&a����Z�H�3(t���V0㬹���Ƕr�h��hɓ��CaA�ͣGA�A2��-����Ce_��bܶ�j�LR�ح�&��C-��6ا�GT������3s%H��k@�������>vt!�R�*]�b���N�^V�p`; ��Z�J��Pd�r7(�8)�����
&�Hk.`C�}*ڦBX�ٺ;Y+~�U�t��5$��e.���E2���ﭑZ�N5C
J�2N��Cm5a#%��Jܤ���(���ki�*�z�̸
<q["��wMe���,¡�Yr��hƙX�b6����&���wF��'\yCU�6��3(6����9��[D�jbb]�\����l��5{�P`����t��cڸ�l�n��I蠅a�����CT2�Ku���H�b�I	�j�H�0Gl���ݧ�Q7I�՘�+A��ݵ^�:�&[{��t�����n^vb�pKH�wq��u��sK3	4�x�k_�״j]Z�����s�B�nm'+B�[��$��Z�b*e��D�btX4��X�٣b�V-+�[�V@���Zҹ��{}6��P'�s�%	��,��+A����n�y1ǀ�D-8��+5� �P��X-�7F� WF�=�jAhP;��74<�����؊�l��e�m(�v�Y�%<ı��ʍL��җq-I�f�ȕ���ID�h:l�[���X����h��MVw'���qX]��V�]j�>ӣ.7�F�4n)#�q�D]�XOn����޺��r��(Db��s-P{�.�RaȎ�6�h���ٛHQϭ�ٯ�/X��JՉ��V$�*j�g+��֨%]�Z�l���w���H��a$ݚR���	�-;(�
���H�rɓ*rnj�Pm֒��̫�d��s��ʶ7R�����2����˰��):Ԛ5ۤ0��˓I�MJ�`�q��6���a��l�2՗J,��A���쬒1G@�w�;:t[:V��P�ə�/���e�E�v�qSx1Y
c�1c�.�5!c
#��IQU�������v��q:Yle�܌c���v�
uz������e6&d���\8 e�)Re0�hSR^pщ��悰�R��s)�YW��95��;I3��x�}�',�u�)�VBn�����c�N��Ȃ��b�r�՜sV�D[�:�q^�f+�b,J����Y��+p=*Heƨ!�NaJ͔���kc̳���楕|���*-��W���1�dWdf'��q�Krٓ*U��5�BbjT�koI��@j�EOF"�����R޵�:�ƈ��(H��um�`��eВQ9.�̆���u�+�K�ٱ^h�e�BɆ��i�.^,:�{P�{Nn��E ��l�r�����
�o)��[���%�wt��k87��̨�dr6���%+D��V�:ݾ�i��ǋl,d�&fE�T�m<�f�f�ې��Bm'Z�z���L�ܚ�Fb�P{a�yY[emHu�5FC�3Xk]ҙC�����XZ�z��l�ͬ�`�B��>ĳ!+R)�СS1�a�)y:�#����^Cn��!nEQ�H,1E�i���;N؀JD���7yn�x��Z�ˋ&�Q�uriqE{pV&SX�mЭ���h��߶6�r��K)�U�C�H^H��e`��Zʼ��6.�2@kA��vSN� 5�j4_s��8�pq���G2��r]���2��G[������0E�@�n�DVV\k��d�i�aU$�*Sڴ�h2^P���`�!�N�,�KFL-1kq�E���4�͂��SD�OHi��E{WL�Z� -I�X6�U��D
���X뮬v:ldDH�,b�T��-�M4��	��Ɗ[��4�YZ�H"!�o��))xp���k�X嘒��T%�;pH�j�ޟ���Z�s�����L�u�=j���9R�X����C*(���C���ũ�ɲ�&.V�"Nm����)�6�� 0d�J����Y��޵j��rV��i����I4�r*�@=Օ�K֋�YK{P���/y��Zu�#̳W.�O'ĶÃW�*���E��C�U)� `�%X�"�	P��WS+q]Y��X���׳Z�7r��d6i��b��V��*O�)t����ۺݡa˿�؀73]o�DtK���K�`T�!g�4kT�^����/3©�Mn9�N��2�M�r�O��!ö.�i�&�0:�Ѯѩ3/$j<���e�-�۸���v6��{5��)F�M�e]�3�͒���oo\�Ʊ�i�*ݡ0��1a������ii�%AxcǂPt⛀��J�4�C#��n���	R���j��R��8�9�ur=Tw	h�b�h9,�V�7��҉{��ݭSvq1y�)l���j���sD���i�F����d�U�������r���,�ʅ�ERE�s6Zwf܏"��Yx�{��v������r
���F��4�SN坢�Z =F�76�a�2��٣[����t�[�	4޺�M7�����R0��+sh�/sFY�&�vPYv��1'{�0�f���fS##�.T����6�[lh�!g{N��{�3i=�¹.�]h�2��I۽f.X,�h��e4i�պ-U%cQ�gpu��عH�DW��X٤fn��j5a���n�^�3F�+sQ����D�K�c96�ޙ��&6.l����/�u�[�-9|$�2ntsb�I*�R��1�`�BƜO!r�� }��9}P�b·z� �n��47�Kersy\jk;r:=E`�c��sT��"�*�鸃[�]n�?#r��g3Yi+�!�>M��B�Ɔ\�Gk������rr�I��C��ƫ>�j��<��t_TQ|�S��V�Yi��1�����G7��4K���}�{S�󡍅ѫ@�TW�e�p؛٫1�
�Zšm�f"8�8�i�����&�*N���[L���K�W�3H�*WY�v��
���r��[	�ט�p�ιNr}�˲mMR�ެ8��4![���,��k~�$#�w���L��!��-�^��e�F�]t�Gf����@���P���I)�G.:��`\�X��!��'�,1����N�{�W���&�RH}�����OWes]*'
啕��o

����8MH�΃�5�b����;�ކ�����n���$���Syb����Մ�Y���]�E�׺�od���%Nvv�G�3�D9n�����x(�8�G�����[̧z#b���-U�j���K�b��LD�6�
\2�>
����zA��6�9a�\)d$n]P�t�J����	v;�Yة�s�Ӏ���A���#�emص5���4U�lX<C��6��y�2i�.RLQ���p�}��g�G:05���l�!GC�즛��ڀ�H�YO�i�j�+m��Y*U���>�x��5gSŝL�g�E�m�^�VZEד�2�-3��^]��
�v�2�Ħ
�]�u���n�ۗ f����Cb��Z���MB^��5�"�]�g�@���n��i�pd��m�r�ݕ��*�iRf����y���Ł��%��m�uċƘr��&L7�v��s*=+&���7|���3�����G��@%�|L o7�f�]�zt#b��@n���+�8��'=y]�:ڄ"^T���l���s�l�u	�9�i��mbb�w�A�y�sI�(|,b6�%�mw�o�Ki��_\wnF"�;��Z�b��meUۡP�.E�zv��n8��E��,���zeq�v��:���a�]-|��'q�32�;��psro`sy,6;o5�]Ϻ�my��K���sn�Bu>��]�Z2���N�Ce��"vpP��l��d���F��e=��ޝ�z��/���NA}J����)�N�hk�L���i�r��K(X�R��XЩ�X�k
�KҔT,�챢8�Y�����*]j��S�)�zI�HUmΖ��b� �>t14y0��]Ղ2�!���ΐX�W�w���
�oL*`�Pu�������l�S)J�{��(W3�;\e��{7�As��S�._N�D�mF�4^���0i݁�`ӑUl�y����*ʺ'��)�n��2g<�'kQˊ<{u��a)7�I�H�s�6�@��4�25Q��Wv����Ҏѝ���v����+��Vj��1+-�P�����WA�I�ް@�X7�BtꏧD㜶V<�dY2M���lCM2B�1�ϳ��)4Cm���L�T[ؓw;�a2���t��`5*�֢�QEIdQ�ھڏ�CR�a.^� 9��TT�IK� nq	P��&�RvR�M�v@AG�s{*�5*b�;Y�Uct�����9�$K�s!v�^��<�;�Q�l�t����`��U���|���;e�}:No�*>�y�?:�!h�W"�gG(�Ʊʻ���[F�}Bt�G�d\})b��T�m�}!�w�����k����7+�CV^��ͤ�b�ˑ����Y��,�
�5-'��AԐd��@E��(fQ̜l��4����P���T��=�8��@9n�lY'����	�S�WVM�< ����t�8]�i�k����SY��6j.C�����{�!xwt��hk��M�r�ޑQ쫀m�;�Sڿ��ھ˕>���3��fj�-�Qs�	!|���۽o5A��i���EX8w�����Y�<�R%kpy�Q�ѭ[]�K����+X�i�JcE0X��9���>۫l�+i'�̭�_`��-�Uc{.� L��nzJR�\W�A�j���ی��3:�tWƊ=��N[=Wyr����[�wz�Vp꾿��6Q0C���$����ŽtGe��q<��ː�b��N�8FT��]�"�BE���/z��$(��7�⫆ֹ�qa���۫0�,I���7��L۰�b���%v��z�4��Tg|�t)d'P�v��O=�̉���c$�I�V�D�)�׼�cy��թ��Ϥ!"��֓�(l�����1cz{�z�;�/]�X+tL��v�K����h5N���r�#����śƞ-�������2Jr���Cvtt^C[A�'S.�p'���)�p�Fol�I�9t�gB�;]jaʝW�L�%����m̩�SzVk�B�Z����\z�p�M�����xYJ�4Z��xVh.�7]��9Z6���@�HU����K��|������u�-�')Z���λ�=y=Z�B�](댗�T�9qV�>�_,���tD�k�;�ذ�(�W"y��nʶ/0Gۡ�)+��xi3���Jkt~4V�*�P^�\�o�gޖR�+:n�LXKZ�&j��Ug_F(>b�E�1�)	���C*�N����,�[�ک�����rB��,�]/��*5��*o��SJȔ�oe��[�؝|�]�ui�M�혛1��U��I�l�d!��
�y9)ٶ3Nu��r%op�}l��\���杌��^�-mf2m�+vpWse�Ͷ�T��,b��m��:l����mu�w���6zL��=�u���S�����G���ܑ������,���NQ娮+[�z���d�@o �8�b����S�k9f]��%Zw-%�V�F��1�;x\1c7w
�LT׺WH�S_n��x�ҝ�w��V�])l`S�TU��j�������b;�U��e�[&��3	��:[j,��5 ���f���L�T���k�um��ϛ�0�QX�|��.���1&Ԯ:@�f-utIk<�m��WD����_�>�.�A��i�-(�gM�֡1��}��77gj��P����cd2��wM��+EnX�z%�� ���*�V�|9qѵ"�5���=y1�mQ�3cNn�'���Q�̭��"�q��բ�Dv��ڎ�m��+��ptnW��J��Ff��E���ԋy�΁i��}����Y��*��Aκ��82K2��ܦ��ϳX14��-
�� q�u���]��;7z�$�r>gc ������	ݻ��V��6�4���惨�wה�N' �[�m���\3��:�L3���P��Hu.�ɘ��5��A��8:JL�n�ƛ��ᆈn�]ܾ{�Dh�x�3C�M`��0��hn��s���ڍr9!����k� �=3��^E0lnЍ@�.`�ok�
ԕ�̤�t+ʃk��K��9:��xG*��Z썒�&9�V�A�4���J�Q�Cl�Z�;�7&p�;�m���g��=.[�/�x���l\ZN�����o#�I�GU����(~ՁCٶ�p+S z8��nȧ���8�j�^��eǽo�5�1�fc�˸m���R2Gn�8	���(mh���$��M���k��s-1q�F~��U�]C�����A�:0��4���I����t�o\���%�=W�"�x{�E|��UZ�h��,�`��R64�K|):�}�Z�h�4��LɰVzN�s�Hw���`2��- ���]�Q�H�˫�)^1��Ú���I�ڙ}z&TK�٤fzg;u;�TnnX�S��!Ҹ&�Wlb��gG6�F��RɌG����k̭�
�3�����)O{��:Y#͕�Q�ۜ,�
�t�y��eJ���.�h:Vk]�qN<�\*E�:a7EN��n��X�����+�m��J������q�v �,Yx�&��kw��wu 魆�Z�x�'a6x(����%im���ˏfCǒ��c����Ν�bݕ���]��8e+�Rc�� e8������P���P��<�V���1/'-k�.j�`d�o��;n���lv�䬭Z��NU�����j E�z���v�ѡ7�6�O?I�������g�v�)KUk5�3do7��L���uY�� �c6�KwGa�m��s�i�6�ǁ)S�r���ua�q;y{Ɉ.��M`8i�Ƹ9��C$�ޜl���X��T�Y��GQ躟�wW��m���ǽ��-�v�Ǧi�c���`VS���S�W��]bڦ{h�S�C�w��v�g7k��
�Q�b�r��[h�����z�7S3�w8��G�>L�J� �$�%��Ĝ!�����Yƈ�+���y�Y`e��r��a�*���<�G"�Q�cC�L�|��Wh�ۢѡGo��*Ү����]�]�yP���
;g�-ʺ&���:-�![ͮ�[ى�/8��z�Yɰt|;�,@��I���{��}&�0��C-ȥ��s��sX�N���]��`�5R/q�f�:��1��=�2uԽ)�]E��K��`U2��;��b	5%��׬�5�ʸ�ӕ�s�:����}Ԗ܏:D(@��t[7۝GG['C�� �`pm��(�ې�6�2���۷��?d�J�@�ˌw��]F¡}��Zk�f�́0��F�lg��zێM�Gs)<�]ΰ}xbЅd}]���r�T����|ek�N��)�/�!��N�D,b�*�b}ȵֵG�^Q��Ą��U�Z,ڄ�R��қ�H؏��)d{Gl1i��\�M������[�`+���;�4��!��n��ұ}�Z���eZ�}w�FC(�>��v�BȊ�S��G���Dn�Ά`�4pt��Y@��#���A-��2`�MQ٠t�f�n�̭1���$��'�n�/���$V��KFjlT�Z3�b6�ȁz�ѧ%턖��{��D�m��:ZJ���坕� ��Q)��(��W�L�;6��݊b�5�ܭɒ���>(d�̤o��G���p����;BY��m͕r}y��<��f��Ȓ�m�
`����罻.?�;6l�{��Qu��W��K��}y!9Mv�V�{bɮ�����Ռ��2�֓�y����z����l�a�Ҵ�#�)���]��kAU��N^݉�\�V�в ���7�S�<{4��@{�g3��F@�8/5,vP��'�B�rZ��N�c�w[�KL����P�sz�:�x�<�Y�/f-�u�Z3��j�![�ۜ"��$�W/���Q�T�������6�-��3F����]�����s�Z���+N:e�\�t�U� Ue46�v@EX'�&�|�w�eX�*l���ya�)CNrw����ۢ�s����Б"�V�"��a�{]C*S�����P�7\
�v�})⼻`A�6P�]���,�+H ���K�l�5��L������1�|M��+�J˼��1�:�R�)����ÇM\�%�y���I%ֺ
+Ӽ�y8�8.>��A��;����i�*�m���^��A��T{�ߓ�&�3x�jܩ�(�+`r�����sf.��v�㹭m� Г]�-;)��k��lQ���LJ۬T�jY���e)���L��3��?(sfU�|��`1�ǃvһ獧׌�r�bo��aT�J� :�J�ZV�-��
��AY�q�s���i�i9�IceJ��l�Eocֱ%���y5���ތU�{i��1���h<t�#�Ԯ�}�-e�&���fݜtUo$���E^�i�XԾ_qOT��v�s6�\�c0}1ԔnM�V�r�]-[���-�ee�<���޶�K�o-tY ����X��]ٕ31f���`m����%o�N����54�.R���,�o��/�T���/m=5�N�Oej��j�Rި콴�ņ-�j�^���{���Y\2�M��]�muI�q:f̃Ì[�r�8d��ݢХ���5T]	�[4/�޷��e� �ok�*�	ݨV0wb��@M��c�m��K�ɶ�+GS�k�u6�淪U�b۸8vZ��3l����[Z%H7�>K�2!@w^�n������c�Y�1Ι�V�f�y�+�|�7|��9��"n�o+n���V�v���Rb�έ�i`��t����(��fC�k�|(��t�U�����c�5*E��:�б���M����X����꽡c@��wR���WO4	[�K5��).|2on�Wmы8��z�9w/jis��Y>A_
���&��W��i������r���˘�΢�2�L�O�u9���\&�'�����ِͭ�Ĺ���sbT�������qY���J�n�V�f-Q3���@ne!%GP9��+:����j��7�ޑbEYY������$���x��{��<��X�9�j�% }�)����Q�ʒ��ZO;���e���\7[��V�#Q_B�t��H��.c���2��j���`Qt�X��H���i*���:���C�C���0P�ѫ�ў�Qw��ed�$�آ^LĬG9a�ȳ;g�P���lR�'@]|'B@
-̖����K鍚�瓭Rr��Ip�VO/f�2ƒ5�J��J�u$ͅ�Ķ��ET��/�l��M[���kK���
aU�֩A�v�kx˓���}�%2���f��]�u��u)��&�7�ԡMf��gb���Qn��ok���s'�򿓒16c|�j�a6��%#dok����K��h���i/�*z&��Ӈ�;�������/qWj[M�lJ������)�M9�Yӈ���Gf���-�4��՗zq.|���Sw�.��uU�}��}�}�g���_G���z�C���aR� +���Wؒ���ؒ�Gu��x�A�w��c�Z�H�Gu�,�`�N �n�c��kWF�9���-|�#	�)P8�Z��-��j�Y�V�6�*��j�7i��Z�|��C �CZ��o�N�)��w�mܳb��\����c�R�
峢��x��O�sfGB�rZ�z #����2��f��nV����}jF�e��Ɲ<�i�HlكF�ڝw��vy���SwX����M�4�'�.�v�V�e� aq�P���G]^�=a�&�]fe���)8rN�9�+��7K8�s��f.e��u��|�N���f�L>�ʆ�tz�K�1r�&�R�YIm!�%_f�{�QT���>ܤ��#ڃ9.�Rb: ����{�><�I.��-�xB�o4�T�յn�353�7mn2U����|���v]�W�`wY�����e��8��7q*y�fp4�#�!l��1)kdf�nt�$���Dk>*����ݧϕ�Au�_H�f��kE�VRp=D�m`4��7J5+&�Kc%���{���gU��j�|��JQ�ˌm���4@��V%��j졘��[mx�������la��P�#pU�
	ҽ:`K��ܫӎ�s��5���e�F��j�vZ.�t�CfM�v��3z�@�㔢]Ъ�r��z��Y�D2k̫w����h��{���.�����cھ[t+j)����ާe$��H#̛g_q]�1�jF�Kl�Iݫ��n���9֔������(%�����ٌ����}�M��9ٔ��VҮ�ΟtN�CO6���	��؝�A=ّ�
��/z
Mʃf����d�U�j����w����N�k�M��U���)g�����b�%Q/	��g#H�(��C%e�r�C�yt�r�c�.�����E�U83Ѵ-�~7��>���Or�8�tG����͔2i-��}v	�Mt��M���H�}�$�e�Au���%�#��Ӹ�.N���1o�K�qU���+{\�R+
wW�A�;�]�����t�'�T-�[�7MG*�K]r�9jp�wwF��~v���@�cRx��*`��@���AG�ɹYKh��l�������y�6Z_L�|�uN�k��E�Y�]t!jz�y-���k=anp� �����d;u��=�܄yԺ����/�rf���[��k��s������/D���A��v��Y��ѱ�$�=(qaA�ȹ�R�30 �q�ƶ�����M��g%^��7�t��������M�����}*B�9�Y[��<�F�yڗ���_fHy�6w*�#5�!�SRf�L����Y|�cZ�Z��R��&�I���%۷G(��y�R�w����&�k��11�s\,me�K�Aq�]W�';$n�D�ʕ����˝�� ��9&�K�N�s;!�q�>z�Ժw��[q���v3��ԅav	�裭>޳��"be����I���FZ��e��G7��<o7�6k�%>�QER�q�{mm8��wK���.=I�&��5P	o��u�mrŐR�W_%�v���sl���4q�������T(�=*�y���;;;��Aq5V8J�kJ�2mg^����:��hZ͡� ����JW�톺�	 ��:�yZ�e�9�w���ҽmV��������]щ2����X�kJyi���ٓ���I��k{V�Ji0	��[�%쫝bӣ3�}��n��\e�N�F����ŝ�4/m���ܛ�]]���˜��93TP�;GS闛yĘ���$��|i���nt@@,!nr ��ACrmd��(.�ŕ�XU���^$� �t��X�|�[�Lq�Sr����enk�4�N�`��G��ۛyO�^������aC{����S(�j�ñ�'�AԚ�-���ޛ}�NY__9����T�������_J鼖��$}�)]X�ȍ,�"��x�Ѕ\�r�%�t���E���i]�n��U����?t�'Å�W���JJ���*�;w��R��ZзFv�Z�޹�H�����������w���ӧ����Ժ���t�ȗg�F�_>�9-[�9�n��KYB��h�c&0�݂ך�Dw&����lA��c��W�6�b��9� 3�7�֢�j`�j[I}��57rv.���.�,��vڷb�6�R�V��s���4w^��r˘k�V�.���/�m0�i�;�y�ѐ�1wj������fh�mn�x"���&�f��ܕu��g�-٩�\C���c1�={ݣ�#�cBw�6���⎷��u��R�S{��(*���Y��-�w��m�Rҿ�l����!��W�@�w�
�]�GB��v� ׫e�	�G���t*8/���+f�[u(,{��6�oX,��ۍ�n����b�lR�+�H�BeJt�N�l<��(��ʅ��`P��Q�l�|����͕�J�:C
d,:�a<�s[CzwPB��]W6�w�f�m�u�FSl� -;�"��w���*^�F]�Y]�y&U��ӽ5�n��`G+\�����4���s��
�I�0)��T��.i�桎�R#�[�u1��E��6�ѝ݁ ����R��6�fP����M-�o�C�x��Ґe�a,�6�)�N��N��)wwSt�nH�,w`�;��{���]h�{Q;@�����p\D�̣j�'.��uI��Nm�	�eaC#�7{>�iʂ�>���/���hT��Ǳ��e��b��rK�T���bcy�����F���
��Ō�����{(�_<z���IVS�k:�l�H����Ņ�s������ ��tC��	��9O�;�:�Q�}�nH���=W8�G�7.�������T�"|����ܬ��d;���f��x8�v�pX'�K�xf07�Q���d'��޾��t��������bu4ϞXU�u�����}�#�1۹�,N�Q�F�r�Z �;��*yp=���-r�ۊ��xYW�hʴ
�2�� �l���n��̖!w�db�P������ަ:K�V�wN�јshlʋE�準��V�έy)l�
5lq��[{��n���������]F�]�G=1��1Ʒ
Nbu�fngI�+ӡ�T�5lJ���g�g��A�0��@:�γ����&m�	��4��T*S��2n:�C���%���M+:��銤�W3.�rL�ƅ���xc`��:�g3��q�	ͤ���g
�7�@����X���Z9JW�hq�S���7�"n�.�3r`��b[�h�[µ��T�Ү��R�p7ծt\P�ь݌��R��Ne�|UvNr�(l�ˑn�帥ȳ��
�2u�%[ɧq��T����&��p����|���[叒oN��q!{oc�A'D,����ƻgX+.���
����)��i]�C����oZ��R�lC�4�$��4ԗӨ���97�w,!D4��۹t�t�� �oe��=3�����P9kSBp9�,�*·\
՛/u=��X�ga��u]f����#�s]�n �|�w>jv�����z������6)�n�����.^��	7�du��X��vˈ����Ҝ�B���,�ٱSj1�=�Vv�G��9®��Ml�aі���*Ҏ����
z���d�]�n���e�':=��� �xEjV23��X���[����=�b�K;HW%�t{)�	/��nV��=�X��f��g��Y�\|1�������!3B�.�61��|8�F�PK/7z�u�ܬ�7�������Z%�aB*��;��]�m�6�@u�e �������n����DPN��n�����`���%F��k����,f�������:��/U�*)�K�`�ñP�P9uҧ��hdCh偶�{x�o�����S�5�ܤ�؋�ړ��1��x��b<D	���j�oX�V��-�_0�H�`��m3@)Ɛ�����ig_6�������[9�SPaG�_N��Ҏr�B39�y�����@��Db�P6�w�=�U���Ĭ�ޱ/JQ Z�ŕu��R�)��5*#:ˍv���h#Rѱ��������B�" ���[�%c�[�3�ش@C��x~���褶�݊�l��(��6��r���E.��i%����v��ݣ�����n�W�8�"�j��Mȱmm|��s1u*��$�ukhulho6]�����vt,`zi�WpU�Z��\�3�mw�s&SԨ�]i���V�Y	���*:p ��\��T�)�i�1�<�ynȭ��f��1�+��@5�=v�Mk]�c�i3�rLq!�y
��a�&㸦�5�艵%�V����f�,{���'���ED�Z9u���u5Q�)�#fK7��XV��6v��л�d��dڐXl=ዃ�����Ok���d�ݧ͔F7���WH�Γc;���r��n��mK�B��W)*`�
x�#��g9�[�Qmu$+�,��7�(]��vP5aӊ2X�J���w9>�8��!�h��՚Q\�MJ�x�zХ������P ���r��m��o�N��t�t��%>�:��5M}4��󻽾�C�n�N�i:��M}�	Q;���y��߅2j�:6�q��F��LXVi��o;�ۦ�Ec��eU9�Hi��b����̏��x�w	l���6��#ֵ͝�c�Ap�����qB�\�‣�H�%�.�lȝww�bۛ�.&t�ù���G�{�י'�g.n�̂ۡ@䂍��(#�$���i�"i��IV 5�^Y#�@�n�/���T�R�Ѝ��6�r��]7nb�/������pB�d��$V��76�����j�� ����A4�e�I��mMfié}���32�'.�>����Z�ǭ�Ҹ:=�Z�|h�%��b��֪5�`Ǣ��FZ����ΰ@�@Q!�;��R��a`���8���ش1��Y/�#tO3Ris��t"u:au ��H8 7�:��`�<)�-��, u(�u��]��+�v��p�t�Fu9R�w3�KtT��t YS�'���99��W	;q�j�=��9���5YqB��-�j��ʸ[ Av����+��f�fˮ��m���%���vrM��ouWe�Y]&��d��� ;�sD��P�C}�VR��Xv�M:*6���d�Kwq��7��řq4I!T��p�q�V��UjՑ���(��H��\#7������NUx
���v�ͻ0%$ΣԻD�لot.�b��͗�jZ �#�7��P)��R�s�.�Y�/��EҼ�V`�2�'�oz	��5�[`
�%�ܴA�,IԶ�.|q����řC��N���{;+�e`�Bʹ�l���e�W�:���rڱ�n��E.fR�%�H�ٖ����WtNՊx���ӵSrB�
�2u^�-�&�
ѷg5��u��F�Br�HSUp�f�N����:ĉ��3����kJt��A�Q���� [���s\�{pP��޾���SY�s��*߫Q��9I3�������6���Lőp�V����q"N�(Un��U�ժt]��v!o�hS�Xի%u �h-f�.d�A�gP��]�Sh�.�m=%s���B�X�`v��I3e��[�k6����dr%+�k�L��b�(Z{��MD�]�ok6�Sd*-���2�=0MVš)�:Z`�]��Z�X*X���w:���Z/:�2e
c��%�De�1�>ˠ�����}�e6���V7w�*b��	���֌�h�4x��|������\W��E[�"Bu���tvG%"�:ɶ!���e�9\���ؖ6H���.�7��l�cC���K5�m_c4s��p�U1����z+��,'׎c5���W'�Sy׵b�ö��5f&�B��\�:�Q�K7s7u���J��6�Wp���Y�\A�ۖ���c�;����t1:�Y��[���s6#3f�Ľ��(s�V�t��5��r� Ah�Cr�+D
��\6�ޡ��(R����[��X���S�3�S/����j�Imm�nk���N(�ȇ�;1R"v٫r�E��ʎ'aNɼկ���!�[-��	C��V9Pg�ݟ�*�+�s�[RKJ�4��Ա>]X�����u��|�׆��m�Cb!Fd��a,.mdw�p<�֊3T�v�p�TE���V)����|�4jڲ`��}�nu�(2,���PTsa���P���C/����Ti:�.��V���t*�hC5I���-n7���Au3��}����T�]4�[����}�h��vnA>�0�qݧ���_T&�����z��tS���T�VJ�Js`�n��ѳ��Qc���)�\��Ι�k�ce��v�,�'RŒ�z�bZ��a9:�B^�/�кeG�p�.G��:��kz�p:/�M���rm���=Ctz_>
�@��E*�{)Y�'M�f��P�)��t6��ʡ�>o��[z�V���i5fĄlk�l�������b��/�`J� ���Y��lvme�R���Yz���d��������c�(F����qK�s0���P�F��ي�$s�=s�yt�&�c�P���&ᅼ�{�j챎���D�;��)��A"-��o��)�J�2�֣L�X�=H�b��cm�N��
 �y��C)�٠���v�z�M�2йp[=c�������,;%���,���r���v�OA3�6r郧3�uW�T�"+I[nIu�v	�F!�x_T Y�{|.ng_;���L�p{u�j�"�5xu즴T� 4���i�/ ב8�<��N�%\Rϭ��u��qb@b�X���[>����}�W��}���7�7�$��2ytUƀUs9�S�ݚ��R�CN/����x�s���n��Ž�&Na������`�m��E��m69{[��W\��o%�듡�����Ƣ��<�p���m�K�����C��$�p��R�]�b�;�^U��2sf�ȫw�n�F���^I��sUbJF��̩\�/�֕@��+��� ��-P�����&��9c�rJ�ßvb�O���1}�oV�f�uYeM"K ����U���7���W$:J������<��a|��]oddv�H���&�P��+�FlBj��\<����D���u2-�Y�w���R�;��c���Iŕu��4�qV�s*%·#o������ �ܖ)�R��^�e�*�g�|s%C|zuo^��h��'�;4q��m��k2_��Ti�ݗʶ�b)s.N%�e�W����6ȓq��U4S���ؠ�V�t�]����spj��.N3�U��(�3��/�3zc�i�d]1�c����x���ƳH�Èk�ǺĹ2����V��7w	=�:j!m���SUb�Jbf�1�P���8ީ)N�������;!J���*:3e1�JV��iғ�^q:���kR����T'8kJp��<�wU�p$u���ݖ�1x-���n�.fC�i����r��t�@Ls;�޾{�ͅ����j�P���6�
Q�)2 �����y�f�FDDT��e�:��!���X{��P)Q2.Pn�"�	�IHL�Y��WM,(-(ȋ6Bd&r4CCD���dsE)�븉�2�B���1H���,%M�
��Ԋ�L�,�v��"e[(-Z�GR�TH�̭U"�CB0���D��ԝr�PW��E�$/u�:ia���:�U����!���+T�-���&i!´u**��s�;�#���*�jʂ���8�E��I9���"h�'TB#.Y)�%�,[REM�\�P������V��E�C=�i�ʬ�t�#D�;��R)Ԉ���ME6\�J�!*�&�a9�=�D�`K(R�D�G1r�<��.xy�Nl��!̳)&����$�fW$4(�D0ڨ,�5�¬���D�@�@���˝e�t�[+�p;}]�)8;78-HLٴ��%s]���N��X�ء������Lcw�e���h_�X�!�Mu_�Q�E��.��Bj�8�pŘ�
��P�.�h����k�%�	�D���c�@EGˋ?	��OP?-#.s��}T5�VZ�]O�pw�A�	**�)i�t�΀to��A�N�SRm.�^�k�]_s�[�˦�IҵA!y�z��rԺ���)���l߷�a鋈��^'LOdmFᯓ��8n8�+��W���]f���ѭf�R�O3,��rQ9x��j���E��֢�Ofܜ���i(K��ۭ�8��o�ӞP�I�����S���� 8?�� �/��"��y��T��w_n���7T,�{��U�3���}�k'��8Kvg��PX�5�)uƚ��^ �<Դ򘅆7������iJ]�4&���Cv֒t�<r���F�� ��\l{=��=��_��^�.�^?N�LźT���+���&%���P�B��G�,r;�K8)����]jZ�6'7kt�R|s�?1���M2��lj8 ���Ot5C׳T�pu�;�>x%�;娏!�[���;C�L�Ɯ[Z�a����;�j끄�v����I�K��x
{K�;�mz���3b�|�c�M�e��t �g���@�}wZ峣��n<��������m(��K���Bb��aU�1\�έ�'g$��oq�'Z\~�c̐dSu������<�ê2X�*]B7�� uwi��q��s��䯽Ϥ��
p �-�X:P���2[W��h�]�������B����'�a`�L�azt�A����9�P����gTaG&�-�'�("y鼻�ɻ�v6%f�򅖀�Yf11� �(��;������ϔ�)Hk�'��T�o�٧{��\����/����?���|��Y��ڰ<����o�B�p�Ӌ9�^�$c^���}��Q��_��p۠9�uCo��,	�zF#"~H��6�t��e?�}�{�km{�t�U�4�W>����ܨS��!a諽5V�vֈ����E݌���}��^xS�-,0
U!���r�����Fjt��s�{z,7�S��;��f�`�m���E��j�����H+#]��gR e��2΃qΟ9��4;�I�Ԇ�)gj�(R�[�K�˺�m-'vʮ�Ϲ���j�:G�L p.t�.��Xx���^�옔V�up�Br��jA�nWJ�k�Q�s��Y]H��z�A���(g��1� 7�[sZ����\�A�K���'`��eʲx����rm��'o:��1��+�S�{�h�Ëe��b_j�v��!]�}��8^ev���2�.|v�$�}v���\"�k+��Ul���d��'����|��T�W�(O��������8�/�sPt �z�[��a�3;Π���w��H�<�%�����,�lS��k��['�%��+��;����Ø�6��V|���q�H����� ���>U��Q��M���&��e�%�=����;c�p�Q�`#�	��ئ���@��,dc/�)o%
�: ��$a�0_Wv!"�T���SF5�g:��`�%0w�d�}m�[���ލb�C�ޟ�Á1*��2�"��V'�r������x��U������-���Z�jJ� [SA	D�9� �H��R��Z^`����� ���d�O`���{��s7K�ӂ9�`)��;�uV"j�(t��@�4&xEDIZpgȚӵ,B��L�D�d*��|�_Q|x��}N�f4B ��K�6�V�&�att��n�|�Z+-셪f℈��a�)zoyT�nxT��杚6��k�1Q����:������pW;$@��mM�a��Yļ��g1�ܩw���L��ۦ/ P�%��a�����*�N� )nV���RX�KS;l/	)$�v�;�����z�a
#v���9�KOU�t�.u�ya�2S�.fZG_CEd����DYɓVE���\�v��Z�~��	���r���p!��w����p�L�r��}��w�\Ŭ�PnE�͏UC �p���Re�n]{�[-]q�-W*�"ֺԒ�n8&po9�7�NR��ȱR�#y�"/������P�(���.���{��c���8�4c�vA��m�0bq����wR�C}?d�n�~�B�2���0h~2���T���]%��	m���*���^�s�8��'��\5Y���1��I×(e@���<����K=Yky�gC�#\�(�j"w�&X;鲳�\cvӽ�W�o�V*C��c�π���q��䧆`� �,I< �ތ3A�F�QC�"Ӗ�e:��&Fq���ivd��PyaN/�(��E�Y�!����R�L���)S"7�V��a_c��X�l�mm916MZ�@&���!C�+L�>0��V�p�r,�?TAI��`�fk�8n�s�����?M`=8�H������4JD�;%!LD�a#��aq�X�w�b�$�Ѽ�O�ӷ蒭��>�9�5^��u��V�T\.��st7Ȳ�����r�X���1��hv��e�6f���(�Gy_>�z���pnL�r�̾5{���y3X�voE!Y���ё!y%��T�n	�M����Y��uޭ��j�.Q^���7$�����v��1�S Ft[vFK�Fv�": ��27&}zH�h��(���!�.�V�1���vJvـ+JE1�)7Pr��2.�F��RDu�V=|`p��Zw-IҴ#;S�W�xu���s��pϋj� E"WC5�LCv�$���� 22˾a(�y)Ų_L��Ļ1Rt95Eq����q�\�!����S%���YSȡ�i�魃��{�wS\>@8�* �:F?��C�R�ڳ���\*G]qQ�����]���{�轵7��7����$	T�4�@SCn�?	�d���f��9�B�������u]R�p�w=���+�+���ؑ�3��mI��pa��,��2~U7Le�[��_-��@b�}��%zB�6��������W3�ꘞ�ڍ�I�`�7Y5�^��:�.�7���`~=�dH���=G�y���Ʋ�T�"Ժ�{S�	g;�~ڹ�'6ڻ}1u�����2�Z
�<�������� �u�E��φC�l�}��Ҧ�Β;;k�w%����'��p,u��z�DfM�vy��M|0(Ǭ*���`+���ZQ��'5Jg.�/��)�n�2����n9yzp��[�=êC�{�;Hѭ�v�v���@`��(T�W㐠�[DR&�WLҤ�g�.��%@�Ȝ�g�Ƶ�t�N3'_����V�% ~��'�DR�^���`@���]� C^R���t����u\ �X��Khm�kI:]#<Y\�#^��(�F*�ha �s���U���o��l�Dpyq���:Tƕu�/�a���$��1�-����Wy|�����I�
��K��E��4&���#��_1����B�Ͳ�P(� h`K�h*Mw�����'6�֒�W����)M�Ơ�x`�z�#��F���>Ƽ�u�h��4m��r�c�>ad��}�d�� l@ �|:P�Nx`�m_�졸�w��/pl�J�m�n2J3cN�=�U?8F�d@}y�Q��Xꄮ#U�+�V�nQ1w*C9l�`�[�y���\cU�Z�yP񬆀�]D%��ͳ��/��3թ�M)+k#�Oc�x�d��H�0�B�N���S�g����A��LYכ�x,0��a������3T��.-��S:O2h�6�y���,	��G����bË��^K7@N{j�T��̀�ݰ�nERJR~��t�*��ᝇ)��n+�l����<j�ۋƣ���Žq��߈���d�#����L������:�c�%K�ԹI���vӗ��96�H�)�����~⤗��udu1��o賰�]!{��|u��m�r��Om���M3�4��CTp͛� wx�WYA�կ6�޹������Թ�*p�QJp���'��١�R��5:���a����X��ys�|�:�g[K�VΘ!9�+�C0ײ��ic��%��y�����s��c7ml��k��1IZ�%�:-�W�n�E�'v��,4Z����Bd�D��ˬ��s9��\�`}Ztj�q2������E��]y�W*��"+ph�	���ω�`���ȸ�L�Iȹ�֔������2�^_�+>��n���d-W��@A�'G]�gE��|��i ٝ�;���yq��ֺ4�`��g�9l����l�|j�����Ǽټ}:nL!X��jO�D1Q3��꧹NDZ��k�>�P�X�j��B��~cB��wΦ�ҁ�P�PqeU|e�0
�E0�D�Tu݈H(�c���5�ìgod�)R3/;zV��Q7n��@�(�V�EWPT{��<��O��.��z�
3�>6=
x�>��"'�2S�Z���Ub����:�lM�^1��^�]p�+|x�$���8'5�6�;y/�Q*8�`0|7}��<{D��}9��M��� ��<vޑ��)M�c���1K�V����ُ�U����&o��\OM�J̳��E'<�8w�*���9�2��&��S� �`��*�nZ^d	�q��Ng4�g�}�UjD���C4��o*�C6!����nw�_Ϊ�J$�2:��� 	�p���V��>�OG�2�Xly,q��'1�����Kς��:�Hv`��MG�?l�x�;ُ��&���X�[f�Ça�Η��yԇ9�Rc�th�s����.+] t���l_�[ ��jz����W�S��U-�@�	}x�[������"�S4ܰ	���'�:��׮c�!����JA��]H5(��0��N����r(�wi2�P�ULC�ZU�]VM�)���t,]�tY�
�~�j��3t�x	V��2�f*�T�4n�`��2���r$�TOGw$�*��2wI�,C�`ۅ�������8��+*��P'j]A�Pw�5ۋ��4�;k�B��d,�;�	����SC�
�V[�D�=s�=�4�����޼S��e��Ԗ3���$WZ��j"cy�e��[<��ݸN��Ӏ0���KNp+z�eF~�w.V��k�] ,�O�(�z_H�n)��{)��R�Mz4!�m[��4N`ɻ�NV�`��_N��:�1���72� ��������o����f���&���~�@��pΩ�"�U�J�B�'�j_h���.e���"�\�{���J�����i�g�)��T �EV�Y5gd���O�1[ia���Q��*����JCm�
�|خ��-[����9���S�WwD�֨H�=����x.�d�i$�~��L�A�b�v|;D�����Jhw={5���\ۘz<ٸ)w�����Z��>��ϐbh�
�*�<;����s:�������ԁZ��w;���X�6\��!96ۢ/iգ6�A��ɐ^�{��Xmt�z�y���ztE����b�����c	�)�X��7Pr�۾�sGq�^k��m���Rl�����hK0���a_�q�+�[amYg	�D�f��\�����!(�bv���FW��^��!_�7���A�U!�{3�橒�5�����*X)�$R�7@$�W��B�'�RvN��+�tȆ.w2���y��ő�"��n2\�����h��)�`iyM(�3���>ZE�b)��;�lWK��9�c����+7R#*��Nא���D�m-N�n�|i�����]Kj����V�M�R�&��� �fZ��@CԓTuT�:�MM����L�GF����R�N;4Х("�qi�/�PM�ޕ�:�n�f�D�ZK:�NC���M�W���΀to�4��N�SRne\b8I�c�O�&��v��0�V�T�xΧ5v��N���h�ү��=1q��s9���'�j7
f,M��Ɍ�ͺ�x|�<��%�nUe�0��>�X�wR��a̺��R�Q�n�%��V����^�����i�`�xU�u��
�x:v�|��xk�Us�.?sσ�l�s���{͌�����Ǽ�����΅��<}g	H�\��<e��j�q� 7�8D�72�\�>zzvq�����}��k�-�*=�k  �~ ���F��]Bq�1���p��grDOX�=e��,�w��J�ܕ��@�c!�%��[a��;�*�g
��u[��,n�hК���d2����V��s6��liA�N.,�u�z��Y@8
l�Ss��U&r)������G�uDd��T��!jS�&e��F�́OWs(�/ ��A��0�O=���#�:[W��^���r+��}�V����3O���s�in�T����{\7{P[aS'{���3q� ��"��L[H���I��Y��;�#m�{PR�8��rp����Վ��i[�~�:����QFބ�'@��Q���Η�,��9,>2���7�h���ph.Ӻ��!��YJ�sݵǫ��Y�Ry�$o����
�m���!x��d�m�=����v�L�}�&3o��d�i��h]�G���m�\{'8�qr�U��ڇSY%\��-�Cj��S7�^��7� W;�p7��oZڈa�tm)4l�E�/;����,͗6�rk��9MҚ�YܱQd���39ŋ� �����;滥fн���6�\>x�J`"�����B�+�(]�͑���C4;���¸ZB�
��Ge_h�/������
��62L��.�N�u�Ώ.�>�6{����n��0��/%+8>�^���W���xFG�NӚk��:�~�(6yudbf%���H�B8mͰ�3�Ⱦ�sk�؂�)�T�܏ӗP�BYQ	q7�&=��Uw3e=2ޖzr�7OصP�|d�׃��v���l���_�������r`;=Y7��~�=����܊8��pg6��cyٚ�tdO �t��u0��]��^Ǻ���}�h5����S�_P�o�OƖ���O��F��;9�>[��3@��wfWxJ�F�9W�)�ZB¢������*��^]@QtWx�s������LS�4P�)���tn�J�#OBA#�4��c�%q7�/Et7����]���jJG�������+��WENK����M}�}��z�>�a�Zѣ�Vv�fG8�j�����ٽ,D�M��g[j���l`b��L�
�)�48lk���n����B�귲��5Y�s�%�9���:/���w{	:\�����GU��$�<ˣ���6��a�؞�CZ�����\����:��j�_b���l'^�2�e��<���nw��%vf��Ӄ��3h@����w���R{�N���^�HK�v`E���l��,�Z��{A̫�#V˸�����+y�����ֈi�(�W-�L��"���6{j�;D	���p0�0|�tu:�x��{iϭ��R�J��!�����J�ްm��o��ϕ 0��C,qC	��`��b�㖮��m�j.Jj'6��-"���=�c&��rS�M.t�`��0��aֵ���4����3�D�*m5շ6-��)�;w+�׌A)H�m�|����-�<���J��؛K�+Y} ��L.���̬��mw�C��ug&^�L⏆M�G&H(m�����e�'�l�%F,u���Udܳ0�[0HMh�G1�M��9'w��e�A9Ε���<��/���)\��ksY� *}\�`sY�F$5�P{n��,�E7�9��m�^_���(J����RkîZ��"������R,wu�SiIQT���AZr�Yz�R)K�P�%�!gT���"�wMK�VI'�zZ�DŢ�j�ITFHHJD�t$+��I�̊�:�Ե�[��9�{�繆j*�f�E��43D��략AwC¨�Y%b�Z����9�dD%£�����Q]Q(�]ݹ%Qf*r$葉AV�ej�)BV�a�P�NDIRU��:���2�$���u=,����s9�hz�TRYe�ffZ��T�(�DUU�3�"51C"�a�f����M+�*j0��F�Vb Ee$�C��W7]�D�e;�rD�����R*��բf��D�9�E#CYhk%qsňvQjTT���t0WGu�D�J�Tʴ�T�HВ"K�ij]4�@�>��������ml�]4���j��wa��+&�|�]ѝ�J�-oM؅uۈ��{2�Z�͓آ�3צ����eA_P!�xR�~�8U1_P?�}�ȡ'�97�*�t��?�$���d������P�?���On���ށ���0���ޏ}x]����"�?W�1��>���1�T9�ސuxOj��z�P�B��H� Gނ��#�x}�;�￼���n�oG�<���L.��ѿ<���9P&M����n�:1;����n<���S�xBw���h���%8#� �#���^�p��
�K�$t�x���B�E}Cƫ���)��Co����<��������S~Bt�{��}�$ސ�w��y|��N�?����7������s���|Nw���ǅp.'�{O&��~��~���|�x�ڽ���F��Dp��=�~���}#�G�߼ohzL*�����������#~C��.�������\N$�����o(H{u����I�|�&�;|O�|�UxQ��y�g���T-�󹻓���s�yv�?��ǫon�p>C�㿟)�!y����}M���y��<�}q�}����ǧ��_�;�QC�xC��=~�}�];�i���HRv����/���
�n��	����ǼdVy`��O@�T��p~(�����>�����v�=������󿝤���x��9P󿿻|B;z=��࿣��_>����zL.����y�}y�o��r��D}:c����a�܋Uo�o#>���1?�8���zO	��!��7;�s�Oh{��
�ㅟ��ra�ǘ�'�nC�A�';]o�<��;zM�	ӵ����ϗ��z��<m�<c�#�9���e�+�p�Ĥ{�b,��|8]�|�Ǉyv�|O�߾v=���?{�����	���P�!��?���Ǆ��;�?;�
�����nB����M� }I�������b�G�f\���Kʆ����7!!�>y���W�M>�����|v��=Ͼ7�o(���c��]��q������v�����roN�|B��,�7��������aw�z����,1#��b1쎥7
���^���>�(}OHs���t�|�HN������>�w��]���ޓ
��k�z�����=�����һ���?���=;xy�ݯ[��v��I�M�(_���*���S�6φl]�vgYW�\ڷ;��6�s��Kޤ�Ʉ���׎cT�Ex���!կM���_Wv3г��ٛӂ��Il̼�SnJ��x�٧{J�F5z8�5-�m
�Q26�d� Mԏ����zY�z/�]�H��o�2֣/��m������}�;�bw��1�ŷ��xL/�1�����]������ɾ�pxw�k��9t��r~M���>���?8������<�?����N>!�;�� ��$C}"}��~ݝ�c7�b�Q[���8��{O���e2���wG;{}��|x�{~&�~pi<�}�����S|M��S
�'ϱ��B#D7�������^��yp������(I��!�����99����x@���ǂ�>?�7!'��ɼ?\��xC�a�����<��� xK�ݷ�N��;���o�<����">��W_W+s<;=�7�VD!�	M�?�p��N���>~�����0���A�<8��������������t�z��M�I;������}���/���|v��￼�����z��Q�p�&"�m@W�i�o���h��1�����S���ǿ�����ۓ�~�c�i	�O�c�_c�;��<[s�< |IӵF����p~d;���<�۵є'}On9?&�������3s^6��S"��
��\��#��"��'��~��P�������9��w��?��/������������G�����Н'�<y�I�'����ﱉ���97����Ύp�v�^�����]�S���kѢ$}>�>��Q����9�������ÿ!�܇�{������>��;��_w���~BK�y��N'�ǄI8����o)��v�܅�������	�j��� L��=���f���R�=�C�a�zC�[�yw���o�������/����|���]��og�����ߓz���ǗxNL/���>����s�C�~������������S@���E�Ò�����ʂ�-��H��#�@�O�,zw�{�m߬z��	����w�ސ������o*��iޏ>�����󼧮��I��>ݼ�=x=&�P�G߿�m�=y�N�o����m���ц=g_�z����7�}C�1������xL.�~�y�ü;]����9�'����]�>8�^8���90�'���8�8�<��I��{q�߾= }I�ݯY���;xM�	�ޘ��~,vT�:���V��"!��!R�ZlW{`Su�p�W��J�.�,]����ᮁ*ŪOW���N%�X���"�$����`��k�k@gK+p
=��i�k������"јv5D܅�]����9Y7�&��N��welҌ���9��Km{�>�>�n�,D���0�~�w�i>���|>���.��!��zOI�Ǉ��=�ɿ''!���w����|w'��h{O)��_�w�~w�9��r��BM��������Y757B�s���z>��1"<�S}�Rq�x����nܛ����P��_���7�<&�'��?�ӿ;I�~�I�v�N����!u��k�1��c�"���G�|a�q�����=��������"G��2>��xD����rz;��]�P�����=&����!�H�� ����}�������I�S�~�cǨ���������� ���s"�H��>���,�TP�U�9�X���#�X�<LP� }���|^��S���>;um����{�������{�>2�U����7��s�;]z�<��~q��������>�#!�~�"��@�Y�C�n�qU��q]���>���>�"$|�1e��S�:Ǆ�;ӏ%��ݹ7�'ט����8s���;}{�o����]���������p�v�'�}����1���1���<"DBvw��^�͉z+ڏ�F{�F>�>��z*���NL)�>��w�xw�9ǣՎWoo��)��o�w����v��'z<Ǉ��ۜz<�P���������E���A�sg���F�>���-���2u(5?��8{:q�}B�U���׿}���4����}�yW��{�(x����X�|8�}Nv����99�?]�	�]�S����~ػ1#�0�}""+�b��!�W��O�/��^��^1;WTv��=p��@ G�;��y��M��G�nW8��< I'�o�_c۷�܄�;����Ҹ߽�v���:v�oo����;�A⏯�)�S{���׿m*��:�&o�{�}��LD��}��^\|N��\ro?�x7���]�=x���$���9����~8�C�x1�L����ݷ�Iޝ��<��&�~Ǉxv���|���;{{�=������>���]H�����[��|G�" ������t��\��}Nq�į�|�$�S�r�~q�|�N���xސ������u������r���?��y>���yL=�=y�Ǥ��v�fx8w"�/��-ہJ`���S��먄L���*���֌�u��z_9K�넸��T+i�� �\j��ޚ��q�<�Q�>���T�tn���ZH�Gb�q>�f�H�,��zGK��[��h�IX�m>�;h��G�K)̩
���[�Vb�X��#��1� ��{q�ϗnw���P��&��	4����c�_]�'�yv��S�oΝ����o	�!}������SzwϾ��o�_#_o��>\s��8���]���$}�o�����IL�B��G� |�����zO�zL>-��;ÿ>s�'�xO���~��G���!Ʌ�wݯѼ!���w����������"<>�9���	U?d��P/�]���{��T�� t�5`����_T�;V. �{��ǉu�һ�����޲ߛ*4ɬZ��u�p�UѸ����Cr���)��ş���z��~Zh��R�p�ř���:.EE,����q����u���8����F�'T&�V�c�N�P��b���b���M=ǒ��ԻӸϗ��߫
@!�xk[7��^B����g5�1=����Nc���:B)3S^^x�{�t�~�Z%a�1�g�Q9yԀ���a̺��R�Q폛�	t�:���@Th�S�^��l���'����Fa�3깬7�)��ϯ��E�����8�aA��{�vy����6�W��۔r������vaQaB� :]ilxUԠ�q��_g=� �osDh�V��/a�1
��\�U��}��v�������Hס0j8�����M͈js"�lw�;�d@|��þyn�d�� ,=Z2�h��'n���ԍ�\��مHkV�on.j��H�m�+0v�]�5�і���v�� R/_t���1�y/� ��pAø2%5�=����^Z�5m�3�ho�}�}��4).m$"�>����<�*��+X�1n�1���,��U�]�<w�sMdR��ͽ>�n��Je.A� �9U�1��e��?1�o�d�/��Q�F��[]�� s�'w��`
����/�I3)O�$tXq��Gy����d��$�EV����Ս޵���*K4���F@p! (�{*8��'\4d����Pگ�z�1���Jz�Z�_ϕ��t���\hqU�ф��q��kG�:a,UX���Mq�pTT������κDņ,"ju�9�q[1<`��u�v�3t�C��$�y״y�bk�}cwL�j�R\&�x�0�`	ݰo�8�~�C�Q��%��ZjD��]c�{b�Nq�7��|o����U"�Y<ɢې5Ù����#��-�6j֮�Rw��k��uX��B�I�?C�Ӫ���t����
�{O�!? �����/��ڂ#d�S��=\l�6}�B�IX<�װ�o�N��"�ʟdg˝~|l�B��w[s^j,��=�N�#f�Cۓ�u�\�][|��Z��[�{nn��siJ��h��t>�yW�a��l�,�������r ]w��0ظX��Yr�Ƕf��ԕz�͜r�s09�u�`t�E[����u����_\j��CY]
��ދ�T����F~�0N�C��:���uKd�c��E��2z?1�;���S�W�%W�W��#7'1�]��_ !2w맊��E���MN.mh �yY�T0.����Έ膲�\=U�b���ی������)��r�
͵�*k��Yׅш�j2g�u��ܩ2�^_�+�����B�ꬓ�/���NPAC�w�gk,4�p��L��*g���NB0����0xm9l��n�ۂ��8��c o����i�B���D�_�
��(�H�r�|���;�����t�a`#���pO�,0>���O�K�ї��k��Pb~GI=FP �*�@���]؄�����m*���C���UVa���Q�Χn���>,}[��;�uOu��6�����A��>rzR]�|S�w�&�S�Zـ-ÚMB�*j8���)V���3Ju�)��A����l٬p'�Ʊ�9:H�lCd;�����U���2J�G��k ���9�[�G�j�������j>�z�����f\N��9N,�J��B�02S��R��{Z�uм�b�R)�%�c��2���&��gڹ�\�A1���`�83�;ew!|�nl]N�t�F+��ۀu,wY��307qodNm���}���7۱?:U�Fi�~�������ܺ���81eͲ^#Xsl�A��(R��H�*.)v�S�?�f/�M��1"�0��i��u!�9�Rb��f��71ˡS֪���;�|������B�r��������j�l��	З׊�[���w�W�-��[�j�q������؈	/V������-�]j�2��Mt��yf����|0S�t�^��N�
T���z-����f���'1A���7�i꣺뮞?q�:WJ^@��u&����Q�üs+i�/I�,C
5�A�Yl7s^GN�*	VS�S�kF��>Ż\�VU3ty����������U5́�Y�y<���ޖ"����&S*��25w4q6�P�?uL�8.)H}:Jv����I�úl��\)/
��ԽWt�Vx�{9�61^���. E��2���Δ$� ��Cե_�-P��#bk�!���qϣ{Z���{�|�=2�>��(Ϗ��*>M)���͊�U��y�ҽ�TV�����S�A�8u{��s�����x�N֜6��7����Ut3�[��jsO�0v�+��d��5� ��Wt4��4�0� N)έG�[j]��f2P�3eg5z(���j�α[�Z�ލ��=8j��N3D��GN����G�,�v'wj�����c1�9;��W\|2J5�%Q����Q�����1+�CɒЮ|��Nf������5.��s��m����F�w;�h�_) oMD��Qӏ��_;k����ER����J��0�i�N@��n�˧V�ڙE��W���cm�G�z���`½I����'#~�]\;"S��a7�"���8�m���@<�����.��rF�y�*:Zg�b��ʼ2�^g��'G��{�<c�1׭jl=����wA�0	�C>�&�h�@|F2E�aK4�E���ȸ{:4<#�i��y!�8�ױeԞZ�j���D�e��PX�UQG7�P�6}����J�jn*8)��9�9���rTT��[-55F-�88nX^46ˋ?	�d���0�S��y���[�9�����8�ʏG��'�+4�Z��W=�7�v�]��A�N�SRneY�#�b�5[������OՍt~����\?A�^�V�Ci"�ɟ:�א���V?�}eq���i�]M�4���]��	Cq��B��*f;��WS{V*,�8,�����X8��}G\y+-�e2e�����SR!0��P"��
od�h+����[��+��~W���<�X�Ո�K�f���7jS�<��%�u���A�5�+�vX�%���	�8)����e�5��UU������MWt!8xi1�!�'���?T��r�[�d0�]D"�8�'�^�-T�W'������;�b��L�F �eW+��n�¸��k�_\뀍lƩ�<��|���NE>�'�{���t��A=;mqb����Px8�ң�{�d"�S����r�W��������X�R�e������R6��t�A��?[�~�t3�����Ǟ�qӎe�qtō»�N��1�
��Z6LL#���:����5�-�
�.1ru�d|�G w]���rb���'�s��^+c��Aݻ�9`obj1e��X�p
J~���b�R���.9봎󑧈"j���n��v땋�Bp�1
�T�]J ltUz�p 	�](E³���������f!�dv֝B���;ٯ�v�]�Bo=룦�6~UPЅV�Bk���<��֎�\Rt���b���2gWjg:A�.�0��~b�'~mցm粝�"��itq�S�̭B9y��j�,J�"�]�Z�ۢ������S{�lM�P�co�v�c�D�S�]��[�q��b��x�G��vÅHT���D���pek�]�
q�;S��*��]��V�|��O]t��]r};y,mˡx���Uݼu*��0M����$�U�����v��b_������ߪe���7ﳫ���f�rju�����4XC ���`�)�3�@#D1�
<��)m�g�</w}퀿�j��Rf�^�q����T��S̚6۠9Ø̓�(�\p�ա�ˌ6_yɊ�q�]�}rݚ#�}G�zӪ���\uӻ��?l���r��;kqң�u���R2B|�ᐄ��ؘ��<8*(�1Y���l����*}�r��7f�{��%bhq�9Cw�ŷ�s�#�'k���]mW���K���/��ޡŠ.*��*����n9S�1�����_*��f��f0k���E����gV]((ŝ�/���K��$ �mu�0�G�ܕ������g	�(��+|0��� �q��z3ڧ�2���EF騹�`p#��e�;��A���8<�:6�c�8�����שG0���2ø������c��*�(�e��N[+>w_fe�t�'�\�^�r�r��9��qcE+	��|+�JW��|�-LP�叻�p�}Q��K���=�:�in&����*�p�n,���࢖�w��co�n�߫�d��Y�Tv��f�V7�[w\)ҽ'%�[���VaGja����M7۸���3r��\u��J�f���-Pgvl�'7K�mM��q���#�0�B�E�	/���2��p�b�Z�R��[�\�,���O��s��K��n��+sT��^��{lt���r��v�%��.G�m0���lfpr�P����{��d�(��$�5��2�l��SL!�{
�r�`(b�R1!O5SWŹfo]X�{J�d���>\�3.�`ę�y6Ka�U��w{xuc��6�>��Ym*�+ۖKhIN��
4�n5�en��93:�w{!��nGA��C&s�SSw�p�=�L}�K�f;�;V�6��]-��5� ���f^��v�o����'vcY�(�<$�{"2i�2�7a��yG��>]��⭊S2�T䑊��}h�sfΗ+���*��2q@���� 74e�2���u�=En��⧴��Z�������{ɼ;/�}�s|���	�����>t���uf�H�m9ksrv��f��ݲ�-�C�������X��T*�ܻM�E���)\�%r�*��ޜo��;�	 �K�[�
A]m�Zd?A��	$D�������d�\��I=�7���b���a�ͤ�;ˉa�R]��ˈ�1��Κ[�8���:-��y��4��0ݓ;��#�j�v
��:�|E.���K�RC������캊�8Ij�w����� �`]]��m��HW9�[f�9s-��X+O^�.�,F�l[Ý�?��0�˭�W�oWsVLܾ��&`م��TXZ���B��:�X���L�@f�n�iw�[Ђ��9,�A�=�f���-�Ӊj7R��l���*�f^��G�//G:A�7wzd GcG&�9�2#T^=�w/eٽ��,Z�V��������H^~N����)N�LHt@7�f�X���yS��S����}w"3�>٤'�޽�麙�.�S��#��F�CWs���%�*M�Bnj�8�Q���N��������%�@4㵀X�$��{lm�ܡ�����R���g��%�7/qd���	�  5��m�c5�.�������X���N����>s��V�E��%�I6P�X�3(%7On��3�C��fܕtEҊ�bbe�f��P��o^�hl,<��g/�dV��Dh��!|e�K���tMm�s�e���Ⱥ����t#8�#/h�w���&��n�Z����%1ar�۫s�	�>~�yya&f��5a�М�[V)���*�,(�uE`�t���B1�P�ִu�^�hjd����[Q��::��3�wi�6e�Th�L"嬜�f�4�s�*�5��ȁ�\X/�ӹ1��:π�IH&kB�(���
-L��RDf�K�%���L�6��i��"ʴ�d)Ed�FOi�'J�#�U��*C�fŅ%�P��Гf��㓖)�� ��ȳ$9aе$h��2��,)J�h�%���B��K"UN��e�"��JTHe�#H���-V�-gL�M"�	()Z�S
�1L�@Ý3
���U$:���F�	*�U���s�"�1A˴�J���D-!E��fL�,AKCH�gZ�44SL����H�(�K*Tua�T�EV�S�9Ap�,-E�r�Jjb�(d��f�CT��l̺YHD���ib%�U*Y�c���Ju��ȵR�L���2�r$1+0�),KP�-J�%�<U0B��2��F�%(�]fR#�M�DU�!�!�<���Ei��\0�\����a����b�$��b�S9Eb'M�P��r��F�Ϗ�w��V�Nʜ���+��Z��
Z�ouД�K�Y���ݑ[�d��Nve�u-���û�"��!���
<�>��W���}N���ոՀ,��:�v9�GI�* �CN��p:�e93��]y��c;��ۉr��(?�g���!�sN�Ë$`�3d�t	�=�<���t+��C^4��(�)���Q)q7-�p�.����3J�0S�MB�*k� A�����kL�ʁ���-w<�ݰ\�{3�?>5�.���N�8\���w6�n�o�Ub&�L��S�,�p��o�`Mk�%N��
��]��%�@�L�i�c+�[	�p�.�D��k �6aP��L�I��|�R�;&����K����^:�iU^��{<����Rb�村��2Y��]�e-�1]��ө�YԵ�ˠ~�@��t�]K>�?���g��c(�']�y�y\��A�������8�f��`��2=��/�t�����ڦxW�Z��v�TU[��&_n�{0 �mdƵ,GB�A�HS���
�"42{A���K*�ܽas��$o�I�ӗ見�[yn_�v��ρO2�1�c����燽�^��f����&$ڞ��[����qG��e7��&uG���mAJ�JX��W�N�u�K��;ú�	-Y}�!�W�!��o;/������71W,,jt��2Y��&�qV��,N��YO�QV�t�㝁�9��8�#�)me��IN���&�,��������nt��*�G�̴x� ���~{^�U5́�%�G��N��}W���S��E��ګեy��8*_��p�+6���ชRM�̠+Do9L�T;���.�ܑ&.n�z���K��5z"�Z�?1[�TT�Zi�K�.C���4g�U��-��\-��r�ǬF��3�����Hd4�cA�L�����Q[\.�_��,B��L�(��1�o(��w"U��+���a��P�:��*�GE��#ę�~���q��
�+O?ğg��kO�gG"�N%Os��m���Tm����U
@�6�&cz�GVG�/��Y�����A����f�3Ԛ���e���8��Vݑ��:�U�or'ff����H�C�!H�'_
�4}���g:��)�f� �u��ƥ��(�{�<�'h���*<�p��#ǀ2� ����^�æ:�i����l!q�v5���4����C�Z޹�<\ɨj����VB+Ⱥ��t�#l��N�_g�3Z�oWr�݇��l�~#s�Q�!�#��7��ڸ�̛MP��V任�V�K0D��1A�Y��BF�Y@<Z̬�˲p,�FS�݌�&��vwY(G�-���76T=�.��ݾ�A�i��?�j�o�.��z��*�y6���$�^n�;:&;��W��W�TȂ$M���Ѻ���G�䩒��偮'����T�P��;��{Uϋ�����U����i�>�1��V���jj�A�����eş����6>|����ȡ��7���+la�<�h���KλSy���^T���FҬ;��^��p]�@�^/{�u.��<k����ˮ:G��w��5�SLsq:��T���UdR���Y�V�5\3M0��<Mc��\"��,���d�gR�q��2UDNk8R��T��æ�"�,���Y�����LT# U|���������[��0��Ĳ�s���O,Z.=��.��	�ۦ�<��ܣ�g	T�&	�:jm�n��0꠫�����X�F������Kw,G:"�s���]H۹@0��[6�J��r��==���O� �h�P�:���]1»N��S���Z6O�!�ˎ�#�IV��IL��@�R�>��R����9<��;?p��NۨN>ux�;�4/9mg�8�ʵZ[{����̡hU��Tq����;��\���5�����CN�ZWV���(x*25�����F�[R���
ڑn5��$������r�(<;*���`A-��Z��]ąx����������-���F�*����ꪽ�P���w�����:i8L��<�ҟ�������E"���0��E��~��r7u���`�E8ss�uB��T�k�����
� ں|"�O;�
Tۮ������܈��C9N�6�A��U�@��X@x	�#Z=r��9��pt���)\KS�1���#6� Σ5��.cȫ��� �#	$uE�[����:<Gם7���Q����q��SO&�x�C,!�Jwl�N9��,W�`�.�hu'z�)���Q�z>�싡��������<K6۠9�Q���d�Q�)�A�KWTU��a�X8X_#�~jy�;�����q�O������~��c��bJv��έ�z��0
q�WC[�fF�:`T��xpTQ�b�'����M�$EOa�i\�v&���Cm�l����E���nt�qd�@?t�"�����e� oT����	�7��T�Ts)ܲ�����sCCܟ����S����c����|ga8;�Q@��A�x��3��F�#��o�� QZ�����x�Ϻ��c���Ĵ� ��ONI9���;`Vڜy�;��e����qHNӧ�C�+K��-	�P��Xv0'/���}z�r)�*�d#��)�I�N"냺��gc��}��D}-�l[���`"�+�G &/�����r�&���{�A+ڰ����e�8Q��hbnЬ�̺����
���*���<�;��W���;�7���m*�v^�Od����բ�i|O�PKG���q��	uXy�6�+���W�8b��7rf�Q��ac��R]��O��3P��(�V�jÁ�\-(�H�r�ʘVw��Q�,x�j������u�v�]Q[c�ǀgi5p�!'��T�8I�TTP>��R��P�7f��Kȇ�6�V�?wu72͌8,?�KF1��s��p��۸qd�Fj*�d`'Q,W[��@W����ٺm�����廎]��	�o�0W�hpO�H� (�}�����ó.zv�HpuU�`�+0Oˍb�������$C��v!7q�f�NI�O��fLk���JwI���⛈& !1'���6S7����]l\'1�����*��f����"n񹔡r�u�³gL���^J�i^��{<��ה���E+�W�z���ht��)�p�y��Ay���}�a�n`9�4H]BrV4�Z�@0@R�SD�=aA]�(�q�3&m�:�Z�N��b���YA����61/���&�}(aqTw�:^#}.���a�ɌBy����aG����#�C���b{�2���LFu�Uu�A�2Z�e�ڨ3N�k��{�8#�!�k�]ɘ"��W��P.Wt`)�nX���|.�,��1������]���dy8,a�{���w8�,ed�o*b����AN�f$lCWDEF�O@���h�}}c�&�t�W��HyS�mN��x{��c�� ����b�T�_�</�ڂ2+ײ�z9��S����p��wt����V	o�t�q!������+�s��/G���oe�uA׮�����Kz��ґ�M�������~��>B[�����<b���t�`�`��8 n`�����d�O�L��z!�t�B34����0||+>\�xS��Ty�]#(��@7�RR7~�}��\'-��N�>ɑ�b�Lh6h
�~� ��^�-���:0@U��mrD`�wUw�v��aQ�Wc�?���ko�\#���V>�l�t�H��@�=$����2���K�#�P�c��9�f7���ٌP�_�)��sg�Av^v��	'اcg&�J�sy�C/��˅Ri�p3�c'@X���'�3�]�<r�b&��B�WFCQ+��ٸ��1`q`�Ӥ;}����Y�F�	+j"ū�<-��:�N��t�|lY���<��jf�Cpltz�5,�a�k������r
X�����O0A�ph��Վg)5q72�f�<��Qm������U�-���-�=غ>�h:���*�@�x}�iX�p��ޕ��
��Z��wO�B����W~(_$x�����t�jb�|��.�\:�C�*���t{(�����\�h�Ǜ��H���EC�wp��<I	A`P��+B�=��X���3(,z�Qǆ>�.�?Rn����^
���鏔�'���{*'r�Esڂ��_���-��!���B��S�z�Voe��6������r���আ��ş���xJd���!;��F�v4#��/���x�߰y	�~�i^|�۩'�u� ��a@��:��
�֪+Tn�]Sz��S6��@Y��2~e�ʕ�!�$_���~ڧy�ߢ�c��>�kަ"�T��,O��k���ƺ�C�TB�z~�e�Fx|�sW]����^��}�Zxd�q2������~9mϟ�����+�q	]�@�Q朝�ǈ����G�:e��9"G\�)N�k$Ӛ��m1%r*NmIH�����랳�a���Z�{@�o���q؍Z���P]b�%J���h��gr6�&�Mb-�j���ʖ�hݫP��m��)�F.�t�_��՗�>k2oee\�|N�˻XbXr���꯾XԲ;d��� 36��I<�d:�G�:���Y\.-g�� �>V��ڼ�/�oL�S1ڹ�;3u������ 3�Z\ S��
�Sܽ�{�u���ѹS��u��Βt�y�Dq��J/c��/�.��1�Ѕ��UL,��@�,��0�K�Yw��)��ž�.��Aq�g�'�^�*�H��	��w��]�9�2���~cn������[=�==��^��Cs6��ljIL��<Dҟ����)O�b
E�	+��@�x�4&=D�\�=�a}��|����M�1��RYP ��(�O=��[2ꎺp�~�`�6
NzRY�o���a[���q7��7*��P�f8��=���g0�'�Z�t��LN?��.�w`�� ���c 1�	���Z�ǑWBc� �ΝΗ$�o#��~sg� �+g�����x<�]m�rju��f�0E�C ���!E����E�*,AT������~���2�/���mzf�]�N�?z:A�I�F�t2c]K��YN�}׮6rn���&����>Y��ڕv�u���,Pܘ�c�4R�:ܑ���1����$k�o�g�cA�n�Iv��g��i2#�����j�"�rb`<@}p�\ �w���E�Ι�ɴ9I�qw�U�.TО�9c�+�������\;��5B����,�vh��>t{�Z�}f��w�B�?r�*v�/���s�T�4����p��-�7�{�u�]�AVf�����b�e���ɖw���lK����C����#!s�$U���'z,5�S�c�'X��`��kХ4�n��*�z�vAJ�}�p)��|�9gA�t��o��׳��zFnJ�N���8L�i��Njc��^�G���w�D(ؒb������)�;g����W��[&�On�B���H���ta��B��!�y�cj'�pj#�(:hp���.��5��7~�"���m���ĸ(A�U�P�'�i,]@�Ф��J@���aT����ea9}cOkgFb�z��)�[����Q�$�+��\/䣂���*�S����茼��D�ƹ����ݎ�3MT=�q��1\q�L���C��U����en�ܼ�]���Ndu��$\�c8-Q�B:�p6S�P����F�0�_M��A&�g<�Z�@U�KϊY<���#��}�J[��*��b}��ἱ�$F9'P�VMC#�0u�D�J�dWQ��;K�OS��ܔq���ۭ��{���3M,j
��O�ɏ��Ր�b�%�Ay�+Բ�{���zeA�4Q���G�}�=��ַ^W29�9<�ȷw��S뉸��8YwO��t��`fB��S�*�b&C�w%��]:� ���ڸ�g�A}м�/���I��$r��StF1Y[�95a��'t�|)z$N��>��&���\IZX���Q����]m.c�1�Xތ�;���s���TJ�6�X��3Lt�.����1#�3�g�5*����6���E�z��|�P�0�u�(�b��s�����vPK�`��5���^�ݝ9*�
�XR�%rs��\ ��/�-5wB�`)����?`����x��*��~�����hZ��h��Ʀ��ȱ����ed����=j��u]�J׺�7K����\ƾ��Y���m1�ʹҋ��t�}!�ov��ρMG7@C�`�����{\M{y��ó��^���A��<@v�B|�D�:C|]����ץsNx�G�8���T'1���3���1�������e�t"��z��Q-	mq�i�:�*r��Wލ����X�ăq����k�w�N)�k�,G����:!k�-�'uZ�_-��0΁�{Z-TMm���0Y���qV��5I^��;2���Bu;�Br�2���b\��w��ȳ7:�%aՖWm��h��I��)ym���.�4#{S��x�@�h�a���	��v5L'����,���DZ�zq.�]GdmEE �6x�������`y)fkt�ܕy%Ḉӭ�mb�L:��i�� 8ck���͐���W�k��rlN����ޥDse�R�X��<r��\����R�C�tW��,PҮ-��]-��c�����Vj�����Q��-�d�yqv�V��厼�&��ͬ��F�F1�MY�4'�d�4�*'j�<h
h�L&�H̗���V�8fGf�*n
�W�٫q�e�}���4��G��� �� ��e#�OM�m(WK�p���y�z�!�ԠY��7wGx $�V�ї���4#7���K�c�n���.�F� ��W<'u��>���1��r�(�0�"�-S�qӟ.t�:jj�r�e�r�e�[M�`�Ш��D��SG8��@'���t6�uվ�nVd�R{s�j�����V��]�^rkX��ϰ��W�W�Q���b��5�H��s��Ne�|�� �O
S�R���R2Ⱦ��p�-L���z��:��[������u�"꨻V����oV��b#��yPo�w�:eve�/Asv������^d�D�m����ܣ9��wE�'҄��w��3w[��omb��6Z�1�hd�#Jl;}���=8rj ���xk��U��6��S�����H�+E]�ZUᵱp�=�nZ����k3�q���٘k�*��5z*���ڠHh+n�=�����Lwmf�b�O��x�|)#��� ��=���I��U�'Dw�R3d�1���^�*�tJ�o:M}yjv[΃���S���	�b�Cy[�\�Ҵ��[�:(z�uSOC�6[J�h�Ė�܂ܧ|�CP�Wt�� G�A2�=�2s�ၪ/�z�F/��^��������՝ƥ��1Y��p&�Wj������KK���mh�\ky,N"��ޗ�6Sx�*<y�/�2ub�t���=L�Ϗ7�jT�� ����ñ�<����Z�� .Vh�ʋ�|��a�O�k�xB9	%Fa��{'*���:��<Q�5�ؚKnH�=�Qɔ�X�ܬ�򍬂�lT�ԛN��ӱ���M8%��/H��]I�����xN���G9�e�V��Έ�C)��c�Q��+bSlmѼ��S�!�e�Փ���n���C�fVA�^m(]n6TVtY�����+e.0���{�`��M�)
��󴾋�"�7�84t�友.�b�.Ǡ�`��j�
7o��um*����t�h�w�;[#�Q�C^��:��NT�Wك��O� ���"���-�wH�ėQ�@���'\rQ%2�@�
2�\�J!7]ĭ
�pr�.Qr�0@�t"u#���L����-	S�Em�/#X\��$�B��*����YĠ�R%e&d���J����[9UiHa�B(r�EK2$5T�:D]R��%"��&�T
�@�L���4�\��UvDA�I4��E�Re�2��jF*X�3��k(��	��L�Bк�j��\�
�"�����+���kLΡ)�qԹI,2e�ei�dkB�1��J��#2�'S�e�P��FVQ�ģJ�	�W �PQI��25-iPAYP��V*��9e�4��jE��J(����T�.!&I�D*J*�Ah�%B�SC�
Nb��������7z���/�7����:�dOz���1m��^�q���}����]��(7��W)�]<gs|�Zɶ��ﾪ����X��=�ڻ8����\cv������U���\-�+O�~LS�rgu�5F�g���>H�"�ƞ��Z�1^g��?8=1!��KKKf��x������ �)�	�}CK�[�N�� F?���S	�C1�T;����U�Z��'�	����ޭ~��urG"�P�h)?ZR��f1���{W^ϼ���9�/��R��"��Qh�y RC�	���	�mTJ�e����N2a�썸b��T��Pw7���I	�:�T
FGAc����w?���X��u���^��b������5��sJ9^�޵&���4E�0o~�v̋S%P@��@:y�кSdqA>P{��`.��(�����?'��gŵe�&-M��)ͻ��F\���!(<Ld�M;���֑��g4����Ѯ5+����?TBn����5�@��叱T�=q �|{UIpq>��y�^>&��VѸ�1�&�3���{lgͪ�63�Sr���)��\Y�@�2�oz�]D�(� «����d��U"��I���$+I�V�k���;*]Nf$�^D�fdd%�Dz��[��H䬭������f��4V�"A��s��<�],9x��u�ޖ��4���Krev�R�-\�r2,(�go"�[#��N�v�����UU_}T�\<l���1��������C�/�͘ѼhBI�ik� ��@�2v׭ː��eu^�[;�hz�#iz�p��	��מ��I�{�x�x��ʼ��~�=c����,�wS����eb�jY�/�S����2��<>Tx�#�ΤFA�M�m��M=��I�56fp|�:�V�	dG;�b��L�F.�@�_���*
�k ���G�t�$x�j�=0�����M<�gΫQ�N��-\���nQϢ���0卅n�;랎=�hV��ž@I�x[��
E=��U�~ּ�ѹ=/���(���5B��ڔe�x��AS���#������%@�,���l�åL%]^���C�c�̗�g���
�:�.|=u���	��w���9�2���Q��3�ڊfV��W�B�k���p�Ûn�PK@��]q�/�FD-Ȼ��nv���sg��R�}���>���cr�
W��A��L	����PX� r�.�l�w�X������k,F�x���ǆ���e9���r��v.�Or�5mU�;P���UҾ�M�����������cBT1Ҽ��i
��>�a�n��EW�/�3�� t��M<�FYz+(pݡ��>���:�K��$O�u-�Xv�q=�V��2�"
~��w�b�U
�OF4��sU�De�n9wb�ɥa޷�`�m�3NP
��[�UfQ�>�J���j�"-Ԅ�}х�8�s��3l;"Y�<
�0 Td��!��Xu�P`���}/�{Vg2�?<8���>�as�IK�ݽO���6�f����%�r�tU츷Y���by��.��g��aZ���wt9m�ƍ��ȟ���khf*���V<WCo4E��#����ũ\�q�Y����T[�v�ڦ�k�-�f-�o3�q�Nb�#��Yu��[��F�s�2�_7�g:��a�×�0\I u`�,��r;;_�_U[���.[땏��=[P�[\�u�Y�RcBe��%\8�M.��Sx3���
�ۅG`Q��61�}���:�����#{엯X�go�x'/:���	Q�r��^]�HD^̧��aGf�(M�*�+��� �b��t�K���9�Ԙ�j�<��[�*�������}"yvg%�{\�QͶ�A�v����+�1*�v���7a�/{N(��������^�GK>j0�{�]=Xz��pUq ꨉ/�"T.��/�
B�b�i�D���]g7y��5��{�~W1��L�v�{l9�CxO��DfL�ٷG�֠����v^(k/�p��M=�7����:`�!�1�R������a4���Q�#aPy2�����WMB��%
a}�����_U���j[Q#[wԺ�S�E���n|�f���:�|������}�3/�$�g�Ɇ`s�	�o×.�ҟu�z�@y�Q��U��l���f$0/|���t�u@�;�7��yq��\r���,������Ό�r ��֤O��K%�y^�;sQ�?G�6��9�&��N��aT"�!#O��>m��rz�^�o�֮%8���Gh���ngZrxV�!.l����K�[Z��mT�,p��m���r��,����_nli�+�淪iѩo8Jj[Q�63�-���ۃqɌ���/�б9��@i�ӣA�iE�3�?z'�ᅮsB��;ax�oR���bt_����Z��"����H��=��)\wbU�ͩm�S3�bC@ǛeЛ�M��	]2W"��W磌ﾯ�9=���=�%O��Tvnft�ȧ:�y�Z�j�#���B���Jjn���8:���5x5�(�ݛYQ/fs�+�%��7�1�� omv�&T8�J{����!v3���O�3D��}=�ڢr�4O8k{2Xۨ�x3Z�\��y��U�p�:��a�b�
��D��P�b0�i��ӷ]-�w ����l���>c7��Ɩ�=�<���m�	��G��)�զ�Q�F&�����/��z�)�.���_=��Nu.��Z�o7k(9b:22���Iw]1}NKu᪌S�|�5����I��W�(,�l�����$��J����Z�/��%F�{k���=Qg�������!�Q��Iѻ��y{+��*�0]=)�K|C}|���]�C�#�{$�x���z�D��[��Q���Uȯ-��8�O4Փ��[��ګ�3ƣ�pE��c[�9�#�[�� �1-(����C��<��Id<5��5�c�I:����^}����.��q�WweLi�}u��Z��&�ѕ�Ґn�8o�X@e��&:´��i��tJ�S�	9�'8j�/p��X}�D}�>��6�[w}��|�>OtTE�2�]3P�S�|�D����ڼyk�׫��Qx��W3���������
��E9�4�3����v�5,�kX��SW�8��"g�}�5#��%�k��p�p���xq�3a�0�OWE���X߯̄{�ڛٜ��6�k���n5�73�Otd���<��:;C�{���̯�c�ś�oVͩ=�j/W��z��^�h�h�f�oye�h��K�hQ�C�����"^eQ�}�w?e.ΔX�!�C��q�m����9gn1�'W7��eD���UoJ�mu�R�Y�
��m.
v��S/E�|�G:�����Ê��|U��,�Wv�B��%�X�qQ��b���i���WZk���gf��v�x��
6Z������	~^^t��a�J�b���|�5K���&f�Y��T�ʋ׳U�Z�ˤw��Z��J�&[}W7�>�Co'p�O7�i�13�Q��:a��o���� 2)�Ml%y�t�<]�j�/s�1d�o*s�/mS�̮Zf!��y��Ux���l�P�{��Yq�B�li�����U_TGѻqO(l��D���@)���:�>���Tr��-\F���զ��!WWa.�3��8wԧ�k�e���C�.t�*��=�2�JRw{V7!����3w��7�\�t=���Sm�@��h%A�CK�>�����5�Y���&�]��j6������,k�\fվM�v(9_oO�P�(S��2�K��jްw��Ż��s��E���nB{�����"|�ǹ�rL��8gA'l��\��Vһ�r����Q޷�`��y�ܲ�ʭ�o-��kX���Z���$Z��o�[�zS�\v�s��7��3l:��9$��µMA��t�.
5\:��tuYZ�_d�ݫk��]C}S��w9�&�uK���>OԞ��>w�~޼?\�__��v��zNvZh�x�j�
�f�����gu5ʦ�X�M|ہ�NTC�dLk� f*��n�I��Ŕ�DGyW��6�I�����v���O����D�� �X��Q<5/2D�\ˎ����H�2V2,�`' �mO_�~ʮVv�}诰婹m�uh�6��\��6��[ϓ{��ߺ�H"��Zv)��;a"��!O&� b㷸�b�^z�����f��������\v/�����V� [S�3Ӹr��g��,_���%��8����{�.uq+�o��t6��mCy�7WqaO^zό��'qxc5{5Qf*=��Z�����ڇ��<����g9#�����Iֻ���t�ޭ�u��C����yc��郪n����!WAH�~�1�,b5�����{���_�bG��@�4}˫��+ҏ��UV���O��JF�^�yp�}p��W���*���)��q'�����M5��~~��Gvk�]��Jyc���-���Ss���@���]d�=�p>�I-�Χ��U=#�{���ˈ�m���<��}�n$Mm۬�w;^%�"����$&��u�)�}���ϓ�ڶ�A��ϲj�=Z��Pؼ]ka,��)�����BZ+��]�]_b�����:Ԑ��x�,P�l�7]�$�kѳ�V�)��/CP�x�e��Zgm]\�Z݄9�B���(���q�S\�Z�kŦ�!ׅu�\�,f�EHS�����P�.���YƇc�erG^��p1>�� ��Y)����HsFQ����[Y�T��OkD��}���D�6_g�pT=��2�U9�B���E���Q+^X�q�u��.h"�%C�O�y���s�W�'Nrfb8��rV��]�>�Z�㸽�����ң~�����W4ø�8U	��u#�
ڀ�230�uj�G�W-��!���l*Ob����U5�mƻ
r�"~�:w^�vo|���up�o�o௫��ʏ��ۍյ��b��z�sQn���gX�]Ti�G��e�;.�kkW�>ФZꁘ�&�����[�ػ�{���땨����lS�ڵ���7�|�x��ػK鹊������?G���='��)������S-y��7���+˸-�}�&��8�1|z�����KԷ�{�at��W���B�JM��M�����Χ�]X�JN\���:5ut�^���BK�ٮTc�{�Ajo���綧:�u���m��!����C���*���y���}ym@rE�&B���e_i��6�H�5bv:��X�>|1v=��V	�-r^�|=o"��Yh�6N�h���t�Ftp�6�Y(��[����,0۩U٭j)ʻ���^J:����N_`���rUQ�菣�WJ+[c�O�us�z9b=���oCYq���I�|�[�HW&dR��m��v�A�|*��}%򸤨�bOn5�[q�l����o!�z�n�Z�^�i&(9_&hO���H�3Ώ��y�U�͋]ؙ�1�Qi��ޚ���ݩ��o>>]ή���z`�?�T@��p9p��L���O��^4�n���;չ	�T�<2��њ�OȺ+�;(�zs��&��s�j���҆�&�_Co"�ۚ���L\g���ٔ����#�K�ή��ɯ�vMf�Q���.sI��7��NXJE%Wb�L�7�����Ì�
�ܚ�%�����]��ig15�n5񩛨��Qn���1-��X��T
p�,���t�{_n��
�;�kz�\$����y�݌���Y�6^������ˎN�r�I��:b�����ȕ�3;ޯ�:��v�dT�W|9嵅��M7�V��bT�Z��w}b��k�/��Q��q�����qv�Q��ҋ'!t	�c��f]��:sn��ծ�a�Y��.A@��-8��nDZ������Xb�+u3���Szr�8)����SFѤ&��}9��GZ���.�Y�R�krH� %,�dP�u*�QC�����-:ق��	�>��XeΡ��ɑ��DTnS�j�Cn5�����J��#)-��s����aS�hx8�Z��\�{�M���_-�\��k*�U�a���$�Pys�����1�(��}�˃�����+v�'dT�L���e�ge]֝���C����]�:��Zg�{Fn�q����j�X�x�F�Ɓ��݀�Xs] ��ˋ&��y���%[v���u׷԰�R�Iu'*,U�й3	�E;b�i��b�tcb�6^����c�o���nS˷vV<}J��r���H����[��ɝ�
�ԏ&,�����L{V+��;�Q��#�؝s��~�XA\6���Yis��Z-���_	���*=�K�EZ[쀁b
�ޡ�Gl���q��6_1�fd��Ll�boìYyC�$R!OF�զ�n�G.�t������j�kUb�z�dZ��E�����:3��b�\y{+q�7r���.�v��l�i����9kI�&����8ꩲ�];��"��:[MV�4�
��*��kTrA|cw���kIX���[�F	��#G^��=��#�Lv}df�yˬ���ctÖ{7�:3j�ۭ�-�)�)�8���ƗK�F���ۈ����h:�:��}�e3*�&̘.Z]��U;-*����nDҷ��ujf]�R�WWu��4۴�6)9�����AF圊�<
���S�;Cml�_O�Gm��![�����V��W�]=U���)�ᚇ�/)�ox�=�=97X���!�r^��mB�7%�|�k�7���x���zvmia�`X�?^5�n��*R����R ):Dz���X6�QZ�yS��G��F��hM!K�W��٬���é��샀���ٸn�IY��MM���l�'�YPW+��ǟ;�ߒ����[
Gf,�A5�6�	ݷfG��s�f���x��b����f��(�e�QJ�p��B�n��J�32�n�٠�����bTL�S�ks�G�J���b�V;*�:�un,C]�����rv�"�^)�1�{x�Wmr�6���B�;c��1��cM�핕-W
�;��/i-fLU�w�.X��VP�^.�ͩS�����;{�G;���+޺��`˩J$
 ���cyΨ���գ{�iu����%tאAJ����C����CwV4���I6�>"��u�y�z��՚��56�s��r�f�S,�y�Hİ������d=q��uc(h��$�ѝ���*"ܺ�θ���'uˢ2���)�޼��v`��O���Y��$��%PL*�U�*Kjl"��
(�P�9QrB2Ĺ�C�"T
&UE��s��(ՕETU"�.QD�E�:�UQ\�RJ����Y���"�
52B�D0�ʈ��)��U�3*(���5 ��6�2�:s��e�F�%��9W*���J*�F�S:K3Z2�ʠ�%N�*�2hI��9$$d�h�P\#09p�D

���\����d{����y�r�'6G"�T�͑�,��+�zT�S�{T�hr����jQ�t@��r�'D�U�*����$码�(��g:�z-$�*,w3�Fz�N{�r!$ �=�2�U����((�R.�I��P+$I"�7w��g*��I9�AUʏ5us�
���'�D:�*�+=�����v��n��R��t*3g���ʢS\�B=�*�q��u���j	�G�
>()^�l-p�y��]��Ɂ���ٸ�Ry��ۘաK޽�*Η��Ö��q�l��u��z&*k0p�8DF�?�W�W�T⭉�\�Zo�]=��s���=x������i�����)U�z>-�(g>�ڸ-�-sD�ޮqλ�����0���T9�~�Wx��q��[��l��g��S��%k�����y�OF��9����|�{+��NN���o�e����*T>��(��v��}�S�� 9P��Ŭ
�H�LX��4=�aL��}R��F)j�Kb����Fɉ���㳷�F�j���V��]����7
�~p[}D����Lm�mש��P��r��N3c�^8[P�{p�۱AJ�:J��CK�b�b�;��	q9�k����vk����������������Z�/&>O��o�ҧ����y��nB{���P��ȅZv�u�B�I�|���b8�Z�-U�9v.7��8��0TCo#;�u�l螫��9a�q�N3p��.Y�jP
L�b�¦f��t�%o�[Y 3MjO��onEom�A)��r��;��2��q�m�}}�\�����]<Rb�۔�mN�[
f6��D*hn̻��1�&e�L���<�V��wi�}������|K�	��r��q0�>�>��V�^����s��m�et�u�U[w5@ݬJR�ʂp;"c�0����6��r_\�5~43����"���|�'(��sBi��\>�l�[Aܕٗ�M1X��p5�ѳM�h��Mk������n�S��Y�k�.�]1:�{1Om\��bA�T�)h[$�=�OooB�j�#��{T�aˍc/P��*�z(��;��V�J����9:�ܮw�z9�}�F8{�KD����2�K������u��\�X�&�1ۅD�|��Bg�a���q��xc�=�'K�	#���
m��V����+�W	O�Ru���s�G4�i~oɗ�֋�E��s����c����Q�T.��3g��a�&�t�k;�"j�n����Zm���U��+k@ق��#�d��S��cf�2��7��RY��w~�ojk1s�n�0�/t��2��k��5��҉��|����mn2�뺚.�U)��C+�N���7q�(��:n�#n��ϧ�v.��YVm)g���x-��9b�M�����	-o#Ƨ_!U�8D�u���菻�g�s����zg{n��io/�p�^8Z�y�)�W���u\���O9��/:-���éԖ�vC��f�O.>�mㅴ�TBt��zaX����V�MB�>N~.@N$4�zWtJ|h���bqx�D\L�����>��z��K2o���A>���wm�M+��b�z+��y�oZ�������:�5�1�P�9����o�^��5���#�6'�n5q���LTbv�x-����r�/����VE���\�X/%��ݩ��T�4ð�c�
�a8���Gh��*��t���vG�o37=�/|�n��'�}���6�j8SPۍv�>F�s#x�inm�Z��ܝ�龸�}G�Tzyo�D��T��^��d
�7�҉��3ٕ+St��C������a�A��{��"�|O���I�L�*�V����@�v�S�4!N��6�}�k.�,'jY�y2_T���7�4j�e�maH�#r�x�X<
8��y�`:�ֺ:��q�{"1����%B_fvE��f�tѴ���Cݛ�(��3qt��*�U8�����Ť��Z'�ةf���[=�-`Q��������P���j����W�����3*�~��nr�{�N�s��i,n�7n�y�=�5o��>�^-���}�Os�,�\�|���!�[q�	��J��]�
ޕmp�����|�sٛ�y�V���PU��W=[�������I�V�Աs]S��RSx����|��]gf��b�����=�9�.��Ƕ#M�j�co����6rn2u]�c6U��G%���Z���%"-����O;\5���
J{�բ�C]�=X"Ӈ���smؠ�}�0T�p��mu'r�5=��gt��S���-j�v�۹ϳ\f���ʗIX��;��ѣ�Y"���f��N.��ә�����w�s��E}m��t�dw˧���T��ۚ���mT��o��."�׽ʪv���J��v�n�a͹�E���Ag�:f����2t��������y���&���m���\u��|����-2w ���L���i��G}�Q�fv��m��WU��&밶�,+���_,��plG4Y�����4T�W|Z���]dF���)��6�;��]����WC5-�fM������V6��Q�o�A�9�5��ɯ�Sԍ�%�S|�7� +�l���t�o ݕ*�7�:���e��ޚq�3�s�I�|ک�Y�K�{o�gVl�oV��g�$�NTs�!.�ka�=w���^-�ޫCi�U�v΍���N�u����=���IC���m|���G�#X�k�f*���g^��ǣ����=��]'z���9����r�
ʭr�� N����f��{� op���qޅ�=N�s7�S�u�Q�N[�je������p�z���X37`�Qŉ"��7U�/1'hd���M�T�;��\+qj}��k9�M��L�6m�Ͷ��(��́�6��Bi�	�J���P������w4���lj�����k긧�/zR��I���:�΁����K�Q��B`�7Q��q\�^%���qV1y�y�ymC�#�2�]�T'�sHo	󌦫����ߊ��kؽ~@��\OfQƪ��-�Q��4j�(zܤ��m����Q~��"IZ�s,P��@Zf�m
�|(+�\�룻��o]ذ΍lB���L%i}���1A�3I{f������JC6���$�*��[%���%�	m�c<M�Q^��菢>��PJ�֠ݟGwvިk.1�ڄ���M�B�:~*�=��B��Y)��y���u�:�Z�PRy|����o�T7Mؠ���/��wv�ɷ��X�ؘcTLڎ]i�	n����{����Ho�\m�|�Q����>���E@Z��.�\r�4�ֶ�<��q��&&�Jg�B�R�Y�=�j�~gL]�HOg�YN?}H�7���8J�����L�i�:�,�N�����@����=�Mzbu7�ʒ���72i�n�����I���k�!��6F-�W�]�V��|��#"u��o��n�}�V�'SK)���k�+��ȟ�z٫؎�4��I�6f��H��3��+;ou�F�b��/��sV�O%��w��Ed�M�>͹�;�޵�9�ܰ�ꈗ�+���7+���^�o_/��e�tǩ�ei�� ���K}� q����aWySﮢ��ξ=l4:҃h�]�%#]Z�\�:���6UL�Z�i=ʣ�lgiC���XV2�gEŲj����s���/;��41d�W��Nt�\�F_a]*3Dv���G�ﾀr�FN��l�^��0��\�x�&�*'��
+���N��r���Px���)i�����˳��2��lf��ǫھ��m��^�I<�'V;9�Dl=�|�C�����x�u�QV;�M�SH�5ʇ�/=����jo�Y���'���D-e��[�zv�«��6Ja�PX�c"�w��X��%.qIR���_���94��M�A-���6�{;1���I����3#�}Ζ������p�(�i�U��e�z\aj�r���q�����*�`4��+�u�|C}�����U;rv����ˑ�S���/}�L�r��ɑ^"�O�`r��ݻ�&c�7(���
�um��������&�T:�5�!OH�*Տ��"/h��Vԩ]�[g���K���Fl��ӕ�>j�|�v��������q]P��]C��r%�j�Tl.s(��Xw4:�5ُTK��V%A�l�RS��66ݻ�&W
���]u�Z��vlW3M��6[%�"�5)�ݗ�Y�՟L"��N��r�V��ݥce����bs����1Q��a��$��9F�6�]p"��_�������b֥�fn�ӛ�Y�TjE�7�5��q�ڹ�~����B�ZR��q׻^���c.�����-d�b�珡�S_,p��q���b��5ڳq3�;�Z��C���^�D�Q/0�y��.m/�:�K��'�}y�e�����JM;�I�KAN���j�9|_����s}��]�T�>�X�݊��[��w���S��#���l�^�}ј�&�*"{�oL��U]Fvt�'c���z�q�&z��|���ok�7������|�_��r�3�b�����<��+��Q������i��:o��f�y�V����h�Ꝫ��nP����ʨ�������ϝ��_=���/=2�|S�q(�7;�z�	��}%8�|Tj_b���Ӹzˌm���INb����n�޻�Xk@У~�9�D�G���0gI�]�GQ.�̭���k	�-��׼���Vnfh��$K�᧘�-"x���jY�y�]��z�3p�Ν�R�)F�{n�M&\�ʱv#���0���rW^�ރ�3�M.L�-�5e�d}:�鴥<����^N�*��ThZA���-��}�8�(�G��bg����T�Gl=��:�v(%��_v��4��+�0ֽG-Dg�l������|]�9ޏ��ڋleD�J�=���f %�������3� ��eVk�u����-�z���ʉt�B!O|����όV�����|���;j�ɕюs�(�p�m�S�sc��F(�p
+wSS�^�j����Jܜ��R9Is�M�v�a�]�T�;���t�}h�@/�u��9)��g-���U*�T1n��Ms��r̮�����$��~��|b��1gz��o�U_���d<S�y/Z�!��B�y=��.U���jځ�	���G��c������N�Iz�wK�Ҁ�y��|ҙ���o�7S�[�S��_��J���=r*�QH:�Σ��獇��7�H���0����Yo�%�؎o��u��9�ٷ;���EX���kj�Zm|�5Ҋ�U���Ed-�VjkE.]�4aM��K��5�����Y}{��R=,��T�-�8C|��R��x"��:��n�*��r�j��]��fcs&T7��#R
	����&hrxxr�q3z�gWn��s�k��^��G�}Q����^;s9����luaQ7˅t��ϝj��t>�
nz<�z�}��N���S&t�Lg־<��į=�Rwҋo�è��#�Q綰���JmHld���-�yL�z}����
ayFS�]�y �Vd����8���n���Zm��:On!M�B�<������H�Ü�aj~�=]���o4�G6jwd�ƞ�k���-��4�n$$���d�#2�-�k*[}�Hf��J��ATJZj
O/�x�g��6����黁A���:�IX7e�P��k�E�s��Q�w�W؟��u�o�>��E�.��иʀ�a��{	\�B>��KE|��]kM�>��||z�ޫ'I���l��8�����z�ʂ�f�ʫV�9F.�B{:0�2�ܚ0L�c��j�y�/u���a¸�銅l��:��=�%�+-���E}~�Z���2m�'2v�I\�U�����-.��q�d�՗&��l��v�r��u�-�tc�L�l$L6�d�S4��Y.^�o�0�we��o����0�&7��c&m���̇�{�ތO��ӛyS{T
�Ji78��wZPΜy�lN� ���!��W\:΃��C纭C���c{�}ͱ�:�'�iY{�L�i]= l-�y[y���'��:G�7�M}��׍X3������("Z�y������a����ڥ��>}��
�H��|�4-8$'�����#��R��s����t1�8\�X�n�)Q��_9��&�	Z2����sH�h��%���Q�&�X��з��v�uet��.���h��6�}�RDs:;O��R�L�U�Us���0)�L��j0�%],C�p�Q:XVAn��Q�:���V$�6�ɒ�=`�����'m�knS�\�:qCf9�r����w`FV<8�a���M���jm�[&�禬Sw[!�!{��i�T/"2���vX �Mq{�w2�.��]��v�%y-�vq	t�@�
#^��=���N��f8�k��,a�좰���SB�
�հ�m�v�g��l�
C�ԺXJ 	�^��),� {u���4(��+m-�Hy��\q�٧z�S�k�	�̈́��.�G�%]z+��t�M����4�%ngtQ�
��#��A�؝f��6�Vm��\�*��[�t��*�c]:˽e��0�.�X�K�=�� <������S*);�T���Y뗎�^BF���&7�䥿v��Vţ��ݳuuԥ�pLt[�3sh�ӣ�6&mv�¶xm��ױ�:]�Щ5RSn�pv� �;]�J��zӒ��@��P��w�X�EsA�5TW�ؔ�t�J��	�p.:h���SΫ�&i��.�X]t�sq��J��WSfb�U;"�u�@;��\2NX�`h�u|r������'@*�� k�d+�W��3�[�IV�n��ڽ��[��ϭهǽy��|ˏ����aR�ѵ4+�4�+����c�TtE8Do���̧�+�EiG���(0�st!��Dd�tmJZw�d�����UB�&o�f���C����Zx���j���wҚu��#��g�-�N��@�c��*k.�����5���wHQ\� ���,�&N`�,.;�t�ݠ-���'k���n��tH�bޖ෹/\���%�x�Tnh�<�X▖�Ve�N�[��x%�g+��G�t扴��P���HZ��r�vw$��Ja;���!��ޣ]�;7_F�m]EeL��y%x 6�*ܸ;�C/,E.�\�}�
n�s��GQ�9�Ro:R�/�ʢ�]�5�,�Pms��oWE�����j�hF�}v7�����+b�c�j���ՠ���wL���..�*v�~��uk�'�E��8_ ��W�wy
��R�tP�����k��
(^��w��s�/?��|��<ǟD,���Q\�*�&[nf��C��a%Bs��T�\��@�Kܗ+���j��q�0��R�7	G<sBJ�wr��.]D(�FiU(�AU\T��-Y\*�"DDZW*�{��Ujj�Ҳ���r�@��]2R�aT ���2��0���vV,��$�U�j�r�N\.�G3���v�EJVR��Qjd���d�,�W*��$#�WMV�B�\�楥�CX��&���Vjy.�r�*+�R��*�ˡԪ١&�qDC�\�9���\�p�֜"�:t;�qZaꙖH�9I�AE�'"6fZ���稝g�x�,��r霪(�M�j�ٝ���g+�"�(��K
(��V�D*�4B �DK�:��U��Q.J�u�/:r��S���(�!���PM8�EU�4**.Rd�D]�<�{�{�� Z٭n�wIbr�	��ќTU@�g-�n�S^`f$N��'�(~V�-��Y���E�����ٞø7������l���߾[�T'�5�_6�]�p�L\r�>�J����Y��G\i�W,������W�n/�S���Ut�t��f����Df�ӻE��17�hL^o'>y���eݔ}�IN.Λ��j/S��H�	e�r����O��:���$Zꁘ;�X2��N�r��)����ߣ��Q��1@�ݖ��qA+�k���?�\���ߧ$���US�o�t���bᾨ%�Y�l����3�O�Iזu=�:�]�Z�D�ʕ���z�'�7b�zF��iPȷ��y$��t�\��O|�a��\����s�a�k$��)kkyVU�Q���u��B��\Bm�îzv�.ª������M��{S��=��5���4r4����>��痎��jOmM��ޚ+�W�陫��^&�
qh��\��)T�{�	;q�یp��Ƀbn�)�se"`���'�ȥ�����k�
)^P�o0#�1 ���u9Gj�*R�v�=̺�C6np	�����A�4'j�%!Q���ņ�Gn����q��R�� N4�	���.F���p��K����۲�
��eJ�����b�p`�DD@�Хr�/Tu��N���x(߮O�#X�=�<�y��x{�sVuZ�ַ�M�l^8��S�SH�=���f[yW<�m����3i݄�8l�#��Zg�+�,��D&�9�9�!Lt�����;yeg�Y�MH�{V,t0���\�^�6�sP����7	Ӕ�b64
�J>���$6$ם^z����'9��R.�����p�[���DEV��>ބoN)�����T����M}�����mT�,p��q��h���͵��Q�Ԃ�>�"y�{�-T�̣;�~J,]�5�c��`u=~Y�+�"-�T�t%���K��3���4,�Dk?[���N��9�z����j=�j�OC\�Ыt���q����_���c8�7Uλ�Q��as+�@����A{}��pO��k�)��Խ]��u�Χ��m`̯��|��p�u9ѵ�CWcU4����̤��%��뵑OE�I�ӛ��x��]�_�G����8t(�Z
�9��澮����$�ѝ��g)��K��oXk���#�q��݉�r��Nn�m��ŁQ7��Z�pH]a�Ъ������$��Rꕺw&����/c���OFs���Q����O�����u۶�u=XzdU��+�;t��Q��u8�Z,�K��e���!P�7������;is���H��no�������Z�n+�����1O`i���� Aϻ�pvm���=����om�|�XK@�*ʤ�Q%�J�e5��vk�Gv��s��j�-�6��

a}�0W��]p�/��͋�ں�o��u=H�N�4[쿹�]�/:�R�+���Ƚ�{K�od�n��dmw\'֞�-�z�<���ʗL�R$����ՉQy[��Dm�������/��Tb㜚Pքô*y�.d���M����_2�},�sR�&��N�#�	s��@f��7#�k�9׋�[�a&:㔱���yV��B."{OW8��zI`���z������Xf�v�K.ؓB��x\����{�VΨ�]{��$��L�Q����U�x���Ҏn)ji��	�U�s�e�m9��T�sԘ�=�X���X6�عoq����_G4��].�Ҹ�[��*��A�ܻ��*(̏D@h��ͧ��wW	��ۍwNV��9����Sٕ���_�'P�R�+���7$O���%�߼T�
it'2�Q�c�Z��f Q�Yr�����#'�/C�<{�����8|��x�;�v�����X�s��⽄o�A|��ٞ��yGZ�/�������^��������y�'@]�z鞮�<��GZ��PU�@\�&�*%1�W-_4�\�sU)���p��#�a�98���m��:����C�
��ީ��DJ��]<����)v@.�:=����ӯ�g���K~~S���]�~�
g�y��S���Zy��^
�yع"&�F����m�ä��]eW�Z��Z�+��<^�[z�w�⚣_boo\5���i��PS��;�l��6���-I,��:��M����%-5'��Q�3j"������9pF-��p�d�N�n�r���;Pr�K�*���Dw�0��X���^�Af�^e����Q�ز��VU����Eq�y9U�b���tL��bXsen5�k���Wr�iur���KB�sdxrRo��P񏴮�]&
59[�:Wi���c*�
oP��ܽ��~�_×Tb|C}����=���l�fm]�P+�`��l�\0.�R�?w˦3�]lO>��s���t�-���xٓ��;SI��+�EG�m�dt�Ѡ'�V]��^�x��R��^Hi'�؞��9�o����+�������+���0V�����F6�����'�^/Vl�[Ⱥ�����b[q����|*&9��U�1��y�.��2o���܌���I�%	:����c�jr�!�1��0�v�X+j�k��Ff�J̩X��V�ە��9K녮�E�Gk1�*�� S])T�_'�a�7�_�����4g�O�r��^ȱ9����]�{��,JDݧΆ�=ͦ�\vʂ�C�Ss���XT= n"V��ZĒ����>u�5�����]�l�������xz�ޘ�YB���m�WѡX���R�Y�:�μ�|��C��?!���R����ng\�j_5LƲ�����P�7E��m,}�D�*����(�İo�á��x�t�eoh�B(�>�TfY���eRI���ͪ�f�t��m��g�n�S�It�F2�up7\��V��u�F�M��뇍-��yNk6�ʡ5����x���u�E���Fq���|C�Te7�p>{\$�Z�M��u�l���V{p&5�����o�9���o	�hy�8j�c�����[#mS���G�K�k�Y1�����ʢJGHy܈I��8kB�m�*�Gf������F��Rq��'-���A�%��һ�S�br]���XڀﳕNe���qE��/��c9V�/���-ǻ'/P.�ԔL�b^��>�I5�=�6��L0Wɱ���!Lt��45;*�RRm�&���|^dw��U;DU���� ��P����deN��7R]�vz�qx�Mmvxrg(��+��R�{+�Ꚉ�v�v��I����Yg%Ak�!С�V�@�«��0�s��w�>����]��P� �Q��)�^Ɇ�V��8=&����xq҄�����䂱�Y7�'�*�l�.�Y���+u��f��@y=.R�vu�Kp�fO�̥�Y�Ԟ�30y���`��bܼ �#��Oa�2\����\�V.�=�Dn,�ݪv4����ѡӋa��1�n���8�^��)8�'���Z��e����OdΛY��<�w�5~����[k��$��[�v�گ�n��:-�]���v���ZI����ޔ�y�])���s��#*����������1�8��y�Ȯq���yu�'ʌ}o�)���R�rs���:�{�v��9aUէ/Vx����Ɣ�Q���k�/����龸u۷	�p�:7;:�7S.)��mua������\�D�]_a��9�p���t�ug,���'���k��q�ˬ�Eh0y�<���uK�s�Q�a�xH�g� t�~�[�����)�AW�(%�f�T��;�|G���K����;j�OvwP�8���oT5�����N+������8*!�M�]Gx�#.^��71�R{��B��x�dF�Ͷ��K��B��y�n�O'<�0�46��gѹtpK�m��c��峖(����\WO+��Mc�N�]Fn70B��Ѕq���ma|�f�ZG�S�W�P�'xq]K@�}����@ӵ��c�,�&K-��Y�q��mB� ��=��u9*_<i8h�������S��銭ǟt}�[Jý[�'�-�{.���Fu���ä'����9�߱�����"/j�rg.9\�V���
�u���ΰ�R����ҽP�.�9��*Ձ�Q��)��?^�~Ռ��xh�j�^�zM��k��
�S�)[=���'"Sɬ岥����,ɫK��u8�ʦ�g14ۍwNV��&9��<���&��f�6+W���}��Z��%���k�5m@��D>z����Z��/����qZ�'�!����-Ϥ��E9��}��s���==ڤ�'��Ufn[\��{��^��~�1��K�oQ�?s�2�_7�s���*{]Y �`�(�;N���=���G].EC��o*��U)�������-6&;BH����L=�u�7�=o~���47Y���a<>/>2�����1�Fef�Ľ�V���w��8-�eGeH`����ZFom�k�L�w]S9v������I)�*����wb.���3�R�g�9Ջ98���U��CV�����8G�r�ՏWaBk4~*]���.L���S�I����Tv���{�v9�䠫ا7��5r�w�+�9�Z�r�����b�������4�A����Jb����6��y�o�YS�n Z��=n��NH����/����j�*5���e�8[P�{jm��A\�k��X�9�o5��F��k���)i	;�k��Y�w�X�B=}h�%��|���%F���T�`s���>4[�O���L���WSt{�<�XT!}3��s��Ld%���˫�\r��npJ��卡q���������Ю�J���m�d3q嫹�t��D��ECov��e��)��Z�ջ�>sM��a��)����u@���)M������;}c�u&��{Q��������bi���?y�S���km�h���f����]=�X�9��-d���饩:��c�-��59�{��J��׬ш�(�pL⸺ɖ3��77r��ϑ���3K�"�jYJ�8rI&|�,��i�-�D��f�<*J�}�v�X�Q�R�J��ؙw�۲������^����v���DWU�I��]#�[��pIM,lj��v���Fu�l��h���L�8�����R��*����-��\v8<�JR�W*�������rք���m�?6�=r��\���h�nM�*��|��j���P��g.|s�8IsY�:Osi�A˒�:���Y����-�z���Z9��§���^�'z�<ӞK�s��t�f�f��w�wY�m��B�;֯+J�uz:����i��������s�oa�� �/g��fk���.\�I�_J����������\�ʾ�ٛ�'V�I�1��Z�F�RL|y��r{�&_+�J��io.1�Yq�m��
�è�n�����u8sz���}%*�����j�ᬣiW�/�}���'yZRs�����,㔝7b_o�����]7C�)92xF�]P3�ZQ���w�����'���2�R��B��zL3�KFG���u��T.<��73	_;�=ޕ�b��L̡�N�šb_�����N����u���
���jf�6Y���VX�V��tu�h0R�C��c�ZR�Fn|��pP7��qcy�c� ����*�b�WӋ��9Z�B� �[�������"�oL�g�L.g{p�N;Vځ�1	z�*D���b���p�А6�W���J9�n�)���Y[g�Vu�V���V��Ҁ���Y�ꙗ����I�/k]�e�2�_\v�D�of��b�s��xk�<�+p�n9�=��{}�e[��5�,p����6�C�`<�3L����@v���N�cBJ�W��U$�MG�T����etV����6�B&��3���!c2�SC�U��i;���Z�M⡘��v"���
���. �X�$�g=] \ƭ��De�-t{�*\r[�Au��՛j��a�Q��eN펵g4��R��ާWE�7�I.ȸ� j��i�+z���:8fZ�D�Ṧ$'A�j��2iRe�V���d�L�x���h7uf�I��� :͙hF��W=[�e6N����N����;*<!ӧI�v��+H  n�*�VŶM�*�aI���P�ĝᦗ!��]ä�5ݥmoP�cs&��l�+G�"�.�T�0�0�R�S��Ѥ������S���;fr�N�����k{nM�� *��7{3��i�Tk�q,���'��ΐM��öeՐ,�j"5�⊠��E��-�;���|���{����`��%����9����-u��dMѽF	�G��s2��l���V�@���ID*V4#��d#���Ũ�%�0��'�tv�A\�y�l�tYU�B���� ���@G��T�:�\���6��ʎ�9�?B��W��Lӂ�ey�o\�Y1 �,N]f���v����WF��۹\�1ޡ�Y�`�����`���s�ޥN�L�E�e7nR�	�;T����~���hH���geSQ4��m�\���n�<)<��&�32�K撼�v�'�d����U[�K�`}�k��D�v�j���Ie;玘�\��jh�}�c�L���w��S�1�6���cz^��Y�3 |�J��ި�������n��3��lc���d��s·o����4
�,��`����d�RKpe��@9w�8V5ۙ��`����[��mAY!�[aI�����]0�Z'+׻�K���d\��0�����0Wv)��Ƈ�ks��m9(���Rjdst�z��ː^˹Sq�|9S�����Į�Tʗ]$,�#&��K 뷋{���)�D	��U'A���QI-���m��R����ʚ�!�p�΁S1n�)�1���S��[a�I.;��fTh��u"�R<��S-���\nM��Xʼ'�8+xH�N2q�fYf�|>Ʃ��	���u��j÷͹k����Vd����N=ԝ�(���`@
�J�]3��AeEwǺ(��]�S5;u�N\�U�T\�+*#�ՑRq�#YDr(�XIJ�FIkE���:jG,���"����P��a�UG9���t8TDQ��QfU�EH����"rs�\�*L�W��˔�Nt�{��T�B�v��8�*��̴J룅E\����r��J=��r�R�{�RdW�ąi�瑥Ң5g�DUEy�i;�K,ʣ�*̻���̭VT9�9�I#W$
#Α:��8X���wK<�E��	J*��p�Tٙ^�ʜ �N�"��G�n�<��wZUU���f�UE��*�St��9�ϟ��.������u��=7ay��-��ʹ�3�d�7Eu�Xm���vշ���uL�e���=���𝜹b�	n.Z*r3��c��)�aޥ�`��ʇU��vTC��co���M��u�ǥ�㹼� g���W�9��\s�5hO��l�Jv�����=�u�Y�kjs�}P�z�Wd����E���M}�0�q�܅��ƫv��\Sk�,
DÍ�;@��W���)��ًky��N*Q+b����Ӕ�Wdr�L�'ԧ�M�{��?o�M[�W*>�|z{L�bL\r���Yʋ������{��>�d;i�TCB����E���i�GN����>W^I�x�Q��&����>Z�������������P}Ӥ虜23���3�=�\���_N���'-�2�\)z�!:�}}�s�dAʫRa��5�4pe���nr�C�¢o�
������fK��M�X���k!���yˊ��ga������s��ua�ׅ!_-M뵰��ѝJ�u��FV��o����.���M9��<�FG/0�?�`Ф�I�r3�#�	��dj4LU1Z���.��+�i��0K���;�Y�u��rk����{|�c+;fJ{^K�qV#]�ܺ�7v�(�_�3i��/k�#�b�ԙc Q��y���Y�+�C�axe9�?m���nY�8J3�rK=\�<�m��Ol��
b���PC�BTw���kE^4�#�T�h�O:5��uS��O�������W��l�uH��<Sn��]��lm�+�M���o��9�]��3j�R�+Z����sѷ�qJ!�K�E�0�I
���]_b}��m+��V�'�+�le��'\("�\��p;_.ସ�6_ϤF��j"V����Wظ�G&��o�5�h��s�`���5�U�B4�fx���
�5+rsS�H�Pb�t˱f$�	�|�V��5��q��
�~N��l�D����0{!_�=沔��,Rji����T<������5SK9�m�>
r�\Y�g�-mn�f��Vم��®�R�1���}�W���V�'\�Õ�L��EJ���o
\b�ze3���7��V;�!䫾�$�F���eK�P�nsP�;�C�/i�Ov]���j�UqRm���ut�O$�\��̴r��!f �"�K���T��%����9�J�F�HY�8j�[%�k~��6;�Cw[���τ��j'>y���gp�{�w?Wە���/�8֣��v��Y��Nn��E 6�v���fQ]#1�{��eg(�������|�4P�3�<�f�N:�C��ZU��7���a�X3��=�z�W	Z����`4-�L��#������j��{�zs�)��m��M���������]*z�@S<�b��)��I&�!�j�%����Vu������~�
y���[�=�%�L��|e5��+�د���6�C���S}P�ʝw�S�וC��bo�ck��.����Rs��X��5��8dGz=LnF��=o��ݐ��<�QRu��򁞃�<mB�ﰲK��>~�E|\��-]A��y�AoՁ{'����4�xo�;JJ��A���/`,�N��\�k�DUa����G�x���:��%}>�������^�*���;���u�V�CuÉ��z��US�d�@ ��<fu��/��"�h�i�R��:b�
�F*ݳ��T���"�����~���>�r��̘8�f�Žա�ѝ��2�ڔ�0-��P�gkqȃ-�ݸ�����Pi}
�qt��Z�>��L=�v�ǳ��s|��tV���mfuR�s43�)�{g�ѕ���A�h�<��3O�����A��x�mh7�z��Ug�\9�X�RZ�=$O��HR���ҋ�މ��"g;w��ᱸq�kF��5~�q���<s��|`�W�E��}*l��^�#���ۀ/}y��ou>�>�蜜�B�J�K��{�^��y]ы�7�4oޟ@�`uRh�^���`�y�S��Of�U�$��s���O�ތ�O���m1ܪ�0ߪ�y�:�x���QK
�sz5���z%�GxeH4���L{�N�u��7E��wSm�	�y�u��oJ9}�f����%�|,ס:���ȏ{����܍��r�qGv��ey�/IӨ���P;�w�J����*��B���S��u���np��rNj�N�L�#�C���i�mz��
�;��>�4N%@�Fy��gΦ���\�ߟ��,�Vqz}�<9�;q2�f�d�`Sbd��G+½Տ/�;�;G��)	M��^�p+�^���}S�~�qݏ׬�ǹ��5[Xu?\� %wkQ�'��@Ϗ��L���V�#˴�`����ƿO�yǮ��[���6�A��FE^$���w�>���;���}�O����S/v��ڛ���\4�YdȎ�Z��}��ز��k��\P�Ŝw�e�R��h�PN�}nk�F��U�盲��c2}(T�kB��z�Sw]�1��YG�ĲS{:���'�仾=��ޘ�J��^ŵ<hq'��{Ơʦ.*e#qU>	�wB���z3}�w��%@Rw'l���|�x~�m�|sՔ��%���$��0�O�ʡ��e�u�HO�[{q-f�����Օ �1.Tw�g����7���S#:!�����!���D���KetW'�3�d����������ğz�*�<W�0��z�ۏ][59�Y�PGS x�.��T���V�a�b�\�#}`���0)�:ԡ�_��}�m��OC��߮�ƅ��K'���3+g��9��v�/��Q'��B�=㰏�Q����x0ϼ���N2^G�F@ٿx.�!FF����g�}�2��H��=f+��W��Qkf�K_sw#������^u�}u�:���������>����<�]�U.Oh2��**%�n��+�v��{���5��eTWv��`��r�^�>��긏z�d@sC{�u ��������[��������#R�kn�s$��v�S�g�.��y޻G>�ޠ=F�3�LOd?vX��9t�F�gC�w%w���.�{kT�7�V��kM�"�Ʃ�gg`��滀�۸��+^p����XU�,�oIK� h����];�e�t�Z�U��Tz������݀+��*-�Ϧ�7R�W(�cg��wOL��p��w׃+xXk�5��˸��jU��;��(�0�*�a��|N���Wm����k�c>O�K�>�UxOg��}���ߧ|gK�NZ���#6��N�{����X���(迫������W	�?d>�g�?U������=�fSp�E��]����e�'3�ae	h�qY5�✁�X�p#����u-��VNh��2V�v5㔺Ñl��=�/��nQ�8JVf�=P�T��9��5C�dF���K�}35��,8�\�\����^��ǞEz���u���5�#��<j"J�2���2���_��A��~1��UQ��]�D��{�U,8�O���\{�s�[��yh<�p�Nxz�e�S�ũׂ��g)W��9�����[1��)q��hO|�߸���z\o�x���W��Mg���Y��9Zg��N���y����|���U/�W�HM��ֆ���>.;�4��{�o���0�hv�ù1�޹��k��ȯ9 �dH/�$Y+�ra(��C�D����>ζ;_�����+:��~�3���)p��S�q7�f��	��]F����p*��Z�/���D�,��k��rES��o���at`�z�V�Ȓ��K}[���������d�n��m���N�ޢ���܏`��� ︄��&U�.I�X�5�>���w�FD�$ۮ}A�,���0�;��u���+ ���E�Dd�)j��ң�������j�vm�Ve���'�� ��
px���h��=�Wg�(Z#���FC㕱�p�k����~���w7�N���qp�ӵF߽H`�x��6��߁�9�>Gb
��謰7�`��iD� ��g���t�7���ڻ�kg�&��ޠ;����PɓP�S_��j#{��D�6$��G��0���+�i�W�!�]���7��?T��*8f����k�LZ�='��u����Oxzc���u/N���swi_mކ1:��ϵ����o��ef�x�~T}���u{�����3�������0�謯q��:ޫ`�*�P�|	��q�z��M[���؞��=y���j�G�m����\ X�bUj�t�X/�,ua� �!���r(�;�'�;�P��=/��Dz�9�ϟ� ��ms���0�d��:��������_�B?���Y�v��<>S,z5�	zW��G�������;�{��F�𸾒OTL���̘�	Rs!��>���-ؿT�s�n^��O����G��������dz�ǻ>sX����,����gv�s,�_��]�Q�h�o�mrub�V4�� ϝ�4������&Qx����Z<rQZ(����sY�5(\s���2�8��vʝ�nf�ŊF�U+޻��d5�\59+���>t����Gv$��1q�햶��� jm���(�X���g�$�Cj��9mՉ���л��cw���P�s��1��t?	ٻ�p�F7�.O��$��,	�R$Q����Lu7�$\K~����Vog����I��A�W�ѾZ�xY~��!:}��G���l��À�,��YT4o_���}����y������e/�~�M�g�Do���d�)S_<fu����/T{��Tl5s�u�k��T|��F�z�. �s��w���������2K
Ijt��]tC3�����5Vυg�W�*w���g��kF��W�7���};�}l~��"���T��ܲ�o�C�wE�/bR�7���
�TN�#B�Ҵ����^�Q�+�1i�Y�q�O�w��\���w���B�z���>,��vK�@���/TK[z2��M_ٴ�_+�7�	�:�u�r�~���V�7���yS�/y��_��+M�����d�0���W�t��E��gu���om����7^;���2�7c��m/$|ۡ�Y��g�����y�܍���;@��6wj�ey�}���f��i�Y|0��kU{`@�`���@��Z�f����/!���daTv�Q)3 ����6-Ģ��l��׾��]�L��c�O�#���=� e5��a�56n8��{���H)�e�7�+mR��v#�ժnr5��)o���g`�u!�i,�*g�$�{�\=�q9�^�v����/�G���w!N��o闆��t9�B�l'�{%t��[n������@���q�u4�@s��yC��$���>ɝ	Õ[��^E�W��*�weOxbN������>��Q�}�,q��
�������^�^�Q��X�I��aL����QK�]�ץ}p�x�x�uL�d2��3C�C�z=(g���(���w#�s|��wqK�9�}Y�mK7g�<?�*���e#qU>	�wB�>���P�#�Ez�fe��X��Օ�u�?[㎲�qD���U�O�C�[;]T��-������m�ۭ�Y��5������ ��{UHۏz����6K���9MD��n�:�n˯[���L�Z}���}j�6g�U�޴���C�=y�Y~��j�s �J�N�ұ����{;{BY|��`W�:�l��V�HvK��c���<s	~�A�UL�\7#�M��QhQ������ڒ1�DL��кs�;�O��j�m�����*>,�q�Ҙ.�����؜����נ��W,^�<�O�U�.iq�3,M���v�q�C/��ٚs٥�)���ՈS�`�{�iL kd2�����`�s��@�ڸ\�5��#\Wm1Z:,�H��r��5�[Vo�*R���٢�r<w�L�WҜwM�yEPv�l��&J����x�&џI�2CWz�T��Q��Moک�\sw#���wC�rc�����˳��ޏg-�Q=�>V@wC�]�U.Oh2�ȉ}[�C���ݸ|Y�DiOՔ���T�p2E{�;��X�CN����P��z�d46�ї ��V�8����W�t��}�#.ڹ=��͑8�;�a\}�q���B~�G>}��o=t�����9���,�v&�ϛ��K1g%?w޵���Z�- ��>�7�\<u5�1�����Do��'���o���в/�����V���R+X��97��ߢg��:���Yd�t�nydxgΩ� c�_2���P�sZ�9�W��z}ڭ;�͘�̩��	���>E���kM�N@�4��N�"�y�<g�O!g/��P��ܒ�����;�G���ǹ��	L@;�^������.��߹�J�$��\\ՉQ���|���ⓝ���<�hxv:�B�ʑ�<I�RW�DUA�>�C��q��Y���{h�*�=�Ϭ�I�Y�������yh8K�<	=Q2�_}~�u���A1��oθeb�۪r�H4�巃t5g��A;�{y��:��9
ZX���F�9q+!᱒�=����<oz�DL]����1��1�{�g&�<̈%V7/:�\�baznk}o�"�{�94S �Å-q8���^�t}�%l]�fP��hJ�n�X�c�h��z������T����}j�sxM�ejƬbn��n&���#�+��hRθ��rԠ��/qL){��؋iv�OE��mQ5�ړ�f>5$z�u��sr����f,1�0�n]�J��c��݌$*7�ݞ�k�N�D7D]r<)�Wί:�T�L�,�8��TlNyou��Vo�4�mG��q��NJ̗�Rؑ�4���^��[V.T1��>�&w@��kGT#��P����{��}J_>���-��)�Z@�V����u{�b�С�ЀWK�U�ֹ'5�m͔��t�����/��kK�h����J�]:�ZHH�7�8RV&}� �fd+�~�wM�/)�X{�/�ӯ�s	��n$@�l���,7��ԫ�K���7����"����4X�ë�=�E��
��l�ta��d�@�5Cyj�3�Tp����2A�Ԛ�uڱY��Xh]�n`��(m>�/t�z�)�J�pv,�
�/d�����xP��d�	a�dl{8fn��7��8�D7���8{��S7ẋ�Hiۙ�nHE��f��eݽ�hjR���Vs�v���Y�nw`5�ָj����RGfi��2S�.،�jw�77�ҵ��2����b�.ƣ�B�d����f՛v���r��woH�6��ו��Uk�o�XIL;:��\j�=� ��&�7��'g+�oD�#M�C�
w�a��oos�ڕ�:4t�^\s�mۓ���YkÜ��L�r�e��Ã+���u���AWD%�v�Z�@ג�-�1��p�`�K���ucB��V�z�:�J��I��Jzr�Ab�!Mpw�M��e�V�t�:K=�7���Xp�v���K=g��M�Bf8ܚ���"���V�q�soe�������W@I�=.�F�Gr��C�}\�/g�[���]ٝ4�zb��L-N⮸W�Ɏ��^��NK��7>qu̧9�6��6Ź*`���`nG|�f�J�� �a�ӭ��6��ˎl�냟r�6t�_wmnu:�� � o��2�l�]��c"��]n�$wM���ta�%S��F�s�о����T��!��P)*�Y��7x�r�Y�\���[>s1�4�\N���t������8�p����u�8�$�We[od�X�tڣ��ȫq����z4�ra}��঺�$�nwS�gD�;��r�e�[�N�m��ou���e�|���^��{�Y�S���ٰ,������X���"���:�e�śVn��X��v��Fe ��[��7��^�9/2N�w=�)�yz��q�
���p�R-k3 �;���G)̥�%�ȮN�T��TJ����	���:Tjy�Ib�#�wM���(�$,�̴��s��r����u�#�%�U�u�\(���ȗB��N��^K��Q9�"�kh���!3�'"��g�yZ7&�wws�&r*wJp�E�ʅB��R�ũ盭3���x�Q��.��$Q�:r9�'gtnNDUW�u=C���]P�,�M�v���ɎT�T�KG]��#H.�`���ܪ�H�%�"�I=q�u;���]��SKMwC�f��뺁��䁨TQ�H��(��T��۳g42SIʹ�eJ��RXX����i�7	��$"�M,�B��B0�S�"�w=<��M���I	QE�g�9�2.���z�?;��w�;,7.R2T�:7w>�+}�i���Z���Z���A�u<n1��L#��Sj�C(_3h���\�;��n�j]�(g~��qL~��M��n�M��߸�GzG���=y�p��o���Y��#��Q��wwt���־�^�(	�t�5�+�Pȵt�r��Bo�����h���{=ꃑh���aw��>1�'ƽTdH-����3ॅq�և�'�v�g[�7'�f�I;�;o�j��d�����~��	g~D@j,�WQ���!L4����⩷�����9y�e��@�(����ɿ��V�~��E[���#$�G2_W���i��7����*j��$��O�$j6ו���z�>�� 7���ߟ����=2����h��5�#Ӈ�޼z��ߡ�o�r��ϸ�{Q�������^&���z��dT6�C&M|�R_�sɹg��م��}��`�@s�\T�:/���q�O������7�cz+�n#=.�롵�:=��7�v�������Њ%�Ʉ�ᵣ�}�ӝ'ov�����c�,��~��'�}������<���e�=��b�~ݺ����q��;��W��:n�`Z���������?�:! T̓��a摲^»)+2J���d|j�h�+]�9u�Ou� �A1��.�1ǯ� j�̫;�X��G]���ֆ6+XR��r
���S`k��cc��㨻m�_!HO�w}�gE�݆:5n��n˹M2h��]� VG=�,[��.�V��Q���\��g�Ctץ�B�XH�l���#s�OU^�P�ʼ�D�4=�[��d<�y�ju�yh� {�;!˗�IG������H,�=�/��d���	Cl�@��]Yr�Hˇ]��e~��)��!@�}2�+�o�
I���o�����+��"���S�x]��x�o�MfAg�g�N-�c��W�L�멞s�/M������}�|}�?O�W��{Y��w^l�
�����V�}����6}��π��h�u*����'4�М~��G����zv�f�	/<*s=�����9��Mg�z(���$���`�ŵ=�����"���z3D+7��Uj�d��{O�{:��z��������ǲ��d@�8��J�U��4I�yT�^ָ�{�ҍ��O���؆��{a��q7�Qq�b�!̗5� ����%��R��Zբ�ɿ+ ����6k|:��q�F�n��G������������d�_NV�f��Y��޽����#ӛX*O#�7�3�h�o&��n=��'�>����� ���:��������(ZSe�<��҇m�+�g����'� �sŅ� ��=�9��֑yV���g{uF��u	��[R>�S8|;ou8:���c+�],E0ʁL��ޥ����蜹���n�%��yvGd@5�d��l�T�]�9c_f�c ��hƤ��"��Mt߯��?�PدJ�K���^��y]ыM��x��ǻ��'zf������B]��P�8}"��ʓ��=��a����dS�i��cz9]�c>o�t2b�$���+��b�uԮ'��eH5�O�U�ɇ�wL>�V鸢������������N�ѱ5��i]����8��<j��U�=9�V/�=ۑ���v#�v��}Y^G�7z���S[躁��<����D��JW��ڿ3>�yz���/]A�v��{kd�)�t�.��ǅэ�8Uxo�=�=�^aM�񑨞>;>�Q����&{�.|�/���/:�W�wfx7Bd�zvD�ݛ��qO�9���~>
�]�yM��huyzߏ��O�y���s{��ƽ��T�lǾz�國8JWg�(���ϑ�rWf���L�|=Ll���*$��}�!gF�J��/Ю�M��e�x��f�T��L�n*��<���9�qw��w'p�'{=�P����<�{}@>~�=�:�A���3ĕPf	>U��g�۩�T铽F�5���9�k�мj�V���B`]_���7dj�u�'�I�����7���\r��LץԺ�q�6��O�V��3��eM'e� �S��v2�ˉ�v��!b�U-��cY)\�3g.I�b�Uu�b�Alw�I#�w�fϾ��q'ν���y�o��}�Dm�{�~�D�r �$0��t�m
��Z���@s�ᓬ��V<�}O��O�I�~=���#Og�DgG������,�Ots���1�_�����}�F}2��`�P��)h޵HvD�[f3���l��};�����O�؉�<$�@^�]禇p�$>��'�+�hK=�O��j�m�����*>5��v�8�"��-�/�j27�����)���������7E���Tǯ�n�xg��H�+�)�7Rw�{5o�{���q��3���0
~���rz�����TT��Ӕ_�խ��[�	���٬�/BG˗[�����}@:��z�g����ї ҟ�`|w㳁���_�x�En�*���{C��~��.~��z���K��t������(��BF:6�F��Ȯ�\��c<�����:o6W��m���ϴ�'���	����?��_���n@���W4�iC�N~�e�P6t;���������T���<�<1�?d�^�eW�+���z$��9�01�������Ѿ�d��%�v; �?��h��s�����Gԫ6$��Q��5���d�8�.���Zz9�+���k�rx�}�{���Y�K5\�]�]��6Km�0`][���;��Qwv<5�!���Xu!A�K9�M%(����qǰ��i��W!��1�X�{ݻs��wl�<�>E��:e�=�%�|���RF�W7�5:o�sޝ����WO�g޺C�����(вR�3|g��z��� 5��>��v��f���jJG�`�DqJȷ����\�y8�Z��ж��u��'��>2�ݖ�)�>���^�m�������T���U0��>�a�t�������ׇd������Ot���A
��zn�R�E��}1��]G��9��*]/�n�M��߸���z\o�x��y\>ϣ�Y��ۺ��'�轍Ⱦ�d7D��j<��p K�g�L(�(R�~3�O	�O�hh����{�aِ�����r���r�p�A~�]��ȁrQP �@��I�+�s"��k���'�v��T)���UE�to�R޵/y��&��z�鸯_�%�Y@@}�;E�|}�Cy�C���W��p��v�s�!�rj��>�"}�Ӂ�q�z�M���s>��FIh��zH�}^�����V�]W^�+s��9^�H��٨��z��~� }�=^ o�������=2����+ًƢ�ɫ��� h�ϳ8����{[�PNd7���sd�8�S%��^�GG��,�)�ŉ�\8<�c2�W�.�&i����h�z�Q� �h�Y(v\�Ρ����v��&/��W-�$ջ)M���3����6����lU�y��^)�j�(s��3gh��2,��H��S�7�/uǳ�wtn��4o�{���~J���W	����(d��G����U賒н�qR�迩�xU�m><��D7�cz+�s��;�����c�2�����;�o%#����6mJ�1�p6�;���t]9�wvP�۽dBu告���5����9g�K\<J.|3'��s^2��|,[��֞'3�3PwL=����:�j� ���k�ߑ��^N�Ego;]>��U���'^^���a#�]H_�v�k8N`0���w�Zk�G_����7��[^��D��LY欋U�~����sS����{h_���Y8Jq2�a*����j�ʺ�Uˎ�V�3t\�����r������e��s�Q��݌\j���Ǡ���- ��Ex��2��3�늙���������{���N|�>�Y�q�������FK��Y��͟aXg�q ��`H>E���H]T�9ȶ���k��p��G���̺�L1�E���w_h{�`����p��o�<�\�j�J�2���H�G�ڜ�u��=���N|�d��3�rr��Xx�n��X����.;�wJ�ưP�}]z⛕��hh�Ђ��ݳG7�IIJa�`���{r���bQ�����<���f�o	Xq�����b�P�SE[4oa�]WY�oU��[�D��K��,̴��V6U�緓��p31w*;�Ǿ��^+{�4��P�=�_�=����̈���tGǥx�ݖ��4�N�fl�j��N��$O�Q��ws�,C��=�?W'=�#;�]��.w�D ��#���5�fΞ�xos;�y���}q���<��F�m?[g>>���>��_�Xz��j�s$�kz��M�Ƴ�tq.�iB�Y>��D��!W/���2�o�h�u���}��O���w�������z�rͳ���K��=$yd�sff<� *�|{Ƅ��5�/K���G�=�wF-y��8pz*4�w�-��߂�ȯ��dE��s��W��ތ���M\f�ʪ�������)�Ҭ��-%���=	*����;��Zo�eH5��U@ɇ�'tø��n�������MJ���Jtn�N]��w�z���W��ޡ�W��zr��\y�܍Ϻ|N�|"7f̺�S�~���L���u��^�Q�N�������W��g�O/W���z�_�s�ǽ��w!N��oQ}��-��3�,�m�����袙(����ǲ$�x�*u�V���%߽���K@P�K��G*!w}�$��Rr���E킜�e(¸P����gz�k�[)݅&�e䭊8��<��4��%fΎ]�]}x��#�z�% Q�]�v��-t���N��q�����el��p�i�\%l�9�ӫ�Y9��P���nFק�����߾%��x,��GE�9S{2�W��
��~>�>�� 6�vV�����]`���;����nQȳ��c ,dTϑ�rW�hydiv��WR�2�Ta�}�V�=���%O�g���g��#mK48�3ƌ�b��H�T�'���;�h�_v���`���X=�'���@z����u���rYc�+~3�*�;Y�|c�Ʀ|��7~�j��O��V�G/�n&����zG��F��|n3ʈۏz���(��C�)x6�N��|=�D���.[��Ý@�>��)��U��Ͻi��s�qߟ�i�����ul�׷.�HϷ��T���Sk �����ϣ`�}_D���\��Rѽj��~��dg[dx���r�ÅS>6h���?���
���	���"���y�xm1�]�����Z�g�"um�X�ټ��g���=����{�뉶g�iL���'��}/��n"�[5q���?��}����-Y��K�+������7^'��O��g��`�p*ӓ���ϲ����k�S��3��3fV�т�J��z�+n$���N��g �dZ
�{+�Z�<��AC��)�"�+�J�f�/�1�]�x�g|�^��8�X��:�}�1}�=���Q�&v�ٹ�]67��hݺ:ºĕgVʦ���_�^E�r�'9#v.n'��gU��R�V�Gu��G7���o}@:����}�����r)�*�d|�/ޙ"y�?v���~��hv�+:_ں����ސ=E箘�~ۡ��'&r�E��w��<:���%oA���VSqS�'M�l��Uɟi�B~�ߎo��?~�����J�y6:�*�c^��?~����|kNG�㳷���᳡�T�J������ꟲڽ�S��hw���"��[SC���z�_�v�3����'�ا yh�J[�1��V��˂}���F�����b=u��z���H_���9��% a��=P�+�H�tW�p����^�6z�j]3�!28?i~��N�exyϩN�иk*G\\�'�D��W��<ٳ�^
��w�[ڻ�ؾ�_�ϼn(����]S>�>�a�t�������z�xv}/-�y����7��d��hI����ID���P��9���&r۫q���x��<C;����f�)�,/ٻ��p�G`P:}�*2���P��2-]?���Bn"}�CB�z��G����{;�M�>��j�L� +Juù�κ�(wKg
:T��d[	��v����������c��ǶZ� ,z�1���F���Py�+�i�����B�9{9)D�@���ְ]�c�e�G[�2s	��z{F̰��yRn�]�G��a��������/�H&�`�����ۊ��0�\�j!A�|dH-����0)a_��hp�nûY����Xo9;��h��W���]��g�pt߮�qW�f�����~+��o�/���t�%�Ss�3�=�9^I��*�ۑ���v�z�>χ�&���h���0��@y��XQ��ҶeE7��_l��c�23NW�UǙ�l�m���_�(G��1��� ��ns�(����
E��(�O����Y�A���k㚲�G�� ��7��q����{+�ѿ��P��k��SΜR�U���z�����S'��������t/j��~��u��o�\a>�W�秧�)��k٬�K�^�o� �y�����<*,��6�9>Ӄ~�:N��!�ڬj{��v�pjp�o>��q�����^��b�=�ۜ/OC2�q�Jy�x����_�E����T��3ܒ\ {���:�_����z�V9]H\{�nF�9�wA�g �T2�e���9�h=��=z}w���� b��W��G�����<9y��s�U'�T}�D����8��z̓��x�af��P�(ҽ�w�d����'wFU��wR��^[��k��z`p���/�48r��M�
"�MV�o B���_}�;��#�`\=J���(0��X�7�y�Fܖ���P����I�n��E���bO�6f���W���e!4�L@V��3@��j^tLJ������WyS���%p�J��n�.V�
��{���;�o.�`�]X�b�ޛ�XW �Q������@	�"��K���E��)�n8c�C:�^�͒��0�L;��X��˴T{|`]�V�FZjH��B���\񑛛�h�ȓ]�-Gpڽw°o-���&��FժQ��s�j�4$��F��)���bw&(p�ʬ��P�x��Y͑���f����@�n�r�#��s젨]>���VWZ�Ioe��+�a����-񑚂�PM0�L-�Yuj[�z���B
]��WdJqVs��[]Y�P�S���f�5;	�X��$Y;2V-e�8�(��ʎ�V92�m�Z#ch�	-�ir��~b�R��o7k�qn����HP�|l��C/"b���:��;��0����+��Hw����Y��s�'�]�;J\�z�)G���b��lD0i��5�!�.��m�K�o+^h��lLU;M���H�ց�p�����u�F�xvw5@����7�h�o3&��}��rV�2+I�LR' F��rw[�^X0�S�j-��5t�ʫQ����*^"a��@>C
�Z�:ì�ΦƮ5"�"���I�����jEgy��5\��)�bP������Em��0mA��'���g;�V�ۓn�g$�A,{6��mɟeu^���������b�b)_���wh���uլ�,���q&�Ĺ#{Ow�ܔ�����]�HAׯW���і��!�R痽0'	��]�G.0V�Ƴ(;����[cD�K�ތ�y�8���c������q�����וա�[t+�>���٠�m�N�K{0��v�C��+��!�E�N����ƺ�C�%���r<��׏)z␥�2Q���ҷ�S/ a�p$WtE�T20�Jw9�xjN�\��r�A�X7 V���3�.�AΠ�{�e=��x�SR��]�Me�2�ۧ��n);�9�M�h*�y^У�������e�� �eJ��Ḳ2��l2���w�6v�K���.���+�]�M��]�zaH�9����}¦e�cB�bWfT�)���;g�Ɯ2�{�%ճ�����7Gp�^��VE��1���@��Y�K��WՒۛ�.Vot�E�gj8�[�ɕ���z�I$��yldAJ��*V�H�i>���\��ۭ�oD�ֈ�q9pN�.���Z�8ţ�;|N�<(�.��\g7���R�\�� ̝Ct�%�)���i�I�0+��8�'`
��R���<2ƾ�>]��Ͽ/�'v�����J��wTNS"�]S�g.r������DP�[���P�0�
9����9M��i^���C7f)d���=��2H�-$�J�R52*�Owt+"�Pr��,�U棻rr�w\�
�wW4r�N���K���u.TR�Y�A:�$��vZa��fVw\p�q'(=�{��*�n�"��e�s�B\#��Fʄw�9F�r�n�'t��NK��Z*�G�㮲ȉ=�t1���'<�wi���ҩԩDG�I�$V��Z�����P(���D��UEI)�P���q\������j�YD�U�9�)G<r�JE�A9rȲ�җ
��aE�)�s��z��7\�9Q�EZ�=��������N�+�tqܣ�ꦟ^�d�u�]�u�����#E,��\3)-��%�7 :1ֹ �[+kt�+��F))��ξ�ӑTpɪ��:���(�3ꍟL���\#{3�
�k�*!'O�վˇ��ʣw��~�}�G*e������z�����nI.�X���O��S�����}^�'��S���L;�R��Q+ke�5�3э��X�2Ϣ�H=Pe�1 �$�Bd�9v�X��~����mߜO:��ZoϪ+��j��[��g�k<c���V�`O��H�>��嫨>�RÁ�bFN�c��W�(�|$�����+�#�'���P��>5���0����'.��u_���M�	����y\Mϼ�/+����p�n3ޢ6��v�[�.k�@J�^/�ә�|����_>[F��|
e�Pѽh�m�~��Nq���mh6���/�U_�W�E�O��gۥ� +=���I��8���䉟z���|tn}�_�ƴj:�W�7���};�}�u��ۙ�'�D�k�ZC�7V�'Ҧ���V`,���+Ҵ֩zuzd{��	��y9��78�g{z�|h�)�XFEDw�YQrz(��>�
%��ϰ�f���F]ʎ�<H�n���Dd�nWU��h��L���(�R\9]��ƶE�c�����D���5	C���}�"��(ڥ*�;�52=m��vui��t�n�j���nj�o�	O�e���CB���6L�:���3�xq �ޛo���W�q�&��/G�wt-�:������ȭ7�2�>%E�{0�U��3;p�i>�'$�
�$�������om�N���ϽCƮ3�a�N?uX���nF��>'j G37�o�O����mf&�%z3Ք��+I�j��vڿuU�'>^��;�Pz�ݹ�����;[v���}K�fV��98�U�M��}N�u�Zn 6J5%��^wϝM/2z�����	I>�
�q"�Q�:�7����?DR%�DBI�}�K��`W�NG��̰�w�zߏ��Jm��ϫΎ�wC�JG���u��z���<�F��ܢ���bI�2�g��>��nujٛg �k�G�¯����Ͻt���F-��f��z��񯌪b�R"��K§}?��������*�ZYb=���{A�9��P���c�q�R�f�g�*�Á��~��"��X)���^ދ��eL�,�[{q7�Kw�+�yο���q�TF���]�{ %��r-�1;��t���r� 2d������R���~Ws�ZG>>��\u�F���z�ӛ��}8�s3������l�Y���꟔�h�W��^��Wc���:�S؍�x<��qpT����+E�򕾾A9�)��p|��l8���kjD�a��������Ds�r���
q���v՗J�wg�9�g%x���[����٩3�9r�eZ{��lU?y��P�>5���(�=끸����E}�R��m��������&OUP����\<�G��uU�C\�f�I\	 ��yM	g�s�)�w�\���8{���(5��,��Z��f�+��Q�=��D�+�/�H�u�R�:^��7L��9.��49���;�o�Gy���\��U�>%�z|���+�p+�t����Y|�/��<l%Yy]�M�ё�r���Ǹ�'���:�7��P���|��w�.AGįrDt\�_\jb���3��
�V鸣�/�}���v�\<��v�>��9�'z!��n��Z�uUWO�I����o�xjK
4��Eexm�R��7��o����S^��������X�C��JKkQ[[����)��?�g��ۉ��T��(迢��'n5S�s�#��5܌����.�ך�;���R��[�a,�����۷<r�wn�ʁ>E����,��>n_����$��y+`n� G�7��;�x�T��y�i�=�G,�)\���h9��'�	��!I6?Ud���_��O`]2�g�]z��]y��;:ŮAS�P��n�5ƪ�^4j����WEefWa
�FV��Rm@�I`}k.]�|"ڃ���IR������\S�(P�j+#k���or,�Q��G	F���s�5{
�B�緹�XR��U��� o�#MPAh�жW��c�^s�C�S��-��qsĞ&�3����Lc�#3�Ew/�>���z�Σ!@L�k�a�����I�{������z�xvD��\w�%�����ݏi��'=,Y>�U�*e����&r۫o���w�x�;�<wf���]H�>�k����9��Y����Te�!J��r�E����Rq>���g܏�+��Ƀg�bg�,�y֧ه�%#Oc�Aί]� \�j9W�@��J�K����q�Mh� ��A�v��w�����>ζ;~~��o=냦�=w늸fK4���	�^����疏z��Ng.{�f��:���,�������J'����ɸ��Z���dU��L���-��2f��zL|^�ٽ�~���!��k��<٘�m_��?z�>Ϡz� �dX|�w�yy�X�^7f�ת�u�GD����D���%��Ǭ~e^����Ϙ�s���{����^&���z��,u��缪��Q�ޞJ��?}ޣ�R�EM|v|:ǧ��i�t��+6^��W�>o�hßV|�@�����al�@��p�AXr�֣%��xm�]�ζ$�Y]}|�������:�Ûξ��-māU�*5:�w���L�0C>�j,�ɱj�OU�Pem����t���x"��l���B��k���G�rS쫻psH��ulU�
6HS�op]�L:����yԌ�*8f���*0�Z6�;���t\S�'we;Z3���!���ؗ-)����%�����|g�y{���{2���Ǖ@��ⲽ���1>j׈�E.���Aݶ�j��S {�Ư�W���^�/K^��Dyu!~�ۑ��I��C�9�׆��1W�����{�^��VUq�<�W����MY
}/�(uQ��!?R�)j���(�i���#�^��p_�ea�"�R7�Qp<��Ϡ(� lBN���c�p�\�Tn�O�<&-\X�#�7��%�y�}�$�q}$�'��&x;��)���������}���3����^5T}7G���V�C�e�!_\.Ϝ�#l�2�q �,ȱT�B�|���mՉ�����7�A�g�:;�=�
�7}!�P��=����Q,�<ITe� �H��l�w�f�����
��k�9�5��BE�O��FB�י[�{�(Nz�P�.O�C"*�0�'�V�GK��^.���Ds�%2�>f��޿+���yb�y^G��F��ޢ6�wlUÙ.{��<��=WZSD��?\fi���InT9,�2�L���.�M:B�ۅV6����P��[J�Q`]"3�ƤqU«2␃�\���7�8ؽ�2���(����n�Ti��i�[t.7]J�#1�q<mX�c�K�WR�Χӷj�Bw*T�m����&� �J�(�2|HFbT���y�T4oZ5p����Ӝ}��Z�z���1U�t�p;y.�oMq$��z��M�zH/҅I|pgG~7���������O�>=��;�ʩ� ��������`�_�Ϥ��f�
�T��^���5S���#�|R�"����9{5{�ǡ/;4m�}��Q�]�@��r����}b}�[X6��Mo����s7e�ع����ﻮ�!�޻���J������<���.d��*�L>��a��A��:�^��F%4�Eg�;���{~	�y}�5y����y�T����:���Gy�5w�;�X����^��YM���t�/�Gm��s3�'���x��`�G�w<;���
B2Ϣ��^]��'��p�*Ϣ��*���x�h���=�:�^ c�W2���<f;�/<�Д��[���6�wfxd=��ne��3�\T����r<��fX
�K��r^�V�"�7�sޝ�Y�|����*�������s۔hY)q�2��,\Tϑ��!���	�5� E�;&�/x_t��ɣ�f�+��t4\�;o����g~�M����ݾ�X�~����]F�a�m���k.�d���Q̀��������d���9@����̙R�ޤ����ӮG6�'�#�.�Ok�M*b]�"l��kI��e�Vt�������*�"�ǩ�����Ͻt��>.��������x~9U0����+�?���)'1~�?fq��ܺ����2=�|��o���Ǹ�:�A���3Ĕ���u�r</.������LDu��>f⺩��ȶ��n[�i�^��=����*#n=�nޙ�.�J�Ȣ���y��@��|�~���]��G)�\M�>��G���)�F��w���9��$_]�[��^.���]_�\9�Q�PGS zCu��~(_-jP�/�ٍ^'���f�D���k[֥�>.wI^�A����п��eI!�⼦��N{�r����lF��U�T�_qfM�Ԏ��?BN�c>>��ӌ���Q�*=�����Ϥ�Hk~�b����7���z�L־�虫�����{��W�܏�����^'�����q�T{��B�rz��0�9�I�fe��վI���~=ؐ�)�ڏi�����]{�����8� 9��ތ�x�Te�g�﫶O�kj����f����[����9�/���\<��v�|����X��E���t�d�R�VD����ޝ�R$G%h��˝�+Nɶ,��7�^7b��a��t6.�Tqk�]ڭ�q��u$�����z�̧H"2�|Έ��r��S��t]I��"�v�9d9�?���8}k���fJ�^k�X[�^�t�:M�?��(F��a��3���6��w��^��~͕��J��u5�1U�{zg��<�O�|)���%Bcه��'���n�;��/�я�tYk�S-l���T��עk�{i���^oy`��p�*��|��̭�갖G��1~�۞8Γ�;��X�3�����0��t��`9��]��{�03ΐ!O����u��7F��.��}���@;�5�0n�cg���z3j󻪷�r��mS7N@J�����J�?exy���Có�u���YR8��c;�npe�����Q%D�f�3�AH��\��a�����I�{��yNz�xvf���A��՝�u����z�v�OOT�~UIncb�ԙ�n�K�^Ң;�<_θ����Iw��B�K��j�}���g��,ӂ*2���_���WO�>�z���R�&�S�p�P�ZZ�����Gv��=�0����W�ه�.K4��ʌ������׽&Pr/s}�sQ=�ϒ�W���C���0ϳ�����&�=냦��~��	gQ� p��;��]�n��/e2�h���U+�k�,��'9�nd��Y��d[L�0$DÎ
V����l�&�Q�'`%�.�AZ;�Ä��u&Ȍ�k�L��R�Y�~˦���ޔ�n�R� �&�4ri�e�;����c����j9�z#�zeт
�����P_n��U{�zt�����z�>ȁ��ɿ{ՠ_�=�W���YW�Si��U`����Q�Oa��"gz���NmC��f�nW�/ޔ����� �T4�9^��5=;�!��>S�g��3)���%�h��~;F�K�|��ƪ�m�Dz��`��^�ӷ�K/U�����SQe�����Zt_���*�6��yp�ޑ�6�yj��=�Z��^HǛq^�q�� ��]�*8f���L5ckC��i�q�Iەr����kJ�-����isX=��U`�,�~�ޜ�g��.=�۝9�q�ݸ3UsL>�g�{��+����x�ׯ��P;q����u^�������G�eneH��Iݺ�D̹�{!go����>+�qYU����*��LQ��"�U�~!��-��?R#�mG����W�8��k;ݷ~Ry܀�����S<r(�`p:-Hʓ3��+D���Ʀ}Q7��ޔ�0�����^��`���$��\??�Pz�i~�WM�Nm�׋�>��'�xgOt�P���|�h9���eJ�l5Bg�*�h%wԶ
�Z�m`^�OPt���QvCx�I�R�e���ŗu}�X�)N+�PU�&�g�����J��f��1[b�u��Ց���712��܋���d����u��tuPt3g&��8�t5�R�-��h�)��G��{��b6��,���z�2��|�R���'-�Q����;}G=~Z��	�$�������=p��=���=�.K4�UA��
D��8������A�I%x�O�UAW^xċ�[���^��+~��=q�Bt�{��d��L���V��w������lz&�<�
;>��g��4u�TJ���!�^W��~�M�Dm��b�+L֓Nϫ�&{Wr-�F���C!9�r|}��*5�Q�����Ӝ}��ZZ<J]o��;i#?����Ulչ�X�U'��D�/�!WR����/���Q��j�G���x���Ɏ�'1�f�mw��Gǧ|Jχ� ��.O���f�
�W��h\EzV���O�W��a�3��rd����+�.Wtb�~�G�>��_Q�]�@�W.OE}�}�+�koG��xM
��,�(W�z%kJ�؍{������xd7�}!ԯ�ޟ z��+O���x��P2a���.m���y��Ժ]3謥������
;om�N����P��U�=8��b��nF��ۥ�<�SB��j̩[��B�6�T�D��C��AK����� 
�1���Z/�{"B�Np[��H��W��w*b32V!�[R<�C[&<ӥe�T��o��[�RS3���e�3��v���Z���[���:� �Y�p��d^�su�
���	�F�W�Ե���t윊3C��[ �丹�7���;��R��\[3-��a���96c��1�َ��7�9��t��]���6WR5��̏S��eʓ��6c��R�ƈ������A�P�!�mh��Lܬ�ب7��e,g%�и�MB�9��oqkR4;N��9
6@B���W%'�OV<��ȥ1��6x��ֺ�^>p��JX�Vc��ZI�Q��)��¥K���f�X���"{<�Cs���-�#+joF2�ՙQ��EveG�x�_s�y�+oe��(��E}�`�AM.*��ɚ�Q��dWB�c{j�JB�h���x���ɶT��X����qH��w�)�Ryr���I/�vCWu��Ɔ�V,�=�(��ɝ�#xT1��4�����+6�Ӏ̦;j��}sC[ujM�M/��V���9�����v��A�F�H��-��}�eȩ�s�j�s��eE{����XL�X�}/8�����c)�s\=)���
9����ga|���)U��DW���q�ʗ*�^tL�e$?e��0��&n�=�7i\яu+]�[��PcU��-SIo-\T5��J�:(���eT�=�f}q�b��2�Ħ���b�:O
Ý�}[DO�m��1�x4Xgb�E���_�j�Ty�OVq4�=Gz�+d�����Q�Uk��l�A�άP��a�z&%<��D�i3��u#���Wu�����&�9ARQ������RL�$��ݸ����CZ��]�)սv��9F�L���d8�����*�%��V�n���� /gB�G�P� ELљ+������y�wRǕ���|�KY(ኝ��I�n�gn-y����Ǻi{o�!�`�*諦�y�M�E��<��Sf�
9�*�������Lސ����ؠ�̬s�%�	R*�]��1�tݻ{ו��Ch�z4U�����wg�)ˋw�oV����W]���m�F�}��vM��;M'rI��v-T�������%!��o-죿@��V1c��y\�R��M[�3��]ݹӣ�A֪&`�^���>.��n 0ZJf+V�c�h�v}�f_ZV�u����yQJ�|���1�W}gX(q� �e����+b��S�E�z)�J���qR$�T�"GH��s�c6C{ʹ5l=Ø\��+�'������g��y�.�l�
����iZ\�2��݈
TQ�1���oM�u]�Xg,�ҹ%�\1��d�@*�$Y������9R��;]J�G�䛘��+��2>x�)HV�����논Kȉ�������E�t��JN�v-������v>��jQD�ڴP���u�,�u b����9�w���^n^��%�%̍WL��\�ˤ���!�N����֔q-�{���+��-�t����뜼�*tB��iNB����#�Nm�9]<Q�Z�yr�$��HB5ܽ��r�`yH�n�W�yG���:!U�23�2C��:��J#���=\�s�E��X94����E�d�9��s����ȷpJ'v�']�W/E�2s��c�z#��UE��B��-ՑfNI:����vQ8�D从�"I�Q��.�S�����<'wO.F�t3b��� ����u:K���O$�Zr��%�V�(���:�#� ��wid�D]0"MB�f�^�N�t"�E�e��ʥ�s�Y����wO,�B�DJE)���D衖IUQ&Q�D�T����(�$�,��G)Q�Õ9YA�\�R�P�hWCR��$��P�s�s2�Ĺr��r4�X�DG���T8uZj� Q |P��P�mGO+GiY���TіIN'%�3d{��%�,�f�3s��WE�gݦ��ծ:����]*g7S�c-��<[X�������f���u�SF�(�I�q�_��ڿ3>�yz��w���,^y��,ؾ�s��+F�g��>��;�t;e�:EeW���(�.���=��ix��b2Vz��
.=�;|7��ґ��/��	g߽{��9�A>���m/�릿3����%��Hb�r|	ˀo;y��{�_��;��������~�f/����8JVe��x�qS>E��4Ey��6/�4���ğ4g��3A{#K�/�q�cs�����]!��sX�5s,�Y�OQ�~#��)���x����X�L��������wB�:�^�>gs��P���iP�)�.K3�Z����`��>�C�Oz?څtg����HO�7����ND/H��HJ��5u�Rr/�[T��=cub�	��d� S�I`Hn�P��V}��G"�����֑ȃ����X��ɟmŹ��_���#o�ulչ�Y�qU2���p�g�KGZ�6+̧Pl�(�z����{�]��Lzb�2<s	��\�]ߍs%��RCW@0��L/���C�s`����vTJ^���t\�T�*+{��nh�ά)��׵.dû9X��u�NW�T��r��K/r�eͨ��V�v߻eqj�q�����3z��M�/nVr�A�������+E�}���3m�.Bo9Uv��Z�i䏛��a�w�u;Km"�D�w%�3�+�jFs�a �Qg�N2_����{=q,I�S$5p'���Jkʇy��P���)��������j��T�G���\B������w{��|��C=��9�Q5�5��N����Z�_�x��>gj�n�^��Ͻ�WF��W�_���憫�J�=��o=S�{��:;֏y�{(��Q�׵>�aQ'�{����;o.|����ޠ=E�;��}�fց�o��to���Ŀ}�t=�je�GO�F�O��:��d���f���p��?8���\�t�rWk]=�zqK�#}U�=������~��9�?�����·T�J�.������h���Ipl.O!uO�!ׯ�O�C�G��1�̩��Γ�;��X݇�U�QXWt�vg4۫۞�>� o�4���-W������x�T��y�i�=�G>�����s��;����z�=G�]FϦYا y\F���4����o��<�hxv:�C^��ͧ��&&���^�������#}r�,�I~5UG��3�n�����T�����i>+=�yL�(*�#�^�+����k��ĥZ:]���`R0�H�����t��E�o��F�I���r��jkYt&�������N��h>�ܴ� ���#���{��`�Lq��r�w�z��ҘNI���8I}g�{/j�k�u���r�G�1�պ:���2�~�p�S����`L*�T�sS�L�sBz!�q�|�Ω�3����xQ�>��<z��3~>P��|��ʠ�B����WOƥ���8��ٻ�W�$�o�'���hO=O��H���\���0��f�P@��[ gj��(�t�^���*�{��r��R��z�Т'�v�g[��]��Pp�}�\U�2Y@@jL,zI�y�.��];��ˣ�P�u�n"�e�|Cw�d��~v�z�>���ɿ{ՠ\z��W�B~v^;�j���2dV��G۳>�$�6\�}��9E�ڸ���|٨���~�q�����z� �>et�0�O6}Mp��wh�9�/�3>D#c"%�h���~;F�t�<���~��k��I����.{�W����(s#7ʎP�SQe������D��
�i�&�g��{`8������E��v�gϽ�7�� ��H͈�l��5�6�;��i�J���<oۑ��A�����%�Ύܪ�Ǔ�,����ӟ}����/�{v�NDq�;����[�Y�Cn�̆:(o�ntf�k���4hU,A�؆���n�ΠU���]�zp���8�VY�}|�E�U���5��ɼo(&�:�ǃL�g��������H���%�F7�z��l�NAU��6���"�dR���8g6e�G��I�ٞ^;���N�����sʼ:�_����k�C����ߚZm~�Ҝ?�꽵�jYg�r�Nߠ�v�0��ʭ7}�U� ��Ցj�O�c��]8�����J������}"�����������p��C��6(�F�ٟ@W��@RN���v{��A�к=2^
l�}��Z��.y�n���b��#�qcK��A(<��ʷ��;��g��-�u<��g�t����[�ԍ��΢������z�G�D9�E�fY�$�,	�|�*�ޏ\�V���O�b�6�G}�s]�B}��߇��z���Pg���{��g�{�f�g�*��2���3��~�ݔ��='Y��U_Ԗ1"�[��ȅ�2�;�4���'Mǽ~��Q>&'2�}ס<���VK�4�r�>3 5 \>�U��4o_���O�� �|��N�'ў�������y�5�Z�%���W�L�5���h��%��n|}�T4n5�Q���#���K��{�#�꜑S��{ڸ/X/U`��_�2IcaT���I�HT��lq��kF��:3�/�i�N�����e��^��s���a�pw�)�+�b����y- j�pcP���Ȩ��MY�c�eιn�ڰ�n��@��:�PVbŊ��
�f�eg ���i��1�A"M�ZTbg7$μ:(t�f�4YR�TÖ��Y�M˫؅��1������sh;�����u}�>d��}9�}l�<�I�3\X*\����+Mv0t��@�c�B��k��y#�ʤ;��wF���Q�O�O�Cβ�O�Y��#)��пa��.��������&v:���/�#Č��9]�a�UPP��Mǽ> ���V���Rt���MV��oGH��[��qy#��:�7G�}��u������N���>���XsӐ��b�^���S����&g������H�9D���pwj=u��n(�'MƩ~7�j�2U{��^��^ٳU\c£6�I�-Emk�����NI���(��z�x�2$�C�1�
~_z�=�e��N�����[Ӿ� yR��[���%�w�ߺwfxc�:v��c(L�W�O��G��]o���yUu ��y*�3�qW7O����u���W�Ռs۔r����2���G��
]�5���sv��X�����B]}l�=,b~�x���t��!�b1meK7x�9���1�c��=��A����[�-���T��E��G�x/p�3���_��Ǹ�:�A�0:�����5J	����A�s�)�o"�J�{�����$�F����z����x�����m�'�8���`�;�X�aq	w��䂉���^M��b(�ݬ�F�-ԕ{:���fu�����\vRz��>3���.L��n�%��W���P�P4����ad�z ja�Q���]T��巷r��N/H���P��˨�w�j<�M�s���j�~!��z��� �>�r �$0/���l��V9�?+���z�5q[g˽�6�n�D��o-�n�a�R4��{�F���f��,�(#������B�������;9���&o��Fo�?Jv��>ζ���'��pv��w�B��f�T��.8�)�fsu@���{��jVo���Q�����\���W��A����l��j2D{�뉸f}&��t{�bzr�`�ڻ��mn�WG���Nem����\j�\sw#�����^u�}���7��Q��[}]j�n���}U�&�	խ��l��29/*�w�G�;W����_�{ή���P��z�%>����n�<��jG�?}�r}
Y*��pvp9������}�/��m����v�G{3y��=6:{�K;�`]Bw^��]
�972�>��(��cgC��ڗ��͕�~��^>����S\9GD�6�Zz7�*��1�'�������hm~�=�b��ZO�̴U��![�"��EFr������2n̩�I�a���Qǝ��=N��;�j��ʝ�5���gg+F��l�G"�'�����p+)Xj��օ��-J_�X8)BT�·��컘�WS�b�:�9�s���.�+��!�Z[�w���q&�o}g�R�{ś�}mn��zS��F����xƮ<�~�}Z�/���YW�ǻ2��C:N���y���Ǟ]\���'�׏=�xz�k�Ґ��L
������]{�dz�����ǹ��>�ؿ����]#N n1�}�J=�������>�w�z��Hh��-��>�χ���������(Q��ݛ{K<�/1�YR�\�'�D�x����{��&ṵ�z}g�{����^�k���gq���C�6��;�C���Z�]|�'�e�#ʡ�L�1qS�L�[ub\��\L6̊�g���֗k�+}�}���:�3����ߏ�@65��`)@���Ѻ���.��s;�qI�-H�﫺���}�CFB���;ޑ������z�x.K5�*2�؟��^�s�O��]:�^W3��|KjT3���h�O��>ζ;~~��n3޸:o�]��%�@�f/ٰ��w���?k��]��7r�}N��|^�P��Y#E�~v�z�>ȁ�����8�`Ӗ!o���>C�z'ߜ�71�=��&���J�<�&�j��f��U�)�ԁ�^��z�ff��}���DN�������!�����P-��4U�d�~k�x7�T�^h�!$o���e	;E��Ͷf^�r���\+���L���-���NҔ��.u��Ġ8ŭs�E؈����b�0gz��3wl'qt�u���C"c�]ߟ�
��7��3�o�}/�E]K��6�_�^ۏJ����lɸɢ�S�^�>�>dѿ{�z���#�Ӳ�X����JӢ�)�xUV	�eOZ��A�7������/z��=�K����~���Gپ>%PɆ�և8z��|�-t9��Kߏ��/�#��Y��[�x'>����>�Mx���_���s���̪p�4e0��eo���D����E_��a\VR�qJt�V���~gՠ��yz^�U��yu �=���u�9�*�߷�������3|Z�w�Zn��+D��&���^��1�F����6fj��e����ۏ�����ߣ��и�:�=�u�'� uW:_�.��_���P롾`_���/Գ��I��'��d�����ϕF����S�x]��z��C�&x;��|�."���{O�a>����5�g=U m�iȇ����[��g�k�Vf賈��,"��do��G�;�t����V߸z*��ND_�X�~������}A���q��sY��%��x�)�;�o�ç�N���N��)JF�����YRV�K\sQ1V]vvVt�)�O"�����渺��Z��z�fe��M�95�F5�[5D�ڏj�E`�a�e;
���˚��7F�R�=��*�`��\�͔U0Rw���9�r�sy7��b$�_t��^`@�$x�|��uT]%�.%�^���2��CO\{i	��W�=������r�v�J2}D�3�1z���J�U�T4o_���O����#�ӣI�|��������%�Y����<CUT�y̕4���G��n��_fPѽh�m��l�c�����|%����~tm���z��U�չ�X�RZ�=$LD�Ru/���_�˥�N������}���.r���~�"|p�s������H���(�k~
�TD��Í};wl��g/Ņ��*�>Nq�!����1���#����f�ǽ>����"��,�_+�'�\��G��5�ͫz�ѿn�>�M��D�m��R����Lu���7���Pu7�O�=�q8|�̃�)��vk�	��5^�{�����s�TQz}��lp�:��8��<j��U�=;��y�kI�{g263��ޙ^���r7!K'j�Ѹ;�Ⲽ��zN�E���W��g�M0�ؗؽU��{5G,J��f}Ϊ�=����rNj�N�g �t;���tW�F�ˁ�|�=�|1צg���W�վn��}��<��Z��=�=YB�2�$�y=��(,����7Y6p���].�[�L5�cV�Cg���$z���Е�4�����k�`Z[�$�J��*�*_r���j��sWC����C��2ޘ:S��-w+b�(l��FvV�f@9|�+>��1׫�[���%�w��{�vg��p����Y�O���k)�*Y�w��{������K��o���޺���Z�����b��nQȋ8JWX�^@N�S��[�}Uޟe���Ӑ��dyv�lp�z�܇����]!�fm�k*Ỷ*�լ?]{�Q�$�A��k�;H_�2����ϭ�W���3�p�3����������C����5�g�JX��6(�>�x��Á?*�qFX��t������M�w�9�<�n��yY��|1j�ܵ``c>�*#o�z��� �.��9MD���Kee����~W�i �M?8]�v�w݇�vs���/H���Yu�f��,��ِ=!��l�nn�~ة����� |��;����Sf�u�v�t�~��ۊ�ߌ��̖k�RCW��<fk��߳݇�ۚ����=j�g|��3�>��<m�׍F@����3>�ۊנ�!!���5�X��<��`��Qߨ��W����T���㚦K�偷����1���6cm������1���co����cm��l���c`�6��6��m�������cm���1���l�����m�ll���1�co���6cm���1��� �o�q� �1�������d�Md�˜�
��f�A@��̟\� �ԅ*�*$���$(�RR%IR�JUT�JJ��T*��J��J$*)UJ�EA))A*T�R%(�Q�Q%��*�նT()D�$*(E *�bR��%J
")UQUU*��H�T�`J(J��R����Q$������QJ��*��]`���IJHH��T*
�% AE^������D)"���Q$UR��B�A�J#�  �r��Q�L( �KB��#Z��W����CYAAH�jR�A�mlMT 6SEJ�0)�  *�JK�BU.�  ;�B��kVhU�0 Q4XptQ�P���tQE (u.: ( F:�� E q���(��( � QE�tQ@P  �UT%v2��{T$"<  k� Q�nu�Cd�;�UF�V�PFij٪�j��(QT�R�V�Et��UkTl�� ���Mj�T"� Im�O  7����P�����iU�6A�4�ij�SC^�C�j��4��ԭTҝ qm5ZR�� [�SP��
4�T�J��J���T"D%�  �N,%���`�jk1` Q[he�U� �5��ݵC��:���[D��ڀ`�I�j��4uGT@u�YJ�һ��T:iR�*��	Tx  �������-I� R�,նh�WE��Ӫm:@�sUZ��l֩�Xi��PnU��4�ڗ%�45���[`	��m*B���U�J���   ��Үڍ�p���Ѣ��)�Tk�G[��ն�j�V��4Z�6;`��X�n�h�S��*̩Z�	��T���IE%$))S�o    �y��QA�,���qɀ�6iQ�� j�1L[i�m�i��
Y���m��Jé�@��+R�����JЫ:��#Z�R��(�l�o   �Q�=h.F�SU��h:hkZmӔ(t(��F�뛄� R��ʛl)��LMR��T��kCZuݵ4��R�*T*��d2���  n֚V����V��S�s��:*�u�r�-��k���ں+iU��
�ZjeV���@�4�iV�E��]�+�T�Xm�CMW���&eRR�@ �{FR��z� 14�i���`"��	R�`  "��zUT�L��i*c
�T 4h�O���?����b����eb�^9����ts�ٟ�k�����~���������$���$ I2B		���$��	!I� IFB		o���������zx����@,��t���n7�2�9�<74���wx�יQ�0��X��������#����5��c�T�捶"Yb�^H0+��!�Y2<���1�dc�ݤ�A���r�ج3JZԭ�j�[��L��IX�gS��"�*�R4J2!���ߔ�D`���2�c�ѦMMЊVM�����7[LmQ����7�R�l�R�����l�J�Ѧ)5U�^�82E�j���O��i�4�I� �]y�cr\�W53yӘ�I��A�YU���-;J5��]��`ٻV�, L+բ	1䩣r�-GZ�3k"擁��Z*惎d�F���/䩇�bӵ�՝B�I�� ��a*]�M5S	�l���q��zSj�v�L��eA��J)Rm0j��ݨ�Ah[��4�U:�˗]� I�[��{+6�(k"K�6%
��Z�]��mmf�7G�M��R�3W�/h��f��sJɕ���=�ՒYS�&;(���+V���͌ص�Z�7Y��3`nR�C�s�m��Е`�؍���n���6�wx�B��t&�{��{�͸,�`�ۈ�)S��j��N��lb���̠Γ�\'���S�����U��	�y������N������/�51H���e�YX��j�Bf;J,���R�j��e�ZA�/L��;���d�S�&�Ut�Qͳ%���"�/#W��e߂wN2f���uuv��M���搆�+@�՗�6���^ͨ�cPa�~�M��Wa*�\�0�V]����ȱ\Z��#��Y�$����h`%-5i�r�n�{�*)���9t!��of6���(D$+]G{�;ɭ�:I"�p7#��)0��n7lJ,8W�F��يL�f�Ad��[R<od���D,�,��ڏd�,=5��u��/6�귍��Tv^M�n�#u�s���"�J��f��� ɏTK(��H�U``Le�j���b�x�j��f�+mm�W���e&c츗�aLXn�-&�݆��kC-��͊�E���1� ��8�^䊮����j�J���̆���ǁ^�I��W7!�@e�Ys(Եt�n*ݭq���	��t�B#�2�r���@� �3��b+.u�k�b��-��;�6�4L�V�$��k�D�31K�ӆɌ�X�W`�-�BQ��K[sTs!��6��yk~�xV�#̕�%�9��4͕"�V+�=��{�t�l�IATyv]7�-�%�z+v�M4Իѻ���P͐M06_� 쫅��u��**�q�F�.#��o�
�u��k���7`D.�M+H~�Z�/-=7���$�Z8�Bj�� b�*<�fƼd8���Gqۆ��ڧy6S���� �t���u���-Z�q�����mbR�5����*%���*�̈��2L����f���iv)q�x'��F��uaSǩ"˕��U�6,�3/�Bmh-�Z)��N�u��l�ef&5�cvŨ��I�n��ע�`��Pѕ�dɢ�c6�;�4�D�`ƅ1}�i���^%W��lq��*P)21�̛K,肖�i6�U�uw���kl���r�
�Dh��pe`�wV�ZT�b��X�QŁ�����bo	Q,aޡrv��Z)�$�cG]�[��H4�� �^eBCT��fm�g�%n��7�,��!�Ä[)�d1���ڀL��IIJYld��3tj�A���r	���swC� :髳*bb����KZt��YH�t��T���s+sQ¤���Yz�B��[6�غ��հ -�5`U��2��4���!j:�J�n��i5��t�d�{V�왘b��1}�E9$iD�	Z%1�7!� �W�r���e����S��2�8���m�fXSJ�۱�S��$l��r0VZ�eMDÕ�eT�[wsV�e!�9�2��o3)�Z6[ܨ�Q[�� �u-���"LJ!��f3n�H��d�(��	�Ĝg3M�[M�C���қX2�nK.3y�dَ��f7n�QH�8��^8β�?^�9(�E��j�U��:GmPV�m|.�Al��a�0\�$�yv���L)mÔ^�LX�م$dn��v&�m��LْmG��N�-���D����cIC�&2U��-�G��Pmfꛆ�2�9��p�:�d�.P�o5��L����dR�x�BS��%\�E����V2��LG�ws� �ᅰk0�aV�k`������F���4��J�����(�#��X�f`��oc�W��0GCma�r˚�;����nj�xk0H�ȷo��eLM��$���X����B�EF���,	��U���Y�V�Z86���f��B[�V�F;okU��:��@�%��&�&Bz1#��VK4�jm����04��1��[�ӁD$0X���0�����g��Gqڧx��f刵\�� �li���U�Tt��7PV�m���c��AF �살hV6�{�ꢴn�N��s��!����?fR�D�{�Kumbw[
�����]c.Fب�P��7Iȳ�.���"�l)�+��jYʽl%>��Bcʘ\W+v�^ȕ����R�-g25ǇKf'D9��W�KU���@��76��ȕ�8�XlR��.5M�50F�(�,��.�"��������Ь�/M�ǅ;Ӗs^��Ƈ�@9�m�nY�{��n����Ö�5;ZE��I���-����
7H��3�!�Kj��u��.]�cIb�۩sR�n��O%]7n��V�*)h[�5��_L fV�95���piaˏ6��0�@��n�C�)^=a;`��[6����)=�f#�:�S��n]�TA�/l�eedaܡN�n���Q0;��\z]h����7�1I,)n�\�w��7/�����;��B��Y��H�6IYcz�`ڦ�iנ1J�4�w�#���Tf����{�Zb14��S,@D�t-�P<�D�k[���i��W�mm��%��≐0l	��]^a�j���0%�V�n�'=9V��af�q�W-��3�v��ɀXMp	���{��p�(�w��c`�J�n�[W�+h�V�0BZsP73ZxCA1$�ջ`�u3[&�a�8V�j^m�H��Q+Z�$�<i��,&d���ѫ#�Fֺ�M�a��i�m,����f#�^�����/Su��n�1�iA2V���v�PV�5��):�(^
_n��Z+-փm�h
�f��ͽ
;*�c�����]�v�30��%z�%n�K��9�9q�@	x��j�:�ɢ�4��A
P譲S� ����)a� +��vW�DT��0�;50�wNۉ�3T��~x]M��k#�XJt&�,d�v�boz��b�5��iH'P6�f&�4�	1�"�Z9j��!W�g�iV�P$Ѭv)@�Lf��nK3v:�2M�j��
n�A 3N�bZaS3�#�qn �M�����ս��[�HB@Ś��<̚���R���a��2�b�U�JƯYy�����LLZr��m@�hg�ɳXHvH���f�{J�˧�[F���S
MN�{0�{j��ެo!��ηJ��h;V���Z�w(�VX:��$/B ��d;b�$��AGr����Cͣ&���{�DEe���Uk��)�&�0�pֵN)2`���tȫn3����Sh�f��!��rH��a 6�D���[1��ͽ{���S	�2��j�+,.ͼ�Aw�P�5�;�xdf�%����L!f�C�����B�@�AkF�Q#+õ����̫��a�[�7dM�����j��Ե�`�j��w�e
�Գ6�Y=uN�f�",Vk��7���a#�Yz�R��N-�m@q��
Ë$�ش�7���Xj0�e"ɖ��������4Q�V��]�Nn�ɸ2�'
.a��
ɢ�,R(��.��6j �F�*���Y`ȣF�!6L��-cN���Ӵ�n�Dɮܬ�1�4����DR�q'f�iG��Mnn���r���\�ax+N��fn�v�D��u�2�1e������^m%Pkxj#�Z��,��R�u5��zC��q�
��t~j��X���<�f���8��֋���"(mU��k)�K�6�����մ�c�t��:�gi��}��Y�t&R&[�j�n�(\4,��3�=���-]ՕcuQ�i�.�N�O�.�s	��>�����f��*��VmZ��P�{M��J�Yz޸]`�!Z����h��R�s��;�j�4���+�����j�ٖn����b�V�>���S�ǗWp�iG�0�Q����t����hBV�����Q�@�ǪASEL3e�Z�۩��V���M�憩�Z63pU�VĴ^̢�lz�FV�O�%X�y�j��#H�e�#-9���Km���˱��r�Cr=��iiXt��L�iV+EVR�84S��5��;� �b�B�ˢ*�$-�@ʊml�:��a��^dF�@��Z�5,�DH�l����!+K+U��8|�>X �g[�r��AV�n�^���֭/���ơ���2�rK�
���ii6��+����u��Y�Q�5����qn�-�˴��.�em�i�M��@�n�2�U��ƚ8e�m��f��2f��J��J.U��br�o9���q��6����QcB���Z��^Wq�P�� �b�W(OP����M����fG�&u.�hf�3v�7M��.�\!�8�s[�c-�Ԏ�v��B�}�A���9��dZl�������PR=D�
�Y��m9���Ԧ*,-5z�3B�K6���r�R��kQ�˺V����^Bl!�^�q���ΒK˳W��#-�h�wp�u���tl���[6�P����Pe����J܉�Wf3�M�b�I�����:������94ò�:/�D���b��6+9+n:[�ƕa�X���Zp�WA:Tr�!Y(J���f���֎X�5���cP��,��[�kf^+��t`_6��ˀ��PL&D����w�Ҷ���5����F��ER}��ihsF6(*"mTa���mƯ6���}��;@�il��KM��"#�I�$�{[�m�8^�r�5oig^�@Kȕ��� l��I�>�����T�f��N^
�+.=�a��^J�6\�#��h(,YY�
{�A�#6�<B� 0�5S����F%�ɹ.]صo@GH�L�(�Pӛf\!��܍��DU��&�S�j
ꬻ�����T����(d��#��'/J6}�>n�E��a`H����SIK9�)y����^�"[f�oKB��hc�q'���[{���rA�)�A���d˰��hB�Ï&=��Vu�{���Oi�<N*,@�J�m˟S��`�mрP��)9�.˷v�:;�(�R!F�Lц[�0��9µh�yR�9�5^���	%��L3�e������}���ʼi�LC�Z[n��7%�6e�ሀ"��U�5�M�/QEl.�P����$��v�V�oj�
*yz�X�e�@�cieb��k&\�R"��� t/AI�RQ2S���0���"
��X��wC8��ƪլ�M�m�㻦ǵ�����T�`y�JX��%���ʻQd��[MPS�%h��1�bfR7i�'eh�U�rTWf�����u	GO�G,F�gע�Ig�l;.��ZN(����eL�S)n�C3�H��2�YD䩌}-f���[����Yσ%2轇U!l�B�b�4 p��r]��Rb˗B��,�(��J;��m�]"�B݄ͻW>�	i+�dEt#T��j�	
2��n���7Wv#�Dِl�U0��+�d۵L��O.�Mܰ���wgY�*�z�2��v��$4c���;�f�Y�P��g+u,`����j�M[*��ET��-Aw�h�n����J������b�[d�ˈm�چ$��5L�ZA�JX�Փ-V�q��Z���4�N���X��$R�4w>��	���t�ݼ�� m)Z,�cf��2�p��+Z�j5,���Q!�6$-�������Ԋ�K�WW.�rJj�*{7[[06�b�J�Z�d��e�+���ۛo���z��VIְ�*����ov7�u��5Xo%��̶���.���y2:�M��,���5cKI�ke֌nX U��A�t��4�JB�1���v]Eu�MQM�ӘV�b�b��ʎm�ɏR�U�u�@$�V6���Iv�$*��_�2�,*��tЖ�nd���G Yw��+2����@M�fixU*;0�
��0�С���)e��V7(�:���n���r�dʻ˵5kv��*ú���y�(�+2Ԣ���y0�"̈�w>8�&����VidWi����,�÷�Lo �nr�ۧ��*]05Su+�7d9��vm��e�{�ot9�ykn(��2��C	��z��gm:��������ӥO^�j���n�
����V�-$�c6�䥕w�I.d}��-�(2�<>�NPϋ�[R3�3�8���E���*b��&f��e�� ���[�	��] r�r���JO$���]���Ñ+r����!{y2rT[�������Mvwz˻��+r�">чE�-T��Y"��Xi͛,���5�u��ڦ�
J�5�qK��d�:�r��pUָ�PLb8͉�&��!,6o[��Ҧ@7�f��&�iZ�7�* �67�'ّ^�W.�m\�v���W>�F��:voU��Dku�w�R\��|�L��s�.�y ]�MT��O��j	j����_.,�e�x;���Γ�,���D2.I���;6e:|�+	p��$mK'^��O���M�P��Z���
��&�[K��U;�;o=�w��3LN�1��8澚�Y�V�\4�v�s
�jv���w��GG:�+}�둾{ki�*n���u��+�rح;�շD��5�aW�4�!}�w5NƤ�ouX<L��͐�^�3�t��B��uό����L&���Bh1�g\霊"���]���K�9V���LN�r/���q���ě�coH�uk{J��a�ќ+���d8����}�����t��B��))�ҷG)ӱY¥��9F�k�+Sgu�s�y;�F�p*��[�>�reϱra�[�-����%�=��\��&T���(�Jy�澨�����p��[V6�7s3�("�:naU�K7}A����|�)���;�L�c/���;�J�y�������d2��RLK\��j����WI��ɺ�KnvѼ!Z�C��n�1@n`+��ڭ��������Z٠����H��z�èxŏ���q7$�g���p遶U�I�����1������N��LHVr��H�guZ��ӄ�C�$me�XD�^ ���U��n���ZXK�m��Q��/��{/2�j[]�jSU#f�|�*�j���k���B	0*v� �O_Kw�	7�p5u9l���=*a��=p���s�!!0��@�{l�JvO7������i�X�]�V�ІO�E�ϖ�G���p|����ڝz�N�*�_ê�.�.�^$#�z���vKFC4��g�7�e$��z�r�Hu����J�g^YR#N^�"���K[͑�6���;�u"�$�.9�IY���]+kѩ:���-A�{Z�,C�*U��̭�F���8b���KĻ\��c<��ִ�n�ٴ ���B0�̬F[q��'N��Z��Rwi�KZj��7�ݭ����u�Rї�t힖-�c}}���BygpF<�^n���o^��/V[ͽ��L1��Sje��N��w�p��&��ڶ>9��[Ϻ�Y5{ʋ�qm!�P\�;�׽�ȑ1�wU�-�l���Ȯ���ʲT�[Ŭo/5��յ�9�Ŷ��$�IRf��l�v4��wgu�؄ j�{����������aʕg�X$�'�����8`��ȫv>�/�����|�-�T6#|���T��7�@�����7�ܠ��/�6���6��x���G��3N,�յ;*�j��aUs9\o{$�\s�-�GQ����9�rl.�}�s�/����t�nr^CpA��`^���u��B[治o�qrwCu�*[͐���_Vh��,ֈ���ںI�$��䷷�����v��G���o$ev˾����ù�ٱ��\Z���fk��D�������O쇂����d����Rw8ܙ. �:}�:��Ub^j��Ĭ�;� �1�I�]�g�f[�ې:zrÀ�dG�Uյ� �Hk��_.ݻ{:�u,�*Z%rȻ�R�:[�9(b�]P��v�PCb��e�짙!;&�<�e:"��ؕ�i�B�a&�����xV�r�bgaW)Ygb����#�;�;�ܠ�{����ʎ��C��{A�B9׃��>�i���0�Oi�'`��烝_	�$�NWdf��qt<�������!5��P9��X5�tv�����r����Ү^�`�V���X��^�,�V�D(��JG7�T�d��S��Ƭ�m*F���l��)�7�5�s��[$�Yw��=�@��:�KmI������5G�yYX�����u��J�I4��ᖭu��8u���������F���oV�k1��op��IX��ӤIܶ=W�h{V���͞��\��8�����T_f�i���{b�5y�;���ol����كST��V;#���E�'\�v�&.��,옷+;6�ok��=)\Ut�4[�͠��b�2�}��-@_h�!��T�>|6>���fW��:+�{r.ڕpS���ohn��6�$6;Q���n(+��u��Wұ:ʐ�D�zu�ۑݞ� ���w7C�&+7��͝u���7/�L�J|�3J���sWw���b�����Y���t�X�y��%�̃�՞
�j;z���BxM�I\mU˝J����Y�B�(nU�%N�;8�$��z�v�]SS$�� �[�"�@����*�z�5!z�] �;��̤��ojs�b��R�,W�\��ȴH�(��Mh�G	c�i�]#��a�M��W`�@�R����[�C��n�t����z:.���ֶ�������w�pc94��J�z�&e��UἩ:K�
*2��Ŝ���8�*6��q��ĹK*��u{)��ۼ�$��U�<��Jq�"�:�0`&B�	t[:�6o�t� �%�&r�(ҫ���5���4�X3XW�ET0� ]�Hgee!6��Z���iX�?P}�{_R��Vبt�����iV���T>V��|��.�c��Ѽ-�W�[�I�.K����q�X�n��)]u\���I�a��-�H�]G%������0J"��/�O�����@IvE��ڑ�v�����γ�v=�\�������\��;w����(��r�g_f1��s�f^�2��q�ss��Gu g�c�Ն�ܺoAc�f��[��+�6���1)v�ECn��iX̬YǘgG(��
��b�/e3M5��9G۪V�O%c�i9ըr+��vh���j���p���jf�&�v��P:Ϥ�4��5g
��,ՎFs�݅���x�{=�˷�C�/aB����M^Mi�,��O3q�EI�)j�t9�N�i���0�I��%�(�&�a&� ǲ��tc�Rg2�F�<�S�/7�[���v��F��]`�P�b�~����p�5���o�y�5\u������pF��`�ML�oY���h�W6���A�V�:���Bj��v�f�9�ޅܲ�7�I�b�K��4������y�w!����T�ޞ��r�J��;[��S�U��p[�d�&J���ܺ�\�u1���r�������	=�s�q%�M�DgE���.��ȳb��=�Ι�(�k�:"^���N��Q�s}n��3$}�y���c�����7r��4ENg�!�cT`��cc�cY[}��� .����mC��a�]�(7�,��tqn���D2�;�@W�ta��&:��*8���3��oZ�c���L��r,[����cJ��du��je�|�K\x��+z�����]��r�|�脹�����@�I����- vl�齹�Kf���뷛^J7�����;�wp�Xᩝ&��OyyH��󱂰�|����&nZ���n���b��s;:����A���K�,�B��V�A�K��ǻ�hMs+34���u�-z˦�v6��mnB+���
ykN���� R3��L��Bp�2V�	dW8���t't��yS�;j�� b:(w6�n�v�&&��v������g'��A�F�圭]i��]�⋫iH3:Mq�1����o�̽¦ړ����+)���K�����Xx�E��;�a!��Jt�Z�Ћ�v	yή¤�ݾᔸb�c{�o����S�����fK Y��OOb��,��nm�%��s�a=��Ȫ��X��8a01 �������]-Z��A���>������7%Ym�-"kga7�	�y�����oPN���k��>F�l�KiY�*E,k��|t����I]vXo	�>�P��L<��WG�>y�s�FY�wظ�-�-�u�h����.j��Z��o4:����gz�V�j07�qh��l��i�.���]���Е�>�Z�|��3A�.���J�q��xN&�R�kC����1��F�g����? Mx�{~z	"nKSe��
�]qH�J�tNV�j�u2,߀�Dw�6�D��K�	�9�yq��[γ��@��<PFt�3Vu���*��t�_F�˲��yW���骸���WV-�v��5tR
(/8��]o,�EA�j��f�U������]��c��5G���,���Ԏ��z iKѫ��ehcf�t�9�t;^�0�c�*�V���9Ӝb�7˕#��
Z>�[y���9���e���9�H���%�Đ�����*n�����F f(F�S�b�X�QnS�E9�UΜP�Z�9�x�;��LȒ�f��{jC�7c�Y�P8@Ybkccջl�M�V6�*e<��J�9�֩8U������	�G*0yUmiF�_Q�7-4�]X��Mh��7F��l.�SdI�馸Zw���4cGWc���5�!�ugY
!+.�#����+w1�g�%ݭ��q���zOWS�	º�Wf��\�|����4t7m�b;j���/����p˃��o�>�E"j�Ģ�+9Q���O����C�h�y��Q�:r���+n\ɣ�q/���q=����,+ܺ27N���:�s����A�N��XT�P'�sX��z�;�=�E¦���l�����^�I0콷sh9W�I*\U�Y���J;�8:S��2�L�]��W�<1���Mg
�_�8ku����G�Ǐ&#2٩�eɼyGgV ��r5��Ձ2��Z&���T�uS��;w�j��I�m������)4�1Y:ݒ	d�X�=3���JN����e�em����r�y|�ec;_ڊn�cɾEd�p�;�jEț��	�OiV�gN\�Q�;���O3:���vi�S��7����ຆ+��θ�h�l�v�l��%J���^,s�Jy��.�^"��׵f��&1.�X��YCAj���^w]��s�}iZ��s�P�x�qV�z�Xꈾ�9���4-Ε/��X�1|�l�7nQ��>a>�C6���3u}�<2hԭ��DYO��<�2;ZR����Y��b9Z�)N��xԡ����uv$���r�����ǏiV�5�B�9�%Fs���W&�󦮾]���Q�ZG��.��唤gC��R�V����sŭ+�;+C{C��`�60�g:�KOW>۽]czP�ޘ%�#"eTUx��а�,A�f`h��z5K��î�u2t�,��c&u'���֮tD�YVE��z���Y��%�
�N��'�T���[���5�n�]7�u�!�����鍉�Z/��>�^�5Ց�gV���:%ȥt�j�h��Ǩ�����.��L/�k!��l�L4k���)�5�n6����*������u��l�s��uj����%��N`.�I��h*�I���e��Rɯ����ҕ�idOx���e�$��W�3)�A��ѫ~�m
%�:�]�w;����
��>Uxh����&�h�a.�_k�h�U�L5oE�oy�c��[���d���A���Z�f^�n����T9R]܆;�;]|2�f����ؘ���Pwtg���/'˰�G��P�:V�Q�3LWY�xq7F�{��� ��B�,�7d껹��k*��	�%���|@�I�"�v����=Q]�gvub�!ƹ�rf,���r.�sv��k��V5f*�y���ѳZv.�v��[i�[���o\tOq���2��
�fk|T�8g[��1�~�]��If�{W굈lܺ$�@��W�6>x���ZX|�v�!PF�fr��T��}���ow��ҟeμl�P�uwC+Hk�Vء�������ᷭĞ�����R����܇qi@��C��z�y��:�T�}�r���˵��=\�>���Ɔ��6fnN,�ne�ʝ��m�t�.
Ԩ�\��[�7qٝCF�<�)�,wj���K.��P�'S��;�=�4� s�cw�'y�l1&ftZv-z���g��b�� ���n��(s����E�f�8]:�@�L,�.{E�y���e\T�.�%�ed�rrD��tn)z]!���Qԉ��G�s�>�։cW׍l�j`�����n�┛�M��Ap�o�T3y�(��KiN˖�"��خ�ޙnG�������J�dW�cS���[׎����m�T�b��$8���!m���uŵrq�w�NV�zwt�J_n�Ԋ{�Wc��u:oV��K<	u����pT>W�a�v)۫�n�/��ލ��������YU�X�^4v�Vms��[�x^�܆�j̢,Yӝ����1�)
3JK�Ąd;:�kzǭ.�V뻛y�.'����k=�F̼��c|]kw�{�![QÝݭ��S����{��R�.�#E.�fe�%^��Q���C���wZ,�(�bJ�Px�
���v���J;�nd�Mc1�@x'7+L7]Jq��4ݍ�SX)X�n��SU�V͠�P[.����7��n�͋��ѻm��R� ���[�V�w_4M����jL<ö�3k)�-���Je���;=B�\�cy�tN|��ɗl�n��A��k!�[���#���@���iܮ VTݜ3�Ҁ|�oo�w[:鶵���Z��)��\�%���g_�N�cEwT��-�D��ʜ4�_vU�6���]G��W�������;�y�[�go+͚E�G�Xeǝ��ho'��N2�6���Wv5�\���]9J�}�5���|�^-�*51���W]��q^���:�[�Ϣم�B[X������?ZQT6_��Һ�3�u��O_k����qZ�Ҽ�R��9%vg@�l#;/z��|��f��ԃ��v]����v`��;J��[�:%��.�6+z�a�������vȻ����V�������=޷�b�HHP$�	'���^7��Z���1��Y��z��3���Z�D�Շ����8���؂* o2`rk�cJ��:=�o�L�²���3����IT�7z�/�v(imb⸹a݁@cZ�U�A"�yEb���x��.�#�'r�9�:��3V*y�:�Ċނ�K+\9�1t�Q�)C���l�J�KK7a�]J9�w ,��ٕ��s��8�wkN����^�m�y���ur���gt9���)�������]�`�.7H�j�mm4)�G)��LV��H�}�$gT�ҡk 	������;��S|;u�W��C�vV�JA�)$�v���2�&��‰i��9�������5�vl���1�?=\܈Ѭ��R`#Y��Y[������f�fU�t_R�,I�R�.�&�{�!+:w7�<�Y3o,�:�M�q�b��n�k;\��(�W=��Y����T�7j,P��7��J�̂��_5(o3[�vn�]�}g�h�ǩ.N�X�P�ΥC���9F�*���˫��M��-V��*y�H*ӆ����AJ�ye�	ӭi�'e�����o7����X߱�m��}��&.Uw�u��k�]X$W��T�N�}��j#�m�2i��mk�8q)��ܻ�{\R&�x�W��Xʒgp��t�`,�a�'��ėS9qJA�i�Gws��8���L�Ks`�k�Y�s�*�8/������;BiwroL�V1�N�gQ5��M�_�1�����@�n-�Z�����[�芢�t��]��ץ�]C(<[�j�w�v�Up.�Ë2q4��Gc�k�NĪ'��q��<�� Ʋ�fFM5*�M��m�űVhN�5
:^��c[�һR�Ǜ���	p�o�+muoL�;j�4j�(˹���1ӎuE����,�u��Y����Ժ2��q�0;K�b��v�srw683��uˬ�{.�^)%�
���b^vwk�x�m�C1K�ӱ�^][K���w�.��l�:LXZ�J{
ԇ�pȸ���o�*�OWY����u��wVZ3�v��Qҡ0�u� !Y�f�nZ]�esU7V�H�� �JT��� �J"J�}X���JF��}�6F�%��C�;�,=øz�j����E��T��]t9=q�S���u{�7�������4�@���<�ɨ,�hd�;n��ŕ6��ҟ���xE$g]r���6M�4sdXW�Ճ�r�7�Ɇ��(䂇H�Ah�^a؝�[w�m u>M��]ݗk5.�%�·U�a�N��nY\���(��5Y��q�unY֤�վƛ:�1�!�vR�7{��j�a_2<��n���̘�A��:}I�V&U�4���u^!�Y�P�PxE�s����gKS,��ճ�Әz��#�TX��.��e�u��.tW*F��L�9Iʼ%ɖ��t�k��n���1�×٠p�?��H�)I�B���[H7y���Ѫ�qK5j�ࡧA0�I��ڛv�6�u�yRݼ�m�Ψc��ۮ�r����U|��I6��v�b�V�v<�3����O����͚՜��X��U�"S�Sj��{Y�]xKD6_1�>�kEʐ���q ��fTUވ��D�gݝ�Ɠ����n�Y�&5o�r������;��*���]ZX��Q�3*�cY�۠yi��O\���_J}(U^��	�u&]8ܜ�s3�Ckw4���T��s�2<��K����e�7/��jAѤ��j�i��r��u�C�sh��Yзȑrf(���i�A.;c�f�	h�W�.���>O�y2��Ѓ�,i@I��A^nܲC�QU�S����0�C���c�I.�]W'Lh��L�g���gO�nmo#��ë7f���%At���Z�^��T�&�o��3��-�h�)�Ku>���o�MzU[eV*�g�����@s�ei��4Q#&�f��s^B9������G�*g�Ke�(��\eӾ̳B�D�e-	�E�$p��;��V]1#�i4s �@O�WS`���:N�o>&�h^�������*�����Q�\ �%�ٍWp+zni�e��AY]���T�_R��4�Qh��w���p\�sWK�N�D�B���;�RC������kYA��'�((k[���6�7���Ra�t�>�$M�U���Jm�z�	�(�*sHĜ����3[p퀁�x!;���@3;�Z�#�w���OF�H�A���=���_S��ٓ�X�V�<�b�F�C��2�������KWn*�eu��vUm"��9��P��]�1m�o���uY�X!9�m�t��e�\�T�W.�W,<0䗭�E���<�^3�\��$��f�<��
ܾ=zqyCY��N14%��i��|�*�R�هN��$컬J/���]z۱��nLzb,�J�b�wc�����L���w839p�:*iӹ6�� m�[	�e��J�'�mt�/�c��V���U�#��#��(( ���v"z�[V#5nl�k���D��PP�Gh*W��쫈f�/"��/1��n �7����p�塦�e��+�}��[뵗+�\Ӣ�X�,�=�
Tm]�Yr�V:��Y�P�]����z)� й�8|4f��ޑ���2�Z��G�t��͋���+Y
�8�,]�e*�t��X�+�[p�%�5�2�����e�\(���=b�嚒�@Wm^�,�iI�v�����0&!�@辤��]�M}˺Z�OA3{o&�.����m�o��b��!ؕӗ����&�nJ�ZVj�w)���0�F�v~�0�qs�Î�X�0G�5V�>ܭ��ӥP������z��Uʟ2��ޮ��K�嚦r��ܡ}z�WC���Ż�r�or �	X%<�BVa#7Y�ͺ�vM�}� �WU��5��l�௬��җ�S�����3�kR�d[�m��R����=S�wa�����B}�yb�:��N��f0��������v>Wъ��j�$߱o|��2�ۮ��t3l���G�G��:��)]vl�2�j�^��#�Ҽ:��3�:���0�V	��PX���_�3�`#�j}�-��έ��u�u�z����̓������M�e��2k����j]�EH��������	<���{C���¶�;���c�v�S��eN��ܠk�0^���D��W�Ի	�DiQX�@U�?`R�+]���C�ɶ�e����B]Z�#�8ϲ�CG�_m�އ(�#cϱ��]�f��_b��#�����U{�����g,	)V��t�u�q�B�:YD�N�=v��hfw)bv�������.c�`ᮄ�v��z�@G��tZu�;qV��H�x�Z�y*�/�b��л{E�h�E��Ԯ�6���n�l����Q�m�.����ڎJ֫CK���*mڕz�
\���4.���bDe
�`�C��	�c:aݩ*�",�m�]�����;�woTh�[1C��h�3-R/(K�����ec�%�m�#MMm�x�2�{{�Y��!˳��W�R��[)�:��<�v��Ӻm��4�=swI�����-I�\�nm�S4�(=em�}2W�9I0c��f�3;�ڮ7�	����eK�;��y`�N�U�+�z������O,d���{�{�;��R��F�s�y,֝���w $��Ejm���8��q00��p�ey��۟9���]jX7��ul d[����SۦOYS*�)8�c�a��V���<�ʤ;��U�V����l���ѩ�9�|(�mw�5e�DR1�gp�[�.}���]L�@481Lq�����q�Gj�$�H[�E��e�n��)�L��Q�N	m��}�cQ��j?����3ٷ�)��x�Z��z�v>W�K��Ic�j�]�n��١�����f'��KcHer��c�n��.悬U�xYJeZ���j��㚖jT*�F5;�*�.l�T�\�f}sa�=�>�-�YĊ�����29�	�*�2��t@��]H:�C�z���7��ٝ[��G���pN���^v�J�WT�90�s ���;�l�P���U���V�s:lܬ��U�H�f�ThP�6&�u�*�k����j�SƖ�q:ZBk�za�0�����B���j�]Mj��z�]�[O��>�l��(�Eve�*QZ�u���Gn|�ݖSխ�|����M��ݰ����h�wD`�|Yy��r��n�A�pA����+H�����U�m��qWkv���wa�2�Ua]�b�i-����sC�a����Zlq�R��Q�セ3R���R�e����ʥ#�)mS����נ�ؑV�d�E�\n��mS{X^�}O�?�O*��[5�唻1Ԧ[�z��fK����Jn��7��{Z�,��;��;Zr�'��ӗi}�������t�=�HS�EJ4�׶�8���lz��S�a/�"7l ���s%x&X:�B��Ẑ��U���H���� v?aߕu]�W���NGm������pfԂR�u=M���V5Y�$A:��>�ݔ��B�P78��Vt�WAx��(��O]�A(��W�,��K����DZw�w��4�d�Ǣ��o+pV�r��ugdM>����X�]�������֤�0%"�M+�Ԣ�t]�I �7y��9�r����j�ӄd9�J	XVV��wt���}�XE��r)w��w�݋�+�róCB�!ᙪ��=I�7#�O7S��1ܠ�-!��LZ��q�Z���Q�:Ę-<�NG�����	�����&�|�����Ru�/�����t��Y0k5:c%�%���FÝw��6�12�Nå�zLU�|Boa0[�G0;�l�B5�S˨8�me)�i������6٫̹���{J�b0�#[y
$���/��s�5������]��4���I�:4��.��9�B���B�ٯxk�J��՚�����\��;��tR!q���0^�i������jw
�Fe���yˬeZqN�7�oU}36 �:�he��f`�I�p���)��w�n���ϪmF�:��^o[�i+����WnE-FqA�a�5��J�,歙�;�pXX�5;�[a�~�8�=hd���*�]1#�|qn�7�䩮�ջ�bîp	l�/i}�N�If$�v-[$9�[���F��t��3{k�A�+M�6�ʷ00��V�0)Ws��nid<
��u&����v.Kܠ�@���&M�b����P��Y�9��0��r���8롴8$����ݘN��w�����gJF���b�.��@�I��np�%bX���ƎFՂ���b��$]eB]����,�E';s���i����1+��{B�Xq�E��UЂ���.S�]� ����F��;{7u%VU�Y�~�Xee�������q)ێ�wx�;y�k��λ��Z^�U�*{� ��tc.d4qN�.�݉��/E�W8*{�r�aC�qCj��tN�r����/�I�d�Ѯγ�r��-Z�ސ��󦅨�ntԹ�b�{�U���/�w,[6P��)^u�i�ǲ��h�N���K>�.���2�+�[d��Ŵ�r�̗F���k�iTNoY&8�.�,cH���n��˳�`�Y�^�ۧF�<�y�9��"�1º�sE�G֮��\M�V9��+�RV�����6�������t�4���&��S/����xv^!(��vhn6�5Ʀ(��Ӄ��Fir�
��P�[�gu�P�O,WY/o�t���#@-ϛ��K/iɨoN�� 8!���Ȑ�Jq�^NVm���d�9�4GTS�}��9�4c&���}���
Y�kf&/���kylp��ҷ:�WyYK}���u�BS���t�mǽ��9\��u�Se���`�{�ɤ���� �8���b:�q0ue��d�i�nCO��VpJӗ��*��J�b��N�s���IH\%��rI��*[�35��Q�9����99nv*{�����e]\|'V(�p^��س�u6��4%*�^#;��$B�ޚ�1*ѥB�w|��W�T����a(�����f�8d��>�q�f�v1��ʲ򋮊�������>�%
A���u��2��T�;���Sm/�-eZZ�;ɔ������B�wa�Щ�&�;Ԓ��n��<���0�a
��V�=\&��yJ��ڹ'���R�Z"�_�8cf@�bv��5�윆�5)�qˍf�jv�����R�>C_dJ�d��:ɦCkhn1]�~�\�YK���Wc��h�׎�]ˮ�h�{�Ԓ"�=lLׅ����ȱ��5�^�|���yW���f�<��q=�EK�`��,9�9������4���Au���ce����WC�@_7����5�YE����W� oq���[�e[�7{�v��,�!��rb�	�tD��#�j��Գ������1˥��u��\��80�f�~e���k�����_@X�nÍ"0P���(%O�y.�El��Yf�����m#��Qd�ש]\����F�rgv�R�!M����y��cr�/���[�ĵvu�(���az&H�J�v旘��PT��T�[��%ݷkA��e�R�)N���t�3 �һ�q�2Y��|N*�f�ś}��H[��쥉���}�j]3��P����ՠ/G�F��+r��B��tjZ�IS��
k@��uF�ʀ:<��2�E�dF9s�M���Ww�WV���ޅ�Y6tw+\�?`�:�)lht�7���,�++P7Օ�ut���ϴ�����=�/�#!��;��8��zFF\z����<A�g1*��Qb�w٫/)���@�9NŴ�u�z�Gq�1��j̊�cv��6���VL��	�Ο,ݭ�TY�tҝK�Ws)V�/]���O��U��W�_}��ٶ�E�y��l��_noe�w�J���������ѵen�Z*,ثiM豞��L�+�p��UMPY1���{�e�uk"l
N/�u>p(Jvk5Q�[�Y�z��˝��;���]��M˽�E�]jͽWw��G��ʝRD��	M���6rsr�+��	�d�Ж��*X�L�-���+����^ҡ���A�k�� ;x���;��+]�:�9�ngVK��(fFz�*���+��c��1H��xx���ėY����y[�P���;0Ҝ5�kri��1淦�F$+6ƫEl�*���:��T-�܈��t�9��N� �J�=mc ���K�/8�f+�w�D��b��GF���Cy�e�$ܻ�a-�c����l�r�;��N�on:�kAդЮ�
wҲ�uG�ĝK����Rs&p�����8��w}f�q��U�YQVb�@�Qu
�6����f;=�jx�g� �p-�k�]��R�o���]w.��ȡ��Q�c�uJg�m���s����{M�� #��P�܊��o1��H
�Xr��7��2�G����vu�����AnVA.r�b���f�W	ƒ�1�د�XT$|�����B'iH���Y ��z���W�n��02��W��ru�Ri���f���s1nl����YU���n�\���%��[W��	}�������_�-Q��f"�(�DQ*TED�F�J�+��,���Ll��m�6��J�&e�U"��LaQh�K ť��ˉQJ�(���1��2�Tm
����3%Q�Z̵f5�*P�H��aU-�-�U��11`�$�h)+�Z��QX


��c2Ũ���QLf ,��Qq��Q���m�����*¢ۘ���c�9[1X",V���PYR�(���(�ٙKڲ�G31�Z[1q�,[�J��K[lE-1�`�j�������G)+�R6�
Q���[+֖0�b&1q����amQH�[mchԣR�U�UR�k�Q��c��h�,`ڪVJ��f&8���G��,�,�猶0�_�m��J�c�g'gG�[����j���tV�ʩtz���k*e�ȯUqjY��
��,����UTTuX�Ǥ�g(@G���Y��.���>L:�J��f�i ��$ά��߻��&d�:��\�(lȽ�u�=�]���(e�.T"ī#�IejY5����ӣ�U�%�ߛ��ja�>�Tv)y懥C��*���>G0�.�O�>�BXE��V�*��>kVO��+����o�0��ͿE���37�
W�܎��a��m��H+:Z���]�{�gAۭO|�rX��@'�������om�駾�Z}!��;!k;�3f���>���\�>�r�>���;^�W-�k�ɝ�Pp�o����냞��F�K��۾�ȡҵb���Gyj�a�����[�� v���nW��79�=Ϸ�o�\��}9��N��\oW�m�}��J=�WI�r��#��s��'nS�t(�2���V��m���\շ��h[
�A}�ٿ7�;��~��ڥr��w,����<GFf�g�u�ou�_\�9��\j����ku"��C�K��}G���KX!�o۹ڹ�O1�(p����~"��ȋ5��IafV1`�]P�YLh�gq��HOFnh�Ns�/��(�yT+��'']��\͗X�I�*r��r���}����e��jo�d����g���9�u�P�6�'����yھ�ٞ�}��au�ӿl~	k��֟�rn�Iw떖��@ؽy�:N~����z��Ί\��__W�輆�H���x��{�� �k�%O���~�7�����"#Y�}�4�j�ġ)�k��y��&��-���������[l<�焱0��x�r�J��+��\��,�=�!�|g��m��5�L�3+4I/������c��V{R}y���>�|*���M':��{Y����[��G�#τT�g��\��ۓޓ�^tű������+�g��Oe_�����=�]�kF�����f]u��N�����?�x2��s��'��Ъ��Ƴ�uh�dP{�����g�p�s���x�tl6{]�<R��~���ûKZ0����ۡG�wg�
�us����,���W�:*�	Mh����"�]�~���6�p��A�/hBP~3�*��w�sZp�ئZ^� w�C�ܦj�j�Ume��l�P��
�$�K��lU�^�wo�*��˫�P[�}��uM/����z���=��0ol�@��9�NG���m�Or��=|�gw]�.n�_U���f���r��2�ɏw�7���)�<�c�ԕ=x=�"�W(7�P3o���;�ǆv�6�.VA{`��{��S��{|3��+�l\�RR�n��C����
���3����nO{׵p5��y���{��O`I��L���Y��4ϓ��l�a|+\7�{{r�r��Y�ķs���cchs�0����zCE��ٴ&v���L۩��aO&�2���r�\ks��[��G9�ӏ���=a������z����g�������u->�����%syJ�������.d�~��{n�~�V�cDȀ8s��s��w�ٖ7��~��?V	���U��ۿq>Ů�=X�m6�9�at:is�+�����G9����qǲw
�/=�ggP��"\��!�}a�Vu��d���N�槀��,p�At
��Ug�(��d��7��7k��9�M�k=�`�F��i�C�J��/����z.�\d��d:Wi��y�Xy����k"Ȅ{;,>��&��F!�ϩ�寓�{�[Pr�ݓ�Y�zuz��B�ym��>��=�N�4���R�`Wy��4I6�X����M�K�B���v�j��fs�说���xe18;�Ã��\��L�ókQh!��0f�v�_G��3���n��홽��B8ą��џPs-,[�e��#�3�V�G�uCs�,����y���3zq��*�ncҮ{�S�ry�ο$����S�&�ږ�?5��{�ڞ���]ާݷ>�9�Jm4��෰ߺ6�9�<`�P�·~�}�GS:��s�vZ�Y����罂wo�-G�f�9��=�9��=�W3���>����Nx�������{n�;ٸ#�l�8\����=��k�Fsl��Tx�76^��n��y�~���ix'�g�7,:��O�v���t��>ۡ/��L�)@�T��â��ʚ�_(!�Ͷ;2���v��V��#P<��hcvVG�IP���i���Z��E�����o`(qv��,�%.��#4l�n%�:L�;tx"��U����r�1��[m�X��z��-����L�z����0����J5�}|�g�a�9�s�}4�ׯv�y�8>i�]�lylw�������d�
V�˴����W�8私�0F-\�^-k�6��ec����zĢ�3���hs�Y�v����=嫢�j�e-��o����i�}4l�v�)bQ�gG>�C�_^��=[�����d��k�o`;�����f�����_9a��ZΚ�W]S�Z/s:BC�w���;0���YI�Ț��:.��G	slJ�C���{}�v�F��Sc���+����{��-��5,t��*v���OM��]�mOcq����\{`~% ����t���<�˿kF��V�yv\=wN�jO�1���ys�K;(��Q�ܷ�ݷ0oA§���h����Gj��յ<�ٞ���o&����ՙ�$q�;.u�!����4S�:̤�vD����hk����qpjq�"�ڬ(2��p��/����6a�M��Gb��3�A\�Y2WZ��	��uݤ�Y��gCO[!{��AB�z6��2e6��\r�m�M}*�I�hU����'^�r�}9�C��s�=��9_���VV'��r�q�(ڬ�����}��o� ����w᛫����{�O�ўO{�3�Lo��~^0]��^>�glY�-�}{P^v���|��`���;}3ެ�^��rV��N����W�^��vྨz1�=y�\�f߬nfco�\��λ�Q~�����TW�||�/WZ[�8k�z;��	�yG�m|��l|�k��\�k���/�N�����+�>3ַ��㕅��EQ�K-��c���`G9��lC���Ύ�<tP;%���q��5��fܕٲr}��k����B���f�[��w�|�o	��͝FP����&��d���j�r��,��	�ޓ{f?�xE]�Yԗ#��[�.f�l2$R�vn��]���1�y�)~�$������"��)�S+,e07y����rw��V5�%���R�/,�N�71�[�<;��g&��d��ս��a#��U���+�<ϸ�V���K�FP���O��5Mށ�@�c�j��(/)iÂ� 6�p�s��37$B�
���{zԬ�Y�ӈgyw��V�Κ	�]�Wױnf�:\tॽաTz���d����{�Վ�y?�\vNk;��{)n}u��L��!��ʝ��G�by#-�:�d�Ňx_�g��?r�eJ��e�z��lןw�鵯{��>ވ��HƇ�����V;;<&�n���Vr{��+�k��f�����V���z��Ku�<���ޗ�]	]��W'��Kc��3�@λ]���|=�|6�h�6ǜg%����uj��E/s.y=�{�f���fx�|-1_^�1�o�������Nݭ*�TU���{K���Wٮ�z��]��k�b�1����i.�"�J���"۹�_g�>�I#�.{��Y�һ�/T;=lUS앑�*�-m����1�ws~�t���}4�vI�`��>>v��]�H��Mk���f��b=I�!v�\В�pL�H*��'뮍�Qo��
fQ���'�#�L��ZA�Ç��z'N^�/ ������i�)�Z�n-֨3vkY�o�|Iw0Q��j�����Y�oiDP��y���u�A^��hg��aչ�'zt^���?�.a��=&Ⲷ�Uʽ:l
���m��u�����v�.o-���s��%�<x�}���zU����(���������u�2�<�g���jǚ~�=�-�N:��v;�d��_�@s:is�BV��{�ps��w�7,�-�Nk�7vt��r����Uu�8`�V����Ι؍G�!L�d�fߌ�7��!/}'��q���r�XM�V%�'Y�/eYgiʵ���g�����c�����2��G�L[��,9�e����յ��]�mHc�{��Y�I_]�L�۳3��أ����>�_o�F��o���;n8�U8>���K�)�w�f��o�U�9�jy�#�{ٚRȝM�t�8��ݓ��e9�G��G���Gk����"�5�aI�8�K�B�3i�-��G��<8���/���NoY��ɇ�+up��ixݻm̮��]�+iF�r�ehJP�ZY��� \��ߺ���u»ޡ�-�pc�N��$��$���toXv�5u|0#�|�uL����^ru�� a�4��pr�Y�����>�o��E��|��ݕ�:��r���z���O�z}{c�ѹ~�;���j��{�x��g�Ov�VE�x.fmo��f�-�w��zm�N]���{����>���g%Fn1��Vۮnߔ�/���n��V���6��N�\~�ټ$ٰ��
�T����^�o���=�u�����*������a��6`.s.u}RNԱV��Y}�Z�L��}�����[%���.�C7���fy߲�{���{ے��}���w9��Ds�gE�Xs��ie朕M;vWn�n�g�k��~��Kd�r��D!��Ϭ!��U�b���w�{O�Χ�\�gM�p	�_��ͩ+k�U,;xB�t���gE�ق��9ӵg�(�[.�O�{g��������%ͱ+�UZ\���a{^1����㲶��L�F�Z�ѡ�'m� f�腺�Z�O�ay�<D���ʷ��e����"�U����=ÉK�X0�mb�'��:M:�WƏ���"n�r�V�cm�vZU!�B�[�f]���h�1�����}ܯ3���L�K8i9�T�*f�M)���Oq��;k�Q�V�H��_��Sy+�w�p�>���<���{����"|/*w�5���i�^����=yx lO_3�.���K��Ko,
��W/�{���8�$U��c1��w*�r�|,9�A�醺ͻў�ח��ˡBݬ����[�goӳף5��~��c��'��`�o��i�y\/�Wuu禽�p��y_���~���cՍ�/MR�u�y�S��w�i,]^����v��pe�ދj�xj�^�ޑ������~c�v�}�	^�f]����yn� ���'�B��F=���7��nZrs��|wg�Z֎��ՙ�ۛ�'�QC||����Ke�L/�8h��p��^LRO��N�W>�|*9��E���s��X]:6?����3m��Z��AO]���ڼ����-����i��`wSYB��Ahgm5@mdZ*qS��
�Ь�]�"�ǒK-$զ"o���Y��C	�7EglJ^�a��hnZ�t�Ừ\�o�-Px�]Ku�*�3s+%"D�8����u�lX�ZkY�ڱ��
��3OQ��o��-�5�N˔�o',:��C6ķ�>ЍGE��uz��bt@�K��J[��bI�$��(�2��/�3QI���S*��.��{x��[=V�`cQ��Y:�8@�v����W�v��/g�o7]ΎsyífԬ�W���Xٜ��!-�eJ�vb��`TQ�m�3,��yj�����*�#�/gMY����ɎZ�����Y�x��`�ފ�Ly�=DSC��B����t�;��m��Q*���/�����5�u�I�W"���T^K�	v���G�C�]����oi����P.��W����GP�JJ�o�F�.��|��QK�6.M�k����䫆���_7��H��Her
 *�M�	��E�m�K��[��N�y:�ny����6�4I��\�����8]��[vvv.�Dgf�4��ɧgVɫc˙vz��O6	&>��yĝ�`��f��ؖs���Wc���b���E1k�{d]�9�k���UؔX�}6�[�s��mi���E2��ٱ���,p���p�.�K���Ǌ5�K֌��S���/������ ���:�p���ܞn_��㧭s��;���2h�[*���/U]�ۡ8�{��ő.t��o6�\^m�f����of�6_EY��V�ĻI6�e�t��J3xQ�R[��E�k���֍���w �M�J5�_v-j����+���ם�3j⏤�p�9a��ٌjse'�� ��ǂ�onu��[o�X�%<�ʬ;�.������]�TWP:�9U���̉��5�Ё8�-��o`�O
���V!-u��
w+���]f��2��7+��S�;yR��Cw�T�ZjH2���*+�IhP�cA���;�][�O��Q�t��of]qsEv��`��,�����e#�^�wS�{)#A�N��iu�(ocG��pr�ŋK�9c�Xy�*�r��9��NU�1]wir�7d�u���T�'`U�����!�NG9oc]7W:Sr}�cZӵ�R��G�0�ǭ�n���	�Q�}o�Ԯ�[42���j^3������W͛�.j���Q4�.���tU�6���3h\]����Pm��p��eڶ�\��̵�\�)��y�T���uX�RRⱜ/e`P+��:c,h�D�h�"f�p]8Ѻl���\{7�^�;�(M��o�Hi�3zVL����C0���}�a9ӎj���-���]ݬ�q��r�v���餦�<����7��Y�ygՉ	A #��J�dm+eVe�VUFbf��F�X�+�UChQYZ�Aeb�e��B�r��Z�����c�J���,UR�T�pr�4��b
��*�b�E��L��+1Ub֢�1�hȃ+XV��d�L`�"U(զ[����h8YD�e̥P*J-��Z�,��%YR��W̑�F��X%+R�L0Z�²��U`���ը��*KJV�*����(c*�!�QX�Ƞ�i�)Sf[FZ�`���J�F�2-.eqJ¥Ab��R((�iZ�&Z��s.J�8�¤1�A�q*�J��p�e�QJ����*(��6ѭ�\�A`����R�mL£�j�㖋��s �ƴe��p��-�ģ333)�anfe���L[,�m�%�F����q�3(�KTE�[k"��|Wr`��mn����ͭ�7�!A���t�w��;��w�a��-���[heg�qf���yPf��UB��p�����!~��*W�{�o��~�zQ֏����WOg3J����%Ǿ���%����󝆼\��������J�^�y����#�;�f��t/�^̰y�w���� w�i�3w��ǋ)RW�+ҹ����u���p!��~���s��"��S�1{)�+.;���ܼ��9���X�%gM5P����b��9G���YF!����_J�u�ES�:
�rM�W6�ݏ�[7����>�J����mF�V��[��O������r��x\��]O}��*aʇ�ͫ>�<�k�s���{6`ވ���18�o��9�����}g3����T�}����z����e_�����{e��*�8�o�c���n�m�3�����gX{t�ަ���"�S��;�w��S�i�>:�*v+345�C"U�l�z�x).��ֶ��O���nu�*n����u�	�ΑŃ�~*�O2t��a4O���'[��amR��٧���Yc����K��E�,��f�
C�!&e�:��DQr8���I��r��b�n���M��~[8,�/��\t-1_^�1�|���K���a��/����;Ϧq����⒱Y��W�l�X��w��*롭�4{�s�h���J�N�	$x%�{*�P�5��C����u�3ە�ۘ���A/�lg��#��8M/݂OK4xx�Έ���z<b��M�חω�ϩʷƳ�~ϼ÷7zN}�n�<^�*�,���0�b&z|E���[�.�S�g7=�F��r��A�cBj����������x펢�Ί�Cz��������}��~�|I�~վOgTϱ%���Mq��>~7B�[��:]x;����S���wR���5��mWdL�\�՟\�r�;xu��Bz`����a�r��W�yOo>=/�nj{��O������bU�o	�s@�M���y��C����21o��`v6�[G���ob��X$��ne5�M�E�}Pէ�fg�p59�y���mt���x3�m�0Œ�����LE���+F��NID36�W��\�6��2�tjx_گB�]�{:E3��$d�
��R�f�Rr����z����4���܌DƇxXs��\[*r�ĥ��_v��=���pA�JOZn���~�K�Ѡ�B8��^�}��_��\�n^S��o.���r�<�U���;;�7���C��t����H���WC�u��M89��{^�9Z/%��X�u~��ɇ�+�n�H}2�NdK{��߮�m�6o&=�=�6f�����vz�咅Ǟ����)�ru��:�üv���|3nSr���o�v���g���p�i[��p�ŮI��y[���ɈT|3�B�ۖ�cd�8��̝�*�E�҄۝�f��;"�i�|/��X�ޮ�mvzx����CD�k*e��"��kO]�ج��]��/K�6�����w�:�ƞ��'����uE��@y�,������m���t��i:�~��������Kk�/"��g��5�`�Pv�ݓU�l8�[�]!�G�J����2������7�G;0m�����.�G&/�Le+�̓�8�$w���VΝԪ#Ԓv��Ӭ�����ˏ��|�u1��Ӫ��iW���|��u����wx;�1��+bi��N�5�oz@���z�g~����h�&��A~s���ץ����������ԴI�婿	D 9������C�̇�{��g?~9ٔ�	���;��m�����Y&����sVA��O���a�O�O'y�ޤ�&�>�w$�xɶ����䟎w���N!�sܒ��<�><�}����Mkf���wĕ&�Rt�i�i�l�g�(m������6�2���'��^S�ַrq�l>@�s�'S�M�����:��}-ܽ�M
����^�W���>���d��$�RL5z�������'Y8�~�a8�����M��T:�2x�����&'Xy7�=Iԓ������޿����o��t?�x�%8�.���]�N �|�4�̝7��ǌ��9풥I>��,������d������Bm�����z��ϵ�d���d�����o���o��1?I�W�7_m�_m�u�<d��}�(q��O'y�*O�9�0��:Þ�+�$���E�~���i'����ì�d<C�ԟ�q&����I�&{;W���ҟ~�#O�q��|�O��PY%M��d�G;��N$�*�AI�O�w��J��~d��sVE'�����I��3����/���?~׺���n�$�i�i��4������/����C�x�A`�d�T&�ܞ��M2���r̚d�k�����@��ȏ��G�[w���wX}Ϲ��﹯3�)1�&���	��:{CěB~�S�~d�!��'�u��/���O��s�:�2M3��a�N%Bx{܁�M}I���>d�'y�k���9���y��ⶂ��y������OgGنj�\kV� K�����v�z��H6�<�J��N�˹*L�[D�=բ�mº��1h=�f&	�<�Ue.Xod��{[`��*�5[��u;]َ�f;�O9a	���7�2ueq�Jz}�7�=�~a=`t��M���N'�RM�~O�g'�Y��Rq	�1�h,��$�d�My�8��y����|�w�:��L&�׺�Gy��3Z�zs���O�9�N�� �'ρ�{�Ld����M5'�3ɔ'����YĀ���q�g�:��O}��6������Gߏ��5�+��|'/{�s�{Ǽם=d�0��L�}a=�0�'i�'��$�I�៲J�a�2�|Èy2�|��6�+$�O��Ad�?P��߈G�6c�O]��?~�3��c�o������:s� �i�9N�I:�a��ԜI<��@�O_�=�~�'N'��IRq!��4�ɦ��d�|e1�i�1=_�{�^�_���g�o�|���e�6��������������<�:�ĝ�I�i=d��L �'�}�?B�M'���T�H~-�B�i�����_�w��U��������8��2?}�I�N'�,8��'_&P�&�Y.�8��N�C�wa��l�d���}�4�'�<}9�$�x��w��b@�y�9��s����y�9w�T'NY�+'�,$�N��&�q7��'��:��yw��N$��g0��'�s4�ԓ��0�f�6��?>�u�4r��g���W���}$��'N����N����T&�'�Y0��m&�Fl�O��Z�q�n�i4�ѭ��R|���_x������{�o��{��Ƣ��}�W�}w��ORq�s�M��M����i������qyd�XM'VO��je$�&����	�O��k	�>�Y��I=a�瑩l��oL�O�?w|7���zó}��d���̛I����(~d�<�$:��<��?@:��{�T�&M^0��}@�2��M2v��@|8��lZ?Vu��cV���"��Q�o^�B�]i�I}=��kv�A�gIbkd��f���%�lq}�����z��ˬw���Qժ����a:1�M�U;Fu�v�A� ��GY\"K^5�V!Ɲ����e��j-Lvv�n�c�����X��	�������ӶO�=C�7���x���gY&%a�|ì:�<��O�8����r
d��N�T�$�|��$�O�}�VI����� w�^��L�}�Ƨ鯧�~��?2q&�'P�2?Y����C��=gY8��[βLJ����$����N �<�r>J��}�
O�~�￧�&2>����~�s�}�Y��G�}��$�=�I�Ka�x����'��u��M������'P�[�M!�sxu�b~��u�iY9�Xq�IX>�۬�����}�w^}�{����:w�o�&2y�rJ��m<7dRz���y�8�u<a�8�{�=O̝IĞ��I�<d���?|�Xy7�:�4�-]Y@�I~������,���G���dӤ�o�L�d�|��CG��>q�L�Or�z�'���8�>J��,:Ì'��I�ǚ�>C��A�n�9�|/W��|{y��u��	Ğ!��3ē�=9�8�����:ɷ�� i�I4�9߿iI4�L`}l������q�|�?Xq$�?}�����߾3������o���i'�(��!�M�g����I�9��?0�a��:ɷ���@�M�w���Rz���+'�ڡ����m�e����:�����w�k����;��kn��<g�$��z�6����,:�Ĭ�{� u��2wvI����q���wN@�O�������@<��IXm�ߝ��.x���Ǽ����oCIY8��T��c&��LI:���`ya�M�`{�E�Y8����'��;�k��M;d�'z�}��x����� H�S�k���ߏ��{���m:w�IX|�,�O�X)��'�a>I��:�I4���m��=�8���>�rAd�ǝ�;I2����~!��/ߤ�����~[��F�̋o������e����}=f{mz{�>nC����1m�g/�c�5JοӬ7woXz�I�5~�����[�������.�'�t����T�V�zGSty� hY�7�?�p��=Tz��>Vi]��S�?�?}���Bu�d�5ϿB�M����T&n�!Ri'��N2u?ad�I���3�	�xe�u�!�w��$�o|�y���?}����\>�`i����l�2~I��rN�=I���	�x���~�@��$�(L7g��J��2��d�Q�:���5l�l��5�߻�S7�������k3\��]2z�!۬�`q'���=d�$�ì�0��w$�xɴ��O;�:���y���y9�IP��IY4���P6ì�=�}�ގ�[�3��N�s~뤕����� a��I�̝C�[��I��{��ĝd��Ld�X�r�Ag�{�:��<;�����I�)++	�K�����<���ߎ}��}���%d����O�4�O�L�OP���m����<a��IY�4w�:ì��i��AHk��(m'�,�h����{��|�|�kW�~��z��$�M�IYXO�̑d��I�$��e�����>�z��>Ձ�u����&2��sY:�1?vP�~�	��ܩ������:�su���r�����T=d�T:w�!X|���=�x���Y'>��M>�~��:�����8�~�Xu��$��y�������u��>d@�힫�����j��ߤ�$��a�'RM��q��5�a
�L�י�I���~����OϬ�O���$��yhx��'�)�~d�$zw���_y��������o�=I��7�����Aa4����8��y�rz���d��p�4����L�<>�	�'�t'�̞'�)�u7qZ��}��zs_���������0���8��8������6��/��a��é�$����N��+!��p�'Y6�'<�z��M￉>`x{���O:��P�ZKgĝ��]���3yQ�:�bB��}�1֬�K��������in&e������k$[d��[��X���R�J�N&,�4 ɰBN�SiY��bґvT���� ��1l�E�(�ܓ�#.a=����*Tuf�e�-����h0Ug���(V�w�����co��9����&�4��P�I�T�����N��y=��8�ԩ��N0��u?$�w'Y7����Ì�d��}��_}��#�'��[}�fPΫ���x��IY?0:�,��h~�!�~d�<�f�M!S��è)&~�:�����d�T��d'u�����I���(~?}5|>���;�{�:�����)FJ���>z��?���8�4��a*M�?�IY4ÈT���=�q�|�Sq����I�V����d�{̟~��~��_]����]���U��W��L:]ᴜz�z�T��L�w��3���VH~�Jɤ�!�8���.2����I�̰�M2��D�v?o��_�z�i��������y�:s� �q;M�����R|�Ԝ;�XN'<5���g���J�d7N!Y4��Hi2u>��6Ì��?7�ZW��}U��?~����C m��9����&�:��ƹ�4����x��O7�r�<a���M��M￉�'P�w�IPP��q
ɣ�����6;��g�گ���?}��ad���?O(m��i�<�Cl�Ր���$��s�u���w�m�ORi�;�u<d�����?d����'��D���}.f�,?�|����������%@�'Y8�e��&��k$�|y���c�C�[�ē�l=��<B�w'6��g;�u<d�7��_��Uҝ�5/����H��~�X��~ߙ%J�`}v������Rq���>�'4��h|�m���`u&:d�O���&'Xo��'RN?������Ͼ�w���˭�{����������:ɤy9�	�4���̓�>��%J�a�"ɯ,�I�O�:�q	�S�{C�䞲q���d�Y<C�}u[NySB��~�4J&�]���v��yp>�;#H��(��ql�v�	�,��V,1~�{�W�7tM�nvj�ĉ>�}�C��:lT�j=�r�;Bn����xzH�gM����M[}��gm�҉��K��nrd,�d]�K���A��� I羾xn���˽�>d�����p�&�O����'X킆�=d�;�!R|��s��<d�a�>�+�$��E�~����I��x~��'�u�fxw��y�������i�ORi'y����h{��R���0�$��}ì�A`xs�$�M2�����d��}�$����I_'<����03���g���w��7��}��1$Ӧw�<H���L�aԞ��@�<d��kxI�:�7N��LM{�:ɴ�Nv�q'̨w������޶G�Q h~,�,��*�-����I_�O�l�O2~J����;=��N�?I�>g�N��OC�rM!�'_u�|�����i���:�ĨO���'Y5�Oy���ǯy������}����ny�݁�&�;�{�l&���&�I�&�ܰ��d�<�:�>J��P�N!?O.����Owd�d��ט�:��̝O'��^�Χ��xwÚ�ߺ󧌞�0��6��M}I��L�I�����c&��4ԟ�|�2��?2u<�g'̩�Ad�����'Y<7���N�����z����������}	Ğ0������q�o�'{M�q'Ι9哉'�L��VO�C�VO�8��Y��&�̦2M!����~��Y�]�o�eUh�.������O�X����M�������?M��I:ÖΤ��	ߛI=~d�;��:�u=��IRq!���+&�t��R�@��Њ�QW��~����~|ߺq�|��������4��6ɴ�����'>������?y�:�ĝ�I��=d�d��l�k���d�O~��D|�����K��_����_���=�
ɴ��|ɤ�La6�i���i��m�q�o������d��>5ܐY:����;d�'�N�@Ӵ�G�X��}�#�6�=Y��t9j$����h�O;-٤7��uZ�c�mwH�������j����|�T�q:�`c%�s$w��*��*O��GJ5���6���Հ���br駑��&V�j�L&uTZ%]�y�	�נ
Rw�5({��r��������3�߿�>����2N3�IPP��Vq
ɤ
�u'Y�m'����	�y2��:��;��N$����!��}"���a��?}��;^;U����w*��}w�k��=d�yI8��;�}�I�<���(M��VM%d�(Iěg�XN2u?Xm�'�y���i� �N�?����duD��ضy�t�~��5��&�Mt��L�$��}�u�2m�����N��'����Y'�sܒ�a4�aY4���(I�M��������"���?���
L���觓��w]��&?$��f��Y&�0�;��:�9֘ɴ��h�r
�4��;ܐ�d�~�XN����*I��VM>�VN2i���u�f<?y�����Ͼ�^����:r��6��>퐮�~a�׬���a�d���O�8����r
d��w�B��'�w��ğ~#�}6���������,���Sv.y�=8E�n�;�O4�׉����!��?>�x��=�w�4βz����d����k��L�N��
CÝ�(q��<7� ��#��ٙ�z�yܿw�������g�&2o�%|I>z�)>}@�e�XI��{���N2�)�u�Ĝa����x��=��u�����Ad����ì�J�~�5�Ǽ������;���5��]~��}zɴ�:w�B��'��=גLdߖJ��u>7dRz���xe2O^��?0�	�=Ld�N$���&��>�y���:���y���]����u��ۻ�p����f���:�������&�$�w�L�d�|��&2k�p�8ɦN��a=~I�<�8�>J�0�0�yO��'P5��?o���=_���Ow\�g��d�2x�Ӟ~��M��s�ē�=��d�VCÿa�N�m�O��@�&�i�9߿i�T�k'�N�d=g̟�쳌���5�Ǿ�8E�<̿k�O�O�oπq`�g�t漽����-#�.T��씲�
��A�'�@*}.�Z����*aXc�Dw38]�Y0' Y��#�ڕ�>fX#pvV�#Uj����\�#��VLE�u�n�Le*���o1e%��q-�����'Il*�:�=A^�o�9K
������h�j���6�}�j_j���p��]�򈍙��ZJ,��yW���� �I�|�u@RyV�N$�����Qo,m���t4��VgK6�.�=<N7��P��m���l�DԚFmԫ°�"�����+r�����(�Ӯo��x��� ���s%s˧^���0BsH=���̀�$�X`�A��Ŋ�Ǝ�.l*��`��B:�����Ҳ��r�P���\uuq9�+������K�i0/��I��ҕ�Ha��W{��&�[u{�n�_f,����V���M�`H:��E�3i�V��q-R"��{%��y�t�%t ������@Sz�\1sc#��\���JoT�����Vh'�}�;>�5��Z�%E�,8���]��o���Z]���v(��7�8� ��.*E�η�Y����]���=Z��-�j�@�qj���y;Nhiץp�����X/�y������=H�������n���^N��`=� ��O�_9��y�zf���}�"���w��Zh�ކ;gwA���ܝ����3lÙ�Y1[A�b�=[�
GZұ�0�����ޤ�h�k�����������,���;kRs>F��(3
]z���`�8)ʴ�Q�Hv��O�{y��NޮP��K�p�S+��۟}h��j�V�S��#Y�+pm�����WK���v�����de>�y�� �XaP�:�3����z���U������N��
76�����w3�9�^s ��툚Jf�����6��^McO �]!vgd��#�U鼤�<���rh(Wn*#�k�$��9k��<
��w\��*]��ژfb����7�ld�zs��s�����lѢ��Ҷ��_>չ4m�O�]�֤�b�µ<�]���wv�E[��z���;;�4�򬱝9d�����q��u��ו19�J�'%+Ip�1�2��s7|��֑�`�0��jv$mD�Ğ[���cg�Bz4��f`p�J�v�Yy��d��;�M��}iY�z��R�=���yz��c��Xv�	�ۣ²��K�܊�����;-5�}i�f���^�q��]����T�y���)�c��1�t�0�ڗ���#��)�r��7ooI�n�����������l��އ�F��JU�;)�Mf|\~:�3��+l����Ś�r�*uV��)c��\�ă�е��r����Ⱥ�W(�٬,R�,2 �$�u�"+��"�+��P��9b�ʚ��wp��`u�.��J��z�i;�w܍i�y܉r��G��\�;��3�x�qj)]��:wqK��3���P��yyQ���q�2���E+Q2ܲf)�F�-AR�eV[
UL�iJ֡m��+%QR[jR�QFƔm� ����EJ[-�(Ҕƨ��k2�,�V�eee�b�i[jQ�
&DD+ijQDs3���J��Y��ҕT��XQ*4(�
�eqU��e��ڹ� �L�*��5�iB����Q�E
�R�,Z�jba�Q̢+%,m�Pf\0mX�V�Kl��ܥ�TZ��ieh�B��V�VT�A�k+T���Œ�)l��TA�KhT����[Q�KZ��DQmP�5���J6���-*�D���*U��(�ѱh���j�UB�jZ����Z
�+YjPhڍ�,�l�iF�JZ"�F5�DF[Dc-R�"7,�ʋKiU���lm-Ad��Z����Q���j��R���Fʉm��J�F�
��K�;��YÝ��a��Dُ̕']��@�Pk��D�W��D���]�]��B�O�gP�},����®+�Γ� �f�O<����	}�}4�H(�ɤ6�Ԭ��	�;�~�����?~���w�g+��'�_ec��u	�G'M���źo�V�7�61�iΘ\~�4�vI�?]�k��=�ۼ����13���u;	k����8G�0����罣o0w3doUO+�ה�gͻ=�t��ߒ�u+����������s�]�H>�ɾ�ͩ&���Y�:���oxz����`!ί��
v';V��2�vK���L����漜�dyy3��s�X�B�t��ևL����`�-���9�����Mό���g���f�侬%ܫ�������ڋ����9;VpOjTu�2�^�ןs���.<���J��T�`J�4v^����4xrQ�Ǩ�]������y��T���P>�L� 2��x<�f��E*S��۝���W��<�����5��{�ɯj|/��������yԞZ��������xu��>?]��B�U�l�V�3TA���Χ�e��Z|���*���K�z���@��.泤텆��#�u��S%�[�A�L�Nս3�ʄܚg�&�f�crg$u%��h��]�B�������K�ӭ�%�_���U7y1ٞ�x?�����|���~9,pب�˔�*oϯmy���ʼ���O�g@�x��B��k���gh	���m���<V��|w=�o:�"W��3�3:ܷ���/�����˽״|y����������Z�����S���	�ޟK��Z�Zu{���v�w�������k�}�y_��۲3^U'-��Ի�w]��V�}LX��Ӝ��g�#����{�`�ӛ9��yn��+�qzޚ��x/�n����ٿ7,|�t�^���;F�Ua�jf�v�zr��@ۚ��{�Vxi�q=Ke�V����%C����%�T��F�O��x��iͱ���ta}���E�Z�����
�Mr�D/ܻ�u����b9����6a�z�:(�xC����ntz��l��>����l�=�ׂ��V}#��H���'�Տ-Sh���M�QM�'h�}*�����c������:�>��X0�f��)r�s�᳇wҦc���u�mv��b��N�� 
D�}V�+��m�e�R�j6'+�cا�m&�o�w�V^����1u5���h.	;��V8���%��EM��cP�K��i�!��|>����ݲAh��~�����M�^?w��rs��/�.u��%�X��y�4��u��_Yl:it�\������^��&���=���<�_�_[y�gn=�W<U�ֺ�����b��5S�m�����2N���V�t�ܛr��?���^�y���c�?q�/��5|�����#G���[��X����s�N~O�[���[S���]��{�ר��4瑯8HÙ�/����W�aǗ�c�"�6��AI����OU\ٳ}�g9Ԛ�>�P�-�Ǟ��'1�]WU׬�垝�qh�a��Y��밦��e��T�=�l`����y�}���*��S݉o\�_��ٯ^[�������?r��Ō�fۏ�u�35q�N�b͹���׾ry���F�[g�r[�V����жl`�K�Ua�,�;�\�9R|���G&ŧT�c�R��[��p7���g5��g[?b��U]�]9Ra=�m6D�n�|t,��o*p�s���wjP壵���>��9�O&��k/�G��ҕN�>\_��j#�5߾�|�Ϳ#�2A����wXN\�zw�s����w�z��������ho?]����%�c��$�:3t���2F@���蜖n�?zw���������䷯�u��#�]]��ck���|�Jk�y�o���[{�3�Â�Ia.k�yN����J��{�f��/o�Q�~U~L�=m6�l���9���/�9���-�o���������ήn���{շ�]�<%�#�Ӌ�_�*����lT�ko*p��Rn6U���E/�J��2]�X���gM �u_���g��j���9��t��2�O�f)q��W{>pV��lT'�����X����u�L�:NS6Vr�Vw��p�r�{Z5�G�LXpw�����غ
�mu��n��R�ɹ��r��=��,��l�ވ��{�a����z�Ъ"Ϸ,�����T��4�VnjF�ˤ6.�~�mvz�Ex�+P�[�ǽ{��j史]��t��n��t�'s��3�g�Qu�,g)��=F��bf]�]��_\]X�ju�@���n�ؙX�&���\���z����C�mV|�+y;oO�W���U��|�ʺ���Հ�oΑʡ8�����oV��;�=C�࣡܋�=T�c��n���&���^��'=�m��Gʩ��[���]#�5!��@-���-��Oi{�������O��zrP�y[�FGi�e�x�ofc�_C�v���}-9~��7<�o�m��m�{h�z�g�F�l��Ek�/��>�.���p����m�u.��$�׏�5�g%y�����
^LwHz�۾�[]'l*�pl�7,':g���_���|1g�7�v���^ϕ���Y������|}�#�}�[��e��`�����u��C{b�wp���5����E|v2y�T�����nnX�V|�{u�4H,��G�T���O]T�~ׇ�:!gEp�~���Tr�yqM���;�A���tO����,>>㦼e�yH��|us��Q�̈+|w��̧	�Z܋,2n�v�S.�v�"��Omw�'+T(���yOL��+7c8�"�r����jJm�VMT(�*�H{�[K'0��o ��i�Ż�j��`^+wu4"U�wV�����f��W��U#����7w+�}b��������U��?~������91��z�}3jJ���U�a�=�d�9��R�FR.��9[}w��#�/��~����}w��|2�ѝ����M�����d��`xJ�5ש��u�ӷc=�ؓ#�0.���d�:�t{���K��� s�����g��=�X��3Q�I���*���	��=���x�]�bzlF}A̹��'�'��t.�h�L@le�r%�1��Οo�7�m�
��8[���ѝ�&���v8g��<U���YK�>>�����^�R�Qޖ5������{ofr���M���5�>��{�K�;�ۓ�vf��i��ǭ��q��o��9��ԥ+�	A���nWw��Utz���j�}LX��φۖ��l���=啯�u�W�&��=�c��)���5�^�i�-��l��plߛ�g��w����Cڢ���+�f��	���OGk�QŻ��Nd�vW�@�����z^;��U�R�M�"�Q�6�� ��]�I�6�:�	L�/E\�_2��	uy�ۦ�ro�ů:�C�#���/'�Rۓ�HhgO��!���[�׫R�Kx`-�|>_>^]�9\>8c�W'����W��#naӮש����[�ze���������[f��nt�\�iͿL������[���rKH�lw�������=5����C9�w;U���l��s}�+�ռf󴭭7GR^����xt/�_�>����͗=�ן\��Ϥw:��kn"=^�+������Â�;!���M�^?w��I�7�侬�t��+LVW��9	��0K�	��(N��y��͐=s�#����x?zz��=��zg�z�c��� w6�`n��0J=�N�v*�5<��0ݻ�KWW��J�V�l���:gL����Z,&ܬ��?���a=�b�m�t�9�M����so^��v�~؎��b���g�]O|�r_�X��mw��]��'�ӧ�=�w���m���pt�[�zptC�-y[�;i�[�����lZ�R筄��,7zf>Zw07�p����Z5�UΟ#\��F�RtFi�A�ˍv�M��%M�(%�/MJ�c�q�b�=�+T�4����Y|#�3);ԗV���Xi�փ�b��S7���R�;��6?}�������uQ�p3�~gP=y;t/�߯)���`>�P��zW^�^o5�-�7��ǘ�_)����p�]���[�~�={Lp����
��ͣW
�O36��׭�d��=���������O����1gl�mhk��1sn"۸���#{�Ms��7w#��v
�������Y[qy+�2������{pO�����'.`=;�$s\�����`/Wy�s����F��9\��I>�+£�|#,c�'Lj?M=���^\���X�e$W�s�`;��v_Ju֟�8G�0�sU���}�{���P��>�ý��εy��5�?-��\�WWZ��y��1syѦ����.�����<����[��ػ~tB�tQ�/�9��;�l�����������Ã[~pV�{ϡ���r���^�w�Yώ�>��|_�ӄk�!]�e�;B_G��V)nOx��<sٖ�i�Y�ܑ/�t��B�V(�-ڱ5��"�r��ne�e�TN�q/rk�StFL-�6-u��Jfg�ҹ�h5�l�VS��ÚV�b�6����o��^$�߇�����ϵ�Ni��o���L�C+6I}yr\T�w�gM.�_L/]��Mf�jy���\~���"����Q�����M����u�� �s�u"�K�3��Hq{�[ȟ��ux@�pw����uN�m}^���NZ��>N���2�d�vG�i���
H��������Us�3�t�oyQ�'�5Y������4��,~Pb��Y����ػ��`S��Cc�=9���0��s�j[tzy��ϻjm�v������tO<�������c�3����y͞0-A�P+o���=�ۛs�T��w�on녏���g�},'/��q��7ݩ.�����竳מ�?ߓt5($=��'�k4��oAy��ͷ�7�ӽ�I��2n�Y�y�^^����gOgG���'��j�@V�o86o��{��9љ��T���C)�xf�S�1��.��v+�U"��6�ʸ�*�O�:�o�.j�N�5��gl��c�I
"�ء��W��m^�YmVq���\��0h_4��tr�5D��캿��z������e���XfsԂ錤��t:R���e� �vK+������ߗSmZ�L��'����:�'�%��A�-�3�~�0�߻��ɑ��6?,Z�rw������sj�.e[�Xv2y���|N�z��ǪM�f�O���͟8�����������:#�р��=�Z7�mtv�|�����wI��,Ͻ���s�ˎ�u��DF���������_�!�B��}�s����S=K�I[R丨=�.�x��ߢ�t�K�lXdA,���������[;�ׁK�>������p`�^�_��fvɵR��T2v��n��g<��]�*���h�n�{��7�ؤ>�M��#�4[snV\ϟ�����	�GQ��j�C+#�u/�naU�!o����NS$/M�Ϩ2�7���������e����|�5�fǻ}�4�}��p�1��D�ڽ�sڗ�_`����z��Y�pm�3^��n"؏�e
�Ǚ�U
Y�	�I�'R��;3/8s/s�y>���kIm�} ��걯֊jf���X��& `��i���ޭ��yt���k/RĎ�.5�f���خ���L83��t�xc�+C+��V��#5��­�-'՚��S�yۜWA���_.��%nZ���5Ֆ�_k\2ܲcy����Kz+sZ7+4�5���n�z5L���_\�;n�otVA�pud��d���*��ΛO�C*���%�+:�r�Ưf�4;�5V��Z�ꙛ�E����\�:gD�P�ׂ-Ύ���U�m��wN�u�T�a��i����E�����XXc�%(�W;F���6w����uъ�M��R�w�XN�k>κ��Κ�/��Y��N٥u�u��v4�ݞ��u��I©���Uۈ9aZ��1Uހ΂���l��{|\�+�|��\���]o��$�	2���f������MX��V�a��ɚ�X�F��ֆCݔ�R��\N�e+�Ӻ�AU�V�t&��â2m�m���V����w��T�' �+UjQp����.�"���1���#z�R�۽iJ��l�QT����f�n�@KK:b����h}*���<=�x㏋�B�=�@������Э1'/O_ͧ�y_fw�c�{9%�Y���Wd��W���x`���̮ycT
n���tn���
�]B����j �e#X~�j0�\[]{��s��sS6�-bUh��Mǭt0l��*��$���[�vӅ[Z��
����{���Ǒ�;`�v�2����ƹ��ҶndӔ\�ߖ!L�(��'+�1\O��6r�5<=��)[x�����f�M��$�7e5�<b��l ^Pխ�F}JS�����]�cN��75<Y�	��tWF0]f�[��c��+=M�l~���^��j�[��32���H_#DWIƵ [���)S�*>D���&+Rq�2q!f�˭�r�e\2���c���p�Й�'G�����^������P��iI(p�����P��;��FT���c^�+���ч}n_nl1X*�/��C5�&%�(�d�υ�!�F����<YK�h�ǺXd�b"efc�-��O��sQ�8O9k�+��&�_ -�,h����ل�.�ob���X�����]BeMZ]�)�%]n�Dp�]t-2(Wk�]#��)��PK޾:��c���ݜ˖D�.��6���v^T�̉]���#}2����n>����@�vu%r�#TQ�A��Ys�o�t�������}�X���%l���r$nF1y�<���y�]tK�q����}��:�u��N6���C��@����b�n�1koީz��{k���Gn�)�,�1e��X�΍%��[��΍�ٳ�vwQ!Byy����?
UB�5�E�aVߚ�1V5�ѨRڶ�֨�Q+-J�J2�KeKmm�V�R���J�+Ad�e��V�l���UYj��Ԥ��m�Ҷ�m�R������n�
(���kh��F(�B��E�VT�*#�R�R�R�X�ҥQ�4F��4b��VU-"�AH��Z�eE�k,�V�K	Y�Z���Ad(Ѭ�T�rɊ�c�*(c�)b�����m��т���Pm����ҥd�*TPX��J6ʨ����XQZ���ZZ�Y+(�e��fZ�Q
�b�L��`�Zʨ-B��h��QH-[[A�jV�U�J�Q(�J�U�T�[*�3&"�d�UB�b%A���Z��+H�\��Fұb�3��W�=�k&�:����Tםݸ��ҼSh���ܷ/�L����Y����G B�c{�������'�[�}_UW�|����o\n�	{__�f���{����<�9-���ٜ�������_���.���Բ<�;�u;��1e�1��@n^�q���o�yS�wk^U�S�������0�����Ll4��������-9~Tj뽷j���Cp��y�۝��;r�/=+(^��¶Ac86S8���k�����������
�:��N��t�L�v��b���.�y����o��(s�0��&	����`ϳ��T�9@��yۜ�b�~�����I=�$��V#���6�l����˕�>w�d����nϯ��>��n{�l�s��ys{+$w�]k�qY�d��Si���w�}����_t���p	͹9����#�׆�񼙮w�����u.K�x%��.�M϶�s��_el���r���X��O#�ku��·]�2�Ww-�ڈ�r�m*�j�X��f
�"�(:��5�E��K�عVF���2v�d�jźk��%�F��B�`�ޛ�{�ͷ.v��^WUot� �)�}N�!���Yú3y�!�����}_}_W����p�gk>���_\ە���u�8��4U��mƶx���˰���Θ�蝎�EO��9=�`?��{-vyP�hM7Xy��M���y���n�#\��Kb�E�Ϝ���'�ۣp:�-S��V��+�t+{�y7o�^���z#_y�ht�9��z�W�4�$0S�^׵4�>�Z��ͱ�=F^\�~����c{Ӄ�}�q�<���=0��b� �x�{o^r��9,��e�v��sV)�G3S$�T��I��9f�DV�I�ߏ���NUO�Lo��;W��[3�mu�I���U�~^��^���r���{�}5��	����m��kֽR�~.�gǧUd�y�wݹ.z2ވ�E���>�C����}��oW��~��F�5g>�i�hC��!;��ol�E�Ix�dо�I��D�W�1w�N�0-�S>���Bk��*�X���txEt�8f�E���lL=���F�Z���Ԡ�}Im5�o�m��H_.��V������k.�HF)�x^7��Ӛi�.�����b��m��՜֜�%�TT�ò��I�G��7,�ܾf�2�D��:�"ݱY"o�>���}U��}]U�V�LD���%�g,WU��R�/.]���4��A��:%���xV	Bs��]|.9)�k�s���ؼ��栓��ϕƒ�h6ئR�/.��r�?"�B3��&j{�|n���׾���Yv���{qZ�,d�pO}�\˯m�6W6��dh$�S�(s��L���<�{�H�˱��z���ڳ�.�DN~��OK~Y��g0J�&�h��h�/�
(^��}n�g��ž�OJs��(8��d�|�R��?�_��Z��!Ã�k}g��\���������^�s�gDz�����c6����ĥ���9�mh�%��%�t�zAu��[�O~8$��G�X)�"�UC֬�)���o;����]�p9D���ǥK��͍�����)5>�\����>������ym�UL����{TŃz]�	�+k�S��R��{'����x������>s*�vR�u,���r𼿛�4����q\>��d��l���{NK;�0�/9ރGѻG�����dR�L���vV�x�K��ӈ`��c�M�d��c���^/��g'�zv"�ǻ�1V�][ݖ�C֪�N��$ r�Uã-����R9�KJ�m�2nM����� �,9���y�˺���Y���p6Gp����"�1��u�Lԥm��A�h��*�9�zA]/Go���2y_��M��}���ǹ��d��[J�q�"Rgi�Wz����|���G^�w/g�X�En1��w����<_���wYĠ��o�۾>�V��m�沜��%Bҹ�p�-~���b�v�L��������WF2�R��*��,�J��;&��H�y�I�L��ܼ9OɃ��#��{|:m;��y�}�q4a�`�ċG�,m	U�x���� ���'=�boy1�Tץ\�%eHVj������Zh3du&�=w�x�a��P��Ӓ�౥Ûp��&�Xg�);-�ֵ�=h�]����[A�:+�Ċ�.���띑O��ۄ�O��.<t��K0d�pL��W�4���؋8%�&�r�#eq��[�ِef��э⫫�x,��"g�s\|ab{�n/OT#/&`�Y���/�ZCu�F^���wV��}����	�|P��M�	�>��O/�O)��yzB?/COD�V1�7s;3�u��xd~���%t�x.�� K��Զ/�ֲ�\/�+�w��x3�Ԁ��)ݻX�<��@c���z��<�Ľ��{���LX�gQO3// E�rR��rM�����r���1�^�~#�[�zS�}���[n5V��s���ob�j�֍�J|ӭ��;ވJ�ȁ�t�un����Xȧ}3��R�a2����K
��������mﱾ���{��?�#�Ik5Ğ:<���ja�zN��y�T�B��D�N��[�GYT�0t�Pö%Q�%	�v.�-��a��dY�f���D�o{'I�$�q|���~_��F��VX7!��GH��Taa��NG��)3��<��'����To�G�H���μ��Wb҆�Ϡ�W�1��E��Y�x���g�(�������ײ%8�{}�9w<W�>��?�7��f���s�#\=�_$�+�rBb�d�'�5>�q�^(n��s��ϯk�ǥ\|LO��x����{́��q�*�Ot>8J���\�bm>��>���8�82E��:)�f�������cx�kG�c�
�]�ܝ�t�����7�MC=�꘡�`\����8��ϩm�Z��_Vˀ�R�_���4E^�{^s8�f�P;z����rǌ�O˦m���3���[j"�{��Gh{,��z�K��+��������,�9C�9|ׄ�Cݛ=�Y�4���3D@���ar޲�\�Y�}|�v��5������l��T5��Ȫ���fS�v熠���;^;-}�������s�����3��:���2טdxl3r����ʺZf�V�TfPL�7�I]lGݘy�^[lQV1X��
�����J��cM.Yu��U��]��'zU��/���U2�ꈉN+��qM^�F+ϲ� \\׽�XdXن�o�.f�-nu��1h���
R>\dYA3,c�/ ��Z�nmh0�'��N\�k-�X�K��D��]T����R"X�}�%���eϕ.u���°J=Y�]�5~z�3���wT�rA\��u���oS@�!t5�X��v
�_�Q(o�n�~~���)3�:�:�ہ�C}��Tŧ�C|�L�vVY,��HB���Z=�Su�i���o/���9�vw6�����F�Jȃ��+���
��>�!ۗ������#���e����e'�u���|�ձ�י��x�ܬ�b��$�V�38��d���]�~��QN���Rus��)�va��#��.�����6�9�.���
ܰ�qc^Ih��3~���6��Y1;��&�!���"�ѳ���*�P�t�z->#kU`���i��ﺰ�
֢h�߳��;wu�+��=})L�l�N�xd^u��/�h��U��}\(���j5�1��z��e�bl׮Ѽ�f+���qn�c*Qb�:�@rd�6 �5H�J��//[�!8�G�Swݘt�u�]O�;���y�![�z��=N����n"�Z%�ԋ�-��E��O�,�| ���ik�-s�9�'�ΜѼD�-�©�w'�w#�M�Vb�Mg������r��u�Xon�;ٽ�F���f`�b������2��	�^�U�),g�J&�2u�=��T�p�͐�Yħ�E�p>�Rj,�C����|Kz�"�s.��U�����.JQ>|�wӠG�~�,LIxyy�ꄛ�Ke`��d�9O˧gZ�F�?Yt��+rd���޴@������I�s�)�L�Q�&�/�9��t0P�,�mU������c���~6|Ė���-�"��N�.�?,	˄z�r���s��}-���R���D���Ίτ�<��}(;V'z��v�dh4�sܾ��tha����U��]v��w�-�ν�K�-�~��OK~Y�'���^$�,�y�I�G�v�6��z�5�nnhеO��yL��ï~R��?EB���*b�p���f�����w���61�i�>P��dq��6��}]^��LTɁ�Ev<q�6�`���kj볖�>��+�bY4�G��U��0ӗ#y%���tmr}���.,�E�s�ľ���8�[���7s�gv\a1�:gT��X���JY�S��:<@ᝯ�,u={�0;�\����.s��󶳮㫸��{�s���W�� >��7�:��Z|�I%�Dm�㢖R\5�/����0f�D�axe��{f[u����c�����0�����{قx=��6O���\}�Lѣ��MhOٖgMKȈ|����q��zMO���&��)�lt�|�U��z�҃!�vz�U�|+~/+xe)���$F���)�n��>\U��������3�s"��d�6��P�P�ע%�V�}tOIS���o=�H����[�}�cb��Zly�i`���ݲƞ=w���K����s�/��3�2���Ҽt����s�ZC6�sY�9�7�J��<���kN����6��&�jgwC�ښX�q��D�d3�s�OW���q���L�����z�Vmq+{�_��GJ	���=O:����ו�8�iR�/���_S��"^�hvHHy%T�t�;�����NmN55׌�r��!ai�͑Ԛ(l��t���%�
j׺���^�\�<[l��%��cL8���q�r͞�{�,�Z�d�d��9ɭ|!��%�?_GV�[�H��(`���1�Z�V����;s�ТwDмx�v�����/u�Bf�6�϶G�I�>{��Gz�9�.�z�8٤�"GՀwUCV�:��Já@��B.�L���W_��x���v}��_��9�<�?���^m?Lsb}�F�������|6a0��te�nSp�/>��E��Y�h9K�$��gs�UPLǓ[����,���u �����~Lr��;�)�w&`�X櫄66�-�=c���I�ޞ�a�H󔼕�U�E�"��4�=6�:�k�=zC�W�qKB��w��	3��5̙��<��X�=h��#�]:��S~�P�x���1t|7}N��u�3��;���������\�*��x��b�ϟ�$5��xS�2���Lﺗe�����6J��.�����E1q��h�pS�L0�$D-�4%��J���~��o)�P#����O=|��(W���.�F�������԰Gh�1Y��hNGr��w��{-�Lp�h௤�V�w�4�*���[��$�
��c"�Ψ�=�Gq=O�J�ؔ=��[̜�GGYZs�ڇsn�ͽ��Gk���Ɣ�+��Vr�pv�N��{sӷؔ��W��!+-b;��k��J��9������u������\��?B��vCp�,L����p���{7S�W)QLؐ�p ��S4��O_�*i��#��#A�7Y[L��
�$���`��-u������ �Z\�>�b/��G]`Z�TV�uK��gp{���ۇu��-�N��u�ڤ�A���\N�π�}�ږ3Z�ў���w;�_��o(oM��-b3���M�e�x�MLu	Vp8�a
r��^N�휂������3���wV�'��=�:rq�Ք��-H0B����&�s���]�r������Ǣ�k�f[������8&�z>��ȵ85N���v���MA)�<�1C�6v��u�� �
k�%Y�Zk>��Y��(p'/��h{�g��*�f�7�tHH�r1��{�V� �X6�B���O��x���l����g�pK����od${}wiMq�v�a�.֢�<=�\dYA31���@뮞�a�/���̖�0�+��iޱ�w_���t�}H�*�<Z^WS/(S2�SJ^;di.���|kN���N��^�[�/�xy�j�����-��P�C��J���vP�z�ʉB��J�B���&�R���ޯ)�,k2�w�����(o��2���_��p$��������d`f����ܝ��TG����뗼9���Ҳ ����Ttt�ؗ��|�G~+�E��yƖd	d����q�㕴���C�5O^<���-Wp7y��V�[�j�(�['7�+[�;t��N�5�sf�C9�-ۊ���Ǭ��u���WN}c��F�JG�<�t�VA��鑛�"�q��<N��芀��Y�I�R�V���X�E=�\P���o-N�7E���	�vn��:[[&Mc��Ͳ����&�G�'-]\���cb#3��v�S���e��ql>�'&u��D�MFx�N������;�[�v\�E'e�<S �6��N�ke��K:s9�.����d����J�� o�e��=�I�8�Ɵ+��e=�Z�V4�=������x\�IP���)ۨtS�5q!���5N��*�*���F�(��p>�;:�j�.-��.��\���w��j��y.nh�^��L,�O����EPrÎ��O�F`{ˠn����Ÿ���"�f-�O+3�y������e�_k�)�mO��&��+WM�L � �:3���EBG�gTT�3�d����n�壏K�� ��ѺU�K/�ﶮ��fv� �j�ʇ��>�%�y%�xz�q萅nW-Z��y�t��V㮮�s9�z�u��#� +�0��8�i���6�
�s���!�ka�A�������cV��l�\/5U/:�OB*Zg�i�4��&*}s@x�,��3s��9�[�2�C�X�n|N���zlV��!��=�&����L}ԥc�~�Ux���zD��Mye:�ac@��s6��z��뺎�`#�oz��̧�5ԗ;xQ�E��v�S�b�Je����6�}ș݉�&���m]������FF,���@X�$��+�E�`R��z�N^X�S@ʳu���]ȱ��Ө-�u3jk������ʚ,dQZ�,�-��0���A�k�^�rN���n�(_u1�}�.��,�Zm�*�m�ug�ڔ:Ln��-W�rt�\���Ueи�K	��yW�Ji���HcL9�򳻍_���9=�U�β�	 �f��񒌽SjV45d̕����I3E��Loq�P���n�����ӝ��޿�@�{�5�m��ԩå�f7/�TУ�Ս=#y�łH��m�4����G��Jm�T��������;qm(��������诗K��#�VU�N��v���Vp�9V�gv�����Ep�׊����2�Y�˦?����W�Hu�U,ߙ�()�N	��x�*B�2���k9ф5NFܾ�GV̮���T��{_eᜯ!Xܫ���%3��8�^��#�K+w��f�f\ ���fJI��y��8���r�Zl���ō2S��#ݥE�	�R��7��7h��A9�;k6>:���[ԑ�B�Kkt���t4�4�����P] �Na"��J�BM��b����f�g���H�XQ>�$X�4([I]"�{�tQ����fd]�}��~pn[�L^cK�+�
µ��F,����-�T�j���j�UZ2ڍ-"�hU�ʶ�DX�-mb�b)c)m+e���Q�����Q*��X��(���H�(��Qi*6�AlTh��e�Qc[m�S2��*���,�b)�(�T��9JcTX�ij��+D
ܥEU�V���X�X*�S-�����Tb�Ub�5�j�(�kh��[h���iiD�Q`�X��Zʪ�J��DQh��E�b�Eb��mZ��b���YE�Z���V�6��J��U��F�m�E��Ѷ�4cj�
%�[aU��TU�`���A��5�m(���X�(�Ub���X��l�%h���,AZR�j��(�EAUmZ��Օ**��"*�Ո�R�"�R����(�kQ�0T��DaZ�E�X��-�U��)Q�*��VV�UU�QDb�"�UJ���P��$˼N��r��E��/�1ۨ$���t�B��珌0,z��cX�����q�h�{"�ҭ���	�����X;����
��^ܿ�3���k��ǯ��|d���K���%�\����Ө����"��NZ����֍�����8l6���������ޕIy�As���G�y�U0�_����ҫ����iG(�{2��6}5x]U.Rc��k��s��U���RF��a{�G��n, W�����5SˍakB��{*[�������;�f"1��E񾅻U�:��xm�+��Y^[M��ʞ\�Z��������ʰ��8Y^6�q_>�ŽG]W����n[3)�ŧ�B�Mu�zwT~�;�Q�"#����]���&F�x��Uiicz��9��L��s2�ޯ��\˄ya�)�5��+rO�9g��-��M��U�Ԣ}}P�y�Keg�tb���Bg��zyҹ�Rw���ee�Ŭ��q3	���_���y=���0�~�(?/4K�.���vt���}����:�9^>o,�����*#� �KA�o#��K������Vԕ]��[�*�����h%�2ľy[kJ���md��*���l���m��:~�h+�a�bW�i�]f���<u��;M�X�r�9���4�V9\3ڒob�7�f��˼��mӛ���D;��|u�)�Ċ����f�%#�a���ϧ�hBW�l�.�V�������k��50
9�2����>�:�Wrf
�X��uꗤ9�2�	��̺��yX����� �f�6�<B��~ҽ��0�m��;�>].{��A�EB��J��<L�	x./`�c�}^�1l�<�e/%uZGR�C;C!��k��;��ŕ2`~��x�r��{��ȮRf��:��o����zp?RJ��=��+j���WȽ4��k����t��\'��Rd�x��J$x�K�̻��P��G��^Z/-�	�qp���s�5}��.ʮ�f?z���	��h�pS$��ȋ�D�]m�f�m,�x�L��f�T�:�kބ������jAЮpv }p6<��p1=J:Do�n
9�>��2��~Qfڈ�|�k��޾�m�jBf݈s�en(=�cb�r�X==l�l����Ҹ���1YGln?ዤu�h_�����rr�u1�P�
�m��S��b����܅�;���lmλ=�8&���9��"���`���~�q�*;&h#��������p��yسyϱ�{X+�Ы�M"��
�#8;=��J��ngw6� q�����]�k.�J�}�ޜ���<����03%"��<rY;�H�gv��Թ��X�v��݆M����¿����]f��nr�w���?-65j��v��R���B��G<�$��30;��`���8؂	��X�zj��jy��z_��`�SH���K�0}}N$s�T�L�u{����~�� ��U����^u��Q�	Ʀ�>WKP��f�#�4P��w��sw[���ko��n�P?
���	�2X��c3��]�֏g��o�Ƹ	q�B����{�εי�}~�;��(Y��	����(�[�\4�Ξ�Y�f���}i�'�f�.���8�V7�q���v/|��OV�Za��~�����MBD�j��vz��#�s��
�}.J��f5��dW�ƃ��X�C5ҙ^<�Y�.�f]ߧ���y�o�Q��v,�����<�<���.�]��U�g��`v~��AX]��.p����gG�_]���;����P��P�;d�Y�i'��<��uja�~�\9s�/��F9�_�]�0%��ۗ�x�_V�6২��.�q����H��y{՚"�G7$8�6y�Z���W���+9��A!We���JCY}{��t���=WR��ݏ�}�J��e�kŚh��=�i���]��uA�mb���E�u�V�խ��u	zV������#hQR��������w_	`+6;��ꯆyMS���3���	�~��eq�z`���Vz+,�COR������z�wQ�A��	���ׅ�GN�T�[��G���zX�AB��c>agV#��w^��>Lz&�+a�|�>�Q���!��vn����=Ly�^��N����r�C
��{ʱ9���ey�sM��<Mt6=Yױ	��C����c����fմ}u�DX�3	mY�81�a֤[�u]kx��z��Ǡ~X�?x��X��tSg�YM���51�0�{Tɘ�w���o�c�;iG�ǰ
s0�KP�Gs��({_�=�:g^[Km	��Wެ�܇b����m�8[��zp�1mgw9C<pMv�=��w*�6��3SH�*�W���s^�yt�ϩP�,W
��΢�Y焲��R��	Ƈ�fc,�@�{�Ev���c4�f.��o�Ȓ\f��#���V�⚶#ϲ�5�<��lk�W��w/J�a�"|��v�XN���ł�fc�-!և|�ۛ[�Lπ�t6ș���6��f�V������&�Z�6�̭ ��d�;�Z�+����o1k�o{�N�E='i�҂V�:����wx����@�fo�	�	�����.	��ߕ{\�E�������[+T
��v=·�4Ϩ�	c}��|���\c�N�����i���D��4K�}ɥ���e�
f^SJ^;di\�C^,r��{��o6�h�q�-b��W�S���B�֥t��A3ݝ�2�_}�=��z=�@=~�7<���!�U�*Z��`�p�K������[HM��ޭ�����s|���+�v׮�>S�k�s����0Q�Ҳ �~NGD�!��0�B^�}������n�i���Z:1ԗ,n�m�JD���U����y7LsB��p�["���Zw�� k-3�����H�!�Y�]3W~�=�CmC�*�󂂡�w�����r���\r�\��@H-�?"r�,xԔ�J��^����Ϸ6���0�y��M�X8�ğ���Ǎ��p���I�W^�p�\kSZ���	�~�mK��ڞ��o�UUN���:���賽~���V�{�����
���3˕C��W�z��af�LF�{�o`}HZ��B�����}�ļs�|�/VMw��^���#��Oj�{GE�� ��S��7�4)C�o3��̈J0�W��z
t��s{<i=:l���v	K�^W�����9ސߩB-`��<��c�[�z��Z�cZͳ�ț���Ej�Oz�ǵ�3�Eܑ!B!g�Y5{ �T�V�R�.���r���B�^�����}�t���r��qĽK}TΥx�
�����-E��qXw3!�]-�}���{X2{�xns�6^;�F�Vo�Ҵ��MhU�`,��	9Ȗ��:1	:��n��Ju����:���f^y~l��x~^�D�k�-Kb\��W�˲�4��A�9�2�O*���Z�a��0�|��+�{Նl�/�v*��X6[��n*]n�[�nO@{�i��S��|G��ɗ�f�'�l�8֣����͚�
��w��+j��#��-u���iU����r�?,	ˇ^�/Hs�e��ߖzz�Ȱ��4NZ��]���yt�M����I�3����g�ߗ;�^�/ڃ����H���27%�O:�gM��Κ�{a��O�ُƑ�%�T��W���ÿ�o�����3�`2`~����ك�����X���H�{8�]�Q�s��'�W��Fً�E'Ip�E����'ך�1���B1�w�s�����_Y���3�<�%/'2�Mm%�꺏Y>:&eS|.�� �U��yc�AC�s<�*�)����sw��ͯWyWW0��![�C��S�0u���Jں����Xኳ9fqǽ�DGY�.d���Y@���}�g>wf\r���X '� �^�ᕵx���o��5n������+�� }�g�-��ڽ����V�a4Ѝ�8)�lGH����/�Ѕq�V4Yy��87r���f�2��B�^��W�O �.*�}p7�#��OR��雂�w��;{(:Qi�}�����:�S>x�9�a��V�cۖ6 �^:����S;�%�<qݜu]޽�9,{C�J1��yևMW��	~>��͊ڴ�4����J���b��8�Y�׭�p��ű�)���r��7<s�a��͋�"U����k��j�K��}et�ܶ�L��w5z!"z�'���^Z��E6���K�A��-=�B������Pel��
�J>�"ӝ�x��h{�8��^3���\����?rM6D�e����ޙ�g���jPy�fo�a2�,i�s��N5�X6z��wh�k�p/����&x�����E|�"3U�wbe;�Yf{��&�'<��+{��}2�g(q���G�Ӵ�͙���L����aL�AY�R� L�è����B��=tw�{�<����
�Yk��	�)-@�`�I�f��3�*H�-���m.��uh�,�������D02�C���c�KB�]!��<ũ2���t�in	ٴ8���`}V��mw���d�$��g�n�]5�	$"�-�̫L�ʙ�n1
���av�W�-��_�}�����"Y���SM�S=I�-K�
�cYA2/�ˏM�:�k����3v����5n�(��u�r�i�z}�N[!/C<�:�н�F��\�9��5ڠ9|��8=B�y��,�����)S/��Wl�R�z�B.U��$(k5�&���w�o�|��b���{�o3;\�ny>ܿ"�U�K�?"a���wdC�?B_�* ��fey�w���]�S�s���w�^�z��Ϸ�
V�j���nCOR������è���]M�9ӫ�AX8Y��Cm:GG^+�U'�񿳖�S��c�}
�9�agR�C�cK�q�缚} ���脡A�Cl9�)��p����s�"��,h�g�矶{kލ�ෳ���﯐w��D%e�G���m:\�z���'�xE�*�ܔK�������<�U��(ܔ�C';�POV��rӛ��Y���]�����Ӷ���R	�t��ŧ�ǹ)�ļ3����gގ�uLP�s��'�О�3J���Z�g����l��x4k���)�uyN��x�y�yb�k��l7�L�)}^w���h�n!a2���|tZŘ����Չ���u�b�F���K����֥�����
IB0O[��c}F�{muX�R���p���Z�ڍ��Zޓ7���������u�]�~�>�����!�c��G|�(Z{a�a��P���]�NeC��]��f{���y]���3*iKq���I�����!�=o@���-5�y�,��NP�u/���C�s*ɱ{�W�u��2ی7�n4�H���r �h��2�#�*�`.)��l��}�olE���ݘ�����i�f*����0��k��H𲸸��f^;��
�؅�v�ը1���ߊ���$:Οk{�7>�|׭xD��,K�ɥ�����)�yM)���qd����:{ux�1n_yv�w��kya����g���Xg��]0�G\l��"��.����N�Z��K��\�����L��j�-0�Z�L�vVY,���$P�O�����]�0F����F�����W�4��K�^�,Qc�dA��ޯ �<"�{��;��o|������t��FGb�J�TY�����QfoL��P��3&{�;:-ҧ�����ȭ���Z:�c>	�٨
�Ϛ੻pmД6�;ҩ(tz�۝ڮ��yc:&Fe��SU�J�,�� ��2)��B���7E�h;�y�[d�AȮD���0ю���u-|.Ef�����/^���_��,���./!�bЪ�S�Z֦��[�=RZ��mԝ�h�lwK���K#�tW���ev@��b�p�����q^�l���(,��Ҽ�{�4�ht&mj�*�>LpU~���;�$w���/gY�}3�}���=a��j��E�2ޕ��yt�b�m�g�WQ�2/:Ы�QR$�^���/�oq}�v��U���e��u�8�x����S���\�Z���~��E��4�[t�/�N�zs�]qq֊z��_Î�}�l��b��/��w�L�;���a�>?�9G�8J0��Kʹ����K C��7�E���d8��̇�.��g���mN��keJ3�����+
	��Q�K�>Ih�~`/���&���F"���滍���;�+{��bΡ��\���L�P�B:�Z���1jc�ȭ)����Ă+��57�ڊ�o;-��>�D���w�D':���w����P�R6[��x^�n�\#rڠ�u�=N��8�|#�G�Q1���h�޼9���V��G�;���#A�:��#�ٺ��+���@(P���L让�\�|��^�a�~��	�o�==l�J�&��{�˓7�4,��Wu�U�nR�{��t�Ӻ��;��;��_rl�����g5���Ӏ� �r4����y�[[�Σݤ�C�㙻����w������f�v��2*j��m�w�=@������F�8�b���L���A�mVC��2�]r�0��3n���ݱe�`�vf���f���՘ �8����7��¨'��&��0�x6�S��ux���Cq�<!+5��,��֦�w�X�N0�f+f򢘂�cGRچ�*�޷od���ٗjWk��QA�����B���S(��5Sn���h���/���g9����O���z���W�0�,"!�6�vr��ڻn��Z{��%�R�vfVv7d�Q�J�cI�p�^T�y�E���	'V����Z3��N�C3�H}�L8H����uq��+�`)�݋�O���jt����W�����wc�a���iȏB@�{�ĩ]l�'w�}*�U����uٶ-��� ��M�f���wQ��Ew�/A�u=��1I\�&������{������6�A��93�EE��#<��p';s��x� ���Wc��
*��S�2Q�gP|d�0��ɓ��i�"˩}Y�-���k�k�}5t�Q=L��Zj;�Y�P]כ{���Vx�9G0X�V�ݾ�or�G����2�uQ�6����P]uԅ�`niE�r��&-�Y)�\���+l�I����lw5���J�v.���2l�f��ub�%��� �����
���"w�H�c�x�
�[�ve_H�lN��b�!
ų�G.��V�A-�������9�4&���#�OfB��a:�T�Z
����|�OO7!�Sx^ۃyb�Q�n�wL����v��Lu�d�S=�	�,�u.��0j 5���nR0�,�uj��4,���9nS��3k�W6�I7�)uZd�U9�0Z�C��s[]�Ef�^θ��pu�cҴ]����1�S^%�̻�QPov�PG�lN�k�^$�ku<y{��2�i�P��z���Mۢ�̮���v��jG�n�ĺS)*��.{�ô�%{*�� �x�m��+��0�q�tp���I�/w]�Ҧ8��9/i31���ST���ݧ��cBŮ��Gj�7���E�x����b�w����8�u�i�,�
���V�wh�7�S/�ShiG�*Y�޵�^�MxEKjA�Ŋ�����Ḃ����9Ii�k�*[u5''v��p؄c�M�p5���¶��8G��*n�0���za��
��,ѝ�朠���o��fU�أlG.�%��z��uc�+ޥ�T�9\�J߬^�Q�ې�gNi�S	9]d�3��������C�H(A�:����&P]M��>���L�H��&��h�~I�w�ם���{)��ek�{�gR���EL=}]](��EAVZQcR��0�j1EcR�R��Z��h�eT�ZT(�аb��Z�Z��"�)�������������eAmF�T���-�kJ��i(��XQh[J�(��iJ��c*VYYX�[j*��AQ������T�AD���X�J�TKJ	mDQZZ��`�JYm��QR�K-(��,Q�h�X�eJ�b��X��J�QTT��m*+`�#�mF�Pb
�Z4���[e����0U��"J�EDF
�i[b�dV��*��,PT[`U�m���։*J#h�U�PDUQA1b1k,A�������E�-�UF�Z�Ŋ,X%j#Z��TJ�Q���"*���b*1�V(�6�YY,��h#l�"��*��,[J���Z��}����\=ׂl|~���b��|�����4M����60����о*È]�|A�E��7��<�]�r���u�1C�� �7oq�,2����'�2x �	���㺰��ת_��_�	*b��f�
�.���X���-�x��x�Y��\8�#@s��$��^!����ͮ����I۱;�I8+�jڸ=)�S��8���vZ3���%�pORJ�R=�
��U��e��3�	d�M��W����(��0v�Ϝ�G��%/+�f	�{@rp���囟U5�)�d۽��-����N<W�lq�nX���w��^��R��"-���S�l�m����-��x���rz�KX��t�{�]��4qδY����;DW�l�7��$-���k׺Wo���n�H������[�{��Q�GR�v��w�+t���O[=�ɄꙌ�EUy���Vs�4v�z�[Cf��%R^K��^*�:=��1�C��Nf��b���U_��� �����}r�l��y{�Z���d1r�\����"U����q��u�ߞ#��$E�3����%�^�2V��-yX#�����L/�qu8��ۇ*�<��2�,���eq�u���L[A���N�B����x\��}�o�_g����%�g��BѶۄJ4_m�* ʤSim��#8��Þ�h�79^��AcR\���
U���y�z\x��n��Ce�f�mK9Vxf���j���.�]����{�a��y��}4Si`��E�;���{C�N55И��
�\����?rLC=�~�g�s���G:C�����x�:i_�b���L��ƘK�l�+5M��{�E�״2�9�2g�vj>���`�:s��%�8�^������&Y��a0���(����8S=�򠮕�ۓ��U���fK4M}Η#eq��!���Aة}�y6����lOs��H��Xѫ.u��=��u���v�z�I�)rV*��g�"����Ǧ�'P�u�d�y����5J���{�>�l�\��VԴ(��*b�x,7���:G��u��{G�ɋ���(�C��K��^0�ܲ�[<�S>ࡖ��P��X��i!CY�J��p0��t;8���y�;=;m�)��W��Vk�3��SD�j-CؗvD9��4'��3����2=������˸�g\��x��f�%f��{���Y`ۂ����;U�7�k�Xu��>^��/1��u��ޤa���yL�̗�xk��3zX�>��_�s>/���w�ڃ9��_����z������;L�ayF�뺱�̓�I�*�ʴ4�='f��j��EnW�{�o9,��K�=Qgι��Z��O����6�+��{v��\q�����;/��z�V�ܨ��_]�ARyeN��ʲ�k��g�~��T����Rtp���t޻؄�APs�!�	fz.c~���(�:���)�[�_�x����W�z�����p�+���C��x:P�����+�q�u1>#��2��[�=��{*o�0�x{��&^��$�#s��(z9}�b��rӀo�idH����Be��Wy.u�(D#-��s�w��s0��a����LL�˞�3��/;9����F�L�8����>C�}C�V��}�2���U9C�',x����{�\�cڋ������w��˾1W�%��(q�AC��J����<%�NP�+��*-u�1���'�\qZ{L��o3�0
�L�˩r6
�"�U\f]Qb��W�<\SW�Q�K��&˩�[��q�����rq{��F�4;D�\���W
	�c�/ ��a[�G�rb�L�+5�o��På��7���z׾jrDIT��M-��e�L̕ݚR�Nݮ���S�h�-�f����v��j�ܸ�e�x����@�:�}�6:�o+|ue*\�^�y���5���f��h�+c�	J����*
>��E�M��é\��������VtX����P�Y���j��]؟4��r����<� �a+���^�����aklS���F���H��P=~��c�>�v��S[�(T.�SI���s�<ڙ�=�L0֣�.ϥ�	g�&�M���~��02H��aH����9{Jf�Uj��`�c�dA�Ev�8����,csjx����rAb����_��G�y�T�\�e�oZ�0oL��*CH� �­�$2������ţ�t�Yj~��� S8l7������XρV�]	S|k��3ƫy�߲��𠠒�§ӌ��OF�]ʷ�a��6 r3�Ye{����x��f��oH�9�g���Ƿ�����},��;��a̷�*�v8O.5��kB��,k`h����v����{!��Ez��[�j���|~���?.�k�) ��3˕B��/\ɨ���2�R�>�^ՙNƬ��`�;rىԵ�B�g�]�4�AX�x���ڕr��r�t��)���՟%�Oj�Ԭd/�`�"�O�d8��s2�Sj�*��Ǫ	8��;ڣLï�{!�f���I�V��$�zS����;�^2�M�փ�eZ����z^�oC��:y�G��VW��Wg�]�y�en�c�6��~�8�����1{�o��:�W,NJs�P�s�ym9�s���CI�̮T��n78f<��Hя'Az�v�]:S��Ɍ�8`�G$/N�T@�����S���_�3΃�d��qL����	�@�A-Kb���\^�r쿯to�����������I���D�s�TBoV8��Ξ6Dq%��@?m��*iJ�C��q7��v�����g �O�����d��&�8&og�y��O������ ��s���y�cv܂�$h1'���
��}j���\�|ڗ�_�s��̔�c��k�w���-���qM���=e ޤI�G� �(;Z}�˝ì�� �B�]ֱE�ݹ���=��r�q��g���>�4�t��]S#�X!����v3o����3��IoTު�V��X�t��x�J6�d�',��x.�%�ґ�,��qb������Ѳ�Y't��r��M�ܵi�7�I3/��`���)y[���m%���ڏm�{�S�ҷ
�4z8x��xl9�W�!��tU�L&�:�m�L�q�>����k�=���:��0vw��W�2 ó=_n�
���Dy	�,mt�F���1=J:DW�V7X��!\/z�q�҆:�1�*a��s����xsel�4�S�����n�pP,_uNB]�9�i�:^h����\l���٫y }�퇷F�5ˮ���\7b1�sLǇ:��&�b�Jjќ��AiM.(U��E���gx(�ý�dˋwvH�fN����Zw���e����j�D�/��sƜ�녳��[U�.���үw�E*��uᙻ�h{Տ����y����\�����"L�Y:3jz�Hc:�sO*�{H�,�Z]��[ٺ�}2_�߼�}r�n���8a�ץ%c!�K��0��=p7H��^{�N���>Xt�Դ�����~P�k����Ǽ/-yX#���R���/����G��]]-�f�[��֑�1N%��.u���{BqS�L��U�J��f�{�)ߵ����pn�Nr*���8M:N^��r��Χo�w9��P,j��L�2z脼����������-�iq�H�j�˰��w�x���l�a���L��W�a��Fڡ��j�y���p�;z20z��@��R�l�!��]H;�}�.��0�w�38����{����B�q_-"��;�U}.�4�.J�S�p}t�e�v�	s�%�-#�i�V��7�7ީSק�+5x�1
8.TşK�a����<��u����uԲ��c����@�0	��o1j���e������z�Δ��N�WY��t��;Y�Ja�OY���v�5ap��Fi>���O>N�:�l���ãX�H�h�� :j)a��U.��nbKX)XV�MY��z"�k�?��3�xu;����v���K��}J2/r�yl��Wl�	k��r��#�IejB��w�0H[Y��{��U3�]���W���{eцZ���U��R� xx^W�b�6��޷P^���kVO��w�2-��a~ͿE����炕��՜+,
z���m�,GT,P.�s�es���|;)biQ^u2����u��iν'�|�S��`J���ΐ�i�a{FbZ��Nk;�obT=�3�����JT�n�k�)�ͻ�xf���RV�t���Z��ݖ��A�E��G�,�Ҽ�$&/���Be�G��Һ\�z}q�Y�~jB��8�o�toVFw��#�e�z��ITG�����>[=[�Y�No�id^��d��r�%9p�w��+�Q���c%Y�s�L�`���s0�Xz�Gs��	����z��S����w�98����Q��)m�au��*�p�4�Y��)��	r����8F੗)�_Vz��{������T�����m<�"�a3�����<%��w�T�U�Z�m���D�p�c���Nk��`�Ռ�z10*���t'-.�}Z�-n�K_b�P���]wꕝ�|r���j�@����yS��e �k��m�̇%�i��ڞbː�rwX�a\9.�Ζ�,(��c�7�j��Ԟ�2=咇�HEL��;����Y{�����5~�ݙ���a�o�Թ+�貪�̺�:�S��qMG��۸��j�zD��7��"潰Pd=�lv	v�Zt�qqe̱��k,�\��ySh���;�jy�� ��_�9�M�%�^�胵9"&˴rh�UzZp��l�wc��U�厯 ��%j[y.�yo˷�w��kya�x���|�o|g��Y�w�:{'��g�uj�zcc��I����biC�cw\�����fx��U1i�C|�2�۳[�v6M�dw<=8d��M��0G<���q��.�.���7u��oS�����tKK:p������Jc��<w���>��h�;5�S�Pײ��=�Q����$ �a�'����0��nռ�}��5�@s�}�-\�NX�L:�)E�k�f}R��7!K=�x^���z���gJh;��IA�
ܰ�qc^K�:��=�GX�v���ECYW�VC@V{8���2�|`����U�xu�Y5�w	"�s-�^��Ξx+�ה>�[C4k=�yC3DWG�r،�G�9�Z)Ջ2T�<@��;W�I4/ U`��Y���3Z��Ws�RtŴ>U��GxB	D��<��"�vX̸�E���Tq��	����6.!Ajؔ��F6uXj�u%jb�|87��ƽ؅�-�����,U�����ݏN^`�_{�臼�t�=~�k�}��A!����d֯��X�Z2�"���`��A����w1i�P�QU�\�q�|ǻ{ʞ�a�zF�2��|��Ƭ�W�LP�V2
�0}�E��!�r�v[���u]�k��ze^ޘu�^�u�	�l�0�u��=>K�Z<����� :�(�+_��C�a޽��ż'p��W�s�@�?.�i�k�/D"@�N�薪-�J�����n�2�U�^l�A�g�
�䏘Bb�:%��;°J�x�q��<l<
��A&��G���̹٣�~�7�_
ֹ���v�ʔ��'.�?mߴ��yf�\*�쩣~�.M��$��˲��fpa����-�g�(s����8+�y*6���?zϥ���&��j�v���=�E��b� Y�v&�R$�_XB����4�q�X;�^�~����h�V�Z�u���x1��v.�w��^�aH��.J�J���ñ�}]^\�.�van�ט�%&4�d�{Mx�;6�%xu��g�p�n�[Us���v���@t���c�&���A�̫�|���l�J2%Bd�qrc���Eݣv����:�:o��Cg�ķ,9�7Ed�0�S����yspe������;�L��+���4�4Ibr�x.Ԓ��JG��\E$���|���3_Ot�2�ܽ��h�l�����_v�q0�������ICl'��߽�=�xX���:G�¹���7�S.��u��>�7����'ʽ�pS$���>�=x+�ޕgo���uO�8Z��)�&�ͪ���
k-e�E�>�s���%j��%�n�V�����N"��6R�n�}�^)*�3�z�!�T���ǀܱ�ap-9����=E|Cꐷ��@�t[��m`Ѿ:ʹmO�U�.K���1/����@���q!�-?k����J��6&ZNy�=�_���tj�u2��q&��tMN�՞����xMۧ�V�3��$�ۦfS��)�1q=^��ǽyk���)���PJc����ī2����d��^���m#��T�g��,';G�J~�yC��ra[s�5ߚL����鄴���]t�G�����J��C7e�Ka��c7U�
������4�+���q#�Z��K�d��ˋ�B�t�u���U�N����=$�݌S1Nmq���w[I���5��}��Fk-t�l+۬���A��	����^)"�9�wl�w�]
w1bt�g]ZhMҟp�WwW����&XN�f����4���Ui�m+�|6�d� �{��;Cr�G���q�ap{������O�ƏmZ�h2�k����:Bր@�θܫ�u���ba��M�)�.�<�R�}x�q�S��8-D;h�w��Z6��i�:��Yn������;w��E��ް��Z�ҵ�"�l�/p���8�F���"�1�]W�����_0���Ѥ������Ik���0a�O�6���>h6��Q�qW\W^;%�ݦ����D�3�����<ݳ�BpZ��m��U��N5���5`��H����cy؆�,_ �*�E�[��IԎ���=�˃�]Z�FE�7w[�u���a�,�U��#�k}�ax!5��6\R�ܫ���tt-�!2�v������k��]P񉸡�f����+���[�,�n0-��;j��n;�2E���]� B�g�D�7JAQ� =G���8�0�K�������hU���J�0֥�K��V^��N&��rƢ2����u;�-<Z�t9m:���b5�][�(��Coi��Y7M�\�|tܫo!
I�n��y�l�� ov7� �0��`4�Q�uZ]���m�vyq|A.�=����<ٳQ��u�1�]@8'5GZ��>�ԏ]�v�r������}�L�gm��6$�auu:d{}�r��9=���9���҈�/3{�&AhQX�V�nu_<��V��f,�ݷ+i��]�� ښ6(�Uω:�eh}7��l5��)NW���l�'p�KCc#�┣�'v-�ܵZRV�]��ne�׍��;L�.�W&-9JLv�Uu�@��1L�:�.t����7�P#.�"�̍#V@�S����8GB{��g�jfK�����ri�ŗ�*��*"�ڡn�_���k��߳mvD6skj���WTɹ@�����n���� SF1[m���R9p�7B���@�``d"�����vlt�9�"�d/����k�g>�˰+��� ��zn��Ծ�R87�q�N���V������������/����BJ.�;9�yW�'V�l�v���t!34��L>�Љ��rmm�U�wH�e(�F��.Қ�g��?X��I�|o�=ɚ��\�y�#�eъ.ǵh�˴ƪ�nc�ց��o�VӮ�GKNMc�2�����q8��X�i��1s�4��:�`#V�kU��6�k��AӰ�cβkQ�ڴ�PT.t�P���y �6У���<$�w���%WTxI��:��L�br�v�1��|���/}ߞa���}YQ�ѭ*�1�b�F�TQ�,b��EQR"��X��D�QTD����"*�UV-�+
+keFYQm�UQb�J�T[h�������Z���qE� *ZX��U�X��e���e����F*�QPX�E���
�"�2ة�ADX�)b�%J�EeB���-�J� �Qr�h�Uڈ��E������TUm�c&Z�QQV,r�m�Q�+AE�1%�jQPV�ȕ*�ŵaU�,b�AEDkL��UQEUR#e ���Z"��"�Kj[�"�W[m�(�J�RҰDAETV+*��TEjQ����E@dDED-�QR�*ҌU�6)Yb��Z�U�++(�[
�4RѢ�R���iG3F"
��Tb��j*�F1*��e���iAJ�*����Um�0QV
�����"J�*ڣ"��J�_?W�f��Q�I_<�7�%�>�6�d����C���9h�A<)�
毴�נ
L�̹x����9[�Wvw-n�Q��]���\�K�vDsWr�v
w�_�,���&9��S�����1�N�֖�ƧՙX�	B�pK4M �.D0� �au �=�Bgp�(a��j�D�z'�/s���k^���^*��0v'<��NR�f5�PL����y9��d�u-c�<��$�^z��_>ǞZ��}=��FT�(�R��/��?Z��<�Ө]�.�ݥ�ci�������fȯ��%����9������5v��P����B.U�����p�[G��FǨx���mϛѮ���U�;��懧���w������C�&��+��w5sv��k����i�?Cl1]�巷l�c���f�3y�;�=ŏ:���k�rh6��u��i_3lV4����O�	�C^z��uH���t����7��4綠�Vއ@�;3uh�~xj5*�Ϸ 8�ugL'M��죇��u6��,��������EЦ��yCݒk�Z���-�7�Ɨ�Ƶ.2��ֆ}Yk�~��\�z����#�gZcq2�ܥZ3{�� /�k{5d���;�����p��yF��l�/0��wr�ber�P�c&D�I8�2[ �z�L�$LX���feV���v�+R�ک��Zhv���:�����S��q]�ɣT������fGV��e�菀�2J�=���(z9}��V�ȳ���o�idJ���Cw��hu�޼�~΢6�5B������Ln[39�w�,=C��ݧ=P�{
�ù��[��������'���!˅U��9�i��l3,S��',x�vy7��מ�*��۝<g���(��Ssڧ����]����ZfUm��Q��c�����Sx�&�a�U�E�W\gn���l~X�;��&����*U?]��t�\�t��:=�Z=B��O���*�|��O>��x�W4y@2>�!��g���M�lvK��ӤxX+�x��~�7	)����_��tΏ8�U�X	���!�'?i�d�kּ>�;V'R"J�|94��bP��Dr7k�$���-g�
�v2�N��#N'Yܪ\�>9���h�3^�k�gWy{��_��7���O��Į��yB��Q(q��Z�t�L�eK^<"���9[��F���ͽ���ܷ~.	w � ��r8�G�:�u�_ׁpM�\��s+"!����Q��͹���_�U�]��4&l��/q�pޝ����2˩� E�|����`Q�������D)vi�:[J���n`���X|{��؀
�f��H���;2��7���M�Vֻ�.��̽��j���Rm
,1���O��S�,��O����=���@ث<0&a�Wva��H�GZE��\-3����~֢ʸk��_��`o���E�$M�
J}Ҹ��&c�ZтKGMŖ��h���@Tp�m;r:̔��.�^�ǻ9>�Z���`t6���+భ�W�Խҏ+�g�(��/)���1�=d��I`������=Rz�m^jǊ}���u>�MX�I�zW��僧�
�ϼ}^�v��'��>I���z�i�s��]c�ⸯ�=JE����Ǉe�y�l��8�����ģw��3f�^=9=�nz�ܹT�o�<5Ա��a�W�l<v(6���b����=1V��t� P���J}2��G��q�>KԦ�C�_� �__P`�΢�^�J,�u�Ë�F�|����w��>
;z��Pîe�=¬�����\u%����S����S33�8z���-$��D��\�B)���)kY�g�3	���>�L��]�JC/�F<�b��3�E��cg�sHߘ���Ήv1��P���Ӎo,<l<TGVX&[]�X���mv�SOZS��W�c*�P��m���o��ww�r�v��,��۩��(������ȧ��7��=����:��P�����f��SoH���������5��U��0Yv,�:�]*��p�^����C�u�{N�j��^�낓������Ӹ��CG�T#��e�2m��7��<�u�3��C�+&*n<�^�vZ�On����#Aϒ�}B�;��L�uO,	ˇ^�����m�!ꗬ�0�5���y&�u��f	���t�4Gօ��A�W�hN�[�؂$/���z�)�Y��Z���1v{&C�%�f�D�.���Ԭ�v��l?l4��/Wۊ%��!�S��z�!ֳ�S&����(�тK���RJ�R=�+���wE_�X���x��L��j���6S���衅�T��(��l	)y[���m#�;����Wc}ө_׺|��}m�/��eC�ڦ,���W�t#D� e{��6��g�������϶�e��-T5+��Zkt�V���R8���踫}p7�"eq�e�ճ�wS�f������JBm�u���x���זo�:/v��8��T����eI��@t�-U6�x#C-���������^�-:�mi�^U%�	uS���o�-a��u����Tt�c�	<5?WJo���)upƳ���*�ys!��z1�hWg=�eV��9�n�)e����+����,�3�{.�[$�q��D	�x���X��Gb}���0��[���Z�v݊!�$,�\��r"��������IN]G�7[^����3�I��p�-�|{�yiӪ� mh�gЦ*G����s��u�hM���d�ۦfN^	��P�y?����q�,V�\u�4I�5.����9���]u�W�S��Ď�*D�z\!�� jw�A8��^��(vyGmm''/gw�a���E�C��GRwJ����M+�T3|6a3%0�Nv3�)��έ��毟,Si���z�x�,��q������\��S�J��g��n�e]�>�ZUyk��#���
Xv�<�$�Ξ�Y�Q.%��+�6�Y��}�p�5]?�W��a�x��E���{�n/��ɘ;9��ϥ����X�f5�PL�g���=2�s�����x8�F(g�1Sפ>�~]��!G.TŒ�Xx�C�#�M�3�vw���o�j�
�ۗp��Z���pA�7�R��m�o�_�U�v�~P��b��{W�hJ=��w=���0<Iey.,�Awy^�w�K�����-3���%����A{}[�Va��{V=~��8dt��7�X*J��h+O�@m�v��S5����
ae`Rv���Y�ʾ��Gp�ӝh�)F��[K�
���۷�#������Y�bʦd�����VSw���9��&y @��*��]LC�-J�Ŕۏ'�gź�#����H�^��f^��t�K�\�X6��p��2�(�,��F���[�f���Y�����<F�	�C^u�m���W󋃩<��-�y{����Z�I�7�J7�������'�	�{=�G��6��S9�e2¯1eYt�/;��gYׇg��l�/q��Lg}����ӌ�b�5<��B}Yk���%�-)����sk�w�d�㚫���2#���3�.�����(z9}��=[�"�Zk�E{�-�;&���Gi^���2�]��)�."�2<��^Ϋ,��K�m�3��3�t��������y~Z��H��uL�K~�8����Km
P�gղ�8i�ZͰ̿���xۦ����y˃�N��1�sWh��w]����ZfUm��$ǔTK��P��Lfd*�8�SsK���l�<霕/��Ӎn}��g��GQ�:=�)%�Ѥ+j��̤6{��7��wm0�����c#죀���{��"�a��.�+N���}
>>�=�d��X��o^J�u�l������S��Ū;�!c޾5�
���b����Fް�ɂ-�O#\z�eʺԌ)J�񷪺�KV��"��1Ho�����D�^3*n���P��Ռup��<SW���jG���=_ Cws�g�X��t]5�Ǟ�d۲�U�-t�6�æd��Z.^���|Ж��Ԉ�.�;�Y�S��r��1ԐZ	%��Xv
˱�Җ{z����&u�j�.&Y\���s;9��;�\�^�O��Aa�J�t]�P�z�P���g��~S1\U�<C�o��ث�%�O(L�1vt��ɗ�s�a,��	!t��\]uA���4��K�^���
0�Z��1F!l)��Yٖ�O�����<1Cؗ��������xg���w1���M1�Ks���M���-��$�V�3."ׇ��t؋-C�����H������w���x��=Z��lU�h���5y��5�s�^s�4Xn:�V�G�C��1V�Gks_�S�i�̿Wbf��mC�>�Mc�I.��Ao-H7Ka�1���q����k��f�tǕ)g��}��iǪq?9�gNyǈ�n�u��>�u閜;N�?(J��9��q����=�V5�R�,�����>���f]��}S�-S�����9��}�j@�N�s*b�P}�嵚1[Y�o}��er�r��V���ek֯%����ت����)@Jp���5�cVR�u�����뵶�)�ܜ�ne�bsP38r5���w:r�Q�}�j*��S�,�_k�v �N*�(f��X7�%��^}��j�u�b?V��՟%�Q(|���_P`��������3�s��+KH�S�s2.��C>�=��Tj��V�Ui��UW���ߕڔ��w��xwlދ ��6�:1	:��rޯ}8�:׾��	�U�%�lH���}}=;��b�g�ԫOg���ʨ�6<��Ήw�w�`�':���o.�h=��Υ/}��S'eyu� i�Ė��N��*��];L�OȹP��ə6���3{<r��*��&�/l=�����jI룸:�(F�IsQ9�u&X���ˇ^����ɲY���t��s�Iv߫�� W�l�}+Ęl	���'_XB������KhR�n���jľU��rg����ޟ/ڄ�T/�$�����fU��z�!o��I�Z��ᏧR�DZ�M�t������n��l�ĦW[�?g��r�8�Z0Ibr�x.���}ґ�&���]�m��w��u�
�EAT̵g�sij�����v���<�0!��Dף�a�⮗V���%�:�l�i�.��T�a5��}���R��w(u*ɯ��[��j��dY+�^���x	=9�(%��u�!\Y����(�=�4\(�u������dӶb1��]9�U*:G[�,V=�;pX=�:�V�.b8�,\ ~�Ph��۶hW�GyK\7��O��Z�F�p&I�V$zX3�w���J�m�K2;v'K�lٯM��]//˪nxӘ��q\>�;㠾���~�<k5�gۖ<��F}n����)�`�^��(�m�u�D���_���9��g�G�`y���j]�n�z7�Zlz;ig����4�踣���9f��TΥd^E��&�ܫ���4e�Ί��7[䜻�*��;��k�_3���U׀V��8��:�9���za6=�OY5r�Gθ�K�n��)��<\���Wx��_�����9|2�<�]����_����4��>���;�_�L��GG���K�5:�N�	��O]o��L�����=�i�L���֡-4��~�l����tҿ1P���&^Ka�N�++���y�̯x��{���{�wh�k�p6��$G5R�ru�pL�7�л�k�{uj�?�>�;(��+{���Ξ�Y�,�4�.F��������,o^�t����B~��5����ziǠ`�,�nm";,@>F��;��ܨ�\j[7��zoϟi{7�['��T^z׎]�v����SG,] w]Z�T�co��P�Ϊ|��˝�2��몯08��y�vnh��ͮ��������$��w;�1hH"���sQ�>�FUKk\�pK�)rWT�h<,�چ�{ߕ�~�����!�C|1�`N���L�/�f�d��Q�.TşK�a�~��K�Ԡ�}�Ln�k�(Z#I:lcKz�Px��f�hήWl�BR�{�דa�T�w���_���>�|,l~�����+���]����0�^��K�hxy����~��X��ow��ff��Kcq����U��
����h��q��c�ӂ����x�;}�����^{<e�e�u}�S԰��1Y�G��Q�U�I��+�'����y��צ{U1�Z��ӂgw�>�����%�\�9��8w�Y�؅1Lu�j۠xK9�y?|2�v[/znte�0������Pu�[�,ny�iz,kR���ʶC��ca�8 1{�Q����Od;��%u2�{/����p{/L��v^��IvF��P�G1����C[��ލ���J�X^�K�f�p�ya�[J�O�qa2<�]ȬgU���crٙNf�0��}�J�瘱�p����0�|���G]oS�{���"���z��s'�;z�ߎe<q�t�>wwO���yz|���̻�� )�M�P��m�S8)R�kUр2�%1�!��hSP37����Z��B>wp̮PK��:qa���[�V�X�1�Z��J<J�ĥ���������#���I��}Ǌ�V�H��wxe�8�f�YJM]�X�[*���͑5�^\���s�X2�H�fB���ۏ��=�u��kin�͡6J�/��o+�X��c��VB�uܢK'1 �ɚJ2!C{�{��``n�c�zn��.��*l�[�1�Qr]B�E��	�O&��[[���YOX'��"'�v�ى@�:^�+��r�5CcpZ[.��mU�ne	��t��x���C-"�dL8�C4n��z�ȯ>���E�\�I�wR��i�t����W/��y�l���sI�#z�T�԰ee"9�y�HcX]�E:xe�[�;�u{ԙG]�����8���	Wr:��K�VP��Jq��\��������#�q�1��
L��&e�P��i���s�J��;2)������<�&�/n�Œfn�-pq�> �YPM�Q{-�
�'�K&Q[��!(��v�D�]�"X��Y����W+y�hz�N>�I(ν3^���z�l�q��"Gh5�3�%��/��D��9`�oR��LE���O
4d�շt^�����.���ڇn�H]V��(��O[��*��gQ�����U�Vh61���v�k[̎a�2:��(p��j���%���H��ZSr�%�l�g��st��9�j��Իm�9��h��*+u�9\��3��jK�Զ��(fN�Zi5b���m.l�.�k�t���_h[0�@yէ�������Ʈ>wW�jʹ��O��\�}Y��Z�u���[j����y�VSǺ�J���Ywϫ+�˱lud��En�q���J�v�	D굵܍��Ʈћ���j��YB=N�e=���#ŀ�����bY�����v��{/�-�a�QǑ��k��t��-��`6�{w�4��ov��S�T'T|����x���@���F�T�>y��4gfJ����+��e�Y���o
���&�q�Ħ���r��2�=��5�s�+����l�i��t���mMz�#�2���:����8aJ=ʳg8���[��<n�����I=�Z3� �u���������I��<�'@������
7���Ұ8�.�F��iwC1AΡ�vE�}��6��|��*�9mu(ѻ�|�<%�����W�dk��g���Q�J��0�E���s�.��ٜ����}�ʬ����w�TdJR��rU�=x�[i':+on���]t
�j��� �8Vk����L.�r��v�!�8͋�t�������ݭQ��R�-V6�j�Sv��Q��lb(��X�T��TA��mb�ciee��$cTV,R�(����6���`�1��**,AEV̪������T+e(�Qij0EF��"�*����iJ���Z�Db�*̥r����R���cL�EP�*+Z�"�*QUQVTR�R�R�V"\�*�`�2�X��feAƪ
1V(Ŋ+m�X��[lUSV1UfR�5��#Dc���3-s��1A�Z�Z�
j����jUTAPm�
�AW(�#m��S��#[1%�PUJт%��V��2��E��pʒ�rʋZZұc�2���G2�#�J�m\��E�,e�fbQck�[JŊ�A[J�.eDQq(�W�T�iVcL0Eq�յeLCm�R�e����r�h�ۘ#�
4r�fZ��Z��E�nLf8e
�*73��QE�V�r�1V�bbb�"+R֦4s(V8�J�fT�2�kD�֪6Յ���Q"9Ki�Aq3*7Hҥ�j��>��u��F���R|�LBn\4�p3�p?l��\�}���V�҃xhD�@��7/M�m�)J�w�j)���]��P��Gk�vf>�����=�:pN5z�R�B�N�+��Vˀ�i�Z��~�}�6�u�R׃�qx\%�����sy�����`�h-5�g�[i�C�L!�LĤ���Y�ϧ뾎x�g(���s�u/���Cۀl��eYL��\���Ȓ\d템���Yɡa}�w�����}c~��jj،L���5킃!��c�R�:G������ًUA$�oM�o���AAx��vfU�-s�6�t�9�s�x�7�\���+۞Qj��7ٜ i�5�6���(S2�R���s]�.x�����4OI�ٵB!c���zk'�-�4@��kR�K��)���q��Y�X��3<{���m{�*��3�V�O��f5��ׅ��8A k9��x��v�xi��U�/��K>�۵n*1N�V+tE.s-�u��5]� pU�����a��=4�du�Y�u�Zg��1Oqv#��Ϯm���O��5��0RV�EXs1���-h�-7Z��yND��S�ߘI�Rz���hp�v4����ȧ]B.�v:��I�5!������]Dq��H�%�䫫m�۶�ܧ\:�Wk ��_Z�6�?�H0��ܜ�R���NE7�٢���;�ʾ}��S�J�*U�^'}��	$��'�Z���u�Z�a�5a��2!�L�eR^�(.t8�5�{�[2���*Em���w�W6�V���g�K(p�v����j�t�a5~w	"ÙoJ�^x�Y�e j�f��V<�5��+r�&X9�}R����V��nbc�v<+��59 �n1�]��8-�</���S��3˕K�ݼ���Y�,j���;$�{�{V��>x՞��p������/N��{|pw��JmT:�@��+�u���%�e�܇{4`3��<�&C�Իd��e�}��=��ʳxo����Zm�D�K<:m�{9��q�/�M��9Ș��:1X���&-�S>��^�L��2�;Ʒ���Λ%���v�[V^
U�r���4��A�Ɖo�
�Bs��{S����Fu���=�|���S����d$����|�ԻL��-	˄{e.z���ƣ�����+�·��V+�r	BZ�޺=�ݠEF�A.j �=��Lன��ï;���Yق]��s�Wؒ|���]�]��U��'������sB���B�V�E�	V��נ*@u=R'�e9��OR���˻Θ:c����o��Z���l���V����w��.oh]w;���y���ܡ�+�\������ļ���t�:6�{�{���"t��Y���垞�s%x��4Ms�I���(8�g���F��=��E*�>�'Ri���Ql�u�R��?�_��Z���^�'�#�.I&GR�1�gF|^��|�3a�߸��ؗ�K���A�D�L�5C�(�џIbrϥ�s��Iosס]Q�!���ʸF�򵢓KF�,u�1�0^jD�B�O��`�H�7������;8�e������1��6�L�	�(����5j��Ͼ=�bϷ��VL&�&cD�.z����w'�K��zB��l?d������+m�5��Z��yt��1S�*�|7��a�k����St��v�=Q�f��s݂���Y����3-<9TϦ^D/6�3��ٰ�����ø�}W��<����~r�Y������:��-�C�e��p�T�N���o#�5vK}��[ڳ�`粴�3�Nf�ҡiO:�us�_�Zn��kީQxf;��W��ӹ\Hnk�����9��񄝤�NU�r�
��޿=#�K�5��o<ҿ�B�a��j�s��d���v�I�@Zà^:+��&�pֲ�wz2l 9�+\`0moGs~ϳ��u��֞Zݺ�J�k���ޭ�^Rk
�@���7�u�

��mV�9�m�+���7)l�rD��YW��s�T����\��^��W_���q#�y��,��E�S�O ]G�1��;�;ِ�en�e�3��P��ଵ�XZh3�$�J�ʨ�~b���Ƀ�zg��Hf�;a�;�w1���[n�T$��U�u�[2���ݢ����O�#��r�vS�JC�Ǯn]�UC[�T��7���d�reoz�$���؋2�'�R�A��C�o;�����r�J{����N�[O��i����盋�*��\�؜�P�H�jQ�7.��#t������N�|2�ԁ�%�ָ��-C<銞�8_J�^*bj)k~������Xt�ͧ��Xz��L�|���ixnZ�9U<z�	T7�鋣�ž;��IYD��=+��u�S���Q���$�h:M���7ᮭL<%�;+=���LP�ʦ�U�r�6�dػ���i�b&>9�>�.�^��¶�G���|<�w�y�EO
H��=�z5[|�~�K����e��=K>���}5�Cm�f$�����Չ��[{&e$��T>o;�Ţ>KM��r=k];��˛�^�ZD���N�(�3�-��OnLe��X����Y]�mqO-:�>�����"͎��k:z�h�Eo8��.GFɣ��'B)n�����J��S{,��+����T�N����p|�=]2G��c�ϵ�aX���"�ά�鿶{���a|��Gv��񥚼�f�@��eq�۾3�f���^#�Acpy���ظ@_�w����Ԧ�~f��{:����n�o�~�ӥ��J��ڶ�e�}�zfIvF��P�r�T����+v)Rw.�CjPz��J�p��Y�yx]ȯ:��|t��r٘)�ù�;}ì���ޝ0k|�ݎ����ً��^��!c=�<1f�'C������)��%�b��r�J�x�k{��7>�~i�	Rǌާ�O\;����kMi�m'��qLP�
w��7�eU��}�%>yGV�݄�`59C�ԾkӍl��YXWR�l�E3�h|���u
���w��Vr�#����<dSW�Q�#�[�&�a�cf*�%z9i���y1�=7уd�< +�υ˱�켪�Z�njχ�?����[�C�5���(�H/ӡ��<X\�h��љ���1 tl.�^
̱�җ�W�k��.�N��9�[�ށ2���!4��<^�ӌ���ʻ\���^]sy�BW�V���f��N���TF�i�6CxPn����v��+�����/�tr9������oR�^��0��&����c�_�U���org(rV�1�W�^�Ԟ��AlV��A��P˽C�!���n�j�طd�:.g�:�םyQ.��$y�A3��Pϱ��X9��t�+49��~Z\�WN��=��B�5�92�ܗ�%���$!���b��\�봻���8[K���;��v��/A�0Q� �Ev�y�Vx`P÷���xu�FP�[G�y���yݥ��eg<����^>�����i��邒��EXs1��-xt���e�^%�mf��y1��cy*v1^H�>6w�.���^�6�9���J��a[�6�5�xt���SnǪ�0r��T����v�C�֍����<i������</���4y�>�M_��H�̆���×�����eA%o.x�W}���0��E�Z���h��U�8:��fh[�Y��yx�"���W��x�^9I	����R�6�ً�9�6��]f���/�F�|��䞃�b<�{;����bk�F�闧uz=�=�Qͪ���P�Zqo�3���K�t-�>yCA��G�YL�����t���E:�+�<+'Ԙp=�Y��(m���v�w��t�ƞ"�j�.�-�r1�\�9KGl�jȼ.I�C+T�[ʈ��2�j+�����,��v2��i&,�VBt$q9��XИ�Y��e�f�NC\}q��ly��5�,����B���:�W��F�V���L�twf�S�C��RK�����SP��F.N�0-��i�k�E�/�m�Ǟ�XB7�x�zW��q:��H��>K�Hu}J�̯����X�9׈����~�\�yM�k�ت�*<�86@o#��K����?,	˄{�l�d��9^���Cݯ�s#�=�+�{ݦ��Fs-��m+���i.j`�C�WRg~����^�Pu�#�߅�^�-�������X���^�>�.�o��V �u�
��  8��(8���}7��������>R\:�K������L]~ɐ�b��'�#])r@�#��>�|H�x��;U�tF҄B����m�u{�B� ����aq^K��὜�����Ǜ���� w\�0�s�$9{>/6��:=�t�����2��$`0osLi�k���J�m7kRjG���$^�����b���(��j=�Q��tU��	�'f����|{τy��/�Ä�< �$O}޷)J�f�t�ie��x^]7<i�T�Ϯ+���+]~�Y�Y][[�(W@dg���؋��lv��a9S�@gof\�ݶ��'sVOUȘ�K5}1��ݛwن<��+�����R�
�w\��ל����3��L�}�ͣ��#-n����I�0)�Ym�OL�(ɱ�g|��^*}��7��#��OR��B�2R�l[��&'�%��-����*k=~��g�#;��<ge<\=�卋�i�9m/L�we,t�(���]�5[��WL�gL�pz���z�A;��)�o6���!�v9��3�	P��O;��h~���S�Mvl��V˦n�ͩ�b�,�Z6T�`.sS��*���i3T9�w�B]��Y�����>]8bh����-�^z��=.$q����N�+4{W�9��T\�x�:�|�fz���S]	�wՖ��|IإCf]�x��M+�Хߠ�͗1e<�a�M@��
N�}8׹`=h�E�\k�'�d��p�v9}�>��oӮ���e$�����f�8L�\���ԴlθF�� 8"��C�(�cݛݽ��x0�D�ڮ�勪4�oÖ�n{�n/d�FV}sb�<��H_m�x�z�]e����6�)T���A2*�Ж�������T����Vj��*br�L@��\i@�oه�ע�ø�9�N�g_j�±�6�t6�w�TW.��eg|�o�b��ee�xF�Z�~��
��s�*�l�~�^�s���!�5ض�Gv�<�dGuαB�p��t�qL�:�ͭ�,޵��H
s.7���kg�9�ٺz�^�����%-�=�:R�
�T��mgg��^�V�T��8+x�'�ѝ��bUu��.u�y���ף�ؘ2�q�P��d�Y�i/��G�^��oQا��ta�3F�츕�M�ݪ;>U�N��"a��%ݑ�hK��w���8�|<-�5�e�}�t�����v�}�F��'���i�a�OR�9��̡�|D5�m�H���s���x�x�;�w��P\��ڀ}갯�c"�ά�齞죀�]�y���}�2�o$�!��螫f�%���{��δ��>���ƖJ�\��5>%'�p��ٜq��Cp��+�l��>��8��R�a,O.�w#�Z�$�#py�e�+���y��ʵ޾��^t[�{�,p����>��v�]Y_7�SSBU��fG��Xr��n�jy������7�MC=���=P���QӟN5z������U��;�xuz�deS�%����g4ڀ;z����K8޷��O\;�v��i�V�x)P�<6�M�=][�/b�v���ْ�޵�NN�ھ?2b#�;6��pe�S��� ���+�G�2���<W&߽�tr���q�/GzQ����f�&4Զsrr{�QfikiE�YI�F��He�׬��=�
���z˲��fS�"M�����K}��~@��4�{:�o��o�p�_�Qj,��Y��(qԾjqC=ӽ�Y���L��L\\��gi{��Rt�͔e�U�ຢ%�U8���<�����|�����a�{0��Un�=�z���O{ً�;M��
�"�(&e��촇Z����æd�7�O_5�WE�q��I�]T���m"���49D�ɗ�
̼���2��\��v�N�� },�}�4����zH+��P�y��g��]jH�]�)��2�P�7u�t�Ue�����s�@ڡ�]�"��O���e�>��K,$�}����4��@7�=
ݙ{�v���|]�ͪk5�u�ht]�^��Vxb��/3>M#@Gb����"��޾Oj��k����pnf�f��IXr�nf0\E����b,���yf�hK��ΟO��yz 葆�0�^�υ߯{�(m�w�R]�
ܰ��+�j]�|�}��C[�n7W��ɧ�q���"�l�V�/��r��~R�:�o<����a5>�{GkӀ���i�AZ��L��'%��4%+I=�d
5���wO�Ez�+=X���i���ƹj<��#�,�( 4�b�}'hx�O��k�-B�Eպ�j�k��^�}���7]h���ʍϏs^!>*}���_t�f�ҷ���>w�:Nd�;&iG���1��5���<��z'ض_�z��]eإ����٣���|-X�5;��{����#�nw���j�-��X����˹ڥ�w\қ��)Ց���\+<�Z�.k�wln#�|o���fe;�wj�-hY#�jD,4�
����v���T��z�7�n���=�d@�VV�9�A&��%s4*n��`E��9d��:4ݬ�^d�k/�8��(�	n��Lw�.�hmgW��'h)T|7��_R���Y���ѡ��W�3(7Z�++sF.�)uZ"�cT�iE��/��Rls����`����hK�G�u2��m��$xY�]�J��H����b�Y��1��C�5|�T=ݫ�9V/�.�F�p�ϔ5����H�d�6޻�1G����5�c��+똨�}=K��V�u+AQ�S���[��+W@���V�Dն#�x�gJU�D�K �����TR,���l\�jr�����}i�s]���a�f��M>�֎������>ՍwҚN����y��7x�ut��_(G)'5�X� �_b���2�͌�݊�D0����ܹpd��f��$�^9�RCe����Xg�AF���n';Rym�V��FnqÑ��8k�P(��뛷��m"���C��AZ���f*h��уDW˹��^�G���J�J^��T�����f=�ǚx���Yf�3B�,JK4{^��q�'�mAOFu^pdluի��
����VP.T��T��i z=�\�Jև*��|�A�5�^�Z�%M��6B:h�2ef���RtN�l�vRڸ�/&4ҡPJU���Q��f�B��B������7�~�}Ԛ˗.�dw��ϸ�z�);���;euͭ8���Գ�D;7�:r7݀�p���V��W��3H�N����\�9N�IQ�y]fO��ޥg���ТM澱X��ZϮ�[jIN��j�lJ�9Gʘ:�����(���|�vև;�c��ft}B�jn���
�}�hs:T�*�V��k��aE+�١B.�s���'�:.�]�����3��Q�v����SN�ĳ*q�Z���]���@Ym���[C�'���ɼ���t9J�̙8���;��-Z���1����(n�r��=CsT�uMy�T0!@6�Ж�K��ݧ�'Df���g����;��N
*�9k>WHK?.Ѿ�9�S�4��Ƀ�E�;;�KG=��fTa\0>�f�.�u����-���t	B�Z]xe
G�]�_F�,qLv��~@��n�Tn;����w�EL���\Гs�Lw�8��9s�]ű�P�@V(���D�E8!Y��B���U�hT�E
���Tʴ�\�j�qFVc��j�T1\�e*媍I�a���-d�j,AUlX�1DE�!�E��VEUL�VW2ʅd�-�j�Z�11���-̈".%R�*-i[���ň�Q,(��b�Uƭ�e�sD+bRص���R�TEƌPDq�#lc�T[Jc#l����U[h��������-)j�.a�-��m���\�3*�e��jܱ�ܶ�p�D�l1.R�,A�-,��ffb�"e��,*bbE��!Z�b��Klrʕ�EV+R���˙�e�"-�����"5����(W-��31(�����Z)�X�k%EE��Z!�*���V
��`���ŨTm��ڋ��nZG(X��jP�nd�Q�q(,DYmEU���R�J��)��`�(�AX�&Z(����eQ��Qd�,*��%�.�~���ך������2�{�R�yWWs��+&�<7��=.5s<�gG��]u�APm�roh�BTƻ%u�I�γ{3W�v���t;�aT�p�Ʊ�z�u�)C��k�#Ԥ^ͫ,'N���f��:;0+�VzM�aT�;���Ï�o+�=U�J�e�C���|���{n�;ٽ�a�m1�rىԵ�5Փ]�7�/N��{|pw��^�-1����-�*]�{��B}�I�V��1E��qXw3!��t���E:���B7*���(�Bw��o��ǌe��ק�Zo�UT2��ꄛ�Key��h8��{�ƙֽo��J�,yi�K�nH<��փ�U��Z�ŕ�e�\^\�/*�H��-tK�s�+���t�uQo	�Ӗ��d���~6���`l$���'��K����xX����N�*W�4���rtNO�I�y�	��Yu�m�sf��+(Bw�υ
��֙IE^��W�O�6�Z�;� [-�z��s̳2WbǕ���K2a�y�I�G��ܣ2�"ͪ=��4�4hZ��C�)��y�>l)~���~X�L]~29/ÀOG{Ȋ�v���bt��חv(y<fa�F�R�E�]Y�!W(�v�cY�l9j���f���.l�����Mv �|�6���jtI�Τ�j�[���˾H���N ��n
�� �x�e[)5,�����S	8��`��#a��zx����q}���������j/�Z1UM��ǫU�ګ�xʥ�08j���6�IBjs�s�m�9�3X�wO�i���U��G��T�"�U3Ə����gG�޺J�P��˶�V�
�o.音?~����0�m,_�����H�:�=e�-��L���m�3��h;e��ޫ]�z_gOo ^8/���܈�޷)O�ٳ]�r\�/-��Q�������Z����6%��S�����y'�v��雂�}�>���Og�/��R�����E��Tkї��'�ݍ>����cb�\O���O[=�%�<z.(��Q�|Mն�!���۝&s��8M�'�9pLo�%\XC�c��s0o��ZW��=�C����4[&b��������=�-t��d1uiY(�_T������N�fp�������KZ�.ypk��:�p�\n���F��6+E..��||���'�Ď�*D�*��Swӝ�-�ֹ��<��9s�	�i� g�:�� t��ړR��>���t�zkqz�~�	���}6Q��n���=�:D�KG�Mޏ�0�{�K���(WSŔ���$^���ʯ�X�6����H��r�|��v��V�̂�>�>�C�l�Z�R���0��s��^�h(
���G�]�d�g��@*]���9~Ys��l?��9��,i�s��}8׸��z�uBiy���:b�Gm2_��8��sZ��F�]m+�ˋ3vY0���L��T�3���؋9,�5�r�嶺�y=y�V�Iݡ}Ays�)2�A,�A�]���m=[�L7=�7�T#+��>s��C�z�g�L����D����2,"��k�M��:�k�=zp����2T�(��G�����y������/m�kS�x,L������.^�~�P�j83����O-��m\˭;w��ë^��;i���bU����}��%t댼�������	����‷Fz
Ԃ��[kh�
b�3��'��"a�Ҫ����hK+���O��]������X���y��oo^�o����ޘ)[܍Y�-0l|৩GH�@S�p�!/����V�\�y�y7���ヷW�ŁɮEᮻޔ5.��=���>[�	w����X�3�ET�y�=vk���/F�V��v��۸g�oq@}�:�,>����N&U_���V�D}W}�6���m�̇ױQ��9@�l�z�=н�Cy�cU�KL�2�Iם�c[���� ���A>����x��oo�l`O�O�;��f����5���wy?���8��\_S�ł%�D���TR��{[mo?,���N`��S)T����+6��̛��N�����!>����U-�K��]�;�m[G�ZdE�^�%Q�uf;y��ze��Mh�[��B6�>[��o(o��}���#����+����:���>��6����n���=�;�$����uh��_Ṭ�N5z�R�@�9{��.��xW��v`�����-`����P�Ա�o[��^��6F�G��3�2�/y]v�3بw�y��zv8��@��Tu�ϼ�m��Ծk�N5��'{̳�^4����r��|��s�KR�`+�ʪ��Dw��8����1[�r�W��~���e�z�5��$\mޛ�/(t�q� Y��uC�����3'<�=�([կ�=��s�V�bx��jD9.�4>���O&^�B���Җ2���s���^*�'�o�ұ8�O[�/���7ꋉ�Wܭ��g�ĠA��J�.k�P�z�TJ�b�w�Z�ѧ���Tz{���_������b�衾GˇpK�$իIA�M@��q���~چ�[s#8J�+��r�f+���� ���u	��ox������R������-0�\��|�0����Q;4m؝m��n��#���W����ۧ�a��ތ� �r���zvk]a��e�x��h�4.���JwF�وS±��} ��JOo���~�zj�.�{��
6:VD��z��<1Cؗ��=4����o�0���r��;���]�}j����3z�V�ޘ)+T"��3."תU{�-��u�:����6y�����]��I��r�Z��FH��VU�q'/oK��k��r���g�35���J�<�s�^*7��U��0��Җh��f}4��������b�1t�j<{�PA��y��.������"�e�+��yt�b�}k�j��c�k�z��b����o���0�����^;�l��<��eym6�;�yr�k���~Y��?V{kRcNz�[�`���οvoBދ"�zw����k�~j��p��^)r�}%����
�`9C���}ؕ��
�-+�(U��Qj,�C����OJ~P�ϺOd?kDoEN�V�TN�c��7`���}؋;),����^@z��&�΢[+<��:�S�7�EL0���62j˜~({-n-gG�����47����wO����g�,pGC8�Ч��*�l�lMZ㤳���k�5Yp��2�7���.���ii�1�I���i�����DP������\�]ׂ*}��n���+�|K���q���uem�\��W*�o��+��6�N��ck`r�T��oUZ%Z���;�`��Y�hq��{�^�Z�t�C���{Wt��#�-/�-�b+GJk���Y��a�����na>���6,�c&�93{<s·Z���G�ݠ~dh8�52�~��	���@�L��{��I:�Wrf}]S�w��K���9��fJx��[9��I���h��"K]R�n�g{w���W�"�(6�c4.;�.���)~�����c�1uܸl��O���QŚ5{E��VM7���#�^J���+ �w!��3o��܃>�Kv:�ǎ9F���6Ma!ݻ�����R�7�E����^��;D�[ȍ���M.��U1�0J�뤮(au������������d�x����:^V��m%��k�E�\+>e�\+l�� m�7zj���z�oޢ��McD��d�:������!\ec@p����t�R�yl}�K,��)�8�>�Z��D5T;Ê��������Y�+�77�b�t�P�R>�mЎ���Á��^j�m؆���7,z �^;�-�鋆f��X4?��A�o{磯&�z��ٌ
kqu%�M���Ů���QV���U�g-דj�L����4�����HyK�7f�niJV�Ƿ����Z@�;.du'�g;R-�&��C�C5/�Nm�l��*V��X]��#k��,=o�YF��]Е2��}����X�M�uD5Z�W�O�ᄹ��bP����c�ϩ����J����W�wivگ.A�Ә��g[��9z�2�ϒ���'0=^����V5�'*ĳz�\wn���u��8O=]{�P������=�yk���)��jg�/�����N$q�"\���ʰ���5o��D����*=��ƞ���yC����\4V��Y�C@7�����]�}�IG�\{}�	�(i�����+5ze#�ݢ̀��a.!��3+;��ئ{������ջ\~���__��L0d�re�W��Ξ�Y�f�u��^�]�k����l�Z�+�A=au!/��Y��m=\|a��~�J�ee����3�qt��@ߞڛOS��C�.Jꙍ Yƃ�Ǧ� �K��uY�맳Pk4��髒p����!F�س�ׂ�yHiK��P��w��T'�Q�[�i�}/����T:_��o����}�&]�\�DT(OW[$��8-%��h��k��L< ��xtuk��k=�{��&�x��x�\9��Bmb�O�}�B&]�#I�u���ˢEL�|9����
�X���4�e��⽦��j�О�d�s~����]�3�K��;D%0��VU���ˡ�Y�B��$Kr^�O��e\}*���^�q��:}A{�t�/��SD�j&}��ȇ�4%�»��>[�X��^ŭf��w��֭_�f��H�l�K�s��e��=K#�t�Tad���-�t_=���Cy�V�]!��H�����9��[J��:Գ\���ȼY�������{9���ǲv/p�/�]��xAPk���>9�L�l}�w�m�(5��C�y�iz��*^O\ܮ����.z{�M(e��ν�L���|j���+��ʶ���ȋ������U%*�n㭕3
��I��(�w�@���|���Kh�)�x�(u�f@��wW^��}gm(���S��|:Xz�z;��1C��{�t��W� ���hr�{��)̭���s�Ƃ w��s���m�bu9C�Ա�o[����ê�'J��{,������2�1�~�;��e2,W
�1*΢�Y���3�<�_5�c�މu���V�y���Q�<8�N��¸Ȓ\f��#���W��⚽��Y]..k�
�ߤ8�xs{�R���6ǏQ�+V�N�S���9�V������W5|zXA�X<^>$�l�Yc��Qt�zrcl��+�\��$ѿ'+8D��XBދ*���wY �]�����0VƷ�Ҵ˜st=�$����kWq�		[�}ܼ��QL6;]�V�#��+��̼we�P�B�\�͡��4�W#-9���k�1=$Uﾨ���W��\�DK�ť��.�Z	��e4��EX�M�4&��̠�u{�u�Ӟ����ya��~��9��o<��@��jWK���3���G�:��9촯ϼ�N��$�f�5����g�{�O�P�#�L�vVY,��HC]-+�G��C�����NyA��x-�n׸m'y/~3�9{Ü�F�Jȃ���8�;`K�Yj�5�.#�۝]�%p�<���I��X-3���s���Qf邒��B*��`��^�ӫ��u[�-{m�ǘ&��F+��a��X�z̑���*׽������t��rx�ݾ���Y+ˎѫ�v/�˃i��y`CƢ�/��8];^���'�o�_�J���9�m��m���j��
���+
��8N\k5�
�z���o ����$���]�{���>�|�Ɏ��<=�����4��E����aOc�g�*��84ߕf.�k�p��57 �^w�Il�%pS�wt��_R�Kx4�8���8WP�[u�.�f�5��V=#G��J[{�@4�uwL�k�:��L�VM�&��[�2�d|6m�a�w1&�̧�p)L.�|�#kA��"�`�����xM��թ��Vm�3g���6�}HZ��_[��G��ļs��z�Mw�|&^�����~��;m0n�z�1�Q�9*��eS:��(_P`���Z�2]��Kz��rݬ��g�ު;��9�y���&�g�X������W�	9Ȗ��<��$��ŷym��9�<�/e���~:ׇ���TT���`��/>�\^�e�Ti�P~[�fz|�����V&wJ��&�s_�`t':��kygOƾI����M��Z:5��b������������~w�fA��I>ۿo����5��VW݃�X}���Qdh4�55^��ΤD{k�'K��_Zゝ?,N\:̯��9��}=-�g����^$�ba�K�.Ӛlu{z��hD�g�(o+8И�w�R��?�_�9S_�ɐ�u�q�륮��y���:�|7Ƒ�%�T��Vgk!��f�WW�:�;
�08j�!�$�3�����kΞL7C�@�Âz�U҈�2���O�k,X�1�0K�h�U�X�9l��
�l}�F��mS׋θ��B#d9n���k:VO�k���7G��Ѯ���ُTK�Ee���t�����:�D�t��z���[��\���6Pǲ�xICٝ��[;
C�LJxJ���)���@�*L���ӓv��6��7eug6����}�eM2���}Z�34��`[��v�mF����#�v�f�hA
�˺j�$�.��������f�-��7���CU�iR�#�|tuY�ޭ�	9F���̛��>8셨S�v-�E�Lm�N6s�(��f��#R���g�!7�>u���QXck�̳�
��R�̽���l*����d8���]��GZN9Z�Bk������3J��:'��Zx�v���Q���Ww!yK�/+{��%s��ʈ����,>+;E�T�Ѡ+�_Y�`�c����8�p9(�ci�%�����\��t�]��nC��j��;M�/��hPҳ�t�\o�l��w��0�B��IvS�"�Av��f��$�ٚp��N	+w�4����%v�hqlYBf@
���9x��`��f��SVfu�*��xT���n���Mf�����;�3<7J��eg4΅#�D�fu���L͓��3�l�=��Qq��^d�);�a;N��>����\��^��6�Y�lMt�U�ٚM vc�E�>�G�;#�5owz����=m�C Qe<ة,��/��N�����ejO/Ģİ֓�T+d�0"|Ⱦ9O��G��ę�b�3�o��'��2����(��e��Ĳ;3zQעơ7�|m�S+0�B�*���3y�V�<��G�{��Szy�A+��{��'w�*���{]��h����_�l7k��{z/�dT��Ōm�\:����I�-�� �a������a�tg�1�����<���١���ܛ��ŜY��xh�Er+�N�Ӫ���
��g:s��".Hd����A��.�y�;(xLtC�Uv�w��!O����,�:s��;�<�.�Fu�r�����#4����˛)Q�XF�o~"�SҞ#�E�ʶdu�R~sq�n�՗Z��5���Sm�3ݭ�CC{���Պ��7��IՐ}`ټ�ͬ�r58�Y�(�4�cU�wh��M�)�15������-�fc纇]<���2�,}2���b��WZ���[ݥ�ZV)ڣ�yќbf�m�{�p�T�k�m\��S#�Պ��i]��}�����;���u����Rs�h�lv�#~`��z��;Mm���Tec:c���h��L���e�l�J�K5k9!P���<�-ƶ�4,L��f���Q�7�v���W�j>SMKH��%�wB�h�O�s��r����)�v�s'SYD�Lp�<�H�C5}ʐT�:ǊV;�����A��ꗝ%ѻ� ����u�v�,�F��%�vV��F��o结,NR��/�z����5��IفvU\k�UE��Kq�h��F֔DQ��A��(��Dm1�\���-�EH�*X�r�Źk&*���QYT��iX.ZV�CQ���Lh�RŌ�V,UU\k"��!�*��4�*����b��X��eUb�Z�TF("F1�
�@eDV(�U�h� *���D����5+S�J�m�F֍B�Ƹ�`�r��ڰ��Q��j�U�+�lR���c	�ISe����
��eb��IT-�̢8���T�Xc2�+�jE�[hV9C!�Q1��f["ˎdZ��Y�E�UXZS�8��r�aR�e`��cT�Q�2�VFҰ�0L�Ǝ0���YRT� ��T��
D�4(d�fol�L�>�qCk�|0�au�ʆU'��v���z�em`����eq�GE�S�+v�ru;��O7/���Ya�ͱ;S��e�>����<�b�sقy���=e�-�M���}��N7�k'�>��P���ɭLƉ��I��mWyi�?E�
�+����5n���h:�N�G3�}ї^��W�Z�N.��}P;��x�1=Kv��77��m�!(�u��ϻ�2��=�\/���_�6�3^[i��=��)�ޞ�{�1On
ɇ��t���ͦ�u�=�Z>�xdK�痃�������z�kK���L�B�a����W�ڨ�MW�{�츇 ��1���b�A��cj��5��H��q��6�MY�$^�,o,��<7\�������]�^^�q^Z�GM#�S�T�*��`о�:&=p�[Ṭ����
�J|���u;�.���~�fyC�+-rJ���8X��o�G��yW�bN�t�ܗ��|^-J}�)��0�y,i� Nv3�8׹g�=h�v�6�vD]�c�s
�z>�������[�;�Yf{��&��(��(oz��x�,MP��-�����=��2�$l#(�k�=��=����̼:�a���J�]/��bm�b�x���ǘI���.��@�g#�4�'D޾_���=`����Ӹ��� b�@��{l;�	�[��>Q�d�ŧ0&��M̬D�]YLq"D�\:�߾���l�$��.��؏&�y1�L7=�7�T#(e���M�j�pޥs�,SPI�p�wHR�U3�A2*��w���ku�[�O^����jx�� �\��{$�A�b��{!�k{=�U�C��k�#�X�P��.���O*kI����|��`G4̥}X���\��)S/����r�Z�p\�E�V,Lv�4�8-%�Z<�7�k#:�1�ۛ���;�,;�]O����S/Um�8)�8��eU�P�»�;�L�ʍ/Y�>�]�S�}��ר�P*�+���x)X{��"R`낞�#�
ac�ϮI����:��ji��׵�yL�̗�xk��3zX��Asٌ8Yh��r��5|�i��xױ�&��,�ߞQ�p�2�Q��)���&S63n��6���Ac}�z>���1��{�Y��l=��C�<5Tog�U�G��m5�ǥ������_\x=�&Nx�G(�[D��>���^���ݺg�Kl��z9�����Y�Y�N��W
\E�ɑ�Wr)���_�^[W��]�ynֻϬ����{e�<x��ܹ ���t�v�a��ϻ'L�=�c��s��IrU����yy���^��E3�:G\��]��r��κ"�8:��X<�J�G��s�Qچm��φBD��<��W+'�/��W]�Wƻ ���;ش�1�[K>ܶf}Nf��,=C=���'��=�:rq�՟R�_`��>�V.��'C��((x�����P���)���u,x�޷��z�ۉ���oS�]wx�w��Ս`l�EB����J�u�ϼ�l59C*�y���׈�0S��/:q�7ïc�Ξ��g��Zl.����q�eUq�uDrO���⚽��1^G�F;��7=^+U�S8�-|�bq�b{0���]�W�t�+���ю�C�\�ͯI��Z>�{f[o��3���'{M�z��b�jrDIT��94�]L���3,e4��C�~\r�(ߏuG��w��!gk��j�W.&Y���g�x!.P ��jYK��u���vl��q�����JԸ�\������=�b�衾G&\;+,�t$�*�˃Lu�k�"7���K(��=XM��^ҙ��Z��(�W}���୹W���+��Y�\��'�{#��]5���𭅣�jS<5��c���f,ޖ).�ʄU����Av!V��U� )R<,v������Ҳ��!+;a8��"��
�q��ڋY�����̉�t��c�n����pL��GeL:ÓT.r�bųBN�^R�|��̖�ݭ��س� �Aa���n����2�Q�}�(��(&n[��欠��u��1W��d`zc>�>�1�k�n�~U��J��t���$�o����us^�k�b��u�E�y-�G���̣�Լ��O�X\��;^��kF{�{��������ڌ����a5c��$9t�V�[�:y��^P�ڳKn8�ӽ_�~�8{��������x��1�6v�{�Y��H>
ߪyr�j��M�( ��r/C�S����/3����}�8���8�Pz�]N׌ ���]�7�L�m��?
�*'n���Oh�a7��	��[=).K��T�ꮡ4�>'�tP;���.��Z��w���ՋڝK�����W�p�'ɇ�E��RXI-���UOW�H���=7$WJy�$�܆� ̧�|��y��*�^#�047����w$�;��L9�����M;�b��O��=`c��X%	μ}��[�>��a�TG	4�v)�`�|y�/��:�e�wd��8+�(����e�/웜h�޼9·Zu�l��١J�p�����	�s/�]�̱G�m/,h��:/^H3n�(�[m��tS�ԝ�=��i�5��,��u2:T*@K�n��t�<<�!Y~NP��1%�z��W��9N��#�E
�SpJ(�������.h��),GP�F��W��
�K!�z(�R�Iɍ�3��VR�;4u�ɞ@�P�����Ü��>�ߖxO[9a�[7�K��U��;50�(��"M�B�_�>��;�^�/ڃ�T/}=g���hYt�Lٛo���14ӥ���y$��خ�����j���YS&C��&y�?�Ʒwz\^��`f7F֎t&��\9=I.���yh����Ŏ��)ծ�6/��Wi�5M�t�kǌ���Q#��Ӥ¡�]�d=�9W��D��f̵��Z�T�����'��N<WI	��箊��L&�3&���$���>���QhB�Ԭht�I[C;=�?N���X�uU�����'��qV�ѱ�:>����dR��2S�;C7w�;v&�*���Ϭo#�V���=y�۰��n&6�d\�����O[=�>�C�V��=|d�&�c����(عm�0���0���1�P�
�īZ�s0me0��śI�s+��Ƕ"����&��V;pyz�1�����s�	����W�G��ݱ���[�S�:�u�������3j����.��+X�يCgOq�%s��d���۾V-og!����F������3�d�d�g1����▬t����}��JE�G`������JZeGn�Z��s�������U��NQ�����o����?��P���������l���T���K�Aqu^����#h.|��l�8�/�	 �)p�u;�u���=t&(}²�!ai�͂:�;�jSY����Y��;��A�c���1P���&_�,i�����/�h�k�E��0����)�,a�7Ә�:s��/Đ���������V<�fo��&��(��ޯ} �Z�<6���j?ub��qd�D�K��\a �/�.�Ծ��Si�߹i�k�qd
��=��`����=&�!Թ�boC��NR�f5�PL����CO�^��\l��og]��O>gݍ��Y�ږ��Z�^��k�Α䮝B��=~�Kcn��!�E(�zom�u̞w� o�Z�L㾸�]��P�\��V,L�?ZHV�\���Ͳ=1�.�V�ț�����h_���J�����1B�T�:����vUQ���p1�;\^�:-��� ��ӻ���/W��2]Nq�ۑ�8���=K>���ı�]���x�Y�j'C�Skv�6�L���ƞMX�WT��k��ff�UJ��Jf�æ�;���eS}�:�.��d�.�sk����t����r���3C�4򫧏z��u��[�y�\+@�����Q�f]";���c�<0�cݒrxVe�S��]�~�p�:�Cm4|6�_�.O9�u����,rY�
�ٌ�f�yu?l
��A��w��ױ	����Cn��,��/3��qh�_T�\��%�I�E�/]�wޗ�F�o�� j��p�W�C>���Be�G��m5�ǥ\|LO�ȮV�0#���pI����|��z{$�#s�;����c�z�����Ŵ���:)�¬��/X�}6gxw^ð��`���-�f'.ϧå��g���Z<���V�,�~�1�{}GM�Mf̗;�5��4'�hjC�[���i���̺w9C��X����e3��=��������/l{��$h�Q��l����J�u��J�΢�Y焲��R���vI��^�oa����+Si���9�3
�Թq�$��TG_�O��x����b�˿k�^>>����o���{F�����ن�`�k����\\YA31��C�"oJ�[w���*z��2���NN�}^[�/]��H�`K�|94�]L��eg_�(���;���3e$-�v�yzBib���U�N
�ζ��	��@�vbۓr�<����՛�N���t'^u�}�*��pɷ�U�
��}�4Yqe�O�\T,4�:�%] ���9�u JZ��B�1b�}ŗ�1�G.�p�*�T��9Z����a�N����;���C���~��LM�P ��j[�g�k��nӝ����SZ�g�r\f7u�9��_���=��LZ}7��ˇp	~�Y}v�
�a�<*'}W�߻=q��%eAI��T'-�L�t���s��dA��ޯYᖏ�;�l�ٙݵ�^<>/��$/0"��G�y�8nU̖;�z�Y��%nT"��vv�G���z��[�y�����GM���8�K�g܀���k���pm�V3�\;s��9<��E�x��p7줣z,)(0t9^k	���iy������xY�������žg4�}���!߫���J�)��j��E����G[�>�炳���(q��Y��S&��p��^�yxa�^���[�j�u������x�OX�]������}^���T����k��j+E���2|��UxRz�P�FE�fg��b��ɮ��Z9,o���`>�)��g��V�{|s��V}�^�҇R��}A�y�Z�)��rOF..}�r<�����躛�r�G�vK�� +�;;�냒-��k�;��]5�)�*�n��v�A?�ŀ90f൞���ˋ~S5��J�h��A�a2�-[Z�YH�ע兕t5�YE��;��Pqt�����dəՈ����a�����˷�;�����_�Wg{Ti�u�{!�s�Vo�ҵ��>2�Z=*��O�5�	�lfs�e�5Swx@����^h<2[�<����8��������I�I>N�~lw]��YV-��������6Q��5�9����^3�����a�G$��l%�J��?�a:�P�rF��_���뭴�i�.T# �d̛|h���`:jƿZ=�ݠA����������ý�ش	I��(7y}j�b.T>������Y����O[8�U�~8�B�y�]{��.��
�5M���(8���A�WՁs�u��Zb��+�M�ญ��d���TC����;�p��Ƒ���+�du/�ۆ��V��j�$/�Jn�`��ӝg]h���ϺQ���',��ᘒ];�E�S���4|[smh�A�w���[�;}�V��]%mC�.�."F�8�sقy���O��Wj�4ʔI�3���E�><U׼6����=�b�	�LƉ�2Li��w�y����)\ɱ�d�0�좦4���w�������I.s4�fkG�sE-��hmNc�H]c�M���"�[�֋.��K7�
�Vv6)�lf҉�N�d�����E���L�r	#35L��'wE�r�74�H�Zo��Mӊʝ�2�����QN�V�{��WX�[������fz�O�m�����E�p}p>q�"Z�$�EP����K����G'3��f|�}a�9��(rm\C@ͻ���rǢf�y�iHn�Y�������t[{n������A�=�ayIp�\��s�	W1�u<ʜ;�H�Q��ja���-����A��%c#�{��V�3��P�u1+�����������$vSW�ǺN���c�gI0;�=����j[����7^�=n3e�+E..�gҾ^zqI�k����w���;�A�O�9�sJJ�WΦ�~��7�=��O]x���\���A�K�xH!�]�k�s5ȡ�lo�t��
�0�c%�0��9Z���P���l�j)�:���;x�D�1i�%�;�"9��v;)�%��3���&9�(oz��o���[�o��C��#��������	q~]H5+�yu6�����>�}_]-���9�e��W̺�X͎~V�;����q|���/J�����$ I?�H@�p	!I�xB���$����$�0$�	'�@�$���P$�	"��$�xB��0$�	'��$ I9H@�XB����$�$�	'��$ I?�	!I�`IO�H@�p$�	'�$�	'��PVI��a��@.�w��@���y�l�����c�:  � a��
%R��V�\v���kB�#YFl���%B@���:T�vd� -vk��v�m�6XF��5�mm� r]�M�i��U�����k[m6�T�֚Z 㸝m���ɶ��iqڮ�[fͣe�F6i*N;�ti3Q��2Z��g+5�kf�$n �:	�Zkm�4���vb�+M��խ��     ����SH4��4 рd��hE=��)R�` L 	��`昙2h�`��` ���S�CR�T�       i��&�&	��0`��$�@�	�1	�y	��Pbi�<)��=�G����|��*|���$���Od �!`?��I$ 2�?��g�D�c�T�	���� Vf�4ÒO�R C�p@Č&3*Ka-�4���߶�g3���|>���! �I�͗y�_�Рa���ϵ�2�:'0O����P�Y�q~��W>�zV�9����x�pYt��&K�["��Mb`�Q����Ԗ.��ؔ��զy7"C��jk���JѢ�n�v���u��;��r�!V�-���W���AH�f�X[��ߌ��h:z�}g.�!wn��qj�r��-<n��Գa�r!�^�Z�Y�=�jؼn�U�b\�`p�N�T߰8C�9�nY��Q�.黫WR�יMj�ɹjVQ���1�F]�W�����Y��mE��	�H�BA IЎ�22�����]�u�[ؗY�(�e��e�Y�l�T�T���ck�I��|j�w�+j��!1��(�?���������l۬nⶮ��+a�B�6�㫻�r�j[܂�f�t%�j��j��CFVlb�j�I�)�y���w�/%�#.��ۺG��c&Q۲��P+Y
9�Z�(Z�\�z�ti��"��ɷ579�3U�]][bfnmf�	�l1��Qqj�v���52f�M�02�r������lcF:���U��媋2:�(݄��n�M"i���E��3j�W2\߉`�?/��G�W
zl:ͬN��4y+ŉnP7d�A���������!���p^r�+k[����5��"�PTҕx��U�Ȩ)`�}�Z6�!�u���b��X4`"͇SMc{���l���v36BVo�J��Rӵ����>�u���N�Ҡe�U۽VM��A�৶2��d��2���S�A]z�T`V�7(5�����ʖغ����'Ȝg��l4f�,��a���F��ͧ�z*��4³��Y*�N��Y�� M���U�,�J�<��y�ʷ٩��F��w-���di�ݭ��©�'��="�K�R��;��3�*Օ�	���0<u�xn�d�É��Y��5�v�J�؄^]f-����sʹ����]��4��S3���,�It�Q*�ܺT˷uKf�[1ݩi��m�Wv9�[�0͙�$��u��D�����7n�ѓE�,|�+U��Jt�U�*�� �(��a�"Q"�^;�j��/-e\���g^��^���F�X7�v��/�쥔CY��n��n�T�Y5cqi�� �����0��f5�n��=F6o ��e�	�V������tM64iA��cU�<��~^�����~��M	g��느s^=��iF�`�5�����{�=�z�c:��)H݌+�s�C�Vr
@{�Ե��aޑM�(ɹҤ J��ug�'U��*,����ܷKpǗ#��kji2jfmI��7:��x�s�鹗)5<n���h�Z����/5�{�:��u�Ҋ�e�s.��Zs�!�s������G7;0ks.7�Thp�Sl)�ɷnw��fC[8�w�c(H�](nF��
Trq�ɬ�N�qR���	[�P�}��*��l��N��l�o��Ӡ`gm�6�kxܭ�6m��q��ak�J[��Y��oi�ӹ�a�"X�9�yҰY�=&��aߍnrU��b)�ض�I��(��]/:rQ�JM�[Xy�e��1������o{4�8ά۳-c�k3H�ָ�.�r��x�'�$�U7z�r4�ZIf໷�k
�V���b�roVtڽ��(D^Ċ�Vkl�`�J���w-�b��72t�W�o�62�.�a͵�\��Ը3t�RHK�5��Kɵ��弆dʐ��q�;�����T:�>B���/��ff��Z ��jtP��;N�yr���UX�ld�n*p;�2аes�8���v"F�u�rs�R"���|���ر�Esr��JS��cH�䗗N{���*��z�uc8}+��y􋞻�]�j����>*��:zX,��Hq5"֤����0E·�aYD�(��A��7KE���F�Vu��x�H�.�.�I|�vŏeK�M���d����O��t�h�մa�.�g�����KUeh��!�mw��5]Gw�f�i�u��t)+�i�������r��R���㲹�8)'Z�-M���(P�(���^��K���-V�n[��,������{��U����Q�\�C/��8�lYt�]�0e<}+J��\j�I�Ǎf]h�s
R��;ZS��UI9�\���H����<"g�8*[T��|k;6KrȾGɘ�w;�y[,��Z���OQ:��:�_��H`|�`�U��'J��Ӽ.I�F�)��G\1I&���wI�PY�.vn��r��dە�)��3�5>�Ɵuj���ѥDΈY�����ؾA.U'Tݗr�5m��h�g5�U�T)J��-�  ��>����{@X\=
�SY˩b�Sj���+���j�G�!zw��p.	ّ_B�K�eֺ����o]oX��������<y�_~2y��H�:�:ɝ$!*��>�:=��p� f�}�3��z�cإ�W�<4#�|b��3�D�و۩�JU��IH�.5������1hAF�8m_��eJ��`g+7z�م�W�2 ���Y�UךLٌl��,^�u�sj�C�j��n��\c/�tA��hMk�%b�W˾�wOm�Ws%a��:��zC{�([
1�5:bP j˯H��� �����c2���t���`���9�B�C|��0"V����v��,���%!�ܺ��H���']�:l��$-B�P{Dm�
��(�����\Ѻ����6gɪ]���ٸ�;�����i����
VX�QAi.Ʒ3�K�wt��r�a#�m���^]^δ�Dn�gRwm�8�8�릫p�5q-L�Ź��Nf��bf��Ahn��+p�\���u���jp�tYnK�]���9��0���;V`:��h��++]�H.i�zZu�]�/tS2����R��ysr.T�`m�hһ�7�bGB��  1J�A]���e�WOn�C]ϸNoY/6�4摪��tL��ݲ#�Q�C�rӝ]�P�]�+���R�I5�
�����b�J���k�������ՅQ��w���W�uN�2BlX�Z�Nx�ԩ�۷soeX�Y�("u��v��t�Cu����7�,ۻa�M���SB�mx�a��)��yV\
��CcR-�E� ��os[̅�H�vݻ���7t	�\���.��_d4+���
��]@���CIW��M�0VS�Q��X�g�+��Wi���Yê��11(�}wX��՝�L �O0��]t� �]J��˫b��≲�
�ľ���]�I�kj�I�y,8��CU����[���B�$*1���Kk0Ļ����U�*@��&5PWR��~5v:�n;�Օd:p
k���Dsg+��!\����޵X�;�J���Q/fVب�-Dd�x��̺��O.���P�� �f �D�K}tv���A�p]6�*�3��NY��v�/��ƊkZG�v�K2���p�G.�ʚPX���ځ�q4�r�^�ꍷG�1���ٖ�dKӵc�(ԍWg�4LQ7VY'��3S��-�xp\.`ˤ�+c:�,H�F���/��@��C�F6�.Yܛ=�ұ�<�È�i7ǇI��#[I]+�:�'1���Emn�9�yI�HE"���j!�\�'�ɜ��۟�\�M��[��\]V�!�[����eD������)	���P;Z\L���ks(�i=��Lbk�a$�����ʖ.Ĝ��κ�I̳�s�l)��(�k�oe��w�u:���w�@�*�#��(�e%QE��RHm)��+PP�� �A""SQ��Q��Lw��Ks^٪����� |.��dC�֫��4̏���T�T�1����M&�MUS�0�e�3���f�c:� �i�p��F�8ջ�ɧhSH�zI�\�:r���;}f�'"b�qf�zǸ!Fu��鴞��A"R���V�W_r蜦���Bv�ޙ��m4����I)���a����eф�`���!�5��(�Zm�JH�=�7�sW�nܦ\'*�IM�=gMb���e�(pE0ugz捳)]�i��kl2����
sY����i�+��4�O���ʣ,���=���D^M�ͻݫ��A]q�|�g[��V�wv����� @���RSƛr�ﮯ�6��L3�XRm3��7�0��l�a�����m"��\��E�]fҶ��-��-T�˩�Ӕ�,�KgI��ɦ)���-!�S
��3)l��-�(��s
Nf�M:t�L��fq�ɜ��e���^Z#ﲗ��3pL���Wz��7�=ˎ�h9V�7�t�C�����ܦ��"<���XQl�ׁ�z�S
p��{ι��a0ɖn�(it��%�U�L��1�¦�R^�d���{L'L��,�t��E'6WL�2��ҘZN�u��zɗlx�����4�y��w��1�C	�8�j���/�+��}�RBX鵽�R�nΛ!}�l���8��(���v3Hv�r��i�(\���e��i�eÆt�|�)����t��U�s�\�l�c��m!��閂���y���+�H�д--�gδ-uE�zr�m-z9V��%���/6�-��2��gi��cT+��b٦i��N9���\�]ߝ�q���{2��cc[�8o:�S��kX��';�������3�V{�6�;i�Ӵ��,�^r��I�oeN����"(@g�F��
g���b��[�c5݆n����[��R.�]�z�=&R�\9�SI�WL��L�6�&*�k	܃F4`�",D��LB��۫L���M=j�!L��l�e���b8B�� �q�g�����4#�[�Ю��v�fn$#�P�t{�VZ�p Y�9ya����S�֝�v��}w�m��TÜ��Q}o��6e=0�-��4Qiγ��.�ꡛ����Ǯ��^x�̧BZa%������N���X��S"L2���T��j�2����0�sM3��$�(�y�]��q��p�B"G�w�Rv��Mj:�TU�J����Z+ztn
�Z��+���T�#���'�TÔP�m��'�C-�L������C��QY�n���(`���uy�b4G��E�.f�AV�DhcѢ �B��/kU%Z 0�'H[L���x/�5�]e�д;8򷌺�FuGL�ua���5���P����P���E��x�?ifͧ"��tAW��~������g�q�im2�gIL/L;�gM[n�i�ч�K޻�i6w���63=3�P�
��ӧ)��qE�NQk��bq&�)����i�a�n�g�J%���Vr�s���l6�I{��cX�m��)kX��o�B��#�!@�e��#LMٓ����λ��q�o]��,T�B�=�e%�w�]g؍;�7�3��-�v�G��9��i��2�L�1��ٶ�E���r��0��N0�IhSL��l/�ݙ�CHa��q-�αٜ�:x�(���!z��Nq�!��7C��r̳<��ծ�L&�e���������M�N�[/5���d��<UOɂZY���g��@V�wEЦ6�V�:ԩw"�\Uu��輚�]&��M�޸�@�62��3o)
4�!zrr�7Ql:^��Q�X���������'M�ɛ[�j@�}�ص+u���Z���Y]���OTg*+9d�]IRy0­����(v2A}��S)u�	��; �K�<װ�q㉪��]�Ⱥ��p��T�rP �ڶn�ѵ "!���E�N=�x�������
��r0�.@�ް��c�a�,����%�6��������ͬu���þ1�Q�)"Ȣ�X��) �b1���2"(��"EQ�TcTTH���*DH�,�|�z�����nf��"���!�{Yz5��'Iy�,Ô2�!lֻ�Oi��Y�]r�y����+�o��)�[0�N,P�8%b�̧3^�����)%�I���F���X�\�B�D�-����z�9�s�������	-
i���n����i�T2�-<�����!&-"��D����{y�]�L:3"�VJ�W�������=7��_�v�N3x(�]<�Z�wSL��I�-����m3	\�a'X��7�oC�8�I��e2���w����d���p��y��M3i�^k:�&]"�z4U�k��y�ˇi�Q�;��JB���a�u�۷WD��ش��Nq]P�;�t�8���QZ�kp��|iq��7�AU��)�g*��d�[K���G MOD�Q.��`��j��B��Ɏ�4�6�ŵ�1�Y���ռ��yK��Db�ҫ���U"���Hs":�z�k~��v�m�]7+:N�� 	P����F���n���i�"/�e���8y�![�5ӈ���o�x��23��ǄTy����\6I��{��bU
8��Y0�����ˬV�nKͼЫ�]T����ȭ:�Ò�h�Z����y�հP'N�XӞkÝ�1��m�A�^:y��
_I����Iq[p����>)����w�����n�� ���|����T�x��'r�����;ݨ�y� ګ/e#0h��%gu�15�P��;h2��[SNԨ��_�V����+f�t^��کIw����j����\!��P!ٷ�:UW�)̞�8�G�P�޼<{p��p��0s���1=tE[󧬴���"�g��cuz�j z�g��Ry�oE"�y�N�;0"�KNZ~�#oJ��,x�%ؗ���+������o:[�y������'z&�[��}�Ů�":n���ȱCOisuu���S���N�'7Uv��b�,�[�=ud_D��n�ܻ7���S���9ϩ'Vwz��(��!�#e����c�`{MU��r�.�*?sig.�L+�nۙ��Ϗ��bB��n��:(^�N�y�H=�9��)Vɒu�x��TT|�P���t����j���ǫΗfri�9�p��ȵE{��u�V��=)���ĳ�2��}�*)�j�`��3�p�:ȫ�ɨY�xn��h�j3�ųW*��}�}�?��K��)��8�:��Vj�U����o[+��3����]/%:�� k.��T�(.�\�c��,3�ʝ4Ү�h�+0�R���7c����GX��*�IG�[� ���Y2�L�:b����r�Y[H-��9oF���d3���4R�1 r� ���Z	��p��o�Bw Q��\;pS4��1i�"@��H	�������ٝk�e,1:�u6튝U�\ ޮf��Pk��k1K�����$���5��κ/Y굮�o���<|�3�#$
�2�"�",H���
`#(� UR*0Y���gyyu���s�cWU�c�H���v�-�D����r�$0�$0�@% [q$��q$!�f��x�}�c5$;I����	8ɔ�W,���H[$:I!0�ᄘa������@8�Hv�L��Hv��'i(U��2�HI
d�Hi$+u�2�޺��y��M0	�Ht�$%0���y�!�Y�2��I$��c;t2��d�I!�@���a! ���RI�v���G��G� �D[�q�y�Uo7�h۩�R�͐�6�3���ޏ�{�b"(DE��I'��$;I&��ߌWY�$:
@�I�K`Lb��1����3�WJ�8>qwe|f�b�˜��U.Sħ��m߻����!�H��B���f�[������=�^IV���+�����k���-{��}��{#�ec/�n�6��M�V����\0�V {Z:���-�gg-F�d3��q4D
�k�}�����#��9Јt����ۍNw����3R)���=�pݱ�h���@�8Sz�S�W�o����`o��Z���\���>A���ޚ�������=M vn�^M��/y����r�0e����&����X@V%��/��]���R�X�<�.��rΓ�K4���4wќ+W���gz�4�k|k��7ݝ9N��aџU߳/�f�1���X#����/��Ѻmo[�G#y�@z�od�����!�x�&��7�L^ �ļ��b-<z#6�~��/o�,��@NﶠM3H`>����O��B�첇��cܯ0�`�G�l�||e�˜"�/V*���]ePN���A]����שK���	ϙ�+�'L�g�v]"
�ET)=+`v�;j�m� oV�}� U��t4�on�&�-?E����*g�ڠ����X�g3rT�o���ǧ"v��5:^��^x�>z�G�O������#�0<�5�����mr���h���q�s	�v��G�Tj���]���2�(��6�u���	�Q�<��:��y�{laSN�|b"$�q4�I܎��;�r�ɋo��zf*�j@k�CV�1e��yo
u~���ʗ{�$^�U�������:��3�i5,�zd�f���B��l��1W]����7��Hdn,
.)ӱ��'!9n��c�=��7��|�C �/���.M��v.w��ޔn�wC���Ɂ��˜"��<�8�Mg�4�ī�z	N��ΑqWCqW���89�V�v�mt����6,�O$�(�w�A:�;v�Z�:��|��W�F���7ԧS<U8�Zgm�(28.e��a���Ym�*����  � *
A�V*��b��EAUU��`�,���J�PX���
"E�-��v�=Gzz���ה�J_��X�����˜��7z�-L�^�͔(�V�酚�1</����,WJP���ţ3�s��+����,���}�I^���v9W<�݈��a�S�6�'*��{�P^����ǷZ=� ��`z燦!+<�����d#F�Í��}�9�Z�Tx���bA�P0�..ֿmy�߆�&�'	Ʃ�W��<��kˎ`!>��;�3'$����3�[T�Ύ�\��-�WXy�9>�\~O�V� ����O݋�"�nz�JԨ�ny�<�VБi9�u�!g�����_x�_"�=��Ϝ��_�"t�@pJ�w���VvB�޷�n�\�4^x��
�adz�H[t��7w0���4�� E��P���bq����AL��h��郣��|L�!��©0k+��&\]v�2�yf=B�
q��?]�9F��{0�%�[ѿ���;�8l�G�;[;�v8����f���'�s��G��]��?��D������\ʘ���ߝ���R%!�n;�Vnf�ߕ�\��ЮXQ�����S���u�c9UHކ�aҲ����Dk� ov�c�3�t�b8w�U�� ���8u!�� ���щ��W��`�כP�Ӷ@�G���*,Ƀ	T3�X��앖�NB T�f�&V�:*�"�f{��i#dC!Lm�9�Huܻ��]�m�ލ��6�~��3�0�j�G�j&���C�ۍg��E�T�å����X��Ʒ}鍇��F��
�k5�GX+,k�gV����Tj��j�S|(Z���`�݌�wju�E~���	��ًs��ۏ�X���O���P�ꦄ�\dn�:�:�G;ݐr�����t�]7I�YC^]̓�	`K� 8��e\�[܆��z�g~�DDBP���r�l��R��2~�����:T>�P����۱�$ҭY|6��y^
��"�EF��1���J��u�p6:�u���lȨ�h\$��I���&g!{�����fSU��q��ZT�i�/(
�BmB
�}�ah���u�~ER��+�ϊ��	|��6#yZ.�muҮ�]�@�"!��Z�o��uB��r�c8�j��)n��+6�p����M�U�T�+%Ӓ�|ڧl�ݔ#U�ݙ�Vd=�������J�q��0l7�${�Jeoz�pԾ��-Ġ�7%����9MC'mЊƈd�K�W��b���k�o:�.�%0Qe2RD��C�R�S��HS"ȫHLc|��\�y����\�u��R?1<�����O�č϶X'-mJHɡjƓ�qZ8���5�ކ�&��_j�,Q��7H��3�u��v��l��b����Q촜C:�L{��W��{ފ������b�_K��P�*r�Oe�9�C�˦���������K�%�ǔ��)ټcM��Vэe�z��ET�^��iv�~�Ϫ6�V��^�;��-��ޑ��/7�#��x�� �L���=~��oYv�K�^��9�oe�勔F���6u���f�KM9����|�b����̎�ɧ�@�S����L�L�����o�65N��U���{ޒ�8��3V�g0H�� s�T��˨?'f,�1��~��Q�r����Z����<�Ӥu�H<�#�:E���6����t������Ʉ�R����:U�oL�ވ�y/�g��{=�_�m�1���ߛ�.�#o�gh=Q�3��|���te��|�˰��$�F�J�jcf|x\���o��D/�D+��w��{�����^k��D{�W�3�
�T����f���w��;O挻h46��,�sCn��SF7�v^�����=喳d���*�H�
֗���ܨw�?v����	q�z�W��{ޤ��}�ݥ��O���Q�X׻|"�P�9���|*g�"*+	��m�����0��Q�Iy�c0_k�dۙ�\����J�w���h]�h�<���=�z"f��u_D���Po�D�sf2�Ȁd�5R�����|+X��3Ǌڻ�Վ���*����g�'߯*7��u;1xT���C��ϝ�7�ʙ�׮ݿ�芙�W�b@Z�1�(�mg�X ��8vn+F���7dED�ڛW�б qL��]%�;�//�%m���e�]���\,M1���OV=J�]C���t;?Dz#Х7�5u/uN��_�wm־y=b���ڝƐU��ׂ�a�lI�!z��p�i���cEb�ॼ3�1�K^��3�֕�R�l��J�!/^D9�'��l�q^�f���e��v)���]��ܓ�c���V�U���F�tTi��K8bߌLV�Q&�����f��d�V�
[���n��L|x�6�t��Ktv�c/M�pR��n����\�i���54���"��(�jg�-�P��p Λ���)� a�1������ڈu$ٽ<2V�W�]�3�h�[�)m6\Ut�"��J7�*��"�,��,L�^5}z&�±�)��4�T�
�ZAJic�X,U�0�*�UJS)�P�\�7�׏*�ޱKz7)����{�3F��#N���U�e��{ѩt��s�+<oAy[f���&��ƒ�D���rn,MřP������08j��N�a�=&v1V�5妸1��O'+v��m�=��=蔨߂%�(~��F�P��ľ7J�g�����gzJ�r)�,�� 0�ޘ/V�W�]�櫊 cڜ��z�OC=ʮ�=�އ=G�b�]<���՝7��{ބ�;P�韦�PG�a3Jh	(�>?+�ŏK�z�vg�և=qxקW=�: ��΂���4��V;�i�V��ۘ�]u�e�`����oV޼�����IU���_�����S���gNѫ��Y�諽��x�y
��V��F��V%y̇�t<�o�T��'w��#J[�u��[%~u�6of9KaG�9�[�����\����ݪ�j�-��b�a_% �Ǹݼ�,{�X��WM�޽�6ߏet��$�pN�����w3eF�N��^J�s��-�y��X�q�/6�~�G����#��@h?L����Y���f���G��x�-���yS��=6�k�un΃�kV����2�V���NG���!���tŗ̽��r7�'w"�}�}�b��9���)�Y�>����R���q��_n��-\>Y/�앷W��[ ʝ;�������f��ա�B����@�s��{$�7��߽�DBQ�a�om<6�}*�'gP��.$�2��E�u�ʪ�y26���x�ST������ǯ���6�n��pm���`ct�A����S���O�����������W��a0B�����F጗�R�C߆�$s�]
�uifhC���*f�@�N{5j�}=��ͥ��Oj�l'F�Ꮵ�W-�ϱ�7���L�_g��R�ouW��DJY�3}'촧ǉ�~ߺ�}w|���1vՊD=��TD���{F	�&s�q_6<��92��j=tq�Y�]�g�y���}���E����j��֪'!QYպ���\W�s"�d�l���kq����|�H�n�/Z��8M�������[�Ox�s��B�x W�N�}���^]Vn	]���O YYE�
dXzR��N�	����b�"[���JN@��f9@�y�y�����.4���e�[a�`%��Vf�cj�n�#c���|�}7
��&�phy�{f^+:�O��.�Qt.m��fY�Ge���|��,��k���[�s�tj��2�H�@S
SH(��-4�%#T�R,P�P���-1AH����&�[�5��F2������}���G}j���u�t��ՙ�L�Z�Ӫ�M�җ�Wh0t�0!��(����ˉ4����f����]E�xn��>}]�z9Iݫ�V�;�qt�����5�C�H?{&�uH{ِɎ��Vv�5�xt���+����ǲVం�Y0|~a]�[�3#�߰ե��T�}d�6i��m�Y�S�t��}�.}�d�J�H~��KOl�:������K�g�ǖ�v�ﵽ�p�����Y`�^�7G�)��Z+l;�얝̄̊G^��;�\�#��F�]��z�$�ϩ�}9�6=P��Xsif�'�[��(O@�����N���UK�����R����)�뙕e �%y.0*�>�#aמG+��aT=c�;}�
7��N����iX>mʇ���]s*�M:�ZMa�F�̬"����|����&��ַ��잝V�^q�W~�܇N
���)���~@b��(k�:'ݒ���\�P^��sƦ8/fLمͫA�T4n��x�C�%�	�V���d��0읾����2��Q�^�w��T�fH�;����h���BϤR��I�=4�s�n��b�����֊H��7z�@�$Dn�	��}c�J�]\=��`ۻ\;���B��4�@�ױ��m2}��8�w�[;�<>��nq؅䎔p�GOl�W�P��� �*~Y��fL�p`P�Ox���f���Z^��f�^�3Z����t��1��vh��:�SQB 5V��b'��k�-�F�4�K/E�y���Q���YSs�ye@���g��F������י�P,��{{�L�a(x�~��׽�9>�/�L�΅g�~�6X��Xկ�.TG�Al��!����ޝm �>�x�e��G{�ʷ[K�L�����Z�����"~�</q-���Ǜv�/�5e�J�~�i��QHЁ}�����̤Oݑm�a�<[mo�؅\����]LY�66U��iJ��5��/@ l������{Z�4GVU�ShfvR�R�jW�Y3��4[8�m)Q�#hύԔq�_jܪ/���cj�gKt+�K�-�¬[�m(��s�ڸƷԆ�>K���P�ٹF.�o\�Ы.�Gf�8�wE��yٝ�.�i�':L'�m������EW�`Vt7r��NZ�&X�0	#�ً"��$��N|�1x�Z�1έ�x�/R�����
S
i�ʩR��AM%"0EF���jP�5B�j���%S)��*���e4+����Q���JU+)�"4ň��UE%]0{��y��z>o`�а��}6���,A��+���-�1k(]<��:J�E�B��>*����=pUˬ�O��lF�]����t��8���y@��|o1v��ٳ��)���4
�����}pի��搹x9�Ы\9�dU���@��v\K쌓�ި��=�8m�)�&���^f��^9���X��oW�jl��Ǌzԣ�QS�C��_ �a�Sq��3= ��#���d)� L`��Sr�����7y�P�����I�Ĳ*ڿ>:��7�_��c��U�FOLa�%��+��s��>�e�%�=k�(�m88����V��ډN9`J6��ӝ؃Ö���W�s�p�tL
�Gʣ�h�P�72�zk�g��;��u��i�:�f�0ao���4����-un\;�x8�G[v5Z8��<}^c�'�+��`3O#���4�#�i�o=ٛ*�+)��n���r�-�v5���<X������GfL��ل��Ǌ�q����|}��"�U����K�	p�E�����kj@H�E1p..sj�>�/׏ӔG�7��ε��qx�	��Zi�k.��U�}#��s�"�~���sk<��"Lb]����G��$��TX/j��i��[������=7����{�_�u�L�����t�o�r��.:rb�`ޚGl�����\��ʔTW�Z�4_7j>*��T�3�~+��/<�;u/)h�
3��X�f3u�=��b�k���`�Oe���̵��Q��rϕv�g�Dh�#��wovd��9�4KFT�P�Jy�ᖄ�Ɇ�mK!C�k�9�v˵�3�w�9�-�Z�"�"�Womv1T���^�*oL�+\�1aw�_�%��}ؐ���i���"�5A;���jY�̆M�:^���땃���Y����an��L�U#��&Jz
���qb�lU�]�S[��E��oy�`yw��0�)�MClcyҷiMQd���s�SE=�w{P��F�Fdވ�e�����=�mڗs0��R��W���ql��4i�ɲ:n�{�X&��&���~N���4_�I� �t�\��^��_Nͥ��+��L��ь�@9+��Ay�3s��ei+W����%��h���gJ��29��3��O�7���3�Y5c�\0�
S�
RAV�4�SJ��QMAi(b�L*�e$bR*�����������i��j��T�����$R�J��i�)�"Ɗ�E"SL* �D�(j��1��)V-UR��2��j���Z��UJ*SEER0��(JJ��*��F���*�T��SB%R�R������^������!wN� ��u����y��=7?V]�U�Q{&۩����q43�2�M��mu8��&R̺Uw^�x��W����.�� ��Kކµ
A��ʬgU���;Ż:l��w�Y��,.���Z�(�6d�iĺ���њ�,�=n�j��H_�����j�����^]�\c��<���~F0<�*�q��BN����9��1��� �%�mM+=�Y��Lbא�
94�Ƈ�en�����D��5WV/�� ��<��d;����<���o�)�
����R����s:��|\�r����Ӈ�2�x6g��dޘ\�5w�t�b<�篶�.&�i�ԛ�E���YUgG�n)f�e�0T�˻����qLz/DG��v{f���"�7�o�]��|l#�Q�Z�7�	�����,�d�2W�K�w�oi�Ѽ��^����}��F�\ �=�o��X�$>Y��hb�Ws��:f��p{��r��Z�=�����'���6�y��'S�>�d��sL��`��;um�(�N����O��"�Q�z[Kc��	Bo��]�����%Ӕ�"{?DC7
�I�n�O�MH3c�|_"�ֺu-e＋Ǔ��'�1l؞�3Wr��D
�-�BY���e{����h�:}��7�Q��� �+��)��n�]��ߞ
L}e��4YxB����i'�x<oI����{�ϼ��@��ʢ���U�I0�]>>��W �]�.-t��kWP��cd��;3�O���$Wn�P���e?�˺�������Zz�ytn]��G3�o,����5�NwV.�FS�7ğKy��7�+"��A��k)l��y���1Zpm(Uk�+ f0gշ��]r;f�MZ��V�����~�ݍ��K�0�A_�{-<~������S��5�"꾍�_Wۢ�[��R�����BV���[�m>�����;L���D�#CXU�2³�Q�U@���6��ƯPU�Ӣ]mЬv��J�s7za��3��}\�����"%���\5�:�&��z�c�]v]}�Tܙq>�Ʌ�mDE�c����O�hV/�u%qFgmL��Y&	"���\��6K@��4��{#} n��;`�R)
���B��K�m�:�X4��Y=b, D z*"-TD����%
�*�(Dh�����Z*��TUQE
�)Z�(�Q�USM ��JU"�PX��Ei��*����H�*���`��]_�V����R����t���q��圪˻C�i,�SYk1k>�@��s���Z�n�㕼q�T��{�K��Ɔ�t[�k�z�4��=���-Ȥr��Q�>NY�^�m�`�1����^c����t�]f_j� u�s\y��і�M�5����rQ{.�F�jφmg��f4��rh�η��e��e�9	��w�=Q����;'��]o������2�`R`Y�7f?\(��6@�PV�_�^�f���*))lа�a�:�"w)o-�Jۭ����U�������/�̾lNBv���<H��ae�Sx,n	#�wyz 7+w
u�ɥ�e5��,u��]BL�<��
Y����� vI��g�%4(���c�YF���j�^�]�h�tq��>�lk8���p�і(b+EL^S��^�� �띴�����=[X3�7W�q�2�G����*;�(nh���i���,����@I�0{
1�Hvȩo�S�U����S�|s����Ǹ�kAV�S��ټ/��:���{1��m]��sJ�$@*�tk��/ �P�
��H����Q�1^ΩFs��&��Dͦ����P8�:��C �\�1]z�� �����x�=�ɘ��s� t"��5|%�zLJ���^T_�"{\3������:ۥh����
��_��������-��go����E֝n��egԼ�Xn��002��u�_��s���ô7h��	o"���q�������]�["�9��9��/6�&rn�@��Ħ'e8S�����v�<\���Z�Pw������}�}z�`�7���)q�������s�tn�^��cx�nr޽z��� EN��!��J*�8�]��\WHS0�{�.o�Z"D�W��c��;4�����]�~�� ����F�_�_�_�_�@��b��)�TQU��D��A�����	 ������! �Q�3P����*����WP�:�+o����c:1;�K`�CՐ&]�  ���X₁&yarz�FC��P�f3�`&aRWT�������C�	��t,�u��Y�<o/����_sǈy�o���o~���/�?��p�ޮ�9��v�%@rY<vfy�W���;������^x��#�@�n�!$Ĉ�?�O�aRY�?��쇺������|@�3r�����������=����$$��~u�����`�%��g�����o��&`):�/6�+�q�U}W�3���4����������U!'��B@ �I>����d�/b\3!	$���$�A©'2J,��Wl�]��?MM���<�����$$S@i�^ٮO���'s���ks�?l��j/���\�M���Г>\@?����3��T�y����_ e�r�t��� ���=?��1G�OMz���P�?/�|��#_G�����d?�zp>�;��5��?y�Cg��BI�0y����,?��yfNr�,S�B��݀���9!�7����럺I��;u�>mB��Yw?"���:8d�I=���h�� CA���F$��Z���!�\nM��}��~}���]�4D����Ip5�>�e��P�frc�J�1$$%���#����H~G�	� �>��������O��w�y���i?�О�Y$�|}�劏�>�B���H}>>3���a�Bq��>�#d���P��C�>s�>���$���TH|�����B�K��4���,�ߠ�:��~�|�z��	g�}�w`k0� 7
*�Υ�.�
�y�3���o��:�����?j�����s�����T=4�|}�=�1��Ĉu�ߝ|0j��P��C��C����Toߪ���`�A�ɘ����#!$���=I���o�z�}:������'�h1�{��MC9��Rp`gw�\���Ԟb,�D��P��(O�s���H�
.��