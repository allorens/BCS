BZh91AY&SY�ю�L_�`q���b� ����bF���        pz�R �("J����UD�U���B�D(�*UH��!(QE �P��@��EU@��l*$�UD�E �UJ��HIB��@QH!Q%(�����D������J�T)J���"�  Ţ��'�6�R)$��X��A&h�T�T�B���J�R�TH��P$T"�R�P"PB��J �
���!*�   ���"��J��6±�Mke5T��Zm�mh�lh�K�څ��ij�DJF�Z��Ki�f���j�f�DD�� ����  ��
��R�F�@J�fK��IҘ ���U!*6� �UȻ8t�Aa0k@YK )E�� �w�BJJ(DI `  \�R�k *�Fښ� 6�Ī����B�+��pB�IԹګ��V�e\���'S�� S�T�� �B�D*��$D)�   D��R��ܺv�P	���*P^9�T�q��T� \�˝� b� ԁ.���)Up�: ���N��e
c$
���@��B�R�  �8we R�L � ,��*��\��ҨR�9�Js]�ӠҨ���UJT�ݩ��Q��;`�p�uT�*PH(*��  +���u]�.ڪhU��J�JX1�@X-Je@ZN�UEt�t)�hR�Ph�ª�EIa0 4�RIA!
(�TU	(�8   M5�t�6� 
� ���j,�Ѩ@l� 4+2����F kZ����Q	)(���U�  8 l�  XS S ԰ 
�� 6�c@�X�kB4� Z�h U*P��UUR
�@)   M8
 X�m#�	�hP!�  3V  ` hh6( ,H�l� �mE*���(UD�   mp �` 	�0 4mC 4�
 V�` �0 �X( �`
��� 4<�    �  ���R� ��L��i�"�ф��(     0"�&	�ji�Sd�!�M11A�����4a2h���ш�sLL & & 0 $���E*4�    kϩ�Ï=�Z_��Rsθ�g7r�ql��s�^�\��gl�� �
���� V� �*oEx��
��<�_o+��@`��b����(��<!E�oG?0�,&�%Nd�Nd�	�`�Nd�a�Nd�a�Nl����y��y��y��&�a�Nd�Nd�Nd�f`�^a�a�Nd�d�y���9��9��y��9����y��9��y��9���s.d�N`�`�Nd�Nd����9��9��y��&�`�d�Nd�a�Nd�rs/0s0s10s/2s$�9��y��9��3s&d�`�`�Na�N`�0�0s'2s0s70L����̜����fy�0�0s/2�'0s'9����9��9��9��&9��9��9��9��9����9��y��9��9���f`�Nd�a�a�nd�9��9��9��̙��s��̜�̜�̼����<��<�̼�̜��L��̼��0�s <§0�̈�
<�2!�$��2�(�*0�s*��0#�
f�T̠�(<ȏ2�(�(<�2��f@�Ps�0���
<�0� � <�̊L��"<��(�*�0#�*M̠�*<�0� �
�ȯ0)�
s+̈� <2�"s ��/2��"�
L�̊s*<�0)��(<§0� �$ȧ0�� �*��0���(<�'2̉0/0+̊s(<ʇ2)̪s <�'2)�(���0)2�� � <�0��s(<�2+̉�2� �"<§2#̈�*��0��C��e0�� � <��0���/2̈�
<��0#̨�
�ȏ2�̓<�0�� �ȏ0̪s��fT9�\�/2s�0�̨�"��<Ȅ�2̂�̢�/2'0#0�s��	�(�)��� �"<0+�¯0�(� ���y�0 s*<ʏ0���
��9�C0+�� ���2+�"�
��� ��*�̂ʁ̢�'2�̂�
<��0�s s"�*<��2�� �	�*� ��/2�̂s/0f9�0�2s2�'2����<�s/0���L���<��<�̜��rs.a9��y��y���I��9��9��9��9��̹��y��y��3<Øy��y��y��9�g�9��y��y��x`��.a�e�C�g2sa�a��d�fg�a9��Ne�Na�^e�g3�9��y��y��y��&9��y���9��9���&^`9��y��y�fa�^d�e�d�	�a�a�^a�a�`�fNa�Na�Nd�^a��y��y��e�^�0��m|m6��Kr�|�ur#,�V�{hbsv�V�N��N�Ǆb��I$M��J�1����ʥ�6����j�JW��y���ґ����4R7�����[	8Un��v�5�f;������I�ΔI����/w-����CD6����<zm&o2�dD��bf�l�U*n-y�\C7�Udc&	������R����"h��Iy�:T�M��dۻ�
���/L�& Ϊ�"Y���-����mBN$�c(Y�V�c�Oe�	�w1MX.=�q��
���k������c.v)J� Sŕm�˻j�d&�b�WC�˗�L�⽐���T֌�f�t��f��[��ʑS�FB����	{kY��6.3R鋧wM�{7��tܑ=�M'*�z�n5��N�Q�o;�7 ��Y�B�:ث�˷�Wx"��ŗ��v��Uy�c�V�A�ى�LC1��ƉE[	����Z���	q�DiكJ�2���k>uͼ�d��KN�C�yb"Q��G`�Y��M@@mU�����DT8�3S
��Y�O3�M�մfUr���ZK�u�!�oUeO�zc��r�a6����ڷ�i�jѥ��Oo��(1x��v�ee2!kM���Z[jL���N�e;���"���A_a�K�f�����\�P�J�ʎ�V�z�o\�;Q?���0��,"�ȓ�;.���&�v��n��Q�0���*Gv�nYd�:SK%���D��GW���(

$m;cv��	r�|v��#Qt�Kh]�ۛ�����f[���̩�G�,^�U\���[h�մ���!�m�$�`����`�+5���*б��Q�'6]3+"[r�GnP�D��]��7�n�Qi{	�����(+&�LU���C4kv��%^xk��5���a41��Wd)yWY%n�`�)��U��ªz�E�l�^�kP�����˲���[�kU�1�Fn�T�#yVle0�(̱�7*ع��x��w^n=36B��:��tY#5�Hi� �%GJ�8�
�m�ˍ;@̏m�QM��Q��w��$s^N;�����%;�I�E�G�ҩ4��a
֣{ki`��N%R.�2��T{wB��*�t�A����f�-���S��q�k��`'uڼ�ʺr��e��	 $x�(a����.�;[Kr�q�m]�
*}&Q�4�Vs�/N�`�bu��⛘����a�a�EJ�7g�r٦uY��k$���h�[̺�/�{�b�N`BQu��p���nK���bݐTӮI#z:1�R�kZ��3Mӻ�"�M�$�Ś�ci�œdlD-�V�,f�R/c4��6M�Y���"�-���eMW�����GR���`��,��ͫ�̅BU�Q¥��z2��k�e��TR��Z�TM1ʷ�q�j$ޓq�2֚j�IWW�$b����e'�[B�FX��KB'x# 圶t��e�w욡��4���("�w[�P���(5���M�<"肕i��UC2�sSћ)��J��W�ʼ��(H�WV {��Q�*$���6-%Vw3J&-���N�x���[�cO.��D-4@
�&�.�,�7wI�]	tYo7���%����%K9C�I��%�W��F7��tQ�D�21�b+�K�!LIp�ɖ�/7f��F�q�a�6*���ݪ���Q��CT��<8���b��tr�=7���3SdrꖝHəD?)jS��^Qa@�:��En�6�no`N�Z��m�^�{37w/Ze�*ȓ�e� n�h�I[��嵛�ո��iȢe��y6�*�1B�/���C1��^l�N�;�vLyv��3���Ƹ���fZ�)�2���c��m�2)��hܩW`�P\���t[d�u�ٵ��Xά�-HFY^�[Q����YQLhE7#�FL�Gqǖ���D��Z`ۻ�ӂ�[a�&CC��҄2��8�X�N�[^�U*�,���M��T�l2.�t
�ɔ��bL�j��
<�PJ��ɖ�i���6��A\��]��L�+(�XӍ�P�E�bJsT-��ͫ�F-;+D-KU# �T�'.�
-7++59�%Gd�fކv���;/@HͼFKܼF�l��`w�r�:G"��ۇu՛�f����� �Dm�B���Ma�)����V)�Z�e���1�y��u�ܳ�7��z�K7�kLY����h)b�y�˘���V��n%�gZR���kT&e&�fSr����7Q�E9藊8�Җ>��əbM�f�����8E<�NR�tF:$}`֨����,F[W�jm^���D�jJ2����ʰm�-nP)äj�}e��Z�����I�{�8/V������9el%�K%�47h�+��#��K������"C#ƞ��3�L����{��Ƶ�3 �X2")�%PXM�N�;K,1-�M*\�y�ǹ���dUj��^����.��^��܌�%:���KS�BY�o*݅7���FV�j��,�c/%��P%R:ģ�#y����,�M�#1����GEc2�qme����E̢�=�4t�f�j���Lr�T���8�M@2L���R����*k���I���GOr��fާ�NVd+a%ǃYF��7F�U*%�r��5݇���V�vѢ�]f,��ԑ��/AVU����I����5�a�a��Ǜ�&'�dգ�Yb�7�v��9�_-6���ƞ8�J�5Z�LC�{��L�cr;���KPd�Y"�(�j��S6���w
1	��E�����VB�<ֳwu�Ml�B�n6�t��n�%���-���N�15��=��3#f(����&��^��]���״�b�qj����i��g��L��e���E��k)�of�z3$���nڈ��m�~YxZ6��VU��CP�!����z�B�&���-�$�Rl#HQn���P7�(���F�Σ���-�,őJӒi6���)�HV��ww5X+(�o5�x/��F�S��4�	Y4�H�ʋ�[��W3Ya��52�D�S&�d�!զ�a��L"�B�9%�wO[�'�{.�a�%�u��u��2����ˇBQ�E�V�J��n%(�mF���)b�VvZ�=����� Pj����V�)y.������yA��x!�X�����-[UH�����B��$���J��'�Q�n��2�����4)~�F�nJ��� 8m���~u�q�Ah@E�o]i��F8j\�f��7nMM�`�D��\���ݺP��Ԡ����SP7!��TP�.�\E%.CtN����op"&����R'o-`�V
q,n����%�Ɇ����Ż����T��E���D7�!��#w�)��V�I(5�ث3������#E�
;n�l˺�J�Y�*�`a�H�V+&F8.��n��z�0��Mآ�m�%��aq*"��)'�(fdBԭ�9�6�w/%�ܣP1��%�Q	]���f黦\	�ٳo4<�����I1p�l'Wu�+���-�(�i7��"1:�2�ӳp��sk>n��(&EJƳC��&�ԭ��f�WJ����Oe7x������2	Ś�8i��رf�m�h��X[oMS1E�b�̧��ل�7!ϖ^J�x^$�1UL��.fޫbY�&�˨.6��	���O,
8��쩃bH�74)QJ6�^Z��˸ZɎ��ǓM��6�л;$��*�Ff�q�,]�{�\d�DX�.���6e����`���^�Ԟf���a�����F�"1Y�K�c�6O�^U�gr��RU����t�7�,zr�]�2����mnR2&�m�7KJ�mf�S��2�E���k;��T h]�jv���g��861G]��	��r���{x�wk`�,Ɍ;R�,r��'�L�iB�y�m�Z*��4e1Jc��f���1KR�&�`��A5P�֦QYkJ�q&�9���{�K�z5ʺf��a�#�A��6ET/k~ʠ����j�n���͐�
�nP0l�ۚ��C2��3<��a*≇���1�;��xZD��F/�]D�uB]%Q��+ucÃ6�:p\l������V��0�ZN��aU1��	6�d�4
��*$� j����
���h][���[��s�q��5�(�gN��L���I,r֠��Ш��f��R
h=m�E��׮�`��=jf`��˺:�D��j�j1��e�E�����U�9��T0�.�h��҇�qYTE�kT�A����U�1�E[.�dl3Z�&���oab��{A�qԹE�
�B05�*}r"�+wḶ�v0Y�)eK��Q'r��e*@�,Sۢ��u����Z4L�9��{6�T�)Z�Qy+f��pLVs�!��hz@$ٕb�f�m��0,�3�͠�ǗF�ҫE�'!���-]ٻO3w�լ�pqr�%CR�e�Y�&J�B��{C��n�(��Q�f�̂�LjA)Ve�	�)^Ēa���r��C��h�*�)�2,��vH��b���j,�S�I݉��hz����*�6:n\5�li���4^n	{R^�y�M���=A`K]�-�"�Ä�W
���dZ��Y��"�D���FPZUĆJ�su)�Mj�=��R`iH^k_3��&�SLb0.�M�+,�7+u=́�E�8�D�֔tNFPXl��9E�s7 oC�R��%S0ږ6қ����7uI��!U�)�@&��B�7o"@�&�Ձ���U��(�����얢��&L�G&�{�����aYheؼ-a{�]�ڡ,=Yp�X5lʷ��W�&�$@�2uu�*�c��ǧͽ�Z���2d<L�w[�Ŧ�qֹ���U�j�V����caY��:�6��4i�J�%�;��ۘ¯	T^P@��+��fKͫY��e
qѥ��[�EC���Od�&[�"W�G;��f���N�a��R���T��C"���~
`��GK�
�Dژ3)݃�4�S��V�Vv&2�hV�aޔ�SQ���Y[zT��S.��WXi<����wR�L��/���J��hb�����ز�V�k.Ŋ�+~��Cj��\=���29��0�N�U��.�nPŕg�!5ʁk��u��`W�rd,�݁�͵���0��J,l�®�?;�.���^�	�M����܂2�6��1"v�*�Ebyu2��=���g��P������nK��+�X�%�͑f"���GubFp�uP��[�(:���<����Uד=A�~��sэ�m$R�sa��r�8��C��]9�֝)�Y�-�����NaH�7�{�������udc17f,ڢ�7@��v�@;зB��"����'j1�qL�e��u��3BU�YJ����,Л*٣���QB�+(6��\ʔNId˔��4 �m�f�B.� ���IT�h��a�����"��mm4�ޘ���,޺�f��.ne��5�,�#��5ȝb�(�p%��-���.�f�`��V���L{��-^e��I�6���Xe��J{�%*6t��*�0t
,k>�E��neb��ܥ�Ej:B�L��V�"��1�xCSM�N\ghDLY{a��K5N)�RiF����&���z�(bT�6F�[=/s|���2E�V��.�n�ڈP/�t6R�FL���~"���1l"j 
!��wwUʷc�w@��JA24�4"k`P�X�!X�VG/h�Ajn��he=;b���n��Q2��,6�e�wKKA���钋vsvFm=�4���v�*Rm/,tN�u#��x�n�5B�ҫ��U%�Qi$�]J[�jӽC�LI�V�\qv���M��x޼�Œ�s�A��19���(7t�$��~UM�e�5R���w��jl@]��l6��Y�J,�Pc����Z�4=��r�޲̥��Q�&�u&�L2�F�Al���+)���X�.,J$�7yd^ڶ��A����4�(��64�үXǫe��O{��7k�V�T"k]�X���.0��U��w�!8��(�Z<�&�pe={�H:Clo���c@( �|���q�--�5e5����.���޹��v�Y��3Dl�VaV�p��{�/��}k��G)p-^v�r೿^O��˹YÊ8Q�r��q��u�]���lCL���y���̼3��ˊ[���]U@���1���a��̃��q�6��046��*�|Iܶ���BTqh���ܦP�X���K;E_>���z�Z�@̚�rӾS!Kۦ7�m�����S.�M
=�H4' �[��1N��wH�_�gM���9�c��X����ɮ�Ǆ;���k�-k3U��sT�Y7QQ�J4i����չW�9t�:(]
l=i���^L�j��2S�^��Y璷Qb:� J�"���$|��9���X�g��9��(K"�	��]�P���Ul�g`�Ӷ*YM.�(d�j�̮a�Pn��o�����9c�C�zT�Y\��
e��;���^�^P%4��/�rZ�	#��nlVtT7�%��Y��e�ԫf��{�xD{���Q�76��PDZx+�������c��Z��H�r�iR8���M*�u]�f��R�7Z3M�����^S�E}}x؁�6�WC��zr���]��HYX�oN�D]�J��R� �Q���U��]��i�76m*	������zD��l�,X�Ln�����8��ɰ�VX��]y'rK��8\$
�Gi!��c3�Ϫ�\��.A�(嵭MG6^�'x8�ӱH$Є�D�K#nU��k*�	��Dt*����͵��q6� ��Cf㶩�Wq��{t딇[gVG����V�x�>�Yt4�I���%@z��v6�YY������wR��m������C{?@����W�ߌ;�}�QWk��m:��hV�ꋹfvV���78�Ks�UN�gQ�\K��G��N#ϵ��;V�Qq�i�+dޢ\���ˍ:���d���Uv�}���<�.}�U�WD�q=W�<bCh���\��`��U��kS�~��gb��i�t�+�j͑Uƃ�*��0Ө2Θ�*ōMA����9�.^mkO���1�#��Ln!�ݛ�5c�\�q��є�6řn���v��9�X����h���څ��c.��fr'3mt�`�Vm
��/���~Ȅ�D�Gn��c2�hmx,N��_2�޸B쇘@����_$�����,�ɛ���=���&��x�A>Zhึfh��n�-e0�Y�$nɕn��:k�������2��=�r�μ�S��Kg�\9|�n��R��pm�tf��ug	�dz�˻A��N�����l��f�Т��/�lUt"�`t�d��ON���h�f�ܰby}jyfJ*��K׻ڌH�V����Kv�r����"|Q7��i\r*p��V;�go-�LW)]$�9�>��];����z��uaMJ�P�F��S�X�\B�$ѝ��Ew]�vl���8lR#��䯨�ŏ^�i�j��x��-8�W:֙�"r����h]]�v{�b�k���(ЇZ�bj��'9&5w?����B��_¶=���<�uR�G�n���y���|�!Ѕ5�^1���|n�����{]��J}c��ݬi#��Y�՝F�:ҧ ��Z��Ҍ�;�6ldܼ�	�NnvU��V�!����kL��m4�����ػ�ۡ��P>�J뮗v:Eښ>42�DVjc5�aR��Oa��%q\�c�p�]	�D=������r�:���z!���v����v+P�[v����|�|�*�٦)wPov���u|��/��O�l��ws[��qB(X���)+��������;�3�8���A�֙�;)�F���6���	
��}���ّSe�!����o��*�n�ݱ��M:�n�w;I�׷Y�nGzl�M�J�6L��f%�)U�f�u�lFǜ�Un�qܖ*M�wf�*s�!a�LK��]�m���eڥ��=V��tR��6K������E�Ұ̤�8S�ú䭶1Q����lLإ�
��V5w
V*�DoX�&>�%��f��lF&�/�6r�����Wc�c95�:Zى>�1n_{m�v�d8E{�UI�;eg	��0g,����{�|A�ۑ���-��3],��40bV�db��a�6a��R��Cc;&�;;��� Դ��O8�y�R)��Ӿ���;(S���#� �*
�#1��8�/nt���1�KI�Xa��u�]��]�E�읹ˮ��'bþ�nt��nv�w�F�w[�"EKh+l�b���p�}�fu�uYo�zl��}��q����v�:k���_gm�e�w���A�S?��yN��i�ck�[��]��8������Ul}dR4��Q ����9;-����GG�J�ȁ�%�>S�z�z�O�ϩu"�Qe�Ц��d��ݙ��g^hT�ґ�:ӹQ��j�b6&t�H��[7�$����m��9ۑ���k3�Hr�e���n�6��.�a7�8��!�n2�h�z�]u��sNj�֣�j�x:�T��皓j�Fv����U	�/�P�]5Z̆�ҏ)R���ԶY���)YzX��f�X/���q�X�Ōw�\���[ڃ����:���D�������﮲��i�z�搆��&%d�R�vo!�_b�<6V)~B�Mv_.��C�̚��{rVշ ̎�3��gIu�W9}��X/��^�zK��r����Φ��w��nQ���Ԥ9���˒G����V0:��Xr���^SO����R�7�P0�Zz�j�rr0�z�2W99f$豈a�S�������e�(��$��S��=dt�<��i��*����n�w.��L5t1�m�d��R{3:�*h�vOu(*�(�X�$�O6\#;λ��Δ����5Č(��Z�`+����j�,֍ɻۮ�W����7Ru�G9b�U�r��qL�C;71�i���U�ͼս&v��o}ƛ��fR��P�v���eWLx��fL���뽫y���DL�]C�u=�'+�[�`�ss��W����/�X7No�k/����F�}3g�]�������jd.Wiugz�'%�\���K�[�����`�8'�U���gg����J�,��o�j[#M�����ZC&���r3G@t�;�����#7l���t����6fr�f^���+'Q]F7\v��ٓq�N�S�L��x�
�5u(�v1��,g,<�N��H��էr�:�-����bL�Ǜ�)S�-���O"��3.BTD����Giꁽ|r�Ǻ��<�9��ɣ�J(�_sن�YyY�~%X{z0�E��V�K��_t�@T���]�TN�m_?�ww 5��,��;�XﺶAL�����9W.���l֣m�\�)�ƙ8c�h��R��E��e�����zh�.³�ҡ.�Qf����EBM&�ݚ�ja»!������I�C6Z;���8	}r�;z�f�亣�˻*H�m��.�.�|��U����lք�X)��MK�z*�#*p�$_cچ�C{��;xv�69���9�6�v:�]l��X�MR2걋.�;�lGy�=��-�
m��,�Ħ��9f�<��1��;�2�I�A������m<{w|)[C��3�!A��kz��k��um�ct�Wm"���=FLɃ������1Y�D��/l��#��((D"�X-_0>A�� ��CG �ݗ�9[I�$%[��_ɘ�u�	��L4��w��P|��ǋ�jn+�Z���\΅5�Ws�f�P�929&�UY��s��_Q���LT��oC32���q�G�kjW��r+Y��GG�!ɸo���vm��p���[Q��k/x#A����[*��Yү��V���n�: @8p��:v�2'�F��;���p�%�z6vp斣�[0/{X��_�8|���楃��=���pj�J���3q�Ý��J�f� rqq�y|�#[�U�u����J.��'�V��f�vZ]yLQ-���/.�n�Ժ8{���C|Xk7���:��{wo;���e��LcOd��p.�9S��ƓB�=V_j��͞:xʴXXR��/Ss�(�7��h-����8����G �ߧ�+�{������2��ݞH���~�Ձ�ݮgR��H&LӘ�!�(���P���b�Ov��v�d�c�+�ɛǖl�QL#xmgwf��|�s����wEղZ++�n�xPh�v�v�Jُ��5�����ZMANv搬�C���_=OV`�qW0������=�yt�Z���)k�5-�e
��w��k;oGH$si.��E�׺9��B���4A���o���;�X�+�ٚ�[D���qg]���9��_u��E���e]�9���7kR��tvG�(�eC�՗kL�m�^����+O�ZaA��+T�,n���Vk��CH�x6�|� ���%<��<:��'f���+� ����U�J�Vt���rw�L�fC����.n�\�*_dޏ��D��;�F��}т�"�T����暹�	�ϻ�dڮ��ffY/w��cn���x�jɁ���N�'��2ҙ%��t4�xARcÈ�ØWW�����v��f���p�N�D2N��O�#1"��SG�Wo�q�I'��܂�n��+z�ڀ�><��)t���0�#[7Z�|נ�<��k���ZΌ�������|�֑ո>{�@��#`�x��ȂUa�W�ET��D�\�n����V��v��Z�LH�������u���h��۬����t��u��3�Bmvmј���g)]�\�.�%��U�`�)���v����A\=�:�D�
�su_v��к���}/�}�6g19��}[2��i���ǜ��4mM�����KE�m�Ჷ�3��1�j��ʫ�<]\r^�4���;�t�7��@�u�Os����3�^K��+�2����ܽ3�ѭ YS7�0.���n��.�]��J���-�zR��:(�-$3�����P�c�-��5gKb����{s>�oȵ,+��5��9A���l�x���\�n�N��d	E�e�1�[�
�x���b�+��vJ�lS��0����h���t|�L��NUܗS[�e��w���f�>3tB k|7:���ۻ�"�e�X�o�#v���:̘����k�`r���(�Wi�5&7C�=˨�ڏl�V�j�f�wk2M����
�uI2�DG*�V�#��4�^L��7��N˱����O>��I�V1��o8��;F̆�Х�7�z�o�uW4���v�|���b4��lgM3����E��=��ʡ06k��FO�����I���g�ɵ�[W8�N�oZrH-��%N݉kv�\��r��A]�j�KY������]���v�!���^��m�p{������r�/�/3X��Cq�=�3i��<�[mg.r�j���G2�z��
�:��7���g	#)ԷN���{�N˿�[�+/+�J�����@u�Xy�\Y1$%�I���T��c���U�y�9^Io\A.��)�S�~��'e��/�=�Ao)��I�H��n[J*ݲ;�Y��p��3� he��wh<fLIQqǖx�N��'I�󕶗f���C9��s��(]�@�w \�g�����0j�w�ꡗ���K�ʍ����HnIoV�ՠr�Q�]�Ǒ���M�����B�p�q��ʅνhWs��t�}�b_)WߵQ�z�{ϫx�pr��,���D�R�z����'��"�Mʛso��I�>��,��"��9r�lsd���gR�0n���f��+n�Ȍ4���}�X��٥�͝�l|}}�mֹ�m;V����ɕ�H�3����r��x��!ZsOǋ�ƺv���;���Y�	�wV���Wc��v��$0���0���g)�6�PD���g�X�_���ݙl��:��3�7oz�nW:+�ar[�w��C�@_gV]�����jVI�Wh<��8�QJ���I��k���P�O�4�Xu�uw|�<�d��.ӵd��Oj�u�oC��1JǏ�;�dD�4AۺWw�uT��J�2�w���,s��&�%��h�����*ǽ�K�n'+F��!*�_d��Ju?��,�^���r Y���iUށ�F����nɨ�7�����#�\o�i�K,�K�Ǎ�׽w-o����ķ�9#���w����A7*N�W�Y�m����T�ޮ��hP�U�*�ɻxt7e�|f�f��m��dU��.9i�w����;�E&�e%������wfQ�ehuQ�9�M�u��ݢ��_hM��2��R>|�����}��^��6�ݗ�b�R��8���X"�nf�㳖m[̴����Iux��V�%z��-�otسw��v�����i�Ǆ}9�vk����X�L�����+Uɽ�o.����Ԭ ���;k��B�9�egt��)�7�Gwn�TW\���n)Ւ�����D�s7!������-F
rucP��2�����˽
Q��4���K\ը�C��69��0�si��4Lx�#�#Pʎf\t��f"T=�c{�N.��n��[��ݓXo���Q��};�M"sv!���ǲ�v訆ݴ�C}ڪ�خ�E�M@����:b�n^Rh�0��	ʹO���1ݙ�x:�����A�7Nd[G�N�U��z��6�P=���m�.Et��=��_c
o�'lp��G@<u�[S+
�\���Tuv�\����&�գ��^CI��}��j��
p2]?�h�wֻ��$�rX�s�}�Bɍ���@h>��n�1bB����TD�{�� O�|�%gF��kH7��|m���_?�{X�����Z�S9f�)�>��6���8-� -���]v}v��`�%��f�F�D��L*لZRc�7GM�Sl����1���B�rΐ���M���c�����mF�_6WO����_7u�7I�ܷ���y�����b;��r_t��N�f)�A��4��$х��Ђ�8F�O�3s̱E�ܪ��$��+*d�	�	F���$Z�nQ��n0`h�T�P��`��J7R�e�)�r�տ�%���	��I�by�ACy�*���ul�l6C
�s)� ����Ĥ��D;�UP��8؇#d���h��)@�z�b�E*�yB.y��m�yQ��q[�a�DB�IWD�}"L�b �*�P)0��	@�E0ˈBL�

ltd�Tԡ$��F�ԳA�����m;*�P��iڤ��$M�Y���$ePr��	p�B�i*i�I�I	��HH3�B��Ům��6�)F_��v���B�Pa�� �DT�� Q�EEV�ʸL~��DҎT
}�("�0�*dD����p�%�^a8�&�$��P�
F�'�j�]�b�jY17a"�뒉�a�������[tH8��4J2�f��!&ڔ]�F�-�b�L��a��h�//8!�b,��dё0cD��B▼�h���&'FLV��K�f"���V'()Y�QQ��~�U@D2ߛ�츧�؈�(����xl��<���;�i�m4�E�E��[�~R#+Z)K�'��S\�Y�rl��T��ݿ<��B�Xs��2���=���}�n���{&�3�yɝ�R�Nܪ�e�q���`�(�;ǙX]�p�T��B��==���t�����t!PmN�T�6^�e=D�]x�XX{����t�4�[k�B�4$9���ۈ�l�Yr8�;r�t�m2�4Ð9gӮe�c�(��6ts˧K#F�V3;#}�QK���'z�L�2�S�ΨW��ƫ��7���
�5`��`e�����1e^�'9m��)��-�}}ǻ�������ޭ��.�:<u4�����T�\�I�K*�j�#�M�(a}sn��yW��pn��C@���i���X;�b>�c����.Ӄ�N 0��0m,u,����>�G^1aQ�^ҸZ�_R�΀E#	�p���T�Sn�=�������}��s�����H>)�*8�k��雷ݝ�[\�e���iF8�B�M�|�^�QR)2f
��:�*�&���ϯ��颉��5�����] ���DZ=@��ӗXK�p��!�k�:��f���s3��
��|�oO\ڱת���eç0�-ĺU�nԝe��������~c|��~���}��________��}}}}}}}}__\���������������������������������������ϯ����������������>����������}}}}|}}}}}|}}}}}~>�����������>������������>������____���ϯ����������������>������������?������?ϯ�����������������wƨ�Q�H�=W�_hfj{2�	�����g��*�<�s�Kv�s�k���ӅRޅ؉��z�?,ɕ�X��}�c	���3��eq�����o�Ь�meI2�wܳ����
u��6EBs�D��K5>�^<�2�2���� Ws8ͭ�bl�3[�4R��F���T��E��%vh���s�G�q��ۖ9�UB���!������� � H!�y�a�{�Y�ַk�Wz�Ro3tZ\:��Hu��^���i��Zt�5�m�����-(s�v������n�UMvք��rr���L�Ԟ�d@���]o<}���p�'(��
5t+ck�f"��a��#��X��e=e<�����N��@�Z�qv�U:��lcw�}���yY*�h�-�4�-��M75�6�:f���cٙM��
z�b[�n����&8�Ƿ�Ȫ�f�@�]I7e�B�x�.�Fe�Q���>�\uڤ��:s�M�u���M�?N�叓�oa���c7�b�����&��`�ve�jXp.B";�Ė�c+�1�݂�u��r��Y�ݥ[J��8��o��p��c� +���|�o]��Q�s�-c,��[?M�VW]�(�#�;�wm��m�X��C�u�N������:�t��� �ޯOg����y�������������������>������������>�����������}}}}}}}__^}}}}|}~>��������g������������������}g�����������ϯ����������ϯ���������������������}}p������������}}g����������}}}|}}}������?�����}}}}|}}}s�����{����@*�>��+:�{��8��O���ҐÛo�M���[-d̚�}_v+��,�}��6*n���BE���͈�;6��U��*�f�7!ζa�����<����E/W['x�C�o^�M��.�h��T�=���y�K��z�ӯE�(����=������*Vókxc���B�:��b]ųu)�O���ĭ1�P��+�\������+-RI�zz�afXqOt'!o���Ǵ��thwT���p4zyFAx:�;7�����t�vu�����c珵����K������ւ.�j�C�|�)՗���G^�#!����5ޜP��H�Le�d�ݘ�� 
 �A!ԫu湝��ٮ�`�	'U%7���J�^�Sq�ʙ�6��(/ZbM�kKLN��`:������%��-0!�xZ�䥡tiJ ��ʧ�2�RX�w�<�4�k$��rГ�J��X�ӷ[�E�s/��֖������e24>c���\�xK̗Ġ&nb)�X��ůBW���u<t�Pr��ꆶ��N�]��vx����8�̻/��d+���gu�ػ�J�!���@,���1�/�����koM3Y�Wp�������]�"��6��h�B�-�F9@�o6Q�ʭ���t���Y1�Y}Nd�����$<I�ݵ�>�&��nf����.�|��������w��������ϯ��������������ן______���}}}}}}}}�G������������________���>��<�������>�����������}}g����������}}}}}}}s����������������>�����������>����������������ן______���}}}}}���������������ϯ������}�w����e��J�+/s�I@A�(��+,!���dq��;s�S����*EC���i���b���YR�},=<�r{x76����vc�m7�Z��-����*5kRT�\�)=��B]�$x҆��#��y&�u�x�U1Rn�v�p���t�kZR�N�:3e]�n`������ToZ&�he3��u��uJt�˴�3ݚ�T:�P�����-�~��x[+��p	�_u��t�k	��+"���3�p�=��Jq��"�*�f+�YCq�}j��A��L��muY�6�,]77M,Fu��6́�P&� ��ɪܴ�B��Y���'/��E�9m�z�Rgk!<��c�N�ym+��u�vP4�{��ׁ;.����m7��.�����ux���i�d +�r�jl�Lu�e:��f�od\tX��684�����Ij���d5�o^�w޳��\j��\��op�����Un�}z˷����b�J�VBGt�[H]�J��Y���|k`<��Q��_3t��EGE���,��]��S�n;�<�V�կa+:�yg��=��4�H&b]�=�A��ʌҽ�<�@�fXn�(�F^k�0�d[an��g���;P��6�mAj�Bv��qYk���u��{��B^G�k�+�,vY�n]7.�˵�eJ0��u�ڮ������
�&�X�.�q���MNͯ��C;���I�d��u36�-5�Ė�=+.ǅܳ�fc�Ȯ�W:�w�H�vՆ@7�|��'w�x]�\�p���F��Y�Uon�Z�o(}��Z'�q���$�9h��ȷ�~���U���/&����o>����n.�÷d���#֚�]��!7ce�̪��Wa#X�,V������5���`�mwx��sB�����*��M��$��v�c;/�h4�##�V�:��n���G�zlA:b}Z#����GUwT�˸l�q[�E�7E�ְ�����+;E{��웪�d>縺�^�Q�Y�k7ښ�:{ %����8�R֞�}�_.Pʽ�M2���%���ӑ
��f,�3-c�+��t����;�^*��W�|Et|���Q뻛�N������n7�8N�8B����t(ɕ/w\y���f��o4=�ɩ�.�9yw^��ʃ9�C)����7SYtx�4v��ohwu��o6��3V��5�����2��d/��u��s5�+rV��բ�;��,��*�CP����,-V�l��b�2�ry���7V�zs�l��v���U5Xk��,}3�z�r �8b�@�Շ��B�����-�41r�[n�2]Ț�7۵a�[�#������׌�����@�Y����.N��be�w�F�-0UԪ\Xv�}|W4W]nZ.ZP�7�[P�F�)y�~�[b /Dۮ7��7����m��}W[c�Ż�+��j�7ʦJn��=ϧ�&k�������*ѥɐ6�=���ð3H�D�1�6*�ukj8��UF�f=��4���̲wmV�ӈP�9QI���膃�U^�룼8�50V��L���y�3�K=J#mh�@XU`�)Ӧ�ފ1�,�l�ɬy���u���9��]��y4�;��v}T��i��Eݜ�邒;}7G4�S�F[�NBX��Aw��Ϋ���v��؍|�a�:#�du�(��w_K8�fF�i8���9������#Gog�N�aC�Yr�(R7��5�Tۄ�,�!3_xK���*S�� �n
&JB��æ�V&�o*L�L�S����у�Tyu��3gp��;U%�޾N���/��bhq��\��vX/��R��/�>�w�av����B�!gE4���vqJ�|�]:�O1a�ά�H��b����9n�"��9d���iQ�3�GQ��[2��۶^��]xIWgV¶��x'X�BZv싓{��J��{�Ͼ�0fא�t�8&/Ml"�:"��5�l��|�9b
�Xn�r�=¯��	6ͦ�W�.�9��n����-Y(Ell���Ysl�ЍM����)��CNw!S�;��q�U�,��l�%���c<��Z1g�Y�$��Uj����6�]�* �J,T�#�	�����jgjMj�]dE�4�x;���E�X�{�1枮�3������(v��Y�I�7A�J٫oIg�Y�Yp���ht"����8/>5D8y��u��[:aR�L�;4Rh;xl��T���=j���*'vgp2����	�����������V7���u�o),}�}i�8g+�_C*���$��]3�4����MC���Gr�Q^n��_gP)`D5�@nB�����rk)�7^��v:v:�c um-ᬄ^�'s�+e�a˭�r��;��*@W`=2�Wd�s���t��W] Z��V�#G�yu���\�c�BW���ŦoS6Ladk�9֙lvՕ�ή�[���s���meh�5���u���6_N�C�(A�Z3��6E���[YB�^䓂�ǉ���n��,�'۸M�Q�h����a/f0�u���,�綹����*V��濔O:��ǂ�r�	7!s)h�԰ĕ8Q�T����O6�U��D=�����p�ҎQ��]Ɗ
����k����D�c�"�c���ˣ�%:Թ��fcx����$�
A:�m�4(�Iqmc
���͔�fU���N��z�8�Q�wQB	�$��\x�L��k{�{{���T��^�@�m�a:�e۝��:3�;o�7ѱ�m��$݄9�
��Za�r�;�9NZ
liI�y�(9�6,7ck^�G!�����ں4x�-bF�)]E$6���t��u^�B� k{7�FH�K��F�O\��׺9XW���!ǵ������I��C�a�Ƀaۓ�g�#�M��=G+#�+B���z�H�Պ�����M�9:f���:�����5n��af�e�k�2r�l��38_�rl�,����������E
W%����w�����b�7�S�1����� �8��Д�FZ�~�F ²�p��V?��i�٘��/��|�������2����	_oܕ�_3U��Uյb��!�gW]���2�oosB��Ƶa*K��<��O)�__L3�f�E_t�7*��-�[fɶ
	�`IRve�=�۹��v�qQ�#���eb���4���vD�9�c���T���mԭ3t��|��F��f��^�����\��϶=�H��ξ�������4��>���9Έ;�ò�N�,��V�L�l]���6�ٜ�A���:�|;R��(1<�����Y@�G�T����� ];�@��y1�0T�i�[vfa��$D�^`�#�m}H-�4�]��(��R�5�af�#TV��af��+�]���aU� ��t]�ˇ8Si��`�Gj&7l�3�U���e����Wu>�6�"cʃ�JlGh����,v��.��wy���ٌ�uXZ='.ya)E�T,^���-v�ʂ�����j�^u���'L`�4�ϔ��V��W�m���kk(��>xM���Q��Ө�[(�f��g�tm�WufFiUQ�5١+{�w@/�>�@�
�+l��K���U�v��h�M-�"K�/(*����:��ݶ���iZ��Hαv�+X���}�ҨGTk՗�V@�Ha٭Y|��e_:�ڝx6���PƬ��3z���H�Yܰ�T�oHٳ�{�J�m����7o:��U�NKqU��ú��X���Ԓ̏vb|a��s����r�;�i�f.��;;��6�-�L����kGM�(�t����1��|���}a�N*=1b�-�9JJ��]i�<�)L�츪rbl(��n��m�
�	L�e� ױ=������t�խ���|���0�N:AKٶ.moLk��z���*�ܤ����Po� �[�ޭo����e+Y�H�V�au/ 6�����I���`����'t<�W�؈��ov�[P�@�2�/&L�z��pA�^?�e���f�
�����5�Zn��7	l���:�*{��=,eoz�;9�]p@�MP��� 
�n��ͧlPPCsK�s���ϕ%wqbf�syp9�Aݩμj��dFIc�yb�z��"И�t��\]f�H\�̓E ��y�$iYN��B�*���|�}��Y�ʤ�Z�!�:�ꮡ��Yww�}x9�!�9w!�TM�?Jh==�g(��&���f�\�E��͸,�(�RY��n����w5+��r�Vb�0ٳ3��)dv�Aa�::4��۽�+�PD�s�Y��A'u���!�C�;�Z�wo��ͧ@�G��G�`��`���Qg<�c/AXd\�ݕ�	Z�h�f'���*qƫ���=�8�Yм����.�s��X|��8^�A,C��h3e�r�uHދ.!��k=��Zf�\�+T�;U� ��}�$ƮQp�̸�edfcÝvsm���S�nQ�*���G0{�5hc�_H�X�w�pn��]o.�Q�^q��<�(�ñ<��^����������t�P^s윯�L�δ�E�R����5�b?g��ڨ�*�����~}˫�y��44�� �"�B���p�3���m
>���E�<�./��p�vL% �a_ڡ���D��O��6����w������b�P˱t��2�V.TǑ@����8sZ�y�Mn쫧o&Y�$+c�Z�����;����/۳�[z����BɅ�$ѹ3N\`����ӭT{��	3��<r�X�չ�ʬٔ�ķi�+z��\p�/u��=(�yd�[����o����W˭uF��6�'x���+��폟�F�:#h�fqydP�HjȞ� ���%�5;3J��5t��qX$�o��I��ZQ�+2��]ϊ���4�㓷;��aS�{|Yʉ;�Ѷ	�����aU��L
E��3[��a��r�������0ge�#��x����wr��U�%��kۺ�@Ъ��lv�J��Z��.��L��������(OY�l�������%�5�eR�Ձi�{z�Ɓ����j��8d��n�IW��v�D�F�h���{hN�ק8H*��绪�=��P����F�d��ã�.\Á���u�1Ҵ���dyE�I=L��;1nb�e#Z���ALV[����������:�Z��}8�
6��1�1a�4�p��o-�������0+w�U�'�J+�'.�������m(HcMWr�҉!�ѩ!�j"�􌛧(�f�A���#L2Ld�|�)$�1(�8m[()U\���*
ATm��^4�%�I�Q��M��HAC�h��\Ll��J"��~mD](������T�Oo_��y��}~>>>>?���>�9��/�T���+�j��J�ڡ�#��E��DD�@U�;4xv��$?_Ϗ�������������3��阊��	��"��((���q�mx97y�N�11u�)�"���EWmM>��>?_�������?���3���~�`�3P�vB�"�`�QO��W�"�jb���	5�'��V��������qɺ:���p���p1���ZcgU���Q�8�+U�j"�*�t��D�:ѱ��rV�ꮵѨX��(��j�3mV�kFƭ)�#�ت,V��m��O��j�
�6]���SV���V6-�j�M!2Ia�㐃mE2�m���h�ó� �]h�ڬO^y���~^OMA_0d��9�뢹#j#JN�)�3�`�gj�[����r �0�B#��B�gO���]��Zb�{�F�^x��:c��wc�/���AF�v���"�1�"��Wn�Qu����m���&�6u���ڈ�����SAE$TPE^A�����k͔��t�GI��+̓o�M$l�f;�(6�W����X�������u��neu�sQ�tM\y�|�qS��B��G���������C�7-7	�J���e�`�#EH)�
����>S��ʢi-�����w�Y�M�Ot&�Z���ۏ���;������>�0&{�G���^{p�����f͸��`�t��\C��	����=�X�3�dv�t���N�Q�b���'���3�K>�,Z �}�<�H;�ov��=ۼB��VD��۫=ܖԄ"���h|���R���s��gb)��h����20�m��w���A2sl����M��"8�Lp�W������tI'b��5wl�ޡ�'hao������׽UB�:��d~��W\-�8��&Ƀ�0+��x�w����\�Ԡ�ɩ瓮r]ߙʋ�7�m��_�j�V@�rLT};k��zO4=�K�O���.�m��qu9����t�[-�.���3��D��z�׾�\��'
��=?r��𭺝��;���s�=ySݻ7b�����7#���`��9��2}l���9s&Z7��G| ��[�wO�����W)�*5�oFM�#�eL[W1�)K�QȚ,gJ�l�[�h_�rE3�_I�S��Jz���n�{{9�þw�h�:�,@�w�ʋ�y���<�x�LL�*OR��o������ ؗrw��^��,��}}b�m�y1-]>���o�7c��m���؞�\}��7��Z w�����f���s�~C³d.���i�ޯf6��۝�;�Z���_ڇ�o���35/ӻ6�t>{|V&߂� n�g�Tm^�*�0ި��ZZ(��j��i�Sz��������6l%|��o��i�e�pɳ�K����{z����!.W��2Uʨ�y}�}�>�� PDS@r����ճ�>̟17!�jD�<+��S��;ղ�����x�Eˇ��f��b�woͯLc%C~$��xUޫ�������Q�u�E�{�ե;��8��d�k��ڻ���x��]��}�U�f��'Gg���>���3��&���Y&�3z��U�,�r_��)�=f�\�Kwʃ�Ci�p3>�b鏄�=_[Ss����ϊ6~��۽f��g�r�gUe>��Lu�N7�3����#o'^1y�pA�rF��+�.ڙܝb��_e^�M �Nt᛽�j�KV%a��î�n��P&�v�n�>��#zܝ�D�3��
��Z���οosA��w�x���H[;Za�%�/G[ �������N`N�Ei�7��}9A�.a�Xe�����������vU�>L|3�z�-���#�>�ؙ��'��OO������w��=��� a��Z����оx=9-��Mk:O����.�}���V����V֞`��DQ
�WӯM�}�o�-X�mi	��gF����1bs��f�w��{R�qA�N��__z������/��Ξ.y/�r=�痟^Q��p���s�=@���t������[�m�|�a�OM�zE�������6�x�Ov�կ���\Rs;��J£�9��<��"V.S��Cb8�잣�-��c���rK?T������M\�9�7�uf� �Vj&�b=q�v���o��8|������P��e壆`t�ՊНG{��A5m��ޫ�GWw)�,WrO 0^٤�u�FK낉�����oV}���Z��Gq�闄9���.�r5�B��Apr�7}XM��c�V<�T~�vr���X�D������})<�V��\������}½��=�=���7h(�����o���7L��L�r\׶�F�jOP''(i�9VM�JI_7�a�)�����Qc\���.ކE�L"-�n|)�C��\��=���y��g*g���޷c�jؗ��\tg�MW�\��_.�|�j��¯�k���_/��b���n�(�UP�6/v����y� ��W�ہ�����o*��|��>��{&����#BRt�<j=ڝ��v�6�}���n���w _�w�_����6�k<Ͻ���k��7�ʦG����A�ڰ��EY������)�f�^�5y���tv�=>�q�=s�^��50�#�tot�*��>wS�v�Qp>s�~�x��ә�p{k�Dk���(��7�ٰ�Z��a�[���>7}o7���𢡊c���O�_l;�K�uE�;�X5������j'���ʀ�{j�/�!�\�y}3fsi�N}wi� c� �G����i��
�7ug9�F�[kI��Aqǵ�S�"�Β�F�ۼ���~($��tY6�!�c=���5��2�r{5�a#V$���6�]OKv���2�i��)�S���UY��T����Y���
4��j�.(���#N�o]���ɘ�lA�!��Ń�FV�N���9����}2cX���i���a��V��CLv&�mJ~�LU� �/��Wl�3}h��+L�v��$����?SԟY�w��O�װ��_o��Ϯ�r��2G��q1�>I9O�ś����0�Vp�hG����6x0_4q�ʿq.a��j-���x��ݵ�u�<Fo��f���e����x���9�T������/WS蹘��5|�Y�M��ܹ�_֑_=�#��JJ��m0�]��m���u{}�+�羆�����B_��W#�����3�����4�v6�����5���vUI��[8y�8tsc��is�uo�ƾ��@�MYD�������[^�@��:��xUճ��>1g�X/����af}�p��W�o��W������f���5o#�Y�Ifȃ+��9�z���,�W�'je��1 n�Xq��r�^�p��]C)���XN�*ǀ�z�Y�x�p�����9��'R�����n����YD�(\�M�q�xj�$��i5;GgsZ\�ɗ�:�.�A{Z£��ݍ�k��in"�qv���Uw7�<�a����a��j9Ţ���l�|�v���'���ڙW5�t��Qg�簃×���tf}q�]�v��� i��	�Q����g�����;��gk���:��	7&`<�����19��nHm%᛺3����Nd<�q�K��C�0��"��p�;3'���~���)��2�g�s�g���D?N�n#�O��#>}p?i�.|�_#����o+E����w�¯�ל��YJ��������1����9O�{��*��B'�
����^a��{�lNuà41腠~��zv���!��_s�Q���H�}v�|�7���%X�J�9��k9�ys��d���wz�.�Yc1���\Jɔjڽ�E��:f.�����	ړ��E�>ڔw���^QH���~*ߖ}�9�3=�Z��6��N��5�o�����姖���0� ��@�����Cz�G��k�%�+Mn�����3���'��퇫å��;��Z��)n�T��H��k�oN����˸Ra��/��&��gJ]�Nw��-l/��Οw�_��E?l5�+��qoh�����Ȍ���l��}��I& &������t�<
��۫�O;Wv}&�	�����N�w���^��'O��zzg�{d��VU]���i��}�{��<͜�	�޼�[���l�VdӲ�p�=��5�n�w��{&�ɸr�����l�����5�D��H��H͑S���`0��6����y9�{}����i⽹�4������ֻo�꒜��>{��C� Ka/�l^���%���v]f�"hEV�����6dU��� ��C�ݨ�]�zy��<{�k�5>U1�����DM�,�������'���[�u7+a�UK�|���e��>���)�{X�1�������v2���9Y���l�=�K�q��=�+ܾ۫�x���Rs�X�u�����-?�����t�S.�i�غ�c̖ Mv��2z��y#r騁0�ҹ��
��(Zb(�[Y�T��eܫ�`� 1�K���rWIǒ��(f�6�7u��__t�V���rʡ��8x�:y}Ywi��o�q��:F |=�Ź���㈉"[Dz���(������|=�ON���wƭ��;ܮ֣����|���݊xWw��ؓ�g��� ����c�o�gќ��(��}���X��^���|���UN�&ڝˑ��[�mu8��u��|j��w�3���:֐#�^���'n�h��'�,B�ۏ�N�S�����{�&�Y,}�T��7��_|c���� m��N
���Q�W����'(��m��e?l'�l��}���ܙ��� �\3ԓ!�A�{���^e����J��ّ\t�̜��=7`�z�a�-�^�dP��#tk�|N����;���u�=�y͝ �͙>����S��#�܏�:��`�03�C�~�Ҫ���l�s;*���������a]�(�Ɇ��zmgT�_X��:�i�Z���Uo����k��,�w>3M\s���%}�f�y!��wV�f���V�g��KV�n.ً34]��9N�$;�%4ʭZ�i;�/.��`L�n���f"�a@�\�p��
��#z��9���k:��^��|6u�Z�^@��Ă%"00b1�#$�U���W�1 h�>���T�����$P}��ښɐ���zt�|���h��9�s=ҽo��v�a7��T	��a�`n{�q���v�(Q���憎E�~ٜ�x`����9us�}tk�Dj���^��|�ӕwgԘe�VK����?�p�n�z�i0:�8�fWu�L��|U��\�ߊ��Hϻ�`�/�t�t�3����ܶ��4m���V><����V�q�2I�8��4g��CP?V�ɹ��}�+�������ÍWG'1܍%�gx�ޝ9���t�:�o�侾�/�����/���J���6^u��;��bG��|�u>��'Sk�Q�͞��h7�oW��˯]���K��^��x>�Ϭ�_�E�f���R������������>����7��.}w�5���s`��C>�>�.5�����oBnigz��g�q����+Z����v۔UΔBJr�5�q9I�3N��L�2�q-\/��~��ܱm��w�2p���S3r=��*�Θ��Ff1E�s���IǴA9�k���,����sG<n
�������hA2��X#����[�R_}0g��T�dq���uX���샮w�=�A��S�.����{�F���ٰ�*��J��''�����{�//KP�����Mq=W�&�������'b��t�$��/�8xnX�۫�0���vk��W��S��.3�O�����5;eT��/k˜=��;�s����-��XnlY�/�-��U����d;��Gf�^�ۓ��#oꀻ�E����ǐ�4��Y�����ryO��<�����v���OW��q�����2�-����ElP���V�f$O3�h���|Of؏(�K��bNe�8�+���n���~��y�4`ora��,�+��9t�\���d�]��A��n�޸q1�7�zu��صx��u����>�{@�F�?a=�n���]�s�V��>�4L��_C����c�3����xx�/�hh���;���M�o!ߙ�"3��_[�	S�:���b�cWL�֬&�Imѻ���Ŋ�և��f��^�RL� �ڋ7� ��ջ�3�i�>�{;2ܙ��ȉj[�E&к����ko
��k��tިW!��	�Gp.�p�\+7IPÃ���A��͵���k��Q�ngW���ݤզ���5��sǟ��G�t���T�#N�l�-���i�����{u���_.���o	����;֪���GX��3��,6��L�3�r ^P��9�Z�Q�P>k���ltmm@Nm!a=�����*�j���!j�GO�gY�rsoq�Q��é^��d#r@����(��e�#W�_7sU�I�weaat��9������\�yDl��j��Ԭu�x�]m�X��i�W����d��\��+�`�tq��2��^]�#,H�(�>ݰg��7��sx��L���b���ٗAS��
�>nٸ䳃6�Q[;��]1B��z�,�~"��w��]���i�=%Ye=h_rCB�e�"0�vPzI�~�B����-�OR���}�Y�N윎�8��#��z�ٲ�vNcxh���g8��^��k��M���n����L�3��1s.�M�-�h�%�c'�[T��R�A9Z��țo���ᨫ�e�k��0�"b�	s���Uh�9E�A�5U�8��o�����	4������^�o&K{��<��&�:seX�0���t3t�>t�x,���.�@�?P"؉�V�\2�v�w�*��۬6���5�'n����W^t�k�����,c.2s�ܤ6_n^-95�y�����\_v�(f���c׼^�b �ժ����` @V}jV��&J�HN�<:��͊ÂM1t���mp�N�tê����ovs�{�!ʬ:q��ө�̋9r�]�Қ�ν/![0�sNh���p������*�]	r���Td�kr�.��P�.�ue���z�(Ia�N1Eeo�*�r��x��Td0�Z�����NUޖMr�����l[�Z�����գ�/�J:g1���2��3cֻ.�����1,�w>|�kи��N�XV�'�m�JRwV�����{̟m1t.���6��e*;n�^hn�;�Ƒ2��\�u�s{U1���V�D��Z�+�LC�WJCM�Ӵ��8̊�[�ZƝ��p�|C�����{�h�vS�9ʪ�x���2�Z:8�E�ʏqkt��$���K�U��|o��"��;gu�x�#�7�\��=�]������2�.��``�m����/Y(Ӯ�s�#ѴL���m��{�9��]�z�� YF*8J�ǹ��V:�w�{�����i��+Z/��楊��&���ב�(#��=��<�����|||~���?_��|}?o�{�kP%Qv�:.�?�v6$�_v:TPU��у�q�~�?���������~>>>?G���~��}�hb
(((���h���]&%h*��m�{q�o�}���D��<��tu���|y��y�~���������g?_}�&"=�5F�M_oǳ^AZ����b:tc|���ST���ƴAAIC�OT��p��PE;c�K������2R�BQG��>l7���l:�w:j���E�SvPIKN'E�l�t!�yڂ��J��U41U%E5�vbh��i�)IM�4�n��	� �^Y�v�K��i�5!�3��:�ؤ�"��"�H�`�Q]yU�tT���KKAITww&���9�y)k�K�	��H�!�,e�nп��Oe�R.r0R-V8�y9ոi)��r/[`wX⢼W݉`�%<ỻBIΪ#��o ���oÞ��mM����f���27���[C�arz<,�,|�;>%�P&3��	�h�_��_��t��E�j$ϗ��z塡�z������9��#~��{���> m{�	Ć|
�N��}m� �3{�|��0�5�}�^�����N�Ce��<0]ha��3���wj܏qwh�e�e���v��P�m6\�v�;�	��>�|Zc�{���LZ1D	�o�N/u/X�m�Ҕ�@�2��C-��ݬ[j�̪=Ϫb�IO���u[�>G���]�D|'��rW���>T�b�[�x]���^@���O���M���btc�r�{����
���;�uvŲ��YD���ȳd��Ā�s��(6R:�Pb��z�ǷDh#�Łb�l�l�^�wEs�褽b��Un�aS���P͇n��@���s-{xJ2���g��R\w��z=�#�d �>_�O�ڃϞg�2�������V%���\nr�.�F	��;�s�V� �AM }��� �[B�|�����ѝ#���GI��j���P��2�w톗 �
*�G҇����*��H����Ѿ����:�G��C�x�Z�ƻ���>.�M��x{�[	��w�r��
�>U�bU�����vK�P7-�O�����zm��_=�@��9F�:w;�~Cg��:ݬ+۹?{�8�2�ϯ�S^��N�ni��7}iv-!�g����ҵ��*T�2�+�Y�����hqv�����#�Q��_:���y����=è����j�d��lr�Tbx���5�q�~~>�>�e�r�Gs��o6��[�=�!�!�V*!fFJ��Cn9cŠ��8��g�"%�]�|0�y��� ;��W��j������雾_��i��=�#IB���Y��gd�	��>��ƀ�:�/��fl~w�f�k�9��B�����������K�&(c�{�z�=ᵏ�S�i�������j��|�XwL�Zl��vXA��+.���Ʌ�L�[��.�ذ��Hn�ZǱ��{dk@}7^9�>�o1\4�$tK5�Q�=[�z]��xU�ՠ>-,��Y#�T�"ھ^�����X�Q(��̞y�P;]��Bem�Ҹ�$��f��2��j]�ʇ(|���&&��?~�� q����������\c�c���}���׃�+$��x��	��h��X��2(�oy䙷u�����ّtǱ�xi��Po+�`�5wˣ�$��K�=��Y���n����1�uE��#6�v����j zኑN�於�Y���U���noqK��g�-E���B�^�� q��R}K'�sG*��5t��3b�ъ~���j��*�Ux w=V�ܶ0�{y%��ZRA���r6n�z�xs�wna��P̮*�+Zj�hLi�����Ȧ��&-���[�p髭n�k�juNb/�-.�}*W+��Ut���\U��O0Vܓqҭ�[㮻-b8g��	%$���>��0����|��}��Ͻ����P��?����;�^׼�����c�70	���K�ô/_��uũ�����QѸ{�"b$�dC�7�����R5t��E��MN1k؏ss3�Oh������47s�{|���}n�K�.�̯b8�ƻ6ۈl��
�g`eْh��lNu����J�nV����{�s 7���O˟�g�ș�T��j���-P	a�������ܷ�*���3��ĳ7l�Z ��D�j�P�r[�ŰlT�]���
�h��2q쨭}4������uv�T>-o`FAם�T| fi�y��@M��q@��y�����I�W?��j|cϮ�@��M=��UK�}g�dن���x`7�0���L�oۨ�@�5�T5L��5���dw8�JKxH�γ��O322��3�bo;7�5�=L���ǋ[�������p7��S�e��2Kn�"��� ��T���#5o2�v�p���<�2L@����UȂ~������P:�<B���~�i~�=��2	�sQ̢r�1����z������]U%��愺������Sȇnx|03�5�ʄG�� ���X}B��Nt�lЩO�.���C
�en�����0q�ӳ��a�v�jF�Qr�e�.!�6�h��&�c��4�ۅ�eIw�4�u��/I$b�!��^^&a���Y�/��f�9؋LCts7iN�<A��7�U\UUٚy��[FU\����I�D��937�C����x���7G7Z. � �Xw���O��쿅3AUE����;�
 �}uQ��^moS鑒½J���fY�k}�2���L�t)�8�;G�!Z��ޒ�B|,ISlA3l��s�Y��z"[[ϵ���ک�|�sto�{ш{�\�o(�݁^��-d^>0
Fd�h����e� o4V���=y�vn�Dr�4�+VL�į�v �����gƦb�sԸ��4�pUSxV	�|L�&U��P�vK��q;�7��Q�����߮6��G�ف+6`V@$�����8���2.G������o��f�#�o�a��<� ���U�=��B�~̤�I���P$+�� .�0��"��-�i�2r9����ζ�upv�vs�S
�n�֩M���TS����ܫ'P	E�G��up<z�=,.�@L�ײ�Ü�f�Z:�)�u� 1����l�f����]7�R�6�y*��~�+O_�-, W�Y��d	*��� ˵�Z���z���C�B,A`�y���<�J�1��.�J}mG4y��Bǟs�W>��d����V��`5d��;�����q�B%��?5�Ck�l�Ԥ���#B+�Ur{�`�m����UʸQ��b�
��`K�x��`�`�|��\Ѵm^�.���1 �ke�]�_Q��P��_c �m|X��&��W�q�� H�ޢݾ�rR�$F�U(6p�u�*�/���R�Z��2�_�QD�����v-\���ܬ�ڽk�=�a��7��obN�L` �; Y��T�����>ؘBK���P	`6E�>jj��X
9��P�M��Aq0�-᫺��h����f͗��h/������ƄP�Y���^}��z��t��|^ <��ր*)4��<H��w�&�;� ���@;���1�@z���j�Ρ����Q����x[w/�mNc��tzX��*u?wHR���X��?�1������N���?u�o�������g�g������T2��g�#��_-%+��}�>���P�^�X(�^����u���խ���gm�^���4�vB$�`*\r1X��F��c�;�����<-���H�TQq����:���gj;��*�#]�D�ę�U�������������qʸ��XG�;�zL ٢۸�t�S�0�wG%�G������L�K�v�W�`�S��e�}�8�*��~�yT��O���I`�&s���lx7�xĵ�;'�����+�z�ߝ� _~�� el�����n��n�tzb�Â9F���hb�r%�m��M�
�^[8�#�<y�5yLؗ�x��1]8ݒ��3�O���`�p��c�*2]��l���EiZ0��S���nb�E��K�0��{=����C��p��=�CvV���Θ����z�H����ξ�W�����殉wj9�"���%��x7��5�V`���]�����<@#�ue��I|�qZ��-;�5s���\Bg��M���"��)�{�S�7����;^Ʀ�YX4�B�C��F��Z�j�i������Gs��U-|Bboʥ�5���ꈉ�"�%WvsU�66��7��4�7.���O��c	��7�%�>�� �w������Z�a�܌X"���Nfy�'kJ�L^B��dN]�R�#�;�Nx௟�U��3֙�`����B=7����Ɖ������Qo�������˽�7�>��)��0�d	�dR�;z�t�f�O?.�{���͠�<u��fj�!�1���f�$�nH�?����P�kđ`%����?�yI�l��;p<�n#���,aμ�5q�9Ѥ_��4���=���}8ϱ�C�wY��"4g��yΛL�"6�5i>gL������Q�%�L�)ŠOPơg�>�5Z�L[9}ؽ�F�՜�;��`ř��z.�>s�2���8�G����4i��:�y\ZP�mo2�)�\��+��i��?׈~_�Eˉ;�B`�k�o��Al�=/����a��o��5Gau�j`k�i�(X�c�3�ό���uЭ�H��4�P�l�����r��!���Raا
��A|�_�H�>$�pM��Ku̕���^���\�l�m��K�j����B�wn���n�l2*��wg,"k�k΍���*뭨��mݬ��ڿ�����p�����ٽ��B�bUig?
��s�A|�ˋK~�'᥅�L���3�<=�=��4�]׋�U����[:\X�,���G3RɛwU(��W��(Cμ��Ș�)�M��N��nQ���ӍW���X��0�mq�,׵N;��f����Ϙ/z;��0���w'ֹ�W�#6�v�;4u��{a>P�m��A�ۦ:YB�����5\e\�K�����nW]U4������m;�~��i�?s�|��F
y��ӯ &���Ly��O׋hn�Eԗv��ʚS.ͨ��ax������͏�-��~%z�iÃ_A>ޕI��i�a�J�X1{���~�s���E�ͳG���!]~�f�t���魝�>d˷d�\3f��w'�8L�64�胭����u2��ye��G�f�|�_Z�x!t�Va�jg������7P�ۢ3f䇰��С�)Hy��|\_�`���I�ڣ�k�J����>�k�x���z������K.P�5�:ǒ��(�
/����U�o3� �d�ఏȦơ���f�/E�������=�UJ��|ȩG9����;aW�r�]gB�t���Htp�ȏC�����n���8��&���i���f(�}O!��6�M��d�;֨����&ZR�I�5X(�d��T��!ʌn�`N�:���5ݫAT�}�;��G�>�9YϾ�π���j^���DDn�K�r�j8��y0���w>y�Ғ���;:�guf�WDЃ,���v�n�&̟�z���ye1[[���EN����F��=��""o�R���]δM���*�1`(tų��`0���l�n.[a0��=��d�
)��a��SU�T빻Jy��Y��'�U%�^�ڨ �����ߕy��<�l�����d�s~�7������:]���'��i�sb�P:���œ=�]|i��gu��%�]c��K_*���t,���[����8���K�m7��u�9l�"E�*m�Ο=� >�d�j��"�i~��0����N��"BU���w���!�(5�1��܆g�W�Kؓ6�!"�j�w�GN<�nz���-�4���v�C"i�;4��/�\sT�l&�ԩ^�zD�E!0�ǰ���m��c��/����>4���!瞝�������P��#�f����K\Yz��WsG�fd֦�CJi���N)�١,�kr�VI���$j���(�~W?1���I~����K�L�L�PM��3K>?��l[�uޗ���*�����.P��3p<s�ݻOAYa;��۲OW|/�g|t���E��vn�=%C�p���.����&l�F�zݶ�9�[�0]��͚�VmM�	W��^:���!�s�R�Nq��{Xy���]�v�#.�G$���&��iSL�߻Y0M�ک��_D
��W�驯 �ƌd�fܚ��v\�C���4ݑ;й۞�u]&'T�d�\�f������͂ڝ��r�j�ַNC����l^�� ��7�B:as��x��36��<��$�8�Ǒ����M啄J�ˠV�G�]����y.��1�ғ�{a`��+y�\���Z���2訆cn,�m��ݭM{��n�]�k�>��Wڇ��������`�!uCl̍��-a em1[�d�C�nP���t�m
���7C����["aG��_�E��$.8�ob}]��K��e�5,��<���v�>�3+��Lk`$\��`�e�47H����e_�f0��4��혞�G��5;e��z/{,�D6�E���8:��'W�t�.5�L$Nm�âX��J���ӊX(|́ü�a�я�guP��1�������3eؽv[���a�\�lRv8��`;9�-~���vl3����451q6�HH�]��J��:��`?�����Gxݻ=�ol�5KI�D���7e�W
�JȟT���5dYr����&i�<G����n�l^���d����r`�5"�j�Ùɽ���;ld�~o����we˒�4���u,���e�ꯕ��_T&l��}�jO��?;�j���*���5�����c'�ݤks;�GS:M��ӻ�um�v��m���fG��95.�����H�ڜK=�/�Q駖�;7���v��N�<��ew���.${���-��S6�^�)��m;	F-�$�=��C�C�"�����9�6������/<D���\S�u:�!�I��1�%�M��)����lc�6�p��5��#:�_���q�U�(���O�BK��p5��v�̛����2O��Nu�5jS|�ي����ڹZ��p�:�̜sYMqj)��4˴�߃DҜaI��H~�I9N������Ķ�1�;�۬�Җ�+��n�T*φ}����.��d�X�����f`WC�no���nBb]]�f��6�X��Y��Y���ɋ`�v�K���o�G��]���glgl^�{��I���~����b�c�VHv���]d��t��o;����l�Y�E%�tj�>A��qL�.��G��<~�|�~��m�߸"��!�Q���@t����Tb�^�	8���#u%fY���i+��L��XN��m�*-��{c���SV��Y���]u���2vUԉ����J�Q���UlF�m���2l˚�s�����06h�ze�������<������8�L}����{S����|��2X�uWwD��U�b�G	�:f���qg���K#���.�څ��9������s����2Z��˹�BwT�˷�j��ٸ�c
�X��K3���ꆁ�+7�¸��@�v[�WN �i��u��Z��Os*��:.�;�Z�H�}Kz3n����4�>����]� �:){e�)!�lW2o0��fqr��_]��."i2�Z*u}��J�n�����e��\�u<ͫ��mx��f������w�͡+T��U�H0v5S�C����.�.��إV�a��x0۫W�+�{ԁ���I�<U�f�Ǘ�v��Az��'h�tBv��ue�%%N�HIYF���mlg�]�s\�����4+%e����>әçY��o�B����)Hel��4�Nٺ2-9+�����3�j�GdR�0�{n��{A=�ڕ-��QXw�9��2���m�o�V���H���ref����L�"�^;9���]�;,��Ä̢����*Z�m�wu�%Rh�5b�����ќ.��6�
��D�����F��)�t�Y�8�.5P]�Q:����A�;�6�]�^�OZ����ZJr�2qG9G���f��iA����4��>��[]�ԩD۬�A%�L{� �1x�G}�$R7}~_��zҢ\U9��B���l*�v���츱f�pm��X�6tXvމ�n� 9�s����0f�Z���%hi�,���=\�n��ɧ�r9av�)��(�w4-�=B:}��cwHQ��L��Srb�Ҹb�BG9@�5�;I.�'��ĸ`��G:T�:l,��w�(�6C�liU�Հӡ�򖢨�v������f�ehL��TӐ�S�N&0�ᥒ��-�s���;֠�����iic��2�eM���k�v]��s/�ʃC5�N�b�q#d�a$ؗ�fM.�;�ʒ�b#:�c�:�<@�
z+��ٙ��`9��8�c��WoU��k��_iU6s��;����t��V$��b�|�]�9��Ѥ�X1���xow+�ٌ�-�sӌ>K-R�d�ċ�6�I��k��y�s���{��*�F�S��|0�9�ta�32��+���`�K�j	�7��������&K�Vͪ���f�呙P<A�V"ݔQ�q�z�x�3qQ��
f������a���/3��4r���l����x�t�r��)��]�]�v�c�K9m$;O�����>ٽ%��r��Ζk�l��/*tU��L�|X���ſ�qopY��R״g5ƔѽZ�K�
�)M/���f[<�у�����k���X��3N���'AG�+�$ER
g�2���/]*�� \��%�!�ؖ�0IUQ�F�$�1�e�a����)r�O�#*TF�4D�%*�xB�$���P��	-���ߖ���>GGC5RP��;b��wr�P%���ڃ�Е���<����������������3���+�1>ɦ&�!��J�&�7n��̑���M
�����~><��y��?_���~>?G������?��:�l;X���X�t>�A�4�SK4�h�����~?����?����~�_�s����'����,@Rݝv5�qt�}��Y��&*�S���o!���E��U)堩$)�
F��MTyo�tb$�hR��j�/����Jt�#T�Ҕ���
V�����B�]8��i�yE4��RR����&����F�6�͎���)�����2!M%	y�Zu��^��*��>]yy�i����\����=�u�(�ƃN���t������n�l��Z4�^I�����:��O�X��?xQE!F#������W ���T�5mCͪ�ن�]i{D&;I�w.U�1�V��t���g�E�t����N|�w��q��j6�L�)���#����=�����λ:Uo�/<��t��z@�U�y�2�'Z�9���y�����l}��m�`�g���wmLw�3 `0k/�b\w�c�y�22�XD��h�n��h?XU\ǵ�:��0u����oO�9_�V��p���O�$_�|�>g���.<�)�NS��oFx�>�j��f�R2�i�4X�"���7�(dk��S���&��0����z�6zz�O��m�0r��鳽n����Pe]딋 rZ�ų���.�YƵ�"%��c�z}ܦ%�T�R����⯆is��y��=��)tmzD[4�tQ�wG�<ܡ�5��H��a�e�,�[�oڌ���-�]�y��v�X�X�ׂ�>�A�KI~��B��k�|�w���Ye��Fn%`S,�u FV@�v�S��V�y2��{e7Z�z��I��%�+��%��}����N��	l=I�Ҩv���u��bZ�)�E����&���L���"��;�m����-�֝�U��O����'z.�R7*O�=�����;3�<I�N�����b~�����n������G�I����]f���@��4#2�|-.��=�s��@�N'�@'sKvފx��S��.��w�����-���-p[��c2�$��qz�|*d��t2�,:�T�b]�v�6	b�4u*㣵�Jۃ�Pa���0`��ܒz�Z�u����'�&�+�K3(P�s���o��^�9F6t��@��<�5]��l����Z��w1z���A����Cd���)�?`*}��P�1W���٭�]2�T2bɘMκ��6�d�j�,Y��U��S	js��뛔�}�=e�=)��q�~h�>zv/��nN{�(ˊ���s���u
Q���"�ɸ��^K���5����j���$d�X�y�'�֪�j�^�czX`OZ��/������-��̻��p��'}��^4��<��Zb>s��K�������Vf���ώ�̬�z�Èȶ�N�P���~[�mo�(G�������;����W)Gt�&�+��;�4ϾvWʽ� �O&4�.������6�M6'e�C�0<���ʺtA�~�c:dZq sL>�U"I�+о��z{�ꅨ}�����ܪ�&c7[{&;�1n���N��'�����,�����^_\)A���佚�cY�`����S�jc`�!
rN8���5�`���|-�7$���?l��0(aSl��t�=v.�#eI��按�Jz��
T�b�p�����m��W!�b�w�pkv�� ����y�]W����n��
f�l�4�k�-4ܽ�P��Z*>��Ք��wP4��X��P��ݣ��o��8������\ع�w)��D��~�mG|�����q�<���� ��ziuqPV5�'/�t͌XE�����N��G�1�m���n��9��j���t! ��8F)EB���$��դ�}��20͠�9\}<hЖ����,~�g�_����{�&�%#ֿYJ�ɬ��Ԯ�n#Z��
x�j�(�4h��K4�1Խ�]gջl�s�Ɩ�fȍ6�.��y��eu�I��Ve���)����˞C���w���}/{VD�n�b^��lz!�`��-:����&	�6Z3,s�l,����Օ���� ��65Ls�:-�.��X3�5b�/^����ƨ<��L7�S���(���{��Lͱ��eKKS=q�;ג�����C��+~�a1�9��k���W8�?��E'ִ�}��0��ܣB׹�����K���U�cyH�g�����p^��שO7��\Ur|ۦd˝���6��^�7ju9�G��1��E���"v�V�mAaM�~��ٵ"[)�`�T��ض+S��3�Y{�_�OE���[-
����e�hh
f�ԃ�y鯑��6f�D�̫ ~����Gez�,Y���w��s%7XX;ӓ�h��Z�ϝ��cUr'�Z�w���m������I�{��p��/63u�[�76h�fk�L���3�����2D����!��Ŗ�Q���ܬ��>�$<B,��� ��n�/uhJ--�-�jΟ*�e�N�+-����&5���v��1���>��Q����4��v˞],)��֨b�P0 �0����w����ad�^�l���#�_~]?J��q�=7,��~�o3;Zf���a"6�>k^��߻��9lt�]�~_r�IE�"��Zd���vso;J���(�k�rr��o�q���~xIϷ2����Cl�H-� �Ðh�e�su��H�h~�s�
��7�<�2��3�D}?Y�8��=���s���������9�~�o��%6��}P���Htj]>vmL�5�=�����O`MG�/hE�x����#m���1OjXRR�ӛ�����&}z:�������kӽ��{hr�Wh|�y���ʵ-�CJ��n��Ӽ��l ���D�m�"��<�o�J"��pܢ&��a�+�F[�m(����[B��U `��	���<,�.{b���M��Ǹcuj�)�����u�Nm����c������5���o���c�(�qA�U-x��10��7ɹ^��彧���8J���m
��p�]�\$Α}��a������5;\:�W�V��C�K1��+���N�CׇV7����s^]�d� 0�j>� ��-��*���1�.�VK#�(kE���/2_m��/���;��vUۙ�f`���b�`�X��U�v:�����02�A�)(h���������Ͽ��}n��2��_x�c��ǣ� o4���=�O��'o>��3G��3@�J��E���r��9;ݽ*vP��ADRu�H��+7]��W!�@&��g,�<)M�����-�M(�]:�;g7*���d�m�v'`,��E�y-�#�[)#�(B�Sa`_�w����_��9��S�FKm�tq��ZR%<������z�,��2Y,g�hE;�����b�uM�F5����P�����~O��צީ��oe�ք�6=[/��5sX [l�/c�oW�G��:O����5�����l4y�ssW�ƣ�zO1�D���p�j; �$�S\��niK>]ۇ��2*,�Y�$
$��!�"N|�0�Z�^Go�m9k\�;Dg�{�
���T�2�_�Z��lC�ϳ��ˇנ��1�&]p�i�8�ݕ��;�]P�{���3�f���5����H*�Ƽ�vW�ť�jcK>��(W�D}3�fW���E��8\�l�<�5�ǜj�������SU~� ~u�~�l u��֩l�\�wc��i�7]pvp6���.��+.�����#u�ɏ�����׻�����u{����~V@�"cJ$	F\н�1���pa�Q����Qdm�kf��g�k����{a�^��k����� ��$�dB������V��L�<G�qz��q�`3'�#�R��@L�#��,I�-u�S��(ͻ��ww�bgDYkb�u\.짺N_��H2�4.��p!�^�=0)�=c���q�	�������S�
�xm��������� ��ۗh�Ql�a;�wy������`�D�ƿwF1���b�7��d�:�2<�{��y���qw�YP��ݵhx��{j-��0K��N���q���oƈ���G{���F���8�"�ț�ǏR��5U \�[㸦�22D�ь-�ˎ���"y�f/�Lʼ���eyޟfJ~/,���S퐬ݍ�jm�(s��f�la�$����c3�=��ɶ:܂G�������e(�`�S	ީ 7��M��y��R��xB�hk�����Oj�gFκ��y6.4ǫ�q�Pd9�_���8�����e+��߾Io�9�a�֙\}a�~��ҿ2�6���燨ޡ�d�(���gP�Q��C3?ل�h��~I��'sx6a/���R*K"�[ �N�C|@�	���ʄ�*������¯���r��?Me��4�&��P����D��]�+���`ފ�zwv�6���񝖲}0�'λ�u|>-�u��\��@u!�����'��u]%1�w�l��~��˖Dx)m?���90�˦�킔W��ܜ?<��?��D���`C� ��J���R��|������.�^�x_�R�"�rԓCZA1l�ׯɐ{��~����G�(�5Dp*9gG�mØ����"�kd!Sf�V5��,(gj�v>��"��A��<��۝���e�W+�r��t����K�?��,+?K�k�A¨b�w!G��ꞿ|<��ڃ,1�Qe/j#���^�?V{�~3 oߐ�1��P�qQ��Yy;���m� �M�i뵣k��D[�t�����n�Wz J��ٝ��d&�5K�P(Jy��b��Gq|~k=������w]l��J�8GX������3n���R�.D��)�8vx���~���b\sT��nr�X"�J�N��T��6V-#!1��+±�ڵ�N+��y��F�a�<M~tm�A����)��톟�E�e�oV�ds/(3MY��簶%�_��C����t��`�.��@VzpQf��*��5�����ಣ�3��	�{8ı�CSaW6�/�f�[u@���R�1�Kp�>��,���/�B &�z��)���5r���酕R��<SU����՗o��Ef�D������B̙����F/;�+�|���eH��N`���[A޵{��4ηo��xz����^���>/�Ľ��v�݆���Z>� �]x�W^�V29M�a�H��7�,�	 ٔ���t�w&)(:�h�+;zǒA����n��|�w���U!�4a��,�R�@�@����ILo��K\9o
iM��a/��Kl�M��!����J\Pc��yO�c�
��w�]��7?TR��9N린j4�+i��&!>�+�[��<2���or0!�[`�i�m|ن�'�nfn5Qt�S.ǁ��=0�����l��k�B^9��"yۮ�Y��,u᙮�{x��U����a4�n>�5䠱݃�P/�����׺�(4y��t�_\HJ�='Y7�k�f��>�42eSʭ��&�Χ�������f|. ��q����I>�������������X9mO��n���b�ߕ�=װ<�ԼC�R�卨ekɾ���w�P̀��wkxp�H�$�c�#e��ͫ�S��275.��"ʷ��̶�T+�N�������*���X[����瘉�9��������5���n��S�m�����_�W����+<B ʋI(���B�)�m��{�k��[ns��w�Ís�7x�%:iڳ����f�	X��˧���)�P�Z���?��
{*��Rġ$�i����[�s]�C��&�/��3�4�q�S�4}+F�<���~ٯW5�i@<����k���]b|�E�݊��o���UҚgu�Nw�·\΄N��N��xA�K�Ɏ�Pv�%�w+��;K����ŏ��7����_�	���C'�J@0�h@�B�F��(���Y��x~��A8�y�͎���3g�+�x�e3j�}����F�_�M�*K�aU��*^�D���/�+�\� �"��`f��@��[�� ũ��@jfM��U7X+hU�X�"Z�_ߨ`�W+�z�A��wֹj֑!�\T��M�[��9��g�]�%2�Z�l����E�JS��ٕ�Ȭ�k�{Z<����r�0d��硯�kO�/TqA�M-{���E���݁檭b�<��X׋�Dz��j�cW��˘���3�*<��d��{$k�!��o���4��r���V2uq��m?v��xTn���|�A��F _SF0�P��K���y7y�2+u�Pt���wezdHީ�u�!�G��n}��jQ�(ׇ|a�>u�:�����wՌiG#ݑ\��xK�#Y"K�quѼ��˔ɭ#%��3�A��61�ڍ�u����Fm�K2k���Z�H�E��V��~��)�$�~k�b�W0�����4�o��4�S����4qq�3�I��C3���Dc42����j\jQS�!������AΡ��x@�̖�b�m��L��u�N��b���4wh���"��sv��z�L��v��ux��si�����v]oNMD�
�CfT�Ec��p�Ȓ�+\����H`_e���p�;�ї�n>F��s�gp#AH?=�>��	 �ʁ�T�
*; �7��F�QI�6����E������Y�#|�ĉ�
��`X�?�v\y�C[�{v6C��ʞO���5��֫;��Do���/+� ��;��`�~u�=YӖ2�pA�4dѫu��y �sT��ݾ���]��L�#}�e~ _��eb��߶�i�g�0�歆f�qv8Z�V�^Lj��&9�=�`?���h˹%ŉL �k�L�U�i&m�W�<ڢ���O;�Gr.����OY"c=��EV�� (w�R �����Z����٢yP���8���ݦ'^y����~;N��w���d�"�"���~��zgh��[��!�<�n%�S`j�R�=pٜ5��f�q���ݶ����l�=�{B�W���>�	���Xi��Źz'��g�n�5Ӡ�ͧ;�/BSe���Yr±��c{\cO�츔��ȇ�UW��.ӛK�-�;�J�ff�
�֨Sz�,̡\�r^���SK��S�W�%�k6�We���k�&a�;V�w�Qx�3Pb������Yc�O�Y����b/���z}��ޝ��-��;EPT�Pʷ�z��T�W�]�����H�6��6�0A\N�S�o=J�xM9������8p�Οs�[���B�شͫҷ��T����x+�F��l��]��m.�������.����lŁ��*2.��8I�����#,�xi����ժp�Z��2�j9�V.�쩧Lz>�q{Vo;e!\�v����B�X;:4Iws��)=%�6z�v:�b�5L�A�ysI���B3C��a�/:Y��ע��n��=���ջ���Ǯ�b��!��Cƥ*,��c9JWX�jl�����H�j�a�z��ѷ�$�8�2�JT�]̗Oi:�C�]�7��K��b�C �uݤ�c�Kk�j2Tt�#��S�*�#�����u:�q$�֜���T���T�`y]�5����Of�i�g�G�����{Sݝ{�3q����bM�"ܠ�8�4��)�5��h�k�gu�\��E��F��0�w�]OH�hy���1�k���(��{E�[F��n�\y��SxD%n�����O!���rv�;��k�u99MqkGoZ����1��9�vΉ���}���Gu]BI�ֹh]!x�t�"pHr�����K��X&Y�A�F컺�a�J��s:�T�9"G���L}�/�t�+��l�/�������荺}�:����n6�ݚĹ-�:�õ;�5b�b�Z��VJ!+�1�J����5���V,��`V�y ﵁>c[\�T��)wb��0m��J�=�`3K�F��L^ĭ\f�&����nQ�����6��:_!y��0�\�i�I5�u�]Fkv�����-+�kCB9u|�����wq�y�*ߎ����A��.R�˓X��;���;qI5�e���SK��U1YFGz�����1�	�̓��bz�n*އ�-�k�4�c�����+2oX)����7X4c}Q��u���K�:�h��_u��	��L��d��w`�v�^d�I
�χ	S7
��4pvk�&^Z�:�Q[�[�29��Jo�g� ����R/��Cq�d���:��3�ʤږ�=�[����K�6sN�.�0�l��&�{���gKJ�pg[�&r�=�G�(�}��Q��;y����]m�7/8=GH�0�aFF��=�����}�R��Ѧ���>�v9�x�6ŵ��M(�9V�j�������grN�hJ�Wz��}:nm՜�8��T������R�][�p��1M4fC�wU���4m�����A����5����t��/>�ƈ�U��w	�_]����7�7��[M�݆�9iܘ���\��k�K�����躍[�DT꺥�3���Ӵ�J2��8^#k�!��s����B�&q7�����T���h?��C��	�Z3$E^Q�5���*�������y����|�������>�_�s�����)��{~��U�A��tQ��EU'��VvêZ���<������?����>�_�s������W�AI���A���6����#GM4�6�=�^y��F7���������~?����?����s��O��O��Qv1q����*N�Q%�Z(Ӫ�����5c�����D����7q��v��.���_9zN�J���1/[d)�LS�&��j��������T��預�I����m�&���sBUv;�z?�wY��l�[n��D��QGF��裶*�.ت.��K�tS�Phӭ~������CK�V���PtI
D��h����:�O��u��N,N�cCDA5���'TUWF-�i<��:6ã1�
�`�X�=L���b?m�^�sڡ|���t\΋���֝Á˭}}��W}��u{P�wے]9\�&�݄[�����>�"�!��������U�T+��������>~��ƿ�������l���g"�)0��-���M��`��m�%+\/n�����V���8�nS���V�;�~�[j`so={S��O"n��z�X6��RFKq�v�8�逳D=�Q�v�[�[��gO$��A�Y:�K���P�^��}B�j�.*q��;S5ͱ�r�.��QN���e��-~j�2i����<�~`��K��jz��S��3{ ���ur���6n���" <0�M�䑡���1�8y�Mi�1l��0m���f�p04Ba{l��A�a����͝��-)�M/:q�>G��[ﾜ^*��}t>�=��;򁣯#qd}=�O1��c���Ɍz���W�#!g��L:��`��/��,��,ơ�覻3=�as�ʻ�~"v������߹�s皯ƫߕj:��dFfc���?�����+�����L颉h�`0d9M��׆�>�3�t�<��~a��o1b}X�I`(��?5o���}x��h���y}K<��s��i���7�L���Ɗ����*�G�;�g6+�����ؤ�xw��=B���ð�,��#��t\|_6�G�by�����[�:_f�:T5�Г*U����΍鏇���wv幢�Y\��+'	�zm�p"Y+5����v�4V��k�V�u���5N>�xm��x|<��T0®DpȨhQ�U(@()� �$�Ncm��;��o�Rm>�6v�KU���}M����Ĭً�K4�j1����ǡ�(���h�Y���AO���2�U�OG"Ym�Z�<�J��X�h`C�/�؀��g���Hf8V�scRa"�a�#�X����5�����}�2�n��^��^�l*��b
/��'��{��֮�̝��a�!j�^z�An�5�4[!�7���{�K�UJn�J��Mm�>�:���QY}ö&�ƛRS����-�K��i�R�&8Bm���=}����s��ϵz��j���w���ܚ�W������
qP�̥���1����#�M�Z_ �,���u���>����0�r��̼��5�p�K�"�G2���A%�X��.�ށ��\��`�黒����c[b0��<�	.Ғ�-5�Sv80���m�S��R7D���6^���T�dCT�LQZ��W�%����Ƙ� SP��
�v�nU�^v�'=Z� �CC0mn�[�cҝ[ۘ�c�Y�����ȼ1lO���k�������w�`o�:��(���L�@�oc8�L����Z�t�1l�oء2����u{Ճ(�\�gUL��-�8�rw_��g�v��0ݦ:��!r���F*$5C�n���p�g]��ȂQ()&���n�R� (��κ���ӌqY�"���ʶ/�t���0"�n�gW4:���N�4�4�+�)ji&��)JVjR��Rխ��(;���i@0��!��TԘ�F>����3���!�^<�͍���&�L	�c�P4k�km��u��5�5���Ô��;�^�)	��j}� ����d��V{�N,������a��V�C�띩�.�w��5Ӻd����M�)�HM�H� ���D'�o>6��cz]�D�M>��n[�i�^$�1\;��x#�ڽl��F�i�k.�l�2�9��i>F����;��Sȝy{�M'�x�=����nL�|J�MG�E��3U��(�����L�����j��aKL�̤�O��i��6W<T��Y�]}���i�.�j��\_���E�⑓q-Ƀ�[2���lRs�!�v�����Wv���{��~@�q+7�Y�B��	�E�ߛ�vĭ{�L��dR}��\��m�Q��c�Pƕ�s۟[�㻯k�������gL{�-��xD�Q��K'c���\LY��]U������F8p¸�{��o!�Xͱ���Ʋ3��t3��>�ld�~�;�t�J7����+1W�C1;͎4�O�37^Q�T�n
������y��%�Wt����_�g����.�%>��:�.�*}ª'O.\�a�F�H]��wMCGq.Ukpb��~�K��a���N׺�L�࿏�m��;�Y��ROҏ��&�&:��}[��)��t��1w",���k�]��mUCk����i)�y1���{�<ARPa��
V�ZQZU%eP�P�߿�����?<��ϟ�/���%��.��JD��I�%��<�O��[i.�8�w>}a��0��t��3�-�O�~��}��Qz#�c^/����2�Ns�U�d�XH�d�9�E��lפ��/F���n蜔]ö@\4����]�O��Ȫ�<�6I��ZӬ�!��=7�P����[�K�%CO��q4���{���}�Z��g0�c�<�'#,e�y�M�K%�;�qc��Ua��%�<�!�tĉ�w����k���\g�$��K&c�f���b/:�B�r��e��&f�����|�Ѭ�l}u�\^�L�I+�٭;v������6;�9��̘�G�ۧʵ�jt�Pk	\����t�߷^���X$�i@����5F�y��5���u��fhQ�����;���"-�|U�i ��u���6 �+q����l����W��;E:����2�B�]�v���k�������dK\��p�z�>�4)ͼ[=^�V��b��H�OY���~�~�
J߾�2�R���%
ޯ#�(v;�q�wE�e�YQܚ:��k��s�e��5��z)��hZ.���k��������2�s��9��\������}��p���Q�,��	:�vF72u�T��0�;��Y��W��c
��tvNv�fT���yM=�0�`?M������=���������BP������)
�B����7�=�I/Ɠ�B֟��0��4�g�q5�\��vl��W13����S�C\Z�����v�3����y��_�� 1m��1��,�ax�˷�����v`k�@�C���|nw���<%N�*��)�֟l;��E>����K}b�~˸3�\x��^6���6-%�[f%�����d���f4V)2�����2���S�Vj�驼��A�~�NM�h%��~��o�Qa�=�\t��K�xny�p�d<�L��N�S7/0�1F�?sP��y�L���7���U�R�e���X��q?�Ќ~;�CKͣ"l�	�\�=W�
z���xcik�f�V���H��}j�����F�P��p��?`��Ǭ#B��;�j�,��[��"�B8�OD��������	�.u����D@����vd�^��jr#V4�y��؉̈́�sI�%�xOyX�&;�?��hkH&-��`�f�z=#Z����cI��n���
��n6�j������
ނ�}m���W������	_%�\��]8�^߽�K����-8
x�t������Sx��tiCK�[W��Ю�ox׬z��UL� ���6F2��H�jP�*�m����]�3��{$�w���!����W�YTxܓ�U�&Z�G���~��%+�;eI�6�=[C� ���H0�h�pʀ�E)����}�����������|�#�������%�pj����ʤ�	(i��D>�����ܪ���<3��D{!��$�kf�*/��N "�-�x~��P�~��B�@5g���/?�I7m��?	�Yf�,�T3�&���[�k�:$Jw�;�!��p#����+P�z��1=ze�ͭi�� ���BD��j�w>F��H쩆�� 6XgU��f����W��5G0�ر&�b�ᦚ�Ǖf�M2g��;b��:�!�WE��O�흡�h�:�yG�9⮲������A�x ����{�M6�.mץ�	�og�s%��V�ڟ���g�s(YeIQӾ6{^K�p[ml�ls�a=s)��*��x�	���d��axړͫs�N��Χ�ƥwP��]ŉ-�8,�����t�Ny�?D����{���k)x��>�Ow�����gPͻ�ѩ��F6ڹ�"u4�C��0�i|�,�V�S���R;S=[u����K� TsiP���*�� �
��G�4ç��m|>�b�n����Y0�gy}���Z���qи�n������n�'j�sc��\��_0�|,���U�/�V\�j7���Xt:	õD���d�έܽ�ګs�åj�Dr����w�sM��z��*¥�@��Ɨ��SQ!��\�0C��v'U��X�r�_�Ȥ(�!	wv���yq�!CH��2(C�2"`eR�����C��d���lp�ݵs{�g*^��� �P�]�åC���ǂ�d�O�;�l,��3�	E���Y�]����6�A����B�Y^����j�(������qq���ͽ!�<۞g:wB��fhJXMD렄TaxhN6K�kLgM50�ϝ���r��Rzu��k�˖h��n=#������qL��T<38V�(8�E�>�z���צ��t����d��p��]Sm�jk75C= T�7���hG$���'�Y�ю��|�b����-�A��0������6<�����l���'D��t9)Jfӱz�/�톞�'��W<�%�̊���Y1M-���.�3��;.t�^@��~��� �&e�����/ގjw���o 5�P�nwOq,��-��{f�h�4��sE�;w��
�0�of�U���Mӧ��N�(=J|s�ш^�$US�ٿ�^$�G|�&�W�)�@��p����^�9��%L��LK]{VS��b� �;wc�1�|���м���+�=�N-����Whh����3�X�{71ǆM�d�`|U��ȡ��UѦ�F�n�+oP��V̕���4�I>&��Vv0j��)�W��t޴��W���ӧ n]U-$��é��U�����4��l��
��#���M��N�\asMA�	M����᷽������q�~�_#�U��`R�AP��
 >|���u(YSP�ͭ�^�ᵃwG�;�X����s�PR���=�L�������wԜm�%�a��!�O���ݚ���[0�/!��Dy��5�JD������ZY\doR��}���!w8c'0���B򼲱��0m�Gg��N{a�}.a���2�Ic�8�6a)T̀�!�^��pQ�1�QݾP杳t6���a#�+�}m�y��&��L��~xyO��Kx&���ze��tgv��ɝ�8��9U9�pQ��Q�'���K���Fu�7;�~�����@�O�2T��r~D~<�Љ�ʄ\{��'(.~��-��L�ϣ���g�g�K�7M�ךv�w�߳�?i�iQJR@���s��C�X��N0��B^S��O��M�Q�.�F3���iRQ�+����^qץ#%���@����[1�u����M�_�+8%�i��>�R6i�q�ET��f.]i^�cU���fu���r�6�35�+~Q�~��]�
�&��N���#�3�ֽR�T0�a�"F�z�o�����w�s%O}@m
I�o��t�5=<�\�l����D,�����v��:u����x]��:����í.4:1��m�v�~�y�GL�{y�>qe���z��⁚���������gl�wF�p���b��3^#��_�Q�i^�p�����/�������/{�~����ģ�@aUt
4#Bw�������������o�C���\3[�����n�.K�UAb�8М�;�Z�:Jڌgm Ԩ���>?�������v~�c�b�9ky��,���"���� �]_�}U�vv۝]ʧ~o�������@��F��{��N7�v��,a�R�Z%�|n2jUu%��0�iENLDoE��0���*ETE��溯Aw��<���݆Ɗ�3��Lm���ff���P�kܲ�e�Uj�k��xy�m}��e��������E�[<��A����ڤ�r��jj̎eε�?sa]c�F]zo�_����˰�ڿBq�c�2������Âř	����yٯ�
D�g)6�^I`�n��Fr��z��zaP�W�*Y�����Q�A�,��&=��4z�h�(:�fy=���E΂%�z��n�!�X쾰�-��:{1�֥7�J<.�J�|{U��P�}��}�~��<\T�q~1R��񦭢x�t{���ɺ�~�_�ߦ����B��R[��Wǚ	����QXnDَ.?�&��<�1E<5~R�������B��vi������1o+f��!��U�� v��4�P��9V�FQ�����l�z1?��V8�2V%>����Y9��p^;I��I#�-j|;|���5^�D��f��r����`]Ta>��d�}1��u� �_ ��Ȍ3��a�H"����INK��L>+��c��1E�� ���@،����F��ߗ�?o�d���]��9��Jī��͍N��B�~|G��.i�D�DƆ@\X<��o���" �;ޯ�,���J��ֱ�DD����|���-�P�Ӊ*d�<u�4MO����vWʽ� �D���ر��b��5��jf�A�>�B��B曚D(Ɨ����p��[,�-���f��<lc�8O��sӷ��k���@C��:R$B���v/�$Xu�s��⍪b��we+�!z��1��+,�~=z�s4��i��i����~a�х��AOC��]��W��6J|b�K���M͎��yk�>>ļ�pL�:z�֨g!��F�~���o�o����{�C��>���ܞ쮥��F1�=n���_�2Gd۸tj]�ûY׉l�Z� rw�Ǧq�w�ٻ��$���pDa�gM	���9B��c_����k�R>V&͕�ٹ�?i���Ֆm�m�mcq-R2lگ�o�M�j���s��v:��*͋��v�]{Ϥ�W[��z[�8��y!��C��;��m8u�+�W�M��սc��  �}+8Ú���2�[o�L4�8"�*��bPVk���t.�E�J�h4�_g7��{vnYv���m�V5���Ь����`��X��\�d�Z��㗶�!2�E۰��V�W��k�3:ج<�ʲxM�o��n7zhElNj�K��5�uIH[[uUѼ����4��Ì:���2�`j��f�u��]��ں���7a�f��ĺ-��i
໔�y;4^�`���U3V�1W�^*�wtiX�pYil���:�c�ͻd��tU��M��	�<�p��l;�Efhvv؆�WI�L�o+N���*s�̛k�)�:�5�i}�}3I*�}��u��op;����|��}]hZ3l�W��l�	��d�)����|8km��GY�%�q������n
ҹ�Rm}�/�s��Văoi����e��C:����x��;�"���/�\��oro0����}�`h�f]��i�j�_ۆ��+����&.�k$D#�Ռ�`��؋ѩ��]���*�껫�F�b%d3���`��ok��l]��r���jm��wڎ�`:�&Dz�����9kj<�v3Q�al��O&;G�ꝴ�b(�y�ϔ�{�Wn���Jtif��&��f�m���9y��0.�Yo��EU赻���<}�ݍ��C!rj���۫�pP  �X�0��7���]��c�g2����������s�[��\He��"��*D9/�cZ`#" ��rU�8�H0�}x����A\hj{��+pe�]C{bj�.�d��`�t*�)x��Bt���N�jq+�hl�m@X���mk��6�oU��c�=b�U��@���o�u����k6XS:p8��J��Zj>�:��7�A;9����\��J��{���s��>�/�j���Wje��}��l95d��,fo y�j]g�{�@B��_4�܌�ۻ��s_g�m�(i�&y'�/�;J�7�����|^����;�յ�8�[�xr�I��}�p	#��uH	{�|:����w++u�.¥��Ѯ"�sI`�X�[闓q�
�#aFe�GΎ��P��Y�Fv8���;�Au#N<X�l�@���4uD�m��9��b���h��3ORu՛Kx5�@�����.�vD\�YHx����.�J�[�Юt��=O3�j��N	>꣝�N)޻�3�=/x1z�SDFn>ʬ��E]�Z
8�=o�6�����I�?(�af�
���.%�t_R$���|��s�/�%�IJ��\1o%�Z5���mKPvM3i���틮�A�Ǎ�������3�,�L�0�
�<j���E�
��F�SY��3�\u}m�,f,�A�%�ܔR��h��P�H���]�;�9D��վ*(�+�7��B�8_E�i2��ꠊ�l�5]��	4U
�d�	��Q�	#A���5H�Q��"D#J&H��4�RJ��j"A���#��`�q;�!	6SM�
�[l��y���i4��w]UT[i�(kw5I�UUGZ��*������|��������}��~����b��F�㎷��cgU��)h48�!%Rk[X5�mU�l`�7���>?�����_��������3����PWX��
�m�������!t`����ZN��������>?�������������~��~�q��E�Qm�%bF�^񪍍F�+�Q&�:������4�h"��y�i�G�΍G`ߝ珗8�4v��Iݫ��:
i5�Wl(ƓZ�I��B�(#X�m�Fv�lE��AGE�A�"(�&d�b���j��1ֺ��`�l��5���kcv�z��Xآ��j��5�o�1�TFb�[Z���i��k��=�N�4Q]sc��:�m�Z(:�6�c��M;f�qDEQ���ˢ�j��8���='0|C�8��ۧv����Kcm|�qUZ(�X��QI4N'U�ݱcl���ݢ�ΜE��ŉ:�g6,[4�i�����!�I�OeR�x.�fX���n�_t�8�O�����̋�%$�8U��U�7o�$h�e �i=��Z��k�F>n�"�F
�="P�cy�:����J���!�Xa2�(!�w����ߛ��w������j����!ޚ�������y��]����2�,�UL��yk�����R�"*��j�٪s�f�KQy*�sMÇ�#* &Z��6U��B�zw��O1�cs��e��W���F�Z��U�������O4�1X4S��ǂ�w��ׯ�C�mAn��]�p�Y�Q���"�E �ύ|��i)X��\3?�����6o���Ji���;�n�~op�}�'kA)M��^���8T�p)�ka���R�c���/Xt��׀�mpl���!��D��Χ'��Q���L�M�i���C��	?7,�
�02�t�m�A��ګ��f�3�3G@^R�ܼ�-���X�7���Bl�ru�׎W��I�k����3k�b�|�QT�c̓�knz��D(�<�\��qͅ������[�r{�L����wzq���d�;{�m�0>5��8�{� >��\o���'����0+�az���lQ��?Cr1r���(Kx;��37�����iz�.�</{�/�A|�|S"�m�����?�;3@#�"�dQwՓ�5�v�wv�����ʹ�?��rJHv��kUMJ���αq��U�r��w|��ɉ�8���8zR�Ԭ_�j��

o�uF��n�y���q��Ը��V�׽�gn�M����β%�u�뺩o�a"���^��/P�ǵǼ�< ��< #�xx0� <=�ozo%a��<13m|��f�q}Cu�n��5_�������_<7����Ea����Q>u5�|W�'ɲ�۽Y��zW�qyaM�[Hy�:z�f�ً�[8���
�Sat��c`���zf��1��,^(!Ɠ79�%�}�i�G6?[X2[&�n<�̧��t�&Ky�u�{f�~�W3"z��N;�����������x�K&�V��.�mU��e<�Q(�q���ZL�r�|�(�S�Zd�П���k�W���y�H����rO��e�k�IE'��)��T�_��@W�*��u�qzkk��[pm)����E�؝�6�/7
�����1S;.���~*x�^,��Ѝ�C���Hg�0���FE�7R��q�X0��25�\�!cd5y�ŧ|���"����*�5z�H�7"۵���`��ްL��d�M������xb�]��|�`ީ\�ǒ��}kK���ީůF3%�Ⱦ\�TC��iP�R3�p2\����j����z�L��2K����0���xZ��ή�a�֨[<�^Me��]YY�[����(�vd7|#SHw�Y85|�`묢2�7�v�#2&X.I�oVr�ɐtYƙq��i��;S�g�:����0��ȫ7x>��A5��i�pI�N�8��mwv�Zs^¿��?�O�d�A����Wn�������������a��|����^����O�]����1x���え�����,���4����}t	�@�c[o��8�,&���_~_~V,z�u��P�!���C��7:��9�A�'h�j����Dl�xf�k��U�@�a"p��K?Aٛ��~T�"t�!3���}���L��r��~��dŰ�E���3a>x���lx����}��n�Ȑ1��#�t��	�d\˵�PQ��ٍ�:^�\Pb�>6��_��l����u2��
����2��O�bۋ���<��d��Ӯw�$G3h�C��Y�?��M��5M �w�iek�o:MP�X�����S�����ϓr�n�٦O��`9
2��^
�Vcs�q��5/j�-dŻ�1S�޾�����y���M�|�EvH=r�,#��e-̔�b�t�<��r�7c�q��˿;�Mf���B�/�r8�C�#�٫�a���8بԫ/#5V�F���,�q�2�K[kZ���)�a�T]��?e�+u��5�����	���3�?:m�S����fJ�@�f^h����˛��":r�ǟcj��p;�]LV�����kY���
<���[5�A>Q�>g\�`�{7��{ݑu���!�p���mҭ�����V��:���Ob`�ʂ���gMȕ[�����/�?��8eQ2(�ˡ�v�_s���8�~f�;8ɫ�9�5�)>iS�M�X3^���$r��r��iɞt(��b��耙��T�P�W�c�����/���2k���2���T�\ь͋7�/V�ZXwj�؁^�d��{hN�s���t�eHyޒ�q;�%�o=CE�+�K-�a�"�n�u���mkܤ�IJ���=oP�t�b`&�z�-{��oL;��#&���]��T�YFKPI/���9�Z�ha,ȼ=EA���Oʪ���Jjf; ���+ЂF��6pFf��C@Jy��Ma(,$g�sM{�;=���Hi��s;l1���f��箹���@TƧ�yn�%�#8�~�}:c��?���3�L��T���Ȇ�Ŷk�76�t���'��Ё����n ��B/����	3�	���Mx�yIg�R�Y�fk먪;�ywM\ӄ�hٯ>��~y�"60�K�|j�P�������Ŝ����7:�T����/f�6r�K��U�^}�g�ֆ}�¿D{c���L�S��"��AO8�#�q���z�Pv7�m~N=tQ�6�kN@ՅTv���8��,��'$_}��^;��;d��n�������_Y��\"���_aJN	U!0��}�5����N���q�*�<6���;��/���g;v�h='Ck�.�;�Fb�
�_r��cS��i���b�ۺ����o7Q��v��
�F�D!��~W^�}��~��~�y�G�p����ρBE�M�i ��t����ׁ�9�������6����L��3�����jҮ�CV�2���CD��Sn��`E�ˆ�y�C:jh�1�oS@�oT�3��s-�ˁK�/W~sc���� �	�I[b��ݹ"F+���sӽ�yTK]���cu�oEA�,�ȶv�@�]7>��E<�)b�1�ǹV�y��B����d�v��վO�k���:I�D�i�+gA��N:5�O�[�2X�{	�`%���
;sautT�j@��aCz-����cC�q��]D�^��4zցޡC9MK�^��]�9SR�8muu��~{`zc�&=3�&�ZVⱶrjmS�O�T	��@�m�Nd�	�|úk�gV���y)6���b)>�O͜T�z�4�+i��=1���-��@�CC�x�3D�O���h�d�c���������oO���T���� 敯�2��~w�*1��s����ˤХ�p,.N_��c�>Ƈ�1;"��~���Of��5{�p�D��v3�`E�R1+)�>3!ً�kvFץY���b�g��^�]JS/�� �&b��{�c��>w�w��̊���7W�ľy<z��{�6�����m̮}�R�f�{Y}�Gf��P�u�s�mq Ν����o���[�??_w���_�%�F���go =�sx.��ߙ�L��m�jD�� %����MR����MW�P�}lF��>�d�;��74Ɇ%���* cC�Hp]'����I���7'��Zy�(�݁�y�fsW6�!��v\d���
\o�)` #����5��u�}#��a����u�ScE4�WPZ��M�t��3S5��\zF�'Ѡ<4Xga��?� _�y����U�?"�%���������(�y~�j�T��Ag< P��l��b�%C��xl`!�Z=�׵ϲ�;n6n�b���J1�N<sDע�v���8p����A���Y��׼G^�ٹv�iy�u��,�!��@���?b@�B��ק��ʅ�d-b����M@�5׮-��&}Y���L�䘖��[��к�lhU5)�/��D�cۼr�O|Pmb�����������^?�I}���D���zj��P;N�r�{�[U�F���x���&s܁ߜj���O�U(	�Z��i�5K�L���W=���S�Tst��S�ڏ	k)Ncݏ8��y˫���.�lS�R���4��ٳ��3s��Q�|�S�$������zGׯJ�'����&��=2�)�@��:.��ԭv�{]l�����)�������|L�8l�ҡ&��j���)rsEp������4wQl��=|v+���9�a�����8�D��I����#�����2��I�??}�?�J}!���(���
�1^����R��%	��"�\�n�7�v=2��[r��K_�]�ߨ׾�yw�xK��q��P�����b ���U׀���nE�Z�0�Cά�*	�޽�gf�B��?yOŚ��@��YƆu�`��oL.rY�����l�R6���On��X��B�mqb��s+�Y��W�	�B��c_�ߞy�v\�M|]&4���#{���� �R����ǈ�
�9|� ���1|`��z%���"�r���y(t��*(��DnV��]���T���l��wӢ���Dű��gX,�����<��bf�� �M�UTE#N��f�()�Y/�-�����b^���.���ݛ 3�wh�f�vQY�o�[��C�(~�Z^�3���
��6�/��I!^_X�s�Zߪ�o�;�ϤNy�w2%?�ˠ��T�!��n�9��ni�ne��`�U�e��L�d��C*d����̫
ճ����OZ���4�<?b�}"G2��0s���8�w�*�Qv����:�\ow5o�i�6��T�+UmMX��:,��B�E̥�ڪ`����c�����>`�C�3�o
x�'�z:2ڜB��ru��Zz&�]/``C|A�y�APɨ�Z��Û9_I����Qwa�r����~��������2��� ��������7E�R����Ӛ���?OG�LOKxEs�Ϥ$�?*��5v��R.��Y������i�Gn.i�%�7!�D��wtb��=��/������Uתּ�]Ks�>�����k8˯�nptb�h P:���/)���_GP�PY���a-�[}լ)��<>{��Y�7'�eaCŖ�������-iP�V�'^��Z���	�tzO�;S�u�Sy�ز���nl�Ba��u1;�!�m!��7+�&n��vEŗ,��S�Z�:g�k0h�ni?b�șĮ��7��0�K��5/ױ"7��W:w𦗸3��T9eՓCM��/�������)�?NHe#7����X[���zQù�@y{�a����喽z_�.z�t���3+aE0��u��2���AΧ���|�b�� ��$'P
T��P$9�����w�b���=�������WYs�ר"�\I6�XY&I����\E���@rԘL�0�<=Bb l�8��ɸE�n���b����1���	��X�c\wN��{ Y�2XH�εa�g��*��h�VZͷ��󺍱���!�����,��0뵓Vp�k�&g��f�u���T�/��&��^���V�ޚ�b���Wo7'g�W�^1y�f�U�	�)LA�u�P������B�D�����)"f��
9݃2iv,��,�-9��r��j.�����ph�)� �`��vX7{�wy�Z4Wϝ������������y� �-��R3^KK�ph����E�|���L�cx�z^[f2Kzp�B�����_���L[9x�g��F�:��ψ��`�x^aL��2�a>�����2i�1�����l�7t���yg��[��>��BT%ۯ`?��>�yI���iϓ��+"XSֺ��lY��f�`�E=3��m*r��.�b����EDkW��d��E ^�����8�*4���)���Ne�ѹ�.*��y�Y9O�������%��6	*��@~���tkT[��a���1��'��=���{��5���D�󆪀헾�g�AA��"�j�w #~���V�>��[z����O,~���,g������d!�3����D���{:D��	<�m�r�cޭii`��"�����5.�Q{�<���.�zkP~-9N�%��s�b���ha��Ȗ[iV��!	�o�/���B��g}�g�����޻BՔ���vc��Ϙ��l��\��7�7̚E��u�x,'�e2֞���A�/K�����t�����ȁx�)݆��&����E���YcW����j{XP�&C��k�*4�T�ꄐt��Y�w�ڎ-[�f�&�-�ÎJ����}�a�i���uX�á���TD#Nl�h^�	P�0mu@��6຺�î�`�7�j]v�/B�b��H��/���׾{�����矻���G�a����{����'g]���D����M�bw�i�\Sf���~ŵK=�IS��:m���2�~fF^��C�gpt��J�͕�+��O�b)>�O͝�c�Z�Ǟ<ӡ�~�6t�*��35l+��SQÖ\+e��<5�G7����?�c�Ur{�u s-�27^��nj��$ގ��#[heqh�@����DsoLCnZ�->kk�-�1䣛��B��u�ٚ�[�gUB���f�>C@H�A�^9�CCf��ΐ)�ء6W�d�B���p������k���5[��o�܄�D;Zށ�$�������zO":2Ǯ�^pVr�ܛղg�3Mv5l3<[�/���No\3�O��
\k�8�8�����7�q	��\Pc=��W��r��[J),b�cP}�.O@�36^�JxXX_�!ڕy�F�v��=��F�������X�	q��c3gۙ^��[c��H������7�\�t^]��Q�|��p���e<&��xd'\)蘶G2}<��vm�2t5C0�%[Hw�h�ef����\��l�"��]��I�)�:72l�J�6�vp�Zh���m`B���N��Ö��+�0��lù�8�� ���f�6y�]`:��n�f^�+x��.m�y�n8�.-,�׵t/��ҁ>8��K��l�a����5���ܹ�5�9Z������A̶_�Nt�=S���n����E�YZ.�k��h���$r\z���#�����j���ٜ��֮��u�JS1��f�.tL�2	����X�gW����X����ԕ{ݜ�������m�u�e{.�'ܤ"LnX�,��z��m�M�(i�*�=ʰ����Q��n��-�t��F��Sz(� ��tI��0l��������z�j���B����D�ӕx'S��2p����J�0\��r:IlQ�'�Ԇ����
.�w:;,JC�ǅ��o2� *�U�nݡ�	�vD����s:�r��2���ق-�\�ԉ(�p0ss;�������L�[�h�F��n�u��3����6m���ٲ�����5����w�R�9�tkX�h�H��v˺���Hn�JN�T��
�־:�QדB:��ok��u*��sxh�Mճ};eh�Ir1Of�gw�pՐF]%R���PJ�T��"�N*�p��IZ�=EG�[ۍw�>籋���j������1�D�O����-�C�=Ձ�!1&UufM}����%�TQ���M�,��5�H��R���UA�NỄ�[Vs�X("C��YY�TZ ���$�Y�w-�'W�6��ȷ���O ��пU]��r0:�&;�������(&f`�7T� �#k�kx��_b�C�8��ɋ't]�j�z�ye�+i@�86.mf(:��-�{ˈ6P�yU�wHv����Z��_{�(��}��o���L�gw��B�T�{���pގ�&��:g׎�}4k�+��_wJD��]w/6��k�̼��f!��I#��w8L
`_]��kV�c��7�����(���ٵx�Ρ[�VJ]je�r �Jj�-'���0�l<��.�NWզɋ���7b�g_`��{b2u���yͬq�{��.m��q�2��L�5:	����qr�t��b�q�e:A�Xw��mK�UN����s�9�W�x.�a������0��!]��H1�	�U,�F�ϯ1�l�t[�S����b;.��75��TSh�]�:wp��̗��;�b�����얕5��5W$��Y��IpGn��[$[�xXq�-+ǲ�qmV��h%�\�W���DP4ibV�s`ʹ�v�#�KOQ�8Pg8���M��Xj�qc��2JXeKȦB���ǘ�磮�M.;\�<�����Ȍ�_��ؘl[�]��h��E,��2 ���y:d\�qf�����G �<A/"N�S�v���<";k��Ѱ�?��y��몙�XƋ�}|||~?ϯ�������_��s>���V�;Y�TkmX؏��׍S���cCM�y�TDtj��FN+>�|~?_��������>�Y���j�/�����ZJ];`��Q�mu�)*�l�n�C]����4�A�c�����矏�����~?���~���3�����l���ۺ)�CMPi<���~N욯5���UP�I��kM��ࡈ+Xѵ:5E������l�tt[h���c�t'yjk�Em���a�gmgZl7Z��٦.����&��F�5Z:8�&��4֣gDlnَ�m�Ӫ/�5v�tW�������T�ӣl������65TA�i�U�65�t�M���I��X�$�A��5���.��c�͉����E�j����SS��5�uGFѦu�b"�hյW\|<�ua[����#HŚ�DhZv�Y�3��S�w���^[/ط3�;��{�������������ʽ�����z��j����'z �3Q�(۷���)z�\S@��P��'��f/�rSѷ�l��}�E�Y[�.�1�$sӸ��<z.ϪEע�S]	���,�	���<��@b��f�[���\�yr�dݞ;2�Ie
��9�{/-l-ј���y���U	��c'A����S�����y�cn�0�U�ץ~���Um������v�H����>R���F��g��ٕH}��7t���]�C2Cd;����w�����s��P������yecmF�!�Χ���WZV�u�]��9��@�yu[�o���߲}���A��� r0ZS��sO���4�g>��קm_r��a�vzFu��XD�%�|�͸�ɤQ2�VcɆ��<��^<��������!�fJê�[Q9t23���G�1�����{��&����z�
���M��c�Os��R��LU-�=��)��3��Setc��|�cO��/%�{����^;�īWGSɼɄ%�Xe{�i�{���=g���>Ʃz�[=�"cD.��L�0ϲ\�y��vs5clm��f��ǆ�i�\�{+r*nۗYWA�޻���`	�D�g�^��b�#�=kI��u�}�U���M���H���$�:��j��skV���r�*�����S��w����ߟ?��Ba�����������(�A�[��O\�dNlqq�D����7���L�|C�!O���<XH����}��z�'y���w���G���"`:�4.=�F*���9B=�މ�a�͗hC�����-�C�G����k;;������LL[,"�~�ϕz����K��?O��q�����{)U��R��8*[�iR��������yw��v͊h��q����x!�*�9ky	���#Elx4.��v��-f��zfG�����w󁩪+����̤!�v��C���0^$��f��3"�����~�foQ���ߥ����! �<�+��?~�
��7U��l�5��{e.L���1t�i�8Ym�^G0�㐛R�y���Y���\V������GA%T"9���W���u�Y�"�(^SP܄ǜ��}��0��������=�Q9EM��2rk�⇃G0��|i��q%0��"�q�y�c:�>z}�T�Q��[��C�w�b<�s=_��k�~A�F���t�T:eՒh��(:��=G���w�/�.�������K��M�٬&���9,u��*�UJ�,���UI�	b��������0�cQz�*�/*���n��$\�J�����o��8�sr��>Жvl�N7ã�.�!��h��:wK��������-��n�=Nc���ձF�lշ�U0U+B5mZQ������o{ޙO؅/�����!ce>}��R×g�c�:��!5@՗㟏��ܱ�`�f�����D��;k�x�<�`�]RX��b�6��;�~�T�8�Q��X�!Я�o����_v����!��ME'�,�2/]'	�\�#��,g�O�E��s��q���1��۹���1�f^����J�pb#�v�B�^���+����\g(,Ь�3k3^�2�0;"��U����!��y`��I�f;�����;\ޑ�}��`'*1��� ��Uy:*M4_RV�W4a�rp�z�@1��XU�E�"�깦L���>�ו0;zgMR�R��\[�����u�MFS�{B]�8f���6;/����TF{��(H�vv���;o�:%���u�%��c��Yu�q���|mu�2�}M�?���?L�}�5�9UIt%P��N&��Mjm�4���ݺk�z�?_F��c�n�ba�r�ρ��,�L��R�;�|y3<��->UQ����\�SQy�c*'��EȦ�,m�B__��s�Sn�ѩv/j"��o��������Hi�Rn2?�b'�j�E�:��YƠF���kd�8�����q�v��N�gS������ b}C���m�q��nK_^u�uۓJ�B�T�����G��a�z����]Rn��].�s��b����@0<�����L�-t�ҹQ�s�=6��g���i��dVO��|W�ݳ�����@c�ǀ�*؉r�{&�5�������6�1~zj�6�R�'?<:І�@�"��ʡM5�j����,��8��ʉ�F�*��M�^'2כ0w_\K׹�Tm+4U���WC�����m���rE1�ַmiu�KUO_^9�&e�1���qd�xHJ/�z�\Pw4��.`&S���3�k�Ga8��*�%��?D�L,R��'׍ș����a󙙝�F4mk��Ί΅���𧅜�=T�Td@m)=����<^�?��O� ��m�K\��P�.�����ix�V�
~�՟��*t	����i>vί���R�a���4"�⫓�u�m̍נ�c_��*�"��Ei����_����ռ:pi��7�L=uR�V*f���-4�y����n�TUøq�����GKq�x��B�p͋C�����G�_��4475��MX�6<�z�Ŷ�Z�,�w$$t�i���{���ӭ�|n	� ����w�X~����W��a�?ދ{�z���
��=�3c5�F9@u[re�d>����c��.�Ͻ x��Y�&�k����fT�����w��P\��݉έ����9���3�!{]�	�%*ٚ�x]a+�u��F:�[���ju���x���25�`o�>`�������{ޣ����(2������9�=�+�:���!KM{�8����،	�LZnka�����-�z=����S�F�llj�K׉���?*e24kh����Y4V���'���k驃/�;(�ɶ�	tf;6�;XW�����H�@��㞢���j��g�U�K�"�T� �3� αဂ��"bە��sF�K��0��׸� ��T�`��%Y����Uq�v��g�b����G�@+�'�V@B�6����>:*)��3��n,"_5*zǳMb�&�2~�b�N���dDO}��W+J�T��ߧ�+p��ώ���=pZ��c�_�[�կGHwe#��S$1k�m�������i��sĬ�?\%�
���j��{l��i���!��6h�4����Ƚ��I��H��Jpc݂�!ċ��C��.�1����Ԅ�+`9�lo���X�S��T���161P��+sw���}���^����˩�>��F'�.1}��f���^ħY��#�>b*�3u�xd�1�v?bۏ��ߦN�;�KmG8w��D�F�£ʎ�{��s��9�<�{��r�v�B����0��>SH�*}�3�}X�� ����[u��1�|��rZ�]A�Pt��ʤv����P�ٝ|�k�:�Xbg���񇾗�.�T��׆7�y���o���`�Xe� ���Du��O2*C������7�Qr%���?2i�.����P���H��v�\�ʹ^��Y��rָ��fBI"�/�2�rȿ��	ћ��?>ˀ�3j~�;��#:;;����-�ۨ,Xv9�n�/ZO���>7��Q�&o=	y�xE���'͵�hʼO���d��W�)��6̶�7�����|c��Gk��[�F�d�pAj�J���aye.1(ƞ|��B��N/�haB��[��s���B�L#�7Wm�vD!Ş%ݲ!����3���U�}��#c9�3_R���Ý��M����q�4�c�	ٳd<׏��^���3[tݪ���0u���3�dx�7�7��2�8F�����^�s�Ak��W���'�X&��ߠ���������C�]<�Lk�J{]O��ѝz�iGU��	(,����1U!���u��Th��yfq��!K���qlnw�S����\��RJ]��5�=ac0~.^��#L۸�_T�9���	4��A�d�i�����*�9SE~uN ��Ǎf�C��Y}N{w���)uɨ����̾d�ͽ�sb�Tt�4@���	q'�>�]�+���̓��I�Y$=M�!/�	�K�����U�6���6�Z9�8�w2����3W
����)����h�w��v�S���2y�=��o{ٗoQ��v���0x�Rn����Y~���A�9�W��Ki�����������*�$�#<+ڇ��_�{.)[ֿ��׶y��𚚀��U�x;�oض�ԥY..n�"pDM�����3:���jלoH����	�2�T�sH"{�J}ħȐs4�kW�<���E��}l�w���-��+.��>{8�5C�[Y ��f4b��|Xٙ�=5�w73z��r��:�QL��<���0~����[s܂��J���O�O%_���0��3{0�$��aq?�<c�-5%���M����y�B�hi�T����<~�[�-����W���v�r�]x^�,�Žs���Ĥh�[�a���˼q�ض�Ź/؛��I�mPԦ#LD-s^���2'�)%� sf�Q��/�),'�֜�a3=�����Y�4D�Hu�%�g��_��S���c'���IP��3�q@�
�Y���oJ�9�А�@���i ���O|����~B��e�w�٦M>��i�K�P�3���C��yj=����Wk�g!�%�����I��M@��U/�:����,�zl[���bR�:���t`��|���O~�9o��%�A�ϔ��M��qOסRጎok��w��X��ggb���d��{��[y��{y����a�oa��G[p�,uޖ\��9���Bd~����ö�H	���=��X{db{]M�����R�9������6�C"�q��8��ߘ�g����T�W���佖�p��P�o����R�i��S�&wO�v�ՙ��s��D���4�L�:�辨}yw�ؽD9ݔqi1�V�y�覚|9��Hv�����Fbޡ�@��6�Q�v�mȘ��}�+�umCؽNܐx4�^g�v�FGk�`�`��3ګ�/lJh&l&�M��Cu[���;���0������3� +���vL�4ߌ3s�hP���}�Z��v^n3����@��ηQ��[0ff��K���>�2��܉���w�5v�J���{Ne��sw.KRvkUc.��ǘ"�y���E�QM�VV0��^DxU�ffڕ1n��*�u|�˝�˫�˥9��q�����7%� U�WKط��%R�����ηG�a�wƯ�,���pfR��Oڐ=�,j�s@��g��s����ff7}E���~l*��U�f�v&�o\�C��1
2־=�gc��9YR�sz#��p�=��|{z��uVIԄn���{��n5�2����p�I���3�A�X���Kٻ.n�뮓�g.)��`��^l=��s��3�\��E�w�9��؉��y������`y�y����qiP��� �����r����}O8��5*�����8�W��U�-��s#���Ork��,�p[�������!�k�BS� m�;�*C���
�$*_�q�9�@YlF��rf�fî�y0��Р_w�A����?jy�b���ף�kLgM6-U��+1����Ft34bQ���瑙�������ȃ�Rio@�Γ���\�hOd��i�yϵTC�����/��`_>�w��� u�2uy��B��2���c�|D�Ցwh�y�Xio[�>����OX��s�l:Ŝ'W|�m�o��a7ޗ������EK����M	7-5;o���<&b��;@�2���#�͔he�@�5Cl7@-��H��n�h¤�}�w72.����_����Y����O��X{�(բ�ܲ=ͷq;��k|���7;��mm���uz~ ���Y�Lۥʀ�N�<���:�lQ��~T%?T�d	lB3�y��r,���Q"�����ͯC�K]j�v�<E�ӽ�v�d�<&���1�"��?A�V/0ao+�_Q����߷������*a��j�bb�c�yZ��m�::t4ޙ������1蓟J�9�*��U�Wp{6�o;�H#όݤV�����;�K�X��*U��Z}j.�ɱ�`2*õ��=s�i4F�[�N�:NnM4�x|<��0�a������[QU3���(�z���P"Y6ݢ��m�Ȝ�ٷxlᑉw��cr:�ۉ��[u�uQ6�R�PE���xX�;�2�zm9́-r��/�靶�����[�Hgtv몺�p�������o2�Y�r���"��;�Q�'�c��y�U_�����6EZ��a��}�m9-���L����L�s�Uä��>g��4�)��x�'m����i�3mieN�k�F8�'�)����͠�_f���2����W�t��>�|X���.CsM�2i��v�|�\"2�Wt�כ3Vِ�lT-�d:	��t\sz5��G,W�ƻ�>0Ɛ�$t3�|]7y�g)����ȏ��K�Hxy8�V]���C*&+���ϠZM��;�����2H��w�Z�x�k����R�7��Q��u�r�|�U{L���<�9��8g�NC��F�l}���������]�D������c�y�2$n�N2�*�����꧎Ї�&^�جx:qg�5�_������"{�ȀF/��D��o��FԌ��E�7���&�zg��L����
������/b`mE��OE�O+Gn5,����:m�n"�:ʺ ��Duu��3w�cv���ܮ	�
m�����a��]0���:��3��tT�6jCj��p�7"�q�5�z̽� �$I�f5���;d���&�콲���f�˺�$�%�T3�Y�A�`w �(���1��:��&���׫��Q�L=eu"*pR�ZWו��չb#�.�ޣG��-eE���89,��۠w�ռp�H�MH�j��{�,�o���Dڕ�
r�j�Vq��3Ϝ�m�1p��h��b�s�o��Ν[c�O��[���즖���a�]*VX�iCz��mrkSaK�KZ��>�Β��IU�jz/gt����:�gsdr���̎���k5��btsn����a%"���.�0Rc/sf[���{���ɉȕt��� f�V"�`Y�g��k�/I���k�A{{�V�u#64�j/&��\G�olnTFBk��� R�a�ouWI�3!I�^8�l]��=��A��/s��e#�M���S�kvf�[�-�TA���5�P�i�Q�^+�X܄K�r@�2N0Ҝ0�C�t���]!��>0�xa�w�0���z��W�ީ��/�1�0�傥��(S��]]v,�Ո4؃W,��g����	΄XV�h��`N�A}*N�J�S�4��J�>�!�VkE�ݝG�c�!�4���Xt`��5Tɤ��F�Q5�[.�uQ��c�*���D�Q3����83v�>�j��DI"4v]��
�c;{�_I���P�MiP��.Lxv�m�-LA=5j���2uZ�NP�8F�Y��*6�]`'"AL��hܒ�f�w^W�k�,�i'�r��f�D,����f�ջ7�Vkc�n���b�`)hN3���7Us��39�����Y��+��gu�(�uo�h/�:������Z9>�ݲ�w��^�ڸ��GT�MJ!\��pSR�sݻR�󶤙9�]}�~^�4*�H�MG���o�N�ub�|��Wg@�on��O@Gq��镥iF����S8��ORUB����wP5��fg����K��뻭�������]S_a���P[:(�����N"�q�ԝA1��������{ы���IE5f�:�Y�-c�8 �T��c r�6�5y�|%[l�ٚ�QN.b�ڮ��o�ņ��K�Q��Ǝ�ܺ�3sv+s�b��,&H7��k�9\8�k�����FZh��-������8S�w�����Ǡ�jvE�W)�d����v����3o�2�v 4�m�ـ�%pZ�3&Q#x�:��GD�p�8�Sȳ�RS%e�sm��������yI��٦<.�y��T�p��T+r�գ-���s�b�䫣|b�W�D��d�P�C"���^�I."�X$�dH�I&�D��\`|lZ����Q�&@\ ��6d��$�!r�1�'c.��$.Pi�3�v��m�;�:�ݞ)����٦�?��.��h�b��N�5n��"(����֎��]�m�f1S�?��>?_�����_���?_��������bѶ1Ik$[Y�_��5��5��]�cl��Tklji�-��/�:�c������������~?����f~�>�k�S�4�؈�:3��kTQ5��#��.�EX�ؠ�س�UP|~��>?��������~���3�z׶֍�lj���Z	��A����Dαmm5%7��ն��v�NvM0%]�mT�7m6���""��Ӯƨ��j"
�.���&��Z�QThu��vQWb�"M�l�מc�/1����mv��9�M�ݺ�+V#��UWEj���A������3���jb�2GO]m��]�]�i��mM�&&*�����Ɲ���3��-�U�Ltlb6�F��e�u��TU~���ɦ(�c=�E;���QŊ5�6�QAZ�=�横:����ը�v1Tu�t�[�@Z�<�	 �A�B�E�A
n�PG-�\�:^,�!7#�q�8�<M�8'z�����(��U�`�	b�'sM�m�W�9����a�c���$ ��B���5:�7�u����2/��~y�����_�K��.XIߊ��a���*�7αٱ��ϏoD�t��[��+��o{��=��Q̼�-�=s˾�x��p���sX���`��ܟ����-�J[Q�*��=�o=��2*0����n{H�f���I3o���<ڟѢ^5�=�;�%��� �[]�.�|Z�ÊcN54[��j�,a�th�"Z�ڧ�B3n�<���R��w�o���s�8\��~yU�b�����(��d�ޱȿ:�3��J�t�wfj���]����a�~�k!�����e���'+�gy�`9�������'E���82il�M��tv)?^-�����nPQ�ܵ��L��YP�o=�]�Ez�%	�]�3���V75���Ρ2Fֆv9=�t��퉃��yR`�6����������ڤ)����d�dhl��g���̏��3U#�xy�ZC3y���0����ж��d+9clSy\����{h��e�@K�e�zN�is#���t"c R��Y�Xt9n/��J�ld��`5(X�ʗ�/b�݇>�I��Je��U��Ֆ�f8�@Ԓ�;G�ɗ1(r���\[[�從�tT�ӫ���z6kޜ�ɘ:��r:k���5ͽd8�.��3ݬ�%�!u��qe�+Uý]�\/�Z�,��7 ��8��Y���Pٝ�3o<ߞ�oo0�{�L-�[�S�v�Ɂl���]�dM�<��S�9#%����POm����t�7N���T�w�7Q��(da6P�kw�Iû�=g�=����S��� BzJ;�e�%��6[�qqً7����d��y�C
P��m/B�ϥ唈����`���c��}e���s�O_T]���������=a�l�����>އ��qh�^]r6��~�������F��<�7��O��Aw\�� ���}y��kϞk���0���d�٥T8�ww�\����\wU��C^���d>���ݖ�h!=A���H�����V��va��Ə�Ԕ�z7x�1�>�40�ƒm��4�`�1[�gT�6���z�}�mȗ�iF��Xj�gӲ,;nD3v���F�1S5c�ʘ#4�5y]�b� ��do���Y\y��5"��%6B{�+v������`�>@����͕6i��V����M�!�ƙ���G�ȋ�N�q3�v�s��U�-��o8�v������x�W��)�X��t� �X�����E:����xp�ΟwVt���]�:�e�38�fN�QڻQp9��WTYH�:��b�.�z�M��U^ ��'h�*���H^��<G��;��$�s*�g��eiϷ�̭��dP[��7U�0X;�r�A]=����ӣ�[u��#��_�)J�kp0k^r�+F�Ǒ����6�һ��jtgK���}r=�	�n�-�����U�����Zè�x*{ۙ)qV��bZ���r�>��}��#�t����c�U�S��)a>���g��-��,+f��[o��q"�ٔu֦�_v}lS���"��+�2�"���8��W��MX�������H�a+��6)O�^�m�����h��hޥ�(~(�%M�לC��\lDj*v�ngY*+�b.��^��e�DN_^9�֞��Z�w�������:X����똼��W�k4�}���a匿 �:�b���>#,fn��J�-;<���m{r���nl�S���"z����yb[����O�ὼK��;��U/1��5���3Q˝n.��u��5|.^NqG��T9M�4�1��z)��7�z�-ǽ�x����om�Ɵf/K[��]+n>�Ϲe���.��fe���g�+��b��н���ܽ��\?���x�驾���ǖ��vk�1�c?����rk�-�m���k��Β�S"L��Sɏ3A� �=�,-=*+���r����m�Joe��qF+4t�d�o3��F�W(�v�L�u�(��ϳ��Љɩ��.`u���:te���f�G{1>�l�g���/N�j���oR��ڕ(��#6	�7�W���e �N}�ѫ��G�^�z����ّi�Xͻ�d�q-Q�1���[��̯=ܖ�ɀ�[�e̕o��Rِz�F��|ו���+Ur�c�ý�΢d1���K���\�>oge�fq���Gt�P���,���F��e��\��
��4bZ4��>��u�k���s���!"�^���j~�|q	k�� �U�����n)�;�3[��0��v{��%��LbF�^'$'l��и��ǱS���0�nzᦑ��A�U����xV�=�wd|R��nY�v�����EҒ#��f�"Ш��y�9V�OE�t�^P�JJ���Ogy�u��<xv)�8��(ͯ�i�*���d��z�̼;'8�'{��]�3PvXA�=�:�x�����J������� �N,�n"�n�3Dx5|�&}ZT��T�w�E�@fߛ'��So4Xs�?r��jen��"/����/kީuevk�qǶ��r�ټ61U�8hN�t0��1��;3P��f�6�v�w@Ӝ6A����k1V3���f�����k��m1M�C����Ż���(�	�Q�r��f���~����D�@=��ja��C���`-�2� c^Ĳ�����Puڟ"gx�1�:h@�]-��s���뵗�
���&zW[['��:��4��2��<q����Q#�P���F��/k-[��7ck�l^d��0��DM+�]�֋E��d�)�Ռо��3d��ߘ�a�;���Z��>D"������rD"&v9+��5�S`�ZMA�8��j'el*v�i�Xy��i�{e�<�Pʐ�jIYl:��N�K���ۛ/��e��eQ
�O�b�k�cS:�{wi]��G*^>��:�\��g�4P� <��qmBzGUsU��vB��pٿ���J]�s��X}|j7a.�R#�Ԣ�������Su{��L"\�¶w���x
7��l(X��Ʌ��n�sB�휓1~��,	���ܧ}ҭ(U��+��q�3iL���V3�ז&u�����U�6�Sڸ��*��SQu`G��y��K����J�R�N�t�Owu���L�]�_�i��`���[3>��똠����t��4�v!M&��o)2fV�5���͓�Ax����@�mT.x�N���v��f:�j�=l�\q�T���3�KR]�Ƞ�F+�f�|�7qņ2�����ry��o��b��z{m����7%��+�]2���{f��S*��dF�bl"J_!g������<�.��L�M�"���l�ɇ��752���v�"-�y���r�40���š�-�H�섫�U{=w�wk:�o�N��5�@z�.��<��r�d8�d���^<�Q�:���xF�ie��^�^A�a����5�on	l�!�����e�p-�
х�����%�)��c�Z��(����;�]���$u�0f_Z1t��F�MU-�$6�����e`�OǿV��C�q^�~���!7����pY�!��W0���ȝҰ����6��LF�h����c��::븱��+uǶ���<�'|��&s�����,Z�v�38�7��(E�qi�Ͳ��]C�*���nY��T�K]��	�k��ӷ����Д�m"���]8�}k'z9�d�f�eM�rZ��m3���<-��~���N&�'�}���x�<d��R�^�hq�9,�햢�v���"j|����گ-��쉬x{�V�w�t�4��y�������Ve��|��%���L��^!mJ�k��nb��di�9���@ҕ�-M�2\;5�J���x�*�=�1��0��k|W띂�����}H���m���YF�����]��f��S3�w��3]Nnͧ#Kz1��;"�E�4j]�w��U�+�i��M<��ތC�'�t�M�e��@�G�0���ȼ�+�F�#����jg&��w���yN�c��	2��ޑ���c`R�O���<GP|�¢�*M%餩�}z�6���Y��I�7�W}��%�X�ه	W�4�m'iٙ�W̧/��3��TCj���7��F��Ϋ:;�A]�.u/�kY:jvj�KX��.i���^�6�S�.Wa�\�P�M���{���M���*n�Ƙ#"7�xD��ouX���zSn����>��DF�����pI��ހ�M=�^��Y>��@I��NǸ�ho5��ͫ�v;�X.�}ɕ�{p�Z��^y<>J����[���t\�C�{�=��?e����A�6�^���{>�qO�ё������>���t�1]��p�^tc��_�ү%�}��f����捁^0�����o\X�y�\�jK�柅Ϯ�M^a-���S
;��B�q�U�;s�T�j(�g2��������m>�$�ES1�d�b���i�D�T�70y��d\d�!����Pf��C	y�V�Q�~��a�ة��v�fi��ׄsv��[T7�zyE���U��@݃R��d�YL�56����J%]վ�Uō�>g�������Wڕ��eVRY�ү���X�m���&�#\d�V�[s_e(�Y�l�Y[�o��|����.��-.|�/��g2�U�J嬫{���J��y��9G�s(��Cz��0�iC�c��Ȑ9�[}��'2���ۗ�qa	�����q0� 9y�&Z���<��S��߿���YM:H�_�wK|��粡+�~YY�jؑЖW�]�W�*���n����G���ݙo�\��[|&xg��ס�9�
�޽����Tn��vrtR����GU�uZx����%� ��S�x��m��3y���Y�3��lk�LX�ܔ���;lm2���q-ʙȊZ��
d��m�ƫ���UM��#�����Z�h����1��k0kF����S��k�B�u�e�j��\�ˮ�j�vR2,Or�+���;�k��d@��^�ߤF��J��]g��<�0��35Z�5CL9�6��e!�h�q�Å]\����yYc�p�J������sz��I̎@_nzV��Pn�Xd�I�/�%�)�
6��N�f��}��<�,��7Y�>�r��z ͺ�mZ�B���<��y=��2�B�S?t�ܤ7K�}y-eᬭ�}��Z	f.�/��n���寫��ٹ��K�mE�a��]�]*��cj�\�#:L��Mfv����]�t����n6/��a�=�{s��SP��X��r��Cnuk�NC�Ge��}%�)x�⩲��\F�,�z�N��/a[��[u�Lm���\��ǊUb��<�/+����@M�ՌЍ1cm����D�?l��U��ei�=Mj�:f4�U|�6�e;[U5Y��x�;ݡ��agw[�6�
�g��[��TW8�S!��=Uo@��u=�3Mσ��8��e�J���cV�͑��w*��M�D=�6rdu9۬�3��aƜ�f�Ikz)D���|Z�Ե�i|�Ket�Λ�f�8�6<��re���o3;����L&o@�ݐ�W[�+U�{��F�S`���}��~��Jn�\�K ��T�4KVrS�G���nO��~��*�f�C���b�s?~􄥨	�P�hB��ۓ�^�F�#@��^K�+����ϑnt��3A�)Wu��Ag�r;Aܮ��Z3~����W���d�c�:�l�Ȣ��IT��x�n�]��-F%� �і�|Y[-zn�>{׼��ԭ���Z�[]Őo^7yW��Dɨ���Vwt�qއǞ��������8�:e;6����8)��=�h\���s�u���vwga�ڷt�g�rU�9j������,\p�Ǆ u��S:Z�x/c��	=YFƅ�[����=�Ÿ�M�;^�$�M���(Q6w\�~�!ӕ�k{ TV�Yn�)Z�:]��l*1���m�Y����황����ެ�8a|1e��*oa�L4'ʛ��^��6K�Kj�YwaЮ�eI�-SډAv!�e�Z�,�v�!W9����G�U��Y��{fl����Җ]1n�@��Jm�Ce���NN��1q	dw6|�,M�B��p�4�C���Ԕ�;C:��Q�voMY�����9L��ܤ��;���� �i�f(GZ�����c�tP��6�*UmsX��-+�{F��;�J���1][g��o*]�F��^ٝ3�_i�Y#��a�z���1SC��y��)��\(����*$���@�^��ݘ���ܩj�q{�n��㻭��.\�l��:���1]�;�NH�_�ŏ6Q��i�z�{�g�x!�bG n�+����ՠ�r�&֓I4�e����{�[�`�cC�����ޘ���Μ�⅍�ta�U]9/��A�F�EZ��,��$)�ٰz�՚mX"����WH�p�w���S����L̎i�k����1
� �FSJ;n��i�l]|y�@n�Q�:<7HC��nt-��z���V{���Jҟ��=��ٟl�)���ZQBꮍ���h�,�&
F�L �v��ɧuC�R��0��uư�����;_s.���(B!��cM�B3s����cy�Mrl�|�8���t]�W�bs�
.��Z��Z�6��ym��u�/�gR��tۥW/���v��.I3j.���� {kz��}WÇ7i�d���&'K���F=�;�֏Vq9���������ї��5�&�S���*��U��괻�%ʉ*�X�wD��\U���+�Kܰ����2�)��(�1tB
��u}Zm��1��8EO)��L�o{��p��{��.�7�8$Ⱥ�dS����k�y ���z6��K���@n�V =��rw�h�-1��'C�S��ʼ6Ȝ�.��v�� ���N`��N�k��S���%Wɕs�pL<��[��3����GXFs�S-
#� �i�P�h��Mwc�yM���Ά�4pT���]��m���]������粁ޝ��u���r;��4��]�}���V9�#t��R���{\�z1��bKړ+,RȜ��:=�P�G)W\h�H.�x��m �nZ��̈́m����LPC��*���I��EE���*-���^F���4ǛQ��kw��|~?_�����f��O}�7�0i1}�=�j�y��G��8�mv��Ӣ=�~?���������?_����>֩֌T�4UFƓۮ�F֎�v�v1m�wj'�7�<�~?_���~�Y�}om�4h�f*�mPQ��z[�(&j��b�h��Zcwc����"�ы�i�6Έ�8��&�5��"����D��v
���v�jIj�a�F"�U��n��&<�q�˹�{�L�y�WE�������[V
����PQMy�8篜u��:�$�����b(�"��%j"����i�D�M�v �h��Y: �>kd������ƪ&h�5UEQUu��-vs����b��U��tQy���"�aחt�u�j�+mJE"%x��1�������Pe�}Kzp�Q�}���G�x�@�7���)��$Q�z��z�Ný�3a�a��z����^��]W�8��0�{�V�I��q>q=�b=�tzR.��Q1��#"+�{��[Lwd{�|��'����Ņ���y\�^Lf
"�����M�u7An�U�jI�2���-�\k���̦��4�FO���v�i�ȁeX����oN�=�`5��4q��m��j'�;�+�����ݵ��(�b"��3߾���R^��s�a�g��2|4�9Ri���D�L�[�q\Ծ��C5r�+Ma�8�w1�ga�c�������2�ɋ��Y�x>mS�:Z�j���πŀ��c�������r(+k�������l^�r���K�`2�u��OK��r�{�\e��)0�x/3t�Wq#afhJ�Z6���~�n�����
a�x���#S�eޛ��v���j�7-ʞ��P�E���v�:W�A��C�̇"��l)��:g�
|^hv��Vp<�	-[B�lmУw	O;C�T��
�s�۠Eu6�O�sE�0b�`C�7SKw���V�s��fә���\ ��7����f�\:Ε�gbʧ�x��&��6h�MJ�{�]����v��猪/swQC��]-5����u���yQU>Zp%Z����P����^[�s,�9:�䫡u�g���p;9��h�u1ޑ�*�j��]I+Q��їY������g9d���Ji�q�d-�ѱNcһ�_"���qں�I��F5�b�uy(Kh9]��s��8|���>��ɍ�`ӝ�}����o6ܞΑ֌*<!�]ʙ*h�f��K��fW]�»:��Ƨ9�)���fFq�yރ^)�I�-5�^7fS�.��!>���XX�	�aU��j��lYm�����^����l!���N�����Vr�!�_�Y����b�����Vb�@��`�:M���2j2�c��k�.�j�Hd��lva�k����U�0.��xp��b��6�{`ά�:�F�2^�H�^2��BL���=~���"�7��Xq�_�������u�AI76��,��S��b��2�Nne���g�9ۿTk�B����Q��<wI�9J�p����>0�ܭ\Ѥv�4'Kco��ƪb������dt����<��N^v�-\[-�Y�K�v�rfoT;�vC�f	(�A>nF�R7�xܯ+�{���
}G	�Ido��ݛ�k�\�h&�OP2Q��_+�.�h�ºO����"�N��Ƿ��7����T�䍳�|e�'����bt0���2k�>L͞`���ӛ��J��x��9+i,�IG��Zz8�F_U5st�j����u%�3�����[���|�-�uwB�[��4,��e�����3=�y�m�7}��[n��i��WW�4k ��7BYq8M�U�%�_s�L��w��yB��M�;��kaV�G�磃�QI��c.8e�zu&�q�3>��{�/+v�V@UՕ�O=���	m�y���l��C�X�k��-�����Z��c�}�Η"�h�w�;l6N_����'0.�����o	a��',�{��Θ"0��d�����T����o��Y>�fgV�u��M��Z����	@DI1�Xfٖ���κ�kG�qD���ȫ+�m�Lүل���BU�ΐ�����O���:�6� �zm+����9���(pz��YH��D !俻���*��JJ����' �l	Vgݶ�����]_N�1�E�w�=��83��q⯸end0����+�����S9/Z�cD2�J���l�~�՝�o��0��U�Z�l���=-��Ͻ��>��;t(�T8����ڷ{_�ڧg�����ϖ���u�j�h�!���3q� bY��/�A���z��A��w6�͒AO������=ʌ�+u]���Yy��z�j/��|ϊ㫋�S뼦�����@~�vb�K���p�h<�t���Μ����Ƌ��5��w�6�`��5J����M�U����˃R!�E�g�x�6��b�\foh���v�fwk��fuP�L��m�zr6k!�NUtKr�����%ڢ}�
�O�����77����L�&hͦ�]~�Ees�u-.��:��'.�v��0s2�vR�Rs�xWu+��-c���,}�=y 9˔C�ݲe�׋�h�g]�ױ�e����7X�q�}�"l@VH
��ܪ���3"�#��;��O{l�fcvX����Η�D��wj����9Y��#zTf���k~`Ş�T?j�>w�)L*��i伊")E4��s�2���\u�L_S����8���-v���q���Dn&����۬�Y�o�_r%\�܅�{�3{{
��{�*�e�Ѳ��i��J�Vshj���WU��]=ܵP��y�殱y����(WY�Q/��Jw��e�f-��mH@�vq{<&�r�O������%ߡ�d.ޟ\*J��u_���:yfh�슓�cy��Ŀ�$�|k�9�pCvt�}fIx��Y���1��0�:�r�ݝm���[����4͑$��AO�l�����i�����6�뜦�m���nLn���K�.�Nz.������{�[cIxhvq��Ŏ��]��ϼ�����}�9}`�hk��zcs%�q��%�A�=!�t��y��:��S�e�E�k2�&�������0tz��Y��5�wn	�fC�h�"�\�7xd�̚l���cͺ�X�	�R�����t�gfn~�)��^����Țw���ֲ�:ʶh��*@��v|v�;(��`���p�0�7H>�� W�se�����8IX�M�V�cM:�P���ܹ����V	*B���zC�^b;j��ne��������o�P�30i4p�>�;�=�7�Hؒ�x��W�SY�ַ�A]s7��UM��>�i4�Wﾪ��νsU$G;�ͻ,W�[͆|���R�{躢U���e��f�2�C7ã���<��Ko�ÿ��מ��5���=�R4�sg:���fւ
��5�B�nQ8��ߛ&�Gc(��N�1�IS��U�����(��=r3���w�������Ujo�RĮ�0l��f��e�掫���ձ����z#�a�ᔶ1���R�y*�7rʷU��s�Ϊ�-����[���d֨����ԺG9�M�U�Ѫy#��绵�q���KA��ł��c��[���3�鳗/7X���s��x�-���.*;A�p��exԾ�vsu�i�hc�WcWq^y$�zo	�GI�5���]{3����k�uMt�H�sv�\�׾��x1TF�b�
�ߝTm[���'c�Uw�7HA�3wM=��p5WX��x���>w��t��_"і0q�"#��rw#*r&��~
r��N9/>5�0n|^鋕���8@�:A@#�����U��z����,2�P��o�_��^֩A3�q����	*n6.E}w$�Dr�w��,�,��/3դ�Q+R(TE�Di�
�x T�0kṝ�UVWIQC��5�Cnl�Y������4��]@cށӌa�c���j�Q��3ѓNw�XX�ф����٫Gћ�/�>�}8uj5�����Q�vy�[l���Sl~��t쫫�Ȫ�7y���?K�u\L�M�>��r7�.�9
�%���l6&|��wJ�+��,.COvh澞�y�i�ZI�sT��H��VU3Z4�{�{%��\U�_M��l���w�d��^��FnG�/>��	��b�R�x�KY�ٳ��Ӭ�S{:��M�52%\-���SRZk�%m�p��噎����s��[6��@fhrLni��Z�Lx��f�[��K4^�ɷ�M=	�]ٚ���`;��㸁]�C��U��_M\�@G��¾������A���c2j�UUv���'����7ki�;��o�I�|?m�?��P�D��Ȭ�ͺy�yY6A����ڻ�T�p䯬3�K����C�s��w��Ho������Y	���8fyw*}�got�mN�)�%[v%�1�Ü0���`���\Kr�H�k#g!�{$�9a�5�4O�#S[Hv��W�}�:OYz��ݘ�b�l��|�v'�}չ1u��KcOvb��7nL�	H(P��H�0/eo\����.���#M�J������)�<��{���K&~ݮޑ�IW���r3���X�Z���m틎[{ۣ�������E1�v^�����5̀ov�]<ih/�Ikn�4���5,�&����>��k%C��(
	���.��F�<��{Kyl��ulLO��p�������W]o�(�M�w�����?�2\��j��tYD�~rgL���6g�h7pÞq��;��1�x�Z�L�G��]1~e[�?:���!㋎��Cim�S
̖��׵�OL���z��M���6e�P�Y'�<D�*���K�t4eNk��k�Ǔ���a�/��k�������<
�_|���96gx�a:�8�ޖ	�'��ks���[O��	�O%wU��F�ݵ�hҼ��1�+�.Y�t��zzR���d���ޟ9(b�8�k�j�g_	�j�^#k5������Mt���v����EŮ-B��|�w m�0A�mG��<6/+��55L�4�pײ`&h=��9���Ld�F?�� nRgeN{� ��sn/T��Q>��c�EV�U��h�R��_>0؛�d���6[�Ov��[ڼvWP���TѧZ-�����6��9�Y/k$������o�ٳ�9���JVod�wr9S�[�{fTr���Η�	��y�o��8��'o˾�/B����m�U�Ի�,���P�nlS�"�^S=�n�[_Ыr�����0���0��畘��e�n)��������5[)BǏ9��7<9��jެ�H�:[�:V$�}��i�\��Y�GyqG�J�5���׌G��ù�n��g��L��X��J�h�h���<�dt�>���Gն�Ǳ
��������\]�7lX�������#L�Fi�":��yO���	/Rn^v@�6�������i���m�a1/�ƭh�^��Z�d�{q�ŗo2 �����������8ziE^�;���k�/����-x!y=�=��X~�r5R����=���j���՞
(���h� ��ǔ7�%Ў��W��v��H>[���}U����~b��^����_��3�k�e��'�$���4�Kd���bN���ri�{906�P���^��kW`�Ӣ���dC��np젧ٽ�������ɕ�<-胆YR,_@�g�ӣ�� i��{HU��l��ë�"i4��WCXk�5wHF�(w�5`_=UyŚT%�&�j�w�픕����Tb�c���X�ZC�G�	>�YQ�{.�P�0ͱ!�+�qO'"H�"� ��By-)d�,a������{��Q�ͫ���Ʀ̲x@�W�9�ʷ+�a��`d+��l�P��0œ���ox6��NOV��a����IzXg_���Kl�o��W՜�|��x{�V���ƪ�#��L;�UK��-�����-䒕���'��L=���Nso0܊�=\{��@�s>kx*pW��|ڗ ����y\��� ��|�@̓�ԭs�+)�m8A�n��wX9�7(��r��t�p3���'����`u�!���̉I^!ʾY�x��K�;|�f����0˦�nHc��V�n��H�I�-3c�x��#���W����9�;#�,��mH܈2�n�Y��76e�����N9�|���wv:[],�%K��fw��۷�Y���N͆�Jr�%���"�WeL��u�d�+^�
�&e)�����9�a�YQ7{�����YqN��}\%�2^_,��ڜ�_Y41�_V���5NȀ�]B�Be��0S:+�e�	*S���'gGD�gv�y`=W9(�r�}8�{���<㜏Ě��qW_w�h�+����6�'}���e�bݹݥ�dabD�t/E�$ ��U��,�}:�S��w��*�)M��Ol侰�ڙ��,�z�1��xYٯt<����{��kk�Z��+˰�p�Q����P��]��5"������e̊��\T��m�}�#=�`n���ŭ�NU��/�=�]1KOsdq��q��=�V$������E�mgF[up����i\�峩�,*�]+�h�]�����f�[�5ԕ���4�Oz��(q�ǋ��b��,ox��Cr���f�P:	�V�Џi(���f3]7��m��c�.�S��X�sv���4+ ��@A�YGsf-D(��.7+%UoV�C�f]첛@��CK�D��e���4�1��@>�Z��a�vJeCE�Ƴ0�-�7dL�vV�u���v5�����Y�A�U�R�ܨ	gT�!������iMR7c��
z>ʻ&�B��t]�-Ǹi̞�Nj�7H��ҳ):���8|��^���׼e�k��}�����G	�d2��ؼ�����Z̻:If���ק��6N]��>�м�*�4��1��]��Ր�_R����^���nʹ�uJ	T�\�ڴ-Y(���`��:��K�rt�<�}�J�9�86�t�Ӽr+��C�m��ѧ���f�E�N� �s���:M��B>JBGRԖw,��WRPi�|���BɭU�hw�v�c�o���刪�t$^E���ͧkhS�=Ki��A��=;���u�/�Zѩ��=��7)Iط�Ǹ�h�����gcOge�|� �G��_����o��l���荡[�2���e:[oE6e%FG؃���;#�Ź�	yrT�:�rX�iӈ?���K��DS��r���=��l����&�^��$@�$��^�jy��N�Ѧ9�4��㬾=�����Q�3�L�� ;�����
����5��k޵W-��U�5�%L]W��b�}Ñ����%��r�+�o�%��bP��.͜����asI2�Fl���WA˔���.�B
4�̱���u�3~�e�����Uk�fP&�+Pm
>nEj\�c���T�u�٤i4ZHBaHጰT�(W�i�@��1`�b�H"L6c�銔��&���Ė]H�^�
@�R〠�O�Hl6�&?�kH%McgkQ}ث��g]�Z�n�"��*O�~�<��_��}�����*��}�U�U���cTE4Q�h��Q�b$�����y�����������?_����H{�DE�2Ov����\Q�MxA������S1h�֭��y���|||||~�����f�}����{���tj�o�j�������#j�����ڂM[W����tF�Clc�~$|�*�[y�TU=b�C�����h;�⑚<΋cU��֝D��tv�QѶ��Q��5y�TS[h���[U�v�(�m���QUT�Ѧ�o����W�c�v7��QUأ_n�j���c��#��1R�V1��u����&��$���i���Vƈ���������]�D׆�ti��Ӽ��D�j�
*��11TD�Ѣ�"����ݚ&<�+�󻢓�	eN6���=��邫��+�oyL�N��]�Kc8ֵu[��W#�����ރ`���9��U��V�<p��૪�����:�bI$�'��4i�C�E�?]d�ܗ1A�4CE﷯�'�̾]�*�5Ih=]!��-~,҈� ��4x�1y��'���HO~�7眹�+:�n]�tHx�e��z%&�1��8�ʶ�΃�ϘD��q@N���0�ԗr�M���Yz�y�.���F�H~�$b��q�7W���X���y��=�@ffVL�q��nF�9�/8�X�o�{8� ��U���_f����)�ؚ#�#��ʀ�r|؍׻�����&�XPDu�������ڽ����n��}��XdXcֲ�a���(LiչP�[�NM��讐�A��z_8�d��M���V�I�`L�'M�������Ӽ6�<x��f�#�Q�ƙH�lL�|�5z�'��=�����^����١��o���Z�ƏbP�;�
�l��i���<d?m�e�B��<3�w�z^��W,Q��u^�Vec�����Z�h��z���HJ���������*��R��������8�Ow1�ki�N��^���I�|��--蛺vm�8���h�'u���uI �,F5W�*��+�����j���ؚ����7�
�(�������c����Z�����dwq{��iA�&^�]	�
�S��8�S�J�Ld4�5Um[y����UNwS=��Mw�<�!r�v���p��-�c�w�k�겯5�;/�9�oz�P0�'2�_���{M��Ҥ+�o�����R8Z��S�!�}�ۢ;�?�o4,�ύ��j�<wjC[�W.Bׁ��t�sb&ol�"�C���Ea� 4�,�ǋ5Ы�g1�w�k�a�+����N@�2��DP*߯ե���ĭ��)u�.����C��6N�N�C�������w�N�K��観�!ʓ(��d�ŵW���촨,�%�Y�j���{��=4��g~j8o@t���7���-7ó]C���,;���nfaԮF;�|��k�m���d�}3���b��w.�s�wVŎ��<JÁ���v	���a�3I���������*��(~�c�*༬Ơa\˭����I�I�*��v}��aw6#SD:*�<���hO�����������i��!������ϳ�Wj�(sJ����u1��SSxv�n���5�m��im���ņU��'T��θ�R�yI�3A�Sw�����/l�LѳR��cFFq��Ӕf�����8i�8��.~��dz�����N�������] V��9�V?`��S^��PPܶ9�rO�i�uvWY���_)�����T	{�Q0����1�'����6�VneU7!�7��x��{e�M��r7t@�ϱ��b�;]|�2��M�,��K�?m���<��s�<�T����Dm�����d�Rv�&ެc�''M��È
��<t��s��MS��5!.��J{y��f�d�z�41�P-j���J�k2BWuf�h�e�����Q�	�(&O]kl���4�Z����q=�>�Q�	e�$NY{B��lM[I�/P�"d��i�������N�ܳ� )��5�{h6�*enߒZ�޶G-N�t>�7K�j�rja��~���ZrR7��x�bҴطG&.۾���!s�o�p�+�^�o�M9V	U�٨8($�N{zW�~��k��p8q���r�Ge�Ve
��:QT�l^�ԫ�I��T���i�S.�ݢ�MOa�x�$w��A?�_Sêw_��K�Jr��᱕!��9q���=Vt�s�m�������Z�a�ۥ�"��.�?M��� �΍kK�ܙ���@���8�~���rkoE IwN�y72N�ď{������/��ie�Y?(�,��Vv�����":<�TzF��/r:�|��H�'wր���s[t�B'��&0r7h��soKN�Ͻ��4Zp��;C��|t{��ֲe�Hf�
x�d��"N� �ci��f���͙��k嗷x(�ݜٷI�;�k�:c��y��|���,�{��'����]��v$�D�R�5�0f=9U�֫�srFp��ԗ�[GgK<y�WuBIz��]{ 鞊�۸�����Q9^�#g���ź�ҫj�l9��D��Nk"�&"�.����&�>�g]+ʌelQX]w�0��j�Y��`Tә����SF����b�gVc��^8��x�ж}\>�ꂾ������a���%�Hn�v����>;7gץv�\#�zQ����@��:i!Fo�S�[�m�r1_=�*�׹��u���9d/��可8��*k�����0�y�u�*vϹ�$���ػ8�ze�-�P"��p�r:���ŭ�ߡ�������՛	�N�I�Xx��e���<O���l9��F����ɝź��\z}�U��-��3�)m��u���gFF���8;]u��*�"|��t���魊j�s����#�c����O�_[O&棜ݥ�����z�Du�oZ���z��Y�y�� 5��Z�_p �=suU 
��YLA��\�sA��+�RW�`<�����3�:��z��FP|j�zWb�g�%ڻ�!z���&�:ݗ$�3���}���\���lU��3Ν��\}KzG��Ŧ�r�t���؛7WW=K���nFY��y�8���;�����):�щ_{�6�K"�wlcb�i�;K��E�ih���1X���"��y㷽�tC C%�U�2ʀ�r|���wm��g�r���SOv�x�1�ٓ�Tf�e=���#�e���0��YH�Sll?1r�3��E;_VC���^��aZT'&5Z.Ǽ͘�3����%�g�9L6�VwNg6S�7�B�]/G�x�iŬ�~+��/j�2��G�ȝv�����p��n��D�x�:�{7��!qڎ0E�c����X��A�w%��0�;�ǳ�PZ�|�A��60&�U�ȩ-�;�ek�����a(Y+�#�͠��E�*��1�Z��k���B#yV5U�n��TF���ѡi@�m�(�}��*ى�W�,yz�a;g2w�b�����]Lk��UO�P2�z��b�tY��(2]�����88�O4�Uγ����L�cU6�v��u_���J�Vz����s �����[ɘ�gى� ������	���h�eP�$�f	W{>�텹�wi�d���WtmYy�q���*�=;�/Ue�*�*ޭ�����*x�7�i��8�/�su��cc��z��Xj�����B�\�����0ږ�®*'���c�m�A�a8|H�V/5�7�Kvr6^V���(t�y�wf�P�
����l:�Vӛs����ᙝ��Y�&|�y��f���)H���J�:'���W�u�|e-��7�v�7zL���^�`^�mQ�y�ڥ�Xaf�Ϻ!S�Y \�ޅ���V�,2w*�/�Jffw��pGwv6�{��c�*�%��nAR1���V�雔G��m�������f��ө� (���I����
��?o����9>kFa�H�L�>��U2�ol�8jK���$��Q����u}��F?�ö�����E��=Xs�jģ0�_�T2XF�`jw��R��IƼ^�{����7�̰ǻ�؎�N��-�m��}����t�?\�Nԃز�g�d��t���0o�����v�k��-o�*���i݃��wg�v���#14j�8���N������!����	݉gY�;���輻�H[��-�7�!���yi*�Y��Gr���ȍ�\����&���Zv/���ߋ�	�Mw?��8�q�aѝ/0ck+�A,�4�M`M�g���=�Bʈ�ۡw�,�͒�O=�Z/]\/����)�be���[0r���&G�^y�+g��������?FA�G?Y�&���qR�g�:[`K�����������׎���7J�]��6�Ws�)R�#�Y%��ٮl�J:���I#L�N�u�&��J�]����ƘM*g�ε��%�oZ�OmI�v�4�M>Oy(�^e��ΨK�+�h�&�8<z�仝R$G;�p�! !�#l���v>�^Y�b}��u�\R��R����e7�e��y�ԣ�)��D�ļ\R���`�ڧ8Ob���J��61VHWw>�W:�޶'_����D�|g�Y� ����~��[_{�>^��-l��o��]�9%�S'~���UTc��6G�#N�S>��\s#���Q-���G�k�^\]�[m[
�g�33������Pݵa�ì�Gv�d�f ��y��	����k�ooį�=ǕGt�ns[�{D�Zg���k�44>�3^જz݊��	.���ԤU�'vդq	���;X4�C��8��HR�s�3|�8�����!�:�3Ǎ���bqJ�z�}Rl�բv�x�N��5��"m�%B1��5u̙�F��=�j̻=W4ဓ�M�.4!���Vl_g�d{_o(k�pł��Kک뽼9�4�3,`Y�����{�.ou��T��7b�f��]պS4��0ȇ9]Cf�����f��EQ)_fO�X��6h2-m�J0�%F�9���J���MY�J�M׆�(�+����w[/;���-/�2p�f��eܜ�k�oK���e�:�:q*��W>"$hre�Q&�iт��D�D���{�C!e[w�/�ߌ��Re��`��m���v6�����<ļB�0� X���n"e��)��l����|�x��l�
�4�x۩����t?s��)Wz:�\Fh����Mu���2֨�P�$V)f���F�aj��ʎM��<T��2�j{���є8�lTe��`QC��/ة��F��B��w���w�J������3qU�1�e^��W�]T��8���y�����-nU~�xf�59v���rGez]�Uϟ���Ugo!�׺�]�����cZ�^k��\����{Y�/ߺ+z���>֚�䶆pq4�Q݌��SvD͌4g�r��m%��8�B�����ǣSOCpY"�`FkJΛv�<�,Ug����]
�!�޸������X��rI7��%����[��C�F�16�6ߪ�J.a��U�+����eW�r�Π7�a���z�5`��8�k�y�6�Z���,�.�پ�����w��i��mU���U4����w��x��WX�Vd�~�R4��ov�)Ft�,2{�=y��7|;���;�D5�t5}�8�e��B-��ܗpt�_�������3q�C�wXpLlJ"]f׷���U��Z�m�OQ��a�/G�La>�<����Cf
�0i��5�W��u�~9�;XY*憃���.�-U~i�:g��R}���C��l���Z����fDj�~�}��5Jk䍜��h�i�6P�~�-�ħ�K�t;��K��b7{����ɟr���=��Cn��>g���
���5eKq't�i5�<q<bA�}�x7�i"�FCe>���ma��	��1_�z����.�+���DmC�^׭ �ڷ9HE�
��f�i���X"�F�-��q�Gix�k
��7��*�`r��뿘�(Y&+j\>�iL=�Qs�{9�sl��ȣl�{oAj髝5�	+�@�]M�b�U���Zc���m^��V�m�@\ڥ���h7B^��߈߼�r!qƣ��~ծ�e4.�
[�Ӗe�����[�%�a��7��J��Mump*otJc1�eZ�ل�0����������hծ�{�������7��x��T�kv�{K/�ɲ�+�]���F���-�xӂf�]؝x����#Y��N�K�<���6�#;�69āCjfd��h�\�r=�<�V�XƮK�&N��k߲���f_8QdVҮ3kx�H�X�x���x�����-N�Tµ1�MX��(�F����zs�k����)v�g�.��lS�tx�I_s,ͱ���%C'�m��ȼ��a\� �����\�gw*�ڻ`;b���O%ٻ��P�����ى�-Q�!&��j��+H׌pk��B��(�*�^�$���3[6��K�e'owL���H�{�{��$ڔXY�����nh���}�˰#��c��Β���n��I��Z���_%��#������vb��d�	Ic��ݫ��
R��Щ[�s�ƎJ�w`92��j���m�Q�;�N�����F$X��%4,'�k��)��^,��ltl��wVJ;.Z�fʷ̝G{��a���m>ToU%�릉��(�릈[��Z7�w�rH�/�aM��s�ƀ�ݮ�T��z��׻)��Ȼ]7���&�	�r�)K.�3(n���	�5��d�Axo�Sz�X�,���n�7T�o#7A��C�-� h�(+���b��TG;�`��K%�A�E�2]��S[��K�j.���,^r�Y�͋V��pU�-|N�V:a8V���&�V�d����#;r���byr�K��)��e]Y�9W���e���Վ�P�.T�O�u�\v��4����W��f��ɢK_9�V���������]�h���#��s[k,S��5p���:|z^����t�<��E��j��o�ӱ;�������}\��@�ӝ�P��YPȦ<��a�$J�Yt��"�[�L9{-�ԏ.��8�«����e���;+.�Q�[����Ԩ�f���M���+8��˼���Y�3H^�AEm����G�(؆��uV�<Nf�X���V6�mS��&ǝ;|-�8��sыf�X�:����u.�ʃso�]j�<x��v�&9`4����;n�]�e������G��E�Gj��2��U*5&'��A�ҋ�4mݾ�EဃG�w{8m%�ʫ4\�#��7��aKr�^ujb�Uu,t���۽�K��l䓣fkɘ���Y�G;�2x^�20.��W���o(�*�+S+��k�R���Y�,�^�M^�<�_[��uvK��DHଊ 4��8E`ncA�5�1������l=a�ߞG���~_��Ψ"?1���m_�뱊-mh"j�3������cA�P������~?���������9����f�&��;g����b���h6�:���LET����<���6:����<�~?_���������}�����܍�o���gʢ֘�b��S�q�t�h���ǟ7�3O]ڢw�����~?_���������>����KN"���V�)��1kUQQUEAD7�w�l���bb�f��<'Gn�f��fh������;=w���"�4P���lb#��WZ����bb�TUUDPA0�cQUWY����A��l��>G^mMER@kKy8��mX��ӈ����"�uSN���=��LF�-4�:Ɍ�t5�;
�H���AE5b/���yI�mw[F�:�"JJ��
�:(�S]�:���UPE��P$3���^��5ݍ��z�#{q��ӺRK�+��m��s0���S��.kU�n<n=��\�+�.c��xE�4q!��~.��h��SiWN U�
�[,_M[W���4�d�B�8/���H�(�<ޗ�+7�D��St_m{��O�ݙu���~B��7�"Za�5�Ѕp���=��"ZYVUugD��ؼ����+7�u�����d�X.���f���[��*�F�sZ�Tn���5��)ݟ^p�W8�t/(~xu9!��u���q�IL�Xc񣕋f�m8��Go�<'"!�h�d� ��N�5�޺��"
5<���.����w
���</��q.P7�����j���l������k#_����]^^N�W�n�����H�3��u��q���c��N�VUNb�w�>qd��v1��i��I�8�8��Fl[�v�\v���o��q(����w@oR9e��oGQ�8ЎU�,Ԋ����'i��Ȱe�V֝�����;MGwNfo���ɼ�����4Z��:��=�������L�1z��Kϖgx�𱧗���Gi\�m�����G�)��GX6+���3�W:JLe���}6�I����no�2e��(l%��d��Ea���]��f. �ٙ̦Xe�J��:.D��yM��M��E�{*�ޱW3us{ �6�s.��s��WDu1��1��0�QR5[22�ڎ9�T�{51>�~����b�wA]ɠx���[q��Т��f:�UC�8؉2�wLSy.�<)GM��7����c�k�L�i7+��E]�y�[&�����t���B�zGz�yF�|��p�.�$@���<����U��V]ҝ����[؛�����ʥ�9e���"�qh��;^�a�V8��nħf��q�kk�������s+���x�M,��aQ�k�&�[\�3�WD="��.�d�*w�D��g�Խ 25���F|��/�1�:�MLmD3�R���^�t��:�$J����[������T���k�3W����o��x�ǎ���$����3����������彣�M�7\Ȣ�'�՛��7����ħ:��<����Cq��+�&���تp|d�aN���-���or�����T�f�g7�&w\Togv��i�:���ok��UuA�ݴgL�:A�gS�1R-T��aM��`B?xxe#�*�i��guޞ Dy�պ�+��zgM{��u�wVZG����|��[M���3���鳻�*���&�3�b:<�݄��y�M�=I;��Oc�y,.r��z�NK£���9���E;��w��']\5�=�u
I�hk}�w�['Xg?.s��q���v���j�㏡�!��O�+ Ϩ_@�F���&�գK�m�f�n��gk�� ��I�2���vC"����V.:)&�Nyݏo���K��a���@����4#�&�6�GCl{�����}���R�P�Y��
��cĐu���1C�z<����צk�4�;-�^:56
7�x��-d�Qz��[U=~I��	���z�������w/�n�E��t� �>;rA΂f��w(��Y
�؁�jh��nS��`ʲ��j�x�>N���Ur��|*K;4�Y�N��$d��*�~1����Z�U������X��X�˾Z,���.�@'Cܪr��V�b>G.��~�g;�"*��^�*��4j|�G����5��t��\i�b��y��Щ�f��t#��hI�m<ov��|�n�-#[���5�$o��r�=ο}U����𹙝�.���R
���iR�0�K�[������!�$lucm����`�{����NZ��w�7�޽C�s��*��&iv�<�7C�g{k~��v�$��k�&����u�\�Y]�*�
KG����:4E����Ҍ�s���"ߠN���W��G)N��5���%gQ�BO	�����Vi��3O����E/-�|���)DJ���	��4ƦS��+�h7>ٽ�<k�Y����ڤ>���b5(��Ι�%s�u{{�iĈ��]���60S_vޕoq���#�G o4�w�`y�#ͼ�Ȧ��Y�V�p}���P�;�K%喝�t;Z�.�j���z��-�dx�\+;�4���6�nśރ&��	7ӑkGOs��ݎ��<�+����=�]�}������~���ڪ��+�G��~6��L��Y�OV߶f���ɹ�{���.a�#L ۃ:�5���Em��v�b�5I-檔����so�a��m�]2IYH��W4e;S_r[������ޑ��K"ФȤ�?�}Ib�S�~bS.\���M��V����xC����pCo��Z�`<Q��W_���Z�o�e<�xfu[0�iw��Tr��޽��ƪg[x^�Ԁ��VXD�X��
�H�ϑC�{-�]�2���wَ�I1l���멝H�UHz�F�{~�$~����s=�i8��|�,�z�(�n/r[[bL�U3�&D��<"_�쎪�j�cqC���V��0�����,��?E�5Q��;G$�7�fQT�V�,���{�Öӗ˧�n4đj���[�,�R/�nsj���;����\13V��Xzq.�m�]�+-��%�fh+t�Y����0*��{�:�u:��<3�6�� ��5���@;Ը�G�Ffa5Z'^2�XeTԞ�!�l6NO���s�9�>���t���l�~��˳�3��ϫ�y��{��l?(�d�3����-�.Q��?AR`�yO���x����&�Y�.��;��ޤ��]��K��&�s:J�U�9���*���E�,�W6_g_Ϧ�Q3�}
���ﷃ��뇿���^X���H>��4�G��|˵�K���fk����3p�v�����ӧ����3�.��Τ+ݺ����^��6�ߠG���.���]d�ea�59��R`�U`�ӕ��&v4�>�aa���)1�D�s�����5�x�t��@`�Y,@l���H�h����OV��1$���q��i��}D�f�͍�u�8�����r��,��϶��n�L��M�"(ޙ��._z��������i��kO���U����s��-V�s
+iV�6�\؃�P�8s
�,gSj`E�iw�M\�]��v��c�=_^�Á�}��lo�Psڱ�<�4��.r�U㱚�I�n��s#��,�{*/�_MϖP''(i�X��Kl5WsÍlj�>�x'�[Ӥ����J3b������
�op9	P��)]��ȋhfp[,.�׈E+�]u�u��ŵG���\�C�V_��v��*�8�4��{�F�Wۺ>WJI�W|����k^;7C��7y�x+���W�>1��K<#Y���6�����i���h��Fp$\+S�ʫܭ��FH�}�� N��QM���L�i�L��	�z��������C�{�6�����U�9�����Skt�#E�L�1�A!$m0���6�����v���!&��V�<��5U��kq��+f�q\Z1O��?-��z[p{gFd�j��l�{�W�>1Mv¤���N:ǋ睳�r�'X\e�������s�A�8-r6�\��9!���cT�y��'����kTm��=i���y�碀�K���V+�7}�D2ہ��T�aj���>w��+�U��5n��ue��v�}XCs������m��g9���Ȟ3�z}bg�bLgmU�'^��/�y�)ɶ۳MX����N����Gר<�a�h�aIP��f��U�3��w�i��@�U������j�����jg3��u�d�d@W�/�[��iGb5��y~ؘ�̛�9s�oܫ�t3�mf�n���Vf,�Z:���^KZ$i1O��IS8����H�9Jk�Ԍ�g��KŎ���]v��7��Q��bB#�Ǿ�e�����(�k�(3�9+H��*­�+x�R����B��i�7)Z�N^d�I&�(d�4���ۭ��l������/}�e�[}dݍk�@���qgC��5��8g���Z/�R��>�ms�98p�Ή��������7}�='y�U]в��g�D�"��P1S4 z�H�l<���s��WV����s�F���i��ܻ��ۄ�}T�u��	縭�u���_*Ev%rc�_w��K�9�lT����⻖����0� �u}��U.�W/��0�pu�5��{�fEc�`*�U�}7!'��k��s�ű��sQ�K��3r8ݪS��;�2�f�,}tT�p�墝owT<���F��R�U��ޞ{��t ��"f���":�j��1���9(��+���{��Z�>��-�3L��� nnT1�;��G\J�j�#g�3�J޾E���I�N���*��̃.�~ǎ�-�Gw��瘾ؾ��" �T���+6|6��&��s
t<��:ۂx�;o�#H�إ�{�=P��G,���21+"ֱ����fn�1��(�zc�	{,n�6����W��,���n�ȱ��m��he�)el�[tk�~Ӈ�,/n�޿��9����xk�>04�M�b�˸��kr�gw�kǹ1�π��j�O�q�ˊ�50�O*uq�������s ��:el�a6򸧩�Z{ז��y�J�u��[�DONglmiڮH�mv��7g�o�=�'�U��;p��z�Y�z���~��6R	��l��>�hNc�Xn��@�l2���4���e6a�Q8�=] �.�g��@�x7�x�#޳^n����������,e��䂉2ļG #�z�g��m�K��;�6����N�,!�E��G�1n�|0f�'��Q�}��Z�}��8g��⊁��X�u�a�t/q�3�YH�8���?~�*�u7�`�|�!trM�#�ﳽ�R%jW����˗�L�/]�ec��n��q\����8F(�[�7`�i[ ܕ��UwBRp��w�V�@[-���w��3�U���	��>~ح;k ]���	+�ԉ��5+0�٭{��$�-"��t}����Z���Mx�ˑS�)�L�w��3��P뷚��w,P%囇6�g;6�}L�TǊ ����ܻ7���gj�";E����7ك�I���f��n���g�cbP�<��}sǜ�Cs2�@�״ �;�ĝ�	L\Y˒;c��Up��gr7�+v��ӏY]M�{ȃ9��)֫����W��&�[����k�ɿT'��1��.6��Q��6 7��,:�-�R��eٙ����tC�6aq�q�))��FƧ1^�ߡsěk�����m#�{�7o�B�{Y��p��c���+.�>��e�[_o	\8���-I�f���bk2���4��6�y��3��˴d����y��Ĩd��0��;��x�>ɝ&[�w��	�����l�]�&G�-j�]t�T7_ͦ�;�Vu��,wi��°�k����9��]^��|ד��B���	������V^2e]�F�1��fx>5�g���nK��Pá�<D�x�X0`T�<�S4'i�Ȟx�6�h]P�� �B<8Ё�1�1�Kն{)K[+�����ẉ�
 �>qAG������AF{(8�(�n��>hQ��CCC 0� ��@��!��2*2� �0)2C"2�!2�4ʀ� �y�2 !B ��%@�� �_%!�B	��"�~��� ��@>J
�D�!Ty���� ��E �C"�l��p�!*�B(!�B�!�B�!*�B(!
�@��B���H���B��"B��J ! �B�! �B�! �B�! �B�!(�B�J�����B�@$!
��B	B�! �!
�B�H$4�B!!�)!"40� �2)@�! ���B�H$! ��B�C ����C"��C2)J$4
BJ$!(�� ������|���������PQR`;�	��5���1�=�S��_��7�9�?�ˁ8�:�g��z�ή�DW�;>��� Q|�0�*� |���b���B���y�_w ߩ�jQ!g`uw�����T	��!�$��,�����I(�	�A �J$B@$��HB$"C(��C��	�2		 ���)(��H)$�B�$*�)�$"@�	2�H$���	"J$�� �$� �"C��	 J%"�BB�@$��J@�0,�#(� �,H1
4��*J"���!��(T(�B��J(� R!�P"&$B`I�A&D%�H$B���dBT��X����[�D���(�"�@�R""F��	��q߸"?�9��c��A@h�5见��K��T�����wjT��@s(xӣcM
�*�T@z����a�@E���������%�ڒj�a�F(���&ѡhv5
P*�*��>��� �
�C	�/����q
��7��`���x`e U����@w���ШD&��RM �'�C�i����� ��� �
�K�D0j���*@P?]�2g�w  ��X	�� ��z�{l�:BP�;1AY&SY	���p�ـ`P��3'� b@��TD��%$*��"�%@ ���"��R�UTQ*T�))P*J%RAUJBH)"B���A%AAREQ)PJ�R�QJ��D�D���*)HJ��"R���T��*�U$��@��T$�Q	$�EH�f��)"� *P� 	B�UR* %BR%J�":4�U
�IT�UTRURA@U*�%T� �"$U"�;���U%n   ��GL��e`֊4�eel�CU������[L�)�mA`�4� �԰�adR�e
Z�)��l)��T�ATJk$Q*T(�  �
(P�����â�B�
��СB�
AgW�m��e��,�M�dAjVl�0V4 �X�V��)K)Z�Ul*�0R)T�������  6�R��KM�ƥ@����UHi�`ƅ)Y�R��jѪieMMeP ������)�f+kVԫam�Fl����%Q*��2�$)U� N��ڒ��6ʴ)UT�����2X�� m`��Z�@��@��(kJ�Z1�����%TQR�*�J�  :��A�,PM��CmUcbJAJ�ej&�eB���0�B� ��0 R�� *��(R�*RTD�(  u�lƦ5 P!IJP�2�EUeLUQ-��ʫm��T)ZVђJ� ��%�P$ZR)��%*��	W  r��Ҙ��2�@K�]�:�:`�)��� ����C�6�, r]�c��u�4�*�!BH���Ux  �=�
p�:��
 �`�Q�S  ��w 
(0v  �[�n� ��e� ��p�Mq(EQR���UW�  �<� Ҝ:�  X�@�X ӸU��;�-�4 GqX ��&)�P8c� kp3� ��AI
Q)JU%$��<   m8���  M09@`@  C� 
`�J ;�`� �n�

�0  &Gn� ���R�! B)�IIT�@ �)�<� i�  ���R�  �)��j�� i"��  �Jeeb.`n=�%3w�+(���E	"%T/S�.�v����ח���0BN�>��0BN�$�HH~��$����� �!$HI$$<���֍h{����C/m�t��;�a��	3BEI�1���͠��.�cZfk��.�,�ڡ�0�Y�Kbҹqt��r�����.g�ka�n�m;J7a�V%��`��sB�03#N�
�#k75H`:��f�Z�!X:!�'�cd�&�6��X2oؖlKPV�7$��֌1�*7z��ơõ�,�mܹ�1�-^�#qY��M�*���'N����<�%Q��2ۺ4m�zq�L��R�Xb�^�f��lj�d��(qXA����HL��%�nd�� ��0��kt`�+f�	uS7z�:!�\u�Z��q��p�f��@���D�$@Щu�푔u�&]h{��؟�N��O~,�m���ͼf^���LS�ۻ���k`a�;W��)��5LF]=s �`p���Ӵė��@�r���T���إ\b�2VUA𥮥i��N�\Y�׫]����e�Λɛ�Z,X��Xщދ	fd�(�7��;Z�^$vqf�[�A/4B%Ƣ�x�AҺ� Md��B�9c-���v$��Cg6RQ�`|�-Z��^����֯7[�����3v��.MOW�5S5��,����l�t�P&l���*��%t�F�@�ˉ.d���W�h��T��-��[8b�X�˺%�]��حLRdIB�ՀE�ʴ)V�5,�CB*j[Jā
J��f�B^S�����O&!��`ˀ�(�U�meA���(m�t��7���b���mf<&[T��ܽ�ѻ�k5,R3�;H��B�Ō��YSiJ��	0C�`�l�{I�Rn�f�Z�%��X�#NQ��A�y����n�N��l��6V����&K�m>B��z�k01��J����s+*0��ڭԒ��%5�yvd��z�M:�̰�q �Ko`s�d!˗�6gݗugv!f��GJ��`��V�ZZ��)�O�b�&��;���:�] �*�Ig
��pf�-!%R��+qVJѩ�˽7"e�
�|��1-�ڧ.HŁ+I3+��TW����� b:�PŃLa��,��{�Y� �������)�U�Yul*��)���N��,�/1�%P[�l��J�������H��ܳYn�ݲ~�qU���n�[��t]uAV�
a�"�d!�1Еj�2"uK��ˡ9�V��j)�IZ�\��i-�e\�Z�a���rZ!���(a�aƲ˙Mj�W���2e%�񬽳Vq;Q��*��4�`���q�9a��hm�Z�*��<j���ib96=�6O��SE�X�eg�+��[z[˙/-�q%4ی�=���y��7�LSc�Sq7j�dn� r�!2��Y��x���,+�Z�3Qj��iv�5a��1��]�b=xhfB�ߢ��0b)͙�&\��M��J�J�Լ�(�u
+)�l�T{����k��#N�%&���1f���h�Mҽ���ĵY����@�QS4�ԝ����kPԦ]�*J�#9	XD.���ط^�L<���A�TfkC�����ڲ#����U�����[�����{R@ª�%�߲%��J�sV(^T��e)[% F: mkˊ*C����r`{���b�)�s6�͒��Ќ-�Di�۬Բ-�W�R[�`cE��2�\�[���X��+e��T������#H����f�k�I�ʹ��K4��i�A=�tH�L[���{�QV�=d-�%��|+��|���c{X�v�0\p����1X�H�,�6�+�	�.������n��f;X�41C-j��)��r
Æ�]6�l7;�%o8�M�z��c�i��*�d�Z��r����C��46�I{Zl�2�����Gh�j���
�n\���K(ѧ�F�8�y*!D��I`rݺ��@)h��S5��Y��^�;e��A�z�ͼȳ脔���%ݛ9I\Փ40.!X�4�B�yo-ժy.�R�N(���X�ItR���u1顔��d�"l�!0�c�.����Xm�,l���� Z��PSea�ƹKS2�����Y:�-�u�:��*7
Aj��K�o7j%��`v�&��J��T��t�MB�^[R�تP����h��eI7q�f���YSv�H_� Q+p��UaCmYm��P,�͠��b�j�������5�%@��f޼�qc��P��/1�d����)4fY�p䙇(<x.����SoY�H���A�{�:9;�dCR���L&�
�[6^l��C%G*!�$,�R��Gtz�ZXEf�V�)Դ��`;ʴ�^BJu.�^F��	8���M3q�,��Y�VG�+ʺf�d� �Q��-�j�z�p^�r��6�c��L!7Zrۃpf��j���oe��CF�	[�ޤ%�Y�[����a�>D6�3)m�9XkYm˕��!#�m�e�|k3n;�T�-��Z�]��D�w@�Z�jP���R�K7(^�6�z44F�)�h��Vf�Ҩ���B�"��eh�����E
�V��whn��ì<k���Y�[��Á�fDu��wR�׻b�ˑ�[�b�U$�l+O71�S���I���((�"+h ��7H:��q,j</B��\)^}�n'@F.�������v�v*�v3�V"��Ȕ̗�e�X��ٔn�ٹO)S�^�T����B��Y@Yil�]
�Y+u���Jn�d-8U�\JTJ�\;�颞2���3"�s)�KYh��{�AI��n�E�m�4"݁TL���[{X��wF�tCGe)Fǖ�P޽*��h6D����KiU�F���.}
�ӡ�m^�jm�g	��7��|����y�۴R���cJ.���4ۍ1y5:v��$�c���a7#a��X�9,��=hӰtΘv7����J���7h¬�o,�j�yM�wIL���9wbR
�T{a�E�L�j��RN�!hn��sm������WSi:�Ĳ�.R�h��]ټ�;܈nXI��+&�n���P�4U��R)[����з�2�4w2ʭ��)u{y�Q�����V��S㧱(Ji�9��(�V��!P��0��X"VqyR�V�j�W�_���҅�E6h#zv��c�H.#-�4:�4.�Y�s`�*Y� �黪�7>�S'�b�cUmm8c��]�ش��n�n��Ԙ���\N��5
j^��g�3,���Q�Vr�@۵���n�WgS��ȉ���T���^�q�O$j��-7kL������h)�n�Y�7a4��2����[��⩚ ��,:��g�P�ֵ���nXn�$B��I�T��8�z���Ժ�)���$פ[SKDZ� [5�`�'�����E,�G������_L��M�e��C.�s�T�R*�(P:�׀��ŭ4�.K���+k2�7b�ٙ)�%��M�CD�[4#3���Ɛ�`nֻ@ˤ��0��l����{`a���)�[�9�1+͎S��,�(��j܀ݢ7lMh�U�E��m���Sn�&�]��/��tk!���8�J3]�o6򠺽��Z5�)�R��7Wn{�c�'��`�^l�n4J�.��2ҍԻh��P˗�x�`��Ӌ\ı��/��ur��X�l�O-h%�i��L�u��g�䠢��%m�"�QM��&kmf��[5�B��o6���R�(e����L�ap'B��H+�'-kv��`Vo"ְ:�Kwn�([:�ʒ�ynPˋ �X{������1�dRtvP40�o+bq妴ѫ�$�vi;Z[l(s$��݌w�i��b[�.�q�[��"]�[j�F��d.f�򃶠/�YF�6�t]��7n�M<����$i5ٍ^3�����m,���U'x�S��"0c���v��Y�s$���.�p��j
'���N�����k�jv1��T��u�N�UN�)��� ;��D��p�I4^n�{u�c˱�Zr���$���1*8�5�i��1��7���w�*�h lBH��(��f�^*����k��n]jK-m
���2�f�`U�J�5��G�-���)D���7Yr�"��)�S������t��V�&����%b��=sk(��:nd��f��GE��hëc�.�Q�{QS�s93XT�	�&��m�t��k[�cǍ�8U�*^^ㅺ�t�ԉU��]�m�6GG~�r��`!KfjZ଑Ld\�xl(�E��6�!�L��ҁ����Q(�K獓�N]�6~�.�r�ѩe�o%:I� ��@Y�'����%��(C�e��	����#)��0�l1���7إZMҦ쁒Plmf�KrzrGp�a�N��1`�ы,�ҕ��5kT1�qG���Tub�Ɩւ��Tx(��R��V���T�2ȫ����(�����LX�"����[qm�4ΒX�wi�Q
����6���X����J6�6��h��<Xں,��m�Z6�sBsToJ˻ߦ:�I�ne�S�o75[�v��aZ"9)�Ih"�f �(k�� ���A	��7�w*��3-�ٕ�^;����K�v�>kI�w@��������0��P�)���r���Q:�,tq^lTځn*�J�%6�řZ賎ɘ�c)a���X*�5�3��ż��JщVh��+Xi��-�8CnD`�yfm�qa�Dh�/F��n�ci�Vj(7o@owju��̺��',ͽ(@�ͼ��BSaV뭵FӺ�����)C�ި��S���X�9Hn=�rӳ;������Gal�0�YL�^I��޵#ߣ��f��2��G�1��'f�{�M�0�ט���+hVYݤ�wf)>Y��*�kP��X^�&�� ջ܏I���^�:W��0��Y4�c��1��i<g],�������+-U��@�:��7km�ۆ#�Zz�`CČͼ�d�v�lC.�6�%j�{�
^kt`H2���[an'0>���Jg5�<���F8���V���6�n�,�v�LA����q��@D�4]ju-+�Y졆%(�x�b�xl e���m"�%MӮμ���I��jIV�K�Af�$Q=�H�����i��H,Y�Ѩq�4hh�sd¶K�ϯ$0�r��ڀm�%�V$�c*��GB��+LLf���x1INL��� �e־���5�t"�LV��z��՚sh��V"9f�.̩�m	JG�ѹ)^n�>Qcr]34=NU���+4�)����C+6�z�p��.�W(nQ��#/�n�ц�!�əi ��L�w���AJ��qVXp��r�)�!�!�46��h�2�Vu�N��0f���7v������ QH�[�B�
��b-�]Yn�r-�#0J�n����G��ح�f�ӵ0��h�b�����������hnH�EJ���+���3W̩�ol��p$'��#v-A��F,�)?��38�2�g]Fl,�,�t���Fʬ`^�aR�M�j`ڔ);K^�����׹	O-���܅�
��c��70�S�n�LVܽ�R��$�v��#�;��2��T�n��/]���Y�H٧x�,j*��5�t�n�Q��lI8,�#�݃�71M�Y�c����q9��c�B˺��T��V�j������/�:��2�@�s�f�l�]���h�77n�TbS���A7���)�����U*]��չ-'��miT�i4v�˟<�C���֋�F ��q<��:-mfIv�����ff/��d2�Y��(�(�?)��i�!�t$��`"�ί�˼{���U���	aU*��	!n�f��2+�LG�$.��0}f��f�ڗnK�V����r��I��(UՃ�R����`�O0̙����'�'�m��&NA�0[����z	Ŕ��W�J��mI������uc/0c��H�B�j̹H��k^ ��CQ�72���Vu8�����7��J��yx,�JƖ�ё�Rm-�&�5�YIdZ>�`����V�������ĬD��{K����F�]���j$Ƞ�Mub��Ѥ�/���(�����YD�� J�n������t:���MXn��Z42�Z�1�֯Z³o&��ƍR����p�(Z�����#hVȳt��W���^�ͳ�kj�U���y�o2'�r-bx6&1��!���J"Ș]�V��iQ��PӹX7h�K��t%�6�?�� �5�RSkv���hZڥ�K��I��f�iҤ�X��CZ�ku�^��{ ��i^���Kf�eA-��E�1�	�q���8wRcuk)���Z�*L�pV9Sv�m��ܢ/V�c��ѓCX��Htv�5��lF��5e8V����r-��´�4��W���3���N��c�aܗxZ�֊U*���.���⺚0�u�ߙ�0�n6kXW�3L���^��̻���,��AEi��e�[ώ�U�JG3C�˨P���*V���\Q��jy��Ln�06��t3Q���	��ު1EN�z��(��cc��@���-x�-�j�HҚ3v�L���*�h���B����`��7iH�@�j:9�vi\t9k/�0�[#�&Vэ!0e�+�V㷐ma�X2�k-��D��t����#p��	�l ��qɎ��:hS&�9�oq��	j+�V��e��t�p؏ ��L�����2G�+��b���ܲ\υ��w����(nn�*en[��ޠ�IQ�i�(��p��v�ܐ@�L����Vgؐj��`�V�^=��*Z`�XtӡQVo�h`Ri��]:�z4��)�qU�c/�:t��Z�wl�y&�s+k,j7D���n�09#S��	nN!k�mܺ�:���^��	N�&n�s�]A�V�xrS8��8g.D��}Qn܎u�K%s]��Փrk}+���r��g>��6�J�]�x�+��r��ј�]��s��	�r�G;pZ5�=�2��9��c�ٴ­k��r�g��v�^�Sm�jK�}tF�9��b�)�Ǽe]!�t����t��|6-����2�;�A��UӐ�l4{/��$$Sˬ��p��h���^;��u�#�nbNZ�l�����
��mu�����u�z����,��&��J�5�U���K*le	��Lѓ
��Ӵ�F\�]��Y՘n��_+����TM��ḋ���|�GW�vb뙮iӝ-츟R��������E,��wS��守�g�*M`�H�y�E9%U�f��˰c[z7)G���o���qT��z7*>Y��o�:ѵw�����ۺ	���\�פ��Q^І��v�������:��
�U��EjLjU|��.�ћ[WqXAYEdH�J�n'�ϝ���q5[�[�0�<��Z0<6�;_Ĳ�Q�.��-0
=�܇,:�0��T�wZ�%S�U�s��v_X/;����ބw]:�9öo�B,���5C��ꗃ9��Ǖ2׹;{5ST�*s1��+2VZ�<���]yN����	g�nӾ��:.�O�`E҉:rͤ:�w++����)��	LVF�Wo(q��w�M;�-�fm>�����%"�2h�guM穡4uPr1J��9Zw�d�Ѿ�Q��v�2���3�'w'��B�V9ͤ�/�Q�ƻ�F�����@��m�l��U�8���}�E��35MPŅṆ{��NZA��k��瀁����7���p>�k+��p��Ǚ�la���q�.�Vią�n���i�=��opP��+ѕ�p㾡|�r�(i��o�L�4]�F���Z0��s�͛�Y\���m��\{�)t�ݡ�(���I��U{mv��@�bg��꘥i��e��5��l�m1Հ�b�t��L����&s����U�n�f�Vv��Wt�(+b�MP�j����c��1ܝ�=f�wl��w��x���_hs �� ���,K�k�Uϔ�7͐�sH�(�Q?KX���7�g�W��GkI�Z��#�>�B�����r�a�X�\3q�OG/"H	��W�iQ�۰�&� �4�:�aֵn���<b�U�����-��k�wJ���7|�)CR����R�U׺&s SVrJ���;�m.�8����P�;#�1�職&bi`/�Y��f�4.��ڌ2;���u 4�g��\*�Q�9�|�ٵ�+5������y�&W:�uݱ<A��PbK�ʹ7�1�ō�vzɫ����Cib��n��8J��
9�(@�5)"Q0;2�4�4���Y�6ɣ�9d�v�����dj���t��J��X,��U�<z֮�޲7{����[�.����}���Fmt�z��p;�oKwM���J�dou*���p��J�2�J�3���!��
ĕ�h#װȐ�^�Ϯ	|qK��(-�شI�Z��ySn�5/L��I�@�����E�n�m*������C/H-v 4Ʃ�q�Q�x�~Ɠ�:�z_t��yK7w��������"8,"��[�ȭ]�9o���D ����0��Fc���1s����Eej��%wgS�a'�S*�9C����j�q^��Hx�i�cf�V�p9ٱ��@��D���ꎰ�y��WZ��X�|VI*�rr�ݕg�&n�Ʈ���"���"����z��V���]M}c��|;5�+���I�kw�%:�0.F���zIbO���m�T ��ZF����̧���}e�h�L[<oh�v�1����La��k&��-(s����oe���Ue,�`�N3��p��V�Q6Ѭ��N��6�ё)�C3l��(b�_ck_sa�<7*�9�q�n�R�ۢ�Ml��9dM-W�,��LfR��	��ûy���EM+B&ok�u��enFp�_�T4׽�5�qL���-�����`R��s�r�� ˮt���1��9�:B2��Z��ڬ��=1֫�:wEj2%%���"�-�	�1�^S�m�7���bԹ.�)F��Է�|����兪B��K��KϺ�0GfC��x���܀��d����fv��{r��k8�]pNg~�NGK��׸Rr;���}\�4�9�`��q���x�3�M(�6����.4[t�������5m��匍) ����Q�f�S\4Y��5�H/�L�"Z�)�=�1X/�P�ľ�W]W�ȉhL�ք�4	��:��vl�uӦeCOj���v�����S�0$;]�JU��{�U3���P����ü V�3+&w[L�����]���^4��u��z�����\��4��_mL�ԘGV�&�4���V��/ws|�t�TQ��Mޖ6cն���Q�j����:h��"��k0_,���^�ouct��|��t�φiMt�ؓ�<��/��XD�,>���~�4]���ݽA�OS�|����y�[Ÿڽ�e�s�\u\4M]�97{K���;�to���m�Z�9p�v�9%�t�ӽ��X��_.߮ɬY���q_<�����
d�5׀p*��
���>pgn�$n�-��/J��1A�1��րJތ����vˠ��:#�ep@�t�w�,m�U:ȩ�[���V)�T˄`W��*�C���خT�g���"��wWwk3�8Um.7��N���iju �����n��u�W\���J�j���m��"�{w.�vP�	'�(�,�X�"�;��_>'�R�,�}+�Y��]��]Ҧ0�2v���NP�Mm���dnuZ�
�<}2�����8�#!f��7�9���YX�GZQh}R�<a��eob�*�k4�6{{��3�#}n������ld#�U�{��XaD�m�TZ�%p��{�d�kwVI�U�E�9��V٭X	�)&�2Q]�A��\�����������	��+z�b,C��tFu���!�Y\QΨ^ea��
�b����υ���h`���eL��s����]0L do���>��v�9Y��Q�:��z���U�P��tg.>���x.6 ��({��-_e�c(��n ��f��WA��L���vg�fS�����0)���wPC��cǛi-��}V�p�p,���V�x�o=��1ˀ�錢��]�ۛjLݷ�%%�]��h-�֤��S���L!��l��|_ru�z��<�p����K+���N�6q���kk��+Z�N'D�l���7o�cҟ]j��ma�ݧ]w�鮜F���� 	j�m����+�\e}�^�l28S��}c�>�ک��՝K���<����� �O��Yr�ׯ~Ǔ,��ҙ��q� Tl���<���'����/*�ؚO{�X|��%:��������sz���ҝg�ʠ;I�V�Nh9�Br���9ѭb���4k�C����zǢ)���k3;��Cn���}H&�kf�M�(4Ե��d9���1.�pf��p"�fb}�o�^�h4�n�qR��Q���^�؞�C]�Hi2B�V��]��Y[q����[2\n����5�c�����U�%���e�;+8JA�{#A��5�^u�,�"8�Zt8y�ָc�:�s����[�*t��)cט[R�r0Eu��Q������B��Y0r�6Iq=Z��|%e�Z���i�6�;x�d&�2wg`�զBT��Vı��m.6īށE�w��nn�n��]�Dw��],Q��7+P �x�n�
�uw���7f���2����3	y3��v�s�-F��h)�+�a�ӕvL�xqu��k��w���l���ׅ�;u�k,�Q�+��v{q0�u��;z*����$|�NVn�o�&���V'u
�G��=�F��NX+n�x%�{�uYYkkY^m3B�6���ۻd.�\��u���D�2�f'$�޴g�Ob�/�@�X���G@�e�����c�E�s�h��r� V}7&�^�3A�B�Jǭ��\��IeOF�v+���u7����ɯ.�}�Z;;�D��4z�͏1�N�e�Sa�nTVb�Ҕ�X����hi���U��N�v�<��a�_[���V�S�-
wS�#�0�m8a E^��K��6tZ�u/V<��%�\2��-q�k���۬Q�M��-�s��
G4�xJ���;���ڷ�iV5mNcbv��4���ь�_G����v�������X���CqN={qcW��1Mg{yJ��)vV&�I%*��V�;ee�*�=� 4�{^+x)1�k�	�9��F��67%���ej�8��K�钇[l��N���R9\;���K:er,�)�;ԡ˭�c;S��_�
	s���-��Q\BN���oo
�wV-� I�������R���u����o���&/�5w����k�xѭ��$�	1��2\�;�8�J|�q���]�ad�B�݆�Ev���MЮKN��7��WQ�2Z�T{O�� :���.��
T�7�:t;Fo=��e^�e�mC���>-�m(�:3���$k4;/�N\�w>�4:�=#�b�߬��݋,D,���]�ʏU34����B
ڸjeL�,��K]Hk	�P����Y����|�ulR��jb�=�!N����=�o�3���5�H�;z����-��'kN�(�F{z�D��t�m�X�(H&�e-�V�9�z&�ڀ���:���I�isY�M��p'�/N>�O:#��3�+YPH���/�ϳ����CM�Mf���8�хV&R�YV��v�)h�4j��j�+-m�#lh3��TWs�:.���F��;���r*x�;jqZ+���U(�ݗa�R"��mc��M��&<Ν���].���â��QIףx'Ye������5k�w�ƼO���cu�4U��t�ӳ{�v�@�X�q
k����-�:R��0��c� "p	[��,]�%{|;��˫Z1�:�:R�SZW�k0��E���j&�Ӱ2M��ȸů�i�o{N;���0��ҫq��x>JVr,K��o���[��nc���̑rٯ��.q��"��Y$�:�_C��z�w�eqc(��%��YOS��I��t�v�5��u�uy�G�]*+t�(cr��!��]�����I3-�� ����pp��t��H�q��DQ���D��gn���9Ӄ�Xy[�G*����r�I����c��\�v��Ϋ�{f�EN�^��W�����%��9�)P��_yǶb��X�4�xO6� �FY�4*{&���cK�_`�����ԫ��Ά곫]��A<s+���C���2dܮf���{>!1��G���6B�e��b��Ҡ�f�+K9KxX��x]ued���l�;6�Q#�햝-��j�Έ�����Pt�f�=Wg8v�U�C/!�Zs��pL��_v�W'��s�qv�˫<\o.44�J�[��Jox0����g2��ݔ�X��k�es��V�MZBs~NWoQ�����1kx�og;h<�r��A�<��j��1ّ+��q�	���j����wj^��k��4[�;7�й ����?u*����NnmL��Fu�Ym�!G�nVau�GRN�����f"�j�0W�l]u[�$�p�\X��xs�T
�v]%wcon�5!w;��U3Z�j�Zҧ �.�s֣h`.��w�Y+��ټ :,���̨��+wtr�|]�}Ԧ��r=�%ZJ�F{���J���Z�Z�`���4�&!D�e��������.���� �Q��Nc��Gls�ѡ���Zv)AY���U�N��-�ōZ���܁C¾�pͥ�m<��-�=�a���(�N��υAKQi 
� 1�\+t�N�y�5]*��sa��7�����d�8szν[yZ���6����xW���T���w*]O�43��gG�+���_u�㮤rg=�U+�h�� E�J�ude �;8�f]>�g8~;�B�]a���imhߟv=teM���G�{hK"M�!}ZV��싆�ܥ���3p%���A�����#�L��8)G�,<	�f;�/�h�,V�e�u��뇱Z7����-߅-�: �.��a G�2�L2�:u�c��-��d*�vQ�Ոl�.�Sa+�e�sX�=��#.��ι\m��/`�C;�v��<��A�#�e��tlaK��,��J|7���vK�i�ۜN�kM�3ĳ?f��}q���Yo��᮵Y���T.��j-t�̏[�*1�N��PGe-9����������k�S�Pn+�Le����t��b@���/.�T�FN:Xp�*��v�7��$�x/3(+�&|̈:��@�
co-mʴ���|++d��O�N�:���|;�,-*�=��ӕ
��u<�5�k/KW�('�.fN���iKV]�oF��=,5jUg�W)z�E�;v�@x�>9�)K�A\�My��g��$��nf�JJ��*Cΰ�́$.<�v����]f��ѩBIO�����oDEw	�ۭ��aI�zdZ5g1�8A$�����8��V���쒛y��4w��[��;��h�;E�(P���"WZ����V[������"��[��mg ��4;͙w�25ǲ�8����.�.=K�2�so��̇�^@�ٔR�\�>��>3)���3��#��4i�iwJ������qpڂ��X�G��Q���m����g>�CP�y�B�"ltK{����a�*O���nU���;q9�wkK�%u�Փ�A�@��a\.��wY�VS�Y���Y�ej�_T��;��w���>��� I$$?8!	&l�O�j��x������%�s���:1�ԫ�
�޴���.QX}����9_k���5X�v�4�Kz��e�tY����4��˓L�𺡬�g*���R��ʼ�^;ן	��V��Co��v驹�5�|JNPi��TC�TN`�~yFm[ƨ����38����q�\��I������	�Joqu.D���2������Y0>
��!�呍t��CB����io�,6�����5�հV�+iX<
���)��ut�H�ޗ
K1I�����+2,	l%B t����R��t�׆��lTw,��v+�@�ܻ����6��4���z��Ҙ̮�Q�'U%V��U��R����#�jeթ���ָEzhR��'�e�O�6J�C�{�9��<���3����C�0�Uwg�t�L0�&q�:���E|5���:Ț&	� ҳt?�����wı(�쵋��ǆ��f��Ł���X׫t!�I�{��u�u^����kUj 3����݇�A(��]���;�Â��f��UB�;X��&]s�0:M�Ϡv�,v�������1c�R��h�S]}l��9���8	ևuU뀗G�݇Q��W��fm�5��mN�Y͛�VqU����PYOc�Gh��<JO��
ݘ�[R� ћHX3Q�C����.�əD��)���,r(-���W[nWh�9�����ᗅC��*+�N�u����4����=G23����s��eoC/#@&�������6�=gc�GI�x7�R��y�V���e9���v)="�i:�*�����!�e���{��a��iB�)╦�fz�s�˱I���:ʏUF�QU&�����ƴ��`�FV�gT
���v��x�������ɯ�2	�W?�-����*��VI5�#�b�f]�}����3*ɻ�SY��ȋh��؄[ۛ�7��su���6���U�P�r�C�f�k����G�wv�m�{��or7c D��}\z���.�k���f��r��MwA7�	M�K��z�b��	Dp�9�c�i�:";9_)�ϥ�#���w5s5u;�`�%���X�z`�R
�vxȬذ�[ƺZ�cv�Xrm. ��)�����:�i᧝��2h�ؗQt�	��ۧA>�Odwg Ѱ�1�;��<gq�[�c��d�x��k�����.e�ݻ�]��n,��h��}x*ru=��14�{���ju�t�Ph
]���1wA�E�Ϻ�����Q���QҺ��-�js�;l$7iv�3I'1�O!7sh��R�=�w١�v.ۘ/�	�h(%8.����s<x�u�y����Z٤�s5uĵG�n�ӂN���Ktv�A��B�J�[碓\���3�Kq
GD.Y�BmIs>��+RkU�q2v��(YB�@��i�N�\�	��`�\B��0;�.��I.�l9jK�!J���Uwg�v
��ކy��*�;�%��d�.gؕ*� qT;��́�z�n�@-4l�ͭ�B9�t��p��f��͒�i��luu
͔ ȉᕕB\��|9�s�����ϐ�vӾa���g:�p��� ��WpzvkG���>�7��x�v�M*
��+j;V�i�3)�w�)cλ�-Vys�_0<��]l���Ck:��63
��s��/��sV�iպ�[�zid��g]6 (
D�ݪ��%V$����*�|�hR7h��z���	���ZD
ߏ2n&1,\��'-ʟCP�|��*y;���c�*�M.T@<�3YdP{�����zr���B���ۄޝG5f��1�D5}�\˚�< _t��;�i�%�9��TV��q�y�wE�*n����fٵN���ks_F�''qc�׽V;����=D�������0�F��,K��VN z�ZH�S��t ��ے+{Wڑ7z�����i��ؖP�v�_7������"@�W�/�:1�W]jy�o�o�m�)D��}J�w��:ݮ��tkEή�{C��ż;p��v �:0�����O3�p�1�7�D�Q�۵1�۠��
���k��8A��ʶ3�fB�Fs^.ʔ���Wr��n���]��)��U�G�֬ҋd�.N�� �s�q1�.�2�3�Jk�%�����A����������fu�(�f�*+��C#Z/+����ӹ."�U� u��r�9J��� �D�t3���<)̥�#Y4B)X���*5j�é�)�6��w�}�җX#ml��о�Vc��-87�գ ��nn�H>K\][O�	SozR�iy�hǐ���c0�!����;b�g
]Hr�B���V>72�e�����t�]�٭�STQ�� ��gVGՍR�����$1γk���V�:i�Z(U��r�+XG!�g�u̺=�67v�nQ�4��^s�l�¬r;j��Wԕ�s{��x%�j녔��;���Z�s����"�ۨ�j�u��d7BS#^sf¹��u�b}s���,�G��$�k����@��[,Ԩ�}��y]b��Lg���u���p�G�TTul+Np�B�7u���g�v�m':����~���/��sֈ`Ȼ^]�!�̫�[9CB��f_G yefk�K�Y�9=@v07��\²�뫼f�]җ#Y(��YSWgr��s�J���4ݪZ��Yf��VrI��9袱أ�	t��Y�^�k)�f��X8�Z��8+��civ ������n`����hp�:���m��~&�Sw@%��.[KhZa]�;a�^f+]����ޭ?+�CQȰ�x3�-�E(��h	#;�ncj.YA��<�ͥb��Eܧ�V�V�y�.� !-rI`���%�e�\���X��W3]V�M؝R�^�����	(�R�͉���&+@��S�x�'�*�ݼ���ӫ��ly�u8Q5�f
C�7@O8[X�7��A��C8�I�ٿ)!5(D����OF���z�W!�3��1݄c�@��Z%�S���қ6�D	x�f,�gP����Gt�|��ZE��޸xp�Y+�A٫7�Kv��p���	�ZӦ
�5�s@�I'�hB�&���h�;#��JެU������v�j&C�Ka��/Q돲��U�yo8ؖ��c������e��Fk:Q����i3d�m�ndj�`�/Xn�2�{6;�z��@�e0�����f]�L-6��ՙ�Һ���r���`�v��$�7yǸ7n��R�А��G�Vh�ɓ(˧zΪt�p�cH�q`y�vͱ���P�N7�>{V惹�:���������C,�lJL h��"�F�Vi����9�k޾�O��8�~̢�-Ӭ܂]��^��L��pjϣ���BWS ��{nw!%as����%_r5w��+_"�t5�}Î2�������s�`%�Փa�Q�-,�4��b#y�XG�6�pD��c���	�ǔs�}8&im)�ss���:� ��y]r��Ŕ:�mUƩ�9nɃ%�6�5nX77�w��g�k�շJS�3��m�'^v�UK-��U�Vd�&R�!rm�6nf�/!������BB��yA��Z��Xu�YX��f�T����6��(�%�)���Z����8����ux2����!�ڒ�V�&7����'�4s[#���)�ݰ&,-6* ���ΑM�WP:��-Vj���v�i�+�' 	Z��LW#44ғ;�>���t�H;�/�O�*Zt�fr�|�pБ8 ��}��J�����ș��%:㴕���ٔs~�N��U�(��ܐ�Lꐳ.�]�� �Tφ�[��,�.�^���NӴYgR����5��uJ�5��2����_,��Ս�et����s��7K����O{�V���`��)��μ� ��
��a.�֡�tu��+^��cx��$/L��̮�Z�v��h��6��}��'���GF���r�ů�6���i�8q���-�f��>�KM	�^�=M�Q�/;f�3����*�8M�u����Xj�ug,�N������]Mմ����u��X�d�u���<�i�������S{*��o&���Ι"��z��9��n��	Z�])z.��(��X�r������_ܳV�ާ� Ew�0����oR���Y��m�����`���c��)���Ⱥf��w���L�[\w1w]�Tȅit0�߻�Jt�.��9Άɗ����6���Η9çf��4�� � ���cl�:�ɱb����H�����R�r��F�k�8^��#+u�C���Rh��{��q �WX�ZB`�-��Xs�.�p���6V�i���sjAy��)h�*��0����X5|ť�E���xS��"f����d
�`"��.Y��SQ��Vu���Y\*i�kv-����x䭹�r�Ha��j�X�VN=d���<C���[Ժa��EB�dھ�x��b�Y���t�uw�X�L2��%sg���K\@{��1Y7z
P*qf�+�n�87������=V�]�s���T�.�nt��WJ��j��vB�"���J�����jq�u���aά�V�^�
��C�s��)J��RT���V����*�S��ݒ���h�*K���5�zN�P�.�hS�g���X�%O�s��B�d�;������YszXV�s	����T�g�\Y7nws�Ѵ�7	;�m�:J����=oZ���_`Id|[��wY�x���+v��>骶��f_^��yՉQ	u�����d��fU��񝡼6�D�ֱ��t��7m,<%�u�C�����1���ݣNwoѝ %��.�.��^�Y�V%�j�k�p�nC�L+A��Ĳ���oֆ(�g��w��/vm�]Z�4����3�b�r���ݠ�@�����`���g)�*��o8��"�L�X#`u�gח9��ô���ds6]5�/��o]��V�Y���1
j]�t���1]�mfB�����&�:Nh�Gm�m��̬��w��a�\fT��� g��U�k���Q�F�e�}6�����jA�V�a�X���W�G{ܲ�8.n�5��l�K���_��*+^�Gb��ȍ��Ro���{H�2۸��f&l�h���n.�.����K���˷��YZ����wZ����K_l�mLC�EQ�p��n^ 0�@���E&��`�Q��ײ�}�S�6�O�ִp�V7]��T�8E�1�زRtн�L��7$t��d�t����UY�}��z8`�jj�V�}�ݫ�[�\�ىQA�f7�֧]�ӏ:��WY�.��b�2g>]ytukc���Wlc�����̒6�$�+�&�u�����͖)h�L]��ncI��m:l��,N9�v
�ҟ�j��a�\'R#��&񊿤�tU�����3z�4�����qW]��v$(�4���pT5�Ep�����	�����+DN(*;�@��/o���z2s���&����Ct%mI���؉����Нݲ8�1d e	�4wrve��z�2�ɷ�:���0�:Yt�,-<^��W�v�׊�W+֚��D��Pn������4حseY=}+AԈWn:��ce0��ޚ��f�g�N��`:�ۢ^�\4��l��c陲�ɴ�r�l�k�v�-���v6¤���77��rY��F0��Y���]@��ܬ�Y��* 6�ЬΘ���	�٫Xc[9X�*̉�R�ʌ�}e�0������Lv�HC�:[�ʵ���<��]Jj��*��5H�`[*Ѧ�$�7b�F�dzo3/���5%+"q���m��K:+���X"��VL��2Fo7w�uΖ��`R��������<��
G��_X�[���f� )u,U��2ͺ��.p��m��>����ܖ�����Of�����|t��7��*���X�n��rs�Ħk3���2f���ũ�	�I���n���w
]
���ݢK���p=��ݗ@F^u�U�<���&��++�+s�n[Ȗ��./�s)po6pȇ;. �V�����Yض�^��_^8����q���n�V�4�}n'ܭE8��T�%��NM��t��|���U��u
ʜ*�����cv����L�N
}O*�k��D�������Gr�>قZ��4(�]����:#J;���r����H#˳qʗV��4��S8V�盀P��q�+(�n��J;�����qwG�Y��9oP[ն�A@�)��lw�N��4���4��Μ�r`]B������}�P�i��r���.�;G�]D;��j�\(��yۜ�i|��&,y;PW@4��M`�����Q� �{Բ,5��y��L	�j%�z��i|an9l!�ebP��ufv�U��qn�-�%j0�։}ܓ{z��69����3ǆ�:�h�i0���ɘ��T�6�i�۾Ok{ZY&ތs0pW��Iug<��5tU�=̿�p�x �����W��s��ғ�&�2$Wx1T���J|���e�u�,��ˀ��v�Q�Ѐ��{y�P{ā6����.��}npW����3T���)ǫ�������pb�W�e_M�@bPەcn�WE�;�x�PSn�h]+�%03�X�0���F�q�N2U��.w���lV����R�r��c�S�n���̮�zG�4���wc���$^gYV Vy�nءM��w8)�#�4���P��nŝY�����ol���z+EH���e�Fҁ&{�j���sݤ�kTy�;l����' ���h�^b��R��u�˭{�#{���1R�����sWC�Y���)faL�u2���% 1�(u���U�!�{1���j3�+㦂k���j�j㹸��o�_]�A������b���;	G2r�ȣ)G�Q��hX�)>�P�V5Ӭ뾻���g��u�n���!I,m��u+r���g!Zb����;��On�,r���=w��;��!F�jus�u�sC|6��Vv��C���4�4�0����B�����u��guKï�^S!n
�}XggVĶ.#�cN$�㋀�9�7�Wu�cgn9Q,��t$�og���*���,'m��k�.�%�r��su�&U�h���y���H�ٗ�]E��VD�[W���_^]&���u�}�Vw!�^˃iЍ�n#}�+~V���2��P�w��@'���ũ挭����]tT:�\ ��lX�c�;�*Ze�Xh�D5`ngE�H����^�ǫ�u��dT%�ugUλ�����r�fhT�dIc;;�|���ХG��Ttb���E�lhǝ�G�!���m	E_}�����T�yl#u�_"������H��*�CA�W��TWӺ�1u}*!���sM'4��Vzs�.�v�A ���ư�
��W�7���Z�����Լ��
�*�T��>t�ܬ�i�{�!GVJ�f�E���g�u�_#q|�w�R�N�LoX%�H]K����f�\���/sd��C]�c3�b�p	�Nj�4,�T.�k���"�ӥ�5j�Y6��%X+��쭀K��R�*ȱQVؕ�B��Ҋ�Nѐ"R2i.��cN��$��]?����f}�}�3������h�*(�ZF0QE������*�R(*�̵PPX)R��*Ub�$*JV��iTs1���UAkil�ڪ�U�AImX��Q�iTU�������PEFD`�T+*���V
��Z0X"(e�H��YQb��hT�)P�4��Jµ�Q����,SZ��(�B����TJ (�.�$S�"�چ�N(����(ȫ����mt�!�UȱE���IZ2
�

�Xc�"�J阊i�"���m+m�c
���"�a�F(���+V5�R�Z��Ȍ

��+*Ŭ��UeQbȢԢB�����D)Kh�R�RT�
$PXb-�
µ
�J�#��R�f��04�4����VAH����IY*�U�e�+
�ES���G2m�x��A��}��y;d����VM������dN����C�[=�)�<�IpHN볭��ֆ��a����ۋ2�[]�!T£fj ��M���f�fJ��E:�����k�'x�nS�n��<��qq�0�D����@�vk@?�3g�}��Kds�爺��|Ί��Hт��{��Y=�v��<Z�@4r%�`����1]9*���<-�Ks�+�VxaK��.n���6�^o<��oK������`3���u��ɣ��H\`YCY�±��p���e���Y�D8�:�ep����k��j�ޙ�0כ�z~��Q������5�S�v�����\V�[6�X6^9l�&
D
�ߛ�
��Xv{��>��5��%]����zJCoO�!g�t��/��\�y�3���"��P�gk��'{m)Ere����Z0>z+�y�Q���h�ӑE�WW�c�.
!�����Nɡ,4s�2?p���.��[�9�k9�8J�w�]֗��׷�M�V��\*�	�s1�n��E��aa�S=Ǫ�j�:�/M\�t8�����_RPsH�t�j�iGUf,�b�~�]�fq[����.��x�5v�,�i��h�xs�AܙRo.��k.���<�H:��7Y]O�Y�t,8ٺUαA��NxFڏ�,�i�ZyÑ�w�5�M���.|I�s��)�sμȲ�q( &N�GUt.����x'�s��J�ca�i�n_�*�}}9P�n(�F���[Bq2�[N%�ii������mMiB:)�-�����㡀/[���A�s�.-.�c������,Rd��"0հ�X9���v��4!_.�i}(Qn@`��̞�@�nyTd�HY/�Ik̻�H��5o
۪k&���|V�ÐJGw���۵
�T6B���I�U�v��K*��MeJ�� C����%I�,�fPx|bT�W�	!XJ3q�Oȇ~�>�g���8�Us��*n@�mX��� WL ����t�[$=���782�ʞk����q�6�� ��J��������)Cӌ`?u�#̖kE⎺�bK�͊@e=[{�T�{=R�ɨa18Xu�d��1�6�I�����ະC�Xu�^P�7ڔ�C�3q���ߞ�HW^L-5���f���Xczg�'5��ѫ0�U�����Oz���'��,u�2����j����)��
�G���x���[�^�4�F��&�V�}.R�
���<�o�5xa*�P�Yc�ĭv��={��M�ą�St nUN�Czz$�5:�zɔ����Z�4�lr��hx�<�Q@�h*�H��Fr�b��t�1�L�Fo�ܦWEw�Ý4������U�8h���9'kp\OB����7yF*���|>�7e܀���Y䈖g�������j�DE��\U��@�ܖ�q�;{W��(Z=X��V�V|�h�����7��vz}ig�{6�7Vf��IouV�aƟ�kV���I��`X�5⿭�Q�h�H�ʲ�Ȋ� =m�k�rMM!��J́p{3�o�|VGL������h�9���LZyE��A�N0g.��-d�ݮֽ�Zn\UXS�@�a��C�ʲ��ņ�K���7��!@�z[{��k�s�pXj�պ���j�����iw0M[����r��5���w��֓sX���<��[�p8�!���vK.Ӯe�����\�/r6�#Q}��;<�GX8�C�x���U�=�u��;��iz����}�n���Gq����M �/i��B���Ł/��i^����s
�u�6�h�]+�i;r@p!��B�$V�D�p��m&�mK�U�8pv�1\���72��/�˓U�^��.r~D@��@��FM?dfH1��f�"z�t�u�yh��Hz�.�CϞ���D�.��WY<��F���<�e�z,�R�,ƴ,�v+���r"�3�=�ַo�')�g�>���鹻���A����O:i	5�C���W��c�\�8S�]O�/)w�㥓�1#>�,n�	C8ĈA-ul�����Z�O�������rba���UZD���eh."���urw��d�aB��+�ޱHp"o��k�ŷ}U��E�Cx���8'�aR�n���ٻP�3i�� �L&R��.�BW��l��*.Q���81~
	u/�f��˨٦�j��g�D1Y��è�Z��_�+]BQ��[�	�B�鶕Q��'5Ȁә��O��Q�mI&0?�@�m[�r���|���D�foq��^3<3�q��JmTD�t���r&�yr�T<������{.�D�ΎJ��Yd�bw�7��(��؜:%�^��WR�gZ R�O�:83a���Q�Z���c|���{���>�j���Y�E
��F�e�W2��v��c����d��n��M�v^�s�3�I΂����Sq&�)�����N��d�F�C��޷���x����Q5J��{���'xj.Z0z��g1W�w��r|j�f�UO�S�]�i�#�g�]���T+�\֍�>�D<�!3����[�
���E�=�0�Q���D��n�uF���N�_(���m�m��჋t{t�ܭ���L}�f�!�6��q���a��8����ي�Q/��]ZbBi�T��\ ˽�J�
�lt�v)Z�Ց�c��j0�i_iB�Lɔy�!
r���T��T��.;��:��l0����=~ѣ�I�F1��3���9B:�E��wh�ց�2ii��\�����-�HfN��#�p���TE�|��g�D'��Nk����D�)D�c�J�p�����O7x�}�7����S&(hVs�W�>���2!|��[w�#�tƨ���\���=[��]��K���@���:�VѸ�n��#>�f����Z�to�0��ۼ�G�hn
 �k,S��<7!_p�h�~V���>fUh�zWl~A�&�l&��R<E����E�� L't��7LF����o��T���x��������&��9��ϵ�=QS�۪��[��uw�p�A��MͲ�{"K�OGw��V�q+իC��x��
��νo������d¦m�]�C=V"��;)4�{�Po�]Ѿ���9�#�h��e?t�"Gs�`cU��5��F�;�G=��!Gu��(�'�y~6�%{`�+��$�n�aA�y ��gudv-.v��.'�"�{}7�[c���V.�<���99(Κ�Fv�X+���.���M��/6VV�Ms���4���T��� r�6w��*���Xx]��fs��|-t�hGmn�d���B�z��6������T6+���`��hxT�@m��]N F��9�r��BnSf�Z���zz�Q�����p5C.,S��E���`��t����S-�u�i�k�	�t����X�w��J��Z\>�h��_��g�Ƽ֩�|WPO=άV��S+�C��ģ7��.� ��|���I@8S��p1\��~Uj�-�ͅ(���B�&Xz���6W�!��pܾ%S��a�#n�Vz�ƹ�m�g_A�[�4N�2jc�Ny�YHDӜ�������r0���<�.�tM���\�7!!��W$�P�����L��O:Cpuѕ��4 ��qL��ۇ�VY��z�� vv��� ��1�A����롈�B�6%�	G|�f��v�~b{v�@4�>�նs��܌�E쭾11�:!��0�tB!�;�8h����3�Q��3o��3KY�N�]�S�ʭz�����>�b�.s���K����5n�1� .8jP��rB}g
!��S��D:xl9�y�J;���,"�AOs&�zn�o��Vn����S|�j ��xN{���JRu͌&=;���x�+�bYV�������*J�����1cܩB�m� I�; d9���rZ�1��ks/��55�����o(a�P���%m�P����>��U��[6���=��7?>7ʲϙ��˒����β��	��w{���Q۾@��A��*��P�4"�y�VJHs�+�jbð��"���U��F���>�5�v����Ԇ�f�g>�X
?xJ[��%��9�%OU�o*��������a�!��Wխ
(�L��څ�����PA�6����s�������n.]�W��	�q�܁���i�"6̥k��y+e�2��U<|<.љ=�`>��Z��հ9�;�γ������m�3b4kYDn��u84\�2��V�'nm����.n^+ژK�cp��?u�j�)L���j����<"�wu��񭥪d�;�bU���ܻ&�i���8Oqj:dJ�l�pڦ��t8��2��#�X��1R���:PU��ы��f����ۘB���9�گzX�=��.�:օ7���/8p�u�\~���}AV����,�Ԫ��������R������[�G\6�(Y��WI��ٺtr�f�bP��q$��EX����7D$�F��,�`"��^
�PU��e88M�x��3w7^*:�TՄ��ڱ�V�\�+��!�V>�)�Ӷ��'>zDU�Xsu`���.�{�x��۔9�#�-E��i1˵8��et�l��yD]lݝ��B�V�Th�����M"�	K% #	����2�j7J������SJ�u���;,R��dh���pU�������		�����D�����v��tf[]�-����ɕ��xW��h���tc�"�ʓ�����OY�D*zJ/�\���V8W�e+V��৻^�§1p�)�3��A�����Y}��]�*q[�t���=侴׉�O���xfQ�x�>����6}�{��5 ��ک��C{xc���wU�*��懠ϛ{�U�ϭ��|��P�'���U����^k=�������R���X�⪆I� h�1p=���W�&��<�ϩ�WC>����Ίyvy�C���9���ق@Єhnf��(ٿ����VvL1���ó���U/
�{[����{�,����O�-\<���dg��/�~ߓ��=h
6���Z�[Fa݇��ɋ|��/ӷj1�������<�"{�۝~�둸��o�H��dGU)����S��ɺW�����w�UPn�AoP���I��}��a(�ԝr�Rh�I�݊X��O�TE�n�~�+���h���\�c�X��9ڒ��[���R���Z��s�a��� ���\�b�tC��0+�ԫ�*����sW��[$<��ր����
���Qʤ{rD�٥����	��&=U�y.��+RU�]gC�_��>�6d!���ӑ��!�ѥV�b�����p��)eW�;�N�k��"� ����$o��c�����Q|T����hΤ��G,��u(�c�a�����Bƀ\����3`3T��j��1s���-)8�f��hyw]1�r�.cp���_Nؼ���+I�Þ��UH�%����W!�Nd� �ل�W�e�(`T���4��,(��w��rP
�a]��F�#)q7�t!8���+�Ð\�q�?VW�Q0���O+\�5hDkP�S��r���oy`�z�q4,����f���2�y�t�8�)�q��u�+�%Z^.����.quVŝ*,�����;q2���-��S�J�uӞ�I���;Z�id�m�X䶯RE�r�u�,��Xt�@B�e�������y�/�=��\���^���(�x�.�VF����5���Ym)�^Pwh��I�}��>��*a�ֆR@eu�B�T��ifʹs���{s�ԩ6�A�X�n�Î<�.��#�/f�FT�� �IG���%�V��;�]�mn��.W�wq��&��}V������tFm�b���-��8͸{�F�߾k.�T'�'CRF�\��T@-K'�`�z��m֚ӿK�n�cH��'��%[�w��V�y,i��,>U_f���Wͨ��7U��3�"���/�I�����;{���8U���)���fǐ�9��z�WN=�M�:ch\R����S͢i;�hp�Q7Q¢�҅�����:��@q�D���jc\�W����E��tr�'3�X��膡;�=�k�����V�+g�/ΫxDު Ԟ+���QV�rXx��X-�Y4���U�=2��K(���i鐆nU}1F-��*�y����i�}�IV��m�.#0����M7(h}bxr��A��P���݌i\���6������[y7��/\�)��
�ܦPϝ�h��Zc/�j�#��F�U(Co�]v�"�͝'���/���A{�l�d�:�����3�!g�������e��њ��{v�.�k��0��OPۦ��5^ =;��k
T��S���}9�z�z���W���1��Ms�7b0u��Y"6��כW.�YzE�h�,0��w�r���&��7k4�1-���X��ӽ.+����-,�b�&��:���w�f�N�U�S/T�L��4�{i�N��ds���9�1�k$�a�f]{�k����){s��j�|{�4:��N�m�W�E����R}P��O&�ބ��&�r��1&�p��fvV�C �7(՝�DP�m��i��ņ�v��ӱ�۪��*n�X��o@2uл�wu�v��1-�]5ՙ�mΙG]Y�)���.���j�L���̊����;M%���e�x����5ɲ���Acz3��m�j���jf�*�@ ����y��e��-��FE�9	A���hĦ�9@�γ�6`���uҩ1�Ryݏ����-��N�V��v�tgwM�f��_i�2�5���52���׻6�{��s΁����a�Hh3�I�㊇�*º����[�5��w�x����op�3mq�(�����L_yx{�� j�MOMi��ur���&U���C�r�:Mf�Df]�%�c)����<d��Vj�����v�HiÝq�^kh�f�q��˫���M'�w ��oy4y��U�����U��;\j���j�ɝ��|�N��(��r6�A܈u��	����r�,�	�z��6p�ĳ����S3�)J�'�_E2V�y�5C$���<�;�X]�QYd�iר3��W_b���K}T̷T�ūf���g!�Ǆ�D;���uDn��˕�t^�㭳uܣ ]s�\X:��kp���q!h�d	��/4Aՠ��#��� ֫ �OA���-�(R�=��zU�3Nc�F��)�o�s�ƖV�IF�#��
d�r,웓w]=58�#zMbVk3�q��}]R�d�j�*�Q��h�\�K����}��dY��wbt)�I�����pGt{v,�l��U�Ӻ|�;��R�;U�fV �ӹ��J�	���xFZ���B��˕��x�@讦U�7u��b�.�c[i5ٍV�<�R�#�h
@`��k�.`n��vn1�Tq",�o[_�;;͉~>��7���i@Bڇl��+��u�2�f�������Vi�O9�$þv�=�ݲ���:�Ê�
��M=���V�΅Ng������4���ՠ��Ϻ�U'�����t�o��u��
Fo.�*9��N�������f`�|�Y��SyǢ@�Yuhh��������Ȉ��#͋��痽Vw^�ڽ��mA����nl�V��E8��P�h�Bu[qYO���'{�n�V��k3�
�/��X͢��3 �ӂF�N��ֳ�q��(Q�P R�� r;�8���M��U]�7�nT+�9Ѽ'��aQ��ICC3���Ş#�k+���,�v6�f�)޻��̚�|�Φ�G��pT��$�ԩʙ}tNL�U��ܹ�j&�9\�JU���%�}WV����]�gy>��N`dn`��{h��J������ة���S�{h�Lʌ�(*�X)��������GI�"5�#Q"��"����,"���Ljb�-Qd4�YmM0*
����ńm�%t��
�PZ°�`*�V#J��f���nZ�b���̴�*�()"�WL*��aU ��G-QdkV"��
�����h�#���*�PP�+""�k
��IR��QH,
�����
ɤ�T+R-I.YP�UR,���X���%tʊUH�ʂ��TU�H,�H��HJŁ��TR)�Y�E2�J� X�[H��P4�Qb0U�Y+!�F�bA`�eb�b�Ȉ�H�XR�,�(�d�1PX�X�MZe�`�*����Aa12�) ��,A`��z�n@����{�b[��;F�Z�2��*����9޲�`���l�b�ՕtSط�z�>:�7�:A�<����'Y瞝�]�gI���g�k�IY������Q'Y�*�j�I��%`|��S�q�����C�8�]��A���=:�Vx��|�������H�Z�R����W�l�	���b��3"��+;d�=޾`m�d���7�qǤ�ϑ��*�yh�|a�t�vn��4�Y_P�i��bO2�3�>f!��� >���z`�C<�$W���~W�~듴�Rt9���>x�:9��6��*c�N��� ��J�ιր�LB��٭B�j��+=�C�c���LH=Y��x«a���V����F��j{�-����\�W�z�L<q'��c�<�gx�9�CIXq;LI�+������t�<哴�%eg��3�i�g<ɥf$�+5>�(T��=d�i��4��@+���=f�W��;��!��VNKb�2t�u��<a����&!ĕ���&�1 ����7�'LĂ�s��I��c:5�I���q:9�h6�R�9�Y�q�C� ����x\��-ǲ�^�R�ݰ} �T�95N��A{C���ͫ;IP>M�k�+�i�r�:Iyj��|�xɼ����!�K��ڛa^=$u9�I���Rj���*���!W(~�R��<=�&o��w���F�x�d�0+�wﺘ�M���&!٪Lg�|�C��5CIRz���'HbA~z�i��Ɉl�ɤ�!S!�V)�_}�x�Rq
��>ɶs�!_0�\��ּ7���>���>C�9>��l� ���%fՀ�{�����Lza�7��1��$�:5�H,�'n=wa�4�U���I:B���~a�1!�lDBG���/�ݧ4 ����y���AC�[槬�Y�J���6��WI�&t���L@�*l����g���_XbVOVM�I�W�OS�w�4��+�v�^Si����r��}T�o�^�Oj��^���O�`_3�/�X��$�����w����:@�Y7�a�Y�8�'��󙴂�z§=��m �CÚ�P��VM��;M��+�xɝ�z!�;I|�:Փ|�gi@����|��}���==T{��s��7@�F����7`\��͆iD���ѬoL��f�]�MWY|RP�mŔc�x&T����^��R�)�v4��n*}`݌ko�:0qYu��5�{[Y��p͍h�ܮ�Hԓy�-Z����i�4�T��z�V�+5�9��01P�3(>�H/'��&��Ugl� �a���h�;a�
�Gf��&'�=L|/_j3�=f!��<�6�Y;��C�1�ϳ���>A�D���&s�Y+ދ�o}|OP6���$���=I>C[�ĝ}Bl:���� VI���>d�$���P���v���$>a�&�XxϾ�w���e��)���|D} .?E1'�T9��/L��3��tn͠t���A�d��LH)�3�%a���I��8ó�p��$����1��gl���ɉ�O\I��;�k��D���;z}}�|�A>��	�\k1�T:I^���M�H,���4ɦT���II��tj��ja�z���
��Xq�=gϬ��f� }}�c�#DE�� c�ѵ�̾SCҝ��X;�T��G >b>#�����"�C���9M�;I~��CI>B��{ޤ޾���ܹ�������5���%J�Uٖ$l�S��1��+�7:��zÉ�8������5�:�Z��ts�{�yΒ<C�bw�
������1���l*<~I�w� ��v�M�ε�'I�N���m1��6^��a_��1�e�LC�>#�g�~���>����r�E��[��n>��y���z�w퓶cT��|�|�w�����C}S��6�Y�f��ĜB�6}���Rz�N��Md�1���z�H��a����>t�G�_|�"����:�;9eX�^O�~����]k��E$��|�����1& hߘiN5��V�*xɷݲ)=B�a��q:}`Vq'5t�ɾSI��5��L�Ɍ�:������}�>�$DEB�94�Ϲ�񚚭���N��ht�C*T��+�xϐ������Aa�jn�}I�bA��iY����a�i$���v[$:C^k��I���q�[�`c=3��}c�>�(G�G?zk����ax;�3��Y�%J����ҐR��ޡ�bt���w��6��z����W��Ag�x��Cĕ ����4�i�1�L+�
��C�yM�|�'h]��F>��} }��|'lus&&����y��2�i`����a�3R6�&��(ۛ�����Q��|z'�K}t�+���V%�o�No����[)��o�=M_uK�_F�6���\9$InX�dY���'KڹI�syn'���
��'>���V�N�kz6���L{���Y*��	��z�V3�I�/�O�.��0����m ���<v��VM���� ��DG��}N���k����t�����18���t��V����x�& t_0��eVx���6��v�x���z�M��J��QLE�ֳ��4�S�N�{5�I��!�0}DCe���c4'��s����ߔ����q��d�bo�+�=�o�Ax����i���
��}�v�3�1:�w�1 �9ε�!���=�Ya�b��K��� ��#�4A첽g�jzD��coݔ��&$=N}C]��Rq���2]���ӌ��:C�{I����a�;�GJ�Ug��0�8�a�
��(C�>La��;��:H,��z�"$G�G��A���y^��~�s��׏6����x�3���j�Tv��j�@�T�&��i6�ɉ���4�+6wg�i�a^���!�*C��nߘ���}�@�,�3�}鏨G�"����lg�R*;����Į��z�������{���&'
u;��&8��+Ú�iY:J�ǭY����͍��R�}SL4��$��c'U�!��I�*O��7+������{a�L�qގ�y����]�<E�L��'9����2l繵`);B�s����~�	��k�i���%gL��&&�.�
�4�o����yC������1C�>C�����qhp�_f.�g��]w�^ t�U9zÌ1>C�1'G����0�g�w�a�%Cԕ�}��z��AC�~�ASj�Ry����.��e�$��>|t�풥MM�iR
�룇���s޻�g=�w���&ߘz���vØ]0*C���,�<M�|��O��>IP>��U'P�;C<9�ӌ*5�nN�>J���I�����w����_X�"�S�xDX��|~��Kb�Suf��]�Ϸ�[���b$�|�S�������� �a�W�
��/�<2ϙ^���}�zI�|��{9��I�!S�@U�iXvs��H/̏7�����Y�:Ǯ��<7z����l̊����.&!<�����h�o���ac;�4w'�
�ù(��_h���	r��X�\��+���#����ht�
V;��{�:��@f�le�ܺ3N��kU���)ݭ+xg�����W�c��n��3�<�����}�䕝3OI1��&2|ʬ�75CI4�I�bc�|ɞ��&>e���,�k:z��i�����w=Ü�����Sd�~���Ưe�����9�{�Ud6�d}/���" pKj�����w�QX���L{�T��8�L��aܾ���,�"�Ȉ�r{V_��]OJ�k�0ׅܪ
�P�KL�Y�`ɼ�֨�1�g~'CQ����9��8f¾�ny��5��ޣO Z���W�{��N��sLX��DèIٳ6��D��"�
��t~G]я°O�,�`v�����#L�k9���??'\&��cL�F�G+���׍E����6�d4`��nW}qU��u7�j��m�pvX�1�u�V8S�,;|�6z���|ê~ũ���zo\�?h�}�����ܱA½�p%a��"8aɆ2�҅�0N�R�:e.;��z�������[ ��	��DS����+��=���¯�����ط]f����<����\�d��ӏ^�͐0h�9M��]p�p���[8s�X��i���O�5~!(������hl��kI��;���V�g8�6��p�I��!j��<�6�gI��GPv`X��%�}[�rj۹ 솣��ݗάM��b�u��%;;�F����[ʃ�����|{4?�w���՛ڱ��,�5vg[�|o�w�X{ݴVe$�č��eC45L��f�u�#Pܡ���Q㝸���L����^:#�9C&[�8�`u�8ٝ?U�|��T�Ve3�]���tſ�������{/�e�����fbүDh	7�?�_/&x;�U��l�pf��9�5)+���7�dSn�^����Y��B5��+���ͪn�f�)��w�c�K��c������n��o�{�Y�(�s:��%��y��;.��4O@YuR)J%�!R��WIGi�])Wf�m��)�����x/bS�7;<���%/�4X�lT7L�,��Q��\�9�+�R;�[�b�3oL���$9`�XvШ�0ٯ��`=��"��t@F#9�e���t�:3�Q�k�[G��q\y��wN|J�\����=L_��qrr%���QꠁQ� .;�"\��v����6!9"F���bu�p3OP0�����O���\�O�cȘ��2��ź:�{������MV��:۵P{"��4��ic+z��,)b�T�v�9�xn���Q y������u�M��u��"Z(ks��� ���J<���Y�E�8ݲ�c�YΣ����|	Z�^�\�Һ�f��J����4�jV�+�]���+�	�8�)��Z7�(u�����__7O$�B�_Sw�l�sH^suuY�xzB� v������]���^r�S�W1)��!d%�+��eV ���?����$<����2y��'�u�~��jŎ�P���O�Bo��w��Rŀ)�X7���hXxHP������4��Dm�T�p�V�V�g2���Y�R����TK�X�kiO��8�3��}�;ډgDh�MQӣ!М�/�|�����\�2�����a�'\�F�b����b�Req�c4����z-Qgϰ��^���-3A�}�z���V�v[|1�j���%|g֓�䪇^�6~�Ζ�d\���U�٤����F�Y0����z���`!���JSpMg�	UiWQ.�}g�:�,V��a��pĽ�����^���5��g��h�`�ʲw�|���_J�-�"��������۶���p1��3�Lv�:CE]<�@Q<_30���0G�e#���{���q|��rۉ�Oh�Dپ{P٫�t���Dr7�pW��Z^THW��!#p`�;�k�������c7�_�,ٸfYcI͗�a�gp��)���9��7=��=��E)=^���p�k�Ə��1�/ָ�g&��Ͼ�f=�S�͆��>>aN��Ȼ+�i��v�v�{��ع�ub*��&���VpW�t�\7h�vs���)(Y����ro�\�����|j����/���c#foJϝ�Iݺ,]�+r��{��o]�����a�����&Y�,tAS�b�&g亸<�T��`8Q鸄�!U��De�w����R$ �sbb~ɩd��Kj$V)cw"4�pa�a��g^��\����-�p���p떎�`����V����-W\VO���C���Oz��`b�#ѩp�~|T���b1B�T�fE���	��Q�5,v�M�n�+ͧ'�ȵoe��6+��E��.a#W�w�2Y��B����\�;�ba���L1Я\��T��M(}'�ʩ���:833�boS�y�k��3�ʟ�����$Ō5�E�T��ud�('7LeŮ΢��ʫ�3�Ui�T�*��~�O�y��Č��Z1��;02pt�m��5�H�>�yW��W�vxJ�*a���cC�>�� u]q�I���݊����B�j�c��(����5V6RU�]g�&�g��H���i� �~��^��^'�u�0ÓѧW�I�	34���M�l��N�Ј�D�/)N���7:�f��4G�pӃ�
�Ռ�qQ{=�"�I�TD�W�T΀������W��ۓ9ꩧ-��ga1�����ӗ�ήz�v�7����T�Lf:#ע��X����L�9�]mW�����;�{¸r��	��k�1Z��9�+~5}�PS�ğn��Vj�S#t��U�|5�۔�vS�8Z���Y���D>����� ��-}L�<�7&�<��ъW ��}�jr���h�;M�ܱ�J��3�٤{>��DP;N�r�9SZ����tgi�U#*] ,�h�aC�:X��S��d8�zp}c"U`l�ξ��r�q��J�<�)���ʉ�O3�B0�(��:����B�|x'��M������􆴵<>��IJ&����<�ER� htr	\c/�Q�ZJ��j�b�*r��8IeV�l�@��w(�<b*����@{�>Ֆ@�	ox^�VSX0�jTt�:U��`���:ПU�K{⅀:�� �Zv@�2�3�nHr�d�UR�i����.�/�+K�ō�0�'�>Tf�#;d	N��MdD�1o@t��0����*�1�8'+�g�͕���(:�b���S����k�sx=~6�*,|��9�;���P���f��R���K[th(Opت֪:8U��ޓ��dӬu���n�6qR�j=�����x��v�a����hl��@R*ع���'e��>��p;F���$�=b��ֻ)+��:����إ�y��8Y�;1$L��eqH�$���졣��8��:���n߮�/������6�7溉y�W�u�X����A=}}�3�{��1ҷ\��
�a��^^.j���X�oX��4J��"җ~��siy�}�.Ǻ��:�������j��=��n���q[O/]=K���;)sl�s�)��2#pOғvx���=7�<9�o'�t���8�ͺ������uѺ\F���!���&��0�n:�4�r��}�x�-�(���p`=�-�������ZӃ�Pu\;�&t�Qg�#j�
��j�+��0�w�Πx������t�nn�.����y��F�l	��dT\�(a<Dj����d3�n����yy8�jr�o�9٫����X���3��;m�����|y�4"i�,���9�;��,�x�(�zr�[�v�eq#k�v��<}B�.5��:�6��]ω�f�z��
=4=��"f�\�ǋ�bE��q�Ġ��c�0Pt�Cr�B�%��G,����N��ٲ��S��V�͔౑r㪁y�.�8��yo'����mM��5��4��kj���>X�[ Y����^�T�PX&j��Ջ-�j�_A��fӳ�#]�i��NZt��M��;�L��Hw���iE��}ӳv�n��H��������O
�������q�M��!��,������v&Cv���P��苅!�*����b���fĽ��B����V�H{�VMW�穋.s��]����`�6��WK���<{�w���PQN&�U�"�?gإ��a��P0�j��`���R�1�m��8cj�]����- �Ux��&&�E�Q׮[���1C�����k��9*N_��^��Vu4��Vg%��~��
�) '�ϼ׸��(���Evk�Z�ay�F�x)�إ5{.K��o�8pq����ꄎϼ��g�?�{B:d�gNE��̿c�~+���w��J#�fi����-���@�r��	UC��:{��&ED7 `��t�9�;�JaF�w�c�5p��[�TS�uZoLF3ZT��Vf�ӟ7p���)�ƍk(��!`��Z��2�d�%q��m�}~����5�g\�둦4�b�uZ�%2���i�C�����񆲱>����0G��W[�>�`��~f��u�2������#k�����h�� �|b�X�]B;h�7�e^����,l�g;����0��t��txؠ-�t��;�;e��jv,͜6����IID[y����q�Waf�������G��ĬҮ����T��X�Qf�*J�ǽ���U%z�����M�ܷ]-�|p���;1=}��c8'n�#-�Zμ�ӕ:k<�e\�q�����{AmPN�h�j��,�*.e�V�(|�����7����f��udj�r����z�X�f�f�m<����U���A+W!uy
���F :�r�R"��s��N��췘��Ѩ�G���X]��W4�CV�
b�n=�+X�U���
@�u�)]�:;�v�	d�vFq˫�d�yN�M��`u_�eAW�D٫z�EL��2��)Z;U�n'�6_46uJ]8��I�8����*8��߀�*�v�uH4S!8�ٜ%^�h�Jeh�F��´Z�2�lK�=H��sU��Ө�+���`���_-9I)2g�cx��Z薳��,�[w�i��]��33��������{�(��sS9V���2@�auǒ��2����=�ů��%-QM�x�	�
��J��(��j[>;�7	���vj��ͤ���Dz�Y<�s]�B�]�\6�ecG1����P-݋��"��gTŁ0��Nk�;,ξ�t�tמ�u\56�ﲐq�e�{pѴs��}ru�
^t���vpv��y�BH���\�:wu����U���"�i�j��pQH�q����#S��D���[��\֬�ꛝus���=�r��n�c0L�F[��Qc�(���5�,Z6�B�u:����@��SY}|^�6z�6��|W`�Y�x`Q.��t���:-vb�-=������a7�[&3ǅ4��w�I���TA��MN�⻩g,=�3kH*���u]��R�E���|uX���T��):�hp�4p�Isc4��Ҝ�UZ�U�1���E�x�d
�x9�����6��a����۩���L+0���KZ�:kr��	xl�Tt�\]k}|X�W��Dt���UѲ ����d҉{D`�;������a<���n�η�{����Ae��-]mE��Ƣ��������U':�S�#_��h(f�-nL�J�[�[ ��oWQ�<��n].�v���a���e� �ʶ
�5_m�i��zӹ#.�ٱWR.=�˖�y��5����f���� v������I�`_6"2��bhvMPn�_*U%��<RN�}�r�,7�/5k�	9V%�84�9B��S6�`��r��@6��f�	WT�J��]�N�/VlM��:��j�wr�-h�]��pq�G�*�|���j8,��kr�6�^,}n֨
�.���F�>��-��h�v���W�N�Ck��GwDEm����wZ�n��e ڎ�_iTi�/o�m�nPV.���`g��Uk�>�3t4��Xi���4�Ŋ��AGIdX��R,H�jU`,]%ABVDaD1���U]S�
��AE5s"5Y++X
:�ST�(��1PPU�*�((��*���Yd�*�3J�"��eTP-�Z� �QD�LJȡ�q�D2�@Eb�b�������b�(T���dX%H#b�PY ������XVQ&!0H�DF#X��Qe��,Y`�T�ARDTQU��Z�R,�ȫ2�b�AJ�"�`��e@���Kj �(�R
EX�\jȨ�"��I�3�FAAQH��*��(�P�*���#X(�U,Kj�� �Ld(�(�D�B,��}��]b���Kb��K,���w�չՍ.�u�wrr�G�[{�o&ؗG�q}՝:	�n��ܹ�5s��W�}v*^�\�g��K(���[8S��&5�<%�\D�o��Y�&co�;�*�27���ɽ�M�(:��&����e��Wa��=���y�.��*�����^����G���끪����n�CB�]�1Qk<zC�?%�q��?G4����G­�o+�8�8{J�P������"��!3q���OK^THV2H�C�%���-�L���k��)���nʒC���b�1���5}�
�Η�3!�iX%a���ȗ����L�fl	�ެb6,ѭ�GG�|��|���<�XЃ���d6z\�B3��/��\��A�>U�)��au���P��h8��K�&'�ɋ��+�;�
]0�0ƙ
���.�L���������Ѩ�z}I���o�t�]y��'�O�ѱ¼�m�e�q9ٻ��0{���F1�"�CRh���t` �n*Q���q���M�u�'�T�I�^U�;4�r��a�g&;�t��*���072�؀�����~��zw�4~����^l�[��|�ߔ�Pܸ�������%�����T���[�ՒKM�Ve۩���`��e���}�r{����)��&�U��I����E��)s��vx�X���R�q�q�;\#Ķ�v���w��+(�]���}��g78�7�k���ٽ)�&��ާp�mU� l2�G���Q��e�mH"����d�WD����Z%����QXve��4�
�IU_wK�<�Uȱ���N��ff>c*^��M�{Ȍ�x�Ss�\"����/ʘu|���cC�*�po��G{n�{��}M`�������!��TQ�����#PV�J�Mj<.�W�~ W>ycLus�Vk���֧�YT0[�uZӭ�p���<��>�<7�u
SPG����=�}�6k��T��%c.8^L��s�ʧ�R�S1��1�J�z����M 9N�nUuTI;N.�N�|��G�
`z9TD���d���յ
9J��D1�m�b*
�lgN�G��������i��(d����T���`U��^:����N�1���_ѧ�s:�_>4j{m>�g]��x�;�c�pz@�$�'��=�S]�J_E�|�W���I1᲎�Z�g9�ջ�g��@깦b)�d¸�1-�ͪTb�'C���\���
�x��_L��S�.x�i{GL� [�`�e���o�e��xh9��N7� �� ���wm���V�eM�+�5�f��ip�Z�
��0��g�2��nָ(ʻ����B��#`i�W�MV� F�'X��ewI+���1���4��k����U\B��t���LE���+>u�*����̣T�|��m����'��X��6�,�9wr�Y���Wѣ-�����5��g>/i�!
 v��Q�܁pd!���w�ZQ]������H/��Ńj�m��R��k�y�����mu�)� �J'Er�2���k���튬�1q}����;^R�=���禧�Sn*t�5U����Z+dr�+�j���t�$D��`�2Z��qp�j���Z�A��o[�c#�
�����q6��m2���ǜ����{��[�
4V�6����< ����^_Ջ��K�T�/v��=7:����gOm��t�U�/�*�X�=���çg�pGW���r�j�8�fۢ��q��H�@�ⅳ������P����塆���&*�lk�����Fj+y����3N��C���p|�ۆ��er����D!3@;��-��=9fo��o&�k9>�|�P�?lY��n#T�W�ܦtc��'L\��ѱ�@:	�uN:f��w50+[ٶ�=Ą�oY�i	H�93R�sc�ڷ�R��a����-�t�\���mai�$�hg���S�{��J�����zR_��&'�}r�������"#�VZ�.����3��6��u���f�<,d�	u�L����9��'ޫ<.�9��d?���e% Mf�Qr��q3��j���
fŵ%��g�;r�	&6�,�S.��X(�����e6)ٸ��@.��2���S]���}���!��Hv��:]<	�;�V�+�� ��;y«5��U!���v0��ʷ1
�l�Ն���K2;^��r�"�U� �_*�);g!d��k讚`���9�e'C<*<��,$��<��8<�O~B�f��l�9��{�8EE��*!
H�j�(7��y���.�d�h�	�C����|
�@Vw�M_�R�c�����@o��#hcȧ
�neّk�\;�j`ӎn�EE�"~v�1Kӹ ���U	S�1��ϏP�fFmX�
��'�W7@T%���r&�hȣ��n�s��c�����y���DKT�d7jz_p���:a��a�ϋ���� ���얎���.s,0��8������[&@�o�=�כZ0z�(0NuE9�N�2ҬW���7:��o� iy������ʧ��a�0nГ����um%(��@�"�����b��YtFt�T]����E<05U�h :f��r��L�
u��e`)�P:'6H�9�6�\3,�����E�����M���`X�jz�`<��%|/�z�k���O�,
���G�%(g����l�F����ٸٮ D��S0�Q���q^�>�,'Z8iג#l�u=&�K��2zӱ��)��ӕ	���l��T����VX�t�_h{[QI��+/[\�k�|/�<4��±�#�EXU�ι��R4�Di��E�X��R�Zr�Ǝ����z#(um����7z}�ie��5eS1�&��������D\�#q�/�Ȏ�Q���7�fa���ͱ�^lo��X�?Q�����̤}�D?J�\�yJn �x��J�8���-A�l�(d/f.���6<,v��/���p6��tiM����?\)P
��������N�_B�Kp�ꯘ�׵
�j��kD�ۚ�.����R��`%4�P�y�z�ꜮIs���/����t<��ڄ�E���9H�$F�q���yJ����B�����p����P�#�g��˸:
UW]s�J�^��f�]i}�X+��!�����J�o��%Tq�*�:�l~��`K�ʕp0t�oIT�W���a���ʒ����+s�jwwmY�8l�Z�˶M[W=�y{Bl7ܔ)�m��`�����]�wj
�^� E��`l�����+{v�:�}"���k7}�9v	=Vq��S�9P}����=Y������kCJ���Fg;�Θ+���V�+&��K�$�����V��s��3Ǘ���:�9?"�X]�o�K�g����:A�|�3/�[���;�����t�#C������k�z}J�?��o�v�u�-�?/���xrХ�uEa�V��g� 9�p�/�0Tk�L\f(T6��̋g��w����G�����~a��:��5f���ģ�S�ڍ����������k�Tγq�h�2ð�����L1��U�4s+���tv������zV��kgC�����N��ڦ��s<c.g��66������=Q:6�.7��V�,��V�+�V�|�yM<���*3���@�___v;#Ϫ��<�0�Z��<�:�f�?�����SMp{Q;<%�S�}1�쾈���MU�����py�J]ߢ;�^�K�܌��̎5*͓�|�A[��u���x8����?cFK�*�llQ�Y�Պ1ڪn�Oq�-��c�]��&��೤J�4i؟�x;�.o��P��:��ER٥%��9��Ƣ�X�s�UQ���ܦc��t��Yף#����c�)&g�C�x:�]ԭ�O*uW}(�`������1c��A��GK|M��,7l�(������7�}�e�T2���캹����]�b�z֒�6{_\۲7���W|G���؏G��g.�C�k��嘋�bCp0�����*�ŉ������꫘�
��ؖ9! �ORg�ˮ�!�.�;t�Ei��.,1*�!�MԜ�B24|�_���w�XvY��dS<�덡�*����_�P�,`u�N�1�K�ݹ���N�u���{���.���t��4�*@�$���g��a���C���Wk��e����7���e���<:�2�D�T���6D�R�N�f�	\c#׸.�8���>��CC�U��_���y��}�2(Ds%�͉����C�~7�7���b{-�+�,�ᙢa�bX�oj�%�<y (u g�]H��B׊�1���TM;�R��
u����HN-V����=�1bb7�U�͛�mP�y@C�̀�xF����b�rЖ#��F>�U4\���轅;\0�����3� 3�EJ9TfE짽Ge�f�Qq�v3�$�F Xn>���|rX��U�"�\�3����yu<��N��89�w=�[	%ג:!�R�f�ڱW��M��ePB�[�[����XV]_/
+1Ӄ;�җy=�-�Qé�J
�Ы�E��r��3�� ��H)f�C`�P���{9�M�7��g�]/9��+f���=O��_������V�����:���K��z.��\�r��w��@ĩYI�Gb�D]���w����6%�D2� ,�)���i��J��,(�O�UU��r�of�f�+ �ELR Wʛ�@o�@鶯���.įv�n�����?�u��אU��+�kw�5��g� �X�����3�������B������mW�]�2��歨���۰η!l�|�,�3Q�@�neB�l��s���t��n��9�M��2����������@y�dA�JŃ��v�ҺdΟ�C�=�h+���2��|�c��x�N����yk��i�g!�e�!���K�2������Y��P6S86�g�C��}	��r�D�Ӕu���W��0�m�)�EHz"� ��� �<ʮ�B&�7�b���{�Q嫪vP��)��@|o��0�v��=���X����m���]ω�����E*2�9�ܳ�4t�3-8��.�B��q�LJ^9@t�ED7L�,'�m�NX��,�N��&�lj�ׇ	H�dm|��h�V���nr���B�?FC҆�^u{x��6i�=�����(#a�<2�s��|�r	HmN���ɵ�5Cؠ��[w*0a�ie�9V+�y�79���`�k�)�O�$jJ�t�|�ʜnu��)	Wͪl�L��e��ŗß];�ۈ1�ޕԩU�;5�U��qp�E�E:ι�Ekx��5T��kx�rr��,�&��f�QxWh�G����諭��fZ�M�;qf���0 � v���t�U�"B��ˇ�N�Z��+�N>[��:6�����n�0��V/���9 �ݴ�rQ7I�х��un�s���<2��[TGkY{��V[N��i�x?�H�mPf!�Pz|:2~�ٕK��v�[��TV�q���)׏p�f'u
~Ru.V0mˁ�\GL�"�j���}Tf��ܒ�>�3�k�U��jVL���R�v%k�S?8Θ�Xy���� ��Ӗ-*�`_ϩ	�pd�l�ct�]�.�`;��:^�r!=�� �g�KY�Vv�,Uc:�<��ų�|��}��M����n�bŬu��D�̝RR�W�S���ԭX�GuQ;=>��ʦri��W׫7��+�V�sL;��*�{y슢�;�u���#!#p�+�3c&(!d�;�/��鑺��mM4n�/yA��ζ������$w`�Ѩ�ꌶ�d���Q�
����SY��U�\-*�f�Ί�i"�Ç'�r��T�W�D�z�1,��
��*8&��N�)�MUvE��:�;�k�s�-֍�Y���n�@�N=x�Xm�釶v��q��V�3sd�T� �}�����S�]\,�}�R�5�����]w�9)R����6X��ۢwg�b2�^6!�Ø
���l�sp������4^V�BD���_����v�uӺU��`L��Q,���-�%.��]V3�}��_}��{�<����VL���kڅp5Tp�Z%��j�Т1�CvJ)����6�o:��Z��{��	0���⸰j.S+r#j5���ԓ���Dj+����ݫC��Uλ��+��B4�H�d�F���v���8�1s5e�ݘ����Bs!P7�1��ldr�hY��yd[UN�p4w(��&��,z�tA�wC/��	���g�q�nk�+�a&��W:������V����*_[>&�Զ�F"�c=�!C��X�Uep'��/�Gl��'G�*J�}*"LpM�P	���gͿi��u�d�Y��G�\�·O�R�Ia�ki��b���P�mP���A8 �n��R�l0�Á������͉p�{�%�
���)30���̴3�Qf�������ِp��u��oB5җ�1����аW��Z��cׇ�:�ͦ*�9�5��k�u(�����
ˊ-�C��筛2��&�> h�k����\�+̫�3�Ui��*����Yp�6a�k,�|�p�>wè�y�6�X9�̘�a�!��}tI�V��ӓ��c��,���-Vo~[���coZvjs���eJ��(�x�G�+�I���Gc��z��lI��+�/1�Wͽ�D75,���ݣMB0���KѝٍN�n�sIk�D�˩AJ���6�[m��	�j��=ކYh����Ggf��>�a��rtA��{��]w~Pua{~5H�np��o��9PN�h�'#7{�n���э,��m]�j1l���׆n'a\�͒+��uF��<�Z���5�J�uZa!{���6d��4��Z�D�,�\�}Z�]�5it�}����;J�J��R���9u�ҷ��6���עi��"5t�)���SL�L���&cgwm�ҽ��8�v]�3uf��|滛���a����i�ul$ѕ�d�� ���zM�
�1Uȉ�
hR��b,۶��A���w�T��@}b#�ojT�sr�C�[���ݰ��U������HcNL��>�/u���RZϹ[��=��[��X^�ٝaB0�b����|�GZή���"�����}�ھ�,
 ���-]\�^V�)u���?#ʸx���;2��ʂ����	���vV��u�aQ�+�S�O������T��!���Z�J�)�Ep�P��˩���E@R9ʭ�.q&FV,��>I�ԑ�wR
y>īc�3�6��XM��ҦDL���Hwy��4kyf��j�#bM��qT�{��s8	��F�D��e�u�1��J\;*v�%��uk�VrЂ���h-w9�v�Y%q��嗕��� ��si�ھ�� ���">}J�fLۺ�#�	74�t['-x��Zƽ�K��e:�H�!ʝq�T	}v5��d�K��s\ȣlr�x{L�Pf��;IŮ�\��U�ݤ���3p��_T^���'s�o�6 (�x���@w/�ĩݫ�Pq�w+n����P��ӌ�����:�ylgyz��n!n������.`�$װ�0 �v� ��k{�(LmfhaR�g��ڷ��|GwJX�VR�]�PC���׫^r�io�w��{M���n���Q嵭l�Plvrԕ ��A�B�VR�!��kM�n���>k�rf��z�n|xkGti$T�5Vn�3-�%o+R��Z��N�k�;�#C�;v_Ʈ�c��ϋ}�w47#��f���9:Z/�*�ѬVH�5��)�u�oF��W��¢��|YX�+����v;9ӕ�^Ų'��n] K��o�8r���)�B�y�k pf���[0���zN�����l}�!��:�H�8#Z��48�[�
�	'T��VMDn��j�+���
-u�ӊ�9�1.��(���5�ڗ�>o�fW�i�]�&��ؿ��� bUEU�RcX��QV�AA�UR1@TE��U"�1�,�E%kZR�Dd*�0RTEQ�� ���"��*�PUQb�X�EEQ@�TEDU*Ȫ(�X����aQ�*(*�*��
�UEPX�V,*�ň�Q`����@�*UJ���T*�QE"
-������(�Dr�e[e�!R)c��,QEU���b�J��q�QEaR��
фQDAB�`�\k�5�6�B�P*T���*
�R*�Y��)���R���ʨ���T�"ŭ��T+aP\��iP%d�"$PY)h�(�b��dY�%_43�\�����s�0����ޣy�)�3��FC�e�Ջw���O:I*�r�u
��U���5�<o/��A��}U�U}U�7�˞���1X���g<x�J�m![=����װ����
� b�Ъ�����/g��^v�`�p������Zr�\5�ò�(�%a�S#��g>E��p��
�bY�ycٳ�Q��\B���\����8bwX6������
�ˢeE�{i�o+�=|��w�Q�H�j.eg>�Uܥ���)��(1Ъ��ϹmR6�v[3���is���/T.�窨��t_)BL�jڅc�-9D1�m�b.HUnn��}O�w^N�3իE��|v{Y���e�6���u*{������T�͊"�oY7�!�^T��F�*�]4�x���ʌ�t,�='�]�;+�n�u��G/G���m� ���)u����6b�#Pܲ�5B9eOL���;0�Q�9�����!.nx�g��-	c|����:w\x�a��'Pq��iv��w9v�{��~i%SĻ�8˦�������:����L�U���9�<U{��h=ƕ�ghn�<��٦lس�s��ey^fQ��
���	���%T	<��g�]ƹVM�&��a��ĳNo��g"��ˀ�0���*b���Y0�yǉH�����L�GdZY��l���v�VV��]ݭb�Ǖ����!���.�;v�.����g.ܨ! ]*�A~�������H�P��L��y��mv�X��
�7z�I�}8r�'I��=Vi:�ڭF��f�����iu^b�zg�X���PU�78�cB��e��KTmN;�l���u��_m�׷���ǵ�A��BP��5DsVI��Ƴ������6��6����m��D[�\t���V,�L�7�w^5��v�k��%�Z��*;���|6m�5�xr��r����Ź��|	Cԯ+[H/@��B�b꯱�:�z�#�[���;F�gBm��5�
�[)]���JƸ��q�u�9V�����D[O�>w�Oӱ���q�H�9#ڵs۳��.�{�W<kؕ�U���q�Έ��Rv��kyQ���b��>��]�E�*�&�5��l?)��7'z&)���jg��(�pF��n1�5+}'%��7�U��m�a�"�m���J+���}��걓�M�:�Ǵ�[���v��@�y�.]��g3ni����r��޽�Nb��]��GYfKU���8�y���Nf��4ECi��gj�4z�].���Ԕf��<7v��u7�/�?)]\7_'��G ��;���o�Q-���W�}_WM��ǫ�F��߻�F���)�t8%�Ά���'f��V4��ֹmr\�;���u�V�LVꯔ���r�q��nYV0%�Lh{��wyL���I�*c5�|e�bu���:ݲ���z��a�輙��a�>�ީ� �>��zX�~F��+��b7�;�=N��e�Z���s��8��N9X��<b�C�K*ؕ�9�'�w�);���3�sz����)�g���3;�|9C��!��`��3���}�ieE����K�������g�A/f���kS|��C6�p�#M�`K@u��o�~ZR�L ��s7�V��@�zzF��bs�۽R=G7���C��{^ˋ��&�͹��?b3��9�ƌ�Y�����M��N����X�Cx0��ʠ���/1��)R V�2��u��}�WR���YFuel���9*�^�����Z���@�]�݀d!
���:���L�z�*��gP�=q��P�rb�����m*b�>xF����h,����PS*8����`�#`���).}���
�+��FË�ܡ�n�����ꪣ۵�)��9�>�VM��dU�ʹ��Vq�F(�Q���O�ڛ��_���.��.Ι�^*wkk��War��`��^LE�*�����>W3�!���H����q�e�4��S}P��-�ֶ%#I��3��̪���0M����i|������;�ޡ�S6���$QbwM�왹se��ǫ:�۬���q�gM~}�o�5��^[E�v;
IX3�Vfվ$R�������%���J�8�KG����eC��t��Ґ���՚�g.��e�8�W^�}�Bz��/L�o�?H��3r�C�D�����d��7�/�&����S��s������;���9���k��ǝNo�^u+yΰ���)خ,��9z��ɦ��}24��Vs|���o��@۟� ��w�}e\s�zR������]3�y]���\k�Q��R���J��F��u۹K����ej�|Tξ�#�⡺���c���J�'>ho!�r�b��	�=Gk��tc4PpVٮT`�&�w�G���n^��0V,�Yy�t�2��9�����h�;kt�Kv��pUMjE&�b�)"������HT�O���>���vOk���a�X�����P�����5�6WFsv%L<�įgn�'������o�.Ҡ��bc��z�:z��f�V�7��oxAV.��/�����,����}�v��r������Dj�qu�ʆ%��ʒ��z���wFt�m���߽��>}�fb�{��������m#s�{_v�?��]-W�ͧ���[S�6hz���|qv�=���~�C|R�QX�s|]�~C��e�TG:{)��j�n`����}�n�W�+��on��s6Pz��W�`�v�F�����i��y��c���%@_-�����}]�j�V9����_Y�Qe�R����k�ވSݗ�Knm�:ֻ��Sˑ���+_p�P�Bۉ�3�O���N�j��/���^u�i�%����C���F������ZT2�ipR��������s� ��1�.��q]
d�V��Wտ�m�-C'#��t��^jb�pY�m��ʊ�C�9�����e_ӭ��w�'�Ѥ��'�oo��a+c�	E����7�T�c�|��-�L���q�H�
��HL(ɽ��1���[	A�=��}��Oe��u:��^�m���r��*���*$��y��\�M҆%K.��E��oGgk�l*����B��Ӕc!�Fj�j��zU�a杢�����O\��ݾI?�,��5۫T�v�h��E�JQ���هusYˮ���is����b_f\�!V�9n!5SM&7�Ʀ�ƃa0��T�f��+{��"�H����eZk��bǰ�7�*�L�C}^��s9�K����?:��ORͥ����Cz3@��)q�����I�|g*ST��f+:h�}5]�����M
"ހ��r�F�ؼ�W�j5�"��
������^1��:M�J��t��NC�{�i�nm{�������\Z�����L�v$Vo���k�?sNT9�Ry��3�=�ץ�t����Qǘ���}崟�W����)MO?�q�Z�����7�'�[������{�Y��\f��b�\n��G՚����u�+N�3������y�nIB���v��an��U����'+ki�7�|@���z�L�_A'<M����N;�N�1����foj65�^3�\����`z�q�6G5�l���{Y�y+��g��Wg]��ˤ����}_W�مa���`��	������c�(�]������D7��ߨ����8GT�}�y����~J���V���Z�E�U�����*�ky���g)w��rosv�5�݇�Ī�6�5��9Y������#\��Ȇ��[���os���dCy5*���ʴóW��c���c��䟡�G[g^�]���q)Wѽ����?'M�ð�p0$�re���1�3yW^+�N�䯱t�[������	<ӹP����*rIY`Bأͬ{J!X��S�!>��.���1%:���h�n5us�oI%J��V�e�q7B����@�Y_O+^_��e�5es�Nv����JtH�oW�OS��Z\�q��,���f�U�bWd�b{�].dݙ��S:��v�Ug^�w�}e\:�����x\�#yiK��~�S�ܾy�s�!�\%�#�1q�� ��
;���p$k�w�������V�F��A���~��K���k"ޛԫ�gV��RDT�wAp�P�}�Fc5�k�j�ʈ�Pɣ�
2nȋ}��yݨ:�ﾯ�ﾁ�b�x��yr}�,��v�!�}�i°9�J�/�K�S�:��{�79ga�׋tOk�S��j5h3ܥv�T�Q�nq�V*��p�&�Gl�{ͮ�Z���ͻ���������j����Ϟz��5UOu�#���2��0t�x�xXW�m������9��1E��Td�(��oDi�H�Whv���l�>����uܭ�^�*�B�B����o�ynP.�Ó�J�Z�(�蛿}FwF�y���~r�rxo�������8f��^$�[�o�pM�/I�F�{��V��5�9�u-�T��_i���@{S��{��C����R��>�z�TO.�]-�BU�o�V�bT�Xq��ط�u��.59���/�Q������]���[�Sh��c�S0q]�E=eҋ��5����P��M�K�}i���t��I��.N�\���bT&�~�/v�rk�>�sV;��y�x']1i�q/��'H���k����,�s2�s˼Geﮔ=<�+	���ʼ�*��l^�\7p����v� ʺʾ5˜�c��j����:�}m�U�/8�Y�N����UW�}�n�f:Ƨ�ԅNl�x+R��rʉ<9�d��VhZ���3�V�[�a��;���b8J���*ن�rʞV���{�,�>f�DS��s� ^������^�oaT[�I������ɦ[2f�[|�]*yl��[�\�o0�j���j��U��1*��q2��>��\EC̛O�ث��=b��9�y�AW˙n��l䧫�qL��S8�9�1:���)��]�me^c���ŀ�V'_C������z�+��\����<X���[kEj�l�]���<�ڋ�w�������o{iBR��V���W˝Y���zA<�b�����k}���j��iX�(ǻ
�0��cT���H�^F�WC���-T]��͟{ݑρ*�qu����_ET�J��qZz���=yz�zս�ޓ}�?CrQ�9��%pZ�vst��N)�٬꜒�8�7���N�:�ΰ)�`�޷�s�;tA\@HI΍�)Y��.������B���l������TB��;egov|�Y#6����:�s�#y�(��<���j�;%��4L�޽��z�v����J��l�m	�˻���ﾪ�؊�W�D����}g}j9��V.n���oT4�����` u�ԯ�WK���8�xi��K����ڥF�{���ꊤ]:]��\sXܓ��X�k�պ����,ߦ���M>J�S�Z�᫲��T��'t�,͗���pnR�v��hYM�w^�"�՛'�
���C���ֳ{b���qկ��o�v�8�n���[�@��t+�='�[���Y�ڷ�ǺN�7Z�����e�Ro���N��Ꜭ�ܑuY[=�D��^��z�;ʝ
��˸�\@n{uR�n�g4u�����r�7M��إ�zL�^K�Rо:��������O2�
���]D>j�L��r3�=�1�׋�sԍ��'.��_D%�}Ú�3��s�ATrf�t�L�K*����ލ���ڣhuBpD�L�����"�:��3���R�{�g�ކ�x����l�Qt�<}��]��������|�=ـcYʥ�i[Z�7�����=g�k�'�/oxZ��h�O����P��n�@B�F��z��J�WîrtWU�O�Q[���T���[0�D+���W�ⷩ�E!r���4��p�W���׽��-�E�Q�C�*[Y(�z�+E�����$�x�84[F)fo�]՝ ���!'�E5�15{c 47��C{��s%��@���4i�N�Z;��O�ܩ Fv��%��ǋ�b�>�*�1�J 5��DͶ��V�0uGՁ�',�+ge�KUi�1��}Ƃ�*-���Uv^�T6�;�[2�d�V�N�Ӭ���p��@�XmmU䙎eno[�l,��%��YY�ʇ2֩^�CBy>=�b%iL:A�Yqߴ�Ĝ�>;�1�Bg���51On�� �6�͍;�����*9B��K�vsP�yLQG��'�x�c��M��:=����X� ��ICN`�J����&�%Yʯ�7�C^k'59�����ta\�*iʎ����TKV�9�%�����eCv�zv�T��=Z�q_6�WM��52V���R��7M���sRt��2��.�I���(P�|��>�J;{��5�*�v���-��O�7� �V�Q��X���Iyeq�ի� ��2�SFvI�v*�}�Xp�l�b�)�CYR�;ZwU����_�����6��)5��}J�(i�W��RR���^ ��I��`�>u���c��2��ݎ�M��<m�������3�R�o3w�m�u�=��ބk=�y]ݜ�uc"�����L�\���{H��. �7��Ix�Tʶ���1�(�D���;���ܬHza��-�)t}O^��:�)�)Ų�R݉^`�w���:7|��;��iRZ��R�w(����)�;��۩�8PQ�b��x8m��F$��3�:4k�䆱�$���L�9��t��9W%@w�,m�V�ot&�}�a��[Y.@��a�LW%\����I�g�1.NFsZ�^�kO45Z�s�@�<���n�Y.�$u��X��r]��Q��������^nC�M�IB��7��hZ�8yւ)����kV���FѠr�*��sc5�)ѵ��QAq+5��Y8��`���Bi���u�:�����kV�D �E�{���*�&RY���D|�ٝkvY$�D�!���bt���6�A@��i�[�Z�{M*��.� gX'`͍�ū��v����ifܵ�,���]���ۼT�5J�>�#�h���A�`H@���Sz7���9� ���=�F��
�6:T���q��X4 )����ۼ[�^V��׏Z\�F����k����m)',P���=ݺ�V����vzU�PD�_2;6�\78���6Ę�%;mn�:�'�oT�W�n[����.�b�)r��њ�Qn������;��6��M�r5�� #�Hz�`�P� ��*1`�VAT&�
E��r�D$W-E�r�1�J2,�c��e�ԣ
5��K%J�mR�Ab�
��R�P�\q��C%a�PЩX��EE%HJ�Kq����+"�X�X%`�J�Z(���,����ĭBV
,P\f&$QH�Ԙ�1Ua��Q�
�[d����
3P�YRT��偖�[�)*\����Z�e��"̶6��a�B��
��b�a�+e�ieT*VT���0*TT�Dci+ X��U��Ȕ��B�+��I���"�S�d��J�V��&7,�
�̳����F��f��3���=u�7ۡ;g6V�WGD��x�j9���Tc̕����Xm����IɎ���S��Lۍa��������������'yÿ}}#^5�ͺG��|[/�������^w����0�<��+|ĵ��������!�C�:����`��5�ۨr;+����e��T�Q�Km���r��9Q��Q�*/����s�ٸe/q��"��i��K��[��|59����qo~:�*#5DҦ��]M_N��L��7���)��Y-^��+��%r�VL\⯬���4��\ثi�����FJ˃ct��	GMS�v��v��`J�N`뛃Z�E�U_+�+����#�38l�}��j���n6�"��5�ἿB�y��{���X���ua�C��¯\���|�k�]�jw��>��[ԏ��a�#ж��Y�t�/.���GE���qOq]�	�f��:�u��`�e�ɬ˧j�>x�gk�1�ě��|��t�[��Ɏ�q�&�#Iew��QId��\*����>��v�6�* 23��2�r<�n��r/3[]�ô)+2�m:L�w,ʙ�B���8�T��+�{]�2��x����Q�5No���B��`��՜�s�j��g�����h��+wv{�㡾9w��iW�8�3�w� �}�3r��}�����6� ��ӳ����@�yQ=2���19��
�Z�Cs��\�H�.r��(<��d�b��p�1�>�	eD𕬫�H�s��"Tr-���kML~~�Q��sY��:��0�\�}�m�����Wd�y�j�Q;����QM+����a\&�i�7_���N
/�J����1�Yǟ(�R���a_c�ד�j��P�OB�&�7�  �PF�P��Ĩvv�"S�����F�~�Na+�q�踶��؆^�%(�n$�j��K2Ql�]}k^NTbzuFu�w	N�|��(^��R{6��>N{E�c�>V����l���qM>ŵK�{i�#:�,���C�9�g�sӹ��+�qs�xD�����*�*�qq��E�!����T����]�t����HW����y��f���0%p�0u�������#\*#�R�v&K	O�w������-�Z��髝J@;����s�]��;B�o����̩�F,�p�ٮiN�S�r���	ěZ���N�֛�i�|��O'$�����yhÄ�����\'a�׊�\��ar�7fG�g�}�>t�6�/n�}�����tE�or���Jŭf.Q#��kꌰ�<����T8�[VS��+����=�"��k�
/w�=������o�%y�������N��Κ�����-=�=3�0�8/و��]y/����g�T���B��N��.�ˈ�����I�.a��ef��(��]
������z`�밹��>���s+�u�����]v�R�ޠ�dΞb�|���w������8�k�CJ������e�Je�ď��d�=�3��!��{
��b�f3�.����Ή�@:�{IK=9���_��x��u~9[�:o����|�]�2��n�UVJ��}谹=�{��U�x��{6���ޠ�9�SN\6�S��kF�85�'u�5�V�5~nH��'�ዬ}�����1�������u�T5؜�
�ECq�r�8�&M�E2�qb)�����Ղ����a\>�0�=��QZ��D�-��E 2�=Q�~���ou;���3��Ժ��u���)k����
�{k�\��(��`{ԡ{��x����h������R��U%��5^�"">��W9�ۍ����Br��\z|��;��Qy9X�⌍�π�A��^���@��wT��{���]*���׼�o��[츷����Pt�f�Â��Z �Pb)�EGs��9���V���l�QP�q߮Vx��ؓg�������w��^�<�}R���[z�v��Qk
�	8ط���+ �W;�b)ɍRE+z�e8����*Ҳ�\�^4��C���kb�p��nZAJ֎�5i¬��K��6�\M�����<���j�P5<�m6�d1S8kV^�IE=\v���g�����ٝ\���t�,)��N�� ��'h�>i)5���;��m�R�u�������&�]�KW Om��`���qp�2���{�׫^U�5��~=NU��SauI�k�d���v�=\���\���}}<WLK��~�=�#lӤj�U�05A��7�X�fˍ��f�f�F+����W`���i�<��Z���fM��,��[��4�R�ʞ�{���!�wgLB�����w{58�Eۻ�봛G�wì}�u�����j��:��f�bz���m�B�>��z��&�<�i��*㭬�����E3i��խ}�߾�̴�M�Y	�n�]\�3��
)��.2w��[m!�jw{+��b��'�W-�9�꯽�
�y�M�;�<L��5���F�03Gs���|�&)W���e^Sb��,{a\��fK�y���3˧hs]�`�s��{�lL5��{CziK����\�O��s�q��?��������wJ7�ge|6 ����[��'&�F��V�٭z�7T��$���v����1��1��}�C����C׷V�n�Xۧ#���xnU�s���$G�=�o�TV-]�5��QQ����w��MBxqZJ���s;��p�Z��wQs���Ub�z��,ꊎT�[�R���梪�u\n"Vk�ng%�j�駣� 厨��s������/a�͋(,	e�[mk��7���y��͇�:�`I�Ƣq�g}e�{&��c+�)#�c��״���b@�}����:�;#gsV:�����X�4,^��q7iP.�q+538E�/�T��g�`Ǉ]y��fWN��Щ�q��X�Y�V����q_Z���h|�3W�4ٶXi�4��t����`F��yK.U�N����x}G�r�b��ɿ@��㚆��S">�C�/^v�a�h��R�xo��R�q���O�O[5�{���ҭ���zm�oj ��p;
�Þ�T-���R7��I՛\η!f�P�bk[Sx�~�x�.��[��u�BV.�j"���̔멧��M8eGmɹ���Qk�Z��>��U޶�z�H�����!�X��e֘�ïၪ�����ς�Ns�:��r��7�d�7{�R�����R���z�Cʘ���gB��,≯
�:���H�[7���tv�2�{��q���r�+�.�4����%nF6);���3���}7jve�תCI�a�}e\:f�Z�x_�2�o�4����e=7t"���ޝ�w��Qv7��|jL^M��E8T@umтs�ё,�*��ex�:L׶��-��ڢ��~v2�9���Ʃ+��fڰ���+�tvIς����9*���QH�5��)��{�6��骉=[�F���/�Ӝ3��?V����c)^:�k՘��?5�2�Ǧ�'��#oU����[p�d����z���8cX8e2�6��OC{ �����f��O�#���&�]]��s�V��8at��+��ﱽ�oy[�[���@u�9�q�[�W������]7q�W8�'qձH]�=��N*��0��r���,�8��v�ns[�Q����*��'�񵗑++08ky�t���ܭ�^�*��������atցr�]胯&V\c�*-7��>�5�5���*r�u�/Y6�r�?&z�|�e��]���q�m.o1�آ��7�ٸ���9�rU֍��ۙ��zU�|�q9��*[�U��-���9�W���n585f�3�����1bqn�N��;�J)�VV��cWu��>ی����uu�w�\a�7�X\��P����/O{�]5����g=W+[�a��ƶZz2�!�P�:[��_rDv����P� �k�_[��#u��;E���R�}q	�x�U}n�M$:����y���1S��b^�_�v4�:��]��S���@�k��������j���*&�j7��֔tR[�Q�f���|�Q�:�ew;Z݊5�V�����R�����8�-9-�Yϛ��r�t3��2����M�x�8�wLg�D}$�{���^:����f��w:s��c����e�"�OH[�򙛨3��A���'	���X��s���o����}q��wk��k4�W@�*Yp��t�]�o��=��Ŏk�Y;�e&}�"�h�C6'/�(�W��5u	�e��}W���X�s���pDTޮ��]^�+��}�z�8IA�ͽ���U�Ж\z|�o���^NTF/ѹjCg������S��:��C�犥���ܨr;*+�z��5�������`3�%{^B�Q����
پ�����W��~0o�y�[<�g��*�9�8���ٵ�F_a�U)��:�[U�1m1�_T=�Y�-�xǿy˓��,��T����Uvo�C���/'��U��un9hW����ƚ�W�`GwN�va{er�,i5ﳫ���s�4l�R�{����>Χ�!�\^{uae�y�f��d�l0�0�Y#0vK�Ϩ��8M��ua��Q.�:T߁��zװg�-�e�z�b�}��B�6&̴�A��.�]ҝ;kv�1�uq�u��|�1J�<�a�:к��j�X.-��r�yj���s�8�_8R���[z�U}�Ճo���9��-�x���q澉t)�U�ME��D�O���O�h�a@�]J�V�xO-����Y��������� v�B��eB��$��J��<��;�=5��6p�૷2q'�<u4���یq��t�u9]T:f���XU�*���5��Twu<]5�B��y�_��]#_5(���*�e�k2wFխgw�+��:�Yo�SU`]�p��uR�m����*$f)wX��*k�И���hC���[y1\�̿�'�
�y�\ں)�9�ycG'�l��E��:�i�q���S1Q�ۃK*-�]�ռ��ov��V���kE��.P���vQ�v�L?�f��Q������8�N���Gv#=\�/qwʵ�Um���z�N6*��U�_m�{��5U�!��^�ײ	�s{�>v2�u
����>��{�i���kk���l��3�1 �,��B���a��NŖ�P<oY�/y�"�w�VV�;#P��}���d������6����U�e�uhAZ_{@ ��:�5lG��4�#�N�vj�*��!�u�RJ�o^��z����ۖ�v-Kmܡ�в�����a~����m����˳߾�O>ҧ+Ӫ3;-E��������2t:O*9���L������P���w�����SO��R�^��Y�}YU<��NIH�#d��Q�T���B�P��x��Y�>8�H^��;i�%�{����p�~>i��]���w=�tw
V�|�`��nkUg�צ���}�){���Gc9[m5���}
k�n!�}Q�J�S|���8Z�������;{�:Z]V_+�V�jyqC��7V���+�L;ug$��+8�a|�彋�O�P~��?S�u<T9w-s��L'M�L22λ�Y:��L�;��っR
n��^��F�L�N#�mWz߻:����j�[�.0ĸ�Xj9U*Y��_d��M__DW{�`���(k��z�$�����:ۍU�J�S�U7������w�����#d�6�ō�����M�N��	�urz�w[�Xr�c^�Y��\Ge\����_�/�21i[�F0�i�ݙ S�D�sm<�v<A�;4K������8�Ⅲ��zR�Ʊ���Y�� Vo�����,U�<�֛ ��L(����Ϳ��6�T�"�;��2�r��L�v���o6�8N��b�x�����qv����v5�����H�	�r�B���k�E�\�N�d��:�t:�XwW�������u�ˣec�*Ð� �[�8h�����cXRP.���������sl�w�i������,�6����g��PMޒ��0g&g.��"�#�WW,u��A��h>]z�-��hgv`S,����h�/gwv���ӳ��@�:�v�����7�gE�ֵnt����Gȼ7;�oC����V���k�3{r�	���XV[�� j�q����o+T;`T��D&�����T���r龨�*�6ՙ��AV��W+��E��yԋ�m��c]66��|y��Ȼ�3��v�8Wv��L�x�v-�|e�����C6b��VT���F.k^�飴�ۘT��%�P�4��9�^h�W���wvo�ui�y>j�/N4ox_V"�hwK��Jv�F<�Jɘ�:�N�MRJ�;9�Z�f:��jq<�Le�Ւ��o��jDdY�2�&[ԯ��Y%�� ���u^`ٹ����j{��&�K;jhۤ�kIP�9�.e�x��Ƭ����t�,=#e��Ń8ul��q�]�/�T�O�	�̿�8��Zێ���wwD�n�pz�����T��T�eu	kB��#�2���U�����T��t����f�q�٩�y��彩�nƪg�����85χ��I��ܛ�OQ��������\$g�����hy��Ѓ�N4�bv#�.�}�ȵ@�F�e�IWo:�;���x�si��8�O C�o�ո�؋8V����c�nvS�o�,<#<uP���*�s��N&t��h�5�/wBea��J��� ]���Y����eI���;�/L2Q9��3�i���`�7K�ٛ��w2��yO]�	|s��=��t��9&�\���T:�#s��w��:�g�=֮H�6F���������*j�C��V��I夔XՃ:��_7�Q*�F��k�����4�H�.3[����V��|y�j�|5D�y�t��2.���K5���W,UzH�0��r���5�2����pCQcʉ���U�f�]�淸����P�-�Z/�I�\���|{�]�ߤ��3U�j�8�QO�t���y���,������=ଠ���Rk��1\��9��I��lr���kWn��.�G��u��6��R9|�	F�EK6���>��\>�]93jP���J*��	������Ŵ�FRo(P��ʓ��zS�(-�}Ub�� �4�i�
�ۍ��m���9dR��HZPih�m*+
#hQ*
H�m�Ȳ�YE$������Z�%�J��d�DĊ5i�LaY����
��²�`�P��5,�V-b0���0r�r&e$�S,�@�%�m��
�
�)V9E�[*e¨�iV
!X��c"�JʅdU�،cPPXڌ��*�A��js.G)(�J�����J0QAem�#QUV���DB[aVڒ�@LV��)Z�c�[l��
ƴ��j�aY1*AA`�ZJեPk%���R�VT�@���5��PFJ[�P�@Y
ʑEQ[k����X�S0�"�>���O��޵������i��`MZ:>�;y55\���h�y:�/u ��wls�T���s�"��A�b�n������Mߣ���������t��f�Q�Ќ��LGM�F����k�U�~��{UFa��,�%�j���7�*IӰ�>
��5S<7�۴3Ɗv#����b�n%G^d������-i�ǎk�y;�Dj���P�A4�.6������K��j@�AKv��TE�:�{Z���+�z�8����Ԝ��7/�S[�4۴�*���hy�m�}��j���������+��ܸ�|�.���$�V5�7�1�4�eŴ�����Խ[�}�V���*��[���b�25���Ӥ����_K��{�fJ��.�+�=����������� ��fd+�5K�LD_�����x����+��_q�ؕ��k����K1�N$;9��vyŜu{�ƕ��<�kMc�MՐ��q�M��C�.c{�5���U')�f���:ݎT���|5;�o�:���������;��ou�*��@&��r3�,*Ǖ.d㚝�&�fJ	��Պ��DЯ���.��D*t�KJyS�F��]3���N��B��I5b��q&Ṿ�K��u�u�7���j^�SX:F�5}f���[?������j���B��-�egO�c��	H�,؛�J.�%�v5:�>�����y���v�G����N���	\�P�bM��.�Zk1p�eA��ro.{�/��I��}�2i�V�W_r���y��鞻�QӖ����s��qʳBկ�y�61�M(��S0��%����w�m��m.Ŷp �32�y����_B��h�p�«v&��T�2��Q�7Ob�63��"��0e�MF'�a^�0��F�j��B��wblN�;�R����\�w�AŵC|ʾ�/c�so�xMs��V��|�:����6�Sn�
�c�9R%�ly_^b�gc1�����d+���H:���fw8�ty�zN�e໏�9��|���j�E���V� � ���=MI��P.���5z�\[�z��T�x2����vW��
��1lX�<bU;���x�1��:��P50ҙ}\c�&���������c���۽G�&�J9n��%���[���K޻ou:��ԯ�9[�1a	D�O%7��qEHԠ��݀tQ�6"�eż�7�h�죍hW��x:�|gj=";�*�V��Nj��
�$�P�����Y�(\�jNq�QkѪu(��x�g�^���#Y��9�=����M���=��]��3y��Q����.ߘ�/����w�߽�?^4=y���ah^['���r��m{�+��3x��ꊾ��E�oh8�f�t��&�_&Tq�ҫq���F�R���Q:�J��F�]<^�l�Q[UJ9��S�{N3RQW���f�~����z��ήch�9YQO��YY��t�G�t��X�8��_�m�wͽ�����<���@�YQ'M�(������.R�vyt�/?w��C�ݸ���n�nU�	˻��DU�ӚÍD9���Ȥ�+����]�[��zCU;ӯɷ��eZ�85l��Pэls�t�`�b9�}=2���2�	�v�:���V��^m_�)'Xvs�]\'��¹S�5��p��p��@W?o2�F9�Z\�\�ؘ�+�q�D �5��S�=;��tK� �Y��k�Zo�I��U��)VZq(����&i`��{�f���no�T�?V�.�.�&��]����R�wtSw�eR'�B����zf��=���꯫ճ�D�?U�O*����Je�m����߫��ر�t8q+�a�㫲j�%���j��ʯ���
�p���7ѐyiK�i�m߳�/e�w��ma[�gސ���ڃ�N;��	��u�9}���vٌ}�(d��#I8��x�~נ�ؠ�=��G)*3�W��M5�4�ᚬ\ӊ�b�F&e:@@�u촶��O>ұm.���T;տI��0��
rz��|�#���A����r�o�҂�qM?��.�����RO�����[6�)P��J{�!�,�{�:������?W�+��9g�qv����r�E]���QԳ�fd�Ɛ���|�6��[>�6�+�=�\G_��#�B�;ɳx�-����zq=eto.��lS��~3��K�>� ށk��a1|�M��=;
�͇�kuW;�V�jyp�>��ts�\C��U.!��6_� ��*cx#|��s(e�K(��^['��A�ݙr���K�^^Cr'����z��t��Z����gerN��gw-��ү�F��A���&��ݜ��r2�i�*M�Y}X����.�w�jt
�*�w;3��%�)ҸY��惘b��KT\��k�#���\D󉈮�w[ٮ��(}�m�{��8�ad`a����'�D�\�����C=\���\+�\��t��E��eq��d�)�v7KR����E�T�D'.T`K�WՓ+�5U�D��׃��93�X�9���'�!�9�jE;x�a�����%���
�6Ƽ{�9~�L�(��\=;�;-����w_7biK1�.�4�%Ԏ[پ����~�,�S�׵S�}�$��z������-�`�+gOdb����],D���\����iZR��3�\�ּ���*�!�6����t�騢F����5=Z�ݕv��H�x��i^{��a>�;�}��#����+	���{
s����OW�75�{.-�.;���I=5����gwJX{1��mn7���1N�_ϑ��a�oW�����8�
3�B�뫩���
�Z��CV���#$���zL�Þ��>����@�#��T���m7�����Fq4H�{��\���R�=��7^p���7�%K��r�_U��o<�����s����U�*3�:���w*e.	��0�����E���Wk���}��c��WA�Go�9�����ޛ1��{_{�w"�~�2�AM��+�a%E&=<��S�A&�R�T_VC<��[��'��R�	$Z��UJ�=�Ua�9s�j�`G-��:����Zj��9�آ��%φ�xMP�W��8�i��{#spbu��ʢ��z�W�S�{�p�1��d)�aΎg���}S��ߙ��y�T,ٸ?JQ?S�2WWѯQ��bҗO,�ф���N�.F~S��gv0�CBƮ��h�wi|����
�gT����ފ[Z�4��޸�NR���U@����X :�ڝ��]�����_��;��[��N�����q��ؘ�(��3	��2s�۾�h���O�@�8�B뽀��wsG�V1���QnBC��kT�(�r� [�q�q�1m��Ɉ��ɨ�Ovg��:o����5:3U[!�P�U�Y�Bm�P��He8r�>L��,�bZ@l�ٶG@2����S |��f+s�K�w�k�����iD��6�րݎ�c�x���hF ǯfp֛̋{����p���9:�G�)���u+�JK��-tx��_}�@�]r���S��Y�`��ѐyiW�[�/b�)�o���(a�<T��Q�L�s���e:
㜹S��m�yQy����9W�pl�"ط|߼���Q��_���u^�'p���%��=���j��b��~{M���[���S��*��z�ΐ��ѧ����9#�t˞��I�彔��8�����ʌq��5A���Ws��k�v��C�GLTl.��g��
���ۗss����X���3TM*jm&�6 �2�g���J���T+����s�8�Ⱦ�Qg[�U�e.o���2������:�����6��[p�CK�;������nvߟ�y�Dc�L]k��+�6nŮǭ5ҟR�Ԩ,�{(�u��Vmq�ukݧB�&�S�:B�in��QWb��9��U7c���ZW̨[���N�#Er�FM5�Q,�Ŵ�27W@�:�k�+S����(�\P�PK0�]I��!Ѿ*�N��9En*HB���*���y�+Q��s+_X�8��=p�Ij�T��OTSk.i��\��'[37*t��b-�Ĳ��erI�{߽��<��][w76}_}����Ĺ�����~�a��4��CM+m�^�9n8ӥwP����E�,��с.��:�.�����f������/�R�8�j�w8�[0�D��2�i~��W��sj��o�O����2�'=���uVѥs�O,����.���)�o��˺E�a�w1�����e�V2gNS�T�M�\��mgK����N���U����*f+l�ʈ��a�z��\&�����af[
���a���CvUè
�ZvM��Piwcxc��⊜�������Ҝ%�c9�!b�.�mA֍�
���u�۷ԧ��x���T���]��җU��נ�b��M�.9��ܛޝ��}�bfuS��ͦ��i��vTA^:|��U.�O�}�l�~����"뺦�a�F넔m#]�r�a��,���}��M��u/m?Rn��n(�R��j.z�Il��]r�3�ghr�|4�2�ʽ��.� 3h8t}^���U�^,6�ұod�s�r�[��,u��>}�F9��Aң�V���u�}������7�9��×�y�r����휝x(��'_��<U^����N��ܭ�n:�YGiޡ�M{�Vҭ��T�����4F�����ض��D;ͦ�m��W�0%js\�\�o�ӧ2YnN-��#NmY|��=01�q��!���*���^1(4g��{�J�."nN(�|��+�r��Sˇ��{G��R�*2z�w����C�Qg@�Z�uS*�Mĥ�Ԭ]1O|9w-rg��bk~�.�q\yC���9�w�L(y�&�
\+�\���՚.��L����|���L+��b%�5�K��/�^I!=wvZ8{��iz��[�}P�[�sG\7�݈�V�Ls������|�t��ZJ<���'��Ya\����'J�&Qw
������u!�3�d]"�z�sN���=b�X��Юcz���t�5�
�u�5{���s�%�܊L��l�;�ȭLE􏆥�d�e��i|������n��0�9ȳlmh����6��f�Ȋ��;����np�W2-�ݽHMy8�6���}�O+5��{ڕJ����&.��ʗ$�i��R3i��F�>��I���u��_L�n��-�2_>2�<d|�u_vP�Cf k
���UU��]��K;��ё�m�|ä��F�ڍ�
��6�5�ܸ卛0�㒜��)īn\W�\8����yE.ߊ�ߟ;��wn��Q	rk�f��pIut���:ٷ����u�:��v���ʌOO rk SʡDS�l�[૷!�e��θ���^�t+>m��f�P\v�(��7}�w�T�ݞ�=]�!�;coFO�|�k����>���7a��E�P_"�^u��If"ewb%8پ������#KʽQ1����o���k�v�0����/o^;��υK+�=�o�Y}+>�8�,�W�m.o1�؝�]����s�v�I�qۗ��v�j_ڡ���_�c�"'m�Ϸ�U��8؏7�N�y/�՚�>��T�>S�[�E1=�Bʝ����+�]���g7Uĩ��gO;]��o����cZ���Q�.�eB��M��>��\W�ܚ�tήw�/d�����G�U;�*@�jjj��vMti}���;�ۃ6��aSu+r(-�wl�53,tQ�@ ��7Zx�A����B	p��[�.л�:C'��P�4��r!�v{*�g�����2:ʇ����@]*��Uc4p��)R�K�1� �8�fg������sv�*�TZ�[R�CN�:ݾ�Y����S�='w;�t�bn�0��otyhi�m���q$)��jK,b�~NR�W�����0�)����H����}Ў�,I���;�
����S��u�KQ�A&s[.�vrw��NJ�K�-��6+zv�w���AA�{�!�#�#Ju���f�&�R���SΓ���w��,��d_-1���	hnpF3>����z�K�+���3�Vb�q�v���+���TҴC��m�1t���Y%�
��/[�'�{Ҧ㲟7��[w��ձ1Ŏ$�Y�l^�^�P�#�;>ˆ�q�z�%waRգ���e%��B0��r��gg#��t�ł�o(۬�.���T5c5r><�5�'1��HS.�w��䒳��(ɜ�d�j��a�_m�=�!rfv[eT����]��/��FV�D�p�qu��eFԔ�*������w4mg"�>7��WP{N��tC�7Ξѭ�C�M�K$���+v�a=�X����<}�mDжr��Ԉ4���-�V��Ɂ�"o�k������9*���ﴎ��m]����ۃ�k-��
��L`;b�ZB�k�)W�k{�@�I���A��r|�`yO3�M�J�c:��z���S�e�5L�<�����V�vtG���7�TxfR�g�����/��l�i��d��'aC���b��Fi�r�C}�:j�:�I�TS�Ѽ�|���6Ս���w(R���Tj�I3D�K8^��2ЙW���.sM^ܑ���7����d�ܬr�*>�[N�J�*n�Tj�|��z��ݙ&�Y;�\R]��e�����zՊ.7xO;�j��� ��P��d�x8Ιzl����.��6LO��os�k�*�Jt�[[V*٫]��Ȝ�F9�̭�h�-U�!Í��n[v�h��a�&�^X�Ԣw-�V\]L�Sy�������{0؆S<#�t-E�X�ڣ���/^�� y5������^
��W@Ⱦ�h3	G�iC���ѥ2��Q�kTV�>�IP��!�:�=׹Cq H�a#�bн�wo5���l�cu���E�7u��J�h�Dx�+k��yq��q�0���R9�.��mf��o+ug���o^�I9�wx�Pw;�c�0ݐ�� u�êgGjΩVm��K^CS�P�k[��`�����(Eg0�`8m���|ڃ{qW;mN�R{9b�B�\���n`ͪ,w�MG����8����n�f,1
�K�PQ�9�/`B�&(Oa�r�a�ۣ�>��H��2��K��N�v��٠><)3u��FP��9Π[d=�wۆ��-e@P+F6���$��H(�(�KeJт�i<�f\a1�mUmkkJ�j���,����X�j6��������aP��TATYDV�,�"
H����.1C��R#1�*�0��D���2,�YR�VT��.41PQKl-�"UjT��`�U)JV�eIR���s,��&XfX*V�Ls,�X�S
մ���µ���9j�*Z)ܵDG0��+���ZIR�P�EUm%mKr�E+*S-�3�r6#�QU����U�R���32ŢT*����&5��R�
̶Q��q�H�*��C)e�1*GcZ\��1�al�#j�-(�VU�U�m�c�*ox���]�z�y�gt��t鼃�n�U�T�-ե�Ϲ��6��N�es�O�*.��+5P�sKo�J�!	�"#2V4BY�X��ĿG_j��ҧ�Z�q��(f�r�ܗs�]�8}'vC��{��7����3[�}p��X�E��=����
�:�vN��S`���}u足�Vy�5}6�n��WZ��u6�*l�֒a�E�j.hC�3xD��fLS"V��؞��W���o���b7iF������o3أm�WP���R�c�����)���c9�՗o(ue�h�$�Н�.�y�2�ˇ�CYӨbyӕ7�m�yQy��1C1.�yvvԶ����B����X�Juݫ�!�=Pv���qX�����zhY�k!@=`���O�;��D��ʌ����7j�qo��z����e|��쨖���jg��z�>r&m^�>ߊŴ����(��jyz��k����D�J�h�����+����m�QP��8�h��Tǖ�Օ<�v��ު�T��{,��:]q��R�� Nj�^���-���O��`و.m˧R���J�eH.VP����0�Bi�8��
���ʷJ�k;�h�9�:��԰���7Gw�*q����-P�s��;2}�c� z��S�z-v����M��,Vh��׷����WՐ����zf��.>f�+��_3�J��fr!{O�v��#�����![�ic�SXs��>m��ߣ��}���	T��뉸?V�Vy>�]b�ո_W-n��p��jw��k�=�5�7��Siz�W1�t���?.�[��v%8ĺ��U�����z�:6���^��G�ಥ�O��+&�ѕR�4}ȥ�k��o�UHʉ����W���aT_�G����@�:��4��� Q���>;qJ���B�gg�ހ��7�ۊ�T�RÄ�}��^��?JF����|���L`�����P;�P�w��!J5�d�) �v)M
����	h����mt�^Z���ٚ�EJct�k�sYG|��N�g�| w�-̹#W���A���1N{N��wO)�1;0�,����~��'���p5���x�7�����{l�z�?S��Et��ۉ�c�3�G���[���}���V��컟=2=�j���|3�
�������),�w��Q�u�*���v��H��v?�K�B�M=��굹��v���?�.+��H5�7E��Y�UH��`�s�A]Y���4�
�ͼN��c �ob�Evw/��FK�p���>�q����&Rέ����s$�8,����q.�1��o�:�>I�΃5�ǫ��VK+�dg���ٖ}�Q"�3.��W���h>.vZ�㮻ˎ�HC��[��u�*�i�&!+��s�>#�*N�N�c�Ƕb૮�oo{�0����
Az	�nd������q�Zn4���� ��e���~��{�{�vM{�n�G�nE�	�^���V�3�4�N�y[p��T�`g�zIr�.<�m���s���ݎ��g�����7���v��p���ӓ���1d֗�M��x}��MݷԖ��C]����iM���k��/K��}���1�/g� �����#x_j�.Gn���alD)L��ɔ��grU>O�������~�B-�#q.j��9@Q�Yվ����g�uN#�ʬb��@��Jf�e��w������*1Sц9ۜg"�"z�����q������/y�E���=�:�
�����]f�4o�0���$g�y+���q���Y=]�����mH<�~�S�Yq��*=2��N}FF�e��{PћQ�$@������R�}�Lz��i~:���z_Em�+���)6�e��׀v9�n$.T���I�w$�S�%cs��8��Ȳ�:^@�� Oz�L�\�j��&��:�@���f�u ��"Y	_)S�IN'u�Rm�$r�.��9ٓ�m���E�i�G�K/Ǵ�����p�U�/>$6n��L�ϸ�����X�e����xVʿT�5�ֱ~̸�u�!�,A��pw�=�ECʧD�|�0P{�]dE�A���:{��i"��['�n���xs�c+��dz�_�2���r|�@y���+�s^�<����L�d����_�&�7n2�11MVѽs�ݟF�cn5U����׍�~���.�(�ɔ��m�2kc�2��BU����?V����~g孊�_�`a��l�`Q��1s�>;����u]�_W��x�|�g��Bq%��W��l{�L>�6����f������z�V�BrLVFU滿T-�����#J�{�Z=�Q�~BJ9~�!i:X���hw�N�˯V�'r���ϸML�<X��Cl�����J7��v�n=���=���%���3n�X剚�;3}��q�ƴ�8}��,��O`_�����v>������F߻l���Ewf�?�a���I������Y�F�l��Uxe}5���ɝ���G��3��**�z�۟~��\�c���U�BY7�S�`�2VC�Н�Nuu��s��u�;�n�>ڑ-�O�U_/�L>b�nYz�9GT��]N�'�p��Z�4�9��}w¸	u�S"����S�\U�q���\���X����<�����2%՝s�����������v=���t���:���>	�T�:���NF����e��W}pD�L�����&{�ZД:�{H�6�1`tWz���e3y2����"~1��UFk��U�z�m��ґ]��� ��1Ч(���DS�sLӑG ���\�9kT��~z���ΐ�iY�>���\�2<V��������ХSL� &_�P�T���"�ft�����̜��y�tw�϶XWӡ�~��g�T�ȍ�5~�p���E���[2����UԐff��;������R}2��>��|���j�X�A���0ı���,E_���-��������F{�1:���ǶeO��s�%���r���禙�;^"�^o�4ݟEL�fE�h��]<�{2�t��R'�� <5�a�>��z_�tvyxO��^9F9n����=c�m^���N���>� ;�ʀ��� \)�}��\b�=~v�Z��yM�����n�q{����o}�b�\{����΀�9.��܀w�^�Iy���q�����3kC��<&�KV�ׯ�7��|e+�n9Y�W�[��Y�R[����I������̻[כ5V/��bB��m��]�ھ@eu\���N��
����6�<��x:�}��I��ÉZ�noW8�@�.T��`N���+�*�rޠW?��i�賚�UO����E��z���{:�:�<qu���R�!�h��������k�?�~���v�v��⳶ٿX~s�}�D���>ki�1����s��@�*r��ݵb�=�{o�7gTb�Mw(��gΤ���/�qb�f�޹}q���Ul�����=Ӂ�^���2�<�xUϘ��碴\6��Gd�YUN�=��u��r��ᷜ���bY9Yʫo<Wwu%�i�ٯ7H+��C�G��A�Ig{�Z4���n+�w�L���fU��v(�z���{�]%����v�����}���5����H-rD��0Q�����R���ul�m�R���j=3����4��^Ӟ�����#n�\ns�,���L�:t�L���Ԝ�C4+���F���6{�W�=���(~��U��G|�z���7�Q�]2�ol��ߴ{=[���>�OP��F��^.�m0�=\<=�({�'��F�jt��s1B��7"2:=w+�@��F���5
�l�9���n�B�K|KG؞׻h������W�A*����s2�"�����z���v�mwWWXKA�]Ք�������Eu���6h�(�YV��)���qU�8�v�9F�^�0䘶���jW�����M�ô�W����]>H�h�f�+i`�N����9[@.[�x��q6v+�M��:���q��%�W����u#ޟ��'�n	=��SB���%���&�`�'�|fn�:�T�/9��н�����������Y꜑B��j��s�waj�	F	��ww$�N��'��4�G�L��\��Iϥ� �=�-��H�UD4{"n��4'io����J���Ox��a���:�d��j��ڟm�'�P�6�����E��B=V&�������E2G8�p��F�9'|t�c˕Y,\s����	鿼��w�6�U�x�{��*�I�(�����L@��p�eyŭ����~�c6�����_�$�ψ1��a�R5�YW|�t���u@���p'$�}�>�J3j��c0�RR���^�y�����ogx�:����LJ7�ݺ���_�{G��ߛ"�>-䮖�tS�7Ϧs�Kb��'η]��蝖6���*�ߋ����G��X�7>^��q��o�tqT�e3@,��=uAǉ���L>C\F�f�y:�u�%��ˑ����i`�͞�c�c�{��w\qaC�[v���Z����ș���Շ��h�m�g����^ѻw��t��M�볨0�|e����0���+Os�=�:-ۭ�������R�]��-��]q�dD�3���ݿ2�=�.��h\��nI�)�ڸ�*�_kH���\��3���t}��~�� ��g��ɝ�gȼ鐪8�y��������ő���x>�_[�֧��&/ƌo�$.�"�\�UpSȁ~)�ɖ���`s�`���;k2IF�v�9I=~�+�|��%e��i��c�Y�2�}�Q�&��-��F�4j/�P�qQ��q����V,�ƙ����kb;և�z�.�\������2��������/o?_�_²���'#Z����>��~����E?IE3�������?W��$6o��ۊ�+-L�� lL��]Y�{�k��9�	T�{2���<�.�`:��z��BeF����<p��8���כ��n�>��~���5��:2�i���^�=��W���>����˂z+'%Ͻ�������dl5�H��N��7P��)��mg�v�y^�C�׍�*���f1��
��^ǵ%^�3�� ��i�>G�&�^V�y��5^�U�W�����b���,�]/T�x��v�Q�4�,��T3�<��؊v�rG���W��`���F}03.�O�jA:28�v�\$�b^���2����K���ٰ�BE��6��r�ۿ:�^_k<WA�o���M�9�,B��j�X���+{OL�7�ݺ��s�v�ܧс�ά����"��ŽEk�7�:��T��w��k �S���\��:�Wi�#�ލ�#�}�`�z��d��yQ��U��챙���ՌO��sך�y�*&�v��Jv���(	Y~��Cs]�}��Q��n�M�6��hc)O�����u����`+��6'�/i�^��i��Zn#}#}7��'�*-W���ｗ��TM}��<ae@�&�WD���>�y����l����ɭ,a;�Ѯ@��G�c:��X��}����(q
\�Ku�|�3�e�"g�3VQf=��Ϣ};����=����:��ςy�!���~�F�4��#1fTL����@߻N��L+��<�8{2P���9�S��Ț�k�p��o&X^E+������ Z��C�}��s�o���iϙ^/��~گS�Y�~�)��i��r�M�O	�~�U^Y�����GMx�w���t���|W���7>�_�m+8Ī����ʊ>n I���=a�v�<-l���޾�W�c�{:��f�n�`�S��
�Zz������HX��ܙ#�)�� �^9��������w��ԋ����#|ꉏb�'ӛ�e�Eޥl�g0�-�'�"�5%q��j���'�p&�AI&qn�T��'8M��mf�:�6����J�|Dv�0����X�Q�i��;���|��,��-�.��g,w$�gz]�kv�Ğ�/�p��
�Mk��Yo�[�έY�Doh��b[7�H�����8KGvGt�6�^QS��^��axi�U�x+kw���0_��\%pD׫��_U���𘘧մoK��ȟ�Զ�]����.o��^��}΀�l ��[�\�p��a�m����V���D��}��3�;^zv�J�w55���6�3zvݩf%����O���7^	����:��C������<�?Cu�j6X�3Z|=\�2G:��s��=��U��Q�q��K/O�_����	X�i��\�����6<z��X���N��q��5���W��뽐8�r�~]x+]*�x��(����ܞ�q1�,Ǡ�����W�x:v ��<��S�`m��@����9�3F��罥j�w�����m~����"�h����|E��UemC�OQ�r���G���1����Ï}��X����U{Ԃ'Hp���C7d���CJ���⪇��;�7	�l{"�(]��io���ʮ��}�i��K�}�ˍ�q��g�TW���ʃ������Օ��s��o?:yb1�jc��H�9YNӬ[&
���&�븺��붺tǶF��X�*kΠ����=d���ɮ��ʎrR���S�2��:��`DM�y�������s����]��t�s!tb�;:/^�Mijۙ��t�y��'����[8�M�i�D[j��nF�r��IC�3e�"��n]�"<#yd� �_V-k��:�U�����k��qq���wpY��+d�;:@�c�i0�z�����5+*}�Mp�8բ��i�"�{v�A�z�ɧ-s!��Ƹ7��5bo�I�0g3x\MoOC� �l9xJ��h��S9є��WK�#.��L����X\1�p�[Ӓ]p��&��@�Z��۾�5�ŗ�+�����fΌww�N�k�s�u'n��R�B("2�ôw1��eӵ�;MLAun)�����������"Cw1K�do�o��2�``h}}X%iD�r
���k�,@w�2��+�7�ᕒ��.+m|��t��*sr�k:=cP�Zz;�T�	�e���.�h��!���Ӽ��rd�B�p��)?��L���&JNwn�����,ؐ��l������Sl���J��S.����ζV�c�t�S�X�9���c�B��W�����r�j�Vf�a4reI�RN�z�D�%������A��J��@P%��2�[~ս���)�0nޔCw'�f�0�i�����t�i��%WL�I�`l�Y����tC��s`n��x���V"�j��Rw]�e_���j�g�}G(kh���K�!λZY�0�l�.5a.��;ϡ�ŚP�L��	��'��{LJzr�ݒ鋋��+	)���ny_��ܶS�r�uzb��2z؟A�X�3�La��Uvx�K,�Y�7L��^�\`�/�T�!g4��z+��J4E Y2G.R� ����F'��Xr�U�i.�N��ȑ*��;ڐ�׷In��ߡ�n�vֺL1�w'k6�F	a�;5=��W���&�m���'rc��yVձ��8˛��,%vZ�0VTv-���ha�TsU�w4w>3OF�λu�2�gi�P.�Zb�}(7��y�fɮ�0j�yk9��X0J���W�P.����.�'eCz��i��((9"��(R�����&�m*�;���-�k.�׹�l��\��\Ĳ�r�y�����0��o��;}�Y��/����{oe
\����zl�(X��Sm�"�Ś	���V,+6|S)w8�.��ٽŮV�uYV�^㬬^��q+a:uh¶p%!,^>�[s��wm����*�t�w_\�z�h�y�m �YY�1�`}b�� kz9Mσ=v�Z���g��X�]<f�n��8 F�a�U�՛S�K�W)�9�$e^����o&O�;�&�k�xes՜VS�ե@��j�jC�X���\�&�ER�Xi���fC��4p�ƞyM���6�L�y�w��^Ź�O21��C`��Pd�U��j ��33�eH�Kj�AjPbřj�DKJ����b�R���2��e�-��UPJ�h����S�"Ř�AV��24�[-er�b�8WV��(R�Pе��\hc-�l����%b�XQ�YQU6�VV�Kj�m�X5,��q̫iY`���m�AV���R�ڮ0�*�����EQ
�4JʕIe�[@�ƔcV�EQUT
�����UAb�T���QPX�[V"�VZ"+,Db"1,"$DUTJ���a`�Q-R�Kkj��V����F�V�LU�2��W�B�(�Ԩ���U����)b��E���"�V&Z*�X\�%�1h�>� j>Fv�/&��T*ڀ䵯0�����o��u`r+�R�k��8�[û]���	��Ys뵋�j�ZW5�WU�P�6�rus���g�(�L�zy�@�^ӟ{��Z;����x�9�,�g��㰐b2v,w�M�l�a�B�?ESb�x���,\d��U��t�
Od����u���Woz�wF:�.%yuJus�t-g�W���mi6@�W��L*�����.=�{Ǻ|f�Ջ;^���iE߀�o^�p«=Y��D�̐�D�R�Gד��qbWF_Cv�"���TW+�֙�>�Ϸ��:���x�<'�n	=��4���9�gG@&�|⢻��.�p�9��V��;g�W�� ��D�tȝt��ɸݱ Njz�ąeT���\b�m��[;�Y�^5���ߎN��9/(~�Xn��B�!����Ŋ����{���8S�>a���/L��mxv�Wܬ\6�Ʀ=�T<��r��̱�M��i�)�)�e��z�F�q��3oG�'ä�:���*�X������΄�uf���V+w.��L���� ��P��#�`J�p�|�d�G��2�L;�����<�U��̨�4�.a�{���@�ڍ��W����pA0��
�w7�\���ج)B��`�S�[��;��N�k�'�����L�z���/n2�J�:�iåގ�3�����};�r�v�f�&��"d�_.�&q�ĹԳ*���ۏ��	�Qp>��\����s�Hz@������#���wo`��Gv(_޼�.<��9qꢎ�ӵ{��6�M�����ú�ǧL��/�zy =����s�w��'���n���po�т/ۢ��y�F��]7�O_�ƈ����*���}7�k9���x�o�p����\U���<m��ǆ}���Uws��ّ�3�V�]؏�?}�X]�L�=	��W��Rף���w�v�x\6U����(����j��N���@�>�oN�V~�n�Qo���K<g֗�>��!�%S�徧�s6�y{y`~SE���r�vO:ک�]j��;ѬU3p�q9U�O�<�~���L�����g��4{1�^�I�[����D��i�G�LqR��V]G?�����`>Ț��4�QjW���q�%��<h���P[�`�v��.��������v�.4��}��de�@��K�Y�w�7��%�e8ml�g�{¡��$n�<���tW��z1̹>��CF���Qx��N_U{=^)�|���=��'0� �26}�Q}���_�s�;ģ����e�V꜐+ԝ#���u���5DWO*?7:�zڮ�~����`׏)̜���~LBj&��9/ U����40�!n�)��K�Q�����ޝ�uf�����PkwW��T;��������� zP����(�1�{]4f^��fV�M��ہ��WWPkS�g-��#������d����tg�Ҵ���G%�c��wS�^���ޭ��Sv=3K�==�=��w���A�g+�]��u��+���5[F�5χv@�3��,k~���3׳�(^����\�\��� n�i�U�{&��en�y��8S��ѻ���u��{&.G�ۿj�y��{�N�Y��P��R�����`_�$���෠b���׏��� ^��n����?�G[7�#٤Ͼ���w�-���uG�_���7{�Z=��7�$�������3�w:n�g;�{��ƞ��+�+ܪ�ޔ=�7Ł?,�d{��3�^G!���n#ʎ�?T��4����z�г�� 7o�}a�')��kJ��
Ӭ���q`n'p6-W������r7���.�1Br�>Ƀ�}���<l�,�}��ՑLf�����޹]��nu0µ^g�;|�ڎ���(���7��_3��O��zf=gъ�ɝf�ɟ�:�1ǃ��@5K#�f���Z���ζ��g�Λ=�{+�[��4d{�)���9rl7=5�z��)����56g��8'�X��|�&��-���]U�6��b���<�{U�c����RW�n�0346�d�z�
�qʷr�U��Z��L�\�'H9���UgV��D叝�+">�tu:瀝�O�񅢯3�\���&����o��=��AiBfD�.����߲�Z)߸��"�lx\:�lVD*��\k��o�̎p�<����[�E-��X�sI=��t��F�#}�v9�G>}'�q��D��~mK/>$6Zd����-1�6=�C�ѳ�)�*�ar�ȋ�>͖D_V�ߩ��e��߸�������>&.C���<�/��#�l�"ex�8\�����pw��1��8Wv<�o�3MG{��*2/�b]wz�3p���T(=��D��>�i�Z���T)�>q��Tp�Fb���)^H�߲e��������)��� <*�&&)�m�/Ǻ�F�;w�l^>J�כ��=�>�#L_�k��/��
� '�ſY�W�܈3����!�[��kᾬ���>+�&�qtt<>�b��s��>�=�D���(�S�蛯Ǖ�[�JJ�oHW�螹������b���K�f���uG���=�Uh�|Q�=��c"f����g=�kҗ�ƏY��#���כZ=q���޹���L	�~���u����yr���`N��hY���2�[��+�C�l�W�3�X���e:J���i�_w2��	(�� �s�;���]-��P��:^�Wv-fe�V�v�ㆡ���z�h�]��xg�7K��c\��X7�+:c��,N�RBhZ��B�yv,9|��4��7��{�����{:���N�<��l֛�r�������� �S����5����2��C�0�O��ݢ�_�z+����uLó�[P���{\��x�@�o�+yNv�3�v�������~���;�E!ov�=��ѥN}E��Wp�G�5��e��`�\}���;�Q�}��}2���z��#{��|��q��G���3��%�tE+SX+ս�h�Teϳ�c|�.��j��d����^9�9��s�i�����}g�S�W�(���	����ee�y��V�+�t�v}U�O�=�+�"���(z���U�=M�Ҵ���SE��g�lm��9��o+S5U�*�wh��q>����FTL�@��+��m0�ӣþ��ZT�|:�ǧ4�v����j@�}�~��ϊ�M�ȁ�[��T�R+Ҭ���f�5(u{jf���^�.ܧ���݆�m*H�������_�F�嚏X�>Sd����)�P_[#S�;�5���3�Ѩ�:%�GK�	��c�}��u���'�K޾ <���\�����p`�c��@B���w� ���f���u�aN��Wr[]�֡����n���]�pe��z������2���J�__�ʝ7��Do>ɷY�k��7�w"7�!Fg5z�@�햞���Ni����+q˅�7��O��s\R�P���l\�.�_~��$�F�H��b���l0�󃠾�m �#ʀ�~�2G�����-���y��Y~��q���\�25�����Ba�7^71�9�_K���^5��3���VE��uy�h� }�H��>���d�G��+t����Z�A��r��2K·����Wy�����CJ�s�oA
Ĭ>��w��=��V�y��=���m0P���s���Vɾ�Ļs����E��rz��"��!q�$�ˏUv���xn#=��j���g�D�����<�t��� �F�s�';�/�HK7�ݺ�g���(����n'e���������j��j6���qmu2]f@ڌ�`T,u�=[�\$n<�\U�{��oh��;_n�@{(��F=�Џ^�{�U�gO���L\k����g�m�_���~n���u��7]}��y�V��<h�8O2�'�EV7=���L�8O�j#�B�>g��S�w����r�,�Q�3�1�K��g��q�yG�9o�S7��\�U`<�~���򎧅�.�c�,nի��=};NȬ�ݬ���[�5Y��V�o���fᐇy��V9��jeE8��(fN�xj��=.(��d��c��6�F��VmF��ݳA�9���c�5[CV]����S+�7�P�E�]�d�Z�q���]C{�c��5٤؋Vq��}�̬z=Ĥ{"�`u��b��w��}s,�5~��
�R�]{���+-��}|/�I�}=��.ڨ^��#oD�wg�����/Pe��d�7��r������ޱs����i�ް}<Ϸf+ﯺ���$S��S9���~�R5���^�'�ax���˯.9��ow�v_�dI��`,-9���j%p��J�F�<_���4��=�Ar�H����[	ƃ���O3f
ۊVD�N{�FDJӹ ��	z��z�_�<r_�o"���m<��p=������w�niI�	�=�M�=���14�m�s�=���xK>�C{5~���wX[{U~H�=.���C(P=w y׍0z*���D�C���0�=]&�����6$E�k��[��ǣ��,V����q�:�!�P����*�N��v�p��-�G+�"2��Fdb�f�r��}��L�Ǽ[��	;��2�9�V�jM�!%���"�^�$ު3=�V�ߍ��������ٿ���q`,�\{a���>�>F��n�Sf���6���1�Tom���)i+�o�iW2�]d�au���4`W����<us��c��
Z"��;�4&p	�l]�0���iu-���k�>�T�/�ki�K'�3y��+�-��؝���,aGP$mc��N�PE�Ö�ޚk�$�t�V���z$u��NB�s]�wzaz�N޶ ��
K�nO�Z�i͡�]R�z��.yϯ�����~dO\˅Ԍ���Fm{+�U'��^� �SX���7r�������8��H�{:�#dx#/��u�iB���IX��a�<��]!�[e�Ǧ�9>�tǬ�b�b�gY�|�l�r=���v�����v��y׼z�����Ḷ�t�$�nnj8
�T?'��u����[ٕ��F\':}����r9�C�ν�#�+ŭ��~[�V�|�(���D�i��T:~�G7�yk|��Յ�=�p*"��y�A�q�|�"���h�z}��W���˦\�XA�KF�~�Qrǀ�>���=슩R��Yc��l��/�Co�ُp��}��@����B�x8��ŋ����|�W�*�JB����֑%�0J<��Y���,몵��<��L[��sӹ����g���Q�Qc��Y�W������H���}MhH�t�Q��=�k��a�^~zFO�)���k���z�y��"����T_-�Has�T���8���cSG�g��e_��l� ��q�t�B��ez����T�ra������;-�qdD��6��tX�k=r�x�=�R����JC�Bݥ�>\��P��D��JFPB��o��}x���S�fS�(���0��Bh)W�B��q��	��\�7�S^6|�{� /z�
~�R��~�w�s}��,��w�M�NV�0Lby�yB����#6棻9�xz�zs�uX=�� �S�.���NR��V�j]YX�Rx8�NW��S�4�RP�Hs��8�q����Cu]-1��#�߮���[��88����60�W��;��tN�?�����+�G�s��@��aO}�:)���2Է�_�ܽɡIe1怞�q꒎��w�e{��5��5�뎦���2�fas�l&�g�H�-��V��W����碻���!g9*�9V�ץ_簌u?kK��dYD�xj�	�mHco��)g�<z���^wHhＴRv�=�G��iS�Qcv�ڎ �3=���^���P�{L�8=�nUt��l�N���낆m��%3KB��DS���ׯ�K�]��k��
�U`z�=q2�1y3��ĝX��w�>��q���U�����Q!�qW�v�הYC<l���+���:�U`y�>E�%wګ��������i����u�N���L�̖�5q���ks�c���R�����1S8�r/��.Ҧj̞���4y�,[�	�Y�T��V�kԤ�Y��<-M���K$\��u2Zv�6��4*��[1���+���/Oe`�z1+�Z����x�4��[��(�gS�@z����S���S�z] �*�eD�d
�+�k#e�_nz�x>aJ��:�p�o���Χts��W=�}�����C{�{ l���P�T�*W�a�%�����P�3���ӯ�K�壳���߇�ǩ�G>~�@������@����qd��� sٿ�MevK���ޭ�����M"G24{va{��g��G�R�V���.e��G���z	����4�\|��n��9�;Q�PFC��?�^k���N��9/(�]ܜ�`̣�{/'ّeG�h>�#�uQ��2ܑ�+L��;��e��V.ßm�_{ޱJg�)�S����H�����(=끾g(
힒�ʥ���u���ֿE��c���Y,e �6r��)1�99�9���{�	�����D�A@J�z���O\<�A��w�������r}T0]8�/�N�G��7��%�����.6V�/z�H���B���<w>��t�ó��k<�=ٻ��ԕ
�{������� %e����/Wx�)bx�v����N��<{"=TFi��!.�oV�tܬ��0��J�A�b`�:
+l��/5�����@�Mu�[G��c�e��O�Ky�4�7�98�+\�Z�P�neu]vC����:�#��Y��濃�K�[���S6!��׻G�kXĢ���ƐG���Q��C��9䞘�jp+�ա�:������Q5�bØ�z7L�N��&�qu'�`WauY���,�5�:����r�����4���%�'��j��е&$�/^�>�B�R���'f��68r�m)yX��q�]�Ұr\�9*���!�% :�۬9]i>��I�g,��irAUt�'C�sɺ.vd�����7�ط��8��yG/����Hΰk
��=voS���^��֋��_Z�Yہ�+kh��Nj]�����܉����,J�.ΊP,���5������w����b$������K��,�WLgE&��R�N���a4����Y K��aÁy��R�+g����B�hsi�w�ނUe3���WN4��q��.	�}���^wm3����Bwi�s���F�^j�Y�D�������@���ru$����GQ�uf�˶�N��B�`.[�ǻ"��-Zwt��@�]�a��� ��J���q��:�p㼷L���mfZQ%aX܌�Ay�M����!�z��ʗ+�@���Z�oB{\D.�v�}�&�tS�R���ïQ� ^%`Z���m��:4��i!�m+u��o/�A�a�΄:���K8rBn�d���L�ko:gS�p\��ei�ΣX�hS�i�@G��M���hWu:%bn���*a�&��7 ��Gu���%+��Ӽ����csAK ���.ukDi�+++F]Kh�jݦ�!���T�L,v��K�M�[ǎ�����a��{[���D�[]�3 * BJW�a{!��81���)/Së{Lb>�y���ܚ�`ͳ�'J_�mγ/�
<U�%!��p�t-��@�D���'c�ּhY'F�Fh��lf��->��s�`Ŧ�kiʷ��z��n��e�e���f����ªYZ_mVv���u3t͉�ѽ�X���Q�B

�����g!w�V��ݲ����oZ륰�\��v��U3�4%�|�x(�Ùف��-v�`�<A�_ue#�՞=|�\��-��	�p�u�f�;��m����A�����`�	��Q�٧.``b��粕���rdw>��[3�[H[�n�]�G�w�OK�z�,s�;�s0V%��X&ڳ�ް�o��I�V��Y[��yх� a�;�Kw�{T��:���4pe!S6�e l��d�qB������	r��Ƶa�p�U�E�j����(�N���iaW�+�ۖ3X����E��ˇ4�����
*#��")�������D���D���X�edX��V�**DV*�"�Em���QPV
Z+eii@�2�D�,idUV*�+q��R�U����b+mTQjQT�d��T�QW)TL�Rڍ��KX"

���A�E�X�*)P��Qb�"�Qb�W2�Z2����#m��V*��V��Ym`�H�1�FҨ�V�b��Z��c�ƋTb�F+-%q�A�(�夶�cb�1�f%
���Trщl�T*V!��U�ʶ��UF��6��-��Eb�" �1Q�mQb*����(���V1Q-��2�JTAm��*�T�jV���UEA���Ռ-W)b*1UV�T��0ʥb�Ԣ �m*���V,A��eJت
��mQF����b
��Ȋ8�Pm((
���]�����!Ag-� >�"<
�g�p�<^a���[�靫�LO
��{�N�+�����5+@^����	y'T��o��1��y+��s]}|n8��g;�s��U���f�Uk˰�2���:.�_��Q,�e˓!;�(�C�u��z�D����#�|��P�,���]�/%B��Ҫ��(���):��VEV7=�����3�_a�>C��12"t�vu��OS�/�{e~�q��G�:�w���g�������˼g�ixw�ը�>������;[�pz{ף>|'��C�{�w(0�Q��]HE ��5i�ע�ӗ]��^*���:��Õﺣ�4��qW	�F�	�]��E?_��!Mm�/A�}��;�������%E��=��|�^�mCF����:��r����A�^�R��^���դ�7�G�<'y����U�4}�H�*_d�@�\�ǳ.;�v�Ka@ ��n��x��M��:�U��ޛ�=�$
�%�p`�{qT��{��JӰ��\=��R�:��&^��
�.���?��T�t��� �[���-P��g�uo�MVѽs���U�c���8TY��L^m���W�BllhB�/3�U���ѳg1�F�͡���λ1o|�`$G�+9u��	����.�+-mc�a�Ե��b�l��pT�=�7t�E]ڬ���F�BڵyL(��ع�p^s�^������͎sM��*MH�������i:=�_�|�yK�8�{� ��@�Uy50����^?/�0_�u,-�����Xy��!ߞ��F�+�b��2|z=�@yd9���K�%��x.�3��_]�V�Nȳ���֯_B�U�<91��y��s�>#�,N����h��7BJ9u�XQ��.�ѕ�(x�g�9>x�C�����>雉.�/\{>fw��w�x���ۊŮ{}������ժ'�����$���
���^MiW>�Y��,�O Z�_�Ay�Lu��exD��2֏(����Жz�����㞩8uL�{5���ɝ��@���#�Z;a���f�Ձ�����=�G����6{�|�QFc�M��N�+>��a��t���׼
������ʿ5�ݮ����ozH�넝�N}�u�{}����G#މA_ϨS�u8�1`d��U�\6�<_��/x�y��_��-�ɟ�x�<�w�ߴ�zO��F����*�NQe�C�Mj�:�	��������x��@�2,E5p*"����f�G��t���|W�K�s���I~���/�Rv�0�V��a�J��{�;���N���S��m�#���of�x�,G&aƄ�Z;M���9��oo`�W�Z+�g����[GH�5�;��:d����GH�cŋwع����@�s7ye�S��Z�e�D��Z��D�?���t��ۗ@>Ȋ�R�_\��}���:�<���0=ëQ��)Mx��U*'٪}|h����@�RX�8%�fn*�"W������>
�t5������^M���+�|���˝�]���(�s��'��(=��LLS���%��w��ɀ����V��h����Z���!ҫ�mO�W=��G���4��q��^&����>��ؾ�wɪ>�����r��yU���<��������w�-Ux.�b���\�y{��*OO7�%���T.h;<B��M�{��N��P�Ùc�=�$�ʭ�l�9��4��C��)��N׍��DNKy���;�:X�3�X�+���ꏦ.=�*x��>��U���W3����bxӌ���{(���|^��=���u��^N��q�5LU����)q��י�7�ʻ�=ݺS��U���)��]�"N3�;P��ŋ͚�q����z+Ӱ0q���$���@�mղ�{m��87=u�#ۂp5�wO��Hë*��oԵ�y\�pW=uh�E�Ň>Dg�W�����V�:���et^}�5�a[.K^�X����:jΛ�ܡ��	j+�b:A��6�Vژ��ƞ�}��:�+&���ܛ]u�x� �&N�"�Y����=r�t�^��$Z��cg^�??I�o��f���S�w�n����p�J��Ǟ����X��RT���mE^�UFC�I���T�5�P��L���&o�Xۆ�~ӛ�~/�>�\o^�|2<��*�Y:j�-�z��Kj��[�5��U�_:��2���ϗ�9�h�~���W�K����8ѐ�ME�O/j[3^���q�w;"�ϥHn����DT\�/&P�ƪ�v:Z:)��pF�y���fɜ�C}�}r��O�������|)ٿK�g�R0���x��aSy�
�C�=뭏c�J3�`��w��4�[��k޿\xaY�q��+�T�U!
�^����?Eב�fvl0/�J�Zs���E�qaϥ"�~�@������N�o�^7 l�9��=�}�mϮ}.�%��������W���s:Ǽj!wT;u���N��<����[�rAC:���d>�ջ^-�(�,[rG��X���	+��F����E�G%e �5k��,x����F�%b�6x��$.9���n3�G��265���źނW����7s�0k៶�Lg����n�J�W��:��w��i�w��+���r�];��J�sn�ޠؤ��D?��y�5���%`�ޤ�vL'[^�@|J�pk�_ 5�c��y����<���nii%V� �]���:+���޴Pǆ��-�Vn�JY|��g��}U���j]B��I�1��лW��?��@��t7u�*���w�qײ[�>�k��^y`)������Q�;]��}�D�ԅQ�)���9�>�͉ofkH�z0�\<������xw��T%�mr�J:R��h3ﮐw��c#�Q��rw�ު+�<��'��ު(��;P���u�z��QP<�-�5hZWz+����_�M�^ Oгq�
};�{��(����p(��<{�����9ו�>l�s>"��䱗[p��T���n8��:c�N�ǫc޸�o�q�j�����ş�H�VKW�_�~z/���x��o������ʥg��)ZP��5��=����m�W���
:sD֤�����W>�E���N���X�s�,a:�dϑy2���=X�1�Y9�9��U���c5JG]���V�7=��7©����.s�b���S;� ��;5���N�~��^/H���f�/Ճ��|��uxr�m�Tmz�p��=SQ��1P*'Nr�����o'h�=��ȍ�h�_���r�O�������^�ˍ%���y���X����YY�3�����3��.�8���?k��nv �i~��@-�2"�,�ǌ�1|��\<yu90�F�s��Eh̃��B7�pu���*i��V-u�XU�b���|6�m��t�VuA-u:��V A�����msu�ڦ�ZZ�7Y�9KwG�s ���~�|��"6��W�P��cdx�<ˏA�?;�{$nvr�H��Y� �y|=�r0�������Ȓ��}�Ndl����î�x~@8my��]}��-�R�]ʒVtYc
�ydT[�r@������H��=� �V��XĽHyy�_�l��1��Ջ����1�n�ߦv"}:��3O�fH��뛨}q��bi��:φ�a�>���0�S�C��T��7��d�C��r=ҥ���Ts�?
@�ϑ͉�����a��������O��/l�aZ}W�~-P�
�T|n<�@yg�U����P�J(�|�ʪ�wO�S3�氭#�;A�^"��=ڇq�^�q��3Q�ƛ̿�T|EǺ��7�Uh�;�F������_N�O5�Nd���g�_��C�����Ǻf� �v/l{b��ܦY��=m;k�+#s�{D碚�8RS2{I��=;Le�MiX|'됝z#L���bl�0��Q�L��6C��'٪x7\�����v��x'��z��ՕLed֖.2g|o\����>�p�m��I��Dx�U�ɚwu��ܺ|PӇ(�=�\�j�S�[�P���Sܱ��\���2�l�m��bȷu:(�1!���^�4ڷ8��oF�&;�v�wʯb���n*��J�YǞ���
��u��'�K�2���W��+*���շ��5�p���'[�,�j� ���O��toG���-��\c�M��'ӺJʨ����ѩ������x�K�w�O�ɝ�R�^·μ�z�Ü�p����H,}L�:��;�&��8{|.�ZT�>��T?F~7�,/�yP��}����~� ��,r���>Ӱ�r,���zw˷U��Y���9Q�&���'-l�h�W{�)��|{�F��˹>sQ����@�^O$g�}����,��G���늩Q.�,yg�,*�����6c����ۇgoó�/#X7؏�ޑ������ez�tKf�0P{2Bș^+ex���nLUِyg���Q\�c�l��zQsq���c��+��G/�b|͘(=��LLS����Mպ���j���n��N��@���=4�|�k��z��ِE}n�n�
�4{>��S$@��K�߫g�T�DѰ�c0�Gy�ǜ���~g>>� z� ~��z��>:߉�\�x���!������o6�u~��Z^�Q����r�P��~�f��t�ȗUc��?
҃4��ԕ<Vh~-`�E$�-�w	�f[�3>?
��.��J��s2Ğ�A�f�����K��p��.�c��?JV��%�r�;�5�s/�ת��q�i�1���d��sqի��u|q����f�)ծπ;��z���"rX�ͭ�'|f�X�3_}��r��{�$�ϦrɆCU�fo�3ۛ�/5����j����������*���p������z�~���}vJ��6�y�ߖ�vw�k�Y>�*}�4+c��:b��{MǪJ;q;P��ŋ�UhP�C6����h�L��� �L��ڴ@����ǹ�'��4c���ǂ{MϤaK>���ufǻ֧�y�Z��[�F�Vw��uH���v|��{����^wHh�-��ݢ�=�a��v/Ӽ��c7Ƽ��e�T?d��o�&n#�\�p��1�rq���s\\�.0�a'U�g{׊�8ٌ���@R�A�L�}�y2���ϗ�>�4��^ӑ���f��D��͘��S,8G���mF{�l����L�rٛN�(��2ej����~�������T��l{�l�h�yO�ܿTz�
��N��.�O*�a-�2ԯM����xN�����o`}�C�ΐa�ΘqBR=��3�����W��P6Ksq��$!�����>r5�y�{�������?�+J9�/��z��,`�b&������m� _f�ِ�mc9���/4�gD%7V�{Bz����ԫ	[[E�P��9�|su�u���c
,`uλs(�u�*ż9�/�Dgr%���O��R+��+�bs{+sk����֏�R>͘i}u�Xs�H�l�+Ѿ����^����P�I�|�쇻�N?2yS4�c#�]��9�P["eϽ9���;�מlt�$kv�F{,�{@Z�%͛�WoA��^@>��6X��n;lM��
��$�}��q����l�O{�%ws�F�4�)��K*�ОX���d�@�;�M�g��U��"�\�@b�����w��jY9�r[��+Nzʘ�N����r��Χ�U��#��o���2|:MDk�y	\�(��sr�����py�Y�F}� ��G��~�,�+�	Xo�>.��\en�z�vL�Ѵ3��OP�����zx��`	�+��ds�>"������BEG�
C���#�E�Q�����o���.�^mV��g��~Yn�KӾ!G���{r�W��hq���5�Jt�뵅g�~0�J��g����z|}�5� ·�U\�ٝn�x��t9��^@"�h�Q����Cj��թ
e��ɭ/	�Lc#���#�5��>@�9��ݩ��φL!�[��.c�1��s%��|��
O3�f�0�VE�mɍ��|�u�0'��{u�w�t�M�Uw<��Ԏ�t!n�B��ai�n`퀗�:���ha���Kv��}�9"�U�wN���˳��ʻ�@т�<�N����L~X�?~�W�v��F���-�98
��:�X��gY���.������؃�n�Of�'���	|m���u>���F߷й�FlCȪf�N2�f�ȩ�@�k}��P#.��3�ڼS�+�n�N��W��xX��?^��p�#��^q/-1N�q��+�n��j��Z�����SZ��:Y�g��n�辟x��چ�}��x��Aܯ�t	�޿[ӴQ���MG����=x���x�Ϻe �r���N�8Z>ŵ�|�֑ȇ�(�r7�:3����y��%O���F]o�r����f���v�dL>��XZs>�~5��T;��g��o�V��oxmn�����(��L���DM~�r@��O�n�U"g�s�:3��Zw 1��z�\z�
�ǝJo���;��zv��r'Ӱ��e��s^���웨{��c~��h����r��ݫ�§Π2�����=�����R�b�r<�@�Ǎ�O|i�uU�+&�ݔ�BY�"���tu=�*0��I��������1|ꏍ�΀�Ϝ��$�^�(��Eh������xM��#zju�$d�a����*�p3��y�ߜ���l
[��Mλc׉�w)v��XH���v�����K}�2R׼7���`.�櫫�L���I&��^�,�Z�Az�!��c-�z[��mҹr��K tb<f
Zf�!�]� z�)uf��mV��אiw(wr�ֽ0θ;m� �Q�>9���H�AQvuq������G�աi�y����c�g��P��r���igW���#���V��n�3:��&N�AwhR�jT�
��Yx��a\s��;��|���3b�]c��*��!B�nY�G��I"��/zB�Q;�� LF�*E��QO�Z1�s3G�.P�|u�S{�/�L��p8λW �]!�1�w�D��q-y�����mY���g+���whN_%�K��gIs+y�k.3C� ���7���ߔFq}������6� �m��f�78��l�����a��v��Jv����U�-�9�l�D�e9��9;vM���Wf��2�1W��`>A��;�3+���p�u�F�묁��<���y;-�WK*�tQ�lP�:�%ڡN�J�ɽ|MmP�9h����L�{�!e�.��2�s���9�c�-�r��+n�gE;�G/+A=k�`z�Ų�l�&��Z�+�ћ,��4R���:L�R"#�*N��o��ʛ�e�����0qE/T�h*�аq�.�`�K�Vڒ���j��99�T�-����[K뻵d��2��J�#��ו�kM��,���P�8fz�D�g[�����_Vu"�K�Z��Ќ�ݏ�x�ntxPks�coH>cSP��}(4ps����Y9�9�3�b��f�1]�&[�N��)U�Z�X�+R���k�-�ն��`v���#Kpm0���Aj��*�n����9�n�q�-���%�q!"��0q�&�V�W��(��ںPe�Oqa��Ѽtn�T�TU��:')�3���ͫL��Eb�I���jэ�T-�jG��e��v�0����4�͑U㙜)��t%�:{���X�����M����G �
VE^����K�����T)��D�l�o�kü8�p�ݙ�)D0m`Un�{lp�iq�"�ϸ��]�ot��	[!#)Sђ�����#8����X�Ur��5oq�c7���f�]laӣ+ǔQ�ض
h�*��'�6p�G���m�w��9G��]nLJԖ����_�B��>�#2�4�C���N� mE[��!�kz��b
��Fb۰���A7�"'�C��0'b�EKU�,C��ɝY��NbQ�ۥ;p*�]���M�Ȳ���%J4v2��}�:Yopf�7]\��rf������u�<�,��܅,M�t����=��G[f�;�|)U��\����=M�t@\��w9�-`�]������c��BF���.�G�����0;��\�fvcy՝{N�򻩝:��rV���07�u�G���|u� �u�Os���>ˡ6�q�kz{k���.�c{ls�Ɔ�ݽy��{E��DKh(" ��"2+m���PՊ�%J ��Ŋ��+X��j*(����X�DEb
�U`�Z""*e�Ub,�(�6�EB�EFD��2�U�A�"�J�b���V@\j�2�"Ԯ!PZ�Q���X��%��#Pm,��D�b��1Qb�`�"
"Q��YEQ��ŊĹa��DV�*
ȫ嘨6�*TUcD��TV[
ՋUH���#+[l1�Qĵ��Q��1dDX3-F� �Z�b�11TU���VQ���-)"�Ub$X�Fܡ�J*,q���e*��Ɉ�(�a[J�����-�K��,)l��AAaKJ��b�[(����U����Ģ+�QDc�U�(Ո*����[J2�!�eH��A�`�� �q1�(�*Ŋ1��s%�ER��R�g1\/T[�c��9����V�Z#�~��q�\��>�x��7��"9��X�� 鈌�t��[,"����GG����~C��{^)�A/�z6���y�����g���|*2��n8����w���a�	<p��v|2�Ӂ�\�tޖ=�7���Ǜ3� ^�j*�Ǜ�wmU�u'6}�ݸ�<��a�'�EǨJs��a�+�|+N�3��Ł�����4]��JR�Եw�V�X��nyDsUq��d��=꓅,��c0Ζ7��>p���j���W�
���G���mH{q�� �������g�8^�x��� 4��2fyxO����t����^�Mt��g�{#�Cpׯ�w�|���z�^��;�Jq��Z���.J�����/ ��>�1�&a��^L�L��s�T;��r#�+Ū�xpP���`�K�=��\_�W�p����)���Ȱ:)��Q>N^F���^Wq�#o���;��\���q��#�z�y�G�QU�^���ٯK�Ȋ�_K�D\��}��¯��C=�ك)�3~{'MH�Ќ�g�1﹇I��z/��|=��,g�D�l�A��HU2�V.W�L�ê�330O����B�䞓�׹��l;PM�'_�������i]\ΗS�b�
�EpX^j����;�=C��+.�m]�#��pA���jAW!�q���d�X�eKΊ�M�q�t�f	ݠ5���C����;��)������[g[���c�f��Ke�)���t@3^ҙĹ�~�:�w�v�X�t������ ����P� ��0x=���LL��eO�z�1�(�b����@�J{����s�;^dG�|��=�T[��*���	��r�֟����0:��}[��7��3����^��G��0l �=�`
LoF�wy3�^��N4��UL>�8��6��}~��Z^�Q�/MG+㟬ٿy�GU׽ԕe@�}�oO(�Ox{(�E���>�������3k�k�4��cܮ���g1��z����>���0�DΗ��C���q��Yzr#�O�Ȟ�ï't��'Ei�s����J��E;���5ܽ��}�{��{!u����vՊ�~�:b��'��z����.2�Ł�����p}ޒ���{8��] o��1j��K�~<�G^�/�G����;�O�a����Ǵ�z�=P�We��%|�*=c��{�]�H�ہ���o�iG�������yh�=·L�SR2W���
ea�/ުѧ�(�n*�{�d��pzet�׫�V�_��]Fi�+,����񚼀䈫�QqwS��m��R���-FКM	e��Ҝ�7��L�ٓj��A�!P���,is���8� ��j���ywh�)�ը��9�,gaᇷ��p`淳��]B�֮���j���:�7^��k��W����R�K��\Ov-Wpj���<�jg�=���ϣ�@S�5����~����S�����2���2���WS���q�Q7��l�_JU}���IʇN�}�U�MO"*�ȱq�(x��̤}�Ʊn�w��kc|�xd��FC��\sޟq.�Q�����g�����"��L�~T��������~ȭ�in2ܻ�_�\���}��`�����zᎃ��z0��=�mLqS������/WV+�`c�Oun%��#j�����ԑ�~�@�����n�\G�^7���tb�6�Uh_�� �>��Ш��g	��\��y�~�~s���^���.\�O/fS�{�.|@���#�!�*�J��{Nl@-���8��*C{�1��\���KF�uX������I����<�*�פ�UD4{&鍸�Q��V��kòc"�6V���Ы�}��j���ޥ71BT�2�z��e�p�}%ѿ���V}9P��oC��|:H��׶��&�}���^ZUW,�z�2�u�z��9��G{΄��y���A����z����n����尼��yy�+�r�ג��(1����}��5{A��(�R��R�ML���Z7�
hs�ʥ�M��k-q� �s�d��;{��WP��Yv1\{�v��}�o�V�V�`9{����뮭y)X$}C+��픠W�7����g��P!@��U}��	�Rܘ~n����x�� J�^Ψ���%n�ȇ�ECBP~bO�%�z��uR�]�����70��1�C͙ú}��u0��v�^��R��_G�v�T�vS�V|í�Z\�h<Ǣ5�{=TFi���c2v�td�\ޖ�n'��6��@M'Y��|�G�	�z���g�v|�g�-<�E�:pzzp�U1�gK��&w��'7�G�o�'s#½�'2�q�˝�{+s}��1Seq�d����vym�m��-�98
��:.{ŋ���AF�Y�E�� �����]�f,^�9�s!W�z�>�>Gr=��nZ����x�(�(�g"M����{��T�gwjk}[�Ʈ��g�=�Z73��K��<�z2=�|�?O��u��C��~��v��P�ߣ���߾���?RtE�W��چ�_����"�3����E?_�����%^�oеqT��2�6w���s,t�Rݠo%��϶��W�P��^��|�%������N8��9q/�c�=�nE�:�E��6`�v�d}��Xml���ꇕ�uD�ˊ�?4��-��n�6�t}����t�t��C�5�Rsk�l�Z�o>�I�.�}^���n�v��ļ��X~��璦d��iߦ7���+��F�
�p��Z�K]���Ss��+,��aU�;�r8�����k�g7�fl����5'nR�����.>��D���z�>ͺ�ne�~^�DlU"i����Ҵ��\u.�������p��a��C�zz�1�s�L��t�e���u�@�T%��un2�Lgez���� ���vz�����G��t؎Ud�m���y��J�8� z� ��@�Uy�r�^	�ܪ�JBۼ@8oޭ��='�O�����E}ذ[�Q�9�fd_��V��^��S��O��+�
<tע]1݆p=7�Q����/��ڇ���xo:��/�LO��WLX��[27j�K��^r0�`�De7�$��d��ge���8���K雎,	Y��S����W�������|�e��@��ΥՕp��t�y�'p�@���?�����Vy����M;ǵ��|�v=��c���9�w�z�����n=�g�\y���&�.�c+&���7���$K�]��VU��=����7�R�g[ T.�~G���C���=�J0��M��Jb����h��c��s>N�ɝ�e���5���u�{}����!�}���wqEMCp~��7�7z�~lXM����]��AY�/���N��\��}O��y�=��V�Gyu:s;�E�$YY���R��1n��h�u|Q��yr��JN���ټ����6m��;���)�VK�j�`wj�OE��_N����D�<�$���y����zs��&+�q���p��I��t���5������z7@�4�/����+��
�*�^9]9�s�G ����S-F������9H��8�/���c����X��un �ۜ��q�@6n=.�}�UHʉt���<��#e�ޣꦢj&+ʯ7�;���$��񍂵Zgc�a�~�d8���#�Z7o�
�W���k��	��Y�N�:��,���A�_Wq��P��\��F{2�,�.��7
W�Yj�g���ݙzl)�J���J%�Аs�y~e���[�Ƹq�pD���p6�7�u�b��<��ؾ=CK7��T�}2x��LW�v�㺄��Q�¼.=�W�<�r��������++޹��w��zTi��yY�Rr�cn#6�u~��_iz}F�e�	�\�fϻ��4u߲b�.�5����-]����C�����n�9�NO���ѓ�3[/I�_ic����8i�����ܦ�}Y�ޅ��TT���T�z�G��6oߤ���ߪx�OW�כZ=-`xl��ndIu�~�o����/-[}j�!ˋr��C�ݶ�B�:q�.6L��u�{��;A���=��]�^W@3�����N���}�7}Ưxv=�����ce�݄v�+h�1r��j�)��ͻ�}�z�*P���r^�Qp��٧�۝����)����o��Rk�=��9�힕/ݵb�=�.�
\r$�;q;P���&g�窰��.�t(�J|���g2/GW��Ul�i{o�g�U���^;��i�����*���Uc�`����st>ng���v}��==G�����y����'{⫣Ԃ��v�	T�{Ww �c�k��ԭ�^��=c�k�(���L�1Db��q�;鸌>�����cm�_���_���4p�RQ��2������kh��P��!�``���&�����Nb�}K���W<f�B�},<�0qFZy�J����h��t�3y�,��Q�ç@>Ȫ�&��|����S���`�^�e�����)z�Y�-G�����˿\z�
��u���zU �*�f��pʐ#qq?3G܃&\gWpva_N�yڗ/�_K��8N�U��a��iup�Ink��Փ,N�Q>���@�2B���@�>��T,���M����=`h�v�F׽��;�~>Lk���a��t�7��� ^ɔd��. ���	��_.�p��9��Tl�m�{�\�x*㬭p���b �ܮkOv��n��\� ����eʉ�$����[wb���DH�TŕN3��w^�.�O2bvg5%��S;���̣�����]�tG�v��r���;:<��n��s��gYS�d����o)�V8×5K��@p.J��:��X��ne��'Gŋ0|2�j��s�TO0H����u�h����
j�2��]���|���u�mH
��,
�u�"�Q5,e�H򋕦EDk����������q��8�;lT+�������t<��p=�3tםx����;ӕo+t��Vi���s�3����J��E5n]�߀�I��Fo��>�����ՐD�+���u�{�')�q<9m,���f���L;ͯq���<�� LBW��Ϲ�~�rz��"���H�O����\
��,[�ɖ���+� �Tv�v��C�zx� l-�`Z��W�H�\�C�[��9FPŚ�3�C�7�|1�;p��nvX̝�]��gC=:=s�*�؏p̃e+���^��3W~o���gk��q��v�+��m�7��sյ���r��9��<��z����X��>N�{�i�h������{��<�J+�%��+VF��[�����6����}3^�if���yi��3��>��
��g��s�uǲ����q��Q�_{����S�����h2|G���N˻l�:�R0�X�H�Ze�p61s7b\��)7���!�]\Q<�u�C9Ҷ�di�t:�s�*��F��v�y�����q�(P{�ӄ�۽��zWJ���QŜ��#}�s�Fr�a�i��L.蕲�sz	��Ƴ$��/0=i�V����iL�&X^Χ����ף"<��2�ʼ:��H1j}���Dؔ=���Wo6�R8����^�*ԯY�mCF���t�ϟ	�]��B�emS��q9�O�U��k��5��g���6O�ߦP�E����h�s�h�_uC��z�-� �m���
6o��5��Q�[�:=oף��KC$����ͩ�0\����͗㵌�lH�DO&;<�{R�ު��eʤϽ3�J9�H����Yn�����7��TFE9��ݐ�y�ڽ�fs�ls�����i�ٕ^����?L�N ��܃o�FH��x���[�I7�g_�ZKB[W-��ݭ�z��{ �Ud�m���y��J�8�z� �;�c�=�qj�`�Q���.D�Y~������0���p<>�^+��c�������C���q��D{�ʶ�k��QZ/�n�:o�*�]�g�y�P�3k�o��f�ڇ�P�e�g:��/*2���={{�}}�ѻ�&Ͼ���<�(ٸhIG/�D-7;,g���s��q�����]ʪ�G�碹{Q>n�,B��ы���ʳ�:��*u����cBi�2�dޡ��lտĦ�j>�"G��b�U)��K���F��G��xG7���1`�����%v�Ob�
���+a̴��v�
;7Sc;:���9�S)wa��T�[��x� xXF�e����=.!�נ�F��'� �H�*)?�[x:Z�ǜk�w�P3��<?�t��0xON{����私؏z������FD~��{ Y�-ʫwւh	�t�J�W��癑�)�����uH��Fu�|�W��}�ï�z���֣��g�����h�~�{���̝S^xK�T<5�u׆�6O�7	]r��N��q�:�]�����9Nb�뛿c��0z�z9P�O��nz"j0	��ø�2�}nX^9���^��+�p��=�]��
�#ιI��ˁ�B�������"�����87P3�'/#f�F{�P�#���~�uO�{�b�s�Ͼ&��9/MDK�~�eF/�K�dUHʉt���X�>o��U��c�]3FϠ�ƬG��v�м��lǐS̽�7�u���%��:%� py�Re�Ï`����^F�g�꺶�׊8�G��,w���ۻ^,?t���l΍Y�+��B�����A�2瞸1�zEU��Su��*g���ON���zwK
L��r�=���]o���BI� B��BI�@!I,��� �!$��!I?���� �!$���$��BI��!I?`BO��$�BI� �!$�@!I? �$��!	'�BI� �!$� �$��!I?��
�2��yS����������>��������I
�
�I*����L�*T��RV���B� ^MT�P�AJT��UT�R���%`x�!�����A�Ҳ�YT�i\u�T�ny ��!��k,�
�����1��makSZ�kV�wn�*%R�(s�sw��4����  �h��wb��*�,H��+vk�]�(w`�ж�4W;:wt�5D*�*�7k*��d�V����f��RQ ���:�U�d���I��@�� �����KKS`ɛ"��]�֕�[m�kj�&��ٰ-��k�mCf��lXԥJ����� 
 h�ʕ)�`4@�FS�	)J�0CF�dɣd��&d`bba0�!�&�O��R��42` �4ѦL"P!4& M�ѣD���G���z5<ԂS� IR�SL��L0!�`CGOI��ˌ�鵺o1~�� �9�  q?X4E�
��@�#�J*  YS}����~o���Xs�vA1�*�����Q XT�X�"6� ��ߎ4��,3��w>v��*��Q;�R��N�$6����@���Q�С	+�ݻq����V�W)���Eu�T�c���[�KCjZ7a��]�B�SS+oRJ�,���z�|n�=[@aˑث���^�6����aYh�1z�b]�Id��͠�m�5�&�-Z�Yk��2��t1��>�����b<����՘^�s�u�^�H�>&j�n]l�m"@j�j�nPTf���b��M�˛`�h
�jݗ��c���K�[��:P�M�F�6�B/*��Ùe���A��)D�(�[�:�Ҥ�qf�/�t���Q�I|�`��ϯ) ��Ĳ�M(��闹ombښ�g�f%E���`�B�w�!�b�G�r�â� KӦ�5j�Fc�l�m ��ʕ�J����,�aE�G1� Օ�����B�/3;N�0�����e�mˀ�*�f��w2�+�frKчV2����v�؍�B��uZoaP�ZCB�Om�-� z���KC.D����Q�J�̨�,���"�f���XLn4J�KU���ͧB
��d�g%�L�L�(l�Q�r�։.��[�Ȳ9x)�Ű�&[��k��Swv&�cIc%τT�0Q�K�٠i!�J��k!��SD��d%�:g�Rg�w1F�-����.¹>��1;5+�Y�M�.�P�l�ճ[��)!1�o���m^b)�)YC#;�����h��n��\T7UH��"u�#�U�mK����V�QY{f�����*ū5xK�U3,�@f�Z1C��B��7B#S��
����������)o�Fy��]�Y�t�!��& H�!;����-M8�mL�h�0�*�ФElw�^ �1�-�н��G���Z5|�3*C�ݙ��3@��OI�@k�]�Tۻ�[�T�6���F2�A�A������Z� �5#�g6e��^� R?��ZF�]��L֬ȋ�-���9�1h���Oe3q9���gJ/	�^Ej�a^5����{` �SIHe����7�Gv�R���O9Wf`7�*(\l@��e�m���T�M���Fl�ѠF՛�A�l���̱&U�n�ث޸t��	�5-�Y(� *E�=;��o�f��9n�����R�1�:.�QF�'%�+��I�E`�'�uL�nC��,T#-ҭJ+k7�ֲ��9x�9 ���*�Xa��K̚Ӭ�Z%�B��Dn�Ra�.��f�ww �M�k�Z��
�a�opĲЧ+^*����$��<(²y��O]KQ+u�P9�����"��:����҉��$�/qH-X����9��e*AȰ�(3�n�F�S��F��yy����t��):�ц��ELn�F����[��C4�	1H�ɔ��;�Z�P���w5Ƈ�Ù,f�ԷH�@���[B�l1Zޱf������lu�,[a�����Vi%g1��+6�X��^'����Ѳ�Gji�x�
E�Ǹ�D��#V��v-H�f�������o	l�����1�kkh�)�&it#GB��2����Lgİ�kh�B�Rie�:�:�ĩV̆$1SDEK-�L�e<�p�eJ"�
K5����9i7�nYgJZp����VS�6�%C~���Y�+>e��<�on��o@4^Sz�R��*��GJ���]�Q��r�j�'wui1�CE,�F����-E�yY��*� 'sV�C��H�ԕ�m�<^�B�Yg,�l[�H�;T���奺��ь�YzԀ����Ѝlu������Aa|i�՘(�2_I�s���~�_�C����[��!ֶ $?/��S�"�?�ᱳ���W�����_�yǞ��Rיq���P��|�k���*��ZqĶFs6����p.��4�j��tT9�Ųg*(�V�C��ga��h�/n�W�۸�)�7Oٝ�0CQ��P�cy�-�T���낁gnW.H�b䩑j�i��2�-���M�WE{��_J޼�9�V���btor����8��;.F3N��*=��2+w�g���jhRd-�ۀۜ�j٠r�2�ŵ2*J�!�mWG��]ligv���v���9:�sȣΑ�RQ�4���l34�kD��c��3Sz�t���y��u��!�����=�	ng=�r��)ʊ��}gx�܁9J��e��y��Rg,��V�Z���&KyE�f����vh$Ê�]Z6����c<�^��5�*����X��Y� �f��i:'��aK��T�}�^�� 	��+���v��\H��,96�H�|	V���uaT���Ν���p乽�r��/9��{�7ë* ����+�:mg6sy��S����B�v����剧T�ܹs���ð�b-I�ҭ�So1P�}m����%��їc.PU�X��T��Η��8�ڻ�U�!�
��j�7�0ou�ua���m�f��S&f��B;��藄E����N�ۭ��|�mMRc]�&���v�嵣���T�꼼IP��*	�o�d��q<�7,)��]���9Lñ��N����ʫ�٬*s4����-�d%u�"{5�f�Lth+M�tqq���V��e�|�m�ʺ��<fv!#si(�2�u����wq���8���R�'��MkfUD ���	j�\f�sw3�*�9Yz�j2A՘�V^W_f���uj�����&8>J�ŴR�$���u���1�W^�[�g�/v�Q���G5�>����;�(��w[J�V���FN���t�J�j�f�s3��kIZ����[�\�Ӈ�rz���_۶��Qph�=�J�z�!�7���[���tYF>��!34�a�q��^�3F��V���@�%�XڏK/���ď�e����I&�f�9�&@����ֲUn�X��a`�ӥ��Yn�-�@�/6��2.�k�]�$�"'K���]B��0��x]�xe3sn�R�l Z�6сh�9U.�9��&��b����\x��ԚxGv�pLGo����Z3���ۺ���j3�(�8��"���&�:���ى��]�B�ɶ�����f�βL�3�죆�B��R�:�{eu՜oBlˮ���|ԭ����r����ܭO�r�F�c�rj�^j���4���2�(�T�$z�<���Q���ך՞��<�<7tU�ѺN+�WÀ�I��u�\Q���7�$���TP���	��[���G�ēs�xm��Oo��(vt�'�|Oq���):����py�[I�)M��26�W��k�S��p���*�w�Ⱥ�>d�2��z�],WGq��+�;:�Rgr��|�8�����"�%׌�¯�]��s�%A}YdĻGL&�;u�9�śܐƦ�����;�@{z�Ny}����ȡx��x���s�j�ΔU*Ն�pPx/,7]v¢B���4���In�v{*�]�h��>E)]�yz�7ZtU.��7�+J5��yc���;�7;��e������7fΜ�ŒXK髷:�|�U�Q���P���z:4K�l����:�'oML-C��ݴ�fB���C���S@�'Q��]�Bkn-��P������ Ӝ�]����]ԥ�Ʒrn���}�n�* W3w���.�wʐv�����_�+�m4�Z�n���P  �$3�r���΢)�mM��ꪪ���:�6���?ɥ�E��J�b��kj�rﲦ�H7���b��+]
e��9Z=q���6��3&(�=�
 �
mq��uڐ3�*ET��*.�;�k=��e�Q��-޾�����u�������}�>T�Y�P��%u��^�<Gn^b�o �G����s���r�K�y��P����]�ϑ��U�&�+�Eۼ�Wq)M��9w+V"��%3��J�	.U��b�.7D��|̨���pii�}[ȥ|�_hd�N��Ι1���R�ttH�n[�`���+XԀ�[��͕
�(�Ndv6�Ő�r�%�PY���Ej���ֲv$z��Nys�:��S@m%}�+(0F�4w �����Q���qc�r����Y��-����S�u���rϯd���m޶�|jb���p���6�:�oi��޼+O�0ʣ{}aNl9����1˥Ih
�d��5�$b̢º�#;rXWS�=p�cw���M�u*�3�#�f}@��J�ᵥ�2���Ծ�\�&�������sU��V�U�U�w.A;3/�Cbo>�WK�E�R�x����
e**��Ұ�>��٣�p������=�ahSg^��P��p�mޠ��t�-pK${�X��G+t��g�;u+�iw�ݒX9!�87�'`�3K�Sջ��7XB��JdY}�a���VGKd7�X&������bN=�L�a)w!ל.����c��`a���;�шDo@ďb���c��(dvI�߇ۢ
4�a��{��h��q��ݾsC���,T�uѵoT�����cǡ�֓�A�o�hQ�gZ[�f����9�a ���b�:AWn�>t�r��
s�ژ@}�U!u��ήv�|��w3�bt������7��3��C�=Wt�ƭ�Wk9�23]�i�MXȅv9mv���;�d�"&JܶI-��V-��ۍݓ��^�,���H�H����<�zFL�򂘊у���nU�!�3�M��jKhۻˁc�Q�X��jX���b�k����K`�N�zӼ��%�_�dp�t�u'h�˭�ovAb�����p4v����lQ7Ci. �q�/����P�I��\�?��{�t5�w`
�-�����<��	��_t��bJ�n�սO����na���;�u��0P�u�ε�>Ƙ�z*n�O&V�^���t���C�ԁ]j��J�����F��{���O��^T����jY��g8h%�CǎG ��۽���D��.�u�6�=�xVu���el�L�e�Y����9nn��WHr��Ƨe�\p���<hL+�7�g�L=�
A��i'�m���]mMn�U���;лe`����5q�D��{��л��-kZ;!�A���H:��>�xj�#�lCY�)�����!,�d��ޚK�!f6,>���kn�^�6��wo,�W�1�R�"�K+N P㯧Fwmmn 㥧5Y	ʘr��[�,L��(V�b\��뗬�2��+kt��Mo@��2������J���6��8��z)�x�ц��������O���t޳K ��/I��7�E�ợ�P�z�c����Z�Xښu\G�xjo"��V+>��}5fW�fl`1ڨ�<U�� �C��vCg���IL�(W4|�^ms%sls��a^��Έou�����G�X�y������U�wS�K�y��S����+�vу��q��?���w�;�����%����U�N��hd����Q̂���E�ZXMw7�0E0�
�f��
��H��4J�p
l����F���ٽ�����0���o�e�O����g{�'��ˁY1�5Ջr��T�1`�����|�RS�]���#����m��vkO��W4q�C0K��xDL�Gw�b/��]�9w��S�_S�E9f(�gru�{B:+��3�ș[�̊��˲		S�-�U2󀗛����V���gpDz�\Ea��1p}X�bW��V%�%�W��:)0�x�N����3)�7ܺ����&���Ǐ�����bz�D��r#J�#Eȭ)$pcH��lU�����v#Q *(5�����V�Y#D�dH"��cQ��DEZ�F�QQ�H˒�-����JDnKcd!r$H(���E��z���讝��BJ�Kkmwp���_���	 L=���kJ���U�bۉ�pl��W+���`7���,���k'���3A�p�U��{�V�(`��ܺ���U.�.0�9�i�l�5V.�у��ߜ]1�4�4�YZ>�NF�t��1���:9�ڥ(_d4�.PJ�!�uה�W����H�� �η�v��8�f�ˡ|�y�1S�ëG6��
ۼ�n⧙þ�j��,k7�p�u@�d��c1�ݬJR�����������5�4y�4�� *z����1_	cb�ո&���毓^]J�\l���l�[�RdG$B����nD�1嗛K��~�� Br�@.���1��[^Cj`�HgFIa)�ˬ��_��.=5���b�Ҽ�\Xe;��f\�;��j���������5Z�\y�o:��z�����W���)���{�b�c:�&��PLW�׽�;�eJ�A�nJ�xr.��7m�ܪ:H���:.��+��*n�Dč8-�7��T�v���_v�,ڎNv�6�ն瘎���ç��x���s=�S�#ZKi�k;ZnI;�Z<�Nv`�)ū��l����5��{H�o��2����w�@���oT�h�V�SV�;�\;���rț�kv���+�)���"�4�v�#)�ח���x��D]�����N���:I��^ڵ�w^�C���K�㋝����G�p8�/��R^�W�����{f�|����r�N�C-��ܪ���y��u�=ѓ�!Ȍ�,	}���X�JK�@�zm �T���c����v�qc��Z5
ܗ(x\���{������>��5{w�������'\��r����ռ侚ңM�F���u�) �S�Yӎg4���`��М¬?7�n7��r�<�{9q8��׋EEcŜ18)OMڃ<;+*.�>.�����g�G�:���I����]�u�\Oh^�WR��'�w�t���;s�F[viXъ�tjnd4�&:^�F�w��1^���M�Dv�����Tc��+��+�,�KF�퍞�v6���=�8[�� ��w���B$��+ö�W�妲Y�Qqg��P�h{2�흏��j�ھ٥�4�{K<c�	�hGI�A`�اk3x�tw��9�"���ٕ��N��.`��m� ���G>�-�c��Ots���ԏy���41O�� ��RaUo]���Q*n^B������fxL��%׿m��B���y�S�%�P��7�|/>�x�DV�̬��wεD�d8�C$e�G�U���\�����%��MS�.��纰��(
�z���и��t>=���_�z�~zʰp[{z��5=�o��E�B�;K:��VF 7�]9m��Eaz55�f9d�]����*Er�F}J���G�B��UF����O�j{?g�����hU�i��۸��l#P��њxʕ/(���Yi�j��Ԧ�G�e=�Hm�ӋB
�ZV���ha�n�rJ�h���m���9'�<]���X����Q�os�I�t��p���R�s5${)�o���C�3G&M�iV+%Y�z!��x``r�Cz�ɜou���&
�V��f�ӗ+"	����63��k�������2^T���HUE�998�2�)&l|F`�E���qJs*��wWL@ 9X��t\�X�cJ�Y�5����[{J��@��C�m�x&�M+YQX,�o�E�x�r`x�Z+Õ�9���,�1I�V� ��к�f�=mm�(�$�����B�L��x�������ɷz���&��܎#M5�+�ʃ"�
2
A�bū.5l]�1��R�id������RB�����-�}%�#��\XSP�q�DRd-1�J�8+Xd�#Eb�)P"@�ϛ���.P�&�0v���W`��T�Z�5GU`H��!w+��T�O��+g���Џԝr�[���+�M��6]a���&~!��2�e㇑��LhW�:�nu��7��9�T�^��ij��u唡�wQw����S ����ri�rf-m:����#�Mѻ]�OV�2�_J䢷�$����(�W�T�ee�c����U�dӿi���+��j��0#���='s�Sd�������0{#�;��������YfQ}�Y:S�ʠ<Z��{r��_��]Y����YW�9.�ѵßt#��G�g�z�9��1u"6���o�������v-JX��Ѿ���堵�C;W303��t�Z�.���ger�;ػ�(�N�������X+�x�r7��ƭ��Q�O�/yI�V�[�
�}	���h�g�� �`�[���9�n�]���.��6�oF�W?c������� �EX�P�QF��~��p�K�>�iA��W��AQ5M`��6���҈����Y�\��L��g�@DLEL�D� ��Ч��ڠ���֩j��q���U�A��m2UQ;*��m*�g������ �-W����F���@�5A���%U�s�I�۪�hWZ��n�+MyҫM�h���	���1��J��k�AƏ��5�(�A���]J6�����}��T
UV�+��+�Q���G�BУ�\B��%Ҫ�j��ߙ��ꈔZB�Zr@�*�MR��Z��T|�h�UY��yϹ�J��1�4%F�j��e%�R�ƨ�(?4~��}�������t��I����f� ����g8��i�:n��O{��{߭*�jG抍QF!V�T[EJ��F҃�����~��GP����x��J�xh�b��Z�k�=�>��q(;�G���h8�u�pY�*g�)H*Z�g?k���*�j��
<�T�W�4VnU!Vs�U��ܪ�(��g�~��k�Tq��E ~h1
8����iA{�Uh�Ur����J�?O��}�+�%ওH�D\@LA/�EZ�o-�1�5�:�K`SH!X�X���j�(�T�����L�_%Q�߽���U�A�%UP�#_%bUV��*��*��j�j���%h���K�wuT9(�HߥPy�Эwg�C?J�??΅���_�#ֿ�\���J�_�D��EeZ�U��@�BN���)-8�6��	��LZ̛�/����X!�L�'������r�X~e�* ��KÒ�6�'L��%v졑�z;Wnf��8�ή��b�)��ݻ�b+N����7Q)=��~O�#�Ta�wY��C#�j	�슝SY���֒�Jj�Qެ-�;K���
�����ں�'*�R��Y����K�[�5�EI<�}�{}q0�9
ϺXŢ,f�\m�TYY�����[�4�������b���iO����ZVu�%�ƏI)j�t���Q�^�<��뱵u�,� 7!��\3[Kޛ�qc��7�PJ̊䒡|Oh��UǱQ�i0*ʗSE�׸�i;Ivl��Wp�uW�w�:�@�h��u�|�����]��7�5���3֫�G�=���r�y�3�&V0��V��A�黲-�.,j��Ɓ��cO�[���Z��fyԛ`]'`��]Q���O�d�/��xzcy�(����ؠ�����C+x��z^_֚4�9����gdB��\�\t�H���c^_�ќ u �k�}��z�*�G=�ɞ�;4;��עm>D��oX����v�!���Г��7g��	]�,�{F�c�1����zbU9>�%�B�k�!+�`K�K�=ҝl�iwjL/~=�9t�HQ���� O��wk?y����$PTU-��5E�� �ŵ���d�ڨ�I����襜�n�Z����@�-��0�.ʼr���#Dj�ϟ�]J���
4�F��yr��vZY�0M%��L�cl�p��*�i�s��h5�[�Q�K��e���3P�\ʃ��z�K��1d��4͎�ԥc��Ǆ����J�Sz9��uX�����`���9��mӞ�+�|������ɠ'�32��־K[�9���,�mv���]�I�K���NB]L��5�8"�徕'vW3�^��`�k��^e�/+��[w䍍ܠ��� ��U�M+9v0`�U� ���YB�W���pL*���,VD�
�t��Un�]X�,PT򝅎�V�5�H
$��PR)�me�X�o��-�Qh�Dp�m	yun
��3f��;5��8�6��T��7m��]�&�@_�@`��F�)�MT8��G ;���5�sM��ج��V#������n�w���qk.�6��V�mEEi���bȤ2�$�!fHۃ��6���*2\�wQ�̫2A��8��ld&36,����-��-n�$�c%e�Ad�*�K����rs���������r�]��S�	�Oq��R�/��'N�ҏ�� b���e��ea��J�b��-Z�e!�ځj���='C".'��4�cN_z��j.�{�	�aD����6��:ڪ����ef�!t<Ǘ���YI<���g�mz�*���������Hx�_wY���dj��if-�[��)Pc4�����M���Z��<��W�����X��������^�Y�(9�c��}�j��.��k^�;'�b=���gE�X��C�c_j�Ep$w9ᙽ���cB�/`v�M%7P-��{K�6I��<����t��$�{MX�4H����߷�|��D�/��/bq;�l�Ϫ���/�]g���S��:��1��;*"�����k�G�Z8g�u�����sm��j�>z��=�z%��mw]ج>��Z��:�@�n�;3**%RQ̰a�>�0&�s���;;W�Qb�����YV�c�Ú�Xg�I�#L�սw㋩�<Z�Ð9����/O�b���B��.���*ɕ*�(��7f��͂�9�[�s�Z��ݻy�8�p �Vվ ���Bm�d�Dʼ��"�_�kV�E�,FKqK�.�n�e�F�dK����c�꒯7Mz7ϵ��i����,����!���q5�����_}N��ln#�q��l�=�G��n/�`��/.(?Q�A*勺������k{���zF��=��NQ��ٷ���dwtn��=�Vfe���|ֺF+W98�Ʌ0Wa����
�Cb�q�k@���͎]1C&�1�e{�`��;
������r_�"p��:��"_w���G��0�bWk��G��Z��p�w��R����@U��d�ĵyv����/�o���D_�q�t�莺~I�����%Q�{~.����ЬŦ�(��B槎�e�0T��R���\�����N�,\�Y`���_;���ZH��3n�*`V��هޤ�Qؤ�n��Ř�ί��wvXV#�_��T![�h_��0��0w�g��iʿ���%U��f�d��xk��s�9k�i��9Ï�(�x�Q���qm5�<�g�h����������^D�%�k���Oc]�Y<Vxe_yK���E�ow��s��9]5�h���[��}[�A�L�3�R�yJ�%H�?�z=���&~#.c>��75Dw��sA�e�O�C��>��m䭶���ޔOM�˭\��R}�]�#�Fz<]]~k�[�署�����0 `�fA�`����&��U��G�󍹮D��eK�f#5ǵ�T��~��[~������ϲb~�m뱷ܓ��
���sC9ˀ��)���
�'~g(]q�'zM�"��F��B��17�7��\���ى�!��WiEL��1fV��q��fOy�Zi�1�*e�����/:ص�T���Oj�����^G/H�O��ι�vZ+'l��f�wT�FZ��{�膞��0dW��~�]V�r���Tz�st���9���t�&aY"�P2o���} ���~�_j9�j���F�qt��s��0T�a) �>��ֽ�ro.�W�y�����OO��|������V���Tn~Xt�Yʰ~�RS����\�1����zf���o+z�M�5��[�-S�`u����WJ�P�����\x�U�ɬ3)�J�(�̺!˩e
���/̦{�αv��[K-�8�B;_qFq���E7L̺��2X���"��b�����$��TS5J�J'�� ��.nYB���9�4�wݹI��+DU��e�,�`��N�J�t�)z�r�ԁǋ�T��fd��/����(0���	n�鬢�Ut��5hM���(�Mb
��6��Y�$lj*�Zt�/ͺ��˂������;�Ve� ���h4q�Đ���K,�]�MK��V�4N0��*9�r�ʁjrs����-~{j�~�N1!�plE%��-n����#V�d&]�b��m%H4KnƖ]ݱ	i!M�6ɕ@�j�P	�P�VKS$b�LAnY��Wv�$��,d!.�ܻ�E��q�H,�H6�2&f(�����q��,fIs,��R9p���3QY�G��M�+�J:�d���K�q������_�����#� f�����u跀t��Վ����Yn��#/�9�nB�� �Ѧ2�wk"��}���ֽ-{�[^�|�g�l�t�~C׻<����i�=3��'����Y%D����޻�}8k D���G��KGϲ��-I�Ca����S T�0Sn�_�)Wg�8�������r�����ߛP�5�cY��Ȯ�L	O��*Ȕ����-�2ɩ���U_}U�mѭ��9+O��̕�_���w���SM[��۶��,�X'ڜ9�{�O1&�ɚ��>pz�N����s�֔�כsp�玳�s��!�CΓ�mBı�V�u���N�\3O�=5�P�[��h�0k���]sܺZ�&�{����)�6�`����j�T	��	�}!�K����+��}&�ݩ�Drm�0bu �ܽC��}���}ٚ1�k^}�{7�/^]����Ug{����tƶ�է����5�������rcƱ4�M9��m׭�߹��Bӭve�ܶ�b�SZ�o7׍|��8��m��2���߾2��\��D�kR�v���y����4k�������ƾ�//���=�����q:�JW.
[����/Uu�����ǂT|��!��\'��r��Z��|���f���%�y���-o���J�3�>�L��8Aׂ���'��(��>�xh3���͝�o���������;�G�i�^L�~����:��$��ת1k܇u�&Ǐ�;.��Ӎ����a{��܉�I�{~�V����(����y7�71�rN�J�i}�=wZ���w��ߋN>����8��y�|�)N5��Z�<�w�y-�z���}���z?>m<�w*�i��/���5n�4}��	��c��3�C%�<G�m�c��p���f�O�`�,�Q���73����<�H��s��EY]���C�zD�����1S���֑��L�]�Z��ǹۭ�F��ʾͳγ�Qi�J�Y!�>�o�^���u���-4p��I����ý���wv�"V��ӯ\�ڽ~{�~�\���Ĵ-�î�g���yݾNM����H#�ZX�%����u�ny7�^�Yt�H�����Z=�~�4�������0|�|N���i�M���ܯ��L��:άq���>讦`��N��aF��mn�Ɇy�GKiQ��Wo,��ʝ㲮�%YKFB��>���{���Ӳf*xkM���2�w�[5�����q��P���1�~b�"�U�ńE㫶�
�DF�5�ksM�w߷�Z���^��Ҧ�����zcZ�y��o���ך�뿾����q�Dm�u4���i���}{��3������O�ɭ���:��_Z��bD�-��#��s�׽5���9�u=�i"cX�ߵ��ӻ�w:;~t}�zt�-�	-s^���﻽<�3w����=���~( �~��C��e������%([[��y6�M��>|��x�a�J;��eu��&2Bf����h��9&{�|�����';v�8��7s|���Û��C�-�y��ϳ�jR��ɏS�S��۶ڹ'�J��%�+[����x4m��:|ֆ��Y����3���u�!��|�MjW��&���˿�iƶ�ܬh�"�J��>��x7�u�u+���^��wn$������x__.���磌��s�7�|魿�3R��(��7�{��g�5�h
LՏ>�*��Ǽe�:bw��u�Y����Z}�{�}r�\��N�sr4}��cI��v�{��=cC�^K�i�uקW�׾w�C�ԉm{��E���������Qhq��[�L����z�w�jy�NZ��M!2S�py9�[v�dX�V�L�usSZ>�V3֪�+�0UA�K
�S|M�=jJcB�NYY�;�".�3��d}�N��J�.8�����޸�s31���x��ǉ�7�wћ��ƿ?&�+�&�d4��)���ˁ�n����i�I&>�2�����ݖ�N?8�!��ib<�]��ѽ�%��y�oQc��B��ݾۨ�P�uZ<��rͪ[l���w}��nƎ'Z�S��O��K��CP�G��O?&�1"_e��ao$J�"op��~�g��s����}
��",��[5���n���qg���L@���Җ�)7�Z��N�K1V�߽��r=����?��z�F1�N����s�u�Cr���]9�>U�+*�N2�)�HX��馭8Q�U�e�7�>��8pS��6��M���5e��k�+�5c�����7�]o�{�h�kh|�Ѽ�~����߷z�˅���e8�J�mґ��aO�}c�0`�1PR�A���8�{dO�j��=Yd���bv�F��*޴F�z;q	���9����3�.^|N>P���խ��QA����&�ueh�Yx+�<�w7ʣ�j;�iT��x�# ˤi)2�i��-�0u��P:���
��;U,�t�f�,s���A�B��tq��FQ����� ��OiM|��1��]�7n�|2vwj^����z����o������io,�k-U�>��D�-̕�=�HZ%���`q�g�J�P�S�5�y�Vׯ�\���Mx�}�F�h7k����+�=��ɝ�L6�U��v(�=���2�b��h��N9�d�VX�p�5d���[L��HG��^�%a�S8д�P���et�vk-o&���N�g9�WHìN���&����j�]>�&:90 ��w��F�`����%����}���ĸ��v)~�i�c�a"[���Ʌ�B*4��۶#,n�]�B��4�E�B����$�W��B�4[�H��*@
G�@�I����E0�ЎKk"�qe�Y�[LI�Z��-�k��FBD�� ��.[#A��rH�X�wli�e�H�~*�T�P&��_�D��k$���dK���\\�e˵$�q7
Ҽ�IE@�f�O$.�?7�#��|�;�V��3_��_C����w�zjV%�i�-`�q/��ݾ/�s��;���ߦ�!�b٬ދߥ����!��C�O��)�<��1�D��F�{�r�j�k��X�Ӊ��}����-����Y�����}��}����M&*f��:�	�F��m&>m0bq�c�B�|�t�]D.3S�.Ǡᄨ�c����YI��4�����n<�P�e���Ⱦ��v�ºn�yK�po;����c����ꯣ�n�z�-��&4g�����O&=J�~�:|֩�����[�z�bu��m�i/��Y�c_h/7�)��W���G�!�Z}=�~�+Z�rt�ɷR���߹Ä�߰}>��n�Ss�3�~t%�>�l)	��Y� f�|�-�ٯ�>�|vU4�N6+I��*A����iv:�5X>"�
������N��wϵ�҇Rл%i7��+���2.���_���~���A<m��ac����҅�CMr��W�}�NJ���5�4���i�[?Y�j�1�o��9�4i0LjS����7s��vm�&@kQj"�_׽�~���o�6����Kk�q��W��y4����C��i٣�:�5�>m��km}�\�ۉ��v��sW���&��c�}�i����'M�f;M'[KL|�>M�iy�Y2V�������^��M���k�߯\���F�u�[�6�\�z�g�g�}}����*��7y�}��9TAȣ��z�}�{Y�~�������_�ȵ�M�dR'}�����Mk=+�(F�6���m��gw��"U��6�=�����>~]¯p!���|�n��%��|���q�h��j�[:j��i;�i������{*��&<���������n��$�.���f�j4�1SEA>~��>0W���{�]v������{p��Ϸٮ�+��?5�5�i���^�&Rz.K�P9PL�gt'R�����;-�久���U�Hu��چ�im1���������%-�O�M8�L$'�^�G�(�[kz�k�f�5n��\�!����=p1�3�m{N}�l�ej4�m<�v���|��8�8�tҕL��};~�5���~���뤭!m_Ӛ�RRϧ[�;�g�~L=C�ܝ�s'l�D;�sD�'}۬���k�o|�P�\!�Ǜ�ϞV�0h�OV�� ��N�_�z�Vn��w�l�m���YϺГ���U]�ݿ�ƿ6��cr�j���_{���g�[k�Lz�`�ӛܛ��~���9�y��Ch��y-�upߵu�,L�=�B��{��kþ�ؕ*|��0g�ǩKj|}��4uRӏ���Jǭ|�^�>��!�8׆��G���v�SY+�f�5i���*�ZX�n���L����vy�i�q�JcO9��y�䆝��C��s$l��ό�����Dg=����u,��-��;�tN\��)s��V(�.�?PUo�Y�9K��߷9p���y\j�+�M�Zu-�駮�RT���ۿO^����:�soS������z}7t�ih[^N�^s���>M�N�ƺ�*�5s�z{5�O�}��v��B�Փz���m;�=�����j,C}|���S��_�N���c��[I��ɯ��Z�uS��־�+|�����?_5�b|��Ь^��a�Y��j�&�}r�\o���Aϧui6�\��,�k�*]�UﹹY�bq��1�+Ojj�7m�1<�m-;�ƿ&�M'^<ޭv�&�1X*(�e���U�T����?��$EƧ�cϡnƭ�ߪ{{���ұ:զ�9~�k�{���q��h��ǯR�߮�k��v�s�u�KZj�HSJZ^�{�w���>�!��W��؜7�����~s���}'O���o���|�#&9�����1�x;������ŌNohj��c/�G9�x4U��Nx`�O���jt��ݢ?�Q_{��������f�f�m�NJ�0�f�W�u�1S�������'��������(]�w�z��p���g���z�MY7m4��bq#��ǈ�x�ۿ���ڹ*F�zV>�@�o,&A�QyV_β�j��k��� V{P]� y2���W�OyW,-TS2?L[��V	�(�M��J�yS:[��]�*�_m���\�}�����ߘ\?d,~"�~�3b��)/x�-��p�<Y�l\�<�K2�#��$qla���z� �U���^�ǐ\*X镁+R�q�8%.pZ�,�{rH��9����=�-�k$��\���u=s=t�u���}c�ѮZn��	���j�Pi"�=�.�{��@���.�8�ˠkt�t��(;��.���=��>U/���/_aL�t�V<�v�J��v���D�}�+C�x�#��b��i6�*�R���9K�b�|l�TҴZ�X�lK�ډ�a �ف&��n�����3sf��jE�����RL�<���Q��`W�����Y�KR̥ӁiV�1����u[E�dj�S��b�N[�ٙX,"�I�ΝnQ��;�@P'Zd3�9�1�9���KE_b�Ϛ[��%^�5����VU�(ͺxU3�a����sH��J��R�������h�Ǘ,ܸ�ޗ�n}��M�v`�"���sTu�Z mnσ#�vR%�u�H��Guȏb�� z��w4.���ڈ�նܶ�2F)-�$n��nŹjM\f8ې ��L��!�@0ZlPt�R	�M��R]�aw�$�9�Z0��ai�Z�i��� Bl�]!� �&]��ZE,���ܨ�K�q��D�,�F��L�ܸ^0����Z2��5�\�w��9-��-�\�p�E�e�ܸK��fY.>#���N�$³|��V�˫9IZ�/D{R\���O�g���V�Q�Ю�9�[ T�c������ݺ'A�}�w@�YýRRd3���j&��S����.�@.�wl��v��~�R��><��X=�w'��]u�ul���u���ϳ���Ó�����=�֜�O��A9��u���vw�>��N]�{�����I~x�ѡ�>���rU��D��D�}�l6������ͩdO���{ޅ�=��&W�H?�L�ٕ���Vu�V�u�X��0$�e\p���l-�������Aj���F_���w��_�g��H����ݕ��6��2��Aɦ�ڴb�]�p����=z�U���e�4�/�x��#����ʆ��3u�K�H�������.mW�ND7G1�p�g��{ۊ�z���xRn�C<#zV���ۈE�H����M�J�@�A��]/*"�_1�n/VB�R��D��@�|��b~���ýV��~�H5��Qp�߳M���C�&�Ơn���^u�.���^'p�{��umj�w�E>��T�c1�c�}�2SQѲ]�{�'t��0T�]1���j9�"�p������^|E�1�������ô��8]������6���-�꯫����_�����wvt���I;d2!U!UYKa�r7P��en��+Å2���/̇d�.��^�KTf��
6�wɵ�-�!���v�X�ʳT����;ˌ:m���Մz�W�C�ډgN\��zo�e�Y{� X~Nv-O�0�&�#��D$��G�$�%����t:����Y�ͬQ��3�`��+���4�v
e`�oֺ�>nE�x���ϒ]i�>���6��b��αW�b/+|�J���K���)-��l�g���E��
���n:�nU�{R�C)�Ό\r�+ٹP]��Z�ɽ�}� ήH���؄�2=���ir�<���k��i�&oࣶ��߿~e:�oyg<}�s3]��.�4��lm���؅br�%���(ov�1ݞOGfV���N�7�5hPp����W �[�;�7.�cu�K�Ko4Wc֯ȉ࣐������6򭲄� =r�� �X�Y"�m����FίY��W�Q>Y���໴��u5���A\ހ)��f���W���x_���:Ε��!���<���c�ݷ�|6�f�w����&� ��ySy���&ml��ʄ��r�-���f����=�qf��N�o�9��{�@�\�U�}�{˹ '��9U��T(1��p"����wk�ep���Z�c��a�����}�t����!��k9��A��Y�1��~��xܦ���캴;������}B�#�����0/�R@_=lӷ{'�rԢ�kV,d�36�OK�z�w'���U_s�6s�������j��s��Wf��JY,yK�ӻ;>��6��a9o��z�Ll	'�_4��Bk�H�lJ�N�=Y��L�I��(�{�@��o�w���)e����b�?o�`<U�*>���"�D��9�s���$��Sc���fp<����;�n�ӀZ],�Q]]�Vh�F�_�C��m`: �m�ͩ2]Z�J�8��yJ^�`������Oi��z���b�q�����'+-X�H�o$8��ז!��i03C�	՝rw4�E'+)��M�r���Vg8�#�Ø��g8BMm=�]S��6�c���&ʺ��
]�'S�b'�O����v�N�8��*D�&%AX"��Fi�V�]'��jY�U� �I�g��VX�˷-�O#d"a�B��Դܻ���]
�.�e���I�l�r��U�0Q���w�
��c�x�<�Kx"4I�W��"8��pE�R�Y �(��M��,E(TVftU�,*9T��#�J� v��+�F���ղ��d�d�iG.��fL�V%�,�H���$�����y3.�$�Ir)r�*[��˹r�j�Qwm��7"�	V�ܼ�G$�Y	!-����FRRݐ�TF�%˒�$%	%Fڗ �4��R�cPG"�ݎB
4�%���w���~���\T��ޮ��l���Iq�\8@�%��M�	���sC'�m=f۳���>=���X[�:�-
�Q���*��n���ue<�"u���Wy�������:Ǡu�S`!+l>�-��/ea��^+D+��37z��4ڒ��c����[��n��Ջ_	U-�9��7X*n&�F�_y߸uӥUv~�_����=��'��+�����y�/O&{{K���� �����4!C�{y�L�}�̝7"�R��ۚ��%G+� �����{>�ճ}hdʀt�t���گ|b>��ͼƫ��^��b�f��C=��wKQ �v���}E�ܗ0������/��?m��oǯuYQ�y�3���.�N{yT��í]�%ײ���4����D)��G�}�{�<�����+��kP�jr�OA<����u��1E��Ҧ�Qk�^d�a1���X�g���b�;�v���։�����8��ضO�W���"��ݪ�J��u(��P�����[����<�l�%��>���ǟ��۵���)�W �O
_iG�b�5�}�PZ��D�˨(�>���u*Y�&����-K�{s�@�.�^;&2/�#�(���9�9i'����9���Ð9��������4�����������2We���&[�d�V���y�il���y�Ƭ�T�>�8Nc��6�QY5p4�Ӈ�LI��IIv�=�1�+�O�:-�Q��Y-|"5%b�������3�d���D��N_=���ȫ�/�_}_G��%o�X3�.�2�ŵ��s)�~�f�X�{!:��^󡅉��mO6�>�M�h�nLV�4��;�W6���jac�lTbpB����b�mE�;��P;�6p�⻅SШ&���=h6X���k-v$�tV��oQ��D5�a@����}U�M��f�o��S�^�+ ��IJ�����W��h��D|����q��DQ�+\睘^;�֐��!�vx�O���������S<J�c��GU[p���D�H�k����^{�^f)o����[c�L��庘��P:�V-�:���.����F_ݗpd,H^�)���U�v��G�N���h�5
g�`�z<�s�fP�_�m�;�iu�Uy��ܶ�[2:]�Me��/U�>a��>�9���9*�u콬��ĕ�����v�|���\C��X��%�wvo<���7�5ε���.K�'�C7]��3-L�;wl���\^�&_�U���]��
PR�c��Z]�Zǖ��?#$��w�1�ܒ8�R7�6�MX��ǈ���$���� �f�^o��Is����Þ<Oj+	Z�X��������NNw�KbYK�o��gr���լ�|���|�`�]�1�*�ށv��Y݆���$\�<J��U�⺮8�ް���*y4B;~|�L29��iߓ��ߟ`]����%+�8��t�.��QX��b�A���.�)M�ׁ�����<uٶI�*a�O
3��Z#͙��p�� ݚ�@gK���7'V-��Z�17t�ɜ��9�.���w� �[w(���m3�1��P�+GV&��mum����+ij���M�TM�h9֌�3��V:��O7�n����#/y��4r�8��Ռ�e7j[�J�N �� ��.���Mb�l�i9��i�0�l�V,Ee��ApR�q21s�+1;��X�vYY���ȑ��b��2�E�+)*b�GR�������7�<"���P&��"�������$�4��;�VX.�0ʉ"j�4^Yu1�!F��TFD)K�*єm��Xă8�J`�R�.� >�)�"cj�5��F�,QDDU�E�@���CJۉh��4���cR���.$UDUG!.UĻq%�%�`��TKH��i.e�����hG6ʉ)$iTiU$����)V�hRK. c�0eȔ�lE��-������ Y����W2�x�v;��b��3:�:H�GIk�f�ju�-��t�·z;�e��t�1鋽S5�z$mgi\��$�4���u��5�Ds�}o-!��3]drVfWA�#����#���#�{M����q@8�K!O�ƌǕ|�U��t}ݣk�s����Yrt�a>���W��̭��7=#��e�m#�!�:֬��c��c�O��@�(
�ٸ��O�5�p���1���SJk���#�}1���)�{|�D�y����WV��m]=v6��Fd�7y�~�::7��/��2���;�sz�#��uM��/����U�CD2�b�̽��M�c��X���*���njEs�"n�:��p�{~z'�qM�A��:,�_�f�O{+����<p�h}&���)�{]�	�|�D6x��;{y'�S����a��b�`D����ݝ��qvӌt���wG$���]�y$��o�;,�:�kw��Ig}0�{kY���y��@��B;���Yp��hUe~c}���|���t8>�^0pU���2&�T��F`�|�����;��&�:�51���<m쐣Ju�y���.i�;�=�+�h�ĂKN,ͣ݁x���fǪ�^-�SƤ���i������/�p4TYBuR�l�n��*>83/d��Ք�s�$GWu���'h��j�Ε��n��]y�_�%fd����)�ĭ�	2���ك�u�}��1�K���X�ϻ,	�:i��]�ei=��~>�F
���`弴�vku�^K �ў��5�t׸��3rr�����s[�6�"��6�W~���.�2F�E#G�����ؤxL;�Z����w:kJ{���%�f��,��`��Ր�@��ǳv��<�UCPðp罷����\c�]��A�'N��t�Xͺ��'��)�]zY ]�k-�a�<J�C����)��s��iȎ<ᗽ�z�Y�Gy��KČ��|��M��4�.��/���k�s��m�/�D�Y�=�e��M�;!+���h%�j��	��n�][B�@�[] 4� ��n�s�!������ǜ�_��q-v-L2�lb��tr�Qv��ȶ�{|����.膎Z�[.5��j�iC�F���h�Y��Tu$�V��i|�^��3W7��Dz����5�^�Z-�p����Ϸ���Q����~A����9�U���٣\�B%�vD�X�mon�b��V�*���*&��<w��HW�`k�����d�M�U��J�0+��ʌ��wI�x󝍚��M����to�3��DR�8[��b�}+n����^�T��V���o1����d}�Ki��;�]����e+
yK~~�6֮�[ �qDQ�8���|E۳�����b����XV�-ך�����8f�|*uj3ը^�� �$U���W�%ľu��F��fV���n��������$��8��P��3;���\X�)���͹�`��2��GZ	L���3s��ܑZ���Mޚ9��t�:q�v�|2�I�b�*櫿��8�Tى'.�l2k��d��3}Gw���'VJ)��Dt�a��RI�E'/v� �|(c�6�]�h��R�l?*�O�P`����)�q��ȁÃ�F�8�1�W|a�M��t~��u{0�̺���$
��K�=�ΓHVX���[�y��A3��0�&����n�]B�FˌVU!�*��Me��:hVZL�d��i�J�ހ�4�u�p���kh�ӥo�U+K���!�� ��ZX������V���Y���],�HQ�쁔CoMV�M�i�5{J�W�y��:TTԨ*
=j$�)\aM+����r+B�*-�%7,KVؙ"��-�*��Y�
�2d���Z7���A�.Kij"B\�j*H� �h[����3.Ѥ��&Yd"*�����KW.\Kh�6��J������}�ϻ�uM|N<�-�久���U3<YN���>��_>�4&���˅�RմWD��̴ ��e�����X�7��Em�J��\s,PD6�p��Z���UFK�r�Pvz�W�s0�Jc�U�⣝�Ws��9�G$���c��gN��.�}v{.jn���Aٝ���[`�0>Y�*6��V��J���c�}^�A�z�6䏂�<�uE�iƫ�?0�Vv��	ng9�޶��k����&�p�9б|6a�d�B�d3U.&�d:\�n<�Ô
�s��Bd5��9 \�9�r=�8R�椠.�mi� &?>{FmA(�q���#�u�@ĺی��f�J��S=^T������wq��:�zG�lN���T�S}e��5'�5����3�焿wt�w�k&�����f�t�{M���:��Y��'-�p�K@^�Ig|�I�\��7�8�ŋ���1+U�9F��G��[��{�X%���O�N�cT}^��ބ;���*֗���k:�s��IǮD.�����౦�tO�y�r$�a^X#aI���N�h��Ly��l����Z}:�[���ӱy�cO��az�.\�VA���F-;[�RĮ�Y�o��>���oc@�e:���Pg<2�jC��O$}��i�x���ƒڽ�}uz)�f,���q5�:�w�'K&2�k]'�sw[��)�sj�]����8�!w�Ų'{���7O(��wv�Z�X�Y���(�9�Hݹo��6@��o�֋R﫱��Ǻ64���Y&�o[��,�|g�A����a�S���7��nfz=-o���YX��>Nr8�0��"�Ȃ��B{O���.�3� @)�j"L�$�}T~�%)5t<���`�g��[�4y-���f��W����[,v7�sRv�>�ls\��}rMo'l7��	�m�ϩmg��.������z��7�J��7-�-�J�:��yj�8+_z�T�����Wh�#6� ����g`t���;Ë�����י�;	�:1��2����Ɍy��&�3�u���]�egO���VGڸ$M�/��+���4�����Y���7T��zox�ְ�9�è��՗!4�;a�=~�!�3o�\ȩ�;�/ʮ��]lb������P�Ǟ{����=7��ѪU�*f��Ϻ����x�c��'ua+'l��Vy��!�G
��._������ج��q]Ƨ�@j8l�ѐ���F�+뵋��s!Tl��H��+53;*���k+^��8��Zr��yW�\�U��kz���K�.Ô�it�Y}p篍?��6)^`��g[só]E�Z��B��+[��{�Xݧ9�G=��*lD{�_��Էi�_m�5FNb|6-�\�o�+F��s$Ω<"�4m����3�|Y��с͈���XD��m���UY�!>#���ā�9�䙽L���\[��=��,>�t�B������,:��R+ś����8�+T&=��"��.\�R� Σ�u]�Úa�qRۘ-���@Uc�Kz^>���P�}�uo*���Մe�i�/�N�P��5���[C��9�QC���تe�Y�[��{��b:͙k)ۍarDM	(\¢��y^��q[���hz�y�%�@���Q�>6U�;�7���`Ɍ����]���"ql�ݩ_�fCv�+��ՙ@����55���}��Թ�h���E�*붊�q�In�C��ʎfu�Ƭ%"�v�,�*?����5Z`�grM��9Y��e����B�nD�q�jƾ��=\�,�FT��.J��\ma���cnM�\P�FQ=E���CI�+���́}��/��jw�ZP��)J��"+H�"�kr�lX�T�ARK������jKK��IM)j�j#rR���[a(F�1H$i�7ubH+rU+p�"TbIM�[�g.��[�qu��g��� �I7��8������4p;���y�/�}(D�׆_����*�ڜ����+c�ߦ�Ymw�\��i��;�/��6�L��OMbOq����v�z��1[p��{��L��U`{eX�#0�k�qǫ�wgS�=��2>����L�FyL�o�����7k�ܔ!C%[&���r���[��#�Uq��n���.t�	�7B�~�KǜwWk9�}̃�o����`p�A,�m�N��x��P�ʭ e�7��K���^+a,�ݥ��4x����ξl�%ݝ�%�S�~���ذ���m;<��讫ה�����<3o�h}Fh��w��ҽ[i*�x���9���^�ո��BNr)l�C�뚗��H��ܯHJ��K���5Q0�5�L�5k���,`v�Е-�4X�b�ׄ:���0����Uer޽�|L��;��D"*��Q���8�ժZ�[=��� �/�|]�����F�>����btJ��0!�l�º]g<pZu�9�R�r�,�u�X��n���s�3�<�^��N�P�AR�;\Zd�U��S��ӆE��Ar3D��Ԑ4�v��1i�N�[ia�ˮt�ګ�}{9�2ϧ���
���j��`��Xz�=�S!E��,�&q��G�s㲝��l( E�	g	�|�q1BR�E�YSg�������e�o��#sLri�]I�W�ɧݽO��~{�zN3[�2�'�*�7�U}.����U=�~�������i������f1������k���n� �uO-�L�{w#�B�������:�S��؍�=��{�D���������	�Ү�g"�N�[�qsI jE�|�sO</��r�*VN�_�s���Pʴ95yJ�[�ݕS�q��˚�=���
��h�>>������3 o&=�{�E�K6v��T���s�RZ;6���Wӕ�D�ê&jP{[�E���'�δp^h���77��\'>�"�]��M-0��w2�'��Y����R�.�3w�R��R���W�lH�aG;�6d@k���V�LeN7V3ɾ�ej[[3F����l�6.����
y�39v��qҒ��B��'�+7��GAQ.�:����'�X�x��	M�	u���)n*�[�״�w�1��y�'�B��<Z`�Xv{]\X�<6ޗ�íKOfCڌ#�-��Z����1�2�릸r>�Wd�*�B����a��#c¦i���l�)�Mq���*��uz��oZ3�+)�+��iwDs��V��K0�/,���7���.}�[Y�ou�ݛ�����Ó��R��e�(�����6�mDfŭ�ӗc�q��\܍J�
�ys��jw;7���sYz� �&.�ڒ�ҧ����ў׮���E7>c��z���f��c��$�>��g���O�_��XT��#U�I�JQUZ������������6��	2iJX�L��2��<����ٟ!��
������X9�e4`4�eUڳ6�1�A�_u@0�-3�|��UW�A�l\���p��������k����L-��ĩ�5�;��fӢ��:U�����ªP:,���k�l�UW�g��m�Wc>�X!Ҁ ��  ?U�"Qjv���c�9P9�G�� <�P�m��W��w����P�<AUU����R���H��LЪ-��0�4q�������)z�
~V�Ҟ��7��w���޳:n,s��`a�W����UViy�-��:,{k�પ�=p�v�A��At�ЩLn�QV��;��n�>v5<UU��@)��z�8�����V�G��G0,�Ⱥ�m�?���I�}�Q�?3����q�P���*���4vP%D��ݎ�?��w��\���~8R��(%}�����c��=���S��ߘz�Wj�=��'�r:`���z�f|�z�A���<��I�6`=tCr �T{�UU��r����;���A�d�P�̋� K��\֠ �$�`���RtP'�f�
 "ܢ2"�`.���}@��P��yE������ �L�ܶuZ�XUU]����xh��9��-�v�����o���6�ߩ�������z��>�!��g�:�
��؏V��v�'�=����+��m2[}��@UUzN����,� R� y���OH*��_2�@�ڟO4<�8j!����6���<=[ �tȃ�J���K��Y�N{�7�C�����>�ǌ��_�ΦN��}ށ�pUU{zג�4�\�rI]�채̇�IB����à���]x�˅�(�.���z"1  �b��0�8�'�yܹu�@  �C��BE�[n�����ف��A/�{��n`�$W�a�(�ݮ�u����w$S�	��