BZh91AY&SY���Z�#_�`qg�����*?���b'         ��    
 
 ( P    
   H  
 z   J    � �  ��ۺ���7�   �   4  � i� Y�  �h��4� )!��  �h 
   P ��
J�(��J�R�TJ$�)AR�P
E*H�mUIJ���UR��
�B(D��TU (���n䩗l��D%!RT�DԨ}�Ufb�7��u�I��C��<T���t��H-P[�H��ݸ�Sw8� P���@ z|�N�:���P<�Nt�꼎���r�r��9�U��\ ;�덵��C�����*��   ��#@�45*�%(�EEJ�$.�
�@^�9�9�8f�O�{���J�,����Xqjq� q�iޱ�Ѭ��������C�rr����  h >:  z5��>A��}�= �9���7g�1��0��<�y4��&�i�Y�@�y�U'vz{0�oHx���Ǚ���x4�@�K�6�  c�*P"�DAN�:�'�@�q�i�:�`;�ǘ���'��(W����� w��cG{:��3@�OE�FFy����     ����5y N�J�9Ч���<�mG �3=���� ��&����n�ǵ���C�eo3�h��z�h  �� ��EJ������*)R%#�Х\mK���`���������*�p=�ϰް<�r��Ay��ӡU��>*�� ǫ��M  ��� ��N����{k���B��S&^�y*@2-� �I)��n���B���{�@(  �7� �*HDP�(����*������ r$: a��wJv: ݝ���:	wR�K 'd���   W�B���}�dʊV�A,�Xt.c"� 4��*:�J'tݎJ�n��7`�C!�_       5OĘ*U     	��S��RT�0     	�h4�j��QJ��     �d��R@       ��i
��0       �6�ҢJlCJz��4ء�=@�4�O)������W���'���?e�I�".�,���vT�h�0���
 ��I��DQ[S�DE;�'�
DAEa���������s������?��}���1DV��$���W�c��R��W������O�"~��!ȿ��� �R.p�a ��\"� �: a �a �. A0��
\ @0�a �!�S� D0�a ���!�"L E�!��)"D0��S D0��@(�a ��\ �8E�. �0��L"��xA�.p� a�@0���E�.0�a�"��!�\ 0��."�a ��C6G8@0��. E�.p��x@�- E�!�p��\$ ��E��\ E�.p�D0���E�0��\"�Fp�ad\"��E�p��E�.p��\ ��E��&�L A0��a�!�,��� E��a �0�0��� �� ��.p��a�@4E0�a����"��!�&L"l� @4E�!�"�&�M & Y D0�x@L"0��� �aC�@R�aS�8E��T0�	� &0��� L"��*�E� .0���*&Q0�)�Q ��C
E�"&�A� �A0�	� ��L *aȠ0�	� aC"p���Q"�a�D� �D0�	�PL �aHAL �a C �D@� &A0��� L"�aCE�C��AD� &6E� �D0���E �l�� aCDE"(aC��@@� &T0���@�*��	�UL""a��ET�
�P0�!�D"�DA��0��P0�!�@@0��U�"�@�AC�
a\ �Y�D �
�@EW�@ �"�E�+�Ap����AG  �� ��  �a�xE\" a["�Up��p�.E�
�@@� E� D"��"��T"�� 8D�p�� � Å.h��"��E��\ �Q�@0�a�E��@0�a�@���6E��\"@0�� A�	�p�a A��\ � ��l��\ D��L"�8E�P��A��� E��A�p�� �
 a8A�&p��0�� �	��ǭO��#���H�Oߜ�e�[g!ݣ+f���d���yh7�V�E��N�t,��9�nlY{w����]{���С1G7!��9��SdÕK�vI��:�U�04�*Ԕg+unH��٧��ܲu,�k-n��`�u�*�1���66��l���K7B�݃~��N�[�$zK^I�rY�Z���9i`M&��.��b�.�1,��e#�;N�!��*��$U��V��I
l7z)�p�7�����b�b�eVɮ��U�j�R(.đ��r��A^^M��0̹nnPݬ�W�g��Z��&�e9%m�a���ca�����`ʘ��PՓ6�a�jVL�ʷ�q�䩫%(�d�7�9x�q�ݔ�rRrjȲ�G�T�oE���f���,n��h�Ơ� �Q�J���G������Y�7c"����YV�ލ����^.ȭ�3���^^Y�Pf^êp]Lf��]X��bw3L����Vl�xr�yU�ĺX����j�={i$8Ĵ�c��$�y4���V����{3)!f�C��YfJ��+6�)��QGVҩ�,��ޜ�� �Ӻ"�,:�n^T�̤�J���n�ckq�Ӣ,�uU�bA2��axė�^a2R�v�����PlVL'v�yi�%��a�[K(�#d:uyIJ��j׆��Pո�� ��gtV���o�t�J�͔Q��K؝�UT��Û{��ݚ���(c�yu/]��]u�ҧ�:C�<����[���,(e:�UL������,�3�C�rS/j�^֋�	ov��ݠm#�j��E=�"�4�e"2�	�J�oc� ���n��m�J�a�a�غ+f��6��'��t�U�جf��zQp�YM��lי�U)
��R�E��^X�A�T��{Fj�k
5�0-�[:�Ɏ�k�36v�Т���h��W2�UZ���I�jӉ��ce�Ъz���bZ��dѺ��T�:^�ǐL��ģ�j5W�P���c��Go,Upگm�}���#e��35����28�,䁸�f5HP���K#�xŻ;Eɫ������2�`�����֪���S1M�`Z��D�gR���A�J��Y34n�YlRs2��k,��L8wov�R�f[SiMT�Y[���cU�4$#!��ٙ�rW���ٛ�{$��5�f')ݽ�;$4�t��+�W��U[h^f�gP�Z7SA�J�6���5V��.���P��FL�*�W�Gzh����ʳ��e�/*ۻ%\'}�p�kt�GvU��Λ
�^$�i�U=U!�j��7L��/�>���w��r���BՄ�F�B�^�"Y�5�j�GD�:��u�+�p�yv�yR%�N��,�6�"�B��%Ҭg]ҭ�i%�*wUh�1�F�.�G{F�ͼ�n��tNh�+7Y��t�d�M�z�J�{�ZFR2��7"��79pPtv�Ș�g^G"Bm&��H�����[���5Jf��yj�0Z�GpCJ�\x�E�n���QŹx��kooH�����v��j�X�ʗ[u~5R4ӵ�^7��lo]R�5x�L�HXAOS��WU��{�4����4�f��(��9N�N^�]�#Tŕ*�ӈ�>vZ�B�(����^4r�^e��`���-0cR�%�]z�f��Ko�!�#�uBӬ��ٯMU]�7e&o wpf;�5&� VzUMVi�4]*̎��b�n����W�-�W�l�cx���d<��9x��)��6V�t�a�Ì�Q�\�7��+ne��2���a�x�Z%�a�:��rS��a76��ьA�i�Y�vê�.�bҕ5t�
�e��zQ��)��6�7ց��V0Mw[*�sm�b����t����t��̪V��T�^�1C���+-K���׋;h\�*�Z��I�^�8ӡwHP�.EG/P���5v��GW�SP┶�]��	���P'����d�խX8.�i��v-�WaEF̷�6�Z�3)f�`���՜��W��,����
�۬rX�Z��n�斚TZ����[�ƺR���+�T�lB������;ؖ�ԛ-��4�͸u�5����r�]m,��=��yR�`Ux�OD���<bܻuF���jCkU�	������HUUf���Ƴ2�����f�����m���wu�6�VY��;�\tYqA�.Hup�l�sL"N��x�[ �t�{�ی�ef�s3]��M��&�I��=��W��P� ��{)a��fAV�l(�6�k7WH�_�G*�B���K����,9�pVC�����cf�mH��e��S�1@t��a��۶�{uG���m\{�)&�JlP��k��ɨ���+E�wy1���\[t�K��Tٖ��*d�wjL�wG]�i�y��q�e,a7��ڙ3��V�,��Z�e,���)�b�Ю�Z�͔�f,[yS)
n�[�N�V]e�uQPZ����0���ۻ+.F�sۯV�����5�&Cf��h��V�b+tǹ݌[Z��f]�/VT����Q&��a֮	�36�
���.���8�C6����lu�T(��ә�d�U$&�MQ�X55+e��å�y����#-z�����T�Y��o&�j��b���pl^���Z���t���ά��x
��P;j�ٛ�lL�EL�+��3�m=�C1��ڳjߜ���f�f�<���EG1Y��Md�Z)Z.���Ahčk���[4�Ү廼��o6��B9 uf�["��t$�[h�6áu����u�r����;�Z
�SA�te��j���Z��"#��um�v�WZ�pf�ӕc�ћ�0��ȯS��6�iU��6��M��'�e]�Z^]��X�%��eJ�q�U�N�/HŅ�۪bY�wU-�oQ�q��mjFX+eQ��+pK��n���,KU�j��/sIU�V�^źK
@v����ڥW���F�n���P8���<{W�
sթ�*�V�F��6mܱ�Z����hP6wp##٫i;(R��mfV�qY�MX�u�����/*���YUnmfk]cD��ۅ-��B2�kp�u0:���Ӷ�)C��3F�q��$vN
��E9-j�7X#l�혵6*�n���������l�@��-��U��$����:,c�3V�Ih��B�E�w�#wy��oo,�8��ӄU�RgV
t�T1�ڰ����Ss%C�(ژ�w�S��e�z�c�Ga���^��3kc�.���x�vA���8r&����7&10�B�qj.Q�aķ1P��Sj���~�B�ڥ�m�meH5L�E�����U��,7-6���Vj��h��a�z�&��x��`�Z�wI�y�b*�-�J�=�,ݝ��+cYQ�31f̫�!v	���,muv�e��+B��rki�ա8+
��0�Y�jҿ'.�p�U%���,�8��q����U�SfY��9���U��A�9�:�]'��L��z]+N����^m�Z�Ƌ��Q���p�+L����w�Q*Ў�zN�]�6m�.�{.իǧ.�Cd���yV�Z._�b����\��+ö�7��QǠK��Pn"t������y��:ʸ�F����zn"IJ�ӗpGco*���j;kJ�36��C)m�H�Kj��
���e�]��{�;l����ul<DuB�ٻU�7cl%`F���ƪ�y22Y����:�f�.�%�!�n��E��Ҷ����LW�n���4ݫӓ#ʹyo72��c��]����+Ɋ�i
�ڱY����y%����d��f��u��P�2h�(�;w��*C/�^��˨셉;!���jA��if��p
��
�:�нJ�(d6j�˦��:m饛J����!Q�	*
���*.K�q>MO������Eڥѩ�t����)҃e�7�t�whӃ3X�r���3s7KF��b��{�]X6)��Z�V;s��,��t���\�A��.�ͻУ�1�r�
���x���eZ���)h��~[��R�;h�uVq+�ͱB��n��5��r�/[f�;^iT�T
��7NNK����;3-�zD'0hb��ц�g����汪�F�^�4t�
7��Y�^1Ua�N�;[v��/tc%Y�:S
�U�F���F���,�A5̭�ƣoje�4�Ye0j��C���G����sn��uy+/Ղ�[lڤ��EȮ���ﲱ�6n*8�ͬgU8��͎��՝a�u���y���X�����Jn�`Ł��=Yz�9r��,,VVU^��ڧm�t�;�F�Ǯ
Ә�Hi�a�h�xv�]�\�Z��%p�.�`�q�h���J����э�u�5��	������T�{�˂K�a�f]��β��������嵙�9U��w������ތ���F��,e�$SnX(M�6�Y2ޫ[A���֋�A�0�ڂ�w��"@��Pe�@��ޅ�[�$��e�ftr��śn��XT��ݱ�Q��*��U��m�V^����{t�i�Z��Sif��%��=���o}yZr)�X��"��I�TK[�Uނ��
BW�_�b�Ȼ~@�
a�7Fת��H.bFòR��˺&se�������3�`��7��a���,�u���s/�hp�S�dmfh{�B��f���Q��"�E���x�T/5S� b����˗��n��Ct"LzK��:F��L�0�����3HDޘ�Ӎ��z�j������f=ʭ��eȱ7F6��z1[���}A��wף�<�c1�W&��Y%c��k6�)4���W���'���|�g�;�)����צ��{�a��w6^䥊�b��F��U,��GjXtH��D�Q��Hl�j���M�J̶!ѯ �X�`�%����w�S�۫%D��X $j��Ke��*�ŉM$����Qe���[3QʦNJ[X�:��B�0n��R������۳�UTGme�S��+I5x��y(��.�h!���%������f�PTvw.V��q=K�ۣ��y�7xѦټDУZH�h�n�m
U5V�fݧw�ovٲ��KeӠ�]</�</Z�Ò՛�)j�q4*颱T��ҧft�[V�Ѕ����#�,�M���J��!*<�U���ћ��6��ieމJF��.��Ǣ�l�,��FR�i�4��n�l��Ģ��ڸ�ɦ��vŢ��a�kci6�{�O0n��0ѹj�x1��Lm��Њ&��m��˱����')&M�p�"����IM��tq%Ftbf�M�L�,K�-�⼽�*��R�n7TuVך/)�u
��\����V.�g7n1���9d��"Ts��"`X�j�hSSB���t6�޼z��n�)`���)G�^ѺU[Ub]fޕ6��X�-<��VIsB���p�:�VP͗6��L�Tf�;�00�O���-lH�ֱ0���'a�wZz]U�I�7p�-�����Vc�f|�;��U�	�be�-�T�ڬ�h[�L*����y�v�	�ĭ:ݢ��t.S�e&-t�z�'nV�1��۽(�6q>��YO�u�{t���R�xn(^�Fd��<�m]n)[����;�jM�Yt��n:�k�#N�7VrV#j��m0� �.�ݝ4B1T:���	�������![�e�m����b;ڀ�u�7��D+�^rj�		NU�b��'�i�]�{*VۃN,nd����5��PYDI��Zƙ�KS%�����;Jb�>�?W���&��7,?4�H'cn,9uK�
{���AmVi�%�VE�ܰ����;Ù���v,�[�;��:��[Y��[�^�q��CdlY��zN/J:]�B����W�ӵ�Z�*��j�.�,���A켉�����pC��@J�����&��G��.���3*���ɻ/F˧5SU-a�xS�%�e�E&�fU��X�{��Qٔ�\I��M0j�Kc�aJ4'1�3H�.]��ə����gi5ovfG�YZ�f$Պ��^�;����sw2�)@�A������&TZ4p�+Ve+�x�V��Z*D�A�U�r��Wu�����E�2�@ߴ��R^�zM
HB���N`5�b�
l� ��U;��wlYӤ�͑툎�A[)�Y���9��5,#Q���"ٹGU�])�&��� A��V"�i�c7M���8�9M��;����V����V�35e'%Ve�㎯hG�$f�9��+S0�sa�w6�'��)j���/��R�0�+%�뽪���k���{4-����(Щ/v!w�Mʘ��2ڠdH����u�n)����ǹ��-fj��f �:�a�;�kl�]�po��Rt/^l�H:sV��/kq�bR����*�y��,4s-*���F�I7p�R�O/6.�zTx�&�7	x�����0�a�nf�)��ИER2h/v��/�x�SE�R�BKz�1��ĭ�P����y����ތ��&U��'���\���Э�v���5Ul3!0�0魆����(�x�=�7dk�ۘQ�y��u�V��pU-4��6jA�g�/F��'+hf�'&ݣLbYE�����XNq�.+8�PL��G+Niǔ���A�fj1�^W��̬:|I��V�~W;`l�Q��[�ѫm�̅�9�CRK)Ce��jL��MсX���8�c�N&���?�Y����nYA/�{Ҳ����U�����Н={��Tܛ�*�K�n���>+W�{���խ���<dN�	8f弼�:(��U�2]ѕ�*��ܰq1x�5�a0�|��O��콧�yۈ��n_+#������v�c%#Tbp�b7��j���<S���]�oF��%w��Vj���4B��Vqҳ���՚Ӹh%uz.����),��*�V�1hߍ��XG	f�<���ȲMu2�h"�/wv�2��慖0X6ʹ4�wVj��u��s�
�P���E^Y*����0
��H�LN{�7{Wz�nn�^�,��*ݑ}�a�P� ��ɗ0�7��'R�b9bJ�5M��f�%[4m;��y�[9��+:��@ߪ�{�ؼ�ٮ�5����Z��C�����6;�ސ�  �(�"���2H�* (H
$�#"	 �"!"�H"(H���"
�H���"�2"H �� ��*HȈ�*�,�,�	"�""2 � �"! �" $�
*�
	"*�$�� H(+"�H $��(H��Ȫ��� � ���"�,���+ � �""�H��,� ��*$�# �H+ �  ���"� ��")"���� �H������� "*H"�*
H�,�#  ȠH�"(H�� �"
� H�H�� ��$���O�_�?3;�,�&�~3�\��Խ޲lԭ���ʭ�����\�(&҈�!�c�����`D�ct1B��b�W���s{߯��oU�X��!4�|�ç,�4i��p�T�A M���xFX7y�ߘ�)�xm�^B�Y����[�V�AY���{��&��s��7ZQ ��wd�x�
�]B-[Q�[>�6�s�,Gx�z��En�t*�ҭ9�<�/��mT��F>�۽47��+�1p����a�٣k�[X=��1]����_<䇉|��oCl��i
��	�R�.D_�K��e�y�{w����7�w߾3�<�&nȄ����žj�_W�<���Ⱦ�G�y|�����0�GS�{׿\��G^�Q�m���!a}Szi�B��@%Ҿ��=�f�}���y���/���s�}gxvލ����O!�L�ŋ�2���yDGA3I�г��\D�2�2���!���5�[�=�N�+��ׇ�Eu�No���o�@@ǿ��ؿ�~����,QA���������������_���y�?F�5�<�1l	��>^\DCZO5�wO]�r��;���.׏�aRVz�PyR�u`�f޻��N�ƹ��u˭s��N���xƎ�<��2�:�4Ʈ�:��E��ޭY6gUK�*y��j�N���	er�[y�[Ye��oYZ��G8�^��RWnlǹ��*wr�&����\}y�O^�[hl�Ngx�	� �G]��sm)�嘲�w^���׳VT���	�����m��$ʚ�Tَ�V��H�,�F��wO�x��o u3uK�+�s2�ׄIc[Y�4�O2��ܝ�����Ǻ#n�fL:�6�,�*S�r��{'A֯���ڗOM��ڔ(�yF��sͮ��+
�/%c�T�3��
X�ǝ���n׳<lj��ݚɉ�,B�莄Dj��f����3�`��Y�B6�:��վ��r�3�4���§ ޛP�\��>r�l�w*9ѩ�-�96��'V��PfW�vU�`&��z�J���#�\����Yx��yvZ��e��9�R�$��X�^Ʃ�9/X��ev��aQu�V;m�Y*�l���j76���af�=Ubw[M]��ڊ�^�9�)�d�-"�Q��#t
܁2ȬYC����ø2��Һ���B�p��}���2МN3[F���5�q�2��e��c��R�:PY��l�ʁ41�G4p�Ä8P�Ç8p��
8`��1�`��(`��8p�Ã8pC�+�']�����tÏ��p5�b�����o|OG3%u�N�X�.ych͈,;�����1'X��t��+��7�U�J�M�7���]l��<�]�A��˺�mKV�vnJ��o]zs��V�w	�[�E%�;ͻ��"�4��'e!��~��9)��Zq�X/l����N&IgI��t���V8���*�v���I}����>ګݢ����ReJ]t�Z�N+k3����K���H�n��^��;6����J��J����K7i�㥲�����T�³�0�]K��Y8w&�>����5ob���k����of��{Tڊ�gC�r�㖰�S���Se]^1m�SRL����K�G��r�&��5�RR�<8PC5�滦K][ƫsZ׼q�\������a�>}�oj��s��_�nv�m�yڷ�I���L��v�P�\�:��٪�:u�^P��1L7]m/Ϸ���ͫ��O��Gk�q���L
���ñ��HG����)'��.������B�َޛ}V����6�J��sL��=ِ�l#yY�����w�W���x���`=�:���1خ�aGs�N�S�"�/�'���tF��JWd'�9���"���
�:��%�`��A.��T-GD�w����R���sv��Գ�s�n���9,�l͜hh���Ç8çN�:t����ӧK,�Ν:t�g8p��8p�Ç�Ç:R�$�^�5�v��"pE+q
�,α��9��Utol��z6����몛�v�XҭV�m��6*B�jp���������h���En圆� ���nz�>�\;6��DѶ�`�"��ֈ�j�5�}Rf�̏f:��wf��ש��t�nB��K��8��p��EroG�����A딧[[o���T4#a�2�EeV�>t�*��ZTǨ�Z$��u��j�R��@��xU]�v�K�u���w�����71�U��yb�d����NY��m��[����'��M�F������Dm��0,�.���7
���;���8>;�z�N�J�Av�o$�F��>E���xr��l�F���{\�oT�{j�!.�ou˺���9�ۼ6��?�̈́�@$�J�>$'��9�P9��w�-3;�1�������k0]�̦�G2�d�kt�l��.�V:�6�J�,��|+���v�������ۍ��X%t��k�吺���݋�b��\6�����N=���6%���j�E�8��Ry^�zMݿv��^;�76U�}�ug=ɛ	{��a��̍ �s�zV�Odqӵ���J�Pҭ4�Ӹ	Up�V.�]wpV8�+�3GL�}dV�ꚏg<����Y��r<��걠�<�۽u5U8�%��kn�N�^��ZT����s�>�S�@� F�4p�Ç:t�ӧN�t�t�ӥ�Yg�N�:t�Ç�Ç81Ç8p�ü�2�%�;[��{;�"��3wV�U�� �#�xbU�A�<ᜨ����`nşh'���-4�ҡ�ފӪ��Ē��d�� X� Uq�����:0o)���ufש@ud�Q�׃[��3o�e1ir��c�aŸ㷽xXx�F����Y4���/f]��cFW[�*��v��6E:��;�����[���s�)w|4�F�T�X����]N�Cї�$fuc��sR�%�Sm]�����l�����8�܊���(�6>K�W+}���F];�̨X�G<�ը�t�j3�b/�2����*��h��uB�쫭q7T\�7H����r���»oE]UN��ڤ����U�Yt{q޸$=q��zV��Z�WY9_���9H�wX�":�R-�G���Xî�r��bn��sL�蘹��V(�1-הH&��¶iT�f٬y�X��۝����śY����ߘ˘�B�K��f�%�J�q������ˋǞ \V������G{�i*�U:���U* �A60����^�\K9�U��ު�ú(޶�]�Q���M0�;v��}H��.ؾ��:B�"|�����k��	EV�4�oy��-:��u��+��ҭlV.Z��/5e����5l4J�1$��/=!�M�,
��/Y֫s|��`�2�h�xa��:t�ӡӧN�:t�ӧC�N�,�F�:t�ӧM�:t飧L0`���`��>�q�q�m�'[��.�ˠ��YY]%l�۝�-��n�nCy�Pt��"�g�iu-!Ө�J��cQZ��+�N�Տnh��6wSYEF5c$�~��-��Ck�!Tj�f�r�N�u2�*0��$i�(��5�T/q�Yz%���Ui��l������勄(��֣yݘsqT����'bҘ��뭬��W�t;���2[˛�;�ˑ��|�N��^��w8�s:��Arٰ�c/���+s]6�\^�Kp�\4�F:��ay����8z�#�a+1��'U1��6�Eoh��͛����3uL��Je�wdxLun�ܖtǞ��Ɣw#�g.��:��6��:�.�5pPT)�C�q�VbQh�f|ᘡ+�v��=�U���q�ޘz��*�nf5��M��0A{B�.��sܩ��8��;,��ܝ]A�O�r|�7���1��a����+ٗ3p�j}�YC��q̇�7[W4�SlUQ�ek���k��19�q��buD�jV�;[���a�)Ԫ�]^̞�w6��+8�B��*y.<̆�p�s���-��ם�Y/v֕X����K-IU{3�s2��ܴ��{��X���֙X�US�SU>�T��2��9�������V�נ�ޫS&J8g#�֬�w,@���T淕+�It���^L�[�n�s�u�y/��e��N����!8h��8h�Ç0�ӥ:t�ӧN:C�N�,�E:t�ӧN�:t��N�:t�ӧN�N8p���սN�pw���:Vڭ|BTtq]\juU�K&ˬ�:�A2Ը4LG��}3E�\I�]�_oQ�ج�ϥ	��QͺӋ�░ʨ&� �D"f-�Vl)s8H��.��s�i�Q�t����#�I�p���ULv��v/Scyj���6�1K�ʜ/x�`��e�L�|�u�6��~��m�/\G��ISo8Y���ȭ����oB���]vqZ�K��70�Ɯ� u��N�{�f����������;�6�;�<Z%��z��o'�rR���S��2BM�ں
�"�zގ������g`Z;:�a�\綻Govv�:w-_ei�aT�
3"�Uy�6��),�E��rg
��o�+&����Qs`�9��΅���Ȟ�8*u��E�}�38�Kv76j�����X�k��Qמ�b�TA�xDٽ`��m==�h�7h�8r�����7�ڝ��r�z��^ګべ��-av���Z^�7����ηD9��v��&������.���2�[�����k=��9h��W1�͛�Q�~IDp���QX`D9r�G��f�&C�ٺ�1O�f��쫘��2�\��/�e`�}�ۡև�Cm�<�*^5�4����`K�n`�Ӷ�P�<36Wr��n<#z���{��y���0���C�*��KT��=�Wvv֌��2��f襝ϧ`�#�h��8p�Ä8p�c�8pc��t�E�4C�N�:t�Ӧ!ӧN8p�ÇÇ8^wR�`���w˯Q��:�%;�.�Ƅ�u�Ɨ<́��*:�sl۾�����ٚ��EK7w��}���^_U�]�K��TFrW�GR�������P����Rm�A�\K��$����.OW�����E�}q�dfn�EJ>*T��v�ЏLzl�`�̱m�~n薠7%�W-m���Or(\�O7� xە�;��Ɲ^�R�p�u�1�oM-�۹�m, {#�)V�Fd�v�J�du3t�ݙT`��3��Hp���L�̸ͭ�gW%D������յ���{����`�t-���D`�G���]�.�>�v�I�W��+U&L�{��X-]�<�y�U�i��V�mޚ�޵�|�ӽ.����6�\��p���g`�� �]�:�ܭ���r��aWj�y���;���)� �q*B� ೢfh���7��^����pu���i�M�]�{'S�W�[T�4���'k���v�hM˕l�]�aF�v�4MD8䱈�t�y�Zx����^�SU���Jܚd�՝o,�2[��Q�[3��x��Z���p����;�b9%�8�_n�'�T,��e!G��x/��^a�X�꨺�BV�=��q��Ԗ��V���ݖ����f�������(WW�5�x!L[�5��8�*�\��(��1�#�T�7�Uʥ5��0�R��U|sN)O���k�u6�-v��d�=���U�<έR��Yp�=��+4ec����`�a ��8pC�8`�Çp�Å�4h��ӧN�:t�ӧC�N�:t�Ӈ8P�Ä6ܲ�Ԭ�f���*�]sC
�/s����uh�y��T�vN>���:�v�`��l^�\\�u��f#C5Yu�]�q�(t����,)m������������;��r��>��`�#+��U�uy䬸76 ;�[�-^a��t<*�(+���i^���A��r�Oo/A�H�2n:�ʆn9�-޷DW��w@W-���e�Y��k��d����Z��3&nuw�y4��Ѫw�΅ۛz��>�]��#J'+/�gh�����]�_��)y��5�T7����e�k���U�Q�=w�t6��dv4�+ܼ��JqX�ɪ�*��Ռ��'EK�J�����Hm,�Y���joU^�+9�x:�/HMѱ�0uw�)ְ��j���9���KKw�»3�a8��$�yo����e;���v�<��巁���Mb�J������8کZ�y�����*+���m�ٕ�&a�����J�˗akl��-$�[�ˎ��Ξk���k���i�PE�����:V��f�ة �sj�Z�&���H�rR>ɵ�j[��qJS+f�M��j���;��{7\õ���Ī��|�1:���';��uhvVWU�[���T��Y��M�|�7s_3¬6�t��`�d:L��ks({5�35�K�m���qn���.��r���.әܳ.��.cڙ�h*�k'�M��P"�v������f�^���Ϲ�~�B41�$`���0`���01�:hѣF��N�:t�ӧN�:C�N�8p��G8p��}�;�ds����l�{����T���WoP����y����YZm���{�-f��з:fq.p{�p����8�5��j����If:W�� �>cI�����ҢY�r��&:
���lK��L`n��h��ޮ��;���\�t7ew��i��8�:�ڒ�Yc���d��^��r���f��є�v��:����y;}��վ|�u]���g���m�Y�n���;n�0e���K�Ux깣R�5�2�֡ۆ��xlu�5en��R��(f^��'iǻڨ�%k�,��m��D�ܻ�{[:v>mԹJ�۽}]��X��F��]�Yע�_5��t��[�*��Oe�u�iF��Ov�ٛ��]�a���%U^�����ǥ����RӖ�T�oK��+wS�C++�μ�G�=�u�����'Y�7Y\w'��\V�V77z��G�f�%pFPx�Ҧ
�o��p=
�^
f�+�WS��+��W'���'J�:�u�+���v�]�l��%ߥc͎Yo-U����4�WXv�Z�^����{�'�I'j�b�PL�GkT8;��4��|�8Z���|�;�N�m��gX:�����dW>��}�l���}b��=�n�ZWc�.a�m�{FP�xm_z�]�6�(�x=��t�x��yCRåQb�5[p��iK�NlYݵ���έ�R��U�<�Z��w9�V\fNY�� ��YWsn]��csh�db�ʽ�;q�����s��w%]�c�NVu�ͽ�;�m@U�z�6!��o^�IB��ml�6̾3���*�ԋ.�0�����E�O�Y�=�ι����6�F��f�a�x��9p��k���Q��rn]!��/1�9h��׺���I/m\}���m�e,���WX���+]%[�ѡB�`C��o.������W����TA�N:�p^s��UL�v�����7%V�sQ��6�ֹyt]i~��A��T�k-�̤�ǃ;8�WC�i����{T"-L�Wscw{����I����F�ٴ)	��+]	�d�ym	��R���z%�VR�Vqu*8��{���.��M�T�m8���C������@ڱ���f���si�Gj��!�a�ҫ�;���P9��u��[t�6�9s��4fi��z�ά�3vRM؈�u.ڣ��o���YZ�x�a=�U�vt��:�'K̭zNP�w�|��w�N�D�ś�pPF������/)�\}���j=��Ҕi�]������;6�t���R��䠤]��ް�J���[��IUv�b��6�ȅV�z�(�tI+�כ٪�]��|���sk����AѪ�n��[���պ����4a�p�.�ujq�?g�DAEH��_������~@+�����e����YJ
Һ��jX?��亞B`�,-�0�Ywh�M0�#]���&��pƕvɪ����sl�,&B:f�C@6(5�`���M.f�κ�dB��ZR%��`Р�mYU�y�Yi�ef��(%�	�)v����h7�nc�Y�uca,iuq�Ue0`�4ĤΈݛu�[��k�8��И�B�RPi
��qŵWh�]K�JgXa�
	lȂ4��5#��nW��Fi�e�Fb�U �6�+�k�l�ڳP�xՕ��ث!�6 �n,��[��1�&t[�G�5�$���i���kr�v5�j񌼉��MM�A�*���[�MKβ-m�	�1�t���!q�4�e\�q�a����\�`��-
�lM5��Lc"X1��j����!]��̀��I����f��8�a�c�	j�֕�-��&l9p��ta�K��S8,u�6�f��ũv��f#��;ui
�
�6�%��a:��bf�Z^3ՙѤ�ۦ&����fkE!1hU�mm�;mRh�r�7B�gg^ę`%36�݉�j����m�a��h�b�M��-�J-Z`�-���,�+��
����@Һ䥍�mT#�l�#���Ϋ)5��tҦa�f�6�]2���	��֚,;Q��vًh���U�<V�����l%݊�<��ZX)Zc/XՕ��^ZJ�`�	�]!�.S6Њ��:	Ŏ4�Jcv��Vݎ.$hs�sI�. �2f��&�m�ң����j$W�rf����k��u��GD�d�9����0L���6�-��5�+�v�hYc��iI�U�5��m3gV#�5$9�5uw$F;3Z�hɭ��`q�`B�-��I�%l�f�LJiQ��34�ٶ9v��!*�j�u�Ʌ �%��Ǝ��Ǆ��A�%]��*9�̆�kfت)9Ż=��B�&uj&���M�$J�c����Mo'=R��s��+,��Y�N&���ղ�����m.֋q�-���iIM��&,5�UL�q45�г[1�!+(H�]xr��q�
8��n4�Y��Xetݠ�m+57�Uy&n!H3$Z�.r�L�m=/�UNluZ9�,�Уp7M�Q��xb�6��4[t����Ȭ�`�VW��*��2�شVYiD�Z���io�<xp�n�vFX���a)���M�	ovvhLl�tP.�X�n�n.5�8%���k�]+aA`�.+%�WX6��g���%��FlP��2��Z��X��5�дFԆ
YjZ^.��Ql;G7@Φ�w�|�4�5NL3�9�ؓV���f�Z��=l��э�܅6�5v�1*A��sc\�3MXm�EF.�i�V��\gܵ]�mF�)cv^Qí�%fi,G0j���^ma���\��i������.UeQ�V������hJ85�e��X�J�k��s������xo7�6��у�� c8���ͣ�1���f,Z�t/�R��K13XX�ԗg+�]F!/f���6���î�t�i�6MLcgh�K�iQG]D�,4a��*L���[kn���Xq��l�J�BM�aq=�R�Xf���6k�%uK0ꑥ��\7P��4��8�R�m�Uf�K�iv3���ʡv�%�ً�XU��.�D�f�l�^��� �[c
�s�k�1�-�e��k4���\�lȁV�<F�<2�b�aj%�l�cY��6��j"��1k�la��֎p���K�fw��$���n	���b�D��بWI��H6R.3i�mڇyW�*A����m��V�`�[-�h��k��R7KfԜZ�@�I��&(�)Y���ĢG0M�T���]�d��R��Y�j�x�6-���DɮJ���΄�i�v�U�5�b�6ڱ���{K�a
ᘺ�l�e�uʰ�ַ�B����P�Lh4t\�RV9EhM{.���ǋM��K0ŻM-����ԨYcY�Kv�1CCm��Lus��\Wk��s�D��,���,�mp[)*k� !9�+���i�`�\=,��'�s\��	]�U��`�e�ׂ�&���h��m��6 B�j�{v�Y���
�u(�����	SQ.��ҭ�9`#��r�fjdl��WG���͵%c�g����k-`K�nY��b��X!�-�J:�%�4�+�:��T��m���BQm��	�a�5�æ��J ʮ��KuGY������q�Py����Y��g�T,�H6�5��R��Ħ�!/;q�KWGCP�E�WZ�k�o-��9E	]���[���!���<��e+���v�&�rB�@��	��N%�R��w��tm���5Kڪ�]��*�[2&fP��3��䃣mm`{5�!�!��Y�TZA*aM�{j����"X��u�b�jM�,Le�3R&�CZ!�ă.	�.%e{W�&��A�M+\�\%8�"�t�oP���V��@�4�궥Y�#�;uͥK����:���i�.�٦va�S��r�ɠ�X,��D�\L�[\�� j<�˺\4»n����i���1��1�7f@�v�k:`3^���Ť1�"�&��fz�1�L�34�B�L�iF�v�7�
���SC4�������^���ڻ��^AC76Bت���@��b޷��v.�bT�1A
6�����M+)rSmH<F��Sn�i��
B&��HŅ��P�K�Uq�/D.Ҍ�TFZ�Q�P�����Tme�f�k-dqP"E�!�ڲ�gk�x�J�8�F��3LWL�JҎ�A,���X=c.%\�6�r��\��1�.70�LlN&-H%qF�9��m�Ԅ��<m�Ʊt/-#�vi)�.��։6�v�T�p����\�Z-�Mx��:r�Թ�)�ZgM���`�xn�)6��VcAl�e/1n���H�4PJbi���n1�	�]c)�ڱ&�-n�Z�a��,50�Sl��J��`��:R��m����XMf�l/�a7;3b���S�r�5�[�9Қ`�ۉ������� A�f[�T��˫�eͨ*Y���Qlф.����j\�f��%����Իej�kڻjZ  �֥,J�e���ۜ��eic� �vtΩ�Wʑ�k-t�I��ؖ (%	���[`˛��s��fkmC��kV�%���(۵�Z�F��k���q�Xs��*�.��ܫ��[.Q���1���Z`	x��V���$���PU�kSs-k��YDͦنB���4.�-�k�@n��	c�� :"�сx̶Ǉ5�Ζ�,�T*��^����5jZ���a�		IJ��D��1t����m�4�paZ]u�fU�j��WS�K-7 ��Ѩ�b"�3q6ـ�����Ѱ:˘�*d؛K�`%�:&�p�
Z�Yv66�,�3i4ڷ��͡�9���iv��=ES�����g�L+��]�R�I|�˧�'�&�6ꌬpe�8����cUXس5i��iH�a6
�б�������˛�K+�v!��%5�(�hk��&��u��$MF��B�C
Z��BQ������R�����2�a�j ��A�V�cYt],�b�b�$�,����ݠI��[��f۵ �l-pF���6�M���n�4�#mP��X�۵���e^aPb���e�^�`F�b][	��͕�6��!B.�Y�k�:��+3��P\��.�%�ݒj*�R�֏6�BP����\�Z!yRnr��bRi�^�Wa��q1mʅ�b���!2:;#�\BQ5�y��R�K5���3�)���o M���4�3[A\�6��	��\v�),BU�]���8�a�iY�Z�.j�6T���`r8"1�A�3h�F�]u�m�/,l[��ص�&+�F�\�[��%���y���6	���meˤn����c9�b��&!�
�3n�4[�6ֽ��#Y\Vi��,�MqX�r@#wi6Ů�0EHh Q(��`���KID�E��,Qf �nU(d���y��#�՚9J�M�#�iB���RP�mf���n�F*fĺK��u�& k-��&$֌�(�V؅n(YYecn�&��RO&���:��Č4e�em�b#vc�]1q̫0cl��4hk�׵��]t�i�@�k0Qw$���6[a�a�MH`J.�Q�`G,+i�]!՘�N�m"8皱����l�f����-��Jh-���Qis�a��-VQ���q�[�7=�[�Y�QP����CM���y�E%�&e�U�fǲk	��[�k����eL�Y�kpY�n�� R�̥�ͫ��3��2LD��۬n.�R��`B���Mqr��|��u�0�\��,��j�!�(�K�%���u��Zb�kc
�,mWjVj��*��ʐ��l�f��z��A�@����s�ڵrn��Ky�%�a�!��r)�f����,�d�ni���sq�a����bd`!d6��ejy�3���Dօp�dF��6���.@Q�M.���ef,��R]Z2�.�e].uf1\��\��֕����k5bCL�qGj�f���F��:�k2���1�)sꨭ�TW,ȹ�TU�lZ���qvR7!��8�`uWX\�s
�b���K	t�mKL��ve֛�1���cX
���%$�����1��cy?���_��c�/QGo-?��y<���hg��w�Sů���y�V��P��r�t���X�6�;l��%�׎	Ia -&�E��#l�si`�b�l<rsS�f�7���r����Ʉ�<?�t�����B^m�w˛e�	x����	1���@�9�S�.qD��XF�=:tθ(r7L׼��UF���x⪇��^D͎�";���w&Ǉ�<:H�n�rNWS���)�ͥ�mnC�y���J��'��H�'����m�q��!��ç��N��Y�G����(�-`�!�	yI�
��L����-����Tw��\E���N<�qм�$��4l�Ä�˅J2�xj�XB�ɧh��[��*F��/�N%�����9�jrn;I ֢���y�L�Z!j�%��U�XS��m�tÑ%Q�OON����l1��u�q��0�N�I{�M�:JHa0X�'L!ͳ;�Ϊ�	���i��U@��l�-C��It�2mhbgI�ȵ���� x�v؏N�����ųa�uu��a�N��N�1�Iٲ�0A�z̻?+�D�wx�K�����ؚ�L(�1�B�2���G���=�ۖM��F�p���	%B�T%sI���	!)���)�p8wd|���byU;a�i ����ho�sa��^�_/7�z�p���@z�����V]�,Lڝ`Km|�Z�yB���8���)� ���y�ӻ���ߕ��Y��W	��*���3�f�\�f�d�;EҸ�Z44h�L��J7Z�n�T�Û�v�ԳKR�KΤj�"��!,�ĦԚ�͚X]	ZZc��O�b�ګC�6���L�;��-�j����*�ʦ�=D�`kf����cV�K��1�u�
�+�L̯2��є��M�6�F��M5�T,�(��Њ١Bu+pma�����#�&�S`��X5�K�
4�ы�]6��
��U�M#	�3Bk�e���ڛ5�Kk2���c��(U3Qb]��W��,�7+��v��7ux����3Mnti���P�)Eơ�@b�4顕������jd�l,����[��д6m�:��a�u�\2��_��V����d�ݡ�aB��;$.MM`k���j2:��g�y-��nG5���5�n�6������h��%��� m16.e؛�qU��<gXцؽN\�ՀM��Z虳V\�Le�8�,������
J��M�#Yu�!u�x����"�J�E�9�Z#�L�SB6md#F����l,�eM,Y�\R�6a�����l��,�����N�����Cb���2�YD�ۚSe��0C5uX�kar#61�T&m��[	m2��ʗFĎ���ٴ��"ͫ�f���j�{-IB�N���jMi����)���7u��ږ��b��6��9�G�u�X+]-sH�vXkX�Vӛ�:8�p�MK��4��Հ��DƷ����+���%����M�v���5�KpFf���S5�&V��dմ%
� �FX�0�Y��4�\V�BQ�CJ84*�*i�S\�1�`Ѵ53j�^�!���m�Hb�u,�Ĳ�14Z��F� �PxPnkQ&a�����6V��Q�؅�y�(�oӻ�'w2;��AT��@��k:���IJ���j���Sk��}fX�,T���jŨ�،�I�vE��V�ͳA�5ZV5�l��'F�t�����)�#� F��Є�	N�:�&�mL��&�:d�ym�D*�������ڜp����T`5-�m4������;0��Q�$�::�k3l��2��ZL� �-�-�V��g�J���X*fQ�Z� ����؟��?����$�+��˳�v�Ol�LnЀ������1wO��^��:p^���O5-���I����nJ��=$g��<?]�p���t%���75_�y��ܕ�"I���Y(p���Y~Z*gl��qI�V��rX�';9J��ld�^'�E�v�ߝVdi��n��{2�Y�f�g��^����ڿh>;�_ʞ������=���-���!�M�����KFP�$+�Ȉ��8Q0�0F*�AT��r�0)�n4\_�^{���د_��aŁ7��t�����;��[B�n!%����ev���t5Vb#y��sON�L[����7�j�������;s�.ܻޗi+�[^J�D�կ�{��j�L嗯����� �Ib�n�Jj��Y�wݢ�������o'	�/���B�T�SV��,�>	=Y$̓��zѯi����� *��ɍ�
w�F����8@fׁ7,X;�Dk�E�%	#��k�^+��B�4�_��9>��B&���wZ����Ǧq�#;��{�����҉KT��P���R��̰�U �Y�-���IQ�}�\����*��b��n�q��oa�3�χOZSqZM<�����ѻ{�wl��No�vB#C=�����f;��#D]��0���To\M�Q?/}��'�7wuH�᧺*��Nۅ:�f�E�şA����\Σ��L�ӱ�cJ���n��1Ӆ s�Or�W�� ���8���q)�ٮ�{��|�*�}#����%�J��2]�3�0��ڣ+0�92��:��@U!�+=�^F�Bj�Th��Miyt��3���75�Zރ�;�v����y�fi����؍��%ޛ��W~p���"���\aټ�Q>�e��꩖ D8H����B���ܺjXR�eu26�)��B(�`�h�P��X����}T��v��t�'�^�����+�n���I.�I��i`.ﯩ,_g���ڲ�hǱ��݈MUɯo��
�
T0v^�D�~�oز�F�_XI�IH�yz���F1+��Z�w8���sp��x-���2�I0pc&�S�N�B�ӵ�zv��9�z�VUU*�3b�T���yFHR�-�*�[�rDF�;�q��MF]��k^|>�0� �R*־��aJ�;�S�2Ijme9m�������p"B��G�͡u�\)�&T�9H-$U`����*V��=Z�"Ya���2����cp��/�A>��-:	B([�!fŹl�X��[��C;,���[�I�|�o��?!���@L�����Z�������/r���
�}2��S(\�om��,n�w}���r9S��7�G^����ڇ�-B}@h�>��[���_uPE؝�ywWP����&~Be�%�b�Fח���µ|�*W����&30NƷn���~�����[mމ�[�T��S(J�T�P��
�	���ʭ�߱Hg�\��t�з_n�^IG>���	;�ܧmˮ���-�ӯ7�X��t`�$�]v
�a��b�#�c9�����I'�3�K鮶���LRux�W��o}����d�4�6��݉$��bo3Uڪ%�\��6h����E�cf�ؑKh,�Fk�J�cjb�"���
B��r�J:���Y�n]ٮ���T.IBke�8��^��L�J��<���Lس��;jb#�:�6HF�5a[�]�7VZ2�W ���Y���::����0c]�lV�lsG �"i��QB4��l\�m�&�3e��9��J��l[~a����R_�%��Mu����Q�ٲ�عr���@�����<�C��HJЪ_
����ۭy�e��7զ����l
�u��|MT?E���� �r7�}Z�E�ܱ;������^O��&��Vi�!�˨f�mx7E�}׺GV���;8e.�����qKX�l�"$�IU�;�|f$����2�|�Ry�Z�-B�}��D/���ϗ�W��ŷ^yI�o������րt�ܱ�'w�X��'b��҄��f�^����6���In�ĸ���l0mٺ�N����0�J6��n�jL+����?r�)��i�n���������S�����{�	*eL��ߧ^,$�)��0����Vg��b:I��W��9�T����wvJ���ZkfXfʝ1��5{<�ʇ>��!����F�}�ۗ�?���4��C:W*N��V��,��������/��|����^ �A��H��W�V��1}W�׬Nݹn=Z.N�AR�"����A�&�
��[��a��zo��I�m�c~�s��aUξ�P~tt<����\�>�z1��.�Y�vqB�~30A��R�Ij����}�1����ڗkZU�(�v����1l7kP����U�r�Fx,����t&|3�B}�]���YC��KG.�9zI9����OL�N��ܷ7 ��g�~x��'�m�cf|�y�k�
���t/��<�7A��"'�+)i��7�u�$4���?Ms��7��vU�F=w�~�R�؋9�u��S\�u�o2��	[˧p=��3-Ri��"l�~d	"���UY�@��Vj��Ʒt��9�Vϼ��n�P3�.���l��u �MG;w���O2|5��:9��J���4s��A�m�-������j����:}��;������U6���L�w>ڟ^��T�?����2�K�� �6rf5�%K`�e��f#t[�)�0�P$�<��@L�������8�Fn��F2B�뭍ʨ��2R�I&0D�5�����sT;l?��&2��eiP�\�r�o�/����$����ݻ�.�օ�+�3� ]ȸ�ts���Q��#�H;v���j��[t�a.G��:F|6��<�-�Rۜ�qO׺vq�@p�5�A+�����++1����Ii	*�M(MwKM!��n�Y~5�+�r��0��A=��0�0�Y�J�쫹�Z2���f�y[�l�yxGA��u��X�wk�h��l��<㛼�}>9V��p�;h'M��S��M��(lU���H�	��4����4���������`�l@�*	�҆�,�Am
ݪ�Y�r���ڡ�j&E�ɭ���X"�^��ʙ_L��#g��W�!f���Q�sN�#Ah�c侙��bG�`F�g���&�"��TJ�
��5J�7�p�д���sq[��D�������HI@6��3S��=B�t������=w~�x���S������b$ޙ��L/��}��+���I���ĺ7�����_M9�S����/�����!��gg+T���'��6Y�Gh}}�+�ۢ��Z1G^Ծ��^�h�Y��ͧ�5WR"Y�5>5T[��>���FȲ̑~D�,�e� h-F�#Y�ͳ�H^G#rl�P�A��3ctX�ܳ	,���n��ռ�[�����ݩc��������ڐol-�ik���B�H�v�E��XiMp0��[*���Gln�6��mcAэK5��.���`ұlq+��Qr7 �+�1Ɋ2�:�3����k��I�߬�a�%,�x�X�\�!c�2r�K��1[h� �|��},��BfғY�Q�����&����#Fڳ0��D&�.�&P�Y�1;�+|TMh�?o}�.����wm�%�|&��wEfC6��_i�w7�ܠ�m$��7+���~�Yr��m!l�##��5U$^c�b����ݘ2��<��|k�A��y��6j����֯VvM��#u����j8��`�a��Ӹ~�X鸒��d�U��FW�%`"J���܊w\�i�3s�}��I1�{���R�e}3w��V?-Q,�2s�4���<��i���p�+�SJ�勫�33A3�fe��{��}Z�T���wOv�{�§fvgs&U]������}O>!wY�[w0nn�խZ����hl"�՗�sF^U�ܛ2�-�˽ĳS���+��tߣ"���m���7N�c"���n��ɍ��ߙ�;�	�o�:�����j����O+���y��u��(��Tܢ���U�(:I��nW�Xn�򽁻�?)q�󵣲�c�����+ӹЇv�mo��)0�S&�])��}�>��ʒ��!�!��W�a���3�ck2`m�C��tt��Bg�J~��!x=/����^�i��#Ɨ%�se������D�G���c�u�ڟ'�_���0)O+�������Wܠ�MI��p[�KD���H�=g):������*j��us�e�/�2�hE�=�Y�G׉o��eO�A��f��(���(?n�B>�_L�}�����֛�ra���
�I��9�U^�ټ�����T�]veJ���b�ꗏ8̕)3��P=��N��ͪ�ߦVB�>����+�YQNwJӭ��v+�Q4V*�'a�׃{����y鸢q
X8��I.����x$/o��Ρq��S/[�v�qi�gQ:����Tv���]d�ݹQ}&�<;�SL��9G:ɫ���qWv]�P�d�}݂�նz�U^��Gna{t��m�t�3\-��+lw*�v:Ir����syͫr���Yy%�Y�+�S9�k�p}|��so���f�{�w�-��7��4zf7��D7�PӸAlʪr��[�'J��짻�J��Uwk���[�xq�7h�\���5�7Eޡ�]s)�rĦ�h��A�n.�/y��0߆ē�X�
o,��\�赶b+lcYtD�!l�㯦���꘻�[��,A�0Y�_p�ʸ�cocd_vN7�(\�7f�Z"bm'���sU�|R�r#2���:�W*,,�,o�qV��Rq��Hd���+���q������n0�!����ˮwZK:٤=��śA1�����;��GefU���z��S�
�!��p=��ݜB4ƃ�����蹐c�hۆµ;8m&6��f�h�쮖T���׷y;�����sU<�|���ҧn捵SnC��.�Ec�/7&^`F��Sʔ`�ά�TR�v�3��e�nڱ�M��V�<!�K�x^`���z6������=�b�M�<x��O%u���8�=���ϷzK��/�Z޻�s�/]��˱`�#������>��vӫ�OBx���f���\|s�s�4�8�<��y�q�!�7��
�?2� $�[�qʟ�yG5�od��O��c�p�bk�p��s��$����4�V�Fr�5L]���[�g�x\�>�N�������U�X�M}��.ng���."v�%��j�����0D�䒄oVS��>�N��q{uG�{��́�<g	{�:�@um���8�6/9�K\�\�O�:|>���mfx�b���ǔ�M!#�ͩ$��I�5Vl�1J� Ӈ�N����䘲�?����1��BC{\�Asv>$8�ja�\^0���p�S������|g��nl6.X��jjj���D�Ύ�'�p�$�d��,�J�֥��q~�91����t�)Ѫ�7�P8x����4��Qث0n6nh��l�����k$GE�g�űs��������KtݧT�TGr�\��g���c��*�\5�"+��C�bF%�"��-���o&[�=�(iJC�A9��tRL�Y͛v*�#bEʱ��$��! 'ϙ5��<�2j���>U�ϝ�����fe3(,�e_57Zgc�2��N)@�/XT����w^<�����j/��À7��#�%�T�w�T�����i��\y�
��B���w�k�{(��àU��޽����/+���8@uSU/�T�޺v��߹����}������!vLڲ��CKq�Gv�T�M,�R���є[Ts~������Z�)���O�@&�gL*�و=f�+�1. {��8�L�[�v��|A��P�i���'9anfh�L�.Q,�{����}H`/!_�/�hͼy����_��!�F�@��}v��yZ^��`����*S�`�����q����P�����w��ھ����y���n�E��9tN�Vyk3,9������ո�;(/F�Y�-��L�T�ױ*�9z8�|���;�}_ ��{���Ԋuy�e-�mR3$���.AZ���9V#�<>�d��߈�W!9�6Ս�(��9�Wbm���X}+Ȳ�g�W�)�����=�#ĀH'ê��=�E���/��m̠��s,��8| {��C<|�� H�<7�kķ6��^�kA�_n��� R� �>`z����fH��;i�Sd�-�v��W�����6�uc����6����}��/z(�@�;f�7l	�vr.�]�^W��>b�C�d�:=>T��8�����©|��_�I�|"}[�����ϥ}"��r���+o\��iw��Nb�'�`�T��괝�_�-�o�&l��ݑ';E�Q�c�O3-����I�,@���_w��C���Z�A3��^Z\�*�|�����y�>r^]rB�<��@7L38� ���܅���{<��}���#�2-��������!	#ؾ��?���P~I�~�3�R�p��\N����˔���W����].�ƾ��Hq_��=AP,6�a���\h�c�Nb|3��4��쯟�V�����ӻ�{�D6�t�#W��5,�hVE�N���3]�2�î��Je{(�Z��V�"�
��4�κ�c�<�4Eɣ�@�!u�e��ܗM%��TU�[��bX����5�e%0��mԣD��J�Vʒ����E�S
F�-�fkȟ0��{J�v��ı���b��	@�pݤ6(��)in�;b%)j�:[-��)e�,ڦ�&��TR��x6�+ZiF�[QrD�h�:+��5�9�u��sv�qc-TU������Rk,���]�;���]���H�Z�4�V��
�q�[��}����@�@x���"����W��v���;��k��;�.�l�p!{�- ��� �%zȒ�����>�R�W��@��	�=�=u��y���͆8��`j�`J���g��;�������W�VO��\��`����*�<�����P��û�b"}���~�@0A�a�~�A�ES��3)��s�9np�$Z9	�Q�o� ������_9��#���p�g�� �����xj�Q���ݝ���;����(̧D̠�L�0������|72+�êv�яz��]��}MߡtC[�D�r�Ӝ������ED�!��0� �-H�m�r��.	���0�T�L��C����^�����?U&@��]�U�h]�q	ϲ�b\@ܵ���d�|�F�jT��^~�@wJ�[�j^܂7�q��(ĥQ �7�J�r);J۪������6��[��	���yS�+rIهq��11;�i<s� H���T�v3M^G��4�\��}��A����5K���t���b �� ɶ��/�5h2��j�`�ESF�Xz��c����k���� �w���Ly �S�TàBT� R��:�z��\  �68����A$�X�ً�d��ݖ�9�_K� ���`���s���G�G��Ҁ5�E��?��H3��� ����ȠN��wޥ�'�cJ��p�es�#�_p���?��ި]�۱l�g���Ϯ�jO��J�� ʷf7X�Q�u.hۑ��b�jͥK���Z�Z�� �5LgM[\�v�3~���U�)+�~w�?	����e�9�K'9R9�n��cum�P���Y�86��y1�d��}O!��_K��� �?�R�{UG{Vı��_X���@2+�2*��S���ωk΍Þ^�����>T.1Y��^z�VIv�Tʳ׸t378�
�f.�U�iDr��e].�X%�5k�jؑ&�ي��]0t|�� /���1�����_W��㊼7k�%X *��|I���x���7�`��� ���սegWsQ�s;�/�ЄG�=�ز�wh����k���uH ��� �?��^����f�_�X�����5{�_Td5>��x� �T�� �����JWEPУj�:�,�&���L����ᱩ��Ks7U\�&��\�V��	kA���*���ER��Uy�滪hD]�,_5��k�x������}��ӪD A���|�R�o�gL︽wYї�8o�ԇ�m��5��Y���d��_?�y��.���w��$��׎y�K+���3���U?��_0@F�w�zL��7���TGny��j� Bw�\#�Zs�l��,�}���ρ��Ts�>14��],0GL� �B���<���wTЈ��X��/ɐ/u��|h%����wJ�"�k��f��ΆJ�s	f�1m��E."������V����`���T��sm;�'hI/X�s8��F��_�����A�NĆ.ׁG��h?������˃x)�8ͥ��ͮ� �p�3'҇�H
��ES�kh�ŵ���l��Qup\�4fe�F�^qh�WWmh+���B*�h�Z����ʯ�M{V�;is��!"����w�ͩ��*2�b\�s�5ޖ�1���A�p������&�@\ wW��ţ>��G�"|���6�����w��k���E�����~_}v��Q_:f��jh�Q��>]=�I�y�!r�����?U0#NIgb�y��[������d#�(�G���xr]��--�Y��;�DT�`�~�	��~I�؛w�ͩ�Ɉy�1+��A�3\�u���l�p��y�%T|���+7o��}���y�_b���{N+��s]�!]��X��oɂ��_0j�8�gqu&z�WS�^���h�d,�g""��i5�"�Is�����x��7���n��ffP/"��tV+��w�nN|�z�yVz��s 1r�/l�v�O���'���TCvٖ��a-��A��M��H����ݴ{%��v��P��R�2�@!p�
����0�u[��iq3m��lMm�
[+-�k��M��Ɛ�ͩ�2��KpG���1s�,:4ã��X�{iβ�˅��q°%Yn��^��q	mݴrXs.�I�M�����c�&IKp�ݠְѣ��6�K3����U�J|������2���%�y�� r�L�����
+"�e��jQm��'���PF��U!悪t(/^�9���w#3�����zT����$��m���>
�}����4�E�v|,����P�V=����d��gK����#1�����̕�=P��o�`��`���H0���K�yd��vJ^�����mWs�|����?���@ݯ5I�a
� �W�ck7���`�Z�b���ܚw����0E�}�.�'��D��ףt	��v���x�MR`���W��c���� ]���_15O{y5/�Vz3�%��u�ڠ�}%�I`�J���/�:5���[��"uw2盱�면pmfZg �E�Jۅ%�A&P�.�Гs�?��v�dU/�R�{����gbgL+�j������{�q�S�&��#�U�����{uW���B|g��y],�0�����Յ����nr��6���ޖ��]i'�Ȍ��p=V��b���8�����m���=�8���;>P׼vn���]V&z�"�]��K���g�-�Nv�����ʺ��^x�g|)w��j�!`.�؆l��_}����
���A?*�$��) A�}��:`DjY�w�wͩY�+�χj�!�������̢�fPYh\��а��Z���;���1�U�u#�e�7~勁�^_�Tn����O�@'+C��!���s���l?�R:<;��>����r:�]�k6{�F.��_��
t,�%%|��u�*V���!��=V�K|0O�І�fE�.�k�˗]h��٦Z�۳Tԋ��+��~;�!�L�����j��W��ەي����Wu����[	�)����SA�A�a�P�H2��=妇۾�F�F����cx�~�x]��/Bs~�����fW6���g�g̦��I��B�ǜ���%YYg�ޤ-��9��JQ�s1�OW��%L)"�%UA,Ɍ��z�o]Z9"�5OY?hj�����s��uW�����4ӥ.�D�5�������BB�;o�ߑy�\�<���R��>� ����*���1�R�!>�uY����kl�.����� ����^gsnV�*�^�J�pYH;������^�F���A��>U0Ȫ� �u���ߜ���[܍����W�X��5�� ݿ�@J���*�=y3�Q�v��[�ϸ�ϳ0���u�b6��6)M�M�ѵZ3lӪ�6�)��kAr�׬1!RA��
�/�N���Ց*}��.ce��f��o��2���">
��`��(aJ�A�*�{�����ϵ?�����"U�r��vb�E�ĸ�J��#�c�E!��9]����� �DGʘT��<O���p�G�G�L���+"����Ô��Ln_�Z��0E�����}^���HA��gPpUL>��z�Gurȕ>���|�4�Xb>:�ϊ٥1EV�vẀNS)d�)�J?��w�U��)�t�K�U+R�5u�v���'w
s.�*!~p,�?`��~�H{MD�Z%a(�����=%}�əVBL�.0�-�s��|�*���W`�v�K;Y�5幊}�*�a&��a�����6�s�L�����pa%�t$u^I
"��J_&؋��Ѽ���͡��s7W*���\��	�_^�>����<:�`��Do�/x�����{�+�X����4����F�H���|��0�B�T��5��gPd��e>Ŏ;��ED�wԻ�	��ȪC�.�
�3�~��?���Q�ƦK��i3�R�~�U�=��gi�k�3�/�*�g|��L�9�-�9�/�Ip�Y~@�-��}Z�d��27[�� Y�r#7��=I_�b�	�&�>���y��߬XU)�5�K��T�)!�Rn�����+X`D־Վ7��ED�wԗ��-�U1b>Ȁ�ً���>� ��m�w��:�^�6!_�E5�[���6��Y[�^eb�x��U�q]=t�t�u����-H���tz^Z���E�V�Y��W1�K��p��d�`�X]DL��)c�)׆y �5�,k�}t��ɷF���U�Y���z��)]
��\c���KB�l��j^eG���Z9si�~�zZ7�{5ff</�u\�cҮ�t�2�=��FkU�{F���R�e醦en��#XU2}���ܬJ�|y3���	u\����C;�;����ʹ������Z�����3#�v��̱3.���|7����:*�5�н�5���Z�@�x�
c�����\��?vn��G+��Ȟ!�wc����׽<{�ӝjF��*9���;��yw�%s���R�nҮ�
��Ї�-_]fi�F�n�;1-�p�ft����7l���uXUT-"R���\(���>������kq�o��/-������;���r�{9]x��N*s�B�r�Ǯ�P�]v�y�����u#�gE�14�B7�;�5w�^Q����#2�]Z�ͩW�[w*�3�j��l#�7g"���u�mtQ]��������V9�K�x�v��.`�͗�3oWU`����;�6�mT�t��)�K��.^uJ*[9ؐwR����UU�5V���7�R�6PF��jUK*Ɗ�K�o�y�Y!N@��MV��`ZC�8L��i�I,���<��խo\��u�Rj^��r�Xt�K��(J���=�2����];,�R]�A�(���d�k2�*���M�}�����ɥ��h*���yesl�@�Gh������޽Q����<�ҁ[�YI�LiD"7<u�3ˆ�^���Ͽl�Q&�W!>6ӊ��7wSP��K.H�3��L���������zw:��$�A�ibﭙm����_�Wn9��k* ̤�&Ů�˂��8K�'�xxyT����
.,����j9�V������[��#y+Q�û���)�,EΫL��RQz}>�;�I�[d�뚺KĶ��"R��Ò�f���j��/xJ�oP$H�(iC��s�H��W%�ܳG�Dx~?���S$\�,d\�3\��QBMdU\\W1��ц�f%W���#�jBb�HG�[	����xt�8w@�>��8��55�X���M�w!Ʀ|[��RW"�<;#c+z��L��u	�8�ç��Ӹ���
�*,��L���Y�Yb�R+AVKg4��1�6��+,�f�s���N�#��W��\k>���c?7�
BV�݉hӘpU¶��Dض�p�Q*Ԃ��"Gj�i�H���x|;����]�����!�9�Nq�ret��\�RR)��I٥�Z�v6s��S%R�j⋚��r㼍mJ�~���b*��DψZ���3�wl-u�H`=������`�
,5k��. pfbm��($��x��-mWL)f�[H���:1�׫-�t1e�Z������\:�p�b2��rԺ���ظb��`R����ZƧR��-ۘv]#y��8у�c�at�&�]^�L��j��k�Æ�s�.Iy�i�)�bX]�
6�+tr:�]K�\�	���G*�k�(۰�1���Wh���iKX�]) C����
җ(�Q.qF\�@�,���L�,qZ�ئ�v��y���͢Zh���0�[R͝��+(ɥ�k�%���Qn��%arSL�e��\�'8Z�ƒ�F]Fl�Y�[5�hMS-�I�˻c,p �Hk<ct��d��G�<�h,���1��aw:�s-�A.��%��%�K+�Lf��룊��ὬRYkn�ke�I�����m��v�p��l�hX�m��8!h�ݥA+-�U�eL](js2���\9HƼф�3�dsB�͌m�m���V��,�E�n�;�[°;9�@�e�u�Q(�Y���v�f[c�(CZ��n��%`:�J��6�P�؎҅P�3m�͙	KdK�;Y������[����d��I�Rb�tc�`�hL,�t65�{u�c 
sxjF����::i��X��<�i����@oi1E�Y1��%y�.he�%)C��h]!a��.�U�u�1�n#3��J�S�Lۣk6��l�a�8�.�6�j����̮T�Pm�.����F)5����-�+�K
��@YiM�-v���j���XYté�u�n��Zv��격qj.����^�����I���뤦�!\��.èE�jѱ��Z�,�Kl�aUРE��	�4ui
��/Zh��@)�_<�4�&�M��fj�h�1���e��b���(��HݠBmsu�5�;h�n{4��A�;�c0Q�X�"4weI�7,s�م.��a�����k�_��	DVBHAa $'w�;��m7zxumsL�hj��Lʖk[.W)]V�$4f�jF�!5�R��q��[L!,ys��T��K�H��	q��ՠ�%���Tư��Dn���B�5̺V�j��4���,K@���h�YC��vSL;�Y�(�-U�V�v�`�KCm��EKv/k�ke(ʱElsX�ٙ��7z���1)]vt+��L�hՆ������գj��L��j�աln
�-��#�VT��[k`�Pb�0�H���>��ְ*���I��3y���.�S�� l;3�����ʣ�	�_�>Q���4f��^�Y'7D������H(ٝ�?�������"3x�Ԗ{�.��ɂ�q�A�O��Eo��C��'�Z���A�@�a��R�lt�7ѡ�'�粝�S������� !U W�ު4�PI�%�*զA�1������<��g.o�s�/A�����@o�>��R8��y��
9�Ð��0H�_:�����Vq���/N�Kh1���'���%�勁�W�+ǥ*J"1�م/� ��0oDP@���I�"�$��E��ڈ�-F�B��k�����M8$��A&������e
�ٌ23و\t�9o}���9w�R�"�+��ۊ���ER!M�?A�
�`A�L`C��l[(���}�pN:���$��͸s!W��2Ί���Zӎ�Ƕ�އ<P�ә,ap�����in����X���1; �`�< ��0�"�! a!!@R|�I�*���Xoﻜ��}�sz�1W���]�`�rPdx��Ju��	���c~�a��BI�4����R�z~Ѩ��ml���i�q3��b�A|�`� �k�^ �Š��?0���=B9C~ ��}��H7l1��|w{���Rﾥ��27^\�;��G|F���6���&&�T��E;.�y>�~1�����;��vb�E�ؗ��8��"��S�D�Ӑ=$�F놷	\�mcL�FLifpR.V���21�v�K�Ů���|���t��հ�v�!�]�'9E��܅�ˠ���sܱ}�Ga���y�{��HFs�\�)�s��9�[�M�ϝ�^j��8V� �6v�kɞf痕�Թ�~@�J`�B��]���� {�۴�A;�f��%�RU�A���h�'m��S�]5_�	Y�n=C��a�����b�ZP��Q�ܽC�+�N��l�-�%q�5"j�����wڬ�U���2^�8}T�AD0
"�"	(B��"(~�U�t?G�^��~���_�)A�a�*� �1UHa����t_�wP�{P߈�/�5H^����d8�{V.��'ɑ�Gn�r��&((� M��a�l0hэ�U}�>塋��������y��#��p`�2YH
�|� R�2gٚV4'����s�m��F]s��ʐr�c(9؛�t�J��t���?������?���7�;��v]?E��.I�K��(+(� ����g���e��(�Q��%���9ﻻn��~"<�|��7�[Yۮ��G��T�!&ȏ���^j��a�|�⦞��0�|��b 4|Y����s&x��7wP<��͈�&/~���2X ��O�� H4��</�u���%�e�_l�!�����Lݮ��Gp^����z(�i�B>#�_:Y ��}}��������$�X�2������1�7�wuw ѫ8�\�rT���H��]��2��t�z����3������","�B�"����@{v�=����ES��f�f�B�߫�j�_���Qjb��!���ѷ�:!���9�X��F�|��� %i��Rݍ��"�}<̪
��E}z�=�C�s
Kwn�um���LL��F���f���5	]*�}}����8�=ydЇ߷�R�L_��5-ș���oֹ����+�ל��#������Rdj� �x��>��'�T� ��`f���z#��� N��*�1 ٳ�����;Byp>�,�v�"�|�*"/�*�����f��bG�	���!<�\!�[�U�W�ʿJ;�zx�9��Z"Xfm@0l��߇�\�F�{�|_}k� ǐ��q���{�����h�G}���w�m&e6Lʸ�8��Ff�;��� ���G�"6�F�Dwfn��*��'�(��3��a�g�&e�a�n�w:
}*����=��J�a��1��PX�z�;9ݼ����z,�<�#u�Y�f�ˋO��{��3�U{�P����c��3e��I�)��m��EMR}D~�A�aXE�DaU�Y��[�J�.Uٚe�m\��4�*���`ql`n&β�v1U6X��\eQ��u�3K�#��Z`�1�8!0�Z�D�W)	���1�7*&`D46�¶ �k�[�4S:1���HѲ�X�9�F�M.i��-��AU�KV�f�h-f�ep�F�&����L��Z�l�cCa�K�MJL٩v�rĳF�7�i������6X�,��)������������s�f�Tk��rTv�_�ע��<#,�}�Ċ��B�����#c;�C�O�勾"�z�c�F��Ղ+!���>(T��<l�v��C�X:.��V\F����u����ջ3������HqB�|AX�'�I���@�����WW��`"�>����%rK�Sa?���{��Z�fn��%C�|���.rrY�_���m��&@�ݱ`����j�!{�#wݰ��O��Á�/�\mi�ݣ�Z�Aq2$RL ~5H?��P|hѥ�K:�^-�80N���Vw��D�_��!��U Ȫ_:TE9�������ػ���?.��#��2�P�
rڦ�4�+j䴕]ۛ�����}�C��YG�!�0~�C����<}�<��h~��9� ��ŗ��d�P�P4����-��[�\߲�����T9(u�ىuRD�AF��I���\א�.<��\%��{))��D[�m��ߜy��0��FL�"�,�#�V���� �AVQ�Pa XEA���;�~�+��|�w_;���\zx��V��(��!���`ݬ皧��^ڋ+�	�?x1�����Ѣ��7Фc>�q^ذ������o����Y���TJ�r�+��s�d%n|�ߛ�|̮B�3�e�9j����{�"7yތK�#�|����^+�YV��1�k�;�>Ak.�]��5L2*�Z���3�]����V���p�/ޞ''�V��g��T�`�&A5J����ʑ��H/G�J-�n57Z��!v�#a�����Y���Fc]ma�AQ�~��. �r��0��a��A�A�a���hX�������ع�#�K��eK@NcV�@���v���cB{�o�r��V 3���݃�y�9D>Þw����@;��Bg���{�2�9|��a�T݂�-6������*��G�����9KVU{ˆ�^��I�t�;_6���*�~��BM}��f}�00��7�f2�Ƀ�� D�PAQ�Da@�\��w��/�o�d��W�I���4f[s��ޒw�_������J�G{�z�����(@#�}���H;���%�}\=�LO}�����[��폳��;������A%zÖ=%-�ɱ�O�S�zgf���y�K�'e}@����@U!��k�^I\;����������|�2=�JG7����8�X��ǬM-C F3f�`�wVe�c��?Bc��<${��eS!v�cvuf�:�p�zx��9�����E��.d���Z�ݯ�mO��"t���}?n�D�6g3����p��8�����	N�� �Z�f���?e�=~���ܘ��o���KS�������_?�R��-��M��N�!�'ky��W� ϛ���-'9E����{�@�>c�|�Or����`���T���Y��=�''U����0F���8^�ķ�����w��FJ7�T��5Ĥ�vj�b��-a}Ø�#g#������z-�I�Rȳ9x�G���DV�@aXD �QE�Tyo��d$���!�O�8 ��d]���Ssߘ���XdԳ���X
XcE����bٮ�&'���qP���A!~>��c���a�������;����eІu�s�sk�yU��0AJ�4s��nB,C�؈
���%2��H�ƚ��2���/^�K��˚�ky�+�<妙#��F$�+�.1�C�*��Eܿ�ԃ �����*\�� ���so�/7Vo�MG?H�������/�d�g�~�en+���[�(m� �� �Sa��A`��Sʎ׀���>���c�jjǷ	��!��j�dU7�R����޺[b�J4 �VC�Φ ����̽{�D>Ë��
�|���,�x<<<P�<��GO��<�I�E�
L0ET#��f_���(�M]��v�~��'���ϗ��J�`�� �puaሙ�"Q��?e���t�h�ٔ�p[^��LڱC+.�)������k6��g;���d��k33gT��]CJ���̙�>pC������X�ENO�+�jꋫ*}DH�0�	���"�B$ �B*	�op����A�J���v"�mKft%�!6?v�
�֜x5��=FT�͉���l� �S9��J�at�5��-�U�ي�-�m���d6��a��Y��ld���$e��5�eѩ��3��1f�FU�i��ga�Ú˃
V+)iv�0��B���2��Q�sDIe ��͆%��.���IC(`�Ma2�k4��3h0H���?_ԟ�+�R\],3&�pkQ�&� ���p��f%h�ծ����y`��C� �/X`���U1�������nߵw�D�Ψy׵6Uv�o+�;Z-�̢�fU�!9ʲ�~M����[��Z�A�H?�F��׼DC�8�}�.�w�?�7l?��\�/,>�������DT�M� � ݡ��ߡn�F�{�*)ϯF?P��V�������*�&J�0����>��o�fϐ���,b>(�n�cz��������c��� |��"���\i6ςm�f�0~�M �"�S=�����	����n�q�8�|0�/��w�F��cە��KF��׸_��__pIXF2hf�,�xջ�I�s�f�t\ ����(M��nDh�gC��	�:�`��� J���n=�����5Z�P3��f1��2��sj#���^�(�1�m����vKs^�It�SK��?~�n����vk��km���a/L��W���RF(�`h��R��;�\h�M͊���v��v ���-*�Vn�~��PO�PA�HD�AaM�h��"�.�g��d'?1�{,�w#k���c��������U1�U�O��;�jb����O�	�_0*��j�@]��mw!���g�l^�y����A;�ƁV�t� *�U�	���nܠ�#vŔ�̿d�X���{��D�]�mq�T�D�����]��,9_f|�4�+̒VW�#eA�U �P��/l����7Y#��_�p`���(U0ȯ7�R��tkg��#e�����!6�.�$�i�`킮Q5Cb�絺SJ�-�.��!8v6R��k��T� �j��1_F��8��1/��x�7){V�� ����*�`T� ��(�UJ��nN~����� �ݽ{��ם�h�6�����A�0j�D�wO��{F��A�$�y()-��$9�?j�@����K������էC�e�s��v+H�3����s*����.�����k���:n���8$,���wU��]���e�h��q!��M�A�)<��\p7���euuva^&����.C�;K��
�{��z�����l�2�ܲV��9T$$#���[ҫ�=�]Y�%�>�:��U]��45k�R���Xۭ�����(Wcs5Im�K^^��ip��xkq�K�܇\����;�K�j�MUz���PϠ����w�]���
։)�yM,V��B��wt\9v�r����$�\�c.��S绛c�lJM��ըU�T��Q�I�3�J\����</4��wۼ��J�֚�a�����)�[���:�@�����ٌ��O+��:u�����;���μ�Z��n`(v�o0��۝W����������;Dd�c�2f푕��z�oos�d�Q�7NqK�{��{���[\MݝҁvT�q�Q�G*O�6�K�8�)�1�8��M�X�=�+���6����̾*ګ�U\h����մx�=�r���y��ƥtm���ҋN�'W*��^��g��n�㼣Ӝ�f�Tѽ�t�z���޽V3a6�+���8Z����˕��WO�������[�g����K�ە+m���PyYr�[� ����M1^��(����9C0��O)�T�jmt<����}f��l<��kP>5ڷ0i���;�88�׮�R�S�+{�:��s�CA�_+Qs<W~XI����j����޺��]O+:�ɯ����˳r�\&�K���S�D��;e�������ya��$Q�4i_���џ�TԐ;�N��OC�����a>�&�T4��q�J� u��#˚jn#F�Kn��-x渜>��i���eXU��Ȥ&iA3��V����:�a	Rթ[j��sI�>rM>������М!0�7C�.�4�E�W\_�X�B�ٓ��|KrN�+�N,�N*��O��á�;��	4��Y>o������CB��Y�R�VI���i��R�|<<>�\S���j�0��d9��f�n4b!3�g�<� �Msq�Z��=8xzw��r�`g��t���ei�h4Z�!	�Xf��Gmm�R��*�,4�������Qz�n:���n����d&�0np�r��G�s���Qa�PWr�ba�͘M��䯐�\($�*7S�k2swG>�Jy嚸4^\wؚP���[N��m�MYQ��ZÀ�`���0����9yy�fg���bM���R��MwX&�s��?"B(� �B($ �B �  B�~w̜��Oy�=&���I��l&r�&�f[ne7��+P:W�R�^��u�����j��p�����q�8b\AF�B�Վw��~��R�P��"-���f ����C�*�ޗ4@;�'���:��}�������m}�ҾwO�ʩ0A5H�7T�ǳ��m84j�\Jh�nж46tY��GB�����0�c��A��@�]��Z��Hd�qK=fw��A���H�2���d��3,���_:��5I���#Fp�����`N� �oS��ٿrw�q�8b\AF�+l3T�G��.�"��2"ز���40��g��[l�-�N��Ox���=|'�8[��k��Ҿ`]?�@Wk�܏G�j�>��|��ֶ]-R����q�;���a��>�}�� ��ǐdz�~��u��mџw�,=�o/��)�s��/��ճ�4���y����e��/O4�朳���RGg���+u͂ė1RU9�S�T�Z'u�2��}"�B*� �B
$ ��( �B
���}s˶s�ϥ�V�B�.���?�R�L#f�TH��֬ f��u��4�n�8���w�0P7k�'�*��=��@լ�%'��7�2QP���镻T�X�،����j���t-Q+�v���X�~�|������4��v�������8�nxg_%����Z��9���4F����_G��{R�5{�w��4Fc�{�Q�a��>�}��b�$�P�?Z�$?m��۫����U A�}^�%�T���5�Ĝ�p�n�5Hsw�q�hĀ�C��@?�,���!U1C�/�h�;=����� ��"�|��D1ݶ�}�'�8+���@A|jW���p|���d��#A�O� 5 �?YdO��E�3F�	�)ޘ��`l@��z��^�=�$p����d���L?��Zjwt��ʇ�ʸ��8����j����*�����i�غ�s:����GW+���Ѱ;"��E��/�j��Ȃ�/������D�]^e�D%�z�4k�
}"(�
 ��  �"���)N�y�����R��B�c�r䰍3u��=P��d��mdpݶ�FhF׫)�� �.�����l�i�P������t0t1��@�5��XYK�^F\Z�+WF��.�\F�y�2�Cm��������f�Ի�� ���IM�{��Z�#��u�9�#��5Qzٙ.\�Pc��:6�Lm*���5ڦ�rD+��}ߩ\����"�f2�lT�Ņ�a��39Y�h(i��9Y�2u���c� �5a�! �ƚcb�
��;��8a\�q��;2�#P��A�h�`�*�|41���p��Ӛy�fy�ִT'���VFw�����hW:/~6�MJ|���񿼻o���&гܘ#�4;h2SѢ���"�,v9�{��J�CD��9�0L/��ł$��E*IH���^�į?I+	)!����&6/���(s�3�� NyVp�ߎ��V�+��̐r��6�?��L!v��f��{s-v�GH�Y��v��ƅs����	�L�E�!���J���KV���S-)m����}��֠����kMK��.0K�0*X����issaM�G9�2�so�4|ERt֋�}����p�w�1�la�4t��7�p���|��|����{ڲ�{ʯq����CjM���/��n��f��T��*��U}�y��t��9��K�C�L�K�U�u�:��+_}��k�d��y瘞A
�� �kR}O�QHD�UHEP�HE �UaW����$�k�����,�(~w�!�p¹s���ѣ���XC:���<�AZ6t�T��"���d��0���z���|U�ӕ�	9�Y����*�QS��xQ&�J���T�s��� G�?%A��O��������dN��8��jMwU,�ur��ʿ~n��y�x"B��	˲��Ν���wᯆ����G�!s~>���xC��"��R����@7i�a� ݥ�L.�MX8r�]�f�\]�8�Qy?f0��E���c�ۂ�ي:)��5��i�iIv�D�v�c�.��I�ɠcX�� W;o����ł�l2*�J�b��f�{�ϼU��h0H�[1f	ޫ�_q��9���mIl�v�����m�y����A�1s]g��J޳����0L,�T���.�~ʪ� |�~ia�i{�5��J�f�0A5J��,̓���!��=�bc$蘕�u�ŵ�Ь�|h�����J���g.����tw�����]>hּ��>�P!XED!B !B O���]{��}�\g+��~�n�Å�@�P	��;��˩�vH�6�?f[q}F���7�����s�����A b{g�8)���e�"NJdz�Q��5H�a��<��K�;�`�l8��<�V�.���0~0l��a�T���TDP�n+�:]���V�ZEkfbc�5���`]��GB`�1.�Ҽ�Ll�ò{�\�zW�t�|n� �(��38-��]��1��P��ìA�|���� ��}��y�sa~���E�2ٲic0��2R6(�o��`f��ox�����|mq��!v����i�zx�׼]��b��gPc�A�� �0zkFG�7��L\��Ҷ��`���7!�փ ��B퇠�������6ioeNTt�_38��F�����cL{4b\A�K����c�^�]Р��[~�JW��C3����+8>�#�b��ص��*���.�mּr�����W�����YQ>��H�H�B(��, �B
"B
� ��>�����
��y5L2*�L�n�Q��R2s�t�G��g�1��/��|A*S��.���&A5J<F��8�9�2.��V3]ט:�/��n�t�@�l���r��c�g[�A��3T���+�2����\��G�"w�|�
T�~of1}�|�,(�����ed�^r�B3��Hj�ٟ5x���yGQ@�c�=Z�p6P]��[2bs���B���h߼{��5��0O! �[`v/��`UW��f��y7�o6)u=��nc<U���BM򭄙�(��m��9V��h��|�׭�\!� 1�I�ESd�َ������?"�De/B�����(X�RV�z��U�*P�ƥm�y���I=�X4�Ls��o���8eD�}�����a�*���1���?7���"�����2���')�OLXmވ�R�z愣u���؁�T���{6���-�	�;���R3�����[�*�*�]�]\$����"�
�"���� #Ӹ�I�z��$�긵��k��F�D��L��(B0�rM���g7C���6aQ��)�S��iGVX5�i�Ae+�]��31�!�[��h�λk+WQ^�cve��uэ# R1u��%�;m�P(�#X6�s3ŻGh"�VسU��厙$�F6���flł]��Tb��Gl������հ�%]+���Z�]*�MV�}����v72�g%y�25��BW��V�4���E��X�յ`���c��0~"�2/PdU0�&�ݷݽP�7��h�6���:�~Ŋ���փ9��QB�J�!^S���X�N�?up+��bD��1�6gָ{��}q�0@"-|�Uш���>�����90A9�~#��X �d���ݱ�g�����w��hVƌ���p`��Fc�*�AX�!��/X��d����p>��X��� ���}��
c�]��u������<�2���wʂ;�d�H��d�`�%�%T��w�G��{=U|#Dg���{��}q�"�T�"��� �!�5�!��+m:�J��mnm��3^�1�tR�iQM5���+�039lDz�����Rd܃�2	�O�W�_wlpˉ��|�H��񱗶��5�&�W�/Sḍ�BQ�(�;��BJ��K_��&���w"Ѹ�p�̼���r����n30҃r3~��3�]s���}nc���H��|
��l�9v\Ϛ���'�*��"	 B�$")�~���|��>�A�~�����x�����jS �t��Wۥ5x+���aH���|�C�o��f��틊͉�Q�P���Јɝ��3�A���>>,��UC4@��+��R�/����
��. ����U�]���[2���
"�0�^���;C�5��> �������#��".c��W5+�m�9��n�!�]:﷪��]��k�RmQT��Q�R"3��с�0}}��Cb3[�f�9�2c����f[	h�[ �k�7��,!66�?���z��z���=T�5OG�����=���x�9�B�ز2X�%�����a���FS�e�~VŎ�4��J�ї��|��X@��:f] �~��nЀ�%�%yI~ݙ]W�e��K�/>̲�ܘw-K����]ci�&^��d.]�u<�nV�U����r�t/�)ԥ�ŷ�wUvo���^:-]-��G�n?HB"0��� ��B �����k�w��>y���s=�_XBo�d&r��Sd�*�xM+��4"��*ދ�}���=��/�Z�b���T���d��>�;��+����՝q���ta���?�R`��_T�f�+��<`�fłj}����6���pĸ��A��a�U!+�Jc�s2t��.z���i�YB_8�
�ˋ^u��Q�#�jH髥0]F9` �v�'�������0;l2*����WFwW���;�CU�"�¹9�y*~ d�߈5��z�T�v�m�醫�u�؊���G 2��ɪz8Dd����	����wӰq@����{�B�p+��~��pA����~�\#Ô����NzѶ8eǳ�k�6
 � �a�T�T�U0���=^6��u�{�S���R���]�^}S��o����}I��W�$��D����G`P�������	}ݜv�Z�jb吥P��G�>��|'����+�u٦�͒`w���V�/��F�-E�W��=��*}"� �"0��"���"0�!��ќ�\ L���(̪ �Z��5HW�����Ϭ`Лj����Ot����P�c��T�c�X+k�kH��>��%�!������N���R��-��<rVc4�BmJFRiX�ɶp�r�w眴��LE.!�T� T����O���8eǳ��!띙c�5��ʻ;Z���N�A�!5�,+1d�fø֟��P��ϽkHu�Ϸz�����_\��L��*0T�w�]z����Ӱ�� � �� U&?U0�`O\��d���}�삽�ߥ�ʲ����3-�̢�b�w#��V���>1��-� �j��}ޭ�N���8fG������A��Ӟ���R��`9Z�@Mk�͖@?U0�P:�x3{��-A^u=��O�b����uڸC+��s��A&�@���;����U����r
A�e>�Kb�k��"U���œ�w���W9��3��Vj�%���P�]��m��y��̭�G���v�������.�|�uV�\������B����O��R��
�-[�qV�9~���x�y�Y�NۡYm"��6�@��71�Z�����R�r��1�Y�F�pf��Je<+"EQ�0a~�O����%p^��+b��r��M�
�H���C�W{�&Lw�[C��+ͱN�eI�/5�x�Y�f
���Yλ'%89�{�*�;�.����L��I]��5�h�����l���7�;M��M_3��b��wջ]Lj)2��`vpJ\#��L�ʏܯ=A��gxΊ�B�[t�A����/� �u���Ȱ=�R�FV�_���.�y6��R��I:�l��3�:�4b�����[��3����~Ό�&�{Z��4���Q��h���#�NYG�u�J�K�C>�EEP�W�r��<W��),\�r����Z�E�UD-�&]�M� �X�]���.V�:�&�3��S��J�s.�t�*�yi7��P�{�BN�������3)-z�U���ӳK<wi�>�+Σe�cN9�K�_G�J#L&TSQY2f�V��<W�dɖ�f�������f�W|�!�)�|6MW9�yf�D�8.
U�6��\"�z2��:h�*�*�ڧ���º�!���jz\Kr���y�T.���7Qw��!��_DB�;�>O^B`��k6�Ҫ4��<�Ry4�w�<����ЍQ�`���M���0D��z��T6�����؇�����%��2�-�>J�p�[�zJ^����R�:����N ���@��k+�ꨢ�ެ�Hn�i��$	�l���Ӣ⏕1UC�E7wy����w^9`�$}�N>y1ͤ<�	��q��:�([v^@d$�͘a��$&��*�J���.�\\xϮ锨Ĉ��b��T��.
�Օ���xt���Ĕip�u|a�D"L��b�k�?hx�C��ȹ�h�D �����:zp����*���*���+��e1��Gh��̕�����"
4B�*"�2*k(��>1����**�%�����"�)Z�n6�LH��=��_�.��:xwz�Q��#�m��#��D�+S����x:*8��(� Qy�:�*�8xt��qq:ʠ�S��G��hGPpDW=�dJ�s�k�Y�%_��l�QG�����|?:t?!��S8����򚞦�k\pU-ܴ�%�qDDZ�Uu,Tv�E���D���Uq(��"".�+�(��P뫳��-r�%EPF���U�l����4�w�M�U-t��0��u��1e�L�@(�� h\Įu�B�V�+b�,)vr�[@���a�u�������Z�eQ�qi{-(���ef+3�%��a�a�m��#�כ5��1z����\WLj�8�+R�,K.�f	������R�%�2�˶��tZ�1��ZgUkfa+h�v��:�SVir�����\�-t#��U��L�Ѷ�h	����l�#���^���n�v�4�l��Me��&-Z��Q��n+4V�޷A��ͤ]�גWRV�ln5A�d�X[�JR]��[LD�j�/Sl]-�z��h�ū�F�� ��QS[6��k�[6Z�2�1�M�7��O-��<kkH�6f����SLYR�� ��/�]�,�Վ�8����]u�-ÊQ%yb\�5���[T!0!�M���b���+����|���[4��y3�����&.���6\�07]�K�R6��[6!����MC[�f��d�F�R�.YKY��n�0q�v�X@Þ�f�r��X��5��ѶiiֳPM\R�F�j��Z��&q��2\�\K�4��+�Z�JUnu���e����av�ckqqr"\�)x]Vγf�sbc.��,�J\��4��1��fU�X�P�+�1��������y��iM.,Y���̭EH"�P�q���3�[�:уxF��;�G\X�к��tvbGM���pT�:йk(Z]G�f��+�򌬯��i[�<j�K$4��fd�p�"��q��J 7�CF�#,̳�)Lvi�]����MK���QҢ��[���I���,ЖX����8(hˎIXJ
.�v�Xh:�-���H2�e�j��ۚh�+Mf.&�R��V���ea�]�SU�v�uCM2�[�:[X�3��1��ls�K��ËFz��´�����굻�O�!DRD� @�N>�z/#,��]q�KGe�[G�2f�H�#vu%͋A���Y��=E��CKeas�h�V�2���626� G.�ɬ�MHB�SD�uy0���DN0S@EIFf��,[����� f�s3�m˦�ņ�ln��k�
�4֖0�Ԋ�1	H�%6��5j��͌�)0a^L�ve����0:R���(�`�%	�R���H?^����X[�9�l�R=Ys3Wu]�%(]���f2�?�������G�'��Ll����㵨��w��p�}�w���h�`{�ő�`_���B���|(hZ?Q���JY�G����w�i�q���{8a]�C������f�{�ú�:�{	�a����p��2.�)����T�xڰ����c��&���r��Gؘ �VGf/��O���ͻ8S�q���=�~�4|�A纝�G'ӽ	{���g@��e�l�>���r������)�d:%S��dp�d� Ȼn�ܫ�+�I���7�J�U��wLh���F��y��4X�&�Y�fB��G$��L���"(�pTcu����D�a5�Њ�7��c1Y�L����5�!V�,/X`�&�۳��y����^�^�\A����˚7�������� �&�J&�P?]�Ց|�A�1��&���]g�ԝmUn5H�6�v��{&�I*�ق����)*�t�,���դ��x��ͭ4j�\[��p�ur��ٳ�W�'u��Ϫ��A�@!a! aHDX@ �����.��Y�������Ҝ｜����@��b�|F=���g��U?k)���3X��&A�?�R`�(�L)���1�'[�U���j�bwtY	��ܬ�4�A�.Ш�=j��5h2A�b5�� U?�����u޹1����12{�8�e�Vb?�bd�R`4�(��%�J*:�f_g¯
��z���L洧G��g����C������Wb_m3���x[����jPm�[���u2�L��t��n�J���Wjۢ�cAP�M��� ���5I�5I�����xZc�F{8b\ExwYߩ�ڨ��~���
��r�L1Q�T^�,�b���A�F��6���彧��r\_WZ\A1���3T��_�vd6��GnN�;�&|���-���4JLGݐ�vz�t�T��/�fmj[��2�\��Z��]�Q
�9vZ̽=t���ȳ����mT���`°32���/�k0���'e}�DA	��U� !A@ﾫ���=�)������(�A�j�`���R��l��׃Ov�^�"�:v��`^���LA�\����i��щp?����
�|}���v��|n�`�+���U�v�Σ��o�o�9u�x�tܵ��֐�r���� ��t.d�y��%�W�Q&Ȁ�i@a3# �Z�t/�0���;$o:�A�Mv��>���e�A�kX`� ���;�VG+^����w�2��n�����$��_�����5I�~�Lu��TG%}y�=��Ħ
���}�^oYLp�g��%#���`�%�"�cs��ʰ���z����wl0ES��}N����V���d9W�~�:j��[����K����b���|�Rv�p���N�!�OK�hw�X�b>4p���3%VF�^�5�W�y�`�g�]-���������t礤pJz4=\o1�n��C�lז�U��4]#a����&���w2�x�������������!!�P���P�T5vt�G�ݺ�aa9�l�'���՟��/�@3�`��C��~5	���������$�8b3f� �P/��D��(3�e�%�e�T�`���%s�(��l�8��lb��  �s��9Z���a�*�tA*!������uԷ��֗�1)`:u���<��x��~�&�F�H0ExBZ�F�c,F�2Udr7�����G}���c"��Rn�z:W+����k��*!���?�=�i���F��v3���g���
�����Gu�0�~ �b�]�CCYӡ����:l�>H?��o���*!�՝g��uԻ�p�u��\�!�ȭ�nB� ��/���6�P�#������/ǯ��Dh��Ժ����Dy����{�F��>�z��	�e�6���Q� |;u�nځ̾����Ď�qVc�}e{1���{.q�.4�Ȋ�� ���~��Q��//��W�0J}1�����篲j�R��]�^�[�W���YW�E�V}D�A@ED�@��y��e��ġp�T�V�WMb�Ŕ�BB�i�Цm鞱���8c.
�\Л�A6�kn�{%�dp%�[j�k�]��cK�tB	{LG:�a5�[3cp)e5"�T��
E���[��	��Jm�潦��)1��[�Bdn��͂ݎ��_�_.��e�c���mx��̣�j�-M��]i�����hYP����g�?\�l�Ҕ�Rm�cȘ.+��Tm�3�Z��ط0b�j�׿W�<�}�/���L��g1h�bgN�r�-�g��b_1{��T����~���?X��]��h0|	3�ۈ�S�M���{��9ë���=��֔�����_*3T�����^&Fbdk@�a�T�������[2�����?�fs���׮�I|���YSLF���%z������Hlu��X�G�S�w �YO�e�K�Ո���P������ ���=(2/P{�2O�e9(0A�2*�FTyc�E�^нw�?�g�Nhꮩ�'�֗�R~#e%#�(����e|�~��$�jV��h���b��$XX���� H���Ԏ���S��h�\KP`����� ȪA�I���#������'��Do�c�
��6�dn��"����L j��q����}�=��qq��g+�u%�ǣ=Org։ƾ��l��J����c��a���Q��s�v�v��j�ٴ
�湫���&j�>�"�����@��)��""�̷��ZLr`~���p~�Yq��]�ĸ�k�A�Ec�!Ṏ�C��7R3�������a�T�
���z#�=>������oF�mM���WZ_w�)|�K��L��N�j>":�g�TO@�9q�� ��g�`�T�͓w�Gu�>�E�`�b�`��{��o �����2	�Lj�I:��,����֦66���q�c2�b]���d�5H�S���q���.|�hb7�&bM��f�c�=t��]�E�-Av�K2�D,����5�0|
�a��o��;������W�m/�m
�:��V��S����&�C�<�_@5����aQ����|bP)��&�4\z{������ �п�ز$~}��o�����_�~ �Ҭ�%�F d� �䬭/�d�/�%�y�7�ݸ2�FDEUa;�mu�c���{�қ��v�Caf�TIk�F��]��m:�+8���B�7Z'��NūֹU_Q��� B B BB)^y�fzw~��3/�%��|
7�2�|v�"�E���=d���M�B�"�w��g�t������^���r��nn&.+�|�(�z�Ҭ$�_��d�(A�T�����ږ��s����Ou9���}��b�d�:� ��c�DE��^��\	�$�`z��BL&��F�[���`������9rl��]��ׯbD ;ؾ�R�^�.׊v�Ƚ���/���2�b_
�V�VlS��I ��~"KD�`�>xpMr���IX�/0�8�����շsq�+����Bo����x��j|��h�����j��Y�.v��Z'��	�A�~L3F�U!U}����&�{�WOk{��u��Of�e�����̦�W!seS�!�<UFz����_X�D?�W�( �*�;�;�zM�zf^�+�ޠ-Q�.#ٷ�=��)c�J�����o�]xE�I�E��7��OD�"�x��a�MM�!7O���F�-�<�X��}ۄ˛ֲ�ϟ3�?H$"0��� 0�>e��}�ϐ��e�2��,s�M��}^s�85��9�xuu��t��u%���D3T�PF��&���T�t^]�*-������K�{qT�1F2���%��0�����X���1��'�����!�H=��h��_hw7ic��uu.�y����}R�[���p�͂����4��R��T�"pzj��U$x��?M��y�syM�G����w��|A�!�h�!FekñxQ[�b�G,�*�T����<�JzN9��2:��n:ez���A%?��D3T�f�1�7�\����@h�a�l�d�l�w�����?p�MpA����s�~����<�4ѕ�h��V���	�[a�L(��%v�x�Lt�^���7ޏ'���~�A� h����H��Z��{��EĄ�s�<K�}�2�d�Dw�]�6�����j�>�*�M�_ܗ�)�
]չ����,}��c309_@G�Г�ߟϨ�S*�d�u�n�ŪkU���A�G��I<�ׅ��j�ij-��.�fX�{Ymm]\�����l!mZly��"J��X��v���R+�cF٤��75��khK)�)jL��C3p�h����-��H,q�����4�����Ô���ik"2�$�H�SSm3�73sm��tn�*Z�˄�E�&�;ggVl����4i��kJ�9����:fY~~�_?z�6�f�����@Xus�c��f2��!��:ME2@�������|�;� �X�]��P�����[c��u\�t�z���G�HuO���cq��;��4
*�"�T������c�`�2�Qc =H2�a��V��f��T����C�Z�&�dU{M�A�c+s��6��IK�R�����p�ż�'+�Vd�(����8�x^��n�d��$@B���_%�o��ρ�/�����'4v������/WR_� ��!c:m@��*o�1��jȪZ  M�ݰ���x<��ع�Yٚ��u��}���$"�}T���c��������_��=�p�pӁ��P�9�=F`��f����6�1H:Vl�?��z��y9`�x�!��+;�9�ҷ%�Df^�K���ƶ��{�wsB�U$�C�}T�H(R��R��ӎo��y����#xt�Z��rfXÈW*�a4�;��ՇQ�bf��sF��X(����������]����<�<��?>�HAa�F@Aa���;�y���~�g��OT���L/WR\A1/�@(0��N��^\�d�|ޑ�џ���7�A �� ͱ&��L9�s��R�7���vn�_�����shX =�$� $��Ʃ0D[�%�ED<��ً� զ
4��{�7zy�������B>0nnOt��:8X� ��<����ݠ�h0ESQ!�!-Oƥ���ô�N�����m%���0A����AU(�5J�ǉz��R��r�R`A 7\%eESnu��`�F��M^Q�b�5���,�/���?������*��⚩�w�+�YW;���[�C~#܄�-y�BL
��A3K��;}_`;I���/�n�OFJ>q�|1."4� �V�7hSR���=|� ��� ���,YL�`����x {|�?�`q�̿�A�wQG��7~~ϦPH��?\r���f�Gw�9v;��}N͉���a[���I5�"�=ҹ�fGeL8L�H�:��{�����y�I3j�4e���=9uO2@�0�b��
\�$�U�Uđ�]�u���ڼ��`�:�j.ebܾKwgUv��+�w2�F�{oD��R�P!l���U8V���pVMTy�L�u1��y���cA�D�Ģ�7o#&�STtk4�I�n�}o7�ͻo�Mi��=F�eCVk{���o.�˭����96��\�R�K&��>���F�*�]�(v��GB٫��4�f��"v��vD�b�"v�t�$���ȺM�����7�R��:��ٽ���z�#��e��h����9�Z���j-��r���뾧U4�ηȝ�Nb�d�uC!.k��^R̰EvU��v�Q��m�f�n���N��3��D�/������]c����z[w-!{`�r�6Nmn��`�԰۽Jzi�#��Ҁ��k��(�a�4�Fȫ-FD�p���rep5S��K$�d��L&d\yn�:���׀�*�9�غj�&�T�Olڪ��ާ�3d�#V(5����}-��i���jV�IpE��o�6FK�ջ�̳�U�����^ga�ʭs���F�ڵvP�d�|֍�]/�ct�}�Պfl8k�6���7��-u�n^ȇt�N��ev^RYG�t�A;��/(K�T�/g��R�u����D�A*� j� ���0���̃K�Bd	r��)9,7*+�?3������Tw!��b���|O�*T��3�*��	9����"�(���L9+2�+1_�鬊���Æ���#�"*�lI�B1(�`Dq�dAr��wM�QgpS�)^�:zxtQ^!v�l�K�0Q�,��9�I���[��u$�j�����Q�9�Ç��çc)�C��VZqƬ�2ݒgH�QQ��E��)����K�V��������E�*�\�W��\D�q�W2�6�bUg/,��<sOT�\SRaMKM=:zt�(� A&0E��{�:8��+E�����n���H��sQu�q��hN���:/i:�TO�n�5U���O��#��8��
*�Q���ʗXgv�M4�x|:tE�븊I�h��##S�8k8�k�� ફl
k�D�����}��e��:i���ӧXW	'��C�.�Ĵ۶L��kR�d��*(S,�&*���,x��\��9ʳ��۸j��+V��9%2��Q��ء��n���a�DdB��z�w��]��^���~@�R`����3�Rl!_R��sz�����H2R�|
����ҭ��)���~�}�b���-���\��V�cI�R��U&�A��LU_M��J��qhy9C�zz�A���}����A�An��R^Bb�sݯ-��;r8`�~��jvc��,�W��*Ȏ�r��E���]�qQ�p�ab"p��V�L�����M�ך;OW��o�ǫ�."4��na�n�aj�9i�MRb(�`�R��*�nz��g�̐�����u�y��k��*������0l� a&�Y��}3�x�E�}�O��_iQ��x�
�xt���n#U�^e�d�>q�z0��j�V��Ѣ���ESv�	F]������PjO�'XdM���GLd�v���Z������1��!Ο����b}w��M�B<��tl����:�k߁��o��k�Ok:�_{��7��u�z���GĞ�'nqTt�D�A!a!�[�G<��!>�\99tBs�XC���%ݙ����6�~�.}�6�f�Ү|��z�Bt�vh�;E�2휮l�L9���]}�ߠ���Ț=�B0�"	Ҷ��0؛n�̆,�p*2��3s���=�}�b`�����������Ob�����T�����+���T*gP�A����5LB� `�T�e�oo&3/__	��y|���w:;;�Gx�����K�5PGe���������+�����,�	"�}T���n�KO��~^Ųߊ��SY7ޕs=��b�D��}��&w����Υ��>�@U.u�V�grhq�z1.��5�Y�&���.���5lP�7�*��"�T'�ֽ�)(��}�n��gm���Q�7}%z�R�~�&A�0j��k�P�c�쥘A�X�ǝu�������7pO�X#(O4�g96i����L\<>B��ȸ0Kv�jlG�d!Y1IL�B7�Ȣ F-%�+EO�HD�F$�!�稓�YȻ\�^�D�t˔4Ɔ!0���M�,�Kb:h\����
�]`ee��-ũ�T��6�]��,��2X5�Ü�V �ֶ��]���GL�Mk#���j�)��B�&tFۘ�:�t8I�FGJ��#�ks�`E��뛄,�f�����	�.��N�K���\�\;�i�1��c<������`���Ϛ^��ڏh6Τh�È�YoR]X$\���� ���ԙK�_w�����5H?�5M�7����[��K���� ����IH���! ���3��6s�zL�ఌ�U�ڽ�~鿝��7�h9+�r��ݼ]ӹ4��^�J5��~7� �C:LY��J��L?�A��5!���A����Ʃ���nLy���b�n=��=���+�ԗ	��ne�9ʲ$�Y�����������!��A�wV�v��Ǚ��[��K���a|�!F��=���Wգ�#>�~r�b�IX}%|�n��0����Õ��5�;]��{4��f�H	�8�6�%��	,n}���1R��f
�����!�n��a(@P%*���%(��jIt�4ל� 	$��A.s�	�A�Ek���T�w�j�R�Z��}I}��a��j��R�A�u���dj���$� � �!��~ޟ���§��*'����bɵg�Dfm�t�gE�ϻ�f𝗏������|���s���$ܺԚ;�C|���>�!�D�HAy�O~�h`�c��;�����}s��c�@��}4�MZ<��dL|���_µ�8��|z���B[`����c^<*�Q����^euǯ}A��fpľ�j�AݿIA}%�!b�`�'d;��tg����I�.�l�HMA�`W~RW־��[���֯��_R_p1�Țy�vo	s�������ʸfU� Nr��T��� b���c�(	���u�����vu���A�
V�sLЪlH+�om-�0���)��-�Q	�\�٠q(���uѲ�h4��Rb:R9�6}|���?Z��}�6��jԃ�Zdnf��z����g���'n�ܞ�^C@ ��?��)��p0.А�	7r*�գJ(3bA�na�j��`
�W�|+]ˮ����>c���[���s]}�?8wpb�<�Qn�	&r�Q��&eB�{g�ĸ��]��^X����3ؑJ��K|X��SO��ٗ��������"˲Av���VŬ{e�6nrL�������y���wP�j���E�!!0#E=�=���}>���f���r��~A��c�L?��0$*I�i�#��wm�z6_8 �y|��L�j��댽��_D�/=����h@a^�����gY��
*�����pny�*�`���Nj��	$��}8��V������̨���H�&dկ���~9��"q�B�tn��y6;-�e��9���
],�2�!�fx�!���k�0&���?\�"��A���v��8�t����a��w��m�^�׽Ɩ����E7�����R�x���r߄���A�O덼�=��s�=��� �$>��bn��DKވ�a��¾f��5�.����]��r�Κ�)ف�q�_M
�\�ܧ}I}��n����?U&ER`���c���?w0�5�3`��;��fY�1u���|��A�#�ʼ��ΟDy�Ɯϙ�ؠX�W���1��].)��r���e"�N(�.�T$��}�Yk�eX<n�ۺ{�|��#�jy����|�͟@�FD�X@�$cC�,�C~[o2���Y�/�uQ���&��W}����������]��s�=���8�'����Z�Ey���E{���Ę��J(�٣fЋm��"J�B�n\�#b�ƺ֮���[��hi�A�́T��<�7{�u�9���.!��Y9���7������LhPb� n�dv��Y�
�fߧ�I�A� ����0p�؞}$/sŠ��M *�|���Brf��-�|�B�U���!l䩲T�#��)Џ(])��k~�y����2�!�,��6J�,�
�Ae����'�X��B� �z�}%���/w�����Jwԗ�ɑ~�'جq�R2t	����R��A�T� �-����'�b�<a�����wb�dz�H^C�QhAH0D��*�ګ������l�dfe�y��K��Q��#�,�77�k�l?�0����M&��96�·r��;W�-��1/�EJޡF�F�u{!q��5�>�HE�X8��� �y����w�;�dqo0�4�psb�6�lѰn��ɪ@f�
Cmn�W%��Y��:�K
��0��
EKĪٚ:�#[���se�"ٵ[����s����!��a	+��#e��m�V6h�������V[��эt������2��o��%�]�2S~��<�l�x.�.ͺ����^�f&q�2��ng��w���|���:���G 5��A��1��Y�Ś.l�\�c���P���|������j� ��LtWv��s~����K���ӆ���@ͪ��4��yE����,��(�q�|s��H��|�=��80�[��×��6�.&�)��]�})�s��v�ч:�b���ip �� ���U15>Zd^-�����Y��>�Ay|� ��L?�S�Ļ��`�{�f���V#���$Z� �j�j�ѹ��{�#ל1. f�dy�""��Wp�[	�Yg��9zl���	g-�w}%��i�߷�ǎ����踫��}I �}�]�@7v�
���:��+.=�e��.���%�(�a�HPM6��jєS  Lʋ��t%	u�tX����?��� S�T�"��q���;��Cܴ���v�5Eh��$gdf���3T��&G:���:4�����||��*�r�~ꜳn��L�.PŲl5%=9��K(^�wo��A��䭢d��-7:��wꘆ��O�|��%U��H��!�BB |M����ƿ&A ���E~�77��(������g�E��e�%r�*��,�6L��=p�- ��dU/�S�geo/�"��}�2�메�.�y?�"����� ��|�������;����3���C�f 禲#}�k��8�2�^����,��=~F
��so�d� �J����� �_���L�r������xdz�F%�6�4ߤ��A�Ŧ�G����}������YfBX\B�[4E��#�Y������\�K-��R���W["G�Y�C����_݇/3��eǮ�S�B�n�y�y{�N��]�O=�p��WHfW�#3(�#�4���'�Fb����d��g��?wNtF\�`���R�t�bA�x��O����E�T�?e/��O�R����]V�y=x�(�P8����,؃�ѧ[��������r՜5�Gs�^oV�d0���֏r���\�r���gy�9���o��V��?H�� B$b��~|�ɝ���uZ���;�گ�w�\�S�VI�Ql��9A73���[�<����O�+3;8nTz�e;�k�&<��̥��W�{ڲ��n��U�3����,���(�T�T��u����c}��N7�:#2��~Ρ~ �9`I^�������ߒ�5�������e�֌i`�q��in��,��s/3A#��3*�pڈ{�\~��"�|��L�V�@��[���8��E�K����LL)��|�A~e�<�.�I9�l��(�Q�����)�DlΊL�n/��y��:r=u>N����c���[�v}�b����#B�!H���$��r�1�"�yA���va�L(ڈ�t�7���d=�� �>��")��?U?�R�7;rng�罉��J�I�&:2�^�[<��"/8b_@��|X�C�w��2�'"|�&��Rr��y�'�ײ�'�wmJ��6k�\��o~�7HU-Gs�F6����Bt�Q��~|�����0�0!���w�\n�ȪlT� �T�"�:㽁/H{o�"E����3�븤�. ��`�S���� �%���9ЭQײݸRC4Ǟ������5�Z��+���RX�
T����R]PJ������}�>��{��S��q���rU\f�K��wrY����%2l�_U��X�T��<`T��Ss]��:�߼0#ɐOj痪���[G"�F%��L�I5o�=��36�B� ���`�g�J$�~����;���RI�d{��oL�z�);�J-0�Ń���_H3I�*�#��@������(PK���ERd��%]�t��8��K.���b�x�K���t�Z�����/�	�u�+�V}��H��w�n��`�SLtz�_w[+��g};U� M�E�Hs,�s�Yr���=���`���my���]��\���|���'gL,Eg��]5R�#7�7�$aY�WY����%�b�(�I�VJq �S82�ˡJ�&���yB�̮���])�措�n:G�vdn�9��w��:�{;MՌ}�;�������N⭆��+#Z���j�R������	��geI���bѧk�v��wZ��5�䁩�%�37R�Pg��mn��Ws��w#06TZf��W6����k��TEf�����j���|6�BV�d��&�7Su��sj���o����an�Q�K5�μ�נ���*�H��%j
�g^�̜��}u�
�XWC�U�YUӴ���ܣ�f�2�q��uɎ�j��H�͋T��tSn�T0�T�:Fz9���[n�Tĭ�Q�DP�&�� ��������X��_���(2nڭ�Vc�7{�Mp���'��T8�Du�Y�,��&HZ�P��s]�-W�Z��a�}�t2Ρ9w"͕u�zwNau[�j�9�\�	,X�"���0m�yR�s��(�ɘ:e��Wv�1���כ����H��e]#;�0�ܤ͔���[��V$f7���^p{ک����]7���0�C���Ԭᇴ�����H�M]����6�e�}���X�^��ՑÓ.�;kt�Vw.����R�NF\�9�]�f�;��,�V�n��)�M {qm��0��X���unT�)�7�ƦN��q|��� W�]��Y�+0�H]=���^x�8�hs|_�jO��7�R�v}V�-GC+.ɫ�%�ty���}z[C�fV5�-����JZMa�.���_��=���%6%�G1j�kγ=�	�\fo����>���o,gS����Du�&�$�Xr��@�py��
䒸��$i��}:w�Y��MgREY�� ��(�T��	�[�tMIA���96)͛_k�KQ>�>��:ʸ��Y��L�skl�qAU�]6J�sHO��[�U][i$�TYӧM�{�4�����9Rq7eVdWwuE��dv���q�6�4�DE5�q�Ӈ���pW��������8�S�uݗ&Eh�FIZ k]�l��2G�1	ÇN�:(��k���U�Ը?0�Ty1d,Ң3�r�X��UgwvcOOON���WSa���J���*"��Y5�ܯ�q��	D����.��:Ʃ	������=e�l|���w8�(�)�HW�m_�=I<�DQ K�$���#4a��g��<�\�!Z����[iY ��2�I"���.Ў@��%�s����gmu̙\>���4aq�S�(�Ck{���j�q�4�֕��l�n�\6&�]2�!�R.c�!�L#�
G4�$4Cb:�ڷ��͸�R�V��B�^��f�B����M�[��s4�X�
җkf��ض���6-[�	M�lN�˵ҍ��J(aD�˨ bg4f@��[���%�n��5ai����!��m(՘6J�K��Щ�����)Y1�H�:�y�ݳ�\Q!�%���Ym�!�ص��DutZ�h;	LB��%15.�T��j�J�-��A�u�`�X�X�0���j��\�Z貮 h2�m�ݑVJ��L�i�YT�0�S$K!)�j����-�V�mm�`&\[,��ˌ�E� ��f0vц�����t]�@�i�<�1�I��j`�!3������,
m�Y�5qT��:в�F�5�\L��,��5�԰v��9f���сrSJ��kq�a�
M��kJ�qp�6�5��ƥBT���[�� kr��4m�4w���5�t�X̐l�!4u�`��m�ڍk6H �ƚ+�v�oh��f�m-,���] �Ż�K��je��i��ea�mM-Q2¶`�`s&�	�� Q��ki��1�����o/2��pM�Ё55�)��m��0K� ��q�y26���ele]|�ĸ��E�^`�q4�ie���kS:�%pa�]��1Lnet�0 ِ�݀�����3�q7T��^�aK����3��fUc�19��\KtZ"K£��F�mCq���H�ݗ\�M��h�¢Y���iH���i�W\:�j��50��a�k�kK�]�B��F#)�P:���5f���l.в�m���Q�(7eMl.�;�K�e�2���iM�����b�lі��*kvo-mQ҆v�c��c���J/f��
en��r30����ː�Ĭef��e�B,\������T�*��)5�c���.0ɳ?����!@���'�o@�1�]�1�Z�̒f�f�3i���X����Bڴp\�.1�c�y��U�t��dGX�f��r�����؎xͼjˁ#��,�n�]x�G��%�R�#he�lM�WƵ%�J���ʳp��lZG\�F�������%�љ���3]s�X),�؎4�a��,�f�L2ñ�ŕ4��^k6��u�� ?_�����Em͚%4ͅ��Z�iZ-, �QR&�����t"�V��{�K4F���c�&�̑T�tV^n����Rw��?��wzw�l޹�y�QzX�$��W����d�=��]�m�~2�d���w��0�{�,�8>{�A�a�.��_�B�҂�})� �;��~�O��L�-�A��/e���Ԭ��H�o+��elyb�gK�"%3H�`�B�2X��J�;�+�R�_E���n�T���ۜ6r&�%��)p �L#CzgQ�9ٞߐ3k�'*~��	ݡd�vD�����7�:��F�K���k&�E�#�0hL�~#%��}%���*��}��X3�?~�J���'��e����Wr��l��0�A�.ډe\ٍ�ɢ��l߇������ �Ӂ����l���7��q�6�p�����q}b�/i��})����od��'5'�1w�T<4�~8^NV�����Cu�Bw�*�R�WN˚m]��2���k4���]�S�Z6E��O���b� �H���>�̦��oϓ��3鿝���7{iq��/��0j�Aoɭd�^J���[�B<��r�����]0���G�����s{7�01��- � �0Ȫo��i{懲xrv�z��_e1�` }�A�N�n���e�a�gK�%��X��|�O^��Ƣ���{�9��7�}����������ןh^8���|/�j/�_b_p>�`���5I�ƩO��p\R������]����5T���5j�n�(J0E0�̰�4	nHAn��a�;�x���� �5L1�2�;c���M�FL|�=WQ��#'{:j:� �03��O�a]� ��Y���j~�kO��D��� ����޶[�����pc����fJ������h>�b���)�`���"�T��_�z�v=ڋ��q�ծqwj��"m��f�<j��u�<�d�!&��h��w2�ړY�~��3�5D��rN?KV/-%�~ GƤ�m�.�5毱/���>�A�O� ݩ��`C1@2-�ꉊ䇈�A��"��.�;c�"{��#&���Z��FrI�Ǯ����u��Hwk���|A����U9�Lu���z�I=��WR��[�s����"m�MS��v�}�����]��߿��֌���g#[n�i�[Cg�K�\�lL��"9q$
p\G��<����] �-1}����5W����ME���K��L������ w��2��'9F�9^!5H>xMp��\��ѫ���P�?���l{�Ot�Dd�,��C�� E��:7�;����?��b��|����~J�.�{z��i���V�3����	� �3^ T����a�@�LN�̾o}^�ʄ#�kd��.�0�v�{�ﻵp����5}�p ��kj��nx�T�B�B���~�y�A���lZ�W����X��n���:Tm��g5-f'sl��� �M����E��{���9S˄'ϿF@�����xL��H
�RRT'o��&g�:�u�ݏp�����W��8���TŀD�/�W����k�߁�*�g�D��+u�m���Nͳl��Tv!��:�S1��]��񕀃�_1Z�`@UJ� �n��ϴ����Y�>��g��˱�uO��)��Vɤ����C\��(�9�-�Vs~&�:X3�2���5׺w��y��H����5K�}�#bE�8��/|A���c�v���(+�![���삸Ⱦqw��^�c��h��- ��b�1p�]����B線oj�hbjH�_0jf�ERv�M�o}fp��b]��.y	������d�#9�M��A��U0Ȫ�1���m��K��r�8��W~�w���+�Щ��	/<A1S��Gג�Z�2����$�*�ݫ+jf'�ئ�9����{�nnA�F�O�.޽�.�W.Ν�{'�qk'�Y>
�p�@�H� APX�n�,���!?��Apc���z,�7q���6�<ݻ!�m���F��t4`:��vG�ɒ1����i�AZ�#aJ�(᱔.[�d�Z��ز�2��\��Sg p�M�Х�Ld�QtI�\he�X��3��������ê�vͰ��Z�Z@����@���P�zc[��e�X�cm,c��ZtH˘nU�ԌmѶj�c�\�~�)%����y�mt&9f�4�r�5n#�YEڭ�b��^,@M��a��߰��	|?�,��JD�� �0���]���=�=�2����e�X�͢̠�#m�L�5O� � *��"�Tl����'i1�x�����K��%���0A�a�T�C����X�j`��~tP&-��"���O�
D=��;]v]wY]�3u+����v|����E���O��P3Z�}`U�(~�a�wPU0�p���=����/�4b�Ք��w�3=r�������_ɀA�`U,�ϧ/}��=��;)�{ܷ���}t�z����A҃�n�`� �?P�"kVOH�3��=��z�����dUvIy6�	A��q�m]h!F��l�tշ�Yn�U�ߝ/y�g��{�O��9�T��;w�s���ߔ;�K���҃+����b��R��^?Ux8����� �$碒K�7�n������%
9 ��;���gn��J۵���L�x=���h5g\��q(���Bu�\�{YY����! �9�O������߰�ԧ����~����A�U0�E��u��ؾ �* �x�!T�f�|�?M%|5����T<��1Q����K��%�@?�S��S �T=B��<�[QĜ�C@ ��� 0.^T�v������:�ɻ�HH<J`��3�W�>�rSA�L�����B��Bf���C�
��ש�r]'o���2>�Z�S0�S�S�� ξ���Ub���s�=���Ar�e,K���h��e�e��4�,*�ra�`����?���$%��e��י�L!*i���{��S륋����v�f�{+we d2�q�
i�ES��|I{ܒӍ���F��5��=���=w����yWx��K� �^O��3T�'ձ��D�mG�}����qFcא *� |��i^�O�)�֥e}�(v>���4	��,����6�5��Ι�Xz�\j1�ɖ2�؋����eq�f��Găޜo��I��g/f@��0LZ�ST�`��S��a+��}����n���x{��H��� �T�u��\�mV5�щq�@dM����Ԇ�X>� � � �1���$ݠ @���&�;���}p��E�����^��}�q�`�t�`�&D���}ܡ0�}���ҏ�����u��.Й{J@�*(��зl���6e����~�%A�t��C��7�[�;�r/sW� c����x��=�;Ԇ~�0� �/��K��O� �M;xX��vv��ߑ�L~>�����镓6׫?ip�����Ie��'!��5�z9���)l�}FUh`"��4fе���I����S%��!~� O�oS���&�4���a�R_�٩B�tYc�_���l�Fj�8^�%�5�b>@�O�MSdpE]�4!��"O��x�=���L0oP`~�a����N����r�dq�a��#6���CԷ�߸�=y�q�p��G �6�r�l:B��0�4�9sU��t擣����;��v�.�)ٿl��E�YU
�BI7��C^R5�Xz}��!"H���='q9�|��_3Tނ��7'��p���6�����K��Xׯ�%�B�9aa9�.+�ѿu�ʓ=�[�>*2z����4ɫ7dYt(^n��ی�X6�-��k+�3Q)�\�׿0~% �`�������w���Uu3"���E�糈�_�V�@r�~?J��+�W���,�V�<7o,xy�wv���{�E���d|�1�1�S���W����;��3�m'�i�(�m'��a���:�������u��뮖*[U�z��q��4��"�� ��`p~"���[;�x[�'XU(Fo����Et�Z�~�L�{�S��/���O�*�W�zUh�����d#���\
���ϯ�Z]��k���3�{����l��h�Ù�D3.�2�}��N{�����N�=T�LEWwRK���^�Xt���syg��L����zkz�nٽ�u�ߺ�7}n�]�y���ކh<��h��gb��?�����+�M����9��WK(kb۔�p��#
i\˛�a
۳
��)��i.���8F�Δu%J��
52�,��HVWGKD���ZY�Q�;���R��]m9"�i-ѡtԉqڸ�@�h�
:(&�ҠQ�aj�@��	,��
�(��[��2e�9L�3
LA�fins����x����,݌�,�FciWT!ai/������hKT&f%6�5`�2��Gh��5f�X�`�J�4v�o�����t!�^�h}Rc�	��;|'ot�J]U�M�ľ��"MƮ��(2S8� ��0&���Sv[���$I
�����|�x]�=�]LWA�8��`|���T���į�AM1�� �kPd]��5K�*����)sY����~��4M��́����[A�M�MS��X.�{�2�\��og���@�H�z��b�,ךk�-����b\tjP׼��{�7�W���A�]��]�˲SV�"��7Ǘ����~x��=�_W��)�8�O_e���� �����{�F��u,�d)����f!��@0�f�e�!m��d(��C	�{��/���d����v�f᧘5G	���1�O�c_
x=]�|�jXdw7�1"T��j��WOþV��~yKgm�O2
�C{[�]�L`i�ͧ!�����^eI):��{��������)ԉ���!D��$!��m9�]������_�v��k�����8�A� � �0�R\d����q#A�[��`����nП��`<,b��B�1f��n�����<��~3+�t�f�R�Z_P���)����#�(0>m@5NA��:�E��;7�c2>`��C���Jy��΋G�xC-�����wj�"K��%.��b��%��ޅ�'τ����X��K�İ�"i�j�`�T�ͭ.�4p`!$I!*�ϸ{%j5�f&ٚ�8ȷ3MV��U���8s��������	�A�N����|��<v�����]LS�]�|j���r��[^�fׯ�J�D�~�P~ǽ�>�L�,{������`�'g��f@���b�d��dU![�[� 3E�V����, �S]�.Аd�] }���njh���أ�ꗑ�$Ѫ�q=�I��`��������݂U�ٗ�U�`��o4[�Q���^��jn��7�/�lV^��1�3*ލ˷��0*��u��ӮƇ
��v�\�[I�8k2�f��T1>�f�֊�yh��ɇ)��[�{��5:�ˬ�^�AM���f�x�7X�(GΝ�����#8摣G{�������F��.��UM�-���SU4M�%�F���Eg_m
]Uϐ�4{�hg1���n��J�N}H�������hu���oI��m��;5VnŜ�\Y�^�q�Εݻ2�Eb���D,�Av_UV��g^-��w�nR��);�4�,�le�U�Z�t���W;5uy���!A��Ӟ�Q�o1�v�G{g���ks8a9;��b�b�f���u�YU�6�Ʈ�vfwx�X#�ິvdU�58�M��}AM�9]MP�������Q��݂�٬���wAq�����r����W�\�c}��n\ׄۢ�����S4ɰe`Y�t����\�Mm�]h�]y�oK���m����Y1��ƖuV�]u}ҳi��Օe�kz�sN:�Q��*el������C*.�c~~���PJ���f��'{qogey\L�ҝ^��*�:4K�.V��v�bnwXG���r@�u՗UyF���k��W7�TUz+�c^�f'���cO8�֗,�ATC���x��z�
'�SY
�x�ޭ"�4E���7��<�SQ�T��l���u��ӨD����@,����~Xy��=r�^D|BN��H{���S��%8���Ȃ��@�ȍ�g_Y�N6mj~3|M�i;�jJ���'5�(��������		��P"r�}�5��i��U�
r��gw���q������Ӣ�bq¬���E\���%�\ER��j�El
o�Zxp���訂yu�WP��W%,%QJ�DO�i��Mѡ�����������^Ђ4�\���K��D��!SYV���%�N:t�uj�SY��۶��e�	LŻ���j�� NInY����p��ç�vp=�rMe�UŜ��k~��ZR�o�f;hB蔉*HSR�r]H�!.�Y�6xBr���.8����k��n�͊�-����B����0�X��Y��t�ӧDz�tgf\�p��,QTGW
�t�Gi��cMu3f\�_<�Լ�\]�p�qpG�DT\Q&5�GbQ[m\LQDE�5!ww.T��ܟC�#	#!	 B!Ξ|�������;N��%��/R��� �U �OŊܱ5��2�巔�>�b��2����=���75�p�ĸ5+���ɵ�]�Z���|fn��g{O9[I�Qk�(U0��p��_Di����g�B��9;���;���HU&*�8_���2k�|=i�?&�{28�lص���U�������ؘ`ࠚ*!�l�����{�
��T!�D�V��z6rӪ����TdLy������R��|�����b�x�:ͨ��z��m��}~����U���L<�U�Dq�g*��ߓ<	���_M*�c�le޿oD��(O�3����t�UT
�W�4�?o����w@���gEt^�.���N��w�%	�Wٸ%R���~P��q�-��ţiLKV0��yt�V&��L�w�{���=����KVݼ��syn����壍����H��]DL������Wk*HUO4}�H�	;����ӝ�b������}Uܦ~=���ܞW��/�o���V��O�]��O�)�ޭ�n+��
��KB0W��J
��,H�]�%-��.R�`҂0&q(j����1��Y|�}U�f�x�+��ƅ��}����)��8��9�Z�_}wo�w~�GL�S�ٓ��cq��f)o糖�͞���߃O���*+���`ls�U!T�U ��Y�b�]�N��tk�������@����U *�	�\Gw��N��>���*������n�'Y���~� �^�@�R���8]�v���T�W酨_���ꃹ�63�i��.b|�h����<=;�0��·��g��n �'ZV-�sxh$Ed�V۳���CaM��+'z�����{%�[Pt̠�fbss}�zp®�S�.���S�1�8�5�P�$�Y���HI�*=mu�u�R��2�5B�U!��T!����-�$F��X:X��SJm�gA�ە��tsP0�GaD��rP�CM�C:�3��ˉ�]v�ȴwF�U��d��f�e0�F�\v-tz�˗	��\6唵l#1�ٺ8�X]���f�Fg%b6�v��)A�Mp��-K{4s1���PM+Hr��a����W׍ItB���~��b�j�E�JYHכ2ْ���5iiv*L�+�u��v�O��}>ɧ��� }SV;���/>�����o�L�8�s]�D`d��?u{wwW��s���{�4�Wռ�����������pw\"�"��~��[#K�T�D 3�Ȯ��~��T�Xdӟ��ڝ͞�,��Ϊ��U"*�=x{���9�4�����»t�>����5d��>�_P���~R��k������wu��FȰR�q���?w���J6�CY�}���a���C�&��_UW(�*23��QW���A���|k5��N �veQ���E��V4����H�{�����{�
�*�����tnM�sg���8�+�7��Y:��B�US�瘵H�4�u�����a�I6�i�mG�z*q�e܈�F�^�Qם4��=�Ή9c��-`�t4ՙ��cŭR�IdK�~�� Ȇ�P� H�����O�u���t�>����4/�Z����]�-f���Ȣt��"�|�
�`U1�#&l���c�s��q�ng'Xq�t�RT��zejʑ���
����+�����g��#���2:3=e������3(f�ڿ\���j�����*������D�hO7_}�}�3��C����ѡ|�Ttת��o�*_�T�(d�{k*�Dm�	�m*�Gj�hB�5L���g>ϯ��ڪ��K3���y���N��Wi]x,�ݠM/���5P�B*��Ј����mޯ���OC�g:7 [���(%�!UUfA�WwCWs��:��=κ�󺻹Ǉk��!�_&z�RVfg��q������f�>�ԫ=�3C�Ig��s�6��9�EKK(�� u����~� |�3�w0�u��}�j���?�^V�wu|1U�Շ��*�|wa5{�U!}�^b<�Lf�'Xs�wI��>��O<..x�\��.��0]�Ol�T��C�Y��\7}����"�@��������wQ[�*�Aa�&f˭ܗ\EEem3R�C^ҷh�9Lj2�g)���[ܟQ績�Z���o
�թ�[��Q�;�ȏ�<n�P�=�&=>s�Gը�7�#w}�����Y��0�w0;�c{J��y���N����2��}��e�~p�~��,��C� ���� �}~4��V��y��uO�����v.��Ż�)w|=H]*�����*B2���^��}��zr>���٫���٥Z1w��
&�Q+Ѫ%��I�bܫX��YU]{]�v��0�Œ�m�����\�Oj�^�tI�wP�c���ݳ����I�pA@�B0�<@�~�J��݊����k�UG�E��ŅOLQS����y������U�I�hT�m?�MA��>d�F9�
��p�d���C����ah�v�"Ѹ�����D}�̌���\�Z�����-�ȥ�5蕾ϱ�&2s�@�T!UO礭y:s���؎� �?��wa�.�߫��Y߾�@\��E�9͈�sv�vw��\�
��H{�%ϖ��LR���Z~k��9�le�߅ߝS��s U�5����K��1�`�����Z���9�[���:������|�s�eZ�`m��𻀅��>�SW��ٶ�̎�8�v��.��r���#�+Ω|$x�q��|�G�r��㼭Ώ?]��A���b�9���7k+���4��#0�z_eJ�v��]$����@��#�9M'�
p�5B5�*g���>${k��_)>\�CY���ӧ�������֥�K��T��	3�Cm[)�g�����q,a�ycݝ��2k."B	+�iή����[�CWm���F�p��Ԛiol�8�s�E,]��
�K/9������խ\�Z*�`�m����e�A	���4)J�����(#
8з�nu�4�=a���m����8�:ʎ��u�L�MՆOo����-�̮�X\�0�n*X31ڻfX[yL�[n�PRl�	A)An2��#��m]߄}v���5r~kr���K8P�|ϳ�q4��/W������̏�b��b$9Q��=��"+/)��㳸Ż����}��U{&���+������^���]T}UV'ZC�1������W1T/C����%zD.K[�f�}���o�P�������~/v���9�<��^�ލ��|/u�/��ª����}�}����k*"q��X����P$��/$K���?������f0:h� M5fq0,֏F�m.��J̑lQ�	C0�8��8�ZI����ַMs�UsD�7�j���|�bU/�U��'Go���>">)S���r�h���-�w^�g�������k3���n�z�Y9��!2�(�c0�̟+�@��.��Tp�B�9��m�5q\�RG�x���� �W����$����Wv|߽�=9ݫ���M���.�.�,r� ��.�������&Dn�T��EF;�U��wv�W�Z6�_+���{�W�ʳT�T���@������:�U5�tv�y�%�sO�le�5�е�m�.ЪUUY��[��΄������m8�!�J-4�ja�
j��t-�eWm3MR��@A�ǩ��w��e���R�ϟF����~�=�;��������wX���@H�9��#UY��ѥܻy���k������b�^�_s������W{�@ѻ�7ʩUS���n�uyI!���١��o�w�����[���{ܣpU�s�7���;¸ʫ�b�&�s���0�˫ܥ�SI������O���{j|>�iUƸ�l,�֧p銥�W��|*�Ǯ~/����}\��_o�N��^�=�(O��L�����g$��J��������X_~�J��u����zй��__n����Ù��2:3'>VF��B��h��&,G��,Q���k�m�6٢r�%5�L8?����~}�O�%U1@�W�U��oy�Ä����hי�����$�$�#�'�9��d�{��y���Iݼb��G�X���X?xH@'��ܤI1*�N�=/���[�sUQ���Tz3 ����>Õw�2�*��v���T��@USH�]0"�OW�|��6� k�r*���y)Ý��9���P���H(Ȱ�j:*�9��j�KI��kިغy>���Uqm��u-w6+GԦ_�>��������8 .& ^.b���z��U)Q��������$���u��>�T��pU��z�V��2cڥW���T� �D"{8�rJ�΂�J�J��"�Q��f�]�R�[�1~�>����U07vq���2�*�뻫y����{�u��W��Hz�4��:F<����J�=��C��Jp�t����0�l��w��c�� ����*���7ޫ�Q�u���nj_;��7��]����}U�ww�x�R�d}��fm��u}_T
�c;g�;]}*b�^��g��b�{#��P���5^V�C����r���vI��en��a��%8s��Qt�T$�$�<=�{��q��.�����v�[Se=ِ��Dw�]O��ܻA�	^�	y�,!�;��uΕZ��r���Q:�KNVK�?A�{wf�C"��8��X�~�yz$;֎��t*mwn��K�9�R�Y���*ǌ�ܾ�./����׀�Z(>��;k���\*�Џ_�	a��8�.)�p_������i��m�]+w�Zշ�&sW�v�6&��34)7_sJ�]�{	r��⸙��W۾*(�7IW�w$�Q\;��&f��
(h�$es5�W;�����ã٘o	v�uЋ����w�s�A�[��ચ��Wݻ��7�rYw�B�[s��	����W�}�ZU��eF�wr}۷�.���{��0��}!{3֓Py��/<�/
��"%2���;ʀ�͗��:��n�N��R�cGE(�;WRrݩ-�}�gI�uu��ӨUed�{�%乽�l���Wf�ZN�V�N��[9`�x�#���������A��ٱN��cڕ���	N�ѡmTub�9e����8�eM�z�y�g=�:��YMl<���@�t:+k�ꞽ�b�Q�U�ȭv$k7Wa�L���>2��z��m�[�n-u7^�b�Pt��X�e�ihM˴2��e��:�b��ꂋ�󘝏�X�b��Yxdu�ă�)���}۽fb��f��L���'s��aUʪ�3�k�#[�W���)6���lOD���o"��j΄l']���j^��&�z���H��L���18��m��4^=of�>�Ŧ��O<���{�f��w�p�B��f�f.��\�(q�����
ͤ�ӕqX?L���ͱWK��VQ˪_?���׽]|��
��6���l�����<�������|N:�*7��z`L�6���:��0aߎHy|u�|����Ke����P��YN��WU�#����8k�A,���T\�\�*�!$%�h�zl�#�J�!����1�^$!���Cv�Q�	�Vu�_�Z󐤋��K�Ɵ��á���㩯S��ร�8��,\Epa*��bR��DRJ\��*8������Q|s#�
���"�%E�d�l�*�*���e1�xzzt裎9ؔ\QMݶGqPU�*+�PԂ_*����BI2��h�0��{D�&�1X��B��⸹�t�7ESkUW�����ÇN��l��8�q����qp�KP\SQq�}sw*��)6����ˊm㛩*F���:Bu����O��7ı��@�l�	����P1j�qģ=�M<><;�����"�)��U��f�8���O�'HQC��Ђ�)9+��Vab"
/��*����(N��`���	�cz�#e~��+�V� K-�.%WX�i�e,i��Pi��k���B�P4y`8�bFVi�Љ�hh��m2�2R3cF�G��jڌ�Ŕ�]�b\Zv��SUm�.�@Z*uA�ض�kxm�@��7g[��[`R�2]bp�j]
ێ���vFd���3FV\dJ���n���J%��т&QVZ��t�hYZ�����W!fa��?���7��5�M�	�-#���2��y��3�&]!V3K3u�,�U���1q*�Sj،�J����x2�ecs�S:ጭ��Ņ�Ƥ�@t{CBe��a�q1fу���ژ@0䚙�)�zQ% 1[A���Gfe���R�	���Kl6Ptv�u�Օ�����)�FR��qt�`��8��V���q�(>Ʒ��ī9�u�s�l� �c�0���i��ĳ@	@��,.F�L@���Q���Yo`f56ul�$̶��1+�r;�u�Y��^��)M�^vf�[��u�v�v9���\8��(`N�	����q�ބ	�K#�F4Y)mGZE�m[���[3D�(@���P�V�.j�W:1l���3q�pji�t+7b�h���j\�F X���v�E��qay,�j�8�V���kXh�Y�(�5-b��а�k���n	s�\��bBj��`Q
����d���K��%��V��e�(eBQ\�%�4�&�.��Lf�mRT��F��4�񛰧m�R[��J�	cF*Y+�tU⺗7gL2]���Z�㈲̃-p��e@�ȳ3LL���-�%L\%����\��r�x��4#�]BX��SP&�������`��$�h�cJ��C:��Sit�UI�w%���5�*A`]�sz�D���#D	��3a�v�(1)XW*l�9�m�ʓl�Db̰�!j0��g-ͷZ2���\mueVR#�͞�bը:Z�q��+����<�o� B$�f�XU���Hy�w��Y�\�JE�Yqqrh��&�qb��Ѷ�����ݩ	�e-se��X��rm Vk��J��V�u��IF��[�K���ԯ�%[-ih�����뮣^Ǯĵ!�SZ�,���vV�4`㙴-p7X]�SCT�.��J����L��X1�!If�V���CZ���F���&�7V�"y������&ֺ�����?J���Qh��h�9�l`�wV�te����v����h�?'��E�N:�=U�e��ޓz/_��w�6l�'���U.v��I���(f�R�o�퓣8�u����44BW<ĕ*����_D��O��Ҩ+�K�o���	��H���OIq��7��?gy���RpI,	(��\��k�U~0�|�k�U{�S���+8^*�]�V�ᾰ8���|�w?�T�E}UNE�PbFx̛1���+\�ɡ|z��T�U���sΩ}T$�0��zIQ�H-�\FRh�$kn3�fnm�c��3�Xm��P5]=І��U�>�c{��;�F�Vo8s��Os��9}��}��TƋ�� �w�[���j���N|BuaW9����9������\�[bbǚGVM�<��P����v��>x����W}��-�h	�����ON�����G� f���*i��1�a�|��AKc�4o�|�=$���οxp}�����I���z����\�h][e���i�W�qC���jWo%�w�lDVoXo��c�ECӍ�t��gv��\�~]�)����ʗ9�/�sh���_��wª�>���k���y�9A+jlt@bl�q�%6p�g��[C,�`f\m�v���Èy��r�@US�����;]}rb�α:��UEe �Bi�T�i��3����ՠ�6�ο���%w��w�*�7�;�T���=��e������DI�$��.����M_c�Y�q9�R��j-�e�LҪ�l:�����|*���n�v�FK�ɹ��k�7�-^V�M��G�,�1��_��<�ܤ�2�~�;�M,�4]�]��N3��~�B[ ms u����h��v��JɊ�t4h p�b�`��q�r�o�Z�w/���/�UUn��ܟ���(
����";��w��7��t���� ��F;oc~������=Og����[K�&t���9��Ņ;X�4��!e��l�E�Q"���敖�����vu'������"��K]Q��iPݽ敖�v����be��2��m��_{F����VLUY�P?��Һ��,���}4�J���T��2�xs��V'�Y�Oe\Ȯ����������I�	)�*��{#��L�% f��V��ϣ��<̯_��w�H_�ǵ}zw�!�r��MⳢ�5f�B��ɗ�j�Fʐ��$��*�ώ�}V�߲�<��$y�>�HNJL��%G��,�|��_u����17{qB�w�z���/��W�]qҲb�΀�
�uHP&���l��Quy+A&�]�4Q�((Db	o�켎e�=e��P������E���mBf��h�_f�W	k�����7�VoXo��u*m���v�κ��B� j�E܏���ý^~��E��˟K�q�Ɲ�T�]�R)UU\���dU�^=t%������5UU�/�G�Ќ>���Sβ�'�U�r���T������t�C�LdаD�^M��w���x��|�7����+L����c�0U���}=�1\�@�H�T�]<��4�r����}����zN�?�d쎿�3�Ԝ���^s���̹m�+L�ن26��$R��O����[�	+!Յ����W��X��nq�yM�Ɇ,��.�B�]�;o4��|]瞱�',�`� �D�`�P1mH+�Ġbj��s�6Ke(��V�`uL�s*��I-H�Y��2UZ6)-�f�	2m�+6��B������ɃM�<�)�7\���!ݥ�.L��D ��Ԣb�3
�Z��1(�z�3O�ŷcAu4&iC��+&p˩���-�E���X�s�੨�D��n;Wj�m����-��[�\�FĚ�ZVD��kf���9Ղ�hPC�}K���| ߕ�A�n�٣W��?n~}s$���5e�vs��yxr�{��웻��C�G�лz#���޺�=���Js؎�x��z;��`H ]�dۃ��:�g��!����%H~_�W�n�yA�W���^�y�W���R�eUW��B�s��h�
;v�쵛}X"�>@US�����m>��ʈ����&��+Dh�쬠�:�l��ȋ�h:����f�_{%dr[Z�"4�� +�*�_U+��^�PH�����m����`���c���"�Ky^̴�jpԛW:�9�+�J�����5d�UH{/_G`�w{Un�Z��뫾�'p]/���U USov�F�0ؙD�F�-�Ga�(Uޘ�s�*�s��ᶾkz�ƺi�����ז��j���
��P�ZP�}�����>�R�_3����<�ۦ/=�Nv�뎜���;��.����EK�D�ՠ��fuxf7Tꮁ�������q`���o�����v����1���]L�A ֿ�Z������N�+��p�P�b珱����P��s��q+�`UTת�{w����J��Nz��ާ���z���
�b�T/�)8:tb$��Ͼ�&�\P�2���p%쒧ffR,�i���u�*�BJp]���B���L1�y^��w�k��FI����ط��
��Ōc�y$BJ�.����_u�bmm�9o�>�������Q��i��UL�S0���~�@�?�m�T�Sb��Nw$gz����-�w���S���7�����w��}���'��x$�;o��#����Y��[�p�ÛA�*r�ƺ�n-��xx^����O�WϦc� �����U��2j�GŚ��a�8]k��Un�W���k3�����.��\S1�Z�G��Ә�]�<ݻ�#vȍ#a}��|�gN�W�����	�>����LUzݏg�&����\@q�p�Co�#��yD�8�Ҡ�R���l�*A�f8Q�BP�8��Q�����r_��߷5~|����}��|�M����:�*��&����}���Y��
��_փ�F�u�|n����E��	�~ �I��{�w�ԫ_���	�'�)�<���E����B�K��{}�/b�qT�۷T{��J��#�b- sڕi��>��{����݄�w\_�r\M��Wk��y���*(��j����>�����j=��n�d{VmB{s�U�&�)T����m�_^|�鵘��q�%+b�>���߭/����U/�S�����~<��{�����j��Ы0u��#GO�l�3�n��l]�@��R�gI ��?_��ju����+���a��M�h�T����m&�Be����{U�]��U 5d�w�����:�ܾ�]S�Hl}v�G��x�'231؏���vOw�=�M����dˉ�pA�y .9���ܣ��~�*����R���}C�I���Ey�BR�_Si�U�+�YC�z��T��S�ScA�o�AOѻ�r���訍�Uu����������o�
�Y�;*�US�LUw���G�77���`�޷q�2�h^����b�������5�^9�3p�N��Z�Y��x#�����\7Ղ�*��2�U�$mv�ov�yܖ+(N_���5fzw�Y�Z6�ω�[����ŀ����f���A����j��F�B���R4a��♌��.&Z��C��, Ѝ�<[.i�if��c64H8�62���%��ic�llF[�LX�t���\�flk�ZT�.R@�%�SR�Y\��.4ɍ4P��V�fkV���6z��,`I�������R����K�ѕ٨+J���8�+�ۜDM2���=Ͽ�~�d��5�R���f�
\RP�vi,��Z��Z2�0�x���k�r]{��̇�>
�s�<F�>#gG�7��^�����*��:����~��������M�y0�(���~�T�p�M &�U^]�����A�'v}�7��uP���|7~ڿs�:��۸̙q7gDB<��_M����L�ݞ���X8G��.�{�l5�U^
���.��ɮ۩�규����`T!UN���\�3�aN����t����MS�=�Ƒ7Kn�>������A�x+�)r`X��,Xj��`�Ѳ��Z�e
� ~�|�ߏ�{�s=��"�;���dϵ�Ǻx~N���c0���_18�H1UP+�Mv�0vџ^l(՜�E�\�*�ת����ĥ�ۑ�.��5�)���I=���k,�u-� �hҺ�����u�)\G*5�Hk����}QCw����[�]�6�=��&��/����p#��Y�zŌ�=�@n�W���Wc����v�$�Wo�J�Q�_]�]ۻT�$�8
��!<w����N���;��*'�p�G���P���7:��.�,0m�ZU5�*x���:������{�6�= �	��&��B���uV�K�+�C<_F_���`��]�e���1�Q&�b�]�\�$ ���;�l�b�{��UU��z��w��E)��˳:�/��Ծc��w[HW4R����o댸z�z��rξ��=ܺ��Y2�p_�b���{�o�H������_�XǷd�N���	���])��̸T|Զ�Jd�]B�^~Xk1�Rƛ�!٪'�b�8�C��u����cmN�&^έC;�/,�pc��[���o�R�8�v+�mq�#1c:n����]&��ˠ��׽�p2d9D�L���td^R��5��ګ��W��7s�h��Y����*�y�)L�S|�6�W�m6I�v�b.u}W2���uPpv7Uyo�k�ڭ�]�͛�޷F�j\�l\��X�(��g���_!�kO<u0��u��E�T�*���͊�`�|s�h2݆4��
�r�XPR��d�әskV�����u�ܳn3b���W�D%�p�ȍ��w�j����J�̏��]�Ckpd����5,���i[	�H*;}"f���F���w)耜�en�WV!uo��;����p^�ܓ���_o�����3�m)t�U�QΊH7w�j��UH2_`�����̥	�*]s�L���)�Z��3��ٶ��.�h�2T�՞��]�T2�^�cIy[����ܝ��U;;��m�S�2�Pc���5�zM�d�]f<�M�wJu��fP�2�,���㪦���5��y��*7��b�P�it��U�3y!� !hW�x����J�;��r�8�w�cԏUdtA�co^��{����kն*5��o[7���e=�j��(���UHy�V����"�^%:�H�^�-l��0PѺqe���Dr�Ru�aK(f��2����,Bk�:nRE�>5v���_"�^n�V�ӵo~x>�\�T\d�Kd��T�8�X�p��"�a*���HBl����	0��H�Ɖ�<x��:�"8./k1QAOh<��e1���t���Ӣ�
��������g��*l�ċ�7lIlSQ���Q�#$$����Q&*$�8�i���zxt^�*�d�2��������	�r���Dq1��hUpAyK�(�8zt�����Ez��
�
���1�n�M�m�����S�|~l��咽��N'9�ENG��<;���uM�X��I��U���8���̈́�I�)���)0�ӝ�χO����/v��ZLl�qS�NR���v7)u!�Ͱ���BpD�ӧ�O�s����5	�ս@�Ғ6�n ���Y|�WY��N���p�#롤zz|><;LL�QE��F)nm������s���Mw�PJ��,�#�ʧ[asХ�xPcf %��l�C]� �oh6���1�Ғm/@�Iu�	�}8��H%������f�];�o|V��ע�	����B�UQJhv����SX�[��]�˿����m�S��c����s%I��n˪C�w��N�>��4���ܱY����;R�(އ�b�
�]7f'{�Y�>�}��kT���f��۲�D�F,�͹�Y�J��a�IAn��������U.��ד�#���4_'M��^97��I"C[�����\j���cu��y����m~_o0cS�~
Oh8#�n��33]�xJ��n "��>UP��{d�f:G��>��Z��NSo�`9UῷF�@]�.����zAq=���Ï?�R���y0�����|+��zFVo��p�����-�Yء�TA7��T�ص��⪮V!ٻ�k�v���i���T9uL�J��'�D�(U[	3zP�
�l�GFZ�D���!UO꭫�j�t�p��J�w����x �����׷hI/�LN>�}�F��v*p1	D%�8(��Il�,l4���Q���C(H �����!(p�G��oz��v����v`������:+"���u���;��n�ݿ���Y:1�G����U�'�����e����;���E�����@uX����8�z�e�|���U:�U�bvj֛8?q����꒿��]8 ����]UL
�.�	��	d9�l�/
�;K�T���������tVE���>���й�~/g{ùgW~����j��X&}P�	�k�l��1̨�'}�����r�ݮ�Y�z2�g?�Ji-xjU'R<�����C$3��妃�Y�:�u�ɴ�q��k���;��L�F��p��ya��f�C(��;ziqf���N�M)4~I��<����kR����m��eJ椵�Y���uxD#�U��)LQ!�Du��$�a���3ձVT��8�] vcM�W0ۋH&��j���/#.	�\Y���j9!ɂ�(X������8B�RkX��([˞X��l�l[��e��.|����b��ic5I�@�d�]�a�5̹Xg;���)Tպ>�����6A֠h\Wp�J�*�$�s�u^GY�`��J!��~��U�{){����"����Uc�>�nL
�Vc�_�UQ��a���,T�R��|37�-E�蜋�@��c�W�������h�|�m��r�[�d��>_g߯�n%ʢe?b�������uUQ�U<n������������ُ1җ�o����W��}��BspP�l@�c��ŏ|��v��v���Z�Np����g��_������$[W����E-�燉>���_wR2Z��Eh\��9e��% �v4!Z�D�j�-6�5
EGe��|"������Ϥ�r����{��&{z%�Do.�6�US���T��o�+f+I�0����e�ԕ��O]���[UPJ5��[��٪�pX�������񡘩+��Q��� mw����)��Wݢ�Ez�w�(]���oto��@1���U/����O�29.�]
����E���/��RP$�>�rQ�bП�ۃ�Px>�����@9Hmgo{�R�z���_{���9���c�����p+�U{�U�B��"%/N��5^n��T�Q�b%�*ת��B��z�n�|����(B���P�����w4��PK��y��u�R�6�)����&�!7ִE��ʨ������xs���W�P5{��(p�4���9��v�^O�D�8�	��Ϝ���}sY��Jy���Ѣ��%�T����(����O@���Z��w������޸������R�f�Pړt&b�-�ҤJ��J���X���Y�������cXի��wd¹+��*dq���ܺ�Z��<�1;���E@���I���j���U!b���1�Q�+�BN@�������������r��uh|��U|U~����W�}T���ݷKܹ�b2�_Fl[P�gF o��uJ�|*�����:�Ǿ}ץ������@�l��J�c.��+)K��b����|B �3�6dR|ꐙ�-�R��y����g�x�ʞ��g t�����&���@�j��/O���N�BsS�<�Û�9Z��g�y���W�/�9]olE��0^w���USE��@���=��2��n�tFY�)�������w,Fx��sӳ��hf���)f���2�P���r�u�>��f*��E�lN�C�ɭ���R�/P�h��f�s'	��Fr�����o&�S[{`�P?N�q�$���wx���V���	~�y����UT���}U^W��Gu�̚Z&����h��V�s���^����RBksqvߊ3a7��A,�D0ɂ���IM,q�՛C���(�T؀Kl����
��ｫ�ww7}6��C�Ζd�8�%�B���Z���n��U^"�� �8>��+����]�K����;6}�=�{��v���bumNvJ��^��n����&ԕ�&�����1����=\mڹ����`9|��b��{\�^��d�K�<&�	�����6mgf�'�,پq�{��)�W/`��+�N�ҳ9�/��B��V
n�r��`�:�����-���}B��5O꣔�=����m���T=s؎̷���"�nY2�����]��#�wf�ۻFM���A���k^���-)ΛUD�c�}�׊z�֪�����7�m����I[�z\-/;@��AĦB-u3
	�Sa��\�y��5�aig�L�C!�Upkκj�Ak�uf.]��˦�s@���h�r�n�<���]�,�]�v�� ���ܤuf���1�M�3MV�4M�g�n룆kX�M���R�l�q��R��d�kemF��̫X�!��v%����ֆc�4
��9�J@�������K�ň	u�]w!�M ,4��
�ːB�Lٰms�>K���p���rJ���љ���������.�+6���?N^���wux-�0l�3�2��GՋ�[X���?m��Y�ۏ���32#���[���2�4�T�����K�/t�����Ke��l�C14{��0�Z���T�U?�������Q�6��US�љ���������/�X"R\�z?�p�}����	d�\�]K4�~��;����n�]Y.v�N�� Uz���μ�ǨwvOt�ܤ,��}�V|�Pk��a"��L�$���a�W�ݫP��g8��"
e�
.7���.�`�h�K��߲{���=�u��t�޹]�Ȫ�w7v��m����*f+j�LuEVY���⹥ܝ$&V(2��2�ET'�������s�9�u�.78ݝB�Ԭ�2�CT˫�9V�|7��[��n����������ߜ .����}����}���u���7jJ�X��exE6����d�[��s��p\/b�j���?g䵜}�m��|������r]{�d��C1t{�JN��u+а;���h1xI=~��$��������}�owx��s<=q[0�/�]JI� t��@S��i�|DD[h�?p��0L�k���Za��.�����
[��nLz��X�j�«&�n�}W.r�N[V��_��������.� ]�.�i��}ǯ����U�%����Oh�3G����U�*�ſq=���^O�]���UHxT�+״YXP�R��q��""�'����]�M������[���M'��j���SF��8�>&�]��Y����83�z�`����?�q�U*�UO�Ol.0{�|�w1T��.���T���VS��DSݠxG��|�o��w����wn���!��J*h��:�_G��;���]��`"Z����E�*���<B�����-O�\��L�H�0�`���-V�)�Eiv2l(��pKf`AM�-�{��U[�k3�*�u���=�켌ױO׺ _
��U{�U��|���B��yT���=~S��p_}��^G�1fz]lr��E_>�X����wl]�w#���{�6NǪwo�;�+9���ኦ�%��!;W���-o��Ew�pY��d��#���8-�W�1X�h��������m�,�����jë��	qf�(1;	�=�(��b�1�+.�[{��/F�b�NtJ��w���e�E�	���wרp�����*��:N�n���#7F3�ے����*���}T��M@�^�ƃ����>}�������������f�	n�m�\�v�ѹ��a�P�P�4��S�9�]�wh;�Z�=�������w��Z9���x��U�o8-�o�-m�N�T��`;B�^v���z�]G\_	���@eӪ��E�A3��:�6v���*��\!�+��>�������UY�r�`�����*K�%�}��<�kd�j|�����/�RgkVǽ�]��>�=�<�����%�c�xU0�C1fO���m�����Dy�̊�|�>V$b��@��?/�^��*��"�(��/�!��A�����U �<�� �2TH*�
@"�Q� (� ��(�@�! "� ��h�)@����  AQ` DQ`�TZ ����, ���*, ���
 D`� E`�TXE�XE���E�X �TXE�TX �X�TZ�Z� �DX$�E�X E,��TX �X$�� 1Z�� V	 �`��E�TX$� EQ`�D` V� �`� �Q`�@j�)!! �T�A�A @@_򛁦��@U� ���������������s����C���9���������ݣ��J��+�3������xI�O�(

+����?����(�C��PQ_��@~�������?tO��?3���Q_g������A���?�c�����������p���,U�E��X0 ��Y`11X�F$Q�AX�XVE@X�VEX�dU�Q��EY $P$S��QE���*,���+�, ��*� ��"� � +���," � � ���
ŀ�*��R"�b�*�",X��� 
�b,��B"ĀD��
�b, AX�`"�H @ A��B*��D��*Ċ��Ʉ������?�AA� R@Ig�|��>�9�3�<�~P�����R ��������~;(����t�#��0��h��(���A����C�����((���(��~������J�(���(�,E��O��O�i66���������|?�Pxj>�<t;� ��������Կ��P�
+���
���~G8~s���������������|
AE#���(����� ~����<,��-�G���]C\�#������DWo�$��_�ɱ�)����gG�AEH���6��b�(�O���>�>?��4>���(+$�k#B�㠨��0
 ��d��C�!E @P 

 ��%  HU*��J�(��D�H)TP�
)%��� `
 (P��$R��$��J�@%@  �R� � � %��(J ��U P�(I����T*Q%U$J�R �����*D	R�J*�%ID�T
�H�*�$�B*��T*TJ%UUHTU@��>@�	�%@�
�JUH�w���������P"�@�ԕQp M�@� g`��� rw$JX ma��=r@
IE}�  p��  r���:
����IB� � �gD{h( { �<l��Ǡ���:*`�T�����:
Q�t
݀P݀���((�  �DP�)EQ! / G� 7`q7}�!���RwR8 28��A\���hR�x�,:�{ w��� $=�   q����w}�缢�8Gs @���җ�����I0��dL�; q����QO�  �Е@T%UJT���� oI� {��9���� ^tD-�(s�� �`�����D�p� �4J� P �   �레��yV []�ϷD���J��B�n���r�&�' �D�R �|  �QR�JJT���R�9�KvqUW�D�nw:	Y�"�I���-B�n�$�05E��ur�R�h�AE}� � n���� � -�T 9 �8@d�2 [�R� �@ b@G=�P @| �`3J��EHI
U�I*E>�gc� ��ް�gz���D�nq�@z�`@���`�r��_l��}��P ��(|= ^�� y]�@MȨ�� �� ��r���� ��!
8�ݏTf #�@�OM�J�1 ��b%*�i @=�L"�� ��R�@  OҤ���0 I��y���O�@������Z޿�$������B�yAӔ~z���4�O��I;�7� !$� HI	�@�����D HI	���Uu���}������魽m��������n�Àg��9�y��uqPDA��!���Z�n*7Sh(&i"d��v�aB��R���{KC/^��׻t܇[f��xƢ�z�di�B��]�F}�^"u� /��D7�:F�Smv��/3hC�#T�b@�n�ȳU�b�!�M�4n�E�^�iB�ԩh��w��&k`����ͽ�8����\��/7�`e�.�X�cN(3��������H��à!`DtMq��ʻ��ԥ+� 3F4��&�K[n̫�����n�d
͜�ݭԪrnE%���nl��)9DDT��N�eAF�K�F�d���^�,U�b�Iu�-�%,�^9�0n���n�n�p"�V�+j��C7-;$'�n�8�����y7e	�B`�����Vk7
�V��+X�drQ��K�����.�#h@nm�QG.7��L%J�a���#o5]nB�}y�����{V�OD!���k[V�X�o#�F�RIܰ�r桀Db�caee�q8����[3�%�nY�m'z�N�@fV�׮H��vv���vd�޽q?���SK��bbi����F^9g�6
F�����iB�
�-`���t���ٙJ���%j�T��������gţk_�졦����CNXƀ�j�^��Km`'oM�4�D=���@`��l�,Z�I kh[�
3v(��̇qgַ@Q�at����	��OÃV��t��g6�nQ/b���(�(�;Rf\�� k��)m϶�ɸ�U�^FD�m#��2���UͶ-˳�n��aa~���9���^7�
��Ĳ�2�޶���k&�FVF�&^������>���7[˴���ۛc�2��<ˊ�!s�R�v�*��Kh	w�Њ�;YJ���b��G�
�RȐ��eLy�	Y�,ͳ01%n�6�w��r��c3l��PY�n��D���7Uk)k(�vm��2�k���Дn�C$P� �.%_Į�)�W��=�њhUռ�����漬ق�E^��u�F�f��:86ĩL���c�/]����.����&�	,���-��F���m��r:fXYJ`�Mn��ʗL5��/.r�)�h]!*���"�Z��w�H�8X�� �eTA��!���U�į5�YvƊ�����MC`b��k %֥z��4c�$b��kh��bb	S۴���� ۽Xa�dG���z7�5r�d��YQ�QeY�A6�A��lӡ�Q���u鵈p팰^�Hdn�y+if�+K�1
��%��u��lm��@��6��8�T���8���A�Xِ�c3ND��@F��&O	[��f�t��9u����
߯$�X�o ��i�v�PYs~�t�h��Iyu���'/K
�me���F����]ŗrΫG�fT6K�c)�"-vݼ�q���6ڼ5l���ۇ	�4v���8.��[yH�:�أ��4��,��fb���̸��(�V��)�{�d�f�FV�M��5�F�{cXY�l�L���lڎ��a2��L]H0�ui�<��
"�th�i��fhw� ��'wVR��|�Wk�z�V��œO3m�7S`�W2�l��Ɣ�kE�1PVh�˶hXRеk2��M��V%=4��rm3)�V�8P�F����@��ĵ;tjL��V�ne9�k���*�G.Q�]���ASj�$p^�cƪ0,vV0b�6VC�֣xN){�2e��Eh�]Y��
�j�c�V���rD^.[���j�C2fm
�\m^���2�͵��1XVfe��1ʆ4ꬽ�"�5��Y�AӒ�@V�!�b�+����k�e�ڼJ��@�܏0��u�,�n%� �V��V\B���X݋-�H�H#LM��N��5�3I
��V��6'[����-��80n䭽����b[�r2`��[Zaݹ���P%�2��@�U�yR�i�l�k�wtVMods5l�B�V07��ؖ�A���6f���m�����XQ�i�*U�=�ݺŗG0�@�YB�dV�Hj�qm�1�r�\[�{���e��Kph��$�"��-�뫽���,i��0��ZI0T�-:pG�bS٨�� ��ҁ����Q""�j�#�t��sb�鸎ZU�[�ڨYǐ�,�ҩB�0^^Ьћ�Y5)�C&^���wګ�gfm#l�A%'%��rhl���@F��`#-3[�D��2���9��0�R�(Y	/���R��l!RZ;��$ǘl�u�`�p&�h:)���;uŲ� �R+�Qa����5z/e0ᬐ��L�����I���#�n�@7wAbfހrŪ�&ͩ*�Ȓ�q20�?KN���nd���n*i˻�go�h �s3:om:����:3k�����@v^m$[y���靠'�i1�����L���e�R�79R��T2�Hb�I)4A�3��nڰШ�f[�p!=�����ҖT�X��ؑ�M�F,���a!x��m��5q�N
�)����t^O6�ܴ��Ð�R7�$���W����{�z�� F0����e[�;��bɨ܊�.��]A��f��6$F$RScx���t֍[l!�+Yr�m#1+�je�,-�Hr����E"j���J�5�q-�fq�9P&�D)��*z0]��|E�����s3.+�M�)Z٨�+b����֝��5������&s*xY��؅�1� �b�B���/+Y��n���&�Օ1�������n����͎�0��wv�Q�f`�ҵRA�	c;��(5���!Z����
��˷�(Jk$^�U�mI@�ŨT����4��2b�}x�r�$)1aR�,<rͅ"�[��k5pDJ�������477�G%&�����ml��6«�c@���60�Y.��*��x�ܔ��X�p�w.�f^��n�[x1�����rqTE�{�&��^S��Ĺ�u�t�u��X]d,��V�M���Z�]� �Pf���N,:$������)T������Ұ�]n�z�n�@�:��u�e�N�[��z�&*Î��J:�eaq��ʩ ��m*�i�)F��]0/pa�X@;�c������eD�b���C�f�`��Z��0R�آ�=�K4��;k��nӑ������y��c�x3.FՍK�K%[��y���B�,tYߞ�b�&���6$U���6�ъ����� �oVn�����Se*�1��Rb����ٰ�d��1�Vr�kڳe�gn�twff	��I��u.�[��q�Y��n�֎
�
] R$��D��5��*�%Jx�����bj���eA����4f���dӌ��T�h�%A̖/�u,�Ot�EJ��iZto�Ti�Q
���]B����m���q�ɷ�c��%��[&޵�K[n�Dk#�֜��o6駳e)�0@=*�x^�´i`ə�@sX�/&�8j^+W.Ψ�ܥ�Z�4���.ݹ�cR��ː�p��a��HF��')LT�gLY�fn�O�]7t3m3Wb��U.+m�W�P���`x�W��`9��Zrآ*V-"ZR�%G����ť�"�EI$�ʜ�S"]������T$�PPS�Z[xeMR�J�*X沰�rBU�M6w&	30%+lI�nA�JYn����+*]m���n��4�W.��q7.��m��	�{D��j\%&!y����k"�HSb�b ���x]n�6/NJ;���.���̒��g(�S��4�6%^���diU�֓���nZY3E��Y%i;0֑v�-u�j�6��c2�+�!�b����]a�b�����#YkV%.X��U�{���Fܰ��iPCl���n����- f�L��tEVԩ�*�v�݃jZ�a�h��@�*�T�"ĂEdոʸ��[��קp���S�.�XR�ҕ�73qlv�1��b��bǨ;o`�n��D,���[�&�v����f3Z$�X��AO�f� �n�Ct`�2���e �O(�V��(@+6��"�D�edʁs
)�Zn�	
p�	���T�MȲ�0 ۦn/�5NY����6��P;��v����X`�Z��};�\�k���)�
�둊��a)\VI� ��%mS��N(�LF	k�cv�̂b��6@Uʑ��ŕ�N `s+[�Ι�P˻�J�!�e՗O�{����YJh[����{�e��m�AG���M"��&��hm�KM՚�7!���]��om�6�aNԤN��2�7 ��⻠r�֩f<M�"@u�ժ f	YQ��٪X��E���p�)�I�aܻ��Ax��Q THU��u����iT@�Z��݆�f�BFJ�L�n�,�������6]��ːnj�
B���ѩ��oa�`�ܘ*k����֠��h��[�� ��Ŏ䫨�T���X�A!��G���Q�2��mhbƻ,�dY�2�Zj�6/%B����1��2
qI�ɱ3jI8�ti�4�NXr�^n@U�r�*U��<x�8.��FnڼR
�kJI�R�ma{�����P]֥��N�Jq:5b��^g�&鳲o˂�!Ⱥ�̚*�D����R���z���RYf��[bAz�Ŕ`�X�8��Ǜ��~��v�Z���f��X8�	�jGT�4�/dV�Y�\Cl];YF�f�n���Ae�^�g
&�� P���l��*�r̖���q&~�T����'ecVpK�.AT.�`�f�4�7��LeD<ʩ�ݽM6�l-��|.�D�V�l�w����Z:�f<2A�����HT2��S3r�R�
\J�bS&�քLz�ջ���R8�Mg �� �]fd]���h�;!�X����jP����/eC>�N�^�ԢZ���Z*΅���nMݪs$Z�n�ƚ��B�V�\��ؕԢ��Eӽ�wƬ+PM���VL��m�Xq�Kih����0�V�3A������J�̰퓻SC��b�ypi8��џ�� ��м4I5�2Qj���Ĕ�$���I�˔l�-�U�D�Eڵ�s@;�h؁�r:/E���F2!�{vH�3UEe�����ӳVSM�
9��-��e�0��da��.�
��Ye�b6��Br�ݦ(/�E��d�%�Nl�v�nݲ	�� ��[ ���t!�p�ԍ=�يY5��A�(�0�U��KhԈ�P�J�攐��J-d`Y�,x)\�B�^i��ӗ-]�����fO�7jM�.��k	�w���#i�
�^�D�6�y$�=՚�	3sp�uf^jt�=�YWyoS��nݹ��̔�D��5E∣H:�![e� ����QoVR�r�*�ԽqqL� �%x��]�Bm�Wxfj�F+��Cw3[�	��Uj�SJ�)V٩@2-��c��i�z�Tִ����?R��S��h�-S�EGY�M+YI�c1a{�'�#"���[���6��j��*ƌ�)৓P�hL[yC�"iW�!�8%&D�F�/Hѧqǚ�e���N�ɋmP,@C���h���*e�P�U�d�!���aZ�ܬ�`vi��Y�X)Vyv!	Wr��X���n.�VTS��S�&J!�˙+i��ˑ��i��N�d���2Z͕�*nȄVN=҉	X��\��$�v���v�a⻭8�d�㵪KX�U�3j���h����R�}����b�[F����ò;�4��4��R[�>��-��o��wtR����^Z٩���e�!1т��K*����:�ȝ`��i����]-Y!���N�9^��E�P��Uic��gq�PMC�a��w�^�v6���ȴQ�>#:5U���E��r�`�X��e�T̫�^L�R�u�Y�f�Eف�Z�̖�7X�A�@*`��� Ǳn�X�S�0�͊�J��^��Uͷ3t��f�+_�J�6Z'JCY�V퍨�ڙsL$�C�ɢL����E�9�f�U�X��YkEnQ�S�2��c�����0�"�v�S�
�SM,�B��XK%7tF�j?
g1裘��.���,M����v3�L��à5�$�x^eZ��:�YX��%E�w[D�6�@Ah붙p���U��EM�)�0�&[�"�z��^��aiYWM�h� ����m�`]�D�s��D�Y���W�)9*CP�\)��c�L�˓'%M`S-\�0�**�-HH31蹜y��ݙzj�2X����p���MKۣm�L�.��I��n���JUTf�ne��Å��mZ3�eȪ�vek�L���I2�;���U�o�e��"P)����חV�x�C\9m���ώ����Z��Z�GgJO�tĠ�ڼ��b=�%�1��R�5�}��h���BX!��8lݍf�$�tb�:h@v���Xɔ�EK�W��dM4U3�D�I10�B� ��މ6ʷ�#u5diaQ^�b��;0ay���;e����ҩ���Z�ˢ2���kF��>�0���*Gy���Yc� �u{�����ua�Y��%��kP�)��vb��$uۛ�0��֠�3���t�ؖ�x�.]��/�	ͣvޜ�!XSy!11��Q9V��nbYw��,4���6�7s�#2�LPƑ���4��-"�+�Mæ�zX�ʃtfj�t=ZZ�1c^��k9��F�DS^T��X�x��gY%ǑӘ0�&n@v���l���gwW6c4�Z�����^\Sz[�h)l��ۼ���2j��$B�T�l��wV��MA��ٓJ9Zq���J �J�q���V�7jJ��1,����#l��?-����K����Q���+����,�en��2اEZ�72�$�4�ol��X�.C2��PXv¶��%��ik?�v���}{ݚ��!��$�) � Y 
@Y	$�@�B ,�B,���d�"�B$�),��@��
�H�E H��P"�@�@��	 �,�BX@R"�X $����a@�� �$I��@�H�(BA`E$�H�@R �! ��!$�E$$������� �	Id�
@ ��E��	"�HE�@RI"�E !"�$���d��$ ��($YH� �I"� ��d �E� ��) ��I$P	I XH
E�BB ) ,�P$�H@��,�$RRB�BC�  BI�>��U������53�(�w=.S�7D����}fv�J�D���Ù����]�]�(r�Z�ao5u���8uA���c�Q2��g�y�e�%.��r���3/2��2��W\����T�R�N@��M�{C%�ڌ��wv�v�������#U��ki�UMV��������U�p�Fu>���C(��fq�^wv�����Y1h�`�:7�p>ц��{F�R�'SY��mᰍP�#%L�ґ3�-�R7yyJ�f�;nNx�ʢ�v�2Qݫ����o��9��V�ݖz��m��p}	\�*_:wc8V�j�d�x�L	w���C[6��㴮v��Y���S��yE���dI"��U;X���Z��5Q;��W��X�J�~���oC~ǋ�Wǵ��8����v5fN8PԲ���ζ;�*��q;A+�/;���V)ޚ�x�oŻWR�]@�"����NY�/5��K��[zH�n�A��0c��o�y]��.��W��8ǜ����*J����:Qs�����F�5͌���l�V��G�/ΫV�E)7[�jR)KLk��L����[�U�2�[�+�5(����Kw��Ѝ���Ow;�X�,vƛٙ]Y,�9 �br���	����e�g���:d�;3f�0)6�R��m[Z'�;�"�Us}�[��ij6i�N�a�×�ѳ:W\m��j�ah��c�]������(�P����b�&őf�*�g�^�J�5��ZS�5/��Ð��kݛ��Ì]CQkgCVR�����9~Y;IB͈��0�Ɣ��}���#���F�<[� �������N�tD1uB�E�,��vn�_.$L.�X7���������[���Mf��a�r<#��i��Y��+���"�lؼ�E̩�kh��g�5�mo�� npn��R��y���z;+1��o=�i��IY=\��h<�f�&��v��vN)9�Y6Z��/NX��dW9�@�V'Y�1_tz��sa+U₷��xQ���]��w}�s��(��ʰ�J�;ג����I�m]$���*��Nр�w�a�fnG�J�$���=�k�b�,fgvR�mn�
�o6�-�D���e��\Fe�c�*��oBHս�Cm�[����g;��k%�JOmE�k���d9˄.�iݼ�A�k2�N���8.���If���:��d]���4Im�b�
�}�I�uh� wK[c4��X�V�b���2\�j���I�X��cnp��h��L��$Z���UhK/<�9Hc���k��6v #G�ȼ��U��O(χĬ�Ų|�inw�rZ��t��Q��̖j�}���c]��L؆�|����ަ��ٖy�˛��d"u�j�ධ���i:̃�cd3���R�)Q�ppűV^��YRLlSZm�1!)�qI�z^�d�Csm�テ�nՕ�Rv>�K������f��qQ��0�l�8et������B��wpɽ��q�ΨV&�gg$�\�j�q6��mE�o�F��K(�����
N�Μ��nk�M�%��?j��ֻ�u�����ɻ�w�6�Y�6"5蘒�
F��YP�Ò.��g����7� 8Mޥp�A��1�C����Y�7"9(t$��sO]�^(gCN�KN��B*�h&U�&Q���� �r!w]��43�=�t`�S��`>D��Z������^�k&jϳ.|�Ru���i�N�4�D�kv���Z6��$r���"`�m�ސ�ے��W0�ެ s�*��&�_Rt����T���hʹj��Ό�I�S`�A�E��<y�w;.�hr�U�ޮ2���eoc䙬��]6�k�:һf<�΅�AiS^�s��s����ƻp�Q��l]8JW�3"�K!��$nj[���{l4$ak+EyF��pK*�C0���.�ho`�P��h*s��޲��˓c�̃Q�6M����P٭0��wm-�w&dR �s7��q
Ф򄭫����9�݋��-�����z.�:^kʁ���M�<$�d_����۫*2��F�P63�gZyz$;uY'=��L3VX��;�3s�nk�)�֍��γ��݉:d]�/1:��r>X�"���J��a�t�1�@���2`ssM4�I���9�۝tLWHE�ۤ� ��#d��N2���x�V`���%�+�r�xΙ��v�^`��x��aÏ崩�!��U�n_n��b�Ӱ��j3����c6t���22���5�3ˡ���{u�2#2�x�[5{�Ax����+6F�f�l��$��VFj+n╹}Z�w%,	ǜ�N]�"4��r�z����^[�N�/v�Us���v84:�Ow0+��ۚ�����O3�z��T���4��uTPVc^%L(��.��gKQ]		��lq(�q���� /1�ɴE��C���,J��i,'����Nj=��(����<0��ۢ�.��W0�+�Xx���u�wcO!���w=�x�JJ���Ls25�CWt��,�.v�^LrOz�z�w�����(b���}Ѽ�M��N�Bc
a|sMYW3����i��[��k�Ys{��(�&�U%��JEi�h
&��\͇��{���R]-�I�H�����w�"�]�+�ח(ԕx2��T�4n�إ-h��)�]�%L�(��YF�݇(%[�^V5��gCU�ׂK<M�k�o�57����6��L�de]�yw)L���L��vj�+Uڷ�=��ݴ�	S�Jm�ϲ�=Qm�v��[�Sm�2��o��6�!nt�݄�7�����*�Z����0�=	��I��-�U�;-Y[��^�v��3PՇ���ß!(��u��G$j����9ωR�	�yKX�6ۮ�B��JYzw�v�<��G9dN��ڬֻg,����;VV�}��y���k[���r�<�%�;�,��{�.�jƳ��<qt샨*�<�N�~�%ա��uJ��T�-ۣf�1f�͹�����,@�(��B�N�M9	��{�����YfGufɊ��5�ˆ���J�K��8���⻕e	�N�_jק�P�*wl�ؕ�jX}Z;�5�B���]ƞ+.w�vWP'��$X���ߕ2:���t�Q�]M�w�p�ˡ��a�n�Ba�zr��ۙ��6���[VY�D��aHۦjpK��.I�)u��,��m]&���Dd��g�k�5r�jQvջU�������`ۺ�	nRy]w4�5t>:ռ�bXa�-���o	���j<S�Y�kN4�T�(;t�jȚ�C`l���;//� ��
��O���yj�Zo�&�R}�ҖW6�m�6��J"v#$ha;����xq]M2A7pcʜǖ�����kR[�=Ab�q,�H�,�W{�Q�h)�m�N"^Ν��Z�΂�(ƛ͓����nѩP�Bs�"kh�s3N�b��D�8�@s����a���Ŭ��_q܇��aA�>8Y;��Su,��P��R<-��A��cL���Hor�5f���{u��H[���&��vv�I�����#TL�x�;�{wF҂�M67�眺]��I���VCW>����g�n�՚zk�Æ��SE��3ZֵX�M�b<�$�%v��m��V�!K}uƜ����u�P�]�l�wǰE��ܶ���mj�3:lh�.�W�9UIG���9C�Rŧ�tsM+̼��^姱#z��7���G�R��,�z��^p�XP �΢e���F��B,��{�tv�XTɚ�O��6c�=Ib����C3'XV]*c;h�x<Յ[�J�m�r�}3hɡމ�N��]Σ��,�,i�5ܚ��p��|_C6v��ќj���B�X���k:s���Z��W����J��P���ޤԓ��>UӖ/"��ss��A�9��;r�1�s�V�Su��Y�Pd�h�y��\kM�	���+�f��}{m\��bg,՚�\�p���M�ں[��dV^,�794�n�"R�+Vx��w�T���1���G��p�T;��uJ ]>p�J���n����"QFC�}y|ḌƷL����m�	��%��ބ�,$m_b�mZͽ���N��Emt�k$��F�f��2��Jj�5S-mٲ��W�@�Keu��;�����'e�I��!͚�u��.V��{iA�Oj2s3B��	��m���L�k-b����0��r��hp���-�k9{��Z5zPV��h��JS�� �Ofvۧ�j�&wr�m�9��ƹ��j���.����nJ�����F�B��Ŷ2",b!aɵiB��Z��Ъ��ѠC�����7& #�5mF�:x雑�:�
R��V�'�I+n(��V��XF����kۏqf�\�Ɇ��_e��Q��YiaR���B�u��	��m<F�_gaVw@T�y�Ά&Eu���㮰Ϋ���ʎ�XJ=��r�Ui�q����j����{�a��.�v���똆�uB�F��][K��C��ve�q������Q���r�Xg�⚵L<���].�gvL�	`��)�����A���`���Y����{u~�3e��[��H�5�D�PV�|�(���Y&�u7g_1���=��5;���S���۷
��������ƨ)��t�u#u�B2����.�*WwdK�3��M�O��@��J�ڲ�Z n��5�b�v �:N�:1m���4���S|��x���ngֱQ��˻yԫ1�٣ח6=�++4L�0����OM8�n�u;pc�J�m,��ؓ�vn0�,��� �M�Sz�Ѵ�#t��L�����",C}gj�\�n��L�37�v�QY���x�Ճt�[al��q1��r;���i˒�׷����L(�(3y{xqĂc\]hsR�v�b�ֻk�4J��;��X��ͷ�����!YU*��-�˜�:�C��"h��r�&u�.9���r�i\�9�hO���od)��w�z�::��˶�B��GG ��ۄjκ�YD �x1`t��A&��ٔ���9��䜛,[r3�X�bWĉȗ�;`��a��(0���	��>8S��cnl�î�sf�	�!`����hU�U{#��ػ�`W3j�����J�����{.2�s�&�l��/�FK9ܴV��[J>�|8�	Q|빝�+�ZGQ0\�Vs�סn�g2r�*��lr�v=;-�-Aߌ�ս����v��PE�����Aˣ6��[W�(�I����A�X
յ(!ٕ��$�B-ٲ�sCa�A�:z07l	t(EBP��[���P�C2����+(&7v�DK���'��W$�Vj�F���E�nvL����'P��{�31)*����F��b���Oc<)����:�x�M��Ę"E�4��[�%�V��Ksr�ݚӥI*���!4���	*�ˌb���6��8�i�r�Zԉ�ꮍ�k&e�a�
��wj�g��Yk,i`��#2�uь����/n�ru1���<��3���6�J<άy&	w�1�v�=��Z30旹�\j��.j���ΖZy�S��L4�w3u��v�2��՚HP��p�e���v�5��3^�r��-����5d���:r���}s���]���E��{��,�x{6Y���oE�[ʙ��f1^�Uڽ����UjE��"�u{ܛ�;]Y�I��M�p3yZ�R�	��r���uY���w���U�kx櫕��R��W�:,ܳ�Ný�E.�5�[�VrY�,G���o���Q�qk��#�O��F��!�W��㬗R0Ue�R�镒d�Ϩ�<lW<M��Q��fC3ws�ں����=u1`��zV)��hN���7s��Q��6&$�jf�qk�0l'Q�I��f��h[kBJ���G��i��j"�eL�WdNR�#��d��1���\��F�EV�����3�)��_�WUC	��n<R��f]�\5:OU����v���� Wwzy�]��e�N@>�ܗw�(]���C���]	�(dx���s�� �5b�ʺ$�K۫��"kt����E�楷��˪=��^���+e�ygoa��t���y�(��M�xr�,y����X\�qQ��4`��k�]ڷ+_��4�K�����3��=5���G/~͕�\�4\�d
&�Z�#N����b�S����j���s0���� 7������V�:�����n�9�`���V�L��^���Pr��~���C�f�t�u:���[h�;�.ޑ���ea@JEA�l+w&�1!�;kȼ���z&����O���W�x�|#I�eM0��Aْ:��!������"-��o�7hC�V�r5J�H��i�Z�U�^_[%�w٘+	�F�b}�%�Z���MV��_��Y�)����w&;�2�9�t��`a���_v�Z]0!��ɠ�M�2Jdl[�ݸ���k5C��"�*��JbU̪1�L�P`��mc���������Ǯ�Q9%=�,c ֹܫ��-]ѭ�NL�%���+-���s*%M�9���^F�b�#->�s�{m��7أxŅ�;!e��k�u�ݙE���vk��8�'p}g���.�;,N���}�>��WxqSn���,�tV˝����I��;�[�1޸����m�y����K8�5|��6`@[Tv�-K�p B�*�it�
���G����8Ϻ�.����i���nM�c
�:+,X��J"aZV�%�[�b���b>�2h5�����E�b٭`
�\�������}�&�0��;t����3b��/[�&��0�:��!?,�3�٥�Vn��n]���{\94�8���/0Y����o70CGp�=G�qJN/;႞*���&p/��7z�;�i�h�NF���֞ΥkN���^�ͽ Z��: ��Z%��[�j<���v��c�e���Q6#� �y'&6���������/����'N��$�Oϖ���̪h�{][�ʵQ��ea�-Kc��h���%2�2��l�
6��V.��BS�R���k�](�í���]���0�B�j��ff��܍5p�Ls�c�:����MT(0f��fTڏ;��Q�]�4Y�V�șm�a0fXc7]6������T6!��b��rb��%�%�A�o��pMmq5����2��fM�
l[+��#l���Qa(˓:�
��R�:b�6��Z��l�-�������l�D�qf��j�&.f�b�ykX��m��)M��L��x�/�g����v�Kc7�p�92i�[Ki�B�H�W*cP��Mf�*�%.�d��0��kC�зi��Ԉ�ي�Qfs� �]v&k"]X��؂[�6,][M1F���3pB���r3D����G�X�u#[3�!u�D9�ؕĢ�q�ʤ3�Y�[*�'�ü�#4��Q�9�A��B�e��hlD��� �u��D\m8���<����*ZkH1�7(��,e��h�X�L3Jm��a4�%V�ؘ�)J�����m���m�YH	e)�Q�S�2��5ݱ-.�(6�ˆ-Y��Գ]���v�Y�:�Jĭn%.��c1t5��n�L�[T�h,E0%V�f���Р^��fj�kLV�-�˵n�W=w-��8��d��(Q�+ta��Y��qX��6�E�V��F�M�3]�ZZ	���-�4��lSn٬�1�[fj�a	nl�[q�q��4�p�۲� b�0l,Д�]mM�H��V-�Al­e���Fݥ�Ǝ��S+K���1y�q6���X�Q��̳@�5a\��5��nՓc�Z���IMv;k��p�\hp�͠�U���)�)�ke�����4�:�a�1(Ƕm`�\h��lcD�7b���Ԅ.���X%���M0�^�j�̛Z\�j�Y��l�PARl�\��ٗVe���Q]�ٴ��v�	6`���4j-FR�a�3F��`"I��q5+hKDV�bJ�ۀ���
�U$�DMͳm��r8�BSL�#a!]��;SD-��NQ�4��[4h��Λ,�b�k�F�n�h�!]s�3�aD�]����cI[�F�he�(���c+��L;�")-Z���j
%�ns\[�X�YCqi��Z�1�HS,�&�k]fmL.,d`�-�s).�%���Mi�,�ZM6�2�<k4Q�90 jґ�[�iGE�8�ЉI��"��V���Z�Φ�sQ)r�R[sb����eXͰ�]/W6�`
�m�u4q�V�k�.١��RUt+)i�UҠ�V���[���"^����n�\A8����\���n�n3�2��N��pB��mj�e�$0��q��b�aVj�Z3>i��y�6���.4�c�B���մ�M[����0��sx�E\l�#�s��n�B����
�0�RD6��i���18r�"::b�bhD�,i��Ƴ�5�#j�&bqS1��y|s����6.����@�56�©�5�k���������!p�7ki���ҍ���ip�l�!l��n��x++53S���t�c
a],�G::݅�r`�*�%(�iu��؉mE��������t�ƈ\љ�C[�K�v���S��v��u3��k���[
�[c���@�n�%K�v����F�a�f���H�U�:�̓�5P�B�����RĶ5j�4�.��gnл%�[)6ۘ��AL\��n/�(����q[0AKhn�ۦ틹�������3��v�M�.��A��	ru��J�٪���g�5��3K�Z�`GJ�kl�3Qlx�l5�%�E�̬���nv�-L�[�J�m��-ͽ�4�!cUD�Ŭ�[)�٤�h$7,�l�����W�vl�0j�1b�ه5�khK��bU-YP�`�5��[qv˝�)aT�ÑJ�L�"7 mPHe�llZ'�ט�����$�&�M �-�p-���;��%�����l�m�Y�:��.iR6&��ٙvY� #m��e�MsF��R	�`�fWV��F�j�Ε��a%�Ե5�y�%��B-Rm�,#T�^W4H���X���-c+������%Ֆ]3E-6���V���7k�#����k�����U�0���!Ld�nٰٽ�uU ��k2��ٵ�t�Mp��;A.�z�tډ�	��6�t���ӈF\4F뒅q�9�kD�h�²޴a4�B�9 �!e�L���7b��2B[�6�n��cTf��nA#�6��wn��2����93V4�(&Hk���!3n���v�0&�WX2�&,�.�p�١EY�[<T#O����y˺�cm�L�m
�ItB0ѮK��l&t���ٖ&ŭ��*6��ږ[7 mjC��#�.3A]��-��w(��������Q`7V2Ѳ�vmҕ�ɓr`1�30�\M35J�*��I�ik�fہΤ����Vә���4�V v���dm@,��h[��A�`�ZQ�[�]İ�ǳ����A34�c�D��X��aƥ���.b�L�YtZ�� kWpj�����t��1l\S]�LW[��i`m*�15f��ܗ�mĸ�#y�ݱ��U�Xٮ�W�3��gG���䖜%J�A�";�� ���ֲ�e�sJ�b����ˢ�Ěl�xr�Y��$�u�Űl&��eah@ֶ���t�0-"D�l�Pe`%�F[B ��hX�
�{Sk�����,O�O<������ �H�&�ê76��K-��1ˮ� ��K#quEHV:�����0�4����k�Mȱ�j��5o7`����fVJ��gP��nԌ�ffb8ś\F�نA{mj���`@�v��-�YS�� \���,��Z���,�\�
`(XԤ%��@Ii�m"��bhT�ı1���]v�i^����x�ha,��n.�Ͷ���Yjƪ	�85f#ka10�j8#�ī��b�0��R�z�jEpL�ka\Cl���	rjF�Vj"b2�&YI�KUahC+-��J��K-ɵ���[�R�Q�m���;&5)sT.6U52�ᮚtT�e�ċk���Sec��i��]T��0��\E�Fi����g��Ƣ�YV�+�c�Q�lQ�G�A��#d���1�ٚ1����])l��Ǳ0���]����Ggd�ٻ�&c�+u� h��P��Y���Q%0�i��m�
ʒ:��C���&�5
b"f�fv�ѹM`�&z�h���3X���ۀ4i����a����rhD�n�Y�����X;g<��[,�b8���!6��2J�2�u]x��h3L�̱����e��̩H�hB�$��Me�+���k�����n��v[�I����6n�q[qvK�jd�kV�BZs�цl\��JMcH�2t�e.m���4�b��Cu65�X�+�Yu�n�Q�ľqIa�r7*4	�6m�U��jK�Y��f��0�Y�˴&�ˈ�M5Ŋ(�M]*�&��D�^0��T�و��pqi���g�(l#6X��;b��TiZ莸3\�;`�#z�ڛX:���l�ι��]	�t^a�^�4ִ����]��Jb�KI��қ �.���J�n����w&)h�b�fl�GYZ�b��H�щ��(�h���i\�+F�.[�ܑ�#Y��\��Ze�6&΢��
ۣ���[+�a�b���-�QЇd42�Y��5�U+.Hu���h��8��Y���b�X��70�u���"l��lj.sSA����T<��	)|�ݝ,��4 ��]k�)Z7����;D՛��G�Z�5XE@v5
�v�փ�q�jش��[0�#yԢ[md�����Z`�2��6�-э�ЍF�,��52l�u�h��2]inke#�,��n�UI`�+�K��nAR�Mqֶ���)�[Q�he��gM6 �B�'W�0�XJmx��S������҈h��سF�S�a,�րl\��t0R�Y��ZAu�散��@<��])�FU�ض\R\�G[V��j���+DVKU H�.�-�)1Z��If��T���"�u�/*9��GT6tf2Zieb��� +�%�B�3�3cQи�,��Ћ����ap9�X�L�͸�3��.�*G6ͅ/X�A׌k+yi���l�w5��q�jeشԀ�J��V�ė6�.��WC-�.��ir�г�h�x�Ҩ�6,��Wi�R@�ҭf[C��u�)Y��9�,#��uà�T6&�m�jVEћ4���Yb�@�rı,�e[x�;LM����n�jAa��%��lSf��z̀�I���O<C9�X�[E�����. m�5�ô���ZB׆υ�&�4�Yf����L�3[�t)r���vq;1��e<_<�ۼ�G9Bxք��M�J�nԵ\Kf8�(�)�]C4 ��S3i�vH��cˬ4���[]Lܗ��Mv �%�����ڥt��Bb�T�%�@��B�oe��왽��c��tf���2�����r���%��M�ټe�l�WU���f�â�j൳v(ҹ2g13/=�Y���s��Ukl[JZ�6R�y�c͍��ljۊ:"Sh�tj!(R���``�*�Rb��U�"��]z6VP�!s��snp�tH�nS�bZ9lE%YbC ��9�f�C.�-zm�]3ó�i]��)aS.����Vn��ԛ��f�X�ݎ��LR�L��F&ZAR�u��w�k(�dk��R;BB�3��J2��0lM�͛X�j�ںU��X��sa��B%�gl99���:�.��ؑ�]cK�a�c l�A85��,�R�\�i�J�Wj�,6�:�&4��!��i�����f=i�T5��)	��C��i��l�`lҖ�cf����ogQ��bb`���sv��F��0С�j�^�/f�L���63hK�K���͠�Ć��f��e٦Y�1j�����2�m3m�m�!J���e���S�,��z^�Ļ��ř]�;͍���+Lc޷�-�1���&�Ec�k���%�V6WY<�o64�X{1��U0�U�E��jc�]8!Z�kޞ���%r�Z�L�EҼ�x%W��lKK%lkm�bYN,%���d��-2�4���YL����KM�i�����K*F+��%R�dXk��y���f޽k�͍���miձ�j�Mb˝z��Ԟ��!�66�J�=N8
�Fس{;��emU�-:���Ju������:I��)�'c�;{מ�޵�Ts9��q�P�{�ro{Y�Sys�����ա����fwy������k�-+h�t3V�&��w��]�i�ܘf���+1�mur[y��ST=y��6�I��`���<1�뫇
�fˣ���p0ژ�P6�J����wj�\���"�j�2��V� 20��k`"F�Bh���lk��1%Ͱ$�P���j�6sq@-�e�4+�[�4h�RV��hԑf墻��̅1�h���4	R����t,-W�F���LIJ���X�WV"��j��`��p9R�m,̶��R&�Y�Gl�:�D�2���u�γZ�-F�T���6$R:��K�J]�2L�5V�&�l��j��d�ˮ�\6�!yC�X�(��s��u5�ch:i��Lf���,��t�"ۢ[%t��`ˡ1ni."�4z���6�SP�D��K��6hk��cH4��0����rYpl�Z�Qe��X\\�3���ƜR�+�:1�b��.a�Y��iW`���hJ��en�,���2`��eF�}T�w�;X�m۳7T�Յv���X�ka�Q�1z�ũr[J
�6e��ݎݎW]5�Ufy]�j�]mj�q^fS�&�јe�Kfak+i�����ݥ�-sn��b�#�� Ů�X�h�`e[P�:m-+���h�l-���-b+��!Ḹ�[���G]eL�tH�B�M�閁ZJڻ�J˂�Y�\�u��|��iJ��M���JSF��mf�+H�S��F=	��).�5�l���n �S�uۗe��DmɃnu�Ԏ����ö����f̕�Gd �̄H3�hL2F&ok-���h�\ʎ�6�˴ե�t�VҚc�D	h�R�T��, \�pfS-�k^�Ų��j)��q�$E�
�m2�� �mu�3Aղ�ĵr���؄u4V�4uΔ&�e��R5���źS:�Vg U�U�8*�5�]��9�3���#M�`�2jpS�(�V�X�
6P�l�sn��4��Jʡi��I��V�fcp�⃵��Q	������i]�M�l]��I �[�9���-)�����k�V(!�cm�cx�c ),m��!��Ĳ����ą8�d)-��yF�-"#
������<0�����yz�xzʴs׼�R�k�W��jQ���Х�k�VJF���k�I��H�R�������o~�����\�#��f������*f���":��3
A0,�ػ$$WYP�| y��B{��3�M��
���ZqdM�B�Ԃ�N`㟫�}\��f�e����g9eǜ�E���!����!e�"�p�`��z1��PD�{� C�9�bێ�+tR���� ̀����{�r{<|�cx�+��^�Ճ�W��ܢ�C����*�^r������SKE��@^ � 9�x�����,�����*���Az#`��nFb�o=���f���dQ�2f �̉��6*2P㾍�~��`�Όs��5J� OtAב̄A�Bo�|���??�c�]
+�ڍ�+�5�5�X��3MHש��!���b^fs����>�C�#2�f �d��s��8�I�51�s�����c�7c�Tw�#�� �Պ����Պ�J��R�;������:s�x�D'���=��� �ge��������"��k^�bX�i&�bW�۳�B��\�I��Omʬq�>Az���_O.�3b���Z� ��Dm̎X\���͘�:�M�e@��D�f@@�B>́�ۛ��x��A]6/��A�"T;�c^G2 ��dQ�o�lgf��]IT?E�Џ��Ax��\.;�H�51� ���	���m��ݱR(�B��� NdA��ȥϙ11�rv�W@X4�]s�ۦlVU�Q�w�m��̄|Fb`�����nq�uԔ�T�4)e��i-��auf#�ZY�[�����[fbPީ�W۠��b&r�r�F<�Mh0]���Cx�K��wa��� �/#�C1̄A�̄ET.�ާ܀܍�_ ��\
�\7Ma�#���	ހ�6�2-�"b��J�T,뀈�Aw "�^G2و]�l�"����e���5�<�U�ز����:b�Ԍ�T����n�w�t��i��C�y�Ony]]�}q�Wf{nBJ�U������bb�z�{8�᎔��2}Dw���̊>̏fE]G'���H��_�9� oc��2k���iê�#x�K�'z ����s��d F�Fd/|s!}��̎��yD�����7��KGq��H�c�A� �6��̄A9�&��cS�tF��p,%��m)c��ڙ��q)a����SVV�L6�	���6ח�d"�$�A���{�
&)��]����U����"�܄|Fb�D��Sj���q?[;T(�W�-�F޻�5Czb R� N� �5�s!��l�=W���Q��d/Fb2(f!�y��eҮ��G7c��8W{���|{�"h#�|s /��иf��I@���s�A�h/]���twqb������Qcb����0�����X�뻲� ݎ��[����Q��6�S���0��t�N�m��|��u��i���|h�3�x�!g!�U���n� ���܉/L�޵�r^�����j�h��b���f��Az Xבm� ��Qqx���7՘��S�%�)B��T�n,�0�P]2L�kXf���il�r�=�����z��/�PD7 &܉ �Ĉ
�ٌ���f�8�(�M��$�Lf�d"_!>;��%�ۙ� J����8jg��S����"3�Gw9��Ȩ�>��> �A�tH�&6���K�%2$�Dw`r$�AnD��gu	�D�άZ�1A�"���z �^E����@��/%ho6��\=xV,k��ͅ��r'Ʈ&	V�n�([���>�k ř� nX�[�%��r��������fp`��o�����8�e�Y�\A�"�|CnDV�F �XY�(h���|���*$.���L+��zx�9��@��B�I�1׸�ċ��X�-��2��^��U�[�H�GP
�o{߽�zo��}Ԗ�],Uu�#`�p�v��/�jh۶0�P[���˯8��Z��)���iK�1���n\�!4#oS\r�WYlH]��ffl��8��u"�ꛍ�h�R�U���H̦�*�hM�X��]������0Y�����1�`������ֱ��.�Ʒ�̖���	�m"R�:������V�jMdTcr�4�TklV*2�֮2��޽�>JSl�d�� ���bWG��ΖX�9n*v�%f���;�W��K(� ��BKq�[����b6�[��w�).�F*'�EՔ:�Yiyx�R-��� ���!�������Wh�F�^>"�Ϫ�@*������U1��{�/C}"Kq9ca�V�V@D]\� ��^ ��mY͡tp�B�Ҭ���j:1��⬊�� �r��j���۟7|L���w�ȹ�ܫp ��"K�^ ����#s8tU�0E%���E�r�U�J0WK�W~�٪H=� n�ץ�7�!֞��U���
�c�q%��UQ� ���D�[�������?=�/�r`ܵ��v��u�%�� ����u,@�X�iv�H����y�=����ۆڒm꾁��GGw/.*Ȩ��B/Աl�f��1� ��܉�n ��5t*|�{��|!w��fX�c	�������kV�f���I��������7K�{�vzͳ��^$i���L)����#���{�M�3C��It��AƼ�m�Cr�([�y蛔�Og)�6�!�@��܃��u�՚�V�\��ʪ���� C|���ȷ 6�H�z��hM�ʀ�q�{Z�m*�'9�D��W�8��/�2�D+���i����l����n M�[��G��׃��m�1xt[5Ǣ��K���1��dףh����M(�Q��0	\00�4kv�5"Q�u�һR���!b�*�\/<b�IAh3A7��^���>!�>�h�������jj;�b�V�]�:�V@�A��_B��"hIn��v�17��.�hZ�{�^����twq��\
��A��> ���Ji�'яY�/.�s���s���A-������ft&��r�aN��=��b�����Ԭ�ɓ�����u�GY-�NHM{s��v��8���ǉ(�X�.�z�Ah��ڼ� m1)�f.Q"���@^ �kȶԂh Cp�(��*3�_O.�[@c�>>mȐj�`�U2������{�El�e���P=��>9�!�2�p�-�/�^u���u��b6P�q�9����&��.Dq�r�j�#�ۑ�1��>{�F�y��I	��Zsm�х.�hWc1Ħu��M���8���^�!�ݘ�={ч�w�Ulcx<*k�EA�zF���j��#6�I��㽫�A�"�mH"-1m�g^d�Ȟ�8-��J��)�'�75A�=� ��D��f+V7w1�G��D^j{`"� [k����ׂ��aG
�*TQW..;������Q��|A�A Cp��m	 �<�iSAѓ� ��"A݀f����cx<*k�EA��w� E���>۰m�ٻ��f��&L���rΆj�z�:��y�p�6���k�#T@	,*�A��׶���s���*����>S��.�ڟ�C.�7P3é�=w��WB5jb�}�iǊ ����"	e�����
��{����,%�����5��rfesZ�٪t,Gm�-KX�#�	B]q5!}O_�۾�#�Y��ϋmH ��Mi✸���M��\
��6�mb�nN�C˴�"�� A�"An�
�+o�sW!#+��g�`!�f]�e�U[��w� F8���r��e-yPGL	WB��H!�qGŷ#�L�y��۸������}YU�=� ��Ȑ[� � 6�Hۋu�Z�d��y����R�SZx�%���M��Z���)T��o���Z,��{"|p��mȓ���6o'e�Ajs�����1] ���c�!��R-�9����0bҸ��,���=.�v�B/8kK�������]K9�k�W6�a�a��8�78�I	���_wU�՜6�9���թ�n1��鵴�%
`��"I4G6��3� ei��q�n�k�	��K�3����X"*�Z�rU Ms�9�5�����WPR��X-[f-�(`�bm��M\3m��P�cA�0�Żhj��*�:�<E�Z�6Ƶ�fa�*j�7�ŷq��Z�PH[d�n�"�e�H��-2B!��B�+�dŰI�Q�!���m�Fl&�1�T���,[����p;翡f%���p���0����]����6���F�C����޾��Yd�/T�Gj��mȟ��]T���'��ɸ��V1�vM>P(�*��=����w ��EoF�(�Q�����R sAMq✜��ޛٸ�*#�%�)#�!�������Zr$�G��6�H�^ ��l����B8���&���6I+����4m_�>m�Cp�8A��L��WF* �܀n(��ۑ �Šy]N��9��'� xܝ�`C!�9Ј ��@��� �Chڽ��yqVg�p�x��8R�|y��n-
��	}�ݰ,� m�<>���������ٹ�H��[�(�,ܙ�fH��ݙC�QR˷!6ͫɯ����Y��[�"��bU�5��q�H1]#��jDN;ń��2TfǑz�����7@�ԑ���狸�h4�F튽ʺCs
Cu#S��'s��ϮwW��B���&h]tL%c�kM�"u0 ��;�:�6��T����Xm�Z���l��-�oj;�Wz���	ހ�#�g�â;�o(�D ��|��� �א-�$�����ll�*�֗�$��Šn8K�RGlCp��my��DRl�f�B�[J��@/��^>nV �_M�����A�� ����4b���ޘԽ@�r�� Cp��mH7�V�vWW�T��9��qH�٧q�n��Nn=�z���� �R_9���L�D��ʈ17	\Ym4�]���!���M�!��eu�(ٺ��V$s  A�^^-� ��)�<\�f��of��7�F�\W�fwy��A;a6А[�A�n�A�}+��n��� ���vb"����ƫ��A��>ހ�F8��m���Y�����:��\F�e��l��j�=�u!*��~��B��Gƨ3�Q���N
��ϵ��Ƀ/��}� �o)��i8��taP���	,��E�-���)h�� R��{0\n��8�Z2"���
�c*�ꓳX�"J�/���Q��8Z��6�H�J�Q]���+^AW��N�ʺ��En�a���n��$شJ�X�ǯ��]6 *<to����̅F�q}�ڥ@��Ҿ4:�2�mI��h;�u�+t�+ͧ�8��3Vl��ꙣ);4x�y��[׹�dź��{	1���XR��J�+�m���9�#i<�x�t91	����b� &V�}f�h��|��O[tO
Lt폯�����ml�m�a{|��C���*�R͝����ot�b.�R;��vm�K0Nfފ���f��j�"��p�
^�c�][cqeh�"��ۅ�m�5�}B��aV-ۍ���UX*�k'/f��[Ul\ܩ�:c'sb}b�
f3�n��!��^VX0�f�4�Ѻ{p�.�XE����E����[-�E�+fo1Rۓ�����9J`]H�u�1�v�e`z���� 5��.M�ۧ�Q�fc5c�5˘t�c�,ĩ}آ�ˊ�R��w�].�PzS�-���i{�9*ҷ:��&`bp<�{˙\��9Xʇw�/�
{ֵѻ���o�����k���V��E�q��{�L��ze�I�+l[�����s��mG��Lv��Vi��㴤��8War��oo(k��Ρ��'Ѹ.���0�9�ˮ�|�l�{�;Z�_3���EȵQ(F���`�s4�^��͎y��s[ךB�,iZؠ����g5��6 ֵ���{�:��V�*1�1,f�ъ0��j���9�1��4Ɲ��*94;={�S��=d�a,*�]i��1�SF��]v��;UU�q4�1&�g=�ˌԃ\%�<�3o
�g��V��,;U�:u�j���4����
�Ƙ�i�k���ܮӮumM�������4[�K5kf:���z7�w�Up�ڛB�jԵ��3֭L�%�rD֭��X�3Z]jM4�u5eG�g�WFg�jՍ�����i3T��Y��yS\��Vl���])(�%�p��5tj�mQҫWC;1�`�Z��:fՊ��8�`WT���շ���(� �M@�:,����:3I���R=)��p4	) ����6�R
e���R�w@Д�Xfe��� �?Z߿UfVk�}��H=����.�)4 Sg�3q��
e�Xk����w��x������i �˰�
H)(B�g�p�&�RA@�����w�s�5�|��A`y����
AH:�fzᴂ�`Re�
H,�d�2�����XVfjH,63(������7��'�5Ix@�A�����G�V�,�¯���i!R��E����.�)4 S̸i�) �fQi�Ů����ּ�5��]R�s(����뚉H��A\�<�k�\4nݥ"�Z/!�Awwa�aI%S}�$���������]��TAH4T32ᴂ�r��{\�u��\�f�� o�Zy����ݚ��n�&��� ��}�m ��
@�Qi4!I��S�w@�RAa��v�R
e�uD) ��>y��s�kz��@R
Aa�r�|�I
���$��9n���Vo���4�[��xaI ��޸i�l���G�Y���R�w�>�޲��~=���ҡ�e�i��3�ZAH,�2S�]�PВ�
��Ci��3(��B�%�2��z������6y���MU�����kw����^�<� ��E�Q
H-w5�
AM�3.H)�3(�Aa��\˰�aI'7���ޮe����k׿�V�p�&�I���M$޻��TAH5P�ˆ����8_ι������5�@�|����R���)��,��/��Nr�F>�G���h�S�鞅�{e���5-ِw9��oa������9����̡;�#.��5��vg�Ò	��X��}��כ�:�X|0��-&��Y)��*���3,8�
B��̢��!I̨�S@�L32�0&���ng�����tMn�=��p�s�/}��� ��0���Q�̸BН�@��{`a�?,�R��a��PLZ�!B�����]m�at�M�1���3%\�&	b�x��$�5E���)�TCBJH,(;ߵ�aH�ZMRAH.�x@}"��n�ER�p�<	��H<;H)k�����o ި������{�I ����i�d����E�aI̠��I%!L32ᤂ�P=˕�����H/ݨ�R�ˆ�ʼ��|gZ_x 
��� ATd��TCBJH,*{��6�_
>@�o��?A��>M��ʧ��ɑ���hJH,>�,6;H)�QiTB�Fe��AM S̸i�d���!�F�R���01����ǳ���(�o�a�����{�$�����A`hi ���
A�C3.H.��3(��$]~��s���o�&>�@�<$��w����)=E��!I ���5?~�5_��+�m������AaW��
B��>��tQ
H.����{����1 ��)��3l��P>��XhaI̠�$��0�ˆ�7I2�H,F��P3��vW߾�U�R��7��i�~����߿}�Ww�����O�YC%?z�ZII�{.H,60��- �M�2�Z~��_7�n����i�+m�����A�A�K7�F��l}ƺ��#0��
�3����u�^]��HR�@���{�c��a�=������������7�8�2�n\gL�:���m��k[c#��Gh𵥊`�����N�l�[�Ԣ�V�ѮΎ8��ΫZ���і�kE;� �*�R�GK���9�an0��ḱ\�s�1��z����[��8�7�<�M�. (�*R�W#f����	�\�*L�N�JR����b�v�U����\
,�2�8��˫+n~�Y�S�E��a��Tep�#��l���:�5+�ԶԖS�{'@������RU�h����RAk�֠)4�L32�m��
e�Xk|�=�k^}~��/���~H-��<
K�m�Y�s��;�\4�R
�v�$�I�.�j���h*�p�Av���-5) ��%9�p4�����v���?k�����ܢ�hB�%2�����jo�����_�~���Ǐ���w$��������!I��H)��fe�L�}G5���3$��P=�- ���Ã
H))
a�e�L�I2�H,4�\˸
A#���^G�?|�}k�0�G\q*L�y�/+��k@������Y�J~��	) ���f����q� fQi �i��]�P4%$�a�v�R�s������/��w�s(���R߻�@R
h@��놙���
!�F�o����������_�����[�� ���{�2m��P=�����G��É �=w�D�AP�޸m ��
@̢�B$��]�P�II�L��6�Xm� fQi5�޾S��:������'�)�]�P5=���~�OW���[���� ��n���
B��=�- ����kP��Xfe�L�%$(C2�$�;�[~�Z�<��}H�F�f�U�(V�1f��WX�w8oTfX�������΁:筺@�w�JC��p�&��H(��X�$2���
Aa��$e~�qo�M���X���q e�Dx<	��8Gw�Ͻw��Io?]�PВ�
�٨m ��
@̢�hB�
As.�(JH,32�c�����3(�����&چ��tE��[P�����.[`�/D�3ta8�n��˜2�f�����8�ʷF+�dzu�]}���R}y
B���{+|��/�{U�;�@R
x@��\4��JH( ��@�<	�U�Y�6���C����,�[�� ����z�M��
�Qi���As.�U��z�������*�\6�]�
@��ZAH)�]�R
Aa���Ci����E��B�%2�˸
�L��y�����A�o�[j�|,�µ���
C�P��tQ
H-w5�
AH,32�q��
�eH,4�v�) ����M��z�`|�~��O���^��$��^���
A��f\6�]��W�u������^��~��
Ag�%?z���%$n���_!��Ì)�(�����C)̻��i) ����H)
�2�H) ���� ��p�9��V�:��ś{�$� ��~�I���>��~ӟ��������[��xaI%A
a���L�I���I����wEQ �C3.H.{�v�����'��0��)h�l���6���wVB3LՉTv�%�����6�#�fm^M~���'�f'�
H,�J{۸
II�g�P�AH(�ZAH,�e9�p��k����s��U�~<~H,+{�󴂐���_}�z����E��
H-s�� ��놙�JH(P�eH) ��a�0���Xfe�L�I���~��������R�I��� �}��u��t�n�I�݅_x ��� AP�O�wCQ%${��6�Xm� fQi/�N]�w��o�`|�Y?��������}�㴂����- �(�$�5�
AMD
a��3pd����E���/}�ȷ��Ws��Ԯ�m�9�j�Wf�1��9V�8s&�U70к��εW��Y��u����sJ:F����0����c?��.������C����,�W.��0����)�{�2lI���$�H.e�UR̸i �`Re�@����|��w�=��q�wp:��
�sP�Aa�=�-&����L�2��5}-g�bw:]|>G�>T��ƈ�RT�E�Q
H-����{�ϝ}� ��)��}p�6��P;��Xi�$2�4
JB�fe�L�e$
3,�A`hi ��p+>��\� Ԩs�H.���Wu�}�>����{��9��H)�d�޻����^�چ�
A@̢�rRAH.e����q�m�^�_��JՎ��jY��k�ᕺ�i�vDu����B����4ѧAI�K������
A@��ZAH)����
AH,;�p�8�I
C2�$��z�k7��ϏWo{ס� �˰�
H)>���կku����y^3>
a�9p�'�RA@���i ���.�~�J33F�ʱ��񏚡
bv�DN��p&�MO�T�t(��AJ� ��@@��y�2o��c+nB�͏/z���[��wn�[c�$�O�����tm�q��!~-� ��CnD�vz����|�^�@�|����$7
��.�Bz:�TЋ�p=ܤ+w�������%�@����!�ȕX�`�OnghV�s&�wkW�=eX�Wk�[��PK��h��r:���M�֙�/r�!Ә��m1�`9�"An<�p �܉-��O��pD�{}�O �\���\(L�	c@6ՐCh_%|:s*T�IF#D��g[ڭ6룦G"�{U����1a��6�]4�� -���|A�Ax��ۑ716��j9�[u�}7e]lB送�{6,��[��Cm	�n �S�*wp�[�m	��95�c�R���8�o/H�@7f3D���y^�6���z�̀�����|�	Sw�1���}2e���qQw������� �VCp��'ү�d��T����p��mȖZ$�c��{L���@{Ʃk��.��^Ǝ� �{�"hO�pǗ�m0��:'���F��=�˚зI甪h+� ���$n�^!�Gŷ5z��=�Ï�UAu��in�ފsl�kԭ�5�/�S��M�@y����Q�o3{�#�d^�w��c6��O:�L�y�������%s2�ܜ%?�PP�ޡ�`qHYp�m�8��S�:�c�n�&�.�����*]�^��4Y`](��E���m�Kc*��1�C5�^,�q��ґmQ��\���HB��Hv)�m���4YD�̄�$0��uAم�iv嶅˨�[�&��JP�����VГ&�;$��6+mi6��*�`MR��u{V��fSHMy`IM�[W�%�L�WL��ʃ�������̴�����FR+c-�S�sS[�y�#�@t�Kl��[�יϨ�����O{V"=p&�MO'+0���&%����)�A�^@�5$�@����RC���A��r�kJ˧B����o����&���ц'n��'��|�g8h�n���=���d׵Os��;7�����౓��4�8���PGͥ�r$��En$��3C�1D��>� ��&��=I�3���1= �{�9VL�S��uǫ�h#z�>n<�V-�����8EOo�3ĥ��p�n.O՚�`9�
����Ȑ[� ��<Ug=]�}yg�X�6V��W6�V�0�kDٲ��l�U��Yi��& 3A�P�[ ���6��!���H�s\6vv��]@z�L�lf��py��H>�A����۟7�ٱ[%��A�����	ý�V���5;����V[�����
B�H�;���;�6�UjDs҆v�Lkyxw 'q�3������п��#���g�M1�"����� ���n [j���T�H���/����z|��Q�ۑ�e�[T�>'��o/A|�`9���@����� A�-��!��;6o�Y:^@�r�m��t���#;X���(w�y��fBF^q��J�V����"|[�A-�@�r$�
��:O]��X�4��+8XR��t�Cq���R 6�!�rX����i[�@c�J��8Cv`حԺV�썖�EK�XJ"LI�Q�q���ԑ� 7 Un�VR-n�j�3��'5��@�%��H�s�8y�H�� ��"s ��/z"�J�m�/�^��/s<��v��������N�)n��!��Q:sLy�f��qc�ٰ ��H-����6A����$czd̲���"�پ�3ّYg����aG}���6w/L��]�H�
\fCv2�;jI�Z�U����xx�xr::�h�Y��A����mz|����VZ�u��u�`��h"3a�r(٘)k�̅Lqȗs�������m҉�i˄}� 6��	n ���mmez	pbS��u�O��h�-������C���Aۨ����>�3p4l����~�S%�Fe#j�nj]��,�k��bU�0�!�i�A2��Bbg��gDw�� "/�y��	n�=eZ=�kȼ�aD�ںn8魟S�UU�ӫ�� [A�"	m� ��ǎ'5��n�nl���PWN=̉�r%��Aހ�"�dIn/]٫�]b#�w`t��̴'��@͠j� 6�%�ɜ)KT����{�P������n�^!�<r$���DU.��j�z`P �_d�=��%�M��f�ז����x��Dg2HӍi��j��,����9=���9J��V��b�	�ȫ�:{"�{\Qc6���oM���r<ȁv�5��MgVáw��fk>���xW/|���7P^!�D�^�6�n(�N���5z���>��PW�}��7��2�c���@���|�Y�k.6����ˀ�L	F�Pcn�a���b\�S��X�Am�Gmfr�5�&�Bɟ)7= ��;cȶԂh)��.}W�&�����7�1ZbB�����~ � 3����r$�A�r縆h��i���'��ѝ
��m�wk8XQ= ��5�[j��H�M��hq@�kRn �|�A'�1�N��'4dw�בV��˹� �� ^|�H-�� ۹ήCI�WyL�-�#�Ԃm;y��j�D��Y�6&��o/u������]@�"|[�A-�^ ��������=TD�`�dh��jL��'���v������}�� mH �Ѐ"w&��j�N��'��i82�P)a�5�g��;�������rM�w/&��/� �^N��c�x��zo ��^,�yop1�`\\ٟn,֛�o��۷r-Z̉�ŸN�\W;�ٮ�U�
�$m]@�U��h��&L�,:\�M�ٽ���ɻN���\-V,��lI�,�Am�"�U����R(V����n�Y�"\�p������9R�.���(Q��YӰ�ۅ�.>�ல�2�����`=}���5.֡��:8�����������"�'h�$P*ط���{e��ŀ��XУ[SR�*���*'J�v�-�9#+R���ã�^m�,�;G��v8ʥPVl'N��U�"ëbl�ͫn�k綮껱}�Ґ��i�D�'�H�Z����F��}u�2JЪ_
�	�6!)��3v]��e��{s9}�S[��O\�f\̌j]�Ä'X�x���ڧ}��g9J���o}"`��Xy>��#o-V����A�w�N���F����ej�.�d�X����;�#y��\H��A
�����([8k�^V<J��*��a��O�^fu!T]��s!ƨ8��k.veӳZ,�O+e�{;��;��x�n�J� jWZVQ��]���.��w1�}��bN+�2mwݦ��&i' �n�ޮ\0n��#�ب:c�D��t���]W*oeoe�9d���*��źN����N�&��~���J�!3efr�,i�ԓٖƾceJ��x��	�n����4�d؛G+ �|0�@5n�K4Z�����N�+A��Z��Ϊ�SC�l-M��V�F���N9��?��Zc3H3Z��Y�<��[�-J�=n�3���G1�,��y�M&�Yik��V������,�id�4�f¶:�^u浘��+w�oVk8����]�CWbj��ގWI�V��8m���i[އ+Y��oW��C4�̨��T�co]uul֬���*ҥtu��l�f+�5hfӭQ���1:��k5Nz�zN��Ƣف�vb�3*�iQ�N�^oOz���j�Y2Խi�j��2��gV�m*���؝�r\q�0޷�+���o{5Y��k�,Ku��Tl�9��t�k4�sW]�I&�Y��vzZ9�,���ɵ�+�׮�Q���;�����5ܭ7U�5�i���{3�1�o<��ui��)/�@8��׿=O�,\ы��)�&K�thR���$QH��[(@�hGb��˫,� m�^�F�piVR���Yn/:il�ڮ.��f���
]+`Y��3E�Ԍs����6Ԧv�$nL�Mn�*1V�;l����Ў�B�]�K���a�;��@N����4�1B.qe�lҭ�R٢��1]3b��y1��e��SCL�,��Ke�e�Ҍ�Ps)N��AٗmS�6HJ���,�Y�Sv�Bݰ[]�%X�i�Y�F̅�F��Z�.�蛇$��g&�e�R��V�w5�[R�u��[�&�֤����u�ņr˩0^�ܻg̳m)���p��\a��bX�@i��m
�Ж�����0�6�R̃wb��.�ل����a��2�Kv�^��ځA,�7��6 �\���;3L�46q�3���73l�f��a��Z0�L�'5[a4�.�EЭ��T2WS���.%viHk�uڎ��R[��*��0�8:�BV��jv�*��.rWMs�x�ַd�״�BQ�Mm�6�c���3.o6:�Fm@˯l��d]J؎�"c��`K�44����z������D����#Rҷ`�+L�kkl��� f�-�q���D�����]l,��>!-�R��&sr�Q�`�Z�H��E��JY�W�N���]�/M�[+�)	d�!H�Ju�c�ۥcH��������n�̱���6���se],��T�ؒlb�{IY�ʺ�h�ݵJ��b��
ŕN�F>x�Fy����d��� ���lU��_5�<��%��$�fH�����s&ڪ��2����9����+�xch�MAn��H��\b�rk5�sDv��
�I�.]+�62��c��Q��)WCM�����ƍc��U�p�4�pѭ�ݕ����l8��2^ݣ%pv����JUM�2����u����K�m2�Xҍ��-�q�BÊ͘��R\Eɛ4�lj]�^s�ڰhlTC&�6����*��b�2�6�`+ke%X�B1�������I�Ќ]M	t#�uE)Hm��7�]�U�'�vB��v�Mt3]7�xy<�DZݘѤ��1��"�QPIf�En�05$�kV�ް��s��[�% hG&�4� -$��"i�(б���QA�M)�+�� ToZ)��V\Xcdit�r�����Rb��Auγ0Z���&l�kA΃��ʎ}���JD:�.n�tʘ�l�ƅ1I��!Q�0��m�Y����!��Ͽ� Cp���l�ջ�V��%��#�#U[5r;�T���l"�p!�3��/0�g�9��Fy�k1O��N�";6�tM\��Sbn;�^�C���wb�m��Vo����H8�xG�:|�nD��A�-�����t����hZ��,���
�8� ��-� ��#��734��VFl}�/6П\Y�+ow.2�}�%�����(wGc����k|�i���Cnd8�nx��.�����FU����^蚹�2��7�^��$�>m�ې��s�EQA�P��b.T���^9�+Ne&u^e 55,DnB��a�]����[��1���A���qdp�5�XY�����8XQ\�oG�5�[E�p �/ u�A�h"�A �jO��W�5˽��!~��w���yy��H�x��e�ع���z�itT��r��P<\��)l�r�Rw[;QM'�{�7�V���>�	��pW[ܸ���}E�����dH-ŅX�oz�Z8��S�-�	��mI͠��@ٵ��Dg]�h���)M�����RA�"����p�F�#�fN@��3��܉z�〽4g��Y���.�8X*�H ��^"��`�I6��mR���R�/� A�����D7wr3j�j�d�y���>�d�}�rk4a�7��y�^ �ݟ7%��99Ҷk/��Fb:D�����h��K�E�Jܚ��C1���l��;���)J��^�?5!�;����m's��tM��0���w������%�/�◸�t �A��AnkU+̲�d����@A݀���9<͊�/�����{`"�W�-�/� �ٝ�)r�NB �suI��r0��e�뫊
G2�;2�_e�Ņ�l$�v#�U�a�Q�����N�q��k�?{	�F<zycƴ�7�'T=g�2�L4d-o.���x{��u�U�m%���V�� A�nȒ� A-�����Te�鬣��q���٪A�'�ͻn��WBn8�{�|C�8�ѹ��F�M�����2��!�*I��^�]�̖'�p+��lX��Ί�/����lA�j���!�,���J��D�w�B_�Ԡ�����	Pmh�ҵW0!��M���UICH�՚��.g+���^�a�Y`��#��ۑ"�]���b*s7�a�q��=���F��kc Qz�I�A-�D6�A����R�(t��9���Azv�@�[{�0��ºq�^��P^7������	��w��6�7[r$�An�����wd9B���7,1�N__	���mO�>��>���f�y0F�΅���p.�]{�Js7݆mǻǜN�ޣ��y���ظ��xxOx=&��]�媝i�}���'a������D��jn�˸f�\4G�����q\#Ee�J�A��lPg��<=�!7����� mߤ[�k���ȳg~ܦ2�
}��V�iT�(���8��)�Z�7�ŷ#0泐�q|��`ZD3]Q�c�JhY��0�f��p�pa8�k5�%�eH�&7� ��@D�"Kp� �U	�rrx1�j��
�+9]��ڡ��`�ؼ��Ԑ|���-����E9}5���n4'��׻��Ft8���x�>��p$Ga(D���D^�w`"kȶԐ[C�f�u�wi;f�52��yy��ZUl����sPD7���"|[�Ge�D���LR�+Z�q�[�����9�Xô�gZ�������v���jA��Amz@m�s	X3.{1�����P�`^��W�uO9������۲$�/q�늚Q8
Iʁ�ө:;{{��	��6�pNݩ<�*a6����{)�<@YӢ����ɵ�yrD�M󝳍<{C
��8t�$�{�>YZ��1f��+�am�W�R�062���j;k��a��X�ͦXGF0�Uem�Y�jv��Xc���li��ex"�eH����3��Al�h�Ff�Ըv�θc�X��	��nk0ʃ6����@�;c.�D��7َ�0�أB� -�[SW �ܔ��k�KW�ۑ�ֲ�r��Qdk�� u�u)i��1���,�fa���������It������R1.es"��"�L�nS,5��m��%�2�?c��P�A�����
z� t�{�3آ��Y�b��]���xnח�nD��H��׸tn<]u�q��6�W��N�k8X*�H ��D[�6�Q�3�t�8������ ��/6��m��pt�TE�k�XB�T�ȥ7�3a��G�΄#�dIn>e�6�G�和V�`�s0"�>j�!���@\�wj&g�E�3��)"�nո7��b�mz<FvȐ[��	n�6�In$����sjȑ��G���Xާӵ�,} ���^@�Ԑ�	ƻ�����Ø�}K�F�@8˞K�T5�(Dղf:�W+�Ms��Yvj��RD(0a�A�j|A�@7|�B}P.�]zv�޳}'*8WY�z+{�ɪ��9 `u�$�D� ۹�]
���l�/d�R�������	�`�nA�n7�f�^V�X�I��"���(�O�5w�W��X\n����3/{j�\r�WS�:���;���o���;�O\d���B�옻�s%�)�Z��-������*�&�� ����"|[�"�	��5{��%)��}w��U�}�[^E��[A� B��7�� _8�j�=�";`r&�]����)��8���	΀-J���q�� � ۹Ÿ����&E�w�w#{��������7r.c�A�) �A�#�۟<��ul�vm̡`ꘔ�Ģ��k��+z�K)
�GL@�����N�c6�o���N�����ϛ��T6�XΧ�6�3���n�<�q��� �܀��`���/Am��!�vQ�+֠���nȢ.�[Zv�m�|�M�{�tA��[���P��*^Ɯi�@�����א-� ��M�ܦfw����̱'r�1-��j´Է>i^6rӥ�oa�}ܱT��=��+;�5\Ո���Ǽv���Lͼ�����gIN�
���  `Քc/7bT��qr"��|���}�Cp��mȐ[�F^�X}9�� �Α>;Ј>-�^�3�E,5�s����8��=��ݛa���k�{�� ��RAm��*�i�h.̫�k�c,2/_M.�~�8���G۫�Ǭ�p���4�� �"c<�+�Cv�;�-эɩfD�3
Y��s�eB�HR���{j ���[jA��7� �hݘ��w"�q�<*�v�s�ҽ��/5�>>mȒ�#��C.Y;3x,�B ���UZb��n�V�9��H �c@6�i& e[�B��#r�'3T�h"1�>-��,neds΂x�����hu���Gx�퀁�	-Ǒn6���Z~��SXw�b�n��oT��AN��;tn�L�;��%�)"s'X�����l؛��G:�wt���fG�헬�M�Yu�����}w��--cC!#.�0-�|{r�R[t���Qy̞f�~��I&�Ý�1>��5��g{E�{�5��
��m_�.5t��U�z���3Ԫ���p�/�[A��Rv�;�e���챉��鈸SiE\6���l��m+��v�c�3e~^{f�� ��A�/���l�u������m#�Bk=���y�z��aw9y��m���/��PSS[q3}qS�Or���D��<ͯE�����|�x:t�59�%L�n,|Fl A��p�n�w����s���޲wR0j	�1]� �� p�mz|^�Cf���[�uY��P^m�7jy������ᴏ�W���x8��B	��� ��Cm	�n @��;����e>8�PB���;�%L�^��	{�H:׃t�n}� J1\���_F��6;s7��'�G$I�+��m��EEJu��Uі(iP�.��Z1(�*�jA����m�oJ�/u���H����Xi�h\��@��u[4T���qui��I�cq-��[{6�tYe2�h��+
؉[�u�\��J��5�[rX��]�+����&�"Rs"4��]XS	��;�����j�L�:�����ڔb��W�VW ��C=��Z@:�ZGm���m��Q4B		k\K����7R�ֵ�Y�
l��j�k,�ge�z�lЋ��K�w�����O��ZJ�k���[؉f�(�6�l]H2����e�TZic�H����z�q>}hH-��*�1H_�c:**�P��Ed�n�Ɉ���S�h |�ڒfEQθ���v��^!�f���WR�v�J�=���D�H��p<Pes�8"컚h�Q�Q�t)�����A-�@ڒ�{#/I�}�=�J��bgp��_y�RAւͥ�ϛ��Z��V؞2"#ט���d�*����s1�J*�H�]�ǜBzє�Å�����k!��� Kmz[A6d��C�wpZO�eȗ�(܍���ڭ*�����}>n,���p�U����qI� �f.`��iZٳ
dIn,շ6���i�L��� Х
b�P�O��  �@@�כ�b���ə�2��+����1��V/��|۟7$7t^�������{^�|�K�Y5p�c�l��G��om��놦�@3,�d��u'��2����G<b�������@Σݱ6NS�����_�	$5�h��V�}Vo~j����f3�E_	�� G6�ɘ��Z��^��9��Ch |�^m�*�E�͘IS��Gl���wU�U �\�D��  ���Ȩ��il��	܀�wZ��	��K�9F�:3<̯E��{�H"�c�7V�G)���E��7�	�ۑ ����uRĀF8S�bۍs1�J.�H3]>�x���mH �З9��n5Ͽ}{��z����nB�5\����v�I]���*�#�7�Z����_]����ߎ�Y>�c�͠�@mȳf�GT�٤��ܥUzc�=���� �=A�H��@�Cq��p"�h�HV�9��f�#\龌K�.�h�3<̡��	��$k�c.�L��>c�H��^ �ŖP!����@��h�x"��\Q����;����4#l�ʇ=�/ b�X��p_7K7���v�l]�sN������p�m�n �}]7�bi��ï3.`]՗y�l�xoU�p�-3.g9�Vh�7\�֨�V��-[;p�ޮ�xXƯ%N�㔰���M*���&N���'��D֫�93jP��I���.�T��+�Yx��J���ujT��c��yM�/IM	v%P��
�X�U�Wl���f+똖�N��2�+�ˬU�6JIK��^=�d�"��pէ�72c�x���� �8У �Oa[E��v�L��vv.�������I0ٜ%7�aOy_*�+8�coܮu�Z�|�yo\��>�Μq�'����p��b�[{�b8��ٺ�a��$ʊ�m±Z�6��vs,�����'|�KU�������[�[��I�M{H�]8�7=ٞ���Ⲍ�t=���c�V��[�'o:�3���
=`�G�<uv�7E�f-5>��d�^�wۗt�x�`���]�a����v�Y:��؏	@Dr�Q�N����}��[y`2�<0rGk+3d�3P-�����)Mbк����#q��$�oVk�`�d\���u�-�,�º���kw��x��%��M\B>�k0�P�u�wY�΢h��'lT��UL̥;;{6cm��;�7Df ��̼��{4D�TsEMJ���u�7Vs��a0w\�F�N��vL��7�w,nn�|�N����}C�$.���:�*RС�1W3�E�yDbj�Ml�C�k��7�����?^�W�s��yU�JJVU%E��i�S�K&V�sd��e�fv�e����;5lbl��5u]Q�s�a�d�d�1:�w��g3����*�iU
�&)0m���8�b��Ù��E�ͫX1ڵ6�lKQ�uk9���i�յ;]�{��5�զ��K�Ӏ�{ךʎN��V�������eE-K��8is�fe@3VT�c��{�L͙�*c��8�wbq�U���cZ�U��J[
�@gf0�t�c�L�9�`�V�Z�ff+��Z��ɪ��ʜuN͌hY��l�˱�Նm4��Vј6Lu�9��W�3g��1�h�h��gf+�umc6Rʮ��h�������[W-�bj�;כ�uF1E�\�889�Wk6g9��s18ܭZ�6�g8�cgMz��{��N���6����xxj��g�ʍ�J5�O8�8d [jA��� e�U��1*���G��"͚�yY޼���<�H�p��X���'�ہb�t��K����m̂n!�B-���s[�Yӂ�A��ӕX��g�� �z/yH �Ag�6�GEgX�GƓ���|����a ��vչ��q�F\k�1��n�-,��^"��vq)�Vm��-�}���� ��"Kp�YUZ""�g8QՖ��@�] �_B�|���;B8�I6�!�B-��ݎC��sA���F�x��"͕j���13�1Q�:x����qu��RD&c�{~�|w`/An ����
��1Y��1�P���t)��������ͥ�r$�!ZP����h1G^!><�A�W�G��Oa����Oa��GL�;ؽ��Og�9��N�V�8�uYn�+"���4��������Չ�&��1��"�P���z7p�T�0鄴d̴G{��������b�|�ͤ	m�Kh/6n�!�f�r꽠%R$lY���:��ETp�z� 7�$�A��u���=+E|�������|�-�t�0]��ױ4������&�xnY���nց��,��s����X3;E�[jH!�/n3��',��	^��3GK6\҉�����TA���m�fG����榶"3ձ��6��E#���j�@T����c��[k�"�ؚ�>�A{u�Kk����mz#n[�y��9*�#jt)ݘ���wB�D��!��n�*�;�};.�@~z��گ�н��FP�����	^��^{�A
�"J��)s9#����r$�	�!���r1���]+��8��]�R��ҕ���.����>xׯ͡��.����]�6�SʽK^��A=�la�c{��r��C'�����&d��9(6��X6�����	<�[�U>Hv_ﾯ�������X�����ݠ�
̀X��P�&�i.����d�å��s�e�\Ui�����H�
��m�gSh�!)��	l�˒�fi�e6 ZD�ibR�bm��:1�۶4�ƪ�5��-�9c�L:�X$���;Gi��a'v�e�	�b�e����٬9�WB��n"U��Q�KF�����&�]Q�`3��.n�43.�O�>O��i���R�ma6�L�f�E��(��/h��fl������������!�������6�ME�Qҳb6����11�E��aa�͈<܉<�-�@���%� �5�f3FDnM8�����k��r3��%�Z�9�P�����kA��D���g��	�ۄ': m�7����!��-��y��EG\51���R��#6 m�_�Ax��5�Of��U���4Ё��nD�T:�.q<���u��~���X��>�v2�^��w@뀈m� �Ck���L�X�d4��hę��)�9�P�A ��> �A�/܎�N��g���d%��LhP`)��-���J�XEx��:�,��qA�F����m�B���C���H-ǑnWъu\Q\$N�ۈ3=��"� �U���ڟ zu@$vL�vQ��j�n��"�THz/ v�ާW������պ4`��t��g$�n�����T�BY�����&��������G���G��oH�U�j>��;��}�"f8w@D>�[��x��wpAn�!�H �Ck�ڐA�3�<�,��ll�6�_	z%Q�_r��@7�nD���<��ZH�n`2b��9�*��ODY�Uft ����^"�J�^�9�H>mn ��I͠�nGN`�;v���1�f��Kv"+�D)� ��@@�{"Kp�Ÿ	v�����/�����f��.���R�t�[�˛�#�`��B�`���	��,�}}#gߧ7�ό��A_^.	L��$M�-G;^��y=J�� f��ۑ ��p�C���gJ��>�y�Zb+�s��\WYAR��df�"�V�H���m�[G��DVB �=RCp!�G�6��"ȲXm>��θ�
�;B�/\Y٥�v�1E`y�63-̵mԜF���lan�9&״l	��Wuq#[�������=�Gi7*�an�ڢ���[�[�A����E
�fR�A�@v���0/o����D�	B�p ���A�����M�)r�����{>n=`�r'Ÿ�=�Ap(����2��"�8��(L��v@Df� ^5$n�ĳ������S1 ��g�3.�Vgh�2�Ă�0s	��T*ٶ��kS�a��~K��	�k����>!�"EZ&�&�9�U���1�8��;�H�3$�72D���[��!�>�|[�
�޼��4��� =��[AO^t�!2��7�P��G��I����[�7����D�ȓ� wB ��O�p� 7Q:�m�f�Yw�gg�Ю�%sC3�B�����ڒ�A��T��u��iiP ��>z��mȻ�5�u9+`��Q���?���_4�y,�U�[(hxV;,�[em��LYh��YVoTjմ�n�UE�^�ó��U7;S�����3�VR]���1�v*o��神��<�*� �z�������ǽ���Wk�5S�AԂ�y��H�y�FH��Kָ Ow) �h"j<@m�v4��_^�����Դ	�n��Y�kfB).Лl�m�D� �^b)�,��5�[�����޽|���,��V��z#���.��S�@��D\8N�@����dW�mIQG�i�;8�>�,���nDݨ7�u.QЯ�D)� �(�P�[�W��;'c@(�@�ޟH>9� �d"�RA�hfu�YN�`�4W'1%�prr&�R��'���� n(������Ԩ.s��sX&M@nH��G��B�LR=����Q@�C�쀁m�U}���ŀ����-��mnz�5��5�{6�D�q��R�
�TB���  3vD�� >-��첪`)T�-�rŤ�ISD�V��ek����Κ�Ź�oj�V��x�uΆu��c0c�W	t�yM�26q�}� =���TaPH�1((P���-���k�S��J�eʹ����2��V�K27^q��-�h�!��tmFf٩-�p5ƗL%	�\��3W.� ���m]2�s�lau`�/k� �A��mj�h��\��QD�K1H�%�2��M����r2���2FZ�[0'�ҫvB�SF2� 2(�R���Ż[fØgf�k˦f����3(e={�����T@�7].n���2(f=��]k1(\A���9) h`��7�	ۀ�#5 �W������F]g�"o�!j8���LoZ���k��mȟ�An"��kc�r�j���[����#щ˞�Q�P���H ��3W��mv�����i�KJA]N=R6�!�@��܊zN����q��T��o�b�Ot��$�x�[�v�j�{f�^@�G\y�RA�hOg9)���J��"�8N�)-7�Bo��Fp���"�2'��7:D�� A-�7�Y�� �GG���bE��>5c�U���֧�i �!��@D3��m��Mx�^�e�;C#~<�$��E�e
�4ZYX������Չ6Xm�[c�5�����7����n��k�fv��R[*/�1���^��U�O'{�#1� �����p�7��J�i yf��_@C�
]u�:/�^��;�J.�m�\��f��L�WڪΫ?>t:��3!9Ι��)H��^0�\cH������u�9ؤ�>����%9���z2U�� ���Ak@7#��:�s���H�s�|_@@�r$�@-��
9·�R,�Z皞�������@D3��d7� E��D�*���A^��#6��n}vbcv��6T_m�)�>Bw;�Y��mв����D6�A-�	�md��N��}�I]?o_Q�}Oi��e2x��S�A�ւ!�G�6�k����ĥ�U_i���#f�`��B�P�GHl�Cb-�ue����Ժ��c�k(��ӛ�ݾ�q��A�r$�@-�^��������� �{�I ½B{�X#� ����� Cp� ����lN���`��G׽u��Q�Y5�e��7���X��u>-�W��x�y3��6�m�[hbj#�.���D��1D��gj����7+�Oa��<a�5����5��V�پ�o	�]E�K�ئRŎٸ:ѹ��pl�< �eF�6j��_z���� �r�A�Ax��x6�In8m�laΉ˱� _Z��p ��/Uq��'!;�=)�A=�"�������l��[^��C-@ �Ԑ� ˙!1y����m9�*�㨎��6�*�p<x�svD���Y޾~��{޽z���fua,��f�nE����u
ј��d�t���Ħ�ۦ]Mٶ,/���@�t�[k���Ǜ%�N_�U\�B�w�th�ޙu�0C��ij<[r$�	e��4��--���\#�t��1�c���BfPQ+۰8��� [j��������!b5 �P�^�AmC-!�#*�ʹ���tD
%7S�QONm�+� �<Q����Ȳϛw!��:^LA�㙪A6��<�q�|3}5s�1�@ �r�\����&��<owG��袗�aÖ72�#{��@���]ۙ{�.���N�L:|Ø��	s�����;���ʲڈ[w��Kk(d�?���y+�|3zD���� Amϛ���\�,�5�����{LDmg��u!3((�	{5yڒ�]6����ۀãDej�� f\�JւC7J������k35,��sV�U��s;z3,��j�'[� ظ��YN��4�ݥq�Hqb\Ȝ�FW@��D�_B��D6В��D�+ojRQF�+=��g9IݨO�2"��d+���=�{��s�@��m}����ND��D��۟7��
����T`�Y,��[HL�
'��@�^@�ԐCh"�Yh]��ي*����ւq�-�l\R�wP��ܻ�W i��G-���ǣ�-��.�(�ϧ��@��|�SG�glm�:� �zy�q�z5���1�/yzs���y����׺%ݯ	q�[[���NX��񱵕�楷p�Ak皩����p�_d�
�˥	H��Đ�CU�j+�GjZBV]�[��n'R��"t�u:�����S=��^R���͋u�,"*�����
�S-cJ&���%��c,��z[뤜�q�+�,R��,��X隓h�6`.��xޖ*�T9�e��j�oKS��a��Kxv�u��|��sM�*f�����H���P�(nsP��5Q�y���ZS�]��.��*�F��T[U�����5�9���*Vs����5��j�U/�U|tL	��-|���^��:��6��pUG;�Z���Ӯ6w65	���1DV=d��'�+��W�K6�C�-�Ќ����N9��p۩�J֦��YT�t28[&#D�;[�i��,1R�,���>����E�����<Y4#��ӽteu�Q�n�k~�r�����w�Sc�;�����<�J��y';YN��J�c@X���V*6�kӊZ�m��ՙ0�Z���yw�.��U�g^��n�] F��`N��%.�p��&��,�3���:�-琳0ݥ��uc�W�++�K����Ɨ��ptU��M���14�x��o2���M"@scl���a�Yw�Դ�ޭ&*f��TFH[[�����b ʳ\�o�1� �-�3�ڲ���X�W�U��+��_1+'+�-)�z���Џuv�Ùp�9{�0�PUy�%���E�D�6ܔ��G;�3I��0���Oo��6a=�_HC�*p���uB��q���Tb�8�j�ͽ�x���g6�vWUƲLs�ew������Z�b^�s��=iZc�1�l���9���g3�l�q�� g4�:88y��3pc�3����0�ك���ij�3oS�����73�e�q�5t�M����68<�����֌�k4�d���{1������ئ��1��q��3�3c3�Xpylcr�rr���g�����8U�9�����5\+�p�{�8�3�~cֱ�{�=���]Z�w��9�w���A������#'L����,�"�c1͆lwy��}��8�Yڭ�%ڬs �bL3ei�9.8�q�U���0��0��æ��9�ce-c����2L�33��˵�My���i|� �m0i�k���WN�����9�|�ڴUk���*�k��4鵩`��Kq����|��,ΰ1��L=��]tE׳(�l�Bkb1�P%#2�a
m62�pgD�����i^�<�I\ ݈�K��T�6�nT�t�.ev��s����P�3 ���Y��i0��vܛl��ݘ(c4�Y�4
�+�Hg*5�5� ��i�޳���b �B][B���i�B�fjk�e���g�ˤ���.
���5�Y��)`m6�3ڮ�ˇl/.�d����P��]����GW�G:oR�[wXE��ceLe-j(:J[n�=lV�GrdZ� �.#�����e��e�����[&ˠdB�p�ً��]B[�6k�aR9�Zݗr'i�����)K-�\���]���w"�%��-M7E�Љv��S�X0Q�P���e ���]Ě�9k�IF��ldQ�]����-%f�M��bh�b�uð"�oj \恒��.���ݞi1rٱ.s�]�55�X˭%�HZ�ڍ��k�34t�)p������r�6�!��,"b7Z�F��	3ʌ�
�J���`����ʉc`��R�լ����l����%���L�%��m�u@.-mL�ZJ�imɚJ�Z.s����u�EΦ�@n�X�Q��6���KE)p�p���Ul�Fj�k40�&"��l�&��M-�R�H���1���Е�Kv����H�&Ɗ-5��L@�Z.�2�EdN���5���4��t[Z����3a3�P�KtB��u\��L��ո�l^Xf��1R���2]�\�2����5��+�ơR�i�k��T��mX�jD�mm�.��]�[qd¹f�,�JCV�����|�f�v9�MB�!,+k�-b+�Q�eش�W�a��*GKb풛m�fJR��͹p1l��k2[Ha�]tn4dMW,4@�.uq��:ح�Κ��"�e�b*,���TjP���s�n����0lXu�b&�������F8�-�����y��o4�f`�Tq:t��\_ ���38]CI��RVB��뱂�e8�fW����f�E���ñ�K`�*���q���4�&m�3Rf��&���\�g�U)`\k��]a&��¹^���ҀRݹF�m!�|��_�e��66�:\�V��,C�U⮫y�k6�
�ti�fX�A�mxe�m���V��.�LfQ�r��R��3��[�����~�k{U�U�#N�t)VĶ���ذ�y��k�F:�pͲ7�}����}�"Kp�%�P��:����]HL�+�	[�S�:�o�=B7���Ah@%����*v-D�m�4��͑ ظ��M�B��n��n=�<x�A��n��um��ڭ�qVU�L��#7g��l �p�E�S�hc#��\ا�odr��x[!]�`��)#: �Z�6В�z�|����f����:,	e�U�u���[]J��3��t�dt[x�x���{�A5e�Ŷ����@�_>d�A��|���xtZΦ�qup���n8O+�ݑ%�D�9S[(�Rx����D�H6(�M#u��a�D2b0������-��� �@���6���p!�!�^n��2R]^�S�Q��vY[�����y��yG�nD��x��P#��<�T�}N�(#��fr)�3�K��q�D�X�����x��w/Ֆ+6�-��B�3�*�c�9�ڗ*�gr�<�p��$ �������;��">�nۮ�FfS�A=����-��*���j��\45@@&���[@2�<CnD��uG�E��	��w:�S��VM�x��k�,�yY@���w']Ś�*����� o��О9��*�Fs�5s����� �z4�e���FQ�9[�>,��r$��qN4�un	��1�����Tf`=>#H@�ԐCheԫ�WeS�2o�z4��H� �	���]�q�t���-���Ykh�YJ�[c�5���v���R/�!��-��qi�V<��xSUY7EE�ټ`�<}�P���Cmy�Eq��w{�T�),�v����`ȋ����}F=q�@���H9� |�\��ͯ!������r$� A�!��Q{[3�b7�z����L�Ja�����P��Hȶ7fN� �ҙsR�l�{�T�r󤘸�Ej�_[�d��\/�b@��b�V��/��������s�]SFfS��� /��Ԑ[A��C%��ݕ����gia¹��/܉�ŨO�⎞�j��G|Gt"*�:d	�qQ}8�� ��6�A-�^��͵�GQ̫���cc�OOhȋ��o��}F=q�{�zq���q�n}���=�������}Tke�*Ssbl�U��6�i��f���aɭ��J�kNo��}�~z��|9[� Cp����b1���uAL��#vq���V�@��to��m��6ՑL�[;{j�g��V�<�/�>�0*��+��ں٨���k�/Ÿ�{��v�Z�Q�5E/�} ���n-�$7E��]N����8��u�kt7�c� �r�A�4>m�r$�cs�&��8q�5�/aHn&�DtTq���PS �� ���V0S{^��=�-W=9�.�-I�wJm���J~��&�V��l��ئv�(���5Y2\��)'q��dj���o]�!!�]�s�>��w�X�Ƥ��#��%��_���$O���f7f6g�����Gtyn��q�!��Q�[F�k�B�9f�"��c�r�4��u1Q��7[��.nԱ+�]QlpM��gι��v8ڟ�|s=qu�i�4o�Ǯ9��X _������~�6�In ��/��lf��=gg�#|A!�*�eG8z��h)�1=>�9�m�bb�&�&V	(/n�	�� �� ��&܇΢�B�M�VEª�f�{5�Gt Z�q`Hn6�C�:s �u&�x����T�Ch!zs=�u�i�4o�Ǯ q{��q��WVrs�
>�^^;�D�q�Cp�6����o	����`�����nwU�
`LOH �9��ڲ�����:�.Wb_Vm�f���w6(a$S���G'���Vڤ�u��B`��r���7k��W�t�b�#ecޡ�˞3�����ꈿ���޾�=˴b;�r�T��������񩰋p�T��3X�n��H4�欱�aZ�5�R�q�k��ٹ�vu�C!�P��M�j��ʹt.xR�*ݲ�+ ʹ]֬�,.�a���Pf�m (%�4ФVdm�lܼ1�\��t@�:�c�`B�����`<[��]�9^/\BV�Z���k6Y�^�J\�Yp壚(��'���A��V�m2���u��"�]@у6,cj�!"�D��1궽�� ��^^�П��K3'����@q�#�HK�S��r�FTh �\�9��A!��m���Q5�zˈ���j�A�P��TT��M�1���A�@������B��`W��qd�A�"Kq����`�A��$V��c�e�fB ��9��ϳ1`#2<2}�d8�{������?*�ܬ��d�2v�}y�]��� ��z����t��p ����KpŸڮS0$�Cr1��ʺ�7����� �w��[A6���hoT誃2]ٺ�DA�b`�l9�#h	�)60P�jR�tƐ�r�J���5��ՐF'ݫ�v�A�j�0N���*�66qfwa�s ��[
�/a�|5� �Tq�Am|�[jA�����=0�\n�ݲnV��t%Ё��G�'f��.���Ǘ9�ٛ��Y�fmJ[��]������m���v�VJW6L?����7���C�>�b�Ns�)�U���Gt"ײ$�ة趴�Yp��"A6 �� [k��SqDr�5��B����Y��1�c� ������/6��ő�]���/��s��|CqU�#��NFgOa���� ��!N�p��؇�w�=�m��pq���*���T�֑{+���U�b�w���7m�m���ݮ�[MΙ�%�$(�]��Zغ\	3-��q
�%���[��s�yq/y}}�|�s�4���U��7�&u�໥+}�3���-�׃m7 6�ҋ��꜉褬M@څW���rt�
B���3Pm�k#f�������nmx6��CkO.�Al�5�9Pj�$__�(�w�y!5-���s��-�0���Ԩܺ*M��e���Bs�3s5[�e��3��p,Śu�f+�2�|;�<��cm�#
{WV�\��]�u�7;iQI������7y�	��x1����y��m�cr��Gf,�%_l�����2�6���"g���i��h���N�9��3&�I���R��*��C6h����)H�+����;-is����;�Z|۠�B�Y�6똓.y�6\*��J�آ��z�6�w��2�d@[g2�z��g�*P�پrDWQ���5�\*ɤk'/8��Yp3u6�n<ۛ��3���Y� �����*�f{�i��^�m �6�kcE�	22�w@�h�b�Qy\�1˞D��w���;���U�Sz���cT��bb8n�i��@�aM��Q�5׻-ecn�+�tֻa���ј�'1͸����B�ݩ��������3m�aV�r d�ҸI�=�%�6Wxn�n���龮�&�[h�(�Dz$A�ij�4.9u�pҋ��V�[3�c�p�*%��o��y��I��nm	����8�s}��
{�N�4����YC�:����n�m�n�����H�Y��}�B�'[���J\� �Pl�pF�!�4r�e���ϐ�i��꺅BD�[
�,̥P��=�J5�l�w��6�m��(o)��,�7�:m	����>X��8��;�R�N|ɑ����y���A��m�p�x��al]<
#z[Q)p�����pwjZ��6�,����8Y0H�yZ�:��(j�f����M��J���Zҫї*S�f4��ZQ]V1��0cK�����`���t���=yXh��`+-F�혨v�2fP8vec(��;l�̮$��U�������q�\j�f�b�	n��-sɩn)�`T�nَ9֛7ZCں�$�]w^�%�8T.�u�h�l�Х1l\Ќv@�7iSb�͡	u��m��mֺ#M�1h�4��ҷ]�L�T5�:&"�Y��Kv�˥v ��o�ю���ĺg`�a��\0��W7Fm����O�HMTvtn�t�j��e�.�[`їl&�[�cXfhW6�=�w��|��@�^��ͳٲQ��ep�޸.s�zn*��3b�W�m7��ջ�j��
�{�{��2�5|�C��1�O ;#5�x����]�(ϔ��sC��m��ࣈ[ӝ�Du��p���mD��������6��"&8����ٸ�ƛ�*�J�,�=�$*�6Wx=��oN�P�KK��A�^m���x�C�|�*��]̅{]s�p�~�2�{���֛h7f��0��2�G10�\f���jҚ��R���Ĭ�J$Y�QleK+�o4�m����q]sGrmD��+\_e��'�7}|���۶��q	�齚�Z���$�/Un����`��astt�����I�m@9�~˴��g.�΄��{7�}|�sb}��P&B�k\(�5{(���������]v��L��3`�]F�w��\<g{��d�b�-w@o�m7�}�p-on���%�l*��;����3m���/�&�S�b��<���ݘ3��؅�ZS��	c.��]Z{�n=m���8�m۬�sJ"=��)�QZ�{Fc��m�����a��m�U=2��sd��Ks/;�њb���HH���).v�ٖ�A��Q�{�tׅ�n�m�M��<��QN�Lb5�1e=�Qq�G���ᶀ�戽�N�s��uM�7�ݘ)����w9��xoruy�E�=%���=��ʹ�@7ٓ�`M-�FN�\�+�~t ��A�-�ò��ԭz���:��X*���nJvw^Ci��2�5�ө�n2���e�!BU[�]9U����w����Q,c���S�`��x��~1�!+7m���pC6�(��-�)����!ekk$�����,�ى[���l�Y7ʬ$���R�b+E#�ɫk�!T���m�r����Ø��H�SN����f w�m���V�S��3)�2pm��K��^"m���ջ����y}wO	���/�c���N�Ï`�8�X�y��Q����S��;��M+h>]�v�ϵ��U�P4gW$�dG7;b�S/9:Tb{X�iZ}�U��3/gZͺw(=�n���ܛ��r�[cE�ޥ¶ˬ4�d�bb�4�x��I�����vo��EO��b����/c��VML��\X�ݖ�k��N6�k��ulfW�������#7S��N�޺��� �i���qz^�1�0�Y�1R0��T�t�!o��{��}����]�������Z����R*�����i���r�����㊷��=g"�Q�:x/��G.v;&�{�3~���U��h�$q׼v�ݯ�Ό��w��Qb.�34�dsEK�|s�G8k��V��U�u�@ ��IJ񉕏�S����M�b7����T�Y�h��ݒ��(l���T%=	���Ժݻ�Eb�Ұi�u�Ď��ɩ�W]ݨp�]ёSD��]OR���������)��7Ǝ��R���i��t�r�fcp�4�g	s337��y����7����=Xέd�]&W����m*	h-V�kuڬ1���p�Z�s�2euA�͌c6f�ͥu��g6gluT�uZ֝���`9�V�M&�M>v�V�f�lo}m���3��M4�N��9Z2����w��]k�������L4�i�T��OQ��c�2�MV4c*f�fɴ3M�a:���Y:��a�by�͛�,�>N��UVa]n8��f�ަz�7ְ��:w39�Q�Gt�hY�s��:�W�z��k�M�q�*�i���og�l�T�j�A���s��d2Z�M�������Z�q�Z�A�Ӎ)v�{��-�M7�e��r4�VZ:��3�j6;��������U��s0fls�5��*���j�bِ}��<7)�z�wF^�f���}��^�kʹ�B���Ħ��0Zn<h
�c���¥�
Ģ����U��ʑ�S��a��m{�Ρ��W��V���l%�a���w��m���='�vfas�=��4J!"a �$� kb9�q^�t�Xj��a1���I��f �DAJ`e�uF>m��q|��/3ި��h����O�>�Sf�5y��q�6�����u��{P��Q-��.�V%��1���ܾ/����˕���6�p�^��0Fc�{��I��:�"��%�0���7y��������l�v��l�uZ9�g�e�>�X^��\zc�xkR�D�6�bþ���|�<pW*n�y�u�3���¯��	��.��L�㭛n�̀i�	n�;��ܙ�������/���m��
���ِ�T#�N�%���p�1�h6h�b͉}���~������FD�lr�;Rh]6�̶�rLM�`!���
�*��$_��}o��m�m�2��e��}�0����A�ϟs�;�ͺh7��mx6#��^�t�H�SX�;`.��8�w��L]�w��{@6ݺηqH�MJO]y���U��+��S¯��۽�	��
�v@�m�phB�'og'&��^jm�YJu��{e50�ۼ�rV�ɸ��V�:m��6כ}к�`�ͻ�ff���U�)k�[�Le�w���{m�6ȑP����� ����X�ylFz\��%�M{v��:��b�5�,�Q6^�F�Ϟ[Q0�ҹ��{٥��H�(:��瑅%��vf��]�i���j��U�&� ������5��]�9��[*KIcљ�y@eu�;LMB������W��I��e�`eJ� �f���#y"6��=���iP�Gkt���r%cv�G�e2$���d�Z�.lsa�.�s2��
�G	��4�!��(�I`%[n��1�͙�Q�X�]uMPf��߹��h�,8]������cR�-�e��b�e��Z�c1B"a����h7 6��X</w]�'w��*���h\����B��������ڒ�.]C��n��W0�}��Q���L.w��u7�'��l�!�Bk-|�7�y�۰��댗�)vav�.�ۼ�{�i����y6]�ͭ����m�Gl�����r�w�`a]��N��A���m �m9
.�=]k���;J�x�ݕ�aw���=����t����ԭk,#��W�=��K(�v�te��t��ZY��B �E0$��V���x7��:b��\5N���2��t����%�`�h6�p<�Gs"�Z��JVOT^��Y9/FR.�Fs5ҽ{ݸ��W_�ٗ@u�0�v��Fe��6QR�Ԭ���6�&�X��_x��W���&�ñ�
k��f�{�cM��坖Ue�*g�����6׃oFh���Vwt"o�J;�V)��or�z�pm6Ў	�T4T��w��z��GLWa�����s�^�d`d�;u�X�/5��my��Ko�p�������Je��u�x�q�K��ٍy��n'q��1wfG&#���j�^.pհ�af�T!�Ff�YY����i���Z]�b"���\ᶀm�wu���J7�V)�r*O��w;ٜ����mx7yn0f|��z�(��A�zv��Ε]��ۚ���݆���e*[�˺���k�Ǜ{ʮ��rޅ�,��k�9R�D���򴹍՚ofC����yH��Ǧ���8����]�Gӆ�ͳ7"��S�Te+U�S{���qr���u
��ꚟ�끘�m��f@2�8��H�¡V�%�����a�����{xo�Wp�5LYkeŜ��C���?I$� �Myn�{*#K�v	�k�ƅ�juO܀n ̏�=1$�E��/��7�Q��6�K�j��RL�]����\����ihj�7Qs'7S��r��U�ݏq��쪮��jx^&>��s������!�T����ϟK][�����^M'nTi�jaw�ǳ�f��`>�gb}�dfb3#9\���Q��&i���jvg����q����Ȥ�9�#a>#��S��L��{��䶭/!׋=U�I���~�n�a'�~(�w(\M`�3l)+s���g�cJ��lkh�-G��áBe�v�o6�gv'+�f)��B���9���W|��J��W�;zw��.�CRSk����8[���9qÇ�ܳs���Q스8-9�������
�Dw6�eI��F��ٚ%եj��2�R�)�j�#�h��&�܏�<k�%ɚ˨�����g,��ｽ��f҇���Iu!��؋r(F�e.+sNf]�܏$v��<���K��MO��{3)�u� ޿�g�ݹH~�h�o��w�n��~8|;�na�}�j�ې�d���d)Kh�N��h���Ō�3W�{����=��׎\��5	*CJK��H~r]T�u��tl=-n�h�p��O�U<:��32�=7��R�Z&R|�3;hC���g>��5��\p֨d������/��nz��X�|{0�	����Ľ�-X�S�R���f��=5�c��m��J�q�B6a���V�a�B���LͰ���]�\[t��`U�k��\v)l	�L$������c%m������Qj�mfi�BiE�бet��6��u�@�a�.{9���-W�%��j͠b�!	�:��t����x�G1�]�c%ҹ�6ʇie�:��݊h���Йt�W\�L�c�]�ήr����C`w����� Q.�]NFD�\�r˝����4���]�����fdĘ��$OLi��m}�31�������mK��q��^���ѡ�C:d��2C�̎o����]qc59���<+imO{���p3k*�o��X'�e�΁��@fF`;��i�sa�sL%\/ML��\<�fb̀3#D>�+�����ݔ�n'S�sP��}	<4������O��K���!� 7�G8�:�����{I���o&�$ff��ܭ���Ϟ����v�
���X�X�6*(X�b�Li�quդ6�EF#�1���=Y翚z�`̅�l.�"k�i��3���͉�R�+�eǆ[Y�3 �C��s���p�& �:E�y F�J#G��*L�hm�i&Zӓ�unڤ�r�����R�voo�\�j�i�ٮr"�����b��ں(?�^D�R�5��M��,�{�`��~���I"�M�q�
MJP�;n���#�����y �d�ffe9�ܻ0t��;�Ƥ�������v�y��fpqq��v��*�v���}̏�C23��:ku�i�^��Vl'n/S�S����q��r�9u�O���o���!簜ƅ�K�͕�Ы�fm��Jcȶ����z�l�m�r�g��w���%�H~\�s�=<p�V��^���Vh.������p�RK��Hi��w�I5,=�����U垫����/�.3�y���H���`�-�,��Ɇ��Էo��� ��L��e�OW��e��t+��}seCf�uwCii�ZسJ�ӱ�J�Iuչx�a�$��q�ݶl��󶚫ϕ�՘~�s%gB�س��-S�ئ�d{2 �ξ�c]L�Y���編���z����psW�{1���IUlf�3#2<31{25�g���C&�sFl��.wX��5��xu�y��3"^�2g���2��nص�����h��̶�ά``2Z�R37D$�IF}1	f��5�̏fb��v�N�Y�<�Tđ�pst3D��V��d2K��g�b�=z�{ޖz�Y-��2C�y�L�a����x7��]�U�p�Q����ff`̨�#�ѯ���
�綽p����y��d�UHjC��_��T{��a��%�4{�^�,v����}����s�QK�u�#Ozk��Ҭ�p�˅n2�n�|�د�����,�us)P э]��Z^U��s.�9�׈��UUw>����\���ԓ��ݨ,�1kGlW8��9�;���&O���ǳ#ٙ.ї�͘-�6b �����\ܰ�։�iSԲ;Mc��KiS���#Yn^
�:�7�ٙ��Eo��d�V�S�\Wn	�2�v
����2f ��8Sٵ׊tz�]]F���/_R:�'���k^̍Z�C���܀}ّ��^a{��6���3^�Y�|2a����*���5$��32�pܘ���7�t�U�ԡw��d�V���]�P�kO.9���n��3�%�!�;�pa���.'+����/�R:�W=�y�����t����U������%V���n�\��o.�i�������jއ1w5t�U���Z����vo�:
[�ܵ���[H�UKD朷aD䩭�s��)�W�:�ڴ i����%D�цC2�qQ��}���[��݁�ڵ�.s!\�{0�8;�ӂ[u�6[?�M88�
���>���zn-#A��w7�f ���}��ӗӶh3�WA�MW��s�����td�LD�3�u��W&�k�Nݙ��3:����R��DIvF�ZءVL�N����d�pGaR�ZMh�QpTUVP�4ETkW�Э܊i=n��˔
��ى�d��#�:������2f�������5__ܐ�*�8��n�	:�]�77�-���6�D��#��M7{�_H��Q°1ET�w{r����%�{G%��i��jZ���k�u�Z6)��/���Nr���4��̈́* ����z��j���*�i��[$Oo��(䬼�xvi�&r���[��N�eÖ��ئ�m-ܠ{aLV�u�ۧ�ͬ�p�������%� ��>��@�
$msB�vކse1J��o�Ji�dQ��o�edV]���2U���كCc���6of��֔Yn�eY�%�r�f�\����*tB*��뾩M����h�YRZ��&
���%�Y��yV��2�\���o�J��dJ��'U�F��^(�&1j��fd�j(;���+"ob
�}ЖfS�8�2쬛��5����4J��F�e�_SR�1o�o0�Ŏ�� ��I��(�ٔI�i��ި�2�����ɍ@���
@ ��H�XmQ�����Fpc��+r�ۧ���mZ��8s��68�z�1����`���`!�:�6�����jZnv60����	��c2Nfs��f�s� �X����6l�����1��f:����Mqj���9�fg>��a��:ս�wo}w�6��fv��a�F�6���Çfc���B�s5G��q�޺��ެT����b���ٻfw
�la�v;�c���5ml�U��Jn�ه=Y���f2k�dccY��3�a��q���Q�m5�llcpls�d�uM��VR���0ʴ���:k�ʲ�&��cI���&��uzyg+���s�z��ޡH��y�9E����%�H�f#a-Y�enn��KXD2�u-�\n�+�d����ql0h�Ғ�.+jB�nba�Z[me�����B��h[�h)�l�VSimEp�,�6��[4k��.�S8l�R� (A�Մ���Ķ��/�e��K3��K��^u��Q���ڀ�+��9�31r8ւ+��m̶�eu	��Ie2���0��R\]W���%t�c���7�[���c��J�m%d�K��j�&�0ݵ���fM����Re�tz��j��Ґ�U�bSuV�mH����f莶f-��k���Q91�av���hYm�g�3X�ћf�ۅVhY�.-uv�. �e�]%���4֤2m\	��P)���.�!]i^4u6�a8c�%H�6���j]J;l�0�2e�+�U�k:hԺ�k�жT�Y-N%N.c*��ĘftIa�ax6�f�uF�7lˢӱjK����7@`iI����cH9�`b4j�('6Tu�ȌXۈs��0������+��d��̥e�IE4!�)5	��q4�@"V���4�F;T6ѧ̗�;X�Z��%W`�j��z򡴤�\�e�b�(�ަ�^mS�֍!3s����$�E�0!f]q3J\�ne֔�M�c�Y���Q��-�g��Y���N�&����,H��mm�"� M6-u���:n�Wl�fb�9%J����ˣdL.�E�l6&L�G4���ìÃm�8�����%1*�#��̮�a�똦%iS\��.�<�������V�2V��F��� bѫf���	p�km�4��g0�Ԙ���Z�K�28$�L�[�[b��(j�p�0ZD�t�1�Jłj����h�ՙS�`�xtq�Ι˙LLZGYK���\��9����8��f[�%cfk� v�a!@[��r��٦q�L�H�<��l�$�q
�U	����N��
s�Lů<�h�K+\��gJ`���v^t�d�]uլ�6�+rV�c�<a煔�R�u��*�Tf�X��Ѓ�bY�n�֣I�[���Tj%��$�W�Z��SP��6�0�eֆ��J6���#Ib�k-r��ت%`�WbY�u���G[L8Յr,��- 2[�vZ��*�%�e�5�ɀ��f+M�k�\ˮ��X���5c�X�-�Xս�����)kP�U��W.,�jPئks�FT3��}��B�Ү�ԅ��Ek��p\�J�-FQ��-���f �"Q�|���6=��ِ=.��s�̾0�{���s���nǪIu!�W������7��>5�#w�U�{��0��s=���a�H��Į?	��U4�*u�I&}$�P���
��,�E�Ԏ���n��h��̌�A�����܁�Vdzv��s��|2a���b��YNOz�gw�<�'�T��It�K9H��g궂7�D�t�E���	����2g��nA�
� �!!H[d�`蕹M���ڍŽK�0��hMѵG�ѮP��x�܁�٘��΅:p7�'T�ځ$p^=��O {231fG�NӾ��s�fyr��r�n�D��w&�w�<EK���wQAΥ�˶��G��g��eD݌�*��.ϯ��UM�.���R�,�K���^��px��|���wO��q��%�d�3�n�0�f�¾݃�R��3ޞ����@fG�!�j�]�6��ۭ���.�<���N���'T�o�zj7��s9Յ3���2K���Hd�e{)w�`|s4�ڝ����Y��Cf@�o:�n���������|�l���K�Uҡ��0�V�;T��ѹ	�u�hD�ƙn���n�����{���Oy4*������-��r4�9�O�����g�I<��}�Ϻ��t��6�]��B�8��N���v�Y���f�tө�sh�2f 3E���2�����e��ܜ�);��A��P;1��/sj]ڞB�R�WR{�Z�0�5��#�����	���|���%bv hח��Kб�\������3 s�:�W����́�B�w����T�lL����R��vg9�MA�W���CRK��ԉez]���jO
��7��4)�M��7������o���wg)٥���Rg�%!)3*@�1ֳ<�SK3r�a�j�x�R�kvu�}t���~�z�^�@����e�X�.��6ą۾�WԻ.������E!h�Z��������#}�w��Z�\3;=��$�;�G|n��}��5Ju�~�ԓ�^��Q|v?<�������绍}�n��3 fbZ��p=����3#��!��W	|5K��^Ԇv�:�D\���Op�*ƹ���T���7���{��������lھ�I��!�'q���x6Ӯ:�W�豊�lQ�TI��}���K�5^�r�?T��A�i{py���y��������L�{�G�1�w��S����J���
� ź�٣�F�UB�G���h�i�4й�+�_^�I��i��2Lח���b�o�q̼:���/%�OzF��C\�:'v�Ȕ����zz����	����܃�̪l�H�� C�L�f�t�$��C!G��p-v3@w�7w;y�-~���l2K�I3�6Zk�A�Jg���T���5w�f�xM�]����5J���S����#NI�!�H�Sl`���{���E�;�~3��Ʃp�w!n=�3;7��֨NL]��Ԃw�&�[(
Q��zz8ED���bpθ����4$�0������h]d��"*��BZ*���E�*���F�c�tQ6�sB IB6Bͩ����7l3��tfGS\��
hV�PX�Ωf��ٙ	R�<f�bX��T�x�L�5�0dɕ���E�`�:�m�kBT�U�
��.����]��qb;	�Zc�Q��N�Z�����s4%��4r�a�e���i���k�XJ��MX�kk�q5�4%���
J���c+3]k;���{�J_��F��2�4�0�I�2���7wkGc����͊2Tx�w��{,�2 r(Rބ���K��Fz���\������H~��REU�'�C'���{ v�K�cˍ8�+eL�nǽ��ft�e�ʽ0Ӫr ��/�eq�b����ǅ��=sj���Q�T����d?I/�n�mm�S�{��X��2�B��$��늪�R����r܍�^o2}����axi���*i�Y������[*T�ݏ��� f{|��z��S��]&a�.�WA�5Ś-�٤y�&�0�"d�R%)�{z���œ9�,�{�3���!���x��6�O}�jCRK��!�3�n����V��� 'įM��,�YX+,��K&���nۥ{F�c����Wq���6���F�z���Ș�i���{�СKz!\����Z.��y�2A�Q�w��_>7��m�HjC�I6��瓍�?1�7r����nǆ��d�����ٴa ��{۵��"v�ʁݷ����2w��@=S����S�ER�I%}������V���ѢS�s��F�����P���̓ۻ+Hw`�� �*�0����uvt#�S��l�KBY���c��~{��zOϷ׫�3����YnΜe-S��)�㼎�����I/�շ��w�d=�.6���&�,����������#ٕb�{�-�����RK��z�B�b����/
Ǯs�=X�����nU���Vvn�&�'��F����>�ФH�f&F�x��D&��I�D��&�����NkѢvd�	K�Y/vh��2�uC����CR%��"�7]�V�8�I/���V[��e-S�ݏ3�������������I#۴���W�L����� F�}�P��6gw���C_I$��nm��f���L���Q(�L�q1�,M5��4Aa�������v�f��A������|��K����n-�C1-~�2s׸C61�3#ّ����8/J-fH��	���t�ue�:q��Ehn�^��ӵԗ.��=�3aj)�Sӷ�6&�s� �篽�K��	���&T��@7;��K��N�R�_x���U�v%w��3�,u�L�U��g�D%QjMl5,Dc�M:���OfH���ǔn���ntpѼpuǂ�s,Zݘ�)Y�PVgf�]s�KO�n���]Hd�}�`)������jk&���Þ�݁��3 f]��Ɍ��5�JL������i����Ě�-��k@t3���Z\��� 8����d��K���9���"_S�rV���6��_j5N��*�gvm������Щ_x��ȪŮ�����$�`5<m���Q�����CU!�kC^�6υC����w�\p߾���͹}$��9����1;��Ru��p�uD��:#
1����dd���p}u!�CRK��B�����X�W����T���P���f7�nr{�V�떍$�dͳ�L=�%y�n��'�yc8��*��c���<]���]ݿfx�|��,��x	�=.��J�o]�*,�1:�@BfJ)�RbQ�u�h'ku�3��R�F�1��Ĺm,͎�-Z��	.��M�j�[u+�..�#�+�<���Y��v�@�vk	Wh��k�s��n���
Ye��^�LBh&�fˡRki������l ��*Dض囈��ֲ��I^���u���usuB�w5j"��l�$V�׃f����ͱ#Ke�e��i�˥�7-ً�+E�>�ߡ5��d��p���&f-[Y��dV˅�٬�a�4қ��%_{9�{\f@���rc��;;��M�{�r�j���ӽn�I"�C��q�މ����y��,qR�tr�\(�s�A��=C����\�T�U$���&,�;=����w��n���F��$_T�CJ����8�N<����%�xf�vw!��eB�;b9��<��ʌ���zH���$sUI�s�W�y
�Ay��\f֊1r�܌��f<�:y��V��
<뢅�4@&�ktm�0$]M�Ֆ�x2uM��;]tFJ���P3s2�dyСK��u}T�a��'ig4��Hd2Fz��x�/r��!�}�9W��},�.s)�����e���[�	�R�����m�-�(�Qį�c?v�}�P�Y,\�]�BQ����N�N�rw=6ʅ��m���=R�{f��DMR����/�7|�;����p��Ҵ6�Q����s2|31fG�ʊ���a�dO��C\f@t(R��-�0pH��3T$7{
��
�F�9�R�]Hj�~����k���)�y'%�l�\;c�Y������1]:�`ߒJAJ@��Q͐m��TL�Ի0�*NqK*\+CV�B.��_�w� _@����ZE�=*�G��EG
�L�^���~����%�H~�F���4Q����ꉥ��{�ɰ�U�wC��d���<���s��!��>�����&&)*J�x�y+GL@���*,���&�`x�W�%��ҍN���ͮ�����[�+��R��/j�#Vt��L�k�ćnˊ��P�^�ڵtV�R�*�%z�M�5S���Z�N"�\{��2�R����+H2���K��|�J�'�6�D.Ӥ��c��9#N�����[w�^>�ӗM��r�A��- ^�VX�y�M�gV�&��-0y�v'Ll&d��d���6G��oo/��y��^q�;J�bцz�#��l͢yVѤ%/q���q�/v��Y���lkŔ�"���V�'hMV�B�ui���F�x\Y�1��A��g˻ܮ
����t���1���g*숋��ܫ�nˏ)����;����e� *�����>%ށo����R�goTZ����9h���E,�=r���Δk�W���wdy��SY{f�8�F2��B��i���Am��Nj�q�gY]kMg\2nԘ���sG@&I���yCD��in-�Cn��;Z��a�n�}[Գ�=Y �`K��Hn��L���0p���p�yrT���;1n��ww�	o2����3��A������,ݺyѩ�v�Pu�e�&�s�a1�om�ȹՄ�'pNB4]�����N���9�����1�*�}c��J�!�w\vd�^pwF$�jbƾ��f$HU�GK��;XГ%��u4�,�
#ˇ�^��1��F�,����;����g[Q�ƭ*AZ��s�~�t�f��B�hAV�H;6�t��m�35�[�X�i�q���Fv�խ;�����z>��m;�����y�eL����i�o:�n�͛��ᱯ���[ަ���6�\fK4��[;�����N�7�s���=<ʎ�����כ���8]w�o'%�Nӧp9�N٘9����[{3�8KV�1���������q��:�bJ@� �F�@$��5�q�f�s��t���Ì5\���ǫ1�4�f�T��p83f�71��{&ӷz��k7����WF����5͙��ͷ�:�����^����w3��sO�ٙ��9���sgq�xu�J���ƀ3�pg;�W��z�qڒ�����3�]�uCv\����4�R5T+h]�g*M�v]�8,߽ƫwnC�Hd��ݑP������t��׳#�A�z*�G>���}^�;��_��Y�YƤې�~�_��/-1=��+���g�~���?1d��H|�B#\m�����f�8r�>���共n�XDmꡦ%��&ڸF�8��ƴ�!�/]�q�ܹ�'����C����_t��[j}^.��r;�7�|�۽B9t���~s�`` �W\�?t/[As ����L}�T��&��9��>�
�������p���x������qΈ͂�R�>#m @/` Cm	�n<�B��a��oI��_}�� �������Fj�~�7�/�v-f��~��]����n��p��ԁ^.����K�+����#���` ��^6���Liɬ�,�Z
�Ǻ�T���i
��f�KCU�-4��֎9��L��橗W�ѹ���B��p� ����׬��`���<A	���=U����7Q������H��"� A������C�u\}�/�W��-Wt���C6hm]i5+��i�2̆�q��l�.ҰfDL)B>>G?��� A���d�]���7�_w��@�:�9�Ǵ�ڽ!�n�ԑ�1*�x5�{B��\�/���z1}5�|�����%�������h�O� G��I}[Aۙ��hD�_o��6k8�U�}���F��f����A�����-� �א/8U���nK���Sr$����]pE.���_��Mp7H ��"):�m}:8����ŸD[jH>m[��O[dwG
fT��[z3�/���O�~���7A�q�F!;�
~w�IC�8f�۾�[����<�Jʄ	t��ӶyS�L�|��sR�R2P��,�FEK��v|���l;�dI/�at��E4	cY�.�]n�hA��f�56G�.4m��)k���7W��P��*�F퐬�Ŗ�e�Z��Të��[����D�ƙ̦V�4��Z7,�	bumQ�&�ŉ���y&��\6��R�ԁ+���U�Q��lK$�j��.չt��h2���;j�.MKx�c;c���ĩ	�Uf�͚]���m�1Rܞ�|>|L�R5ԭ�ь�M*n�Ь�"8���������;S7<"��	��}��w>-�����V�@�}�}1{�|٭��}��ث���tz�mH!����/R����g�IFt蓹|�=U�k�o����5�7	��B ��o�w{e�jM8{�h k�Og)7� >�m�����/>��-z%O��C�Fi��W����@@��dO�p��������L@T��FF4�z[B���� ��ᮘ�}���$u�/x�u��Uf孮g!x�~�^n� �nD��^o@_r:Y_h1{�'�>�����k����	��@��n��6��؍I�B�%|%(�2�AɅ�1������h�-�����a6��[4'��u���x�[jo����8����|�ߨ����}�}�@�A���q`���@���A��{�vRs?7���G��]�ú���Y�³�M��$�It��9�~�;.U&��y�^�/�ȃ׼�*`��v*�rb�0Tyb�j�e��g��3~�>9�!��?F��~��u��|'~���A��~Q�ݠ��Ԃ2א'�A��� Am�[��T�������1{U�w�5���$�B�"s���7k���Y����I�+�#�/ڻ�K���3��W������N`��Ռ�:0�B �h"s>n ���m�/>��@��U}����ހ��	?|	��b>�����W��[i��p�K�)o�D��iB���5�Ц���t؋	\s�c.�]��0Q
`Lx苁���D�D��x���k`E����5�������H���;�0��`=��ӈ���Ŵ-��d'Ro�ұ��Q��u�芎������U���	��n��n2�WBT6����1ι�A݄ 6�!�3��^M�ʼ�1��O���FX#���o�������h���6��Í����f4z,�����l��S������K4h�zgQ�޵g�ofH��\;z �u��|'�� ���-���Ԑ��)������! �B�
��"�|c~��O�S_W�}��X{]3}=;8 C�3��Ax����[^n/��@�1/v�-�u,�D\t�z/�/���O�@����wdH-Ǘ�@���'����[(_�2o�% ��*lE�)C`XЭM��-��fK��.���R.���	�@�� ����_��8��|��?P7_(��#�b�;��:Mi1{�(�[j|Ci[�#:����^����qΏ/o�*�"-w�W�_Q�#5�5k������l�mO���<�y��� 6��Dښ��~߷ϲ �R8�Ժ��|�<�?}@��p���,I돬��>��A�A�O���Wq��Q��?`5_(������=���'߄8�<93���S�����D��b��a?���N�07�J׵wY���⍊���	QTnR������@�~|�������A�nD���֨�����$�Y�����k���f���${�@�7PD6�|@m���q;޼y?{��\ek%Z���nɚ�9��/
��N�((LDz&A���^�{�G�����n(���R*��=���5�W鴾
~v�~���r�>��?}��ؿ[@6�	�p��}r�f:���@���O���]Ɵ�)��A���D|A=�) �u��}�9��ͺ�~�U6�c�L�!�p͹�� Am_]����E�T�-_�M?�����A����D6�O�mp���0k����y����������Kq�k�����)�{��������c�j�V��q����	n�����$�u�c��{�A��~ʤk~��������}�Ӻ�-�>m��{�;?\��Z�e�L�n]���
�;]�h���]�����\u<�]w}cj�k��g}{�i�g�n3������s70��*Y�x��bqm�eh�t�S[�.��Fl�����ʪV;r!��BWe�ŵغ7��tn�0H��K2�K5�m �Ѭ��4�ڱ,R�#������5��m�.5�ɨ�45�ܺʹi�S��T�rA���B9�GS.��))��%ʂC�FV��멜VrU��:��@nJ��̭Tv��B��i��0����[�Z2�tn��)�O~w߼kr:�:����)�&��h[�7��s�Lj�5���i�:���hC��4'���[��+������.&b�������[�BF�=�-�|Ch/� A-�$WvLC]\ٱy�}��	}��`|��.Sq��W���>=���$��^��?��8�\�� ��6�O��Vū_8?UK�ۚF�u�U�Q��o�H݀�q�mI�r:*�~̓w=�#�����݄A�h*�-}�����b����� E��gMV�[Q��z����-� �[k�A�O3Nfɤ��-}��~v������r9_��pS���ۛ"Kp� ��}Q��<�I̒�d�2e	
$��Vb�1 �[���2��d-W0h0��%�h�.���,7Ё�m���������Pk~�G����]�|�`�Zk���m. ����A-�$6�������ae"��f�Y�����3�E�ݜ�L�0d��M���n)�b�y���,a[�M�U[j!F��E����s�=o����"rV�1}?G}��a�3�5H'�5�D6é�U�3ג�v<�׫���y�_\���R��aLy����y9�U��)� A� A��[� �s ���Q;�|Tw(`�؂w�"|�Ud}MA�ߔ�5_%=�)":����:>�1�v�����?o�Hm ��-�[����BT
��b�}�_|2Ԩ���C��Ёk@6�|Chn�뿣{�d�A��"$�FHP����c)�:��ٖA�hEL:9-�M�m	L5)��W������E�@������(�����+��S���n8�����b�Df@@�ā2=�YcH��T��*�}>!�UYZ�&w`�~`���|A=�/N��O=�+|Ɵ��G|�>;�mȒ�y6��ǚZ��	����5�D�FFo�nվ��I�5�z������t�,y�����,�1m�u+�Ns�R±Jm�v+�d}��� ���"5�@�����-� �V�N������ݟ/Ubǜ"	m��;�&��L�u��1?	�� ��"p�֚gp?�x�� ۱>n ��!��m����}���Z�3�t|���(��ݿ/N��qD�Q��]�>TF���"�{��K/���,������G�muf+HV&łKb�DL
�<"�/}p ��Ȓ�"��[f#쏗}���.%E�_�(/����j3v~�U@�F��Hm[�A����폇�"���l�4����"��Bkt�G\�s������$�	�	���B��Gn�	ބA�w���m�����+�ϰ#���Ў����Q�{~S���q^ �ڐCh!_&�Q�|r��:;聤n����������>]�_ò�T_W��B"{>��o�1�f[�q~f�:���]z�����K�NmK���_���t�V��<<�{ݷ���m�-z1#d�鵙~�c��|����A�	m�!����vْ��rT�p�c���럮b~?=� ���$��6��k�1Ϭǭ�Ϲ��{UA���\��R\�e��獠JĦ�����l��J�u����BGߪY�Yi��y�*����e��=�k�Q�SŴ��聻4�����Am�7ay�����;AO�;���ﾁU�c��V|>ˊQw���мA�@��kz�ڣ�����$�^ ��|�����Am�޾��W�mFJ�S��;s�g��=��hH-� ���| qĔ�}���؀���p�����:[3'��_J��A=�)#v�Do
�X5�>W�K��@�r'Ÿs�!�kwFt�d�[��?e�(������x�5��mȟA��}�ok"��ؾ�#c33I���������p�1S:�w�(�%^�AY�B�3WqQ��:[�� ��Σ� ��n\� d���*�uN��K�U�y`������7��G��: �s ý���d��ze���Z3�h;w�0o�a̩Yon��s3�xKw��޾��ԅଷ�`Y�[FM&�'f��EtiR��H!d��^�S����;��q�ڪM��Zo)��m�� M�B���v��%dwS��d��U}����GJ�:�����@4t�ɸGu��Bo
�)@-��y��:���v�]K/�gNK.k�5���ܐ}f���6!e�hx��7��pu�zb2�z���L�j���sl�w}�;{��+�
x��������7��Z9��)B����]��K�Vrfh����e����6�mk�e17jn�y�1�P����5�t���k� g^^|������4��X�	���f�-j�X�5	�
�C�\����ﶛL�;�5����������DH�6.�3uٴ�D�S/"[��m�O.��U�I����z�ڙ%A �%Y���{>	M'k��{;@�㥣ai���5da��5E�����n�q0V&g]���a1 u¦�y����ˁe�c�p�_q�U�����J�,�Ξ�9V���Նl$Evmws�<o~�s	F1nőy�^d�^r9z�b��asN��Lͽ�|�Yr[3w�����^e�F�t�ֲ6�Q�kY�g D��ݜX��po8��F��veݓ�v_��5��{�yv��R��ڨ���mҕZ�b�#4�YiB������w��]�U5�g9]0q��j�V5������]豜V�yc�sf8&^w�VK3yv'OS��gc�3&�x�u���w�f3b����2���O�f6`�f��V�N�{�da�i���{�랬0٬�xǊ���yW���hy����٦�]�}�5�2���m2hǪ���Y��.�^�ީڴ�������ZsՆ8�odt�Uإ�5�1�k|�<��1q,8��@�7�lذ���h)%����6V���WP�W�0�{^�9�sV�Md����y�y�����x�Y�X�y�7��g$7�������-5)����a��מYT�}t�|��T����l·�xl�����1���Ugbtؘ��`C�^cӘ�hl�	�u��ı��u&�+,eU���j���8�FF�٫Up9��8R�c��j�� �؏Ps@�e	B���-u�Ƙ10�8ֵ�YTZ,��,�+�A��J�f4���t���cFU,&9��D[v6���HAҍ��<��0қ���[p(��":;�Z7�у��6�=c��g�+5HO2-���X�@�٬6Û�sq��5j�h�sD���hr3�3���m/Ä���8�j�6f�Bne��M`B@v���)U���:፱�C%�B�1���YL�t%���֎�IVU�ѐuR���e���n�1�Uҁ#��M4���R�l��mĵ�e��KZ���`�44�Ѝ�4l�R8m�t�(�&�ccl׬s� q�ea���X�`�K�ڔ�&f1�I�`��C�SQ,Rl�	y�]tM,�Q4iU�d8f͹�R�qUMl��0�G��Ҫ�P�9�Ku��
BXcv��Gb�Cb�D+�����"���B��ʜ�PsU�]��,#�if�&���Vd%�ZB]�р�΍ջ���Y���-xQf�h%�����9�ɪ���f�]��p��6�L�Š�4�Q�J��AlYe�1���lcF`z�mr�i���T�{Y�h��e���9���Д�JF�lƍ����I�6�4�턫,WX쒘�ZX���%Za,hƉՃ�7@��B!�X��v�^u%��j��u�ښ��Վx�-�B�� ²R��ZniI1�n�#4�4�G�!�jk��X�l���W�-Y�E˗�s�͡��V������[��23����.�55��5��cP-Z��-M-�8m�	u�r%�!0��d���a�3�G@wW�cX��f3,,i��[*٦�vH�ga[���\3dkfp%���66rR7�Yn�h5�L��Mu �L�j�fmK�!@4ڑɨTz��c),��M���`;	knr�
)U�P����5���-�GrB�v���Z��Vm2Ř�٩���[�j�G1������v� ���ǖ�U4�q$�0�՚�K4MiM���	Q�[6ЫbS�,�ʲ��+1h6�6knckE�0M��v,�����:���5(E���WE���RYse��r�YJ��^�n
�m�Tn�d��*&k�m��/XB��3]+5q���áK������/s��6�Ɣc6���jZ�\���]��Mڔ4C�A~���?�Q�K֤���p��������7S��k��L��t�;�^MEe�������<�mm� ����E������t��"/�z{�R*�E�N�fd����Q���~R;�"�uT�+��������5mH"�A�� ��H-ǐm������"����e�(�����/�W햝�t��l�{ڸ�����
w\��/P@�мA��U��s8�gE�|�>������Ҿ?``�p�#�D6В� Cp�m�Ԏ�Z�w�l����yE�;陓��F/�G�����A�	m�jξ������w���	���Y�Z��Euiyj�R
��Ԗb�t6^vD����.q/��F[������,�|�����ﾷ�����]T}��y!p�<A�Axod	�mp�|�RUY�'�@J��GR�#�Dc�Y�@;r�Qn��v a������/Zs�J{��2��u�4~Q,w�e��"`+��I�?�����(9�j��N5ʳ����~��� ^��Ȓ�wwՙ_dE��Ax�����/������oD}U�}�Y�ו3'l�dt��v��F���mO�m:>.�2�v�(�+�8����1�H�w�[���_���$�BC?Ƿ����q��du}"|u��p� �Ԑ[Ax��C��O�T���� ���n��jq�Y��|%G��|#wdIn6�v���_�y,������H�F
7W�F�b5�Ѓ��@��Mi]Z\�\W%�b~���o��v��!����w�_c��S&���*=����߳cui;A����@��"(���]�to�\"7�![f>�.ﭯ��_��� ���<A�j���O�t!�ӝ��n�N��Hm�[�A-�������k%�
�D.�`]gujiH�t�N~Eg��S��lnv��[I�Xf�zr�D���'C�^�/�;C��%�aA�e��=�3�?�W��}�."ff�=�\Fw�Zw�ѣQ1a������O�hH��/�.���G�D���o�Ag���N^}��ep�{�x�o�RCk�[��A���D�P����ML��O�;�}�^/��_�ա����l
���6�T����t�����}&Q���mQlֵ���+����E�3��ְ�S2���|���}q��n ���ݞ�Üu�]������CD��=�}j��!��B ��^!���Y��!k� 콟v����.n�)��>��L}��ߔ�wPE�p���{V�9֧�cH�ۑ �M��֬����hLȥ���n\R����~�f��!��#ͯ7Dt،��ޣ�y� �����ڑv{�9�Q}u���J���۹j"gb~5B�2���I��<l�h�ig3 ћ�b���4���J��W��S��������VϨ�FW_Y�#i/ٞ�r��v���#�գ;�#�Ѣ�{�]����B��������1��/H�Ax����4�/��ﯦ��yf)jL
ʬư�u��@U��\��j[Y��S~����|�@���7A��
�_!�}�^/��+��+��/�{:0��h ���>ϗ�6�-Ǒxԑq����Q}�4?�^ ���E��6�E�W_]G�W�~� C^Ȓ�} ��dut�%�l/|����Я���w϶F�3y
wnܥ4ɍ��L| ��^��-� ��S�@!�#=eJ�?
���A�H���^�Z}G�}q�Ⱥ���e|$���Ϙ�U���|4�s���y���j|Ampg爫B屧�T֧�쯌/���*=� }��'Ÿ@�hZ�*�=\db����Y�*���L}Ň�oC7\5q�"��8*hX$�vo��D0�W�6`��]�Zk;��O[Գ���5*˜mҋn�����BZ�VgKm�lf��V�s�uE�ΆGc]�q�V7$%�����ۻ����4#]SV��$��&��[T &��W8نxۮ�;���m�ʒ�`b�	rd�V�Q����F�cq(#A#�6�ܹ�%6���q.�Ύ�ę �sr���郱��v.zٲ�eZnV�U+�2��7Fe5S翰�~غm�5��qږ��ƅ
�e*IN��r$��ig�����߾��'�Ax�܁>n�7г��JS�L}�����.���͘���V�A�Ax��A���7�����R��~�܏!�B�¹}��>yw3��>�?}��!������~h �����Ǜ��h�߾@�Z��L�L�=b�2���Q�@����"@-� ���:����
������!4o䳩���&>��T|A>�z����9X�iޏ �5 ���"nD�����%�ߐ\8p�]˫���e\�«��>�\Ne��u5��^��y���Ǟ�'�����Yl
ȭ��ѱ2��q���.�fIs	f��s���<|�o����篙'��7��ڛ���Rػ��~ɏ�/�F�|~e@��$�@���@��� � D�?|&F�ܔ}շOsim��͇����cB��𴱂�����)ǟ#K�K�X0���t�E_]�k��X�ro�;<��	�TY�Fb^���(���O}s?-w�䥃��������uy�т�r�{I���TC�/�ۑ ����J����DȲh?�|���yW3�τ�~� ��!�"|Ch/��f��蟮�ug����A�-�>�<�-�����1���@D$��&ͨϹ�<wax���6�|�"�h"u_)^\m��B��Y,�������-�~}��"=��fQq�j�E���y
��瓴4�(�%"P�%Vm�tc�[e�V ���^M�����+�K��܀�;�"An�UD�+��.���q�u?
��H�&.r)oۜ*:2;�v�^#�ϧ�6��^ ���������b��b�H3�y��:}9�箇%�Lp��@��� �wg���ٞ�À����-� ��@�܉��hv�ٓ�����ﵥpm�=��i���R%`і!���N�f�]&��n��Ge�<�� ɀ�.��!-��C"ِ���%o�ٗ��: [P��7���b۸�?EG��|���7A�m�!�6� >���t�}��H9�y�*��W����}n2���Yh|~��m��᠇N@�f�E�����^n2s���JB����
����ع��~_FG¦�?}u�-������\PU%gP�RjM3+ca16�mc:\$�z��j�@�d�鄒�Pg�~�A��{ CngŴ*�����,o*s��]x�飝���E���z�m�!�����,�����㗗���<$���TO¹}���������V_�A�}�����d�}�L=��#�m[�"�G��j�ު'�y�੮�utd|*~��^Ȑ[�6�!�"A��m�up�A�m����U̙_
gyS���|�>���/cw3�fX��TM�.���q�3�љ�����Qw~6�ߡ~O7������8VK��Rv7O;j��}CK	s�8;:2!:̨���������i��f�6���n ��"|[�۵i�g�x|��'Ef�w��_���O�k>	��Df����m
{o�ߗ��տ�����L�&�M�)�c�#F͙k�V`3�c��4�����'�,���]:��p� �ڛ�o�lL�Q=_FG������<�"^����$
̟oE��h"r'��9;T��Vk�o�\(����
h�dʟ�{�N~����{�s���)}�Uez�Q���v�`"nD����ڙ��<3�O���ߨ�f�wS�Ϥ�Ј9� Cmz[A� EÝ�nl�u/W��G�"	m��g��8��u��d|.~~�!�cRd$�~�\ƃy�� ۿH ����W)1��:>��Q�}f��S?#��i��SM@ܾ���|[j���m^���O3��m���q!��G�%CX����RĠѾ�w+�͕�"s�.Txw��2��}ßb��'�V�E�^����es�{�i��@eAu�3r�5���kb�K�K�â��^��W��uf��׉�&�-�"%Ѭ
�n�X;-s��q.ô64iv�Wj�����my���.�ʐ�Хf5☰kb�Y�aPF�M���n�jV�h@�7c"��ۓ��1��m2S0���!K�ڛ:c��"�f:j�[�I���	���4�Z�}��?�o�H҆����+(�͸��6\�2�1��^�3�qm�bL��~��&�o�[�/6��CEr�>�?e�����}"��DC��FG4�>�6�-� �ڐ?1e{w=�A;�M�:/����z������~�n�-�w���g>6���Z�s�$�4!��>m������2'�WtL�I���N���Q�� �����-�>m�!��R�@��w�p��!��C��������s�Ϥ��衼�>���W_0���^ϠYn>m��6����9�΋+T��b�c3;ͮ�����^,_�E���5����POgM�<>�IY �1�+�Fy��/y�����39�KWB�t���B��X���7���&��ɉ�/Mb�Q�x>�A�߫�b>Ӹ���p� �ڐCk�[������'�{_�:6Bt`'7�B��C/�� ��N�<n���f����b��-���rX8�_t�$�A�	Kp,�7^�Y�Țn	��"|�
*;��Q����s�k>�O�G�h"q}x�`KLͭ��)��;�I6�-� ��N���Q6}�;l��
�����{����'Ÿ��h Cn}#�4g����� ���k���
h�̘����n����=�ϾRDO�ޝ��d�o��� �r�H�m�%������oݪ���9(+7���7]�1�?Y�|~��!��|�썀�*���̸�:ǚ���7�լ�P�A��	��.��5��1QP�P���&�T�}�/7%�������k����#�s��{�f�V����}w�$�B�!�r$�x����h�=иh#�ϧ�6���e�O���۩��:�> �s���������O׍{^	݀�͹�q��^r�����q��S�z����)030��W1Ɏ�M'����'��mo�vBл�jGV��Ip�y��c�j��/v+a�`�چi�s����-��4��aT�W�m
�����oQG�k�TXq�U��W6��Ɇ���W@��hnIh��Iw�� ��Ut&��t)��Yyj$�M�Q���W�v���r�>�X��UfC�i���n+f-B��E�zw[�λ�u�6�E�}�ɇ+�I�rj50�f��Rr�H��\:��n�]sp�Fc���Q�|�Y��[[��=�+[{���݉I�Xx-8jn<Ǝ�e�c\�ZΫy�u��Gc}����,�e��f]K��w����I�[��9�((֐�&ZL\7p�2�cD����oS;qlGL����L�ϔ؅bT���f�����; �X]�a��2�mJ]T�;�:cv`��xr�eC��ξܮ�s�P2��u�S�O.�k#kX�ŉn/瓊�iX���O�z�-<����a�o��袸*R��IM��Ȃ"��;,9��j��o3D,�5JRl`)�÷�T/Kڰq�w�׾�{\��aD�$��E��B��T즟gc�}���A��%W���ed�B�T*���,]�=r:vGA�PjZD�{h��+��ݓ�5v{���=DEEu�9�>�7���H��E�;T5�;�n�A��"��ˊH������U0�hлC!7i���ܒ�)�F�K�v���w�+�50��b�M�䵁���[�]���<�C�,䔟��7��zf���v�C�Zrk��M�]�'�0¬��WB���7����V6v�m��NcG��&���eh����f�i�ռ{[��W1%�xy�{P��Vl�ֵ�#-��S�,�D�kz/�V��V.����i���v*��*K��a�µ�[ك3���vW�oTWk� ����{�ޫV����Wei2k�];0|���Q�����Z�7����o[[��vff��gղ��o�5m//��u[�}u�>�Zq���I����I�+��q�}�kc��w��kHlsּ�;CՖk`k��>��|ѝ��o����f`�MS_=�U,��n������ف�o{-j�3%6>����Gz�5�Ide�Kql��4{+l�9)`�*��i;�ĥM��5N�s��#��k1��e�{3��s�5�L�l2h�Y�SI��zڷ�j���b�i8H�}C^\l�S#.~
��H'�[Ar���E�DJ����&��x�7^8��ڟW�E����"���o@�]�%�W=/�:�^.�x��CnD�[��m�qF+������$tX�&'k��6�}SMG�>Ͼ^�=A� A��������9�#�A12�Q�1�*0jC2��1���1�
�Y�U5tDsm���������qd7
���GMWI���D��HX�b��߾� ����gŴn ��RGѻ����΍��>.�OcR+ע�Q��p����\�����u	-����2�:����e��G��D6�O�h>���{_}_�Ui�mV��UG� �������Ŷ���C�R#>�:XL__�'�:�h*��}5C��k'�_H ��G�FOڍÝ�a���r��܈O8)��䫱R�6^�s�j�!�C|5g\�PY��K�[R�-��so�]�v�32(�Dܸ\>"�g�ﾀ�n<�-�>�E��n��S����m���y*}��W�]s����{�+��x,Gޢ�=�А[�&и�|sL��&�FI-���63��c�S]hc4.E`�[��L�~�vH>7�y?�@���|@m	����}U��'��Q�#m���Ꮦ�n ��>-�>!�>-�^#/��Ζ�<KG��
���GL�����_zA���D�Cm�_�ٺ����47Ё��> ��Ÿ@���R��ˈ�c�q�u�NL���p�a�K?]�����Ȑ[����mȑ�
j�L�}s�/}p8���m5�s&>���6���>��� ��/Lݻ��UF�mI����>mȟ��{>���%��)���>{�o�)�G�5������Ј8�@����� Mr���p��-<B�Q��(��6����)UF���wY�/d7fg�����
�`B��s����%2��8���;ط��J!�W`έ�X8�]�Up���]h�V��W`��JF.u����] �a
ԅv��i�D�L^�XFl�2۶AF���k��32ѭK�]3�4.R� ը�e��h�Z�t�D���Cs���
5������]J[�祆�ј��R�M6-mJ�:7��e�$�35��z�X饰7#�/,�8Ү��e6�S��k�<ua3�sE>�ϲ��
�fq���D�5�n�ҍ�Q]SU5j]U�4U]��+�u��2����kq�ԏX숿�0���<~���O�[W�}��ek3v�"��	: ����	n�ߟ_t\�8Hg/@�}>>z��q��}F���êc����> ���-����eП�.z0�Խ_Z�� ^�[�Amn3$��H�?|�>��OI���L� ���ycAۑ>-��-�e;�+�k�\"��lQ�mH;"/�:��<~���O��������p*�7�v�3� CnD��@|��6�p�8���`���咝��l)���1��?��up�>-�~��~�.�d!P`��▤���kK�s#i�٠LaA�k��s��\�ZtԬ+ܹ���}���k���od�GG�\%|*�����#a���G}�vlz}��39z�h p��mI׹;ޱ?m�ό��p�`�������t��B6�1�m�<]\r���Y�f�)Y�\�u�
���.v]�Qvc!d\K2�a�FW�N>��56>Ȋ�`9|����S�@�����n��t���c���2	{�� Cng�6��Ԭ���}YG��X���l)�3c�In��n ���pн<�u)ʷ���O�ly6��'���>��W	�U���$�Ј�&�7�����Io�x��3�>h [���mI6��#�M/�$�׺9;8�s'��Q��&>?	�������y6��=�Ub�6����d!���B�T�8���eAr���⍷LCb��ɦ�M]ч}}�ߪ�3ݲӽ�j0m	�W+�����L�:f> �����D�ԫ�{�ڐCpn �,�=�.�o	�/|�TO���GH�s𫯄L� ��Ѐ �9Cn>1q�A���R�_�P^?l#���H-��n������%�|������x��Cv�~<�c��=}�n+^;j/#�n�6�KL��N�*k;���H��W��+�ӳ��6¥3v��H�j�,Y�!����L��@^?�	�n@6��#����*8�3�Dn�����R�[�3���|s�RE�en�#�y��_r���[��AmȒ�Led��+�*�A�6��\xe|*��?	��A�r���М�?v�YS�*���HJ%H'X�,���t�d�+����%�ln]u���-�o2�H���ϯ9I? �p��mO�_�6�(�툎?�c�S�W|��00�9��v<�CnD�p�;�	�gؙ��xP!��>#9=q�%.}��U?�c�A9������>����?]w�ݝaQ�qu*H��>��܉�n<�B������;k��+E]|"g�>��D�������ۯ��_Hn+쿯>^�ϡ�mX���A�{���Lp�� O�@@�â#�������}
h�ʏ��
�Y��g_�'�n߽x߅#�) �]ю���U�]��lm��|�����S�J��V�J��udO��q� 栈m���@�h"x���Ъ~�m �����}pvUO�����R;���-��=����݇�L��ef�&sK� L�SM�.�J�-�6QE�������#-��F�>��$��6������'�;�}fn�3�/�s1/���Q ���"�@���qD����R����A��^=��A�+�"(p=��q�&8T�'� A{�$�)U}�'~��\R�p�A�9�΄Amm����>�W2h-��E&ePw�Z����|&�T�^�7 �כ���g��G�}"O����D�����p��M��&~����g��o�u��|[A�x�<[jHn�n(P���Mr��D['a�>��{�cz����h��Չ����|V�&����g]��	w6H������y
^��RQ{{�F�٢�bs��<���kT+om����'�e��*Ho��T	�����>5te)���l�����j$Ы��%4�5�B�Zb��4U������BP�]i�z-��fb�,.�m��).`�C�X�Lu"�n��Q�S�ɇ7Qe��᭔�ݢM2W��.�驨14���M��wX��
n%������*��[a�p��Á��j&����֚۴IY��'�3<�[].�
,�C
:�Ֆl��2?~ϧߣcH�3�ԗ,���K�-��]��ژ@��h�Gq�6����i�}�p!��^�6�����m�p�U?�c������8�\�m���@�Ё�mI��-�D;�5l}[�k���5�~�E�?B��r���� �� � �m��Aj�X��ml A��$�^-�����w/��tgFũ:�ts��]�U�z����X��f�=p�n m�rca����ԥ�k��/� GoO��6���@�_���*���1���A��ft��/��3\>6�xA��$6� � /���7bwdWϢ>�lpnPq�V�Bh�\��3���s�^!�"|[B;�D���	8�HT�LJ���C81cfE���.4���Zl�g@�\Y���;�{����@�6���b'��˅�3*~Uv�΍��|����\�/a[A Cmy����Ze�s�g����a3.��f�i��4ECMq��mp�kEja�"���*n#`:��-�������Lyq���:��._�FWL�:��8rW��+���0�}��-�q%�@��A�#�ۑ ��� ��g���ϫa�˛��~��B � �!��q������J�5{]�]j�y���"�mO�����C'Q��T��=�*e��dV|Fu�~5��>z�6�H%�@����=��ʧ�h=�:nV��|�?���ڧ��-�>on�W���g%�h'��� �H#~"�
3^ieu�˗\M�%fE%e\�:d%��%���@���! ���U�WЇ�|%��|%O�HW�udPW�Ѥ� ����p�p� ڒ3���X����ѣ�*�ꚱ�"/����G|f>? ��� AvD��s�5$ح�Z: 
۹�p��!����f���D�ԏ����n��sN�dۗ;Nk��� ��aI�67j�Ҝ�$�T=���
���q��8\��[�����hM�|�/6j�����Y*��'G�1�� �R݀�n<�m�!������_ٰ8�������UC~E_��/�>�w7_	S�}�":���@k�Oǀ���>#u[�|�S�h/���}[8?}K���䏾3*~�Ǿ���DЗ:��L�3��t����&�.�9ԛp�0���n��TK������%B����c{�5���m����WF@�C���:$�:�>m���~S[����A�@��A�m�7` Kp#~Fڽ5]߽�ߪ��Yz��]_�o仾34���S?H � ������'�g}u�#���W��e�@KmfP�05Oµ"!Ud��LG����ޯc��6�������"b��#���>!�*���nW#ݑ:$�:�> �|���oxt�q��Ef}Q��j	�x`�s-	�41r�sD,G�=Wd�7��!����bW����'�
�L*pC�,�FTa��x|}���)!�� AmȐpBW�������f֮��ʧW
���?}�p���Z��Z��ٜڤ3>� ���)�A�dA��8v�Ű]s3
胪Z_�疍Ԟg9���C ��R>�Ax�<jn��!��G~3
����?n�C8W�8�[�:�}�CpnĂ[�Cx+8D��K�z�8-=��6�y�5тJ���O��q��R݀�n0|����7�^�~8�"nD��|�
�)x��\����VV���5.��2����!�>����>���U9���V ���͵>��b"��D����L����f����G|.�q���B�}�"s>n<�m�o��Ϸ)W|���=�o�B�7M�G�*�#�e�N�C�U��9�O���  BI�rJ�!$�P$�� @����I?� �	'��I?��@���$ ?� @�����x�@���I8@��O�@ BI�I?� �	'� !$��$��!$���
�2�ʜi�Qr����?���>������9�@ 	 h    >�   
            �>��� Ϡ H 
$AQ

  D�� � 	P*�PE7��dAT��"��P�R��R���H�TR�A�J*��(aE ڈT�I*� |U�(��KcT�2�w��[�SZ��T7�k
�}p�.�%J�@��厍b+/�}os���P|A� ���`}נ�;�����ϯ*J ���*�5UP�T�T�{_,u��:��}9��W���g#]k��g�;�Q{�;��c^�@��_L�T��vҹ|��{��=WM��ͫ�c�ʺ}t.�ρ������7,�����$ ���ڪњ*I* �U���\�}�>�/.�S�y'�U�=��4�t�jٯ�����*�f�g_@y��E@0 ���������I��x�N�U��r��髵&�¼�z{۽����f��W���N�I� ymE$(�J$ K��{:wa�(��;�U7����v�w�v���]�]��]����ε(��  ��WZ�w�$�;�.��A͝h:3�kz�5�;�z�1:��:\�ݺ���E{�U �*�%P��5��ݺ��v�g�:+7�@��7n@{��oC����+�qI�w-�J�����^]t�Z�y��;2�Z��Խ�:�zRn���ƪ�6b��       5O�%*� & `� �~F"R�I�=M0y@�0  � 4�j�0��F���C �l�"4�P        ��(�Pр�  10 $jS L�Sڂ0M4�L�4ؓĞ~�_����{�
q��tcN6f�ۛ��*.���0DC��@hT�
"�AHT>ˠ�*��H����y� �����o�ҟ��}5�H���(;آ� �(Xn@= ��>G߀QC�yЦ����%A
"��!Ȧ����{��5���G��_�?�2��ϵ�	��ĒI.I2I$�	$�I!�H��E!�I#�I$�A$�9%I$�I$�I.I2I&I.I&��MkZֵ�ּ
��������"� �+���@�wCpU�Dwq5�WqE�D�V�p 7q 7 7]�Wq�Qw]�WpT�SpU���*��.⋸�(����*�*��n(��(n!x����*�)�8�	���	�)h�� &�(n(��n�`�n ��n
��� ����`!������x"�(��nૈ;�����x��������!�����`n&��Z&�"n��
n*������������!�����;����8��
�� ;�x(��*n &��h�n ��n ��n"�`����"����;��7��Zε�[Z֯�IrI�I"��$�C$�I*I$�I.I2I&I.I$�T�I$�I$rI"��$�H$�G$�)�I$�I$rI$pI$�H$�G$�)�I$�$�I$�Hd�I$�Ir�I�kYֵ�ky�m��GU~�[	����O*?U��>���y��,�p�CO��  ���C��8e��ʛpi1�囎fc���B,���re�6�5�m,�y�#O6��)=�71�JҢ�T�2
ܬu��d�C^�E�Zn�/a��,�f��j�Y�,[�R{w� 6��!n(�uPK)0�:0�ֲYw��ҭvuZق�wTWw���n�=Ul�L�Kv^n�:�n}��ލІM��v���%��������Z�2���:f�@ ��'BJE-ں��;� ��B��k��R�m+׎z�N�`��p��de5Y�.�:�t/�:V $�c�"V��%�XZ�Q��'6��n+�[���זoe�:K*�Ү��E{V-=��ym3U���w�l���8$�F>ֱYj��Ly�u�I�2�Cz����z5X@�H�c��rP����#"�L��R�h����eʘ��z2;��.��Q�Ŭ��ݕ[XyD�t��'d��6^XV[zJ�xo QR�n|r��ܖ��r��1V�.L�xs]�ô5��KtDF�i��%�YS3by��w4����s�i�Y���١��kAM^�.��8&��;?%I�t�]���5m��������+[[��Rq��.VHټum
����FM���:.�7�3�Wv�	ђ��"���Ӌ yH*�-��VhY�h,Ň4����vr�*�ջu�L+yH!
��6�+�הw�+r��L�)��A�6-�b��y�C/
+%f7zSh�ܻչ�lm4n��#���v���{�mc��=�v�;OF4�\����T5��W[�mXA܃��أyy���(��6�;(�mfX!ԕa::vū���
������Y�*(uDT:;��hG�.��Yhԋ�Ù7J f��%k�h��FѢ(V�.�FKY�w��9HKR�m�t�ޱO-�*ַ��V%	�j�Քi-�0]��n9b�L%����~�6ަ��uW�n����k9j����q=V�llr(�h-����)\�嘕�y*d��ǩ��dZ���ow$�����f��(��i��̽�W�'���L��05�B5iY{�ށN\P�6�0�:<�,O4�;����u�8Ka�VJ `������Cm�.��+I/,�3a�ްm�'�;u����aJt�r�i�W�yN�J��4dyv/F���Vj�̭�Y4��$��1�a�A���<kR��$޺$�5j�N��;�l�ktճOǌ��[41Y���;�ֺ2J/�mFZ�-ޙ�+ϴk�V�lsX��ۻ��ؤ�,Ւ1�W�(Y�B+kҖ+�h팔��T-���@��ب�.k%�i�LI���R���+#�E�qK����"�JT�A�&(��.��o!V5��Ż�"oV��R�u�H,���k"�-̠�LN޺P�PރS0������F8M
�:�u���C���=Gy��)KyP��2�Y3y��6ͽ�ʖh���=�Gn�k�SE=���8�kQ@����hF-mh�,�İY��ڸ�� �m��є�M۳�A�&^���w���]fU�j^�_nAg*
��9���Z�T0��]�R�IV��b��VUn�;��k�Ad�j��ѼDb;�l�Ͱ�Q�/$z����h�HZ�2�Kώ7��)��;�w{�B��̗"�@��!#�t��c�]�+*;��U��re�\Y�i�L5iܻ87ne�J�\�m00�)�h�/-J�ŗ	�d��6��ٷ�h�ׁ�7%ڐ<9V�I���!�j4D��i�A��6l�n,�V�.��t�L:FQ�Y[����Z�Ul�SW���)17YR�f�������tXeV�x�����\"/.����gq2�k�����z)^V�n��'P�ˬ	�n��dlѼiR����n�K,���ba�˃ٝ�����^��6��ԫ��e��S;30P��$�^��Q�[��[Twc*�r!L�f��a
�SrwɅm���V�{Q`ʚ��̊���a��wZUM��HU����V����(,�y�F汊92�m®56��FBwedB]CsI�
�pS˰ŦXߵ��Z�r��6�b��q��1��[�ʸ: @XŃihf�����%-�9,Y�I�+[m�m�ŪV�*�7���*c��,�5��Y�*��Ñ6��Lĥ��e�t�Mʏ 7Y`Kop,.*6�.ac%��]A�r�d�I�2�+�x�*�j��N:ǛVd�L��̭����䴋ַ@�mՈ��au�S����`��(�׸e$����ަc�g�q�|+_p�c���:�@Y�-R Z�.+�)\�Foۖ����nQ��C�VD���fBRT�BB^T[���7�6bsn�vaU��Ԭ�Ѳ)ql5[��	5��^�꽕y�cq}� �($P�Op'����6��Fȣ�
cu���;Ƀ `��ٛ,(^-Â�YKiB�%
��o��e�dw���+�v�vФ5*03{q<�&��,�E�ȵ�^=��Qh(�W�P�ce�� �wf���6�Y�	W!-�TSVV �.] \B�cT�+E�jNO��k�՝��%`�2�7j�@�0���.�1�$��]iT�'�1�s4��ى�9�(�=P1�SDeCyv/oV�����+�%�U1�MLWZx˶�n�p�y�Y�Ż׺��w^�@��c2�S���4��U���������̥��ig�(��*��͘]�ۺU���"�JK4<�*uW7U���.ƭ�	&"`��bF���,��f�"�b�c��X��d".� /P��]�EX�F:��y��k3B��H�ܭ��7�ćdyCK�L�(e�R�8THՔqL��[�E�&���.���j&YT��-F6�m�T-���Ma8��r�j*N�XY��P��wP}�a�v�ͬ�Fi];/~B�e�U�{7Y��e�2�켏u7�qX;w�m%��ɪ^�V�@Ś��M2'�v��pP�/�9��.�e�x�-&"f�Vl�V�&Bk�3	�r�ٿl���q-1�R	0���ԷV��ê.]N�i:����H^k�FZU6�۹��}��o.��YSn�[�\�x/��Q�Kk�,J��h�Ѯ)�sCv�c���ի�C(|
�2��?IQ8.�� 7kfܬ���&�p����4��EmAf��U��M̼ջY��y&� U��u���e��o�pV���wE:f�S�E�������9+6���eXH��Un�mVRe��d]b1�$�+v���i�%�R
nW�A�V5�1�9Z1[�vv�2sqKŹyFeV�s.���r��l�d��Td'o�L��-@�#��b@͏wIR�m�Y�`ڻ�������ӕ����Ī^KH���2���fn�n�]�(-3�r�9(�L���,��Xø �T�4�怵U�)��Z�խE�C6�7�n�9&V�0=Y So�!O`�WJ����iD��wk!�[m]J7����ڎ��-�Œ�e̩�W��k6�Z�����B����;9:i����,]�ñh��[�����Ó~R��R̰qB�j��D�H߶�b�lVں�dک�B�ç0]�)*�g#[y���Ve�[��<�Ww����qeң*&>�3���m�V��xj�����qK�b�{������7{e���E[������Z��W���6��pi�ʰ-���[H8\�2���{�lٛj�j-;����e�-R�fK)�ڗZ�#r�ܽU3p�u��Ԭ��h�,_۫2�aw�t��,�
ƍ�m�l�P�I�w&m"ˤ՚W�rŀ��5w�'2�fiZ�Ov��Է6�a��	�3�[xVnn��kGh]�n+̟nT˭��1�]dMS�ʗI���`�e;�&�u-�������B��c�,bۼ��/hK��cR���$ ���u]]��sh�R�cե��M%����6H�&e�*T��w#�4ayG2�ZIVB��¨c��ho$���/
:r���o%*���*汮�ȁp%���xr����ܧ�MCg(;wqȀ��n�*����b��CQ����X�7nGX�Cx�Ձ�E���e�W[b�f��Yb�$InJCw ��Z��a�1m�n�2�]ݪܥ�bJ�L��c��s6�Y!q�ɖ�$u�Ҩf^����f�kr(,�8N3������fZ���in��gY�n��Uj0��w���5ĭ�+�o���*�|�y���Ώ��
�Y,C&�Q�J���͓��0�Q�4U�r�4nU�V�C�Pَ3#���`�#��x�r�K�G���2�珗����]�/���7l�{|8n��v�s+t�<3.К=� �ݸ�n�I�˽�\.+˻ļ'���ڦI �V��|�w�:�}i��}{&���F72����y�
��2&����c�5Y�L97�^S���[��S3?8Q�����O��Q~O|������$���k���ܷ�'U!Kj6Y��x�|�_��GF�hTW��QdPBDRDdAVABE$@BERA$EP��@�U$ 	D$Q�IBAQ	 T�RAA$F@$ �T�$@Q�d$ Y	BDdQdB@�P	DT$  �DE�T$$I$AREdUFA$IQ�ADT�DdU$A�F@ 	Q�$T�Q��*��EdT
�O���~���ey������%��DAxIn��}��[UA;ϧ�٬���O���	?�k*��g�~B>���I����z=���jJ���1�$Y��9��A��w��`*���سc�#�|�R��]ѡ�C.��
׍�s�͙��cΌ��f�� �}��YΚ�*�2T�}с��F�;-̕j\��(��2��ӲM��&���+��Ӗ=�f �[V��_�GWTnTx�ze�gb��G �l�V�븮���f�Q8Wr��</vj�Y)$�Ύ��oFk��ky9,f{��U�;Eǣjd�����ۚ��ֹ}��1����t��>8ɭv������t�kD��	C0�趒�������pv�J���1Y����M�w�P��D���wM;��r!�]+�Vc��j�lv�����$x�����i먬� ��l���� |����Mo$�+�ٺ�A��.1�o/k\bɶ޻�wum��=m�m6�m�i��"m6�onm�m�n.Rw��Y`�|�I��8W8�54�r�R���0fӔ�΂�W�2.-��ao:Ӗ�6�2���UֻDYT#�h���7���9v�py$��95ֆyYZ"�`w��Fgw�]��KRm'� v2�b�khq�O�f�F^u�ܰ쏚���WL�G*<bM�`��ج�m��v^�2��h��[ݔ�#�^�Du��Oy�=n��6���[�o�Y���|]Ũ}�v��+)�V�pY���ܡ�a1�/���»���%-RJ��jko
�Jl=y�]�}��xb<�஡wO#���}܄�zsj�U^�T��7�ָ���ެ�Ӭ������a0�Y�ڱ�m�k�,\oY��"��C�ȚS�����ֺ�T���/5��+ e.�)��+!�ʣ�׫�4og^ğfEHv�9C�u�_1w˷���͑�:J�{��5��,���oYm��z�m�D6ۆ�n�m�m�m���"kfK6��֬�o�U�iB�Y}�3g_F��7뷝ݷ�B�ni2t�3ѕ;GA���P��>�$ۭs7�Ĵ�e������f�b�*�zG(�$�
�����}vR�ٙ7ú�0���|�kX�7���v�����ڸ6�C��M�qn���u��ذܧ���n=�óhZ�$��vR�f��6���S=��H`�Ԉ�j61S:�v*�D��0���p���:�b��P�;:�F�轵�J=Wn�[�e�u�l��-��L�G{��5�+��N�/j���I� Źp�w�X�	��l�);�,	��jn��TVj�d]��i �n9�kK�V�'D��k	�*{�R��f�b�	��n7D��y��Fu=f^a`��c��oB��R�����}4�C���mT^G2d�.��Y�z�m��m���q�n[m�m����r�vW�wr4g��<j-��!i�*i�ye��[h��O����K�;�72�=��Q�.�mNY�jܳ���NXX�f��Y5��6�;Z�C;3�Vޛ*������=�R�u;*��Dd�z�6n,��sb�݇e�Z�;�|��;�����c���v���i�n���FK�WGJ�W�I��c\ޫ��<ה܂�i�S,[.n!/�׸b��Ν�P���m[�D��Ep48��*$��vJ~�.E(`�"F9����V��4�����x�K`\�Y�,`���;��yT��uo����S��vU�5 ^���χh�� �h�\����71�/�(��D�ݕ��)rs\�hS�4��P�*(�%Ʒf�@�6�r �C��C�=�����k/�Q*%č/%Y�yz���n��l6�m��mÙ�m����oM�����doh�����ΗjZ]��e��#9��\0@f�k6��l]�]��2�pǼ�,�obU�G�n�ws'c��=��W���a�O�Ѣ2��F=ޛ�9S��k}*�C���ȫ_c�\;W�35GN�w�e&*�&����W�Wgݴ�ַ���f�TJ��:�ԤƭTV9�F�щ�'%h˗�uo��#r]�>2��o�������k�v�ڃR�˼U.���2f�4�7B�vm�����t�F��}"k9^�jl�vv��	b��{|uؙ�7�����3%ͻ֔K�4�$�i7���d�!ܱq����S�9v�ev[�����n���o�'�S���b=�\��F�WwLx����2`n˳D�Sj�tTE7gd�V��)U�������g+�(VQj��(ӎI{St^�	AZ'Iٗ)�Z(U1��<��Ц+L��g����m��6[se6�m�i��m�m�,�փjy�3U���֙��p�"�wi���!YN��\� j��]�{�,��{ׯKSle�J�z+Aq�M�X�W&V�]o(��u�J�v��q����X��YY\ZL�d������Z���tku�>q�r�kwmc�q�8Բ��*T����j:ɢ�����ET�4~�n��8�٧b���mg�J�P��4�m�e��@���R�B��ՙ���8��)�	
Z��5��ugA2�;�B��6�����c[:�]���sF��]HEr�e:6�[�Z��䡼a��$T�M}��{�^ �郍�)�N%B�so/$@�%��!���&����f��6�X�Lٽ݃���.�4�=G�sOv���j0ݞ�ĕ�Z�>7��Z��e�����;Kn��ǔv���6��!����ޛZX�ݝ��RE���3!�f]�+��WY5mcm����ݶ�s0��m�e��m�m��U��}�Fܬ���vJ��]�H��wZ���rT�;�l}�Ke��wv�)�5�{7��}����������j�N��'��v�k���"C_K��9T�BU��N v�l����M���#n�����ZF����:[\�jl��Tq.��2�t�{ٷ��zo����00�2N���M�
���6���]��}��>�g]<]1=�ZRĬ�|Or+4I��^���ה�m��o����@wz[O3+�nt�3�-y�����Z�r�_47��%hyY��ڈΙ9��k��riѬ�}|:')�^X�����n�f��d��n�e$!����n��أ@a):�K�y��'^+�% &�kr�}�.���Rgn�Ҁ1��H˭���v�S�+&�]�Ї�X�7����ޝn�GNJ�dL�T�ubkV�-��ܶۦۇ30�m��l6�m��M��xV�l'Zh�yN�X��#��-k7j�,���Ř3R*F򯥛d�r������7.�9�̬-\k]մ(�t���OG�C��Dn1��#3�n���3�'�jz���ق���Vճ����yf��]���B�oV�����ʽ$����8��ǘT�R��JZ�w�Qm�x��+�*�6�f�D_i��#� y�a��SrJ󈕯��Բiz8V�ĵ��s@��z����=�}���6i�F�C��0��K��s/��[�%p/[W����
���t������^f���U�vft=�m�/I0(L�M���Ѳ���>��'��?ѷ�u��ޡ%�|�ǵ$��g,L�%��:nWe�[�$^h�q�]sDF�b�o[&�%�!�-�ZEmvQ8�V�P_�iiX�]�v��$Jø��F6���Ęx����ݶ��vۆ�s32�m��m��m�m�.j������FWs����.�Y"�,F�Ηq^�`*K�N���P��Fّ��fM����/��v,-wZ��whѢ5ps6�J��4�.�r�_V^���$M2/O�t�>m����_!5�E�t.�t�]|�Z3���(������y]��*�:���iތ�ޕ]{n���z.�I����F5 ���A�;ǷbŇ!����٤���]^]i��3�T�e<�`�V!���Q�޴f�\SP��(ʇc��M�;٦����)ͩ9���N�]ay0٭�q��\���fA����F�N�zo�C��T<�#���N�p��7�Ms;��w��)k7Jә:��n�i�R���׶-7e]��t�^�.'�6�ú�U��_B���9�c����5��"����L�#.Av1���[��K7��jCM%`d##�k��	�iҶ�`�6g[J��jrv�dӼ�ط�'�6Tq�GV�np���Xe��X>d����]u����"LХ�jX����g�c��+��Z��Un������*�޺��(r�:�N�I�6L�o^PQ��Z�nw#bmݜ2�!2松�w2O�ƸeA�l%�� ����e���ѓl�T�J+������>�N<�r_E�:���Fw���b��ؙQ�Cb��ݨ҃�W�ڭ�9����}���]+��$�BS�B�ͳ����HԤ�].��*�}5�sP�L@�����]�vr\'�ir����(�7��=�TFJt�L��N�H���Hr�Bf E�Vv"ZZ���]��n�)٫R6=�k���~��>� ��I��
bKbTI�п.�����H�̧��@@�C\����r��]�Z~���E��2g��p��5\BL�5nd��KT�kå�r�l�i��M]�զhf�C71Q�l�5�&�֙�l\Shˡ�S$�L�����&�j��C��XB�]λF��`0�35v�������3�<��� ��ٷS9[E�4�Ma]ر�6(P�+p��6l%%����Ŷbk,��R�m���P��+���\���;X����i)����C��˝
�����E����R�h�v���h���{�;ҧZ�L�4G��[�my<�m�)c�`�K����h�\8� ��b��pN�R��g�8�0��uj�嶸q�С`���B�t6b�v^�֡,�ѱ1�4��V^qn���.%b�e6A��c��,�K3v�aXn���s6���B���#E.�Ût�㙛`L�:��д�8f�ԉ��E��-��,� �;��k�1��a
B�ĵ��Av�3��*̛d�*\�Q]�V��)��2G�n��`�vi��T[�k�n1/:h���+2P
ڮͩ`a[�����K�A�SGE��U��;�V+,7k��� Ty@L\��Gk1cvYe�372��Z�͖v��E�t��J�h�K����t1�ͫ��x愈�E�L���ֱ�mj��2k�5���[�-ښ���
4�!�U��'6&3�qVƻ�{���f8Ǆ�2�B��mNb72�	�M�:�UٖQ���&�� ��ν�	��`İ���4�mb��Z��5��]�L�[.�j�mc�W6P��.�Vض[S�Z*�с`l�"6 �\ˍف`��K�0LM����q h,�+KX�c$��XmPC:�KRf�3i �e��9�1�s�l�)*�
�q�I�auV�MJ:��t" f�v��������SF3&��T��4�6���61	a/)lYWF\�s
:�v�Zۃ[UX ��"h�9)��z�r���(�m
`u066dP�\;�V$�l-�9���ɘ�iK��t�ƍ��V��)�*1i5A�i�85�]A�®��+���&T�e	�\���7 �8 ��l�5�����7�nz�j��W�3MQU��+�M���Lö�+%�Fiu.ch��SM��-2�s]cl.�dBX��
赋��M,r��5�k�;s%�̢�A풚Xx�>���#j<�B��*�Q��atc�.1�g	�5iR �f$���ї����4�Z�Z��m	�)D�b�%�r��[��I-�d�
]��6�5���,��,"�Jlm||�Le��K���vˣ�pk.sn�,����;8#R�Mh9t�Y���L��hm.��d7X0Dn��B�ҝ�-��tKMv�ѸN�ּU�Z2�Ɍ����| by��[k�Y��9�6����m�S7e	l�6��H��4(g�@T�+�U��6�o�4��d3�t6�����%�C�����R4�V�ƭ�%ɓ9��F��̳d��B�%��fȸ�`괎l�%Bk�.aZ�0�]��]�k��=v����E���$4z�&�b�X�®�b�h�5;5fj�k�ؠ�;&Fvp��m�$�ˢW.@�ԦQ��f	�!w	z͂�L]��Qk�β�M:��R��W�Z�L꺖8��\�#B�`�j[q\3-�A�t*�Sk�!ڀȝc��3 ��B0���Jb��.w���O�h::ƌ n��q.��ɂ�I��-4��)3]H��KUW`���C\�c4�vp4�#ܙ���q@�$t[m���U*�-GM��sP���ҋn��l��"�5]
�w#f��-Д"И%�&WB��f�P���A�]RI�6��[�jӊ�s�slkft�4��-�!]67��Sjm�ԛg�Z;����ZKɣ�3;3ic���./6��Rб��:�*Me�a��٘i�.˒Y[�;�V,Ĺ���P�̠B.�YMt���kb*b�-��`B�9�b����(Չ���A�]칍Ҥ �B�γr��HgYK���dmߛ0� �xFղ�4�]HH�G(X�2Ě셦p�!7�n���]� W(.#�Bf��ɭyEU�[*5&aYh�Q��iX���q�9����ױk(F���9rihL�\�B�U�a��L���k0M������L��[H���]�)m׊J8��Rգp@Gc@͎!Nvl��)SD��Ⰲ�is�0�k�R�0�I���aÂ�	ìM�َ�����:�R�lG"ܓF�d���qZݨe�%#E���i�볝�ՙH8�Bc�쩠�
�W;hi�W*m[�j�n��Wf�mYv��H�4tt@�������.��F�M頭@����4[,�"\�B9(��Ҙ"孕�k�l���+����1
�gF���� ��4�ˋe*�f�B@���
P���L�fin�Àɱ\���q��ɡT�-"8���.06e�asK�KIrOU�_�V3/�:��1q�K#+�&��2\�1�(�*�X�2X�ņVm�1%���U�@..�G��<�Ka3�����i��F�j�R�wsj������c�L�kYe�,�&�ؙ�j�n�f�ЦsA�t�n��R݆c]��p���-6��q5v�ћCh(��p�аm&e1�8���l�u��膄Ы�qn��MW:	5�����,r��]�lfni�
�k�6-�3Rݠ���<G-�K�^�)��X+j�jY�WG���Ѵ9[�����*�����ܭl�q6����*�21��͒#�+.��ie�a-;���]c,�Wa�2Ui��ۘ0���\��UW"�Y⯑��[X���.cnR�\�l�!��.kt��d�I�ô&�(�5�@��8��Zl),��WGg]�l�9�r�UUUUUR�Q�UUUUUB�.�@3�*V%��#�4h��u�f���.�6*�t�m(�b�3ku`��u�]�92ۈ\���[��]]�*�T"J��v)�2�ZŃ� ���v��4�ۘA%�U�|�D���_)RD��b.!!"
Dd�Դ��\o���V\���wG�e�v2�*"�"Im�A.U�.!.Z�&m�7�n�Oal�� ��ւ��:�V����fe��e�(�����N�(����iR�q���E�d��4�Iy��ꊺ�lahJZm���Ym���̗�ia�ww�bvMKli9%�nYu���jBH�2H�B���9���F��k#Y�J���,��	�p��\�����!#�**d��"�	c)�1.�%��7SnY!*]�Ǘ�F���EinXݐV�q��#j�)Ui�I�I�=yo��z}K�
D�*2�]s�P�,��h�,lڻGc<1X2����aP؅��`�c%�:�p�V��aNU�����D�ųeɢk.3�Ȓ»V^x�]�в�i1i#� kmh��R�����(:ky0���-�ur�%u���1�9�Ҡ�楛�D(�źZ�5�[��mr����a�qεML�a��7:/!�B��f�u�?<ZK�+�Ͷ�I]���f�M
�����v��Z�������b4�Z�SQ���FS�F]Zq�M�m��Z�v�n�Z;hj9��Tx0��9�����)�εGq����i�b�����VK1T�!������ h�Zd��ء����캵1�[� ���E+S;h�FDt%U��Іc��u*[]D��3b� ��ƥÔ�d�51ck(�-�.���6.[-�k�����طR*�8"8�l��j-nik��ZE�mt��T!�.ٕˉ��Cb3b�x˸"�7F��U�P��Q�h�U��=��x	�cP�3X̂,y(�s-م�+K���4eD�j[uy0��)��a��Z4�b[�����B���H����2���6qt�ku�w�Rj�n+�uzN�6�-��4���")- ��D�Z�Ҋ����:��­�l$-A��Aj�,�����-�Q���x�	e-�ӆm`���)m�YZ��X���m���(O��,ʖCa�a���Dc�bbP���r@x}<���R�U����o�d6Vu��3��V"�T4���]忭��$�<��h�yR��]���m$��|k�[���|���{��4û��v���j��UV�G�;`���#��r�h�t�6ئ�s�z��{�ކ�:��ۙq�������ѣ�����ۖb�A�(����X�&&`D�[\�У
�-m���B>���Ӯ[�L��^�eٺiz��.��f�B�U��AgP�X�z�j�r9��'���ݽ5�WW��5�U�ݝ�[��}vc�l���`��g�yA���i�������{���dn��G�[��ZdR;�_�"KLK����"=Z�3�y\����n�4�RP{v��[�N���E�<��{����F1u�Dk��I�ғ4ZB�3��`^P�9x��i���$~�?=ݯZ��xbc�]ܐ.��|��$'zC{k�&������_N��=ij��p�%���e�U`��K�#g#�GG���H�t�E*�7�]�n6�J>s{�rs/�nb�7ޜ��h�gd}�L�o>lu��P��$~[���W�?2=U��d�'�SR�$�U�F�B���[�ٚG��v��>��{���w�ɻ߿_=�p��k�6��+�@fU�#.�fY&��ޞI$~Ë�ޞ�=���y�Ԍ� _Ay阵���	�?n�Z~d{���x�78�uJ���*u��T@����+������b#�hl�i6�8�f����g9�c�=�k�X��ى�C.6*2�8��}�Y*�^Q1��f.�ƫh�X��ygg��-����M�׃T�ɮn�}h�-���iUݚ
�Q�t8Շ��Wv�R��[�6q�j���^^evn�����-�n�٫G�����n(�g��~�������t��{ƓZf$Z����pRE#I�=F=}�llU�Gwf_}v�H�62�q�u��v���&:Zy6��_2R�$P#ޞ��~(���zz`��SV���"u��{��ô�&�Z�ϡe(w����:Z�r��ݦ�{��sw�8x�����)�8�cl�35���j[ґ�x�-d�Z��Bl�ų\*:b��a�]�ȸ��rڅB@r�n3d��J:�\��&��"R�Ϙ�6���-���`x��	f���8⭁��-Ԣ�A+[��v]W�����efJ�+���9CkZj�11)L���4}󘾸�o�;+p8��#���zy��IoER���s�FK���"=��7��u�%�"��������c�=3�z��ɪ�H֦)[�<볺ic�۵�Ȍ}]�<����g^����+=�;���"87j�S��u�2�T��VDDl����]jV���8�3����rj�3OVx�E,���zt����Nm���OK6i�����+�r���]�	�����綸�k�������̵}�w��f��RWSU�0����~��:*�h�m2*��\�X�EVi���5L|�v�a�OMٻ�"=��T�����3��vc�����̽��w��g����qe#�[��,V�*���u�}�6*ݣ���!�]��u�w-^��ϐ������̀�ZJ
�����T�3"&"s��ܚ5H�����$@�Ԩ������1�|��U6h^�+s6�C4�[ٶ;��w�K�OGi֫�G͔������>���R|����λ�MV�9��]�3]�������8�T#{�[i�#}C��#_Jn�v_�5�K)�"��;z�[��{�.����/l�ƶ�EX�	?P[�t�\}�{����L%�]���ބ����ySw��{+�,���ff6�e\����9�x��=z:��#f���MЪ��.���/��L��޷���ATܶ�qo��`��4�G�_�M8�컈n�������n8䶠r�?!1��í?3ﻇy>�7�^��ͻ�3P���!�"���nRQ��@�խ�%�䊷{q-���p���&fE	ڿ��O<��uT�|0��	�����~���[��37`cPi��
�J̣J�&fP�����Ë{����pW�F32���ͬ�.Y�-}8u��pn�����bJ��Ui��\�:"(��N�7n������� u �$��v"4䘺�=�~����^~�F��O��)1&r�]n�;;���Om���Q�V���9���K�s�G11����{+�(�b�7z"�ֳ�.5�2+(O;|�$�G/�O�D�J&T�Bc+����Ւ��1���L�R�8��in�^m�!l�"Ü&���S7+GY�ٌ�\,�YF�٬R��tɋu�s�f��b�Z�sM���Npv[�(#����u0J�a��J��.���=���v���ַ7Ų�����e�]��~��DN�׾�>I�~RV�>�۬J�+�ԇ��,�i��=7n���,�,�t����2�ܹ<�e��U�q=�{�|���i�L�4��g�߱{��NK���>X�����e5�%�o�O
�
�v�<�|�����ک�nm⡘d��H1&��1�)�#+M]�(�dD���9��`N�V���{,�l�ֺ�*�+��I��qU��[��c����Y��x��ؤ�JͶﲤ��x��Y�j
���7�|��)�3e����^�ŏ(�ޗ{���©#��Huټ���3���V�f�ydp֙.�o'��/l�l��8��K�)�n��r��=�w4�"�`K�.�M�F�֞I!��jF�S%�,2�n�1�\��ġ9�=�5U ��݈��rL��s�w.?L�	1g����ۊ��e��Y�ꞡ�&��X3S����u/}�X<�ҠZ |�������Q"�r`�};N��b�&d8�b��$��&E�k�R�	31�\ȴ(��2^�8Ñ3�eX���m���g2���WU�/wQ�l.�8*+V�w>�wvU��]G�6�ڮ�t\�L#2�kά�ݽ������ˮV�ӆ��7S������7�֞�\7�C��P���YB`�N��嬳1��8��z�VAM�s&���f�ǯ{�y�V�P����u��͘�����	3�恹�����h<v�͝eK��Pkft@�Wdp��C�=��oM^���/ʕi���]mB�&e]ʛN,�۩>��2D4mq�G	�����;Q����şqY�-*T��������W2��7>����t"�م��_r�ٛ��`�� ��]��+f]�lӿiY�=�p��ά�r�v[�K��]��&��;�pF��z�f�bd��r�,-�x��<
�n�s %��Nһ$o�;.��&)ʘ�J=�N����m�$�E��^��oB��g�2�z!�y�H�w�9�Ϊ���HIR+$�Q��KK��lZ�9}�6��r�)V*K�Le[�-1��[�i.o��4�Y.�K���`�Ȩݑ�F����_^�z�<���;�̠]y�X�Qy���S� 6�j��E�I�QK�Q�kd�8RJ���u�l�[�z�tc$	�V����p�%��.ZG��C28����b�ȭID$	-R��B*�)i`z]N��zv�_9���Թ����P�Ym)(@i$e��7L���kl�Z[A+{�֥���ݱ������̍�Ui��w����&��=�b`RB$*IG|��}���[�q��O����,�m�ha��*P����	��+����M��|�M@S����zR>�v��R	10�d�b,�ŭ�s���U����o��*$����o��&��s:��һ\
�r��B�]lG��:t�h���#��r|�ٕ�0�[���UT*�e�xH��Sg�9�xkC�ܧ(fM��o�2�wcM�;��^y9�^�L���Q�鈹=k�o�
'^V���w'{�*���!Χ;�t�Sۮ�Ñ."�rӉ˄|>������Upr-�Ҝ��~��vԖ4�Uʫ-\o����
��\y	�����1�Z��U��kE�ƶ�,c��U!�R/1���̳�!)�,�/�ǹY������#r�VlGӯ�������{�H��U~ʗÝ�j�C1#0#�G��;��|����2�.����S#�njz^g��^��=��1�e��
Q����f��X���{u�M����K��}�E!7��>���+���Ҝ�,�0ڛuʶ���S�a�p3�na�	a�EFV��F�J�M�Pg�*HR:C>	���mM9{2�h�s�f������o)��!) ��[u`�K���Gl�]6c��ڦ���Ep�C$�H��SZE14% �%�r��Ƅ9�]��4	]��3���8���҄�*��v�*;e#+�}��/�LW���B��k]��
�{�`6�������JȪ�S���;�듎�����ERKꔖ�ɝ��2}��9�Fo��ԧFp�֟���c뻙�5B�^�~�c琏O�AJ�?�ʓ�y�.
�?ZV1盈�o\�x/���ī�(��U�Jf)Oo$=æ�׷��ܺs/��{�R>�d5Z����Fr�0gزa}1 �"\��(�����s�(�>:o�T�*:�ۍ�<�q�c]D�p��tR|7t��� yO��3'�-҆U�R����%����6�뺘@U���XϱZ��˿M��}U<}Y�$�8�{�/q�C��z��ub���h��5�L�%sݗ��9�|<_9� �N����G��E��a`�Rq��n��� �� ��8:�޾0�فv�2�%Y]*���g\��DZ�5���Wt]j����rm.��3{f��PL��S"dDL���v�0�UO��v{�әg��}�Foؾҍ�G�EG]�Ib�o4������� ��i�B��Y�^��*�Ut+�_�:^�91U��y�Y3�A�4�h��~�3`���	[$�ۻ�zu@�����;]�m"�����Dkι���o�*��V�+����<~�nY�̾�yzd��w�S)+���t�H%/�5RG�=�k芫o�ާ��USX�E���϶a�+�s2�-n�\A��39�]��}y�׽�z���{~�~8�W���*���G���鮈��? ��sAh� �{޺��r�� wŨ@� wncY�]ۗ�s�@�D�C��DN��bf9�;�i�І�P;����1�@1�� U��K)K�����w�	H| ����n�b��qd@�Q^�vc���@� �a@Z-U�$ g4�k��s�^����P9y�G��_��y��G����5u{lݢ�-��f�CC�]�Z{�qM�{�����V�s�(�|�~�P��N~]���������j������QCG/�g]��1}g<Q-�D���m'T�LG
���9(f�;ᙯ���91F��fI��P�z��pы*�;?`��$B� ިR� ��� }�^�=��;���f�j��x���5 9������9�pALU�����4Dm �!��@�t��w}u���9�o�@�U����R�����zիD�� �h.A]�h�����G9�.D��}|n�;Чs/6�e�| D��>@؈�AJ��fh� g4!ct����7���pS}�%�=�Z��5�5��������/Uh�Dj"pԙ�;�By���h!x"-�A �����3 �Y�:���' k�@����W�x�3~ T;�����8�Qq -�j��KqE���:���&�@���K�N�΅{���S� �~p�_I�\�W�4�'���oޓ;�y�HSlB�ݲ�*��5���͛��4��i���Ye�r�]�)��и��\Z�i���iU���(�Qk�nu ͖h�P(�-(.�J�m�\rb٦�^�+F�5 F����JX�A͌3s�ͺU&�Ͽ;��fT)-��[4\֙暷5�.E���Z��B�AĈ�� wb��!{���s:����Y�*)��G}u�뚓�7�QuJq �)(1-!��"K^�|��Ίئ"��� �s�oY�|�V�h����DN���P��U�| �(�;�o4��1Jf)h�`�I9�u�U�^w�[c���^��:�� ������ষH����hM���D��������#�&���q(9}�=���k9�D��m3޵n�}�Nt�LGp
 �x�*
B!�DLb�-�C����|�~ %y��߽N3� %/�H^GP����� f b��X�g���BS* L �(����bR6ZL�%H��u��:JI��N�Z�lAHЁ��h�� Z��;�Z���ۀ�6�u�N�/�-�D�t u@���mA�"�#Q���yD�AO�(���s��J����|T��Ύ�:�u�ɩ�mV����/}k��J������9 �;�"�q���3���3��<�"$ w@و��u�]@-�cS|���D��� ��@�E���x�օ����Y�:�W�h�DI��#f*N��@�G�1@�DNw�;�Nﰠ<6�%$�<�����_�sV��r"H�"5&�c�.:���q*)�RsAx� �wlj�(��4�y����	���Y������* ��u�h)7B"`�1H�q�s�ќ���^�ޭ.j�a����n��AΈڭk��#P;��	��k� b Wٻ��S���	K����V��ŀT-��7�$D�3(�b���@�"cS��ԫa0^�-@����g�3{�j� ���!��,�IF��,@q���j;�&bf Q7�DI �'%D��% �
�hw���;w����[wi}��V}�v��i�ê����5�Ҳ�/F5�'x�v,���f�w{�}��'ĒI!E��������� ~"$]�mҁ��$��P����[��]�wH=ua��x��ֹ������N'�TPDy/�]�~��hQ�8DA1��lALDJ��ջ�;�<��w������w3��G��������p0@s�#���=�y�'�3�CSR�@���"�T��GT.�8��QfΛ?zI�i �ȉP%G�L怼����O;�5��g�x�P8��k}�j��9*#�����S��w`���q ���� ��"j W-�����sc\@�R��"$�(����n��1��q��_4�$1H�Dq ���������k=�7�;�V��Z#�"�]R���"b �ȉ�u�g����|�� �F�D��;�.A�P�@��~��]��3�@
�<@�� ��Vz"�xv��}����u<�u&h�]���ј	��lӾ���m�����y�g����s���#J���"x��Q[A<j�.@�� 
�>�u{`Һ����.��k��)VNnBow�<��({� L��D���u5MH�,���"���K_a�F��N箧����m���~���*�)�G��̺�j����穏}[ڐ�[��īMjW\�.��m�<���{:�#LϪF��Q2[q��3{����X���� ��<�_1�B�i:|��m �73[���1�����?�~�| H}��(�4�:����0�؁_��Ki�+xU��[�(�r�$3�p�7���`�#�y�ҬW��Ρ�2+ч4_o�M�+8Ñfሑ"ۛ���m�Y��//)�������e��zNue��;��h7������#�uE ��9�G�N)w��P����D輝�:�0������-T�j�y��]��39�ugcm�d"�f��Y�d4���xY�.����#]��Hf��-�.K�;ܶ�q� �yr�Ҵd�l���2��+un�'N�2w)��غ�GL߳�mfm�Rݕ��:��W��P�RtѺ�)]���WXa��Nȗnʬ����cZ��X{g7�c+�as�����B�%���]��Av$��s�b)��v[�7o���ƍ��,��y�\[pÁ]N��WC�O*�z����M���nV>fdZ�R�P��F�Y^(�JN�b�S�[֢SR*0��m�ˢ�3J�@�Ǟ�0sby	�	b���&iK܇����V��
�<�I"�~��nv 郩��1L؃�b%s3&L-I/>���ͺ-�)AI��XRЇ'�^=���rZ=�wu%r�ڲ1������ۨ��I2J�����Q������6�P����Ki`�Բ�v�ד��Ԓ�V��ݶu3ę����ZK����`&9h�{��u�$ذmB�h����vZ6`ږ$��{��5��%!F�Uh���m��;re�%َF-� ����wZ�S�}]��D�q	P��-�mf�X�9�겊��܏����߳��!ơM`m�[ފ��BR7��	.c�Z�q)ii�����-,����"F�X���p�B�&���Z1��4[�K�L1��5��#{?���	囓A@��f��&�q��G1�u��R�db.�ZG:2�`�(�ur��F-��+����d��E�Z��Khe%S&ļ��������	0W;��F�#E��Qf��
3l�]K@-45�(a%u�Ga������A�P�M+1���KSA*F4�-
��z;��b���V�DI�!v�Mf���@.R�#�n�ĉ��t�e��9u�r�ݖ�$٤"����&��F�in���M�a巴��3&3]�u[�hU�(ĉ,H�,h�K�U �Y�b\�il!rf�U�$i��2��t	5:�lՌ&"�M��]4�L��ң,S2��T�V�i�.�3�r����7CF:i���yMp=K\��뀴X��Z�)���	�h9c�l"5q5H�׀�P�%�ۈŁ*�\�56�Y�k���Q��RX�Z�ьs�&6�]�/jH�)Y�<�5���n�[(. #
���i��m̵XW6�hTF[-e]^�c������814��j�v��t\�s۶�.�m����]
�ET�37#rYPC�3����Z8nt��a��ԭ1Lݮ�]Z��'��$� I�H(T^�V�r).�D�Iw�f,/Gbۡ6�E�S[�(h�fZK���Mbm�kH�d�������Őب����limF�fյ5�Є�5J�+�F�V��ا\j�b���W8ōح�C],��p��i\;��fq{�����~�s(٥5ݘЂ�A��hŕY;�Ar�~���w�K��]�h���R�25���2;N�d)�C�g�Ž��Sϲ3��v2N�ǂy�]�F�	(n�Q��������UT�K헎[x��Ekf����� �d��q�����]�^�>��s����}��vn8NȗY,'Gvba��1$�RAH�Q-3ͷ#����M�2���Km#H>�׻��S	6���m��V5���m9�{�
�tΤ�f;+nC{�Ҟ�^k��"�����D���w�WV-�#"��+ �H)"+�_��r��u�w�����;�~,�� ���g�SE
����{������x�2+���3S�n�s(-�.�r�]��Y�x����r8�>����D�s���E{׵�z��t�������5A0���ϟ�U��\FP.�sL�K0��$)���Kh}��3)�Sͥ���7�D�:kEe�̃�uƣs�}O2)�=���=�]�9��t�IܜA"��'���^2�5L�J���ݣЋ왰����[+�T�}��"Q'�3�U�3Y�m�Z��� ȃ ��2

H ַ�u�������u��!#�
��U��ۨΏ�-���{О�x���v3�	��.�Eڋ)`9]��{v{�k�2fi�{��re��0���;��t%��Kv��լ*bD(�$ӮRd�C�����3�I��?!�z�ш]��Q���:Fe�V���b<T�f7F# &+gs*�Ue�=.���nu���hl�3�H���5��:�9Yy�o��#�q�;�vD:;=Y+K��TFۖ�����qu˞߾��4λ�:����P(P( ���$�,������fe�	~
�Jt/����]�B=���Ii�*��ޠx9AP�O�J
DD�!��ц3\m1w������(�s��_W���ѵPp��'�+L��П�O�ae���w8�;uVm��VD�Kד"�'��G���z꺛�x|ȼ������5�;��wuN�fK��u�vxkU��s]��B�g�UW��5(]�o����!�+�z:WZw��a(�-R�C��fU���];��igu�SU����TEٛ�k�%ZS{��!�(� ȫ"����**11L�B�Z�I�.!��]tjTf���X�s�X�4R[Jr+P�v`���\0�������34��)��m�Է\�8��K�Bf��+��k!)pkr��T��U˥�і��gh�g8����h�}�?l,��Ɋ���[R���_
 �����"g?�ɫ�:�-m��ַ���[�9��X9�����}^ܳ��:����e&����x�nI����{|�q;3!Vݲ�a`��"f�8��sM�a=��~�vΚ����d�׽v�%*=:���nY�9S7�~՗���<��=j:�U��v��a�.cfv}�c�_|'����͇��qy�)����	,]��_r�t�yt0]jW��y,�5@���lB^���1<�й��.���q�#/rw���-���X7�T<DRDBA@BADBDE ���7��^3�|��� ��̪y�y�nP�M��H̘���{�r�.؇��w\Y�t�r+�jK��{���<�FZ�oU�4ҙR~���c�d��gou۾���"�L�=6�߾���|����*�,��9����-Y���,l�S)��~WD�����[�۔xұ:�4#�7;��EԼ�z�g�g1��y8��"f�P-�}�s�:~�PD��P#���0���̭&��%��«���ֺ�t�vԛ��qA�""��؅g8���3�d�����VEY	I	dA��{?7w��'�(�.�j�4mr���x!�r.�{b��a��3���!�R��_��O8��l��{��b;�t�/������n����˕*4ѺǴ.֙NhY��RV4���}�}��T9]>�vﬥ�T�a��_Qu"��������-�F'7�\�)�����O_���1�1LЁ�32���伍�k0���L�W\ ����[b�B�4��|�?0=��$nv�5vb#���A�PR�< R�ϵ��{u��=�Z�_��������wl`��*( �
� 2 2(�"/��`�L�o x��?7�{[�k?Tpփ�'য�� K0~�]̑yf J3&(����4�t����y����������})�R�W�spob����q*�Y�ߋ��뽿Y>�h&�����cB��k����(��yX泪;�31�ԫ�+�5��Χ1ǻ�r��iR{k����P��Is\D��ؽ�}��;�'}�ځQ��z"R�����H����)^�)vi'���j��Ъ�4m��uR����ҝ�Ar�(� # � + � + �$�:���/��"�X!-OKi���kM�h�kRܘ�#���t��B$ ��'-�N"���vD�]L8��Ȋ�u�]	��,%�����nnmA���$J�3I�Zm��c6�`X�qe��Z�ٕ6J��������#�����mU֌0i��D��0"$i�f@�Y�^��Dvv�Ę�Դ��Q�*=�46k�)%�s��x3���Wt�̑$L��7:�%�)�ys���UM8*�fWP0޶2s���Y�Аy��y�Cs I*��t}+�r&c/��8�'����������~��g���#b��5�
����Vvf��v����x������j��������Yp�v��o�F:"O>��it2��Jy�M&f�����\�Z���ԭ��;���^��>���		 II	BG� /��|�;鷗ߪ���k@?����2��&T�86�E�e�{�f̋#MR+i,{�OoD�Ԧjr9�umu����il��Mk��̰���.]�s�~Jt�k\GR�À�%S�g��BH��&�1�5�֨\�ftKb�jH����k���5��i���'�Sb�u�w���s�Qݰ�k���g��2-;HU!_��ߤ}� ���߇�J+�'eT�I���#&ln��
���0T�%�۳�eه v��q���.�o	�X����yt��*�,�wxu�a��W�W֩����h�Z��Xy�����?�b��8#��w�θ�Ki�e��ms��g�Ͷr�I�����x0��N��g��>1�#o���5�iq�LcDS�;Dm#�aRp�eM[`ѩ��x��ULBEnUl@���Q�E��b[�B���<[Z��a��9�,6�o+"q,P�<-�e@hW_<vp;ܫX3Inc'��ܫ�S�*�ki�	�4���=��D�#�m*�Nc}���E���^
�Ԓ{����}���Vk_��ul�-]hl�u4��'/�gwEdn	6�d���j-��7!�$ڈ6�&Jf��\��J�ssD h��-�n�nְ��Ŗy>[)n?�t}����RP�����"& U�JJX5�v`�Ϙ����(�$�Ir0c\������jy��x#)HK�.\�)l��-ے;Ϗ��ެ���,*ؗ�Gm��([�6�I�
B˥��]�r�-�YQ3��wmY$T���$�Y�[%N�\[q�����,/�<mwT�n����>z�ש�Y�:���V�2�cH"���↹��,PH)�d���������oXX�㘪d,��"�2_l���ݜ����E`#L��	,��w;�P�*v2�"Y X���alU��7�m��Q# �#'o's�B^��7%�(��A��{�R��u!)`�A�HH�wy��;4D�S�����_66��,ck{%���F�Ӡ:����9ף�)�e��6E$��Bt�ː<Fy
�k%$�m�y�攍mj�i-�W:�Fie
�XD�P�����֪��Rb�J���"� 	 ���2
Ȩ�u�﮳ߣ�/C���X�)�眾Ζ!�	��������4"��NK�u���)$l�Ӈ�Ō�y�����p���ϩRV�Ѯ�vY'.��f���s�v+lȚ�*WH� zf$�ɷ���L����g;�ލ�R���Y����P@�1��w�����[���zO'7=DM\
�x���3�t��{�մ���D���1�f�GF��yQ��%�����r�w<i:|�'=���;V#k��������WZ�1m^�j�*h�[yּ("�"�"�""� �"�����׎cf���H���u�X|���x����x3f�����y��ߵT�M5�inڣZ�2��J�c5ک�|����=�r�����ݷ(ouJ3X�~�j�����/�����gUoO���Ύd��^7
�"W�j�=����>����s��{羊�*�>�/K���������y�M�u��ưh��(�G+ا�U^���L�!��wq�嶺��$ə�P�����ܫ��a�k���1��P��K@X�l�1�:�ӧB��g8r���%�|aZ��W��_�@�RDd�VE���ǜj�ꥥ�kvL�#A��4��M�Z�3p*70�.qiT���#n�!�k����j-�6��U)-6MB�@P��X�f��3���t� 4n�+C�XZ�R�[^q*U��2�V�X"��­t���~��S�O�ٻ3AЖ:.q�Z<#-َ�ٟ�w�y���w��>�gK�9��k3�?6��u
��ɘ��E�nF�M�lܾ����-�� �f�`�8�Y��?,�̛�`��"��FG^&���bH���ݞ�9��̫�iF�p�����}�������m�a<ϛ�D2/_�6�o�P: �0YWu�f���&�a�j���5k��̉sV�:gzg�$tpN�2�U�铚s,A�)���SU�!f�
�n��?�ͽq���A�Ga�u��[4f�c�z  �FEEY 		dk^19��=k����'�d32���3���5SJ>����|�g��M���@7ۦ�r������,�葿�jA��[��n�wc�"'�pq�5 ��$�Ȇ��ι�}��n����}��{�;�������RV¦�ŭfh�Hin]͙}��:~	Y���������5�[ӏ���K�c@wxH��[�:6k=�g\�|9�,�e��	ޟ�AY��b�3�~+�³��V'�t7a���P�u6�P���|��&����;�I矡U��E
 ��H� ��s���V�I�&z>�V��[T����aT<���ƪ�r�װ���,7��Bϰ�"eIfVf�y��z2��:gzg�����Gz�~>~���h��.�4R^3��/ �jZ�Cfgg��c��`���^��l]�|^C�-�Ց�3.��+6*�����=�����l��zP�	�i�4�e��v��bž�7�U�{J�Ġ���B@�Qnj�\��Y<7��dEO`#̟e�՚'p�mh:�\ݚX^��[�U�b�����of�s�����@BDY		d$A�\m�#-
��<w�*�P���{o+�]�;�h�d\�ob���0��	L���f�1v+of8F�]�����}���Fb.�z��t�tX��*g�{ު��|�Y���A{�ݟ����F����64���Pe &s�*cj5��e<'�#n&}
�,�fe���)[5�^�Ι�qI�1˯F��Xn����ڒ�OM�욲_a�^5�H�r^qk�LX��؞�f��O�CI�gk=�C�tܢn���]U��� ���*H H"H	JAU|8��m�,̼�f]��P�����3XԦ�����ôk�k[���
 �lFcm�D4���\� �AH���M�jdvl`��pM,ۉ�[e.�LH*m֐�B�H⻮�Ŧ	�l����]�Sae��nX�(,0�[K�.�v�Tέ��0a6N`�#��f{�}��/@5	r��=�S̪+�)gF�>s:�?r�ft�sZgc��S��jdP�����ja��n���{�ɘ���	:�;����"%⭽y��O
r�i�t�tNV�#<���3x��L���ͯL�L���$L��̞�;���t��31$���/e֩���#-َ�ٙ�
�2�[�ם��5d�(���Sʫf<s��㱻¬@�55�.s%@�\��s'>æՕ��,�C���YW>���e��5эڱ^|@AEYI		B����5�k0����,8�8�b0��8�B�]c݌��nw��g\Ľ�'�~���� �P����'�_�6���{����>�W��;9���{;';	���p�_o�~�?�?�_Q�����IA5�.hcch�����$���f�k�w�Bw��T�2���GCN�&Om2�;1�vM�<(���[�#����dę�2�bj"�8n�b�nkdG���@�	�k'oK}za �ٗ7mg,z�Z��߭[=�x�+�2(ȠH�HH�H�H�ֻǎ���}xԞ:��X>�CcyR�H�2b۽4��O��3zg���0������UU9p �)���u웲x|�� Mv@�)��?=��1D�&+Ih�ٚ:�(�3fbP��kW�(	�Y{��9�ep�
����J��4�s�Z[�?!Д���������kFL)�9������Z��$�m��{�WLoI��+5,�X#\C��.fe�V��Nv�}�u��u:6L����$�*��M|\�5�-Jy�vpER�P��{t�n���}����� ��2"ȂH�"�n�=�o�݋?\ȥ�7��Ǻ�_L�L�wt�ߍd�	w_��E�f#* �2 LIL����Alp�Cfgg��;�$q�r�7_�y9d���]�&A�e�3qV��_e�_g_Nv��b�Y���i�UM����[�}{3���ܾڪ���^JE�]^0��۾�����7'��p0��),���l,e���k���'�eҒ&Á��
��.����ʸ������Y��+D!mX>�׳F�-�>ѯw�PCA��H�?�����ݼ�������1-�N��Ad^�2,E�k�y����7�6c]8;��֭3��"6�FR��Θ�\D��,�Y��I�t�L�I��{�;1ӷ����Y�;A�H���]�o�ɰ�,�G �qW9�U��P�=�e.�6yf��d�L�'�fd��HЋ�nN�Z�;��c����go0N�Sк��֩bt-�}z+{b7�C����*�@Of>���;$����d�}���h���`UaY�6k��{A*n9/,�hA�h�t�R��ӮÆѡ����n�����ת7Q�i�)>�s��(gZ\6[�=�+���t�CR�M��$�9��:��F�6tH|.�h���y�33Y|'uu��u��Y_hU+֣�(*�#&^���8;ڻ��fjn*��K���͵\F�S>x�!5��U��P���)v�y磽W�� �H�Բ7��|Wf�~�z��4�$?ii(���`�AX�WBˬƁk���ڸ[ѱ[������W��cˁ��S���fkd�:A�SHT�ÍB0J�{��׿=o!t�Y�۽.�IS��X��|����Q���j�Ë���~z��X=lK�k��J�f\g�����O&!��h,Fw�owz��aH�j��a�oU��i�Z,�n,ԇ�=���gK�6�&�ۆ�^1�awE�^R-�iO��b���m�s֫}���k�����v\���p��c��bKK@ËKw���n��[�6[p]�̍��n�BѧfŽK6�C���Bb3���w��D�l�1c"S�-i�H� �k�AV�bD�ƪ�q�E�b�������%�/6K�JvX�)eK-��%?<��!��C¢eu��Z�!-����r�3j�l��ЅҰ�)���l���4�f`\C$GF]�7D)�VX��{1�0ݓ�F�èm�(Rk*��%�;vf� ,bj����f�.E�4�ų)�l��lv�%̬��j�-u�!�lR[.����g+SK.�ґm��E�`�1�� ƭԢr�u�u�`]��7J� �x��\�)�an���s^�ȸ%�A�4������5�K
��8*F��հ��l�7�5	�+��`6��Ʌ�hnl[���)*��)�nl\j�/f�{F$n�v�)Y��p�䴅��|_��z��C-Jػ�	�s]	���\��Dv[f���`�,��*�j�v�1ڮ�;�!c�5+c�q�f��C�K.I�lK��8�ڌ�*�ť%��Ja�F���hMa]\�VS;��s�����)M�^cK*1�M3$"�f��+�8Ek6+3A��"��V��`�Q-6P8�ݶp�rШ[��9�û:9lp���M5V�7���8�-���B��X:�3�͞#ԙ��yxU
]��Wa!�j�Q��T�VSj�*��Ƣ������U�UU]�V]nĺٶ]���!�6�\T6}���pD			Id@$Tj��xK��ɫ.��5
n�MCp3��^X%�,�@&5�̅Ж5F�J*��S�]���X���9��a.�b���s�s��Wf1�k�Zk�4�-m��Bۣ)��*X.�b���Gi��Ƭ�Q�m��?o���J�1CE��ر�1±Z�~�y=y����{��N��L�7��G5H]!Fq����U��Yu��}�x�ff��u�P��}�[b��^�v8t�3��k��ó_^�����k�}��)��)�^���4�ߜ�E��ڽ��|��r���ٝ��r���������k��x̦,�&p�ih�EL	�)BS'�j�@�눾�W��a=���:���3�r/�"�ϥE��2bb�j��h}=�d�V������y�Sl�ۋb���Wj<غ��Q�>� |`$��"H) �(=gǇ��_��/m~���:й?P��������k�K�����'���eT	�L�"��x��'��B5x��-�$���2������T��td���]��}�_:B_����{���3����������[\�PXM��n�v��>χO=\����-� ���s�i����M5E���p>��Z���b^��/HG���i����zɚ�c�mT?_M���:���r��zV]6�
�~4��17��otys�}����;<�7�Ҋ�B���$�$A�@��{�}�V��&�>Pd��+��1,���7k�Hޛ�}�Ns	���e^�gJ�j+��(�Y[�>��5�Y3��}]��3���L�dE�\7ϟ,�}�xO�-��TwX&��H.6��&�����g��~c.N�܎����U����~�T��$�x�W����׵��<�0����+�Gn�C�Zj�&ga�:Ȅ�����=���A�X�hM�ՙA���{��L�y��E۾��Rޗ�uf�b,/�+EL�.�4a-�8�|n]�yQ�W��Hw�Űx�	d $@�@�RAWX/��^k��|W|��z����"��>�yX�23�ޫ��#��j����V�d����m���!@��&f%�5�G\	0*rj��Vd��:����x蚥�bBM��y=�^�ۙ�����U!Fc�g��[{��畈��3+�"bi��360���(#��b{���%��������d
4D��P|�:��'�8��2����wtw�8���)^�#/��6ܰIK�:f����v8���6���E�V��1*�¾"�� H�"��gt�wI���,��Z�J:��0�e�m)�2k�su��D��D1���WCK�ݰC�L�$�E��.�7l�hX��2Z�jФ
�4��L�1��]�Z҆yG0�,!�%-�Dn�Z�*Ua.������ɡs�mY���x����/��cn5r����\���{���Q=�[��M�����Y����۰}�խ���O�2~�<�.9�x{����$L��*��`�|�<��N�$����L�I�KZ~�)�U�t���x?,�^q���Gɪ,�,]kn[ܼ�kyI�����<?7��<'��'�{h��LUD��˪4Z`�Lݶ6*�ϝ�O��k���-�)���tt���C��hW�m��f����ݜ3M�L@^��\�ѻLtq�\عVѳ��8m��]��:�^� ��DdVAdBA	{;�{�*s��O=�G�hdKU*vb�&>���2QM_;��{��$�������f�p�P�8����������9s�]=��?)�E���Ni:��� ���y���\"}~��b�A<���}{�x}�5�a�+)�*���L��]m֯�I����#P@�ݡ2�m�S�̚��7\ga�:怹_\c�b�	���p��I1C�Q�*"����r�;���<D�}�{V��'�`i|�ʪ>~�Hz�7�솺*Dѿ�h�͉f�K*�	�*.�@M-��5��ȭȨ׿��x�	"2 H� 
��:޺��痓	~ 2�8�B�@Y�-|�l�����(� h�T�j����2�(� �5�^so�w��u����1�$rx��:qt;�뮍G� ������ۮ��D��^��L�&DH�KmsE*�l�ɥ�1�?�&�:D�+�%�_Z�k[�{��	{�w"��M6T��~�j��'j���-z�f|�P��WY������/[�mO6Ý��=�+=�h�bq��t�ˮw{uѢ{�0� '��N�5�Bw��DL�����=����{r�a. ���]�-By�ʃ^5��n6읿W�z�uxW{�o��K�s���o&�w���P��h�Z�R� �{���br|�5HQ�F�]5�o�A��N������8O�/̤|�,NJ��O����G翫>)�kG[]�֒���0�r+.t��=�����!,<�
�E'�ۿ]z4I�`1܊�聢9+Z������'=��%��w����G��g�7�MV�
�BEe��W �Db��oP��0ER���5����w��>�?1<�-9%<�<��a�_D�P|��( n�I�ߒ�������Vs��}:�2a��<.6�r�'��D�W�����.�R�A,�AY�PA+���&�=\�r��i�v�-ݴe�v��5�9�L�.�F�7U��zy<�����b`�L���B��R��Z�)@��泂&�dɊ��VcZ�4a�]s�8Y�u�eX�9�qkvJ7�0	b�T�p;;:�F���MU�!a�k	��^vέc��Y��5и3,IK-0EVV�"F0ډr�n�Z��ZM4hYST��Ω����r�=���>�YZ�^��2.Ա�Xit�b�L�y>���ؐ�ف��Z���N��o���.� ���&��9N���������ۮ����Ψ�D\�{n�U��<�y!��ϴ=ٶ��bu:6�� q�C���o�Ɵ�s�o0�a�C��]X�� �e�db��mA���;��+�k=��^]���y�-v!�%OЎ�� ��M�wfe���\���y�ݺ����� ��~��;uhv���=hd���nm�EС���ne�w���|w�RS�u�۰�@Ԃ32��O^]̤(�LU�.?I�X#�YW� A�Bz�通Ț艴
�*�-Ṷ�pB�ۧ7q�woM���9�!�jD��T�1�FԨ���� �I�Y�Y�\��3*�"}w���yt/��#q}DZ,�fv�"*��	6���/��o�n�939={�}N�D������Q��h
�;ޟ��g"n �HV��mv��yw2�@��uа[Q���(;��m��i$��P\Pю�.��/���.@�(��$N�p�C��Q�"M{�ƙI)��K��+Q�8:fݱqV�x�C��<�����������,`�v6�F��|)��|�,�G�ktWC�F ���)����z��e.Zd��#���SQy|l�_�@w����P�%@�A���ϯ=�䅥owqMɕvf\yI~���n���C(���b{j�]/E�AۋV��p�z��A�wU�ZU뼨X��S��ز�d���Z��y{�Y��PG���:J�+�.���I��� z��,V���4"�;[1��vT=��˱��Վmi.fꩂ`'��;Y�y|�#w[)a>T����e엁=,<ɳ&�� ������8&®�A�����k���-�ņ�����m���R��N[gpcw�uE���"�s��+�9��Vʡ��⚡d,z�ٹv�2��?��t:/ab��fv,������^�Ua���\H�����L�:�1��
�&�#�,g�+V�hRX΀]�]>�ve2�,j
����;����'�ɗ���ӂ�d�]�ڬ�̨3���w�.�ڥ��T��Y��'�@��]\��i�7�%I�*�N>�(��V��+�e�B����v�ɖ��o2�,�]�����~�EEZWv�Zd��,b4ң��DV�/��y������F1���УQ���H�!�7��8�M�FT�1X�0d$R��Q$�D�CswuD�H�� �QQ�o�M�b�iDRH�L���֒I��D��mԩ�D�"���`�
���B^���l�n��!!$���im��4�/6�u�D�I �r+J��F�-,-��!)�-",����0��I"�$$E�"� ���"E�pR�ƕ�-D%B�w����0bDX�F$H4�I"�9#j�e�I$!�$�F ҋ!JF�(�H,c���*��(Q�I $A���x�:�l��u�A ���E����8lM��b��(�V�@ݯ��fE��^vZ� �@��y�ooׇA�)7�X���u����U>��>ϵN�ϧ�.�R��'��d,�fg���Z�����Bɥ^v��*�f�{GgP]M���#�3U��y+��X�o\�q�\ǱE�H=4�h� ���/��!v��	��+�̈u�,��8G�cӷ���e�����ʻ����)��5���^������n�8�d��0D� �8��OsϏK�;��M	Y����P�s����Ve�Dp,���'j�nÇ�e��Ѯ�ꮊ��tnl���4P����ru���q5m�o�x�"! ,�"H��d~����A4Q~�]/�X���@����w=�쵢9}�$�?Y�T�V��u��{�מ�Ol�E�2�,Z�٘����Kvc�6l?l�y��BxADDv��}=yw9QF��}Y�0�(k?X_�Ѡ-��V���Bm�_���\��꼺�Qm�&���fF�a2�>k�Q6݂���752��5���;-h����A?U"��p��,�
���8��U3F�}ޮ���HQ���r���W�r�	��������-ד.H!8��^��ƨ��xV�T���Y]6�6�����On�������V⹐���{��s3�����9���{,�(�JR��(�Z�[���� �����ݚck��p.V8�5�e���ZU�7�*:��f�6�,ڇ*�s6�v�L��:1�j�ku��**�Ea^��:�K����ѡmb+QQ��%Y���&K�B҆ms2]q1��2쟯��JK�ck,^&���ȹ���i�6|�o�e��K<������;1h��w�s���^��$���?U!����?�ʵ�Uv�;a�)}�,���}U�w�����#PØ�`�I䍯� �!_Q�T#���os��:��� ��?m��(�� ��9+��i�ex��A�R��E�o3���A{�-'��m�r��Ͳ�!�1����FT_���~�����>>�|�������_{�Zp�o�F9x�&n����R���a�+�^fS�@\5b���4�x���yMj��f�����k�#�)/��9]�d՟�y����9zj"��{4g\jE�C#5��c3lP��e��b8��'/������«�)JQiUV�|?yA��+�؛�ߞ_�Ţ9��|F�;s9�����r��OO[�l��R��doj�����yw2��{�� �u�ɲs�e�y�"i�A�g0鸪��gVm�\�e"MNqc�($%&�9�"ry���{6�{�}��r�b��}�B:�F���G������X|�2�-��J�]
y����:�f.ϩ���O	4޷}?<���Me�8�컉K�
vc�4AjH6��El܃(nP��R[ӣ~���<rk9��Vm�Dx�������r�\�ߒ��u,�Gv]"��o�o�ٓ�c�ffgr�?dhU���ٷ	AcD�m���G�Ͼ8���8~~�Р���'�@{����+ՋB��9�8h�D�Gj	*&2���� ����#�������%.:QƠ��/m�d�WH>��j�5Hj�0\iC�ޠ�@�]5��άۡ0���n! ��L|q3��篋����.�S)ԙIx����@��ظ����^���	j��f�ub�"����-�+ʸ"v����7ek����v��6W٨.���]��u�M���&�	ˈ�)O�S��!Ђ.Ѐ�G��B.�XSYY���Y�Bc�@ ��?n@��4Cf�Q�[�#6��4C�H`7
Z�}�*{��/���DԨ�lX���p�|8��N��rۣ��b[�;c7��b����p�q�S$^�ˉ�?IQiiW����0G���M��`ӻ�Wr*:����/������e�JBOk��6>[���*��0(�
&-�˨b�G�K2]�L��R��X\'�
"s`A�3q7��:�n�������\��\}�����8�&~B=촖�Bo�ts��������E{����<�6�ۓ� Y���X�b\�_Z�E53߹��%��cG�z5xO�-?A^�&l|f��+��<GB��E�n.�\g�6�Lu���mJ�-L�u±��`3T���;A����f�F�]s�Ȯáw�FrAy�"���c��)��N8�*�JV�WV���3�f�,o2��;+s4��7��%ݬ�2�5�����U�U����Sq�CӨ�h*�]����L����:ݠ��a��)�G�-�Y�V&qQ��Fՙ�����qh��e�1�8�&�\�b�M��r�)�Ѭ�X*�A6��!@V8�rܓHu�U��P�%.�e�]����÷�k-Qb�CX-�r�*���f6���\~_��o����2�W���{o�����%.ltʹ�P �'�&�AB�#}��g3��?���/��=�W~���g�*Ow�_ÈЗRg�Րm}v����0D]z��q]�B?SC�/#�2E�["@��"*n�-�'��4�����gv���쪉��?�Jܞ�F�*�vNCy��������f���!g�)��X��>�wyt"�� ޘ�Q��A�mp�h�ӂ&�e��~cb�$1Y���ذ*�u6+����O�[����o�g�s:����5�:!���	k罈�^�"n�bn݈���o�g�e�w���r����q����eNٺ�m�^õ�""��D�T�E;���:�	�Oē�?G�dc'����:{o��uvUD��k� �Wk&�LN����A������Ap x����W���Lu�>�k¤��iЄ�
�n���� �� ��b�u�ێ���\�� �z��A?f�"� e9���L��e}��Yn�w��UD��M�����˽ϼ���}�ɗ���˶��+,6��S/�'�>�@�-� ����uW��U����j�a���.�,��A� "�T(��Z�#=r��j��5t���hG�h��g�~@7�w!g�f!]�|E��иeŬr67�������˽�b��Y�s�9Nm������;����r��Yf��s��{�~��R��"H2$����]N���1k�xc���:�1G��PF �O��N�ѩF���A���N��_D��.����!q�53�uԎ춷e��;���!��9�J�����5�t.@�|�� �@�wgs!��}۷���&&P�A��hE�����E��!��G�q��e^���u<�������s�%��y+�����#��_�?jRA݁�n�D�f]	��H��� ��/�8V�ֻV E���?i}���Dz���3f��~���{�j�WI���/m���ӽ���.��ܻ��n&DV����*4�Ӿ�oQ���^4�HUe�K�/|��چvp�P���z��[��"_�	�~?��j�����K�]��G�ߵ�Vjn�շ�'�2�Lt����������D�������>gZQ	��1���e�q0]	C.��i�6��=���}���-�u�ێk��^��c!�>@^!�(�w�B c�T�r��*$?AJf����^��,���_@���UCT����P( N�A��X`������'���ՙt&C#��{�������q#um
��Ӄ���s_�v/A�Gˍz���WnQ�B ,�A�2��PA?V�3�f�cb<�׈<y[���M�����}���vmp�O0������{��ɚT彑u��Xw�e֥�wF�<Z�nd쑧�6s�hI�F����h�'�7�M�-���v{�p ��{�Ep��V��6�o7a��G$�de��CDuY����p;JK*��v�chK�P������2ru5��͘Z�V��U��d�Ja#����#��G��dٳh��S;��>�����Л�R5]O����k╲~u���������_v[�.-͐͡:V�ܙ�q�5Qy���}a#'�-N�S޽�=�4�������g5���ХIb�+s\�4�t����d�2��L�{��ݬ��n��G�6l� ꢜ���fH&���3��[J�5EA�݃�a�f��n���K�:�d�/qȜN�<��ɍ��pc���<�W�GV��@�G6%Ӟں��d��؁{2���x�m���u��юܵ{mN��CrS�?Q��u����h���&�]��Yi��j�����;xJža/	xk�2
	*$$�E��Y�ѱd�+%I����vRʐ�0�#UUFI$"��L�4��wEvH�R#q%ihY)$`B@owy�	F���KL�*6!.S �
BI|���%"����"+����A���0�\�ZP��^n�u���������IQTV��-�T.�w��쨋d�cH�.Ȫ2FIJ��Ԍ�F�{����Z�]�5r(H�,�n�B�cH��1�y��9$�6\XF��J��ڥ�^�KH��YB�`��޵�Ye��-�
Kci�\�$�-HA���K���_��`��TŹ�2�鵳R����)�R�	�vÍZ��AmG%[ac\��Du6m�t�!�����4.l��ٙ#��cpB�E�v����6�����lt�3�3ͨ$c�f�i�B�,�f��vXF-�Mt]���iԘZGR��g�v��,lҡm���:�%0��x�,�$�R:b`q�aa
,��Sgh5\6�*���l۵1]0��B���H�:��aLk�C������5��y�SWe9���4��� �
�-��2Fb�� 9IIvZJ9�Q�DҒ�h	t%Ђ�@E���\6(��l(��X�[�Y[{].�f��b���*Ĥ��u��Phj�&�;R��a��*#i��[h�+Yve� �@�6�4X\����q��fmH�XQF��ٰ`�mk�4�K-�qf��vҐ�&��4J�S�[c�L��t,��R�Ij�4`�1���#c)vR�����%1�"˙�1L�6ַd�.���A٦]v�DCA��MtKb39)sn��v.�4�j�\�j��MP5Uѥ�\��ռf�5�\��"�pU]��-j�8Zۣ��ei4
@6�����sA[��v�ML�{Q[����! �������MhlP��	m�i6��Cc>ɷ�,O@
]l��5kmPTѼ噚7M6Kmv-���Ph�3�1�L�ns��jc,۶`.�C8��I��&s51-3\���y�R��Ԅ���V����Gl�e���~͏��s�CA���!6���6�����{Ͽ�#�g�W�Mz�3_L��.��:�#A'�����M��u�n��6R������K�uF�f��s]�B"y_ !�6g8��D�[�	���,P˫aǢ7طj�ژ@S\A��7j?���s����{��P����h�ͼ�g�Ғ�Lp�OAё��r������"D/fG�r�0�v����b_��B\c�܎�á���9�����m�v�}��?+>~{�|as*��XJ5tR�h�ę��W���/��_D��\}d(��wU�ژ_2�dip �����Y����� ��>�(�=�B�2�&��ѽ����d^�{]q{fau�����q�Ѳ&v�!���H?H��O��~?��g�'�Wy߿]VeH���D���ʩ���>p�yA� ���O�v�J�l(���mv�����+�A�(Iuvi����g�n��i��K�����]�nmL/���U�f��@n���nЎA�+U��Ϩt�ȝ��WUfL���O9������vȃ�Zf�<'���5�2M,p��`(4@˩6�&���H�:�w�߲'1C�޾Վ��B����0�]�3*>������܈�`������(��G�j��ܻ��ژ_q�PA�7j�3��葥��� �́�]���Q�~
ÑeW]��w|�I��J�Q�S��=����]�tM��wWD��9�Wu���ĀL:��{��Y�"a<g��n���K��՘����̇��� �H"�@?]�j3�ڱ��Џ����Ӽ�>����وH9�+ x��oϘ��Zwr�׺������_@��ږ��J�魃�Wۤ�]$�"@�#�k�Ҽ�4m�[�.��3�&9 ��F�2N�e��=9�"c�}���`�]��Q6�ɟ�/��~7j��_���ّ�����F�o���u�й�F4 �Rh��%�#��(�.�A�W1��@7�����3�}����뿃0}!��*����2�"�,�t���n�w�zo"D�@'����Y�'�����+�]E�͔W�/w�{�m4sɆaڰ|�
^�}�,�K�ɪ�O���I �������a�A���|A��_��Y_�N �QN/m���šr�!p �@�7l��}�������qr���^d,&H�+SK��(�>��g�xu܁�-
�o;�O��qL/��S�1������}V&�?v-���v����=5�"c�}�Fd"����}?^��W�u��bdn�<Qm���tO6^7x�.�s��
 �@��ݟ��ӱР����7b �"[�|�չ�0���ծ�ȧ��嶾�<����������B�I�������q�Y2��>�IRj���Hxh[w�yxq��[
#+�6���F汪��`p�8պi��֜5��[�:4�te��Y�Kg��-
�%�_I���kkP��ĩ��� �	�`�٘�)�K	HC:��Rbd��ڴ#�a�l0H9#����,M����b�5)��].�+KX�,mJ�X�e�6��n&�mZ���]
miP���@��emխ��[�����ƖoC)�ײ�΋$dɘK�e�0|��4��i�GvA�v��1�����]Q��-����w�X���C�������}�ޛI����C��q���0��|������+4|�M%9�!h�n��ݳ������Q7���uZ�1�<��@���_YCg��2����B�?Fp|��j��o�Z!ŤA��Hbҁ�E�� p�À.�c�T���+�n��=�nq�n�� ������RA7kdfO���������_q[\�G�lX��A5��00!��>�e��G��1���2}=]��ܮ�R&8D;�GL1�(|���2�ٶr�͛5��έF`������zc4�&g�Y4^��ؘM�ͩ��j-R�kfAY�'��	�z~y�?n��Q�~k?vdh\'y���F�:�����@h^LYFNbDߤO�A�q�������R���o��5n�M��0�<�B<�rC(�3 D��^yٟU����K��#q}W�j@?]���ŵS����t�k��^eh\��Bc�"�b���7�ϡ�>�.eR	�Z5�b+�&#A�*���=?���d>�7`@�Q�s���R�q[�Ll��B������I��b:�ݜ�FPf��.�/9ٞ�P&8G�Q��BH�3�i�����r� ��x��1	"Nb��OL#C.B�Q݁��M��Wy��̧�qN�ݳ��S
��5�'%:���~?�=���F��"?�hP6d����B�#Z��G�t�#2#�"7�O����R��o� �	RB�=��a��M�R���亰�]�v��=�W.��y9�g�7Y}x"d"�P��;kwL�g/AT��f��,�X�)Df��K���/!����^9��,� ��7������g^V��n��:�!��3���i�e��������i�����ejM����*R��j����f$�{����,R�?^����0�.�mo#�=�H��f\=~Y����Y��_gnQ�V�wU�G�|�1`��Ǟ�έ��/����,�}��K�*cw.�=sh�����ڨ�~�y��NU�gk--ɪB�=��O��^�����fG���F. A�c0S���1��s���d�K�?o/���ŀ3^�d��Ϙ`�ߤv��2��4ܰ4m�[�ɕbfE�1�AP�ev�}3������P*OM�{��Ԁ�_Yn���ԟV�׫�0���O=쎬��@��A�5Ι;�u�ă��^��(|��M��5πڜ�W��tyxMT��i��v���r�|o� ����"�}1ۗ~c#��I�C����ѹ$Vq����\j;�e�?[?6T��f����.�;�:��.�{�\}��ݺ}~�����1z4�� 	"TŒ�<*���S�;$�G�eR�.����ݾf��=���}�w�10G��Q]����԰�%0Uv����5��J���M��Ea��7�VU̷41�8YX��e6y�T� �m��̵+34��h.n@���H�k�v4��Z���rXjY�K2L��rYXPƷv�%p��ù�g7ϟv���fu��L�Й �;%�M��>�#���(�+ AqY�Fu޾��˘���3/�y|����Rzמ�Eݖ\5-݅�Z�MeX�G��"2���������n@�C1KX���d?,�$�r� �6j��f���Y��B);1N�Q�#���w>y ���E¦p���(�-}�/K��GK�����hR�"(@9��j1#��Ц��2ԍ6)#�R��&�;���>���eǌ����2{S�؍�ޑ8y(�J)\�(дj˶.f��#�
��@J��qt�;�T�����{���)7a2�X�����J���W�;+eU�Q(�5?\����.�1��;���n�>q{)���$�O���$��� o/�G������빁)q��#v��XQ�T¨6)?HjѣN�0hz��zj�������Y��� ��t 2�i���̅���A��� �7�@�ݮ���V^�I�BAb��Ls����K��u�

��7��k���9�n��e.�� �#v��n׻wˣ���K�x�ŷj��e%�Ō�(��-���_%��}�f�=|�����M�wS�9t��c��/�������v�.��ȗیq�_A�U]���p�/�	�@f�@ߐ�i"=��C�Ü	��B�ݻag�U =�y1�:�����߄�B�S��-T����EfQU{�:�[�m�F��>*f�	�X�_{�䈈Ւ%V�pԎ[bv�h<�m���7�j�[�o-ʽ�2\o������ce&�)���+U6��J�׸9U�%l�wd�-���6�eb�4�'
ֱ��ж�q3�� �5��."��ֈKfQ�t��@�lC)w׸�Z�t+5;+�1S��Y�̵g;H���S�7�9�WK1f�����)�s/���;K��!N�M�megcڭ�jr+%�x"(8y���e�X�@��߰�KЗoq9��S����N�
�����pj��+���2�2��7�]�0a��D2��Yd,��z�WI�3�*/�&�іʚ�������;�u�ܭ|lk�C���k5�^�XU���1}/Jme�JAu��ҕ#C2d��hik;+kk~̓3���Z�d�kB���׆��A,�ϲ�ʷ~�s@���;����\N�L�R�
�M$;��u�[BR�y`�u��Q�����B5/y����n$�G[�ƒF�4�4�d�e#L��F�^n�T���ŦAXDRJ���E%�YH��/wy�����J,�2�K���T�R�!B�w%\%�����IF@dv����2A��\�e(�W���!$^n�ʑ���H����I��"�$�d���P��wu�5�1��IQ�Tbԩ ����)!)K�E�BQ/wy���e�,cHŹ�U�0�*#���!&���0���dd����,ZQF�iTUn���1U�PIv\�](հ�#ci�+�xC�[d�J�Y"��Ӫ(�;�ߛ�}���n�d��#�����we[�/0�Ry��B"�|p�QWp'&��b� R��Glw����$O�><��AݨA���Ӕ�ԋeG����Yx	�Bf��d��@m�Q�݃��*��Y��̳k�S.�Wf\�x�r˼��,_X���'{*�B}]oޏu]��]�#���c�D�_e��ڀA�@"�s�O]�� Ӂ*��sy�@%�Aˁ���H�,��_Q�PA��P�j��4n��f���^��{��l ٔ������^w�o�s|���^�yʿ�X��v���K�<�p��8B������3���s�r�Y;�:�� �F��ۙ�dm��S}�7������_���n��y��u��k��l��g�y���X���&�Y�-	"�#�h5X�T�=z={|o�}�>4�#�`��6a[ea��8���Oi߫�����t�(|f�/E���~Q�>�Gn^o���������u�#�e�n�`��^���4��"�;����Ws2�|~澍C�b�<�� ���ۨAfG�~��=9�����|�G^@��¸|j;�¤?Dh��8(S��CA��f)����V^��r�h�\��hf��m��-/��T��"�!���2*��[sW�<��fR�A<�Ѩ�$nןW�gz/!�9g�f�$1V��ᶇ�<DZ�Wn��V��7|�wG��y�A�y�Ҋ._�*ۈJ�$��v\�cqf`Ј���\�����2Y�tf��m��Fj[[�B˘�,B�1�FZ&�e�+4�(�\�ؽf���+��r+J�,{;M�(�*PcZ��;
ma�%�Ըg1���,�t��M��s�_��h.�6P+��Y��c;U��+=�(��z����^�mﺦy����t���9�R:�u�ka���C�͊�U�ۄQ���`��{�Ӽ��9G�~����k�/g����M���Yu�=�Ӭ݅���~�<-���(���}�M��̤k�����A�QHYH��@��An��(SwW��{�zK�%�P�E6�]�7�4�_ak��ځ�0�9����!��9��p�/�$��j�wQnq� v�ޟ�.��xE�p�-	�d,��ً��oϲ>��;�������z��U�L�G��>����~O���Eݕ�݁��+�u~��df�ŐI��k&��J�<��k���PH���Y��Y�&�GV������x�V�GM�[�}�WG̢2бM��;��f��(|>��~l����$����}�m{6��^Fr�BЀp��#1
ny�K8��@�C��$�h!Y7��O��&R��5�d1�cAv���A��9��2>�l׍��U`p�T���<3ِ%!ŕ�hAk�/��|~�~��Zf�V<�p�5�bPah��ظ����竉�6l|ٴ�N�(�H�k~��|�6����>8N!�n������
z��A	sY������Bz����,�Uə�;r���{�,u�&��w0t��&��EOe�`�Ӥ�S:�=�5�o&t�P���Ǽ�ˡ��W�}�'��d�̑)}��e��?f/�����H��5NW���ڪܟ_uì��'�#����4wP�7r:Q��4mXu}3�~���7�ӽwq2�O4=!�يA�����n9X|aY�R�D���%�3	���P1&l.�}؄s�A�8�d	���o%vd�K��3z����6 G�Bv#�A1G�3���澦���z�v�{�Q��@{ƪi�1t����];����ЧSj��×��aS���6��{+Ʒek�>N�g#���`�<�������琻3�*�∸�,��74��
�#ؘ�"��T"��V��v���	0�p�C�']�v�
rwy�y~����]]5�%\ݘ��������%����G�w�9Gƅx��>`A��p#��9�ٚ��"d��*T�rV]�V8G�].V.&�8� ��}㖾�A}�[���]�L��/�L�O��׳���Sݗ[)�bjAl�ЮJ�t0����I�oB}&VO���5ݺ��Cs��wƱ/&y1��C�(l}�������n}]�ӡ*�6�/?6��b̂��hn�,�g�,���Z
r�7ޗ�w) ����]m�,���7�����}g��mEu`b�dO�9[��Ļ2D�G��w ʏ���r>�����z�>���V.�u%��O��U�F �bQ7I�`�3��0�DY�*!%5�/Qn��D��wQ�j�9Z�c�Ը�&�ѧj�7X:�l�VM$L���iLVYn�q��7gZ�m�F�]�*lZ,"�b�f�c����`��t��c5�sV$*c��ݕ�4kU�*l,.���O����u�ܸ�SPm��[����g}���.�}�����UIl^��(��at/�5_!������}�֣�)F�"ȭ��M����~��wd� �{��D�v���{���P�@����Um��}��v����ٮ|qve	\#�~Yp ���>"�H~Wj��a�A�5��ͥ��~���8D���_�`��<�X��]k[���qS�e�0ѓV｝����@w���#v���Ҳ*F�����Yߔ�
a�(�Y�]�H�Fص�m2J���n��e��5W��qve}+� ]񩒀(���_E�d��0�pQ�a�`����sEx��W ��-e����h�iĩ2��']@�ϺU��>�~�zm)5���Q���5t΁��ͽ�ж�"|��(����d,C�J��q��뻙���A�B�<H;����]O<�9���!n�n�dT�x�.ˡ+��Qb�hn�'H�s"~;�<�@��5v�zG]�.ܶ���+0��	�B> ���A���#^Թ�����LJD�P$�T�-	�s3\�W�ذd��m}D_ѕ�ϣ���e.p28`=j�n,�5���MyAB7h�@51�V�>)�\�r{xC�5X}t�@���\��� �P~�P6�7j��n��Qf�dY�<o���l��7�3��j�r�SPD�K��j�7K1^`�q��w�9G�hxՊ6��/{�#�70=�U���?e8F���me��w]�̤5��xf6,�)i_
d��6j���Bl���Qg�f�>MVUС���w�6~L�nߢ_��~Jh2���c+I��L�c�H�L�AS>+�¾�<n��x�����r�����œW�]hh �p �ݲ�ݻ�>Ǟl�΅�W<���󻣝���\A#y#��s̡&'�+�Z~�B�;��� ��ˉʁ���g'��>���17n��en�hݕ�sX�͛���=���|h���j�Ւ�o��9��~�b]|�c��o2��[��5q��f�c*
�����_y�T̘ `"�7z>����Q�O�T�s��y��)}�>RAuA�!{���5;�{����Fhk]YD�̢ٶK�1�ۼ觯���!�u���g�׏u�]7BR
����V$0 ����}����-0���b�ZR��o����Dq�@@�Y���fhH��W@1^%Պ��z�ԭ]��O�ݎ�a.��}��;��'L����n�E�f/����:_�w^%�R%!��3[��ЪcH܏��4 ��j�߯(Ti��w�s���ŵ�����'��_�@����Rn��,���������zQ͛����Kr;j�슅]��v�:�2�o�PC-=S��x��L1ױ���<���X�j�`^_J%8��K{ibW]�wZ�%���@i��R��X(+�g��7٣�����M׽�'7��
OS�]��)*:W��p�z���}
賁Oo�v�o]��zٗ�Ƕ���\�$�ژ;Y7���U�+Ov>�� D��e�a��bF�)3��O[N�d�0��J��_۱ns	v>�t����{���L�Í\��Z�`+�����A*e���wIj���I�U��*W-��8=�@˱��C*J^S*��v^�5f�/Y�L�G�9�� ����T2��/��j�4ݢֺ�a�NUB�Q#wuۑ���)4�����5�4�ioI{�iG�/\� �����@�Rd�(o+���ј%�'ef�7ʞ�mu�o������=#[��"w�fMe�n���4�_,�o���>!�R�Jg%�g�.���\�>����� q>R:�9wm�x���	�e���Cۼy|�M�FHҾ� ���2�"Z(����EEc*FR��7�<H��DdD�$�-A��Д�RE���#���i�j䐒�wu�d�(Ҵ�,�5��!r6�ciC!$V����wtG�.Ј�-�	��Y�G6�m�R�H��,)iZ��,�r7y��V�xl%�J�X�%,Xc�sr����Z-��L�I2�������$�i4aI,�Di$�%�j�kn�%G�+Ld�Iy�ͤu��*��iԊ*�j,��\�R�P�m�(���4EiGd����6�ڊ�1B%�6�V�T\�n�U��"͹l��@�$��Eʀ�B4�"���ӂ�� �)��B�cl�\��%$!m�����_a�ĽMM���mҭ�
V�p\��l5KXZհl����1��^ڒ�Q�7)�E� �[Y�\k� q6 �x�KUU4�l��P���T��YQ��"$�����G;)M�8Ut���n!.��a�Cf0�3R�\=Anjk��Cim�e�`��Չ���]#� �%�]�D���Q�-)#�SfF�
�K7rR��Ύ�Иͩ���c��-)m�R\��Q]snR��P,�kk]A5qC4�a��!��:UՅ6��u�5͢d�%�--��� ����1��ٺft�%� װ�mt��yE.m&�"�uc4�5ڕv	j�sl�[e�H�	���9�.xU�[�;X��v��j&�Ce�1*V�B��MX�j��z�F4��*	*�ĩ�.6�bچ�CB��[J�V�� �w[�E&�Ґ�u���<�Dq �EK��c�,�5���̍�ƌh0ʃ�궍^��![*��Bi���7-�0���nR��.�Z�ƕc�^сF���f����KU��U��ͭ�^ҺUx�u�31��n�ᣬ����ĶgBn+�b��ܛl�;6�Bn��pʪ��kfP�K��2�r�V����|�V���g,�_.e�i����6jQt5t��K2�bh���1������+eleҺ�X�W[.�����VkK�E֥J�D%�f"jZ�I��X�[� v������v��0�
����a�fQb�eM���M��Ϛ_�r�F���3K6�g���(�\�\O�-��;��'�g�=��y���nn�a/$8]FfD��IZ֨ ���B�#9r\%,����z��Ľw"W((����6g+Xߴj�� �^�����'�k78Wpi����\�=�U8��Sf�5b7r9;'C� �~���AO�{;ގ���K�\"C{��i
&�D.�k�f���z7nȦ��n���.��)8
 �� ]����1�q�u��Y���41�����&�B1�I�Bby�j8~�\�*������5=Q�Ơ��`��M���r.,�2 p�<�u��.�g,9Q�4�9q�ZB�.H��6�ދY�k��@Ҫ֎ F���e_[�7u0�#y}!����V4�Pt�-z�
 ����n�"�E�&�tU�<K�r0���СQ�p�`��g�m�~�
5,� �A�SY�Wܩ�^��7�8�s,��(J6 �B����3*�ق'�AD��=��K�'yAUn�K�vm���ϳ�>S���c&,ʒ��vn��#`�A�n���1�AW�dn�FN�n�Ļ.D����
�ˇϏ�N��C���^UZ?	\��_I�P&���򮼼�%��j�`�����{���X4R��_�`�a����
\�<eCY��Z6�(��k]B��rXL����ר�����z��;��K���}� jɪl��c��kL֊_�`����c�ǉ_\�N(��L��<yҷ���������|��Ԡa����㔏���1�#ՙ+����w���HMV�M�:�\EґÄ�//�{勬>��vU�	}�^>莻����e��*=Aw=�D_W/�6o1�����sȐ!�(s����7^%���@'
#1w�w}n��Y��}fڂ��ڏ�&�	l���}n�*��5]y~�_w�����f�?ɼV>0ԡM���_�<��]�n�?o/���m�@�ǫv�mᨒ�c�(�k�~E�iJfO]]���g����L���J�����ˤ�P]�Z;���@��A7:gٽ�ő�"��ݙ ]���r�zֲY���bJST�(��j��̀�G-6��Xz�p�~�X6�ͧܟ.q�>5t}�ʎ�(a�����_a��Mйй�
�d�|#�(���w�:��$5ȇ��엿k{�k|�N��`f����J�����b����?!�qv/��+#GMY���AA���5~u|}N��#��8�����Q���ߘ�y$7r�эn��w���uv���Ǚϡu]�K���"M��dq��%��w�1d���g�e���-OݰN����6,��n��ɓ��ků<|��:x���}K��^8����tf�V��*1��٤���a���[2J�,B�0�0�W	���;�S #U��0��6K6��7:���56�e���`"C�)	�+Q�r��js�b+JZ`���ک�(�U6[���{>}m�]B���]YG]�٫n��>�O����;ݾ����Ӻ��f��{G�D.�2����~�k��C��t�c���*iϪ�v�W^��q|�� 6T�v ���J�E��-	��`��M�'��Н]Ǣ#��_�Z��Iݨ"��$�׋�2E�#{7dG�.�A���룰E;+{\���V�#h�@�-}v�{�󤯍'=��S�����B�*"�����;7$�o`_seMX�h���^3!Mt�+����:Y}}2z�������B�Q��� �s�s�뚢 ��T��M�-��Z��ǝ��hɑMf�W��ع�}x���{e�]Y���&g�O���6g�f���	t}��݀3=^��ߐHF�K�d�AF�v�MT;�U��m��(w��A�L�(r�b�V�U����T�(� 5؏��Y׽Н]�K�Ҽ���3����q��� � 3�l����\��u�̞������B�U�~I����F=���I�1�̆u���Z�e��;ρ��w(#F�}��5�s�ޛ���\�*��0�C�=��x�)�ý勭{7>�~maڂ�?AY��{��Gd����
�D6\͑t���*�_�M���M�N��v��ۘ��Ø��wV]�]�V����d��r�mb��e����|UU�v�OM@I:G�n��3 G�B�z3ɧ֯Oΰ��� �jd�����}W�ZoS�����x[�ﰱ7n��у�(Iub���q}����7޳�~֠�G�b��b�x�,�'�K�n�V:�E[��B]3��)!(L�̊h�z�|m���������zjE
q�g�ѽ n�|~�[����UP�F�kH�\(�u�����`\ϐ�A��7�Y�ky"��Y~�]cM�8�'�m��g�雹ݸ{|�9˄���4����i��9��|������&�-����y]5.�A�<W��8�t{a�FP���m�4��47NW]���[u��l�}�<�)3��f�͟��h�l�éVa�:�5���r�B�;�U��.5,�R+Nu���]�Af�h& )�)��-tKx�������X��X����;�sq��ӗ	.l�*!U�����qD�ꏝ@r�%F�'�Fwo�~c\؝�z�+��$����N�3"�B�x5�[�Kk�J�aݕc�=�9�\TT,1t�-��S��>}R<C�d���X��g~/5"�j5[������/.��Iq�PGcI�_6��_\���B7p<p�I��M���;n��4�\#�(��9�؀�� ��N���t�ҫ�ä�(_"*}v��˃7�_�Fd9�%&�m�`H�?#L(Rw�Q��ĺ걁(�m����M)Ef�K��X�(�\)���1���lDqs[)5en�`�ʍ&�h�4m3�e���@�l�1�tQMi�a�Z�R2���5K�,nn��T�p\���O�ڲ�+t�)6&�.l��-3,]�6Ne,}!�
��
Hn��[��uδ#��pf%o��Nř<W�����AR��Y��j}�מ2Fzc��	������m	<u� ��يT���ivi����X��X`��:�����ι�C���̀.�>�8��Du
C.�j���T'1eGK��ܷZ��q����w��o;�f�?1�
lՊl�vu�� n=�_�� ����}�l�tq�y�}��m$��Th2���Dx ?r��p�(_!>Xc�0��S��%�奒>�4�Iw�h�!���^�t-,n8��qc�>W�%�SX��CN"[gUgLغ�5)术�U�)��}w<�#��@[B��#z�NB�x�x�x��_Q�s<�ntyGm��:�̌��|A1F�	�Cw�v�C�W/��jv���t]��O�t"J��x�D�U �A�\�`�A4;�->���ڏefϮ[��q|�С:��Sf����f=�ڼ�#b]+	��K�q2����@�����������}d_e]��������n�W�@��++=�������!i��C�hI�4W���1N���]�@ ���B���G���s}������?��Z��}&�p��w4����P��4��9Q�	��U57�0+nW
3:�vU�aV��U�f�(u�;(�����n 4�E=%��e�Y�+�r�1R=]9w:�fS��ɒ'+[�G�]�G�t$1���Z��v��嬳˝��"�N#s9�Y��Ssp,&����7w��x����ѵ`��ͷn-;�]�(m:M�7i-[];�5�r���6�i�K*]�
5��n�N��gEgcS^R�H��=PN8��H:����Fw�SK�5:�뛒�&A�v�����УY�jؾe�S0�+�s���DY�b��ʵ�N!p�m
8�!9g����oj�:=�6���R�?�S�%w��o1lkX{8t���������r~�ȉ�f�Hr*_Ϊ�|�v�hb��ɴ�r�s�r�U�yc��y]��r�h�^�`��9Jr`cEε	�q:b&qm@é@t���^g|߭,��S��S��A�V�Z0%��E�$B(�"ߜ�ml�U���%�a�L�5��KNd�nAi�Ơ��n�ZJSv]\�TU*ب�lR�-F����Y�n�B�*HPQ7��
%��bXYm�B
o7y��#$I$E�H
R[$$�HI���	R����K�AE�8��JQF21� ��ˊL�Sswu5�	(�,%���K���)jI��*R�h�(���4QD�%�����aڔ��&���Ai���s7w�AEiXƔTE$Hq-,b$b1���%�V�Ѝ���"��e�*���y
ށ �� �����1	p�'�^�WƊ0В-��Z��Sy�<����:P��A����(��AV$5t>_�d�u�k�iy��E�	/���[�b�7������V[�����_����%�.S"aQԄ�R-t3�L￰�g������P ݨ����g��`\���zޮGɜ��[��7l�u�9�'3��	ݸ���7����Iq���~?q�~7�;�گ/}��T>	Z^TB����od��G�k2�RUUWEE�O�(f\���s�n�{$n�(���&gL�mW�U\Z�u�^��
�빒�6򂵟]RSOq.�½U�h��a4����������OkA��*�����������D�X�%��KH�kI�B3����-[�J����9�t���<�>�'AZYY�p=p��+��t��������폯=¢��]�6�A��G���ᳰ;ķ��k �x����Uγy��Ķ�m��9�d�������R�osv�B����n=�����Fm���lGWsG�� �PH��pޛw��.�hn���n�\t\u)o�C��*\��b�tb5g�Ah�nb, ���Բ�P�bivІ��;���L�"[	c���%Y�W^v��QX�0����;��n��wgT��-�]V�C��b51����0��5�*8�Ɣ��A�"����&YB��v�\�j͵�����}���#I�6�P�3L\��S7Z�;_��՟^��L<O��o�����
ܐw�ȑ�$��^h��-ݗTyo��}m�B�R}�%�_	��wz1X�����~4�]U����<�i5iRG7G�}uӗTf�e�^m��Os�t�m�U�-^r���l���!hOfr���������G��R%��-Z�~�p&�+2�����5r�Rdf��u�Z�����|��)K�f�4g����յQ�(���*t��fyODN5(	�U7�ϭu��(�;B��Э�<���&�~�ނdo���B=[ƸRZ�碶o�+���F���Y�jb��}�u��>�ّv��m����F��>�%����|��#�)y�sGZ	�T���Ng�^X��l�>9{~���G��p"� �}�u�G$�K��-e��U�Q����usLH@��#��ꊡ���w�i�I�N�Ơ���4���z����(秚�}��B�U�]o��o��V��i|�gTZ߼�4�r�	w�f��e<x�8�R���}��[][����5_*$�Ԗ4�̎=7:~��ߒ?$3���&d���E7�~���g����,�l�1m�H�I]�Vwze��ufm�ڭM[j;��yx_������C�Z��ɾL�X�c��K6��ı�HS"b`DL��F5Thx��_[S����v�S�׮��)Y��OLۋ���v���)�o���i��
��	���r��U>�ܙ�Q�����^)�cD��r/�Z���ȵs��mV{�5�=k����I�r[����w�J��)^�L~#�n���*��,�ҥ��4�Q�U*�IR��m]��z�M"��s��z���zm}����jf\�̻2�r�2U��33�E�W�G��+I��w=;�z�=�T��<��5F�6۽��6Z�.)??��B=����RCn��e�n1��g�RY�o:M�ɽ��MM#�q�U^�g�
���!����3�u�u�Oa���v��*�U���p���6�^vz�/�UG�M�.!x�-��@ŵ����-�uҮd3J�D���T�ͧ0@�D)g��xX�,c�[bE�tsR���*ik�;��%#tfĻ�.%���Kة�eG*gZ�֥Rڄ]R�.�H��g��ֵ��eRbܛ-�s/*2�8-n�ZY�6RZ����[���]��ԕ��)�#vs�h�B��_��=��b	���MBf!,و���̡/��QH��nwu5�Qq׵?{r�^��V����B�@��ꣷf����n}9����ڪ�0���!I��gE����z�vis����]�����>����}T.v{uq�G��t�^im�M} Kq�ސ��!ŝ��D�9���*�bE�a�s^��A�g��;��5JLX�.��odm˿��3yF��5�[v�뛽�/#2/�uH��}��_fy��s�%����"���#�iX�7������w��5<������7���F��������7�{�͚Ko#�e쫇Y���I8z����]�=������%"�|hTv�VD��'�Y{yx�W��{�!�B{c��	Ԫ��wq΅{����\����}./ ��)��:���z��|�6sX9wn��5��՘h#5(십�)�X'UU!Jy���g8=؇�ޭ�@�̟��ޯ-��C.��g�+��y�T9��6��uU뻬̭BO�5�j��F�/�sJ��ㄔg1[g��ncF3DF��L\,�P��Y]c_l��/��M���Ƥ-�A(Di�h��k*�R���g��}7|(�Bv��߻a��1_$�e@�:^�{g�ӓG?Dg���M���H�V"�2�F�]3�(P���l�[���Dq�\�(�"��_�C�m=�$��~�c7�GAWj�MLR��#<Ӫ�S���;9��}\�],��8ڊ���n��_Sֺ����o�U�b<_:@��
8U����*?{3$<�c���I<4'��/`�z�����&cKMhs�KvЬ]���Te��ԋ:�E
&�2OVVT��Qw�Y��l�-�j������|�У��ww�1�B�[����L�A�f�)6�����Ms*�e��~���YJ�{���q�̏yg��<(?��Z�f�[=~�O��}��K̙�q�ns�j+�x@̪����d����T��\}*��c�����>�x��T��=�L��u��x�Y���g�gZ<�Эgw��7�U_�/(���XwX�w��ƭlT���kY��L�|y�G����X�K������bb(-
�t	
(P������(����� ���V$#������M�,67FK�Irf�@ym��C����c�X=@�T�J�$�@����� ���@@*��U *��A�� ��@��O��h	�ei�%B*	H 4�� 4�҂�  ����BH 4���p@��� 4��   4� 4��\HH  �Ѐ� �  ��B @�@��$�ظ�Z-�G��PJ�@~\��7�D��1�C���II��8�hP�DHT���PٛyJ�L�c:�v[�H~>��ar�QY���{�`01r�eľ��x��D�Af�X�ETO$h�Q7�J\,&X��n�PC��x�����_�}`wS�B��* ��dA T!��E	�l? =���V>`��"�{C�����lC�$�����Ip��������Q�/��>���VQ��� 
��Ծ�?E����{��D�`��%�!��)���>.�`�m�4I��j��q$%�}v?߂~��U��x�FZ��4������}�������O�)�؟i�X�'vAE(���N���E����_D.�TD.�VvK� ��T�����(Aj�	YlP`<w�X0}����OI�h/����0PC�
R�S$�B �@�� ��c������ó�z�^`�����hF��~E=�����<>Jc�z��!�|��,���E��~�
/��B�Z>����Ϡ��"�*>Š#�d=�_�#'�'���	�;.~�y}TX��캗�b����}��i�|���̏�r|�'���<z�	�0���:?�>_��{=g�P�hu���A�8{x�������ab�����=��5JI��ET B��A T>���X$N�d��Ol)������������`3G�A��)c(A4z,
*dr��� H�"�5`��B���a��
X�
\�`z��=��t�vr�xL�(�U��hCj�ψ�֋	���-��);C.Q�N�t��" 
�
:�{?���p��� �QϸP����� �z_��S��h�����������ڐ_p� �|=����{ĸ)�>A�_"��'!�����@�O@}�����q�ؖO���������?a@ 
���}�`Ϩ��X2"�	�����?�N�?r�H�0O�Cm�����������<�OC���'����Md�$F���^�"��nO����
<���!������)���S������3�~s����e�S$�|�  
�����&t�BX��́Ap��4�D���O��I� �O���Cb�M�FJ=�F����H� Ͻ�y'�#A� ~f���~�9��������=��_� T���{��� �pA��|(r3�h(�!��ﰟyk`ʞi#Ƃ�=��@���WǓ����H�
	���