BZh91AY&SY���_�pyg����߰����a~�}  @   �A��   �L�      :@�P   c@ ��    ����    �0�������,�+�I�CY�8Mmhޅ�W�Q��C��6ΖK�^�{]g����Ƿy�nm�:w�� ���lͽyt^^���a}��   q� xj��lNv:v��r8���h��v�9�s�wFg8�w�_M|x�:��n��8xr�Ǹ��ڲ��<�v�ûs[v�wu;@=��5�  ���|��ww9�]�9�q��:n-�a�u[����``��rw��7����u��5v����=����wnZw����t�{���K�:�  �z^z㝮�;.܃��8�N����F0u�[�sN��To]��n� �nwWN��w]�`��ۻ�wW)�u��   �Ч��l�61���ѻwd�L3 ķu�gxx����f9�.vݷm'p�띭�;nv��                B@  @           �O�4?R�J�` 4��@ 	L$$�Q���&i10�#L LL%6�T�0F Fb` �i���5H��zU@���M4  4 4 "HT&�DdF)����S�4�MG�ځ�꟤�T�
y��J�2da�4�F4d �|ϟ��Td�e�T���mE�˯��O���#��no��1���.����lcz����f1��oŴ`c}��e[�����[���y��n���G���P��¢�Z������*	RI<��UU��)������ ���-B�j	��W�?~?w���>���&_2h��sBw�vNh���RxH��Y6v��z��n$��I���txS�keTׄNx�O=#�w���A&���rD�=i��{�:Ru:{I�g�����k��uͼ�w�zw��\�K֤֊w ��ܜI����������Y�<�N�N�:�:��J��d���Nt�Y=��d�;ϋ���l��'�?$�zO��%�z�'��i��8�RҏPp�,�+D)!��IZH�N�B?s�tJG��JG�:"?{��C�'<�`��%ȝHu�'�R>&�H��<?t��<�v�}_'XN�:����ģ��Ed�ߓ�N��5�����Y,ѧd�.$D�X��%�'�vO�3d�4DD�"/	EFN}6O��;����"x�I��vO���\"%�'S�I�l�4���e�8�")�	h�䲇���Z(A<�����e"%�"x��'t��"$�K<'�,�|YF��7�"WRp�_i8���(~���$N�xJ��Y[<�P��"_�|��,���D��<M�~<$M�ͤK�N�s�6O�O"�',�7ĉ�:w�2���z8Q�����D~D��N'�'���R���^D�c���h��K�<�=��y"p���Ή�ޤ��"j�lG�v��zX���\�_'�;B?_5S�S�oǆ���L�h���<��(ntM�OF������6�萦C�l����7�7D~�Mۈܡ9�A�:B����OzpY�Kj��V�#VT��/f�q4����6sGMh�O����]�'	���'yu�J��|�����=Gh��5��#˨�N�=�}S�9�p�^�g7R��LN��R�%�f�p��'c��?x�lu,MQ��F�Q5�"Q#R�˴�sPn;��Ӳp���D{8 ��Q�DG����|�7>AUD�B�g*",�ㆵ>�2�";��� �;S�uU]DFD���'ȋ���{��=QzbhӪ�#����8P�����gQ)jP�ڛ4?j",�6J��ߪ'
�S�a'��"<$DYV�#�TD^�ObP��R�>�':�Cdʈ���zjQO�j�"���TD�ږA���SŎ�#�TD�#ʖCZ�"<�DE�D�Bs�K �|�4�˨���7��d�v7uz�ꈜ�R�<�#�zMF��H��{ڈ�D�%�M�Չ�=���,}>~=�>�7�_hބϑ��!_2~8�#�G(GҏP��>��C�B��c���pE�O�J��c�!{���v�?,�5<wRĻjh��S>��^Eg�Y����>>��=����:u$O�>Cܟ �腳�3�k�SDD�f��Q�x�<vNv�w���:��Tf�O�S����)�N��NßQ��H�*P�|�|�(㢚�f�iE�����G��3j<�y�۳�r�&��;���Qު=�D]Զ�_�R�K$��z��un��Q�=�D�8%��rw�(��Ի���yʏyQyS��T�N�~!�,d��HU�=��Q�N�w�)���K�蔋U8,�Dp�tp�ԟ���߇��Kǯú{��>�psNԉ�|Ա$Պ�i���q��k�"�������>�Ǔ���y���yN/����_E�4��8����9蝩�7"n�G��ݨ��OI���M!�59�\�C���}'j�rK�܃�c��{6>�OrrڕG$���K�M�x�Z���>}'e�/u*H;�nA�{9�.���59Q9R�NT�K9'#P���A�!�Bɸ�[&,��y��w��c��_�=S�.D��<Vо����{Z��!߬��%�}ϛ�:�钇���8��Rt٧�p�p�P�IĤ��#�ݔ�_�i>�!��GmU���.�B��G���y)��؛�V�7;Ț��Iõ,N���zW��eY��D�$D}$���D���C���M�+�}�?D��Dy�_#�&��H��M�Ҿ~�Jؚw)��".�p�[�{��R�/̮�;�#�J���#�D��"=�C����H�w)��u+Ŏ�+��~}+bkڕbo������7�W��H��Ny��G��X벾~YVh���c��璓Bk�{�"hw����f���pK����lM"&�JN��+�q���Y��M���q;L��}rK)�#��ғ�m�C�>�O�+ޗ�d�N��E��*�|�"pK��<{�WO9����ԳR"V�rU5>}:k�;l��	� ��$Y[(�j�����'8l��"�Ou��[���x�vy'��&�r�y8����$���8�W�$u��}�w4>$O	ڏ��IӬ��d�\���rw�M5�Uq�]'Y���t{R�'��:�nG��rxsr�5��fs{��Mɫ�q��a1�����pK��z���'%JԤ����i䭾��FNi����s���/�����ٯ9�ּ�lו��檨jF�i䧳���g)�^�;&�����>��/��U*K�%j=�x�ҹ��Ԫ����y)8꫇�,��G�u\6^��Id��n�\���G���;!}$�_�ৗO��J�N����sF�´�5I8�O"/�;��Iy'=��T�K����:���p��_����
p�)P������f���}V�߯�X>E,`bI�ZY�&��j��:�g}�<ޣR*�[�D�l�|�f������.�y������I6^p��l5N*��uM9����|��=��Eu��U�ݛ�ć5����;�{y����4�;TOל�}u�/uo�4��O��:�?V9�|���qy��E��7\��-'�ʒ��z��ox������c߯+�|�]��AZ�\ѩ"|����{ժE�{;�Z��������ݩ+j��pO�T�i�.���{�?Nsu/KԶ":����9����۱SZ?"h�b���wu4�l\\�����R*�b�m6�y�,��Y6h��)�T������z��-�WU�s�n��κ�ɻ��Z=���z|u��?}�?C�~|��%j���*N2s�8�ݝU��D��������e���E����z���9�٩�ݟ#ӏyG�'�'�v�E��U?j�q�j�����'b�}���s:�S�g/׳��[��߽I&�o}����G�/Ϛ����Ȼ齒���}���7���/��؟�)�N��}ӻ'~��ӆ���8�H���n�'�Rɭ-�D[��ؖ��U{W��wb�&�k�]���>$�r��wڼ�gE�}�{&����^�)%���bi��*��k�~�[R}�o9gˋ�~�߽vgM5'�<�jk����#��n�tsW�ټ;�I��VL���O�}ž�"�W�M�۷x�����>������X����$���W'��4��\�5o2�[�f��B�{M5]����D�(�pG��q�ؚ�$�:i�lR���v����{y�ݙԺ�P��Y�gQ�ޥX�ěU٩����2.q;��uC`��W��jJjp���\J�$��ڜ��K�9�8���q�~����V؟�ey6��)%D�ShILrK/�����<��ZO�T��WT�>}�䏇y����7�xM3�!s�(�<����N��/4v�U�4��ƪ񙳢i���H7P�/�?k��&�}
ny��$�}���	���=�N�,qA�^�=o�ۅ���[�NQ�~l:�;��A�݈�G�B�Y�d�VW ��b�7KA"�	cՐUe��D���orD�����;;����!�5�ć;gw$61"˝�7�4��Ȇh�EAU�5�#��c,����/�^Yy�Я�5����RG�=W�\[��Ȩ9MJ����Β��أ�8����3F�m��76��[{T���h�,��ϣ7uA���R��m*��e�:�^�R��(�>+/"_�"щ������Il�<�W���G���Fmm�]}	�u�=s��D���>~� �ŏ�'�s��b�v��uQ��Y�r��g���-��#�<Z6��h��v�W�GP�}϶��<�����#�y��f�k��7Vj�X���|}�E�?�E���x�F�'ت �$�f�O"��&髣�'��!���/^}�w/h���}�}��]����8_��R�,o��LL�7Q���-�Y~����bGT;�Og�2p�'�'���'Ϙs5�����Ơ�����l����s'!9��ۛ��ŕ�Vf��4��1�N���3�	�M`Ž�wM�'�mX�x��XR���i�5���ȉ�W���E��[��f-Y��K���w5��>�Z.�g}Nj=�q2q�֛˛���/�ʲ��.!�s�_"w��{��j7Q-̰]�����G�;��>!u�X|.ӎ�N�qe�Y�bY"I\G�#*�벙L�V�[P�7��:^�5*X��6���U��E��x9��G��}i�ߞm��c���tt�Qx�梽/�O,�=�Ŝ�rgɯ�sF��#ı.����nw�&.!��y���!�7|lC�7���E���N���$�k�LK5Y��:��v�F�W���nTU�F٭#k#һ���E������h�G�#dzF�����g冣�|x��z�������y�zMm9P�Ď�5��1v�^.���C�q��<���%��|g��}��.�s�%a?S�e�=Cy�Jh)�s��ۏ���'�E�Â�j�, O��Y�mY�/������^���H�Ws���|'�泅�K5�}j )�Qz��bIJkE��x�s7���;�:�����>!��(�ŕ
�����^�Q�F�R���7��nNk������}!NL��s�ӏ��w�=����po��?A�}��!o���5��%c�2zү�s�7�,:��٭��o��l'�Np�Q�q�8s��8p��{�ut�e�&��Cz;JSE���k�7M�Yy�\�Ɉ����
iڍ�N�P�8qӧb.��>f�����4N2�st��V��!s�&��Yl-��ΰV���w�=��G���j:���b<{�;D�&�棖�r �r�*n�-$��h���G2 s��B�9ٝ��q#����(�`����e]dl�t��')���̼�7��h��s�[8��8�i;Ó?q��=�O��~]o�Ѩ5�.�5����<�:��'�K�V8��Ss�����Nr!�;�+��d6�,�oCI�9��{��k q���<������$�,�'2�K�p_h;��8�R�lZ�����;:M��{�Y��޻�{�ϸo�Ӛ�7T��j��6��*˛�vN7k�̷Z��w~i���Ͽr���d�?֍X�X$'���}}�N)���K��oM��of��w���|��]��\n��$�o�-�$�%؛f�iu$�Wy��x7o{z��Ө�޹Ԑ�Gx�2B���f�'K�͟�|�ݣ�����7$�n�y�7��E�M�w� �#�4u���K�A��N��9�o�vvMʻH�M�{�J�����K�b���bƚ7_oyl�篍k&�|�W����=�n>L���5�r��t�sP��=I{���x�^�w^�]��S�,B���;Zı"����g�o����x�u�kK��>G�^�}�b�'���7�'$Yy��v��8���;>�y�u�q.���^�J�V$���l��]��s���i�j�9S���I��M�_sx�od���b�3�Į��N9??/|��ő����i�Yyo��ݩ��޽�抵}������7�&��_����*��p��������\,R򜸥OV�Kme%-�$թ(ӕř(�V�TК�%�v5d%��RlHI�4���^4)E�"7IG
�.7��*�aQG"i�KGlYWm�cdBM\DV���ImC*b����Ȯʐ���Q�۔IER�ƲJHDϦ1[�Q1�k�"Hq8�mVA9!"��*1��؛�l����M�L�yTL���"*V�y	.ud�Q����Ƥ�:�"�̍X�X�vbM��������z�%jT�	1&�v�Q��5#L�cQH��U�����SVǍGe�<S-uF��Q:�WU�����4�V��H�MQ�[V�3�7��
�X���%�7N�M�DK\��6�?]��d�F�+U�)Sc+�nbmT��lj���T�(��q�"�k�=ш�2G*J&�n�F�65UL�����e%��6���Q%�D��z�qc��/6ҟIu�ۥzM�YnX�Q�[c�j�iD��H����U��O#X��uGJ�!2�j�JEcm�	"��YQ�B�CM�8�!iR�4%?�l��D�r{��i&>F���b�;k�V�,i�S"��h�����5����׶&�P׆�mR̲�.k�:�Wi�pc�p��Il��QY#p����Ɔ'��0M���E.<�(�q��#�E�٬i#Z�IM�M��B�F����uJ#T"F��b�F$��5�p�n��,���#��D	����rV)b�Z�w��W,l�&�$�h6[�3Uʓ+����^kݛr��,�&�A1�r��r=�&I����rxcհh{rWT��2$�L�GjjO�nĢͬj$2��([�֯ˑ���UF�(7�*��%���R�r�������V��$-���{!�����Iv��Q��yn=5Ƅ��PiJ����.DKƲ�(1:��GĹALK���l�	��$�"ma�2�6�央��D٩]{����䔸H�ݻj�����I��ݙ��+|��}c�?��X��� s�ϡ3��A���o��~��G�y�������������O�O�$A�O�!$`O��������9�"���U|�UW�Ҫ�X���UUTUUU���V�U괪�QUW�J�j�V����UU�Ү��zTUUUiU^���t����U�]���9�s��9k�*��B2$����efUl�j�7&gv�m-��I���-�՘���9I�[e�i>�[��_*�Ux��U⮕W���[]����b����Uz��U�U�]����ZUW���եWj��UUX�������U^*��t���������եUUEU�|nV̓�1�����i+l����V�&��� ��H$ +�DNs��5�yU�ڮ�V�v��Ҫ�WJ�j�Uv�ڪڭڭ�Ҫ��*��t��U����EUx��t��EW{߮�*���UUQUUQUUQUUQUUU�]H}��||M��|W�MXZ5r9l�,�= O��$'�}y���W�J���������������ZUU�Ҫ�V�UUUUU_1X��u�t��EUW�U[U��[���1UUQUUUt��UҪ�ZUW��U^*�x�� Ȥ�"A��j�ۖۑ���ڲ�Ke6.s7����ĳaX]q�&ܛ96Pܶ܃r���"r�^*UP~����_h�ꊠ0"0/����o��U��  ~?Y�q��>�&O����O�:'��tD��<"l�<t��A(D؈��� �"hN�bxD��bhCblК �$,DD�(A(D�D��"x�6%��6hM	BQ�O�� �6 �"Y��'
���4&�x<C����<�� ��"%��<"xN�%�(A%�A���F�M���U}�k��_̉qg���%(ی�9+�l��x�i�4BlX-5D�I���)�5W*+E������N� ��*��3G�cc�	:!�U�[q�����h�(��r��E
+h�ePQ�B�Y>�'�rnҎ�h�N�V��d<�#u�#��L-�j��b��D[P��J�-�]��y������RdD�r�*Q��-��IZ$�[pH���Si�piX��ǈ �9��X"���VL�LEv���������C�/a5CK(��h����I��c" ň�d������TJTWDɖ���F���j��1��F�eC�/Ƿ���$�\�*ވ�T5���$N)Y^2�CH�#�wBejc��2(S���#r@�P��*��P��Vc�-.@��AAbZ'\�,u��L���nX'������J�*R5����Zk$.F�"�	�-� !C���1�V��=Z�Ski �\����K%P��1̰m�!≶LL��,!H�0D���Ŧ���QZrإ��c��q�!�9�"��V��C��U.8Уiԫ��)P�iT2���� �iCBv�[ibv6�N�]�J�֭DEd���J�+U�T�A�jjYYP�MA'��:褣)!eH�!��e-V�6��&��Ua*���.Ul��Zⵤ�iƁ�R�-B�8�RRE"��:�lM��ɑ�D��U��&�ER��9$,lS�GV�Y:M[�,�M�2]�����	Z�u0�iWbD�#��K-����KI���x�#��	�b�"��E&�Uc!J�GRdn�ڑ�mV2�L-eoF��j�R�ݼ_���W�wv�|||fL����,Uywwk��}�fL����,Uywwk�}�d������W�wv���@>���:p����(�#�4��=���MbbB/A� �W+E�H2��l�cpxF�S��1�<DAL����6D�
�D������#���Z.mBBi����dțQ�b!r;Q6�ťC�t�l��v6�.Y)c���Q&T��"S"�ȓYn�M	�826�ڮ6$ۈ�0��I)V%�M���W�v���!�]Y*W��v>�O��'R�(V_�.��nw!A��f$�	`(�wۊf&�93[��27fG��$���e�Xrmvu��
�&��÷D)�=o�IU���54�:�l䆦�$2X8\ęl,��	$�;�����1ԓx����LiƔ���R�S�y�����:p��F#�Q=�I%��Ra���n�875����a���wp����c�j;.�,�Ζ;D�F����N��88B�#���6����1��Ա�I�q=�L �v`�Z'�}�;�Ζ%�ç���x<x�N-_ �^Aa��m$��΄Ɂ�X1�	�pٔ�3L�1�/���}�Z%����R��%�K	d/ �Z*fb�p��f�ٓ9��<��4<��ˆ���-%8�j�Q��P	W��$nh髦��r]4D�CZp^e�y���Z�R����(�!ӄ=����1��$���b�g�ɌY�4�|"�n�i_��c���e�f7%Vت!�;Df�3��V�~�V�O+����U6�n�PM�������ݳmRWl��U� ��x�L�B�L��4��֤�9�u�1��q����O<���)jyO:�R:�M�sRg[orJ�rY,�q�"����oZ���̬B�Ls]Eg �S��b"�����,��y&Ɗ��h�e��[�Z��f[0�����dm�I$$O���sϹ���{R܅<r�HSނ^!�ͣ5�l��.�Ny4T�\�إ�
T��.�nC�oLՋV����6Wf)���jI�(��[�o�$	F�.9p7l]�Ce����Q*����=�E\��l���c�2p��x$����k{�D�{�3��I⟡U�e-MiS�ITbHZӷ�&��r��`�]%��jy�<�Sμ������-3�Pm5)�ܘ��$�cdL��k�"�ٍ��D�84^24q�eɒ��P�b����`�e(����(nLb>�NX�B�%�l_Ac �i����HۛI2�d�"t�r9�pUTX4��7l؀Ga$dvZNQD��vO��eſ8����u��t�CI1'6$�H��1eǈw�)]��>�Mg��P���m�##�;5�7D�6ؤ�S3'Dzֿ}Ȇ�W`FWr�D8�ء����ϰ�"4j������w<^���HBl|��ϴSy�b�C)�~�c<g��ܱ_ї�o���|���(�#�����`��Ȣ~I$�L��!��݁wo���c5lQ�\��\���s͞�n��:v�Nt�k&HD��֩�+�D�`�V�|�;\$�2;M�� h�W��;��Z\�ڿ<ֵ�Xdq�a�)��j$��?<��Z�Sμ�������{�"��%E�Jݸ��V\)nL�b�i21�J"bP�T+ZHHI��m(�X��6B#\I�m��U6�(!L��U�*L�V��!d�4��I$2�U1�՞;
h�9YK��6s�8�G7�5F�&��	knH-73��w8pY��#�WW.s��ړw�L�
\��	2I@����9pXy��k	�p���R�Ai�&K���p���Gr��%��� }|�)aȴ��dr!���>ጙ��\������?-ǔ�Sμ����Ӝ��������7*lłFݜI$���Zņ0	�U&̽�t��m�:�D$��1�1���oM1&�&G7 �CM����B`�ӏ�9�9�H&?�|�����M��0�UZK㡃�&�\�FC#�K-�#9$݉20�o�VS�K0�>��t��쇴JzM�4x�d�y�+y�-���iǙ��Yp��a
Hx�0�TL&��n3iih��[��-�6�-����O���N�o��>[/�iճ�NIl�-M���gh�Y�?'ȽI�|�����'�3n3��ZZ��0�L8V+���ɕ(�rL*��L�D���D�='��'�K�򸗊��Kē�./��<�[,�1i�'䷙ŧSii�q�Z:�Oɵ�M�2�=�L�L�ZZ�)Kn�i��s%�[6��6��g�fҗ�-<���8�fN-�#�jKfy�[�<�K��K�-◕��~FR��E��6�V��}��%�uLHB_������}W���U�ʖ>���T��S�q��K�;ޜ�Y�p�l~ֻ�h竾��Oy�|m��^ϸe�w�v��U�����E�[r��=�K�.BY�Ͽ�|t_�5Z���߹��9����~{2*����Y���fVfs=��ə��{ڸ}�ٙY���{3+3.���8}񙕙���\�]�?o{��c�:뮸��O)�^Ot���b4ڪ��a74A�8b=��kUV�	.�7(WL2?���I�Ң�a��Ձ�Ԕ���	ј�q���LF��B���γ�Q*&"��Uk$�����kE�V��L'6Pz��l���!��1c���$#)��(��a��n��[<N�[�ht���E���XA,����`2�B`bs�@��
Ja�)���Lس!c���B1lA0D�S%.X�.��f:p��/>uN��,��E4�m�/����*�!
�t������$�!*�ƨNv,�	f�D0h��F������X�,!�iB׵`v�L.	��H:a�H��ؤQ�8d����q���bYAST<*�-�D�CO!�3�Ha��2S8 m 0�ht4`�^	���'���	�0`=�B����a���������1���Zs2Sd��e��6A0Z��Y�eg(�v�1&�:t��'�S�yה[�"�u�s�<�:��1�&�%g��ѱ���F:��
����r��d\B�:�+�XrkR�F���͢�j*�lCSQ�q����wV�H�,f"�812�����%Ω#�q��vH�m!�YT��89\*��H;l*�$�uF��9q#���p^x����F�9r/͂G��u�4[,��u�.v�1�����׼X��gI�(�}r�q��F�}n�%�P��Vu%`����)���b+�����$�Ƃ+�B8��vEut7f����xbbpR��[SS�gm9���t�M�wQ�qd�Ě8�o0i��ԐԌDD�~��B�r0����a����J@��%ن�4:����El�&ʦ�1J�F��@	B�tl��a��eB$��� �����d!2�&��c�=2ߖI� ��C��T%U�J���t��M%	��fŝ���W	F{4�zJKHB吆UyՂ�l�8��8���<��)o	��L[�C*˚UUQ*�X5d,ĳLC�$D����K�H��L#�E���,��ju��O��g�mƟ"z�h�<n�3�y>tv�B�r�7V�i��804�!�A�4��CQ�(�O2K�ѕ��k��r�1߽��q�m�m&�����t�no.b`�$��;	0�9-���v��g�N��|kq�s&���q#DkL���[i�p+�mO-n���)�u���8a����zBBEh���0�x���U}:�U�;P4@�A�㺔y��D��ܒ��l���)3#���0$L�b�j�.7�=i����Ό4@�Z���08�����(0��ޟ6Ą��Q�)�rL�1����$[������Θ��v��N�>�rw��S��[�7��)8o�[z����3&�HSpz�݃����)��,��Z������A�m� �8fU]2�x
"\��c�{��n�*}VL2|O�[�|��<�μ���2�[m���! ��VƲHe��j�7v���Q(%P�\IB(�gHa��`1J(5�F����<P��a�"Ѽ&6��Ly$�[g��E��e�����ld[¥J+�|9KAtE�C�N�˖�G=Dj�Yv0ʱ�IM�8 �hM�K�C�He�u�]�l��AG<IE������B���Ar��xSa�Y�f��mg���
�^��޽���XI�Gq���O{۷lJ����=a��, Q�$ B��EN8�t���<p��Z�y�^QJ[*u�TIy�?rwd$kr�,V�R����׷V�5o��w��!�����11a�B!3�����7��p|�G}��{���$�jԅcO)n�l$����bJ��������}۲4�q,��M��79�DE0nW\S�g7&���2Xd�X��9 ��7�t����ђ�b\zؠz[�1��T#R��W�A�B�[.
*�"U@�J1�NQ$���E�d,���(
L��(u�@9i[�$(@�] )M1J�Bhz4��J��p�X	��	Px0=#0@��g�B�M����$&,#r[QnT294U�JУ�W �)G�y�� �mѐ�%�&ɏ�G�-O�[��y�yAӤ=:p�U4NJ�$�Z�\�p��UT@��J9R�)+d��9NjXn@t����`7P(*�f���f5�N��B>,Hq�CdtDɲ�fd��JK]1�J��$�6�ӏSb#����1��k�\��_؍e���F�ぶX�1l�B��4p �iٺ7�T���M0�������-w�Ǣh�]8@7��I���bo,Y�3�;�ㅶ�i�����ן>S�<��)H�:�{�������r���R��Q��7�� Q��{�B��wd��Su�Ջl���u�D�TjU�!���T��.@���cƛCB�e�D$b$h��a �Z�5���Ǘ�fQ�	h	�\�*��@��w]Dc0��@>(S�+ւ���eX0:���r��W$1G��F*J٘8KX�e���5,�r`0���Ō+w��E°��
�(h�}U&t�#�m���:�-Ky�^QJGV�l����LH��Lk1�����e�w��UUH���vо��ʥ�T�s@��F"z �xB-�0��B�B��<��;��7P�伌���M�%C?���� 5�UU`��l(�]�S� �{ZR��i����&�L}�1��cX�!�C&qH�Lf1�Z>G"󽱪�T�`[0S��&��IKb.���ތRE:�L�(HǄK�f�ŌKq���8��r@#z�"��8!�e>�)�4O�:�2�Z<�[+y����eh�0JI��h��a
D��VaDO�im-�Kq�KKKO%��)ii��il�.~����n�d[��c�ų�NIl�Ke���ii�e-"ٷ��ե��ճkg�n3��Zٴ�ٴ��������3���D�������0��F䞒�mfE��#W&q�I�Ql�"�"ӌ����H�2�#�)?'ɏ����|�L���Ye�6���^�ǙR[Y�ͯ2ٵ3kf'����m"ٴ���--8�m-��i䴷�ql��\F�IiȼI-$�id����و�4����i�l����s��y��d�}��4g���}�����"կH��[�m_w�|�g9d���-�e�T�DH�^Dx�8�ʭ�oQP�Z��||�^�o.�[J"G�����S�Y-k�V�u>�ݓ{�(ظأ�;�N_9�Z�v6�R��}o6r^]�����;ؐ���t�ի�I��&#�ۉj#�Sk�����^�ntՠ�$DF��,U�F�Dn�TMI�i��[�9�$R�|���M�M�;튛�i��N���� ��KB���)�|�T�瘩��ٖ�gۃ�9��g8������޳t���~.�SO�������]�ުS��+GN}a���n	�)��)
~_v"_��f�eH�Q6�~��q��Ec[�ݜ���H{�K��e��G�(��|sa�N�#`qD��wD��n�;Q<bͩ��`1�Q�n�K�}!�M���q�S��,;?9�7�y��Ͻ�>�6��^O�9x��ǎ��J{����-�~9�{�_/WRK�s�6N����rz��O��tBX������R���W"F���(��&�+h���Ee����ȶcI�=�����)!!\V�h۶Ƞ���l.&X�1(�+a,,V�QB�l �Ȭm+$��F�Y�,qT�rE�e�&�V��t�Ů�Cn��<������%���KSX�j��v�ڿ�WM���_j��d���������ӊә���y��33Y���V��r��3�ffk333�ҹ�]�f{���fffqWK��.�3���(㎺�ZԷ�u��un��gъ�AL��UJ�cD��ML�uԖX�Z�H�t�1R%�#��Rd Hx�h�qh�4(8Kk+e��� C%�n�Uc��W��	�����U�eR1�8�Pk���k{���[c!�*��R%TqA�"��ڔƫcA�j��7&5L��6��^J���)�5x����}�>m��m�uS��H�i��w9��:�j��)Ӻp\;�Y�E�q��y7-{k7Nv�uu^w�C����`�b�L0 "|A"�0S��@��Ȥ5H�86BB�08�[("E��=�-�4�n\���BQ�jt���XN�,l���R�R"Λ����Lw�����\i�BwħdK�y�Ƙ�`�E��X�:�S�~df�&�#���j���	b�H�-��(̰M6�W���b�݄#���	]�T��`n�?��hi\�@�!H_t=��UEv�Ob����|�N��μ���y�O�N�������ۿ l�<�UV��dM�,X�.�� r�5�8HB	�&P#�x�%��q�,�=mEѡ���Cl���C��5"�c�{4&n<;q�M:(u��X�����#d�əBt�GK�im� ��E�*�d-c)ī�Zո�t7؄!0?�� d�x�^��>(l6,@�D�� `����t��ّ�p8СO�`{�u&$~�)��x<��|��:�Ϟ[�:�R:�[cS�Z�MFf5"#VI*kJ��@5]$�@ℬ8��.a\�������t.X]�!C]!!~I���F��l7 5C0�
T3�26!:���KXf>��c��4+UxB�ȇc������:�$��i�X� r4y�|Q3%T%z@2���ÐO6�Ƈ����
q�z��kX�M��<�CP6(!RBJ]��w%���K%�47u��'��=� J=F����b�4X��G>uO>ykyהR�պڮ%�l#m��UUT�{R�P�J՞�̵U��t<�l@��p�i�g�#=r�<}�vDD/�Z�1�E�[*y2�-�%�HBB�L�1��Nz8��1qƍ�..�L�Ʀ5�j-j2=,Ga�Jz8<=@��p>4h�o�#b�h�w@�u!#(s���zԕO\�L`�Z���Wp ���k/>:,I�s!��Y��
Ԓ����N8pٓϝSϞZ���)H��m�J^:�&z�B'9#��m�j���P���E&��d �!D59�Cb8�(lܼR�b!�S��2�Q�B�n;�k#��"�*QN�6�0M\.]]�R��]$X,d��:����n-�&�^�7�;ބ����!�aQ��*�y!ĵlw�9ǉo6e�m��sq	bI<��<�y��y7y��'}��t߉���%���l@#N:�Y��
R�&�J��	w%���ИD�@hH�cx��IcX$�q��ꒋ`�]�2]��ZI�&�IPَ#r,n@�A�M=��>t�N���Z伫\�Ō�!�6�ĥVڢ���\/k��t!�,Ӗ8؁� ��Q�8t���B��6.X���N���yk[�QJG\[o����*��*�W��YR�R����鲋U��Gln�p��mD��6nPh�}�x��UV�8qOKs~8@8n�. �ō�)!��s|#�ҥ�I�kC齪_Gm��Hq"K���KF����(�{��򄰨��	f�dQ[���F�46�7 ` ��86/��!�Q	*��g�X3օ��44@�cKTI(8�ѡ�u厼���q�>|�ַV���,���J�	��UUHd";l>2P���l���\�V9U	���эG���h�d�=#N�:	HI}̺l4 ^�"_0������e����j��J��̻W,r18�����GꜾ>�
gL8g�%�x\�ڐ6A�I$$�8����2�����%)�d,8|�3Kw^�!~7r@,%ǽ�4Q��N�X6�Ua�jnXH���lX�y̻����>�������ϟ8�^|��n�E)q�ޓ��3��\��q�� BJ�n�a/=UUR�s�����;�Ǳr%:�*�i!!��L��6�e��19f]��p��Gv���5�Ny��i�1�hl%�=�]���!�����n:����$��Ǉ��8�W�f��ʐ�H,a#p�}B�e2�N�.�pqG.ۣ�i�ޱ�2��ƣ8�?c9[o-��y���Z���R��o�57�p�h����Dj���`��]�8�1j�\�m�D4c�s"4����*V�ı��%�F�s|���kQ�Q��*�=��Ԩ�o���d�UUT��Cy�m	���R���ir�+�n	��lN���|��yÜ�9�M�&j�x��táv�f���4�MzO�>s��=��1�_��I��2��:I	�._%�{�Cq�y�d�[�#d�/�O�˙4A��Ƃ���ZG����D�������=<�i��^��mp�Rj��x�G3:w}�<XaC��~���#Q��_����<��:�ϞZ���R��f٘�q!���ԅ�1�趙5ꪪ���ꕁ�aW\y	.�,��#f����<���ৣ�i�tha�o���%�{^I#wz	hԞ�Ir`�h�%��5
�H0���a5;�- �3s���b_�!Ao�BF$�DA�LG��C�l�K*��B�Z����]�������s����S�C�ó�06|�2\��Ɋ7R�\0d;ys�!�{!]��7��u2�q>L|�KE>eH��D�	F	XD�0��a0�+f��y�N���KK[:H�m-�m---<���KE�R�m�ii�-�S6�$���ٓ�d���ߙ~JO���de�l���ٴ���-���ߙ�Yl�Zil�[�j���h�-mG�'$�%��r[-���L�>|���L�H�dy��֗�Wn%�K{R{^�q��V�2��Lu���JF�jg)i����>&������χ�=R�ͥ��o�e-"ٵ�imyl�8�m�e�O%�����ql�1��y���Kx��)x��FR�i�[l�[+F}���k��v�z�|�ˈf���zM�;+Vz\7��~iK��o�o>���}�53��B,������K�Ro'�vw{E����N�o_\�u�>4��p�=z�O�!Y���???-WKy�]�gs33y��j�[�r�3;������U��s�y����V�t�|���w�q�]u�����KQGHp�g�	7�UUT��ƵͱI#��%]t���	����֡D��W^��NKݭ���¾�,4�̡�K� fT΃�uD�"�l��dd���	.����F����\�&�!ø6�6 dtmɐ�3�c,�C�ŧ������S�6p��gΓ�ɀ���6���s�[�ߊ~^2���m���:�V����o�uƚ�5�M&糜�9�� A�Yۡ��pk)��L�g�k�p>����dN�$"�)2����c}
ҽ�q�Һ��w4�q���1�J���u�1���k�i������G�1⋄2v;�R���B�͙�E����w�~��F���:}PC5��2����a�,@�9�bQ��Y�k�I�'̨�b2�=����V�o�u�V����o�uƜ���ӂ���`ͳ)r"b���ٷU�Z�n͍lkvc���魆׭Mbz!q��3Fd.\Eg��ݗ�PZl��Ҩ�O)4�bZ�q��b���L�[���Ě��-��ܕ�*���!"��D�e�2�e��c��UUT��+d�DuO�׌Y�wxM�8��8�i��N֧;ot���Ҥ ��*�l�#�Іs?�_��ڑM����I=���=|�+I[�as�.��2�t�6��� H`8�V�h�$*�07��I��á,62vX�ɉ*�^TlT�A��t{���|�cԼ��#%K��ׅ�y�Il!*ܻ �,9.KFGbBJ��J��UV��4��,80�#,\xx��G4p�Ե�j[ǞE8�g��D�?~������J�*aG))0>�Ї�%�pvd�ҹ��S�̎s�~�Đ�m���y�S��F�,����'I6t�h4{�\�ݢ^���Q�m���Z�rs��p�zQ�ך�9�I�������~��x�K��>e?>c���6����庵�yo-j[ǞE8Җ��DBE�-H_�#�Hо*��
�g��h*�kEj��UDLɜ�b6[Ɲ�?-�l��M��,��h�����6�G,�']?�I:�81�e�Ȣ�2�,S��Mh�îK�<.��rύ͜##��F��*%���h�� X��Å�p`�q�͘;8�e�dpd ]Җ�Y�^���H�i�κ�T��-疥�y�t�g�\q���7����Û$���ƛ��!�J<����x97�EX�Ϩ��`C�^�"K�6�M�ے]��e�'nIgi���2�Gi������b��F�?o�����L����LGp��뭱l��ۍ^F7(�(i�ϋA�R�G]&G��k,D��I�h���,��+�?>b����)�qź�o��ז�� �4m�[ѸjV�SU�Kkҭ(�7���e-����pYG��4��J�^!q�6 �eC`��eJTDŘܴ��3��:�z���C6nF�*��-�s�s�9Q�t��o ��w�\4�r�bW3�9����+�!?
����*�>O9J ]��񆶼t6\�\��*���aD}���繍)�2���u}c�b=	teJ�b�op�T2tᓨ���L&��ǚt��c���a�#!vX���%��R��6�2p|Q˞abt�1�w1���>Z�|�-�kR�<�)֛*�m�\���UU��ȸl���u�#����
c8���X�@��4x����4s2\�UQ���,C݄!%<l�Á��0C@u���^Ǽf'��FQ-gc����(�7�D�÷Ňaa�F�p�b����rȅ!b�ӌ����lI�����=<)�!baZ0�d�Ć��Z�ls����p�,u	rn��1��ǆ�~�p|���:�Ωkyk[�[ǞE:�[��ۙ�UV�T.��\9�V�7=���r��F��챙��?��ZLDE-�l�8+���GA�~WYS��p�W�p�!��Z}���\�����Ft��fԱ|�!s�6�p�B�3R�2�H��@��񈈱�4Ct}
�XCGr�Ə$zpX��Fj�7!c�i���_������|��yk[�QO���bTG�������$k�ʎ!p�瞪������bK+�/�BE�J!q��!.q��HX�/h�,��+0L�-Qn��9BBBHq�\�_{=6X�*dl����f��܄��D������ ���α�4����lm�w�lԶ���ؐ���65��|A!	M=��D�L~u��8���lg�Hg^5�~��E>eH�Z|��d���Zy�*[8����-<�i�[(�[6�6�4�M���ͦ�3iiĴ��ճ��ZD�[,�-6������iIii��8�]KGd�_���q?&��d�Z[+j�kf����-�O%�3���ɛL&\������"VL(��r��GD0�k�BY��Id��z�#�.9�UӉx��Kx��'�V���Zc�����R6��ǂ��WDN��N'����>/�L����Z���)�������-�~f���^����ů3��̺�<�������xO	���)ZDZ,��4�K�lܟ���2�}���������.l��K	�5�iY�EP��[EQê����,ҍ*۽�w6$�ydJ��4D7T���e���'�� �R_S����7��䧬s���%������;򚥗Y���{�J�6.����~#����Ӟ6��j1B�YH��;Yu���)�}|���8޴�k�]��+Q$%��|���Q�k�%WsfUCM5�m��mf�V3x^f��<�3���<ro4>�'����K(��!ӥ��v�����{�>�6o�|2���|��B5�y�-}�M"�O�:<�8[��Bh�2�
���	�����c,!i^A�m�jN��E�j#�(��K�B9	ŇF1	�T�h��gi���VůWw�ϱE�:W��k�}��x�ovv)=�\�=뷩��N�{�q_������k��n��G9��=�����;��sǱ��}7���sn�9�ש�I�Y�S�~�NO<O�R��JI��\���\�P�eV!���%e"����:I���E���B��A�ňCyd,�R�����}��݉�[q:U$n<II%�If*6Z�I=�.=z7�[n�qF���%V�j[u���X�^��ƑrK"�6���Tğh��lYF�(�����h��jk�yY���f�t��.�3�������Wm�s�����j�Uv��9y�ff-��U�wy����YÎ-խo-kyJ)H�?o�Τ� �s�,e�D(+"�5Q����$*��h�Ҏɪ(-��[ �\��e!q�*Bt��lR�Q쪼W"Q@�+pE11,�"c�%�J�	rT,&:�
��1,��,"!2R��u�%�V'#�*�(�#�ZN*1Ti��ڝ��%Dh��4&�!h��qKV,�:1G �I�fG�*�}UUi!�C+H������KQk��	�f��S�,���*��ó���4�,L8!>�b�C�a�ѕG0!AE1���qI'��#��I�q�J��$������[0���n�����.C\8�0�'�6�W�6!
hp�x��0me�%!���r�O܎��>��^7I�AO�o�!a
�g�z$XHUY2�?��~��٦π�h��V[�<��gM<yן-�o)E)q�w+��m�{�ՙ5ѣ\�UU��0�U�����B}="B�������b4I$!�˗���x��چQ�\�"�қb�$��͢��Le�̞c�#�ec2�鍞F4��K>=����=��i�ʁ-n2��Z�l�BHF��C�6V����<!���LnB��zN�C,9z����rI8��L��m��[�u�<������u�ǖ5D�v���A�����C��i�3U1�?8��yH��O;��(�-��0(ȕ񡲟�h��BPk�A!�'�M���F� ���e&�6�mj��پHdk[BČ�㓧F�F��Zly:8lBK�0h�����4B�^�+��:�!ƪ2�($[K�I3m0ox�O�v���~o��)�]R�<��JQJG\i���W'�|�UU���������E�%>�m���2�=���_���� ���6RVU-%(�J��KZ�ՈI�.�9t�td�7�5�����ta���Tٳ�,X���<�cY�*L���z�k��%�'.��I1-lwc��J�܎Q�!�SX�B!�e4�C���82C;�b�>8ܸ��4��mn<���jR�R:�5���E��R��+�潃Sc��U������t!DƳ� �D�$N*"D�
@tJ�ȶLo�v��"֝H�M����%��V�������ƭP�$W;⪫I�U�����Η�g�������M>��p�)9'���/��t���ߩ��Oi7ɲ]������<�j$�>}��6�cf�m1x�ď8\<�%�iV�QE��d.`�B>�%A���1�c�@�$0ߣwc��HN�0@.Ṝa���[�u�2�6mM)�#.F�������%�I�X�ˑ.g����4˗!��&d�y
�!E�~S9�1n)�>yo:���ֵ(�t�.�ʓWe�D�⪭4B�P��ǎ�NC$:_6D��Ii���u�M�2B�# Pǭ��Z�Z�Qp�vxr;�`�t�cC�rT�lrh(��͚a����sh�rT�&ƾ�!�m�	[b9j^T�&K`4i�܄8���=y0���l�>slM=���8�'�!���d ��00�4j�z'��O�:��<��JQJG\i�~\Ͻ��2�⪫I��g+Et��	P���ۨ�#o��DR1~��j��/h0>v�t�rܢ}���R�{)�F��$�Lӆw�6.73~���(�6l�pB�hoc^(���IQ��9:�F82�.�zI&~mH��ߑ	�e&d�.�����m�rx��%�E�q�i<�-o-o8��uư�R�Ia$�Rd�ڪ�I�-�w�g�c��Ј���|��ۈ���A��,c8�-JMn��%��#NIIC�ݱr!a��q'��L���r�X�d���rX�!,a�\���/2��Hz��L�)�BFplh�����3}آ� ����������i��u��ϞZ�~R�R:���;e-q�kV����[%ȡ$MD��D�0�#�����b����6�J�u9�F�K#��Z��&%�H;D�����Ͷ�o�)�ۣ���|����9��Vquݻ�9� �>�噇��9.���͋��y�v���#	!!\
 ��d�<�t���@ƆCw^;	*di��i��`�����Iй�x�������+���À���\!9XE�6���X��b��1bAi)Q�R��l"I�i�l���p�Ƙ���B�N�s�Β�_u=0ܹ�g��y��[�qJE2�5���b�D���e�a5���6���B�Y(��������|l|`�q�ۘ5����`���M@�f�(�60��rz�Xѣ,D��L3Le���i�Ա:Ab>&���^ʖ��|%L>�I���&�$�!�h�/7$.#�0h�d���UQM���C��J�+x���d�)32��qKy�^q�âxO	�<'���xD�<t����8���BP��btN��ň�8&Ĳ͚D ��:"tЂ$b"pD�:X�6$4&�(J��2|�!��bhK,D��Bt�p��l�d򖶔��jZ���yy��xN�:!�ĳe � ��QL��blO�ɽ}��9n�_4�9��~{ߎMKoUD�A�����$��/����߾ٽ}�w;N�\�����7��ﺸ#y�ruG�ӟr�v>Q7��?t�c�F���Uo7�u�~{��+vp��%�z
n\K��~��_Y���5�d���9X���������z��ƪk��za�����1ҫ��󗙙���WJ�ۻ�^fffb�]*����33331�U[���fl�f�����Z�S�R)�\i�X����UV��SMn��ˬ,���^#d�y>_���6lX���-~9��y9��{l;!��J�v�j�MAH2��F�b�,��o����Yq��<���s��X��3���h:87���cr�(n\��s9��xrB����\������<q|����-��-o)�JE2�g5)���yYʪ�����ަ\^ʬ�mzIWi�����(���Z%�h�\.��9$�V#-ŕg���I$��i�XF�Ι��=�E�$�A![焨(�0���e'vI�!sa��&N&�,Cj獜������$�\x��\px�A�i��M�ѢTx@��ƷU����i����	zgۈ��y�bz�����?<��yo-o(�ǄxgNd���1�"��֪6��SmL:ȍ��[P˔���B�Q��+̈́�9���%�Znӈ�Kg�RiHۣ��Aڝ+��;pv��Zq$��ݻ�ڪ�A�l��^��o�y�8�{����o�=zL�ʑ���jo��ټٽn����ٹ�x��'��xa�n���EC�m�F�r�#����*T�xْug����<xω�����-)��ڥ�^�=u���rm�<�	32�q�m�c&q�8pk��p�����gGΆ�C�CD}���]7rD!�kI��YAh��5l�$B�ܲc8��z��_#H�Nl�8�#:��4��0D�0�<Y��<QӇ=�V�J���KǼ�UU���������1�����`p浫S
cV�b7��"d�8(x�"��&�CGYGK<ё�F�Mǽs�T$���E�Y�C�N�Qrkmxd�Yc��dn�Fr���SU���d9� �-�>��T6��#J�5q���q%�!T]0�r4��h�|��qo�Rַ�ڔ�e�	��o�ⵟ�jI��/VJ����l��UV��)=�5�JW^��d���X����q!D"�,т0�'/�p\��%\�Śs9��*��ҮD�!!U�i�&Qŋ<�h�7$b������i�G
"d�о!=L�l(xl����^0Cx�d��Uh��j$Ѯ`lh�X�u��deS���
��,������M�8d�)k[�mJE2�*{9L��Lg�ꪫI
�{C����|1{[!)P���&�$�[���������"��� Ȉ2
֢/�4�5)%�����ϳ��������Uގ��������т=+ɂ�X���=
k���"��B�l3yjK��vl���M�3�.nxr��HIQ۶�e�[+�c��<��?6��<����<|~?!��<3���z��LnG/v&����͊"�)��PJ�*o&�Ѱ|aK�Z8)�x���:1$�,�$�h�dUL˷#�F���UU��͙�&�y�n-}-�>uS�i;�w7�����T��U]�83��'��;�S?g��h�̴C|cX}�$�L�ZO<�/y�_"xv�eQ�%��c.ٰ��D<A�ǽ1]��J%[E�@M��h��>ç�����a�[�i�p�0��MȀs�K8p�!�G�#�!��V��T���D-b�*�r������l��d�z�_�e��J|��-��ykxt��HtN8\��'�eH��UV��,��J,���[���=�Ģ��R·��ݱx`�`�G�w&��<��C;ra�⊬�(c��Q�h��(��v���T���[ʦn�������,SUUw�~u�RJ>2B���\p|-�d#*�d��C�n�11�8�x�n�/�6��-N>?�`�4x�t�����{�;UJ�Byʒ��U���\�&� C� ��|d�y<$��}�}��h��������	7h�a�-u+%N�I��<�s?>�w�i�dI�2���a`&��力OJCt#��I Y�<Y��6��t̄�,�:�|i�I#4:B��k^c�����>R��|�Z�SJQ��g��M�y{�o��^�b,a�e�Y�S^*��&r0c<��q�g���Z�^:M^�Dz����/�T%A��b��C{��Ƌ���w�A�g��E˹�� ˸]��6��z�RI����ӥrO��7djIs�� >��~@�1evJ|���M·����ẕp�bvŌ��`p�����&�6~?C	���tD��tO��:'K(D�"lD��N�D�'��%��ň�BlCf��d����'M"A6"'O	�N	blM��4�BP�%���'� �tKbYb'���%�?6AL0ц"xN�!kZ-kmk[�Z�y�{O�?(AADJ(DؚO��.���nICd�z����x���Vfd5��n���I7�u+E#�I�3e��F'Z��>p�a�E��S�d���Jլ�֧9bl~�z�4ԁ�ڨ�Gw�7{ӱ�T�'��V��Tb+n6���#U	׏S!V䍻^OԷttn	F�c#-Ej��?�ۛ�>�rp܉fŢ]�����B#�!�{���*��x����P�q�LC!�Aш��wI���SQ1��BL�2R�x�KD��(ٷsfb�!(�I���P�"z("(��X�1Ҳ�D�ő�ԥ�F:L�t)��Ǹ�\�	�XR:L�%.L;Q�٧�k���~�᝾Tw�Ϛj�Z�5N��߻����yqCR�:�ml�T�XʕU�ĥ+HUlv���jy#�;ݪ�4�����(���Q�+����qZ��J��&*��k.5-�*J�y)%^�4k\SGH���ˊ� �ȕ���]��X�F�)S�N�MRH�~U$��h�V�7i,"��5^�z>=t(��ݰUl����N���U[����ffff/V�V��󙙙���ZU[��������z���wwy��Μ,��0�<&'�<C�:p�oq/�L�`��+-�Ƣ�����mQ�rdwC��3�!MG`��s[���� B��)�>i�����Ex�.pd"n�PY �%i��D�M׻h�pD4�LE��uF�5G�9&�MB���*�D�rN*�CN��5�T5�f�n��Y��u%�L�3&A1�����&������ξ���Vw|t�N����)��^n���^��#�M���	�s�9ڤ�t������"EL0!��u����Q��
.��<t�]6�g*B���M��$���$�����ot�hn6
2;Y��رM�kJy��x;
��	:�pgL�"��<og�J�.A�;�e�U��H}[���+�Дךɏ�&c�<�:�ϔ�:��<�o,����
&I�dv;UUR��-��h��cd^���<�A��09޹��G�&��šH��a�����;�xc���\��<g��߾)]d��n���N-��ޏ���L�	��7p���$�i>�y�ğ�;C�~?=˝<2[��0<f	în�'�p���ߛ~Z�Z�[�yky֔�tN:W�FJe�PcRU0�o����t{�I4��p����M���$3t��/�n�S��J�*���s�xyr�2o�>8'8����XZ�Ŧ�4a�$՚ݑQV�uH�6��ݯt`��|}����	@�b�^=yyϱGY5��m&á��F��Ƈ#��KG{�	
ct������[2H9r��|X���6�6ˋeO�S�:�����:t�D�<�"eݒ^�UZtӗA��:a��)61�����2h�H��Q2�"Q"F��i�2��ٟ^���F�&�lsy��<�g�,.i�����lI2C�e�D	��&��6TK�K<h0Q�y�Jv��k'�w�r:v�83��R�FHL�̋���K��e�ؘ�`.eB@�$���M��h�R�)n��<���JR)�\s:*؛�?\\֫C�r��n���C)�&*�r��,�]o��rQ��V�6�(ݙ%{`ʘ����/y"�+ℓ���:)+�jڪI=q�GF2,-�T�J���m��x3��vx~G7�����&Yni�7\�4�1쬵K�^�|�%̃��d�㭏4`v����r�:,L�J)(�t��p��Ft��bI�?��	1�LH��DLi���ѵ�����,�gqnD��Ne�t��?<���o�z����"�Yi��BG�/�s��2E(��L�X��1�u��8��yռ����iJE2��u33Z�#ibBsW�UV����Y�C+4	���}�&�"�/�N�J���.HI�+�v��Z�D�����q/�d���x�Q��|v�Д�P���!R�0۷#�a��ɟ�Х�و8s�pB�ʄ�+[��Z��!p��M�}t�0uK�;�-��k-�(�딠�q�pǌw��b��>[��)מS�>y�Tt�D���%C�D������r6Y�F�d�L<()�`�ָ;lw!�T��	!�pN�IFx�h��x?���ڣ����VLlicI�b���	�u	�n��<p�Ɍ�*��
�\��p�s�9T��L��'��O���6��wƅj�ӁÀс�ʁ��J��>y��y�έ�<��eJE2�̋�����hD�1��7{�6۪�J2�h��`C�ح	`��/l�c��[��Ȓi1�IK�e�42�N4;c���]r�7<lu��L�01���`�fϜF�7c��\(���<��|��g�V1O��v�m&�t�p���7��9��͝Ɯ���Ɩ��[��S�)n���e��̯��7��pe���"�m�eV7�7�|6��N<4��.vJc�aA�2q\��!���b!DIJ
�؝Ӟq�W�I�=��q�V%��A�RcJG���,��*�אrIve�%�~I�CZ϶zj�'?a$$�4�M�N>i�T_E��`��o�aA���^������^{ ��~Յo�p,��������\�
)����7hʢ��;0;�d�$�6���j�\��D�#V�����w�$G��:1�0�3�h ��w_:��ileN�>yN���)���<#�:pD��j�<�����&�UUZ�_��W��g��B&�BCsH{r�8gX}�����l2�]���2y��z>�A��"X,5��%Q��=�C�p8p-��Z���Pp¹HY~y�Y��.[#�F,�h|9A��$5R�9$��.S�ǥB�rHBt�Y���-�<�i�ξu�<���P��xDD��:YB$b"'DN��Љb �<'؛blК"A6""tD�H"&�D���<��,M��L�i&�ДA���<	� �8l�e��:'HYbY��L0ن"xN� �D؈�0�Řaf�0AAD���"hJ��nS{w��j��n��W7K�=�yf�d�4������5,�ߨD�4s�O��j�E���>�{ϣ�aݨ⣺�sY���<|.����>�9�^�gy{��i�;�s�o��u��mzZ�3�?�����u�z~�o#��]�M�{�Z��g+g�ܭn�﵋�[�wu��.vW�W�T��g>��/���{ϥE˾��ﳓ]�[�����>��w�V���33333�U[��������_1Un��������|�U���s'�-�qխռ��R�E)ˮ<V�j��)kU�k�+��Ew��a���l��ƞ�$߱��Z|��ć�"���%X��B�d9�	^��2a���!�A�]�
��<1æ<t��������W�̓��,�J2l=�����~u��|�_<��S�QJ!��6�[�^�\��RV\󞪪�_+h4$�������
�v����)��¦�J��6� ����V4�φL�	�7��+ye���K
s�ᤰqՇ�B�wM���~���#�ϸd�4��L,z9䃰���%�*�φ��E�Z���S�)�"��q;�v�_Q#tn�팒��M6Z��Ar��fFɑ���F�CS[�%�)�:l �CV$)��bT�d�<�v��+-�)E�XХ��z��m����e�t[��L�.r�Ã�ȫ��C�P���'r[x߹�ø�{En��%�E;�s��qa�6�w����4�73�O.��^�m춁��]�'U�Ά�O��yF��+xz]l/�Ȕ_^�
���C���&�@�/��c"4t�!��%Q��"�Eu���l�'��?c�K,�ئcks"ߟ)������[��!��6{�!�&A3�z��ѭL*圻�t*$�����z��MV����Y\��r����A�tm�Vd�>��N�c�:P���bRH�!c�)���7?`i�r���q��c��UF	U�c�Tn4�K>mZ�|8��1��/�|��<�<��R�E)<&˻���I$&E�f�UZ�x����q�p��cq���'6�`�jT��}M����铇�8��$�����*�b�8���V�Q� ���� �x�Q;�Jl]��������B�*�����GA��K�=�׬f����8.w�Ħ���M=�'a�f�iO9�u�:����u��y�>u�!��6`xB�$�*��j�ep��jp�1��`��?�D�s8�������A�7�¤�D�V*X9bNx��zs��XwÖ��C�!����d/oci&\4l:��g��>p�P����$�t�*h��m�8p�X��c�y�2ۮ8����<�:�R)���o?(�K�P��	��+$U!�� �*�����Ү������ApDa(��a��LF�E\}5�|Q!�팏VEY*GmU����#�bwlq�8PS�UUh�\9�<�a�kI~���C[�;��"�����y݃��[�9'N��/��DUkj�;�CZ$$9u�Jc4r�ۅ�zi�֛�i����+̄��B��ӽ焝h6��'n�S鐜��FH�M�C�v��^y��DH-A��h�H4D*����Ж�H3��8g�|���8�иڄ6����Ŏ�<��y�<�:�R)���1����;UUh�
���*�UZ%F��6�s8t9���i�3�y��g��ܙ����'�G!bL���zl)���1��:M	���Ux�j�EGIL���n���̖������X��:wߌ�+�D��h��
��V��M"�E�_|Hѣ�>R�S�<��R�E)�S�VN���#(�<UUh�\�*j�gB�E�a���k�74�/nɒ�wŃW����r��gL��'aҋZ��,�!L���D�����q�J��<SA�v91�\0t7i�9{L����	<h����N��������;��[�y�o�|�V�yKu�S=Fg�&2R~�jgPn6�̷j��	d���`v��Go���ф����ܹ(�����A�@�4%mQD2T�(&��Be�Ӝ;:j̵�`.æX�ns���?����?��FRhf=�Ȋb3�c���M�?u?1|�y1I�Ac<��E���zŪ�kI6�Gg�o/���8�y���O)׉�<'��<tN�P��"lDDDN� �%����b'D�8lM��E"A��"A��D���<'�6&��6hM�Dd>C���ADxM�(��D�,؛0�	�Y���"A6""tO��8a�4```` �"%	||S���>��)KTi�_����ԗ8;#E�d���a+J&��E�`����x�F���$Z1�m�E��q���s�|�)�UtI7�2uũ�Fi�ƒ���-�RD/��f�:��q\+d,T���l�^�KP�6�Z�*�W�8����'>y��SH�j�@��B?R���u�ɡ � ЙM���L޳�B�gr��	�N�;���h�zmD}.���7�E�4��2�e4�H�B��#g4�6��Q@�<g�-,m,�FY	J�BX��E!<����G�
%�⧡�`�.<E��d5e
,�!��%�!��y�J-�s�8r���[�����ٸ����Bs�1�V�G�/9�Y���%N֚�BH��u�l�R&�ZZ�T�:�r4�Q����R*[T�J�P�d���`܂d��BH1J!�j��uLHD��T�rԒ���Dj�"!��k���$I���
�� �H֓M�&Dᬂx��H䆱�ˏ��o���'fJ�ժ�R6A6A�lU�V��Cs߫��^����EU���L�����EU���s33331QUn���33333U[����:p�ӧNa���R�E)�O��L�OD�Y�o:52�BF�h��k��F��d+."��"��ꨥ��A!����I�6*̍�h�$�1,�m��6X��5\��,ԸA�tF���%�*��2>m�����ġdjX�LX�R:)TuJG	U|�ro=��4���tV���j�Lv�z�S��UV�n��S����O�b���Cu�!s,����u�\����4�B���醭͟������; %l���׆@���!�y�@0x\�M��R��	C��f���-ia��:Gc%U�B��\?����o|�3!�7�PJ�Q&����0�T����<�:�R)֙�"�E Ʋ[1km$���X.S�H�Y��d4� ����|���0{�c��{zoĪ�����e�/I8��i�*��t�i3
B�LyE���,��Ҷ���*Z���������G!��P�k�I�`�ظ����ɏ�e���y�_<��S�QJE:Ӹ���ա��$�6�	g�݉E�96�z컢�vI��`p9&dI����r�g�.|�?5ԚO�H�=O���
��0fI�P4��_=n���\��8˰�7�Dˆt:d2r��ȼ�d229n9=�~b8�O�)ż��S�)Ŕ�<t��@��RI,?��Ǆ<��hLI/P���2/�d��-%yki4���٢�6�H���xϲ�N᳋�,9=���������	F��Cm�*��6Q$�l.�xrӵ��HBJ�2�#a��<�$|e��I3���}1"�����c0�F�OϞy���yO><p�<#�H?t�ľx�(�F�Q����wV��ٲ9=%�N-t�TBk "#Td�J2	f��҈㕁0[��IP�͹!u�-DUCI+&H!`�[#rwu$��MJ�I$��9�;�>=�l��]�qvn�zqsoy̛��H�ӵT��mҊ�<hl��a���HHhr`�Y�����/C��	��%[CO9l�<	����W06/mh/M�s&K�8��4��g����//��#	$H����O�d>>`$J}�zIZC�I���Ō4d�[�y�8���u���왉�nI$Jh8ӗc��𒓎Zr��cTWN��ŉ0l�2<-�N6�$as.D�AAô���d�<݉���N,�E�� "�����������Z ���ħpi:���5Xn���L�1��8{đx���揟?:��y��)���<#�I����u���k�WRRD�N��=a��iu�L;�C�!p������{�<�3C���ΰ�&N�9�"��#_ăl�q�ɻ��qg���Q�A�~:f��M�����BG��d�}��j2�� F��$�'|i�������Ι��P?g�̔�B��8�:����qe)�J㩘ra�54�I����$��4�������$L�?�@���j��QTcU�"E-bq��	�L�z0���s]rT'[#�B�����v:0c�K����t�᧹�xv�p�T&���x9�d�T�h��#�I�25	Ғ����!�	��9)�1�Q���iNBE�S���?<�ߖ��uo)���P� ��6G�rR��uA�6UZ���:�Nc�L�P�)�G8\�!��1*�8�E����"
6!2e���Ǝ^UĝK
�B�t�(�LNKR��(�V��*�"\�I%�����'+\���dg�f�=������p��H�%mK8.MP��4�HD�X�]ʱ#aq�kZ:��M2�ō���nHdzqt����X68;�USD)�oc��R:������3^�����#�:S����Ք?-Y��KD��P�'�R��U��f�.�^��pz���x댩����yO<�R����{!զR�Ky�$���VB�9"BE�؄)��jU��B�tΚdj������N���p6h�%;)��C�xtQ����a�w���Ү����a+H�ʒy���Hr��Xh,�OD�
���h;�/"R�BN��GL�eCg!C�B0ˣ��hՉ48|X����x8`�֧��|��<���S�yBxDD��:YB"P��<'H ���M��bxO�ӢpK6lM�d� ��b"'��B"5"lnDG�'��%��6hD�BY�4A���8$!��'H�,K!�Bi�R�kZߖ����e��<P��"tD���:X�%�l4Ye�Ye��<�O4פ�m?D��!y��|��h�����	��9v.��~����~�|��]��t�|䫿{�
wz�c��N5�����{�w�ŔI|��Ov�|_���r���۱M���o�׼|��o7^�����=�y:�IX�����6�u[�-�]�������(w�O��}]���˒?יvqw�8��|o�����;�{��/5o�w�l�}_%/����|Y���ʺ�z�����G��y��E���q}��ي*���ڹ�������wwv�fffff"���ݮ33333Un���g8p�Â'O<��S�)H�ZkrI&�d�YL �Y�3�AN� �DH>����}�C&tLA�9�J�q����$&�c#u3�C�bώ��B�u���A���%87�	!0`�J#UXhr�l�d��-��<���\s��o<�����qe)�GD���I0�4�?H3��%ْ�I�a��Q�L�V��O���Z��ݭ'�ĲB)y�ų�).)����vw���`����]�Ɯ���yӣC���p|h�Ȧ�::4�cDD�bV�:D?V=����	��e��$4b&�ٚ�������ƵR�b�,ˈM��e�o�m����u��y�8��"�i����}�崚�DNAJ;+�K,X��A�Y��5]+�� �Waؐ�I���]��44q�׋�!cz#l#nۉ��!��$�ӑ9h�+C��%aԒK-�����㜧x>v����9T͋�u���3Uk���ʹ@��w�������|d*�GnY���W<`0����x��dlg���=D���v�q��86|��GP�P����d	���8g�fS8��\/�e��D��$ZY)(�n(�N2��FD�p��O؈�I�፫y��-O8�:����qe)�X��&33��9TQ*C�I�<,4l}`���$N6nRp�,e��\+R+"� 1�;A$�|�4���x�������aH|*�·�X��a�l��}VyXH���\,C���m�,����(�4Ş��ܠ�&��V�xA����+g���n���Jx>�����ή"ag�b���n���8�:����qe)�O��cR5���.\5�9�$��k�n�>�:���H=:a6di߃����z`��M�0:8e�_$!����G��v��MB�(�&f�韲�30�SE��v�_ewpI�t�����,kE���:IPl��Ѱ�Q�:�kR���y�<�|R���Əb=&�D�A��I$w�I��$ �aI��Ig#��� S��~�p\7��S�51�i������r�LjM2ۖ���E�{����G'�	Fu*�;��hr������! ��vB��:a^�H7R+G��9���"x����k�����#q�rД6,Xn�0��A�\���a+GI���J|��q�[�y�Ie:��ҙ�}$}rǍD������F��cz�ku�ep��%1,53q"-���1GX�����r6V؉h"����\uD�b�)dVVU�m��|�Ie��;�ʮ��uq�K�o��Nu�o/������ը��Ǿ��ܩF�!�8:��a�b�@�zT����CO�!c��	$!TUT���uB��ܲ��7;^	Q�rCp�N�D�T8U�����-E�EDC���<�����9��mEx�2!��J&��ۊ�8ft�,���\[�>q�[�yן�:�dK3Y	b ��$"2$T�Q��L22oFZ�Rur�3sI���'*�����5�r>
B�
jL�MĄ��p��KO��I����PbB!�(4G���$6�����.�G�=E���[�$6t��0lec��
%UVΛ7��7���:���:�S�<��ye:��j�=�#	�y�$���������s�6Jn�n4X�$�
�]�B^2������q�C)�<�`��f�`���S��5W*Æ�Ə=�[#G��+���X.�4a��*92C�~�Ԝc�^G<���R$"b&!�&���~c�Skq����I�<�����:p�8ۉ�H�<�q�RRG!@���bч�G&�~�x~��~q��&"
��j2�JˇSg�L�|�l��fàs#�t��&Nu�s�%�Ga$�y��^���v�h����*<�M]�<&́mu����D�$6���f_�/���$�R��UR�Ti�m���������?y[a�g젓���kt�DQ�A'�ݽ��_E�\�q�����G�c�-,KI���I��M5��E&�D�$��KKD�F�M���h�-"ZZM6�M�MF�ZZM��M,�E�i�%����ii%�l��-,�E�i�$��DѢI4DM2I��&�$�4D�I�#M"I4DML�i�8�4h�h�KKH�$��4��%��&�HKK"KKG��ۢIiiKKiL�IidMK$�$��MM,��L��3�KH�ZZD��-"$ZZD��$��$��L�Y&�I��I--2$�KI���i���p���%�idkKH�I��id�Π�ZZD�im&�d�I$��I��$$�H�I,�I2i$$���RI2i	$�I!$ɤI�KI$�I	���ZD��4�4Ȗ�-$�Id�$�ZD�I	d��!$��	$�$��ۄ�Y!$�Y$�D�I��$�I-�%�%�KM	!$�D�ZY"Y2K$���I�I�I%�i$$I��%��h�i%��I&�&�ZI��M$�I4��F�H�D���8�I&�Z,�Kh�i%����4�M$ZY"d��M-$����4�Y&�Z,�$�D�I-$�I��MZI4��ZIh��DL�4�i"��$����KI"H�i$�%�i$Ii%���D��,��ZY"Ii&ZM$��D��I�IidM�BI��"H���L���i$�I�#DD[M�""ZD�M�&���n0��B͡3Ba�mhC!l�F�4,�cB�BcB��d,���	�B��#mfжd&4&"�;u����V�:�s6B1m�3!f�Y�FІ�mlG�2�&�X�FЁ	�d!A6C��7FB6����f��B̂�h[hY�����m�� ���ж!г!6��, �!1m!fBLB�d# �И���[������7Y7�㛂h$-Y��E�Ј�M�h�-&�l帪�ZBE�E�D�YD�4H�hMȚ5�E��hւh�$H�$B$YF�$B$H�Y!F�-��dMD�h�D�D�D������dH�Dk4DZ"!,���V�MD�D��"h"&���"""ѡ�DD�""����"��H�h����DD��!���"��DD"D"4DB4"D""h�B!!"h��"��i���"h�h�-g&9��&��"h�4HЉ�Ț$Z!	��i�dH�Z"5��$Z-D��D"�d-&�F�E��D$Z-A"ȴMdM4�d&�"h�&��F��4H�YD�E�MHZ7]p:�B�D��H�HZY�Бh�h�,E�4i�h�&�"�h�&�Ј��DD�Ah���-A4&��h�D,�4$ME�Ј������B"Ah�"$&�rr.�Р�i�&��h�E�M	�&�4i�&F�BhH&�Ѧ��H�4Ѧ��-Bh&��F�FM�Ѧ�;�t�h�DѦ��4Ѧ�Ѧ�h�&��Z-дe��kFZ��і�h�kCM�4i���4-Bѭ	�Y�9�0�B!4-4ЈM�4	��h�4-�BhDi�Җ���4D�4w�8M6���Z-F��4ZkF�&��4kM4[D�� ;ۢ�Gد�Z��Br?�|�������1��6T��f���1_W�����y�w�,�i�|�.D��7?O��Ϳ8O���u����1��7����-9�˙��7_����|��s�~������>-����#�n����?O��y�?u�|�U@���r������F~�1�������ߋb��~~C}뿿�ϱ���|�%.b������'���"~�����ꊠ;�E?�?���H?j�����Ж���D[3�?]b���7�?��II�S���F������ܧg�P��|��X%�i@?���׎�?Lm����|lXQK ���?8�������0"
�"(?���0 E6�8Zf��(��*��M�G고���(��L/�|G&���1�Q&Ϥr%��h��Q#cmD�AYR[�~F�$����Z�8����#�:�J".ߢ��=��<�U�?Q��c��ğR��?g���뗛s�T��h�,��`>u�@6����w�����|�������?���# ~t���)q�"A���O�����߄��G�g�?����~�b3���z����������:xl?F@�|G�nϹ�@������?a��b~2����9C������u���t?񰍋��W�P" �p���{��]�0��g�TAi���}�aL#��KJ+A)(��%4}�f�-�E�e�����6�r�u�p��Bv��UP\������_�g��ʢ���&��F~���}�O�������k��}� �L��d�7�>�T����i~��~ˣ?��"��(�H�����c�|����TU�����&>�_{���/��Ejڵ
�)���B�[SR�L��V�L��X�
Պ�+������5eej���j���Օ���+++SVQEej�Օ��ը�[VQYMZ�յjڵ
V��YYEeb������V��B�mZ�+(�[VQYEe�jՔV�ի�YEmJ�VQYE2�
V�V+emX�V(S+)��b�X���m���+el(V+jeb���B�MY[)���eb�V��c+�5b�F���m[V�X����Z��l�Ejjղ�2�Օ���E�V���V�(���ڶՊj++)�+���6�L�VS+S+
jڶ��jjիV�j�ի(��YEj�+�իR��j+QMY[(�V��Q������j�Պڶ��ڶ�)�mE��jjجV(+�
�b�����V+j�aEb�X�V)���S(V+�Պ�b�X�V+��b���b�X�V+��b���b�Y�R�Q�j�jjQM�+�Z�j��Ee�S+Vի++VԦQ[V���QMJj�Պ�e)����Z�eb�jSP�Jj++Q[QYE5e)�P��Օ�VV��MZ���ՔP�2�V���������������eeemYYE+++j����VVVVQYYYYZ�j�����5mYYB�mZ�Vթ[V���ڊjS(���mYF��(Q�P��+l���B��
յf�����EmB�B�L�����5
eeej�e�������mYEj�Z�V(�P���P���5����՚���PV�R���YEb�AX�PQ���b�X�Sj��b�X�V(+��b�F�V+��b�X�V+��b�X��+��b�X�V+��1JԣV��+jQ�+e+��2����J�)��J��J5(R�VՔVԬ����)�Vء�YJ)�jQYEe�յ(R�R����+Q[VՔ�J�)B��j�VVVVVVVV����+++j����YYYYYYYJ�j�VԬ����YY[
(SVR�lVՕ�VVV��YZ��b���YZ��ej�j(�[P��Vj�(V�S|���?3Ο��'�DE�(�����e>��������8��X��H���(��l}(��� ���Z�"�|G�6����$_�~<?���J�wC~���c�m�n��~�¢�S������d�ALO����?!��Keo�+�?o�?g���������~���VPlO���6:T����?a � ��b?�ߐ�0�#�O���>/��	�'ԅҹp�*\��9�i>��u�`�����_���T����O��9����)�m��