BZh91AY&SY���?�y_�`q����� ����bG{�        ����fMT���WVlli�i�mb"ٶ�ز��V�Vmi�6v�v�(�Tpm���M��m�m�lm�6hƤ͌Z�  ��{ږ�i�ԲER����Fڍ�j6L��;[U56:�i��F����u.�Gl���V�v�����V�wn��lm�m�2 iZU2Ѿ��X�d��q����1n;�6���tg��ɭ�1R�\������/b.�Ff��]u+el��cj�j�7�u��C^#U)=�孵��[F��S�ݚ�U���  <h)��P�=�=wS�:�{����C���z�yWn�{��wN�9�{��{AԻ�ޭ��ިun�hi��1�A���íEC�
��u駓���ٸ��FF�����_r�4�*�ϴQ
6}\� � ���((v�8����J R��۩�@���*  =뽞C�Ψ�FЪI`����_^������Uj�C+0m�,����z�=�  );��:J�ު���K��dP }�l��|P>������ ((�]�O������o���iL���>�4=�p z��h�Y�����V�2�ހ����|4�Uz�_O_=� >����/�hi��y�uQ�����@}h+���ڪ}�{ק�_�T��>x z�_^:󇧠�Y��P�����b��Q��T�[5kl�   �{��h����}��������ݾ�B�����@v�wվ}�^���
��>�O�����B��������B���ʈ�c���{C�T���k�Y�f�f�X�m/vK���  V�� .�o{Ӈ�@	�_g�4)�ϻ[q_@oa���>�� \���Ф�z�.�x  S�s�����ox�U):��=�O�]��2�Z��a:�]�� T�9(S�Aj���{4> ��Oo=�������=G�0 e{���/+���(ggt Wќ��
�oI�V���Z��B��mm.�   ޾
 -R���;8u�(������� �\ �v��@{v�� m��\����k�� �Fmz9�۶�M�n�JVգ� � =��t��h<��@P=�{xzL *�]n��J�����==&�g ի� 4rukO���ж�e\��j��| ��m� Gw�ժ���� 
/u8�I� ;�p
 �ќ@]�qT .���6��� (�      �*R� ��0�&�A���{FR��h�F�212h�1���%*��@     ��R��i�@    �� %*��4� �h  ��L�I4&Ќ��6��I➓�����h�?����R���#�S�{�{��>���ߗ�=��¨ ���_::�8����(����@@U�h��#���g�����?�����A���1PV������PW���&��?� ��������?����_�9�}d?����02Y|d<`<e�����x����~�x˙O|`<`���.`<`<a<e�����&�|e���|f`��_|e��|n0�����0������2��������/��020�3��|`<a���_����|`<e������ό�O|`<`<d<e���e�����C�C���,�x�����002���3x�0��x�x�x��/��2�����/����0����/��3�<`<`<d<`<e<e>�0�1�O|`<e����/�q��_|`<e�_|e��_;g��C��������������/|e���O02��x�x�x�|c�C��C�S�_N�|`<d<d<e��x�x�f|dOC�#�*L�0�x�!�*�(0xȡ�*��0� <eT�G�OD<eP�C�TO<dP��� ��
2�x�	�C�O<d�G��ʯ���2�0
0�x���"����2��2x�	� ���@<`D��A:a|aP�S�>0(x�!�"��0�x�� l�0�x�P<aD�S�T<`��AI��<a�C�P<`�#�*��0�x���� 'l2(xʁ�"�l*0x�� ���0����2�x�)� '�POP<e�C�Q|`_�(��	��"2(x�!� �"����2)� xȯ��` �_<e��@O<`�OBe@�_E�_Q����D<dW����0�xȯ�*���l��/���ȯ����	� ��'��2+�|aS�_|a��|d��O��0���/��2���/��02����x��'|d��_|d<d<d����C�_|e���fO~2��x���!�	�/����_|`<a����_|a��x�x�x�����2���/�>2���3>00�����	���2���'��3�<d�<a��<a��_<e��N�<`<a���/��2���/��2��Y|a̾02���/��02���$ό��>220�|���iߞ�r��������K�w���?����cmP�N`�{!z�a1�K��X7�yq#qÍF��,��ǙYa�Q]�OHw��3��Yd}AW����
���݋dTwU���Y��neZ ������c�cLQ5b���b?�uu�m�a^T�yY#e��݆C�o(����ݠ[:�ϭT\=כ�\0Mf:qd��1e�K(����T��]h��[K>[�h���ᤥ���4�t����e���Kc��U������M��9�]�!�8ۆb7[�����y.&��$�ݺ��͖�`8���n��C�f��4M٥Ȱ�1n�h���H���%)C5 ����(�R�EY%�@�鱊�yn�F���Pp#KS�m��jQ�l�n�d��g+hB����h���g)��6	���. ޲܊�-
K� ;G�f���Bm�1�N��kXE(L��]�B��[��9��lH6���w"�{iʽ�T�B���zʎ���1b���n�-��C���h�1�f�7a{Xճ���J�XyݓE�i��$8�J��o&Ҭf�Kin���f�*ɔCj�vXN�͂���
n��W�c���M��I�[���ܼ����4St툵���)Z��4����5�5��/P��h��]0d�Q��
[ܗ���oת�Ә����a�r ��D��b4�]n`Ñ�R`0r��('�3�k�E)k&dZ�[�xê{w����<�v�V�n�Scgc��TK������ì��vJ3wlʻ���d5��f��v�N�4�*�s��ի� ܭ5��m
ؠۨ4�7*�!V���ZR��3V)���G5扨iO%k�tuh6��&f
�q���V5<֙��mY�M��\�C����#�4�C#��Ł��S��0��S�k(�S� �o�ycwpFe�[E6���cjP]m��);X�Mպ��m@H��6(��ۨ`�1������푺T����.	u��ݹ4���"fZ9J� ��N�II�JS��h�_JS1��\�ܵ�rWRν�9c9 ����!��v��v�����0e��a_\р6]۬�ێ�e��0�&�i*J�	|j��*�cR�+zK��5P���a�!��,��6eL����b.�Q#D*5T-�s��QOQF�E`�t+B�5
�l����4�ۼ�H!Ư ��j��i�oMn���oj��@M����I3F=�v���
w��70st`[o���\U=���KM/HVT�m�؋o���zebw�U�b&	�-��N�{�ur�P�QsǏ��ҀF�y���D��B�N���4nY�͹}�ñ�w����VM�������Y�R/-< �Wv �͉�l���U;̙S벖S�u�9�Q)���{r�gt ��]#w�h�I�û��6�5��͔�m����WQ5�.�{��n�+��v�)+(�^䬺;6��,2b���z��!-�R�ᕆ�Y?R؍6E�v�V�����TDZ�R�ͱ�m�:� �/!���|���&AJ�cv-�Ћ��Y�qJ�ΣMjJe8@h��V-�ĭ��: ��aA,4\�E)�˼wXY�SP�olL��a�D��h+���Z/i�u//s F�1<R�j�m$��a�4�b�;�5P͎��X��Em��#t�*;�A��&Ck6�ķnB���kPqf���.)b�-��!ssP7b]t���í9j�4�c5�D��)�0L�؛`�
�ݽjV�Q�P+)��Y ]P�`� /$oI̺k1j1�Qn^ձ�e�A���Q�z�4�7���l�m�ȗ, `��j^|J��]��a��h���KM�B<%Z�� Ǆ����Ճ�j	h�B��&a
:E�$�m���z�LV�wNL�̆�wb���V	1���Z��l+�4h4�<����`���ur�uZ��km��e�I:n�Q<n0٠0k��]H4F��K�nh��$�ia��(\/KAԵ���,W՛��e�.ڂB�v�E�N���u>Yx��/2Im3t�wu��q6S��ۦ��5�2�#�n�0Ek
�&��r�<95��/H5+TZ�n���	L��75�f�蠭�1�׻��2����޷�Bd��e,{����u��g�a���@�z���,��
��p��x+b8�ȍiE�D�D�g%3.l�Z�2��bk�ԬU���e/�{�6�r��@�E+6��Q]⭎hFsE���[�N��i�`X���i�WWt�V/O�fm�(K.��rY4tMEৃv��_G�p=�Q����K��oB��$�l��8��6� ���BA0C7��UL`%gL���:[1�`���yFR,�XisE̘�:ZK!�@C��>�&/6���J~G2a���R(���R�4�����޹R����Q�Q�D�F�0�
4��6�}����;�h;7���W�'�k���*��2+ʱF�ٔ�]lm�^|nFf��]��)yt��d�J�z��������e<䠞�Q
A4M�[���rY�X�V,#��q�77��$�.�v�ȹ3Te�733嬭@�(nֻjj�X�ӕ	�6nf`Ѱm�{$t�m&M���IZ�9Fu
v��x�۽G5�D˷�7#֭���C�۵�@�qd/L�Ǥ�8� YWZ�ԛ��ZN 
Q�"��K=���lXn��#��-Kcj��LM�B;R:�o�6��gTN����15��U�&�e[I��5�f,�����Y!ƞMh5jU�� �AdT��0'r�&	�6�L��4�^U�*Εx�Q�y��AF��bMTο��\�3V��cb1�r����1�u1`C��kN���%["��ȍơ�X�Ԉf��(`z�V�����d׬�ZBQVa"��2�"�lۥV.�d�s7ɒ��&a���m�Zc�-���e�ceTj�=jiR�ѻqn�b�6�hcbB̰en�nm>b=�]jVjo����/f]�[�.�f����tX����XC���`(U�2��Z]�lT�Fb:�5@��a�
��nL,�Gv�m�ZU^�6�����ou�j!�4�nU�]�D�M�����v�����3p�e�EVZ��ّK�f#7l)��*��ҽ6RN�8�NK��D�aՅBc��Xfbf��M{�-�u�B&�d���mY�Y���M�r�{aM"�����'Jxf���hf�x�kcn�-����\�*�Xo
�P� ��@7� 	sq�!nI$�U�r^�ED�2��)��ӑ2)�^�A��I��p�v�B��ce�X�V؈(,G[���X�ۿ��nTa��l��<�B�)�.��6�AkPݷZ�iјX�)�0i���Z�U�*;×3&G��@]��*ō�x��0��$Ŧ6��V�$�[D��M�p���Ev�:n��}�8�/v<�E��pLDW��r^����pQ�-�x��wL-��v��M�#�4�TӘ�	�¨s9��qe�M�+� u��5'�:i8а�� �;���$w��2�n�ա���y�]ȭ�iŭ��cYF�n�7��oUsKin��('1Ϛ���dդP�NSz�ֻjZ�l���#-�(\��Imb�q}�93�N��B���Km����q�{l1Vнj����Y�W�$x�V�S]�&)��É�g)����5R
�(Խ�h��i^du,I[�fը�y5魤Tw4��[`��QQk�-լ�`�8(F�Smb���Ȭ�Dx�G�3Z-nY[�rF�p$�JPw�9C޲�0�XU�<�e��j®ب�[J�3:ugl�&�	&cڷ6
��ə#���M�8�H��w��]-�Q�qn]��VE-�t1تV�1�&��K� ��q��ق��ġ�g	*G�&bf��V7XE5PXz㷖f^���J��MէFk���h	�Rŉf	4�����A����F�ֺ�%���3��p�܍��&K�&d֜��ɀ�N�M��M邶۩t���=v�fn�D�ӻ�
*'�[џZ�j��U�����٬a�j8NXĨ�9 ��>��$��E��^������A�YI�Z-�d��̬�BF��%AHDI�FP�Ԙ7n����#��!R�V�C�J*�c�e6S��m\6�d�_-HC�F�Z�^b�V2%,�����<�7m	�Q��I�)��%X��lKQ�T�w��W��ݚ233iS� ���J��7j��6��Vұ��on��U�i�o�U/t���*�ķj�U��d2��m�����\�ʴih;E���G2D�J&�;���Ǵ)�6�"������C�C��ݨ�U!.����"�$Vݼ�T)�Y*9 ��E�͍��m����X���˸�ع�atL����%ޣ[���&�F��n����Ȋ-t3a�
9�>�=F?����VQ��t�q�b�Ӣ����o
Hޣ���u���h�IKi���h�{N��J5�7��� ��0a�����o3.�YR�yeQf,J��w������X5iR$4����˔Dx �A��2nȩ������&���=QJQ�!A}�(�ɻU�ָ-B:�����G5����X$a+Rl��6�4�j�œPǨ�+iA��u�l�.�2V֜�4����T�67���A�6�f<Vn�P�J�?��&��*up�h��iT�س�ۡ+2D.�՘�H��a#:�6TonC�H_Z;F�����ͽ.<YHӃ)9��0Άp�O3��e�Sc,_�XܬQJQ��Ť�ޙ��Q��պ�1�^��[t��W�Ld䨦^]Mv��Uc@�-����ϭ�H�m���Y���~J��d��]�ճDe�(V4�x��&:W�o2m5��v�фJ̚5���;ۢAB�8�a;	e��Of��oh���Q�MQ-xFPP`9�X��t�%�7&��:�`f� ��3�nn�Ѕ��v�+Z�7y;�F����"4)���Y�1�7,�Éէ�ZcJ�/!�J�0G��D*UG5��i��"�"�J�0)%�r�6h��G�������Rj�n�'K]m�@�E
6���RO�Y��n*W���694��cE����K6�-#�s$��@�f$�JNڬ��"D�,M����:T��R�'��)��9oj�ƞj����7��we�v�E`�hG3)���l�-�y��D4^@���h`��X�
�G&�a*�
�,:��r٪�jFJ�Pۗy�$��%��ۗOim�{��1��d�פ<���L`1Xh�0�*=���na�7��$�5��v�ke�ː�d	e�j5����z3\644�ٲF�{[$�mk�6R�ˈ]�Q���[�%J8�VrjU2ܻD�Һe����gb���6�S�m(Q�����gw1�J�NK� ;�1��E�����`n��i��à0���l1ȋ�`�.��,�BAuD�kz�U]�ɺ6��N��P���-�GCȥ�?m��VRekTеF>2�d3@b3�c{H�g@x�"B�&�,[��
�0j��W���L�W׆d�,�J����"f��sRz�i�C��%Bw@M��pVa(&���� �C_׵���i�V��fǬB6aԊ�F�q�	�S�A�v�|kE�g�m��j��=�*�؊�[Zf���F���5��]�[��A)+v�44X'[u���-a�3`�ʴe��<��e4��/^��(�`&�1�x��S˔d��!ک4���-٘����2A#�ZN��3�QU\����f�c�Z�U�)��lzѕ�%A�'��f�,�yI�CUJV@�Y���T"w��A���Eޭ����o6�Z�\ĵ�ȫ3 4h�E�	Yn��R6�5�F�ӑn݉&��N���X�7B�(���qB[xD̽G+tem��f�3��cQU�#qi��n�V�`��b�fl:�
��s)cb�i���?�YlM�(̗%,bi�M�۬VN�Sd,� ����i�P%������e�<�c+2�F����e���¡�ځ���Xzn�@�˨�(ML�,`U3�G��F��f�b�x>ͣ(@L��ա ��i�2�R��V�1{L�+�F��N\�z[�R��ȼi�5�T�ܫ�0�Ț2U�'#�J	0+�Ԫ'G��td�M��	f�,�9�L'<^3�fP�� �$&�ʇ��<������_��W  w[z��د����}�V&;2�a��d�2X �Hk���B�3�c�rW,�AIVs'�p��4�&G
hvM��☃�{E��0��e93���K�tvz���VP��
�r0�WGBl$��.��1��\X\)��p��tX �uGK��=��g���ɾ)�dxf��
�Xk=�����2�g�f/t�9�
��/ad��W��h;*�Cp�)���B(!�p�&��d0�,l\]�&��,�*
$�8H5����R6u�f�з�IxM�C�Y�([�Ш�T�;�$�=�٬�@��v6pv�'���5�)��p�*ΡhX�,'J���^%1��!<.Gf��(
%�p��aA��('�"a �Y�A|{ =Eజ$�����xL+����*�b����.L��p�1��f�S��*7.|N�	s5F
�8*:�����ql��%�y�P������l����,.����sZ\�D��H]�f`S=H���t67f��(f�l(C,Z[ ����/K��x
���H�L�.����VK6f*��
Y���m/b��/��vOq�`y�pB���V).2�r�K7E�p��0�[
aT�����/I�L��a�O��kR�����0���g������'�����à�.	\�e`�M-/�$�\�j���Kj9�� a�b��^fЎ7���bƨí����0��#mv���얪e����t�w�H�&.�nHݎWn��i�j�N�%/pL	f�g���:�l��c�#�y\�и*����3p5>[ҝ��uXeȥ˭��1Z�y�����T!ŞIUnj���A,��}1�2�^(�^��$�����r�.os�L߄����ϲriR������(:�F��f� �9
SsF�27;�ǽC73���^�d}8��u��r���̽uY[|�)�h�����<��}o +/�{b�&q��Ԇ�p��}ۿ�˹Y���Y؅9"�j,�弲����[�L�uaъ��H"�$�u����/[hcg-���(��nj�]��eZLN��1ӄ5qv��q����[���ǯ�";���.��|��!��鱻[��^s���m�H�}�c��5t�t���B>�x���Qaۋ�n�U_ s�b0��5H.R����j���̶`�wa6u�-�K>���_p�-���zdO�Y4�����d	r��Ɔ.�f2\Q�m���/ 6
2i=E�0.���LY�3�j�M�ehs��7�jE!�17עgQ|�saDOzY�;��jz(���J뺃���s�Ht�+�fc�V�Y[�΍��Tū�j&�L�ͤ���{�ÏX��m�=��t�{l��Zb���N
���՜.��7����L��f�Ln��u-�pm]��/��:)�8D)J�*k�Y��qTQul�*�
�ҭ4�4�b�c���i��QyN�F�Ŝ�׃+7���(KQ�:sI�YǁX���{�V:ԵZ�z'^��P�I�xI�Q��r�4���8rh��'�<��:�Uͤ�K�fK��������Kv5wA\�:�Fj�
���,[0+����6��]_8fB�f�e�\�2�8J�O1�ֲ�&@-.���<���Հ͈��p:���7�ħ���[��o.�^��uwF�ǉ�ܳ�7ZA�f��$Q����1z%�醌������cO�� t��G��ú١�sr���:�2�'�ݳ���*�d�23g���2�˳W8a��pX�C�����b�><>f�|n,�v�Ą �Ѭ�ӆ��Y�pz{�wQ�,��@Jo���j�8���5���|+S1���Z3Q ��Ъ�6��s���]�4�����������j��ޛ�	�h�*6���3r7>���l��-�ͥs�=������rk��fP���HE
��7i��{�e]�a�#84�;2ҩ�V�w��j�]ɎQ��>�fõ*6��Lalp�Xe����4�p���ϬNW��Xk��G���e���v�:�Eu�S+`�9Y��\�ֶQ���'O����Z�O�hv&�9�u:�I���r]�vզ2���×����,��2u�aH�_}q�3�2EG���ƈ⺺������w��������v�����m��l{��B��͖6,�V�x���c���gd"+�e��2&5&gt���5���(wӸ�&S}6�z;{��]�}��<&����zMy�y�7[A�9��2��O"{� EvwN�����.�3#�:-L=s�����=O�"���j�A���CY����X�:y�9��R9Ǳ��/��X�.�rԜZu�����$�ү,���Z����ʛwoR�u�\�����h�)�f�w:�ז,�&�5�D�Y#DY�l��9�K;�A�Ї�	�z�����e�B�¯X'4B�(a�Y[g�on�O����쀬;�CD}/�M�y�3�!ӣ�!���D���n	2Z�Ηi�;C,�Aփ8�Ԫ΋�!��DM�ҭr9=}�X�(�asz�m���9%j"��K�r���~�2eJ����:�4�6�.&n]�m��o\V)�J�g�іULN}R*�4#�
X30�ZjV+�+w�� v���D�$�r^#�n�a��R�E�_H���r��-)v.{�v�+����nO��2g=�nڹ|�=;h��9�c�Y-�Ό�v��9��!��f*��@���k�[3̮����,��=[P�/V�H�<e���=�9�Q�S�h� yp(=Pύ_ee����BȠ����f����=X��K[�v��: yƭbos��:�J���FM6��2��5��OQ�:Ynt�"#�/]��k�n��wG�J<I����lzL�c�$����[��r��VڋNE+*mS�8k�Qf�Ph�:���â<Z�ű}6�>v�ZJ�'Q��u�Nx�1�>���q�ꜯ�g��+���4j��w+���b0V˲���,�HS�+���!����
(G��S/ ����ަ5���kY~��J�/��i㬗���۶�ُ��x.�,-mt���s:�t���Z���^)�1)��A�N:Y��m�ט�|��9E��	��r���pVgM��ffҪ���s��U'',pAѻ.t�.9���6�����7~נ���:�汁�^�ݣ����t �jn��bm���������#��}у T(��a1�b�_](#�ֈ��;ø��א���h���d��.�Mķ"��+kw^�b�;�;k����Y���3�mb��Y��ƚnge��d��3.�b!�6���J�5L��e,�|N��"6.|��H�m��ۣX)܂&ێӔ�՞�pW7�*�ŝ����pP���L�;l�yz9����Z�W8�E0���B�Ĕ@7��ʽ���H!�Mm�ϻon�K}G�i;�N�e(���޾�;Fns4��:��OY���+��l�G�]�.�]�]\!�����+������"�p42.�a��Hy٠�lV��&.�M��.��]f�	�		،wqڙb��-���^�n��jy |�V�e�3U.}yP�X,�]ml�"�����v�,�;p��e�\��r�G�]p����n�Z�Ѿ��=N�r�W��1�N;#��4y�{�T���sk>s��}�w	�ȸ�A��D+ݓ��pXΣ�#9�+0[��o&s)�&�\�_b�Kk��,Sn�2�;�K�3����l�59�ۨ6��A^M�/S����Â�{�����������Z�l�
��>�Zpvڛ�R�8��F���ď�t Ŕ{���k�oN�"Jc��Z<Ӌ�:S�7�Q��^c��>5�u���֟s��8%]�:�p,a&&�u�%r{�U�u����;��G	�O�zifSb��t8좐�:��[V��v��i��ݿs�:�V�d���u:�)�W)�]72Xw�k���-��r��z�K5J;�����������u5j�]�<-�mq=°�l+�R>4�,fR����^i�m�QRt�3 )�t-j����7�=H;}�fwp�J�la����e+����xB"�'"W4q�웊;����N�BtT㧻d��gwY��8T"�*���{W9f�:S����k	�����rs1�����L�7n�U6�d=��F7k��f�,<��Dh��t��a�d�������缋��[z���O�|qG���E�{��O{x�4�ӥ���r�X���u�E���MΡ�9�Zל�E�f�q�W���jbdƯ2�}�3�L#wv��0wy��F��@��.��Vr��oK�
Ӳ�ђ�ȍ�u��0���Aٚ���u1�=��5��Q4	���WY�h<1V�y��2���9[w�w ��n�u[˵g�d�7�4��vb����/�-έwb�^�fR���,�.tʸq��s<4�_
�X����5�]� ��"{Z3^;�,n�b��>��;���7k����p7ɋ7��t)WY�'�JN�#�s�y�2�X�E���oA�A%���m�ohe�o�ka�0�����-ۡ��� +_ٲCS'|nG�V�Bi�:#��B��:\!�� �1�D�':�*ĳE;������6]�+�+�������e�����v�<�}�`Gf_9μ��]M���`��h=�[Rn�+#�+�������\�gTLR5�8�Ƕ���f���(�7��Jc��HΗ%k:�Ron 3[�~%�e��MotX�ժ�)�h`�3
@�P��	��W�5H�CO��a�˴�V@�t�ԨE�F�e�o=	�g\	L
�qC���A�k'v�<��*�b5c1��՚����I�dJN��k	�,}��/V�^N��'Um٫S�(���1S�����i�S�qcnƵZ�&^ٸ[��p�o3�i��K�3�C4�1n��w|�q�*}�έ�˅�Q`w�
�D ��&m�\�ȴ�l1��_S�tx����JN�1�9�jD'����ݼ�ZH��J�@����I�w+vh�b�^6��;B��ͨ�L>5�M�es�E��g@>�;r��۷Sk���L��n�=@��C\�C,�OQGmD 4�	�ЇNhҮBv����ug��Y�9x�E@�+T�<�2f��s޷T
�qh��On�9f�ZO���1JC��L�<sL	�$�&�[�P��Ъ-9}ך�R�i[p�#c*�n�]R��2�1��fM��j�
5�5�������}�.)3hش,VT�
�s�ȠY<��e,��ԤN��7�b�F[d��:]�hf�2<G�3a��1c�ĳ,��mъ���@6D0�po/��F��r��g<W�����
1Q÷&rұ����wy�~��{^��!@τڷ]��&��s���lDq1��hܐ�z�d9\�I�T�7�Gz��sl	Γ;�� =������F��α�
]�o#�2!�����)���[d��nq�\a_fM�Z<$l[��=0NyK�Gy�OTE���ڰ��Y(�wP���`N�.�:�|嫓�]���3;^!.�e� byR�"4ԓ
!�()���G�,��%�T
9[���)jHU�j�Nm����|Q��Q�ͥl*��A�ý�%i����q�L�'V�QAlbgon�kS��e��0{��I�p5���g�z2]	Rh� ��J8�wg+�E'�B`"+C;�+p�Ew�N$\���yn��\ 0o��Z��|vK��`w!I����'�q��L�q	��]6�;`8w�P�3fŠ�/���'�ذޓ��s2�6�h�^�1�f�#�s�T&�w��زBl��GWb��6�V���t3hP�a��ɢ�ĝ�v����1�=�X�*�)&%�socv;�'us��V��so�B-�:�3������Ε��Α�˭��&ƱqN���;j^��(\�@f�h�q�0�j�0>�u������n�r�8S��s�h�%z"��V]�2��q�n�㧖��6k��h��[�>�X����!��LwQ�js�7�|���n��Ol���I���g+3D�)ca����U����ho$Ҭ��`Os*�,��v��i�e����9^]v�ҵ��pf�b�__<ߝؗ:�5q��5���u�1}�(�x�M�s��ǻ��j���z����=]tm���n�vT%�~��ʴ����f�� :�����L0F�tX�ue蜨�l�[����gS����T��h�+xd;;�D�[\u�#�f;}��f�[�˯��#�ҹ1� @�۔��fIݗQ����tM]Yw����v��q���tu8�U;�K�h�[z �}1`�C1$tY7OJ�3&[Mwv��ֺ.Jv���r��M��x����Y5tc��nW_s��8D�ܡa>�A��]bq%A��o�2X����M�[���6)��T�жk��6�noN��JJ��ql�M�9�\i΄�Y���'N�nt}����\�jBQ�^N�ݕc�.M�����tF��L,��x�#[u�VU�;J0��c6��=&�W&r��]+w�K&�v�̹�|�p�Kw���ܥ�*�je�r�y�YL�2�j��R۳�Ҋg+�J�c�puwf|�Sb]��ȼ���`�� ��㩔�7�&_=7l�f.�\�ν���xc�W���GZ{���x3��D�U�ga\4p�:2��yO�WN쾼�����N���<��/��Is�wq�uӠ��Ӎ�wvs�B�Xa|ւ��K���V�+�u�9vS�g���3�wvj.wovwww.���\���}}���N��c�@'R�'T��9�-H�potۊKQڥj⮧�+�֞[ͩ�����>�� |(�!�� ���q�̉��/Ϝ@��:�z��<��|�G�DiS�C��!� ~�>�)켞�>�y��{�z�� ���)�N�>���r�\�|�9{ז͑<�뀚@�˨S� o�>����?ު�*?���?�������O�?�z������_�����g��������?������Tx����:��Vrv,B����o%%��+ճ(>�ռ*�\Ti�}T�k��p��e�*ƠC�gS�u�o,�+woK��on9�!'>nC�@+;���^Ik�5U�$�����v�v��ͺ��wK����7���t�������Y�b`Ӝ2��.��3/���tKE�4��ɋ�']h�̞֐͔�tj�3����J��Z�֭�A��ܵT�l7ثg6�u��c�L5�fN;���y7��Y���BC�4���oC�3sVʻD8:���u}T�F˻~��fHnl�@o�Ō�x�.컕c&Y֎14\ɴ���y��  ���u٧�4\.�V,[�����p�9�{uqh�����M.�nP̢��i��$F�ȒX�e�\�t謴��{o��z����W4��W�z�F���,W��<S%�[:��z_^Jɖ�����X˰�[��f����EU�Y��vPx�wDb۪
>
���{���(F�A"6��Ζz�����᤹Э��	�d�U?V,���E��ە�^=:Kbtڙxﰞ��*M̶r;��T[vt{���P������̉m�e�q�E�d]��B.�=g�8.C-ȭ}�i&Is7H�;-�o��Ϸ�}�����=>��?____G���������������s��������������}}}}}}}}}}}_______~��5�1���@)�w�]�2h�1��V��^9u}$W��ti��̭�vg�zA���Ɇ��p�� W�Yz$���w�ޒ�Q��Iy|8f��
G�0�89RC��M�I�ם�y��}5�n�Hݨrݤz��L9�HCJ��q��_L}y�¤�P^�f؝BLQtj�g�X��ޣp��%��Ft��YǺ�s��J��5��ÁN�X:�T{k0�:^Ispαu�,����b3tO���7k��<�|Ț��[��EM�v����ݍ�gd�}sJ��t\�����n��Rt17s��N�֎塅��T���_K�S� �<o`yS�u⮬&*��j�%�U�6�����ٝw��^E��(�'wܫ�3Zx�e�g�b��"n�܄i�tVE��~�ΏslUA�W�mcu:F�'�l�}����f���n�������1��0��1�aL�/�LtTےt��*捰ή�N,���EO���F�rXE
<���;t�Bo�]���M��>����l}!���e�`85���R�%R�6�i����ʔ��Sf04�.�˙�vA��n�b���Z�5�(���l4�G+q}6mќ��7c5��aI�T������'�[}Ò�,9���ۥ|훕�\�o��E���*����c�[N�����__��}}||}}~�����������������9����_________Y�������}|}}}s����������輪�}�o=��~�)n�)ό )W��`;5b�\�ꊝ��yr»
� �!�.T��t���v�b�	�!����0.�U�a]�m7��?5��|���9EN�����H��<):��'�'>��b�W�5��b9�����Ng��Az�W{rp�ǫ����^M��-�T2��M���ᝁ<��	-D[Oj�h�̎�f��Ž�:)�D�U��^�K�4p�yVSݓ�\yRxhuư��rdP'��U|�k:�} �]q�c0lm:V��Oj\e��ȟ3��]/�0H=���&�Um�QT���ʸ�^v��j+�^l]KeHf���>ő���Sޙùn@E-{���Y_0����knP8�2uk�ł�M�f�x��u���T��D���WD�P<�T����yU��6�6�̾�v,�X���/O�"I(@�6��{�.�w����7��
��{r*�H�a��3fc]����A=T�5�
8)V	��ҖK;�u��|0�.Z�:���R�}���R����r�Ϻ=�Q�Y�W1�Iҹ4��y��L��|9s5f���?��8�+J�8�Dы,���<�(�� ����8�^�Gc'o-2+:�>3v���ٰ��r>,[��Vg(oM����������������}}}s�����������_^9ϯ���}}}}}}}~���������������������������wy�}r�ӽdෝݽH�V��0�E�PHc�7M��֞�����c��5A�7�7�pۭ��JC��x>�&<o+��z�_h�^�O#����֬��*���]�m�;跍�yPc��SNH�"vm�m�I�GY� ��V����4����	!�9t�!*n�!��Q����Lb+�׋;O� �2�|C��nݬ���]�Y�Q��݋�w�2�pQ9�W�~ ��T�|�����ӆ��M[3�U?fT���ڧ����vm�uǥ�#0K�+�VW��V�{yū��<wf��}q^�G%:�����D�����j�2�2�����C�Ӓ�3���|���J�kM�aל�<�'�'�K/��ڝ\:����T�v��yKIuL�\4w�b�@��By��
�=�Ւ�Q�ZP.�Ʒ��y�VwR������N�]�|>-�+� � 7��6q���ۖ��;��� D��3���hu�2u�b2�Z}�7��.��c���m�t�L�v�b98�� U����#/&�P.�b�b�p�"}Í)����gu8.��S�����kN���¦�/'�r��@S���q��S�c�G�4��2[��������������������������������׏�������������}}}}}z}}}}}~>������___|������R�4�fֽ��=+`���Q�#�Fb���#����%��X%�#*dsn�3N.%Т�;��j
itl ��6TA�{Ƥ�l>��1tG��GU�RE覍
V��z���9�+Z��l�.ۢ���d��c���5ܦ�w޹K,:,sZ��.WG�Q��vP�;p�����m�ڏ:Lƍ�<r�|x\�-���\5�<.��:A,ok��cNZ��;6^\9����6.�I30wr��w��������v�9��9)�"�B:2�y\ݲ��O��_|��_ �2�S��t�[�u�n
�۬��RY���V��V<cl����<ʕ�hk���~��K���p�	�u�bnG������կ����xZ���N�՗SA\�5K'/��Ks�����Pe���Ԧܲ�#��`��2��s�a^��\���R����}q\^l靻IpLN��`a���s�A�l���GqO�]̕ڕ�Wt�B�%��7n#�VP��P�Q�*�.�*)L�Q5�1Yo���:d}�+$��,.;���J�M�d�;d�tuܚ�ћ;���2���(���xr�;�k9�K��r�B�!�l��؃�vJg�st�x�}~�__^�__^>������___^�___^>�==<}}}}}}~>����>������___^�______^�__>_~g64\��.�]��j�Q�b�*�(Nh�y{�{ ��C��<� ��0�}U�.��g���^��H�/�z2�j�9�k��d�we)Om@!�6����6��+��^ʆ�Y")sb�����3z�X�ᨸ)6>�n���D8��9Un���q��P<�7;��1���<�����G�U�����r>Y|���.��l3�Ւ�6Vl���a����j3��ۉ-*\��f
㽵��<A�pҖ+%t��*&њ�Z���ۋ/�xڶ�pk/3��6)݉�7�(���w����y��]�&8����Z�Ћ��_��������F�N��a�f�3Vo]]�""�v��5(!�p�e�k�����rc���p�Y�K?W�bD�B���ɕu�kXd��9�����V��U�!��_]���d]3;��tl��AiX��ZT��l�+�Q�	��-��6�Ѯ�=�8�hf�lp������e��W �VTi-��^�������|ݣ��O%�Z�teÅ�}��C��k�C�3a2;�[v�ʬ�.C�I�XWPe4�}�� �.��˪��^8���d��A<��������%��RS!���ū�D �n��~W8�O3���}�?����}�?���>�����������}}}}x����ϯ������o���______^�__^>����}�w��}>P��d�ׯJ�4q��T��c ^��2��q;zw�G/!�lak(ʏ~�99�ɹ8�x��gq�S���ϕ�ބh=����r�]6��i�e�6���f���Ҧ�i�E (b��]��̽o��'loZ#xH�v�ev�����{y:����N"@����9隠�v���ɯ���į#T��d�lV[���[��J�m�#�s�զŮLn-Vam�m�{p}T�{�����+ř���R�-�hm��_����*e���^\m;׻�ND>�&�-�hդ_PO�,jX��,U�|�1��B�X�|*&r��5��Pxr��^}_P�W�h��3y.�(o�M�����j��2�$�م��{^5�,#t����8v-<3	�R�0�\��*�Q}ʤ��������b�S;1>��o��g]`��������*;�2�#����P��s����q\��syn�l�lL��^���	�ʯ�X)�����M��rv�&��� ��ٚ�˖$�Z�M���f�mf�n�U}\Ѡjlg���H�M�ķ�B9�{Wp�C:�{iC�8�b�ܰHlo*}��:Jo�E�ܴ���6zn�b����&�.LL0;�u�A��\>������D����/�U�Xe�b��wn!,���sOed\5C{�Ϛ��E�5`�38��R��s�䭖hj�	M==ɫ�,@a�=�o������������������}}s����Ǐ^������������������������}}}}}}}}}{�;�כл�V��jط�Eq�w��_}�ue���]��r��nq��P�]�Ǡ��ҍ�.��+AN�:�h��7���C&�_
d���Cz�R�L@�-r��&��Me�Rc�S5�n���K�:�r�����;�g"��	�g%Bi�M�tGk}u��뢌�d""��M�C��(�Zx���PzYu�k����Qպ���S�cRDj
{�ӷ�x#�.=�$⁽�f�|���'��ۇ+�_o#z�S+��P�0-I��j�n�ĄX~�ϫs2f�}Wi��C�ɶ�:�Q��C8U���Pm��U�k�F�,��S�֛��7�l���e}KiU�lv,`�60h�M�Ej�:H�b�?�^��5��+�j��-5t]��I�`!���&p�����T���6	�$�M�KP�̚���2rF��H��+��7�Ȉ|���e5��h^�̕e�q���*v>-�)��,1&kT�����6����� r���4��`މ�ŧf����N	����V)q���P�
8�R��{���u.��WΝ��yM����H�������^�}�}_������uu��њs4RD���udW����4&�Ȣuc��K�pΠ������/N����.H{��v2��|��%ڰ��	�^2�^D��������2�J��:�uf_b��?RX{:�ϝ�^��o������������������___^<x��}}}}}}}}}|}g����������������������}�u�I���,���3x77���KN���E���T�r�eʃQz+��[3sn�7\�l�Pq�{XJ`)�H���ZJW���2��f�O)��2�P����9�@���.��5�*���^]<���6��=�=��tK�����-�J���m4�����s�m,ʼۆU��֋���novuh˒�} hkN����$/B׵�n��Ur�Mf�aܼy��8��D�\�j�]aIJ��̏�J��:�_�q��U�V�u�+�fsO�3�d�����2`U��u�,�8�.֦F�V#���\�?U�l�:�-�!��*x��04ʃ���b Xu��9�����t��ݎ�*��u�2��C;���:�D�4�=Ү2:ݝ1�Y'�WvWt٪n�T�X,�\U8�H\��9q�
��;��Y�0��j�}�nq5���U�;��Xt��D�x�'j�iңٳC�{���8v��|a|�����\�!�.)�p����Z���!n�DQX�{zv�ʂU�>�L띁�u�ޒMm<}���ʶ�W�b�NbJ��:�UY&:���*��^H��cq���&�����tF�+�H���T!<�.d^WK�;v��:�R�fn���Uq��LSwj���n9�x�v,��ʗ�T
�H�:n�8ݽ�&#��W�R���L]����vu;9K�F$:S���r�5:��X���agP���P��J��gS�FZ�D�Uo�$	��&������WM!�b���w�����R&�e��]*P&��B@9k{�GLv}�{8n�ـ�[*'m5vp�)�ՠI�C�\N���ҍΡF��`�t��4��E3l�[�I��h�Q
�AԮ���+#�Bz^`5�MeCD�qF[�(_s���������W�w�u3���R�s;�Vj��i�e��µr��wq��h�V���C֬Yjڷx��t��L�B�w�J-�Tͩ;f,�*���{�p��P#���$���,��ø-��7%��uG8��坻��
Dj
�R��В�7:J����ۢ"2���J5ЃF��ַp�yvQkgv�=N�M���7Y�0��W�Y�|��Б�O��h8�Q����R�'t�@Ñ v�әJ	_}W�Ç�-x�`[��\��?Up�����b�p=��$.�Z�@a/SO�%up��8�f�c!�r�tX(���t�L���c8].ͷ�p�3H��*܄�M-�F��Q��X�/�|u��
��´9�rC��l�8�=�ئ�Ϋ���+p �ެE�v*.鞓O!���ב����䖹�1
�fc
�;� l�09��]a	�¶-r�7�L�a���J`�f?0/(��ǫg߸�����_�� U��s������?���/������?�/�
��E Q$�PDۅ$-�l��r�,�p��0�1�TR�	����F����a�H�E~M��F0B%�	B 1	ND`2FR0D$G���%������E��("b�4�m�􌴣��[�$8 �|�.$A�
H��H��?2BiE>N#���A
MO�d�[!�"�I�E(Ҥ��0��m�_��^&*�D�������B��G�H'`�!x̢�QF荲^�{��T����j��<ݰ2��	.r�V�,��xT���� Ի��ĭ���o]�b�{�E0�a�C���ﯝ��b�l����b� ��U�<�9Gc��x(V�]�������X}Э��Z�Cq��vav���X�^j�4�շ��x���sXaHw,�D-�`>�g7Ue�W9�S9]rHYU�5G
�1���Û�՚_RA��X��#W��"��6�c�K6��o���G�j�,���E����X���D�
c2n�\\��c$g[h�}�SZt�|4i�W���%��+z����4
ޅ�4M��7��ݘ�}0k��|���y��u�sR�2�欺k!
�u+UL���3@�vQt��h$��ⱞ<y�6/�c�f��{*
�ª��}ԟ-���w�a�CU��Ʃ�'p��K��y�gC�Ʒi��E.��R�$�ƭ.�x�����Ϋ0=ݽ\�F���� ��e�a���M.�ĭ����a�u-�G�(����璧q�cfi|�jE�L8N��⺒�݃ؖ���H��]q���4�e
h��OR��*����9��7�{A 1jB#��F4̀%)��0�-KNB�q�	)� �¡F"�e���K��%��nH�h��EA�*2� (5�m�``�D�����n)!a�B7('�ԅ�q�T�"X�	�!�B�
��C,6�i�����)O�!T�m��}
h#D3he�"��X!H�D(��GJ6bl@�4�)I�D��L�"-6I�Q#*�f���m�"7�@�0B��8	L��q��L$�2"ؑ0�.F�M(!I
P�q%LEDĦ���̦�7�RB�-�$�'��P��q�L��%�҅�f!a4�)?�28�M�p�Z�ڒ5R$'�2S�1&�M�!��*��tۀ���R'0$�P\�4	,�
#e��Bc*�ޣ�f5�9ͬ\ى���"y�I�9&j+�n�=��:蹊��mZt]bz~?^ߏmC��D$��_Z �K��1 i��Ds�ձ�#��7lr���������m�TZ�\�;�s`�8�Z:9����3Tsuu�-�^���y/�����{~=�Ov5��k�����@	2JPƅ�_$�B�a�c�=�UU:���sͯ���������^F"�X���\��X�`�m�	.�L!dx�$E|L � ȅDBg���A$H�RsȬ����~=�9ͣg�g9\z���9}���b�5�����z�s��M$i0�H6A)��`���'�?g�9tE;�N9����Ύ�j��������m��k���Y���G79�n\8H����হ���R��uns|���|�����<8V�v��.�����u�9j1�1����-���������;�g�-�7�upS�s%k���ϝ|�tUd �F:�p��s$/�ɨd_܉/�P��L����8�Z���.�*�s��~�^���qo�5�������bѶ9͝���W�X�o.T��b7u�r�ת�y��ww~c	�� %��pϚ����0���H�A��m�B8���$D�F|�&�G�P2�$�R�Zf�4���R�˄� (P�%�|�w�E��,�ME>,��& �$��"
i��1e�F��@��Q�i�x}ܮ�}۝����޻Ԛ9Cq*vO<��'^�K�eo{T`,s�*��Y�����HbF��'����1@�!�H�p�̶�PE $dRB"KQ�QL �d�>AF�@�,@R��ᛛuțh;�=p��|�c�n����HeQ�d��I��if�E�Wg@/��"t�r�.KV��0Q3˝_��@pL�ﲧ����ކ�%{�0g!'�};x�F��>�Z��p4�}Cߺr~c�|o��~�yU6�x�҆
�~��b���3ˏX�}b���� ���������'8��q�{���oǛ�c�㞯zE��S��i�[Cޚ��Q��	�v汷q��wܥ'i���H��{��*��>�'ݩ�dgz؋��^����%pN3��ߤpoooP瓵�wr}���3���YC�xx󹄼��
�[�z��%��WԱ��zeE݃~����r1��U��))9=c������X7}�rcH���~j�^�;��J�M�Ƕ��'��^��%�I�e�-�-��Tq'�y�� q��w�o��+t@�q��{�������y~����Y�R�"{��de�b)r�J�-���4:������ٕ����7�$��p��3������և�z�\��(��mߩ�ӥ�#���.�a�Ӱ�
�\\��j��0��&��9��G;@��#]��ɗܗM[v��U���Q�}��X��{�E�o���9��vI�Wd�'����G���l������z/��,���t�3���Z�K����h�����ut=c��_��?����%L�����ݞnuu��5�߲�w��{t�4�W���#���L���|����}uv5✓]�)�=X_mf�#K{(����S��j~۳�7�7��Փ8I뛸��`F
�����V��ӗ�6�Q|�	��9�;�t�pm&�������H.����נU������G�듑Z}]�i#��8��q�o�y1=RM~���]͓��vߕ>���42-��?%7���zJ�i���x�k���������,^��م}0y�����Ǽ1W=��l�_	�2�G�e�ݠ�NP&���y��7�c�c�]1�[�E��$:�����v=LT�z�#4���p+0r��7�Du��"0�~����o��ZMDn�pw��ǭ�Є�x{6��w[
��vxB��'+�w^ݫB��w$7�|��V�q���l���LwNwʎ�Wӳ�\�������O|��;�~��ӥ����j��6��9��틇|���Kd���e�ߣ��9�ֿe金�x�c�+�3��'c����%���*p��
��X��5����n��}pxV��ov3n���ƽ�X�&=���L�?�^�Ջj+ a�>;����{�&��Y�/1=m�^�+=���e!�;��.�׊�������X_x{��r�	�d�|Q���ݘ}C�k�j��;�o��;�Ƈ�P#�I�˵R]��'�����{)?m%3��*	�*�t'�{j�ս�l��\��{cm0��4q��ۆ����T\��x�v��>���L42�9ۯ{;��z<�I%|����0�*��ڕ]sޤQ��zs�9�/{םy�z�{�}>ўi�5���r��)����*Hj��V**cS6����C^@Z��K�js���*]�,r��k��A������jǙ����.��;*iY��6�`V-P+E�lWc�>S&�us1VB)�A��=���O�������/	�S�"�h{otez|�[l]�x�Qܺ�uN�T�����r��R?���Y�\�����P��#����P-�`�i��f�見���d��&�4�`�YL{��+E��Mw�;ñ�j����,U��ߚ�G$ڃ�d��^�B���i}S��8/��(.��������z�G�Q�.�$��g�~����z|����x�}���7'3���*��?6:���"��׍����N�h�sD�q��������\f�WW2"V�����V{(�^����pJ��s�s��������x�zd����;��j��k=;VL[�ĽK1p�S���zt��;7���w���&U/V��wb��P�p���=SgI�ݧ�"u���U�ە���')��N��VH�fǞ}���'y�����&o7��<�4�w��=|����,����[����[�V����)�^^��i�����!�p��M`��r�fk���5�m�g2�L���+��[�m��aY̹Ǭ�|z�`!2Sz���w���w�H����E�s\�Ⱦ*���ﰿQj[���6+mgP"l��#�"}�e���r.��_<��,8,P����O��+P�rCM	@����nG%��1���D}�oR[*wG�cq�u�6;�r���=��rO���Q������8��ܘ{}>c���O����Q\��X���jzצ�h퍏�؀3Kz�}M�(9��.潡�磫�&���曈T	h��p>aێ2v�x��i�~�,q�]��v>W���y��y�����>��1ui��\=�s�O��>�ȗ�3�=�����q�PL���<� FL3��1T��'ǽ>���E�qך��?-�������3�������	����]�K~����/$9E9�W9�<�({�N����O��;�1�ch���H=��^�A���I�$5� ���<�>�W�!T�^__����N��⛠��=����B�V��o�^�Oݚ�HW��F��`d��}��Y���WY�!�5�]bo!���:=�ҕ��Ϸ�D0��L�벮��ͪ�����*:���?yJ��B�@W�3S[�z�d4�t^�99��wR������*r�ک�ݰ�ӓ�ˡ����fp�g2�\�;�i�}�ћ�p�ܛ}XwϺ�{���N��9^����fנ�vdq��o�Ur.�k;�}���~",fM���o�Gq�E��=~/r}�����z��5���>��,����o|��za�ͿLd
��nH't�C��������|s݉7:3\�^����o@��7�+�&g����W��ow�Q�f��M��n�NcQ���Ldw�a��`����1��.q���-����\}|=�}�w�j�^跔k;s�j����s�e�c����׵�*����'Ubm��ɛ���`ս>���Y��&���|�kP0-�{$�uӐ�7Q=�M��m�����ԫ�oZ����E��4����6��zs���~�����fI����X5�S�������o��M�+�^��3����W!��쇼V��{ٕ���~��i���=����<g�a�9�
����C�ݻ��|����T�dǽ�x�_G�
�ٙh(��VE��]�׽��s �u�7@���>G�Bkv>&�_س	r�4�8QV'9KH]L�#�!�i�F�qc���_f���ϵI�{�S�k����_�ލm�}~s��U�������j��52E;w��wT^q̪q�(���K�"�8�B�tϽ��;���K]ٰu����n=C�d�n��`�cR�iGQ�ߟ�y�����\���1��\���x�N�⾆�8�����oM��6�����F���U� ��.>��R�%��\�NU|}��Q��ʌ-��{��>/�����]�"Ω�{>�/*�s����y����vw��WH�&�{T������ʔ��|�pI���w%�a{�]e�4w��_A���#u�,�I'�c~B��z�4�]��Q�E�3��Y�����L�2�_w.ǜ|��>�ǹ1����|(������|_�<��֧j���6K��79ћ���&���w@n��AV���sF�旆�fD6���奨#��nL��a�{�ȷX�q�y�ݾ<6�xIY��hzB����gU���*u��O�C}N�$W����[�+��J�Y��%>�f��՜��u%�YϮF�V�[2������)ô�J�W��)�)�ve��쨟o��\��J��wM��<ﶭ�{uW�+�Cx������C�÷������ulc�������WǸPO�divW�x�����W~���o�ptj�,5�k�g�GDئ�[������o���uH$���J���Wq�mJ~�����A�,	S�1�4r�'�ӫ<�o��(�Hz?S��Z����`͵�r�/zή.7�7�B��D��y����>s�xm)��������3be�ϭ+����mvg�U�^s�2�WٻG�*�?o�yg�{�>^����,�y�_�����`���zs���<b����/��g*û-�NX%�{��[@y`oE����^=�9$��F9�7�0�Ͻ�/��|�=�������|�Ι��{X����YЩ����`B�ޛ�Rj��&��e�������S|���r��?f�mJ�y�c�*��N�Ƴ^��1ǈAis{���0�}bv]�H��Dw�S�qqX��yC.��f��X�G]��)�o5�
�4��î�x��-�杍���g33��!��	.���7|l����/"�iC�B�	O�!�p���ԉ��;�Mu�n|��{�~-d�U�{c��}9��y�r���g�~;9[&���N��q�}�6<Ք�o_s��|=���%~6/s�ܖx7y�$/�Ov.����G����YwV��[��:�3D�w�r��Lf|Ǎ�A��no��{��Rw�W�/(5�g;�H�dJ�p�=5��>�e^ό�_WK�[�U
fm�mg�T���dC�޴Ou�o�ٽ[����/��M�!���y}��j����oȩu���_��To�W='��ʫ��^�8w}��]>=��t�?&�}�ޜ��&s�Ӳ���p����V��xXc�A���k9�3|:r8k�o�y˻�{=�QBPI~�H��������ެ��U��܃�l/�o��ݳ�&^դn{�;úV%�����'}�j�ߺ�s�e{�L��e�Np�ḧL�P��l4ZYx��b�ݾ��*��v����զ#S,�N��?�h4b�!���%w:��:����9۷��L�ҡ�}��鬊+"��Su�NC���p��s�U�dgW,笍Jt�
N�����_M�o5Gɭ���|��M?W==���YV��V3w�/E{�Hj{q��ƥY�ݰe5��=�
�g^à�}ã��nڛ<;ns;:{���	5��0s�VT������C3�'���x�{���;�R_�9�}��]7�_{�ms������_xe�"�&c�-.�]����{�ƞ���(s������<E�ԡ��9��U������yP�*�l#/כֿ��l�%ݠ�z{|$�����>y$)�k��7�����$
�s�"��6.9�U����~�=�zA�׹x�̣jqx�9̔������E��:�ψх}��7����^��w��7������N��^��[|��,��κ�J���s&�!���a��t|�'�O���$�z�1������ᤎq��G�����߀=պ���E�kf���9XQ���{.X�o�����8s8ۖ��XYa�k��r����%�C���jm�[�q�1@}�� ˻�zf�~C� ��҉�X�5]2.�neev&xL�Au�d�����w�#K8�z
y��wy|�u%,��JM�A\+��� ��ʑ��7�i��MqO_"x��9I��@��)�i��f��E�U�<�t�Q��w�I��L-�Q�y�_'\�J�8L�a^C�8Nr�̊E���O��狹���V�am팠��xLx�>�i�p+�:;5hû��c�K�W�`�kd<��o幻��}S;c��������Ρ&^^jW��<�do��6�>��	F�m�v��~b�kO�}G�~��KR����&ChEh|�-�g
���jT����L��0�MzT9�ٽ²_}&ͤ��Yݟq�أ٨`>0&xaW��m3ù#��w*��ϥ��h,Տ��')��r�,�y��1��{W��G��ژ9���	�v;�K/:e�}�v��f�@Ӯ'�ӣϷ�F�)Ue�'����N��T��7A.)��f�)ki;J����P��+^*��@-X�����γ�^'fnZ�J�B�g8z=��jE���ifv��Ł!F�a��hQK�x��ء��qU ��k��㕔ɝ�����$7_$�̣Fnǣ4'�����UNqu:h����
hmN��l�n�.�Ih�Y"��5aÆ�1�Q�� 
��#i����	����c����Ϧ�'ݑ�ݽ}�ݩ�g�1,�pЧe��(�-[�	�/]�8b'`ܺgul��Z#39:�Z�ʎ��c�N�1n`�3��
i����)u2����VdI��Sv��l�'�/Y�\�f��{M��Z#�H=��U�EV�)�u�uՀҸ�[;�����@h�ڬt~ݷz��:zDKqN�x��4��2)����x�/tfT+<��J��Rz���q�b��Tӹ̜��3&��dX*�:v�ȦrH����@�z���9%��t�W,�ީb���1�Od�ܮ����Uâl|%��
W�X�Ί���l�Ŷw"�:��\����څ�Ĥ�Kl��r��o5We��-\�"��s���-ˆ�}t �:Uͧ/�UZ�����	�a�C�T�A����]�M�>'�d\u�}˧r�s�*0=6��l��X���N�=�Շ)a�X�倬{�Tד*��ڶs�e_J�V�3*[�_mS��,$�r�MdrŠ���N�b��K�c/u�$�ˡ���?��thk}WfN����2�`E���:�T��6�]�9������^�a� T�Q��5�p�X���\�n[�)v0P)��9+���h���:�R���W7�����R���g����7�+򘭪5j"-�{�q �D� ��<1ࡧ�p�#�� �(dAM�)�%�gnO�׷���P��ɶ�����K-��!"D � B���U�_6"/���c��sp�Z7{�#�nm��փ��������+[�b��nX��]\�)��|�u'*�wd���]\(�\�|ξGW	�w�,u�]~���oon��_ B��:nT@$&�M�R@� l��@�jI����9���nI�p��\7��Ƿ���ERk��Dr��#�rۏ�	�%Ί��$0��_/�F�Ÿ\�)�;s�9���{{~=�7 ��|�<�r���o�)�h�Pؔ >P��1�(h_PC�B ��1 �,0��8B%����������G{�w#���Ϋ}�W:y�<�j�L|�|�]F�?3�Dl�Xƭ:�l�m���1� ����>����[���}t�"�깊cu��[[�g��Z��ru�>m�k��h�ˍW�s��5����OoooomX�>P("���`τ�k�MMգ�1�����㖠c�dC}��M�	|R>��:�JJ�g;�91�r�9�%�1%�i�}
 D H�Q.���Z��}�1BO^g��,AT;�K��+���)[�yӻ-�=�B�Q�t~��]V�ѨwA���in������<x|��#�7��ܳ���?H�O%~[�t)����DX�9�L��ov�T׌�wkzwh�C)Qr�%�%�͇2C��t��x�-A�6߸�$��p�j]>�mP.���۶��]\�����&r}�5���ߓ���h���ۻ]�ӴP�(6׸�7�3i��&�Q�{Ihƥ��|���v���
i��NxMG��\�I�z��xM��;_T���U+n�+�? ZX$;��*�:���*}�D��o�%~X�����������P];���0e�1
X�����Z[/�5M���,��d��d�m�Z�ˤw���1���1� eDu8����gb��r�﷛��*P	�i]�^@k�c�dRuϚ���o�m�%9�eFC����?��+�'Z��y�:ίs�4�Gl�md��Y�oNyƿI���E� ���֦�kh㓐�6�[�j����wrC�޶�R�E��<�}��4����5�,����}��\��Η����J�	y-��8�t�R΍�۬�v��^���#Lx_SF02<.z���"�4��m�S,oE��qz���K��O�X4��4�p�����T����6��xt�9��Uݣ��=ͬ*���JD%]�i�k*��$l�7����{F��{/ऺ}�� ��K���e�4�¹���\�8�:���A�[L�܋�i��AK���NEX����w/s �ot�Wo�H������,�hLw�^�`X
y���w=K�]��?1|���|�ߪ̂�f_�ɾj�.x�s� y�zy�cǞ��7X�$c`(.xD~{�
�j��?gy2��g%�r0�y9Æf`;���0���.��g�5�M�#5��x;c����M����奅p�x�;r��L>0
\f��c�w�[ٝ=E8�Ү���*��4��Aܵ`�kHM��t�v\��ڹ��f(y�v��Қ���q�?�,��tq���m��9�6�͗�ͳ=�s*��?eX/`/ߐ,��O��Z�#�S��}��1��>��-�Y����|4�:v���J�R���D�?��4�P�@gܢ[��bj�>ޙQ�ۓ粚�n)�n��RT�l���7���Hsٸ�i*��ъo=�~�6{T�=s�!�Ⱥ��O^��mV��d]e�7B�骁��h�'C [�֝��"X�� c��3n����[�!�`�}[��[m�⅔y�wq Z*`f^��y"�M[� �}f)8�Ȝ�8�[1@�b�Ң�ZaRk)]E�M�oN��zƻ�<��;ms;H�C~vD��a��*��x��s~מ�����ѓd�X��%Qm!f�3�kF��X��jU�[�{�� ���r�A��G8͆�Mᣭ���V�����]3q�Kub����9�$�{���	�)"C��q����3,+d�!���$�
d�BL! 4�W���ߠ=G�'�U{�����<t�/���	�'���P��r��𹹳R��Uy?k��m��;�� ��o\�P�I�[e���b�NGO3;���J|�I}�rzv������S�����K2�ͫ���jZ~��1����v1�k�3o�@^����I*�s}����y�S~�$��4���b�#9���z�,/�ܨEఐ_��ڧ�Z���,D��!�d��,��L�� �|�U+��;7/B��:n���E���h�z��Qw����j����p��G6��������FK%�/N"g�m��QD�%_���yט��=�,�K�dm.`%LG:j0��q��zhUw*2�o�g�Нc�8�	Io	�!s�H��\��8�K�x��E>�w�47�Ρ�3ܞ���� �S��,=��W�w�����=|��*�z��+�����Y���~�=�?i�ߠCR`��\��[�&4%N��t���5	�;ٍwyH�p�E�/(��F�
��({ɀ��n�v��6���oH��/���z��#�`nX9d�T��
�y��d�����ۃWtBԯ�Dqd�0=����A������ENz3;� ©ز�4=jF���R*���Ҷ�����^���4p]�J�O*���o8�ۮ�7��������DR^܊پ��f3]N����Fs��hA�'!�o{���ӯ�'$������{����X[2Q�b���Q,�怈�l3�`&�Nۆ��q!\`�!�{t�]v�K�L��6���0\D�E0k&m�?C��o;C`֗8elZ��-��YF�m9�mC!�L
j ��x��>̐�� ,a�ܡ��"r��j�^��=r��m�f���W��Q&;f~Ln��@<~�B!Ə�R��?~�kg���.�ςeI]xV?nᔏ�e�6�+@�9M��K�J��,?p ;�]��ѐ-�C������ǋH�SmC۪X�7��)BWz�N�e�jw>��K�[����L�)5�K*k1O����o��P`#ֶA����5�h��;Z��U��������!�2[8�,��g��b���ײg�}�w��r2�@2硱ڟ!��Y��{f:׋Xd:�C��:;�z��t��T�� J����m~3�laM�{j�k<��)�ڗ!h���Ƅ�X8#YV@-i�X=��JW���{s R~e�ͼ
�����]��b2�0�=n�--��R��ޑ�I���ȖS�RoOa1[�oĪ8�Z�-���H�vʢ}���_mcu�vD�_t�C��ʳ� �ziI�Tn�pL)H�ͧ��Ժ��]�1�P×F����4 u��]�̘�q�Z��V��,�b��������ū�:�NY����kl�׈��[�[��}�zq^����;{�m�׳'�i쳭�	�ע~�c�V���D����ԇs?O(��g�㍅
w�6�>u��v���ٖ��B �p�������ky��`8O�o�N@~,���t�U�+����=�v�t�7V��ב�M9j|�$��	�o�-ۋ�k`z2G3�`��&p!��'D��P��NN�>5\�}L�V��)��Nd�q}�c�Noc���I��3����������Ci�e�)P��s�f�x��x!!E������3���"��"��1�a��I�����n?�����˔���+Nj'asb�e���K��1ـ�7���@�����-��cMy�h�����.�M�/tbU]nkʴ��%����U�L�9�����<_/e���U�07��eR�j�k��և�SD�;�S[d���L��J����Ժ|����R+5|(�Y�\��]�F�ߜ�Q�P�����Yf�I޴���If�l_�[��n��N����x��zw���aT}�}Q�}��'���͟�!�>!�t�+���!!�oB�9�̚���M�YT�emkw�Ӯ��/`:��S� �(���HΛ�sUM/�K#���睉�5*��A�^�k���aTl�3\�j�=ݺ���r#��J�iK+��$�Be�Q����mi���Ϲ$]�����na�pv����S�Owb⮛z�x�:�ޠ�.bb�1�WMmmC��=�xg.�U_E'z�+?U{<G�zGs9��yN���^K��ؼ��|�#����4~��Ɲ�_˗�7b�c�7�b��Իmd&�4Q�$j��)�M ��(������z�O���Z����8��/����:��
N���K������x�K��y��ҕ��g��R�`��.b��wU��a7O=8�Q9g�Nj�,N䂄��a'��������U ^?�Zg�|��}��>�c@6_%:8��f+�Ú�\��m�
��h+,��v�̶�k�hOƅH�th��U��u�����t\����x�e�bG�Љl��;�l���X:p8�u���XmHwՔ�:l��%�=�#����@`��B�E,�o0yC�z��9�+��[�O�=3|U^��A�/�M�7�J��N�/�,1�
O"4����)��F�5,����&��y�x+��8�������B��W�����6��O��:��=�w�w?T���i�0Xlq�p�ܳ���w��N����P��j�o�}��#�H�r`����f�=�>�n����t]�E�v����w��ٓ�!co7.���)�F�BOA�rig_e��xlwV=�L9��P�l����e���E��]��Z��npi��v�Vw F�X-�}OeGܹo�I�>���حv�)�7����wf%��˻�M+�;�U����	��e��&)!���k�}صd�
)	iHK���؉ Q�JS�q��/���D�5��
Ί����%�����Y�����d��`_N���ٲ���%���9���Ӽ�,k���琂�4���g�f��z��`��>���:���"�юS�B7��^��T�/ʡ�6S�W��
�A�={� �C��Kf��o;#��P��cQ��/����vp���^����˭��>50.�)�c��y���K(V��[�,����׭M�k��(���.]�&��ޗ}��?D�P0Sȹ�n�xL5�L���i?e,���5a�eH���(W��r�qi-oT0�y�w����[e�g�}`)N5y>��n{�~��ު�/�1ܧr�;��a�A+�B�e���[a�b����/V�0!�eՒh��2��*!�M���Ӫ���?L���Z��H�H�rƙ�����-�;�E{�	�<1m�l�}gW�$c�	���e�a࠺fCȼ4XWL ���1R���<sm�cy��s���V;�����s+SH�ŝ��{y��$лd���:�g�,�<���cX���d3�G"LC���v‭p�H�ΎkN�׬U�x��=�\��ν:fd�_=��-D�Y�K�K>�0T��udl��h	���v��wvK}w˨K�;�R�x=�+65`�ЍU�]�s�Q�z��܁p�ul���HNe�[ZmN�r+�4�>�G7��W���y��ot�0���K7��9����	��s/��U�|�Ë�sj�{�ť¨`v�LX ka��6V`]�B�1f|�פh��t������7QL��h��wC����;1<�p|�˹4�_�p�A^�A4��gO]�z\3�"]�?��m��D־���Vɍʞi\�3�ʜ��������r�p�Ƶ�3��&��Q�G?���VF�?���M��_ȏ�@��x�]n��j�L�� 9N4�@����9'�1�Qʶ�&�;��h�4Ǚ��f^q(�n=4˽O.:v�޻k��v�#��_D�\D�E7|��ͣ��4���j�oE�'�7������@���%��_����~�b�]@d�g����B��H��>���@�i��*�%�Q�û]�����wn�x��/���ZCb��� 0<��C�Կvd&�Bw�\ISgF���J�k�$����hT߷���'&�ǿ(Y�f0�o�l)�t�s)�]!n�_2k;j{��c��1�����+2��v���W�����ژqz*Ԥ6��Zw>�*��<=��^�a���L�zU��ML��3h� ��i˞��˯0��jC���*�lг	�s��G�醲l&j#,u_x�:���=3��h�4�uˬ�)��yC��64Gpܫ��\Ql'_Yj���������y���o�7�7��0��XriVj�x,'��e�䪙9�J���N0��� W�!��^�i�F�k-��ؔ��Z1��ͷ�;u�}c���i��O�%���1:�l�S��~�l��nf�Xj�pk��@���ʹN�-h��ö4�ڰ	��4"�E�9�\�A�V,�g	��J�����5�)v�s��v�RX��WڒŇ�ή�p�|3?W���^�"�*��/�T��j�t�ž�Ѻ��szm���.F673s���1��x��{<*e�E�-M^�F���}��2R;�\��F�����&[�������	މ�����}�����P�m��Z��E�p����h���6�I�IΎ~����#=��)�܈8w������+�A�Sx��n�Y���%sqgz�Ɯt!s	�}2m��[��ړ5��
\k� j�l��ל��n:g}[���{�z����(�r������C�!�[z#���09�.C����y
�].���M�,n�Nݬ�wkL��D���.0����́ݿP
�%nLx�_�?<Ϻ��<��fVY�`Ĭ�o�vNᾑ-w�<��[g<��ƕ���I���>"^Ǽ�W�ܧ�S�+>��e���R�:�/2����N��:��(pA�҅rUq�H�zMt ����p��:����^��O�30��L�y�<�a@0�Z��^�*9w8�]>=�%� �9�7�3c�dW��W)��^OsE�;m�v�ю�Ǻڻ��?�9_�?;l�������%��15Bw�	��Uz������8x����A���a.�f�yה�Kk�xv�fע�i�ƭ�G�)|2��L�'�ߦ.�LR��U����Gn{�Ю�&��RcЇD�ȝ��t5�L�,�m�������xi��'��o���=,ѯ�ŤGwQ�B�GS���5��dg6�;�����g�q���=ٕZ�O�}L�sC4���wH��p?��Z���-�2fu�c����J����U�Y#��Ǡ�WA��c{3V��@�����˯4c�Z}"2x�]���Bŕ�����+ӱ�7�皍����+�A8�ղ�QT��^��ém�z��z|������J}Ȍa~����5�n�.��T�.K�޳㲇Lkj�v_����kH����T"��z�*ک(6?E�<jB��>�Zr��ߺ�4'��{d�1�ݼ�wv��A��{ߨH���M81qN��=��5��.��f7$]���d��ذ�U�����O�qW�i˱�=Z��:n�h�ڡ\̼����t9b�{�Aһ;)��"�c &�NXcs6�g�>ɉ�+m�bf�\��D�����<��+�Í��QBh�%ӌ<Y���H��M�[�����w�]�,0�o�)o>�es'\�hT��h]M�Q�����J"��GىU����f��o���ƥ�h�GϚê�π��@+D����ͩg
��"A�7p�8�k,BUR�kz�`�(V�� �ӦV>Pmͳ������L���c��h��}0�3�nHm��V�]("t���5��ф�gƻl��ŝ|�fkX7%�ڎ�ޞ]-Q���D*+ݗ֩`���Ų�b�蒎��e>\�z�����]7��WV�L���7@v̅�2S��G��-SmWՐ7z�m-�u5���k&c�=��Su��s��e�L�ܫwˈe��$���e:޶��5+���6�V��7��8cΣ�q;ZCG7�W�������v8�\��&�10rqx9��i3m�͑��c����u�+���\�NQ��.ޗ�*�˔3Q���.^����FP�|e0�C-T��(*q�wY2��.�@9Y�m�Kp[X�\���J6�ܨ:������z�"Z� ��o�r���Gڲ37�bÐ�F�wQ��
�˹��vA�n�icf���i�A6C��^�|7�K�x1��Gֹ�F z�<U��̷w�(3@��n�y[�♈7zC�5�7�B�[.�u�jV_h-��9�%ض�n�,��(�Dխ8�)�`}��t����r�@�ۦ�׋Zeǯv:�N:�{7�����s�u�ƺ8m���VB�V��R;	D.�U}�.G�f��+*��Ffk��ަ�,Gk������c����s�ߌ�yV�,�a�"|�Fi9z�9�gYs�ͦ�N=������b�j���mk�ucp6BpqY�'�tR�j�η0����dYG2�ԙ9�U�5�%a������ޙT,[�M)� W����b���C�S��'��OHBv��]���R�QclvU�
���	��Κs��5�Z�53�;@�q�d|ٺ1JR;ϡŴ{��t[��1mm�c���4�h�V�m�-��u���|�u	jgZ��X����V�K�n�����(e'����\N����t6�Df���'�:�
��Nf��&^Z�ɖ���6�|F���|sㅙ[��&���f���b�|�YD&o�Be�'؊�qb�j�}e���ͬ�'NB�[A����Rw֍�d��g�r��4,+�N�۴۬�-��]������J$��ŪWf-������) �CZ�x7�s���-6z_ZMv;�S�[\�᝝w)��vn��J�/�H_�SF�\��H�*y:ӣZ����Q�s��[cN�s��󞶝���u�"�1�&����Ƿ�j5�cjqM���6��F�qȎms�y���j�h͊���Ͱ�h�jB��}�g���q�1.Aʘ���#{�r��9*1[Vն"b�h�3m����nZ��E��������j-��E��w�U�MrE� A �"?"���E�Gc]c����V��n���ޞ��w�[��k�r���h��:�u'�cUQ�B��Ξ�n��Kǧ�Ƿ��Iv+�1n"RC���B��(!��3��E7Vy�u9����{
|�@����4'��˔��m�k\��n�8tW"�������>w�Iu���.Z���+bأN�Ӵjձ#b�cc[mD�EQ�x�~�^ߏn3F��5��nMA��uj5���p�.ᱢ�GI�EԜ9�g�t�"�x�ry%k�3�UZX��F�2[[f�4j�LHh���?8(���mb$����a� �0��h�`L�DB�B����	3J��ޚ/}{���O���K�Sn[����N�K.2�h�xқ��I\�[/ik}�S΁����,�DR@�!�DC
8BE��q��&#p� ���bq%��B#q(Df�)|�A�h�jF�P�����:���u�uÇF�8ug���G��̤�L,��+0�ȏ}u����.5K�o��b��+D�F�R82(���P!�$���i��-@�\�i�T;�v9�9fϢɞma��G�x;/lw$bʊ�9r���H�tb�d��Y�~j��8b��<�4����aE8��#C�ΑBMk9��L;v���5�Yڛ%Xg��`������.��`�2�82=�qP֞�;u��/o0E�M��J�"䬨%��.b��c�C9}hw�O��8v��R1U����֊�蠤T��z�n���C+�ٞݵ����ߺ�2�W%�����o@�ƞ����*5�Eŷ'{�ٱT�8"�9��{ڗh25]3c�Dc1U.�hͻ����j���yfE�pS*��T�kp��xi.)��}.Ր=��j��6j���tۼ1�|sX�c�Tm�ޝwQ{�[��5"�!R���_�0��[ׯ!0�/L�~�+�;\�Se
���R������1R��C��x�T#�@�8~�%����F�߿%�\��Κ�;a2�b�O�6�Jv���c�wr�s�m!6�U���N�0��v\��c�6u� ������b�L<hk��~8`�����73ܱL�QQ�%���ΣeQ����{�p܉?>��{�V�U���B�;�I�:v��+fȜ����&Yol����N�}�V�o��D�a����y�H�0�	�';Wv�[o3A
��l��AT������?���e`�	�	�e���m��Q��U��y)�&�X�{Wr7Q��|mw��0�ƨr�n�!�E�A�i�.L�]�3^\d�5����ͱ�e���t�9cl��DP���zwƉt˞w����*��Tt��ᷝz�j���o�zC��)�4����S.�Ш�Z��?3���<��6v���os��PI9���������k��A�o��4.���Z�a`�%�cý��[m���#�m):�����΃��h�(�4&#]4o��i5p���Uܨ��݋�G�C�_T�p�xz���3W�X/r:k�D�]D�o�	��X���O���;w���;��E�&���8�ޮ��,�uO��3������.�z���tW�}�Aމ����CW�:O��!��yc�6���sSf�X����,�i��~�^-���v�g�?�g|����ȉ������k�}�:�13�`����mkS��}�s���K�f����2���Z�M��.�Kdǿ�Oջ}XDD���d��.��m�nG'ֱ��Cu�R0��6Ο}�"[�4�3���3Z?�d|��5u�V1���c�MP��[�~r�{2��E�]w�Z\�r���'�K��¢�#q��x����F�MB��+/���⓯T���ld��%]�A�)4�ծo�[t�QwoR�|��r*��<�K�~�_�O�̃00$�2��y� 7�{�کް��(�����%�'�ؔ1q����n)��u�>��D/16�=#e*�B�(l&7�q~w�U�\0�wmL���)��ۙq�RͰj!��Y�@W�%4�f�n�ȡ����3��b�<��e�0�_4Z�6��9�����v54�7\��ʍ���O�tb�B�Ye^�n������n�Ɉ��	fJԳ�\~��}vC�D���t��q��ļ<:�U�ݒXx�ux
�e��cB�+�:�{���jb���#��n�3؜�WW��8��l��plvC��'���It��9w���U���u��M�C���=M��Oc�g��d�mAڐg��	 )v֩Bu{ &�d�y�,)s��2q�� �6��0[��N���Ǽl�YJ��G��yT�9;�C*È�vO� �k��Ĳ��l������|lҤ��Л��K� ��{U��ǒ������=�>!��� D6�-L�Iy/�9zR9��n�9��O�2�%���PZq���ͽcAk���߃�(_/�.v���3��q�k���4�u&�o�{�t��ە=�{6)�cYD���JÑ�\緦�ww&*x�u���:�i"I7M}Θc�WV��I�7G$��9YI:%�x����B,p�v�Y��z�0�ؓ<�dj<0,3��͡Q9�_Ϫ��2��3L�2��� �x{	kG��O+[�ķ�t�M�I.�~��XM��|�`�|`����O� k7�q�9f�{���X10�������+�"+��_�f����qA���w�$;k��e�<E$��So9W��|Q��M�
�Q��_��
�k=�P�{��#����lǘ��>���q��Iy�g�|<"Q�z軤w�U�v�e������pX�q�E{F�P�{�;h�9Co�m4��yOW(�u�(~��_ �=���ZIG(|��J����偓�hp�Tm� 5��uq����	!���am���Z���||�}T���
i�\r�E��=�Of��qQ �S;����˚�{6<O��fOI\�y��m;	]���e���^T��.�k7Yxb�v�{�ׄ6/L�"��QMb�b���M��۶��[:�^[8�>��15dU��gn���<ܡ�@b�
�-	�_��x6���s�yO�b�M�PJs��ٵN!�=KW^v*�<�.�C��}覶�BR�282�dk�����Z�T[y1#��㼻B��jKƋ�km輦���(���=fV�pL�OI�.�x�S�}*�s���o�H��6��sϝU�7�&8Q��-=C����?O�s��C��m�09gi�� ���*a���t+��ge��4v
�;��%=:v;���1�r��X�:N�UU>������e�	�	��I�}䣣&�Rx����~|��|��(gŠ�%�d�E��X$�:R�`Z��%�����������.���3_G[�8�J��%;����+U�"Ћ0��\�&�/id��+(CH�/��=���ʢ�<`����/7S�״2�6��}�׼���L�&�Y���]:c[
7@ǹ�s���Ơl�g�x2��*��, V�N�oD훇%
�<��XH��;^�.SJ{	,��{E��[�vڈ���d;��=lƗ�X���s�QIս�z�dU�I8�]$^�5}q�}�>=	B��{d��~"и͍�WӀ�=!L���)�zcɡ�a���Q@GT����I�o��M!^�S�FZȗ}P�r�N�NV�Y��L�r�����%����<��`���1���/�i�;C��~�uP��P�/�y��4���:�Xm&�\���0�{�#^@v��^���f�r��Y�b�n�rdM�?[/!��\�iކ�i��d�k��t��N�	ח�"'ҧX)�e����HL���6t5KA�=.�g�����	���N3W��vtb��a�3��5��B�\������
L��o\�7z	�"�Պ�t5}�v�1{ Hv�-ÐU�\dlk����=-��?b�_�L��K��(�Oͷ�_@���~������	��iR��jĊ�&u�Yo�!��|��5F��,�o���	�aFaԐ�LL L�L
L*����{��?_<�����%��QV!f���7X��w���0��E��	�xgt����{�]F��wc���G����De��Tu���J���A� ��+_o�e
�ڞ��JM�)�cNHӣy�Q��~ʈm��3�Bw�{�Z���s�\���-uElnu˺�*��6��n��C1e9Ie�F�\]�چ/!�S=���nq��)�6Ҝg/�\��bg�Ö���\ͱψ>D߆+�V�3���(�t=}wo54�̑)4cHbv�a�	t���؃�u���)����v؂��,��_PJ}��G,m�S����r��]���:�%n|�pA����w#*D�~��u.�Z|��S�!�̦T���b�2<�͜T�qALs;n��*���hC�mF�<�j-�x�ʚZuy�n/m����r*�Yaf�_��Ya�r3l�9�aU����/N������W)��t��$0��a�7��H���z/� ��
��F\iޘO���e�Xl���ݸs�j\Z�*S	�l�k�`݌�E~`�����f59�Q@2��-���dXCN�e�̺��Xv�������yq��"��dU���̬�gͻ��;���vy�&�"]>���Q�Q�Iu����'R�9�$����Q����\1�P��4I���-��������yr�3�O�Ӄ���s�Ѯ��v�w� �Ȭ�,�,ʌʤʣy���y���<�I�m۳h_�ʌ�����6�U���.�Ǚ��^��L6�su��K��s��ϥ��kkfM�2�%� L��6�Г2Z�愣�9�w�|��y�����n���9����{��z����ZD��쾘g��褏h�8q�Eo�bS�\�^W���h�09�=M������&es���jDG�︡�ya8��h������K�{��
�`�,��6���ڜ+k���e_�3��~�,������i߱�߮���>r�#ϯ\7N�L]�A���$��AvTD~�����Á��'���R*)�a*���®����_�M�����*J�V=�Z��+n^G=;�3[[[�j�8�^�qǼ�GF���!ߚo�ة��d6:m�ٽ,��Ĳ�J�������D��u�*����&B�� Q��z�ɌS�Q@	�#i6�i�F��Ɗ; ��H�L�)�\�Smy,�`����h^�s�E�棍���Ϲ�AB���"n��A����睹�`�U)��H	\6թ�ܦA�N'��v����of̬D�R�*�a-�9틮Ls�V�"0()ގ!eT��(��ηW9q�:;��C��YS}�>��c�MYΤ������D��=Z��J�mr���8L5�WfS_�eu�,oet�h]�u��u������|��؉�`e�U3*� �"3
� $��s,dR[�ñsT8'��1C��!6��M}����C��^����Ӭ����Mod{f�y,vw��&7�K�s�
z�妄�uAi�G_������6����ߍ�����wڊ�@&����[�k��M��6�AQm�C�û��k �ڇ�D���m�;���z��"7(M�w�\��ke�C/�aA/��!ӅhT���l�x��"qr�鷁����]�,so�������C�Mo�o�6�u���Ժ5��E˴�C�s���ߗ�ey�Am�@�m'���g>&��R%�=z�}q�����L���������wT��5��Eb�O"�*/Q�����;�z�C�,&#��ύ�w��~�a�}ө�$dt3VA���U9q��7w#�D~��H����g�� ����@��^���Cv2��:&���G���|�)������C����˾�	3��ə���@�߯'ӗ���m�O5L�Jz�y;!��N��6�)f� %cPz7.�G;6O�tиy���oߎ�,�;�C��*1��1k7�N$R��{F���y�1Zɘi��~8~=�{��?O���b.�U����9ǫ4Ga��	a�|��Pu}�48��=��>��Rޮ�>=����rCo
|�͋�(8|����k�u�zŭ�k�:�Ͼ{�DO�(�22�00�0 L�__u�xn�|���>�=�y?2��&8�b?�D����G���ǡ�b����r�ͯID�PՔ�zx���e��|��]ɀ&DjB��u T\�k�&v�+�p
uOb�41j���o5[&�W�M�9m
[��g��{���qU�,�H1�N��-Z�'��\Qp�V���=wBe�cR~�J��D�V�K�ts5a�zdNL4�u��mJ�؟�f:V�~b�:��|�������K]x��ͩ��n.�#��uS^�j���5.��z;��°��H��h\�=<�}�
fg�;P�.�-�B�is �=�f��hR5�W]/6ࣴ!�k��'�sԹ�	S8��$ZY����a���.���]s?��|�E�B6�;�i��P�֧m2-w[ЭZ��At%�k$O<�0%�m���eBd�ts��׶1߄?y:�P|���:��V���{���� t��B)��򇚴����o7h����g�@��l�����M��f��-��H;[�����CG��?5K�F(zO1�Cy���S��cR�E���$%=t�Z����CZUǈEo�ә���E�N���h@l�}Q�ޫ2�T�C�m�[�7�5ֻ��zt��R��90m��`�}�]���OV�]n��*����x8N�*�bÛ]������\볏�wvm� ��3�`�D&E	�B` ��{���ߟ���UۨFA�o���r�Y���iwn�D�uo�.<�ƷVh'h�TÚ��z��-��B·�c�mz�qA�	~z��;i���=p�H��D��ԇL���ҥ�ld�3i��Й��j<�mP��ܘ�MA�S:z�}4�>zL�EoSUS��c���WnB�lǰ�UP�9o�<8��^G�UHkFm�WG�Ti�]�x��Z3W_�i�
rxi��NnK3�Ac\��P!�5N;��5��i1n�mWa��V�3��"=����DY�/��)� �J��!�?Q����+:�u�F"l6�އ��)@/>��s=8�����ڃ����VnY�?��h()�&5�Y�[_�Y3�����_�L\{�6k�aɇÚ�}�<(��ncS.�4[z6��}ŜJ|�v����4��cK�e?��]�&���*d���"qP�zWr;���=[㸦���1��^�L�c%�f���}x�.Ոt� ��f`���+zx�Ni�e�R�gR9cOT�Dl8k|��<=zQQ��P'�b�v��Y���6�[S:���� ��XO%.�����@Fqӛ���8/;c8n��$�/�)��R��v��/��΀L�y�Ԯ7s($����;v*J��i�!b��'���6J�ۧ�Q�JR�ɓN�@��WK�d�C�]25�,�Zث����	�_�(]�N�x�H�ꙹ�o,��<��}���{��P"�����	a���QәKT
�"�־-���0@��oy$�d���لv�lj��Ŧ^�kNì�L0ؠ�Am�o��@���;3*�4�1M?^d��Bm�`�ڷ[M��]�z޳L9�a�\�6��0+�y�=�T�y>�g�^i�J��
�vN��Td�j�ܯ�n��ӽ˅v�8L�׳r��g�tQ�e��oF����+�r��.u*���x*$�H���(#K��9�X9������ףͩ��Z/��� ��_"gllB;�m�T��j����
W;��D]��k����wo�5�Ұ��|�W3xn[������4p�j�=%�o'%��@�����TO7a��k�h*��P��S�{acvf	�˓��V�!�,�7��IV�et�����7���t#A�R�զ*�y�c��_�尞�TɜD�8�wn� ����0Y �%��	�ie�+%��ρ�ľ�ۈv+f�ف��gv��Q'�`�t�q>����6��[%ptЉ��k��J���cq�HBӻ��1`��l��!�.0�mD���#yV��fi'ȤW��$刌83� 9J#�ȃ�)ѳ�(�F�BY�������x��8-0kP�CyPECNʼ)�Ȟ�u�կ��s9�^��&IY�6�7W�g
�Oa�\��2����vйt��.W�qp�d����#"o^��)�%�L�<�y�0���ǲ��pg
.���_���$R]���>��\��9�>X��^�����Eax_s���Ufr:���T�ioK�At�hL�hpn ��X�GO^����d�
%�����G�9�Q��Y1nR�w t���bΙo��Ij��X��N�ڻ��#Ӯ��1��5%�K�=�$rn�=iC,�΅ԙ�ͽ�]�a��V��>���L-�n�K�D��+s(૧&��)&�݀a\+O�2����A���+��f\�|��)`z�7�
�	�y˯o�d�1gvl�J};�l�H#A`=���g�o�x4]v�t���k;tp��A�\'SG��!^�FPr�s�����td<���	hopC��e��Y��`��Ֆ��9]��i[ӋO�Ɍ��|7�����7EE	�%�fXI�ޠ�1���y;E���A|x����q9����[#׮��,q��7KG�/��|	Һ��D��N�z�u���sè9
�m��kPImۄ��5���� �v3X��V��_���ۣ%��4<�����5Al����61E��hؿ�*�'\�#�bۧ������9�;|�r��E5AG-964b��mN��F!���*1��r։ыb���x����"��#�ί�45�=Z�q�����(�u?'��i8kq�==>=>=��ͣm�r�M��jcW;�QA�Q�[gZ���N�T��������m4SݬX��\�(�h��<��<��nq4r+Tk�%'�������s@Z�4�P!B�B�	B��1�Ul�b�68c��3\cݗ�6���ק����%�w#�� հkZ#[���g�p����cc_1˒��b�ǧ�����.cDN�(�;�8?Bu�ꨗ\��E�g1[}��厏��S��TM@k壢�m���4�I�k�Yi!}
$ ? `BP�����" @P�)�`s������*�?�=��L���l������}��ov��Tmd�iz�U�`d#��)�`�^o1϶���?l���*̨̂̂�#H���}��ݼ����W�Z��|S�9hL���I����n/`�Jm�j�9���Z�*���S��l9��}ĳ�b����9��m�yO6��xhӋ4���ͧRG�3�Ee��r�������pw�C�w|��	��ߜ@�����+����F\Qݍc��E;��ݷ�C2S�L�,%%��:k�;��ƆWK��*���C�����C����𙻆�X�g�����wp�5�ݙKyI���]�zY�x��%圾}�Aރ\�a1��#�lP׮�/[�9�iv�[4���66y?�/�Z	�h�S�ğ���b#���$N���ٰ���q+w:d�����v/�,6���?N���Ë�;���?z�ʏT���.��,B&�s�u�Rv~}Q�o������A-��@f|�A����~����t=Q���ʦy��چ���Sl��:a���$5�lf�<T�o��3"��@��!�rr7�j��T*���ݵA�*���&q�<ٺv�v�O�4�ڂ�Ú8TS�v�(��+���мfߵ]���d㛲B7w�Y3t!�)wj�o+^�NTݶ)l����ñ�m����c�tV0��$I?�$I$Q�v��qd��W9Ct��콢�oK�.�ه5.1=D��x�}^��5~��f��E��;������ Q̨�*� 
$Ȍ� {����������G��p�h�d&�
�N=M!��(Pn^kœ&��f�n�~��}��߫;��A�5�D�6�Y�bZ�T�z��m*���wB�-�xy�f\���jF����i3$���wf;`�36�[,��}��Q� �ú!2�	U2/x��i,�a)8�������kwm9�s4�{�Zsp�Ś�y���,y�k�h��7:��ji}��b�M݁*�ދ��m�T���RW�N^�mEN6C׵ŵH��(˰��	��&�_t�����j��/�ϧZTCM���6{t̽2K�1��ҝ��*��u��w�wO����s ]���Y�Lë���6����!M$��9�Y��IE�1nw�C-ps�)���fj���KyaG��C���Ώ]ݗ��.Խ�"Zr��Z� (P��y�:���f�e���<=l��!����0,c˶�F:����/-�>�3MW��7f�7*+��$α"�����P܂�yhL��既9���ye�@K�bz�='�q�ccg��1�n�DdtO��g˔:��3�l�ǝ:傸�núu�3������.�+-٫S;Nb��6+�´am[��3Y����t5ȗɨ�;�J��>:��]W��0^�;���3omQ]��>;E[TH=�Ȩ1Ո����]h�ȸ�LXk;1��T?l�̂(�*���Ȭ¡2 ���˕1^�?��s��J����	|-���[��m�C��a$�����O? ���^%��	�>�!F�c��#�8���tG�|�B
���Y����n���-�N�}�o�DA���I����X{��j!�ߞD�ǔVRm���ͪ�:�{�]Չ�ո�9�r0ISe�7.�����_<4'M�1m�1�2����&�_v���	��y��o7,f��g���Rp~�I��KH�t��qHq�wa���{�8��T���U\S������b���3k�Q8��%�J�8�-���K�=L3~�����/����7��J"�π]@�ԥc��A�HbY6_�ʦ�KhT�Ȼ���y�Z�#}o�zջ� �2ؗ{k�_�Ը�0)��������=Z�O��ѐ��4S�+��}7�Cb�c�Z��B��c �������.�o��>0��;�NI_������7���=Q�N�d<3=ډ~�-���Xα��5����Yx�K=��)��� �'��,މ��A���O��]�3/m��P~�����R}�J�4�G(mɿe�h�s�1��/\�����߬h_��f���l����L�Az�S�z5�F������C��Ӷ�v���Nu�ŹƷUC��J�̎l�P]֔�Q7��`��J���x7�ͷS.���joV���O�syiݶ����ν�κ��� O� ��2�L� ��0L(��^=�6���������[��ީ�R��g�[���(��;w�C�g���X�Չ�6WqsV�����~���C'<�_�ly=/]�)�X	,��E��'�2wL�V�e����|��s��4�^t#J��ˢ�G��#6�Uw*,6��4'��>��|2%�g#nK���5�ᆶ���"l�q���ZY�Z�y������+�w`Y�Ӝ��7w�8��6Y���:K�yt���
�$b������c�$kL�Uo����:�:�e�k�X�~��Ǘ��OK��kV|<��D����o��:k�^�n���'��+�$��3��x���w��j�%��B��||~~t��G�?��K���P��9e�.ݭB"c�(��\��N��eF����}�F3R�R��u.D=ƽ�wYwz^l�\�zǗY"c ��z��.�|�����9c>�1��D�L�kf���ʊ͞Q����*m�Nw�c\��q��Uh�B_�枘@*�z�e�jK^'�T^4�R�V�[�t���VB�8�m��sJY�sF6M�����O��C;�<�J�iᒟH�{�j�PC�y�RY�:u�;���3���`�C4�zmf���k	�3.��Ls5p����f `Lt��w ���}��A?l����)2�L  ���2
�~~}�����z��[eЬ����71#���k�~O�~�4���!���iL�˕���n��-L��c�xb�߻<�(iQv���G�Qv~{N�k�P���o��( i,iӛ���F���ml}�����=>=ʕ������
K%���C`{����N��f泞�4f��h2�C��C'ÃE��b�/Cf9=q�e����"��f�2 Ɔ(�
v��KH�p�n�񥭧�D���c��d�y��L��_���ݪ9���YRH`�{:�e��^�?G�x�?>u��c��G�Z~;3��8�M��>m�8�J�x\.��-��/��?0,�-E?�C	g����r������b6.���de�V��zÈ�Ւ�x�OIGs�����*5�����h����>��}O��zwS-3Efk���[]Ag����n�=q^Y���l�1L��0m:zG4��Hq��5rn�\I���i[�^g���ԗPp���Ό���8%�<L�F�I�^d�C��H~��{�ߣ��:5hO�r��E��>�Xb�)�)�]�Q�齓gT�'U�"��0��9��}�8�������[�aR:0�ӱ���:ʠ����B�z��[���5�6�9v��vd���m��0)�̹]��7��|>ψ��"�Ȭ2!�@` ������ ��؞-�_眑"2>*����'׿���ͤ_܅���[�c4���m5i2��S��uu��=��גeZ�o�`����Ϧ?~U��K����p5�tAl�k�T�~�'$f��vm�d�B�����s�,�Pb�?��0���SQg"�ǟ7\@p���ݘ[i�0Dkmv�<�k�@.�h$f��������g���9Y���%?<~ҢA�TNlg&Y����f���Rە�
��+���^J�V=�V��[r�Ϻ��ᦞ�a�"э�9��z�
�����f�q�����Fm�_�ħ�	N7��̱k�`����u/y��������T�LS�-�����ֶ�x,$��p%TȽ��m�,�aݛ�ٹi46�b9ս}j� %���]�s8��,��5-�F�<��K�U)��]�D�?M#��t���	�n�r�wƢ��e�f�)\�	��h\�/�CϵN�3�����q.����1գ��#vV�A�W>�/ͼ
��>�p�8��8D:}g�i`�կ��vw���]k������׆ɯv5x���*��g{s��N���N�Ü���;��ؘw�iU�S�q���v�u���@���G*�&���g_C{�GU�;/z����|*S'�G{�3�Ҫ��+~�r@N�����i�U��[��g%����� ��
�,�,�2�$| �>����da�m���W��?uQhlL4��nD�So�$K%3�4JA6$��\����O��A�����̸������L]�6�Ϛ�Լsx?WqѶ��s�;�wh�iB�[�̉i��j쀡E����B��*FV�f͗����7������W��<�R�\�6�]��:i�n�L���AeyڧI�9�Q.�L;0O�(��jq0njB7�-�D��
z�sa{Ǥ��ٵ,����{~7��)�����"v��TN�/!ʥ��;��^�6~a^��X��T1a���(�tt�!5U��u�u��)���#�6���^AD_���$���	��a>�q��>�l3m�=�*K��z�g�����3v�/3��#���J�M��%���~iw�������j^Q����jA�rf�;4��O�E�;B���q�v��Cmq�a�U4�n�=s�j��:���b�<S���n��>KYk��?2�����N/�W��p;`����׉�)�= �Kej�v�[�4�����ީ+�iP�x����U����^E5צ��u��}K_7�ƫؖM�\�eu�X�{Y�P�nΌ���&��zv�h���e�ɣ30`���ʲ6�vtMDe�싞��O�}ݰ�;�d�e�H^���"���˻��ɕ��7<�Cx��L�3�Q�UǶdq�SZ���(��-�}�7.�����}���Bee ��Q� &@	����_�R�gj�S��HỢ]�+�aߥ�'	�R�^煏�閻��l��&�t���|A)�H�c�X+fo!�����[T%,�q��ԟt�-�4ݩ�wg�������}����&�Ef�U�5�#������l3<SO��,�s��63j�KLWLi�Ռ�r���MCW��H�y�R}�	P�nF율a��<ь��LN7G�	�]�km'�R�4�o�"+�;P��R��tO���}k��-��@w}}W1=[\�P���ۇ`����r\���%��?�U�{ |�<���o]�̚�&K%�'�줎��x�̕3y���i��Ɓ)�Y�,It˞��L�΋���"��Ia�k:)��T)�a��
k�*��L�dZ*y��S?��C;��36�a^o:O͒�Q�
>Q0:+5K
P�:G��n.��*�5,��'�L��tW��N$N?�[�?A>aտ!���k<G���F?k2��:�gӟ/TT{����(�μG�TI�h �wЃ�jK�u^<yۓyW��:�-f��-�r�a�d�zԕ4��f�����VO�{h>�@q�i�Y�N��e�OgK����c1�'��6�U�g9�Uq�t�E�;#ّ�2��ޕr\�ֻ)-i`���X�j��o>��=���μ�{?j��Y��Y�ad@�&U~�X&X�:|�=�H�f�ɽ�F�m�x��^&F�%rZ��ފgO��	���κȾ4ݪ�f��
T�	��-��z2����y�W�Afנ8��b��gT��q�2e�L�k���^��>Wo�,��\(��)�_1ŵ�"ԻG�!2��P�n��klM�ŚԺ���A�/)�w����!��]�F�AT�["�R���z�7-�����g-�oWKWch��P��n�Ka1�WB��V����&!��|�mr�?��Z���:���ŠP�=�y�;�Z��mY�̹�R~�b[~=������cq �ݔ��7����ou=�.ʈ/��/Y�V1=��N��z�u����R���%�Z�J��7Mn��`b$�T�u�xm�m�gdǢ� �\3Pu��g��q�d\�{%uP�n���]v�[Rl�ý]��!�](���꨸?r���_��}�[������p�e�6�gT��m[�M����RS�� ˱q��]�!���	��n/X�m�dˆ35��/�"U��R�g�*��r:]�/.ױ�Oa@�a������K��\�t*��gd	�=Fb-����yٛɨ�Xyݳ-լ�H;郪s�+T�{�Ъ���3^{��{���%�F�\��UHtb�ҿ�}�W��Y��I��I��������&�새N�R��Y&1�8g�gM{�gӡT������� m���ؼ��=�ŕ�Ԝ�wf!�ǏY����䣹�XJK	�ε{��zC����	?���Ӿ���uW?oM��T;=��B^[�FI`Z�zJ����ȥ��q��K�9|�6�8�by`y�6�^L�ْ5Ba0���bӒ�Z�c��$-d�4c�ԉ&��t�Ƣ�������B\�������3��x�(�ʧ�}�u=7S��5 \�=����[��;��۠i�N�Y�}�薌r���D(���AO@c�8�.��/#��lW���*�n��Me��q�[�!	=6��6Ξ����v��o�0C��T�\�\^8�>p-һ�e'�k����d\kt=�A��!#'Tۿ��F�;	0톞%�C:j�=7�TS���W���e��j��0dj۟ne���8�!���a�ݡR��<0J�`�<=FI�p�?*'��.����B�;k�'�:�i��J/�L�_b�ol�f�ߡn�����%�eՙ��u�:��K+5q�z��X�2�5�z��+���_.���iu�Ǚ,�A�WPb��,����*�=[�g.:�V�z����@��yO�V�Go w�*�d:�ʃ[�I���e�>T�u ��"3��n(���:�]\o�}Ϡ�VK�Վ�*�Kĩp�z�99�M^l�/9�l>��ft�oq;&=@!sp����fDF�]�%ϊմh��]�L�wz:E���E���vG'�ͳ��"�g���9��*�}�R�h�:+i����2GW[���S<q]ӐJ]Hbl��OMJ�\b��O\���D������g�\UcUr��Y-&(�����i��1uLY���m�}λFJs��N}g2��J��%H�Zbn��h�\	r_ٙe��5]
�Rɇl�\�E�g;�Ef��$��l���v�B��X�&�88����9)'O'�9��`'rk�PVn�^�C�V�f<��i�Ԗp� �5���-�me z��K�l�Q��T�)���{A�v
$P�Ǫ���[�K�H��i"��[�a���%��n�j�r�h���>��*��p����t�T����˥α�8oF���L(m'��(D�j���5���-�1�1��r`w[��Ճ��5;�jգa��s��k��.0��ξ��W]�-�V`��M� ���gx��^e���@�ġBQ�Rf�5
� ��eE)����`'{�V\$D!$�i9��u�����WĎ��ჸ����i�WR����4�����F��\�I����ZZ��;���=u ��z�@��l�m��ܶ�ɌBf5�g+�V�,�l��:�Z�QͼdCr�8Q*r桺�-�J�@v�.8�S�|�|�ז��к�
��{f��;�2�(�9��y�cc��+��;���X��>���$���,�gT�wϥ�PFGو����Ұ_��,d]��^�э�B�h2�Nf�6�7���IDtAH��D���/x޲��r��nsX��m�K��-1�h���2Cs.J2l��u�ȶ����j�4y�Hk#L[��"�r�7xLۧ��*�U��Zr���Am�fAW�������Ns{{jĸ�����pGk_7ct�w%�2�0dέ���AP�Ĥ�W�q��WY}w����m`��|������i�mŏ]���.�wL&u>�V9��;�O��8�s64F������.��Ԅ�c_R�y�26��4��x5�_u]�p�6S�v�,emod�8=1.����,Ǭ#�$:w-v�љ�"���#�),�Sin:��.��[�]հ݁N曘�(�ow�%������"�Ըd{���<D�?|���|�����?'�Eh�3�r���`�m6b
��9c�<#�4Q�[n���������{'Z��N��xpb9<����Em��:6���m��oOo���w<�*#E���.a�T/&��l8d.Yѣml�	������ۻ:4klR⢃Am�T�V�I��m�;ᡣ���j��6��"��������q�6M��Mk��ä�i���跜NW7�Nq�f6����QT�����=?^���|�흝mX�T�����Wv&�q��h���3���K$�p&�����������ÁUWͫ��:�Z�r�#U�� ֊4b��E�DD�x�h.m��[j�U���5�������h�>j�[Y-gA��jh�jb��g�6m�Ul�Ӣ�X�;�L\�k4o��Ƿ�����.�������,j�m�7�f��Z
�g��\�֝ѧU����_'W2j���M�*��d��'Y�ۗ��yrk�.�I�X���b�!��u�gAD��G�$Xa�I@���	��
��"�'�F	H��h����,f^��WO98xK\[���+~��=�M4n�u�X��'Ig[hQUjF��ǛvaI䴝_EM�W4!� 02	Aϙ,4�-�M��A�>���d����6�%�C)T,IL��4��I2)"1Fa� ��T�U��U�T�T��{9�������\���U��DD�
0��H�ІD��K�#�;?�4��ja��u��W��6�X@�)�Ī����+?w5!-�	�f���N{:հ��q�}����C�q�k�_��M��Pyٜ�a�Юg�i��*��Rש*��gho��{�O��
�`�0�5�@|3�)�i
�-ogަ��z�y�	zW���#�IJ�濿S��th��K���uh��4���묩9�Q9;Rr[�70��T�t�ky�n= T[sW��;ǳ`<(mpBeZ/jO�Y6�C{�����)������i�]Rݎ(䣛�çhT���l��Rh���h��ż^а�B��y�-���-�uJm����kk��!)�S�F�8쬪���>��3�b�.���Dj�4�o�}��c cO�6y>a3�lX�R���Dݞ�����$���[���+�~�����Z�9��H��
az�ϱH���hS����X�S����(�/D����/�b�;wv�Ǒ�v��!�G4˄T$/������.�o��#�C7x�9�۽K�	�N�7�4M�2�7�B�r�YopC�'8T#E.��8���:k��mR���uV�g�o����������.�����|f��xZЇ&�G���I�ϫ����JL�L�L�LH 3"�,ʩ�}�y�~�E��=�W��~<���|�mD�T�q^sr��]���/���
S~��
u}U��~=����z&-�l�|ɧ2�ݸiڀ�҃u���⭧���O\�ڛi���9'�]E�ڞ�~C���
i�(%�MG��X.-�Ζ/ܧԙ�μ6ϭ];t��¥4	�§�v��߁�k����&�mU04�˄�S輄�Y�dڴ��(����m�Y���%�*��;�O8e��v����@w�v�U(	�ԶGW��c�D9f[TÜ[{�v�l�%�W�Ȧ�*�1d~�'V�����Ε�ߘ�΄�uW�h\]	�.�S�T�;����|\�=&\P�2��%	��b�{V�kR99@�z�{a}���MO- ���/�6N�&���f�3���F����/)�4���g7t܋i��Z�/��z�L��o>�`��,z��}oZk�]��H��R��g�[�|��b�זiJ�ߨ��W߳�I"}a R�;���<1n;�'�@�Z}�����r�Κ�3�/�H��1��.���'!W��<��s�|)�9��E����߃��a��^޹�r�f'Gb9s)��[I��� _�G���W�m�uwu!Ն��f3���8�'��b�]v1^�˜���E�	s�;_,p�	a��ܹ�>]r7;�}���T��0�0�0�0����"�����ϾXT�}��=�D��;0�|}��8�&7������~h���ߺ�Ya�k=];g�!�>G]ڎ������ ��H`�_M���ΰA����������y��hgw;�MUx�"�n�^^'i�ȶW�#���zĽ���.�����ģ|
`����?s:���-ſlq%hy�;�C�=�(�6�Ls�A�.|�6�p|.�U�:@<��6�����@�A�)����b�ö�6{??��3m��]��J`���Ν����^��Bz~7P\�]��^Z)Z�3�%�ʘ<���$��͞�L��
��R�Ɲ-��5���6�����2*m�5�|]�W��#]�ӟ�"�Ek�P/[�8�9>��Ӵk�Y>b�؁��K���K��JsFχ�~U]��H��4�aR�P�6d�2��=���s�c�Va6ג��5V��[p�������3�w���	覺�b:�ʢw�qW "]�Ưe��[^�e�e�>n��Eۊ�F-�+t��n�/N�����2[�2)aZ�XCƍ%˺�e@�L��������Oeb�E�Ys�7R��7�ؐj�Ӑ5X����Ӛ�Kv�eԵ�#xg^���u��gz�m��6��뾚4�r�ׁl��GR=-qF���̫
Tg�7ח��q�Z�ǝ����`Baf�`Be���=�o���:%����l�@��h��d��a�;�}�|���c����.D�s��l��T����7txY�pY=���8�K�dˆjz�}���/L����m�x��2:���̸w��}���y����j<���'ܳ�a�<ۦ�0zق��B׻�TX�S��X�▾0[JVO�)~gg��}�D�=�a�n����hȭІ˪7���R
��j�wr�p�V���⌖I��8g�gM-E4��@�	����3�.����TQ:�1�������֨Un���q~�مB%ό���\�P�fޗ��?0fS���ҟP�m�=ΣL�k�Cs���uc��<��X���rk����6�sh��_�rnle�[���,Ѱ6��!��W��2O@	|h����������ϯ@�R_��U'J:��w2���Wi�v���mmd���"?�,+=��`�Ŝ�L_p~�Ɉ���f��7��3q��l�gt4hÃ�^���x�g���V�R!��վ�{ݟ�c)vp�����뽬�B�C|�`��>�Q�\��H��tˣi)�A=��ŋv��F�Sd���s��wCo_pM��omd�+���������5�bPmqƜ�[�]��߿�O�
L�0���(̩0$��뮯��\�k������ߺ���r �~iH�(@t��1�W��M��H��S�f���L>�d�}�Q~_{�L�{����o��O��y{ڽyt�YC��1�"Fo�dџ�� 2!R�Y]hr���~��B�z�EV3Wk�����ʦ�e>�2�}ZD���!6���5���[r���N��7��.������ql�45W�6��k0|����Ũ�2ĕe�=�#A�}�/	ڹz�[>��czk,�7�5ě>J�D������TG^��N��c�f[[�� ��ȼ�����'3*g(mIec
���;���ƚ�u-z��ֶ�qI�xmh��tN�ZF+��2�3�6�&i��[-g!��,���.�#�&ڸ	���[=/rD��!}�믷�y�3��:3���R}k	G7QR����f<�p3�bD�'��RL�ԧ6���w��uݚc�xe�����v�Q*�=�Ds.�bF��Qm�E�� ���y�U5�x$���]y��'�O����Hw>�A���}��CHS1J�[N×�&�ۜ�׎ƽ�i�q��\�2�!y=t�4`ҫ�
'��ԏsx�������_�Z�1��h���t��T�?A�)�.n�]+2L��ȼ��g`�Ү�x�d��Q�p�D�V9�N.�pS�}]x�o!9�]�[�b[եNu��������0$�+0�+0��SϽ&+C1���(4y�H�G���^y�P��֟z3���u+�ͨ��T>�1\��S��a�Ν��r����P콕�p��B S6���/ͅ�>��������K�n���M���������>�v���d~9@���o���x�1�yB�������'��+9ͽ]H6�ke���t��l����]ݬ��6@e���6_Z'���m�zG �0�ٱ+�~�4���0%6]��܏��Ã-�X9��K�����~I���MAi&-�^O����wi�R�ܡ��f�JƠ�n]<r��!Ϛ��1�ݿ�Ӳ�h���f�	�� ��*��ڰUG�EE0�DǘH��b�\�ͯ���ܬ�S*�;[��;`�Zv�Eσ�ֻI�U�W���v�6��o�ݰ���m�Ǚ�GN�h��=��!��������ne�#�)l[�6pڡ���1���%8M��G6��Z��gqy��g���v��DƱ�9����Sv��z�T�CM�;.��������sj�yLV��}����$2��Kz�@:wUY�?9lgv�� �S��<�	i��m��/ZB����:�Ŝի��F_7;7SS��cp=�ǯxn��S[��z��:��O[����]���[�QS�_=]�9��Ƶ`����=��}U�`Y��R`f@��� �Ǹʅ|�4���s�8��T��	��"�mV0֠�K��&�3uz�3�XԺ"�����y����h^v�ӵ�!q��,ȟ;���s6���P��V��R5�ԎP�9"ٸl�[M��|�gWh�6JH4G�r���gjgd�]��7�D���K?��>�Sͧ���e;�u]*����!zS��1fj�GP��������K���}]?���sqz����UȌ�}�`g�����?����k�H�����������ywߊ�O͠; +Х�4f���Na1�ݺ��/#)��͏V�g�˵3�Ƈl}��K3@m���sP�Q�0)̘����mt�&���'
�8�K�[W�Α�i��+��D-"q���1��?~?���!�A�]��!�Pk.��>~�#[GF��Nz�I�O0�9n(9�/�\�G��X22��K$��/I|A��;3Å��D[J�z��}���]
�촓CC�SK��������zj�Y��XV��~Q,�Ɩ~��=0��ߖ�p[Bu������5��1cc�eX��ծ~�X��S�+t0�缱��g*�2�f]�-8����"���j����2�JJ4e�5���`�UO��R��} `�c\�lJ��\Nk޷�>]�N"^�u�LO%o�8
3j��<qΚ���Dl��u���6��������޼��k�aI��I��[�����{��'�I�^�T��WA�ݲ���㿞���*=z��fZn퍎y���ޯ\9�n5e��������{N���o�B�Ϭw�)����/ca@�"�"���K�>ݶ-	��V֥��VG0T��oW���=Z�Jm��P��8�Ye����m�3�\�3�~�X�E��95���5�Op�k�kj������x��co�N닿bچy�a�U&�c�f��<d��bj����;N��R�b�P��;�R}ħȜT�X��^
�7p�V��r����i�e��ơYu�F��f�Qr����˟�
Ȩz�b�WJ���ܕ���=�>�6(����S<�[��b���Pta0wnہz�Ƨ����q��wa[iuJ{�e��-���q�R��:��!�H���ީp�y�y/�Ǣa��3MT� ��G�yo��q�Z��,�9�a"�Nk�QD�&�4���	S��=:�j�ݣ�z��VU
�s&\P9�A1������d�Vt3?l���7�{r�8�0�����Pތ�.�*o$ԇ�b[ݮ�YsLE�*r�e�kt�I�����^��v�Zk�	1���?e��e��ŗz8B������ ��[±���g:6�uI��.L�%����c&����j����&nn�~��2	0R��̌�_����c��C��_�uݲC<��D�6$	�O�}�'�>��G�U<�޽�U��%&21l��C�F��r��0�m�خ����F��g�<
h~�����}n:��)VU�y��j��/k.��5N�g��O9�ür���ýG}����9D��1�<�?��}aY���f�,����!�^A��$�A �I$�P�Onf~��T]�1�ug��Xsr���ϯ�"=��tkZj����� �����ٓܕLA�y ��0s�2��ƾ�M��H��M�l1L��t����KD؎a�P,�S������"�U��Ңj-�!w!�<7!1��Q^A���H�QN���];	f��Ķ)��u&F�-c�U���M��Tf�	q�T��eL���%4?���^J�|ׯ��4�]r��5��sg��.�ҡ�٘jb��M�iF.ȟF���T�o���1,��.��̥:r����qǷ�{�h�cpf#>������2lK�&
��HR�1�ŧ	�dÞ	�t�e�Õ>��T�3S�����#sV5���(�	=�@�g��8}5"� &Z�1�4[>�� ~�Y�=�s�^Hத���I��ௗl`�NdmM�Zz��|�����y�=6�JT���}c�i��R9*�B���5'���ų��P�fG�;��7�5��і3�i�d�9�3����&�i`��!9U�3�9�_�?L2)2�L�(��Js}�J��U���Ir�8Ԧ�>I�UO��y`�> ��{�!���a�8j�/qw9W�ì�-�Y����5?8���������%�EJ��*��=մ� ��H�y���YcB��ئ����lW�<W���gz}��(E�������<��T?~��<k˒Xx�m!��O����\�W���[{*@�ٳ"ZF�.�k�j�J9�ld(
&U�6?>������+z�!�@f�/CC��1d};ɗ�C��(�����Z���EfᙕTN�t�/;ZJi�a�}ȃ��WM��L]��S�u��B.8^��<���5�c-H��J��T�vmv՞����}x�o0wW��)������5�t���h��O>P,��1�����s���͕|����]�ܹ���k��7�7�U�t���>^���dW��;t'!�i^�n��N���;�����\^}�|��'�;���c8-���7?N[���C�KOw]L>�v��0�l���3���K ����1|�ʠ��S�'A�}�Y�4�m!�#�xz��������鬚G����fd���#�0��ʯ��n�⭷}�-<&#q�N�l��ݘ����2:�;�Ϧڈ�4/'g.3�/�n�_g@�:��,��zf�aI������v�Ē���;.�@�U�8�X��Ġ01B�|��gFgW��:]�����Ѩ��x6,؆���U�!��u��&��z�)�c'�ۼT+ax�KC �-�Y���U ��-���ʹ���q����X��t��K77Ce=X�a�҈_)i�Ș�`@a�X���8e�N3i��]����Wd	S.޷٫���B��(/e�q�^ѱ{�59�\���+��b�Ӡ�
6��8y�s�|k!1�_l�����
���CKM���'i۷� �\k���¸�3x.{��]�ح'G*�zZV�&���/S�f�]S\73xи٘Ik�P՛����.����X�޴b�CT2G���k]e�����wt�P��:���͉�$0���rX�t�'-�:���)֋8�vo=��kc�q�;�%n_dQ��0aʍ�̇z�X�,u��R��t��%�V��st��6�Q6KPj!>v'1�9w��h���(�ST�����,{l��X�f�����|r��.��[�]�<:���fF�r�c�n��l-J��oY��BvW7�[-�9�f�}��+=3�sn�>��l1�f��,R�e� �"HLD(�uM�h��6��`�_8��B8�-C��~8n
TA`?YD�S{_ LH~�|;iγ��
��/&�,mR�;��7DF�^�}��n0;8}ktD�=v��գgV.ɱe'8G���4���88*IC���@p��]��u��LTp�˾y̧1&�A̮�&\MЀĮ�&�<:fX����%uC\�c�N��vf}�r>]b+6�]lA;m%�d�1+��oV�y{�k�f��p�*=�wb|#V�e�S����3]�9����h�S��#�w�38S	�N�,�r���M勉G�v7�5�:��-L��k*E��nc���17	l+E�<��WM�ڌW�<j�1AZ����m��ݪ6^����]�\1�=qo%�1<�p
���}Gi�W�u�u"rպlj٘���JlŪ��Y���W|�oI��`qL�{���V3w�r��W��K�s�|�ׅVu�|�6P��oS�yh�
N��gYop�֫r��yLv�jm�)���D�"�ہh�,���42�-v>�b�����0,����B�"�Q\;q�2��x��6DY�S7j,Y��ktf*
�4kj�Lq��b�i�8��nL
���w	�Xv���@�nG�"D�_c�O��n\_w fܓ���Ԇou��s�wv�''3���ܿ�j"�c���Q[b�5�1�p�Tf��^Zy{<��k��է�;YuY����{{���.�.%��ӪMZն����m�Y�4�F�ܫ�1m���5AS����O������O��Vߗ**"��h'`�F�EEZ��A�|���6ձ�"��G"����9�3������(;�[�71��ٶ'j4STUZ>nr*���[i����o���������l֗s�E�n�E3���SG,F�����cd�������z���j֯��tp�9�	������=F���I���l��~=���Gq��k��1��UQ�W1�lEu*nk8�I�F���N�9Ƿ�Ƿ��U�a�I�9ȶƓ}�͢����n�r�1rMD\�V1���g?^��׷���j��j��s�9gl�g�ːQ��Ѡ�nG*����WaIa`�~���6H	?�ngMA'!�"H$��h*-:��ڜ����[��ضe�����O,��Ѻ��b3����}�ӯ�z���;�|��د�O�#03#2�)0�����~|��ʪ��G�N��15@��1��y8��]�� 7B��P̠��L^���d��'��ˬB!vl�5�M�o5SR�Yn跈�zw��!�9R*����SKϖ\�N�㡬��a���o&6��6�������1n�s-�\�º���aK�C���cr��q)�j5��ڛ����9�o=zE �m�q��>'����m��n�g�k;G�\;.������jˆYO0f�_70�����������5s�,�s�����ܬb��^еV�Z���}<�r�ȅ7���:��
�U�G������=}!�2��f�8�S������An�r�ė�g}oK���я[�:���d�yM��E(%�K�Ŧ�Z���_*���-0�1r��
',-ssw��ܱ�_�,PlqJ-JXB/��B���O?���Cmll��`�a-1�p��u�6�IId�����Ccݡ�@u�aF�Л�E�|���:�D��^�
�n�}u=�j�s�vy�:͏V�g��6W��ْ"t |���/�߷�������c�˲R}�'��4�����\�vCk�ǅ�,��T�aeL1 ����i�-�7�%�ܑ=ޥ�T�k��]�
L�\��P#�>�ȧq���V�c��^������u�Y�=�V���uUݼ��������&I��O>�������~�~��\������,.�)��H�C�^Y�#jMc�W��� 3�u�~��{o{���X��&�{��S� �C�6��&qP֑��lX&6ܗ�f�3e���Sc^����fwg��7���S-��\���?+�/���6z_����6�<�߼���oHb���I��]����:+Q-�&4���O�?���c�?��Te��@?��rc�5�Ww�S�Ѧls/l˺����wY���:�W�#�����U�F�pm9�\��D՛�*�jfG#�c/��q�� �\;f�Sn�!�q*a���`*�E����QR��{��̾��,؛z��(z�	��`%��kovJ�aMAnK��������5�E�7:*��f�Z�6�4��0�^[n�c�e�>ٹ9�-�vZmEH�l�^�B2N�����Bo@ʋgm,���_��V)�-[�hWD$�a),��b��s"����c�eQՓ}J;;%/�k���q/�O��(i3�A�Ǻ����s���d�ʺ^� ����Gڐ�C�Ū�FB'���c:�Lma�]��-gj���$�p�7w��� 3pHT+�{Ec�%qxT�»�����F,\�z[#��0�b��p����]&��Wu�wE�s�����Տ�vi��O�����}i0�A0�!30~��~�����T�?W��غJ�H�i��hF1(�|�	�����w�������D�+M~_��:�*0�����~�80EI�M�n^�����Ԗ%��&�\'�J��ᮦy��F�c���	�&�v�N�I��p��;j�~���k�J�ZW��v����(�֯��4�?�f�P_F=�����w}P�����b�zG�8Ȝ��f�^ljzJ;�e�%��S�ks3W_goD�q��{�Pmd��7��{�^��o<41�<ޟn���R3��<�^~�ё��#��~q�۹�ʥ��9��Ɩ�@����>��\�&���Z����gX���E�R��/�Un�h�` ̍�������Z3��3�����TcF.���Usk�d�q�}�-�x'����ّ�,\Գ��xx������S��S�N��M���A��u�0fS�=�e��~l�D�SO �*m�%Ο:a���'�q�*rƩwŝ{��5v��������yL~�b��w���H"������"6�!���G��ܥ��F�i���J��w�8p�V�[}�i��n.`�s�nWwq(?fEV�y`u����N�,N����d�di/��X�_F�[٩��OG]�>��bSx�{c���;�+��%b��E�=�Y�x)����j��/�Ɍ����������y������^*%2���ž�#%�\���F�ʖ�6hBl���}���Z����^Es�9�+�OuV��O��Ia����4��
!��w����/��*��;�F%�Xcݎ�9��u�P/3���y#G����j�i�i��=�	�� �<'�&��%v�����RUL��1M��q�O]2�za�(;�jEЈ	��~����Vn�!O6��O��5�5۞9�
�M݉U���n/mP�\cC�6���e���S��n-���Vڪ5��{���qO�x���R}k	G7�����t�d�L�u���E�{��� ��,��!�D����|Zx.2>���������΢	S��
#�u��Ǡ�i�>���p�9�oZ���į2�������r�7S-�,�)����������f+a�[D�V�{x����j��"`b�:|�h-v��yTS��QC��(����e�\�\���ޝC;VǞuyO��Wէ�h��p���³��o� Y�@������l/�z�B2Iړ�²������N����pͬ��ħ��Y,^�_�+Χ�{��<P��#�*k肾�>��>2�x�:�kO�e`�o�-���X��&������
/�`r�R�/E�3I�c�b=�]�������bi�����G�������_�P��{��s��=M��ɞ��t�;�pf�ff�e���0r+�P���]�{�C}:�s�}#:F�tmnw�䞑��7E��Pga#b���c�Y�AS}��x�.�	����ӭ
1l�k�ez7NP��<x�$My�RS��5.��.Dm<;!�	�mV�tw�fv�ε�z
L���\k+����v�Jq޽�k�q�a�g-�y�L�g�=��y���aq��@�J�g���,]�����19@��0;~��}(S�6�J·��{�9	ꓷ?/=κ̤D�L���rn� L[�H�{/P���B�2i�2���uk�e��o��.���ڦߟc�ss7��bK*��+h0�k�s�]�~v�`s���[P.�s��T��|Ԇ�����)��6@׎�oP�˞�����m�9�v<T�8�we��� �MC*.�>> �H�mӃ4m�,ke�Y.��} ٝaC5I�d�״�18�Z�V�����#�����;ȧ�c�o	�2��a�W�3��i4��ؾ���}��%:�`r1cʿ-�ߠ�@^U<�.`�Rbr�οݹ�;S�hT#�9�LX`�������ð�Y����̉2�Yɢb̄7k?
�꺰k�Ɏ���.���U�T퀅�Z_Psl�G&���cm�]V�q��;8�����̥p�������o���n|�w|����4���ķ���oi�z�՜�O�B}�W�_�$��r@��M5�}P�Tjw����}eB��H�k�����-��NX���� ��_����T"�{��垵[^l�5*�椭��&;�q�tܪt���d�F#���Ccݙ�3'�
7���t��B�>��ed�s�^�C�H��l������l��<��$���_PЎ-��#W�����;�n�qwr�|e.3TcIz�R7\���ݛ�1���;��C�� ���?<�,؟����w�z��g�`�-��o�z�������3C�q	7x�kC��6��갞�y;6t��W�bK�g��x�S�Rro*� i�m�sŗr5B�<�V�[O����{�Pe�z�7=3����?-����	�dG����U7j��5u?Uf�'��3��mz$F3H*�4�ZكSê��j���v�юS�E�PwP��q�q8=���j�~���Cn��VD�]K��4��٪-���q�kٌ|W�����?&��)oo1~Z.�iw-Tý���]\��3�ry�����H[Uy�"�MgOp�޲�zG�p��v���>�Eq�_w�f������#�ig�9�VV��5u>�g�h��I3�m�wg�z��\��{��~ؘ�!�"bg߇�̈́���h���~��5� e��P�	QS�� �_�q����O�Qf:ޯ �0��0�h%t+/Uk
e��P��ʖ���ӍJ�'�m�[��(kL����h��:��5�{v{;��d�ҧ1ž��Fh�w��S
:�VOb�	l; ��l�z�n>!��8�{���>��李����Q��xk�q>ᷞUSÎj�Mܷ�7쨇�|w��=���2��H!�Y���^x�K���<����W���c�ؔ�f��`ԁ��*^��m
��k�f�2��{h�+�qt3�c��A�d�	jd�/0��)�s�s�Ls;LdW= ��C�m�OX:��Z}���z�9�V��]cμ�="{z�8�L����k%�x�E��|j�9vxȀ�Ɯ�qCS��]�v�n��/���LF��DGs���
�Re�x��'I��_���B�Z�T�T�x�j35Z��0O�hD�t�����{�LRxheQ��������\P9�p������٫�;Z���^��^���!?�����(��F��G��xf���|ϡ��|�����׎T۴�aZ	���6j��+���;&��\��E�KS�3��]�9v��
�rY:T�"�{�1���o���c�3�m.���,۶�]�39w���E��8nf��;6�ʆ��77v�;�e�������ݝpXDo:�7{������|���y���=ı�h��7�5�%:ѯ^�PA��"=@s�'U/ށj�,�#�c	�����B,9~�F��>ª]�b��~�����œ�u�+:�-gg��^22"aq��ɥv#�X�c�]���.��1�>��A^{�
8A�e�fzY_��j�3�>�Mfo�m�+z�e�̤�/C՘^k���z�q��neld�(A�z��B�۸yG���Y.���c��oכ���9���ɥ��py�g�9��[��<0�"F���5J�o?��Rx��>r���#eid���}
>��� �k����k��P?�T��r��[�N�7��ݼ���Y�#~���ޑ��۬�U��!�����@M�Aɕ��1�v�k�rή��T�� :L�.r(�[��)�o��ȁW�����^�	���͋;=q*��]�ݓ�Xi^� ft�=s�tU)��%V�V�xŻ�aqm!��S���ܪ�����Н���h]�3;3؆�=!�B.%�N�����؟�J�o��\�3n���f�!Ë�Uӌ�A*��-��D�W6Y|ڠ�'�n�W3�,@d��q�N�Nk��Y��L�o��(��)�9�)������FQ�f ��vv�/:�NT:���13�k9[ru(���R�^��������$��'�έ�?=�������������X��������
5����(�5�W'� G2��6ުR�WF���Na��:��>;�t�u�K�0�	��
���P�Z�uC\���׻Z��Wt -5$T�l]�;�.b���B¤e^�J���z������j�k�L�jۢ=|j��ɥU�Э�oV��,��믑�sӃ�.#"H`�ށ@�z���챥�ӊ��`-���:��oķLB�JD�iC��W�c���,��O��={J����P�ƻK)<L��>a8X�y��g�P��� /H����|0��14�p����{(�W�a�;�B�Qm���{�X{Xrߝ���Y�i���)��\o�c�e�W�M��g�H�`��c�9�ͷ�r�xԪ����8|,�?W�еqŇ\�QAߦϹ��#�s��_�B�-���M��Ҕu�aL�V��K��vmS�:���"��Q�>�a��ݮ��D�e��4&�x騭�M�����k�1-��)�;M�T��W���?*��F�㧫5{���'Ӊ����f_b|o��*u�Z�$Y��ɑ�Kh����8�<E�2���B�V,�gy��԰���j�4���]�WHu���I���uTiSPt�<�E�sU�S�V�辸:-3K7M�:��;T�K��Z�}F�v]���U*9ο�W�뙘�&f&I�y������U���~��Tz����ĲmIeSj�Bɷxi�x�66cU���D�:�oM��t���T8�ql��y�[�t&\���Ӝ��R�Oz�ghp��Qnd�NVGw�����F�%��ץ.G�������<a#w?�?J���BbP��*��t�`tŃ�Һj���}Z�.�Pkl�[�i���O�.9��s�jؔss�F'��>V6���б�b���=���2r�rǲvS"�/��.~�W�x0L�2���i�R*���_;�������^@�u)�ܺ:Z���+��^�cXu�:��"�.���<��4q��}�چ�<v�T_��jH�d��"e��1���3'�
7�}^�;C���EҦ�Ր�]
~h��U{��a�v@���g�^��/��_A�[xN{�7?]+���f���Yh0h��>�TW�輁���炜ey.���Oz����֒b���U�G�v\�}ʾ�P����@g���K5C9�v�t����̌����#A0S�3�,7|0xQ��/*6��~��ɋeG��4>���b�f�d�A�:���3/����p�`Gw]S.�]s�'�2�m���6=�W��+b����x]sw�Lc��.r��i���F���˝P'����O`���G�9�ɮ	K���H�b�yNd-��1���ۯ�:�d]֝o�3�,^ü��ܳy�r��ݮ��Ϸ|������Ɵxњ+����V����Հ�]t��3�Ž����G]Àө�;K��z^]d�*^����6��Spyo,��%0��.R�\�y��C��+�s�l=����77�%e��;�m}�i�<P�1���Ȯ�C2�yD��V�i��i��o1G�ݷ�]K8�&��go�RF���1<����`�7x�[�ι��t���{ޭc�ާOʯVi��Fƣ�N������(��ᘷb�έ^��p���5�`��EQ�#-yֻ��%�&n��(t.�n�X%1ޡ�;mߤ�����{�X5�_�x�
��b0��-a(���*w���f�q��?B���o�8V��7E��f�Cu�5�,��aQڦF-�oIX�̚�`a}#[G	�v&�GP���Bۋ���-%J's{����Sf�l�y1��aJ�gK\�w#�D���j�s$I�Y#�qru���:2�^��j�n��]f�Yl���UBuu�"��,%4+w��.�:�C7����
��B������	m��2i,,��#�U���Z�]�+s��;�j�-_Ij�#� �S�!��j�����2n��7K}����.�&g0e�D��$uJ;]�+�*�r;��v#�o�rM�$���kG��E�4��}�.�e�[���Z���*�[b=ٶF�˂�(+�,U�L<�r��x�	�|ޡQn����sF�e�p�g���׊S�%��ޗJ�;�y���w��G�-�+k2�Mi���K��7�r̷�Q��4{�&�KBf��n���dY�H<ws�E�$��c�u�[S{�X�\cph�Q��U��\sv�����!�q�cI]��tbz��aW���an1KŇ5yg=�':�9İX�'s��bZVu�Δ��6�'9f[R����o*�]"ފ�Ӓ��o���=�j�ȪͰ���m���ӭ��d�q���x����vQ�8���&�R��r��C��Ѥ�POl�l�%Le��	�lJ�������v�b�\=L��_DDE�N����7��3׺�eo3H�r-�S�����e������Nk�ԝ��
�V�6��[�����Pm�ϝS���&������©�kf���C�0��t�$vy�6_J���;���#��ctu4��ӳ$�G���!7��ɫƟOjݻ��I�s�9�˞k&h�56>s�:&�ybڮ����(�j]��=?�����'z�F��xQ����q�o��ȸ�Eo�s���/y��F����*���p��]��\:6�Q1���������%�lQ5�ڍ�:�V�U�;j4�j7[�{|���{~�^ٻ��4��"�w6>c�r+i��Ƣ�E��5�1��E�8Y���X�ܚ�:�H��������������I[r�͹��s$�T��JpA���N�:_(_ �������\� ��5��~?_�m�!B�@��A�G�F#�4�H�*����y���1�An����1�g������;�	0��L ��,��� �SOv����2W7�i&��pMku��3����~=��*֩�j֢�m56�(�ڣZ�h��TE��rvɛV~���~��^�ۻQ0Qkkm�`���E[�]�p��j�[:�������5�m��\ڮZ�u��b4��u2l�77*���"���d�Z'C��$2H�(�6�A?�ԡPC$���@�$z��L0�
�$�ځZ�f����4��G9.-���iu���:�G��Yb*�	�4I\)�rs/zU�Y����L^d
C��P&�"��z�0�� �%��!����O�M�#0@��$�j�J�t����L�e�T(O��!4.U�,��$��"".U���s����LA=�=��mM���2:��cci�S��"2؟Y���e(�Z������_�r�Ȟ�`�?�F|��&��-�m֣��o[�<�?N�Ν
t?�^v��RoOc�w�C!���z�Ξ���ICm/X �?�H�v{�}k�X�s�3�~���v�2�tf���� �A񚊺>Fm�W�<ڢ}:��$FAN�^�T*�q��ek^d���qL��{�e����G(A��4������;H_�X�A��u������"�Z��˲-D^�`:^�7�BuO>��CޘM��D�S����[X��O՜=^��b����p������w��Q薪c=fT��Z�a1.}��I��-���B�D�M ��7z��r�qh��ax�{�d|��vQ����������AB��ݭ336鵯j[,�7W��y+�\٢?y��`le���>����?_�.A`3b����0m��V)�mC��Ӝ��<���2�)G��#�6�NdEs�����^�-xBh�ޖO-w[��B�V�u�9f�f�;�k�z9�<��qK�Y�H���� 8ꊶ�<�
�K�L���9�i�q�`���_$ ��b���8ju��
��.�3Y!ݳ��>�f��"���<u�Cw��eXD�8��ϔ#�h�Hu����]gJ�ss2f���nz����'�8V�	ˎ����K$����uٜ�ٺ�OS�O�$��8����ܝ������A"d��	��&�}��G�����{�Z��k���zӾ������U�,�%��9��	����g���ҩ�����)��vo-�|c��Đ`�W;��}����*�r�.+�6a= �w8�'���d�8�\�B�=��U���a��!C0fr`È}O>��S�<ޝ�U�����Q�K6���)�f.�t��N�|d�P�.$��&4�ށ@u�"|[dI��L~
�^�*?���+�=�N��ۺ� �kY1��&�I5��v��@f��!�^"F����{$m-"R�Y��p���:�HY��S��=�Y8M�jjY�u��D{1�iR|is/܄c��˪~$;��>Г�;c���h�d}��X�����E0�y�6Ο�޼��0�\6���������5E���@�{5�q=>�ێX��FPn�jFO�M���y�ڛ�벥rf�3g�t����VF�6�*CDU����q�SQMҔ�	�a�+������Rn���w4���t��|��*%ꞝ�-Z��6����=4?�~?:���Ow��n8�.�0�󬉽s�no;+��.0H!�vVs�Or�@X�d�bv�h����?,�ݙ	�͢j�"����|R͆���'6��2��GwW3֦#p�)=P�u�/7�X"$fֺ�C޵��#h�������~'�@'��3y�,3��Jԛ��K&m������/�l̹�;ݼ��[H��/��g͗ܩѪ��b����%��QaqYe��z�����Iec
�Q�(^CדE;�5�w�7�R���d��y�;_:�CE�Ȑ4���^�;�L4��bp$���:u��7C�q:�Ic<�켚��I1���vK�B�s_t��\�G��^S�jQ��B�欋��	1��go��L�r�H�(��߿| 6o���
~���K�:��L���@8�;���W\��G6(;p��5��9�yoq�V��ţ��gƇ#������C��8��O��ԇe��C�~�z2>�ƻr��^B�1	섔&+aӍ��Y;m���� \d�J�v�y؝�Q����ِ�=�{�r�c{X�6�����|H���l̀��
<�΁��O�qI�_{����O{_>˖w*�]�p�� ��9�[J���HEoO�7p,q�����4�=��xt/��cf(�
^����K��d&��X�^��p��iΗ��+�8�ud���f�օeox_������6�����=U)�Ԯ.K���ϱ;w��0O�X��;�ɣ�k3�5��;�a�yռ�`Ȇp�(W��wDl�(���������=ȭ��:�������S4��4�x~��>�R�m����7ƥǱ����6ۗG,7�8SVs�Fى���& 5�tf�������� �l>U���l��V=�g���&��^��vm�~�H"]���������] ���w
���Wr�f&槺��5\�0�J��3�{e!�6����/2F�����z�UK�U�!�fLR��!��Φѐ�o.������nq+���b�m'��l��gr�w�%�|�>�����'�-�Z��d��w
�U�s5�D�F8��Xw�cu�O�f�_KW5�1wKt%��g]�b�xC��!avt���������o�A�v$f8���-��~�z1-�6�"�LX�3!������D���V`��wu�|�K\�i�p����F�ĳ�0[U�;�Ӷ��j��y�%�:7$�r�^�ܲ�.\z�����m�nbƞe#gp0��j6��&I.}�M&�n���.E�WY�y���3fb�[M�$y�b�8:�[�Өu5�z
Y[�Y��ȶ�]����6��I����o)�Y�x��\)&��^�]����F{&����S��b��y��=� �&�i��&w�G��λ��æV��)�%6ď�������+�I�P�9#�z�2��%�l���37a��w�y�'^��wO-���[�nִ���{���0����,�X��_���j;���Z��-I��]�V��kc����mz�M�;�����?aޫi#�j`E�͆�]5��-���\�s[��ds���;8k;U��6�c<0�1�$���JE�6��ծV%bۺu�jۿ���&z�g�	���N�������7���&�"�+1�}�s��q*e���Sr��d�̃��4��*��e{~O��:<�[m�k�ōg����v�代�~�g�r/�_7z���$2w����,f���k2f�e�0�ū;��z�d�d%_����.gdA���%]��J�&��*�}"Jn^�M�c	�ζȦ~��k���¥�Ϫ� &�X�`��r��ߩs-���*�i�>�W^��[��:�+�/cG%�����.�U�Z�U��E�v�f:6�:�>�u8�xk��okp�C�TO�N��n8���T�F��jɢJ����+ƞ=�S�ٌJ�7�7���67&��������?������y��EKE�����sH�c��f���C��7��pv��'�N5�2���Q��Wh�<������J9���7��py�Mnru���2��mS��rV풺}H��3v���N#���ȳ0�Z쾎�������+����H���^V�[�<�%�r�n�k���v`�f� ��1�g͵�#��w˘]�Y^�"�_&�g`��f0���Q)_���|W�0��(�v��}�۬]w��ɍf�nOE�����b�wm?�2����V"�5��骛�l��#;�v>mM�����4��Z���n:ޚKr1\\���n���Ii���*s^:�����>���/&�)g���֩�t��S����L
�#h���_.zszC/w&��9�a�H�������U����!��;�4$4b���@���G�l`F�c!��p����{�Yxm�%,&[KS�������e��������s&�謜�X�d��1EPH�ͩ~P:��̗�o�I�4FR�u ^�{�<�=Dv�a8�T�+�VX��sƹu�'	��n��X9V^*����&Py;���(���	�&Bd��{��=�w��Զ�f�"�[�zi��5���>g-�7�xX�T�I�M&Dqۼ��v����l!���pR��7}�L�zLW�!�EX}�ۥ8��׾��r{�B����_��}�N�r[�|$�=˛����N��"[���L��y+��-���*���K=��g�w���V�^»�ǽ�}��$�����z�~����[�uX��t�M�*�p�����늆�o6b^3)g<ds�9]]1��Wt%�B�1hv�%��x�g�~�GtN�E��ݽ7mʳ�����=�di&.΂`�7��mؗ��b���w{�1<�58R1��x�!;��(L��t�ӽM��Z�Ws&���lm�3��霼BM�����L���fk������#ry���Ŗ(αӂbE�&���N�ӧ��(q��c�]ɿ���N����"l���
���Bf��Pނ��Y�*
O���s��hx'CE��n��b�m>��j�ZrW":WQ�B�P"�=�;o�"���� 2�\+�=���6�И��$���bʜ�p���-j.��Q���a��P=V��0ӷ}Q1ݑ�K�Ҧm�٩�#_��xa�2�W;��!���(:�;��ԣ��#1�e�8e�q��Kx��53�=��-����q잗<�wE]0�t��v"�z��+ͼ��lvF{*��������&�����D�l	$�y�;q�<��u���z����vGt���eF�e�׭��;���ֆ��������nҜ�܍9���㥌�44��j��͚��sa���^Ϝc��8~�~ b�W���5��{�f̥�0��s�݆3��9�� U�@s;�'�ߓ��8���zz�6�uo�"�]-]QO�[8�g�,*����ff�~��`5mH��*���d�r���*�\ �a�QY�?/	����#L�KY��b�iu�]Fn�cS�wk����Q�	=�.4��Ou�8�[�m�*�Ҳ��6�݋=x�f�o�E/��W��}E����ݩm2c�Vn
��}ɦ|e�a��[N�n�kP���4�X1���F���Hl�詼&�#> �u�Ԝ��;��J��UMd��n��頾d�W
�@T���V{�k7��\,czq��'���ҋ��eo)�5��ݴ: Q��N�nN+sv���o����Y�K��ߍ��`d�!Q�+)g^����"�2@P��D�R�Eq�@�w�ئ�ࢯ�G:G��flPiܱ�w�6�Ic��I��8�d��̵�Wc�Bٻ���d�Ʀ��r�WM�r���+�껻?�-��:{WG���[��;��	���,㪴�:U;��^G�wn �͜���oX�ܐ
6�^��7,���E�yvn�T��������;��F�OH�5ZǣGJS�[���Z��3� v�{m���-3�N)��5<��gv)��<�<�v�otY��/��Gz��a5�����3��/!�fn�1^Z��f���wR��i,�by�9�t��b�?<���������en١3��aw
�|+��[��k\��z1���sv�v�	�|-��Iyk�GWP�h(���8�d�����Sb�h�7��#6�{�����r]ٹ�I�n X`�[H�N���]���g4P��
��eYg����gm�%d6<4��	���S�ͫ��YynW���"���7s��J���/�ӌ`b���蝝��u�kR9yXynvF;���jq��]�׏7r��"���WN��G?N<uLNL����7�f��u�v�;6&����3���Sy�$
� �2���3�4�xS��EDD¼�ս�:�Z�?���s�ӄ�{��C'yNP���~���w~�o�^�a�9�u�e�z�4ϭTn�;+��	�Q�f�����x�/��j�f2�4�s��[�ν����<�^EEE����^�#��`�j�OGz�:�+!ۻZA��n���e>�Ş���p�ܦ"����1�>�z��=S�'v�5��g`J�F��U��k|化����=�кo�IɃx'���gw�fk�ؚE���l#@��.�{����ڭv�������V��9���]�q��U��E����g%�'��:�w'܎*
y��,��Q�\O��]o���g|�r����{`�=vzxt�T
�)�vlj38�����ut|N3�q�� 2Θ}f�6����#�!�C�c�>�ɼ'���������Gۧ����K���2�2��S�µ��iB\�1��t�b��mc ���[-�2��L��}�����Oz$Q7Wь�ڷe'�r�L���)
%e��]��� 癗�`�#����:�!��-���6�}������t�)JQ;�38 �|7;��F���M���[wDb�;�A�:��eBl�ϳ77��-\��=֐�fM��/2S]!������������kB�V�[�|��c;2�-�H����d�WL��;/MA�q�6r�)c����L��wՙ�C7��8���TG)ګ;;m�щ�\�pu˩jر*�z�b����ͭو�R��ʷ (���ۏ�as)�|�[6\�՘�����J�6��J	��fN�엗�ʩ#��n �g-B*�in�m��L�;`��r����v�\]���u
�;c��Km��J"�֧NM��N��rH��|ka���m%���^�v�-78s|���yo`�q� ���̩��� ���n$��ʺ�FQ*H����������"��_����X����UXԦ�r<ϸ�Thh���s
�0���v�� 3Xײ�vuÃ���)�.GY�WO��zi��J�)�fL T�Q���ؤÔ�Ubg5cF���e	�=&�^H*��!C�S��ʦ��3��Hr�5��c��2S�i.<t�?3�����~&�2I)4!Nc�>	�P̄�P�9*ISm��_b
NK��B�I�� ۆB,�F:��H3�AA۪�r�r2��a�V��mL�P-��ӄbpʀ�Rs:��=Sj �`��N�xө�j�{�r�]:�4�o�W���)j��x�!�4����^�.Lؔ�l�޾���Н�/[i�f�ci�u���o�Y�Oe�ٝ�e+f+ƈ�����L�����
2dq��Oz��wa%+�p�p3����<r�,���t��kn������E�t��o�k��X����0�]K�z�-[�zT�݇�84F�9W�&�l�"D��<Mc�սsqwP��C�P��p:{+0�p��V�(��3[+�x/nd-a����Q�S�S��+rV��u��*��bԲ��u)������z��� �I��I�S3��.6
���Tm>ƺ�t����;\�iϮ#��`���LU5Jƞ9FnI�C݉�V�.b�اGmJ��Y�u���Th8�RCPu������&h.�"���2�	y��>=?-$l�ʕ��e�&9���6���A/|�g�gY���2f=��q��F�#K��Ss�wN�b���a�����M�@&U��.�[�Y�(ږ��Ҿ���@��(eN�Ц���1�R�g���+�<LE桽�]^܇��[ʲ�D�|{(k#��p!v�N��:{w{1&*(�!}�d5�l��J����D�TET�u��1������_����h��A0�wncE�O9�ڴF�S��cQ��U0F���3������w���p��p�AG�71����Cb����h�5u_����$���������4i�4�F��LG{3�Um�Eb�DEm�b��(����TT������ETPE3Q��TlAh�5�m�[j�gL�kT�9���~����x�Z�.skl�Zj�N*ӱf�*�b7{�-Q��������DDT�V�#PSE-TV�.r���(����mZbѩ�"'Z������IQ_1�QCMU\�Ɋ�i�l���h�c��L���m��j���p��Ƿ�����|Ή�
�j	��1q��뚞C�h�y9�(�"��V��E������h9uG-][��5T4^�qP�W�>G*I�<��/8�f�h�l���Wkx�� ��Ql���t�կ�����AJl�-v�s't�e=�,�ڷ�=a��}�u���fa�5�k���W�|����o�|����1��-.��Ѿ�>����
[����jj��[fEN�.����Gr�4}��Š6%0:��&�hjhw�k�ƾ�1���P-�y���	�.L���}4�]�i���l������݁�)?�J�ϗ8�rZ��� �j��elsMؖǺ��L�m=����hȆyH��>�s�+3���9:E��3��6�u��	�o*��\�YW����sT�&���k�c9 n[ηZ���ْ��y�	4���v[�<>0e0�H��W�4�q����l4�^S��r��nA�G��NPՌ��D\�w�T��J��\!��_!��miv��P�uh���T]^#kh�U��Am�Wy��(]ݑ�YqI�c���*�:ح�IRR��f0F�R�����u�ߑ�\��7�J:6dȜ�ką�-�dE��H ��ͮ�@�W��W%� �l�qp�kN��Ҧ�q�0:/s�ھ��a��~�A�>�7�Jol�zob0sV����;:|d]�iuqbg)��r�'\���Z�D���i�xΧ}T�<f������=���|N��C)O�FZ7@3�%R�iVH�y�-o�N#�f龭���ӵ�bh~+V�m��@c�>n�j���{/]�~�Hok����m��AI�#�5ו�I�:��"��p��9�+�w9��%�s��S<�A|���s���͜��;�C���W����󡏖�n9{�1�j�v���S�Lw�d�a�[й��Ua���͟l0t5����?��o���Y2K�X���,�pW	��yҤ��$Sw��-��Ձ��7ux�:e��ló3A��Sͫ5����O�������Dw4�e$ގ�x���9��1��� ٛ�k/_o��φI�9L�L��bb]��oI��x����b�{�3���G"��g��{1��7� ����ˋ�]����+��*��)�^0_=	C�r�f{�e������]���&�4�w�%��4�N��'B鎋7g2���<�\�nu��w�yF`�b=�;�G�f�U�޾mM�.���%$���k��:�$��{ѐ����0p��u������n���곫v�s��.��0�,������i�K�z���l�d��@0�?Q��P��)�Y������v��?d�l��+1G�0Q���v�ue����TL���Z_�U����'�qC$�X��G�/���S]��-�j��P|��/J�;���J��6abUAKj��NKv���K��i˼�qz��\�-����q��P�Q�vʭ.ٯ�b�B��+k�v��ۛÿbugv i�̂�,��{��ba>�0���9,pK���ᵂ�&�r��kQ�|:Ե� xo9d_���V�����m���>n��}�����2�o�l��~��}>�	l�r�-Så��ޱ�]5�m���6���6o{�-WϸQ��Am����[�/ּ�	���ou`��ݡ�tFDJf�y��������~�߷x���c2x��=TD^�C�@Tf.��`��"�AF:�a�ݔÖ��G��n���"���+�/��f7[..�����U�4HkOf���:b�vᚻ�ヺ�AV�㲸
O�+�`� ��P�e^�s�K���t���u݋O�a�Vm�:ӧyA���T�ݔ�_r����8�/o��ݭsջ��rɮ��7"���4�)�7"痼���U�%{�(h/l��K.�GNv��&<;e�{���=�˱k�Ɋ��δ�\�~��6��6|N���[0h���`�0�p�<xF_H�����qb�V;�̤4����"�Ggb�i��h���{���sa|�����@���~3q�t�M��6g��dx�f�6x�S-���Gmc]Fƫ]�X�&��&�U�춱HԍHd�S�5c4�=�9P��չ�����&e���+��׃��٩�ꚪT��
����x9�C���0z��_�'�r�+Ok<zv��i�ܹ��7j�
��c�uMD��4����t���ܯ/Lv�Y[��Y�>��Sxˤ5����mHc-U}v'1�w=�7ݛs�� s�AX���r�+�UV���E���E�&��[��zi21��*���=V���@����M\�tȄY�eL�@�f"�u���4�`Bq�z������X�R�DW����|�I���}�q;֯�:�ɋ(��VE+b�6�.�5���Z��%�lX��u�t��7�� R�w7���wN1���'>���h����!�9P=?n�+��ͯ����rWmU�]���zxm�U��wh��h�O���-5n��8��C5��2����4��bf���}�S��Րoַ	���$�fۤY�6�7Ql�v����Y�iq�Ѷق nΘ}�r��u Z3#�xlY���۹㩷o�������Y�8�؅7�G�|���ސS�
��0�\�y�+�����Bz�Sy����t>�->�#��u�TLBqh�>�N�pi�2r |����Q9D����zCl�m2n�`I�v�v.�1����;�qV �^�k��vwnh�c!��3BɁ;�Vsc^m��9^�e���4'!H�}����i������"F��G�FH�1s�$�mؘ�l�mV�H�T�&���SN^�
��¸���@w��^ҙ���ll��l\�]���a�ɜ���WO��[��Lb�bwwm��YxeT�E:���� �H�H(�� �I ����z_�=�o3��
t���;���H��;�}Ԩ�e��ƭ�P͎����tf�w��ޓ;4m�[h�b�t.=�L��L�o��h<m��jߺ.�����d�-��k�\��ѯ�f��o��kBק��j���Ǜ�K�֦R�Y�S�չ;Y�f������}��х�M��VeP[��]��k6<�掾�O�ي�y�ns\Oa�~;ЖP	E�@%��d�I]��5AT��-i�g8��:ۍ�|��3K��f�pz[���lrV
��iV��.�$`��U��/oz���i�r�E:,�pVEj��h��~᧥л���)�Y�F�K���uB/��=�e�6�Е�k]�j���;��hwu��wqW�m�ݐ����Xs�x��ȇޟD-�;5%��&"����֓�.�vj��A&�u�N�Rs��e�;-!yn�-΋����.���gws���S=O�u*�u#��������}�9�~^W'l��, ����u��>ݲy.gI���Fg���6���s٭��U +��J6���Ę(�7^��:�p�Z��o1He+{Z�Z�b�1�lHq�V˂��h{��q�I^먶*W+�����u~�Ĵ����H�o����"(J��`�1P%�D�!RD	>�b��������p�.y�w��=f����#^M�Ev�[�U�f�uVU��޷����L�Xd\z�ŧ�ӛ^�=}S�'��p/$��|<f�oj�)�9�χ�ۜ��n�FGk�S/p:e�SM��S;�xK��	���e����g�|��J+��ķ^�|����ƴ����,^�k�zC>�<P��$�f�i���e��<X9�*��5�:˻,��.c�O�R���_9!��^+e(�<����k��r.f����
��L,�*�EZk�oԯہ-��r��h�U6;_m�˾��~MؽOoY<��{<9�H�Kl�w�{s�M=�z��+k��Lf��g)��*�i�hc�����%_b�M��s"�#��n���h���^$ǀ�qf�� Q���s�8޵���[�!����Y���P3��ʕ�s2�-����`_$�@�mp}��yR9՛C��S��L^.ձ�y�ۄ,����Z[V���~��>�(��W��<��\��<o:��8�-t{J,���5ǂ�����@���vc:�S�24�ɩ̦5�������~5�U䶮F��V퀎����FҶ�Cc�\2�����i��Y��f:N�J� V�
�E�6V��AK�>��ۋ���Qj�Pd_��v�Y��|���}��+�vGF��J���p>yG�
�n�,��9,%=�M5�vp��f#��w)��DA�#uϙ��ڹ��u �����b��1_c�V���{>���M�<�/InFO8��3������:�].!-}~�a���a�g�Z[ �WMrK���`�����u6�V�o<433�f����v#^����d7O�0`>L�#/���P����5_P��j�JTy~-��׼hW���}��Y��,�����{�&�Vv#�Z��<�-��m��h�'���,1���Q�H�s����Nn%�����6Zc�[	Ț7W}���<����L�N_2}���rw2r�[_�S}�z޿x(��d��S��j���Y�w@t�3K�,q۝��!S��G{Q�W�pPh�u�]YĞ��e<w�c��|����T�#`=����qWˑ���G�+�t�t���Ϯ�3y�ܼ� &�Gr���Y��M�k�u���Lt��ǒW6�B�S4�[Ҙ���'����W��;�7qQ�g���Un]>xꐊ��|���� m�77���{bwv�A�k2|P���.��ex�tw�u�v�l��n�K���}Ĳv�����^�N���$oثd?�*��z���IӬt�����R�gz��Á/D���˼�����W�K�,�]yC�f<�K3�*�sӛ��ѝ����4<%���wo����9�y[Kw!Ջ07X��#&��#���3O^v��������>P�[���Fz�D����!��&�����:���^s�L��ڸ3�5�ǳ9�hr�Iش����o4E�O7��XGm�I%���{�LC={C��l�?�~_x7�"��~���=��e���
F�+�O*�����r�5���~��vZ��П���cf��2��kGӮ�������=P�o{t�b.Z��̰�V`��u��ձ��n�y�@��	�w�g^/o��sm���\K�d宫����t��{��0�,ᠫM�Cٽ�%䇐�����pp�v*Y����q�~\�1��O=�=�Ʒ�_N�;�O,�wz+7S��Ѱ��05{@�d�c�h��mN�����?Q�|B��f<ֿ'o7�-��bj&RI�}�^�u����Uy�~T�v%a��~��Ta���OSM��0��I�ݴ�Chk���� 
���Ö3��LobSF�3W�1=WcMEo,�D��H��L�z�N�y�׃�C!1\�7����j���'�b;�1��M�/��jK+o��e3ǶZ��ᙙ��.��kz�cqa,��ܟW�ȼ09�v ��vVٵ�J�v4�}�cm����)��ۭ��r6��%[r���#_���Km#K�sW��Z�ƭr�ܮٚ����os4U�����U 3٩���i�ѯ��.��&3���g�5V�s�Fp�gz����"�
h��Y"�E�4j]�
�����a���/��m7�F�'�غ�V $����`�4!5�A2E+�Y��=�`��3/�knT�_*Kem�9*z�S��Y�6�]IZ��e:x����v��%[�`{o�m�|�W�5+�3��d=E��Ǭ�(�MU�>2Ѡ�m:l�3�왚�A����R6��(�*�L2k��:U.mE���P�#c��|m��������W��s�,sw]`�r㥬���%/�J~�ך�����`�Z�+�YEo�%�|��,J��+3����ח 7RQ߷Y�8B*��D�3�^k9�`�d����Q�ΰ��v����J�Ň����a��+����Nc2�jY݋�;���l��,�}����T��	��ͺ���-��E�3���f�"���vwS����J>c���;I��>%ηr����SZm�'�"��o3��rͬ�T0hO���	 �@�w�M�.��uP��]bPΩz ���Y�"�6���l��]�����2����2���UMSV�����z�9�ƩH�#��eh�ᗛO6}|��Q��V���9S8R�;����u�&���ދF�ge̺5�ݭ-�0����._wK�XJ�W��e�T�]�G
�9ٶ�B*V�v�p@�W�^N��bC�C\���Y��&ֳgӃ옛�Ǜ�uAy�K��n��03r�+��0���(D��#�e���E�(&�#,��.�
wj���tp���s��Ƥ���v�둾����5�(�-�hb��G�S�+	F+q�o7��۶���{�ʁX�i�j���4$��S�P�OoeE�V�*'N�$h��b���|
��6�k�EU�zܙ.�'���؋���5K0©u�I�u���f�փ݆�%���@����������T�v�Ӷ�h9�
|{�#�n��D����U�+a�ym��1�.���%��:C�f�o0��/�z��nc�0Ψd��+�]'b�V]��Sn�a]�%l)�ǧL/���tg�L��wJOek*:�4J�p�F�̡�5zȝ�v�(�Ri�i�JK�ə�����n�6z���� ����j�7"����ȃ�:]�KK/���au��Z0�J�x+gc{NPǃ��z��: �����fK�t��<b�t�H�=C�f��$����	��g��J��}ˍ<�f�`��p�N�Z��a�|sBS��+�\���ީ�)S�����	j�D��W����rT����q}1A�Ke����m�;��9n�ޚ�/.U�9���&���:��mj�D�����Uk-]��6��KjV����nR�����*�]�����f�f�����j�7��y����8�=�����K;D��I���\zI�i(
iъkE��4�G��u:���`�|��TUU�\��zO�oǵ���31G�t��Ȋ�gwj�b�cQ3l���F�j�RM���3������5CM]�6�E�ES��F�r�¿6�:�8[ەsj�$��)�*������{Z"Z �ţr��UUQ�trm��cZ.X���F�g�oooǴ��*"�
:�]�-����ų���h��9�E[h�U���֦�(��Ƿ����;��F�ӈ��P��JBL��g��H(@��3WS�ʊ���Z۬q�����{�DQ��b��j��D�V�Q���s�*�a��ˇ��خ�s�+���������{	&���i(��j"�"��/��+���G��&*;؏��F�Q���TW/C��������+m��9���th�W.b����g�G%�E�ǷDLu����N�-��5�u��%�a��z�w<�L4���<5b�J*�kd��fncQT}�	�׾5��p�˛�96�"��Q�f�H7����Lٻ�e ��G"h�E'ò���5��9� ��2�ݲ޺�={l�wnl���;�f�8��3�QHi�j^����~
@CbO�n3�F�`��_&��Ip@[�2� ��ɍYh$)�a��%�
)#�@�-�I��!�U")�]=+j�Y'lI� I�4���q�S&�<WG�M�{�JY��z��Fn�8lN����{���"[s��H"x��\�̰��2|J��y�>�2�0��o��`1w���#�ݧ�"cb�=2����*�]�,���M�!�L�/���q��L��Vx�����-�;=Y�|��:T�RZH�Щ�"�<Xv�o=�C��H�Y�\�Ö5��OQ���p�z{tg��4l\M�u�n0>�-�T{�фϠ,3�vcֲ7#N����ngp�G����$�v�fyX��-r'�@���)�8u\���`�>����s»�]��,����%���Te�������'�ߚ�af@=��b�w��S��!�3�oo���d s�9!��^��F�H1@x�����n��7u��WfI���蛠(�b���bCi=�V�<^�����T0���,퍜+����}]hWp��x��^Q���|E�X�rE+�������N��-�*�;g�Y]�6���kq��\2U>�H���{{7�\5g+8h<�34#`���r�4|�{���r��QǻՓoW�j�����z=Ė�k��6��)����	LK�l[!+�\�������"s�o�����޲��=��v��L�MR��o[*�H��I禫�3�a�;�vgpݩ^�䦴
G2�9X��� :f����^�<_]��z��a�n�F�kO�����q�Vk$
6��9��o�\�K����VwMg���m
���2H�c+
Y�W^P��u^ޏ\H{b[,sb&�Զ������"�����\c6V�����:j5�1�y�V=�k�E�H'nC�5ׯ3�`ω�	���_��ѯ'\��IE��G\�V�v��lm*��;��Y��/��(e�l�-�w��b�8�|F}:�fdn�;`�:d�ª�;=��Wې�2U��z�y�������vу�%��Y=�S�q�/�ֻw`u6����V��}�I�����p�`T8�zk���\Χ�~]�����̧�k4:�K:�e���L[�����o������7�C��|&:���x\�i�GW��Do�k�]W�7�Ǔ���CM*-t��H!�7�Ժ	� ��[��y�z���]9˞74���N/s���3�k�v��)���ot�x�;ѯ��9{V�����ӛ̆2�p�����~B��0�w+�,`M�{���
��F�͡ϸXа���N�(m's��En�G��}['�4g���8�߭�����#x�P��x,.%��xV�V�ɾsY��M�Ϩ5�=�"&���[��8�0a��q9LF͙=Y���	mΗ�z�g�q2��f�.��j\�*��ԁ13���˧���fd�����˲{�n�Ê�n3Ǻ[`^�:ߦ�%���QmQ��7��u�����.�-;	G��6Oߛ����ګK*�e`��Y���g���ܻiҫ���vmi����	e�)x��zn��y�i%�OY�-9n��95Q4p��G�(˞�"�\�Gsͱʀ=+vɡ�֎W�n�r�Zbq�u�7;N^h���	n�p]j薏g%=�x�/+Lk2��8�~��1���C�V���o]���^%��YZ=��M��o8L�5�=�{�-Sǀ>~9νw�z��MP�}�]��_:ǿ<����u��B+��}z�Oe�I�
5u7(�㱪rGۋ���,_N	�x�|~���{�7_y�z�U�wT:GG�g$�G3�#Vu{ ��{0��pև����!��e� �$4�)�wW���`o@u��/��r��y���2�Z���3|��v�UŃ�Ja'��4�;���	�Ya#��p�l����9m)&�3�gL������T�Y@%�s�m1���ʹ#�����j���6��N��&"�f�QΙa�?����C��1�'���d2�!v}nc�:s[�-�o�M֜[�]o�@6g�b�f�ڽ�ݜ��m(�o��-�7{g�s;K��̯�ā+L��T=�r������³�s=�dwuw^���6|tX��i��(�x����0��W��տEd��z��`��k]=���ݺ�l�����3�V6[>�R���P�l��I��/��ʧgnr �}�V�W9^Սn�D��\D���kޖX�>FkIٖG�w���v�q�9��H���ݭ^ֵ�G��Sz��o�;.r�ɮݛ�v��3xi�ݸ�����B	
LX����@�8����n�^TY;�/9��uY��R�Q�g�MLR�bRwS�z�Ɂ�'��ؑ�(�]�r���S��w��v�#�(�h1���no�Y&���A��|�m�B�8!��3;;�RgO@�Ƅ�q Q��	8�]ºg�ffYn��3�7v��kz�𑷾!�Ǚ^Hrm��vh&c��֧5�a5v�Sq��H��k��l��k�Z[>�K�����k���m\�mp���;��N������y�)����M�,�Z��b�5ST�J�;����-��@7I�a.�,�x=[#��e�ޯ6�[k�FdS���{�W��N�0��r�U�c^��%Wh#�6�Xf�yٵaً��,�ws�B"�*ck��W&Ƭ�(��K�b|�"�f��1g8�j�~��=�|֍���&u���R��}ҬM$�;�e�s�!J�mvh�X,�
�	2|7춿h�����:��l7���	�UW�C��v)���׌�z|9�w��A��FB��n����/-������'��'z;.�
��lWZ��HSiG,Sl��+PFPX�G���N��z��9�2��y��|��ة1�f�+Y�a�R	�+��L'�<�¶w%a�yl�J���e
�K�8v����^wg�>�{���=�����!�t��dl6 d=y�<ə_Tb+Z��׌��Ox;�w��ۏd��P],�0G��,e��6)��C_;Ɖx�)�?e�n}�=��<Ve�&�]��-���-*٨����̈�3_�����wV����o]zU)���T�N8���!��:F+eq<îpF�^�N{�;���$E���F�
��y�'�.U>dq��i[���Sr�7ٿxM��j{�c۹�$���g�je���!��x��*Zs��q��ʧ���ڝ�w�Hff�̊�/TV�+2��xl�X�j�9M\.��x��=n&x:�{=O��5 szX�X���Y��6����'v��}�P��2F"��n�k_����V���#a����%ҍc����;3�4����q�F�y�N\ƍSpb﹦�F���d�����(ۅ��ݢ�fp�Ŝ=���e��p�:,*�P�ʇ�0AX�n��N)��E�K2�U�&S�&#��E!-:���2����X�����ɾ����]szd���:��첪oL�
 ܷ*�8�����Y|�c������t�(gK���S����xu�l��h�2 >�O�>��<��d�ڋ��wM����bn0�ɼc,T;�r�¦���D�0`p���`�LA��X��Z��Z=
ڶ�3�+�������ʏjEe�S35 ��WQn��e�"鬔2�4<z��	��q�d���=�l�W��>��&[��q�8��0�8�!/�1�\��D�3�x�>ժ�ܰ�M�i��2�n�f6���Rm���<^�k���B�"{��F ���sk�}��͈�@���_<�g�1j�n�m��1�~�~��T0c��q�ݕ�Dl�q&\�v�����x�ݳ�gm{��U�� ?%�c4�rz���ز��%�\�׍*�9��W]���`a<�+��M�S.�YR_��U���)���~�o=x�_����(�v���$
�	��qG���g��s*��~��`�ȼ�3�`6������~h�H���u-gO͓�WZ��Y����ع\�򶢷 �U�����$�]�3����b���f1X�ݒ���r���9�Vx���E&(�VJ���gs0�s�U}S��N�\y����-�vWW�fU6�hL/t��;n�)�Q/�c�oZՙ�i{4<�o�s�n�XJ]�l���5Nب�H���YҾ�D Ag������=�Ϭ�Šb�6�.��iwX	"L�ַ4g�ro/3FUݨ�t2��q�ළ����g���!\�JO3�9���{{z���i e4>�3uu��� ϩuo7/���|<��e������s߽������q�/�Ǖ�J-��VO�@���t�} w+��r^�-;���B�P�t�:�wm_�1�V����!��������Y)d~۞�x�ww%�n���|�n��ہ#������9���ol$��v,s�F^���ţXf�:ԋ��j���߽���8vY�U}=���+�OeXi�׈8�da���@V@�X��k#|�y@k�pR�뛢��<�/�`{8�+T���b�^霕�K��ܙ(<��zt���z�:7��y�B��ը��$�I$�wϞmn�V��O��YK�CD>S��+�m���fJ9����Y�"��%jVyh#k�b�cT�R�8�]߫��*�(v�N�ݘ/��{�l%M�D�)0[4!m0��%�&
}����X;��c��^=/�0����f6��7�5�!�0�N��3V|�wƓO��S�� 5z.Z��?��MZ�R)ߡ�9n�<��=��8��8�����K+-��(2��!�"p��(������������Nn��,^U#��xR�w���d̺q��3�����K��ڢh5}`��'�q>�(����Y��M��{����|Oٔ��u[9 ���[%W�a�~<:��R��;��L�}\r��N�^Ti�^�&��l�X�e���52����&��;��o/ɶ��wv�����s�{
�N7�W=���L5?����� ����CL!ڞ߶�Y�h�/5y�ӡ��Y�w8��^��k1!��M��A�`�i��d�~���<�g����fp4�;��^����8).xb���r�8��.t��B���:7��/:B{���|���_���rPށ�A�5�f۱�:�W��������)�w�bWm�S�#AܤqV�2\7ϻ��p0��|�h=��=N5����]a�>�.��y9xe�`a����wj (�ޡ1�(�c���N�-Ӗ=!p���0t=A���8�m���L����؋J�ζtn�Wݬ�ƕG>�͸���5�����8K?���ڪ�Ƅ�y�n��09#_yh9СNq֮�����#uZ	c��_�Hn� 0$j7Lǂ�v�<���ٻ��Wlum��Kr�φG-�mt�2 l6��s��i��0R9��j�g�<N5Ks�+_��$`���e�ذ�?��~��D�(l�?v��H�B�m=�x��hv���-�/x+�L���(t�el*�/ٝ���rEY 7O��"n��`�L���f�ޜ����c抻���!�q��6ϐ�͞�bjC��Ɯ/����8�%rD�MVl�^m�ӽܺ�$w�VCIM���ǘ�3�K(�)���#��l
��0�y-<1����f���-
'6��"�ݿbγj�Eγ�V!�i��U3�2���3�2�
��+c�L�
?@��|��l���uY啦XiL*Yg�;)7�l�
h[�x���j���c����sz��3D�T���:c�הmW��I�+�9㚻a����j0>�/�H^�(���!��6Wf�K��oUt3܆d�rl�x�4��)��������>��{�c�Z�r��%�\�殍��t�^;=*���I�Q�j��/��1�=��E˭� �G���jN�}s7O���t��wZ>�ul;�6�n��4��u<��S�z��ػ��퀆ʒe����Yy^����ǉ��N��Gxd�R�g�M��asSr�pǞј&�/�O�L�,L�����X���k���
�����ө����o����a�s��q�S��=x�lV�	2��ײ�Ѷ�WQj���9�A��T���=r�6&��bX!e���c��=d���I�X�u\U�¶�;�pN�	����i���ʲ-nc���˫6�Wiآ+���pj��qk�vۣ��7l�$2\嵦�!"�'ٖ�B��Ƈ]\"���.�E�����.JY�.�G�:�XYQ����u�� �ca���\�lS�{�3�т�����$es�(«��tm���� ��Z|}?H|��) �h"$S�K�N �ݸ)\��Yh�C����};�����nw	]���x��5�Q3ُ)K���l�7���}��依r�%ڱ�O��3a�S5i��u����P�6�D�ه�q�%M�B�[��CB2��W�T0v�r��V�sf���#[�lZ���̷�2.#R��j5�/B}��HD8{x;�	���K;�:E����&8�Ȇ݂C����u]����O�3���\np]2Py���W��z�Зm���K:p�8mdW���bF]�_^��i!h�3{��q�N啶;#�]a��(%X[��B&^] v��yeܽ;Ǆ�w�a깻�jdr 9o��/�ģ٭�΅�7(�.wh��҂���e>����=�!��9z��c��tq�2hĺ��RR�>ÝXk��h��g�(z�DL�I��}�⦾}X�&L�p�m�}ɨ��:�R��}�7ţwwS�T����F-����JQ�u�4��_=��6�ՍJlulcyT�cK���2�@$��u4>�u�߬.T�\�в�7@WJF��*\	.Y�s��04���b��W:�/2���fZ&2!�a�[Nw��5�2.�N��J���K:���\8�-�Cy�7=����3�;{�m!�Bd5J1DHc���\�2n��9b����M�l��Z�c�6�=>������*fd��Q�i�"
��F
*96�UU5s�5lW�gh�q����V�.l?_�oomET_-QUl�;���("�: �F.Y�li��#�cF�b ����ק��F�}�Ir+r�Y�j71Ö*��r'#\���I[Ί�Z5�1����~���]�w+�s�o���p�����Z ѫY��g5�h�*��:�1��ܧ�������7�=c�11WW8m�]�k�)ֵ�*��c@�l�	���&�G�R@�Z�����~?٦�Ƣ����W޷��TVɈ&��ˑ�:7޷Fh�X�}�t�o���x������m�Ʀ��Es;�5Q��/9γy�/{y�K�%`"��|c"Q ��I}�
h+�����=��5EAsk�:؎�51S[�F�}�ߝt�9r�����M��θ�s�K���9��QN�:c�ܣd���1�N+���1m�����1U�±�X����k�G\�J},���1W�}����ʥ��H뛏{jp���j���]ťVۣ��E�T����5}֢8�����w�;46<�FUnwR�����<�L��mfwZ�Z:ge��l�@b�j��m�ܭMyy{�r:�D����	e�aN7�Y>�kh#��������:`L,�q���{d|3�,��LKn�6�V�%u�GZ�8KQ.����ͭ����Ȟ�%�Ղ�@���aos��ܙM�iqb��UU�6�.!�48g�J�h~�?�B^��K�9'=q��Jdm�D��L�
Y�5H�C��f��o"6���r{�5�^ׄ 7� �^��5�с�#^)A�<gm��J<_����'�����X�6ߚ�����*ih[�h��ks��j3���=�O+Y� ��������Gx�����Q?ݐN���s�f��ñ��oX`���j�bm�5�6E���uڱg7��jc�w|^b"F��zN�/�ok��q�~F��K����9���Ϥ;�{�m�oG@��9��L]�{�: dˤ��\��_<Ȭ��g}J�m�Z�0��5�.=�.���&;kz�)�����B2��muF��[����v��&�ç�G]� �՘{�����CjK�����M�<{(���Ca��-<��|��+�9�T���'3�	�Ђ�߷ҟ)�	��,lL��!�`��U��]SUyyϹX�v�Cv�w�o��+��y������<�$j�h��k2� ~by��۱yUm�\���[K˒��O�׊�F��*�����5T�������:��c]�ݔq�Ξ��Vvܙ�U>�D�9+l�璻�9l�-�N�݇ �>F�^dn�Y����Z�Qö��],�J\�b�^е��j�����{�k����ȿ u��c�,��dWz�?��������&��On���aQΈ�؊�,��6׍L���,�M�_�+^���Т��$�Vcn�}���|y�v�i�&�ڮi�zY�c���e��"�LMT�>m�f��:��Q�\���g�Z�HC:l�$f���ݠFt�V���4$�#y.��x��h|&kЪ�v�e4���Ӌ����Ed#k|��7�rN�2"%b-��Α���L�f�Y7L���Zo+��wvL�S��kCf(:�*�.�n��� .�T�]�����&��D�]'A��>��)&Y�F�(D{�=�{��KJ���1$��2!Wє8gk}�%tz���oH'ue�c؅l��ͼ�iˈ��ʞfMv���2�N)��Z���Uk ���V��;��^����	�2&�x���gm�����>��m��z�ƀ�4؉�N��a/�Pf��ϛ��}q�S��s|X����gi��A2�t0mz�}�"Ř������I�S����=U�^�����5`��2�C@.֕;j/eM���Ú&	�qF�2�����_�ׇM�2�πŲ�t6�>{'�}�!ZZNm��Rv./�����t�I�qT�촌W$7}C����m�k,���ei��צ�=�8�VD.��)��d'�ⶒ��ՍYL�4u�X��[Uɪ�^��_q��-e�Dͤ��)k^�Fz��:�@���4M���IT�`���`���糮���x���z�3ն����@��F���K^v��?=�w��qh���w�Q1��%zx݊�1���捆�(Z%� 
�I���_Hx����@���*���P��ء�1�w`�b3t���9@�,2�bkI��l��<8J��g9>׽R���f��]�ƛx���s�y��O�gg\Ci��#v���qxݤ��/T��~Kk8g�Z�i�3�Ӫ��y[�N�6�r�q�Z�Js�m�뷑��]4?�6bi;�aB��v���m��Z�ܷ�7Jėox��P��'���+7����"�yޛho-=��}2>���>��2�
��g	�|y���qa	p���v�9u��� ��Pn��M�A�/Ωl`��
��YaA��P��Aj�	졖Jl-��l9�1�L�t�Ԯ|:��7��\��3��+wu��F��$��Jy����}y���"�g�l9v٭����w�J;m��tA�W^:����������yҙ���aEI���co�r��>�n�]d��8��Y�I�ѯS�3��e�8��6)��(K�q;Ę|Q�wP�l�j���y��|����&/a_����K����]ky�l��g0I��7[�}v�%��C�\�֏)���j���bmP�M�s��6��o[���ar�u��8�,o^P�5b�{�S[�H�v�L�pO!�fW^�{�Smp�~;�f��أ��me�X5oS״��yQ}�g��o�h�~�x������n���#Sy�$�f\k��2���3*���W6h�/)ME񘛩[
�H��a����t��ѽ��2|M�* ų���s4P�UƜ�JJkr���i�;{�Iۡ^����U�+>�[<u�2�<�7D�D����Z��S��acX��z���fNв�h�T
ǌ�e��z�򥕒�b���b"��7�����	e��fo=F֣v�����22�h�L��(ׁ:sxu�@2�,������2�l%�+�-�Ze��E6��mk��i��ϐGlx�1P�V�Ejͅ��s����)5/��dGUg׼ʬÖB��"��=0�۟uN���]�i����*���ۙ��y���ģhFu�cXvW�oHr�r�7<��a��oa��u��9�Y�e��CeP��p�˙�Ӣgh��%E�m�yH� Ad��Me�|XĆ�-�}A�3�G�;�K�M�u
4��'�N�Wy}�|aƪ`���:�M�t�{W�	=��i�[w� {��y���'��r� $��Τ+ݺ�+�q���ހ�͡�dK3������O���(l�y���W�'�,��f�:L1��-��A5�5P���m��w`�<�ٚ݋^��V�% y��{ǲ����lu���ir������sc(�����v@7+���{�oŤlc���;�Znsӷ���nΎZ�=��)�?4�$�w�銢l|��*i�kh�𖧹����2�b����c��3��=��Q�k���W�nuY�;�;��27P#s7^��TՌ�#-C��˜�1U =��9Bju�/^����페�����ܑx�yVI57XqU-�x�m�5R���+hF	���e�$�5"���a�XQ�%*�� ����ʮ�\\�k]ҝq�fq��9=�/�+���xJD��~���6�s�P���e�F*�Y����JQ.���V��1���A�w��P�Κj�ฑ�-�YrJ����P+z2Wf�#	g>D򯰞��ś&��:Jc�L��X=3����\�Z9�s2CP��w��*9H)��+a�_-�5�Wf�v�V���[vT0�`� BI��g���Z�F�HHP��-�Z�$K���N���������3��l�����d8�-�v|��8r�;b��/jd���w"��l�^ f���UBW�,�#��{OD���s�C#S;t{k��iwOw ^o�mwl���<��9>g��V�M����IB)���s�Du�I��6����^UoH+�+e�#���v��:�@�Y�.�1)4�3�Os��w^� ��\�״�R:�VZF/
���d�h�&��W���{�W��̍�Ͼ�������������8����1x��	ۤ^�>��ȴ^�R m�ܨ�O��h�͗��� ƢZF�m�����gru���d�p�m���ؾ�|�������iĲw1'�>��1�Ld4s�{6��@d^=�R�һj/Ci�;ӄ��xj@u3�j��:�� r�ҋ���֖c+�I �����������o��$֎��'�}+��yd�{mST6�_K�-�l����}�V���i��8t�/ ^ާ��W7y�B�y�Svp����������-�o#0���8��гq�ͮU�^��M$zJn-��ԆL��)r��ۗ��r���A��߯���חg=T�k�P�$4���R�zYd5�$E�S;�����u�;tD���P�Ϫ�HN�l��Eq��
��Vј�]��Vo���'�<����=6��8��*�w����N���e�?0|�;L4�2>t�\OG����g����2ɮ7o�ҿJ�#_�����(m�ۛ����N�{�Q��9 �ڠ�{2(e2��3�z���*k��1�Tٰ�K�v.��⬪]���]��ןq���
g�X��͉�r�l��O`�3 ޭ���y�i]-�{�b��
Y΋���Z�Â���l�?'C_.@���b�3��T<�m�ʅ����p8��Ǹ�9'fEbMW��V��0���!q���w�4��6�BKz��0����W
����3]�H���(��?c�딈�J�v<��;�b�n,wdVHqy�#C<�ƽ���tv���ns�7�}�y�W{-k�+wnF�<�z�����Wfd@I-�WN�7I�Vv�<S��r��5,냛덱Be��m8�,�wwf+��ц�ׂP��;�]�Г��ݐO1�Fm�"SԀ{Q���֜͌Q��f`�:��ta��܋��9W�=ص{�b;���9~��t���vq���nc"|��v|۫��h���o��|�ټ��Z�O\�5�t��&C�P{L=f�@�=�w�{e�����(��]���xA{D�cTd1�SF��u%ۨ9�7����6�ǫ~�\��7~p:��z���GrC'x-�D��]��Q��m�f<i�F�x�Jj/���eл�Ð*�q�gV�1z�3G+��Őv�v���`7\�yF�K��G����;�wCa�9}�wvŐ;xr� ,J��Y3���t���49�4`��ٷ�5S,�r�LNur�����^Բhɯr�k�fU�����Ǉt�J:�ݣqvcD�mX*'mP]��	+R^K ��S������s6�����	f���PC3�3�뗦� pY4 ������*�r�2q�+_M3�d���M�+�ܼ��X��|�
�H�+��$4���%�2Ξ[(Din��w��F�\�� �6����i�Oլ�"@x�tr;/�%}߾������I���\��l\�fn�@Kc̈́�a�g�w<�K3n�̢G=�ə������0mF��lql�#L�����\�l~r���"�t�>R4zz��r���j"�<����Pu{ad�R� �Ee<��]q���R85����)7���n_d�v�;��:Br{� ��S=�W�Q.��wsdN�M��Ǜ�Fљqܷ2��2�v���m���>�b��},�%�B��f�
��fi;��s�^�+\��#}�����t����|�qT�>Í7���q�F����ȫIP�~~7@�T����O��m�ѵ[ۛ�g�A�W��>_d��u"{�o5c=�n�T�^��gwp������m\�D=�?hR���<�3|��LG��c��O/2�C��7w/Ȏ�-��q�{~�3%������QU�� �{������/��.��G�� ���EQQ�������DD?�H���;⠁��[��4���x��8��p(� u*�� R�Q S��$H!�e@ �p�@ �~H��D�  �  @�  E)�  P�  �@ �@ P�  Du����4� � � 
 � " � � � 
�a@T ��eB�T �a@Q �(` �` �Je@hb`P	
VRbD�	X��I�haBbV�!�`��a�s�<�a`� �s�9@�8�D�o��t>�����b���"��L�̟��7�����������������1��_������������ ����x;���g�_�	�XT U����!���?�?�E�� b�_���@��t��'�������PW�������q$߁���?ڞ���"y�����b��p��(0�0�*�2!"���K
 ��!0!��P�R I(�D�*�J �D��R���$"�� �P�@(� �@ P
@RdBe!BaD)�B�		�@��I�		 ��	d@�X@��RD%	�$BVD dBT�D!H�`P�I$�a�H$@����s�C��o���?�"��� �( ��?�����?��G�
��Ht�������u���
�
�����������N}���g� �߶;?��O��b��G�J����}:���@H����(6�A�g�¨�/_�?�y����@g��0ץ�<	��������:?cѧ��8@t* *߳����(�����@_��?����ǟ�/�����������O�x�>�U {���?��@_�����AI������������A��??d�y�� ~'ډ����i�?�:�������������_�EEQ�~=�8:EQ�����������O��(+$�k1Ƶ�X)+0
 ��d��H�|w��UUT�UE%TUE@")R��U*�J��%(��	T��J���*H�PB*�R�$	UH QDR���((�XU����UPP
��TUhh�)(%J��DHHIE$�QB��JP�!(	U
US�E�P� �R�*��B$IJT���PJ%
P���(��JT�$�����$�QD�
BIUMh��)   ��m�JFL+l-�6$�h+U@�ATUR@R�SSXj2��kZ5�"��+i�
,��l��i$�I
�����{�  ;�  =
��p

(P�ð�
(P�A�� �RS�mlJڭ�J��m�ZJ��`6ƈj��k`Q��5VJ�SQ����"�R���jU	DJI!�   ��SZU2�X�@Ͷ�eVV�,E�Z�H[BM�kP�k �´�ж��-��(ص��U)Z��݅2�i���6�4X��U�TUQUQH�   ���@-I� [[5��* %���Tm�41PR��ʱTUQ��+X�4� 41J 6
�$$%$U�EHQ�   琅UUL��-��
�@�5�-bU+F
j��
EM��Fkm1�h"�L�PJQT��R�� ���Cb���L�T[)�4h& *�����Ef��DT,�"(��RڈZ��UE�EP�
B�R@�   {�x5����M�Q@�2�����0  j�`  -+  ��@fFh  U�� ��`(�f��5)A@RIT�   �*� YK  � � �F� D� l�� &S �4� 4 k @Z���*���QB�Ox  <  ذ����P  ج  �Z�@3( 24�` �3
� �� U�` (b(A*)U�T�(UG   8  m�  a�  �L� fP�j�  f�)� 3S  V  
��  E? 2��  h��$��M �M��e4�  E?�(1 %<��&�Q� � $�A1U� �YE�&��k�)��� J {�栌3�3�V3YLsW��ήk�I5w���I5 $�BC�!�~������I$��/ߏ�;�şʓ��L��V����na�`l�]�9E
/��ҡ�-�U�)�J�f����"�ۡ�f'{��e���������d����3>°�i �J_0�G/o@���4�AZ��+Qܓm�5��0�.�L'7�+1\m]�p �{S&Qѻz&9�5YGn6�����j�C��f:ݠ�F��8Y?l��x�0�`���ne�GZ��\3,S%
���cA�ON�8)��BR����Z�n[L�8m��$Ѡ���v-�Z%h�j*0=�ޝWb80����+�h`�Y��1tJ6��ZU�b�"�~��To)�1����2a5�fנ�h�l��q$���V��#n�i���m�oV\��H-z�8]ܬ�f�)��YX��u ����H��]�	��t�d{�R�U,'oX��P@vFel�Y��{2��!J�B�b�Kj^��7,S�@b@��-�B���٣V����¤dH�
�3�YRm�A��fj���/&�dV���C72=T�Ŋ�5sa-b72�d�)�tt3�S�]LEʱ�"3�k�W3�om�p=����y��u���[����Z���#6âe:L|5J�kl*SL�v6�ʗՎ

V�b�bv�^\0h�I�?X�@����QDV�����K�٢m��,x����YX�V�ly%�06�Ⱦ��2�*�L�3R+V�jI�'3(�p �.�Z͓��3�2��a�wq$���ղ�^5�]�م�5�L�%K�E� ���	���Z����f;
�5*\{�-�v�w��zI���Wy�5���!�/RQ���B��rSOȯܢ&��Ӽ4���-K��&RǸ�ıY�S��j��-Fѣ���
�>.����n���Ә�3i@k�d5p�;�,мV�7�2��r��6�<�r"*�;�u+�0�N�5�u���̦�6�M<_��A����2U�f��&��ʶ��B6��gT�y�eGF�6�Jv�V-!�nh��໒�JݙSnӉ��ܠ��n���ו%^m�z����j)��U�v�\5n�ƒ�Z�£��)7�a,�f�|��T O٠^]�� eَbi}/v&-�E��3@��`����mGu�����-c@�P�h����߁�G���<��m#OT:7&kI:h�*P��j��[*�ҷ&n<	Z�[p�x�:B�U�c��K+@�.�[%K���j@�ܪu���r]�]tj���O%E%Q�\��/&�Gy��t����V�k)Q������'3衄�kt:]�L7����QL�vݥ� �T�M��/v��-;L����{�NJJ�MM2��&cܫ�sNմ��Ǵ���������C�l�Xh�&٪#2.jŭ|�=��L�B^�Ub��^�]�;�v��S(�p�������W�q|�����+lm1kTMP(�RT�Cn�]�8v�M��(���VK����qEH)�mG6���ɂ�T�E�.�.=ZpZ��w[ �j� I�꼌Ԅ��X0�>ǂ�K>d������S2*��^�wl)�ap\.�R9xZ�� M9��f��j���#8�ԩq�,�E�Un�M����?X`f���]���e�5�&�q���V���+���a5	���G)K�n�Z3�(n5b�2m'f�3)��s(`�?[��vqͫ��*�-@���̨]'yS�[��,k���4�Gur[2A��.����V�66�:�f�uo.����e͒�$������&����,?�1[��^5�f��$�N�#���ڲ*�Ƭ}��nXD9��ۑe)R���� 2�gq�.�@�@*�Yr -M���h��jPյ�
{{ғ2����� �J���#(�Э/I�ˬ�+`�)�8㙔�<td/�*=,��M�)��Њؤ�OEL,�\(�J���ޜwlk�Ր6���lK����[���V�eh��fļE�����h�wB�Fc���8�VC&�tt��Z�:�+z�<�.�7A\�(QJ�%XR�z2��:�L2�2�u�\�X�����a�v����V?���,z�B�AE�a�v�VD�1ޡE�^�̱N��l21��v���$��U��X�%dH)�jP�Yb�2C�^�����(�4ܤ��V�a74m��nR�qi���7tZ]ٷI!�[�x��W6�*�./��a�x�I�JTڳ� �xZouՃ`�Ma�V����Pz1��	*��-B���zUʷw�μ�Sr���eˉK�>FJf�C����[�jhM^L׭��c�1LF�̊�-�MM���ݡt��3(�j ��t:7̚���w�l��hF�X��Fں�(�i�J4�i:f��a�[��-C��e!�jٛ��j�����C�.�a�ݗ@��f�W/fJڻ��6kT�M+�0/]`T\8�F��vd9w`bWh�u���R8ۋ$�h�(]�� �Ȩkv�4!c�CK��81���&�E`��n�J��&#w���Ÿ́�!b=W����G�ݻyj��A'Y�%*
��T�r/��m@�ѼEj�85Z�u�S��d�J���96�=0��Y@�x���࿖�cV:,���Udy1�����7kr[I���S0�\5�YI�46XFVk4�|��nR�W7)!�1'o�z� �7~�b�靽���E�n�L��r�����p@�eӸ˸��"n���lTצ��w�2���٨��1���\Û��z�N'F�Ќ���^ +�qۉ�� k��w "��ņ��[[V�OS�U��W���x�3|�ܨ�G��{RƴX��H�ɡ�����m��ݣiaW1�:.�V�6b�&�wkh���SR�DEk��a=x�R�OkvI��v�]�N��04��6M��0��S���h�ۏ�b&n^�� �ݡN�q��f�Ҝ�ګ�D��� �5��àt�Ή�p��d�ٲfCp���k���:PKZK)i/�\�*�e���cpa�A�dSN[��
9,F*BN\��\�و��872Z+��ѷMhՅ�o�(��YX���&�����n�7]G��b�&��N�J`��a���y�T0��f�[lb���6��:�e��<˓,ə4����f�����c1�/ۚ�~Vf���w*�����CD%���52ժ�Sw)��rRU7놱�f�eZa�H�ٛ���!�R ��ޗ;{��!hON�gr-�Y�Z9�S5YA�+^��B�U]���or�#V�oC����M�&#�k~�+�h�Wm����MkT����/nf;�n��vX5�5��F"�k���Lҁ4���P��b36+zU�ct��Y
��Ut��M���Z�0;��5kܣ,&-�v��&�6�0f=@=����d����ͭ'��J��+j��a���k�b���̍5qm	�4���%���Z�����`��m5{��R�C�fKI�YM�IH�����2�����Wl!h+��dX���ɒ�K5��Ѝ8�����NZ6�<����ا$OK�`�e�v��Q��n�0�/��%�Lc�³"sU�n���	��àA�E��k���L��6�eF�Ĉ� Qݒ�Q�yw�b��܆��i��,աA���7lHf���x��זY�mI4�L�
{�ǔ�W0-�0��vf;�Yx�͚j�i��%B5�m|�[ypF����-]d��]�-	2G&�h����B�� ���7v����i$PM��;�dPn�2�P�K5�5 ��+�cW�5����
V����7�������4��e�=I�aKݧ{l�?<�aWK��7W�WHRT���b����Ьl�E�CRl���m�M�m5�l�C#��rT�rnZ)-���AZ�YX�'!{�[�["�b,��v6�{�,�Wen�z��zF��C�ZZ��I]in����H��ɋ$jS��c���� 8Y���:[�Ô��H6��4����
��q�rPԅ֊!RyJ���\V�u�0��T5.lcby�&��J�]�z�B�A2���X;$n&(��(�:D�p�R�Yb`�P�A���ch�Ȟ6�,��/$����U��$��YHRb�`����1��:�ef�����e��-�ё&�=8ĺ��:5,Tեz�n��h�4СZ��5z,^:T����4r�Jyp���bZp*��Z@ �m<�7g*�]�X4-�f���1�LM�Ҥ���Y�j���Igș�x��;0��$[Uz��ԕ-��X#�1��؉[J��	�*�
�ϝ��+����S��uz/2��(8��̫��t½�%'[O$dV(*�jE䶰fc	�+m%����0�!�QP$��5�{L�yY%���8njQ���e�z+tX�Z���iR�C��5�h�[�J�����y��#��N�b �[�7BQ���,`�a#��u��6.�n&\7G"�T��"^�7��nnեd�{��	p5�n�XVp�K\˔�R����)j&����2��;F�X�	��Ӊ�p�nT���1&��x�M��Z6�-���MY�N���m��0I��ԡ&��z�c7o"���n�{>�F�N�4��sc���bb��3P��(��{me�h�IA\fQNY��+�ͺ��b�rӭ��,���A����h��\�����V5��tF��Y31AJv�<��۬�F�eC���
r�)U��!��YH�� �.�X��d4��/�;t�,7)l`��6�elq�� -kG�m �e���K�Smڗ��X��9[*A��6�� ,YV)ʼC1�����IR�J]PPT�x�vu8��:���+	�.��uX�	<8&Ky6�*���N�A��5fh
���Q;J�4Y�"n�,��B���Kn�#��	������4t�������C H]F����j7���ʉFf�(���QWIQ�;�~%��.��6��]��wOv]ԉZ�l�"w�+3I�$���s$���FB��:h�wDӤ�mlϚ�l%\�f��ӹ7VM�(D�k�n;��ؕm��d�k�߰S4tA�q�K�ti��H'GV<ak�K��.P���im7�RY��� nBI�Q،h�̻�o	&b�G#�QI��L�7T�X�d̀��d�=�*���-��x��3ʗ>���̩f��i�2,H��Q���$�8�wF	�4��,���>�I.�U���DXE�9�����Lc5�X��*㘕�{O�j����5�\�N���T�������Ս]�&�]P�n^�h�L�7�V/-�N����7Is^�$�Z��AK���&m�oC�L�go8��0���Ǎ�����V�w�Y3Ssmi�`�X]24ʴe`:�@�D�-GA��� *�D4�p
�z��nAF1*9g(MB�D��e5,5Ok/h��E͗ �dO�S�c���]�{�`��8k"t+h�ܫ�VCףD�v�u�+�xK�dm�y)�<6F�9(�J���%Qh���a1D����o�MS��[4j�/��-�S
Ѳ���j�m��A��	^]cA�ZƌՌ^,���t��ShX����,�~(���hE�x���Be���sf��̽H<V����7n���hV��E#�lA��׻�� J�m �.�!��a7{�Jg�����*����Z��޺&�d�*�ꎡ��Z�ܢ���[j��LyXe����/�EL���8dGk�]:���H������71Ȱ�\��f�^lF�
�𛡌����-�V�>ܫ3e������:���Dj��7ef x�m��"G,��Y�0��\r�33l��nP��p9X������|d�ʈV*�J�m0��#��?m3j�4D�p�hМ�A��:��Z�5��n���0�5�jk�T��n�4N��IӒ�sJ�5
w� T�]�QIcv�v쥒c�%�iT��R�{lS+~X��0\,��X�c�jl,;�B�Q�Pyg*d�-�׶wsܘ�b�J��*U�yX�]�8����*�0���n�Cc���Q�5��3E��/f��+4Pӷ�e#��7��Z]�t���L�t������Kr�D�:�G���6쓦=n�VøT��U��n�ԉ�����`U��>w��l�w���N�Sf���Y1��Z�#2���)1h=t�O��HM^$c5��WP[{��GG���n��u�n����Wt��+��*�B���A���YA�,c��z%j���`�zUj*��og�S�,5wMU����3oi��QvT7�vT��TrnainL1Ag:j��������xRO���(k�����[(��h��`q1X���@;���T)8�*�Z��#��[9��E[���c��.�hnі�[
��2���e$�⩠MXs,�mk8\�ض�ı�(��!�E��2�t8���dCV^���Y����3��%��K#Ҋ(��G�b2�tU���^RA�ĕ݄�
���b���\X��(Sj�[!�%.���A��J&#��TF��Y������u�)|T�\�Y�n����[O\��SC��E�y��t}{jM��QU�Ol�N#�m
�/��q��B��D�U�?��7�e20%q�I�U�0+���������R7$�����{�b�f6��p\�P�쳂ڹv���S�1�xund�XZ�����v�s�,,	i�s� y�K�Ca�qA�6@�V,�ӹ[c�2�TyR�n`���x��[7���K��\���ov�D�u���������|�I�u��t��6���ڹ��tL�}N���4�9B)o�{��1S͉Vu�Iڷ;� 6�!��ǡ#���8�m�c��L^l���|�lm#Ű��o.�#h�u�^�ڝ��mP�O��sG*Ҕ/O��I�qV��cc9d�G��:���(��3�p~��Ҟ�H����{��x��2fECOu��m���N1	ܝ���&��4�^�ӱCv��ݡ8��y����E|F�?C�=˖f�^ �\�Px�iu�*�w;����U.��U�/���
�i���R��nP���,B��m ;Ugq�جK��Rۣ0�b�7`V��;�X�B�v[rӬ�wP�P�v���x�[V�4شw���%���Y����]�	������s Lb{������0u�d]{i]�U�D�WWB��Q��������9�z�K&5OZ�[O>�"��]��W9��RŋA��gM�^�`�0{d���ꌪ���އq�6�8�עc����B�k�F�s�n�I�W�c��@�jB��7���F�Z,wk��;idm����t<����S�V�*i��� "��� us��=���r��j�`���5{N�@Cr�]�ٗ[[g�c�޺�J폳ԦY�xG8<I����b�����6��B�����$l���L���u�v01������o�%r�u(�u�{u��U�pkz[����ùչ@�YS{{Mn`@�
`fkO��_ϸ����tK�4�;uj��ffS��N���e �7����Ѳ�[="}`���{���)���u�8�+o�}���:%m{B����/	���<T�)ҭ[u�����#Mt��wݱZ�,�lMۂS�]X,(�7�����T��V��X=*�Z��#��
�n�_r�;P�Qv���;ec�fl�-�g&����`t����ť5� aj�FR�|bL.#2���G�N��:�f�d�Fj��ӗR]���j��^T�3�K���H�."�5�gQaR�gn����+W��V�@WE��r⭗����FV5�Zvk*_u��;
�s�1�T٘wk1\}��S�7:�R��3GR���`J�@i�@�|�L}Gr!i��}0S-�fAóS�@�[֜cyU�\��k[�6t��Õn�򱡦�C�&Fn.�/�6�J-Zwb�{�\��L��C����������T�]��B�i���0jr��3+�}V�Pb��KF	y�+k{4�v��G�[����%�	F��i�����/:�<،����k�3�=�E�^Ƭ.�����=�ڰ�jm7C������Ќ��g���X��E�|	�Δ=����(/���6Nb}�%>��r&&�R��;��䙁���P�0,�+fPͮ&���㙙���1St6��b����g#O���n'}��H�qYIw\�6v`U��3���;�V�C��R��WT�J�=Æ[n�1��>(�8��e���T��0��X��n�0l�X�Ѱ-��E�2�÷J�al�e����	¯��'���E���i�1,�������1r��c�+����i���ٚb��w�J
�,,�X�T�
�M��ق�.�\�3�Ù2�t�r�,W���O��,p}L*���[�+3�,�.�]����bQ��]��!u���pJ��#{�^Exs�,�v5�Z��c�~��~����(���ӨXyq���������yO���b��i������\��=ަ��p��Y�N�}I���wX�(�r��C!��7� �P�GbѢ�i�Y���s��M�阀Ԕo�#w��E����Y]����:Y�z��n����uX��VL�KY(|�+nvGс�
�sR1E��c��ʝ0fq��,�ܾ
ť�bk�M�x�W�L�4�,�i���dhR{Xv��eL��M!�l;}[PF�*^�]�W[�ݨz±i��T�a[�=�u�qjƲF��|xz��u^(�+��R����-�[Ӊ����f���(�Ͱ#���g/��U��gokͦ�"���3yu�r9X3z���%>�	@����n�X�� �!1V��	4.fE���4�:�b��x�LT��ܚ������ȵR]4� /X���*�c��u1��r�RO{�"F5Omr���ڦ]�}�6�)���	���m�GQq���,B��ͺ����YoQ�h�n��1�9qz�B��Y�Q茒��27wJ`�s���.yQJ��1���^U�-��P$��	��z�Q�4�!��\	Yc���:knźz�[��-��eɖʖ)0�E�����M�W-Z���{v���貸���4A��g,�W˚��� M���ƸH;��ϖ�]��1�z�䇒X�?�&Jѽ�F4��/o�$�³*���`�ވ��G��k"�Ժ�l�a�}�^Ӗ��M���j֛(o�q;*ZՕ5Z�[�si	=���Mj�w�����$���e<��1HE�d�kR�^�L�g���ڎ�}�u�R%�r���XS�-,��j6�ָ|��A[���Toc	u������m�_ctq�j�����9Y8������6�ێ�.�ȱ�<��޷Q
Ϟ�BC�c*��mZ�.�̧�7>���r<��;�|��=L�>fr�9�|֟xB<��U����Z�Nt˽iu�-YNu��r����%��s�
)����W�@Ժ6��1o�9�ܘ�M���
 �-ܾ(e5T�G�ԯ�U\j݊�v�b8��=�7-진:53yq·sp_Iâ�����t�6�1	a�n�9J�E�svX��+��GW ��wunpv��� M56��7��nJ6��Cd��復b���,|:�`��`�5x~���3�*��.��jwd�6_Io���&�[���),��'.��J�r�.��
N�/i��=�Ѭ3h&^��GlN�h>BY�s3\ڱǮ�͠���w�z����Z&ew�� )Gh��ei�w�r<�V3�M�����aN#O��,�k�� 0
�F��=��i��8��'j�����}�c��ZV�W�V�q��Q7���=R�=k�,.��)}U���LT��g�����:a[e��L=Z����v�2�zxG۱�2���]^j�`k��%2��NYCl:8�)p�g��y=�Z%R�<�E,A��u��Eܔv5@n���r�}�U3F�"�I׶����d�l��0e���Z_B��9�P=/b�봘�O�R���!Xwk�Ɣ�{V��V�6�֮�Ap�䡀��N�����Y�R��En���|�L�ёvf�t]aL��4DT�
��BilL'�TGQ��jgVDMeչ��r��LY��k�\lH{�>��[tu�,�mn��`��K��'8����`�e���l3ސ["tgv,��j�H(�XN�5A��0�#�w#*��M+jj��*�'p�^�&����[wF�֧+ls�zz:�	>HT��Tpf�����iQkZ��u��yw_Yc����4j�U�YЅCgf�*d��BݽtKc��>�јk/x��ۦ�&7�:�su��q���U���j���op�ȃz�ƕ�>�\�1� p����&V9U�mD��Q��fX�V+�[��bT�]�SUQ�em�.�q�QM��z^��]۽L����[�7���gF��G���\9�2��냬�����Io�v���s��V"�ٝ]vX7�'2Z�)*Y\x��-��7lu�!S��lX�2�vVa�V�c�h>�Q�0��x���:n� :u F��ᕀ��#/�J	f]N�����m��X�#,)7��7��!r�ot��dE���'�MU��s����]�k"&�s�[�}l#J>s{�vnK,!�4kݩ}�Ёz0议�p̟f-k+�-.�Y9��}�k�K0��=�w��]�ߋ���v.S��Ӽ�
��+�z�D�.����p�h�ǳuWM�ӡKo��g
F֝83������{X����7��s�����ً��z���S�}���=�Fm)�($�V��b>#+Mgq�Cib[��[6�	0�46��%�:�4z�$����J5�E�7G���������W/�U3kT�jr��<V�N����xq�
+Q�m�Y��	s���j)]�D�F�ad���A���7��8�s�N�*��$Kes�O*�YK5�%v�� eٵ�Y��B�/���4�f���j�&��n�-ʀX�%>np"*
��7++\�`4��r��Hw1j�ql�w�q�hev>:��Ի�]v��̵ΣH_(l�շ��=���:��)Wɟ��k6J���w�w�Ю�9�p��[Y�,��	�Lc��ܤ�2����G�w��ǰP�wZ����i��7�v#x�Vium��!�:e=Ǧ�U�Yi��(5µj�lK�A��*�I�-g'���@���ho��Yg��lgi.��ڒ%�Sz1��G���:�+�Z�!M��f�Xz�u�)�6w[���H�W���U�
ݡ���wu�͠�}�
����뵍7�EX�q��\q���2��� _}��z�df�C���d�/G_+G-�PR�����6Z?f����7��Ʒ�Xk)�лsmo�m�
�#{E3//�ֳ���B��t�����/t�a��.�:<���wةAN ���ӹR�Y.
?XXڢ�bw�U\�w��u��h�}��:����Tݓ�̘��9mٮ��C�L�4�Q��~�,�uK>�V��x�V��E}:���=�y���6$���\�����t�����8���-I_�*�*��|�SF���^Q�lI��gNT�q\��f��.����Ԗ��<��VRzy	J����`j����d{A|�s
�����r6̄0$.�]v��gt�^b�e�u�z�E1�VF��e@N�4�rv�ٙ�ذ˭HJ{�:�b�J֥t�M�棸��p�8-����d��9x+7A�Ya�n���3a��P��T�R�ʲ���P����y��(/w�'z�3gR9͝�����D)��za�I�fs�Q���Uo: o��á����-�Yh5(k�>Ͱ�#:���2����9�`�S���|�|�7Հ�ܪ�94���;��(��W�i6���*eXg�*7�x��]|����[�mծ�tVή�V25�Fj�;x�U�<Y](��p����2y]]7�*L��rL�9S���'lݽs��1�-��"^�'�����P�jhK��Gj�=�J��7��MRp��j��φ���f�(�ި�{a*�V�@�P����.���g[|�94-��,���e��l�b��SgsWԻ��[Ahf�c��FK=���ock� �߱�;L�%#��7y��%o�eB7��V�)l����F�͢˝t��	�G�ɕ�s�[��+�&��o�0�;Qa5����^H_��t|oZ�Ӆj2���ju�Lڼ����24�0�{��--Q�1��"�4��tk2Y����\���y
tƞ��ݜ̠�u�X�(	���nM�t���oZ�����pgg�M�*���Xo��l�*I����=wGX�ؘ���d��U.6����T4jNӆ9��Vv���k���&T$ұ�v7�t������*�t�,m�Sa�!�/7cٕ{ �&���P��޹���5r�rRLl��M:oC75��2�+��\V؈���+C�=`P 4���6�g*`Ɲ��;#hJ�,�]Ά
����8�]�Zc�P���|�	��Am�pֱu
U��so���.f�L<ήˤ�9y�V0���1򺜮oX�kr\�}[���N	���..?������ގ`�t�<�Zr�Vb�O-�x��a������f�sO*&�Z��+쮹{�o�U�x���
)�~�u�M�)��W�<��v:���lu�w���Š�u����(Ҹa+�v��'|@�8�;vP(�]�ff��ň�VKB{sn�E��F�.#{��(m�������+�YRm�������p��O�[˂Z�4or=���Q���'u��:�b9(�PhL���m�v��w\������s��C�i?kU���z��ۺFC�=Ǳ짱�sp�[�2wUCM+E<[z���3����L׭uC8Ax�=����� �9e���lҺMp��x�H88�wv鱶$T�2�}�֜��1�9N�P�ޝ�(Nn�7�����7)˴���멖�s�-p���Ma:�Z5�v�#}��3=�`Ŏ����x�e;��
�g<��6�l�˺��\��\���8)Y�HPhr�9.&j�����Ζ�j{��ΆgR�f��۠�=:�)U����&au�F$c�`<��y�e���[���"���W�v*��ä��8�mo5kc�1���=˻&`
t{3E��K��s4k�1��s��=/;�W!�K������ʗ�P�E�JAJ$cUe`�\�».ۍ.����"��+�?u�HYڼ��/��n�����o:���ӑ���5lpR�i����F]ޏ��Ȕ��F�[[�	�t�wVV����R�����U�Eׇ�t;g-����wt���U��������7ݺ�v��+��ʀF�*W˼�pYݧʺ�]'1L5�����gD�Yz�n��yā���p������q1�I��I����Nuzwk2���䱶���V�|F�y*�O��ő��t�H��zia�2lh�ƕW�W'.��0뺕�6�X���v�Kٽ[��z2� 1�Z����U�>νΕ���쨷ut�t�.��	���4w9���˹�X�o"�y�3��!��k���u;(����:�M���+x�C�"g�t\0�u�����uN��Av�j��Ռ'B�'\㹝u{�Z��&�Mw.��ʾ�����!��@�$���9�kU�u����xm�X*�yF��3W"�V�}vQ��:�����Y�2ve85�ux�ytw��R����(��幋+�\Kj�� �C�\=�����l�y�nЦ�i����_�� �
n�9q�4l��y%'��K�h�|T�.���ݙ����UL5{�.�א�rm�9+��v�a}���{!��
��zA�i�t^�Pb���s"Ja�V�=�K�νY�\��ŒQ�/S��}��ve�ƻ�ל�iM�J��l�1e^��=j�U΢���!V'E| ���|7���,=�o�h���+'teƕR�64 ]ɩ��VK���� �U���r�X���<�,�Y	%r�
鮻3h�/�;m�f*�7o�2�mҎ�}�S���+>����>�MnԠwwȧ���j�+S� ���-�:]�l�'N���zD�Խt��':ދ�(7�|;�h�87�n�V��6�IOj�3E(� l��i�N�֡;�*�0���nA�)����}��Hې9�`�)�����b�7��^���+-�+#����q7�ɏ�r[�������}
Ɂ�\��1üT��k�EC�^�d�>�N�n���w�ec�J��|���ռΙ�i�әLt�],��NQ��>U�̇�gs\�cA ]�r���᎝��+��qm��zM쭓z���AJd8���I�ẹ��A�N�_�u����ނٷ-y���
��Mu��x(L�Y�U�I��1mt�[Ǣ�T���R��r��[Ӣ��[�L�ޚ�d=]h?�hw<Y�J�ʑeqd
��hTxz��S���f���GJJ��z��c���6*tS�%����9��� g9yZ�Xy�p��CPP���'����5��6
m+�k�����[��i�ֵ���v��o�q�)^v�/���8��pK�{.�!pl�\�����nվ�uр��C�F�F����|����b�<\>sQ��]4a��f����sHI���P:$m��7��G�y�^����/���i�`y��N�)D�n�4o�&A�f�)Ҡ5����Zk�qr�K7ɗQU�ܶAؤ7�����r��%k�D�:���)�W���)�2��C��8E��k��j��K������\N��VЭ���ޠ;$,M�_�"']K�B=Kn�މՎ.WgJ�z��(|*�'��(�\v�8F��g���Q�)��v��D:�� [3��gU��z�M���&���T���`
G_���z�nZݧ�.2;t��񷩂�5�z�5�&]@�>S-@9-��m��#�r��O(Vs�F�X�Ŷ �6��#�z�F�b�	mf���eJ�H��j�|N�6OW=��AZg:���^K*!2�`���E��8C�ҭ�=�[n����� �ec��.k:����ؒ4R���U��<�ٜSέ�s�a�l��bEle�F����u�.d��X��[[}{�*�XZSrI�[30�]�CwWa��EtD9��+�������EN����3�X�K��&����`��!��Qlnud#Y|�hP"�K�!��,�`Լ�C�։�
��S�	w�E؁¦�>�D���+xu>�{B�p��'��uq�H�8u��7���
xe�2>Xɗ��qC4�JO�fJ��]m�b��E۹�S�]V��I�\�g.[��^ad�����vw5�r�O��ѥ�M���uy��nX[aѽM]_.��Gai�����J�sO�|�'M(0h�[B��x:�xDU��vS���0�c$���3#\�`ށ�{�*��WE>�䵘gn=��e'���Y��>�Uy���s7��<Ǵ��9�������m,�^�yr�,�2�ԏ�8�$Jm,FE�XVg
{Lܱ{�����!h4�-u(�%�\)¯]
Gw�U��
wJ�V颁b1�KU���D����Zy���bO��]��m�Z!���_;�ηU���g��]�?����կq�jgt�+���[LV1�����ԯ�Z��9�_s��_<���[8o\}������ӓ�4�Š^�®�R�
�Bs�	ە{�˪�*���	C�ƅ�Q�7�ʸ9ik��"3 �Gb2cNf[ws0t����&
�F�ʔ;���^��`�����tY]Za�6P��1�8!�NMczh\�ܫm��&�"0�U�\�c�uI��0�v��q\����ʘ��m-����������D�v��t����X#p����6k�qT�VZ�̡bI.V�֟M<UXj������i�t]D�������Y��B�'[ٓ@y ��ސ3\\�\�W-�������a��uh��cXw�
�4��4WE�_@H=n_����/:Ct�rmr.��V/Hz�Y�K�ק�5���7֛�=���+��a��h�>WF��+aPq�]xó�e��}�.]t������s�ҋ�f��;�.DMWmZwb�[]��r9��VFê�.�m��yk��w1���l	���p����R)�I�:ܙP��qB��I)D�����U����Ȟ�<`���ي0s�s���[�9�����Z�0��������9Jxg��0P&��+ĵ*�^5jcZ�!L����V��cR�`��&q/�R6��xE��f����^�B� P�VtZ�䐠�}��@��9��4J�Y�եF��7l��S��˽5-â���GW�u*�:���Y�q�l�R�����Y�n������x�}��P�6�u��ԕ��.�<��i�t��"��tj^Y�5i�Aeե�p���+�;�T��ذ���(bq!����j��L�@j����xJq��]6��Uب9%�q-ZrbI�}qbע���jy�ٽ]*{������v����i���\����Y����J�WK��EX�qQڵĒur�}&�U��������S�3]��WxґYO�d�ho�^���u���q:�J#
ǳZ�n���˼�tô�GωE�u��i*ʓ�Reǡ��:�m�C+�q���=��kA��97�:�z⾭��M<������s�۝�=�b�]؞ݾ���V�Rz�ulZ �c�ODm�@(��V#=��&�sh�N�X�r�U�N��d��v�"����w	r2$굑�]Z�]��b�?i�dc7g��ݙx�MB� ]�v�ᬌsr�q���t�
�5�]�+��$\)!��_w,b��␾��5g��Y�!U��8c�*[�5���r��<B�e�P�5lWe]����q��[��7.;�7;��:��PE��;sZ�.yQ�}����V��'3��̸inV��ތ��.���b$�Jq!��;2�JCJ�@A#����+ڰ��=س�U#qvrHl}��871[��-D:S1l�]ubr�_s��Ҟ%\"�PQڜ�	ګ5u�gFkPT�iJif�u��;r=$ճz��P�1@"��n�����Vc=L6�'���tѭ7���Se�t�XqsVY�D�H�b��U�5l��aJ�wb�m�cZ��&�.|V'#��pI�	�����7,[p�!�0p�v�]����ˊ�k��UnS).�m��h�hv[;��Ԟv�c�q��ٹ�0ՙf�r�j*��q����V��%B���du"|�*2�ݦWkvbr�ث������}0��9�h�?]�k�=75�:Qˏ���.�˷��
�瑅*ڥs[&�+��?q�͹��a Fk 8��w ��V�B'X�R>U)����ۑ�]YO;�8ݜ�o.k�r� ����&it�α�[�N7�c�~�r�W�2n
[�Ne8$3��G��v���=d��:���Շe%X���ޝi�`gD{�zٹ��H�r8�9���^���Hv�b��wxyN����I\���]ѾrA/{w���\���b�Q[:͖�ǘEu�܉�PT����k�[�����Z�gT�J��^9����x���|_3�G4���6�&�p��jƌt����݀���ivQ�J��V�P�-hH�Ѷ*�a�c,,�f=�k9�� ;*�Q�x�ar�S8n�㕚�xi��qs���V�A��R0�~��֐f�v&$o5�p��׹�lu�v'�in���]y;��P�#�EU��ŉ^�p]Z&m�M�F5P���<��96�T?T� ,�R�3)3������Vk&���\�«�`�`�iu|R�v#0��ɝ��!V ۻ�&�X�b�Dr�Yz��آ�grJp��{����.�_��ʚ-�����5�3�Q�����]�v��i�\��VP?tG3��g�r�g�T�;�i��f�۠�WJr]M#4��<u��Vy�^}�!:�v�v��!��a��]�#��z��ޮ�p�3j��&��|Fj��H����.�H��R;��2���n�yOjc�d�
�8�VO>�X���,n�Z��#�ݥFX9J�+R��J��Ι{(6��hm��O�\�_w)� 4���ֹ���1p�[���f�[r�]Z"�T��G}�+�U-s�v�0����s��N��}�f�k[�	[�/�C��D�p���`8Z���%I1|��-+�۹w�����"ײcoP�K<j����6ya��|"ἷ��N(jEb��Go:E�ݫ9Y.�E�:�A+ڻ
�4�ٙ�����P��ݹȱ�r����-�sz9���${v:[W���e;{��ތ�n�cG3:�m^V�5N�Z�n+]\z���9�X7�i�����JN�b�v`�:�s7�gL�o{@j#jw����� W,K��`�Tu����4Z�h0��k�q���S?�/���B���=b��;m�1���)�N�`�]b�j�L6;��S8E� ���v�]Q��݂,|Ks��M�C�<7X!.����EЕ3,B�C�K�WO�����ݸ��T��A4mnt�p�Ų�:�&����d��]�k��n3J/&T����ap�r��墔�-;�Z6|۽���[X��%���V��ݚ73�l}Z�T���{|.�bYu�,�%��%�@U��d��V;i�{�oD�!�DżWw��v_Vh�8X.�>'�C�il�Nh[w�)�:����<����W�1��gKE���t+���������)�;ʶ94���ͮ����{�VfZR�C)��Cb�*�Jj=��[�Gq]����{�Ev��:��AewW&���-�M޴����4�|�Xұ͹%�JG��}���-��wm�G� ��Ifjެ2A#p붩���S�W�c;����"5�Izܮ��^2��M�6ew3Os>κֆ@���M`�عN��,�| ���:lB/����}�S�t66���Ai��#BX������G�TK"m�q>I��)�eIA�d:����Œ�t��[�j�ƍ�9���ٟLt]
��v_&���$6�j��ovv��(�M�k���M�j�y2�%@_tS(m;3V�.�J����H7`gi+��Q@+�6�m�
�jmM�:U�;���b�΂�<ۏ��R�i�&u��z;
g}�ǚ�`�޾����-Π#�5'L[�r��j�w�G�Z6�2hw>�������d��y>VU�䋫�5fq��J�M>��(i�o�U�J��d�}�b�[*�]�;0����Y6�-w9�<h�T�#�馝_m=�X�تg[T�_R�fe����q��w�V�"k�Wv�]�<B0�4E�d3BBtj$tL�)�q��@�Kpi�DJVV�\J�szѮ�$�M2�q˝nIWS0q�l=�ǯl۫�@�Γ�}����'G��67k	Wu[���a�,e"l%e�6r�Ve�L`u�`�a�Bͮ���d&p��ơ�i����N��6`�ξufP�euʡƷ�=��3"rD����/]�F�: kӡ��}�n@�e�V�{�}Cu1[6�� mN=�5r>�,�����y�epR>�b ���_rV3�{� ��\���*;ʺ1�s扬dMu����nGv�^r��6���_t�.mO&eK���bx�Q�S���WL�X;3"5��1*��s0q��45��>�oW��c{�(�U�Y��UŞ��1�P���� |ǧ����y��W���7�f��y��l;������Mm�׹]�*(����q���5�x-�UÝo�ژz�������{:�I}ntlwp���{�ۓOK��ѣ�!����B�%p�z��4�U�4����j�1�C��Y���c���&]�	&��+{#�E6L��V'R�b�n���y��E0T�N���e���6J�^*�N��ǅ�֋�a[h]K"���R9�i=כ���7Ckg�>"U�P�[�`E5� �RԘ9�6&��^_�i�.�f��ds<�m�.mڧL�F����5f�v`c���7�Y�gj����A��f�k*��l3V��.��;��>q��#�	н�&����G�̏r��%�Gv-<��p���t��jmN�I�Z�Ov�����y�l9�q�=5-��|�[�m�VW* ���ˑRupeg_͝|�i(�BM.��f��7�e^�8-&�TM�)"�'6�K��� X�^�1wuѵ�Y7ן^�g�U�·n����=��!e3S�5.��tF�Փ�TH�����2ż���S��z۬�C%�
��-e�V�wo3V�Xe���R�<���wW*�vX�z�I���r.��Oc��mC]ό�X�"��̹nm��7C�#N�ՓM��q�(!d���ʳN�k����9�N��W�_'�����s;ÛZ�J�V������]
�jSЦ�Xo6�ߢ�]�;$gy5�E��6�4�-U&���L���ѷ�X�})��şXl�j�0���ue[��P�I-��sS���bNQ�����[}�b�β�K���dG��oW���!	'�]�Ο�:YӨA�����;!gQ����ɭL�ߘzh��q����be<V��t��رô��Yjr�7�]��ӕ�N�hڒ�=pur��,���U��8�<�E�j��-��D�y:]k�e��A@�k�s�Ԋ7�w�T�ČXz��m�C2�)��|@+~��^�*��1�ol-��jN|ėٚ�|3iJu�e��{:�sI����ܰs��J�b���g�i���L|�^�'��kT5�ν�δ8�I@��W<�P��2f���f����ܦ�>��֩����Y�.�Lj�3HTZ}��uQNuٮ.Eg>�M�=m\���V�R��@�B�s���-���y��|9��S���5���\�S_@�F��2u���w+���i#,U�WN�
�r���Ƿ$s�V�^�mT	�kZ1�<Y����ur�n��R*�v,'�T8$�X�-�;�M�X�o���wؙ�3J�|-;��'�yMT����8QۗǮ#D�bէWgV�O�j�w��2�o|�.�,D �ż�Z�[D�������L6��Y�s�+�!��9뾮4�3$�Sw��u�RM�U�׶ }Y�b�з0z��o_Tr�!�{��K�Y2eR�.�2�vt�K��[�ˇ��k�����*�*�xh��c�ëI���7u�^�E#�Bە�^���v�T1tn�t�K�o���o{�@?
P�Ҩ���(����]�(�hYs���I�eqDS7-*�-����TT������H�۞E���ft�,[F�I��]T��	BT�D�jk����Km9��B�e����F��iIa����d�;
t(��.�5,m��\�$�hڕ�n!����fӑLӲ3� �e�!b�]��ۉ5t�74��d��<�,�<�t�I��D�lZ�DU�/Q���f�F�llX�jb3�͛���Ɋ�Xٖ.����vf�v]��dei2nkjaV���fԣӛ\T�
)���T��IJ�I*��Ĉ**"��Ehŵl2N5����n��y�^M�K�ui)V(��h\JQ�LBȖmRgn�Ѷܦ���%nt&��C(��D�Q��GlD�/)ڞz�g�y����U�2KM��x�ð�Q7L��2�#�X�D����(���q��M�������ْ��1�j�N>즁��n�8ݫ�͘�{Rt��q�ʰ����qOL��Ӽ��ǁ��Wو�A����b� -���Y�
�n�T�ju�mrνሁ&�(�T����'��V3;�t2������p���9�<���{A�)^Aw\���+:5���x:z�k�/R�9�D\�	jY+r昬��q}���<0���mĩ�7�����$v�z�������~���9�/!�40�rZ00��.ʙ1ɣv~u�zb�̔��s��bBR����{�d1��n#YGg�ǵbo��Θ��������Z�mv�y����S���N�V�ZX�'F9�D�����֎�?X��E�����}.ֽ|�=3��r����ByV��ͫ�T}��@[�!���T�<n�D���LKj©C�ft$+eX��W
���QGs�vn"�����,�3_Yp8T�\���rJC6gi��Z�F�s���^^3I�{��c�ĸ��]*���DY��^ԓ�%�zJ��5q�&�le�s��Gm�p�]1y��#����Pn���#C��O\R�K��|�.*���R���{���Όp��b��l��۷�9�b���a%IA���vԵo����f���}M���)tU;B<�Ź5X����S��Z̵}bVG�~��N�Bs���Z���s��
h���9�}ǝ���(�!��R���}2��N��/�����n�����îa�Q*���Kae*��d5���n���c@G��l��h�qͫ��	�;�9�2b���}Ӭ��7q��2�f���=S�G��r��4:��}� ����ʅ֪8��w��@����F�7g���+��S�X�b��~��J�XP�N�Vu������?Y�{�e��˺�o�U��;'��r'���^��Mf�S���=�2!���*�_�;� &s}�3�U�O�N��}�v�-�џ�^��/V�� w|��z��Ev����Ny�kl�Gp�뱗�u����6х9�C�Xv���a�,���s��j� ;�(
����f��V��Rn��	s��:�&�N^�z��ױ#��
M0�����P���9�Ԃc~�u��X��Oaʸ��+��U�#e�K7�jRC:����(ݘ��L-5�A���Xc��@a���D���Ō���{w�L��/��`1��^X�ߵ}�R�Xv{��| P� =�:�:��S����R���{�����+�E�jM
x�vV�n+W�Y��v�l��,���of�|$������Z�^�g�׵��=���+�XcwFJ�·l�hl�BT���[S�gL��{K78���!FA����k���cU<��[�t��Ayp��c۫�,��|d\㡇��ڀ����kق��gZ4����{�;�>�������j/2��]*vr��h�p_g�JS��`o���n��4t:��+	�?��{P�m1�;nv��u0��V��<��vc4�j��}�x�1�7���;uH�0ݲݻ��٘�v�Ɗ:gx�L�+#�$*���#���d�1x��g�{iyzƋ� [�{y�κ�bI��k4��*�W3��2������bӗ���S���zL���t��=W�k*z�ۆ@��ȟ��Q}<ʬ�!Q����_���`�ZY!�j�R,��o���-ۅ�Q���]�H�1�~s#��Q΃�S��TD����ݤ��a\g#J��H��"9��pT[�r-��!\a�"#�1"J��,B���7�}SZ��mI��%��n_[�3#�B�S�d;�÷l�.b`���<O�h�J�/WK�K�WE��!�����y�[��p�rb;Sˉ��4�5Y+;�2Ʃ��`.��(P[]J4�ώ�c����孅�-�"�u�qߍ�3g|�2豝J���u�+1�$T�Bۺ�%N��v7[G[���g��p�)�1N�c��̝�R�]p��U��[�\�pVz�v>�:Y��):#�@�d��B���=]�
�2���zۡ�X��HV$�ߜ����k����XFa�O�%�{��`��߼}R��%�����;�!�F�+��4���D0����Mq�S���nu%L�Ltj�Cq��8 	|$�S,v�A��ݨW�O��g�L�%�l
�i�j�-��{�#��uQ+d�ߓ�cr&p,7&��΢��V�+ر��)�o����S̸�9J�25�j srx�?(o(��I� h�T��i�Т-�qܝW0�uT7y´�#:_T�5LFD��s��u���OVD��8�B n�RDwV�4�vg�S�ASa7�)�t����:k���\��V4=��g
���5t��m��ó��?rˮͺݭ�M@�V�R5kJ�Mj</��ixWJ�HVTv˴η0�]:a�-�Vn�Wئ�+�{K�qO��^R��j�g.O�+<�\9��9��YX�^�>��Nl�i�}J�j���9H�:T���S�Dd�y���n)T� �:�L�yp�;N�K��)�5�=EOg�V��
�X��74C�=Kk�z{� �R��^�Ru��p���<�,���Y.�{�.6�ҩ��RS�4\9FH�Ԁz�/b�G����X�;���j|E�bf�{�`c�Ю�ДM�Q/�t�NZcu]�wc����q���ً&U�8�3��aqЄw�Zv�GN3ǰ+��@m�G��>-�ە��+���ܭ��j�Fه��$�#I���0S(Bߙ�rP�"��B2keN��r�4s���8��h,�\�y,u�����g����N3��w�q�F��]��Ӯ�Z�Y��69"��am�S&&����/`l��!oY\>�L�`��z�#2P����Z������ =Qh�Fꖐ��x*T�����ݸGs2���U�A�غ���w�.�	.iX�f0 ��y`TZ�D(D��rQ_p�-��y�8;��5b7[��A��s33*��H�Xn;6nH�uU�,v,��4�h�~��oݧ�n,M�Qe���'r>E�*��e�F����ȍS������9���6lp�:�C�hŝ�5���P:Hn-����1OAa�]z�α������[q�9=�46��:a�aK��w��{5����\&�$0Fs�C�tU�������*:n�#3�h�׷�wz`t8δ���*�!�[�� ��|b�̅�כ�+n��-�ky�Vu�7[X��s8�xc�<�90�6:��L�K���>a����6 ���G+��&<�:`=��M��M�s���(�eݱ[�vv88����+��	4w�>ʴ�k9�Ͱ�1!�=W�i�&�cj��\꧞C*� /�cC�`1zg�xA<]n��c��7��)y,B�E�E�?z�8>t��8�3�ί��
���7���U(�E׊x�Zn�i��K:>�AnDK�Z(`��G�g˨
Mn*���Y(����7o]ԝٚz���엩Պ����eqȋ�Q��F0[S����%�v@���@'t[f-V=ʽPK�v��㈡&Xw���������=�ӗ���������#o�QJ�b[��l�9O�����,Ǿ��3R"��hQ�y�m!�'Z$\o6��㣴�9f�ǐ�w�8��[���u�x���Ϝ}g����*�p��t���FT.��W�T��'ԁ��#�d�W5�[H�����"��n}�C1Q#�̃.�爔pm^}�Ϫt��<��#]��f��f����E����\9�t5$K.��/�2�T,!��S�rg0�H�0͞�iL�a��n��q��}QϪ�s8���$�Ol	�u 	<!qˉ�B-�!|�7ۏ���V6������jįaҨ��f�m��a�s0c�W�.�A�gh^��<R�&��{�ov�x�MWMco�vP���B�x��mb�k���E�ee�A�RS��m�77�P��Qb�4��V�Kg /U@��I��,V{��o��:su<=Jp� �Û���?:9P>��,���#��2��BJY����K]u�D3���=��Ǝќ�Ů#���чqF��9鴯���;�V/A�oU���R�jA1�ņ�� ��=��X�r4G��˷�6b9�=T���r�+0��k�k� ��a�S%�E�J����j�{Y��cz!��}_Ou�/��=�@�M��F���� 2�|@M��k�����=k�rX�p��Ȧ�\�0�"��Ӓ�]-f�����*��y�s,y��_�){E���P+qP7'�#ծ��1�u�ۜ��]���7JՂ#��'g�����a^��e���v��K�7!�?,��؋��E&7��.?G��p8r��WF4�F6
�7�-ЅE��7�L�/:bB�����T�ݴ�b��W���~�Jsq���n�;�o9�+UJt�ɞ^o T�x��*��ct}>�����c�|b�9cS�bN�*,<I�:����<�h�U^S������TG� � l_O2�6��I�C耝Bl���	��n�����yqJ]3��6]
��.,6��s]e2�fWoP<��u^f�����g���������sĉ�{sw��'���Y^�+���V+Y`�����w5�.�����ѷU�}v��v�^�EwL�MwqJ�]�%,��E}X&7&k|�X=�gI7��Pq�H��@Jh�#��,o�:5���L/sw��_2�ܮU�p��n����!�O਷}r��a�7#��LH�0�/���Y|�:�|�$mt�5i+����l�cDp���V�.E��$��a
0a^B0f���x��Y.��f8`�ҰňB�9܇ŅNb��*�������j�~D}eݒ\�;=]��{k)v�(���牊}1#>�,n�	C(��I�3��PjpH�;bUvu\��z��'8+%�o�:�Ky��<�+�+���wY�9���WK�q�z��ia.� W#2.� �<b�s,v����n�+ͧ��ƈ3�	�s%�Zq.q�;.U�����4��b���x���a�U��I�.�6��������~<�yN�-�s
�W���p�d�,7�o�okt�8L`���TD�!�7�S�&��["�j��(�*��֧�a���ޛ�(��W5��΃��#|�\M�w	�ԁ�q��l���$8����r�.�vV֣Qu؋>E^n�H�9�'��"��=*�w�r���ux^�%+���ǜ�L��2.�/�rj��sX�j�N^ �wD�����ʲt������28��ꝶ��q泸\"�M`l�xzҭ�	�[R�gM� \.Tь�����87AT,F\4kӊյǌ�Ez�K�1b4�L�@�(U��72�-$E�ݮ�9��!����ʭ�O:MĺY��; �q�元=�m7�R0w(��ig�t�F�q.�k�z$�ތ�����Z^��F;5�t���m�����f��<��c�˽\�E�b������-�Ð������x���i�{(Enؼ�ꠊ�����^UHs��䮷�0L��Ҡl@q��f/��A_ǆ�I�F�I��h���;���iegA֝	ۙ����R�n�8%�h�0��FKV��(ƳÓ��I���j"�S	�g2�Fi1Z �B�T����W�=��i6TЊe�M[�v1N�J�޻�y���F�����(zs.�����մtC��B'��b$�Z-]�3v��D=W.�N-vw5q��kS ��<�-[�	�78��e䐶�l�Ҵ��Ѽ�X��{YD�:�۩'�<����1�o�۪!\���f<�U"Mq���+/&�}�p8y�[µ���+)���s77�2qIc�KK�����Jq��c<IW+9p�%�p@�`�Ы��;w�y�\�k�w���hq�Ɏ�wT�z���Vt9Z�y���&b����+%�,�=]�*�ְ�Ϛ�uT�XX@�jY+Q��ӳ{~��o�v��U*xE�+�N��|�}(#3��r�ϯ�S�ƢN��<�����p�:�}��|�B<�L��9��jո���ؑ�f��@O����u���;/�Pڳ�?��<慫Qjd	�\	�TNT!_YzP��p� C���{l@_Ok�������"?]�?C3~�1c���;�9�M��lW?��C*� 1TmHb/T�W�������[�kٝV���L?�͗[3�2ݿI�r88'U���D�j�~7K��Dz�p�$��b���[y�'-+�-�7kNi�\�MW�p�=����X2X�q.�zW
���v�⸏�G�_f����o��2��s* +錸�P�{@R'�z�[�n&�>淵\�K�*"�qb0�F�y��
[82Ξ㌽5*��qpGנ���t�nR��(�ݲ0���B&⎳�6���N�H��o��yk�Wj����ߤ���S֍}M����1�Q\�A��sv�}k:kX,𹏷)*��t��[�k�`�6�ս�]<��^���&
Z�[�M��1�6C�HJ�x˭�]c8�/���Vi�W<Ĩ�|t��N���m�w�J���Ĩ�-�sQW������S�]�]M�/��(�ܗX��>ɱ��%r*"��w�l��ھ�6m�G�.T]������@\�[���h𬙃 仦�ϲ��	jw�Y��+���i+yP�{��B�tW ��D�
��u��$����ٔ�y���岙�W�9j�k#x�������X8��������VGw]No����[�C}L�f�'���|�wƯn�[�}�=n�L撒�2�1p�r�ꕵ�ؒ���Oo08GA��c)6�υ..΍���t��Cu��j��Hq*�=�1ř�0<�l�L��w��+DP�ﻨ�y�S9�+W,F,d]���9��S3{1ɺ�+���q|rX��$
wY�p���޳M>�M�:�؝]Л���Z�0]vF�_b�R)p�6K�����23F^�d)�IY�Ŝ�z7��˕0ݸ�)1�o2�(_S�k�c��D��[�&ᛵw6��Q��т�غ��Z��`�N�җ�0I"̉��p ]+V�G٤T��dz��mR�U��,�]��]�yI�j�G�edz��tY�v��Tg�w�2"ӭ
��znӬNu�ؠ΍�\���\�͒ed�O!WG�r�)Uڭ�5���;ѵ�C��g�)g���њ��Ӗf�u*̩
�9!J����� ���������A�$YG���y���n_�Iϑ���m1��஍v�}֓bkbwF
�'9*����ٛ�@�:�N�s(^CƩ�je���]�^깟.�9n>Yh7�\��T0�
�{3Z���f&t3�{��@D��6�y])�t�U�Ν`�4��J�dX�����ţ��v�%�#H􏮌���.��u��t'�R�I����A�����1N�����:R@�Dw'��*Ý��Ө��϶�t��͵[�����n.��G".��d�pM�zM�>��;��B���'8m���Js�Wy�5��n�짽@�.�.�|�A�;�2����䶳s�B��j�قx�o��󍃥�o,P�;>�}���p��s(�t(Q��P١��	ќfU�_�뫣Va�D�К�:q�D3����� ��/Y�6���ݶf��ﳁ�]����[j�꺛*�Wu��Y���nRk�E3�nd������k�~�A5�R�\��v�we!Mq�u�m��ȹ��١ǅ�sd��v��؏gۈR��qm�j���0�� �J�+;��m�#�S��E��#�Ys�/q�G%`WW��^����Z�kL�Ik��4j�U�Ф<���D���^�J[o�&28*ڕ��{���CY!�E���j��F�i�Y��}k:�7tZmf��;i�w���_dc�v����1�݊Y@�b]�b��*��kb�Щ1�t�*��W:��+(C"��Û7#ɭ�TM�v7n'm�"��T�
�e����εrUٝ4��b�G(�l6vs�^UEy5�s�$g<�Ix��yVU�eibW���Q��q �U<�ɕ6���nMRr�Q5SJ��,��T�Q�)
�+4$P%��b`yU��^�xR�hF��^�"����V�!�����)������[�
��e�S�ëg��f�W��2F(dո��X�u�\h��+J"��R�H�t�s,���"*"�%D�]2�Br)tC�O4D�L�,)��USH�t���*�Ԣ���RK1B��]<It�B��IP�\�D�B<L$2�ԉ�����i�e�b"{0��[F,ۤ՞TcY���7cP�&x�_W�"��p�ɪ�JB�.��s�ΣBv)��90ռ�ntu�[�R���Mۊ�EM<�%�.��]���J��t�u�~Ƴ�q��3��0�_��pN�̤L��DI笴��~@ZC���aҘiي8�!��BФ��q�'��7a��ڇλzVq% ZRg��$���%�y�9�����Ʒ��y�s�C�:���O˔�HS6�_b���0�L��g�n�:��ᄤ<�T�
��:�L9�a�����&Xy�KIHS:�Yhm6Ŵ��<�~��e��ݧ�<���=�WU�_U��P��Y��ɣ���R|�%�I�����S)����`a&�������3'�s(RKz�H��,���V�Rq�+a��1�I�[�N��=�����z�7�9�|Í��q-�\3�>m�=˞��a��-'����q��KC.[�s�',��gWڲa%!L�=��+-%$�b�t�^�̗�5��&P:��3|�5�y}�k�ﾽ���r���8��d��|]E>d�j�q�'öBߓeT���S�2_.f���ΰ�{f}D�L�At�1y�-��In���}]�(����u�����C(Zr�����]�Oew�}���x����U���=�2�R�Mn�U�IHL�bé)�0�i�����U�!���S�J�,���RWy�L��Β4{�&����2�V��)�皘}�6�J�Pʕ��>Jgу�|D��)�}�KB�,8ϒ��(�Ρ�Z%�A���8�j���hZAz��Y�KC?Py0��)-��'P�µ9�a�$���v�Xe�T"DAY{4�Ϯ��[A\��"��[�ON}�2�I-
�5�)�V�r�!wA��凱A�-�ͤ�t��e ��6ۭ�=��fuA��M�I3�z��Z8CGՔ�2S�j������~k�4G�#�"���j�Y�gRJw�\�Ai8�yXy%�m)2{��d���%0�kha-��Փ'�fZ铉n����:����c�2�Y�p�=D�a��^w��WnuUx/�ޟf���ϾV$Ö[��o��M��%2j��L�<����>;��AT8<��CI����
V|��2w�������Kً&��IWT��Ii8�3�����^mqa��Vh-�s��hM�Asd8��q��@���j�^�om�毑u�w��7�J�T����D�h�S�Y��\Q V TrYz�[�q����W�Vg�p<��c]�쳧x2kU�v.:Fm̬*������6���|�U@�f��Ĵb��9u)��J��W�P��c�\$S�<Ʉ�:�Vg�����0y6��)����P�Zq'�oMw���8�C�ݞC)��r�����v�zYש-=1¶��^�7��o{���ƺM�ZJx��@�B��8�uL�-&�A4�C�|�!��l'�d�I���q�q�f�{ra�}M�p��G�֦׹��˾���&Ъ�k-�B���E0��R�"哉l�a3��@�S%3qs�-%!I�e�Ԕ��V�A~O0�����(<��4��Yl�i�d�d߮(a�}�
��ػ�t�D�<�Ϳ��?Up&����~�&�D)$�}��&}F8���I�,���$'�f)H/P��GS�e��Ϊp�3�_h�w�L�aX3�C�4�@�~���zO�^�f���;�}:��z}˔�C�)�|�}�IhR$�þ�He'��k��$���ZM��L:��n�g))����@�����N���
m��0β�G��������x��M� �he���凐�AC3����N�l�OT��)�z���&m
L���Y4�S)5�\2��I:��ن��[��)-��[�h�C ���{�uZ=f��@��^��BU&�lJM�]�6�u����a���h�u2�Y�9x���{����^>JI�)5�Xm��:��o��2k���:�%��+S�ċ0"���1RS;
�9Ś���[��}����8��C?PZK@�g�aN�ͲS�u!��&�f��Ru
t�r�&�0)�I���^�k�a ���̘���6b�h
)8�ﻉ��" �n�]�˚ҹrZ��,��2�B�))=n�\3�qN3f+He ��fj�;D�- ���0ʳ	)���u0��S�|���u
Chf�ef�RN�O{G�1����1���<���+}��w�Nu⾾��u�|�IHe���
AH.��C�i�aM�fsd�C�l8���&R:��Ѽ�|�!i2j��a�[���)�0���e�I6�g����2��S,����7m�E^<�k���an�n���M��M�7ʸԘ[�;]m�7R�GQ���4�3g%nh�MP��}֯q=Jm���`Vg`멕*F�i����xjh\�]�Qk�r[ ��0,����Sox��XR�@�������&���2���%�/w&e2R�픆.��-Xd=�$�ʓ��u�L
C�>m5����Ag]���O}Al��KVO��ZϹ�{��>��z��/��zֽ�o~ �a�-9�6�P>Ja�цa�|��Rj}�O2��$���	�2�_&���)2�RM�KE��3L2͙IhRq�m�������CɇL
C��8��p�ݽ���]�����C���G�fG͒�D�a8�J�D7�Y���A|����!���I]��Yl�������U���2��дOv�]BеCi+>����Jv���s^���~�Os����~礴�B��q�SI�{U�y��[`[�ty�@|��IL�%%!���piR
�g�^0�y0Ì)����>C�l3�����Af���KB��- �z�9��r�>����J�='�#�>"#1#�}��D�m멊��䤚Lj�&]�ZO!N��0¾@�fn�P�
aN�P��P�JC�|�o�����)�����T�e�6g�L$��}�W�j���n�������׳���Aq����%�R�
:�$��s������&��|�- ���^����Ԧi-��oR[���'�JΡ��0�RAw��}�̛�O2[f���a����~�d�>�� �G�}l��,2��Rq�X��X
M!O�����
C���	��3�0ɬT�i��D�ъ�AV%�P|��H/P�t�N�h�,��3��Z��	���ln\ٴ��X�b#�} �W,�N!�-&���P�Vq��e�H|��c���M$���q��*�R}�Xa��X��p��IL�~p�3@[:�II���eS� �؎�
��тǎ��]��h�1>L0�������<���Fys��i �ɺ���N�h���O2��>B��!m0�pϵ�ɤ%$��a�����ɭݘe2R�@�7Pb"��G�B��.i8S�|���UJ���x�C䔇��öJE��ڬ$�ꇘZ��i:�r�%��o�
C����I:�KH;�q)'\��-6W�+&Ҙc>������^�`�p��:���>�Y�c^�|S����ہ�7;��;��	Ki|���9Z�dK����_;�V:�f���v�y�f�����f����	�e淊�]��;E�}��姪I]���F�����Gc�hֽ�^e��K靝
ū��t����r �3�!#Ykkg�~�y�~�f���P�O�JͦLPa&�]��d��:���I��,�i�tn���B��9��J�R[9}�x�䷬
M��L<d�ц=������=�6������g�v=�9��RAVE�2O4�$��TE�:�B�d��[��u53FS�Z�\��)<���S%=C�-Y��U�u)���.�BO��z�X��ٗ_�𚡙:��	U�)�z���"��1uՖ���<'���w�p���x93ZqnksPq����#j�_�;� �<Р�J�3A���l��X�~v�9ٜ�k��1�xc>�5ak��Z��6��8�DXX@�jY+h��E1o2z�:���ɿmׇZ���ު�|��
O����]g*4�3�P��N�E[Tl�h���� �1ʣ�q��+�ꂶ�nQ���C��a��B1�c-뼐�W�T��T�8<��M��6�|��CWv�k���C�Ev�����n� �𰬺�@W�*���[���C��y�1��O�ݽ��S��c̿��]����&���}-W:�y���X���[�E[��k������Ӽ���Zqg;��<�1�
��eZ�1Z�~�\O��x/y��=���4���rxA�gm�=��N����VkN��R�,ń���0���m�����Co�G@�K�T�W��t�G��F
̘�[���gz[K'��v��v��U���c�0$��Ef�����ǈM��5�Pu�W$��!�t�]�b�`ٍ�'\1�/�L��z��2��*ޖ!�����5(h�}�x�Wk��r�o�ծP��g��b��΂U۳���~���j�
���L�v��

�c5Lw�{@R3є�d�L~�i2_����@W�:���%����t�pg9�9�5);�s[Rr�v�mݾ��&�S��8�]?R��:��H����	��޺��<M���~���1�^���Q��ŚTz�ɗX8��՟��'hu�m|��K�+k��b�vNŷ��0Ru�/5���E��@����/�(�nY���1U�i��ã��f��9�:>�y�)n�?Pp�
���a3P����@�2�
����P�0X��#jᬺ3s���}ҭsR̥����8�� ;;ɚ���b��"�⭠:�Ol=n����8Ža���b�;����r��!�����ǔ���V�X0�*ss�͚�Sp�����$>�/�rn{�l���>��W�&�r�*0:��6L!�����(\@R�]�`����쬻���g^�M-�b\{[n��l��\���*w>�U�=�<2�cyݏTlp�0��C3[F���#�6Sqe�7�MR�h厡�']Ҏ[�_klZ��ˡO�zI<�ˣ]����d���sֻ��JY�J�:*�Y;�������J>މ�]o��궈�~�b���p��&���F�d��Z�A��� 1�L1	\����CR[�z�5T��C�t��0E������͝8qWC�~��jó�8��G�=�ȫ-�f��;w~�7��}0��]@�Qۙ܁�����.�ق��Y֖=�Eo��.�5xd��H����f���2�U�Qg��z�_�+��&Έ�<�:2''�P�=�i<��2C�6�3P��c�T�/�h���l�2�Ћé⿟d�&�Qs/v��	<�{�[�j
���E��fC"�q�&_�%QBj7i���Դs"��;���d�Jd�^�Ii܃ݭ�������eU����5�@sʸ8�g�֞��| �X��ݙX��nN�]���G.1�xaWZ80p)��n���MV�_uK�����ǝ�c�A�ɓ�Ď{�BS��1Ɣ����C�a�'�O.�7'��@]4J#�e#��M�Nr=V�c�R��Mk��L՞��)u�S$F����V�\�n�W��a��s�=bqJS)�f�y���9�C�e�8��s2�D-�W�u�	�Se�i�V�!ݤ+N��9:����c�����L�z��Sʿ��1n�}w6�6\]��'ֲ�<̘#��Z��������ڧv�F�Z��JP.�M@f9�hhO�J�$����˔Xg'8��!���2S5i+��:[7�UQ����+��ݹ Y{\>�;b�bN���1Na���!Y��u��V�3�p�S������Y���ڡ1:�a��$�Z9�D�}�Y1+�$v)cv6P�1"��[;�a����U.�9
iP��h�x��Wg��e6��mG]��a��,E��f�=��zF��R��Ku�=�H\¾����k8Na�'�T9�;p͇��v�f��}l^��L�����v[�ֲcAq�Ʒ�!��K"�a
���zP�gL��J�\J�)������Y[�s/�㺫Mƞ�o�Et���Mk dstQ�Ә~���8n�L`t$��2s*�%���0�z�\�LV8���_!�SO���T�k��h;�^{�)5���י���z��bD�^���<�7p�蝞Mxe_ /�4=��p�ӹ�Mk�t�LSǾ���3=��6Ϯ*�B8Q�J�q���*�CY��%|eZ^ұ!V���у;6�[�]Y��:��V�1ĥ;��n.6Ň�1��Nu�5ѓ��V#�P-���ڕ�V��^�T'�c�Gۈ\�VX��Π�����q
Ě��Q`zi��6�eXŜU�3Y���ǫ��K��B7*.�ךtTQ��ف𐨳�}�]�x���z�@�ʖ�ox��s�kޗ�������r��G�uҨ��|��\y�ە�Y�m���n����p�W�Qxo�s��dS~%.��'$^}�0B��>�� i����+N�"�{�`����u^��"�H|u>�h'M����7�P�.���٤VDi�!�� D̺�N�r��7�T���H@��A�P��H�N�1�:[60F
}0�(�a�xt��U=��v�8��Ԥ��x�ʈ��1�:�F���:�W��t/��⦦w�v�G;e^��7���4�[�u^�(������<�ER&(hv@\b�A�v+�,N��F�@R��t�{_HHC�Aw
�
�fD��,�B�y�@v</�k�g�k�2��/k�p٘�-t=������1q�Ϫ��.���1��O,	��3v\�ߊ�|�0��15�{ޝ�H�=�
����0LoD��N͞�j�l��6"��@^�s=t��o2�K�6V�Py����m}�s��FJ�d�A�,���T�f6���0{ۮ�^X4d	$qQ���Q��:-q�ڱÜ��s�=K�����H����޸+v��v�,e���܎�|kgT�8"��j&]�|�����n.��i>,)�(k`�T'Ws9Ӗ
w�j�7�a��	h��駡��5X6��s�!�Q�8���Q��꯫�J�3�?z�D(�#�k���!�c��"�Kk��@W����;QԹ��3�� D��-�:�;���v�Z��L8�p�V�6���P�	B²��^��Y���X=Xx��A]Z����}5�@}գ��׷�pV�Oi�Rp�]7�
������gÀ�,����Y������C<�@
��:��Z"~\�h����x�b�(ΏZU\[�Њ0�z��emٞX�iq���!�\��0�fK�i9CE��<n!l�b����)�:UW'�9�J7��.�'��d}4P�n3��\��q�Բ�F��7L]Bn�2�Fe�v��31x�m�Hh	������t
:Ȣ��L7�_�4�ls#�i�N_a��|s�^grٟ��l���S�gd٘y�L �g�oZV�Ds}_n�b�3���Km�Q�8-iNT���1������v�ܦ��-��*�֏I���z����8���YNo�8�U��r�	0y�A׼�eu�}�ԧ��G|�dc�J�i-�] �*�lO�k��׷���Зq�k�&��_p]��Z����vuq_勬@bn��;�Իm�F�5�`��F����:�}ȿljZ��	ZaH�e)�� ����.�Y#�݈/2�����8������9Wnv�B���U`l~��>����[������~��$�'&a�P�V��	�p���R*t\�jC(ED1�;�����Ӊq�>�=�g���Q�*�86��'_S}L\9�����=��yP@�K8���-��r����ҝ�1=�wČ�~�)�����aTbV��3��_*��H�%Ѳ�+�Ⱦ�Q�;�T���ҭ>M׮W���8�1*<��(\!�f�9����4;���M�����!�l���vY4�:�Z<Oו7fxv5N�'�B�b��qK�F�O/;0p��gH��8���HR�v����t�$t�|��Y�~_/�R��^ҡ���臩������T޻��5�*;�C\�áۙ�*��+�2Ga��%Ѣ��[��{�Z��ڪ�"��P/3z��,[;�	������~[N��ܴ[c�N׸-��i�{w�8�_��.i�C���Q}�u1�0�n�@����B;�y_e�]EE���t=��Vl����nnl��s0�3��L�+��e��j_���ة;��t ���z����������,oܽ�^��QC��A�o+U�x`4c��l��A�� ��S���25�{��*�}7<��s�Ca5x�{�8�;k��vC��t�D��])Űh>�V�� ���w<{��
��+H��p��5KyVY� �p&�k֭��h�B�+�r�U�v���D-�����Ԍ��WD���r��1��BBS=�0o^�Mؗ{$�m�,V*@�À�)�Up�/�t�xtQ�����(S��H���²�pv�^�l��g�х�1Z���9W��e���x����t=[b��Ǫ�����6: ˺�wE/���{o]�9&�vv[����rb�̵%[��Wm8�w%��mov��6�U龡�$�*s6�v���1�7�*P���e�u�x�N]���-��ХL�;u��԰�
v����5�e��*8���(��P�O�t�G�h���5� �Fj�����k� �Bps�}=8���w�1��,�|{,aJ�AjtQ�'hPc�Ij��C���X�2�֋+&�!yJ`���G����ŭ7Y�m>�j=�^tZ�[�;R���c�S�����b_2��������8t���ݧ��g�	;�F2{���X\*v4,,�VQ�1�{�y�/�mB9�5�ƻ+r�˜��T��*�v����o[ͫ�:�Pވk1lT4:2�}��.S]+�N3}��{�E�AgU�����`����&�4��\�W�wNVG\��>غ��C{��� 9��nc�0����:���>�xK��<xuV���;7L��7o6�d"5���{bj�׫���~YW�R��3��L�
K���1�xS���u ��/e���n�3��O�#^�hCvE�2��u�&us�R�C�Y0nӕe�Esp��"I�{�x0Ջ¨�:k����e�� ���������7�Ӳ.�ל��R��\ߴ��^�B��Dr�.�R�s�N��)�᜾�u�X2X-ռH�Xb�+u�Ղ�"�k�뤈k���4˄ͫ�4+6NE#�	��N�����y�\��9�6�W+���O�Zu�V^J���°W��E�&�"�&���p��
�l�Dt[Fv�����܋ޱ���DaCdN���gKb8lҠ��dgjT�9`�9�;���OB�)�]���s�B��o�ov��R��X���$e��Wk+w�)�ͷ�p�"��*��3���]R��w�+�/�Γ#�,-���f<>ΫT�n
�y}���Eoo�Y�.���0�K���iJ4�t�5��h�r�3�c��������O>��4$����p-�UԂ�,��P�MmɀRa��n�kT�N�2��(j����P���و;��zuŷ�nN�<����[�����ѧy*�-�&�]��uc��#'�盰��мC��$.T�A�i�hB.U���
֥�;�+��s�9�߁�4E\��E"2�/,���KM��ۡa�*�QY+��E�j	QF���]	�a�ᵇI�S�r�"(�����E�����Z$&���aW�I�i2J�0j�O47$팫
�m��R��t/RC�$�v�m�4W;\�����YYe��MlM���/=(Q
�1F�QLU#���ffzk��➊�N�Y�b��
�fET�k��H��,�0��"���B+3R��I���&�&(�����J�$�F�nL�&�Y��i��X�bA�e����$ضvS��	b��F�g�k&&����izY*�n�5t�M�	�P��R<��B���uЭ��z��l�4 �W<�ۖ"�jP`��Q$D���������e*E�!dDhE�6�F��b%�.YU᫳�2��r�*+�Y�M�]ED��O"U]B�ȃ���*24#1E]�v�ujq�Gp�QT��\��p�J'2���H�4�7$@�BڲB)4sL�K!J8��"h����b$d��W�J�>�m���_G׷�Hi��b}juK�XU��䊕���;�ۍ��h��췳��0GC/�k�j��h�6u�TT���������T���cۄk�`,R5ёmr��{B�M�|�xө�\!5��O|xw��5ɦn޻V^�uy�o+�]��8j+�?�A�J�Є1��
5�1u�O� �OuQny�'�>ɡ�Q)h���f��U􇫕���B��(v��	�Ckc�O��:' �����=�h5��D���hӜ^��$lp�$븶�L�̬zc~O*�G�ۂ��q����2s��~ܬ��𭫩o�E3�i+��3��NcDpL�+��\�3M-ZH���S8uM�3Q�Vm*��wK�����/�'l�@����!�?#rɽ��r�'wZ:E+���kb�qԖV���]��/�S^&�b�.�=;�\�B|{�b��;j�8��}�V�ܯ��������3AI{Nj���Z>�rNE�!�<ۍvs��L�Wu���(C��'Wch�I��@z�#����W&�BN�;�Y�o�S]#7�*]9R		�[�ۡ��`��X����&�L³S2yF+h��ǃ�W��3�&�})q�;SU�r�qj��Ӏ�N�k'i[��ϐ����	�دJި��b�u��r�;�Չ&T���wcf�Z�^�t��{�9�wh�*�����n�W*q�g�N���N ����5��B�IΜ�5��J]����,6���ϔh]�a{'kf�ҙ#DE��N��SX� t�S��<��r��sO.VU'o/�a�D�0��TNT][���X�8��=P�"{�۝S�FFt��ny��-V�w	0���o�RDf�Mh�'f�O*� N�Ƈ�U��@D�U}�zg��`8�䦞Ǆt�滊��8m�3Ƙ�D�o�|]gC��q�B=��a�5Ї]fnᬶ��E8�W��s1S�چ���m���R���o����b�Ԧ1M�a2����=g��Z_L��rR��5K�')�Lh���#���@�Pg@ޚ�we�O	ݷ,��9�X������IX�a��j�\<�'LX�7���Ӧ8�ck�k�U��U�8�6�S�/@��9 ,�#�� Q��E�Q��:���?�*BP�P�T������9�&���O��1R�4T�ID�qk��W�8��
���Y���X���� �³��Dj�:̈��&7�f%� pY�HD����j��ʾޕ��c֧|!�����v�J�e˫*,�x����U��g����Y��ny���KGQn��g�wޅ�f6�s�^��L[��σfE���\k+���D)�޾;�*�
�Y]#Z/���E���{���D�a�%*��+Q��ӫ�^5o�ꪯ�"L�b�r�-���u�/��@��Xx�$m��B�ܙi�dR�{�tT��cZI�2qT�_���u�8k�U��9�#��1�����X�D���ߨg�̯���`n��~�9qp_t�' ����UC�HJ��� /�W�8��s��;�5�껂�x1Q|��\]�;^Ru���Wt?���]�S8ew���#N>�Wr��U��đb�����5(�ᒍ]� ���S��l����ݪ�����J�{<���1�mX���hp�_M�!Qe��p�
�u�:� �8حi����4}���Օ���V�!�ca=�\�f�/�T��y�"](�h[�3=]�B�v��Ӎ��o�
)�x����yR��^|��Z80���h��P�8X�:걪O�k�m|���*��]����n�i�P�P�(�Z@A��,J��婣���7�`�`�U�ZUrd}?Q��n3��\��7)���s(m�Rr�x�Vj43<���v�Xk���]�OiM�7p]�@��ʀ�T���OM!����l
�.�P���*������e�������R��7Ls��ԟ�������k�Ee4([0�M����U���Ntʉ���7������ﾯ��x�޼�a�B)��GE[����Hq{O
��ץV>�+3a�\�"�`)Ft۹ZE+.b,F��R��f�@sں�
_>��G��I8�{�s�� ��餾p�Oi܅0L'o!���_U���|N�츪���(la���U��Ͷ��jfq��"�[��|�+�X~z���+�+鸣���Ʒ5���̮Y=��g��sB�0����v�+��x�ŀ��zV�u붃�"�Pe�M����1�'�˳��E��vy���@Vw���#[W2m��ԁ�<��xr�{7��.�5G��Π�0�G���B�����x�|
G�T�;1i�ψ��,:��8���������v���iV�����V��C��
�4����q8�����`��m;ݥ9ALU���n~ɥ�A�"���-���b����#�Ȯjr�F���ǳ��W�v�5̔G;I�P���_S�'�۪<vR�]f_��{�8k���Z��ױ��&�fc�5�u���v���e=���Yǝ3B�N�33��BE3�e���:v2���ݯ�Gz>oyة��j�V,����k�C�f�bt��EW����|=7��zz��9����+u��N҃�56s�gR������ꈞ����=!�?B+���� +�H��:�ƺ���j�R-�Ѣ��%̑�^����9�Yˈ�ӵ��k5���hߐ�>�U��ݲ=g����/_�5�خ��5��<�_�gg>8t��/�����q;>��yT� D���l�@�)L�9���.2�������s�мz�Z<�+�Æ���˘a'�^��bD��l��͞�Y[��!�S��ad�������{!>�U��xq:o@Mg�9�\J��㊈�%1g�ז˖�����/�RF2!���<�p)�nD�&!�ϥX��n�p�P��tĞ�i~�\�֧�&#Sۇ	� ��C��F����(����'���B*V�f;+���<y�p�:��l�ϣj5g�ғ��'$G#C|kE�*���(�9o}j��J�܇�7vغ���չYy@=1P#��w�I���B�l�ba9�ü�X�3F��լ��c>�}&�v�i5��U��5�V�o�xX��4�h��w��Ω[��=S����%�\/�8%+�V�n���ڇ]��\��Qp}y��K��v��K�K���ܝ#�n�q�$Pg|�i�&Y�9�@m:#��!����K`n!F�4����[�zW3M�r��>��i�����D�>��%�x�X���~����*�W��~N����U�}r����-��v����5*�c�_/�
�`�>�ޚV:N�Uw^K"�Pz�\�]!��,�w�Ծ�O����5G]����_�^P8<鹃��L��&�z��W��TTiBMHyMP�p�Dq��2�n�������4uXz��Ts��
�L`�70٨���CT�3p�1*�(���1z�M�T��-��wy(�t���ǰWZ3Ʊ��Tǯ�kB��y	Mk srx�ӂ �N��A����$��tn����J�^"MX�D�n�,Gm����s��Z����x�>
��@v�=h�����R嘻ɉ�f���yvg戫��D�ө�^�����Z�����ZkI�dWVd�����O+��5�Q���D��IV��·Q+�[�����v}�����	�U˅�m��T�/j3S��d����. ��ÍA��@�3�1�G-�&Q���n-����9�1���9H�dE:cE�+:�I��J(2��sj�߬!yt:��r�����},u�K0-���j�J���j��z\�e���x���]���l;&�v���ۢ%�$B_K?L�>҅��/b�9Hm�]�b=�.�[H�gp��|Jԧv��$ܡ�N�t���_dj������D�(����u��>���51�/T�|bG3Q����2��c�C��̡.�0��]��6�c�q�$�ꖀ��nShs�s�A�U�4�Py�Q	;H�|�T��q�U;j�^��hF���6�G)IC6bR !�2�����6yW��U���'�_�h={~�Nd�<��'ْ�	g��;=������O�ޯ��0t5uJ���p��1yT4�����-�f�a�Wv�9j���ph=iހ��ā�(DL5!�ܙ�my���w��M��y����*ˁ�E}�K�ճ�9�b
S \�vy�A�\3DP��⫛k���s��}���!W֫d�iz_&,N�	'F�} >-��P�1)|���j�7}@Λ��tg9~���Ƌw�󫗦k%35�Q|�g�@f6袏m�@��ect��CW!��$�H��|b�Kf3
����k::[�y�ʽv��O#d���=�_��:���S}�=���ف
�m[�a��e���1=��L�zz�C�О>o���U���z��:��u��������c0�2��|�@�^���n/&*6�v�}F��ǂ����.�j⽬9�ڍ��� �Oz�]��|���"��3�+i�.��c)g;�钖S�3Rug,�{���#�u*�W�9�w�.^)S�����$���V+-���E"}:�q�1}=��=����7^h��K�8lW;�j�)4�]�s;�j���@u����]C�3�:��tHOtWԖ
Ѥس���	�Ӯ��sm�eWg,����������^|��&��1ۓ���P����9�M��8�,J�]�R���D�԰��6~b���U���;:ܦW�ser��}����--'�qZ��Þ�`>3�Qh����!���t7���ce3�)ժűz����bS�rp#���J�p%⯯�a��[;GP�p�p3�;׏�wS�t����淳rJ{��:�����q�`Yϓ�p�}ӡ_ׇ�A=e�Hb�*D���5
0.<H�YSe��^�_t5�����W�N��|��zH���̽����&2�Wӎ]9��^dgϦF���:�� 6r�~aEb�q7���nn��:��wR(t��c��ΛO�����7<!�`��P��K�g >9�erj��s�[��.NC��sE[���Tf��4X�+�ƨ�5
�&n�z�2H�*��R�#eb�į�;�[��B�BYO%��p�	^�xl8�W��R���N'՘޳��J�������/�kOo�sgoN�9'3��C�ۍ�R��a�sW�I �ow�Nﵷ?n��?`V�Dw���"�#���/N�B��
���fP��D��3����>�/�g����O����G�x���Z2|���n�+,l���+K�3�_RJ.��H].��t��$���銎j�0���> ���Ƨ�ȹ�0�&�k��p�Di����v&Ō��b��d_Ţ������?��ȏ<�ӓ厺ͧ����k���C��/+v�w�+3���f�b�J�������2+����^+�%v�;��{uTkI}�lY��cδik5�,uLU/c�����wSƙ���
���v�_�&�nI����B�N�g˕�pl�z~U���w������.���7bIɋP�3�x�v.|\�/��w���h�c$nnl��:�Lpu�6O��j�1�Tg4<�}Kr�,��G纍$t0������
?lC�ӳ�T���u�.2f�wN��Ea����z�o��)}3��֨Ic�T���,m�����c�=*$�m��PXli���6*��>��������^ΩV�xcj�H�3��S�k8���"3�Ӫ�f����:�=�F���/f&z��k�3S�s���>W2/!�^g�G�f�T/�zV����d�ɜ!]t%�.�E��y{��ө8�����o�IYn���e"�5]���>�q�c�|�K�+#��چ.�E\A .�5Z6w���>��绠i�'쟊�����ݘH���~��'I������Nt���Vz���p�;�^��9B׾C.��Bxdj�}���p�-{K�;�Ҕ��L��T��;�F�����%9����\x��r)b�rX�!+�W4��#�!G뮿gӡ��Iϭ*���S�ʤ_k�qd��:\�s��\MDZ�r@=#��MK&&)mD�����̫�y�k�)e�٫��ȦR?p����{T����Ҩ����2�~ӗJ:[���5���=�7)���{�R_�pC���+��!������|��k X�1�E��e�ڼJcv�R+����PG���{���i=��]���qe��ʨ�q� #C&@��F|y�s��'ku�n-O�Q�2e��&ڼ��v�t!�3�#���<�5�����G������k���`��޾��À�W�jǀ%�|.Z����i��*���dl��RN_��vʽBD=��VT5���k f-�vQ���]'B��i���䴜�k�Tm���6��s��T�E(�۷�^KH.�;�-Rfj�bh�y��Ĝ�܇^��	d<�U���]wS Wn�Ҋ����#��=��oW7�ɭ����]�'�{�8�:�P�ots&X�<p���ʥCMZq�yN�֞�֓|�9V�#��=ZQܧְ0n���R��0_],�"e��Ĕ���]��,#��+8��	9j�NL�A��eؠ��D"2e�x��S�]ۖ��ZӮ�~����d*���ԪS��ggu����..��R��������u�ܒ��C3uuk�M"��ɩK�����Ѽ��m)�����'�:������n�U�4��V���Mz!��6^��]�#�H�Z޳t(Bz:D^�d}��u��L?J�ۼ\��+@�2�i��sYƣ.����s�Q�r��1��;®�]�v�TU���(ڭ6���V�#0�&yYWg�=�2�S��h	B�є�%-�'UY�7r7�;�Ƶ�wͽt�6��v'����;8\�Ӎ��yQ@N�i�ޢ"o�泹�<����٣o@ʶ�T�E�
y�v`�M��S8��FV����p���,wuW+�j0yl�&��|�^: ���\b�	r�Xh���C!wz��(sW�-�{��.1�
hn�^�ZV�m�.;��̩�f#�	�R�Ȯ][�6���H�tg:ɃR�#��%�]oc�Ի���8F�h��-�)b�&��ƍ�[.8�)��՗�ؑ
e.�Xol�0�A�����'�*�U���1v �v�؝�OI��c.6z�j�3�[�(H�B���y�o�:⩻�+m|^�싫�����В�
��5�9�>̛���E�^�I_�����W�9��V����cP�r����y(��h��Ϟ��8~)T걵�+M�И�uVĮyN ��� �SV�6�4�k���!c�����h`�7v�Uλ�0�����A�++��j㈸�w"���H#�0���#]��v�Y���1��o�n��\�h���:R���i2��9`�-n��E�-;���h��4h��H TgL��gji`v�q���uChS���w-wY�-+��0|> $Cw�,32E��l,PB�uى�p-ҭ�Wu0��#9�}: ���C�efR+`Ļ���Q�*��7::�� �Ɠ�B���z�V��:��W�0�5]�]�"�6�1�;o��v]��+Kf['j6�y<�-���C\@>�L���Od���,\y-/\2�a��3Zz]q�Ԕ�to�H]� ���kx����w��<�r~�m��9$G��G�%����dD�����0�n�U����%Re%ѵMD��0��<�(4rAB$=�����b�b'�E��J"'� Ԡ�%�DV�:gbPWt�!=*��H=*�,B��ST3I�!��+Eۥ���Dzz2eʠͩ��3g���Tnh�z*"F&EnfI�F���E`��f{M�j�e�J�f���jV,�����^Z����F�螆�����Dz�yy�RI�[l�jjE�)J��I��Ah�fD�F�ѳ4��s"J���L��<��M6w8��yE���<��&I�z�&*ʛ�4��d�e�b�i��zs۞1W6vE�J��"�I��!EnE�KΡ�hICY9�5R"��\��7Sҭ
�\�t�V�1L�R=�fB�5:#Sْ���V��V�hiy�6�tʢ�!SR�#�Y��W-J*�֍�XZ)��l��!^%��$��Pg��(�I��F@:�I�z����dÖbYb�Dñ�l#&w>D�vo+踛��K�����s/b���t6��gml�ui��磌꠵�.�鸖��c�v��o�*��V����e�c�я+��N�	W�L?����;����:w��o0�z�����6P�����v�ƥP���F��t�o�����dFtP�Y�T65mH�o�/�u�̈��I���P��E:��e}�a�������u.S�X^w�}۽'�}h�xj;=U��^�}-�숩a��U閪t�u<c�����3�2k��s�2��d���LWTD��V������	�ӃDp�7�r�Y���]:��5΍�Z-��=�@�dɒR�����tΉ�j�$bb���.�/q�5�Ghٵ�p�)_��l}��}��� FTLȒu�D#U�5�*�)����GwE�٩��م��x�P�O�Ce��KF�����������]�'S\�*l�?�J
����],E784�� �.���"[�|V} =2��E��,8��U�.�8\8���8L!�ba��i�����s��b���_Z�r A�qNM^@u�z�L�⼊|=�dX��L��. 2v*dJ�LWXT5T5�k��ͼ*�_�9���:��c��Ok���t��m(mP��C�Jhy�]���ǈEC*�U����N@�F�ի��-�}�ɭ�s�-�-k{rܙ�h5:���l\�l��%��������R������3�������M}�i|r	��@B���ٷ�f��f���/5�#�1�1�!+�_ ��]D��+�`a�r�������
N����b���0��*����v�g(sj0�oUhYmc��s�R�ŝ�4FY[8��\�3Q��XӼ�q��ThK�2�ݹu��V�������͵45��t�,�n��&�����˄3�Y��p��ųz����x	��q���3����"��X.�]�"I÷���*k:&\U�PY�G��j�R�pm0^� p����~�*Uw��BU�_.�g.��Ņ��	Q���=��r�;=���=�Q��:���1���'�7:X��Q	� ��F7�=������sֆ��oE���`��^�wU����5��+w�Y��2��i�6N�ckj�v.n�E����9��l�T{��;�?S��u��}՛�ͽWѿ#�2R�U��oj
�W�m�uy�R����J#�wq�>/�^|r�vv�:zB��Zi��qtI�(�ެ��ugm�
��ݝ7ݳ�}�{S�����:Ѩ����$�X�u�i>]ܳ�`��X�6����i�5k�v�d�Z1��:���s����t;g�D� ��iOG)�h�ѻq];���vL�HAխ�ܹ�ԙ�kV�U�������}_R\��Q�OUO���\s��n��z2S���a*�	P�YR\+��N{Tn�o�\��b��ݜ��LR�4��&;Rz2b�"�ev��}��.�zw�$�2y�,듍t:�9��j!N�����yG�E-h�����e�L]���']��+�>�c���^���8秏�o�x)�|:�:g���{|a+�u�mb
Bz27����y*�q�t�+NPIGt�N�W״�������NC�pֳ�~�}��U�*��9]q�1=�^o#[���[���
y�n\)�v-�N_m���y�:����)��wkjn�����$�S�C��ڈO)��`�|]9�L���Emي�$=�����K^NTbzkT��o9N8���v�G���ؓ$E[ ��ǧ��� Zy!`�Y�\�W��+�Q��gVl���o＋W�틬e����k6����'ކ�p����D��1֟�qu Z��go�,��ó���ؿ\&S;ۙW+�\����HEҬ{���Z�c[};��p[��Ǻ5�o�Y4�:�:�� u�J��'`}��:�-G��G�OJp�k�٣����[g�e�q�8�~!{j�R�c�K}�3��Jey�ogWOZ��gn��y��째6�f��ڔ����[�Y|�nT����EGy&�<��E��ž����[�S|u�7���lJ�5�j"TN�>�N�)��z[��Z��و�]P7�4���&*յ�ՓGT@y����
�}׋�ol���C�7���qַ�>����;��'�n<�_Av��p$�X�A�N���ǥEԪg���B�ޖ{�O7�1~o�Ժu�U�ۣ�ha|��msh�\����Zޞ����t�4�3���c�7��#��������C��/}�4��j�B��p2����F���\P����I�
>Y�Rɽ�A\Cp����Lz�,���+rq�S˦$k�]���������r/a��2������&)[<.&_h�i�'(�;�*S�j�#V�5�0GYv�<�>�S�����Y�(��֗	��\���N�ZSD`D�!T~9�9'a�����iYHvh���5�=M#I�R_tI�5} �I0ooe�̔���A��\�Ǣ$�ŷ;2v��fC���[3vs��j,课��u�dw�l���iTk�R�������jV�%k��\����k^LGuZ���MCY�ɥ��(�O�Ǫ�|��L���������]�c�q<޻Z�}�@��9m��[�4��۪Ύ�]�!8��,�O����^c�������M֩��n� �]NA�Yα�v)ա����7��P��r;*ϭꢱj�^ڧ���=�)s�����9�{;P5��Ij������m{���zc�9Tqv�=+�z�
��B�c*v���=��!����z��v�ϴu|��T4�x���	1\S�S�ؚ{C�}��t�n{Zw�4�˼ֱm��ֶ%O2]���aN�5���W���I:�<���z�F�{�k������v���3�\�U�Y�'�&�s��G���;ѱO����5�q�_=�ز�d�6o�l��f�sx���1���.�ڕ
������I�Tc��HdN�ui[tw����-��Go�L(�QKOwPg�iq�
e��|�T��L�] Z�x��S�@�*�*D���4�a����ڈ��ze˳��[/�4PoS�T9���k�&����6A��/��着�2l���%��^��iq���|9�b!в�ƽY���p�1Ԛ�k��ܾQ����e4��K��<Я�f)�0���TՂ�x^f{u��Q�����ֹ"���iN�3�:�=�P��)F*���a�������4�[�a�ve�̸
�3y�m�4�f��u|�@�y��//tY��qЯ՘�?�~=~͈ebǷ\��A$��jU��ɵ�6�����J�UZ5�\.�:27���~��c��m2z��ut���{�*�6������)��X@U����y�����k�x|mU��lrٌ��z�(��I���c�6����"ީ@N�"O�8�#�v0Ӽ��Xsa�S��x�(��P�����p�^-���t[��/ݭn	�|����R���,����o��ɿ;��V�'MKѽ��mޘ[���0Y�A��T�߄%e�� �ɓ,�Ӿ���S�]�lU�.d�))V�[%�z�«�:c�*���]�Y�A(�Y�~�ҦrNN9[�����]͋���[��eԜ�dު{�Ů��K0�y��z���9J�ݲҠ�l���W�U_g:^�Y���t*�zZ��,�����{��Q|�Jkk��˲^�JsC����&���w�Cr%A��j�����W�W�}史e�c �����Z8�V�6��E���BwIP�'z'�|����b���Շ0��,���/[����E^���:���nW��eJ�)E7;X��:&�dO*֫roS����'��E�Cз^��黎8�0����+�,�ԧ�f/.Nx5/O��WLސmvzN�͍ܨ�(�鞫�Q�>��؜��^�����d̾�5����ސof�C9���ƨ��Z�5�H(uY��p����]+�:�+e�?W�>/�|��rʾ���m��-*kV���b�|yoY���}+�j1=ۀ�迵��7P���7*��ʬ�.��AC�n��{����/nJ����~��ez�=� y�	��y���J�*k�m��ߵ�6oP�<�|�n3��i�w��v:b$+�"���z��}g�C�������l=���2��H6r��G#r�xk]���gn�aB���i�z�qQ�2��㝱�T�Wﾯ�����F"�ٛs�ܟ���p�r�Cw
g�X�6�X^�i�]����scR ����[Z����w��1���yN�|���7��r���KZ�biRCk����)�b��0���7�5�ڽ^����nC�"A���]SK�ِ�׀vW��vn�+��O+w�~y�joR�{��ɑ�j���V[Xj\�ۻE���X7Yc�8��Q�T��kMN�rP�w�Osz��zf����r5[<�/�\߹+�4	����7���dk�9I=��RZծ�Ηv?�9���}�[�S|tw^�n��\�����1M
�bw�!��C�ؐRǅW��Uw�2{�����]-�GJ�W�+n�Uj*��m���c�q�{�r3\������\d��MR��J�p�)�mi�����ݚ�b��v��
sj�T[X;t�=�Et���$�|;Ui���2I� \
���R�^Рۃ�D�aZ�z%J쑜�F�9IR������l4�W��i@��ǆV��N�d�]Ef�����[�@-��ܯst�r���K�Dcg�򸞁	YV�@8�օO�É(o5��dT�����ﾪ��_{}�ŚV�����+�n�-əsК��'��x�k=���ZY���O��y{�e�Z��٘��⭘j�B���k��.�HGn�m�nDͮ�К���OS�s�'�����a�]��LRcrk��t�v�e���o�~��[mQ�z���s����*Yѓ-m��ޮs��Z��<'�JѼ��
k��c�5�cz����mw��f/��ڒ5]?�������G۞�#ym�J�ʪ\�#�r#Ơ>ߩOz�Z�]l��{|�T�O�*|n����3�=�/1�ד��/�/�����w���y�C+�C��ë�yF�o-o��[츶��|�QX��R�bN�(<� �f(��&yez�G�����QvW?(3g'{�DP�8��0�,��p�}��s�rQ�|�Z_����~�ryFk��߹+�A6��m5�q���.����k���G�\����k̊�BZr;g�v����wgqڤx_<�6�����jeh�E�qt����� Y̥��0�V�Kx�T��PJm�Y�
X��mۥ�Sݎ�l��5;�dQ���v)��o���Ыc�T�帨���C���ꪪ;	}���'�6�{�QΣM�kN�Ykr#^�D4���h�qJG�:3�M�m�)w\T�5c�vjV9m��Q\5<��]�޹�+��x��ϗ���|�I·0�-���e>J�Τ�:���%���w�����v�4����3�ڷ���B�P�B�ʑ����;�ͭtR���Yn�(���i��ݷFO��wq�a�� t,���Py՗������n�U-w;Z�9������7�\=4��-�+5"5.���}�.7YWZ�J�����λ�\�9wS��3�:�=�O0�(���n,��{Wi�=S��aw3��^��O2¹�eֶ���B��Z���==�S����:�CED�v\yl=��3�,{a^�	1]�nc�1�p�[�׀�)��g!��i�ˈ�}�U�^b��阌X�&����F�J��ro ��{��u�@�2�!�Gw��fl���{|��"���)
�
��0J���ː3H�'���iiI�����ܡ����t�V .��:rx:�2��������j�Jʓ,ebQ�^N���J���]QvF7��e�>���5LZy�&8)�wfr��Wf�䶅���P��IQ�u
Ј�j���ƥ�c��GK/eu���������pJ�][��T�>���&qup9R��.�j�E�]�ւ��^>�6�X[K�HEfuʸ�aDVni�z[޳N�+YS��<xQn�S��FA�+'"�u�N�*�x� /�ҹ��C�u�ܶyQ`V7^N+9���)��ߥ>�z�{E{KN�Q{�=���j�3�F����YJC7;Ѝ��`��S˼�f<c�l)�eԦ����z������:
�.:J:��z��.�m��V���P<%=.[,���7N;
� ��љV��绺g7<�f������v�n���aIP�+i�D�P�4�J�|��X����e�f^�p�YS�[�щmu�������8v���H���8f�)Bm3�������$��땏��et˛wS���%���H�K8�qu�s^V��/��h�Kۤx�(hEl 0��\�����.��%�F�T���I���M�1�+_r�o7��}�m�K�����p�����(m��j�<jp�Y�q�%22ԍ���{��`ݤ��7]|�T=L��rjSͷ�'[cv����+_F��������/ �]�;�H�&+f�'�;9���m>���ӵ����7.C�H<�Z�(6l�S/8���Z�:�[4�[�B�P�ݪ�4f4:�A"��'���I��ܷ}p�α��C.뺸��Zt�HV�Ô�.H����𗧬�rty7�;~����F�Ɲg5���),N]�Z�Vv�ۤMo=.gS�ܻHÓ�A�n�fJ��y��@�Y���`���Q�_^���w �� �Ad�,�f�h�&��滃�Yn��}���)*�1sn��v����I�r�q7�Eʣ��C�����׭�c��Hx����lڈ��:��(ȑWq����l�q�<�fq�{pr�.-��ο�����.���E��P�Ӕ%�:������FZm�J�o�u`ޝZ�ek:���v}f��}���a�+qKu̫���Q�F-��	��BM�y0{���2'�HWϱ�@N	���G�V��[g3枖�t��y[���o�";C��0/�"kEε�����a��("�����*O����M���+(7T.���7&�h�D�$3
r�/��>�:̂j:�DyN���n�N-x�[�o�,ڙ�C�
�)t�)��|L�8F�!wQ����ЭM�A��%�ݲ�v�M�o�N�Ȥ��n�'wz*(%-���Cwk�ƍ-Wd_qR�O��jK�WR]Oq�f��G�5N	��d�����4�s/:��ON
�i����e���quy�����bj�O�QYB!L����$��a�A�.V�Zh�&����7J=��D ��Jy"nV��g9Ԍ�YːnՇ��DufJm[��E��6fMVbK�%��^̵���	�I1.�L���Ш��;)vx��i�a�JF��atO=����m\�fФ�(��M2���pPI<!R�I�{v,:�3hE�nR{mb{0ª�H����N�$(b�^!D��%�g�����P�Ȧ�f��R�a�z�jBrNHy�J�!'�Y�f�4�Ě�"���z�^�V�ᴎ���i$e��	�Z�[����{]J��C$�63�J\��I!*SS:��D��R�z�g��֭l+��zn�V�3v����Xb"$��b�g`s��Ԉ�F"D�]��I�k3����h-�2ĽKrB50M�0*�3��|�����o����]¹�i�Wjg1DWu���Zו�C���;3�"��\�J��׈��;�ṸH�b��,����""fq-ʥv��X_�:GT_5�!�p��mt9}�^�^b�ǰN9�����.x��r���/��[K�o�p{��;��Ͼ�J���� ������p�Ș>O�oϫfu������LS�^Im{���G�択Ԕ���ZѻN.sm�ڋx\[�QR��k�#�q;�}45������#�զ���9�2*���7ck��18��:���KʍM���{�WWv��J���'feM�q������䯸�m�gP�_���Dzq���GY�Vf�F����wcqs�4��&8��~�t:�mgP�r��������ə����T\6�m��j5;磻Sx9�2����v�!ԍ�۞ZVl����\������FZY	��{��:����rs0��n�K���`J{���ٌ�rJ�-s�Z��]ơK�Lv�F*��Ǹ�����U���� �%�Q�7�R�鉜�sU.�&]����m!@fQ�o([BU:p���L+Hɒ�|^0/����_���u<��I0�^�.�BfNc.��k���;r�:�GSNR�tGQ�4n�ԝ9j}�Lc:z�"��i���7ƴW��>�� �u\�CTy�#P�YS�	�d�w��׼2��ٽ	������f�qO��X���t�b�ӫӍ
�l�Y�ʽ	w�|ۼΠ	� VNb�i�I�s��9��E��˴J��һ&���VH��*75�����v���IX�mѨ}�u�]@��* ��+r���6�GK�Km9��%�ꚍ���T�����q�X@ud9}�r�37&�R�=�#�{=��\�󱋽��O�c�E�lm5.�x0`�Y/+\���qh�����yq@��ci�l�ywb��nD��Ѥ"�|0��]T]���p��.-�.;G��Z����Բ��ZRf[j���:��NM.;��OQ���c�T5�p��!{iu.�<����n��jCO&����'���^��z5�O{�3U�_�v;��c��_T�ۊ%W'u�j�&���k7�R����Q���n���H�����
Zt=o9�y��t����L��G5��t��Ҵm��r���^��&��K���@ۛQ�Ӿ��r�9����� ��`:'���ާco�-��{B�wo�qs��W\���D}�}E��k��Zx�zZ�#�W\������{�	˚��;�S��BH#N1�7Jv��,�|�U�uu�O5p5<��K��
��q��^'�����7��R� �QqR��ʉ�1)���%uF����ȍ��qV�#D-�ʮy�̮��l���1���0��ʒ�­5���"�iI�YF���	�Q�k5۩4��>|�LWRW�6ʿ��U��YS�1����4�'�ߕNud�=9�,�6{9�O�y���噥(��P�s��Z��Q��V[�K���|�z�3\%���;�g8u����f"����]�R��x��E������J��/q��5�v�
�;�t�S�eC�!t<��������z�[��7�F�k5�W���Ŏk�Ž�V�<���>Dۨ��yС�P�nM��mߵ��~�Ό��[E.�+�+��'�>�����D�����p�żWбVK�^ڵŬ�����5�0u��2�u���FFWY�V�N�3�F�Pf�m�xGx�U���w��DI�D��X�@���4'.�f!�Zl��F;[�x�bͮ%e�L�s�m蜨Jj]�t��i�3vm�Zҥ��着��gn���!ը��u��������^c���^qC�K,��V)9�1]�R���8jqE��Q�(�7�)���������X���L7����y�]�z:�N��׾�����7����[�V߅鎳��ۺ^J]g[���>~����Թߊ���g��k���΋k�[�J�ȄĢ�Z��4�/!^a�T��*���ʏ��K��j�����Μfp:Mۈ�N��s����m-t^�t�E�ü�,�w�UO����e� p4��3�-nPY�)z�/���yVM�uE��>��|��5�m�N�\Ms����׈wjo��X쾎�:;*$�����+�	����3wW:�q|�rҸq�)�;QS���h�Q��$�l���;�#Rb���L�[�kX�wq��w�K�
�z6���ܲ�0�W���@4�}���H�h��H�Y��ˣ"x-AE-� 3=�8v3�@7ףM�~��t2ԃ��4Qۜ:�'L3�k,i�K�Lx2<gIv�m��N�]˱K�:+Rƹ,�9eј�8�9Ji_u4M��[��GN��`�I��r��Uvi����[�_UU}G|{��ls�#3M���ۿD�9w�ͱ�9�
��*qi��)2�s���*�{�A���p?J��N�f��}N�L����������oJ�n�#^�f	g1��RɊa�a�X��
���r�2V:Nɸv�ͷ�Nv�qy�	g�r��m�ׅ��ƗTE�*�zf1`=R�v��*�?y#9���[�=T�/'J���t`.�63�n��rk]�4ɞ
�_���t�=U�������5�[�~d���������쀸0q�v�PԸ��������bzkT��Gs����LF;�_7�2U#������t���tZq,��~8��zn���~���[7�Ǽ��@�g������>��Qj��i��yѵ�q�F(�_iy_&�Q�U�f�o�gNȣM{yc9�lOg�?Er|�W�mJ�Z�Y�V_ �d�!O*c��5L0m��,kW�d0'5
;1�,��������e�%<��(��\�s�챙';�50�uO&���)�����ͮ7�����S�jw@`�W��*P	A�Qnn�����ā���z�}0S�K�j����r�:������ϚO���q�t_�ޙC�^�9_y�v���Y�1��AaZ������*��j��N����5;磻m7�_+�m�����E>�5S}K��]m��zѻ�1X�\F.�O]��J��[��e���,CbRs��Fht���i(��p23+�;1�
��<�IE�^�}޶���in�6-7�٫��$X��ATa��F����`'�pe�'K����V󶔥r^潣w�oN#xk��Y�Q����&�Z�����+�m�ozT�^1�n�U��Yl�F�.f��k�Y_>^4��nB��O�mQSݩz|����c33�Cdr���6�UI:w�|����g�̾�*�^����sP����w�~n�˳i�eIq��6�r	�V�@u���j���w+z�rU���s�u���җo�G���b�gܮ�����<��]2O�0�!�U��g�����ei%��P�����s�u;�8%�j�Q�;�hm� Z!}ܥ]d�{��u�*�����_��hv v�57�$�>W��!]� �������˲�,r�y�y���A����9��������Wg着������=�'���r;*;�����sñ�+��\�\��ۑ\�ޤ�Z�OB5���5�.Z2�����u[��Q��Td��b�����m���}��Fq�瓟?(<ͷ��[~�:��s���>��\Ň�I�)���k	�=�*-7�I���9��3�,$:���	�iݎ'�=�m�Ɵcޞ�4���}�1y܇�g��#F�zFv�s���|^��5�r���TC��7Sǭ���ԫԷ2�j�Ǣ�V������N��3�]g��Y���O����;Ҹ��]�E�G5ct�I:�N�Ff����ᄨtvT�%v�;�r��>�<��k׉..���)�N�N5�����[\�=�9O�5*������w5��}������|��Y���֞�WF��嘘�HuC0�StR�~�N����=��:�p.�k<���|_�j'\Nݲ�X^.֯�b;�Z���n;���x�l�N僻��]�i��D���}�U��[�M���[W���l��؛}ۺ��t#�i��6:�޺����h�Q� ���������TCt����5�����Čr�S���ށ�2ƵK�ӝ�p�1�	>�c3+�Y�з�r!͉0����M�s�9lo8��w�m��T��t�SaC�S���y�)w�4-U�{�\�v����Z'�/�xg9��Y5�a\&&~O��&���F�jL4j��e.�7�jV�� Y}�_gט��ŀ�y�w׋N&gS��%��S�����z�z�9t��W����;��xo1x�];cyS��d����,:��sCm�8�|���vTA�uoR�D���Lx����c����.ߜ���d�������o�[f��T{n�m��*+�����x��5��O�oǞ����<������ͪ�󆼢��11G�Cy���*{{���i��
�Z���v1��Q��;Zx��QO7�hRڪ�ыu�ҝ㐶voi���{�hڕ+Z��������Άw�=/(0�����Qs\�H�=6�kմц�Ǉ���N�m#�^y
Gg|��F�R��&Sc7�=H�o@U�(u��p���i͠V��B�:9K"�떜��q�Jʵ�¸��}ܫQ�Vm�J�@�\躭�?g3xں��9ui[��n,h�7��W�V-��)��fs����L��5s�(lm�J���D�>K
|�k) *o����'^�w��z.��s�x֛����������^�K=�K�*�����'���J>|;��N��9�Ʃ
�ەʦ7'^�-�Q�%�:��ۻ�]1X���Ұ�B��#.��jQyU�N*�U^�ۨ��`mc
��e}*d=wave�9��Q�����	�-�AE�ӥ�U�/ ��{�h{��^���%`�}�p1�2�؀�cy�_6ՙ��;j[ک;]=�d��VZ����8:e-�K*�u�m[΀�/�����O��װ�V	y�UsP�����\/sџ��(��,����1�1�n��2�^����޷�U}��.nZ��l�
�l+���ۃ�y<���@�Ǘ�@)�ms�ImF�qGt����c��5��{@�-,��Z��'��1�=!�׹;��U����\�H�>љ�mI|�}��B�Co�(2��x��ը�Дy�j�tfI}6���1�Vl�ի{X{�\�O$����HJ틜���/�.�Q�Tt-� =9����֦d�L{��f698횗k:r�7R���������^o��էjo�sh�K�A�>���痺�}���fY-�"5;���K�B�hv���u�ߏ���^�~�_VL���"�����$��V��C3��I���V����?P&؞�y���K�s�
ݵ�o�����y%��*��9���=�mm���5����Gr�$�h��mjt���*��_ͦ�)����ʿ����%T�%BS��Qqq���k����ga�$�3�-Z�jyp�>ۄ��Wˆ������=�e�����c��b{9�LK���Jx�ȴ����FO��d��������iy
r�x���*�<���i#p_u&5�RbzSU��ڏ���i[�Q:��:oUuݕt��&Wzj��"W{>ސ5p�x=�ާ���mV��}#mc�0����,�(�D5u�ad�����َ>p3�$�6%�M.ʱ���1X��۫��B�����wx�2��Z�W�j�S�f�0���6i��g�A��W:}ͩ|k�s���u�3�;!rU�����Yn�V�A4;�Kڝg+��w�\!Z6\�]�pZ������ԫ���x���)
8�$3��GX6�+�uu�܃*�p7�S��pCͤ�-��[}a݌�ɕ+�T�v�	c�NPUum���ttR�]݊�u��^r�YLX�hnX\��F��5jz�R;7+R;���9�Ր��7�P�������ށ&;�bcbw3 �=p�|��#e�� G����$��*C�5�};W��Q�J�4胙R�q�����u0azJcE[����·2���f��XM�Y���/�6��9�9S�e�Z��<�u��sT}(�y;�C'X"���l���B^���_M�G^^�N�YY}X�d8��o�S�8*PI�+w�J&�+4/�V<�53u�Y�6��%J�VZ[�V�H�j���+-�|U7u�r�Om H9Zs�;Ou֣�&U���]Ѽq!�֋P�G�G�r��Q
�Û&�8�fL�`��t���!}ǣ`�zt�Wq'�o�W�^���ˠ|�
&��;����;88r]X�=�4Wv�$����c��K5�;��ED�TT����׷2�\췖�/�H��mֶ1�V��y� �m��ZVR"��h�����1*Y�(%���kpD�H�؄�c4�j��;��A}y[t���橕��W\�*�7aoN�o�I-�h��%(3{O�:�1α	F�vc�mێ�S�c�*s?e��wsY�ǹA�p��#%vV�Բs��%O��Ʈ�\y�6��]�/�/oR�˰:�Q� Tr:y��m�P]�5�u[;^�ݥVA�]&��FB�B��O���3��I���i�Jtc�J�Z�˾D�nKDf�!�2Tz6r4�ܔ�l��]]��{,�7���yL�0�&0j�v�.�48_�6��pZZ��E��e�pws0]	On9F�%�v��Z�R-�Y�kF˝�� �����(���,��h���úh���1u��W|L)^�T��HG�����i�KM؛]Wu�����Ӥl�����]�W�/��K�E�'ٜ��_D3k&���ap=��*u5��8�&t��_�j{�����O.ÃҞ��M�����������J��'��:�1���d��a��7�,��os+��W��\�����˙ٯ��t�W:[�:���6��9M�m�!&j�d����c��2�JD�����X����G���{X�.�n9I�3^��t��/�'��!��ZIŖ�n�`�nv�:�R�*�g�I0=r�C������l��
���[IR�vh���T.8>��7J��ܮ�b4��ohq��'}��S6�M�ҭe��Z�4�[�{�ar\1;#*�oq� ���K�:Q�\���G�r�{d�I�Ad�Te�j瑢&�HxF����K�yN���"Qs�L�
$���BE�"*!EĬ��Cȼ���3
��<�,,H��B,-MrJ�s��T�T�/(D�	�BDJ�aPE�zezaH���HW��e$jnzE�xXU�%��B������9�<J<�f��XU\��T[�c�EAU瑞�E�^�k���F��h����Y����xM=OHO**/�ԯ	UsB�,\�V���gi2D�"�D��̩!r��L�������<�W\��D�,���)�<��L,]�)0"M�2�r����b��Ӯ�[О^����f�
j��AWZz��{�$���vź��3���(Ry2)�Y�iu?�����;��_����S��3���|�9Q�	�LF]�U��l��G����Ocs��g���\8��ow�ŕ�NC�QmS<	}������:whrѩ��kN�<sQ�'����!զ��)��#EfT���*vWr�]��pieE�:�{_j�g���w�C��hiʍ�p$�/]r�=��9�Lo+a`��uj��Pq]E�Uy9���Pb��y]%��c!]��5v��T��(��w�5�׺��\Zgض�R��]F�߰�V8��׆'������R����]���=��`�dU�ī�����4�o	O%l�N���IkJ1��ϯ}״{�x�]��w9�m�*�ό(��<�mꮱ�~���j���޾Mc�n`�޿���-_?�ٍ���������@D�E��4��'bu���ƽ��jyx�]�ގ���YQؠ;c�-i��ܖf�S(˼�����ލ64\O՛l�w`�53g��XJ::�����I�]�S��s;��7(^��rY���,�������u�{;w�u$�d�ך�>}25V��� �XFxMϔR��۩:��i�F3�ﾏ�%Ô�\�s��)���J���Q*��+�]��P4�5��dRQ��e��v�5;;��O��0�(��!��W֚ˌ]�Qw��%.�sJgqi�|;S�n�%l�*��U#�6;��^��^��Ҕ{7v>8����-m-}H�Л����#�_3��jEYs�����ju��w���d7w�9�]��s�ؾ�	�*�a��,��\���&�2V6�9�N�����1�1\Kܚ��n���]�j��o�N�D���Z�c����0V%��O�s��oPZ���h��Zb�z���T9��M���ZaeԾ�4�1U�8����ש!���M����u�J�6��p���˘�U���_��F�6����E�=����8�'^�~���ؽG�yF�����r;*�4D�_:�$�GY����u=1�2ga������,oD�վN,�Op+���+fA�Z�itnB�5*��M]�x���u���[s�u��<��#�Z��f�M8�Hwb�I�w"�J_]@u�][��O0��⻸J0���W�7�	2��na1آ��Lb[�����nw��.��q�Z��Tw;zS޴��I�m��y&u���WFd��܂s�		����˩s��}ק����~-N�)��r�%�=�W��6��+��&����Uqێ]�9Zӯ��{�M�[�/�֌��g����I����t;�������;h�O>"-����:ǔ�]�.v�]���W�z�.�{�J�s�Uc��[���g�,��G_�+vզ7u*Wn7�w&�o�97��m���ڌP�����[nFcv�t��k��f+A�O.1��zZi(|;�ތ����8�*��QJ����X� ꧣ��d_9'๫�.wq���q�/��'�yU4�}���1WEe63����R_s��`-w��'<��:�C9��6���3�l1{]�]��8R��t"����[��,+��y�;���*lE�����/��y��=�r�����mˮ4�����h�Y�m�nwh������\���Ta������m3C[c(�3�ow 2�µ-�y���D��VE֟&P�G�p4$L����`]�_���.�5�.~!�f˂LU?C�2������-�5�f1c�:�η!�g��h����s�m:.�eWɸ}jr|����R�o�K*�:�-��^�V�zl����ϝ��&|�ߵ�I���а	���_9}�hCɢ���֙W[�Sx���s�c�z1D�S{�8���U	����o)�W3�1�y�ۢt��,���6�뺝�����'��A��Q�����d%�)����	'zQ]b��ݸr/*˜���UF(�Q�/uC����h*�](��&���gE���r��v��'���!{~]��.�}m���\�jk)���_[Ow)�k7��:�f�ݍ���C�8%ۚ�ᓗ�L��Ĺ�+]�C[�o�}�N:[�O���D�A�ǀ�1���8+{q��7z��5���?�ȚZ��O:�����y;������8��x��D� �n�it35�q���W��q�m�Ibo���+So�^���5�3l`���9�m�@�./U�[8�lj��y�z�ǽ!pf��K����d�ũk�K1�kl��>�u���l���q�]%zҎ�����h������ni:��s�.2���zS��˱t�'�jZV�v<g2U
���nΉ�S�7�{�K��wы�)wR��b�9��6D�=�Sao=C'��E���0���0���4��P��hF��v<랼��X^�.l_�p�;�Ì7xG[����(^�1P�e��⢖�wkr�^uk�u�����S�s�f�<4�09nq����΅��CrG�q۽5�vf���юT5�9�3�6�j����|2����r���S��ZҔ>a�����Rh���[��>D��mV�Ԯz�Ft��m�;]���~)q^K���}��ڧ�=]�)���z������{���8l�o�~m���eŴ���o�b��a�;z,�c=��>Kr��@�)�Q��x||{�-׸�U�6پ���O+?V$"k�QQ�iD�@�}�&��3Kdf≃��cѝX�r���	�Ιu�-�۬խ�C�[��4�;��Aa��3I�����9�#�/"��.λ��F���1O����0^�
6�Zn�q��1N����xB��}W��綊o�/n �w;�Zع�q3wh$�=u�U�eI�<+�.���F�)N�;5�Uk�5pm&�wa�θ�V�����F|M���`���^����v�[E�*-'۔�S��}��`Hb�}{��ԕ3{7�]�;a�|{}�B�~��(�����[��I]�Sٷ*��sJN.v�V��b]A��R�u��ʾ�:��]�����k�O���.y��{�1��v�����o��UD�¢�R���\FJ����аX�d�T��~�s��8���������eS
�(T�L�`�#��;�K�-{����{A�]"���s�Ng�T�n��ѓN���,*�	T@�Xx���}lT����rO�U��izej�5
u����Ѫ�-ؚR�1i��/{cc%u��I����W+��}�Nw�OTZ�ܞB���@%=To+����8˃B�E{��u
���k�7]Y�˦���̨}�b`�.��.����ּ�e
�싕�3\۸����Օ�������&:����;F���~Yl�I��/�j��C y��e��(�*8�Y�D�/9|re���`V���o4q�-�0v��m�G�g�q�E������'}�78��0�yy�I�vrT��V���UU�S���g�*���Y��k3ё�����K��_':���t���{I�&{*���Ԡj	�V��˩}�]�^b��fc�`����qS��'���%~����r�+O�K/����m�^O�v���V���d��wX�R���s�8_t��Oh��s�̨r@<�X��sU�Ү=���K]E��F8�Z��]J+�����#^q�{�-���⮛S5��3̉���<���x��=�Ի^g�o���r>�{�긍i�ɘ��9��	�^\ߊW塛{��Tf����T�GkO������T��1�-Wne򧓧3���ߧ�3��C\�;F�{Y�5��Ŷ_;N*��Y��gWjIn�K'v7;q��7�M�J��X��"z��¢���z��Bu]�Y[��kq���j|�sY=�i�����m�(Ufy8%�Bm���6��ſ٫&��%#,��+jdBe*�ƥ0�XZ�����ջ3Pr�bث�)��{ ����$�z�fu�5�\u5sX����wD���t���,��ӈ0Tv����t�q������j�T*��hCr+V)���A����V-y���p��K/Rzu��h.��i�u��V��p��;|hn�'�*x�6��c0��k�p;����.�_)}�	�p�o*YYJ��9�!���T�:�i
�ں|��\���$j�{zE����&ٔv��ų��f�W �L�{5u��NHw/)b~j+0�k��V�Bwz��R�p���k�沝��y4f�Jh�f��rwJ��s+�J�a���Y��:ֱKq��Z-'�I�K|����޼��J��8U�����GL����~R�לIo�k��f1`3�?oPU�:����8��%�sS�c���j��Ң����O���N���]C�7�?=�.!���j��bw7��4����d*�6�9�d[�Q�������Tw<|+i:�����=K'^#u.�5�G�}��+o�������4�n����6���4i�>^V]Nn�v�8Kf�J=lvd�����o@Y���A�'��N��%O�&��v%�f^�T�ڵ��S�	r���w�:�{"b��l�g<��Y+&e6G�"=��g(�q;�;h./1��Xx����wY�w���^�ʡ��(2��[��o!�c[�Q_A~���+Ήjr��,�=κ:�u�i1m<Χ�_'�o��:�b��ݶ���������'���8� ��C�V_+�*�kym��)���X�k��;��:nN�����9 ����f��5���7����תE��{B�݁�h�2�gs:?T)��)V��J��+��T��k_+�]I��ZV�-�cME�H���d:��k��N��gX!.�B��K	pϭs���X��uKV �'SݦLo^fȶ�M.q�����.����^K�r���'�av\�*z㥳��[!>�F�u��sGZcS�1�I�����0�k�]�'���yr�2����cVe�w1����Z�|�39�U��eK1G{�:��%D+��*���n{��qf�{����D$��*#p��܍�5j��m�٥74-l0˲��+{�4J�{�v�2� �@P��+�k˯rR�?v��͈]�h�*�o��ն�]ѭ�T��D��]�����ܠ�Έ��n	����+r�n�	�kFt�oeSR�:�5�3�X�^���p]p�S=fL�J�[S��F�����fҭEi\k^	gU��'��l��R]��]���qc��ǽ�W
i4�r7-�<�?������������A�)}�]��*�ǵ�A�Ҫz$5�0�<*+6�ݷy��((y�6��8V+!�l��8���o�b�]�7y�����G�e8��Z��z��3p�\�lۃk(�8�}��y�|��>+�Tt�~r��Y\��ϡ=�yƞ�֬nl9�%�w��^�թ�3:�ƿQ�Q�ǖ�ZC���'�P�es��m:
aOe�*s�e���q�t*����}J�⨲�_ڧis{x�[�M����\�U��w1Vy���U��y�v�� �8��D�����|5<����:vZ��+'2eo8�Ck�y�ƅ��OT�*��+�]�i���W��KŹ%c��лn��.۾8��	P��.~)p߾�"���${)�����G؈TE�ճmXe���D�0+�t*\��˶���K����c�n�Y���zЙ@;o���#:5v�c�k��*�Z�]ڜ�c����S�u��.�pWI�Tgzv5�vm�vj�ѷ>E�[� 5|k{���,P��U���B���v.��I[7���Ҥx���_*���o�o4�Έ���B���E�P]Vf�Ze��� �+��tR}+�R�b�F%,��۸���p���6�3��ثe���#����l�tK���S��ǶbZy��L;Zb���&R�ɩ�] ��k���w\��^(�nNjS���U�G]�˹���*ʳm���7�<�_Jy��c����-��y�r���������^�T�eEV[�������� �hnecf�h���@فw�R�_Y���"����D���h
"��_˒ȱ擲��+���7�:$��<,K���/.�c��Ǟ��gh��0	�A���|�U՘q���2M�d�
*`��+N�g)�v���u���3��R3��+H]gB��
��5��������U��]��3��ęÒp\!X�|[��sׄ���*Q�kw�=�=܋��~{����M�[��Z	���+q��U��7)u�:$�	ؗn��W�e��d�љ̄�,�Vx�S�*�4�V��B���y���g��g6Oc��5��>���U�w�a�*X)(�]i�Ĝk^rZW�I:ocum�
S��g��aU�s��|czm�֋v�w�V+���H���Q9�;N������Jj��-�ݺ��6��u��3*�}�*̩o�M��6��rִ��Gw ����H*�N�Akmg|�uv��vp��N�6F�+Cn��t�|o��H� 0�9Y��V�3��i��E�������B���tqF"x�.�0cl��V��*}/If���#A�϶���`��h�f��[Ӏ�9@��mc�e�e�,�Zt���Hv���gc8�a�.$���P�*^�(s��AkRtR�ՙQ&`\���A�Ә"k1H��˧F>��W�����b��!��m���Q��$)ǖ���<qSrK��Y�9DZ�wX.�Z�6q��t��i��_S�r�����Գ!���1S<����W�����6�.�$j�>�����2Z�t��6槟.�+�����7�k�Rv㭝p_��ʱ�f"B�{ӰT	�<�@]��K�,��{�c��Ī#�Ү۳|��']u��F%Z�]gh��γ��Sr�T͋mA�-�*0VqK-X���ow�֪����r}Զ��bAc�8Ir+���dff	+�U1F��4�� e,�ۚ����>ё>���][��-�H���-)٥�M՗zVкE�������k��#}�m]m܋/D�F�1x,�<��(em�N}֎�|������	�tYSU��`���Z���B^b�Z���y���28�;��?�����V]Z����iR�i]\�/79�'/#{&��e��'����Q*
�E���a���W���{����z���*)T�
�Q����#§)����"�UR��6�ʋR"�p��*(�"��h�<L�1(ʔ��
�I�*��**���E�u��$�BH�3r�IDWTܓB��%4(�;l��(�H��*��(�����C���P�3���j�9zTE�G.`EEn�A���G�VI��&�yJ%yFXU��g�fQU�!*U$$y�xUG�.y^T^T^QDUWWk�EE)�A�����DT�EyV�yrF����D	�[��^QU^TP�\"a"dEU��yQxF��%ȅS@���Lt�
�I<򌐽#��� �J#��Td���ͫ��
SR��-US8�X֌q�����ֹR�J�ܶ����s�%�3q��4Ƣ���l�#b���Y$Jr+R{L���:��c�޾���9[���.6�U�ѭ\CѓN����_%�5.���F+5�Ox���7:�6��R�:�_\B{�\=��v&)J=��/)8��y��j��f�й���� b^���2�'<���o��M��>Νf�圓��`�k�YT%H�
����5��{��s.����t��� �fT��$�}S}����|�x�{rU��X��e|�{6�,��5/<�a#ݨޕ�5��s&��KL,�����W����%;r}�[�� �-b��9c��zuݫ�!������c��Yq�����ͣ����e��),~��P�z�&��b߳�8�����8��ZQ�����2�|��M�	���<��7��Bc��[X�}��{-EG<hk[�k� B7M[�H����<�Y��	�`�r/:��vq*>{���kE�\���wQ"8o��1������MZ�Z����v�q�qە�*���v���gh��H�Uۤ�=��-+���>�J���j��߅9g@�4-G"�!����V��[Җ��K�&LfUw�뽬[|*���0nG8���|Gp�כ7f��˛ʳ1�������������Gsy+�:[�5���z��]=^{��[S�i���jf�1s֛���5\����[���P~�j��3����A���g2ӎR����k�)��7�7�SؕP]E�� �� �W��J#�3'ycu��y��p�����N��a+�P��ڒVj=���ܯ���R~��zz���Yq����M4����z2~N��7ܷ3!�ؠ[���ͥ;2w�<1��I��U�\���J���}��/4.�V<�So}��{�4-��H�LA�DW���gL���u�&��q]m��6;6]f�j�k�sC��=��̢�t5u�y?W�2���l�6��*�x.y�]^�"]j�ͩ/���d'p224QK��[٫�Ӈ1��Js5��F޽��1�AT$�&��D)�u�W1�%�d����m�ڜ��n�l��\�4ͅD�÷N�I�_�X�fL;v�]X�L���ŇTX����
�0˙�ܥ[�L���Os��sw�A������L*r�8[���,�v����t+��Z�a��{^���<�h�kqU�3��Ncz���A��o"�2�K3P};=��i�j�2�JZ~��R��W��z�T��>��m�;S5.��q��㻜\wv��E��>w�ٳ۾S�b��a�-�լ�[[9��ݮ��94�9ގ���/�cm�6V�\HQ�}7WR�������i���5i����:t�'���8�=��	`ݳv�Oa��|�2e�y:F^f����ޮ�[sbb�7�O6��[���儨��G������x�us��z��^��=�ꃱ���:�=�_���K�q����߇����̌_y^�t3f�(����gT����o��]����O�zhc>���p��H�C�xu
��D4&�1�Fb����d?�k��{�~���8�V{�<چ�[�\z������]1�Rk�/ʫӓ�ϋ�:#E?_��>S�Yy�Csd��ё��%�@�KG۳7[�����"�x�pfE�̊�N҉It�݅VxJ[<��us�7��){mB��% �j�Η�]�eg5�U�y�ط�)�MEt;_[Y�r�)�v*i��a��0m���9�e�#ՠ�>�#!g;������Ñ�r�ڳ��mǸ��p�b�8�[�ɫ�gﶝ�9	��/�{�EG��w#ޙ���L�ٳ3�J�|��/c��p����o"�+��W�g���Qm+��u������(�?I���n\��T����{�}��޹��n<��s]�J��"}J{N��ÜQ�և��U+��zv��|�t��lϤ����<��V�!n��x���#��&�;o�LO��[F�\�wd�6��VK�^7�P�N*���ep��2wǽ7j47ǜkP��T�ܛ���en�w���Q���_�^)+4�9��s���u"=3�w�#x)���5C|B�$lCbJ9~��]�l{M�n�<���������~4��j�f2}�S�'�Ԫ�s�{ʨ�4�����ǲ�8n<��s�$,;;,e�z�;����o|���}�,��kG�e��oֲ=�75� w��+}�q7�m�7���~�(m���MK�]
�O��+M��F������`vϳ���~�#|�G_�l��<�WqZ���g���}��n�.*�㇗��uV��U��g��z}��/g�H��ב����~�C���hAӵ~�1�0m��MhN���	��̼�umzqU�r��廎�a���<�ub$z�wZe�\x�XgU+_�rΰ-3kںN�P��Ԗ�\.:�nw^���ܧz_I7�ŧ���Y9�S2���������+c`6/;k��@-��^���^6cٺ)x�vOmT?�WLa:�FL�'��ƾ�{O��߼Q����}�8,�9�b��g�o��_Ob��M���j]�q�S8K�}����X��L:۩��Ǖ��x��<��˥2�z�4)x���S�Y�z��qPf�&)��_\�9tLzG����y��[�ޯ1�}����+�����7������o��\R�e� &j�	\UH�?C���l{�j��f<�'ЧB���aT[W�m�[f2<���{�鯯��x�zK�ٸ]�o��i?d��%=��c�3��V�����r�sO�Vա7�׋m"�>�.��.O�7;}��f�gM�_���i�hقǶ�1O��v	h��@�=I�G�#Ԫ�sӴ�X�1{���Uw6����p�wnD���F�\��#�2�W�11O�h�~;��xj���9�w5^�l�ˬ�W��ן}�J�oc�\ w�@LW���ȉ���c�6�u��5^�QG�97�������S���T;��e���Uh�@z(�����-&��/�kC:6eעgس6*kWpzV�b�_VAI���6^�e��4�tX{�F+gl*�����{�,�L��'j�3�)^%1]bқg�����+7��$�{�eX4�;�޽�r $x��@J�,{��M	����w4�{�Q��MO^o�4�i�ӫ�W5F}҂35�(+��q��T}1q��Q�o�w��=]�?e��'�����UҴ�����{C��V�a�8w\����~����[�ޖzTo��M��gL������ۏH�W�f��>��,�ه{��,f�Ì���`;�x��^D��C�s~����lytV߳�_O�H�-��9��ߤ�YP���ÿN��� k�����/{���������uZ����9�:;�W�.���,�L���!lb��d��pze�3�;:ü�ʌ&�}�k-{7�/Г��!w�|_o�7�G�w��D��d	N�@��0&/�p��P�#ћ�zv�o�~w�S+��9��:��~��������U���+=�3q*@Z�oN�շK=/HX�lR�k�������\��9�,~���`S�tg��qo�t�����=E��y㫓�ll־�ܵ�TL{h� ,�UH��ex�o
�{���w��8g�鋏p�����۫��H��4]���u�٢v�Ѷ}HT;�2<���n�B+԰�����j�$ds�RD��z�Ř0��_�r2z�+���f���B��VwG+���{Fp|�R1�a�.�^�	��%�k���o��J�/;^��A��Ņen�7�����e��uZ�P�'r`-4:����`'^�"ԢZ
��[-�}���'�s �I��P���`���o�bV�3��)�ױ5{�o'?@{����[����5dy� '����A}^�G3���9�qZ��u��E�^�ߢ}�O�jM�<
�~� ;��ȯ��9#�G��`xc�DM9�:c��9�^x��|�����^������o�3�}'m ���*�W���T�4xԱ��:7J~1�uR�������/9Lȯ�N���W.Ð�9׻&=�H;+�X�:�/���]:����w�o��9y���x��5��Z��<:Nx�2���r�%��C�����顾��֦� �Nz���Wlψ"��T��}��+tÿ�k�o�<��L)_��>��ψ1�J\/AM�E�
�����M�����r�Hq���N��G."r��ʫ���x�X|1�. "���z��
��e�����~�εv!z�#Q�ι���q�x�z���s��^V�+���Z�T�.�5^�«f��s�ps�Coܬ
��犬o�gj��=�ED=�;M��z���׽�@}x�W�t�����$�[�s9�2�����G����������6���<��6�t�Ͻ�~�f#��ϯX�������(;��4��#J[ϺaR�5�_�n�i�Ȋ�jl>����>�G>��F@��]b���VxV�+�sH��&�v�F��נn���G�a]n�ǣ9��� f�V�;�޾9�q^��΋j)��5eۨK�ӆ���"�»���{1]��l�\dγq�>E�s����<6<�{Ƕ��5�b�f��Ǐ!p�;���v�f���7��g�)M�U5�@u?Je��B�|X_A��ћ蔏:�l�D�{;>����;�8/�;�;�Æ9����}D�D�8�h�J6��Qo�q�ʔPޔ]��G�̬�W��o͟4�0��z��q��x\��,����<sqFG�t�����23����ދ�.q����єys��|��E��y�����[����.�� 6o�0y���UCr}\>j��L��})���YP0,7���8��tC��x�w�G�J>����e���w���g���������ӄ�)Jg@�Xs�c+��dz�_�3Ӵ�3���
߶�b��T�����{�)e�x�i�d�=�)�ɺ����bi��7������To+�X���Ҩ{Ҳ�٢j�t�g�����e��K	�L�z�麇ו�a�z�N�����ᢒ�L�c
��kC�Y��{׻Nr�Y���5C|r�DW�bJ9��fǴ�n�;����/���J�rvɝ�+�#g(�
����}����p��5غ�z������x�/���#&���Ќ:��mT�ۖ�n�w������݊	8����a'!2�3�h��@���Fӭ�)��*�5M���z�rP�^=8*��\[���j(�3�B��/FEw��#>��t����=���$��������hn'=�u"���uc�p����}��g�bռ�g��o��E�eD�{�gM��Ӣ��P�7�O���������n��w����aBp��F�o�k�O TZ�g��u��+ڪ&�=������#��v׼S>�Z6s���V�	����� 3�Z�}{m�/�n��W��j�I����x	��X�O���^x����Q��w��XfW�mT��ɝf�g�<��ю�k��'���1\��c<d+�N��6}XW�� ��^�c�Ƿ��C����Jn&��1]�xe3y2��G{}|M߫o	F}:n�a>Y�k�~��Zrl��S:V+�ȅ;E�Ͻ��(��X�7p"¸�>�5�>.���W)w�/�)����q쀽M��t�W�t�7>�_�|�h��*
���U��T��mV�c�����o���e�_^��NB~�x����Tx�3�w>�[�����zy�F3?"�������<;n"�Q��^+exڍ�Qա7��P��\�{��ts�����[���P�ޔ�ؾ��k����R\��v_�S�ep��^Rxc��*�⳦�I ���lww���#�K�f��30���A���wN�TX���*��o�^N� =�4,Ӝ���t���CrR#v�������5���Hأ��l�T���{/��u���	��C1-��ͪD��>�i�%���	cԝ$|3��y&�cHͮk1��t���]!9�����"b�x����@zo��E>��z_�v@�x^IiM}R�;n��U��VMC�gz���ə��~���Q9U^�͆6�6�w��%ǉ�����V���-'<��Z?W<���F��Uޭ�m{���Up�x�i7ωyw5�����o���#���͉-m밽�T���fk�>��Y������|�~���y&���%���M6�������jRC�㲆���+�û��3Q���V��	�z�8�|��{��]��
�2FL窱=2��a�=��g=�.#+�X�٭7���u0-M2D%�"w5�v���\�mr��j}7�B����?��vk���W��A���k�j׵��&���uH��y��r��'.�)eگ^_�7�9ǹ:�ވN��~k����%���xY�������ig协�[�|r��};z�^P;�z��No����������*����3c������!����o�#�ߔ�g-�����ĳz ��[N���zF�':�I�:�6gp��;��A���S�jVC@r��]ʱm5ϧ%j+�!�Z���{+7�`.��l"5���l�B�˖�`�Sn���|��A�)��eQ,��j��&�������Z쮑�K���ּ;*M�3y!�F��7�3o��z:��0ˬ̫������������J�O+�2��㑩�yq�EՆ�l.��\���3F��)��wr�]�C.Y�؝	�{F�2e %�*���B�,�r��(�B4fĺ��?�%�{vU̪�dqڂ�B��۳�z������ZG��yטkh���s��[<ʊ�,p�)��Dr3n��*�W�� �l�BDLԶP�k�Uu��薞�/#��瀹ltQ�uf�h��4�m\�q<�=6�Y�Ҭ�m���u�i��T��;w��9ZX�k)o.u�u(P�/�q�@���O~��e�MgS�ӗ%"/$�Y@os�����c�]�!�f�H�t;\l�<�D����Տ���;�ij�S5-�ΰU	@�ۼ`��Bȹ�ӧ�^4.���R��a�����������2옓�N�|���;�S�:���|��82��W���"ۋ&YOr=6Y9��B]�O�J^>7Zx���]��K޺���+LT;d���u�����/c��X��YΠ���;	�o�u5L�պ���ޣ�^c&�g��mh������m8�X�s�;+����Ɛ�k�Q�y�q��'uv�ξ���I�V�T�VC�e�d]��Ύ�먲�l
u���VQe�ǔ)�;J�^�pj�� �|�x���
ɵ�*w*y2۠�x���]�6�k9|��9Ý��޵l�c�.J�{��yr���iS	��%�R�[��.���zkJ$n�TҎ�O�,bp.ٯr�=+je�Z��a*���2%r�M7gRX�j�'��(K�s��<R G��Vreٛ��ܧ_�N��@Yxq�4�>g�����
�<ym��&�T�׮��,�3���39��að�9w2�*��9�(� ��o�>��ۆm��O	�)�������ycq]�f;,iS��ƎRu�v�f�v�t+��t��X/�;sg.�oBG�9W���ZS�7�(;_,�����]G��jY�oc�(�w���+��ӕY�fXF��@9oix^_���]������խt�o{��Ը%s#t�� ��c�⪛��#�o�Y�S�/�/(@�b��Z�d���v�KF�E�e�B�cx�7[����wZ���:��{�S����o1�Nh�B���9�m�������gc{���o�	՘z+��4�α�4Q�Pl�P7r�Hk�l�	[��78��ǮBBW�^N�����r�:qhYԣ۴�}�[��*�4\=\�cYNCx�<�;"L�,NR2�m]�������2*�=���x����y:I��xh�;���H�7E<��)ʤ�"�
�����@��3�3�<(jTJ�$UF�jfBx�U��ExZ�QT\�"�lfyI�^UE�-db��S<"�4�<����Xj��W�QRJ5�(�j1	2�<�<�"�h�'VE�hq)�8{�j�PUz�Z	
�r���c<����!^��T���QE���$�����xQ�W1C.K�TZ��Yy*QWQ�Ib�A�T�UTyAI3&ITP���E�U陇R�^L(�����"�R<�3p��*)7x��IIYj+o<o=�R*W��������+��AJ��zbF!DUQ��&HE�2���f��F�����z��dQxy�yܨ�H�Vs/'+��9�xy䞞���DQ� �f��1ug��C�tC����:��ҳ�Z���{���<-�7����ӻ.8�u�)S�L���VK��[�����}o�!<C�(�������G9���ν�!�_�Gm���z�;!�,��@�W����^;9���w�Y^:f��N�+떋g>ږ=w�h{"�3�#�.9����w�n�>�b�Xr6_?�N��Z�+�?V���w����L�Q8�Ŵ¥�؄��,8�	���O�:=Gݕ}��R����o�r1T����r�-�'�7qR��W�a�Z>̍�j�ݤdW�My{�Ui�̮��^�s=~l�WR�{���u#}��y�G�� '�R�_W��Ĵw|k�0k=�������V��A����ʕ�rxp�~ ;�۷ U�d��:/�L�$NEfp�J��^���b���ExGt���5�������#�:Ϥ㭠���[���9�UCG�;<}�8�/���dM����K��к�vV��_�Tr�p�����.1���9�� ���BL�Rվټ�Y>J��I�>���g�uo���댟�Z�A���=\��b������zD*�xz�u\���תVuV��ӑ�ka��A����>Gz'�=�[�l�OGzx�� ����w�f�F\��K_������z���K�^t��ٮ7ʚ+��x^syO��Z	3��!0�ov<zo^^5��#R��]�kA��F!��l�.�����^��u�X��1��y:V��o|�[�2�B8��5u��ӆ>�t�!Z�����aŪ���Ԛ`�=���~����##۵���I�ꢎ��vw��T<ٜ8��Yp3�\�����ub��!��X����p��,����g\�~�Z/�h��L�xvvX̝�P�����R���G����>�>\�P3s�`U�Y�տ?\r7ڮ'ݔx��t�s���l����{s���]���7�k
���1z�'7�G���<z_�ivq��W>��(�Pw���Ȣf-����:
{����&̓ު�&.y�/&u�ɟ"�̆�O�tg�����~�#&� r�`�v'�W;ki��G^m1�}Lܛ�e��T� U�S/6�����3�٢��W/�5�����{8y�mJ�Hx#a�>�z��o�Pnj	�n���J�u��������M{q�[�Jq�Լs�p�g��#E?_��!N�e���J��Q���%�@ǠXgtϳם��:ښį����.�~7�Tm��$mϪx�;�	�Q����2����ѿ���������7�l{dvz��C�vu����s#e���Ҹ�u�����(�C��/�u"�˒G����ݗ�^��u�!*,^��g?o����Xl��/>�	-����Py��t"~\@��R@�f���Z�X*Z�]�|k e5J櫚���ۦ��k9˳��������.=+�q��;+��tKv˸�}�����P�;5{n����|�	���FiĩQ܉��5�4W�ba�}tɯ���Ҵ�@/o/[��;�����=���Ɋ,���X�����k:;�c���*6#�7Q���1�MVѽs�ݐ%��Ud�pߪ�}t�2�]꼯;��B�Lb�uN��. ��@�Uyț�{q��a����5���_W���ަ�ۆ5wm�ʯ]�����g+���� �u!��G��,�僂?�_ET0��&��i=�����疮����&}Q��w�-��T|E暑���n���M��!%��TB�s��X��Cm�Т��0n�����BUZoJ�o�b��#��s[�O*�/ٕ�Tp�zI=�z�3��=j2�����QҶR���\2�kO_�>��\����w~�^�O�;�G{U�������G�ˣ��ۨ�+�k�^����6s�X�FMib�&w���令{s����^���N��9�nϗ�#ޑ�����~V����-�������~5���2gY�|]N�v׽F;o�{>�V�������>֩����W/-��C�ȕ.M��桁]ꇱ�S=TO�uK�����Nu7֘�9DZP��JJ�����Ձ�X�Z��89�6�����q�� ��o]e�.�F�foc[[k��d��\����p��;����R��*�����3;�ycI���L��Kq�Z"w��9αC0j�-��Q�]�;O�u�p��iБZ��lx\�V�����;�<ٸ��~eU��]]�]�v�������[M�f�#�ʣ��M��t�W��/���=~�Z� 6C�p{j}:O��̡�����l��ET��t�M��w#e�V��o�ٌ��v�v#�i�S�i8�	��'�뗺�I��1-0P��R��+�a��x�}�୪By�w��(��c/�
������k�ȫ�����EE�F�1̯��A��T����W�����c��t�����y������O�V"o<�������bە)ύ@Q*�S�2�__�����7���{��Lz1M5wF�m����M�{��/�}5�~�P��Mh\{�`M[��M�Ux-�6��!��u�^�G���w��)����0�>�q��k���|�f��=�C���h�Qs��r�9W����}���=�G�/>�
�u���^�&�K�Ż��:��pq��������s�4�����������Dc�n~�"ɾq�Z=y:+M���Dm0�\xo��|��O��ط��꺙�/�:��٘jL%��-���Ax��ģ�/�xb��QҤoz��s:��;���srl�t%ևܓ���.�ң�[����'�e�㞶�}iU��poVli�]*�N9���/-��O�h���CW/;�f5�5�Wnl���0�vʫ�r
�`�W{1�@��m$wv����׶t�ǐ�}$��;P��+�X�٭7���Sb��2�c�yt�ٞ�}Q&|�:��:CEǻEh�=�s�'���xk+j�i~�A~˷�ܧ+˗�+���Iv٫叅��U�����v���/e!���R�G�6�+uFx~�n��ԛ�����Sܽ�;|�����s>��cm�_��o�?.��q�����x�:����`�U�8�Uؙ�O�5��:sy�/uü��L\d�^9�h;���s��~-����1�s�,�ŭ�T������ ^�������$�����rJ�nпJ�3�=
V���ƽ:�÷G����|4����Uz��L<��5���#�-�M�a^/si�o��Gy��U���O��~�6���H�/_�<1N��<��!���P�UHB���Xr	h�3j� =�-���MM�}y�����,>�2=�n�:}��y�<��r7�r�G��)�@of�Т����y��r����ڭ]�r�\o}c���J�o�]~����R��� �۷"�˒7�:-�&m�PQ�gO��FoZ���Bv����Vح�u{ڒ�7�����&�a�p1Ttmga��G�n0�o(̌�Nq�F6���҉�I��0{�F��ы�7.��+-��qL���Z�X�-]\B�;6[�a�{=�l�%Of���8I��Ժ@���G���˧�����ωxj9x�z���ߎo���I������]I㛰�o*����V>j������*!���"��;����b��>51�?:S��`{'!8-B��~��[��Z))� }���+]O�쉺��[��}���k�s��F��SD�_s������u�W�%<�*}��c��x��"�� k���L��-lW�{�	�K*�����oscU^_�*��J�6�Ι<G�����/�=����2x❨xn���I�����#�\J��{'��\w��s� ��b�7��Dw�;�ꑱ�h�����+ftf���cc�禽��z��z��;:<9�>���s�-9����F��\M������;�(��x}/�{�L�tZ�Y��W��XgO�#&uLk!9Q�|v�����Ϗq����FŊ�3}�S�;�ݼ�Qg��[:J����z���s�,^L�73�^s��O�td{μ�^�B�������"fAS~�>�θ�k����tU3rm7T���D
�Jnsjaz�i�bTT�׼���JˑG<��ɴ5& {�6�z ��*帷��L!I2�Eç*ZV���=��X�V���kkEEd�OcWI�b���+Z�Ԓ��V���:�6��g\4��
ΜJ��Y}t�)�]�3ޒw
9}QΩ�u>�������0NҏŴ�m^�N��;(����#})��7�=���Pnj	�)��^.�z�l}S
���R����Ѷ}O�����އ�F��z�~��2�4�nn	��ё�`N}kn{;g_�_�l�}�PѶ�D�νi��(�s�'ED_�܋�ު����@l������}�n�xwN������EmP�*S9�Ndl����R��M����_���ۗ"�+u��/T���{��c�=��Keg�ڋVDӞ��<V�X���C�����U�X��\�,���rNyK�ߟM�����Ț��R@*�ޛ�{y^&&)��7��{>��į$�A�K�����!_�kw:��3��U	ٴP�����m��U�{>��{q��a�Fz�MF����ز�����Y��;y�}�ǡ;5ý2|z��j����H�1%��W��3c�o7j%����u��uK����G�2�3[P٦�/�#��>#"�9~۸���8j<��s�$,<��es�}��]���_/h~��G�'kf��/Ǥ�`m��G�3� .S�n7۷q�m�+������+UR@���*�F2����C 9����'ӱt�0��8JWS�~���q��_:��T�: �v��3"��X��1N���v7�ޫD���.sou�S}%��1]�-�C1������6�����x�<#$Bc�)�a-u�OMs���Wغ*z�r-���G&u�"���q[���(��ޕ�dL�8϶���g��2kJ��8v5��M�Kms�>�J!�_���|�g�QU6{q�]�5�^���1���}$�Je�Q�ZX���� k�#ٱ�m�7{�l9��P�����,�7>h�t��B�����Q��%�E��6���خ���gY�|�^O�w��������1~����������������=.M����yU��^G�ftELc�q~I��{ǽ|x������χ:���Ke����p����ȅ;E���	j �l�C^w}�Vg�oO��x�C�r��͚�~W^��~T|Z;���~����ʙ0���9��~9�
�_��>��۪��]y��3�e�Qm_	�o�ُ ��~�#b"ڰRr��zO��^ru��h<�7�c�'�|'Պ�CKoYd��S��gK
�xe*�g��SZǼ{�q
�8�������ʨ��!�5
��#fn"����	h���=�b�F���yҬ�랼�d�����N��� S�hG�r$[���*�S���M_��9�G~M?Vq�+I���گwgH;4M����c�!r%���n]��ݏ��+�u;e�ŀ�ꕴ��vٙ9��h0 �����kz�Iv3Q�;��m�w�ZC�`rx\V��k;/�e��d:V'���%=+�E�'g������_kL߆}S^7�T���t?m�W�i�D��>�͆:�`����p[���L�qy�!wJ��+K�q��k���q��l��<�}�σ�$�yω{|�r�3�
��uu�pJ[���r��ٵ���g�|4��i~5�,ˇ����c<�N�~�c��T���CYuأ�t|Y�?�QZs�T�ǲz�����:'�k���}������=p./Nx�֞��������n&
��*}�V'�(����3�G�E��r����*��3��>�`;/ux gzd�(�nJkӤ}��N����g����Bply���8ug�P��V�;���u���Ջ!6cgŀ�ܭb�9��
�GT�6���7�<{������^�C�yp�.�{&pa鿨����	����z�!����/�q�F�����cm�_��o�������>x�G��P������nV�U��ڵ�\�%�р�}U�[u߲e9������BN�Ws�i_x��"/��7+���G���ת��Kٓ~:Vt�,� v{�1SȊ��-��ږ=q�Z�����pT����懗�/�1Qy���kJ��:�OI�n,�����Gӻ���vi���yt���[��'a�a̞R��>CP�6�.�k^s��r��M�/�Fp�h��XNS��S=;�������a��R�Ĺ��)=��o)$C�~�}2���c��OU�IEO���.R����>�s�c;G�;\K�����R=Q2�D�a^s��l��7�	���ڽN�n|'f�Vr��biy�9;�x�~���:�ǲ4�nl���HB���X@h��_�xl��U����_j�>��&��E�t�ϟ��/#�u�¢�n���.ƙspH�n���l,�F�]��үn�;-v��Z b9��Ly��Ҹ�t�zN}�ԁyՠq�DO�꜑�#��DL(��F�n�cγ'�Ǹ/C�"~�+N�@>��9�5�ƣ��+��γ�8�hp����^�yn��*��;z���MG#ƥ��Dz�V�����,m�p�!϶�.��!O������n�g\ׂ��'����3#^�֣�d�y��ׇI��s����4K
�e�.���n{���^m)����@��/M�@{d^@J��>Gzz��q��a�Fm{�x�2�9�������n�@D_v<��G�\l�.��f	�N�$�Ι�t�ó~ن��;bsʬ�Jzw�s�}�zn:��:!/V�����g\�������t�䈖UUm�Ag�96�׌G��.�%	��O;+U��p�hۅ���}����'H��`z�ⲧRc{Wm��mav\�+��}Jܝ���Ԓ�-���a��m���.�/]�#��dY��XLz%rO9wY���$���@m�ojZ��P�Z�����7�\/������Vaב/]�EzQ�Z��_J���P�|t�9J��I��W���,t�ĂwéE�u��a"�u V&��o��_<2�uu,W���1���c�ʵ�op�{ݧ6��W"�l��93��=���TgtU�lG�u<��{ӟS�j��:�V8 �y�N���{c:����W]��ޚ�x���(�����\{��;D�eЬ̛\;b��6��A��_*s4��ZY�_0@�E$ɳu`�ц�/�HU8����7�U�hJ���;�]�p�9��E����hۗfmvV��&��N�{F�F�!]�Y��[��Y �iU�֍�	oWt+8b,I�4�ls��;!%�-��8sC*nяX��GycW\�Cv?,j��3-���2�S)�G��fZ��*��� �'S]Z�t�h��)_����Leui�|嗧Hl|v���anu�r8u��8r|��
�ՙ#qMȨh.k���A���3��_N4Dm���N�حЂ� �#>Jb�����}�Nժ��Ӻ���lv�ɍ�T�A���.����W;u>�l�l�����W�$�t�$ �+�͉�6���w#�e02��&(�S�e΋��{`�y��ѐG�^�ɷ�"����e�΄��u9|����f�3�.Vv,`�'F���P�6l,Kf�
|�ų,sT�_�C���v��K���v��� U��7wj�ut��n��t5l�1|V�� ��mI׬������9�A�k� ��)�B���$�m�TӭJ�W�f��X����&"�C���hԳSa���Y�ہ��ќ�)�r�o:Z���)��)���q��^|����%P���RBľ���=�� �ׇ�H��p��i����~}�m���Nz�ܱr)�M�S3�t�ү�=��B�O,�yt� i�Lzl�͔�*|TN�v\���TԒ�K�M��h����T*��G�+Y2q�][Vc�������:L���#��!�p��;�R�x�F�a�b���I!lŰu�i��;��;��h��*��i�.ڎ�0,\4|�b�b�20v]X�3�w¥ڝ�u��y\f-��^c|��=��U3 ��V�6���1e�K+8϶��ޝ�Y���W�g�z�8�tNҡQ�+�mi���"�<����W�n��R�݄������o�[f������`#����V��(	��Z]s��}y�3�b�*�J�--�6"��L���BQ���AQTD���t�9�
��Ȉ�#[U*<�=<��1r�Lj�B(�$��������I*���>�yL-�Ł�_-/<���T�yI#7"��	I�A3(��𝝻hDMr�sD� �ȏ���"� �h�7"���Țv�����o{�$|ܝE�ޡL�(""yⓤ�����nu��뗈O7v��w7�>�sEP�+ʏ(fE�1�ݵ�L��M��B��B�S�*<��US��ݮ�-)����L�*P��ՒX���iE��(��<ʨ�9��J��di+�]�PQ�,>���s�QPE��k��I�Fr`Eg�R�z	��\�"�%U���C�xW9�<��J�*I"�v5����$��}}/��S��|��ݥ��Il���U:}��us	��]a��_ay|h�:�u:BZ�I:��R��%�9˗��:ۏa�ﴸ�|}s��n'{⫡�㑿�Uy�Tv5���Bf���Yϧgw^�����cY	��#����W��~=�oӼpǢ�ً�x�=��`�����gN��_YG�p�ʜ��*���x���=�L��d4:}�X�7�n֑��O�ۥ=o�
���Ҳ����㼤�ƯlU#rm�7T��ȁ�~��٘^��PϮD�Ϸ^nI�c��3���z3\JG���Ļ�G���P���(�a�Ȧ�W`��wb�^mnU�糎עG�k�X��-�[/�%���4W����*r�-@!��x����`)+���{���};A��`^��@����mCF��W:��r����p��_�܋���%��?=��Dѫ�r{;��-�`m�A����*��7����l�iTN������%��O�;��w@Y�튃}62_n��r�m"@�J%��10��,����r���C��~�u{�;X�M�)�h��]^y�ϣ�t���[���/�Q-50�c+��5;Guχt/�CCO*ɿ^ʏY� �,g�!T�afDƬ���;*�G`}���J��݈��.�G��j�['����7U����T�R-��&�S+�h�i1�R�HX�h��Ԅ�9b���n�L+�u���}o*R��r{�۔��=ە��c��$���V�U6�*�#��8��=H)�l������y�ĝ���
�;�EUy50�r�L;��t�����7E �w����9^��p�Q�f���T|n!��Ľ��/E_y�(�Ǫ�d��7���Q;P��o$r}��q�+��ڏx�y��ꏈ�KOC�vd{b��!%=���#(���^��x��t�~�U�^N�Ώl�Ip&#�z�����q��7��v�[wC���Q���ڮ��>ݙ�g�x�=�}���%,�ʴ���_��3�g���,������t���'�V��%���nמ;��7���w�~��.<�Wq�T�:�*���&��q�;�q�@��G���:�eϣ����y�<�t�'ډt�w�8?e�y��YF-�l��z���b�b�gY���= z �J��N��R�|�t#�w�;�>G\E����C!��~�ç���F�):���VP���۽�O;�g�E�F|�������yp�O;��^���o��/�J�.�^D{�6+=3��z�٪�����ӕ������=^w�|�/#f�F�9�\{ /Sg#�%��=���O���2�+�ފs㱕�kM��efa�y���ל7��
=���Xݫ����բ^F��:V���`FS>9Ԇ�z�Mԭ\�]ÏJ��?��cw+5�a��ܭ�{�9_QL*���1u]�b!�j���E6��n�۶W7\_j�7mJi���#�]�WTg����1�s���w�UHu.�&��c��F�a�v�C�����D3�K3;?eq�k�����Ś�}/�:8�,(ɉhق�۪Tk�W�Å��̍�QmZ@�L����2�.w�K5����=��>�F�����3p��'̈<�D�}O��r	h�����2�ދ��RȪ]���:�7���U�>��{n���nsbd��\�)~�>�K������T|�#݂c�j!&k��S^*#��,�5�p��[�\�r*��tbΨ�"������ns������u���5��i����_r�P�7���ȇ�P��̱����&�'�x��Y��OZۚJ�I9~��a��r��ٵ�ד�3Q�ƙ��,z�噐�̟L(�8���Z���yZ㼪�v��:|�Gd�>��,�9��x���7�'t����Zn5��f��	_�<h[�o��0�Y܏L��mu��>~�7��1_?0+��l�ɇ}^����i�� o���g�n��@Ϋ�α����ܚD}�[m���w������Z/�=�s�'��vw+j�k�/�a��������o��:ja��Z�rd=Jh�K�̬�[ �G5ܩD�N9���-�VJ�n��Me�7���]k��+�
��f\�Pe�c�49����8��ҳ��8�oݔ���W6�]��eH�R����/1��߽DzfG�Gz�5�����h�{�p�5��}�%�'����p7������7�9�ބ���L����/��cm�_���Z������-��{)���K�`U�5ޞ���!s��~k�f��x���;ɔ�.2g�ӑ�h;��߸�x��"/��]�U� Ϸ�R���lף/v�=��3s�۪`O�<����-���c�����
|Ή^��H<-ј�9��jtﯺmLe
��3��}���#�Y��qN��Rۈ���l�V{�<�i��{e�������Ϊ��#я�����8���O��S�7>�!��T�R�^������Y�y��}��7�U���H�s�H�~�@��Y*/��G�>5i��6H	�tly�ҁ�>��Dz�]��7�=wiaȂ|��~=&���κ�����V|߱ =��Z*-�9"�&��t����^���Ѭ2��LV�������_������.�����o�L珤⭠���b�S���Go���5���ꄎ��u��#�+L��;���,e}�\;����:�(�%���\��^�욵�Y�F\�1��(��Zָ:�g`xl���n�q��.��e����L�l����h���-��)�El�ʅ�H�L�5��\�Y�Cd�څ^���mv�{<[�\�V&�HZ�!INL��`��W�#���&�T�Fd8����x	x�#uW7]�:���?��v�ಀ����#��k��Qײ[�>�Z�5�y`*��c��d�*���YQ}Y�~ʧv�
�a,5!T.#���>��A����z��E�k�XЯO���f����qS����,���}�ϣ� '�j���T|E禎���bG�	���$���QGo�ڇ��	�w�����ah�g{�˦p�4��OK R�v�W�|F}��gz�\?h�{G�f�$�E������>�Hg��>�<2��#'������M�@ڌ�`W֝g�V���#/j��W�<+���H���wO������y���t�X;)�v�J�����	��q��~�q޷���{��MU{ӕ�39���̩�N�|�z�dG*(��d�rrp���\���:��Z�uA���{����ە�y{�ekT���y�x�7>��ό/tL���h����T� T_�3��;#�����}w;�ލ�F��xX���ё�)���Gޭ�*��w�g�z���+��p3���ו����c��q%��<�[>����5[�\z����%���#E?_��"�^i�ܴ��lH����"H��؜1��V��Vҝ���_�o�<#w�v�W\�Z��p謿n{׋҆��)Z�$�-���x��<n݁�r���و.�>O[-�L��iY��k���l��Ɔ����e]��*ٕɞ�U�}Z��N�ͦ�͙E�0�GJktj����3��FF�KW�o%��ن���W|���ߏ��L���߳�#+yO:�e���̏cx_��Q��/�e��x쩑�ϑ���͗�VҸ���_�s�;ģ(UY���j��=�ր\:�r޽�/ݹr*-UzH��nyN�3N{�@�Xs�c9z�����x��l��c׻�q�׳J�ә�T����ϯ�u$���x�����11MVѿ�χu?
��r��nN_w��ĥ�SRxyy���ޗC�rN���ן� fg���7P��+t�~^*���+��*�u�J�յ�=��}R}�8�����j��W:��?z��jj����=�C�Q��W��9�E-�9x��7ӻ\V�-�.څf��q��3_mC��/Ü����0x���~�Dxꬹtz"��cy�]��e�����#��<&U_�J���>�)A�k9{c��x�q�tY�}���O<�y�β��>kl�M�%q��Cnv��ɭ*�2|+M�k��������{��������TTq*���V~u~+��?Wv�7�{U������;����ՑLed֖/&w�Y����=�Zj�� F�K:�[V�*t�낕�b��1Zuh+wG(��x�Տ5C�\��U�V�(��q���r�:��ǽsr���D��ksj��\J�������C�Q�A�g`F��kU>!X�l��7���o,�]g
�N��w �1}��c�WV�j��)v6���E��#�87����]e�{��9'0�����_b�aV�a�Dɨ3^�lўi6��̱�Ω����r7μ�m���/-��C��f��a)�!;�$=�Ρ��c����_�g���ax�Sˇ��{No����o�G������z���j�}j���E�.���7�b���'-F����~W��H�{d����>����3�t�xc�<�_��qwd28��d�w��o%�3�,*�j�K~��?j��tj'����Sa{��N�U���,f�Kd@A����3������X#7�����fV�J��rk�'�>�#��\���t���\W�f�g�1>f��R&'�}^���Σq/�ۻ�z�H���T�$|2#Ԫ�|rP)C���۹-ύ@�QMș�&ŭ�D�,d�^��q�Bݞ��ҙ��0��F%�~ί�=.��R������Y5�37�!z::�w�'n>��s��r�x/�Q��Miz}F��\�T;��6n��q�V�W^G�g��s�z�n(徐���i���u�|i�h�	}���®�d!A�8��7Wk7+�
�v!���;��{o@�H`V�$�7&�=׊��=]:hd��Ǒ3��G�����a���|^� �&T�.��c��;!-S�o�z�Y=�sL.9r��Fmhw;�:X�3�X�G,̇��ݟL5ݙ� r}���Vn<o����:*=��#ʫ�\%F�{��^���O�=?��d�\d�%�?�f���Eq�eo���Z���Mnq?�V�1�V���ަT�o��M��gL_�뼌ۃ�5�kȭ������G���F�����7{�*�4������p�י=�W�j��я���!����&�]U
���uP<0E[X�i�u���j������ᷜ�F��������8g��{�Y��g�O@����o��ʥ�=�J�QATc��^L뛌>�����cZ>�aQ�/��S�|��y��U�Y���];n�$6�P��ћ@W�����}�q�)�\FL�zy�u�9�����?TN�Gf�Y����{96W�=��w���]e������ -�`g�<���|�g#jX���h{�]C�6
�~���7=�eH*\}ޟq��~��ʜ��=q.��9\ET�TL�@��)���ğS�.�q�w�W�W�Vċ��������H���ó�U�P��2�'�=�������4yp�v�����*��T�j@�K[�����uq]X=٘��CG��]&wz�̄�P�7JUq'�z��헗�<��wf�R���H����Ğ���iN�{��|'��LӘ | '��Yˆ�9Q<�Y���V�ȏ���r�n��{�o�	�ٙ�o���|?%O�{ƣ)#�ϥ"�~�@���Y!�m��gޟ�xdyM�sؘ�M<�ٛ����qO�f���@b�D���ި��u���'�J����r5�{���18�{��ߔ����s���Z�)�Ӑ�aD�5��n=�U^7-�I��`����T��Lͽ}N���j��b۩"�Ly����I�ZdV�����V.��5�k�\�^8ع�ȥX+���T��H}>���Xy@Ty�zJ��S�{"n���n��ä���g}��>�̝��&֤]��h���X�FDy�=4�4�� �� %a�T�j�m�a����A�fg0Y��Q��޴R(�m ������T|F�Y;���bE������=2Q���Y��^�w�s���ш�亡�ٵZo�>�龦 �N��Kվ#'�p8�޿T�y	��"�}�%��<+0ٿfV�[٧�i9�e+^+u���Zug��u��-���z�ٔ�3K+A7Z)��盗��k���~����27Mҵ`��~v�KK=1z�'7�G���<���*�H�U�~\M���w��;jsc2���T1�n.)l�y�eo&�zdW��ln�N�j�qP�u'����c2�>�j�2�>CN����/��� /�=+,/���o�BL����pwN��.DA�r��\ȼ��N���3-�;�"(�
������|"�{�^ב��E��[+蜜�*�s�,^L�7�>E�ɅB:i^���᫶�+�+н^G�7>gr/��7�\nC�Y�n"M��e�'�Pc[��W���X�V^������k�)���Ѿ������yh1��C�����f���6�^�Β'3�-��Z��@��+�S̺ͨh�n?,�k>�x��Cw��ޯW���}�;=�T]�f��hp�_�\���7f����@�KGۛPѯ��q6�֑��(�s�'B>}'{��6�U���9ސ=��w�@�73���g���,-9���j�Wq��I~���/՗��g=�w�O�d�4����DO�����?(�x�0�"f"������ZZ��M���~Ud=�I�O,�;?����s��3�9w��q5nk�@����S.|Lw��m���t�F�LNr򵗷��3�3��z���~���P��^��� W�|i�qU^�"n��R����Xö�tIK�ʌ%Ҥ�#J����4%FX��T|o��@yg�j������1%߾���U-O�7�Jw��:*&�1w%����#2�Ýλy����d�$��B��Ю�ۜ�J����������9n��0u�.���#�(ꬱ����*s�һ�f��o�k�s�hR�a�C����3V��U��nX.Hw
'B��cټ��nn��w\h�]�F�ٮ*���rg|Ħ9�ۺkn���D��/��uX7k��(p��X��b��� m�A���آ�V#��oX]: �Ew6�ƕo=�1	�I�a���8��U��rK3�ÙZ��Z���Q��op4ٕw��58
������;�S���N_ϤIj������z%D��V\�Eԡ�HJ�7 �y�r�9�}gC|x�X_$(޴s�l�8&.�ں��>��7���ap���s�G����Nԅ�:�Hq����Lz�v���l�1]��I��{�� �f5���a����D�f�s
���/pȎ.��,v�"\ݝT�%AV�m^nvfl�I�!:�����o�h�b�%f&�ܾX��^P}���ε²���Vm�uf-��:9u2n��&���솒[WwW�ō�e=�ٱ�ElZv��5�p�󯷹kh��W3����Q6���Am�^ջ��$�Z�tHu�u��A�3����{1���qǻ�%c�ؘ�i(�]�$nj 2O�%�3�3gI�p��%f��&���Q�Wj;�N�C�R����5 *̗wǲS%U�RY�t�'2n�k�na�9(�x���T����s׉��iѳ��H��ik.c��C������G��nv�)9���ޞ�;��}���y^]�9��k��Y(��&��U�u�;�D�֘�;����Hvt��U1�ߠg�B����N0�-�k�󭽠�+����4�i.����
U;��>��C�r:\gQW�Al�{����c��F<j��;�j�����.���q���JU3br+Xw:���+� P�B���V-�������X�ڵo{�*�fe�0/FZ8W.H]j�� ,��ׂ�z�t�9�R��lh�(���Ʋ񭗅��`�ѕ1�W�}S����h �&�.�`��UgTszS=We�s���J����9��U�N�g= _|���.����Y���;����],��4^�N�iˀ��}�c�j��܀�!��oh�w7m���.cA+/��ҽ�v�;��C��O�m������]�N���o[�\�i־�ܻxfd� d*k�K��P�c��1��y���et&��i#Թ �ReM5�/��8Ԓ�V�3��ŲP��V�'D��>8Pp;��9�z)/6��3���Y4�s7'%����
WR�R���)�K�$�YŃ��X��&����#Ď�ŐJ&%3�5�Fh��;���ɷqi����fƴdM�ն��jt}E�16����+x��vMŴ�Ev4�p��{yBgP��`��?�{�Slxs���P���t�w�թ�\d���J��f�M���B�F�7˵՝\�yݜ�d� ��R�e��j$��H&$!x�Z*�9̙�9�B-�G�4\�R*�Ժ��J�j�Ȩ�U&I�e�dh2���\���$��<�jS!v�'�Q�$UUQ�A�fz���EFKY%�`A{��l��Q��Uy�K�B��۰$��!�5/
�R(�2
��J�nZ	E],����=�h�Q�#&*Qma����+m�tH�&h��Y��،2IG73�<�p��kr��U�5ج�6؆J��yF.������NI�k2�Tk��E#k\��I����)F�d�ֻ"�c+#�y�.��y�z�"b���f2�򩱻*��W-<��\�ʨ��"�Lإ{��j^F���:�J5H&�d��u�I-��b4��s��嵌T�dȪ�$%u��	=)*Қƪ��VxR�` U I@�B�NV���-�sHW�٭�jK�7�=π��[\��ٸ�*8/S�^�I7��I4����#��K�wgzsS7�����s�V~����n�;�6��8���ڇ�P����uG�^���~��~��:����zg�H��I��x}�챗���+���Ǻg�b��#��s[�\m��W�$�e+��Gh���Q�̨�ym�7rON��P�6�v��3�Y�+�r7�|X~��=��k�*j����
ݥ�<���������aF1��z��K*���&��d����Ҙ��y��ī�~�ꐶ�֙"��#�����hvyu�b��l�vOlET?��G�-87�mo���� ��G}c��>�&XO>����s�|��߬�~��2<�����)�����Z�k&ֽH�'uל��/$�X���=q�S7�,/�uDu�9�l��~�ڦ.�Ò���!Ws���Ѯ3&Ǵ,�_������@���٠ѸI��Z��\{���ѕ������������۱�{W��5�WU#��D�d��w#e�_[W�|�5:Ga�>����u�Z|f/%��f=��3��:j�n��x�zK1-���$Y=�̆W��d���j�vtяf��7ÙrC&���2�Γ,���������pI�tZS��+�^	���6�:�P�����B��zK�Q��n��_ �^���S6��ޥ��|m@�����4%t�����waԱtc#�3j�>�b����N��#�9#��>�	�Wi�7�(����w�̃���'̈L�c*��j�a������t��s=|Bt���R���N�c�����D��^7��A��l^�E�w�)^Y�7��1��h����@�xk�k��=�W��@y3: T����~��ꛞ��j�a�s��*����C/$�tE��MF���o��Q��C���6_���3
�NQ�Z�~�]�3lb����Y/r"��n|6�kC͟	��cL�F�=\�2��]��M�J�۶�6�笹�މ:|��|=�6v�ǿIe���S�ǲz����>��tV�g�2+��b���Iټ���N[w��=��G�N�������Չ�~�:b��	�7�(���C̟qag>Q2��w�~���T�-�b>����@M��@�����N��pW�w�Б��8<�N�_z��Վ1��e�ү�Ot�{}����1�Y�� k�#�7��v�~;���뽗����H	$��O;_��q�/�L����(�:�Wq��&w�q��7�,m�ׯ�s��K�}^��>=���O�]�zo����]�����r�v3�͔��Q��/Ը>G{\^�y؏9�j��ZvOu$h�W������s�d���7F����"�4��0����3�7ݢ�'xwqx�"�'�=��]oO�-�Ȟڙ[�u5{}5[�9����ɦ�´L�+��[%t��z7����uN��@��T���\<%9�ɟ/NG9��s�q����,����oK��YgQ���n%*����e��%�*@[qT����EEϑl�=��q�׈���d��,���)�:2K�������Ǳ��vk�vn �m�U#�-�=�T��s����5�[�9ݴ��o��=�g��|�Dm��q�Ǚ��-����xc�7[Rrk՝�8�g�!��	���6���i�RE�e���#�_�܋�z�n�8�x2��ݏk=ѾO����4(���p���@�~5ɷ�9��~�y���^����;��哷��Ox��W��B/}0|Z�&���Ȁ_���^�^5��W�����hE!{k�LߴH�Sma�;9 .y@R�rG�T4xԱ���=ei���kó�X��EF��l��33<�����U��71�{�M��z�}���Itn�}�g�un#6�;�����R|vM��y���Y>�g�ZGz��.9����?:��zho� =�� %a��S�x�ǵ`�;���'Ϩo\�/ϐë�A��Wث��(�w�������
�r�L��� S�������Vu&띇��?4���g,�3Y	��OJM���oo_S�{�����BL�����Vz���u��}]������^�7)��V�ۧ+s�����p+k݆�����<�� JW���uG�\wz�+��Hh�Iӑ2|{9�u^-�~IS�z�����w�_�+��ڭ7}��q����v^��遦�n�Nװi��;�n�]�(�F��y�f�"�ۢ�~�ik5�~��Ǯ��?M�@��@Rs~*���O�F�ar=BǱ�>.k�:ns��#ϯ�ǲx迧����a�/rg}1z�'7�G�\O��"c�1o\JS�?��%�X�Q�� ��4���<��/N�S����0&�X�ɝgӋw�������u=����_���;����9�;�~�xܼWy��W�f��7T���z1^��fy�y���6Z8Lr�٥��A��ё蔏g����/-1N�q��P�ϯ�~Йx"r��R�u,����dEy���W��چ�}o�q���ϟ������~�_��^�BCgg={=��̝�Ӹޟ|J�7FG��n�7�����4j�W:��_�G��0c�Bo�kus��������˒�i�7����P�.|�@aa�/��m+��/K�^�ۻw)R���mK:�؆�:��)e-;���-Ʀ�.d�#ck���8����7�(^�rY�C��5������6	�/���gc3��F��'Y���)J*���yY����L�_x�9Wn	�R�?�E�yܠ��9��1�e�M-������������}�u���9 _�q>f�yN�3�tdJӮ,R�����"]�o��m��d������s�鋏NW�3����nD�E�� T�����Cܟ�<������^|�N��{Wz�����Ԫ�m������J�S�z��. �<�EUy�o�r�Dm����wN�r����[�㮓Q��}W^*��lbuG���z����+E��^L<Ǚ[�ތ���sIXXC:s�T��6��7j=q�^�|_5�Ż���uG�\F��<z��yHz��8�+���cW��K/�<o��Zo��c/Ӂ�L��,{�o�,	���\���}��2~)n��ճ9R^~ ~��֙X��n=�̒{Gޡ(m�N�q�ZU��V��r7�k}��z��A���ٴ.��^�y��K�:�\��{U�߻l���]�=Rp�ʦ2�&�� �a��y]~�3������}}R�u��.#9��+�օo�h{#�b����9��ő���E�W�ӛ��Ei���d���L���uH��޷��^g���x+����y�u�6���_~twqmL6��P����[��]�ūmr@K��:��m�i�f��Ҷ�C�mŠO�3��Śo��68�G�ʷ,�����ϖ�:is5!���}|��wYwCxc�r�yQ��E�E&�t\u�o�5eR���$�y�r���{�.ͩ�]O���M��pި{�L��2��ϒ������#Ų�"���Z�߽���N�ٙ�P�=�����΀��Q`M7p*�I��l�h�s���l��*�}�W=�[X��Jv��<΢��'����S�Yy���eHn*�x�h��c��l���x�Un���-o���/c�<�3�#��{#�E��Y1-�0X{2E��<�)�Z�*}��uU=W>�=ǃ��hM���C��s��9�F{2�,�.��3f
@y�R���D_�/�v˶��.�Zr	��w =P�$|3Ԫ�r����z��PG��&�Od�;��a�_�:*��}����ք�{�h�~;�a���=�*��=.���5���{������^�Ϧ��}�;�O���&ꩅ��y�C��ղkK��=���	�Q��l�y8;�|��g5������w| s>*]��xr97>y���FN��l�&Mic��7�'_�{j�h����2�b�W�z�z�����<m��G�=�f���,�9���=���u�֏^N��#y���tO��H:�N֎J&Fƭ���8�}�e��˹SA^��q
ī��Y��2:Gx%L���V�EK����;ֳ:��\PE�W;v�l�u:L|����]#zn��S��g�P5IHt�J��:%ꦹ����{MtJ�s/l��*}��;��NrG��>U�O_�l1��=p7�˕�ڱ7{�gL?0%iQ'ӳ�yE^��vvܸ��{���g������j��/佷�N�W}�$\G�Eh�= �E�Y���cq�Oc���9�P��1��h�} k�#�63��_v*��G�GTw����׫�Q��x����Q����~��g��%bΩ�3�ί��O�,���@L�L��z��Do����{��9/l��zvZ��Y�S~�������QEc�]�̈́\U0&��	Nbϧ�_9��oi����ܯnV%���8�"��-��7�Tm�VYY����n%Hn*�Sȋ>E��2m��K}�sG��ڝ�|��Y�ѾW����p\{G��������\z�Mc�5�;6z@[qU#�k�MC�6�Uĉw��Sي�x��l��mx*�~���y	\{#�DmC��#�!N��<�L��\�e.��w�{�����$`��^�Gֶ��X�#%��>�@��4W��W#�6��ʕ�V{ksfס�e���o��!���{fQ����9�ws�0�i4�&�u��=;\
+�=�f,�t��3R��~��&�~�����5�֬��YY��eD�R�jX�30��dӃ��t�=N�r���������7gL	�.�2�ԝ]V�Z�CnQۧ˶>y)��Y�8�>���}�sD���Td��4)5[������΢L�j�mh�p�#wnE_U9"�-�>Qj��s�w>��%�����x�i�k�՛9ڬ����*u�iH
����s�#b]CG�n���Q��ZdTF��5����ے��[Zgo<��g�݊�}�f���t�u;��y@9�*�]O��S.s�xz*k]��w-�
���(��ATr�'Ó���C����Cjڲ������|��U�0���[wEnti��j�c��i�f׸��=�� JW���uG�_��d����bE���;��6�9���R��G���mQGn'j�}P�6�N�㳦XB�v����O�l[��n/g{8�@j�ד^C�����x�:�1����ۅq��f��7���2��2ѥu~��{���V���>�*�G+�E~�Q>ܣ���7K���P��֗q�;��!9��*��׶k��u��r�h�����4���{~[E���l�`������5t��c�߭�kM�������握̾>�2�t��FG����������q��Y�{����6��	�%���ȝp$���gr�0�)@ݑ�\�}��\����V|��<�1X�mE�5��P儨R�e^F�V)�-��>�i]�|��ѥ;%����%G���b��I�W���_aL�	l���/q��?��2�3�f;?<�%�@���8U�˓y��vyp�5���@�9��*-�x�L�z�٥��~����ޯ���_�h�G�ç"�rtM���.�k}װ�^˺Y�� `������+��mCF�-��=�����,.ȏu���y{}tj�{��9K��p6��/�T8�y�A<ٿ���n�;�KGۑ��q�Tm���l�w��57~�}�Pu>,�>��f�\{o��#�>���Ѹ����FAs�s>��26_�uS���u��+댪YW^��Ӿ��s;ģ��x��n\��T��̈���Y�tND�N���27$��>f}��D�TF��o�*�1q�t�3��_�ۑ>�MT�5Ah���8�	)�uK�J��"c�IVѽR��} �e|�\��׊�K��9�@��x��y�h[k��o�f"c���[� �aڌ���q��f����:�4RVi��T|W�r����vS���ꜯp�u�d2=|$��2��3a��ڇy��<=�ƾo2�29���mEaU�Λެ���][`��3�en<��r��D-7;,e�p:�V�O��FUi���f��=�v�R4���I����M�OMj���5��0������L��g]c�{Ma���7���\��F�#�՚��u������U�:����b��r��g㠫�x���3���d<αֹ�bo�9��訮h�|0Ef��[vT٧�����Q�ʉ�yY�~rI�7�(m��1�3�w�>�ߠ9���y�{ϳvo�|*�G��,�V�私�����*���m�1~z+��I����ʞ�S�k��@��Z�2�׹��G��{n3��F7>��Z9�����V�pKg��_���gr3괳٤�UB㎧�c&u��&|Į�u���~9��;���땖����{�gspyU�uy���7�f��)T��U'_�T���K+�E�ax�u<�x9״���l�(@���ݼ;�W���U7��֏C�����P��l�`e7p*"����!����dyu�oQv}�ص����u��Ey�;�>G�j'���>��(�A���m�T�T�h��c����5f*f`G�U���k��zVĿz�0����{�騿[�u�>%�1-�0x=�����a��6,��V*�D�[��7��vW�dl�*�ڴ%˥�ǟJ.}g�UA^�n;<b|=�Ҭ�
k��y��v�y����XLLWu-9�wpL>S�X�SL�s��|����p[�H@�$��B!$�B!$��!	%H@�$��H�����I?̄BI�H@�$��� �@ ���I?��BI��@�$���I*B!$Ԑ�I?I�����I?I�����I?i���!$�H�������)��	gҀ���),����������0���� (� �JR��@((@�  T�J� �@B ��RBQP���R=b��QV��R�$J�R

�*�T�JP  ���ҩ%!A*U)U
��I
R�U)@�%R�'C��)HD�P!I);5*�Q� y'Ml��V֡� F�i��1�Ĕ��P͉J��QJ�i+lF@�U A  ��(��!����
JR�JR�{�  = ��pt�� Y׼�=+��2�f��X�D@ �p 䐠D$��kU6�ii����Fk"�ֈZمe5�5J%( � gR��(�E�kj�-6͖҅��V0%�j��Q�2���Q�Z��l�T�6���j�!QJR�  Gp5�SV�*kH֪V��Xm"�Kmckm�R�5+UlTڵ,-[[	1�٫J,��mQ&��I
"�� ʫ�m�`��M�SQUjS,�����ٶ�ݹrZ2�@��T�a�������mjf�Q*j�@�Ap �ڴkJ��eX��UML�+)��Q[j֘�R�kFl%6jL�*���mm�f��M�
aQT%@ (�  ��TYU�՚jfT��f̵M���SV���e0��STi�jʒ�e��Rd� [p  �Ҥ�Y��
����IU���٪������� ��M*��P�UP
RJ�  YsJ,�Cm����E�PUDV��Z4��R��z@  � "mR��4h2h�ɠ� �0��0�)U=Fbh�#�4`��C��L� �LL&4��)� �$�4�4��42�� H@����ʞ�2$�L#�bha���i	��       �m�9mZK��)[�����0���)x��Zu�+;R-zV��
|a&tP6?8�ATx�� �S� @��+��������G�@�� �5P	P�'��$�L���Q)
 �%�9���ε�~���ۿ !�����Y���g���VYJ"���?��!�yG+?gX+Ik+���V�T����w��Y����T{�7Y��zƲ�,n�)���av�ϓ�����a1j�Vc���L*���LZ�%��vv9XpnXJ*�K���)���l���4��ɬ;Y5�!�'V�[���l�/9��E�C.��f<����`�,����Y� ��f��0��JX� �6[5/HVr������
�
���]���j�fT�dϘ'��`��ɣfk$H:.�ͨEj����Îƒ�"�YO��|�chv�3m�Y�j�a����,�w�M�vr��4��Qh�:F�ǵpe��6S�KC:#�T�l�7Af�ka���(������W���P��e6�u)P{��ap��3`_�0Mr��EϮ�ޓ�Ňɕ4��1Zl���İ3Nn�kV�e�2����6��N�y����K�(X��yd����ZAdˡyZ�z�)��"�{Plml{X4*5��`��܎uVmTt�KbZlZ��9�ޅ.��Z�[2�x,8T���SfB(l�UƏe��vz�5���4�[$�jEJUl��ef!N#Ouڻ�ucxsa�
�@`Us�w�f��[5��	����(�e�D��Z���yD>�t������j�Q!�ly��It���,]�]n�?o$��e^�&��VΡd��alw)M��
��C�WX)]�" �̸)$ݭ�48e �ZD)�xB���nf�h5��<Lb�r��̂��j�m)qSЯ3r�=�Z觰�����A�HI���J���j^̳�"X�ܡ�Xɤ>5�L�]�A²��&e �VmS[.���#��b̚(�cq]��c"b[��A�Zh�م�f��ŵ��ŻM��:Ӛ�(��<�J5+J��Yj��Bٸ���V`l���R�=ib�(�M��t	��3ٵY���x�^V�mr�]:,�j�Y�:��J
��ͭ�nT�F!Z6�=˫r{�mbޫA�E�%Vp/8��nw>�vh��n���B��A[y�+�Z���+j�\���Vn̠U� 2�]�v�ɔ���oP���1[�(|o�����-��kpS�\r��e^%b��5F����I�o�F�l{4���(C��ȳV��U�c�*ˬ{z���D��Q"��[1V)�\��y�:��ՓE:*��Zs�4��zsZ�W�x�t:��p��ޚ,%���^]���­TN�Ѻt�1#��^��ZU�3]�@��
&��â���H[��;*�V���R�
�wU��*�ɢ�^P,�6`2�t���eܹ(�CXG�90��V�wt�/Mk=l��W�Bïk@��9��Wj�V�*

���03�@Z�YKf�ǻi;ө�wyi\wSH�r` �+�1���
�YYVv��8�p_"�
e�s�b�(�靺r7w�yy�J�2"B�LX���g+lL�M1�/4,��t����YX�˧����V�#��ed_5�A�L�&Asom�,�6U%���Ў��!���0l^���sq��k��uL�[vk�p	>X��(��<aK��
w���<Wɣv�;���s��l'�CghwǷV�c2����ƩҸu���o%[w"��H�EVKU�#sp��S�]9�<�\���_�]%Xmq�y͢6���W�Z��F�"�2iF��+Y�).�t��fnn���	WI��}!wS5	@%��J���X�;W
��ȯ���H*�: {JlJ��:��4>��f�d�@��hTL?�]�"���#��Hڂ!��s@��62D6��	�v�~7�T)h��ԉW*��7��Q���R���U�3wP��f��n����G+�[R�����=�n�����wn�[��I�*�i�5���O3�ȡ�+pB���^Y��^kMuun��/VD���M��wN��ُl��[�ȴ]���-\p�so6J��#�|h�L��Z���1Vb�w����UX���(St�!Z��Vel���R+h��"*�tl�S3*8&������;X�-'��a1V��^���LM݄��K�����(��b�!�(�-�8�l��QI�-���$�Y�&.O�=�պ�U=e��yI<f�ӲD7bQf�����V�}�Ɂ�1��XaS-�ئJ����	��S��ʙ�-�*]YӮ�3��ph�6U���$u������9X�YD`�o*
���"��`n���0ę�.�{NK�NS�7C4eKI!}�-C��4ow[�x�8�{^��Jԡ�jt�5����y���3Z�+8�'��|��5"0�f�q ؽ۬�ۛ���.��*{�a��x���T���p{���]��d40�0�	=zM��YR�8�H��{����/��T� 
��ڸ�_Ѷ0��թ�*0TQ�^V�sh��ӶAXA{O5�ڷpaN�Ы5��P<�[�)+�e��CUv�睟^��-�����E�i[��q��콫)��)GZ��
 �V�Ժ�K1GWQ��m��*�3lm�M:��6�[ba�jV	�^
ͣ)����ë�b��9��v���:ݑ�n��c0г7*�;��+�]YRԷ5M�Xͼ�4 �gJ���@��v&�Sr'��m����.lXiXK]��jB��Gv�{�%�|�	x��2p���ɳK[��n��A���ԧrѬ���
����Ww���(����0#JR�0�Z�x-��0�қW�ԗ�in�����N�p�� �ڷ�fXu�ګ6D�CZ8H{�3Q\��k�J�
��OU�Y���i���HR /2�ݖ2�,8�����B�"����Se����,<{I�a�7I�甹n���ZzV��\��v͔��s^<�c�]�j�3�V��O1��Y9�J��eJ�4eG4�LR{r=X#,��֡s��MbL)i֚%��VQ܌|�� ��V��t++�S�X�>�yXLʔ��)ܗ*�iҳ9h6,m��{Kh���j�"��Ʒ0XT�!�l,-J�݊���8 [CM9gv�yZr,{Cl��LZȵ��� ��d����~�ō_MV�B3���H�4l��J���=ʇr�0R�B�wW.Z�Z�k���f��=��բ�B�Ӂ��r��i]�N�[��N�4���4t%��2��h�������3J�>{�������N��j@�t5`�X���nއ�|�Ci�W%ؐ�|YV�Ѳ���F]��֛�w���7l	�{!�)z0m��M,t1yr�[b�\۩cu���D�a]�����-Z[�H��:�x෦�ƌ������ o-�����+�Oh�sz�6p�)=����lBЅG����d�L��d�:&��v�X�J�j�%�`'9n��j
6E�a���Ă�!6�1mm�oK��������l�m�a[ٽܣs5�5�K�Ӽ��.!�t�
���[Zˢ�h�����*ʸ;P\�)�#���y5�xn�Z�j[5��F�8N*�B��T�TJ���Y��̞w������>*6��)%�G����5�n�����=��
�7�l����Y;X�k��]51bX�ct�[��i�&��U�ۥ���H�(���#�7U�a��5���F�)R+4~�w��]�47k$CS�����t�L�7�+n�ǋoZY�D�m�U��o�0- y���e[�A�9z�Ҧ)�K_-V��v226ɪ5���4�;Oe=���L�ʚ�7+o6:ѳ^��+S����#R��zp�^H�-+5��VslɁ%`�i�.f�ni{N9a����h=�R^�Í��H��Z6_#3���$�oc��(��G3���M4�C�,�� �iy`8������Q�sF�&SCc�t�Im�SA�8�3����c3q��Ax-�ܭ��
8�W,����j�h��V�%u<YL�۳�aY!�m&�M����^ڼ�bߡ�Yy1��l:s,5�:^m똦�xm^f��YF��������T1�@�6Ƙ*��G*��	jf)��5h�Cn���l%'��σ�E�70ZQ�/�KZ�ڷR�6�L�7o4�w��n�l�U2 �����V%�`�гYT�Na��7nP�*�/E$v����9�7xrI�#�u�3�7^���a�:�T�D�t��s�=S*i���\X3.1�bB�Lֶf1yJ�BZ� �):���R��
�N7O+-�"�k^�u�՝ɫ-fS
���^��2��ln��^���@DU�v���zN�:F��}b�0�^�W��޻-�|/"��z#-�[��O�a��ۈ�e��d}y{d�-̗Q"�\��Ў�;l�k�(�Z�Q�7��� im� ��=g�������X���œ��ZK��O�4t#��qύ����c[X��sd]��f����Y�`Ӻ�kVD�i%Gd���'�h�(�9n��y�ڬrγ[���dz!j�f�W�ܥ/x�ΨľV�X7��Pн��ã�Ե)�k2f���g��*�?{�5X*�S�b-�DRR4ԃR�۰��q"S·R�n����wc]BO$;%;�Rܽmg%��o��[sb�`FN5f�B�{��JT ��^
A�D���NV�Ol��e��
jÊ��]>�r�w�a��n������ �o8���䉕�6�	�^��԰b�������u%��.��5%�0�RS�a9|nL���`j��,�����5�5z{�l��oZ��l�<����J���Bfy�\��!�P������2��;4��dF����GN��B��Y���3�A@����d��\�C	�}Vn�H�"Y<y�+q5��t�z�J�8N�N�I�9�W�>4�$�n�XDT�EDtv�.���n�`O_
���ô)3q�ٰ�}6�7}��_J&V���E�xF8������[W��,
��H��m�]�7j:�wy�*�����cq�[ǵ\�v�2�X�k��|z*{r�1�~�_h�m�C':�.�V�4eB�Y�t���3^�C��7������O:�� Z	o9dƏd�5�gl�(X3[Cs����x:��H���|���Z����s����U���3��Pu��faf��txe�!Z����S�oc��Sm
�'�q��j�Ec'���sH��=���=�c�Ɨ�i�N_cZ!�ɇ��]�j��t�%a��X�:��u���)@�$�phO�j)��9�Pv^�0�@�qg,�Γ�z
�Y�rc�"9�ٹ�o"�N&�\��q����Q�+.�ۺ-w]���J��p>��D&�)��L�7�1K/��;21Z��充����k������9�;H����V�<��7�H���9f�ޠ����v�ʚE 6��R(�0؟�a��i���]��-E7NVLLb����`�K�f�x��Y�kE;�'|4q����z8iw�rpEevr,-c��)�n��(VR��t{9!ǔ�u�<<O]!�,tx�Q!�K��Ǘ�2�뙻�����F2��b���|�P0+�VɾҒ���tQ�@v��;�v�w�\*��xu5�+]��ؚf�<?#r�v��B�սV�͵��=�6E�\�\[���į7w`����e��*0��#K~
ubo�#��Ƅ#�뽉��u��a>	
��֒��mrLu�K]�u�`�S"|>c�}T���̝5�yk��P{�媅�h��A����n��P���l&9f��R�j�IR�S����	:��\������b��U�%�́�=|t�ҹ���Ļ�����Z��d�/��5(F�ʂ�f�O����Uu���{`�=Mf�y�r�c�"r�ir����StX4���[�*�+��Ʀ�_8m��t�]	ӵ+#��Ҭ\:kXqհ�2����]}c�Ѹ[1�kot7Y�q`�����ʳ��8V��<�	������F�Ւا���7�Q��Y(TŶ�zo1�V���(�wƂ82�S���6=��ާ��!}�X�𴺝�UqwTkt�����x��Z.S��������a+i-q��#ӱ�Z�c+*�h��j��A�>Ō���*�Wd��5��0�|n���IjZ)���5f���S_|�A�v�185i}�]n�u"g7w��U8�3F�R�n�4��:�[9��@ɼ2�Xe�<�ɯ���*���}�mZ*�-D���S	�i�L�S�l�j��щkG:��c����i#�t��'WV��g��X�V��J���s)���ȸ$�9�%r�2�jT�0�pA}Շ,�gq���=�͎.8�v���\���IQ������e���!����b�s�i�Gb���4�cMne��b�*��{S�v� �f�ikͭ��h���CK&�[��7SЭ����y��H�MXkr9����լ��vܧ݅<��U�J�V� ���Y���S¬�lfӱ�r�MSnvTT�3U)&1.%RrR����}ok!��n��n��Ym⁙ʷ<m&� 룛Y�5���A
�kCpq���t�.m�!�Y�(i%��aK�wλ#�*5̛66_ҍ��,eZ�9	t14�sdݼ5�,�W"rkR]�ڰ��O#6P�����$A���M;�M$W:��8���̉��}���ii�5�Y�:	nfw=�,��W%:Z�e[��9󠌬�1(9��v��?N$%}{���2�KU�L'�v��X�� �AdQe2^����zt9�K=��NSVP�M�( ��2��Z���]��ʮ��gTZ:����X��K/�>��}3����y4tw��*Z�^j�r�rJ�t�R��N��N�W�eJ@wk�%P
�(������r9N��m8hXi���`��gU�A��[�TI�o�wJ��vR�X�����xz�x���r�Y�`V�l"uet�l�p��K��/���[���(Z���`n�Ά)���0�pU��Z�o�Yǧ��[��t��RX[�=���V9,�reiS�Kɔ(�*�إs�r���I6>B���g]���t�z���V=����� `N��N��;����)) ]օoTԣ�{�q���[RE����g��ד{�)fّ���`��^�Y@��_e�[��d��ߟh�j �"-��+�xĴ9�y<���Wqu=5ۊ�9YF2���إ�s��V���-b�˻gf����O�0-��H�dU��:���׋�dO5
w�+WV+'��Ǧ�a[�" !�C��^�ծ�9˾�C��#՗�ԓ�Z.�E�~���т�S�{un�b��U'7т��}�� Ĵ�6���p3kL�IR�v�Y�lVpvQ}�]1�tNc��k��}�p�2���F�+��5�eHﺸ�Q+-��3�'�wXM��թIa��31q�0���I�r�O+��ۡN�<��ޒ����&Z�aWP�~w�z����f�:�M���f�י6�˵i)�:�tF�E�q�wz]���OMW�k�7ܷ7�ZѼ�Mgc��oM;<��J�]�X�Ѻ�k��/N�m%�w�b\+ P�H��:L��s�s;��&�ww���9i=��Ն��lv�H�XwW���F��yu7�C�Y8�Ĭ^+��3yo�u�ʑ�EbyӠV�ř9r�����Ȧ"�2$�Q��%�v��tm|��>�ca�p���`
��h
s2r���UF\��� \��b|�F�ݽ@Di���*г���#��E�lG��ޮ�A�.bk��#����6&\��!Y����;{1��G���܃.o9/aɭŝ�W�4[��!�.r��7#(neaJ�$%�V71�V�5\�	V�6����|�7� ��"�g�u��kU����7D��e�mI�X�Z�b�#̻�[���!Ic=��w��4������	wd*�ap���صƮ�u
+<��x�ι��W�"u�n�"��4[��t�齍��0�����ׅ.�����xxf�e�'���6��t��E�Nc{�pk���@ͰHW�nY��
U�E�2�j5��xw\���Ɍ1��:wU��%�mۺ���8S���O�s[	�*K��L��R�ۅ��k��sd�APW�WYxv�j�KD�҅8�#��l�0��{�xc:�:����O�ֶi�ĸnt޹n�\''VjEJO�
b�š���K��=[�{1>O�H2��ZĔ��w'T'����eX�/WCH�����ؤ�3��57i
�Tcڀ�C	�H�*�ΐ�W��̑��,�jP��^e>�^x������V;ި��#]���6�8��n�4-��2�P̂p�1�}�ma�5��Pm�7�3#<#���(t�Tw�Y�yD�F�����B�\Z<����{U�9}�R�9GZ,t���C�}`��ʰ[�d�`��H^ܛȣ�`W���f����m��6���8t����%c̎��:G&*=FV8��8s��"��R%b�������4�d�U���f[��Pö�:��a�<g���s�t�s��`I[�ť�5*E��'l5�n��P�lԅ��Gc���D�>�o{�c2<ʸiY��;h-�n�޲/�֭�$w[��hȐa87u�Ї׆[�{۹B�����cs�ޭo�E1n��Tγ/��t[2�\�l�ȫs���&P.�fk�9ѹ�C-#��3y�_�&��6�m���bdc��sq�$neպ�r!%n�����cU;8�dѺu�$ѻ�I$�I$�I$�I!J9S�����Kn8�.-�eJ��| *̛�mWX̻�[�h��sn�dR5#̭�ӗy��M�Ȕ�ͨ&���'nq���'Z�c��f��w75��R�^QNaRQ�k�̒	za&I$�H��I!2N�y>Zs{��o$�k��������ɷ���P9�ǆa�P�O#)��)\�U�A��fT�X�{�.S�������Q�pL��*��w(�v�Y�K6V�Z��N�w|��os5T2�ҽ��<�}x�\3q����"z��p(зuw5wh9̮ɆP�+�9�6����`�>��8T�[���l-�D�e!GS5���17凕���m�W�q+6�P�R�Сe,��1��9�X���R]�ɖ4�m˹�u�ݼ�R�k�Ms7{�U �$���E�֚ z�GS	�( �@���G-��[]����/�IP�)X�M��nRmd�m�g��8ɧee��+����T����nzr�Y��OR�8�:jtsʆ�]ȧ��]�zY{��z�5��l�I��0ٺ�+ZG�l�A����c\�[e���]F��o�v�Ǻb[:3MLX�6.T'>]Y��<��ָ0� PU&����}b�H��wC�v974S��L��l�K&�u�eK譎�9\�Z�+#s�Z�}� t�+x��ܭs�E�M./j��][l�wb���*<
3��*SD{�Su/9^gt\��%�M�PQ����=1�`��hn���e���ܓ9J�:���]��Nĵ�7u7Pn����JŴ�����J�qT�[df��i6ml�ޣ�����ω}�����k�( s:6�C�=+s��>�;d�U^��B*0"��Hp{.�+Y���WB�95U�wj)�m�79�N0Ů���e��C��n�σ�6��Q��]%�b�t죳*Z�Ƭ<�y�E��&�L�%BY�r��)�����mK��`���{� �X�Mi�bc��hW!�֭��� ��b�U�8�2k����#�V[�x w����av&�4�Ɲ�&�\w�5!��C���������Ua�0���}B��e5���m�!��w�@��v�.wKE��g�l�����+st���M�ioT���\N�����ޛ���s,^�7}��fm��8S4Ĩ���r���{��@�䲕C�c"��&��i���ZT���`��M�;i�T�������=�:�>�9hU��m��2��wCln�G� m��b��ޡ�/��%]l��nbÒ�]	��3�ͣ�s��.i��m�R�6W�\6	�m-�ފBnp�KF�S_l��vB����̩h�����:�87�i�3�JՒܝNm_}ua�4]f(�(�����k �rq�̛V{N}c�K�p�mo
�7B�ӬB�	�Μ���ƥ46���V\v��r�r�ز���s�lk��E�'��4:�o2\���}j;��J8��tv@ٗf�@��2�Xbݶ�N6���P���faׅS�W7��Lv�˧Ovo<�;�\e2Wb�s˽n^s��OV�C��R�r	bK3U���t�t���RD^*逗�XT����D'\E�zr��KwXy�r�V*�ֻ�`��6����4Ճ��i,���/[�G�{RACf>��{��Ә�m\�d��nY�m)^�p�2�`ҪR
q�f�����
�g���
0�#zl�>P��$^�V^��"{[�y5^��Z��X�1Uw���<�EԾ�[�3���TLd��np�fP|y�h�/�ͻ�#�5Q1�w��!�+_>�VڐZ�a�Ьl�v��Pu3���q�
��1��Qʗ���U;u���׊���_qŐ3���^o9��E�aE��V��V��ە�F��׋v�!���ԍ!U����P罳�V�w�c@7�fƝ���iv��2ڲ�%�sT�(�YD�57=�6�qqC���mw�d�@�����iJ�V���b�h�ҳ�l���7o$�R�6B�����!���{���"X�(�-N���C-��Q�5'ol}xaDfm�/:�%	G���)[iI֋W�J��k]��!�����z�gd|�И�h��t�X�ц"�಻������3v3&��e�1˒>O'U�v��ⱇ��^ྌ�O>`����dln�Zݚŭ�C$��GS�]�[��ǯb<xn永}:��U�]��L�*;d�&������GyΧ���C2��8^����R��ʲ���G,\\�1� �,�O�V����ڇ�+w3�oa�@��Z��Y�/��2,5�hЫsL�%l�ō�E�xl�gu�G]*��G�x ��M�eT�DF���<�*�MY�9 ؽ�@
�ń	�h&E(�%�0�^���[�r��6b�gZ�0�݅�4��v�u�l,�Sk��F�Cp����eœ��7�(ցhw ��#��ǲJ��m���f�u��Fl�5�ntY�֥qó�?B����E���;��yXJ���h�k�L��VhNZ������]-^�4�M�r���u��'�=�2=)�m'z�]�3O�)�{��]�r[��!�Y�M+X7k]�b�i��g�0r��R�ΰ�0n�2�w�����G�e)�ʇG�~4�CFD�~QY6�4v��Ax�zv�5�jX��ݜ�\Uݬ�8�b�M	�5ZMށ����^&�,��q�� .���a�H�2��R�a����Zu�-E�D�6�O�vЖ�.���fQ�vԫ�\�ͭ)%�*��#pi�r��4J|Ow 3��us+-$O.�6��ö�B:�J�lj�T�o�Cu��K3�ѧ}̵*͡���=J�ڸ��J�r���4�s
��K�[C��+%p/Osü^l�O��X@�SN�c�͙
�v�T��:������1�ʾV*��*Jw�B覻@�X�1rػ��-�b�i���*�7Q�
�wh\OY��-��\EN �'2�v���t�6@Kuo*�T�>����Cm��Y�ځ��N���asvn�w�M;Ӑv��71�P�B��N��;I���,c+Um��.�<�Rws�֑i�����]�7�`�>��H��jn�V�&ݍ��-�yiҢV�g���&��]��2�z���X7w�f��6e� ���5^;q>��	q�;��r�wt�jt��m�ܴ֞����̕4���� ��������L����s���]��cu�G;F�W�1��3U+q8�?dU1�I��|�*N��\�6yCW֨R��f�)��n����1H�z&]��jv25}�z�լ�q9��o�J��9�z��o{�:��|��=����{J=(��R�eba;�x/nq�umv�
�}mK�j�9�wX�a�@IQ�}�b��3Q�f���VōJu��B.��RRے�͔Eܬ2Hk��0�����S�Ĭ�GI�LVLo�R8�L��<nw����*���,�3��\!:E;��[�W\�fq����'Nu�0�'����Au�,��Y�{��#b��v(�osW0��[��˨R(`����n�_N��H���
�!d�S�m��t&	�6J�O%�5Q��|k�0=�����S|3h�%fK�,��e޶���W����q���g$Y��	ѿ���i�y����ރ[XY��չ �4�h��;� ��K/8�k���fJw�v����P@�q�/s�|�w�I��3h��u���d�0�!#F�v�=��!sR�F�v���n�7Vu����������$�ǀ�|R��un�b��5kz����y�5�����2�|.D_�_=��+Q��I����97J�K�Em�D�[Q=�7�ΝJ����Pf;�҅�H�v8�:"���O3�$J�ѭ���ep�p#8�S�[�k�lna0������1=��P���5�����X�Rr��=�ś��64���Q�:F��ڿ�aWuyx��6>C�/��$���T�ay7�7oc�m��K��@T�xV�������b�iX�ӊ���9wP����N{-�h�p�kv��H�W�k	�ʅ٬�z�Mh�����U�E���o#wJ��w�Q�SN�����v),��v�4e�\�o���oQ�z�>e����e�R��J��;f�+T
�7�{Ěj��N����~�����R��u��R׼�u�m>�����)�칷���L�)l��4{�:�Ǔ@���x�P�x�T�+y�ks��a �*�ݑ�E`z�7:40�;o//kW�-�0�o��A[�Q�Vc��n��
�СS�����ѧH�c�OklV�H,h虆R�%���0���+g,�j�����%o<���o)��2q�,������8��v˶�s ]��=	u0 �z�qܛ*��&��t(�Ca��:��p;`S�Ю��d]�L���Ϋ�`;��V��W�O�L*�䓕YfmX�z[�Q��a�j16KďPWr6���,�X�q��.�:WS�6x�`�0g8�5�I��Uܻ�%�#���ќ�ʼ�:^�h���lh�f�u�G���Α��!�6�;^�2�5\���-��dXqeYxQ̔+-�!�Q50V���l��\�\���w���$�u����^�n̅�:�3dT��w^�UR�:�l�2����9�:��f+t���������8Đb�Zŝh�ڄ)Ϛ�Y�����{�L�e����hWG���`rZj���l!��1m�vb�ԭ�J���5�4�#"Y�ge'ytv�T�L_o�p�wX�d�I���Y�\��K(�h�L �m*oA{=ڃ��l�x���vQC0PA����ٚS�},bw��(�2�d��:�i�Qs�*ݼ:�0�Ij�����|S)1*C���]�gXϸF���8��i�-��ξ-�=`�7Ci���f���G��V�G�W�[yz1��sNV=�z����AO��;F3�mzR#x��	BD{��g���l�~�g*���<������&�]�l���4��.���֤�ڜ�;%sl�lZ8��R�� ��fe�j�tbm��NN��EL�Ri�17z����L��|pGs�b5>���U'�:�Â�^1�ƩM�/H��+��v(�)a���ĂW���	����l6�ٮ�$*w}�X�(�V��=mN�Վ�/�wmtEBo�#ΣA3�)�.���+Q��۴N'̀4�ܽk��4Uc��^؉¶��r�_j�(���S;v���v��kj�@ ̠vSb�ޞ:⭘�q�	l��Z�!���Ն���!m[c��p����G�{��VS2sW�sD�:Ċ��B����n�8ҘS�?OU$:�@�J�ٔ��;v�:�\GV��Ai�P��;��WfMh":��[��3�3��:���V������5���*�<$c��Yg����P㳬� �1H�0�n��u�d��o�<7V�a� 8�,ٵ*PP��*
K!P�䉨.�"wD�����u�\���'���
�6'�U��3*�m�K[\ʮY�b�5�Uv�T�h�eżpC7
����mUr�V�\�UyLW�n�b�q�mUE֕�mu�u��r�.DX�Ѵ��ek,IS�A���:�`(+�(�,�+�X��[��q1�q����Qd�6�[f�*-J�RЭ�¥@F,2���U1lXTs���V�β��<��(�9M¶�S�-�s.6�e�S)nSE���b�b�QS��k�ET��SF]���V�r������Ĭ�n[p���6���۴��fPp�J.�Y�wb�4[e)ps9��kqis����mJ�L��&ܸa�����[v���-kAL�W]ʺ�-Wu��u�j�Jb�`��^:�Y��'{x���.˷�"�z�D�1j{�W`�:̑�"��݊8/�g��>qM^}{��b�w2#��n}��;��G��gY�O���<oDf��|d'�Z�Z�_���/+��C�$���;[T>�}S��δ+�Λ-��	�F2r�S<��")��3tl���v�ሸmE���lff#���O�5�>�3e�@莻ڝ�~��œ�,j+�s�N
�J�t�l`�ƟM�\����Ko�Ș]7��5��:3U��m�7���s�ޞ�f��Yx�/���l�PQ���bo��r�1=K�#���1���M����(��v�fԏn�c0���-���[�3I��z�[�"��^Hڬ�f Nu���94��
�e�5F�l��"׫z�Kw��nf��S�7;8��73gu�F�)��y��%��~S��RO���Sp,���o���
��8�6��*�(�ßr�hFG��e��)s���[Y�RG:�E�H�q;�Ʃ�X����ӻ3/<�;;
��զ4�7^Q�'�ѼM<���T�r�C�Tr�Gs�j;�A��̓�+,��aGG�v�c� �n��pI�����zu��I*ˍ>ӳG��s��D��;���+Rky�R,�*�;vB�S�>�
�߳��>Q�$���+;���B�K-?j�S�Q��{�%��^�*�^���[����Sج�þ
os��!�������76�I�Y��3��zzN����a*w����l&׆ɽ�蹘�nf�C�s�uϺ+c4sEҵ,�s_>%V��/FU�MfJ6M&��&�˕���%�V��ՙ:��뮭H�p�
y�9�V֗8���=S����u��yf�Kٔtl��K�IV�HVTў��C�/�c����j}^��a������*���:]��EWu����X�5z�Z)�wk=*���\�#��2��Bu�	�����+O��nỨy"7U��n��=����C�{�z�9~e�mL�n�ncl^�m+�P�<�[�.�յ"=�'��ҊR��}E���G�h���'��>p�w��ӈfnN�(�X=]�Rݳ�����K�������8�%zM5�R�f��J�v}�h�\Wo{f�^k9�@�ev���Xݭ�p�2�N��{f��k)L�{y�f�D�$����)���,�$��#+�Q7�M��zz����u�Ľ���Ԡ�ߨ76��x��{~2������<�0d"�j���}���;RJ���L�l��z��ǓA��";� yaӖ�i��4݈�c$�d�;Pz��P
�W���ذ�3�
�<�R��i�r��2�����t��I*��=�V�����]y*'[^rK�����3�Ҹ��L[���ƽj�M�����.������޷O�]�s��j�齾�^��ԝ2��SD5i-�wM"1e��e����h�P�ҧ$��5�3G�to~��W��F��!r��hz�geӭxɀ�wE2ͫ�W�8Z�ݙp���3�.�v�Y�/\✔�0�/8��p���oۊ՟>iV*���g��vo%�.�Q����vj
����������X��{[ ��*��Q�4��X�X��O���a�=�>�����1�-�- �eo����h��?I��T����j= k�5��Z�c�2���e�����y��kc�c{��x�n����s�@�߭�YY�gM6ℇ_��N�r��]�|$.I?c�O�(3�:�_=��a��*Q�n_���J{]Q8;`�&\�U�6�8�#=��jK���.����Vtឝ�!>� U�X���i��� �ĚJ�@�ځ����u�t1}=�UԞ�zl�/��排�t�����rƴ:Ԣ�tvs+�͝�Ye��&�I��Ɩ�Hqh2G��G�Wﶼ(�7�M�TAC1�6sv��z̚����m�vSʍ�2EomGF���њ�Yr�lMC�X�p����!�W�|E����{k�g����3M �1�Z���0]{<���(WR��G ���'!�wl=��GodRuo5j�_�y�7���n�}o���T���kÎW�%.���T7�wԞos�Fv��S(n���cT���d�5���Fg8���+����[�����Ok��Uブ�m���u�ݍ2(����@ʮ���*�;y��*�\<��M]����Km�d�Ɩt5ݢ�hg؅���/#*%u��Z8���6V��dZ��p�1�LW�M�Wv�{��aE������X�-�9nd2T�`��Z��V�7B�]��]q7��++2��8���JK�=X�<�R���>b����Ug.�	�A�7��v��ѽp�a��s-��w��6,�Dp��t�F{e�R�UO�E�s�a����y�k4�|��/�m�y�X��#+{z���$Ȝ;}�����ltz#��ܪ��ξy�`��v��'|Z���2�AT��5�]�eE��kkc��X�S܍Nz�����;��P3j�5�)��pڞ�G/�`��[����L`Ű"�9�|��s��N����F�. �Z�t"��/��U�Ƶ�m-���ߙj�S5Wg���-��@���7HyJ�)�����;�h��6���Gl�%�궑�L�ɖ���.N���3MkVҨ��L�����#+ۂ�e��J��sU�)q���Q�Wdi�V�[�E��=���%�y���=gI=ɶ34�8��?W���]��qG�V�;�>��>���y�^l�x��Q�[je�j۩�S׷���{X��}���bql�S%:�揽�g�Y]������ ��7�����n�^N�,����tӊn��E)<^F,��>J{��Ct2[�`�	c���{3�҇GQ�4[���ǧ[N��U�YrM@��!S�V�<T>�Z
�q�~񗹝O��e��Է�ȩ9������n�i^��gfT�W�Fc�/����{�5w�7&�v���Y�Z�{�J�@7SN�(���܇ّX-�d�N�d�/P�/�]�s~�Nm�V<�n'���	�׀�{������n5ZQؓPq��T����rzkϷ^Tدj�o8�[c�+��֚�4�A���c}�}��%����B3����gg4��7��0���enj����z�Q:�Vc�>�!�!+O��!�.̴�:�y+ٓ��Q}�!e�t�V֚����--�|uN%��pW6�t���d�8�TOvU�eՕ�և��s�sA�^�!���Ozf+�ݩ0v�
�*6[�|p��L���VF��Z��H��R{-����F]��ոq�\wnQ��z����+�L8]ķ�O��� ������5!+���s��I�]v�5�ٓ���ۓ���T�w�.4y�nGl�d���w�)��]f�ڡ�ܬ��ho�EHk��:�<w~�+%����(:��^[5kq����σ(���a��Ӹs� -53��m��3����a��OH#V�\oO,�l���O��M�y�r�g7L�����^~�{�r����6�oV�GER��4��zV�a�F�j�8������Ÿ�R�{gJY����K��v��o���G
]�p�y��$%�9�]F󈺢k��V{e��=r{m���+��	�u�}uj�P�ܫY����^��EW����u_�R����9�&����e���y>�&��z��]l��D���C�d������4��mv�a�c��Z���Ծ�vV�guȫQf�U���x��\����@�4�0)yW+B�;|�]I�4�3��iH�y�1��V=�/i�ܕ(9�IntJÃ\��M��E5���W�nW�]^��u�_#��U��}i��4i��+rEλ3����8GK3OV�8m2�$���8J��k.�
`�	��3�G�%��iv�Q��,���yW��4�,�w[�M�2,��h����-��޹.��a�S�)�5|3*�Z`vb9�8ghkb���P0�a�4�+p�xi�\���z/Ir�dI���������v �ywl���(��:�̢V��`bڨ��tC��k�[W���	N�\X/MHZ{7����>�*�)j�j5�)���n��|,ʋPF�c4Ú!���H�+���o�ͤ�R]�^<�MT��]N��r��32�k�[�u�uvr�+����������^;�ѩR7Q�yj��p8���d�j\�x���
v,Ҭ�Ђ�Sm�wV�T,�t1m�ępc����B�2�	RPͫI�&�4��P�)]�Wn��4�M�rF��"R��
��N��A�T]��)�E[�i��%�U�d8e��Y�V.�qc�6�5�1�@.����]LcˁL���@2�<X��a�&�?B��YZħ ���0DEbX]B����p�!�Qs,dQP`�0�s畋s3?Mg��"��!/Z
��
X-[[��1]�����VX��@�O��9��Yhn�ˌ�u����s�Ͱ�L��͂��)sa���;Y]��.��@�H�k�5Efe���Hi�{Ki�N2��|��ұf��¶�-7m�\Ô�8HP��[����G��x�]��J��nʇ�9X�.H��,��ܐ����Q�nT)�������4//mKm��1.k�u�b�fw���Tm�Ǚ(�٩p*֙j��n\�̴��Z��mݳ\�6�DUv�nc�eSn���m����f��nf"�,bb.n�
�]5�fc[j�����:Z"��Q�U�R����T�SS2�u��M�)�FjT�cS�R�����M�DDq[6�i�]�B�s+�LfQ�UUEUw0�b��
��T2�]�ݦA2�J�b�Z�뉫j#^p����FZW"��W[PmGw�5VԻ�\�d��,�2�+��1�n��e5�Y�Sv����es*d��V�ܵ7s�3rf������؉m��ppG�v�S:~��s�˞�39�Œ#}5=���cךu�!�L�[]ƹS�rsT���ۆ���!+����l�dv80#��#���-]˓��Vq'ή��u�I�\��OE!֠������Q��u0g��M��C��4����}���ʺV*�����q�~��ǟ�����||)2��n�ow��݇7|-L���c̯���MbX�Vsy������O���D�����;�m://�P��z��cɿW�
�.�	�{��v�$��Y�,9m�ĽX�
2lބv���5�zu�M�~�=\ؼ��OD�d�$2����-ux��Wp�[�s^��%�ٰ�b���\%dv��}{22rܸ���~O<�^ѓ�!��f�N�v3�"��%S������9=;��Ӝ���M���en���S��j�[Q�E�`��}q����e�tS��*�V`��L�Qts���띓p޵~G��w^y;�l_r��;ñ���lgf8�g(���z��TJ���N�ULP	b|枞�6��f=\V5���`u�,fS�o�Vd����8�[��{��j����Ǖݧ;�diqz��+b7&x�7�> �ٶ��u{�\M'�rlG-�}eeZ�L��-�A]�/W��<-kY�w���G�:�u����h�'�Ӿ�Շ�py�֪{�Z��\'��?y�bf��]��v@�)N`nY�P�ws/��|K�@ik�*�B+�	y�{種����+0�ؚ�>����v3���̳��"%,Ps�ru��${y/�*ӺۺϤ��C�s[ݑZ;7��i�.6]>֖X�`��V�DZ�'��Y2ZU�Ih��4^��i�4�Jg�I�٣���:�s�޻@�+yNg͜�;��&vn)���=�7
:B.9���£���*1S\�t���C�tH�=��s[��<̼��+넥T)j,��{U+6���2�]{rt՟ o3^���e��=���5���k�pVc�g*QǞ(�ɕ:_�;e?.�װ˲xM�]]f�a[;Ͻ�s��s�Lx�@�����R��s��'���]6�����^GY)�`s}��U(��ݖ��]��B�#8�y���z�o~�����/�%|�P,�c3.Z7�4�_A|��"���p���v�q�⓴�%�2'��b��8�4)�*�e��e�}�E���U��lnj�C��,S��A�G��O;���������I��'N��ORk��!��t�����t���O��z����'�p>������{�w�߳��}�_�vȤ���;@��!L�!����:�'l���y?2N��t���C�=�t��>Bx�و��#z��=y�4�/�S���{ގ���9l�[$�&��z��vO�}R|���g��x���u���u}�Ͼϻ�z3z�ߕ�s�N q���'�>�r���	��2tɹI�'hys��?P�t�zÝY��L?'��'�;�ξ��`q���ԟ2e x�=�2Oi������́�J�ɻ@;I�P�2�ϐ�U:����B�q��S�D�@�D}�>�z!L��&KO���	�"�̇�����z�3�2,5;a=�l�2w�Ч��k��|q|�ӏz>����ǣ��ĆRE'��O����~I
��'��G��O�O�'�N�����>�X�{�\�7����6b��Gޱ��@ɽ���3P�����=w�H���������!�!�'�u�L�#���ؖ*c����BCʫ����EM�5��@"�yǱ�����t���o�#��<�:�pY��H2�1st�d
�����4uiy}�鋥��e�8�����ۑ�|�sO��>9���!>z2�t��@��~Bv²2t}��O�I�x²J�z��&��GFy���μ������O��>B�NЕ��~�t��'-	�2ot=d�Ho��~`z�ΨO
a���O̾�����������_��@���2}N�2~a�'&��NІNX$=Cr�qd��I:�GL{�c�b"1����7�δ����0��~P��|3�ԓ�7���>d7���3���t�;��q!��t���3�<cDt��ُj�����oܹ��=�q"�ԓ�'i��C����:~H>����!����~a���+G�Ǡ�z:}'�>��d6�~�Vgr���`}�w��$��O��Rk�>a|���O�:g��T1�LB�C��DG�4*�e���KWܿ�:gI<`q��P�3s$��_l��~��S�Hz�����!�����x�z��yϳ>�T������w��:C��Hg�x��жI"�������A�I��'��d�����5���R��q߳���~�������!����z� �]��$��OP�����E ��ז����8��p�'�q��3�������3�>�������>���Cԇ�6�c�~d?2z��Hgv�q��8��䷄1��T�sT칞9�y��3�L���0�z�]�ŖR&�^���)J�$a>����-�P�+Q:Z�l�){W��Ƽh8�Ҵ�}�+�ޮ�[][8���O�,`sѸ�.R�"e�5tS�o�ԓ�=d5�0/(�������$�z�����@��d�0��=d�$X���:�p����}�=w���~믤�����?2��2NNP��{~d�!Y�a���4��z���C�Pܳݡ�aw��zo�����y��^_v��=���f@񓴛2�x�f�Bz�uՓ�C�$+����<�	��blO�B�A@��Cy����w��5���a�	��"��E��5�d������X|����%`{�)?'L�����{�z���~~�C��z����'����!���!?%a1���@�7��	�%@9�MI�޹����=�z��?B'��bIP�;���C�O�1=C�`z��~BT��:gl'- �&Vz�8�2�����p��ǭq��mɽ�{pi䩹�s�A�{��yϢ!	����<�@���q����`z��>���S�%``y`v��ʄ�d��y�w�ܐ���^�|�i�'l<H)�P����<a8�O�x���'=�$>C������<�9������9��y���|�ä�L�d��v�;Iϩ!��2,�����3����2{C�䁿S��O|�K�9����_��N����ߣ�sE�^��iՁ�"��'�NwOXC7ܑd��2O�<`t�~a��>d;`z�}��sQ]��|��bf��GFP��$�ۂjm*�(0�Aaξ�Y���˩�G�]�t��ۮr����E�6��;��ʮG��Y�6�K�b�<k�<�W\�[�.8��e�t�{�y��� x�>�!�$�8���=I�i+	���$�|�wh~������x���������4ޮo�B3��?!?$ߨO������:?RB���hE���$��;@�'�IJ����{��=SU�ӓq9W�}�8�1f���!�~N��������0�!��@�>9C�I�4>��!�X�3�L�GLD9�7����%���s荬��z@>>I�:��I�|����̇�d+!~�=C�M����8��,&u�?�s�y����~��<d�'�PXjl��'�wd���;�gl�����I�t1�9�����r�z#�ѿR��r��O��DB��֫�M����&��l�s���zI=CyI?0<2NЩ�d��X~@�����>>���u����}��
Ȯѐ��3)�!�����	���;I^�6m$�%foXćL���,>Bg�� )|κ��s�}�޿���v�l>H>�2,3�C�Pܧ�'���Rc�Iհ:I�&��x�+6}d�?S�>d=a�y�>�ڝgׯs�:��y���>9�T�3Rv�P�������Ot~��5�z�~d�}�d�	�8e	�q&�� ������u����}�|CN�P��$��ߔ!�<d�~������k��X'�3����EG΢f#'�1�c�C����]�_S ����F��n��=h��bP�\�W+T��2��4>�Z�>��<�h����BS���+w^�3�[>式/A\�-����X�A�ܔ���l2�Z#8C
B��ҷ�q�/b��=`i��q����k ��z�a�;`x���:��?!�������7��g�w￹��HJ����H�a�:��@�́�I�����	�"�݄�SN�v�t��?$��!��O9�����ל�<��]|�N�k&�M~?S�!����Y�(2gt�����O)�0�
�(B�^2�kZ�Xi�����f�!Bg�3!r�+´�KLd�Y��$5!���ԓm!�O̞'�C������Y<d������{߽�������}�	���i���@�>I�;d?=�P���I�~�rHg�Ha`K��j�\ mz�<'���<�U�k�L���{����'Y!�>�Ӧv��'<����a;a�ĝ����Ɉ��S��xk�9��F�_r6����$���	�I�=d�&�0<�z��t����8ϒ������� T�B��ݝ/�)C`g#�ܲ���Dv���2)0����ϳ���>�����g.wS_�׮���p$�&��]��ۣ<�7�Z�b]���o997�oT.�j�5��n���5�S�^�Q��S�7��wў�j��<3#�"����l�v�W!Gp�T�3���W)_�=7�2��-{|f�ܮ�����l���QT'��2s!γ$QI��I���O?�ǯ֝��ҋ�{�s�d���{|�&�����W��M�u������5y;��UiWS<K�1p�<!-r����M�X�8�X#NU�WR]A���kιSQ�vm\�=��;Z$����������&]:��Q�z�ZĹ)���j^մr�g\�v��C�S^�͠f��_:���]zϤ[�q�ދ�x�'xqr����7��gzڭ�J�ڑ}�پOR�gN�:������[q�g��>��r���-=���y{gW����ap��Y�x:��$��]���6!z	iW�e���搠@[W�d��X����}�9;]�3��Ƽ[�Y�5�+)�fWV_3���b�7�n��)������s���"��x�ʁ�0�>�
Ӌ�7mk8Ȣ޾V%'��uJ��;�oem��wTwR}�����~�}�uC��&���Rj���ߜ�R�,�/%�5O?f~��������Mt=�yV�n1V5��kyK	�E����P;�i�P�'4�H�q� �6����A{���Z��T�N������\��{��y��gj)�%��WW����)���(q\�5S�Y���;��h��T�c�~��iQ�)J{���6�)cvy���ˊ��&q��"a�.y�9�S2_��7�����V��gAu�h^���ش��̛M25���ɷϬ�Yպ-[�|oc�r�β4e�4�w@Y���R��NVFۚ>��W\a1�Fi�i�ҕE�[�mf]t\���}7�ݼ�˱��ɇw �>�jᴤ���ʺ�u�3��i�&;��7jqI;���*�d���S��˝���5l̺эW�Ge�o���O1�5�\�.b�y�trb�(&�9$��3�zD5f�����Ej�Ce%B;��[pt�x̼���5M�"v�Ȅ�ұ۶MfpĨ�ŝ��{��7�d�O,�ٙ���V��Futm��R��=p�I �"���~�o*[��u�S���qp!���a/�M}`��vU�Q�4:�$���j�ɼ��7:K����[���f�����ViX_��o>�YZ�f�6��`���\ԴfX��P�5�c`���\�
����9�t7e���&�՝q愴�}@�2���?t�M��J��)b����diw�e��O�F�=����~�І�u�d1^;fbw&1�\�c+�k)0�b�8�`�����2ŕWn�RS�Xl�#����b��ݪ�7��9��t+Yx�;+#����>ȰU�V��Q9��NR���yt�ha� $!It��`�9%��n�bXʅI15�+�SىǆVTP2�T@ �XpfR9(�ؖ���7��;��˒�f
$I3��`�-řh`�����Uv�<	�@�Be)O��^r	R~�ONSF�X�T�M���ݖ��J�"�5j�:�A@���4��e��F���k�!:	�buB���z�J ֩�J�:�[q���;mԊ�Bɩ�9(��JV�%��UԨ��ukM�2���]:6�i�ݔm�~2� �ΐ�:ڎ���)iv7���!Y�)J�c&ʇS�X�4�$\�Y��7.;+�@Dۅ_[�v{����������;J����}w%����k����v�#�Qo��m�����`��TL�J�a��,�\�kG-PW(]�������p�QE�۹r�ڙ�0�nQUƪ.5EUe.;��Fڙ�`��h�8��"5�T�U�ib���DDA��5��h�ʹY��%˘YU�¨�R�G�TR�PU1ԥ��F�k�R��R����q2a����D�娪�V��̬Rڪ�J��!mĹx��*�h�l�PQDQkQT�������m�����QF�������iC,�(��j�Yk+ˉ�ƮZ�������˿�.z����W*$�e�1I�:�r�k��j]�VѤ.�Fj���R��=�Du.8�y_�Ǯ;1�=�q���~u����>����pTX�y��7��w�`�.�U�
�f��k��U�}�||sLQi�,� ß[tz������h�'<�����u�(��ݒ�g����hͻ�˔�9�S"8�Rg�9�Z�5~�<�[\�bз0�l)�n���-�R��3L*�S�����%-��}�$�[��h�O��YVh[�׺=�ҋ+V�ݍ�,3������Q�_<+�eT8��79P����q҂�s�BM�Q�yZ�QO�;�������d�}�F��`Բ���w�5��ju#ws�.ʸw�t'�u��|XYD�Z.E��W�X�y���(��z���=�5})�*���)X�WÖ��P���4�T̓lt�ؒ����oG@�-D���=��Q:�3�f�k$鋆.\��z�p�]�p�O-���#2�M ;�mYi�[�.J�ʘ���:�����JX��QG��1���u�����&�:��s^Ԥ&�5�%	�����I°�p3r��=�f�ޭs��C:�������qjF�+8���]��n�(6�³��4��}k+M�Goy({f%��W����;�ߣ�����̵GbB�w��7�2f��Z�X�q�o��X���k�v�41ss�;�i����2�3���|�{ͅ�wl��ro]��N��&��2�u�Rf;4���\t�>$�v\c��`e�,��t&�ٜ��Xi�nR5ffw^Yȥ�T�2����o*�I=#�s�/�z=�Ab{���~xtT��Ι�ך�v��fW�e<�lf�}ۛ���g�eA�q{(�:�9�u����9�[&"R��y��n��& Tbz*�iJp�i\��W��E�ge�mCow[R�9��-c�n���}/ZA8��+�Ӎ{�׳������Fgr{�EwO
{�L����kC)��Gy,� t WB��}.�3��ꀗ�����we�;ۈdy7'[���{itU��:Y��G��)�S��S�:�v����0��x�9�~�]:�Qǰt�.^�g�m�fg��k��r}y�_���L�P-�_����Т1��~���.T8��y�z.�|��iV9��	��V �W����Ɉ9z_k3���"z���i-�$q9�꯾���o�fc�4�v�5�����zH��W�������v����.��b#O��3�e��P�uu�7z�(����m����UӁ^V���+_:��.�ʋb�e[z�\=]ˬ��M��,Lw"�k6˳�
�k�c�rw'<�����n��g�����s,4b����S*%��3�rn��O���7l��#Yz�rk�OϓU��Rsk3"���缴�k�����z<�ܩTl.k��w���#:�:�٨����w]h��d:������oïs͏k���ɞ��R��.��iWs��IΘ�kV�ǯ�]!����D���XL��e;�)�.f�K��;���&�ִ��E=���Y�F7���Vh��ұ}k�f���G�!�|�"k�U�^l윊R(�����Ta���ʠp�����sy7oN��5cd=TՑ�d✡o*ή�0\c�ty�Jb����K�y�=���.LD�O�^^��D��sx�x%!��l��򤮪G�F��P���*�Z�oW*J��l�=����n�w�������_`��i=q�>�k���=Y�m�>Yr�x� �*"ң�,���U�c�gr��V�Ԝ:{f����E8�y(��Xٱ�����(��|}��sr�`L��uu|�X>����-���f�xNC��x�nӝU).i۵p	X2�,g5���J����Cܵw�;�',$�m_ #�X�wiEVk���]�\��fhjm̵u���|�	θ�I��r�����{�㺛�~v�Qg�j*�bn���va�كA��|���YD�Z�@ң4��}�<�{=��b4��Q@� ��n_��Ĳ�rE�f�c��s�y�>[FXh,����l����-�bS'R�K\��gq�g_��7t�+#M��w��gYO����n���H��*���9A�^U�h6��i��ך][������lwM>G�tb��c�Օ��.�j�S��[�Ey.Q���Q���ԯ,��z��;�]*Z=�'{��!�8N���l�׌���������Yѡ�w�u��;��K����&���2Mj,̍t�y��z]��Z��9{z��,uP��f�U>���=�2m�Z�ըu:(�2NY٫c�VN/i	��FI������%�{�׵v9��;�O��9�A���J(Mn����%�pۏ[���G��T{�)D���n��%��,�~���[��/YJ9���U��K�S&�w�Xh�s[:��aOL�\MTsA�w�ܤ��Y}g��3�"�>=�Q�sM�Ζѻ�ӽ&��݃���mP>1�b���&	Ƌ\�Ò����(F��J���i�h������.�>�8�"#�rw.ѝ�`v�5�	���׭�s\����=.mQ�&Ӻ��ӈ+�O��E{Ӟ"���O_��*oS�^o>��@�wag��3��Y�����>�NS�6�mS{g)9u�ݞ�������3-h�XS�q��s8l�L�v\B~+arv���3��e@vܭ��|�oQx�hgZ��-�re�s2R�B�c{i��JV�Kk�������o%�����++[v!b�nW�9�(&��G�J����*��^{�h.���iebqq]���2;a�OD��j����J�|����ޏ��)�f��헽��ċ+�35�s�I�/�{��86�	�7�Zi�z4vh�IyN謑g��g�5ë׍�.;�,΍Em��F�{����D�+[ۉ�D�s)���/m�>��Ш�o���	�؟�򖄗&�5sRq�WF[E�/"9Z�����)ĝ��B���,������^�|؞��|��4�KMqy]��ڕ�;�Ȟԥْ�9���i���Un�K9�	�Ʋ�	gGSB��PB'hA�)9�>h���o�E�+�[�$P�R侏Dz=�)������]�*�h-����_9�ǎĮ[��l��]�y���^����/pѐw��'~Y-MGݝ{���m6�R�8LXA+�e*�3N)e����
[3=r�7ePΆ{-'BT�;!�ѳ�JE����P#���7.��Mga�=��R⣺w�ӑ[��l�cʚ��N�8��{��tG)�RU�SFn-�v��oUOfN�)
1�_X�3V{�r�~�~��u&R���CwGs[��Δ��[;��3E'@�d��p��4Qꞿ"����͞��nyt2z�H$m��X���w�$2V�g}$���%��
 ��n��u+�kzOq9U�1�F��f�����Km2\�yŌ�Yl�V4�9Xm�ء�����U}UP�m��f��ݑ%� 86G]U��SY�s�q��zq�~��)����m*ʳ�Uǘ=)��&ʞ���{�c�?DP��m2�ov\\��gs[����^qn�zqwZ�����0_��񯫎N1�}q��^�+z5^��l:Ʒ����ޫ_i)�S��n�b:F.��FԔ�f�Id���
ۓ�UR������5KeҾ؇)���,l�,�U�i�����>�{"��M<\��2�du���t��ڵ�o9w)���7��Ն�5�(*�`gI5��f�f3wm�:�dZ4�u�7 ��:���4���lm�V3	Zy���M4H�.&CʘN���t8Zd��J��eX;�J����y���b��6�ˈ����W8��Wxݸ�P�Z]���l��Մj�NĜ84�G�Ge�KX�֦��Ɲ�����Z�*Y�K�V-A|úd�]����̼q /r�d�dR�Z�c9\�v�
{�J+�=�Q�2%���W�mr"F-N��f���u0N�g�Յih��oSx��¢x4���a�+�B�F�E�f�}]7�q�%Q㬸���]�ن���n�M��Qdo�6��1�!8%�Q.5�:=�ʺڵ�#��r���	٬�]�m�y�X�.���(dP_^L6�)�R��Q!_i$��.ݵDa&,4��MrG�	A�]�v����=@r}f{���\��h�����m][T�#�K�YH^���ǅ�iHfA��{����q<�P�l�R���/�X�����Z��
>t"���{������b����ۼ�n��ﺃvϰ�2��i��D��/C3�B�0\Na�Lxs/�x^VHݗw�N]���B���t���I�����@z~�C��a$��0
�ux>�l����k6/��ɉ;���:��)U�vp�I,6F*Y�a��:i;Q:͕�����YMx(j��L�jIQ<;V%`���h�FFo.��HrWN]�+e ����50�g�QCd�ZQ�JZ��h��pM�N�So�6%�t��;˰�m��pX�0NӖ�,�i��~�g5=Je�aJV(�vx<t�U�a�O`l��4��Lg&t&-ޔ�������s��Ms��,�G�'���4�r�ya	c&er;��T�X�6WMO&[�c�$�ȀY�ɭ����"HVL���"R䮘�]o�}W�b5�-T�EUィ�XVTm�1�cmDYiEV�UJ��u��S-�EqR���,MLUqQ�jV�UUj�f,V+[s1�Z[UFV��8��U`�[R���QFe8��R�+Z�U^e�V�lT�\\�Q�nf6¦e�m[Z�S\�j���ZUm��+�Ʋ�7n�lk-jj\�̦+YFҬ�kPZkm��s&%�%-+�&DLiS-��[b��bZCr��\S
6��
SS҅E��I���`e�ɃR�(Q��D �� ( j��?=��3Ln{��eq�Z�3
x1K�œT�ϡh�ӛWm�
��#.I꯾���#F?x��� ���l;��tOt��G�U8"����(�n2G�kw�U@��(R����]#w-�.��oc5�9]����w�4Ou[<T�-�J�a�|���`��訿��J�17=l�3M[v�Y���:��̮�5Yi+�3�{���_�"�u�9�.'U�l��Q���f�=z�Z�Ou�WZ�o˖Tgnc�u��vz�S�9���5�ض	�qb[w#gb�e�&�ӡu�d���'��gH�{�W �/'	E/M
OW��*5][VVQY��0���JV��eJ��JW�ξ�����^�Ӿz"��]�@�ś�_SQ�z�ϔD�%�-Ǫ�6�3�_a���f=ot�b3��C�P�黋$�R���kOj<�Ij�-�WD�$���p��)����WBF&�1��UUU�fx^����=c�sq��z�sm}:���4����͆0�=��G��tY�k8�&��co-�9pK����Z���Q%�Q��-���M8�]y¢�Vӛ.�]\x�&��e�,��~������F�@�G�T`t+���V�8bn-o"�Z�
!��t�V;i5qaUhx�� 8^S��$��+�+�*Q^W�/5���A�-�x�t�p��wn%���zq�=�_R�S}�cgW<�;z�ī�.v�n�(�IҘ6�����Q�������cՇ�x�;�*'�C֮@��WCͣ�Q���)"�<9t�1���.@2��}@�{u�{9���eca�y����|�.JRgoo%��#��t�����1��h$���}�)i�wy
ߟm�K>~�{=Is�������i�z
!��;�q���*�n3�I�t����H䱛��9�����Չ�U��
��V��J���;�0�mf�C�q�+S��PwW�Kl+���+z�zNs���}W�k',��N���3�U!0t�UʺfQ�޽�u�������9WC��cDi�JrD�u�S�v�{�z��=��X���(�O����1�yn��wN֮�>+^����[�*/R�����t�[��\"�
��~6
J����^N��X��ihc�)UC�/�2�a�xT��t��0�2��]��Y껩n�V:���p
�3�݈M�q�??�Uhݧ�P���YC~�J5��Ra�xN-�P>Wԕi�ص��9'������@�%;0\��Lw�����J�wL��[9����NM����:fR�x�q�ĵ._��DG��q���5��'��\1� m����pߎұĠ����x��w��oi_�v���ۨf|Պ^礱\�]GB�D{۝Sd���i��P?�T�֍��p�c��jt�����۝�TW�v/�%�ɾϳqh�D|��TF
z�P�0	V�0�z����ŋ\�o����(9���\/�P�q��N� �Z�y�=�2����p����r��g�p��᩵�D��z�ϲ�U�!	^���z���f���s�f�}P�t�ߺ�9���9�P�x�bo�m���˨��\�+�=����T[K��53�ɞz<7��9-6<qh�	�H�r�}>(S�8�\5'EHZ�fX�VQ� Ʋ�fgfD>^�W<��'F�Pd?
�k���yj�"H�	�eZ8��=����&ӧYP3"��S�`��C�^ռp����N,���b���LF+En�EѼw�TW�S;7MLq{kVr��{����x��n�d��ُ�+������6%Ҝ���M�CBC|j��X�ksp��1U���<�)Q1�a��ђ?����	����[&M��>�O*��i>�þGF�������,&#VO�w����<�d�޶�{�n��h	~U�g��x\8j�����k3Vg[C�b�>̼��X^��ᩭp� u�
�i�q��&�x>hR�cݻ��rB���+�h�ǆV�����S�r��Q,8��%�2�|����^r����x�"?o@���.��zr���q�R��2�u�~U��D�{�����,>,)�F�!�fo��=W�]o��-=����ÃI�]j�
������޶�@�|��{p�qі���A�Fa�sdT��˫��.�P�`�yoQcm^��^V�7�P����FpPŒ�Y���t��.J R�i�/��j��֊����=�@<̚�};r��h��]��:XT�4��+��bm0s'^�QeHN#��M��t�5��Қ�cr~��着��8Ү�3��G�:\NX���=^=�=���yT�q�c�lE{�ۆ��_mfz��{�>ϝ�s��xTt
�0Q�>��:�t���#��+=��@x2D��;N�z�93
T�4���)q�'\O<>>63M���q�(�@�>�����l)�R�}	J�:��48Gk��
҅���-/MXє ����[)c̩��)�/S��0��Y��7Ѭ���ᣙ�H��q��zx짜���-y�V�z��Zo�8X�PA�T���)`)OE���vB��~K��8pU�A� ��`���[;1�,�������Xt��0�^�4�hk�MX�Ǉ(��H�p��[�o�I�k9[1�&%��5P�	���rZ\j٭ų��7E[�QɌYҥ���g6�E�.�T��Z��t�P�����]r�ӹ6�zO\]^�H��=K��J�UU_US���{f�^$�@~Wf�#�/����լK�A]��]J��0�=�n���|�̱j�p��3��G���pX��P0��g�9��{-W���Uʟ1Y�q��p�Q�������E�ogx/�pb��&�s�i͜��瑭Gæش!��k3��t�����\ܺr�N1��5V:��-}���k���LS��w��iG��2$��ʒ����&&����h�Z^�&sl��w�������z+���k�LR��PUlEQ�Z@�^����~�b�n��,;�Y�]x�gx�7^U�Z0J<��s1Wy6K^���ۜ;�7خ_$�]2*] 3z����ƪ91GH����76e���Ţ�c3�8��O9p�eyW����M�;}�Xh�=<Bb�L�����Ji��]�j� z1B3r�k�	����u[[�dT��3���r�� e�{��'XO���NZ�v� �Nܟ�����f��<�:��.��v"��P��X�h����h��2��n[��n+�w���)�|+MiU�u�4�#
ӂ�P�<,xW�n ʷo��j䔈.$9ɵԤJ���QOj^� 8���x�|)CZ3�'	�B�s}�p�
�]�^��B��݈M�hl�h�<��y��V��ٷ9"w}���Pphp�\�����lu��=����ɱJ��o��܉�c��g���\�]K�6�|�o���A�S���z��\��f=���������B�rň38�1~HsV���r�ｐ����/�ʓK^��X4�Z(�7{z,\�=���������G"��h�O�
uW��Ϝ�����߷��!���yX���C�Pd�X��A�P�eg/��7ak6צ��$�ԭ�����^�yK��}-��<�s�t��s�\;p�j�. rt�#jp��S�ׂ�r�vۈ�I��4\���O�}����L�Ln]hgR�Y]*i:sӚ9uC~;=B5'j��F�)���C��rP�p`�YJ��v(4k�^���/�����:7�r��c�A�F���[������_�Agu�љN����%n�NEۼ�N�v�Ƙ��6fQ�����}��sKE���e�ĺ�^^ɾ�؈�CF
��U&r�*��d��].���e��7 �~�W_^���]�ǫHV���U��X!�,t�2��0�TV��nW9q>< �c�уGH�֒<>��Ia3�B�̥eowjd� ��]7���:���P��8�9���MEu)]��YY�3V&��»�k��N*�|6��`0�1SM?jat�f�;Ҳ{}�a��<<r�I�<)x��P�`�P�P�u���Ճ3$����S$��n�r#0\���#+r�dz2�OjPUԂ��S�g����^_`�^�ۄ�u���+�:{Sp��(��pS8�5�e�}��Z�:�*W&֮ē��z#�i��nd���o�R��x��T�-x�ƛK���I��h�v)N_CN�Z�M�N?7��U��F���M7�`����X
}���n�f�B�թ�u�E��PS�Ju�7��f�� �g*����u�i�A��f��1|4\e}���5���k�K�PW;�WBK��VX�Z
۔�h�mQ���W�����"Ws���#w3�]k`�vf�����ӄl������Y������F{{}�E�?M=��� l0�c˖��b�,�S�Z����oo�箶ջd���ي �͌ё�Q<)�.�+N^�V���	v�qЇ�&5�Ύ�
j�A۫�*G�'.3��~8j_��]]Xzb>?^��C_�hZ@?U/n{}��h9p�j��+�n�\����	��7`w��ic��,o�o�*�/%��H��S|ؗ�գضf���5a���C"5���J ���-	gqV�SDp��uX��R�V2�(v��Q��>��;&X��w�Q3����a�O+)�V+���P6U����0;J���܌=7�� ْ��͔
#�{��X=�G �ZK�E�ň��-�7a�fEm�&�)��e*�,M��H��]:�3�dV��`G�n��ZRb�_\�Y��BU��J�9�BɃ���3'#v�f�H홌v��/�Oz�M�{bGk2;/�5-z�Ri;�QL����ٝ+9�<F�Su)]8���V_5��v��{��j�D�{%����	e+�j��
9�T�3*`�����Y!��P9��MD�T"�J���k�7�~c��ת�)�P^�xrE{�qJ�k������Li��|��h��$]�kmt�˧xk��V*{P�-�$�\J4�108�/M$��!�.��ct��̩EM�p<�ܷ�,*���n�Y�z�,���{ݥ;�(!j6�ܩ�n�r�U�)�齡r�Hc�J�r�]���euph�c��Z�]���4-�q픢���D�FBr�) ���	�5�3�%��b�ۡ%��,��V�M�����b�3[<�fj,�I��{7�Y7�I�����NZjc&��wJ�YK�-\�1sa����I��*�m��(ƘѯeZ�]yd\�ަ$78=�.���K�h�[���Ù��dGn�:�v�Prϲ��:�j�T�����v��s�
������:yٷQv*��,��WLA�q���5�*:7U��b����p�V>�pd�Em̮Ρ�u��j�9�űj�x�t������}'05۠qp2�J�&d�B�����)��;��/3������f	+�6N���Z��ūJ�-�-���dU���S�k��Q�%,FҒ�(������QJZ#30�0JZ-Dv���h�Um�V,���Lh�QNd�ں㕋J�ڋKE+T[X���˘��q1�&�J��ז�̩�m�5E�V�cmm1�KK)Km��dĥ����e")�Ķ�Wq�VGrd�M,���Kc˃�"(�ZZ���j����\�ԭ��s-����J!mq���6�;�A\�+cl�娉Z����E]����2�1��Q+Tm���.RW���j`�Xb��绋Y�ȍԞtز��PW=�o��*�Q�r�]�̼쵅ㄷ'������0��
�4o����7�E �F@j86�� UU'$��cxq�z�����lx�T^X���5!��+�U��^����0��7��y�N���/7O����KF�Qv�Z5��������S�q�^d<;��FЕ�[��^χ �T'%��Rf�/�
�7�q������޺����� m�� �����:Z�������l+���
�ZX*㢽��7��ظA��Ik/eڜ��P����{U.�����U�k����T�����q|z�V*w���ŭFޑ	���,X��Ga��*&�*�q�#�ѽ��3b��\�s���:b�(�tJEk��jm{nl��3�X��k���q���3�P�Wu��t(��/�[���|��߯�Dr��w�w,�B�40�Y0H���>��Ρ5��Պ���PB NnU�=�Eً��]����-�� e[�p5�>O{J���"�oވ���T�ph�z������#�>Z8m�,p���3U@�}�W�z�4v7+yԀ��ؿNY�S6�T�嵳v����ׂ��%���W7SK>v{���Cm�F�y�J��"�-[٢�L��w�5�ՠ:�p|���σ��#p�]i�|� Gg.u���=y��(GXeT:�I��NL�/�+1`�8�{gY��S�~ם�K���A�9�WJn �]X��_^ɏ���B���/
��6/ ��GE�v������C�Ty�,ڭ�e�`Ӌ"Y�KR�Qr�M�`GK��VQ�<tTԴ ��j����߮]�4tHq�O�֫�Ȕ�K�E!2#�)�&zq�5*/2Ҟ�^<穑f�S����&0V����Q�-&�pz|��	0��u8��l�oNe9ŕ;1fD��L�k�[ǧ|%�� �,�+d�$+�s�J���/0�����撈���㵚�L��c�rX"e+�W5Ir�ԗ�z"=WX�$��\��,�4����j���ܣ�kZv�_��Xғ�j��WW����)�����4�zυe��2�����3;��S���:D90����N\>��RhT�La�j`�;#\�/Suy2�]�s��T����}��٬<�p}��O
�~Z%�Q㉬�&&:�[�),þ�6�9�P�'�ڷ��e�5����Y��=-�~���"��uY:]ok�֧��uj��q.��e�X�^�&|��-���ok��{�ςߎ;�2�̥��(�B�5ī��6^
��<j�n  #��4���Ȯ�F��ɾAC�����V:Q���
zi�Yy�Ʉ�t��;N\��pݩ5Th�Ә��Ý5�]r�Qu
�e�Ό����aѺG��F��W&p�o�L�yq�^^�F7�]K�T�ט9�^&�᠜�����^NE���{w�!�kS�g8�
.�I}��$�s�`�ޝ`���J��%��W����ܫ��o-{��� �z�E�V�\�:��4j������7O`�V����d*VE�:Ў��l�1�%��L�u
s�9��*m���j2���i�LV
�	�FS���:� {�����87�f����3c�&����F��*p�§���p��f�)E�[Hů1r��{N&)�&UzzS��^/	H��i2�`���Lɼe�M̛�ma��o6������u��ȩ��q`f�b�o�j9�//p��mx?���Ly�-o()�]:���u�F�7�*�OSBM��g´z�4�uX���c=�ø��\�V����w�n�;�ǳ����|�8.��+��j��OV�ce�T)��݈�|��)�oe9���e�
�
���b�DӬ��s���T�G!��D\�Ap�E�P^�"��
iY7���n67
:m�T��\���^����V���.n\��12:c�vr�)ŝ��$�9�8���}�W���^��6�8�H&?U1Lz`݀����U��9��ׯ���Ŵ�}�]�9����~���`�BP�n��Y{��<��2]�)�j�:c�I�.rU��K�ۮ��1BݫykG��'���#n�J�Κ>��._,���%�6}�R��5臈81�l���������2�@��ε��pP�^! �V�ڌ��/����C��&
�_��E��	:P:x{��iV�s|^�����U���2�7O����豋�k��6QAy+��oc^��p�/ؼ9�u
���^�����|�S5�GV�}��a
�t.ep��������P���Ǣ���G��N������+2.d�a����� F��{'�@Ы��o���M��=�xи���	��qɽu1��R�j��j���	��4�(Jй ��F"7�\6��X�:q��|����&B��]Ct�R;����6&j ��a�����8�'�ꪪ�c�L����9���7GE:��ڨ��E��QT�zK���|���bic��敆,X��Ga���P��^�s�D)foF�},bQ(�e*dFgQYQHS
��� ��`�U{G@����ˮw��Nv���S3�Q�Z�}S;;G�\��x޷V�q7-�u�G��:ポ�k�i��=/Yw�.I/BUb�m7�A/�z�������G^U�h�2wY��=��z���}seݛ���5��-�ЯԺ](k����Ho3�>�^T�[�@�}&%��h������WWX�˧��Ȉ����i����hL߱WNW?p/��vi#,������/���L?��\5����j�k#
ӂ�ypp�<:�zb񫸘C=�x��#Aw��K��uu:ת]��74R����W�]eN���$�sm��P���#ƌ̝�y2�f��� �Vr&��:H�s��W��{;چ3���?(xx��<8/�˃�xs^N�a�])-:�5�H����7kX���X�}�BQ��:�:��@`�>9M�͗|�
��\ؼF�XR/kʝ9�<�P�Y�X8>G��Gm���|��=;ow�IHx�+Jb��IR�ԫ�X*��8��b��O\�wp���h�${ƥ�JJ��,J�U��j�K���޲'\��o�����N%�K.����&������P�e��7[��nF�j�w�t)�i���.pR��Ή;����V���e罾��W���[a_�L7F��Lw��Zs)���,л�ukԕ�R�̾�%z����U�Z����J�9Rp>����K�����=����=hOԩP��0h��Ѣyo'�{�yÒ�^򚡣$����N�pZ��&q����ۍ�7KfJG'p�[��R2�X��/M_��Y��ط�>aV�	}����_he��W�^ܩvuZ1P4b��1��꯾���'��Q#�,������[����k&S�o�磝v����R�ӃN�7�eSy׼�:�p ����9�f����q�Z*���8���h�N.�1�E\�J� )}y�Ʉ�n�����Zq�`�C���%�*z]�Z�9��te	sD��2�	W]�@Gg�к7"roz=g*��x-��ߕYeh��?��� Z������!����m^�`6h�T�������*\�Y�k#�>Y��=�{� �
�Rb�Q���B�.k�l�E֐(��So��0zYx� q�iP�!�}ǅM<.�����f�˃[0pոp���M��ٝ{Q3�0�mQbg�"���O�*��*v�m��R���+&�ƚ�uX`�$Z�Ѩ�;�[7����*Q9e]s�~�r���^��'C�5wܛ�h��f�4�x2X@r��|�A��rW��:	.��'[��Q1s%0ni跣�<V�om$����Zue�"m%��==��SyU�	����/C����u�-x+�u1�{$=��
�[7��ꤰ7ʰ1�\:��M���\e�+ܼ=ƞ��x���
XX����.s��˨��R��0ڨ����Ӈ�w��/N�����;�in�V/E�r��b����	��D��+���7����i��.��V����t*i`<U��캵����7�4�D��Y��y/�W���UX8mڰ�ʷ(�
P��I�Jo���K����f�9��Pt����~���W�G��U�V��޽�@
����α����xѠ�UN��J�y���gpz؎��aTPv.VٜUR58�\���ݎ�,�����"��BԴV�İIj�ō	т�^�^�z�S�~GZ��`!���y��;¦�r�8u;訑�#0-�'@ґ��n�<��˒z�+�y��J7����pVY�BS+V�gr�c����.�kJ���5��
�n�Z�:�Қx�2�*)���W�CjuXx��.:�����!�tJ�,G&�!5� i�>�UYP\�o��:��TG��|>��� {PC왬f�b��2�P�n&S:�iؔ"�s?x��s����=aM�B=/��ujx��3����w�|�hRg�Sʎ��tk�[լ����z�{S�6�6��zՊ��Ȃ�ZVvlt��c���g&C��*��2Tc����3��F��
������9V?�h�ō`�wy���~�R�R�ah�1=%�j�\ ���r��i~�6<.�S�;�@X��z<<��G�X8`�j�V���L=W&�����f�����^&3]1/�p�o��U�kf��9���E�����������S��>�
�6��0 ��ⲫ�>s�SJ<ƍ�Ԣ�^Uݱ\,l�6�1U�M.���m.��Uf@r���N�K�E�v8Dˋ4��Ę��,יs��i�ս�d�68��V�;���]=8V�fV\��{"�tܱ�ܚYI��w0͝,�Y��䨎�+oKyv�'VgK@橧6�On�$f޹��j�g^�Jg\_%h�S�.��$�"<��H���$=\�B�4ފ����Z�6⣆��92r�Me�v�-1�6��p'x��2��[�PM�V�hhI�w&�2K��QY��5�6���
c��ÇV�	����[�.u0E��{UsC/�5�pX��f"�TJ����P2`� �9�:��2�n�̧���WŻs [�PWE������̳ʷ�43��nq� ɺ�g�kA�se�9��;xYF�1GB���W��oV���+lD1	9�`M�WZ���';^6��n�zA�RT���zV�����u֧s4�������6�*�
8�S	<�G�b\픵�5���v���Y��Km��7���{0��gzda:���#kλ��'q�]9]F�����]]LA!�.��ý���A��W7��L7������-�����4uk�OkM�xQ�X�Ӌ7k^4VR��D�<L}�>�� �f������<ԡ�prЫ,�]�h#;뤂^[��u M��;�v�p��w�n��X�<��u�����"�^Ԩ��Y��F�����76׹��r�S�T��كi�9�!�Ж^P۱F&z�����hKj�]$F��"�PN;lR�_�Zt紲��4kZ�%,��Y\�m��,���[n��h�k�K������6�U��]R��#|v������7���𞅰��㷳�7�:�s,�6��vm頴��Ŭ�6����coQ���㕴�D���e���c�)�n����e����Ⱦ�1n���d�{M���T�Q����K=]�j�2lLphȚ�Ԑ��ͮ�z�vs_)�u���MpI"���ɸ�DϨVVUE;�:��V*�t�`�s
�V�X.���J�K�fY2�-[�]����c[U��V�"�T\)Jʍh&ePr��c��m�XT��rk�,��ۮ9i�L����j����9s5*���bъ!��.Wb�W�)iQpT)l��m�r]�T������s3��;Mh�31\���ͻ.ҫD��w01����ʹK�+3(�ܴ�\UjUE��ie���0���-yq�g�5�1L¹���Iy�o��嘹q+��b.�ݴq12�m��)l\���m��MM�)�ڥD(ɩ�]ZZ�UVQ�G�Mwin�ijV[qkH�Hh�EQ?�������~9���d��V��<"�A5T��&�A�G���K`�a��ܗ��DD �n�ȩ3� b�`�Y��Z�?f�1h��k��6��ƭ~35M��Ƙ�z2iuE{U)��>���ρ��Z'i�E���Q:�\�.,T�#��n�����6L�r����LA�Wbі��������v.��)��
�X�׊��Yݓ�E)�m�i����_�w�ņ͌W뗨)��
���/jz���aZ�J-�>���M@�q�V�A��4pц�Ӭ�=�� V��b(ߪJ9��{��G��U�4���g�ߩ[�9"R,(־��ᩓ~��1犼�X8�aqѻ�j�p�n��>�7��Lǲin�RJ��X>!�@I�p3Uj1Q�7QY���R���ٚ���I����Q��ӓ*�8�3OH��SS��Q��=���E�y�@l�2��5��f�1Yͫ�E_M�T��G5��{��c�՗Kl�Ԁ��Y��\J�s�s��W�tH��������-���R{lʘ����8�꯫�6q��Dk�z���:n��_@�K029�2P�Jz�JNR.�iWVLQu3�;j��o�ѿ@�Ty�;��d��ֹ��ؔ~pf��t���u�V�4�%:�RS�.'4Sڅ3�����2�K�����`���uh��j|=ڝA����>[�N܉�[����7a{�E��޵ZNuXd���-�����~�5]��)�+)��s�/1�:���|k�{�N �	Y���PWS�w�7/=��@Ǭ��G�<�#V��WSU&U]aKH��;dAwOHqK��b�gA��0dLtR�(�(��aDÖ);��~N���U��E��?��o�}��U@�
zT��=2r�i�z�C�A��,&6��N�W^T���41
sH֌�Ί�x�\k���J�C�g��DVV�cg�ο�gg����)���՞%.��Z��:��`o���ъ�s�q�)��K��
�n���!�D��Օw��hԻ%Jޣwϯ)��:��$nu�W����q��}�Wzn߷�dp��pU����z�ՋIh!>�Hxk ���آ�3DW���Cu\HBX�-������+j�ȅ0CYB���۠�w��á�b�h>󙎖�k)�~S')�DP�!�LT(r��n֤�K�e\�Թ�.㪤v׺r���
��WH�ox��}<ۅ�m�e�T���xX�/�D[��F��u�is�q;e��9�1�l㊬��`cEN�f��3�\d��|(���߶����y��8�����r�:'G[�C�U��PUP�{��s*��Q��,>���F���1U����z�
���X4�~�BO�B���=����o^
�A1�=�^7��
�L(��)�KS�W_z�+뭣���9�l���g�X����uHB��$��/m:
�-��Y~��W�3�3��;�r��H-�����7\hvѺ�4`�9r����[���/�	U�n��7n��A��s�E�Ҟ�.zD�\uخ[�̨�1� kWޙmfw��X'�y׃�=*R�O�p��� Fbk:�0?����k�2�*N±��x*�0ed��n��<���%�,��^��:4q8��`bƇB	� xZE���6�Q�k�5�J��:���$�v�ACK�1r�������֖�dܸP*t�=�OT�1Q�N���� �P�|�bk��f�o���
#���4����~ŨشV����z�L���.��h�V�Lp
nm�>Y�;��[��m�������|�p��63�.�qՊЅmeyS�XM)ht��s�������olI����D��,��W*�U���Dx��SS�s�p-����.���bÇ+��!ŷw��+���?e���ə�Z]�	^��˗;�L���N��鞅��;�-O�#����m���F�c4F�_y��5�4�f3�R(*�X�Xk�S�Yܹ�ܙ�y�*�[��bZ:LOIALf�\������3�RRͼǽ�W�˷}����[��q�W�-AH^*`�h%��w��pˬVЯ:N���E�jԼ�������پD�Kj�K�cf��X]���L�.�+�st�]uԽY�B4%����g��yˆ�������P�<1���(���(�eeS�swp��ܔ�F��̡ιW����)���X�.^\e�
Y�2fg�ʠ �;ԗ���ݡ~�v.��E�G�
��p/�a{��z���Y�^���V�xh���	��lKڄk�esKzwS����z���=�=|x�3����<M����z�-�*�wyk�(u�v
����(9۪xÜ=ZV�qfwd8�{ 靮"�>92��P[��.���*�哃9��F�؇-g,�����"��vQ��ت32l"���nLv��"�u�3%�%�K��nL����諃;KD��@�t^�P![<��V��бٕzf�.g�j���zRy�8��8]��(Q9-�b����4�H�/-�=bt�rg��J�y{fj8yMLUEb�;ɽK/���y��x\��&�q
O�X8ì��>�缣���m59R�L�*>*����*�u����Ӄl�wF���E�
KB{ض�����=��cf5�/o@��
J>wҥ0�a�.��z��֩��kU�8!<<�d����uGp������4�b�+N�l_s�գ�jrX�a�84:Դ4i[�z=�v8o	���� Þ��+kkN��aAT�\���2p ������	�稕���:T�n���B4t���LB��[Ww�-p\c�����F��ȴ��G�Ou��Q�Mŗ6�)�q�YanS�u�X�޹h�b�A(.�*Hof��}zC
�����d,kt^=��y��7W(�.H����� ��u��5�:�j�Q�Ш�p�Ն/-�����%y�p�>�`�|<3��וj�B�x��%�2��t�ٮK><��fUҾ!�ߨy��-p�?�Udyp�'�8?$/="�߻��ԅ��/Ԗ�Փ.��i��%���&kB]S��zSjsxh�`�p�E
��i-8js^*�x��p�ɷ��
�_�.Ŵ^:K��	��;KO��(�/.�`�m�ݥ�;7��px1�ϐX�x�
�mW12��b�T�m9�1�j͘��J_n�+�p�<H�>0kԁ_j�f�����:�d���N���6�
ˆ��5m/
bx�KZ #�bс��#Jw �(��˪��U����Mh��4V��*i����Px�n��s;���whY�U�ݽ�A�4j���mU1�0T<��X�Cۉ�h���J�nrk�u�]��Dz9<<����������`N��yh��P���^nA|��knnL��)��F����{vCi`�����!�&{o�ov�����Fd��*0P���&7��
������bǖR*{��}��}C׷]��;�B�4����"�{)]o^��^ܓ�A]�@�ʶ2~�y�^�=Re˜��s�*�F�%Wc�Ѻ��⪐��]lc��N������+��v����15��������ּ����+F#*T�+fx�����2���(����z���%a�U�y.����G�N	gBt`>C�ګq�pM�25�@��%�.�*^�SZZ2oԪGd�S,�M��z\Ls^0*k��xk�/��P^:{�zA��}�=���J𺿯�Y*�yÌ=��dDҋ',�ٝ�e���J&@�9�L��5���z
��ܱ!{�_л�Q4u�[;,9y���y,`�h"Ä����U�7���G֪��7z�h_{ �HC�����Ȇ˲^-Z�fa�:�F���,۷1q�JL��u B��f����W/� ��${�o %��b#R��։���g�fyV
��MN�5;���0^г�s~�7�l�@�זzܧ�f�~g�WY5f�$c�/�Cͣ�P�*wGh�,_QX�FNoW���#��Ya�̧]�ß/|��������e
�գ�#�8�T��v���	9`uz�A+�G>Z8:�X��#�d�f�{��0�v��F	�]x(7����z镎����.��Kk�x���6������ 0n�ƫݎ�n�C��jbC�j���S�r��liU*b�w*[�@`��4�ρ������~��rХ�=�u�J�t�Ҁ�p��G]����G�!�M�ۨ�����Mg^ltu+X��pu�75)Nը��) ��u=�:���f%�R���y&N��Ξ��!ʧ9%1��(���U��s{"�6�q�������4$`�Ix.��+A���m��~��E�|�jMw���$x���\"�g�
J����p�+=B���YB��9��2���)؎*��b�z�Uq�MpЏ*Utp^��>�`~�f�YDP4x�7`f#�7�}~T�ɑ+UD��y;�ٝ�sK�ٞ��������p��ұ��#M1�7���Mau��ܿg�x5��4�����`��D/�}�/�5J�J�;I�w�oA����|*+�n�(���5H���5��v��Z��R���WO��xR�k@x��^Ţ��x8Af�c'%Ϝ�Ͷ�����d�5�Z���K^5h�\�U��ZWj�}^�R�"�X,�Y�Dz���A�?�V�[��3j�����&��Vp�eBr� �x�Vs���]u�p>]���#�b�i�x��z�1���eY뱛yV �����;eƽЎ����Y��jr@a-������wPcT,^uU�N��y� 6��.��*�j�˦)�Fvd�Ό�\�w�V̼�:T%ɖ^������I����1��9��������+�{��O�I�h�v����tf�M����4ˠ/z #�݂6U�����U�~�,)�D�C�Y����Hޞu�M�ZJ�Π��V2T3*�f�G.��F��`���}묫�0��_uk���Y��JA��T���ǂ%}]yo�����TI��pR�y�x�Y��a�Tٵ(���m��Գ�t��(��SV���o*���#J�Х1�R�]cy��g�)��]B��U�>7X�{O����=��Ɋ�;�ILJi�^�5�fau˳)��Q;{�*禶�K
��X����b���@D�u�����R��'�Zo).���VR<l�ڕ�)��CS/ܗr���%���l���Ql����*9Wh����lP�9MeL6(&U���I��,��Xr��)d�b��3,���B���l�HJ.�]�ȧͻ�H|����6Ѥ��1x�+hf]�VM[Un�W�nJI�O�*�42GQa�X���n�yC���{�n[ l�.�,��U�9F������h�VJ�Y���5�i擮^&���*%�1!��i�XNY�t0�v�P�-5�e72���bT�~�2]%]�lZ��maXNV�)ܻ�O�'F���*kESI���g��Gu�he��B�wb�hn]�*��7!Cf�m�&�T��#]�����+0�t�
�Q`�m���>μ���Nn��ܴݘnT���$U��9gM;[�o%����Nns�B�Xmg+�4[���`��p�z=�}:��{��̵�al���B�!�a��DKV��r�Me�L��P�E���j4w
�U]�Pܪ"cmD(�u����4��32����b��������[��P�U��67/ZQx�u\B�Uf`���
kTqܪ��ܦҖ����W�IKf%b�1�1(�Ws8я��:��#9�dKTms��5WYD�T7)�j�4�53Z����r̥"�̉�ʭ3
�LlX�j�:�������`�B��4��\�V����
.n��1�\AAb�J���7�]n��m+���6�M�����Q�Mnڎep�j��V[QYei��m�f�L��q�Z�Z`�Q�K?5EP��_�;:s��S�wc�C����fhf+͝9�nfQ�|E42Y��}�ζ "�;5v�A�u�����K��7�}E�F�n�\���_���EZԓ�ؿע����ur����B��xMp]�cFx��kt��r4�ֹ$��*uӓ�#��;T��U�|��/�{�8tl�=�_n��k��}j�����>xr��E��C�b��:5�z�ް��[W=���YC�i�:zs��1��ܬi: GW�#t֎.�7}��G����/���}1YJx�d��1��{ǋ{[G2� `F�a����'�z�W�%�.`��e�ڞT�E��IN���]���Ό�s�>�X��YEO%�{o�����:=�$��<NѢ�8��F��=쫵����]L�PS����u��xx\8:����Ԙ��jŪKA	�J��ˮ�o����3�8=r�,��4�<8_�i���,)*p�¯��w��A��g]� XJ�,9�umk8�$D����#F���{�f�/�S�k��؟<.��t�P䛻�o;9$��CE��x�^]T����eN��e���:q1�u�Pe�dJ�ͧ3�\|soן:���<'�H�<�$���=���e2���Ӵ�JOqf����u��yRixSǃ�:��pt����ۣ/t��qx�$k��u�+���ޕX�G�PB�NX�̇9]���ߗ�y�;��|"��.?����Ә�)�b�nE�dJ?nP՟;��a�ZaǕN
&��^��ۘ�^�V5آn�ݳ������=�"-�!1&rSx|+PLlyLws�_?8 �a)'Xe�V��S�U93���=�f2��e
��)q;���B�
(!��z�'ǅԚ�'�<z�*�Ã�LZ��e ߼�n���h~���8e B˝��:Y�.���Ц�b�Y�r1�3vU�&��~�[%�5vbܧ���rUX������r�-퓪Vh�G'�cҵ�7c�2�\�WWS����ڴv�j�B����l�c���?�O�L���������r��)��^]�y�Uӵ�ׅ7��>q�A^k5&/�p<R���C�uJc�%mVȘ6c'�����^��n�>==���J��hxkh.;��t��'�b!��n�Gجhc��R�
���Y��g��=Ax֪�t�9&�Ó7w{�tv�����*f�8$xADj�@r�T���������[�OS��O�X�zҖ_��­k|)x�}�H#�QYF��թ�<��77L�z�j��ph��U�5�᭠6��T�vć�7mI��p�+�d���&��+:�a>Z<wQ���3�m�z%L!�Fu��!�U�t15��n�{�z��{�\�qV�\ U-}��`�[o���: �8��W�����6��+ƃ���&и��i	�+c�J�]X78�f}����\�`_����l����)]"����2ݗ��1�7.���ܬ�qnO�'�Rb䉼G�L�ׯ��89�x6R*k�d�(��\�78eB�J;�O|��yU�C�4��k�O�S�_R���#����.�Wd�5�wP��ڻ���aX���S��ƅx�]�H��k�?K�u�)�լ~����;5&VS��������h��'�5��kq��t�qU�X< ^�RlT�!�؅TΡ�� ��֟4Fܿ+v8��Ϭ�.�l�3�P*D�z�j�V&�ذ���-�M�U��::ς
�*yV%�PKX%�{�����SӺ�@�[�Ӊ
��
vkB�B+ǅG��G�ٹHu�Wu�g����=ёHxpCb�$�FE���;rcJB%�Mэ�ij��Nd8�3"<��J�
xt,JV*�S���bb^�=��x�RTv�����f���l>�����
In&���`y��Vj���ު9�X�c�'{9Jz��+�ZgsQ.ٹ��|�	.�d:�h�D��8����ľi����^|�@0뀨�S|.�$.�K>iV|��N����o�;����k%ʛ��*+�n�(���x�U���L
Ư7پ5�EL���K:ꂬ`r����c�����o��^f���v��(**���`?��ێ���&�U��cpv0S-.y�L����ؘ�L�U�*�<xK�<'J�w/ֱ��a~q�-پ!G�<�ǹZ��$)s=J*!��#�:��|+3Rt��-z�{׏��i��Z�e�Z�' �x����^
BI�yqSx�cȜ����֍��k
��u��-�p ��7ZÊ�H�{[��ke��m׶���,fU(՝��<4VT�F��k"(o2�x�e
��ܢf�S�;N\��p�ʼ�x*��
K��T;��^��k�Q� ʾM,ˈ�݊m�$v�tX��m�V�#y:�i��v,�M��f�d�	�Th�r��̼	'w���w��6����W�*�������4�[o+zM�ύ(��р��Ý&%_��§'�UA:`�ل���D`R�%�:9����N�Ud�8.�ʔ#���P�K+��d�*�8�s��sl�F�pKWG)1[(Ջ'A�Td���S�Ѹ��f���p�Dֺ J�7�L��U��gC�da� U������٪���
��r�;W	6v���/�>DL�Uȟ8�B.�Ь��3�~�c@O�3Z�v�f�u��yoF��JW\�^>�3K��7񫦗
t'�g@LZ,u�(Or��+��X٪�|�R�b���8*�3¥ʱu�!���K<[o޷J�����{UK�_��Դ�'G��Z'�h&V��u�I<���e���F&6z���yN�T�U^$Ĭ(F���~u��`Iy�P^�ɔ&�Ug_�Ӎî�h�rxQ��g&�V+�]����KrD��]-(��:32��98d�ñl
f�fέB�c��rD�s�UTG@kS萎�f�~[S=q��==A�A[��Pv��S�KEk(L�Yx��M.���� �|�l��V��L`�l'�D'V	�k���}]�
P�f%C�����x;�:�<1�
�%��p֤����v�< ���M@4�\mGM,���ѥ^���+R8� 8W��Ё�ú������ш����e�y��oP�
(Cb�Z�. S��t!O1R��d�6D�����D�ؠƷ���*�m���,u�*���)PZs��.�V7&��GA����,0p�Q`�F�J(- r��X���w�yF�
��7���d��q=W�r�=T��pl�7�Z�=�{��~��ݻ������F���ʅ���V��\uR��|���nf�)7�1��ȷ���[�y~�ؽw�⺐�n�eeK��DeH�R�i{���4{�>��.��5/���;5f���[8��2�̓��UO�L^��8����b���H��`��5K�Q�x��*s4ѳE�S�"�Uf�����GU�d*��a	f��W��8�N�>Yxe�V�Nˉ�p��\��L3�����b�EaK�l1�w�`�f,*�QpL_c��g�x��h�Z���3m��yݼ�,��f��x.T���ޮxh�壃���f�i����f��b�1z����P��]zjŕJY�S:��,OQFu��#��xh�V�7ʼ��0h��,}����*�o�>�=%/A�\�J���4FTš׹V��,,�½��g�I1�@r-
�|ԛurȆ�7QQT�BU��s9��x��Z)CYH��tJ�&#���
N�/b�=��#D(|:�ee����f���A)f����Z��t&�Fĭ[�f��6����"�"�1I������5_HJ9Y/dglA9�ٔ_ol�=}�l��.�ڼ�m�<˅7'꯾��[�����}Y@��}{&Ss$)�Y�T'��Vr��wt\ӳ�^=�L�4�D�^�vz���؆/6])�p����Kw䒡����ƍ\����Q�n��gUO}>^>�"�^����:�9؜�F���k���T���b:�P'塝�ܠ0�~�R���|͊�M`}/2��ĉ�Rϥ%PP�:R��*5X���m.:9�ݞ���S�e˞��*;Cn�rU��w�H��[���;1�9�7T��%�Aݧ�tm^�=�As��\5� �9�yr$�����
�sJ���3ގ�ݻ�g];�`9Ț�;�;S�zp�R�;�x#D:R�����
cP�Q0r������z�.O>8��sFrq�'���N�P�ʶp�)w�����Kyy[�":n�8����U�k:F���z�T�K�M�U݈"���7=��c9:ͽ�^��sy,N��/�c���{N�q_I�~����y�����n����TO%��:��tF��X`�'�@7������{�K��D�P�p[�w�fӷ�b�
��]߁Cz���R���c����:� �Z*��ː��$N1�	r��;-&�
+���vL'�~\Tx�<)aʥʼ�xV+�������#8Dlo�WC�+-_�v�}.�V�-I��B0c����_�g
��b��
Ѥ�c|~��,&:���T�`�񨅈�Z����v�� wk����O �pખ�(�Z*	ih ��컎Z���j��5�Z S�ʗ���4�7T<8*��3��t������5�o���ú������0p�z��B-�Ta��l��I�N������g���Ɠ�(pUe�^0n���J�XOn;�6���
�����\�+&���k/�³th[��X͋�o4��X�����pl.����k����q9P���h0��X�%2Z��Y]Fݷ[òN��ձL��۽V�x��WV�f�9��3h\���t�;�P��ǬQ÷��V��[*���Y�N��|��yܶ�bh	�9.r�F�]\����$q�����1|��W�Kp���ɳ�K�Fw)�}s���ǌn�=H�r��%�O�I�鷿]kV.Wv�Ǐgeq-š�6�\���z��^iV�]�t��Xk��κ$F�N��*^Kd/veȌˌ��a^G�DѮ0�8��H3�w��L��:�g�'�Zt���eZx���ݺ�����7��z#I�ٱ�z�r��b��j�Mj���XӼ�]a����jp�$4-�(���XUf�����l�qj�i�J�ǜ&�]+f
Go:ӵ��c��Z��b��}n�K�SѼ�n�-Ko:��7�Wj�q�vd��d�ȫV�.ù�����V8�7YRBV/�
�e� �I�^�j(3/���
��ց3!AU#>�M4��@⼋����˻0*8��e���
����Ĩd�H�����R;�(�ʄV]�̻�%2�G󗐧k��}i�#m�r4Mc�xF�����yi����͇����J�g���NŐ�U�^�[��F�F��#��)`�*��B����s�G q+t�wc%4�H-ŉ4I��`�{�2�Sm�9�٬Y1���v��9%M��Xu��J,fV�(�t��+��$�wˎ�u*"��X�P�tg|�����+��mm�m��4l^튌�+p^Y �xh�kS�@�y���9��d�S� ,8 �lzh�G��R��ʆ�e��ޫ�ɰ�dp�[�㓛��1���`ɖ�
}��M�o#66�ږ%�Q���A@PQF"��9L��i��.S�(�3]U����YF
)�10E���Dv�*eT.�Z���Յy���r��.eFm(����E�ʊ3�.8*��3%��b����Z(���LsJ0�bԸ�HV�[Y���F1v�ԣ��n";�1]V���IT��M� ��`�QE�E̘ۚ��\�S"�Kh���2��Q��v�Ź��x�&�h�e1(�Z*�+ƌU�֦r�U�7,Db:�����bcf4��QM�[�D�Z���[-aR�U��Y�45�\��͸�e+\��lU�S1���m������ט�7�Vl%I��n+ޢ��ʚ��.&��Y%m��U�r��z=��\��Rѿ�P�SS�z����d�1eқ��5W+�Y5�%a��2+dʚ�p���^V#��Jb��+�*���K�=@Zz+�Oh��jo�@`�K�x�7ޘ���&$�\�.o�tɅ����|��B�ܘ��zS�^�\*�=��u�	C���g��lX��t< f���D�ʖm[/��cc��gM��x�ݻ�WX����X�.X6W�����-��-�ʣr�9|�T/���:�αAOyU�TNP��%C�qа�z�ʦJ��R�C���sl1|P�`����h���d����8�KD޽+՞Q��?z��t���jd���9�#���;b�zl��si�����_��CɎ�b�������u���pGn!˳,��2�j{�a���4��Kv����|u�+9e�w�ftgWIۻ�q�4��څ��������G�1D���+��
�bFS��}UU�{�U�R��%�ҹc(�K~}��ke�Z>��t���5[6�0KX'��{�`kʋ�����P_1w2�K{V%�S�*ϝH�S��0|��Z4�k��!b�-Ĵש�����b��yq���TMqŞ��R?_mߨ�Ϧ���t�.����G��t�8*,9��m��a�n��OU�Y�C����v"{���D�: ��{k}�֧�*��ڽ1S�k��@�b��Y](��ۣ�:��Øom�	�m��j^m¢�F����0r7�����:�)�v��sYp9�ֽ��qIoH7�e�X��)e� K?e�`����a��	�3��w����k4�&=B�a#x\�A���Ц�ʞ�Ӭ��p��k52/�ܙ��j�1K5T�V���k�N��O����Dz����y��Z����r���\�ʬ�?#�̥s+�cݥ���'�LQ�m]ے%�&g>�:���@�&�A�SB7����,sxK�f�;��wn%�[�'?}���<���;u�1ڗaʜ��9q==4d���>-1Յ�!���t����Q�!�"���+B�8�J�H)�G�����<>�J��{w���8TF|�������V�Y��X�BfV��7r��\�ѳr�s���+����Ds���P#Eh��6w�Ke���p�V����R6�!J���U��+������H�����f��6��x�諡�BX��&�n��Wo7��%�s,p�D���Sv!6-�X��s��+νݷ��<��'�.0D�K�*%L��Ѿ5�:*����Ғb:����X3ki��!�K#����/��^Z4�C���t� �p4�^i�ӌ��AEK�FM<��ѕ7]"pH)��U��m0������10/��9ݦr�h�n��)P���k�7/t��)ݵx�I����LMjh��;A͎�/�6�әY��B9ΥF�tz���m��<�]��p�91������1g+�d�u�~]^l��-v`Zg�=�W�3���FP��E:�@*��kԥ���+�n�����C��r��wn�R��G ��ٯ$�(�=��ǣ�
����V��A>���q�S�K��&�\s¢Öz�k����W������K �b�8�Q�w�����0�bc'�uWM��l�����#d�ft���<YAC\��m8��c�� 8&r��
�pxm�%��6X���B4�)c��̬�
�Z@�^�
p�9�����B�m)$,���vV'�`�^����\��E�)q�]#�%y}��-I��~��r��bhT^8�I�V:Ԇ�n%���XT�`\kկW����H��)���Ұݺ�q�J%|�/L�8� �sֺY�M��܆�8�IP}r����P��_V����/$�fT:5��r�I�>�d,���K+ ��[5��mx�zx4����P��`����*��=�@�}����R��F�b��#N��xT���u�}����4�z���h��p�P�׆��/k�������_ʠH\�����_�� �^T���4����`�υ<��c�C��_�Q)�ߥ�C�lt�l�Ɓ�5�")�#f^,�ҹM����:u�9��\�A*�t�6c	��(�V�P䓭=۾���ׇ���<��r��wZ�ibT�âk���t.'C|}�@�\)pu~�-��]U��0��R���L��g����ȥ�{��������	z���v�Y�Q�&�j�(E������M\�����$O������V�Y�k)o�"�1<��Rd�ٸ���˾���Tᥢ�,�MN�W��W��tb��#��N�&�����VYfVWv��fn\/;g_j�3�uT�Z�(\s����珛�
W�Fm�B�0 4h��Q�HK��רV�O&� �>������֭v�*�U5�C�_h� W]�d��7��l�wo{v��VVל��1_I�S�<;>5AbT���Qy�F��׺�ߝ�Ċ|ur�~n��F�NK,z͙�g��\R@��d�{f���C�*Ы�X$��kB�5��t�������>�M%
�:9;B&�t��N����"[��O����Qmj���N۵�/w�z��������C�+ǄF��@)��j�"�f��:�ڎ7��+�V��!����t��j��5�� !}�Z�w8pc���jY��b����Z�o(A�70�*�b�hF�h":S����䩡��_@��U(dR�r��Nn�+�X�yRŎ�T���bx�����(���K����{��ܘi(1�v�L���O\w������嫛�(�ۙ7S��Y���@�18��� �"�Ns��g�:��r\�=V���&+�-��1P���֝�h��	�����J *q}o�V��r��/g/"n m'��ݛ�Ȏ��g�S'x�Z@���=pAx��������{}���X<8}a���W��t>�#./o �j���6]�z]�TZmPT.���f��_��:�d��D��,Y���[yt���*��3�jb�����O]0���T�����Jؽ�����gB��ٱ���4�	L����2����	-z�w�1پ�
�����LXUH�/�σĨ��e��lF��#�q�S��Dφ�P�/�RT+���'L������Z=��IR�!f�|�HW�h�g��#�P��Z
�)\)U���֞ܒ��*n#��=�{zN�TJ�9�PMV.Ε�ʥ�Xn<��xmö����p`�n^F�#f��.�ޮ�1WF�\�D�r�dsv������Z��1��koo8�,<%�W83@�Fur�}�rvu�s�&aOOú��J墀��Q�n�!8??����"�g�.igU��ū�c��]ڥB[�f�*����Ġ�Y��3�}ޏ�e�K�o�n���Gx���乃ծ-�4Ee͸�ut{J%�1�{v��؎����
m&�츋R3Dڣ�����=��GC����/�<�����^�)�W@�Z\�AL:�=m-Jo)[\�M;�b��S>Ld7N"%��������E�X�f�����A|�m<����Fq\�v�}ټ�o!���@�(�ͽ8�s��Po:{�G�.�F���ٗ2�Z��7�s�I��g$�q�e�����ӗ�wqo�	�߻%JK����bW���ݓ4�kY��Ego%��urj��S5`Ku�)S�{�U�Ξ����$ݖ�ˤ/=Y���ˁ�H{]�⊎j��y���${Uw�v�{F�@�O�	�{���N���n�:֪6��D=��6H��I��8����\6�>r�*oS��}��F'w��T'vq�� ���~4���1�&Ҧ�<�yCޔ��ҫ����t/ֻa��L��i곋q�V��n�Fj ������!����m�3'������g#,�
��yh�����&�+�pi�n�N�M��.j-*�c���CSyȵ��򔮽<,z��%l��NvɫfVS�jt�eM��o�iIc8)�M��s��[�g*r�dy�{;w�d���.(�eㅍ,ns��nH��'�z.Yvm՗����mm�-9f�"F��u�ڕS���̨*��<�)��y#d�LZ�0�]��Ǣ�ʹ�Pi�:�k�I������mO�Ю�g�t}�k�/+�0%N���Ż�{�f�:O>S��7�	�ev�D���OS�x�bT�<Q�7<���~�#��
4��)��O������{�u�]��n��������v�7-t�Tk�m�Z�dV[]�����mR�aL�?o{S�~��}}{���Vǵ���N�F��(�a�h躞>\�"&��J/4�ܘ��z�\N4 �Q�ͦ�}F�o'r��5���|8nL��'#}ti�pPiU�����Mpw�%Ko��OEY�B�t� Ms�������vuhj���t���,V��|f;rm��KS�lf�v v�&ѭ����H֕�mI�m鳬�sC�p����:�Xb���;Y�J��(5�WA+"ȻY��n��qr۴�u���G/s`��eJ�*���Өaw�M|d�]�DV՗I%;�6��"oNø%Y+z�wH�c��\/T��t��A8�����,�7�"2����Cn�A� ��.}�rP�(�ٯ7�˳i��2���<\ڣ�'r�L3\׷��I�ە%�{��^���bN����s���m�y�g7r�K������;7t*y�!����\(���� ���6��}c�	u�>��h$���}��!�#)wYǃeۣ��W�N���s2���i��͡ˋŎ�[����� 9��8]�K+-��	M�S���[�I� V �I�T�T��gaɶ���X����k<����ʦd��¼�r�Y��/	���C��:2�L�$�:�2)e���t�CgfU��LD�7�6�A�]��h]E-�h��� �,�p\�b�V0���6�(џL�Z��b�f٠odwt�8r,�ÂXU�����A���Vy�J�� !3V�Ѓ�J��[ǒ�-�J�w@�� �MY`�ƽ�3p4`mKA��m�-ۄ��u�LK���.�7�۬��Zto�׀�h���se�&��ir�*¾"�
����F�{״:ˣxw��m�̶kU>����`�BKt�7�cibo���������\I�����+%t�hT��4����sP]@J��Qr�{F66w�ׯ}�z�������`�D���,�ui��5�v�5�ʪkn�0��Q�(�r���QQ��f�h�4R�օ���J;�\v��:���^\jX�EZR��
ъ���Q�������*�r�Z$�f%iZ��b*cn4�(�ҐJU��3.5+�.f �q�.9�hcpE� R�m�v�QVe�V���SE��.��v�c�+m����b�Q)�E2ٍ��*��TaW0DlU��2��f˩Qs%˗b����i�̢[h���dPƈ�Eԣ1kS�8�PQ���Q���-�"���Q��F�*b�h��r�([e`��K�J �8��Z6��Y,B�Rƣh��eR*���g�:��Ӯ��M�e��M�4�
����`3y�q���K��<G&ͼ�2E7��K?ύ��7�`ʳ�w�dwQ�#�˜æ?K��5B�C����t���Z>�>n%u'�ƈ2=�^�I��T�M��w�9���pM��r�q� �b�7;l�wg���k`�8�52dNo�N�H��ӭӓ���po��A͊����r;*]m�iZ'_-��)
e� 1�����_c�it8��F�x֭9c��g��3�&{�yk�pј��lY]2I{���̲��>�G2,&2�n��07'p�ո�����=�,ө�in�]Mu��N�uw����7���b;��hGbێ��d�ࣗ��u����q'c<�Xȣ�����>B6@�X��y�������.iѻysB㦎���e��T��-nͅ)+�w�^�Voyĵ��M���D�,:l����
ήgzT����Y�4gv�����)����{&����u���%����%��~gv�oH�ojQ$�U~zdTt���A����M��k��2f��-����rє�S'�T=G��S���)�Pv�I�飶�.��&-�΢\ۛQ,o@�ݔ�@�_vw$����Ǟ9��s+8�/\�qҫ���r��dW=���U��>i7���({�-�[���9V�M�h���z�ŗ�v������/��[����O"�lv�tB�N�Y���Z��D�y���q���ڇv�a� ��q��y���f��n��H�]GB��MQ�����y��/YU��%��f�,a����Y9�V¤Q$dr'�nj�z�OE��
�fZ�T�׃&^��&�pzDE��K���٨�։��vr�����^�}�iEۻi����Y�1��с�y&��\�gC+rN�45���{sG�3$���ĝ��*L	��1J�׊�4�A�����g}If���9.��}�*�� ��}�'�"���/��'˪���!u���h�xS�Zo\;��-��8��z�%���J�ς��bJ����ª����r����'^o�;�Ô�oG�¡�߯j���͠1�W�T݁�5�dG�{����|���[K���$lEh��w�A��j�[�ఞmO���*b��t�M���`E���#M�;"��y�Kw+k�x<nL%���ӎ���nC�#��ҫ`��ٛ�Pu8t�����v&�0%�>�PMrQQ������B�ݙd���.�f��+��6x��Y}�kz��g��O^h�I���D^tص�3%���i��n1Y��jQ�|�;ˎ/�-�9����r��O�Ս��G��߼uVֳ�⹷g�r�aRp�DTؐ�ܙn��`�7�uZkc��ɽ�3�֞Mش짻9�N�B�"��Kԫ;�!r^>��ktm7"��VQB����~�.r�'���<^�i�[�ccS��MV\�yj�@�,�\U���o*�$�9=n��2)�$&)�sM��ei��-,+6�G]ۨ���h�u`R@z�^�Gp[���پ:�s�*Z{�#N8��&E��n^\U1��nƝ%�
b�4��k}�?���Z{��0t���[f�w+�B6��>�*�48�}Qpm[�3�m�Ūj�Aד�'�m������ˡ��/�(?��G+i�5o'���1ĵ.�ީج�V4=Tֽ�/�V����W�_ʚ�FN��X��T�2����������F�	ur�Q�O4r9vܘS���˞ԷspWs\ϲaY��(�M�*��)���8e�"��wJ3���8�|Bf�H�fHL������9�j���Sx�~�=w��]	o;3t+.���� l9��hڀ�f�b�BbP=݅զ����s0�o��9���\Xj`N`�Dݨ~[ҫE:0a�O�)��^�)}0b뮡��Q=�d{��y�����Gx�}����t��AaC�G��)/O�E�w�Bcx��0��:9�GF{���J�N�^rm*ӕ�a1�3p�
� g+�c��<2j�S}���V��ʑz���Gfi���~���-�ڑ��S[	���O�~��5��N�>��^=j��p�z�)�ծԎ�ǆ�a�*<��a �}�u��h�����W�\]�@͍�
R^���D8��4/�dr�� x�-�+�Qׅ��\�>������,c�w�C)cOc�vO��^��e���	�Ǐѱ�}��@���U����^Y*򃳧� Z.�
W�\��9�X&��;�2t	��W$(?D>�h�ك��>r�D�ND�M3�c��Ô��6�ɤUv���Z�W�m����fk�Kqg��ޫ��^�]�]�-h�Ӛ��{yh�f��dS���ŋ��=��򥛧Rs�ڋ�N���vټΙ�ع�Ƌ����G55Wv��f��ח˅i���}|9�1�������=�/�'�1a���#t�$bY����[���&�vo\r�:Uʥ��gN>]hM9f�X�����Ӎm5��U�l���I��ʑu�����|f36�-q���I~���q��E�b�z}�
���n��~$��v3ARM72Y��iʚ�Bwy�����<��gĿ{��.�H��.E�q�r(���u�6���fAۥ6�^���y	��$z��:H�q �8�gg��{�!m�4#�utw���!���h�f�G��Gj��K�a1)��,�2��9����9/��^�h�~��=8pl�0����>�Z�k�vy�M6��N�ڷJ�ˮ�и��	�N��v�ja〹�� ��y�R���6��>�+�G��z����uk�1�V=8��,�������<�:Vʫp���;��Z<�Æ�B�p[�W��4bN�;gqiF���/�=,�4m�m�8�*2�eZñ]��Zh�7��6�Q�u"���K,�wt�\]�q�fK&�e ��f���ju���4��������KC��P�S���]�jd/������[r�Y��F�tыc�&�JM���P�S u�-S!��?w���R�FA{��V6����$4�gLP��W�,�r�M�f���p�Ѭ��VQ@���ϮC����{3�W�ͷ�����;�%��(��ۺxv�y}q^O=�Fb��vB�;Yp�� �]��m+�8+�˶�5�R�����D�lZY���wSQ����ku\�2F�d̄��{���g�sȫA�����~�mT8%ף�j�N_D`�U)����YRl�V��Ο9�.h����X��AF�J��t���J!���sw�s�mc�H�V;#v�ҭe�s5�/l6q���,�ÛlJl�$A�M�����2�J��5-3yrm]-z�P�&u��Ą�-�j�rbFԒ�K�������̌c�9nSrN�V��g@��l�ȧ���On<�QX�CS����Ǳ����;�2�u��w�x��R�e�d�=|$G�60�P�9�j���=>x�i��T���-8kV�ⶶzyTb��r���p┙��g�M�z
{��Ӊ�Q6�fwA��SY�����X��syq!t-�$��!){���Zx��V��O�ib�L�ŵ�y뒖����cِ%���
^{p�#���������'����W��^�~�v:�
�Jp���г����g&j�mf�7"r�:O����
�S�����d!�Hۏ �xq[�w���Wp���WS\3�ڜY�%p��IXj���1�ۮ>�+Qܻ<��N�[�R��g.䪝Y�r��g�tC�Yb���fgV���h��I(;��tW5,姺ir�J��� ҬhW=���w]j�����]����l9���6�Uo+D:���c�Lee��.��3l9,}������ty��gE��57k��4�����etޫN`sW!)��%s*.Cj��[g�)�����D�^���T���oV��Rq*�b���5����뗐�/G%A�����nL��&H�<Ʃ�tpX=�΍x,�JO:׻.�B����7agZ�Z��՘�m�)k,��\�f�%+GGo�3oHi�V�묭�+>y��ω�tm���z$ܱ�o,�Z�$����ι{d�����0S�3�9d�v�۳v�m<�G!�-�0���b�ѩ�u5��Vz��B���ip�-تB���_N�¥I�4��$��*�{ ��U��nj�8��w������3J�q𒒷2�RK����X��;�}���A��i�6iq�v�(#�OO���Z"Ns=�-���݆�ڙ�;�.5(M�3kpZ"h��V��1ʃupa�7efj�y;7]^��q+��%�jP[
\��2���{�;��bk�^m�5R�XLh�8:;Y�ZݴM�V�Ճ�l=��;�P5�W�V�@Np�MntǗ6��|֡�F�&	]X��Ѧq���%p��������\}�B>���9�ӥ�-L�Ž�(�
J�k*�;bsI����"J�:��ǚ��K�t�z!6��Ş��s��lݍ+{c�56�К����c��)e��![D��=���fq�վ	4��/"5�ɼ��t��:��]�;x�����!j��?*�e���ܴl^�}u�"����V���4I4�P �6�-J)�am(�a���[Q�"5�5�*��T�js
eWK�*&n*�j��nmũM5�fm2�J����Uj��a�m\�r���F�������s]0wnZe�b�-�̥�W-��\Ey�,7,�8��^m��Q�LD�V�s�S�e�S-���A�S�sl��CR������m-�˓2^5Z�kE�k-��i����U�ջwe5(6��J<���nѧ2�Y�u�b�l�Mq���s)�m,q�)Z��A�Q��h̥/.J�Ub)Ƣ��x�
���X�Ƣ�QEUQ6�f4QQ���yB���X�Fү(�VQF*��5��V�GX���R�U�����B�|RU9�»����:�)��LL�F��Zx�p�:�����p��!�wW���qlΑIs�j�I�^��e��M�c�/Z���&{���,N�X��u !���j�U�uL=Ӱ�ȝ'jӏ���N
�[���=^ލ�R�/K;*��s�k-�b���=�=���o����Oӱ��]l�]�.���k��uT+�5�N�Wk�?$�s�fnB1�k�T��綋��b3xx�9�����=�m�B(m2�ps�ٖZ�ik��hE�u�0� E�Z<z�n������uet���Zw;]��gC�3�Ȍ'6+��7�^����#�R�u��B���k�nmAl,Z�K��q���rQS�R�G����j�.tUM�t�z�;���;(�ڰRS���GmZ�܏c���"�5��,H��=��#bx���t;��̼��6��}gqO�%�t,}-��~Yh��*L�-esT�&D�~��D��@�Dz��YtW1��gj��˻�I�6�K�s*7����D��̫�.�ˠӑz-Ÿ�#<�[~�)��\ci�2\�v[���՞�]+/D~GD]���qv��]s����2MEa�YL�ׇ�B��N��x��QI�B�wR���h2W{VJG]MV�S�p���}FY��湶��Y��Ǟ}�͏�wq���#����j����{j󃚊�UeY��Կ���� ��MMY>7�5�.�q�7ޕ�R{��Q�vцu^m{U����p��Ώ�[7�.7���k�Sj��v�k)=�eG�.�C��H�q�ŭ)Xsj${����F�G ݗ=͈�i��or�n�Gq��W��(y�뀲�=�Z{u�9<�z9���7��c��:;cRgYӥ$��
�[����(_f���۶��Ud��i� ��*dg]hܠ��U�#�lUk[�X�Q��|}�y�ocDP����]�A�ޔ��{[�<���wc}�����{��Mx{x��l���9��)��!��O̤*��:��z��>vh�ts�Lbߜ��U��N�}�<r���W5�ʌ�w�;*j����{v���&�����b��J��0̄��kFp�qS�2�N��#o7nާH.��댒-XTS����B%s��<��ضvj��V��.�!R`��z���u��sC�M���͹%����s��HBn���#�	c9��^'�ª�˩��y4�Z�;}���a�G)
�������d��:�U�"ϝ ��)`�@`
�]�/��:���Qu�b��tH�w!أ�J}]�kq46��]�.)��.�.�>[^>�����Ys7�v��sn��C�9�l!��lf�M�쮆��'5��z�[��2���n#������)zMAz���}y���s���p�t��h�c��W\-�櫎.+;u���=���^����ˠ���Y�'/RE�ټ�7�Kz�%m��ӫ;P#�CX��������"�mv�u�L�R6�-]�֜|�Ł�|%aKtNJO*A��N�_�Ľ��&S�1Ʃ`X��Gy6E:�wvn{6������f�_A�z��tRj�w�h}{ٽ���V���k )�����N[�U�";�b�p߇UK�Ʒ/�w%ҳ��.0����Gk� ͍�h�,	c���J)�ܓ6�y�y��?E"�_�L(w~f ;^�o���^�ε���o��}��'�-��^��^�T>��.��}d�F�qr���=oW.Yz�L���GG�3Z�uJ�S�GX���2���j2����mE�N~N�B�v�;������#0Vi�����#�q�:�_�J�@�Y�ΨE��%�Ӟ�;�r�h7�1�,��*��.lGeh�urҼ�K˗;�L��y�\�m���q�"bi2Kg�4�z���+d�n�P��1�����ߡ�|闿q�솤Y�ܯAZK���F7 ���@y9��Ƴ`DY�՛h��~1�UskוV���2B�jW������s��= ���z���qt��7�+`B[Q{����� �#�I�|�'j�mDN	�S�����7��A$���6;�}<K��^�5o�F���XǛ��^_��N��Y�6y��(��[�*ǈfdm�����TÔ=�:���������Jg��L.���RYY�TL�&PX��,��,�}�?=^FՂ.i��V6Y��u�4��Z�[�®�R���)�.���{���v���	C�����={�(ۈ���m��ރ�8[n'�8�egIe�[(��ي�v�0�(���h��6�o'csD��'H����v;1[�{M|�18P�j#�'�c@��ʌ����sC��J��Me7o\u�/[����Mm�g�n���Rk���-���T�N���S��zF^f�����g�L��ny<��T[�Z��~�4.�	�I=��#J/�>��ᶼTo��^�ynof[Q͇*Ƅ:ۜΥ"f����f%���Y��UE���ˣWzn��,I:��5�t��Ĭ�}օ��L!K��i�ՊAG�{���SK#:p�-�(��N����9�m�n�.�T��:uu���N���ڥz����I�i�a�.V�H�awH��:�Y��9]��*t��kee:��H��.r�5�(�Jf�� ��Ϋ����t�kӳ=��,������n.���F�{��l�I�u�����j�V_U>OY����ә���R�mcϣ4o7�3�m��UG6�^�s[c�7��ꁵME�N�
DQ�z,�Q&�b�l��`:<��T�y�*�6߀����.)U�n׍�����?*�<�|����S�)�2WtyQ�3sۉu!7=BǢ�O#����`��N����q��˜|�U�)=�Y�C�(�n�9��6ҡV��Tײ3v^�cE��yY��|c+��:<V 8փ�F�b��-G
ƴ��fRk��U@�E<-�xθ�q���'�L{}�NrD�#RBzs�g+J����e��_��XnP���ړ��T�gn��T�i�z�b�,+�~-l�z,��36)�����_J;xr��F�k��a�<��Q�����I#z�1��^�1��o��s�b8��.�fP�֐�Ь�=��U��f�Vh{m�^����0/�+Q���|�U3B��)�l�Z&����c�s[r�>���p�����p�׍Uy�%��'�Q)ל�vU�{o�Gו@��"R�ql�������x�P%%�Ow A��n�����(��}Tq��P]��޵˺)�謨r��]Π�Zo���R��c��&M�Ωb*�;�Y�ͣ4��h�Յ&M�{
�$�P����ԭW0`�h"Ä�#c� 7��b�9N��bJ���N���ڀ�`g;}���a�Q�HɮAv�g�@�h�Sg<Һ�n�V��F�{a��U�m5+j�i�X֩�����(�䛃�A���[ꔧ����I��}Q׷�+d��u�*2�^�O"�cuݍ��y�PK��j�K��HY��,�FfMo�ޱ>(gL�(V�[J��>u�]y�4Y���z��^8ܪ���E<�ݒ�3�ֻ$�
�dUSl�'���w�[��\�Q���=U4A�=�o��]������.�_~��_�_������V�����l�� �4���� �ؒqP#6)3��>D�F^^��L���������}�J��4�$�"!$$ ����7��=��d�hh!y��WY�`�%�R��I���	� b4�I�o��lm����0ٞx������B&qXgI7�a�Z�$ZYݙls��a�$�Ra�E\+�L1QP>���u�Jr�����UP?P��  	��bK3���E:��k�X��#��w�f�#�W�W�H�⢠_���s}]��@�Q��q�%y� ,��-�� o��F)�%Y���)@���d!����<:��Zt��fJ}��1 1�eP�*K�	X�(�� s�D���1b�
^�"d�������zT�6*�f*�
* &�������lSG�}@�$�7J�LbS^
��y�O�dy���<[~R4�d��W������rkni�N}��2�$}Pn�	M�d���˯gBޮ�T��{]�f�����|Os���"�n{b�|yC���U/v��D�$ed�!��U���* '�����O|'|�D��Ɨ#)��s� Lʏ�c�M�X�8��p͙��c@Z��.��Ti�ĞY$u��`��{ r~�@�T�-����K�$i@U a���<1d�"�E<��>L	���q��>���ˁ�#`����L�n��$�����s^Y����'�=��zO㶆O��$"�z��
�8G���+����}* $�ҡn�.��=�ǆg�zyd��G�35^Ij�6i#�ք�	�㜺k_��![t_ߴG���/3��]{�j"�v�J�=��)�\�Y.A�H�v.� ��A��IvZ[\�PY�T^��|	
� '���c����<��{5UP;c�oH4�r�!�Z�fKr��7��Rɩ@<��!{���8?�]��BC��