BZh91AY&SY�ci��_�`q���"� ����bD>�    }>̊HIEKm�V�KCD �FUe����"���-��ViV���l�Z)Jk�*���%%4�٭�Ub���-���M�Z�}d�[fl�Y�l1��E��fT��Zб���Z�l�h6�*�k)Um�e�Y���am�[Bű��f͡��mz��Z6j�ڶ�jX�YhlD��5��fԕQ��eQI�il�i�ȠT*�
i�V������E*��f�Z�[e�ڬ�i��l���z�U��6Q�-�  ��b�U���l�{4�{ׇ���x��.�-Z�9�z�]�n�W��w+�]�u�*��k��a��j��ǻ^�gTݙd�[C����M���ժ[R�fm��� t ����)JRޥwM-5�^<�T���;ӣN��+zYҪ�K�xw�<�R�{����!R���k�Q�^�ǧi�%�m������JUJ��J3V��8�͵�b-�4ͯ  ���*�EW>�ԕJ�I�k�m5+m�{Ǫ��*J���ܽiRT��{�W��J�J�Q�I�ԫ�<��U��Ϸ�<�T�K��w�T��(N�իRL��k[VRfVV�π ��|z�*oy��r��iV���{_)U �}��}�/�h.����J�*��}���{c}���������ޥDQw��޾�E/�U�r���I�{�+�]���Օ�Aj-c�&|  ����Q@�k��ﯻi*��Uｵ}�G�٬�n��}�����b��o��R�'>�w�YTS�+���T��7����Q��[�yo�/{u���m��TB�MgA^Ձ�Z�2l���W�  ���R��+�{m�%T�*M꫻�R��%g�u*U5��;׏={5R�)o)��7L[m�z�ʥ*��+z���r�����\�W�R��.zR]iR��W�,��[mk-V�5�������  �#��h�}�{�k��*�j�W�J^ڪw������*����U�fU��z��j�z����W��V��
����Z�����ti�^�ֳed���TԋiU|   <����ލ��ou��޺� =��ާM�ּz�S������w�4QE޽oz��]��란Wz���� /%�d�UCf�	���[�   o{|k�`w��� U�.^�V�=PD;����F�,�=�֫�GOz�Ǥ���qZ���w�K� �h���J�9�:�M6fkh*Jٖ���W�  n�TU7�.z��z�pt^��gEP��w� ��^n���w��w�QC��8���åz4<s��E{k�  
   50T�J0C  &C	����%Abha �2��RT�      T�URh �i� �@O QT�S�S�0�P��L&�R�ު�dS�ѥ���聘�d�?g����?�����UV,�\1x�u���ٕ������}����ϟ��D U��y�D_�?Z� ��"�
��p'������O���
��Q�\� *��>�*|����?���_̩�Y���p.a�W�>_� �dѕ���9��!��@��=eYC�@����!�z�����������!� z��I������0����+� z�}�=dY��W��@����=e}`>����+� z�������������������������������|2���� z���,�� zȞ�̠'2��z�"z�(��ف������P�������P��D��P���eD=a=aD=d=a>EXOXQYYE�AC�Q�C�PC�C� C�Ȉz�zz�(z©� '������������� ���م��P��P���=`T=aD=aA=dQ=dA=aQ=eE>��L���(� � �����������ݐD����T�PW�P` }`E=`}d<d�ES�P�TS�U�S�PW�ʧ�	�f ��=eYC�P��=`Y�G�S�A̡�z���'�!�zȟ,��'�"}0�����L����L��}0'�� �����
zȞ����0�����(����^��I���_o���T�g�2�ͷ)i�`C��e���
.d�Pڹ�+%Ů�=򧻠e!��67-+p�zު&���d��͛I=�(�GH
ڻ�/0�{�0���{N�����qmf�?�+ ��3g �N1��(;R�2��Y���#!bd�4j����&,�
��3oq	��ʿ80��U�����b���Xّ�sP3mR������aM;���ֽT4��K�*�T�;2Y�7�hْ�h�v�PqVY�� ^ȝK��eh*���8y��6��1p�ҵ�[V�+UJ]�]G5�$�z�Q��+i0��d�p���$���q���w�`;�(PYqk�!K&�eMr�tm�:�^0Q�C�l\�Cq�29*���QoB�A�*ֻ�bs%���1���ov�3U!#�pjt�Õ�[�']CsZ{�z7E{�Yq��� �u9&fѹ�Hs!�n�l�[�ӥ�=w^IXd1@���	�чm�X��S�)R�@ݽx1^1M�wj6n�%P1ַ���(٬�Z��[IS�	�4�-;x��Qr��6�\�ӛ�N�ۦ�F@P2��ca��56TL�/V,1�M��y�i���i�wF�ib�z�jJܩ[@h�;��f'GE���@mf��-ъ�j�A����0;��2¦ ��XYu�L�	zè�w�,f�׈v���:��s0�Q�D�gp��T�P`�4���(���#WZ�4��̬b�-h�cY[K�сZ��3eLh]t��d�¹�J;�l�t���4��F���6am+Oh#�=Գs��1}���BtԳ#�;�zL����Wl��]d4n���u��v�fG4Y�]���4�V�7X�-�nѾj�i���Ǹ��o"�6��^*3&L���Q�sRm��m=�H�xfDY2�d�*%��D6�Չ;�E�u-�:�\z����xڶ���A���U똜z�����2�Z��cx���ّ����A$M�9c[�4�Bo��h=�*�-��E��Ew[1i3�ث�9Wt^)R3n�ɂ`B�ط+R�^#�ݺ��;�׻V-d�� 亥�0��Fm����&l���+2:�(f���LRzѭ_��b����K-��E���V�<Y)d�^M67f�5���B����:�f�*��"i:^!GT���'�h���F<��^�&������:�,-m���������x�+���`@ԗG7F�e�ԗ��t����e�:,hZ���\�+��{��}���$��+i�V��h�d!��b��D��S;��y���e��w%4*��pf�D�6�?����;��aw��r`�Nn��&t�"�
���3mV	��n��Vi:*"1�;��Kf�b�F�Y�wl��j��Y�aK69�9��0qD^[���:��wuMc��.�p���G*��i���4���\��[5�z���`��q��ǀ�&7.��� ���i�h�4�GS�n�[�)�� h32�cP��;3s%��D���B��q�4�e�V��`4*���m
kKȡt#i�q��J��;ZE��ɯc�yb v�hʓpm�r�жaÄMǓ71�TX1�:b�U#M�����@M�ŉݵ�#����%A`��h�֑�̩��Hf�u�֡k$�nЍA���E?1��c�,Ôu[R�F�5��D���� d�.�#������wFB�M��hțR�U%��lv�m�*:��k�+չY��C�	{��ݽf�[�	�ET��:���7p�\@�F0ml"É�u*JYb��(!A��mb;L+j�aY�U%�Z�Xr`��5�TG{`�յOبīRv�%L�ˀ<y��J9M�P�$��vX�ҭ\I�׊�m?��{;RB�1���Ռ&;�w������f���IA��2���
��΍�[Z���f��:�6���fe*ZnL:n��H�-���a+uU���)��̠�-�Ѕ-ԶR��wW-�W7��3hѧ7P����`�]P�ڀ���1�I⬖q�f$R�+rIP�8�6s+-9?[r�,V%��lq��md�p��(�ņ�u� Y���A��_ݨ�V�eU���qh���JA[�����v�!M�� ��f�'Y�R�-����=���W[�IKj�����p�VI�e�M�v�ZON^�+$���x�S+f40�ű�i�-��K��$r�j����ԕe* �O7�u1�)օ�o���~�t�	��c���2l�*h�L�a��t-y7<3V͖-M��5��X��*@��^f�MS���
���ҭ���In�
�Y�^Y���"��Tsh�̬��ւaí M�&&��wI�En�;mm�t0��JR9,Bøf����	њ�qf#��q4�l��bR!��N�x���,�KC�""�����:;#�LYJa���m�¯Pd�����2S�tib}�ZnR�(��fFV�ͻF�����V9�.�mD;��w3�̳U�j�1���"0-m�o/�D��D�6d��Oikz]Zd:ҝ�cQ���Vm3�q�Jq���˨�
�z�Q��q*ڻx4��r�̡�#��L tJ�j���ɩ&P�0C��m�Kt3m�/.����LnR�
e�ɂ�3�/3�-y��II��j� M�2@ov����ő��ֲ/C��2j�.�ܺʙ6���"�7^:�����CF�ӰÕ�nClV퉹G(4)�n�X	�{��>8WޗY�K=��4�������%REfr�F�v2v�G�V�J�v�7m�,5�q�Un�2��f붡Ò�;�;F�[xcW��	zdZ1c�46(^$�&�mH�S�5o��[���̛d`W�m-���:I���ܨ�J6�]'fjdx� �P2�*њ�%��֑�H%�r-��lcd��d�ֶ���MF2�n��̭9VNRtkxS�r;%��Vc#�yc@	�:T�����s&�ú�X�o�;��M���$�BM�B���u�b(�or�2�9;�˵%���섨�+��u�f�Ph���1&�:����"��"���!;(kd66��{y�L(�r���[6�]o�b��m=tM���U �V���Ń4�%�N`KH�ZQ:�VBN�tB�R��f�ؤ+4G{+e]M� L��dՕ � A(�Iza����3	t�a-!Hlm!d�ŗy�V5��7j�{��4���A��+;-Qo2��]�]û�;˖0�Ѱ�:�^��J��Z��Hx+(v�Ti;fʋ2��Owb���
�A�Z�D
ĺz��°,�/u�rŊ�E�KE�A�_wT��fn*Y��n�z��Q�ئ�m��f�fG��R՘N�T�G�̲O6�3<���֍d)[J`6����yI�9.���,�/�J㩳q����A�̡R�Z�;�tJ�H�F�p�����h�*�,nޝ4-m����/q���؈�1_��[{{e=[�j:06��^Ѹ4%m��7��)�c��9Aa[�u��t�R�'&�K����޶&�ۻl�W}���j����6��6w_[��zFb-a��p,�`f�lƶ٬��V�M��Z� 4��JY0հ�±�^�����:D��.��X��d�N�ɣ�-����o�{�X�Z�I^�� ���8e�XstJ��;���m��<�GGv��+;j��;_�ŀ���^Z�Y��e4�K-�t��*��ˎ,�w�O�{uLֲ5�
	�4�Է��Hz�fm�f�hܒ;˱-޸4حf:��y0�m	"��!�X��|3F94-B�K���)S����r�aT��Ke�]���Y�Vө5
6^d֜�7��Cu�Jv]\�J�Q�Ȧ �/)ӏ'�O�H�@�%7Q��P�+pm֌ƞ�T��
��0@N�T�f�mʀ���y��S��se�n��I��ͻ�@�Zk3cyz/��mt~�Y��1E�wܑ���CK�&��W�	�͖k-��k,��,�FЃÆJ�-�ׂ�O�2�;`U���q�ӮcU^X�.Y��I6�C*<{7���c`t
ה��76G[BAvlQ�7V�b�M,�g�1M�U���#�3c�t��f,�Ox�[O�n;&���[�J����]�b��'H��mn�Cr��m��hQj�.�3V�yX֘]C����OXS*�-7d�ڸ�MX2xYk�ػܭ�f�mK�6��7 �6���P���ش��e�Ҹ8Jyf{�QD�Zf��3Ia��v��2cg��f��a�ї�Z"�Њ�{��,GW�PP	��јP�#F�f����*șvP4KAR;t*��0Ԙ�ة��e��N�Qۣ7k�Ȳ�˩acq���!*�i/�Y2�t�DfR���C%���b���{AG<.�mۨ/\��9�J�en�2�y�@J���j�
މn��|��6-�8A�B�'F�3����b�g^v6S�ۄ�$�x�suع�=ai�����6��6lP�m��ͦ�b"�E�d�7��#m7̭��`\���tNbѹ����i��AqebǺ�

�(�J�g�2JH�7��J�[�`�"���K^�#"
�]�V���Wnj�
�m�f8!�vR#���oz��0B4t��7N"�a��35�)��RI-��b�	Kd�����-�ҤCB���͋�c��n^'����ɨ�!X2���#-*������V�n�W��y)[�`dұ��!�9/ ��M�-��jU�6�T�*(-7��oQC������p�x�EfT��e-kwl�׬*u��d�_�+�Ǣ�T��*w�V6��(me��n]M��{Am��Z&�&y�v��t-���Xؚ�1�I�
���yo=��Tb����o��fms�Y��7j���jbm*�;yR�j̚rCD(a���|�F�]�F��+�cu�[�d;9BHYc^f$��(n�O!����b�vh�ܨBݖ����5I�ݱB���mj�2�b��.��It���n���8i�!͛k+)V�a���j���� ���p���A��H�n�+#��aL��cZ"��&����]S�'�2�#X3`650�U����ҽnLžn�p��`�"� k��k��)�3�V��(�m�a�Dl�+L� wP�i�n�Wԩ�n�c�2�rbp�eKU�2ޜٴ��4�=����IU��ݻŻ��oFT[R�{h��:�h�KtbY�sL6�:BT���C�5�oىㅁ����V�d�n�eX[�jښI��;9 ��r�Ȋ3*�_:}t����w�0�S�KH��f���%<ʍ��R�Ck0�M[�BR�aB��{�m�I�GUZز7{.(�z�Ke�Y1N#,�p��6��(�ܡ�[r٦�iɯZ�uM��5�,L�b�`V�QF�B���r����:�-Lon6�q�o&K̺h�㛔[,��CV�u*f1)l����@��M�=BXù�5�c�X&ҫ�ku�b�rtB$�z.�ӐMx���M!q�Ļ��d���FR�;Z������$G�^Ie s)N����n� <9��D9umd�Y,�'��4=Z�Sc8��r��cѵ3D�ٴ6����tҵ�6�=� Q��x� �*�^���0k՗����ӹ��X���g:�(1�r���";�A.Ax�42-$÷�*+�9�N*�2����ҭ��0��nи7��[N\m#Z�wf+D&���{M�ڧB�[֤��{���4�,:��u�f��/t����ڻgr5��eR�zuV�[�3۪4NlK8�E�R�G`Ti���E�"	cw硽����7j���W%��RZV�l��HrD+��hz�/`]=Wa0��5�)���>hP�ʈUo)ks�����G5�2���5gT�`�Q�d
�{vSUmP-J��xj��F���n��Řƅ;`�uo�R���0�.�j��O&�N�:�V�^�dKR
���%Ðt���+Y�m�9+h��a�J�`7�a�CR �j  �JXɺv[�N6��6ۢ/+��4�27L*����ڎ��+e0��%+�eT;���	�&�����rC�vܴ 4�]�n�T�0ﰧ&@���k���lb�5aj�Cs`��v�ѺZ	�����5*Xo�i�أƤ�1���*�̕z�$*9Ĵm����x1֊L�;%4pV�4�i[��P�3MvG����Jt�ZX�v�.�&<�H��l�j�#����{��r=XNE�y�d9w�b�e]��w[�
.[L!@h$\Х����E7{��/v���[��R�I��UGD*g"3oQ.�OL�u-���%���&KY���Ŵ�0--�Y�^�ƺ[�ݫz�*�AV��XNc�葃� y���۬��z̲Xw�j��qEh8w$ge�`�F9�@�cn��lǸm��=���.VScKEE�7{0<�X)�X�ሦ�5gi�ѱ�lf�o׻Z�)�u���qF P�t��[M:sR���n؛�q\3��wB���3*�d75��T���֮�6�:ۭ)��i	�r�f��-*�gS��"Lc)�4�492�y�u��g2���3.��1n�N<U�9M(�7gs1<r��U�:lj�T�ܛ{�^[�=xp���t=�G̒�἗{����r�9�\�3޴LR��S>ԛ]Q^^d3&��!���tRK;C)�i�^B����.����p���r]g�nP9z
�h���r���Z�9v����=��M�N�akώ:�x��/�W98���[ݭJR��u��ɚ2r�=���n0�5�wd7�eK����h!Mԛ�M)��	Y��N�j���
��M����&�v�άx��|�3e��X�(f�a�Ou�uv�]j-�Se��b�����`̛n�Q"m�Ӝ��c͑镺K&���:٭�Ѷ�i{��٢�������^��� ����C�/������mۿ늓Ut��肄
ڻ�wg��Y*n�U�NBX�'Cw)IƷU�qqB,����U��w9��S2.���EF
�e^��'GWj�#�U�Εֶ\a7�6AÒ6�T�b�FY2�,y��T���Σ�&��p��Zz��uu��Tp�|�Q����̑d���M� "�>(pt�r��$�5Y����y�QKh�r���$�\��s�ޛ'��������F�jt4�^��#�|]��X<]7۩≫���W��c5����w8R=���ʂXռ�	6�lƜ�wX�,)s��Ƿ|�맠�����z#�Չ#b�s/�u]k���m���8m-�P�tp(��M/��5Ȍ�E�(>���B�-�`K��6:�M��$Mut�%j��B��u����D��m�)a�ŷI�,0�6� q��/���C%�gt�ݭX�����9�T�Sy�}���Z�\�cF��st�~R@@��	u�����	(���<\f��\γ�\�ӵX���h������wֺfTX���a\��5�B����v[H�Ņ�ul�5Z�C�.uY)-�=f��ua�y56�y��dG�gm�[B椛W ��mun�{%�8���{�)PԖ�7��=��k�,��4Gt2�r�T|qmX(�q+ ��b/Cm�6���тw�uo�
!à��𾉌��m��D��`�Y�V�鼦��u:���*�QU�w7���2��Ӧdˆ[�1�Cu�P;}�ŭen8Ņ�\8��`�7�֞�Qfr�S����V�X
���ur"N��𥛈�4#N�P��4�+�����:�s2��&�KI&��L
y&�ָ�WgC�{Kݸ��F>�]�v޳2������c�ms,η�������:89�i̫�F��#R(�G¸�wd�;��W�9����5R^ΰ�4�cx�J�;��h���������u S����]����"bA`�ίq�[���7:^:�1@�a묮w�J�voB� ������q]�m���uW	�����3�G��*9I�ڪ\�ɁG��zz��J�ľ�[\�W%p����+|v���"�-�ёuhYW��9��j�%8��;�Y�3Q�Ǡ��i��W.�W+F�N�8�P��H����6[���
[ۍ�0�IXZx�%_:�.n��(�oc����.e,���<�������}�.;�����ܨ��ɚ�-b;� �!��+W)xv�t�q�3lh���HҐ��`
ņ�I��yN���-Ǵ�(�Z;{Bst�n��nU�t%[��z�d�Ž���N3ݮ���� �+�[Q��Aܺ��Y8=�Z� ��݃-����ejEOk٬�t'n"�ڌ��{����!�	���.�u]�X��U��r�`���ޢ����{G��x_���n�u<�]@��q����H_52p��ܐ���(j�yc�#����
/ë^���*L�Lw�l��
	%�U���I%a��]�;ӿv�3���ƚ�U8*�vVv�ǩ�	X\%�},3�Gk0G0>ݷ,��ų��a��)�l]a��P-�Q7���pVDw�em�鲧��BP�qR���>ɇv�MVg�z��[����S���@��.����N�ܭ�G_<ڇr��4n���.��3����\��.�e��uj
��]*�FA��!z��V�-�v.^�۔lJX�wU�b2�kN:P��D�e���:^����R�Cn�c}(m;���ÿ����gb�颺+#%�_�WP�r�^E.�ֳM�J5��e���yf)E]k����,���V�&Sf\�S��U�:[�?N�yۂd�3�����7�:$O��ns�.es�����řʡ���5l��6��iW��ͳ��7��k!��+�J֧+"o��#G��J�.��SPһi��U���y��c���q�r��t`�ͭjɳwu]&��w�k�\���2Y�	}�n+Y��!ە�MD��,�;y����x�pWSWpk��1;*S0�Uڞm0&^u�Ǯ���{����Z�*T�J�2��Ιt�2�.�sr�]�G��rfk]c�^��c�;��\d�[ڕ�fՙ��J{���'���^������rQܻ�z�
�S���]��M�x(��m'��vd������B���B�̉o!��]rG7\U�Mչ�-���dUmA86�D�q��9Cja�o4�����f��`)�2�ܤj�)��2Q��A�(�gQ`J�7�#8L����y(l~�Wu�J�aұ��b6���HO	��p�8��,6��Kn%@Mw1��w�tV�-v�;�WL�K��g5�r�Es5;���Vv�'e�0+Kbq�d���J���sfm�oc�i�$���3P�)�&�ДK�9����GY]Nֹ���s��-9-�u's[ջ5寈�Z���
�r��l�4*��+4����|h>��hͤ�ն�ck^��y}k+Wڷ9��x��_`��븨c�9ņ4��Wck��Ϛ��էl��m�ݎr
)Rܴ]�/�z��/��m9ǛWF�����v�������*̓��}a�sX�L�%��Y[�X�sMF��i�n�	Hnm�Ɨtz�*f�����Wc۾��I�V;|7iᣙk踒�*3S��RyW��}AD#:�I��q�:@Z2bR�dK�VT�`�Sk�b	����'.G��[�4,���ϭWy�|��۹�6�%@b\���Xf��j7Xs:�n��G�P���W{�Dݥ�"악Pɛؒ&�&vv�%c�W;��B�גZ5��Z{u ���3)�X��7�z{�D� ���o"��ܢ��W۴j1��%^�<Be^+��+h����k99������k�G֭�U��ڷ���ƕ7��"u��;%�x��W���=�`���]��{3�js.F�|n�˚�"�BV��P����$�)	���K�k�7��X{H����2R��m_�;�o(�%��n?i ���4�J���3Y�,SC�XT��c.U�B̂���38bX�_frmZ�
�)&՜��x�FԎ'��yQE�H+h�9S�q�P��˲�V��`��R��j����R��Q@���MhΔٲ���0j��*6A�+R�oT�,o
�lRJF�i�z��H����ɕ�.����ұ���G��CPV#R�{V�2�Q��Q�[�k`�g[���x]�j:�2_]�����oo��<{��U}�PL��[(�ܜ��J��8q��,
��j=��4=%[��j��`V%�/�p�Q铧-�Da���n��9qv#�ֱ�ú�����R����j��q]���ث$s8��N��Vұ�Q�L3�fk���� ��t�MU��j�����;(�Էɒ�Ԯ�*�p��;�������:��X ��(��B���"���=J�<U s�L�5�f�8����c냫�z���0KW&9��8ll��h���n��ϙ�.��*�e'tՕ|�2���@�9q�
�R��Ψ^Q[���^&�.�Ӭ<��:�C�܇��cK]�8rG�v��$�KS2�E�{4{{F�.dƫ�<p���ڞ���==�ϩ���<�o��5��(�֩�q��Q/cI7�^Y��9h�
�`q����I�v������F�k�,��RۘYv��vԻ��;?=�.؊b�q�La=�y������gz��o"�z��P�iΤh
�d�e�t�&w�}tѮܛ�v�̬\�"^�:r��w�
v����e���\����-���\��e\|�K�me�E!�%xͰ����V��Y����4��h�M�77���ż�,�%gҽ��۽�9"Ӡ7��6YA�����n��nv�N^�^�}�i*631ޣw&�5껱¦8��:�[՛.0N�J���9�I�C|�����]�	��v`���T�Ji�AqL�U1�����^R�hQ�'����Mܶ�ĸ�����	���oeݵ�L'&R�[{�*��뛑�d�2��@z����sQN�͊��+��:�G���0��7�gzķ,����;(l5a�'9�����D��J�Vt�(=C��q>&���u0oL�������p�Jښ<�XlY���ŜBj��&b��X�qP	R�Y�e(5I�ݼV�={xP�n����;Cc���`S�F2u@#Q�{z���P�u-�7V��Y��.�sVΝlm�c�)I`�sjE�[k`u2��	�2ߵ.�uΦ�w!*3�j`W�[�O�&~;�<��|�5���Ú�BU�$�]z�<d˘p���_R=yVܵ�����02�o
��E�8pT���d=ڪhţj��z�8��|�k�Nd3Ka!S���i�˰ծ��i��4;z4_\�.���s�f�/�+�ٜ�;.�6e�5p�١l��J�
�tݫ*��y���Z�Î7�o
u�K����[�9)���Y��z켮3J��m�MT���;{x�:�wj[+�ɮ��l�ԭ�,y4��{sr�u�VE�y��<��Sg̂�u�빇O*-�J���[#�h�{zD�W��Q����E�m�Λ�6�dzN�խ7
T��#쥎붆]��B�O4���Y�h$Z� �F^���U��{R�ޠ�Wz̐�3L��F�G�V��U)J�/��5D�e����w���s%*u��A�T^��aQ֝�8>�k�Dj�$�욄�����������A�l��g�j�<�#�f�);�ᆂ�+������}6G�\;ϵԣ\�0ZNn΋ W�NsY�r�X�ZS���J*�ृ��~)$�-Z��%$U.r��9�X�/�(���J��G)�"E��E�*>�j+��tVS���D^���`p�: I�@K�Q��n�9��B.:RR��\ح�i�:f�of�bǹ������!�)EO�-�2}���:,�L��c��3�Т̛,Fk�r$h��ɠ^g QGP;���(���w���c&E.t�c��=j����8�X�I.�db�'1��('!�'�	uv�!�[x6p�0�Qfov�x�X��Sچ�[��Z+�Q��.�s.V;Z%��@jATW��'%{�R������`�t���W��Jk~O2V��^w��Cїj�MI�tqn`�E���Kk*N9����	۹bLy�}7uޮ8;����)B��tE�K�E[[�#�{�IN:����f�)95�=�
3Rl��;v��o �Y�s��B������5)L�}�O<��cĿh�Ơ�8h3���^�pUy2wifJȠ5�Bu�W*��#���6�kk!��c��̰�2��f��6QћX�ض�Su(m
�+*�L!S�f,J�e�Z]M��j�JK�w�7t��͍m��)�=b�r�=׹b��bS��39��Es;u�*���+�c뺡����v�ᨙ
�qޤm�Ky�E�|{/��z�"x�~�x\s�_ݾT���%S��0�+S\�k�+*T7�v:��ORG����A,Z�1�;��y����
{R��I�P�tz��u����9��$T�,�2�g�*83�.�<n3HD5�򺤜�ܫ����C)�kӍ�]n$ť:}w7�d|��+ش���A��c�s+a�K��ø�̮�hv�vhV�e$È�ܴ}x�5����G��U�\�dt�u��C�b�y�c$����K��+��%�5��j�\D�xTL��h5>Œ��x�(at�1:FB�Pf'/���+/7���!`L�T�s��Lrk�b2�m� sY�z�Y'P�k�A�63%X��K�l��$����} ZI���^+�V��j='�Å%�'r޽��qVa�c�ޏUl�$�L�v����w*�����V�,$\�0��Y@Nh�]����;̬V�fs��\x򚬜�MYc�\���c����&��5^�XP9�:UҔt\(���V��ӽv�|�����b�����S���V���m��rE2��[�s`]@�E�
�Q�ͭ���ތ��Lv�2V�G9\o�0Kw#*�t��7�r�����vK4�i�{y��w�Q0���.��W��9~W;�lԁ���U��u�J�.�L��q�b5{5�K��2���۸Z�v��T�ё;�"��ʛ���a�oJg��xt[�}���4��?J�V泆�v�M��&�\�y�䤮�+.��+;��bV*4���ŧ*b�GU{]]�_2��R�VƩ%'�B1�����AJ�U��p�>�2�z^���p��iL4.�C"�[u�c��K&���G[��Ǝ�o��avE��*��#����5����bü�S2�,��^WR� ��]Օݽ���r+
�Nd���G��՝tL���&�������}��3R�������An��ue��ƯAKu�B�-0�n�x �;/h9��r<���0�ag�<u���ݿ��tJj��F�-C0n�\�7d�i�,�/�is��7�t�ǝ�30E� fd�5�$�+�7}����/��@��֠��Sz�f�g�����=w+�o9��++V���� �a%���P�GL5��� ��kl�M��N�`�L�v���9v���P�rJ���5C��n趎�G��%]n�sr�C���ǵ�{K��B��E
6ep��v�NԲi��54���J{�{r	q�%��jÛ�e�e^��,�h6���Mf1��Ȇ�-��L�ٛ[
;���4�Q�-*t�!���i�@C���	P���7
 (" "A"��2�b	~	Tn��R��h�V;
@�wwTUD�^� �)��Զ
���ܺ2�Y��H�6�,�̫���Mq�$N�E"� QA���F
�k�����AH*���P���j�υ�t	Q&�j�l��σ|�|;�uz��������� � ��������􈨢���o��������������@_�����?�C� ��c�.�&V���x��C"f)z�m ���c/��jMw�<��^&��8`m���1�FrU��.O������7�`�����՗�Ԧ�n)}_����FC�oD��4O�F9�1a��j��y��n�8z�i��x���G���f��[ �¼��A�n���۳Si�8�� ; S��T�X׌���"�8���Zs��Ū�f��-T79Sځ��M։j�ݰ�( �W_m��_JT������Y�l�p���r��5�!,ZW;Ժ
|;3��I�<���JnH��Oj�<�������-y��.���Q�.�U/]ԳtaF���3^�����9�C6s�j�jA�'*�ݛF��:9���*c	dI�γ���
��_b�K^���[\��|�T�cɎ\fu�&l����P�͈&ȥߑ��� ](:=u�fq�t̢���$�tn1�N����`�0�n,-���9�L9C�Ukj��x�p���%���;�))Q��&*Kק��܂I=�z�5����Q��/�ޝ]x�R���B���wn_,P�#��n�="Pb�� B��-B̧�Y3j�K�z%:�Df���IP��{n֙�)glOzL,�gv�YX���f�q\�zxnƙ�,���A,Y�v؝(;S���������[�.X�3fi��� ��VCk�O3'[�VW=�
ΰ�ȹX��2��㠊�/tᴥH��I:�&�Q5�q��Ն�r�a�;��F�uD����n��P[m�z>���ك:d�a�Ľ9a]u �8])�Վ�c�K5�-
o���.ޤ(����)Ӷ����M�۵t��sj��.����$�m�c���"��h��vdlݫ��J(�r��������:�_^�����-����
��Z��n�T�@Q��Y�ꉘ�댺����M�x��c.�Q�\0�[{(���2���ۑ�W.�l2����nSU�3���Ե�<ڣo������8(Ɔ<ܫ�i��t��·���=)�B^p�G�g�7��ܘĵM��j�Y��y��88[T�s]�l��u����v��q�1G�'/GK�E�n�;����g�]��*�C�ы\�D�%��T��&k5�
7
t��aV�m�}���gy���J�h��L��Oc��wc�V	��ԯ�مkM����X�7�<����U�z�݋r���^[U�@*�mK�*�_��[������O�����y�}�xƔ��\l���P<h�!ndk'CY6<��\��noЍ����E�Y�w@h�L��`Wnh�tWj����vⴝ�����F��S���ʀ�*k{c[]�$R��u�6Η��������q-T���Y���,ѷt׌/4t��^QI�^����u�r���ʋ�/�g�83�'0���R�:��|u�etә�"�X�F��D����ՠZO+��C��r���z�m�����7��k5�*�f�2�7څr�c����2�m�̮�����"1rk.�7��b�tu���5�i�7�p���)����e:�:|��[R�ҵA4ৼ�u\O1N�M�u��p�5��֎a���Z�u"x+����R3S�E>�Kdt{��[��Vꦕf녝���aӔ-��J���(zb�B�oEm�nH�����7fs&���*���/9��t^�ΕjfZw���1�N�������փ��jm��a�\(֥�3�;[P��y5D���v�gir�]8V`��[-ζ/�.��&)�'�*�9HW������ō��u��3;�;I�w�w$(h1��[��9�f:ai
v�s��=+h1�Yt��/��vܳ��<�j'0\w�oS�LrY�C��h4��gQo+�EBU8�̷|�u^��u���݊Y0��N�GO-V|���ȳ
y)����ɼܶ�=w0SuUe��P�I�u�z�����#SQ��2�t�Fn�n"#aD��2��ؙVݷ�mKY8��oJt�C3�wP�1�C����R���,��⣏d쨳����������02��r�Ѷ��Af+��+�,�uw�=�YJk�D���Z���y]2��[�g=rM;�t��1����L5�WrfҤ0e�#p�Q�5�t�vl��9}�>4�.��x��Ӈ��i)����YUM󮳲j�5�Z!m�{��/�8�}�͗]��Z-���E�B2vL��-�o`b�Q�q�3��I}�h��Lѕ�&��f	��˨.{MVT�f���ÙQcJ���g`!P���=3j;:;)'����w:�N
+igT��a�I�T�|U�\�Se���k5X.��S��cNabp�}]�o �y� ���v��,�bT%�a��I_�!�F$�^�!����;צ���NF�.J�W7�:�f��+ ��u���.��M���ϜUG�����M���P���,�Ve���V���aqpy�.���ں���5U��fO�[y�f*`��r)�&4���f�=H\�j�@)�/pF��y��^��/���&���V���S|����������-��5n�N*��G���[oJWCu�+��n�f�h��d�O%��7��{&3W�mzt���U�:���M��l��ja�t9	�� N�Ý]n���jF�窈��LUu�䩅]�h�[�S(��Ƶu���yІ�'R��vX�-[���w�\H�W	/�Rs�(ҭ�ķ���;�|���qZ�T��WL٘��U�m�x�+G-O�D��mNU�,��o_gʵ����@�N	5�a�f8��z�9y��c��ɍ��(�g�TS=H�+���Zih=����-|��(r�C��f���7͓N)�-�	�bãT�];{�����s�ZӢ��}�)��6�+V	?v���3I��0dm�8ThU�.�.����*��W-�>����{��$vu;�KJ�i���Γ��Q+��L��eЧ3�be�]'J<{kE"�R`�R�� �2I>����k2��m钍�zK��%
j�xI�!�B�x�Z�J���U����6�Z��ۣ�DZ2�\�x�v]�쏨�F��2�L��������ٛƝ�N�$���kCf%pW$�6��B��h�M���ηB:�5�|6Jg��D�ihȖM��8�4S�z!�ڕ���jS�����k��yt��߭�olX�ʮV� �<�{�o�M�ս1mX�9_��V�2���2��m=я�[�ʗjV���:����	��)y��;4��e��!�e�t�.�H9�ʔ�Fb�o��1�@��;y=�r�U���j!�*6�fX�+�du�ibþ�)>�;XG�� ��s�u�&qz�Y1͛ᙂ��Mn������ͷ+��w!0��pkS���^��St�C�+j�J�QI�vv�!D��o^V��no֨��/�4軈�ŇcF"�JA���D�9��8%۳�r�(K�$����������҃[�;�ͩ����N��W�{��F�[݁��E�uE����|��#�2j��J��w�����|��VYBS*�ϣ<�3z^h�0ø�.�tk�cÌ�҉�̞cu�F�wj弈V�+���Yɝ�t��ie�a�j$�/�tyZ繑.Oz/���h��J_<k��ծ����b�N<�_�f���W�8䠷L!�����%���v�t�Z�Z`e�(^���:KT�=���c���}#TM���C1�t���ص��qfS2�=N�D�V��5��U�61T}cinq�e�F&�Ip�U�[&���DڦU𼶦�f��yF�f�6�S�=8eI�yX)o]ؒ�ج�w+y�M�j(�7�����B'I���3Ya��|�Bы���7cu�+��{d|�m�~���wm>0]M�t�Q��&F��5�iQ!��M;����T�P�~ځ���%�
k��hu)��E�Zwe*dT(#��/^��T:��E`��l�ٝ���M��kǤykA�8˔z]���-�=l`��wއ��<g:"��;s�M�>/3@9�?�qTN�9��e��S�䲡a�h��NRtlh��t�G�e#��m��ɋ������.��j�Y�++�@�ַz9����ە��b[����aY`�f�7��FT�=v8���vܭ݀��yW��#w����h��iJ[�`�6SY�EZ�DG��rYՊE{x�(�;����(��9z:7nJ��c|t����1��%U�6+2&��G�\,=@���2`�d0���3qTTҰ��{���<��6Z'�܏�����k:<�j���V:�䍌-R�|��ɑ�D��B���I��wô!Ϧ�dd+*h���^7+�m��+`(�7��6:b�Vji���T�Ѣ�I�ol�T�NiaZRֲdw�ܷb�L#M[���ŧxAAwh�.!�ah� @�iՊ�+��]���ɮ����5Ğ���`��L�o�n�xv���-��K����'fJsz]������������++#F�AI�#h�tJ8Z��Sv�3kY�!�n3%Is�-k��U9�i�$�6ڷֻj�T�!��t#-�t�O��\ ���)�m��ӵ,X�i�O�`�|,������J��c�޹,w(�6d�E�o���mm�y��J�p>�"��R��,�Å�`K�k$�Y���5� |ct�:�K���2��L[�su�@�K=R `�s8�n+F�
\�0CS*ԇ���o�F�$���)��A��啨�S1�]Xæ�=W]�ES;*u>�@Qt{):��B��V�!�tӤ�Z=٤�in��r������L7��;:���q���skTľ�)��n��Y3�0Vuv;�A��^	|��{��#)�=N ���o��Tڜ`�z���|�T���b�����CܨK�j�<fU��MIE�wY��k��<�h�|�[Yٓs*�%
BK�4X?cQ���;b�-Mj�'hɽ3��WZ()����gIy������ph���R�X�oi�9�e�nA���θ���%G����&t�[ˎ�Wn<ٱ嚷I�"d�@���æ����)�Q���Yȭ��Ƣ��1�of���;_z8�ν�����������'d�3k/e����/�}�9�#��*�2�K����T)�]=��h�ﴉ2�M��G;u���%3�R��E��*t�I���U�qVV�u)P����V�]��� ZɎ��-q�R7ӕ(�tR��������)�-�s�[���JЉܫ� �.���)\�kk��J�4����l���oXZ��F2�F�fA\�Y�����7Ze�^��5�H�H�|
�n��+Cwy��vT�T�K1�[S^I��L�%Ef�g3��A;����q9���3&J��w�Ŏ�@Z�_J1�>�˒\[.��F%��sts�Xvo5�W�T�E�V'qӟ��6U��f�"hڡG���ZX����3l��-��I��&�*�z�ԥQs(�NjZ�Ô5��r���B*ȃN�ۧ/$=;�����r�����G��J���{�i2�j����㋱ȩ����-^\uJU��ۮ��)E 8�٢�f��rw����v�>͚�ݴ����"7Bj�f�
`���S���#u�oT��$8�����9(qY�܍�.��^�[
{.��]����ۿ�#�NVt����c��0C����0u;i�[�>�X��&E�-i�	�%Ӏ�5����9YKM3�F�G&�\1��{�;j���E֌n�,��-�,��\��#��.:��Hl�6�LW$�^Q 4�U�BJ�T�fÝ׷��VF�������ʗj�hU�g1ѻ��Ic��J�0�-�o+����H���$cְ����&�v�S�DT(loD�7�w�x�>uݖ�[LE�rS�2`ŕ��'[K]���
ښƑ�� T��4g,��יUy�i�씰]�h�c�A�,o03iu����Ek�b��h]emkv����+�vL�Շ��&ok%nl�$o�l�B�
U�*W�Q�z�\����m�\6���b��ojR��,,\}C��2�z%,��t��u׻�C�@q��m�ɋ̊����S�w�NL�[���j�:��J������콩��9�{���FS�]Jm��R&`�v�%ݑ�Un8{5=u�h]�S{5ǻp�.�N�2�F�(q�4.�Iƻ���x�l��t�WRe�$�sr������hIF�1d�A]|}��a�ŮŔQq8dҨ�6/T�īi��nR�q�d7ƘI
����}(e�r.�pZ��X��LG�e���l|��*��ERn��d��R�E:E>x����M$Z�	J�&^��0���m(J�O��E��;;���^���OtUՅ	�	c�N���:��.������
��,��sO(��e9f��p���-��̼��͌>{�X�qҡXQN�Er�˝F�Qu�!y��+��$]�܃�S\�������\M@REVk��i��o>z����'����?k+���w�T�byg�������;"&�UY�(�sh'���p�=8wt��YoVYu�57[.�������Hr�tU^��'�u�R�4�E�ɵ{-�4��f���x&���ҍҤ�K�̥�<8����f��s�O���\廃��`���s�5�#��K��b�W�3(��3��A��y���*u^L��L|�Tv�Z�Cm*tŉ��h\;D�r�z&�Y�9w2��<v'�rżC"��=��� ��Ww��比��l���uenoZ�8nq������GazI˧��X�����������< ���:�������O��_��O�'�s�������|||x����������B�<I��7�rN��M(6i�K�?���H�㷉g���=h��+7����dK�J��/�o��J0-�=��J���F�k�ηZ��z����G]#��/Yй�\6elKP�(`�F�;��;f�%�WSoSU�;^��odkfY�}1T�q��,����-L<d,T���f�w�`.��Y"��K$�DVv�b h�͡��{�Z������n��6�%��J�VV<���v��-[�H��o�b.\�08�u�V���R�h<��[mǇ�NfKðā\�������c��r�5�q*I�G�̾L��uo�Xh&�Ij89��L9����ݨI��/�ʖ��L�j]�HV1���Uږ�x�l�C6�J7YnT�(Sַ̀YF��
�� e����hV�GVv4�;h�xy�oer���h��I�a5�^C9����8��.>R��޹Xk�����o#ʘ(�$�Q��1���ڣ��[�P��T��]�L�Ύ�b�v�ܔ��)w׵��T�ڹ�m���s�;��w����<Z�1��b�Do.�{� t�Mk�(�$�]�kV�;��vc����M�:�\��2Ԛp�Q��vU���tph����r�UM��\�儞�*V��wK���f\��b�4m�,�j�^�r�K�g�֯7.���8L3�,�-��4���D��A�˩�V.&]�x
�<��H��Űѭ%�����(:6�c4L�E1T��l��7gN٤�I���ن����h���EQZ�X��s�iq�h�lb��֩�	�֓Zu;j����m��b���EA]=D5G�F���6<تh��c��'N�&n�&�OZ�kF�����f��4�;�����;��j����Ѷ�58*�F����Q��4�m���bAE63����T�EON5�lPPE�l8����53K�jb��"h��í=���%h��j)�b����y��bk͊(&h������RR�DAUkR��jhjb�q���w�$KAU]���Ϊ� ��i�MDT4TUv+&�tttltlcJ�:"()��'l��i�~����y�8�O����k�ٕ��oPvղ�趀t�c7�l�������×��o���q���J^���t�Z&p)� QӦ�
˲�0��G,�a7[�R����/�4۽���j���se�}���������i��u7���?��~��u��w�@WX�bԄ��{#/����}T>n��y�d\��W�W��c��K����
��+K��MzG+�d���Ww�xoUt�%�1'�_���I4�]�/���B����&c1���K�f[��3��}�Ω�[�+�=�2�[��5s�/7mOgN���$�xG��/�sב#�`z�>ɍo6��=��
3yE��q,Mq1C�񯇟���G��ӳ�E�x���*ؘ���;�ps�3q�o�	�t\Z�z_}{Nzz��S��ok���Χ��t5s���N=˪���~^'{���z�	�q�;���@D�>st0|����8��X4!��Mi�ܿl �z��V��7<�R���>��Iʽ셧�����7�Ϣ�s�9�/: ^f�tX���Jheo]Q�f���f�������u���cS�z���
�,iIөH �Í����u�00B�n��ם��Ҫ̗�k���L;ՠ{/
t��Z�'���|ua 9������|䵻�r����PpR����e��y�+��U��m�{:k���s�3��W���re�PW!�tWL��t��d��96�p_kx�������wO����O�(	��BP;��g-.�y�:��d��z�%�^��(��qQ��m{���K��v��{5j>;�,�F�a�s������us�.�g3y�A3��f���]zo�#$�x��Ӎ�,Z��Ȑ��e�p�̗�U/]�r�vJ�}k�(T߳so�~��%��̕�ْ��E����M_k�W¸v���:�2^v}:��4���}��u�f7G>��1�{Þ])�����8�S��yw/�d�#�����>��k�s�n�w��������s�~O�.o����'m?W�`5i=l����`a��Y����%�!<�lf���0�B��X/HNhN���܊p��g��`�b(�����t^	7�V��e ��z����TӮ��hEؗ�K���$l�|�p����%�V��4%�����*즂��"�'�e٬�
�P�&�qųku��Y�H��+
3.;bS7�����Yn��L(`��׻7�\[����_U�$�5� ���]�k���f(nv��5:
Y����,�m��z�XT޲{͞�?s1,�9l�	��m�Cx��z�ec��@��ܥ8
�N�����s�\�`�jv�n�F�M�E�Tnܪ>3�ϩp
ʣB;��3�鵘��FIkʼ�:��M��C6sl5rz��{����}+W?���B�.W���v�<�{~z	'��B�����g�j�������{}p٬COq�+��p�f�ߌ�w�NL��Q�ʌ��i��z�W[y2��/*XR��2���cs�u0����\�sӸi���A�T��k'�����Qw�/lC�mu�4��	�?c����nH��f����~����pY�~�o��3>-Ǖ)�u�%����x�UBs�S>�+��Ӯ�>��އ��v�=I�����MS�Y��-_I�ƸV[��*��ӕ���üg�9�Q�('ݚ�h�HX�ؚ��bj<�r�-.Yd���j��Z�u�Am�`�mT�����|��w���^獵��%EA7�X}\T{OF�Mu��5����Q�ׅe=����s]#$���V�{l��&kΌ��ft��\�)�C;v����A.u�9`o�&I&��컪�+l}�$�z��|D��Z�Ηp��`PڤF�=�Zx]���y�yg�������������W�d����s�e��"^�٘4�X�;e��d�OzM���o�3+C�.朿�r���V�k���~-s� �z����X�5��x<o�d歉�PE�K��sw���W�d�T��wne����>;`W��d_S@��8y�^;N�� ���+�s����:)�c'M���I�8���]��zE��>]]��-^W����-�<�9���/6o���jN1ߗ�<��
�I���	�~����}��'���]솻��t���1'��ߧ�ϗ�C�8�����8��z��]����2��+��L�U��v�S�{'�G��_]˪އv���Kj>���Ob@���2�sw�^�Ec!��H�76��p��2��/(������������e�	]i>�`s����9�w,*��\zH"�N�0��6H��	j�xgv�$F�y��mlퟶם�;���-�M�꼗������A�u7�*ZeҡWVr��-��E���YM���4��V�<��ogXU#2���;s���r��'���ק\�[^(S���q�	��
]N��9����p��~�����K�%Z�S�R��yP�UnY=x⪗ϊ������z���-s�N�Io1��xL�և3`0�s��m&�3��9����<�����q=~��m�H�{ԟ��W��[�UV�'�U�9�{��m���K&s�w�_'S��uߔ�V�n}��dާ�}��ۜ�Y���� ��⯲�9x������З<+��������wW�>_M�L�(�(1]{��������ES΁�)7��k<I^q��4�F�}��rC��{�qYd��/|���ݜ�İȬ<k$�܎5q"��d=�u5�;��Q����\�}wd�m���F����2sl���6�����T�wj�Y�=����Ԋɼ�-~{��۝�o�o����> �U�j�H1���{�Jx�u p\��d{K����p��i�[�Zs9�����W[�p�Ht��[|ٗ�WZ�SJ�A���W8��74�[M����ơ��ܒD�p=����{S#�4Yʔ-(�n�꿽��/f���'��2w߰��0[��y��ف/0+����]Rת�{���p_Ϥ�矠��}G��y�y�`<��ђ��yb�S���~�6D80�Ș2��=�Lf�g�ߗz�iѱ�
^: ϲN�HV��;�(��������ҷ���<���נӞp�RZRg77܇�{��M�ʟ9yb�������g���z��V���;�t��U��ɽ�}�L˙re	��R��?K�+�}u�֧v���֊2L���|o4���O���{K�ܐ�ѯ�aH͑0�L*'Z�J�q�z_e5��k�۶,��ƍ���"ʭu	�z��������=�l���u�Ϩ\'>�+��w�������V'�xg�9��z��=ݲn�03:�����������dȉ�j��&f��~$[l�����K���k�����zK��Ԋ�[ٱ�A��6�gr]zii4�s)S�ŵ�d;��sQ�ݻ�oNQpcs�;������+�ܷ���Ij��nJ�i1v���;<ȠlGa6����rƨ�hĦ�:�p���ڶ�Ilo[ޛ���[�����J����d`sb� 5F�N�ί���Wop��Y μ���u�ta&T�/8M���n��cv�ڮ��o�^��U�:��<�|7K�7C6x흓�b��n�\e���N?*�kh��T�gEu����1>�=�篌�ӆ�cF�/ݓf�(�wo���y4�A�
�=Gx_��\Vk6�=���_�cf�lcִ���r�����q�����?L��3�������!6�ó���(y{ե�m��w��)�z`��y�.���Gຢ�V[ʻ�_S���9�Ǿ(�r_a����`��Z���ץ�Cd����{nW�ʫ�鹍Rƻ�z׷<�7��5w���g���q����h'ǾL`�����V�K�3G: �6�F�lY�޳z8�^P���^�����9b��Z�;4�/�Q�u��P��b�!�=�[�]iM���O���U�OpP�tL�q�!֖2m����l�μ��x�O{v�/���gg�i�Z�r�ڷ5��#vN�8��=�Z̻�n���=��wSY�`Ul��*�=��N��s��0^��[d��4�s�+�z��L��t�5�.r}Bv���Kٕѝ��oVΕ���n�[b*^�֟��c p�3\H����>� �aq� (���/�XiU�ǹ;q�^;�Y�^DO}Y`ԯ�і��+d����4��to�'�')����+)<#�h�S����j��L�s4oI�4}���ɺ���>�vߘ�81��O��.}��\��9���e>q|�E,�k�h_^ҿ�#e�{��[�M9^&�\`9L�6G�uBO�f]�u�S��/�̊h{��5�n�����ᑵ!�����v�ͯy-ڪ^�<�6��X{T}!��^��h䊐N��g�쪞%�p3#���u��t�K`�=���Ono�3�C�L�,�C/��_�e���R��6�+�t"~�)8z�bz�ӻ��.�ضg���ö�Wmˢ`��][�Q|����Xs���o1K��^�(�גfK_>�O�o>G����&R�̸&�帜6��3��]��5�,i�Xai:#4�bE	��[�y�C�7d<�e%�1��z׽J��������h���`%Iº��X�ń5gj�Q�����'����O2I2Ns��$���������|�Ϟ_��7��^���۞�9��"���d��Q��i�e���u����7��K/�j)Py݋%r_RZz����]�&2��n7�\oNM�;�ެ/G�\�U=[+���~�X��\q�������{1z��Ck�ͥ��tKܴe;�N�F����w<��*rD=eߚ'-�;BR��5���]�.v}���^�pq�V7��w��L6�m���x�o!�Q����|��vj���6���eC�|�Pul.��2��t���0�m�^�g}���w��H�ER?|i�����Q���'c�w|3x�%��3��Co�^P�xnv���D�jp�ժ���eW�?id/��;�8}�6�]��3ݍæZ�O��LNȲg/x��A57@�`f�b���v6�q�g�Y�����+���6<�8���mXPE$r��������ux8?_Ǉ�������Z��
 #���s�cr*�ԈND��=�����+Z��Xs�4�{wj�K]k���u+����FT���tͶU��Ʉ�Q�u��%u,6���A�&���~-�Šg?��Mސr�Oײ	v�n��ۼ��ڈ$���nd%87lH�_C�'Q�o���z��_�r����_A7��I�ܢI�,	؝�j�G9���Ե�S_T�^+�M�Ntz)m�3ѝ�����ۮ+���L߾{N��8���Z�<��^��ܺB_0fĹ:~\)_�����|�zh�?h���y�����B�Lmp�km����#y����E�r���c�,�O?e|<�}F7��š;z-�q�N\��la�8N�.�v[߳a���z�v<4q�9�ϗ�����L��~NK�[vN��`~�lP���.8J��v���j����h�S�+Z$���d`�ӈ?}<2�<YN*|�XA?�3����|����n�Q�S�/t�V�P�\���e\��L�2��0�{F*�< ��������y�>�G������/w����q�<��f��ڳr{[nU��Z��FW��L����M'y7��<�K#�!�3-̙[��N���~�JwJW��qlw��V�h1�Q�'��sF3�̹;B.��}��"Lf��Ve^�'������,��VTz ��[\PV�ou$2V�)Y�F��Q�+�vR�VS���]���eL�4铟�w�������YQ�t��(���!x1�
����9S�ASx�s���H�H���v2�'z^*&ά�C{�Q�VU�ǭ_roc{��2�|�l�𻵛|:��Wyu7�t2����>����*<�]*Vn�)i�������I��h��u�*�j�u=u�E�O,3�k�}Hh	��Y�����
O@�]�Yu�=��㋑�Gƕ�3"	zs]m��ǲ��_\��0-��;L����!H.�oή�l�_�]�܊��a]�Ք�r,3�a�Y�'zq�mff�#\$(��P��F�:cy��\�=%���*.]���KUh�(v��ٹap�sc8"��|����L�6�eF��˂��r��P�[z����u����,O��q[dQ�A蕛t��t��Q��ֳz��<CK7���4���
��厶�\J�x����mD� ə\w���gn��`�(BfC��\���.q��A\�w�Y'��ߥ<��L��R�,���2�:�<�����n��S5��7
4��.oT�T���vh�j�9�puo���6Z.�ʲ��,xY��Yֈ�����<��L�fO1����>�>�ÝVL��P��E�9��i�Z��dDc�I���NRiI�uˉ{N��(Ҭo��sy�@�krs��)Ң��p�F��B�dIoe�Tn��R�u���&�ٯ��T]:"��u٭�X�����gM��v'c��2���܂�h^��&�E �O��PF�`��-�x�N�}��Ae�Oj�1�䗘�
��c�}��t�J��q5V����(���������)VV�eږ��㢱.7պo*peS�v�[���"�eÉ�F�L�!�A	���ņ��X�@p�o�]ڀ�>[���Cvl�9�zV��S.��bZx�I+����� L�W,�͵e�k�����nNS;Q�Ý��J�z���>��'.�oe+D�|6��b,[S�nlm��Ŏ��qO�f��*S�a��v��y���WG�"��;��nr��<�:t�{��X/C�s�C��{r�S#;%@N����7l��,�]Ҽ�6[��5�*��\��Ι�*�MA0��4f��
��G*>����,��/i�:�M�:��N=�����6V��,��Ύ��{��άI���{n�R�AR���i�f�#���V��Q��lò��m�#+���2���u��z���9]]ZE�2e���v"u�h��\X+n���z��g{��j
�MWD·�S��d��u�Ny���4|J!2���H�Z�6�U%55V�+F�g�v�ևg%_6�i
���j�:���JH���"�F�'c^�`�E�3��SRM0�$Th-����0����^Eyy�(�����AZx�N3�&��Ti��lݢأ�+�S��o4wrp���{�:֚�b3�l�lU���+�ѭ����jx�=�3s���F/<�ǎ)"�Ѿ<��
�|x���G����6�LY�H�T U�	��R 2U"R
��8��e�����ݞ��z8��>݌d�lh:;�
k���#���y5ݓA�d��0uF#Ag:�5�"
~1�����`�������A���ȣ�ACk:��|��ر�����>2yh��Ͷ�۸:��ݝAAG�;w?qI�H��6(��A�t�\�6�vN��N��ظ�ו�y��A%[&�cDS�n�d���Z��mc^[Z"��=�U�m�;�3��vz�_{�j��L�]<�[�t�P��0�6:0��R�1;G\����;bԺ�:�u�hA�]t��=V�M�fʷ��������.dk"��5;ׂF�2�~���R�z�Ίyl:�vTt54���e���ib�Me����D���`3��;u�0m"E����13	��x�1(U���6��,�m%��cNm��/�yS�*;5O�-UQ 1��tZ���!��9K0����%D4���I�nWb,���K���J=����=�T�/�^�=U�.&�ubS^�_d��լ{D˨,[2^$"'sѰ���yTW�"��v/ZY�K�:�2��.����:�� ���j}����cN+�0�RҺ�P��k��ڮ!�R�-w�r�=�II�;.(�d$d�lF��OX�/}sشK�1��M��Wo�ΊN��tRsx�(��{��!��6�SG��θ�o����X�ﺔ�|�D�*84z��0����)8�Qi��P��Z�1������C4�0K�̬Ӎɟ���5��_�Q�u�	�g(��ĮZ�p��u�w
�K��D�-mww��v˶FU�>�&�Cp.+�4F8PαW�h8d�/��Y���n����^ebJT�����G57�ڝO��sZ�\�ٴ�7%[�{����|�2�x��Xe^��=����f�bn����˷e�n��U֬ɱ)�d`v���Y�щ�K��}��X���`�fd����\:K�'xM�{�����Zj��uf��oe��p�ǚ3��B"��r�icw��f,��c�N�6&;����au��t�J<��fȇ��/�I��}0nF�đ��c/�u�H������l�P%�)�H�
�KX!���Լ�s���)�r��
�Ƶzc��K���.���0�Q���Y�=sC�W6�����a�K���+ߝ���y7ziGHF^Y	q���[�|��qm2S�]�Z�P�bUW= �XwL���	�WM�- �4�S`�-���R.�-BC�uC#ؕx��f&��7��e���;�i������#�zn���wp20�Wjt��&����1�0.;ڰ=�Q��)��/~��w!�ͫj��wW{0�C� H;�/F��H�'J��kX4�8C����)����)����[�ʶ�j�s8E�qO�	 ��t���)v/���8fE��S�R��-�r��6Z���r��"��IL����!�:d�@���NC��Sp����j#�T�����_*s�'mdd��Mǆ*���1L.���� �_�����Ȝj1�)�j�g�E{v1��_���`q�'K�]	����NB���(
[���F�
R� r�6���Ә8�@jjQ��+�������rEA��Ru����
=��%��}v(�V4:��*WBUFs��b��ё�i�f�+k#k_-y��V��ՅY�f����Z&;.�uq<��o5�$&�w5R��;�+�x�b^-��T��(�}4s����ȭ�r7��xL��kaS�-޹U{qcE�~b;����|��Kр븠�V��쨲��VFΒ�j���oL�ҳ��d,��\�Ý��^+2��'n5��X{b�U6���T��=��q���%�9�^�[o�iU�c��T��~�:��P=��ځp^m�=�J)QG�b�@h=ύ	��b�I��>Uw���`�dx.U�(���-/�7W���(���R��R*8�!qʮ\�S�/�w�6E\ ��w��y��U4eŚ��3���{ik�iBVhb�L��`q�Ń��\t�)�]Y�c�vl\`<�N�ǻ/�ػ`J�.71u9u�����,$B���Ω��Uy]"լ��ڞ~�����G�	q\Ae��+հ!���F�oq+hbI{���Rz���D�읪*�8\In��sQl@F"k���e��\D���䳞;y@��^��16<�Ξ&��U�`��υJ>�逶��5�7�� m:#���{y���d?�)=��|�H�aZӌq�Uܟ��N��ٻj�nýa�8����B��뮕ӣ���xd��w��FqGd��#/�J5m�%�Ա#}��ܜjf�T�����a��߳�2I����8��!�Q�����끰ZV-�QP��5[ۛ��h��įz)�]`�.�gR�Y��aXV$���8��4:�Ϯj#���\Dʜ.9V%:I��z!g��Ym��uZ��<���L�]�jV�c��f��
;��d�;�V�cGOġ�Yg�<�/�}��R�Ow�}�HFn�s�OSO�Qۻw,hM��ey��o80i��褂gL1�9�y�5��#�ɜˀU�L56Jb0��y��%]���Bh��R �+�X���0(�J�����!���}�P�?�BT_�I�w����*c�o=3�i�ny7�ǋ�;���}��ט8�#��Ok��.ڈ��fRi+�a�Rt��2u��&�9,�e�*�Uuȥ��;!��r);��-��Ʃ�s��nYsl0���4˥��Q��F��Ïb���i��Vm�O�Y���ƎHu��H���NXZU)���)���:�*�qm2���*S@��ǨBk�_Xk]���ν���6G4�b��Ɣ��JJvO)��P���Xd?0�)eA�pw���J�ƃzx޷�3b�8��E3�y΄|��&(EqU��PK�����a�XJ�wl}��1�:5 ��=���y� ���K�C&�N}�LC��Au�r��,ni]�#$+._v�Ē,�O\�� >8��+����3��n�Rm�i�fh�>�v�^���|�])}F�X�]ݛ� 4�b)�@�ɛ�dʃ�
Uo����2�p��˞�$��
���+�@;�����
���D
��IkN5�O��;�����̶�,�n��ևdn�0&���X'1��͚�bظ�cf��"No
��~f�OO[jo�&/O�4��qJ��.�3�3Fj�����r��8uم���p���^�*�w�T憦���r���wT�6��k��W���g�͸Ǉ֏?�a��:`{���͡9a���i�5�Q��F2�����4�2�}�l�XӉ@��#_b��jAD0�wE�����;"z/�Z2��>���K��>�t+9��M>�Ԃpfӣ�u����C�����N�K�l��3�|�=�Y̑�浅���&4�*y3H�	=MF02=�w>���ov�	J~޻o&��{m�U\a5}�:)3=�)�����=Xғtz�B)�	-��P���^�v�.w<{vd�tr]��,j��Y��觊����JS0�9,�m��8+>5Q%u�~2��Ͼur�:��U�ͪ�4������h@�B	��3;�}�C&��ɯ|�]�)�ƬQp���x:��%LiqG���a��{[�3,��5�������C��a���+yM&��3q-�X�R�L]��RWI�����,���W�n�u揧u9bd��m��ۭ2����|�4��i
�o�]��.o2���.��3�����w�n���c�g\G����2I�ZW@- Y2:��N9%�I�\��NoؤSe�1��S������Ei��ё�'soN�ݟ E;�mR��mdph�y��(��bU|*-?S�Y޵X�[3^9�|���8i�|TNî�oT�E���|�Ϩ��6ә�ȸ�� k�EC'���(�hjgQ��/��c�t/�(50�<z�w�=/
��`+!�0-1����u�Y�,U���&��D.�)�ݯ�*cexq[`��Đ6E��X����,�`دl>Ta�vٸW��҅2EI��,N2��=����K_��ЕG��$m��`�\�C���F��R�u�ٞ%���뜾�[K�uCq�T	T�m�S����6}C��6jg�u�\K@���V���l|�Ǚ�y�z�Y�W����V�z�r��q��^Ӎ��e�.6gb�9x�u҇7|��5qO$L0+q"�]��-��2=����]� ic�ɂ����\�55;�٩���l�1L�q��i���&�-`�5���qފrh���y�'��}����d��y]�n�-�	�>�=������s��P���;N���q=s�]�l�s���	�b��hn�f]���=T�i�Z��Ex}I�އ7.�,�wG+x�wS3��U7ZbXf�O�m�2�HvM��4�\AoY�=׍�d<��_'ظZR�j��f��<B��,U��njH�s� ���������ӥ�V��*�p��3���>��"UW��٨�zn��r�m��J�G��OZP���������b�ݯ)v/���:�q0��ʃ�f���]�6a��C��K n��>�J�h:�7�����cK%Y�,����#���9�t+�)�4���b�.���\�0���-|�2��J):���j3�%��n^��6l��r�@��Er/�[?��^:�'弬S�����ƌ�7�-փ�Y"��M�H.��isᎹ��v�p[���v#�}Nǰ*#�3d�u�PyZKM�K�3����G�Ef�������F仟nbJſ�+��L��qn�R���R��[Ω1�{,S��2��ߙ(c���wEt����%�u2��e˟��U{�a�bzo&+��%Bf����A�\�q�沨�}��O[z�d��.-!�n����b����pņ��i̱m=�L�rL��֘�iM�%j�ӏ��[P��|hO��b��0�)�-�l�\�a���wA�����T�ګ�~Nܒ��.���T��2~z�.��;E�#+�V������.c;���Qˠ�d����u������\��*ǝ?{x�Ԣ�G(�%@���p;�:�r�XX��]$=�)Yݷ����W7!�R������	a )`;s9a�w��|Y#��YcoW2h�n�1��f
su��8'مR�@Z�r�r;�e�%�Nu�`b��y��+���P�!�:�D�L,7��	a�x�;���<�d��������������
���<޵"Z�tD03�r�D�n������CFrY�<v�:0�F�ڂ���$�웽s���8��+5�}��`:>���h�#�*Q����Z)]�X�91P]5�x��T��gt@����F�
'��hrˠe�e�m�7u^��l�ճff��8"o��޹���m��#�A��$?s�o��%r�J�4���C%�����w�y��R���b�O�9�ʥ8�֯	ۭl�����k��9K�!��͵��Z�o{c ZeCf�PM�c�I���������r��̚�f���<��o8�Y>�a�3�{��G±�}�"�e�xY0i0@���F��%
��z����N7=d.I���[_j�=���|iG烷5�G��3*���I��3(�&��T�������(��ս�q�8VY�FY]��p��S�mU�A��7(�ygw(�v���ī�Z�lkc~��^�-�w&��+� ��F�^��i��&���ј*#����yi�F�P�*��ހ[r��MůC�c^����-�zP+r�:���D��y�9zJa��gy*�E�S;��V��N�W�T�G�RХ����
錦��ųKl�l�K`����D<q�_��:a�j�M�T�t�s��s�m��5��,�c��tҫi�]7Q��|�.�YO���	��@~�+�9�E>=)����w>�^�59����1[|g��\��H+�>flV`>1���g<�:Q�z�nFoFr���U�5/A��"e6�V_Kӊ�-�ip�GN�%��B|v�/�}	���2n����g
j�y:�ٝ��;v�iC_!%	���PY넺7x酂�,�	�<٪<>��O"�q��O;�-_b��:�*}L��M$�znPY^v��kP��.ƌp���Ye��9��P�7ih��v�Du��3vB�J���9tx#s��ʧ5���ʕ���7�z���Y��o�k�s]�jn����Cr,��U��[��pagx-lԣw P�h/�1n�]�œ�ܨ��%D9�~��m4�V�E"k_�w!̭�D,�����A7`�åݡ��y{0��F�c�L�v�Ks�m-VU��϶�]n�!��Ӯ��K9�Ǧ�GS�з/68�;ʘu�-3�nv�X"����umI�:/�\���Y��_.ˮap�ם��&o�-�T�4�u�
1Fb���fm�i��]Iݳ����9�?~�Ȱ�,�Ф�DEg�<d/����m͟�<�������&��.�՞M���b	K0֞6�O{!�ʯOt������k�\~ǉg�x���t�n���0�ƶo�D拇^$�cƘ�lt
���մ�'\3?�BS��Ky�ǚ�A����S�(S	���������饏�2�҉<zGuD|�S&/�@�13*'��U�n�B�T���9��Y�y�a#0)���;A\<z��RxLg#8�u�5h*l��Ucl��Q�1.⴪�n87H�c[ż��BRa���M���la��P��D������S��:y���9��������g�a"��`�%q-���䢌{�d$:�����m��Mn��3{����Zk�/%A���d�uHs ^0R�p7Z�Z��d�+y��m�R�gj���uS�Uʙt6��+Ֆ���j7z�l�I0*Ȣz}n6�&�P?,�q� �9ݕz��7-9�rYB.A*E5{�*{�4ra9���:�o�Е]1I�lAC��
.g?w��~���?/���������9�����u��W�X�tȬVΛ�%hb�O��*j˖jp�(Iv�7��^F3�j뙤l�@wi�����R9�vh���2#>�Y�Op�,=����-�d������Ӝ���N��2b���F������ct7��^�٪�;�o� ��ݭe�噝Z���ԛ�,JKѽ���oF��&�v c�R�+2�)�U��#׏��,�ewL�ƚ�+���+WMv2��-f�͹r� J&�.BQ�:i�KV�O��@����s%զ�>W���k�h����rɭ���EFl�[@b����fڸ�T�v�����:%�4�Dȯe���Wq�a��g�#�kwT�^fr
�ޅn	l��s7:�m2�g������H��Aut��t�vp�^Tfmm�޼
� m\)wLI����༒6������(kY�f�2Pޠ4����b��)�yQ�Ѧv��r��Qb;YN�Z��h5��VqyM0ފ2�68D�Ϻ��:m�Վ�M쁢�s�����q,�yja?d��bsK{C�YSh9��ᙔS���ŕ*�h���; ��K�{�k�!�Iq�8s�L�r���r�bxĚ�1a�*�6C��"�5�5P��8"�\s�e��ʹ��.���r�c*U��ţ�+AN���F�Yuf�/wxe#�/(�&��rܺ�O����VVR�U��@$"�)�P=�ڱga�e�u��Vec��dF ƌnEf3oaR�� ����M���Z�aS鎌��q��D�\�Z�Q>���m4�,��f��uw\��-a�9����;fZ.�e�L�U2q��t0~���9�3*���ۙ��%��bٻ3-G�Ӿ���YX�K
d�|�-���P7�
�b`�����-��O���m�1�""����h&��Zu��J���rѮn߳��o[FY�3*H��W`�7Fc��@Q�`�W2�"�I�NWW]����K8�ku��H2�����<Tؖ�^������#�K��2�m�(�7��ޟ����Ɗt;���0��,F��8^���R/�0V�.�q4:��GUbcT���(�c�e"%]+'
޴)�m��]*p�o��e̖�j�3�1vz�J��X�;�����X���Ed��w��N�]��(��\���7ni��ܼ��-�2N��cy��U�C ژp�TXHf҇5]�����ݹ��蛭��t�/bg��c�ح�َ3՚r�lm.�Ȳ:�+�0ġٜj-�՗�E�wy�����k6S��R�����li�u� L�����ƢA+i�*`�(
՗�ȍJ�֚�=�.gGh^���xࣚ0�x�l��u��M�fd��(��.��\��������ۓF�j��NE��2�����Ӧr˟��gs�V�N�sN��4�Uĵ�C�@��S]��oz�-�u;s��'E�{#9M�Dek����6(���A�V�����VSE0U�0��<h�z�3o4Ku��s.u&�F��ZQ�q9�P�#�\�dc����\�[�oih�fd�Q�]� U�J4Hta�BW�d�*K�R���]����}��L�i$@h|�"��N�i��n�<xc�0x^cP^d��4lb���5B�Fۣ�h;b��ZCICSEV�h<���Ŧ�C��v�1Q�<��S��G��t:|�l���hth(i���փ�:
v��N�A�u�"����������V�z���I� ��h:K����[V-[������5MQMCE$N�D����Dy�ABU3IKw�=y�M#�3�K����i��*���h*�h�;�kF-��cuܚ
Z:]S��jJ�Btj���8{wf�F&����ABD�Ĕ��������l5[)�X�ŃTt(6�A�k`���A�[`�U�n�4ttt%��g��v���=i5�:�▀2Њ,�`Z�5�Fq����$i�.��4����Ǻ��4��V�96���zpoJ����
P�6M3]f�	@�:�^|�o�x(}�������S�<��4.�*���lO3���o��x��d�`&�D�Tm\؋�b^�������C-+��V`:Z�J9OO`��N7<
41�gH��3���z�3m��㝔�t�v��bSc�����uԶ=M��/�a;�p31��<��_��s+1u��H��1B�N� �ʽ�Ҿ���e�/̜v�P�q*�K61�v�zi�g3e��[�U4�ߗ�5jP3������f'J��hl��XG��ۓ�б���1SH^�&&�D8��3k��"٥+�g�f��/�Oi��\K�I�=5Y���-���:]s��$��auV��'n2��~�`Ɯv<�N/�Y1�J��ƯN���ƛq�ݍ�|P�ETFR��ꍧ���0�Z��2��k���,�;��0�7�q�\��W�w9��6Kz�C�P�z���u2O�y+�G+q��n=�Bؤ���u����r��j%��@��Bdʆ!����|/d���.Y��j��b:M���b��u�d�-�Oٓ����)Wuro}�}�����/<ظ`W,>�����5�b|�����G{���q���SF���C��:��b�Ǌ��C�X�_I8mu�8�b�NV:�ti�j�Op�	�d��V��&���Aۛ���nQ���c>�{���&�X�{Wr7{�-�
V���XV�*T�G,��	F3&�^�x热���f�3%IR��t�K�h=�7�ׂ;fE���;@ņ���Ǳ>=Be0s��Q\�m�=�a��B9�U:O%��4��2�o�Ԧ)��J`gB����c����!�+�&�m�����2����۷Y�_���l��%�`��0.���iO0�$d�8�y�'jg֗��݂�7qe�ukөȼ,{Q\�rX�q�w�M�&S��@��b�ĪR�7o�]:� �ƕ��kdʫ�W��U9u.g��-�(�7ΘX`
�	:������[�U��-�x���(Ƿ]�6����%�]�]QMõ���؈6lf�ucQ5�f�V�f�Nm����9��ܹ<�<4����dY�0����6�_tc[׸����N�dta#Z����v�g��S�ӼX�N��&t�2b��^�qe�p���n�p�Cl����iQ��K�t�����T:%�\�G�%Mm1�;)�Xzy�Brt��y�e��|q9�%��5,R�_A��q!��H.3�r� G��9�kqsҠ%�q�%��Ea��8:8��!DKpl���wB�
��(v@����H^WsU�g��`��^B���E��?
���o
{��siZ�y�o1gL��=�.���N܋2�F�Lc8A�����"�ƃuf�,g<W&�5�W����f�QL��ꅩ���;w}β(��N\��P��C�P(ME��ʌn݈jj����A���Ӄ�WM��{)�'p�h�
��:	\B�3p�1��6"��1��O����}��Cn�M����y;ؕ�mn<��ݥt�3�v`E)��.
UQ�%z�Q�D�a�����֕=Դ��1t�6��8|�������oWz�6dH�8O�a9���H���^���Fr�^�ك2"�򤗏p��e
z���+�UE;x��6�K2��x���*��>ji�=4����ﭯ�	WS�d�<9��c�hǨ=xG*E��"S�	L&����c~�:�)�����-���Z�c�<� �Iv�tlǟCqȦX_���i��S�v���v[�������x��N�:핇�c��t6D���(�����p%���t#����P�⫓̊y}������q�,�m�/.qػ�65bI���ֆ��C;7덍���@M�}�J��/_�齼���d
���x�����w��˶��o&,�8�٩�[�r5SB��{�~�F����Y����1�ME�3����<�6�1���G|i��.[��0�-U%��~�jV%���^r��#$�wn���������J���H�.���4'ǲ��L5�V�w�r�gx��%d�+9�2[��{���{��>G2HMM.ko�NU��S��T�{Y>�rb1��d�71����`=o��w��B|5w��ur�t%�]j�R�X����cc�*ì=rVn2�2��k��3�6x�gz��	��u���m�p��8����c��?5j�R4�����F?��ܙ��~;#���(ќf�t�Q��箈}̪�3��̌�&��A��?	L�{�7P��Dwz�Ct���sf�Ve#�c#+,h�[�0�؝+.c@�g��z9��MF1���4feT3-����$%�J����ȷ��n3\�%�d�	��0�at��J¦]���<7�^(j�k���/�$��	�P��I^{0�'�	JfO@wK���tE��f{ҕj�������䱟n6��x�^n���%�L;jx��Z�ֵ��2j���M���m峍Y�'�Xׄ�s��Dv1�<�fo���a�~�;�/N1&�LH�X
�N6&�M輛N����kdSe��������j�n/E��.뇻���z�(4�΍����|0�0���bUv�%���1:VLyWo���7B�c�w�[�ؖ�䶒�hc+V��feB�c��0��zA,�(ɐ�Q�+��_6�;�9�+gX�sToy#UVvU�kw\hJt�2T�cE&,���R%hx6r��z6�#��ɍ�SMj��TNv������v(����� ���B�������̭�j�)M>T�l�p�Oú(�1��v���oJI��/��O��3�d��5��Y%�(T�}���*���iy.szGs��e�R!�U}����YS�g�8:����y���ټe=T�"%��	#R�7(��Q�v<�Ƴp�\��a� l�0[��鳟4������cf��tY�sj�Iy�׊'Ǣ�ܦ���W�ϡcE;�jIp�`��h��[fd��=y�G���/%�~��1�h]�.��xnz��Z�u[��=��=Z�J�6<=m���'@����Y�Ru:NOx�aN60�v�zO>��C����.;|��i
�GMui���M�x_Y���A̾�t���9�j1p�	LU�E�s�8]Nk �����V	j'6�uq��}G�r��X)��ĸo>K5启lZ�V4$���;̣ύZ�£���-A�*cMp���Ygm�C�xwb�c]�1�Ģ�ɐ\wK��[�N��&hְi�dkyRn6*#���d�����¢�%��kt����ҽ
	��0�?k˺��>wQ�.��
(�A�j���'��0}��k��u4��yu���}�،���]��õJ`e`�L�K�{�Φ�w75jm�a�U�N��vq�.^��)Ry]�񒫱�]ʃ���X��p�B,�rᖎLg���2,���ޠ�_��S�_^��L�� � |�x3{���^k�'���xi���O�T=��:�������Gc�$�<�c��i؎�-waJ���-[��zZ�\U�����ꎷ�ya�B���A��QI\�T�r�-K�7[Ff^,k�g��eؐ����8�g��GGE��~{e��E���D֊���&�� ��;�9�[B�ҭ�cVT0�wmZ�m��e�î���&E�E�7#2�8{�l<����Y˝�u^�Q}���x�/e�Tˋ��u�i/�jq�R�GA�⧬�LS>۴�4��{�\����E���.�yc���+�t���~�9�B��F�pb�Ẓ7Y�Vg���ޗA�_9�@~��a\jS�-#��w?R�$��az��9���j���H.[N��5_�>'��pɗ,ڮai,����e�S0��̼ͩc���Õ"�$(�6�z<��z��$�����2$�*\b����=I��U[�Y9��<e�e8��S�
��@�A�t����Ys^(�|��QL�:Kx
V�����	�q�'�2�V�p���N:A`C�c��<��o��)���F�v��u�	rz)��Yvb�+�ʔ�U袱��b쌩bT/��i��2����Ow���5Jt�Nc�/���]yӣ*�ez��y�v:BR�Z���Va��/ Z�W����}�W����x3{�����K+���� �J��ah��l�jj/�Ƣk���e��86�C�
��<�l�n���ܽ޲��Y�a�ջf��!<�
���\�/R]������ާ����p�o�;�C�0�&r��kZbqY!I�[`c@:��^z&3HJ�5�l�W��󜬁��T2s7�P�VN��������G��G�9P�e*LR�%�m�+	>�UǳC��k����El�x����&���θk���1���F��T�Yȱ��ۻ2��{�=�қ�ζIH�%�L���2�XC1�!�ȼ�b������8+yI��Sl�t0���c�뱢t��*��*�|�g���i�u�a�{:`E)�\Du�&O��L�2��L2Ls��7�9v��Mfu-�3��{���@�O׊i��*���UR&@��fRi.�iU'(2o7���}7Tw)wo-h�;+!����3��	�$��:��yfV0�T^LxP�h�����Ǌ��fճ�e������.�@v˞��h�=Aߓ�Q~"S��O6�蓐:�ma���'ndh���Mg�k��-MqV��k�\$���T?���s���m�2�a�j�L�O���n�2B��y����F�l{]wX��=i!2�ekλ*�u�;J�����LJ5\32�\�f�]�{2�}�:֏G^�u��3�ӛ�E$�ו�*R�\<���������T@�$�Z��� 7�4oR�5�kL��ŵKD[H��F�{`��RjsK���͞t5����h��v*��I	"Wk\�����0����Ϭ��X�2M�Ir�>|ck �c _R�oP�^D
��(�i������@-�k��}��~L3���l����B
�C`3�τG������J�陧iλ�㱝<��v�x��6���,ǣ�R��Xs��76�f]��	�t�C7t	��;o���)�UGiy̗[
�x:s��F_M5���¥�c���DY��N���Q���%�q��p���iY\�MX���\�rc�0	�[O��}��^9�#+�Lׯ�M�;��g��y��NK������Ӫxc(��#̺��U��Z�/�dZ�F�u+�=Cm�0S(jhxȻ��e��s� �'�n�w)�7=KM:��)Z�۹��ۄs�]tGc��M1HvU�NY�4�h�\yDf�j
5��v�(O �↿��%8�z���zA�6��d�[ی�eƧbl˴wG�9K0����-v\��Sی�8������V�f��v���+>Z�]aZ4eNR�٣ox�o����9{ϋ�*_�C��7B��ڠ��,wd�[�j�Ӵ�I��W#x�Y��d��<RP����&�ˠE���1�ǜ��y����Ht��k�q�ս��Hjkp48wf�o�<<=��x��>rA�e���b���ר_)d�EOy;sګ�l����~w��!�{�l�l�Q�k�2�N��n�b�Q�)��0;�@����$�}��&���6ZYT�imk]���<�窆��t�Cl�m�N��yQ��.(�b}�8�����c>ґx�˱�8�Nqr�m�u[[��Gq��mqe��m=��V�����BRa���l���C�\X�K_�cҨɕX.�U&y�PR+$
5l1�\\��VS�Qx��ͬy\U�K���QܕC����m�F=�,]�=	�M��� ��f�]>�0ߺN@��hkڭ��ڪ#T��{��ˬ�Nm�[�]Uʖ�W���"���6��.��ǻTX~�ע��6�8�dQ=l5u��ʂ]S����^��H��;�n�\�r�ߗk���*�jIs5�F7\�����;�4.�x�D8lm��R/`V���q�TO+L;69�:�=���c.�S!Q�u��㪨s���xhF�;5�<�S����t2������\f���phc{ح��R��8N���X����Z�[4�Y����/�n>kpMcpȶ�}]��p��!�xt!�2ValP�tH�]}Qos���"X�:�(��z��];BM8��V��P�̒�o���s��x,G:���n
���v��&���ꗛ%,ȷ�
H��7ϵ7�{�{��������]����b���?<Q�3A\��p�H�b�.s����d{����:1�b&jMw�5��&P�ߌs�l��&����J��sY����F�Qѽfv6�rl5�b��-[S)��0����L�lZ�-�&�;��ƳAnXY+��`��k����aPD'�]��'�\r�L�&S�޷�S;t��	�.&���_�a�p;^R��'����KVĄ�������.�p)zL��/X⚮�^ݩw�{����o9��v=2A�&�e�2�T骱t�Ҫ[�u`D{!�Ȫ���b���E�0���,|�:��<�X�՚��o����s�}�s�Rv�$�g���\Yc�n]2q���F����XΔB��}�S��Κ�:͗5�-��.��swO�)׸�����+i*���ѫ.W�I�
D=8���`:�(<�$d��C57^M����Qv97k�M����9�I�%>D�+���7��K���qM!�©��4����6�O<U�]�d�*��e�<B�V�)�lO�|)lȹ�b��/L��@`��������z}ޏG�����}������{T����R�mܶ�t|�c�C뤟]�(�S�s��\���Ÿ�7���P"��Ԓ��7�F9X���WgQ֌�;��sr��vJ��tޡ�]%}�bm�A*�F��RA��`�	溥vmu��j��5j�(�ʢ�lW��:�Dr�0�e�,�	͓t��޾&ɨs6�	{3\�4�o�Dc�ޢ�	�eY���W��L4��w��!��v���6��k3�G����H�*�o��]bF�9H��8�<:�'�u|+ �j��c��9Jn�кWV
�7,���eRQ7��*�ؗ:jhk$����o�T��%���Z����i���˺܃��j��0�X�b���Sf\t]Z:�C�sGR�F5N}:k�����xa/���+�oOT�������a�����|���cEDO��'�ޤv5�bR��{3u�{k\W�����B��<����o�;��s����]���^v[i(�s�
��3����\�5�c��c�����s���|~^�Ƣ�6��F��uu�����f��pW^H��Eڬr�h��|�24.���hi�=�hSv�{n�<�rQ-�-�P'J�#����M��oD�*w�s��Ǹ5�G�f��V�{�Y�ۮs%鳲��T�tU�:�ΌT7��"�'Ãݧ����!��[Qޥ�M)= :[�N�VjF$<i�(e�,�
N��>�"V�t,�h֦^R�GN+X���<P6b�1�˖�F��zuV������@��[!:�B�DVQ��u+� rֲx�?{�O�RW|e|��}��dV1�^��<6����w-}�	�Q�ux��U�rJ���khU��S�4�Z�N����|����v��X}���6�I��&�r�kv��J��R�KQ`.{v	ó3&�tQ`����vd�������sY!γ�e�UQ�U�h��g$萜�A�<Rέ��y�,�K&�oS���r��]��vaЌ{LԺ�1�ؙ�V����iY��N��?',�\QM+��ry��5�Mͳ�^A]���i�z�0K6��=���7�!��mϯ�O�-���)��]eޱҳ�8�L�F０��`�#�=�]��:͠E��鋨�wZ�P�W&���a=0jq��p�37*/���y�ˋ��nQ-a��*�k��O��;VJ�TL�t%�e?h��RXm�
Z@�Bo�g[�ś�c�U��b�,���P��Hbi-��(ŉ1���ޠ�a�<DQ���-�ڇ4�6��u��.��C��������2�ڱ&%*�Vce�tY0*�o]�nel���\�v�[vݦ��+]sKC�gp��v)f�r������m��̀t���՗��)�(\�&�����P>�P�[.�4^�I���m0��	�jтj��]uqT��������ހx~O �*�#�u�
:EAQ�·�n������q���4SQOC�[�� �4� ��M��GZ(�(���
4u��A�B�DDTAIq�:)i��lE�Ihtb�m��b֎�i�(�i��Ei7X�j*�I��4USEd�t�PQCZ1%�7m�Ԛ՚t�Zvƙ��()��lGm,KHt��7e�4���K�X�)�d:]P�ۣ]A����k�:t['A����ԝ��.�jSmU��릚�b

bi��c�B��v�TQ�LU���::u�[�E�k��"�h��b탤���j�J4��f+�d��Gv�Z���v]&����'R$�LI��%�}�&�h�9����FM�?N�xBmw^s�?k��;ޫ����Ӭd��y�B��.ĥ���x�B��m�q��I��G!CU�
Oo��xx|��xy���ie�4]��o�-�<7��}ǔ�|ZC���i����=��1�x��*V8�ǧ�5�&�8��5�id�+h�	��C�ӌ���t��X�hӋ4��R]5�~=!��ly۬(x:�b��n�;y���=���R������_�D�'����6.�J�.4�y���DV�u<wx�2���}.-���\ ����
�	`��2�[q�do=�qtMn:�����"�y��ַ��n��$i��,�h��֮1�����pRa�_�ņ�u���`����y�A���K�*�&s\_�*=�Z�>�酰�	�V[T��;�Jz�Gp�f�7{D[�L���B��묋1��l����i[�I5�1�5��.r��9�؂�3�7rE�{OEj��3��sc3�����>�mT踻n�qHZ��채µ�DE����3�\��+d�bLj�6��y�<E����>�ڦ��{�;)r�+O�z{�t�E���؂��8�{&׸�C	���J)�t|lE��!\I�x��y�s`|GaKkw����B+�U��fXoL�wKMB)�4!7jK�S9^48�ἧ&�v���f�tLzߊ��^�%��9��{}��9��Xy�@; P�α���AghV������Ǒry�}�B�UrM$v�-��}_xxx|����0���f�Ȃ-K.jo��ŠN�9���_I`���BT\%&K�g<�F9Q�co_R��5��%&4��Amy4��6�7��~�SL��{5uT��]P̤�]���R��G������<���)�f�7�i�̳�>�^f@]XP�)��UM!3�Sm��+�s����B�����.�CJ|1�Ty?��шv{Z�gm��5g<�,0�0�%R��<�[p�ܾ��eU��4�������Y��Ո춃[�#D}K�ҽ�@�-!��.-�*)������|����.�Tk�#�S��U�E1�Lb�,a� $������c�Ȧs��:������D̫�,�vV�nf"݈J�.{�%�2���F7g������؅�t�C����z��#��f�}����[n`�5y[J�kZ��ڕKU���sa��ͧ��#u�	�t��`�){�F`�zW}���l�L�?	O ��M]ܨ�;�۔��H&�Z�>�dzW����n�~-�������O�e�\)��Ș�K�|/^Ǥ�]R5�������9��}&k�l�c�xReMZ=������ٿ��W�q�g/MJ�$i�Y�����������hۥ�&ūW|(�ou��7���Q��9��:�t�!�Pwn't�s���
�|dn,�&w\�c*L�e-oǰ`�W�8���yᲆ�
{s�nn��j����Vd�gA�\b�H곷L�vwqߊ?��@ҊP�� x3x �<�"����b�w�lYD32��v$�<+p��W_��h�L�r�m�zG3�1��AVD�9)I޹l�0"�P��1�3H,C�ّ����ե�?S�b+y��3�2�Qm}8�g*H%�)��-���T�5��S���ԋ;�y����#���Lh�Źo,xj;O��84��Iꈛ��MQ���,�t�f�P�l�`ZB�y(��$�%|Pc�20��W��O;H�׫�=�1ӓ�N���t,�c�ޚ�z�2|���mGt�R��tC�_c�f�Q)�R���'1aRL�s[l�r�c�K
�&O"�u^��σ]MI�	r� ��m+'Ga����LץDQ�ˁ\�C&5����s��Ƣ ��H�H�z�v�x�T1?.�֟���_��heM2�M��ncE����Re�)E�򶣯��T%%���S`-��|"s����l����unf��M@i���u��-?J���E���:���H*�����ᵏ+�Ka,�����=�!땫�d;�(��{���T�)>n@�X�Gw�]l=�)^�֠x�h�j/�oe��у�Q����x1	(h�B�{^ˇw@e����%v�0V
f�JN����u]�fVn��ñܞ�͡�<o\g�9^VnsS��+�i�2+��R����F�s�_ee��1��]pff��Z>���?�D� �@f��f��x�ʴ��7����'�-"�4�H8UKP�r���ܶ_���$��"����.<��*���S+�g�_z���|؀�y��~��I��#%��s>�,h�|���\�R:,D�Y�����-�$g�� �����@���O~O��@��^�����.n�%j��g�c��ĸ�R�y�1&Yq��N��<�n��>���qA�t�C1x���|��:�ڻߓ�hf�K��=ݮ8x�� n���ǫHd:>H�b�R&�6�uԶ)�]ԛ��n��<3D��>v-��O �gdex�=�Z���׍CS�lU�N���@�e�`�Ӌ&�pK�tI�����`���P�Lɕnϛُ�J�c^���rd��`k4兒�(5,�$��k�ʝ��љ��Z��v���
��L踺l҄��m@��y'�]��v���Mv5�cy�n�9Q|k�wYtj�G=>r�QHI�&Xb�UP��~a�r7κ�lت�Ԅ�̫�!�=��QX���~��h��b8vR_�2*�,��Tu���0ġc�aR���(������@˝�$z�`u r�QW�<'}�7����ِt���� �l����S���Z>��!�;|����!Z�o�dY|(ީG���7 �bJS�5�(*�*v�Eyc]�86��3��0G8��5��5d�Tˬ�%�gXU-��s����D�*���C�JQf�)QJB%o  f���ڲ�A�7!n��-�}���L}�n�#��T�`���EsFL �ݘ��F�@K��_sws'h����c���'�Y"�)�qX�a�*���h���엣u�Pǌ���U����w\.��I�X�PY\ɪ¢�b>瘧�MGH�Q�U�:��@�i.�h�>5���}���k-��#��٭v�R�:�w#ٴ84�0�vr�/}0���Ys���4�����̘����Ӻ�nxȕ�w������j�ͅ�.=�<�A�P'�"����2�o��> �2��Κ���8���R��&�3
.�{eW�%E�����j�f��V���8樤��Ugxd�j��ؙݩ�O39W�O6L�4gQ�:�G
�2U�6���9Y�vkY�{P�͊�t_q�t���+ي�}�0Mͼ#.-q4��dw?���0��b!�m���a�U�C�_-���<ۓy:���S+Z��\���Ɵ(;p����tC�0kQmZH9���'a�����T'hܛͅ4�cM00Y���U�fᨘ�qC�c[�5���&��4%��c�V�yUn.���Mkm���R�pn��2=،νy�9yM�=W�5L�f{U��=���e�v)��6��z�B�.�<rϞ	{����e�5��n�#�L��]�6�z�_;�ܠ��ъ��7�A�6����Pk�c�ǜ���R��
��{�0��Z���U)@�� O��e��d�ھS�w��P���Y�д?��Q>#>�����<k��wLq���&X�غ���a����r�Z^�\��ϯN���}�>���UP���iqG˨g�sY܋�x�ώ3�]�ڑ;BG	��Az��ث�.�m0�����6ZL���r��&q�=>����駙:���hr�3	�]Y{�S����1�����B�y�k���9�;1�E:U)���}�S���6dVh~-�8�t8yW�X>u�&YJ1�
J-��ZIփO��5Fj���{�nTw@*g�½��q�v�d���F�������2T��F��w���	�I��<y]�nuQvijd!�;])4z��4#�K
�)��UL���6�^Y���	�Q���G3͜���z^�l������	C���f=�#Dq�U+Ai��
:;V���	T�޻Ψ�%�x�⎜��h��[!����;i.�΍����a�Ť<��H��g2GT{�Ĭ�MV�躎]n�E'汦9�����r�g���M�pɏ+1��ǖs�x�i�a<#���S4��ľ'F�q��u2���˸Lc�`��pRt����[�9[�t�R,�Jċ}��x�m�4����4� �00Ol`�0y
Oz�R�D�I����}�w+]��QZ6X},��h�9��j�J���i�r4\}�
H��ng�g�+G���z@�$�?Q�eA�iU������!�;{�$�P�%W'd�<����Sʎ��I1�ֆ�t�B�8/�:
��gZ�fmY��x�:����5J����Q�G7-����k�m��M�6@���ٌ���(�ő�w�6j�:}\X�������W+�_>�]O�^��f7E::��1Y<����L��-�eqKpf[-��9o��tqV������N ��X�l�X�k�c��Z�wt�g����އ)a�M��bm��	�>�BB�/X�dJ=,u�1/�K;Ȥ��⻩���Z�T�=����{]�V� �l��G�C��0��P�Tn�6�b�l�ȗ�M&qu���=���׊m�hp�s� �^!�F'J�(�3��?6��ݱ�D��ΐ��6�:fL5�|ZfUCU�6���9�_�S����b�����
y�\�P�:�i�8�ps�mX�<7�b�m�d%5��d�!)L���\�e�v�0��o|����!�R�ۓɝC�s�sQ�W�%C0�f�gas\�?Z���l��ɲǒʦ�۵}�L�5mQ��݆�'�&��Up�d���R����}�*�FP&�2O��x"�aP��g{)�K�s�79�.�8�쀏���ʭxI���@�^/�����cs�2��۲+8���me,�����ScI�n���9&b����
���� �)�T�B�B%{��EC=K�*l�)�xi��$;�XR©�!#00�UɆ�&�]��y�؀{/�i�kl`z���y�w*"��JE6P�D]�47���U����^�%&<���], ���7����n�a�l"��L�EE<"\s�I�IE��Egj���n�Ө��z�D-�ް�Ǖ�V�6�HSWF��u�%c1U;;Ič�_��"���}Ԥw:��5	WP�A�����s58}��W,������s��K�d�i��l���s�q�/غ�����+6��ڑ���%��|z��D��;@@�s��u/!g����t݊���f�8~y�B��&<�7)�:&,^s>k�7Fw��<��#�\9�I�Ú�G��aka�٪>.�0���l���� sYX�5�@��ڟ�:�*��䰹�蟾�kZ��c?�gg~�fj��|�K��=7�p�F{݌Ҍ�Qr��F��J�q��C�Α�U���r�H8i"i�W�Uϥ��Z�:<������K�L/M�FƧ�v�XcN����)kF�Z��@�hI��2S�>���M�~��Qh�+��i�Eܽ�N�;�]�U�]����C�A��iw~�q@����mn�&X	.#4�v_&~NMyX)K�Am���[�����'�e<����͌ո*Y���+	�He�"�t�f�WXy���'�Vy��/��מ_o�7�����I�R$
Ei��
�((@��=����x>�]u��^q��|6Xǭ'w|�{K�ԯuɐ\wK�ԝ�?4;�d��j�(���'"�p?)����o]'O炚j�|o(�|�!��5=��M��$�wT�M"5QX�z����ن�d�t%�9�k��;C'��%� ��ê�$��qU���m��(�n�d�㚲�V���:�j�����;Ϸ���uC��G�hDY�~��y1L1(T�X%T�ܒ�;U�qٖ�����n�����u@��z!́�.�8�`Tj�6���'Jso+�K:�f:wj�9sPg1px:܇�D�ư;���-�O�0�����B"��P�/M2=�Z��ٲ^��Cgu������V��뎦(p�m%�<�tǣ�Qkҩ6�F��͡Z���߹el������L]�K�w������)7͙�u����^;ϡ�-��E�!�OE�3(��ڦ�:���+��A�le��7��v��uh��n��冥@L�_̴�(u��*-ʽ5�`(�~!����P[֐��e�!�J=<��i��umi)�qQ̱�V�h�G(:n9�q�Q�O�s�	�2e���a���1sy�����n_��>���9j��� ]N��J"��L�(�er�s���1&�C�oN�\m�ө�bbP��\m$�X�ރ��\%G�n�k�!�2�s�x;qb�o�%X���U����S��Kme�VE�d���ę�b� {���|�	���������X��UpaWY������u���c%Y�V�$Q.y��y�5���;[>�Ղ��K�[5ڸ��I�gxԀk.�f�v�brGs��%��uj �A�(X�#ɰ�]s^$���mS���/6vZ%H�a���TS�ʢޡ�걸T�ȥ��替*�mn/m�]����?O5���튫~���d�����i�I��s�o2zt�֫B=��m���4c��-�hK��-��eyU����������{X4?=r�����]tY�f�f�'J�BI�~�|�ڕr�Y�ն�B����Fɯ� ��R_���p��x��W	Z*��.�5,P�^��2m��'^�/j����,ho3^�9��k%K��͸4�C��P(	��q~�Ʈ�{;�KuK�v��7w~�b��x��+Հ�xgQ��,�y�t �V��g4�o)0�eB���s�э�<#�Ԃmt���ll]�4ȥ!2���c�G��ؽ�x�G3%	�`���+��Yk��|������V1�8T�u�;�fMx�:�l�Y:�F��g�q��Q�Y��{���z=��_�����z�>�O�{=�>>�p&�EFĩ:�B��>��e�ۀ�O#*�.�V[��W#czI�p@�ev;���/�]���i�hJ�S�K�ش���=�l�yl�������M<p�Fc�32�Ig[Y-�g��T�"�+�TT�vƚ	\
G+Hu�v�P<�f22��Ժ�6����� ���7ǤɊAd���RLy��*Ɩ%J_;�V]+5���7��K<*Q��+MtűM�f*���.�����wk,-wC��<G���^R|�O�th�fE"�OI�<ݙ��H�3�%��h_�{�.i�!��H���J��%16k�N+��kw�:Ms/fϻӌ|�Y��* ?a�˚�����5$�F��Y�r|5�b��{��A������`=�����iIZ�r���i*�S��_>+�J��� ��R���f�V�s�4uJ���M���������)��u�i	�L�56՛��ѢἛziԨx,���
�e!��ղ�lt4J8w�^=L�aw�ֳ{Z�v:����n�!P��'.���g1W�\�KhʘN޺�W�:�s��"�[!��x�i�g<)kɍ�\|x;�pov�Uе�#;z�JtR�R��e�o�U�7^�?��*y����o��;%m�^J�9��ڲ�ctI瘬��d����p�6XT5����:D$'A&�5%yf��p!w)+�懊���Hm���L��X�
�0�rKG09��;��P��J�F��PGFv̆�i8�����I�'	��<��X��q�ҥ���J�+�ø#��֨�Q|�n�aݰ*�^s#Y��+8)��[$w�򮶺����Kʼ7�j�C.���򧋨�űdɄ�t���F,ls�|{L�;i�����ek�[]�;El�ɂj��I6Q96�x�;�7�:���;�j�)z��H��d=��ŕg}߹i�k�ir��L�˱�+25�S��Ɇ���432��N�5\hh���� Z.\�b{�C{{�u�%����m�;rca�V�Sw�Ү�6PR�s����O�T�R��m,���	�&�昞j�g`��5��)���ޫN��a�W�qP�͌�Ӟހ�^��]6��8C@7�֙�w[���{b��˱;��'7���X����[�O��ƕ̭v!UJ�ꊁ�K���.�����[+nd����W�i]���D�X{m��4�,��.f 0��*j���]�X44S�e�Nx4o����ZgHT��@�r���"%XBlp����;�Yn���X��Ɍ�5
��"5],R��5!\������b���X��=]'QMT簛z�y.(��G6��놌Je����	�
U���ۏ�1:nR�s�8u^7٢���7ݺ
.��u�)u$�Z$�^	R�l_l�e����sU����)n�c�/z�w�"���'�]ݸ{Wm,E�w�w� �E[
A6
�)�@�i� ��":
=���b>"��h��M!�b-�OM1[[��{*kI�GlN�F���f��E�QHQT�0]�qZv�&ƵmM�D�%%m�:(4h�wj����F��h��`�I�aѶi��4F��#�B[m�8��Qj-�h
���ucb�[miӢ��64����A�kZ6�l�֣�j��b�DE&�h4k];��tc`+�U5]��#�U�����vh���ėq����r���k���Tv���U���h�t��vΪ�:Ѣ�!���T��QEEC��8ƈ:�v�kb$覓Z(�щ.�]n�Uͦ�:�]�"ږ��u:+AA@ti���;4u�ulj5�MV�AѶzcILv]���hcc���)�y���̽fɜ���������B��	�|؝ qi�ѕ����̾���3��
�4ۛ��e�g�(��5�z^YX���2-�"'�Bc�È� ��
R�L"��"�}���W�}��t���/0��w�*!���D<;�S#�U2.uE6�/B�{�Ѳ����xT�#��/!մ���5Ïb���N�ac�W?j��r�!\�[��
�۠��'+3=�Be�b��$��m �<��F�H��L��U��RjsK�k��td�%;��(����K��e�N!��h��EJ��?0�)���⛼GC�:��me��B麜���̉�5֭� �ӷ�WbQ!�o>r<�nq����<���$�E8A��6�����1M���S�]�iTg9	+;��s��4ɝ��s<��n	G7-��<��˶�@f��D0QD���T;h�KS�mC������f�"L��{�|�Uu?�z݈�uN.���2��7��T>����7l���ڃb�U�@G'�>8���ʀ�f���f��jӔ����ON������~x��Ô��mk���ͤ?�^yT�_'�<����oҺ��������:�Em\��̝E�z��0W�͗�b$!ų#Y14��m,\u6�t'y���K�;UU��VvE�C��������������Q��^ͦ.��a��t��z��+�z2~I����K=�2�F�[2mKהCd��<��r<o����]g���TTz5��lx\t�-�Ž����sHIh�ʝ<���}����}ͻQ�y��o0�i	P"��"(!f��K
�*|!3m�5+���SǞ;��7�$8�y���!�ad��I�:��nũ��� �bߞ/���_��*�^��ۗ��l̙���U;Ey#H7_�h"Od&
{f(�+셃!`����� �.��Y8��^%��.&�z��#݆Y<�ERf�R�ֺ�dk�k�VUܞz�U98��f�r���2�@8W�&�A��4�R�#�u(M��<�x�9�Gbb�����ݬV���ڡ[Z+kZ�ۏL�����̣��R�H��,'���tI�(����fg뫽��\�n��/�\�G��.��ke4���7�^R��dl���#�V;�^f�S+���=��8g��K���c�*-:X5P��Z�"��zul|EH*��������jJ%�]�Oypt�~�Z��:(�f�i�k@EE��O��+	=�[#�+�m'`��� �.��S�nt��D��g<�����y���g=��l�j����v4�ƳtV�c[_Hj��'6����Γ��M���ˊ�B�;���՛b>.�[a�/^�r�ߒ2q�\K].u�>Tk
m�q�t����FAﮂD��Ă���~����Ck����+h\��Gkx_8��zEfL�d��gwn;��.+�j7C(��C��fɕ�g��[A	�^fnS��8�R#�ia��ۓZ���j��gf����.q��VmN(�R/�H�H,ʕH�#T�3  f<���b�����Z>����w��i�5�qa[5G�>.����dU��ͯٯ/�&��n���N���{��1�׌1ZƊ��6�٨��
yi��j/�(�N\h�Q5�=��7]���j�u:��ۜ���w�"2���&qO�ZAZ��pג&��H�5����Aˬ0ӗ����9�Oov8�͡�Bڸ'[e-��&�^u@�$5�;j�CO����m)�վ��p�C=H�`5ʇ��TB4v[��f�%r[�%��]��u'-ʦGv�'�ҷ�5b��O�(~;��=�UV;��R�f<Sn��3kϹ�hcx���JA�^ww/B�/P��Wo<�P1�o�=�S�&<�yC��$����^(ϩ`�[�5����|5>�߷$˿}����;�9�l�"�O�}�ɋ�˳-��@��Eс�Q��,��l� ̜壝�i�u�N�.z��m,�Z��	e��=�h�����>�ҏ+%��?:]S��
a�D���ݴ�a���Ǝ=I[�>/a��
��q�.V�c)��o
��O�zb��E��rҡ��Z��3c٣����\ޡr̴��a�VS��CF��t
����;�:8H�rii��i}����/��o�A��	[CP}+*Z̄P���Xf�����3�u15��(��z��α��i���̄�����UȲ[Ħ�꾯��徭P���e@�U��)"P@� x�|C�[���3r��X�> ��^y�W͍~��E���/��ț��9�f\��YF\�G vGY�C;F�4�'��>>z\��Y ���>�;���L��E2��O�FLdr��O�����R�!�>�FD�._��Q����؜1?����(�p�mlq��w����-��5�.�M�E-ceද+�~\.���X:S+�Ѫ�w����_&�[��I�1�0�Gr-�Սu72������H����K_W1���Uy!D���r
6���q��&v�v�ѷ��x���Э�{�T�Ë���Yφw�Hz��@�A�~g���*i��5�,s>�����|�W|�H現���l}"|k7s�exr��M#��"*&���~�'�Q�#����_�cn�CO&C�	��t�h�d�X�B�y�'3^�-XT+��bl�r���Mjft_]hh.9�`MZp��e���oZ�:<��A��z��3��
�E�/\�(��\s�:�,Y̂WX�6)�,�c9V�/\����G=�-V�US���={��L���`�Ɏl���̜˹R�����D�a2�<�W�����m�;���8�[�W��\�*� �H_�2�K��T'�G��ƙ&��:�Z�4. ��wX5�i�Լ��L���k����@���T�m��ym�z�b��.A8�
����L �?���d@���
Ph~�Wפ�ۻNs�?Ρ���"�QL�)�ܣ��I�ɦ���v�(��'���M.-(zנ�v�ׯ̡���=GdS �:a�q����9�+yIe��I�rUWKn\��ʦe�;!pt1�EL�޽���Z�r�(Z��h"��ڡ�n"=�P�8�	Q뜙��`��lj��ѵKZ�,iջ�q9!��(	f���{�N5o)d�`a�e������e�Y��X�w�5�m:��z�����V�)��!�����5��.ٴ�^lAÓjs�d��mMP��5ͳ�x�����cKS�e�����]��8�O��`����y�*̻eN6�[�8)l�<r��T��	*��`q�m������6��=�I��K��tl��.�q��2kJ��*����Ζkb*�^<���RS��������Xd?0�)����ڒ�g���L�����ڛ���4�j|C�YNa6��'$G:]:�]s(��I���$-
f��雷9�@���l`�l�^�{�H��Κ�p��d��gp�kk:�KP�@�P��i�� �iZ�.�kҶiP����9�.�M21Q��疸Aa����Xq_;�~�l���bC5��9]dǕ4"�y��i���rE�c��@���Y������gjQ
�}1�X *^�57��1'�n�Զ��qd�s����e�]�sa�R0��0��>��}B�BR�Zi�$O���c҈�����x��[����Λ%�ϭ@q�'3;�/�;��ncê=��Jد�t�t*y,�燷�:;d�3#e,�	�m�T:8�Tz�rq���\���m��*w��7���`n�Q]��p��}�r���`b��Lls��`W�(��͎���c�&��FM��q��Pt������\�z�
 �ިY�!���bhr��r�M�3U�AU{
ꭒ�vLB�'fH��k���z��J���C���Q�ܫ��`ǖx��F�����C���D�2���MF2�>-3*��n�h>��Pm�R�-�#�A�ç%HӢ��y춴D��w�7D�	6r`��.a�����5뫉����%�����,�k�mz	\����)���F��l��5T	�Ť�WEZ_��W��*��LK�U��5#�:�m��&>��S���h�h뛅�h�v�A��fo��1J�����,*�3�&c�Ì���Oo���2�I��ky�����4��C�Rsϋ���;5H�q\�Jw�M:��W��#��$�ȮdhW��~��u��n݌���ƽAT��W=y/e����?ltC��O��
ct~g�N�+84y��㷌m1��_ݓKK6��}��[��:e@������qq�]�*���uV��YMu� ��]_��f�W��n���U�[��WZ�a=Su��ﾯ����x�xx|<O��U��u�O�:�(��bUv� �Z~:�Vu���NLc���U3�0$���.���8$n�)�c�h��Zoa\{3�4ϵ�v�J�|�	P%�b�a\�iۗ���i�>%3g0��Ś��tqA�p�&<\E�wi��R���XG�ܺf�n�lK�K������b�F
w����� 
�,�Yn�@�dي�����]s/��e���hO:A��%n�tm���x̺�	:��;|��%2Sj�F�3X,���DJ�o^��t^�O\�#�иo+�j|�rU5E��;�[W�XbJgOK6}D�p��C����WD�j�]/���k�Ŭy���f�����$E��u�G�pK�	��'kK��R�n���i ᤉ�!�lt���)?��&Y3��øђ1�_˼ ,ձ�l���e�1�W#���u���םCS�mU�ҽ��L�B���۔c�K�.�d���P-9�.������Z��U�?�i����fߎ�<�q�=��T�y�Z�jt��j|��3����Nr�A{����f�7�90M�z\��4c���l�T��m�wg*�+���.�7�h�,��������bgU�����=�Ow��]a��k�C٦mlrM�W����RՒÙ��I����i�ͽ�B׻O7:�Y�"��u�V�e��k���U��RX�o���rˎ�x�7�do��U����՝ȪQ�X,+f&��ݛw����̞��N��O��΢��e�;%��"�P����ߐ���׳����͠��k�����Lqҥ�{$����,�ᄺ�R��>t���z���d�����^�S���2��QI���P���Dr��z�d��@�,a���68�Bq=��s"�;��G'�ڗn�x-��閿-�O�-�{~J�\]�VT0�yګ��AϝT�-�c׹�+��m�=�Ѓ��b���6>ƙCHw�W^�vl�I3j:��Z��TI�b�>�h�%�]�r�
XVs*T�A�s㠴�f��T���"��(�\��o{���6�p̻X�a�z8꺡��SaÎ�3QGOb��A�T[���x���n!4�[��r��(��˦�M]V�趗C�J�1�+�:��~�S��A�L��D�@�;[;����dPȢ�9���ϵs�K��t-#&O�U�,"d�9�3�$b��Xڅ�n��~,N��f/�Z���9_e�V,�1�q�_ܨ�83<]J�a[�N�]�Yͤep�V�-�+-�{�Ή!�{{��ٔ6?'�=��R��H���n�j�F8&ְ�m�*`Ø�25
ǻ�G�T2�ɾ�V��s3hsT��vr_��ĥv�̩3�c
��9DWs�ʗ�iv
܆�%1*9���V���΃��hlnGl��l�[R������^��zc�L�4>,7�폼�xLŧ먦��ORoW��V7<T��X��[�UM�\c���m@w0T��G��n�1�Sî��-"Cfr ���`@xX��Մ����1�ɞk�O׳(����P��X�K.���
��Oi�a�Y�]j��*!�!I����a�Vg����V�a�.�N�����(��}45��.��Z�޶5�E�G=��o��ѵ�z��Pڛ/��Q��@��g�ۊ�(\�����C�� ǆ�����R�fr���1��SF��*ۅ(�S���X���ۚې�ڦ��/`���T �\����p����d�!{~7�gwڥ��[����#q���ފ��>��l�k�q�;>���g)��HM�T�����*��<=��=u	���G�-=��*��`�T�P
Ǐ�zUV;�yK'��)�[�m���X��ۯ�鷳}���e�sԾ���b���0dϙg%1�4�a���}";�S-Ÿ+6{'b�(�\Oۜxխ�����L��i�a4S�ʋ^ˣP��������l-X�Ȉ�F��0#�1��n����c�;���m����n�A����r���uKCyE�����0m�`% P~�|f�:k#��Z|��u������'R����%�^u.5�-PM�0���
��]\������&^���i���� �v��|��x���)�.�M�T�j�6��zm�\���h�iT�k�=���EsNfM�R׋��c�'H}0y��*���'�����J��/����F�����bsH���l�����A}d$�'U�,�_*v���[7�9W�o���cQ�Չ'�n���
C-�w�G��q�!/��Bm������KSQ�J����7TRQ��c(,k��m��x�`�T�$��f�]��	��&	�`�,�űqbƎ��ȓ��\�E��TƂ�b{X��Merj�3�F8wDQ�x)��D;~fY��1��P��QJ98q�0�[�{��(?��Wn�튑,�^�S��s�FT��I4�-1���f6�si��XC�j�\y�Yd����O��_.�,�z�)W�3�dײ0�֝Kf�H�k�ꁬ�i#�����1����uW����=�U3�������n�����$~\C�^<D�	E'bf�<��+I{8�����R�4t[˩k^�o3�SW��F:����fFE�l"�;��A��rD��� ���y�>�W����z�^�_��yyy���_Kx::�Q�E*�{�b���zҀ�@�6p�G������K�"�)����Y7�KR�ݬ�{k���ٸ�M\���]������Hr���
�+O,�T� ]t\}���>,��U�������^_=�HGOj��ȋ&���"I����
��ft-ŊR�\U�T��⣴���f��V{3-l�GzS۟�� )i�����ʐ�}a��ƹss�h��	V��D�./y7�0$#�S��',H��ƖXm���Õ��-�;;�d���C����Ӻ�J�_���$d�j!'&�F��26�p|�n�eV=�;�m�X-�ۡ(ޚ��x%��V��&V�U�"y�i�ή ���.X�1y��%ӡ�����N���)�k��X�����8XQ��H���4��5���˾Z��9�N��ҙ�ưk/�r�2����3^U����Sk�����o&I�'M�T�6Y1�G�vK��v)�[�`vZ��t.>�ͧo��=*�Y��]�~�ـ�gۺ�2��RF��V��$"}��<��D㩚3�ޕq�{O���DVf0��-(�#�eEcͼ�}sk2u�̈Vgb$Q��7��|y�(�b���M�-��6�Ҳ[E 7r��	fnj��.ِ��h���L�ێص¹+��*[[�r�VM�0�i�f��F�-S�%�*����S}������/�t�\�䔡�V�_]Ǳ���
�Eiʶ"T�*�`	�)�*�E���v퓙 �n�QI�[�����%X환K�E��nm�b��i�^��7o����V�,>�/k����4&[��(��_��*1i��u��Ƕ�%�8`��Dzu�xDA�TW���@����g�6��^G���]:t�Ԕ�N3�	�t���Z��R�|�����5��uChT�f±��qIU)��1lh�G�7�6�ЋyUa�|Ɛ�z(����f�$W=�����u�zU����\��\G�2�:��Z�`�q�#���*��w��jJU��vͭ(VgX�"������Ol�Q�b
����O�j1ô�V�ǃP2�� ^�M�����F����%��[h�w!��;jSZ�)V�\��~̬��VpMtL�"l�R|�q���VU��z�����m�4�b����)�^T���u�p� a�������`�2ݚ�tgM�H�6V��(�8���.�)9��W�%972����F�9f���E.3���t=�@&m�Cul�z�1�EN��M�ϙ�m<������@�	��d�꼨��cOw�3��n%Y�^NyК��Y�p�|)[��C9��Y�h*r�6��y�r��2�4�{�ft�ӄ���\��Ԭ<^�Z�ة�ޙ�b�XzS/i�ge���y�g0\���d���$[ܺ�vl�Ԋ.;7�6��
����F�i����ܛ�:�DZ�6�|.�rb���PF� �cPִի4�/7TE&��X�c��m�N�;gm�6�]ں)�4W�qb��ӈ�cl�66�1'��OY�l�ڏ-E�h�AM�UAZJ���c�Il��5֝i��]V�#ɢ��@h֍Q���Zt�Q�N�h�EZ������1�أ[19�mۢz�۸��mw���[e�����5�&��lUնi4:�;4*�U5夢"�����l�4֨�Yֵe�1Q��k�WY#h��OEV�5��[�i5�l�Zk���X�NmAlhm�AѶ�8�1��M�UN�F�h��A���QgTS�1$��C��iъ-�M6�����qj#EQ�u�,AZ�1V�ٶ���ŵ���<��͢�"�֎�T��x�U�5OZ"յ��3b��F퉪���Lh߀���|���ړ��]{]�r�Է
�n+�j���j�iXa�b���V,�Z���s5���[)|.��<=屲ݒɹr��M��@�y�)��q�x��S]Ͱ�J���<O��̟wJ��vv�)~ˌ�E�'*Ů�=�p�=cK3at��UI�󉆧nq|����B��f��-7��rR�ͼ�ʙ\Y$f�6��^}�(��ra��=��	I�=.* f�H�{Xq��`�;�dl���חC�y��[׻����E'�P%��9�k�1�o!�XP�Д�~�,v̠����nknnAT�Jv���w�Z�����؂�M���Ei�kW������ްM�/�Z��-W��n�ESO�E�'4�f�/z���u�V[=�.�"�=OI�ZT	z�Ŵ8G����%��LՌY�mchEz����n�u`�q)���迮��_��EՀ�=�b��g�PO�'p�B�E�Mp�ˑ���$XKY��[�6z;���9��H�~�[;�t&xjػ�3�2�7��δc���Lv��-d�^)I���Kp�٪��j�Q���p�ҋZxD�.�0���U�΋^ERa�)�t��g�u�f��a��p&�K0���SkZ}�����z,F�Hwe��:�q�:P�﷩ͨh����+�ʴ�dCN[�_瑵�;��+��y����h�#i�Zӝ�F�z�4����ovV��h��j���#��A̔bqU����!�x�6��</4^mrJ�	Z����z�^��IܺM|.O?�+�u��u8�)���B�!�<��f;�AZ�Q���.����&��K����Y�b���Dܶp������]��O���m��1��@���(��&�F)4�J�SM�g���+�R`e"��S�Zw����T����'$1�.�	�n��+*y
3�o-wq�U	�s4� bt��0{Ns�w��;�nO��3"a��	�<���,���5�1�Tn�iwKI.3f��)v/�=�:���g�E!���I�j�E�W^����2��	B��Tp7�#:;Y'�yd���*Z��o0{n8l���c�T�9v���R:�)���c��_����ie
�gKj�t��� ����=}�Mm{�Vl0��㉒xWK�;Y���lw�Fo�s�[�lb����q{P�z�T��%���r�^(�H�#xN�i,wJ�S�.��S�m[=F鯦})>�	O��T+�1�i=o,�'-n#�Q^y�|ڠ�l��!԰aYΩ1�{.�h-9�	���X�~��zU����&��K@�J:g(�~ϋ��%����Q�3���N��yun��Y�o���=���+^�3�e������Ϻ]t��?��b^uʄ������ ��58���>RY9����ݵ��1˞>�nX�4]����yd&�ya�{�X�w"Gq���#mt<����@`�<A���UTx1�y�[j꺃K�-���\k����1v͇���\\{ �A�QI�Uf��s���+��Ɔ޹�z�Ȋ�·�p�<1�	�-�1�@�Ԅ76Iՠ�h�G M� a�5SC��Xy9���'Z��ӥ��U�J\Y�<Ò2[�x��\�J����
%�泑�h1��-Z�̾C(-��31������B��N761:#��X*K	�)�Z�;y�����E����J���� �>�OS0'2��OQoP�uY�v�4�gظ+�I�����l�#�g��.:|�X�A�t��`��'6�B��K��=Ԩ�9��8�ky�����J'�a��D����ۆG`{�8&�8�&Ɯ3��j�G���)9B���c(�~�;{�۫�C5��l,��h	U&�b���(�}sQ��a��2k$��"e�ښ�5�m�n>t��0���
-.����GU�|���<��9�(������-5��4Y]p�*�5�ܓs%�.��hnmSc^:c�EB���S��'�C��v-�z�^�=��o��v�8b���fV��S�3�N����<�kD�^T�R�gT�C�Fޭ�e(�
���꼝}*N�ʳ�be��jjqifC��_
���#��Q��㜁��O�G0uoMt]���aY��بbuÅc{�v�*!�x#;3S| ��j���'�c���+1��� t8��w��7�0p��n/��ҪD��kȨ���k���h�ia��ٝi��p�	I&L�V<�d6
������ɥ�飜�*�<�v�I�s;u�1�ҍꇺhS^q�@�b�ћ�����Ri*0d�,Ԧ8�XO[���XM�O��r]�z��TF.m��b\�<��\�	�Q}0(�up͍���ϲq|QKA,�e�� �B�sWb��3�� �Е.r�	��f��mY�u�C��d��,�`�{�F�.��وs��+�c��x�:s�Z�e����\1�<]:��(v�j�n���~k� �<�ENt�(���d/f��{[����{�<�*"�T�2s^ȖS��Nޞ�b�P�ќ�-�׫�f(�j+ز�o@�����'�bk:��T�=���XKM�z�['ۊ�[Je���)(��Q�v��.M�=��R���2����F�J����:/�����_��X���K]�u?b�3+�4%���:ϷO����x���^� @���kp�B���9�ݪ�P(�dza�Ů�#m�F���{{�����l�nn21�y�19�w�2ʫ�.3c|�{�=��N!1𫐷�❽&Y-�R�Lj�[YV�Quu�(���Do�W��Q��tH4�i�L!�'��U�&�vN"G��ᲩL�X�m�{!�{D\�l> xVf(��C�m9�\ϻ���2f� ��w��2���M�<�w���a�Ӝ_.��rgf��o|�f�þ����`7;#Z������]J߮?��)A
�V�FW3H�X;l����N#+7;��,y��[�t��˸��ۄrN��q�3C��N����켊��C��r�4�8���)i���1�����QڑM���ۻ��&Y�BRC.P�)�_�1#ytm�{��z4��6Z��U���=�U�b���{�����1)�P�Y<�f�\x��j�����܇X�NMDۮ;0Cִ�3�P��UI׽��U3��j�ʺ[��h(���e�I;���D.�X����<f;� �u="���&/�@�3����aU��)v�9I��ݒ�l]��B�y)
D,)c��n��.�K$W8�P7��L��Wղ=[��h���ȗS�U2n���c#sM`�+#��*R��ҥk�*-99���Z�a�@�ztgzo+2�!��.��	�_|�����K��X��Zo!_3�4��Qa='Ϳ%@�`'F�381Q�3j�j�7�B�\����c�X�&s)6v��L�mQ�WYp׹�C+�P������5qJ��
qq߫!�R�)yᵀh���P����Z}�cP�ox8;B��DCgO.�1�
h�.�g[HN�O*I�
�s�U�W�5�V�D���3�'�>��h�p���N�а�q3xa������^pOZaATM�f������7\�/��6�$�dQ=l6���P?,��8|Y_*br�}^���ֹw��ޘd2�L(��e;E�v�������-	U�I�3X'�nl��j4K�zenO]��|~�&]xd��{ܩ0ձ͉�fϮh{װoԽa����uA�}������'M)ɼ;Tgh#/,��W��{+���L����(У��<��麫Y�-7���[q��֝����V���Fla�-��� ��_*�"�2\\i��ț��D�t5�dl^�,��7�x�R�S�W	���bY�4�o8\w�S�G\d�ϳU����U�T�*]|w�*��6�.',AfX���R�q�ڢ+ک�u�T�?�
i��{�fd�6�+.u��B����Dʜ(v�i6�B�hwL1O��@��g�����2����y^�]�i\����0�[�b)UC޿P�
�y0�Q���>s�&/�ve�-介�#�/߬d�0`~S]5se�/@��+|����~�Zih��,y�ҩ���t�z
�c�ˏv�)\q��4�ә��*���.��{���W����Foh�m˭�Z��̾��{��CN�ӕqT�r�YYv�*9J����{��t�4d?�	A"�A����L�dV��=�r}�o \�0��:���)sj)>�r'5���/=P��O@�+f]�N��Ut⺐����cg*eg(64��vz.{[�oн���1]ϮN�~n��̳o�Gv2;q�OG��LcH�8�s�wU��&�U&�9�\��>D��i�[	yg6ܿ-��jCm��T�چ�z��L���:�{ T���f�P��1�̚n�Q���z���v�n�Q� ����,��PY�clI�Ɋ�Ԣ�nb{��'����񫕜z�l��W��Å��!�ERa^&�1O�s�#�e���gdst��ͅ�p��э�/	�8��&�\��Is�z�o:ej�d%�e�T	�Re�u)��Y���x�J��8 �k m�_R	�~���z�ͩgQ~vl\c����${Fd�R�qt�r�;�e�%�!0��{��7���fC���(�a!�\|	)���cK���S�]e�`��2ʞ{���R�7�S�DkMT��Vҩ��Q����G5��m���=�ɹ�Lk�W3� 9��5���.#Z�Ϭ^p
�� [Ǐ5R
�3^�*�s�t�l�vr�o|Q����QR�W����6�:�G|��a�}�뫁Eq��o�eXў��ƺtg2#; �S�2+�ԭ�	5Vr���̧+(j�pDI��M�T�GSk7x-�&��5s9�[P+����}�9��nSG���δ[�I�-A�	v4:6�p�����8{z���*�5�1�_@�:_��oNK_
M�xt;�®�k��<`d�S`1R�ޅ`�3�ۿ������_�WXFĩ���l���we�k�A���E��5,S൴��H�h(_�����3�4t�c_}�;���Ճˢ}�ul֍g��9��3~����]��cgN����g4;"�?�,�4+]�TG�'2��]%�6����1t=����LF�C��ވ6g՚�@�q��wL�[�<���h@�׺b��3�љ��˵BT_�)2\��a��*c���*�=�7=��9�i9B\6!�N�j��9z�D-פ��{i,�x��mRW��^J��-�f9ƱK���j�&����u;��^�)����UL����n:�(���M;�e�Е���!ǹ�7�]�P�K�)V�Y�*���j^�^S�
�M݉U�ǩe~�3p���ql�4��ϴ{5�Z)m��&��;g#g��Bn��������Qq@�*���f��b~n����5�RR��;'W=lS'�5��[�c�W�1��^ԕ������=�:��&��bEP@�k�7r `a	a�f�黒�����/5�����q�x��1y����S���kU�F�Y���m��kX]�R�T�}ݦ�ꨧ����UW�n}�o�H߃���و�}jT6�V0�e��pޯq/"'��On`�\�k��l:p���.����.xr���(AYhs�X�zbsg��.��'�6�jB� Z��'��e�l9B�iZ��z�"����	��͚������Wx�L�(J���{D��V`�z���W��T�Ly|ȋ1�)���:���{<�\'m�^��s�sTox�#���S�ƍ%����{d�֡Ф��3�z:FMN�y��R���r�qK�nD5����H*%Mf���_ @��t1�#�����C`a�Ju(���@���(��H��ݾ@�عCr���k�㥮�n'+,Z����
�h�MF�\�s6�7hc�x�^lI^�@���W�hU̾�̮�W)]�Ғ��g,��:���T���>�̪���Ɲ�(A�s ����m+P�Sv��QBt�'��)�{���1BW���S.Kg(���T�g�2��|�w�}���pͽV�ה�ͯʢZ��؅<�ZJ�q�玣�]��b�-������JV�p�C��~������a�#q>����0\���E������ncym:��T�ϧ)�_x��w.�X��Ʊ�QXL�+�N� 9a�c���DnI�6H� �ݝ�^�N.��}�+N�š�vk���V�sк�n��2���M!�^:���N7�64dS��o��ē��i����TJ׳��&��ɯB+n۰-�j�SL����)2�츪pEOh�NOuE�N�9�ݥ��ւ������+����|Dͧ86��J��'��}���P�ݤh"*gY���/��夙Dp�mia��vn�!��O0�?)EŹ�Q�f<yN�GGH��J��{Ρ�44����D��(�s�9��ީ��C�i?�X�5��KU^J(�si�f���Qʯ.�riFO%�s�5�Rn��o�n������^@������sx27;����CL؛3�wz鷗]�PeG��tY��ۑ��1$�Y]u���f(����[B��w�(U3��m�:���A����S�T��1%���P)�(lRH۵��'��f�.]gk��ln*M�m7������A2+ %Ra��p�P:����`V����`F�%D�Ź�EgCjk���S�+AUKl0똬zO#���8��,���@�H��U�f�ڋ�L��dۨTgS��L� �Б0�f$Okq�il )�Z�/�f=�ݡ��1t�@�,3@��w���������W�{=�>>o_�Bݗ�LCN�4�.�fih@�s-p�mvh�I���%�M*�����m��(�������՜;�U���SZ.Su�f��m�LY�tOG�߹�R��a&��P�lI�����;�)`�y�!����ɢ�7Q��	�n��x���Q�f̀ڄu�XO��N
�ŭ��R�e�z�-=��%�;��8�m�0r������2Mv�ķ���S$�l��0)`�����n9�$f�c����g5]`������V��|�����t��5�ܕ"�]�R˦VfG]'�b�.'>��`�I�˲�9-oPg=.���v���p�羌391�J�K�odi:��l������kv����e����4��Uۺg=��h��,:Ј+h��[ ]'�*�ʁ2T�7T���7yß]�qy�e��si�v�'p=ky`��"iN�;�qU���X����ݜ)�	ai_mJ�}���U�+�>%�ܷ�mZ�"�V���R_��4�w�՝�t���`�$<��9n��X�٪��X2H)͕�F���]�,.u�:9��gt6�b��3;�'<l(I�J{�"��n�L>C�-354F
ˋ���pucK V�X�+���5���o�Y��ُVaf�G]�3�pn[��ws�CkV�r��oډ�Y%DM�y]'B��z.dם�T(���l���nX��v���j��2�Ր���at8��q<�ih{R\d������2I�T��ST�v^fE�r,��e�:}I�hmJL�iW!��i�D`��Ȑ��7D]k���IlV跇u�=ǂ'u�uµ29;΍ia��SMyK!�r�����k@��ǍnթZ1AS6p��[$�:�n�2HHl��W�S-�/3�<9�}6�M��xd��ܹ.�w(�S7�.��.�U3����α��i	��w8�l��Ħ��YyW|�iVR���k�#uK�;�����1/�X�u���Ug���P�&�	pf���V���À�-�9�V
��[��u;/���ݳ��,>w��y������CP4*^<z��J������V@�s����
we�le	T��r��]��{3���ulqv�W�
��If���Z��3u�X�q�鸬�\�
\T̊n�ǝ��� N
���Mǜf2Ӧ0.�U��p����f͚�V�1f JN�];�o<�g*4�3��:����&2�rnv�{����X��C'4��R�lׄ��Q���<+��hu7\;���,j��81w! :QZ�u�����-ï�c6+�Ӈh��
egS��N��|M�y[R��mQ齁�r�p���iQ�����$�m�mʳ�N��.*Ͷ�ylU��o�N��H��rY��� ��5�Z������N��Ӂ�M�rN���l�kA}2赹Q�7�E�C�޵F���uljV��Y/.Tz��N���7$,���(+k.\b��㚜H;[)� c�t�&�S� �RϏ���ž��v��u�wa����H|��DM�lF��Uj�k[T`�ӭ?m���ءӣcQN���ۤ��h4cllm��;E���ň(��l[kZ+lLy��#5��::�1b�cf'l�6�[c�$�Ƴ�-�m����1���b�Lh�l[TQ��cOm]:�,u�Z��kgV՟1��m��Z��hԕIF�GZ�1Ql�3��t��[��v΋:����(�/#���"���A[X�ELV�kE�ն�Q�`��$�5ۻCU؈��1hlo;�6+3i��PZ��h�,ƍO�QD\v{N+�V�;j�E�1��D�q�Y��1y���MUZ�S��b�h�ƚ�����f"*"+Z*'F�Z�� ��N"���Y5u�8�mT�QcDm�����j6�E4cb��5w���v�WgQ�Ub+hu�SIti����ݶ�;u���!y$H%,I�2'.��N�A�Q�gۼ�N4Vͦ�V���A�����V��+	qP�y}�o�ۣ�k�ur������l�����%o��|���F'J�`m0�"�5���qz�g`]��/[�l�"kvI���d<U_`�iT瞒�w96�6_L��P/��,��4���:M��S����������s{rZm�z#��jvA(�P���mFpi%�t��ЗV7��8�!N0�ur�l�����_��t>��:��:��L8�F��fav�Cr��s��+��׶I���&/�ʖ�`ޘg�w[�9bZ1S��^�	@l����o"�M��P��{�e/Vzl�`Y"v�5�)�뗇�����̻5`d�<�[9W+�൝(�m�S���Mƍ��x�mm<�k�����br� �Ue�fs�]����?�w�n���e����-G%ܦ�ܳVڭb�&�XxRX������%�g��]�b�w�+��M����f)ֲ�LC�A[Ω1�{.��Aiͺ�qI�ᖭ��L����9@ ş�t����)��ħ�*�Xۓ7��͜tݡ�g����	+͗e�SN�&8�]��n��N:ii׊�a1O~u�}��p����M]s����h�G
�оզ���]˫�"�Nc7�p�r�x���F��+�dcXwxV`ۮ���v*/���hS�"V�:HKI���B����'�u�;�Lȋ���4�L�?[��(F�.��m�ϱ���!�V����m�����IG�Wϡ���WgTrGy����u�}�Su6��=�[&d���<��U�hˊ���"Gv���[1�q0U��h��������ӕ�����'�����U��T��G�x&��%R���ӕ���,%� �� �FҷsT�ltn����!r��j �=���ĂP����^Y_N�oqP�I|��[�;ؗnU��i�3�Z{� яƢܣQ4�mB�p��"CfrY���v��hz,'�\���*.��/mN�ƹ��'\2;����ᑴ�p���9~TC��e�p�+�(h�2x���
Zױ*��pY�	·u���c���F3���_���U(��7���o�|鍌f���k s�4���D��&бUN����+q����C���Ag<����0��s�s<�LL��ڶ{-�7	{`�e}���5
Tc ]Ôr�ҙX����`ԉ�]Ygs��@�p��f��!^D��c~|lE��P�����c���'�q��m%l�B-z;�Օ
���-�_kȪ�Q#���%&I�h3��d0=��y��_1�(��tl�Ҡe�}r���9|#[Md<&���0��=Ȯ�r�2�G)�S���N�}{|�PmjKy����������:;�,]<��)LV��6�� �O�A����j�^�[��Iisz�՝��*N+{��u��x�NO����M�H%4�oc{i%��3r_��'0����.���W�5�a��Ͼ����x�9�Ė�Ye���'85M���Q�7�K��K���Qk�tj��e�1�Ϋ��݆"�v�u�Fy��ʨ=�H���Jr�ʩM������y�<e@jh�,S�Aރ�M�*�UC�v�.�ص	Bu{ &��-^^e5��5Oʎ�Ñ��K�D;aY��*�c|#���Q�8��?����me�K)ʝ��LH���On����1m&��^UKF�x��"V�@�qhP�
�C`:l ������������>�0��m����|ٻ�-��i���A(��lJ_/��do{J���s��˼c/�t���=]�,EM��}{�̍���zOT�~�5Ig�Y^v�&�Z�$d�0����0��5�smڧj�����lL�,���U	���'���J�7dF'�1�dy�ծ��׏n���mk�3n�+˖����Q]���l�X !�:�"�@��*R��q��6d���N��w�Q���*�g׆�S3	��
��m4�s8�����W��4��ҶJ�:�����R����%Y�l��L��Ҝ�i;B�򉦵Ln�B5s�#˘�fn�砐��l˱-*qǶ2׏�	�f;���ǩ���[�d��.����fZ��P��aT#��	�ۻa��҉�����O�0�4���v�@�i=ڭ��8-�Dxp�ڙ�VnL��(昻��S�)��z��C�J�����S���O��%�������O�&:�ɟ}�OJh	����H���Mk��^�id���eLJ��ͩ�{�,�F��;�PcSWcc�6�W���j��0��\d�k�R��W^�>�D?��Y��xCJ�5jF�_�)@FH���y}�]�mfe��M� u�P�t�����&�Q,[,�M��4Yߝ��
�%��%׈�ۤ�͟�N����Խ�5�_l��=u�Rsϋ����F��ߔf=QS�����ȗ�'����Q���-�<Д����,޶1�T.p�A�g\����U���L�؄3m����v��E�l�][[zZ�j!�q 7�Q�n!���|(���6b*z���u�*�sme�ʍz����X��\��y�^y�1��x\�P��ǋ��tJ�F�wK�U\�D5;�"�Rs�2�r����(�b`s��>���\-��,��f��z{*�ޣq����
�v��B�C ���&S��Z�hQ4��%z�:���z5,@�c {�n�g���;
�b:�fS����)Rk�-����T�U���߀}b��q7+*L����;��k�*F�w3����-�}�oF� ��.Wv�T���4w�u��qJ��7)�=�����1�@X�N�[H�J�<��n=�5��*vk�coT��wu/:���zyP��L6�O3���>i���=Z�J�X�3z�	fvj��(�Q"n����C-+�52�fZ�/I��:hu�3����thc_�@{S3�dN�_��|�����}pZWj �o$M1r]ٰ�l�X�g�hj������c%(/|�w#�z�����׶�D���/���MOǥ3�Y;�*��~TBZ���tS�͌wݻ^��傪=��'g�ݞ;s31=igx�W2�3\�����h-�'J�`��V�g�d;;'9M�-h��u�Xn�S▀�hW#W�Pq�\�O(Y��`wT1N;^R���g�ѝamQ==�V	�Wo������5	3e
�xcm����W��jc�K��;E�>~�}�@~�٧�]V���]S� ��x}n�8�U�E�]�v{�-z~�A����(%�(�F��5�O-�����O @�����o)��T;,�f~!��:>L�<��/�<W���M+�<1E'�i,hG%4����q=�t�?ct���LهRY��g�Xm+��$�Y�>�w��"51��>W�RЋ=R�hp�ID�Um��֎��Wf�5'cK���f[JӶ�������̎Z�N��wT1Gcd�o7{�'�c��Ħ+\�q�~靚�̖�i��_����qw��$^B;���|޽��a��i���{:`[�m����V�;��VJZLVe�.פ�gmt��2⯥����� �
XV�*Ltr�^q��&����&zX�e���lqkv�A�y$�M�a��.�̢�s�����ڑm��^ņ�j!���|GJ0dZ����c���]��Hh��0r�Jn/��Je�D�v��J��ھ�,�.���ȹ����X�瘳�������k@��8�z[�G�ڮ`��ːs<��3�<�qR��e��{��v��#�+�K�ǡ٭q�L�'0��4+�Uq��ө�dw>4�og�M���΍9m�A`��e�90��a��5�;����y��'O�aH��̶P����\�^�uk�U<}��
�zH4N���g��!@�ҥ���l&����'T��s[v���f��e�`BD�j<;Zi�&��Ԡ>��:�̶��	�N��`�\3��jU}\[�������ًK*#A�]:h��1�m��P�*�XQ.;�8ƴ9e�2�2ض�yr�#�x����*Y�J(q��9;����>����Ыm��ĥ�iiM�.����ڜ���Yc��3�}>�����Ӵ覥��c/;x���y�f\e�d�l\n�Ym mۂ��n�n�Y7bu���t|J���;Y=�o��˺s\���Gӓ��=6�D��aUN���Kykh748�"RqL��ܦ��i�H����mǥ*�����39�4�B5�v�E*8������,a�t4D��w1����W8w~�
F��}q
y�����N�ٮ�n���U���=۹������g�Dmc��(%t+^�8�ȪÕ���I��g<�d(��7����s�L�n�������4Ӧ�I���1M2��}q��"���<�K�@�jd��L�x��1�^J������F�Ct�"Ja��g%Tȹ�w*��r��ytKS�)���%$���-*e<��_#�,ު8N[�^��f}XkƶU��n\�m=��.�\9�D���y,�;��Iv�.��и��Xqi�ix�.8�*)��R}k���e��^س�y���@�ri���0`WPg�)����=�ٱ,w�zo����*�<X�+����tGtf�k��l�z�Ps�[lƭI1�˭p�&����H�ss�����s�)��҉;s/�ƽ�1Ql���e*�*P�m�$�������т�����}��1h��L�XHAC��X��,�F6��&�� �}�YS;b�T�ͩ�Ւ��i��W�h���>t���ѷ����6GX�b��&��"[Jf�8���:�[����W�g����������9��%t��-k��v�0	�&-�d�y���U��3b]�L������cA�z�\��T��rY��j�S�p$[�����Y��'u��ziu� ���e��2�7a�����f�cV���/�v5�Ƀ;$�c p��j�����z[7SdO��9s��3%^7\��cCYn;�=tf��ff8B���]=,���Ƭ��ږΣew�a��h�8�^n'OR\��X{-�^D3"�&W6ƹ�j�n���;0����N��X-QY�o;;j�oY��q���de���>x�fk�|�D�Y��N�n�[������ʡ�B�I��n��u>:��|e�K݅�r�v4��;=5Cp՘��6�}�E���s��h%~0�|��RY�Am��mO;1���؃
���qe�qkd<p����ϟ��{:R�d�x�*�fV.�vW�L�S��N��c�na�&��Af�+���@t�(A4�()Y�n��Y�Y�Z}��G�ev���6��n]T�ڹʹK;B�mJp���������w��4�b��X�_	��m9K*L�wB�U����J�o����)�c{R&��O߃�@����o�m �S����~8���6��Q}�C�%avPJ�vd�����u�%�d5em�8� ���r��["�8]�>Ի4�>9�´4mN]�3u�qH�^lT���B���&���}���z���]��"�f�7��x�A<�u6ܹu���%�y�P׌}�t�t�o���A'������<�=a��뒮�:1 �t��~K[/pm^�uB���\��έ����f�;�>�܊��ǕfE�Gh�+|��i�ԫ�IR���@F����l;�lz�����[��<��vD"�\�򚌞��|���I��dw0e d3�,�L
���#�p&�fi�WRw�Ne���FT)`RuG2�V���_ֺ;���W�HEN�w�OOs;[�ۦwv�����_6��|��X�M�)u��^�|�y��������}��'��+(y�^�b�J$W�W �ӧͼ����!N����T��8;��U���P�yi�֦�^�m����C����)��T�3+��8��ڋ^���Ǯax,�j�1˫�~ݥ&��P�y��ʮ��������2fa��=���Ź$3����%��Sj��8e�Ѻ����SE���֛��z`]�f(+8�Dd�*r�7��9S�����-��8�9��cVa�'"\>���Wv%�;PQ"�`�Km�قv�m�vT.���D[�:�9l�dd��U���jE`��B��)�O{,`�~��=���u�wl����f�ϴ�@�mR�p8�d�Hd��I�Ѣ]��y�*i�z<C�=w�ǒK<6uT�`�yxǭ�e�M�!ԙ���t��\�12��������q5L����t���+�˼���Og��`<O�~{O�������g4���
����ͷ�h�H�d�R���M���֢&4u6�Es!�m���d3�O��ϡ5�=jb����W+R]�op[�.�I�W<��+�؊���X��fvX 2�v�w(���g��%(���H�^���z���O�����=������z�;�cAk�˨��G��=�[�;�+�_��h��t�i�ζe��.	���c�n-eP7��jXF�)� ��K-��>���8��`����M�x�L�ճ[O�S4��w>phs[�C ūf!S�o��X�9Ȫ�A����<�0%8��բF��	+����r�N켮�SB�����|�1�]c�;���(*�����Ӏ�M�N�ef���q��>L�ttfē���9�d*tk-p�*�����u����{�rP|���i�yL���ѵ�᭚Q��
U�n���������aEY@j���S���Z8�|񉚚�f*q=o�`m��JuO��BQ�w9%�� ��[��N;�r�CV��yiZ�\�}O�s�U;�sTz����ش���nrS��;g��6ot.��2�]Y#M
aʷ�L�.��P�Sû[��靫�O&wU��;���̻�3��E����Uݘ�<jq��T�B��ȅ�Ƴ�P���]N���T"��tޡ���Za���q;���S.�(��Z=��T%���2$�K)yh<Qu]�ym�[�,���s������0�:�vo5��Q�6h
zp��eLP^5\�(�[�y��^��Qw:�6��rQI�!c����@�Ե\��u��U�'�(@�F��e�����ƌ��0M���Rꍆ9����2����5]h�(=TͅW�CoHvuw�\9S�
7:P[�]3�g\W�W�f"4'\/n�{jl��*�������P%��(�r����w�\�c�}ݬ�d�y+���Goir�4{X��R��h�c�wtU�B�[��VB2 c$�	m�肯������֠�^X�3�⭸2(����L�q�Umq��qvqsi�7Y��vem��o*V�N���n)�܌�a���{��cɖ�n��d���Ie��D(gkK� �d�A�R�r�5��e�s�y�ѳ�:3���˩�����U8eq�3��\|�>��)��1]���n��k3��frR���.
�nL�,Su��^E}��WJ�ka����\�Ƙ:+lM�=�M`���h93�P���+q`�<d�y6���@�/��ph΁�"���ܔ��#�:m	���m
繻R�tu�>ە�@m��ԛ�$X��y�@Q�Y���i��5��'a�K�O.�6��E��s��v[�R:�ZC6�N���F2����;�cS��o�uph�{39nV����:�d�[/�QM��5��Aon�L�7���W��������]�^��*}»nכ,�mۘ����j)_Z�Q��]�̞��GǊ%����k;�
�9�N��0ҩu/+I$o=��ν�ט5�;;3W'�A�u٩�$�xDn��4�*�����&<�wLZ�Fa�ї7y�P�*Ka���\ԗҞ�h(�k1ج����3=`K���$�n�8����-e����T�i�ky-o+rL2�H�ͮ���YtCkm[j������gkU��kmՠ�[}N��cƒ������E3b�����Uˊ��f�f�MUkm��N�6�"i�'y�t۸�[5EF�&���(�l�
��]�Qm��#����-��6��
�ۭGX�mY֢v�[f�NI؛��K�ݭ�A�&<�#��(�:"*�65ME$h�gv1�n��h���,SF�6�M4�cm�V#PTD��m��IA���5��f��b'F)���;&
���*1�lZ�A:5i�F��kڶƳ;8�j�(j6sE3��k���U�s����Ѩ�������ES1QM3=�ة��k����3�|�ꣻ��+��*'[wjq�ŲF�*�j��t�8튠��,^q��j���GF���mQQD��F��v��Eb�c:ƝDDĕm��u��
k��ڠ譬V���tmbњ�N�(�V��;Ͽ�ۏ�[}z��V�d�͛2*D�])���ⷔ���"�����ݼ9�_�8&��(�ەR�o�����TS�6%�F��}�D6߻ٰ��7�-�#Q����$MU�$Oo=�TJ��<�`u����o+��>�Ƹn-lJ`m���V�3�c!�J�'�U=TFO`Ӗ��r�G�^95�P��d1��ک�?�=u�Z�T����O1�׍�f����m�cil-'H�%jK�u=�2���O�d���cj�6z(v�h�DN�q<Z6.;}�w�uy���$#)�pe���tƖfR��#L2�F,��gyWu3��)"q��*��I���N�쌬�s&.���?d��w�N�6�OKb�<d+�o���MH�;�V�g�t���8�?bs���ŉM�K�,2]u<u�w؛2� nT���a�jȋ�7��7�?B):��%j�h�S{2�S�U��f���D鶮:\2���õn�I*�u=�T:4T�X��U7�
���u���-x�N����]�(4�}�d)j���\��n����Rf5���C���PzL��k�g=�Q"^���pp��~�M�p��r���@��WU-���N��e�veq�]�ow�J��N��7�I�n��0G*�*yM�7�!ɿ>��,�Κ�:���Y���^�G��ߜ��{����R�!�4�j]~g<���)�[u�/�{V�Z�3b���B�El:ޘp�p�Y��9"�@�����1�h�QX��,���12�l�t�73NXh���Q7��8���pا1:�����e�����Eh���<�N�|5)�w*ͻ�����c:#�a��]�@LlRF��aVV�Y�խ2A��>�I�	?,e��Z�6n�0p�8C���D4I��~�	�~��Jd�r���Yg[����ܞǞ�h��w��T��x��W��#�w/:��BθW����ز������m�a�`,g�r����)���{��
5 V�6fn�ں[{_��i��ZW��iUg;���Ʃ���N��Hq��V\�[�{�;N6�fT2,s���g��x�嶼��{�//��c\�&�q7�w0Mӭ�z5��%^�.�s��(^.�G����Wq�Fۃ��'�}ʦ
�r+�3�� VK�w�@I6��>5���c��sY�$(��A�ݟ��"3I
dw>i�_����>��ofG��T�O��j귥�Yf�ү���΢�.F�L��SWR�0�o�陌]x��t��:��4#څ �6����;����K�rN[H�$mt�J���]��<d�v�댩F��T�5��M�Ku�y�rG�h�HJ.B�u<�� �k2��K�d��}[��~�j���϶�%�7*�+����Kj���6�K�a����-7D�kCx���׎�%e�R�kҗWY+Z�Va�)�,pw`�nݼ;�L��6TIۣ���� F�ř��ѳQ}/9x�v�M�TA��q�ʻ[ q��;�3-��69����>"�NO==��9R��y�=`1��ij����Q�]����F���$�{w�'"��)���޽^�,�o:}�'��)j���p��r�!��YA�����z��ε�n$�͆��"�M�����I��7	o���ܵcSf�6����ͼu��0]��~4Z�G�Q��[����"�Qe��K�u�I�]�y!�V�J��1�# 1e��[ܙ�Е-�η��Q}à#e�𭏮58i�K�8,���:��\��E��}�W3����h�R�Ms�l��v���寓5�goU�d�E��Ow��1��	��h�\����%�kxv݅�:����'���t2AϙU�)�{��̨ x#ۏ��G,Jv��q_݆�\��y�WǊ��v�u�\]����!K��s:29����������suX}ǲڻVH�FC�F�8�����	H69h|��������`��S�T���[�Ќ�e0�����YqWd@~q��e��%��ל�t�I9B0dzn�(o&�H��$f�G�9.�����+��đLˈ6Iz�*	�J��}��ܗ�&�\2t��]��׼T�ǆ�<���a�^܉��.��H{U1��t��B���K���ֳss�i�������ov�/Bi�r� ?KT���5�"h>\�zM7oY��=�oK����efҺ��u"���Y>�IM�A>n��7:��Ύ%��wK�3���{	H�1V�Ww<��}+Y�T�I��Ⱥ1L6�L�y爫����1�d�}�U�2fv]\n�m+3XhgkJ�6�^N��Z��)�B������Jm�X�+vqCh�C�ѽy�Xĳ��jT�WR�h�+m�n�`H�W[���؋��k\������l��E���Ө]3�	y[fnO��gw���J�:>���a�2wl�����\sɠ���Uvl�e�f��q���R�Wh��%�QE��Ź�j���v�c�z�z٨Y՞�8��}����ʖ��4=ҵw�$O)�0AYs��n��ݜ��.a������j�x��V�sv)��Fp�G����5G\S�y���B�t�Ս��+
=�B[xf��m�Cz|���
������ͫ�;�ȸl�G��,y�#�.��GQ�{����qa�r#�n�,�.b��ފ�"�F\�H}ҫ��I%��W�Hn�����(�â���h:�zxd��ف֤X���?a�l���� %h�Ӌ����wӹ��-���o�n��-J�#f���֐4����[�(	��'�Gs&o��Gn%���>H��Z�L�,�v]ܸ���Y�?�R��h%JkeI�Rڗ���R���㧂�䜞�ۖ�����a{���;��H�Z���#�@��_�F(�+l������R�g>Npnuuq����h�B�Wdko���˖�w��S��ho%bf�T"�>��o^B��B�*�s�`2.�ɚ~t*o�V�	�����$oz[�[��d�rk˱�֩�6Z����R�&�GlƯ6ɚ�ǉ�!�2���� ��oyޥ����K2�b�x�����m�6e�s!���FI�~��/>�r7\Wa���7�R���n��#[�7�ZDF�7��-|e�@�V�pq\z[R����T��%Xe����C�����ʇ�N�Ȗx�:�T�8����1�*�	|���ט�Ƣ�ʇ��sG����||��] �w�\�bn]��2�pؼmB׮9�eUVM�\��2�&����Y�����#�=A�����#�Ρ:F"8=Z�3u�A��I5�G;E1��δ�9����6��&֭���@��V�_���ʶ��x�{��ٹF2�D�*��Ǫ7z�rW"�6��O\�p�M�xz��YL�������;u���K:^K�w�E��De�w,U�����5�=Oݞo/��`=�2R�c����'.�k(��YG8��%'{d�6|���P��z@�\hl��f���� Ef�J[g���H�Sԁ/q��9һ@jnP}��L��ZvGDHZ��	�ݵ�Y�W�SC+��u􋓛�_w{X5׵�X��k�f�<��������82���Y ���*���Xd]�x�{�����q6�����/&�{�s�4H��~��p�z!�9^��=ٝk[��:�
hl����۷wUx�X��FG?�B�F���8�����Y9Mg���s:k;�,�B�⌼�҄���B��V쌲�;�{%��n����&�ݓ�_z��-SzEu�=;W�'I��\�����)0�3����eM��΢��+^i��G�f|�*�R���%e�
�R��J�(%��^����tu���,��S���i\��ހ�
���m�p��Ӕ�	ű��Uxԋ:�]pު��T"Ol�q���
j�S�:��'���A׋;yٻ;�e��f�#r��5��z���vq�!�f� ��\��jX�mz'��4����	����z�)=0u%�/�N$:���kr���C��2��5�������qp���.�
hGf�Tg�|]7r�r��t���:�*����&��!�ݒ����fJ����M�X+,zS��G��R��)�6� Z嗽(kl��MZ��l��Q$��o;Z����bdwwa�l�fߑ���\���q�8�=�	�D;��찛���1[0D�ɑ�TѶT��\l1��`�	��!y����j_|VۿX/;|�uy?d���eU{���W��TTJ�t�%����W"���]��M,�lz_t�4Hf�!j�Dc��t�"��Z� ����p�-�����3s0��L�ڱ�;o��ڍd��G{En��s�:����ŭ>+_%L����ia���h1@u_$��U��E����D��pw��va�;�̆2�0����e�8�{rA�0��n^i�[!.���{E��L�^���_�
:/0�{�^n�����Kё��EZ�"o�����Cg�[�!q�BU^i��<4uu<�4{X�Wz�rSŎ�z�D�]]�1C����#'J�7�"�<=3ɸ�|��f�4	5�9k;B�j�ߕ�ý֓k������gt[8��gRQ�W1�qkU}X�T*\mfi�N����j��r��
�.R��)w�K�Az.Nj��Jg$%\m��&^���'���n.��;jt�X�r9(ZÂ�|}�o�k�u��מ�fߢ*&�Y�5�	��g!\ʹ����;��c��wTaأn
�sl�L����㷥c�S�3'��[�[7=v�[1�.�"�h�H��+hW�UMٷR/t�����Sc�ׇ�ٸʓ���O�q(�GI�s���b�WUc�=ձ��[;��N�Z�ЫCg�A-���j}ܫ�y7$x1��ή�KyW^Ty0w3����Zg0�p�3�="rR�,Ӽ��4�Xd�M�؎z�ٰ������Fd��O��:13��P�[��z���D�ұv�ɋF������M�=u7r^�m�X%M�׈ۄ����l;������v]�Em=���{�w���r�%�G�g�08Ņk$�3dL#������L�l�U�^�Uo%�~(�H
��wFN�ؽ�ְF:<b�B	;��&L�e�'#�F�n�?�M#��C�S�rN9�t��J��Z��j�u��m�"ݢ2��L��Bc��ӧJ��d���r�K��k�F���*2�*%��V��>�&�,@R��=eU��=��ܸ-Er�N�n+0��:>��ٽ�!_��FFMǶ;%�m���y�@�0y�ǽ7�m��R���f�u!aF����ڐ,Y3۱��x��=b|��~�0��rO]}y*�����ra�����}�:�]D�s�1�Y���?j�Y�z�d鞌ʡb�t����v�Լ��0���7B���^�r��ъ͈y��$��D��Hl�i��u>�l213Er~�Uzf�#5Q�z�W�=yz<L�o�)my��ِ-S�l�{�nU�G[=�Ӊ�(b�ޭ�kȨ�;��o ���R��ԕ�Ѷ�1<-���l�$�ff��!�l�苑��,2c��Ko�<�Ȩ�Z��#on���R�������1o1����"��*(g��R��u%+56�K�Տ$��z��7Gk�u=�+���5y�,��{���t��q���{���O����{=�����5�[$��.���x�a�3���P�) �Z�<Гݬ9N��v��Q-�ef1,}�B�LͬV����lkTm>ŀ��zS�6�Q�3RT.�k�n��.���E�[.U��ݭn������ݥt���puu�ux�r����z�'d�e B��0�]\�h7V.^��lac�é��77�ܱ���/K|��C��a��KءZǉ���2Mk:��.���C�^�&H�xy;�ɢ�-e�*�����y�W
L�f܃v,<a��s/z�MgOފ\رëG2gcCCov�=y�����,�\���$ֺ'*N�dF��f�6�OW@���3�1v[k^{+%�f+OU�����V�v��CiU��"B�S6���(	p)X�ۡ��ރ�D­3��gki�sL�j�=���v3دA�r��&gd�W�Q�;��w�5}$͇l�s��46��rK�� �i]��/)�.;t���
�:�3(D1�OIYM�����Kr`��_x0�-�C�dWQ�W��y�x��X��]9�tr��2���nӐi�K������0biR*ջ���u�vp�vV�$�Q��Sj�TD�@D2Am5ub]'Z�;F�m������6�^X6tI��vҷ��+�J�*��Xu�3�X�;ƀ�o����hGC�к���>�i�S��h�ƕ��m����-��r�:��T����X�S�~/o2�2Xځ�I`�N�f
�Nℭ�ky�.�0������[Hme���63��7�b�ǕoV�gfuu��¶�T�3��	�Q��څ���
�����fT	�W�jΗ�"U�d����]��A!�K1%�5>}VkU�8�НW������Ϥ�rS�7�{��`kE�y�Dn�V��lڍ_cr+�K���qJFi�mv�ە*vT��X:wKC:9 Ν��(��Hs��+��*ǺI�����VR:�4H����3/��s�o^f�%*�S�(3�r�Iy�Ȟ�L���e�a����� ��mor�ynW{�r�8q�1[�q��N]�9Ӑuj��2�Ǳ��E\�ܤ�p� ��8ř���Wb�*�ة�ksx��ԧp��E�z)#���u�׽E�5�VBhO����*aR��q�y��a9w�2Q!�Ӗ:�k����Nf�
����j�������#����Պᵙ9�>Ý�2;k@*��*Ðe�ُ�����;Ugyb�Z��<���n�������[�tk��Gj�����G*���+z�b����uw��N�'��R���@�*���n����lJ5�L \�]5Nf��1��-�����56\��FK�\|��7$P\@�9�]��&nPx�R��ݡ�$�ϝ�X�EL�in�{�D!��J��X*���j:YI���%�4皙�6�퉌�]D�����
v�p����F��l!D��I�n�C�I�*���ԑ ���(�(���uIQ$�Ό���[���=����6�wsƳ��m�ES[`Ѯ�b���ǘ�GOڨ"-w�j���[j" �N�����F-�F��m��.9�pST��6q��UQTM�T5E��4<��e��*��n�wi�V��&��j�k�k���0Eu��h��b��3�=�ż�]��F#K�4���y��቉��6�3��Zb4��ъ����[m���To8���k��d�kcQ�vv�� �Z���լ�G�w��Q�j4h�h17f�u:��E�:ŭV�]�ۋ�%i�5X�h�w]m�6��J�
LJ���)b.1��A��E�F�G�MN6<��h�j(�����	�4ղ�GG1��<:��cHPklh�m�Y�J�G�||��((�N�u�b�)8s���������K�}�Rg��+�kd�� 6�`ɢ̺QLٱ)y؈֫�Dnh�y��	%�`P�DQ6�H�U�-І�F��f�_��J��6�:�5ǎ�u��"�9X����^�U������#.W.��y�2x��-�a��lٖ7�L5,&����f��W%�Ϫ�/t��g�\���s��N���F&�ms⣧�J�6�ؕ�kAz�ٽw����]�WGw�h�gd�L%�i��Ta_Io�s��;��ˌ�ٛ�cK{y�eo��u�����xjCr#����M�&�{�@8��@�@�b��:wR�/��S�PO�}Jγ���T̥h�2���b��ű�t)x�K��v�ށB�ռ�ڬƸ��S_oÆd�ζڻk��R�^�O��d�wH�a���F%�k_t���f������oc�� �:B�Jݡe#�(s���3[cD�]c�4qއ�Ffȉ��H�Q��'�x��'�[N�ܭ�G���F^�c¨��:U�'��5O��1���,$X�МoJ�٧"�l���ms��W��;�w�2E/��{Y������[����Cm^,mΓtD�gAq�uҶ�uenv���v�M��nr�e��fY��
s姨d��6��R�sT�f�
G3B�j����Z���{��uG�WV�YU8,�D�ʮ���{��3�4��.��pT7CL�r�*��=º�^A�Uvf�%�n����n���@�'2k�U���u ��-s�	�qg��K]��n�.�SY�C9�$��5r(��Wq�v�6dy�k�-5�uS6��e<�_2���"��kBZ��0Fu�ާa["��Eiic��]��^L�>
�������gz�b��G�;i��Fq��c\�F��h�W���$N�&aq���J����4�%�z߻&L�g��F���1���-�$�D/`� ��H��]����.b��SU;�yz�+?62~���6p�m��އ��;}�?j;�����ĩ����V�ǝ���8��s��������0`�ƇJ�t�<�a,�kJSe+��V�1қ��m����G��γ�oPR>�.�b��:_{�ыT�ժW�١��C7YT�����:v�����2.F��e;![]	���1ؾ�y4�hڵ3�+�/��ԛ;�Ib8�@7Å.we#ȓCW���h��7s��)�1�7,�nZ{��A�,d1�ba�d2O�l@���!��%���7�τ�X���]�[�e�u�>�R���Ns�v��҈�&��Yod4S��(�՘2b��-��R^5BT.9{�P˜K��2�ޯ|3]QZ��{Jbk�揻F�<N�Ȍk�pi�^��Q���֚t��T��|i����S�1U�>�ɗ��Ii�zX'�a�����EX�$��53��ڪ��g�-��@����|�j7%��[�u:���I�Q�ujԥB��wUf�M�.����[�jZ�l�W���n��B�i�?B��]���|u_\���lH�i:E�M��<�nZ��}z��m��پw���$g��T�=+v�%t�9��ˮ��i������;6;o��]�k��!\Y�n�K�TYJ�����Q��j͗(���.���	�+r�u�:�~&�H� �x��]�j{8=�W��[ʳ�=.�ٗP�餵��8�ӠD�k���.�@��]�ThH�Z��uiCV��M����jK]v4�kzAǎ6�4^�7�^��wd[���*�ǟ�3��D�D���4��0��֍��gi��i��;��bw1!丕~u�8�����(7�^;+d��<�~�%Qو��%�2�t��n�{�zۏ��Ye�%�xf�|��pz��v�U;\��W6������ê�mex�k�m�t��k��a�Լ�ہR����8Q��:�l�s��}>*6H�h��;�y���ڦ.�tNg.+��\�O]1����H��}�V������������;e��z-Wڜ&�ۅ���[;���\��q��ךs��9;o/cB���7S9�Z04��4@j̞1�y�c��Z��R"l�\t���w��]��"܌��c��H�Bl-�h�N����g�~��U{���H��.s���I֏2
�v)�A\�)m%s�����EM9p��eϻ���g%��>�������Z�je�`���βmЭ�5t�4eL8�\ �S麱*�x�`ý����D���=���>9\d�K����JMY�p�����l'FI���<Xltɣ�pYפ48�Յ��������H������ξ���ly��f������1�R������
�o �
P�<s<�ܙ�+w���AN��J�7���k&��z�x�ty�BT��}�=ЖqR�����U��Xb����Ll2S��x����	��E\���G}��us��jf�c�4����7�d�κ��q#�܇{��z
f#�}l&�z���ў�I�lEum�ǌ��%���6��!%}Bs-����`�{��l�vDԕu��=W$��{��q\�y�٠ݙ�_�|�ag {����j�y.���r�ԗ}�M{o��m���R�VC�
�Z�f�w|��D�Vf�=�p�4� ��[�{�ﭹ�}�es��SL3�4��U|���Z�����;���,�I��Q�S�g2��ӳ�ܲ��fZ��M�U�vec�e
�*{�1���pǺc�@e���u��k��j�h�[�\TG^Tfy"[����j�w;\�Nt�rȠ)����(�3Z�D\uw�Ln$l�b1L�p����3�$���[A�D�ņo�h]d�Z�*[�$��CI�1C��B.1��u8�X ����a�"�r�<�SYssST����O^�p�R:�Фt�юgo<���D��eue�j��j�N�-ˍ,@*��qP��ߟ�~�<�����I]���<��\��*��fK��)�"2t�r�h�G� ���0,�UOyB��b)�/���Q�s1Jɿ'��_��S��t�ԗ2���W��L���C'B�����g��i�zڸ��R�ĕ� Q�d�6^Ub�3'w,��<"o��.�q���ݔ$C��3��-o6t+T���ΐ�j������ê(���i����� oJ`"O[���eo�����j+��X3�|��g4�4��bN��Y~����4�G,ȓ�Rِ���ɠ�
�0J������a0O��'x�t��Y��򮼔�|�����t6�������v�}��м�#%����2U�f�'�7�q%�?n�H�k��u
���ʶ���������g4�8���a����׼�ouÑ��o�`h��Tʠ������b���Q��~�3����+��
�1�*<��wi�6�G[t�1�nc���w{��ݒ�s'e�q�Qh͚�:q�2�c��,j�ؼ���{���j9B�Z���g{�I��?5!�)�=0x���SݺL�%�-�i�-�g������Ϸ�U�1��il��0;_�6�v��zR7���7e��Hu7;�lc��-��鼜�X �g�W�ax�s�#p���f�1���/ss�E�Uǉ8p�V�^ϔ����0���b{c��#��
,�Գ�T�wc�j�8ݚq{0\f^����-�u�R��(�Rl�3�c5�L��w�� �ז��n��ZA6#ți�m�*�	F�������7kH�s��&�W�6]�z������(U��s&G8Y-����)uP�h�e�,[�#���h���VEV�q��듯�s�K6�u� ĸ��A*r��zf\�1U!�L�0�"'H�	�I2V����y�UN�<G<�^[I\�2��[Ls�1�CU+�\�u����}g���%�Վ��?����r�����z�or,�B@F�	���=�i�Zn�9�T8V�Je���":���ȇ����������M�����.f�{Gh��K=���v�P��:ux^s���r}�T�*-J����nqQ��ިUk����j�R\u8��Uh�o�xa�S����l'���S:��tI�>.����u�3��]�JD�*�
��r��惾o>S�+���}6����BM��Iy���TEo<�1�k��ݱ���G"�|P7ɯ��;j�cv�[�b��;Cg�9�mKn����*�a��Ʃ���Ux�ULkCdfN���y��o�t��K��ong��&�k��\6�i��gj&�g�3p��J�"Q���S��g�fe��Y���b̭�9���!N1��jN��;|������ݕ~(�!-��:>�b�_�'���|�?�u�<�+�������w�1�5Wrť�ul�t��,�G�l���s�Ʃ�yx�v��B�����Lg2R��������_��N�E�s�ed𬽲�\�3\�sY]���ȱ}��9�Xc��<��je�ބ���b�F�iR�V���1z�p��]��z�_@4	뜮�uzE��Y6E)k�p;�$�G'ę�w�і��4���]�K��*T���-�w�����[ʜs&��5>\���颇V���رvkIk�,+ u9|B3�V�㚁*qp�qh.� hhՌ|z��v�b�J$}�;�.�d��YCu.�Q��L�Uݖ�{E�x8�(�{[��j��6�ǌ�
M&�T�z`3���EdM��לO��U���f�l�&_1Cy	���i��aǌ�S��]�����our@�ՙ�&���֠���b���mi߽*��-����]���w��g�n�:���P.0����Pn�6�+���(4�k�7�U}���e����UA�\��5��׆�x�BYA)Ici�b����׋C��^嘵r�����wS�[(�Z���amgֺ�.k�j���u����'�(��S������l��=W��S@~f�`�t�w# �M2_���3B�)a5�X2�9�:�miP� �}B	s#�����gv�|��QK�7D�uK	@�K�e��Cϖn��c\f��}��;M�P��z�^��~��,&�K���ˣY�h]^����lg#u��{��=��U#�Ȩ���=4�gc1	M�<Gi�ɖ����K��oPY�VA1Sq���a�qyc�H�?�B��v��wN��h!-B(�ꮦv��7���$��h��ܞ�� C�Ǫc`m���s�C�u)n��'�56	P�ረs�<g�C&4�j�rw԰L�>�U7rYg[�Ҩj)�����k�>H�y��,o<��G4�`Fٟ\�w��\-��c�ڹ骆����mi��������&���an˺}��X{1+z�q.%��90OQ ��Ùۃ#uƍl�� alkSG��A���Y2os�zqOB�ԂPs#ݧi���H�R��R6>[u�WA=zr��g*ƍw"Q���4NǄ���2^}�ŧ��4�r��#,���vX�N��Z�{���Ց�w�J�9���|���O)�Qo�&�������/Q�U;���a��cR��W3�2.*1%��%G�� ]����u'��u�:ɸ� ���m߶��n�{�j�L��@���@��y�>>�/W������y��p���j`���Ȳk�h�U���6LklN�uK+Z�/��E�wm-n<o�F�i@�"��潑Xg��J�ʻ�]rb�l.Qņ��q�Z��@�q�{ЪYX���H����]t� n�	Pf�<s�X�a��5K�U�p�H5�����X�r��%�(csP��u$[e6�O�\ۀ�j�V*K& ��sZ��f��*sَ
�[�u�Wh-F����Y�rW��	W�Uҧy�IE�����QR�$mr�{��ƚa��W���Z�#q�y�kj''����]I\ay�_nV�)���u���*�
����ұѯڬw���(]$~}B�F�k�{��E��}PR;�u�Gt�Kj�q�Ѫ���m�N`Y�q�K��Y���w]Ci��Dd�x�>9X��S���1��n�1Ҥm	]M��p�C+�ӵ�i�����3e�u�`�4]JTv��{��6�]A�������H��zJ�u�/���ax7v3|oXЂ�����@�V����Fc�oR{�VdI]v�{EX]%bzrF��5���kz�d�i`ݚMr�k.y�peE���]z1��*=%t��5�u����7&޽�u��D�\�l9hF�VRR�w;*�͛v�g'���t1���mp�mE��K�������"���g�'}F�eG6�Ϋ���[����f�����_�~i�q���1����AgC�t��������D�Y�)bx%�r�����R�*��%�S��+���N䚫���|�*kn������H�/+jvu^J�)U���\ׅ���aI�C�Nt�a�ʡucr�۾�k��+p��&������3��t��V�9{�=1A��E��)Y�eL�gk#u�T�;w �}5S0m66�ɛ��S=D`�jRbU�����-S��xWt���B�+e�v�Y��AI�[+��n���`'\�j� ��S�^�]5����t\���ĀYn���nK�f�ԝ�3r̷�}é��_-�tp�F�ů7���Ÿ9ʺ!�$���ӗY�t�5��OA��j��}f��9{Ƶ�fɈ>��� ��V��ɀ�}*K������Y��t��^b��j'B��J���s��=�!�8f��s`��e�%]��м.�caw����S	��[�+2��z�@4I6	��p��c;3�u�"A��I��/)��Q	�.��]ַod�6B���cV՛i��͝�X�ҏiz�G��g7t�9Wk`��-{sl�d���l�Ү�U�p�Uhİ�9�9��y/^�䆅����[{f;�:�o2� ��ȩ��[c7m��Cͦ.L���U����MN�
5ͨ�����8�z�u��gK�HSJ���*4����Σ�+l*�m�m+4�\�s�&��b�7bT\M+�}��6r��bci���G��f.��4Vܫ[��f�rР�6�m�iw��F�cˮ���k`�G^s���k:�J=�J�j��km4ѵ�Y؞�GDL[j|��u�]kWX���F�g���Ej�cG7F�Eu��]h�uV��LIڊ���7n�"��cAAF��T�v붍�S�i���vi��*��&�b���`�cF�b���e�����v�;iֈ�mӘ():+D[`���1kEk�:4�5�1j�Cثlm�`�*�ͺZ���T��F$���8��;:�1SME�mN��ED3Ph�MSQ;Q��&���v�l*4V$�F�Lm�"+�:zj��[b ���h��Q�Dm�Z4Q���>cZ�5�1�gml�sQV�4k���U8�gT�D�P�n�'���NccE媪j������Z�l��b�Z�J��tM�<�QRyv�Wᗚq��>U��%�䨣>�(9j�'�<�,�'t�<����Y0c�;����5$�j���+�J��,�ͧpB�q�v�M���?���J���x�`�436��4d�U�i�J���[�luֈ�irb��]O$e�#�K���ȣkhr�ûً^�)	�Si�k�����j9�����ZF�]��"��x�]yQԠ�ձ5�g�]�{'C���=@};"�"�T�S@��U�Ƈ��U����8VcMV��9rp'|�%��.�Xzs��n?�t{6FF�ZUC���(�M�{#)��yO���ꔗi�з�h����(�v��f�؞]���O�f�bn��v��+E2���E6���>{|WX��^hdEAn4[9�e�5��	��"�}�N�T|������+�=z�R���������'�#��z� V!��P�;��z�:�����"b�[�jj,��Um<M��W�#HhO1k��P�d�����H�b���5��YVV������q�5ε�\FӖ($5i�キ�<�(��;��f+M���s�+7$����.񾙛{B�1�xǴlo\�O���M$r���qwc��p�ۏ
ݲL� K䳯{�l�X� �9�A�ܰJ�:���p^����A��7#�J�-*�6)�#a�<A�"&�V��/�[HH��n�[�+];W�F22�@�I����U�t��gȯK͸�h��i���SY���;o��0�Q�[��O �Y��!��oѮb��v~ﯮ�����f}�.p��[-|BsՈ������g�:[a��7.�M;��s',;;�޽��������9Z�V�f�����]�x=�u[��E��1�u������ڔ���K�&�?�V�{�5κ�ĥ��Vʻ�m��Q�淪�FwH֜� ʥ�96_���.��H�䍆tQ�gCku�f�v�g۲#8��p�ҩ�9��/Y�Ǹ��M��X]�vV�i�����"\�K!�k)�����9���彫�9�d�=,��dƭ���a�&;7,²X��r;���Z�u-��ok����!� V�����أ��U�֫����R�2���Km��7��r�&޺��*��Ώ���K�6zm���>�Y�o�+�����g.�j�!f*w�n<�A��h꽌V�Y��S�b��\iΘ��u�r
�s-�6�}�I�oA�ڽ�cWz�V�f��h?�z��!��(�;��]e��]�6~���[ �5H���9��(��������5�VN��ٻ�wN_��
�B ��P�wP�8��	�{�+i����Y���,�=ٱ
go�plk�]�cG��6��X�Y#_V�c﹮�1Oz߽ӳy���;�#7��!�u6��p�}�"�b�����=t�=�[�2�A�%������U�	�<�fC��%�2�X�����D���t��k&�q�m���B4�yUz;n3��E1���Ի���똈y���w1'm�Ϻ!��[��	�1�X��$t���k�8�!��auH���Jf����R�	v-��B����nP���5���y��:a�_��[M5�Ւ��߇gJ��J�h�Zd�LLj�3��6�9٪.!��&��܊`5TUm��S�֙��a��T��x�T��1x��uvn�R$vJ�������5�yA����(�����˾
��n���T�Z�A�rT�fd���غPp��e�D��y�,���z��e*Ƶ݌��c[Y���G�jA\4{��eo���dK�Q��-f*j�<��Q��MBz���o��?j�v�����!�0�D�9-���<��F��su;�X�\ws>�@XR޴�f���]ā��|T�[ż�u4�~L{Z�\U�+���V��h���5θ�c&Օ�)+�E̳�e@�"�T��;�z-�0�5o�]H	��R��K,�ݗ�⳨fU�hض�Qm�&��<���^��g?�7^W�0��ا�:7��uIw,�::�Hl�0��m�����1Fs��a�˳f#R���|�um'^����6��k�p�F^X{Oh;<E4�n�����u�*Ɲ��la�S	��4�U�VXs�}g���P&�t�}����F#0�|ȱb���i��{�3d��1@�=�߳Q��Z'�����g0���&鋊C����v��X���|{�d�.��M|�zq���%,i�e���t"M�J{p��[R�����b�7�:�����ط+q����;�0зh�ۊ���mc�w�%_��"e�ZN�;@�Iz6���g�9��3kyn�η
˒��(�y�k��"�Mo����?:���z,�lq�:��\�]j�#L<Vu�z�!�x�Z*��P=07�s�{Qr�u�L9;�]����͇�/�� 5*��g�7F��-)�Bҳ�gj�9O&�ſ{���&���wS���K%��7�������]�J-B�~�n�F�33rL\h�Lu�++mdB�g�L����5�ҹt]?̴<�	��=<�w[���7���;@YU��eO���'�K5�rЦ{)MH�ӓ��6���=�>�h1���G��a5�io+�9� �>����V��w]�=S'�����7R��l�f�Z��;@�׸2`���գ֛P�^O�C��.��t,|�k�9�x��'{��}d��y�5��*�*����Dy�r|ݝ"���7 l�FV�6>�`�f�*�ڨj�
�v������$�ab<�6a��2'�|��������a����1{��%}��v�z���):Θm[��������lZ�o(���>����������|Q�Q}��R���H�:�^O��փ�EQ��V��x�m9|x,����P�[x��jx�[��槧����{O�{��˥���KաϜJ�J#ߦ~=�u�t�'n���F̘Q���3�F�ՀX��(,��S;<m�}���킺�mx��q�}xp�s���a��ۏ8���L���&��8�Ӕ ِ�C��2��ޱV!�n-c����mO��q��31�#��ZI�՗7�u�Z6os�up��5�����7��<��u��:+<�K�$��W������3}���D�i��{{�Pޑ]��u6�f<����Uug�t�s�y󺯻p��2IǮ"��8���<t5�� ���J!hj�bZ��N�@��F���8��ﺣ՜9��MM�qU-�~��m��%����;ͽcw�':H�H2�"������� 6��)P�y>J�ͺ�d�|���]����MN�y{g�b�Y�Гe�b�i��{�v_�H��*�g�ӊ��u�h�ՙ�Lr�y=��o6�=�Ǯ���:c���E�6��e7+M<���:�l�8U�h�Gq���J_�xB3Y�KD �/�f����� ��0�LLE��}2�N�\i8-Z��Ζ�a&����;M����^�����W����QS����M���Y���4$��"��3{rJF�n�޼����Ê��%nY{ųܑ,�ss�C�(���=����F�9s�������K��j�k��s�(4����a�k�ɬR��V���fc"�$��mbݟ"m:�l������o�,Վ�*ʖ��æ&L�]I9���e�8ꤳ��˺V��6��C�g���3q.�l쬥�,t匿Ҍm���ǥ[۫,�,$j�>Y�l-�meA2��Y�v2�`�
���K.�B�����k(�k�+i�ӑu��z	��:L^�3u����ȅш�Sl�M�)���>X;*�v���.�����c:Sմ��þԱ��4�6�;9�m�;R�2 +3b�=��j:L�Ϊ�jΪ�0�Oy��4!�^�X�}ˬIV�H}f����ȼB�",�Q���#�Y�m�i��[w����#K����g�����FGoV�v"�pg� Z�9�����?V�i�މ7�$,-heկ,*̺G���+�B��ʊ�F;Y0��	؆	���[p3�&�{�
��uۼ�BUř"��z.]��7����
��z�j�4��4����*��;6��2<ĬQ�2�Ѓ.u�[]�Ƿ{��_e��w/#1%�#����G��C��uOT=���8��l�v�c�Z|Zf=���P���R�y��Q�*�(oQ��xM{v��F�rt#6��s5�֨�W$��6B����A���@:c�'�C��ζl���۷�m��J��P���5�N)a��mԡ.�dLֹՃ[�r�'v��u3s�7j�	�����M���u��f�m�ji2�n��C���1��ypR޴����`�c@��]�H��S��(�ﾐ�t��S�M��\��&�
]ҕ��u!����#	�dM����'��ێP�?l��i�zq7N�(~+�Y�[/{m�ۤ���ZOM����Z�<;�}Sw�	��^�����r]֖VB��l.�o���o7y���.f9��ƹ��#��-�vk�{`��#3��{d�F��db��!fXR ��w���e�xx4�l�Sjoq�����Րi�W��k��4�k�����zU�r�Ｕ��%�9�L��Z����v��/tl�29��mT�V4l���ٽc�{��
Ư�R�c��C/\�g���Xo���'L{��yL�\)�wO8�IOS�t�-}���m�1F|�ìײ�k�����r�Wwy��ZOd��z�M���d1�����b&s��8d�-1�7z>�����IiŸ��oH-Bt���q���,5�T6 l�OM�e}�5���b��+E�1��>Ӎ���Ɖ �R^�v�᠚��f&Ymm,Rr_!Ճ4s���0l��h΋=�-瑺H����b�Cz�m���ᘭ��b~������Gt�}j�w��䣶��貤�q��.//1tp٩�k@&2w�Ԏ6����5�1�S�r�t]�%�^gOMV`"�����9P�N3֡)j�vS�����=��`v�g�wh��v��t"vzV�TΕz����,��	fU��e��d)�34�ӆ4XNv޼~i>����2�"Au����Y�4���� �:��2�iA�k�c��U_`�Ѧ$���u��ͽu�8�a,(�,u�<�﯊X�i.�A���H�/"n�l���L�>��^_'�k��� RWdt�H�[��[�t��V�0����H�ǕV\R�1\�z�5�iX���Z�m�1e9����c��2�p�a"/�]̗.d��[�x��Ϭ͛F�x��,����q�8�S�kE�.�k�\\��ZIt��cw��E����|���p��t�W�dv�����t��iU,���&T;��z��j�뤙&Fm�d��&=�+�	�[��x���p6�f�մ���������Zܕf^���sYY�+����Ղ!S�?�_EFY�3��������OZ^��Yϒ��m�x%�ʉE}__��c#�4Wp�ɢ�q�85�)$�v�&���4�se�ג��2@�53?'uT7�0�V�g�o��<�7t�J�ZwN6�^�5��i�[w��3n�#�ϻ׋�'~��h�b5�-���L�:���S3�@�Ԯ�yO�x۹�UU��$f�d��cB�ֿ�@��^���<\�?��?������߹���<< w�B
�/�߻����_��]��q�<3�v�(��"�*��*��*�"̀HB�*�00,�(C(C(C (C*��"D(�UXa d ` ~{�| �� �� 0� ��-��@��a�T � C C" C( C�� � ��ʠȠʠʠ� 22�0"0 �2�2�07�*�eUa�  e aUa�U�@ �  � �ES�2��ʪ�*�  C  C C  C*�  �� ��2�0,2,2�0,0�2,ȳ
��Ȱʰ��ʰ�����0,2�2�>C�a�a�a�a�a�eXe`X`��s�|}����?8Q&Q�|@��o��W����������s����0?�����/�?�m�_��������h �������E�ݐ@X����������'���4�`�_؇�( ��?�?_���$�?��O����a>������o�� ��"�$( 4�H " A  I*�@�  D*�B�� 0 �   K*�!
 H��� ��� @�  H�?� p�� ��c�xb���������*�-*�@�!B ��?@o�?���������<��}���@^�������;�O��?�3����?�����W�?$?�?w�~i��@_ւ *�Z���UEw����B������`�_������������8 � U�?���_�A  �%���~�0�����ϳ����	?�����W����H ������'�o�1��`�'���G����|���}��'��� �
�	�L�������~ϴ��/��O�W�EE1���x
 ����?_���?�2��b��L���(��� � ���fO� Ċ�ǽ�IR��_M$�QH*KZ�R�(�Alb��̤�HD IQ�T"D�B�¨�%@����QR�Y	��**�ӗ5�Y���k����V�MRjb��Yl��Fm2mmYFfYP֭-�D�ʄi��5N�G"[5i���U�(Y�m�Ӫ��lX��j�VV�M6cT�ڙ����ٶ�ͥ����ڥ5��%�Qf�����B֬m�m��fi6ضm��f�6��SY��K+m��ee�������  N�vuе��������]�ݕt�m��Ηv·Zuۺn.��[��N���\-�dwZ�;J���pe8��EFKn�jt뭬���w[��u��tۣu�R���Zm��U�:��  �a�P    yF  �  �A�CB�
(Ύ�
:;�[^�]:�Z��u�k�Y�7.���aZ-�r����)4����]����u�T�!�R��Zf�­���J��  3y�zh��9��ݷv��˴�u��wC�����wZ��]:kX�3�N�m��fv�\���7r۹�Vk�hѦ�7U]V���S�A�nEUv�[j��E�j��մ��  w\�v�A�in�:ܵm��:��P�m�ڻ;Wv��
�ݹv�˝�m��u]�m�[4:�E�pm�ZմܝWZ!X�0 �]�v�@�m[[��5��m�l�USL���  �T��]�� 4�w8�S(��\4 �q�qN��EjLt-wuU[��]�c�tTW'V�֤vV%B�v��mZJ�����U�   ��Z֪�������9U�k4�6��Q�
h�5MMemF��n��!jӵ��unwu�]��S!�Z�8�N�@�F[6SZO   �ꧪ�5]��u�`5ں�m`:���dӤƺQl,E�UJwv��R�m;]\ ��s8m@:� Bhm��U1V�Ll��Y�   ;^  �N�@v��t Sv��  ��  :v��
 1[�  ] (h9�(  M� ������Slf6�K�  ��M 5z����5�  �  �àh ]K
 �n�8 ����  :3v� ������v��՛[0�h[m��Ŷ�   ڼCB���TVu�  ��r�4 .�p  X� �rb� �. 4H-�w: *�m��  +�O��*Pa2 S�0��� 2 S�<S�=@ �JR��  5ObJR�  $�D��T  jSdD�`C(�P��S��<��R�&2d
g��Ͽ]o��7�ӎg��߲y��IOٜ��2@���HBI	�BH�q	 BI�d$�	# ��BC���߿��?��ԟ�F�����5],qt���CϘ�1\�L���F�ҩGwE�˵�Q�O�ъ���6�����֣����!J�cj�n�6�P�Z0㣂m�P-�Vp9�Tݵ26\�x�!�<zY6�\�-�C��t�E�V��Xn�e�`�wd��Gf�%����@��oc-f]1y������le�'(�V��n��{��BC#�%��\��vmY1����@�B�;�����q=#�/��f�]�t2�	��z���*�u#��Z2�E�{���V���%����p���IJ�
aͬr��U����t�ZV�S%�S����
⧎�iЏ��`�׸ww��-�(%��[Y�fj��RV�[�R����l.$�^��ZU�����ol�A�wC[7"�jd�J`kC��EY������bp�5V=��r��2[� �`i1)�l^�)4��m���7ͬH3tM���T��D-�$�\�T�[��}oC�;�K*Tx=���v�+D�
�L*#�fLj�b�fm�w-�Y�5+wN7�\K*dp�ڑv��P������{&�B[�W���[J��,�I'�wsbJ)Ld:D�+�on�j����0�ZB8lEVԡp7�[6���ֹ���lP�aF��1���*����V��T�M�Y�!yt1*�ۣy&*2d�9�U�!�����mn�}+U��`�F���Fq���n���s+r�רԣ@1�ٗ��
�[��ޓ���*�o]��vż�41��k����teCkE�i8a�����4�����Q��T��-9b9Bl ���F��ۍ��(���ŚA3eE��`�j�<$(8�WV�p' ��f�PKN݀4�Uӽ����4ͩ��kf(t���2���SwK�y�5�$�n
��l1tb��X��z�r�x.��]����}����ڎ���먵{���M�[����j�����U�p8fM�q��n�J�j�YMA�;ūV�gmk`�,�u��,��0�����ur�
:��U�`]�M_,�rZ:Sw�����R㩮�fL)��K`3{krX�Pn'��Y)l�ױ ̓��0t]���4м��H�w��F��$)�Ъ5.]��8	оz�{����=���sf�x�F+s6 ��,0P�v���#�*`М��S)*o������ӸΠڠ0hm��h���s k+"�卭cd�rB60=�@�I��e؎�b����,0��p\5&ǘ1'4����-j3����mc��\h�u�Ƣ���%�U�l�[��bG�r����c���,�4,+^[e�Q���2n0� *�)ɹ��F�Wh6ߓ9���K���=̻f�����zn9)�`:vhc�I�a��Ӽ��c(�t��6�Ěk#ה���oN����f+7!�@ku��2ܺ�32Y�K�eɅnf ��@+�G̕y0���"h����J䔠 �M��U�.�?j�+�*����P�FW�(��l�F�N�C󵔴K�Ґ-���ګG����w}���Ш��ʻV�+Y�ʷ����$a�J-�lLY���,�2�\���;KP̽�j��V�B]E6���w+(�(�la��1den�
��[�T,l�֦�yf�%AZ�¬CfQ"`ݥ���gc0�L�ː�v!��Y�/�l��*�f�apAh�ȴu�`GeyG2)y�#W�٭a������t���Vk{N8����[{Zi�p*F��l<hh`J�^0Ujp�v~���$��n��H��
�k6�U24l�'M)�Kik�W�X��0��,,I�HD�ՑU����\Į�y��کci�����}�n�<�
Y�n�^���׀ �ee�7�����44��^ ��7KKŀ�ݡ�B+õ0�(��I���1P1�L��/�a�mm(!�AE.*j� ��(@o�Vp���sb֪�ukwvt���N�\;�GB�eD)����^�DB�	�(lYt%�t��w��W�̔0ԴҬ�+�6/�M�LM�����9����,T%:t(�L9� H͸U�ͽȶ������$��ݑ]��n󹾾�P�O�Yx��Op^�Zq��p�j�V4�Ca<8�ˣ�+Q ���K�kw>��x�&�y�J��F�$�W�\daP�As���t�G5�;n�[�I��vIS�h�-�6���:�c@ǣ�kɡ�X��UGo��8��[e)�r�RM��{z�#B�6H�
1:F�>�-��s]Et�$�@��ӛtb� ��I�s
ʟ,���6��5d�0��}))� �Ͳ��(jz����5��^�V��ͳk	����	Y��^S�M�q�i��#@���Fܰ�x�@f���轧�m4�E�a[S)f<IP�aY��QE�r�Vv֑uv��+6��jt�T!��F��gRn��*q]�48r��Qe�e�m�x�j�F3NL���bCe�1�ڻ�tt|�����"�`V�.��$����j���%B�d�	Q�Rl����v����R�V�2�ZQ��)���`%L�y��b�w+OR��M�r^a�_h$���`6̍4]I,�pJTK�r�dʎe�t�;���Yv�]B�*Ty��Xb��iR&�V����ݦj��Q�R X䪱�1� �5/����2�e�v�w[e�8���6AܽM��%٩JT�XKp���N�;V�%�cJc=�r�X����ouYYY%�KQA�5��u���m�Zn��LQ��ūp�7�4S��@v��$�&��lw�^2-����:�L��Z���f��22�;�[si�3�i
t��8�[EmV�#�h�Q�v��8q��-]�nOl�Kn�X4����:���I�;L��r�v����hљE�����[A0̬$YW�Z;�(	F���Z�;�`NSկbS��Oh0��L�{Y/a;�q�%Kd�5ֽTۥff�cLp��u�@Y��yKHJ�1�'�):�#�Q1b��m3k4h�A�Y������@V(M����m]LV��J+�O^�j�p���묥�Za�]^Lv�\�(�/t�WN��\���[:E��VP\ζZ�gp(>�o�7u�f����h1��H�FP���똥-��a-�m��]�ԛf�jb0	�\x���32V�V/8#Ya���i�ԣ j�*�B��ݢ�^c)B�ac+k(|j�%-�B�F1�L�69j�]�rս/Y���[�īR �z��d���ڀ hV^�m�v��"t��u�y�&Ѫ�Hn�E8��%2���t�\;���̓D�J��/u�%ܽ��mȊ�t�����S-��Q1�Be]5�R�`]Kzd�)M�t��P'*Q	-���*����{����s̭yP�mi0<��	GH����O�3x`��FТYI�O h�hv�+u4�/�F��aZ�"j�-�����]���m
	��԰&�6L���ֶ@:Lf3c*h�7n�f`)�ܽU"�wi�7E��aDl�-��e�D+a
�G���J�0'p�xu�,�kIkcf�$ѩZ�p������`�5ہ偦�n*JQ�ؘyshI�t�i�,����Аὰ��Ŷ�"F╍Qb�X�[��IE@�Or]�47a�ІӌV�$u���4��:�U�s�,�� �Z�G�Q�OjʕcP���ΓK`�A���pb̵Yg�;HT�Pm�R`��KU4(��� +�h���(�ic��r����d�x��e"�$,i��\�· &��Q��iּ?d���N��.`��4�Ǵ���N��y�f�!�̈��ֹN��ݐ�s�pt�����xk�#����*F+^a\N��h={�-]] "�m�C��0+�y {�M&sZ����*?��zGn��͌�(�����/&U��6=�pYcdm?�l��"vbW��*IV`{��
Lk�.�o0L��w��rۼ�6bFd��J����[�lK,J�ha�^�"��5���"*,��Pˢ)Y�2Q����j������'vʈ&�G3�9T�'���;��hV�A&�"�,�t*�[/`�����.���lX��ux�7� �A����7�hXdE"���%X���ږ�4/L�wu1k�yR��+j��c	�n'*����F�����܇tR:�k2�oVPb��[J+�+Yɷk2E L�/"����<e��7k3v�w�ab�Ӕ�5M�;-�+��ǀ7z��4�[z���ّ�Z��ki��9pf@�Uj¾��a�"��ʗW��/�X�ԙn�"�ӕ�F�V�����w�n����-kY�������Ywmɐ�B�)Ȟ�N芍t��`�hvUk�V�Ư�%�M��^��u��2�E�st������ B�ص�c��l��R�)�۶*� +.��T��qTK	�Mf�H��i�n]�V6�"ՄHT�O%���t���7b�Ym`k0��8��B7(;ql^V�ݍ��R4�)��f�#��1,�w���e�*����٦#��
�jV���Vb[��h�ᆥZ�%�ӪJ�PچA<�{IK�`�HR�r�r[zE�Kq��J9�U!���V�'Z�[;2���:D��H,��Y�4�f�T2�] �6��X�F�e�K;��6��Z-��VJ�1v�w%��tPHl�%6���ӈ�&m��lI������w�e\��#q;BD�-��$�wo �j7�/�k8EE��q]42Ҙ�ֺ�0�$��X\�NV��nⲢ��{��IUۦ>Ӯ��<Ѫ�v�Z��R� ��JVpTJ���j�]X@ܭ��U���Ǥ*�b�W2��`�v� �8�]�e*�H���V�˽�i��m�Dl�x�\pCbY�6���ĺ����YG~�3&Ew5T���%b�M�G\�W�7�HF�
cԬ�+,US2��sH�]k	g6��f46"�4�C�v��A�6�3\�mES,��D��2��a+�"���ӱ��C1Fͻ�ƭL�Ҵn�J�9x�	�aM�0�:a�SM-�3Li�jXg�]��TT�9����u�J�t K{�td��a�����#tZN��x}���oT�4 R*,۩e^<��B��tDm%�@���dSыM
m�I֘(8f���MNg�(��@b6��X�Cu�����eC* j��Fl���چ��m�J�tựf:�`Ś�e�pH�)�rRgaa4삍��7�I}v�JEWX��Fa�,5��oJ��Z�RmjQ�5X�T.�2�Amd���b�E��sV��"��a*_I�꠱:jJ�[L�^�u��Tt8�Kk^�/ԝ�xUf��0[���ud�F���e�����;�i�A�է3e���mL�����7E����
�r��'u��J���Gނ���iB���UVf����r�M%��U`䫚f���/-eFjwV��߆�N%��bMG&k�$+n�a*o.e���#�4�B^j�)m�A��b�ۢ#HVbt���F��v�����PjTՎ�i������b��Y�W��޸�EE�kZe�WQe�BƜ��>M��D텊���i�*�DØWѡq�Q�8��l^-�����0 �|1����I�i��E����V�ܸ��K��t�a��[�f�Ŀ�n`��	7V�/]C�|����f�B;j�5����M,�^�gqT��b4R�X�@p�T��+�I�S��g�%ݲ�i#��WVa�#)�yt�����T�i2�I�6��;"v�R�'�2�g/v��Ta�3ki^d����\Kw��V^��U=V�v0��a^�/i�R�]�^���x��/N�m�{�銚K�V���f[��#�)�ca�R�3�hn4Ƥo췵3M"�eJS�E�i%�e�J\�2��c�����Pj�$mo|�\�l7L0��&�8m�c��H*ā�ᱱ�޴�^�Vr�އ��^H�bma����z��z�a�F�Ѝ"�F��3rj�Xc�ˊ�lB�YM�*���K)��[�V뭚����e`f!�+��n���\��SX�̏ [VEB���˖�Ԉ�SFQt���)�+hFj��U����d�S1Qv�ۏ4=TL�x�pV���a6��[.]��:G�J|�7��TN �]ⰱq�];�ۅ�Q�Y��+E��T�bk5(�˃ �$�k���M��W�i�V�GoX%:T
��Y��*)
X��5`�����,�!R��؎�oSv6p�+�Λ��g �xr^��v�dN,֑�h��y��4��<�q����v%��۫H��gjգ�	��)Ŗ�#51Z�޺:�V�Á���U��-*%u.%#�Q�J��Vvm��>Lֲ콚o^?����1͎^���cP��
��Җ1��\�h٪���Fj�&����ޜB��,���X��9�ث5�k*�wTW����n0ť�m��!tӁC��ۍ8v�+7x�
�(^]8nc�NpL@�b]�(˗Z9N]���.�H��sm�~J����J*�����ǌ�B�NA#����9���[zhEwjȵ����l���g%��T��2m�KJ�0aW6�8�Z�kʍǸ�w=�7p�uV��G�<{R虎Qq5rJP��iob����nfS����d{E����4����Q�b�S�۹�c)�N}
�A7(��E�T�-�P�ZYՀn	{�ۖ�J�'2�l{��i3��koQ�-.�j��z�n�R�D��M��"�@VEv��v$S+h��Vt�����mAj����q��m�V2�ۖ@q�ҋ��b]o`��V�n!�&�x�-�z���el��&��FƆ�wo�Ȯ'Qp�+�՜�.Ң	��b�+��ţn!�����Ӳ��u��9���I��9�J_Z�X�S���������p�ef�;� ·�.'�t�m�Xų��UJ|%5���Ͷt)Z��B,�4�nEݜ�3tƠsʚA�.S{Yܰ	��j�3e��|2�8�-�n����TF�nX��˫�#��u�`H��os�h=��� ���C��r&�n�����A���x�;�Z�b�pҊ�}R�V��(���I/>m�Q6��bN�3fb�JC5#4b�TfN[����[�<x�.�Pnm^��)3�)�9��N�Rɏ���7�.Y�
��X|-����q���{�(���r,��"�l��W�K��bW]�*�G� �u6�Ĵ��*7��d�ژ� vf=�*�r}����O���n��3�k��vS�u��R= l�Eɸ�
�z�y�һ�H�&�\�0et��rŎΈ��i����pȍ�����l%�@������� �M:uN\~���
�.fcsѺf�_X���i�t���²e
C-ӹv,\p�1KH��]�ԋ��:\��j�"��V8[w���pʘ�x��,�1'5Aa��޷�9�oj���w[��� �a�)h��M���w[�����L�Bd���צH�I���F��&��](q�2��ռ�M��qE��r�v�VЯ4gF�J��u�ˠ�f�;��!Ӹ�M���GA��(a��>]��;=��%���Y�j��Ý���a;��+G�K0ĦR�[L��e�{]󠰸��l�[,��YQo�W�
ݨ#��������b_(v�Ǩ� �yYC�K��{`�t&�Ʋ�S���Ftڻ��M�4Y
+�Ef�����[��[���sFx�+�u�{M%��Ӛ��ښT���e-7%K�3N4��Q{��d0M��S�bs�Uf�0�t����\�UbE�3Xl�]+%�n�P��Fo52�7�wYv�u����UԜgXF����aH8v��qA
��P/G�B�Uגvd�b���O���cc&��®����[V:@tCA]5r�u�:���Wt�N8Ы��+�k�^���UN�F��X�P�J����Z�ÄkE�����W�����o>���P{�(��Ҕ��r^ZZ�\��5�om��67(�4M�h9�$�^�s�Xw��gQv��.�!���Kbq��L*���S:Sˠ��X!44�4����Y+t��z'[�sX+R���J�� nV[$3�5uy�58�6���1�j�oK}e�Uڏ��UǱD0�h���R]�D&<L�p�/
c5r��ax!�v���f�Ҹ�n�sj/�  ���r��ct��M��&ýx�gB�Ǳ5@���0H2��\R�pR�}%�I�k9Dhq*m�|��@�Op�<���ZIf�n���&Y�,�����r��*��[�*�	:���6��D\��h8�����p���(��m�����K}�RK/N����L�R��r-���%����)*��/:	�9�y��4;�mX\S��j��W��SƎ�d�u�bH�Ci�p�^ou��$TpBn�X���k�*��n��|���3dC6�ֈ����$��X;j�/q.<;p �>�?;�9�IW]�N��l���2���^���k��z�1C�PCv%n@���xk��틠�=��%��<��Y��ۙ��ķS��B���u/>�BS6V)k)���<�Y����U�g��է0���Pkn.�n�DF������/&�aUC���/1���H��cV���m�K{{g9ܝˬ gbl���	+����t���&�����n�� �ٕ��0� �NW`H/���˺R��T�h�Hj0D�'���M���f6F�o��e�BU�=�ǰк�v���hۧ�tU����3�d)ɳ��� ��������)�m�N�N�U�sjv��i���Bޝ�l�����B̺z��,NE=U�f�X�S��o_ � {���uص֎�|�GNNױ���[�$խ�W7���Y�*H���]��P�a�_jO�WJ�3+\�V�;D���٬���X�W7�a����}jVf[���NL����V�!����:�v7�F*�7X�(��ծ�h׊�K�Ie�ҙٹp�Ё�}�j׌��24�BBPqi4�A�rq��9v�
�E]Eׅ귁��T˖���U+~�/�gL��n�#�i� �!7[�o��6uJEZ��u�s8f�%K��w����L�%�\����m����0����ܽ����T�n+��n9g8+��.%�J�|4�2e�a��PP�ds�t�i�lY=O=�hӠ!�$�±��}f�We�nü8��T,�j��X(�	��m�R ����]��FM���u�zut!�
����w#��0��i��OyN�s�ܦ{�w�j{�k�S��fe.W��$�t:Nev++)�1i��]����Z/����ՆI��Mn��ހ��+�8�z�K�h�zg�5�~ͥ3��H���gt-����v��Ư�Vun���30L�ůGH�ŭ\}��C�o�q]_M���u�k�q�@�KtCR,��g�w����w4ٷ�����D�Ƚ���-��ׂwwQ�+j���\S�H�4Ϸ"�w;*��t]+0�O�ZeΆ���顛�c��1�y�ʽg�a�u�ss��QK�;�����f�O%ll͸�N�O6S[ח��lM���w��T��ؾ�<=�A��d�qp�="M�y+뺾�!����8A�NU��C�C����:sMQp�ԃ�kj����y�d<vX�Sz�y`�K��t�p.y}����*�����k�V9r��AÅ�Y�
<:��������wC� gE���.�4��x�愹}y��6�Ő���1����@2�E���K���<z�rA�$|�i҄�h��x�rjӑ�y����j<����~���x����p lWţ>@�;�w7octd�A�˺��0۹l�[,��-�����[��d�Y�	-J�,�K*|]��O�d��x�]Yq-�E�XU+[�il�ctà�����%A�l�sz]/�Ũ�a�M��V�s�v%l����H,�sq��V2��9ciۋ�.�޼��6��ں]I��׈(V8Cc�<��0��>����ړ*\&��9F�r�6*�t>�ͷ�(A}�q*���ML�ɫ;͇{�v_�,�v�p	���F�8I��!�e7�N���mRn�ޙl#�t���'��b��^Z뼥H��a��D�y�]1�7$�wR9k��bZ6#-t賗GywT�Z���*��C$Gc΂!��վ�J�Za�Ru�h*���
��K�K�ۮE�յ��jb����ѡ�z~�8]DV������A,b%7_5;c�P�+��)4^��v���۩�$S/ds��T�b��iy�D�-�a��Af��.U��ɬٖ�"��8��4慉2F�v{�1�.�$X��J�Ś�������h�s_\�tB�֚�R������>�Kb�v�F��zmpM�*�ڲ���Y�2-�k��u�+, B��Ć��i��|2 ���\$\z(Z�$
qֽ��{b�Hp�B�Jk�$�"��T�F������cT�`����<-�]�VW:圲�	�xG͸"dͻ���+�4�sx<�]A�J����k���r�J��t�Փ@	:�d����^�؝�6��K�{a�_�3�;��ʋ�0B��N.������De>�Є�t9`��tnզ�<��C㏰�Qv]Eg�`�osw#�E]�ބ<�/9�>�l#rb��*k{��|�l�������z�T��7rG�fl�ܣ&��+�o��S�&%���7e:���.�uNO�ʝ��F�V��Ln��+������sJG�v���G/^+L��CVc�����ٔ��_'V]f�\�=�g#{yj�K%�z�����N�,��@[���f�&iUp�ǘӃ1 �iW���C	�;��X��øĤ�@�B�WL����`H�}1;�G�!jĲ0mv\n�4�gAZlc�LM�Q2��ڝo.�DU��%��F�b���bF��$�kރ:�Hn�Y;71��%�:\��m��㓯S"�@��U'#�4�P���ə׶��6�8z�+E������i�b��4~�N�]�[�	:�\��W��u	h)�� ��`��	��}�nQ̌�)n��7����?��[�^J�|�A��%*�[���k;�f��L��n �9�u���z�Y��u�ʱG�w��Jg����-��V��<t�&]��|8>����2`�o�lgkW�u��ӌ+��J�0d0���\�� �����2�ئ�]�c��Ǟ+�0�Tof)H���9��hq]a�h)鰈�ӼU6n.F
\x�2�M�:݁{�c�7�������hw�e�jh�z�G;JU�t��'IVR���2s��E�����������[���.j.����.f�Kh���k]&��H��G��*l����ҭ�� �ǫZ�ˠ^J���:BL��=8��3@P5�T�j�+�VjqƬ�kn��R>����E����L�x��}�����u� -؆>�G;�-%��3%�u�� &$z�3{��b�a��ݽ�J�/�:��{��.w��ϋ
Qb�r��-�A��'�36��+W)��<�fք��Ղt�.��T���k,��1��c�t���P1�͸ՇR�H.���Nw�TZcwYK"�it�ݐ��`R�9��Q(�4�U���Ub����\ңR�؅�3�5m�m�ӂdq����o�:��O��ˆ�d�xOQl�Q�#���^�
7MI���j^+Z�教7�adM�j\��z.�	�,���S��U'62Br���ۭަ�4$lN���q(����n�q�������ZD_@���ݠܽ�<;���|�U�hY{��Sݡ�+9md�=�/�'ɨ�I8*��QwD$%P��5���vx#�������;���ΘCA!�����nz���U
;HE�Ǜ�RS��}�Q~#>v�\�jح�U�R����S2,�շ��9RR��f�zy�ى��^��.�w�.�	���#Jͥu5�k�o{S�x���Uy~����y]���v+�t���w��<S�	�����[j���1��4�e�j�L}n�淍w�z�nXu;y�C���n�q!#�nA����!zv���rwM��6�)!�NU��c���-����6b�g@T�M��3���zo��zBV�ڨ=F��K��;��m�X&Pݴ���-����.=�����pc�)d�Y[�s*�k*ch+���ȞVݭ�0�x�oOL�*�Gf�sy��K�V�9T�\������s
���+]���Β�j���L�+x�ʗǓ�J�2l�I*���Z���4��wI���/����.� ����^NhXΗkL�����r�A����]��쒯��f�O�M#[6����G�^�Y�:�
.	���Z7V�����s��WhٳtLu��č
A��:��8����3���)��gfդ�YJ�Ѵ�,V� ܑ,��f��yw�4h�u&��2I�w��lͨ��[5�	0{S�F��ؼ��w;7�*B�i+.2��2ۡk�h�0rW ��P.�F�҃WZص��#{��vӎgT��n��3B��MP��ݹ|��:]��Le��Jȓ�aDU�N���z:� U]��wmB�=��<�u���Vv��N=J���V-� �Y��S�.�v��f>�J�=%ݒ�Q7a�/r0/:]bӢ*j;w��ut�
d�9c��b����a�D|��́4�]r7O����F�n�|�Cʦ�a�m��#f�|�m�Bu���2![�puE6�N��w���<�MM���h�𹷍�i�"^jTk^E��q%�J}yf�+����>�qa���u�d_^9�M��K7&:
h�us.r�@�A�!X�������uL�L�g��D���mWgB��Hɻ�ӨfW���$�:c��ǉndTIV�1�VUի��3s�u��P���Q��K=f��etwh����k.�N}/u-|��]�e*;���vsu����{z�5Ε
�L{�2�)m�ō�M� �v�yM�egX�!�td�t��<Qq"�3[=/��A������1}M�+���U��s7��\SY;6M��S�sjG�6�w!WVD�ޢ��˘´l�㜖b��9��Na���`�Ő�����ǚ&@�J�eh4���J��r�-5HulF݃�MO��ws�:>D\�+/7�t���Z�5�r��!�l�Z��u-.:�M���ϹNZHk��Q:��l�5К�p��k�ݡڏy��^ � �p��qe�>)��E�%;q݊z��:kE';*tQ�@��V����_;Ê�0�F���_s�Y拑VV�M^ud��Z	Dp��V�o�mE]���jf&���R�Ugq�:
R�.�M}n�K�����e��dq���բ���GZݾٴ��MҴ #5���5H6���en1}��`��C���͗�ݐ�+0LՖ����ȝ\��H���O,vWAzl�M5k%GyrV�5�8��������h=X:-K3[�ӡ�m��@��Jdt�l���Y���*�yb��Q��݈-���Ѷ-�skPn��e�B���:���`���l:�sp��E�n��!9R��f�d�U�㾼�Eފģ%���q�n�@��r�O)9źj�ws��|u��ǣk�>���!$���$���������g�׿17.��r�YQW(���M��ˬJ'�0���ha�n����.���8(Ό����x lv�J� L�_m1��9r��Xsi�cG �S�ݚ�F쑀�
wyn�R�6��]�,z�b	�������&�D�ܙ,��E�Qc�*�顀̾�WT��k�<��L-�1�[�<���GEf8j
�V������+��Ǔ-.�(��m�M�������&�x����g�";r�bB�t�V�4{m�]vl�������P��s}ì�:9�)d�����.��vl����9!�ƕ<�MY�XۓR��`��"5��뒯��{�e	�dZ��l��W��i��e�K`�B�����n�RF���V�r�����{���48ŬS��K�gr�r<n�OuB���v,Vs���TR#+=5X�xY<��ćٯ.8�R��]��WV��Ѷi����)�Q��6[}���ߴ����K�j��E,�.b��\^�q걬�Ǒ�O�SI��c�g��ك��!|���:�r]7v�T��s3�æKT��&�REZu5�%Z0�.c	)�D��/l��ݼ�uZ��g+��lG(Z��)�- �_k�z��)4/���n�U[hR�y��P�MeT�f�	dN\�Les���$���Ό�C۷�17��o ������24�\k_vS�]�ZI��
}��!�N�:[lVO�eT�N@�-0�'͏���䭬�O����n�J�sR�r�]�j��Њ eXf�ؔP�u�Q�wd3�(I\6��#�����%����a��*xx;�4J�s/�Tm��à0a��ԡ�}ځ�3�˱�Ho7�Y�C��*a�cg*���O���;"%֬��/��grB,;p�؆�|jPh�m��t�w��;P2����[i=1A��QȗN�ݰ��Z���_T�:���{x��U�Kw/���D�e��Y�ێ�3-l���9�R]$�*�g,9+*�Y����圑
tۥ�0-�/�u��>d�4���A��$St�ORU�;��;����ڽP5j:�t��6�����D�NW'���ٔz�0�ᗊx�ÛV6As)�y�������2�WA�O����PY�Į���\]�Q��7!/t!ʕ�N��2����|�v�"�8�Q�E7�́���v���gd��\�y;YL#�R�D�Cu5k�| �C�ҝ���a�v3֩�&��d�	6�Kə�Y��}�Re�l��+�p}�)%!.:J�l!���;jw(G��0�L�rD�����2��)�N0`���� �}�=�+�T����6���ta���6�7-ecU���3�y]�L:
j�w�t�%�ꛜ��aչ�g8UG���dRd�,�t`	jNȃ��ٳ�5�T�4�Y�tH;C���3$g9��1��k*4�kK�;�}���6�`*}�ᕩ��f�]����Ft�PS���2��n���Zn���̤̣+A���=�����8�A6�e3��w)u�:���m�����H9Vt�E%g.T�_<�[�AU��9Y�W���%��23�fb�*I!ٓi��5�P5Hy`=�uՔ�/�'������aT��9f��\Z�j�h�p�0��)F'd��ܾ�F���g)s�:p�,�b�e��Ȧj[��ڻ��zֽ�:�6�m���2m7��ڕ�&�Bź�m�("ٱ�J�}b�K|���2�A�eb�,և�Qq�ncF���F��t�|�.�ݒ�n%��`�:n�����o)�ŬuE]z�0�������H�\�c��*�Af�Vv�{}Yl�;	o>T�z�#k�g������|,f��R�@��:�]7@��.n�T�K��9���_E��)^z�t��p�B=�����.=έ���*vy�VmSȎ=]7����B���Z�#WI��|�'#޳Ê۩w�ml��/�@���[���z�K�kk��+�����wHL�����]�v�#.;ɏIyjRg� e��,@��Y;�ЭR���}v�+�M/�i��/	cJp��K�б���`�ң�(�32�Ĭ��{*t+���B:�<,��t;Ǵ`˛���+wl��o���{���YPU�BÌ��^k� ���0�YG.;���Ĳ��.q�Z��Co�t��U��ⵠak��#0U����U��A�c�����-v�m9����{b�(�i���.���r�mo'Ѭ�]� ��m3�т�Fड़ڳ9�ݕ����]�*�%ЋN3��$s�4iݶ&����跌$�oy��Ukg��e;�P�{�s@����f>�u+�G$ыN�FU�d栐@�(�����(<�pf�m�1��
+-��9Вg�y��V163� �0��:6�\�FL�}��`�\��.Х���vTĜ+/F�з��m�r�D�����)�0�{�n���wغ���N
�t�$κ�A��x�J*:�Ӳ�`GJ�ͩ2���/�T9��2q�(�!v;&��΄�\�s��
���}�J*`+�.��t�d��Iw��`���mg_&��CrQ�%�J��RHnq9���l�o[�\V�� ��G�>�w�M�W�����Pv��/]�)�*L�n��V�8v�;��[+S�̏E��J#T��ͦ�gwI���9�ܖb���2/�9p�(@���j�+
Y�G�m_e�npm���o�_l���"����ńԸ�1u������;	1�z����"�9ϒ�/��d���e�-ǻ2͉�'9L��|[�o��D�[�D�v�J}�s��otM��ڃq�M���=r�N�xC=1K�笝ӔA�ƭu�a�%�l�iA���w�+Z�/����Q.�c-��jg!n]EESuݭw�[ˑ⥽�K嫮��e�A�Ret} K��붂}9�nY��ʾJvވWI��F@[w>.�2��.+َ�,N�G+�9ofdP�����g'����n��8e�ӵˡ�����Ϝ{F�9!L<�������N.f�(?��wV998Z\,Tw�.
��q��Ʒwi����]c2j3�i	-��9Y��	̮]�;�n�Ֆ���5a �*(�7V$�ѭ!�77+>Uu^(6��ä�1Rl��|�v��	��ٝ��z��V;(�8�3w��e��|eJ��֙�s&Xt@�z���ԣzh�zJY�\G^�0j[�m*�ܫ��r�Z�p�f�������h�1f.������g�&v�s���c%)h�u!mvP֞Ï�<�ѷc��V�n6����3�A���|2���/2�>j�gzk&�2�:�	u
�#�J7qNMջ�<��&�H���*
oo��NT�
��<�H9��z�V��7oi�zD�[>�Ò����-��0)�oH�IűH�	�����UCbSE\�{xxl�i�k5L��L{'̫�u�p�6* _FY�a�H��9M*۔�)G6�\�@���NάV����n���SN5����Ik�:;�"�������2Y4^�
Ggn(��U)\��'����Qr:X�K%�xl�ۻ`-v�uoU���1+rDt�R�\�>�+G8A�9��3~���ZR���;�ek�nG�\�t<[�Ww���*�[�T.t�Lv���	�*+��w��Z��4��l\���6�v���@��a£���ܻ���)�[�i�yc�|!]"���[����7ղ���U\��D��hEʾ�4qPgl�}3��u�S��ѠP��u�Z�k1��N����\�yx�Τ5�t�'&>�SH�a`J�N�K�V���<�W���X�sl(Ӯ�*�C��KÉ�Ɋ��;QT*�*.�J�ܙu�%;M�r��]*�R�n�A���/Q�v��Ð#��НT1�un��ܳ�i�n���6z�͗��u��{�є]��ɻ(��tb��x�S��x��C!�!r���;�lX0��Y)��@�qWx�[x��&����)1���%+(��Oо��kR�9g�Ue�T���O(��ne�;���f��eb�2�q�$�.*6����G;����5H�7č�ض�Ʈ�E>� ���V�.������tO=�C���UVa�M�c����ϯn2� O.�f;;��E��D�[�����WM����R�n��U����B�&���6���&K���3:��.���D���G�:D�69�yfOZr9&~dͭD�V�0��r�Om�a
%rmh�|[O���;���㯻�PЪ�
T�+�������������ü2�6S�+�iR���}�`1��BqgX��Ẅ́:6;�lR�gu^1��$k"ܤ�a�#O�5��b�Ѧ��[W؝����w�Q0Bie���I�v	�����[�<{*t��KS6֜9�2�lQ�-(Б}s�)n<�i�%C}$�\L�����c٧�;(2VF���rէ�̻�*u�d���� Aj�+�3Q.���A���B��V7P���-�������U������%+ �d��'���+���u��vn�=L0�Pբ�<�T��m�QO��桸��W����]G��L�M��c5J ������vʮ�m*3n�9��[׽�=�r�Lt$�1�BWgu��J�sj8�dt��+��V�B�z+��,QvQ8ܾ����E��Z��l��;k]c2�p��A٥��Ft�{����2�K.���N�R�M���`اA���d�f��i����z��O+*[���H���e�����Ϸ]��c�ؾ�@-��6
)0m�b��{�����F���W�%*�9dlV���=#acA��A�k��]@�K�J���<���R!o�,�d��1X�R�9F�6ɤ@�DˌV�RKXv��E�x��[�/��p��S��Sw�,��Q
GNtS�u���d:�1g����j�R��k|R
��,�P���8�/$�zӬܷm���X�ZΣwVhkU��f����LP�;Q0!On��T�ך�f�|>e�<a��Y�Sq�:����-�n��������PXz��|�91�%*Ϣ�b��� -�k�n��67�([���uȘĴ7�l�+n�*ޗ˽(@j�s�ҷ�g�{7��\�K�(�#0�V�Y�����t�a,�x0��2q�
�A���X�Jv���G��y����7�R��B��R�;��k��ɾ�/���'�A���P�a��w^��WeYෑ��*��uF*tn���w�,��r�Z�)rbq���Z*�WBi�^@��o�z�
�JODH��K����LV)����F%:��Òa�b��c -m���wm:�Z"��u��W[��Jbt����M;��9Fd̓)��]�xx��L9K��P͹v�g
!�ԷLajELS�D��h�h�%�l��_#��)��[�/e�ޙz��t�;7`M1u�X7V���m
�c���zf�=���9t��6-'Y0�/Z3�뱟/5�-%}:ju1Iv-9��e�+N���Q<|����3Y���i�	l;RL�`<�Ol<oop-��WVPv�M2�<��@��\3`D���nъa��>4����x��<���$����0PI�B���κ��m�V�x��v�7�	�s��s���Y�����sGi�wxp.4���h�<8�x�6����/f��R^��-�I[�f���Vic;��0;r�*�܅��2Y��n[e[h��Xl@����fNƣ����zh1k����J����Uq�VX�2��1d�.����Qk%<T�9���f$�kR��b3���)>x�#�U� i5'%C��V6�{˂ð�	���`]DR�}nB.��3ݏ��\]�≱{ܫopWf-}a�r��F�d���إ]A�Z��D���[�@�.k[��#��W ��v�}كB��	�Oj��}q-���d޷0���,�F��i�]��A�������m�/b�5�����s�˔���J��su]�E��������7gQ�#�@�B<�%ʓ.oE
\25�py�k���1nA}�p�3v֊����]�i{^e�b,�l�N�^F)�v�z/9>X��5���t.���{��6^�!ܥ��Ԯ�6'�ΘUP�em�y/��5��d�q�WE�#���z6�Ī%�S����`�,Rm��������;#x� %-)�ыﲰzy������s��\���7�YZwNn�t8ַ%�S-�5���Z��w�T�t��JvcM*�E�dɷN3�7��ut��kbZ��t�+�U��oV����t����R'��f:u�����Ăs�i�J�7K���{f�5[\����{��z�pɒw$�-����X~c��.Y��耵��o:���\�����#^��zƭ�����9�uЅ_X�%l���x���I�ړW�Vr��L��j��C��f7+�ɢ���U؛��}ɾQ�Gb,j������ic$
�M�+Xk������N�Hk333�y/�:H؎�%d��(B�{`Tf�q7�5�I��.��u
x`�/��{��t���\�b��°�K�TJ��o���8�s��g��qP��y9��Y\n��aњ-5:��؝p�s	B���EHkݼ3�^#]�<�fm�#���oz�2(��N��e��)��;�0]g:ɝ�G�/��s;nG�V�P`p�sH�b/w3o4�Y���P�8Pn-��LU���b�e��1�IZ�]ws�1E��/��Ub���G���P6^�j�V�+̛�I��Ba9�����ΦӰ�G��/~f�ɽ�M�.*��g50���;��6�}V�,U�\�"��S7���ֻ�m�����3�����sf!�4�H��O_��禲5������}���ި��7�v�/&O,��xNNTm�����4hźX9ؗ5M]F��	���RQ�Ӄ�9LP���C3��e��c�ѩ�a�ҕ��F:ʺ��A�(W.����xOֳmnW��H΋��$�V/�v�I!G��x)��2���Gn�n�����Td���,OA�q��Q�npb�h�S5Q�wr�(ُs�U�PՊ��:7`�Ѫ%�䇓�9nT����h�'ݙ�7�j�V�бu��+����r-e܊;I�	؋�A���B��	���VD�:[!��#=�%�N)�0�1��h�����h��ƀ& G]O]���H>U��u�����PQ��W�w�&{-�'���"�/Mv�[�Ze_[F�P�p��ҙ�����cw+'f���dm����� ���}� 5���e�w��j`
��b[kwH���#V�)4h�ʣ*M+]��(�r?B�Nw�����;�~F��岯g^B��J�l�&��8��"�-�/o��:-n���5�ϛݻ/�u�v��Kj"��Q,��:J�pG��n��[}A�]P��=� �����Ų�s���vƌ��Los�ô
�&N�;�D.]��/u2EfL�l��n�,�&��,�2>�/�L�eb�+�{f��Ӗw3�XڻfUI.������{�3��i��8�\%L4D)�E��$���fUi���m�d$+��Bj��K"��H�"�(�TQ�UU��R��TQUPF�X��V��b)V�QE��)mZ����X*�*UA
Tm�eeQ�Qh�Hڵ���e��*4�T*�ekQE)J�1�V6�5*Z�E�b�Ub��h�A��-Q����m*���Qj��(�ie`*�*���QF(�jQIP�	DQR
5*�ŭEJ�QD�b,Dl��(����)mlUaZ���(���X
KR�X��Km�PX��(��J**��U �mH(""UeQE@Q�Ċm1Qb��D�aDUh��R����-iTZ�TdL��A�
(��)1�F(��(�Tc&#J��U3(�)TQEe�+�r�"2�H���FE�m��1T+]���[��y���w��qW�v
906�v���=<�>-�2��&�fۛ����WNd恐9�x]�R��ֵZ�{�Uk�JE�{�P����5[��!v�g(J���:����?�Ȫ�m��^X����>;h޳w�v�(*5�u��u.��['B���BS+�@�8q��:�9H��}�k����0�˾�՞D�o� �E�f�+�6��]�^?���Z1Jғ4.Vf9����K7�
�/y��؜�f*1N
\��V=����f��00���a�*�����\�����b�[倧���k!�j��4N�U��ol�Sב�X*Z�E���w��:���q�/�p�ؤu�H
�����[�B|�p��z��KpV����s%�cfCѕ7�!���XRȊ��X�-��! -o˞X��k�Kl�ls��$�j��S%[E��8�\._����I��xY�*���}'���;~A�j����xⲮ��:�{_gN��ީ7����c����=q���;qT���w
�&Q�.�&q�[��Ύ�TI���t������(v�g��1��5�2g:v�N|�^t� �o���i��ʧ����0���x��B��}1�9�r6wLe�i�ߵVx��|-[�~��*�u
Zg6�Z��3F�3�����d֮�5�H��_6HUųS�s��]�����9�<K{*#�/`���V	ܟf�n�NBb��v��[�2��͵u��ˇ����q���8����m�\��
%Q��� ��j�0��z�q�}�H� F%��quI։ڿ��q=�p�L7o!���o��gpd�eOoM^_r��qU�`5*��LpwknZ��F�:��w璁	VԈ�o�u]̥�`�ޖLJ�����P�`�!@>�V�Ä�wq��M+��U	���Js'��]N5zgM��W��()*zM̡���G,��a:��]<I�zr�b�}{�>)�u��{_#�(��^��%�<�/⫴�Q���!T�?l��0)ҧ!ѫՠ7�����.���T��?==
�ø(�M/4�Ȏ�i�9��U���0>��j�[�AI�0����a�r�%��d��"�v��]�7a�YD-��0DA�����	�=�=8��YMk�j&��}�,1p�q),���E	�P�4'q)1z���3!P��Ж�g�f��rzo�VR���x[< �jY6��`bˀ�����G�ߎ�6��bSX���u5p�/
�㫦q�i��!Se�(
�<�Am(e�²��\&��:Ԏ�d[O5G�b��
��c��379&.�x�dAܺ�u� unj���=�fC������b�=��cb��[�kU,#� ��îFyF�,˧�&�	gL�k�m}BKH?���#f��x�2�q펱��Ս g���[Z�Uc�J6-k��K����ϝ|��>���^V+�D]�K��:<�vzU��Tr������zg��u��I�5���7L��=�~7M|�+��e7,Gqt�@r7�>^%��zg��-�?Su1s��<Lą�v�?d7�%����m#]�G�ʮ��et!���]����r�	��œxa�P���SM2K1��1�ܽ6��.+�;�H�Ѐ����=�^e?<���U9�?0~������+s�\>B�_\<�c���3�t0�/X��R%�mt��4��g��U��(ԉ�eT!���!�/���hpߨ��^G^�]��q����WQE4��E��5��pU�W"��aTU&-�*;AR1{��BWa�Jx�]7<�Sse�Jf%�S��ƈ��l��j��8O"%c!�v��׍���6a���o�m1��mm��2���s*�ps���1�T�^'I�#�pt��>�׫ �7��N1\.�EO�,��9ʌSg����T�+-㷹�Ӿ֓����A�{0ٯj�u�B�q֫�"Z��n�W�ٌ@�vn�ճ�	�a:�}��@0M��<7F���ǐ�INW����$�u��B�&�>�դ��*y�������2�F
K��;�M�#�s�n����%�'J��;��ޱ��o���/x�R�'^=����CɁ:�[W����C"mHr�k�*����\�	*���J^��08'-	<b�cr���o7jy���U,���'}b��y�ڣ�S֜�-|�N�ܗ���uU�h�za��aa���Q�����iC�3a��9�:� ���v���ڸY֢��nN��M��������c8eD�!�P���ڻM���Yo�Ֆ���-��.#vF���@r�b:���s�n��U|h�
��]�7]z)�Ĵ�}�;;gR0��k����*"+\��b�b �x��G7u�T5�Q��"��(�&;;ZOg����MC	��W3*��_V����(F\-�k��se��5�'I+}e;�����Q�ה�l��H�o"�|��:5�<b�02g�\�o�+���m���D(������^�^B��#o� O�k�	SC��"�Lm�./o{�����ט��.��6�يT�ñ��Y:�����,���g]c���p,'�{�櫵)��縎�saT�Zck��S�3{��gu��[jU�]���uȆF��E�c`޾��Y�Q���;��;�p9�&1S���W��B�՝�\ԛ��8�M�c�&q����g� �r�+@�ȧt* �B��B��jܕ�����U����|tO'I\�W3���NP���C��H��d�e�_�JM<�#C�
����羾4�����K��A��~�[�MVogQj&�nu_��ҍ�z�����þ!%�Hϙа�Į1��4�ϟ+!��B*���N��Du�����Wd�����(�a����<*���U��3%i�B)&kE�}V����s`�:T�U�K��w��E51`�o�Q��1�ҷ/�`_���4��!���2V9)^c�s[���jDS�|�ٶ��Ļ��Y$����{.��1�\��8��g�v�o;0')��[Z/Fg��s�I�ה�F)��'�p�=����f�����QY���G`�݅�ٷ)�n�p9m:��V�bU,��h�h<��0{
��̆*z�Br���0����oTŎ*awJ���� C��)�)9#a=� _�V��ח�hJ}�94� ���~3{�m]�iY����.Tu�c�^+O���[�|{Ֆ-Ֆ�&qip��҅n䶛�}E!�8�3��z���Wwan6�ƈ�/����s�X:���H�$����z�ҩݐ���`���˅Ū�]}ʶI��l{,.���u�7�
�y�3����������7f5���2�P�L��Y���ޯH׏�˖叱XveVg��3���O�CW��^���j��Ũ,*�E�0{�M�a�#�s�n�;ˆ	^�gN� D��r7�/�zWY<a�q��N�q���T..:���
�[+�����Ҙ���]��du(��ͮԬ^���(�c�*W%���T<������-�{M�/���O�1\*�s4���N�㷽�6?.�f�7��GT%��f��f��-�]������w>r0���ް����q�J��3���7�_��>_�~ݚ*�:Xp������W��:�9� A�Y��l�"�];1��%��ȑ8�{��ؙ��� HWϓ��3_��!��)}��a��C��^�!ϙ�Q��&���py��+C� E|�H����72�F
p���oAL�PYd�j���0�0���h��'�m#�������<�,��7>Q�S�_)^>˽�1���js}7/�yn!-�i�1
C��K/�C|K%z�={t�_T,�A��pr/v���J�샴a���\��☎����j2l[��©�.�T��ʼa�1)���VۛIbO�|/�n:�7]�Ɩ�1j\��[�pvp��m���%�ُ{�����r��#�@���5H��R�s��*���=�&�d�6\���g��C�/mK��|<����,l�`"{e|��b�fJ���T$�}�+�
�2ƨ� ������n�ވQ�|��v�Z�������gA����ݔ��J�7`�$�a��'.�.�C�!R�}�)���Y�+�k�~(Q��x<-��*>jY4�OQY؊>�k
��gr5���F���}�b6i�<'�V�#�-f�Y�8��q�^�����&�f���c��M�Ө�l:�D�]qWX��".�\����U�}��[���c��_ ���;1�B03��jv����
�H?yq���@n�ԃs��dx��[�#-�֝�X����ƌ���S�[u�duTPW��h�m�h�v8خ1��~l�}��Ywz���jz���[>�z]W5:�&��.[w�;A�����q/�6Xʉ��= �p5X�pws��۬g�5�U`�7�}(�U��enD����'�uN�1O���4*98L�/����方L��^rG|e����m �#[ԳV�%J�x�f�ݫ��*�m��ե�W�p����s�#%��7�?���ZF����s�EԦ��$�P�do��15W��
���;h�ޛȸf�jz/(�T�m��FQ\Jh�,�$x��\^�낌Y'�,gl�s5�E�c��<�O�@���aX�����B�Y;0PV`�����
�򣡫ɷ�eu��Jk�������Ҽl���<M��g��?�7��Duk!އ|t�D�*����ܹ��ZO��YV�0��WT�ힵ[��G�,c�)�U�ޒ�����&Ż�!)�"��0E���a����0+*�M����I�CB�����[!�����}� �z)Zޣ��>qI��neq�S�2�O�nvNiBwS*9X�-)�4�y�S������ϗHe�>�؉��V���(�mX۞�{\i=�
wC)��#�u$z���������dr�q Ӫ�Q<>���wwڜ7��0�³�a��M�Qs����硏�67]�[�sEl��u_c�p��8�&ژ:u��x�D��R���+���&��WXO�Wj���tV��#z{Jz!u��^X�v{� 5�\km��U�A�rKޘ&{<'S�|3�|r�ܣΛ�;ء�KsD4G[�<l��FmX���c�k�草����=G#{�._z�A��YCPD��:�e[L	ʢ,�����`���-���mXaŢ}.n٩�\{�Z���Mܱ��3`�+_�X�'g���C���ȅ�L@�S�F�SOs�:ŝ,f�&�ʙ^'�z�rC7��A���^��"�kHO+���,����4�]�/���&�g<��{
m����Q7.j������o�:̃~����A?��o��WC/[��~��j�/>�R3(	
sI;e�:(�g���OuJ�ѡ!�;��[�a�T�1��B�B�����\]�'�4#����N��鳣�7=�"�ͻb��ꠊ�@��6?F=�4䣜A�K��X�ð��v
�F.9��Q��c>�
�������rP�"�EW*!+M��8:/v@(9��W��[L+���AcQ�m�qR��-d؈�Z/ݶ�#ի�ݵS���F��s�ܢc(�xn	\c/���t�AʚW�%�*W	��0�;����jWB��xg��,�GP�g����~�s��i���`���W����H���egrGie��P��dW֝������^QQn�MF���q��h8��3lgv�ޖ��]�D�-�6o�)Xx���̊𐒍���JQ�ћ״�'�=���Jh���1��� �t��o���\qF�����~�
�*�ֆhG�+�'d;�3W1*�m� dt9�@�r�`��y�t�.�i����m7��v�N����{�$�%Q݂�)!�c���RDe}���-����D�ԲV]�X��-}�u�ޚ�\�Vl�9�>��3����Xw�y���S��i��ǻ�^�p�EWYh�!uQ���'l��o������I�8�n��r�SĪ�~���G�:���c֝'��1��ҍ�݇�4��JE���b�+u���|%
˵�
���/�S�".9�1���4�-���ֆ�'>!�,��	�7%ak"��0Bȷ[d� ���ݟ�k�L�8 ��|�D��W���[����˭��L�o�7�i8!��8��쪾��*�K>�R �+;N�a.B��Lk�|����<��|��s�4[�ò#d	�(p;2���b{ñ�yw,�ԯ��	s�!ׄ�=�}N�<����l�w�*!��hqͫ@--b��w՞��%�'h[����+ q/�M�JEBʩ�9�Ϟ@R��������*�h�#1E��K�t���ܛ&�\|��%��!&��2�Y1
�h�ͪ�k��;��,W������X��3��x�u�س�+��ڨE�N�6A\�%k�W65M��C�=8'�9b�u����[{P��������h"3谑Y\���0[�G �:&rɖ�1e�P�S%'V�iרB&�wZ	hS.MI�Y�4���;�kp��v���#�����X��Vѧ���̟���O����ש�7�vQ]5���>�תŅ�-c.�$B��U�Y���𙨫�S��s0�I��|�"A{ɞ8�i�w$"�ŕ[3&����Sd��	�\��=�Y��Gf`R��Ly�O��|PN6.&�N[/���bCt�����`�L*a��u��j���>�u�����*���'ͭ��ի`հk&Wp���C��xrN	�z-w���s����	�f�����wx���u�h@y��t� z!X�/k�Ve����f��ݝ|�2�48���giKF�cJC
��N�:���c��9�΋mX�`�:&*�C
�Ic�0��פ���4�f��5y�g�A�P���H]����	����������`��q�t�Z�;�׸r�W@�q�,���8�KE۱�kw�	A�r�Ů�mk�"P[�51R�#]��-��a��~5�(�#6l,;��{���\�nqQt��K�A8<��a�-��+i��QYԸ˨E��Ne��P�l�;�R�	�l`'�v�Ɂ��X���ܭ8��\/��т�����H��e���׸�F�C��*K*b���t��3]�TH�]�3P����ɢ��A⻩�|���Hl����@�Q�d2��.�Y�r�����}�6���ζqSih�.c<s�Kw���]i>=�;�,\

�]�8u��4�q���d�U]��v�Et��8d�<�c�fK��U� x��'C����SMu�s"�p�fJ�Ԑ����̰4��{N��³�\e'��l��Z����Qe�pǂ�/��'�����_ٙB�D�蛪�r�=mt���л樑�N zek{g ����E�kOV��$��Qv�3~��W�����s$�낳�"e�mk�s��Sh��L�W0_)�Y�nI�e�j��.�B�Uc�1tU&,�@��n���R	8tk���sz��H��knn`QVoMj�z�!R�}C�4'|ņ(�M�J��Oj�������1��@��{7���][��N�������|��H��A�R�u��1��
�h�͔���ؙ5
b�nt�D�z\��.ptL"���+���1l�]�*8�ʱQ.�]��s��춳ʙ}�γj::'� b� A΃���.���9�����6-�U��d��/!X^ST��N�N���Hqs���0Z2��k+s[��d3e֎�������I�ǂ�U���|V.���9���z�P�p�"urkO1r:�p�b�s�<:\;�g-%r�=��������Y��N�mc\�t%b:��m 
]��Xx9�١y׸a@;L`�����X(]��6ֲ�E�Qb"�U`���-���ES"*�iJ*#ki&5TQD��*)T�
�j�dE[aF,E`�"���VTU#-��2�`�-�YAeJ U�ұd�-(PEb"֥-� ���h�U����
"���Q�VJ������Z�Kej�QT �&%�1"�X�A�QE�X�������`��
��m@Pkb�aEF���
������bA`�"�ҵA�"��AQ�e��q��,b"
�f2�X֠�"�"��*�UQ��J�B���DEYb�YX
J�m��,X�T*��F�"�wV�6�R�A�9[�ٲa�w�q��}(��G5�e�	3[*�<��ZU��o���|H|�s���=�d��qҌ,���B�۷��|�Y��/��q��ATݲ"N�f$є1���q8�M3�LH/���N!�C�T>aS�~�{�����o�g�ϒTJ§1�Xb����;^�zխ��׵>��߽�qP��I��J����.��|��4�Y�wz�\|H,�,*T:�T��ܢ�'�����:`Vxe���u��~2�3�q����&�} x|G���9[�'1�����{|�_e��m��{�i��$�N��~M��
�����I�
��U���b��5�c�Y>M!��5f�8����lY*N!{eO�U`,=�������d�׿���[���߾~��t��6�OS���̀�䟜g{�N��a��z�I�+a�����u10����'��J��>��&��1d�혬�/)1�ˤ��>dϩ��&�8�o��;_��o���w�~��޼����f2T�k��������?�|�>���I�:����ɻLH,�ܦ�I�l�A}�u�����y��|`T:�^~�m���3L�1N!������2��w�;�������z��*z��CI��iY�J��vy�$���LM���~Ir�5��$��'�sz.01��s��a^�$y�d�J���I��w݇��Rm<�u?z?_��;��7�}���>�Ο3+�
�o�E
�a�?&!�+8���?'��iRu7�����^>~��w�&!�hu4��*c�7�2T�B��.��kOP*N�S��L4�OSHb������}��4��s������
��N��ޅ�d�4���nJͫg���=I��b�z�Oɟ����$�ǁ�ÿP�AVo��I?!Rl�C0���������Y+*}�}��/�����������k��i��!�t�?h�V|��I����� ���f��Ԙ��*n�%k?2V����?8���bN!_:��k�@�I_����O>g��v������1�������������Na�+~v�{ϲ��*�;��!�:�</앟��1=C�~�sĂ�|¦��y���<���B�=IY7��4�$���ɞk	�4��-Ld�>B��HN��xG�PN^����E��,V#�@饒��EBy[���r�ӳ��m�N^��P�������]bg2O�^��<�2<T��tPlJ�jb�y�']��%�DA�:�1��̗h1�.���pkj(kq���
\�q��Cz���owj���|���T������I�}��u�Ĩm����C
O=��:�0�
���6��b|����23�=f!�{�Ad�{�M!���ܵ}aPY��LD��k�N�ͷ_o3�����}�>@�%t�Ձ�����8�q��<������I=g�{�a>OK�d�$�9��d�����!��o5���ĝ7��ֹ�W_��^��3�ߙ���^��ğ!PԴ��'Ɍ�4�ݛ@�VJ�M�'��1�C��C�/,7���$�����v�Rb�}�2u���Y��ȡ��'�$��������s9̾�}���3އq
퓧�y�g�������k��Ag���
i'�l��D��M��Ax��0�8�Cl��&!����:�r�����R!�պ��#��ύ/J���&*��٬�}��ٶ��$�;�r)�>I_����$�T=I{�膒u
�O���sbO���Vx�yLg̕*f+�Xu$5i��c�Wx�3�>La�~y������Ns��秹߳o$b����`u�73�jq�!�����1� �׉3���*i'�*l�k��$��<��Ci�'v�°�9d��|ՊL@�W��E��Rj����;~��Ͼ���t?r�����Z�����1����C�:�O�é�� �Hx�=q';Cw4��T�!SÝ�4�'��8���bVM�Y4�:a󤘅�!�|��g��s�R����;���w��P�Av���5�I����'�g����!�������T�B��o�a����䟻���O;M$�g4zɜ��iƩ1E'Ύ�W�#�DD)�{�y;�To��j��>����~a�����8�'��hi ��?O,�i1H:���՚IY�߲M�ԕ�>OKa��B���s�B��
��&�z��)��X�������*rc6|��쑚��o�}
�d�P�;y�)* ���C�Sl>a\g���C����W��Ag�����z�$ߖf��4�0���0�/Y�9�6�ԩ?!~�k&�u
���y�y�o������-�*�;y1�.ƽ$
G(���U��h��F�v�D ��h��w]�':���Q�ѕܱa��E�.��A5W�.o��n����Y�f�}��fz�Ȃ�V�;p�xk�}�wX����u��>� �Gގ�TaXW�Y;��ECi*R��$�,��w�T5�O���fPĜB�d��e������~��z�H,�����w��������I�w�?_acǢj����ԇvF�z>��4DH�Dya����J��v�f��Ę��'�}�H*�R^wz&��Az�����C�J�ȝLE���SI8�O�?8�k2��W�x�SO�
��:2ս\��~���-/W�~�CG�_�1�v}q�d�R|�O��b�|�3Ă�'��N��8�3�13��D4�g�bl�<�z�$C}��Ci�~C<>�v��C�K��:�#�4F�<��*�w�ޞC����1P��|����kI�nytϙ.��>��MZ�]!���&��J��g�<T�B�{q'��c�+�ݠiP�c������Af��g��1N#��r�NI�7꥕��1T8�C٫&{IPY����I�k�i6�dĜB��a�z�Y����1�a_ܰ�wA�T�ӟf޲TYY+���q���1Y��L}B>�x��m�����z�c�h����C�:{�u�LN&$�~��WI9���Xb�x�'�3(L�4>v�8��<���m��&=C���H*�!�u��M�����n<>�|~c�}Yvu�q���Y�';^�aS�,4��YϨi'��'u�mX
O���ڒ��X��Ʋg��'Ƭ�q�򓎓�]�`"d�^�i�C���1�a�w����>���G$�Izw�4/��yb}7�Hq�
�o�u�'�~Cx~��!����@�T?$��7揙<I�*�k���Հ���1������䕕�箓H�d�S�0�� ��">���q��FFWh[���y��I��c�;9͚�P�LO;�N��� ���Y�q8� p?kZI�T=OP���i�*5�<����R~3�&?2bN���Y*�@����aXW߬�k:g��u�/������~g���bIRt�x�}d������N!{a���� �LB�Cfs'���CL��ï�8�LH?���}�����d������Ci�'��6�]��%��o9��k��չu���d�=+)!��s8���e�Ξ8;mK�_#8�����8�y��^I)����eVV;����+�O3*�����c��922E/���S��HT&����r�o�t��f�Z�ݸ3�3�r�H��%N��T�U%kr]��P�Hb=G�"4�U�Mn�����R�N2g�<I��Y8�E��g���p�I�*q����������<�~d�c�OӉ4�ɜ��xg}�6�d��q���u�v��9����~.��\ק���Ys�'�f��t���z�!��1�bAg��{�6�CĂ��`z§P��3�,���b��y�`i�P�9����&$��wy8�~Z�P�d�f�oك�����{��""G�>���N��O�%ea��������Sg��Y�ϙ*��XbN'Ɍ=O&��X!�f��u�4�Y��`|͡�ma���'YP�=O�4�V>�" 9����:��κ�^C�%&�6����jq��LI���1�aU��|�I�*~��5%M��*�P�i�J�*2�'P�Y>M�Ұ�B�M�S�M�!P����+��!�������Pg���ɣ)��+�L��n$��gO��+'�Y�w%CI��g>é�4�0�;�h�%eg^$Ǻ�!�6�U������I�bMw�z�ɜ���t�Ԩ�z��M��">b �B's��(������t��;��?+I��~���>K�Cg�w��%~d��I�����%��w??�� �'�>�BLz�H;����|Ci���ﺇ��Af��y���?!��f
�XT��;����wF���������u�=x��1Y��HJ���& �%�N�Q�|�eCc����V�p����yV&�I�Fvj$dՖ�ۅHن�K�q&8aɄ(<(p�8j#��*�i�	� k��N�C*Y�x�W��{��_���5�`��=ɿ�R�t��q _J���~ӧ�������lR�*��q�3N�Cw���kہ���7).q!��}'�U���r�5=����ު��Co1���X�c��}����ܣ�=o*
�Y~Q����id���&��D��p�D

�(� B��b�l�ĝ��ϖ�f�U��.��<q�
kq��	�Vn�s=W�:�w�l��܊�BgEA���3���h{�������?���_b5�P�>�<{>�D�(p;7�;��v�K���%dy[�l��J0���a3q���ȀXXn��G^Lm8_�61P����q����sٗ�':k���
�0�3�MK�&�'��fC����c��� s�+�D2��B���eZyޘRS"��0�x,��~��MXޗR2	�8���ev�V��N�H�m_׾��΀��>�{ֲ������o�G�[Yq���o�$@�	g�]F*:Xl���;%N���#������n��6����� E��F��J8*�n}F�F��U���s�d;�@�IX�C�$�w}��&*:�s	�.��׵T��`ʇ�a)]A�A��ꈖ*����z��HH;]�zq�. �xk���}_7�ŗ8�������;~B��D�f�eRx����{D�C�n�Z��?!�����Vْ��x�8x�٨�Sp��$����2Kz"�s���l���.$�SU�*0;,l�B�����VK̕0ڑ&6�16v��@y�ڵAK�=�R����r�i�q�f�m�/y�1cȮ5F��E�H�����:�8l(,�Ӌp�oe-X�C�7�M'�h5"��8�y1��F�nl�r�C.��ui�+z� S��҇Bzq�6�ŗՔL9Ͳ�Θ�pF|�C��C�P[f#�rR���TWf��z�g��� *��~���a��x��������? ��a��<�).Ӈt9W�K0]�����Bܽ�0�����`�d]<K���8��\5�̄�3�NtO	�>V�\�������$)�]w��4s�?eS�5U���_0�$t|~a׽6S�`U�F͉K��c�������n�����T1�M#��:�.'Ubκ�/����L���v�_ϲ��)oF/�֥����y���]gԼ�9��xpD����z:����~���>�:���iǐ�W�q92�fX��z�GB�c��������yg�ʦw���0���]�aKE���0}l�\�k�s�br�8�(k��p6��)��$�}#�ox�;_u{���A�:0 �Tb��J��5;�3�n���t	o2ጃrx��BSD���?L��W��5kPun�a��I��\j,��
u�r!�5z'�U#{����G�s��A��W��փ@���My$ey��^{�*���k]
�0Mv���Lk���ҳ�U\���+K�,��>�7�Y&<8���A�1���ntɴ��ܒ�x�(\6�_L�9i�]�E��ȯ2h�t�	U�����	�en��F��HFN�Wv�7DE+o��:�i
��	U<���U�gKf�:�n��wDM*�'��v��k��.����̌� �ơ>(C�=�.��9:C��+sNr�/*�O�36Q���"f��޴r�=P�O���k��^$9�*ϲ/V�qr�|bD`I�2ru����<��W2;�����s���I�
�Ƀ����D�B���?[;'~9��Ɔ3&sDF���Wp/��"4Wͪ�7T�� 9D�R��u�7��K��C�%�vJ���u�a[�1 ��Tg�r�P�K<b���]�%{��}�Z!<6��*��1s������[�)^֍wUi�<L����u���Ķ���Z~n���ɋ��u\�7'.'��HkH�L�������E��ϯ�g����l��W�?d{Q���}�0���b"����5%��M�q���K��a��8PφI�+���s����◆;n`�5�Ĕ��S�-ݧ�/��M��3)HM[�	��s2������_ڄd_o�8�W7�`a$l=p[�'
6�/�巢�ur�d)8�r^�3�3 �}�9�ƴ���l�*�|-��j5�.�Y��������aqĢ�tYOqvy�&u��^w��$"��;�	�z*ţ�+&da۝\54(�Dՙ�K骶����-m��bϛ�#m]}���\;6D���Rg�؝lK�C����Y5���:���8=<��Ʋ��c�f;!�1��U��X���|�Z�<�<g�99w���s��D8�=��9��r}p� 'M�����{(EC��$dGd�+>�@�-�VKڸ#���w���}�=7����P��W��k�2E��)됏-�XqK�
�UFk�w
͍�KZ��W��z��>J�{ǰ�z�l���|YcQ�p��3;Iw[�ޱ#��=;X�oa�)a}zD��b"�d�l g�C�ŸH@3��6	�F_+�	��P��Iv�\L���[�n��������X,��J���M}~����݊З�?n��a�����t�Y]58|}�T:��]Us��BӼȠ�xm�+��4Y��E�K*�Ǳ���v�>���B2�����ذ��GU�p
V���I_O/Ƴ=t��'#+i�4O_WZ��������O�Qc�J�����A�'�
�6��Ç�lؼ�a:�Q���ߪoi��:O� ���ͩ�j.R� �)}Su�и��j\T�K��9�lo2�3�]ش W`o!{�B�`�`��]��v������y���.̛��h�D�j)j� P!�zZ�4󬍙9,�5Y5g
�ӊ�vcU�!+Z2&����IO�US1G'C�80*����,�Ѐ��yd)ʄ"���Tay�����2��.2�۩v��{��"�KV냇�xAaYw�
��|�S��J�{�	I�߂�^Wv�=��fz?��A�af�Y�%�S&��$ ���Z�c#8��6m�'����R�%��wzp�|��1��~��<r�e;28=�w��,�Akl����Uwo��tv;9�B����������5�9CE�>�<{6D���C�?����7q��T��V��f��ͪf�0����Xy�(<7:,�v#��S����*7�{��C��K�Xz����*@�S,	��jM�O"�eT�sw�-��p��*�]B=�|'m�Gm�d��_Lp���K�0���U:5�ME�enDrXDT[�/�S�o��L�u���;Jٞ����\05���3�	\Uu�Y߉���˳3j.F�lxRP-���C�'�ooi.�+��L�n��P1�@����k���g�ऽ���/rة��K�=,Yp��t��|'.��U�P�K^��N��$����=Ew��w�]%+\K��"�J��]3���ANY�����d&�����
[W���_�f�d�A�:=��<wj�}_\�*���zG����=ԏM�婪�W�F��P�o"�f!��<�`��J���L��* �Aü�ڙ��v{jg�B��Sx�J�>�,5ɚ���7��q+(n蓶� �Y�I˦بkm���Ccu���\۱Nj#�m�����,j�2�0jok󊹟�U*9ʥ�V%Y��hS��G�ӄ�}qx��#�ZlN�1������Bϣ�Pw��a�T�M�3��7`-b�S�kڑ&-�����Ej�=���x���n�U�/<�� �ٍfi=܁o�<X��3=�_�P#�<���<N�v��,u�e�_�Z��7v�R��eoh���9U��� �JY7�a�7\5�w�"�)G\�1��|bε�3ެZ�ϣ%LF�\�{�9�T�舴ut�q��c#������i�=n�?�".ə~^�������ŵ��1��ҭ,�G:B1��n.v�xT��U��^,e��Vr��9��8~���J�n*�a�(�N{�ۮ�bB�/�ɷMQ�^+.�hڹ��!�؈��R�X���;�����Eѹ��ͤ[���1$Ѻ=,�Pڰ4�{ɾ��
Z�́��d��&���s�	�J�7�e��V(��x��t����d�y�:��A��Eİkf��h��N��٭Sd
7u�����w��/o�L�\W[��4:���q�b�\J�Wp���`�ei�ig�^�l7�a�H�{���Kp����%DҠ�N���L���������z+�h�+i�D\�\@�<C��:���JdE ���("Lٔ�Vm��^S܀�C�����iR��-�&	�.�9�����SN:��"��M]�IU���:n��-�[²í�IҀ$��n��k;ؘڦ�T�ܺh���CJ
Ý��yЇ��Q��]�]Rn���nh-�b=�vh�CQh�n�2�v+��9�N
�ݕ˴;6QE&���s�nb��p�%g�����oj��tH�m�J;�]�͆�>�j�KT:"T#�ǺE\��7�գ4���,Wm�}�*Y,M����P8�����%�G�냁��];Ӕ�4�k2DU	A�3d;�:�)}�ɋ�h�&^��D�RE�Z�:���94<G+`jcM��+҅��x�:�zU���{`>�x\���u%�넧�>X�ˁ�$�	[2�a�fa��'�ʜ�����)S[R���}�2j�hc��K6o5v(ŉN������6�Ǩ�5���T�˼Ôuӧ�p=n���G6�(<C���IU�m*!k��8���&@�vt;�Yf�-�	�92�{z��X��Ґɗ��:��l�#M�֡�m�͚Ycycx��1@.b�}ՅJ]쓦�F�WV5��1�q�Q�#l��a���5h3t��Cw]�%iPι7/ �<����}OA�+����`�1�R�Hَ��YY����,L��wr��R���k�A�y��e��6� 6jtn��j@�ƹN�'�PV�B���՚�炲Y�هu�@��ʔ�c�D�Q53�͌d�	.bݾo^�Gt؅�!��9K{��.��f�H7������5t�)cģ�ԧmh:n_)���;-���dAtN��TB�I��F�uy������m�M���ZՐS�K��RE���ofu��ǈjY�c�ۺ�Ha��l�m�j��u�"VID�eƂS.��h��F������E�'��Zu,�w�����Lsq���KoL�7���8�1N.��'-��QE�r�c-[��:B^uL6Y���v�̡	��� ���(�t���&U���w\�Z�Z�&�t5/V�A�2Q����rV����_Y� IH� ��[˷4��ob�#��y�)�;�Մ����� ��gm��I|���1�'�l�.�+�����6�7J��O�4�3l�Mҵ00���P	gJn�]"^�\�-�	��)Cx���_�z�5�b~�)�{�C�E2(�z��V"Z��h�����������Jʬ­h�Q-YR[K������ER(b�J�,���-���ZV
��X()ec�T�B�
�[-k��\�
Dbŕ�Q�ڸ�d����5��D*�X4�#J�X)"�
�$PQTS�	��R*�(�"�Pm��E2�Kl�����PQF1`*�*�-�r�TW-E�ĵ�����aS(�T\J�ˉ�#DD�*#iZ5TV
��0�hڢ�
���Uea�fD�
��TUUR ��LL`T��UTa�*��a��r���E>Ӷ�FŴ[�^o,j���5���<�Ld� �ᘪ���=:�Nj��7rSV�@��z�jn��K?�@6u��Hr���]1�e~��1��Ǧe�;œFH����⩢~��V�jcw)�F�r|Gk�~�yop����#�ڔ)�!��J����\N}��[�s@�<b�����T��Z��3W\,��B�%܍v���lq��L��?�y}�5�)bۻKu�h��V����j�q��t�I���̬
��73;A����/9r�7�#۱F�ւ�yt z������D���L�1�8Zrp��ydv����;�����7*g��.L1�7]DlR�c�\�������z\�AK+�,�y�<��*�x+R���0�xY�.�+Q��2a[�X��BuD��/N�q�6�
#F]n�:)c��9�ʵ{�Y}A��"�p� ��'A��l+bu�{����j,a�<�_�J&&����`HXp��3�dC�n�0X� �bO��Cr�͎f�v�S}a�~�+-NO0޾��\=\cD˨H�[��7U,��1&���#�8x��2��������*�k���޻���L�[IWx�X��kn�,�MWy�9�e���&�_x\8.�.�N���7z�<��V�|�� �#�-�_pF_o&f���+,6�ӹ0�)���oL��P2)��N��"���y�x��ч:�:�4��Ͼ�놭d;�N����A��Lw	�1T�>5��c�x�<EiY��~�3�4��
Y.����e��w�[&�V����[y��ٴF9�(�b��:s�dBG�0&lFdgo=���X~��!�Vah�諄�Y�v�x:Ü@κ�F2}��(���L�+�ny])�x��]�#dW�*���yh.RQ��{��#I����ZW����>�&>�N�QE����hț1���k�>un;�6�U��.�\;�\�J�hO�~[�#I�+�63أ���јi���ʒ��V\c��v;�4_ʖ,��&�j �3�k��я9h���9{�^B��z�TY^*�LP<j9{�'-�����7��B*!ͻcLG�>4�
�z�Л��5ME���6�Z@�1:۠BE��[$u|WQܞ6c~�����������f����y(GS���P9�1?)�� s=d#R��¼j�!�G���Q֩�>��=���1xz#[��t��	b��v�w���!3��5S��W/��y�m˞cy�VrJ����s�"R�r��t1��הDN�N�� 2�N�͞�dU`�.١S�]N3E�3 2�k�6�Z�en�tSL�	��nR(rQݼ��ε�$1��1M�(�,�O-��wTM_.�d�A����؆��SFgR�}�|lb�f)�)R6=���\G���
�\���B�&q��*���D`sU�w.o�t����j)S�݋�cDrFx6����tu�� u7�ȫN��Pa�V>�sꩽ2n�<|��;���.��i<��a�q4/67LIΪq�]�b�J'�Ib�©��*o^��내x1������+ҝ�Ru7_x߽y_����늝7	��8D4)ڍC;��vM�$Y��ꭲќC8�z��1k)�d^����K���W��6�͹�a�6�Gv�[c�-7��d3S|�ZkE�V냨}���aYw�
��| �c���m�{�j�J�^�<'��`rʌg��4��<�e-�#,������s�y	�{����ݤ}4�x*�@��,}o]2m��wr9����v���@��δe�������~s�[\�OW�v`#a��x)1����csC�̡���=� HS2���d���)�Y]�A�U�M��w�(��a3�����ۖ�w1���i���G-����}z1�"�t����pTH��v'-0��>s'-�)Ec���@�<��.R/x�U.�]^of��.��$��+&�t�7f6u�Ɩ��ǒ�����?��G<2�����-ڐ8�M�����U�叻'�[˨Α+`��?�����8��[��
�=���4���&�x!	mUЭ��jǠ6~���w<1��x'{6*ܨ������%��\�6�Q*� o%�p�+���E��h'<��Y6=��&����P�Guq	�yk��'��`���1�ٯ�|��vW�WQ�<�aω��j�7%V��oGA�޸BC�N�-P0T*�+�ظW�!����$f�hB���F���Y��5�R	vqpO#����&�D�͗���'z ���i�Q�	J��Y�ڎk=:I2*Mm�EX�l}(��#�@�g�3�m+�8�I�HQ��Nnu̒�I���67� Ypf+N�}7LE[����F)�wJpU_r�71p�����Ql�9����UQ�w#u0)�2K�4�Y�6'X�Tb׫Q�Pu��`�97�ʮL�������*90�y��1i�}4��"u���pt��~��HWY^a�;���T�5�i����n/� �Q���U+���Z��åO�)�����)�N�,��v�*�־N�	ޱZ��ZOjI�8.����7�Wsv�v@#���Ş7�����-Ɠ:���7�����>\ų�*���ݬ��u	8#�fWA(�3�Vv��Y"�$�:��	��5��Eʻp�h��@�G�����çii_�zÜ��G���>�*4�����_��4(N *�U�L�l�����80u�2	B�W=�b�S\�,��:�@̑�6�ü��tD[:�\��l����n���_\U���R7I.�*Z�;�Ns[JHH��N*$��.k
�u�R8��?[�)�!�gt���q�&�':p\��\���A?����7R��ĸkÇTJ���G��[�:W���4S�k�>��`�m:Y�3��;�l�YO��o(���1��ǧ"*�
�� 8kF�ے��zy�u�t(����d���Pg���qIa�S����n�EQ��$�_AEH���w��.~V3Ct�تJ�2��_!1M����B�%��`h��(��BS_�!K+E
��C�_�t�X�߽e�`���]pQ���~��w����V��U�Ӫ��/�^NF맽4��j�1�mU��\Š�|b�EЕ�n���L�F�*:��L�1�8\''
�k՞�����0Jq��E޼@]�
���&9�]q3Ja��a��pC*9;C�ӗ��={0wUd���1{�Erk�� ��҅s�H)|�q^�L��st��2��h�b��'��+%��j�To�Z�6s��u���N��)��s�����v�iņQy��]ˁ���`m�P��^s\����)���f�ծ��3|�|>.�ů��z���_�@o��.�t�FC֭��|LgԺ�F"�f�7aL��8�귗{LhE��WF�Hn`�Ø�X����:�U����yb4}��yz���4/|z�]��d��Wz�8�H6���.���&x�|J��s���eԮ�zD�М�o9�W�S�Q�Pٵ˷d�!>�)UB��G�sdߌ�.y�g���z�j<��_�ab��L:�h�+ܕ�������N�ܞ:+O�֪��w�5[R�Gu[R��es�ϸ�5a��V�.U�+a�Pݨ�|��2���c�$՞;G�y�A�9��=;b��Do�����|bk��:c���
��U�(��ү� _O�}f�G�_��R���G��t�.���L:83a���5�Q���"(F��&hu*.g���m��(b��uK��<����o�k�c1�1����������Z�<7���������)B�/xn
X���E�����p�)��@�^�;ƶ��	�9���+dVO� ���R�b�N�;Zd�֋݄��4L��t ���x�w�Ucc��D	�C�ֈ#==��уz!�E�w�[�=��n���~�>�<���[��wu
޹J,�r�r��T`�j����G+����u�`�{`3L���bG�V��F'gX�Ww��W�W��:G�Tڹ���v���=�EY�U�
b��Q�\8E�ˍ��;KG9�xŘ�F���jy�(�P Vq���uG�
�A�I�q�5��F3�*�r��_N�g����}�g(o�{����!d����=��ǫ3���BϷ�>�#J.�:U]k��[*������ymo�'@(a#r����Z���xn	\c�u��*^y�n:ZlUg;a*hG����@X���E��[D����������B��G}�`f��l��8n�Bٸb�{V���R� ��e��" �7j��ڽe��{����'ҧ��f��=F�K���%1���#+����j@|\���+$���ckc��En&V�;� υ`a�꥿���p�\=>�n���"���V
���㾓p��K���l�B�Y�3�g�Y�1k)�q�X3_eBc��C~x��#&knrP]:�F�Ӱ1��M缴!N��#���+u����,+.����t�@����S�����ή��#1�IM�o��{<:u���}�=�����@UVFc�Ѡ4�U*����lݵ���nFF�J�I�c��U��xuL�u�����e<Xb1�݇a�l�֎�x"b�M���c6���r��-�AWpN�w��DSz��9qn���)�XhVw{��#�b�^�oFA��(��f�Ǚ�^�kW��_3xmExؔ�Y�[A���cNO=�2[�֒�Db�=Uj��mz��潼�K�jq�O�����r��%��'*����0�w��j��#���c��P9���N�}0�nCw�q��CE|������,����4��r�_�3� ��w
�eb�����aa��3!����)Ο�K������I���J5�ۈi� 9��y�%�*��|��G|��C�n�w���.T������<�E��g���5�?_Z�؁FY���Lp�X�Vwкȃ�DGWnK:��v
�}����(9��pu�,-R�c~��n>H�;+��09ʳ�������hC�֨��n��zV�*%:�9� E��H�P)�Q�7���b.��؉�m��˗U�g6�%�����T'�\M��L�����J��f�'�E�d����Hf"�bȓ�5[�4@�C��Ð9���Xk�5�C}Pŗ8�������2.n�{�_¡���'8���8<�Eb���e9���.���}ځw;�p
F���p�֖��0��z�TSy4|�M�����Ƕ{(0��Cq�ܝdBS�k�J��X�����6���J=������W�W�U��p!���Ҁ���4����1nHB;٘���ѕ��#�9�R\ZϒxY[�v>;�Qp�n��$�s�J�Dp�	�:�1��V�%e�ڥy^L�3z�-�/Jc���ѓ��cy�|�,f�=��l#8�����a�o��}�|n��j�2�"��Pb��%&���Y�LX���uY�pȗiÊ��KO(�Q��I�yp�{��혰��,���\���[���0�;HrR
��8c�
9bta"���9�\�8�r��1���j�@����[|y�&�s:!��L6��.���7��}�w�H+Bd��Լ�F�\N�Y9鎝T����ˎN�6��=ǯ6���F�)��f�jtd�����ϲ��Gqߥ�Jo�QW�Wm��ƴt�[�8rlў�Fr8��A='eG��S�����pX|j{�2��,��#��!�騪@O�;�Ü��4g���J:�٧�K��T����cK1�Zc��cmU�Tg)F�Q,$��+-Ԛ^F-
�Xw�@f�t޽Q�hu�pS
a�#3j^�\η΍e�3_M��z���@�g5�g 3�K���Fw[t��u}�%֬�Q�L}���Fp����r�MJ
�����M��N6(�q�C�a�lC��6l1�`����u�>����u�1��e:���R/rW�����u/K�΀О�C��a�(Ԋl񩧗'�׃rv�h�Ǳ���G��3L��Z�n	�.�q���w������V�\�Y����˞����7u�S�#`��` ��1"J��.!�n㶓8�f$��.��,�̛��Z�	��y�]td��,�S.HF��&9��1Ja��a���ɞ��3�VcrP|;�zzwI�{��%k�~��7
�<Od=+m�0R���5�7'�V��9V
'��x��T���H�P�1\	��@�a��ikc�*z�-w��Sr�������#��b�:��&��qB��� �
˰�b �hI�����(Al�N������Q(g۵q�O��c.�3in[�T�,���U
�m!��9n��saL^����k��A?%����h��~v?Y�k(���R�Q���r��Q:ܞ:t�x�X���n^�W�\�KF����(�A�41�)[�r�1Z��ve_!�R���W�O���wnVel�T[lь<|usUh��sh���BP�_��ڡ���O8��1�M��y�1�[��iD��V ���˥c��w[*��X&^/�^Ьʋ��h���U^�M�svs(r��1.=I�ǜ�srol�>�N7�9V[����@;=\>Q�y(E3E��e��H�C�2�5d<�5�;���X�uCm�=C2%ch�8�Θ�[��;�қ���m�����v�$$������c�Sg@1JF�f���T��i�b�'��e_@мW� �[�o�u�H�Z2�*��G]Y�T���	{$��ɻ��]��l�;��&����RW��\��S �Y�X#��X�&k�{�8��Nd��],]*�fyz쳾Ø=-�";~ǔ51�g;nύ�j�`����G�DѝVj��&��5���<��Ybi�ύ.l�|�sgVTΊ�,�m��rֽO3�\�/���X���ӊ�4h�w����{x��m�]#��z��/mJ�`A�ؕ��d78��Y6��](��9|����˗X6p1� E�ݬ_vT��JM�.���cY� k��j��1˦]v�2���Vgq�rbGYLu,��*8��?j��c��5��u�aO7��wa�`<����Ҽ�S���66�pu�*;J��0vF�A��^��pٓ��e,G5�UJXX�B�P;Aı�cj�x��$����|����V�Bݦ.�� �58�0Vѽyw�)S(��K�ż{J7�buuH�
ތ6$gu��&l���g��1U�N�����,Z$BLJ��O\�s"��f`��Y���z��g2�ㇷ���S��f���ne*�3*�bӮ�WĘ�I��F2uN	�և@N%�:%F��y)�ס�;E�@0����4�b�s\��[j�,4�Ӽ�K6��F�ƀ�HQ�\��:��ǒ��p�ՙG �]l@�%����ѳ��W�#��KrXkdH�J�Z��mm��o�«�h��R�p7��.j��'+�r��N�;C���[$��"���H��hM�PŶ��}ԕ�Z��H8s.���<�'��|�ދ����#q�b�t^YN�� 1�t�y۷��%���8��l|�`��G���d�b��ݴP9�P���f�~#��1�Y�gH��k0�DP��s�����G��K����^-��z�𳂱") ��d�Rȱ*Z��8Gn�۠��V��P�x��E��193p܋���&K���B�@ګ6���c�Xܨ�|W�7إ08�ͩp���U���o��:͔D4��������"�9�uӶ�(u�:�f}��&+V�c��u���j��ֹ��rhV��&IS�� �bK�emC�.K0Z�ަ��z��-����*�((�iF�UH���E&ZT**�X,Z�R����dr�"�dP���J��h���`�bb������Dj�+RJ0������#R��[P�i\�dJ�
ʹKi*��G).X�-�DFE-��%��W-b3*"!����K��+���ŎKq�(��R*�����TQX�2�b�[J�7(�r�q�\2Ķ�J����q�%F�ō�UJ�l)h*��`嬕+
��((�m��-[[X��2̎1�eŉJŊ���PXcX�XQe�[B9L1�"�
e1)�,j�*�[LV�EY*��q31XV�-B�b*R�D���bcm�b�c#i�c��*&- �J�~�DA�IpIYs#��}BF�D��v�3
����8X�	�:ڕSF�	�Ӹ�
ɺ��Uze3���}u�޸�wW�W�W�^��f�^�x�6?�l����F͖)�Av��p��a����0�DU��5��l�L��n[��=W�[T�V��
���e�v}�a�JCat5���W3�蒂�<9�b����O�[z}j���9�㏝G�wLj���d7��vhK��R/^��/1�:N��-	�Hl��P�R���o9zr5�f:Kt-,����]1��k:GXNƴ�T�h�P�G ��1yjb��Q�����6s�?!�^�# y\�*t��5&�9�)p�
�qw � oe;�PT��Ph8:��j'�Čhr:s�S"���=�.p�2�91���
Kg�H= ��s/�Ox�1U�^�.�RZ�׸�9�c��;�O�x�=����1] ��;�sPC�j;�W��Gk�fj�y������RR%����+�
�aˌ�]0:k2۱��ѻ>��"�ٸ����)b��+��y]t��]�o���-��P�T7�Ȩ��r������귧�|481p����G0*�@�Y�7�y@�=I����vt ���|�D�u�/�(�l�]b��C�����s.���5|nU��x
�W�&��ܩ&�-T��׻(⢯��#fo`�2Rݧ�R*ˆP�����uW'b��o�c~Ѡ�����ft2��9W��7��f[��_}_}U����N�ځo⾱n[#�T爺��>f|�Ɗ�-���=�Rf��g7iAf�#0�����	�'�>2�h��W����1k<S�+JL�+���f}~�`�����Y��cj.h��n�Ç�a����_���tmp������)�|�c5muܯOL==���mL���v����]?��m)�h�̆(���`�
�n�[�{�aY�*�δ�!^�<<{D�N5R�s���J9�Ѻ�#���Y���ݭ�]OQ���&�S��s
��n���,�":�}=k`�)sƢ�.��w�Z�/>�x \�}��� m�޼�}��mf�-!z��}_Y�F����!I�����|a��?f�P�U>�"�M��ޡ��"�w���(z��d�0��ل��ԝ���,,-����r�;�SD ����.�A�x���Ӟ�@--b�����%��9�~}��kh�aT��o�M������i�N_U����؄#o�̳�Ԉ�Mh�]x�d�(}�}�<��̖�.;�hMW�,�
�q��@t^�B�?�C�7}z�Í>AaG3 M��鬪�ڢ�%h.:T�ty��%�(:����L�ڭ�yB�]ey�^�,w�^'Hm\yT���\uUr��m�"�`�ۊ �.BN�Jy+�Wz���DD}�5N{�9NlY��U�E��Ϻ�a���Kv��b��|N
��|�å���m��x�j��u�X\��=�j�9�-��0��a�Jd7,�.3�g-�d�gu���ؐ���t�k�p�C�����Ҹ�3	�<���:�LS�"	˶�����5��ۜ��I��."gP`�c���p�@0��9J�\�����b���.M��l��y5t�w8��@+V��WP�r·(?���dv�E��GCl�2��S�`m$�8�ט��l�ÍS����>��d�R�ZrMhƛ�����΢��_Å�X��;=�/:875��̉�+�o�~�t�c���(�+��Oa!q͝����	�DА2w_gQ��'3{��x)G���ؓc��UR�N9�6a��)���:n�	N:��g�5Fעڣ��{����˳���j����T�뻨�m��PaQ�ƾ
�dRR��^�t�K0�}��A^Y�!�]-f�~Y�p�T�����m�;d��#��7p����+gαfP�K��U_vb��e7[n{/d �Q���<{��~S�h�|�s���:��Ь��,�(���wm��&���HC�ŷlr��0�r)�M�5f`F.�S��YL���A�� ��2Uv^A��`�%�Z��������}��3�O�Z�X�fR�C�<�·6���D#]}���0n�=6���w_����u� �=�SO����p�PV�.P�7�/���.�*�v_;~�k����dY+���9Z1����m�GvS�p&�c-���אcB�:�|k4�*�{�p�z��y��+��e�]q�2��y�q$UHqu���clpJ� d����i�̃{;2i@1^o]S{Ǧ-������B�%�tn���������Y�\�*��^o^��=�nY,1S���r�q{�.�(Ք��')dH�Ax+I�;��vro0��å�j@qj��0(�I��Tv����E���ݴ���D�:S6�����ɚn���{��*Bl���k���5V!Z�w���*�*��٨4p����[����m�)�*{�����[��������GO�˻�+��8d2�V�����¯z9/�B��+X�us����p�l�^� ��g��A��(�@L4�p7/���u�h�p�S�wPapPX�Z̳z>�rX�X���$)rŦ�uɨ�B�[�m��3J�/�e��f�"���K��-�,j��k���[b�-d�
=V�����&7�hY |mg�=�ǁ��iԓV�ڂ�w N1��Y�g��g)Y&��KC��tSR&}U_W���kӠk���U.ΓQ��*����	Q�6 t�b�5`4��
� �hI����_=sn��u��S��
ok�{�K�t������> `��n�*�W�c3�4�q�v�˭C`�Y��_�Y��xGS��k+�L�ܕ��l:�Ǯy=��>�oc��J^
�۞¼b���V}�,H��já�ڷ��U�+a�P�_!�Sqp]WP�A��5U*�7a�z��p�ba�^���q�!�����H�LU�/�vxY5�"���S'F�͡�7��-�r�����-�zb������sYEQ�%"DP�ɘL��2�iw|��q1�
z���Ǳ-����U��ϯx�
���R���[?v���+�q<����4�_�!}4��[�>ո���{��9�kn�3�)���]��'�j�,h��Wu���r�!���c�;�O?s���Xj�3��^����4�������6r4��i/��}C7'fz�Q;Y�P�x=^V��
�� 3g�чJ*��Z�#��:&P0��>Cݬ4�IH�3{*lB�,e#�Mt;��:q	�8c}h��Y����7������.���D�\��Fc��t���c�4f[v[��e$�{�x7S�Lz�r��^Qǝ+��c�σ�L�jԺ=2�ƫ��c;�;齎�u�DN��|�3���磌���
��
��enq�QӨ�?`��;��:(a��d���d��a��Xμ�=��r�w�FF�SxU{,}��<;����|Hƣ��%1�@�;a;��p�����\\���X���y����|3���Ԋ�X��<<Zw�,ypFřf8@�:�`�yJ�l�׏����X&$>�Y��Jݿ��(1:y_V	���T!�B�M�1������e�z�]�@fy_����}j�M}�itR1�"DZ�s��m��"�D�)��*�T3�Z�m|�
�&b�Oh,F��6[���)mn��W{ٙT���3΢����5ٜ-%�"t���S���z=lٔ0PG��6�z�<���1X�v�C���L���{�/,D��Z�C!�ێ�8m�Д����Oi�1�+�ʄ*�҆F�ԩ������sw��q�l
��Š-T�ȉ��/�\�\�\��X���#�}�d�W��p7ഞ^�3_LaQ����N/kl���u����R%�s9V�Q�W\4gϴW�,�:�.�5�|���w,woC4/��Y��E��]�m���o��^'i��؊sy�u�D���IoK�pf�&������N�����[�qߎu�D]���A�Q���h��Dۛ�3�t77��� ����ek���d�Kr�
�m"t�L��f�W�f1�����<�cu:z\i�^;��uR�!F�Z��ƺ��c&���{"6@�0K̠+]B�x��&o�V��1G�pj��f��IJͦ�$�(B)_�6
G��W��	�Gê����I1W�zL�����"�Q�\�jkr5�\���X�
f���>��,,o�!�/+��i��{�oMG6��ݼq��w��W���l.>b�����[˻�����M!�Y�����O��z���_|�nY�5��.�f�L����i�h�pY�NOR�-WٗS�M"Χ�kW�a0�6��*x_L�T�'��j���"���\J��N�~�m1r�ӳ��]�v����({���Y]�|�|_k��VL��K��i�K��weV�q�Dȗ�
�mC�j*��;/���S�^db���eS��2F�3z�Z�eL�뱝���ŧ�h�p�I��|��#+Y��ѓ6�w��R�:3�s��������7Ɣl�mV�.c������F�� u9ܚz7.�u��R��7,N�o�7�{�;�s�}��fђ�e����������ymX���YEy���s�{�X����ʈ9��k_a��rժ�|�b�o�T�=��娘��%h��e��j��k}g\^��ɉς�=����o�.�Mu`�G��蹺G�=S�_�'��z&�m��<f��N)��uu/t�'����V�W�B-L�ެ�p��V�k�[�m-6�����!{~�u�a}�Ք9�#���o>��~��F׏Hj�y��r�roÍ��k_�H]�-)ِ����p�q���^�8�ˌJ���ݽ�S]�p�>���^�P�R#��ϖ�4�����e�cB���O.-��\c��m��J�OQY���Mj�� }��%�t_�S���+�w3y>����Å�n/�����խ(͉���Y�Cy
�#^Kꓪ�z�mr���3���;cC+��<�;B�m.躮u�S��`�=4@�v��^�9a�n�1��:�Y�Z����ՎLBN����[���<���m�}�����*��n²�YX;9KQ�+tLݠ��}b����'U��wg*m����e��۹�����!֩������� ��t���a�]Ϟ�;��]	5�$A�B����{�l�t���s/v��1P��i{w�f$�ˠ^k8'	tE;Jx�]��?}\�ya�d��Om��Nn���e�2��ۈs���d;���E&8o�vT[VžZ6��'����Z��ܾZ��+JOdB��n1�j�����i�_g&j;��W*UF�;���$��mE�8�ή{IQuITڇ�];��7 [����`�l�V�R��-�}�^[ؼ{Q�A���5e��8⡮;=G��3tq����I\5㕸j⪟�5�Z�����/'*#��(��n���zo�Cj�����;�݋S����V�W�>R�^_y���s�]��;)pox��Ϋ�U��ih��~�9G*$_r��g{�K}]���F+|�n�)�{��چEsI�6�}Һ�q��^��,o\�놮�u�H��s���� ��M��P�]I�tA���%�
T�\i��[r�>75���{�Sۡ�<�K+����WS¯������zt!غ�*���o~���h���o�NuA	0jV3Pn�����$���>������z�pկ�}��5d�iOs��>�oW�{����q�����g@��s[���u�\_��:�DY�m&9�A��zt}^>j��\�F��d��l���fh����a@~Rz����&ړ��Z�����݇+]��js)��ɧ��y��Е|!(Q��.a.����Z:��}M��Y���S-�⳾�=K�8��G�1�LC�J��+��	.7�X��DQ��k�%ڹ2�7��m�7����
���Qn�Ҕz�.ڃѰwh�w��R�w���nCw{��4���;��\'��-�YᴪI��0"��I}�[[�������7�q�eD$��i[�
U����_��9�A2D'.����3���sX��O�W�3Ɏ����N�O3}u4��xe��w�:���y�C��\/���ޛE.Ҽ3���T}쯦\7u�[++��+S>C�
�]���>Yu(o\�|�S�ie]d͹���]��Des;��R��T.�k��6.B���U�7%f���T*�,T}�n��e�G��fC�s;:J}��)J���9T��aՀK�a�2'uÊ�Fh;2�J.6D��N#�*��1tۨ.)0졝���`�f�|�Q�-��D;j�J�q��Kv����pvL���W6�\�]�;vevۉt�q�����;K��z���X���#���Mn�m���;���\Y�����WV��8�$v!=������Y��&D�����3�a��?ĩ��U�EgM՝�����@�՞U+x�r�l
w.����|���cn�Cջ��Tַ���IYWp}���D!R�[��ka�������ؼ��n1lDzЋ���Of�q����X�DoX�>l`�r��|I��c�[��$r���
d^�YΕ$oM<�yk6V��t���l�ؐ�g����3��<
3�ֳ�.���d屇��M�ON��us��U1_^�`����:��4Eݔ�X_K�݁D��b�U�ubp����o��;�$\�qas��S/���9$bs��)bOjv:����/a�A7g��CͣD5]En܂��dC�sVNS����/Ѩ�=�B��՜MTh�\��L��e*�	p�U	·2�8�h�-8��Ŏ���-��@9NU�>�V���;k:v�4��*ں�a�ٜ'!+���d���E`v��ʕ�"�1�]��v���-����g��R&5駫-T�u���<�28u$�9�:ؽ�|�4ۨzٽ*J�/N ��ՃP��ҁ���U�A���q�EV�TE�����h�ޠ9�3&_8h�0�6�b�7]se���o[:M[n
��7x�$mŜ�u�s5"ۆu���|:������1�I�7����c�G�[�%�:�tFѠ�xd���hM�HK�-���m�g�N뷗N�7��$�|�Y�V��%�D�qY�=���7�8`�A��2~촰M)�<g ��&u� �b:�e__#� ]Nf�4eG*,5��YQ�x�ܼ��6tH>�g{���{��uth��H½x�:U�8����`���(�n�b��Db�Wm,�R�4�����z��c�;��V6��}��M	
�vf����+@��ܢk�^]*.��t�ٳO���/���_`[�]q�R�<6�3KYǻk8� �W[:񫓪z�yq.�6:|�=�G
A+�ؖ�'L�H��ӵ��oDe���3qmm̩Z�t�%���}��9v�:5s#���tw����r����S�V85\��5�;r�[�Ӣ��z7w+D5R�)�!	��!���M�"�1���k��,�>y����1�>�.t+/3-��J�}0/��%���� e큗��&�x߼u;\wS�7�DX�C���|���Q��;RD"�U��%��M*�wL���RT+R�*E���� ��hT�P�b�-��mT�J�,L�Ę�*R�QeeB��,q&eB�-K�0����� �ʩTV��Q�AG,�UFЬe��QR6ʊ����L*ԊV����ne��mim�Z5��F$Z�VE�J-j(4�crT@D��b)KE��6�ˆ+��T*X�kb�,XѱJ�H�X��-TA�Z��V�b6�n8�R��2��
Z[m�hV"���J+j����l�R�B����0U�ŖU�kH�V#PZYb��,��,��YV�
-�1*8�ԥ���+%kRU-�m�JŅJ�l�-���[j���W������Z�\nYb(�"�ҍ�����A���&0�Ե-��Q�-�6*�����QU�)kW�@
$�$��yfY�������o(�(�n7a�ʗ@�Ym�Agd,�)�o_�)��L�	a�|��.". 7ԣ����DDG�|��w���^����(�t\-Ѯ]A]���U���	���DM�5����x��.7��I�.�|2?c�5���7+��m�ZK�{�&��}d��;�=�ſ/R�T�VTG�f���Y�����WҮ�:�`϶ʕEJ���\���m:��L��K�wL�'����Z���B]�.�%��j8�q�Tck��?_R�����7��8z�n�WO�WN�f�M�Pd��sǌ~��5n��w���F,���5�_/?O5ώKM���]�þ�Q�N_c���dSs��j���BeOè�9�3��eq�S3Բ��t�F޶����wm���M�7�iB��Q���Y��L.jB��1.{�����ͤ���n�����Q��CWS����0����|o�5�5|����71��>���Ի��S�󂸇�����xO3�z��u�e+���J���Y\���
��3v�P�A��3�ro7�4���؎�h���� �pǞ���s'Ƙ�t�(ܫ�e�jM�3Թ�2�t7z#Eb���Z�ް��@��؄��or�K��rw%Ɲ��K\������dLv�R7��h�s�?��.̿��7�k�q��rk�55����U���<ot�a�A�6
	���`'���6E����l4�(އ�}���g5���:���Lp؂�(�ڶ�a��cڡ��١2�ෙʱ��+;|ت���n�&��)��`��v�3�.#���9�j���h2�.R�ԕ_6��G<�q`��ϊܕ\�n�sz*U�?�4�����ݙ��65h3��{��ʙZ᩺�1���Ku���5��kgs��T1_�	��ЬZ��k]YQ��+�f6T�������OF�������E[�"�:��Tn��|�'���]s{IحT��KK�Wpm��C���bv�T���6�w����9��:#�LV;7p��=�g1�$�<Ow!^�t����PU��PkZU�t��y��+)I��5��u�M�	o�2�mZ�3q(p^ƣzq����,�E]Yv��S����_4�=�ۅUq���̇k-:�<�ai^��%�,�2�9R��lcr��cc<3��7��p��=,�!-!ҽ� ��p�E��v�	̾�c���| �w��{�Oo�+�;M�J��k*mnC��]�y��8�L�Bg�y��@�:�s��8��?Sn��w�o�kwю:3^���l�P秼���#�g���՝�\�85��O>|�-�I�	6�6�n8����5�J���)/3��5{P����'�I��w���\��ř���J�ؔ�У�>�r��C���X��3��w�$�D�����S��v�!��lw�4�ױ�Щ��k��x,y�߮���N��'�T�eۥ�W��Xjuj��nwn�6�6�\C��p�s7�yP݉������4�+�wu���(�/v��%/k�7͛�8�3�BN�����Y*E��u��:�$T�g4R�v�1TE�3���{ЕHڨi�낮����E�S�22��o��_Kj��r�m�ی<��Gy�cf�ϑ�mw#�U=���4@r���^x�@�s3�����y�e��e\e�Ԋj��`M�}cs�N�Cj���oj)8yZ�}�{��U�ͳ��(^$��.�_f*��T���9�-D2X�t)�6�\�F�$Gm�!t�尹���}X/.��Zs-@�o�� �nsÌh>Wt�ج��K��u^�Vm����P*��\,ʻ�C]a��͞g���mΤ3�Lc�-ؼ�cr�/�����.s��Io*��Ɏ�Φ2�kq��1Ov}��������Cih��;l�4��VD����-'{�Ғ�1�%�s;[hy��ꆻ)����uܓ��6�:I.e�X*�/����k)Jqg|nw�����O[�ϝ��5؃���PQ7�;Y5/z�Q��.\N��y+K����5���X2�Ì=;T��{K����r�qn�F��Pttk*7�I���z�>s��3�6��I�i�v�X�4��J�BR67��s!.���������i����6���6��ƥQ�e)�'���}�>�"�m[�/Щ_?�dx�E�C��oZQm#_Az�������
�.;�m��WN��^q�j�& �JT|�1�-+͊NI�K;�.c%��3�81�8�H2���T�r�wB��2�'�`k1u���4�p�9D=��N���ј$f]���R�"�^�5�tlk���E{��+g�K/�0Z�e_n���K=��5���� �;������wty���_�]�,S�ˎ)�iu�:V��p�(�{4��f�0��wm��H��)k1�1L[�_b{��$����8j9���W���4D����uu0gc�9�<�O�g1k�W�ʂ�ʭ��fa^c��qܺ�s&ap�;/�D����x��.V%}��NUs�.�������a郔�8:���]l�����[��4��( ��-y�]�'{}�����w��bC!���eͼ̭cr���;q�<��츊���u"���X�u/k]Y�G�f���ڍw�m�5������V�Bϖg��<!������|�~�u.�
���<���׬����E˞�y��D��EsI���lOJ3{H^��8�}��k;mJ�Hj4���<��C�+\u��g��ErB`�lu�����<����ை�k�֋H������Y[O����ehݟg�V�[Wb�(�k�[�AYs�S�m�O��pօH��������Pc�̐��3ܸ�q�	ɓ�}�j�]���׎�nw ީ|�r�6d���X�=��%b�Z�-�}I(�G;+���}#��9S;77��p�Z���Xdʅ;�u�Q�T��+{�v[�̷�}_Co����wm�=�b+������AѼ<���2qKxtO�wNn�����u��Z�����m+�q۷��j�QǙWSqw�E��]�z5�#c�Ĺ�u�\���xb{���B����.b�wtkX�'�;���sk�(I���o��Ṉ�y�=�6�����zl E�3N���N)���~����I�U�;XO'�T��=w(o\e׷Ϡ�$�S�y�w�/��sO�j�4���9��Lh��4���ʭ�:쫠�ڇ8ߧ��^��zE�$�Sj#P��&c��������<<�WE�o�c�+��S���8���H�
���+�n�a���]#y�u0�[��{�=T=�j�^�+�[�f2�Ou�mI\.�����Q�f
^[D��M]��j?��]n�=E�ś;Hn��� ��6����v/S1��ަ�J-��*� ��dy)�(���ͺ����2���eN�]��u5�a}�}t�ߙ콎�N�\�r�.���.'���P�b�	��g��d�ﾏ�"��z����7V6��}���'ϥ�P�0~}B�ߓ���t�t�:/��Y}��=�k�L���zY�Ѿ�J���7�麺�������Γ��4��^�S���ޓݳ<��P�Z8ޞtmo�q��"��*_eN�`�s1�3z��lU���|̫wy�c���U��f����ϜVe�u�ܛ�$�Yl�Q�_Cm�ϝ����e�x\d1��������Z~�+��Q�ꬔ3�+WuΠ֧��ou��Q�º�XĻin�V�%�7'�n%�lt�����R�Q|�Z���'��&��8]��6�L���i)}]���}�ǽc��K$B�H��u`̝�������29S�989�N(���r�tm_8��s���)�;>��X"D%S�wS�圉׊�z��F�a�ɱ6��LӝN����b>�K{lV�h�/�z"`�n:��:�euU��I[�9��4:���L�w9�	�
��{9�2�_�մ���w.�]��MԳ5O�Λ*�ǔ�Wl�Sn$�xз|�V/+g��Q�C$������^V�9b���lmT������ gO��E���@�̸G��К�;M�l���f�g����bX���e�C�����{�ĥ���pV�*9_$��j\)�t�:V�U"C���Ċၖ�4���E�8����	m˸d)mC{��GUrή�����tNӀ���/Ms��1W�x��V�?e�Ie���+�Rr����Ӵ�Ԑ���-�wN��_{��Z��|�ſ.��Y䇈����m')>9�[i_Νb����M|��cp>�8���9�ȩ����Ӣe����#}�ѵ����v��6_f��չ��������`%X�3�=��R=uܼ��`�K��|��O�J�g�=�Sl���^���tv孵��3x��A�@Z�����^>w���L{�>]��I~�Z0�oԨK�}�Bu���%ki1Ϛ�kyRg��|+N\_�9K��#n���E72(fg4�׸���V�r�#��B�U���B���K�) }ިc��	�D|�A���W�X�w0�A��E�%p�}�;���'o�A�\ �r������2��޻��)���r�6k�����s��W����S���{��w�����֦��Ѿj'���t�/b��_���\4f[��O�-�����	�ǳ��+����K���oT���|-\9���k���'d�p�)�}��4�5�j��;���*�%0!p\�$�7V����ӭo�4O��q?-j�Z&�rW�9�_��v'�<Q�F�k�5-M"u]N�,�����SVX]�q�:M.g����N�T�� b\��9Ewvh�Y����ݔ=�տ)��d�p�D�1�zZ���sv\�v�s�{�m�R5���Ɗ��	[�x:i�X�;��ԙ��c�8�>2%��j���. �����F�Wט�����br�D��P{/
��YP$��m]�F�D=N'�d��<��
��㉹G̹�<��Xk�3�-�G�~O����n��������7�+Xܐ���T<��|x�ҥ�)��x��fM����ʳ5���MWO�\�*աufo�}+���K,��H*8�iY��H<s(�WKR+f|R�X%k\o{u���"�j���3�F�+���	`��'<ѷ�rs� ���z�Te/�{��o>�ѩ��7ނ��׺��r�c���ؘ�O��Z�k:l�S$F�*g%��:�oP�aeAv��U�şA���y�LMw\�K��_��t��z6��T�vW�Y�R�z+�D�W�'�ŗ�}n9SkubYr�C����p'��u�|�_F���w/3nEBgå����TY��^�)��H��z��J�}.�bW�����S]�z�v@�9ʊ���Goj�f�+����=��!>t5�\b��p��Ym��Bڅ
E^�51��ӣ��em'��Fu�;��s>���6�Ƹ�یq��7�w��Rn��{q���A{�!��P؅h���9�`\�h�/��mpM��8���G��)�}`���4Բ�C[Pa*�p���{S��.�=���OL̶��䐻�h�o!U�JQ�pWh���F�������Y��)�7��#Sx&��2��x�L�rL'��jp��uD� ���5(�aT���a��PY,��)R��5�M N�yN�.PQ	oܧ;��w���;H;�R�4��+���A�進K�R�Y|�=�Rm�;v�'��VXf�Rrj��i�"s&����mQ�����Y��@b�7HU+1�K�Ċ.9��[�:�:JŃ��.R�&�����ެv]�����d�q=�ٽ�-��OQK���N�,ɸDT�Mf�8�i��[���i$���Jڷu] ���&`��ٯ\�Sz�]5�78v�����`G,�� �7��/V
����[Y�:�a�]���^L��5��vN��k7�A;!ghVs���3��CXv�- ��]ʲ�&����s�r`�?R�׎��j+�z��L"(һ���)�}-\�b���6vփ9i�L㼰�!�'2L������ҷ�r�6�з���O��K�ti	�	�j��0���:,���)���x���)w�ص����w^ު�aY:ӥ�e��<�4N�-n�i��ng,�"웬�D*�B#���x�/:�m���G��N�m��+��{Hһ�#Y	J��"��/���s��H*�gb�c�W���Ѳ�9:�������J�Y��oB7i������T["b93B���  P�BŲF����V�ooGTi#����+�f�F�^ 3uqw��N��.0�[�3�!5o&�n+�+qC�/�E�Z��;��ӻ�F�P��R#Z\������jj7B�Y˫�Z�y3�W�-�wJ������T�}biְ?��/�2�:u��{��dZ��� �+-r#;-㮳B�+Ҍƌ�\8�ďh�u�\hT5r���];��ی��+c@�	u�qT4mк�ڙp������%J�'��D�t	�ō��0X��#Ѩ���G!/9�U��]�r�`�u��b�s���K'�he�c�t�%YzA��v	���6�FJ��9w�qBq�]�9�&�ט�*��3.�ˆ�
�[�8��Y`�Zkd��*#1�hNT�ٕ�c5����Ԋ�n�ɽ��+Jŏ����7�#*i!!NXޭ�z0d�vwL���e�k�]�+M(��CN��'���9D���K�Z�0�t��V��m���
KVp�)aʗ�!�t)�L4GB
�/.v�#;O�٢ܴ ���J���j�lHMla�Xe�Q�cz�b �ε���H�	bu�>5�;C�R�zd�͎�(��c9���P�g���21�Dc+aʙYx:��v������0�Gnq��"uv�4#�Y��@�Ԣ;�X�ֆfŷ	J�����}L�P�Â"4��%�	�L�[B�^������w~����=�����`���pqe�[|tFضo�
�v�x�j��ӗ�S�o�`8x�a�^Yn��9H�;���xL������3��a�4x������3X���}�)tHy�~�P )�Q�[Z'Ԣ�Q)EQP\j(��J"-��V6ŬF֕[A��R�Q����D�3
��+n8��n1f(��ED[lUQ`��±�ʨ���#l��m����ŀ�c-�kZ-�(�"(�%r�ХJ#X������Q�����)A��*�mk�H����-
���ڑ����5�mF����؍DQ
�0�U[ZW,�5����jQ"µR�E-��P�V�Z��YQLj+TĠ�#U�h��Z0R*,Q�U�Ym����V(��B�����ij[j
�	X�*U���)���ĵd���q��6TZR�"��R�G0�J�R�D�D*R�bԶѴ�Q�Z�E��*Q�����1F��EDm)j��3FۈV
*
��"ж2٘�Ŋ�EQU2�Em�j0m�#Z���Z*
0U+UjV1cE�Z�U�E�UU#T��1*QV�$(�PjJ���RŴ̔UP�TUTTT(�ʖ_�}�}�c}}�ߨ����K��J竦��Q�x�CYp9O��}K�ء+G<x��oHpͮ,���+�r@�(��b?�ﾬr�*���*�}|�Ri[�����:�����
+���Km���G�.��s,^��]ez�ᕕ�e$�Wͨ})�p����}�����ޔ݊Pz	�r��敓���9Pu�9
��Q<�Z�jU�%u������w��"���)q^O�c��(��mq/GC�O˷��uK�T�<�;�"��a�=[l��Kw��c=���Q�J%�\m�Ȕ;�BxT�w6���-�J�|�.;��4�n���!%y�c4˔���s'�1�օ}t�W��ݳ����Z8�ܞώ.*�Z���@Aݬݴ�v����cT�&����-�{Ǚ�Esh��Gj-��^SEF�t�����:�ʳ�\NW-*T^>�����7?B��n�ر�p��a���)�uS���s��e4j'��뉭��a�hkyc��6�m0�7n���g*8Z��Q�׫Y��y�Z:-�0�y���<�=�C�e`��ޙ��˫i^��+�& B�bn�[~ky0�Xݓ�8���MM{�n���^�ۋn�=���x9X|�����-ȶ��`̌j�]}�����Cv��f�g��_���}��]	��~@b�)/�]���gQ��U�5���OԞ�JU�Χ�2����Nv⥻6���)O��r_��%�%�-s˅��CN,qPs ���ϙ���-��(�NQ��ʸ��K"�g��\�q5��;j�zg��)�i<�3��t�	8����<b~K���5�S�X��\b��c�~��ѫ|�����rk��Sb����:��JY��h��ܧ9��I����k2���욌ow�����o�����Bu�lbKܙ y�&8D�w~�𗣢Ѽ�1�|�.�5��%E�RV�:9,��}c(u����:��z?O����6:=���9��/�ڴ����{yk�e�����J�E��مҨu����e�}1������0/"*~�>�6fjq�gVpG����Ԣbݧp���46qޚ��eG1�E�Q�oaԃT��8���:)�Wݪ\�T&`5fu�=Z5"��.�������t�۽C�?Jr��[6;�[>�,�^��Bz�48][�|5��}AЬ�MuGy��1��"�^�*�C�v'�Hm#˾{p���Vd7�{��.���J�rȗ����ow��E���ge�ЄX��z��s.���)��w�=��_}��s��&Wy8���z�j���LR�z.%�֩OFp����a���5�=.>��F)��p��к�\�:!kb�x����p)+��w1O"�e��;�/_1�[����*��ҝ�����c����^���^�ve����K�A�ܙǹ�fw^����o�zq����z{N��i9(ز�y����gͤ���S\��6��v5Ԩ?D��E�@�ݫpI�7�j�	|��q�4�'�k�����~��H�H��y<Dq.�اpo^ћ)H�x�`�K��&���V�ۺJ�_.����h�-����tu��O8˙�n��@|���m#���x�q���؋t܎q�3F�V��o;�zlہ�F9�W+^\a]��O��9�wp�7/Ê`5H��.�'�̤⇪��`����
n&2{v��I��r[��xg^m���]2佴�׻�A���R����.ȶM�F�m��z��0T����\��-���r�8,�a����f	VzXT��׷����&&v8��u�5�ƃ)��S�vM�a��_W�%��������൐�؟�1¾/�Jڱ���رȚP�0�O�,���7'����7s�Ӈȗ�X1������Ti���23��[���Ϻ�V1�o���#�ۿ����9��;��]}�]P��Z��_�K��#�=]�RO�H�E��b@�e������9ֆv��tk��c�w5������v3Z2*�y_۫Z���ʌQ��Oݖ�O���K����Ө�]�H�����1'O��v32�u�-Y/ڴd'��*�++ޡ�����:�F��U{�6t[^jޓqh�1��*���~ս�ޯm�m�D�l�W��~}�Ž�<�W��*�[U�C_�����8x�����T�Z��	�.�˨�\ci���'�W�pY�h<���4���x����/>��֫9\�YE�7�9����cSm�q���/�-kQG�v:u��s��ۅ���]H�v(�d��q�9�6mU���obҸ&�`h�S�����U0-ͬʓƥm.ɇ�$��Ir5R=�@��}�X*��bޡ[[�&_�LE�}&�3{���KKZd<�3��S�i�t��O� {�Gf�=����uc��\�_дt�O��i_�5eB�\Kڙ���oK��ܞ���y:@��ᐕD��>���Ի�AO��yj���s4�8[5�E���T�φLE:F��e_��0��]0��@]�qN�(V�*���
��h3hT�ý�h��D�����'�� )���S/(j�\>%;��j휪��+���o����&B���'����4�}�&��~��\Y1�;���F �qʿ��7���mCL��>co]�E͂�g�YNq�g�5�k2��E�3����9Pu�B������4��ԗy���w_+�.�[�v�kB�iK���~vȾ��[����P%���oW-U#�foa�nǡ�p׊Z�����j>}�V-�w�ߚ�e��H���t�^۝+��W����������F�}>���Q��
���iW����t�t�WNx���88�:gG֥JM-/���Y�9� ]���oܟJo+�K�}��;DL���qWl��b.m���yDgU��%Xr�F���,���ia={�N��u�T���T�[���6���j��jL�:��V{p�X�{o��)�z����n�Il�u_�8�gS�f[z���{�v����{��bR���A�j>c�ݨN���J��C\�&���{��v��[o�u}v;�ʁ-��F�A�����o��7ò��������X�^���L��p�����Z[�bx�����|8^/*��uc�t��>��>���������x�H�r��&{�!f�����R�R�|�Z���'��D͝#o7�=~6}8�.��M��-���N�u�(q�ܔH
��b��MJ�z0�ª&��-�Ci>��u^8ɇ�b{�0(I���2�g�Y/�w�,-�׌oe�-n��F�Χ@y��1���(�r����A���D����K:���{VX]��_jk��UK�g����׼��/f�i���,>{�ۑZӕ�rk����T�O�ݿ��r3������n�a�14�0c}y�i7ա��,�����$.��Nȍc�r��;(4w�F�M��N�փ��߲T�+6��.��Č��H�Qo̼�~c����f�XkhTs��L�� 
T7�z"��Iy]u)�=>!pW;��`����ڰ�;�3�ca�����ݲqC28���R�)�5:��[H�;��c6b|�<��(�ڈ�Ϋzgy1;�Ē׮�tsڞ��!5{el�S^�����?C@u���k�媷��AM�x�:*��m(-s!G|�d�V;�ߚY��������C��&-3 ��B�z�y�k�(W�7�~s���bWmG��|.c��\�n�Ԫ�S�Z�:�]]H?R�{LŴ����N��^�.��f���V����@�%U�:�u��	8���J���c�Q��u;܍M���{�����S��~w<���"$��)�DܛC���w��7��t8~Y5;�gؖ��k�c����&�G�k�����lG�W!�Bgä�X�ȉ�y�{�*�Qu+:r���$VJ���ᩭ�|���KO{E:�pG���
�՘bg�NQ�� ��l��uwN��m��,p�9���o�.���o�wzݤ5���[����$M,e>�g]�dkae�4����A��]�6���T�X�2�^�$�c�Ȓ�����E��ì@��ˏ+��K@�<����9f�a'���T��7�4�D�����yʕs�M��$��N�Id��U}�u��v�y<n�@��Qx�܈��]���J���s���R����a������ ���W�]����=�k���k���wZ����sw�<Φcem�;n'v;���!�����쯌s��bV�������[�v��.J��c��UP��ܭ�X�鰛OaXÖ�>=L���S�7�d��3��ܽ��ՙ�iY��u��.3z�����q�݁I�������goww}��<�əqݻM흴��7����uK���fv�s��7��C.���n��sպ��$g;��[��v�椧�l'���u�Z�u>��Qr]�⧽k��|}5�dw�OQ_e���n����\m��r�vbm��2��mL�����B����V-�Խ�uO��i�OW��r�ji\�.�s�W"�ך�6�_>��Q�����]Y'1��2+G�.�*�d��MI�_x�*�w{̃V�ܬ�[s+Bz�T�TO4��5�E�Y8�VL�G������gjF4�f�]9��`�{�iP�#34	a�O��[jv[��:�n�Xf�����.��4]z�ܒ�j���V,�j�J<�{��S��U^>����4lce��1��*�k��J�@OcP�j�'�t'$s̺�����m��z�n;��K�ݸ�W��C�6!U��5Ѹ���A�Ng��\��'t�w1�m��󷨪Y��f.���{R����A���Z�����K�+���w6�sW�;�5�i4���5X1֗�1C+I�)�T��`�h�"Ewm?w�_�k�s�{ޒ��9��9�[5%=����3]�.-V��6ʿ�%#a#�9�t����f��K93��Y3�$͚�;��3�7�� �/8_������/�%�Mw��p���	��bmަj�w�y��=����NJ�`���A�dC�����Zl5kk\�w ;��L�m�6�S,�-�}�ѐR×B��n�\�lM�{	,��"��<{qVRTm�x7�u{g)^�KъQl�Zj܃��<%]�"��{�6���9����XՊS����e�5c�_4x�dE�lt�u�j�f[�+m�8���5b�m^W+��[Mӣ�����Acs�M}��黍�&�ֺ�U�U���}T�����LV��T�u�f^��m�K.�sg �n]n-�f;-^7W"3�f�j.^��:Z>�ѽ6���/N,>������|�OOY���6�3x�Դ���P�
�)L�����uQ^o�êG�*C�|�����E�X��ܘ�9�0=�-{�;���[(tZ�Ь[��1�u$��f^wSc�KTz�5�g�K4��S��Y��-���-gخ�M�����L��׻~�pd~�Q�ا��s�������6��`T6J�W�c0�=�b�t�N���s����Qʎ��M��Z�|�uCKj��=��K$���u��:T�u�.d�9=NW-*Wk/��[�;{\�35u��{ғ{�Т�xf���}�XP��{�[�r���u�&��J�!��uX���z��Nǲ�X�����7���\/��Z;�Ů�s����ʫa�O�,�F�s�k�c��Cэ�{l%p!)�l%_K�����.�!f�XMwF;40��ҽ�&�a��k^�����C���E� �zZ�D��("EqΚ��fV��txe(`i����mG8���,-ˇݸ��^tQ��Ւ";q�Q��,�)w�a]uض�
頛�4�Xi��8n� �T��)0��<�W{���q+t�����[��Ϊ�џc%�E��B�|h�%K�f�'�2mAO;@�xm5~�.��c��yC�ϖA�x�V�5D`���/�0z��g��Yis^Mh7P�m?�Y1��*8��Ǹ�U�G�ɦ�s�G0�A<`�:b��Ƕ(*kCoZ��>�/9 ]�t0f�L+j�b�n��L����
`]mWN���E/��bPn�R��4`�e�:@_@�j�����r�� x*�j[��-ǜh�Nu*�e#����0jd�0�t�#�pgo8�7AN�]�{�۶@vj�aQH'9�8-mEM:R�ƶ�<�Ԭ\3l0+k"�ӂ��CXv-�vg}k��k�`�ԎS�;����Ϭr���u:��t�B����=�EiJ�_;�AGB�Q$�X�x5�8�6E4p�|��eY�fPOsLʷ7{{r�򚕈�Wɰ݇�����]���U�P�, ��:�t��f�4־O�诨ܢ-s�[R��i
��7.V���{��X/u
J��fh�I���ڭt�n�3�+8Nz�9����MP�{.n=��Y�G�I� qN�7������t�E��7�];k����[j]n��3��V��7���m����nV��ʼmVi*�8Q5ԙ�&L���^� �`7d4��zf49,/0�s1���)=�נ���;
��7#T[�%�Y�2��/7[���5�ObLR8��M{cv�D+�2P���6�m)m����k�� jD7�x&x���u Y��71뛍�5�����=�l�nV�4s;zEt��6TY[;�d��;��QF�����Y(՚�q5u:�1�q�]���!z,t>�E�ov�Ep�"�Ky����HȈ�o(�r��I=������|w���p|�'��L:�l0�P��N�	��ˡb�c<�v��&��0=
�ń��[weu�{�-��1:�P�m���>z�nҋH�d\ʵ�%�'�i���'q��z#Z2���3�U!t��3{
4iwѱ�J�[v���!�\v�-qr���S�Re�����]e<��cɺ��6����WeZn��b������n-w}�k�[�eډu�E,`|.�ūި7`�{ܠ�4���Hf�hށ��3Yx'N1�+�r�%��u���z�a)S� �,�YnKi���FY�w���So�.�� Ӽ��5��먖��d֘m^ژ��y�]��J��GɐY�����6s8�Me��D��T�ڶ0��
�	��-Ŗ�0v˒Z�I;���=tyy#��4 ��'s�z�d��i����X�4�3 ��;(�T)Db#*ڊ��TEUDVڢ�E��F�R��1U`ֈ��Җʢ�Z�Zƥ�4AY��[�$D�V�b2�%��c��+���
��R������(�Qm(�"[J�F����*1c��b(����E)h���Db��1U��D*����V1QQEX,eh����DF�"� ��"5*#Z�V �����ň��5�T����hc�ƍ����LJ�[iJ
���J����V�"�(�U�Q��j�*"�ڊ��H�Ҩ�PX����+-*�U�ER��T1��E��
���TYPF ��(�0�TQ�EDAA���1V���`��+VZX(�BҖ�Ee�ڃ-(*�*Q*�j��m
��""1H��UX"��QEDQ�)YU6��TU�+���1�,Z�1�F0Vբ��Ue�8�R�(*�V�X�m�-�iZR""��EV�ҍ��D��������}5+��]VR�GvC�}��#��i9-M0�`Ӻ�Zq��b�٫�4fSa�lS��׺iv�!'Xf����Pl�����8��+�-
b�Jn�n5+qn)�5��Wu���Wr6�����u�>o�}#�M��7��ڶ��s����LZ�bb��YE>��nH��J�*�Zy�h�I·+VC�
�ܚ놩[���9Q�ppص9"�cA"����8TA}��l�Y=����#8����@����1�n,����o;ی�
nD`O&xW�݌5�g;��2g������Wz3S���㫠��'i�P��Ah^�tsZ6{~)v�栐�;���j��B���/�@O]��*�{k�]+����,��-`�U�@�����X�3w���6�^������7i�.��Ƴ��%=l�������J�˷�P�w㋭�q��r�n�a]w�k��r�9Y���|�(:n�7C��m^�o��C��]e�+Ũ��:��kb��{��5;��*VlC��kx77��Ѻ��7]-�*wa=��A��4��v�K,��<Ç>6�hfz�N۝��V!�_Dӣ{5#ol�oV3h��?kꇀ}��ڿKW�*Y�׫x��g����;�B��3u�a�H�}}wYˋ�rަ7s#�r�`Y��Ϣ��ܛC���#7����8��d�͚J*�ne5�+a57�����h�rov@킻�P��0,��WAb��i���zO5;�Lkyx�.t��)��Z�vA��R�v=�]��-�\oݷ2�Nwx��7��pO4�������'_q���r���;MĜ��}6���ϭν��܏:��i�� ��c<1�rK�N�/iȓ7����ɕ:�j�ܮ��s�κ����竪y�F��{�&��g�[+:
�4�e�}�c��p1+^_�vg�K�o�:�}v�2+���[��8�<�֞B���Y�v�[1L[�X��V����+Q��rS�b��{�z�5SP�������Ɗ���*�/����_�*�\�D{�Wf�跔����j�t�0��v��Dh��fb_Y�_�$*���kɤ�Z�%����h\dVs��e�'/�m�N���0��]��*R��7�)�l<���n�ia@�<�݃��j8�+��u�)45bӱD(&`}���m;�IS��F6��\���[�
���6��ŀ�ju��ĵE[n��:�� ���Ύ�O�z��FS݂���k���_^NV&娟�����"37�7.�% ���uL�/���`��r[��c�{`槨o6�o0_j6���84��T��5�=�ު��*?v�hZ���[� �a]ͯ]Z�r�)����n).�;w�퍮��EXډ�1+�jHȽ'�\�ZJ���r�;��r�7����o�3��J��9���^����H�:{�e*���^ʥcˆ�N]�t�嵁si�'Sհ{���Ke�J��S�zD�B��Y/y�q��(���M�i�;ņu�굸H�����ЦFF���ݢ��X�wR{_si�q=.���0KL�+Sѓn1FO��w��P������fU\�ߏOU��>9�P��Ul��U��-��q��#�Sq�<߲'�[���e,��i�0�=���{�I�����&������ݻ�B��(���i�")�4�CO��3	�]��\���#W�7ǒ�#5�k��z�L���׳"[���Z�$t7��R���A6�̬�X���U�w>�I��ލkq����+�vI��ّ��
���͋�B�-��w7��������c���[���WmA��Onc�!�
)�r�rR��6:�m�5fX圝�7��<�l������׈��DzLn�s̷�o�جda���G��`]���3�r�!�򊺇�O� ^S~��w�U��e[y}�oL�[3ڝG*��Y�U;�/�j5���y�&�Zۧa��am�ǝ],�ǵ�A�c����em�D�מ-�vTi>�}/�ML���h��p��v���ӆ�"�=6�wg�a����靵`N�C%�I��h7����M�!���tJ��V�ϫܜ~��>>��M�޵ǔ���7�sV��9� K�Ӈ��r�����Jg��T/�(K\�&��'���[�ny6�,~��V�]��=�VkF9�ocR�q�Q��}�a��iޖ��V;�E�2��̵w�q������L��s�����2�X��3n��* �݁p/Q�2-G���l\j��˹y0LP�[O�K��c:��{2����[�m!�9��܆�xi���is�/��g����2����Z�tÝ��S� ��wk���*Y}��zN������s[g3p�_=����g���͝/o���J��d��1W�����L��I�́o;��ڞ��=�������9��`�|�aܦ9��ɧ�CC5ӑ�nkǣ��	�O����c�ߩҤ�ʱ	n��NL]�w:��|.��1����<�����pI�S�9�O'��w^c�������|!��+^Xۺ�ι5��q�����B����VNل��e8x�T��f��!M��̞� ��鑯V�kR�S����\II�	/A�f�~|6tak*-�Θ�xf-c�]F�'f�����=�7,u8�FbeWͨ}pUӿ��%�믊ܣ\��C�N9�i����[u	�����`�+�-F�cC9k�]�p��G)k�u;�F^u�vkq��gTD��.�c�����Ud��*U0���/.֔�<k!��:��d߲t%ݜ%�I�_-[�1h+|�f䃻\#��S���_Mgϕ���>��v	�v�.G��v�{�˸��������A{=��l���������X�IH<�Gu7p���CCg���X����5vڻ�R�k�F�;CR+���x���b�{�;q0��`n���9ެ��^=�]��;7�ʅ�T�~������:��ǧ��~��h��f��|��J��Q/}�Ϣ��D�ʾ�ByQ{6�^��̡-�^�v�=�u!|2og%��ە�=!���*�	},����cՇ��������q=}n�/�s
N�_N�K��S�͏��:��-��t���s���1�Yߵ��w�M&�;(��^�p9��qۗ��M����0I�K˸Q|e^biЕԻՏ2��������w����n-
u2Xw<D�S<����0����*�5!)����s��oLE.�E5��3�9~���ۡk�c��]���J+V0�V	Ak�r�s�L�n��`���'6͉ZQ='�e��kv���{p)�o@aO�e�V*�����e���R���]��Da�w}�4��1ZS˚����lXth��7:uI�N�]ەskU���=��$�^�{12��a8�����eOl@��_�5�%k�]w��3f��}*�n�͖���X�����9;��a�)(���L��t5w�%�5��������*㛠3�Lp�;rg�x;n������~p��Q�g�)�yo�:�Ͻ�q�I� J�;+��;s�8Ȭ��԰��c�9����U���{ޖړ�������v��(�D�OA��{{�<�p6�nQ��/*�TL�P{��䩡_}�NN��E�ڮ�{�)eѨ�����aߏ8P*�,�FR�\/*�ǞY�Rp[}^M����=/�&Vs��2��1����R]å���w|\�&2�.��[�T]������5�%mS7�q��d��9�H�.������������97O�U��v(}���s��+�Wf��*��5A�u����N'�g�w[O+$T�ZIw�9���ͷP*;����U3�F��ֻ�����β��ϣ��l����
����H����S1��:�onʆh(a��p�\�4�÷Ag{�U	t�Dea��r8e>��os)++��K�v���E�벹iR��Z��������.h2*/32zrq��K�<�c�%��(r��5<���v��=k��|{Ճ=��긮�U����X����+ѵ�/�a\nB�Th�����R�&���_t�"���2l���N2i�F*׺jq��^�|���k|���z�-NQ9M�%7^�z��-c�}��B��o�V�)M�A���뉸�;H�(s9����n��ޯ� ��L}}T+E(��K�'![�V����R�燠h�>�*��y����~*�x�r=�Wh���eʒ.!C,d�gAZ~�
Y'Uì� ��:/pR��~��zUz`{'�3�N@W�e�h����W�}ѝr7Ƴ��LV�r��&���x�bu��HO�"�ȿW��i�����G{·�#�f����,������� ��$)��#�7P��+t¼�t�=+i����.��5y{EGy���x��w���~˱�	#��=q�]�o�-�����= �|��
-Z�u�uR�m27�V�w{����k�9��)k�V��J8�J藭�"�⟑<����Yʹ��X9K���!���I77N������1K�mZ��,5Qm��n����|29-�9c|{g-�4�"��G�3�i���;AN��Z��>�P�[�y������e��L��^�X/�%��ai��c/=P���g�v�[zz��t�u]^ys�B>�7�����/��Q�q�:j5�\M�{gJM��s����tԾn������������O�����,�\���g����V�Jͣ����6V��y2���A�}&������,o�3�7���yުiי!�a���Y�� G�'��5��`��ϫSh�)	X? !ݯ^Q���Vc�����.�?����#X�f�þ#b}^���}��������/\��������,wM�Bk�qQg�V��7���m��NՎ����VZ�_���ZsŅ�����Z�nK;�@��r(�&"����	�q�+�� g.g��m��ꂏ����M���Heq�����nK. z@KHn�9#	]��Vtӱ�9;��A��}D*����ש�ӝ|��#׭�?\�>��g�������Itzx�}10�]u�9O3���\g��>��c���ҼHŔ�4�^�UX��6��{��wk�Ut�ض	�3�����Тf꣼Fm)u�V`�����aJ�c�HA��xGg�����Bx�M��ո3-���&p��x�r?9�P�^��k��ksc���ن`=IwB�S$�]���/Z��/��\���¢�H��t��}>û3�v
�N���{��(���x���}�;0�Q[�}��<�@��"�>5���g�&a��Ӵp?��5϶6f�O]y���T�u����\��p��X��X�3��T�ng�m�f�y�
�;&��.�Q>�c��.=�j��7I�;5�8��?X�}�n��=���̀��2�q��C�,�V~���ճ����t�iCL�b�_���G�<��\{��컇�����/O�������߷����|9�=���co'���'Ei��>���BK=�������u�*	T��QySr��y:\�uW����/M��;q�g�P��֛� o�������K����H��ۤ�_��w�
��/��ݢ�P9g"K�f�&7��T�� c��T%��������:��{��~�w��~�:�ΐ�~���2J 1Gg(���XN�]W��~.(g܀���eUE��v��{��+�=�*�^��z�*�d	Te��X���")?z��O�;f��]+��v�_s�)S�P�����
�A��h�4(����LY�t��p��;.)�����V�B���N�b挋�%gd��J�����1q��P��Y��k��U�L�V�����ٝg9�z�� oҟ;^ۓ��N���]ci�p��5)���_fp�*�ۏ{�i�K[�8�NnNn��D�QT�����C�I����!/1���[�f��/�r�,���xN���jx w/ϡ��;�J{Zݛ���#0v���w9(��+�����7wn����c'n�r+J��T�a>5��V־�Qs�Ȝs�w�0�t���NdώF��c��ʕ�-L�7X��8ث� ]��v��X�42��JP��Ai*�h�"fٸ�������.�N<�8=�ԟu�sNP_4dwӸ(��K���㷎�!����8JV;F
��ub��,�E��JcR����C*IF�*:���Y2^�wy6���&��D�t�3���
�8��h�C,�[E�ZI:w�zf��q�v���.��ʘ�sm(�(����fU��l��^�6�����E���LV�1ٮ�B!�c�@/��{���w3E>}�Pm��Xx\NP]%ǩ���^t(���`��t�n��|ދ:�h�y�����ӈ��g=��
b�Rk�K��gH��[��]�q��Y��蛪�e�\�]��o�*���\�x�V֗vpNT���q��.p���C���k�tC\��4�=��n�u(��Hin�X�7E$��X�hQ#��:_.�n����	J�E��%�4@�5���<������R�n����Y��T�V(�iܟ^�bͅcٟcG�/H��Μ̵��{�+��yt�q��J�`h��P�=�]f]��!Ƕ��Cqa���� �"�ղB6�������*>�1���vMe&^��;Z�ޮV��|O�ߒu7e�#֥ؿ�+	L�R�`K��N��ee(mc!�!Y�]5�f��:P*���ͣPJY�mc"=�Q	�njV�D{h��6�]�lz�8���j�'R#Kw*�<D�rNM�U׷�j�k�FۡJ���7ܠ��޸^�ِ�*���h�4%Z�0��&�����z�c�JC��Ԗ'Gz^��3��a9��N��(X�����~=X��s�!�b1�!d��5n]:t$�"�7S�T��_[;�-vv�*��m�0�������zX���K��ۙك���KŤ�u�{3�6�438�t�>�$7A� ��E*�f뾂N�z��J�]^��X�Cs�YA��fC�u�5��VB��oE�U�H��Gf�E����v%$���z �04"'^������I�ď\�"gz.-^Ë+!J3W-���GM��`���V���2�gVa"�tH��p�D�YX�$Nv3'Y��v1�+�a�8I3d�w��;%�FY/#�/i+��c$m�m����B�"�����֣��DU�J1ej1�ܢ�)e���J�UQP��b�+,[T�iTX*"�D��YR��E�KT�F%J�T������Ɗ�UX�Q���e�U`�1E�Tm*����¢��V���
�U��U+V �e�J��VU��*�m�*)QH�UX**������"��)����EX�YmQm�r�!�Ķ�ʨܱ��ƈ"��1b�)m�F-��1Q�*Vڊ(��S���1U�,�Eb���F�j���9K�ȬAq��DUT�TPQDDE[hV����s1X��-��TR[Z�m�ĶU����D*R�J�ETb�$P �+Q����eAH�[Z�iF"���*�b�fb�Q���X#1(��U+n8ccX���8�`��mH�-J�Qm(���e�EԶ�X�j[�*	\r �e�EF��D��)R���,���
�j���
�@���1T�t����y�����Ցs��/4Q�c�5��˭]��F�5q��)o1�`�����Kx�sn+�b��j�Y}��#����Qu��
�zJ�c��Ys㐽1��o��Ͻ�^-{$�P�ž��\9x�=�5B��+�ً�%�w�~{�\��&��-���?Z�����Wi�~���Y�{�������e�;�-XJ_��G^��n��F=�A��[�z� �D�a�Ykl���K؅����g���ݜ�3D��*W��]�"}�z�!����<��_A0�|�Q��*��-f>�Un�23��>��{�+):�6��m{������~�#!z��,5=q2�S���	h��nf�:%h���fǢ���^��ǥ+~;e����g��n�Q2�a�����G�rr�� LHWeU֜0�����u���}��Oƣ��W~9�Ǒ�y@+�{,�_E��Rnf8gNw�,"�e�wB}��Z��u�}�F��k��)cS�Q��znb�=�c�v$Ǥ5D�������8+Mm�F�M��N��I�=q7Q���`��K�[θ��=IՏ�����r'g{T��$@�ޚɇدj�	/��")��7%�۝�^���1_^O��>r�Y��y� @����"�K���߻�d�.6�n	��Y��0Ⳋ��٦$��!�#�pT쌾�NW�=2N�qq���l�S%%�����n����5�c���(���+��	�T����T�:�5r��*�S%��&iV�۱��W]�k�cq��s0��Nu��/����#k�繂��'�zO%���纡^mV����r��Q#��s��n��P�t����,��WMo��E�h�
�ӄ�~*vX��ۄ�ddt/X�6.秺{�5�>�:����X�]��>ӌ�����⸫�m�7�N����ziVi�y�̣�a5�>��e�q�zu�Nr'�V7~��o����{خym�|�>��踼5���������%�����z�{ŋ'�r��u;��ϙў�����+�A����{���%=�$W���u��Д&�q�[�Ryf�e��?(s^��<���B��8�<*wz��^y�G���<��*Pc�S��6C���;�P��7H��+��ꂈݭ�/;�Lg�]t�Jp��I��;V���_{���ȅ9E� 7<O ��zhQn�7�Bܻ�5N������~�4��"|o��*9�R*=>�Ǚ߽�:*�~��'� mɀ��!(���U����u�<���s i�]^��w~���ӼJ9��#K���Y���%���V/x"����J%�ٹ�)|�,��v����r�֍�O�*4��n6�δ���w�@<y^�N(���H��yJ��Q����U�!l�X��r����`h��k���+.�Z���9nM��Qڂd��ـ�+�s�Cd�l#�A�7��ߐC�ۄ���x�`?�Ӹ�6���-�S�����u���D���罹�z�����s#�}�Ģo�)���u�x��j����|;�!cn�����_��n/z&w1�k�h��UG9^�s�u8�{,��L�����;�g��֗��m_�	巑�gw��M�sP]�H����>��ɻ��p_�"��ヂ9������i7��I��<σ�1�}4��� �T9�g�k��n�/�#ΪYG>�<_��=�3�8n;�Qˉ�����J�[�����ܿe��}ûfp����L�`r��G���Q8�}���Uĵ&�'0���|�'��,�ε�j�;�>н���e�MiW>�|FzwR�����>�,W����,�?M���Y��gֹh7��=�'�o�>��Led֖/&w���t���ك�ϼH��:��>���n���~���;^�V��F�絨��`�������*�7&u�U}��w��7�Sȇ���	埭+*ت�Ti�Dw�6{~�W�9�C��xr�����Sq5	��ÿ�S/W�~�)6w����&�-�<���('���S�e���e�Q�G�y���<�F��(Ljw��$"��TL|8`MO�w7����WH�P�V�]C���L '�,y���k��H��X�ɼ�!��:"o0b�]�`"�b���;A�0�/g0vf�R9L�B���q��~��2��/���իb�Uz����;ӱE��Z��S���kP��f�9`^�}�E߶�J6��ǲ�6w�3�W��|n=Y���9E� ��7��/�Ω�.�`�6s�t�H��L����;���Um_	O�ه���x��=~�p��o�o�;'6zj`v8�K�S�G����똘���WB�%x�9��x���Лu]⇽���5�������b��3ہ���v���[����-�����D��>�iωkgP,y?Se	V�A���]:E��	���}��{k�Y������
�^6�%��2�W�1?S��7�i~=�u���P�Ou�Ӛ�����3��|}�ݐ�� ��Y��T�o��f�Fm�׳�w�܋\�g�O��ito�_n�F��>�=����=䓾s��r&|���{���-G{�&d�'��尿���Ưi(��X��ݻ؇���:��m�{ =��ߠr��Mo��%�N�w�~��C��Ӵ�����:'�k���^���dxg�u�>rt�r���@�Oc|���4��P��Zj�J�h�}��~�,<���V0c1��l�"���cO;z�n�J��X������ �Fq��4�\�;H�亵ɼȻ6:�M.���{�q��x�(y�2��P[�éʰ>gU�7�w�ޮ��:r��fdK��6��p�$0�}��p���M�h���C���.3f��k�7ݴ�ŵ��C��2;ֺ��2�;Yϻ�����r�8>�85`��r^,��xrva����7���}u���g��3v0�ǲ�vP�i��F�l��l�v�Z
����墐��(�̱����WpᏫ8��4������m�-��tK:�c=	���;ʟ�]��6���3��U�H����O�td�\U/�x�Ƚ�_��o&}����OįM(�zsޗ����O�۫W��l��3B���(7S���y�[����T����98Pl���H��^�1EO���
V��謹�p 9��yF���rS��GUi�p�}Di��W��ĶQ7�x���B�~�-{����@�U2'�C�NENw��mOG�������#�+��8�BS=&�Xp���\�=�~��Mۇ�A�'ՆG�Rv��N��ޠ����e��Q�y˹�5���O��o�x��zm�S��xc�͗��X�n=��&����G�x�X ^���n�ʒKOD�c�X��ϯ�jhy�N��X�8}�r�Z��]Y|4�8к��+C��ސY]ܫX;U֣Q�.m�6A���uے��B
G�ֲb���L
I����o^��	:ˊW��u�IC�^κp�itv��;n�GfG:�U;^�J���}ژ����<��п��T��t��lq/'�P��U�Ө�O�Y@;�L�N|Oc�4�8՗�e����[��f���u�o��i�Q����F^��Lf�^�����t�S������נ]\o:��|I�ד�V��-50��a}���k��:���<̓��y�wJ���0�j���)���.]x�}Z��bV����;P���a�f׸�zxܦ �M
��:'�Y�9���{�)O���ꥩ9����T$g�z+E���ˉ���N�<7�{�<~Ou����t&����T����_��Ͼ�l_{V��;�̣�PY��g\��oEh��Iӷ2�x�Ӳ�K�r'֬T=�=_��10Y�ގޗG�|�m���ޯ�8��Gq��x�*��g���#t���	p������|{�c�2kK��gT��:�''�43����>���v�5�w�u���u�<k/N.C��}p��f���{ōͪ/ӛR���v�x����^g����rZ}q�!��P�ӗݜ��{(�*����f�(�I�*o�G����=���s^Gý�=�ŋ�׌O�鹟��E߂��y����+���Ojd[4��y���Hj�����
�G�,�Y&��m���ɶ�b׼h:U�u\ͬQV���.�Խ*)��y��F.g�d�K�b������鎉�\�;�2�`5���#�����F�ɛ7x�`��w����� ��)��;>rM|O޹�b��N���N��x�9�H��~�yuۃ���;�dJG��X+����V*�˰CsPN��ό��������fg���NGz��l�o�����q7/֑Ͻ��9�����EǽU�/ �R��W��
ky�P+٪f=#��T*
�g0�2!u?��������x�zF���#�F�he�E硥��g3��jN�F3���~��dO��tdA��;�����Dz�_�0�izgކ�>����\���Vz@~��d�t�D��Z;q7P����11MV��}�z�5�WGGg� �U:]@T��϶x�f{���q�u�x�=� ��?
`�ϑ�S�+t¼�t��/O�:�y��d���Fj�^��Bǡ�b���7�<�!�]�/E^bJ9q2�m���o7j�&�iN�wnu䍯կ��g�M\mCf�o2�3������Gq~���>���J7�,-9�J���*�1N��#����2v�o�-��v���<�:�����}�q7�̆;8?v~�|��׈�\C���ޕ�]'`^f�Dї����F�}j﹵�ё�J�4���00��8�+���O�M�ڐ![��x� lVf:LO�]n
�Wkkka��� {�������ڍ���碞�w �s�.Rv-�-��Z��UАv��:�u{��D�ڇ;M5��Sٸ���}=>vX����댖+Mƹ��`o|����@������>�:�)yᕹ���/۵�b�	�7^,�c0Ζ7�ɝ�t��k�c��{Č�/"aV���׏*�#���s�}�Z��Q������,��~5�����}��p����6_�!Ԃ{I��IY㎰��!t�|w����l\�z���C��
�D��Ia�3��\4���`=�^�5Y�aZ�y���D����;��;�\��_�uj�ȅ9E�� J��<zz�[���2w귍�w���/���T.�x�^��~Wϗ��p��<Z;S�7/��jr�*���c�G����=���f/-������H�>����c���!(�����l��B�g>��}~�A�r�o?7�a���z��u�����������ز��K�����gQ���
Q���b��?7xaS�ߝ�#M�h�r�B���_�.�14��� ���ǥ����&S��� ���Fǣ�U��d�R~��g� ��^6�șh�����~
��c!��䵯#yڷlL	�7������9�[�9D�܀���$�B]��o�IwycG$�<��Ӣî�QWNt�q�@��j����'_V�u�:���m�^��SyБ���[xP��J������Up�B2�tOZ�{f���a�?x�S^7|�{!�`\{�,����D��>l͆;�΋�S�TA�޵2g��/ߗl��sF�)���c^����t��yw�(�Q�>%�-73g�پ�W\U]\�l_��My8�u��4��/Ǔܸ�}^wr�3�N���w9]���P�===ΒQ��g���ӑ'�����g0��	µ��gr��{#��q�-��ػ+P�*5�y�Y�gt#�2}�̫~�����Hh�ɇ}�W��y�Zo\����G�vO���;l�]��=+���IO�"r"��g���P�
�B�;��g˾�������g����>��=��j��}�,�����~�[&���v�����-墐���(��2�����TO��9K����hgkS=�}e#s���Ϻ��nB~�q��O�Wo���/^<��8�-�%;�S0��	񙣕y��Hy]C��Up~�^L�>�_��S���ޯiq��_YzyU��ݭ�-_���+��4�7<|h� }�+���LT�����6��G��Hz8�㧴�-L���Y/�[���1�{HLwe���8�\nW��+�l{joI�ƌ�=�!���[WA��W����r��]72��+*�{�W$	bm/IJ�.2�["�9��4�^���o%9G{b.�<��#{���XÒpǹ�����sO����%���3�;��#H��^�_A-�M��yξ��}�B�tj��GL�F�O��^�5����#��wސ3ޯ\xi�sq��Cn�Q�+԰���	W^"��S�[r�vO�z����g<�|�#�d�+��#E_�܁p��p��G������4Y���R;��=>���}e3ݢc�/�TOD'k=g��/ z� �<���T��D���TO�lv�̬:+��ށ9�G�YrG��Ӱ9����p��G\{���>>�g�K�{�D�^�5Aٸ�WRi�����'O��3��߳�G�.V��|{#T��Y��s��~�*D��{j�b�MP�$7m��sd�d�7���50��n�y>&�\�3K��Zud�^:R����e»�l�����{�P������"�;�%a�/���B����a�m{�x�2�<=���e�G_�e��� {罯�~�>rs�B��n`���pڙl���<7���#�$�S��ש��R����}��Om D-�~'��G#�����Z�����u��'�x_⪩�ok8�{����z�}�S��ȡ�JC����?dw�}#FѺ��62��+˻h�0�}�w`NX���l�{)���U�ٲr����:gRy�G"��^\�ގ����v�'�&�R�-ɲ�3W�^v�޳V�XKRM�շ��[�1���QsZ����	,&�,�@u.;�\��¢�"�*_�"g(���������L��q���;�θa�k�vNԓwTyY��$����!��ם L�w��erCoV��9nV'�/����K8������6(�J�D�	헷�v	��2�l�ι3o��po�(ʪL�y�1�y,wZ�3��5Iۭ���������p^����M��°�|r��{�Y�(�l1Z۵�]+lhU�UϢ�[��c���{��P��f^��Z]0VLX�Δ2u,��k����+�B�����4��	�t�A�w�g]����hh����P��n���fr�]ټ�h^_��S2_����� �x��"��s���ʼ�(T��E{�;�p�ͷ��>��F�%$�J��u!!6�|�])�d�n��#u2�ΫZ���*���՛���hN�R�*�E<�\����Пnƅ���[���M�AI��I���Ѷ�[g����$��+�+�HC��MYi�[P��0i_;�t�NY�;\6#�M_<TK�����H��Ԡ��p�Z�u����o�y��l�mAN��������0k�� �o���٪����B��渻��\%�-�ms��,���v-B�Yq�s����і ��׉�a������D3�^Z���QK��N!o8�Jk�ypﵰ�E��:!�!]_�z����쾾����Ϸ�9�vB�S���B*o]w*���Cӭ^����`]�Ǡ]�*�t.b�m���m-Ҿ:/8���1�(m�%p�b�㻋#�ٝ�6óv�-�^���#W�L4']V�3��*�m����C��ܧϘ��b]��HDbwډ�F�F4�{�\(�b�A�r.	�wTV�5��l�9&���ڸ�Ք��s�m����տ�EN_'z��aʵCc���l�XF�ԤU\#s/T�-,亰Vn�Q���Wh$CC��+n=f��)�������i^d�Ԥ׮�mҜ��)�=-ŗ{mT�V9s����m�b�|��\ଂ,j�ܺ����]�,;8���=�up�bg� H��tI�>��	�_GRFt�녤0�vڊ���XE��}׀�ų� '%ۙ��pѥ�@Z�7neV��I�=�c�@�G��V��[�)�݃�ٝ��^�@iȕp�s6-�Tq�h�:��ZE�w33!�VT���2Go�ɦ��N�AK�ؙ:�h�x��4[!پ�׼+L�*�1Q��R�Z�Wf+�s����{N������"�[TTXV�DUUDeB�lE��(�����R��*��Ke����[jX�(-����QQ�֥
�T*��AU����(ђ�P�X+���X��
��e�l"�2�QV3�"�LV(�*%�(V��U�,X�,F[ecl�X�őBصAjQ�(֠�E��[
�TUZ�E�Q(ĕ�(���b*,�V-�eq*�Ȣ�b
ť(���X9h�QQ"�ŀ�e��U�PQ�Z1r�Kk-�*ň��X�TEV
6�Qb�m�PFE �"�V0R**��eE���hX��R���(�-�Ub*�*",��b*��,X�J�-)e`TQ��b�++cX���Z���"�(,E�
"ZRVDJ�ʩ�
�b�+R����Ŋ�6�kj�b�h1-���Z#Z1TU�ĶU�F
�
��R�P*�F����G!��{��.��s+���D��2��4ͪ���$���c\�_�<�8%��"�]�c�[����w�鉙��hIRu0����=��wnv�@��j|9w����u��pѿ�U~�ơy��U1��<��6�NkIx�ϥ��U��&��ɝ��κ	�Oz�n|���߶��qד�ot�b
�tB�T�\�o��q�> /�?>dp( ;����+�Sn{Ō'_�R�#�Pwg��-�̍��\]߬-����/m��;n��;>��G^������U �c
e�=���Y�!{���ع�/%���CǼ�FF�%#��{���A��S��v9���D�11M�&m�^��f�wpUyW����_��D�Ke�X]��E{���ϔ�^�����9�&����%.��|��w�=qV�q��^�C낍[J�o�~��{��s�'E_�܋���%��E��س�{tyπ9�`!���T-�XZqt��n�o�RX�w�'x�n=���|k��0xs<�����=j��MĔ��LL/U�&i�x���Zw )co��lvG���c�7�=$ru�9D�����a_f��"\�
���6�Ģz$�v�n��O������q���_p�[�O�o�S_�̘T?�%�;�dCUj�a�d�;pw�ޱjx�zJ4���F#�?���sDȊJ�Ɲ��4�7�T�V�P�V6q\<�{r��'��h�(6�LF�ѥ�i�Wڵ�5淝�x��sy��B�]\2�^_ j̘#n���Յ�U�Af��E�U��G̓�Ä������ӕ�v�J3��H�c�g9��ϝ�9ߤ��VA��H��;q7Q�{�K?>F�x�b/r�z�&�{uZ��Q��с:ǹ��y�Y���<�<mL��fl/޽�7מc"�����C͞ӣ����Ǽ[˯9�]%�T5�ۙѓ�{ģk]�A��;=�s]^(��w�b>�Kyա��;[7X�L��R�Tg/\{=8�&��N��g\L(Xw�������g��v:�h�%鿧҆��xfһ'´���o���5k�����X���5v�_�f��xW�h�K�s��:jWXY�|����o��Zx|'�Z[�N�^C^��3��Ѫ=ӛ>;[�QKP�x���SG��B���<��1y�R7^�0�w��L�>��ܟ���@m��W�o�O��nD{��9�W��exuë�6��Q�%Ir���`��j<�����*=��H���ϥ��=�I�~ӱޒ��}���J�.!NQe�%-�a���{���S}�7�F�V���˸{V%O��������9���Y�����N�>���MJ�Q��*w��|�dx���xd�&.V�.��I�*�'KtI��!y��ݞ��z��u,��i�c��7V��LN�N�v����J�`�${}R
�8�*�1�'H�X��A���v��ϓeW�yG�r�-�6񺃅ܩZ��d�ݥ3;�_�9��7��:�ޏ�b�����<Φ���3�����6}|����a�O���>�����8�O���l��ba���F�%x�!��k������'�j�� ��>}yḟh��C��>��$k��ِE}n��P;�LL/\�c"�W��Ĵw{ݗ����y���i��ﳗ�����:�7�(a���˂�?�n&[;q2�__��j�{��Vy�X�X{����>GQ�ϙ����gGD{ʯ�>>t�3`�G��ȧ��D�L�-��/~[�XMO�ǤS���~�:��l���=�R��7f�oZ�N�{��m�G��*I����^Y����Z/s�y��>F�nPW�Z=d��F�fjKN����U.b���x�ROM;�ѕ��P����+����_��8o����9'�����g0�d�7u��ge��BW�Ckft��ͣ���M��f��U:|��bo�GTw���Kgn'j_�^����5�Y=W���[�^���r�� �@�:Ƥ���h��~YhP}�p+0����f���z*��ץOuT�lc��F`�����'Z���jX�E�ۛ{�yx���_�����ZҘ��ԴA�C-u�R��9�sa�m�1YM�jeg6s5��s���|���`�"{A�od���`��ĩ��7[��^�n���]At�d�ں2��'M���=���xc���ײs���Z
���8o�ݤ2�C7�0��{�3�8�Qҫ�t��r@P�c���u�D䰙Ϻ��j~�i���k�����w�#�h���}�]�^�m̹�IS_����7޸w�)φ>�~9�V=�7�o����_�d��L���LJ�C���rL����XE_� J'H����5<�&�%��۩^�!��������f���r�K��g��Ҵ�#՞��%���ĺ#����k�[(�¼^��!:�n�s�����>�����H��+c9�)���t��� ��P�!�����ʓz��ӑ����!�����ꍿuG:���d\K�$r>���/=�F��[��^����$ͫO��v؄�U�T�V<��[�	���B5�~n�}=O�mp+"�� ��ا2�����l����$����}c��郃���"iOi��;�9U>8׍G_���˜�����x4F�{;׆�v�{�H��s�x��c����y�!���"�\�g���
��N�70'��T
��w�QYet��q����n-�ێ]�9e���[}��l=	�R�n�S�����6p�`��t�`>�WY���jA�r�{�v��gel���Gp�h7����x{*5A�qvt��˲ �4hi ��M8n	��˔�du����s� �����֨.�����Y�*&ޡR3'7,�Go�.T����D����+N}'����5��_}���u�v[���6�y�)D���Į�����x{ޠ�.<�k�����"��V�G�v��'��H�����v|&������Ǵ{A�>�]�?c�󪖤�yQ^�]�z+E�ޓ�.e���Gx�U}1 �q�����w���D.��z{Ǧ���`
�]�<Nק_I�z�鯷��Z���k$������Ҝ����uy��D���r����sz|�m���]��7��$����ԃ����֌��fE)?yG����\�=uHz�&��ɝ���W;�;�Co�O��o��[�H�'�]P��R���zOvn�p���}�{��%��%#s��z��`M�x�y3�ӑ[t���wa�t_m]�TK�)m��j���Z����^�p������m�[��|���T�>'e����=��B�]��v�^��)~�	���z3�R;��1�}v�ѵN����N�޹�a��ܭ��ˡ�t����z2=�y�^�}�#�Ͻ�~�(��M���WѾ�4T{����9E����1pN*��&���J.*4M�Q�x��Jx@�r�t��N�64����sj�)�9�@��ɭ.2.չ[7��6�I�u��݆����1ʄ���)W{�VwZej;8sN�XB���{dՕ�Z΀�]K��B|D�J��FW46��=���ϡwue�l����+�ՓB��0o'��r!��F�U�-{;�G���^�{({k|rm�Ҏtn�>r{���I���T*�#��,-8�_��7q>���?��89h���o��I~Ag�y4L��Y����ȫu^���-���^��D�9�}+N�b�~�����������/<ُ>���=S�;��3N�Or[;su���SU�n#\�wc�$�ԐNL�n8�9�^w��?p���8�	����r ���u8���"��������}y[�����{E�=��<��OD��}�}�����C	𯗪�7�������m�p�J9s,v�r�k�e�?�o +�q��Y��j:�i�/��ʇ��{��uR�9W���G�ڜ/�(��m���5��^3�f�2��t��h��N�Ά=�6���=��eqRY�B��ڋ��}j+Gb�v�'=慄�F՟�����Y�q�g��n5��M��,\���Q���
���0׵ѥ������ܸ֟FDy	�7%��Ȫc+&����}:�q�s�uu�����3�LY��gSk.X��K	�ٹ�W�vF
x�N;�V8;���"�˻����$I��co��f���wV3���������}�J�ͥ�=���yA�v9��ƙW�G�RD�a��v:<ݏ`���/��w�R��[<��F�5�d��>�=�9�������(�)��UƢ1]1>�Sc��:Kͬv�|��ӧvf�tӳ����9��y�߽���j�����AdlL�_Ia)�T���tՅ�y���h���nx�>���_�G�ý^ӛ�L������ڦ/�=E�O�'�~l�#�&�or����Z���b����Je�7ׂ��~W��H�#�t��}�L�ږo��wG)6��d�p�|��`��h���t+��n2X�;���V�p�O�ُm׊ o��������g��o�i������^����މ���.��W��^6��x>��*S��T�5�f�f �s؝�h�G��������Nў�������w�A	��p�����y��=Oz�n��s��2��>4k8N�nR<��>>�@����q�܂-ύ I|uL���'^G��.��osܺU�q�ޭ�q���Ȅj�צ�/��_�z}@OZ� O�(��y�N�Փ���;�g2}�~����A�6�h�Qn�N�i���񿛳Q�z����q����s�K��d�� 3�=�ڗ[�t\ahT�����3v{�ˣqP���]���x��t��h�j�gpͅ-=C6R������qih3jg�3y�}�d��7�_E�&1 0`)V>L��uԕǯ:]���Y|��k��NƘ���|}���tW�i���:U���V��N�_���է��	�d{ws��Gep�zax�R���8���e�UEz<���|��G�Ν�ד�}q���޹��n[��}��VӪU�r�y㐗H��p��֬@��tx���q�m�1}�=����wѕ�,^l֟b����3$��a�w�'�m��ul��k����ɿ���,Uv���Z-`��Ix|�*��f����:}�z˺\�z;�UD�x���vC�_������/R
��<�8dyh�/2J:�oM�]�t/�i>a��y5>�����Q�'�ӓ��Ȟwq��W�������c5	�^xz-c�Q~��Զ�n��p^� K�,0z��O�޸w�L�>�>�~8��c���SӞ��Ţc:��W
���,^
�ڿp�U��j����yl�(�OH����1<�&�i�}�8=/z��e���dK�z��:^Zp{��;�z}����X�>#�<�g�WKo�,�M��x�������z{U˕
Z�#=�Бq�y��+N�d�{��Q�^5������&7�\)s�3�F�EW��Mf2�yՑ\GSy�.5���+nm��VW'���:�1Ӷgs5�(ŉ-һ��rs䮇(_	��p�E��L��{���V�'nѥ:(�}vd�yv�ݖ�H%�Rͥ�x9!�������r�ll����n�ݼ8P��wԬ�żw_E��*om�ŏ���5�.�<."_�#����+#E��Z=��ơ�<廯xݵ����{�����qПh�#rhQ}OA>�ơ��&�q>��⏶��X k����vwi���M��b��NI'�08?Z�&)�i܀_���S/M����,���l�L������F�aJ}ͺ����d��r�F��GMK��!��+L��;�،��Ш�w��1��L��Di�����f=����M�t�I�9�+IGz>��j�2�K����5���f��9�I���Dǀ�c��=�%����3�A٥�V=$�7�V��^��0��������!���x��%��3ΪZ��TGT{�v(\y��<p��Z�Uԥ�A��N�9��/њ}��G�3j��i��M�� R�w�_���G��N��_T��Э�`m�Ӊ�������}�U4�i
�ʇeuMf��f�J�l���Gq���p��k���m(�v��q$��s��z�Td֗��:']����t'��<�2A�~:h (�M:��:Z.�~z����B��f����m�d�Vs��X]a�s{:F{a�m؁���{}|��W���Xɺp[��$	�:�ww�0Ws�齇�n)��c�PV���ck�%�ٺJ��nrbno,��]���5���2al���������{��׏#����8JD�`���{ŋ����ȭ�A�UĂ\��"��	9�Ҥvsi�}�3�=��;뗧�U���~�>0�퉔H�*v*��O#�\eFn�1r`���yq�<�^�6���ޚ�>{޽��H�G�^q��a�{�������b�>6�3�����q��FgV�q�x�����Y������c�}@`~�W���}�&�ʮ�K��jf�M�vbk|%O�� �7]4(��G؟\j-�q7/֑�zB<ϸ.41�h{bUԜ�n;w��� {��R%� y����jdas�s#L������UН���؜s�Q�5�3߮���{��,�2��+�	�o�QH��e*UߝGĶ{����;�,mU0���W����s�T����S��m/L����
��5�ĢnKGn&�_�^&)��'���Íi�T�Vw�7���^�C���������OJ��<���o�X53�Q���ٵ�M(�����y��:�q��T�iz]\CW��ӱ^�%����r�xd���1%ߢ="���P!M]��Z�ۥ�=㕜��n����Dw^�U2��,��S\y<)����.�J�5�ve%�m��Nb��!Y�X��5,���Ґ��w�y�z!�%�U�L.�	̣F��;$�@9]z��7�ܜ�t�?Yl�=\X:o)�f��pS�])c�G�B�Ep�u���^̽��^*I(n-�{\/kH�hؖU�v��������ԫ~H��+��*�Dd��;3hޅ a^)`\ *�0v�����.�D]M�f��&��n��Ʈ�:��F���ܮ�7�<�*je���G1��@P���1<�9�Z�f�͏;NRʢ��n��n���DE�������s".�	��in���_	g!�ٝ� ��qi%�ċ�cF^��&"��z�Ȋ&.oe�u�MΣ�+>l�Ȏ�M5���Ρ;�l�������=�����l����Eٱn&E��ֱ�6Ю���>�YUb��Y�Y��t�DՉL�2 @���Ho{���p�<�&<�? ����G:N��y�w:�m���#!� �z�N�X�.�7ct��W{B^
�t��A������2_N1�*c:7���S�Lں-Ի�d���KFpɿ*ˡ6��;~@�V�f�U�e+�ust=e���8wjVic҅b��wq`z��UW��5��B!H=b��$)��w���v�R���o���.
	B<�ë�72������Glq��I��{�⩀�V�����Gi��hɧW<7t�*�6]0+_������e���Wc6��pN-�=1ݨ�u�X�Zf�T��!�E�3k�jj6Yp�R�ߢ�*��X�]��,]e�8���MQ%!E�86�j�+�BOF����������&� і��U�n�#�[g�i�[:3�,��c6,K�D���L�U�gk{^7BQ[cD{vp|tl8/��M�
�Waz�䫘�r��Ƀ)X����j&39@Нk7�y�iNn �l��m��&�i]R�Vq��,wH�v\л����"ؾ�3�v��;�kM�ߕ���uk�Z��{�P�jGk\��E�)�z�ms��[׋M�VÆ��;9|����1t3o[�5VFP��=<��v؛GX�U�CwdGIDv�5�[��Y��IYJ�����p��F�\n�Seԅ��X�4k�B�$h���_�^o=�ĩuݹip��$ƕYV�2	fM襠"�Y����'O�ث;��f�noG�����f:�h>���R�;�{��U��+�u���e �.�������f�����Z��Zl���O|�޳K7G]g����Si�&�+[SK�G!���6b�@�-�twY�f��� ���*ګH����أ�'�Mo-�Z�������\�Ŗ�Zl��^{ܘU�as���SΊ�>�xD�q��fgv0��];q�wQ�!�5���+�ClNU�8�+Y�\lN_R��(yh�"�**Q�
,PPj�2)P���"��E��eEDZ�dYkDE*Z�Yb"�Ҩ���J�`Ĭ*(T*#(����QDTX��V[ET�"؋BVIEeem

�+�R��VT��,b*�"�VVV�E���0X�
U��Tid�mQE��E"%�* �EFЭj�V�R�aU��TAFҊ�ڢ*,b�V��B��*TP�J��*���F��aU��m��H�A-+Q��ŊԨ��
�"��bȢ"�
�"�%�DA(�kTb�щX��TY[m��*-J�lX�Kj1EX�QQ��`�l���ڌTF$��������%#Y+F,V�1���V�"mF������֊&�0��Fu�a�.vud�:'B_c�,����u�`.q[R���ͻ���`#|��g��ίO���c�T���m���|�[��ͥ���&w*�{�~	̖Q�uF�P��2/sr'&�٦k6�ʱ{�nuX��d���ς�D챞6���Ǻf�X�=����x�����m�u��m#j4b��'�3n&��l�|zt3e���!��O�o��=w3,9�����j��������(~���%Qϲ�VaQ%��Ȫc+&�����w���w <�e���X��W�H�����y��ޏ{-�-��^`����~7��l3S�[�0]z�{�=�)gԻ2%��N�m�������p��#����BP�1R�׆��n�eW�Y���$\��G���MBb��=q��]������=��^ӟo�2��/Å�:�lO��j�^Ω��t7Ѳ�A���Q`LSw�n2S.��X�o䟞Eb�6n7�\}Bu<D���n�x3��ޛ�б�r�}�e2� ���+����N��w>}D+j�O@��}�ۃ���}u����c1�^�\���=������Q`@l�LL7r���V.W�{�;�v�ڧ��ǽ;�/�e��UǼ�Ώ�1��i���>�C5JZ)J��S��ƚ�ޥO	�Y� �v� h���]>�q��_7����}�6a��3��R�aj���V��ˍ��в�e!cQ�d#�T�Ҧ��YF�s#vG+
�S��;-4,�WR�9u����Ñ��w�7�V�cb=ҋ��l���{2lL.�Z:`���"`�+
��y�=�������y܆k�������m V?^�����V���92��y2�
�hU��$}�bb��������5M��\/�yU��ϝ�� G�Ő}���]��Ϯ�X��JyΓ����A�߳h�U��5����7f���=�<�r<�Ѹ~
j�졾�6��N�/�Q&���/pς�Dܰ�3kC͟	�4��j�=i�dz<�vb�S�M�nN�W���^��[3�Ͻّ�Öw���Ӓ|�5�_񥍏�;��X�s,�
��*}�W��ޠc�a�T���5�ʱ/�Ѕ9��0j�{�?V=�"���FѡX���w�Fe�o}l�l����B���#!���r>�q��BE����X't���E��M��s�+�5���r��ή�q:�y_��d>�_������N<��1�Z)
Mk�K�OT�M�H,�L��������w	�ONO�d�����{���߽�ŝ���TiG��H��J&��KA�����ҏ{{�n?��K���N�e˨KM-���Ĥ��wn���ʁ"X��N�Q&b�ۘ����G��rk�}f�P�������ҭ�}�o~q�:���a�����^ژp@�X��h�,L뭙.w_;Mշ����8��хJ�@���mV�
�>���z��ٵIφ�T��Mr<��w:�]D�+���w�y��㦬�<��q)Te��,��Q��z@�]SjyzM�d��{S#������S��J��\���O�џo�R��}�C��ǲ�,�d8�F�H��t(��%yw@�Ώ�]3��F�~�6��<#��w�3�tƟD����k�~��ȃ��z���v;�lZUWnyz�t�lǠ�V��.�>�*��FE��$r=���Y*�n�\{��p�s����:�κi�.��5}4*�xp���#P�_��\S��+��X~� ;�Y���x�f��z=����zp�tvD�c�j��{No��Ӑ�^��f7��W~3^|&˜�S3Ll��EעF<x}:vO���\{�d�g�I�a��t�\Fz�u+L��{^��4V��]��O�Wy66Ǣ���d�G����=��䛈gļ7'ȫ�n���������kǦv��sr�YP= Ͼ]z��>t]Ǽ�N��M{���"��%a������//z����ӃL��,�z����ZLt�V��o+���d
�y�J���>B��Ve�yRpW��b�2v�������=FZ�v��$��|hN�Uot�ٛ%cP�3��uURS_,Lf���Wa�������u���8(�jK��).i�8��W�I���d���� L%~�j�|�盹
߲�H���ޓ�7ب�'��MT_��n�����zg����;�g��Rmx����=�L5Q� �[��K��x��:w��"�U��Y��q@���'��o�Ԗ��Z�5�<2��_�>W7���m�����>�l��X��U�z�K����FѵW��mo�d�:.}8_�H{�{3����A9Ȟ�X��^��Yʭ��
a؊�b��%M���7{��;#�l�a�R2����x�-�|%�����[�P��e��r����^�����������^�sJ�+~��x��%�>�e���r��u^��~�s��>�l�Dqh���p��漏��z�/�}��z�:���b���S]��gK��%�k�*kՎ���7�5+T�v#
e�>�(տuǳ��M��~��kc�*=���5��@Bz<��5E��F�Ǝ��G)�x���@7(�v�>펨�m�Q=/֑���#̶�I���}���=x}�WX�Z���U�/���,;S 3�m�ә��~7�n�dc�.�a��9��pL\�,���:U�>�f�ZC���tQޠz%��W1�Q7ip�7��ǈ�������ԁ�.��:�`����ӫׅU�Gщԓ�����M4$ڛ��׷�#�Ι�2`�1k�M��]c�[u0,�D�����z�ܣ�6��v��]���}ӼJ8��>ͺ�V꜔NIh����&b������Zu�o��m�^s��^��m��^�Dk����L\A�W�3�O� W�fA���x�MĖ���C댯��
�S~Yz2�g�v����G�e�c[���[�_����pX�YW�� o�#���͜1z�v6Et%	�{;�6��Di��U���p���?L�r�nr�x�H�����ux/���{���Dσ��͎�ݨ��m{����F���or�<�e�+����x�&}*�sfî��q~gjp�?IG	aa؝�2�Ӂ��W��Ǻf�e�Q�����zÿn9;�s�Qw��}˻܍��8}��m�7���s�Cnv�ˌ�ү�
Ӭ���c}(�
}�;+,�p\����Ƕ�=��7X�)�Q��N鿤�>YLf�Ĝͽ1���r���WW{��Ժ��l't6�י"�5�"�΍^�ZϹQF*�JF�K�{�+�J/�;��$}��F+��;�9[u	�M;1�������W����^:�CF}�h��(������-�w�A�KQԥ~Yg	�\�hb�е����"�tڍ3yj:�WMꭢ
&����|�u�<�ޙ����{rӸ����o����}$��SѴBɭaǇ4�<��|V�lf��IoEr<�7/m��WsXCK���e��{!��E�'�Ic�L�"���S.�]���t��''�~ӟx�_g�����9Q-��4��*ػ�TL��p�H��;�!�-ׁ��)�Cڱ(��Q�z�.*�^��;$�}�;Yj�}s�ƴ�t�7���d)�,��@l����z�T-d��wQQ�t�ا׷�i�.tj����n�y��o��caN+�w�a�z�q�.O����f7����YsF��x#v\խ���˚/�R��;bo�Us(d{�H��t����fA嚅�������~8�c)vv��ߴ��wmv�ٟ{�� ?JG�G�U��u�\zl�<���׍�+�c|]z6U�g�{�s/{�%{�3M�1�R��7��x�!0��~5��S^*��k &�Q���������H��E�R����A���!T_�d֗��o媚.A��k�6M+S�����D��O���g�K{�����>.r���H�ܰ�6�<;�=���:�;�u�55;/����v������=��Qq�S��~۸��p��xT�3�;^�z����%ޯퟢ-�SY�g,�� %C�p���0�/p�Z�i�t� ؼ�]��<�w��KC�=h}~Z;`�Z�V�P�B74�<k�1Wd'jm^�Or>kipy����TI�w������_���p����oI�k����.��[q�Uh��C񱟪�(�Ǒ�:��TY�\М�{l��	�7Z;q;P�ne%s�$zs0{�C�s�j:<�kN����������#!����l�j~G�,�;�f�^6I��5��<�Yu���U�����u��w��j�f;z�M��w�]���v�	;w�0+���^d�Qz�!��d�v�&X��tP�b��f�N��'��n}���9�⻽x��>b����Q��FQ�}Zd�=���&|=2���\;ɔ��"]?�^�AF\켬��M	���Y��}�l�w�g�q�j�o�j�+#d	D���T����w%�W���B��f���%:���|������.o��SA��� rت�>�Q�[n������x�D�8�}��!T[��/y��ǲ7�����#�>+=7>�Cs�0��F9�n�/ؠun�>�]ꬣz�<��|�શ�Cz�9r�w�4U�W"k�'r<�\:���gcw9ʔ} c��L���4�������#P�m�����u�>��U�o��0�Ow����K�'#*�^�0�&�̫�Վ�=)R��=]vY�#
[ke���Bc���^���TXN�!�;��2�fₗ=����kh.D��Q�;;դR	��puv�*��3|�F�7x�s�\�Z�+����]8�W`t�|���˖;lv�� �e舷U�Rre����TD�S�ӹ �ӅK�i�M��鼯2���BB��{*�������w�I��{�d��s�Y9�t�\g��_\�2*5���w�r�sJ>1>���r�yY��~�znb���)rl{��$ל���$�����+t��#U3�ӻK�Nįu�'��R�����>	�>��9ҡ�j�[TAށ+	�*�=�<&��9�~�5Ҋ��ot��}�O�3��]0�����3/��*#��{.����Z<i�v�o_�:Z���~�g�A�Y��a�B/M�ٳ8p?��V��߉�e���D�cf���϶dQ:ϥ�����v�[�:v��c<n'e����W��f��7�5�����3��\�h�O�
S�*������R��.5�����=��1T��Η�d��b�']�N��n)��z�o*��g�N�9����q�8����y|��5x���.p����\��F!�7V��H��g<�O+����W]x{:��yg�����^g�#�^��F{�G�; ���f������Y��?
�M/�.�.{A�{o:~�k�~
v���/��/���[a����V��CO+aq+�7];MT�3O��C�(j��f���*��c<�_K]m�d�;{�\��s���o��V��ٸ���b'�wy�(h�:X�	HVA;��fk
�.��;��G��.}�I�͟{ӑ�0�nk�|2?^�^�h��W�\�A��N_�y)'6v�[��P��3���x����	��5)�Q;�x��}pQ�����Ϸ�,.����u|k)cQ��49½b�ꇋ�y��77^��@�FKGۍ��f��J��_�#����>�w佉ы��xY�}��\.3���zg�\ s�0Xuj�Qs�s>��2S�grwfaC�_���!V�f-
��O�:���N�(���.��dW�꜔NDIh��L/TZ�&����w��=�r�����*_R�wg#O|ݱޙU鋃�K�9>�_�����I�(��}^񚛤=�tBkߦy_�����z�៭�����W�:S�� ��e�Ey�R��=C*]glP~��������6V�+���i��U�~/��W���]�|��^��T��S^*R�,c�N�秜3�4����	C�~3a��n�;����/��ܸ~7�{���3,񨢢�R(_��݇<7�d�e�{�&l�'�����vX��Ӂ��WM�i~=&�X����n��n/��Vr�E�XL��?�#@��?:��w���{�l8��>�

��b�\��!�J��6�r ��t�X�d�#�VOh��s��z�-�� �җ�gz�UE��3{�,�G����Wkے��[Ԓ�HC��6ݨ1����wv��G�s���O.1gT��}�:n#�����|Oi��JvX����'´�^xS-��/5h{��:�����׊�>��o��{��n<�\U��<aX;��gܪ�ļ�� t�1�Vm9���y_�S-��w�����;W�H�k�q�y\:���C��Z�^`��\s�u:��U�&֬��>��z<�������ׅ��:ϧj�==N�k�~�q����}s�
��к�3a4=����NkS�{��.j$�����޸w�������������W��o���B�Ϋ���JW�=缅DmZ�<nK;�9U|g��M�`Su�l�[{V%�[���a2<�<�L�e�ܞ��*�3;�<V�4��c�(�� 6x��}R-�%�3��e�n.��ҏO�e)���}�Л����c>�B�g7�4���ì���%���10�EҢ&������m�O��:w����z���t�:�+Bn;^,l?m3�pb��5�f��X��G����+��Ĳ��k��c��H���0�po�!�=�B�(�s���@���~��ﾈ����$�	'�@���HIK!$I?�	 BI��$�	'��IO�BH��!$��	 BI��@���HINHIK!$I<$$�	'���$�Ą�!$��$  �  BO�!$I?�	 BI�$$�	&�$�	'�����)��r�� HU��),����������0N�y�$�I��( %%ow*�I
� ���F�Q@lH�""QR�*�)IQ"/0�`=�.� (2�l�3j����p7	�Z���� tw`-�5CT�p9�R1j��U"4ГF)���8,��V���e�E�gn�:۸h���.��C ��4��n�E���7wAwq�vvܒ�IX���m�T�]gtR�U��ҙ�7[�m����JjM��j��pw4im[j�#[L�V��ʙ��P�αm��m	[UV5l��DT�P�\��Q�PV�KM��Q-hiw� P@ ���T���b4 h��ɡ��x�%*R� 	�0 LD�hИ��L&��@���Flj�jB)� �I(�`C �# �`20110�L�L���J�Q�P�=4ɤz� M ��^�Ӳ�ֶ��1AUW��0Ur?h�EUT�
 E>d
��Abt�ϧ����?K� �a� �5TV	��������@$#%����8s���Z�1��×^X*
�����d�ʟ���]c_��ed5*T ����g���~o�c���Bjˣ���vNHVA&M��udL���;�Qr�V�����	P���e�$��S�KlS�AFS#\U�蔣bH�fX��v�j��W+�(]��jʕJ�7B��c����(2��1ޣ-	4n�V�7�-�U�+%AC���֩��c�Hf&P.+��MQТ�Y��b�{&T���HO!�n�J���ѹepj��
m����#���Q�F
��lF0��$ɚ�`�V�(WL���5tj�!��@;����5��G vs�Ց���/m�[���R����G��]���R�w�2ÃK��X�C]$��ʀ�Ha_I�,,��^N�M��Ȱ�W4^d* ��ki1��:� ,-7x�QKSi�{u�\��W�xi��*\.��u��@�A�kT�E�-S�m�w!��Jـ=ܦU#�`X����h1��e**�1n�^w�#R*���Dmf(	
�K�C��Bnb5��Pe���*�7!��Cb���Q��Ǹl�0*��[��\��+wYU������ b�
�!�z�E4���z�S&޻)V�L��bSRm�Qˑ����2iq7DQ�`²ڬ�F�7E'Z���@�݂;jذ�De��%��W�����i�5ZT��ث���;2+ɭ�R���I�$̱�Z�zn���:�gb�	VV�G]�ڼd�o2����ڂ�#���i4�N�׈1s6�f[�q}x�N��4�0&�o"x�r��,$�^$�P�V�h9[����r��	�E�V����Htfd#��a����p�]�P���Ky�e0I�����rX��/ql�w�4��YIiF��.�R�h�e�����Y��`ύ^R��Yhݜ,-;��xh� ��&�W�6ʥO3A��>׆��p�Q+�: F<4����!Ô
����a����ѸTl�b��B��-�ӂ�p%f���.8�Z���#����ǳ�a]Ve��i�S�٩>WRh�ݬ�"5�
ϭkV�ح^��[��b�Fj��Ь��1�J�"�[u�fmj����M��TS��p�+K��rԳ�4�KDVi1���];�-H(�[F�	����װdX�ɒ�ɤ�a�*"�+D�w��Q�%<$@���ۄ��Cs^�ij�ܦ�n��"mY�]�,{�[V�B�Il��;ZU7y�֊��d�PEG~�ue(���x/�dn�:��0�!$Y����cj�P�%����h�5]<*
ӌ"/2"�E��ii5�e13(�&)H��%��h�k5b�y�TkA�l�.��Y�
�n�t�:�VC �
ҕ�n����È��$�wK[7#Dn�&,^��	v��6�fy�&`T�B�If�6�<:`�l9viN'���bG(�l����^KUd��ut�l9t�kU�Kj�Be6�r��Ip"�l���%
�B-M��r�4�o���ƚ��YYk�R���0�Utv��pU���c�U`=�F�b�����1�(�Y�X������d�C�l"KZ�]&��+Բn�H?-��8�7�m�W[���7&O��2���d���Z�pn i�ͥ��\�B��ݼ��ō�*C	��44Q{�Sɇ�z����[��e4eK�iv9lf�Õ+�hH���cB�r����jZ�����I����M����J��4��4�Tw5��Ƿ�R�����l^d�Z�EK�t��F�*fmy���|�xֲ'�J@}�h�k��[�� �2���N])qim����o0JD��V�V��/�������������BRC�ݪS���~���?d~����Ow��$���B�GopG�A�g^�zJ,��=�� �z;d}�Q�k-b9]�[KU{=��e�^;�za�}j>ƅ����ål��z% �����R���YDNV���B�ٚ/����]u��l�$��r�:2noƎѽGL_;0���s ыL�h��_q��.�4A��[`J�����j>�H�ۥ�jZ�%��z9Q�=�rs.�iR=*R��5o^�"�8}:��Ԁ�
�[�-���.�ܲw��0�#ɲ�FjӤ����u���J��5��臱3�w5c|��;�Ђ�1j��L{3/r��ZSB��ĘY�erܭE�\��-���M��.�̾Vbc^��'�U޽7zىk#쳈��9O0�\�٧OCm�ѕ}C%fT[��7��hgq�gt{,�KT�f�n\��9�����sDM���v5
sj�B�Oee3lbAb�c��	y�K�yn��L��!�{[do|�:��vN�3Un��m>��V� wd��܆i�o��Fu�#æ��6벴���4.�5�_wrԉ������gy��w(Z�3Y�.�w���v'�_]u#��[�'\�W�r��,��o��2�KuuE@D��Ե��
QwJ�2�U$��dr��}�Y�)�C6�v��d7Y��3]L|�eF�ҙZ��v�+�5K!m��U�����YQ����3x�a�Zm�Su`3���X�q�7B�P�9ǩ*��	��nKuϤ��Y§l��

V&)3��e�����ÇZ��F|�ӳtSW�����e��9gs"�b�K���ى-H5U�;�&kz㋎ޖ�gwr�k�󊉏p
u��W�E���M�W.��M�nʠ"o�q�adU�3K�����1�bZ/(*�!��l�S�A��:�1{�R<2����:�ͫ�Ŏǫ��0U��6�U���g�U��q=�+0NW�7o})J�YuȽ�4�?���3mT�,�d�����n�t�
<�϶fp�-W9P��������&�E�C�Y�|+��ܮwwV-jNϮ�f9S����޿�j3ilǴ&�­[��!�w*1q˓s���D�xe&j<�Ywg�U�ݼӮڔ�t`�p��w�v�=��U��_o){����4H+J�D|�T��v�`"Y5̻7���M����Ҥ(i���B�}*1�۪h�a�.���#�h�Liu#�q�0�#\�����m�\E�o�v�v����eSHW�&��� P�#s9vA������,���n
��i��n+�J�΃�nX�~V�S��e�:����a����_Y��}��}����ζI�&Շ[ �[���`���j��� �����M�r׍3on����+zi�6�Y6��\���j���(+e,�ܶ�̓���*QVU�ܩ9�P�w ��?c�,�mwP���|�fI�/�vmp���-��N�ޚ�K/X*��U��k�V�kjݔ壕�|TVtcM��\{�G�C�ht���V�E$E潑.F�&�'5�l�bN�tM�����H�t"} _]���#"�\	Wb��cFhj>o���U	qr����oS���G��)��!a�s��WF�t���k��2�h��w;n�qV�)���s����)I�@�}*Ꮺ���|�S'����4�]�~DV��A6v�Փ	k�͜��#�Hq��p}a�R�h[rC+4�Tn$��`uIMqȞ�v����fg���ښe��y��s�*�X�}m�m�C_!C���L]�'%B�����SS�E�4�a�j�֒��s�̡�	�d�E>&s����x2������3~g�ӏ$��c��1���e��ze׬灛<�1��� ���	�SUU 4[
"���aAUw���ݑ3�~��<YA�]����Z�[�ٝ�zY��ΡU/n��Ǒ�n�Mc���1�)Zػ9<}Y]�/:ݷ/ۘ�
�K-RU��P]��P�����m:�+���˵�\`;vt��A�b��Hr֘@��W�m*��8Ц���
��g��VIC�w�ayg;q�XS���!��1���4�c�C� p̈襘���n�Z�����u8o1�L�}��Ĉ���"^���1u����e�eE�3
�[<�]*���T��KB��Zv��J�V����n��}/kH\�'�y�lR�/u�NЏ��ʻº��߭Z9c5�R̭�i��ҝ��kV{-�^lt��P��7�Fe>K��XKx�_9����M%C U���/��+b֯+(���yQ���95�s�Wq��%��f	B)��c��[�)nY�7��8e�U�Uej����������B�;��*T��b��bZZB�*�<5¯��30�
����zyΝd6]L���:��="��TP�A�uR�`v��t^��,��\�;c$aJ�A�����oi\�8X�^L��0����*���C��,wb�%(�*@ԙf�g)�[`.���4L�P�F��Ck��[�u)$�9�k��uB���\�xm]lzR�4��ƟXi7(�����S���/�n9��,�k��Z6�@�f�$d7v��g\�ݏ��\��%U3b���s.��y(�|���{������������7��w[Y[��F�K�ݵ˶�������xV7���X�'���Vʛ�f�,f���b�'$�	�CA�]�z�]e�-\ܠ��n�	kV;�*��x�)�,��'Cx�0+���X���-��y��r�6��P�8���Z���B_ob���0�,��Ż�+�9,���t���t���|�8����f֢�CĊ$9�vխ��)�^��M�X�E>�;�!|L�t��u
�QIt�c��;k��Ү��ЋL�l��T�ܻ&�p���AմVp�a��y���X^K{mރ)��t��i�*��޴zl�M�.=��5+�Y��f[�Wuq����{Z{вXp'O#�Ӯ��wYJ��V;i��^�2�v�����t���@�۔��Sz�d�ms6v�ox%�]!��f�,��`p����|��c��e�W��t�y��OWR
�\lgZ��
����������2���Z�ɗ���u�c�^�,I��Y��άk�)n��v
��_	��C�����Hq.��sg	�csg@��u�;�÷N	�r�Z2��r'��\�(��v�%�]�c;�Ø��1�6���
d���u���:�EZQ �{���̸�ä���t���Oym9B�Y�����S�Zdȝ�`$>�w�󖳸���|N�}�\	<F��l��v�ӵܻ��q�9&)Z�AnvE�0J�䘲c��>���;����<�cǤuK��4��<��
�yV��u��o���x��ǽ�`���kVt۽2���cW��-�v��a/9^�����S��ec8JK����o��G����Ta��J�j�l���S��)�8�Pw�l�)2�y)t����o���[:Y��:�;9��M�v����bl�j	��ٛ���o�mf'�W�a5"�r��ھ�Y�7o) ��l���i��Q,�v������9H������v屄Lok��afD^���Dc��;[%������'2>ٻ/it���;��K��u�!�=^�뾕
����U��t��;E�:}�۬5����Nb�)�s��PS������/��6�����Ƨ����*���"п��]P�Sx��zѠ���3o's��6��p6
#Sq�Jn��u��:��c�o�T���>ڹ��άۉW1qwd%��ue�rv�b�-Y�/��U7%��i��N��Պ����=��8�삗ץݭ����{�((�P���L4;y�(��]f(�Gh�;h�sNK@����JJ�K�Ѩ^0h9ٔp�Ո��Ї76���DN:{@%*PM�Sҳ����wv^L�۳����t��k�+rQ����#��a���.�6Tp��."fQZċ�0�VU�U�TZ0��5�ih2���j����cj�UQF�����F��#���B9��.���@��i�Z�EW�5���g����u�+[Ǧ�oa	\{}9��?�Z�S��8_ }߳����+I�ފ��m�j��Gh�Ec�2�n8���j�:5"%�V�����
4/��<w��}�O�q�G����K��U�����yzp<oM�:5��~�#�g�^���z������v82��7���se�o�ݩ�Ը�ص��WFDY��˕�x U︎8�Vm�T�.pn��.B��:LҴ���.��+����E��Q�qE�SP���*�1|WI[�~BZ±�QP%��s2�gH�պ�� ��e-���3���p��N����,c�K/z_"ɸ���]���f�JU��O{�c��=��^i�U��E<��q�B�o�����% .}7U��)ƽҝ��N^Z�`BԞ����om_\����<寫n�h���?1�Ɂw��+��+�ȰqC�N���;5�^:==�6\�,i�h2��Z�!y������������@{\���e�dA���ZW��|�0Q&��Uy ���/�̲� C�L:�w�SZn�IOgU�Q�V�X�����cܸ�;�JC2���0��z*wԱ0�$w���ݣp��f/=���4s/���ynD�E�h�f����ܪ�/�RoM�ې���ٜ��*xV��M�{�w��+E�³9���c��=��\�|�Y��KzE�{��1�c<d��sUm����?mJ�4-v�������DYE׹��׾��P5&��۫�A��Qt=���0R�I>�}�qC��������a�Wed��lMm���r3���ո�]4X�'�%�s:�)�++r�vqW)��k���ů:��.S��/1���AaSƜ�'�o�ʾ�[EU-������$)��e��;h��6��aޢZg�\m�'�^�Q�G����4�wZ�ٻ�Ȉ�'a��T��-�U}�¡�TJ�,?eW]%�G�����<�r��$�xʛ�Qs�.�j����~燐�.���NU9f�:���tǘ'���Ŕ�/bV}�:˟��<^�����"ɠq2s�����4�i� Za�{Pv�m�(��˻놂�<�Jć���Q�W�p:xs�6����oZ�JH�O[g������l����"�q�*Z���P�U����j�E��E^��'�Xp���1�����<���+w�}�s�~��9�k�3;7��0]��i����^G���f7�G:�:���wQÓ�I��算��a�M�׭QEg<�H;X�R��f��@t"zQ�.rVm[;�t��zg8mS<�w�(eEښJ�%��,C gKo+m{e����1^�*g�:m,�8�u+�^�N��9P<9����LlS�t��"����F�_%�>�6�XP�)N1q�_���ƱQ'=��|��g�[K;[W/FU{�[��U՛!����G����eo�f	�������õ�AZ��aU{�}����?���z��M-A��H8/�����i�SU����9Ƒj�ޱ0���t���>�����H�/�J�h����4>[�)��t4e�L���y�A��MX6�pȩ)�a������oL�r�o�k=����5i۱ԖV����I�4)gA�5D2�ق���w@�V��Om+zێ��|��vD㒹�Z�:z5X��V��U=����o���m�������>�xm!e�ͫ��0[�Zd�$�s��x�"�YHeG.VT�<�j���h�0�,+��#�� T�2⁐��m^E�tI6T�r�*4p�7b�y8ڊ��5!��eۂ���R�T�o�yNb,2}(G2,&�Z)���q�J�	r:�g&]�����8$���kN��DE���3p���E�E�*#H�-IQKB"�4� ���lE<�\IH���D���J�mDUd%�
�#$��Z��(�*�AB�m#$�hBI����8�W���6����<�æ2���d���B�n�U}i�F��~]��~Ȯ��ݙ�K��	v@�ɨ������������w]�΋������ʼ7�盏v3Y�
`��YQg��(��t��r��}#��rm��Y�4����[�@�k*���z�A�QWmV�
�"t_��]�T5a{I�Ys��n��k�3X��"�x����<��ȶ|�N�Y�{+�(���A�MdC����fݳ�
��bh��pP�0T�hi�EgYd�c���������_������j���M��9!���yu>��P�d�!��엻&a��t�٭�ȸ�u�H=s���8����f�5���ٌ�Os8^�P-Y���O͆��˹��O{(6�Z�j�w���[6 �jR���ٹ~�Yo;��b�kR{�f���<)�霷A
���6 f�]N�U��U�C�=ꜹH��3�8M}�+�v��b��ǼҢzk�oW�KH;�]0^�B�WW��ե"&P�/S9��T4���x�y[�n�@��>��=�R�?W�
4|�h�[h��V�0�T(e
.�������0�Q��mQ��@��GZ��WZ"UkHQ���w�Nws{*���0��+-����QƩC��8�e*����3UF��5EB�J��Ta+��UGZ6�-Q�ܪ>j��(6�zO�K����?QQx#g4��Ę���'s��Vܠ#R�H��ڷ������s�L{މ�(��R�r���Um4�[h�Pk:5��fs��G�Zh�W��@+��XB��h�5\k�����l�<Ѵ��[E%QƂ�ڣ᪣���L���h��T�9�4Q�UGkR���Q�(�P5TZW�{�:*��KUG�}�5���Z�6�*��U �@�S3��Ek��B���*�����Q��ꪴ�XԪ��Yh���w�{�UQ��E%Q��U!檍%�*�ä�:�GO�����
��젬�B�J��T�QƊ0�UJ0�X�9��Q�J�5UZj�r�:����j�� h��+HM�5��y*��U�5DB�vUj���3�m_%m���������1�1����-��:��'+�gs��A-@;y���7�뿊 �+�UU�Vڪ>Ԫ8�m��
�Q֫iUXh��9�wlު�TQmTj�!TM�<�e��T|�u(8�Z�Q5�o7��6u������TQi@y1�]D>B�![j�=�{<�\J�U���U�[ED
���=*���鳮��J �m����_�O 7��u��W)efQ4�I[����3��qݯ=^\��n�~Q\W��N�%�ܿ1Rc��������%�&����M��mn�|&�J�:1E����+i	�PB�{�ӄW�y�u��߈Z���[�변�"JA�,�����P;��w=k������`�YI�~u�s���y]�%+��zܯH�1sֺe;�T�ucm���ȏVx#�xp�^G���w�N�׉��,~�^�G�!��,	I�}N������Z���˨CF�Nc�����,Auyy��7�J���EgX�vm�
� ݬvR�J����٦t��=ѯ��G(�{B�,Nr+��0l�v�2+Q���s2�F$c��Ǟ���!3
=��ŕ⇳�Y��kM?��P��⻹��K(�<җ�gIM�;��nHb��8���3x�}yX��?d�{LK����gR�������>��A�t���Ys�1Z(�����CH��v�u\j��6Źb: ��Bt��/�]�P�z%u	�1Ϻso}X����O�F��h�]��d�?���yxj>Ϗ}��R��c^i8V^���|ד������k_��ϐ�7!�Gk��̝E�i.���Ռ���a�YF��εg�}��:���W�0���.s �<��$6F�,��-�_�IA�j� �KFS�ߑ��+u�PH7!<��l<ܫ[��.�\:�v��6���*��7��
�+��S�ͻ���7��Q!	��&�dZS����7��Yו��i�!E�OaVM>O��J�k��<4�w_�V�%]�Z����STW#����Ƿ����V��]ڣ^�fwi���"2��.�:��9��]<PB�Ȁ�WQ�ࡕV��U�y��XY���a�N�u�H	�YjCLP
�W@H��B�����/��7�@��pR��an�!W�� 2c�R�ęgI%ʠhĭe���e��e�b�ȝ�.P�pa�3(�t�cIըT�� ����oy�f%�o7���'��{�0-���AH"�j՗#I$Ę��8K�b]Z[r1��ix����$UXŻ�m��ض$�`�܈�A@qe�B(�L�Q�U"b@Z��V�%K�+`H�$�,P�{�^1�����j���!t���%�t����u~e���M�C����)W}�h�!�ѽ{p�
�I]�D�sU=����חo�a�ũ��#��5ϳ��p��\��:����%N��/W��mILq�� ��#+�b�e������i��^ܸ���
1���֣��\{8�`q�bt�=ڿ#����ҭ*^���@�J����t���*+����
�zH~�S�ܐ�RQ��Iۼ��9<�8z��.���<p�u}Z�x����u__u��B-�:WF��	zԼ������"�_G���9$��>�B�
�ԫ~�;X�����FgT�=3���?O{����������ZJl�'k'�G]Ğ��zP�����P^Q�
怋���b�e�;.��t���FV�0��~S�zs�Q�*�N�$�T��p�3�-���G�zu;���G
�.-\����g�7��,�v&�`$Jt�\	5��n+����h$q�"#�X�17�-�UHf@8�!�To94?���O=��[b��8�5-B�^Yx ������]�q5@뱑-n��\9}��՘.%����<CVcӗ7fR�2{y�)nk�ׯ˘s3<��~>����j:�n[z7��դ[�3jV���;������,r�7ړ?��z=|t�,Y����
��:�]�⼳��^p�R�(o.�{�u�KI�H�b��VJ��rU�e����+$~m��ԯy�[��R�-�t���{y`C��o���9RZ�,h�qج �[7���t��v�%5�կ�izC��N9}ݙ�C�5��ޏG�sV|�t�_X>�Ύv��ٻЁ<��g��#83�����wEк�X�O���"���)rԌ�q+	�u��P�_ź���ʧ���e��X�Ъn�uM�:�'1pɦ�en+�8��2K�]d¨涡���r�-dQ�)���K�e,�{-]�%�~z#���M��/��1��r�/�Bq���1N6e_{�Ë�2c|$�+��4��� �S\�巁���q�7^�Ν������ZNQC�Ƅ�..�#u������o��pk��6�Ҭ3d@޾/�;���𩊕��xU7cչ,���=�=V�Om���.o\��au���F�<T���V�ᗴ��"=���_�������ua��+���$�Հ.��4��^���u%�8R��L�󛸚�Yq�o=��GO�{%^��}ٴ�%��a�>�Ag] �nQ�ޕ!�2-7���g���a�F����<��<"�M	�q�n�9r��	�Q�H¿#�#�U�t���? ���)��m`�7/���c��}����e�_�p:Rj�֜���g�)Qv3�����8<0ЎL�璽�SI��x|9�yN�Z�(�`�&��F�yK}��k��l<ƿ<�����ګ�(vQݒc2h�E�t�:�U��4������y>}�ӝe��zH\�ت�/��s�y��|p����}0��X42�ݛ�s���AP>�/��MW���L�9a����ٸ�e���ܤh7�mla��9S�l�sQ��6�E�V�Z�,7�#��5iwȂ�.��y���Y�}բ�j+���5YA-�DN����cO��:�)��ݮ1�N�-ј�e��{[.�X�)��a`�u�t!Q�	36Y�`!�j�f���Zʷ�R��P�w۶:�M�{;fEn���\@�p�\��J�N���wڳ�{YzD{銹"H:�*�@E�]pn���S�w�i�[nF��4�z9fevm�{΅��y�_
iԒ�2cT���,k0P��[�C1n�^"�joQ�X0�m*thP%�R���F�][ȣ�l�u�I��XTU2cA�!�%��B6���+�L����5R�2���B`�iā[1d�b�Լa��L���(�>����$�&c�V�r�Ci�wQ�u)A�,�4�8��#,QK�#rTQ�2�]q*"�*,�ibciKLK�j�[$T������TETiR0X~"�� vw]��f�w��#y{̮��UUU�NO䮽���أ��Q{�?EI�������� &�3�:��51O�sFo�}m��v�+po`%h�7�M�
�����γ�2L������c�Y�����O�b����]�,������p��\��V#@#bݗ(T�=%���7�c�U}Y�5�ޡ�4#�B؝Ĉ��̩ز���Dz=�K����M����ל��0�1,Q+.����لΡ����q����n��{;찄�%x})s�Mm�^����Q]�pT���J)dwc�f�it�f�]�]�k��^gΖ#�4X�[E�H.��t�Q�&e�v}�{��>�����3�V�!�u���h�L�G�q�;:��H��W��J��`�s<r�}�J���Լ����8.Kz]e�<V������_�^w�e`�v�s�X;0,7S�xN{k�4�2�_��!�jO�}��;/s�}Jf�O�%˳u�w�攰p����;������/��NH�p�~���\eZ$�v��L���*ȷ�sw�����熎���qi�V�k�e����ʑ[�]�^`������Nd�5"��68Y��V�fٝ����#�;v�իU�Z�J��ykIu���x��]I�s��~���z'�H0��u�A(���@����2��w�o�����L�>��u�ާ���{�1Ъ�P�UźT_6b��)շ����Մ�J��7��4�(1�Z��k[A�,]k�z3��Y\i5�o�ka0[�un�Z�{�)�����9=��7��e��z�9�;1s:�� �y�����#��_�����=�	��_g�
���3S���B/�}W�f�u���A�7��Iߥ�%Ӗ�F��d�	�\	���qu���#j�j/M���3ޝ���I}𙷇���|O_S�hT9��o˟���Lo��"�?U}�}Y�J�쟏�����WZε[O��8;S��WM3��;�]K���]��Jy0�m�F��ٗ����s���gZ�A�a�YT6��5��7����&ZP�~���ƶ�{a���`��Q����������]]�6~?;T�Ѥl/���b��'r���c''�L�@W�1�s�f�� 8ڥ^��\$��ٗ����|�;���n�/��wz���a�k�҆�i�]�R8W^q�(�+l-K�z"9��aM�e�|5�'&�K��n���fWLBj��[}ۮ�I���y�s�0:M�C(G^���ƴ�]�Η;��Y�t�%��a�Q5�u�^M�o������Zчm֯���O&Ŀv�٠G��@�hzjՕV<<��`��n�b�4[YN�y���k\�0sFy;�p�o��ߜ�1�xƭ�r�j��Ø��4G�|�6i'SP�{�vc�'-f�t7��߆�:N���#�q��rt.��TPk\��r���y1�u���mq�}���f��G	׏��SOS��fܵ�O!���a��L3�u�=�q=�V�|�O;B�,jrg��]��/����U�V0`����&Vݓ�k������qH�>kY�&�25�v��n�ȕ.u߱a��ե�Ֆ��t���;�n4a�n�^�f������:p�8U@EP�j�6j�h�	�.�3��%#6r]J�_,��%An�6qFr�o���=��mv�Ll��u+��F�[ǟ�N��hʹCޛ��h���~���K�� �����Åg�풔�!�>�mZo�	����&�ۣ>1{ｼ�oSMdr�be�a��zV�O��U�S��jf=��W��I^�������� ���0|��Գ���P�D�L�SI�ݷ;����Z�yb�q2�0�F����f�z�<ֵ`�b�T *������(�3}e���r[���4�F1�])��6��^���ED=v�epeG7V嘷5��+:�`{$��lP=���2��Q-���Zy/5�d�_SP���Y��d����=��<��`<B5�h�e��I���F�3�o�H��L�n;�/r�:�3�K�!�(��N�ٽ�g}
y�]���j��e�r��
¬������S۬\¥Cm̮��*Āy����*�r�]��}�
y��`�Iz��}z�D��]e\xI0֮�݀u��
�uy {ֽ�X�5����k�:�f�#>I-��܃7�V���Jzxl#v
��j�mf�Dq�];k���nNH�cy�|�1@]\��t�IhM��8ɛ�)�s���].o/��w�j�ݦ��dwrgH��3[��{�s���ҋ	% �$ZbB��Ȃ�NȢд*��-�Aثd�����B1nD-��B4BH(�M*BTnB�H�҈���"J�RH�j$a(�"��2��2LB)lĂ%�U�PUQ�*(�DaT��H$)����������Z��GV��ﾯ��������߈��OF���o�m����*��V+@!��խ>�Ct�)ٮ]J0���j��f<��m��9�u�m�0�t�ׯw�^�]5���y4��{��I��Zs0]���֍�w���xͺ�:H����<��C[Ŝks�r���y���m&�����v�&&�Jʡ��<���w�BӸ��Gԡ�E10���c:�)t��[�|�b���{SuK<P��*�k+p�V$P]���we��!��z=�.�qFvWЮ+E�I�-*�������n��L�-cP�an�vV\���3}ޭZ�ᇭi�Zo�Om�}������J��N�x��Э_e+=Zj�hB���h

�0�&9�^�����\ܭfh����ְ���O~�MmÑ��w{��n���z���ڥf������9�G�p���x��'a���O�y���c�4#EO�Tk�ɍ��1��j2&�7<V�̠��M��hJHu_M��Cn�W�kR���Dw~����~k�8a���;�o8k�C�|��u-�ܗ������KCD�W�>�3}�`��5���o3O��㻼�]��q5�G��&S>����";4l�[kܔ�ƴ��e�z�k�·W���e����y�r�S-��սѧi��-D��5֌8fqux��{�����]>c��޲�5�P�g�B�C��fOr[a玮�d��o�p�^D�F��t�Y}%s�]��c|g7�g{ȧϡ�v�u˨��r��M�ph#\Nn���۶a�0"[Dk�Zi�3���4�8��B!�
�Au�vz���3SOP�8V
�V��kf�*���57U},����Zhk����;ԭ��!�q���f{8�Q�&[M8m�5e��X�q���x���k�r�q��k9ƫI����6��_
�J�`ݯ�9�euN���v�b�,;ֹ�HI}9k{	�ӫ�x��U��ݭ5�ڳ	�\5���˴�V��������^�\�Љt��\�jk�&Z6}���-f]��y������	�L���=v�cG=��������4�K�ۂ2�<|�R����$�v�v��gp��Qh�����&}f]'���7�cR����w�W���~����J3�Us;�z�D�[C��\��D�\�,�y�1��aN#x8a��,)�̖2���:r�0w�_W�◪�1-�>k?C7fh�Ӻ�3��".P���LY��;���˲�rV���Ǝ[��η���5�C��+��l4Y�����1�!��/7Aϼ*'{5x�{+N{+	�ܹ��e��o2���e0��'!�dױǍ[U�@�Gt�b��f������W�M���h�>c4��g�)Y��xb^���]����Yv��=�<��|����;��0(Vq��,}O<'�w;0��S̬��I_f��V��\B�<񭵍��]�uT�
�)���V5,�T����	Y������6�w����tJ6�2�3�Nw����y<�N��4�>��K�����sOF��ӝ��<�a�f�k]L�|�̭�56�04cxƳ�J��^O&��zCɤ�a���W�5���U��):�֟L9�M��)�`�ݞ0rc�ۃz��Al�� �7;&�H��}�&���b�������
hԶ�3܆�L�I����E�=�,����D��Ƶ�d̬5�˳�;zuz��V�=L�]hj3�'1hi�A���LA�E[�W����,���~��V0Áe� X�
�
���#H�3[
��#��''��4�qx�̛׮�&�<�!�����;���osSz�ާ�<�~�/�]���
����]+��k[y
�;
��9h�#������eI���ַ���8s�^�l�:�k8�w��������	�9�op��>�ѴОb:��8MLX�~�|�Y����[Ƽ�Aw���}�9r���Dk�n{�^���}A�2�ډ����6�ɖ�'�se������{y�ך��k����{�ÞƂګܮ�I�����{��Zz�v��V�S	��=�w�ߵ���q����i[j<��)�!�睘�������G�kj6aO�m:��M�R �z{��o9�bt�t;MnVP�f\��Q׌��o�m���(��K�FZ0��q#|ݗ�ǈ{�Ƶn����k��4�y�{�1��:ք��]p�_&�d�7��k�Z����5�����f�9]Ngo��V���o6�îB<|�k�՚�#�g�oW�n�	漗�m��'��OP�9�ޠ�S�|�����3r`v������Rڄ�OJ
�� u�Z7`�!�y������Vܘ5k�n-��L낮��}wW��4��5%����U� M��9w�i�f��d�ɽ�AݑSq�k��I�8�����<u�L��v�l��#��b��e�,�.�t���Mmn92��1�h��l烓���-pl�G۩s��P��Ld�X��H��i�}읃���k�-4l��h��%ި,e�ǜ���0%���j;�.���h�P�ܱ���:ch�����#�e[b�N��J��y+�7[w��+�ԙI�,�tVlǪ��Gn��=O�8���'/Y��i�0U+�����<����l�b��Fm�+xp�b3�+0)F#݄x�4c�(��/��2v�e3[¶������ׅL�hf�5��MP����]�[��D[b�!F��Ҋ��"1�0�iPDccn
�"��H2(*�(�im\dpƛ���ҒTc-*)hȣ��7)�+p%HFD���B\�TR��H�[X��d��"�D�_|B4h�޼>����XR����Ԓ9;���y5˔~�&�O�&����Q���/aʗ9>3�!^��x��U��^'��L��k�V���}�i�cp��B�5x�]�zVʦ�&_<Mu���Xߌo�5�8�\�k�Y��䭵9�o8a�i�4i�^Lۜ�5ƶĢ5�;d�g�ve<��J�E�Z}^�����{,����bB�Q�+�����ڙ��&�M�c��K��ju.�V��px'#�_R��]��Y~�������ҟ5ķ�ɬ��e���W��=�Q���OJ�|�K�,�u㼝׶m�6��X�16� /���]���pC�}��,�8�⫭4r�A�4�*Qg��4��Q�h)�J�W��e1�[n�5��˖��[K���u+B{{�^o���k��5N_�]��ʾ�Q�������o�T�&R.��u�D��|��ٿ5���7~��V�#�`E�9��ܻG7�_	�r�;9>*�����Yt�p�TmUW�I���h�)��}T	�����-k0�9ji����i�f{�漛v���J;��B4{n��m�B;f�^cW]�8�N]�z��\E�x�H�8p�Pߝo=��4u6#�Gm�n��k}۰�ƸVF��N�
R>~5�G.L#r���a�k͸p���!�����5�>@�$��U:ׁ5o�NoD5���G⫞�ߓI��L�߮�̣2Vo�&$rd�M����Bbk��7�
�}�pP}��)u��*a���玓.���$�=�Ʉˤ��OCI����Z�ލ�u�������桾J�A7����[�6�2��m��w*���9���GR"��l^��M��V��>�\(����a�*��ib��ƩY���D�[k�釾���弳ּ��ꚵ�8-�{���;�R�ʏ�Lbk�G��ޅ�9u��>Ņ�|��:L�֌R˕o��|��Ul�ӛ�J�Ka�^�C,[��C�YL���^Ռ���"I�x�L�lvг��7�=8`O�_�r�0�TQG�-�g���a&�Od[C7�����!z�%3{;bQn�/'��A�v�ܕ�N��9�����?��%$�n�a��}cO,Oն�
�y����,��W�`�Y�Q��߮�j���``�n�����/iJ#L!�N�Dd�,����GLP�
x�~D�O,ԍ�x]�f����]��hn ��cat�zF����M��)�eė^ k�V�� /�Z������M:o�Ǆ��&�N��P�aa���gM�������h��b�o�<ӿG����A��{_7=�io]����lM��hB�-��7�1.���^;�F��$-��#�*�=#t�buo��W�;�����jС�@�$*'�wvI�W��U����e�M@5���*���*G��"�{o�V�'�W�u�2\�6�-�>�HX�ew�@w�2F���W �6C�|����􇒛n.Kx^k��݆`�q�Y;�2�E��U}S���3��T�=2�n����m���_�N�d'��t5�S�9c�AG�Vl�B�/�Q;��*�7�-��d�Y��pǾ��)�g5Jx�Xͧ��õ���o_�^Yu���e�� Ʒ!�/�H�<���*�w�������~_&��ʉڽ��<Y�S:W	َkܓ�4�d��^.64R��U���'6m��hj��{��.��a��J�[�����}���p���V7��;�}������ٵ��9�Ká�B�R�9�%m�dy�)��t�U����LԮ�+VOY�`��w]��\�Zy����ۄ�V����+���ڍ!�kb*8^�x�^�o���M�
�Z�R�&%��-�	�帲�h*�%���&*7W�vT'���M�q-; Jav�0�2�k^�Բ�$9*��d���n�H�����#Yx"��dVe91����\��$�B�3����vF)Ua`��G2ܖLܩFdp�r*��x)�V*�Z��̢�+��-H	*� ��J;v)��+1�F+�H
+�(e�A]�@�r��ċ*�^KDYX�W`��Ыݟ���.��%Z]�����='YOW��u��Z�#�G��]�Z�$dde�qF��իH�1,ii���hV��a��F#b0�.֕E%��j�6�[Q�H!p�.�T��TH������Q�I�K���]�ƢH�jأ���Yho^"6���I-�۹-��v���$QM��yJo8�k�v�66�iݙJ�������<"�7��;؊WYG�J��	r���}.
'{��]W�8��q98��حP�q6���@����#Z=������' U+���n۔�S�
�sRgMr��J<�sh�|�����ee>�ئ������L���Kj�J�٘N��q^�~���#[�6��K�M#��b�9��ҝ�p5�mdHt�i^�%�[��WF`��B��'�tu�~��y�Ɏ������CfY�+��VEFL��a��q��Y��t/+�w��o	��{^^#P�w^�,YI�mEЖ���9D�ݫ���}�~}�8۴�2{��Ǐ7�s��O��O��#)��)��!w��I������$�P,�yw8СĉyW,Ǯ��㗂r1��n��7�m�pǫ:n/,�{�O&>�u:GJyFT� �F���D?�p�\]I�#��p̆�u��Uj'߾��Ie�g��5}�䘱�Q�Du)b�W�-=8�Y���K�n���yE0���|A�5|���Mv!�Ҏ�_:s%X�wN�j��]XŪU)�h��8.(��w��,�-V�H�u�6��_\����K$u�Nr�p���靫8�o��\�����~t��aᄚ����t�wI�{�ວ��|^.�жjtowy�G׃�]aI�a�2��}�ں(F�6�$���e\H�-��o|�f�֋����[�i�s8��H1�fR��i
�he�����4Γ�#�t�TW(�ծ9�m�-Phl�r4�r�7˗ވ��uv�b�����_�L�5j?{9������3���Z�,|�]�ceo0�;�#Y�Må*����⤰Ho��{���*d9�q��<�M[ƳA\�v�K�%=�ø�+o"��=W�AT���43o7}�;���9:�Bq���css��x}tY�,�����N*�vY���Ywg���ou�2@�����,�sг-�e�<���J�O;�����;�Ļx�H(O��	5u"UmN����yXX��o���|mb?zg�R�;�J��egi��{�����](�Ze+��d�+��|ӌO�W�u{����t�;��֌cL�,�_��~lvi����/��b��00"C�^W�^��PQ'%��O7CY���1���ڻ�C6>��y��-��ز"�!��/�+�Y���Y��'#{uS�zl��V`����{l",�E��A�a9#�3�^������$�G ��}_>�Ҳ~ܧ�6�h�t�\�΍KX�?.�;w1F�2^��B	�q�Da9.Ҝ��S�^�D=4��c̎���ͧ[��͈]��~���U� =F2�n\����|o��;h�<A͡N;�]�۽{W�B5�u��9ۮ�o��8('着�OO�3N@enB}t�O·U��ٸ��`��گ�C)����]�AqһudM3p+3W+z��Ob&��[܅=�ܬ+�-�A��D�3�n��^���F5�����v�w;nEۊ�x@���h�5T�Ί�b�r��f?t���bO׮��vE(pI���~�7�Y��)`6�f��Ս��n��'K�ŭ,k7V��8���V�����R�k���wn�^�2�6�NX�g*�Y0�"N��ܛm�-[꩛�f]�]2���M�wŌ�<��m���d*�V����#�%��хS��7������\E�Xh�Y.e�$o�h[r�1�V�hc��}�U��h�U�rg�,ʉ!�Lr�"c��c��E�-�]�Ұ�I�*R���N�ɘ���t��%f�0j����Y�
/�D�I���0�ر.��L�Ӥ�YM������+Ǌ&��a�wz�VQ�Je��e��v�"�6�]0��A���B]�H�.�T�ʅ�Ceݥ�"R\�Ĉ�FLbY�rZ[b�	 �`��n�"�FV��U�jƭQ�����h�iA��ET�.�Z�1s	#L�v�H�� !IB�  E�/�EhW �^,[�".%��F��ً.��hQ4��)�0���܌�oyr�ކ����*h�f�}V�M흙�*a��yIn�Z���:yg�>��LۃoY:�b��,Q��ʄߵ�a��c��6�]�6��w�K����[��/5��c��y�PgV��V��!Z�F~�9��$�;z\���̮��w2��Ք;���Ϧcc.I�#�y)�}�7 �l�Mb��ʰ��|}\��i]�Rk��J7�!�ys�1��Il9��"������y��«�Jg�:��8��0�s���F�n�i,�����|��슼G�ֈ��VX�A�eo2�.�S�����vE;V���ٝ>�(���}�r�v�9����g�fΈ����^.�A͊��N��TεG%���\�K3`�j�X"�>�6ò�򾀝�<�s:�#g�`@��Εn�^��F����wL�҅߻NE�������ѻ�@FGu��	�F!�ӞwZ��#�Ngթ��_f8��j��t�ط��ϙ�X�*ɏ(�����F���]H6 �p+�vr.;�~��غ��[t��Y�/����?sƻQF�X�~���@�ؑ��6%�+Ua"Z2p�
-v�F���&툹�ȫ��s;od����Id���L����&���+�]�P���eh�γ�5�R�n��E�V;�S�+D��=��f���R�{2N+rޅ�7�{�r��+~4�i�^S��>��
�j=���� �:7�6�2rx�1X@j�U��H�藅���P(aI�C��.�2���`�ٕ:6��W˒<�ừ~�/7�&�.��n��'�\�����ٚ3-d�9/���I���<�T{=C��1;p�훘X��頍�Ġ��|z�\h�l��ʥ��O�j�
����$OE�t��=��1s� 7EC��K�ּ�㋷�dM�bk�t�np�cEZ�<Ӿ�#n*�A45QqD�ؘs|-N��Ȗw��ڝz����g�x�䥃�)�ӝ���#��#�6Ҿ�P2m���j�^$�%5�"v���H+�egm�u��s���$� V{��:Bϧ�s�h:H��`��k[c���}���eDW녾��|�f��y쥴הn��f-�n��%^���x��mQ^�]|���ۀ�s��Ֆ���Y���A�O]	�hq�:�p���t)�V���+�u��7[�xi�S����q��U� �<�Tp��U��!�-��=�T�e��.y������Y�v�b����GF3"���D>�#,VU,wOo0ثt�P�����t�/$�P��ڑ<�;c��Uǌc���޼�Ɛ��2�8Q^�T��t�y.X�)Gm\�e���|���"_�}�����ϞN�ݻ{l�2d��D:H��p>���2/g��|kDͬ7�:��ާz��d[f���t=�5CS�ȗ�{pW_Y�ա^�]yC�=�@"�Q�ԝ����l�q�Vmj�YC������\�'�u�gLC��{��+��ϊT�ں�Sޱ\$�V,yl{H�YJ����"�@�{�E=�m��9gP���5U�Cz�����y5>�I=�#F���g=���kS�7ò-Ω�fk�Z�[�{2VAR�!�̼yx��v|}�;?>Y⯭�b���8e�e��l薌7���C�ath�%}�1s���vp3n��)��M�=o*�+���1w����Oq�]�q�\y��liR�V���Mr��Kl�?,�ш�&����E�e[����
G9�8�5�]B�6*��$���c���,A�0�X2���(&@�1���F�0�@��4�s]�rf,ϔ���I'z�Re+�R9u����n�m�U�Ȏ9��� m�?A�h�+n�Z�Pq%���x�	$��+l$��
��"F�e��%�w)�.H�lW�+�l���D����,q	$1F��%[1wxeZKn�"��Km�(��!Kj�E� Y�P�-7r���2�6AЉK�DZ�h�,��e@��j����^�_^���:�쏇tv]._���f[�y1����Lt�V_�N�M��R7�*׸ĆlS#8�+����p��^����fO\^?�Zs/8W��w~�opn����T_���S��Y��M,�{�s��Z��f�'o܃�� ��@�a�a-�Z+U�v�6��x3룇;�wĝ�Du��]���]/���{,��6ʞ��!���X����*P�f�#����$D+ftO:f�����7��8/uk��F헮�c�ҥ��R���.eO�j׆��V�,��>�YY�t�y�7�Kp�!�,�N�c�!Z�>n���ld���
�񥶟>�4q/޹O�L��6:�� ge	Wڻf���d��[�9f�$�uq
�q+9���I�暤�AU&��wJ�8�����:x�a>��i�ʐ�N�n�+{O1��<ݺA��YAR���˃���Vִ/�]�L���ٍ��n��kcC���qآʞ�末g�k�M>s�V�x����*-]�J���k�H����h�%fWi�F�����L
�orvS5�AS31��ׇOr�{L�Y�O�I���٣����Ď�=��=�J��3�^��tMVqL=c9aW�+`��NL�o��w��c��*L�"6{R��� ln���=a{8i�YR���#���-�K{�Q�x�ld�)X�s-W���{5.y!��ҥ/f���'���oŢa��������[�ܛ�k '�^�K�zT�y�"����m�O��B�Z4r�ތ�μ�oR�1��u�%
�ٺ���(=9�����$8_v��=��I�c�YS_�v���ws�A`	�5���.Kqe���u���
����g��7/�U���e���HWb>��iߑ��?=Ssνվ���av`� NU�i��"�U���:��.���ܙ����wdf��d��L��,��]���W:o����B}b|�M5�4ճ���$bG����;'�[��>M9���	�2&�ʙ��ic���`at�'���*�o�r���[�t�d�yha�Ս���.u5]R�,]\8(do��t-�y�4��]�4��*�:k;10�������5��:`���w��匛�%r�B�-i`e��%g8�Y�5dQT���];ѹc2e�m����gwD��3&*�Q��� �ǌB-텍VC��+�+�^���"P${�fu�I&�\]�M9�1��Ν�#�D�-���w����f@K���¢�Xi�e��Z�K�GV�]�}YBn�J]O��(�T8���WR��Bݫ�P`j���jf�K�j��ۮFT��ՙj����k8Ⲳ����z�#S��Z�[&�he�e�Wi��Mwj�T�oo;�GY���J��Y5�=%vk�jUx�ud2���Òf�0c3ԃ�R����v�O����6���A^�\3T�&N-�z�/��|UJ<v�V��X���3�y!/g�l�3+�h�l׆��^�����g�7�'�9ׂ�)Zd����"�ŖbZ��çoc�z�G~�.����I�Q��6��+ �$��f���K|6�ᖙ���n��]�E�-m�^��IB���ᝬh̩]л�aqˍ)L�,��ô5���F�Fof�W<�'Mӫ]��0凒�UÓε�X�.�)�=
��&��Z=���İ�i��+�)�ƽ�2�*%���;���7 �k8��o	 _$&����u�����+XY3�Գ�M��Xv�5v�V��!)N�ط� `�#���j��;F��i4��KuZc�:�.k�F6��\殲����ݼ�0G3{%5S>D:1=AG���E�;�K���5;��w��>�j�(H5N�4�4�%L%��$��0ČI��MIP��i�0$Ăb��I�#WũcWl�>4ZW�S-�_	?B�)�@01*�[���Zq*
�lai���&����h2[V�	.bL`��o)�0A��B�w�p��70�;�*x'�!��P���١v�\z.|s���7(^'~J�K���tp��A�G�/��L.�=Z��zNvB$L���RT�DzS���N,����zGn{�*�wk'4�^���)�����	�aG�Ik�~����tKg�]0�gw�#u�,]�S=�Y���e=i��e�ûm^�+6�>Μ:q�J��,�S��a,߽�6��r��!6��;�n�[^52�)�h�D!d�/$F����fZU��g<U}���6L+�L��O�����s�^��]h��{���w���,�Y��g��^K2�/�q�WJ�;�KA�ˉ}O��c�;S=�A:L�ݺ{9�~��sSu�:��)s���y��ݸqkM��[�IP/Df�%��M��}}�5��p������}���:xa�l}̜��yO���E^^���~	���ّy����T�x���z��\c$et�{��]]/f�l�fWWI}.Ӹ�r6�ެ�u�ӵ�^/Y�C��"ۉ�h/#N4�����r�����)��TJ��Ԣ5�DPua���P���E�ױR����p1-G�Cn�XW{6�;��6�l'��1�Բ�u�|5f�T�̞�Kof��B^v���P+z7S��X$�;��25��.�ǆ��@aU4PD�*]��h�`B�\���C��]gS��#���oy�HKnDѽN1;�1wO`չ��Cvb*.�ٓ���z���U�w�E�ސW6la�<5Ѱ�ӧ1��Ê�q����o�4�z��2���+y_r5͈p��jF������M�V$��~�=�ACͿ=��c�^`L8�4՛u3Ŗ�I�^��T��mŎ3��r��|χ_X�.��fwD��n�t&E��C]��]�זx�GbZ�2�p�d�=g�}�/��aY��9d��H�6�t�l�z��މ��Ϲ�)W'����v�Zz�޼���uv1ܐ ��W��W�G���=?~R��e/#
�\z����}�f��nY
Z�Z��tFE����O3���w�������dz�p%c������r{�s�o���j;�1d��j�/=TV3 ���ɉKn���	�&fX̊��1./<��ھ�@�E/5�P��r��"Ӵf�>���촕rL�T�7��b*�#��Ϻ/X�˝M�H�5��o(�A�JXKl����}i3�Sݑz]d�|/���,]Nuǳ�|��W��`���*+���u^��yn��t�g.zu{F�4<��G��4-0��6\F��K�/�.ǮR&*�u�ޞuv��#���V���.saВ�K��[��E/�ojX�Q*�k���#���⮤�Es����;�c�jwceZ��1��Y��s�g����70] ��d��+T5�I�I=�p�%�eaPp\��3�V�Џvwe��|ރj��s(C�K~�-�������֘��i]�2B�}�1f����H��~�G�~�*~P�UU_�D�QUUUl?_��*�^�zK�PU]�{Ag��a��f�Ӂi�������h(�����ٳ,7��i�ͅ��!�h?~�~�5�Y�Y�!�␨*�i�_�5�gfkj��Z>�W�����z�����U5x��Q���\ oS�U������BU9,>��wX�j�*����3�m7upc� ��x��� *���bV�G���&�����`{ڤ�-4���o�:w��@�8w*
��������x+��g�%����U#2yZ@��]pL���C]{��tb0�n�G��-4�@����*
���.�I�q�M�((�-PU����ӅZ��(Mq��f��{T�6Lt�ƃ�PU]-��$�-�2k��]���h7$��)pK��@�f1�_�����}�'���_����N��@EU�[.yb��|pO�p���,]'��e4s��-��q�������"*�-@��]X�iC�o=����sTWS���0���1�y���\(DzI���C�GUj�J���?p0ayBr�bW*�����^T$AQ�,�
*�`���0?�B5�G��q��UU���M�U��4+��~��1%	����Qt�?h5mQݙɎX@���
*���4��#�0�j���w��V�O-@m��?#�h3�i��l�rJs�4�,zP@P��գ��DBw�x�i�)�Ix]�~$�
����]fQ�GrL��>�0�#ܨ*���B�l`��}��͖��<�3����C��:Z�y��I��K� ���8O<`k�<�4f
ۘ�{~;";��f/sg����UAUx�6��B��R)��`A�xI��9���2_�ӳ�p�	Qz��EU���`փ�<_w���n�AEU�;	� ,i�uuH٭X�+�V�t�Δ�dĂ ��БyhҎ����.�p� ���: