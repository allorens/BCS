BZh91AY&SY`S�d�߀Rqc����� ����bH/�T    ��QJ�XR��V���Ҕ-�e6�J� �J)��*� ��hQ�J��M�$��Zƴ(&��kj�llҪJ��M���飢��i��m�"�T�6٭Z�Md
���dڨҤYe	dQ�T�d� �UY���4U$T5�"S6��`k%�� ݶ�ު�,�6ll�C�!�\�U)GRm��u"*+Jje˻*ڭj�k*�+cZ�k%EB2H������mcmV���4��ԩ-<�
�Ħ��A@ ܼ���c\�vwu�U��t���K�����d�U\�����4n,��:t���&��5��AEnՔm��V��t�թe�+ej��mkW�Ҥ  ���� �Sq�eA��k,T6ԭ�\ �P�ʔ 	�ܠ��TRܣq@P��sF���t� �g\t���5(���af�Sbix�QT&�6��U ��
J[��v�����R����ԪeR������y��z�h�aol�����n���v�y����v�kZ�5U����ֶԵ���ETH����JUu�=#���(z��� �K�릊�/8R��A�y��� F���҅ =�: S�/r<��z���@4qWa��m�Tֵ��j+mm���*AR7{y|�= ��^�B��/<z]����o<9�S��t��cC�/p:���U׼Wm�҇��{ޅ =m��x{��f�{ހU
S�m���L�&�V���Ԋ�����}�J^���(:j���=( �K�� n���H�E��Ѥ���]�� =� wK�+���۪pk�+e�U)�+Zi�i�d5�杖 n���d�R���]��f�q�U*��rwP�*e=��(
W�{�:���n;�� 7)�`WEw;\  v,  ]��U%�k!4m��$�����|@��p��4M������ �6��FwW  ����ۨ
��� ��`h��;��hY�m�R�Xf���7�}( ��>�]��)e
 ws.�7V���� �)� p� ګ�@�`BwU�5��h���**dU>� �w�:(��p ����f,( M;p ��E g   @ �w4t4�� >  �P�%Bj`�J�5F&�z��214�2 O�1JQR�  @   "�����L	�� �2`�0�O��%T�       e) F�4�AG��Ѝ�A�z��TjSICTxSğ���   4?O�����[?��M?��G��f���wu���>����׼�;�u�G~Ú�9�UQ^��**��G���.*���  
��v�����6����߁�~�~���w������߼�X��"����U\��
����O� Lچ����6��|������_�����L.�͑�`q��Ge�0���1�� �\`ade�)����@�@�P�@��000�\`aeeLdcL!�����C\aefLa`ddL`Laq��W2� cm�q�1�1��P�`1�1�1�1�1�D�T�.2�0��CCB`����D�����P�M28�ʛaedLaLeL`�CGWCCM��� �G\aq�1�1�1�1�0aLee`L`\eeada�CWG@���P��&0��"��Cl��Leq�D�
�� �2 8���8L c ��".2�08Ȋc ��0�8��*�0���)��&0��c(��0�2*��	��0"Ȣc"	�&2��"c"��UeA6��
����2��Ȣc��	�Cev�c!���0(���c"����Wd@6�c !�(&0�0�2�2m��L�����.2����#�.0&3�Gav���+����������8�L�����La22�002!��22����+����������.0�a1�1o7��d�o	o]m~��`?^�o�7w
��*���˽Z�3r�(��۱��&)��B�Jf��/4?�+��|6��>(�e�@�%�O9n���u�a��PP`b[weƯ��vX���J#�Vpᬖd$Yr���L�{?d��h�{��s�K�p��b�:d���/2�8���D��m�a�����������K�t7v��7[���(��{��Lk
Q����E������5ZCn
6�V��e��n�$����i�]�6�%t�f��"9���]^�7V,��oF�nY˖Z�����B��1;;��&P<����-�ǂ�A��M�&۔�;��'��8p2R�w$�;H͕��;��3sLK�hP"��R�Sȣ�����N�j��pVSWt�ËI�\��f��us��Bi���f;eRQ,�'㗵#�j+��22�V�0ŜF�n�Öva�ś�v��F��T�c wu!�T��\��Q�x�R�1�l]^V=��)l�9�I�r��=�s�wWv�ä٠B��9����[E��V����YOr��8࿯U��r�vr�Иn���b+ae�[+,��T������H�X���0dm�N�^f��+�s�L�G�eLU����N��7f���{���yͥm*O0a8�m�)��M�I�Ȭ�5�if;Pm�a��R2ʂ�����Z����j���e�wZoO���&r�]� J��Lk"迵e]-�\�R�Y�[E���"�H��⳹�Z���0�Bmh�d�Z��b5�5Xkhe�F<2ջ	�� ��մw[X&L��Owږfe�gA-^j���CT�cś�*���YgZ��Y�N�S���͠�v��0�A[q)�&�4��$��"�؆�6�_���s!"��1i&�{F�Xy�1{�nlu!������4(�pt˙o��CD�6d����4�����J�R�dW��n;�t+ZƑj�c�{��̦7�Tܘh8vI
��q���g;b���m^:��6�jl���0�O]�s]f��{T]bl�-��<���`5a�����	V�� J�k���C��/�ʼ�X�i�٤]E���b/p�s(L�J���(fY� �@�P�o��4�,�;����*
��+nMUKp5��]K�F��5Y��Rt��aQaN��4�+�X�g����AF�ރ�c,�eAY#�+l�W��`��+��q�P�-�*[�����E7�X��sY�0U�V�U���"­5��f�����R)��lȔ��,�Sta|��Ѭ��7R`+N١4�fHּ�z2<�0��{gt]<%)y��̔�([s[5)�L���K'^�kc��fi�
`��R�B���r��k��T#�yq��3JNQ�9��x�wWt�DXj^��7K�Y�w/%�
FjصJl���h;Ӭ"�0�Ց#knTәw+H�/�NfR�&9v&<!ks[��J�P2Fo����E2�c����	e��

��w�7�c�+]��6�N
?n�8.����)l���o4�в�^�.��v!�����������Q�t&Qhz�Դ̛7Q��=a�Q6ޔ��K�����;���ʝ��LU��{i���՗��a����+"�ٌ�PRQ՚p]��E31V�32�j�S���c���*-/f?�����7*P�{��vm0�X��O���E��L�R˦le8ZPͫ[�0��MP��ݓ���n˲.�y.�Vɕ+ڸ�AJ�1V-P��eRo���'x��9-�`e:�8�L�-!l<8�ݡB�������6���[�"^-��aF^�O(JЙ��9��/F�3P��z5�i���Nj�-%�@��525=�;	����5+�x"{ �*�\t3wVVeY�&e$D7��D&mCd1����#q��b�m-��=(;n^CX����r��qL��yJ;)6x�ofK2a,�׎�-	j:��f��<��%J��C��=����騰P4�
ϐ��d�����GsVa{�A�gJܽx��KKT�Dy�����cڟH��ئS�@�@�Ψ�[(`��R��ZYd$U�qU�@������hxú�z��2ɷ�ml��E��2K�W�ZR'��*�!(n�ï2��xbu�k�QA�=��s`���oeJ��:iŊ�ݣ*e���d1&�ۘM
�ut��陴,���PR�&&�[�61nAWv���0����7鐧�Z	�v���\-���rnY��n�("�o&zn��ʷSn ^L@�*�:tqTV+Ƶ�KF�#�M��-��u��o���{��t)�c��5�2�s�R���
����so��4Է%cS�A����'���t@T�AU�FڢQ37������D��T\�&��e�d�淂�ډ(s~�n�MڷBhuYB� 9gvc;SCB��W{4mʘ�3l�OjG�Q�x����{P�v���HX��f�9W 7sJ� ���f�(�*d-���Tv�İޓ�Bn�]'ccr�F�P%tiZ�m��)��FE����3QK,�GsP��ѵ���+T��;[n)��b��Z7A��s@����>��D�ne2-�)aFk,�"��Z�2��jvm��n�5�z4ZN>����#u�Il�Q�H@@�`r��@h��F�%��hV�G@ԋ�t��~l��4K0�T�Vfպ��>�\@�wh>�t馰�֠��{��v�sS�K+.,��dK&)T����Y[��q��<�܎�'b��7n�f��<vkf�� f�e˶�tU܎�k~-9�R�+n�yAn�n�u�\aide��&èv�-�P�+��-�#����2�ś��a�ʂ�m�Z�M#�yL�v���Qe6u��w��)������gv��࿋��! 6L����И���iV-n��[
���xnQ�Ȉ7� #3�kj���ͻY���d'PҠ��C`�Ř���bT�V�nR�\�ʷI�e)�l<ڧc`��]�B��6��[>� wy�36�l�X�Yj��+)�=�h-َL�Ho�Q\�6��9�"�7hV'���+v㝏�!������V�b`��MÌ<i;v�V�ӆK�����3^��.d����h+u2�e�u*�U�P1�S�.l6�Y������
��e:e�"��eи��J���� ��m
��ķj�:8��d�?�x�W��AZa6հ���oL��Q�1ޕth����q�\-�D�ɫq�[V��!���z �j�Gs��9,yZ-i��3J�+@X�i�\S*�T6~(nC�9�U�X��t��%�A�n��0L��myW)V͔	���j��5�6��'�:���+&�֚�C��P�,��M5�������[�`��@�� ؝o>�+l��NJ�����2��a�X�7D�*y3
�a�h0镲�u���hf�["��]ۙ�]���&+�����H\�\�R�Y�3,,�Q������6<ų0M�W-���ƥ��U���9m=��[�hF�Pj�u�h9M�iIT�43Z'[�4��fT9�N��F���b���Y0"�f�<Z�ɦv sm
m �i�����+����S̻�4Xɪ`�f���#b�I���K,j�Y���\˽�m%mI��J֪wm�*�l��u[���"^cpӖY��!���g�1�i��5&�Fӑ֊�Xݩ�M�Z��7 ���O]f\N�'
��Ci;m��e��\F�/w4P��ޓ�r�j_�9���s^�Z4A)�L��CSt=�*7L2�,X�r�t�IhM��XU�@�Ų���6b��ԏj�(f�c��pXv̐�<X�_��q��.d���k]�Z+^�� 1f
NVi�{��,)�+�teŮ:E'�m]��ZOd�h��,K�	-0�b�J<�t�ilo�H����IuT@��H�X�}����D�.�b0��<�XR�}3u@�C����K;vuM�6�V�.3��Vv��R�)�䉽�Z�]��l �Z�4�N��ؾz�;֑jދeMm��}�%�˪ͫ6�n�����R�N�agV*,����l[�0�i4�[Vs1i���˧���x���Q:�.�,S�n�sB�1*�Q�(c���G���:�د����z\N����in!oRdV��/^�q9��z]��e,�ܩS��2S�u�7Yo�m�&����8�r�*5&��]���8�L��֓XD�-��	{+&�U�Oe"S
�8�2�{5�z�F����Cm��j� Dѭf0%J����ڊ�K���Owk%�EV}bi�4��K]���z�.l�kQ�;0kY��0�e���+(^:KZ.��u�0�;��)�lX2Jw"�_ۧ��n�NG�9�Z$�6�6�цd�*�:�!���V����[������F^움Rۨ�j���7���X��X��(Ym���a��ڻ��ָzm������Y�u�k�4n*|��<���/5�&榎�y�ŝ��Ҩ��ݔn;X�=��e۬9��	@̀�X���g#�4���'ݻ��f�Jۏ ٧%�ܰ�]�Եm��Zn����N����m�52��td�4����r�ޛC����h��aXc�8�ݚx��̠v��2��J�P����,D,ʷY%&n"�騍�F����V����E:�C`Āh%G��؄)1��^5���5�sV@�T�[�BŊ��!����n�m69t��P�(�C1ܠD���R�%a��*�ŀ �b��Y%������� ]2��M���v��<�V@YF*7�ƺ��C�Z%�[If�ϭ'����P�f��a�~f^=��7n��<:��;�]���6��`J�@�Z����t�5]+���R(�1�����;g&؁P;&����<�	��;�X��1m����+w�:4��� ��w�����NŪr�q��b�z�[?56�܊΂r�zs��M݉d��f@��I�e%[�K�cчff�6���O�,C1,	- g����p��gu}j���S���(hsL͎�����X��y�<"�A�IM�2�/2�J�YV�wj��Mk�H4툌gI#��^ަ���ԩ��N�W3h>mK;F�dfј&�7g���^�{�r=%�kf�U�������R�26Z�D��˱��oT ��#��B�KGhaE(3�Ʃ��,X7L�.����ӘpS�2�"��fm�$˩r�H�Dcv���5�5m��%�� o.���$�Ok�*�$�S6h1ˤ��+V7�F�ĥ�6^��p�v�q�T�*�����iٛ�R�a�t��t���rɁ˲��`>�R�)5���4e*Ԙ���;�&ɚfC�i�+h��JͼYe��V�,�q<����

�;gI�d�S��]�gNY����r#w������2j�X\���<�z1�^ ːb�
�Sv���f�ե�,熦9���׊�����u��U������:j���n��mR�����v�����@k�8�yV�M���4��Hɐ������w&��B�]G�(n�,��J5[>�n���ޫ����=�9>�Y�z�hH)�fe���I�F�2\�>��׀��,�m ���Z}�)�uqҋd��-1
ة�oV����Qe��jl��P�YQ�b�M�so2�+a6�\�JembͭڟbHB�ڃ�ȺGX[�ҳ��9���ҳfc4e�Y�XFHږH�	���r��ZL׶���-��
H��O.$�a:(�<��ߩ��Z�X�&���S6�B�E�Rim~��e�J�B�1��u�p��7]�D;�5�m��cN��Y�e�Q��湠�/Edd��os��C FT�e��ǒ�Xʷ��jB�
��}�����d[��[��vn�r�D�rFkpµ�V��Z6*4�䬷�	����ic�M��K��3G����ٙ/,�G~1�3L0�Q�WOt֬�-�%UPԱ��Z��
��f�3١��Q��h�`F�	RǷyX*"0��������I."F��']4�]*�ua��B����^���� 6�bc�3Z��hd�����&Ό�n�]#2m�v���p���*A.�WKE��6�m�+� Z���r��l%Vv�#��ȥ�D�P�О6��ԮJ9xmŀ3�6؂Q;�X�35J�)e֐�hS�3-(ʴ�+))���n���iʒR��̋%ŏwi7������w��1˲�y�b�Y�n\�����C	�T�RU���rM6�M�zB�*y�!�[;�W�t��ɘ�C0�ޘ�Y��)�sn�D���2Gmn�0P.�DK�0h&Ö)`R+���n6萗�uk��mE�]�i�����zh�Ĳ�,���_gg����aR�o�2X;���k{��j��7���w��I=�x��v�-Ņj�������WB|[;�u��XF�p=��l�Zj�,�Q���ji�W�;���e'z�K�zu�"lT�Y�"SYчe�7�������f��mY*P����j۪��p�Gt_���e�ZWf�It�Ә:��(��-TJf��N��Ρ��u��&b-^KF�:[i�'Y,�V���C����e�آ՘��Y�Bq�}�qwuή���H;�&7��b�����AL�#��#��.�걝��V�����"�)4b8J������Ԇ�lRf�����RJ+�igE^����Wu��δ;uj%&�Nܴ���iu���I�whV��]��/6�3�����!��26S:���s-sp�Qщ�L���Z",9ݑ�K����M���s]�F.�b�"Y;����mc;'�vR�]�j]�3����r|(�a+;�ֵ�D��0�C��ޥ��9}��N�x�v�������
PS�?h��T ����Ū���/������p*8']�C�Č��r�ͻ���p�*Wi�x�&�|�xf��[�aJ+�Tu�Zq����b��R+жl�3`�?�n,����]�~�%����Z����x�G�-�Z�Ć�=z���]3Z�5dBd(^ryK�a�Z��)���7��ll�ե��uʇ���T��$1,��[.G9*s���]1R����;+����X�H%۬�VV �@�֬��`�73���u]s��[U��w���� w2�W:g�WD��r@�s��E�g���ݦ�/2<��Ը�#��z�WZ��J.<������׃�Q���Y�֦����s�V��K5+)�͚i��ar]��ʏ�Ĵ�Ǌۛ23Q]&_uڀm���"Ҳ�*� ;#�M�@\ຳg\�Ȏ'([;�v
j h���_8[5o�������%s&X�8��բȷ�BXE���w&��x�%�b6�j��՝�	�V41��Y2�W#cH7XTr��ft�� �E�l�:]d���LT�M���S�70�Ғ�z>�y4tR���9��-��ҋ�j�w#�FWB�;�tv�m84���uƓKE^"����,6�d�h!�"X-��ɐEeO�$tlW%��3R��WW`!��תU��A�ٗ��"RXr�D������`�������N=�K�Ñ�\��6�]:�f�Ju]� �λ�uK*�'Jd���n�m5nOj�u:Ci�` f�-ˆ����:^f�k�.+ר񫵶�PK�,�Ƥ���o�i�gT̐A�\p�f������e�ޥ�u���������j��=��~���B�kLy�D/�����V��Xic�ަ���/6��2'�(� ��c�4�ua��V�P���iF��ɲ�;�7�����$M��3���5�0��7Ok�R'L��,���X�g*m�ю��;�)��X�����`��,�ƕu�R�r�/TF�x���̼��λ0�]V�h�y�M�λ��[q~:�lO���1�wr�{Rd�¸�FS4� ��9һr,)+H�5� Ä��(���_�U�_�<c�/nRK#�U7p:W���NN+G���ix�9�u=dt|ܶ�m��SEd�����R���̠_ƬK���};^��b�]�ř-r1p7m;iAsU�;&���rP�WAR���!�w1$7�>1�J�ˮ���r�"G��d����]%a����V���腚��mN��ZZ����z�����X��Rrۭ�.^6k3�D�lnwY�L��d��+R
;1��5DVg|&�_e����B���ټ���G��\ ]��쁅V����q)�����ec�ˍ4��r�pfZa�Jܕ&�_�orP���g_'/2��r��p�O��u��Q.� ���̮����Y�ei�ٓM���p����X�RZdZ܁Sѱo\5z����`U���>oYbr�V݈yL4�;d�3�
��� d��X�3B��.�p+�[ю�kD���4����^�x l�74�-��,�-m�=7C��)ve=�Գr�g4�h�H?��y��s(��C-�0�!:�"_<y0_"�,>�C*���'�qqڲ�XQp���ɸC��x�T��'^d��8��qtχL����a7$�8G��"�mP��P�7n�5q6z[m��,WɆZ�\1�r-�3�wzݹ�m:T���q�ө\)D�E4��AORX�mܮ3)3��2�M��WN�z�ո��e�4�wkeζ�6��AE#���c�9 �sն�8	q��k��іn�P�_5F��zFsK��c��γ�_9�ܽI�	r�
9/�Zy�(P�]6��m�Ĩ��f�	�����V��N�m�(M��t�l������@Yݎ��t��v��ٗ/x�k��S.|2ZgS����-E�D�v�1R�-:x�uL�����_B��Z����A�Kp�89���EƱ��.,�];�e���D�vM��H���ړ"�7n��Vo����܃��'NfZ�E������*uZtv9�pQ r�:{3��ޓ[��	ٷ�@����.Z�fu�6�k:�ݸWAORەؾx*�M�(槢��p����Ĺ����ivv�x�im͔�W�z�A�$�6�Y���rP!�o�gN5�{��v����pm*J��ESn��+2�1����޳±��ﾒXݬ��\f^u�v�f)o�y\5p>�dP'���j��m��=�dz����k�͕��'�k���Cp�����ܫz���+.j�*�;�4�'�xhO2:L_�����3��������1d�ǽ�t��~���zl���K������7h3���K!�n��α�S{N�#����%�U��E��.�˸,�_>��4��km��ڔc��Q\4:��<�VP��r%��o�m:�wЌ�6&6J9X����J�>ĭ)����T���֦��0_u>�T����Ɣ���hNe��v:��g&�)�Ž)e��tSh�N�IM�EmCX�]�S�˲M��*D��֦	T!�7{�t�[\�i�[�P�R��X:�f-Ǭ;��nJ��.B�U�Bm�{�.� �ԗ4�b�1��;r���ܦ�x��r)�ʹ%
ǵRꛒ�����yj\	���F�sbu�9(OU�׷vN�ja��f�i�D,j@I^k1�U���� .�yK�d�W�s���;x�Y8\�����eb�WAU��Zb<9��sp噐�ۡ�V���Ǌ��;�� �69 !��_b|��2�O��{w��]w��+{�����xFv�n�r�J%��8Ru��,ɚ�+;4��Nb�����6��������Uq9a�$�h�s	BT�ɒ�)�{�)GR�/����+u�5���8$7N���=�q�R��T6�ԡIgV;��Y��9�n3�4[�n�ݺ��j!gHse�3��y�El���������T�m�{£Q!��۬�g��uq�ϚV��Y���5�x�:i�'��r"�z� �kw5�qp�L=�2%A`�6����8z٘R<�ŵv�"��{�����l��0��Ό�J�N{�R�5uۏl7�)��B>;W-�ճ«p�x�j��8X�dy؋\�`����:��<�k������0�C�ϻs�4m��'(�웙}��R����#���\�Z���'���M��l<�&5ƻ*;�e4�>=�R��ڹ�:��ޔ�oH�a�K�\��i.���/.��u�7�-9�1�@��ʡ��v^d<�4���L�mZ\ޙ���mv��L��'��zs{B��҇`���Q:���+2����Ow��\�^���/3w�x�{���J�.�}
u��\�3�+��Ki�����:75�H�J�t�;5�,��F��}�`��2��^�ݎ�G2��z�D4�(��˯{�$m�d2�n�WPy�^��엕�G5��'=����\��R�i�j:�-�|�x��U�����=m]��f+"v%�8sn��[�3�y�:^4\}��%l�p_c�en��Ϧ�\�����&9]b�3
"U)��mP�ƦQɏ����A{�)�͚�\�x{]��k�{U�jIQ:�fw�%=YhKb\ї��������E����H�j�c$8.�]���O	:}�g!G��rIT�X��|�	"�R�LԕA��
�.p��MrQ�옲�p��@���N���1ʳZ�Na�o^p^��;���n�"�\ �ssPw��>�Q8Sz�͗���MX�v��H�HoC[�D�I���d�ٝ4ܼ�-e���5��u:!L��U����g1���%���kLFV��D�Y+���g�{kK� '��D���O/���qg]ҍ^�1�3ka��SɎaH��Y���6Qjf��V���8��6\*�(���.1E2�}��=ޏub"��o!��E��Tt)��v��Mm�����];U^�L�
�[�{2���U 6�؎��Ώ>yWڸX�)E�[lH�S�$T�338顙�tT�P�xg	�ŭ��'�!�$���W����e����i�-����$]�&�	Y���ݢj�&삡KZ툝�ŋ����B�����"���T���;����+U��Ȕ����g��2�Sj�$yG�\���&�@��Z� �u]%�85��Rc��顧��1P��U2˦�6p�@�7�$]*G]��j�9���ϕ�.��
���i����x4)Σ[w9�͋V)XX5s��L��{�&�O��٥V��Ig2q�;�]�
f�R;#����J��'v=X����
��\"K�.��{�3�o:7�b�/����c��ܼX�/��gn��Ol�۠R�x�6��8�`,0�n�s��$�wk�F��ۘ/^�'{�}��I*jNe��Y��$8��ˤ��w2m�6Y�Ibl^�-��QtՎ�#e%�Ah�"k���F�nM[�p�Sjr7+B�������;J ��Q6�ɴa�\����M��m�hc3�V�͔0U�{�ϑ�Av]u��պ7EK��P�yH�Bw�������A���vom�8�W)��kC��<OD��hS�٩����S<�6�v�si�%��%�D1�/�|�f�uf=���D�2a�U��%�	)S]�zV��\R&�g6^X;A�wjT��b�T|M���*X��Xz�8�Tʻ톒 Zk&m�7�Nɽ*���	;���� T��$l�-�[wk5k�Dz&��n�v�k�'��K��/Xu�-o��k\<�3����5�kiG��"�k��{(R��%@�K�Yǽ��=��(L;��_mk�}��[ػgƵ���)C,"'t�1����_GA㷿w��]���+Om
"]���X�P�޾Ebwl��:_.@+�"�C(��\-&�Iv����b����y|e�z�
ÙӐ��w��t����5���}���=XSA�[�s����];D}�oH�7.��E�$\bmu�l���Gm�wq0ݡ]E+��0�_�ä��/q��WaوY[��榩-e�[�����K����;Lnm�K(=w�n����)te�./�{ݩ��k�,�m������Ё�j��P��S��ݼOuGi��ѷ����JK��}+-Q�vuN�HWq��Xx)W%����+���ںa���m"��n�((#Q�����W��}�Q�FT�r�6���d��bZ���>x�Zμt��ж����3G`/�+5i��Cd������b\B�iȍ�_G�śH��C�VXo�`z��Y�i��~������x:�,n���ڧ׫�V�'J��}�WTl����Q�bj�&J�o �r�IA��7��?m��i�<D2�qY�9�q>�։Sd�Ŕ᱓f�'kv(�d�x \��	l�W}\N�e(����'(h��������	�3U�,�	
B�o�aw�)}��z���K��H������;Z�u�,�H����@e�C�Ҟ����suhj,��X%�s-ֈ�q��-,L���b>Z��)j�ú��{@�l�*�dI�v�ùbL���]̕��˪ֵH%�8K���[��#W��l;,�77p����`���G1.�s	���BL�e���b�,a4��ɻ^hv^u�{�n�>��n�Bv�kWY���t�Hp��onp�/�Xe�mP�4��V�H�:����ڙu��v���;wE��dp�s��h�tu/�I1�z�1�7F���"�;��0\�����u������V���V��Ew�D:�:�b[��h��n2�J�&�Ã9��)o:��MJ�T�(��4,�X�����Φ�֐�®��8P�nG�<0�n�Z��20V$L���5anƻ����r��u�P��/M�g�9 ܓ�E���JIӫ�q��#�4"���v��<Ɗ�8 ֢��`�<��U�3�K(��1>73!�(��{z�p������sWk��q7;A,5��<�>�-n����
�1*� �틽�̑�x1f�:�h Ӛ;S�,'OQ1ܥ{��z/�:S�/�Ǹ��yC*�Ӎc�/�v���o6eU�v_sl��U9�T�a'*mM�1�+�0ܶe��,���ⱆ���I�.�7�"QX{�[���r�L
�2X���(�ũW�:'��R�ғr��aFM��g9�(K����s�鬷�O2��mb�as�܁�Wm��.�����O���9�[��TQ�2��v��7E��R�b]���`33�S׬���K ���#o��]s&G�Gf�G�������Ũ�DS�0��
O�6�ٜN�V�G$0��p�{\.K�;y�uc�����{��Ttf��4���Nu�r�+�����Q�{äu�pwBl�!�qMˊG6�N��O�\�eE�I|��b��H6\�7�{l�)Z�d��8t�I���I%�$�$�#�I$�I$�I$�H�2I$�I���8$�η���u��$�'$�I�k�f�&C?�������_�m���ӎG>�������y:9��o,.ܮ�$ζ�9�^$��ܭ��%՞�&��|d��.�E|>�i� �L�E��*9.�:�#ď"��;�w�Hb$O\��T����\b)���EՏ�C�>��L�DY#����!����9܏�����y�=Ix�6��(�ȒAS`�@�cN���� P-�Qc�D���Ms_�$��P�l���PA����   Q(1P)$*&Y�#_��.a$�L$��nA	00��*� �I'��yu������0�F����� ��_����>6�������=�}�g�6��ߏ;�0�6�����>�����������o�w������ߝ��cgR�%�!�F�b5�oe��y�&VV�-,1��Y�V�d�~��oY�A\]��̧R�i��8&�7ӌʍ]ky[�Y7U!��K�}����W�o	z�!�`p���CfIu�'���nkI�f���ǷY�R� �)wB��w`��K���a�>*�т�ԧf��]�1��s|��ɶ;��=�G]��zW}ԝ�e��b�]D�C�@L�|I��n�K�>�m���Z���k��d#.o5�˰��jzzܲ6,V0p����tN�N�6D�I�� 7���W].��@����*�;b6y����G,�k�8WNkso\\�Ж:�W���μI�e>!CgHp�[�YX�w���f`	��ξ�r"�)��R8��u`��J�U����2�j�&e7d���S.��eK;�n�i����΅�������m�[FԬ����O#��wH1d[��
�^����<�Ysxoa������a�r1�k}9�ά�J��b����Q"�#����Dآ�-��[<kD�,����^uY4����c�.�<E<���sdc�F��ۺ�	P��w:�*þ`�c�j4NMgAB�K���u��'���ۈ�ˌv \�݆��6'N93�o*�&�=с�:�
��Vb�%J����~ǷǃǏ<x���׌��Ǐ=<x��<t��Ǐ�Ǐ<x�����Ǐ<x<x�x���ּ���7��z�o����>a.
�S���Ί���t���n���{(ЃH�G�uᵬ�N�� B����6�>Ʌ$����>��z���n����R,<�b�TT	R�G���S�}��z��e9�2/�۩v^k��7e�O�X�;v�˙�@>ֻk.���*dw�p��{�m�������ug&��E�Zu._6Ġv��T�A��*�|�o4j�.(�y�(���+��u�E�v<7�̲,<���'�Oy��8a}�O/�4ݫ��5t!�Ʒ��w6�jq�[��ږ�ۮ�VѮ��b���BȠ���K����Rͻ�5B3:-k�������+Ot�k �!jb|)s{�%��of�zn�ue�)Ke!ۇm�w�]���&����O�7�c��5B�#{X��7ͼ���:/�2�cᛦ�C��38�����H�o��H�JB����y��	nL�����Z��sU*�W��L����fs,݃F����C���n��N��s:3s��u<th��Оh���<��D.���P3�G�!0i�Hen���D�D�+�*�̽��h�̒d��־�+�e�g@�v`�E���z#�Y���Ɍ��|Zg{V^Ј:�6����ҩmP�-�E�l����fɶ��/�oiU��
��m����r�D�x����|�_/������>�Ǐ<v��x��Ƿ��<x��ǎ�:x���O<x���Ǐ�Ǐ<y���>�O�ˈ�اIkn�Y�Z�i���h��N7�v�mm��;F9,\:�U��0��}�t��fG\��
�w6��+���?���&���}X+������l�8zh�W��+� yo+�lɻ��>_\N�=��@����U['$wl ��d��[�S�	�"���������ݹ��o�n��m=�Y6}u����dU����p�䁗O.ͧzI�*T1�}��K��[ۭ^r[\�q�ۖ��AF2���.�mZ�FK�wav��%�%��Xr���*�&��_c�%�)d�5g�$l�Զ�����oZ*�U�b���h��\D&�٥�;�xM��B�y�Ћt�QcPv/d�ocW��td;Lt}��]��V�.M[@�h�W�F��5%$�݆�]��el��\h�f	� L�(��O 4�e�3�H�aVp������Ӳx��:�[{�(�C�C��H`�uڑ�Z]��μ|��|�[y0��kld�W\��ƽC5Hi�(a�uj!ta����&��=��Md�Ef������W��6��~D�j��`� J^Y�I��33qM�}�`�����!Lc�aցJ�M����.�˂h�p���3�:���Pi�i
����>n 
�2仝����gv]k2�^N�^
t�Kۼ�)jG��w��˦�㵻��3)A�}�?���>��׏<q�Ǐ=<x�<x��Ǐ3Ǐ<v��Ǐ<x���ǎ<x���<x���Ǐ���s������[nK���1�Y,�7�/����w�ňE���_Av�W�dhV��>߸�ԩ������P��D�nj�	���Ό3NXߕ��HkJ�0F�����ť�m������n��iu¦%i�b���ە|�_��$"6�0:�S��%|�	�H�Hs:*�w���G-T��}9@��-�]�;cT�#�qyc���\1\�����o����0M�s{d�R;q__'`�哶\X����X	NŔ�b�x�X8����oWj�����:���7�¥0�%-�pr���ƺ߻@��	ܠd��Y�`o��m�cR��Շ��!*Jr�/��ՁL��S彖z_t$�WMQ�cg%������r�IɃ��ք�̉����y4iš�gi����*hmKS�R��cx���[Z���IY�v�a��s��RZsy�Q;݇ ��4�iЧ}��֩ ݲ�ꮦ��d����˟�<�v6�˘"��o����T�-�;-fg5�h��U_��a��qqb���:��f�Q�o��yϨ NMS+
��V%�D�H�fe�X�8�Bo��nb�N�톥`�\�gM&��;Ӣbԝ�j��j��][����g���{*��e9sm�.�-	p�K#�3�ÈA��os]��mp��.��B���W����/�#Y��TFҧ�B��O���}�/���^<x��Ƿ�;x���o<x���ǌ��N�<x��Ǐ�:x��ǟO����}>��������ǭ81ט�P���]�ߺMJ��NeՈ�Nr��#�͖(J��d�y������:���c�P��T���^�c7���n���񍼇�BŨ;
v��^�\ŀ.]-Z��a��XՋ�i;M*g^��X� F����mm�S7Enm�������9a���ZP�d�"�b�p�.Α�����bM�c���\�vG���m�
B��.��u�9��N�Ac/;�R$�}	!b�f]�����7֔����2���[N饏��fgǥ�q�p�O�xd��բt%H�K��l���
"Y=��:gY�"2\ne��(^���V8u �n��`���4$�Kԛ+wx��r��t��O)�c����M�%�}��}��y�c��\ˬ ��v���*���Ҷ�/{�
����:�8�Ŧ:3:�����툞e�Dv�$�Ν�Nm\N��W]Ff�3�:�;)Z�^r�uL$���תD�{w0���:�����m@w�_n����B15����Ծ��:,���,.`����\��.h�V����>Ic�S�4�8#ܦCM��n�j�K��wp���'wӻ�����LΓ`ݖɼ�^$��)\�p�V���o�$aΤ�Z�����Hiv�Ǉ��s9Nmd���ܨ�rV��]]1V�,flR/ ��VfN,��f4\���;P�Æ��k
,#�з���K.%�3+��V�hi�*q�'�I����������[x�i��w1��4��m�[S1��W%f��K���l�G ܣC6�,��i��H;wm�Z��uN��3h^+l)fX�ZF�y��}BP��͠\׹�"�V�����n�3��VU�}�4�{�HH�?6�=���y�i��;�v;ϑyz�I�W�~�"�q(��u]?��/diGh^��&��=�yr�A�'T�	cyغ,���!K2shj�ؘ���tYB�:�Qۅ�0;����_IlR@2�9�k>ͬ���t޶i�;[y������4�B�J��wCA��&��.�n��s�b$eoW@�����)T�K�;tV�2�2��CI��iE��P�:op��"�=���&�{/sS�"f-"i�v���9¨�ve��j#}巚Z(�(&��&��v/�����{��G��}�X�/v\މ֜I���+���5���(�3�?����u[Q�5->� �7�5��.���p��Z���Y��aձ�&��Y53lwt�D�*bˉ�:�*q�6�D�m�O"2�#:+B��muu�'�	�m_=��PȘq�����/4'�.�J�x�Z������������uA�f�����Q0W7NhB�%�lu��ҷ���7���©]���u��҉���7nEb�:IkGr�\��U�M��s��hT7\.�o���ak�1��c#��ފ�xem4���Tm�T]�P��F�z�HK����oY?16��Y��A�J���s����E_$�l���Bħ�"�^�/`q�LGy��n����X�O2f`������VeE7!��E��eb�x�r�읧t�d��H
Dz�l�a/U��B��@͑oT(���"�ܭ��b���$�=c2m>���W�����RaD�S��|�[��|�_i��i��ɻK���C�E|�
����	��YA��6K�]�	w3��qt����'J�t�V�^H�t����Wf���J-�⡙�L��f��>R��L�{�i�#����w�wQY����M����E�L�wi��v�8�]��(��X�j*��n\��d`�����|��7i�"��\�o�ᩝgV[��m�k��0�b� ��7�<78�׍,3a�r\gH��,
h�#�ZGh1kd���
ڇ�m�*Z���y��%�on!��{l�zyl�eۻ����g5�^9���B���r��c��/(7�[�P]:7������upnQ\��S�.�_0�M{k �����[�A��H���8⨕�뱝�ղ�1�7I����5�y�Q�I^�7�Ƀ)��ל)Ί�H���6E�Oj�CN���%���$M3�N��o�{(e�Ͷ-���u:l��%����p��:zخ�ȟR��:�A��Y�>�l�7m.e��u�<���j$,��ٛ4	o6�f�n�C>
�bɆ���Ƭ⨲�SK��ͽ��}n%V� 4�M��n�i��r�Fu(�e-���1�󰀨�)]n�Eҵ���{��*WJ���4%zM.�M-s�Z�W�h)�.����x䋨��^��7�$�6�L:��i�ɷ|�o�.���M�y,���;���&�E��m2�}6�׊\.Уs�ŷ����ڙ�h�4R���$�r=��x@���כŜ�kn�T��J��v��Ц^��F�I�[��,l�cі��4�4u��:���=���^Mѡ�p*�N�jk�Yѻ����gGe��NB������i�k�p�����YxԩqsG
9�x�9��n؊�qN��O����x1W�P�z3���G^��Ui���*w	ț����8�5���wI��U���{Z5e
���T��r��b�J�3��
�[��^���ZeoA�B�B�d�\��f8h�Я�qf��X���Z�^��0�(��L��P�}����CEA�Vm�O�+�����9��4 ����Vj��7��,a��m^�Q��A�ٓkYZ*�EQX��x��b��R�D]�D�6w�Q���$�{-���6r�(ݚNH�B��yU��ګI�uǻMu+��뮷s�t�t䴺�I\�Yv�1ΫhRn�R��}���m�y�\m�i6�w;�;���k8�A�1B�)�3Lu�V=sZ;2�F� �g&�uV�{Ɠ	���d�1�{j�X��՘�[���$z,j̾���ʕ�.K5�eN���n�9�f�G��۔�rm�B�mC�T�.-�iU����֗y|���Ɲ��m�F��_U�ڱ&ῑ�P[L_�L�ք�}�r�0��6+N�7�2>�Uj�/2b_s7�b�aC6����W25���E��ݶz3�)k��좂��jjT�����,YkJ=Ł��Ɲ�p���-s#d����w׶!Qi9aX���o�J��gl�����L�Yu:s���|�j��U��ܸ�b�YyWN0{Ol��W*h�D���|�z��%��{3����eH�-���ǵ��S��g;ں���"�1�*v�b��V���3�,ZL��ms��-F��v��H��,r��I��q3\�Z�����Cw�Nc��2U�ҹwwȢ�m�l�r*��t�<�]�5��΁����q�o����Sٜ`6[|��[�fjK^��Fr�}���A�n��wD��$�8�R(R��JC��O��O5vN�a����2�.��
i��ۊ�wq��T)��ؖ�}cb���zF�������w��oF�L.�pe�{O-83�u.��7c��ƨK�@�S�)1N���<X�`��W�Gf��"��� mM'\X-�ZǄ���I�V��Y��]m4VV�Ѧ�(�%�v�3Q<yy��2��[��U�Hl�&P���L�YϘ��e�X��]fVf������s����g �;۴���a��u���6�:Darٓ'QX�`�zcVX�æ�D#��Q��{	9[׍�]o���
.H;�bc|j)���.�W+��Q�e̶�(�{AZ��m����5��6E�<�b���\;3���]����}m�X%g��Q����4'.��Ð��c��GΑO�ljN�� �Ko.K"��ߐ� �[�r���R�	���d��j4�ƞރZr�&N�qH��j��ˬ3e�D$��z�1�5K�e��eu�,�_<��T�����T-l�)���n�6�]czF�ofL�Im�wтe��&�o��K��
�d2���V����&=(��Wו`�u���ĩQ�5�vc8F�}|����̀�{O�oMMԴ���1�{��TW]��"�̈r���:fSZ�7NJf�ы{+*�M.e�����r�N�o�:�v��R��q����t���]V��f��0���a䶆c�]�F�܈�h���4��.&7 pLW7f*Ƕ��h|������D�=��������u�V��z�倸�?H�/%/��w��v�����r�w�����~���p}[�~o��}��L�O7�v�;�޼�_���A��P��	��2d3��I�b����Q�_�h�3���]E��%�;U��:�~W*��8��Q�]��-{��}�6�I��Ȅ�9����nY]�s��nRO�|k��Z���͂Jg�X{;홷q��ը�T8Y�8�ef=�<렏f�j��BKΌ;�q�5Sw"}y�1Q�B�ςI��Zv�]�f�٬|�&b���N�wbH�q8E 12r�^�܃2�hi9���73##�w�4(����'x�%������wi��M�;X,M��LE�Аd�$B�V�lVM���9zͫ��뫉�]u�wR����t���ܵ*�q�·:���������4�:n;���m���X�,�v,�,k�-ܺ�)t�}]�;�	��r�Ҿ2�m�y�'u8�#o)�j���ܼ{�d�t��,c��Ofnib�Ve�	�0���v�K�6�-���E���`w-� ��<�_gx����g��s���N��Z�Z��j� o+�ז.ћ�7�١�Mغ�R�a�H���Sy͠�
e��P�Y�6 :�J4.�w]s �S���9�E0���cӯ�,��5[2[y�����.���n0�����bNP]����;����	tՉ��SDBD魝��F�9ǲ�]%g�]wW�Y�9��Wk�4Ȯ:уg�f&��k�G�ԕ��Yݬ�JR�$�N��*N�}[��h�i8��4"��MHdn?� ɆH%�$$�a��k�JPE)	p�J,�"I��!�BP0BY�����I)��m�a� �O�	L�D�����TEP}kLQMDP���w�\{��Tp�,�F��jիL�Z�(M8�Ǐod�_i
>�PAQUr(#�-J*(�r�Y�"�P�w'4�̨;���{���ڪQ���$QT�ʾDMC#��EȪ��2E����KN�E�ۏooo����
nd��9s���HFQr�Dp��2I�.S�!$�r*T��y�7�����r�����R�G+�Qr���TQr���
����E*��WL�ȸE�9\�"B�Թr�1�
���dGp�+�� ꔢTvS"�@�*9�Q˨`��p�V�*�0�**
��&$�j�Q�r��D	)G9D �)�*Q��"��Õl#�A�Tft�Ȩ��(x�W	͔js�ʪ*�$*$�e$ҹ&TR��s�N\�Y�Ȯ�"�T(e\*#:�IUl��
����*�,�s�,=J9T��)���J	./v���(#2���bS��U��d��������[R�i����Q��A�mu6՛�ŕ�	Cf(�l*�]l��Ò]}�۴��-4aD���\O��H�����J��v� s'�U{qot[:�S��v��ʱ��6mE��&���g =�`;���dl��n�� Q��W��nb��y�����ߗ����v�H���v#H��tr1�I'��,��j��֞1U;Gז�����1�ǫG��͂M�x<E�؎|��⼝�n׈ֽS��5��_f��}�\�gY��װ����i��1�Ϲ��	m�������Of��}��@��0=^��&���������mBp�%������5g�������1z�)����S4+��-V
�a[�{�N��J^��&�v������ߏͺ�c�+
goR��|{�.0�7;xyV _����d�����ӓs��9C�uD�jF6ge�z�"^�.Q��o|o�WS���z]^��]�;��g#�����b�9��זMK5��iw,�޸e��Y�`�ݬz4!��נ�OG�z���]�{b��_tᗦ��:�4)�x�t�^����}�=5����.�ۭRc�����p,Z(�Ǡ�X!Δ�X�gZӪ��Or\�ea���v�u�%L�wR�bXys���X����:��zY��iey�܆|��A���tn�k��֛7�����{}�VL��##=P���>��yxOA:d��YV��K<��@g����p�7�����
c[-�Q#��p�֩\�:��Ev�[lg98T|�V��W˽W����Q~`N[��^�G-{q%0TR����O����ȼҿ*�mv��+���7��z�o,�P1b�0ͻ�v�%��v3���T�@����3xz�of�2e���/q]w��M�^󸤲�>53:O4�*pW�ԫc��{*����c}^f�����U��m��ބ�U��2Lq�ɭLc�L��� ��&(�W�r�r���7��ɔ�g���W<�������x;ә�8S0�[k�tz�O��G����[�ޥo���d�����ѡGvGut��z����&יC�{a馶!q>bn���_7����[��i��H��l��U�|����Q�%��t������EN<��7w��O��+�$'A�Ǝ���v�VY���!�h;�&�<\o��R/���t�0;�����:���$KY�R�Nى��~��g�J�L��O��/'����%/@�2%��8[F���U�x\�3�Vk�yx�`y�ޞ�^�Wa�F���A=�������������:��l�Vx<�#u�C��ɾ]��������]G�Ռc'H��rxtv\N����/<�F���X#rίq7�s�а�_	��o���7���q����.r����*`���+����(����Ub�ܼfW{ޕ�s��N[̂�tڝ@�U0g��ue��A��c��b$��|hG`wF���zp�ǘ���`��U)=�1�6^�$�8��i�"��x�u��z�"';�Df�aj�?U�V1�������w���U��z��o��k^e������դίc���<�C�U��@�ɷQ�]V�҄u+�[6��\��O�����m�
��&`D���	�a��c�{�R�tPzgS�]���k1m��&�
����df�xJ�s��1T~a�΍z3�Y��6U����\ow����֗8�,��Y@�������5m֩��K��Us�٣R�O�#����[W�Ǹc�q�i�,:�m���^0cs�qe]ʴ�l#oҎg�s���w8g�uƵ摯����L��s�Q��vUnʀC��X��ǹ�
t�W6������\�\�z�����Ʃ��n��u�r.�y�_��|�e׿,[[����� �ׁ���$�%�zA;�k(Am%��8��L��O��@ ��"�c����*�����^�{�����ZS���~�C�^cσ�l�-��o.��˜�%���k8��D{��x��)��'�A�x ��k����X��l�ǌ[�`4V�qjL��;�����{�|߮W�\ݥ�E���Rv�0U�3��������>�ݛ%�F��[@7i���`��6�l�vA�6x�Ɠ-�X��n��22F�Ӳ/�����ih�������
�j�
N�Pg772�Ñq�7c%�t�{|�-�۶�Ѣx�����k6�}}P�.1�vGZt�AӖ3����`´�>[D��R\;N��n<:�F�b�&i�ˎܤ`���nm�Ԉ��#��jI����/�������)|Uu�7`B������o�����ӵ���l� (�Rs��W�g��Ð������f�uӦ|��Ϝ�#��;��n�$���E��WQ�Fo�^�(c��n���Vth+�:�3���s���v�N�Cݥ��^��t���W0��꒮�3�x�M�4� mL}]��go����X��$q�$i����b��5�	�9�<kZ���[q�շob��t���A�G�mT�A<�f%�����^>��1:Gi�G�Ký��y��oDi&}G����v�"Ͷf�tOsN�c��p0mA�>�DV��m���|	���$���{Ƶ�����]i�oչ����8�Eϣ��Z8V�k��U[�s����Zgo��	��s=t|u{���ת�k�f1�Ͻ��L��������M6{��K��<o_���{+<�{;&P��]E���8=���:������l�C�����ӿl�
��^X��t��^�~���9F4+��NY�8��Ѩ�pv�>����*���hw�c���}T��x�(Ŋ�2n,r��;9A�sT��'Vk<t�.�Q�[����5N�r����ڥ֛$Q�o:��0T��Q�{��M=��;�}��㢥�-�����{�b�=b�AX�xQ��J���:�g�m�X=��l}2�Nݓ��|ܾ��|�=���OF]2���(���79�,I�@|	�WSLR߅G�Z�����=���{�ۥ���ַ=�al�3������;��S���]����=�^w�v�)�"^e1�z���ymL�B\��ʽ.������TP�<�k�U��f���M8�*FW���r��#����ʺ���XWX��/O�������z�q������7���;��жWß���VV���nz[��G�E{��oo��+�]*�l��g�շ��x���Ui�)�k�H�{a�6"����O`1���oS�Fvx
7�O[w6]�a�r[g[�����}>�k"����"����7�?<��u�~�H��V����61�k��;�Q���r}k�I��ق@�%�rt�b��n�g��^˚{2�؊[@�Nɂ%�s��h�cq̐��1�7	�V+���mj鷡�ަ)���Ȗ����Yn�M��K�Z��pZ�x�>���-.��J�w��;G��}^�*�ΥF{@�rwI���5c4Gn��DU=���%��4�5ci�M3�q�.`q���{D&�	1�+wv0x]�U����P�&A<j�/g�t�u��"�M�4&KNOfў�z�0����7g���y�����7�l�	�ۧ�<tMbC�tl�v0Ȱ��ёY�j��Y��4t߃��m�,��:�0��3:}z��}t+�J`y+^�l�S���r��OzX�@������S�����,Q�p5^��V������zU_����܇]<�٬���<Y������,ۈ ��a��o�9N
^�O��xkVT7�1�Z���*�J��Ω���o�<F�ߪ�yA�?��%zn���Kr����^O��We%��n�{�hzf8c��:ۓh_̎�i���/e�w�������o��cמ�f{��f� �^�l��{d�����\�[{]�6�}w�*},���Xݗ	��d�}R��I�j�x�\`����r޻c)ծ�s���۬�q$:\���6�Y�8�Z����_)Ztz:���)m��6�������9ۗ)��A�c�������=��c\z��4(��7y]`f�U�����=TF�4������ͮ��<ǟ?.�}�&�^��eG:|�Z�"�$e�k,`����h��b��A�t
�O(ǯP4몥�����}�m�V���ru_�ތ����E�ҽ/�{p.�%��P��;�W҆n[6�5�E\v�M� �/��w5�7[�MY2Ltf�ؗ3M�!��0�N��;Ǣ��)�s��F֝�rO3������C�������l!�\���^���I}�oו�s�<����^�{6I7�6��d���y�=8v�γ˯�ŕ`xp��<�OY��]V���=���h32����N�xz_�L��||^
�W��M��~{���l�)Ȑ.���\ގ�
j�(��TvG�	w�d��,���:�3h����]�`�Y��9e�V����=��S�<������4q��Ѹ�r�l��#(wQ4{6�YuwYeqh�C\n6S-�x�=&�n2kuGvt��}�:�&�y�rbVJ�椯�7���zL���W��(r�^����m��h8��/J�+e�z�v�f��OL�|߯~����+�F��՜�e�D��mo��MǳD���U�2�5��o��U�z#�OI������S�����>Z���S~�|+j+5��T?,�)�6��v��r�±&���h�	���Ŷ����!W����k������Ӣ�.U�t�h�����y>E罍?`��}`c+Û�|�r*�X���|Y�bM�"e��4+�X�N�>;�8����ا��D+�����E���n�^��w��ݷzDN���ȑ��
�3�NdlǞ+�0��踛�ң�j���6�q�P��$Ћ���;4j;=Ǳ�ٵN�z��{���^�'ی��aY<	�&�#d6�7^�L�G�נ���\1{oY��wb�`M�>���F�Y��c]�2;+��/01�;�fnPP�Eq{��Խ�j�[�2w���y�۞w�=i��T�8��[�M�$c�zite����a�&��b:,�R��Y��r��ؗК��X+��vaҨ4�D����me䆣��5��7s{�M�G��������l�r	�rgN�e�m�s���{�x,����U�+��X�^��u�O�gT`>���#�������'�&{��T���w�R�^�pسX�XE�6;���|��=sƀ�'��ɟY�����;	pAf�ea�r�>�{�f��f�wOW��L���4k�}�3��W�Q�h ��=-u��{`16 ��g9�"4ϣ{���<;�D���S۾���pˑ�%5�X�_$�-�ݚ M0q���ݛ�&p�oQ��������z$�h!�n����}�_�d4�7ͣY�oG�a�6@��Vm��ʷ�I�ǯ<�����W�������@������@'��A������vX�݄�p�;5��6z��-Y>�pOH���$s���'���������/���ws�d�b�˗���XZ�,N�]f��í�������j�5��	n;�]�Kg;-%��v�u�1�_G��J�Y+J����Ri�eZ8�9K�8ֽ�Ù�cz��0g\:g}�G�]�7�a!��1dxU�A���t`wa�iԥ�F�b��ΆL�¡e�Mo	q'��
�GI�6����������s�k���R]�[��.�'�Vq�_)k��R
{�"J���7���GW�b�G��෮��4j�Ժ�<ar�աJ�v:5�96��'-C�����(�67]V��mquy�*/q 0�tǕ˒���P������dn�5�����W�!s��b-p}��KV��V)
�xUc�[�ku�8��Ԕ������/FKv����6f��� ��Բ��4���Տ��;	��\/�!�G�s�6i��t���R��O��W6�B��y�=(�fk=R�۾GQ��������vR�h���Q��xEt���j%���ݸu>���Z5�`�v��V:�l���^]ڽ��V�ٜ.��aq]��X�6ܺ�E�;/%e����i:St���vں�خ�/��b5n�h���-�czsw�Yu�$���0�F���V�-a���$�Ɲ"�/k�e��n����<i�|[ĥ��k��]鵁H��7��ތ�؞�,q��gɷ��f�"�m�.���m���W޸��OKs�X�^AZ�j�|��v�$������k���X���O>��'���"[j���(�lh�������byz��u����;���(��_�Z�]{S)�D�{V�TA��>��6_u܏.�i�{\��uЉ4���^坉��� �K�%W�' �:�0tĵe�w+3y�w���_}m1�
�<�D�;�&�n��3x�����>.�i���p�]G1�7i�ݧ��J�7E*y�aՐkr�iX�~�o��+5�N�uZ��������۽˒;|x%N���a4��\�͂�SW�U�j17�Q���,�3JV�Cv�qFM��v���y�ц.�!�WҠ$�1}��}u�u����2q@�n=��U���Aok��x�6��a����k���QǪ���F0p\B��FF���%�5N.�:-��1ku�~88�3|��G
�m�^�7���Goi�up^�^9���-C6j�WA���rRͭk�_s���K]�N����Y�9-��
*�o8������QXJ�\nHf+��Q���'�v�ҴVM�]̧Xӝ+�&�^�Չ��R�u���c�K�koJ�����nV�WY@��k���bw�.J�r�gM8{�l;7�]P�V�P滑�rq9�P�S�8�R�T���\�H�L���M2h���b8Tr�0�W3�M���\"�:��^�A �"/>��* �;x����ד�:���b�f�(��"�$�ô2rr�_�.UPB*��E��\�Eʊ�ě�T�����ە�^�[{I�Ky)��?\�RS14S4EE�4EDkV�n�)�7�ӷ�{���w	�.]V��&�,#A(���"�s�8z�U,%.Er��]��Xb�+
XB�W�>=������{�|�"�oj0�qj���r��!e�;��:�T@���ėwp�RP��/�prx�`��ӑ�Fy��V�������:Vi"�9UEH�|��9I�Kԉ\�,�Y��#�	r�^YULӝ�<�s�[�NR�QR�ź$,��3Net���e�Or���y8z��/8�ղ������c�㬉L3�I�UUDj~(T��[���[����!��	"���/*N&Ur�2�+�p�7L���D�"(�D��Q}w	҂5�#�L�$�B=[��z�}P/Ke�S!-g�9���VE:U!�@q2?~IB� 	�O��s�j��{�t0TzZ]��۶����ڋ�X�Ѷn��ݲX�n�o[u�	6fu�"�9��,������W�z?v���d������&����4�!�q�^��{��������ݻ<��@�P� �cڠdV�<��5���-�0�ܞ���g;�Y�p�4����YA
�%�<�{6�i ��p�܎j��쮾]/��LL�J<3���O�a�^��|�rfڗG�vm�vPej/h,�gT�jqR����p�j�:�)��V=[�P��Xt^b����	�];���%6�LDi��mʺ�h���iS��	f,l�)��k���a@�f=zޭ�[�	�2�D��2�[ ��f9�ʚF`X�Rl��i�T��p�����?��+�I����|j��:y���(���c�M���,�[Q�{[���r��xF����w=?D�I��NoT�eA#I��F�� پ��Z*=f(�sR3Ya�k4*�^�|M��z��̟���a����+P]�9X�"�U�9�����E��7ǫ&dF��枬>{A�k�G���ژ��{�I}T�I�M����N'+C\�_]-�5���%�s�L��?�p��-���~���^�b�~�21��V��E����+.�2�oj���#���6��sһ��'|��TZ��~�Τ��6A��v���;ݛ�`���n�#Qg������dB���W�&����:d�S��qdt1��n��#SveJ���Si)W�8��Yκ>�gEh�ط;���r�&xC��:H��\���*�x����'�(�cЅܣG�ƺ�W:�X��n����.��,՛���|���0z�%{��n�N�V��P?J,T���!���}S�tW<��o��F�M�uP�aԦ��c��b�b�~yD�Ƞ�1U��'������Z7k�q�
C��]��s��2��Y����:�1\��-E����>7"��Tb\������u�)����� ,s�vF�V;�?��t��8���Ũq�w��S|%K%S�r���w�U!������4"O��/n9�'X'�m�{c�*��4�G�C� �du�B[���z��C�/݄eqB�qt��������?yd��������T؈߄���5|\�n��kS~�[2W2]�sg7�[:~iw�\]�Iݮ�X\��v�,� ��V�{\��Cqzz(m.B|n;'�,�,J��r�Om�Qp��3` �^��rqms��<��֍m�d'h1~�ş���,{&)/C^%^�U�^���\:��w�'�o��i��`�^ ���D��u9���!O+j8�![���N�ޭc;m�z0�y��n�W��ߪ���
�zJ��������Ɇ�N7z#�U^��:��jJ7M��Q�l-��b��kc#�w=�CVr��ܝ�a�R��w;�Y�E(|�Z<~I��#��t�Y��{�
�ǖ��koW��v��qN�(�-��L��1��J��RS������D!��r1U+�+ض���s�z$��9�V�7��v�oR�"�sjs�n�_����d�7;jN�$h'1e��w�xa3�>��4�O��Na���!�٘iM��`�Mˎ;s<�^v�.aSz�W�M�Y�09�-瑴Ms�w�~r����"jּr��O�g����N��악���'��h��%s�,j�^[ܔ��m2>)"k�صW�������鍚Q`t��lY�hCg:Ps��YB̓qŒ��6�y�ں�^�>�{��<k�����Yȫ�:��B�|�����@uH���4-XQ+u��\�
�Ix!T���g鵌4��=7�^�<s�7^����!�>.(����?m�,9�aJ��m�ܡ�pKc8Q]��&b�ܢ���A�����V
2�w�\=h����߯*Y�u{��a�,+
��������WN�v8��H���g�1d�5Eߜ�6$����������2(V*�޾�6�v�;��}[G>WX����YV[���.nDx��Bz�o�\ł�J�ay����0P�Y6==���o�z���hW�ˌm���H��sY�afO����ު�n�$�kr�|/2f���{�bn=4a
T̼��,^��䴨d���@z��?��g��v��yoVtCג��O :]�l��m�lgxLzBe�T��3��ǡof��4���[��T^����ƛ�H<�c�Fx��E��k�"�m�P���3�2��mqG�{��@T�P~o�h��Obj1���Kcw���Z��`�:��zm�1
[�x^dӶ��s>��(tS<{DƓ��5q�tcj�ډ~`#��M��BeBҡI�5�57rz]�fg���1��ت� OԬ��x���C�%��#| ���G7:c����Ȭ���\͘��,�B�F�c�m�'�o��[Rt��z��"|����}�fc�Ҹ��mf�����;f{��x�E�7E1H�g�w���~�*ե��$x���#�GNPl���]���Y��ub<#�et<�Ȥ酁ʥX�ʱu;qs.X`���-�,�0)�P�����防��a�7`�U�F������z_�E�洠���K�5'��.zwn���;5�&�����L���z�0�Bmj���P�g���-C�NP�%Q��j;��J����͌�����'�G���Z�݇)���vn��L{ �b�B��=�7U�d��ovYn9t+�6\5�u��R(+��-�V%`��s���po��yW��GҥP�'��杳z��-�;L�
�qg'5P�*Vs�ʠљ�ہ�s����Kx�`-�áy��O���ga���4ڬOQk`�J��q�Z�7kN�k�,��9~�/w{VE�s�>���vB��W���y"u|o�FN�{����xjEC:�ER����k콠8ϧ�8��P��'�<����y��hz2S���JW�4�:�fwzu��S�ݐ��fI~�Ǥ���qh��(w������>��ğ�x��{-u?YM���iߥ��f
���ŗ	1���A�l�m.x9�q�v�_Cz�ױҳ�n��=1(�xv�g����B�O��?K�=�u`$Ww0��m�o�gX�B�K�}΄2CF����
��$�\���e�^m�^Y�:h`( a4�22�ߪ���[�6� �3m��A�U����0��ዢkz4��\bYA���z���WH�x���X�^�^�W�V�+v+����it1Wd&��h�ai�7Acj �MV��{�q�x�f=[ռ�|w��7X4���C�;�O�"c�D&�W��5�!�ޢ��Bq��K$�3L�Q��qo��L��N�Ăx�Y<�_܉�ć�><��>}{U��ƞ���˗����	B�3�O��n$��h��~��-`V�����;uPjܪw@5�,!2�k�w�Z�0eN$�b�cr���=]|
-|�9}���QN�� ^0y��L�k�(�^4�z�ê{n��:ݳ�M��1N�Jcl��H�>ҹ۞�������e��?�i��6�_Q������?|�\3[O������}},�H�a�'��$�E'(t	o.l�g�ޜT�Pyƍ�;ӵ]a���O���=�����"m	��/g��߰�v�0����Qi�d�牣fON'���{�8�j.���#4D�@C�==1�A~?��ޔ�yʵ��c�6�L�y�-�a�iSO Y�y�*��ćO��$XׄCc���UY�y�t�����|\��&iN��[r=V��
~c�ɷ���U,�Z�"wQ��<y�G�ʕ
��}�����>s�����BՇR�è1�?b�t�Z�� wˬ/Ө4zs ��Vf͙y�V�ۥ�wXV�:�ŧ�鰽N�����Ga���%���;+�b���-�PL1��l�Q�$֞XsM����C�"e<J/����6A��^�ӧÙu�Pnys��hq�.�8˱n�{�\���/�.�]CF�w
�oE�׹�~��D�z-��&�*�������O0�������"�ػҡ�v��&.��n�	��1���	ք�s��Ѥ�ˈ�V_u��b�^�;��Y�SM��a�P����@��#x�ׄ)��nS����Ʒ���SpNn�g=�ׁ%�^B���sU����ǇRōv�R6��0n��"R?~�[�o%ok~�@D�C�#�'�Dõ5�'�<���l�w�������������a�$J��ĳ���D����A�PK$�3���6ʆ1e|�*I�c�d��~��3�RI6U�r��Ւ��D��v��X��'ְvOAd	bWN3��{k��r}q�͊�숭��cKU*����qhZ�\ua5��/��|�vz17c���R�M�j�����8�s�,��r�m�٣���65�Ĉ��Y��0����Y���})���2N_=����Z+����y�>�Άw�!��'c����1�� �H?�Ðʶ�6ޗi��*L���2S��u�U�,v��n��ר5H���@ߠ�����F���y#a�O�0�}YfdS�Ү��Z!w�Z��0�}�h8�]`c�η�F�=5�Aߙ�=.wb��B]0YnN%4��d6�q��R��;�)X�I�R�dâZ�d��a),h#�$'ٷ����im��sZ�!خ���mT@�IԼ�:$�6I��T�Z��S~WZD�M~����(,OB��W����@wm��:Ƶ|�n���J�H�j-U
BS[a�e�n��s^{ʞ�7r�S�g�V�L�5�MU�R�qAQ�yID[U*�iY)�:�y}z��Zc*ow�<�Y2D�*n̕�O����w��<�4�b�Wq�ݱm�~.\�)���`�{����s8/��O09��i�j�J�a�J粠���������4����d����Gk�:/��B<̆�5���f[^΢Ú��^�.��w�����9�ք��p�Nӧ&�,�j��.�����omו	��������$-T+���y�4���C��v=30���$��x|ז��V���)�i4����) ����7P��\�F�N��{���@���].��T: �xc[�}�W���H\�W1(鍮�
1��+^���^�o!�����B����6���b�.�y`�vf��л|��C�q��D�U�ѓM�\�&���A�+�<���׋)��M�Ww�UD}�?�5�5�L ���`��4#?��d�f���MhR!�X3\*��]��d�]��r��];��4���{gh�-��Đ�Bc�!>��;�?]�;���v�c��+s�܉�/��V��3��S����-�?|w�-�'H>W�	��io(xe{{��.��ʫ�v��A�Օ!�g�9�Oݹ�v�dNϷ�F�V�}O"�m\�Z�YD�E��i*�cqنiU�м���a�X������᪪��N�-�\�fܩW�ol��WC�7���Z.�V�]��7�#�4ovI�7���,a��Ć�hY�^�3%:��,���Li#I�(?E�{������]���4^���{��uWZ����"D��P��{Иg�������^���ۨ��3�v�{W�+,d�q���\��ak/P�f�" �`�ƅ�Iz ]���z����J��.�����Hi�r#eor1(k��p�����k?��xN�`�a�r0ǎ8��2�j;��e��CP��FY��6��̀l!4�a�[�v4X��(@��
=p���6��M�z�[+R�3�+$;qȟQ엌G��jM�`��{�s �a�pt[� ���@���$O/��d�.Ӆv0[1PS��$#����{�vy�Q����"�x��z����K�jx<h�_s�2�*hӵ��6m���v/��.���~���8�a�zN�/�Zӏ#��)�WX�c#�]�[�L&��B/P=����@X~�->	��~o`19��!�i�C�$@"G�b�7���k�j��V�g^jv��W��Y����2H��I�uE����CZsp�4�����(|.�=F�P�X�a?N�n�ʭ��'[g��N�O.�3���ޠ�����[�ࢇb8�p������J^	����8��]˹���jN�ĠC�莄��p��RuS�Xӛ�#u��n�{]��_9��m[뭉��I ��:R���,�;�����{��l{��g��:�6��ͼ0�^����%55x�C*Z�lm>Lǣ��͵.J����1����-S���Ł�������g�*����RX�V�J����,��,<�(�����GI��^�n�/V�l��Pd�-)��t�xz��[ռ�a�ݏ��d����j��|�^+�dJ��nB(:�G
����'8ĲN���+
�&���|`+���Ȫ�\<.6���\v&��P�OtB�㝛����,!	��E���-�� �D�65H�T4���nO4E>t���>C���zg~��򺤁_Q8m�Н����+�;$Î�2/�1*
���T2�2��u��9Q~�W�V�B�By�Ȅ�^���7��s�a��a7C����[�I��v\t�u(��A��/Z�H�Fi����a�Ϙ(֐!����^�zi�>G3�I*̇��K5���\�^>���ct=x��zO��ûk�Y���Q_
=�U�����Y��9^[�ą���6�[Q�V�{ғ��`������l�6 �vm�63���<?Od
����~��:���<��c�.���{��
�{��M,�;��35`0²��Ys�g=wd�ؠ�C�z���8%�f���d����Y�e�p����<� ���H9��M��S$w'�zĮ���-�� �eJN�i�:��;�al�I��@Nz(�Œ��nY���o�T̚Պ�Oyk�-�ׁm�
���A������M�ǆwNA{&p�n0� RA��/0�yx�7;�g��Q�գ41[x�7�4�w<�:Jە����|�X�BK�Xʌj�(ҵ3��J��vjU�I`�PMߦn�8P$ ,Y��i��8�x���ȱSua*��N�W�cU�Գw���b�OL�5�ӭ��|9��u-�}�6b�n|��sڮ�fh�fӱQ���n'PMع!���|�ͅ�݄Z��sT��Ӵ���m�7w�
�.�G�l/�[�z �4WV��Nt�p(�]�:���f
OuMߕ;�[�[{
���h�2�=�/R����C���s��4L���Y��21w�_9�[���2��W`�v'cAVN���[��Ք6�JR��A�";�x31���Ɲ�ˮ=�\����a�@V��s'T����%����9O❇.tغ���*�L��F�8CԚ;�d4�m��°�o�n0}k#��o&50���76��,^>v�.w}TV9>�I*i�+`�3n�[!N�;��Kޚ.К��ZnP��dNM�$,̧��Vʐj�{�m�Ns��tw���䴭��"h��o��3��2�[�� �XJ	���G�+�Z��~��lu��.��8�u��+5�Z�M�a�$H:���r4�^9s�ħQ>�<p�]I���v�V99�KJB�����l٩��D'P۾�tn�Qҟ�X���-* ���ir|L�%y�y �E]�pr�֗P��]�AP#Bn�ϭ*Y�*j��Z(��:��t��ܝ��js��X,VX��}�m-���a]�w�9�9aٔٮ7�i���bn�<$x�4D��V�ۢî����0��ja4�m5��:�щ�G6��j��ƴz��p"mK����s:��}۽|'�v,��{Dz��ċV�JI��'F��\[]T��)�׆;%�	Υa��9��� �F������Ϋ[St�c���6�:ouʆoKQ�����\��W�FНNW	q}��E��ۖ!v2��;-�cW�S���鱝����U����r�IZrp����f�3*��v�J�6F�R��&~�۔���֝
`�0�s�\fV�5; 2ͤ�%c�6�(j�1��� 4F�=E�M���wo&�l�/��ck`z������<�h_�o�+R#$�7��[�n�l�¼�lM���E'��P�f����T�V��c���b�#J][}�b��/�����b\Ln��L��s�-�|CApҾ�=�d��p�n$�J������#T���lT�J6%L�8�y�����W��}�qa������EQs����J�TT\��3(�DXi��=?Oof�;ޢގ���Pj�r����DUx��$"���EE�dE~"U���։�4�>=>=��w��2$z��-i.�s��
��"ʫ����A�z�EB�U9�ΕW)&����OootLE�����"�**(�U��W ����oZ�M�T1u���ù*%˽�P�"��O��֏h]c�>�x��r��P�	\����t������-l�P���EEQ��E�g�W"*�ʢ�P����g*�TRBL�V�z�x��&���Q!!E�Iǉ�S�c�U���u�+�DO-�˗di�
�"�B�Ѩ�)(��V��*����"�F�� �RyNl*�T4bTU	���¯8���|yS�Q ��XNfo�V&*���ͷ��q6ַ�m���4�1� �ˀ���` ��Tq[Q�S���Y��B�E�M��1��pxݕd�b�ɢӄ$Y�cF)*�|�s��v��K贳��^�$z��/c��~��?
��cYc�`���3������C�ۻ:ȝP£I��*�G����<�ňM�"6s�V˗��������0�ƧOc'��Q�S�9���6�w��-���;�#���,�xu�c`c%���(3��'y�"�w��:y��v�s�ӻ-�]����q+=�p��ͼ*�&>��`������0�f��,U�mn�ʖ��o]��E
��3��5��à�����ʸ�jz��I`���1���E�%�lE���X�E��W�ݨ�֞�(8�rb�VI^(�3��2���PK۾q��鸪�x��2{�n�T�����L(D܌V'"��� �X렜��,h��g��|`+�Qp�C�:���D�5^e,L�md$t��'eLJv��u���!s�D ���):ĤJ*���{�L�3�A��@�'�xUU
�6�t�\:�dc<	���,����f�7қ��!2Of"S��seU����b�6緃lJhR�N.�gv=4�������2'��R.���5{/�َQ��֭�K��vކ�lw���yy��)�}}ʥn�F/]�����X�B�F�5��Z������t�04���Z��Aܱ������|��G[����n=��&v�6���򮾂[j�C;+�GG4��;O��2�\���_�;�W��\����CU<�l�q�H�΂\h������w BF4�r�	�G?vwN�z�SJ��cEv�s��6�/z��q�N��Ô�"�<�4�o(6��W"x�XV_�����2��0?x��VҐٮ����8�`4�Q�\���W(��RX�GjHO�ێ���}&�v3�uy�]�0{`4��2O=uEs�7"��̜qvJ�­t��u�$�o�&�ti��n�%��q��*�:�1���B��������3���Bպ��:�cҵ�r^�GmF�L�lr͋���D1��E������wS�?�G����g���3,���X�J����D�l������Ro#Ӝ��A�UyX+��D�yCC����sƏ�/����x��x"�N٩ې��L(�����]����P�,�)�%�����,jj}滾	��ݞ�z�&�d��ب��ݖ��i��_	�1@A����f������-3��	�e+�]t�y��Q� �3$����{k݌i��C�v9o1r���4��m���a������[�i�oT���=3��gnsJV}+lXq<�ˊυ��
T�^m<�M�b����o0S�|�Q�/Y�F��l�����wYtK�����sk��[�v�&TZ�����5b\�\�� Ʉ P���z��lm^����h�}9���g���W�J=U�J�D�g����XЁ�����`� ʭe
<���d�M�ST[����0ў�+��[��P3�U����4�����\ڇ�/�߃z�}���Z��A�ж�	�%��۔/���[�8A�z��U�K�Y�O�/��Uj�zd���CخR�u�4�e�����l)�gEH����Ǡ5��c�	-�$��:��[��ɗ����xq-м6E�W�oL������#p�7E1H�a���

�?�~է��x橍
ʰ�ܻ����g�z����vQ��y.�r�\�k�.�n�`ӖQ���.���|���B'/8�� ����@���ZDp�n�0t��У�S��8����Z~k	Ab����Y���q��魥-�mma�v��Gy����Zc�kuLIyM��,V�,�&^D�?hf�/�V!�J�G�vF�q��^�<�}a���k��M6����B���KvQU�.���X K�<�T�/b�sJ��m��:Cp�C�wf������ƛn5�ر�	�f�t��Vijs���m�
m�ݢ�#���FFΜt|�孋��y5���h�k��Dp�Tˤ��{7�t�� n��:%m��!&�ȉ�˫�.4Vmd������W&v<5���\���3����s��m�x�o6{c{�x������J��)&�Lׯxb����1�GS�(�[���>;r���b�;3�����/+TTC$3C.��8ۗ�z]��u�s.���n�f��E��Ǥ�qh��+��)�mv"-�Ķ����֘�k�[�\x�u��Xt�O�T�x׽t��7^M��>���D'�R8�ky픶>J|FԿ��Ԯ�c�P�C"Y�!	��!�Za�z�ǳ�#73M{ݒX�N��Nm�g5B���߄g��
^��_�KL�eW��i(M"22��T�y�nL���N�n������m��w��Lڂ�!�Z�`Z�G(=7�=���z��C�S�{�h���R��Y롣'm7lp�8�r5��i"Se�2�&�Ji:��a����ޭ�[��+w���Z��J@P�]�h|܁��β~��/��Fi��(l��Pߪ�,c�������Q��`/"Jy�����w� -��A_����+����~~�N���NoڤS*H�kh�VL�\ҽޚ���l��\:���a��D,���_K0R;$É��$�����F��]���b�*Ky�8��"�)��s��ɰ�T�7d�Wꜛ��:��990$���b{r�d��R���>oo&J��{T�0�ys�&n��9���֫Alͣ��vmk:�Kwm;n4˛
M��̒�v��/$��s|݀R��߈'��P3YSФ����@mp���&	��G��+"|>��_������j�k"�5Ym�Fr"vE>�ff�.����c�L���@���?`a��Q��,���]���� t2�?��i�~�R�rƵ�l"�J1�A(�zO�}���|�"��D`�:��9~#'|~B3d�lB�ٸz�C�)ơ\�a�8�Llɬk΄���GS�W>�U,�C��Ͳ4�8�F��m���#*܍M�8`�>'�v�<�:����ȥΥ0�cYc��ϵ�{`;�G�6�Sۉ�؇�x�홝֛�#" �2�K���|g�������hGP�I87�Fi�-�[dЪ%��9Ǟ�u���0K/c�o�\���ɕ�qG��\e?!6?}}�(0�P�<�\��9W=��_��S�+�d�#���$3���~U�Z~�V�tZ�D�N�zq��������6
ԥ��8�����U3M3��A)�A�r2�6����Z~��%��:�<#�9]��K�j��m5vo_I��u5s���g�l$i�A�QY$5$g#�3gW�����I}^X.�����v�;VSt�[�
ι6{+D�r���,Oi����je�Q|`հ��m��mؗx�>����w��R��R��^^V`�z�n�ro�f�%Hz�+r�e�ԏ*�4~]�Sr1�AY�U_.��
�����䙡�!0L���n�}׿WϜ��ï���1�����ȣ�{�t�Z��	�� KukދN>��j�-Xu�Js��&��g�ka�8fC�:F`xN�m�����:Ū2?;���G���)��Z�e�/�5��]^��~�L-�+�j�T\9��|�M�Pe��L$�{�2��)����'��x�1KB�7�WS6Z�{@�jĪ)��l�	�d[B���	1��$;˫�����X��3�^KE��6�'d;k���ߤ&+�QzK�pgӾ[�	��AƘr�zw�r�vT��m�Op�-|/����fGeJOW�Sl���iy�7��UsӘ8h�E�_̼���f���F��WԄv�ǝ	yN�Op�a<rW<���^y),i�`��ٻ�Aa]:�:�]��GS'�A��\���ـ ���άI�X����,(Z��3j�`ڏA�&j�9��X��m���Tk�!�n<1�tYy����&=09�Fq�jéX㭏J׹���by�j�����9���S���X�j/aܗ+�y��~j���k@~ל�+���E��y���Sp�I�Ou��K�.�R�VV)�DGKm���ڗU���.��_��>YW�u�+tVc��&<qm"����2��Ua�֭�\u�d�U���s˨��#e���F\:��� �y;����ﷻ�����}�p+04��(R4 R�	�.{��|�>�u�͔7��Ǿ0��l�0��z���g2=I��	��omw��x�'��c.�k'�LկK4�����¼8ėj�b�ޑ�hT}�Q^\5D���I_!J�,M��o���y6N��h�7x��]�s��;��E�Yy���� �@A��K��;?W9i�eׄ��gO��S���	n����&pB.'љ:^�U�m���/!�����B9�s<��iB�R��<�������)/���sC��<���!ܯ)��4~ߘ�b!��u���^�އ�{�V�iu-AW��dO�㦾����/���C�?4;H�8�X��L�s�-��@<*�p(�7 �j ���"S���g�u������xd%�/p�!]��98A��K�x5�����F�)���5���1~�����GYh��Q7YF�p�����]�7r�����^t}��_8_z{z!'<�y�n�cIL�����N���={*��Y�W��n�eC!�'� �I�n�_	�vQ��vEL/�J.��T.�n5ȼ�Qw9S�1�QFn����m�ͬ"��9Q�-W&�� �ޙ+����>%`�ө1p�Kf�N	wV�..k����B��oX�ĵ��nXv7�F���"��s�zzn��5t	�&��.��j���w%:����'0��lQ��'򪿟
���ahI������>s��{�R����;������li����7H�4(�N�⮗�Qi��a�[�==5��Ӏ�mP�n5ܲU�=�e�{��6����+�I�=%�j��-
{y~h�����H<���C>��>�t���u}�1�*A>����s��K_�ji�Yk޸�31���f�ܡ����aˡk�PKܽҎiWR͵�l� ���ѿU��z?)�"o��މ2l�OZh|e�ۯV��U&!?KގS�ǯq��;P�K�gbLl�a\���k��0��$�B�ay-."�콁���}��]�K���-���zN��-4^^���뫴��"���
�^��pr�(>'Hl�k޺]���kCi�A8s!ǧ4���b�uc�����mY/lz���|�6%���C��{d���������Y���tS��������1b�W����)>{�m�^Y��sKJ
>>K��O>���(<^4����ׇYM3m��P�8�� ��Y�����o
�H�x���,:/�Hż+��l~���Sĳ�5�&�^8�������#�gHmc��}kr���s��}�-t���^]އϱH�:��EB�Jݵ�)D�0.@��Z�����=ZY��-��i�tX�yZ�/n_��S����9OW@�j�;����G\����UZ�U�aBe`J`ZE���(4L�u���V�L�;|�׿OQa���W�G��I�� ��֔�{
�q��zi���-�ݕM��9[�
��:�Kq�qh]��"hyvB#sW����I���+
�,��	��ֱ��ކk���6+/7�o
�k%����k���t�`��_I���>x�Js��Q1`�-w<e��{�s�Z:����8�F:����Ǚ6`}~[b�8a�,9*H�I>��<��2�-y���bޱR(����	�/O����G��M�遼u鶢�'t�����՛'����W��+�]?���'����@G�LkÐ��X
���Bfh�K�v�u7�M��խv�/6�k(~	Gs�}w��v�lc;l��\�`ܜ����GX�
K�@v�R�*�\��rhK�j���'�>�d�ͫ�@UR͔6-ݛd]wb����^k��~�&�0>�����K�so]P���dR�:����b5ָ�����6n�'n���0���SR���B��0d��B�}l.��D;hGVI��Fi��(����6D�)��y�fj%���ft/F��7�U����5₡�ŠJ�����#3d�16�_I"m��[,mwI9��e�37Ⱦ{tz'�y,^�7Ĕ|"
�pt�
�]�[�trO��k}�1]����Hڛo1[�xk��vZ�9s��`W�W.~����*�L(�̢�� %ҠP
�Ϯ�s����:����j	�[�-A�_<3ǽ�9�����X��ԍd���sʹ��N�G��,0׹�z�w�	݉.˂�b�	������6�hl�w�C@�q�10��\^��t�mW��H{��]���>�eڦi���)�A�v�����O�w�\F.����"�5^���\c��ch������zynִ�v^h�(1jd�ԑ�g͋e� [:{v���TuV�Nf^{��0p=�D���t���Y���.z�:�}̄���	�� K�]Z��X�n�gZ���uy閁Qp�W�����E�צ$�H�:ūѐ��:!V��1I�a��j��C^T�����u�C�fI�ӳ�N���?��?����u�?߈Ϲ��,� ��)���<�~KX�4¶�tD󢔊FU��b�u�4.��cz}@�3�AŌ�e�e�1�m�YK���L�~f��ft�O�Q��ax	���].2	�8\
�o$n@�!8��uX�LՄ�K�#[JF>�&�y��� v*��ʒ����c�u�
�j��y@��z��Ϡ
�ѽ�.4��U�$U�o��ٜ�ԥ^�����f́�E����{�!��m:��%����Ջ��GY#�YAf�.��HIdb���u�:5wh(��:�Vf��c�A���"��P�{�I��SztWf���X����J����)!Ro-����vvSB�A�ngm����\l�ౌ�}�T�5(�{(ع�����C��իFɯ����U=� ����s��]�YZ�=b;��:s��ү]��`<Kl���L�TQ�-ԙۓ"�hI�������BZr�m6�"8Қb�Ǖ�,�t.��c8�MޥMЕ����H#�L;(<r����MS��w4㧸��s�u2X9%�Xv^��T��QH+�zPN:�?=v����*`�x�(��\u���Mb���VH-S��j�M�f�8�UXNv[�Y��z$W���7��ͥvS�:Һ^S� gqkq�ph��w!��5�.n����1��7V���mt��rc
��R��1��a��1�`	�2ڭ��0��a�->��F�ͭ�|h��;z��k�oJ�eT,��nj|kv$b��+l��.����;��|�Xa܂�s�d+�6��7Wa����k�:�k*�)\�<���{�n<�cj2��ҪY�Ϗù;��M�����+g���eX�~���Ш��W1$�ڵ�����|��&�7�B����2vO����s�kE(bq����䡴�P��d#7~*��곛��<��X�b{]|�s�&��xɲ3/rTH+��EPn�n�r���0rYY�&�2!�ŕt2AM[�5�`;�j����8Жp�;W���C�,K7W�k �d�7H-RO0��&pɌ�L�ׇ��W¯q��n��)�� 'z��Ņ8��ҹ��Q�!\�J��6�\[��MNK7{RYOH��z�Eɔ��4��XY���`���އS�v��*��Bff��sV�bvBZq�to�7_P��1�&>Klm�\1n375�V���n0��䷏%$�6��X�9��d� ���}���J�	�G~t5�H��*-|7 {)���ਯ�_W%,���NV=��)[ѽlM=�<A
WM��U��3��Uсmժ�/\Qw� Ŷ�d���E0�=�[K7Jp��f���+���dt���qf�Pfk�����$��#y;s���H4�0hu^�^Ϥ}�����oL�Z��>��
�M����N�zé0�C��Nf�*m�yw7*:jQ�n� �)���Gu�V����|v��@m��\�e����3���sQ$v��dDٰi=ج�#��p,�8;�/6��ԩ�8Yg8 m��P�(Wv,�Y1��|�IO~=�վ+�6�.!�>#>ܨ-E�b�A:�p"���hP�p4���ݣ*��p�Oi��wSK�۵B���O5��ù�o}��L
�p�s��I*�3g)٭|��< ��9��`���U2:o��Wd9�3�mkK��8����I�>Z֟ Ȁ�ri�eʎDPP]�moF��R�B�;|{|{N�)�J��@U��Ag�s��v$%r9ɔh�q�ŧoooobwQT�BQAT�ݪ�"j�֞��U%LUDD�����8������"��|J1n�Uʈ�(�IT�A���JR���6PQ���D�d��x��Y��EU4�̴D�P�8\�GeQɄ�!腘p��*
���;�H)�0���Q�2��w�Џ���TC]Z�jju�(��A445H�S�v�*����2b�*��o��z�8�(�DOI�!&=0�#�����T���$�7���kv���;����Ɓ��[y��J�щ�뚕߻F������%>�.���{��x~��x1,T�Ѵ	|2�61�c����2�0� ��P��*
R��^����>��Wq|��0��r'�%�}<hV��L*���yj�q(�HJK�C-+_B�P�<%���#�ԉ��@���/�FǏy�^y�0r���s']�U-O���R��qqQ[9b+�`�f���ߘ�8V�A_���� B��?1���ꃎ��4-[�X㟈8�����R�1��<�'���^:���*9���:��aߤ�B���5�@��ٵ	�g��D�D�3Y��1w����p��5Ι�t�?|�wތ��B�xyX+��D��$z��(p�ѽ�c\�g��א�I������X���0����¶z��OY��^�����c"��漻��E�(�QbbH�=Ϗs����/�ce�?{;���e�z���8A�l;u��K,Dq�}�=�Iu{��<����}l�k|�#2R{��Ƕ�n�4��	-^��+'��{���w2�K�?6�5�gt�u2
�5�Dw=3�r�}a�p�q%����|؂W߻��o��{���l�y;�ZY�(��G�=oM��skb��M����~v�S��>3�B�B�#�.W���z2�U.�U�k�;�R`�~T�D����rbN/BW��:��GB:�V���]sC}u���NS�+��m��j�dyo��S������m$����Ln:8<Û;Ӝsf��fG���NZ�m`�i���p�3�K\���/�V�J�U&Q�JfZA� ��B�X�R�B�C��>����w�\�ߞ1�y��	�J�'�+��߹�2�9J�/��f|���7�����$�\�K�!̯hc�����6x��Ғ�5B*�߄l�=}Ǆ�-��R׭5�S1�L�/��)�?����7��}��):,�ȺA�)�FS~��1g��ӫt��.�}���u�r�$(f����ݗ�D����]0�0����R�mtx�i��ɝ>���G~�KĐuZ
����~��T� gla��(➗窽\]��KKt���Z��֩.�ԜD�P[d?��_0���9��N�#�i����Q]���������-&����s$R���@�^�<���;��`��Q�g�'��O�����K^��MlmJ�a\zW=�����*�Y0�۱b�ɔ(�.��3��D�ݦ?aѳ�/*s�aD:�Zza�q����X��2��A��*}8��dj;r�k�,3�R���It��R�8u ̬L�b���|罨b���v�Q~�1�I~,��s�*+�v���gfT8�l�l���lg!J���Е�'���Yt���@��C[+[�k����B�bw����%c�M\��L��R�z,]R�J�r�>u}��F��:x��.i�8b
��[��*:�s����Ůw�{�w�~y��޻�kE:��(a
�� ���H�H��"%� %*� ��ƾw��ҋ��g��aA[s|��>%�<C�4>"T�{���K	��6q�6�	��v�5��D(��m�t!AR4�E?�@��uY���ԆAi���|�y}&�+H�E�������W��3J]<��r�r���)>y���5�LX|a�����Y����h�!�+O��k�n�t͵{�H
���;(2�jq�d�����l�zǫxT:]��Ƙ�C�|������
5Ќ�OGN0�ޝ������eM^ҚOaWN0<�o��o�x��oO,���KY���u��W	��5�[ ��U�^~����=�f�)2�����F���皪5���b��P
V��X���Ȝ�T���&̞z�)�|��M
�Pg�0�!g���Bڗ�*Mm~���ȸs^�����?��f��+�f
��1�\�SA�Z_�a��O+1�1Ζ7H�^[\Ú�1��>G�d4[A���86�HJ;E��9d�]���n"�γ��H�	�����2�K�9�ܧ�N���h�C� ��-��bll���K����?�,^�_:v=�.��P�o�v4�kʧI��3<����,}�3����S�Q�;)^-Ve���v�r`�C�$z�#A[��(�P�ޕP��_��!����W}�o;��;�ַ׷Y��������"}�L�P�*3  �4�+J�0���
�"�B��ͱd$�u��C�n�wD�v)Ʈ�\�H�P�Q����I�wm|ga���_)�5�X����<9��"<Վ��Ρ�B���L�cPM[]�zR~k�d�ͅs�
�Y�g!�6ԓ/���#%[�4!���`~`�"�!�]�uCs��B�(L;�ƲǴz}� cY�!Ը��&!��>Z�}��b����QhZS��sO�8�y�-������%��$���$�!]w������
��?c�x��Z�^ø�xg�����
H���ojF�GS�*���^����z���ʫ���Ҽ�揎��>hA���r���`�B!�E�3��pt\\lg���h���v;K�]XݎtwO��)K6״��gJm�m�e����<�dLVȧv7���&/�z=�8�1^Ai���|춑㐐qAd Ŋ�!�$g�ٲ��WU��R9��{us��:]���r�kӼ{F@���}��¢nA6'"��.��t��%��,+��{������ݦc�}�}��Xr*kr�'��.�9�2����ɴFB�:!X�{)R9B��ٸ�	F�۞�X-���G3kzWc�M����T��ڬ̷�]@���7�b�If��+%�٥��&��ݢ�]������n�-���'n_t|*���]'�$�h0dO9����=�9�[�G[���~J)2�L	�0�@�Ȕ�B��{���f�Y���w�W�{J��ZU%��#s�e�e�3�rޯ(2�u�Rv��n���/*y����G]Ȝ\���s���M'I)�Ҩ�s=X½�Ш�oD���y�J�y�J2Z�\C��.f$r�֯%�CH��v�oR�ȴzb�t�/I@������w"���:�I_���������������%�a�m�%=_�M�.��`sO����s���7�~V�fCWA�o���
��Qv�-/��>� k��*�yu	ޡF��aG!s�u��^o�Ic�=!����᳋�ӻ�u5��'�ֱ@������D@-��g\�:�̡f���d�,#Mn;c�aZ9�l��H�⵲���Xtr��>OW��1�7���5\5�y�?%��~!�W����ܚ��q��L�r�������'[���`�C��O��(�{�^�ԯ��y��w2�K@�,׫r�Չ*��U��(v��ƥ����.Z�9��w�_�ЇQw'b����n�����f�u{����;�XY���~*]���a��D[�����)�j�j�?6F�cI�K�j�k��+���nZ��}b�+��]�N�'V��Z=�-������Mg�2��2 ���U�T��")��%��zvi4�dֆ'����ɲ3 xQks?���×���ok/ƞI.U��F�ۺ#z��d�;�}���Ȍʴ���L1L��
R�J���� z���]�0T	��>C�|a�Q���f/"������G.�j��x�z��[�K��.b�&�+`38��L�"ˉ�9���T^��k�h��C�W� ��"��"��t�|����0�(e��/\e�5t�Ú�|XP����\���p_˶�D0�Tx���-���=e���!�ˑ$��p�oM� ��V�i�����|����ޚ竹�z�kAj�Ϻ�URū��Jl�2*�hR{�(]���{��
{gd�i&(�ל�q�H��+V�l���p�Wc���P[��<��ħV��	�T-�.�[-�9o
(�X�농�ۅ��w���>T���@���^�7�Ru��K"�s��K�F.��iM
��M�T��Ϸ0����� ͒"�Cvz�H�]�a�K���r�@[�y�n��d���5�(ͪڒ�Nʂ�NZ�Ç؏-�B�li���MzBn�g hQ��N�H����T�C^7]q�g�W.�z/\������\k�"o�����!|t�����/��>��ځn�?��9O{m����h�F��J�đXγ)�B;seA������6Zs��; �v�	�����.<o������]��)@��rX�%�)�X��$�Z�����o�G%�U�M��vn�&U�icރ�k<��Z�;����߆����ʄ¬�R��*4"B�
%(R�H)B��P���O�$���=��km���F��Z��3~�C��,��Z\={��B5�K�0MM�I��#�TDշvwX1��{*i��J��~u�R�aXzV���%�^շ��\�6�k��
��� ����Բ�oq��T"��쟚@Ɇmǡzf�\I������>�z�3�@��1���8����M��}����gߩ�Vax/��z��v���{6C�ϯ��c�^��ٜdB-P�	�|��D�=m8��E���!��1.�r�Cap���f�Y�b�DPڬa�T�C1���yb��I��WAg�>��H�<�Z�5�k�)��3�2��K�$�E�ޗ��+n~�]�n5�~�-�wm3M{�S@���(.��"��g�������>$���PPZ�Esvv5nj��9�Ws�ס�ɛl�J������S�W�9A�f�'�z��C�S�
ɮ����M������i !l�?�Eǧ�f}��5��Jl��Pd�iM'S�l��OM㝷��������^�h�W��?;Ǹ8"X\���yV�"������z%�s4���7�G�}�����z�]]*���k����І:�Y]�������@Cc�g0n���+vl
�{�Ϭ��/q{��t�n;�R��}wX����\7g��_D��8�fig޽}l���Km��aɆ�����A�A���J��������iT�R��R�&R��ej�Z�A��F�Q���(��U�o2�Pi���5s�9y�FCȠ�l�ɢ��~�L�� ����A�%:O]hy�<��v�m�X�v������{��,N��s���>��ПT'j>��Y����nNZ��/���Gn�Z�8^ή�/�"����)Pk�sQ1��ϸ-� �z�M��P�iō��sY�R��y�:!��M��9E��e ��E�r1,0��-��/Qq���gcD��Ҷ3�����C�N&��N�������"�J1�^J;��O���v�v�_��;�3�ޠ�$�w�N��X�,kȇb����s�dS�V׽	>������}�^w
�[-�5c��먇�&���D��q��|�����*P���dR�S�1���ڒ�H�A�	�Cw/g_��t��u�uv�zp���U�VX^6��[�=�s�I8Q��)�G*y���SwM0��:��W5.�jy�HqEV��4|��ؽ�^sM��łjٱJ���z�%���h?<����37F�3E��;�c��e�ܥ��I�gC����|�]f1x�R�Tnf&����a�˫���KIS1�$�5�1W��j���$��R�uծ��i�7���A���7�Y�C�o�a/� ���5�}3�L+ߛ��s��\���`-��E|������P�u�oWEt��w��C���}y��*��)2�A L�(C ����)0����[��J}�tc|!�-�����m�ޏw�,�4��ܔ� ��˴�|kO��u��qd�y�'s�v���B�k�X!0����{���u��Ɛ�A��K�d���Z�Ɗ�b(vqu�m�]s�2-���Ӿ�/��|Ǧ ����\�'�㰂~s\�ټ�j�"������h[RZkY���=�^ʋ�Up��(}^�5.2�'��Ӭ��!uD4x̎:k��v-P�"�s��׎��r^K�"JU�\�t�C����|�ɶ��!�zd��t�V�7��V��!{<ū�$�b%:��W�J��[�[�hU������9�&ƃ[ݕYhֿu���|�+��C^�v��T�g��LU��&%Ɓ�2�w�W~=a�ߪ��_������[cD�P�!��P��}X��5�0S�(�H1�� -瑳s�ף�A45fn�m��=n�����N<àǞ��Gw&�\J/LF+�/7׹8�ַ�d��<3j��-mC	�xwf�w�`�ۡ���p��红����l9������R~�yp�&^��G�)է�J��)�v٩�Q��7��Fˇ3��B�{�^�f�2��:Ko+������+ΰa襁�f:�3,s]n���r�@M��V�ͱ����\���aq+Ǻ�m�-o,ך��e�<��O�ow���s�{��W�&Z�Y�d�dZ)�V�))@)T�Mw���_>Vw��|���̀�����}j��<{\0g>�K�� �c��w���Y&z�y���1�f'4��B�dm��˥k�*=�e���m	��XK��`���'�Wn9X��=$����G�g��zCjY��Ja��l�k�C�����z��{�A�.�!�߳�x��۷���i4ȱ� x��7�,ڜ�C7Y��q�'�'y0���X�U�ߩN�qڍ��ʾ�mH[?:�<�Ǝ�2Dbwh/�,l��#���"�,��@$?%k��$�S�̖�T(���I�"-�3X�����F��B�@��i��Qx�ۯm���$<���g�fޏ3R}��C�tc�b�R&���ۦ�WT�:��L�=���8�,3*�̾����i�HD9�F�4G���$	^��A�,��}=�.�Ȁ\t׫] S��0Lg�]�5U�v�e��>Q�4��Bm�v�bcf��)����ҡI�J�vN�׆=[�O�흎�焣`�R�h���8�}���'P�n}�!��k6���)Հ��	�"���u�!�x2���--(]/�-�n�7���d�$�f�d�-]���b��i�Nkj�C�Sⶹ��5׮�ǽs��1ӭ�kF��e��9n͖q�g�CMZ�-��9N�ۗ�o]�0�L��L���+8�[�.Zro'���{�9���˫��ͥ�I&	��v�n���kc�4����f+�؆>L�C�q�rHC���&��YU{��x��Z#o!�T����{�$�ی|ee��tm�`�أm&XWj-�Ϥ��C4�t9�3;lP����>|1�}.HńS�Vl74�t{t�`��&�z�Pk=�fJ�k1�g_i"��J��� �19o�	��-�:��zڵg/�|�5��#�|@�y'@��9]�-/�7��X{�"Ⱦ�m��ݎ��)X��QsKÜ���ŀ�g8�{���Q�b�#��޵Kwb"�G�.��80T�!Ed��u-�b�v�NY��r�����������jb�S�����w�
LZO9*	8×iK���2ޭ��,n�nט�wu���i�.j}�nJ�K�c6[�
�[结�r�5�A�:>�K'5]�tӏ��K5x�DM��7��g��^w}㎕ ����M�-���y�ݡ/��zL�����M�����ئ�.X�i^�JI�$Xo�v�q�ի��˳����t��BE%z���t�#�C�����uf�U���T�n�Y ��d�Y�Sso.$ĥw�Y�*f�<��!ŕ����D �퐛eu�݂�ځ�D�b�h��j�����'6�Eն�e	
�x���L�-T��`]+��t.T�"���t��C�:0�t�w7.������f�T��}�9顦o��S���"�����SW�vv��h銕������y+eǡ,,���QL�ѓ"�w�����
Y	��.�5��nvn0�ԙ�Y�ց����Wر��"��;�����+�<����w�$	���=�ڕԨ�5Ww�`Z�'�!6�;;���[Z���-w^	��I!�O����X�W�ҁ+�]nu����.vŝ�#���x#��-_Q�N���n���������4\�cևE�vrC/k���ή�^�t6� �j��xVE�nmǯl��.�R��1�}_P3E@/2-ΫvЭ�RV k�U�˵��&#y7H]H��v�[ �q�fW>��' $I���6!��L%0�칯��O.��W�}��Ï6��`l���q٦��U��4��K[�2�a�٦����NLo;��1S� :�c�2ʗޘ�+h9��T.'���ױh��>�6��z�՝sI@��*{�]b��'�x�9B]F�W�v�����f�I.Ѻ큙�Y-���7�������*�q�����tԲe�S��yvڄ�>�oC��_O��e��G_2���y�F�ق�l� ��I ��s���'��c�����tDfEe��k,,����i��j&��ϚwU%M0e�i�����f��-&��{|{^�����'D.Q�G*�\s�q	T%31D�F�
�'oooO���j�/����i:���B���B��W�r��
�2�&+ ���5��v�����Z�5
	�UE$��΄d�N�Zj�*�ܚޛZbL�ۧèi�j����jY����h��NQdk
)�Օp����$��hT\�����H;ז�Z�c���#�aPR�	��*9Pʋ��Qp����QE�:q��L�Z��h)��(�d�tx�Q7��\�N�nS�SK�:ji
Ԛ$*�����RRR���$>�Z	�x�u�\�Rg,�e\�]�
����iʈ�7��2	����<�a9>�﮲��k��:�t��{Oԁ�u.j.�vY̊[��ѥsއ���B�fen1�Z�g3�I	|��}3��#0�,�x#bP��jC�f�h���J�
��L��ȩJP���?~`[�?	}��p�[n��N�w��'�!�	��G��oD$�����"����UA�G&�h������о~�>��t��5i��9m�Gܫ�V�X1��H���1^��e���mGZ���������]>&QLqt�w4�IU����̜3���=B1��}��7Z+e�6����zSp��]�/gut�f-?2NX�w�,!޷ <y������\�bo��;�(�	X��+н��V�Q�̩�К�`Z���vJ�/V����*�K sIzp�|�q�-�)�����{j�we�>^p�\�54���Z�t&U�+�J�)�z�"�sHWR͵�`�4%کݪ�D��]��`�`� �2~k�L3n=^��*S�:�,r�N=q��hʵ>��
�}6�<���Ԩ��@ߵ�(�������jj�+�g�՛'���E��s�e�_D�U����m�u2�.��\"�������4>����f�X	��8=�3���{ȧ7����,!�tj^D@"x�;H/��ӭR������c��u�wO���מ�m���/k�A��j���Z�q��]">W�넬�fN�>��a��!�ȹ�Weq�Q�P�
Zج�>4hM�֮�Y2@�5B���A�Lz�:�Õ�oR|��S��E�fM�gwm�S ���������
��_|��{���Z�f@i�)fA(��fV�&�(A(�Z�����������#Np�o�p�4�d��VPB�).���~/��­(�|}�}��:~��@�~�����!�eO�T�S��͵J����3(2�jq�j	��3g�ǫxLXaQ���<deR#����y1���".=*�*��Q�>�"Z�A�P��{WN0D"�h���Nu��.�R�Z|�ZĘ�s�2.��S~�<(F*��A8�8ĲO��۬T%Ќ����Um\�o����_�����<C���=���26���fʘM���A/��7J��[�i�g�_�o���b�y���"�RF�[>�sh|��\�� �6��N�|ʩ%x7|<6Q�����7ɲ�0ڸ�p�z�$��S���R���9�az|�>�E�� �z.����:�Yu�a��4�ɀ��jd��uL5�M���-?,�)���3L$��9�:��-������#�c�"|��5��H�ݯ^����8�r<�jF��I�����I��!�jm�o���c�O����3��`0>��<�C�>��:�|�΢`KaoA5mw�)?5����dS�2��ء����3^�� ���#pZ�so)������Vv�Xu��n-��L����n�O�p��3��wV�ATJ��h!��#c��S��#�e���j*���uW)h�k�^v�c	s8�=8��VeLR]���Z{�dL;���������J�L�@Ҥ�4(̀D,­"�Ĉ?Y���f�{�Y�f%�ݘ���:���~/"��zP��@g��I�0�]�Y+���5k��R��t9_��{�U[O�P_��_�d�q?��i�*a��OPn��ˆP���^����p�t#��N���aC�@��+��
r�^ø|�Zh?B]���=Nơ��8��3���A��ͣ//mf��o�Wv-$�C���sͷ�$�ȗwUZ]T�5w�R�w���	/���y�P�]d��l�X7�ћf���t�v��� ܌;m�5��=���A~[U��#�y��I1�X�|¶�Z���������V7yt++�!-Ed����͚���wf�_-}�;Ю����ﱣe�%������f<�x���V5�B}i�N���2Yv����Ǆ���n���(��q�A��Ơ�Sp��� �d����nby�Q�ne�[UO&ui��gT�<a�qr�pb87c߸�'V1*�*��\�P�^r_�5�=>���e��H9��7Aըf�{X����-�^K6��76��L�و���T-X�E8����e��/e���Ĩ�=��=[�Ѳ����f��oQ�a������՘���ʭ���4�/H�l���K�n��x<�ib�Q��A�j�I���i�[Ї��v�������mZ\c�����r���ۡ�3�q�5��!V.�s��C2��+t�s���}����Lg�#�*d�(
BdJ�
)R�hA(ZD~�����n9!�o���!�6ȭ�doz]��z�+t��&*ۤQz�\hg��"��e���&��$������#��"�S �y��,�v��ʒ����"� >c��1�ה�ϼ�����1�[����%y�`AY>�^�TS����t��_�.�/�O��\�g1<� �jij���z/])�z{������%�ƱK������D�^��W:�r(ڭ�P�K�g|]٬D����E�z�O7��4��Zk��Z�>OP!i��&1]��U�Q�[]��E�ۘdW/:��:�ǥkە$�5ʊ�8�-�6���.��_�b�5��xZ�����>��>qa
��1�i0桉*�t�=�1Oe����|6��N�)�̭g��ȸ�:��{��L�[�L3$��f���� Iv��]��D18�\F&��i��F�����3t�sj�Ϗ>׉?���hy�S�W�0����^E����ًRU�dS�6+�p�����/�Dg��rt��~�	X<���ـ�3%'�
���=���5x�Ym�x`�<�P6z3i����<�n�n�4�&O?F�^��W���'wY^"���96u�x�#7��Ɩ8���ʑ�zZl*;��ᓅ�Ek%^��ʾ�J&<{Z�\��9��]&����j,���fS���h6���|��ڝ�t)�j\I��:�[��햐��	�	���J(
@I���~|�)b�h��CX-��� ��J�!˧�n6�5���\�ρ�
������b7M�0ќ��t����K[i0?;(2��R�`G�={zm��sƶ%�<�^}e�9�Ml�YMJn�vک���>i.��u�\�K�����d��It%v��fz:w_iᶠ���ٵ-Nb���Os6�,�tss/�09	��CH�S<����6ħV��	�T-x��ݡw8�S�UJ�s�}ǆ�N�ǘQC�x+���?ZoW�'�����j��������;���
^���Ç�<��������K����4�<}�;��L�8&9��)�3��{��l6ı�,�;*�NZ��mvM!��#�&�	�͵�����䥈�?g!<��E�U,U�����֔5�K�5''���C�̅��S�[�x_�0��ye�vw���5�zT��	�ٞr��е�fºα�6����8G�\��\؍��q�v�\z�I�f%�l��V�a#�J���K�Q�!]K��ֻ�Wg}0A�A�2��4�b�x�s��a����rɕ�Zw�
�R2�ݪxmg�1��=�ޖ���ԖL����,�[:Z[ϲ�
Ъ�t��i�.���
Lew�Aw>����퉓a�1V��黰R��
s���ȅ ̰J
�(����V;Ĭ`���
p��s�A�|�!��q�^��+��1	�^�r�N=X�v{�u�,����/b�e��0G�B���(�]z�+�Sߺ����l�m�_J/���h��cּM�wCη���y�r�(�O���-���þ��h|/K����3巚~���x'��P�Q]�_w�I�ǻ��CH���D'�z���E�ڔk��%��������y�ή�%M�M�����/X����i���h�,���K�y�i�m�^Y�=�d��������@T���Ai22�X��Jz��͵J��� �����/,���;�Mc���Jv�4�%Z[ٛ�jP�JG٩�x�Ň)�Eǧ�N0K��W�o)�� Ɉ�����հ�&�	��s<S�i�ꕉ�%x�Z�OUX���e�p����S~[#sS� ��
����te���v��|�m���%�
�&�o�\�Σ�"����Oٳ �L�� �����I��;0nz�e�Xy߆R4��by���NoT�eA#I��7'��}��K�X�a��B��_��^��=ѯp����OxaR�
�]����/o�¸a%�����&�pn>5s=����s�s���h�\�:Nne�u������.���+�պ��w
�e6,���qѬݵM5zC{��u߳�t����v_p+�D#1�n���/�qo?����>1#A0R�*L�BP ג/������C]\3�vOC���|1���n��Z��l9�����}��`m�F2f�9=p�C_-n���D�Dhm��-I��h��M���-?,e ����uy�p���O����ML����!o�=05ÐEj��(���Z�ge�Q᭪b<�w<U3��p�z��5h�/��u>ii�~���>�{��v/ƇU
�P`K	��������U�F��8\L]��V�~��?$s����UBr��D��A�x�<yF����#�w�ƅ��m;�wo�n!G+�z_-s^ipFz��k�g}��ͣ�M�"c�@�����ӞJNTV�1���׬�[��[-=>���A�T��l��
Y�Esװmx���o��5\G����!zl[�ly��W�[!]Y�ܬoP~yÆ����@���-Bt8��;�j�~��+E�����t�����u��4PP�@��Σ��i�oO���3Mi������˴���}�f�/5I�or����Sůl�w��E�aXC�k^=�7�}]cv���Aƀrb����/�z��ǀ�&��쫷)N~�`��	��ºb�On���{(�J�{}�������`[�Ŭ�0|��!U��Cϰ���En�L�:,�U:����C��JUmZǓ��Z���{C⎫���Q��M�",^���R6{;��y����{�F��}�p3+0���;S=��)ڷU�b��6q��@��\bUc�d�)���DW�.z�:ƙ�ε����lz�cX��.��Į�g��|l��s��;�	�Ո��+�by��y�Jv�M���v�]΋6��M,��·D��E'X��Jg��S!sEM}�[����L��_){����i���Tm�M��p��M�^��=��Jt��H�TS�~�a��ЕWN󩴟l���rշ����>��O��2�[,���v��T�ax	���^�\h�+�=mڭyu[˧f�V�۾U��`�`BF3�	��#�o�K*�5>�WJ�@ȺC�䇨�f]6��9YB�mBYh��^=5������p�݈n��%�?G4��I�%=�B��z#��Vq�h�v���'K̈́����4�H�VQύ
?�˺�'��6����0�0���Ν����']��k�K]i��Zk����A^O@LA�4+Գ�&j�������?�O�r�u-T-_�J�B�)���zTsK0[Bi���]0F`Ϸo�P�Q#�PM�?8����e��ɷ��ct�sh��CG�����_@̱}tc�L%�VsB3\�8��]��W�䀣��ǖ���:w������I����������-,m��C}�,�ζ�#��伌��Iy�czb:�t�J�<�s}�o�4r�V��_b�lR��3"L"�B��}�=ߺ��w��������<�^f��Ai�}��f;^��4�ƕ���Mc߹C��q�nj��^��6$.��S���l3ʩ�6/��3�[�L3$��G�ۨ7E�{�g�ߧ���s���U�<�/��/3�+��x���ڢ_ �,�֡���(l���wBG^;�.��}�;[>]3ttnvytQ�v8�`�xc[���`L�!\O�2R{����3iUm���ya��L.�x���m��,���VHB��M�ۦ������K����`�'V=���Ǽ�[P�z�9�lNT��xw)^��A��B�Ru���PT���Jm�xn	o�w({+�w8Zּ�b`����3���KsW����|d&T��vл�u�2æn��	܅[��v���!���:-��ė�p��vW�i�y���Jce�S�	I`�OdR��=�U��]�/�i�M!
�=s�<'�o��!ŴH>W�+�Bz�xk�7�Ru�-�b!�;��y�Q����6[��+�����s��`������;M�E�~��=��	��|W��K`��+,ޛw�;*cԏ��w۴���Q�n��,����)����lM�+5����s,u�G�xQ��'w�h�����{�t��d�,�'�f�5�D�mv!h��k�m�t�&[j��<�\�K7�����wc��厰����R|d&"BdfT)}��7{���
�������xE��tS*����`����TX�|��?>�ٽ��z��=T_6�ء�KZ�B��4]�S����� �45Iw栜K�k��#�X����?j���*�9�hb�F�L�bK�	�LV�.�*��Q��l+���!0��{p��j�*�l��.���8V#Xd�
<����mM6��Z�_�*��=+^ʂ^��ԣ������;f��u�/�"m�_S4��܆�0e�:�B8����Ɖ�X7:Y�{����ϩd��9uq�n_4I\9Џ5띈�^nY��}�	�ah@}�mMY�{L��5�tO	.L�ė�,6Q�i�Fߗ��z���;+�W���-�b����Q4�������]�:�l�&�b?����7�4Nmci���	�ǩ�Ny��(#t�V8S�������¶�ò�(����F�_�9�^��X�파�����i���YA
�%�<��m=y���/��h]�L�W��=�y����kh֘��~�U>�zܙ��.J��� �ڜ`Z�9A�_����M5q�UR�c'Q4�w�l܂)����ڊ�ӻJ�^ r+�#�	RόpDEZs�7t�)؜E�������vJ�7���1�YT�6n�˹6��A�y�-���Wt�vuȟs�}��gi��4ڲSNb�@�u^n�?Y˭�	��-l�\�w��k��4���ò1E���2�s�t8���s-u;\�J��0C�w�>�N��\�A?��|��|���ms�*��TseN|voh��1�������%,%|9�ҸÝ�m�3A��B�yD�!ٗ֙��.0���f�T��o;c4�,���69��lm��x�\��3��Ӱ+j��yW�r�(!}�N�9����V��{pt�.�t�2��O���V4u�C �m����@kj�]���Z��C4�]�-.�m`lw�va2��"����H�?/e^���CB��Z;�*�*�)}1�t��)`�]���Ԗ���v�LaBn=�Q��b،r����)6l��W"&�A[�m�%�˃;9�J��ԛ�2 �>�gu���1���D��^j�\��z����Lyջ���l��m9B�z9�M�^�x�of�z��(����A�9�&ă;PR�4a�PhWO5\��-��rW:ޤy��󕕔V]�ó���p��}}�n'MfMiS,���9����:3�PYˢ�n���W�R��í��v���	����C˕`Q�Cv�(-��OuqfAY�ۈ�]B�X7��P���v�O�=Frg<��X�/�p�3� r]�:�NV[S��ns���Vz��M�fe3�q�x�1&p�40joY�ܣWB��],�i$��t���Ɛ��rȁ�F�q��ݽ���@.�{goc����ڔW-�n3�u�u�gu(6û���kU(D��(�6zΩ}��v:)��s�r�۫W��R��u��M���K;r�\���7�ݺ@f]p[=�r	����!�iL7�Y��Z�Bjݬ)�Z�]aɫr�.��tƪ]B�Nɛ���]�
�3r���뇩��f7�+u��`��ݩE�!�V���W[�s���Q&l�H��@v�յ[O5�'cl�����ڵC���զ�=1�%X��kt���Vd�x��V�u��mNҲ�p�)Y�j?��٩�o�~Wn�M�A]�bw�%�0>�*��ih�[�R��	�0�����t�o�ִr�ۉŚ�z�)�w�Y|���Ȕq����!s�����ÄG�E"2�����C��b�����nsV��$*d��,v��6��g2���!�N�ҫ��Mh휷ڽC&M�U�Z�Ɗ�Mu���Z��fumH�;�,d����Pip�ZQ���u���rt/�q��u��pK�c5�9V�/EvWZk:��.�$��6�ܘQ�����bˌ�PBV��{9��}`t;��b�R�I$�J�{�:�s�y�����h��QE%XC�U�rA�DTBn�����oN?N���;����z�\U�\�r��(�x�(��֝D������ȱI��O�oo��op�S��DUU�Ѻ�CI0��%�.�{{z{{{C����uj,��.� QN&L��PU<���f�ą$��������ި5%[)5^�L�)��G����AuZqQ|Br��8\5�fP���$��Be�s���\"."iQQ�)cឩ�W��R��Ng� ��*&QɑQ�()�%��j��`RĔ0ACK�iGe]�)�Y�H�ք�8��|t��'Բi$Fp��Aj�ѹܘ�I�k2N'U �AA@�E��	Ep"zI��Y��J�h�5:��A���^^�f;��Ӑ�8���,��qwVw�w�]-&�!�q��*�c�
�5ufv�ĩ�Z�쬨�߾��
�+���,¯^;�}s��þ�9��Yַ�����h����o��X�(ןf��,2� �jԾ'��)�{���dݺ
��
S�ǰ1�з�xA@�"X\��`�1W5�tX���aGU+�Կ'���ej�&���sz�+�%�y��9�NW��}_J�Ө+�*�����!��7���>)��L�$i5���6��.P���0�m��9�ŖM�V���)3r���"̳>�L&wY��E+�R�'�T�Z�ߊ���}�����w�j>\}}{���k�#�&��cs$^�5'��a��6��9E��e"	����N�{�+���D���6fes3�>ϘE�R(֘r9ó�ױ;�@7X�����/6�k(y��0IjT&mc�k78	f���k��5�^Cc��@��w��T+�\�ƄV׻�Ԡ�by�挊�E��U���&M�ߕϡUK?�5�ܝ�����ZC���������[��U����w���� ��^PȞa�F�״z}[y�����@����Cs9���;���C=o�Wb�$��U~v���,���A�\X�vg���U��׶Awr��:�Y���
k��^��;��fd���]*��:���F*��]e[�fm�uؕ˝N �ᬸ6�U���s�b�n�;Pֻ��k��2L0@&���><����m�_��}}�m�X�\JN	85l/Ic�_�θ�\-xו����n��W���\��t�L�Cb���9ͩ��Hn~���X�5n�v- ��q'DY-� �m|yJ[��7}��"��ơpD�Ѓ/�o�~�}w����^�����4�5�O;W��d�b�Q"r��<PZǺY����=�o
�E;�e������Ww���B�⢒��Sn�hg��ɮ��'ۋ[+Y$2&-�Fl�*���=;Ǭ��|�>c�
�M�>ݥ2^��c�0��]�k���=���Hxs�v9��Ɓ]Z�o�YQp��fA>����(���a2:��U����~ޣ�:F����x��o�~�c��N�)��QaMAvN5uEê��3ױ��V�����L�{�C�?���O�G�����?d����$�����T-X��qӌ#n�R�P�VŶ�����:y���usz((֑�p��Y�4��z���}j�,�:��7�kK�h���1�pi��������.n@��i�!?T�#���2��j�`��Z�2�a�_������n�۹C&%{Zyx���Mi�-fjP�μx�kwӝ�d
S���om֊.��ckV��ȫ��3�gٺ�$j���z�:k�zM�r�h�3S1t�`A-�����31�����=GD����¤2�>�iճ�Uл�����|�&R�(/z���>�|���9�n�+��L��?]x/��V��'œ�� a^a�n�K�~�'�ƅ�!�i�/�rϗ�6�"v�aHgOs�U��^l/����}���&�/q�P ��/�$><_L��ϡ�yz�z/H�3o�w(Yc�V����k��ʩ�^���sۇ�<��5�����u�!������e��d4H���q�j�J�a�J�)�zc*9���'[���H[��CSH��K�3u ��<��kH��_�mK1��_�9�� ���c߹/L5m���,ge��svч7J���C�ր��@�z(�	���p:�']��݇(��8ėc�I��I۽�u'i�Kfa�-lk����חt������V��29�LìY�S�9�A[wpV�]�:�����x�4�].��U�:��e���!'�ә�'$�o�:�n��QOL�=�y��W� ��
�W#^k}�M��$	�u`tS<{Yɳ�-�����_��[��HP\=�M���jV'*wύ~2�-{aTe
%Oj5�q�^�z�9�}m飶��{fsPv��yS��M���JKX	;P�FΌ�T@���+ 	r�엶�e+ "���)��/8f}��r��B@�觶#��Ė����R�3Q��Ih�n<���`Z̻W��i��!Cn�h�-�x%�B�E��]����l���o0�y�y��H��Eeڥ����:&5�zBv�1N2W�ږ�.%6_	���'��"�e\ꮄ�l�ԝ�I��s?�m�6C���0O_�Y	��=���?!)���N��T��>v��Z�>�aL�%B�6s[m�@��x�����(Lɤ__�gJ}�ͣ���}%�a����[���LJ3�9s�@�7���Ky��|Gܲ/ْ��k7("�������,�10בE��R��ˉ�W�n���@��T_��N��í��{�׻��ـ��Ln�dI�4��P8���֢��ZPX��%ߚ��w�p�U��E=>U�Fm�he2,J�`��΃�91%�t�>�*�J�/^��f���zY����L��ې}S6nV�{���C��#D!��G�9���ښmW=F<��Ҝa�L�~*{�Oklt�<aw63�m-��Q�f%郕���Ç@x���C��iɆmǯnt�'*S2q�%I�|e��w�s�R�|^F}8��9��nY�z�p�g���<��{ڀ?J�YkS`��餝�y%�����c��s��).��zs�`���>>Q��c��-g_h#v��& �6\��^�o7t�+:�M�p�;ʢB�\v�mu�F�V*׏�Y�zU�ݕ�K
��&���X�!Rĥ��A����R�W����\�^�����2LHWg_9��y�?>�c�vOί���Iz���;(=�P�f������г�b)@���S_v����]�i�њ�s��df�0��i�C�$^�i�[E?��Muc�VK=�����yլP������#�6hr��j�|�u;�~��CL��Qi��,:���W).���m=�;9�ý���u��]����
yg�����:H���31��ۈ�й*f�;(2�jq�n;q��خ&�r�[c^��t7Cz��F=[�WH�x����"�O�����	_�b�;�JlT��uN2����;��&7�C�O`��z/��/)�����2��4D�Ɉ	��GU�u���i���;={��5S7>���%�t�K%=%����=������01<j�Ml?/�yX��s��\!8�ӂT����^	$Y����'��Nlj��3*H�kgێm|��U�8W�J7����8=f.�|k���5�|@/�#��<Н�i'�b)9X�"�-�a�D���e���nr�jZy��
�d�a�!������y����i��ڞ��q8�Ny��y?1�}���>H>�Q���42ql��tۤ�q����oW�\�{ml�2�N��%;�YI�Y���:�E��\d���CO:�|Z�E�ps�`ք\�S�PV��`]�\�n�љ�ӘL�����N�W�	��4cu���Pٝ=�߁��7��]c���*���Co�X|L�a�Iv����`�[5�z%���U�vvQyң5�%w4!o�����~Ģ���*�bC��H��
"�0~�vOƺ�W:�X�	{����4�i����M�~�<���F<�+�*�f�طvm�`�~a �����#[�8�)�̖���{y���Mo�f�S�a��5���]>��&��l�����Yh\Uz��]�$0Q�~���^�.�zX��0��^�4#�a����
Zfz���E�[���8O�>�z�SϾ{�ǆ���Åcό?b�i���W����̽��E$<*N'd�*>���~f3_�N�f�� �E�5�&ubzq���G���:?_�]����
Ϳ�m�%g=�C���FZ�|�R����iA��|ql��Uϫ�v��U��([^K���;:�/��2��Y�CRFq��l�*ŕ�$�y����?5�������o3;�7hn)�m �	��M�LJ��r�Om�*.��f� �eS�GA�Ƿ|�&��ʹҹB�հ���{Uq*uaж^؄�M�CJS)!���L6������$f����'\0�D�W��+�C�|U�|E��#*�)���Z��{;WGA���Ă�e9�K*��Ϋ�>N;�̺�
|G7�=�u�xD�Z��bb$>u��qw,�������+����v�3�Z�#y���,{���ĨR�TXS.�����k�8rR����g�#�Ѱe��cS���Y�vAnm�\Jd�D���IW���E8�Ọ��m~��W��33��A^���	1�C�h�2��f��/z]�w�Ze�/2M]�ϝ����d�U+�[9{G;jN�#A_��^���xa>܁!�B~�s��	e@v��ӱj�\��3��]Ä\Ǥ�m������0}���s��.+�+?>���	���?��e�<���q�1��yv�aK!s�u��^m),k�Ӱ�'>�Ƀ��D=�_���ߌ��I7�	�2��n�δ%���TW?X��,�d㋰Oy[��Z��2�u�j���{p��k��Ӯs_��Md��ͥ��Bv�572��^� ?0��g�Ԭq��=+^ʂ^��G0��'[.�CO��k.-#n��X��p?���3�������3-��,9�aJ��˦��;�\�f[S�չ�2�&X�����{�L�w���	�y�6߯*Y�u~�n��(�nI���Þ����һ����۷�rc���x����'�y��F~ڐ����ak�y��}~���s�mo?Ml��и�]⺢�-.v���4�:p��[���Z՜w)>?�.���}��e���{��{qR}�h����*H�o//�Eof�~y����a�q8�2����WNǠn���)�i��Ƈ@�r��اy>��0�~P�+f��E���,_`#g&���ϸ���ǚ�^J �iڼ�E�P�xcC`3`.!��pY��dL�#9>��i8z�an:Qz��;cE�$Z� ��
�W#^i��t�=������F�̟B���'�=��t��.�e�h��2i<��J��jm<�-{aU�G�o`�<����Fi�CS�e��X�t�}�[P�E3ƈ-�8&I�$�W��(ن��8�%6!&Bd�H���TbV٭��H��33�hf�u�V��Ol� �ҜI|�L����CH�y�����`mMP�2���f.͘�os��,���o���	�|w�-�$2`�o�61M���Rd�mgKt6�/ ���3�it���W�4�P~u�Sd]��Xե�<��_!�#O�~�昊:q�#m3wRм'��������0�UI.�<�ዩۨ4��6�yü��Rm����vU�Ԍ�,v��b�Ѣmz`st��B��4�ך�mWK�{Si���Ae��ߛ��K�P�;u�}e���Y[���}�}w�>��/n���d���Y)��^R|d`k̋	#�v��
�q�+&�+7^=����s7S��\�U���4sc��k�l�NHܒo�5��Vo
�N���-�}��7T�@�J�g)]�������o7�;P�I���=y�>b��G�U��M'W�,P�r��%Q��k}<�f���uZ�ޢ���j�t�|�QR�C/cӇ�^@q ��
|ã���οPښmW�=E���	V0�=+_g_;�lC7�􋻃X#�\��u�]xW=0}u	����� @�ØO���h�������nt����h�ؽh}�;0q���M�_e��}8��g��ܳv
>���<�z�H�@g��gV��Jo�V�{��C�>�;�� �ƚ�%~��c"�I~���@����:"��u�������/��~\^��̓�o��E�n9�
i�I�I���L�$�Ư4��$? t@#�K��-� lEC�osJUVa���U�OfC�s:��斝
L=�'�uE��ޑ�yfY���K�VPB�).��U�ɺ}8Jq��4�u��/6�ӫ�M�.�^@�g��s3�}ܙ�\��g�t�vR�-\�T�_�u�{��[����+�����ߓ��ռ*"��0��Xt^D\zz��ӱ^��̗�<�٤U��n������pb�ҚOaWN0��x�oV�^�o��
7���_(r����6���(�
�CS6m8��l'�oC��VVgr/Wgb3�R�;r��dQj,�Ӣ��shy}�G�!�L��캵��WU�h#|bJ������B��򻆋���6��(HD��As����]�Zj�a�j�Fd�	�ΨI�G�������y���=c5�] �p��z�W�������wN���2SJ�\Du�5s�:y��x�mhӍ�tU5l�ݷ���l1x_f�8^��zs��.�R)�0������'�<��輊�vn\]�е�(d3cLq�m�1����Y���0�{��N]�9H7H�Kk�sLW>�v��;G�qz#����s?N?��>�h�"=r!6צ86�������i�M��Z~]�D��Z+��4�$ͨD��^B�f�p��a���+�q�����ژ�����2�,��K
%�s4ٻyK�kt������t��^� "�k�ѳ��WU
��U�9a�����y��Ν������5$d�-c�o6�|ja�/��ͺ��C�!��Wg*�]����>ou���u����J��
%0�c�^�˧շ&����u�lC����u���S���v�mz�w`V΅�-*a�Н����wyX�{t��l��
X��+���-�Mg`�⢺�+w�[�XH}�&S�`�	�D��;05�#��s��"t3E����-4`���C�ʹձI�I��"	��X6 �b��J�	?^f&�6%�/jf�<��uu*�+�ZR�g�wY�-�Hz���b8N�˝0�b��Mma(o/x�N+kc�gh�ڙ?3�E�֑-Y������M�x�M��X���������w�3#���T�!����g<- �1ڛoz��T<���|�'g�L�r��H,�݄l�g�7ID&D�Q�=O\7�+r��Y�`P��+h��Isd�v!�
}��it�|�{b��Y��:���S���ُ��5y?%�D�J�-x����1c�fMC`-1��*�H,J�?5B|�e��*='���{U��x�\��\�6]��yAlZ�uܭ2��*��2m��j��sQ���;Y��g���6ܺ�v�Zv�ån��>�j�{�N�Y2d'vX��oq�{fgh��p7�T�aRK9�9^�
U�|��qꥴ�U�i�y�ɉgc�8[�[��#F��)��+Y](�(���+Z-6�F^Y|���C�q�=].�\���ٰ��GD��᚟�5X��*Ì��ື�����.f�'�d��j񁤫��g� �*����3
�cH��)�o>v���1}s!��17qRK�f��r�N�h�rݞ(n��^]�.`��E־v�8H�c.�bvK�XZ���'K��e;X�ĳ5��)#:��)k_c���C��@Z&屩���[�d��R��;2�N��\�f�XF͎"� �(�
�;��}����My�zCD����#�p�Ԁ�H�d�T���fi��m��N�ɲ	�W���jS���\ɿ<3a��+n��s�颂F���-giЃ�F̵}d�Љ��ܺE�-�aݓ�%c���.=�Yrr�+1NoluL��M��K�#�wy���I��
��U��������vip�Dr
m�o�)�.Ǖ�bt�l(c�ή>'�z�=�ȆP�������G��8�9�͠�u��Tk�a�;�^rn��Z���,v��+�XL��L��1�ƞ�ĶQwtʔ�t�"sk7�͡2��9�ݩ�,��TY�;Y >�{��86TGtpٙv�M�H���6�=չ7��ek��9�u������I���Y{D��q+t�ٿ���5�ξ�M��b��tү��mE{�1���m-��L��I�s���T�uB�i�/i��,���#8B���*](5e��dBH����Gd��{J����	�n���i�G�J+�AY��0C����Ma�>ojl7X�;Is����6���̋�k�9&�ԁS�-k����H���w������A|��A�ҷcB�d�w�^qZ4-.7�o)�wmo<����՗���y�q�ѝc��8*�>͘�7G�iY�yٯ���>�3^�n�)�E��w�)*W�˶uP:��}� �$�H��w2^E$�N,]Y;v)���-����4[7eҦUFw���G���Pju�5.�.$=��1ZE=�G6Uwռx����R��%15��M�*�\�^�Hr9䬞�A��Z�F������V�R�HC��Օ�®	%gk��.�9Hr��r�Sh7.��$�������5���N�#�˹r��p)���]�뗐�xW��ƕ�������������<�V<��{��T�t�YǺ�Q�N]�USx���*e�ҩ�,����<�I���SԤ��9�.�p��HM��.^t��ړSZ����� �޵RS���T�{���O�!�$����ꓫeӷ��Չ$*��ű$�w;�P��4M if%I&�'rz�{�r
,��'���y������N%}$��<��y\(�]'3�A(�p�>��ҸD�DEZ�T#��E	nyE9�NBL'X��^����8�x����w=��΋7e�c�.+�V��H_�VKqష����ݴJ��'�V�Zl>�o�ynI��.�s"N�+�o�e�-W��ʶZ֝��{Յ�����������4DK�)-臎j�zaF���N��W����Z<e��N���i�{z}yfY�"�51jF��9ND����N��v;�#�5^Z�9������"W��$��xCV���b��"�!��aC}�����
~w�?}%�Gi�,��$2F-�se{]� �xNZ]����5>�4
鎡�T�eR�9/L���'"���A>����u�!��f�>������	�/V�χ��V_�k��܆x]��9��t���T:!X��S��P�bUԻ'��vgE�uJǤ3_����杪[K��!$��?Br���`�����|x���d������T-gEje��F���9�e��ӋB�	��"�t�z$Ƙt���2��f��{��;ԩ2�qp���]�ⱯO;u�mX�)^�����;�0��B1�C��y�0����f����[Xy�����{��r�d]`o1���^�\��\W(Vk��}�C���fJ�Q��A���]�Q/qy"y4XQ�\��j�����~ʆ��݋�kTAa�����j.}>�C������6�cʊ����w8^�s��N`TD��ƹ����ƥ����r<�ŝF��ZSu���i��%XY����G������}Ң;����.��OCA)�=�1[��i��<�޽�U�����7j�?>�7�������I�<Ym"�OATRsbNP�`9��.�TXW���c7வ���}j���md�P��wu�e�k�z��a����Al������4-Xu+u��Z�⠗��Q�.���.��_[.�sT\�>�,�ǰ�ٰXB<��7Ah���f��΢Ú���t�<
�2����y�tpk���Н�[�mSk.qE���^�?�K��Z�pM��	�����Od��+_�b���-^i�SI�N����m�����Er��c��$����P�?2J���rk�D�	�y?h����fy�kzA!�%�].��U�Zgځ60y�;)����/�l���_s�U9.�a^�B;e�UE��_�b��/! �ݎA~�Y!
�y�\m�j鋇X����{��us��>��*�}�}�+�<�U�ѓM����u�dVe
7���n�wŜٞ��_���P�����yDo�ضx�G66r�;�k�-�>��a�D&��!2�76sV<��������m�M����L:w_mᗶ��^�l��" $'��COb�kI�n��x�^���Wp7��1�֎�pʓT���fݒ��XVn���/_0ŀ��fk4X�X�!��ADrv���{��h`��1:H^�xTM��E�t0�z�'#��4�d�v
�̶��P���觵��]�Gw�6��o�>�ݐ=r'�?4��vg����>�������w������	�"�F�cֽ���{w�Hql���ԅ3#��vv$p}�A��!�{3��zd�X�M4���/��)�sP���?*�� Ǚ6���y�*�3���G��Ys�=��#5}��Ǆ �5ܡt�yT��tS*��:�`ۖf�Q#,olI�U�1������`� (d3�	�Lm�ޯ
W�����z^�(���䠱��K�6?M�Mq��<�Gt���5��ad ����ㆤ#��A�����#�g}�.�Te�>��,��sB�2M����4�*A=��i`��?j�SM�:D��&��zv�%Ǳ���=��ڕ|�#���q�T�6VŰ}��3�a�.򁣫����X�.o��٣�oF�b�:������q��m2s�*���P��'�����˗I�b&�5>��n#ء�]eCk�R�}=���鿕.,m��C	�E��6ő3d�O��<Ļ�� ��MW�+�S���}f�ƾ�$wPn����6��#�h@28�;I}�΄��}Sn��D��>�kd#fǁ:lt���<��vyUu��$Iy�s|�,�D��f��^~�v/�w���i.L����0�o,��-+
ܰ��d�:����5��k��b�e%�'��n]���M�G����NF��V���o`Co��?<���o3y��o�i'i��p��.%���[���r�={�/�oW�^Y�i��%�P+(!���CE�����~V�����^mᱡ�z����@{�Nf`[O<ɛj\�3R��[�i�!f��:7*�e���A�hT�O-�������@�zXa�{�\zg�f�M���۷w��UV�Cn��xO6_A�P��E��t�
���M<�f�|>b����k�.�Y�;�������u��#�3�������I�#4����*�}kJ���r����)�Ϙ?S+��2���~vnBcXl��!	���A�$�b%9�"�P	Mmq�!�W�׸BKj!�V^oC���{Cc��
��K4��i��f
@ܞ���)9wM�l	<����SF�u���.{���߭x�QW�c]�����u7��
�_�y_W��޾�����j[0�d2������F-�e ��瑴W��G0�����B4�ڪoJ=_PB��k"���v&�;|�!�=�5�2t���>;��8����c�Q��zY����Y�����8t|�}�k�ou��9Z�ٜ�6�Q8�]IQ>��}�ԡ{�ޞ��� )�@g*�C��c��4Pܚ�?>�
#/C���4�ۛ���k��unQ�FW;�N�p ]�}ӕ7��b5�S:E��v4|�;�;� �|��߼�~s:���e�&��_7��)�zнC�z��MV��_NH�TeU��P�y<إ>��f��Ż�@����,[	թ�J�
gkz������K׍G6�q�j��A�k,{�}Wu������;�&�/��VXt1�H�ۣ�W�?`@�a�t���ySZ���#�2��l�f�?&��)��n��&Ѭ������>Z~�$�)��~ghx�o�0${�7<��B����/���43��,':��v�Adt8�B�,�e}�4���,`��5���zrS�c�;���Rp�{-,r'��4�.�.�
��H��� �5��x9���2�[7�<�Ȼ��2_%����6�2z����N�r(vAZ���!�$d4�Ͳ��-�<��������mi�ZB�5!G;���7#
�Xս	>����u�!��լ�c�ċ��s��FW)���'�ݫ��ARI;#���9� ��$C�v�峌Z�!s�DgX��*��R�	U�)���T�������I��qS_R�����ǟЛk�U�Aúe75tBd���t���3�`�`;#;�y�;�a5k6tB�^qO��[ǲU��]R3Yx��Q�����C�cw�r�{s3��k�)l�^\z���ӤG�˕������0�c��5���ט�꼁��������{�I�yuz�k�m�jml�V]��R�>��¨|�|��+�ߔ�>��)I�ߣd���k�u��5�&�S[,�E�H7���|�<'/r3Pj�����d�7H���Р��N�o$f@@�Ƹt��`��U�����ٛ�5;n!�םP�T���)�t9�n���Cl��;��`�҃��T�rP�����4���o[JCf�66�t���,%x��<�W(��(,hj4�;�5�|}�q��=�1��X��߇)c�|Vv~��ܨ�\��;�N8�T�z�O1��XI{:k���3���������A�`~e>`�8�Mյ#YW��V�X��R� ��q2����K�Gc5�^��m}�,.$Ad���
���3��h#c�D���(^�0M�)�_e&h�����mC��N�"�*��:i�S�g`Yz�W��'������7���T'�f\3d�4��ED�±�m��ۻ%�9�k�z#ب�ht}C�����h���c;P��lð�n����it���È���x�3`�
��<���'[N�S�u�̽���-�!H�Y]�,C�Z�V��F�ֳ��H1޹Y�����"�_��¤ȟO��ѤD�2�ܪɴ�7�_��՞�}hVcD*�U�]�Pƺ�B/4t�}�S��9����@co{J �T8-��Ӊ�.��mn(;y�n�P����k�����<��3y�1Fq�L���5!X�a������U��7L2�<([����d�9m��t��Y�q��E˼Ī���-�Zƾ�
x�|yܯ+�T��Ɇ���HZ�]��~P�nP|Ʈ�Ct�7M[Y�"�dl��)���?G	�,J�0�Qꆱ}��mZ�Z��"_1e�0P{�_�i�z�� jMϜ�������כ�%A�[�/#�ն�m�-��׉�UO�s�P&���#*�=z��A��D�c�����}^&�+�xF�ɐ8�T����n{�)�J�8k۸޾l;0q<��ch:� �24��G���M�`��m��+pg�Mwii�MK�1��0^#��
ͽ�6c��[4��iݴ�Yݽ�"��+ݮ�چ�P��}J�a�iܧ��W$�T\R��;_���W|�0GMK�;�mt�L/e�7�-���:TfS������A�k=�=$ȶ�4}�SQ�c(�RJ���M��Y5�l띚O�c��/�3诜�C=�R�W�w.�̩�L���I�|������ۤNŵ��k����_��
+��kSfȵ�u���e{s����3y��/c��
��oo/�I<Q3%?�zd]��g����G�D�4���Y0l4���[°V�k����v��9C�s>�ڿ�PwN���]4-�~�Vv�5��_�-�̠(�gyyW�M�uN ��=7��h�������Xe��e�U����0��b6���J�0# <+4#gؕ� Ͱ�9����$�$u����f�۰#���4�N7|�)�m�^�Y�>����9�^Y@m��mr0��M0�K\��^KVN��:���c��A��t�.{�7�ޢ]���;�C��vٕ�3f�����l�Kۖ�,��n!c�Q�v��л=�tB�㙫�]����HY\�SJ;���z�E�9�)���[Nыn��6��2�' :�����絲P+�%�#*���Qy�T��Z�d��n�Ϯ�9˳��P���Q��Az8_���<��R�����XI�O��)m�o8:���c�y��%e�NP=7:��VԻBrY\�k�uC]�V�O�N��˓w��VT~�җ⸒���!���`6�ճ��j�NR;Y�8V
}P5|]�
]�]&9\2=�;�2��ok��}EKv7���L�����Cs��a�o0U#���驪y{�����mәϗ�H# :��(�T�sǇt���q���}�m���s;$fړ�d�A21�����`a�{�H��V�#�]�De����9�Ü8\*�G�J�Z�_;!n�����o;�|h ����d���#r�����)�������0q�� !�����E�^4�r����rg��J��u^�J��)����=&�)����Oc��m��
`8K���}zb���]L{ܺ�D�B����#ь�ۥ����A�	�~�vC�%�����(�9Km�p�a�IG9�{�<��p�d���:�sG�*gW���Ԥ����l��P�;N=��oK�T����ys��G���3�b0_G�m��"��[4]���Ý�~Ź�!o"'��Z�,��NsCX1
=˪.A��3]U�.�������F����V��sjf��j�$�=c5���1��;����W!'-��$�����˱�SL���.�f
���ά�E�-vִ���x4�â�a:�p��H�wfUժw���fu����+��W����AQ�5J�c/���v\v$:�� �VD��+)N�u=,�cCC^�H6��<�f���Q6�FE��++��>Ԛv�����*D1T@�e����ϳX�kS@�r �
��v1t�s���=DɆ�9�pn�ڷ�bzU�Y�:i�M1���\�H@���[:�$�P�X��-P�l`�ͭ��k��*��NI�|�ޑ�n��#�-�H\�
+G(N��U|o*�bZ/;8m�#r7z�ΑV��K���j�9���t������Mzq�Y���sY���	E�K��*��W�J�}���0��	�����ƅ�/�����c��q��=^�J�N.�R�B]�y��`ڲD�M�XЭf�GS �C	v��j��J�ٛ=uC�r�k��*݅3��g���,���Q���za,��,�	�z^�`Odn��)�4��YT"98� �bzXa]㾾�S��C3pY��kNF�k�:�;��n���#�/��a{N/41

�c�y&�^��P���Ix�F]��"V��������m�v�+z5��,�јލ�Kl�;r�ņL� {*�6v���wfvWt��B�YCU%e���z!���w��(�Hbkp+�,*�7�t����wӡ3��Ii���#��Qq�0q�[�����[�����5	�OH��z'�e���#�
�0 ����J�D
�����&2��^����L�ll�h����bm�}�,�ewk�"�OS<�]�(63,T!rD��Y"`WJ��'[y��f�L�ZWh\�����f��z�>!�w:�FզS�l]��Ts:ձ*Pv��z��	6�R��2�j�ؖya��1��+♖��L�;�\��^��p)2���F����|��$�5�+�9���qe��Yt�L�cc������k�9���m�XeIf�\�eSZ&}���a���R�ɮ��R���p����vtvfE�aB�-��õ�e�4��h����k�vY|�����)�Wr.J�L\�}���ik@pޕ93��8�+��]�G����ݹbM�o����g�d,hҫ��m,W!�X�K�N�MN��;��&գQ�0�� (�3D6�jv�}���CE
���r�z}��w	���1���YPd}��j��u:��xgV	ikW�U�n;��t�TC��*&^��\�3�\.u7�ЬU6̨>?�=�f7�!T.ns�
/�:�ٚ655J�<����PB�ݼ��}��bsv0�uC��ެa]A��@,LޞRV�λ*�C&nm�^����$+�v�>�9�����*oCvޘk�kgF��p���Id��c�t�:�^<؄T^bK�[OZ̓,�bԩ;�������ݷDԿ�:L>��*h���Z)=CU�k�\�c��\��H�j��T����;� ܝ�*ۥVj1 �<���ARWY�j1
<�;�BM�cfl׼s;V�w����i�ζz}��q	#tuWd�q:��U�-���T9Vu���ڝ��PњDU��ɻ�	�_4�Мk��n���V��*�r����]$D�����,��_;�z�Z.5�r��쓶X{��or]L8�@�%�"�e�T�;����S�3���'!�=9 r�Y{*�ܳ��Lʄb
?=]�u���.�����	kuU�&�;N���B�5yj�G��ܲL�Ǆ�A�5�e�֛��aPe��4�f�Qu����T�F1V��$ٵ�����et��䚷���^w�S�����5
�f>��m�B���k9W�6npoRku܍N�rT��r�.���J��~Uy�����N��뵺!Ǳ�&��q���)�R�U�}N���ݻt�S�9�$�H��3"�i��C�3�E�Ƞ�.��ˊJJ��N� ��;{{~���%p���N�^����Ü(H��r=I�ɔí���z�| wR�(I+r�ǆ��Sx�nM�e�4�����E8�.�-ڨ�Q����q��Ƿ����>x�y�I�;���-Xz�:�}��A�B��\؜H,՝�z��{��ۃ��"�I���P*�ɼw<��&PS��j%e�ȃ֓e�8N�"�(Ts<��4U�7��z��)VPQ�MV�4�q ��\��Ӕk)"��EBw�Dy�y���4�3�M4Z(4�ʣ�TZ���Q�
�n���p�$�W�抖eU�В˘$kI"�_�ǲ!�(s�U��e[)bA���r�*���E7c4Qi'"#��
.�
V\({HNM��h���+аC=0cj���%�>7����2�]�M	"�P�q���*�qݔG� ۗ�ֈ�G�Z{6�d��<��o0Rk��K"�t8���'�6F�St{|�9��a� �
泹W�oi埧���v M=f�7��vn��\����G���h=��`F�_;��*�v1���ٶv�17=`�#1�^��W"}ź�q��Oi�<�75[�KXy
����f6l����:U���ז�3{��Iva<`��k8bg�`�ʥ�c�Ο��B�;�̦F�Д=r��W]cw ^"z�O+"t�h�N�*��F߶�Q��������ƇP*@{�53>ˊZ��:�	�|���ơ�������g���`����u#e����=G	ŉTdg�[Q�6��$n;��<&�^n�)b^��B쓷u��[ n�M�!�3f���N�m�nc�v�+�5�~!Qtw��N���r�(T��A�݃"�Z��ˇ�ӛ���D���Ѣ+J��IYxF�[&x�M��t6B�/���pT�Y"��M�6A�z�W[�S��{��X�V)��S5]��$+Y�K�sdYG��=�Y^����MS���^qH]tx7^�w��K�֝�l�×2��Ֆ�r�pl5����7�w���©i�7+���ٶ��
�RE�]� P��Bx*�ì�{vy+E�a�T���C���Á�,+�:��U3�y�l���AF�շ��c�SA��:h��if�i$7
|��t���{P�� ��6Ϧ}�}S�,���T�3����ϟ�j�H�g:�h�4��\�iy	nϕ�2·��s�4��1�?��}�z��y��;�0�+K�ҮEm)�D+`E�R}�� G?��P�7j���0nbw޶�=����Aa�NV�n�{�/}�:A��ҙ����F�8��-����C���,D����,���=���~�黰>Ϝ�����s�v���:������}��A	@x6j7�]F��$��h�|X*�Ŷ;�ȭ�h�j����?��WZ#�y-W�s�U��0k�s*�9F2M����Z���%�%Xا3�p,t ��T�zg����i��ۻ"[�C=Ӵ�y	z|#��T�ևϥn5钨���G�]�K�mgd9ߘA
��r�<]5�z����9׫�2�y
eK�	j����P�-ї��0ʾ�٭�zv�^��Cs��!rH�� XӋ%72��1�;Z�49K��y���7z���1*&�w��>l+�"=�7ey���:n/w_�����H�O�mM�-��(��2�Z�q{4�z��mJ����\gr
�rAM(�㶏U��9��<�8oUʫ����,x�B��T���F�Pe*	)T��;V#��1�t����/������p��T�����d����*M΋w�|��W��S�Tq���n�sp�9�p�t�y�(��9�zRNWTֈY�b�z�}Ļu/]b��g��u�d�x��N��^����ι�E��z��1��Z���v�"k����.4�[-���=������a���F�})����ǰT�p�Þh�/+��#�du�������۟����:�W�����6f��kvX~/������]�OrJ�銒�����i��\d�Q�0q�ow�?W����)��zw֭�����V֮�:K����J;���I�ܕ໸�h��J�/��N&�*{�E�7aw���<j�yլ�CT{&�N�r�c?:hP���L�f��������2��G�����N�#I�:Wg�����b��o��R�S9�l��u'��b�-)q�>���^�{׹����2�0�/2��#��[�����=A�ʝoX���Ȧ��Җ���h�㑒�O�/Xw��}ρ;:��\�Ky��E�͗g4���>݂'Kj�<��2:�ǲ�1�}xI�b�Zew~�%���c���gh�u^Z��G�u�r�U��ng����7�[|��I��E�i��T ��*f��f\v$�A.��7(�V�37ǲf�)�-%MQ���C`�L±}��ȹ�䲻&�v�:4�y�fzụ����a�b@}�Zlv@� w!eω�-�rW�$_*����UDYm��|c�h٪>yU �3�^%����},.a!�#mn��9�N�����0�1�TI���S�n�vd�I�k��&ӻKtH���\�hhB�`a�F��E[t�	q��[!�S>_f�^���i�r��0/��Ҙ,��y�F7A*��}�&�3_^m�r�v�ڬ���InH�4�s4ӑL�6I�Ǵ��֗h\�U�1,�m��֦�}ǔ��!ܖd����|�fǔA��cr��\K0h����M���Yo,�Jw�v�~�dc�<MmE��`��w��;��oIT5J�5y�OO{�[�m�'m@�5�{��L,a��.�%zq������J���vd�9���t���Hl��+Z�����\��GTҡ�ٞaum��j����P歙z��*8�f�K׼a�[/w�5�%ӓګ8ҧJ�[3m[tgm�<��!�m=Y��B���=MѾo�$7�Ĩ�
��s�Ρ�T��LVaGs����.�������6h`��[2�h`����wmF-���vS|�_k����z���S�ud��^��A���T�tSϴ}�OA���dV.�׋7��`��� ����c/U�9�e��n����^��T(ZǤ��u^Y�ݑ�Ą_c�>����wzcY�-����m=-I��F)�a��BMw!���b+C[�3ܰ#�c=wc���cY#6�G��S-�>!���x���[>E��ZF���v��ڷ���ܧ��O�jx��Lm�svk�o��������[�a����u�^��/��5\��=ܭ��橴�A�Kgk�E�q�N��s��Y�����x�
To�Ǻ�E��74�vY��;PF_���X�����kyhh���tC����7�K.K{��U��4�E[:�d����a���d#-#���ZwhnAO��4O%P������+MNUvE�;i�{�tJ��r��\�q�wJJ��זɞ<U��*MW9��}������@�T�]��ࢸ)8�=�'W)E&�QL�+m��ٝ}�n��3��2m�0�@���5l������.���5N�z�mŽ-��'��[�����a]����lÕ"7���\�׸����������wtO��<��mv�Lی�o{y��롁�\��������	�������J��[EQBS��s��g|�vD<ǟO�R�W�Nz�G� !���3$nu*�r�[���u=s>�ڿ�P~?�-G�E���|_�|�w�b���w����vC�C�ڱvXy����aN��sJ�ie�~���݁�/w����ڮ}�G�N��{�0�q*��lU���ؒ{ُO)뮓!�_N�ko)g�u5Ou���	d�l����ZW�uu��3dw�<@(��3=�Of�8p�f�a����,�T�A�;��x<���4zfS������`;O���땕]w.7���� `&³O���6/�ƒA���y���M
���=m3��J�4yh���N�ڼC����t�Q����}�g��3S�N����%�H�VJ��s d��y)������;�F��纶�jC)$k�M�@i(7��:M�A�>͵t)����5��D�)�$ٻ�A�5!���;����
�$��t��mQ�ɹ�"���!Mz1�.���vÌ�0B��B5j�=����@�0�y%*��' piɧc��뷈����j�O��=C�[�n�e�>"}���k�Y`ggY���˘�[9�6�fgip�׵%T��s#k��2�!�(��9�cET���%�['v��O7z��Cl�����@lǁ��.��4�����mצ����ڛc�s�v0'�Yb�l��:�V���|幋1�Trs����teS���o���J�=��|�M{Ҡqc���lrɍ1�f1I�vV�n)ʬn��*���]��d��mk�or���<-Fe3��Õ��Q��&(����U[��7>��|[z��⢂���9��岧��ޱ�����n�vu2��������&�����ѻ�\v3��22���w����]���bQ{��j.�rjb�hO8
��6gM�F���W�w(��jF8��'Y<��;9چ<M0�cT�=�zw֯�eu1Ք9wU���5�j�j^�E4<��ܵ��8ޠ�u1�a��E�:4#Yl���D�l���م^Nr�7����_�=�M��a�X3Vo�%j�����b�#Em�0'hRa��^�I�~uS��y��*���i0_/ �WCu���|�WB�j;�kޔ���K���U�1%zU�F���^��졊�\�0�iM�[������0���eW�,�C���%Y������Je�,��R��w���8 �-�(P�ꧨD���k��� ύ�='��`�͛��Q�@�֫��εE�W�k8�eu!R���~᭺4�E[�U鎯n:�n�7p��K��ͣ�3i)��emU�����+�&�t�̏vݫ�P[��nuD�֦fg��xL�3��F�26wK�ղ�S��F&rň @w�e�/�@�!_�;ѽ0��mq�L��$_5��UG�'�4�MH�\�B+[�*�\���ݠ��o�;��#�w/	RIO�� ��[��;2="����)�F�H�t볙�����9�I�H���3��ml������K^ol[�dw��k��1����xP�e��������Y�R��K������K�����_V��zy��y�0��-��t�W��*������wWGpbb�a���n�1P6���`����;�ӽ�͞����KV��Y����t��d�A^�K�[�����x���4�8g���j7��<7��7�����u+�l�:����9���k?���t�B�e�BZ���px'�(�đ�2���z6@�v���č�Yc2�"}�]��L���W;Sm��kG�^��¤���$�*��W�8PyCo5��b�޼���@��Q*�L�1�J]]��9���m:�\t8�F�n���n�MjW)��9rMKMr�w�imf�ɌR������i���Wd_\}��rpr�.ä4�2;�^6Ej�C��#��1�*y��nc�2���<Y�/1e�����#o����0,���;x^[����"Gi�ઃ�7m��*�oS�����i�Og8������+'�w ^"}�z����!�,�p�U� �Ͼ0^�Nt�C��}�Ws�#�,��W�T�_%�sN��Z� o&�%��gۊ�m��GS>�qA~����XhYG�<w9��s����S��n��4�*���f��zˊ��z-�׃}B��jз����ӏ�.�GA<�B*�W���\�vjf�ʁ���l��4�d�R�#�ʸ��{�%�/
�mD���q�m�\�i��V�jj�(\��p�~KhO�GYxݞK��!�:�!u���V4i���#K6���z�|ɷ�!��c�ܽ�5e0��K%F�jڷ5*H=Y��M�W� �X(.yKj�����n[����M���&c����Q���H�Լ,u͸	�u�sh���	�k+�gQw%n�Z��\�[ʜ�-ec-PdWvr�Ed���o��Zܸ���z�����^��1{c��%,dk��x��*�KT�ٶ3��;P��R�T�$�>��&^e�
�ݘ��6^@K+sk��Kw21�H(�X�侫���p�;kS��7U�i���e�]�(����v�+iv��ԃ2Fuު��0%��I��wQ�;�;���h�������]���AfOE��teIe���K�+O�I"�_Փ`��PX����F�a����D�����j�������l�e�43*�!�y�a�E�Һ_'�˾omau*lG�+��8�6�5c����b�*Q���<׽�/	B��#,��ީ�/瞣C*n\j�za��Gx�ڳ|e ����ۛ���')\�4fKp�f���d%�U��,U�+�
v.k{�kA����j���X7�bj��v�8�@sjܳO@b@5��)���cb�ԸkK�N˛jD�77�!/B�N�_'JP�B���Kޭ�,fG�.`�$sM�}j�&�����7[k���nM6���[Y�R�F�U53��s�-��-�fTA&3nƮ�� ��Y�K)[�7�0���V2�q�����W���w��T�i�Q��h���`��*�7���5�=�a��Wc Y�v^����V�KA2����` E��qv+�Ln}�C���B��FA�M[��	��nF����gyH���(�&>,��Q2����dB���\ʀ�0�Xx�����&�D�'���5�b�%2�]�̆�B醊n�32vr]pC�,ڷeC��
1F�7�����r�3u��-�Bn�솛ݐht�-��JH��Q�ӥ�[�勳�cLJ�L��K�p��pW�luI�]�b�0_U�s���XĞ�mjZ[W.�.��̮�`�nJ�|��5�u4�94�Q�o;^[x��} �Ê����n�nv0]@���e.����5̮t�9.x���>�o�eL�����n�U��3d���<(��]A��C�����驔�<��53�N��I�m�v���J���S���Ækz����$9�˳�zNƃz�wuU�=c����WS[rt�E�>Q�t�%-��H&P���|*�m��}v�Z�5�:л_�-���z�c�8c+���6��(���S���r���P��:��G郤K�� V,[Ko7u�tb���o�/�eX)�p�%���5�8����VHҝ�7�N��YY(N���6����S3�]|�i��n�����m�':�*at�����t0��v7/ A���y�ݑwH&�9ܬ@U�N\g�f��Jo�o*�O2i.�Jr�FI$�IF�\Ȥ[�����JV�?�lR��*i�Ӥo�}���ܙIDB���r�$h��{��ff�2�e4���� ��+�v����oa�����9EU��X��a�q"���9�C3QV��YbŻy��{��e}�1:E�$4Ҹ� ���,Zm�#J���J+zw�Ԛ�i������vP��JHB�ҫ6\zMȂ{|��D8D*�,�;*�fgn=�����n��V�SA�h�n:�E�#"�#$H"
4ҤD�r�!2�T�PDq��&��u��RF�*���l��\3 �����JMSP���g-���$�
�W/���P�%b'6! Ql����u�W�Z��;��(���Z2��.�G�s�9���.r�wnq׎!8qL�NS+4�HUr�����rr�*��H�Ζ��U:EȊ���UT�E�k�*�,��@��-#wn�;�Th$R\A>P�|��y�M_��+v�J�'o^r52ow�b5���Z��[�׏6�e`�y�ӬRC��v�m�KP���J"�$�X[F(Cqô<x��vsÏh!����G���"gQnF/��WC��k�ܫWYqOEƇ�������;�RH�{�kba�ݟ\e�{q�7��1�upx0�q��a�zngv���b�-�Nz��9�;I�}��ղK9��{�����"���{!�7�r�[�����@:�\�m~�'��G�E��nӄ���]&э@�a��rB��-���=;͵��Zħ���sv��a�e ��+$m�d;�"Ϋ�-���8qW���Fag系��Mk�	�}ʐF�{Z�b��!�t+�?$�t�Q���=U�!�Mii���1���9�u�H�Z�U��s+i�����mn�1�y�K8��feM���SrBz�$�:8ٴ�]2�h�P׽[t3n���[O8R��7y��tE�I�P䂐)Dsq�TL�3�?8����K̼�����ɖ��f�v���+�8�R��'b�b©X�@w$ݔ{���"j�ߡ����e9+�����c[w���,V��)�4r��+l˨K��ӌN�6�3���:Y�A3(�P���J�`$�o�k�\J�Dq�^�z�iХSn��\��ө�nk�Uq��%*u�p��qI�m�����I�j�U��V� �NEL"��p�|�F�>H�e�p�d�ϙ�A{���,�suا�H��>�{��H����HG�B����F[����FT��h��@�V����cĶ��:�	�!�۠��y����Jb���v���:��z�Z��%8^�1l�f�vB��y�q(�[6i߬�ڞ��Ƕ��c����=W�g�lH���	wJ�z.��~(��ۺ��.m�R�7���ʲ���7}���y؍X#�0n�w%ޫ]�%+��[uC�{gJvNNkq�[;��_o�/,�#�$z;.��j婎���4�B��6�,�3���Y���~`������F7���Mܦ;(38����4�����*�Ż'�t��g�1���Lp�_����jb�}�.5�u������]0�".k�mn�@����w�����u���=�Y[�W˭�oI p�L��Z��U[��+�)�O5��wGz��uwOrJ2丗'eѣ�θ��I������;KyZ
�jU�F��4�+�Y1��8���}��"��A����b_���S��޷��� �=Lc׌%�
;�Ӵ?[�jY�^o3_e]���-�xs�"$i$HH�u�Yj�E����mX�My3&��n�dd
��y�&j�.<���~ �tс�z2�\�7ϧ����V�zY�a=��ꧪ&�>=X\�UE����h]�$��y\�.����ĭkO��G�3�
���qby܈8�@F.�/�9��0TK���Mм=�h���}'U�9��/@4���G�s��Ѱ����䆫�}YޯtR�k�T�R�6Rۧ\fD��|h'�R�݇�o:��[�Oc�#զl$y�)7I��m���N_+�����_`9�K��ݯ�26�C����a~�+ �+������ޚ�̨�r����y��gh��a/���t�Eq��䪎~���7���og��C�-v��Z�%�Tƽ�1��u����i(�����s w�s:�'޹��H����X�⎗lO;Sy*�� F)�{���Ș���.ۙ{�w�h�mZ�M��Y��X�gb�L��}� �la]��8�(�pŗ�ʥ�f[C�pw3k�U�^0�q��p�ս^ْ�6l�N�l��m����,�sI��(Jݐo`t��a$fǘk��]9=�,��E�`X2��b�14N�.�� 5?6e�g^��uB�жF��n�N�b7��ʨ�N.�7csWX{�s�y)�n�E�>��A�WDI�ٴ���zı-@xVk$j�x� ���^d�����K㔸��t��e�9�7X����z���]�ti�ѽ��lw��x7}�/�<� ��%���κ�ac���X��P��H�΂�B���&�F댗	��?.ٍx����Qs�t���0��$�M>����<6�w �UA�3']�U��X�O@�yZ	.�y��܎�AR�!.���D�ѭ.�M|�c3"S����n�$��nws���(�׷�Tַ}*�f�]M9��[zdT_~o�ݼȫ>̮w�d֪���!K�y�,�ͭZȆ�a(�%�g�"xG��z[飮D|b�𑵋���u�$���Tې�k6[=wN��su��B�t�W_r��bsn�f��Z�[ab8�8��J�s�`����Q�%��$���9��E���3BS���P!ɑ�3�e��ݝ�&�-�ߧ�."�=���:a'��ESmV�7L^:i��Z=�/��&���<2D%����#�RV^[�z)���C�����1I:���u:��8T:+k��@�
YxݞJU.0ʝt���]+����[��c=/e��{��C&�aN����w����1����6\؍���'����ȑ�G@V�25�Fc��Wyey�k'�-�=�V��4�hC	ʠJ14��A;�mt��Gp��i���M�\�T�-c���rå�L�fOW��O���o%�Q5)��������~�)=P���ӷܡ��lc�`�T����5삺������9�-z	�ͅw�Ro8�TԌ�w:2�I�·3��>��6�g_#��VM��ڳ�ųC+�cu4a;
|�Q�:�8�b;�2<��F�U�6�̴sR:z�V�?��	�0kЯe�+�W�:�v�T��;��b�u5��	>��l|�߆x���m��Q՘��5�Lʻg}:�Q�R�����-�j�+v�k��4��(�m��54U"�q#�`����9k8�vj\I��X]I�(^��%t�_`� j���t�`w,W"+�jhUXxJ-��4^iv���Y��"$f��+�r-��;�@���0��2ek(D㆘{�Kch�-Vn�2�P܋��xG��$�T9i���L�C�d��/C��3.$���{������ɋ%��B�W$'�9Ju����Od�B�F����]Dl�����#j*����<#ǗD��l�U�R�KSȖ����x�y���촨̅�s�ndU��p���EH�"�tL\��k穻��M�m����U޳�aTh$US�Ǻ���@"����};q��G��K6XZ��b�=�%+�\F�{���F�ÆCf<m�Aj4�9��`�]>�k*��`
��e�ս��+ܩrw�5d�;gӸ����r�c��T��9�څ�rH��ޞ�|g�lm�R]7�%�l�u�hX)w����Ks 8��e��ß�^�׷��{����_C�K������^'V\�P��l��f���P�㋟]�ϻ%0uu��m������GT��e�L����-�[Rch�~+sC����\n�c{H6�e����C-h�W��|�X:���zs�F���F��t��K�k4�nV�;��5�4�;�]!fGI���!�7�$l�ɽ4��]t�4�g��﹞w�s6�Փڪ�l��6�lo�|��<��ףYj�-7�ʋ�{��w>������*�7d�1�ў��:�h���,��S�0�o
��wOo��N��D���]m�8H�m28���Fz��D��U�3�x��A�n���xޟ>գ{�</,����)N�{�Z=7E���;u\t�ddZ�bh؄+�5uY�+	޼0�ʲ$���3�j2r5�k�1&Y��h���,	S�OW�l��Յ�fgv[���8z�'0�&7,Ur�Ӷ��xs^��+�b��Z=1�u�u�����w�������丢d�UG�'JO�P�{����w�������+s��ߛS��S�P�����V]z�!�:��Ɠr��k�<�����d�`��3u��*� �v�>cVL���>zgMuu�+8\��r��V2�x�����,�w8KZP�t�oq�r��]^m�0��݂؀�|�>磵��o����MX#�vu�J�]zY$��/��r�H�Ò;���4��rYֶwt
@N�R#FǫB[ћ�:EX��5��m���iT���D��/�L7�З[�C :="��}I𾎹�c�������a����l�x�0��y�p0�OHa�K���!t
�=|�����͚ƞg)5ս헝��/RF�<�;��a�,�>���Al9h!-�2rߝ��g1כG��ʭw�+vA��������ކ�]��Uy���n��/���Th:W:ue=�R�+�l���q�+�j�Xh���ieEa�rnû
Ӱ2�՚�)�+j���;��^�3J��T^���8u	�P*�x�8f3x�5�1���uϸ�m���Ϣ�c���諧�j��v��Y�ʴwF��{;�?�>s	]���Cs�_c�vA3�a�RN�r�	��́�.؏bθ���DVk_b7&��m���H�Ӻd����:��/��d��,X�m���2Q+;BĽ]q��g^���+wke�k���
�N;�g�ACq�D�܉7��F>�DSl�vU�L��¤8�m�����<����bk.���W]{�5U����2���nk8�H]�?{�᧓h��#��=:�^ �܂W绒Ê[8�15��9��Z�\������g�)�w�IM��,��9�������U��Ok9���jC�'Ѐ��U���H�d��n榜�o�S���k�u�m�H݁�n_P�XD�.���i�h�J��G�By����x���7Lbi�
��0�W+k�t$�:3����ܰe{��8�;�;�I*��t�ә<½D�Em	ࢸ.��=j..�s(�s:�����CM<ڎ��W�d��g�����
�G�A�pT��|Qg���ޝ���G���1s��sW�zL�����Ӭ��E�ߴ,���"�^����l��'�ub��]G����6���|{*㣓˖Y���~=f���=��������Rz��\D��_cճ���|�ѫ���<��oug4q:�Wx���|�O^���3*�<�/Z.Zݜ��e�8��U��kj�%���bw^�˸��|�m���A$��:��M���gWl��O^v��ʰ�"��C�vgUxGJ���w��QR��mB��ءb:��c��x�,��q��ٟ6����n�a��F�^=�������;��e��z���`{�8���`;m�!f���w���͵�s/s��w�C�+D������=�h3�]���xVj7�������c�p�9<�73!� �cN��Fv)�FC?�wB�-�ժ��8t�l�3V�y�|�ml�ѱ��]!�Ǩ�r-���b��1ʉM<"�U^�߲A��y��9��]�����Tʕ[�ӕ��ց�M�$�K|u�{��P��Vmky��ww����φ���
�N�&��$.>+�
iG]ӝv��pѥ�1��zj��y \��Lު�b�K����a��3�m�Bf&�Q�<M;�U��M���V�E[/D��������~f�zt��:������U-t��50���M���K�ݔ��[��7.*�g�̔gN|��;ϛ��{i��v���'��ی���t�}.��YH�'�/{��Ξ|㫽S�Fԭ����o	��ݽ:����_�as���6�Ƞ��Zx�jpaM���-qThb[�:����U�\�ܧN[�r��z�={.��آmò��oQ˫�]�+���ȯ�t����ڸ�[B�P���'{8������[� -�UŔ�2���*��G�a�^�,T�tU��u�o:ʹҺ�YN�6ĕ�y���~��(�&%BD.r�5c�v�!	4je>�7�a�WW�;]v��J�tև�c���4\��a��w[0%r�F:I���j4���^���Y�%�/Ƭ��.ɂ�=И�O8���KFd���lx/�>��J����T%>UEL�'�Xtf�mݪV� ���S,��Y�qXZ٢(�PʝT+j�w!�E�a
�U�����k0�e
|����{sz�(��TǷPe7#X���uw&�� �$]�S��Cq �L��]W�l��з��7.������tn���o�8�˻f��I�w���|˝x��a�����]XA^��26���n�&�4g1�.���r��o�5��9�|�_R2�B�[׽E�Z�͊Wc$�wo���J�5r�a���$.������$�������X�����C7(T�d�n�o�s֨}\�yu�Yx��a�8�ҕ6�A�#����e񭉈�5=�]��ט���;��ꁱS�&�c���̽kR`�HƋj��2��V��c�e
�.�M�Ӻ�|�*ۼKsB�Wl��#7��5#���ބM�Q�Zf'�����v��%���+�2#mj]�� �v�9X��Df;�)˱��:�'���ȝ%쵹�'�m-�J�{�=����e#���̀1|��t��j��cj�;�xJl;}�esW�+[�j	E�0!V\��rhhre�T/D�����ö�dv�w��vr�NT�4�J�O��|��/��e�d�d�
�i�	���ɷ���'��w:����(N��E����I%.ݠNY�C��k�	�;���jL��n���C�*$Ŵ)�}7��Vj�E&k�oL�TX.�n���W.R2����aJ��i]3�7zK#j�G ��p�ws�l��Y�<�S�a�sM�����Ո�ns�ӎ��gq�i��%SF��K�t ��[���B9��"uZ�O\w:[�y�Ldܙ{.YMa�(K�K����_6�#z���nc�Z�[j5F���5O��=�����G�g�9HP���>���v<�u ̦��T��v�Wqhz�Q��Lܭ
q���Z3��yl��v�Yڇ��(f
y�A>k�gSvr�ŏ�UtK򦅂TbQ}$�I&�dΒL�@��0#�G�BZ���⑩z$QE�S$��QR��TD�4�������z�T�jbt
�J�!3*�Q$�� �֎���I�{����{dI�'*
D5.T��w$"���fa��"�^�Z7�UCj�N������A�]�����,�AȊ"���\�L��
*�E_m�ih$�(�����{���q>���(�I��]M�B-����9r�iagB��10�H�H�0"��̈"����B���\���̊
�XA#�49˅��#��"�]ny���r����B�Q��J"
t�W +�x���!\>]�9{���rN Ez��̣*"�jQȢ��H�UG""�Nr1R�9H�)��&�(�� �
Nqg��5B��)�I��*+P���"��ĔWR�Y���z����{�g�����l=��X��^p����Q��wQ��x�{��I���
�Y�Еy)E�ʗS~E����ْm�&lu9����2�W�;�����T���˭;�E�ϒЭ��({~y��m��(��-���xҒ�uƛg��]D�6cힼTy�y��WPk {|{>{���A��[
v�֒�@�K���#�5�}�)���3T1iٺ���h�fO�]S08�*X(oA��oOU�6�$QH�y.��̮��UG�v}�N�����ᨌӕ�1x� ��j��F��u]�b�s���z�Ѓ�<:z��S*q�6�>y��#z����M�kMD��=�4z�'N`\�?�BH���4�����=��0a]�7b.�,;j��Ζ�l����B�<��rn��'h�Pc�g��f��C8wö+5��p׼@�G��wk3�1�w�L�<�D��6C+�1.m�����b6��'X��=B6����"4��Zt���m�q�YY�>�b�k�TF)%]�`W:Y�5��d,�as�(�Ӎ���RB�E��c�N�y{g§�D��*�[��\{^Be09�.i�"��.N�q����^�sH˸�d�+��*:����5b���E�S�1��WO\�t����
 y
0���oU�j���-<C���Ϊ��
��Y"++dj�3�q`�����"l�ȸT��M�[�Ck?[wv���z�c�4�FȢ����=2��0���,Af�B ��)��ё}���U�$#x�n!]Hȣ�k�uQ�駉�t
��J
���s��Е�+tF��d�����9�T-o�6[��Z7���>��*Ӭ�.��n��C+�EV�[ٮ�d���2�w���݂r�����&vj�(�S��# 9]"ح2�﫛�Uj��0�q1`�mS��UlN�mR����v�a.+%�.����P�J����p��m��b%�.�mg?�� Q�K��q�k�+��9�~���Z� (< ��R�G��w��yP��b�w�X?[��շ���9��?���=֖ľ�p��74�!��af:6`m�vC�xɯ_�Z�^�g���Xd���$��QǑ� ����A�9d̀�Y�Bd�t�٢t��80a�r�ڬ�X� )��=h��ܨ/���]M�\w+fU�`��>�^�޿�8���1�������Ͱh��W�bT�*ӊ���Jj���c@>`�6�h�;�;f�`�݁2�e��r+*R4t槬Ѳ;��b5��t�:��9�ok�W�`�!u���쐕�f
�ƿw������`7X݁������Y�a�d��M�9�p�}a�Q���lw�yn�Y�1Y�	>L1�᧦7*Gb���v����H�g@�ZRѳVv&�mK�B�!GK?]��&��&A�"}��M�yz��=���v�!��sU�ڌ��S�7"�4���*Tp%�)��-C��\��c���T;pos� Hހ���b5�ȁ�B��x�U�o��>�Dp�����>��!��1ܠ��3�\���vKz���]��:a�<�HT|�'�{�fʗ�=�/�K�j�i��<e���)�p"o�$�,����i��P8o&`�v��.���:��bz2��\�X�\V���Q!u4���-	o�z`��ɘG-��L��0޳��2��-�jm��<a��7%��Ws����z�mO*�1�m�CB4�f��8`{D�5"K:�wl�CfӜ�Rr�x�9׿������C]:��)�[�N�\[��x����u�m�a�y����H�n�6�dwWK�T�o8�d�J/�o<��z��nCT��&�d����h갑3��/�]�e
|}�Wy*J����������r@�+��Β�R�}��6�A�f�i�D{�&��7S0�Z��Q�����*|��ho%�
&��*=b���U��{f5�÷��_D���|�B`���Δ�an�m5�q�6C�u�z�8xPf��[�L\�u����C �>ٜ��wk73��޻
u8�O$��O;��!���z6}�+�uk��� `E����
�yJ�E�uUcn�Ϲ[+tu��3I"}Ō{N��Fv)�q��,���Tц"3Os�u�{!֬F\^�h�p*舜�=Ib�E��t�lS�y>��#�h��o������b��ƆHbW��W>�6m���ޡw/�귂����t���퍛�J41��"ٽ.��v����A}!J<Dy�jE�\��oo1֨I��SOO�]��I��/�uԫ_��?��!��Hޮ��xf����S�2?T���}�Н�0Й�;�X$'�>&Ѥ�w�k`�|�Bk[Wj��}�Sv�H���-w�4"�$.!erA4ۋ~�e����Hjڒs�P]y74�S�"�?]�<#V�o8����l���h3��AT-/�U䔪S� �\�SS�x�_�ȧE�x}��]��0:j�������h1{��~&�<�*�EO>�\��. k$ɤ[��Uu��9|��3z�����xҒ�\H5��f���'�a�v��7��n꯹�]�aC�����l)�G�7�TW*\�2���|����ɽ��4�[h=���m���zؘ[����f7���oZ؟QH�Z�J�DNk]��k�����ǂ�e��f�̸���h�0n����u>�=b_0�f����� IPjFH�`��7��#z��3"����p�:�:����}"to�5�^�*�`��,7d�ތ��-��m�{s����V�Ɛ�nU���]et�V����Q�i�#�kS�T���[�����`�u�sP4�6�벺(:]�z!=VO+�wԦ�5gM�ٮˉ��õ����j�����_� e���w���"�{/�k������j'�HN6ݥ��(�1�\��@�v}��1��Xy������6B��k8wP��SP��z�w��5�Ϡ���<y��Ye�9s]��yTGnݞ6�M�a�'"�<rכDf8</$��o'�xp~�ޭ�uT��9)C{|��3�#�}������ѡ3WU�k	\��1#���^�Y��;�(ٟ_
�9�nl�8e�	g��y��Ũ'�v̖g)k���#�� ��A�*M WcH=P=Q.g?�Wa�)^�,���9��ާ�7��gt� �
��M"�I�:��fW��V�*�NJ��X؜f��p�t�R�9��	-���)+�xF��S��W�-rc��"j�N�ec��T>����R.�"��!@��V�f�F�ΑC���ی`Vܵ6U7S�Mk[�l�lT�(��wůX/�,{��c<Um����P�ul�l]2zo8,��{�h{�v�]P-}�&����
X듵;c|�6�wM�SWmn���TM�;���(z�Qcm��0tn����y#��yS.^f9ټ��}	�h��j�7�]*!~) �Os���+{���ź	5�9�U~����a�W�.�.�#kL,���*=�*� �����m��v�z�!�2�������ᄺd��D.�W�)���(����n��[gwDѤh%�#2����6@a�,�ս�3�`37���q��Nދ�9戋Λ��<����t���`��`Fn154!����[�9U�VU�hA�wH�]��WyҶ��Օ�z�.�-0�=M�(�ck�C2��4s�����8�v���75�Ƽu"E樽��ݽVY�`�~i��Ӓ����EMK�ն�x �X2�x��!+�̭\hq�l���}Dd�m�\��MAȃ�o�]I�p���P����î�x��t�c%X��F[�j�����5�"	�"F�D�惂�^_����IV�yOY9�F
ޱ}���cR���B$u��VD�<�}{j}�Oa��r���)ţ4�h~�=VU�-���D��ku��=\�*��A�`���Տ�~yޱ�W�F�|A��Wh3����a,1I���&�:1B�pQz	�2�-�j���ԋ��ݸ��$�r%��bnm�H�����\^;��WBz�l{�S5�k�C���Mצ`�ˊ�)a�
��]m"���ӕ4�sr�U"4wl1��~��
�*�^�!^�$�(N��k��w�=�@����&�gd��M[:pr[�"	5aغ[�S�0�]�I;s���F�Ѳ�x)*�f�i��@�FH����M�L����1h�m���/Wk�4���x���t�@�T�:+k��TԷi٭�{��ǝ���x��_*EXn�kw�t�I�uT��ςZ6�1�CsMc�3�a�D-���&�m6�$4u$I�g��F�nM���gTdUB4ƛ��c6/0���(w�>��wu��%�x�v+/#N�\Y�,�uk$�Ǩ�`o�i�T�ٝOаtu�u���ѣ� ����l���6t
�:�w��#��#>��7:����"Hz����MP�VlC@���[���FlQ�k_+~�	$2��.TXn�κ����wP7��B��V�5�2L�t��{�t����X�RX�G���� +2w��r���0NM5�Y�s&>oؐǚ��-��m�H�O�ܨ�|��a����m�V�R�S`�}�;��}��@u�`���'�٬������y��FE�m�!�����7�3��r7�{�gƃ8�mՁ���sk�!V~����7$V��m9�Ӻ��$��{�Z��(����!�"6�%�sh�C��"�5��Y�����d��s��#;�PK�ȴU�~�M>�^��w�y;���
�ĨU~�!�y�˟��\��	�ZA6���8Ɍ��%�v��V]������S=����`=�ʛ&�\d�.!dj���ѷ�iv�1�b���v����rޚS�u�5j�;��O��C��W���%���O��<l3'IBQ�Aڹ�n���NE>�5\�5���
�-߶�f�:�x4G��O��5�x=�I䊪�t�t�6�v���]"�[`)��w_��qE��_�/=��*F�<�)X�.6l�yuy(z�u�z?�-�{z½�)Mz/���O0H���&�wV��ov���U�V��C�;Fޑ����DN�P�e;g:檺Ӧ�tMh����eF�^;��S�kr�]bhk͢y���Űs��nhj�=����p�2��r!;.�g�+Aᓡ����}�ޫR{�1
��G�/��w;{�ح�>�OĨ�+�Y��������������v+a Kt0�Ak^ѿ�=��/����~~��� ����{��p!H}*|7����9�!䵡�lC�����=g-�Y��f\��UZ���3����Gt��H͖#/8�7��a��tST��z]�U�f�xo^��P0W�4r�t���c|����RX�Y�[���]iT-�@ny�; YG�sԬ�8S��`h�ƝJ��N�C/(�Y��k��kjwq�)�t��mz��y��3��#ݼ����773az6�+;���Ӎ̗����b��*ثGt��,��o�ʓ[n���fa���p�&��<�V_W�-ԍ�F�{�jf��f]{����M�@�V�Zv���r"r� �Mp9^m��#��>{ǨI����|?`����~�{�ճ�@�EQ]���UPD_�?��F�`"-���f�]���Xi�efD&RDP��D `Q�@t!CC(@�"2 � !����0�3$ `" 
 M!d����U��P �� !�� &�� B�Tiq����� �� 
 L�32�14� ��� 3M0����Ƞ��1!�fk`�4�0(���2(���ʠ�� L�(�M LC �@Ȫ�!" C���:�BP ��  ��  d 	
d @�U] @� 2���� �*�  @� 0 �0,�@ʶ��!����(5�l����8��@��{�7��D@�D
T mќ����a�O����W�����>W��/�w���;����? �}o��a����������/������Ϸ�����1����������Q��"����%TV4���~P����G &����v�F�>������˃����oɏ���������z���}�ޏ0�~@��^>a�7ӱ�מ��꾃������_�L1��E;�`6���c��Ԁ�� �+ �R H��  P�2*�*�,�
�֐Ъ�0 ,*�, ! @ ,��)  @ ,��� J���,*����H��a 	�U�@H@% 
p�A�   
�/��C�?�~�������1��@` (�?/�o����O���=����g�u������������%TW�� �����~�����|~���~όy?����?�=����v~��J"���v�_�~�g�'����C����'�@UEP��+�P�'�4����%DPW���6��=�QX?��4�~���vy�e����`�~-�?#�����=�q����m���������c��o���v1���� �<��n���??W�}_�?6�}��}G����}$|[����������o����k�]�*���O��g�QEP?�?a��=N��|&����B��>��?'�>��|��%�����ჇA'�s���TV_B����t!�[ ~_�݇}�g��������ˡ�k�~����(+��������|���c`�~��>�ן��?�=�}���~��~/�}!���e5���`J,� ?�s2}p$��ϡ�"%*��$)R������BTR�(��A
� $�T�*��%Q@�� ���QR�)!U	J��U���	�E@E*J��"�D*�TQ%(	AJ��UIR)R(@T�U(�d��I����)*�� ��*�$R��*�ART��QD��R��"�$T%���*)!"$�J	HER�ER�H����J�*������  ܢ�V��c[nVY:�LaVkMj��E��t�Nv�&�.�qۡ�Z� ���)�V�u�:��+��;mtt�Nu@��4�n��t�$��
��EDD��^   Gd����MhhUHo=�Ѷ1$D�$D�ո�^�D�$6ǭ7�a�"��ob��*�@� Tl����[��i��Z��f���5�wZî�N�Ui��Gu5P�5ӺPED��Uф/   k�릨�i]��w]�ۮۺ�t�eQ+&kT몕ك3C�]����:�]ٷ*��P�hMݩ�
�쳆��i�Z�mK+�;m
�:�J�H�AE(U(E/    ��RS�R�tZ]w[�
���t���1r�l *5j��[]u����l��Q��;�vmt����ܫQN�ZW#�Ƶ[L��$P%(T�%�   #Ïv���]�V6طq;�]�˚���*�G��m�u��\0٫ٻ:E�k]\��S-%A�q;]��]����)t$����
����   f���b�ut�r4�j76�ݫ�0��W[wK]���kۭݳv��;���E\ik�s�α���"V�\�5k����j(�	�U) ��E   {ӕ�]� �Z�M��H�kM���TΚ��U�lUj�:�]\��n�w`6�@ 0�(i��+  �*���(
�(�W�  k���[�mMΣ5� �:�tU�  \:wM�@p[�  s��U�����[a:%D����"�UQ�  9�@:�4�N�ܝ��@:	ƪ tnҸ�	]�M�` �e�  wc���  4�Mh�A��ݪ�@���̉TU�	JJ��R+�  Y�2  �o@ 4�;� ;��I���9[@CL� N�0�c���\q�Р��� �� ��JU#@24Ѧ�S�0���4� h�"����4�  E?��   jy �*$   �)PLUP  6R�Y�V���HQ�22�*���j�d�dF�<d�ʌ��dd(ɍ��������?�|�����l��ll��l��m�m���l�&6��
���������Xn�^�ǲ�V\iJ�vhU�`b3R�b΁�)t�t�pX64R{&i[�B�9Q!A0]�v�]AvP���ҍҙ�6c�Kp'�dhBI�K�[�]����o��L=Y!&��R��w�5�2�wVol8��� �.=ݽx�@[n�ܕj�T�c����d-�H4�m<F]ثZz��T��5�Dq���n1z��X�� uRU,Pѐ�D^e'p1��Jt3r*I�qYI�H`�+t���ӗ�� �0�j�Q�x�~���l(/+>�F�
bV��&�HQ�7�5��3a�6�)��Î��#U���dE�����򵝽;o#��h&D�hzL�m�����;u�p �ԛD�ncѸ�ˀ�{�����+1Ų�҄��fd��k_H�ٰ���2����^3&�0r��J��������9�,�7�I����Xe&��(�h�B��1悘��	&fԉ'��	i@�+ �T����������mcnM��VT-�2�5��L�r��
����D�Eb*��V�^Lx�Ȱg6���mҳa�t*-h��iM��F`b��bnwogZ��Ě7ʬ@�M��V���M�
����sJk��CQ1eJ̠��r���Y"��¯�ʕ�Ҷ��1M�-�)�0,�MI,�YH�nB�e���^h)Hn�ZQ��û �=C8ˠ&�7m�˲#�n�A���b�y��n��S4�Ҵ�t iY�vѴu�-��M�t4[)����6�!�6��6k1��~�9�3-��\GIY,�d���\e�Yu�V'H*
2
��]��nLh��f�7ȩm�5�)D��JOl+��me����{�)�V���9w�����2��Z�e�ē/.��F��`�5�Շ��`P�?b�`lk++�&\i�0�l����=̼�u+i�)&5��2�eٽ5&<Ҷ�E�S�Y{e��Ė�V".�}R=V0�ʀ���a�fU���Vh���a��+��e!MlU�kL̗������c�8ƅ(X�
x)�M�hVպӮ ����T��ٕ�<�bPI�-7�Q�RKn��[�=�ɐ�_R�Z޴+	"�dG�vB84�v�:]�>�[rg�S�g��h5�J�pI�fɸ)�#@؍�5'x�ݽ�� q|�ôCS\�x�K(��v�Z�hRحX�ܤD
����xvn0�z"����&�+�.*YO�l��7%�R�a��:: /dW2�{B۲5eX�1��K92�N;Ce�kr@��,<؁�Uz���X0�bŶ.D�����shi���1Ԧ�YTji�����mZ��i�Q�ܹ��F��و�F�9�-�y3���@/qX���˴qą�M�]��_�L̎���v�O6Ҡtj�r�Cs��hj�`g��H'p��D����3F�Sz܁�z`K74}�b��>��~����Z	h��l'4��V��e��(P��3!dn�<��6����A�1�A�8qP�� Cu��w�k5�X
D�%A�3%G&�A@K�²�1DkhB�
�A�s7�T:VC�S r�f(� �/"�n"�*Ƙ7��b��;Z
��ކ��	BqnR���9N�SD1��V��`�k]ݨz����%[B��W�A]%�74�"2�7�	J��?M�&�MH���c��,#/%�Vn�e�)�E���APa��WIR�Cc7���Sr�-`b�yb�ۖ�B�^P��Q�Dm������A���h9��M#u%�^j��Lo�8"%��X6���ۼ�|v��F��6��&�B�f\��/u�E�F�lm�wH� <we!hVf�����n��Y0	��|�(�Q�v��"�ՏMĖ�+1�����J�c��V2��l���ڸ5�6��	��}��(�S2����˛(]��.+���۫����卬t�� ��jݥb�B�.�n}�ڸՊK`�ĺ"�b�+�j6�FT��O(������.��Z��Ama�NąQ�pFi��QL�ܡY�咱]��B��;v��n��g)�f��fceP1��Ɠ�sh�-Y��]ˎ��I
� ֝��'���0�ƣ9"�N�S�Ԙ������b� 7]�����B��1��7��+U5V�+_	Im0��VKn�S��v��6	�X�4�r�XH������P:[Kf�
EX�Y�I���u�Qx(]��[(�nTpj� 8�F��x�N�c@��eѤ)�W�E����j+Q����Lk�v���jK��ۖ*m,F^`����F^چ�@�3�F�2����$s��{�Q�yVD^ǺD4��z��I�b�i���P�[Y����X��� X����ݥf:�BI�EC��v���K2�w����Cj|�kLLP��%k;eY ��"n�e�;�t�V�M�!sd��~W�,�D+&�m�]R���̀8�ֶ���G#���,��K�n�3sM��KU��7��0\y+44�]^M�Jwn��6j�(���tl�//4 �ձj���)�+a�.�۽ܺ�((*M�ЍZB�\��U�jgVN�v(H���V*�NfR�D$[�7rK�ު�A=��	'RmK�J�e��w��>33VD׭�֡	���Ye^��EC��S�-I%צ��Ae8j�����Pť�b�PJd���l���GJ�f]Ķ�;f�w���YC�yvSU���Ya��57,_��*����h*��w#�&�����K `@t 1�M2�5v�i���t�&V.P�ƍ���v�����2m�wV�M�af8�el{k2�A���n��+K54�.�M�n2"3e���5>bS&�E���G\Lf�F�*M��kH�e@��oBŁb!�H:�Yl�EY�V�ѣR�n�j�:�wV셊�^7����	�5���!.6!on��Y��� H���vJU�+Ֆc�\�k6�
�FZ�Lh�vNV2�1r
�>��ȰP�@��f�r����Eu�[$#�w0l,��G���uI��T�w��r�ԩM3)� r<�wD�i뷫ueޱ�E�L��o�����횈ܭ�ԋV���!�-��ieR{�-jˤ.�6w\/	w�����f�-�h������1�����(b9U�'���l��auq��:�$���j��c�ұ��#`�Pn3�\�q�V�ۺR��Q���T��K�5ث.���
E�T�b�oc�4V*i���Ǝdn�z/#�V�휬�S��2�H���k��*v���I3K�Q�n�.?���^e3ֻ;,�i:��ׂ�"e���Y�X���2�ql�1��T9�S.�Q�P��n��E�&��Ir<�m�J t��P�X��l�v(C!�P/m鱢�	b�P�@К(��)�i[��&:�t�n���[����R.l<L��31-�2�_M��sY� kz�cjՆ6Pu��"2V:�+]D�V�BʕU�#)��]C�U�e�	�>�9�e�nM�ۭK[XڙB��lS��vU���6H�Sܢ�ṭ��^?���"\��l͢#س��e�"����qL'!����n��T�����.�Ď�cIug62(����z	Advރd��L
c�J�j4˻j`�eVҰ����]���b��+N��{SPN��XmJ�[tT4�]]dWzs@R�D��]�%:��9k,���U�LƓS���vC�,�P��03��>�q���LZ2ZU`7 WPj@��K���2,��]�l���[`�Q�^\3q�X���K3j|q[���&MM��������v�a�����9lV
ʕ6�+vvX�P���gW0Eg �gc���J�@^�E���&��*�]V�*�M(j7A��SK\��g�#��j��G7n�'&Q�@Ў��+&��CIJ݇u()�ͼ)Z"��bƶ����I�њsp�GE��e;1(�3.	���RUej�ΡX��^&��dm��)DhUy�[�>�l*�.�F�yYRں�\���cA������zH	mF(M��P۫z�dosJر����E���5��l�otZ��HH�o�6��Z�i�7q9�Q6v�(5���kj��Ҫ��6ۺ����,a'�W�2�Vn�Gae��.���:J��hn�G1�dScۚUX�!��|h�$��NK�@4���qJYhC���$��ž�5�k85٬Z�c&n�H;z�f��l%��3v�L���A�Ye��x�'��3]�F�5��	�X0%%jQ�jm R�(]��׊�婲���S�VZn��&^�E��1�B�è6�����n�l,7u�WH<�0� �$�H�1mXe5����+�snh_,�m=�`��ˣ�,�ۥ�K6�*ha�ߋֆ���,��ciR�.E�R2����O(S��twQ?���ՠ�e��s�+c�[�`���jb2��v���_)f]jՇ���Ir��a�%FT����^
Ѯc�q���G��Q��Ų��W��סnH�Mv�\�/j� �C[j9��Tw��jЛ�Fl0�e�w��#-�4f�b�4��&��[R]�x^�(�,���!�:&�= 8��T��� �J�
}�V�v�5�f�yt��$˩�"WJ2��T�������v^�a��n�+H2+kaB��C1Ɏ��x�$�i�#�X$6��{A��.U��H��Ј��V`0#O2�̄ڂ�/�kȬ]�]:
E�.���aP���-h6(RB������VB�Y*VJd��˪�VU�yR��
�n��:��OiPթSk�i�)-ּT��[����/Pt"�IL�:���O�nm���VbH-��t��ҹR�7�W״v]��t�+h�ӌ��e�+n

�#n��(K3;t�b��m��V�l��u���J�8�����Z�h�̍�qX��bo)�0�b�=�L(�A�"��:*�[�ӧn\��3A�wf�MԽ�i�.O��ZN����c]<�%��@�S�y��ҩУXx6��Ք�<W�M�K,Ѷ�a�L� %��V��vTU��ʺ�
ceG��,�?���va���QX�ի��*L,,��K�nM�O��P�0)���ó{O��Wt�82�\j�觕yj�u!
��	0!V�szW���GS���B�U����h�GC4mnb؛���ڎf`z�S*��W
6������fnPɖ�hِ1����3L
�^�nF�&�ZU`+�����7"��*+�*�&��)xn��R�ۉ�
ߜw*�]ҭv�%��<���9z�$��
��9�}o�XV�f����C�v0���7v��W�������L�$��%�7,�XKQ(iV�Ne�[pie�j��JJ�CE!�sQh���'��4�w[OX���P*�ҭ!5$�B�B�	T����se�)��P��ԼN����6��5Z(�ͤ�X�l˄2��1���M�li�6��g&,4at���a�[�U�Yf�VN���;/VV�KB�h�6�J^�A�T�M�WF�І�sY��*�D4,ȉYz��Zv2��6QR��Tgk<z�:
kF}���B�`�iʉ��c���:;;��د���t g*�!���D�a�@6y�;��t��1,���tu@q��2����fC��
I�	uPD�;˱�h���/p֫{q�փJV���T̭]�A�^̷��ږ�^�D�c��
$�K�ĥ��U�5$�Kٕ��[� ��ɵ���p�f]�m�;) �h��ʶ`�6��H���r�(��1`�����p���9��(��h��u�].���Gx��eͥ��Y�����Pp"��l5OPm�9�2�&wZ�@�b�my��H�ͦ�,0d�s�=N��Ipn�q}�ݢZ�A^ԅҦ�sf!Zl"�R�-ռ�� Vǉ��PƭlX�Uc1(Vi[B�[���a�U�7�#aT����˷$r��P6%�M��AI� ��GE���*�&9z�	���5uo�WB�-��	d�u�E��c����,�\�A�#]�7��)l�n?��2K:��kU$�V�a.��[	�{*���X��33n�U;{;Lf>�V
�1���`�i��4��-m�t^��:р��"�Ǖ�+o2�!61I�v 3$��S�Lȵ<Q��En)g#4�K+�1���5;�*��4�xq�b�6s%����M�H�G]Xm�n%���L�f5�2���:6͵W��K�aU�eX����J�����aLdFj���] ��f�
܆!�Gx�G�e���ڼ�O���[�"�U�x]���ĥ\%��1�������2�J��z*(��Qů,��`S�-�5�X �Qf­ʏ Ֆ[]
��5L��+�#�%��.�\Ǡ���G�H)�:�1�{ql{���Y>{����P#M��iǲ��aÒ�����d4M�i[��:��(5��Z��8 �fl�w��M]�Z�p̐bi4��Af���X(e"���5(E���U.h�5M�t�e=�Jw⤑��˲�R��ܷI`d�f�3R%2�Kv�ʷ��Y�G����s�	�s��J�lۤ��5��S,�	�(�t�̽ݪ���ki��#Ǒ��@)���l��9#2�QJ�^�;u�]�e�#����kr�p�ci���cvj��VQ�ZT[>TUeM��S-��Z�b7R}�[KnB�%�f@$�e؏tn�$V`�0iGFʼ�n�.��V��N���Ԉ��X�R �f������;��iJʺ�Ӂ)In��Ҧ�[@]`�-X��X�z�n��9� ;���b�eI׺n_P=��:p!�sNnq*up9�I��dml�G��٤&p���!���폲�[�0VU���$ے48H��wE��Z�`�ۇy-'�V��f�MV�\�����<�JVog0�c���c��-p�����B�땜�Y�tPd*��e+슺�:�Q�}�+e�%��p���]%�2t�+�nE'T�\N��#�F����8֬W:ȷ��qku��4o��v�KF�Y���d�J��6P�2`�6��eڤ��@L� ь��H����m�i���:fҳ��v;���@츲�(����HV�Q��Fe�i�)5\V�_.|�y;>%�t��v�뾵ǹ��q
���d�z�:7�El�`���9H���ښGN��6���u��Ԉ�{9=8�єf�9a6�n�Q#�$�n��B�Mfx-(�i���Ĥiaε�8�FݥP�]
'�6�j<�ׇ�ؙ��a�yC�c��[asǛ���\Ob�
�*��,Zd���rw�5�I�MrO�沖HvsXo�F��n s�%����Z+�su}�ԓ��M,J^tb���.ގ=�v�"��M�Mν�ó�Bqy���:lı�[�����,��좲�I�(Ѹ�A�l��Qm񭍎Y��vU����\єwX57H�EP�T���-J�.-��]�7��`�I���m��9�6��T�Z�I�$�b�Ih��<�����S��[��I{6󘽢��e�X������sk�rb�
�0l=tƵM��]#�d[d-lΫq����Z8gQ�,q4�G�\�lt�c�<�W�����峷A1縒�x�|�Y�%S!nT����z3^�;�̯[v�Z��Ǭf'[�5�q��\->8������A�y*^p�t��yݬXbi��:�jc��>-����ݣB���5e-w��t�gu0o�zN���Ď�K��GI�;��U�d��^�]2��A���7}\�b��Le/��e�YH	�n��*�hs�7��c�F*�9�#R��jy�C�h����b���ɷ��+k#}��8�� l9n��F�WV YG�z����!�*��WW+��p�����{,����K��Lo;���%�n�T�uH�Lu۳��8L�%ˆf�X�tK.�=��A|z�r��ʖ"E���h�r�ѭ&ᝫt�T���aoݜr��0�|*|{w+���Eucr(ݪ�c�<ݞ�f�%3��V�gk7q�]&k)B"֞�-�&��GhLā���J�ï���k��s�EZB�TN�k/�(�s���u��l0�(S+�fw0�Q7$�r�������>�0c�U�kgX�V����C�1
�)��d`Q��)�5��aw[c� ^&��{À���.��ò](d�c���Aq��6^�d�+7�y�/δe;\N�f]�FZ���6�]
3 ��h�AUwtm��r�t��-��e_k�t�za7o)��1��o��,�+E���չ�u��n��b�إ�m�8�.�\��1V��A��s�Ȼ���0���_t5��iܕ�\���pN!�{�m�+bM�D�%����g�{mb�<�i8JV�6�[a��F�eӮ\7�9.�9��|�;��J��>.U�2��v�i�{|޶��DF�81WEY��n�.g2n�V(��KH�ő��3%;o����R���{�c�Z��wP��;��ܔ��w[����Ж	�MԚ��.��b�w����Ygb��]�a�kr�!k.*�,�eh|9��9kG'J9f����kX�7���VW]rw�e������V�9ލ�G"$���.���4��Lu��Q���4��f5Ռ}m���C�Q*.��e��
�C3z]�7M]|&.cy�İ��MY}w�)c�y�&.LzH��WC9���#y#wVT���C΅��t���Z`\g*�`v���b��Ô��\峹Ձ�/�j���� �J��^f#[���p�-��$;�%����N�]������A��(���q^#���m���0ul�u�v����w���\l�,�T�����{.�F��;�g(;u��q1�z�d�(ֳ��k���\�8��NgJ8#VN��L���4��A�`8���)�M�s�}W��2�4Ǵ�̲�o�-�)�`.�ɋ�V��nR�O)]��kϘ��i��ł�c�tZ�7F��e�]�n�IwL��y�O�' ��v����n쯆����������H5᭐ŦF�ӥ{PSR+�s��/�#��0�^q�}�٫�:�9����wL�`��9�j���]+j�W��6��{�T��.�Y�g4��pc�ś-T���� C��,�̫��*��.��\��Σ8*��:�Q�ɫЗn;�O��C��3]��!.���튮� ;o`z��YA�P�{�t���f����~�Zw���@Fq~���Â�`b�y���{7���Z�=M�iw��2�� 0Sg����Z���zƣ�6�r�`oQ4n�y�]��ֺ�0nn�F-�iT7��W�C�ϓ�T5dcoZ�|�63���t�����6�r��gM�:n�Q1���\�yy�z��Z����L�MB�.�m7�l00������A�#z3�n%�ĉuحU���]`V,��<1$��Χ��X]�vd8tV$�ײ�Xg_i�7e����Z*-��"C�Wl�Ԉ�p����؊�WҌ��凢yR��yAN���o)n;���Z�h�ݼ�@v�Zݬ5�������n�M�����-�u�:�z�F�������J�ۜgu��Վ��y��%��*���(1t��E�=�lt�8��_.K�-5h*��vn�p�t��y�ys7�ۚ�GOk<߭�÷����R=o��ӧ͊}�,?-�vF�q�����[���7H**���w��U�n��NS�7Nnr�ԆVrބou�8�N5(���}{#�C�q�b���;��F�쌼z������t���4GsF��(IhTGos�Z:��]�8Q�W}�6v�㛄��8_h]rͧъ�f|x,gL�v��C����<�����u���K㸈��m����g��F ��ǻ$:⬑8+4�k]voeɱ���-�Y��jkq_.����\f�|��
7d#����.uaL�y*��-=�X�TV�e'x��tZ��Z�b|ѩ
}���z�$\�7X�p���t4f�񛈭U.7��IWa�0�Y(�2-�¬��B?_P������)�����r%k!o2��.�t�3��Wmfr���0�K_\�f��4Ml�.d������y�vf-�� n]ӓ�I56�]�[na��p�!��\�m@ő�l�����.��4Y����{dA	^$h�H|6����p\�Y�9ZEN�vʜ�Q��f� ��c�<i�w#�Yћ�k�L����ٍRu��F�*��epk�=fZ��ɶt�(�O��t���R��ctVs� bԦNt���Y��弒�g_��ͼ�d�k5��J�-㏶b�L��}5��+�ֺ�	,_uŵ:��X��T���_p|�{64��x�{׫�j��n[���u�O�Wu�����=5��S�b��	��ۺ��w�9f�ˋR�b��I���J�I��d���pu�b[�P>�Ttb��<�8�*t-e��"��󮫬�՝|�@DD�t>�CH����&��l����̧.*�Q���L����)��m.ε��<AK9��r�,ɎU��);\˹ue.���u��:]v�H���QLX��o�*�C|n�ч�.`�x�:7�uL�U,�A�*@���%�J�Ⱥ�1��/9]v\0���S�Q5pc�� \��m-\��d <�K�w2�wo3k�=H|*� ��Mpǹ��)��)4S�W5qS7]OR��rV6흗u-�6^֖�/�VN�G���Фܤ˒�P�qGD�/;(L2��g�{�@WZ�c�ٮ-�.�CNtn�b������o)��v���w�ƾ�޳3��:�l���V��5f�F��>�kEdF�VC�볳h�7ϫ��Gʥ��6�ܛ�1(L��7ǐ�"'O�2��T�xF�:�w��/N,�*W!\���jjpa�I�`tG��n1�����j��%\�����
-'h)����A�����Ӂ�\+�t�v1,|Ͳ�C�mb�-=&Э/���4�}�29�(�%��!h���T�4n�2�&������|���O!|��3A\&�q��4�J��ȓ�"ι�JK��5�
�[oR=Q7}���=��l$6:;�V(����6ܺӽ����L4��F(d�׎��g�Z������鶹^ �n�q�U��}�4C����˅DާؒF#>,�������^�űX���;�NN�뛨�hs\�t�t�[l{g�U���/�1�mƾξV��V-��=�f�뻹:�ŬL�a���K9n�:`��ք/u�.����c&�dy6��h�(��A�P8h�E����CHr(l7y��ΡqI�*s���Ļ��N�.(P�*]��i>�7NEDY1q}Y��-�O�nJȱ�[u0+\!�?��=���%_T�������<���x!y�j���f��՝�T�x�Z(������tv�*�i�܂�A�7xq�P�����#���à��Pd�fRA����&�I4��V���(�~�v����J������p��WV+Zͬ���B�������C\�o�5x�w�q+��W�H4�S�:���z�w�f}#��I`�p+�GS/�����K�J����o�.�,a��3}t�ɝj��ز�%nR��يr����R�W��t'9v�{a�W��	��vѧk���&��KM>o��s���kg���݁�P��L��\�쪼�[B�jaI�ԙkDg��&���,��/E��Z���m�wa39=�ގ�3�,��VYB��-%C����y����W΍�b��;�A�%�V@�voe��Ug_	!9����n^;�e;�JO�D��Ú�˺³��&[%>8����h�*U��_*X�w'|_7}��&^'A����Օ��PRv�>*�l�dRKĬ�wES6R����*4������g'wU�d�� ���R�����ٳ8�5�)mE���'>�e�x;9���Cs��$��9�X��5�v9��S�/�sw*\���ݍ��,>\����C�/������=���^uI)�T����R�*���wfp�������]v�Mu.o����n�V�\���0�^)n֬fAƺ/��Y]o�jJ]�}v#!�]H�ܧVس��,b��j�t��B���F��t�����=!0��X�S� ���i:h"kE��uҖQ��6����c�ڨ�f�7E%�L�u���P;$B�y��z�<{�wwz�s{.M/	䠅m�n��%;:�&�1Yy_Q��[2�}���$[��X��v-�
���$�Ë5>�J_d̡������1���J�/T+|9��L�'<2������R���oR�"�D���7c-Z�Տmf��g�3�]�ù�Etb*�[���+أ�C�5�f� �ͥ��o7�W�Cz]�ۘt��k�+����\���V	?rU�������{��R'B���oUf��CIQY�NK���1ܤ��P��2�+�T�Nju)b
�Nbn	ܶ��Ȉ�k�h�[ե�����
Z���hM|�b��="�O�p$Nחt�,�y[�|��g]u�O�+�l��U��&>��w����qj3�_sՋ�:�N�q��u�W&l5ڊ��p��cXΡ�YT���gs`v�V�#,X�DJ�v���[T&հK隕�71'l�"nb�-�b�Ҁ����� 7�Z��Rnj��r����w)l&ࡴ7Aߦ�k�祉�5���C��k��(�ˢ�E��"�`�z����Vv3�B)���Vl]�t)�:��a�Ƴ ӽ"�LZ���~Zz�7X��/i:�����ͬ���땦�rJ&�]����
]��V(^�r�X���w�1	ǻ&���]m�؄H�7;z�3c]��օn��������|9'٩<�i�M�{�'��b�6� xq� t�d|����'���+�cHs����V�������#b@�qn�e�N}|6�i�^��ق��2aI*�zY倞g�Z�h���
�I�݊�Ųl�vQ�p7Hs7���@j-�SX`
u�h�Wj��0�<��ȶ�tm$���˲Pp��S,�U��3�[��a��ϥ�wL�=�-�yO-c��Ӧƃ�J!N!���ۼ)[Ϩmi;�we�{��]S���KX��!͵�;!`<g �=��d
�W8���@c��j7QLW��ы�q,�4�9%���Dc�;�p�k���7f@^��5a����ӚW��mRFc6{�%"h'mА�{)k�{�7	(���c�.���	ea5���,H���JJ벟=x����/a��i�vb����B?�t�C����찹�n�cٲ�6�m\�KI���#1��
S��t��֜G6�4=+g�hWc����Q�Qe0e^��L�9`В�[q����U�謼-a��'dS_[u��ͣ\�qʻ����{�:*�B&FW^g9��OU�8�������˶n�?����mtԭ�dh�[���<��Ő��X�����o��S���r�Zc0��֒g���k�,�tm�2R�����ч��-S{/�����" �j�o~�'T�8̴�P�ۃ��%�M��[�go+v����>�g0�k7�h�.n���d0�mh�ö�o�%񤲣��f?��Z�*�����XӼ�����تZ�.�@WN��z�Z�v��L�/�$�i�}4U�>.ۅ3:�=�;�.��M���NoIx�RWK���j��Q.kY���3�3�s�����������������<=�%��o�,С�N�~���aڽ�Ê�mF�]�(}뼉��͠±I|�/�:Ť��,}����H� �m�[�Չ�Mǧ��q2
�\��E�Ԏ%++�o�]��ͪ��$�n�T�{�q�H��P#��;7�<������#va)�l��ǋ�@��������
����u��e�v�*2s0�ػLz�7C����U�]�s�A��N������+M����=6���[���J�3������v	$m93�ۺřݮ�Ǣ]đ�n(��S���w��;f��jQ���p����b�׽[)��|9�����"eLV�T�3`�GS��ܧK�9�fe���S@�y,F=�cw[�L��8S�	�l,_Fmҕ�dpϯ*����3������X#x.y���L�H���@d� S���N�J9k��k��YĚ����N]"$�6��}(��P�m�+s�������]a7:9}�Q*�R�e���M�wmu�ZӍ��E+[�9�ճذN1`�t9Sr�2�I4BJj;�.�t�}W�R �.�FZU��5k�y-�eu��em���z+���wWĬyT50��vp3I�n��9sy;��A �ͻ�z6η:㙰SH(����.|!v�Z��������E|f�M�t�5��ɦ<���c�[��_u�W�P�De�Ӱ FV����[ٻ�E֙�B�"�s���� 锇��=��	J:��x���m��>K�#����F�T�(�ŵ""U�^8�^_��C���*����R���]:�	NUϬ�`�ڴK�kM�sw:��	��f��P���L}�rjنf7T�P�<3�Ym*�N7���V7��b���������w�K/ON�b� �3L9��ӎ���i�|�=��4���w\�#�fd�ӏ����+�|��]�J�k�#��'fkY��E��hs5�0�qWV%�̴��F��o�C�4�tֈ��tѮ����\jiZ����4+D����r<է��I|��Y ��F9v��;���F2�/2C�oi0�G���8�ݝ���uZ��|̫��:����*�SXw&U�R���r�G��kWIf��}PY�kf��9�1�V�u��b,�:�$�ڨ2��C�5;
�L�F�mY�@�v\�CK�[��[Ѵ_-8��v�����*^��Hޮ�CO�>{[cS)�[T�Ա�qy}���k�s^��<�Q�.�CH6�\O�����wZ�R�լ��W՗!�� �5���sh��n�U�+-a�Ƭ����LK��
�V�m5��k��y�F�(4��L�'Z�n-�BR �u8�GB}ن��jf��Pn�*�F�νk{T������RG��%4�;.N�Ȭ۔��Ŋٺ�V��N��L=GN��,W[3�ws���mr"�
=��˫S�(Wn]ak������K�)]]���0�!GPpm,8v�C�3�hs!�c���Vf�56�]��p�|8��Jn=�����Tu3�/6�+q�wb�Z�=�d�I�t@]�h��ń�KR���
�	�}E��Y�n��17t�%k��� ��)}b���Y�w3�@Hܻ����|�p�֧r�w�	 P�_(�V��xӉ0o�[�'�gf��c��ʔ*�9@���Lu�oO�>i���J&��s]v/(��uݧn4Te����(l�5�Ph!�(�v�xgnF�C.�:@GQ>+������f����sMuwci�"��K��B�(M���X�2m=�p��hq���\��>�Zzs���u���}/��hݘ$�9S�iR#������qԷم2��\���dQ�ǰwN�u6��B�����Ǉfi
�Y����[|�]wI<�L)n�Q�E1Ё��AkE˚�dw:��T=q�!]�ŗK+E����^���}��M]��b9D��;��$���=�R�,V�W_��)�s��i,����������e�oJ�^�E+]1dꚷ(�:.t��K�X����Ru�9��ghԻC±��@enX�};[]JVT�W8vgSq�F5n;���ݳ23��)њ������y��0s���������KW2�f�;r�|���ۛZ��.�"�TͱYY�q=]ox-t9X�W�1�7�s���<|�i�a��Yf0l�#w�͊���E�O�"�� �N�����Bo��YLP&D���sG�	�m	x�L������j5�`kM%�i�:kv�����W�A�uՊgo*��δFSK�.^;e]���okFk��
-ܸ���\ۈHKRi���RQ���ԙTN����]�#���q�������h�o*oD������|٫��̏4������=Pq ���؞h�3���CX5AhG�B����s+�W�iKQ"�ů��ANhUڰ�
��W}{�o��m�<�#Z�m���5�H�ĩc 9�)��Y���u7I3Ѱ�6��]��7�;�Mn���L��:W�f���S�Ė�BF�V�����	����9�I�4T!aV憎">�W#z{s��ض�5_'�C��rL:OuwK»-9��z�pᲱ*ʓ6��}3���k�Z.�u���@fV�wD q�_u���眆t�,��Ã%��v��[z�:I�6���k r�Q�X���kevK�����v�|Yu7��r.�&tO��Z�(�YE��\9Cٻ݃��^���;(Eնk���l;�[M2ɹׁ��]�J�l&��R��4�`��)&15Y�7n��"tM��i�4kX�����LY߯��K����ne��ɑC�e>.Z���4� f�Wո�yZFe��_����7ۜ�|XOa
œ\�-��Iӹ�9��kd�
��=-���p�'4�6Ĭ0]é�|��K_oA��
�tc�g1ܔ-p�7�����Yb�Q����U�K:�c��D�I���o"��l'�W��ِ�Ceu@,"��7.�U�C��1��#T���G7���|���a��q���t�q��\J�O���=ȭ��j�uns�R�$�J��q[�_2�?k�S�Ҿ�Tv0^�5+}E֞r��h���K���ى����#��yu@�Ja�샬�Tr�Xu��/*�=�9aAv�`��.������t;\�(�u�;oc
<�
me�+q34N	U�n݄H�L�Z%<q�����.
[��^�}��|���2�B�S0�ޛ���K��������v3���(E�9@$/ �7��[�ܯ����ӯ,����[г��X�5І��!0
 �tb�W:��[����5�F�����'o�_ؾ��Lh-�'i�nF��B�
�p*v��Ƶ�`;�.�Gv�YB����a��tK��`Sq�ZH|d|�+�\�9�u�e*籫H��/���ǈ\�"��\�'��¢�t%���i�����C�j�0Q�eҦ�c*��:=-�o5]'R��&�X����A�^J���}a��k�6��N��hn���d�R��x2��o+P?"Ns*��_{��%u><0w�ze����7���v��Vg�پ��wY�B�kQJ����0���uo�}�q�廵+�gts� �����eM��S�	ܓ�}��1�����[�'f�*BM���2�`���e�<J�l$y�����Wus�]%"�w�;"�J	-�A�Acm6"CA���Ekv�5[��Zкw1��5�
�s��g@.Ft��E��o��VNt^<$�U�Q��BV�%B���!f����Sk6��:f[Ł�Ǽ��5�묉�j�Ѯ����v�%�<�:��/&<����@���3xnr+�wY)֋*�[�g
Kqq*'D�!P���8�U����ϐ��c��|&Q���%��W}�I|^_m�E�}�;C����&�8���;K��JQl������A�Zs�^E4:�.B-�98Wp\tK��j�w��c�V�km�J�8�W���T��m�b�M�}G��o0&,����չ���vһ�D3{�נ�� �Υ�}��VQ�t������ms��W�����{� �[M⧭��x��{+�^�-�7;c�V��{(���n"���Û�]5�i�M,؊��} �:>�v�{Pd��.7Zngv���taB�!�o���B�.^�>�o�ve�������P��7:��DyR�e�о	�n��g�a��M�c�T�U{�	w�j��a�i���L!ݫ!�*٣PE
���n��13z-z��(TbpT�}�c������<.��7͊@ч0]��K	U�a	Y��:J��ʞy��soF3�eN5��-�C��1W4z���FƐh�1b��*ԭ
� H�4�P��)!X�������2c$�J�Ù/� ��iM̠���e[�O^*|�o2' �&�mZ*�ܫ9��M�+��QQAn��gc)Y��M�o*�_f���˛v�+TP��rz6@]*�{��:�U�J�0)�]��qT�Ή�-R�	�ޮ��4e��W
w��n�o[_��͗s&�1;0�`o)E�v�G�j�\�8�آ�����ng
4�U72��:A�V[�Va�i�;�F-6s���;K����%\Ι�(�¼8���i��t�|Ʃ\6��T���TbTr�;KUem��Ҥ�ul��g��Xh�jΪ��pe�!\}!��-eh1�R�ht$��ʛ��O��i>�ƺx5֬��sݫ�6��{��cc�;Y��:��`7���傴���'�,�[j5��5	R�'+�:V6�b�v���v!N�6�s��n�u��v
�l�6ۮE�5�w)��b�h�9P�gI]�o�GST���;Z�P/̗$��P��j|t� ve)��lp�=.�4|��e
G;��v���L��{�`>��J|9�Ϊ+�J��n95���yCs�kg^L�kR����VD�m�N��B��DD��V�t���5f#����jw`Ԗ$��ďۢ����kV2�������tJާ\�B��q�ܣWuc��zV"4���72�l��d��J��������\|t�U�n<��g6����`2����7���5�g(-�?s貺��T1Ә��]Ĕ\jU���LM��d�]s�������o�56ftB�n�Juo�
�p����ީ���'�H3+7Ov���+��
v�9I������9
Q؛%ͽ��b�9�!'����l�E��4K�+���I�����Î_j���&�[�d
�ˬ�)�U�B�K97y��>�Y1�l��r@	;�(j�(�w�v汀|D��g&�$����9ſ3#�6�
��AT{
W4њK�c}0H�_;\:��4�^�X�>	@��s�8+���Ӆ�{ݼ��ܣO�	��M@��-5��e�`���#ǝW)w]�uы��C�/B���ھ��K��\��v������M/~Щ���9(�n���JҤ���na�S�ʂ9���7�v���=Wԧ*#�RJ}��C�}�-ޫj��6G\���]`waj2P�
۷����v�Wy�zz�I_
ѵ]��m�u��z�ɏHXř�\�y�F�iv���9,���`�z�[�q���EK�()�����#���c���M��ܧuɩιq;��7�ڏ���ɩv���٘��z������ϕ��h]�@�YUd�I�Å#	L��9L��!��Z�k8���+���/:&�9��&�� ��d��Θ�hrժ�bv©)uX�Y��tݸ f����4z�rh+�k�d��i�����n�f#n���gm�9�0D���ܔҮSMfש��6�X&cᘃ��M�nb'p\��*�{��d|��vN�
�pӑa�]P�˦���sZ��}ݸ�%&4e�W�a��yR�5�ºӵ�A��J �QXqX�ʺ8S�pͧ��a�H΀k���7��&�;�nc�R���;��^f�\e<���oIgQm���K�!-�ϥɨ^�Kͮ���@��J�VYz��U!ӱ�i�C����$6Ov�R�������<E���@���fb�Ԓ����r+��=�y�/�'ؐ�n�9t�Xv+�2.�����2��͒�ua�&5j�#��`�3�/�д�>wXV=��81ۥ��Nմ��:5�B"�W4��`�핋��۴]��`�ٰ"M�aY7�q��C����t��z�}X�`�eCX�&�X�4J�,�I��Q��R��D�"Lλr�<����[Wk��3�/�+.�����J�KA"��ڥ�XBO��Ѻ7k_P�t��&�ھ���鴳�4]�ˣ�Ű����ů틟(wA7�lG�F���F�o-g�B��1|a�;��eM�n�u��>r+H�J�h�]���5�s����1���V���
�Dl���hP�yR���G�|�p����v�hQ��uffrP��z3��q��km�$c���h΁;�(��Hhi+u5J=]���Z�'�v:�P�h>)ַ�[}Go-�z:����ڔX���[ǉԎv�
��x7]�[�Q��Ӓ*톕�U� X+zWw${z�woP��kUi/#�;���z��Ol��.��a���I:U���%{gJ5����7�+�t��x/M�C:�;.�&qj3��w[�0�$�����CGo�r�'FKq��jӿ]�W��r���%b��I���\�2������_�]gk&([�Oh���ӊm�H�J�}+*�Ы��ɜ��*�"�D�eK8e���S�v[�ge�;�ќ{��t�\�ٜ��_-K�4Wv�E�v� �Q�C!��ۏ�;G3�E-w�|�v��L&�U� c��*�S��ݿ�<�R�.z%D���=�{�x{ޟz��{��<[}����uo ��/�`��%��x�N��q3�o,����A�e�hʶ��4�.Q��oȕ���gt]�war�N�Q1�v-d�A�]ܣ=�_\R�`
��%�__i-e�<w9�9��s��<.�eu.�A��Cgg	�N$�
����J�\�!'�Sh����j�4Fs���`�X�XfvaE_��S1.����dW���_m�5�[�����/3K�o����u���gu�Y]��u'�A����|�Ǯ�>/)	�y��.��բ���y*̈`5k趚U���
]�p���Wu�<��$���fL�	ר�}�AGہ[�����)���XL�ⶻ��ft=YOFt#���ǚw\�:ҝ��F��wI3:M䕭�gb����<�OT����;>�:��sWA駮gl�n7oS���E�7Pw*{JӘhJ�icz[����.�/��ygE|�����wp��$R�${+:�Ű��w5*�SX���)�u���q�����ݸt>��=�c���M��'�S�jEC��.ޏ�%Dnޒ9Yzp���]�7W�	kF�L�Ũ�%y��L*�Rų{\�٘��(6��W����7Z)��;�r�f\m����]�p�WA�ٛ�/�f��<�e�,u�)7(prel��F�����g���}�їP�vc09	#��H������/uŅUE��	�k*T�������ww��P�;�;5Î���(#Ⱥ���^-�<�3��t'u]u5�vN�Zh8���u�/nឳ���'/P��1=ݻr�G9gsܱٝ��̓:y�N衄����K��]�2O<�<�N�n�r5�H�ny^�	\=�<�5�#�u�(�ܜp��=���Y�GQ�\�/H��r�=OE��srs\r&����ba盹d!�+����NU���j����Y."�U��+u�e�k�'��j��w\<Mwr]ݎ��x����ܲrWu��R^���B�{��ruZ�;�䚮{����y��Ouqљ��nxW���t���2+9bs<�[��*[�Xq��&j^���c�zUܮ�yYE&�T�e���#Or��$�A���rYL�<��5����z������N֘4������⫍䓹�CA,�r�]�ϋ��ٶ�;n�V�H�ۤ��ⓧP,�h]�G�b���T{�B�E�.V�uY�r�wkA���lӽ�:f�[��N�e���������~�.��6S��2�.����*��u)�r���8]ݫ�������*���ϵ�Q�b눺q�딇����z����8<)���M���ش��:�H;C[�7:Dc��7�y
*����\�=��;��ل��~a?48}�a��)����̀�]E����h��}Y�V]���!�׆I`�<��}��TCn�1J-Z�$�hq1[խA��u�Ne����b�w:X3�nD�ќ���C�ܝ�g��E}'s�഼����}'�#¶7�7�dl9{x"Ev��f"�jK݇U�^Ə�R-�d� 1"�!GO�BT�C�Fn��N^.#�8�yv���y:f�tm����Ԃ�5p�}`�4�����.k����L젹<�����\i뜢q��a���V�v�����{�O��$�.JգB%�K���Q]u���Z	�)�y6V:�8t���\;+zĩ��乨1؁��B�O	�Z��TKn ͅ����5i��㻄1��wʞ�9��6�p�*l�uu'�.͓����oD3^��q��K�}Z�M��!Ո]�9��k;��גּ�.W[Fwp'm��i���2g4[S�t��>{N*$f�|;>�����
�D�ݢ��1n�p�r�t.�{�Lґ}��8�#Gc�:S}>��!���wR�-�k�Q=4����O�����s�CM�A�&�ld��K���#:��#�y���s�
gON@��c	h� L\U!�*��kn��SD�`�l��>��R/j	7���g)��D���̸Tt��}�1y�v<9�x0.��E?�q? Gx�:�G��p��8̪�]�����uPș�/c�uY�����֔�ܓ��\��!%C`rȐ�4��="cm}n8�&�P#(JJ{'���,J�\�.�0��1����s��/�c���:���s�>����@j�E]�3�q힭��Pc7.���Q��Z�>�s�
�ˬ�6Y��{b�k��u��,y4d�Ta���Wv>s�=q99ހ^�g��2��)3e]��'r܆hr���X�:Ч�'1]婎�j���F��u��n����F��r�s!U�G�}j*��]�v� S{aZ��}޶�B+����ϓ�&�-'%`U��{��xZ,�e�z�Ż�'<�EY ��5t2���S�U�`)���Ss]2�%ej�4�7�.DR�wHJ���o|I+��ͬ*�-�ۏ�����@_t��^'6Iw��Zk3_R����FӒC�_݇Tع���>�9�+���J��T�X+�,��h�g��Iu�Ec����*ڀ*Ȇa�E�D��s}��n#��#�v��;AƑ�A�2/b�a�z�BZ\�b0�$�&��ftʫ��Ve�A�ݟuNYE��R��]n�{(y	����g��q9a���&��g��}���Vd���<�b}��V0��L�Y<��ҥ�e+D{�:@���K�]�׻;ng��c�_$d�� gT�u=צz:�Byo�R~�A��ahcw`�	=�Io.���
��|1�P8�q N���=���Њ���T�YʗC��s��w:��o��4�_*ߛ�O�H�z@�Ϥ.�«v����7ڧ��Xw=���C�=�1���	�1]O���`��a4�!@脻U1ܩ H洊��t������ٷcrh�Rz��ԛ$2|�ӕ�!�	�4���d�D�#� ��o��8�������Źy��i=ۙ`���b�*�`�4�!:�ҕM�딊2�JurZ\�x�?>�z+9u~Y�'B�{����:����[L0���ts��J�p�ELk2ed��v+r���S`�:%�2�J&���\����p������y��r]vi�D'�{>C,Q��U$I��z���́]�Ԯ�qY�� �L��cw���P����C�����*��'���پcUPw���?q����d�F��2aH�|��
yXެ�7QNQQ�VX�@��YRPl|��Eڡ�C��ݦp����F�9-L�Z��B�������64i��b`ZԮJ��W�d��7/�0,�4��?6a��������+6�;�t�2�Rcv}���".���5���U�uCЏ��[���-o�x�=���S�S�al9+n٢��i�A<�����s�?6j�q.�	}��HT�����Y'#�a�����3U�%�;�F�ָ�Kkl)�3(u��VV)���%������y�{�w�AZ��XE�Aկ�=c�"�9�(s��ߎ��T0�^�X��O}Ѽ���n.�ԁ#��۪l�Bb7P�^��ڢ6�M��n�nI�W��[���[.�j��}6r�� ϘG�:��ZD6ٛn�����ʰ�S��NV�λ�X��Vs�ߵ|����u֠ؐ!q#�da˶�M�� ^�b��{N�R��-�EΣ/�Rv^����<Q㵒��Z��#}�6��[C���ηw���>'�kh���S@U$������c��X�����8\���3r_=�\33�c���X9�$^�Ad��k�aF��F�[�9���k~�4�w�83�
|k��
>��*��rKg�"�4Z��8$e7(�8�Q>Q@iۥ�B�������&��ߘ��Z�j���ocNo��6�3��w��n�R�L�P� ,�x����Iq�*%n��n%�іO�D'U�{7�Y�_l�L$+�� ������̌�t�K~S͋����b8�2��ב!0��R*��������d<���ZN�p����_t6� �8�swS��}D�UHDF.KGqZw"c�s�@g"�)���WI�#5!pC܉�y�;����D�VM�m\ѯx�^06[%{�?��5ye��"�>�ܫ��J��x���)=��'�����M�|��0[?[�\�a�J��C�j�~���c�Qc��q�� �>�x��WD�V�'Z�����."J�����.�ȗ�L�Ō ��3��S�i�+�5�]^�>�}a�e�d8W�4s�;�Vr컘ŒZ���o����_o_�0E�f}5j���͑���Z���^5��[Y}S����rH)*��{h���>ﳹ+bȁ[=C!���Ė�=Y0z�w�(�n��OmɕkΛ~�U�z�1���������B������h(�����Ԩb�e����V�U$���;1�!�s�]��78}��ˮ9���Y�DwErE�zҋ.wJ"�HÎ��&�P@B=O��*g��T���-���"�/WT^�N�V�Vlf;J��r�~�u��۔2E��$o��W?�5�.��P<_��%Ԟ�y� \�Y���#.�^�����2hW����"��T���%�G���2g/ٽ���v��h{��T�1I���걮OU���r���Lr�&���@�D�� z]y��[��q5�`9���>_!�pA�|�O��a������0�T	X�.1��z��N38���MSPJ�bFr#_F`�D���N��W���C9�3�m�X�"�{j�:9�ݼc2ި��HP9wd�$ F��U�K�0/��#g�7�W�p��/:=���vݜO���'=j��&+�4�D��� �w)Y��r�A#$�^O��k����D#9���Kt�(بN�'�v�I�@�z#�Ej�j�������;!�6΃�o�$��"T���W�Q�%�M��X�˟"���iJ���:È9�JJ6,�kH��B#L�g�Ҽ\��CM��
5Pca�mͧ9�&��X2���P}���^�W]j�$3^����ޔӓ4X����U��m�loP���8�l�9!r�.�]��R��D{�����Re����
����riǏ���Ү�cC��9pǲ���W9��v
ͤ1΄V�G�I>Y��C�ު��=z�r���cd��ٖǔ	W�2����X�U�@�[�13Z�`;�\�1�v�<�/�����fF�N$+28�l�Cz^ر���og�$�f��9��2�D�w�F�5�!1���{����x��eU����9nC4(k9E��]�*l{Ӷ�aX���g��W��;��4����*�ˣ�5XuE.�Z��Nz���v���)l��rj�����2'c#י��(>��z��Jih�Iu�Ec�����U{��ߖ�X�,�M�e�݃�)��4	*
q�]y��i�P�"�.����&!�!Fx�����<�g�2����[B�Ϻ���(�Z�[�]n�{)	���h���b:M0&t�t�՗P�qf#'Z��s�P�3�3�Þ6]�>�q�D0�|e<�W�t���"r�;DL�آ��,j0�+u"H�X�>��^�5�١����pmd朸9[�p����wS�WxDx���ڨ����q*�GZ�S�3|��&�i��r���j�<JBcN��[b�oF�W]28���t�ws�e0�e�o=�2���ѧ����������)d�F�_�S��new��6Ln�Z��h�f���ژ9�����=]����jt�Lo:�n�t��o��r��o�E�T�\���Fj�l�J�n7 9�1#�F�O!e�%�8UQڞd"3R��2�Pۺ��[�\�t�;�U�+2y�	Őڰ�͕C��&��!GD%ګ�c�R@�5�=<*���)��C�M��.��Z���� 7�\�ha_��i;=6O(䍎@�ڝ��(�TiL@$*�&3]48`�ö���W� �ƙ�5�+Cp:�"����BU}�NcU�i�����P�Rw�B(t�6���|Ư�������H��oyxE�Y�]�Ug�f��Y��B�}$Hj�:Ū�a��+�6.���v�&�~�&��oM���p���|K%��	d��u�4)՞&�0o��U�N߸ϋUb���;׭A~��s�Osx�2-7�H�=��i��ҹ]�/D�TDu��٧CЏ��];o
�-��\l��'�Q����f�,X���c�'�i7���q��ڠ5WD�W<}�ַD���E�b�-Ω���3��K����Յ2{�HdO���eXu-��:�es��*��8uK�ӹf@8X�}�ʘh��R6��v1H��̛ �M1�0�C��N"�`����"���<���e��]zL�5J�y�-|�������To�.V��St0�Y~���/\n��r�}s����.Ⱥ�-�R��JhuJ̲j�-���Ty�;���n����Om�W
�ꢠ��ixS�1ǬbsG�bs�dW<Ep��u:^�0�V����5��[/s1���j�@��ϕ(��^���@�푳�Dm��a����D
/��&Nd(�r��U�y`�&�l��������i�����ܕ���}4��x��Oqj[�;��X}���՚��~`v~�FJ�o٨�MWÕxS�5�zҕ0��^^
�x����A�LN�"�T@gqsD��St���DF�um���S��劂�*�劼 ��>tD^vNע�#ts�д�r�'ȑ��W^s-C��@�U;��6���Q�I�:s(�ߋ�b�;.7�3����O����[�M?$+��τV�zf����w��^_j��֡�t���6�G�~���"�l�u��4^�z@���s�tH�
��]V�9MS3�&5�DF���b���]���*9yC���tʇH��a�ԛ�gu�r3�@���������x��Kd�v)Wve��؞�.�h	�{f�� {��&C�I�������vZ^<�U�9o=޷G�o6ā���z�x<�"�K!��ws�W՜�o��]u�N�⚝n��L��2=X�e��w��z�<���uv�X�e����]X�5:A�c�wȖ�շ�5_3�I�F�^+��n�U���*���ϵ�Q���"�5/ιH}��kG�N��a�{T8�D�,O��[�� ǪL�Q�?���u�:�>��#��QT�$.gE����E,�m�8�uݢL3��*b� �4����N[���ˠȿ9���h�U^��Ve\���f�O��g�������^
�v�������,� �oV���׍2�Ɉ�PL�:�7;�ۮ�7��ٗ)�7&4K�������Ӎ7��ץ����D�~�v�� @�g3<9��7���޺�̗�S9���9B�X�е�Q��z��r]ܯ=�&`�%�.�m��66'7jY49�K9qS�A���)+Ȏ&��e��W�+}.G�v<��,Տ}qQ���I�;�걮OU�������A)��U�A%�Y1W���ʽ�����K�q���(|��mk�>�M�6w��j�pqm{����꘮����(N�����T��ū'��t���ȍ}��D�9Ӧ��z�u��_9�H����(�E?r�S9JK�xc��R�{d`g;��[e��O����
��.�T���\��\c��K��b��;�W��5b3��p;�� ��l�PC6���\ۦ$w�_i�����`Vj�G��������'8�9Wc���ͮʚ��r�9y�y���&Ҧ�t�(sj�(!����|�[Iu>;f��³;�vL������o����/���I]��V�R���`��`�%nj�51��L`��"�u���+z5Z��t�P����t�V0x���ɴ�=� �y׹�[�� �qx�1a&�D�%BC�ӿ@^�]�E�,�2��b\��^r�m��2e�'w�o�k&��ζ:V��w��\{uP���r�g;c��\Q��J�=��ք�Vc<8K9��Y͢\�Zw;��yj���JQlN�Xq��H�2'V���`�S4�.7s��z/|;fw�m��-)V��r�挮ƦpY�(�\�yZDj�Ae)�X��W'�>��ȧ+��k�޽�����&���Cu�s/XR��'	�ifH-S4�2��]&��������&�]��U�:��'c�����cTjF\t��.��ciMC/N�h�I�9��]K��'��蒄-9k�7&K�4��L�#��>˭U8�H�U�� n���CCݺ;6U�	�e%a���ik����t�+�)�*[O[�k����Gi>��ݜu(AC�P��Z�g�`�ڷt��3�NΖ�}�W#\������`�}pǦE}n.��Zt���]NS���`��,�;e����Y��9�۸�<c�r�<��!�t����Frm����A���ܫ��-RI�`�ł���+�Dkhp�S�-���s�`�e+G�޸��#�ӻL�K�|%�S��$��fZ�hq[�����]ԙr���ק3���#�tS��v�	���(DMe�7r��d���w֗v�t�O���9"�/P�����4L�bwX74��l<}{ʺ�7y<�)�� ��Kb�������L�#h�FΣ���0E[�b�� V����t#b�������msV����W�!���=�&�h3,��=�㫱�D����Ρ���vn�T��tY��jx.�Wb��v���kKkS���Xc�LM }�c�c{[2��,۰�&ƭ8(F:8����du�٘�Yް�;�(Ak���HXU!kd��	P�}�aucY%� λ|i�1�}�M~�h5��W�ү��ͱ��p��,w�s{�8���L���^Z�!���ܨ��cs7�\����bl� �-d�t%�"��Pc�͢�;ۧ�Zk���2���j��|y.��5����DP�ۣB<u$��F!�і��k1%`sΦ@[y���ݗ��B���I6\�F
��l����P<����ܹ){�I�WNfeAOf,}�ͩC�T��4��e5m��u瞙(�>\(ԧ����]��TH�R�������u�k%ww:�^��]r�²w<qh���%��w*h�Ď�ʹz�Ѩ+��!�jhV[�����G�{�gp��!<+��{��duԥ�T=��<]�q!\�;�y�W�3(�������[L+B���sV��{��E9���t���g���I��,�'+D�r�FY���sGu�5#�"�,�'.��9	��Yx$��::��J9�⻆��NI�i'������n��hS��QOUTw%�+7]��ub���[�S�yr]��e$*�M��Py��.���W��*�T�R�y��
%��D�n�Nbe�E9��Y\���B�����n��.�Ip�t̓�����hEE�"hh�X�aw�Dr��u�R��*�t��|�s��|,�+�a�Wλ9G���uB��р)j��a���HxI�;"ȶ���ngl�i6Cc�v-�x�*\�6�vp��G�>��G�	? �Jx�c�BO�ro ��t����ۓ��<G���~F�!�|���q���{s�@G����]�>��" �?��fϙ���[<�Oձ�s����=�����ʛ�|�&��v��'�߼����j������0��y7Xz7眻�4r��~�Ϟ��oG����$|G��#��O��A@��n,�I��yq̀�B �ή�\p����� Qfԏ�I����|�'�|v�ߓ?�	��:v�����I�!$�`�����y>[�מp�|��M�?':O�9\�Aɑ�Q� �0s�14}['����}d>�(�?wG��� q�X���HG�$�_�9����D����ϗn}}��~O.'|/��xBv��|[rrnw��xL?nv�O	>�� !�<Gخ��8���O�՚������M����m�ܮ��σ;�����{7���w���8��񽧤���
<@�<	~tϼH$��}����t����/�o)��.w�v�!����w�Cf�I{Rz^��$���O0r��{����~������ |O<G�oo;۴�<���')wc�H� #���&�<���Z9�{ߟ��0��ߟ�m���.��x��ʸgv�hg[���zs�T�n��¸�:#�]����O�����yO	��!��nw����z�	�]��Ϸ����=��	��;rN��;۵����;zM�	ӵ�?���������n�1�y� �H�ڊ�+=S�N�������@��y�����<;˴��?��|�{q�\�{����P����<;��C��90���Ͼ�����®�G�<&�����8<}��N~&�B>�"6���i{f�^��~��ȯ��߽;|M�H~=��x_��S�s�������a�s�3�Q qc�}G�������ù]�$�����`��$���0}B��"��'�}t��Q��|ܼ�]�о�3wn�N���e?���;��˧}k���ܜ����o��ۿF�����&O�������$�������w�i���9=;xy����������9S��nM�ك�y�Ғ�=P$�Ł�qQ�7�c594	��j�D�X�[<Q,�CD� jLhT�l���Zǳ:���B��t��-\<�a+eW�^�]y��W]��z�u��ڻ�����N��4ا�˹کKP�}�x(H���u��v��a3\8m20��q=Ӣ<ͽ��~�;P�G��I���I�A�oo9w��{o	�7�����ߝ��z;�N��O���>����~O�9>��޸����n��q��8<|��G��8��A����b	@^_l��%���������v��>�`���ސhH�y�#�}�{�x�t�A����}ǿ��>���ӽc
�������Nͮ�سduKT��SK����m�˽;��S�A�	7�$?&��r��C�����'�q���ɹ	<����s�'���������r0����HV%���#�>�>��=���{�����F`3������1�뙡4��zO�|���N���|��˾���ﯢ��xq��97�E���:�~�.�~�Sx��9wq�}�/zÎ#�G�>��*��q��2��3���-�xE�ſz�>��#��tzȢ�������G���z���ri	����S������u�?S���s�j���/�?;I��@Q��yBԀ��G#�=�7�⁌١s������#��Q| �̀ ��0��߿~�o/�P�o{�v��	2�O���x�yw�k�������o�'I��y�I�=��	�۞����ې,���B�>G�D{�$��MLy���?��ݹb���ς>%A�0� aX�#�I� |}���<	��9�o.��(s���!&������x����Oa}�y@���>����ۈ�C�}�"�>�+HqR$N̨�j�Y�����dxV@�%�>� 
�${����y��@\��>��ޏzH�>�z����}��:��"�|����ӎ|��z?~�x@Q@�>6G��k�$N�������\E��m��/��M��2}�"�@>��X�^��]����|��L>O�����N���>�����󼧳��y���k�G�#̀����޲.��G�����^�2D��*�DV�N}��ni��?'�}���#�ȓ�>�#���^�������7;�s�O��raw��q�q����S�x�ɼ>�{C�|�c��&_�������?$��k�ʟa���|@G��' �}�����tA��X�cnL��*������cf����x�H��gN��k�ͮ�e��O��'t�*��k)�wE����tvr��k��KZ�u��J��drm>�{��$�`��%�]v�fִ9�t�v��Qp	#ks��v�bwwrQ�nu���_^Ԛ���H�G��@����c|Og�<.�� s�����w�ig����ˏ%q����rr�y�ޣ�!�ܒ!����7�{>��b*=$� "=��꟔d1qy5��ncX�7�ᲇ��}�s��8�x�����nM���xL*׽�C����eY5�Y��y����nt�N<����[{w/��G��� P�> N!����%_�� L�]�y��_̟����抉��A���F{f I���7�G,����:��3��������������z�����
����ǏQ�!���zv�w�k���xNv����￼�3�3�mnn�'�7T�ۿ{�G����NNW�ۿ�����w���#����<!���þ�To�����.��*��{�o���~v�=��p]�?8��슏qG�>�4�����@�<
�VF-s��U9�.Y�Q��`�a�g�e���u�Rw�h��v�ߐ�^c÷���]�����Rv�������� }~�w�\.N�����ˏ�%w���7�ߓ�r��v���0'~}?[ț�����G�@����!���q����yw�}C�z�c�Ą������!޻��o(Rw���������P�¿/z�WH�=dG����=�>�>{a�トF}W�������3�����}gߏ8<���['�וp)�;���ŏ(x��N��<���9���nw��㟮��U�E8��|C��½HA��2��>�{��Y�~^�(�3%��,��}wLzHG�$����oHro�`�>�r�ۏ��q�I>�<������Sr��xO
�S}�|�rw����ӵ[~~'��@s��T
>��󴩾{~O}�~����L-R���6{������{�v���i| ����E��O���O��q�r��x���~8�C����Ǌ	2�'�_�x��$�n���x�o�ܛ�y>Ǉxv����I��� �_�{{�&_�Z�����n{s�!T���M����p�]&�\��'8��~q G��">���<�!�������v���]�O{�pǴ'~���yL=�z�S���!ULQܾꟶu����@&2����,=}��地=����>�[v�*��|�Ԃ���n��^ʸ��R
ţj��.��P��ʝΫ<�+�*ڼ�Gj�.WQZ�3F��TƇ�G쏟_fF��<3 ���6ns��]G#�����.3^��G����_v�����ÎN~;s�o�yC�a_�<��𛐐<o߯��ü�O�6�S���ӽ�7��xM��������p)������I�!}�I~�&��q�����wx�>�>Y�����.��P����.㳅��#��}�A��	#��eo;����M���xO	�߾��G����Ʌ�w�����z�m�c�}'��������׿9��>�#�������$�@�ǃ;��졝�s��Lcܣ��>���q�>��$��>����N�>������*7���A��Auщ�S��{�?&��G�>�.
#H@��n<$���:|$��(���Ӊ迩}��e��sa��u9���2 d#��>�Z�z����Ν��������N��~���Ǵ<�Ӵ�����y��t�����rs��y+�����������Ǩx#�"�!��4��A��Ϸ*z|��EK9���y^��f��?����2�G��|4���ۑ� Q����,�?��ߟ�\N$��v��{�yC��^��@E�� "=z�����D�a�t�}Hv��<u���o�_ ����9�
=���Me��̓�{�}�}d� H����� ,C�ú�|G�����"����iW�D7`jf��@�#Tѣa�L_��#��KZ�x=>ݽ��M̘�Т��Yu1r�>0�%t/g�����2�2, �3��9�&�z淧-�vwO(y�f2�yw1��n�k�=\g�'f�	f�Szo�ӽ>a�1 <���}��ޖ�ߛ��Yq�@~���B��UΏ���s���>�$�3�L����"�E�� ���;m2��ᇣ��$/b�N������F����q��`,d>>�Z�Qڕ�������d���wC;Se��p&��8���T�v���j�g���j\���N�w�9X\T�ɣ��l�o.��ruU�[t��sDyݪ�-�K�"�p���gf��v��Uk�.\�;;[��r.:$u�'N�!�2z��V1y���A�(9�g/�S�A�jV��ipr���W{k}k�cڞ}����/�jA�Rbs�����-=X}�����A)���Z�2p7n,ӷ��ot���L���)v(��9�Wd�4�ǣBmi�C{w,���>���vx� 2��t<˷�<D�0�Ha�Q3�C�#>ȍ}��ic�:n�����襮�<�V����c���ﯝ���^�*��{�Ą�;*�9R�����n䭩���{���~9u�r������ݖ��Y��O78MyӡM���G#�\�ڎ峥բ�:`c�,UԼ�7%��w7�����#(7!nt�`,���'�:j佅jB��Y[��1�����'�s7�L�r����^�y^o�RƔ�7$�\ɝBRQ�9ddon_t*{y��ڈ>�'�e/TmΙ~��:jG`�u\���y�8��)7�w��"A�y���u9;�F1�*��T�����Y�mt�B�#���&�5��{b�k��]OR�Κƣ1Mo���������ˣ��e�8%�죜�=�w��WJ�ɾ҉{�ۋ���*��c�-C��Vp�s��M#���蕃�5f�Z}h�'#�_I�Ӧ�RS7��:�vi�! ��/^�V;����e�LkS_p��J4�|{�=���_$ȻA�o�*͘���b ١�{,$+�nW��8�WB���>�r}�/�;۫8�C���{6� ��+��x��&3���[i5q9���,���Ea����ϲ�� ��¡L'K��7%�$�N[�h9���ϔxj�vˣ^��=Z5��XySG�s��R���ż���=�ybLГM-��<u>�Fa��P��^ (.7r� �T�S���׵d%���g@��&�q������	j�{+�� M��M��!�w#�[훒(���H:C)lkYU�e1��tϫs����S�	ջÝz�{#����'QMzA��j��\��C�&��GK��^�%.^3�[�^��N;�~F<<`�N�A�떭OOH��\���J�:�%\7�g4��������׊��wq����	ԽY��N�^� ���ณ��H��?�s�y3i��Y����w#U�:.נ;f�Z#٥I"!�i��U��@8�tB]���r������p֧�N*�a��9���`c~�/�.��S�xԥ�����G�ԫ�+�����C�;�\h~]�Q�t��&47�I�v�Ko�pj�Z�*��p�(���5ِ���|����}�o�#N�S��gIW{Yʤ��^;a^=��¤���])�S��C�)���/� 9��`��ũ����sCK%�乀zl��H囼�����k���$E!�͕�3�3����Y� �q�a	�ҕ^n �2��ţ��y�l)��m��Ć�pj�����i��ubU�~�����w�d��lpx�
�p��跹f�Ȋ�d�c�Y�:�+K4��@�b�Ë�[Q�^�o�\��!�N����s���I��Di<rZ���+�'fb�k��@��#1Wk��>�� �=-�^r�Yǩ�m:X�ڡ�[L�!<J������Jg\��*"<\�d�6'Le��|����;�n��s:�)��r�� V���t��M,Nr����}�@"��5e�Rɯ/��4ǆ{dk�b l��<�#eY1�^��G��C"w��eXu��RP\s�ׇV��y���z'�M�VV��F�f��צ!���yv�bsG��>�x�^ˎpu�4��N�ː��;��a����*��Q��U��in�H���d����� �v'oU�y��SZ�	��F.��"��Y������t�뾡��R%�+׈o�Jx�Ц�	V�1aʳ�\,#�� �4\f��S��ɰ!�8.v36�l�dAg3��pM����<��/�A4k]N�õՑ.7`�1s����6=/��tf=��]��u����ѷ$�W:��Q1�kơj���]>Q�^���&�+�9x ��:7�:�',E��Y�қ�kZ-�rOb�-죕��	ml^�<Ll��S�u�O76G�n-a���W��� ��V�����-�4É��(��s��*!��U�6�������\�_-��xWx�9�"�gN�s�д�r��<�P>���u�)�yx���נZFY !�����F!kؓ[]!���t��d��z�������X�n����aW���[����z���OJ�r�}�4�E�A�ћ��j>��Gb
��$�S������<���vg�Ls����e��Pl]�P�%��7���@{]�빺C�˭<�&W m�x�8d�w�W4h�^:�[~+݊|�(�H@ǻ:Y[����f'�c��q�A�vS�������&��w��h�mO"l��.��4�]�����;�:9��m�~;S�׽�:��+۔k���jM���UՆ�S��5�TZ+=��=R�R�i�jG�����G1^�)���5�w�	�����;8<7�<�j�i�n�zn�`�o.����v�����=Q���\��D�]K2<�Z�^VdX�-|:��v���ѷ�wQ�h_ö�f�W��k�*��mi�`�Q��v����m%QD&Y[��8���hs���=Ş�p�~1��w���[��s.�"����G��A�S<��ӌ��q��-�C.�1W Mܨc�=\b�Z����f���ό�<2���8���Μ����__���W���=�ˏrG��43��qW3���u���-��ڰ.�γ���z|�_$dS���;�F��,�����n[4q���Fv��S}n;َٹ�O'u���CAZ�������1y���6���ob�׊��j�{��𡧰3�ǉiyJy�˿U��Fb9hm@\��)19�OV�Zx�/q�>����8vu��~��ؔ�� J�'��8HխFb����Ɯ��h	�����N㕾C�v�y��G�7���r��#땤k3V�N�(%�C�#9��3ܣH�q��}^�n��H)ܬiOf�o(�8��S�@/x�`�y��yV�t���#\���//�����ɨ�>`�`�%P�~���֨{��
�<��np�� �6�+��G�"�~e�F��*;AM���t��������x�U���X�w�K���u��#]oC����摃e�*.�!��lp��e�Y��nGǩ�nz7�G�vMR1;i��/;���È.��]ؘJ-�w�2V�c
��9������`5t����O{Ew�֩�ح��f����ܺ)�U�:.w'����D�Q����)�.Y'4L{�zO�9/G�9@����;�ۈ�u���d��$��?&���
Nj�U������}z�4�ot��s&�l
I$�δ�m=��ޗ�|҇�B������U��io���C�_MH�Ϋ����	��b�&DU=m����� Wug&<�C<*�Q��؃�fv�q!Y���l�^ޗ�����zO������
>���{�U�<����3�eU��qܯ1�Z��(z�߯2C]�7�7�Q���hߩ������^ᖐ~�~�N�S8�jS�􈨳I"�g5��^bzV���}{�b'	,z��#^�rJ�{;b�{����z%^�F�>'E�K��ϯOu���k�n\��O'{NH��s:�P��C�&�R7��{�w^gk�4���q�s~�Vp];�'u�/�5�^�4�1r{6�L!7�}�\2�&K]j����J��mը;�@��X����	��)��"��&�dqKcZͻ��C���g:g�1�<m������)�<���*�Ģ���m�"Z�iV��`F�!᷎�4XxI��R���l��f���_N�ʔ��Ѷ��/����oϰ\�l@�mq�f�+Grr�n�J �ey�#d��.�/�O��+�����7�z�<��u�f\��4�W2$�&v�k�ڜq�T�vvv<G��"�p�ÔqR��쭵�!�۝���%�t�+2Q�P����,�lqz�T7�|p���qɟG�i]}���V`n��K5�'Zgr�U������vF�Ǣgs����qx�3N���$��X*KN�/2���^o�mѶ�X��>m��A���{v6�u۫��GV0��R6��E�^h�E!�1m�����~�7Hu<�����9|q˨Qy�u��Qq�H��k�g_#Փ��I5�3B[1�*Y�tn�t�je;8�6��mi��VAK��U�"��.�MZB����q-|B��GX͸�,�O`8p�Qf��YQ6(�+��?v�Ы��������ȩt�)�z�:y̾�t�l�'>H!}6��ںU��D�S.*eP��Y�1�h^�/�U�����&�L��9W7��Bw�]K��9`t�m�Պ�U�﵆���Y)�{],�K�p��`<+`H���i���M�3���^^���c�1A��/r�e��Xj�h}�{���s"�1���E)wD�Uw}�V5����PCf�RY�u�p� ��8p	��N4�/�>1���{�ee������t�$r�A�]e��|���T/+u�X�.�޺#��}a�V�����'ζ���� $�Q圣�{���Շ���w�x`�V�k��.��Ƶ��;gb����s�ڊ���֡k\A���\)�. |�whj��[\�q���Ff�	�(�4�:x�}y���FN�`_+V$ i�Ļ{7K���38K��S$j=�{C��oN��b�)�uf��>Ɇ)w��q����Хܞ޽���u7�d��o�����5{���bsB�:�lb�xtUf�<y����G����û��Bi1 l�6�`��WC$��oD}�'.�;���Ӱ��v[}7X۱�y�L�T��zLn�<g7-��+ �i�2+R9���L�GBW�3:�����/��]rU��{�0�Gh�ֆdt��G1p\�I��o��+[b�`�}�#f��7Ld)�B�M�gf�C}%��v����	\M�sD��-�̻��yV���Z��� r1R��iy��śiq[w�u`�՝�N�]9��.�����d�E��w��R�De7��QYFig� �w��sX{qA��[�n�;�B��6in۱#��u
�-�=B\���kh,ʏ������ɚ+pE����Q��A�'������n[7��\Z���p%%�<$v�J�Z]�c�3�����D�]�x�J�7�'Lva�gta�nvј{ ��*q��6�w�[t5�[�2�mÁ�fҎe3PC�

"�F�F���Q"(�OD��u��w.y;�� �BU������{�ݸ듔��q�TԒ��qQQ''vn��-s��Dt��Ks�9��e9"����k���jI%�*$!&*�
rs�	#��Z�)��(�iNK��Ny�^��Q)�f��Ije��Z�H����T=p��QВS���fԴ�s=áATh�{!2�0B+��rP-�j^)�J�:8y�*O2�̈́���r*��Ib&d\S';�.w]��("�@���e����
;�'�����i��n!h���囮X�D���p� �vb����N�!�$�E�Q�r]sܲĢ�9B�4�뗮�醥f�H�R�(�����u(��$��t�<r]+b�h��/)��PY��a+%��[S�Y�EXa�Z��q9�Sh�HE�R�t�N�*.U�bu���wMG3ĕ
D���m�K�6DF�*Y$��h�E�E���=fQ�v�f���WK�u����i�wQ9ω:�1�b=��dym=�W�� �R(޸�hWig%]��:v���o{����!�w�^�2�e�#N����&[�Nj��R3�{���͏��k���{R�,;}f�B�V��ҭOOH��r���p�<&�������$Z(m_���{�wg���X�Ρ	�uuKՙ�t�V�&���It^�O/3�Ws�f�gN�q@��qM�c���`�poˠ߶�9�V�Y�	��\��-I��	v�͕��`>[4CIW��ڜǀ��rD���Xs5G5�R��NUs��3^N)��ElK�s9[�"�ޮ�H��	���fa�f�L�!Y�بg9��Ɔ�:�w�g�#�|��D{�/�&���U�Y�T�R(O��J}���n=�Nk�Չo����p�����ӳ���(���wU�cu�f����r!��
uş��e���6�WCx��x"��]z8��2&p�<W�7;2�M��Y��%���Eb�p$϶�`���X4u��u?`���������~x�;�c�7+�Cr5����%�X��+�}R#+��z�`�-��,3��ǭ�g��5�����`+ά�n.\�O��CIfa�$��qO(�O{0Ķ���-�d�v��H��I�58U��V��"/z��$�f�,�j��v.-�ng-s/B�C7�ņ%��f�fd��&@�1�h���-�p�[��k��d�b�]�A��{�oa�O�7(�T�a�_i�ng��.[� @�{A�LO4��d�-�s��5���)�K}i�ϣ�5�+��m'��֗���=�	�;��
�0PN-�JCb�!��(��NڵS�znmǙY�W�++���+��F.0�v�d�r��sm�O��T�^(����
7A��I��/�v_�`���s���$d�h��51���dw���J�K��<�a��q�oVa5����:��@D�����It��v������1�ªG���k��|�uM*Gb��?Z�k��ʷ$�*���WL������%�0�L�*r�.u���΂X7��C�:�9��P�
�G�gmoyY=�D��|V���a���g.wi詽���xk��5�n|p�k���f��:us��~J�w+8EX{f6!�Y�f�i��k!�'�-`X�̵GB<]W4Es�b!#��Ĭ���.��B�{4�.�a�mA��1tl��Ŗ�X�4�jN�.|#�"'Tt,�5�1���8<��i���z}�3^�m����h������IMT��D��gy`�CԪ�Yb�B�S��h�⓱���R��+|GUB$�B4���w6�4�_6�l���Y��c/�iB�]沐[�A��Čb����m�x�������1�&��5f��0��W?(͡�����{�{�cT��jT��!��|ɏ$a ��N���}D󀈠5rY>*b.�\v͚�{bj]��B�/o����q�R�7��3��-�L���<ᓉ񨓀�^1U3�M��1>��e���3p\Fϱ�NK.���r���M����ߜ�l�}�s3����[͇��K���Hf�w~�bQ=�t��a��g�~þ�aހ@����5��^B��X�N���fd��>��UW9j^�Pr���ER��hq�7z�1r�>1��u���de��͹�A�+ sφ�v1��.g�;���3m�W�g�v�J�@H�*�*�<*��_0Y�-%zOة��qN���(S�ݙ�6��2��Ɯ�k:c�k;�5�ܘ�!�=Ҋ� 0WCി7��97����K��'1�:EZ摾\�gyܲ6W��ᇣ��$/b�N7Ɲ�-P<NA�;X��ؗy��57�T:�59x����r;����n*p�I[u� F9ڍnWvv����H�o�b͊��ø��wOi��8,}�eN�Z;)`��.b��U6c钤�����a�ήBW��Y>ۙV��j�iŦ�����7RSoFK���\�΢�Ծ�L�0��X���Wn�{f?Yɘ�̼�΃c���W��w���6-%��ro�����3�����C��K��}��x96F��*Y}ۚwm���]� ������l]��TW&	:m&L�j(b����ƯΜ�'ɵ��o?���4q�*��}�9�x�l/|���.#�%�A'wB�\;22#_F`V�uW�z4U�tSK@d��>�:_U��;]r۝ԭ�
֘k��P5{��a4�o���֏\�:�?F%���w8�uM�4��p��x�M�%�d�Y���Ȍ&��^�S吋��R��{׻�P	tm�ِ���fɯ'��D����nt�e�$�Ɖ莅��}u�Ft�Nt�<rw�Ԗ�6�`�YQFX
N�����U���@�Ա�)��{n�_�m����W?S�K�QQ>JI�0q!\i�=>��^�\�S2��s_>(�.�½����X�mi�93�o�^�wϷL���L�p������`Y�;Vdmt�C1q}�&��=Ǳ�����V+�����P坆�'1ƺ��k����H�9�'2��7f���!.6U��ڪ��3�aap'�ax�k����Hf��5����:Ч�'0/G�oȝ�&g �\����%�\q4u�277D��u�$��{��5��Ò�����CZ�RP��^?�Sw+�,z�c�E"�v|���HG;�o�7���f�>o�)�W�C+��p4��RoZ��ּ�N�׈s܎�;Wte7��n��wMU"�^ΣfE|���+w�b-�xxa�Df%��Mol���>I��v�s��(>��^�ł�G���ufL��~xd�;�xGHڜ�j��ܫ���Zig���{����Fe>��Y�^_\�z�pu��9���p���K���ݮ�_8�h���ɒ�Z�p��ξ�"�Ű�ov�w{�s��F�^8(��ȃ���|+������\etT�yޞo=���Ƹ��g��9˽�{����NHo�=*Z�x�cښKd(�`�ԉb��Bv��ztJ�������^q�$�Ll�ܾC4�BgJ���;B�<�����KEԂ�Ѫ���ɼk5��T�O����P�'���q'�p	����豨��_�.mM�8�r�Ÿ�R�p\
�l�-gD�y�r�'Cjӹ��su��qD)=�Os��=�v�s/QD���
�N�v�9�TsXu!x7���hi�N)��d�V*�s[��/8^�,\KH�ꀱ�� �ّ�4Y�Cqu��shz}^Z5�x\̷�]��o���hw]��5�n�*7��/2�GO�"���+v��d�`:����.��񧹩p���kF����x��I�z�b�|�w����lԔ�s��z�����Y}�E�ǹmMW�r�rn�۸1�;�O��r��Z�:)��}U_}T/��vÌ{�r�J�� �Eȡ#!҄�j�MǲJt���f�ڝ�=�Î��ծ^��o�&�l{��:�/ ��+:�[@�^'X�]�,��^Wc���pVa{�C���qq])����nnވdoc���V)�I��SO�rW>*���˼�:�;���;�kE9s��)�dY�nCj�+i�K��i�숶djZ2��z��p���wa���t�y-��� �|#B�~Řá�H`�Z��[�( ��(׶�L*�u���w,�2Dv-y����T\�(KK�A/���lB��j�ĸ��ׅ=0PN

d�/c�U�a���HN!��o��EZ�C#vTq��Q��LC!�e��TǴ�1WW.��3�[3���˟�N��mgy��{c�+P�YH0���<h	��QQ-aa�..Y������7��.3&H�17Xl{���[�{(u�BøBէ�\W��r�c\^@Jٮ�F ����D�x�ؼ{��֋Bط$�+{ގ��O��!ͼ�˗��`����*���aG]�!Y����^S�;��VS��Z<q�i8N�ɥ��vv��f���^�`S[���Cq�9Y����;N���@Pqh��d�VP�|4��v�Ϝ��彬���s}�Y����;��ؘ2�]0�1��D\�eU��y��7����0�v�L�|!q0@�$b�P�9����^P��.���s�FH���|���z9KJe���L�
�;B`���Wtx�\�Ð�R/�t��	��1+&�"Iu���)���.[]�j���r��.[	��<!kؓY]!�����Z=�̖*d���''M!�3-����MZB�.���GH�+�f5�1�P�~��:
�I�zr�3}.>H��᝵��cӯ����vg�O8�Ppj�_0G�ױS��h�����%orn�qȯ^Pdg:�w��Ԫ�'��p������l4�-m�l��bȝ�P�]�="�`���vk`�9ڻ�r{.,��7�V��Ir���q��MƉj�wu>bs]�J�0�#KU��9*Y���Kb�ܮ�WD�kb1�N3 �׹O����P"X
��uƠ0�<M[5�ʅ�)�g������9o�3�M��˧��k3o��$Ӻ�M�U�i�{��F�[��P`�	�i��N̢��ᢕe���@����|x��̽��.�{s)�V�!��}ܚ�w}�y�>��:�tי��Z�ֈY~�t�m-��3Sp�|M�/hmf��'�t��{�����BK̔�YKU^��F,P�L�V�%��U�黽@�,�*�W���H����G����'�B���vآ~�H�u%O�����]��W:���*����� �T6#ۼe�ڻ\���{k$���2Y�M�f�9��P���������]�q�Ч�y�z�#�7���M��;	�>�C5O�
�7�T:�9x���!�9�K9b*p�sٽ��ů�[/�Ҟ�bɯT>�t� ��T�r�ڀ��/;��֋O��8p�I+�삺<��oH��O���/�����x���;�P+�z@ۙ�Μ�kM\Λqa�Jp�h)�]\��"�s����ŵpϮ@p8��0�N�N��A.
�ȍ}��i.e�L2aI�g`Y�{\�bǖ�҇�.�Y�m�Ab	�q�� �O�bB=�eo����v��T�����<���Y2��:ᑼ���	���Jy��h:��(x��?w���3����Zu��L�u�ȥP�ٲk��؈��be�)��L8d�#���3Т�z��ÕW\�{�ꬽ����G���= .ɳ&r1�`�6���H�CύƠ$S���Y~�'�ujn��.�f�P����e-v���Iػ	���O -JO�j�vD�>�ͩ��y��	�>�wZ�[���Q��g�[{�;cǦ@�xc���������j�D|��֕[0V��],V8j������uTvؼn�|����3��iW��6/�V�t�WF�
c�6��έ�O���󎷻�'�(��~��hvW!��f���Lux�{Ő~��b�(��P;h���՝��Hg�#���Ρ�/i7�w�4��g�Žry�=߃��{j�-�f�}�	
��>����<cy��'C}���+Xή$��r�r���_9օ>�9��ܟH�j�s!U�z�xeg��B��v�^���8p4ϔCԶ��Y& ��hl��ׯ�7��t��t^���7⑵�	N�d-�D]�e�I�"���C"=I4ҝ���י�4��]b<��=w�룆�;�X �
�Zj�Bg��=S�mt�B�ǻF',�ˠh|3)��+"���	y$ܜ�O�[^�N-8B�b\"��&�S#�����ݵ�tT�����s�u��fU�E�?_<n�d����ڊk�<dV��ĝep
��$:��]�9�|^��K�go�:�I��	X��.����Z��w/�ƍ+,�T�t�P�=(p7�����o%��=�R��܃�L��At�<y�0�No4�p��R��s�<�rx�A�"�s�����W�Y�S9�Ǒ����i��W]N,'���A�weL&`�{���n�;!�TрbK��p��ռy򹷣�WQ;�F�"nwg�E�Я����y��ʎ�)�f�r_�j�f=�}|��W�7CI釪��ލ&U�P��|�-���gC�Ζ6v�y�ϗ��«ء��D�նtO��T�
vH�m�x�X�m�Ii�����X���C�s \/��YG��$l�jØ=�9��2F�ӕ@s��3��.��[W�d���9��S���!�EG�)V�P�a��^K��*1�)���BA/5��r-�s��6fw�ԥSp:="���J�5r:�Z�>��˵ՉUo����mpzM���-n�޹��:ʯa���I�L���pɅ�Q�㹂�d4�M��c1z5Gr�x�����f긼�1֟T2;ov����w�n)��QX����B��&�������ݱ����bJ7�9�7=��E��j��[L�E�Rڥ;"-��h��ּ�ҕ7<���c���s�q�`���7�د�ڷX��p�2��M�J������m�����l�����K��8�̬0{�E+��#���K�iy��cڰ���
5Uowʽx�}��~���U�!��Ù1\�+9GLuq�gs��(f�x���^�:�ݓ�vT�l��]3!�=3pŗ�5rͫY��B/=�ݕ�z�'b��~r�f�'��|���k�J�EC�-�]V	�����KAt�ޠ 6��:ٳY[�˷]�R]�R�Dw��R�u�h?�e�2���8[|i}r�L�N�X�6�� ���]]�l�ٺ{Q�K U�F;X��|�l�{G�q{<]!�l�KTBh�s�κ˧�R��`=
ݧ\HX{l31�>;��+�5Mg�;�d�ʑ�Zk��kx(e<�'����~7�֣r��N�EgA�p�܍��}��U��H��:.f쾬��	َ6�J���;�vԗXBu]�'=湱m�`��d\ӭ��ǳ��M[�R'��.
�I��εOm�q�J�S�Rc���GZP�ۻ��.�QT���&�%V��
�-�����C�LC�_wF���^�sGl��Å���M� �j�LZ��2Z�amʾ}���|��s�[�]Pݫ61�P�,.�ЧX��3E�Y�)��&�#{�iޥ��Wu$ح��xݮ�wi[q�B������cJ=������2TK1�n��)�n��&Z�v'Uн���e\�v<�ke*%r���#���/(S�+>h���+��mv���X�<�6�ivgʨg=��g>s'aӪ�]��{���_'�����������Pwͬ�'A�� �����ct����h�%s�ݵۦv�c
�#��"�a��=yJm���Fu�[�9�3�/o'X�pȥf�v�@�`��76q|�u����B���;v){��cT�<��$��S$��j�kd�Q9�s%+Y����\�L.d�m�թ�w�uBr��%�s>�,�xr���,v���rU�q��m ��k	��VY�mlB�i�VD��e���g%�hЂr:/�MƳ�Ί�X��VNr������
(�Û�kΠ,C�E u��PFD��˼pKO������v�C��&��6M�[GxDr�,�6�GP)K���&:�:���+��(<����Fi�߉�0���tﺒ�'1�5�w�SS��}.0���ͻ޲�3�Vs��x��]���lN����q�5p��
ZG��Q��Q����d�S�@]p�6�y.������sW\ԋ��:a���Hm8*}���8�Ǯ�w�s�/C'���tC��ی}c��;e�x�b�\��*땄�w�}l)�^;b�[���8��EHq܁B�1^oU��\���4�yi��j�0\z�8򞒧N؋��"����yz�|�y] �@	u{u�&�/���b9\}�y�-��Q<�Wv�TH�d��\t�T�S�M����m�J���O.��*���5S�sr=����;�/�"Q�-f�H��u���i��=X�˺䯺�QTcÝwTv��u%1Zvf�����5	pK)E����[�!�Uy��t��DC
)4�g��](�E��f��d�efԋ
UP(�vdJ�f�;�Tz&�a9�C-�J�G"t�Z`I�r@�2�b�f��ԍ]�ȩJ��2S=S�,�jE��N��VE��H������E�+V��	�+ݹzj�$�rEZ��q�<��*�{�TQ8:�[��/0�V�⮕yEI������'R5�JC=\��9BlȤSLڳEp��pƻIE�QAT�:9���*�3ݞ�%fh`Nx^T[<��tr��*<$B��JJ̥A0�*�*�RTK6G��Q���ʊ����
��QYUa�ځԣ(Α�5ww+�H���%V�R��J �C� b$�U�c$Rċft���:R:�uY����T�Qd�	3e�V�K+9�d��Ȋ3R�Ze��ՔY�Ѧ�UH�e�S�)27ut<"5��uԬ&���j�[Nr�$!24��Z�Iӑ
����I��U�&�(��Q&�_�4膞[��E}�2��U�J;����fr��:���YYO:�|sv�;@�3�LebW���x~�;�˦���磌�����"�F����}��T6
o���Jb���F�(�@�\lLC"}��yw*��L]յ�1�_n�ˬӯ�ω�L9�(s��۩����0ۘ�T�##���(��hs��]��8����|���₳�y��17Xq�8�rOeu犣q�5��mA�x�S��t�Z�V��V9���|���yDMg���hwk�z�2�ִ[�G+�}άv>�.�(����k��5D����0���;��w<�ہo{�a�g����\aW8$agu��k��]��W�{8b�q����DV�ujp�Gt��\���j�Y����IsDK�8�Jyܣ��e^�Wi��,��X�Pg�)�L"9�D�����^q^��!5�7-�l���V�LVeif�o�5a!\�P-�J�s��J�r|������ȉYj�#I*6=�h����iz���Y�3@�����i;�p��`Ϩ��"#W����[�9(�B���7&��Q;�s��*���F��t�����-�x���N���x�^7�M\��U�{ՠh�����IZU��.f{Kj�}�m
�f�AR�c�4%���#��~O�$�tm��i��uq�aG��"�UMwVM��xBr�:¤:��CTڹ�9Ƴ����Q�ʯ���V�<7�N��V�X7Eʝz�H��{�x��mK�ܩIW��sFԜɉ�zp}�N��]q��`����8%҇}����]����^�������24�L�q�U��v%�@ݎj�r�x���k��h�f����[�١���Dc�a�R9
*��$.P���j�#h�>&m��<��O�u��d.��������w�m�^��Q�����@]�*�*�<�'g���Շ��L
�e=��=շd�`bLW:֠٢��L�R~5>�Uν6nLh�Hύ��l����M���>tT��n�?&cT���_X�2Y[H��sq��r��s:Y����������T����.��9��{�-JJ�3Ȭ�8A�C�\���T;K�k�y���A�)�K9W�(��&�ɧx�^��^ګ�+����GB\�;(.CuA��OV�Zx�;B�s/���佝s�e���_�Ej�If��F�j/�w/m�sN\z0���j���U����n�[��'���`��g՞p8��0�HЉݕ�"��{�̞�p �,������1F9V,t��a�P�����g�v����V�N�NAo����8��$ٵu��1���퐗YñFo*,y��k�.Ӎj�����{�Ɏ��!��TpL�j��
.wwC:�J�֯��1a�/A��!t;Zqb67���{�7z{+���SuD|/2x�C}^��#�X�;�U�Ab�a�G yi �Y��7�Y��poK�����)�~������ϫ�n9!Ś<����&�:(&�����]r��`/��/�h�EFl�ڂF�3��-��L��%)��r�8kǍ�t��m^����m�����/b+ּO��F��c��c|q�[�ڨo<�Po�A��ҕ�ȹ��tDdʹv�ی�&郓&�RJ�kbj���y��]o��*�9�:�j
��t�/v)�[6o+P}��!�p1�β�N�Z���@��HAڳ>�3�2���R�gK�, �}ÙWj�M�5�^ؾ�'��g�M=UJ�%vW�v�S83Wi�<���3�^E��;6l�b��&F_Hf�CXUk��+�6�
�=�Q;�`�N��;��d�nW�_v:l��c�������'m�7����!��ǳ�+�N�^}s�r�^Kg,>�ǫ�w+e�:ϳ"T��F� �VD0z��M)ގi�;�3� q��pJj���2n2�ݙ�S�6�.��V�;�,��,�Eu���#�"?�ؠ�mi��Ig+��[\�K���y ��n�Qy�Y�v{���������u�[PtP@��\��c�8���9������]�%�;�?�7)�S��z�����}U��K�|�����*�������pd�I�4z�ti{a�L<�YS㎡8
��� M�A3����^��$eJ��pG�c��>�DtWC¸O�ע}�5��)y1�@�Yr��{��(q�[����a���<�y�����$i�M%�ࣉ��P������z�l�b ��N�r�It�oMm#Lvr�5����x`0��[��`�o�MFh�]���Xq�٘ ��2Q�O���L��"�7CM�/V`�:u*�r��.�&�Zڝ�v�sY[+��D�B<p���*�Gjy���S۳��{�j�mQEa�n����_�߭vp��KBԒ�@l�ܨ$	^=��'f;V�Q�Pũ��r�f�K-`�������q�D��+Rvsd�D�FGT�@Q]x�ّ�3�L�!Cv;�޷�Ǝ}F�#v�1[N�*R��v��M��/!�&F�Kd�{$�!>��s9�u�׶��N��;F�M�l�j�g�����T�����
uşN;�*FCKE��&�}1�9�����9�52�M�+,��X��]հ��V��\n��"`7l�ܸD<8��MD:�o����)a���ՙ�ȳ��Y��Nn*ي��gdn>�pҰ���ZUp�}�s5e�B.���) 7�gTj9Zo�&�oH�����3�������ζǳ���}��b@��u�C�wKz�D2�����%Z�p$�ULL�͗�{��3�ؔON �՞�7�1g�IBȳ"�9�̭�l��*�,��������3m���'�q�L�?�v��{��
�$%ԏ��EDZ��7�Xk�X�IA-	D������yt�we�7K�����ޙ�Xo��r��o�����6!|ǵ_ؗݕ���E�Z��s%E��"�F4�M�Ѯ�#��l�*���VV)27d(�S���NQ�2V���^]�19`��r�}6��<�6��N����	�T)FB�5����%P���-�}�׀F={�Hu=�Du�n��� q��$�s�;J�k��$wp�¶/4J8w(HG�x�!�%F��S"�]�һ�ڿk�����'��E�/7o���6�ߟ��&��ʔ�|���d�A���;�W�&��V�����^��ESpSP>�B�{�tK7��*z�oB.y?�R�#VȈ%�G��q9�}��
�vF��H����R=�/::7�������Ɛ;�2��غ�K4�m�jTk6р�]^2�j����ҢF��	�A�Z�7�X;�M���z�;��S�ǧ79�5���k���%ո:]/9M�&��w}�V9�ݮ$0ι]Q�N�aj�⻕Ց㓧(��꯾����z.�m_s�H|�Zէȑ��WA̵�<n��+��
��jc*�D9/���td�gs�n0��^��:_�}I���zU?��*SJ�r�}>l���R�M�������]���-��BB��4���,������d�g�Ls���\�=�4�S� �;��4n�׌���r�߱�mS'�'�i���{ݹ u�� scr����]�f�̞�}�QQ���nz�{V�ER�~��NmEҧN&P5�DŠ���5��(��N�&G:U c;4�M�*ucg��fs�2�[+�d����[����s4f�sC�-� ��J�ʭ.�8��'�e+&A;X���B���ͫu���9�n_C���ފj$)�Jr�ӭg��	AQώ5���'�|�L�W��pN��wݱ��D�����Y��9N#�ٚӹ���&�#Vyk%,R�s�yK�u������ᵓ&g\>���Z�74�!���(�Mq�K��(��X^��nk�y��\�� �kf]��N'���ͬ;��̺=�Q����Z�k���*Xql�ʷ�w�H��渙f��ǲU����ZS���.�d+�n��(<|�f��w����U_W���Xa2�;b�S��ÍA��d�Zɞ�bn��}um��hɁ������3۷��uv�OM�8�[�����B�u�L����u5��Óf3a�w��8vM=젧�L��o��\�#w/��'� �u���5hy���Y{u������6kwI�Ѿ݄=�\Ĵ����}���<���}P9��!�u)�zVc�OX��k��tRt�}����rͼ�p:�W�F����[�����7bC����p�*"#���-L��}`�j݊�&tX��h�>Y#�\O7��l[��q��9 �s����.��C1��x��9P�.$T�����g;t�LVG������c�q�r�Y���x��r���=|t�F��v8�fvD�9w$\dm���k)����;A�'������}��H�tWm��N�V�Ʒ�a�*�����ṛW@昖f���R����ڹ(9py����=2�����gp�2cӲsk����X�^�6��8��wTԮB{*�����q-'
g���Xn�K��D���`=^�����ǂ��*1Gn�姙���y��I�1Z��}�a^ֵzp���}9�\�z��iu�s��sye����~��{���畣T�VR>�=��g����Mo��Q���2����}�w5����#K�4y�\�X-Zu�I�N�(��s���P��NJ�q�-a�fK�ς�q�>�>�,�6�l$��%,6 @�8��z��Vǐ/}K[f�˶�A�w=V�_���P�]��d`����<Y��>�[~��c�I%�
���Cg�]���P7sI/y;�(��b�9sՀU��v����>��;$|򔾐d�k'`ÚǺ��F��Q���n@v7W� ��pH%�v�q����.�Ou'��n�����+4-BQþ�@�o��Q���V�!����y��>������v3�ᎦfY�*���aˏ0'pWlFm��y�W��o��W{�l
��h������p�(�*�ܖ�Y�o�ӕta/�R��Xu3�����k�Qw�z���32�������h�B.7@��zX=���ܛ�PHu�붘�l�m.����tpR/'}��KUpn�����dP�b��^�*��Z]}K{��������<�]q��֟�k�.yG#��t��@.s6�oF������7GI�_�L&���.��]� �06y`:��.�R�"Dpg�����U��;�����-��b|7��m�zz�c�cx�����Y��O�v�4t��g�篶�������<�Y#]�:F����H����u�ځ{���r=���˛U�׎&Q,��^��[,�K�h:Q�����b��L��v�E=��7>kҲ�V��,zmKQ:�N͕��c'��)�=�#w���~�P�������ڰZ+V��l�76��Ӳ[s��qm�]��C�t���3��KhqϬ9 C��בF���p)4�'0����3Kl��;���Li{��B��ɵC�U��y���Byy���g��-OM�8�Q��]ƴvր�{^u�yNF�-�'�~[L���3����
y[���b�F�]�-`�	��Zњ�T���J���)��B1�;^������d��c�������}4���ܩ�:��Kw�c�d�ЌC8woV�nt[�'瓛ue6��Ҭ��u�4a��y9�T	l���{��Q���+c��T�܈Ps�L����dh�����a�:�-)�� �{wڛ�xzMV7�ߘg�Uz;�lJ��jdr�1�b�9v�Κ͌��|'��q�L��v�{����d�ף���^�e��lE�e^7�9�w�7��y"�7.9G#�>������]jkv�R�Xu�^�ʮ)�fs�Y�Q�͛i��j=�p��b�ݦ2���e��ȶԲ5Y;T�&E�Y>����/���=@�:9F�Y%jjɳu!��$˴#��s!�8I�^M�O�K���c���bF�e�l[����-w�ƖD��{��j�W:��.��(�S^�­RFbY��1%&ŕ-���r��ǁ���H���tcV�E-���֮5;�:f�O�P+̬v�N>�42���<�L�t��/4��s�Õ�χ��H��;P*םN�θ1,:@��nS�v��46F�B��lMO��Z�T�B�V�K�7��r�%u�"Sh�!�y���)�C��J.��g\������="��̇��:�&襪��rnۡ��_X8�v��O�o!9E�no���d�3�n�8��/�V7]�(J��mZ|�:0��G���y�Z7��;h��;�i��Sv�@E]>,�.h����v�b���V�V��|��7k�nR�����v�U�V�J��4�R��|�x4&T(q"��/�U�aM�jb��J��ݷ\��t�J5�ݺ�@ʬ&�������t�rzo<yD�Y�B�g*�SŹ0#���!�9�>z+m
]Q�.	��m�лZ�y׺��R�N�g&��^�b��ܣW��I�wS�>�p�ۏV��V�X*<��s!}���^h�ls��T��hm�H�Vch��N�W��2��h]%[����g��m�L��b�*�D0?�ܻ�t;�饶�L��+k���#x(7zd����O�9��:5�S!{�����Ng6�|�H�`���q������@��]�w/
�X��c��`�7R�r�RDˉJ��xR-B~����߈bQe��U��Ε���[dLj�X�j\�����[V��Ù}�\��em�C�7��9x�0+��[���{�^St�(m��!Su�3�$�S䤕�mط1�Z���>��'ѧ]�y֜�;��[;��\i�2:,�.� 觺�֎x�Q��#X/�T�Ι'"u"w܊��Wt���]P,Z�glǻnj�/�L�WR�5;90���&L�t܇b�k�2���ĭh���NE��ں���<ˮ�\�_Z�	Z0���A5.�]Y�h�u𹘶u�����m��g:U!̻KV�k�]2�����}����@]�W>LPSFۀԩ8mm��n�]�U����qI�}��DnA�;�һ��96 ���sj����'V�9�l6����wr�e�{��K�n�[���^������ ���ݺCyv�Gb����/^]����*[��cr��nD�w�׸���0H
���}�m����b����դ��nĲS=�3dڷ�L��4�>�R�A�WP6evbҳ�-v<K:܏�{��9�]�sv�˟a�x�MKfn�X7�c���-�u�[�
��%�S�����rn���2��NW)�vnqv�_4��Dh�y}+z�IS���J�5ÝwQ��)�c�Ge���)��PafWZƈC[aFF^]��Hȅ��κ}s�Jn�e`����r^�����)m,�������]m�XZ�Q=3#���s��k� �eѧi�s���8������;U-졆j�vV�:� ����t�Q?cwYر74�(���1W�)�T��bA[����ځ�X�@�ʽ�P��Z�]N��@���4SD��n���Yf�E"i��URFU[C��Q��b&�"�bYr+5���f9��!zh�f(X��N�p�c���	)���\Ԏu�'*2-0�Vs����UPS�C9D�a��T43�V�]+ �	�<�y�A�bAA]*XH��l-R���w/K4��%B����+B��q�z���aJ�D�hȊ���z�%I`��܌Q)G$n��"�t��2�L4�V��!�-d�T4��B�h��t�<�r1:U�U!e���+�	f����#��=HjT�"!,�T�J�3K6�mD*��f%��C���	�X�X�U��̒#D02�M3�T��hd��ʢ.\����FTd�2	EhXJ%ԐCAf��L�P���3�-CT�͖���*��˗Q235�mjj���Z�Q(��,�D�W,�IT�D2 �V��b��9ffr��0�Y]:.g@� �m��dy��-�c��Am�ۭl5P�ʜ��,<���}7��F�iD�:�hΥ;U7�ۦ�����ڼ�%�g�����(�Y�j#n�k�9I&�ml����j�az�`T=٘����EP����ɋY:��}��^�Z��b
Ojp�x�̦e��2.�K��4�CƷ�.a�驳�o=�ɷ��R��:\��$]U�=�6�D���U@-�w���D���Z^���L������i�>��[��ƻ�^T�ҽ�qòvb�:κx#�_��k�}G��tc�Ez��g�ʚӽ<�wE���yANl�;Y9 .����jWO�OL7F�=�a�r�/6;[י�}3���(c�E=�)�v��`.�铻��/g$CVrl�N`���2sb|�ۯo[�b�}M�k���n�:	VVs�6��Z��"��͒阃���+sBDӪÖ�f<�Oh!l�9x�6��iQ��[`���I�ӆ22���}gFiD�t��)/�+i�e�h��,�����
ɶ�xS*qQW�=�Cݝ��ޕ���:��&ю��ʓ��/�T��B�[�*�O7{(�r��M����i��Eݝ"'�QǦf�O�NF�ψZ{��ιf�=THL3i�o��AEx1 z8�T�;��������E4^Z�2:�
\lzN�܊m�����y�/*}b*�	w�����g4T�Ѐ64��9+�ɠ�.&�^D��ϼ��c�x��E�u���ksԛ�m�c���H��]�˸ۻ���Fӣ���)�'$A�Qz��{�?W�C�$s��t�q��k�M���C���-k��}����;��͙�,�skHY�8�Q��2|��̉���w#Bىx0/�#nʐ���va=�1[���W���j���;5<�魞�>��Ʋ:����j�Z�ܧPo*W`�v�	ӎvI�Y�V.�>Ҙ�e-95�DԦ�I��{����j�9����i�Wj�����R�p��}�4oq?T=�׶6~�.P��ݼ�Ua����{�9�6�͵ L��'t�9Oz�27^)-q��^��[>��.���.�2̼|1
��ԊxU�߸�k����i�4�Z�v����Mi�hF�r5a�aڏ�����m��g'G] =��#�w=(<����#������1j�����)hfa��� �|����_m�@;���oR�����2Y�֨��}���31)U��,��^��dd�ʘ�E,�b�����<���'u���P<��kR��i���ז��]���t���'˹�v�o�������twL
F	�;��1}y�]ޘ:�3Ϡ�ob��|�m.�=�+��N�vW] ���f+����󔅮��2�>�^��z�O%\��=����W�Y{4M0����ݢ��ݙ�� r=��bv{s/�{ڴR�1�}r׫q�K3�3S���кe��}cg�H+\����f6�`��	K���6k.����JxH��U��:ӫ<�a{�\�h�.M*�E�ɺMs��Mx�[ѯ�%���l,�k��c�A,$�ʲ�[���N�f���{m)��-��~���ߩ�^3���\�^�,��E��^ә�@�A�?]R������LS�1�n�y�˝u�K�^/�������VW�\)��r%�~p��
�Q�T�}tVd���C:��e�pČ�t.��+ή��*}Te�u�h�[s�.QB�1L�F�7�}����*��Vr�i��u��p�f-}N����.Vh�!����T,����L���P��Ts��_������ez����^��e�䲢*w��������a?\hu>���nL�.x}�	��3��{_C]�׹MD�=d�j���Y+--�7E���Fv�2�i�u�����g���x�Q��4���]���]VI;͛^�t�X$���F2m�fWCm�:򂜍�[݆u��5R���e���O3�ɀ�}�&p%ul>��;$|�I�Dn��3��
���۹���c���.����ڔ�'�U׵28�X�r	�'R�z��S�nC��ho����=��.��݂�#i�K��z�&Ѻ�k"je��-y!yM�����v>}�p����x��|ʙ�V��'�OZJ\�O_��W�<ٹp��6t�/L�K���Y���_Ov�z2.��i���'{_P-�t]q��X����,{ `�niɹݫ����/���Z��J�5;�eq�LD���Ǵ��Ba�۩��pYʊ��7W|�j�<�̣Z����%�$N�9p-�`�����t٦7���ݴf��E%9���5�͑p����a��r��j�i����r��EGC|�f��؊�;�ՙ�<�7b`��效��l����&�Ni�����P)�@X�B�{}��o��G��y��C�<�Y<��\������^��Z��Nvy�v$��e��O}�Y�jћ�Kio?I9sZ�^߾y~��Os�=5{�J��T�]�彌�������gҒ���_`�_�\�ͅʓ�'!3�e����`�����
�}��.��O�F�}im& ������.	/�a>w���a��*{͛s��]���T�xH��^7ӷK�xf�G���ݺ�6�	^z�4�Q�.���{����������teu��wy���nl��C�2Уg͒X�l��O�JYl�-�|+5)���i�-O�z�.B�v��oD}��}G�r�g�lj耛i�;�ǻ��"�\��W���sj�nN�v[<�L�%l�7J-<@�����p���a� �M�|�y�K}z6�+(��]����I\{��9�}� ��t�>>㽨V�sW�c˲�`m��Z���ʚޜ�}�M�RKYZʵt��Թh)\w��}�K��;���������E��I��
QWJ��������j��b�aVQ��Õ�L�W�1z}9�ݵ{r}���o��"�O�oOf������/bBon����r٧��A�Ѿ�sH'.D9���w�Oq��:3�u���l����M�P.����l�8j�p������鬝�:����9��:��F��'J%��E���Q+ZUD�El�h�"�|��-b���t6ٜq��O�N�n�q�N�"F�P$J��jɘ�9O��u�7��vu�N�W�5l�5����'2B쭍l@'#�y��uY��a޳͌c��:F7��5���j;-a�e�V3��[[qxn�V�T�1��%Ya�U�)x���؞����u����z��í��T�mܩX�^�J}�6���q6�l�FO�\���x������8#۴����{��o<��:�O��<�tĥ�an���+�07uՇ��f���_o+���[;7�����G�)ɫN���N���n5�&�2u�a�m�	�&0�p�v��R�N=�;���%z���ש��rQ%��ø�:z���>���G厭{��2���?��2��m��Q\Ղnt��g�w�����v�(��蜿̐zY(C�������\W���{U3��]v���+��_����J���~�r���%���]P
͘q�2x>�Lq�8�/�XJ�o�ީ"��}�/}�\��yT'���~���Lg�8��{�������������<���[NZ�bM�w�Ĺ򺺦�:���K��c�S�����P��:�s甥�&k���m䍾�=y�۞��n��P����V�ԅ&ND�U׵Z;m��%�k� �b�ðm7�8�]���`ɸ~�p@��85�#6Y���c+n��V�^�z�{Q�U8X��r��F��'�����K�j�l��3[��;]��,��~.�χ7b@r����8PElKl�̅E\�Z(��S�n�>⹼�{�$��7��tˣ� tq��Y>'}Z׺�^Px: ����_�ͫ�WPmG7�6��y�s;gz+����n���Z(�lԌ�f8!��y�EY��J�P;��[T�_n����Ž]���^M����<���;`hc�
=�U����[�ѓ������uigv�ʟ�ﾪ���6jn�Ɍ������

Y-��%<$�z_��:ڨ(�=�5s|�\��F�z��M#T�y���>�ǻۛ\�]�9��|5ܝ�S4<��α��b�s�/զ�,��ZSj��l�~���k����c!S�2�����W7�
�o�R��)n�AR�l���~�鷜�S��OXĦ�i���s��t���~��r�v����&�y�储~�(]�<o>"˻�|N�Ѵ�rVݲ��P'*p�d5�SQ!l���8չq��{�����sۍ,�Y�c1c6�����l��dI�w�j�=���RKk�a�������S���w��﫸�7�#������oiμ�8"������Yy"�lŨ�'X[�Z�쌙q�'�{u��#��s�q��F/�|zi:��W�����o���^�]۳	�wb���޺c���C&��c[�2�L .���"��:���u=ȁ�|=#�=.�ѭV��3j�4g&�+�2^����;6���a�.<9VvT��{�S*:�ĒS�)���v�&>w���_i8�K&���/zıI6\��#`��3��gt�7����^�d��Q�F���Rײ	Ǘ�m��>%>{&�Nj�,X�9 �]����u��~Ⱦt]���/$Sf�����c�݆nxo%&n6��M������M㷻�>��wX.�����.�C�'	T];ck�6ntJ�'C�F�X�Յ�,ִd��Y-tY����W\��S�L�)b����>s/Rj�T��qĊ�܌�v�sof$k�]ط�K��E�-��v�^p��Q��[�t{.�\�ȼ�u���æj	�܁��}�-�Y���pc��G����j��Kb�$����9Ӄ=/�~�ܻ{hlX[03�\��t�k����-�t9�κU#�4�A���S�!	���37A5���ͅ)l��^1+RmF��{��ă��-��!V�G`�QK��Y��[�|f8� ��u{�.��K�=�}��lע����p��\o֯3.��U���-Z�=��bx4�C���)[�3NY���Y���o�����"�y3M��u9B���jt���(WR-_v�����`W�ۙJ��2�P.���	�B�wm���D{�v�Sⳗ7ջ��ԉ�:��B)Hn���X�9vrb��y����I,���/���ʟ4El.�l�=S{FV����d繀���7<jQ}t<\R3�zP�﷮M��|4Уg�%��턞l��a��+j��IH9r	w펺 �ݴ'��f܂��$��Tnc^*sVda���z]z�{A�<��6A��7���A��ޒ�uh\,��0`���L�p
M���,�L�W�1��-9BI���߽0u[���7{/�����<�V�sΜ���on�޷�x���f��t�d��s&���Ox�������ů����A7�@�����f�6��nY'|�/��mt��Z�+ws��zy��:E���}�[��%ڄOXU�	�؊ͼ���x��~�v%�.-m��ᆂ�q3�����~��b��c?#����C�ņ�=�@�� o�ɵ�q5:��KB�	ӂxє�dGh��R�!���r���-�u��o�+�7�ή(�:^>F��#��*��;:Mh/wSWr�9�������O�6�9�e/��G��{I	6v_�e2�U�ɹY���ٵ�Zkx1��o=rj���`KD�
7����L�e3ë��#Ozq��9��K"�"`WGը���wh�*
N ��=xh���'��!k�9泑tê�N��Jh�]�wƐ�6�6xܷ�!f���1���v2��D��ڊ�L��s��������*o��P�\2��@>5u�z�
�U�6h�f�o,�iv-�H�]b��0�0��1bɛ;�zY�B�,t�5|ź�{�����Ϯ�L!�{R�
Ķ�#mj���F�y�pѤ"(�W�gMl{Rb��v:��Պ���Sp����V�=�	���k��U�-�{�]��m�8_R'0KVBw����n|�Ya�N�%o[�S�������.�5��k/�����"���䑵�]�5�"!&�v�֔ʣf��S��Ͳ���q�Os��S��r�,oX:\;�&�t�뵌ܻ�A���r�wqS��0�5���ӭ?e�
��/�us��V���W���i���}Yc��$F	鷂�KI}rC���:� N�xQF���5����%�e��Q�"�·c
O�r&�掺-��.�η5���9(Vd�1}��΍԰��w��ݗFt{�ң;A���
P-1on��9��*ӎ[W.Jp?u��U�(rǵ�U��͗rgs츌=;86÷�a�Q�����';�.��e˫}���ޭu�6��6�L�V�Z$���\��vr��H+G8J.�&�)�G��3G6��[�32Q3 �8�r!͎����#���b�gWS�B��J�ϯ�W6�^1��֞�\�.��+~�;:ew�.�I��RɎ^��]n��U�G[n�<�(�*��J7YX���:��E%��et��/����j�..��� y�d����T��<֮w45�V�7��]Y7�Sh6�͔lX-_fF�8N���\�-��b��ǬֶX�|�g4���C^0�x=�u��Iܴ�K�9�j�PE2$���D�1���2:ëk+^=��&s���)�I=��K���
��ѷ�΀�k(����[x�wS [	�}z���Y��{���
���W�gRJi���\�](R��9{Y��Rh��S��(��Y]l㠗�YϩG�(�_W`�-����n:ZGϬ��on��a��2����Z��PI���í�lX���/�U�'*�4���u,2z]KHM�4�u0m���}�ˌUq��YnJt��N��%����Zͫ�^=��-�g:�}v�cܻ�u�uG���������.���C�oTj�6�=��b���*�S6�ӫ3O��T��d�b��]��m>��u��mV�-�p��6��l���� |Q)DM�a�$ȅ
Ӭ�PI��$��9X�JZ�*�(�$�aRY�����+����G+-�j�]5.����SS2��* � �9PFb��aTjTr*�Za��4ÅUem0Ԉ����##CK�������UZ$,�ִ����
6���!QR3.Uf�UZfr8�*UB�R��K5�VfR��H��[hQT+��4��K�BE�Q�Q$�YR��Bh�e�dTgP"��!TA	���9r1jHY��Q��p��!&�p��*��R�%)J�B�B$6�I%t��IJM.f]!20B¹W9
"ZkB�AD�2�M�H�):)VBduH����P��Qa�eAZ!]E���Y�U��r̊� V^��:!gxou=A���}��#H21�2����=�17qz8��h[W���	+:���kH�s���)8
7��UUU�5Sχ������J�b}׬Ďlc��*F;F=�v����=�ڗq�mה=�����ݾ���'�f�1*v��&Q,����W3�T*}��~�ޱ.����[�����ݵ���J���֯�������W���y�ޗ%1e��oو7�b���.bz���	�xݵO�5Yî��臇]�V��
t{�r0�Fj1Z�Yi�,�Ț�o�-kӖT;�!�gK�x�����8��.�5�k���E4<��(q�o��T��ܔ��c=v��r��J��!m�Z�ג�Yl�-�;�^F���ɜ{y�ʰ�!z=�9J���[�zZ�:��z�6g}t9���R���KdO�38�!��y�#7��~=�"l������"��&F��i�KV<"��H�S4|�^^�%;u�}S�j���xgD�mHRd�9*��Z;m��8Z��$�I�ٞ{���{ugK��evzޘ��^�Hm����r'T&�#��q�Z��0u��
[�Fׅ����ٴ�B�_���f��+�Z�0"�7x.δ)�_s�3�+m)���Ƹ�]/��ŭ�w��/�����a�t	�古��ʮ���fՋ7bMIE��P������Xy�ǖ������k+D��Q�a�666�m�Fopd�M�9�>����.���:q�N<�:��Fi�2iE܈5:����]��S�μ]cw����v%�P9��0�\�XY& V�\��ș�⅝��ڤ�i�Z2t�f)k��N���A��e����hV%w'��!N�$Ơ�����V���%���SĲI���~�p_Ĥ@ǽ=�y�Y��eK3�@;w^�K"�N�D��f6��I�ѷ
Q���1�p���Pu�O2��߭(<����I�5��vzdr�u�&�b>|f����|���T�V��Z���)�]f���"cg�q��|�[�r��F�Pn�Z��#%}y,ʈ�������nS�x�(�+��R�v�s6	��|M�Z(�Tb
N��iGv���H[=ih�9J��xǫ���0��Ew��Ӯ��<$�ʇ+2}���U�H;�L�9��7�.��u�^ط���u�Q<�)�����t��^�m�>N��Վ.�"������z)L\�����x�Vs����{z���a7�)ѬV���dFa��T�_�}_xco�ފΝzr>��0=����^�$��)e1�̦*̵�$]n]�1ɕt������L*���g$�8�e�s���tm�yμ�/bmWM��;���{y��qX��T�Gu�7���>��H�^�u��}��3����fw4i�k���wY;�p@��v�ڔ��݉���UaU ���ܣz�3w���z��
znz;�;�{ap@�3���fͰ�͉/-	"�&N1ݕV&�f,�nӛ[���i'��#�9��배^!�s���LE�ݡ�6wu�$��&�]�I�BC�:�eda4wEڬP�hD�S�L���앫,��ִf�]����uǃ�Ff�_'�����e1I�m��Bx⣶�7y��9���{�ls-�"�lޣ�Ox抑R�*���yV9����9�V�<O����l\���pح(�*����c��|����m٠��t����Nq(m���F�T*�5f�\�,���l�@Cֺ� �O�Z����������8�=�6��*�>W�c(j�Q�D.�'2���P�_`�nmv
K�����Y[2�n1't�=�������v{�m��ё�m�t9Dt�{Y� �����'�&j�۽Qtai:j�YQ�۫.�M�[���H�(sɝt�q��=-k�%�as��b��\�c;����r2�]�yC[����y}�E�M�}�;n����q�]]��k��� �3u�� ]=|�㣞v�9̧��KHVk�������,�p,���`�<75�(�������7�i���lp�E̩�2����T�����A����ەaD�^N��_Ql��+�
h�wR��幵:$oq?C��/v���Z��	��~el��ޒ+�]x���Ε�A�n�t��}U�m�9������� ��2e��k��=���.�m���7���a��s�{�AOt�'cC��ԟdM�T�M���zѸ��/:�c��dό��F�/tT�I�|}G+�H�N�<O7R��&U�zپu+��3�iȗVp��T]@��V-�%Jަ,��V��m,ފ�(u����7��+�-,�SaX�-�gr��9��!�z�2P"�<Mm��֦��f�H�gfYiW�+Zs!W�����)&¶ﰰ�̼���3x��Z�!U{���#Y,zl����Y[.��F���j>LQ��b^����B׾9n�w�5d�Wdf��y�(�ˍU�Q57j����`�i�݉Z�r9 ���Z�o�z9;���F������Ԧ�,/Q�ؖޗ^-ۯ���� �.$-��$�kƵ�#�4kn�w0��Df�x^)6*��C�i|j8I�KCn�g(�i/��)�of+�l3f��3�i�IE�O����A�Z���D���b��8wBJ'��ޫJ�������a��vz~�C^z.�jo~a#�s��@΃
b�H�n�5]")�f������Ҝm�����iF�v�����Ǚ��$�=+�Q��,� �VyD�`�*�E(���,����s5ٹ{�v�H7�!��/���%�(��2k�w��3FeJ�g�^ס��H�YLy��=MO?[�;y���6�X��h�I�#o�
�Nq0o�"&e^��KӢ�J��e�zVvF%>��XFŗ�����;y\wtDWR�ü/�6�>���S�N�u����Z]y����S�e�&v�1`�2�y�R�)e���ҔA��x'����e2�����t��n�,���5�	=F�������t2��KÕX�J�`#�%ޗ�z90ϲdl��ve�J�2Wi����m�j��P�^D������d��]`r�/`'ݴ6�9��]��o��a:��k����T�3rz"���[��8�+<��u�ů����xF����,4��{��(�Jn-޸z5�g��k~��3낟�U���ߐ}�K�5��hh�⩹���N���5N�W>R�1cWs�v�c�+���&�K�q��O�&�3�:x��k�9�.�uǃ�}7�����M��hI����m���ۓ.�-H�ל�o"��f|����oR����PT#���R���,�?!��r��K'�D�R�<k�ۛ\�]�9�����!d�h$4�w�����Ƥ�.�[��]����xرva���/q���W�0�&o,z�D�1���8�j�pu�0v]�FR8\�yG�E��TAp�M،��o\}��bht4,.�������_�^�i������O-�bQ���˞u�/�ݭ*vl���;�w�����Bv:�z���������yn�6�R݋���^Qm������U<�����t.���=b3���I\���}�0�H��%(���-+db��eDT��T��f�-���8�G��av�SCz�� ���:U�ymd���/vn�7\�W�8z���&z�G��m�B�Qҟ=����R��̯r�5�V�G)����i؛���5�2�[9%�?1��u�:#^��9ҹ\
��>�ͻ��-ߨ�]����h�9��}��;��,{�.Φ��핹�A>�ftm��e�o[��N��+ǂ/6}u�ڔ��"�q�W6���G=�wt_������V�d�{}���=���`[5�����wT����3���9��V�P�}���גԓܨ0�\�FV���U�8�7B�k�r�*��w�����L?uȮWnF;��8n�m��d��	Ej	ӊ���%٤q%&�:^����k��"$�Զ�c��w�����#f@w�z� �F�0s+�+��#��׷+����N�Ym�g��M��S�>3z����V߸?z�ݦ^uXh���)=ϔ!V��#f"�
�\����}Xԡ�0G# � ����y�\o��$\�kkzv㳅�MP�{B,��8�[d�En�8��qF�o�*m�.k�<��5mY�����k;.ܴlOW��9����#��:��~*�	��f��L�F|K�˦痻%w�OƹD{#E�9r�N���ic*.,�V�x�{���]�Q�ҧk�(�+����ݧ���s,�-}/<�54nߏ<��z�Աw���xf7#.\�C���ml���˃2&H��w��AB$�q[�D��Tc��|n�x]=|����ms��h�Ǽ��%��+ٺ]�w~����Ëo=�P��:^���p���:����F�G�����[�}E�ϼ��C߷�2��r�ǯe{�龐���(N��Ռ�ָ���iB�h�Q��&,��3��ϯ�[���/�F�ʷ!�k���GL�uU����<�;����<��}bZ�[�n�I�	�}�2�*B��NY�c0��"9�άᎺ(��k ���P�P�Y}X6��Ņkw�Ӣ�p�d���6G�b/��يK�gwe�oi�ܾ���k$N�] W���IY�z��ź�FM������ͽq���r6N��9\*�Hӓt� ���A�ۄ���sg��z��7���0�i�������L�U��A�r��y��s�����v�	��:�~|�`J�4�Zj�I��X� ���њWg�]��2��}z��N<��5�3g�el���Wo����;�c��]��:��,Aq�%u�<���֟.��gq3U��K�ܴ�d�;]�7C��܎A[����F�ngj�Z��ɢ�3}��,��v�}�syj�K%�'�-uN���9q�〹7;���MdE쑖����s&�܊e�%�
IlF6�O&^�ާ�/'[�^��1��xuyΐ�L�jUMN��r[�%A��	�,1׽n� ����X�yHvBP^������'���V��2��i+���
ӕei��#,�6:�g�{��e�/6�=�t���܊�̢38�Lo=H�Vd3vK��v��·�+�P���k$�F�E�Yr쮮�YcMң�!#
��ۤ�':u1dz��V���Jny-��̷�ֵx�����W���vہ&vr3���-ȱʖ=zn�U�"�O�m��^��z�eH|���K4�{�(r�e�G!��յ\�O��T�x��]P_G���哂�}�m�9	����v헧-K �N������j�Y=qh�a���y����VӎSl[f׬&�r�N��JY^3���h���3L8�L�}m�3z���F�දYRi�$�E���ImyJ�a��7�8VӍ�q�-��Z��d��;�D-�ɕ�6v_7[�l7t-��T���{W�U7�OM���\��r���}�[R�9J�DI \>ͻ�
�7[�S6p�znGGt�(g�B�n��_p���Uk8��q�cGgd;������.����g�r�z�ڀ,��l��!���#��(+7�L��㥊̷V���ca�rs��u���},���:��j�E��]o4���l�b�4��d����	��5!��W�7�L��7j�����h�r
-u��U�a�ĭppcTH�%��F�u4)mJ�.�>���#�jV[�4M�ؗw#���ui�dr�'�$�����}�#=��f��#Q.��*ˎ�9�",�£�q�����BK=+Wdݾ9�J�o���0q�;&���2�r��}�*T�̎�.�:k^3�RR���p��b�@Y�[T��J�e��fFh|*9U$�%�PbZ�%�eoXͥ�x�♁)�����;2�>��/��6�	�K4�֓q��Ĉ1k������x�}|r�r�=�aé"5.��SY�J���u��_fv�VE���g�7* ]�i�۲f�u�r7O����/kL[�`�֥so(�]bpyD�yΒc�(����{ �v��LQoܶ��I�d���V�}X�7�H�31m�hj�,SgK2tgT�}��js�F�\[� �c�/J��v]��p�f�Oa�$���C���+�]y�g���	Ѯw��9n�z-و�)��Z!
���cn���*V.��[B�.7Z��x�J�a�̨RԨK���C���!�����a�,���+�ZS�����8�3GE*�wf�r��u#��NK�gCVi��Gb��O,��MFɴ���AD�G�q�X�j��=�Q)i��$_Hjf�����:�!��s�.�\-8��Լ�X3lv췕��9
T����ChJ�s���(�,��{�ou̱��� �sH.3����dd�Hl��y%��E%�m�{��]+�.�)^
Y[[;��U1\�ي�꺉Y�ݖ�c��\���������._KH>�oD��&��f���i^2X�֌��%�Jt��k
��g�����ɥ�sk�?a��]��D���2��,ǩe=��2X�އ�w�J��= $ �X�ӎ��4y�!&���/�r`%��-=N��wx��̮s3�b3e^CY&�+��V�	%��&1QiK.�j���-�v�g*�mNJ�P�mh�P�ٗu�f6*	c��*�piࢻ���{0��v���r��y�`����<�p��th&V�62�ͮ�]����q��y�4+���˯~@w!oX���Z�������D0��3����G[��NԦ�7w�5�A��lɁ<��`���m2�0>N��n�� +,wwS�=�ƧG���.�Ț��
�"�����͑2vR��gy�SV�ܘ��3(�CL�}�eD������ei�z��珜�NSw:���4������x���(j/���Ð�<�Z	J��dr�هq�'�`�<v����[��oN�Л&�h�mQ�X�Ѥk���w-�J�}|݁\%���n�2>\ J���鮇u�/*�I6wϻ7-��B��׷�L4L����,$H� Ȃ�j�J�)�JYE)5��YJY�9Z!�u* ����T�	V%�Ĭ�*�.���.��H�Ȋ1Y\%�Q
I�GCM*ŉ��4e$�L��±hM1AC
�f)����D��"(�(�"Ĵ��0�5R-����5 ������V�T2�-�d�.D�fM:t�*��U2�(�)g*5�*p��%TDa)���B�KQ9e�r�T6T��:,MTH����fːf"��difQVeY�˚�Q���R#22MZl.�6*a�E�UIA�"��A�s�Ш(�TQdV�̎ȫ:d%DZ�+���[MQڅ�(�CeQB�-D��e��S��QEU�RA$�,L�3dDQH���,��$D�r�*���
�ʊ�2�Ul*�T%�bu�BrQ#@��׏?�x���y:c���c�/����
k�f:�W����c\^�V���pmW#:ȵA1'T�����W}��͊�3��2�NF�'j�#6}krt�i�Vl���U��!�{`�����m%@���Y�B����NB}=�4�O��09�.�uǠ���.��r��m�wj3��v�s/R�O��c&��qQ��^k�3�r��N�f[b�F��Ų�gGM<�Oz�^p���yO���_�4���5�x�����K��c�6�W=���O=�����h��v 5�/l��=�o�w�(
{=y[{�☉C�����^��f�o����ы�z���/�k>�2��Z5�:���\k�tC�ޣkdd���TEKkU9��khL���ۼS�1��_�2|a��Z���lߵ�5�o}[�a�Sfx?Rv
�đۣ;�e�P����b�[�`�V��JN��^c;�P��dV����̗0v�V1}KdN��:'˞�p�ъ6}K��΋�[�{��~���+�Aɧ�d$�^�R`�����}eSƅ��2�+�������	�Z�m	��v/����٣�kogP޽د�c�t��uף��+�K;q�9}Q�:Aw�#k�Y��t�n��n5�wC�z���;}W��TH�u�Y�f�WwtR��!��.A=����5�F@��"{*Ú�� rɓ��	��������Vb2yއ�V�9���h�Q��y����)Lp������O����O{��}�lvS����d�{|� ]�ʹ3��nMA�p�r�h�����PV��[��^H���q��B#h�O+��s�e���˲;������E�ޭ�`Q4��vdsf��)�C����������D��F��7`�:�(�ז9t
�W>�o��������ͻ����Ů��9:X�k+���ڱ=L�?f������~��n-�e���V:���Q������űn�z�t�n�Z亀�.j5�r�O� U�Q��Q�[t��Z���(�KF%�U��R�B7�X��zu��/��hO���Mx��^s���ه'�%Fk1��%��9��:U#�$b���2��aڥjȮ�ҩ��`���jȫQ�����xK��Cl���{��i�:kѮG�,�~���]������Y���N}P��+0S�Ϲ&�����[Oj3m�|��S�J�;�
,�鸦�h��t�6l�����-wT��m)�P��#�)�̥;՜��M�l�M���^5;=?T�z`S�ma�oVl*M�9�=^�A�OIio�ݖ����r�T��KUx�, �Z@X�(-x��5�j3L�b�ɮ�H;U=ih�^��Ëo;��l�r��Dv���7��ܙ�/�7��fk����L��zk���l�����л�i�rڕ���ov�`R�29�yn��s����E�N��s����3@�,��^�5ΰ�*��i27^)-�)+)��6����Vl,0,�q��)�;sB�W��V<a#�;1S)ebdn�i�U
Z�d0eeif<|"z�U<N5��#w3��9���V{U��ؚ�^
�.d��L��-E��.c��'pj7l�f�Z5�R{Ŋ�-uV:�'�<���2�ӛ��ٶ�q=���+˻������"�+Ew�
9P2��(�{b\,�'c��4(ht��vѺcz:%�����|cޗZU{�M߽�{�=��#�QkE�?��W��6�r%݋�[��J�t㙮�kX�%Q��My����T3�-�J��gV��1.rU�ʎJ��͕�*� ���8��[��~��W�R��(Au�6ώ<
ؙ3cd�"n]j��ڤF�Z/N(LR�Tꓪg4 tq�9`���6!(����s��c\���˅�rY���-��m%<6Ž�*���5���2��]fr��{P���m�n�RȬÓ�l׉S�i�K�`4Z"Y�k�^����X���ZB�z�}Vy�ZPy7���<��x���˭Zϳ�}V��������O4���[u[!����7΅�5=���*���{{����ـ��.̄������tж����_Y7�^=Շ�Ϳ{+���l���nF���6j+V����)õ�{�0�����=ioÈ��1�1k�׺��ݝzr�&0=�\6E�fw��N[�����;���C��k3 ľ�/K��/V�UC���r����5���"g{އ�<޲���M����$V�4�X��n�sv��O/��q��D�
��:Ty���J��k��d!�0�/M�x���f�9E;kgK��j�A]�`�֞�O|�k01ݙX���'	;I'����[�������"��v�Z����}$a�q~�wo)>�V��ݜ�[#ggi���n�g��*}�y3=�xZ��m�̩빕C�y֙h�{jB�'#�1"�����j��=����e��kLrZ��ɂe��|�ωN�dPbpd*�!")�g	}�Sbh]�i��=Os���M������n�e.q�������޿}��U����n���:�&�����R{�G�r�rwX��)��|����_�}�>�z��76�d�{_���uǨ���B�2{-��"�ީ��4�ѓA<q>��ȡ��q�-���S��t���v�r$B��[�sEK7B�F��
�]B컫�y��6JM^F����w6(�[6�0�y�b[cr��v�g`�d�u��㟙��굗s:�{�'4A�z����c%ܫ���:T��;�E�ݓ4�؜M��}�4H�/a�E�e`��r9�{z>viF�2K���U�|�X��a��i�`
�0��JsS-�[W1��AY�܂��#nrbw%�hTK�	2�Z3$�ū'�E���\����^��&�]��i�tЍy]�':���J���M�6���:�w��|�Sd��fj�l��LbV�ڊ���*"�ͪ������1{>�]>[�7=V��a�&1��� ���Dsf��ms�����ǺM�c/{^��oz	\�p��;Kh*c�����r�էP0Rs�)e�8O�o������й�<�u��Z��k�ÙO�u��漵�>��r��[�]S�l;�͇Û3У{���|����n����}@�4}�Q�A��T�7����yu��g][��-��9��)͓'cx���{�z�E�;��wr�}���k��5Ԍ�����V&G*�vOo^�_s�j���^W��Nc5�<��1��׽��7�\=���o���i'��p�7�ӽ����,�����k@�xgص���>�{�o�����vsV�գz7z�FV��-���C�6��Ǒ�# �#��҉y�� �L3��"�̏5Ϸt��޸2�_}�6��	&���Eݿp�]�k�]���a��R��[�8��.�n�<������.�8�;spI�F%I��kw)���F��7�p����mE��Dm�qmw-��[�7t��C9H������s����[7���^�{�U��j=ɭ�Wp�Av8�6{r+w�p��H��r
�5����1�3cfl$��t��|:R�ĭ��{�l���/k��6�h��ٻؠ�.K�4z�����M�rʼ���^9�H��.���L��h�2�.�]�8ԛ� �۞�Y��/}酣��k�ov{E{Ue2�����[�="�!<m2��ͣ�E��5��F���o'���e͑�v`�ǣJt��Oۓ6���Oke�.z7���~[�'��.�S��z��:~w1i�������Aצ�P�8�0�ws�ƹ��V��5V�w���3O�u+�]̇!7�@P�H���E���x��Uu��k���0��j�w�M�;0�
Yq�(�vdR����s	(�l;R��ۖQz�i�8��l#e�4���m3��Þ��k)B�g{�GlAu�����M��Q�ݶ喜�h��� l���QMBn$v*ʽ�͔p,u n�r�/�%����/��+ˣ��Tݶ"�Ib�g���^g���6�e�o�f��Bwv�ƅ�\��cΨ�hݩY�.	��\��<WuE�S��f�ݲ�o^�Z���)��#P��/E�)�`έ/��V���Ϥ���nS��������PU�0�Rb�e`�
mf�����/��S�7 ��N�/��'xg��4�IB��� �D��j��׿o7J|·C.Tݳj[-�}|���h�A����4����HL;�R�ԩ^��K��Od�'��U��p�I�1��>��5�ұW��:5	��A������b;�<������4_i�)��ܜ�Mfc'���F�wN��M}�:!<c(��|C�����q^���/o�{,*j���M�U���-��Ԑ~��!�8�wV;�Ep�e"��B��z=V��C��`rm��yɋ����B�^�"[i�5� pLâ�eP$!��е;-k�85�|���c]�~�y��D�z�I�$��}����̆�)u	������K[#HB|nq�{�7��(� sP�9�1�g�a���V=�)��	𶪬t��uT�2ΗS�^Ҙ����xb%U��R���+�2���vL8���{�[O��ON`�5G&���r��֮]��N�q:ue�ڗ��8�.��nڷ�˲i���a�.-�
��u�k�-{	�:WU��ɋ
�0U������ժ�!ѹ��lCFU�UN�;���A���,[{��;����	M����f)�͸��y���{��]Έ]q�9�	r���1뱕�#����L�R�׉K�epQ�ʂ���@��*�ѝ�9�:��v�k^�fnasg�d�O����ǥ��T�ǷZw�qp��X���_FC��N`��ܧ굡�c�~Z`9�"9�}en�1+��Q��[t�����<������e�����B��b{�^�	iπ��Xh)�Ot_�D2z�'\☩\9��Op�Ti�m�V ڰ�Jݟr��x9�a؛��/`#�!=�8����+iK���GM:�����t'��{��V�+��<n/,����Ǭ����nW��ĝtU{����K�϶GK��b�}ú��[w��c�Ŝ��s07F���}�����\�=@ � fɞq�T%Ck�u��k�S�����#�Tͽ�r܃WQ�<ѹG���m�t��|d��Yt
���'ɀ[��C��%��Axj�R��֪�|vi�ƚ*;��l_�t>��{�B%�C�%��rf�TJQ=y����R�q̄"9��)�.oк�l:��ã0
e�L2��3�5MqmE�Y�ۤ���؎v�5�l��K�1�'�����ơ��5Ξ�q���tZH�F]�[�?ʳi�E~Wf�-�We���ӷ�aiՔ�NI:�p�.b�¸��k\��q_Fk�𒺵ZGm��(��)o!\�mf� �9�i�98\f�\	Y��%�s��\��.�幊J]}���ϐ�5W$"[6�͐�Z�67���x�*o.7�s�\��P���Dt`�y�6���2�؛f�)��yT?={��K��\�h�-��rgn[�`��c]�����uT8�0���u��u���.A�[6�h%�_wZ�tLD��s�5>R������H���wSL���G[!sO[�0�X� eź�C"����.�05��Ջ5��K�5���8���YL���!oC�HM�ʖ��˧�
�.���,.��G0c�z�K��fkJ��_�맧)�Oh-�v;�nQ��S���4�8�4m7~�)�Zb���~�Z�|����w�U��ep���1�=1r1���2��S����Q��&�@��|̦��.�R�Vr ��e8��|�w0E2�a���'�M��*]��`��>�����*]\�5eȿ�o�x�w%~P�3��
���[�բ��w"��?L���j�v1n�V}�wDve̌1(?^�J7=�<�o�����N��ۘ|��1����+i�[]�V�OH������x��MS+f���/���[gSw�Qυ�z:	�������_k�G���41�ֈ��]LkfR� �BR���e��2b݊���hMh*�^ʵ��R�^�dF;�X�<�C� �{�2����V��]�_er�u�z�6�du�0<����f��.BWd�f���6�\���7�9��"K�-��<�n�c�z��N�9��,ܬ��7�.�䲐���:k)�R������*�������n4�����oh|�ԅ��g&j�9�V��_n��q	��B��!��P�jЭ�[ީ����:W��`N�,�K��o]?�!w���X��Ge���E�=4��-\5m�YG��F{Kǽ�oUE�0��uͣ�>*��c(L��PP�ָeL�I����k���49�ha�3��@74p�T��uӫ�/�v��p�yN�� >T;1=�z�RN�5{�+3��M���1яD����1�F�o�����E_[FB.�k��	'V��u�\8N�V"q��>�X��u�b]�|V�^���SR3�jvw`ғ��ƹ�J�(MU���[�0�Ud��EF.I���Uj�#�7�;7���2��²�_PH���v�1���i��2�es˲��\S���ki":�\
�U�zI��s*��x:����Y��f�����Yn��`������ԫKu,��h"���#F��
&�'���jyǛ.��GS��l�%��s;�P�Τ"���VD�&����WP�;L�u�nw.{��&����Ō(H*W,��h]�i�$F�kYԵ�wL%r��=E5��{�v���&h�=o����61�w\�t�6\Z��F��w��WM+<)JsZ�@'l�;1,�la�p:�9������iT:��rQ�Ba���Cպ@�ڒ��j�v�vq�*v�9�:�]�.*k���.��=S{͜��fv�70Z�'-;=q�NMW���71]*6+5�g�ci���S������<���e�Z��T}W����
�J`厛�W��7�Ku���g5��*;G�c<����F�7s;M��԰ؤ�>X�w��L��r�%���uf��xs,�h����X������/R,N�r���\c۫�vʫt�p�kZ�»�>��x�X��͘9�jq�nelḉ΄Z%���|1J����j�5}0�V�WJ�rs���;�R��G��1�`Gf��m�tj��v�2��.�L��2�q����2+���6�@M5�.+���V��u+o�ݮ�ѻ�Q{�f���.Ū�M�|�%�+��嵐�r��Ө8���\^� ���L�mH�P�O�Ӗ��CXy��G����'
uk_�\S���y�W���.J��0}����3�3�q�@���Қ�[��8���بV�����4������*��NŬ~�5�QK�Q<t-�{Z���҆�I��H�k(����H��]D?��eA�Z��;Ϗ�[7�𠻅т�1N��3�Pa�M+��+��htȚ��jI,��"�U�XbTZhҋ�Q%�!Ȣ�"���i&T�ё3( ����5$*���hH��f\�+�*��Da�i��RH�T��2�QM%$L1iAE�,�9A��"�B��"�e�Ȣ��t�D
�8$r:a\�B�u�(*���!dj�N�5(��D�FlL2)N�uIE�d�UA� �.�G,Ί���Ԥ1e�IhETRkZ�FM04F�U�TD���Y˓L�	�"(�+�"��K2���IQTDT"���H.�E�V�(��9�kNEʪ.U�d��T��*9�
��NY�s��N!˕jDTr�4U(��(9f�P�2�l�M�$�,NEL�JYE$hR�"�8�mh�t��TT�����I��*�2K�\��S)$�P�%{���߃ן��U��X����y�iӦm�v�S�1�*��b�]mZ�U]��X�x�텙}�]VT;�i�C�U�h���Fq����/� �kں��M)M<SjU�/z�ќ-|i�؊AW�S�!�:��/,������n�wgh������7Dk��9e�;��K�{���=�[Ԉ��|^��a�ْ(���虇�s9�e�����X����Q,���%�t_�_�u/l�ܩ=����׽P��h�.�ٹe�^i���9��0�Mҥ�YIΓ�Nȭ�Dv�!-����00Y$�g�蜕:��������n��]ӎ����*#�8t���g�S�F�,�2�%���ͦ��!���t�e�%�_����:��ۼ��%� 5������VJ�=�埨���-N�-�O<ƥ�-��v�m]��~�UR)dE2�}�Be�G\@�d6"��kyYvTϷy�;�v�{�bߠ�쥴�o۲�Sj��V�Uַ�zE7d&x�eՔ"�����`��5ړU�~#GX����@��t&>ņ���R���ۓ6~:�Ok[��dW<q�28��P$����T�vl��n ~�8�W~uW���o��E��9u�< e��������z3?nZ�,�Q��yo�2�S�L&�xvҫ��tJ΄�1�t+�k<'6��7�޾��K�@�i�N�O�Âr}����-v�]q���0LbJ�Ń�c;]�Q����N�e�[@�۩]�U� ����8~:s���;����3��goj� ��r�}�mݏ�H���/�
�Yg�:��v�Z��
vv&_*�]M�&��w!m�w~�Π� � ��ñlR���e�a���8���Vl1S5�t���ۃ7��q�#��k9Bٶ#��{O^b�p������n�r�O^�^�[ ��b�Y��|kw��c&��}�~�1�	����^V.�um���U����Gp7ԩ�lEh�Ye���I�㹺E����9��|����>�n��������^�y�S��K��ԐmՍ8r,vm��N�i)�8E ��! ���H�NAީh�fT�^^���4� =�G^`���Ȯ��T��������\H?v(�jW��y�5#yM���E��]woJ����n+�~��0�t����[�SĨ��X�wJ%�@xhJu�����
�}���e".�	m"����b��´wòq�.��z�Ep�e"��@ܵ��71�{/� ��TX���H����6�]S�k�1�3���b�t�]@�l:/��u6�,�P�ŏ_�
�W����Ǌ�T���
X�'B��!)�t;8bc�l�������W�&��Ʌ"�ډp�e`�g��}�{�x1���[C��꽙w�4�mL���P�]}w�,@�.Y���R�Narw[�4��Sޚ���Ό��Y��zL�����U?J�5�%���a`:�a����Hb�H�Y�����,�W� S�H\Fa���5�
� q	�Z��o?![Y�e�g��U&���[��K����*���aO�#k2z,���5���@[=��A7�4���t-W��X���
�Z8�<��G�k�|��ʛ��w*�/�7zߛ6e���'W�j�4R�pN�h\��q���e�^���&Ѱ+��r	3������v���g�����/ǥ�Fa��]c�
�Ga8���hz��XU'��7b�1��w��<���tP���	�Z�n����G mr�&�VM��#ua.N�s�Yf+zwr���/���%K��D's^���S+�8�uOp�Ti�o�4�����[em��f�4u4#��F��1U�%�~��.�/��l},�غ�
��q��f��6;4W{*K�q:��� ��8�N� �[U-�h�;�iҾ��l6�I�̫苞O�ؚ9�������گ�Q��P�O�4�4?vײǼ9��y��4��v�4޹'���Wy�����s�QG(����z�Xm�"���f��;L5�����R5�xv?_[�e<��J\ʙە��k���┚���v��j&-��=Q9j�F�֓7�}@R]���r�]��\Xz�T�W���2��-�q�y�6:�5c�,w���M4wW`�=�6��.�E���2ˠU%܉?t`�Ɍ+�!�}QSQ�[u���͞N9D+ov�>���h�E�Q|�e��6����7D��Q���rmeNga'��5�����+�Hxh;:�D.	�8�-lk�=$��״�~`k2���-�u/�5=�ԯ/��B�괎�y��d/��ܘ�iI��G?Sg��(�:{a�hp��H6�����I��Z��I��f"��c�6���*B܉^�)�yL?;�a�71:]�T^�T�Gb��K�dy�9�>�]&_�PW&���š}r��Y��˧�����H�������W7�pw��Q{\��S,�wSK���u�sOM���yź��)�-��X���]��Mw�./�,ʣ�DcEnVS+b����ޗ~�M�Rє{.���+����pF����!]��0�ܳqm���>�~����^5+@�y��W�(�u�)��lW4���4mw՚>�g5�M�-2⯾���V���FFTG:���U1r1�I�-��y��m΢W8]S��j�_��kh�b�����ǖ���n��c9vMԵ��o.d��"��/,��)ҷ��e���sRh�r��Pk},�q1Q��XUw �����)1c�z��[�0WC݁�R�����[ήe⾩���Mir�;;"Y��j��jḥ7FwvN�e�2ޜfq�+����˶��?�̅W��_��Gi������Jw�*�uSKy��ڻ���t��;�R������d��Ó*� M0�V�F�q�G,NIm�L�Qr'�ۿ��U��݃�����b������矍�Q~}�4T����ʨ@������ ��;�]a���]T�����[gC�Y~Φ�1ң�T�y ل�f�32��^��9j���]LB1�ln�����)�*�ͽ�h��t6��2�a��9��.��^#Un���j�G[��`��ƻӘ<"�BA=�ڝ�s�%�z��ߊޤFoC��z���tԠ���O�9��̠ʙ��ܜ��[�b(���]E��w*OV�u���P��b�s"I�����늝�*���
��h�d !$;:S��N�����~��A�����D�9=U}o׺k��wI��-���8�M���,�: �8�HW��x�-���&5&�w��}#��F��}޳Ȍ�e��
�B[i#]"�����`~��9��6L�2�D������T��qB���nk���]N��	���;�`�J��O7��75F�;k4���\l�z�7�X�jR�u�ܦl=�{��[�����0V��j�P�w��X	�	q�:�(�}�J_;+�����%.�rn��^�=Te�E�y�;n��#{�:PyJw)�x�ӻ=��;�^i��H������n�S2�A�%S��'~f ����|K91m@-ʫ�P��{\�.�u��-�4���^��y��Z+Ue2�K��k��i�ݐ��cf�N�Cɭ��
��`�#��'�p�.֬�ı��g��X~<㶛o���p�ձ�M�n޹ɋ���[�]�="P��
���,�^�����^6N����E�8��r�/�mu�dɭ";�x�SO�/�Izl��{�@fSebGe�v�\�q���S�2��n����El��0R�l�[űJK�W%ϰ���j� �TB�k38�KۙS�\�2gIj9:u��Dh�*���[lG3����S�n7]7p6�F�vۖZz�^'�[�.�������yr���<B}���M���E{M:����*�_��~]��u*n։�������T�ۻ�l��b��6Dx�!<����B�)��m]\����ҟ*x������#���+��v؊A�=@"X� 	���v���/��ס�$xB8����H��������9Q:���=D���
�yo9ʇ����`���.Ͻ����r^�^sY7�oY>�Wj��0+܋��g���Tp���J��$e#؃�\ٸAX��C3���N>�;2mum�:�]7���CxyY�ٙ��r��]�Y����زy�ޓ�o��k�!׍Bk���� &�@�؃�a�v�D��B��{U�_vT�5X�^ꦊ��e�+�#qt����!�Y�q	��$�䎅�S+�����6�Rq�Fh9��-�S6"%��WRA�V���vN8��X�M�\"T@�暦�խ9A�)]��g�Ne����h&K�xԢ5��\+��Kmx�]"�tq�����۽�&������tuP�8tH�di�f�p���JN���+F��~>�5R��2��'�v �!��Ҍ��u�%���c�@�p,�p�i�4�9X�*;�ݔ�Z����j.]c]�qXz�m�z_��L�����x��o/��0�G q�k��}=9��j�/qVc�����et=�y�k)=��!oC��x�UĿ����@d��<)�d��ֲ�b̂&"�}�܋����fc��F��L�hz[Q�djZ2�n^���u��`��a�̤5I���4��ka�':dp�O�73�����^Ds<��4�l� �@[*�@�2�LM��a��y��~�'�����q�
KD��/����<�2�����k�0�5w�Ҭ]��.���WbǫL�N�G�������Es���K�<xO��c)X�Bc�EMY��&޾K�X(^u�F�޾��	���t�C�i�:�q�ݚ4͙��t�z�G-���0eD�\��Hǯ	R�bٲ!;�����8M�=�IV�5�����ީ�۽�XCV��MC�&��'�q�Fm)t���um���>)��̭������a�����/�b+CO������e�DO]�l��a��U{�-~]q����_�W'm�`�X����3:�ԟ�[EF��=@"|B �ߌ2���V���M:�S32e�c�����|�uM+ƻi�%=c{�?8����_�ހ�YtT�O�	<b}5��q�-�,b̜n�Ù�����n+�B#�l��=��M�H������6����7D�l%d2��;]Eelt�#�6�wN����|�#H�b2\�.��_�^�Ctc�7���k_(���m}z�>aUD> �b�3䇈�}�gP�������t�p���A��Zw#�qe�W
�Ő9���(h�
3;� ��	�}+.����ޖ~�b͔�F�7'c���Vt>�^�T�7r����s��t,���ɥ�
��P_\��4;}�?_����^q�s@�:����YCP7�A��/F��f�$�}}�;ٹէ��~�c��
XO"��B��YAV̌+;,��)���I���G^�kZ�t�d�9щd��U�����O�2Oq�b�G��޺�ۮ���7\<����j�;��|�5�f٧7/���޲2we�6����Q2,�wSK���u�!sO^�ɇc�,��C�9xX]@�Jzv�It^��N����&;E{r���:-�w������B����ǩ�����q��S��o�7<�f���.۔i�����+�7��h��H�3�6��e���h��:>����������1�zb�c���	����Q��G���P4��Q�ݺ$U����5�5e������W/Bzq8�.I��R���%C��Dԧ��dR����줩8���j����%�Lh�4!����eM=2EO3�@F��ǟ\�<�7(��;��h�vV��>��)F�7\�����b�^N���T ��xl�'�;�U��;Zg�82�tS*��1)�E�GO`��~/����:TsኝsL�3<���i\�uT��BIýN ��D'v����9����K�{R��m��h��t6��,h��A���� �旻�ힴ+�S�'�;�H�w�0xE6�H'�-���=�^+���=���DMs�c��\��nؼ^��x'b�YX��L��w�����)��~Ι�T�Y��m4I)�X��&�0	�P�ZiiݣQnO�0͈�1OnQ J�n��"�R��о6޹�O8�R�j���멲(�����T*��RzvT�&�{H.���>x��t���UϢ�ʦM�<S�;�8!�7���Yd#\�.�����/]|���js����d�?xT_q��t
��a��zZ����gJ^4�=;"����2z_�;2{j�N��e6�����f����w*Ol;�����@S.��z��h~K�](=�(�#N���k�8�����͹�R;j3F�e�o!-��˺I__���'>(�̸Q=-5��ʷ,,�U�~�S��Ϳ٢���k�(�~"Ʌ��vSu�*��"�wK��(��Êii���M<i���-W��tT@��(�p_X�u�0pcײ��<��ګ)�]3����OH��.z:�`P����P�X�x��U���d:�X��{�F�'/Ʒ?0���� ��M���u_�X�2T����9{P�:���R�B�q�x��mc��ws����(�Y�8���.p���g~���k�4?+v�E��?����^����=Z�.��W)���$�e���x�1�*8�(~�(;N����=�c���&7@7�y�嬣A��J�*�ñe).m�e�l1p6�8�>fẇ3�J���D1VM��.�	��D�7�##�yW]��M��Yږ�뙜*Qw�\�
A��yy	nY�=������N;���>�uܞՖ��dYS�ӈ�J��{ٴz�ui��%BH�IJb�y�e!�*���*����Ci��醩q����oQ�;�R�o}6R̴6�=b�	#a
���[
�q��MY&��A�F���U��i��Ό-ۨ4fb[p���o=���ګ�J��Ѯ��9�ͽ�¬,�H_�0�^ۏY�e�9^��S����W}��qv�J
u�fյ�8Q��:`�hoRv�.N��(��L��n��4���d�W&_QY��s�`k���[ëY.�J�%@�o[�%�l&�Oc�ʰk�Y9��j��bO�k32e:S8�Ta�f��Q���|��ʼ�ܧJ��Gz�c�Ѱ��� !;�F�e��5e^�޹����e١��-ۡdb��a8�eb�8j���@8������A���i�J��3/Hs.���48NwϷgm�#5h���i
n��I3LY�:��H,�kR�v�d��s���^Ր�����#޴����>�������%o�w��s�E8oq��F�C&�͘���ώBZ���\�o>�Iv� �%8�ٜ��+j��t�j�9]�9�ݬlTI.N+;&�3��}��X��|v�lu��Vhs�ٲwn43��ƨ�ZY�r�4wg]f��B�}#Չ����H��I34�V���i���Z�" S��u�P���j�\�Xjh�%�������Sw�����v!r�K�]S��YU륣���(�K�>��uS��+�!�jϱm]�A_X$�0=�{�>��n��"������-��1�[Y;50�u���u��^	]�hL�l	�	һ0D:6�@f	�Y��je�k]b\@��6ۗ�v�mU�͏x!'X��3c7�gw����f���$�u#΅���m�TT�s������峛�����1�$�m�W����Ռ�z����+�C�N�ok
}o���δ������
��ǖng,]�9R�M�0d6�re�v	e=r���+����%n�ⴋ�3D�.ڊ�K��fJ����=�1���:��]6��Dg(H�:�;.��巶k*����q�碧vrn>岭;<B�FK����r�<q��}Zƫ�s�N�;�<*���c:#v�{㐸�(7s�0�`�}ʟu�2��nd4��j��ky�	{QYe
{����)��8L�̼�"{Y�O
Y�(�׵��p�[��@,��B�Voi��cX�=̺Y��v�sx�wtl���|Иo�A���& �iD�Ζ��z��Ndk���T�u���o)9sk{�I����VqW8��yw�]�J�n�bTx��6��!*ࢥ��O/	��êv]���d'��l�m集ܔcҒAr!qOcgm]���K(2�����XX3��t��|��2��w�٦�`��]�8E��-�w�}�?��T]�S�͖�e�,�(���+��e�\F�b��sr���U�D��Uf�d�XUTj����w\謒�����"���r4�f�Eg.V"fHTi���kE"�1*]ۆ�9�a.��;�
a�"���<�*�R
����gJ+,�C)S%)imde�E%�*�eU�G�\3L�3�s;�J�t�º��5T̫kBU���t�U�I�]r(��)Q2�);��Z�3̤�z�n�z]Gt�Ƚ�����Ua���瓑�:��9A+S#�ԭ�4�H�M���%��W���K#��,9�aC�圂�d�W$�M�̐��h��N��Y���K���!+��be(��ܖfQ�ȸE�5dPU�Q���VP��S(�)ԯ�=��Gi�����5;V�I��``��Fؓa��9���i��vM]��q�Y����)G���Z��נ�Θح;�d}�[i�&P�mG3�-�b9�V��T.��M��um���~���1�������~�ڟ�G�� S�K<F�SLGm�
7غiն��qM}/�`���Sl3���,��9�WeD�j���m��T�8�������O7s)Q/8ں���h�s>���a+�Æ�r;^��]ʛ��WU������ <�N�oT�wK�R�8�2���kۇ#����7c�wd�]���[W��X�9r j\H?v�	�Ԉ�1�p��U������.�9ڳU��|D������~
��]:�5�H|�t�x�I�lҷ�N<M�=�ޢö�����}6␄Gbxl"ֈlLWRB�E����Wuc�{��E�685v�����R���xhJK�1�Dk�1�Vq�LQ��^]@��+������F�%E��ΠT�����߮'�yb8lK����УxK�]):'L,�!�{��Hd�o�D��΍���|�$w�Ƴ�_	kmB .��g�e��a�ЎV=�R��6ͻ)��.p��\o�ʙ,V1.��v��[5��vi�����}p�	�[:���	G{�\)���4�k5nQ�����%b��^��'\�� ��Ego���Q�$Ŕ��6ͬ�h�S��8���y��\��U����º�+���e��}���}�܃;y$e�E��ٙuj�s2��x���^==6�L8��g�e�����='�i6�/�n1�tY�F2�.nS�Z9���	7�ڷ�˲ỉ	u����~%�4��w�M6!=�+gQz�i��`1��p��5�l�g�f=-�Ų5-��_|n.�:;Ġ�:�O���Ͻb��ж�u�g0	 E3\Bg��[�<�Q�eʘ���,y�&�ꌊ�͒ ���n%��{���	t�ѯ���E��ܯ���:�q�T��h R��0�,vh���\�[M�~]X�V��/������%�,NKOO�%�h��ff��Q}���������������K�߄M4���>�ĝeW�W?��+��ICD�D��Bۋ:��X9�����;$��ns�;�[gK���.����\מ�,B ɜ\��� ��Ty�ឝ׋;�s.i�5T�G+%�BU�-�C��wZ*��|�)��P�Y�p��3yE{���wz��4�ۑ�5���٧�.Wh��E�Q|�]�k��A�gM`G��ًe_�T�--A�Fv���ֈ��_eJ���\�pL�5��M?aTś2._e^���l�扡��24r�]Y���+�� o+w��YWh�L��>W�ɛ5��T;7r��Uˢ>v��i��VB�gn�渶���82�	,rrΏ���!�	�s��C�`Cs�iO�Ͳ�S�x����Ml:���x������O�7K�Q�K�BYDK<�!���2����vq�}�iw~Z:��NO[����7U��hl�-l�KD�
��W~7�
����
9�S���v�l�=���ڔ����_/ra����T�1�?%����s� �L��T=-�T��:�f��%2������Q�l�m7h�]��}�jB·u'˫��rz�|�ɇp�6T�)���6n���#�w{$>
uc��B#	���+)��]TE��w��Rє{.�Gׄ���L×��o�Dodk�%��9�|�~����cR�ٰ�nI���b{C���Mڒ���kˣ��+v̊抯����Z*�����I~�CJj����'.��w���m�PPm�5͎�\Ob�7�/U]�9����%�7�a�Q�.τ2�����n'0�.�tV�ʇ��v�ۻq[�V�r�+��t�C9T�����FC�%�*#e��6�:�<�׵97_��x���m��F3�׽X�qA�r�!9.p�u�ARpnYΰ�2�{����C*�y�a|6�
�W�Wce	H��������v:s}!Z�uhRYvL+�����$��(p��5�b)�[�dN���Vwq9��H�y2�r
�s�����������w�_h�v5a*Mf
Q����m�E���*v��ܶ~�� A�ө�)��u<SҸ��-u"4������2�{GO`�6t?�����/�O>�T�+Y���o&Iɝ����Xu�8�����u4�%��u0�JSOڕv�m�~E�C���;����35�T�-%5g0�C��8�%��2!;��^�H'[1�Ot��n����������6���*�(��ȹ�C�T>�_u0��4��gw$�w�M��bq�z���J4�e� ��R��0�~a״�qt�}��ƷOKD�	��-όjBwӲ�o\<�W�1dS#�l�E�!-���n^��T��wI����K�q޺��q�C�.T�Z���0d�a&P~�Sr:G!���w
���I�����~�w|�QN��T8V����n�N�B�e�un�;�b�-�y��C$ah���M�ܪ�W�A�$.�wΌ��ܧF��h�-
ޞ�#��x�tmp�C���]�����;�oUk���7�W!���MkAܺD�O�ݎ�L����sF��q��k�跎�W�zV0*���a��ӵe��;���J�'>�/i#]p����M6�Vu){��q�z��:���v�'y��ws\��X��W}��J{Hh�D�֧�c�q���S��y�:��=7l�l1������b,Sh���#L�8�;9�n���n�N��l)G;2-Dok��F��z\�.1/{k��Z�14�((��:s����3��@�����ۻ���Z�����5�l�z�]��|���_��a��xC+�`̣(%�n�Z�%�aDh�1�l�'��Z�4���J��l;(��ܲ��a���ɭ��w�ʡ�=����b@c�D]���-�&d�m�L���G3�l<3�nu�w�e��Ga̲�?NɻuU��ܧy>����\gRKR��1]1t�h���Z���K�X)�L�)=f�v�Ed䇟 ��O-��
�[!C&_rbS\�������������D����ɳj�?6&�O��.��.Tݶ"�2i �#�D'vr@z`	ؼ�O(�q�*]d�2��V9��wl�8������=�,��\`�)Rʙ�� ]���W��=�����o}��I�9�� @:�����4W���{
��]:�_t����,��O�;�Vd��܁��$T_�F�^��{�Ѭ�m��mV(���ܭ�y����z*���l@G�Ι����K��7��qV�iU1�e�N�|�b;|�qn��Q���fI����ɝʢSI��W%�jA)]f*H2�ojQ���j�V��ׂN�;����=g\Sh�!bxl �"[i��H_�E��òq�3.��z�q�cYY�KE�T"��x��l�]%��"1�H������k�W�tq���=���KS�Q���F��B�ٷ�Q�%��I�7�V����~�{o�έʕ��)�Cw�uP�M�Ͻl�����X��7<�����#�or��Kl3��-u��[t�҇���V>����.�)�G;���ǧ��Ɓu��<�Z�l0�d�EN��W^��Y���݃�U�x�O�[���l�L����I�ڷ��&������6B*������.-��i���v��=��R�^��E	��`�0�W�(�:���7ǥ��F��)����N�#�Y7q}��9���{`���GX��ng x)�!3�Y�M��1+��n��h������3��MT��˭U7ͻٵ�V��zc���Ix[����~g��1����x��������{��lI�y��?F��:�0tg{��n�����&4SP�	p���hO^��"���	#�=4����&j&�75F��BhC����h�q+WmO���!{{�S�����"G���!���1����j1�P����Eɽ4n6��A���Β�<�NNQEe$�5��m��4��E���y6ls�]�n����a7C0��\^w��2-����H�9�lN�9u����p��|�)��Op=0_���b�v����p�S��������Q֪�E,��_������]t�o�uc�sGp�l�w[L����#\�=@"H@Znp�P̮N�u��ӗ���e��B#�L�!�T��j��lz�nt;���|�2�_eȕDL���J�u�*�GH���%�k�%���
��>����E�Q|���|G�4�����z�ۦ.�Fҕ��p|�B$�8"K �t����\k��=�!Eb2\�Ґh՜_�k1�WlOV҅JM�����`���+�xCϔ@BL�%L�!Þ1/~4���B9�<�:��o73u�/�=U}}{�_��q���E��K[:��!@�x�=L�-���R�ly��^�>鲑ț1�y��C���}<�����o�.��!�UH-�T� �֥���Y=�a���s�~�߶0���&���:.���5"����M.�w���\��odÉ8�C�*,����os+���p��njL���;A&�m��eeuQ�����,z����/��_O�,[�:�C�j����e���!����]��B�hQ�B��깕��ܒl4-�D��X�d{����{ WKz��u�+��}�e�����Ҥm��F�ۄ9�+�L�����\�ŉb9{�1��]N�wRȔ5b�v;��/S���`9�:m%��{��>�ɏ{���<������\EюpD��sO���ny�J�4^l.۔i������n��݊(\��v�5���E�h�n��Ep�"��#)�9�l�=1r1鄙��2��M���c��e���F�k~ɔ�8��@�.�}�3d1l���LB2�2�x�ň�9�CFo���2����3h��6��{T����Op�eR_t[.�/XrcEz� Me`��Xe���M;�vZ����sd(��T�ߖ�C�ְ���(�n����%��º/^dra�P�!�O8�ʺ2�΍�u ,s@���Ԉ�6Bg�7�ez:{�t?��M�c�G>&cu]ȻKk�;���^�� P� nz ��?eM1	G=���B�x�J�E��?�CF6�:��M��H�؋F�E�������b�ߋ��N`���	���xt���-��p�3��xf�Ȫ�t�ط�����a��-���@�tP�{QR��Yݣ�фZr��2�T�͛��^�R{{I�t�W�L0tt4b�!��a�2�����!�,~��`�F�Z0{�H�ʜ#�yh�pi�/Y�ȿyV��@f_�:���r#^�m��~�,� �^�t�C�{8ܹ���:�����ᵎ#�f���O�񔿼�;]�pѧ��^Tι�u�{;�V�����6���+y9�r���)�)1��q�Kj�b7�LW*O~a�$n�]ӎ��]M�: �5^:j�ѭy��:��9����������G�!U-��Q�O�[�˅7r�L���L˺K��g�����U~�wH|J��z���d��5�	�	���[�v�<�]I�-����vSu�3<)dGws�ѷa������[X�.��w��闖#� I�ᱴu��_��0��^�7��,ז�1�ՠ���-U�o}D71)�H�	�1t܄�:�X�m��d[#l�`ǯS�l�~���ߎی��F�P�׵X��t�[���{b^3��X����b��=m��W~���qu�C����|�}o�G	��m����Ѯ{�)��B1t�
۔���^��a� 3�\�0k����x=�lPp�4H|�l����&7�6�%;��F�ј)@�U-�`��}�(�y�Rl~�t�:vh��5�#��T�Ȉ�d�.gUeG�b`��6�(e��Hk]����b��v����J�R~�����`�����n��g���qC�E����V�.�$���C���3b�Q�����v�:U \�٢�&� ��&v�i�ȶ��Z�������Tԋ��	�%}&�����+����Pd�uf�gp�{�����p�U��q�C;f_[��;0�����c�t#�΅wKDWa��s
��+��\�o(�WDT�}Ѵ?^�B@ߛ�Sv؊�>b6�(�;�8�ך`��f�a22/[lN�Q]��6�û
��<���'׶�n��y��m.TݶW�:5��_$��H=��NX��7�r�γN�ʎ̩h����xz����d�7��m�5��eL���Ƨ��O�]. =��d�Q��9��������Ki��4W���wUF.�}��=�t�xQ���9S9G��Nc�;��>���\Sh�Gbxl �"%�������<;'l�ށ/R�߳��}	X�-c�w��A F	����!}%�Ԣ5��\q�E��aݧ�ĩ���݅����`b�o�n��Q>$>>:���J�5忋�y��u�� ��+��r��ɝ��Q�e�2fCwr�+�9�zЖ��� b��>�$C�7f�/����T9��s��kk�	�3ϵ�U���.���Y��b�G;���ǧ��q>����-~s�����Z���V�c�t��L�
ꃣ�\���Y\��L����I�ڷ��&��[���M\�9��E�;4��kz��._u3���宲ķ�)K,�����f_�����9���"�13R�U�'4tc�{͑�����l��|�!�\E�����]�غJ��ȇR��SxM1�֧��Kn��N�c��{'V,�kn��Y/�+�=�p����GE,��Gպ,j�]rvv�� ��<B$;}��N�I��햪��B_]��٤�8�5|w��YU� �S�����ԾC)�V�����/8`6;'8ܓ���%��U�}���4�r�@U���p<"��]V7o��꽆lG�F;��wnMp�o{~��"�;+M+[)J��u��cɎ��OX.�Y�%|Z�n�2ge�Ώo.�Nޙķ9�:���K��˦n�qYhm��ː�����������;�Z�[����%[d�_gN��2����v�b��[���J�������^�63B�{Y�]��ej����K[�%��@��5�chU��B��r1�]�}�ıä�M���������L�vՙ }A-twx��A�V꼁u�ځ�ćB9�@H�oI̲:���Ű+'��ز�F�������t��Η3ft�4�X��p�sl�f䉜�f�>Z;n��`"��<�x�������nd�pX�H��+Xzȴiͱ�f�)eG���!���W�6@���%��5ٖ����;��;+G�N�h;C��ph]�;�T��Qy�&hNT*�qZIj4�b\��6���I��2�l�3v�,f�l31hw�󻈧�rǖ���j�#��-���h��l�U�K��f�>���;c��B�g5gW_<��ړN^����cdN�c��=�:�w�`i�/�#�J�g8R������R������&Dr����U)R�M�fC8��Bp�-��lf� ����w�^�٧���}���m�V�Gv&���Y��ˆ1��X���6���9�K����&u̬h_hvZ�rwjoh;[��H(G�oT��-���0	ഭ���Q��c��]�M�\���k��t��r�)7j���om�.�\-�Z��A�-�*[O����/,�v��<x�7�
��u�I��I�+���+!� ��_v��v�&�$���A�jm۫!t�:[�ҏ��]��@<�̮���+#��Oz�����Y�R5땰T.�&ԕ}�G5'��u^��0v{�-Lҥ���N�>�C��6�=��YD��ϓ���_ʒY��˽���ޱ�={u}t6��"}4-t��~�ۏY�1^nk�Fr��)��6ul��
��^el�>Vk|��x����$A���0'��u��x��p��-�obYw�C��� ����ފ��T5*r�<L�=(��ju�:��a��Nن�a�}0ܮZ���E^�L	r��9��s�q��jPѬ�]�j��it��ح��`c7v=� ���57urh�މN��D�D&�r��xK�n�q'q#�N�Q��Dq͇�z�5:ZQQ�#�e#%��r�	dEGY��eQ
�]�]�EQ�J�Opŕ��5��IDRdgu��uj�ܗq�*��/:�[Ė*H�̢��֙��Y�;��xN���g3�t)
.z�np��s��ֵBC�2��p��']Ђ�����,H����rK�9�"2s�<�wt�P�E�R����D�bI滎�Q�G2�9p��.��eT蘦���af$���y�!U�	�'3���T�bIN��8�{uu��L=K�K��ԏP�")ّ��:'��R�=FI���Ը�r�Wk�:N�g�yDU�e����W��t�R���Ͽ�{��>�����(�Sڋ��7��)�99�LgZV�*��X�|�]��,�؎uf%ST�6��4mJ�z�H��Rwv%����8Ǿ���s�S0�X����*f{@��ڌ#0�py����x��SǆΓ5���k��w�*�ߎ�Ί�"��	�Z�n�S�p-oq������vb{�b�n߉{�ۨ�����,�#�'�x[	h��_��(�1���^�<@�z]�����~�ۘ��Χײ�N/�{�ڣM�l���aɍC�&�B{��=4�q��7b4�8��D��ھ�X�l#Y��7b\��p���=����T���,v�����N�ȾA�_uWU�����9?4�ʪZ:�Ѻv6�uc�6sGp�Ηu��?`1���06`[�棺7 �'� +�1g{P�l�!p7�uM+ʖ�MBU�/ǡ�F߳��h��!��<��r�'_7z
���Ygf�=s� �t;��Lw�Jy�6�H+[4�D.2�}�H��踎�O�
{;�fܚ��5�j��k*��tO�Q�,�1�=	N��m�'�B4�lFK���P����C����Mfc:�73j�f�S.�a�� &a��}�� �z4������y�J^;�?��!HgC&rZ�wq���:��Q�wʏ(/ơ��Pź�J��U��Se;��Uc���� ����R6+`�>5��0���a�ň|���'��H(��nݭ�l�w��Kl�O����]ھU�7Q�1��a��������Rqb66t���׸jo���C�{��:{Ƈ�H_���"$r�BC��h`Z&�jR%P{F�k@-ۙ�#dfdO{zS�o*���32�ǔ��9����;�����FhTp�"���z<a��i��x������Pxl�m2�M����ԅ��J��}l��9+h�l���a����f�^kU�g=9�,,��tW�E��ON`�ʅ���ah���dWL�+z]�E��,bZ��lf�-�]��W4W5�]=x���М�	�3�c�i���5+@�{��nI�궑�4��';oj��m�Ѥn5M^�4Sp�"�~��K>F:�L\�z�?�����S�f��|��u�v���:۞ۦW_8�CJ�ݿq�!��w1���@fP�W/Bz��b�5�������G	�wӏﾲ����K��_T��R_t_�d��91�_�'n�s�A��y��8S��]����:�|=.�_�L����0R�ι��m�E���]�|��*�T�֛�����jD&ԅ#�r��j�7T�=����e�Sw71l�W�&z#�u�#��o��
��r��:�=��c�[X]��<�Ņ:�:�ն�#�a��-|�A��Ѧ�7|�=���l�l�i�eT����no�kz��X���U����tPgK��*(:��&x�}S��oJ��ˠ��yBXy��u9�y��yN-�Eٽ�o���Ղ��RZ�$}��1���]L5B[�x�J�E��1�����j��܎y��\�����i�*��#�'�)�G���p�NYmN�[�R<�4Ђ�c,�W}/<�9E����h�c9���e7L�ʙ��ܗ��-��GXbL��k�����_�dj�׷�F��b�.^�;�'�{I�tf Z���
��h�!	b�*��,%5���2�3���ۄ�@)EH�P��O��#p���r��;�����
e�8�����'8c�ֱ�u� �e�)���8��6�A��j6M2ἄ6k$k�S.�.:��y����v�gjO �ᘪ�aj�w湞��8w!`Ÿ[��Rxl�B���Ywr��5�Xvz�z4���E�P���n#����c�a���H���x�uF����[�óL�תM�[>��[��u���5�S��y���y��SvBg��Ք5�B�����uB�{�ǃѯ�p3����^\�����A5����ܪ��*x�Zޗ=����v�==2���X���&u�2&S<��̇�5����6A��*��8 �����NR��.Lt�3/�����Q��M`bF�{]|�s)��3]����{uթ���Uo\����R��Sq򅪱'v�Ż�%J����\ղxs�*�N]'Z)�7-���y��fZ��ǝ56wxG���a=8�-��wyf��\�#��ˤ�\�_0o��Izl��{8&4���)RYs���.�p�-��s8(Lw m�Jwy��0
P�^�"��<o�������ft�ws����y��:Ĉ�cFmBg�/b9�c�pT.�Z�8���rTls^���l�e�i鳖#�MD�R\?0��F��U6y��+M:M��pۏp������/��^ˠpw᫩Sv��F؂+Ԡ8�a	����� �+�|sj�q��R&�#7v4��9��us��7B{^ΗCk˕7m�EpeOP�1 3�	ݛ���m�v��&z�O<+�����=0��ҕ�Ä�m��d�=�/�o����T��=@C5�J`Li�O���T�?��V��ah��6^¹�7N��}��OF��;Ck���1�kDrx�\Bؑ�'��p�nt���ٍH�+؈�ҺRt^��ja��,4���4^�{�\w��c�tR>Q "C�x�.��^5(�}.��%��_����Cp��r�'ߋ�W�V-jcˣt�@Mg���HP���E�OI��Eq��|'+�X%`("H�s�n�a��a��A����6�J�nh�K�o�֔��U'|0�u����]Ж�a�|G��8�b͹�Ց�Ӓ�Gp�mԝ��O}r9�cP,t_����������e*��k��yo�����&���{
7�`�}�w]�/r!���T��]BGp�|���ɶ:�,Bg�p�k�a���)�D<eK^V7n�D^-�x�2���o۲�i�Uc����^�gK��Ý�4����\C��� nڻ���1܍��źwo�'�5�Q�0�v�$�>:ܬ�{b�x�e�/�M����B�}�7�.�dˋ��a�7�qC�f0@�g�E�n�i��+�a`/.�F��Dv���� �,6��T=���;j�sEs^e�T*h�/|���tW�����L�x�t��:|�율I�j��u�͹z뱠s� �)m�3z��zc�p��/uA-��	�~c�({w��J0&ۑ݃����E�.�Ü_���m��M�k�jÓ*� M0��>q�N�}����k�E"2(��Z��l�>����N��t�Zn���;���/�b+EoE��� F�k��gl�����i�Ցzr���a6�1EmT�f4n����{�h�m�.�i�u'���!�߭�؏	��9+�m�d*��u�(eY[BV�t�-"��m�cP�Wqu��m�����s_#\���x4�u<#�@�u`R�W���bx\�|��]D��[U����ջ�Zq��Ee�o�5J�qW�*n魛���Z|��M�O]�z��8k;��oRS�\�P�@����uH��52��|�m4�%]��~Q�:]ց�l���ڬ�1;Sȴ���)��@��-;�:S�)�BA-�| ��M�I!s��rvN\O���1b��m_u��"YD8B|X9}!��qZ!pO��n_!���ּe��u}/}��3�l�0���wS���>Q	3�>�x�xĸ1{3���.�#���d�e�s͜jh�\�߸��:- ����J��"`�w�P�;�{�Qc%Y$�!�Qr9��9lN��弪����T�S�u��9�:�S[���p&�{�{��&��h�(���H�!�
r��[9������6�h���\���5!gC��˫��p�I�%�ߜ�eXΤ)a����̘q>1�qn�S0ȷ4�Ә2B������+)���Ddo{mLiȖ��MN����E��E������:�/BpF��Ni�F@M��+�R�-W��j,�2������ۄ�Ř��k�ɉZ����\fZ0�}Y����G�����c��;������Xy�k�r�֪�s�0�ΰ��;��(5���
�G�_:���+������_�wWM+��5�x/���OC�D��h���Vn��L�����[���"��j#7���չs�m��cy���@[+��]c������zG�E�z�H�w(�@;����/�79�]|�=�:���O�|kjf˹��x�\��(Mw�`#+y��u%�z$�a;.�o�'�嬪<!�.�ql�S�6�I}�k�Kװ�ƃI�s�A;�Z��MDd^��o3��!�ĈR�M&d��Rh�v5a*V`�������>�'a��3�ofE���,7�:_�dÚj� h�X�,��GM�	��Ī�[h����+��:��Z�1���6mGml���N���1� وD���:����~멆�KsF,ʝ2��{�鳠���dو�Hsb���/:�k�L�Ġ��)�Ń����`��p�N�IU�l�Qo�(�ݕV:�v��y�Guǲ�����j���St�����ܙa�rڳj�p�=Q��9Ɣ�(�Tfp�sKz����T���y��*���
n���d !�w��u^ض������G��ί�8�Gl�m���ګ�}r�Jt�;�����
]ӎ��q/���d��u4^Z�3��\�!��#�zE�Fͱ4˅6��^H�H�.�.:����pSfZA�{����޶��Vu]��ŕ0P�b�]���K�CWQ�;��/*��WgN��n�ߌb�6{:�G�6W�q#�;0t��&�T���2;O_�\���Z�}b��=����GW�EnY;k%\7t�@�+�ܔ�d��?p���u\�"�r�:�R��8�p�q�����ѫ�[���XΦ/U���jw����T�f͍@H��}�u2gW�����k���,�]��e=����kU@m�Q�۫.�,u�e6�x�U����;g��Ք)�u��^��f{�F��q�OvxDNQR֤m��qx���v4�ݒ�^ܪ�粧��އނ�鼆�B�ٯ%��c�7X�����[g�H,M���<b��:(I�q�g����{S=Z�.��Sr�}�~�]J<��e=ڇ�j�5�Y �C�1�f8n�~�(��& o�w���0
P*�ð��f��`���b��շ_#7�}��r��\���CDl���6Bg�lG3�l<�羭a�2�mV��Ӫ���n� zL�g+���@ם ƈ/�����0��J^H���c����6c���\�y�l�}/�`�]��u:iS�=�mG*���H?rg����=�Wj.(�:���m��"�t��j��׽��O��.��.Tݶ"�2��O��%�f�,|{T��|N�쁂�n���j�Q�z��MK��|Y�h����/F��D������V1���{�u>��x�K4+�mbw� v!M��i�����&����$2h��a8v���o.i�\��[ۓ-( �֝�Տ�yV�*,`�x��aơY!��b��IܲѸr��� ��-��0С*Ǉ^hK���!���3��K�
2>��M$�yժ�b&�`p#����H�,���A�<6qq��f��e�����u��7_;���7nI��h���8>|̳��}Ȓ�H_B1�ΕCT>�ᰃ�DKmԐ{~:�v.��u�nc����rq�7wV;�tW�Q "(L$)��p�ͱ�Dk�x�\+m)Y吕S�|��U���MU�k�^��@�a}�_X.l���lMlJ���3�
7��S^�Oi�
�{�}�f�pOi���t��q��ǏH��n��}�d%���:�,Be���V��~pI"�U�G���X��['D߷g�kڪ���%�R�����2��x�c׏OM��
����qH��:�s'��g�e�3�9���v�$�>>\���S<E��~o���D뻦����5�N�un�V+{DWc�6]�=�>K$����!Л��PS�c:
m�5΢#��uW���i��n�]����Q͊��+ݹz�n.׶�A;G���ΪS�\�";�:
�7�>��ב���D��5�,"�:�aT���:�rp�K��B��<�$���E�:�3oN�X����ήQV���:�-I�u��	d.��D�5&d�&�A[�:��e�RI�`a��d�+��k�^���G#1^�*G��K9Ͳ�v�������1)�#�˽+��zg%�*��8rR^�Z:S]#�u�0x��&�A�go�v;b��`��B��T�Re�M�׷�7�p�OQ����i�W�#�d�4��N�`O�HR��,~�r�O8z���O��{��uI~�����4�v��m<\F�e΄8�Π���%�צ��"�j���7N�ِ�{�h�m�.�WJ~���aF��Y5����h���z�B} ,�(��T3�6��P�К�}��ǡ�F֪� =K	���+�6"��'}�޳�+�S�� ɇw�ӽ:S�+D$�-�}"�Wh�x��'��ʲօ���-ѝ��6����B3�!���9!�Q�/�!pO��&=l��dUϺ�o��{7g���H3�d�8tfL���St�t @�d����L���R�ݛU�W����J%��Α��9���C�1F��߇q���E�t53�-�D'��5qsH�R�c.�km���N�5���qwj{ʽ~ևW��}����?{���x<��������������1��1�����1��������0lc�.�1��������M������m�o�m�o�m�oF�`���m�o��`��6�6ޱ��1��Cm�cm�M�����m�o�m�m�ɶ�1��f�l�{6�6��1AY&SY�?�{�'ـ`P��3'� bH���)�) �Q$�D R�T���E !	*
�*!($���*
IR�H��**R����**U��B�$��I6e*@IJ�I�eJQl�N��TB��U"����@(R�Q"U@�BPl`�5IQD
(D�DIJ���EI�5RH��5U�J�!*H
�RJUJR�*U*H�T� �*T��T�J��()J*�T�J�!"�UI �   دyv�m��8ss��6�ڒ�i���[��ts�����v�4�UE�5���a��V�N��U�3�C;���V���I ����  7<���g;٪�uq��]�P:��G�E�z�P 4h�G0�(�GGEn�c�:@ ��U�    3�� E�ѣ�� n�T�B��(h�UJ<  �QяAz��iE�9T�+�p�]ڭ��N�B�`�&ؠ�ùCkPݷu��kaAr�v��pn���l���U@RT���<  ��̐i:1A]S\��T�.�76�PvR�Ҙujû�k0]�k�5ݺ�7W]��7vݔ���Z��&��WM��k��
��*
$�Z�T��^  �kV�[��:�9��m�F΅��
��kwmۣ���]�6t7.�;s�vݳ�ݩ�R����Xʻc����ۻn�f�-[���H�n���Ӷ.�E����)#��   ��yv����Wwa�ĭ��Ի��5F۵�U�]�vջt�M�0�P�9�u�)n��U�vv�ݻs[m���YuB۳���U�9C�]p�wN�����R �HP�)*��
�x   cw�mD��kbMMnMZ
�v�vM�QwUlj]��֫�n�Z�6�uC��v�B�.wmݝ]�]T3��ֵ�;e�ݻ�]�n��nG]�ۣ�����D$���)E)
	�   �jZ]c�.�]n�h�[�j�k���k�����g[n[����\�kW]2v�[s+X;5u9��M�]���uۻ]��F븭���mݺ���ZP* шR�   M:�����Ӹ.T�GSk��v͘j��]�۵t����7i]��]�sC7lT5�[c��w3;wi�Y����[��Y��Nݍ�kmm�5L�ն�UvC��v�QUT��E]�  �u�vծ����0�ָ��홙u��"�Zƨ�]�W8�I�]C��ۭ76tm��t붡Y��:����5���:UT���J�m��1�� j��I�T�Pd21�{FR���� )邁�  ���R�  ��~D�UJQ�  I���b�"I[ p�J0p�"P�$�Y�5d3���L�Ai>��׿L��ky��}���䄐�$�Є��$�H@$$?�	!I�HIO�!$ I��HHs�9���uR��_��JV�T�RJT�ݧ��\Z2Ef�f!������Ձ�i����6���| ,U��yB��i�A�P-Z��t\W(��úL�٨��ZR��B�1��t�Kem}�V킱�Y�H�3A�*����
���wZIt�Ôor$*i;8�fۖv���o+$���sR$\1�wi2�)�ɀ��&��⦵�gl��Ƃ�� �ͱxF]��6*���DTQ�b�t��������R
�Ħ��q����)m� м/u^�,U��wt�;�b[�ưp�� V���2���ٴ�g�hR1����b�m�'sX���i;�F�`��[��rͩxJ����@] oZ�Wi�x�*WJ�t&�I�ٗq�y�3��7��U��b�1Ԣ�N䣒\
P�����I��h�r�o
�z�#i�!Vl�tf��G$Ab?-��o�5�v�+3D�J�h���PKr�j�Wt8n�F&�cq�B�*Zn��`Ւ�he[HUڕ�f��Ĵ[��9w�Ř���ͦ/Poc��Z�{���*�Ȗ��q��Z���n�u�>͘!"RV��)*aM�g�Q��Ƚ��.���
<��wwk:0��M��R\���M�hٮZ�%�d��*�l��iM�jS�5>7D5j��r]��;N]�αjE��aC�`r��m��)��:�`B��1�V�]��/M�X�3&�En� ��{R��qj���&P��[[��4C� 2��W"�~2Bn���GpAi2�:��+a�����2],�h)��nK�6P���X����k�/3%�`�h�G�CAݷ� �`+t�ՂLː���ػ�edk_-��V E7z�P	mc)J��P"ٵ�kV��`^���Y`P\�4@)�,Mœ�e��tV=��A�ҝ]\��vr:Ke�:�aٚv���7U��R[{��j�I8QM��+^�8�Ncj��Y%"�J
�ë�D^W ͇a@uu�y�Ғ,�-C�!���A-���=�v�j5��]�	��	;�4��m����\�?�4QW����LX�s'R�F%�\)��Sؑ��jkJ��;�uj�KBKk�2P�� 4�ɔ�˺n���l�0V&()RD��"-�;o�aebNөd��C)�� ��ϝ��]��Q��n��B����6���]dUz�D�Z���C0���	���KQ�H����F��oRY���%Q��(Ī,�`Mq�����Uyb���V�Q		��8,� -A���PC;�̍;��U-��v23�L;���5��i�҉r1��*�k	�EP���v΂� V]#��L_V�z�!��)�t�����Op 4L�[V��ʲ�l��f�Hbc�
U��ơ�c٦L�r���wt�n�����"�gM<Ż
&����Z��������ݔV�>��G�h�IJȅ�2f�ٙ��Fcӳ5lQ��ݷ��[RJ*�+z�e�0G��/-��M�\�^�t�[� �C�2�� ��F��CDZ`����u ז)'%����ࣄ�gp����e�n�X���z*���7 4��
�r��Y�t�tn��l��ٸ").V�^����_L�bD�;��u�0�2��I%���A<cdn�\����d�t�6���a,D�H[; ˦L��*�e�v��R�͛r�v�D�g�s��!�Y���Go)ܴ5=�Z)��(��0�N�[�Y�`�j�/4e����u@�L�6��p��
&m�=�c�ƮS�Zνu�E��w�H2��sf*��z���u�SM�J[z�����76�EVEbz(�o��Ob�5\7�)<�X�y`���̽��4��Hzꁫ'���6���z�#�+	�U��f�XͲ�/�Q15�j7���zbIQ�a�T�Z��w um]�VM�7>���N����tʥ���P��e�/r�!tM�Uy�J���.�ێ]y�6�gt:�f�3d�@K���A�&L����fR�Y���v��H�sr��t�Mn��rbD�܎ ������{Z���+U�<a^��T3N\Z�U ��	$��l�kl��F�v.��:�0cT);�C!�
�+�w4�J8��m�FK�j
V�����Q�h�[�f�y.*Ub�8bײ�d�h�-6�n��;#A�����
�7�i�J�vj۷V�c� ��6ehW>B#AU��h:5'j�L�n��@eb��ۢܔe��P��U���9�.m: �[�/n�3>)�*�M+��i��8ɘ�EiX�Sj	2��3 7Yjm�����&���ͬ�Uu*���bD��VX��"��f3/MPR�� ����v��۠��"�f�,5[D?��]��'6ls!���Y��;L�o%a�ZC�l�6��n�� �7N�6*H�@k#WC�����X��{��ɘq5��ʖ�HM���*$q�Uw"�e��$J�j������uً�:Jv�:�"!zF�&��P*jL��.��5�?�k���hff�]�J-7���G@T�2�X\�%��
��A�Y2|�\���� nC,S�[DU�����b�H��sd�*\Рv����tƍЬ^��ةP�e+�?�w�j�޳5T��M5@��T���O�&	�a�X)�.�xl�F�{j�cJ�WX.�.���4*`������介���V��E��������y��Jx���ihl:��щ�ĵ=�+t�dɐn��T���z���.;��*� ��,���ޱ4>�-[U�`̺���t�������)6q&7I��=����FлCJ�S�R唂�K[�vS�E/)�NR�8L��4�|ц��Cn���0��f�ݱW�)���N��l�twYX�{>h|Ӎ��z�HӽbR�L�h��ʦ1Mb{wMv�ͫU��N]�p=623�^kc(�r�u�j��C,�r�"򤬺����Y2�����R�h� tw/ę��dX��P����[�c�D��l��ӹBՔ^".'WDS����G@��+]]�,dx�\��,阰L���'��0����"(:�iM4el��n��5R��k ���ͻ�eA
��5d��v�aR�RcW����B�46��fD�CcTj%Qn��i9x��LU��*�֠]`��A�dձ�w�����g�)md	MT2n�A�6�&hҶ��D����v��MՃ�&s��`�a��#�ν��u$@�Th�2�<�(�{��V�W[�"cZ���9�ɕ2ϘZ^@T��Ѡ��Y��c�x�Swt!����h�L����z�)��K : 5���k��`:�V0̼�RЁm��c5i�vc�q�V��qeH(3cak1j�$v1���LmSݧYZ�\*�c�2+�L���x�V����E&�0B-l���<��FN7+a��!��B�;�Kjl�:[�X���<T��t�S����
�w
򉫫
�6�5+���X�BMf=v惌�X5�3��A�Z�D"%0�T�ȱ�2���2���
������\�p�����bN[u6n�NG�ۅ�V6�nEV�f���s5��c&���῕I����=���m��� $m�##��ETtiޱ�iU�#�J�{m��Eyl���F�O�ORVa^��2��]�߷n�v���V%P��-�:�4� -�P��l��В�l��*(���t%��0�l���D70/h��v�d��abN��(kYO/lѻ��7H��A���e*��ޚ�R�n@vn��%��scw��,|v�,-�l�r��yw��۶qe]�J�r��۫�&�ڶś�Lubҩ�e�+9G�Vi7d��p2 ��uۻ�s,�Y�t��LI��J��r����^V�{���d[�j�!
` �D= 9YE�q��u�̱N�]��U�޹eف;�d�M��6ͪ�[�T���j�`�9�l^V��AZ�Î��K�-Ȅe��<�`�v�TA�J�C`k$���q#+]��Ae@>�9jӗm��-x,�0�!�Y�H�;�iMf��S^+Cs�t����y�F)U���1M+�YN}q���c��X�T��6��n�t5GZ�1�,���i�p�Y���g���Xl�S5lM��a&����`d�E�a���n�t��˕�*	y"4�F����bښ4�d
P<�6�Y�k��#%��\4�
���h�/O�ŗ������	R�lXY-@�Ã�������j�0�M5�Y�j�mѽ�R�(�$�Qg��a��0�&��D�V��)�6Ly&M�Um�FIM'Z�v��4ve����h{�Z��gf�xnP4�L�����O3F�-���^֫Y�Y�K�/6n��� ���Ǌ�B�5��f�b�
��th�TN�Q�n�nPB[�:52)�(�B�V���G��Gc��H�0[	2�eb�
�
m�[6��I�i���*	
�Ub�URUԱ�zkn�R$Hڃ#�Q�:͗+������0ra$��X��M��Fi�WLFQj�T7�bI�DQ	I��a,�/���	�ibeF�%ɖ2�YJY�i�F�;ٜ%av��l�$wK�f:W-�[xn�7�ڌ��0�;���"�bM^�XI��m� Z{�F9�:t���j@�o�i�7Y&�b"��nXl��â�RM�{GTfl{1J�V,6�K��2����&:��<�[�):��0(�#Sfm�"�'[R����♌�;�ŕ����=ki�u1m�7mf �Õ]�vaB�r����;���7Q��L�1v"lǚ�y�]��F��b	�u�aP8oCʗ��t�WJւ-*��q)�<��b�8Ѕ퉷00F��vn1��M	n�f7^]�ڲ {����6��3u?�ّ����\{�ɷ�^�f��� �,��F0^X�ՙ��n���$l�Le=)M�3V]����U��o5�d-�ݷ�4Hؘ��}��b�n�FZ����#SԵK �ks�5J��g�6�"Y;w����ܽ���H���%�Y��4�6��@��Q�(�Zu^7�l�����J��a�X���]#I���0E74I��k.�1����C%T�f�{��� ��)LL���q�E���f[��T&���ݥ�n���+[��TPd֩R�]A�*�y׻�B":�Z3i��b�����c�/Bxl�5"�6��S<��YJ�fK�4"ҪJN��ഥố��5	�iJ̖�e�X�YB��Ǡ�q��6�bu��cu,�͚���۫�	b+��2ţ���X�V^;�k��$T��� �>�/��ؘ7̵YwQ`7�ìa�L���p�+6����}t ��9i�Z�Rb�8�S���U�bUm=�����"���u)�֦��5�sT0�(���/p���ef�I��-�M}���P��w%�YR���6f �3�t���1=Q��6��h}��[j�d�5V��U�۵�{r+�.DvZR�]U�
A0f��S�m�H:/,��
 a<S�)�afc�E�m=�G"7�b(FX����S%֫{�f���kYc鶶�&3�J��kJF"U�����*�6�ʡ@f(�ٚ-�Q��n�j��cV����La.{��vRԳh� +���߃%���A�6����:�#�n0�S)�F�ހ2���"͋�2�F��4�.Һ� �mM�I,��YR�wf��YH��y��Z��f0��J΅��9`^��ܠNWu=����ĥ�y&<1�45��Q%{����h7kl��h=�/ 2�Y�(�Mjݗ��Sg3sk\k�^�jZ�
��A#�*�b�?���i�V��{�N���E����?1ݐƀ� e�F���	C)��P��l`-�[.8Jc��V闤���P��-)F�%��4ٽ3*2&�R���V��4�%��H$�o^ZEV�T��5KNJ˸N�Z����Iy�D���a�4d�R#s�-���b0���N�A֫�Rk3_n��YAӏkr$��Y)8q=�ɻocO3T�д��+��0�i��`WZ�?,�s��Y��L�S�eˬ�lb����(VH�C
�Ç(�Bl�&���Jw�%X�x.3IF�nXÔ�zp"����vnU����b1�Ksr[Cu,m��c]Z�IR�맚xnH�Z��Pn9���(��eZ�"��t���/` ��T�ңR�,@��0��[��ї3n]#ݖ6V7i��yP��ڲW��4�V<@	z1�l$5�f���e��7B�>lC7Ba���q^�I����9n��:fV��l�)R '�̉Ab�VV���SɗU{�+]�tv����1�=�Ƕ�=&'/��N��e��U{���⴦�e3F��p�z/j	�<���@6Vk�.���M����4p5�&n�x�F���b��EGr�X7�Z��N�V��?B��e�Dpbƅ5��%�V2e��)�Ӑ�eF��������.���5�d��[���Ҵ�8�k"��N�|��[���b�V�ڧ��NΔ��v�nS�H*� ���M�Ɋ�ѡ��-�t���--�ux���h��J˩�m���e,w�*X���A�dT�`3U�mn����M�N0h6pK�^+�-�5�"[v��ݡ�	f�7�j}r�:���+B��&cU�V�N�׵GN�ط�����	��u�B�oeBEEG�U.enI�f��1����.��p���F�q��H�Y@켹%6Q�VΗ��?�k�s�8]hS:�<����uɒ�]
bZ�v����OZ��T	S�zgr��c�X.l�=����:Ò�V4�b��` g���c�|kj���_CA�7���[F����r��!����n�:���]M�,�����T�㘳3kz�-�}�9vԵ�ZJ��!���Swmպ�37�D���pio(�d=�c7�E��m���.�T(mvGąyNݼ?eI�-�JGh�>���x� |S�U�l��ƺ�ɣ��G�=W	�Wk[.��yS������p��+vQGA(>4
`��E[ti����D�v�r��	Uok�����>���`4� ʁ�v�T��0)on��U�b��G���ut�Z�����Z6iݖW:�z����/�!d3�νѻ�X�����V)٤]hv1j ث�S)���iè5��_\I�V�u�v� sټf֊�Y' �2SGp����N^>��\��8����e.�3�D�W_�{�0�0�/gWJ�^�,���RPU�dc�����φ1b���r9�٣S��Z��i��K�8o坷�	K�/7l�UI[��㣆:�gn��K�]��u�4"t�����Szj8ŻKQ]þ�x�����g$��r)our��b���ἲc;U��Q6x��shs�[y���Y���.���4�3@�j��ܑ1�%˻�oY���b��\W����u<�N+�[�q!�捦:�i���.���U|j��.jT�˭��80�v��+�n����U��X#_����-���6�o�o��ȒY,}h��X�Nfȶܱ����*�%HC۲�&���-��8g ̳�$��C�W���m����U�-vm�tc���vsq=�Y�U��z8īV1c58�l�z�ѫ���Y{}��"�NM�p�]��c�b�uҮ�����"���4M��r��"���9Y@���$�����yJf��V�^��rU?��c��	���Ɲ��w�G9�G{�Wu�r�[��nT�+f�|�3c:7s���j���B�L�S�+��s�{F��u����Ӯ�;n��Q���['Y���A[�}}o���kc2�c�N��i�q�q�=ܝN����d�)�4{�-��u�e�]|2�ͧ�vR�H��QB�
j-�m�ٻ��1:��Ju+@�'.����x�z��o��Q���.N���K���W\Ŧ�ֱgO]�A|�9s.Y�I�I��ih��i�6է�&͆"\��l�4��v�z5���kr�o+�쀊�[�{�<���ĥ�{��˚Ͷ�T�DHлݾ �g2]�We9�/el�=v��u��0�fP�����3�b*���B���j�Wj��s�Y�^hj��6��a�
�'V��=�t�O�n��zv��b�%��s��O���E6D�x*j�=P��z�N<xu��s����I����斂��ukz�rS���2ғ^��mY	��MƨLǵ�l.����ì��yV��j���t���د�ݥ�>��݂��ͮ�U!�:e�J	�lvG�y���A���\� �zb�p�L�k��d}�d]��{r6��1v'gjK7�(��wl�����nI�j4��������hf`XpsfNK0��tlk�մ�h\�ج�6�٨ɵF���S]��oi��2����9��W<�¬�q�5�q��Á�t��3���ٰ7D�l��X�Q���V�ԀJ9���:���Q�{˝Ս�j,�cn�>#�R:x\�`u���C#��Wq����7A�y��X�c��]O[,<�
��ߡT��J�-��v�=t�cZ�U����dZq�5u��u�n���y0d�5]��r��ʎ�4R�;�n�]�k`�Ć��9�}�����OP�C�2���IaUf%�|S�tGC���F1��eTRq��1H�����q�{���|�� 4�]��7F�C�*m���v7N���klsw�ڻ��ў{}�&���龬[�k)��g����Zt�e��x�g���u� �b"��Mg�tU�f�TT�]�u�Cj�UƲ�n�K���2��f
��� ;���I+n1�r���8��AV�R⍠P9��;���P^�	-�C�s�U�f��s��(��g7]+�}Y` ,��aC�eY��w�ǋ��њˮ�-�;���h��K[�c��1�:z1"�,m��*R�GM�+���ֽo��Y[�F6h-i��Gn�7���M%8�iF>�_UЩ�����o���Q���Z��<�ǉu}4q[��f
rP�}��b�z�J��_]]��sJ�p�իU/IXx+9�&vn��C}D�X��֗��F�@�坙+��fLm������5G��e�.۩��z�u�}˻����[���9�M�X����˰���H�:+W�>��ym�����U�U�U��+���zsS���{]�h�J�wc�z9<m;�F�o�⮓8t4i<��۵k�!'.'nӔ�;{�����Y��x���̼�@�Ǵ�}���pZ�ĺ�+\5n���m�3��\��'!�p�D�dR��5���zK��s6Аh]nu�G!GÕurG�r�j�_]]����%�5�
޹[mU�up_اw �n���c7��]���k���C.L���ޮ���ޡ�M���&�+i;;��eˬ7��w8�<p���U��_en�:�$m��#�"Xkk�\YI��*�x�$N-9���7J�7{LWʊ��#�i��}ۗ5�ڜ��jl�8��Ev��}9+�+g_���0����K�ĕ��`Uo�G�����c��P�v��V�\q�T��1�xpk�;2���!�X�h⧎���k���֧����ޤ�;������NAh[w$����A`q�"e)��ae��-�!ƃ�@���U�u�V��u�@-rt���7W\�T�}�|��r�-����Ct���1��n����p�)_s�<�u/g
J��;�(Up{N�e��[�V'b���+p7�M
htj
��:k�1�H��1󫭤7;�z�L�"�%fj4�:w]��Í�j:LlH,�o0����=ޮx3��o� ��Ic9f����w�.rS���$V52=y]��w���w{ڻ��(GF�o:�ˬ;[X��^e�LmL1m�ح�Dݣ��i�YIs&�}�|NԲXhP5ӡ=B�1�h�����	�7i"N�asmh��j�.�Х��4��S;���Gx���r�2�u1���[ڗګ�x�����]hl�d����e�k���^8�[��A�6Z\7o�����?�L��(;A���R}R���m�/�2�����UgV�]=>��u�7�Z�AlpO��+և����Dr��]M��拹���c��`�C��r�)����g�7vv��hr��ݳ����ST�z��>�9.-f`�z���[��e	'���Q���IE��N���ӌ���`�)��|�)\UCj\w��Y��e��u� �V���Rm�5�_md�U�>q��ʖ�l-e�"��=��J��ꦦ�>�r&�n������E�Y�w��B���h��X��X!�E��h�&���*ǛDfu<�<��i�����|��ᄆo�Vn�HV���mp][0���X��G<�����!ҥ�k��N�{K�����y$�B�f���%4^��FR8�,���#vx�x��\�+����ݬ�����
�lĲ�q��͖��N�3�_�1a��O�3X��hP�u��ȭ���6Fj�Y���e��ɐT\�F2�0�	jϮՉxm�=Y=̺�y:MB�׊��E�[�is�997RY�öfH�/v�1	w�5ʌ��r���� ���M�;c���i�E�rsaB�&�Ы���ĸ��ҝ2�PY��ɒrAD'�+�L^d�v���jrV1�gUJ�tm����E��J+�2vή��/%�Ԯ�Sf��`���tsm���j1�"��O8�G7�{ۭ7ܺ�E��WG�eiv�o3r��i���G��K2n�z��7���U��ƞ-�7Nf�\�+��T�G��-�\�T�]}���xu�^��/[>4]d��_1t1�"ܾ$�YF�战��'eaUmSr��ں%�n�XF>�&	��Z
�:��!D:�o5����\S3t��b&�yic� F�F�S�Ο�_���)/c��iBF.'I[:Q�.�_P���dZ�7tEҾ�ҞY��O_}X���*�\�J��{��f���#]r��OK�liqt�˨�],���k������z����$�Xu�ҟִ��%�e��Uu�!/z���&-[b�M��gR��u�+�֚9�լ�F��;Y/rĖQ4͌����T�j�O��vW#!I��/(�m�4o1��v�r�)���Cp�ɨ'3�g[��C�\�y��٘��T�w�+��=*�(�N[�3@#��� c����D8�P/2e��C��>���P�v��j���Y�.MB��d�������Yɸ2�O��/{���t9J ���.��Z���N��3V��Ja�мGBE��g%wc��.���c�{T�yۻ�ֈrbW��t3-s� �ƪU�t�ҹbK�Vp����g%�f�Ӂ�f�.a$ܳ����2�gVۭ�I���0�r�{Y�(X����+��#�9��s��c�VvP���jU�V��ڜ�o��v_w  Oy�3��d�T~�*�v��E쪩z�k,��<�C��G�k�8!Ke<M�:Ӫ��@��Y��!�{l���{B݃�C���V�he-Ռ�.��f�02޽�+*�N*�m!�`J�iK�F��`�H���sucX>�5=��Nn��۹y�����F�.k��r��F����Q����4Z>j�}.�7>��
�s{�R,��z�}I���h�+��ow��]p�.Q���I�ιQ��҉L�v�zi�njfgs����"ޤ���յ��]�;�\�ك�v�Kh�s�I8,ڴx��u{�(�T�t:�i���v�����GVyzk�#��V��f��=��!��ѫ)����v�"��zs�6�eKSg�Īq�k��m�z]sg�Pdz�|˕4���u������ހ`�:��1�"�:��N�f��z2u���@�mdW7RQ]��̍�M�c���ΗtC�6]N+r�-���"ߒ�h�������q��f�8Z��e{ϼ��0n(OyY�YV�n��/��I�k�X(���N�*�=;vCt&޹CP����:Wsr벋��}��:�����kz��Ӝ��L17VgW_
W�Í�%e�)��wd�U��u�\�p-�-P[;:�*ˈ&�� ���D��xnn�z����'BAܑ\�gu�6��|�ɜ.�<�wVwL��}�cu��[�qg"�6�2��e ��9�����>�C5�k8X,�7~�B>�Uoa��wy�L���@�$��u)��>xu7S�����9�<w�ш���6_t�[���F=�[�d[��G�Eٽ�v%�$ε�9��EgƙIL͹]��h�sz�	ATR��X��tt���]���j��Չ�1%����U!��v��l��P��2��W���9Q!+�l_)V�t[�Ԑ�&bO4&�v���z�[�K;_:�w��w'BZ����C}�rL�(�hޢ�V�����shK�x�j�/ �L��)C]M-��osݗ�b\h�`�ߚ�����K��LyB��d:#d�T����r�gQ-��Z�oK����V%6rY�[��(G�:�fW2j�NY��[#�ǵ��@/��}X2�3f}WW,��*^�Kq=9]�ݷ��uI�hd�֮9�<���ɫ+pn�L�GD؟N�K���iiJ�ڀ���b����pʾ*��Nv[�/må��P�Wu��cA�F"��� +6棙3����M��I��栀�M��n_+��=��^sx��x�G�oo�r�� iP3yq*�֕ul�*XF�<窎c �{�j4����['��z5������Y���eP��=ɸ$��@r���r��e����<\ʉ���j�����܆,�z@\u��������#����=Ćv�
gz�B:�|��t�e�lv9ݍ ����n��<-����dG�����W}Fcu��-N���:t�{�W;�$����K�Zo��]|Oo] vl��*���s��T���S"3�)ef��F6k�fht%�#�o.�G�$v��K[����$Pe��UiU�|�*�_d}�lHN���Ҳc6`��湀�̛��gK)��V�Փ�s`���m{�vW}!��DU��m�֨�C���]̋��*vtr���d���q)̮:��7]�+���*��%Z�K87�m�L2.0V�O�����m�ʱa֖��q�6��w!��#43 ���+nPJ�DH�۠M�h.�줙�5���pT��t�E8X^�Ǧi`���rtg&HOV��h�ٌj<(��)��}�"b�G>�0m_|{RuZ�O������8��ӺQ�#�)4a�Cx>�H�뻹�vvn��pd�"��%�;6�(�89��]�����f[
�p]¶u�>�-h��:	���9�+NN�u�ϩ4�S��\ͺV͔�I�
���W�8r&�����s�ˈ�%�z/J�f�����v.�h^WB\b8��}�ތF�`Pu����m���ս*vfXW_wf7�D��k�4.�[��.�l�=;����E>=ǸQ
�}�gs��m�6��m��5��m��t�o���|�6�sm�M�lcm�mߞ���������H@$$?�B��s�Ǆx�ގ��JN�F�����^��v��l�[M[�\+[NP�e�Cz���IL��+���U���E��	�΃i�b�N�t������R��s],�]����.������!�		��3���l�%���p1�ņ�T^5i^��T|k��� N�:WT�Klo]r�Z9��ф�Z��ˮJ��u�����V��S;zX�r\(<w��ՠ����u�xv�;��=��`�%��u��x�q-̱���)�6��<��ܻY�t�6w{>18+X-�_^vIH�H.=�D�%.n�����N���|�\06���멧�#��7y�5R��q����3f��BkM�yR��['���o�#�ݩy��m5t�;�[T�@�]�O4�jc�,��ɢ�_�te�W���vG��r�<,�73�Ve��/�9��C=�[T:�������c/5g"H
�=Or�Lׇ�\J��KjR�Af�:��"�m�YJ�-��Cp����[�������vI�an���j�3i.�����������1fȊ�3bںv�h��N�V��|�wwb��6�ky8U�KtѺ�M1`��۹Q��,�᫮�6�_+��p��70;����{м7N��sӕ8�§��-�-�\E1VX���P���[��c.��9 ��k=-�i�h��q��E��c���\�N��֊L���Z��ƅu�4���/4�����M�3�����G��v�Rc�̵����	}S!�ʸѝ��Ϗ*5���ܶV5��#x�e�u�*}��u����=�N �Ɩ�n�2���[��;C�weZ2��&�N�����*�商Ҥ����{:�$3��1b�?��b��\.���sg�	mq���g$ae��f��56�ݭ��@��,�v	:=x��Ŷ�-��-xq/7��@W��K˼��.N�X�¤c�@&m>g���u�����et�VZ'��4tۣ���2�\��bL�uY�s8]o�]X�h��ּ������d9���H�'_do���G�.��D�:�˳%`K7�r��}��l<j��$Z�r]��d�onNc6\��μѝC��m'��2���+;-nv6`�OpC)Z�ʴv������8+J��]��W���V%�f;-+Y76���S���
S�{NЂ9F]H$��1|W[�jjj��9���V��ʙ�zR���HǤh����5�X�M���hnS���f����LUi���b�r��Ѥ�@Why�]�q�2�/������6��<�r�+�!+PͼP5y=�7�WҶ�qv2�]�6�����Uf�N�����ks�D� �)\�3��졨^ *�Wj$#���s�U��q9u�.�;�n�Q^���u�Y[�N���u-1r����I�(UKv�\wM�By��b}��\cF.��n�8�|����Ѳ��`�i�(_vC�@���{���>��]�Δzm,����[T5��Q���I*U-\�����p����	#�����m�Y�[�)ǅ�m��H�2��k����A�P�{Y�ʝ�DI�{��Qx�%��>�m�:m�s_���F�����f��y|��[�,W>;z�o+�9�m(�B*�Mf`�v�[�硻�}K��@�d?>{ r�����'<ٕcI��&�����o�S�����J���x��;��`M��*�]r�WS�:�`�
3.,NXه�[�(�%�37��+���&��K�d�{�����;�k!�/�4{c�KV�m�/�e8T�w�,�����Y�����I	���s/��X�ٽDwXZQ�>�ތ�S@:����/��]���s��ޓ7�	�n��NZ�u�9��1V�`����!�AZO�W �C�[͸4O"��]qɪ�$�=��]ގ:H0�"��אK���q�����ʭٕ4Ųӏ�"��ͺ'o�+���
�]��-U��9���lou�D�1+��.S��,F�7nʼU�N7��1e�4vIm�x�v�j�O�T����+jZ����swMn}7��э+� ��;�h��	l�X�������w���>�]#�}�)6ʏ���hQ�̵t:ۘ�n��䧻�)�v�{vЧ�����:��e3B������A[E��6��5���潱���mosC�����8�]Y[��V.�$�F�@���f���2�S�B0+�w���]y�ͦo������:�}[k5Х���D�jY�����&)&n��ЪN�*�+g��V�q��ؠ�/�!)�U�㔌;A5��y(!Qb s�������}vž
�w��3v���[�n��U�N��!%�2šs�L�������;2'�cw�9Nt�wQ��bh&�j��ӝR����r\ݭw4�V9QW���H>�>�3��V�Y*ϫ&�J��a5ҕ�g47k
�H ��󫼭U�M>��
�`7G5��5ֻ�"V;�� �);H���4�ٕ�@ފ���M�\��	�.'�����;l٨����-V��s.=p�*��ml6f�k�/�f��a��N�7�ݨogIbԀC��}�9�In뤽'3;�]��1{;eb�{��#�ڏ��� n0�
�eKb�ס����6���h��D��'�sLr'�qLz�3׭CS�D됳����1��k Xm���uy��eGb��r��ё��lՀ�m�EB���&�;U�������`Z,M�.c�˸υ�i5�w�o
]��I�;����0[��)zͣ[�
��.�����Y]�r�h� �^to�K���\/��U˘������˗ڶ�u
��ш�Xb���nҕ�h<Ѡ[�*�0�:�jsR��Bw�To{�S��G*D���x��U8J���sSv�$zM��1p��
��n���ȓ3��GJ�=��ڛ���fK���x�C������t��˧u���c���M�!�P��<�9�d����c�vI��s��pʾ�-�ʼ�#�nD`�<hp�L^��H�zHk)��]DS&��r���D�u]37xc�ᔜ��ۡ[[,����3#��%��L���M_4��o%��O[��T��x�
�w���
�{��b�SE��]"E@�yƞ���q
�6��U�cF��L���>�C;q/��4d��i���RT=���+�_8����s�9��ֶ�J�u1o;id��벇U�cT���z��m��v#d�@=4�U��bTܹ�9ͩ��v�wG:��v���E��F`|��f�VYXh�%m���jGC����&�z,VEҝ9<��є@�x��3nwvd.�l�pA�u8S�uӭ�;����\��
Wuζ��,�*�0��WK���,f�L}� A���@�͞V~γHV)̽�s��*��8ˆ��1N�,.��LP��aen���▞�]pP����닭����'�7hb�&��ط�6�Y��Rqj]Y���������n��bڎ��X�=Γ{h6O�J�ռ1Bf��ˁ6>���������aˍ�M=}�.�ef�ʺo�ׯu������3�v*M�q4�:�eu��:�3YO4TB��Sb|ۇ��r��N��P	�{��չ��/����m�-;gUu�sY�:���Ϯ}��Q*C��:���X�+�cջ�Ku�H�|���	�;��h5=;Mӡ�.���v� �]^�S��H�i`���a�?-���#��.�&=�HϚŗcz��Je��䯬I�^�}œ�s�:� ��b�6�*����weJ�����e_^��~wv�.s��;�}J�A��F��3l�Z(Tg[4���� �ŷY�Zx�鷻g&l}�S��*��	I�]�V�bBLvF=���"�jؾ���C2ApKD �v�K�]�{\�D��P���/+O�u�����B�N����6oNl�Ӎ�N�"�R�f$ŋ�w��gb�Q�vJ�L���y�ڷ@�f!��:C-a�¬�`�ܳ���Z��]��>�e�p@�H��ձ�J�ܰ���RQ@.һ�t�[�����ME�Cy*$��.�k�m;w���H��f���Uru�w��#q��޺ޘ�J�<�����n�݅��^�Mp$�1]5v�j��'��YJn ���b,��[d�hJ*v�U��®�醆��TZ����¹>��%��u�P߅k�{����;�Efc)ݗ���t��2���}ӯh���%�ru'��mDy<��0Jj;ӁY�#��5�k)ԉN�N�씵�a4��P1(��/�u�F6���-����rr��q<�93/���<�+���G��i^uNB�PA1.��M�&_T僫@F�f,z�u��ì�ћ$�g"cޝɝ瀟��n��vNU�Y��k\ɖM�h���o�p=Q�OP ��T�`(�wǵgذ�uf�bW�7��+>`I���oK|�4�򭓈	�K��P�b��������Ǖ�8 p�Z�&�b3B���̩��r����;�����<ܤ�I�)l2�ۨ���H��@���5l}�E2��e駦��ⰞӔ�Tu�2�\xV�Ծ��l�$Eb�jX�X{Q�5��49��Z�ҥ壵�v!Qa�b9�
�L�{����\��,p�(,'�����Qݷ9�$���@�M'}�C`/��-�Z����ig1ϳ�[�9o_5�0q�q��k�9Q��r�Ec���BJ������
�{�&nWf������ZHB��N뙛�1=���
��\�kjdO`J
�#�Zv��i��ȳ��R�3�4�Jk�76����0�O�3HSA��
��lH���Y�Is�5)zf��L��;7��J�/��4J5�+J8 �n<<«#Dcchu��*���{Lp66L͆�l�D��9�&r%�mN�LK�#T�8��E��<�Ჹ�ݻ�z�K'(��b��3�xCW9j�t��4d5�õ��z��d����2"w�)]��z��MāV:E��طVcit
W_�3{��O2�%}iAٱ�ȼ�*u�F]hF��y3��'���|�}{{��\�����R9�
��S�N�:���+�J���ǹ9Xq�m������ųO1ww#Ƶ��b���*ն�NX���Vv3��&�r5��U*Ю��7�Y#�u�.��K�7ՃGTc91����]�Zј43n,ϱ��TT�⮺��#y��j$�H@+�&�Z7uvؤ���ۮ�2��c�0-��s^�����]L�C����1�z�V��w�B���d�nJ���styu����R���a��՞;��ӛ�� +�r�(�|���c\^[P�*5ux8�s�u�u�
XSs�t�oZ6˩�+Iw*����̝m`�wk�6/8N��h=(���:h�
�o'W��8&h(C��݄',,-�L��a,���al�K�@���pR��v{��vjY�{�͎�r�S>y��r�-��0M����=8�����Ӵ���	��n��o�'m�4o��R�����9˰Ny�������0梩�>��E}uoo	����l;�7.ڶ��Xrk���>���G��Uw�r�ŉs\&q��W�����J����Â�]*�*���Cc����1�od���N����C�����S��B��W��<%O��z�V]���ֺw�.�:�q�����C&@se\=j�Z�6��*�'�Olio�WV��zr�v��u+U��n���B}A����9�+
�y/�#�hƦ�O*��oX�l,ff���v4咹aZ�[��nV,Y4��x暠�Z�
e��Ù�Lol�v0
��hiәb�}lI�m������452�V�o�ܨjJs K�f-�bvη�7	��)�O,�C�kOf��sYF��0Sћ3V����p_,��
4t8�nոp,�+8�ۆKWb��,�F�1�P*��r��k;�i�,����}�|��:��VGm���99�<��_u%SFi���P5��F^H�s�46�
�9MW�[}x1�0���ަֹ7X����w��֝��Ik5���v����(�U�R��=�J˓�V��cX�=��J��E��3�1;�wқ_^Ә���B�7Ջ9ss�5ΖPބ���\.�P7��Q�	KO��V�lg8�i�t>��"Y�8_@)>���mm�";{���mL��j}��IYFS'zƾq�u@��utS��ɪ�-����R�蜾̫OA�˵ә���]ڙ�F�g%RJ��Ӝ\�k%��I���D�X��<����G�09LE%����A��3�9a���T_
���	)Ӷ���.u�[a�#�E�c�/r8�[[Y�#�ݵie��C5��������WV��pt+xϓ<�Z6+�����+���n�b��ՕE���!-�o�ʴ;�kU*k@R4y�1W�cU��Ŏ�P�V\��㣲n���J��$7��q�S����j�3qu6yP�M㏒e&�^o�e)ر=V/8��:�Հ�;��3ΏAV:�CT�9լ�7�s��Ҵ��ǢWU��{v� �0p��!��"�*o�f�̳���R���'A����Ul4����sR�]���}UÝ�D��1Pk+��+�v����Vm��_Vq���ȣ��wR4^��T��f�w���%e����f��;l�[��߇TR�;�ݱ��l��4�YP@�D�˵ڭ�������[ֺw̅qs�AI�v�+��1s��6�8qn��q�g{�}A�t-�]f�ekE}\��_	���4!՜���L�]X{mְ��0���Sn����u]����ɶfp]u���8�M�N���U/ ��b��b�G:���"�a�<�{�o�+���꯾�}�^�î.:ie��N�_7�[���y�1u���Ǽf,^�S�d�ɽvs��h�F����ӖkRr�����v�EA��l�nfJ����c1��N�E+wJ�oAp��U�@Ej�GY��3���8o �.�w�j*+G�*�8��� ���o=���$�q�ɋ@�u�A7an*\����X����j�V��*�w��C�n�
��WI�cz���>���A�qI}[N��u\�^-vVO�1ΔF��v+��r�#;c6tL9����e�"e��P��vUծ5���R�]�WΫ�)�-3�eϏ[�Sr��"��7�3%X1�*{K��b���=<���i��rꏉ䕡	A$��7\�㏦m��^�-���e�76���,���3_��gk+W�À %/�����@���[����g/Zטɗ����stcMf������3�
Sӂ�f�(+�ΝPӬ�w;�
hʗ.���Z��{SBZۭ��N����ȥ��v�>�봽�t�_)�;�6��c�$ivf�x�q!��d[F˱A��x��5{YK�t�ћ�ώ�u�h�<�Hj�m�[����xz��%�h=�ը�}VlT�\�����pݻ��Z����Lڕq���9��������޳�H��o(u�w�rT�G�f�94M]R�#�hy�p��C�[s�w���{�#X�ŰR�-�5
�iU*1m��[*�V��KAm�Z�� �D���km�D-��[ZڔZ%�2�mR�J�j�j�*�h�ʕ-mmmm��`�"�Q%eUAE���m#m���V�UZ[*)QU���ڴ��2�j*�E�Ƹ���Z�V6��*Ԣ�h�lk(2�eDTF(��b�Qc+Dah�T+ZZT[V������Q�A��e�ֶ����Vҍj���j-e�[Q�*�#Tj)*1DQT���F�Pb1k[,U*�"�e+(���j���T�bV�J�jV���Vڢ����)�V�Z�єQ�(�X�F2�E̦"��E��JT�Ee�j�6�*�1QTU�-J�J���+X�j��+�L���b*DE�**��)��+�nE�)R��*,`�j�q�k
V��@̫�m�
1A�+
�P�J�b���e/Ē@$�'�[�'�\w���]�7i�y����*�cF���N)�b�.�}�/yu�%_k,��;K���S�v�1uK�}�a+��q�5���ǆ��,�<�1��*�hПf� ��/�:߳4U�	w�.5ɺ�ӳ۩�G�D�Br���~�^v���%�˄!0X�����7�^|Yl>���f��u�m��"�J^��B�Z���F{�<�b*h����|0��*���]�n�{h$�gs��nQ���|��<�J�v���z`�C�#�8%"��=I�N��
l�L}^ʹ|P#�Ȇ��!֝#�,��S���r������=���o��?��>4��A���o3�����Qӫn����5z�S,g�2���*"�v�\O�N��^}�N|,o�s�K"�Z�0X�ɏ�e�F�|�#�m��g�����������xVQ�-��b�$�#7�P���-�yX���{V�qxQ�M��A6�����1$)�w���h�>:d��2�a�F����m��^>�A�Z��q�״yM��/�p��R�B�t����>�8S-{l3JuC��<rk^:c��!&�Uc�Ao�j�V�\��D;j��r�eD��1a�U��F�^u��iw�n�]�C��P����|�U��S;���8���mM�g��'���዗V��A;����L��b�Wdݾsk>0Eݶ�WS���,��ܑ�H�s�'�Ü��K�\��}�E��b�R��*E�:��f%x���x�o�(r�z�^�=o���x�Bm�C^�
�y�6�@�:8����I-3>WdrɳX9*mt���B�Tյ{�O=g���V��j�0�ϧ
#CmݭV��b�\\Hf�ݖ�r��f��ܬ���\2>���n�r��M[��Ǘ�, ��\D�R�@j�6S/����`�n�ș�_S2���u@驵�sʄa���ut�<q�=<�	�z�C>�r�T(U��%l:���k�D`�ۭͻ�f������*Y��C�.��!�İ�ux���V�^^�t���z�a"����5�g6��IΗt�]~���r�	�]f�`�����I�yc�A8�v��ݱ��U�llp�	8V�����_B����x���J$��瞛�=_qss��a��"�.�ғZ0:W����S>�$a�YGE�I�|F���{R��Իew	~�n%o��V$���+�j]���|�X}5xi��R��:��ov�؛��5�-ܩ�]��.��U;���ꐌ<,)��4M�n��	���s�L��s���ͥ7��*x�n���9m�M6y��[
��z�ԭHjq��6�n5lZC�\�3k��僖��vG%-�ț�ұ6��epԺ^�C�����Q�8����׶!-�SO��J�Ϧhy�I�1=5��W.�8��Sx��'������1���i5��VR�@��RW�ܰ��Ŧ*ώ9ʏ|����[�H�+��6
27�[�#>�6�˾���6� ȵ�&�eA����4�V�P���܋���i�k�g�b�f+M��=v,t	���T�ULp�R�\,0Vu�R��d9B���W���ͨ�t�:9����ͯ d�u�d�ܼ+
���S�w�:�KG������
�-i1mv���r�߱�tOq�7�� d���v�CZ�H^�,JE�]V_�W�5���I얎�N����V-|������b'x^	cz��56�L69U���� ��4=Y-H|;��lo����ε
r�.S.��ɡo/yY��?a�J�e��ũ�i��(x�s/wז��#���F��P�~���n�.S.fX�of# ������d�1!¹�n@��Ó��'�����H�@�/�
R�6��ݩN!��,���Uoh]1�������v0�j��ǹ)�M��:C�����>[�Q\���$��%w+c`_o@�A|����@5-й�l��$�Y�eZ��.���wdH�� ��� �GfCׂ��Ն:ﵵ:���z�at]�bi�M}Xz�՜����yA�]����|e����ғI&GRρ�l^:�+4'�
Bn}��5>TŜڀ^�`��9%ү�����P�I.���T�"�e���W%[�gg�Z^
���n��&�2�����$����J���ăϻʀ��C��(�7镈��2����{�䆛/=�dv�T��Vk\D��1�\	�w���V&�Z���s�fr+ݽ4��hq��L���V���,��)���X}p8�{�^��_��P��_��0f>Lu�i�j��510MVg�x�->Sݮ��B:��/WiG�k4���ƌ�`�lU���r�r?�iܽ�߯i,x�Fl�p��� >��As};�+����e�)��S�����uK$P�R~� �7�6Z�IX�'�������x�c��}����*��B�85[3>j_��\��>�H���,o
�X��aez���LT�q�w���na����J����X�A���y<Vu�?�����Otl��Ի2�hB&*u/�_e�v��I9`��јjnov��],�c��%Rb�g7<��w�؄ŕ�Ҭ�2��%���hNX�:�Ԟ�V�&��E]�,���}6�N�d�7sV�����VJyM¸��X<U=ݚ��ۭ�}ݜ�z}�T�_U8��:�6P�{=�&��n=3�����g��/j<j������ﵲy���qy㛰K�޻��(�D��S�\����=���4vò+x�g\T9��g����Tʢ��Du�~h��ê����ݗ��x�g%�����a���P�k��4��{=�P޸{����� /����L�	�j�&D���E��=:��o`YK`|�q;���F�)=%����I/�\ƃ�4M��X.�+�����4I�7����<���.�۵I���|e�����Mِ��N.�����8$��n�:�(y���eY��ٽ(��t�&/�;Cje��ď^�Fs���R0{��9[C����5��N�d���)�4��ת;�����	@�p�5+~�q�g��k�6{~�{G�ߎ�S������h�y��j��.׹��2��N���@��w5y��-/k��,��Su��uY�TG#�r����nF8�a�Q�AT[�_+�Ks��l7s�mv^ڜ���e���X�JR3�5�7�f�����p��}}�3��`숆�T:g|%�5�u���X�b	��>�W�ed�Ӂ�j�ة�[�^��}{�6��z��ٻ�`��� ���6�h�-󌼎v��w������62�j�0UDnLW~��q�ע���p�ڜu/=:=��#ۓ7�������zn�>���XͮtwB��U^�����w:`���{.�p@�M��엏P�v�>-�^���ح���(}�$+ �kG���u�-�|e��v��ܾ����0�k�h\�B���"Lŷ��_��z;�4_��sN�]'?N/e:;G��\�9�屼�֪�]�=V���k��{g��U�q�&rȭ�_{OssÔ�"���ٌ+9r��X���n}]<�8�|&E� ��<^
����d��K�tZ�������hn�gI�*,�.^y�z6U;�Y+���`C���=��MũrⰦ� jwm��Plq��Ogj��˷���gtGElE1�{�����-�2cn%�s��j+6��м��.��\:��+i]�jwT�n��i�ԡ�����C���3�Z��ow>���Lξ��>[S>�۰�x�	Τ�=��z:���=.xڽ{�7��[�a�y ���M�S.'�ֳў�&��Oκί5�چ�"�:T�q�s�&f�W:cd/��)�;��q�,SY�,���<��G9׶���[^��zQ{xGBLzs���+���CFzd*۹D�X���6{bU����z)�끍{}X�8��ǧ#��[��o��9B�FO�gg3}P;���wZ��<��cW��-�<�+&M�˾���f����'���0��IX�9��xj��LX�l��m�ԯE1�U0�8p�seW[����=�ϳ��+���i��0����8�Uf�L��"}��ڷ�z�}�I��M�����n�S'fSY�T�f��nmN,W�|VA:N���8��i�H��"�Wge��y��y�9�F-�a�#�͛f!X��v�ufˢ�\�_T�*�ILUX�cm����w(v�m�����:�+�J}O���Ǣٺi���=k���e\�*�򛍘3B��WR��p](2��J����Nۆ��5�\�0�R�t6�%'��|����o���z��������q���2	�\���\��_Du��{�����7=�^D�ɿ��عv.�<�����u�8�}rev�'���{�tg<z�2���W��wL�~y���9���
�40_ּ�Sr��Jn4Ў��7�7\��A����rp	�y��ݹ����MD4�z�纭r��z��ܿ.
D��r���Q�ɞ<C�G�^S�KɣӎnowAQG�_{��$����:�,������$CI�fe��X���2I��$=�t�Y.i�u�x�A^�oL�c<q/K��g��{�`ޔly�lGA����}lk��^�r��C����}�6^Ӥ{s��;ٹ�W�p�8��
�s��z���i��.m��~n�-Sa��P����w���J���^��m�P���	�WI���:_#ر����S}�t�4�o�J� �n�2�a�Q>09��f���}X�>?^�v�t�t�J�7.���x��U^�q�BS݈}���+�ܺT5B��5m�[}:<�Y6�ov��Eo�j��n@�{͓����'���ǘ�ݬ�y۲{x[���+��?�Gk�1x���qe�[̞��jc���jsR���}$�����~9Y�����'�՝0�1���Y��$�O`������wϏN�${���Xs����L�I��@�l�nyg��h\��VV�\�n's�Q�Ӟw�;9_Eu[��wtfG��֎@a�B���Pw���bOg���0���/�$<Ey/H�zsǲyr�����Ъ�_*��x���g�ms^���h�Ғͺ��ސ��gi�o(떇:�����N��+8q��˗����H}��}8����9 ���0�s�(t�V�}�y�e������Tro��s; ��rf�dZ�dJ`v"��%�2�/,t�{�ûݐZ*�_m��S@`��t��t ��c�h�=�`�R��#�D�{y�`��ŸVdR�e�D�^ݽ��8��͌�������/�
W�"�(��t��PT�2<���$i�#�������D/�������-�����N�Vf�༲:1�M+�����Q�`/�,�a�O*�N];N��Ä�;���͏σK�oT@9��[\5���b�����g���>G��d�o��Y��0���'�s��{��g���0<��z�98�^����k)�hvkD��3���&?or��ꔙ���y^�5Z}�k�Vs��ǧ:�/E�q��C�1<P�����u���-�z<��6l_>�W�g"�{V��=��ez�@g�	�i���eߒ�yKSW��^�G�e�v��}��������=^�A������JҲ���Z�l,�p�����N�}$�E�g�F�.g*O7��y��r�V1�j�m
�l&/D��86P�q|�tM��X�GB.0fz���'On^sB��>1���-�)�����j��*��g��f�l����\�ޜ}��!H������u+����g���v�Y��^e���P��.B��31�v��V��kˋ�� ����N���wn���beu@��/{{�fP7��D�&u�Νٗ�Z��Gj�N���>W��a\[��m�E34���4��["�J�T�{(�pð�Gd����Et��4�ecv�$�+7s�t&� e��ʬ޸��:T��ם�(����Gti���*��Z�?]�\���d�2;�6(��[}�w��43��y�����e���]��Q,`�	�.h��c�ٽ�P�]�`�В���2h����e���/�+���'�,�{m�)m�b 9��l�Uw��f��󆦻n�G�[��9,h��+�b8�U��`� ���H�hҏnl�ݝ�=�Wx�j��Þ��j謼�:��w`*=��C�ue��7�牨� �v�1:׻��nY��Xϻ��cP��E8�>�b��r�8X�3�Ү�4�x۽TN��:1ov��;{�֯�n]>J��R�	�ש�;�͋Yco��R�{�[�Ր�v�-���d�պsJ��b�e����1n�y(ފ�)̕&/<�s}ڄ�+�?�@���j�xIc,Ӎl�4wE�b��z�i����;\�jO6�i���R���[SYW�9��gi��7)�){�k�R��`S��Y�dY.��N�3�-�f��6]۫���q�<O\ox,��e�R
歾e���C[ӛ�-W��f��b�ӊZ�GJp��d��6�]f���T�����Lbtc�.Dr��k��OyJ��F��mR{2�s9(��J�dr���9�E����­�IM�����@p���"�k�gv��z7M+��|���ڵ���1^�X�] �-bU����:��q�3�vj&7ʙ�'2�⒛Q����m5�|��� :��=�Ÿ,�k�0����0v��L5���w�(ͺ���s���1�N�]d̨�%�����:��*���>���*��9O�v�LI�����R�p!ݐ��W�YY��5�ӵ�RP5+
��kb��q$v^b�\���{��鳽��`�uV� �ڴ��N\îT�� L�74Ԏ� c���a[k���{��{� aܘ7���S�q����Ӫ�U8��V����%��.@Ļ*�>�1�!��E�W2��e��j�3m�ww�-ܼ9��!t�bf�.�o/��6��5N�ܧ��s��9�8�|2�a���^D4�݋b�'2+�,�2咊#�2�y���AU�Ԟ�s1Ȕ�V��.^��s���n�:�ֺJ����hWr�'S��E)�b�a7���	:�w`X\D��[q�Nݽ�NcW$�96�����S��m�ަ�t�菖ad���݊J�x�g!1t���+���X�f;�;C�`K�c�!i�e��ѥ-���H=���:m}r�p�>�Ջ��U��1���}~$P@#�4�mQV�.b��[J,QUP(�+S-�j��.b���)-b�Y�.7-+q+�e�e��,EX�e�J���c���������R"řl�����LqAlm�PWLJ(�-�+YX�B�[�ȋUq*���-E-F����,��LT�m����YEQ�V�mR�iJ�FeĘ�*U�T�X�!mb5�**+��(�-E�b�0C���D�(,A��D�K��Т�ZfB��iq��b���0��1�ml���U�UVe��jZV.%Qke-�占���T����J.QK[S̳)`�Z",PX��Lf8���h�Ƃ��PF(�DE�lQ�cEW$�,1U���\j�6�QAL�X��+
�����)"�1�cjQTk(�B� ��k[�_H+J�%$�U�ݗ�mi�;����3Z^�6�۽3z�6�����<�xsyi(8���f��it���ul�{�e�}m��3ݏ��S��'<�^���gG��w���e��u�m�]�������{�l����y;8��C#Eت�G�`���Q-�P���(l��}�7�n
���<إ�E�B;�ɽ�X��������7�s�(=���k�n�g�&��������|_�7��T]�ܽ��==bZ��W��׹ ��x�Nu'���ToGWmN�Y�[��x<�e�~,c���n{����jc�+�g�
{-[��{�S|�գ7f���{��}c��'���pbB�X�1�~��2���<��9ڂZ���~��鳔ޔx=����I�Lg4y\�S��q'�{��{{�M]
˕3V)k=�5z��{�*��8��=8#��,�!��8e�bȹ�9�����
�6n'av�<�(3W��-�����UvQ>�j�Y*��N�r�8�I�L���&;�V����ZH��U���B�w�'rWz8V�i�t��6�Lج�yx��iY�Ŏ�H�i"��twv�W��vV
���������RdG���LZ��
\����\�9���E�ώNl'��}�Ɍ�x�U�/��ڎ�c;dS�"v�y*�J���aos���w�O�A*����N�a��ZyMx�k/��g*��ø���:�N�9&��3����й�\�'<I�E��S��E�F�nw�J��YB��`t�0�����|�k�Gl�ȃW֧�M�7&MJ"�n
�r�����8G�0�9���{0=3���Ȗ��ڷ�tBԑI�m�}r�e��@Nܙ4Or?U��%������U�y�RS��CJoK�;�K��py}�Vhc��9�˭�遧���3�>w�u���ѯs�i5pvwb��x����'»ٲ�!��jh�q}��^��e;[>�Y�c^r_��s胶��g��L_g9X�)&�ư��{4v�W5ztux���!���TB_���K��K���Lu�����8QyZ}�D�g{Q�!�Ie�Mp���&�!���:�m��縸���ʮL�7�z�xXS駎���sZ�w0�����^=e��:�I]����g;5�3�/���n#�u=�{�m�F�t&����9!٩�Ýl���wp-�r��xt-�OIl $=ྐ��j�y�*��|��\�E䰞�p̺o=]5f{��Lޔxy�lG_8����/ta
�S���W/LI���q����t�jTw�J����}�{]=CW�3_n�Ղ����.ݙ��Ӄ���/E�aƻ<�S�bv��=]l7�j���&h%�<�� yON���N��>=��7�-��;��T�mF%�����k�b��TR���66�u/$q��j��7�eRW�k�/#�v�������
��v�^���Ӽ�v���Ȭf'����u�'O.(KFW�P�ͦ*�8W�����w:gΣ�	��x�Bq�1^�v_<j��V|4���ڪ؅�ֹ�����=�&�)g��u���~���������>��gl���w�U\й|��(<sWڃ?X���/J (��1c�p�'vR��g�5F�a�/5l�"ޯO���XaA�U��_G�ׅC�6Φ���Y���Kv"g�F�x��ዝ/�9�vZ�.��J]�kuV�r�w#���S7m�>'q-�ɊC����ܴʯ�3f���pel���~q����Mt/�Gl;"��������.>�"�{��N㭟,���<����\Q��L�a��ώ�����!\�Z�ߕ�۟n���p����!�Lإ�p���!�<��qҏ���9��ɫؙ� ��u7�f���gn<���e������6vwU%����}'z�6wF�1�7Se�{����4��Q|�F%1���2W$���=32ʱ�v��S�޿�J�u�"ɽX�I�O�?>:�Xu��������'��a��3��Bw����E�^w��ּs���ژ^��x�bv~�2m���d8��V�0�I���k'h߹%}d���"��l(q�i�5�2q��^�z�GЏ�ۤy0���������|#��C���a6¡����LO'�ì�A`h�p=Iğ2���'̞~��$�dѿrJ��9�y	��������0}�t�G߼��Ƀ	j�w��d]a���a�i��6��X��N����I�CS�è,'�h��:�ĨM�'�6��T=�r�O�>��$��}6~���BeYT�~���[o﷿|��&>�x�2ì'l״4�hMn�3�N�@��'�:�����O�uN�'SL��{��u��P��������	��?}��0�pА��/n~_��v�����iAw�1Ng2�E)�u^G�G�����x���QOp;J�ܪ�)
Wgt�����eY\��A7��,-���pQ܄N��Q��zhY�Z���k���
| Oy�Y�J��Ʀ4Pnv������4!W»����B�g������7�������#��ԟ���N�d>g<O�Y�I�+<���ɭ⇌�Ad�vO��'R�����I�59�N��'�{;�:�����d�ڽ���.r��=����?}��ˬ�d��3Y%d���M�'�8�e	�<d�k,�	�<���I�|`u��,�=�IĜeOܡ8��9�bG�ץRc��d������v8��:�zs�8�~~d�y�I�����X|�{-̬�a�5�C�x���e1�|�S�	��7�:�����w�G//����}����zo�Rm&�S���'�7�u�I�,���|�ϛ$�����I�i�5�T�$<�?2�q�O!l��'YLd�!�׾�/�3���j���w{������~{��>d�V��������ݲ'Xrk�m�'<I��x�L��ې�f�4wY
�>O9�IR|��͡Y8��|u}w��}�w\�޷�;�>d�;��m&�ɫ�����2q��yCL�d�?r���y����L�2w��v�Ԛ}�p����ҿZ�����>�]���=m+�����ȧIPP����H,;hIĝf���I��V�I�y�p6���C���'��{���O�&����OX|��:���i�a���:^�K1g���ߦh�ս�OS�N��d�CÚ�T'�RVN�d���q&٬,'>O5�C�$�f��C�1�'X{���I��=3�4~����x���?�Ҡ���rk���DOP:}�l�'�Y�<��2w�$��k$�XL��aY6����N u�~S^XN2|����ĝd��}�}@p�����Յ2�A�+�G���}z�Q�OLg�;>�Xm�l�1��=@�w�
����Y�����&������9�%J�|�dۤ�d�'̝�������E�l_�1�.�w�Na{�����A��U��ӗ��;-ί;��È��̞��2�' �6�]|F8c�A��B�X��;k���u���CQ���=�|)�o_"���SB?n6"�n^�+�. ���.��]ތ�4���s8ݩ'�;�W�5���E�N:d������Ax�L>���T�>�p���&�w&�q!��!P�'�o���ԟ�5�ē�57�I}�N:��|O�~> ߸�f��~B�Q	�{o5od�	�I����>d5�2i�R~݁�<d��y�I�Xs�u�c���ԜAHw�i'?%a�y�*O�<��}_~|W�%f��7��=	k���9��J�$�����6��a�I��4{a�N������I��{�>f�8��}�$������$��=�d�VC\��8��V����q��½�y��?sw�~�~��=d����I>d��%t��M�a4���}�:�|Χ�<a����ɦN��O�{�m2u��xI���y�SL��4~��]g�Ι|>�۽�|��O�}CL?2~$���>d�&����������Y<d�V�<g�,�$��<ՇXq���I���_}�����¨;Ew������9�+��~I�:o�>f�O�}�q���'�ì�d��O��@��~u�rJ����m��0����d�~�g'��j��Uw_}� �t���ثI�f�_�/T�w�P�&�P;�삓l�J�C�p'ue:�N����m��s��a��'5߼�����g�%d���>Jɉ�?m��?#�Ћ������pEm���s>�;��~C�t��)&y�P�&Ұ=�"ì�J��� �u����:�w�u���2wm�z���Y6�m�����??|4y+�,��~�K�+��1��8%d���ve!�<d�k)�'�1&2M��y2q+_��Xu���=���'P�]�߬&2w���i�9����ő���o/ҰA߂��[ry���+$�w�2J��C�Ӭ*N ���u��R��I��<��x�mћ�u�������N2u��ݲ
s�g�_�u���}{��}�����S��*�&��˹K��c�<x~�-�.�����(<���{�6k����>슆%lP
*ǣ��b�:������/�����hݕr�5��j�Zڀ�/�r�:G�!�M���lWJ��JM�tc$]\�/�֕;��j~1�'3��u�J��z�${����������6!6�?���+$�<9�IPP�>�hT�AH�m':���M��xj���	�k7��N�����q��l7��F��>�mR��ֳ������ߵ�,����$���N2z�O��!6�2k��Y'�J����͡Y:���(a�M���M0ݲN3����7:]}��_������i���O����I���p�'�&�B��i��g;�u4��M>���d��`)'�J�$�}x��m+'�P6ì�|}��׍�R7���4��{��k���}�p�V���0����Hh���d�z��w$�$��<d����a�=Ag;Bu̝;��u'���VV]{�����ֿ.��{�[��w�+'��I�'�M�&�,'X��4�d�'P����&�h���$��y����Nz=��N �5��*I���T��9����^u(}�_�=���|���C�?Q�}߇_�d���):��_���d�!�p=2z��?o m:��O��I1�?s'X�J�w�u��)��~���9�g;�o��Ϸ��~�1�IP���!X~dߔ�h��$��'t}�,��Ru1�&����d�!�׸~gY=ağ��rɦN���gXM�P�{�߻n=ߦ?��k�����Ǟpٮ� �������&ҡ7�4�������0�a�����̓����$��N3hM?�<O�Xq�z�5=���a5�?'��aę�����y�}��w淛�0�M��9�$���4�Aa>g�YԜed6{ܞ��'�Y?w�̛d�޳�I�M~���O�:��3�ﰌ���~��?Q����mG�L�ׯ�����y�c0���a��'PY='�`!��A}�kq'Xk�a��$���Τ�+!����N�m�'5@���������~|6��h��?}�o6�)�%\N^�ʟفQ���� ��ثx��*��\���J�\�Xu���Y����Ys)<:e�nryX9��m6y�/�Y��*;z���]ȭ���i^�����jv6;�ǽ]�:�J�y;{��;�0���p��4m�۩��?����X��3���C����T?$�eO�ՇX�L����Ad�{��8�ԩ����:�G<é��=.�u��'��d�'�y��'Y'��{��o���v}������Y�Β�c��u���B��:��gM�S�Xu$��:�!����d�T׼�N0�e:�u���u���'��|���]��w���}��߼�yϟ~{$��'��Y'Y'Ό���!�����:��Xa�N3F\d�!�&�,:��m�ky$�+�,�d�7�� �u�y�k7�y�z��X��鞞ﻶ���$�����l��s��'�:wY
�>g�<�+�Ka�+'Xy-!�I�hˌ&�q5�S�I�Y��q��}}�����޽�5�=���~�~��;�~d�&�Y�삁�:k��N2x��}�>v��ONw+	��&��	RO�̲V,&��m
��ZC�8���I�g>�����[�<�\�������;3�C�M������d����a�M�����I�'����'Y�OXi=��!6�d��p���<�*
>�Ь�J�w��>�{|�7���o[5������I���u��i��6�Ϭ���u�z퇦s2z�h��u�OR|��Y:�2~a�Xx���d�C~����=��7��{�����7�����f�%AB~t���*N�P:�l��XN2|�=��2N'�����n}̜I:�w0�$�rxɶ�9�'S�O�,���=�y�����x�������;?{���$�޲J�$��ԕ&�Y<��'̝|q����߲z���N0�9� �d�?}�l&'Xk��ԝI8���~�����x�^���~���zq��)����|������2h�x�:�A�rJ�����&��<�N2|����d�!����&�8�����M!��>�>��`��ڨi�*�&��w�4)�`ǽ���n�֘^� �����s���_ar����f^��h��aB���Xt�v.���Mm�NM.��;�u�N2��&]�g���YSo��=��K��N;��,k|�wW�ء�;����U�lΧ�?�?}��������?A�a�N �59܂�>J�Gy�*O̞�2N0�oܒ��Nj}�,����(q�i�6��N2�s������ˡ�����#,��C�}�}�}�	/�i��}���}N��LN�y�Y6���s���O�P��p���O?k��N�oVJ�svO��L���y�>��g9������y��=I6��i�XO{��i��I����'P_ܤ�����Aa>C_��Y8�	�l�M��ʇ��@���&��>I:��y~��g�guow�����v{�q�O�>N���&������gǴ4��Oo��N1@�����:����a'�:���'SL��z~�d�T&��� u�R>|#�G��o�������d����?$�O�Oԟ���O�S,���&�FY�I�+<���ɭ⇌�Ad�vO��'R�����I�59�N��'�w�>k��{�w|B���NBs�g��t!��~����k�'Y'�Y���i����mI�N2�?&2u?e�a6§���I��d�&��IĜeG�w���V��3�{�t��w���'�>a�ߘ}�$�y�u����w�8�~~d�y�I����Y%a�!�h~ed�!YɌ�O���I�MO(q��o�������M��m�K�+y�u G�E���'m�4{ܐY:��|î�N��^d��d�'�rI��'|�q��}��*O�KC�+'��[�:��{����~ ��n-�������i�~U�����yC��J����P:�ߨ~��'Xy���d�'�{�6�'���a8ϙ7�d+$�<y�T�$>�F��~�<��?w﷽�y�;*�H,;l!���х�|���6�2M���u���C���N2w����$�k��OY<d���v�Ԛ}�p���M�����_�&�$�FMf�1Nt��3;�:���v�.G��x�"Di븈s/n�#�v�~D7=�ƃDx��|���&�r�R�:l8t�&op�]�D��'J�%��c^<��4�G��˕����x����]���,���}���~ߞo�u��
�z��=�	PP�=��VO�XyhIěf�)&�u4�v�8�����'_�o0?0��!wgY=a7��l�a�����������{�����:OY�&�i���I��&�{��N��5��(L�^$��J�P6��6����'���uē���a��?��~?}�@��\�buOk���?�Wݜd�����2i'�Ns	�i��,�y�	�>d��`,��xsY%J�g��
ɴ��e':ɿ)�'>GJg�/.��}��G�e�����˞�{����_�|ç�����p��Y'={���I���!P��4s�!�>d�}��IԜՒ�I=��d�b�������h����S�|=��]uߧ�޻�vC�N�~ɧ�OY8���d��&�j}�u�T�<���Xu��59ܚI���܅C���Y�}�
O�<��O�<�������]Ǩ�?z�w[��G�������Z��O_��d��i�4�:��C^٧�&�u'���f�:��o:�1+9�Ad��w�:��)�ORq��=�0�I�'|���<Ϟa�;���������Oud��O�g�E���N&���$�����L�d<����u�Ԝa��r��'�r�~C�6sxu�bx{�:ɴ���ޙ_q����{�o�w~���0�Ԭ:}���Mk�$�d���I_R|����	��&��(q���MOl4Ì'���ɦN��O�{�m2u�}�	?!�8�^���a���=��;��sק���w��l�J�h����'��7��'̛���B~`k�'�x���XO���4g'��:Ì&�XbN �}|T�{ߜv��t�#��~������� �b�}ԜCG<ì�I���d��	�i�N2|�I�,XO^��$���y�&���!����'SS,�$��:o�������������PN�r������m���l�:")�Vvda�T)���E�������6��y|$���6qy&^V�x�JD�^��������E>�Wi�)�'j^z�y!VD#k�N9n�6��k�G{9R]�I4��ձ�JU�v��VK�]��s����SrV+3fƤ__nv�}$�֡��^-����P�}4�9�O�?=������msq+wRj%;t��^���
ڱm]�����E
�-Wo���ݖ(��.e*Ut'�bƺ���fYns��*N<�ح����u�w,F]]b�����T�\z�{;X��/Y��ʾJ  ԬIQ��Г+�����կ�1
ǒ�V���P+���4�u�P M�`9 ��wG�Z����dTgeda+��Y�P�U����3����e"��5�z��߳�d���d�B��J�q�׊�J;�5�qj��M��ʃ0�I]Z�)V�g�=\Q�ުC�΋�+5rhky�A{��:Α�	V�q^楋[5���F&S!^�X�厛�v�1ݗr�t���B�5d7V��
��;)�G��WY��.�?&E�ݮ�x�خ���i�͋C�IJ��
iTW� 1�9�/��;��G�7��b��D�s�.��f+�8���-g]�$*�kApe��뭉uۭ���������Z����@��-H+ni:qv����w�X��C���l�_Q��mv�;%���z�U�D�y�q�{���esʾ�RǩВ�r�LX��sc6^�:�K�7���[}[�p|�PͿ�v��\�]!�8�4���V���|y�����clm^��^
�J��܉�tv�`=͎V�c�A�x��h�WkHen��(�[b���^r؇})r�i�vd=��݁�u�Z*�����<���]CB���{��ՌԏR�Jyx)�.�B�#A]A�mp}&by!G�K�����,����<��_��i�o��MF�Z�R���w6�t�$v�0|eJi��{i(+��4ӹwfb5�v� X�6C��R��_J�ƫ=ٺ��7/�C_�\�U_w�D y`�
O�.77#re�C����J�(N�dM��d�]9d�\�S�F�A�{OW7&j?-�4��O���Ѽޝ�M=��[�-�r��ˣy�hx�i��84u�B���&Ї{�t��R���꧘����ך�b+��Ž�
�"�=f�蓔��k ��w�ÌZ�������:Ai����L�H��Z��yrɳ�z����MqK4=�+O8Wpu*=dV��P0�U��������
�ʧZ������f�]��ӦL2�nsО�D*�kn�|֫���7:�R}n�(n�ծ�y6s����(fv�'J�Qa��G)u���e�.�Yvt%���r�5�6����Z��{��N�Y[;9�Hɉ�ݠ0��]:UK��a��X����Aq
*�QE�ю0��Ʊ+�Ԡ�,��IUc1�����c��� �PU�"�b����
��EX"�,FJ(\a�Y�TUE��Q�(��6(�TE��Q�1�+"��؋Sm�4QAEc-��U�j�Ef$��ҳZ�PX9kT�*b���[Z�F�30��,U����k-��Ո��TJ��	r⪵TEfP�a\B�E�P�cm����̹K+R��mY\ɈV
EQ�E���F�+Qe-���Z�"Qm�l�QT���+�`�UY��T�ڥEQJ�U
�i11�%ˊ$P�%�"�2"�9a�iF#��X�1�2ƒ�Ŋ�)TR(+i�,YR��`�"������԰AH��Ŋ(e)mb��S�s�8k �P�w|��s{�o��NZP/q���[E-�K���]�#w��]�ķ�#i��y�w3���m����d���]y�|�<��?�b
I�����8���l�d�Vn~��N��y�Y��=.��&��'��Πu��?k�y'Y'Ϧ{�VOX��VOq���ukw*ĝ~�sՋq����}���O�"?q�z����RL>��q+P�xE�8����A@��N��:���:���O�?v��9�����~�߿WZ�(r_~��{�M��~��?%d�O�ٔ��x�ԩRO��?C�O&�L�C��J���ad��ݲ'P��rw�	��;���X��ΥAV�~���o6���;�	c��o�:~��N���$�>d<��
��,<���u�����i8��P�<I6�7��'?Yo0=d�'~��Ͼ�#�,�m_�pH�U{U��س�S�!o,�;�����o>�7��ݯѝ�����M���yqF�	���d!�a��>!��ڰ{b���}kUv�sI]���ާ<��; ��E�Ȑ����x�X�6�v�yf��ׇ{��Uܾ�r���u/������ɨL��[g�w�mx�m�bXO�J
�W����	�#��!�ʪe]I���Z/*d׊u�8��^F���9���Q���.x^.�I2���ًo%�aؼ���m��� �J�2dz9��1Z�c`�e�C��0E�z_m�҅�Rf�|��ux�X;�c�rM���|�������}�y�3n-I��̨����ᚧ�6�u�2gj�2.�3������&�]��f�����<��;˘7�/� A��[�
�c|=����ڹȧ��y��Y��sT�r���9E�Ӿ�N��i�v��g>2'�̼�Ívy/��X�c,4K=��_��z�SE����L`�H58��&v˖�=�WyxSެ�ۙ��s��5�wfئ��dnw����9$�py��x|2���s�U^������ȷn��W�
�C;\858��0��g�H��+hR�(H�듔<�q��P6S��,��{՟^�
g�79����|"�q���Gt\��t��ӂq�_��ڳ�p�y<
�!pu�l��$�v˷]�����)�rtz��ޓ{ہ霾�룸��a.j.66ʵUm���6r�fw�n��o;�y8{g����x�g\\��7�<z�X�\���m����8���}�k��sˊ4��o������0ɐ��D�A�h��S�W��^���V�W�ܿIE_�{��FX��(CC�t�ma��<�6:
�+7b�Y���MQ���΄v�+Bn�=������ۇXC6pi{)=uX�7W-��@�䦬]��.=�U�$��,��u��>�}�6��Q-�Q�w�
/����\��k7�^�j�2#�>��xւ�I�]9�������=p�}t��6SC8�M�.�[�@��]�Io��\$���O*�݊R��	�ս����;G${i�˱�I� �:����eh�����\A�2�89��ag�����������c���Fǜt�L �}�y�aǢ/}Me�(]b~t ��v�ɼ�r�Ϸٹ��g)�ӊ���p��=9�m�z.Î�L��e�����+�˟T�_b�Y��51�^��^q�2gi�緆`����Ad�p�R�{�=��{���VYx�'k����^h7�gݼX�f�⫞B�s��Y�ޅ>�
��=��v�+ϔ��\-�v�sS�+C��[��d�P�-��f���M��ɖ��������1z$�(�ڴ�w�bg٠޻aL�/9���	�Ԗr��7.��/�B���,:yqV��v1�� ���@V�%	�k����+�VŹ�����B�M<��a�;���&�k�:�b��#�ˁ�nӴ�B�]�8R�;$�@�muI�xg]u1��}�KS����ڦ;�﷣N�Lu����f��>1����ع��ɰ;U^�=���c�P��K�s�09���D�R;`��a��u���/7�H<ɚ�z����\��;�����E;]�d��Dw�������u�֢5o�9��g�s���B���NF����[�5�C�3��e�7�å�H�8�fOa�D-�Ş|GK��d�?_ȞDZUd��5�
{��k'ݜ�c�H��DW��7\�
u�s=�x��$���
�Y����=�Gaӕy���9/B�%òW��Nu]=}>�P>�5�]�T�g����8��e�Hk��تy�5��{/5>�2��8s�:��rb�Ri\����?}�E�	��L)�_t���J���-u�-,ݑjXWN˦���f{��Lz"���,I�!��xw���\�|KИ�/c����䦳syM:��NN��Ք�
kuG��nںġ�N܅�gm�ݎ�=E��'�i�p�t��!�+q[���u��x���]�4V��Þ�5qp�H<�6����8K~��v���q煞k_�����I����&l����ߑ����+F'k=1�����/�AUʼ�]S��?+���ٝ��pt��[�漬�T�,N�]�O�P^t��|�5:�����~�)���)�z||��r��֤m�؋��kw+=*z��/�5˪ab�~}�|58�w���zI�����r���iP^'�i�Ʊ��g+�3|(_	�g	
����)���c�k�����'�Z�o<
�.��9 �P8��Loס³�e|1��t����q�i6im�;��/^����������kʕ���͌bL�� �ɪZ��o{����S���Pn�����gl,X;"����U���<9�E}QW�y�)�t�b{}��<}�j#������<(s�����y{���V�oA�ϖ`�ٲ���<�#�^��;h��0�N��Wx�=�o8�Ǯ�S���ے�`E�Y��
���/ �h�P�4�-��kt]��<�c��$��J���ѽ��V�#���>7��W��7��k�P���������\Pg�kCZ8�4�^����&�M�݅J���{��������M����������vO���1�Qgaq{>r-X&D�4J׷�Q������}�W�3�S޵slf�hg^�q�Q���� ������ᓺwb�|wF�D���b��_[���{�kv�t��2��&��wo}�{��׫,Zֹ���D9�k=�U����'��<-z���w�V�7���O���D�=*3�j�"��{"��C����/P��㳦,�!ƹ�;���c�tI�NϬyzr)��n�>Y]��\Z�I�nى�j��K��nrc>��H5y�r.��M�ҰR�=�pL�S[�b����`S�.��d�N/����P�'kY�IK�q�������ٯr�F��+ܕw�c�/��ßjq;�`=;��c�|~:�sd��}��>0E�3k��B��VWB��ecs���>�y�!���]J�:�%Wp��__|@���Z&W�cz�%�B�2�v[���a����hR������s��w���|7�O�z�Ӕ���q^�B}9Ʒ�v2�os�SA��c�gz���۝�Mh**���)���ʪ�꯼��H��$%߿>彞O��=
�����x��ysf��7}.%�i$�{������6&�/{s�r�gl��`�d��d��@�k@���Ɋ��O�͇%���o;�ys����vF�`M���T�Ͻ����{�F�R���4�;\哞^	�⋭���ޱ����-�QOs���^�(��
-qw�gMρs;5�oO�}�q���z�Jƙ���	�51�a�@.�I�{bv=�f�
\z��e��Ӕ[J���6;
Oz���~��h��Y�S�j���͏�>P�k����M�h�^Y:��l�~�έ�޹���UxL�ò����.58Gm[m�$���vb-�d��7��q0��ϯ歡�q�e�:A<���O��j�5@<�afL��q��8��^s��<��t��H�曵��*Y[�M�E���u�����J�K[㯴⢁罭�^`Hf�6J��z)t�=���`�,/pR��D�%��� ���K�\�P�C-���3ݚp��4l$-"_7D� �՗X�N�Lu*�e�gh]|�,{jwL�t������Tڛ%��»���!]��v���51�^��^q���W���oG�������+a{�S�Pp��~�����av�0yl�o$r��+�W�*@��Sptw{w:��X�a�al�O�R�T1���ns#x��K׍�P�y�˵ezm�Iۗ&_����,�i񠘼;��ѷC�.�'c]���x'�w�s������^o�c��8�e;yR�T�����΋u>�%��O!�Z���d�΁�z���_D�
GSr���~�wX�]���m���B��-�*����7��Z���Ny�q|�Vw�/r�戩����2�z}�r�<,�P�u[2m	�F��y'��p-�8�雜���6O�ҟn�ђ���ʇK�.-wOo��h��H�?L�ەo�}K���|=�پy��� �;CY���|���O*~P��,�ZQ�5�{ �Z�W����e��U�<��C�9|iT�Ս[�Y%(¶�
��k��f��m-A����>��6�\S�l6�W-c��&��]�|�t��,�L��w��4;K�v#9r�WO�<�o���������<��A��U��[וpr�C�hϮMQ�5�7Nu��g�Ce��o1Y�{sGW}��a�G�)�xo�M��`#@*Z��VQr^Ouȸ^��K�����b-�OH�|LH^�=}g��fe�W��S��uw_A�8֎�/0�b�z7�M�E�
�8�E;��R��/��vl������}c�+��r-�<���,����Lk���:�<>�*ǽ U��1P{}�G�N}�[<�ע��}Ob��mɗ��Z��}������z��%L+�b�.�^�||��y��k[�WmVĩ��etA>�<9?wD�� ����o1�S��^�����3"+�q���ۗs��l�j�\�e�z�eA�^��88Pn:�4��c�k�7�E�kN3ӝ��ܛ3�ʃ솺�YR�Z�Tz9���c��:z��F5>�t�p�x7��
*&|�+��-5�Y���!ZT�}�:m�mB6����C;�bV��'��t�ٷ��7W!��=�qAx�v,��h)2�l�K/��o�X����aN�s��n*H��aӄ�³�:M��2��\]�:�)~ >�o{z"����y8����%��N��]k�61�3 �Sw^�N����ϝUvW��I�r#�������>�����j+��~��s�{���� �(�޼y;��4o/��!C��Os}���r���y~�$�j�߫��<���\S��g$�;�a��Q��}���=��e����
���e�lTY���%�I�D)�zY��f�I�I�W���8o�.��f�k��{��.>2��$7�w��]�J�4se�����#O&݊~�ts�:�zt��&�I�O�k��
AnvT��N����C���mv�D��=��(�'���e^��f^yB�û̌���A��6��@F}m\C��Z=��n>[�v�u�Wc�,�1�sr������+~�8�&=9�g޿Ovk�� ,�A9��vᗤ�|��ž|Fen��ΐ��X90���&z��3�t_X��&����e�IɘSY�%������:6o�7����m�8���jD1ܕ{3t�j�H��T��p��	oN`�FϏ*��`���_q����]o.�G��mu^��b������m�O�ؓM�V�Ԧėj;Cp=�)m�\r.�Ctd�*���@P5,�\X��vx�v��%���Z�w���5qc�F��a�3q�ڲ�� .�-��Z�וU���U�z���%ey����"�ů+���1�F�n'����ɻ|0��>v��t�h3id�+5��K�T�i�r���h,e��a���T/8���Y��v���z�Y]�l���1���:2���Ě̵w�Eq�{��L��N��.�w$�y�s��T�r��P�b��t���T�&U��*�ͻ��	qb�֟�iղv*tU�{u�L�i|ڼ�RQ�q
�M�O+�ǌ�3z�hj�YK����+�o�d�V�pN<Z<�0g��7��0E�쩀�%kYmΗ+^��a='�\/A#e�n� ���)[���!�-.���e���';3T���me�]�5��ǺJ܋�S*�F�h�I̲GN�t'C�5ݽЉzv��q����I��U� ��s~-mX�P$NJ|�h�sY�E6��ҷ�Yi��{��.f.�1��ۯ`ߘ�2���q��3���զ��6H�c10&�7�f�I:�k퓮v�ƠZ�R̋e�F<�c�JؓW��J��7��t8�����X��$5y�Z�;�쀷�8]����1OLZ6!R��b����/�T�e�.�4�p� <j>��#PN]Y�bݧH����WO�}q�`gT�C�3��j�v����އ4Zr��4Z�-��'T��k�r���'B�|1-u�v�&H�e^e��lɕ ����qYz�7�n�v���/���):[�7�����X������%��vjЕ4a�t�>���Z��sy	v���D)<���Wz��+�=�L�V�5b��+�*�אA(������C���n�})�f���W*JV;3q)x�H��a{�kc��;�ܐ%H�i绎C|w�{V�T��g,�4��9�ʎ��<wa���Ѧ�������N��"�̿VE)a�z��t�K�����0SBwJB�k'��o*V�Qe���/	;�=w�yU�F�B9n1Բw2��|���D�3{P]�.U��JS4�SvV��:��z���G-��' ��}�:�9���g�r�oR�ZwZ������v�w���3W>�r��q��鑻�j��]n>��H�.7z�ć.K�w-^����{hb�T�]�Y�o��w6��L&��4q�Nw��ʓ�Y��\�� �b	D�G���y�P3���zM\l����E��[n��+@wHS.�A������{EQ`�R[j(E ��F��Ơ�%D����
@c
�!+��-�X�!Z�J�I*"��ATƲ ���VVV	l
�I1�%��m%A�Q%V
#"*��PRXJʁV�#[��"(�*V1kQJ�؈)EaX*�U��Yr�� �� �E-�����+�ʕ�T(�ib,e@�. 1����@QDAV	l���"��P�cjª6�&%U,�bZ����F��*�X���"5�(2Ъ���1IZ[P[l����TXV���Tiks2LDKj�Q�J(��K�G�{{ӵ�wf��:yQ��l��ڈު�W0�|�P�j��˷�n�j;���f�4-1vý�ec��Qv<u�;[���|���isv%^����z�p��j�_t�|�<2gn��&�峉w��n�N�}SN7�3�u�S��]���d�����^�g$��L���n�^�'�<�H�į%��T�ح��p���R�O=��,�tQ���Vȏ����6o���wg���b�C�86F{�^Ħfh]&ݼݯ7��A4�k�����ƅu�U�Aκ�:�+��x�}�8��c�� �rl{9�bY�tv�(�i�
�4K�1k��ڠ��B�e}�o�	aM�y3{08_(����*p�y}���G���;"[d�~�(l��[C������xk��Nyy2<Y3�J�������R'�6sN*"��<��:^��y���v�s�.���"�&��7���njC�KCY�zu���͔�q٭�n�X��Uײgg������9�7YW|��{"@����{o���^�62�\P�y�	��{Fv�LP�k4�9?
��h}���&��]r�i�d�i���U�WQ�*R�T�fH���+ٸ�v���鷨o]⮐a�2q�G�}���Wީ
~?T�^�>n-��%�Mk<n��B���͏��xuxM`�Kx�x{ӽCvk�Ndy�2�R�r{~�q�gT��q|,��]�L��>��E���3zQ�����L �~(F}a�hvuZr8=��9��y�c=*.^N�Y�&��czq}h�8 �=9��6�N�g�����WK�݈��p�/�=��C��Q���Lf��>�|� ��Ji�݊&w����ᲊ�.j(>?�j�//�5�lo��0j��c!���Ǜ�ݪ�0������n|���W���L��t\�c{��uxa�S�<y��5�`j;��G�$�˓/�f��y�ʖ��aw>�|<㔳�ĭP�3�B��N�L��}5�p�s+X:u�o$�>x��gj�=Tc�����}�Ns�|\�ޜ}�D����L�zq��ò��N��e�����	��L�%#���ŔGh���R����:˓!�zM�,ø� ���k����6wg]hR0���6�C�Z�Ӌ+���x/���C�bj�,Ɉދk��.�bwS����t��~�磌�NQn7�nz������֮_l�I��`��w�s�쫬��t�#�wѣ&��̃�����ŝp�~�u��?n{�j��e���Y�����6�+6�v>�#��d��0Y��P�aqv>]�}�TD���]z�d�gby틻/��b���94�"��a��ʃ��Z�{��Vut�$��n�k��^}Qgaq{�F\��A�h���op��W֌���;�t�W>�דk����S�s#�l���ٗ��~~{ѓ/���%��Ø{��c��"@n�o���L!�_*� �X�U��*�	�.�[��[�j����8:~�{>�Q�NM�s�����	�3��������F):;ۧ��Ks�U��E{~Q�ZW�&^�]+y)��c�u&>����U���|�=8#��[�ׂ��
{'����%��cf֚��>�0+�G��w,,�|cd:J�M����W�Jվ�X�
c�"X�I򷀙YR6'}�{���L-��y4{k���jW����i��iU��]O� �.�=��M�z�e���(L�ʋf]p��	��ʫyJ�7�e��� ��hS6���-,��2&3W�r��q��L��=�9o��m��cJ�հ�r�G�;�����w˨�ݲ���:G�$�w3w�a�=�y�*��ZxYˋ+KÂ�V��pp�7����rM| (��]yv�&�����3���ǽ�/��Tms��BP�T���R^�evT��|k9�r7j�rބ㷏Nl6�#���W[']J㯋bL�u{�~]T�f��q���G�����B#���,�m8A>�����,#�)�{���>���-M�qo$�\a�Do4�d�=ûr�q�Wcn��N?g���=�9�/&G��M�s}��oͫi���%�w�
Z�/��g��<��^9/�L�1�B�w�˃����q��<C�b���oo��MgK��eE}�{<{j�;�x=�osˋ
�&�.�C�bN«k4�9׉��n�41��]ywg\�)�trU��ę�1�� ��(�ھ���uY�Ttk�<��!(�������T}r�����GWV��AЎ+�JӲ�8ں�Q�9L��I
ΐ� �xnG�y������t˝ެ��[cG��� ��Dֳ�^˧�3�d|�К�ĆU[zunҸ1�Z'C�	���{ ��ez/�d��ʜ�8]��/e���N�������V����F��k���zTg���=R��|�
پ��9��nɛ�No�gxnj�������&=8g���a���7)�!c|�^�R9�wYe�@1m��W[W�����(d������tԳTr��1M���:{n�vml��$)���;�v�0yl�6�jW�GK%'4f������ʫs�ۭ����+�*~6z#��js��;��[8b*>0f�o�מ�G�
l��/��U�T�i���8cޅ��Qg�o�۞�c��_Gs�:��4�,;�h��.�%���V��Ӷ]�v�mP���Y_z=��_�M��z�r���$�)׃��Y��"W?q�w�'��b�0�� �3�����tuȨ9lSh�>͔־W*1.��w��6�J�dMW^�k/:Y�+r�e�;r�b�M��.s�kJ��;A���@�s弫�����>*�f%M����p�K}�B�_�������{��g�cxO��q}\�^x���_�o;�&of|�},�xL�ۿ	�Q]�ѿf�"o��v�ڮ�����5M�rdx���wK�d;3}��}ِ{[�+������|^}���qum�W%F�Mvs�����W\�F�����`y��_k5�].���l��\�9T��d'Yu�k�ˣބvJS������ߌ5�˨rL�a���F���^�uA��\4}@N]�(:=�}�;o�cC�:̬���^JK�Hm�,C�LHÁ��~�@���.�8's�uΔV���|�����^��ҽ��`�����s1���.���2��1(x����&d���9B����cP�wը
�Mk���=��P�P�JԟAB��,p6�y�II^��@���_����w�!ǐ��*�����s��V=��	�n�����Ǩ͐]�$�;�n��{�f׏�k�<�9�zF�ߏT��ۆ*��wcG44�:+3�����s����^�t~��H�T+�'ٌ�b�;�w�J wHQu�f���J�η��uįx
��C�pM\�����ʰ�!����{F5�T�����K�y()��f	.��t�S�V,���A��c�v!:���?\�~����������y���~��m�4�q~^����y]6!�V`LtK|a�9Q�!OG�j����K��O�æ4��f`iL�<a~���P���7��h���S��&�_�*9o1��[G�S�X�ŎgY��������^�t���L��¸�/�-�'Z�rM`�׭�dO|��Y*��/US3�,�a��N4L�vJ1:��\�i����5��k7���w'��m�|�U�p6�-��˲��;�#�,MX���}"��i�OJ�ԄQ����pi���/�C�Qi.I�ikQ���;L��r�S.�a�cA�;%���G*���p7��]�E�k9a�S.�Q*Y� 7Uλ���L�|7��٤�Z�Ǌ����kRC�-�|�D4����;=ud�et�&&&�|�
�ۃ	T�]���A��3��ڮ
���v(W(�Ox��xe��.eh�p��0\(L7GV�_����[�'<֝�Vb�x6���`��WD]f��J_9��9�Uxg�!9$r���nϽe��uС)�����i�]�)��xYa�~�u���6��7r�1�ŗ�Š/G��Pn+dWW
{e��Ȅ�
�TT����'c<pZ������S#�]�72.�n�S��%q�����!���E�O���������wIb~�wW���$��GY���Rt�
�m���<`��f�P�h9��g2��aӂKܽ�/�̿)��1.��u�͟�m�]/.�.�7�y�dv���K���p�;�����~��������=ȋw��B�V&<=�[�i𭢞���z߳�`��zd���]��+��O���(��e=�τkHZ�}�/K�w�2%�|C�^��3(Qڙכ��xn�xq�]i���Z��9m/�p�붝˖��K��;�i��j�{T����ia䧥3y���:� ڠ��s��D�{$�_+�Zw=�-{#|([�.罐�1Dz�-d�+�Ӏ���RQ�d�Kv���X'�.'�.�Zh��S5����5�`�x�Ƣš��K�F����MuOiw����L���_j��ʯB�x8O.�{|w��k^�WK�Ŧ�7�I���q����ט��ݟl�kg��n_��3X�U�;md>��gވ�~l��f�7�\D��#�"����f�G�(j�glf!8i�6��@/wZ����z{�n��u�G�x��t*�,E�����W����æ��Pd�[޷�=�O��)�Odw��Q>g�jW=�I�T(MyG+:庑�Tya�D�bq\�n��u�1:�x����.��� ����j��=I�߾��k«3�لNx,��/{מq3�.�#d�;�DӊP���nc\�<h��|�vԤ:��V �cZ��o,U'�� �����[=��qL���y�=����ց�oRĮ�\Pz��T]P�)�O^�Cx��2�5Ǭ��~�-fl�fu�W������;�G���8߆��tG9����NV}s,�3Uu�'h^y���rmK��,!1��CY]傝p�߇?�����:-��{2k�j�V��k:bu�E@�W�����􆞣�(��!���Mz*b�I��˹V�[/<B��)7΋���⁺d{�zxR�pa��a�OR���:h�h=G2���S8=��̕:],þYk�l�E�[hc�5(Ab��HKL����`o��9���#�xH�����z��=�����\\��Ol�0��� ���<��JƸ�k��yNCA���59����
�H�vi�xka�[O�`�<�8p>"U\x=�/펼��6*��ɽ��W����f��S����o���tKPw�0�͆�Xcw��[��;%Z����$x�=g��*�W{�����WV��N(�����,�#�+��Lԭ�96��f�T�9��cڛܥq�S�y����f��UǱq�%���f��9��\}\?W�UW��$t��;(>}}��eo/OR�c%qxR�,�����`���T0L����g��G���5��z��7c�C�9.>��p�VZ8l0�+�����jC�b��1E�|��@�u;˕�ŋ~0o��A��)��cM�>σ����Q�i�eU=��P�eޕ3�o�V]e�!`C"q4���Y0�Sj��\�xN6=�3����jH��'��v��x��G��U�H�ϯWq��:�^�e�K#R�>��p���;=�ֽ�[�^�]�<���|xȐ,�<�ͮ��@��L�����o8�e��kv������"Z�.�$��ݠkW%���~)��қ��di.����<�t6S��V���a�h���38秒(��@{��7��������s2��m������&�c^)�F��b.霟L�ED���Դ�z)c'f!��׶���p�Y�$���*Ssn5�����t:�8$6Ό�!�&$aϟ��߾\
�,����|B����:�='���*�<�Jwx�2#B`��u��;z3;�݅\���^�d�R����h	��*���2ﺳuZ�}W���]�������﫣��d�~����w&�;�q�4L\ʻ�]k�i��b�slcm�2��M��0@�v�� � ����AR����Z�(.�|��YV#:i�q���6H��;��o% ��+;�ژv�)]�GR�꼭��d�8���2rb��z��5-a����ۘz��Ӗ,���n��J�d�w+
���9�$���3���-9|�+ <�p��t@r�+�	Cv�ME�	�/��{��Ԧe4o�24nZ����,�JU����E�g��G��GE�Ǫ<�w��R����jj�\���鷉9Z�˴)t�,��ś�}�W��=3|ĕ�%��y]Ӈi���ý$�.�"''+���w٣@��-�F���2����̹ܜ���ւ�YJS���A4�h����$�6Y|CՒ����0n�fW}��a��$�3�:��&k�.�+c��åќ�TnU������K"Uud�3�E�QHl�ͤ���7'>-\�Q��f�o+-e�Uۛ)�g_L��iSZk_��ep
Ƿw����Y���Z���[�i�Se���MM��r�QR��q������)_@�f���U��.��Pu]����]7�G4���\���}v�>]���:e�mL9}�=���!��t�����ۏ���wko@�d�Md�ꝣRt&�;=���>�<�v)vg��,/0�p��D;���)Bb,��s�:w���d,P�ޒ";�����3�El.�%��(:���Z������*v�ٜ���\�D�J���8�u��\>�2�`+��R�sD��!1�(�wK�p�o��v�d?wgJ����q+'^�_nw"kh�6��������ٛ���W�Z/�*^���!q�%ؗ����D7C�d�B�'�U8�6/�u�v�E��˔�\���@��0��U�k��8���f�}�z�̽:v����GyP�G�f�}�>�ς�eT�on��DR��gt�}B-��q۳n���#�s��G8L�2]7��u��	�[0l��H2���#��SFJ�_K\�;hi-_��i3]�-�#�7n���Opi�Sh��G;Q�2���*SO���Q_r�}ۻ�����8���;�s�-o�,,�F��T��o�.k7�6��S� 2PQ�&*ݺ��\(N�f{����pW+��.�*��k�L�@���>q��
T�/ui�N&̤���;uo*�CX�S8������H���l"������!����k/��P1t��N-�,:�Jp;Q!ð�B�k2��F��r��Q;}R�ڑ���܈�٣O�#)��tF�������sSzN}�L����mn���Gʐ����_k^�[�y�Gۄ�ͮm�c���D�m%OP*(��Q��&&Z.1�[ATr�\�����eiFŬ���P��m���EQ`�1*
���U1��\B��F(��QkP��m�R)Ym�TQE��X��.4
�R�V�V
,�5�*��Cm��T�UJ��QUjUeEƖX�.7(U��*��Z�
�V"Ul��b�J�6�UQ�A��*e��֙h�(��U�mJ[H��J2�[U����*6֣m+�h�*�0�-)e�@�0TE(��e��($m*$�
�-��m�Qeb���X�Kj��Œ�(�qpQ�h�ikՅ@X�lh�!�H��UQ�$�hR�4��jKl��}HUB��T�;��fw]ۄ�.�e��n�bU�\%S�K:m�vP���
�z�������(���]�������ұ�U����o?E$�5���F�ƥ?.��^����J$�\"�I���.�K���ɝ�ѮxpRz@^~��tu��}�}�K����9T87�%�/D�p3�z׍X�Q�,q�6z�̸��\p� L5�yT���I��_m�E֪�*��yi��^A����Ǥϻ�I#~��¯{��^4֋�@��m;߈�*[��ux�{1Oqr&／g[e�u�g��gO�8����Cq{�a�|��0O�c��x7Kάɍ_�T�̵E���IPD@=��;��n&f4�V�:��zK�y���#�oE�t�|�]-�w^���(.�����-9��k���u*R�,4��zxB6�'�a�~UB�;;^b�Bd���*��UU�ꈛ]p�����g�ve d���0wK�X�v凋{����>)�,U��X�6�-�Ԫ-ӹ;�]���J[Dz���^.�X$r��lګ��=�`y�X�aQ8N��>�h�Qs<yzɃڦ�f����3q�=�՗eW�9��å>���¦���ْ+�r��7}^����y�Tv�{fZy���g��y���J��k��&�څ�z���oT�Vj乙Xv#��"�pK��8�o_�>S�asP>��W�}��}�>Ny�7�|��.e~������*��Wh��E���H`�[� �G�{��_�����<��G��b�eì�G9�0`���O&s'�0��&��$l,n�h�L�ې��`��(o�}�R=l�"n��PbP��r�V�(��L�U����=�����PB=Y��/뿝U��מu��Ⱥ���0?8�^��S1�冾��۝�u���PnW���TJE��J�)/�+���Z2����URu3��~��t�[�i ���Pnϩ|$e�g@�RK�E��u�8�ګ��:]#VwFmʭ*���Z�z��_x�<[D���d�#�>_<�&}�U��*X^��J6硿ww}9�˛��-!���{���L��\������(���+,C��;�Y��t{���Q�u11K�zL��Z8kʚ�M��;k�A�C"�(t���-��C�8Glj���6.PY|�z�@�bķUʨu+�Ρ���|D�)�Hx�\^H��_\�}T�ޕ�b�w{T��s
*�ge�܅�+Y�̜����ʸN��c&��EV�.�]��-2)S�0[ӻ��I**VI������񂺛u�Wna Z�,�>���	�;WdR󯡮ũ�<\;F���;&A��`���Η�ݸܩ�\��?W�}_W�A;�y��
�ߪ�����e�L���99����G���홟5	��uW�{h�(ft)Ə����>�O�Yk�F�\��Z��L��L��H��*D�Wt!�i��_�}��gO,��ƽ\=�Zg���z��t��p���J�ʨx������mV��l�|]%1L��f�z�k��� �tz]���B�6*���Ӟ�e�������j��!�-�g6��=�6a0��s�g&^���[/'�*#d�	o��ϯ�b{\��w�|��(a��aԇ-w10���<g�9��T��F,����|���)�s]�[l�{L�=H�K�I�֊�Zhu���ڙN�ֲ�����u�l�G�����z��n�г�Yj�U��FB��G�/q�w��O�rq{�{sʆ��:b�Y�����ʄI��_<UT,f��w�,	C�{���6VA��J=��=�7�aݩ�D��"��J���!�����uD3c�M`h���>[}3������b�I蠸;ϱ�-��gL`�����Aul����8�����xF. �={��?=�l�wo|��k��;��<z�jV�+��W'ӗ �����J!S�����j΋���e�Ga�gn]��w����^�����#*3�������>�G,p��I���g]�`]p��(X7󂞥����"�C��nVn���"0��E&���@��3닄�O���5{�XN�R�7��C�kyGL���d)��}h��[�<�ේg��|l�5J�e��ԡ������ Cpy�u\1��3:o.�mk���6z������t���	�"e}��:9�Zd��؄�P�^<���ͫ�7���9��wС�2I��yf���.�͒�g��Ί����<���{-��+ͭ"7��5�7݃���C�/S0�v;��;m��{��☫��H�4�*���~^�ٺhʆ�j{u�hP"���=�Pf;��;�X�W�As��z:|�#C8�����!,��j�Ow[������C�&�yD��*g�&�mC���Bq���0iVYH&��^�5�y���e��W����
��I	�TFح��x�)�b1\�t����+��m(���޲�a��O#b&��E�qr��3ƑU2�hC��������u�+1^;hF�]��oᕵ����ŭX<t��z](&N�L;�L�I]>�xx���cP�@ݙ�0DqJ�ߥc�#n��v��L�K6�jmh{id�S��Q�{Wqs�.G�=z+��[��a#%k��h�X�n�1Vo�����+�ܣ^ׅ~~\qPg��4Hn����~]L�P�e��R��di�u=�v��gl[;Vv
��$�:fD��	�(��{�J�=+���l��c�b���{;�:R<2�.�H��T��������LP�	�G�K�Ո�ǆ��y��Pۜ�oQm�b���^���	�]f��󗒃�1&p	��>�!�&$a��������n�^��M1�����b���Y�o�:Q%�������i��f�'k���x�~]0���[���`T�u�0�U��2�{�<^��9T8��_AB�b�.R��3���]cB��*��w�Ġ��+o�iZ���!�.U,�R���<2���"�'���IVFT��L�ǏO�����!1{��^�gճ]zUe�7�U#,�Kΰ?�zr)^�Yzl\�+ �o3Tj�R�1;��7�ƨw�۲��E������V�rݗ�1�/A{*�2FZޚ�I�ޚ���yE��G�<�������/Ɍ��R��eY�lb8<�\�x�X�t���=zԡ�����VR��^��:��ޣf��*&\��vn*����Լ9􃱌�o�o��ݪ�4�E�/,�{B�]��`� '��Xo!}mՎ�S��`y��;[\������R��/;�& \�d��@tS_� | �C�͛)O^�~z���I�ŋZ,0Wٶz�`�C��j(s�'�ƙ�.z?%��{;;$�wy��p
�t���ҩ,����G����Sl��g��H:�^�Yط�=�����Ok�{C��KMn|�*��|ð]_�D��mITs�'���ގ�f��fq���ol�*P�H�8ޕ����4Ըv(�k�q���b�����76�>�̣�|Fyؾ���3�����(;W=H�uH���KyH`�ص!����ߕر�j�����P�2ǈ�9���L��g��g0O"aS��izP�
�۽=w�d���d�
%�Ԅ�3�?�L̵�az�˙[�<so*_������g�7�a�7�:M+���J��ȮϬ��}��Çƹ}~ݥwE/̗Mn:Y�IY�%��2�x�t��^�V��b��I�Tm`>�}��nO`׼��݀<��k�R��q�j\�Dx(�x<H<��������O���WˑVU�ҽ�:�yb��?V��\����w��2o[\����/V^�puO�}��n��L���5[u}���)7{�E�����[��>�����f�-q�"��۬]�e��{%2�x�vrb�-��ꕌ��9Ξ�/�B���M:�����fk��������7��^k�>��ܬ�}0�,�D��(Gt|�yhL�*����\C=��x?���3rպvX�,�}[�13�_ϮGv�<���_X��pw���~�4g���n�M���LC}��d��Mu�g!J��~��Ҽ�u^�l��COC��"*�0��=^Z���uo]"�}�g[�
�P����0jA�����J��-�ut�s��,{g����qF�+�|\Z)֕�D�",c�	7�:f1��R�>3%F_a�:$��ا�	5=,f��X��4��R�U�,���[�G���t�.Y�J{ӟ��c���UA����v	�]Ƿ�c7��P�Z����6F���lܵv4�P�׻P�X�V��6����-��f,zX�,G�ڱ�׾��zU#�P��T����ݎ{<sӠW����[䄮i�XY��0�VNx,�������2�&Z<uߖ[&1�|a=H�kc�����`�KQ3���-�9l��Bu�3���-�~�X&T#���W��8��!^��i�SF��gf%��f��ՉmS�����lUp�!~�ʆ����U�թ^"/��}�AV��k�#(u{�x��9�1�"��qM�';�տm�O����ƯWjJ�%M����3u�綁��wZ��[��׈�������{{ �������}l�Tt�V*��z��
�C�-;6�u4�O^=��ו�r�C��w�ͷ(�k�Ű��/C=t���yĵ�Üw^u�oR9��Vc9:oLsm��K�R��3��l��B`��U��B��P����DǗ�;Gf���vZ/P�7�̼�L_T��n��!���G�:��%�h����۝9;���kgg.��yY.�h!�۞����37����CE	P�Pp[ڬ�5Ca
�r۹>KQ]`OJ	ɻϱ��œ�չ-0i���>	�B)���`�S�"ZgƵ�Gi�`�5�w���^D�c� �abl����V{s!�;�l�!t�W����5��w$��zLPK�����ZX�p��V�u<�A�q��^������b��{~v:kH�>�����|��j��X�%qxR�.����4(�s�7=uv̝1����ġ���>W�Ʀa���r(��'({��G�:+ţlѫ�a����^Kg��a+L�0kc�z׽+�����d|��A%�8�&Wq�X5Q�UEf����*{l(��w�S�c��nٱ�6������{V����O{̚X��>�C;�OC�����1�s����c\�J�21�QC3��==r�S{��������|>q��bq��w�������q�������Ա���x}���⌍�4���i��2v�=����I�J�"��(i�Q/4b�%����K��	�j��Y�$4��<W���G�,���Xg������IW�HV[�h<}Ճ�b�u)y�lIUEx'7��]"8}J��6���H��+��NH5����}�A�'�>�|9��l>�3�ݞ+�ɜU�T�!�4�Xt���å*\<��|F²���ᵫ���u������Y����Ixt���q�L�6�GP���D�R�$�ʲ�oj[��t����Ry�/<ֺ\}�]4<:K�=��.�Zs衽F]C�2�G�J=�yMY)�g9���+�BiݯA���x*���M?q\�(>1&pHm�%�w���U��5@��;���m��W���0z�n\�p�R/v�[�
��L���vͽM��Z����]�g�V��<�ʚ:�l�+e��"���ʡ���'|f
M��&B��I����@{ܚ�;G���v|U!��R��f��\�
Dq@s=B�C���I�A�ث"���m�U� Ӆ,Yn��|�u���Ug��y.Qzf���m`�m} a{3v�X�"wSO�bmS�=}��{�ya<tFl�;�G�UUUU�<��PA�,_���8㭪�Gkʡo.�Ou��h^*!Uԉ��_4��[:=�w��c�i�.���L%;����c��Ī�mx�֋���S�Y�!9�@�4��6^����B�3�.c���C��Gxm�]��}��S@�b�xÃ��	��H�yՁY>.J���F�Y�/P��8��w��eLq31�2��j��%�7.X��gs�Ch*���������5gg��UL�d��Ab�Z,0}�򋀦C��ˇ�uKx���V��GS=����.k����1�c�f2�`w�`Q.�IY�Kf��̫JWw�\U��9^aO$'��@{W���W�|��IP�|^Z:(�t�J��ʹ��~��uM���r����'c)�%�u��zTFƠ*��Ij\��)�.j���K��,��Zx��GE§�<�|��ib���O��}2��wt�C(qn�^�j�d�1����,X�X�ecjm����s��R��9��L�a�| �;}mI$WMH�t��q�F������gp����}|�O�f��q��ݼ,���7cGdl���Mj�q���RYJ=��p�z���u�uaz�r�s3Lxz�		A�/0�e5�f��N���Q ʭڻBh%8ٵ%�JR���};�j�Z�w���#)��c��������՛z}(7���U�5��ӎ�����\�U��]6�r͙F���c(�wIL�	��WVR���ee�{$(=E�ɴ�N����MSSy�{W�Ķ�]�n�����ps�o��e>}Y].iæ�U���Zs7c�� X�n�aQ�M3�6L��f�T�♮乃��}���a��i�Tw���qeIU�[gy�I+m��ڧWkF�5��2�#�ְvU���r����iq��/5���s��[M�����9t���0�m� ���Y�{�p�I�>:;G�wQw�'��<4�������j3E��R�xD�n�!��갅滭`d�|�8��d��3v��Ϋt*���Wa�U&�eu;��v��cN=�y��s�K����۸xq�F`o+(�s���薯p޷m\k}Lt!��)#Gi��XZMbV��[)��$_^&�P��u���D�����G��z�g���5_VWb��$�����p��˅ M�t�^K�>Y2)+�oJ����%9Q�-\�֮]=�9�/7Hax�<�G����\�5��j����Õ8U�kd�&��˙,���G۷c�o�����u�;Nn<���^��z^19�q0Kݗn�Rg��=���ڱV�;�WZ����rU�Ź>a�l���g}k^.̫r����;7�]��-��XN����e.�_sk��z�Tݎ]ҵO�'SU�t������;�n�ĵ\�yS�5�s��
F��ƾ���"���B��5�\4`Ǐn��ݹ,��Z�5����%ۨ����!��k9����7�.0>L�r&�G+�hM�Q�v��s���X��9�m��֨gd��V�xRl=s�e$Ʒ�2���K%Ѽ�yF��.�W�t�9ܚ�w�&N�,�]'�x����ԕf�GaaD4�9�:����6]����ں�wH;��Lly���{+5gh��2\
�q�7�9	��E�J/uE�o�q�mrV�w�i"n�w;�9b��[!PJ�9Hz��'vUʃNf'�ު���}Emc�J�~8�4;[���o�w־���|�hN3S�F���Y�f̫)9�*�l詇��o����za��9S"�Q+�'�4���J�B���ښī{E��ôw��B�{�V�ܦ,p	���}�v]]��['  �M�X��Y��g�����oU�)������9���)�<�c��w"d��p�����,��lFL����׊��sU�7˽�ҷ����m�V�O��������e��(�ws+*Z�#m��5��Uh���B�IYQ���
�[m�ԬU"��,+Ek�m�����"VRԣiV��D�Dƙl�"�j���b6%jQ�V+�e+kJԶ�+��)D��0�$X�l��J*�Y1�2V��E�ڠԲ��Ɩ�(��("+#ZV�[TA�UZ���YEh+l������0�)K"��J�J����$D��k+im��-�m-(ff�֪�ĥ�QdV�id��EQ����+
��J�(��ʹV--
��Dk+*�b��6�l�-�Q�l�TXT�&Z-���j�TZ����Z�.Z.)D��[k%���֭���Z�¢�"J�F�m)h)m���km���b�F-mm�,�F�P*E(���il����
%m����-�Dcu`|/��#�z.�ԧ�R��͒郖!�lt�i����K��-p��orY���m�]շ�T푰���Ƴ;�����o"�͎^�x�O�J"� ��lV�5�{��ׁK�*�~������=ཤ(aE/�8lX�d���$O���/��U
�j_��~|��ΰ�)̘q�]C�:侩ݡ��xi���^Bug�z�_L����#��^Z)LZ3ǳ��bf>1���=^Ǜ5��u��ÇL��>��
rϩ<H>ˢ�;����#ףcSiޟ�g�i�(�~������+���h�'@r�&4��?U���X���9���7bU��<��WX�ɫ6�{l)\7/r���1�eyǔp̧�z;�P�ɸn�Ud}~Jf�9yPx�;`7ՙ/�g�#5��M]L�?	���}��ߢᙆ>�^�՚�k��k�93Ɋ�ٺ��~�p�g[���i@s���3�H9X��e���|p���C=��t*�Y��\{i?^�ఌ4,WV�&��tO_
�c�	&1i7l>w�.f��ǵm�q�_�ρrެ�H��̞�K��+�����I`󪋨\|ǫ���w��D*�ec�^�5���l�z����k�s�7'������=g*A%x�����}딳_v��*C�F:�G{p���դ�K�����W9I"xP<��(��*�<�/s
�i>j�4��8��	�/i��2�>d<v~��>���ګdڜX�ď��K�%�]'xL.���Fkx�E��-4,�b�:9��E/`s&-mߕ����N�Y�<��7b&1�"=��p|n:Ϧ]Q*<f3,��||�زq7�l}�-�h�S#W�Dl��\����,�xl�a��=2��~r�r�S|�%����e9Sn����<`�4Md���BA<u!�e�G��q|��}��l��ZU�.�fˠ�jĳ�D0�����y�B� }��J$�1����(qӳ���VB��u/V��V�0�0϶��V �̠�	�2���a��Q�wE�+wX���
=x�nIu~�zc���lcgԎj��mz���]��4p#D�,?ZHk+�'\e�����"3c#�;�b�F��{h3�%s���&Z�B�e[D�Hi�>�B2��!�`����n:���כ���$\8Oq�=+~�l�����CGD�X(8-�VF��o�)&<��Z���dL�������nu����^���d"��mD�Ab��s�ՙ��L&;��5cx�ը^�ѯ���hVԬ�z�P9��_�Z�M�C�w�F�"P�,*����Ň�P�����uh�m�9i�ٽ�o�|9�wk@7�"�Ō�#�ˉ��֦z2�+�F�'�kA�9��1[�����Ҟ�{;�٘��g�fB0<��JT�\=+=���=��������rN-f��+��|�D�2V5�O,:6[�k����D~\6�����ν�<�uw9��ڊc��{��8���2��I<�O,��Ա^,J�GH��q�6���&&�m�"��w�w6�!�Z`8=Zy�`�L���r;��Q��NP���Q�LU�ػnM�J���o���^*>� [C��h�g8&Zz�1����96�����}ʸ�|��v#鳵�̫�|b���H̥CHW�[|eR�̩���Pu6��qs����5���2zD[Ӟ4;'�(L7�
۩E\d�v"��5z��`'���g���m��s:\�Һ�IIn](x�^��dw�����F��Ƹ�X�f 1�P���Cvb�3VŖ�J�;�|�|��*@��}8��^Zϭx�֯���@�����A3{P������C<S�wu��wJ�T���a��^>�3�xO$E�;:�AK� VP�{�4�ٓ1�Ce��S{���靏t�v�X���(�%:6h�����#|E_;ʆz�2�����|��I���ܹ���/kU]d	>�+��������{���k^�¥Q����Ѹ�?ȸW���H�b���J������[;[���iKٯ W��_�|{˨xzEn��~��;>.�>�
�9����D���)�w�Q���F��	"ˬ4�]����^�RT�.���YN^J�$�!�tW�$�y��;VeX��,d��G��j-��ͬ/ùY��U ��.���oH����%݃uZ�p���	֍�J�@�pb=��K��;+Um�O�Bpp�Z�5��^���j��%���^kRϺQ�{�|�)�Q9���
���J�Bz��b�RDZ-<�iy���cL_>�M���$��]��{�bT3kƚЄ�X-J-?/�L�\�޺�f+��;k���X`�b�2��t���<���Cv�K��}tp��׌�/�����K^���'�}��q��B,.	0G��L�o�v�z������O1��v%�nT#w=����cC���
���&8�G�/%�,X\,0P�]J�-��/�jfB�JL�m�e�;�
|ϗu�D��zxB5#h��J�]�N���07�\.Vu�١[�#���Wm)���Զ|��먟:WmJU��������ao[��=�[hT6���^L`s���@��:�F;MPq����Э���f����1ͺҶ��iV�l;��:#����ȜhȺ�ea��3��Uy�۳�,�=���8\r�]�W��'���tf�r`�A�@�'	����1������G��{{��)Ӫ2��#��/4K�����sVf����ƇXTF��%�0o�(��l�vn��r�_O+����+�\r�Sk§�#�,�	�oR>��xKR.���`ɯ/�}���£�ݑ-�BUw�pX��/���mM�S�{�D4��گ/o W����*�fb�^3~���ycg7���4L��$�#��(Xr���a�,k�E%�l/؃�e�r�`�t�~�䳏��~+�W�f�8�	�����I2:��lW��}e�r�CWsK��}6�a�;Ōu�*��r4�9�z��*�z�T:R/�J�*�S5��Y�c�J�&>�7��}l���ʪ���$��%�|�R;ʪ��fUJ㞃Չ�VVt
=�رD�nW�)�3�����*ƹ�U��h���d�#�>O-	�����O�����������WN��}�至h\]���\U��q�<g�Խ�v�����^u��I������4�/R`dq����)-�zG>�h��n�hk`k谁���*��gn6��@�/��49`����gk~��;�A-�̇��8V��9���:�9��	/~jr�$��ӵV����^f�����dS��_*���L�瞬�����f&	��LY(,��uW*a��6V}*�.���Hi��٭��a=�=�ӹ{Zppuv�O��2R\0����s����W�A� �!����i[��?E���C=��=%�ܷ�o�b�0�,WO«�MiV螾":��/>�g۷1�'m�v��L�p�E�x��ׄ�%=��g�ee�VGMX�����|V?A��o;����.��@ǂ��>� ��K�/���'�w��{�̸{2�P_V�O��kN�3
�|�X5vW�EV?����gZ?R��=�u�����k�H�(k���]U��vH�6���J�l
�"G:��$_<uY����ل¾>�k,�x���0jk+�^^����se�,�,�49҈�+�7�qw��A�t�՟'X�ռ�!]'�U�pS��9 ����%���P�6:�v�\�D�
�c^��/�`.=6��:;����է��b�vـ=�~�=�udʞB̵-l�A�ց�t�J�:���{�~��4b�w��ޠ��t����"X����pV���Ѿj��i��.Dw*9�ه���Cs���1�N�=�s8U�ءK�8w��pwː�Lt����U�۳��S�c�p�P��ƼZE�Y�Mm��E�7o|�c�����K�Ӡ�nR=����z���v��Z�s�_	��A⪡cY�����"�r���m�٤���C�z/u}�y{�tc2�x��{G*uK�!���{�����M�W,�qy,%�p����Mn��m.P����j���5G���p'�nخ���:�kc�j�����,k������2�.���N�"��{j zz��`.�bY5V����������}Pt�:V�e*u����/��9y'������j��ҟӫ������"|,ns���X�%��Zv��ѹ[H?/��WN��+fͲ�U
��Sk����˅�z�r���c��$���+yz{Z�+�e#����h��%	�yOs�Wd]O/JC�x�i��>���$r:�?�K��G�\=���F�{eg��p1���q���]�#����/�]B�^��9�ˬPf&����C���m����O��L~S���6�ՇE��T1,�8R��]1C�������Qd�}}~c�;���z���i�>�0�Ma�͊T�W��GY�{�	;_��e����w�|�K;{����`�[�^�!��@E���Wǭ�]��R������F��л� sJ��\8��\&rjJ�p-����Nho<ŕ�\�Ҹ�ƕ�}������u�_��h��q�[��	����Ъ�W��(�q!�������F��-}���x�T,�|�9~�޽�I�Ǫ{2*��Dhm��֫u"�<\Z(&e�ݖ��á�]�9���!�B}]��ޙ+�Nk��e�Y�jD���@֮Jk����#D��S�-n��v��m�W ��pS�þ�4�q�>�zfq�}<�V;v!>�Mgv�xP�7�j�&k*����p�9;�s�H��ϺD5�)�a�.���a�G��è���ޙ���m���|��t=������RW��e�gI�����A���島,�=�U��L����4E+^��v��u�B�p���沞.��0u��7|蓜�{,�@�s�����){��8赢JG�'���)b��p��!�B��{sŧ�-�xo,�{=%���6�������%�^kR�ҎY��L>ϵxi�U-e����߁bVM���}H� ܗظ�g_�9�P�-��my�I
LOM{�ﺳ����Y]+vU���V�j	�R���C;I7Ru�F ��`��vVL��+cP�%*q��Lv�j�VP���v`��ޜea})�X���y�CMŠ�e��@l�u,F���.�-�lۣ����n�u�/X�k����>�@��q�s��{5v��Z���Kvs~�z�J��qP�]C��I^ʹ`v-0�Wj�.�k�) �{�����r�R݀��P'�Q��ј.�+0�m,A�apI���ʃ73S+O�u��f��gK �P���a�v��!��x��5���h�z�e�;T��,_˅�
β�VS!�e�4@��Ak��~��@y�-m<Pȡ޹b��xߏjT��i��*��ϔD��p��T�[h�t�=��K.��*�<���'���v�#65�M�U��K�xWU��U�ξj�W�Ýچ�~��������#�!<�%,zN�o>�9��v�ƇF�y&
<��1cLY�&ziޞ�,��H��P��3.��M����"�5��J��R;E\����=��i�Ώ7+؁�H�`J5<
/�֙M���eï~����s�����~�Κ�c5f�WR4�u:[�ZG.�ͱw�`����܅R�H<�]�=�ɃY�����y.,e�*Q���>��C��[K�t��zR�~����.��Z�����P��N^/��ڱ������1P�1 ֱp�M�Y��r�3�ݭ���u��y� \�p4ƪݘ��<��[��m�}�Z��Q�o:���r�ܾ�jh���,����(Ԇ��.L�g���������\��Y���v���]A�#�_}��7��MYe�Ռ�Q}E݌>��6�x9br��P��$�t�^,/��.�u�g���T
��:�E�x� ޲׏�����%WDx�V�v�e���
b'(�5j���i.�س���o�M��k�|7O���Y����Ҧc�S��%Gt|�X�v�nx�7Ì~N9z�ͬ�ы�S�����%�{P�Z�ʧ
r�����q�-<K�9���r��.��6�h"��-[N�V�� ��3ּ~Z|+Jd�Zg!I���|=V�;LFɓ���=���7iO���ݮƞ69i��01��d`���g���ПU�r]z��f������<��o<\)A�ɦ�w ���lC�e�Ҽ�78�b�8;9�������Um\��8�QL�}�p�N�fpw/�)�b!"z�d��Լ��SV)e�A�
R�����ݎ���b�g�£H��b�K�%�,S�%�^�Z3�i�z/�(Κ�I�2��p7���kr��a�.��bP8Yio��C76x�~�4����Y��Q���)R��ln�KW.�w��
�&�Y�ik��Ѽ�_.����f|�=��0'��G��f�B��9i�mU�55eޭv\b�T��[5�VAID/�iţ��u�rҮz�P��mDu����x�pV�j��f��j�a�+!y�kUgK�3*e5'd��|��r�յuq�L�5��R]%��>/1_0�a��:��7���XE��� 0m�Y�x��>�}D���b���,�5��G��b�uLq����nSfAC��q=g���x0�닏��L�OQ����"�VKwPuM�]B�g�v�u�v=��7�����JQ�Ί�!���U�@Ӯ
��SߢK�O�r�v�L�,��6VM}w+�]k�j��ƅ�t�-IO���*LޭD��4Ģ��Ӽ�kT����X�-RՃ[M��cz�泓��a�r��ը�t���an�Q�ݬ���B�E��k �rWVwb��x�]0�e�P��[�*y�`s����OJن�a��Jh�7�_7`4�#W��tv���rr�s�x[�*����
[w�fh�C��ND���:��(v�N�սEgc�X�!�)�r�kV6ZDց\)�\Ψ#;*�C�)�������v�;�`�R.���󘄬޸i��a��-�����g$p���X<$3���t�t�u2�����P�ɨ��kw�o	x�R.�a�!\��i��EZ����4L�7Ut��������H�!�p�R�
�ԅ��u�Tړpho��#��x��9�V�UlK�4�S��W���Ud��}�X���N�&{&���j�\	Xz��r�`�R̥�\u�v����ip��
-wY���c�� �Y��,i�K3o�^�}N�e��q���Rޅ2\���+�J�*��_�N�&v\vrN���R؛!ت� ��gJ� ��o��ù�*|[s+i-�^����Lr�c��N9O�B�(Z/�,���R� �w��]#�:+k1�-h�ae�~=����źK��J�7�޹����**�[��*�г��|u,.���:����O�kT����7L�S2��Ŗ����S{<A�z5{�����j��:�M�]��¢��zì�<SZ`kw��.0�Nfw��4i�h���G{�i�mu3Wi�Ĺ�����c��)������KGPI�x7t��'P7�7A�O��e���L[���k��&�ح^�R�.�t�+�v[��0�ӗz��.�|��QڍrT]ƻP���AGۉa��Ek���m��z�s��kN�[a�P��w�;b��Q�@�h&����(�L;�W���7*�E£���
4�q#�y$\Kn��Ƹ�aj��+�K��
�&,�;y�B���Ӛ<�K\z�8��U,�@�w�p��#���U����'|yq��V5�oC֩avy<|�K�.����j��S���oU�� 1��v�k^�*��uK�4�v�{���{ہ�²��b�T����E�P�*5��6�R�W3[��J�T�J4���B�����+�j2�*DDdb�U�J�2�
)iLnV�9L�J�-73��������j)Ym@Qls3TX��lbJ���-�Բ"ƌ����9s�ұU�P�j3(T��[*%��m��R-TZU�������-�Z�Ũ�ٍ�-)UkE�%E�UŅ�mR�Kh��YR��
�Ԗ�kPmq�3�6����DQe(�`�[m�"��T�-�eb��cl�F�E�X��Rť+RV�SLƕb���`���Q-Ujʶ���UE�0�Ĩ6Z��J"�TR�m��*[e@c�-��(6��2��Q�+B1��@X��*�TQ����H�[,��̮Z�TT���T�kW����Jԥj����ְ���-F�2㔴�Qm,ʕ��s(�b���X9B������9F�\0�/!&ٲ��d���/@l�.��S��K��`�Ս��ԝ�-,��֣rM��˱�]�ܵ���Y�lH�?|p.����Eo�W;i=^,��d�sz��L�!���Y�t�l�|����^	��FɱΔF�\a��Y��+���ךx���K�Z�u[��൲��}�'�vyS��I[��.�4o#�Z\=��d`�49OG��w�\��7���SL�\��˔�S**Ϧ\��'��� y�Z]N�vV���j}�sy�V����+Tny
:�r����:���$�{�*�re��`��UC*v�o�~"+�G��٘�mW�����g ��]��h�-B�UȖ$4�(a֞nR,]�	�篞��4��4&Ӭ�n@���+k����vu�.x��<�:��k"�<P*l�I��u���F:���D5��!�X�äs�h��ӳ��綠�K�I�S)y�8!p{w83�ߣ�:^L~APs���xe\\%�~�$�hG�f�g;{���;t�0`�u�>�m2�ǀ+ظ@+�+Z��)�x+�����c�^�tՄ^(����ƅͫcƕ��x�yt�5\�L���^WqP8��|/&�ct_1v9��F#��k��%μP���w�(�R��7̄���H��5��wb@�7xkoa��Ջt�Л��e�J]w��їԛs��l� и�Ռ� �Zf �Dny���c�ߧ�z����%��0��?4�Y��m)b�V��Ҏ����K�Ln&f|��;�h`�>����;o�s�A�x����,�dz���5y�x)|&T����@s�p�]`���uB�X��.�}�{)��5��i������6R��'J��j��E#)�}LĬ}��Q{'���4:�xxw�R�+I]��V�{B���8h,q!���1%�Ѥ+]-}���Kޏ���"��/9g1�6�*oY��>ȫ��βq�����6���GS��+����!ޗwWx�|�Z���z��19��J�s�ɗ�g��������J)e����Yy�|�1�w�Kǖ\�i�24���ﯦi�\w�O��g��yXp·)^%I�k�z�����kU� �7�R�uL�l�u˨xzEn�t�k1,=���Za��E�1|��o"@��~lή�ә�'�6Il��]'_�H>�=�JJ�E�c��e|�������Y�\���m���K�(��E���%�X��^��=�W��L�E���o��r(�sJ-x��gf1cX�3w�;�ژ�*���ϴ%�Kōbz�T��;ԧW��;�8��:�1�{ ����Κ1�:�w^��Y`'sF:��l/��3��z���ͷG�xc�FǄ��"�[�xg�Xxe�����Y|��6�5�e⍥7�.l�kP���"�<�|�Z0H��_LJ�?]z�Q!Q��C��]H�緶�E�mg���r�s�让>�_H�}�)�	���au��������� ��TvϷ�TI��u�Y��}h���̨{��,�|:Ƙ�L&ך��"��[���	�+�y�����`��M�`!��F���-u����������u[;�?#�,n��p����o(h\�^���Ɏ˞E��m�˓1p#�LnW�.	0p;*���4�V���xø�KtoY�����Uq�PG#|���z°��И�3�Ixa.�z�*{J�7��P��u�=�N��x�5S#9mb\`�i�	*kɂ�/
mҧU��hw�b����P�~��(I+�mN,z�3��d��'P��x�q���6�v*��N%"ϫ��7~�6&�g�[W�-bC=K��H��U�7�RnqPK�}8�ud�c�YL�[�..�qZ�c�W1 ب�"O9�;��b,�{9�z�0�Mԥ��;a�Yf��rmީ8H��k�U��X�
�7�S�N�Y\2�s�,Xx�On=���_h���/�ZU��&1T\k,s�ՕLo�i�_[̷;WU���{J�N�O����V����+$� m��+G��s<"�?a��\#6Q=����g y��>���5���-�R3��<��#A��*g�(s�u&w�n��L�u��KE��1;
�z:�;�m�+1ed�|��Șnx�5�:D�q}a
/o*�X�j�&z2�`�����OS���T6|qS��|�͞�OJ^�"��x��Ԭ�w��{Z;	W�����}������V�{�=<�C��ix0�9O�=I*�H�^�\E]]�;殰v1�э���/(�u��F��=�꫃P�Ī`ȑ�G�]���i&v�y�(�L1���2�?mW�lH3`,����=�2�z+4�����tJp[$��:G7�]�]١���#�֮�ɹ�
��X����g�Z|+J{G��q���i�|�6P�(�>�X�5ܽ��xϹ0��X.�KVԳ�wʳ��ּ�|)�S&��3������"����d;s{�T��W%>ǖ�v��0xe�8}�2%�	s�����t_���f�bgϥ&wQ���3�eg/K�̹K��t�[}�ư�Ǚ����fQ[0��GG+�ʾIm:�U7���N?k׿`���L��z0s˛|�j�#ŝ2�i����%2���>6�no�]�[�j��p��:���{�u��>�����ǇCu*U�;���R&���wW=�=��X�����8�`..�r�j�g	�v���q$����ts�EŒsU�05��������ó��X��8�k�$v;��,���C91���9꽔H���H��\"�N�����f����C�h��Is�3����ʴ��CC�m�_]Xׁ(�S.�y��n�L�>�w�#���o%^1�����f!�ъ%G���+�!��9�
$:��K�������a��qgR�C�PW�uU�BΪ�˂Cl����Q&��B:<5���Q�-��5�?p/
��g�U���va~�]�4�Nw�]�*9�+a�apsF��Gē��r�p5=R�:�����tmu~�c7��|��s�NVmL��#�e̬��A��<�-*��B�4����V���:vAh�)D��=���TvPn��j��bL���b�˄)�ģEsX
��]�-y�%�UB}�7���J�^ux>���n�3�P�2ӢpIy�X������ܕ�Y��W��v��,0~�jlmӤt�����p�q�W�8W[g��5N��S��چ{�ݕ��W�J[��S�rմ��-�ta-��ә;�3o�Z�����'R�g%ݎ�v���_W]�=�i�S������]�x��N.0�nש�]Kߙ���Y���=���?�(W��vu�;���Ѫ6+ld�<ǹ®g��IpT2�ݓ��F?�pu�C\����5��ʫ���~��o.��b���K�Y�oU��:�:0��<�0p2���:��L~�=P_�^�U�� Tl'�bV@�i;�ʚ--����)���[�,o��<�ȼ֥�b�c}��m
�>+rˀ��7it������f�{g�n(W�ZWQ�=�L�}ش�q"7����K�S�5O���W��{pW5�v���H�YR�e��K�e����H�=C�$����̭^�C�ɓ���x�Yh��*��[hXR�+��*�.�-1����(s/3��j��c�����t�N��k���z��kMC=U��(q)�ɘ��O���Mo%�˯�1��q��t���P�/���c�g�^�mӢ��2V]��vGS��%d�����n��ϒ�P8붼6Y����"�|a�Y8�dtFƦ�j<�c>+����y�9��xW8�:��m�f;���,<��wb� ���^�+@������������n�y���%XZj�f����I�Vb���N������| ����+����3X �ᣲ�����D7��H>X��X@5j�U��m�EoGV�j	��Xԗ�v��v;�=�~���9���\ru�z&-��W�f*_J$J�hQ��ݍ�A�3d�r�k�^X6*Z<�.'κ�
�>11r�zxA��>�zfq�O'�}��� Gg?<�#9��OP �2�/}K��=��r�>�/8Q������*������F����}:��P�Uǃ&��� �U���t�]~��w*�9�Z��I�GUcW�}����+;����U��p՝�>ىq����TYد��>(�o�^�d�77��.�����{�N(Ehs1��Yu�K�����S:�l����U.��z���qg�����C)3ٮ�-an�a��-K h�_��C�辦�	���Z/�=j+���GʦJLx9kaᵷ�q��y����P�����w�Tº�oz����a=Qﳕ?TZ~���R�t�㪤���v-39H��8�>+ =w(w��s���Q�V�U6t�ݴf]�VT�Ԭ28.	0p��P�����$ T�_�|<���yM�I x�֝�U�K"�I��L��-̡��h���J�ͱum,�y�f�vYX8����9���\i��x�ğ8=�U���WnbU�r��>1���:�}܏�CT6��i���3�/Z�̩��%r�|_j+7-Q����V���u�=\�3��^%�7>�xp�a�63�Yim)��JǠ�__
an�Я�x�"���~�r:�G���������'�$�}��!��°�ۥO.��2�Z=�-z�a�bEܽ�F��=]t��~�OB�1ъ̝B)���3cZƻ��d���[�A	��عr����ҠW��4��jJ�����=,�`zN�o �9��v��4;*���.@�2TG��=ͫ#	:���,��\^��i�}N\ՁL�Fg�,�y[��|�qVn͖@'�n�$���zYTH�8/��hG�`��L�C��_Zg�}M�ՁLP�ߪ!�b�Π���2�>��&�0<v�{�g�L�a��D�H���ew����F=�� }%v��ܛ��d�'X=�.�b"�△����=)x?�!o��Z\+Q
�Q�{5r3�eL�X�����9Y����je3�z����e���(���	���*i%����kf#����udT������J-YwKI[P��e��R# }�,���sƧ��|�G�	�oF�vf���
�?'��"mm>J	��w.�m��D�FT�nU��}����35�v���Yn��m����>�ح�<7+����]Q���g��VS�3��6����Huh�����N�����R����ܺ�(1m�˷(��ʷ7�vE�tz���k�˦��8���t�/oK���sīLƉ��I��I� �u����S����Y�#�L�Z�5+w�I��
��L�#ʇxKU�`6F��oh��y�^�+g1v�h�r�f��Jݺ��"�ڕ��_�?tS&��3���m:|=��Ֆ0���.M^~��9Κ\2e�ݲƞ7�L+�z�jg�ﶳ�;T�K��.s���B	�y4��x��`.�H9Y�{�i��h���?�=�,�_ ��.�fSN=��ǫ��'�'L�w�jn�mp����	85[3Q`����׫½��o���8e�����xV�)���|z��
�|�g'˟�.���.�GR%�L�Ol8����њ�^�VWn[����}q�U�e��� \h3:�E�P=��J�nl�2������׼����+��4{��\9�>Rz��T�Zj`%�;H�j�˱��#����0���w���#�yߩ@�:f�v8���~p�/&*<P��<҈�+�6C��ԃR�t�+<��W�"��>�����3�w٧�R�u~�uj�i#��{�]gET��9->��Y̽��>'x$�u��B�������Y}cl�� ���ˇu��V��PFU�ت:Y��f�Az���W�x]�,�w��_��f��w��Z38��y��"z��S��N~�X&T#��'�;���l;�4�I3,�<���b�;�x]PƵ����~�l3���^���9Y�2���}2�VO|�P#���]��P"����ȈO�r��/��Dy�dg��:τX�~1&{¡���p�e]]��K�l����(w˺ۭ��tYK� W�P���y�3�>��^�h�<�x��仭sO�b�z7}�3޳Uhϖ�;�˲P�»/���w"��r�x9��D��`�/F{,�'f�a�Ufm#��)��Dj��F�+�=k#\/�����<_��E�ϮoC���m61�kt7v��I�!h}�1��e3���(nj��0�:��`���Q�e^���۾��	��\Z���n��^���(t�"��,n9m'�Jƹ!<��/}f�ǂ���Y}����읛��[��<tdk���D���E�ǃ���7��P�%��2���R�:��%4�7q�����y��@��r�È�ZRR��=Z\����Ʀa���5��v�G��y�u��it��k��۫��շ����՝��#{T�Y����N�Xքn��%t��i��Z�#��h<��Vm��.��Y����6$��SɎb��WC��F��D�ә(mGO���r���������� t�?slu��s�7J��ք����&Y����Z����┮[i�T�[׫��J��#�{�CS;W�(@*���%).�
/W@-���rU��L
T%;
���:�7���S���:t�]A�m��s��c���|���0�ҬMmv���N�Ǽp���7�pP,mR�(��lM�[$��jvB�W^�����WKTt𡻼)Z�4b��v�-�V�x���Eي��KHԢGO���j��	�������ݎޙ���4����X4� ׶K��2�v�6̷�bBr�S:f��|`�
�oW8`�>���wmw	L:k�sa��V%��%�P]h��:c�j������m%�bc�	�^)�q�F���rj�T��Wr>�����ζ�D��v��k)���fJzEj��F��Y�\���M�C��<y��y�4���1�)a�[���軲Sq���9�,i=��Q�8/�)pvۦ�k�!�O�-�Fm��A�[%�D�*��wG72�8��%�՜�h�uGU��Ҭ��'�olֽj�B���:[�[^3\�΀9�E��#t���I_a"��M�3r�g	Z�F:��񌶳�ч��L��,���i��}��_)]"�v��P��ݴ��L�s����O	bR��E���{���|�^��f�okky���������J�>�*�fk"�o$'ut����5s�y������e-�x������l����7J���e�٫����t�4��;ti��j`��,�YjJ�4����.)M52�������%&������o���ٰ�1K�:9�~�2
9�.�Y���2�l�[���r��:U�x\��](H:��\V�s��E��ݽ�$-h*��U�,�[�ୱq�z�΀j�3B�=vcھ��-e�^��-��3Q��08�5txH���R)-x�9�Q��Z�7BouǦ,=�Dm�������yR�,h��Rjs{�]��5�Lĵ���]���"�DE$ލ.���ݸ���f�A�[��}��]0��Y�!�F}be�2�o˺�<;)����E�ܲ�w�҄j�F�wr��ض��fӬk�:��d�9m&{� �\�c�s�;���L�s��8�B�����]���] kc�ڂ�4Mi<۸��=��Ƶ �E�)r�b���8�	.���T#�;��N�N�f+�����Q:�dTũ���u�����.t4��4ѣ�v^R����O��Z(a}ɞ+���d�]�Zʭ6D�{K&����%Md�f+�+x!�3�;|;�� �Ɓ �,�KF���R��U��h�Dkm*�T�Z�Q(�"�c*�m�E�r�e��[�*�V��l�aU��iQZʌ�[Z�E�Q�Z1Q�V+mJ�V-�bb9B�J�T�E�b(��ʭ��E���V�*ڴF�cl+V4��F�m�hƥ&8�KPKJ�cX-�-ilZ�6L�c)e��QF؈(��ֱU�(�����-���[D�b�R�F�U*�L�"e�m�[V,PDTb1VУ���Y+TE���X��bԨ�e����Kn5Dj��TE++P���"T-�QX��֣hU@F�UDeUT��h��(8�-�E
ʴ��YZ�Ʋ�m����jV*���`�Em*���ҥ��
%���(6�m��UV�YR���[���B���XQ�����E�iE��iR�h�b�fQe����m�Qm�U��0R��UUkm�R��62�B�ڈ�([Q�*Jԍ��UU��U�&5`�����2*�Z�-��h"�Ղ*���*b[��xVS�C����TBw��a�٣t�������93���I(�F_f 6s{}NeG����o\��w�vE�\���k�ۥl��'�����B�K��g
e���3���Z!!U��q�uO]�B�L�V'g;t���J24:��xzU%���R�gVT���e��r~���(�=dk�[-5>��Y��(|r�����}=�4O�C8�����������>A�{���:F/V2�55`�FRdT!�I��B���ҭ�]tX��8��<�!Iv�9��#��]H��m��<Nm钸���x��γ+��2�@�c�S�ݷ�=�	D[�۾��#B�(:;ԩp��Z�VDǺ�f��xt�OL�9�qSW�G��nz	9wW���6|�B�j%t��A3�>�R��[��X�1,;�O��j�r��<�L�[U�mq[G�̲Y�l���qV)8��v,�U"����kP�4h=\�����/�7�
��O	Y��%�X#@�;�v+�S+S4��壶#^}�b-��ɼ���邪��E���r˭D�S��ת`d�9f.%�Z�i����2h�Cb���#+:k�^U����6�^J��ֶ���ӡf�.��+�g���o���@���EtP�|��^�v�[E�?��������J�K�E֛em��w'>Uϩ���A�E�j���V����=C:e�R�����^���&x�צ��f��6�,让>�@H�}%㭪��,�j���䫥mۥ��+ϯ9Z�þ���uT���Ӗ�g�m�E֪�����I&'����݂��1����?mu��e4p��`LY�{�¥���X`�b�2��t��z�;3E�'W?P|��U��63ճb&`LtJ�a�[��2/�S><v)�b�˕^��9��<����O@��<Y~��#n^�
ëИ�3藆=F����3���AK�vK�oK0���p�)�d=Rߩ�*��!�^�v�*yw�ڕ�Z{�����&H��r��K�J�P���&3X<��FN�0���5����;C�>�u��m��-�ڬʗ-Ϯ���(�x�%Q�(O/DL���m����ƻ��Нh����q�W<j��訏bL%�DW���g�S�5`S.�6Y6򷕜�V����{<��x�A,֣|١Hh��K��(s���L��b�\:�Q�n��w�Ni��F�Fհ���d!d�Vu��-��d�};S;Ԟ�9��9��]��q�B-�j�mY}Qc��].Ɨd*�ړ�/8��utd��Z���'G���	3#��a�e�w�N�/��n+R���pa�����F��H��g{�Y�ȘP�l���&�_*�ެ�\���V�}K�	I�������2��c�2�=�L�B����to��.��Z����J��^^��5@V,��{g�N��J����(�`ߜ�9xL��IakٳFu���9�.�^-X):���o��[�8�7|�V�0�*�:$�FrR�ixa�rE�¢�;rw�j���*��Y얚�낧�\0n�C��߳� .�q�J�:�o�vp�K�j�n�D�>̤saͩ+ΥcC�}����´��x'��P�Zh��W'Uw]�۾��L1��C�f�B%����dR�n�%m�x:Ҷg�i�)�]o�c0e�C��<Ws1�;v��@��ϥ@t����=<������p�%�d��a1�"
�j��c�I%�����̀�r��3�/;���R&��Ip�+yZw����-r-o���`Y�ػ�Čϩb�^DM��;�	>�� E�xچ���.�bͮ��'�w� ������ne�[�.��	7�1���r^����ra�Zn�oˤ}��؇1�҉���:��1!����g[Xt�4�{Q�\`H��<��o"Y����b/_e�{�/�9���%9\l7���q)҄X�"��������:-���
ti�s�����0z��Y��òX~��N$}�T�{%�,:��05Q�q��Ԗ+��G:YoO��b�o���Z���:��J�ʨɖ���<L�q��w�G�W�V��$�xዝ�Y��Q�OR=r�6���!��p��n�?d��T���S��K���/Ǐd焲�s�g&^���e�<l	f��G\a��\�wW�����~���|�ޛ����3T;a��/�N~�Y2��v:����.��QΏ��n������o���W'Q�uJH���<�;�Zʞ�,��	�A.eL�y�}�;�B�42)�sد6��v�UT�bД<��Qhg*;+>-�u�E��I�0˯�խ�N�M��Ǜ���ܼDP��UT/aZK��G�o�]�5���fk#���ΰs$����^ɥ[s
�h��k��:��"b 8_z���՟%%���J����}9@f[���o�ԝ��Х>����Ֆ�=K�t�p G	�C]�z,Ƹ^W^�w�w��˾=�i eFۼ���#e/�gX��=|�VK��X�y�����L��67�b���̢��C��ПSk����#
�Ǩk���|�,jvq���"�!� ��0���;o�.�.�q��xorn%����
����ءC�o�v�@��U��i��e����׭�춗����7�U��B����2��=Ќ�c� �9������{��:����0�!h��L�~E��U����E���[I�k��f-;{P�n뻯j�g��&N7�f:Cb��uu��{=p��n�+񒎫�8��j3C�E�W���Q�t�����:y�O1�^�2��/L�tSuG�Y_7��P�g�Y����S0�����>��|7}N�s��8��ܜ��~T|S�jV]j�����z"���l�=��96�>�z{���s{v���ʅԱ���v1E���dhg��K��U��Z�n	��b}[��z����)��\������'/�'��*���i4l�E��ӳ�6��5�}|��Yxn�#%��,䩵�e,��*�0���B�#cSJ��8���tƖ��8 4��P<bwe�h?Pϩ�soL��d�+�ys�exZ��S�p�v���q��FA�P8eV��]l�ų�uQ���[��Y<]�{�mX}�a*v�g�0��.��p�4"P�<�y\��R�{/UG�bݳ�ڝ�C�'�nl+��
���X鮝B�0�C|���&�ыw�s��ڴ�&��Ɔ�N���i���r;ݡ��Lkt�3�����S���7��j���m�̂dZ��(W�r�B���2��:h�ܩ�)C�]4=�Ic^���b��7+}�ǉ�y�F����5�˗ˢY߁�H>�,n�kv� �xOQ����1����3bGV���FܯDv�g�GF},C�bF���Ge/��دP����-��ϟqGu��6�<�7ú`����-|�c>r˭�'J��/()b�6Ov�=�~�W�g��C�3��Xf�ۨ^�WT�@��A�"�X��qc�����dծ��e���a�V�/3ʥ���Y�z����4������O��o�=�2d�4�&����Ǫ���"xJ��#�8�V�㴤]���w�Lψ�Z���&�s3��10��=��?P�Z���6!�f�JJ�d��X_��
T���
��E;�G������ӵ�L����-8�/W�K�n\�8|&ÜU�Um��:�y��٢�h5M�w�J�'�,0rQ�u��r�jfC�螛��랕�Y)@��%�")�C�U׾�����h!���.6Bv
�չ6��kl�*SKRl�,� �L��R�w[�籇�eJ�h�^˴r㡒FYs��v�P;n�r�\��C��j%��#�]A�1�u�Ns���8�k�����=�8��Wv}�����#6{;P�m� ���&Ǻ�l�tbu�Ų3cZ�����la/#����}�`��j|/m����
$^}mITpl'���I�ex	c�a��N6��^Π���,���;ؠ�¢4�\���h��/�L带תyB=��L-a��ݵbe!��͠�� E��ꋸ�+������ҠE��0I�S�Ŏhb���j���z<	�⺤��ɝ�gby|s�v4�s̳�d���&[>�d�`O'�D�����R����}�yj���;��J��ܞ��'���K� �B�8���OC���P؞4�t��X�SE�d��ԛ"�>�����u�A������YU�創���8������Bz�sqbX�}�H�/S�E]S4v�E:Qj�����0d�#�gpv��/ǜ��_�����=�$��
b�R���tiu�c�9�nX�}�v.y���M����E�&�+I7�JG,�=١
�A���L�>�=��3��
�o��g��MQ\쬭�����<�z�n�05�R��b��DK �Ks[�v�$a����{�,;��-��h��]I��v��=�$�yn�g>�ݴ۲�Hӟ_u��-L]Q�r��S#�bq�:��iT뺳���N*Fi�c{-9V�uH���JA3��v=��y{JwB'�0v+�ȫV��`��o�^O	2Ԡtf{���)�^r���*h��xϟ�y1�C"��c���L�{�X���w�ߒ�ǎd`�s��Ig��r�S����U�L̝���ܾ"ԃ��5=ḤM/IP���o�b�0���
�`ʙ��Oru�i�K���W¤G�c�0�����?|y�E�	�[՛�,B<��s����m�kԼ�#H��R�O�/��S��8��:�,�jm����oKH{+pg��/;u��oV}2��������e:�uce���2Ҽb��(��wڳ^�ۓ�{�Ga�:���Ô�v׃�q�2��Q�i�
�����t�Hu��99�w�J�b���7-�O��^�7�\�ᕼ��]9�H�88>�*v���̠�uj�&+��J�Duۙ</���uT�����h^Y룧��#��u��NuR�$��'�����.���ԁ�+J��k�S�u�.�YqZ��[g��ؽm^�GptU&ǋ~�+���2uZ��� @�`ض���3�O����ܢuͽGz��4��^b�h1;��0!32����Bv8��jJė(FQ+��̝u�lU�:WqĘ���^"��C��,�V���8v�ЈTx�W%�QS��b��}����ɞ���J��P�𻇬gXE��Ge�:b,P�g���UW��Cuө�3�GE�Ň)x��"�����I�Y�i-r�旆�^��\.�P�n��^��Y�8x�;��p��Vv|r��>=G�CĈ��(N�]��tOջ�
�\�^�{,�s|�9�.V��dt��
X�5G�����.�E�ń8="�z�F�^,�,�r��o
����,�}~�B�s��S��ڮ}��� fS;X#�:P�����%q������&]V�ˊ���r^������=V��]t�e'K�Z^%c\�1i�k�����E��f�S��k�J?Ki���z}q�p�|D�w�_C���̺N�o��)�"��{F�u���s���	���3q�L0�/
\E�L�U�܋����[t�;7ٯ5+�
����X�3u��ք�%��sj^�|Xzj�𥶁hr��h�g}<A��ļ�gUsԘ���!_4�T.��<&��^\]+���PĲ��R��!�Y]������ɓU�Q~�����os�w�XTK4��U�k�ڐ�-Z6
��D/��x�M��Yf���Ɍ�B=�.�4H�j�(d�vI6;�]G��'d��W'Ba՝|�h�;aS�:��.�wj#��c1h���ҥ�{����{c�ա�?2���d��^<L7�S�>�:�l{�L�x�7�V�:2%�f��X�2<��L7�yUUx��]��l��9*m{e�K#슄<�9�D�������&�յ�'H��K�@�L�we��g��9��J㓚º��gB����i6�(���t�,���H�T����`��e��3/�Җ���m��Og-o[��ԡ��J<zP��ѫv�7ݙ�=��yA�A5��].k�(S=~딡��%�@��*�T,כ���y:��{��<"���E���eI���4��r�`	�%/�t��^�=��#�Ne�&I��^J�$��5gå�u	�sT8V�$��a�yc<�}����������,���~Ԟ4 �]c����Z1�N�1(m���b��c�2�G�����%��1Z~�~]簽��u�w�R\�bK��eޔ�~}\{�-n��;��X�2������K�I��-����8��U`����n|��-�nh����u���ۿq��p�[y	�]��V�����
Bi=z�����SЪE`�L�q���fa�xq�O����k��۷p=��niCs,a��վ;z��}f�Y��Σ���r�o��|Ť����ஷ�̡�m��v���.R��O1b��,�[��^��d���a�暀��ls�4�,�T��I��imE������:
Q����Z�lgN�u�ԅ��_\@���]á<mVtds>��a�Z1=pp�Ӆ>�X+۔\6OjWsa�u��d��7k%-�_.�^�����{^���fq5xYQb��

��6��Gf�ʌ��F���H²=��(g.�� \u��]���&�sOR|~��:�������ŕ�k�m]��������F2�I�4����6!Θ���*$����xx��Q��x(}--�I�d��Z�.�s�C��.݉v��c����$Sx�;@��q�Y�h�s���k4Q$�=iT��H���K2�<@�[�B��u��K3�O�=���iF��WX����7�Y� �:@�J6�npS�;�V��&f1/opQ [w�Z�eyi�aP�wV���X��VQ�����Q^vˉ�Kr�rK�:���!�mm�'��-��׌��������O(܁̙��Oٻ7��yz)sF�4��4��N�
�6d���kVh8ɥNZ��2;K��l_h�`W=ہ��v��vnu�`:��|!̮{��ѻq72	{�2ޣB�Y�'�e-�T�XZ��t�;��K�2�.뉢�ϫ�K��2�f�� x�d���ҹ7���Y�;xcy:��ޜe��W�e]ȬdgZ����Y�gK{�Q'�*�r�w�R�E�gA:��Vg@�XYj�@�D�.k���pQ�@�ج������]��g+��mv���h�9G.��)_W�c���ʼ͉-� �0-)��sT��|�`��kѽ��t�r+k���.��&ի��X"�x��|�=�����$�V�$�@�?�����m�����8�oljFȂ}vw��A0�&vnS�-�5�˴� tQ+���R�v\��)]n΅ԛ;�mh����:]��w�>���G9�n�go���gW
�+;��w���D�s�o���뱏ni�][b���u�t`�qg����oil�G�����,�U�$��Is��{�oKz)f)�y�_kT-ݼ �*I�����3��sM�p�[N(�to`=6mm�f;����4���Y����z7�m��l�X���kd��gu�@���ͻR�^���s/�}қ���#��j�!IIÎV�s���z��t��EV/��}ǢVz�3�Z�e:�s%�y��%u�\�@�Io<������޸ W>&��Й��+n���O*���AP��GC��fK_M�)������j2��.N����l�Q�l���E�
�f5�P�S-(�j"#TU
�QU-�+Z��kkcmj
V�*T�-nZ9J
�(��XPB�|˂V�Z���k-��VT/�Lij�YQE
���h��%�ڒ���Um�T���+[m������
52��m�Z�IJ�̨�l��m-�B�Q��D��L�F2�ة�r����"�
��̴��hբŋ*V��bQQ¶�[h-B���Z�խ+h,���X���"��UR�-��ڹK�XŪ�+Q��0U*U��U��J�"�m
-�[P�Z$E�Z�<j�R�XڪXѴm|f.DA�Ֆ�� �4�j(�DKJ�Zڋ�-�ҥh�[l�V��b���R��V�j,Ko��V�TE��jU���Kh��Q"�ţm��h��Jؕ���j+h6��bګE�r��D�KQ�ҔEDU�P�ҋj�1��[E�j��ՊZZ�UZ)j)mV�V6�Z"�S��(�j�̘�U-���QE�Z�Җ�j5�+cm�jA~�B����Ck:�a��S2��G+]�2��dw.9{vkX�_G���Es��e��|�����s9�ej��)x�Ĭ�녹:�]�~��:݅��H3kŭO�0N{j^�F�o*J���S�=w��y�$����7sà�vj��"���l/�{�PÇN�m�~��q�1C���/��s�y��ab�>:c�3q30��ӍB�d��r����Xlg���Vڗ��w�UY��ۻ�:E��*��a1C�]FT�-�� �����L*j*��P85	:1�^9P�N���Üqd��|�L��\�h_
���Q-����aϋ��v����̼;�R[Wǐ7w����h3�'	�1jc�+C��Eඤ�9�X���LC$�2�ߗ�����Sy���d�ˤ`�7:�<6:���I��)�U��t�߅9sQ��FS"�7��/R�����d���z�ɑ��Pv�OR:�#ǈ`�K��YS�L~�;FM̔fN&d��w��G}\s�RƑa�y�pL��{>�l�O"a_L6M�$�_�����S{V��]��@7M>�qN熼R��1�'�������¡�R8t�QVE0hV�ޠ<��!�^/m�5w�\k�z��;�TAu����1�}x����w=��ڐ�g��9��;^ǚ�<����7�����:X��]��^���Lv�[�9�f��-\q0Ф{Wv�3#����ۃ[�gS��S��͝�خ>f�.���W�*��h��]&:�=+̘�c�eW�H���&xu�sI��Ѱ�s$�<��i�{.���GY�/-��pUC�^��0M�:�N���0{�������yw����.�H�C�m�g�U��d���m�Z��y7\.��P�>�7��z�ݥ�f�%?nEw����G�#�6t�o��B�V4<w�I��´��x>���k�lE���'	�}��;�J{L3~G�E��(��yb}�r�����]���U��y�k�qbN��<8��Wy1�}cb�P8�4�&[=�"x�:�¾����˶U���M�����P]�uHd�W�c���� ���]m!�*JuY%û\1����K�lzz���H��ӻ"�1D@�[�J��*���ɾ%��Nj�f5	�/S��J�EK��<��7��|}U7:Vڶl�Z)qh�>��AuPT��x�}JD��.U�ջ����(�v-��2yp����c7�X&\=�^*���a�u&�2����ɖ��b���y��W��ˑ�WSy�ʸ���*�M
,�{,;]3
pAj�-a���t o��fg:�$.�]��t):��	���/�>��u~+���Bدw��`��9oS�N�Bάjk�c�yS����G�sg�	J��%Y8V�w���𾰺���Z�o����c�{ 焵�0�	�����ׄ�#�.��`-5�����KsƵ��.N�W��nxnܕ'׽���f�f
9೟L��_�6��1Q�6O:�D��Ʀ�ǽ����<�b���GN�C�XR�w\��bt�s��};N���z���55\�:����bΦ/�/��~�sj�+�dX\l5\zm�����U��9Y���A�C����+�Ǜ��eA��*�]T����	C�{���ʎ��[��X�m^mn��R�7��%�t�yG����C��뤐�Y��_[�1`J^��ϟYyk/V$W��nS��W�Ӗ���\��{G*uK�!A�6"����}t��]�Az�~�+`��,��e�wn����<�:���`�෵Y��R(p���CֱFl��Pf~�rbs�V��8�h��'	���m@:z������2���Qҷ5CNʿ-��:8��{u���mCC%�#�e;�c��P�H��X�c�i{앍r\~��]b{�r���_nf��[��pwI�׮e�>jw��患��p����t��:���[�^>��>o�f�o��=����a*٫�f�V�U�!��D��vv���`�p�	/��,�`�Y���:�w")_�:|ԩ�]o��6��ș��
�H��e�F�|~�����?����k�K�L�#m��_�j�}yg�ڎ�튓��=^X�5^3q��|`�[�I���E�{�Y`���J������Ƽzr�þm�=%��Sm���G�|���Km	���E_����mN,[�0oe�j�JuB�X��Z��v�t���=�|Ֆ�ő��\�u�b^�_+�"^��\.�;2�z"a��uC���Bq���	���7ǵ#���@�~�No�>�$�L
�WɳX9*m{e�Hd}�P��)��o/o}y+k�2_3׻s#9�A�ԅK��|q��X�b�/>����9��J�Ny��9%��E.�T�#���yO��j�$J�����W[.�34e����di�~Xw�,Y��]F9�=���t&�rL6�r�2ʡ<�V;�P�nU!uλ�g�r�P��4&�і�U�ޜ<�Ko�'������.�V�	P���(w&"Y�d��.)XUCS%R2�+�鵱+U���5S9��7��a�l���:CU�_Q��pl�l�K���j!F��#.Zݻ����13s3�M5ao!��1�$��t����q���yL]u�2�j}����,�a�qm��sC�X��^68���ھ��޺��g�S��WI�F�r�b]�WHm,C��1#?��6��^���[��p���G�R�.�3k�r2�t�UH9p�q&��Z3��'I�G�Z��-N�}o�uv�p�L;�@T���{����K����7���@���A���z��n�4
�lq�6�=9���;�f�`C�e�b��;����g�V޹�^����y>���z�*�=&���H��zk���gg*���OX綥��6�[��`�3�i	2y�3��a���ά��w�*�n��׭`�ڕ��K�m�8�,x�i�>�G�"IPDA��8�z������*������(F�(�|f��=��l.f]��^�a�Vo;IK/�`�.��R{J�A�C�^��'R�һ�ȡמ����S��FZz܉W��<�zk�R7fK�]�Zn$�R��|*o�D�W�:1Y��L ���*����T;$���M9��yCm	u@�Ĥ^��-���.�N�H�O)�J&h���`ჷ��x��G�X�&`@˓�G��rd�)�nzR�(}�r��}�6ۻzz��c�k|:���n��Н�ٙ�hR��.�۝�w	�4��7�(7fmu���T�F���Y�ȣ�7�w�e�Z����#]�r�u��⤩:�������]� ���T���ޗ������%�0m-�"��N�>��Ng�:s��2f�م��ޢ`<�����=���)�GPiP"�� oZ�[�t�D4xJ�N�{��u�L��z�L�u�RƐ�?z�L��{'�9�O"aS�s�$���+}{�����3�2�N\����Y�_Vun��0k2�P|e���.enxd�p��p罄���/y�.۝3�^>F�X���K�����+8�|�Y�u�zUE|e���4�7N�������t������,-0?RK�E�eJ�)&F��SeVXf^ڄӕH���n`���)݃3i���K���Ԓc>�>�ז�����qK�·���H�k�ӞU2�ֻ��7ʞ�w�G�h���l��wG��3������1EI�Z|>��쿊�DfLRm�/�h��k|�����\��q�|"�z�t�ڥ�k�j+Z�ى���˭.�xy�Ĩ��j�Ag�0C�/���cҺTM���ɖ�v���<lr�
3��Vz���Ձ��л��%�#�a���nd�罆SV�&�ڑ�@�u�6��8���l�ԛC+���]�\��\��k�;|����4vέE�$�w�h��G���]�d���2��%vT��n��*j9I_X�1�1՛��i����s��tG�Ok*d仯_W`�~��L����r�N�=B�-�ĩ��������=�3�ǫH����d��c��+�y�nCY������%p�(��k�$����Z-{.���������B4��Og�m���.�h���#l�|��PT��x�/�{ĩ�n}4{#�l��锹�]=��f�G���7�Y2���WPU��(��j���	@x�/��gƖ��c���=����Pc�n���Ja/+qv�9A=H��v�M@I�\z.��i����^X���-�WOG�֐�q:�XY��a0�慘�ۗ���ތ��0�޿�&_k������w�|��)�6�e�����u�=�3h)��S�d$����^����;�m��=��H�rX*��z�dPƃ������kO^4���\Qe=���W��G��%l���!��#W@�;�ꐷp�wh�!E�3���~���"��V=$����0̾�M/�����EPe��b5uT%g���G���w���ޟ@�t��q)y�X�Zے�]���
!<4u��y\�'N�*]�u!�jGD�4�g-��p	��=��1���;�-�O�f��Naf�X+���."j�ü+���"D\b�����B���j޷��GCw�E��X����}����c�^;�s�_���ʶ����|0��%Q��Мygԟ-����P;��(�Io�(��i2����3��t�����6X:෵Y�j���#e�%Pz�y,�R|��7����ef��,z��җ��gN{)�+���;�N�^g��s"¹ť
�GtX9�=~	d��ox��Y�77�׈�Zu��e��C;/U@_K�Ac����U���r��m���sa��궃��q蕖���r��q�p�|D��{��z��JOi�L&�vd��	��7},Q^���c�׌�`����]n��J�E|
�0nΩ��uranۤ��U@�B��a�}hg�Q���9C޿2,>���G�G�i.�jüڲ�v�+B��<�8=�j�ҝP��qՏg(/~v�t�FF�p/g-�.u�z�<~�q�*��\�C�)��S1+���<L6���r���	Ɔw���f<�����ߕ��/��/Gݨe��u�A�ҷ��1]��_&�ag%M�}�̤2>ȨCΐ�j���֫�oD�Ю0�Ҥ(r�՛e���D��ا�ga�3����p���7�{θ�/Nc=�3yɊյ/��\ʆ<@e�w#���zx�������WgQ�	�]]����j���b����n,�Z��|���m3��T[������"r�e�s�%�PW��^�����r��f,i���0S��ޘtў}�F��ʰ�fƊ�~7ˍg�]�I%��rP]L�
̰=M)o-���*|�[��寱<��צ�25���%��}Wq�B�p^$��b���-+�<�ݶP���o�D���Zw6����gw㣓���k��ñY,�D�C]�~���yN
4"���gd]��@�zu'*uKcB�^JK���!�t`�:�$a�14�1��PKپ�q�,�*B�Ѽ�P�R�a~ѕ�t�UH.n$��(���=����D�<p<�^��p�K���l��)��pb:�?.�X�C�C�oEuI�B�~.�f5�ᢼܤz�}z�&��au�������N��Qg/�s;�u[G��e<Pp�0g��U|0�݄�� ,iw�x>��>ٮ�}�͝�e���XZBT\SB��w�܊�)Vz���ac݋L/�-Y�M��i��{ɳi[n�o�ٓ��ݫ�1O�0���7��KZ }H�:�ǵ:)���*���L�28RTj:���!8<�k�i�39K�����U�տ\w����ɭ�����Y�Y��k�<����M��'&�i�KjfqP�fj�#���pI+.֤��:u��>�خ��RGLƻ�̼
���Za.�n&f4�V�P���(Fܼ8f��3@��\�321���c�s/NAU���P�W�(X\,0Vu�R��RL�|+�{^2T:��/�i���w���w=�~�K��,&=W����\s䖏G�{K�6�l�yٔ�2u��߶����1}���߈���~Ъ�����4�aUD�?�e|�0�J���E�r$}�P��#�Z��W<�T�g��d��{g���7��Sk��U���(�'�2s���V���3ì�8�='U�;{i��ʕ�L�xlD�~[ԏ������!2��iP?q��Pc�L�]%���b�&+�cT�W[�5b�p�ߔ��[��,��o��ϰO"a��,^����.�E/k֢[f�'�>����B_�ܷT�s�^)~����>r�V�c��j�v|��^��}/9�p�3Ƒ���J�S#���l���z�6�+.d��Hx�m��+�$t"�/V{�b��k��H:~���D���R��I���Ȧ�Z�����G��%�����]e<CB�y��]{��	Vp��A�v���D�=S�a���G�*G��n������ý�12z��6�� љv��Q!��Q,�r!v�Dk�*�v{u�m�CHq[I��_\kK�T<;"�m�{.��6�_'H�}Z�խ5�nf�Dg^���/��N�o�����s}�{4c�S�8�=���yS]*v|�M�'Z�Z��EL�	r�|Y��#G���D�~������m�v��n��<�+0�{�n'"	�@Z3��v�u�[�u5٩��Bv�ǧ1�֔-�էo�BaD�r��X�w9j����8�sfU�����}��)�-��)�1�{XT��3���敕F�,?%�~io<�E[b^�6�׹�]:�o�/j;%�I�f���c;i�\��vk���)�j�0:=��6�C�Q�h%�&�+�t��5�FRڧ�����3+���w�W�2�C�V�^�W�^�Zml8|�ˡG�ӊ���~����r���5�sr���i"~�ì�t���v�߅�)�lM�3�q�M���FQ�6(ڱZov��*ќ��£��9H��rr�����ۤ%�e^����/�+���.��A�KE��w��]�k�$���|,�]X����6c�{Z�TJ�M�F�H�W��x��nB��Z!�6��wS�JaG�W�㊕	W����j{�7*���]�{wV+��Dj^c��$�論[�deEN6�޼\g���v!�UJ�o#z�^�'[E�L^.��X�����#����X�o]�{����켜��mT�A��ݯ(A��m=)�3��e���̢r�Cz(K������#G�vV��N�k��0�Vf:��H�y�*.��Y�F���T�/�v,�TZ�ꔓ2	Q�`��0h|�-��7����+l�¬��GgC��fI����ۡ�V�q���Y=T H�k:�0�{Q! �It��WNKEݞ�)�³�s�#%ޱc5������H{HD��0�_I�>�5M���m��sƏ	�t8Gt)�Au�#�:nh���z�g����\7/�k;)e"�;V*;���}P����e�rT��K;6�G�ö�7�3V�W� 銡�}VW܏S̱mmم+e���u�KO�B�����c-��+XFa�7���N�+^d�6H�g<��z��W��	v�r�$�R�ļ�$����$��w;���^v}��H� $�'+�ڃ2�*�l�B�
�et��<5v��gW�tT��S�P�)ٻ�m�!��X�v	�M�k��N޲;R��derBȩ{�g\&���5�ht��DQ�kk�ofa8�����f���/~V�632r��#C��`�L�[��K.����+��?4�t\��6�}���xw�gM*�/��bqS������k�k�n�pfy�o�����@$�A�B�Ub"��Z�Qj�T����
��y�R�`ʲ��(Uj[IiV�VѫQ����F�X ���(�Um��CYh�f\�F�Z)V�G�.+l�Ԫ�kEV*��V��I�G+R�m��r���cKR���iTkm�XŋR�il�[����y�.-e�jZQjUb�m-����eeT�(*�0XѨ6��Q�0����<�̲�e���RԬF��[�YEQP�F1m�����Db�U�,AD���
�VTJ���̪���Qr��[_)��2ڢ�"�V��|�y<S)|qƴ�U-iDDe�V2��[.Z�Ѷ6����QKmJ�mXV��[V�[)n5r�\pPWZ�YZ6�е��hZ����VZVmg��E��Te�j��X��ưC-V�k+�m*�KZ1JEQcZ����miV�m�W��Ke��r�*��DR�"[X��¢�Z�""R��ը֕�H��h�a��8��ҾGT��{�V�z�mc��j�(��S4h�9����3�9��w����}B���Qi[�ױ����Ԙc�l��p9�K�<
�����t�m�xmB|tKJ�u8���H�!�����r�b�:I7,oϧ�E��:�I�#��	�����x��i8D�t�SG�S�ͭ�C�ݛ��Л�����T�9\i|�@l�ƨ����^��YB��lmt�z8�l�}�s&!��3֡�Z`���d�Z���1�}cb�����-��-��4�Kw{}ojTKa�"y�޷~��1�#~�gj�T)�P*� ��r�53��g��y���j��sac�<<y츍��b�^�Jǡ���0�^��脝��ޞ^�r<�[���<3����!>	՟zl���^Y�E4�R�*_c���	ĉ��_^yw(}[���U&$�w%7�a��	���hN+ظL�f�]A
�a�G]5uc`.��1`X��f�V������S�[3|�&!�0�=]����.�!��
�pKJ�[���d�~�.U�I4��i�v�f�l�aC'<re�z��^L�r��/��`QY��Z��+1�gY�%�rN^@W))���!�Aoy�γmz��Z�j�KFa�#��l�u)o{��(Wz��e�9lƥB��]q��Q�#9lF֣8*�h�5{��(Z]D��kqrYk� �u|�_Uށ��[a1oz�ռn�vȘ['���lfj-���7+ǉ��b �d�8�]H;��z���z��A��9�-g�*�Y�"z�����ώs�nf��HiD���׾���x��<���)����P��þ9ut�?Q���qp�-l!.e`���o�wE�/��-bR�B�E��~Yx�����O�z���q�|bL���U���p�&8�5��k��9M�l�pi��4LPB�*n�1�(a��f^n�2�T,EM�COQ��*����4%�8Wb�z��bq���Q�~^���'�3��oÝ2=�,R�ʌ�+,x�t�4��s�,vz��ٍ��3g<�xU���w�M�R�^�gE�m@t�!k�c>3)��Ԑ��k��黚^C�x�z���*u��|&����nd3@�.ʀ�����!�9�!M�*�%�З#
��)�ug.KŦ��c��q�?Kh�쫏���%\x=�3�ҁ\���޼�9M�;���= �.�i{�z�^3q��0���	u��)�x绦i{ig�6S�������� �\�����ǩ�ں���_y��eE[�D�Ș����ˆ�.ƋV��b�EG�6��N#Z����������j{'�0��&d��Ŋ��oV�9���v���������	L=�A�n5��t�N�Nô�6��
��#�W���OŌG��n�>�L�jf����Q���p�x��C��	�Fr�����P�~�o#��-i`�W	\}�*���fX�r�+��X���cZ;Tdh��5u�n{,R�s��-=�'�Yk�J�!0�rf%�F&��`NP�'/�'Ȟ���*$�VlQ�3�jy�Z�x�i4l�E�U\g���:뭲�7��e�����Bü��C���K�#�Ԯn��vhk�Z�u"ł���,��H��~��S��޶=k__�*��R�f����-�̦aj�҉��P66������ųn�h!�	b����Wu�Wz3�N�{�w-K�4�Y��d���&[�xCY�����Od}R5�qײI�t9�n^��U4�%�x����yiτPޣ����eI��K�5�&{ϵ���z��s��NW���Y��-{�t�\WbUv(ʣ�	BC^���ž5^�U�$����U�0fD2:�0���7��X_��efwLT�\"ә��HN𗔮�jnZ�>�cebu%W����D��媲�u�*�u�lqp/w ��KW�"�Y���ga�V;gٴ,����8-JU��=��������gM�+.黇8�Ot�<�8hQ����⣐�zja�)��sqQ�Iս��W�ד۷{P��>�FϦ�*817��%�K��~�#P�>�e��vWQ���e:���}[�0���J�FϦ�/:<�YC�V��C�x�;�۫�i4�{Od��	cO/�L&��P�����w�X;9W��hBx,	�~�mKa����6�W�;����Q�?�/\������0]�"���i����0�N�7y�ǖ|p�k��I<9vɊ�ߩ@/P���apJ���Pf�f`)����/k�\#�E��Ib���
6:B�f��t�!p3Ԗ3��\0�=J��U��Jϭ��;�C�WD���*�O.\�T��=�����(lx�E_�[��Ғe����¡%u٦<���OB�ٷ%g��!<�z��]��5����;WU�+/��W��Q"�[R$_�^�z%WV�y�v�������;zP�^>MNR����O$��[82_1DnΤ�[�cu�<F�K�9sV2��,����������(;V'���B��;���1v�2Z�?n`�b�+��;�0�5#�'j��b=��=է�=���:CX]�mi�j��K���|��
w-��E���E�t1.Ns�*��T~�V�Wva[�1W����T�l��ӳ���;n���T�5�t�S��X�3�k"��c/�-��l��/ʕn���ܽgO�ì�!���d�O՞�L�	�L2�{��h�f�n��{���+�DϷ��6���
+����Nxk���x�x��<�˛ҵjm����k���uo{7¸�)�4�U2:����~���^T��5�>5���ʵOr*U���:9����N^����~\��-�F�zTވ��%YX���&y훍gLN�S�Zx���`�IH�Ĕ�X~�ò�L���b�q��v�u5����Y�^�{z�2�כ~0�yY��Z�J���Nd��K'ˎmx�Z�2���">�:�__(��zv�=P��+�=����G��	czo�����"�z��v����ܮ���;�q<��7�K�S�K^?->�E2k�|�B:��/	^�w�.��y[=�A�B��~+z��S7�5p��	����ᄿ����o�7"�P{nË�������E3�kt<�nl�P>wǹo��ńaÊ���-h�J��d���\a'�3Q��oq�N��Ts��{3x����Ǣ���wE6���}�[�Fs#ѱ ����ww�+1��T���c�-�[v�2|�:ދ����#����{��V�����o$�C�'�]�rN��.�]M�V&�n�����Ws���\��roU�����)�q	Հzl�����+#���R�QJ���ZV�,k�2k��߭n��Ō�H�ܔ�p��`��~���~�ɖ��/u�i�ʺ�:R�_u��{|}�qé�b�R�����(ZXg�&X�����V���L�<�J�G÷K�~)#]okM��q$tT�-w�a��f;%�2s�g>/{������mSH��ݔ���}���h��K���� �`.��O=E�4�?�NBǧ?e��G�=�_��Yꝏ���!���I]�p�����J�.َ�X�E�6\��C�֠�0�]�{8�"k����a�k��k���PG˙X'����9�;#�k��8߆��]��R���vC��6h�ڀ���(_��$�xKV��.��b'����]UN��]�m��f+�gIb�{���y�1]k�/�o��<�~U�L�<D�A*���(L��Uyw�a	���z�vj��������~������3>ޘ.��ug��z��C����y��*Ԣ�n�]+���c�R�nھЍ-����gy#�����:�X����B���G�ODn+G5�K��I$�h��y;��{��8_�r�}�EL����t�ř����N{f:��θ륩�jhyb]�Us�Bm^/P���5���e�/}zt!���y��Th��D5��Cm4xK3틃���ӳ��N{j zz��w��Д��n\]r����!�G��-�ג�8F�^CP�֏e��ۙ�Uc�qÁ��˩�M�N�Tc�� ��� �Y{�-c�\h|V��b�w�Hw�-&J�*�v���U��w�i��o0�Q���#|�3C'5�}^��g����u��VT��R~��mQK���I�T�n�F��<�[3���c��A�H��R����Q3wR��P�5���Q�ʣ�B ��$#����p�]f��ws��8�j��l��z�5���`�y��h����=ꭵC�Ϫ
}LįR��	�S���y���2HT������(w�{�¬�'R��+��ª��WdrɳY�g%M�l�*m[���{������V�T�u��Pd "654�i
�� �+,S1�"���y��y�;�oV��~��\�6���� ��Y�]�I�@�ڹ(
���,[2�Wh���K��}t�hn�]Yi�?�=�T=|�U�ېR�P�rt�o+��|��ı�EX+@:(u�;8W9��Y���`��y�����0|�_I	}z��Ϛ�)�Wc*[��cN�Vv��\���B�\f�g.5R�{\#��c3�O���;\4-3�[o71`����˥��'ý�^�fq�O'���!���V�r�b�P����\���~�����cR�Iv�>�~3<x:��zT+h�Ɉ�{^�Qj��:��[���׉"�^*��u5����)��]f������2���Y�v�u7���	�FBQ��p�[�bz�c�l"𭅣�<ԫL��W�������JÕ���*fh�٬&�\��$F�@��=Z2DN�_z7�:ѳ�Z��+�o���y,v��P�B
�X�^zd�N=�IM�-6�	/mW�Y�[�C��^��u��4�<�\�� �&�g�8������b-<�iy����b���m5	#k�w�������Tք'���5��B�"���ϫ�g�e3�`ö�-�U�6�<�3~G�2���Ҵ��{�4���V�FS��l�v�V�]�2�K�_˂L<vT���ҙZq�^���C�-��q�T��{�q��k=v�W�1Ғ�zR^L���a�������r�S2j�������Zq���l�S���7~""3s���w K����v:��=Fi�}�N��o#�o����>]�A��1�\kU-��\�hCL�(Ҩ�yX�@J��y�u������R��4��c�,��DzK�&/pws�Oj��r�`�Ã���l�w[S��3��Fd�ܖ�|�����{G����bF�%�^{�+�X�P�B{��]�3cZ񶃺�uPK�z���W�.�9�n:[���N��o�Չ5����L�I�+҆����MN^ƇF�y&��(�6��ұq{~�rO+�{N@��q�.z�˄db&�O/yYǑ���OR;aݠC�^�)3�#c7���[d�	;��b�ŋ�2����T9���'�s̳�%�^��m�.E���0[��w���|`�'ґ'�/�
/qA�^度}Nxk���~X^�dw�;���p��ګ2}��p���8:]:�.�t�go�l^:�+�8�����6Q������'z��=v0�wJ�3��X&�H�+��#��墓K����k����?p>me=��k�g�7��V�0�|e��IH�D����?vZI��+����ʠ�k�Pd}�c�e�f���[:g'�*��5��3%��'zQ9c�9��QhB�}���{�f��l5�V}>u��ڔ=�]��]oג�rz��םί(F��jYA)SJ�C�L#��%8���om�ʙ�V�]S[\�7�rGl� �1����{���K���K��V-���s�Qw�,<3�''\��t�x�j�vR��n���r�Y�V1����R���ίg��r�ԋ7վP���}p61��a��-��u!��]�D5�k��m1Nƙ�r��LL]���7¡L��L�#�3������_y�9$���qz�vo)��9����cO奛̥�%ڭ&q.zT6<�>�T�K�S̮���|(��FĦ1��y�p:���%�ܷ�o�`XF�]8��C,�9��{K�"ۮ�+������w]�x�9\/��q=�J�Og�mҶl���������m9`�k�/�S'c\\�Ԋj�m���%_�8��B)���r���}8�j���U��,,4�ur��zo`�i���n�Pݫ�V3�&+�]RbᛱȆ�pS��^��Y2����,����t}�^���^��Cz
ZD_UΗ�$;)oN&V8{/= ��t��,�H�L��o+���_4dӞ=��7P�#d�J"y8��u��V|�cOVi����7�.�3;,�`^{H.�g�Yk���{��Z44p���2�L<������ΐ�$��BH@���$ I?�BH@�RB����$����$�bB����$��H@��	!I��B���$�!$ I/��IO�	!I��$�	'�!$ I?�	!I�B����$����$�H@��
�2���|�����������>�����&�@�� ј 	�N�VI٤�&�u'lH�h �����&`Ab�]��0     ��L� �LL&4��)��R�G�` ɀ �`20110�L�L���J�)�b` �	� �  f�4`� �� CM  $ M#"14i�5=B~��0i5)=����(�Pu?84 \A�Q_���J��T
K�`���?��W�?��d?��
F@��D�@6ڐ�%� \`$�� �PN�V]U������v�t Pt�.��
m����IL��j=y�=�������d��1�g׫��)�0�쁆�df��L��2Ԝk)���7�!^2U������97�F9	̣�9p� �Qbi㘺���8ba�]�FL�T]�Jg���O&2B�ڋ$���1�WP#%77i`T�PүBff'*Ѣ��s�b��E�S,A����(+�C(�11��U��0U�S2܂jC*J˩�'Ix��[s�U���&����)�1"]�@��J�DX�3.c3I�5�Q���`�*�ܑ##�*&	�n�T��-���NI�V�(TK�H�wF	(FH��Y�f����˱&�#<��±W�GD������W�w�B�̪t�*�9$�D����&+��9 �bȤƤ,�΁��N�ty{�O�Bj<��.�OE�,њ@��DGO+[}�"T��U�|�����s3p�����,�y��ػ��=gV��қz�m���[MMXM6�Yi��4��a°�m�Jm��I�������mɍ�*�<¨��f�=y1{uL)MȻv0D�s"K�ցM��m��M��m6�m��m��m��m��m��m��m��m��m�ۻ{����la,X	<�!������U�1w���j��U[8qCE�����zt3m`�u"
ۍ��t�C kƲ4�wA�۝�DmĖ��G%�icW�R��d@�90&����պ��xq(z������2����i�wl������FY(�Rպ�Kǅ��n*�nضl��5X2�e�1S�Gd16Ԅ��
jd)3vHV�6o^�sZ��W���?cy��{��eǉ�>H
�8$1{m�W�Z�Tz��n.����:�^|~DJ��P���Q�j��Ç	+I�n[Tr,�0��M���7B1
%���dm0@����Ǉ�#��Q�AcS �li��V� v��(@+[�l�D@T�,�򙘊�j�
����O]i������rE�'b��	�,����"��D�P���Te*�kbt�f�CA1R� F�wX�o6�V*p�qJӟ�3U����F�N5Y�f�)f&16c@I�0��r��6CB�����ZC�d+_�A����@$'�B2�0RbB�1�!����CgZ�)�q�H��Il&�I�pD+Rp�$�2!N�4�� )�t^����4��IS�%�ySIl�ŷ*�H��$5��4��!���D<��}�����q��l�i�ښ{�:�xͫ�(kDp�4�7'��L�q�q"�]�m'ַ���tn.�^Km�*[}3Ӄ2���D��7<�ؔ<������r���~�I��n0���u����Ob��ѱ��΂��)���������vI��̬'���ssƻY�gkm���ί/�  �5}֟\gY���|&��q@��:@�t��.��E�;�u�e��D��\�B���d�R������g�6Բ� ֯��5�Z�� p�CH�A�i���� b��	���� L��H�j)hF���em�X���Hm 3ʍ�c[�CH�mB��֨������Sh���`k����?a��"% 4�$|	� ֝���j��	�Љ�6�!PRB�t��DYZ����z�h��q}�ն+��8$�Nw9@�!`gyZ�U ���#5��v	-ˡ��[�ܲ�x�e@��>�#����88����'`]TW\�d��Vٍ[kATq6���}a�Q�J9��ؾ�b|���v�w{ﭴ�2�m��6�S��݇yV�$F�� Y;��k���+�\F��6I$�b�7W�g�L��E��F���w��N��<&/��9��k��P���|I�z������u����=O�=3yV�8]G	S�A���ѪK���a�1�K�Hzk2�Oa۽��o��S�r�
DϽ�K��v�҅q�v��C�y&ƣ�=�0�>�(\tq�(|v���aJ�3�GĒ���؉����xQ��-���Tb}Jl^��n/�-�`e�O�nL�N�͜�X�.&B�x�	�}�}��cړUљ�����œ��OGo�{�G�y>�����oɏf,9}��8)�b;�f=9c��W�1y�)�%U�#��S1���vv����JvK�8x��3}���m1�4�z5��ji�x�=���M��T�������#þ
��"f*b���$�e)Jo�⥷�yő}��V�r
��T�A5���@Z�Jk Q�*��GMxmFp�4��-1Kχ��W�:�\��+�a[}˂�'��Wg���jj;�fN{��6�z)Ι�s�A~O���>ʟg�ϣ�C:U���b��Jk���X���0GFM�g;�@m5�p+c�<�R)�sѧ�cGY�&�N\M<]���D0�su(Ou�@��P�Qr��u��tН{eF�OOcł9�³��_'-+
��B4�M�3���q؜e��zP�2C$橍{ή\��P�s?1j��K1xo���~�켲xp����U���.v-ԉ�(^`��J����۫���F��s�#ϓm�����m��^k�'yw���۷O3]�{E8ޏ�j܄hB9+�sLWZ,��Ao��}�l���v2QlV-6��q[�w:u�}��^ݷ�1xy�l�$�7D@�{�WD���9�`+d��c�FM�d�ԁ0o:��-�Z�DҠc2y�+{+8[��o�l���Ul�C�u�����p�e�^tF��`�F�J���eU�O������Ϋ�Ls��c [W�T#�~uRx�p�;P�O�47oF�cޜ�xE��v���f����Z�Ox�ZL^P�ݗc�t]l���ql�wo�&�#+�6�γ'��O]�j���u�eo�&b��Ay~�E� ��Jn��fR��3f8��])��Oa���W�w>M����OM��wy�Y[��a���Y'we̷v�k��8B?	�pPD&Uk�1�0�7B�}-J&�Q�RM�Ҫ��N������Z�)����Mm�G	�f�m�m���g5���@L�6����'�4�.=R`g&q�I<b-Duؠ�2�ݫ�}���j��Ng4uR�nɴyYaI�iT��"h��������3�ۡ�;��}��u둧�x�,�IŹ�f'�R��<tg��%6������_���q�lHҰ�j�[XA/ܾ��Le���R��'�VV�,�c`���uk�څV<.������D�t�8%�W�F�h������PC8q�zrG��#�t�Ҿj/i�u���GM|d�*���¾ҵ��8յi<��@Ȏ��.�ʅ��g&JMB��]G5�el
�c�
1�J~c �]��zn^���:]7q\�csq��[���Y%׸;,�M��&�OAM�۫�����e�m�p�cu���9ɉ�0@�I�I��l�̦��(I&Ļd�YAn�q�%3��)=��"eᑲm�n������MR��|�E;te7l D�ЏKP��F��8�k�����W�Փ#W�qa&|�	TL%��#ك]6�N����|v��2v�dq&N?+�ů��)�b���Lv�r�Qu[����4)�D6��R�D��ύ"PC}�4
�H��� ������>6|�uтB�
��Fpϵ�I���7�������q�r�C��Q���F�R}jK�'ǋՒ�*��כw]Y[� ��S��t�gŔR�h9+�A�؜.�Jz�o���b#ȉ��{J�H�SK���>�5��+$�*hV�f/.��3����W��_Mi�I����-=�=9	k��ٝ�"7.�g�n�p[34eXx*��3	:vj��/MC�wtO�w�W3����mc	��cJm��]1!��YKD�Lc�o6u9��umP���/����Ă@� h �����m�u��l�7В�δ�&	�&_s�cVB���(��4���1}���3���z��'
��F/V�p�w]~�"�JG��94�x%��ģ�pu[־�A��(^�7]w� '�)ώd���Ĺ5��^�ȐvJ�y}z�f������ �0��W�!Rz��f<�w��d��l���Ɠ^Ǘ��%��)��}����a�v�3�ĕV�&���Ta��7k=��H"����5�B��8�^L���iAF��}�s7� E���H�������!��it��L����{�OP�������B
p���Z�F<�QD��HR+7�����eqT�����6}JH��D':�O�4D?��(]�\��\���v6n�U=��P3�%����jʛ���#ibm��X�i�Xԛm�Sz�D<u��d�9N�<L��#t��A��@ B@��6�Ԋ6 �$J ؤ��-4�gw��+��8���;|��A;cI0V$�L�B��e�9�ڎ��}�_Q��=)� �o���0���c'�2���*3��L�x|��z�{��X��j���<���(Z�CHXg*��k�]N���B���Pd�L�ۃ�H��0�Z���c��/g��L�?�^0BkN/lw>0�=ac�[�����|>;�C8��m�Փs*T*+���!�S��[l�}��"&�)/a�zPw[F�+\��Ydy��� ���tI���7�Ue��:L���v:�����<�"=Jr�S4�m��(�rgY�s�ќ�e.�K��#��\��{���z����c�g�
W���n�F�a��t��u>��X�8`nҺ	;��"�+>�`��X�m�X	6�Og2��T�ru^�����I{gv� �G H4�����!�R5��C�B@�0@	Є���	 �@ ƀI�H'�k;�� �?��-�n:U3�}հ��[m��y���.���%�9 
�С�Ńﯞ�Ϸ��Ř�3�8�*[΄%��Jd������|�f����Ū��Z�܉���Üq9�׳>��@S+7OB��W���iWT2@w0O_"�֗p��S�7{�Y�8�����ս��՛�o��l��S�����g�A��T�)��s������x`��~�J:�x�u�;�����(V�w�Axu��IK��uv�I�����u�#h��ˬ�0������4���6��Ъ�^�)��&�m2�I��ʷ�wn�Qycm-�ͩ[Z����~ �#IQdD�* T@*��+\e�Ü�vkУݙ�o4��9�L�s#��b�]ccmr�q���F��J�dbB�������b��d��؝ݞ���̀�M�w��ts\*�1bP�����'�7ݨ�C\�ε�v�hE�����T^Fu3��F���>�h\2.MX�q��a������u	9�����r{b�d��OI=�ui����Xz*����8T���_	�Ռ���l�C��X"&z�;����w�96c���Aֻ�lBR�&����p���rz����1P$�r:�k�x�Gx'Ǵ�tT�H2I'�J Pm(���(>�h���(<��v$#�y�6��f���Ф�ʾ�\��"������l�-�e��)�
JHb���a���3O0�ݍ�jq��	K[�|Θ���N9�:Ή�Lq�ۀl~"D9��A�ܢ����u%=@�����|�3s��<�ͷ,h�U'^Vk�$��,6Lx͸g�"��o��oG�u���Z"���\�g�P�)lv'W�����A��L��	��G뽃O�OI�^��!�(�{���)�o���;��|)`�=�R¦Q�r	�`h��9��j'ģ��K�*�e�V:{�ë�3������6�;�?� (0���N�Lkj��Zy_"�\A�2��U�&$�C\���3�U�����d.'#$8��\�� Px�JdFI�fA܇ q��_pz�	��B3��Q�t�'7���=)�8 �A������?��i��2��q�҂��᥎Ő�8��~�vw�����p��C�2�E�d)J�>=�xz{̺�C�Ɂ���ѠA�-���^���>!��w*�<�=$X^�/@���#�C@�h!�`zt��)~�F,�����!�L�S��Bs,�<ƃ{���!���S����l ��h@� A�6'M�4,��"4�pR�s
s:�%��jmy�2�J�@@=�3� `�W,�}�A��5s.h�$�:\0����Gi�z�a��5:�Dp�g`�� ��׸[����܃q?!�i���y	`S��9���g�z!��z��p�n�I�#o�R�˞�_��D��厓��B$��*�;�~Bh���D/� ��V���p5a�~!���	���<}��&y�4�!���[i�A�q �y x{u�d�
l@�N�7�|�,����#n���Dz}"u	�_�3��e��z�pDЇ�0��q�G	�%7(3��\�0%�(�
v���(DP�1_�g���u	�=��~'7_I��A�_A�I!�n'geA�3 �tb��6C�k`�N)#�!�)���G�'7��ܑN$�Ft 