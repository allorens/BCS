BZh91AY&SY�k81ߔpy����������  `����n      �    T +xi!TT�D*JI%U(�H"P�      �@  }��  ��qy�6���j���l�uֺh�4�����o3�Z��7_�W�w{7kf����Ꮅ���Z��y/o   ��y�����돯���Ǽ���z�������T5�U�X�yկ}�{��k��)Vk�O�ݦ�c���v�]}g/^gw�  ��}�˝�v�Mog�s�OM7{�������zz�ׇǾ�����}u�k�����W3�{:{��:�����  <l>>���-c�v��y��k���(�wϳo��=i`�|v�m�;�'}��ӯ�����{�om˷g<�} }�����C}��ojٷ�����:�o� ��}���]��㽷7v����=���nT��ܫ�    (   
��L�5!���O 4�T� �  �L   ���%JQ���&�� �F&%6�&%T�6қ"b @�@h�	5	USjb` L   	��"DT�SI���
z�Q�=G�4�h1=@TI)U �111�z�M ɀ�ߙ�I	�$�Y���'�H�Ѕ��� ��O�5?���D�Gh@���
~j�ҕUQ!�B����������wG��_���`)I�$�DY5N�뮳�����gHGj!��HN& ������h��ȇ�����ğ�������~�1���?��$����H�$X� �&5�a�l�N� �$;$1'L�5�.��%�u���7b`S�m�vN���8L�d�@6Ʌ����K��	n蘩%��M�&	�B�*2	�d�M��e��y>f���Tfj��pR$E��k �n�q� ��AƔ�Ζ�͇m��ubSAؤ��&l�gYv]�Y#)�0)�6ҫIT���@�a.�VRf��ތpTZ-�f��t����v]��)����%�������.�U��(3A�L��eT��TK��vSf�)h$Ⲕ�f,��?il���h�L���U#-�.��J�
��ݤ�
�/0���ʙ	��e&R�+R����[G�����$�t�%�*�p�^�ʦQ�l�2�ٻ5�S��
vJ%Q)�H:R���zS'C%��p���E�(acHl�eS2l��UVI5D�)ѝ��%���&	�h�7O6�"X%��M'��Ka��-�ٖ��s�YT�'"�"�K��=)�:I�eD��Va�1v��J�%O
��ΪJ��qI8����Ri����ihL�$�"�6	H�K���·4oZX�I���V#-��zTjZ�-��딵����4�FEl�m��ĵ�Ol���J��l��RV#���:�Mc(࢕�v&�RT#�*��V���=����͇�Kw��P��5L�s�1dk�Ι �5Ff�)��.���2��N"�$�p����������:�)��E�Fh�6f����v]�T��N)���Wi*����_����=��k)�vId�JX`,)Q�e;8�Kd���Ƣ�(����4�dS>�j�Q�%�Rɗe6m2��VR�lŖ0��&��tSD�+�EZ2�[��tv�D��i���ueM�P���,�%�L��եq	[��8�-��M'	�n�@�	Nil�2���Ku�L�e;:�$�Y�eXR��8�-��M�V��͢�,/zSf)�lղ�"s
�2��
l�&	d�8b�)���2��6K4�''�9�����L�2�:H��	�
�d�&�٫ec;���vw1(��`tu�OI�ԥ�	dBN �eYcX�]8�-:i4)�M��sK�k�6����-��-i-h��4V�m��pS&|�%��i&�Z�i,i!G)ѧ)7	<���d���%w%Z(��=+[0ɬeqjYS����A���l���2!�f�T�9�@��[Ҙ�IV"�:���26˼J���~�AI��2Km*p��)
`��1��4X�ikғ6VZ��t	s��I�W�2$2#ɤi�% �ȇ�1M�Z�ј��eP�$���Ʋd�/	4ZN���F����#C#}���*�t�:)�v��ǥ0�R�����J�)��H=J�2M��H�!JJ%AԤ�Q��aQA�^RO��C$�TAA��6��)
`�~,cIj:��&�m'R�.|\bT�.,�HdHdG��)�(xS�J���)��ʡ�A�IcY�N����
�MX��*CZ�L�0�a���J���:2!�LS���Lc����~,H�sLkĥ1-]�l:��aRԚe{$0ȏ3��HT�A:J2�b]�A�c$-�L^ZV�-�V��/QX���'TR�Aͤ���H�N)�b��Y�*�4�t`h�E1�^�xl1l,$1^b����2��}��"DHS	�Aѐ��a������'YY%H�$ݼ,=;��%���2L2pN�&��%�m�@:�F,�,�,�����4,�+�W���l�Hl�ct'Y5�5�sH4 �8&�`4�Y �-&dH�C��Hܒ^H(?`����k$ΰcBx��pQ�O�bN���&�^a��#@�"��b�x�e��JC��#�n�b�ҷ�1oR��1�:��EPu):��0�������I8d�Ib%P�B�&���X�L�&�E�VR�.|`5�4����,�y4�e ��
b[J���3s��2�9$�f���0HaH��I�A��	���]@;�T�rHӵ�������]�&������S��,��X�E�X�d�0e5�2g���T�����s���!S��i!0X��m�wE���'D��F0X�`ة���0D1������l0��01Z�~�"XI`�p�~#)��1��cch0���H���,�bC�C��.�A�C���0�h�g�m"�)
����'�[ ���/�$��6��g��gF�em��E�EiU&��.L����3��VҶn�W�VM�AIZ.RO�K[Ԥ@Z�������,�LǄ�=V{'܀CdnEr*�9�Z��*p�Mp�:��71�ZR��4��4m�]IF�͎��r���������b������/�x���걟�W�%>���LGS;����_*���s��8���r��MƚŤvs �03�3;۲@���?��Y�Y�3�׭�~���ڜ�Q+��̻񗝹���l�Y� �1׀��֌H�-V������m�9l^ӧj�����eϫ=G��sl��7�f�ʻ�Y:74X�ˠ���:swn��V-����`�}+9���]WR���̉ӼF���?C{�J`��e����O�~��}���b�x]�E�G���k�)��/nG�M�����f�:;�l�!�<<�f�{gΛ�<N�6_��틭���j"^d�ݎ1G\��2Ix:>�n}&u�B�����a�1�e�FeXc\��m����aF
���lTx�,�Ϸ�z�=,���uyϧ��4�}�	��!ʠ��{��_�/�ߚ����Lr����P�X3	O��>��;�Y;���B;��w$4�3X�}����6oza�Y����З��Ę����F̫��y��m�5}�uy�A�͸
��<\c3�fM��R_EOBt�~O\g�ɝ��ca��܇m��*x��X�[�T�-��.��.����:�i��&�y��&Ѯת�ۆ�
nxc�����/N�j�W�N�ɘ)n:Í��;T6��5�uEB�50�2즚0K艼̫�(��6qE��f��u��m�7ۋ~s���@̐����M�馌�]��|?^�2'���<86w�?L �f�fL�_}�r
̬ˮ��EO�����
����"Փ�p�����]EImL�]�iY�2���'a��;�TQ1�{쉲h�b���*�Nܝø��!�8�~��.g>q~ʂug��ܲhB�����^�d�d��)�ᖔ� ��=�]����)��7�������9�</�<���ߺ��m�ӊ|f�&N�[��a�fJgmȸ̝�zb�a8��M�T��W
�,�e�j��S�B�F+Q�4�%�wGd�Q�Y!sVf���L��`R؛�׳3;�3��ȧ	��L}��Mt;�n����Čn`�&�������f�</Wsqv;�}e���z��3��öM����S~����c�3$�9�ei��W���]TOƲ"��*����}�fd���q;���Mf�S����ɉS�Xt���^��܇ķ����90���mMۇ	U�۽��̻�P*(�ɓwN&(�×56sD��wsfR�%b&0�Oe:w�,�E���~�|��h�a"�������K���k��7��;�n&4�1�̛��us�br�'"��nT���:xj�g�+s+.�12E���I�`L�YK�fN����ݛ��܋����֮����`��-)�~�i�f�NfFa9�f��<���tL��a�a!�(��,��3:�.��;*���n�LЕ���r�����]�s���,�ӵu�W�UHU!G!�w4�ІPt`~}��{I����t���M�{;���?̃�
��Ҧ#���a�ҍvd���O���y?+�%�L����1>�kg�9�~��apJ��Ó=���\s2��w��,�q�g�.s�Y�?O�c�m'�c��y~;��T�.s][��#72�Y1k.֥;F%�]&\�UܟX�Ңw&�Ĩ�Q���80r�ꛨ����';r:6'
(o<Ǚ f-��b�C��7:[�~�������~G��t���sro�0�z9����<�vX~���%�1yi7W��d7���&�^P�0������qvY0fUgLD�7[����4�'��Μ̚��1�|x��O�d�v)�Y��.#r�a,Nj��e�a����ŲSI��y��QL%��4g�<WM�9�߾���tа��%�~�=�R�!M�l�,�"�f���ڨ9l�g����f����ѽ?gCf�*��:d�7�N#����䌁�p��;St�T�Y��cxo�����L�T�u���)`��ͯ�EeV�Ǳ*F����$�d(�i�M���=����:SP⟙��l�����ä�;'����eL~�C��~�m��<�e��'S~�$Q�����'1l�S�I�8xŷ�1��(��33&����lXU�ӧ+�F�v�}�Zl�l�ܦݘnE����חE��ڥ�%q�3e��×���fAi�c4�S)8�rwN\lF��AM	����	�2v����3��d]DmjͽYR�;T-s���q-�qQ�^�?m��Oه�����ś���6w�N̘>��=���6���]��x�mp�s=*\�B�2�Òr3b͑��}Vӣ�=���f;���-;g2^��}���ι�4����7�Y�_U�N�zww2oSW��?M��0ƣN���[���"�{%1vi�(d�Qzﵚ�M����c��TAj^�n]�PҚ�w^~�����N�4Vd����C7�	���߈,�Q�.߷V;�T^��ٓ;=�'�+}(X����'�������o��+V�3�.wz��Fd��y�5Բ�ӆw�Xw_�{T��誨��԰O�Af��ܣbư�.d�6Y�]�{��O�LͲH������s�m��܀ί�bձ�-G�C?�O��	�$/�|>�|8xQ��+E}�����!��$*I���ϟ�Z��!n5����&[��i�p�7:E%u��3),����EQX�����2�?[�9�\S�EA��h4R��B�Z�}$�j-N7u� )����1N@�!��:H"��ݵ	�-MF�me]��[�\��4����J�JL�u��Ƣ2�Z�q)��tc쓸�!��H?{�6��8ߔ�US�ϕRy��=X����,'޷p�s�Y1(Ԃhi�G]��H�q�1e����>�W�]�YR�(N��rw0�G��@����Q��.��������-��ovgyZ�d���Bu�ť�d|��t��w3&����0�w�rdV��1mb�}���"u�S�u{���KTd���dvQX����a���!�6�Y�Y0�[-*��y��X���j�F�A,v��66�Ԟ[%߲J��si�Q9-�i�/�ۍai�A(��jr�Z��ddN�T�8�q	]U�8�R�KIENE�0x�@-��+u*�:J��O9JᎧZdlmBG��W��Z7���U���UZ��"
?�&��vƃcpM��ūUJ�uA*U��-�[R8�`��)"���l6_CM����ަ��+��q�
����⭖يZ,k@M�ƙSp�J��*p�M�0���]U�S��T���d��Z;
8�c��Ʉ#S�Z�*# dE�*)�1L|�1~C��˪��LMc������ "�Ȃ�X���Uf5��G#%���u�UTN�"J�D��fN6�g�g�U�p�b�TǊG`�q����[y!e��L���i��-��5wqy����pŷq���m?���}-~e�!�{Zw�w�I���?�5�d?W����|�}��|��U|�;|�O�����8���m��6�m��m���[iL6۶�m��6�m��m����m�a��vۆM���m�m�m�m�����m�a�m����˪M��7���$=���-$�oy���{��r�n�nm�m��m�e��oXm����6�6�v�n[m�m�m�m��ݶ[m��,6�۶m���n[ݝ�[��x�m��&e�m�m�k� a����m�i�ۦۖ�r�n�nm�m��m�e�I�m�m�M�-��6ܶ�t�r�m�m�m6�oa��6ܶ[m��-��=�����ۦ�m���33,6�m�g=� ���8�wEwwv��m���9m�m�m���ܶۦ�I���m����m�m6�m�i��vۆۆ�n�a�۶�6�6�v�m��un���m�m6�m陙��m�޳��� ��\6�a��m�-��x�m���6�t�r�I6�l6�m�e��m�-��oYm����m�m�M��m�m6ۖ�n-������m�m�m���UU6�6�wv| �G�> 6�Ko^6[m����m����m�e��oM����z�m��l6�m��m��l6�m��m�M�-��m��m��嶛m����q��n[m���s}�{�w��s��)"0"��!�_��A�����!$��w�������>W���A��?������_����6��zڶ����+f͛;m�zzzz�����n�m�m���|�ׯt��;6m�m�n�m�om��=m�ͱ㶝6�o=m�;m�o�z�m�h�M�[6lٵv�㧍�z��n�m�ح�6l�j�m6�n��>=>;>ri�z'lIG��luAAF�d�184ȿ��GJe��pQC����UV"
<��.�,{ug��=x�͖�х��A���9��.�:�q�n��薭7�3�rٗ!����)�8U�G`���c���j;+"���5#�E'fD���Fc8ĉ$�1<Vee���$p��Z���7k�A7]RQ���9���㻶���\g�q@��>\�_�1��<v��WHM1�����p�\/��]��6*�\*j1��9��FT��u֑a�:Lx��dM�ʬ��r'Tp�]m>�	И+M��Q���u��WȾy���^QƣV��d�/�����x�C.(��ps�4�jrX�R�2(�Bi8P$���i��2�d]UY�m�	�A&��������	Ҷ..r��^�L���C��{����˻��g�>G��9��9�}u��2�s��s�����ȡ����w.��A�'��޽�s�c;νm���j��DN��:=�O���l��%�c*�$�&,NH�3$nW��j���[��"F;@��#��d��	.L��$i�|����1���9Q�*�bU��� ��k�Y��yN$M�T�0�g��n�����T%kd��)�#���ȗ�I���kL?Ɗ[bK �EN^WM�������`�˿qG�q}�q]M˹�ȗ�vS]����	�����Q1�"���9�$Ky��71מ�N&^NmƄ�����i����õ7�"wϪ>�$��������xb����j��Ȃ	��4YE;�ux�]����Z��W���%�����:i�L�є�E֊�J��1̵;C�`g���IF�.(��z͘וUq�7���S��E�tx�mU^<i�c�uc�b��ɿm����>�I{�<�9�g;��-��2�2g�`����������ev�G��6Yߚj�kx�[�����Cp�ga��-T1M�v��^$H2�A��Mz��I���i���������U^�i�c����i��Y�O.
��ek��#^j��=��m<�e�
���]RTc��I�a��pmS!DdU;+�V�Qe�3��!E�>�mn�Ki-pMa��E�$�n���x��������)��r��r�Ov����5N�s�4�L$aY��^�g����i6���t��l-�-�T8����I�H���b'B"&�4\
�RU�V�)51
�C.n�ɡF*l�)ĉ�Si�8�	�Q7NN�x�M9�ǩ��]*�(TKb��G��p�ɴ���v�{�z����29�((�!�,DC�䫶����+u�{���$8��q�j�&R�;�z׷�z�)��e���B���,��컲U�L�󞤳;}���U+�����a��}�����+j�U*x�<�k}����փd�e�Yf1���II��m+n�8{��+N80�/KJ�rH8UTU�)#���䤴�w�Ě0ۢ�h����ͽψY�m�z�
b��9�f����8�`��%��3��e�W�����$/�(��(�?Gƺ�"d�!�zI�8(�ʇq��cM��%� ��a����ʚ�֓6Ԡ�lk��i�|�f˸㱨P�JD�V$FJ����[V"�<
��+8�wm�#��f.1 ���
����$"{I=p��c�����"y),.��0��h�<�5eorZ��Hh�Q��3�޳���r�å�iD�Ғ�	�NL��&(�*�oH�()�6���,��c8џh�kͶ��t�,����a��ۧ4��BB�F7�ִ��s8���CHQ֣�.�Y��a�U5b���m0��.[��rq�j��Bu10?s�B�Ø9.U��q�'|�Լ��+;U����0g�5�(����?�GCCC�8���v"t����k����{^+�Y�q_/��ی|����X�Z�+�W�UǬ<6?	�FtQ��JZ:X���g���������q\_����l�	��6>z���G�t�+��1�|/����::ͱ�G�`��RK,�WG��%p2�';#�t��j�����=fD����~�D���kKZ8_��'GYbt�I�Bt��B�^1Ƹ�/n3�����Y�j���D���4c�/�����ɱ�r4ذj_��٪�'ENxŕ�ӎ��j���&��i���=�g?������@5�K��.b�l�v�\�g���q�US,~��}���U3ß"�;�����xs�Wܻ���xs�W��뻙���.$ww_��kYϏ{�UՑ�,F���<Ye�Y��K�����(���&Z���)��B��q)L�2�� �2O��a'h
#���퉃N��/�j0J��ln k�Z�j��1�X(�V��t��&� �*eOc0*�EM��ٙ���AC�Ԕ|�d�m��H�pfx{�T4`$� �6τ`�O�'��u))<�6D%J�a���q�aHh0PYb6���e�YfC�(��QEX�����$<c��ʶ��Q����53�����(E����#�p���:+( \P`-��<ݩ��f�P�.���Z�T��UU[�' T��R	DE��B�����'�&�Ģ)�)B����6�- ���4��i��}rAr\��t��0�ਕ(X�_̞�(�TʍE�=>a��mv	���,�̆9�O�}�Q���P�N�Lyb�r�U:�W���Y�"d��r�4)�Ѐ��	2d�3Gs*BQub�#�댕��N�����:E8� ���cN�� @��A֠�BSXU�CI �E4��i���ޒ��Ax1���O����i��2��񖓚+	�Glp�(M�9i�������
�ܠv:l؋J=w4:J��~Y��"��-�����N>m�X�`��&�-#�&�e $LGw��.��k�i"���|�1i j���.)���$�t�mab�R���&��d�'��݁�%�� a�dR���lB�!,�
<t��,�$�-�M��.�j(��(A�h-V�eC��+Q1�ڶ�SHi�2g8����F��ι>bʞ�pA�������Og8@��5;u�vY+;���o%?	�3�Q���B]T9Vrp��.�	p,�)V�k:ڈ���E8��j��y!E��S��2�+�R�Dç�cI�0�``�)GsMn��>��,���M,��,�g���c\�[�����QEX�.0���%UTRi2L�Ի�OS����.怬�ˇ�yT��J(�1�$j����V@N��qcf���QAS90a4���(0�9���y2{_J.�g���{���-�,���o{�e���ڪ#鉣ET*F��
v�z��N�H��L8<���0�mp����|�M4�N�a�����c���+(��	��w��s���;�~�ZX����ݛ��,h�xY��ⶅM�T�N[ͩ�"�`vq*֦Rk��p�����a�D�.&K�t� B�7��GY��[Z�c���=u�zj�$�(��@�&�%S��m���a�4�p��4�M:M�u��o��EP�Ъ
D��U��Z�`x��ׅ�U]DR����[H��dN�d�MQY"|�y.+31�J�����ڔ�Bp%TV<�Nu8�/�E�̒��i�/��V �4jy󧦀�w'�^r�&�`M4m!���3	iI�U�/�k|P����#;dۛ������v�-O�|Σ2�˥>�s��F���̤Bf,�\�
0�I#�N)I��G��Q��s��aZi�vi��Ye�w�a�%�+r�rR麦8վa�W&��rPn�M�2����`�6�k�2�G6ձ��=t���1�()!4;i)�YO���CPo�4��NQ�gW��˕b�n78s��X�d�u�Ӳ�!t���Ҫ��[J���96p��!�bC�O���,S�95$���XlȔ	e���?=cӨמ�v*�G���W�ܭ�`�;�i��MX���S�F:b�x�w�^����0�i[�V�����Jp�%�j�V���&�����n�b:>��
�LJH!G�N�e {Q�w]L>��:��>~7����䌐/i��+BO��t�Xx�!e���:"%����B��<Ǭp��(J#|���zk��)w��ն,J��H�B�:�.�c�u6�C�r�	�܁��>|��}U
�P��8"@�!lS�_bJ��Qf^L%��'�(�Et�p�X]��T]\�����CF�4��(^��a
0��Ux�|"<,��xSlDO�_�?1���ژ�^׊��q\_�����[�t�X�-^�G�<p����z"=:U�l��'�
>�#��+�x�6�;ck��g��Lb�j��HC���+�:BΎ:�����pm�&�K�8N�m��#���gG}#�p�!ӣ�t��������s�q�8�1xv�-^��s��OG'��O	�d�p����I�^*���x���\_c�̕�xU	ᱣt�>�GGBܡ��N�/���ީ6��<n:*/7%t��f)�ɘ��f-�FᎢ7�&L���
�]�q�2�m��-��\y��N��n��Y(��"T����T�<f�#�Z��Tc�Mf�����\��{��N��e�g��f�;�P��*��`4�as����W��6�)�as^Y�d��<L�5���,�{S&�4�%ABg#� 84�����F X�d䱑V���D[�~�@4�w{��{���#c�9G����$�:fl�ݾ�&r�,�|�5�ϿL�o{"��#��`��L�>�?Y�����!�����d���QF\�fY����lB�"�{���#�i��LdDu:�+%u1��Ьv;��U�5�(���1�;#N~��b�DcDX�v:�V���~�����M���a�8:ڑWPOc/0M3������3�lD���j0 ����J���D�m��U4�tQ�X�bq5m�ɎW��������?�I3����ww\;�$�wwOe��p��=��=�wuû�L�wt�]���I3���՗w\;�#��8p"��N��:"%��gu5�8��2[Wj��JIw"��j(�PQ�����nU��1�ʬm�bdRr�3.6�;NX�D����ǀu.)���U$$�H�%�Zڲ�ğ��t�<M:L�<̶���1�2�n���5`=B(,G!�T�=�+�F�'/c��4ЃO#���jv>�:�Q��]�Ӹ�0��~�U0]�����&$����{�fI�7��{��v��h��ъ��7��ܗ����z�7k��WޜGMBX�г�DD��y��0�q�h;�l�ِ\��o��\ʕ�?B��
�n\�H�I���Iov|�%���bXp�iv�Jr��
|�S�D�� J���{$�&�'RE\"i���'wS�
,Y��5!��&h�e��WusI�v�ƊL%u4����UU�/ut�1Jp�y�X�M�2X��Y��,�kھy���ll(��q�~ESé�iU���``/*�X��Fj���Syަ�T({�/ ��4�])�j���B��45B�B�P̠5���
,L���=L�pd���oN�. �}�5Z�ss��7�H�z��p�L'!�d	�2g�g�.&۬�- m�4�?x�ƝJ�{�=3�+��x�������i4j)~��.�G9E
�9a\�W(�QX)��*����i��|��,�.�EG�^-�,�v�	Y1yr6v�;Na�;3b�Fp�`	��-��t�l>M&���%�	2B��+�d����4SIN]��� �Գ�Mq6�;H�_����i�f���aX��;<����c!�V頻��k-��4����כ��E�;=[�9(�Q�ŏ#Q�6��#���-'(�25�r�U"j�%�T�4�UKCJ%���LÐ�f���M�%-&Q�SzI3�6����9i�ͤÄ�E`�=e�%�5`n��%�R�5����B��I�˄�[�Οr�n���YŘ1�,�bU�"F�O��� �t����V-��l��	Bh��f�OT�5d����Pri����F�G�5�Lv�<h��h�KB���R�a�}��U,��M��gh�t�i0��7��xL�K1x��c�%8�TS���jv3�E0e���b�`��FZ��f����0�U�5��b�U�f/�NG�ѻ�a0�-8�?Uf<�y�?<V���U�!`+��EX%�2�aô�P��A�,Z�K5$���?Q�t�!��=;��*��j��%ߵ3R�OSi�����8c�}D�>�v�~�'o���0#�3h H�UW�NdR�hXJ��|w��4R6��N���䐛G k����g���|hJ�4dD�"'Ř����Ƶg���k<f�S�9�=Kx��7q��V ����(�h����rp�"�"9��n�����Ze�d.���c��0�m=Ӥ����z�|t�`j'��j�(�F���F���.�Y��i{5z�K98+��-�|�8���e���ޟ6�+��V�*�i��_��7'�^QB+|�7�E�%�&�Ln`�D$�c��,h�����i���+Y��!D�僲�!�8W���T���0f��c�)b�楀����t�y>[dd'ɷN��{�M%�II�I=[��.�!�"a�z$����n�%#�'���D�&��9B�;���+���L`S1U�5��\�>2ͦͩ�e���!�ĠJ��|"t��N�s-���c1���ʳ@�L��{	�Xx�ɔ��u90a�@7�s��5��xi�a���ut�S~��iP1 �-�)͝�V�g](�!We�K�K�`�LQ{,���8����`N��>-:m6�S�rB-0�� �G��Rʟ
'E^%��J�'���zq�\^׊��q\W�\q[^:g���1x��p���������3.ا�'J��G���?��<l���8����x���j�j�^
(�D|3�xl�G���tW��Η��ӂt�8=8;4���:x'M��Ӄ�p�'�t��ta�tt�8Η���V�/¸z���c�0x>I��'nE'��d�_����~g�����\~fƇ��Ĳ�">b�ӟz��X��>s��T;Ugi��&�H`a�I��I4�i�i
oU0�LBV(ڮ*���tm)X�S����!��m�U/ɔ��i������N\!�-���ߨ4�C�P�@�.iha�d6��iY2LuXe���(�8�E���mR�:큤�8a��ӗ^��u�d`2�ܦ? ����˻��������՗w\;�#�����.��wGOwwuV]���<����ꬻ���y=���U��s��}���b��ZqU�N��[l;���_9q	��&]9ls�to��$�*|��������c���^5!����ֵm�[e��u�i�f�N��Q!�0����:^ �.eS�BgVl�'ws~{��y���t�4iⰬWoJ����k��a�1D��!M��D�{F��X��n��/]y7�ܗ�W/����H��KZ=����Ō�0fjjV�Zih_��rȁ٦��$�xڟ�	'rN��O79
0;�Qf ��L�g�*�|*�drv��g�>���o��b�,B^B�U#?�?5`M��W��t���0�S�H��% #��Q�ڊ�fk�l���A��2�A[��
��{���&H�tT��E̶QF�_��y��K���W)	$�:�7�ru� Q�&��O��:�1z�t�rB��]&��4����`�U�+p��*��s��w0R')>��Ǌv���xI!���g�>�%��+$�qYH����ϼ�<O}6�4�.���c� �҈P�Wo�?1^:ttI��7W�wg���е�!���GU$131�@�-��N1+��i�樔a�GŁ{�-<��ӘL%��`��i�+jnA�*h���US��G��P��森C������u�ɎG������.���^)��7�g�M���[[��W"3z����|b��wV@�W�3*71l���Q�Vl���T�������o����^��nxǽ{	S��/�G{T���d�3=����G�Ѱ�'. b�c*�k'0�*S�b�:����<j=�?nko��1tۇ��Dk|�	D�h�������1�+X�'6b��y�7N��gǀ�U&fd��)O/�m�'������3WRIxfH��TT��Ѵ;��/�?�A�����#���t��o���E
��5\= �6B�А�a�U)a
�(����tmj��$���S M'O�%�m-�a��+����7ei�kL�@~N'�nx)�]��B�'��́��)0��R���މ��"�Gs#'+
�|�Zc�	�Øp�t��r�.T>�xtUZ�j��W*g�7]˺D��F�u)��;i �-i���&Ȫ&�7�c�k��*��9�X�i�FΦ�ݺ?&�:����u�h�j>H���т�2B�"l���R����l>��&d@ �<�$,�^̉�}<ED�a�B�o��/g}�@��b7�LDY+/"���,nZ�dJT��&�S�"v@<�����ı�n8�&6���
��D��������}�#$?d~L�9����{�V�l���A��	rImJ��:O����^r��z���anlL�1�s�N@�d��(7�<�$$-c.\�k5����sP�6C��2��G��	@�'e���=%�2��m���5WZ� w�O�Ｊ�)Rڽ�\o�d�$�ʝN�H�p��Kx��k��;>�cIN0�N������,�����Qo��_{T�2�`�s��WE�j����G+}&x�6�+��O�8��Z����s�*��(���t����O�I���,��Rx�{Bm�F��t{YS�c5G9��ʻi����G@Ä֓l����e�2�"���rC�0�ө�>O��ߍ�� S���^F��pZ|S����|t��+鏛V1�G5=h�M%&@��?	�?�6)ϥg՛�go1��,���"&a��o���IZ�!�G�4�tա�Ϸf��%	���h�{o��ݵ���S^h��>̻�P���JZk~l���;⏡��vf�
��(G��g�#<*��O�t3ŕ���v�=g�q�qf׋���yո���p�/lg��>N�)�����:Q]��~'���=�l��Ht�:'xu�$OS�Z
7��Q������p�Oap<0.���C�,�����X	�D�x0�����<:�1:^�gG�,�nE'Bt!Н	�p����6;:�3��`�^.�Nun��U�\+�������|3�E��+bP�lhN��!~���:�g����d���0��vwYj������^��B�L���>'�;���f߭�[[�����G���Ic��L���I�b��1�J1�#oC%���>B��LO붔Qۗl�vn>~�ZR»=)�],VW��-�h�O1���s�����t�X���+I{��w9Z=;�aa�����(�H��F���V�p�ƿ{T3�����ԶWx�y�WٰB,}�bm�[E0r�ӵ�B'7?[�St��2�֙�3n�qdT+roe^p]Ӈ�a�͗.Q�iJ>U	��>efF'��%B��;����l��z�ڏ�JHp�2�bC�(A?J�(!�%Rz�~����%@��Z�6�T^ڽ�]G�s�6����U%�~$���U���˃S�}֚�Nʿ���ɩ�Y�B��P�Ģ+��!���Ṋ��޷�kg�˜������i�UQH�*b"�c�$�u�W�wø�8{����.�q<0�wwUV]��xa�������{������q<0�wwUw߾y�9oX�±\1�f1Ƌ��:�/�Ɋ���'eku݁�Gu�URLlN�X�ɒf6���%#őZd�L�P��4�v,#.�œ��iH	5��.�����N�gP�-?'\4�7.d�
�ʀ̜E�
,�5%B���y�f�^6P�D�ID�i5o���;1}�T�jy4!���KE��K�w��r1�>%��m9�ju�C���'��i�q���^�/���f�W�v�w��1ej�1_�x��>h�~+D|p��}��cm5:��FGL���z��ˊt:��W������g�US
��]/��U愣��n�-���c�.�US�Y��S��wH���h�|~��f�u�bt��Ɍ?6�+h��:@�LMő��BEB�P����0��h��8��;qT��nP��(�T
ϖ��ތ^��>�8M֮&��j�1���oS��ı���O�*컪�,���X�d�6=�09I8�ߟ:N9�"C �4"'�{����͈m�vZ�(��^���2���]��U`.��*�
�F��!�?�\�2����;:�j�?\�{�{x����K�P���v�!I��N�;O<x�"r��I')��C�=�������uY���z�i��c񏝦�kP��_��.́y�ʈ0�99l>���1��D6��M�ke*�MWZ�$R���(�#U7Ï�U;�F^A������>*�Ԓr׎6V:&�-�R�n
i���E�_f�D�r*V_{�����zY�:�$a���(0�n҇)��Z|@�����j d�(=>SJ�\U�����GR:үa�Wj�t�cj}���FN�Ш���Q;a�r�ý�O�d�ϡ͆��`Qrzb�DQuV�(��4�"EFv62A���y,Or*�+�5�����a�r`��Uҷ����`z<8U���ra���qU��c�O)-�,P�C��z`��xv��gbr�lQ},�bj��5B�E� �FR#L$I�ɔ�?8�D���,�Rz��sb��槏��@�G���/�[?%7
�V]X��"���0I�p���`��Ƥی1�ګ���O#0�R&S)�OD����Mr�S�7b��G���B��! w�q�V*\��;3@`��q_O����l����ug��W��cI�gjI�V�A䦒�)A���}Z�u߭�nz�u7嶪�|��mU5���B��>�6���G]X������� <E�8f:Q� �Wȣ�WL�X�:26�x6���8�Ԓ�*��a�|o�
'������J.QA`�"}ڗ͚=R��z��J"v�Q��C1�&Ϗ�7�m��J,�&9Q~�����t�[�~��h���c�Œ]Yw*�*��$t�r�����5/'�NGo�a�Wj�x��⧼�̫n��Ǳ��;�p�0��Pe<Q|i8)�if�m�q"i:�(r�0�9���A]���=%k�,�2���!��5P����󄴡4�,'a)7�ŕ�#�#�D�
�]�=*|X�z"L�zD�=��}!�����(��֬l|(��G�&�b��>(���E~W�t�����?1�~v�qv�&�Ñ�Ԩ��H��G��ΏL��h�'O������4q�&�f������fD���9'G�G����'M3C��t�>�������t:/�����.�<6>��<R>��\g3����g�Uګ�=(��K(�P��8�Ҋ�g=�M�4`�R֪9��&U�B'd���/u=�����n=äDꑴ�q�Q��oBۺ}�SFN��DBnc�ؘ�b	(��b��X4!=�UT��|O=���UYwø�{������q<,�wwUUe��xY��˾���;������q=GÇ��'HC����=b�[%���xǩg&�Q[t��݀`�Ԩ�?�x�������%�Y?�	���q;-��:���{��Ϲ�qn%8���NpK����Sx����L�K3�����ٶ�c����9[����2(�`s�̸��Y�U�+1���*�=�j!�o��ܓΐ�c�,�q���	��7~(��bX[����H�q��۝H��SO�1�ګ*�x/���D!��(��n�5!��"�m��L"u̷2��ev!7�JkY9�!�dx��h�)\jGȭ���!�ds��p�8ƢQ����B��QM����S���	Uw1S2B���aE�Q���/����n���'��*�����iԉ���o��.I$��K#�m�8�H�O@͵��*�`�`bs^i�����9Q_6��#�m�cmX��N�N��L�I��}�5IFG)�5��&D!�M�M���,d�.̠޷^&FL9���2��_��^��+ ���oI m//��Zc/�̭�d�{~N'ia�������K��_�]�v���kv���%�D�����Xy6��{IY!]�SD�
�F��"CB%:ps�_���+��˛�LQ�V w�0�𨝎V.I�i�k��w�����ļ��S�h@�z�I���n��62��u���o���d�\�l��
��4��@<G��]�0N�i91�����V`8�CM.a�ɞ��*6C\Qf�ndw��m_�X�U����7�cA��Z,<ֲ"�f�)�q%�K<�fS�ħ�?k��>�RUZ�e-�ɴ㤦�6a生=J�ib�l�鉯�8|*�Tv �R�b0m�:!S��ѶѪ���FnΕ�6t�v��X�U����;ʟ���6��\�'"d@�s(�˖`'+����rF����S����,��"�Ek����'ÕJ�$�D�jhLS���MD��IWS�Jr�Y9$��o���.�{���}׽KUT�
L��B��C۴y�<x�8�:�K�;�����y��9B��He��ć�!��!�p�gu%��p/�_����O��ƮS�j��-*���-*)rƑ�0����>�NG�}Vf+7��+�~Ucj��&��X�j<��5��y4�a2�/I��WwWeՕw��a�u�r|�Hp��;2�a>i(+���dC�F(�F�ju*�7j<t��HL/��r��$�I���gfՂ�F��L��3	�6`(A>b%8h;�iWUK�
�f<�k\�Ma+Z�| �'-2��8O�&��o��ڮf�k����ľ�:!lO*(D卷����'L��}	&�É��`<��ƽ���:t�m�d�6��5�va=tx�v��X�Uǅv���E��wCa�9�FY�!�e�&[D�?j���H��1>g1s˔��s�W�B0�Ȗ�m����b��9C�#@��
)(j�����D��Z~�3UT��ͥ:"��G�D�*��W��O/��+Õ�G�F��+���m^���^4�.�e^K_��	�>�N
�W�Bl�M��D��'�=!���=&��q[q�������[W�Uū�Bt�d��$�&�L�����L	�G����Y8(h����xj'�Μ��N	�rN��	�c��hN�W����ʣ��
>C�����Y��i�G�,�l�q�x^-^>W⳥�/�ş��DMң�8QS�e(38���ӮP����dSw���0cv=z�lnR�R���3V'��F5bq�&���5����.�u�3�!>�֡���&�M)j)&�K��k� �T	|�7ok��1���"{&(Ƭ�3'����ז��^k2d�n`� x��B���m[%nR�W�ˊI!1���$��4&ܰ��fn%`�D���&�`tV����v(�^w3W�D�n;Pج�H����YX��&_fe��>^(E���5D���&'X��S���pVL��d"u�ׁb�I�ȭ��X��*n�h��*�Z��6�m;Zt�����L�6�H'8�;n,�ZM�H�����Z.r�T��+���>ꘅck ���&$F`�����
��X���9d�8�T�[d�-��#"��c�;�2���v�*��dR���;TD�)8ܪ�����=G�������w�{�����/�q3û��ff��q3»��ffr�w<;��ffo�w<�� �	���4\�{]��P�y�.*�G��#�,j
V���B�B(�j�k��c�[�$8V삎��-�Er�M'ȟ�V�+��RJm�0�)	�I8�,�V	~�'%N8N%�Hi)2�t��I�ތ��(c�'��0��sׯ��^�|u4N0r�ݡO3$�i��oקk%{D������oWwDl���YVx(˔���J:��빼b��w�0�'F)_�����vĮ�J�@�u,8�:�և|��O�HC��b�S���r��M,3@y�@��YFD�Ub""Q�&�,~����#'J�$����v0ٰ�?\,���9�tA4&�J8"h��c��N�2ZG0�!����<|�NA��Qtr�s���2�m�ݫ%��<4�j�ٹ�\����2�M�Fe�%*���^��5K�=������F�N��Mj��γYn����`gf*����6�׺�H��B���Ø�SR*�~>�r�?C��;{;~��ιz�N4���_	���U�fb��ZOK)0��ښ��&�K���=%��=����j��a���/aS0���ݚխЗ�1�0維`�����╴��:w��$�l��^B�bƣ�c�.ffr'����H�`�ra�;2s]��!>,t�bd�����9,EP��^���8򧞳Y�+#��aqE�D���^��~�W��cK2�m0�˨FH�e�->���:HI,�!��S�l��t�2y�Q�hTW�.;=�h���Z*��k��{%ł�ۈPk���8�\�X�?Mr�|v<:R�S�8�1�:�0�}��IJ�g��Q�m�N%��g3*����4�p���q���,��吤�+N���&�=�e6�Q��C�!OSM1e��Q��(�gP��&�	�4;�FO
���s֍���Q�=<��n\�����2e(�i-:!��0�X�����e�5���a�p�����P�j��~��MA�r(�&ӟ���ɧ��na���O�j+�e��R�l�ƽ�BopN�i��/e<�k=�Q����Ah������(�yU$���횋߾On��d�����"��n��զ[zȂ�M��Ԑ�uI���p���aL�&A��j��
F��N�3tS�Wk��f��C�;%ț�ܻ�p�.��}�3[���:x���>�x��*)V5[,����UF�Q�qHZ�nud�E�Ln�j�R����."(��r�F�̕;XjL��&�$��
�o���8+r0�f��"pA2!�QGD$�1sY �2#�	7MX2�I�a���uah��[I�-V9�7�2{/45fy�N7	"�-*�	*���p�~��&�g����m!�k#ԁ���&O1/6�dm����`�c��i���Uҕ�1�� ��p,l-���H+)�"��EZ���N�:�V�D*+"��"�Y	YX����8ܑF>Q��u�\R�V�Q�t
�piC��C� �!AB�QT4"�UM(ȥ���1�,q8D
�ʻ�n�	IĢ9���'��	��=.NUj���ŵT�]&5f!�D��u0Ɋ�2�6}���ܝ�u�]�e�I����I�����j9S�W�V��X�8�z�&��U��!��x�.]�wwV��d�4T9�Ed����,b�U�e5�=TU��%q�6m>,Ä�m=�}*��+��ww>���٧��5L��dUZ��ؚѣ[���֏6�O����j3��:x|q�m�M�Ӧ�i�����<m�x�f�6l�ӏ��OO^��t㎜q�����i[6lٶ+m�m��v۶�x��m�m�<t��z��m�co�|���<|�m6�li��6l�]�i�o=v۶�h��f͛6�f6�m�|x|l�!��Hj�QT
ήIL�BT����n�׾��Fˣ�O����'qGW<2�	l�fY)�A`�(C�
I�+4e)���'�a�VC�Rj��)ڹTRe�LX�B,�'R[%$�%�����u�	i��a[��Hb���zI�o4eÊ���T�M�t~�5T�;�.z���#�j�g��n3d��Xb'�0w�7rff_���&8wwt���p�&8wwt���p�&;���33=�;���wwL��g�c�wwL��g�c���+�q�1�q[񕒱�59l	Zf'���IV�H����������c����I���Q�r�W)���ѭQ�G�g���G\�=�k5�ws8�&:p�^M��f?j{+qSҿ0�ʪ�1�~u��me��{1ų4�0�+�%�f�&�3�w��[��_~tQ�_���5v�'�s���OLg�]�r��Dӧx��HBe����gowl����^�ё�w;��Em�<"'
6QE7z��sm�u�m�ht��n��GoF�bQ�&!��]Y�d����ە�O�<C�Oc����cN���($�[��2��X(��Q��7eb�eG�r<�ʾ�Z���*��\�Y��'��L�4Iԉ1��KORe6��q��o�&��N�k�UT�%�O&즒�i��C�*����E�Y���*�GE(�a|mG#�YR�1�IRX!��mf��k���N�JW�+�Um��Av=`�ǽ ������p}���0C���_""Q�ў�UرN�͍`����'��s�c����m�7΁�i�ӄ�Rq;�%==��*fͤ�ui�)(ƞ&4e<�4�vGv����U_�W����c��V+WF	�10�|ZZa�S�l�����!����>�a��T�_�b�8SIU*�鹉Pf�K���y|�S���M����!�/CE	������3d6�նڇ��N5,YqN8`�ˏf��;����;I��S��O'gR�19���%Uֈ�I�F�S����߄�繋չ3	T}M�M��v���0������Ժ�n�L�FN��/�K��u��y���Zcx��X�Mugg���[h��J�\
�Z���Ҷ�ؚ+,����	Sӊ ����Pn ��9]��|T �j��������84`�!"(�HԊr#0�V2|��%$~N�i�y1F��i��-��i|J:q�i�;p]�r��Nn���͞���x�m�	�۽���x�"�����vb�&rm��K�i��+�Q��kU����U|�⪸�lc9��C��D�u7��*�����L>zZ{��4���Ou�j�J0\���8�F�J���7���naR��Y�}CTdm
أn��%�EI��%SI��:i�;�$4�B�F����&72�1��$ ��t�!�=i��^�~�^i�w\3��bx��y�%���da)<m�֓=s\O �g�Ғ�[)�.ros�.�i��0zf��9�ڎ��zU4��OCM�tI!0񉇉��2A�CBpDN�]�����e����v����*}�>>�gx�x���o�W~lW�e���Bs\�;��H����J9X�(�{�E�{�.HL��OY���;F�_�Vd������$.!����;G�oiE=M�9Lk9}!.����T�&SI�e&�\u���N�ǧ����mnݺm�j�o[V�<mҶlۥlٷ����Wk���n8��i�<m�l��m�M�m�m�m�o�>z�o�c�m<v�m�v���6��o�|�����m�ٷjٳj��N�x��ݴ�M��lٳfͶ���m�������B���V6��W���a��E}��3���Z�6a=��O���U�x�
ݝk3ź:7�֦a�7�uw'\L�ג���ֻٕ�keo�k�}Z?!��ݒnq�f@ܤ��7-q�I+c~8�C�9;\z5��ȵ��6-��+fc��Zd�V��c�c$-�̚M�����k:N��D�IΊjae�@A�(4��Ux��������SZ�C}�g�fv�.
�J�Hn,"��N�SG�.sr������L&Ku�{;lA�Vc���]�>U~��K�;#����.mz��#�VcǙ3ws��d�"�z���d87�[��&����e�[ډ����{!=L̪ 1bn8�����o�O�M"e��ynF-m&�j,]�UT�-�*Ѓ&b,�#�.-�Un2`&��5Z���U���ʤ
��l��%GZ|�VmX .�!Ev�Tn<�gc�2Ѡ�R�A�'�EUJD�
C���M�(�R�8�jI2����ə�p��c�wwL��g�c�wwL��g�c�wwL��v��c�wwL��v��c�}�{8�1�q����O	AG�D�G�M5���_M謩�l����Le0�6�C�؎���(1E$F2W$�%x�j�J�tT�m�VT'y�L�BrƬH�S��{"���k�%jdM;c�![(��.�$�	���ԓ�M���&��U+��u7��1��Pz:[�!I��[�%u'�Z����|Li<B��Hk~��%�hwF��Fk�>W��Y��B� ��=b"h��w�b����x�"ұ�Q(�ӣf�V+��ʥ��V��i�^�ZrY�FMl�8j�'̳bl��m����*��Ÿ�ˆeC}�}��|}��'Y��fgTU�����X��h��<eC�4ac}��Rc�t�Ƌ%��A��]&ᦨ�W��%g7��E-�x�^rI0pd����;�oj�����R�l�!�v�{O�˙3G5G ʳ�c.�5Z7(h��B�<7ij��<��\�y����񾪢d�5,�,���ݗM"U�CP�	9��=�=�`4ͼ�=��M#+<Ͻ�t�U��.b�>���6��M�駞�!��$�	�d~����F;<<a�<UW�v��Z��S�-��s8#�&� ���[y
��k֚p�|��w2� 'j��̙r��ئ�6�RHL�d���X'�ئ�Z&D�j��C3w��tK��rQy���]��e��*���c]��s2�Q�h�z�V!��o'�R�GS�	��y4�-�0��w��r�<s&�G�yuY�K�]5b�Z�A��;j%�Y��	���=�+/�RA4BȜcFg;5n�����i�x`��M��:�6����4b��჻����/��\����r�-�n�#�?{�G6���Ti�:�*��W��Q��4kG$�"���U��B��!a�DL�2'D�:n��px���6�|��Y'�;v�]��HA�e	Ee��w�Rڥ�׃܍�ёө�32Z���ɐ�иpB]� �L6*2��r�o�:C3
�y�Q�OLf(�*�x �YC�tDM����+Y�mUV�x��|"��C{5��Oq��Q6j�M8�E7Kl��.ۣIN�d�t��sFS����C)��1F�ߜ��x�w<o�]lҊ2�.��YVSN�)e���XNg�'�`���Q�ǌ0�J����6�2�s�{�P�+\Z�pN�s�pO�a)$�r��Z3I�f8��q�w"&(8	�0�
��Il�K���NI9��[qJ�O��bcڵӶ��4KKc�-�O����3���O$�Ҍ��4��6F89$1���%B�8;��-,��E��jTg�';M;J;��a����6�1�+��(���vQ9uV��m��vR�჆�@Zs/6�M4���*��vIvcK�g��'��AG^MW��\bH��&��R��
��gH�zb�������Ǯ��F�z|~?vzxx�|ڽt�m�m���m��ϝ�Ҷl��fͽ==q_��Wi�qv㏜q��x�p��m�M��޻m�o��z�o�c�m:x�m�t���6��;m��ݫn��M�[6lٷ�x���޼z�m6�lV͝6l�j۶�cm����^K�y-T�y�}��r��s�X@��@8o%�j��8Uq�E�V@�ҥ31�#��K݋�e���q�h�(\a<�����Im�.B�iVո��Z���2��YsUS3;��ǻ��f{��ǻ��f{��ǻ��f{��ǻ��f{��ǻ��f{��!tN��ӕ�T%u3��"6{I����m��.v��I7�h�]n�S��eJ�P���7٘bz��$�Io�"o�s��N�m�6�m.��;�<�ml����*��(���1;����M"Vp�z���błZ�ݥ�-�j"ʘ��G��z�r����![�9��҆���0��ڻmE���p�u����+��s��4:����C���z�
z�qU^1����9��L�Np���S1��n;�B���.<L���<Pb���\A��[%B��KlV+5A��B�9kq�&�y.;��Nrƣ�"����ä�q1]��&4�G��d�]>�yKSi�$����s�m��uM2����yH�O�����mU[m�w,�a�p~���Uy� �p�!�2"&��I�f�(�Mܒ����	��>�j���]T����6�l�s/W�ظ\4K���>��Ӓ>�=���w%���4�"�ܪs!��Id_<m����8����vs�:�jn��;�s�N葔����N��4&DF��u�q�����%xE��<gk��ZX�T�e֝���)�������W��_����Q����j�V�hV��9�qL�nEH��*�5�.�h��]�ԩ%=|�M���� qĐ�U�������RX�)�1⪻c�1�.}z�x�a9(LB�ԫ�wt�>X�젊݌�P\J5"�Z�"p|��uuv��S���Y���t��S���.�(��QU�:4���4W=urˢ�^��<�C�˞g��9�5�]����Hq�<� B��b&�B�"{�0�۽�zpcL����<SS�j˳Ř��,7r�H��aw2� �9+@���L�::V��DA
�c⃏30���\�X(�b��V�,Td������'S�%�t,i��w㲙&=oGγg���y1ӎe�г�`K��B��]�,�f`�'R�	]��U�C1���Q����{"����q�7�C��E:Uh�A�m���LU�)B�5"�|��|�������m���a�*�F�(���UT�<p�ry2��
�/�ц�T�P�c�G0�C����s�=TYWWuvP�<Y��f�	��w��-�q��m�Y}�kP��eZ�4h8(((���p��'t&�O>)��[O����c�����;�a��MW��%���1RM5jj`�@Bu�IN0I!�]Ė�m4���'@��$fM��Nyt�B�
�C�8"'�b3+SA]�v�|W�_����q��E''hS�9�WM\��YzԼ�6�h�{jz��˫��5g<�O�8L�&��-�r�g��a����`�3���I�j���FI$���ڟ�?D�b~���`I�����$!�(����)D$� �&_���.&t\o41PEgV`��$�H�I�C�JEHR*"�R���TE"�*K�,Hő�*"��*J�*J$��J,���J,�(�J=R2BQRE$QBQd�E�%BQd�EBQakXF�J(aE��X�3�*Qe(��*FE���T��b�(�F)Qb�E�,���Z,�Z�4�YE�YEJ-(��(��*FEQb�(�EJ-Qek��X��,Qe(�(�X���(�����eQE�Z,kY�:V�:�uX��,�XQb�Z,Ql2�d��,��,QJ(��Qb�R2Qb�(���(��Qb�(�#%(��(���QE�X��Ib�(�E�(���(�E(�I(��,QeQR�QE�,RK(�E�X��(�E�TQb�YE�,��YE�(��,��Qb�(��(��QG�0YI,��(��,��,QEQaau���X��(��Qb�(��)%�X��,��,��*QERKE�-(��(���(��X��,QeQe(�EE)%YE�,��QeE(�I,��*(�E�,�eJ��,TK	$bF	��FF$bFTKX��Qe(�E�,Qe$��TQe(��YE�,RKYE�,���T��,Q�2��e���E�X��b��E�бE�YR��J�T�Ib��-%(,�,T�K%,R�J��Q,R�,��K�R�,���Q,R�K%,R�*)b�)d��JX���)b���K%,R��)d��X��X���)b�J%�K%(���)T�K%,R�D�K�QK%,R��d��Dȥ�RQiib�K��d��Y)b�JU,R�))b�d��X���)d��U(���b�JX��Y(���X�X���,��K%,R�KK%,R��b�JX��RR�,��J�X���)d��T���)T�D�K%)ib����K%�iT�K�K%J%�Y)E,R�K�R�*�JH�J��R�,��K�R�,����)b�JX�)e,��D���X���*�K%2"$�A#"0F����*E��V*�UV*�"#�QF#"1�A�"#dF�����V*�X�R��S"0I0FȌ�#%X�"�J*�(�!)I�$�TIH���R%B�J��J��)�DX%"�)$��D�X�R)$�X�H��E�A�Y
"�R)"�Q�)	H�)!H�
DU��E�=��G }��1r��(M�c�	���b�,��(�F4PUITfz���O���ɽٿ>����(���k����3�>��~��~�׌�]��+K>�!�'ɿƒ���g��M�������o��oQ��������,)��R~���x�"���?�����?��_�K����9! ���bRDAhDD�Xb���'�'�#�������������Hh��)K�pO�����>?o���4|~>��6~@������P3�ğ���H��RWٖ�>j��Y)*/��'���?����߈�M_�Z�������u�����1���?���?���LDD򢅵�D)	?�@2�$�TD��d* *�����o�\�U�x?��?�.������o�'i�N��ER�UZ*��Г(!U �F_�?��P�߱��4/�?^�7�?��p�Ò�D�������?���#�?���?����EUD��6���������?�:�?��;�������h;��}R��鯬����C�d���� C毈��~�������<?����TO��@gW��O���_�!�<��_�?�0O� UTO��_�+�g�k��E]���2����8M���M$�(P��*��+_�HBBZim��.�8�NXH���������2�@����ID?�)�Mh?��������7���r��^	�� JP�3��I	����߱~�UTO��P��)?�?���?+����~o�Ε������*��}E}��i��������@�䈟��G�����G�~�<�UUD�E�~B��0 ����~�UTM���?M�������/�����?3������ZWI � 0����pI	��-�������R�/��'��_����?.�K?��_��y}�����i?��M~�����$j�����?����1���c���x�	�$W�`H~���#�J^	�G��МD�/���?4��*
L��H�c�~����t:O��T��L-@���)t����I�;�0�����C�д��s�Q��}��.�p�!� �$