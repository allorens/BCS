BZh91AY&SY�Ndۋ߀`q���#� ����bH��        ��am��P��S4��@�*R6kmJM) ���+Z�eZ5%H(U*JV�L�KYT���j6b�	&�󑡚��&���:�̕a��mj�a�-�ɦ�ؤ�J��ZfVֶ�h�1Qb�l+B�KJ���+,Ս�4���m��$�-M�|�����իMl�׀�F���k�	�&m-m�m��[*j�5��Sl�+mm��@����V�-V٪ѳc+J��Ĩ���D̥d�f� wVm�����    �絕V�a��j_G���z �2ص�*����kbY�ݣ����k��Z�Sl�:4�mUkc���jUUt�ڀ*���m�����t6ڭ����  s��A����J
S�9���*uF��{׵�SB�w T��7�@	wWJm�.������u�
(Phsr��i]}�R��`mm%�!VU�l��� �{|��:{��x �=���=� ��{��@�\@){t�Y`�4�z}���n� v�;ett���l*�5ew� ;�h����kT�ٶ*Q�  so@(�y�{�}�o�sJ�(=��������hi@mu]�J�Y�P*���������� :�i>�UP��+bԉ5�����  ������k���@z�7Z`:�wW�
U���А�	η�4�<�T=���t ��]A�ZP�K�Z��5���jI+h�m�o� 7w� }���v����=�z�)Zv�\ ���G�)C����z����W� ��  �3��/cCM��h/�j��!��Xfتđ���  svـ+��y�z�Z�n� �ƽ� t�r� h��� uq�^��� -=�� [�q�=�[l6Q���4�)f�  ,�� �p ��  �j� ���@Ю���j��]v ��ۆ��ػ�8@ѽ����Q�wkFҙCl3�]1-�6"|   3�|t �p ��� �0  {���� �Àנ=�p�\r� ��x �k���z��lж��4�U��P(֟    �w�P��;�  7vv��@1�  Z�� q�� �,� �� ������� Q�      �   L�)Jdi�i��Oh��E@&LL��&L&FO`��T�@      O5*R @    Oz�UThz� � 2   !)?R��Q�j1'��F�6�������'Bww�����/����_��<2>�[P����B�oϹ�������yL�� ���x+��J��AS��@_����QU�����	���g�������Y��?�����*#�EETW��U_ǧ�*����}	?��?�O�*
��������_�����̹��&`3	��fC2��̆d3a��f0��̎a3!��0f2��̦a3	�L�f0��̦ba3)��f2��̦e3	�L�fL�0��̎e3)�L�fG09��̦a3	�L�fS0���&d�3	�L��S09��&`s)�I��fS09��`s	�L��fS0���ds)�L�ff0��̦e3)�L�fs!0���ds�L�f2��̙�e3	�L�f2���`s!1�L�a��&a3	���S2��̙�e3!�L�fG0��̦e3)��0f2���e3)�L��̦a3�L�fS2���̹��&d3	�L��S2�d3	�L�f0��̆a3!6a3!�L�f2�̆d3!�d3�L�fC2��d3���f0���&`s�L�f	�09��&a3�L�fG29�̎e3	���09��r3+�\��29�3	�I�3 ��`&L�2���e3)�L�f0����as��fS09��Le3��f09��r���fG29�̦e�3	��f29��`s!2f09�̦`s#��fY��fS09��.ds	��fL�2���e3)�L�f0����.ds���0L�as �f \¦`dĄ9�0�AL�#�s
aQ̠��s($ȣ�s�aQ̨9�2��Qʩ�U3 �a�C2 ����s(e̠9�2�f��3(��S2�f �)�3"eA̢��0 �ALș�a�(��0"f ©�@s"&`� ��W0"L�dA���W2*fP\ʋ�As"eT̂9�S0d�s �d@3
&dA̠9�0�� ���3*(�`Ëe�
9�G0"�Q�f���0������0��̓&`s)���2���`s)�L��09��̦`s)���2���d33��fS2��̦`s�L�fS29���ds)�L��S2���`�3)���S09��a3)�L�ff\�fS0���&d3L&a΀���]_�Ѐ����7o����L�A
u#�㬋VZ�j�Ѩ�a{b�Wa���0S;��uYy��F�@R�t�SC�]
wgr��
j��Y�a�a)����%CJov���K�,��j��c6���ٱ>�\��"���oa�e�L�5�0规[וP�ӗo(X�L��e����dɺ.��)L��i]���LGw
؀��0�lf��5�����0�.�ͻ�֍��ّi��Ź�]视���[�4d����&k�	�ܪ!�s#��R	���x�q��Ն������\�"n�C�+�l�l!{2��c̖�z��E^f������{F�5B��dv�i.Q�Ʋ ��KX�ʽF�i6k�`A�6�[+h^�/s01��D�%7d��v���7!P��r�I7�i��a��{!˔��8���%� ���&�����6����k*�s,�t�e�8��r�N�p^�"���ǘ�	���t�$���[kM9�XR�%K3q�ڋR�Z��{��3Fg�����5��r����a��nيP�y����ج�8T6\�� n�N-���55^�oj��C*��5�/6����Ȩ6r��3+ �3bV�N����LF�J��y�nͼ��-a�i�ĔD�N������*o5��W�쨥�igibɇRP,-Y�fl50Ѳ�R���gC9C[�+cj� 2XY�hՍE��n�.5/[4��̩J��H"�wKT��U�w�m̦�cU�M��ݷ�Q2�L�U�2��u�,+v+@�@|�K��+x��y�q�O5:VNE�Ƿ�6^
���^�뤅�4��, Iң�LZ��`Ƿ��-��xj���2m��W��t�����C/�V��u�x^dQ8���pڹs{ WVX��a���8
�]�vN����3١[[zt�x/oj5�k�yD��l�i9eV9/65�ˊ�(a�Nٶ7w0]�0`��M���c(�n��f�J�%	��5P͈,͛�s.X�e^ހJ�����T���:r���ز14�Q1��+%��v[�5 ��ך(ɤB��SZ�)a�Y���B���2�Ń1�
��`�{�u��xृiT	7�g�^꽳[cN���H�Q�q3�hʊ� ����B��-l��y��p�aJ@��s	�W��,e��\uV̑��'V��>��T�+m/JQ&Q��@J|u�"=���9����l��tLۆ�U��hܦs.'N��Z��l�vޝ�U��r:Z�
Eԡv���r��7	¬j�,S,��:4�9�����vf�*#Pe��j|n�,��W��k+w�Y&��
K���bh���d���&KG=���X�[��n!���7(ĕ��M��U� �C1'���V�1x����#kcͳ�SW��I`Et�[f�=n���d$(��!��(PX�w[���e�2S��2�Ɩ�6�4 5���$���6 !B$�^�l�	���d˺VC��u��Z���� ��8l�4-��i֝��c �u�pM�!�!½�%��͌��GVf�ys.Vђ!���f���t쌷����jk�Ě�Iӏ���a��G<7�D��㽧6J���J�sGoM�G3+o̦�!&�$�
:��n�S���4���e�5A��75�`��RL`��GY�Ep�U׍�ҳ������&.e�p�5^�s�x�2M�P�2f�2,ՐǛ2҄L�*ؙ[��
)M��P_p=-�͕4ܥT�A�-����%���N;��lM	_�/��Mk}a*]��/9fg�Kb�5Z����{h�5��7^4�m3"nD#,����:�� �t�SM]�Kh�+��1fJM���A:��mC\?n���Q�M�q���#>=�SD̸]Jr�@#�^�R�2�y�on���xǏZ�;h��6�YP������K�2f^M���m<�6��àJ��*|N`h�0��`��q�mM�{�i�!R��ĭ�dXE�퍲��y7(e�%Vb9���6�l�X:`�o�����C���[K#�t�;�MKI<#dl��f+Z-��U�9H,s]��⚦�T�]��4E5�Cь��f����eԧ�&q�rƇ:�(%�����7�?�MF��з�jY�!�Nf\.�V��*¬��q��P�6��t���]�w��\̺
��Zu��{�l07)&�i�h�d�cԋ�Z�5�j^I��V�F�Ѝ�d�T��Dn��l�5WN[*�`F7�̘��rm�O(Ā�m�g)mD��Z5Q�Әu�M;����Å���m0�1z�^����gt�a7��������X&�3BǕ-��"��e`o�E��-�ǋ't[׶s0�D��/F�d���W���yKJ{w!���G6�F�]�����z�3Q$�)S�]0F���e<A0q+'5�޻[��,�
)�ki%��1����RU�:f<��gջ[�*ƪ�z�h��e^�dVu�m1W�j�w��-h�/��\�"{���@��4�[10�-�c.V�,E���JT���U�c\�e�$�%*��dYS6ݵd��Pе�o�.�����SAiAJt��\�ŋ-$��s����Ysڡ�*�,c*�<�0^1
�Lܸ3r�FQ$�x�����1�5%a��:e1^�j��1�iѨ�m5ȢZ
�&^���3(�Gmʒ�l�`�L�q�ř�v�*�L���08ƦFA�
��I���5VS��5{*T%��ܐ�+skr���4�MR�a�q��0eH�9n�W��as$Ɂ��6/b�<fF�V<'<j:��l�!ZJ
��ʒ�	蹃yyR��w�=��hOJ1�qfS�ܽ;����5�g	`��C�ј[٨�ö4+b�p3�b�If3g^o KY�#%��S%e��K"��ʇ
F]7d�K�N���:İ�Ӝ.�����o���<�����e�]��ۯ6�d�FQX�T�(M;? d��0 f)�@Y�U�2,�����WD���Mm��,��D3����]
��e�,�P�71�ߘKr��@�dq
J��@�\)_)�3i�T�E}����y�hX������ω%��l;�Ә�[r`cu��KZB�2���:�N�2�EYgd�[{ev�B����yt�����B��ךP��gaej&���f�ۆ�n ��Y0���n��C���ѫ~w��V��@��F�9�6�K�cص�a9K]��7L�!�n�l�����T�t�]}ְ�o�猲�Qښ(����w�z��`�z�Y�e��kl�S+`���0�^[�(Kh�%��Å$��ꌵJ���w�_A,Y��
���}D��xt#6*Ǘ�'L��'a�j��ȁU�r�6�������hinc�(a��`�v�:8�i���
�
�gKȬR�fU�i٬8����Nt`;�t`����Q�P^�`���j���^k�2��k���x2iTȭ(G0��f�h��4FkM�@4���U�(nV��D�\�*BR���&���ɡ�1K�j�=��t�m�L����;��Kx&�m�e¯>{!'e�x*�<7�k1�&zmX9Wp���Û,����r����;�V���ܛ%����[I�m���dwr5��B���17/7+�r�x,�-��æK���(���$���\g<é�m���Y���h����>W3���(YP7o`��mmH�Q�K��m���Z�KF�;����um=���"KU"	�WJ�̓�E�'h0��aSY�a4�IӘ#u1�⣘bd�����j�$9/qib�-�7�BpniʅG6�y5aӈT{ uyrR^aǱ��k@�k�"�{W2���$$:�ld���"�]ÀIu�k��u��-eKř �]�:d
���{e�BeC�9�����Ѐ0�m���moF����$o�V(��e��6�;�v��x���
c��f����Mb˩����A$\:�G���0\Wg H�*1�4SÃP4*;ܬ�ܵ�p���ú�dv�.�T�0*{�CzqRز�ј�aT%����O��)���W-U$˄5�X%����V��X��D��e�j��"��������bt�	�42�'yX��['�X�N�(c����t��K�m�.ƪ�Ln� ��^�3��rmM�+�*�%1o^����l�P�(�J�0E]>3i��%�ZgvV���P8��e#v.i�����ђih٥R�ڋŰ�n�l�7��sm����zɸ�"�d9��h���C6�~Z�&]�wV�K6E��N���I
p<�KD�djP�%ƚ1z�c&�e����Wt�.�]��q�Kv�J����k�,LN֌��ժeF��%�i����^�N&�S�2��c�:ef�-a�ʻ�wv(c#��b�zh^��)=�j	���fm*7�'W ��p%lkr�)zs!�gQ>2&k:~��N���>�\uV#U+)c�Z�"��6p��L;�`�ٔ�VᎬC�
�t���,�P˦(ڒ�w�,�z�V��Y��Hi/I�,�j�rK���O��0������Y��q��j���*�x$�Pnj
��uO/%� �����v'{��aۛ��a���/C�[����iJ�5J�pK#T7[7kۼ7�GF�I��Kv��+[���)7�3!�L7��j���T%Kln��&�����N��.V%�@�K�Y�l��+t��tf���T��1ov�!=RcXc���'م�%
w�`xN�!r��n�7u��F�T%o�(��b�ٍQ�'K �̆T�
��-mf
�!�V wE�C氬�٥ÈfA�
V+u���#-���VA$�"`V�Dl��&D֊h�0� -t���I�ޫl.70��{*�5;�N�-���Ӓl��-0�Z8%�0�0)�V1�$�՛����(;�������#5IH��ś�c(��6���ɰ��o]̳Z|��W[+��E�g[�]'�{e�w���1�J����PH�4cCW�ƛ�cP����K��ZP�3v���s)�)�u�7^�EiL'��R�Y�僞Ln �t�
%F���XK�a걌̤��{�G��ۄf�D+P�S�3m�.���f{v�h�틺�H�)vƑ�P�<#oT������ʴ-5����L�r�f{��1�n����QYYt�,
ѲI��
{Z�Y���yY�G�S���%����.�
*��X4:�n"����в�d�r�9&6�#8VL�!��J����T!OYÁjOr^
�]:i�@��'��BI���Z�!��%TW0ߍ4r��[��ե�����Hk]�xLv*޹�@�}�mި6��E��{�X�V��S0���U\�3��ֈa�{�ԡVƖ�hu��ݜ,2&�6������ݦ1Ь|U�$n���6�ZN��#�Zi��w�+0��^���Gv�v�r�R7��䆱
�]��] ��H�h�r��K�Ղv�����8t�H�i�d\!�z�[d���`��X�ɖ]��p �N���r-c2�L��Ec;��ŏslɘmơlQ���k�mT�V�8���s���Uګ���-a?��J�ݴx�O��:�%�X���
z�k]L��Q�)BKhP�4��E��!U�\9�쇚F[���6�֡�$Lxc�aM���&�f=�Y	:��`��&�Î�CWVp��F-��![Zf렜�:�އk<z@�BH��x�˱�3-�Wwa�a�'����%Ih�s	�����6t���	� �֧4I�{��61�\�f䰚��VA�X����ڡ�6��/5k��b�j����֋V�[R�۳"+S��u�@F �Yt�)̏/~x��+�%ȴܬ�w���sxQp�WkJR�^� 0��ku{LJ�jf̿�����8U�&\,C׺��0e���ɰ�R�e��4߈�{%[B�Q��|�D^nef�'t�Ө^��xӹ��Xv��VX�ob�&݊���ը@Y��U1Rܭ<��7�l��B0�N���W@��l��IZ�ױ[��kHM��n�Q�i%��|��Uh�W�\�Z���m�hS��w�8�)7��ͫT�{�v*�+�k��V��#�t\���&�N�b�&d�Dms:1LU�4��Øܼ"�^�ifL���Z`�
W�����1ZL���D�Ł�o�U�aX�H��h��"Ņᘙ"E�Su��d�ь��EɴHi'�HL  ��1��<Vup6.�c��� �uk'C�M�3lJ$g�0(y��PZ '�.Z��|^nT�: �#������J
�hЌ6���B��K.�!A�*�Ȁt@'���r�]� ���q�h��(;�C�L��T,#��p���"DZ٫(-�� �$*1m��)��!Z&�%"h{	R 3H��(�q��h{X?��IF��W4 ��m��8�xj	�Ap��r�6�"A��:�[#��.c82'����|KB�X�W*���BNӵ�0r��Z�L�i i*��ĳC

ֲ1
�g���@�\S?3�È��>�	��cW*��D^���P(E#p�'d�-*JE�a���4D)�$"7(�t�at	��^�E���0���5n�D�d�M�P��P�Jt,R ��GF��Yr5<`3��YL�YV^a�::F��q0F"�u}ê���#,("B��ly�yC�јBlhp\he���.�YN�Ab��[``���-�`A݉��Vc{��;=Q0[F3f)�����e��v�
K����cwCF����HF D�1³8$�˅ZM�
	�2�ʱ��\LEL��f�Yh{7�@�o9/<�O�M�k���H����ߛ�������}��3�|��������zq�w3�W�o[Sw�u�z�8/�]>lU��i5�sZ�,1��a"�Խ0t�u&��h%����=��O\�Rƚ��-�ecJ]d��i�	��y,�8���ڏD�/�9Zv�5q���R�^�f��t���&R춺�w"�,"�QB齌;���V�͒��yn���b��$�f��gS$[��Vͪ�$��+��6�vƱc��+�r�Xˍ��}E}��$y���!dQr��\	����:�3XX�tˍ�U��6��Y�}��篂8,�yR�V��#��[�R�{g^Dc��l�����eq|��Z$��~�N�.+���8�V�1����:����v�{5F=�<��ºT�mK�»3c(�vM���9]��Uz��J�ܒP�V(���[N�V�]W�3u�hm�(N��[�]F��/��'���ړ7569�&Ⱥyٕ�vGv�d5vb��֢�iF�f&�錽�v�D^1�E�v+K��C��7װ��ԡ"��f��?[+�!ӎ*��R0�7]�qat-��Y��}�]e!M����i��f�G�j�<{e��V�(��[�A�J�����:���5(��W����� '>�F�"9���-F!��n��Un��J�"�-��ͪլ�o�B0�X5zc��d�����S5۔�j��̉�ȺW�t�I�}*�Ce>`�3a9F��	j�;�O/ov,��1��M�%��&"�^d[1
5v6�N�7v/{f%�b�����HH��L�jҷ; d�`��j�u�m^��ٙG(v@��������U�u�fockfۖ�}�,�*-6�
���ʆ�n8��J��d�+�6VR���k�"��R���ش�{9Y���.��Ⱥ+�����]͎�><���H�ݎ),O"����Wr��R��ai+�7I��A[�VS��!/2$H�.�fo{ޮ�3��X"������c/���[��!�]a��+ݥ�K�D�6���������Xs%=E\����$JH�� -�&�[�[�);Yq��;I�v�>�٬�̬}p��?rUt2a��A�r	GLF^�C��c�D�A���Ķd�on��AÚ�c9&ڢn��뛱ͩ8����L�m�]����q`��v�(�T�a�k$t�s�v�����CI�"�w#�W]["V^O���U�8{��J]����N�\S��o˽� GT�C�#�F�ḊY��\w�gN��u"�qXdsu���mk���3���僵��B�vv'�4�׆��ٸ�ۺ�&V'Z���e��YV�:.:J��}n˳�+[���z��W5�6&*5�.7�v��뷋诋����s��a|�iB��Ɠ���9f���Ӥs#�,�N��<�.L���6��p;P����*M��z�
K���^�(3)��-vo��f���ڧ
\A�n�2�
x���Z��G�&��(�w����Y���γ�,��򭖻�e�������,Z�V��0ZR��U�P>�z5ڂҘV�ǍHo!�D�C�X��;�t2��p�0}����r*�`��I�����Sf\Y�����p�51�A6��s�k�{ƍ�]V��#F�ӹ���8���Έ`#3���9���1w%ԗ*�L@��0��Βk���Y����s�����;���nV�k�j��yX`�A�����Z*��N�ԓ�4���c%5ۙn�e�P<Ge�]�G�p�m�j%ΐmG{ia�-n�l�ϱ�Y�eN�;���vbj�gn���tͲ����r��t�i�3(�2�fqtƦ��l;*�BxuE�E_B�)��z{@4�D̀�s����^�}��;�u!S#���Wz,%]�iv�h��,ܷ���sC-�����'Ov�_Y+�cw�3�,�CիX�y%5��I}�s�ES�p�e�h�1ݵև6ְ�Y�(3eq*}�%��R��#� ����&�fZ���A0�ڜl�zUN���է�*��V��\��z���u�p�&����K��]�����/ X��U�X�7�O��f��|{k,�K��5k��B@MSϻ{�S-ò�v���&�\b�K�^���gQEc�8�f?C��� ���uT5�2Z�wo3s�����KS���%�2K嘕)R��m�t|�b�:�N�9��M�F� �Rs���%���)�U�;2�,-�Wd���(-�8:��y��T�u`H�ٛ�y���ԉ�|.*�e��$��W�"�0m�6q����t�CG��m�7K�9rU8���S��.W&M��g8Ns�A�YM0�e�O	{9-b�#��U˾�b�p.,�W<��}�;ζA�i�v
�;TO)�u�!��� qRu�ĥ��w"��:�/{M��l�-��z���C�T�,NVe3��+�4L⇑5��*ͰFٶ��ڸ�nb@E���ֻ���[G�k�d�-S-�,x�a'�MV:ڋ	�s���V����:sC�>�]�ƹݴ�VN�/1����ûת�c��4Y��\�ц�T��rr3�Q���Q��������
�5mڥ��.=��n;�W��}9����9ZvvWLl�z�������W0E�Ֆ��Q&�� e����+��W/v���j���^��Xua��Jz)��.�h�uA\�fc�p�f�9-�Cv�MoGy��3h�P\�h$�imqǥ��_@�CV�e]��ڻt�&n�8�@�̃A=�Ip6�˯V�MB�bnEz
P�0j�a�<RӶb�M����ąm�j�R:x���ٍ<�z4+X�ҏ>�5+�YO�=c��Ә��\E�[�rh��u���fݮO-�;Mʟ_	�-��YH*~�ޱ~�2=K�n��ȝUkq�u�`��ͤl�!6�]Ԛ2��K��a�;t�NHyw���k(*�yv�����K�Ю�U��x�ʆ�P�y4��+�LWlHU�w��l���ry4�:9�w:��y�9=��9��,U�5wn�[\w���srޑXa�d7��ݶ�.Q[�������¤�k�+\6�|[k9qv�Q7w�G/-��f�=�w�Z�տq�	��6�u��8�J��=K8�w�󮬸�X	���O)+�q�󭅁a6��3*]��7H)Ȫۼ+�^��r�P���$˝åDQ�k/:���]�^�Nm*9ޝ2�m���r��+����f\���ӊ櫩7��2���r�Z�=�],����EE��!Z4턫�ٔB:ygj��̎�Q�ƙ�7b���_k��$+�A;/��zFc烋�j-��F��m��s&�
��P�5ƭ?d�i�-�3|n+ܢ+Fi�N�|�02�gڴ�}C*k��5���fVI���a��N�nh�v�Vi-�E#q����K��c�|e8��G��{��.��k m��Ύa�:�BB�Wf��S5f����Ƶ|��ޚ��0Av�8+��x����L����.�JŘ�i��Kh����҈7����-�Vt\ ��^L/�̈́<�/ ���"T�N��7̌��)Ȓ;/o��v��c���e�x�0 ��9�M����'YJn��tv$I.�ӫ$��lݒ��V-%
ʹ���ֵ�M��i����MG������TZ�I�HV�c ����4F-�@Uܦh��z���-ؕ�vٛ����D�:b���1f��J �nU�CzL:����@�2w1�*=K�"�|Ou('I�n�;z�'lgn�=l:�smZ67x?[���u����.n-;�X%��oF�頢���k'+5 ����{oR��Ԡ�y��NW�[ )s�D��<���4ɛ�'^T��u�V�V��Sv��u�������V{\*q�J���Yy-�#�C��`��t����	�3�K��_0iغ�ǐɄ;�e6����wV�M�u���*(�nq�ۡ��N���8�z�dŁ������˥S:��@�[t9�Jٓ�okXB^����ʆ�&�MS8�
q�5z�V]&�b��>ׂ%�4�:oktm(�x�Z8�q�r#z^�u��5cY]bq���]���V�L�nR���H�R��\ n�wR�n�7��m��.��J
�6�o-�z&jM8ӻ�q��Vo&�Ĥ,p��RP���ъ��j��J��1u�,=>��_+7��ę�h����g0^m;ݥ���� �P��>g[q�`��Ga6��/.�K:hفy�v�nA``�&�z��:��ԧkڬru�
�2�r�l�ݫ&K��ѭ�}Eے��Um<7�V����5-��0���d9�Sx޴��c9��m���m-��~w��9�О����\��_йwu�9��h�u-��0�w
�ZH͜m=n�����G���B�db�3�:�zv��d,�<m�Vʼ�]�r}2��E���փϕٸ�ݪM��X��7��k���=}��WÍ���ϲ�0�}�3rd{{��*b������c�r����XC]��hw�΀��J�ؑw5��;�F�P��л�Z��+8�����v�z�1���֞3u�@�*{���K�+�5�x�S�=�	Y�e��Z�gϸ��x8^cNn�j܆'�RHn��+$�1h��X�������{�[
�C^.�2n�Y��q�8Պ�-�]ve��@���-E�&�	E�o������D)�clc�L-X8��p�*i��S��v�Be�ӎ,���
��:��o�JD�5u/)k��K)�y��!#yu9�RǊ�p�{J�i�j@�P�S���M�Mws��i���hrx��{ۼ,l��Ǥ�Э�jj^C�έOn�����M�`Ŭ�C0��ݚ����ct_��!"L���š�z��P�|�暢"�xͼ�Ԗ�/��Y"#�yj�ڛ��l���X풕��f �/���2��Ǖ���{Q��Վ�d�z�x�%��|F˨�h�"�ٰ)p;��1���~��r�0D2��X�����Ii���̵g�<�w<X�){t3��:��ab�=�ۭx����tk�uc��kz��AѾ��6�3,��噎l���s7´F[���+�0۽SE���ڬ�ԛ�0g�nZ:Yng^���ܩ�N�
�t�'��a�K�&����N<n�T;��S���M�}��G�1+���Gq������4�r:����H鷈2�"�]kz�1u9��{1u���q��< ��[6Y˾��fG�{4���r�Y�N$fk�5&$�ӓ8.d[Ø�޺�{%E��}Z*3�/;C�I)�l���90���vY���2%Nꞕ����Y�]����y��m�*�]��-�7�T͜z�$�!��6i��6\�܌��+�V�۵Yu���;eEF7��Z[|�؇b6�:�&e�
}�{��n
�ͫund��'BE�T�{���;B���hWZ��Vpv�&='�c���vI#�z틵��#�(���Ў�7&aCq���!��¦��hbq� _�u#ˉ�D�����:� ������z������Bͽ����EJ�N�kk�7�^Q�;�}�XΗ:,�˳f�F���(eUVVD��u��id.C�S����{[�.��}|U�����2��^�p�����Q���iu��;N���&tu��e�t�Z�**�J�%uY���鐊��N 1����v%��{�gZ�ar�C�>N�é�:0M}Ղ��s�J�em���p� a���=�:vR��%�����9_f�X�br]��Bv�S��5�+iQä�\���5�93�M���M$N���-g`J����YZCn�j�˖�5��6���J�3�_2kvP�::�v���&�\��%�z�Ṇk��Wt�Uٕ	ٸ��kD66�<�m�ڳR[��2G#&�nCSHf�晰�I������CBJ�d��W�6_6�'Z�|���;%I]ٳ:��t�,[ۊ�vu�TzN,c���%�5ni�h�.Ŭ�N4�$p���.�G]�j���sԧ�9ܽ���kM3��\%ά�|�|o[u�JQJ����$)d��sa:$�\M��e������a7�~�zE��KV+r�JZ�۬)3˧KN����!�9�j�$u%�P�q=�ߥٽ�;E�,�����]�l�d�VQ��W/9t;&���,���)%W�̔5d�9v`c�r�b)*P�-�(ow9��9PZ�QɁ��R�hE"�z�E����%X�).�ܜR@23%ʗt3_bss0�I$�I$�I$�I'{����{����z���0��'�g�<�o��(y��[H�ۼS��A�J��b���;�'���:~Hy��F���������I�By�/�����W�̆�����@��Ї�vh{!Jꏗ���Q�O��������S�o����#��K��\/��:�.�ᤥdx3������~�� �-ȯ�Oy�{(~sa}���<��9���J>G���?{ÿ�@E��g���PA>��(����_?����L���������C�����~���S��y�W�N>�e{r?5���ƾ�D��y^��4W9�g-����\���FCv�.'��ͥ������3z�fU�6��6rq]]�V�/ <��Gݓ2ޑɉu{6T�&��ݛ[��R��r���q$H9�+��_^�ȫ��(���l�T�A���c�����.��-����%����R�9�SY�Um;Y�Y��sC;�
#���8�I�@�8����ms�#�^�d'Y\+�P��J-7u�{�@����Hg�W�Hr�wF��V���1ww���AN!e�eS��JRug�r3��U3�R�;����W{�1Su�&�w>�ェ9X�>�5�ymJ]�Iv}w���<{���L5�&(�V��e�C�<��i}U��}dY�+AB�/7O�rF$����^�B#�:�u�����?�<Qt�WQ+���J�rK������m m��*x3���v�� )�����8�gw|���u���wmQPǓ�7���C7�5����3ay�$�x2�{CV��۰n	��g�Ѥ�<�]��[�آ���\Z��n�lWe�M)�p�ڕ٬g��T峮A����KW�oK]\؅�3����XMsa����s�ݞ�o.d#E��"��jvJ�>��⤪�U����b��q�t�:��\;.���<M(L�t���?�������ׯ^�~=z��ׯ^�z����랽z��ׯǯ^�z��ׯ_^�z���׮z��ׯ^��^�sׯ^�z��z��׏^�z�����z��ׯ^�^�^�z��ׯ_׬��ׯ^�z�=z�^�z��랽z����ׯ^�z��z�^�z����ׯ^=z���ǯ^�z����=x��^��z��ׯ^�z�랽z��ׯ�ׯ^�z��ׯ_�^�z��ׯ^�~=z��ǯ^�z����ׯ_�z���ׯ^�z���ׯ�^�z��Ρ�cyM�Zi����+m	�	���t���«_}5����#:���_k+kw���w�3JΊ��^F��3r���Q�"��uN�$W�٘_J�/xq.	�J�����)F++��Sy��{fRuB�׼�2�5�jl�*��i7�G�6wl�ȶ�״��X��R�T���ؙ����C�����̨�ѫ�ٸvd3d��bm����G*k,ػ�	
��]��x�kKW;�Օ{�`u���u�e����e�`�!&e��%іL}F�W7���]s��6R���.Ku�;q7+]W)MP���,�U��L͚�2J1��J��uǚ5��1[a-���Y�]��9]w��F���ז���������Z�fS�:N ��j*��Ε�9; |�D�ЮU׃�,uV-Wtw��eb�л�*�	��A�H���V�wł����6_ 2�t�ڕp����l[��+�:�O�pr������m��kFE�@�q��Q1�Dz��gw/�Hɪ�W��S�4WXڹ�7 �;"����Л�H*=ц��_
Q+��\/�qb�LՎ����*��r��]��ٖ�Gh!�8��J�8�5M�gFkbJ`��{f&��Z�����@C,���/�9�*�<5����e۩#�6���q�o�ם�%|p���z��Q��f�ҧ�W_����}����z��ׯ_ׯ^��ׯ^�z�=z��^�z������z��ׯ^�^�^�z��ׯ�׮z�����=z�=z�^�z������=z��ׯ�^�z���ׯ_�z���ׯ^�z��ׯ_�^�ׯ^�z�=z��ׯ^�|z��ׯ�^�sׯ^�z��z=z��ׯ^�^�ׯ^�_�=z��ׯ_�^�x��ׯ^�z�=z�^�z��ׯ��z��ׯ^��sׯ^�z��ׯG�^�z��ׯ^�g�^�z������z����ʽ��F��	�(����!���.���+�|�wn�Ys/$��p>�9�kL�^pV�n}X��6vM�
���[�^a#E����;Ws-�$����"� EY���g﫠:m_,z����n7��u�ԥM��M�-տ6es��[�re�QO�`�����5ڛ�Zo�Ь�a�x$��;�(i�[r���iZ/�"���gv)���+�b[rv�n�YRf�!�;r��V
6�;��,$bA��|[l��+�����Wvv#��K��I֮��L��+�}�0ٰ�u9�c��U^'�������9}fR;�̥x���}�RWX]�F�o]�ۧx�)�S�Q<fw%�sn�p�o�ϸ���f��D�_,�+7�l���˨M��f �u<�wp�l�K@y��.�oZ��l��j:�(�.^�a� <ZvJNnV6늫���Xk]
�*F��"K��:YWf�q��b�)�u��M$ �k�����wS���oVl�ԡopi�g���>vf�N
��Ws��+�du�^Br��m�沮�v���� ��I
R>V��ˁ�߾���f�8xZ��n�^��l�'���"^ol�ח�&�]��lu=זO#��p�@��md�r)q��YQx���l��*�;dްh��)�z�gn|p���킧v|�J�\�q���So�bx3�t,�[yj��R�f#��WV�
�\�r�j�H�kP��t��KD<����C$�Mʵeش�Vj�>�E�5}%�<��N��j]9�᳜
6�qWĮL�k�f�n��*Z��v9�
;��˧��v>�^gd�j��U.��˒/�LC��
��/�r�hN{���[���ޗ�nu������n:aQ���BK0�-�D�����1�OvJ�>��"�3;k�F���x�@��_[�+F ������������	*���q)��D�n�Tу�h'�宩.�Qᗲ�jn��EمIݷ��O]n�s��1�N���7�)�xy&M�X�t�P�-�VMUY`S{�9�5�)}N�:t��k��
�l�G�﫡�Uv�6�Z�+AA�������M3��:7�A����j�{-奙�.��hQ�`dWW�9E�א�O""�>X�1* ��lgu��.SZ���Jy��=�}ٸB޶��q��:6ZĂ6{ukJ	m^�3��v�vs�ڽ��FLpR̙���Ôm:B1��e�di`�W1<�2�t��U�?[���c�;8�����ݨQB�Gu�I_wt|&ɇ,����{����_h���7x�ր�0�����G.��t�D	��k}��/�[k6�S���C�f��+�9ռY�[n�o�P*�K�ͫ��7o�N]J�������J1�[ۭ����fQ�oWQ��o�(�ʝ�s��عu��-YX�2%#�w��ou}S��*�'�,-�T󖑛��˴�tĥ�:vU�j�ŌbmG]��Vƨݱy�2�[<P��}�9͒�#�U��E,���7S)
�o-MV�`�>��ެ�[!v�Bm�h��X��9b�yv�稖��f��O�MW,�u��X��`�N�[�g�t����8ngK��˨����Y:�!)-�Y��@�ⶉ�*�>��p"��6�F.�#=�eae#w.�Ã6�m�w���b�҈�M�4����ªY0ΐ�P�wM���������1��x�ǹ7L�2%[�Ukxo2٨f=�D^�m`�3[z���=�y�W�峀ݖә��*�1UVf� �3b�$pNõgwN��װnG�	N�1��4F&�;��+n�H/)L���t��$7{Z�הR�|ldڠ��^[8��>%�w\��
�'	�Q��0j{뙛R�\r���C3549��c���u�U��J���J��`d�V��F�������p���^��w�hA��Z2��X�x���G/Pdd����+YJ&K����K\�gXꗗ�M06F놃Pw��lF�ܕ��աZ��'L^�k�����,!�m��ܦY�k2���-�gw�����v��ʥ3wjA׉i��@��l��]۪��@ư�N����g-�$��SQׯZ���Y�C<��r��,��yT"2�-#lS�S��,f�T�����X���4�=W��N�z�<�.�u�R3i*_T��3E�W��؆VҬN��QΎ��A�ü�=��y�X�b��\9i�P�ҹo�3�^�jL�9�.���Z5
;"�.��2j�!��RfIE��uoe*s)�x�lͥA2�Մ��%���x��ٺ�m[�i���"y��0�+6�4�k�B��B�Q�\hWf����@�;�X����jU�k���I+�e��:�~���	U���a����h�[��Ц�c����m釦��m�oR�'XR���V�2�B'qJ(�Iǌ��ٙ�zV+��ʧ�0��w:��*�p�`����!��i?w�\S;�v0ep;H�.��@ؗl�WXmÎ�k3�!��/˖��X�K��]��Wr�"XEفF�g��0uC�0+��t P�u��ݨf" a���//V�w��& }}W�b�G�ڱJgpߧ���KSD�|�b��8����pq���bA`vIs�#g��Stv'b�n�$�40�z�h�Mj����rarj��f�����B��V�Z�.���p�t�;Y� ���N��5,���/��;[�C�O�e�1�~��DӺ����(�˳aw��o��v�{LًM�X�["M�dE<ǻԴU�Qٮ��kd�%��Y ���t�yPX/"�5���	W˃���d�J�@��%J�����ݛ;d�V�	1� Ι���Ug�G�iif)�1�J�a�� O^,��]�v5W����p��hgs( Ԓ��Ut3�_^j�`].5f��Er+c��5���OL��Ү���h�ִvڗ�M �;�s[]jb��-�Ŀ���h�y�*i�R5��>̺�X�G�֫��b��j!tY������Uj��2 "�3��U�s�:_�]i`��7q��
's)�X�#X��׹Y��ӭU��\6.14Ͳ�$>f	Df��j��󯱰��Y,�0L|��0�@0,�tИ�)ɦN�k^�t6��͖Nv���A�w�#���K�OA�"�u��/i�e��X��1,�q���u,w�'Q�i�9^�e�Î�a���k,�x(Ʀ��C]���Y����OF<�f�5��&J�Z~jS�.+��Ɨ:�nJ_l��9�\������{�Ȫs���NZ%*��)�!HD����+Q���"��d�����
{ڶ�Vu� #�Ms:c+P��TQ9���(q��32ɾ鮐���Wu�׹�2-snRӥ�-�os/n�I��N��d���aZ���7K�6��ݼLx��^�6�X\�f���XWհn��X��L�j�{�蒯�J��Z��D���c` 1�9�O-�n��-�yt{x�W{�&r0��c�s��f��5�
�ma��8��4�U�^x�V�]D��n������^��E,|\�������t�+N��v�l�%�"'��<Ց��z��k��P�m-��b�V����&�Ann�OmL��xPK��5Z�	���yƳ|�\�2�e�����7�:-ar ��N�K�+WJ[��O"����<�r9]�	���w�R|91�Vn,��mY�6_ϔXw�k���f̡{Өi��V��5�txކv�;cbXk�cu��T���Jg#ݔxI��6Z��e+#��X� W�r��Y�U�F��ˬB��Y2��`��z��$%���G7�q�8�o6�#/��(�-���g��-R\�u�ƒ����m�h����W9�t���Y�*��3!�e�^������j47��p9ۆ���E]{����X�����v�>��tȱ�M*Uy��Z�����猹w	��Ub�5��D��v���@�a݋=�T�Ldc�Y�c��)'u��fQZ�v����]���0Hc�W�����Z�&=�D��-�S���t�_C0iįY���G*��n��0�C�|j:����|Wwv��]Ρ��*��L]���J%:�Xj�7�$��;�(��Dax����9�޾|ə���C��Unq���k�U��uB��z�鼷v�ﯵ�D��A(�� �PV�ֺ�t�$F�U�8���������/aY��/3A�p7V�jڰ�[VL��Δǐe�����	rg(����*��lMQ���Q`:zM:!�)n^7���eK<*�A�˾��J�f���zF���M��ڠp�ǜ��:�����v�`��.�ᑱuL1�����N9S)p#a�,ˬ�NYΏ�Ir]Uf�2]�Wǈ6p6R���%�.�S�c���S�����l��!V�S���0��6��.�zvj�5�"�o[;Z)*{bXI�h	��v�*������k2)��_1��`�fh۠AYA��s�^"��5&Cᛵ�.�ZX3Ĥ��|�(�Rr���T�b�:����&��T2w�:!� �8�%�[R
F�yYX[�c\�a��/Em�&�x�Q�t^ �:OxKX-������#k��R��a�;нd7���e�2b<k,�5�+z��vS�;��c����*U��G�3v4�e"6؀l��g]�=a�z�b��0��8�L�R�f��b7�>b��"Go��Wv����B��DU��t����B���61��)��:����r�Km��^b`�����6�qgmj�J�]�d�3�^�X��_;F�ؙ�t�7𨳧M�N�i)t�n��ܺ#�0�cʻ�I,	XR�� L����G`|�x�2��1Ѹ�
�f��}Ys#t_MR���89T�L��/	HՊ�H�X⣺��>ٜm<c�Ks��39�l��Ct���r����@�8���9sVIcqwS=�ӢQ�F�=3I�(آ�w_}����@����G-歔#�0R�%���du�]�"V�W8d�<&��씫�0�w�}w�nH$DU�jj�������g�R��˛�ٺ����U�8(_b|$]i�wV�<�<^�ʪ��d��֙Ν������]�險8���v�NQ��E�cq�[�����`�hrޮ=5�ԑ��P�zN��80T�r����?��������{�������w���5�������5�������9y�p�4jD�Dƣd��В?�l�T�ҍ�!�Tl#HQ,8QJh�h&�1�a$���>��)�)�l6�	B�DQ
1�Fm4�p4"i��Q6TD�27,�T_��0I�c��q�ԅ�?ьM �d"m- B��vN��":q��,H��Q��-S��TI��L�d\�"�3��E�a
=���Z(_*:;��g��K�:�m:�A 5�/��%5*֐���i8��`�,�ȉҔAfduj��(s�K���k5�'>���.��A���E�&�o����5���r��ą2������,��̑���l��̆�U�)��+��ԛ�ep8��a��¨ԫ����|�u}����KQvmX�mr��Θ5��l]�쮖+ʚ'E�������V�U��V��Y9�M�+L[R+snj�9Λ�U��ش:!�Y�%�K13#�e�@7���-/��q�"���ק�bF�'Te�[6J�R�H�c�"�w	�jW'D�R
h��֫z��\��͔��PD��Sg"t�2�h}[���
�O�X�K��c�r/H{����{�&;�J�6kY뢢չ���)��.C Ι�GE(��)v�=�3�����B9���8�h��,��y�Y��{B��.�����fp�V ���MT�0v��NK鵔�r�.��'�(��`
�L᫠�]n��#he@�=��f��5�6^[��}���٧}���,���ݞa����Y�f�U�#�� �蚷��N��v���Qf���;v��˩�R�[΋�,,B�Zn뜂���%�	�}N�E������<�lW	���:�	F�)�NcL�b1��h���-|�D8�!��LD��C$N�����8b&�j�n1'F�x�#�
QG!,�CD`��a������(��XJ)䡎,H�9""�0��B�*|�A�0�
j��D�N�(�'�b@�3�3�FK!6R"C�-������BD�,H.KB��(4�B�f�"��D6`Q8��T �K�����$��B�e��j"QHB�i�� ��T�E"�r�y�~J�p�PD�ߘfEp�A(mB�%�`2�q"a$[`����[�̍�L�(�J$Ӂ�0�m���KLD��d:a$�%ፔ�d��0B*B1d����<�+�1t��4ƴS�LDCE%DL�34U5T�� �F?}�
���Q���_��������ׯ^�}}}}}}z������тj�!���Z�`��cELT�9Õw�.⪣ͨ*�e9�/�x����ׯ���ׯ^�}}}}}}z�����Q�E��4S4�|��h�iּ&�9i* ֩'X�k[D1QU��Qr3Z
�����17�<���O����pX��(bh�*)�X��MkI������P�a��<�.m�" ����E:uQEv�p�tb�1$S��Vن��׶
�����*�ڢ�"��*��sh"�+F�����c1U����5r��r5Tz%���E��\�T:�DKW#3��*��N�ՌT�sX?��-Sr6(��9�-\��ت�7�xp�j�:(�E[���`�gѨ���h�V7ˇ�51d���cT"��uEL�"u�r�kb���j��j؊F��m��>x�j�X��c�T�-B�ш5�Lsf-��-�U��)5�p��{ϗ�Z<��<��F��+e�X���4�4hH(!�BQ�&�0��z(�	�Q!��p �Q5D1<[Mw�~`�~�塖jN��.+Nd;��-|�_pAVJ�S�%)����e�bޤmc�5��Nc��ooV�ĩ3Ņ!�!�KI�&H�-��$3�D�H�$�'�@�!�x��ߤ�&A�҈G�����B�"��a��JzH�L�������{��eۭ�x�2�`��KKH�@mB$��NO9�ڢ�=����^��g�4E�~���A�o{2߱>�����O|�����9+���ޓBO[��np\Ӎ鍖4l������W�WfHw�^����@l#��m�$�c�9l�s�f�{6��=��~����Qc����;'�J�Qr����{���`�{=���or�ȹf��a����uy��[>j�2d�N��<�.Z��u5eo��������%<�����s�g�zXc��l�� ���,\x��>�ߊ���OA��������=����C_��!���Y`��n��C�=������û�wF���W�sO�|٪���j��M]J�o����.k�ȲxgPn,%�`I���=F��'�N�3F�aw�5���6�CD���NV�y�P,�C��?�Ț���A���؛sшc�����yR*��]�íSQ�/K�w���a��/m�NR�K۠��֍�/Q$��H�mz���d�U�J�4�U����Sj�^
�G��&�/���*]��!}��1���h9l'�S��v�P��z�����1�h訝��"���ū��~�����Ž*&��D��j�:f��Xِװ�~�{�^s�}���X�X_���}+��ȫgW����^��N���y���4�;��]�͢¹�i"N8Y����pr�9/�u�ƈ��W�%tS0n�K!G�9'�՛�qv|�d͢�6x����vV�����8)`'g�KOO@� �0���9�����#(_�n�_��jd���>S��~�q�&�{�6�:}�c����c�q�[�qs/x��<����y�sV�C���FoPPT�T�2�O��������C�>�����2�6���y'mȣכ:F<�rM6Uh�R�)ݶ�F�ֳY��CXL>�i:^&���i�`s$�ܞ�o��m�y��θ�$c3^���w�;MG7yژi�f���~&�n����=>ݳ�]-m��,��|��_��v�8r�B�0X����y�sK5���ЏES��aw[پ��ܾ��.�)! ��t�=�&As��kN�����7����6���WS���.�*�dt�Gh$5��V��$�4pĶ���y����s*��]�c�;|Va>>>>8�~���vMel���F�4���_A����lH�P(��E�3�+�y.v���M���G���z`���u�ӷ��u�p�I��'u��}i��.�3�}[���o�˅3��f�9�Qk�T��}������Ly�&i���k׫0����O���·��s��s~F%���iƼ����z+6;q{�������=��=__ʝ����w�R^��z�uy�����CjϷ�kk��x	�S�U�}Pի�N�lk&PV���ӕ:Q�I���/o�R�}�ړf���r\�:#�=2��v��o/\�u�n��^�C<������rS�3�Q�/�|����RK�NH�&n�^������n�G��EF�e�$`�"��mO�p���}��ʛ%�d�ҵ[��W�hH�ܩ6�Y�[%���I��3���p���Fǭ�B%֮��Fb�e��&��t�(1���6���P�ۮ�kG\��;���1��V�㻳|6�uE��ّ.2�t
)-��=pTl��U��b���*����[4��;*�qkv.�s����>��u��o7�ȗ����Bu{x��$�����l�/�]z�r�d��.���\&���xc��n��N���n�y�wƙ���yQg_)6���g������h���z�xV������K�&����l5�����q�o����[�+!��Nh��͂xooo��	$��;+�j܍�=%E7�z�]}t�vP��}V��W�N���$�Oi�	��
�^�r��I?V�~o^ջy��R��S}�絓�����ܞ7H�������S��K�������̺O*������1xZ���t��糯��p�I�q���I^����]��_r(p�VD��t�i�r��1�Ff�o��y�*�鐏kϣ+Y�yT��pX��<�:��F�����O�m�_d����C�?IX��TfV��rz���g8���5�e�k�0A��o;�w0C	%���k�q�W��A[聺�٫��Џ���V����M��T�����S�곝�enK/���9�1�2�V�>b�u%ٍ��J��C�y�	2�N�:0>ˁLy�����t2vF�]n���q8�f]_�
� m��*0w L&n�a�kkrۆr�&{��R���i�_KɲSX�<�u���~ٝ��:��
�L`d1����`׃��L��˖Q>w���Z�٠��׻ʤ��uTU��8Dڥ]Pg��Oy�c�p)-�\��م�u�{�f$Wp�і��j��˛,��sP&����n
��M�c5I��Ջ>�C��߾��y�1U%�ފ�<sDگ��o=w3�����D+sެ����A���L���B]v�v[�U�u�G��z�8M�MC�1�j���(�ÓjT��z����D6R�f����OC�>�9xIfA�NY��ދ�>����Q{Ƴ����tu�N�q������M�=��I�d6V�g�T�q���#��l��.���g��G	��,���v�h'��q�|��=!���;CQ.�A��oƇ��Ѻ���x�#�s*T�z������W�њ��D
�f¯��k!0�=�<n��R�{'w:�&������څ6[�WH��h
�\��L���Ɗ=wq���+�.c�Xs��O�seN�m��0�s��.���x����_�Z|��%~�<���7i��l��@�����]�q�pᜆ��u�h��z�u���b{k�t��u��z$�� ��~��&ް:u^�_i�����"���E����{)���K�9ىm-��'H����K;�h��I��_^�%���m��=UMӞn�<F� �y�T	������5F��yT�v���!�.�̪��+��VrI꺱�[aіN�����^��*����tI�>�_}�_��<7$wGz|�+�Cu�7�ޖ�A}a�k�p4m8���4˶��fm�!Hl^[�������:��皋e���s��Pd1m�mOM��ǘv��sRk3"���{ܪ����J�K�5�W9�U�%4wQ9���]V��tX9a���� NT>���%}�3}��e,���c�F��o)�i�/�X�S��:�!U��������~��{�/7��/O]��e5�[��m��x�z�m!�i��^s��Z�k3���D}�z��$� ����0+��>��� *>���S�ֱ�n�I>3���B�M��2��x\�U�M��s/�iӳ�)zuAS�_��l���'>_��]��%�� �"Q �l������<���W��Yܽ���+���e�`��ܞ��=������;[�c]����7��ُ�۹�c4�*v{'y.�����5�ZV�W�70� �/�n���3�	&�>^�t�u����闒f鯢��X�us�>�
/����{�o�����5�^ԝ6��h�ʞ����l��'�;Z��o��Fx;}��a�4�^Qq�7���&��5l�ק��^z$ى;����W;�|-}㭃p[��^�Ћ���'�_f枧��<J����_��_�3��y�8�V5����{M�+��Ƨ�z�s�4��4��i�4���a��qk�K�r�U���nr:��G�{�B)��#���|�5�����ʝ�J���o|Y�N���&����ׇ�7>/�;�}�o	�%5�#��w�ի���,xt��X��-Υmc<qT9��3�r�<��s�ZC�e
&�����29�y��aU�cM���>�� �pWS)��}N�x�����0�&�+�q;�ٴ%"w^fˊu.��Vw�Ol���ȀJl9وN�-.�7�����x�r[��6=����8�J�s�&�M�˙��吝�KW��+�g7o��e�r�_P�|hd����{a��Q��)�}lU��E�Ѳ��yY�~��{V��fd0]����spp�K�#���v�Û���9^�"~U$W��q��=�RJ�������}�����E37��������A�F:A=m>��U�U��{~:+YU�ܔ �F+�'7"�x}�qQ�>���@wI5�&d�0v��^�ǫ����#y`{8����/QqWuw��$A�����'Ct$����A�-��V���!����o�F�'�.�����8�����sϷ��x����
~#/�݉����;�d���:ہ�op��<'5�������%�Ob�x������;�{����lZ���>�{��D�Wǎ��@�|�w��f�虵�t���]�Fl{��|ۓ�b�`�����a��V^޻�(��)m*�����X�}di'�����;D�;u�޼����ҬW��d�U�Ȱ�Һ��"����X�AF����\c�'oӻ����|�||T{���7�I�ĩW�Řk���[m�
�����
���˜�{������D3=u�?�m�yu�~���ը���-��/��{��;'���74���U�ҵ�]
UN�{��ٖ}����ש�f�� �{/h���Qѧ,�TgX~�Pm�E�_��/sxK��~��<�p�����>k�������;D�L/<y�B5Y�۠�Oyw�nN��q�V�C9���7����{}��ޝk�ަ�5�=~�v��)��%G����e��St��}^�T4�W�a�{^��r�89{sLvMT�H�4$a$t�_`�4�����,�x���u���r�Ʃ�f�U���i<k<E<"���S�֭�WQ�@���S��eX��,�Q����Iʾ#��v O`�W�~���q{:�̥Ƿ�#�a�߽^X���zI˘ɷ�r��L�&LzD�`,��b�E�`�r�;^��|=�t��Fy���c�+�9�^�y����.�����	Mw4lɗ�]��q��<�5M�2ۃ5#��ܢ�8�ov���۳�o,Y֭�}JN:[�r�]�[qv�V-�U�%�$i������M	��Z��h�i�H��y���]ew�S6�ڕ!���$��~��l���ĿP���~́}�K����Tz�^�{��ow%��Vf�#%�zZ�a��@מH$�S�ďjYS����/k�{gG�:d::ߏK�,�����I�c^z|s�dv�y�}��p�ϗ�uw��q�5�Y��{ǯ��}�o菤�������e��4��h�䟼ш�S�WT��U�ߤ�ۓ�Y��8���=�͞/�֣+�v����ܠ�|M��]
5�^�\L�a����H����׽&�����2��v��c���6�������ө��ӭ���3�K�X���g���賑�8[�wYwvѝ���}�G���>4"�WZ�^h=x��/��csCȮ��]��mAg'�IMl����̧�>�P*�:�X�ў����s�g[��Z��FI��D\��ZrN7{�&���]w���\�B�����b�Ҿɠ�V�Qeѫ��.���=%��T̘Q%Ǖ��Y��i����ݑ2�N-$nwWA0��95�S���9ȣ;����,�y�-�*$�'N}w	lX6 �V	X�3�c����G4��1���\��6�>Yy�M���t,9��Wt�OQvu��eAXVc7�Z-$��f�DJMїٳ����j6���D� %ɺX@:n��	oA1]\�;�8(�\�Ul��w�B'Z�gt���� {c����V�9�c�v��1F���:��;�<�����YFd���w�,47�+�;��y����$�\Vhy��e�5`�F���bј5�M��V=}#�q3����+7�lme	x&��n4#7�j��<��N�xJ��I��8�ka�Et�ze���K[co5nm���yQ�l�!���ܛ��y�f�b� V��@���#��Z�������Ûr"�����eU��n40�"]B���L�D�<�<r��`ޚ)Ryi+����)³.P���$�12-v���w��hv��
��L�@׬��]��;,��	��a�Q(Φ��"V�ù��[-@��k��]\U$��a�#
B����$�^X�=)��讀.m-ﮖL�8__Z���R�`��-�� ���S��i[�%F��[���H�^6��vP#��S�UL�E�]4�Wf�Q�M��FA�`�::n�>[��؀�;�8��>���N�mp�Gg�ճQ�.��������{��j.sdu�wX�t_I�)��ܠ�ha�	��aiפ��(���Q��Zub���t&�<�Aa*:��g_��6<*�9e�>�{a�Ԗ�KN=��<��X�}����4�Dyj���=�9;��k:���ݰT�Qʈ��a�S��%ݜ��x�Y�]�$nӜ@"��st������A�;#G%#�	�Ɛ�W[E�ɪ�6�m��$��x��4�krO�f�{)n���FEy�*á��WЎ�#�z������̇�.�x��.gr��O�r��\�wwZ@�R����*Z,%)ɀ�:�^v��+-�2���n��c��cU]f���F9ι)F���oz�+�3�2)�K��Y}����Ź�˾�r���
�1��S���Ϻ����R
�E㸓Y�pl����}�,��ȅt^��ܰ^7��nٛ���Y�_}�pl�<��3�b14
��q#��<�)|���WM�Ԣj�?6m�[�����E�#�t��N�rs��$����.�z�nX��ie0sqtr�u���2+�Ӟ����M����3��ƟK"0�٥sP�x�\4���'�$����<�BS�77�Z)q�v�}�7�� ����^��(�6ۜ1\Yն����ٌ��h��.H��Ӣ��V��rgE���
-�$�-��^mx���RXح�Ym?^>?�^�_����ׯ^�>>>>=z����������Wtsj�.5VX����qh���DUGgZ.q�
��hl64Xph��Æ�4r&g���������~�Y��~�__�z�����ٓ,QTh�TIvۜ"i�����/)���X&�b�9�kW�rh�m���.�
���i��/��IT|���
 ���)9��r>���b�ت���"����6�5�j"����RTUZpMG�������nl�Z�%T{�r�E�1ʨj��#TQ�U�Μ�I��EUQDTME12@Ak1U�խy|�AD�1ULY�jx,gmT�y�Q��"=��AM�Umة(�}�sELPT�m��*�+�c�|�Mr1QT�5|�Ir�O��j����ETP^�/2 �@$�G�$�I6B�ѷ��E-���R[+��D��2��k�\'Z�d6tH���*=���Y�s�=�X���ıL��J�~�>χ��������F�����v�	|NVu�ͬa�侎- ��GNŴS��"��� �s*1�gj��s5���ʭ���:��5�0[�({d��.[ѽ�ٹ�&�%]x!��}�i��)i ����/%����:���xdKG���x�K����r޿K�9�/��T�a��Y����O�ս�W(j���۫���7$:�d�z��Ɠ`ȧx��������1�W/>�g)���E[�Ds\��uid�G<Ćx�6��3Z�'�P�tx���/Y�z�$�����������t|W�#������X�~��f?w!꜋e����O��Ji�%)��Ga�^�d�'�2���>9��^�Le�Qu�V���Ї���AM��8�]O�1�C'$r�M�J�[ ���k{�]�:<�k��S�^f��<࿁e�͵0�t��`��.���4��s��n�F��a�/e����M��{�3;�~����R ~N���=b ���L! &�7M�i�|��E�����y�?#�R	�E^��G�3D�j�����@�\?cE�R(֟C�G8���O@�^��y��0�������}���Ɇi��r�X�v��`UT���"�eqA|w�����]�|�$��b�Z�*n��ŋ=���F�x{�T���bG\��*_^p-ڕ
P5/�c����>������#'z5�5T�||�?����(��q���ܨ���?8��契bc�.�����#�W�'AG�����-��n�u4D[ F�����t�<��y���J��2zW�S���|��ۜ��.V�6��e�+�Y�H!��ghZ���2[��̵�a����U�������:�G��~e�ؾ�K�ѽhy���H�>���.��#��}��I?�LbXi"m5� �
r�P/a�\aR��,�T^WiQ����ѡ坨��͹�ġ�A����hM^�.�=0��1n���QL(�J6rsv���ՁW����M��&8 ������:���6�ں�CvIv
}��)���p���S�����6��^�y���|�#V0~b|iQ�����u�{�[�s��Y�q���S�L ��
o\�CW�3�����U�-�<���ô��մ���x�;a��FS�������P�Î�22a�׆�x�ځ,h$k���F5���s^�΂�,�!цȊv�R��������%�)�O#�ZE�&���A����^%B��T��W����\2��G��1Am��iamgmesXvl���dʴ�s_|n�+L%_�������sp�*�)T�PY{I���@�>P�/��^�M���]��N��]^Ԣ@֘�I4"C�ۻ��m]˶(|��c��L�5*�wj��U,�m��=������xk�?�%�ߐ][Q,�ݯ��I�vFr��$8��<�����{��_��{��_ޑ��@��� _I`9��$�^�IP�
R
:M��cm`ncH�ɣ8xvk=X��Y�h����@ĳ�O�`�C-�����K��R�ɽ�s1WVko��p�uN 
��蝲��qt1i�n?L��,>�ȃ���
>{b� �ٍ~���h�?V�G���u�+�q��yފc�S��-@.O#��/�K��V���~�P�|���B��W^]��ŀ�GC8l�m�R�W��U�=��(�XH���#�%8�#FC�Ƞ����sR��K:�Y�h���w6�y���E<41�"�9��.�*�xR��~=_������B����!�w�OX�r����p�C������,B`kf�K\�G�����pr^��U�0j�X=��Pxܖ�;G-j���=mB<�}�h�_ό�?/�ٛ�XkP�rT3�<��5x�L3==�ì²��ə�A^���B�(_䲹�U��t q#����Zo�~��ߗ�7@��s��v�øxv�r+���j��0��I�u��O��Np�Ay�>d�/��n�)���naΆk7����r�&r�tw'3�je$�G��7gZf^i��8��-�_���b<��M/%kX�n���������u���b׵�j���;"��%[S4e� �`�ʧ���AK3�n-���-Y���#�Z2������LyRt���~�Dz=�y�_�nRC����8^{��PnF��Dl�U�V�Ʒ}!�)ײ�~�X��d���_E�o	����䇷_��Υ�=5,���&yk�!�[�W!
�y��m�P1p�*ϴB)eD��~�=�ۻg��;��6
2�ܾ0�몆�q�d-{�A�WB��҃����1��/�.kjD���s7���Dz����h����È���VUK�Cc���%�&W�P��2���O�f�Cәs�vw_iᥩ��OM�?��ʘ	Hf>!�w�x����`8�oa��*�+&�[�G��k�?/j��q�����2:f-�.>��W�bN,��I��!<������J�fsS�u�q/���	��X�%���9�
cI*����Wq���j�?1x�`|G�L���b*��d+�؝��3�䔉o*��w��酣R���<S��R�}��k�C���[�Ko�����n=e�%�J"<�0�F��p[��f�wl�q;f@�rr-?2Ng�V���A8�p&fz6l�x�֞��W!�wPa��`�O�F�T���FS��K(]�Uz#�x�~��H$za�K��\�Y�h���l�\�G�_
��c�G ������Y-�������wݧ�{\��\���f�23UL榬���C�	���%X�68$���כ�<���`�݆W4n�)S��t��L��-e���n}@'�صuBU��y������Ǽ_w�߲b��1ݛ$[[[�۰��
��0e��&%�Pڢ��+MkxP'�k��k��=Z���Cُ��N�7��xn�lOtØ_~W掯�jy-�B��^6����D<��d�n�C�3�g�{C8׫��r9���1oQ{�y�5����,��8&���*��w�����/8J%�Y�2�������>������zK�"m�D[���~�y����NN���[��C����˅蝞.�/x�r��ٳ�!��%�qh�"x�v�_E��b*�m��p��̸��ե�ySS:"KN�d�!�Kսݡ�9���4/��4U�B��%�;�S���e1���/����؇�|b�}�b��Ň����7�%/���ض��*f����ͮ��y1�79U��C�����[�9a����R)���8���|�����q�E�9���
3m�1�v�C�E���N1^N�-V��xF-�4��{����|w� �c{C�	xz�nl}�ƨ염���H��\�@��,(bY��y52�)Rk�Ds{��t��� ���.�q)��+��f��}t]�7�wV��z`���I5�m-��W��oR-�3���|5R�	,^<�J�f���,��̬�2患������Iө�%:r��m�n��|�bn:�Q3@KSđ��ҹN�]r�ܬ��և��~�߼��������vJǂ�;m�G��Q,�28_B���8�%9��E1�������>Eè;l�>R�[��wo�v=h��4����G������������7�O���Oo��n�F��,9��LI�h53����y��D}�d3{��I��1�}�1��~��k�xg䯐�3>��.I�NQT�q��4��Ǝ�#ۮ1�̼�\lP��3L$��h�X(��R���LKu��1`/N�^u��+��)�5@C��/a��e�~���bC���j�jd.� �~q~i�J�D�M�s�Te7���G�*;*�F
}cMz��} �Ky���N�ۃa�?�~a!���5�T���x���^3�Ds��D�C���Y�2[è�k,{'��º�5U�z/��9�A��v4f,��SD�̼��3�zCs9M̡�ap(K�>n�ғ�^Nf�W����y�h�-�w�I�]=[v.�m��=MA�/K�;z�k;~�|�"ak��n׃k�u{�& �����Z����װb ���w��������Xw��5KO���_W�:-qM}���7~�y���l"��"��wgY6XXi�瘪�{�ITXw���� f��sG�;����Jp��$������T�0*��UX>�d6���ʻ�ۙ}�	Q�9��U6vm�r��s������r�Ov�.����1��v�q��x���������xxE���-�*T�{�WW��*��\�lROY1�araQ�U���k�ޖwo�t�hd�za��~lO^7�I=���	��ğmY��t���N���{���4dVrC�_Y-�A�*��ԕ�A#:�C6q��gO�.�,w� �Ԋ<(��Z�>�����{�Ǩz�[��� �����O�~�7�U��#6�_m�@z�-�`����V�q�-��ٜ ����PD�S�S��4��Z�2C|�'W�W�+�0���'A��$C鵺m�vc�0����~o��M�EЕ�nv���})���Й'�9�f4��Vh[yk)�|qrc)]^iڝ�̇�_)���{�ǅ�]0珄��L}�!���W�},Z����lr�����	k"�yfG�57l��V�>�3��μ�"��a��h���#�(-g�YZ{����0`��Rw�vK�@Zb�?��N���c-/�D�������f���A����!�m��s�ouu)����X9� �&D��z����7�r��	H� �� �|��{r|���ڤ�Hp�O�JCF�!�[@���%�?W��o�8��RX,��ҩ�7��i�r�ῴ�9��oX5U���Kd�4~�5��)i*|����!����K�9N��ьD���S�G�4o-V(�1����;5SV�sf\�D��*KW�ݸH�L!�)�9OT�7�U��\7��P�K4t䳺d�꣗��
w8c9sG��}���<z=�  �ZR"i[�!���DƦ�H�4-[� �-б�~�J��nn3cj�t�ͨz�: |-XK�X!�������N|�7ffܖ׭�Ò~�׾��/��n|�WE���Cӵ���}P�k�hm��>Uߘ
��~"�5?
a?h��덙'T7e�Hb���ۮ]���5YD���-��*$�a��虗iD[�{�[,y�h�����<[��/�^vۙo,�_r�z����z9巒�v/"�������F_|����+�m���Cc���j�KufݔF�C�󇬃��퇱��ۑ�7���P�p ��
��B��[�:l鋇F����t��C6s���C�x�;�΂XF�\�b�k�p._z��[J�!k��0�]
7)Y�43�}N[���n(z��	��r}�5Q\7��04  �����ʨu��Bl�	��%�^0��M�[d�m���O?���v1��[��2�����q%�B�y�CحS��Ӣ�9� LJ{�t��pE�/7D��uy���	�����l�={_q���-��$8���>Tǁ	��p����S(k��4Ǣ�r1��j���iw_6��Ov,�B̕�+����"���E�}v��l����Y��-��{��a���xo|n�K�(�ޠ�32���zR��W�.i|��F�8lU�Å�!�J�X]�U��u�ӿ�{�~�����????{����ܙC�%�z���>#��Tkڢ
t����<S��b��7��澴��de����oV7g*�=�'��!�R'������E�xXF�\T?}��[TC� ���Ï�dz�fOh9�z��L�C!�����&4&n�;�T?���s�i��rĮ�0(�t�t����7g!�an�	�rC�_���=�.�S���?M A����L��K�n�Q����普٨���oT+s���=���</�1�dӼn@p���:�ã��Z�^����%���	�a���J6�,7<���y�\dϮai�H�~���=��C���}^�"�/����"�ȇmt�O�ٶ��f3�\����{���#�W��'[�>ˁy�z��Y�i��cF,3��� v� _��������PW]��vI��y�R�H��l����~/��H��D�Ǩ��b�l@߃�@�>
փ��ލ�sJ[���}���5T����%����#6��4���qhO�p�PO�Ͷ�xK�5��<W�d\�^Ȗx����PCb���'>�
�ǻ��������,���k��_%���~��fd��5�"�ڝ|E���dv:�ց��8���`���?5@��Mv��6%Ցk6��gD!3b�������5b)Fq5R�Q�{2^�g8�	�U�:7�V����?] ��9��(�������;����� W��y������{����ݍ:r�=x��*+��y�}�,�bKI
>>K��K�9��,˒�lL�Z�=�(��W�4d!���ڗM��5'k���6q={��W�|)���������1��|n�4�;Q����\���<ssa0CV��y4#�A��z��[�z���zPP*@����T�)�L?J/�wot7!�a�YHܧ�j��`�ʟ�Ji��[���&v#�ם)�
J��CP{����EUf4�9f��^y�C���B}&z9�S���bS��S�ʓ[�Z�OF�������z�����yoCR���ڽ��j`gٓ��e�w�F�|��ct�,"�*L��F�Κ�M�{u�M�~?����,~]���$|�9�hLpl�q�%�_)v�� �CђǢi�R��1��y!뷪}��_̋��Pu�DW��@�x�#��>1����-z�-�m�b�׶�7+�C��r~���4��*��
Y���=Pk;5����H�b�r�HinV:�:�ۮ���zX}BrA����f�;�Nk� ����Q�T��l[�6���^�/� �1ߟ������K���=yLß���ř3D�Z��-�ط/����:��)�`�p���PY��i{��{���dͷ�]q��H��Ж$}R���QvZ4�抡E���4�T{���/��4��iT}�����1���oJY���᦯�`'�,f`uŗU��M�βn;\p}�q��Z�$#uv��)�Et��X����6ƺN��F�+��n�����ۄ�:Juc&���[ŹQ�	=���Uָ�����'G&��Mv�"�&1��͔��eoonD��K�ŝD�������ۆ�q�=��H94�B�t��ȍ��n��ڛ|��K���Tj�ɳ&dtx�x���K�i��6�K\�7��g�U�"O���q��]))\��@b�zi��&��U�PӚ�4�s�o	�6QV0-̊��|��� �����yf�٣#+���َN�;���d��Rg"�6h[Å6:��L��aS8��@'�ӷFu3���ה�����:�[����t �ꓑ�%t �����CWd>�r����7�l⸅`��FF{B���8���D5P���L�Qd$��'��K�+�S��'X���[�h�<2�CT��V����+.΢GdZ�h�VH�9Y���Q)��*or��崨��{��ǥ�ز"uA�{8m)��n�\���dX<
��4�3�(����ݙ�*1(F�9N�Q>w*ᣣ^(_3 ��6�"�uc�e=�p�&.��v��7��� �bN�W�Vr�z�7�������_��f�12�?��7���n�giq�kj�	���=�Ny�I�󘮂�'Z���S;!��ar�@�xKQеʰ^uh��R��0��Hd����]��t��[B�>.��O���-	՜9����Ĳ�_Z����c�`ѷ<N�d�	���r�L�5���C��k�Y�M��2u�=�!�;S36,� kz�i�Vdf��Z��9�T��NͰ�o�ܚN��p�Aa�����2�Z�S�q�p��u��eӘi�l�$#|e	�ۃ4_=�e>�W(�ro����ɔ�nme��m�Z�U���Ͷ�9��K)/3Hл1��	���u2ԓ{	��k������30�J��AA���N�o^eg@�UV�~;l<�1_=V�`�7.E���j:u0e�U���Yd��}h9�B�#���V�FbTwېp,m��L�]Y
Tem��eiM��eTw��R�aW8�q41,3�{qX�t��JRZ������㬍��X�Wˌ-ƍ^���)�u��G.���߭j�6�',���|�N���\�oQ͗�y}95f���	��k�̘{�j����ĺZ-�z�pe��MnP� 'Vo�3�njsY��ҝvRN�ʐ&ğ{�O��#Ȅ@<߃����UD{�6���v���݊*`��������'���������=��7����������||||}��EQ2KM4~�55Q�i�Ӫh(�f��Q_�rt�4m��'>��~=z����=z���������~�_������\ΊJ
Jh(*�I�$��k�V�٪(�C�N`�q''I�4�D�MUUDPQIEV�j��l�f%�����C4D|�s�W��b�"mLT|�"NZj����s\54US���f�C��*
�3��H�*Jo�PRS2�����D��T�ZR"�j����9��M��$���l�T:M5MU4�%0H^��r��4M.�[��\��ִ��{��bJ&3@W$��AƊ&
��U_��AS?���̮���
&m�r�{j&�T颊�9&���E�I'���,�)r#"N(�D�Cm�d%516���0�5��g��^[o�6�&rM���G��j���9�h9ij�U��}k��0�Q���z��� ���I �A'��-��a#%�$D�9!,�J0��Lf7 d��)�YDj�5M�$2K�bכ�/��8�'����"����ӟ|<Og����Æ����`�"[I��_��w x�?>��?�M��j�����x�Y]ھ����M��ja�}ԽR`+z�sӖ���=L���KD�BkL:lOB]������I���i�;hq�l�6�g��(��Fɶ�C���Ő��~���}C���z��'_lLd�n�i��gQ�5�f�ĈF̽�ʨlu������N;���c��zO��{�"]�`�#E�4�& I��b�)͌��m�*꨹�h�@�������{�� D�I�Bo�\�����}0�4;��kM�����|�S �x�_~��G������]�xB1�������!��R+{a��fnjJ���g�f�2��lxZHSpב3x?��r}3�|���|3��{��a���s4ֺy��^��^�c����c�W����E�wވɳ+�vF��C������<[�^��t��&�s^�؂��&):ħ�T)5��Q����㟭������Ŋ�v��ۯ�|���8�:#�~���|�xH�����2O~bS�e*�L�C.�o����]ǁ*Uo8���a��iYӭ���qb3�C*���/z]����J�,i��N��� :�m��X��˥��Z�Z����<���>�FE��p!}9�bS���l�g�Lx����ܣ�S#�`����L:'���U�7� ��>�Y����t��g�YI��xX��hqa������5�AΊ��>w�~����R}��)Ǐ*�:�|y�C�Usm�y�b�@��&���8�,}��$v� �p�'��0#���e�\�R�q�j-�/]�1�)�iZ^F����~c�065�^�УN_��2�қ�N���p��]K�{�3�=^��¯���w�˔^�%%�4om<y�$}'��r�P��!Rӵ��=�����[�DxI���ϵ<hYc�Q*y�ΞcW�u�$����،�Wy�l��j��#o����x`��T1����Ȑa1�05�wo'0q�bS�����BOlC��Cmgƶs�q!���U Bz,;�p���g^f@�l�f�uBa��}�E��g%[�:�Ҩc/ٙ��]��D}��K�E�i��>=��{�GO����`<�{hh���?Q�1��ris�����#�]�M��N�h���nנL���
<#�����C��7�C�v�7��U��g������"�17�N�/"ˁ=��@� ��;L�0���@vǍ����r�7{z�P��qD=ۄfJN��=5�ƛ�%�_A諟(r5曍�M�ޔ�A����u3@��mc;��|��˳��Xꨴ��8�72Y�Ek��^q��`�ѝ0�eS;H��FGd��ǽ%o���>�uF�Y#�v��� ��N�zri�GFm�ٰ��]�.X�z�	������-�\2ۦf�/������2�d������P���"q�ǂ(��?7{���z��N=C���3ƈ�����5�A{����ҹHZ�X�  ƭ]
+mLf��Q��Z&���Yz���:̜a"��. 6ƺ)��?�q�����n6�{�9*_�~��5�x��*z9���׈�ß���֫�����y��(�T��G@���� �G�5>��ohm򝻨�����T�[)�$ca�I|&��a*~�����n'��x)�'I�t'�XC��7��R{��h#�>q �	
E�׷�
u�bY�oJ��2��i0�ؾp��SJ}k`2�������XNZ.��!@.�0�t'�3υ�T� ]�K��J.�s�1Zf�u9m��8'lk=��gUW���S.͌�fL�G7P�	�lȞ�'��;.9���PX���Vָ�3��j��\5N=��/[�w�1��!�yG�:mi8F�TėQ�X�Ѥ��*���]�-�S���Y�D�]5���o�� 󯗰�0|�'��'��1R�\�lY��˄�/UEѺ��z��$y�"��N���>�os]���@�@Ű~��3��������馯_��*L�7BԆ�w��~v(��N܅�Y��M��H�ÜBy�ŖA���W,fS���t賱�\ݰT���[�aZ�]eu��v�Gw6��@GaA���CWL��7y������/L=C7�Cƭ���n�|I��ѣ�ã"u�p~~���x
���� �<}����q)c!�fg��^M����ɍ��������N�/ͧ�Y�z�{�y�5{�����gkѶ�,�nB�iݡ�M�Իk���7���g�I;h��I�Ũu�v37�����!�m^.x�=u��H�)ʪ_p@i����G>��略�������!�wA/C�Z8�v�g�\�cqy:�kv��m�o!Qx��cD ZZB�b�!�u1�x[�CZFn|�^����KV���bb�G\�v$=�����Ԃ���*����T8�Nid�����p�^�JzьplŲ�_�0D���M���m\e4M���gH������O��T?h�y<����2=%��>�O6���|ʴ���~w�;Ű�2��8 lD���)���[=^cX��x/B���؀l�Mh��W���,1DO���g�#EL�֭�@�%�x�F%�%��";��Ӂ��zT�<��Uvv�W!�>C��9�)�T�`o����y�%:N��?�"�A%I��]��ݧ����7�vn={�L��Ú�����*q�e�2��ٔ���Q���'*C���b%���%�έǌu2�*�nh�UwIB?�S��ᛚ)'�ul��u`^]����qc��zhb�9(�-g�m���b�Z-�VOA�mʋ
��M����A��U�Q��)�Ӗ��݁i��[]"U}:��H�p�L���'a�����x���ZA���@|
�o��s'J�m��t��C��^�5��0��Lav���[ͰA�;��La�m��w_���P�4������Zq���V�=���ކ^���R	z���:�Fi�����>dY��X+aQ�0�m��S����tj�㧱!�ۗ�5�v)E���^�J;��>X���ĀcVW�"|5��.�ʯ�ӹ�C���n\^�-���C����D�M���;����'�>Zd�ի�� �H�b�ٶF�}�YM���i$�f�\���3���8��<3k�n�9�è�k,p	�������fv�2`?��ĺ�t������|����T�C��G0"D-"Z}�,S�{���6#�m�O�S��	��=��f���.�ܜٽ��݋��ՊXkڬ$x�eT�E�����X�c%�>�۽�Ċi����h�|W�*u!�Ǟt���`��DYz�)i���$�2�[�C������_�ʾ���H�����Wگ��Qi����Ȟ���쒜d�}��<5��9��x�� /�³�t�q��mD�+��%x��_����zr��4����.�sw��!�1���8ʆ@��B��r�ě���3��5��׭l��_}̰5�]'X5�ר�s��n�z��J�i��%�!��C���v��#������B�Y�~D��a����:���g�]ے��R�Җ�V��>�.'��9�hB/�C^�,�H�����Ⓦ��Y�X�sẦ������� ���� xxVn�J
{P�	�F���������o��n@�P%��c9~����}1%�_n��#�oP��3�a�)V"K������t�=�E��z�LRu~ĨR�nseA5����>SxF��d���_U�+�ABa�
��I�.5�M���5�L��2ݐN�bZ�ۜ��p��=��O�ڕ7*}I8����Ы�q�!���A�Ðʟ[�eмP�o�3 '��h���y����w^e1C�I}�H��nz���v��FdW�B%��~
7�6����N�zX8�A8�SY��"����1L���,�^���[��I��\<RU���_��08�C�mשr�>g�z��0��y��D��bW*�	��I�z;5H�f�x�]�O!�w~t��_��ōDݏR�]Gp��d�,)gO1�
�X8�k�y�j��W��j���T���0g>2�k
�@�W���w�K-�4.|�A���z��;c�ő�YX��҇�������'����9���J�k��P;���뷝'���4�s��\4�֡�i�u۔��)��8u3��Z��������~���ڢ�^�F�;W���l"�wb�#��K����jn]4��-E�	�e�C��q�2�$���1���Cz�/�9��s�y��??����+Ǐ"�����[��.|)KË��3Z�z�hsI�^�{�3p.C��#-���JW#�k��n�#���oe٭_N��и����I�cE?N�S�/�A\�j�+Q��;P�$@Cι`��ط6��^E�N��\��8�v;��s�3xe��V+�����t(�p���'�>����"����TUj�ǆ}y�Z�}��B�ך�����C��w���_�Ϳ7�N�Q��m��i�W)��d�{����˔���1�eܝ� 5�T�=w093��`��@ �mJ��)��������MGΞ�a�����I�b��I�(xՈ��	�J�'�nF��f=z���p-��ҜK\�"�ĆT���5mF���]q(z���즯>%�����JK�!%B�F��Z�ΞE=��amwK�7oH�[2yO�����'�y��*��fj�<Ĳ/z����0lz��s	�v�,H�om��:m���0A
���<79}!H�����]0�jQu��Lii�˱�JQS,F�U�u��ܒ?F��i�vu]'��@>���g]i��L�,`%n�|֪��3{�|�#Z /�{4M|�H_gF�Ih��C�7nes9���v��?2g_u�T^H��w�km�h�|�VA�#�ٙ��L���{�����1�<	��z=���ae���vrƻy��C��f��@�0`8:m���"�A�7d�q�~+$���|���d�[�K@�������۪�_=k�ߓ���C�0B��<{DkX���7<Ú�����)W�mY\�T�ݼ���S덛�B�&��ܨ���*���X_�u�9����_�b[�y��u�e��\jCώ#������I�z�!\S/b�>��`�s����B�����l��Wոr��3s�!̓π��u�8���S�>Xw���I�i,���p�*���w�Tm_o4���!�a�az�n|��!�~F�����϶�O�I��tc�W/��\��}\q�2��4�!�P�eO�a�����_%񒡻A�:q�7s�s�- ��nv܆i�舊~K�i=y���
^Ĥ���L|e�����2<�����t���kv8X���S{�(����[Z��8Q�.�@��O^�xi���ޖib�38����5>��2�wa%\����8J2��-�L�,�Ԕ����z͜OC��z�P�x��a�u�i¥0����X��"�kR&��D�e���d�,�P7]t)b��J�C�V)ý-����@mu��ԻݾaJDJT�WΣ��W;���6밋�X:�&�wZ{�bV��}�`Z&wZDj ���_�2�Ѽ��?>y�����?O�A'��x�x��"�z+�������Z��c��}�݁p�V�!V����hzW�g��s�>W/>�D������}H�8���W>������B��L��j�{�S�HD�Ɉ^@쀤�Z��\P&%�{	)�V*J:����1����WZ��*, �_>h����.���G��ҹ��2O �ӝ*E17��ڲh����)��u�_��O��Ć�G�Us�����Bc\��􏠽���z���zW�"�S�I>���lT����ɛ����0��c�|�<�aA�"mLpm�_�/Q��>,�W��:v:��K�} ��^Z^F��&�H/ ��>=1�Ð�_�eos��ٕ1tڎ��BLK*�4*�}+�(��\
��ܨ|�y�=�4�~�Ȁ|5�Ú����N�7��8����L�O��%�Hz��M��G�?C<;�Ϗ����l!�Ke創�p���wvwL��#�>��9��}l��Bչ�è�e��'�����M���sN��{N�kg{�\��G���
�(|��y��_~T"3�#�[f�׷�'�1�'3l-���vs�z��z���Ӿ�Z�ј�y���9Չ����S���3žᶚf��W\kAw�;�����i�U�����U�dY�v�5�n�s5�z�!�X;f4���^��u��\�r�L.�J��]:�}j���R-����4:>~���T?_��x��x��*����Ͽo�b�}V���4Zy��5��#^�ѡ�����<:ǫ�	���A��6��']��5p��A TN�r�ni&�:��=����l��EE'A`y2ِ�r���J�=��kW<�(��f�9� �uw���J�Xj2e�A}kO^�x;���������dJ�"�w^����󇗶6�O�@VM����q|�77�Hd��ɶ\���m�J�m���Q]�Vk�+�c��`u��v���qrP��i]	>�@���X�f���m�ަ�ȧ��]��$˄*b��{`38��.E������S&�\�ׯlGZ�L&W3�NTY�A�gc~���.����Y|�"Sǃ��Eפ�S�O���[���F���z��3��w_��㶼ԕx��3�I�>Ű�;"�F7�H{h.�q"�:��ڟ��vOu������1���$}��L���X�(���^~�秏E��
�  c�ʶK���,�n�/��Ut-��0Ol��oS����x�/,���9�����MsӸm| a�C�Q�a����x1��|9�xluؙ��5��֮e+2�Vq�u�E�.vP|�����glݷl��I�e#YΤ�8�J�n�ꗼ��6wn7<����wd�����(Uل��R�_v�zq�z���h�npg0EO�Ӡ١��N	#;�n�N�����-�Kz�Gm�vG3N¸�@�N�s923�+P�y[�1Pù�:\麒��F���0%�ѝg�ZJ�ږ�c�뭡��xl�Kz;pdeZ����ӧ�$��gf�B�+�4d^q���h0t�ZnYg	�
�;r���u+d�3�2ɸG�E�5�N�y�X��ʇr�).\�g%���C����?���޸m���������2�8��i�\ۡc$�曍Ƃ��On���j�dQ
��B������4Uū];!��w7c��&�eFh���hiP��v�[��t:+v	�.�s�?�����OV��O��H33B�,�1uJ����l�V�'����x�|��j��\Pt2�]��E�ײ�=1���NfP��Q���!G���:�Ҫ�eq8B���u$��kF١���Β���z &.� ��|/��t����N���U��9'!\��]�ν-b������*���3jMLH-l��p]ӏ
9��{ �F��k�iV=v]�lq��Y��fA�+R���l �iF.w�_t���q�W֟:B��Y�)�6���Ʒ�����_Jb�
GB7rP&�3�-+]�jވ�&v�>��ϋ�h�=�}�C��W�n8���5{�n�t��O�R��&e��r�*�X��1r3�eQ��ޜjb��}n��]�D���<�����7�̢�S-�:^i�_ Ԛ�ɶ��؎���ʏ�à�K�:�d�K�Ҵ�F:�ާ7ut�41��sn���W�aQ� *��kw��䢑xmA�%曻v�<u��t����͗�kT���$��5sS��0@���b�,v>�b�984�IV��[���^���I�v'M=�c�P-���A�3N�`�=�vٍg��o{4�P��E�Z�k���*"�:��m�Y9�+���n�MICח}�-���8�7Y���:Y(E��F�*|o"�.ť�:�upP�ع�޽]��l��sv�y2��%���J�wI�)�Z
W�Fbg�阝����G�X�� ��K���1jA2�Y �=�������ʾ�r�i�6c�=�����g�p,]x�J�{:��G���*�SY�i��r�J�W�4��#n��:%hz��Xaܭv6\�����RQ��m�F�tQldUw��c�9fA�7�Vܶ0^80�ȹ�m5"}u$"2ou���.%\���.�B`�J�m_=�\ �)���H�W4f�����,�Z�=:��s;����J�SW_����ݢߜyQ2��AQUA{.�)�h���U��<}~?ׯ��ׯ\�����������~�_�ښ�d�����������"ӧ��cTU�nX
f���h�y�b���x����ׯ_^�z�^��_�����������Ԛ�Ql8�PDSݨ��&#�����9��hh"(��d����rt��Ql�J�8�-���F�+��TG-Q�45DM	qLLs&!��N����9�������5�o��KIHP�%���#lURQ�\ �Q��S5�Pl)JfZhBd�.|^'(������jZ�lO'j�r9"R\Ί*��E�4�)Q%UQT��CȪ�&��Z�f�I�=� �G�EW!�"��?#@PEKH�as�J���K�����

)b�$�I$}�A�3���üp��0��9�'�M掍������oQ3�&�f��!��R=j�&V�o^�:�5�����{��|��Tz����<x�"�-�I��S~y�>�!��K��0#��ԘU� y���/iAcK�C%k˽�J�}�+4����,�
�/���|���L@-��D��O�<h�']�U;g�ع�8v�%ݙԿa[}�i�֯<�4� ���
���!Y���&2�n�9��ٓ�,5���;7��Ӗn�i�Om`*�a �ε{w�p�3�69��yeu����B������#\,a�z�G ����q�]�f�@����́��p04B`�%��o�4ҩ��]K�sK�; Ľ۳Z�I�a�&(ݯ^&@�>:"��@�r��ywF�ͪ)G�S��gl�fa��({�&b���Pt���3i��݁�y@!��y�����%��T�놘�9���r��p�h�^j�#)Ĉ^�t�/V�ՙ׎y�_A/^*�!t�K�0�W<�����ׁ��U���-yg�b�Ă'��ɢ���
���B�&�p�
$�x'V�tټV+��	��6-�z�*�ئx�-�'-bG<��I�iD�b�.�L��^v5C�e�]S�}���!��\�+�� �N��%�f���*�F�6����Up��mV�X���s�IN�-T �W5�5�="�͊W�fե�=��7���.�z��#eWR[�?T�ٯX����A���y�Y�ې�Z2��d������7�<x�	H����~���Ϟ�YP-���tImJ;̙/e*�ģ�(~瘨Z�L˶�/�$~�~!�ǥ�k��֤w���S��5�:���X��^<���wri�ъ�)�	�J
L��M��=��J�Oj�t$t��`�s/S�>C�ς����oHޙI�1,�ߵE1��&6/�YWy��gm�҅�̓�A�m�Ѭ���SyV�����]g<Sc���**%�q\f����C���y�6� �Mf��m��+̛o:D�̥$3��3��/ �e�<����.P�����8��;`>ߨ8�w�6Ϟ�<#�D<>W�5�\mA�m֦�G{h%?F䳩������\�ydk�%C��8��^��n@v������s�S���cg*763g	�-S"[�i�a[�V�NK�9W<��el[�!�9���*}���VpѪ�ق2������m�V��+�r�şSޣ>�S�Ƽ}��	�]3�����
�e=�}��9><�D��S�|sU�� ��^�/�^=-#�@ܯ�Z>�e�B��r�D~³ӡP,��]�rģ)�Ӄ:���Hr_$-~�f�o�M���c�5nc?�啯A�<�Uq���Ң�'ĉ�+rWΥ�U�Q����.�Վ\d@٣�%��\`�A��x�!�Z�u۹B���5\9u(J����������~~~` �}k�~W�%�g����v����r�V�t�]dld$������v������� �R�ǆ���v�\���ci�_d��f�2�������o�/jT�f�W��3�q�"<]'�/v�o۵�ԃA��E�SJ�3ǟNMJ��S���B��K�����񖙡��>0�>Bջ�~�ա�s�9��G>���=����+�i��50�uy)�����ޝ��{gSӍp�08��D��nx�P��Jc��L���ё鞋a�@f\ߩr�m)A�Zx/�������o�b��
L�,΀ѻVcLWz2(��.�@�yYMʭj��\Q1,��JO��J�4��ӽ��x�y�v���QN`��1����B�������U�ݒ�z�{��!o�'ǘ��Z�B��^��W}�[�ds9<��F�Ǩu��� ���B�=�//����}3g$3�>"nkt����i���쿩^�s���"�%E�5�3���xض���iD&꘰�i��u)������P�rv��1�@����2��+K��=4�@��1l�(ְ ��0��љ/�-Y�w9bҍ����QW�n��ɳ��*�ĥR˙wۇ;����6�{�0Lm�⬲}Z4>�VJ̼UG��Q���rU��}�*����L�9>��$dʷ�`wFX:{5�ye:{ژn����7-e�V��������`xy���� ̫��:��p�=���TKm�H���D�Zo?#޸�!�X4|�@E�㷵N�4��uk%p���=�Y,��h	����MX;�'���ի�W��	��ʩ��s����`�N�̥�3���t]ً���}l��B�� �0�/ޞ�:��=>� ���'hj����k1����=�${�`@���:cC�(~��Y�K�	���Yoٷ��W��L��⨷c�9b�ōxg�h�gk�![�8L�s7��Y*s��;��6:Y��x����0��$�wtE���l�bd�-�5�=���M�N�-Λ�v�mЇ�E��l�Q��;�|�ځRim�!��c׉m�ؙ��^g���n��(Q"1���)���Ȧ@�C�����W$5$d4��k?1��C�<%��ң�n�iz�BY���|��.[��ڢ)�uu��?r�����G"1@�5�{J����J޻}٭Bjյz�1j5�5�W��f>C<���+?�G����_�|��j��~�g,7�ʨ��M�{�1���D3YWrh�	�z#���5�%c6f�O>� ۵dr1:ۭۙ
��C��F|m�,����H���b_L畔���(�)܍��v�0�:�	��V�ғ�ǜ������꿀�_����~~~c��M��fZ�8����p􉿄���j�����=��By9�w�>���p8&�H$��e��p����u�=��o&64B��]����ML{��$hK�N�؎x*��w��
 ҳ�0��7��]"dp~��>��H�"���~�/7�o��-κ���u/����9�8�{���|/jy=�b�X� ���7OMs��zC!�D���K�S�6�C���w>z]7H�"z��0���w��=����y�}�����Uy7+��%����Ri�s�B�#�!�bm�	�EW�*��S����T��Q�g376�:�޺�Mԍ�a%�郕 ����a�����ǫь?H�k0�cr7r�+�@�f��{���!F8C�JװUzI|l���ka{w���y����p؜�K�an*��d9i�m�h�����s!����m�`N�#�|z�X/���t�g"ݡD��v��"�<@�no����f��RaDė�a�����:"�o��<��{7�e��~[��W(�3h-�S��><jP�r�"�oTJa]c�P��JC)up�X�r7���`�ɹ@v|���{�'ٛ/��)^���t�WW=���vP1	�K2�b�����zvB&ٺ��)`�$b��n�PV�rnΜ*�0����M��������>���G��� A��;�O*]�<E@��σS�dS�g���m"��݃�*�����h{��&�����^.:ݳ�S!O��{3�"Ə�H>1���fZ���x�/ ��P��_;9,P�^�q��:ȗ앛�. ����<e����lu<j_:*`tC�/�A]��d^�m%���c_m�YlxKՖޱ�h_:a6�A�%'*� "z㦿P�E1�b͏��m˺�i@�:��[O���RUK7�F�$�߉��W�*��g�9�x��4����O�f	�/z��#c����"BL�C@�S�O�Ib^�JK�	*q����{gOT�ۆg帷����3�&�A��t�+��ϯ�7ƽ#ze'X�%�{����J���ou\����;6m\�A��s��`\�
��~���Fg��aX�8���0ЍJ.��B訖�0�'����_�+ض�Q��-A�6�������;^�|v_A?vO�����q�EZ�_ڪ�y�2(,h.�5������~$O~�&s�*�|QI��ZfpByІkv��K��n���zi�T����jYt+=y��鋨��BI� B�vި��΅k^LW���|MK��:y�6�`���CY��SE7!R0P�ee�pYxn3W�M��=9]�Ϯ���[c����y�y�=��{���m�oB˱��My���o;ٖp����7v�Y�$o��8��E��*2�F��	P�zY�|^��r�B5�{���ݑ���H.U��ڰ�
S�Q��B;�o(X��^��8�U#(l[�!�4���R�J��殐�!� ��0�[Κ�-ؿ)��P�ǣ��'�Y�(��Lm�����fb�lk�S�c=�9��Cj5�?*�L�$nW�;eN�/�ǥ����ڳ�N-�
N<̟t�闩�����O��O(˼�a�q1*l���$۲tgV����ո"9Ү��V��t5sH�F]���k���5Վ�2������z*��/�8�5%�/�����v�0c��P�����WA
��zzE��z�m᧱B�v`�|���4�&������D������=�]Ӿ�o3y3�f�0�rQ[��,B��z/�q�H��=�I�?]>A�ţ����켃�y��O>{%�Q^�	�)�ɔ5Q%���{_��p��}1O~���t"3j��s-O�3��6y�����#�7�,p�w�N7��ߝID�̵��E�j6����htW;�T2*�L����ުV�<GA��'*�~����љl�=�vYV�K�]�	 �@,��3K����P`���ږ9�F;&*���P��l��{��"�@�5(�7���ή��l�N຺������������=���)_a0���C~u��>���:y����Bx..�{�t-~�'$�ع�[�<�Mݖx
~\�Su$�2�<�u���z= ���	K3��+�V�0v�;3+X�N.ީ������̗]V'd�M�(�%��s0�>G�Ű��@r!6��!t�ɋ�Gz˴'�@���կ�a�0��n[ŤmzOU����"�A�:����{�졨��a���8P��^�n^�Zg���#�}��z/I�`��@"������U1�QW�D�'g`��K�:n52']T�n�Gu[]�J>P.3��Հ�|���s�Q޽�CEӸk�-
�H�^��P����o(���������i�zKe�Yc�Ea��]�U�4��{��?~[a{`H�h@�� &�E�o���Fᡢ1�<��7ȹx�Vau��^�s��s4¼��v�ʹ��rŨ;�׆x��с@��V�I�3a�&�QSv�^��t����#*�и��_��knƊ�t�96&A�b��ol���׹�7[vn���nm&�w�]u;s�1X�F	�*VE'|ҾD������R��Ù���b(t9؄A�\���A&��_�/0m�Գf����m��M�t���Xcyx*����[v��>_m���0���NJ.�]��[�C�E#ViZuW���>_����z  
���B��ٟ�3���=5���6}�hMwo���!�F]�kR~h���iE����܆�nOO-s](3��6!0k{l�ɸ��E5��	/����Hj	m���b9�6vO)y��?��e~4e~�
�|a�s���:O�� _���D���K➾�B����g����T:��� �]������'�Mp�_��+�k��ln7�θ�˃isom�ZT)7�U��ֿ]E�ȧ�t��(2.'bK������g���s�n)�d�\�/��J�A��PJq[ cǦ�����`�;��G��_�W2���1^����/T��R�pc1W�7H���4(?E�ם��1B���M��s��:�)�?'4&�n!�����i�����Ͳ��X���.ב�s�GÖt���vs8��_]��@�a*:�Vփ�*���_�3uz��
����9r��տr������7��ת���w�˭� �kAÍ���l���B^K����w�d��������R�9朋La��l:�þJ#6��|o����d�-Vu\���(UG8����w:��hR-ͷ`�daGʃ�z�4��1�L��U-���୧R=ɥ�$[���E���3��I����L����4;$�M{_�?��8���
<;��{�����2}��~xi�LiT�/m�<������>�K����M��l��9�wQl�,_e���@�gu�"|is�r^��Q�A��i����0B�_��(\Ϡ�X��j{e�Kr���22�����Û8���r_�w�j�4��e轆s=!�'�nĴ��3��t�3� /s!���8��1�(�vmхW0�bK�&�^�L�:����]<�y�TM�osMt�L���<C�w>yw�T[#m�"|g����W|��WݶW��7����
�.�A�׊xe��e�����̵�<2��蜔3�2W���"oz�f��p�]b�	3��t��Ցj����'�;�^ӟ&C��F]+�1֭M�\Vol!��ݐ��a��i�X6��@fǧP���5�L��m�7�LN�y̛��=G_9�n7 B���k*�����L��ҡI��J8�(�f>4��X����k�;��;�Wc��*d�Kk�y�}��W)��Z��NR��1��}��@ óh�?�lq�~6��b$��\T���LBʼ�lQ����X�eN�+��xN�VV̸�me����Lg�5۝��5�2�LC'�e8g;81ZN�43A9����[���A]8c1ӤR[����8�A�v%҉벮 �Q�pf���tB֔�;+�m´R�����	�����ZK��ō����fB��Hf��_V�{ZФ�����h�r��ѣ��%���(p�4E<)�5�΍�)�3�(can��D���Ӳš��V��8 KO�x��v��`�0�6�1f�R�@b�^
�=u�5����t���B�o=��J��f�{ס���ݙ��RMGX&��3�!dGrЏ^c����s<�yiJ�5E7>z�ʁ��Ǳ
��1���]�˧��������W��Bf����2w����2�ֳ�Ӗ��U���)j�m]XW��Kh�g��j=���OM7muǩv��|�d�jbѼb���{�6�/�螩��fR�><�bbܷ"4Vf����l����l�mT,R�$R�DԻ�[��M�\�wJܫ��3�ڎ�ѣ�AP(���װ_?r�6��:�v���[
>�'�5xj������U������/T�������$���c�%�	%L� ��֓p�g!��w�'Cve�l.���K�9��ehw
:��κ�@w�{CV�s����ȥ�g��o�
�t�6aww�E��~)ت!��#w[{ ӛ;�w	Kǹ�o\u���A��VFB2�꥔/8�mS��.�['{9ab�m�˖vT�AH�-�ehUs&ގ��k_M��wpx�iV�JoiY��F�nsc"Z�}�-���j��m�&7De%ِ���X/�ڰr(n���&>�+�B
��c�Ӹ�tg�������AMoh�����G�A;9�S0e!�rJ�+�{�}ǈɱ���41�7|�=rX�����$X���h�BKy���o8j���G�~ ���J:r����qr|,��������R���Q��l������4'F�M:�|� �!�X7�cj��ۧx�r��=uoo�o�]�͓��H��u�%�����uդ.�u��˔��Mjۏ�t��*�N����N[-n��z�Dr��G��{�V4nt�6�d�<Y&Q�"��!�3]%��XUH2�;}���2��Ӛ�O�Z��(�����1��kWw�� ^N����0uk�k̺_<S'[�����0#h��z0Fv4u��Ll���c}�{*P۫��u�
̍C�N^�ܛb�%iX� ��TP����b�s�k�N�'6����D^�0$%NCyw�zr��#��)��]�yr$UV.<[������.��V㬅|o6�&9m��� d��nRD��m�nV�{��4Clj xc��AQ� �KN�������^��z��^�}}��������~�jZ��~߲�*��:���>�r��UD4��z��~=z���ׯ^=z���~>��_����>��v�X߇�!M4����ǰ����+ݘ�4�+����h�($4[?9������̕T�M%>��r.�< M:4i����h"�uIA�Jv�	���+��b��Ko�rcJ�O�d��4�i�4:R�M/�����U\����4kT�o9�+�*xAAM��9&ԗ�J=�G����|�F��4>ZNmZ�8�my�#̓M4�:)k�w��15E%���{�ߞo/9��z�{�WU@�h�FYi���0�ͪCV����!��D��w!���.n}�Щ&aWԸ33*i�d=W��+r�'XcƧ���^�me�0�GZl��I4�Yq@b��<c�J�@�H�YpLm7��%I���.HD��^)���N#	Dbm b��{}~�`���=����~���"��&(�ގ�σ)���J3r�VQ�Y(f]�o��JVG�^/���k�:/�逓Ⱦ�D���ze'�,f�����%]���n'����|+�V
���f��!u��#�U����}?%=��h�[��Bhf���WlTr��Z���728���;���4y��:m���թ�O���'ъd�v�����p���������%� �T?5�Z}���?s/��״;:�}�{_��]��7����˔&i��~%Q����e)��di��7 <!ú���gM��N0�����Ĳݙ�#���{x�״���)�\
�Fk������R7����5���7H0e�4�D�����vl��Λeqʆ{����>�z�Q�P�&c�_���,];���P��=v263�A�{����W��>N�l��E���ܡ2�U�^2�_/p��0r:Qȡ 3��	���:�;G�XD��L#���E��/�>Kv�W��2	����r��2ak�&�g�~�`�<�Z�kv�V��'��_�_�������x�;��)q6R�̊��Mx�j�S:��V*��� ���v�S�xc�OT��YӸ�y'
�����,�_�:�|aG/	�T]��Y�.݋��GqO��[Qq�i���c*d�gDn;PZ�1��Z�fQG���e+��/o_x|=^�}��z=�xz�J��椧����}�ʽ��&�t�����R]�����C����O�K��c�~�Ff������ ���,Lz9� �\��o���E0-���3g�ǶtHR��m��m��κ�߆5��#��B͍��S�y�1/>�."Smzɤ6'��}���h?q�G�{��3{xr�(�=X�!àf��ɘ����#k�*��lA`Y1,��k�ug��\�ԟ΍�_�}箛��e��,x/��^4S�qp邭�Å��{�c��S;c�86�/9�Jּu���u�7�o�J�[9�EÞ�G�A���C5�r��a�ev�:Wv��F�Խv�P�)N���f�w�˦T6�3�5���/O��׶B<v����-bs�Юi�=]�C�Ɯߞu�z��Þz/�2�PgW�M�ݪ]��1�=���b^~�}uu���U�S-�W����ۥ�z%��H��Z��' &2��w='�q���?N�0{��ԗ軃vu}n���3��@R���r���+�A���.L�Wl"��<^�����X�?Bz��yVe��2�$C��H�ь���-�R�/f�u���v�Wڂ�{��Z��<*Ӎ��� d���|l]L�2fr��˛��̶F���Mk�W)�������u����޸3��$M��"��0p���ӏ�����G�����7��#���-n~������i�����<�y"*��!ֵ�]�������V�!Z�r?�k�~�t���}�M3ܶ������+|<Ǎ~�O�+��F�q��n~�o:�-Q�Y��wP����6~�a@�����NZ��w��Ihm	��ܱ*\�ǫ�z1[KkL�b�z^�	����׬�T(���8÷1.]��,�{����w�泑�TzUjZw�u��!,������֜�l���D����T�G,�j��=�p�������s7�\){ >���}�����e��R��"�m�,�C������!��fN��eQ*�ț���<��σ����a�{�oL*.��[b0���m��T���*���͛��cb�-����s=��6㦲��~!v���(>V~;����ãŻ/dE�s�u�@�"C������^�Cx��ZT)\�,)��8�#�拇�Ol��	-��#(oQ45�5߼!����'��b��e��x�b^Ø��]^�)8���$nE�*��ǿ�;�exr�d��Ѽ�",�ȋ67j��D쎵�
f�U�x���o0��"*�K�&�c�;��ϵX��H��t�G����&I�\33V'Y�x�8{86 »�W�b�T�Ǧ��l��]�����D6��3m�eea�9j�g0�~�����~~~~ <n��8��L[48�zf�Y����4�c��Xn�E�D��?E��[Xյ���j��UJ�xa��{�h��v%��L��N�{S�옦E����K���S������Ste:V�/��:�J���!�p?r�.�fD�z��
��<���ʉ��S�2�TW*�U�����\�&wqCr3�� 8q���l���RK���`z歘�5W���3;���Lts*�X�Ӝ�� AC�Xw�H������P�\�Ȟz���:Vp��R���qƓҵ�r^���a'�u�{w���y��)�R�,3N,7�f�?d��̮}�E�j�J�����	o@���9��/E�3犣�ܔ�cC��M枆�A�p� �gun�0̓��;e��Qa�Iz�0���	�
�rf	��kz�
�W��h*b��;><�^]�`F��� ��Y�����6��zY�7`�
�e}z��{j!V��S�ᴇӐ�hvt���x�(|?1'���~5���*�Uj��#���T˾�E����WC<�����ηg��]A�]+?A�03RS3+����e���2��c�}�����tp.�7n�K���打��#j���	T�Ժ��v�I&t�p2�+p���QS��O/�5��Mt�I�Q��60Po�����G����xx�I#-�	�⼸�rl:�9��N�]E���@nx^��GÑ�4���M��z����t�L]�u�a�] 6֨Q�4�^�*�[o(.�����p�����V\����Д�0�߻�|���-Kv������E�C�N������d�L�)���@�ǰi��T��{����^u[&A�5ĵϢ�>S�+T�P}"KQ1)̈́��MP�� {��:��B�ϖ���b_���e/�ڄY@Q�翖T}��U]��A��� G7�^[�/9����K.�biuZ�+V�aA��9�.!>�p�@�"+Ҙ&���i�ʆ)f�=�`�ݸ�v+�Zc.�Uol7�g�}Gz��/>�����-K��!���u�'�i��4��fЭ�Z�P�^J����z^=@����9bWJ��������C�2���}t��eg�׿m�*�d�gg.P�,5���`��c.�m��e)��di �;���ŷó=�ffo3y�0f`��n�a-�A;�£���uS�k�T)�wN0�w)Z��`��uN�.�9k���[C�*	�)�	={�p�G���TՌ�T���@�d��T�u�~u�]�o�Sx��[�Ɍ�j�������R�"�w9���d��G1Ĝ�o���k�W}��B�K���B��M�(vs8�fМ
oh�w]��̨?��O?7���>�>$3zr�{�B����z�¤0g:.������oY�E2��C��j{�gӮ^�5BK���p��fK4���;�66�Ǹ�������b�U+z��ڹ�Ȫ��}�Λ*P)�=�Cw���� �;<k��"�.-*��W���)M��|d���\�M���{h� �rm�2�^�� q4�[E?�b*=�ψ@��.-��ת2���W��z�i�B^���Uё;��q*���R\eY�~�Q�"\�w�`��~��'.�{���+jd�@���\ǡ<��ǒ�m�zPc~U6��$v��͜N���g2~ox-]���*���I	o�i�?AN��-�X}ט���E�F��W�ˈ����/Vv�Q%�s�s>?l�g���7���i+1cǻt-��9�ݙ�0.lD����V�d*�U�]���I�i��j�<�Ά�4�Ħ�T�����Ξ���A��ˋ�L&
}{#�os�����e�Qژ<+�J#����r�xKR����'�.Pq ��t���zz��,�H�Y��[��f�t�h�q�<+��~�=���"&k�r�V/.��c�:�V�2؆Tc~�QX���ܮ�Gi��IC�uM�Yl�.�R�K�:7C��0q��:��$�]�W.3�w��԰k�Q�F� ���2�_a���;l��mn��G����@���1ԗ;�wdLKC�H`ɽ����^�w5R���b�7H�IQa�@]����l��	�N��N��Á�P|kS6����Z��}{����ŋ)Ӝ�i��q�m�)�0�Vb2�,���a��8�xe�S�-��H���<P$&������q�JJ��(呲��)xw�∯p�>����|{�H&��1.�F��ғ��.��t���5��H�fD3���?}���v�9�Haiි'��Ǐ��c��R4��%�,�[1
�"0(�e�ǣ���i��>h�u�v��.�>B)����ļ�V�l��t��t�ǔ���e΂����	�vf�Ӯ6Nyf�qcF��{v����^R���;Xr	�3\��M��h6�v)�bK��~�nj�w3DYz��L�s��7Y��VfM�c(S�!�5��D��tX������^_P��(�)�C!����I��'��oE�M-��n�%�[ͧ���6�J��{�0���ߞo�	�N���5i���=�ܤ�np@ɰ?/r��-�:���iNB�)n4�vh�Xod�Li:�6��_)Ez����{3�N݂��~G��t��4LJ�:q�ݏ~���7V���gXt5��Q���!�A�cu���O/pӃ��YX�wR3^[��/T���������z�j��Ƀ�n��i�ޛȶ<���3��,�h��DH�0׹�F�<Sc�^��ښ4c�[OJ���2�����l��n*a�3R
F`x.��D����ي�y���ڪ*ndƧ�1����a2�dJ�TXSP=��^ꋇ�{g�L�E���;�c£�U�VC���5LRv�p4Fܦ֧�,Kۘ��#!
Rqw8�q�5����˯s�>t�o�c!��q"�)���phށ�zU&@�LRn�k.��#3��љ�ut��i�6�]x;�xg�Nd�b�D9O���z`�սN��ڞO`��E�zl[|��_5�VsF��v��c�^��T�p^}a����;�@A��v���ѐ�n�hW^u&�()S�l``��AQrvWS�.7+���5�ʡ��<;���ˇ�M��6�켗J�V�,���Oc�4ָy�#;�.�J�
:y�Z���Ӄ� �M`��$<;�~�;�T�v�y�x��j��pX���c!�v�o�=+^�PK�_�G0=Q������7�5<�sC��?�(Ѫ�����<�=�����em�үkr�f��V��'��*�u��w���[�6��SO]�lfz	,�r���k^5���Y:�:�0��*T���䠈���5�	:��׶�s��͏����d9X1g��{�???3��,Z",�1�m����ݥ�+�4Ft����<��"���r�Jf�2%��7�4�S�;2��]���SlM����O`fl���0�<�ڐ���6��gp�a��2���a���s�<����'U	�.K�v;u5(P�Hr����qVᬏb0F5���A���@�S��LS���4��H�pb�32)�Ř�z�	��\`dI�iD[k<�7X���kU��x�M�>�c!g��f�u���ϣl3\�NE�>�����U�B�#^i��thtv��
~�$W��}�eL���Ғzl�읬�\�K���-�r��� ƽj�JN8z͜a71P�)��m��N�3w���bd��?���h=Ps�%Y@g��P��%��L��ґ)�Q�z3ܑq�OJgj<�t�6�*�ᖿ3�
-�'�" "$)��S��D�bS��%E�n"�a��k�<$�!Q���5�*��^�����HqlY�'�} ��>�锝�\�L2�1�17k���1MԓyR`����!>�\@..��L�h ��"<���Fҧ�5��θ��U\�v��x:ݱ�-�]OyR�зv��w��W�7����R�3~�˱W�z�C������{� �4��dQ��ݝ�M�W�,���5B0�I�dw3��:-e�u��[7[j}R���]4��}�Ҋ��]��V�{�0������'���������>��*�]g���Zhu�Y�6��zhs0R�$9��a�5<CL�Uܭ��BP��P �{\�~j�B������JС��'�;`>�a����L���)�w����2-�s;9}�,5�^�EQ�X��{�P�z sH/N�:���d��{�Tv�D�2�Dc�S�Z�S�hmP�O�6ùB�IA/t��g�mvhvF+�Q�U��4H\[���~/0�aٲ�k:m��*ޣ��y�9%��b*�,JӘ}���f��ݾ���Cy���|ZŬ�����3�ŵ�n=��'#o=�C�c����iH@8�Ow�ǽ�af��GJJ~�c��	��z����6f��r?����}A�F}X���/ŜqM;H/��ӻ雗���@�86ᴇ�n�0�l��.d!��<4��ܟo� �BhwIj�e+�q>��N4S�nBf8��{ї����Xμ���0(��a���M���ja�Jm�j	���7N\�5U$�:~�k$Kk� hz7��'#�!�J�L�Գo�86V"��ݔ�ˢ:T�Z�m�	��G��k���iRF�j!ӥ�Y#�;f[ӊ=��
ysM��b���N�dR��H'}�{5c�ЋgY��{p�V��Y;�2'K���WJ���ع���f:��-G2�
ΙI\�������r��[��T�R�������9��q�pؚ��w��l�n�6m�Ǫ�v�%�%v�kN���1\v͕J���s>�HS��g>Vl�-8�\���:$ed�-�|ZB>��'ݝ��D*Pޗ�t��Y�&�	ka����\"�ٕ;7��D��J��1�)0g6\(r�;�{�[v��|Z���hE5�o�d�Z�����D*�|�U{I��U]4,͵h����z)Mf}g��7Nf�7�hCJ���4�AKt��vRm5�V���Z{fY�r@��o5v���0M� �:�)��!�%Ĵa3���j���
��]��[Vj�K��3�l��]�:�R�Zi6f�T�	��WY�:�]��\8r��Z5���X�=�0���fł��h4�ܺ���B�d�&���o!';���HU�Y�����r���z�8���7�Øz��4w��Tbv��
V��)�(�ڽS u-]�U��Xm�݇+uv���T�ni����lz�`El�O�e]A��ʬHv&:?��#l�Ex֥S�Jx�j�����y;��.�d�i�NWj����ڿ׍^�W9��w M)���nv�]۳á�ˬ#���X��h��W6�9�|2t�H$���_B$�ʝڣ#��U�M�d��ln�wb�Y��=��0UB��̳V�o^mYQ��X,��KI����k8g]im��7
_�����c�b4}}���`�����+Rr�+8�h�����NHm_a�Ĭ�7�VjX��7�0��y4Kƾ�$�����_r�
�m�0�כ̭��F���I1����W��8961��+v��L��{�XY%u�bf&[h��h�E*�Ԡәs���Maq���ma}���_	Cd�@����h�����i�s�i��\Vn�0㭔�͋7�=떎�%K���]�q	@k�m-u�t�Yֱ�Z�,�d�x�t���*�6�B�q&�M�"��]t�+$^l��J����ڼ��)r�6�]�.��yհ1�*��܎%	1��1�ڨ�{Aha>�̙B�*���ຯ��ۙ��:���力���/m��U*pT�"c�Z���(�@�<���1��5y�Jb�����2L�FD����u�jW$EK1��C�҇�T��JC-�LPi��8�^���J��j�Y�V���aޑs����}#�qNe�y;�t-��N�����"K��b�f:Y>#���~ܛc[a�<�'��>�p�64�Hm��"�N�3�G-hǎs�����������ׯ�}}}~���_�����i"���4�������u�퀈���袍������������ǯ^�z�������}~�_�ߧ~ᥧ����Ӧ��>���W���ɍ�'�y<�I��cl&'Q4Z
CTQ�5��r��cE9�ca��5|���p�'T�I���DG�r��~^ǜ���
hӢ�$5�
l�
�m[^A������\���#�3��s�'�F����#TnX~O�6<�(���9KkQ�1ͭ�N/�˛$ys��i�4\1l�n|1��"��,���H�	���J�����u��Il�����5�y<#lE��Bh�kmI[cZ�lh<�76�m��V�Y��F浨�<�w�������R��5SR��\ǘ;�8ξ�j|pL�-P��'#�/XT��ZF\�Σ,���nUWX?�z{���7�y�޶�D���<�����Ԏ�Pgx[G�Y�qw�o0�
-�4.��>\D�����/n��뽸���
-xgo��s���0D�c׭���3X�\�,.@��|���ZղF$��N�:�N�g?l��5Ꮉ&%��>�����t�On���x..��,�����0��L޴=���הBd��ħ6��cI*Ml�p0ȸu@ty�؎�ڸ��ʬn:k�e�5��3(tH�L�N�zL���&*�t�4��Laz�@>h����g��a(�ޝ�ΥL����,��cb`��ӯW�]�[�I������s�e5�L8�l�^����I�/Q���P�cZa����z%���U}+�(��˸��[M�������u��t�Q`�̈́5��ôx~��ܣ_�BA5}S���.w^�t�����6�m�dj��-�q2�Ն�_t�k�Ƞw��nc����w��C?��ɹ��S�q�ۭ��� �s:��w��_�s���M0r��h4vk � ��s\{�Y"5���SX1,�;���I+~�Y��̮f�qӚ��j,�ks��2����Ee��Rw���C��;>vlV����+Y��)��t���e	J��0.������Wq����V,��u�1 �c��5U_���z=�����9ϛ��ŕ�4��.�ԛ�ŉ��)86���W�;k�s�r�{�5᝽�y;�`BУos��ޝp����u�������#;}�Ś�/\aۘ�.� :"˨O���˙�e/jxY��]<��+g(\�w�hp��[ү���Yϗ������B�v�*Bs�]���i�um[�ݼ�*�;,{k/\�o
������[{�dO�m�9{6� 㯵�q�p޾I��S]�5`njʌ�&CH��e]>�m	�����a�wj�� �K6�5z�UE\Wold�5<{^��^�Ϛ[t%լ�	���5���X�.�nUnZ������F��Bvw#��2)��(�z�����a2�[#Q�t�����8��4���̪�y�Mu�RU+8�ӌ7��^ƩR�n��M�^}�Ľ��N�$h+���2qv#g730aA�;��y�ʥ̴R���,�q��2�^�b��dO�L�p���Qz��j�mE���=�vh�7FT ��n�T��x^49�C�Q��G=�vW[��"���ی5ߨ�eޞں��-3"�4�Eq�қ̥v��sOohe�֘�^����MƓ9&�S�U�I]�HD�P�G�z�w�[J�o�s�YXT�m谺vc�ڭ�.��lc��R{�O&멉����N��g�U,���y�����o0oX�OLS�x�Ǯ��w�*��:9zxrH�Y7k�Ag��s�m�~OAIy���<���zh8X��?���y�k��m��t(�|V�o��5g�����'��\�HO�9�[Ո!̅�����*��/�=����5}<O��!4�,�6���X���2B���kH������>�E��l_(�M>�|�[��ϑ`�dk���7Fԋ��h�=��f%���G0�箵�9�d?��l&~�mՑ���^*H�����J)遅��'�̺�	�9*�~�ǿ�4�������5AK�Y���$���Τt�g�	�Ƈ�7���~�m��3�3~��P��Y� ���#m��Ͳ��0=1]��}�7���}�N�)��y#��eՌ#�å��Rƅ�B��E�CM�.�tE��x�����(E�	<�p����֌yP��x3�`���˔�~�-�Xf�W#�{��5�Ӧ�z���>�,.!��W�;�w蒟����{�D�zțx`�9"�.R��0�U �Rq��͜a"�*�PNTۥ�J�E���vyR�\e�]mjC{��Z�*{�澂��J�a�u���.WB�S�'�[���s���E(�:t���P[g�W�Ō��m��i���`�
�'m��u�d�P�1Wiff�ᮮ .�Z�I�zo-ҏX=�.��r���}�����`��y�k3��z�V������>��q��%YU,$8379���H�K1P�����N�;��}��]�w��:f�Ǽxi�ۇ=�aY�H�����:��D����u��������7���<�^A�1P�e~PR��[BtL�*���O��y�G3k3��w9Ʌ����Y��ǂJ�
}���s	�\<�!0Z�/����|.�5�k�ǲssM������c]�Q\��~FeX�ފb���1���6�^�g	ف��~��O=O��k��;����&e"ו
60�wt����(�$.��2ac���Q���mwi� �H�x����Mp��h	��ZoI�w�J�/K#X�%��*�~�i9w�a�g	�ԭ�N�x!02(�:�bb[̉e��Xr��iA/t�ovA�O���=ާ�����^�?f�`��:x�]ٵ�\;6[�gM���r��}M1GGR��-Ǵ8ϧ�K��f�s�gn�գ�<�������k�^WE�o+�)K٩[�0fŬh��orho�+��,+�����)=pJ�Pz�]�����]*�v#M4^�?b�ZNc��o/��W�KaR�m��vء@faR�p���<�p�;;�M�AoK�Ȯv�ջ�dҍ��-�ܝ��2�ris�������|����A�6w�˄���;�l'�KOp���>��"��
�C�{�.��%���D����Br���\)'�G����f��(U�}�@��Z<.���-��(t���<3�(�"C����t�'z�`!,������З�^E����k��u�X�B).2jȯ������W=XMv搱vQ�)�0F4�	Žŗ0�~|�鶥�S5Y����,�|�\D;m�mq��W|(U��:�����3�]�X�<�a����((�j꼸�Mn�U��\k�sf�Ple�}-�D�����ޭཱི2	�PxaN��p��x�%�M�cW�3�ō�9�	D�.��dU*J6�}ys��A����p�/s������Fm�Os�bv ��'����DI��H	��)ƂJ�=��d�틇[�>̹��*��L����_�3e�@g�7?��Y���H��w�F�|s &*ۤQ�%E�1/e�en=��3;K]L�:��u���C�����:y���˜���P9�޺kf=�%<�wi�;S�.fdfͺ�o�����ț�W��g�J�o&wn �?xO9NWen�B��B��AxQ
Q_��V�۴)9b�fe�4r����Q�'�t�B$�Y��7�N꽥�R�X����]��=N�ˡ*���w��^^C�`������m%4���S��y4�F���l!�9!ߙk��Km s�����xXDk�OF��{���ުZ<����I����zq�[�p؝�h�����2�[=6��:)a悦�;!߳s��7#rS�Y���R���]��zwf�`؃�>�2t^�_�zP,[v+cS-��)ڤ܊��������hz�L��_��;n������3�ǲ�֍m�-�>6��vO����L�pO���
��ƹ������?����9�ӆ�JY���`xgi��<A�70���^�N�9PޯFt���MQ�?IM�����I��D�v�Ӹi���?3�ߤO<�l���z�g��s�٧��d�I�܏;?���IAp�h���m��42NK�ѷ<��Wb��i/�Q�DC/��c�`eͱ����8��.®1��[*��ax75�Hd��ɶT:���p)�,a�wk���̺Q'{���v\>X�ψu%Um��|ma�P�F���v8���ܹ����(�m�������o��7��rMV�z�����۱�e7Z�$g���f^��� �ҙ�����̣�8���z�`y6U��GwD�v���(�qJ�Vs(�殷��'aƻv+ܾ0�����.��]ʳ/fM���^�/x???��@ .qB�_�����s75���M�2s=/�$������!�v�+?q�נ�1ײa2�dJ�J��}o`�N5uE�{�����|=&l���ι��~��Ƥ]zcS��6� ����LKۘ���F�u	8��m��D��r}����0�ר�}@l������O5�9)��g��H��^�i��0jj�~�ƅr	�&�v�V�y�����&v|F	���w�|gd��`��q��]�2rKS��S���,%e���s�� K���aq�τ|��޲�g���>�nE�suND���c��]���V�s�Q˔�1`%��0�3��܇Ǘ6M�mˬ�,Glg*��:c�g�f�t%��ꄓ@�8�� ��`��cJ�/�֑�=;�8`ֆm��U�5�3�'b���P���D�:��Z��^��U��F����y���Wfn�v�6�=0ow�p�X�|�Г>�vpڝٚ��y�kԤqm��@����f�s'/;U��,�9���x��a��5{���x����<�C�^�,(���:��-�퍭�ěx����0"8g �s/��2~���J�a�d�!A�g�?���jw	W�h�E�x�@l�/�i�K��,�c���vD-��K`�ѻw�Q�.l累�JP(�dW{�A$7��0A���B���0��O0�����~z#����!�=��OqȢ������^�3 �zc�����x��yOl**-��EWw�4@P�����wQv�t��^� ��M7����i�����p�~@���bq�[Q�v&y̚�yZ�3T�%�=5�� ^A/-@_B.U@C}�ךn6�5t��z'�^��uf��T�_�����
� {N&.�ߥ�*��~sc�0�U �n�6q��Yb��/������)T?7�=cč1�`PZa���l��K	�%6�5�	��T);�Q
�U��74���̌ǫz���S�;A
-�����F���)��'Z�H�Ѽ;����%�;�ea6�+xU�C3yu���q��R�o�v��Ο���CjN�� �'��v·���vT5�=v��+�l���������nm%I�?E��s�`��5����^�L`�*���m�y��������t���F�� ���0q�Pw����9�ah�Ulj��0�L���B`پ�&��;��/����֔4�T?5'ٍt�y�]��z/4u]�p6�8)^=�H��Sz�Z�<UĊG2�x�+�i��''�%���t���c��o�S��p�6p݇�a̻�usd�i��N����i�ŵ�4�T��s3�u�WoT;�EU�G̛��~�@///{��ѹlx�/��9�����-0�kH���9����`�����3IP�~�����h�.&���ٗ�j����u��>�Xdz�Z��գ��2rf�0ylOG#Z�ܝ�*&��]���u��TZ셳` �ß��~�@��fx1��ؗ��%��w�����"�u�@�E�����u���i�ۧ`3>���D"�!�����E�
�a�3v�9-��̢_)�6g����KOp��C���htx�Xh�IO��:?��k�E<���3��%�;<{>�m[Ro��Cwt"�ŠM;H/��ӱ�.z��N�kKt��g��ځ~o_�K��q�j��37k�//�MwI`ht��p4J�Ğ�G]_�����l�[�M��Y�������-9���νW�jR��Y��tU=ͣ�E��!�mS��f��ӝ��ٳ?*��i�C��
LY~�輈��ʋ`M]P�8=
p���%��禂��8�Z�D�HŰ:�o�ޭ�[�?�P.E��1 ����;��m�^����^^��=�Խ���\���.��e��(�C>�z.�w.�2������*�V��ȓ�׫c]o^�B��7kW���0b�:�)��b��pwI�T#cL뫕ƅ!J}��:���i�ٵ��po����������=�`��bkg���OW��Qo�D\W�1,��J�L�¥^����?
{w�Do4�w0�Y��V��q�a0R,��>�����~s��I���j��K+�f�B��FX����8�G��q�!�fanv��Ϊ`��YɆk���>��
@��w�J�|s	�N�E�3�F/#��l�4^�塚�gM��O��dX#��@r!6�d\/Z��jnd\����n�R�m��bh&�؇2qA��(�;�]��>zc_�!��#����OD�ׯU
��s�j��U���q{d�g&��=�ct��f��v�[��.}�MƦD���z[�S^k��W��,P�ڶ�	J.+�:x�Z��{�T��&�"
���ූ_����x�=+�6�eZnx�@K�S㊅�s%�E�Yc�=>�3:�+�F�����s���-�m;�]F�^w	�2B)��C�E�]��w��I����
��ƹ��S�UzS��Q&����:Up�/�XzQ`p����4>?}���;?W�x����__���v��et�ބ�׺rB�����u��S#x�t
A�a�.���Bp}W2��Mb���{Z8�3*�K����;`I��7��Y����-�J&XU���P��\X���y	���P0��N���Ř�C\$��ڬ�3��(_):8�M��b�VD���Ad���T�|�R�����1%,X7l�S�)%Lԕ�s�y����2��*�E^ߟ.!�i��lYQiɪ��w/��,�L� �ǀ��m*ǝ�mt;�k�,2�H_Z�R�)�I�N�l7��CI;WH4Q9X��r������2�o����
<�(^ɑ>�⊍X�����S��j�B��7��j�3X4%��o���s�s��������%����E��mu�`���VtnMx!9ąF}�5m�)�]�tʥ��Pt��(���V$|�uH�J�vG�ux��F̷$�I[�Ht�	���ufG����qv��O�(�G�+r�)U���س�VҫaftǇ��@��̬Ԩb,�˻;��B֊-�t`�N�vmHOTE����,ޡ4��wT�7.^�:3I�qݴ�.��o�rʴ�&&euX�e^���Vb�S0��z�"G˸8Vq:y��<�Xm�,Kx�U�/w���C5V1J?`�(0
��w�A�&i� �N8\Ʋ=N^��;�4��c���;�N."oUn<̾�p/[h��
iw��:�;*\	`L*ݷ�훁ϓ��bۑV������-����A�y���~���:;M�2���t��%�˴���_�@mrlP��&_dj���M �j��>��(�K8�z� �A��j�vKɵ|.�C�k�v��f��j���M�AA��wm��ȼ��-&�T�]G�;��r�W����K�[��.��eqC+��^�V�����s��z�
�s[Í�ٯ*w-���*�j���\=���[��o���m����,C-_��W&*7�(b���9f+s.Y��A��&�h��޳��b�b��GrɆ.�k��@��(O`ʺ��ϕDn�0��'�+��ͮ|K�6���FT;3Tm\�Q:���-��&��`��핚T�&N�\�6�I�L��:Fc�Wv����ے�֤2�5y �N�fʾ�9��E<�����.�LO�A��ص�����R�u����n@�[\r�wyp���/wqB�r�ӯ��;I�gv-N�<'F>=N䍅�����U�r6����&����z�k���������7����ks:s\����5�u[�-*a$��5[u��2Uͨ���j�t�������~Mɖ��=�Ձn��_9*S8#7�乖i�-?�[�a����7S���H�e�շ�t#%��i`���V?��w7��>~]��l����'��gN�>@i9$5]ܗ�Em�rC��珏�����^�z��ׯ�_____����~��z����*��9��Ȩ�>D{�������}~?�^�x��ׯ_�����__����߰PWy�WT�����KnCs&��W��=�$�i�˖��kmA��j'������s`�y<���Z9h�N�t�C˖*4i��r���cb�m�.oyb�E4�bZthӪ""OS��hJ��<�yd��r]:4��b1>mG*�<�!�|��'���hh�J
y5�s�_��<�TK�X��Q�a�u^Z<�<��)H�`�΃��m)͹�,@|6N.p�%PR6��Rŭ���c�����AF��[�LF�<�ލMi�LPR���o*��yL�R	��d�-�6���	o��bbm Ẍ́nb&�7z4^D��T��N�$�[�:�� �Ȅ樍��Ź�V��>�}�T�.]X�@�A�fD�N���q@H�D�D���S�?���A�!%(�\4�r9�a&�1��!��B(� ���?��z=���y��%��0����pO���۳g`f#K0>���E���%�e�n�.ӄ�e!���>VWA�D�� ��5����;9�����^Y�4��Ę�a�z}n��'5�ȫY��T�#��b�ԟ<����0��{�^v/~��H�l��I�*�FEn����Alb�@��5��K'�PZd4�M���l�瞝�X0�k��Oq�h��P�W�'N�F��z`�d���ƯGAO�c ^�j���c=�q>���:ᚷZ���C3��h��p�]��h!N$CƼ��ɮ���pe�d�`Z4)\�,)����X�X��^.V�4�Y�!7�(2.��I�}p8Fܦ֠�	�x���-�owY�T��}S��ч)ƨ���e���@����?"����ozF�)L�C�����z�ا޻"[q2�~���'(P~��{���38k��.�#�)h3��F��]\�X�R�gN�.��t�YH7@������yO�τ|����&�Y����[���{���.��nAt�T/k�¨_J�9P����g\���!��!ÎՔ�c���n�e~���`s�ZÉd
��VN:|s�쓩�$����|D����VVjDZ���{by�C}e�?m(_ޚB�xɹ�=zZTx�C��UN�$�8�0+�q v���R�I�E�s1v�9�6��1 ������0h�z �����o5[[?=1��K����h2V���WE�,��4�u�����s�|�z9�e3�}Y�M����@0t�<Tku	��gۆ���:�=^���J=���[f2:IP<��_Q���!�5B�T��d` l�?��`�h��o"��.y�k������_5�HT������kj�ؗ��-#��!���3�����X>h���e�_��y��l����2٫H0ҋTIz�7k�0lk�[9y�x@����C�{a�چ�B��Z&9�k+:9��o$i�E�k�5�"���!���c��^)Ẳ2�W`sS+Z?���G�b�{ު��&s���T�cH��^Z���T7����Dm�n��wP���K�n�{T�R�t��k0��*3&�ؗf����c�t�ˠh%%�����D�뛫N�ߙ����'�#������O��zH����@>Xث*���^��)���L��S8��j����B�"Wx~�ѣ&$�/H����)v-X"*<CO(�붛3�"۞�^��:������\��DK�)=�����]�I��A<f�k7���Awd�h�3��ā��fPક�g��۹Q:]h�*�ˡ�]��~X^����G`-����M��4��Xz.���)�$�d��3�����=��|I#�&hT�8狫�7�dJ~����	��Z�_d�c˞.Jd�S�x�,���W�=�[O�D{�{;gFFn�Q�7�>�K��%�{���4���_8���OZ���˂��$�te�n�f\�XN:�2����]�oEM�d_��=��Ɩ�@��-A�6��A;�%Ȝ��ɳ�S ��0��	��6�@��ԝ�v��r^��$��]
����Tޑ}g��vn�������2��4:liDkO��T�0֑z����Q����f��5����1S����$n!|��>j�u��� V�� O��ޘ�R6eH}���8)	�1]6�WF7���5&LE`�������כ\��m��2�D˦|]9��j�٥�����}X��h'��!�9�G3����be��]�:��Wuv�f���hݡ��8}뢽߭.��ׄ�)���}��u�I��|�����'�C��u&��{XjA��x�v1\��{}��������	�8Jbv*����JX)	��	o>ލ�	�w��ozG^��\z��n����4�����ǟ7��&Ѳ��]8ƐQv�t�Z�t�u9�y���*J���rϳ�W�k�>�Tλ�͖g1�=Y��9���=j#b�_W2����???2� ���e�o?$�+���]�7�
0���[�W]��IT��Hl�8��jެC7u����I*�e��9,�@!g�=�/o�+mrB���;�=�}׊k����fm�1�~[`�֜�St�=��@�2D�{4ve_iF�FOor��Ѯ�띳�(��0�^D�ޚS�OZ�{2ni�
QB:޵��bԱ�-��Z"sst�f��~ �@�����|L��8R��L���Ԋ���R��,2�yU{�+N0�k�lޡ�t�i�Q*� �T�W2N㩸����^�����:��W���'���"8�~
wUj�}�F���=�� ��n�Ea���Mє�y��F��n/��6� �M���a���z�߭���웮w�u/��
,����ӑ�Ƅ��Vj�ϙ{��1ڷ��H'K�6�������]�m�O*��/���ۇ.�� �n�+�b]:k���t����q>R��}R����V�_ss�&���r�Ŕn��w9&�-�}�Ek�D7J��a�t v1Ȧ4�x3��1l�����m����iYc}ՄM���!���6�Z����~~~d  ���Nm{�	ǫ�c�p�s���v���K;*z�!��z>��1U9��J�ޓ+<j�}����o�gFQ���q�V7��9qy��+�#s�����u���d���mf�m��7q��d5�M��v+��C�<�wT�6�H�K��*��7<���h�x���f�vѦ>���H,��u]^��$�te������Q���ϑ�����Y,��Vy��Fz��C?�1���h�j���~9��
��u�вj�7�k�N�h��{�ϡ�C�ov����/�r�M��F����K�����z��*!.>m��=��zY������=�t�s[q�0�i�OW�t�B��QRR6��� TK������qכ۟�:�FYL������}�Ã�vz����x+�Q�^�;�4�a�!��i�������w�gb����4����[�/�V��m��S�I[JK0`��cmk�D��b��XE�:�3��C��c�̔�<Mۏ(��Y;�)�Qo?���\��p��Q�C�����4�96�;'�m#�.;��&e4R���q�d��1��y|�y�nlB�C��we*嶖�fȩUğ���g����@�{���3����R�u[�וA���n[���d��IfB[�w�eU�3j��3E���.ɚ�!�"�7IH�0��k�R7h9�L���v�4�s�p��Ǻ�.1��R�]��4���+K��T� V��Үe6蛩8���s�}������:;D��i+�fn��b�C>�`��3��x��Һ�
����W�3L��˕ygq���7�۱Ę�T�xF�U1�&(#��\�k��s֬9;"�VQ=Ԋ�6�.Lrל�p�]��`6��G��a����g$v�Ȫ�|pE��׬��'�fD�1�;�<;U����/B�|�*|V��x��ά{�����+s$�ׄ�Gh������g,�`B��O�6n����J)#�7E�n��$�s����|��C��w��s!�؉rVw���jT3�H�\���L�,D-Z�L"�w�x�R���[��f��t��Z+ʽ�<�6���,	[������
�.����/ ��g!�#��ΓgI�֌��d771���4nf���nu]���j7F�����x///{̒	 u}��ߪkaSl�&���v�>����3/FW�$`y4��JIy}��ٙ%�35=J��\!����a�$#�*��NP3��0�e]��(sMt1�rlݑ7��]ڟ\��쳂*�y�ұl��L�V�-l�l�7��O��j�g�&�������[?�5�O`90��J�g���񪷍�KKU	���v|^GI�&�	)W�G�z�ٝ�{�ht f�Ī�AdL�|�|�m�n'��[�w��a�#�8��o���N�h<�]H�v�_�	�����������i'�|x��3��۷���а]d>[�j���6�+|��(;�"4��*��GY؏Ou�W䒌��j�T�v�w[wUd@f��rn�Y���T�����g���SES����)�B9�T�2�3�H����l�;�#�;0��l�DG)䵐�kO�v��� ފXm�nt�4;�D��mȹmE4�!�V�z�m�%fh�r+=���w�
%�&��\2��h�K�]U�]ս��_!8E�G&w�q�ei�Y��+qVU�A|�?��FDGt�'E���)v�[u̖W��dws�אw������{��|O�}�!�:�+�,�r+h�����L��z�uw��9�o�F��-	*\��wwiD�+���<�l�yFh'�� �n�,�j=z��"�1��[�8o[�v��!�:Dp2�d�Ժ������WO��q�-U>����u^rx�,G��P0#�Y|�rG�"5a�\�̎,t���OמZL@_ �vI�q�|��~8Gj�}�W@~I<��qW]�&$M�0`�MQ�r���1���VWk˫��<{� �*�x55�0_2���Y��׼Ήm�n����'Ǎϑ�	�<�}r����@��{����3q�fZ�l���%��	@ȥ ��@�܊z�a�|����S����Vw3�;�r�&|�6.κ��4��AI�;W��646A����.����Q]��njc��˳]"9�h%Q��U��҇Ż:��ݭ�W���Tt,��A���;��[5q���3:e������c�e���<e:��ch�E;)�~j��=�}���]I��؊	��|ձNC�N��*�[l�Z���fѦ�ǩg�&����[$X�;/2R�������������I#�:��e��idgp�����WD����ܶ(��.�n )���~ճ�����~
sV^�F����ܸ���l��1N2���I���]kQ8d6c�۠���6=�s8��
ͮl�n�~����=���9��^�^����r[�=�e�.*f^��]���=U�z�Vwƣ��	���˱�4�-����T�wz�v�÷�kQ�r�Nz�q�e{�<����L/}gc3
�7w����N��m��4��=E�ex����mcR���`v�ʼ��0�}Rc�̽�� u�Ѐ�6�M�]@�ʠH��QR�3�]Z��ٵ�[ۚn�r�(��G��`R�s�K0g_Y�,�s��a�盟��ȭ���ix�/>�du1����|ΓD���5S��n������ot�ډ'|�Fi�r�]ދ����+F���}#�s�e6�9�x����������8��SI��l�_3vc�ؖWk۝���,��+ ���*\aL��j�N��~,]�cί)��x���ˣ���ҏ�h���)]:��hS�+��&�ki��{`m��Wa��ʋ�3F��.f���?����//!���t��J�3g~�S&�b]\G#<K�Uҝ�&u=-�":�v���G�aj�OIo�����={>Ax��2i%���t���fh3'�����bX"��DW��H��qbyߍ#�+F�W��f�I3�]�\Iզ�� �����ffN�<�W�\����2�HV fN7��$�7�Л�e���[yo���;W����l��r�vd
�W"'�+���t���K�#�Z&<N�i��W��+	���L�S��c���K(GGX֚��ݾl3� �46ǫ�;�u���&"Q���|zxo�l5o��)�������8�3�1�+Q������]�t��5���l6Ձ���Vg�����;z̖�D Q����F껏%��J�ޘf:�&���r���U*e�0�1C�]Qاۆ�99 ���T��%�T霝|v0�W\v�H��P�h�V��.�i����nG��PJ�P��0�[�8Qۈ��?6���,��=�(�}SU;!
��d�r�m{VkXX���a]�̔��θw�m���Y����-Ho��f��hP���)���o��w[�a�J=,���vJ6l�xD�]X{�J�$� X �n�-��!�K0LV	����
Y�\��`�\;z䡀�S�Ցĝ�VE�D����ѳM��]��ͫ������L��[u�����l�JRc�]���s�i�P��{l��u��oBn��Y���|���tXx�,����*���Ȣ�b�;3��FN����RQ����i����h��aQ��bg�v���pX��,o^��h�sr���B��8c�8yX��ev+7��f4
iLDҝ��'��O�2��\�Qp���9H]l9)EG�j�������<x�E�b��̧H��]]�"�{����#z��A�O;K�	����X��ɥ�f�}4�cs�͢���MZIuB7��i���c���y(ہ�j���:gG@2ngBp�I��ޣ�iŗ��u4v�sP{��h԰��:�5�j'+B��n>�t*ټ�W�r� 2l���;U�Dj�̫��j�"8B��sN4����Vz�0Vc�|��]G�b�B�b���pk��a�ި F��
E���=U����.��^��Z[��7ۧ �2��>��~>�i^\Ǹe�UhT�ņ�q��Iֺ��J䢊��r���{��D*���
�,Q�9�VU���7A�/q�5��Y�;�<*f��5��t�]����S})�I	]��}���Joa�4�/�]9��q���o�q�o���M<�o��� ��_Q�J�-�2C�mr�9,'lvs�����8M�9pS�ܥ���0
�8ʝ�j�̮�0�[�3X���|35դ�*݈kp��-V��p���x�b��igM�ik�և�G��9�]�=���5�*	-t�9��S�v5���y��5��ǅ���ѷ�Tpl�Qj1�l�=5	��0�	�Q�iUٛ�Z�,"4�݌1�h��1�J��hݩhN
Ow���Y�UeZ��|�)�E�l��sk-�̚Z���f�w�+%*��ma��،�����MV8���-
�'2�eΗ:��e�3����=���R}y�X�7-76�	7d3�\;�Z9�.��\ke����� ����.��2M��۳b(�M
�'
e��$�}�{*��@u�����^�W)������No%��8���@��te��ͻ�*1�z�F�Չ�:��,6z�|�6ljt���R���u}�i�h`��W��cFh{���j�1�yoa�0F�%?��9�L���������랽z�������������~��b���֍:;�r�(4��A�j��rKtܤ�mb/6*��F8�(��3��������랽z��������ׯ�������(�ˠ���l֪&����@r������&�Z�y:'�<����.jѶCF�V�U.�1݂��y���1?!�-m���73�6�K��/+�/3ɋ��9����Q��U̜�y���F���9g�m�����EF܎CM<�.s��5I��:�lh+c[%��ɪ֋�s��Ѷ-c��Dyh���,�N�hѪ��+K����N,ZtQ�f�"��7#���{�W6�F���F^lZ�44TO�$�N�[<F}�5UU��آ"��Z�$�3Ph+T[����� �H�B$����	k�~�uߏ�a'G%c���(�я��6����]��J��PQ77S�A2��+�O��䚕]�h=�Z�*�@�W���������.x��W{:��zc�}mѾac��9#Wz��6��Wo�"��TѺ�w���rU�M��x��dq�>U��J�^��^F^f��	U���7���n&���WSY��$�׀�{M9�@� �U>扺�����/���-ѻyot��5~#�n��s:]�Q~���\x���g���2��F�Q�犎�́xz'�Ǥr�'O&�����--w���q�'�%�����V{{\E��@�����o
OT�35��L�t<R~�6f�[�gf4����ө��SǠS��0��nV����,A35�"����M
Ӽ���w��v�\߅[8@�Ȼ��D��-9u<����gpΈS���y�h$��)��w#i�	�xi���)6fL���]�֜3=͑g�	���Ҥv�HG�)�$�O���N���na��m�Une��G*�>aF���Lea8�|p֋L=��MC��<��e)6�N�%��t���^,��+(�WuE��]�w9�,p�'q<V��B]G_ge�N\ߧX�_���2��g�	J�n�=����$�'*��w���}������C0ٞ��V6t�pQ�p4���8Z=�%m�im���}k���&&vv��;:n��k:�,��}�^'�m���Z�Z�fݖz���[+L>��ѱ����y̌F�w�����Y��Gg��Q���𙋍�Ki�8�d��;�Z��]��hoK���b1l]L�T�u�5�5ǻ��bG�0����9�S��)>���e�qe4���;X<�'��e_y�*Jy��i/�(#��	��(t����N�[��;e;�N᝘�e�����Zi�^�]�Q#���;Ew9Q�<�k��Y{���}2٤Z^��</i]������;
�l�j�i��~Y��®��FX��.�d2WC�J��KnW���躪�Ӳ��'';5�ij�z'Ė�YJv)̌�{��g����Y~����b�R<�7x�-pOe�[,))�(]����Od�����ݝ��~~*\�����=o��7�,,�F��b�l�̜��Æ�w.�Dժ��b���.�R�ۘ��	��0��^c���ةE[w������3f����������>��y��~Ɇ|�~�{�j����Y�f"�	O��[÷��4:�3mM�(�g�k09#��ػ՗��5En���z�&).!e��J����#�2ni�hM�M9uUwLO�$Gv8�$B��-�WP��$��R�I�jȖ��1a�gok|y��zޥA�V�<3	-�����o���ZG9��3��A/�w��3s*zO5��*Z���s>��ϤDy �n��ѽ)&�O�L[��?_9�};�NM�e��rGs{�Q6d6c����m��Ј�����y�p,h��ř؝YД�E���|��S��.BaȯoNigf�i��뭎�ϯʳf}Zu��3�.���]�e��f��|m19zV���ѣ{!�7Yyސ"�����]w�W��e?��NV�en�3T�}���&��xMW��h;���>��f�?q��e�U�gB���W�����GJQ��Ҕ�$��s;%�R�6�[o�k�6 �����s�R���N�
A����%�����	%����_q��{x�u�щ�U�(^�v�f������G��=6�����;�VM���X��9u(J�l���{�?���oG1#i_?MA��1�{�́��G ,��rE�W�,�7�S&(��L�}I�Ʉ7�R�I|��pe���3����5ᯖ,�w�`Rh0׻��Q]��A�@$�g��(z�b0_C�I��SN���G-�6�i:�,����ӭܶ�=9Ѣ����:�z�r�O����9 �����@�����_/ �@P�	��Z�ok��9��d���y\f����r�UE��sP�,�C���z�M�<�0;o[����S�^)��mub7)G.V�m಼	@�fl���KS �**z���eUqت�vd��xL�����$"��#�K$ԍ抝�a��S�.c^ �^���d���K.�wfD�t�Ȃ@���3i��f]r�o�ߗA��a&�&�wȫ�g�J��]-T�Ff��E]�3�C\�[;p����70`��վF��|�H-��b�cV1��d"�.�S����fJ&rhԥ���������l��M�{z�
ɂ΀	�)3w��W9*�-�C>�0P��N��b��X���.`4O"v�r���Zۚ�3^@{x<˭���>�|���жwQc�Wd���A��gy�V�и�6�!i}����?�%�1P���8n�:`�����"��\l��Fhvg�I�K������vZQ���x� W]�op=�t~M0F�Gc_v�D%1����Kū�;��e��0���UOU{��7%*�,��`����a����W��H�Ҡ��l�訽�٨�98aQ�.��i����l���G3�F��®��f��?X�Ξث��k�f�	׍e�cdv�5�O�;��Y�#T3���K��'�/���/���M��
�FGd�b=�+�i�3��}�ΨfH���wY��θ�,�(k�n������uB$q,pL���1���n�����Q�Z^x���fDZ�������{0�G?Q��p�o����o����U����@�x��=ܚ�95娭�j��^��w���cMd%NR��M�x8^.t7����	�u�D$�{��?~Z;\�$���^v�|V����<�m](*��<b�ݴU�[�QQC1߶�^T���EٳE�ɧ�Iu"�7x����Whu[�1nWD��4���ϑ��>�/}�@�j����W�/�o��ƛ�R.i��@�^���t�iGNO�W-���%K�s��s���%B"Ҕ��ʭ���[:=rU��Z��8�e�{�7`��V����>=��IJ�Ҧګ>�S궑G�q��3�a�"���ot��B+x����t{�IT�}o9�fz�?�'4ٹ�0o�]
��Fd����ţٳ�#^�Rj�ʐ�ֹ!�{fW�a/ѭ2���?���U��g�E!��rDjپ� P����gK[�4��kɕ�S8���J�W'��oy�9�eKق:�'���:�\�i�ӻ[����xěΉ'vM� KS�4 �Uә���@}p�|s�{��5ҳ�8���Υ�_q]~Y�-SJ�b�S���7�'�sn�X����U��!��yW�����;�ϝ���x�!���G��9�m��2��2}��C�i���@��k$�����"��fA˕-��^V������Xe���U�Z�4s��wQ�ƾKA����������୛}������2��l����"�i��p�ؗ!����O%s*��xE���7��h�y�!�)���F�T��������W�r��XY�N������e1$���Lh�5���c�co'ר���#�o�7,l6��WQ���'�z�����h;~xVj-)�o6@�����>я8Ң�*y����b�u�f
R6)�F?��i����J�1����>n�?#�����X"a˥�3���
��@bȴz����s>�g��z�#24�]>�>�FŌ=��F���Er��F�H�O�mH���F�8�o��V��>�Z���q�ҝ��Z��J�B��H������9���O�o���^fA讑è؅s�(�Y�G�))u;3�vգѹ�սݼ�;}J�dU��s��EM϶80�\�Ds����Y��_7��.]LK2���=���D�}r��� �H@~
=9�oy��Y�c9�e�&�`^õU�iٚ�-����'�Q8d6>F�
���4���a7�66=}c����^qt�����`�[y$��.ғb��'��>G
0�#6�:�	��6�-EC��bЮ�Gv����=ܨ���C�����e��p71�����j�^`�I��w0%���������#����L�E-S���kETU�<�`��g���\� �Kx���ӈ��ە��&�ckTej��(�y.�]�����^�m͆˒�(ҕ+�%t�=WE�����7�	˺rS���@Ҁj��kߢ*�'���ԸN�0�a#Z�T	�w�j6�̬�z�_VQ=��w7���i�����a�û��T��A��|�p]�F�dm��乞.L��d�$����G�2 Kچ�òzC�X7�3y��p9灡ۺ��$��uM�f~~����i�?L�7��g$؈���ی1�7AS�K@:(�S�@�k��Z���2��&R����Gn�Z��)�����9]�)�0DN�w�^p;�I����R�&������l�΋�d���� %DO�\ UҜ����ݗ\m�f�0��������c��h4�+�|��S'��Y�x}���nؽ����~śQrwR]��ܦ'R�8���j����k��,B���ur���t�βS��eV��K����1r��mNi�\��V{9,�(��8�����_-o���,ޮ�����_�x///~��vs�U�y��U'�(Y��ݦ*�)��s�ֽa�yp�,*FE�yl���6���U�c��]�6ټ�6zv��ܪ�o̑�OL���R����N�ںh���cI/�/g�y⨆+J��	�rMP|�;��@���p���g��.���w3�G��́�H�\�R'|�[!���̯B�U.�"�#��ͧm�+,�ʟG�Nk�V�*=+���Z_d��X�p�"��#����y��w���@E�F6kQ���=�K��7����d�v{+�ͷ���Cg6S���oTAO���U��\��S��ө������/�[�-�vOQRo`t���̀�|WP��>���կ�,hu9`��~}�;�$��$q�����J�����n�my���Q�T1]w���w;:�3��4��&��wx�r�6y�;�i����087��z����=��Ҟ�NF�n�]���D΄ƻww�#(2�Ht�C&b�zp�#:�yN$:��e9���o-t��i���㐙���-�'.���+��JB�:	��yhv;�	`u/!��m�z�
r�qm<�=�<ơ�".{����3�������;�8i�S�i�lU��bF�L����1��F�sU�R���5�jۜ�U����@x4y�sm��D��N��h������Ss^+R�W����v�~d"Uy�n�_�x���癆g���{�'�θw��e���g\�v&�{fGE<{a�w �Бy���X햭�R�Q"è?N����W.(
�|h$u�ٷ�sNv��PF�~�I9���k��:�Z�6I��$vWrJ��*�#rv�@4ә�[8��{eOu9��쁻�Z�Wpqz,�%�����Z��OB�JFUO�r6=N�2���6�wb;��]��
�ʸ���	 ]u��	%%�ͪW6TYUݵ���ٺ��O���M�nL���}~S|Zܔ��V��V�S�KU�n���gtyY͟u�K&��n���d�ճ}|+�}�,p���?p:����CL�d�H���ї`����,�}��˙aJ���3�v��//�pIp@а�]_n�[�(u��Mx��L�_8y�3U"�)�u�����a'k��.��������&Rf�����ν�/hh��ELN9ϭ�����vl�B#����.ѡ�d�S`���'*5�8L����]}�qf��@������utsU܀����-p�o8a�i��×�}�j$*o:�-�4� �{Oi!ncG�H?���}��C�1m�S��{;��xC�J�Ft�<q�އM��ďS�,R�֠��o^�u(�w���vOc;��Ѽ��ƥ�Ө�ͻ�þ��k1�)�t4�+�Z:�j�����r��rH�jU�k�zv��05�Ƭ�8�/:��)�A��q����I�:�B���P���j��9�U.��#;�]��tNnK��of*�"3Ud4t�ӂE��AI匃2��Rm�o1�����ͬ�������ٜ��M|Q
��=P�ښ���3s�hs3�6[!L�e��FV�Sŗ5I�sTxC��z�s����
᳈ǒ��y�"0�A��:�pw'��_ch��s��U���\����E�e����wu� V����Hq�gv�iD�QO��Ê��NZ�ܞ@���+���k⤩y�[݋(vʈ��]Q��E������q�N��m�
|ݷq��V�
��A��l x~�xǤ�V[_J� o5W� �~�9r���̝�H���s���`U�oh7"8F�����ȹ��ZpmJ���#bO�{#U~j�^�*&�A_㗕5�X.�՘@#�wm��)�d`�MCs�W	D;p'r
We3��-�V&��Ote(zs��B!�qz�H���|�c��aA2�[�J�l������vq��`�$<�g�-d�v�a$�'�fd�x���FpC;^u��nq�N��n���3VC�9�Z�fQ��Mc4N�ެ1�A�����0���P��V;j�:����}��l�6�x���'^���&�q�j��U��]�yX!b���8`l��];�9��ܝ\�\�۾2�wmuI2t�Uu�%��)����
�hK��0)��*D/�u�\�����7���7oU\]����l�\�e��uj��j��p���rڸY�@ĳ}Q%�0ΗzU�:�2�,��S��su��|;��D�cY��22k>���樔�Mt�s��&���-Ìl��˘�#�]�]�]�>N���E"-�I)R�v���B.ԲG@�-�Gp�b�n�"Ә�������Bۧ�+�X�(�{l΋�.|މ׫8`�y�.�3Bw^��m��f8��D`���54i�\0R��;de��1]��r^f��Ǳ���ϟ�����;l�$ME4S^��r�E�gi*$���m�s9��������Y�ׯ^�}}}}}}z�7���қ���l�4cjs$AF�k$EU�֯�r�؊(孱���O6*os�'Ǐ���������z��������ׯ_�ס�*��Ѧ ��m�}ڮ��j������ocMSh1hqV�UTEQ3QD�T���ɚ���TE{8� ���.m%�X�50�Q3����"��٣�UD�ƀ�v�UAQA2L�����"v1i�2i0���ѱ�h4y�i����<�LQbϳ���HQL�m��5TUP�fovj&���|�<��堢�Z�mT��L�DL�%DDD�D��`�d���O9�"��e�a���`��61�U��i2�3Z)��m��`����h����1MQF�TI6�J��ӈ�`���6�>m�Q4��4S�ˈ�h�O��-"�&(aq�iA<���8)��(��p��L(�L����gi��5������|�<!Hٕ��#1䦴��3ְom멇��ո����=�z�	q�`a�	O�D(Jb&�m�$m�$R(�$�Jb�	5!��E�����uP��Q��I"B����)�	,(\0��\E�;�߼�>g�e,W�&��W�{�����8�W&�e��o�QJ�<5��L\�y5p�t�nWb(���>Fc��Wye?�r���C�5���F�m����#�T��ff2�n4�� ������oW�oB�����Gug%��b��}o���L���Uܖ�D��
�t����w �/*��Ȼ�ZZ�Cp��/S�������t���q��x���3le��v���7����4�d,kp&�l�q�[&�-���Ԉ�	��\�M�`�H]����h3㳍�`E�YzKs^�B�1�M��(ͪ|=��:��y�;��I-��O����a/}p���rj�ͽ�	aݺ�1�����谔J�%Zȴ
�S�Nr�> ��̳��(�ݪ�ו�� @`�����\�>�=�)�5���ͥR�}��#"�Ed����:��JYP��ʯv%"��Ai�xR�'��hw!�F-�ܳ�_ _�ƶލ+��b��`5У���.����rͥ�Ӓ��(S�Wش�O�L�]?ΐ$a��lڥ����vr!��Fq`��u�&lgR���cr�3[*�^�^�n�̏gr�u��X;M*��7y^~�����L=n��QSP����j=Bȃ�qEB��9h��P
�O],0��6w��4��ʩ���}
�N�R/x@�e��F��x՚�Φ�n�x���g���*�䧃���U*���r!�2��N���3�D�>kS�$Ih���!��*�t�IBX�6cǶ��b��˻�y��Y׭�my�|��a�17�d^��)�G̶<��'�S�{����'%��%%�v���m�Yc�>�ك5�f�kϺ�3A.���
��Jܨɬ��v�C3O�R]�`M�0����'_�껒�+�n�Y�/9|�g
�����8l�I�`���8�oC���ی�I���q}Y��U�����=,I]�z��� �d��<���.n�p@Y�r�fc��8����K�E�:�'=�c����xhR>Wn��fT�CM�����ЗO�{�B��k:�cO��[����:��LL�P�_�mv�7�Rd;R��K{\�Yza8(���7j_�EI{���9�m;P�����3�.��e�$����w���Ga��ͧ� �G����tP��J��P�������wݢL��ó�g��i�HtZ�'���i�<IhE�c�P5�\O3�\s���a��|^j�^(��>�<$Di�崹�ʍIDT^m�0��M�s] �����h{�ͿM��`���:R�%.8��h��6���y��z�YT�K���,~�s�znj%�|���3"�H���Ѷ[��+(r<�yn ��3���+�,Af�T���m������Cv6���1�+N���hA�T�et���y�=aAY�y�
�"ڢ�SM�s�6l�r$ߘ�T�R�^�ܙܷ]��Eջz�p�ɓx��g��ʏB
+�G�T�Hߛ�*��>H�k&��:3�پ���;�{�2��[n��g�"��H�`R�5��[<����Q�����0�F������n�uQ�!�� `W���T���kQ��=�rR[��`�
��R���>�v������]��h<ld��������wz�κ�7ӕs���>�=��ը���=�jS�jl�X����%���U�Ӽ�3w$��m��M���U��D^X�N�ѵ�"�D�4(��u6�봞�����{M�ga���'Uv:.ո�a�,�սQ>����&��j����n�ݔ�7�2Vv��n�7��|�Flv����v�Rv/�s#�ڸ�1��H~���'���] �l��ǟ�}^}��'��V'��}��ꃯ�Ǯ�ks��k���&Mϊ۞(�~�<�ݝ�l�a���]� ��f�w���:�X�J<�l�6����d�~�b;������9a�i̚˾��枅.UC81ȵޘ�uQV�n��yo��"w�_=�Nϛ�e="ok�
�k�&�\ϭg��hnCں�*�݀/���tVv;U4�Ѯ͚5��Y�ܛ@��#���8��$�pl~`c7SuN-i�ٶ��������p�J�2�k�YsNge�
z���/��Nb;�n7�����y���J�)T!+�w�{������6�dm��"�G�����-��ޜ���Sw�qb�K��E��6�2��n�K��hzp�ᶜK���q�)Ξ��V��wdK]��Զ9o1Z�ܦ���-���.l��-l�ma�e[@�y57���v�'�H���g��G��X/�
�R?���o�W]��۬�Vh�R,�Y��n֑ʖ����3�������a/�sh8zR0� ���u�K����I���.�x�
����@��q��I�xb����@�e-�ٝ[�K�*���q�_����W(�sx����1�N����Q�w2�e�l���Wc&�jtp���j�S���E��a�^N~�VY�VO��'�'���$L��>��D�nu��᭦1�k����d%y�7�����%>�&��bB��N�\e�n3����H����Y������i��q|dD-��Rv���ԉ��O�7>�O�nm�̯wu��iU�8c��f:��2⳩S�/qm���'x��z��m�:�p��s�P�`�5:�}�"��-�z������훃����Ս��ئ�A�tJ�u|vt;�`F³@E�#0c�͞�\3?g�g����4R]���V���q+�:���H�s,����Y�ۧ��������f��b&�v��.-���&�k\�"����=�%x��iڏC�'X����V�k7|��}���$��_s�cy��ɌN�n�h���7[���!}�&�S��%j��;����}4J4U�<���Z���K8���#p=�F�����q�V�Q��[pO�/��eH�f��.�^�t����P�e���LA�0-k�U�G�t����D�d
Q��.�IJv���u�\�l{�GՆ|t��|j�t�(B����EB��q�e��R��t�9�n+����c_�)v+wg�!S��g
cU�E^�����fj����C�S����U��h�����]R�F����0�E�� �R�U�r�ɽ� D�{��a�q����f=�m�
��3��٪��st�s��0E� ��|�֪��(�\����|�W��Oss�j���'Wu��	��S�":6kTȭZ�eKu.ǭHt���X{���L*�M~����\�#n��hK��̀HH��<��S.�a�&��/Yw�t%���鯓��(�Ӳ��X.�볬",��"|t�fJ�W5�R�\�X$��z62rrIݵv��iom�Wj�vN�]�|ܚn���N���LŘ���bK8D������N�d��₃0j�7����ǘ}�x����ޮ��^�N澷kM���6���<^,��UR���~o�7�^d�cn=�[��NL��`ͪ�ޚ���
�r�Vv��gc��d6�`�(y�� ���� -c(`�[�C{muFE��Gt���g�l��M�H;fEg�9��\��P�0Y�LMus�\r�qݙ�٧I#�6�ڐGH�g���D�~� ϦoYo��s�l��9�fvT�]ǃƩ��Hȼ����:(������?+�����i��o��1ުU�V��	=�Eľ��a5B��!* ����0�����]p�W�*k�G,ra�XǠ�w������.j%���0K����&����׆h�8T�%�˪�%��g+�X�w�T��yw��'�����ߚ������L�2\�|:i�i� I��a�z�Z��Mg�Q�fM���L[o�m�����ˆ�"��+K4L�U�f�ٝ���m�tWS#�Ces�ȪX�+����XZ;g�;��h����Х_[�am��[wE��1_R��h�-�ٺݓ~����Wq��ߙ�~�|��l\M��%Ię��S�n��+6�^u,�g���Ӫ�C@��=
7ϡ�P�[�3`�9"��g�-��妭�v���8i���w5�̺[�4v@tz�^�6<,+��V�*�q��m���?ڙ��+of�Ste>����3c��!�����1���k}�L@�峚�U(r{�����l�j�p�'�.�(m����[�{=S�$P��z"��L^3Meou��<t����q�
�d����I��v���u:s�V��ȩǾ�XF=;�)�+�����>Y`��V��N�Suk��4��b�C����^/a�T]bY���^�]���W�oݽ�7��.�
�b�o�t6e�@q,��ɝZ��k�D�&L�M�`���c�]���=�Rlޜ~١<E+|�l3�\h�
�EZ5�4��绉� �f�7.�U���ڲ�����H�.��*&��L�H��ej����#���(u n}3�s��8�)��n��g��u�����Wu݊ ��l�%��]������/X&�ޮ�2f��p>b-�
��j��|�j�x0�٥����J�����4��S��Q����w�8�C"˗i2R�r��~����m0�#Uk��老�4=$�Q����F�Ϗ�,����L�y����ɤ^ڞ�)�X�;� �]��.�q٫�Ncf��t�GӍ�d�@�+K�(+�9�%���Ĺ��t;�l���6�`��ͽn�<ø����â� V����"��^��+n�T�Ag(nV�{Nk�b.������p���v�n;�{�'�˧����.�JT!%O�l�����t��k��I�l��@@\�+����z@�-���$]`�ܨ�Ջb�M^�Nr��}>k��^�#`����W�>�Fz�f�P
M����j�l�RC����&Vv�u��������X�۾qr�n�\)N��0�͞�~�ؐ;���S��=���=��`nq;yY>W/�*��3=���`���+�3ܺe��)�k۴<q\� c���t@�vce�U��ߟ��)�_^�ԲS����_�)љo�B�)!��c+�L^tA���LQ�M�	�Zb�&/>_lEJJAcJ��E���dd��#;u���%N'#�r�nN�@��dAn�iC�����x�^y�H�l��}��z�6�'x,��n���	7���;Dl�}���Kk�SAWL^��b�y�����D��Rz�P(�a�#02�?9j~�?b��;R9��<K2aSlC6���o����aT�2 +��gϕz�3������5J/���C�WH����wG�#
�E�tkS��(ǵ����<�A�Q �28��<���)η�#�� 2WJ�g��ֻ�j8�e��u�.�y1��z<�F'u�E�<�@��`��O,N����=����Y�N3�Z��U��
��}s�!>�Cd�F��g��.Ѫb���K�{����MS���/U�vY�+�������j��XK�.!?�x=,�=��Ӿn��Z.��t^�7t��>ݡ�W"�
��u����T�᱙�4����.X�Ͷp�:�u�o%���Οa3�Д�]��SV�B�sS�EK���MQu�4o�7G�p�3Fm�].}���*�:�E���d�B�(�y�M�!��Q�@P<yQ�]��関ڣ�����A�+]��oy+�:��-yu��]t��W<��7|��z��[s*Y�g]�̣ηR*]v�
��k�����l���p�.�N�:#����˘B�o7��J��D�'^R�h(A�x�;e�;F��"V��'y��c�p�:{�ਜ਼r�ι����uJ�6�ELW�`6��9E�kʾW�ڝ�IR�5c�뜲�:�lhT��=��]z�z�X�r�YttKݣ��{P��o�S��9@F\㴣M�l���v�#�!ԯ�`�Y�'[vf��ԟ+eAD,���w]0�v�Z�-у�&���2
u�J�I-�^�6fY`��}2����[PoR�h��J�;�7�]��7��L��0<|�v�ޙk��
�=v��@�.s�zƞ��kw��L�k�޵�J�b��S;N�ڵld�,��M�e��:4�t�cip�V�N�h緷.|�� �Rc9}87�;yɡ�l1v�6q&��E� R��Y�+n�'R�M���]�2l�JN�L|i�]2�:�Ly�u���c@9�a��W�k3�5M�jLtV��@�M#� ��8$Hp�Uɉ�۟䀾W��]���e��]�T4vK��Ȏ�.���ui����ĳ4�>��'��#�P*�4ɸ�R
4qVl���|R�)��lʝl�V�wYtڍ�p竰!DY6��BAUs��VP�I�Z��ܧ���ټ�����i�V3u%.�H
�}��{9��j)7��u���d�n[��&�=�{2��� �J�jP�F��ݚ�v!��v�L&�Zy*X�/��lݻ�^��x.��؏��mP=�2��\	:f�((�n"N��f� �`veq����~�()r�9%�I'�Dm���p�Ŵ��3�
v��\��+��V��J�	��m�r�=��wsf�4��t�٢5�p�u�x"�@�÷�֪ӆ�}+ng�˦�ە�ûZzEs�
��BUӝ/e��	H](����݋(�IK���Ïs�(����=��o8����I2�������"��O��6{��"��Z���o��v���a鴅g)��L��{�	vqvΓ��T��ʑڽ7�f�fi�Sy?�^{�������\���#u��Rt�Պ�l��$6U��/��&��9lb�p����k��ī��5-�vzB�V�0����d���o}վ��znA�R�P�����t�w#;��$�L3ܢ^i<YH�u7X�&S3Xn�j��+�yY����Y/q,��;/��$���"�ƌ{���2�:�S��
6���-�9�9��0��pK��!Vk��x�0�N�Q���r7mZ�2�^mT�婈�+gU�-��PT^Z�{�T'�3�ح&ƫ�s�^�\��b�'<|}~?������z��������ׯ_��{�j��"�+�5Ec\�(���0`���h�b*���AElm6����5�fs������z�z��ׯ______^�z�~�+��1kVƨ-�i���E_q��
X����&�����
��s�ܩ������*`�*�-T�r�QQ��((*�l�1�5�h�E�W<�ɨ��&g��y�l�3��Š������Y�)�3���<�RPS-�A��E{yr[X���"	��51��\�,6�r����b
	���Dy�G1� $�"���"fk\�.s�-4QLUr6ڋmDLhu�@�9QQD�Q�I���gL�y`�<��!���"yj%�NQSIO,Lkr9� ��`��3�b�� ��<�r96��劼� �77"*h���EE4%SCG5d�cks������#�RT�m��J�Z����;�y�)��lf�b�J9cX����glD5��C(�|H4@F$I �� ��}�q�,*�V"+-c�0��M40���9���W	�;��z�[8�h��lbnvYqX���͚�߿}_�zY̘�1q0=�4����IU?\�u��m��$2���Wpތ��{˝�v�Y����9�����$����񷌶y����\�G$�7&��w3��=��QD�&�l��=���VmP֨w���j��f����Ϡ�N���5��T/�<�z���"OVT��Ή��ܾ&�	v�@�k�2fϞ8Ȉ�1����q����0���4:���'tׯ>����L+���ò�dF�cJ�M44N�;�lE�v�&/���8�Q��Ѵc|�C3Ok0M/��Gl�\C-�$H9���3�zM��<[ah����mK4=�-Խx�xߌ�r?�^r�J���U���F��1w��=��;=���[�X�}LF�RӢ/��mu��玘c�E�l<.��D������DHKDi�����o�⻵}]t�3��4p�撾"c۬T2�V@v"Pe��~��ш�#�1yC������ʼ7�l��r�M�\��vՔ�q�5܀��U�ի�V�t(���}�����D}���,5�ϑ��8��ʺ��Q��>o7Et^�n�=X�-�t0�b<�ٗ�F��d����_U��ʹz���z�������E[�>�B0׃�P�S�Y��:b��Z�������H� �j�A#�z��\��B/Ӝ�+'��L��f����[��x�v?u�W(�K�qO9+ģD��A�D��D�?�/��*,눦���u�Ndt-m�0H����7�HlH��#@$SW�DnV�:�QE��!��NUޞ�ΛH!��{0O}��o@̈́��䊾y2�0�i�s��b��4�����!�;��u��D,��� ��S�*�z��輮D�+{u�1����8!��5�獳x�z�>���Pir
�~�Q}��k�5{��4K��*x*����Gh�>:_����cZ��9�n@}[�A]�c��^h���V9vE馽:[�u^$���!V�����0r6���j��:�T��U��mA���
��fd�q�(֍q�J�5:5lv;gU�-.ױO������b9N�����7�vu�;o�!�@K\.�1j�Yk�]b���5�ܾh��(�����+���'�W
֘a��o���kxo�|���݋��y� ���k������ʩ�D���'�QU�O��
{3����ΥA��=�({�XU��ճ���x�W|�XsS\L�"������u���7��9#A?M�]#�c�ٚ2�d@t�����}RL��g�T���_8��[]�"h�$ω��/"Xi(�e�d�U��*�\�R:���ez}Qo����ܭِ��}EI)8/�=��+�:�#@>8��1��pTk���3�!e�ҿ97"��k+�9����zK�3��?q�$q��{jz)�a��;���ɝ
�2fۻju��ޓu��:a��ab�o��dtR�l���4�a�4UE�Ӌy��"c� f�δ�\��u��╁��:5�;w�"�oޙ{�<M�M@�YhW ,��F�"�n�B�$�s6[zTC:`n(�ȍ��s�UD�14� +��O�(�"+x�����{�w���r�W�J7�^�qn��o�㡱�r�s�dW��s��3Ͷ27�,(�"�E��S��G�';F�,㼾�1���P�u}Rɐ�.�����;�����Ο3Wm�I�N��&��fW�dP
��?����Ӑ۲�9�;t�����7�ё�s���r�w��V׉��>�������:+hOL+�L�ɦȪ�*�U��f���C=1=:�[���t��������t5�b[�ÑI�p�U'q��v�`��9U��Yؐ;�ԵbXd.O���m�ZL(��ߥt��ѽl:څ�~dr��F�F;��Iݟ\@�&��=D��5%1���r���㔇y�M��R���ܖ�Dԩf��-Z�O�.ͱ��f����5I�F���=遪d@ˊΥO�y�P�����UnU��5��2�@`�㻺B�!�����,�}�0�Y>HD;���^;:��3[ĺ�<�m��v�h��:�8�g�#�c��Y�w~9-n���j{5�~z�CPسD�����u�˹�JF�<x��� �b�Wm@��7[a�]jʊ{��Uщ�$�Hr�5��b����߸ٍ; [�Ϭ��������o>�I:�Z�(�Y�wil�6��z�]��yǸ�.�s%�ʶ�p짘te����"�kgjcOa���td=|�:��-g	�b���`�)E]Yɦ�8�f���Z�����&���y��ȫ����tmg��w�>���B6:Em��zk��e.]��xt�.���l@��'���z��1�iǬqk��+&������<J�q6޾b\��2l�N�ܽV��"�P�P~^̔b�حԈ���C�0{�����b�ޕ�䔪��;w��Mc��9��A�d�B��b�6�sN�`A�2\�9�h�P)BQ��G<�]D'�`��zAǈ�U5�{�Վ�O6@.A��z�=;ԕ�r�\�Q$��'㷱�1���O�y�ums�V���9�6)�8���F�I���'�
����3&��wG[VVe���<������T�&�o��9�"Ȉ�NНSZ����ty��XxřI�-&_��� 5q����m��Ͷ̬�F)�5F%W~�4!��'�]��?b[��2��ﶘg��F��ۚ����h��e���W��p,(rY�SW���òs$^�;Y��<$��o	>�S���ߔ���a�A�vm�M�M)r���<m;�� �����.F��}/GgcV'B�m:/��]B�I��۝������>���Ks���h������{��{{j�u�Xn�W�|B�e��:�r�U��^�^JBŲ�]E�Ux�� �;&��`l3��g�!�j{V�����pϥ���]P��(��z̎���p�>��tQ��5��ˁ��Fa-�-�a�X@<j|��C�#B�/�=�xC\F��˺�i�����¯�qf*-�F�	�
-v��ɪ�����:v#Ii�����ҏg^t�^P��<+��K�]��n�g�I����g�ᛒ�e8)�2*�S�:㬋�EAԎ4���\�kC|�}�^;2�~b��^�M�c�7�@�ݑ��<v�.��R�Ч���3C�{���=�[�~��!Z��م�=HN,��Ȑ]����j�-5^��&��O+�6��bo	 Mxy��*90B��+z���rEsF̄:�3�d[��MM���T�͔&)�皶��3i5���ɽ\.�B��Wa��cGz^K	W�;�����T�	��-��b;��Wo-�����<=ǰ�{s3��N��;�v�R���W3Hot�[�Xj��;�uACzԤ����}������������c�y>��a�W��*��Б�7���ҧ�y������6��­李DQvjQlո*�9�0�ƛ���]t���v;Xk��޹B�Fjh��OFg�?��T�:���=�m��t�%�'H�Cn6{C3y�ս�3�J�;W����뺳i{wTwS�����O�!����5������DS�;3�7�ΘK�����Yݻ%yWA�u�KuԻ����v*��Ä�������X��W�W�'��F0��R�b���5���?M)*�;��	��8w.�%WOu�� ��^x�9��c�Ц3[�:��\؁��-�j�������:�qV��5�U�u�'$����׻��'.�i�!����J@��r�pT{^_��� beޒ���ݴ���OsT�C_�͛�f��d�$i��y�3f,�ǀ:Ń�g��I��my˼?�3K��-��?؎T;~�L��x�ƺ�m�SP�)�X�6^#H� �E��i�m��a,3A�k"��W0�˗7�;��~����1M�ƏLL%�k+q朴�|�])��N�����T4�d������9i��kN�����軽,q�0�^Y7P�r���Ko�\tR�l���^ɷB��y����am���=u�7���(:x�V��E��E���"-)T!11n�,�/1]������DT�BqV�7}�v�C��d@�[:��Э��EH��o����4l�˵(Aͮ~�Ψ�g�q�eʏ)�@�d�I�l��T��Q�βc*�l�X�]'	T��ucY������M=<2pF+0������z'O��VyF�t�Y�#��X�ǚ�A�cX�>[=��bn�U�,4N	+Nd��+W$L�.O�<��km�7a�I����Я�ZtWC� ����z��Y�o�0	ݓk�T��|�"1vgf����^U������N�)��ݮ����~���;������&�̼|JQ��̙�O��� �+�G�oCy���@]�T?����C�r?ojJ�M��8wV\��@�m��&^��@�%�%�E3ԟ���Qɪpe>B��k{�׬+:�{���S��uTk8J���2�2��q���`����J��ʍ^T�r�����T��M(3ys��qw�ge��D�Y�|}������wX�����	��J�)ѥ��`>ِ J�둹+��M�WԱ#=�O⿈�������b��6�������Ɠ�n!؃�y�4�ON�m#9��ٍ I��f���ùXǆ�h�dlS�;Dѽ�4�nw���N����:ԫ�W&���U�D��IT��-Y)��"""�W�WԿn�'7ʺ�a,���`����5Q4#����rB�&WCE�۫l�xc�sz���w˾�m���(+���RN��\B�t��
�-*1�{w��=Wyx�f��,������G*��̋jsb�yP(G\��/����먊�S8o��9U��jA)F�R�Ќώ���n���x<��R.n�e�Y����8a(����g���{A*�$��GG�|;-�z}���M�pQ��yf�oS�}�������hޒ��.4�= ˉ�����J��W������*k:���X�Fs��
l�xH�4����ש�n��(�Zk^8r��D�k��� �l�����e�ޜ���Iv�̴�GC�k���ܗ�&�(y�E�i���;����Ȉ�����������{��_w�R�@��0�9��"��N��%F���nV����&�g���z=�5��c)�0r�Kt5����������K����3+%�-Ko�
%�U��$g�v�k�Z2�\j#��\��w�0�\�L�S���������7��e��:�>��!xuB��w�4ܫ��;��e�B�)��
Y}O�{�j��uCN�mf�m��a�B���e��Y���;+���VھK�A��`�� ���g�A�cfq��1s���ò������^���[ota��gf�ۛȹ/+6�c��	�S^;N��xJ���ߓK6����i��O��پꜦ�g%{BӍ m��3��xQk�pGz�i�3<Cj�ʶ=.ԛ{&y�6x։:��jL�2"�D�{�w����������V��p
�+��(����{�g��( ��dU ��Ä�������QC2�0��C�2�0��C*��0! �2�2� C
�(�2 @�0���Cʰ�2�� �0 Cʰ�0�2��ʰ�0 C*�
�ʰ� C ʰȄ2� C ʰ�0� °�0��C �0��C 0C*�(ʰ�0���C"0�2��C*�(�2 C(°2�0�����Cʰʰ��}�� �0ʰ�2�0,0,0�C(2�2�0� C*�*�"°�2�>�2��C
�"ʰʰ�2�0�*� °2�2�2�0��+ C(ʰʰ�2���&F��DĘaeddXd`Xah`ddXddd`Xad`�$Xa`ddXa`ddX`Faa� 6G" C C C( C" C C" C #�p��� �� ȀȀȠ� ȀȀ��.�``P	�e	�@�@�`T	��PBi�P&&�8<&&A@��DBI�Dd��Q�Pd�pC(��0!M0!�M2��LL�����2�2�0�� Cʰ�2���XeVV@� !�aXeXeC�w��� ������Q�	�QQi��Ͽ������������������@����8��.p?Л�?��������?���ETW�������PE�_�J��������!�������)�O�����C�⊨����!�����Iw���O���a��O� ���C��د�a dPfEU
AP( �@ ���@� "E@��E�" D�� @ ��,�)" B� $� �    )" J��(� �( B�(B�
�#*���,�BJ���$��$+$�A(
Ш���y�����O�(
*4�
B���?����o��XP/�hx@�A��_���+�����������?�?R?���c���������O横���C���?�?eTW�UE؇�����C����<8
�����:*�+� 3������C��O������o�����O�����zQ[�?�i�C���C�w�Q_���i����?��;�X?��O�<��?�?�������?q**��?~�?����ETW����x~�y������'���?����?������O�Г��=TUE}O��?��L����?������_�����j��/�����8���*�����?���o��O��(+$�k&�r��96�0
 ��d��H�>v=P����MP��-�*B�h�IR֨V�֩KlJ��TP$�(�	يQf�R��5��B��R(U*�Z�B���kOn�4�����%�-��֪��Ӹ���j��l����4)�-����Z�F����km*��mI��(�fڶ,�jڶ�df�Ģ�ZW3P�[`��A�2�̖�V*�,�kY4��Sc*%�l��#lQ��S@6V��Tkbl��Sf�-F����l�l�m^��,�1dfh�w9�I։;Q�   ��wcJӭ6��vU˚�)�k��u�n��<8봪�t�:�v�ҥR�wa.�wj��t��뚮덻�ۗB��wX��c׋�)+�6Y5kVle5b��m��  ^�E��Q}��
8�a�D�(P�C��<�$>��CT��mxz>��h+���Vw*��{��v7eS���˴�p���m�t�.�U۲]�:�(v��*�T;�Zuۭj*��Ͱ�m5����)���  {�4��s��`S�s[n�ݪ'p���mea����p���
;�)�;p��.���6ڃ����v��GRUΎ�c��[��j��$M�Yl���6ڧ�  ;�C^��7:�����4p�j���JjM�
��z��m���MD� �J��PjCKu���ֵ[�8PwRɶ��յ�V�lmhd�cP�  �V���i0֝-��::tJ��B�;��jͬ�����Eu�M\�Ӡ��QT�N�Z��w���嵕Z�-�e�j�IJ6��   � u�ݪ7t���Ӫ�ޏ]:tRkv�V؁��wM��ָ*ݧ�)��+������k�"� ��&���%l�j�l[f�|   ��(��ҽ�Q�5�n�m�F��A�WuI �W�t�D������=�Ǽm��RyåE�����)+P�)D����V6-b�6I�>   �R�AKܣ��JV��r����]���m�OWz�J����JTUR/x7Im [ԭ�*Q֋�z��]��)�o��IH{.�MV�a�;��m ��o�  �ϨJ�Z����B�Sp�q%����W)J��އ8P�d�;���T���n]�{iT��zw����03T��O����%���-��j3�-��i�Uo�  ���$JW|��z5�fP<�(��)�xs�%J�oJ�(*�*��e�zERmz�8�f�I{�Υ4��p� J�D����4ԗ��O��)P  "��b��(����JUL��  "��4��@  S�h��UJ@ he)!��� '������_�F�����{&=����T`�-�u/��6<�1.���K��}�W��}���.��l���0m����C`�6�����l���������������Zy���uw
�)�,.�|��M�&�+UϝE�$�kv��N��G�[�V�z�ꆯj:�n��3X/R�N8�\ǂ2Zp���x��,e�q"k~�&�J^�cVښ؛�[�!Rڴ%�K��Nd���,M?��t֬Ƕ6���j�d%
ԶL�䲎E�Yb��M����T�gfh5u�!��[�iwy��n�Ys35�W�!t�-WFċ`��P��sq�8 �����(P�X>�&�ӥecn���j�kcљq�%sV�#X�"��t1o�vn(PV�[ͻV��o@, .�m����La�Osp�{$�N�k��Rᇂ4�����K,�
�y�gn��R���	�\�9=��Vm���V
(0ZT�23�Z�SЀ�&��/f�vM:qJ[�JQ�Ky�j�:�Z��x��`����P����olfʷu�n,.,0Px���[ѥ�H-����Cmbѓ�M�/"
�V�f�%6�=H�� �N��۰���yvNV�)X�N��u���g��� ��@4F�B�V.�@ 
5��j�M��x�b�ե���Z�6(Xu/s`i���y�8�8tϜ�A���#Z�b�
ʗ`E�Br��C�S6��u�v�m���8!˕%�$,쒣hS���B.
�,��j��d��ʺTM�ү)]b[��V�ۧm`�@n���02�ŗG3oqM�&eb�K]��Um�P]�)bYi��1�;�uf%f�,SX
Q Vܰ�ӽD��YiPڅ���� 2�#vt��q���i�u�nhR��"J�m�
R�ҺMc��R a�KwX�.���ybU�ZAi7��]���mV�jP����K�b�c'Zvˑ)�����$l'�v�I���T��+�Q
�n���d��A��V��SŸ�!��Z�/>��Zr0(��ޭ�����'�o�	ʹ`�.�X-���+t���Nfds`O]g�&�5����hD7�	�y��{h��tVn](6]k��$�Ă�&~���O�b��5����fX��l��8
D���u�  �4H�p5F�T����(�]��Y�Z�+˚;�]�f"�qV���D�\֣9j4&T¥^��m��B%v��՚����P�]ZӫOh����v�u���fn��
�
�ǹ���[��By[Wu+v�.,,Rl[f��/��.탐7pS��L`(��qX�^�}fůZcL)Bkq!���W{�Y�Ue_�R���ǅ�u����V�).��%��20���Z��'����x(�����I���:�z㼴Ң>A�h��Pa�ed*3
y��ya��P�����3��K�b���j��a(�	��MF\�앑j�h���
�:�b�tj�{r�����l�Ni�n��eB��$V&mE�Їq��.<����u4�3.VВ�4Va8�4`V�ab���K)��7����B�һ�S�Tt���hIv�T��������-�(c�*����@�CIQ�.�'�B���Y��0�횰^��ҙ�Ĩ��*�J�R#wJ̎n�E��b������ʩ�M[pj�T�D�Q���c^u�/�1��;h-\pv2]g�u)�d�Q4�T�G�X�$�Ζ��jH7����T���D��[9��[��f
�c?$�J�[��t�	�����^��V�Z��:,-Y6��q5��v/I܆hz��4�	+h�J��f����jݨS7md�U�Nv�څ8�^�f�clݛ��Q<�4~�B}���y�h[�k5�m^��D�E�)*Rh%7D��j����)�y��"���ܨiӁ�
�����'QU�
6a˅��hj��e�+,
ۙ���He�!�ŦL���6�h�ź�qY����MG&�M��d�����NɴS���f��Y��+ P%���!��#19�g�\״ El6�3U�l��Yn��B��[1�n�h��jw�oS��n[�n�$�Xwk �Oh�j�`V���j����w���`�${�|QӢ���!�,P�EJ-�p9a`�B����FƜ1�չp�濊TI%�e���k�)Yͤ �������	4�X��;U��{���Y|Xi#�雭 ��DtMF7o�@�ld��b(���q��ڌAf�~Uv*��P+ZO*hЫH�=K6�,�f����ٱ��Di^jorՍC]�`���:�Խ�!Y��c�ж#s.����6������f�x��n��V���P,��[��Yg	2�Uj���v�n�q�G^5��+��YeJ�ө���)T�Q<YYE801�ŪJ�h�2˽n�%��K���VAb�â�}��㔇:L��a+�>Z���A\�����;������DBY'I�u��ʂ;q���ãfL�hE�~{���O1�ù�[���֋1�rcͥ�7V�37R�Cd�mjbf�uDAS՜�(�����t�#��,n���0	DV �сݣ7V�I��k˳��Ä%PfYw,$�47Q�Xˀ2ށ��V�*Ε���ܴm�w#�N#R�A*����#�asee�B�v�Ϭ8�z��t��K�*J�sq!2V��Y��֋x�X˺,ĝSv	8�n����{�q<4��64�#d�E�Q������	��E3X��·�v�9G!E�j�86ءkPqQ���^�z5`�|F�W�����h�
J���St�S,˧�kos3F)d�VΉb���tw���´3)�Z���C�����lYnL74��c�����$����P�
�)�j�pV�ɸ���iE�@��F��+&2����g0���'�4�Y	���tpB�e��b��YV��I��l�b�R���3pRL���Q�Am���X��cS�k�H����6�T-b݅,�*�6��c#f�Cӛ,��8ԴS52*�*�����ɻV�t��I�Ⱥ�_:{��)^�Q(.��Y4)D�ѷ�I�}m��j�	T�i����0���N�F�M���Rn��0�aŨ�|�&f���g��U�R�B���A�-F�,V6��8�����/oU�m�f��a��A�GXE��fDޡF�x�U�5��2tbw��,��[oki�X T�)��pnk%,vUF��E�v�Ѡ򥡫��CrQ�P^�Q_n��M����m]]-n��h�&���jV���BL켩��+*A�z7i�,/�&����w@�������Oh3vb2�8~v+7�@�
��ʸ�imo����%��W7i�Ͷ�'C4��h`�iQ*I(�0��s&��¢��[�)�Z��D �z������v�R��Δln����)�-U��'�=�P��9z �R��7%-Qn�q'��r�@$
���R��Z��6�,H�2��%�e�D��V"�iVH�A�E���h٪�(��L3�m����7U��k���p���
u���O�y����B�	�c��q[�@��՘m j�ъ�f�^ijJٴP�@)+Zgnㄚ��ٺ��V����4n�LMv�;�n��m�[� :*M�*.&jZ��e����ѫE;ux0��� ܫ�+È�L����d��{A��lw����ڏ��Q�����	U�A HͧGh-j@��8hV:W{je��į�3m�R��z[���Hn�L_�^���;���/E��(��tR�3:��8�2�kj��,-9n�>�"�ɒڕ2�4�7�v�6H�(�BiǺD�[���xV�P�W@�*����2���E�[�xťP��3X�r�%B!�`tf�]3�J&�R�)#�������AK�ˊ���;�1-r=[X�r�e�gqah,�HţqPD��f����uI�n�@�,H�VecFb)��^��	nm��W�w31��nVc���
[!�R޴�賌�qIt-�ڥ��;F�ȴj����I$�505q��h�T� ��q��Z��Y,M�M����%-�m�Xָ7nfiq `	5�곇����)�D�9�ĦK��^��F�` Q��^)0ȂGl���:������X�*��ȨC��^=��C@��I�`��(��㕅���jZ^���,���*�
6 �l�$7V��9-�?A��P�L��ۃ��<X3jf�w�	,]�Ǘ�[�`�m�,�x�ǓH�yP8$-Â� Rv�1�� Mhj�⵫Uf`�=�H���n�k�2��Mm�����cq�z��g*�캐�A����|1v�J���%u�r%��i���YCBIn��u6˦N,I�u�����BRڍj�K���k�7�����qG�=��ׂ�P��Z�l����i����݃N4.�-�-h���g�J�� ��,��bvJ2���0 ���Z�&�-�L�pZӅ�9tB�Ѻ� �����l,^�M��B��	�)��V�ź�aIeVͻ4�q��������{a�l�+o!G-cM�Iu2,4zTûF�E����n��f=X�,LMc�>r�m�帖�TJM�gI�.�ɠM��m�{����;--Gy�M��_.	��QmR�.��t�U� {��t��+����'q7W�D*�m���a�16*G�7&�sNcZF5���di���)��oe��͉���´S�[�L���M,#I��G!��j�E+�e*���0&�b%������tV�k^�RV�@�n`���wt���U�2�jkV�"�X�՛�jb��eM�n�
���1�S�1�ĵ�ծ�R"�Q�H�6��e&1K�n��r��X���G"�z�nZ	̤�7`)�PD1N�@�
ߣ1֩[׻+p�n:R�C1|��.���֥�>[��1h�ը�VQI�(<u`e�P�7�ȱ�Ic���Uy+�5��1�:�V�O[B�q���qZ��f�.@��m�+q�HKi�Be�X:����5�������e�D��'X���kʹ�lZ٪��NL�#n�K�r��l�N .�e"���cͺ��6�܋)���F�E��+N��<K,}�)�y�:���=T�i���%he��Z"�W�4�7meH�!I@��:wK�(4uf��ml�̙�V8�0�*dǺ�[���]O��h,��m .��X1ݺa]��C51���bj�S�f�X?l5����(�oJ�n����;W��H���rN��%�!�އE�+�p]�-'t+h
i��2��WX7R-a�0n8 ����@<չ�*�e\�9y��;�n�%��CԱZÕerQ��di9�S�gn����#2�VX�����V�G`�)�q���� �@����&)H�b76	J�K��p("�����&��:@W�V����'��r���ІmP'2�^^�V �;�D��P�[ �n��ʕ���U�`2�˶���XѶβR�H��	���+-
��)�c��ɡM`r��,)��R��JݻW3�V�.@3@ˬ&��hQ�um���ԭI�*MÈP��m�A���&��s��,LŌ<����v��v�H -�j̠f����Xop
g6�K2h*���q,[h�KS^���5d��	e� c���`3j^��ԙ�볁ùkke֋4���-�I��&7YR��.��{���`��&������h��f<pؽ:��N�T��f�kdY��YӘ�Ŕ�i��KnYf��Q���i`��Gnӻ�V��jlȘ�ع�)��IZ�Z �SwV��eL���E� �}A�Uf�����{
�0��\�!;���RD��32�4�a�݉�sTF�\�����,h��7[�7*D"f�P�J�Z��"3l����9aI��]n��R��;�Kt�2�t3v��N@p��`{@�����
z��c��wD�sD.����IeGv7cwv��`�����
�,l�i��NEIȠ(���Ķp��3���w�4�U�ձ���Yëe��Ű��j�ݓ.���F�M������P��6�t�9�C&�YqڣN�Z�Ս�[��--��L�4u��ɖl��wv��!y4-�kr�0becWj7Nk��6�^µ �y�9�y�Zq��֍崲�F�&F��A�}�2�X��^=����Zr��'��aw��{{�^B�*O[t�����#O�qV��/�S2D �z�[��s^��+#b�iW�Zy-ܻ�[�-����W[��5V��̃f�&�\A�ߤ�WN� e�J�duΫ�ק��+ܡ5�$� �婃b�B�N�������zƻi+%'����t�AF�hZ)�M��󷲙�a�-<J�g/�/~�:����U�-<-�Ɩ=�N	1��ܥ���nGt��bٖ�Y�В�6�0ul�vf��� rD�j�V�_Za����Yb,��#�Z�	�1Y�5S0���lYU�Z��ɔ�tS��˰槂U��������=x�����zqP��<� ��U�s,%dhۮ�L]�}θ�j�u� ��|ʥ׼�=��1\O=�m�GY,2\ӳŷr��Z�"��O-݃W"��\@f�{��T����Z�\B��͍0�"c '�lf�n��٨�m��B-ց�Ê���C�(T��왶%�p�ܹ���56�z�&���7�=��ң��;u��ZԹ���GAPV�������9�k�-���R@�oX�����4bd)��A�����.�Skl5���6sܦ]"�q�x)؎����5F����e�sb`x��oh<�uV�Ў�[Pc�j��j�iե>��"�NΝ؟?-/ׁe�����j��wS1I�I��o�R��vv{�⃪����5Z�K� hW)i�ZZ���1�9M֏7Y�~��A�lj5��%�J���L��2>��	e����}ҭFXJ/fj���W�2�Kgd�1U��;��m��ƶ��E�.���uqv�;��mۼ���<!�6���@�ֱn�\f�#m�Ptf�xZ�	s3W��������R����Vǵ�k\��"R/6�p�a�!�㨴*�k���.�{WvS�S��N�wZ�G�v�3�Z	��9.��;u����%A �$
����[����î���oD�V�3�\�Ymi�z��i+$Ztu�(lጴ��HNK�:��HpE�W��\s�����SK}U-.'s��'��esH|��U����iv���#�h�u	�ۨz�^e� S�8@`���gk1�]����!���7S��ӄC�����,������k�}�A����!�s*S}�=8Wf�Zk�j����H�b�V��H*�`qr�-M�P�[.S��n�g,K�l�����-����H�f��{���]�0�m�yY�T�2�2��e-k��C�A�X�򺽻.���ذ�w��/�B�|ۧ�e�����G	]Z�5����->�Z"ZZ��ϺK�,����|��i��뷼 H��]f�׍�X�5A���2�L�AJH�S�����$J9J.��;��_vơ7��k�)W׍��j�v�`���*V�d-�ZQn�GR|Ν|�T]�s�Z�D���+(܅��ݗ����Ҭ�}�Gi�AG]��|�k�J��=Eˏ��s`��+��T۽�`t�b�z�q�հ�V�8h��xY�e���)N�)+�G�]]h�.>�ɹB�Z��S�Y�)���2
���2mZ2��.��y�U( ��	�_=���;�n1%��b��2�wJ���qů''��=yuyee�ep�y�'�o�	���ZrҊ�Kw�>vG^�`�룓Z�TaV�<��%z�[��h$.=����`}��5��v�w �bo,�l�J�@̌e_mrʣ9���尻�{9�i��ٕ��n �s�@����ي�"!q����ڝ��ܳc�]��l'��U����!L^��Oi*\rZ0݉���E�h��W;��he�i���|��k�F�T����fj�s�����۠��l߂Lo�Y����_i�0E�:�ÉoT�Eپ��K8�=nX|�<J7�N[m�M��\o:���_f�N�Žky�n�V,�@�-V���[nm�ꕸuV$dR���,V��䎋�^��c������FN���ʔh�7t���N��/N�k���d˚V;�'`����u�}�!�ޠ�R��H��m]r��ۮ_Y��o2c���)%Ϻ���`�r���*��r��\r�e�PTeC�'Yr���x��'n�.5vOcY1��Vͯ�AV��/pi�]D]v�1��E^�פ��er���%_>]�Y�EGz�,�Z�M|���N�� �WktK�M�{ۙ`ǛK
:�
�taXs�+b�z�ޙp��t�t4Yr5�_��r�mEv}3������NM�;R���U+ڢ6���ӊ��JPn�߃���l��&2��q�T/]\wy�����A�'`�<lt�T��[ԇ݋F�ڜ[��rlb�i�H��EK�hO �s���sf��y��];e٩���+�]�ܦ��6����+m���)����q����
���ָ��m�a�*>SU�-�b6.�tę�V�l%@���T�*zcɳ�c2J��)���� 3W�ى�J���C;�T��Sfr�/;p6���%'��F7kk�W�(K"}m�h�w�������
�h�dˬy���]y}soM`n�z�f���9�E&�NK�m>��@�嗤i*�]RC��]
�8�8�4����i:6aݛi4���N��6�ܚ��뒽m��n����f��R�S*�-��:���Q�Ӻ�CXP�S9$�ɓ1֙iA�o��z1���>�6������/�/P�u4��^n0kq� 
���2a��֪�t���m�{���p�0�B*�;�O�#�
�h�GtZ�c������f���!qm�ǵψ��4�]�>^��>{��V�{1��wVV"�J��O*#69}����$^Mz|R|�;6v�n۴���ů�R�X�t�������dA�����\qy�7����n��Q�Ug2����f�k:U�>�B1[\�
���`�"1N�*�g2�@*�����ޅ�*<v�pP�k6��Ϛ0�f���qi��.�w������6�ġ���Ӆ4h��n��QON��z�I�X`ۛ�Q��[+!V��Y6��- �D�e
�75�@�I��!���*�[R�"��iN]���;�R�b�u���]�NѼ�w��r��-ڢa�f�M���4�XN�&�x��ZKF�FMCB����V�ۏ;r��t�[M5�X��`���Be�A�/����)�<s�y���,���$m_�P�7\��!�jj�8��n�p_`F�,A�2�a#G�r�;h�wنդ��K]��:1�A.�����-(l���Y�j��t�NZ7%�uҭ^il��ul`�&ZTh2��
��r�ɛ]`KT�������KHB.�Q�.��N�>�78�c���6%k����r�����l�t�n2�<�Z�keF`5(�ܽ�:lRD=ov�ݞW�J��
�X{!�i���:
��`T���K���S[��=ӊ�Y\��)�-ZǛ�v�CTxz�K�M�%c6��)��I�S�S��`Jt�:��E�۩�*c^\�]���*���}�u0��)�d���\�|�*�T���E���s�ȩ��Bv{��W٬>��!��IF(��v�=cx�xXo�V;��@k,5�bb���[Ztv�n�c9��-&�5�9�jPf|0�W�11��/!qT�[����݂��ݴY�Z�������ą�kB|��=�a�O}++w�/C��f,L����vk���EeA�,[�4s3\[6�d�oa7)��w���ֆr��T.ڼ�xB����-�غY�z���)b� �c�u+�q�w���N�I��eN�ᮭ����<�\hI���0�Oqj֩�rď��\o�9�w"���T�q ��=���E��2���j$ڗ��ر!z�ۮ�ε��H����kN���WJ�S"�$��|��W����蚘
Z1N���"�5�K]�ds�d�A���T�o\..��:3��ns�]*�ue���iεu���:�8���[��p@0֣����,��H+燛�LL��AU�pzപh<C�S_K0s{R蘷��
���kB��'�P�)s�����-'0:�l]�y���/�r�ù���ʵ�xm�����`q�\�Փ@p�V-���������W�aoN)�'�OJ�{"��{bp�K쥼X��W�`L��ouAC��2�i�~1�\��G5ֻ�&��SPTsYì��gT}7vQ#�:�k��%b��a��җsw �2S�n>V�m'��"�!�مg0Pg����v��&�ᇵՁ�̕!J�w��v+��A,5��V�`�2�j�y�� ;�%�7;uj#�v�su���j�!5RV��RTG�մ�h�2rzwz�̝����o��b��e����Yl��N��2�P�Je�5pdʳ{���1Ģ�������N�H�k�i�u�����g�k!ݵ±.��#ށ��={���-.��]9�e��3�v�I�͛�z�jpȭ+�;�c2��-JؽHd����"]s��K�o{\D�K9W�F�p��v�E�T�����ݽL[+�`���oq��U���i�;�}�Ѿ��3��sA<�+s�V����g5���v�rQ�ȼ�	��x��JY�¾_^�B��×���@�O�!��X4���:E�.�Xu��"n��1���i^�}�E�w����ݷ���fC�Ҋ�=9.�nM�u̺4��Ә�d��u�t��lv�x7�$l��\�=�\��&��	�ј��h��w��J�������Ɯ;�M����i�Wz4WS�-9�|b(V�M�y|o$��f��[�Q��Pv�9���f��F,KE����c�*0WR]��6�݊�[�Yo`n,!3n���v1��6m[�E���`�e#`�Of���� �����99��Z�glf��<�P�����WSxU�.w��Aur�&4]�u����~�Kf�n��A�gv2���,�j�)w�m�G �J+�Zʫ��(g ���q�&&���]&:�'r���e��e�Y��� ��qī��Cfc�M�W�Ӷ_U���p��&XCt����ڝ�9e�_[�N��	�
�m�C�b%B��_`�6�~���i���
��*�4A8er��X�r�kZ����M�]{��H������yI̽c)�
j�lj�4+c��Pn���e�Wj��]�_D"�r8OZ�t���KN��r]��j/�]��M
�[����Uu�n�X6����n�pJw�4�X)��io�J�R��df�k���=��3;�- L��C8e�����M
\G1�p�w�U��}H��fm*W5Q���+e��t��(�J{ۘ
5�*����[�"z����������FX�Qg�<T�X�hn�˥�e�*��5ca^�j�<�R�#b�,R����R{/�]�k���
GO-�2�M��3#5erJ�m����)��t�E�u
���,����G�*����\ehW^�K�e���v����Dկ����*��p��_��m)N��xX�6�Q��{��h�v�m�sg[OY���t��in�$�І������v`���e���]�q=����S� d��&�aU�5*>���`c�&�gI��-��Y�A�"�Ͷ��x��k����O�;�u��H,Z����s4ep|h�c3��ؘ�Y�5�x^V�7��� �ⶤ�s���͍=��2����J���ᴅ<�h-��۝ђ6�M�I�u�.��� V�Sk�`X��ʽ[[D^p,l	��VP�]h��\n�Vܶ�_5al43���zxK�S�Z\@�< ,KX�؎�ː�"6=��U�.�崱\�%�pcҶcnW+��ɤ����~�o*���&��I;Ne��bA���73*�՘�)!Dp�.�Z\�T�fH[!���<���܃��sdYW@:|a6�$T!���ц��,1(_aVQ�4��J�\�d��q��ͩ�z��D��gj�xv��Pp5�33�B�Qe,����e�P��`�N�,���hnpPF��E47[L�N9_<�|`�(~-.6�v��5X�S����1+ܕ�������g^��z'��aY�]��Qt\!���}կT.�!n� ���R�O�=Qهpڭn��)�eM�8�-X�J��&�
zqQ&|�8.Nuњ�o,;{��\^Q�N`ֺ��2�\xe��t��O22��i�6%��oL?�v�y��VwĎj�Q�k��
��X�V@��K1�ii�l�N��С׵���:���B��k��ެC��&�	iE�v+��GG8��,�X{%e���{��nF	��#7�;�,M<i�X����*:��]P�ج6�����H3�-#��ޥ���v�wf(@���1��4�:%�����բgv��\]��� �U>0�܌���A;ꑷ��X�:
�.�Q�s�Y�����6�K����
aM���u=�E\��&�
Sb_#�H�iհ�v[�޸�wr�=d��W�+@��nbj����*S�!��Y]F�Ʋ���,Ј��Օq���r�jN���I��|l�W�9�7ط�m�쳎�����iz��"1r����� �:X�h�n��D�ep���Js��ܫJ��\J��w�Y����ɑ�Y?qR��/�el �{nG~
�P�H:����r��yt�Y&���Ѥ9�/W_N�ڛPݞaZn,�7D<�-�!u��9�8�FUu+�A�c�M9cqiP�=�f�z]�L�/@�(S��X�U�dȖrgA��PwRa]���[�r���d��ޛEՍ�5�M�9�B�bf��6���OA�6M����l3jд)o<�j_E�h���;��0ܐPR���B���=�{�9}��i�(ˌO�s���uS�[�[c ��F����ˡ�8�}�����N����۬a�E��eu��Űt�%�h�eh�-��6�������7��e�q�j�}��^Q�mֲ���n�+�a�+�r]�5�/�\�@9�d�)�-�⢐��)�"#��+�gsY�g^\�u󠑵%�Ok�%�Xk�_Z� ���}�N���R�Y-k�W:e@�-�����b�����v��ŌX�a�Gs}I�r�@��ݧF�`�\r�Ckk�1H������&�}������u�x���a��E<�`yz�b5`�5K��� �LnV�p�Y%"-�f���w��BskLj�+8���j�n����2�.n��[X��zvka�	�4wV�&��t�8�Sx{�6���ہF��N�(opZ�܋��d�Ҳ��gsV�lZ^�c'EO���Z\�ZB�m�s����u"��J�7΁zj�Q3�P�E͎�*Κ����DnF�;Y]iͻ�s�
��"�g��؎k�g�<�L�yb6��'�b�7%d]��;����v�I�v��ﹶ�cj��z���W��c�����	�����7s��uwA�a����k�=v���q�d��ŷb����tn�s�<�&�Qi�s�nc�v��$����}�U}�}����1���l���ϟ����O������ח����`�՘U�@�H�Eê�|y���NgqGd���[\�
��ar�*L
�
ɵV��5;
��sW;6t��^�)�B�t2���s�����zy�q�I����@,�=�l�E�*�]�Z֑5�Wv�,���]2�3:�]���.��kB#J��bQ:�)��1G*��ݷ���t��[�W)!1����Wa��y�C��vt�*�?*=����4={}�"i`�^͋���O��+���CQ��Z]J=O3(�m���v�p���Jת�n������r	�4���N��`��J�)�xuXA� 3����iJ�G���Spb�%\';YX �Qw�;h��Y؇F�`S/��']��z+ev�����`Wo&����v�F
Ԡ:�M �Z��k�rJ�g)I��K��u�e]���Zݥo-ӱ�x'����Mn�':Gx�Ү��![N�wmtS�Ѭ���l��W � ;MԅVj�g���nk���Ru�m���ͻ[ow\�C�G*N9�|�� Z���L�x]�]4+��oV^�è��I�Ι�	��f�keq�/+T��.P�wM��S7ۉ`�Sv�m���۾�ُ�bsE8*3����H����)���M�ͩb�L9�)��\1K#�=��k��C���S�v���yP�+�(��ɫB{�V)�n'�CV�jٗtVӧ&!v�\X�yfg�һ���n"�ݠ���Y
��s�(�/L1s�Kr�1 ������<K]&n�Q�X`�s,ݺK���ݗQ.��y% �_��v�%�RtD��ޔ%�}���YЭ�԰���]�+34��j_ܶ�8R[}�˪PW�',�5�mY�69A�����$�p��֙Z`tr��t���|]s�y!M�˓�րlY[�b{R�[�Ӷ�yj��&�A�eʝ�)��ۮ��'���[4�!�S�qɺ�Y�ہL	R��	��A�ѻs*� �;N�v�y�ţ��L�w�����x`;��O5��E��w����)��}Hw �(��`��XK��#e(�w���[f.M�
�pm�]޻횷RN)ŉ!�������{عs	�AIu��/������bĸ6c6(+-26��^n#�p:[N}d8Y��c��JN�}M�,>����=�U���������'f"U��z�B��YzHvS�R�I�ɡ�-t3;���k+�|Y�fc�!Y��i��^J�Bи�M-Z�!���Q�9g�fn���ȋ`Rɔ��j[��G�w,�$&���;�T�*�t���
��N��Kۗ��Y0�� H�M���(���Z�Ŝ��Mft�)��\�Rt��٫{�2�01���ZE�J���k�K�V�ϳf9
�c��$�u�6c��V"Y����R�i{[����&u��j�+yvS�e�H����Y�M�@���w}����]z8L����b�$T�|�[Kw�+��>�V�e�렓p����B��ё�}�����K9��ַs#� N�(�X�.���"4�D��z��,>������;c���i�3E�ه �5y:�y����v����n)��"�֢�3�sz]�5����1�"���;8oWT�_4G�n��Т���n��|��kDQYj��	���E�c�cP�n]�Pu7m��YomN4����9>�Es���F��i��#0n�vۢU]�%���I�����.�N�je�CPV�n�Y�����2���ן_N�7Ox��JRV.뷖u��Y\�U�7���0��E2�6�^��,��U�C׋!(tԹ��e�Fq�ʵ�ȵHL�vQ�3(��M��ͭ��ǭ��v����gfp͹opp�e�� ML�Uu��Kq�+5�4�T�e�+j�|5�<=�a䛾8&3Q��1*T���,�j�f�߷6���Wcn�=E�o�Қ�v����:�kX��4��+�kx�y���Τ���WWEu�/Ptl��j�#; � �fvRxPb��	w��l6'<���"_��Np�3K8h�t�<��u��R�7e|���{`U8�T��]�͙B_+�J����N�9��SY�N{���\�Π?���X�g%D��p��+����dn(H�Π�k�ަ�����ow�,ŝ�?�P]��j��c�b�VM���n�e�1�C��46�ح��
���qˮ]�N�2+�C�VR�lc��}n�Vb웴	Aڕb�T�i�Q�Ԝh�RR
���.
�^�� �\Y�q殼���Ҿ�Si�8�����z��x���e<4��I�n=ز7�����Y<��Y�#	X&��-�J*��U�M���u���냆�VST[�$U�霧c.�i��*�>T�����&ZYf���،��0�9�'(�p��,��%jr��l��=�Q���sQd>69�*�|ݠ�v�m,��7����ʐf�is@T�=��r篃@賆�T��Gv���5�z�sv��ރl�	\��2��dӧ;vC'����-uc��D`{���ů���gyX��Ob��#���tkkOE/�-�ֺۛ����јf�&�� �4���vCI['���P&Zݻ�7 ��hS6q��y��u�f5s{,[" V�c�B�XM&r�����"�Ey�s��ǮWf���K|j���eƵ��B�o5}N|�P�^�w�5�,n'5������@���C���q� �v�n��\�����+E�S�Vo�$8�H����;���m�4wE;��q� F�脢�Ũ��oz�i�����g��B���PP�6V3&�$�l�Ϣ���:�y}Ƀ����ņ6�[*\Dc������^d,w2f�X���uչ�S@�Y�&`O��T�z����ѩǤ��
t%�A�;nn9�E�m�qܮz9��<�՗B�qZ��@�E��n�-�+�|m���	͸(��:��(�k�վ��,plX�Ἦ ����j���z���1\x6��4���O�ѣ���G.D/ J+;�A\����Н�G�;ヲ�&����G	�9n-�b�n��5��R=л����:Ӥ;�!��+�����5������$+&�B�W���7k������w\�%-���@���]�YPJ�m�v��k�܏o�wS�q���#���)Tኺ�=SS:mJ���4���7b�t�Z��eX.iWBV�Y�`�i�toG����.��%RPWot>���c�| ���� �\�{��DUV�颜�I͢���"&N�H8CQ�9N�jޣ <� �0h]��Ρ���b_a�%��Z���\���ݾ�(��8bڄ��*uL�*[�XΤ�+Эu8,]��i�ېfJ�o����U��Te��:
an<�L �����M[�8����4^C�V��䀥\����wV�b�v�k��+N��c�(����u�*�h�r�1��!���J8�9 �Hf[�3��A��/�㭑�p�J�Ii�)j��2Df�R�n�'���hSO�ӷ�� H���Am�Pim��ï����O�у6žsr�l	�V��Vn�4%^N��C��q�����iJF��I����k���| �4�j���gQ�m��ޗW���5m9���=��n��!��崶��| �B�;y��U�\��J�ʙ��;Q��/J:��w$hM'����CwU��1��0���EJ��w7�@�o�]2<�	\����H�j6wjz�`�jP&�mc�e�gh�dQ:���m�Ή[\5��B�����+��[%��`�o+v������]ilk��uK�X���]v�v&�t��9��:�f> ��dZ�n�V`��aq�w���sU�jJ��EhA;�*�h2\�ɬ�4��1n�jrԩ����_V��QeK�v�%�!x.n�Ea+JZ��@�ʃ�Ix⹄�03j9t�oY銥Y��m�y�r�W@�%����A �녇�E��V��0[fwe���{�4؎̽u�n%{zkjp���F����KD�o��X����X�t��Ά���:�)k��r��I��ڢK�5W-��R��x�%v(�l��K��]���d��q���_LT�eq�U�91�$��ٺ[Ѐ\U�{U	G(���Ǒ��LΡ��.Ҁ��՗�>W��2���S!�����ܞ��F����F��q.�BW-[y�O)]�-Y�U�V��'�5K������8��v֨�f,���CP�/N����鸊HV�O]F������n�ٝr�WqU��S��{4�wr1���8�[�d�q�J,b�O6��-���4��Vb:�4_P���=��*��B�uuã�b<���ٕ*�mx!�V�r}�-(\�����C������8(�@��-�n����30jܽ�8����ڶ�Qh��o��5л��j���ᴦS�y���E�]��Ea3-�[��g1��}@x���Z�W�,cZ�;����/ �WES�D泼Xe�Vx�췻�����0��+�GYc��K�n�6�&_.�튏X"�miD#;�����i��i�|��5�W63WD�5��G��m���.۳4gm�nT��w�v���}�zl����v���[�Z{o������cY�:��M�d㋅�cj;�7^�u��TTWX�!:��������
U�v*���C��ۼ��Ƴ|,�3�SчrSPsWƂW��]0�	o--Nˮ�x�֪�ϛ��JVNQ��h���4�XX�!��r6�۳��gGA�f��Д�W��M�:;ۼJX�(q�B���\
�Ѻ[����ꝩS؟PTv�YK(WX�C~:0Q�:��@�xF��O��a�J�
��wֳ��np�&4���
q�e�M�v�j�T���-t�U*2��ZKv�������aȀ{Ϻ�ݴy���n-6v}���ޟ4��5�������w�<@�Y�;hnG���qIR�u�ә�ҿ��)��[:�N��[W�P�M�N�p�' �{o+�`/w��(��i��a��³u�T�@'3<t�A],�m��wѬ��YGWUȫQ�p?��̐���\���I��i��r��va�+��[���n�2���Ѧ/j:l���8_�Ԉ��n�2Ւ�T�\j+\>�kOv4�9�9�|]�/��)b��1R��E�>kuM��J��(0����v��̼ܖ��a#v�/z�t����4c�,\��	[ܳ�km����`� �p��fI��]��IQPV���ƺ�ƭ�6|ʨ��RD#�_
��.�*��c������ڜLk���s�e���F�[Kq�igH��P\�d�� �R�`�*�v�|�9��65�'R��wE$��HK\��]����T�fF�hj��O�*��܈#p0��m��,Vv�����%��[�.�`SGRYd+p���W��m��Z/���i��u�t�vD�Փc 3S�d��H�juB��[�xz��s	��Ղk7��R8+�WJ:�;`	��vt��sV��m��uv;��u��(�� s��1�d52�ݱx�nF���2��]��=kR�˾�]����1����.��(�+"�b�Ԟ���Ic��8A�����A���Vn��0Q�(ZG6L��[}��G��f٘��t�b3�D:o����L_N��odQrt%n�����|�1��dqU��!����f�oo#���v�Ab5`m��3Qɹ��_b�ޡ�F�u�^�m|����R�M�}ί��2n��{5V�r�� �+��Hق����e
$���@���>VU�7fJ�9vr��Q��n�B>�$룽f��p�%[��v5��T�M=�V�u���hiY��6ј#a`Kh�o�K۩�#���u_c��+R�-f �����j���ʉBw��%��b���z��s�Uǧ����AJ�V_2����������[��f��W�����آ���:nM�`(0
1��fh��l@VQ޺R�A�i����Mo>�b�魛�T��n�0w�g\�d��"V轳��@@�A�V
$�O��:�^ˡJk�:F�r�,Ac1پ�*���
�r�L�Z�Kݡ�M�wvg-�{I)�����i}�6/�a1r�b��Mv1N�M+|6N=ԩNvl��h]У��tH;}Z�c�i]�Qξ����mpL [I�p��y���h��rܾġ�7�S��5�U��h3�A9{���e2,9H:�x5W��b �e�;�!�̱K܉Etᢺ�iV>�Y-��ڗJ��.|�X�����YS�^9�D�
��I�̷��{�O5kƒ�e��;vdR{�8�\2�W�mD�ӛ��;��co�հ�WxU�D��w]������G���]_k���u�,���[݀4g&b4ng-�7��D��<6�-�T]e.ܠ�a��4>Nq�؆؋�؁"�+#8-��>�|0����{.l� )��Yh��5v:z�u�8J4�鮒풏e�k�H�@tRWi�UxC�Z.I1V�=1�D��Ck3�X��m�,nS[�S����7l�(�ǧv��S{ѺR^��2�l�{�Bʐ�f(���;d��ULЀ�u�n�7S���Z���퇫6�Sl�j��ͨҖy ������N�4R�|VEEXG��G2������ne ��l���X�+k�6G
��V'�vv)o+�$�ۆ��M]�<�Z��Ues�P��C/nEZ�(�u �ab>�a6v���,p�3�;u���߆�u,q��B�ˎ|k�oh��M)�EeF��1Qʽ������G���?��a�F�,�q��ף$�\#��9KU;�6ի��2UL��iK�ʈ��ے�A�&�Y�W ������m����!��;ڛ�}fuL�:����g	��
�6V־���m]�v���K"�tw;��4;Tw�Rձ�4dޛٜݖh�!^��!��j�UM�V��ve%t��6u��2˾��'�+��'v�w�Cc"�f�c6��1�	:ͪVqV�;��&�5"o��޳w��{yb��y
�lp�N��t�K��j���G3b�u��K�fͼ�V"�FЋ6��K�奓�ef�F�JGV���N�y�\�b������/X���]�d=ˍ�w��@��ZS���9���en,�è�]EcL5t�[�bQR�ŷ���y�9k��k �E�sE,+��]���e'��ԉ��5��9r].������e�Szch��(�[Y[x�	m����������y#W���Q"-V��OĹ4���֔t�ͱE�<��VNm,�ӕ�a΢(��g����/&y2 �|E:4]�}�P���*ι!R��S��)+��U�&��қ"��DP:S ��91VǸ�Nzj@�S/w�=��WӉv�=�㊮4�kt�(�u����Vv��޵|B�$�s���5�<+(�8�x���|�gۧ
�rU�+�)�W8�Ӹ�.�%���-�������w���33��Tt���Rrʫ��֓ݮ����2L�"=�ȩ��Dʋ�dR�,(�.($Y%��E�TuZ�Z�M�+1"��U��Zf�#R
�(�B2H�"��+�t��.\����QQVs)
��PQUp��y&�E^g*Y\�0J��J
$Vr"��CA*���**rؑΊQU\"�Q$�8E\.&s�Rfl�S9Dvr�4� ���E9��s�������uiDA\�DZ�
�9T�Er#�^(�ő^�QUg��u:UUd�4�L�a%fD�"����Q�OA�n��*I�+���rԈ�#��qTQʨ�:'��1#�s���PUl���PT\�ΕE!
�L��*�����s��~yG�~�=�0���i�͒�5�	r�(�I���;v��ɦ;#7],���;��Ѣ���wL�CY��~�n���y��W�}�5�7����Ì�N��
rv]N��g�3��"�6���x!����zA@a�F2�Ë&U��m��Ј��]+D��SŚmf6*m���7Rm��$�]���#o��2.ei�#���:�Oʢn�˩ZN���75]֓�Z��6��+W�f�߹8���ٵ����8���Ez�U�w�
�����Y~2�#�=�J�p���ˈ[LԮ.z��]c=��XK9�#*��B �}.�ꀲ*��ϧ)2*���/�=�e�0B>�W���y��2������OXg@��َ\��N��!}�8{G ��g� h�pX�2��L�>�@]��K�t�(��WQh������tM"f�+ީ1��V����#<A���tWP�_*AG9ve]�ԅ��>`�x3�����i�C����;����`�LL,��G��"��F¼�V�OS����R��"Yzcp������\���@�}D�E�u#|��ܙY�8��+P3C��u.�[��7"��(#��E]����s��{6],�� {^�)���4������ݐ�q�;V�&!����.��9����H0T�A�s��W��+W`��T�U��D�p��Y��9���[O9C�{��{n�q]|E�������]^uf��ΝW#����P��K���h�T����k��U�J{7*bj�o�x����o����,�Z TO'=��P����p�t��l�7>n���z�'���?X��$��[Էy8��ۨ��$uA�|}���kG����tF
�I�C>r��`d�M����Ř�6r�L�Q�e;�G�(hп��Ҷ��V�_�V�j2�T2d)�Y�;�Dm�Wm�7��`�'�#�v��������ǧ����T�v��f1K_K��7�g�"��u���V�9�����L�7�6�x�P��� ��G�aB2���a�W��÷���D�X�Pzkz���'v�g���ME�p�{����U�������EGҺP��'�\��ڃ}Tk��o�	�������a���jt8��9�\c�-<ۭ6�"n��z�[�kkI;��� �Ra�,ܤ _^��/��%O��s���δ�NXq��[=�U�q�b�U�Iݺ*�G��ժ���,*���,��<��	a
2=~����Ԅ�ʉ"@z(�
dk���Ok'c��ctw��j�T��/f�#� u���/shd#��~�[Ӯ���l�;w�qu���+q��R�O���n��z����RK���n�xD�S�
o��XVl��I,��s��{oHrQ�n�=)�����]鐊D %�����>'����@i�z��Ni�����Qx6M wuj*���r/�n�P�cU�xg��I��3�n�k��K.=3=�U/�*�^Jc�X�Ls������n�낆q�xAF��H;FPY�ܗ�&����%� tF�3t��T�s�jb����c�����:ڨ{�Z��,B��w0
�k�l*����I�g@�q�+�;3�wb.T���k)��N��� Ƿ7�Zm�MM��h�Ɵ�����Z��0�IJ�y�\�}¾���o�N���)�����]���
^�X8��yQ�c�u�NT>��A��� B������)�S�Y����(z�[��)���;X�uX):���4z+&�?�=�dW��I��Vn�lvJʛ��D�W���7�s!�M�_|�h�c$[ɂ'�aEUp��|���|�}�Tg��v�H3Wѻ+M�*���2cRN̛Nb5�#Q�_k��
�'��dh�y7�.��q�y���ڋѾ���R�h$`�n�dR�ψZ�u,u����DaƱ����L��N֍�6����:�H�v�#lۉب��p��6A��3&�7�in�}��#v�b��56��4m
�֪�޻� �&ke�3����,�m6�l�w����B�n�b�ᫌ�Ckz��.9;�!L�X*~?u�	�~� ޶�N�}�*1u�lyʾ4�Ք����%ז��j�J�ULE�'A��'L��UPU�݄�� HS�Ҙ�_s��id�|��n�����6�`�髼s\~��L-iޗ��\m)46�q��!k���k�s�9md�~��_Y;g	B��{��m�������z��Uz'�%�s d@�q��oo��9ǃ�4]v#�.�ᎂ_H<��q�냞�^��1y{����F���e��LFGs��]�e�T������b�\�7,GwO75�*@�{;��q��45�,ษ�"��g�#�}�U�B��l�v\�O��1]�0��\~v�or��j�a��@W��*?iHo�mxW]>lW\j�ϡ�C-��D�N���j=��%}�\�����|�P1��h�F�xs4���<1x��7$���lJXs���D-6��F�w;�U
@�B�
b$0���� ��U�f*��e��b�e��yR^��n��e*W]��=��;���C�(�dՄ˩i՚�F�N�(��T!�&lq��#��s�
��׫kU=�H�H�0m�%��Ѻʕ �t���Zy� |��2��H��FY�N]YZ�`��!�)��U���bxmBk���x����B��n���HR��3���w?��I��A�7q�>�z`W^����'��*vٌ�se��f0ECn�v���4-L�.��*�EX�yy���6���@z��dп�fˈ,+�����[g�Z��l����0�����"�-����gq[�}"K�)f�:<�g�������b��?RJ�/!�`s�s|��w)���򗈊@z�S�U�Dv�	�z�gҺ�NEc&�/.��t�&���D��U�{]!M�~dj �ܾa]��	��ş�GK'�����ȧ[��(�/��*���
���=K�a����J 96$!۪�FL�G7,ta�l�1��V�SH��\"ͩ�̞c�Ԣh���gZ�����/���s]Sδֱ��px
f�z屢Vv�6�{-^�k��g�8�T~��r���E�Yg��\@Nm��n�r��|�^��:g���T
x������5w��K?]r����2�la�b�|���Ree7���1U��v�FзV��
W� ���J����dn+/-$��Տs���É[��1��jp�v�Z��e�5y5ݻ� Tֶ ����AV�r"S�y9C� ��Z���A�A�:���G�o �A�6��{�g2���{:�E�#���gB�����Jg����Wu�4,����&	�0x�R�U���������'�=�5����x���^3�cݟ(��Ҁe<A���5�X��8�����N9�SϹ��u�d�b.��u	�R�1�+n�d�q�I֗ �z:릗�nL�� ;�Φ�G����K�������v��K/K!��p��8�Ȁp_QD�r��:��w���.7�oh�=�?]uSeӟ��r�k���Rt��3�T:�B�.J=�j쭧O8F��e��5��;�]�S������,n7]Ľu�m��:�Z�|��<}�\�^����+H�#���0y�Q��p�K��pF��&�r���}T-Z��)�9�숰�Ԗ�=����к:�K���g�ڸ޿��H�e��]wH_g*z���P5K�]��lK h�c ���6���|G�ٱ[�Jgh�O�eJ�:.i��2�!�+*�-r���MTQ�2d�n�������0�Hd,>��7�9-�1H��sΚBG*퓶�^�+�E(���or��mj��,���/䝖����~�c�>�� N�ы�[�/��&�NВ�B�qS���Π���l���}���0��&������'��atx%i��Y�����W�*,\>�,WVpv�޼�y��1���M}n\����r0��� tN�Z�UV���l�Z��qa_�8%&2/'�&��%O�3S��.#���w��^�ㅊ6^���ŖR��/�1`���A�߁���������v� o׮��
\�7	S�10��[]r��'���Nˉ됪���~4��6�vh��W0h{��V
���=>�]dT�FmRB�
hk���I��Rk#@q�_l�su�/����K�!-��`��5���DUz�ƅ�9i����m���� 
��i�N��9|_ݿ��B���<2�I1$�yVJ�a�4��[k}���W�~�H���B1Q�0¸���6�+��eey}�p��p'pX���g͌���~;-��(�[k�,��L�S=x[s�����*����&�Ten�O �ثㄝeh	���ڨ.��r��e4c>}'s��Ю�_�=N��x^
�0z��u2�b<]|>�������0�T��_�<�K���P��D���¼�J��y��m�A�΢�k���G�~�ӫ�Jĩ�8�sgh�,�!�����h
��1���i/'=��A�xN��q��K{)��;�,�Rfc��&��8�eH�V�5Z���qֆ-��0�N���La\��4����2�:�����a��4�%�3a�&�L�5@ď�0R��Z^!qx�N�֍�8�jUXk��ԙd��ʇ;X��z�^o'U���=�@�&p$��Y2���ö[G�����&/R�ro��8Cg/!�+�_��!B�L��:�V�p>���Z���N0m�q.c�,1�^��R�|jL$�<��k�F�#\� =٩��'�6�ۓ����8�Sk���\��٧JGX/���/p̍�çz��9'���0�R��\)������L^�xL��Vuc@��^&?�*��t�זaTG]{W�W^ګegZ��}u��8K��N��l�����f�⠣~�~�ܺڤ<5a_�Ct�"ϸ/��t�h�F���>�ݮ���������1^��9q��p��1�g�٘>�
�1a����u�z}:x����CTV>�Y�J��@�,�<�W��s��/+ڜG^���J���\��!v��Nɰ�����e �4�Gs��;��Ơ��y���Z$���f��~{������tb�ee]@t��2�V�}A����2+*(GU��]r�����ԝ�)�WcJM�U���M�'F�ó.�4�8��{
Uڋ���;Yj��=y&�禹�D�W����]H��rN�a�\`w ��#32IK���B��EX�@�0[K�5�q�3A�iW��:B/�n[=��[�#�����Gi�����P�wH��@h���Y��P�n����_U{����Y+&;4�����p;dY����ߨ����� �g���b�� �%��1U��F�՘�]0�i�y=�M�5V����p��Zn�H��;����ϐbt� �����0��K�Ϣ�R��~���"����y��^2䡎ӟ7$GW�����Z5p�A1�F��w���G\�`�7$�sm�3�����B��oWϕ;l�@9���3"��Q;n�١jd�)I����;6�	^f��"5��㚦�������+��P�[c��� [%tC5�3?4; ӽ�R���!x�g�`����.M���U'C�_Q\bs�ѩ\�.�?SJ�-��x�ֺVK��{�`r3�bT�V���k���g�����NS5ᘙ���<ׯk�]�V��\��V9:��健�#46ˌ?	�d��у��߳ؐ7��7���ԉ*�^wS)
AQ�9'����ݽo<���K�]v�>�!K�̝tHM�W5���H^�V�m��PS}��^-C����f��0��٫���nH�t[7E�3-�]�	��Ԫ��h`PAE�.��N2��{ko���{X7�54f]��X;��Ρ���j>����oA�~���ϵ:��!��n�W92� ��Y�1}��yk*i�h���^��{��{�8��ܞ
�\���*w�o��S+]n�U�a����Y1�y���y&wf�����Kk���������k!��TGAN���n�r�Z�-��wX�c���\-�L�q� ����QW5�Q��	�W���i��>uI���z�e�U������/�����Mu�9g	J��b`���<e`���Aw�~�?P2�9.i�����a�+�2]M>�~��bߣ�m*Ҁa��?i�2��[�AS�@�N�;�cf.�89�T���4C/�w	�-K�+o��	��A'Z\���	V��e��Y�8��������Ѹ�	�ĭ��jK/�@�m|���y�8
5������'2} �ՠ�sޟ�+��.��=X��v��jN�g�)�B�o��<9�f&��ɮ(� n� t�$��Y�P��xh�t��3�X܈n��}V�0Y��kV��߂�r�[}�r�Nsp.o�)�I�NU��Ӽ�`j��h�Ф����ܭ��Mݑ׼��I%b��KKk0V�>ղ��[C2�:ɢ�$��-��譖Q�#:�GF���Ӝ`9>S��&�R�	Ev�g��D���է�FP4�q��b�]L^P�	�D���� !i��*���;O�}H�[�(.�hU��������i9��|�V��.�n�����% ٳn��]���H���o$������m��hw���Uo8������qPAF��lPA�����ꤢ��Fq��MQbU�����W�iP�6�v��N<��f���vT���X�hZ��ى�1�������z��ke9Ѯ�t��Q
{,���}����S.��s���
7g0u�T1���H�7��\�"��ow�X/������Вk�2���M���s��i!a�n�55��G%m��ݟ�yj޵�m�ゐ�Jߞ2���\��u�f�('J�QI�lg�[%�ggƧIe�f��n��lW*Xt�r�*�#��'@V�ϭ�UfO����5���@�J���ԫ�d3�������YL�����������h�K��"Ss���� �z�:^vKLWdpk*`���t/�\[�d�=־����T�8uS�����I��.�u�[��h��@B�Ts_+��c2ug
��v��g5�Ih�d�q6�@�㱔�b����<�`%
8�_)�}]�Qk��Bo>�m'��,J��cxG ���@"�3v�,;��2E�\l*`	(���BN��V��}�Gy�w��F�ۋe�ܦL��b���5�������C�Jn�т��[���rwPuΕ=]q,
ō���ѥ�>}1��,^7�+�噦�(��yo��Vs�7qQ��
�R����YB�[QCB隵������Щ���oc�{뮾j����h��S�8�[�pS*Y.+x�r8�S�v�C]Ch�1,� ��Z�ug�@�����2W.�&V������z�Jݴ�.&������T`�RJd|7Xim�L�R�b�xjLݝZ�+�A��v�l�S�9O�D�5:���8K�Y�u����[�U�gy��L򾞅WjE����9X��m8}X��Z ��h~��ݮe`Y�7K�Lx�����	`���(R�[]&7O[��X�$�{W�öV�ҩ:�p-�cFU�v0$����K.ڶH\mű,5�Ύ�ݮ�#Z�%�V�P��),�ح*�������`Es4u��˘7���+:[�U����1� ���:��b픰�)��Z �yG\f�}�Q�H�n�l�&�)K罬�V�)�Pu�����!�I���9JŁ˞b����`&�����0�6�Gm�R�N�b	�:k�y$�C�E��H��2ew
��jj��~���ک-_bwQ��]tM��p�c����� 2rz~�Ut��iT�r����QL�R�L$�d� �ȶZ%El?�=B�r�jY�g#�XD�R�����@p�0�Qz+*�5FRuYDp��7+9��e�G"�k*�0���IhTQ$%9�]VU4�%ȋ���'$�
d�U�J��UP�0�^M#̢�TTTT"(�Þ���*�ԣ��$0�L�ad��s��Qr�B�����ʜ�E�T��`EW9Qȋ	
R��I�`I!UfJ��݈t%��AU*�
%J�
��TEJN"��94h�z�ug��Y�TUȱe%��tY�J�G""N�^dx���2���r�*9�-�A��T��j�)�V�l�?������L�"��Dx�r&S�i.ܮl3%0r�¦���7{Ғ����\^T� 7-�ٶ�t��G
)w3�3j�)D]l��G� ��т'���ǄE©���ȡ'�97��:�];��E I;:|�m�{��C���?����=��������.�|DDh�!�O�!c�>����J8�j׽�-��O��0}�}���DAm�ޏ~�1����oϾ�?_���]�?7Xz7ל�x�d�=�ϣ���ΌN�Ϝ8��SzNM��w���",}��} ��|G�J�&�_��%hOt�˼.���B�}CT�W�p�v�o�>����n�[�o��o�N���~P
o�$����_#��-�~�����p�s���{Nw�t{q��>��K�,Dh��������ˬ�a�UG�o7���у�}"#DE���"��D!���_p��@ }��M�NG����o�rs�?�����zq8�������zM�	�~o~vW��&������oi�z:�v��C��E�����_��aO��p���}��Y��v߮�p>��{w��7�/V����w���8����zL.����Ͼ�?�raw��<�E��s�oϽ��m�N��?>�b0DE�#�B�����F>�"57z�ʅC0��k�ج�qS3~�!��L&����߮������߯;��O[���v��C���c��П�ߛ��xw�bw�k�|����_i��]���mD��$||�7�@��">�c��j���hzD�"e�do.3��4}c�1����~����~�!����9�'�ߝ��aW{q�\���C����&_����z�w���C׿�߉�!:v�?���M�	=�<�o����ܗ��?=�ޮ���{3�Si/J��O��b>�ǎ{�w��o��N����q�}߽��?�����|��!��?���7q�aw�?]̟]�
���?�7�oG�w��P���o�y��#�#�"'sٞ���cw�Եr�g+D�ᷤ܄�q�_�	4�;�i0�^ݿ��ϟ<�]� {HOl~��{v�{߿{���zw+���ߎ�{B��,;�oם�tx����]�߇����z~1>��3��������Y<<�e9=���|�y�l�w��]��HN�{�����>�w�ޝ�}���©����������ߛ���w�i�����'��v��_���<��ʞo���*��T~���o��~+�/%�v��i���+��U��8]�}9��C3���ζe�}��b�ᠰ1<G)�����Ǒ�WY�����A��{v�G2��P���i�ҫ�N��=����:�%͓oכ�k�f�ۃ�$�+��O���=�cwc�=��������jTZ%��u��_����$}�?���Q���7ל�����x��ɾ�x<w�k�Ͼr�>�����9����x���'��޾����~�����8=|��e�����o�>{��c���������>�>���G�O�>�n+~ ����o���y�`���������Ɠ��<�����bO��������`�na������;a}օ�M.� �F�������@�b0DI��!����r��C�[��8�yw�nܛ�����7����y�ސ��z����{������~|�7����#���~�~?|��#�Kĝ~�ٱx��8�Y#�G�>BD}�=����M���{������]��(?S��C�z�PP�On�u�a�l�I��M���o�x�m��oO�Ο�G��}��ꏐ��@�=�R=�"�=�9�Q�f��h�|G��S���}�7��x����ۓ��q�M�O�}��/���;����O?}�:v��r�X�C�������tl�b$|�p�$G�}�^��
;qW��V�]ʝ�`���F�D{Z��#� =o>�oO��o�n��L�S�|��'�~�]�~��o��Н'��]�_��7���x�;s�#�<v���o��&$} |G�u{�v:}_�<�u�����Nq��p}<�7�'!�����;�]�|7�{�990��GϞ�ߎ���߷&����|����o�rs�>V<@�Iğ������~�rn@�#D}BG�|xo��;a����ef��ސ����C�o��߮����<�:w���+��~�����m�o��y7�������bw���}�<w�Ʌ��>q����qψr�ϼoP�O���������+�煥f�1{7��.#�|F&�	$��c��;���c��<L.�C֭�#~!ɇ�����w���叉�}v�yޓ������;z�����0�����}�o���1;�}�n���'�>�����VJy2��G��=��>�ѹ��}��&�>�ｇ�N���=F��S�r{q���0��{q�y���raO[���������Վ��~������'~�G睽;x��}�b\�Lؤ�}�>s.�O7�9�=t�3�R���>�9��W�E%wi�u�9֩�9�.�NI��X<��n�2�BkH� �]X������L�Lv��})����,EN\��զ��Tj�X(��Gu�o NXt���z ޶����#���;����~ӁM�=���zI���@~��ޝ������������;Hz��������Ӊ\!&������]���n��:?��OI���տ]��]�v�ǣ�>�G�"��u��Aqq#v��)�l��}�}�"D{�����}�y�>��ܛ����H}M/�����zC�a��?�?S��]�޾}��=�:w���&�B�o�r�	7�zy#"$ǄEi��������.8U�-�F�i^�ܥ~�CF���DP#�B#��G'���<We<��������|��;��7 I|��m���߶��>���I�S�=����_ѽ�������ܣ�|r�F��>�D����w�䷕��.{3�O��Ǿ���A}�b�P�#|w������w�bQ������<C����;To���޼�aT7�|����9�]��ￜ�}O�9>����oi&�>�#=��p�b"D}e��^VMw��w�F�����F����A_����@���8�Q�[�ۓ}BQ㷟i���<��<I����~~����'�����������}|��I�=8��W~~�M�>�!����x}���U�Yy�-Ń�?����S"�L������h~;�x�s����+�	7���S��P�������N�=G�<Oo�nq��^�����m�nb�}b ��8w���F�>���ַ�l/˖^p�5�8�}F���>#�>�'0zM�_-����Ҹ�]���ϝ��={�N���������;ێNq��u�aWe�G���&�=z�P��#��S>���x�����y@�F�>��]^ϥS���G�"$G� �J�޾F�C�~���y��ە��>�G��|v�y����nޓx��;��='�p)��9�v��_/;U���<O[�w�j�O�9L*���������߿�~�N{�N��s?T�u�B�/�}��jj�����'�_x��aw���}����� ~<��w������}��:	2�O_~����;�ߘ�������7���#�x�u8�݅I���p~�����Ѕ����^��Q�����G�|I��>�.I�M��Ӝ}q*��">b8D���T}h��G�Dl;�}�#�#�ɇ��ߨ;�}w�9?O�p+��'���zL>F�OϿ�~'��ې=%飬؟R�f��FW� GRܯ�M���O[��7��)�}�<��)+1�LW���d�5�X��;\&i�����Oe;���k�8���<�٧<�.v�{��7����w���|r=']����ʁ�4��-s��8�g���U}�=�߽�h���W_��s�۝�=��!ɥ��ꃓHH�����<w�i�V����~��{�x���o������S~����?}B�����7���;�s�ۻ�\}bG�!�H��K��{�^�J�r�O��aWe��I�I�տP������}���x�Ν��=��C��y�;_cx�;��m�#۷+�w��|���ƥ�D1�>�X���z���3F�&��L����TȬ�J���r;��������Ez��u�57ˏ�����$\]��O �����>������}��������/-�8#jɑ[}&U��?Ć�lݟ{�*7.��z�O}��M��m��P�r2e\b8LA�c�
�������h�m�����X2�^�����l�gZ��0���qZι�'TmFᯓ��8s�81���g���_k�MOQ��,�����/�R����2%Ҹ���c=��X啚���ǎ+�''E�Ͻ)�!�
�Ԇ�>��!p!�B����qJ@c 3��|����̭<��M��M�<�Eu�qg�Ǿ��-o�#����C>Wz+���� :hHxV�����3�5@�#1{��Sh���Q�~����( �Q3��\�t�z+g8߈��I���F��2v��j(qU�����M��jR�m-5�}5��F�p7�	��E�T'#�'����8���*a�����}ǎ�c)�'�vأ�d�÷Av�c�6��ѕY���a(��b�Uw+�Бˮ�w)�*����ɶ���v|�\�Dj����<9D0���p����d��pvP8M.:	:�.� �|E�i^���{X�iVy���T�����ĩ�椲���mCθB˜e�8
!7�oV׻2vS�d��^ǹV�Q8,	9�b��3�����,5�����:U��~Ȕ��55�����ض�v�hF8'��^��� ��edq�"�:��>t��p�iC{OX��U�q��P�@ޓ���o��UƇ�"�G�@h_��f�{.]�[�Dh�W�����W!�	���d��1��ۜ|��N����s㨅T�_�C����D$�������;>��/A��S����-C4�.�a;�
6�b z{�����S- �dң��loN�����N���7�/��$���MQ�2d�ͺ�3T6��c��d���r �r���-,��[������}+)
��i�޼�Y��1���M��ߛ�F�q�UG3q.Ǐ��B�4a�x@�\��xpJ8Le��wh�Bҧ���3��b�=��Z���z�O�,�Bn�5��rH�+A�Tj�NT������{%��:���m� ���ԵQ4�%�8����R��Q��v��J���r���RJ3�ե�rp�972�=3�HB��h��������35�{*�\n�RNp��X�ꯪ#�u�Ϻ�c���z9^��6�Nqd��Q_E@�릫�]9��{�^�-��$y�/8���gV��w�UH};)�a������ɣm�h�+�q���f�w��<O=��v��w�^��<rn( �l�����}�q	:��L�T��H������5zz����,KՓ�7���C�����X�v~|�2��|�"���p�59G�}}$�ʱnlE�����n7�.Ƹ,l��c~�!�a��]0n�eal�zZ����S}̅�:��&���n��<^ y�Z�x:J8.�^����L������t�c���̷��0M��Z@\�*cm�Z���L#���2��{��W�Q�93�K����>��^�5��SÜL�F98z�����p�����lTUu܀��x�����U�����������-R�b�NS��!���f���&��S� �g�����I�٭�}带��}~FW�R�H��F.5�BN�9�9���s�����z���Ru��"z!L*�ܶ�_�Z���Jչg֎a)��f��p�{r��'#�������1K���cV��`��`&���M	Ǉy�=�-����47���ǽm�w��%��4sN�U+G�ly��0���U��!�@ͤ#�P�3��\J�)���>�����38�,4#�'4���l�oOIu�7�pa�l��ցP�w��9sW�n>��,�y9�@�:�_�U2ꆼE\t<&sWi��hz�/�I���'���uA��{ӂ�=t�L�R��W�Y�Vڈ˯�������tu��\���*�7����'��L`���ZI;�̽@p�(]��?��Ս�x��*�an��/,�l�ni�v<���:[�Ҥ�랞,(p�+􆘋�n�3(9�lč��yt"�K' X|t��+���QC����.�d���R���R
$�xM�!�s0oae���H���T��Nxh���v�w5V�g�G�Ј��આ�To�J��@�,�=�����8�/h�6�.��G�ΞR7Q�8?Q=}�&~u.����}72�W�����t�`���qS�7M\)�Yۏj������[��Gm�3�/N	E���e��t�uM/
t�2�=2���������	c��ny%Z�m@�.����1]-.;f��G��EG�!ߛ^���M֘1�e��W1`y(�O����.�m-�P�G�\.�l���QP#�
���;�4.�m��c�3�(f�����b�D�ř,�a*��w�s��Bm*��
��8ܳV�ݩu(3N݆;�-X�[F�M�*ܛY����.(5q~�������\�v�ɫ�<ؘc/�Cۆ�礫�
P�x�0�̯��C\�]�X�sj�ɋyU��;��UP�.,�?Q�O5%��{D-7�ީi����U) oM}%]���V�����։�^���]�a�ϡ[Wpe��jf�-�#z;���w��r@���P�̎����:T��76�a�$���񂮄�	��m��6X��0Sn�u���R���C�1�0�,�~D�1��f��A�f��)�2�t�WǴ�u��2!�VY�/���t����
���.9��1��Ӿ+ȿ�DwXPR��E�=������U"�V�+��<�m�%X~k��/!�`s�"0	N�'�Rv����Ax��.�E�^�o�>�owy.;݇em��!����j�Na���`iy�6����D�酟+�F��ǌ�=��nv7��q��=��)���k˓�㚝 ���a���FF�3���ݫQ��P,�+��zLKM��~�>���	�O��#�����w��>���5�1K�׼KI�Z
e�K��d�^.��pnaK� ����v����@1�Q�w�S��a��6g���Vg-�m�^.��k�f�׈M��'3�JTth�SC�?��o�{�ſ,�����v]l
��J��po��^"�n��������v-����H�GL`�; dਓh�_OK'/��@^�puQ�N����¶��-�Z��*'�GP�q����7�E|�v!b�sXd0���د��|W��7�ly��};/W`/g�︔99�0�7�����G"���1�X(ec7~~;w��z=SW2ϙ[����� N�����q.�F\5��.ʐ�����2�?E,]��xY���x�cp��_gU0����!�w�'p��Ա�eh_#��	;�I�7�Tgn�r�!L�+�[YK~�o�@KPm[f���������!��\!q�2˫ކf֧t�zT��6�� �#����������R���R�.�i���Y[O�>-�k��\����
�d�(��
����]���;�|��ӗ�a�DZJ0�sX���!=�t�ʠ��}PЅi&����UFy�t�h�����4+tv����q�N���(8��V�9�f/�c%����=��WU���_�yy���<Z�w�nW]�Yot�����dZ�q
�9H�4��H�L⺥�p��a�݊�LVk8R���R� Ԩ` �ٯMNfUa��{��|��R�]ut��R���f`7�tրd=l�6��T5� ���U���s�XX�H^�g��6n����:��R}���">�1f�p{)���G:�\f-)�Km�ؘcG#�������hX�.S']�8���39��n}�>�\T�v���/��	:���"��ɓp۠'��ֿ������E�z�T���rw�&ԈӲ���E��;g�n��8�޼�\�P�g�%�ܸr��U�a":�\�o0嫬%!o��CL�g¦��C�c��1W����6�J�da�uOP!I��S:*jl���.�ԡ�a)嶯��,o�x5c�ʎW����mCY�"�{sk��ٛ���t��y��0�9��~��.�g�t��aX����[��֮�����6L/�A� ?�_\Y�P��?_l��:��k����x %�Y��N����g1ȼ��W(m�S��D=93�6��s��_;��W�ۆ��j��]�V�&׵{��H�f�5�%�a,�itUo�1}0�X�HS���nS+)�ڬQث�y�
����az�g��]�A�UE@��|�����]�~��{oǭ����N��[�A�N�,[�#��[k /X�ż���B�oe>]Em<��;i�6L3���M�L`G���	
%k�v��t˝V�I<�h<�/d�N�CJI�v�gQ��-���"[[\[���[���h��u='n���]4%�YT��Ђ�3Uh����B��8H����v�L^hy6K������)j`��xck�����Lٳ�Bwi��i=x�H��n�Ҽ��e� �cy��ъPچ�j)l��LN�D3e�K9kwb+�140�`ժ�,١NQ{��t⫳�ts��[E�M�v�6���鋔���j/��#�z�E��"x��<�.�j�"d8��J�-�,>�Ο��S��\tp����_a�l�L��d*�E�oc�gN��Wy�D����V}Ţg`6i��F[N����<�Wh_q��r;k]@�"D�|�d���3 5���}��b��ofg�'��C{C5�U8�؇Z00��P���Z푒��XŷgK(N7�yy�"��b�=�t橣[���Fn�5���b��jf�	tH�/��&�:޺��K�����&�
ނV���,�IP��Y��]bYq��v
�@!ŷ�|V� Yg��t��Ǻ�ۊ����x�gh��1���-��V=|��û+�M����9��J�O�[C,�B��42+�E !�F�jp��p+�;k�4�n�_6�j��<���6)�jD⹕t� $��i�NPC�@�5��&�f��]��4�N���F�QJ�,��e�8�E봌�y�23:�$0���GE������Y�8��U���N��셑|�jfnIZ'T��0Q:�����Q�!+ui���j��x+��r���)�VGX@���aGlH�W����v�w��u.�[(�+i�KC]2����"Dw�<}����=OpnYrS9)��:+�����ZjVP��[7M4��@7Y(��Ņ�r��V��W�/��N7tb����bcs��-8�Rl�Z\���Tz��϶]�C�+V_B����"g�v�����s9��+k��V���W���[�Q��T�7/��uo*Iv��f��4)�Q��ڛ���9o�-�:��M!�$�b���Ίb ���ن�Z��;#�"Q3y��vG��ᗴVsi��+[�[��$q�u�[�.,��C��z��®=ɛ��\��ȫFǓ6>S�c|N$^�m�)���V%��]dd�sX�nĞ�緧�m���r�#@S]��4���y������S��$f1L!CW$��I䔑��+̚QE,���C�{Ǜ��&�e*�kliRm*�I�gU*����,�ZE��L0[�nھ��͐$.\���T�i�c�v�kK�/�Tݡ*�fҖ$�%��q�[}�`�*�m?��֮��Z�0�_j�U�+��$Go9^�묩�B2y;�R�W[Q!nK����=3��376���t� U 
'�p�,���E\9��UEQ�2@�H*3 �Ȣ(�)ZT��+9�Rr��˕�E*��+�t�P�&PC�W��<�/72,#ir��U�.�D�r�9Ų5.�t9�*�I4�T2s�EPEedz�T�H��E�Qh����8Ze%��*�\"���H����W%Y"�W�S��r�J���ӗ΄�J� EyhP\�%HQEU��s��$UE�T�'��9DDG�^q�J���Prx�C�BjN�G+�Ȋ<�*�\4J""��.|�8AF�HKB*�$���z�\�9�:��W(��'�#dQȝf�%EU�A莥L�N��"�FDF�Dd�'9��aT�$��J
��Mgu��WT���ɕ�<�u�e^�N:��kH�^����t	j�[9�;/%F�n�g;N�ut�N�N:��u��5�ʙAX�O��>�#�8�X-�["��ęG�ER�8I��P@�R�R��%�B7�����Ͻ7݄橫?�)l��Q�sN����D}���;�.y��T/���em��@󹯬;�Wj���NS��u���#Y���J�� G�Vq��2Dۼ����ղ�t�����b���t��3�9v�m�s���%��m�Y�;f��>�����l�& #�2^3�gG��[�s!�M�W3Z{�r�/����Bޱ^|hY�D�{Uk0W���B6�ngw�Hv_�	'dB'd�X��i��V2�ΐ�1p��q�� 9k��@��3N�k��{���LF뿐&�zX�����V��&�dF�:e�r�����AȎ�OPɅ�'G�\ݛ�(C�U'&��I�gq=e�훼���N������(9ٸnb�sʑ��� �|F��-S{��a[(�Yv�{���g�C�`��Vc����C><5��c�����TH�F�EOߊ��+<}�B�&]D�]qc��.[=;upI�W�N)�r�:;����2�\r���ۅ��W���S7�аV{���Ղ/�r�t��jX�գ� v���v%��:�6��V�sX�K;�k6d�<{�8h>����������������^q{�k��A��x�Ձ�/>����{^�s `�q����u�M�v�kƺ����ʉ�Ee�q;~&��l���eJC��P��'��e����gP=��V���(�RlD�޽X�鿄X��EAn�Zh���re�Lzf����a~���x��s��J�-wM���?8=�EVCN�cA�4b���Ek��	��u:�aI�	{��e��U��c	�2��=�����epY2J5�d��zc�]i��8��_Z�]�{������Ϭ���.�D�����=ꍸOo�d�R ޜ9uR��f��:'Tp��~.�r�s*����xRSv�nH����e��Eэͱ5n�{k1s#����!�#N��n� ��(h�5�v��ة�f2͖-��e�&��1�ZM5(����&ڻ�hq'��� զ{S�W�X��3O�'��
��X��ow|vu;�yه��K���.����W�\H��

_�ȿ�Zbk��A�D�V�
�����-�W�n�k���@^[�8-��/��]ov$��}��Y��h� �BtD�����on��8$N�Pʦ1$��qgww�G7$�����o���w1�E�Ao
/8�C�:���:�Rwt�=BP���z��4W ����د�/	^���t7���}��Dc��Ȧ.��D~���Q�2^3,yDF0�DOT�;!i�/?�tu�/�wU�w�W+��X��A�->W"������0�7,/��=\>���5c���RȋW㏫ް��`��X��0�3\#�tƄ*I͎���b�Jd^)3���rv�n�����N�>�Y���}m�B��O���vcc���s]S��.*�id^	�u�#�0+/˲��	���\v������E�r�k�^�������������i�-N����܃�Nfۏؠ��� 	��0��O���qE�+�0�۴��Ko�{���[�G������7�/����m�p�k���8J�����8#��:b9pQX�KS]�E�PrOqu��@�@��J^��bs�-���˲�m�Βt�I�G8�ޒ)�J�=Q�����
3Y�H,�鋈!�w	�&j׹�i�pO��5>�t�쏷�+�M�,�ʽ�!���HP[���=�xW}j�Z��R�;옳��P�볷��>9	 ��ՙ���^h*]s��S\�x;{��H�n5��h��-p�Yy�;)uň�>�h���׶���=�c	4�;�g58�����b�\Ya>�2�F�g*��1<�M>593�>��}jVN�w&b΄����ꪨg)%/RB�A��V:�L�I`H��`4���/�J��Pb��Z�#<#�bw�fվpy�#�>���QD�� ��0�B �ewB�>�M�O//c�����E~wׅ���9ǆ���!7��҆�?_�Ѕi&��`s�&4;�7�y��uX9̭�i�;u�X����5hg�g�����mց�~�{F�����F����ȵ�cOO�)���x����Y�}�����Pۮ�5p�c ���(ۙ����CS4E
yU�-�f�O��tS����7�+�������JS&Kn@���BVn��gx(֫N��oZ׷N���U��8��C����������v&���N�WI�>�.�l�����ߺ�BP9��6�҃�����vѬ)ٱ�Fي��x;;F�j@�n7{������n'I������a���w���y���T>']�_vk��i߄1����:��Jw&nb���,9s��*|�Oa�����U�M|��`�g�ː�1r�/];�c�n�����|$-�p�o��n�����x�,*�~Ew��uw�Z}x�{����-�B���v!B�Owo:r�ck���auZǼU�	��{O4=��l��
vqP�`�oh�G�2O��Dɫ���5B^n�]G3�����=�l>ǭ�5Rŝ~��wx�EJ��|�������{\Y���d��a4;��G�:)�u.�^����W��\ʁ� ;��Zw_0��1��B�o(�V��hiQ�FvQ��0bgC��}1qJ@��v�1R�LVnS=����5N�ց�����֍x����*��¸:J8-���*�S����=�B���Cg�d$nA=�*w�ν��=HT�8I��P��|j^U�C��Y�i��?aԈ�w;���C��C2хd��c��I۸x2H��l�t	��P�`�z�]uoa�͜۳��|�b}q.]Gn^�q�j7f�d!8�J� �R�����3�<n�iG�3�V�9��[��$�"��v���q��D�<���c�K�uv��l�P�P�'r\ B"��3>)����R]l\71�d�%i�7��B��y=cm�m�N�I��<��b�!5�x�^1[f�ۓ��9����?-sR�#�b�Hx�:+<�:<��U,i��k�3�$���I�z�*{�[�j�5i����M��K�;=X�*��`��>���v@��j�j|���*D�>חY(ܝfbѕ�l-!7�V�.�T*���z�[C��j��0m���2�?�����=���h��UY�1�!����a�-r2���i��X/���]�/�Mы���?)<�y��E�MT���%w"�6C���+�����q� �t�z0����.n�BP�2n��3w��KH�T"�����W1_w*b/���b���ni�S�Ч���@��4�s3Jڕ�v7zW;��v�o(�N�TI�b�r[7�m��������c���s���$\�H�T~?V,�����Z6��tÂV�����M�y���t�LV>�e�@P%��{�},$��D�D�n���3��?<Wx}��p�̱���ș�8%�p��U��<�2��auy��3+R~���R�{�Ki�S��Ycn�����l������K��/
cӗ
>sS�ԩ�kw��D�����hD�ٝ���\5�tƴ�Y�+W�~�*����|Cѧ�:uk��n\+':dF?�7lc�0�_�i��礫��%\a&:+���$m�פ�=:�����1��T�G"ʣ��/C�,��=��{ԇ��D��3��%Y����P@uG*���z���6ͪ,ҽ��J�WW&{)=Zn�T`Πx9�E��� ���#�U��q�D��_`<Vu�iNVP2)�O���Z�ԉ�dv"wMry����'�ɔ�l�ю����Y��o1�47y?�ﾯ�����%r^Ǹ ��G ���;�\�a3�ڸ����R0�ҡ��P�܌��tr�;,;�ʦ��J/�Fb:�D��Y ;	W¾��8.+\���;l�/eἊ��3D��eAQy"�D8��t�6�X���@���g�1R�c/�҂�+��'���t�q�*�S���N���rɨm���:��O�`���
�F`�Q���]�)b�w|�y.�o��܍�3�nx���<���9c�W.OX2=�
0cB�*ăȫЩ��Q`7[zw��ש���MUɸ6X_#46���C㹀v��NEAO#�O�v���!�`�L�Ҵ�]EN{u��S�w�6�0mCuBF	�Q5����Q�F�B�ӿPY�)��s��Ts�	�O
?r0��b��sj����s�vm2u�:��UG��g4�c+�t�������T�9q�H
�k!��|�LYCq�Z��a���7�PE��m������xlc���W��ݧ���� g.��8(�ٷ��N�lЭp�29��0����W*ݼ�9k��R�r�� �Ꮥ��s|kYY������*�5JX��c폜b�[���c���R�D�5���X
3t< {�;�wFU%N�5��}y�5`ډ�t:�[���q��ұ�	'��������}�'�����v��"���C��{����=2���<�3�yT�E���xKm_��ݲT׫�W�=X��=�C=v"�"�O5/a�1
��\4nG�u�Q��mo�P��xZH#�%l��얺`֗]}Rai���v1U0�:d��,��0Z�3�V�� �����Z�OIX0m�tpUD΁��8FĖ9�$hMF'o�5%��4B��^�es�e9�G��IUS��@8/� �O �E`��}n6|n�����b�et�N��#�^�
�M�3uȸ�'J��q�*!:�!��ʀ��@L@1.�����K��/6��/�/P~�KWX�Hp�;�g�t7]��=w�&T���Fx�����J��z�܈�k�`y-�
�l�5q���	5h3��cFPۭ�cȫ�!<`�L������ǫ�f*Q�x�����㻐:�b��ƣ-*�M}��^D3Z!�3���+_.���r���h���"j�֏PG�h��<�`m����ϧ��5)L�7	���C�V2$���Wj�ʐ0����Ff�|����z�g[zUf��{�(V�[�[ν�}����Z�O���c��E^%���Jj�Yّ�UT#������U ���ɤjR�{1�x��qc�]Ae�}[���'R�
�Usrff��?z��~G?UU}_}V�5�~�'Xʬ_XkN��8��C��\�������b{�S��n�O�h@�H�{�B�v��T/���9�`�R1�scJ%�4T-Wm�X9�k�p7�<j�6P�NTP�4��mfrx.�f��;��FF�@V�:�`���6�Nqd�U����Sky��{��咗��0> e�lp��B8��c9����,�{72��@%�����C�^7�dC�6�v�oO��S*Kd�@��[8�����v���J{L�O��&]���vHibY��ܮܺ'&�;P�V���C�_dʁ� ��:L����aY|cv�'� �1�ʧ�A���FMzφ^#2|-��r'�V��ĩ�����(�eY�90��w��o;��P�@�9�������_(�t�u�W?�B�:J8>��_*c��$�n���f�Jl�X>$1��;Pڸ}�V������'��$�	&���Q��^��u�Q�%�C�.L`���-��Q�s��p�IE��b�*��XJ���A��C��'�nɣ�7dDtsw6)�����z_H0�$$�`�ٶ*[�:�»�o	��}9!k��WE�L�7�v9}�L�}w� ��h3e�Ǉ&���p3v�u����2,�{�@I �^�ҳaNB�ts���Y�J~�����-�����Z���T�/>yw��TO:w.�>:ܑ�Sق2��&�L�;��g�`���p�,�Ͱ �����7 �{2H�Ɩ�_��)t�d���96�����ӵW�`�#�_d�p�<��7,$��֌�ɠ*x�W%ic2KF����R]m�s1�Y���X�����\fțD�ցQ�<X�%D(�t���ʼc��O髼��VI.�}h#s�o_yX�ra��e�s1��Ȥ�a��'��?m��Jڌf�pλiu���'[/n����p��Wr.d9�nX�@~����62�� �F������RJ�ڻ��p��le��i��~��Vz�BN�E���fl�A��f$o8ʑ=G��˱����qj�L�Ǿ�{j�)鸣#E��9�Ԃ<5�'@C��~y~ZF�4e
UW}�%��@�������,�
��GAQ�X���J��@��3�)�nN�V��%���}I��^h�j�q;~&^?�y}Β�p.#�J�K�y��Wxf[����YBm����2����B�g�"�ǌAXyա����!��J�R����(���f�fj�"����nj�1���+e���k�ݑ�Ұ�����*EA���m�����x{�9�VPei���8(ՠ:P�9h4@�\�]���&��df�ǳT#��#*;�/�;S���ծ-Q��6�ybr�;z�n���\͵+�j��ߙCK�h�ʃ1P��(0v�:�g��^�svQ](	��{�6�,��B4ެ=�n�,���[����}-uLYI�>��ܧ%]�v%�+J��c�u�{��J���ϼ��{�� :�R7�wM��Y��#3���(6��$F�x6
zUޛz���YQ�2��:�8�W���X���gi^N=���ߢ,�z���?!�*�\�yi� �ֶ�'#��]�Ěw[�s���7�c+�7�aK0�gVT�#�lvϺ_pIw6�#�%`�CBS�|Uu��D/�\j�"jcq�3�g�m=<0^�!�;{�����o)ge�-��D��'��a��S���7�T磑��V�*��:y�V��2A�bȺ'G�"�T�V�X�m��X�﯍;��8������ޚ�5���u�R�4p=�:�n�_m�y��)ԝi��Z`Y�\Y|�L{�Y�-���t�<,�+�&T���[�HС?;��m��Cl��iT�KE��Gy|�z��Z��fڣ�A�6�f9>U�\�CF�u+��t,��
�j$�t�C��4Tժ��i� r�w*(��b[[���]�Թ���A���Nv62-#�d�Μ��0���y5oT�c���GTC���ܬ䬤�B��~"���������؇,�+^G��cJ�{Q�oL�[B�J
ͅ�-V-��ɺ��{��7��De�_J��Y:�)e���80��l88+�je=��W�����B�ư����x5`�b�N�Η��Q�����2�4u�P�WW���ٰl8V�VM���x5]�#5Ǟ��}٦�����n�p��މ%�Qsr����1BG���C��I���s8���`b��jQ7]٩�4�T�xӖ�p�{�=�<�n�,���=�Rj�/��9-��,�8��_`�h�P{6���n�,nd=$ck`H2`�0j��9j�j���<�ٱ�M��NB�ʃ���l�Sy�Z��1�J})V�t�S��&��q#���okP" Ƒ�f铐��[��{�1WAҵV�]�jQ{oko6ma۝�8�z��9�*���3�$�rTe�����$���y����h��\���tk�*�rR�]�x�X��j�B�wF�r�̚�u���Y�8�M��ӎ���f��h�;�c��1N&F6Vum�ڇfDx"���(���?��O�$7��]��a]N�2��#��͍B;u܆�������vT�ɬbWU����e-OU%r����}���z���$��r��P�z!r���'$u�U˔PhU����s(�K��BeT�Z�dr"yJ��%y%j3�
�tТ�m����̇4D�@���IZ<�]˝�8��r���m
TO\�<���x�0�aI�9��.jG8�,�·#�NU�Q�+3S%NW+�������TFIr�\���#t]MZW"��!" �!�wK%D�"�s-���Q4� \�\��+�
3Ԣ����\�����-("�'yr��h�z��"�Jםr�*8s�n�=]Ԣ� �#��V�NS�{'VD�'QMZ蜢�T'Zn�d�U�wR��6�
I�j;�eQ�fF�tH�K^0�3ZRdUTD�$iwy�/�6�S��"�G�>D�("��
�=ю���/�jh2DI����b��`ԝhbuc_8�ז������:��y:�,�.m�u*��󕗺L��L�?�����U��Sr6Ԛ[���e�O�n��wѾZ?1Rm��+O���:\����N�kXw���_!��.���lFE9l���pk#�1�au��س F����z���$퍈���Q���n�dgU��bV�>e��A�}N�|n%epY$�H�'��%$����Z���}�3�p7eDQ����3�eQ���zs��Y�{$</6xj�^���=�Bw~���s=�}I��'=��:F �>TH��eXL�;j� �=��)��0]C�r{eXk�Rd�Z0�Yk��f|)}(�1�����g�;�B�\;!Ӷ�m�j��|�k��T�_�<��s"�c���wv��L�j)�jߑ����1.(�s6��8ʇJ������A���e�c%�_F���� \�$���12t99��!٩��O�:GE$b\'H+�J�h���~��q-��� E���>�r����.�wA�k������6�D�[F��d�u�����\��
�`ah=V~�j8� ݞ]îr�\T�6��2�EuǪu�X�v��V�\w��z���g�u����]�Bɷ��"��հ���>u�V�tk��
Aw�k���)C����#❠�duZw
4���sf�w7f�T�i!�X|/\��]�s����?W�}�}T'��^�ڴr>����>)#��1�I���{1J{.�F���wI�"�����z�IT�%�FL�b8I�c��b#<]�s�	�O�k�_we{ENTpwV3oo��T	T|}S��S+]k.�ʝ�
�x
f�z�[�|�?�Vv0��G����,�7��י��w[F�F�*���ֲ���u�cY�.�3(�!��ћ:tA�bcv����eM��# {��q<�φK�g���x�s��{��h0;l|o��B�_�n��nN���lR���� =/K�����'��K�7>�������h1��Y�)�r�nJ�Ǩ Ǿ���~8+�5BG��:d�@�,n�3
%�c�=�@]�!2��#�7H���gd�E�'���E�D��qIQ��7��Y�Z��9�L"񕙺���T�t}�ذ��t�_w
.��Jٳ��_@"���B��]h��5��բ�^�i�v,9�}�%A��H�a�Ave˙B��v�o]��zOt���V�r�_+C88��괐��M��ᇴ��l�^t��MԽ�a#Zd��qR�K�I���K7�l��&�P����j�g.�qQ�u���+Ȱ�����0��$�{�[{J���`��M��}bS=Z"�sP	)����ﾮ�MKs,zl���\�B�܅���xι�8�]�����!���]�˕�����w��Gظ�M$�kle����4�"
�qյ�3`�l��a�y��Ac��9�j^�\iOKYm����9�q���Uٖ�[�t�Z6����u��j_d�j��B}F�I0z����s�u�v�F��#�1�.'�ف�h;��k;�'�~�Wc+h�]�/�	�a�X_s�k���s���;�����՜����ﮔ=޴v>3��j	��m2��m�8�J�w����=�>�o
i\��a��2H��T�V)l����vT�����n;��;�ˎ���g�渝�-����̎�}z�Ō����;>*y�[i>�y�R�l�̩�ܞ^�t���n�FZc�r�K��_aQъ3����D�!��A��7G&��OJ+��;֍�[i���<e"��@y���n�f���X�:�[��5�˛n�Ȯ���h��w�ZG���a�Im).W=��j�<\[�"�1X���zQ����۔fpo&���/�R�!pv��z���_(����E���U��U}E{���`�`i���yވ��ڡ4�P_����^$!�p**c]S���Kq"�\B�1���������Q��3WA��4���eJ�������e�i����b�t�_>F"��ޛڇ�����)�ˉ�FXzAl��.���n|�IYr}��]��Aũ�
`�$���K����}k���E�w�4��!o����uJR��klj�����wyH쭪~�q4��T��r�]�J_u��jX����D����o.����B��d*��u��ȋڪߧF7~K������n���uZ��@�%P��8;�G!:s��3WT����J욎���Ǝ���X�qw�TS�%F�����p�D�	���#�
��̜���>�'�򔬼>���ޞ�:�������\a�t���T�M�M�����W�e���(���w�`��QЛ�a^24��e\^ov��C*���ǋF�`��>����퐋
:7 �`��L5\GC��2*2��Nq&����
r�Fl�
.��R��Lñ��p�k���w��	�w��EPU�Ν���n��G�}��+�}�}�
�+�K9^-K(�������o�}ȟt`�����J��+ԫ/��1�-�2/n.�ͼ���/9�N��ێN5�9Lԓ�X�g��
9���g��cU=m��[|qc9?[3z�����ᨓ� �Z��"ť���n\Lʷ�q�V�c�Y���49e_��c?gW��eF�<&�f���H�d�����8tM�g�R�r�v�ެkg��v�WUĹ�B�XO
W��ҷjq���l-M��/���P��h9���qC�W�Tc���8�n�G:�S�1�oCYoS�i��Y�Ņ�D���tqu��y}���-���DI|�)*4�=�|�z�<�.o^]�{u�|�:�n�k"�?��r\�w	�.�ܽ���\�љ}����}�[��F�rpn�'�X�S�׫�EО�t'G�魶"��n����,m�F{�|���/�3��a��Vb���VH8Qqh�g��,6+xUb�����tm�Mm6�K�>J��t�lt���{�P��%��..�j���ZvfT/��6+%:��!f�pwl΂�7_<kL�X�Mj����W�W�}�����	��DqƵ=���2�"
_ћ�O����0a4��a�;���*94����8�o!�r�fx��mݺz��J�k�W�Jkop6�ټ�5#�˙��l��h�LBv�+g�uѠ7k��A�ǒ��Y����Q�k���MQ��&6�Z���b�%���"�.�.",��d��I�l����>Ӱ�_N�z�����[}���BS?k�=Q�t���3�69�uI����K�f+�C����|d ����Ã����X�֔�zS|��jt.��k^��dy�צ���ǂ�'�ds���^�:��b�`���^�r�%ݻ󝾷)Fnc��q7�`q\�|�r�u���9�V5��V;#�.8�ܱ�_l�\:����NOW���FP1D�w4��h��ֵA��V浓��jm��[�h�{�"n�������.�\,;2�[<gVa�g��w�[��;Ѯj���r|q���Y�iq�QR5�p�͍fl��*hR�ON�������Oe�覮�Ǌ�9;S(���5ܓ�+gH[��%�O�}�G�
w7�cKѠe��+ S�] �/��Q�k��)�kOa:0�2�^��q�o5�O0.��������
* >U'���b�����p"�
��{i�Gr��H�����Ol�n�XS��:`�0;��iu�PqK��ΰ���9<��9�.:ye�ֻ"���N[���zJ�����(M�Ԫ�nK��Sx�e*��>5_u�8�q��O�2� ���u˓x!��/[+%+��kn��1tae$ҿ��o��oa�s�cb��Y��Eh�͹�m���b����z�	쮌$����Ű�g��ɣ����T��{���@�X�ʷ��^9Gώ5S~�eO<u/b�:��t�8�kw= �
�_.�w�N����Cf-���2��ވ����n�s'�������IQ�����s��0��:b������pH��4�yE'vW�69���\n�urZ�)������>2g(p
�9�Ve���V�u��/���/=J5��"�;�f�ĝ�c���^��[�o���u%���gp,/:�3�U�v�u��r�t�#�W�g\�v*�|:��B��u��Z���UU}MzI<Jaa�Uܳ�^իJ^�bp�E�go������[�襏�^{�[�X�ɗ܌��ok��Q/Wku{\� �x9<|����m|���ߨ8O;��3׼��նFs��3�y���c�󲧜Z�[i>�q0�}���:���ͼ��w�3(��z�\�D�}_aQ����66����۝��W��{%�z/Q�.x��늱�X:��/�T.�_-�=7�mV�<���3m+o}������Bsʏ���v�	�a�!���w<��ۣ]��~ʉy^�]^��e��5��=��Я�@��hk.�w��6z��V��.ܝU܍AI����[P�Rt݋�r`�ɊSyϣ�^V���t*��OM��Yހ�="��5׽o�!�9�̉)�->��m�j^���k��3-�V�9r���-+�g5�K����b��ǕMnТ��z�-t|�nd���{�}z����D��u�4h�-5�� ���k�N�r�::�JÔݣ��y~뫨x*O�[��][��8�b>'x��Xu��
�/�R��Jr"�V騖��!�ܬ�u��?��ﾏ�v�4��-�s�T��q�Z�~dE�v�2�1��s�dz��]�W=%Y�5����?'njfb��ڪ=�Mt��,؉����p�.��X���	�I0�!���G"a8���G`-��_xt�Ԟ�;��juN��帗�7�6;�;���ӆi���g+\a�t+���Y!T��D���j�n�s*V-�Yەj�u��'�E�gm�����8�g�rfmu�.{r�x���[�ֽ[|���l�<~��r�jw�Z��]��{VmqDu�"�~Y��_�/��f�>�լj~�oRy��)%l�=�w-����u�5�:V.�N��^�F4�W;l�U����ίB���x��ӛŹ�۪��wh����[���ݶ��=ۑQW!��o~:z��&�[��Ff=�Ñ{`�p1!P�7�M4_=Ⳬ��[�7+�E.x�*�}�F��
�	a�c�:,�L�������m#���ٍ�PP���6���ʜmz�XB�|mP7�<WZ]�)ru멦�x�zt@��$���9�%�K�����}6&7�5ii��`�s^	�*�ڥk�}��}�]�kwM���@9�v������;����i�i�AY���^�E̎�����8pX��!�As�)TI|��J���|��uCeS��{�T���E�������~�&hJmٿH����r�ZP�=y��|�B�S�E�'�1�P��s)l����@��]3,4�jԸZ}�{a0��-��v�k����P�s.q�;��#y���E�9fmn��HpK6��6�&��b�m��snk�Y������N�Y٣1R�ʗ9�9���k�2���.5���L'lf�j�N���w�U�&�ޝ`���;rs�o&���w=i�=���m�1Y�zt5�%#��K��	��Y�&}k���x�Y?g?a�>Ӱ�S�eF�G�{�u�s׽/�|oX���:�~���վ���S}���g;e9�W�[�K9�+�^�t�GÜ����Vнq+�̮c&-�Q�{w��^�������-y��PRԷ9t�-wɁy����y�Y���`�;��ǇbI�/S�*��!X�&���i���w�B;�g��C��n���_%6��U�	���}֊��I�Ñ�B�G����AEA��ta�ڈ�5��&�6�h�KK&#o*�u�4`޼�(Ѐ�v�'���#�G�_
�v���ݻU�)�l�v��kD�G9�{X�Ee+�\��m
T��J�|��$�{���V.�]�FM��d�D*���Zf+����F���Md�Y1K3�\A95�:�2���۹��ڙ׬�E�V��V�;]I�t��*�f�������Nzw6�
�ܷ;��wH=o�#H��ֿ#����O&_
�6Z�0��t�=�]��l���X�Ý�ɻ�+x��������Q�%"ļui���n*k�Z�����
�.H��"�Hp;�fԥ�M�ns�w�������8uvR�������J�{�� :�Ոf�LL͝��V�q���R�;%�bML������-P������M�e�m����@�{̡锐���Lԃ�
˵���G���[cw�:�[H0*������?LtE�y�[�V�k :�-�-��� �u�]�_u-&�&[s�Z< 4��:Į�<E�*�����ʚ*��+�/���[�[h�"�iS��p#GW��G�3E����b��h�3��Y�h� �U�Z��!ȝ�O4*d��DoH+��&��G.���Z��vr�HK�켕�v�Gz�V��Q�暧Y�ɭ��˙K,$u�c6�����i�m���H�-�M4D�Y����c�<�]�RunTf���t��+��ʘ���.v]u)��o���ڜg=�bA��h�"���p6d}��wX�3$�U�*������2�Q�2���H��̾�q1ɺ��Ч��&Ҡ�Fc�劖}p�N�s�\�ܩ��aF�T�v%z���En*2C�3Նޚ�C�*�ZZ�'���,���M�[�@���o5���f���9��+�j�9�K��s��->�WwnΈ�-Tq��\�k�Vuz��/Z.�"�c�q���Ը�L?B��@2k�W�x��l�f�䲰ĒAi�X �m�UG}j���!�i?�nAP���i
׮ŗ2��k77�n��Cj��^��3N���[ʤG��c�y�=<��v�!}ۀ,�5YK�mV�<�ڰ�L��h*��ɡ����m��Bo�&G\�Ӆ�#P���[�6��nl����u�]U�f-^�U�i��M�'��[��G���p�޹���JC2��3��Z�'�[8|Z˧|�]��G aȱ*�⾢1��k����Ϟ"웢"�V��b<�K;u�8���zo�MF���� ��P��:{Wϧ�����Np��ؿ������A?YU<y�G�'/S!j�Aʢ�*\���v���˞o���;�w�>R�DC��Gt��R�ͯr&DUj�B��y$j<���J(��%�:TQ�����e$���$�0��w��/�M��e:h��C�:T�x�8jJ�*V�^��̇8�\���46G5":���c"N���ZhDy�����u�'"�v�U+-�����ȭ�--2:r��S��nr��B�haa!��T^�W �6��H�(Z�ʽ�j*�j��db����b��t�Շ:YD���z��;��W�%qۄ�E��V����wt8jZBa�iQd����=ՕP���/eA�f��c:��Fe̂�q"'
�ɗ��E|@��ݬ�D��g�]�@���Yuo�7��v��Q�|+!���@	����imT3 `a�=�$�"h�V��7xO꯾���9�u�p��t����w坸ǵI�N^��P_H�F�ڦ!,�qj*��ݼ�G���P��[��/��ֳ�o^��usyeAVVħ`�6¯o��+~�}=2�io�Z_aQ?E��Py��v��[��#E�M��z5���=���J�b\o��]�8�<\=���g����i��۱��Aʩ�Kz7��w��!]�b�|�z\��K���p5�_=f0\�Vc���0S��#;җu�yԻ
��d�0*��Q2�_ԕ��r��8X�V�4�ɽ3V�A����[P�{ecw�ۆ��dJݟ��#��D�����|�r��)�s��o/浮��9��齽��f��7o�u��~m/e%�wٝ��_W؟r���ۍ���x��Ϊ���6�-�*���c�n���r�w���*�w�v.8��l��Xm�i�)�R�Q!s��w������v��ޥW��Z5p�A��f�WT ��ބ�/l9� '!�K�wAVj��s%]�HU5󎳔�mݰ�@�0,쩅»k\�;oy�,��$�7OC��[��h���h!"Z��ILV���j�^�dv���+6�W�}��^��M�-�R�#m�Z��gL]�HOetgi.f�m�cbr4����rOz�Q�"�O�r']�P���tu_�k���5�{�j�΋]z�=��,j��k���M�>��qQ�f�[Aܕم;��Xr9���]��r=���µT�Rp�6�m}�s\Y���kb�U�qZȮ�蘇S��{�4�>u�6H=ϧ��\��䯹�Nk�wϜL,���ow+�<��Q6��^��N�y�R�\rz�O1���f��/��J���)w�pfQw�y�tb��|�⧜\)����J'�諮M�n&�M͸��x��v#�f:=h���uz?��GT3�re�O��k��$��Frv�o�|����/ݹQW!�����:�k���E��5���^���91KCY6�\�}egW˰��d�0)�y�.ږ�R'n��6@}�%��0�s� k�m�v��ʀX���N��\���X3y�#��T 0�k
O�*�@���}kd��n\����-Κ��ܴ�]#b/o/�rGP�j���*`V������I�A�����ͩ6�b�������Y�_u�[�������J�kyoCYoC������W����$�}L.)�a�S�U^�p{�`�9'��jkг��N[��nD+o"�����VM/�f�	D�]q�K�|{�r���q��Cc;�У���u��T�����@�삽ûC��u:J�n��O7N���u��Lբr���\��2�!��ѣO>��Z��5D�͞4ܛə�P���sFz��=�xy�b�]3�)ۚ�f~⺠m�Z�j.z���m�j΄�_��ԋ�O���l(��Ȕ��z��gų\�tI�X���6�ٗ�M�͎��5Fӆz!�����FF]kՙ=w�{Ӻ���c��W�f��k9��~��=�5����u�'ۖqjVgf��,��܀�Y��S�0�o�eZ�j���s��9�T��C�ϫ�9G���z�z����称GTjÛ�kz�C�9�Ѫ��b��Z2�k�������]���9��v[��n�lH��6
�i.����%ƛ���T�D����B�]���P�ǩ���uG�sҶiV��O�a�W��>�w&ӖT�Q���}��+9��n�^�#?�����-xfQ�H�U79Q=��j�&U��Kw�]�u�oq��qp���n��^�F;�ۅ�2�
���M�=+2�v��=��=��J7�A��޾�l9K�K��o{�须(r1m˂��a�uo�S��W��Y��u��a���Ă��*i��|�+�{I�ٳ�7ն�M�v>{��~�D���q�趛�z�i�i����d��K_�ӯ)!g7�^�?%v�G��D��R�������zC��ݨ������Y{ݸ�Ņ?/��
����iu��w�N��5.�W2�K5XQ�f�8K[���޺���??�4+��W����oe����E�����jn��{8���k�o�<g5�9�D'�}WZ��k�~䗫�_)�=fk>9�#��\q&�e�w��ب�6櫇����<��^5��tI;�g�Z-a�p�����Lo�S4BL���nRbᲷw�����40_,�<�+Ƀ�-K�^jt��Jz39�:4XIs��+o��u0��Ĵgu�����\4BE���%��V�)]o]Ǵ2-�;.^��y&#��G��y?�����IT��ov��	�SQ/rj>�N�R9\��m�l8ƅ�wK�P|5Q���5κ��U=�eX�*ޚ\p�qƢ���ߓTms�}�]<��^��	��!FoXO��wL��o��#g9���+�ϏAeo8N��k+uG��k��wԄ5�������y�����J\wY�'�܋�Nμ܉fͧ>��������pf�K�ϨA�n�*Op�)��-s%wd���|1k��\�.Ƥ���[ׯc�X�;o)��1F���h�V�}�9s�1��˅Di���u�6��9��3Ӿ\FL��)*R���þ���ʠ��O/�>�SU}(��=�힖S�n ��

�q��N��Mͽ{��5���p_���/��Qʑj�аaF7�j:�!-y���zH��r눟O;����X���9�Cy�>q�F*������:��7. Z'�l5����>�3$�Cl�n^����=~ǚ�[*N�]�U�����Wm*oT8�<Nv'դ�sƳ����n�r��W#y"�k+�޴��ޚ��Ǩ+#�B?eۊ��Yu+�r��1Q#3���)�j\����GYn�@�'�꯾��+�.]nV#�Ԟ�˃YoB�m=����;�	�z�	�Q����G��M�WW�[U��v��p�<�kZ��:������Xk��j��e�$��֨�Q�a�݉���+�>=_r�:�y��^&+������I��,˞7��oD-u�j���L^�����l��8+���g�͛�G]~����"�~���}5+s4'ы���s!�6�^�Vkg�&��C�9��#��0����6���=<�@ ���V5�z+~��w.zIF��&�]��D닎Cr-���0
�����eUmkr[�z��Oj#z��rz-8F�p6���}�0��c��ksr��C�� �=����k)5�;��c�ם�jҗ���6��oj��w������a+"�G�g�.�-T���zv�Gju{\�x9<|���K��Q�fF�߯2|�,W�]7K]�WX[�ձJ.�|k�K��u��o�O1�;�}I�+U���l���M*z��zZ�wE�֓;w�ީG4'���Z]�g����l��"�c�r_�s����n�@�����#�T�VP�S��괯�r�Ō���V��?O*_�a��㝞����Fu��6���:��b�*��Y�*TF�7v�X�R�m�x6MF��pC������ٟWz"�6��M���V��������P���;����-e�i����Vr�+k@ق�n;��:j�k{���a�D�d�{IR������=9����b�I`��d�=Zz�v�R�(�-��:�{����h5��-y��c�����i��n�\��>���.���r����oZ}v���
^���L�L�@.��ޟ�2�_��t��hw�0.:bdo�q�}��
�qƞ3�g5�9�D)����MJאk"�m�pgo��R�M�?���Ϛ�e�w�	�����"��6Ō���꽁\t)�W6�4�&�c�f]&�Uu��VX�f�[˙����(��w�t�]�\|.F��o�#;�u�Z�� ��-���U꒻l� �9Y;x%�9ԍۜy�ʔw;��ߒ.;��*Vܷ��iȎ��/f�:X��Y�ң������֛u��^v���"w2wy�ڑt�Q���eƻ����m3��Xc��<�x�T<�ǒ��:���\�ɨ�[]����Zp�6�]�8��.�Y�7M���[k.�.",_�[�5�[P�sc����5Z����NS�`V���|�.���J8��~�����)z?����s�S�+L��N��y����%[O����{����Z�̣���nr��2Gݻ\_�7�y�d��<��<��K�����l/�����ސ�2���OUte�+��|���sM���q��{c�<���)�@�w�K]��F��Q�1Z��.�}HR���4�ľ}qg5svձxr{1�Ҵh�76?���u_��Sэ>����Ɵv ��:�*����I[o�/;��1@�*|��)�oԕĞ���m����vЀ<�:6�/�9���Tyj���	WS��&˷�_�G/�6!�5@��#2���
:X�|��k�H���]�W	�^�M���J���V�%��W1Z��kj��ͬ��⎷vA9����sH;�N��a�&���Kmsx�E�]@H'����3'/Y����/���[K9hv�}���QP;��_�z�'��_Nsq�a
d�;���;c����gS�q̥w�����]5	�Z�ʼ������T�f���I-}�ZW3��>o�S�v�S�D)�D�
�LSQ{�׏�T��I{澹�Q��TBM&��)���9���\$=g�_yzrq�<ŵ�j��p��;S��H�G.f�|��Y��K��3Ur�����Ff�A�W=���`uq��".8g��9R~�mOLo��S�j�8��U����3����&9����S?g?aO�^y�ӊ����<XP���U��2�ہ��Ƹ���o��Fb�y�c2�Q����5.)���/�^�$���'����w�N�r���/��I1�b�=�c�Iki5�3�u�5(�c�eK�i=k9����w��q�f�ڍ>�ۘ���Mj��i�]$��S�P��ꧭP�]w��'.s$_e>ܣ�u�
k����,pV���
�����8�Õ夅��Mv�a��]+=9���Iu;��M]��S�������ئQ�n	����\䒐�B��}�E*��I���r3�\��Ss�)��*/�<�c%���nr�}Y;w��v����/9��UE\f��^���C�\uQ1��>���SDN_3%G[�gk@�U���z�ik�]�.��NG�Q��}��>���>1���+Rj��	e��}q->���vU�hQ_Ȏ뎕��̉PF^�������=�oR����=;���+��������Nc�r�!r#.��PU��R�5�j|3�q��黁a�K̫��j�Ъ�Wg�o�`fD�z�.������}��h�x��%��	��ɹI&�^ٽ�ԅ��E�ȯ*����N;I4���ԕ=y�:N
��z���E�A�{6��]�@O����)�F��>�ǜ���ɵ� %���߃�gv�D�lTB�z�]P:���}k�c���,Ok]L����� ]v�M��CU؏%
чV.��J�@��,AK�S�w}��Y�˖�4��&��n׊��r�j*��Vͅ$4:s�Ja|��3��Ndh�A�ѽ��.��v(�;�8��2��A+jŵ������ٙ���.1���s���mc� �v�K��/�qpdR�-�@�F]�m�[r	�k۟?p~�=@���D���<eN«}ҵ�����]��Y�,VO7�i�X.;��zf�^,�O�9���ќ���g����ф�/t��Ƀ��p�ΰ�j����2%��qT��maR5d\;v��>�/���(*n�v���ΈG�Cyr�e���R޲�]f������t�T�..��q�j�f�����j-Un��b�;E��Ұq�~�<�����Jp$ �em�Z�9�1��ۺ�/��ˋ��t�a���tw@�@�5M򧗮�:�T���*G�e>�|�TVs��U�An=GG�ѱ2O�z*�4��6�a�4ؐ6��*�%i���;�أ����ƫr����g6VY	'�k�c�r�q[��D�O�E��3��h�����v+ a�Kl�1q[�J��ݒv>��������z���@(�C�M1�c����A�������7a2��/�;�եKGQ��v�X���a
=OGCh�j�[Y�u-�i]�Z�Q�ۻ�uVܷn����w3in .�X�C3)�J����f����U����V���y�����x���bv	�3sr�r�ι�]b���m��iz����S�������#�<��u}�	U���lԹ'�,`�I�`<Er���x
���r��4���%iumu�d���t*]y�.�oP����"J�u�Tg��=x��'�>T����9��uwiݣ9#�19�:A�L�2:r��-Wt���BR,5{��gc�	�EC8������4w�_,q@ԫ�ٟ"�-����.�m��|����*�5��AwM�r�.�h��s��3���ۋ$���}b���L�{��/VR���%��h{��e�̅ʳ�;x�
�or�̻�\/-��P�(�{~t�_99��cS�̘9�&�W��;��Daq�*5+����_L�0�wm��D�`+�'��ъ��[ݺ�-K��MN>�k���L�=;8-p��w�>�u��**GvL^��ݠ�U�r�X�ִ�ŤƗ7���4In���\�gv
|A��v.�֪D�-�CP���������*���5Z~���y�m	��f5i�#݁�v�����v4Ͷu�_;�����忖�D�G���͡2�����J��[�j�Y�LwI���Yk�7��\M���m�&�De֌G��I��c�j�h�cw��� �^���x�Fƥv"P���S%_9v�m�ۊK�9��MX�c'>��k��/�3lJ˕9��o<�+B�Ȝ�^��`P(U�����s����g�kJ�č�V��y��UR�9������Ts�R�wvm�K(�����2C�r�BT��:+s�D�֧C1��z�,�7W%�'uȉ$����2wd��
� �S�S���D��p��<�IM���Et59�ʨ��q�rJ�;������酡F�S�w'8Gr��d���[�����
]s��Eh�Xx���KDu��OC�InA�]h��s�9j1EK��G;�U$J���He���5:�,�s���Uy��-$�����99u�Ou��$4w+�]�ۗ�Lug��\��%E+G]֜�T����)/J"�IM����,Ԭuʼ9	�p�6�L�<�%����#�g���I�.Z�:JUZsnHzP䞋�瓸���
w���x"��.y�&�YjD��*�bgC��kUt]dK0��B���m3R�:r�4L�r�]S0�U'IP��A&�"0���нY���H�#���ӻ9J�oh]6!xp��9-u��'T�8�t���.k�4�����lt�Ĺk�V�n�~��y��p[.��f.;��5	&|��v�D닉��6F-�E��[����c[R���tk��ףs
˗��mF�[�N�Zp�Cn�s��q�LF����Sc/0�]ZSӽk5�u��eD�{y�of�E㏱8f��L���,�9��Ee���SN=>�ō3�_��3D�ꕃ+�:���pT��>�o*���\}���!Ցe�H�g������>8�����}Q�z����Ekknp��=��g*�:ֿy�~O����]�}�������H�*y��~׋e9�۪�cz'�m62!�j���=8�Y���ڰ�z<)w�D��Kw\�o`/��
���m>/���gR�31]�w0H�r�y�E���5��;�$���+��T����5�Cچ�ۂ��l&�WuB�(ƒ��^����}u��#PRym�ޅ��}4���7nS|0,�+Wv�&1��>F�謧��G��[d�.Ҽt�j���:$�(��<�P�C^f�j����L�O���W�i�\s�A#��rv�dݹݘ&d�.;��T�4��s�%ˋf�WD:���Id��Λ�G�O��M���(׹R��x(ДO����K�S�_9��!)j�����ţ;�O[��~�a�.&Ez�W�s�v��u���+�ҥU�Ҝ"��/N�p�kY�
��~o����tcA�3�d�}��������8%��K�K��e�l[	��	ۚ�Y���X��Dry�w��!���F�[r�{&���ԋ���I���]/K�Ɬ���W���[�K���PO�^Pۓۙr�M^-����������(�l��K4�j�	�b�"cX���i����l�s����i�eww�i0�ؔ��ovu��q��Ȯ&a����=&z�[�V�[|k��v�'=��f7m7��ډ������ypӍw�e~x���Z�0���܊��+"^}qix��e�R�w�˞�P�lOі�y�)x���}��'���t9E�\�Y�B���O=YO�E�[�(	×�*���j*f���WW�ll	�#re��E���B�B�D9j:W{�n]���x���ޏ-^M�;�2�V��9�Τ�k�^`�E���{�j����٪����5�AR��p%?���������B�i�Y�.���t_.y��:m\K��oz����_l��f��zT���}��n�2�,J�W�p1!_-M�SM\�}�ݍ��/r��Ǡ�!?}������ʁ��F��<S�1��5w.3g5t�,ve��)����ݸ��V,)Z�*��I|����5i�Ui�O��хt���T|�`V�P��邠��!���!�l�b��C��5n:��/�Rֻ>|3���:�6��&Ex�6d�y�1��}OQ����>�����J�g5�{��8�S�w��E0�-Y�;Y�������Sq�e�J���*i[/��q��A�ҁ硽�|�O	�B�R���E�z�nNj}�����o����q�M��ɫ
Ft��9��b�[=PyoH��|g��9R~�A�`���n��aޯY��.�v�%uk���5�Q����-u�ȣ�]S���R}N���na�=�Vu��s���34�IP��j���.��rvsj�k��F]����,�D
{�o��|mN���+3v��{2�6�i^�fY����\����Y>��of7��8Ma�w0i7�!ʍq�r���n��̩X��xFe�ѥ�uyy�X㓮��j$qEq�t���1P�j6�3@�i�2����޹�W���ڵp������מY��Ƕ���â�TE,�M�����Y\F�����J��ڢk;��ค��s�'���ٷC�W]Y�����T��z��T}hzsV������*��Q���\�ֆ�/f�~��(�����?�ߢ,��ڴ���į5U���"��	���"���/�����&�4��E;Ӌx���
eQxe9Sp@���1iɬ�	���-_1ɊZ�����+:�aU�hP|�i�͛���K1nݹ�j������_�B�m=�+�����9��0�u�Т�Ld?����i;���RҊw�ֵ��gT<㔝6aԨ�Y��� Q���Q4�au���}�ua�.e�*�~V�����Y�����\1Z�<�r7Rh���	+],=�C�[6�^�Äކ��j���-�8=؂GM�	�f�Q�ٵ����u��΍8���y:��,E�ߩ�v����{�9�38���۲v@n$o>��+�1>4��!o�����5���ӛ�����~�ŠL�.���T����I�k�s��gl�*�9]�#�����(��UZ�By��!<��nP��љ���9Il]��4㻑��|��0�Ȕ�V�T�:�
�4�M]ܢC���JΉ떗mF�.��4�`�n5�q��.&#��Z��d�i�Y�@���+Z�. ��JY5x����'&��)(��9Z��t�ǚ��Wַ�N)#ו3��ȗ�sVe�$����ᚷL��o5m��Bh��*{�XJ�}��Yo�!~�3D���V��N�k�Eؕ�J�{��.���z_[�<&e[�Cj1�W7��2��M�c�(Yw�q�K �E�b�cN���7��=:��r��w��sި�'���drϬl5��+���V�V��WI�<&�����U�8,覽�Yn��)igf���X�����i�S�h�R����^�X�=��^��	���r���z1�ޜ�!n�>^D]16�n���6�es�q`bf�
3&-B1I�����s
^O������6ΓW/�m�U�l�Վꏊ��"�Ҿj��w�C�(m���}_a�щ�����O��|�+��T��V�յuu� *�Y٫�Z�����i*V5��zˇ��Ci���\e$GRw���Mہcw@Y�Pb�Q%";��%��O-�֖v3aV����������)E�\AP`%�iu�nG�y�@v���N@:~E���s;��t�Vr�d�f��R)�{V��|:�(]�z��������qmC�6�3Z�wCl�C�sP�S�P���Yݔ�v�=fk>��vۓ:1�?O\A6q�l�'Nqj���ᭅ�u�M�n�� *����_d��ڑi�����иwݯ�33��.NuP\DT=�r��+��2�<��[]����p�#���e�u�|k3]ԓim`�]`�]]�Bŉ��4�B�5������-��*�ĝf%\z}�m)[�ծ�}��\j�T��n��P��F�dT8�Ɲ���	��BA�TދA*�3�3��G&�WI�{�客>��
�"�d
"��5��n�W���
339Z�����kkᖋ��X��5mF�Z���N�w(9��	���s�m�/k��g����G�*���/3�s�R�[�U���vVH����ո^��_����V��,���nT?[����et��]�x�X�
��[�ܥy|��eB�k�G\z�t}^�6��}�zT��>xH��$���{V�c�Q��G���Q�\w��y�t�/�7���] E+��ji���Ѯ7HʛucAW0��d�]_a��1!_-M�SM\^e+���pM�η�8�H����+�!��a̢<��)΂G[�z8e�L��엨oq#;�\�姷g+�aJ�6J��!,�/��̹$nK��;�'eS���_ړ�\��-��rۂ�a/�����p��ݬ�q��i��ef)�6b>��϶�E�υ�<g*RV,)﷨87�F��7�E�1��+)���W\�U�g�b�Z#N��Qy��GطP�������,��|�G��%�Xn�r�+��LS�l��YG˾|:�n�_:��3S�A�M��\F=r)�rZ�z#�/%ͻ#6 NPa��R���~������g\p��ݱPw��k�-+g5�|�h���s��vDmݝ��N?W2���|�k��#�/u9�쉥p����3J��=�Y��t��y��Yx���������{|�˷��=H�r�D�U>�;���|[Dޒ�sG�Z�v�B�z�}WV��s�lU&����m�{UR�BJ��`�6�|��}H\��������� Ҕ�'�3d�Hh����kz����׉�6���b�p�^�[S�v�]���b��5q���ܼx�d�P�����^2���_'y9@L<0�ر��Vv�q����pVO�1TM�+��ڢ~�|� �x-'�d����${�;���~���Lx1y�x�pf��ӝ+X�xGXz�\����z�9۬e=D�7О��,E��b��_�r"�3��W�V{!ίG~���h��0YL����RV�K8]F�g+��.��ul�	�p[�9:�ՙ�H�w0�Z�[�7���f0��1ҥԎ}���ˤ�Fv�8���	�����"���r�V�up����}�RƜ4I!|`�rR<��e�h����(����:�^���=^���-�E2������{��2��:��
���)��9[�
.\j���kb��kOT��s��;w�:�ۯg��M��g�X��)9���%F�7��5�B�m=������o�(uꞾp�VV�l�lO�'��KN�O-�k��Χ�pB�12`Z�nZ�t���XŎߵ�Ap`%7�M�]X�r���ۚ���M�)�~���ޫ�d9����d@KD-u�j��cr�rYaWݴ��Bk1�ƞD3�y���"�����[�R*�͉Z�ypy*��c֎���5�o��q���D'lR�z�|-�z�/y[�ؒ}��|�ӯ=Y����mo"��5	&Bn5�9��x�
͞��DUjf�'jr��4�����M^-��z�\rtjӄk����8⁞�	Q)6��n��%��G��`����@\.�l�Ҽ���n��d�֍z��ΟjL�潻�f*a�[�
\��8.�v��-l��EreM֋Mp
&���)Rg���0pu�wb+Vt��TUn���*�%���u��f4�R+w�ȷa��i��*1t���e�������͎~i���]���vhM㪹{�F=�y�C�dJ8�����x���/GV�^��������nI�^6���um�/X����i�离���c�}~|qc�)qHdbT�� v���x�s�3u�+��.�?G�9����y���hrϬl�T���Mn"y��E���ͧŏT6��F��4_fl7������ԕ�Pyj��vO>�nq�ޘ�@/[�.Ta�����[i��K��Vt��닥 f�W.ǯIz4n���:�=�2�JR���e�r�;!�_JZS@\�+m���A�� �?ʤ�Q{��RXk��)˹���_.�q"�>amB�8����_od�_4���wfZh�[�Ԫڒ�8�çy4q��c:��9_C�SH�1�oI�BZ3��XE��^�^�����t,
�֍��xMC3{u��u�턷.E�H����v�j�u>�+Fҥ0i��R��ﲁ�\�Ƶ��6�-&t�_�i��i��R �� �,�2Z97�S`�h���R���6����f��AQ�o3�& �F�d$��J�]L����D֮��6V�z�V��
��l+��g1�� �#���e��XZd�絭����HT�m���0Rs��+	h[�(�fM?\
����(��&V�{�GZ��g:2*˭:,�r�%�_M�u�;�(i@�	�s�>7RM4pۻl'+���T�h�6�l�q�k���س5
�	s�E���t��_l떸֚Uְ՗�ֽ��'��z�@�w$�WW��:oQ�u�B�ܯj+��k�`��-������@,[��溆l��W����Y4-Xަ*�O��Yxv�KJ@ޡoFVgڸ��Z* �=h�F�h�n_%�:=紐�/^������}��T�N�.��8B�ع�]n�p��BH��j�(V>�9쓱A���BLU��5��D
�F�0�na���U���:��ݕC:����'�ͮ�q�gEN���j1�&6�vwpP%g��+ �N��r��k�Ȋ��E<��n�a�e����� �. ��Ӥ�YV�ĵph�2#n��*�k�����	�"Ft��YB���	;�<w�h��4�ٛ��X�ৣ�y[<i�^l�����0�N�i��	�p}o6��,'q�e���m\ٴ;e��v�M*Xʗb(в�]"w������J��{vn�MVax��� ��7N�k��f�JY�=tα��� �@3��2[��.	-a*A\i���/��*��9�4�Y�&���x��o��e.���P��s'Q��Ӕ�O�N#Ś��f���0��BQ�I�J>���
9zۺŃ8�t�6�Ġ�ھ��Ğ �u3o\�S��y�Œlj}�Vrh�ȠX����]G);��k,p�A�hL]-�����(�'��˒���'W	q[�KQZtV�.<{�m�J��oaK�ݬ�Y�e[��֜Kw���%B� 	|��|��[���ZN5(,mʓL=�j��*^>J�q�,t]b��]&t�s��U%�U���^K�y�'mp�%Ͽ{�y�u�Qc�<U1�D.�۽hE;4�;�:[�/�;6�ⷖ���&<j�
몽�:ϽĎ��7���'�|i�E�h`�[[v��to�E7�X8�/�tL��_45�%�E4�R�oU�gTL���{[����(�����{S��u������<�KP�:<!�W�5����]���tT��,�������j=��Q��L��װ�shmb�e���:�S�*��/�xI�eb��Lju��f�~��������c~�(в�*�HЉTV��U��^!dQ�:����I
�b��v����UI!*�����W�t�DU�R+�r���R-+*0JΫL��dh\��J�;w\��:u�s]J;�IȪ�(�;���'�T�Yģ9��C�Q��Ii�UE�Ie*2���åS���Q:*�aFpĩB-d�Z��wC2C
���B���͑)+4-]��$��H�F瞙f�|I��F�u��Rl�s�usn��:�U�y�*"�
13
L4)6UR����B3$V��Q�Q\�V�"8��眪�V���E���Էqܬ���$����9�wTH�U� �yNsM�9(�),ʝh딣���u�"�0��=N�z�^DR����*�s���:=zrW<���r%RunIG��SK2�2�9�f�L�R!V�.�y�$2���Jun�i�+rZ�T�h�J��+3����A�B�U @	�)�ݝ��k�jNh�����e�CP�O���Aq�h黏�<��9k���y���=ā�]�}�o2~��ƭ^ؒJ��\�*s�|��Qi1x���)�u̹�B������U7���P[v��J8hg�澜ז9���K��e�v�0���푘�f�������rQ�<ž�X~zJ뜎��R.�>�P�a�2�]���LU�q`�!�f6eO^I�q}��hڈ�̸��j/�;}	�8��u�i5~��A�/l��E�Zw�Wd�y�c�ŎI	`�R�BX�5˓u��1�V�Pd0w��գ;��u�u���?"G|r�9���	i>���eWeǷ�vp�ma�9�V\k���[����۾L�m���S������؅��t}^�6�����>M�������6Wm��Qx�M�T�}XTM��G�lc��}�n�Q4W�vL�fc�^�5�����}����*�T|^Q����Z��Y�ؘ5fxE��04�����έk���Z�Ee����1i���ch6 笕ٕg��q��땒W*����o��j����=Y)$�s���Xn���p�|*ͅ������E3nv�}y����֥&\�xn�!�
r�nt�g��*��Tcoh{�T|b�V���#�>2���d]��*�^�]�r/7�Ӝ;&�4�y�=/�2���,)��h�y�DIA��Y+=o�Vj羸=��m�IQ��on���ڇ�����XR�ޘ*�R3r�6���$Fe뎺n�>��/��-k�!�Χ��:�����vQ���7[&�����[r��=�Э}�ZW�k܆�E<gM��� ��W"��ѽG�!l���WH}o���J�qĚI�����D����R����ob�m�|�3B��ek���=����q������r��:�ak��2�]��D���P���_T�q�3�T���خ�|`]���M����t�ƥ�i�5��`�n5�#9Q�0ۖ��,�����~�)�1���Y��{�yٝ4�ܝu�pͷ7��+�q��5����@��b�t_6�)��/�84d�oM��Pe�m$��ٺ �?J�CLd[�Y˚� ^ݚ���4�gT�tp�#Dc|
�O��$�b�u�2��ڵv�\i��'���F�Ir\8��|��)��I]X�s/.E0��ur�c�	����ޖ�I$��1,y9Sp-�Q�_o?:՛6C��Խq�Y�y8Q��ةZj$KO�!\�x�2�r�_L�m�����&޵K�p���Wf9�BB�M���4B��;����ƹ�dr����\�:��j��x��0��=�'��g'~�Ύzrt��}ވ�ͷ�T&���%y��-�]Y}t�b]�1����Ui���r��j����j�ƶz���~T��C�9\�o�����D���ԙ�3���C�;�\��}p�>V��W�P��qg�nA�,��7��ޅ��= ��*�_�RӜ���޿_�!���~#���h☇m�z��J��u�b�U�Y���"�ߎ|Βz��"E�]�Y���vzjz���ʞ�7�!���d�e���*z���>���,�d�i��A�p'�� 8�]�4o_��߫�f0~�UPF�ِ�)��m�/�B�!���T���ݱW�.k�@M|H�����ϑ�h뗵&8�<S�f��k[Z}��Y�DpP�/u�(ҥ��o*���X�<��WV�t��Z7�7�<�3�py�D:�P�C�-E�F"=�(�.��&�d�p����w�z����^�{���4��U>�kW(Pŋ^I�I��J�Q�M�����]%g�ի��M���%�Ԥ�x7T�*�mߦo�N0o������=$L�Ro�����|��8>���u�h��Gv۠�z�L�3Z?Vx�q'Ҧ���SV�#
s�ӆ��N[���x�d��ӭ@͞�@視���R��Ћ��b��ΜO�p0�Ǚ@٘hUڵ��6��5�z&�ߺOx\ǶY�����dW��j�i���w���y���g3=Up�9����/��
��!�>Լn��m���=L?NT?_�I�,�*y��}>��+����%��k�W��Լw��{��9�O�q���f���x���S/D�Q�t�4�@!q��c-�����F�1g��5j��R��%�3��ϟR�f�5��wXF-�!u]��t���(`&�7�ꦥվ�JeOar�D#�7T/}.ix��C�V��xc��Ҽu4kӟr�����r��\nb[��3|����^�Tx\R��7�̱;q��N�a�N�1�^�{����'ȝ�^ߡ\�&V����,d�+'3�	%���2�L��ϴ�`����{��<ೲ��=@�ځ����V�g�p���]��f�{�]�X4�l��Bݴ�L�j��b���f�@�`�d����f���K����<Opm3�g'Y�.����o;���'�Wy"�D�YQS�[Anŕ��1��*&����oe�X�-��6`����{wjx�Y�OW�a�
�3�H�T�'�[yb@�z�g�O�ޘ��͡�4`&}���y���y;aq���Ie�$���8ʡ�l�(/���v>�27�l�,g�֓��UE��A��?Q���U#_��<��[ S�X�n�T@��W@c��U��J�Ѫ��s����1O�.�FGU&7��0{ZwR�پndj���*�M9��w�/��*��8�ç#C����]�}��ÝW�۸�[���U��=uͿ�*����bo7wk�=��Q��Nh\^ad�9��v�J���������3�T����wpo�����5���5	)�G�: N���1Oődv�7������G���m��>�-�������>#:G���Ɓ_w�.B�rz����1]�ψ��c���V�>|��U�ǹ;���8�fg��ۙ�y��8WR�L���d��e!qr���a�_��35᾵b�`^6a8��w�!s3.��;.k�߲�X�������`e9ۉT��	���ں��(�N\IS�����M��d;6R�u�okD1��Y����ᔏlWw&�q�r�ީ>Ʒ7'�,�76�`_ ���('*TjST�BP֩�O�:�5T
�+;o�+keb�1ԧNt�#Of֋�6�]�զfV��]G3���B�^;����� �!�-Ќ���s}U�=������~��,~98~��_�?%��9�<�U�X�G�O�A�!Mh�1F��ɴ�!���q=L�8l����Dy� w�_���5*�L�~��Q�f�K�d֛�r��`n'hq+���w�M����ʓ���gS�;v��8��/|���������s�z������x,����9�=F ������%�)�E�A��Z%��L���O�)�+Lu��_�tN����Cb��>P�[�������>/s�����R��y��$�L�#�a�^��N �_�����O}�s��W�Ϣת��k�~���������w��0�FH�z�_f׆��ε�TJ����΃�>ܳ�c�vM��eNGw����`���'n=wl��վv߸.�hew�5#���ŕ �A�:A��HyM�,+}�Cӌ���t�n|���2F�yC��=o��(�������W~���2Q�D( p��]FC��0ӈֲF���;`�a?=���fP:r���i��P��q�/%�-V�8R�&�NEQ�z�����)m�;s���`�K��=�G��������ف�j�Ӕ�`˝�Y7M�b�ᕹ˫2�͆�n�8��yŵ�5:�x�F�B`ͮw�&TF����W��v��<ƶ}33�"�>��d���A}>����q�p�_ؙ�����]~��ꏢ�	+rn�HxO��ր�u�u�ze����X�*��n�!�D���bl���0a����<�ÿ�����`P�ٙ��5Co�CfM|�SG%�T�zzD2�G)\b���b��,1������E�-�
͞C��ˎ��w�1s��\c�#�ٕ~fP���ދ�
�����1�fӠ!����]KӢY�s~ͤ=y�x�n���JuН+O�r<�S72�\dy�`g������J�C�	��΃���`
��+�ȗ^��Gg=w;W���+g`A���FW���Nq�e&�b��P_T)ɝ;E�����	��Ƃ�Q�P/��¤�ĺ�>}B�F>��	{i�u�VD\�(i.��Ez�|.zc��97<���J���Q��U���fd��2���1���^�}��Դl�^�O�];�1B��4��^�V6S�L�c���T���.E��!�7\��}p� qZ.8j½wH��_��N��ҭ�lv�Uhֹ���)"U�����9ӮM(�Ĵ�ヒۊ��'|4fp�v̂�ε��n34�[s4C���ɽ(���Gm��Rq��7�M�����\%i���=*í��gS's��pp����w���¦mvA��$�b�ԅ�KNi��=����<���Ͻ�Y���Ǹ_uHMW��=��7Ht�g�I�_q�O� π�"E|}-�ϭ]A��7�$:�r|����V�緎�{f}�<<1�t����Ǣ���DTf	��G�x�Ba��_�ī�Z���75�a���Ƨ�+t'�����������uP�@H��-�`�>�\^���È��CA�����R���Bzz��w����^*E�ۿL��`��:N��>w��zg����]�pv���~��{�J�+�Z3�W��_�'/��h�X�����mN�=ꧤ�=3h��GWvH���x䘯W����C}�Ի�t"���b������;Y}�ۥ�յ�\G��=�.N�]َ���џS�i���c�UXc�?]ȸ��g}'��b�y灠;�l�\Nw�jA���L>�;��w�z}ٽlp���a���!q��w�*^�MxgE V�3®1��^��o����+>�0�FK�cv��O���2��]TW�Eԯ=N1�,�w�+��cZW�]=S����:Vz��_MpԆ	Fl*һ|�_eK�9	�+�[���ݛ]�4�t^�b���4�sW	)�G`��Vv��7�� 8S�*��QyE�ܩt�Ek������*;Wd��]�=vZ�}�^��������v��r)���\��-v`z�Y鿣�B��RW]��Jz�S=�9��v���V,��y���p���ĝ]�>���L��YLjm\n�g��xiOG*,��I�;��=�|:��;�g���;GD��)�`+���<Ð�wA{q�cw��W̭Ǐ�6�P£t��VE�'}pe��g����w�rWf��iv��z�܏z���)B�Jm�{Kr�/=)4���Au�ť�,�Y�OW�a������H�UO�y�[yb��GXT1Nɐπ���ڢSx3��W��_��Ǹ佤Y,�3ĕFa����C��2ٺ�Ax�N�ۥ����`[~�[�VV[�u�|�}����>�������߇�%�|��j$�'��@Q7cѸ{W>�W�OK�};�����g��U�˽��c��7A������٫�̂�|��+ц/:p~^�=���Q��w�Հ��|/�����Hv}��p��K��(u^@6�R�;�`��Б�Zw�ٜ��9��<�e���c��=�42����S������x ���������f}�W�Eyz�bp剛o��y*�`,&��s>�R�6�A3k��.��p_b��TqV��b"�o]�h\C���7�{�ev�0\7�E �ʉ��T�;�'Z렼���5ˢ��}rе(h�Y�垨��B37f\jA�sv<�*w�#��o�M+�K�n;�q�F�	{s^���F�[5p����w#��~Wro��E[h�U�$M�)�)�k���ƁQї�ӓ�|G�c��n��+�͸�	�5�y8�#�yz�]����wq����Vݹ��G
2�<�]H?m04���
�z�)r
R�UH�+�����g��q�O���}̟��̺�;.k�߲���R���NF���s�@���y�^�EG�A�Og� �R��M �����������12\ײ?g��MǿNx֗Y�����u�?��>z6�׉�^�e��:=u9GD��ql��G�}�^D�3�{~l���7�V�W�t����qԚ����L~��m���;�ǯ>�.�kMӐ<�M01:@��^~��^�O���Ygs|N�,���Vץ �_����}t�E�%+�0�ў�w�e���T<(��;n����]G�6M_��BS��l_��9�!��^�mH�<I�B���:�=ز2+ͽ�����~�Yp�'[U��2�c�9d'q�k"���]��ρ�]9�I��e���|(��h����ޗX۩']�ֶ�,@�B��]�,���a���i��fl5�U�M��Q���zGXf*���ٖ1=F�i���Mm��η|��,�.YX��ofr&�Ch�1���[�l}����Ww!z�pg=��7�
�RTna�:�^�n���p}׶m=A�Bs��\苝҅<ት��ӫ(A����99Y��P��x_MT:x$�����<EdP@�bdV\X_&�-�s�K{��c�r���79���6pȉա��lR4d	�M��rb3�U�\wL��Ԉ>1Q�
U)�;�F�	zU貖U�e������VTy��rYw��ur�J�@f��-���=֩ �yuƮG�-k�zo�+�Cs&[���?L���*7u&�^urMD��/�CKq�e��u�d��{O�c��v�z��H|�e]�9��2���C[�����O�V��|�$ofqI�D0�[c���;I��`��|b��l���uk��]%�.Ȉ^)�Fݺ�Y@����7J�y�e{�G���3[����bu�[X����i�Ƿ�OR�ͣ�Y���8:j�w���I���=�7��v��M̥"��ݬ���(����i�v#2�6���u2�rge/�	cMn��[�(��9u��M�i�t�=ҡ��y�����]G_n11�W*D+��P&(�Vpz�N*;�>֕L�H�Kp����)��Sq���K�fҵ�P���tD5�w���2���V҂��Zpx3��\�	�]�N�WQ����Fm%��FK��1k�kz�N��;�)����n�DҢ�m<��)�Y�\\���8v��V�z(CI��ۣx�3�-��R�ڕ�����cS#E��2k���_m>��=k'L�������0:;}�"y\nG��Ǫ�R˄9��K�5�NP�뺲"7����Dȷ�c����8k
P���v�֪�6<{W1�L�T�Oi�ml�֞Tm�=U,3�c�؋�������r]�q�B��+���#f�{-t2a�FM��k�,\cH����,ᣩf�\��n*�ѓ�z�oX �,��p<l�f��۽a�d�[Z����i�I�닫-.�l�m�"�X:|�����n�p�}��s���:c|Au��S�k�{D�;f��-������@��Km���mG*�3Ȍ���Li�W��Ң�cb�fԀ����b�����X�I�m�RS���g3n��=��Vm���+��i�ڳ�v�U%/�L�Z��;{��6�
êlT.]�q��r�X2�^�(7�Yg�M,���f�r^��9LL_6�c��Ґ�/рY�NV�%�v�޵{u/��E���:��V
�38N�Y�nK��u%��5��e�	�3)�����	�Ɇ�ˏ`�;rq.���6��R$����\���z�AMUSNu��¨�X�L�B��;�Dz%�bꛉ�D8sf���^{p(Ī�5:h��U�L:\���I�M��a秹�J������i�)*k0�g"������W2J֘�V�EEb���J��-�=��$Q+�"WH�r���C3�K+f¤�Q9\��8�4�9�	R�!�D�
BL�,4��*M,�*��\R�:�I�>Lp���^��J���;�vfIX�jfPU�C�.���L�0�JV�Q"�r���j9;q#'q<�P�H����L��U:̖9�mp�����bi�!Nl���Vj���Y�jbb�X|���TJ�3 �O<<�D�=�HO����H\��$M>w�+J2u�M�I\�̷q�������SL1B�)�>wuws��T̏��+�V�T�D���,��y�	R;JČGuӖ&UQfV*��TYuB��^{�AV�3�AAu����|����wj�d�N�K�5׶v(��X��i'A����	��dȒ϶� -�7&,�+��B�G:���Ģ�ֶ���!s�7�}S;�R�3�mՉ�����=��xd'S��i�[L<��8N�?\X[vд;"�+���p��3x��fO��[���.��G�ԅ_�ֆ�o�oB{A�i�Rz��ឃ>K��k�}�;��3�IF��@��H{��9��Zz|��cS\}�r&��1���9�D��R��?���x\Fݻ�|(p(�P�8��9_n@U޵�43x';Z��Ĵ�졳G�����R�mҙ�3� ��h�;E�P����d\���x�w��{>��5}�����l쇐�s3�����-Ⱦ�u(Y��6T��襖�8/q*����jK�ME�����p�9��έ`P��ٙ�骜_y�U@��p�Ʒ8z���{�P=畞[�|�%�Ƽ�������G�/���\vF���S�ю�H��fRS���<�Q%$��N7�zpW���D�j�Z�O��s��l���u�3��dg˙�:y�x }�Z����ǅ/iRe���3����z����΃����|��G<��
��( �m���.������� zM�&�k��*���AjNt���s;νxFx�]��si�[�T8�d���UaS*�1Oyil�|�qR���T���/e�6���Κ�䢫�������.��ܒ&)-�i�,
��Rq��fv[;�2��1~��(gꟳm���<��'�̬��W��Lu�p�/�9��3�K�o�w�~{������߬�K���g[������>�����O��XJs/�D�P�c���>�v8w׹�4�J����Nܮ3'w�0����1�^W�����u)J�Ľ�.��gug�W�Ϝ�9Vj���u:��]E�ȟ2�\?�!��1������������W�.ZJуݦt�"�H.��G��RU>Nr۫o�~<��Nt?ǫ�����Ҧߖ}3r��G`S��xd�g�(�)(�[S������"�t�z'��u��gz��jq�r��S���Bq��������|k�d@�Fa��-���^*�������ÿr��M��A;�nw~�˖�9/��ޤ8�o�F���d�;��$x�n�����1�s7�Gd�8y���0�\.�c���c�^���Hm��7�N�,)%������y�x���
�~��3Nǥ1#�\������lZ��vۡp�=�0Md�Ds8��ݏ5�� G�zc��:�W��U�ڍ�J�*�r��7��ԄC0O3��uk�0�Ut��5(p�Т앚r��aw�՗�D��Q�)׹����*圹�p�*)���I.xz�^1ձj����e�%�lӭ�,4�f����(<�r��9�{��y�I:���Y@��W>9#G�P]j�|{����K�{wB.;�ء�8��.�U#�j�پu[�>�W���Qt-WK��a�Kݷ�"��M_ٴ�\r���'��U������v����R�鐽��teT��`i��*;��,�*y��}>�Z��w�=��=��]���%��M�b�їJ����}��Y����H�z,$c��@������fV=��{ë��:����׷ӕĴo>}Z�@Z��M�<(��m)+���l���-�+�o�u��p�ɭ������]~�OnP�13q��cSj�wYZ1��JM��k�kEP��wB�]�,�^���N�I���ze� :g}u���9���za*�=(��h���P���X�ǖT��-������%+�3� �.�|��NC*��,�.�"���1��z|Λ}�e������ ���1�mK7g�<?T�$�3'Õ%t!V�?k�Aq36��Z�;&��y�>�܏u�z���Phd�i� i�TtM�:���	E��>��7J���W���v��f�y�0�E%p�ͼ�R�Mf����%����B��* �����L�oRg�ݫ���Fw:r1Q�N�5t���铦�������'kv8�+{H=��%P�˱��AU��'�!9e�	\4���B��J�
��}��}�↲�z!���}D>7��T���@�^� r��,�9��~�彍Qq�����
V��hyM��[.�F}�I��_7Ai���|��U#�6o-К�b��B�vb�p_�d����/�����J�z�1���|:� f)I���n7Uv�^4���!c�H�u#�����{�&-�w��>kW#o���1�z|��������	7�7�{wL��U/8q(�;f�T)������}^�qE���]Lz����'8y�p~��3��Ӱx�H]��l�3q�T?F\R���2�+�RG0�� �[s��ޥM]����{<����f][v�|G
2��H_m06''�U��ߺͰ�*2n1�,�����\�d=�^�Ǖ����w�32�^;.k͚�k�ʮ�S��Vo��A�=w��{��R>:�u��l�8\��M ��b�={q��Z������֯߯��o����٧O��q�G��3�YT�s�%R��XB����W�=2~��!�Eqב9�i�0��v����nX��H�t;
���a�Wbi�0�[��=XBy�F:=u��>�/��v[�z��XU������]B�۫�G�$-n"�������
�jH�Sb��㥳�ӓ2�{곒��7��UJ����2�@��n]�Y��s��S��rTJh�^��������U��φ}� ����GMX��e�a�V'hr�W���4�y��S�M5#ohOd?���Ȃ�ϼ2�ٴ��tdY�R�0���+�H�S�͍��q^�}�}/�n���tB�M϶/�ǞW���п�ڑ�sĞ5%x����ꒋ��7����Ի�26%𸅤���c~~��,N��D�ϲ�^�D��xz�E�s>p���K3��E����5O�,�:��5��o�!�;�>N����kn;�L=�W��œ+Vrhm
��
�h:��D����O�!�;&�w��;��'������Qۆ��{�.�������ю�%P@�F@��d �Z�p�ւ�;c��=ת�-�^��o�h߀��<�����C���qV̖P� p���u���aL7������S�%��N�V�n����[�t΀��,�����8� ꖊ�X�	���Y �O�1���B���w���-�.����y3>y���^���f|���r3����2l]{1+�`�CB�����c�pi�;���L`3�`��g���9�l�7����y��4����k5�q��hs��C
t��|]�Af[��򲥖kRpX���T���9�jK�U�t)t=s0�9�����W![���;
�j��[�^�Q�}��>U���r����q�j������uk�n�S��L�zFV7 ����N*�7|�mO��H��xt�w+N��mxVl�=����B~�F8�C��N$xǧ�d�Z3'/�n��J�	l_���6o��T2c��mhr}�ӝ'o�ͤ=y�x�n���4����β=~��[�^�NOS�Q�Z�Rg��6�O�{������q�s�� ���3W�3 �yw���Ժ��H�e��(�n}�<�vm<Vep�3��=1�p�=c&#p�}k_�U��\��Y�VANW�_K��ӟ7����7	��E�����+���e䦗�{|�~��*�����n6e�Q�@�I�0˳����ǽ����i��:0m,��e]]��[�����'	���3�\T�mEp�����O�r.�c��n��������q�}�[ى�HK62s!辒W�P,eJ�/��sM�	{����!�cssB&/E�e�c�|�[#��&�a�o�{>%���$��,	�R"L]�������MNB�j��5��� E�U��(ݯ3��z:�m�CjRu<��/+���$�^��k�9F�!�0/�j��'��u�]'^4�Ɗ-��a��0L���tUP�G���D��lq��CNmK�Y����1}�贍��#�e�Y�Vp��S(�Ό�=�
�a^�n����w"���*��HN�~�\{"I�9TA�p'��fL@�kr�n�����L��qx/}�)�{�<2���Cgg�[L���zJ�̗5���G������{�|���ut���x��F��޴j:�o���9���u�_ͻ�˪� I��S�T��f�^��ZE�T�А��N}����O����.�.��t�2R`<���>J*�lL�f^z�9��ZG��Y-Q*��5�Oŋ��]��t~��~h;�t"㻝����m�2B�Y��':Cp5�1��E�=�rz��>�>�/U����7�#��m�OO'�*Sܸ�6�hw\� ����j���̏\F�����ԏ��*;��,�*y�.Sf�7U|�W��V/��m��T�7���q�ܺ�c~77�Y�����z�#�̝�cn �j��>���C#4;�X���T�o>cΪ{9c��9�D,��!4��N�;wh�o�ث�x8�;pp�.�E�]cSۇ�g�@�T��+�ʎ����}1�D�??Hr�����X��>��#C7v��Rv>��Z�'�.X�q�x��K�h�OϷ[�e7HGpHþ��/�*F`oG��*'s��,qֆҾ�ݥ'`�[J�;�@rl���n�!0��^6���9��88�;v`z�R�Ji��;��Ai2��ह86��)�X���Izߏ��]{ǲz2�o�N.z�;B�~w�i����8JW�2��,]L�d2�L�����5;���ZJ�VjC�2ԑ�C��G�^�<���b�kjY���p0�r ʦ,�n�&��]���~���Z�iX_Lk�s�9�zi�X�D�\7}/�+��육��ĕPf�0�8��Z�w\�����ԝ����/Z��������>�c��ߵT���@�^� r��V��9�ك{��WvoQ:���<;��ϲU���l��1�l7Ai���;7¢���X)d�{���ґ�[^�Y�8�L��ޮ��`Rѿ�*C�׭����;��6>f󢩥.�vuv����R�m���D(����3��Y�,*��#n>I[Q�&�g�z��{���z�4=�Z�I���G
t)L�����F�[5k��_?#<�0}�WEZ��<��n���n�B���xπ�c7}��e��t��>�+�RcqM؏�my�;L�d�X;V	�F�^)kc��(3��<<������4��W�	%d���W)�E�C&b���=�K��̉T��m�V�y��mԜ]�P�Y�GP�D��u���;!�,�76���k\pᚚ��K�jQ!Z���7I�4��`}շ�4Y}��{�[����^s3.��3�����F܂��Zř��<����uz���&e3�!dj�!z���ח����32�_�칯cvgX����Q�\q�-yy���9��B��J�;pp�Wk�^*�/����dEu�do8>c!z��zk��[�p�j��Ka�r�;���?��Ǡ�:��@~��~߰�f�9Ty�&�܇9\u�H�؉ӭ,�h�V�����˦s�Մ�;�����Nb3 �6+&����+�M05vS
�)_��.����H���!C���,��������9p����Fz�ϦQ�J�m˩�5��/'B���P��}@R�M϶/�ǞW��/m���u�sďCX�k���H��~^��c��T�2+��c����2�c�9bw��+μ;%���p���mQ�o��B+ݯ�K����M`xg���1�>��7&k˺߆=��xg��8z�ێ��S�=�tc���:2yF��s��<k��ޣ>`)@�>nP��e���zP��Z�S�U�������}R|�杚Y��_�pg.����K��%�o"q�8{9�s�HmC�f��םb
�U�r�q?9��%8��|�`�/����ے*&(+2P����Oz]dx7+T8��2�:m� �������昦�W���]�0���u�l��.���㞄�q;p��x2K4��ʢ���|J�K@���ZW�yJ��:��{]z;'f�5/iu���y�;��d��؆d�_|���	��W���|}��Mzׅ��
���czׅ�pUn8Or�M�>���t΀܌��m�L��pTuSK�'�v�D��M��o/�|K;OL;����1��G����b��+��to�� }�> o��z���Pz�.~�Z�2��bG�md���*M��a{�������}wB�X/�ٙ���L��܉���+.Q�w���˧���=����C�9��i�qOk®3i��6c��>�\��ǧ��/x�Y�<���#��}��H�4v8��_�j�mhw�O��t��ͤ=y�x� ��X��+�=7Y�u&)���~������J�C�	��=JB�Tǯ�0n�?n�Բ���ϗ�v]2�H������ϴdy���x��ΤW���ע���pT���Ia>�`z����z(�%����VE�+ԼF}.�N7���п�κ��d���D�Oz�&��<���l�^�yu����7����n�,GVW^�Z4mr2�;T,Wu#�ﯚmL.ԫ���E�{��;�z��;��T�j�1��J�u�u�H�@�w0qn��]�ch@OJr�w��ΖM���#����Y��I_$%4IN_ga� 9��Gq<x���KS����E�{y�2f�7ݭ�(^��z�dt��+D]�g+yy����g�7��Êfa��X�Ut	[sC��X
�Ar�U�`M��̼�!��_4�����qN�A�{6���+�ϐ��ӵK��vX�q�5<�K�x7$�h��YWJ�%���fhe]��E�+������q�;�-9�Ȃ�j�&^P'r�-���M�81̄��J��.�Ϻ<�����B�K`����̕�����฽�� �7>d����`5/>�jr�@\�}z~X~��PN��,�K@4�絽�`r]�餆��se��g^0��iQ���W%�8V^�X�6b{&�VbĔ�r��Ӯ�Z)m���N¡�ܣw��(_o�S�3���)��[in����rͩJ�gu��+9T.�E���x3�w�r8�$�aɺ6-A��o_|or��z��_��]A�g���.�YT�پǴ\���D��6ڭr��_��imm�sD	ਗ਼��K���VM��zR��s��U�a�xr��u�x�Z>�9��4�.4dZ�j�lP�u�l�r^��{���WՄ�MmiffJ߹uV�
MK�v�nkg|�����Y�EWT�0��7�Uw�׀r�Z�9���s~.�8T4Tř��������N	��1v[e6,�ks�ne���Cf�-��5�gG-?�n����:1����QR���¢ �bI��gd��K��!t�ڑ���sJ�M�����Ŷ�e�Vݛ*���n����	Ed�$ugT{����3�6��ϙ���c�ΩC�	;��t�˻ӧb��Ջ&P�Q6/��k���i�8�kbb��
nS퀠���&��J\v�Pċ�x)G»���H��JR}�ܗLqn]�Ѫ��# <�\���4§F]fϤ�!�a�V6���SͧdG�9��K�VV�AND�*�r��\����I�t��e����`�b)�{j�I:��t�p�K�`f�}XEڤ��\��w?��w~�u������0kg6�0�-G���A�,6T����_ز���?M��]���R�Vh���֑${w��@ĺ��֞V��ѽ[F�����M���	�S2�� �+dMN	8��"vfc�ܞD^���M�4�bY�ݭλ��5t���S�W[*덉w�w��Aӗk ȶ�N�S��h�c�抰/z���3��1�ms��|ڨ!�V�D��,�2��冕��L7�eA�����[�7bK֢�w�֞$GٳF�(W���(Q~�( U�W@�[E��f��E䠊��W0��wr
���G��KU��Dh֩�e��T�*I(�<�"��s2��*���� j�S��볢.����u3ZU&�#ݹZ�r�T���9V��\�	�ds�4(�C�p�"�L�Q-J��(���UIȢ���ez����*JE����4��1V�)���YQ����Q��:RY
"P�P�I��N�E%A�I=�t�\G3�dQ�\�EU�A&fZ�JQey��9�Wwr����,�L3#14��ʴ�CNE�E�Ue�Ҩ���,�ˑZYUQR�I!S���X�2s�Q��P��M����C"D�0�GG'*���{��Ir�5�)��­b�F(��EZ��F�D
z��B碝e��8A�Xf�A�U��Rg��*�J�r8H��:�(��
���p2���ب9�^ #Pw+��΅��rfI�a�짤N�ב�ik���fs8���[Np������2*C�rSɧ7zB�v򿵏�L�_���q/Eªq;q+���W0˳�k�a&��Ӝ�H���Q���緧KѠg��^�%���3��S>S�w��Qc�'̹�1�cu�o��`���z�����,�%z;<}Z�����z��$"��R���|��sBzz�8/F��nz����ܰg5��IGSU}]o�{ d�k�x��`X)(�[7^&�6{'���:�]�C��,�y5.�z��_QHCm��H_;w'(0~d@�8��W�k�4y�)����\o��!��"�1�.=��Oogc������W��T���]�nd��� 57��K��v"��{9Nҍ|WV`�/6j;F��=}���<��H���f��N0T�{�(�ҟ��ҩaxK�Dgh2,�엛��+]l��ߩz�ݥ����c�L�[���Li�-^.R�v�O�Dj��"�%�Dǖ�`�����.���C��j]�=���0l��]��b+���Dޒ��O#�5�1��E�=
���s�O��DK[z2)��]�	QJ��μ7��z�%�dM�1ݵ�h�)��^���8�*D�'s*pC{2�F-'�ib	|85�Y�+����	/:��ʻM32zn�.V�<��a���E	��;��ޱ�6�o�t����]ΰ���AldH�@k�$#<�H9�N��{/�wI�xٞ��n���Ƽ����5 ���ʎ���B:�,��Y�kU�0����J�����c>n����y�u��o���^+2�r�+i��+�-g>ܵ����8��x\�o�b��s�W��Ϙ󪁞�X������SheȮ�<}��Щj�R�O��ʭ7�~%��Y�Q���e�Ư�W���K���F�p��Ǫ�3���F��ڨ �*�ᚯN٦B�=S�72�W]��K��|b��d~���z+�˂p{n=��]��'ȝ�X��2�@<X�|�S�ʿ��.������x�>]E��5�z��~�x���!�֣d�=��x��f�DT��L�C�,�n��s�w�eE~����~������3��D{�޶=�%� �d�X�J�3�=!�Ŕ-����Y�݁\��8L�H\A���}��qx ��~"{���R��wn^D���D��m��2}ں:��nxy>�:�ځ_)���7=� �ۊ�e������6o�;�\�+�޺�^E�C)g���Q�;��,TΈ�����/QĪJ'�K�*�Z��&��d�l⥫�t"����#�� �^�(E�Z�ʊp��قq����܏{bTi���6�ˣpV,b��H��:z�@�C[FI"�kz��y��֥l��Y�!Y�������Z�G����2
= q�������}KF��9ϩ�ӽ~fwi�����Z�*
���O�����K*Il	 �^SB��x�|�=j�g��7uV~�h஥���R�G���T��Q'�;�q)�1�B{`x��dT���KY���k����ӹ[f��N<��vn;��E�ۯ���n4
��2�W����C�=s��]�e��������:�y������+����ns��g32��P{�
2��ԃL�7؜�����˼�Ii�����s��][��ᐽ]�q�����w~��f]�v\ײ�+��M!����{������ʮ{]#���s�*�����\A�@!x�X����eu�do8>c�>���AL�OGY�'}���n��ƴ���;:O�&���S�������,��#5½�������G+7�=�޲��갖w����	��W*;M=7(�g�e�6
�f+�b=���)�ۧ`guh#��s�!C����ϼU��Q>0���k��L��D6��Ec�A^���u�սڥ�q1kA`�{�+���ʇ	�0D�
�9=55�3�9��yTy�P�nm=�-�T$����N:Шb�'�1��S�����켣�;1��j��e�+V��	�q�XZ.N���oK�.��Of��Gtu��pH����D����ڛHf_딼n�Dg�]t��}=>u��o��\]x���rq+Q�QL�܎�i�����YKp����;������yӰ�n8N��A|\�"%��:�7t9Q�mWb��%`��'8�$�t�=$�1�>��E�V&��������<�7(�.*��B���N�Q^��DZ���p �X�(�7(+�~>�O
�z�hhr�baہ��^lz�����#]7�1X�S0��ʀ-� zd �_�{��&�˾���ns �G0���0yRv�/[�(������x_����C���	��WQ�1ɾ�^�Ոv�xt���Y����ʕ7���Xu�>b��-�}2���_uS�� v�����o����Ng��_�O��!x#k����p0�{mп�gd<���<�L��w~c>��~"�kÌ�>�K��	�CՒk|T�4�D\o��/����}wB�:��B�f|�x=厽Vo��V�� �o�#������\NIZpK����=��w��ވ��`���eC�����y�\h�1J��jݢ��L���F�޵3����6Q�3+��tDҜ&�C���zWv*��}l�ބ�����NX��^��@˛#D�|�G$=� ���߭\���-��)tX��[��D�I����EZ�|Lǜ�s� ���t6��4͛��U�j�Z��N����;q���c페�hQ�H�žדw����������BtX�L�3����+�C�4�����+=^�J�Ѵ��ëG��}~�����ӑ\]����(�n}�#�ԅ�n��'tvr��� :��~`�V�ת�2��J=39��O�Y�'+�f��#��N�k���'��n�J, �Eߒ��vg��n��8���V`��N�!Ľ
���.���y�W������+���V>�ҽ�[uݽA��/�2j�|?U_"O:K��T����ʯ��;�p��t�l?� 9�������Y�R��!�;)Tw{���o�ei�n/���e�?�X�����sM�	��~��&Ӊ]���۫�@�OK�\�~!�7��S��� 4�
隑�-�t�ǋ{���Ngdgq�u\pwq�M�Zݩ}��{����[5��f�I�`@�a���_M��8?mr����7%g���J����7���o��ybe=	����3S�������Z:L{���+>��*m�W{�5��ޱU�օ�[4�`?R9]����SE��r��*�N���	6r6u���O�C���w-�W�x^,���Eԑ�  ����VJ��TOT�Ӟ�W�y�n��=n����ӛl��]KX�
�������E�������G�����qy��4n5�c����T��^*E�ۿL߭���g]�yc��#�ƽ�$�Q�%)Hϥ��l�x)Q��j��m���0�?;�@#�z.|�hڜԕ��͑�d�' �w�<H��O��a�
�TK��>+-���Y�ew�}W�,�;���#�*�uء|����G
<�lL��uA�SO�rQ�h�[U�;��/{̪j�)x��/y���Fs3�V�9��אP��jA����9Q޹��uD������e~Z,��M!S�	5���ߕ���w�b�e��F]*�7�sq��Y�`(�m�ӓ��w �7��y,>��8��/E� ��s�����Z#x����0v[�7��7go#>�7��n6�exHd�q�RWO��eR�	��>Ǧ9�ubg#�)������<V뱱^�����\'X�z{ �����ӹ>����򛍙`+�.�O���8�:�*$�K��N^�-xl��w�d��7|�\o�]#�p��b��,]L��!�ʝ��Y��㗙��C�,�����K�7*�)_37@�ӯiW,���OR*�k���k��|p}:t�uN6H`<�t�Wrw4��.Т0��%�:u���G�u��u����-��5��ґ�Y�����Er#szmep��t�[c�w�C��c7��ci�����GnUp�X���Q�H��;c� nԽ�#U��=�_f����e<�WB��������=��[㑞���o�� ��b���ߟ�eD��p�\#pE>j��}��qx=����|�D��[U9�wn\z�q0+�O�F1��ϵ0�Md���C����x	��@���ȅ�a��S����H�uRc|7A=�Ļ�m����n��-�w�����u��"t���������E�OS�H��c���6P�S�1��Ӡށ�^@^�q^d����T�Չ �^SBY��
|���E�>�#+{zUJ��"���<3�S�d:���(����������b��z��y�
-c���s�͜ӡK�T[g��#��R瞓S��,�3>���ƁOї�WNO\!�W}7�[ŕ�������Ԭ`��z'ʷL��F+��{�[�����\g32��n�σ��FUǜ+�� ��,�4�^c��Ίͧ@'#�Д.uA␿�h?����:���7�9�@zM�z��y��bAxNyӟ�Kj/�?h�0z�uu�~�֝�l=~�u�l��qμ��Y�.�Pw�\�����7 �Ȱ����J�#0
�ۓ�>��l�
�0�������w\��L1��BRV�s�`#z�:��{�/��N�*��)�.w0��'TԌ��w@��.�H90�޿��|K�g��a�����۩zN���^9Ԫ�5�"�M�����ٿ�'}�5P�Ω	����O��<�㳷3�*:�NQ�qJ���P�؈*��n���]"-t)���v������h�O���Tv�������:5k����v��|eM�^W���}hr���B�g��,�����O�:6,`�*;���^�U���y���Ү�U�,�,K yti�,�
[+�}�~�<�ԇ�(�{h[[R:F'�VG�����߳��B�"���)迈q;�uWOBt�r���9�dA|\�z�<	�'�����#�7H�X����؉�50�*e��>��[ubn#[�q�)>/�5�=b9N�<0��G<��\=9��ˀ-�,	��@��A]K�_z�[%���"������bZ���v��������z�ه�$���`��[ T���w�:��5�5]�;����8�m����������z��6w�_�;��~���0K:���D	�}3x=��yan�ۂc=�-+�ӄ�c���Ө�'qʺ��.łoۀ�d�As�  &�X= �u�����.V��&�Q�`���l.J����_8�A�>D��W��=}z��7w �]q>ǹ�TJ�7��d�&�9�N��6��iQ��i�0<fw����1�צ\.ܩS}ϯ��Z�)K�m�L�8��S�׃��]�J����lx�⵾�^�$L�FG��f�?٘΄����6��y3>y��U�����f����W�6�tz ̴n
��&�s���=�j��Gi,_�լ
��T���i������eo0L��2����*F�;~����E�Ok®3i񿽷�T�]+��,�&ǎ$�v�`��q���.1Ӊ�n̫���b�P2a��Z�i��S�'}�Z5��]�wϫ����ۼ�9̿dd.f|�1LW��&{�+(g�R�T�!
+Ы�Ly�q'�+��ӎ�89^����Ϣ-vۜ�.Ԍ���:���FG����x��Ϻ�	k����_�k�3پ�g��>=�u�Zn(��� bj��^��2]F.���\/u���7>^���W��X/�F�h�(�UE�B�Pc��C]ʓ3��)���h������� ����~����� �R¨<�ϔ�Ӑ��F����^�N O���*��:=���ж����9�¡z���	X)��OȌ(�v��/-�]���'{���0�ks�s��h�/*Ǳ��[JO4v*�!��<���j�0uG;��(���]ӣ{��Qd��(���\��P��͓;���qЋ�d����"��{�^wA�"�a�]��z�2�����5υ�k�y�X��q>��y�8�i�����l�ұ��=p�\?d)��G�$�L�%Q��)
c=������o=�݆Y06��㚑��O��/���!�V�`�;w"r����v-
P�{dU�$��=.=ǼfO�+�3�v���n*�{�<2������:�^�w}&��w��qFӑ�����>��Ј)�G>�p7 �>̄j7��z��p�T�*�/gnzo]9S�~���y��w�w���V3\I(lB�?��$�B��81��~:ј�m_�����\�d�N�o�&��;%Nq/�ցO՞$;>���a�
�{Ɔ�W�i�]O����P�(����w��n���wt#_2(s��0����2~ۮ��";�i��]���2Y D��	���ˆ��^��î9]��Ȅ�w"������̏\k�(\y�5 ��~�ʎ������0e��:���0��<��H\A��/[�M�^_NDw�b�e�����^���k�=F�UW�`��3��N�iRk_�Ч:&��fnޡ���ݖOwm��1�j����PV)Q�8�M�f�6V�7�^��\�aL9�n��v���^�,h���7�:�?7�%5�۹���ڦ���`��1h�O0�tC��[{��]oY��++�5���ڶ�灭�(�hs�K%uF�0���I��z7�>3�mt��H��{0(u6H1_T\@�ϴ��Ȯ�¶�v���}O���eڕ��BV1k����3��.����\D}������2��WK�R�M����M
���S�x��.N@l��dCn��$	%ZH�xF0
�l\���.U{)M��̧ԋx��v��\x�v�g��b��ot|˨N��a�]w�J\��,9�q��]���:m;�]�Q�Iv,=N�995�J��ׁq�8�{�k��X��pY��(�N���v:��A��l���K!*6(�6<G^Ͳ�$Y�����O,�.��a�{8mǤ�\�n.��z�Z�m��T{V��Y�mP�pU�(�9����b���k��}{X�Ȥ����sz+�o��&dFhcgݻX�7�+l��|mB���<{���:�=}���4�I�E��܇�P�0���R#��˹�ă�r.m6�5�;��m�KJ�fQ��r|c��6]խ�G�jy'�i�nP}�*���wv��5�bw�*�cl]����4~�%� �'j]���K�u�k`�3H�y�*���{��`�AY�0
!��i�Հ�|��=C����ε]b�S�SQ\$���7�>����n�"�a�����	r�ӐT����W=
�>ujtIVrsͲ2r�EN�MP7��+r�g+��2�w]�]�L \��D�ا�=����s��=�d��֦�y��ύi.��W|���(��#�Atuk�o�%�ހ[�6�$o+�fʾ�sx\,�j;�R��Ӄ��i:������1[{N���C[�m^>�1�<[Ѭ���L��'��s�%�>�ش�/ ȁS3��z��T�(��B��]z7��KN�p�ێ�,��v(ܹ|���K8�Lʶ��5j��K}�	���ݐ�r��֣�%�Ψ$�sAT�b���7��ek;"�F�+�8u�B������p����xeo]:�=J���8(^��uywm�ͱCv�=�����bSVf�ڗ.�Ff�N��|u���ݱb��V$��;�����PPn�\2�G���-)`#�|_X��C�1֒�h�Ά33Y�+�Dan�M�]�V*�"(L����M�~t1Vꥸ�+Ĩj��k�Wtz	��p����I"�,-����8�,�f��sgv���j�l�Wp�D��ZfՉd<�V��ĠF�|d\����$�7� *��z���_]l.�3O1,7�tu;mwO�aV5�B�ф�ܓh����<�YI�ނ�6��=8f�����[|HS�b`P��W����9�`hTh��Μ�R�Q�rYUTrRTqВ�4M���ε@�����b#��D+C��2�r�EA�9%�^#����E9%˕F-
���-2��V�-RG;""Qc�Z����ʃ��9b��Q$�8h$fj;�p4�W ���A�D�+��-K$'W	"*�Q�Ά�աz�t��(��̎���u�\/�����\�g(CZ$뒻���'"�!9��\�9^�]nG�HH�ܻ�j�����i�0��Vf�,�K����
2,0�8M3E,S��S*-.)9�]ZE���l��MR�QUK2,,��Wu<0�i��QE
I�adAfB���f���6�a�j'.s2�B19.E@��N�XZ�(IIi)�P�j��������(�
V��U�m(�����3(�K.�Y�jh��GD�ĉ�營��k�:�2��ج���E=b�$�n���z��b�D�%z�n��B�]7t�Z�9�l���9�/ p�����Y� _�XW߂YSk;?A�9 ������^ۑ�O ��s�3̘	xe:�]�Q1�zr�/cu��<��
#x�8p;<\�w�eW��J6v\�UQ旈	߾=ɓWg�R��O\L��9��o�O������（Am����v��Q�,�)�`$슝hNA���;�J�.'��Z6G�]�	6��"�>��9��% X��O���y+W��[�1���45�
3�b܉���ұ���u����������£�P��ZxU�=���1�Cg�=S9�uR��D[��o��{��8��Q�z���/i�(p�GJq>�P&Mb\ܚܿc�1P�k��\A�_ƫgXȾ�qW�m�>���Ox[ZjV�(��٣�r`�Ir��(�"���'��ޚ��'��@��������~W��$Y9��w��]�1y�~�G�ͪ�<�wR�6��7�Af�PGH��u��~(_-��:�91d6�o�s��!5��S�����yp۸�_���3}T8m=�驞�he9�����L��ǷFo��������� �;��<�s]b�ͫ�������>�.�F�<���]�-�y@������M�;�х�eȬϛ�*���"f|��(r��U`N'�x�9�9Ct�#��
`�\�*��l�\˺J��zb��@$�n%����*��OϮ�\k�sӎ��cR`vCI����)�;T'��k�#M7�l��U��������G�d{ʍ�u!����ʪG6���<g�w��n4�.$힡�4�:�g�m�^���V$�R�q^�HT�>�W���|n��32�۷3��8Q�Y��O6^���tnv����6?U3 U}q�A�g�B�#�~�]�g�.;#���d.fg�r����`�+���9��"|��c]NUuǩ��`e9�AOx�r�r�;�T��^��X�ՙ�bJ~��d ���'Q�F���{?~�����k3����3�(ӡ��9GEҟ����-T� �������{*��ϗ�q��y���cW͛���h�O���J��馋�z�\8}W���=���W��}J@׳Nej��q��9
�c������vn�Yёc �e�{��ykS�O��/��f:�(�]L���e��3'Uk�k�g��{.w+���[K�`�'�t�ǋ҇)S��q�] �P����OE��;��q==�>e���r�N�%��h��+-��0�a�%{i'iRwhv��S���Q��حW7W��{�(ED�����)��2�o�X�d�*�ě��1X��jk+��1�ŝr8C��tY{�����u���{������՗O��#�r�eY�Ov���j�GNDʌ\�]6��{{�g1]��r��p��w�'��'�e�0<�����O�3M�	�[�q�Ij�.=2<2����8�)�BrY窡������P��ʾ2���@>���5�yS��G����h{���$�;}*s_�����pӸ�n��GdNIf�9Q�=0d�D���sqܪ��>�=����خ��󽝜e���C��s���pӸ��v��
6f'�;�qj�]��+���v��L��d::��>��֮F��3��D�<gG����˫w�P��2>ץ����n!K%�L�$����D��Q���o�����P�{m�m��}��Ϛ��eE1ƺ�T�����j��78�P�2Ѹ*pTK�RhsB�Wx\n�p�9����2I�K���H��|�>MP�&Fw�aQ�h�U��Y.����<��x�x'���o���W\ߍq�;��D&��N$z۳+Χ�#�J*z�44L�aJ��T���e=�Ox,'̚J\���뼞����dd.f|���n'~�����CނV�`�!�e)����#Niw����i
�Q��E�����-���r� �ޅt����7�:d����x0��NSE�Ee���5�q�x�m�ԃW(:P�G-Ѿg�30fU��R��	��[���Y�Y�*	�[�)\lԛ*�R��:Ҍ橊8[_��<����=�̟�=�9\]��_�r�n}��V��x���
���1���a+8��(����Tz�+*���_�W��`
�ՐW�X��1���t��9��2���xo�[���z��<����"� �WT��u�n"���n#f}X�@TBN����2�⡫s��g�ȗ�z)����{���󮢆Z�J��aA<��1�NBsk���Z/]f�Z��ǋ�j�@�H��h�������~�V��W�$y
�$"�Ԫ@W���7�ݠw��Q>}rw�f���n}/e�N5C�p�\?d)��@�,�ĕ�X��մ�7Һʰ��$x���/i,bE�~�{^eo�m�Gf��Y��9A���櫫���evx@�2�;� Ex��F��z��*ᗹ��)�Mץ��R�uu!Wݖ��@��4�f��_��t�S� ��!���8���j7���o���L�x���qHeF����}� ���~`�{��)��s$�P�KR8��/ԅ]K�r"}\��.�aW8���I�A��q,�x�E I����W}��� ��uN��a[��u)HԮ4�g
�a��e�@Ha�Pʆv�r�&�޻���*~�|
rvi����|��IͶ�Fh��pV�J��Fbݓ�ʥ.��M ��7����\Mϓm���Ү��M�A�=�dq�ԫ����l�5+���Ω0}����3�	��tmTv�D��5���Z��ಇ�]y�c�쭳e�<����=����P�t�|��@�r�����\@�a�r��_��y![�k-R�俋� o�Gg���s�F��u=U�ә�אP��jA���ۮ����puT�mJ�C=��y�wu��"�����n>򼾜����3,U�7.�Y�~7;��}��[Wy[.HǺ��.7�7�Х�� ��#va�ey�- �齃�����Z"7��1F}6�c����Le��~Jˑ�D�{�<�p�[JB
�v	aOa�|.���*蓩����<nL��|꼗v���ׄˍ<W�=��~И�5��r����&�ӷ�
l�K�uo+�W�⫻|7kԬ�����b<��B���d��C��1o�]#�p���@���Լ! "��s<������q�)Uƙ��iv����_{���W�,���b�ږhx�U�4����ľ����R*nJ�uR�y�+�o��d{���Ͻ�G�۾��\��.��=��z�}k�k׆�v�b�ȥ�eQ�H�G��cj����ݮ\�q�-���p�^P��,G����K)5h#aEV��uw��	Npْ��:�)WlT�o_!��:���mp�Z��ʅr� �Y.���͵�ǔl�$Q�͆���qkQ�\���[�c�M�!�׾?T ��i�	L{"��n*e���M�w�9�'�{#�D>(��oPSb��{#|�T�����X�r �5%�!��P=-��,���\U����sӛ�@8Yx�z�Oa�)�|�'J�{둷�f�̂ʀ8�@�끰_��-0�λ�>s�绞�����S����K��07	�{����9��*�� +�h]t'Z==�w�^������Z�p�m�N:{a�uI��Q<�*#�:6�OmA�)P����g�/�C��pG�Q��.���R���u7�ŀ���n4躁���{;4�ߵ��&���C�EKB�{���F�1\w���~urq�@���޿��R�46:��i���� �o60ԇ���d��Rr�>���������w���ELȇs6�5ߤ_>��s�Byz�wн#&]��h��+:�Y^q/I�r3�\��2�7��m-���Q�IN���B1��2%�{>�~/�_��X�!���ZO�̴U�~���z��^�ď�_�N&��4�C������9����B�i�٪��j�\볜#c4'M�����l�}��B�>�s�0-������;�R�ɸT{�`�����f\���Z��z��װ\;Ûv6��[D���c��(���s�.!��9�-�V�,> �|}2m=����"z��=�6nws���/��Y����J�Gf��>����|�K�5�X�Z%����\D�?g�����y�z��9�u!{��H�B���37��_w�O%������#g��pz�{me��tD-��>��1�Ez��]/��>Zf��^w�xo�!4�ZHԻ�������:ȧ����k����/�{�����\^n��V�Ԣ&B���{�p�P�'�`\*�qS-�I��i��9�0�T�?x���[���5����0��൭��g�L8���t	�Te�!J��r� M�0�v�����`q�ޗ&���S��w��h!��\N�����$�J�� z�z]�CʮJƔ�\u��� �+�ς�޴�S���K���;�.w�p�����C�3�ڏa����pT�7u�}�8IͧF���/r�n�Z�/������>�)K�Jf�c��[��=�گ!6��Tc�=Bj��"��mz㙾l�jj�%{ޤ���x�/Y�VX�xg(x�s���� !��g���+�,�!�3��%b䮹'Y?�:�C��<tu��*;��{�kw!���'��r]
VEM�s�_��.��ӟ,�a�f�����=h�:I���o��o^�Δ%�L��38��
��`~�k@��e��9�.ϑ�ȗբ����.�����y�����b���[��#$�>����3>x�P��!g�ac\@����JӢ�ӓ�2@^�{�؛(�- �l�o;���B��t�G�58���b��`i��X���)��v��M�R�v�xq��^x���Gq~�ȅ�ϝbtX�Ȅ��s���G��@q[#��F�O�K��P��+۝�ck<U�z�}����>�.Ԍ����k7>��d����=��'���z�j�H�g�� �����0��ʭ7_�Wi�*15d\�R��Z��f���:a�+��N%�7��>���:�+"�	Co闆��B��U#Qp<�������=�c=��ˌն����^v�{F�/n=��Λ���x>$����0����T�Gy]�<D?Y[�o�x����cQYo�k��.E�x�9�u�m>0֎+GN���	0%� �=����j���嘷q���՗���������]9��C�o����d��}�%|:3�;S����5A�O�����K%��y��/P�}���6B��{�o������4����8^f^��q���rx8d*y�}Z�@�p�T-G��<*�t�[r��޹�ɖ�9L�8�7`Y�>�����@���c���>�ͮ��`(�W��ː��L{@�=��9>f뉁�w��w;S���T=!j�k��n��z�{hN��*���r����@���@Q�^*������ybv��lG�Hq>�3FHI{Բ����]'}"���
�J�D ��<d�\�/���h�kF����KvnQ3*����k�j�>�))��o��_q��d�_J=$L�Ru/���/Ƨ׋��fb�t^�X��}B����T�#�S&9�`OXt�Gm���5��4D�ݞ���;���Ӊ��>Xi*��k5.�����Ec�W>�#�\���s��K��1s4�}�Qk��u���m�ȧ/M_ٴ�_ܮ�1�'뺛��g���s#��
��#R*=0>ظUg�߳:+6� ��ꆮ&��x�,���B���o���{�����e��f��N�v�tG	p��]瘀�}3�Ϙ�yU8��0NKЂF:������/={nr+�h�pa/X�|*l^?���d�q�Lq�gO;�#m)+�`�>�ⲫ���Q\��8����y躼�R�*�¸�<�)�����
�%��ά8Wˬ��q�7�`�K:^WgBc���	N^Dk2�8m*6�g�n�Ňu�w:��p�w���=�.����1e�Ӏ�v�P2�����*Іn֐���L�m�[!t�y&���X5~���>�.�c�m\n�k�hL^��9PA\}2�W�g���Q�ң�PY虍����.�+Ӯki�uW�}h;�?n����;"ۏ{!�����t�7}�ql�V�+���*Ib�{ev���#�_�f�Y��lq���cr#ޯx����E֣�Գx��*�[yW���M��� 1��@�g��5OE�M9�Ⱦ�1�)�����g��K��}/��oq�1˚�8?nQ��(�"}�=$�<I�|f	��P�"��Q.P^4�TOKw�9�#��~�Ħk^a�񡊬�֗*���q�B��L���߇�%Ӑ)�,n`G�e(YV9��*���- &�r��- �j���-t֙��;7��uT�iAUDL���7\��PΘ�����,�2.�T��ۡ�V��i��qw�#!���	�y6�+���7T8�B{lH^��Q�g�۽�m��ԏ_O�)��g��
Xz�H�m_�������(�����9��1�����~
���6�]��U�!G�!Q�«��R�t'TED$����e��
� �1��xl��� l�����ck1��P�1�����m����l�����co�c`�6�����l���6cmc`�6߀l����`�6��1��0�1�����m��6cm���1���l����(+$�k t�����0
 ��d��H����bm� �F�U����dԄ*����KmYUkoN��ҪR%E�KZU�*���jd͕Q�Y+f�`5X�C31-P�٫/�"%GV�iiZ֭�v��Ʋ�m�U��Ŗ����S6˷nݕ��il��Z�[����JmJ��mb����״٬�jՍl���2جR���+1l��M�hj�d��f�Z+&��jk��)�fZi�U��KK�V��m�)F�5�����m�eo�;f�m��d�   -v�Pڻ�#u�
(�F
 �[���#LR�@�� ˻3�sT�� 
�]ڢ%�wsB��;U��l�Fڔ��҃m��  -xzhUa��sT
:�t
�Q���;��F�(J-\�F�(�(���hѣF�c^�QGF�4h�7�xt�4QF����4�(�;����2ɋU�U�ڬG�u�  ��A@���D���[ 4�t�h���� M�]�tur��TM�b٠қ:p+kh#�T�uE����Z��2�[��H�,ǀ x��D�l�֨i���Pҩ�v�ݻ���5T��m\
UV��4�h��9��J�t��J�t� w6����[6m,�EUb��� �oT�`���C��Uvӳ���P�Sn�í�*��9��j�u�Ti۔=J���uv�E]�m�C����taֵ@�u��mκr�QCZ��d���ku˾   �y�U�Z����B�Wu��t����U��Zv�J�n7 *�V�:���[��T���V�v��eE-��9�;amE���v���m+��D׻uU,l�E�¬�-�   7s�M]f�I�;c:�n����V�f�� 饫�� Хr�v�h�	׭ڭ�6i[�';mm�����t��/Y��\;a�VT��Se�l�2J�m�%�b�_   >��_l�֨C��lh(�s�t̦���r)�Cv�����[���]-�5M�)�#���5���S���l1��+m�P��դw�իf��6�MS[�'|   {����1�kkF�Kj��M4X���UN�5�uì���H5���w)6��gV�CYevꑋR]�d[%�t�:D;�LFTٶ}���VPk�7�   �x-{���N�ꦅV.�ۊUP�t7V�56Sf�avSZѻ�#8�hvu�ݷ#Cl�Ҵ֕K�]��V��s��m�UG��T��̪R�  S����  ��S�aOU*S@�O��P   �?j�b`  !ILU5(a)���ƽ>�W���5vz�¦O	�qm��D��x~����W�߼������* ���aWB��aW��* ��QeQE;߼���_�:����?w�������c�G��3��12�,6���f԰5K��ޛ�
�I�p�"-�C7S��!���a�ou0U�IH�d����q3��2�Q�V�����=�[�H5Jne-��{jj!t�;�k"��g-m#�Y6K��_n����"�R��Qʷ�m��{�"���n�J���!���ӽ"�Ԏ����@���~��dΦ+oZ��<��eJU?�gG�V1Nc�[@�0�A���{V�:�3)V��F(��0�rZ�wÇڬY��e�:��#t2��*Sj��㩹�CƳ|�cC..݇�D�؀�>kǑw��[~������e	sKۗ�a��K�=�r���t��F����K
�����G�sm�������R�׬���em+�k�^�h��ʊSM7.8u�M`��춉	��kw21��jЎjYj-��rȇ26<#Xv�U����&�ґ��n�=�s8�/�`�V���1�`��"�֚Ɨ�
�<�M���̦�)Y�b�CE��zU���ۭ�i�Ɉ��ؽ��]��	T���x�H�A�Ln�+KTq����D���(��VV�V^4)]�0�XAR�J�+Z�[HS�w��8��,m���JQf���Js~Y�PP��^j��4�h
�*в��G
�B�;��)�[����U��ǅ�Q��3f�1@���Q�3RZ����wlЉ��F=�>C��a����*��9z��%t��h`s� ���[����of�p蕶)j�V,b���):�7ZB�bk�yQ��k�X����A��/4 M�t���P:ER'ff�af�J�R�u�%l*�MQ<�b+NM�}��[j��8{G�S�JLd8�4V=r�^ѳ��V�M��Hn��&� b���W�Cj��á���dL�ıwz��� �w��vw[�����n	������
���!Kr&�u��^���c���G���M�^��Umf���e+m6c�!&/q�"�a+^6q�`��_F%Z�u`��5�+�D�$2JB:��-5+(�q��)�h/ �i�4qR������c��Ԣ��������v��W�GU�K*��ʒ�f)W3"deM�A�B���/6�f�'a���fm��㗚Z_	����G#h�Xج,��X���F�խ�6�A{$oe�Mb���ʅ-�b
����H�b�l��9�B27�+�n�B�$�ì�b�-Mܴ)�a9z���Ҙ����v��zQz����W��-1"7svA�a���@�U��Q�Eu�Y�:����̱�Ձ���fJ:3Q�f՛ԅ�GPKF�j���-�QS�	��L��� \ƴȴ� r�X9��m�L�P
D�Y�X��K�U��+�2,�yL:g�R��5�%��b(���R�r+o*��Ѳ�Σ�%5f|N���e��L�O���L�!��i�Ve-�tf��.�%���QƱ����_E(�F��ne]f�2�PcV��q�5�d��Z�dh���'�k�j��� Ԓ3�"5Z�&��ʓ3h��ݤXG:�������ʂ*mj�Ɇ���Q�r4��)@5MJT�r�V�4T�qV��YL�(����L�۶�~˧J��n��J�����2 ��[�^����>v�ʁp�K���v*x^�u1[��l$�F��^�זԺl��e�X��l4#�����(]P��`�!��;�<�c������-�;�Y��%�+H�*�Pb�v�!�>[�2󽌗�`ܫ-ҀZFD�F��aPm�C����zG�[�S4��V�e K��6I� 6��GRn��A��7��6![D���3~��uC +VZӄj��ʰ0@��\;A���ow6��ղ��`�����U�َ��L�Z�������W`Q��"�$2���h�Hq`8�4hm�m��J��@=��#��L4h*�[����p,��4���U�6G�L���Q���;����Q�'u�H^����wnV"���ǳn�VVl�2ֵU�a�,A[�#�%6���EG�kr��D8��l���� f�5��c�l��k*GOj(v�Ӛ��iU�<u� 5ԽN�b�J]�-�9R�F��ĝ�y,1�h��3K8�J�\5z4յ���ƁqV@����X��kd�%��B�{{ sv�K���T�{���ukR_
f�Y�6��7C.�M���R�
�j��V�M�N��`ϭh	Q��Փ�#s�n0/uV�A���K���6]*7$���mօY��B���]��W�k/+-��kA�������nE.j�ɹ�"*5�/N��N=�u�B��i[q'��f�Z�ݱXvܢbT�nhVA�G׳#53&�Щ�[X����u�r�`�I\RTse�c�saw���knL�Z���+m�M���pT��dN���T�$��s��äF�Z��S�hV\,��pU�\֩�tm�F��R�P[�Rz�F�D$�I��k̶H�e6&^XvBS[oPd���Wƫr`ߋ�RdV�KqU���j�<����n�@�x��I��+l6u����ߥ1�� Fˇ+�j�J�5��CE�қ���qH�����7V�ף%�[Yh���Ю�I�#�4��d�z���t]��+���ۥq���o4��B����l��.a*��e�Y�J遨�1��H��TEL[M��tYAV�{Fء�������2�����FGS�,ZRF�nɘ������;%�l�D�9p�v��5�`�(����s6+j�ԃ`P�f��1]��I�EJ��8c��m�H�u�e���X�]ӈ�@�.�0�X�,�K�#2�Yf�$FkkZR�Ţ�m)�Ȗ�y���ɭ[�v�;s%�nV��:qɗ��l/8a���;�_��Q�0�z{��j��W!�����;���<^�Ė��"̢�����9�@��8n�Q�I�K�53����V
d^ŲM�PY���jKG1G$,+]i&Ʒ�Z�+�P{��X̢�:�q86��Ķ�5-�Xl�R�*�*V�b̘	���[�X��m�2��[7l*J��\����4mV��IJ����H�N���	�5������X�;�̵�e�f�a� soTfj6�����8�p�KvU�(���Ɏ�";X3&�:&݈P�uEN&��Z���l�@��0��ũMȎ�e[.����2C4M�wk2�1I�6��t�݂D�%������q�K��z�ufȆJ��������kMKaF`��jԸ��Cv] ���(���P�pܑ�5&�u6죣�����VL͑�/o,��ն���i|V�h�`�җ���leѹ��Gbe�U��a�:4Í�*�Ð�N�^*�R$m�`㤶iA���6����lLԤ˩u��2�x/D9�KjP%x5C�]�ix'x���Z�Z�Ia�(�)dd���î"Qz�����6�U�@(�
6�M���۟];�
5W��`��p�pZÌ�mj�3LW�����v�B�8���s�ͭb�]2�D�&��d�6�Mj�c��)ԡ�s���R�F٠\��cm���Uuyv�-��]�$����2D�q��
&5�W��`���*l(��y��0�8�=x\��$�o��-�u�
w�\_C&I��6�X�J���n��!VCb�ȶK*��R��EѐN��7Uc�w�S�ݘћ��a��$/QUd��g�r�q�U���GSw�E
)D�h�E���[�׷��/#�1�X\`�O��m闩	R��o6]i��K�Y�'v�P��cV����h�M,2�V-ɘU:�ED�w4ݧ�VQ��S�Ļ5>�XP64<X����ҁ�b���"���Qhc���V�կS�X-�� �M͎i�Wt��l�(�V"��lh�:���iJz��0�0 %�q��`D�W��&7&�	ݪKa�OUn̨�%�ٹ��A�����n+Kx�C3��gP�� 1�:Z��!���1����(8��b���R�a2�$�3�e(p�{�
�l$��{v�2�-h1l�G�0�^�R����x�O4���pCeMu7z��j��wuQ'j�% !�	P܄AQ7�F��;-S�:�*�n��J��-�iXd"à���q�n1a��j:�Edϲ��v�<j��Ӛ�_pP��ʊ�T����w��gV��	�c--w���0nI�����{�VȦ[	ܓo.i#+KP�6���pEKkr´2�!,ժ�D���A3F�k�xS�N�`otҊ�����()ФV�P�礃&��`�����Ȓ&c���f��{+]J�]��5�����&X�ڕ�����Z�J,9i��l��w�A{Q��&ȯA�p���>=0$��Ѹu�wP˻ �q_Guy(���� ��9`A�q
b�7�/���&	�4�4�,n`6�b�G7JL�k�!4U�h�Ye�̊�*��U�����l�u �\���e�+,	�6�-�,7�kQ\�P:��q
)32Bw1�M^�N m�MɊA�I�b��5SF�^<$���̟+���1-��X��ʔM�R��_,�#�Q뽽�P���b�(�IL���"�MT���(��ko,�[�
�kX��,��&gcQ��\"^���u�b���4L2��;H���-K�ݟ8����G����0�ᨤ�IKÐe �$�k(c*�3)n��L���صV�Q�-�'����طm�ʐ%XeZֆ+
D���9��I��wJ�z[��ź�#��]2�^�@�Bkn\�z���^��#Ӷhm��'1\���f:���N^��)=	�M��caݑ�lh*�Ǭ 0�Y+J��yn�$�l;0�8�d��Q"�L:D2�����y4MIY���Q! ݦ�̦�.�6���Q�(��L[�jj��m֠�S�X�R[��
�����ǔ��HJ8M�e�I �]Xu3/�	H:���7ڶ��`�p���)�5g#�y�y�������k*���j����H�����B�ܶ���ܰ)�ɸ�6���6�0c�,+�kK�z^<��.�@��VJ����ĉ1�ͷL*�b��B漑��X7lb���+�aڠ/D���eֻ��咰Ռ�ٯt��
Zi[im[�6B4�V�
�$��Z��č��Pۢv��%",�z
2�y��`Rث�X�z��`13��f��&���T� )è(�J`ͺf�-w��v	*\�iAњ$���[u�n9n�TM��0h��m�h%�[�<y�j��,�z�S���u5�nJEK{"��¹/!Kj���%�K��[�v.y���,� �Xղ1����0���(���Ϙ��G�*w�����I�3)^L��dr<Q��T𚻼�#E�:�a!�2����S��4m^��M�T���$=ڂ��KK#6Mb�$ť�w(�z���ͅK�N�[w�LiL�Q��B�����.����#�i��Ih)��0^1f�d�r^*c2���ۓfn��Y6��9��U�����1�q�6m�T5��J�R�HR�LG�1К���i������#�wS�C[Y!�0e��i�I\��Zh*��PTS�b��Y��-%ǵ� ؈Z�/
Hաx�I�Qa��@N!z�����Cj;�*um�[���'�FI��7v�VJ��NQ �6ͼ��@J�hM;j�	���V��]9�̶��P���FU�%,�V�X
`�W��[��_bڎRwX�D��H�mv+fV�M�֞ID;Q���-)�(�;Ce�T����/�1$���;��Qu3{�u�j���VԢ��jn̬r���̔d��V����-�dĥ�u �nVVa(\���G�y0iR��*�t}����֤�3b��:�MW[���r��'���Ukj�[��֥���yC2誺�J�K�m�Te�z�P:����6J�S:�o"�sw`����cU�3T��HVs�>���Ѭ�9�=]�N ��.I�s6Q�5#Q�^�����S6���%`�[��T(g�V�&��O�V%)ܗI4Z�W�"u��よ���BЧ�e
�
����v1 �Fa��Se���wo0#d�&���XK%���U�ӳz5��MX�D)���WRPa�ҳT�;T�!�P�柎WJ`�I���F�vv6�o/w5#2�r�jI��@*|l��r�e�ZoaAEF�j��U�
�`V���0Q+ja�T�+�OM�
O��`����ag�&�7��e$�͓si��Px���˭�j�m]ZʅU��6Pj�*��C
"\L�+��ݚ��)J�&�Kvj@U����&�V	t���]i�r4�Kal.�T&04�P�*y�]��l��)��q��-�S�Tօ��]�!����e�6>է0F��^��q�q�K+�,�eC&֧2�Ry%����eiO�=��'i%��O@fԑm*���m�B���#�1hXP�L�A0d醞����f�%��5`y��7��ꦐ����x��6�S�ҙHV��Hĵ�VllP��v�/k�,z$�ͩE���t0�hH }�ƌAlm�u^Kq]FM�:�+������-*)U�,�Y�^j���NU�R5$�ʵQ�c��7]]��X)j؜�.ؠԻ��j�5�������u����Z7s�b,��d���`d��2oI�w.��_<�_e�#�g��B�bW�r.���7����ܦ�7u�~��	v��Qݑ��묢~H)��_�I��f{:���f[x<�飒�k�(�6�vk�5�P�}���O(q]�s_&��Id�y,�|�ޑ�|�,ȩ�X����O4�}��i6u�ja���NBȡ�o�e:��y�	�㝉�^1��2���=�w�)W^6�W�;�Iۏ��VM�۽�b���\��K`�>6���{�n(�Sg�q\���Z��f�(���U��z�Xp��'�FP�a�xo!	��\3[2��M��c-
��������}'d"���B�._\�����S���W��3��{��9�:؝ܞ��I��Ke:�Β��z�R|��p���ʏ� �Z:�j����,�3VY�"�qj�r`+��M�Wl��hIZ(<j^��YY �m�nnV�1,|���)�R]�n�ӳ��d;
��!�^������<��ɚ ���Ws����x�G��x��9j}={A��J�,C�xQ�W����{��д[��#�Bݣ�m�����m�����?k��涧]�,�3w=}]�Py\�������7�6^)I�H�����o��O���9-=�R�\ t{��h�Y���<�t������R�cwG�G���De����J�P��lu�8[�\�M)�C����=#�|.՛����g�nYU�'#�0dI�T���B�ճ�{R�e��j�@��w��m�|�L9��.F�!:��n��tL�EHO�������]c{w����R��}��kn��y+f�m�����#�%6y�Z��Ư�䩩>nZ}��;ݏ��be��Z�Խy%��.ݐ�֎�$+�*;��6E�yڽ��ִgg��Z��!f���F�����{-�hw�S����텍G��M?R�󳶜zy��|��eme�q�S{������f�:u��ԝS�]�7�l��u)b��4�[W*�_>���i�Ef-H��Yg��FxGX��]X�pҲS���ݨ��l��1��1A�A^�M��i��]@�&_W�6qd����#�j�k]�^C®��kOQT�Rt�D9*��L�@�[�M�(J�9�#-�9K�%��}D��w͜n��6�n�W_��rs�,�%�s�����#&�U��2 ���:r����h�uJŹI؜�捔{��|�d�e�{\qX�s�tM8���Me��iX���툃nL����w�����L`�Z�q|�C&���4�8��;�ep֦w��,��t1)��e��	a}�t|.(�v[��RE��U��Te	ڣsCX�6m]��^���}�nm:M�]<ʹM�AA'�<]Hs�8rk.�s��>�%oM���o&Xv���kt45^��1qu ��;��2�/��	b�t����G��(Xb=�;�q�6�0�]3׻_�Ϟ�ߪI'qW��rԇ� ��~�0}��7!d�w"�A�[t���3[�Op^A�s$����.�;��o;v�z���w%'�F��^���0\S=��N���q�h1���$ɣ�(rW2n�*��r�m%�1���nU���d�Q<��h'��<r�@���[�f�e�ڒ��l�|KkcD����nENb�ܫ�L�}�2�\���*�]�� ��`ws�p�۔�s]l��y!үD�����o��)i��y�^R	��Z����G��q8���Z6�dg�2��x��[z$��]�K���6F>
��b�)�&nG/G�'uU�1;�j���^���<�-��c w{�Nt��
]���:6k$1ի�)  ��c�����&�w!yC��:�dv)Ը.�0ɦ�[������U땉��7;x�,�Q���#��aO�3�x�!��v�Oa�Ws^�Ǵ<[����]��U����q�W�n]t��A�z��X;k[y�ǻס�8J��/�u�N)�����@�N�A�u���,��7۸t�CȖ+Z)����x89֩�Ġ e=k��LKy���}�u�˸���͗CH�_a��l�c��|���^�b���`]gA�^Z�׻����e���D�h5gh����Pۆ���Ϡ79��άj���NAܷn��AχR����D�:Ej�yjkƖWM[�vC]˲�#��SO�@R��`��?Y�ﯮ8$�;���bu�V ����kǹ#򆳾&��V) �}س��۝����ȗ9%��(�
-@΀�Y��Up"����Ƌ1�V�+�j�7�Z�O�4\��,$3j<]�W��N(TN�S�;B����i\�q��/���-J�WقDH�k��nI��N��<���U��C'T!'+ox��٢�ۂ)�Ys[��,Z�L�h{���Zb�p�r���x�0���|ax������m�=�]]�Ի�nN9�F�ܸA��/C�n�v`��o(&��6��;I��=�I=���/-��
ݝ[}/sR�(�,�urK^o��2�h(N"YX�Ѿ��4�Z[��NԄ���a���c�V{y[C����g�5,s�<�!��γ�ݏ�F9-��ޅ!S��w���G��!éQ�����s�}���Tj��W8��x�j���Y�4,��[5:z��|��7��������Gw	WUcdU3��͋d��۹\�h������,��jM8R��)���5E�©{Xn��|��"���a�7�gG��8�WɊ}�Q�f,l���BL�����|�FNOB0[�7�<����:��k��Z�oF.+z��mbt�(	{�m��Cm�n�.he1��4ӷ/��;�k����uPTd�����՘�]ڝwn��؝B�7U,^���a�y����vP��p�E�ٕ��d�Os\��� G}f>RM��Qs�@�L�=��� ���'2.Վ�1�Nc�إ���w.�Em���C;Ll�{!���݆�w6w{��3l�)�ƹ𺎔[��������`�VZJwd2I[[�]f�ʴ�Y�y�d��	�O*�D���l�<2����{���iէEn<�j:������YX��X�h�G���W=�X��rЌ��eqㄑZ��{4�dwoC�G3䦭	��"�ƶ 
���E�m�_#
��Vx��W�KqR�H��p�J,[$NΖ�����[�eO�XC1�O�Oo����ݷ*RE�������.���i4��}�u��]M:@X��gwSe���uu�g��1e����-��e)F�<�+�}� ���o7�=��X7�7��فZ\��w�3�ڏ�{�B��o�9�)Т(����ɯiӱ�$�K���������g>]nOwv�WFn�|o	��z����Vqk�ͅwc��4�es��0r���z�r�R4
Z��:��Bvv4���H9��,�����8��-gall]{�fo�]k�y�8Sx�+�W�+��~r��2�-�q��X��.�N�9�5LYK�V7�SZ|�;E��{L�p�޷�	qR)]n�78sV�.R&���V{�i^�LN(3�S^����v���D�)m%����3�d�"K{��}�pg^������A=�����t��}��+9�r�-��p~�Ƅ�U|��q{��=�s���u�w�&rɢ��]�&�tx�Pl�G
F
�V�����8�ˎ���e���{0���g%�xR�;�.�d��E%5�nM�r�Ac�kb⨱�9�7iVr������
�pJ��B�VX�Ot,�5itק�_]`�i$vVs��G���N4�JZ���>�xwu���'��oM�#���~�E�Ι�(WS��0�-���T�Y�^7�S�.1�b�����t�nJȜ��ڒ��p@i�1^��n���}��p}�TPN��.*�p�i�ש�^nfW��߉�'H���t����LY1,s3;Sp=�kD�	Y��zJZ3]�Mϕ	�*{syn�9��B!��顰�&�ܮt�ON��K��� o�ܫ��C���@b��%os�lٝ����4o�'{�Z�M&�C d���9��ֶtTD��o���ylҗ�Y���w8{o��&�f
�$s�천�>iZ^I�|������_N�A�)�mum����K؝�6�R���k���NCvu'ghB)$s.$̙K�|���i"����vb�g+�ͽݧ-�9m��0�q� uR�n���0��FE'�;9v����`�}��s���޵;�M�U"�r0�q[�=��a��Wyw�����w�������(�.��}1hcO.�u��oה4�׊��˜����d�r,���*��u�j�b�%X���0�姚�%�倮׭�龵?{z~y0	����'�N˓�m��}�u]�����B.�5ݶ�5SaI��F��K^�,4�>�(Q3�a��OK��l�P�� ���pے�����uY�tmJ�����>�pWr�y˫���}S9���^�:oK*�欽|mdݺ�%���˩�mbq��E@��_��V��Jl��뗴�Ѧ˾^|-���p�86���q��K�&f>�h�m\}�����\�CA�$�`��8�X]�w@t���Rٹ+Ed-�f��8U��8_h���:�I��� �V���?���Y���GA�X��.�EՊ�ҕV�yoO*3 ��xUu��scx�L�^{N�Sٗi�Bͤ#P�����쮽�	RI����v��{��"�	0��l�W%�۶��w����̀��k�h�3�����6�!q�vP&mC����ܛ�)�,�sE��ڹ )Q7���ݾ�!%}]NL�&]\6��b��p>㺹����`����`w/�+p�un�\lQ��k��N EW�X7}��H���yA2xE���.�s�kOt�"�����E�0]������N*�댮���4�y�[ZPޥ�%�r�t�j3��/"�8��ԫx�<�E�n���Ƚ��vʳ��^�4a]K���K��;r�X�����K/���$�v.��ƭ�.G��[Xd��t�ڔ&�
��v9������f�U{���p:��u/�N��L��3<�D[:��>�;����շ�5I��tYyq�
v��3�<�!�D��zx�C߻���ICک�&��x緽�F�Y�h�^6Q d�Wf�ҙtx����@�g
��J?I]Ivf���}��E��7�%�T����M9"Pn�։��w���Qo>=�]H̏&n?z�+�4�i!�5�=ֶ�<%���l�gZ�N�ݻx�IˑQ�ޠ��#�*7]�]���/���;>}
�5��a�U:6�!|���aA�GZ75�R�[T�ޑt��/�^�-,_ndX���r�f�G�m���7� :*wo��2�׵{�}�kbާtk���|b�G��d�}���C�f�
�1�s�W3_��]��7e�K�+j�X�r �J���r���9U�n>��H�-��&��r�Mp!_��ܬjk0�X�ռ�>����M;;�`��⊅�鶔�������9ǔ%)���fNE^�����1�nMZ��:䙔�j7��D��8���9ZǪ��}��t��A���ʳў˔W�vq��U�{Po��=J��=P)�]L��@���_����aC+��ת�{^�>�<��hY
��e�n�,8l �	�Z*c�௸D$5{��*����O;u���8��t��q�U��v��R��
Jzid��4*���f�S�G^���ýcB�w�5�8ߘ����]N���gl�����V�-����R����{���x+|��f�X���B$��T�[F�'.�"��Z1��z���.���O�T7�ʖ7Gaۮ=�!CQ�R�z��ݡҒ��_ Zi��F��y�'N�6���|�]ȫ��xk����QA�842/T}��#���,�^q�N��|��L��r`|�
��^�n��c$;�^Wl=:S��c�f����|ҾX��'w��E4��͜o{�F�u�IȆ����y���Q�NgNޮ����>�-��O��77�!O�)�9��l��YCu��v ..���7ǲ��b��|��`v�dh��b�G��\.�R���бAgU�5�v-e�V�y�2��Y�;=�>�{��(Ԕ5K؉��wB�䄔�헺�+U�H&9o�Ew�p��Y�nt�7�����r�y�o'�kX�T��3s������WD��&��LjI�gY2Wz�ξ�Б�9��Gqߛd��D�8�U7���$�Wa��Ӵ�C-D^̹�.���sd�v_8�^�Ra~ELdv#�qK�a�;e�!,Z��ԩ3�D���U��t�摦�A�܅�_{��\XV\!t���d>�_����|��bj�_r��j���c�[�{n�����{���}�۝=���G�5pICŷ��V��a�u�ҙu����ih��2��:�p�}6��� �I���^���,�f�.w���;�
{h*�d
�Q��\�Û���`�gxD`�u�$�Ʊ�l�-���4W��E�4l��t��3V!zi�-�ՠ�2NM���U�)"���:���l�o>�K:�M��&T���2��ހK�e�P��dIp��ڽn� w��9���E�P�YOT��UZM��m��NvtnJnRy���*d|	��e�b� /(�T|뮬�˵sc��Z��-*��P|��(Lꂮ6������8y޴2�q��[�J��9*˲���=���G��oT+��&j)8�x��=�v7��ߟ�ϵ�>�f����w����D�	�����r\)%&��!�G߆p��(��Zsk!5������A"�fc�S��K���6/2hD�)<�u7���1rk�/�L&���Se��;jW��#N�ky��>[Ǔ�]��,���ԉ�:�\�jբ��i�:f��5>�"=��">G������rQ���Y���K0"x��PcWkb��Х(+��L/0�Y���RSk�u�����nL�.�S�xm�M�m��s�T]��N:�&��U7,�l�e�<;y�AU���%*[�Qxr�wNk)���t�7��S��\H.���+�*����sw8���^Վfd=L�r��\��Y�C�6�p��1a���6�0`2�\H�y�{�^=�����׺L2��ԝsw�M۝��F;}%��C�*�>������Y��[to��O���)X=�E
ܼ��rcctqʛ�4��<�ă2|-39s᮳���DN�q@sw��0C��ιƍj&���̫�X��>��#�'(E��`����g7xf�]x�9i�y��j�N.�:v�V�	��[��J��A�t��3`3<�$j�����ӗ6���i���l]ED� �8��B���2�1�1�螻��߭�X���ﰞn����v�jd{�h\�jR<i6@Q,�KzM՞�]�.��$z|i�
�B��e,����b^�s�u}��ǋr^C���kvq/+$��ʭ��Z����Ӌ�@
��Z�9Z�ގ��p8>}��5�8�z��Ri`�(A5)��H���T�,��\WG-5��)i�Ս]�+�.��q�*!k*7���w�A\�o)��I�S�m�1���k(\tdj��C�/��9su[ݬEҊ�)������m6�=�B�syb�о�hTƭ�a�:f핥#�:�fǊ�%d�NT��an�51��X��;���7���s�/�t�n����;!ءu-,�����
u4'�_D���˼�3�]��^����%3�j��o�]�M���7JΙ��7Q�.��{�Ի�0�� ,��.+��*�d^�>�83��>�FA�aƕq}[��@�.1L��3�Y۹Ӷ��n�7��Z���1
�t��4���#�|�J��vY�w�!Tg�Cwsh�X4�5��V8تI�+�T�y�壚Po@�0&��dG�v����[D'v���g-��cFC�)�?J��3*��Ւv�D�r��V�B�Lhsz���ɻ�栽s�{G9m��Z�z�Ȕۄ0ܒ��}�i5��˘��`�b�o,���{�p�^�Q�!��(5���Y���ڶmҢ	0�Й�w�z֙͂8�E�-����
^rN�x���D4��w.+��"�*�[B����Jw]�8����Į��s��:�����2�Jn��1TG	t(V��W���Z�pwY�RR"��2�Ǻn�X�Gv:-g]�2�Y�9]ڙ�����R��6�v�N8]���	ޱ���EmfWj$�#�(�'�����]$�p�8���v��R^9�/u㭛�97h*� @��`�-C8.u���s��
�vk��&��nST�{-�3��Jٸ��*� 
��}�$��EK�`:���V�eK��L�{���k�X�.�ǁ�mo]q*.	��u�o��aJf�7��mЉ�a�/n�VY�X���i�4YtT�
��F*���5���@a������X��;yt����U�tj	��)�Xu����"�6�E��z��p=�d��Vƙ�N ���R�����靗�}; �o� UX�K�X̶�ZykV��W:V�)�4�hbFYVw�W8���y�a�Ξ�ͥq�Y&�~��QYƉ��o��q@�=5�#�V�oZѹE�oO:�՛���N�v�!�$�.�ƨh�zV]�3K5+db���f��l�]ꗌ��'�8�}�퓾����d�^k�l�*��/;M�Iپ[�5`�LY�c{� �X�KN/!�T���<���9�CY���u�|ڎe��{w�̤��Zb��*-�/q��;�&H�m؁\��H�uG_r̋�ʺ���%Ԟ'����R�'a�ޓV,���:�2Q:s�R�q��o0�F�;��x�Ҏ���g^=#_�^Ǔj\9�+�g`B�h��h|Ў�ZP�;Z�Ջu,��Ѧ����r�N��M̲�p{S�e��u���z���V�l6��Y<ji�o�̤Yz)f�=�*ެ��.�γN֌�6�;ծ�\���#��&��g�/���Z���Z[���o2%g&�!ʖ�*����$�	��vE�vA�|7�\ˈ��Y�v���L)�xm$��+'w�q+�{)xg��V4�	� `����(�c�<s���K�7��OYo�y�H���y)��a\+k����h��{𪲎� EwB�B4p=�3- ��!;��j�t�= �����;�5jT�]c�9�
�R��^j� �)qH���}qQ�JxlBq�15�ֳډY9u=�m�W�.����k5�%��t6���\�[Z��h�dn��@{���i�!Qnn�S� X.ܲ��O�m>��cp��U%iH�ɸڊ��Wmm$�j{\��&}\�۴%I*m?kO$�Ϸދ嵁A�R��bs
���2�l�:����r�W�K�5�#�l>۝�#e�A��M�c8~jj���B�H��S�8Y�P�3+@6�����@Ʈ�M� �ͧ0�M��z~��K���gdu�(V� n��-�f�y���,7��HI�Nԝ��i��R�(e�u**��83	z�)Cy��L<%�3a<&e���o,C�M�+C9z��y��;��22�޹[-.ܢu�b�f<{nn���x��[�Y�`>s�J���ӽ�`OB�+�`�,�P��v�Q�)��YV&fԛ�Q�0�j%�/d�����V�љbGڍ��|q���Jq9�e�̩4�o����do{��fM9m7ɪ=r��nY|������ô�آ
sT��2������D�I�/��3g�ܔ;�7	!Zy��{k̦�u5Q�orE�txr�1���h�e*� "_�D1�I��'��6T�m�$�ˡ�q<ܰ��;��-��MS���Nk��#8�.K�Ol���������o1���Up7���� �ۦP]������j�������h���;�EG���Y��Qttou�������{k{w�A>��lgw(�<Ot�N�2���)���{�\r��pwn�}VzQ��7NyE�0�r���EG�ﺦ@�RX�,��Nا��fh��w42�V���'3ϴ⽏.���c���k{�x�)iTܢ�J��b5�.�iV��{1枮Z��a��Xja"��<�^�ᝥ�D�]p�Qю�vQ�cA&��t��srwh-ͮ�G��Ԯ@Z�;*ڊ�F��R_d]���m�=(�zP  e(�םez�z��#��t�8mZ�Z�W{lp�_��o)ZP^��<4�ͱ}�g}k�3�Fd���\�3�kG9Ϧ�^�\��}ʿb�#w/����Uf\��a�����<�C6+ܙv�D6��JV������p��P��u�y���7�̶N�$\��M����8_m�Ḕ��<�_x�x���˄.��	�Kt����v�/�@@�5b�h1wqY�ski�wܪ*����m�'Tɺ꺾�&�ȼz^Ꚏiε�w.;�'ڣ��q��m�k�j6���n�����W'�[�kv�t���Ŕ޳٢�JK;�7�����߄��ǈN+�VJ50�B�f� ��
��<b��y�����͠��̠���{g�f���6� F�����ltO�}���KwT��w+i(��\h[�>ܼ��]5�����g54u��&�&�)���7�E��"�����0���d�=Y�0^�xm�4:Ԝn�0��z��'x��o)�
6���ɕ���N�%yڥn�W0�g�m�wc
����Wkt򑽥a.����sۆΐxļu�#���rb筅�jf����#�s�R��hOtW36W|�ʽ9^
��T�Oh�+�ɠ��d+�5���S��f�l�{+���[� ��'�cx����o:�G.��ӊ�Iۆ�Y,K(ԥNՙ���5��0�Sn���G� ����ܬ�;�69}�¥iS�:��m��
Y�b7F��\��qi�o;dh�/^g~`�廔M��2{/����u�� ��e}+��/u�y.� 򹎺�Owe��J��3׈$z F>�Æ���`&Pi�`廧#�+kd1���V��[�e*���7O��3t�8IW>��/�v�6�S��iv��q(�	�d�O~�Y����Y�\z�� ��:��)�i�V��*f��DQ٭^3�9]ppj�|��]�\�)�v�a6�4�Gov�����ٟ_��U�|�׌j��&EkC�.����}��}�˦!qm�ؐ�N�"G}y�i9s��zl�R�:�6�[���� �3[�f���1�K�T]�e򛺣͹J���8:m������	�I]�R�+Д�r��S>�%�~��zc�w���u#=�v����X�p�",�5j�.�v�����W�3^)�뗜���b�X_-�?)�G��l�<�����jF��8$a^��n�9#�=Uz����G)�\!5�⯶=�ԯ�R1�;|/l�u��`����(���ڑ�Y�ț3xN���A�y�Fh��18!�溊�����`b���Mo�������&�B���`���wj����w�Zl�26�׻5*<���zw�~�y�O�>Ԝ0��J�8����W`d�Ȁ��.vͫՓ��8q��Yrf��;Keދ��f�<��/���ݥOCas�� ÓP�R�ڂN���������l�@R�F��w[�k��]K6Z=ڧg�7v\�ۂ"=P����qna,O��2��v�¸��6�`+�k�ۙ@��0q{���(Nd]�.c��wq������)P��L��Tx��h��  �����O�hJ����E�ث�cݛ$�o�H���!�1e��mς���]ԗmG�:E]H-L��4N�J�B{����?��X�8+�f���{%�~[�9U�\�L���o=l1��G`���W�^���M&�2wI%�=��{�Ճ�{YObP�y{����x�휪�7�<���,���Λ]�š�f�z3U��8e�9���B��*�h;�iT���C�[M��@�v�	P̋}D� bw�9j��we��f��EP�
[}Y��nL��7����Ҿ����KgE�Z���y<�l���Y{��V< eX q�LXoL����0��̜�"ջ��c�`Oa7��Dmq(g���Y����̫���r:q׸��� Z�����v*�����l;�������}.��"�������V�7Zw��F8�
��r�	�5��pn�I��]k3�mլYr��}mu��T_p��J�V���霹z$�ZC#�{h�~��|�ȃ�vY���"r��{�5����Sd�(k�Sڗb~���5`�"�ɴ��$�%�@�5�ZNav�ذ,�7$3(��"dX�8>[������)G]����E^��tL+�[oKg��F����ݗ��#�ݤw��y%�; �f����f�_���-W4&�F����7��[҆C�-Ż8Ԙ���=91��E�gJ��Ю�Y��[Ԓ�쀝L}��N��KG%�h�����v�x���x������~����/u�E�lB�5�*�q���P�X��b��.vo	������wķx5�:��)[���Z�&�]OtB��k�X��,�g*~crQ�J��w����}�@�K�{Z7��f��:�kh^��u���RK
f�u3�n����2w��ow�ų���t���yz����-E��&�C�Un��0:��7^�}x5&�ً�L_KN���P�R'Vn��d7��4��������){z�������N؀�v��:&�wݗ��-��gR�P�X�Ǉ�Av)�A�3��*ޘm�nx��>�=p+�f��$����z��:Д��K��m�׳1S1n!�أf���]𻝥J�G&�̷ �14���4�;��G�3�sge�|�����Q��������Fk',�Y������Ϋ'_5O��<�.le1��-�����S��0�'�B�,���i�y0��HâI�(���s���{8NȌ)j#�S 4� G��̱#^�R�S�Ϋ�Ý��w�7�.J^��c7���{���{����Ƨ�b��z��R`{��"Dg*���i�K�7��G7F^�l:,�r��z&=&Y����c+�t����y�w��!���tb9ה�=�\��>].x��87�q<0���]��cGgqf~[ު�}�Ͼ'C��a��|.S�Z����N���(������ޑ@�K6�8zy�����B�R�wd'��Z>.�ڇ�e*�e��u�_*�ۊ#.R�x��TY[n(S}f<8@���M�F�{�t��3j�d	}��@�l���
-�5p$��3�A��nN� �{�����=v���Z���� ���3)ӵĕv���/2�#�J����d��(&�73������Ȗ:��O�� `�LTt��������"ՓǤ�Q��sӋ']�N�9ٸ������8,`�|�T��-�v�\�Zx�q�g@�0P��[��!����㞯K�9�)�{Z{T_3-r��8��nw�W�}_U}瘒)::��qtB�7�(z�V|��c��%�]"2��)o!.rviB��1guк0C�t%�)��zM޹e�GK�k7+�
ʍ�LL�/[�35^G+��}`fZq�վM�\{xU�ݘ`��Z|-s��:-H����D�eF�)����3��b~gʩ֪�{�:�%�-�Ӱ���i
];&����ǻ����*��g*`+oL�:�4|n"�R��݅]v�|a��.��'�D�q7罼��^`,t�{�nv\쯰���D�n>]���\@�D��I�;=�V#��qS�f������w0��Yٯ�{On�N >��.`�������8+ї�.�����+�^S)�ڴ��j�'�'�ڃ�����^I)-�s�2#ձ�٣��1Y����Gu6-L����2.8s�
��=�.���p�C��'d#w4�2����sdK�Ԥ���6�b�lix��Uӥ�rR˶��bp�Z/N�,���v�{����@�<���g��MɔE�9ʟ8{רۧl�ЏwT�ߍh������`�J)"�ݢ�3��t��:Q�^{Y����}�Ԃ�gG�\�]n�Ns�x�j��`���űT$�m˶�j�g�h$�@�6k��Rn��#��B-��-���1,ˑWqV�w�L����-�6E�q�E:ߗ�P����3���""B*"��#,*&�2�H�&���JH���̨iriʲ�
����L##	����ȡ���&���b*a�����+,�����1ʂ����&��H��h������"3,(��s1����(���2ij��1ɋ,��$�����s2�H(*32(( ����b*�20,��Ī� ����������
�����"k'(�&��	����3���r2�0�����*���3
����$��� ��3
���**�j
$����� � �i*"��(*"�J������
��(���	��ɪ�02
��)����&h�(��",�"f)�(�h�"&"j*��H�*���Z��bi���b�(�Ĩ�""�� �&��Y�)�f�"j��"��((�*"���(�������"���$���������iR�CΞ=|���{z'v��	�\Yw�wD\�%Q�u�y���ゎWW7ZWV�w,�$�;�8�c�q,�N4ŭ�R.�ڇ�`��a�����])V���Y��4pۥ|d)R�2�k��Ed��ty^��E�Yז�3TΘe-	���	��H��a.���du��u:��.�Yw�`�f�9�@�V{eј%a�©�t8)�80�˻3=��3 ��u!W��7��&�����X�+��7vf}���l�Ň�t�Nت�Iz�kY}�3݂Mj���؏l�������~����B1��q�o�=q�E��z�M�=ԧ���`��jZ��yu�^�N��^~�3ٛ��-�|�,�q�~�t����f�y�8g��e�{'3k�Q���>ggH��z>�U�+�X����r�>{��n��h8�po�\;�y73Cgt!vmUl�ؙ�ݱՍ^u�dO�󽇽���o�E�ޏj���
�;�Ž�C����h��m;]��V�,g��<ܰ��G�y�h��[7=�z2N�=�!������##
X�p�sީ�\�i���Y�N�+gvΉ]Z����S���������B`���rň�ӫ�L������UW%��ͤ�[�MJm��N�դb�ҽ8ghX)�P*����+��F��OK���8O���|��}�1�n�ٰ����.�.kO�'T�o�+���A�zop�80��;����]a>4;�M�W�����rZ΍XPcޫ�s���m���t`:�9о�*�f������_����o?{�;e�s���5��q݉�R"9����
Y����߮���^>X'���z�{پx�λxK�]��{[�9��}e��7|-�]�v����w�K�K�*{vo1��>+='��7�:��վ��'7�:^U��"��\�y=�����R�o��}�i�y��|#{�%eǄ��g��{)>��z7D����7��/NA���z�Z��úϷ�k��~�u����������߶t�������{�gn{��܀Nh�ސ�,1���m閬vv4g�KS���={;�Պ��&�����c�����ͼ��y,]T�^�j;i�M�{��(��C@;B�>=�jJ�3����c�d�ۜ�K�v�@T�����*]�7:�d���/"򐁎�,��E��
j�	�ó�u쀭(L�b�O��R�ws��ݞ�K%mozX�5�q��ǧ�{v{��a��
�}=J���Ď.�t9z|��S�T�~�c6��n^�q��=��?*�������ް�ku�{��z+�:�������b�A�m�N_�G�6�f纼��y1v����k^����7�M�����(�l/�c;��c���y(rj�U_���nzur�C��#��}a��4�/S��_�����w�V6]x'��wnsi�<�Pnt<�����gN�]N�֓�E���ovw<��0?=�K��M��~����b�{�Ύ�Qռw=v�y܌���.�f�mK>����c7������9��}��zgW>����<��{��dJf
���*���~ �~�:��'?\�.��f��]Ž���ѧ�Y���a�s�D+OV����y��+=jv-mרl.e�;��Yw���u�s��k�+��Sx�ii�̫�il̴][[��F������='2rHԷ�ݛ��(��"���U��aa���vt�3�8X�5��))��W�9&ī:b�G(s2j�Y���Vj�2�Č�=�54����h$��獡�q<�"}[/�L����x�r��Y�@.�I��W�O���~��������y��]m��Ю��Z��X%���D��X��w��*g�t��Ɵ~�^x��y1n���s�3�YfQԁ�\ϥ�ޖ���(�_�}����י��F��q����zr��Ai��v�?{]뎵��s �2�L�U�)��\ޞ=��?N�<������sn��_��ٱ���r��+��s�n�����1~����K�6��B��'ۭ��^�R���{�~�Z�zb��ێ����z1p8���v?/MY��Q�J}��}��9�k��x��j��\8W��
�FA�v����]X���϶ܴ��ϧ{>qǾ'jx������~�c4��~%�gB���ڬ��U6^pl��rӝ0���k�9���a�8��K��o���D�ޛ�[P���yP6�I�v`w�_]PS&�U���azzN)`}�ڋ J����FL��p�5�i�7��ZO(��-�s�z�=��
�Ѯ�w�Y݉��-��4d�l���oT��1:;"�{gZ�N��7�.����So[�XO@�ۦ6�����M͘\�i�5��y��Þ�_m�N����{�.w��:
V��;��Lvʥ��پ��O��娠��^�fz��tQ�,!΅�P3n�;�=���{R��%}���mdn�j=~�Շ:��"5*pwBtύOd}��dp���k�J�1���;�%��^`v��7Fzj֋ש-3ۤ[�'�ϱ��>�y���;���`�6Ĭ�Y':�dR�K�����dS}����~�9;_�w3�Կ���EM��496y֭۬����E��A�Z����cn��:�]+/��v]�kF�nEr[�,�֨Vd���������G�0?�ò���ԧ�ݹ�z�Uɼ����2��,G�N�hM�_u�z/��.]d��ɅSwZ�f�{��_<
�m!���8��@Á�Ǚ�T��YK�6��ϓcg�P�c��̫.�&�`[�q$)AGfZj�F%[}���V����ǰ+�����K��=�mv��jZ�t6�@u�u��X
�9��7�T�sQ��=�gw�#��;7n���y��| ��\林�0=���r����a?N�ǵ����ծ�G*���r�\�Vz~6������ld�����no�\ư*��ݔTR��t:����н������������q�G���y^!L�y����eF�[�ƶ}�׬/S,e@�ы�f��Ǜ���m���.��^�����;���VP�;/WXKe�L!N��tw�a�n]�)u�dy���꬀��湍���N�c'_�J���VF��A�5<��LZ�{T�%��}%N�;u���}�'���& ua��g
N�r�]J�x����9�3`Y�`Γ�t����yx��u��G��Lѹ�D}ܥ��r�����5��P��ʈ�����g��m�Ux�<"txJ}봷��ސz=zȔ!_,ݰ�:��u�ۼ�7+=���$�ۙ]/��o4�����Dt��md��+(���� .��w�y��HV��[�D#��]�,��pU�W�A�X瘃��ۼ#R���7�2�O���7Ҁ4E
Z�^��G��ў���=μ��+7�>K/-�J��Y(e��Fj�K(R�L�_S���',��~�F�	��P�z��;����w��o�ػ��zY�������xH�ܬ���}��?^U������W��b��6�[��bF{#Lk���̸��:��K�kh��z�JY�Ckb���;n{}��y����1aǦ�A��̵vw��噵=�������6����_��{)�����C�9�N�^��]_��=�η�N|��ك%�Qк�yQ׶�w�y/����q�ɏt7[�lg�y��ݷ�'A����?_��Y�g�G����w�|�'/�
���������Vת�o�SމVrok��6.�f�!y�Elc��^�.���ϱ7犺5yG�\5�@q�=�Xr��5���C��ī��{��̿_.�uuFl:��JΙ�rziy�祃g�;�mu?+���
��w�֭!�BPwD��E�穩���[|8�ě���tS�"���WǠ�u5�$��ȹ�%���6��s׬-eһ׷��t��r9"��=闦���_v�_#���v�h3�}7�o��F� .��*tg �K�>NS��gI�Q�b־�Z�I��9�}8��v.�G����grw��{lvNoAr�SlS���P�n{ӌ�3e����gH���{NNg.cv}ӪE�l�!}4��7���ԙg���,I��ݓ:Q�Ե��~�5���v;��,L#�Ӂs�&V����<�����z��Z�ݗ8l��:�nvנ�_\�[+��5�4�u]=���ݱ�=>�q���*��$}�*����q��nM�+vN}��{(e���{M��t̩��{�7��}s�n��W9)�x0�9�0�g+�^Q	U8�W$�_���7t.�&���F��q��c��f
0T�^Os��WF{����{7��U���;���ǆ�����n���������ֻx9K�.�rh�u��=��~��Q��������n:��o��^��m�FK�O��hD�Qc�pHm�nY��-8� ̦ظ.�W���M�bv��^U��g�G\�����P���������LN�w������ƯQv>%�gy�Uw}�����.�V\���$#E��	�%�ӈ���n�E��5��5ގxoo'�M�Yur�=�ٞOܾv��J��}C�=�W�u��M��	.Tr���͌�v�[���䲖���)��-������[���|3٢���pm�a9v�w�8��}rv��+>�:Ι��kO��d��-I���9��>]���V��ٿ7,�@���M~�lܽ�k�ƹ��n<R7]�eCg��K�����4p��~.�nlNs{��:��I=ފ���<����a���D��[�����zr��ZO=~�t~q��&�\���r^��Ͻ4̯X���`!ί���b��ͱ[����M���ڭw��]�'��庭u۞RģF�	�>5=��j��;�����b��{�{�~�y�:������m��*���0k:e�;�r֐�/ �#�kW�O���>���U�9>�%h�snV,��,�nW<;��̺�V�ӂ��c���n5�.̬���R��qE�uytx��N�s^��=~�ɓ3��f�V�e��Vz��Y�=x��y^���5ZU�?n��epڴ�F9�h�D�r��wLY��|��Z�	V��5�k�y%���V��mga�y�>
�-S���&
�	��¦�{�r��5/��<S��z�����:��cnq�ȼ�q�y i����3��ż߮'�W�ȭ�Lܝ�*���ݯ�V�X[X ���#r�{��r_�o/ꎮ��T7�U�ڕR�޷�J����Ӆ��OA훊�ͻ3�^X�~.�S��Dޢ��|�}Q?y��g��u������9��s�3�6{����٤��t��E��|�_����|_S��ۋ�U!�{�=��I�G�s7���(�v�/��yy�q����*qJ=�.:�ý�z�@��7��q�&��,~�����͍����/_�Mz�^���+я�:�p�.��F7ܥi�5��{�U��oI��O6�����[/�b�;g��y��ߥ$���z&�Aׁ�wF�vo�.;x��y���h�d�Qt��Ud��[�]��z�����*I�\�Ca�w	��ڭJ@Z��`M��ά�z��x��>���:8����U���U�.���ǻzѐ�-Yc�GT�s�sٜM�c�S��Fl�������z�ƈ�i�1N�j��� �*Msȥ����گ�cqxy^��V-�d|9kض�٪�*�7��<�n�y��{};5TAtˇ��M.��g#!TzqB�%fp�p`0�&�n^F]�[����>�w�@S']�)��F��)��m�&��X"뫑��,d��ku#']��8�1*�E3[Z�R{��X�cKµ�{��+{!횽諺g<;��qH�921X�U�%W�a��Ur�z���Y����@QS�K�l�y���[�q\n��M=�<�&�0f���I,����n�R�z�\�p4gV�ćư���g;[W;:\��ĸ������(�)/:�mMXzx��s���t��m�~��r��)D�v�ꝕs5�$�T��P���)���]���sdO9��Tx/u�]���B�hi	�ui��E��b�����e�aL�6���
Ե�����ۤ���V��@�n�V`�����wn&��#V�L��y/�ۗ;�q+whq�J36������Q��/���th��ˊ�ΰ�v|�W`���7�����3Up���c�{6�Njud���/2��=�8�Eb.�{��J�˥R�S���)V9�c�R����R���+�S9𳔖��RZz�|f���W�;�����=b*뻝��\A�ҹ�GM�L3|Z�4��D�Դvn�9]�	��J���X����:�tޜX�l���˷�H��y3w��8�&�k�nV���Z�{�=*�S���{\/��W�}����%��h��jD"l�[o[����$47�l���s�56��\{	���՜l)�=/n��+�$Ꝉ�s�[�JB�K˧�.V�"�IVɷ{+��V����r����VK�^H��L�a�r_n軼���δsE�T���������H�=�a���t���&3n��>��lv�H+9v���^���t������3mS��P�cE���Z��T1U��rv�	�5��oѩK��=��;�R��ҏ[1*q��C�R��i�+���oN4�؜&!���v!߰�� YEa �e5Z�0�^�UeGw1r��y�Õe���Vd�Γ/�r��i���u��vΥ�����WX��SY��Mq�fH�(�fVZ5r[��T;#�W������>j�QԯTz�𪸙�uz�⤛��2�taj#�3[�B��v����;z^]Y�o8$�Eu{8�{�5�.���n�Z^6:�8-�p�Ytx^o�N�!W���p�"�P��d�=�K���Ovmt�뇁����{a�϶bħ�}֌מj�i���J`�(f��b*
��( �h(�j�&�"&h�����*"�(����"�����
(
XjBf������d���&� �)���a��I���I*��)�bf
�������(�&*"h� �$���h���*j�( �b��)�h������ ����f
" �)�)���f��j�`�
��!��
������f����h
"X������&���&�"��jF�������& �	* �i�jf�����(��$��&�"h"(� "�������#<�Ύ�׺t(�
'���7�)pC�-�W ��Ӱ��ЦOd/�rn��KӪv��;�BT;7���0�X[ڽm�Q�l������ڶ�?zq鴷�:;_:(�Ǣ�{�/mLӵo��ն�垎{Ӥ��r��m�s�x�J�pE<W�nn����x���GB�'����^��vl�ݏzkp����$m���R��N|�v����p��:x\/��F�~���K�,x�z�vt��k�iOv7�݀7���w긮��=�y�pS�g�ɑl5�&��K̓��t��}��o�Y-�+Yܴ�U�Z���Ƨ<�G6\��oڌIILX��pz�s.c�î��������\%�by�ɴ���ۙ��^��#C�c\zz�s-_a�4B��@�Z;-���x��t=C3|�L������z�41�6ǧ:oN��M�yƫ;r��o���[{j[uG�|�*q{����J�=���T��s�����-�V ��v<��іB�x�ӽ�y��+�����9o�:���`�ݧu�J���+o,q��ik�֜�%4������h§)p�/@nz�쑹��5��n��K���1U�<ўß��&y6w��Ը�7�ư��v�|�j����)�-E�N�Ϗ!u���Ս{�<����K����@,���lx��������>r,��͎�S��8�7��/N��wq�{s�~�}{WFN�'-����q�I�ϫP�5ֽR��I�8�l{f��mr�y�~�^�Z�W!�o��Q΁ɜ���d�g�����ʱ�v:�x@���v)�ӧg��\��z�4|��y69Ϝ��]��i�f�vx/s��|�=�eB _�ik�R�_g7=�S7���q�f�eܤ�=�nt}�����/A(�gF��{])2�7�zL؝��7��<�e��>>�漼���M�B��y����<~X�g�D�����:%;�\��w�>n^���d��;xW�Κ�U��xV��ǵ:nau��R��f�v|6M��q»���J�/無��8���eU����ܮ��&������fyC�X������W�F�=����[��f]���i��,�8����dT��b^]�=�]h�\�����ۈ�N�"�����}(IA�wa#���}�&�JCD<��9)����
�{J�gK,���UB���]�ρ;����x�<����#�"�,8��S�s؁�]��k��~mú�d�&=�Ҁ��y��7�=�8Ã�����w,WS_+�Oj&�Z=����?���dCԷ�o�O���oM7�Ewn�H�}iܞ��݃�Y���>��L�}�+E�.�ӬQ��1{r��cJZ�>rK���mONc�3y<����=�����������/��^���j��{*�����r�n_���G5L����Y��s�;��*U��'�Y���ˍzT�,w�C����ӽ�8��\���?/���s��Sw�W{�sdm�gˢ�h\
�L����0���_��YɟpǌL��կ`�Xl�Y�a'Iz]1�/����m�3ْ�O.�k��?����v�.���0JaS�>�'����i�7�&��/3�ki<��9_m��YA�]�XOQ;�FN��u�f��+'vC���ϝ[�r�,��˘���e�u���Q�'
*#��&s;��z�3�z4Ԏ���ո6�{ݠ�ث��*�M��2���G1�uɳ��pf���+����}�ϧmIp�{�����N���ֺ#�Ί\#���x0�g���_�}%e8�~�{�_LwV���������q�H ���dK��E�o�V��/���y�;����z8�Rjx��풿G�Oeߘ�F}�>���;~��r�#���������_d�9� j������@ϧ�� �>u6����~J�jz|~�{Ρ�NC�Xp�/#�b>���z���]���}^�t{����}'f�h������@{�iyK�~��>�@�>;�ï���_)�d��k���u��
P��Z\����9���k�w.��C����{���?>���9{/pv�����9'\ގ��}�����1��W׃��N�n8'�&<}�-{��(:��)���~��zy���R�������]�����d?K伿^��G��:���w'g��NK�N_��}b���U����㿰2���w?�O�p�=H�9��:�pR7��ܾ���Д>K�7��J�N���˹^u��������q�9.�=���aB>�~����]f������#O�ps�k����h��G��G%�
C�|�w��r��P�/�����_��Z\���^�h{�����B�w5�=�@�O3������,���h~?C�9g��#�~��~о��:�z9 w�9/ѐ>�{�p�9f��<��z}矾���`�.㳝�]sz����ζw��>�ϵš�ԾFI܏�����Q��^Jy��/�r]�]��h^���<�ҾO����w�w�!�|��oHy/��{�Z�7�����eg�����\ͩ��s�Ou�.S
g��ۓ�є�8W.��eׇ�q�P5��D����ĕ���䋛��6�k�V'T-d��O�J[��mE>׃�[�uo�+�g������u2���t�L"e�]S����M����������^���ޗ�.�h��d?�<���=K��5��/��ܯq���!�W�j_����_ 伓����:ޞGR�Of�����GƄÂ�g����+��gsǽݿ������u��=�ˮo�˩|����C�'�X��^GZ�p�`n
WG�4�pR�ߺ���t�������~�����_�71��s�c�C��FY�]��x}.���_���/w]ir �����&���)�~���XjW�9?�7+����d�^oo��;���x�S%K觸��������K��G/�y'y�<�p���7W���~]��;uޗ!�%���!�b��w+��<��^�κ����umZ��b]$���!Z>��?Y�A~�����@�^y�����.����r�G�=ޞC��|�ßZ �_�=��jW���������}���<��#\���Ǚߝy̾�Ͼ���K�d�P���5+���7/�r�9��r�^y�ϰC�m�z��]�Խ��|G�}?P��F�����(��9���
���ˏv��\" }��_B?}����`C�?OF��y��O�w?��=��r���r�/����	��{׷����;���^���}���y��vus�u�޺�{�>���;��;�R�A��z����-/�����?C��h�~�q���B�w��`z����>[��ǩ{��:����7�7w��s�o;��g~~���Zq���qK�w��]h)_�����d��pܙ/���u��_u��؏����$Y�|?�:G�~?-�k��&�O׾�����׾�����Nw����ݼ���`;�4���
z�Jre��!�}�r2�rd��@w�]���Z@�q�����ɛUo�?0�ٸ	�X`͡�q��g��kژ{��s>:��#euv��KN�a�CB��{/����j.�Y��߷ҟ�[���㳱�E/'O�]��S���z�*�y�����`��G���\=�!v>�Efp��.�w�fDs/ׄ�@�)�~}�zk�o���;����A�w�����N��[��d������s�C�(M��r�>������yf���/����w�����|����}�����Ժ�w����4~��ܽJu�C�仃�ߵ�]FI�����_��<�pP�o�Cr�'_sBP�W���>��}c��Mqg�n�w�7����{��qr���hw!�1>��=]�o�N�ܧQ�r_��'�������ߴ/�rN�w��R������?���?}�#�����tkW�7������ }/>��Խs�.]��:>š��� ���O�nG�Xw��;���4��ԿAv��^��IC����ߺ������g�݂���/q��<�Aܛ���|9�!�K����:|�C�}��٬G��z��c�_##�X��r?���;����{�����Ѐc٦�����w���_sڦ�kh��9�h�z�������G��hܼ���|�zC�}�۳|���t���d��?f)��/#�c�_##��|! ��ߙ�1~�7𪘟�ݷ�s�,�PP��)켌���h��:u���w'a�h�^H���w/g�iy!�>]��K��!����C��k�KȻ��y�gy�������淾��~p�5?��
��������C�n]�OF�Ї ����د$���似��9�7����~^@,��G���
�)`h���,�k��|��0�/�|�k���:5��y����_��7/ђ��C�r]�A�qL�po�y�p��r�˹y���zG����)�e�������]������G=���9)��Z ��`�A�w#�?G��7?�~��'%�S��7.���s�)��O�;׷п���^��� �^R-��O��56��t=�_�
�\j7o��xv�`�o\{D̋&9q�{��<7u��:�}Jo�_gⰬ�m�r��;R2+)��W�����SpN��3U���>��vÒ�"�IaU���+�w��,������_cr�]s5A~=�⨁��{�o�f���?�j�_��oH�~���y�5+�to�� �~����a����~ъ���Τ~�`r^]�tg��n��*������c����q�?�eq����P�s�/#��W:�~����矄9\�K�P:����.@}&����������|�ʟ��p�q�s���z���ۄ�oO���py��;��^��G%�O`;9�/#�~�����AԽ���wF������|G�AD}�Y��W���0m�p���a����{��p_e�p����A�9y/�v�����r�~��<��|���Od;�4��}�����=���AH��l����ޝ����ۍ�0z�w��r]Hs0|��w~�H�/���W����|Е�I�~i\�A���y'%w����]�Bto�J������U1��?ws�Y��߃��Io���>y����oKK��C�a�|5�}!���Wr�.��=�H{��=�7��;�<�2=���#�U���Iw+=��{w�Y��H~�� ��Ҕ�K����u"tw�α]�{�����k�C��w��w)�����p����:��v���#�QJ�/)2��?z�.Y��gӔ����T!r<���c�?K�d�����s����^��K���������7+����܏�<���MÞ������v������>�>� ��~�>��9'I�����ѿt��Ju�4���^��@y/���<�쮥����w@�y/��X!��7��o߳���Ǔ�ڗ��Ѫ�d{������~"����w�<���v��I�{���W������Ju�4n^K��>u�����y�_$:;��j^��z������?:��:N���5qՋ�0mުlJ=joa4�h��b�!�j�ވӐ����x#sn�v9�j�9�YV6�v<g�Tf`�]p��T۫g6.v�ڝ�	���s<T��%p2M�׏�zwL[���1c�a�H�S�U���ǽō�v����|*��o8s�߳���R��`}���u��!�����)z������߽i��:��r:�:��y/�b=�7/%��?�����#�;��ާ-y��m�`y+f��߾�޾��_d9�-.��αN���NO�>����&�t~�A�y�i(w.�#�7�w'$�[���^I���������e�he�������x����}���}/�����ԯ�z�C��	�1=���?�:��w?�f�|����؛�����'��rC���JK�7�}���Q�����l����4��~�>�����}����u�����o��{=}ޗ$��b{/�RP���w9d��n>?br?J�u�M��������ܝM������n��!��~���	)Jp~�z>���/[ގC��|�ßk$w���w�u��s��$�S�n��)?f	���ӣ�M�,tG1I��6���ߗt�_���}����~��3��似��}�=��<�G���^���m�ܝGf��wKϻ��G�{��\���7O�@'�~K?C�W�;�?)q��G�/���r{?����_���'���R�r����r_dz9�[��~���yK��Go;�?OP��矂}��U��Z���cs�k���˹��"�W��;����a�_��F#�}��`r�]�����C�����p�_Iٿ�:��~�ܿ���|��:?|��{�ǹ?o��3/��v�� i{���J�:���^�sp�>�K��^K��Ԏ�<�^�<�G�?���9{/pv�����9'7�P�wv�ֶ�a�ο�&�E��|��ª�bPj_ ��7�y��]h�+�<w�#!t���~��X;��y~�����:���w'g��J�A����6rbT:ɾ��T���7xYUae�qmaH᫬{��*+���ތ���5�J9o�n�J���7���.�p[����ֹ�+��}�eɬ�� ��ħ���	���,Tq�5-�t��ԣ��W\ź���!��np�&�qk˻;������_���o�yכ����WQ�]�G��GQ����]�Hu�i(7/�S��4%����R��}��ԯ=�KK�x��X;��{���br^J=:U�<�c?*ps���7�^��!�au�t��ԿA߿kr�������)\��ގK�)�|�w��r��P�/�=��ԏ�z>�K�r���KC�䇙�ƻ���ל���}���~�����~��Xy>�ԛ����Ի��������z9+�����F@��i����s�_%���~�D^<����O����L�˜���|��>��h{�/QѬNH����:��?���K�9}y������Z�7F���ԯ��p仌���/�+���5����}�����}7ϯ_���ܿK�����}���4>ڇ�w��{����X�W������w��>���������%�߽h��:ׯ�´}��|_��~����oq�9xת����G�����]���\�K�>�ߚ]K䇾��d?��z��~��Ѭw+��~:����{�仂����|H����#(o�V�8rW����8p�������Gr_a�~���|ѹy����^B�u���/R���r_�n��5/��ԯ�r5�	��D�uE��ߺ/~��Y��y��~�s��<ҙ/$�����/$�7����G���Cp�}/i�y�y#��5ޗ!�'�0=���9A�@d?}��B��߽�s{����ٟ����?F��5+�y/ђ~�C��]��ߛҔ��}��������?[��|9��|���}��ԯѽb�?BY_���D�~�C9�s��D}���>�ġ�����<�q��O����Z�ܿ]�u�h7.����y&�w�o�ܽK������Wf��wK��v�h�~���3��4rVm���Wd�y�1��3}D,t�N�V�p����>/f�^�&�kV����|Y7S&�'��k�zV6:��&`ܕ�Fc�V�w:��@��jx��,�.��S����Y��]���� �fꤲu]e�*���蝹��]Ξ����_g��hr
\��2_`��9!���;��{���X�˹N����>_A������o����?|���%���ʙ߼����>������}ޅ�u/O7��y\�C�P:>�pd��K�C�~�$w/#�O�����'��y)�h܇#�0�&]��}W�w�Ӯ�}G︣�=�K�>�w��y=K��]��@������+�:7ޗ#$t>�2_c%�� �K��:?b;���NX>��*����x�?�s�,��g�VC���'oGҾۓ���u'%w�K�>@{�i(?K���iNA�s����=o�.FB��7&K��F�w/���������h��]p�:�~y�8���y�=[��~����?����rWQ�~��rNJ﷙��;���|�Pn_`�|�({����P��}���}���Ɩ���7�-9?l��e�s_��\��b�/!��w�ܦ�c��^����y/P|{��+��<���˛ǐ�	�|�Pn_c$��h������w㟿~�o?F�D����5��r:��}�r��r��u�NHr�#�؝K�O�a�r^�ܟ��;���O~�$}�$�xr
W#���︄~�W��y6L�{5����^�C��]�I��%���}�Һ�����w#������z��`nW����'RnG��G�y��:�K�K�/h}�?��~������FW�!�w����ߺ�)��{.�%8=�A䛗��|�4���/G���Խyއ�R�/#$z����k����9&�t����� ��o�m��6W�|��}�q}��z��ο#�<�7�'�/pxsz9.�%;����y�oHy/��v���a��u/#�X�s�
�?x}��Q��ٯ?{��"W��d/񦺲	�����OlM��E:!X�GA����FM�����]�!�ڰ5��
Q��N����Q5��nᢳ 2q���5
�9ctd��B�wب�sUXG>�oo�P�h^5�/�K����v͊.U\��A�ѹ�D=-�^7��z<v�m%����K'g�k4����m�d��@��%��+5V�%7�uT>7�Ӆ�AnZCn���N��5)����U��j�|�Ė�<�m���vx���P����F�k6��|7�W�eSuC٥op׸���!ZkY)���f=���t��di�o�,J�,9��zk����<�����C�k�hRμg��2�t��%��|ޜ��7�=������r[�<�d�cM(����-�ܠ��!�,��''R_\Ռ�1�]������YUE�֦��1C��f�W���ک0�TKQ�Gk~�`c��륞�ήh�?�3g!���)��Xx~>�����
��j<iN����C4C-rQ��*���T�˒;
u=
�y��:�Eᨉg�'�VD{�ﯠ��N]���Y�h��?w�q��.C7��۳�D��K�U��r7&�����B�^��K��(���Zߗt�A����#}��-�����&j�χ^pE6]�{H�7`�GH]�� X��;����m����t��yc386�E�en`���Ni%L	[���pU�^{}�w�����K�0Mڈ�����]:Smi�Ǧ�b+*�����K\9r���<��c:������.Rc�-����#t�ËV�#8M��|�ӆt6������mx�dԳxaͩovTxop�0�]e�t�#�u|FG7|��N]�mV���۬�x�L�OF�oDg��
=yryJ�\�Aa�H6>ޯ<(|tU��<M�c;����fm'��Pݽ=qoI^�'!�u�0��R����k5e�c��rc�Q�7lv�g
�\->4�m6���s�&��]tO.��o�3N�+>�����	r:mvT{ǖ�j�q۸>�VsK�2
K�!+,9�͇ü#��"��~˭7��֛�������kv��d�S�{�W-��EK�FVs�t�Xn��<����OE�*�x��ɠҗE��g���ب���Dj�_&e�$��w���O��v�+�F���z0��s�'R4o�′����:6�!��d�o�ـvt��V��l9�r���dDha�G϶�-=]s�ԙc%D(�jnR���Μs�ᠺ��F����h�9��3�wcK�m�t�Z�j閶��\,p�rR
3�]Xd��h�r���H��S���)�p���B[��K�|��=a��IbN8b�2��W���v��7���]3�o5��d��Ef!_!���DT5E4QUILTD��EU5U2�Q1-UPDTRPT�5S1Q1DPS4KL�5M	Q1DUQIQ�T�SP�@U��LULA1ESCA0��XfdDE)@SUM)TQAEQ0E2D4�QMVf)4QS4UQQIE1L�CE%%��PDf9QQE@�Pՙ�RTP�A0SIDQ%PUP�1M4�DEL�LBQDD@SL�9�SQ35UPED�IEQ4ED�I34��SUE��QQT13%��?~�׾k����M;x��]X(Cc8R�� ]�u�M��cP��i˨��n�hw!6��Α�w˪�K����C�������y����w��<���g�w�P����ϻ'�O�0�w�?�=�7�Xv���zvH�:9�Q.�^���Q�ތ�����-�~r�Nt���}4�v=4����r�csط���2�6{�����k�Pu[�C�c����&��>�쵽69�G��9m6��Ov-�G������WX	��n{��(xCF���v�\�9����W&t��i�]b��Ί\�9��3:�'�[������I�kW=U��9���$˗ա�)c�D/��4�����|�f	�����<R��OY��{�'�������.V�	�����Κn�^�q�~:$}�uz���3��㯹�x%\x"��K�*{@��jV��W���6�c>jM��>�|ɕ�Ru]M����۰3ܝ���T���z+��0k�����2�9��E�{�~��T����3ʫqokoۿ9�Z�x΋9pK��[�X���|�q�K}�M��*�<����Az����rڤ;TTѬ����X��֘#�V�i�e�W�]U�]���e����h|�S�i̫]��L��s�i>D,�/��z��l�f9-�Qj �*y�Go���&o��*?v���^+����}��}�<u��6������Q�յ�|{e�O�S~}71���u=u���sٵ����\g�C�8Xs�N�}/W�a�|3��Fxa�Oz�z ���2����^��,pk���zp9�{��g��-���陵8������l[<�������B����,w������w�t2/4�a��>q{�gs�N�N �݄�h\�/����}]'�9~���	��%t���nf���O%o����az�ha[ ��ٿ�ܰ��S����x�5*{�Բ�/S�����D����⯰�쯯�^w�����J6�W���:�������{~���5�{�ذ��E u�	k����]r��3Q��y��Q�;��l�vՀ���z�L3�9C���(l�ˑ�^� ���9K��Z����'l���f��m{l�א�}�U�`�6 �|�lե�u���{���ś�-��}���>�-��q��5=^Yf��ebo��6-�&� �'uF���ڕ���l�ڍݨi�ᵷ�.Z��Ⱥ�fO�`R\���mh�L�D �/y�ϰ�NS=��#�\wdOgL�;>�η�:��7�?W�|>f_O2H�x������2�g�7�Φ�����}y3��w�g�,ߦbw'^�t۬d�!s:k�'ZnU6;�y�i����c���W�)�\�Uɕ��WZ�`���������7����5��?��We��3�],�ނ1Z-ɱ]O�V��'���V_���]iq�3�e�R�7��$�ILhp=�z��s��c�a}~�9ڮ#"X�*�c��_[Ϧ���G|�a�~::�7.�v`���sѷ���ů�B��uʿ;~��7{e���8ۘ���=�.Tӆ��3_-���Ô�����LÞ��=v���t/�&}~�c ��m�ױ�Ղ���5N��Kk{y����˗�s�5�Z�{j��0�Y��X���oªO<�<�u���}:�s�����Ǿ��������az�������uvX��x�j�]�]7Ք��!:^scNe�ik�ob{�ۘ"6��}m���[>��츁���=��U�-��Q���7�ged�Ү_:�(��.ɪ;!����8l��h�Xl�ˡN��3e؝��䇱m�uuY�h�*F�-%�{������nM�w�w�x]���˘zw����>�=aY��N�^���[�����SQ��_<��4���2�f�:t��������e糼^2c�'�]v8�T{�j�|�O)ƻ�?`��M��~�szv.��h����z߳��zk�T�gӟ�],
��
vY��'S7����������
�Y4��ݦ��g��l	D!�诏9!��k���_�^{L�Ev���Q.�������/λ��	s�t���s �.�X���'����.M�;�45/d���%�Ұ;xJΚ�t꿩���,ym�ή�'��2�����&��U�
�k��_�M�%`�����]z�=z�p�}���)��_�gݣ���n>�S����p���S����WuӺ-��&�������}U��홃z#C�B8Ÿ�����.�H`z+�|��f�0�B�)]�b�wz�Ҭ���]/2oWu�M*\K���{r���³�8O<�`���p��[g�ͤ6�]Ε�=!,�}�|g��oX���2(ݞ�������6���Y	�{E|���e�F��u�@����Vc��n3�c?<�sK��_�s��S�>W�}b��Iz��<s|���F����7��u5�eM�*[tzy�|����՘2&o��>�;��6�y��~������<�Ũ�V;����Mtt�D�+:o�V ��c6�Zr���o�v�߷p9�ct�9�H���R�7]�ҏ9�.2�!S`���!ͷ-9o���{듷a��_J���֫q�"O[�Edm;]�V�o��l���'�	����a<}�7+��u6��5�/c���Y�au;Ke�Pu|k��1��A��
k���
��ŝ�M�ޭu�Y�_�v.�����c�\�q|}�ss}2ǅd[l��~���tT��_�9����.����u�wɢ�>�O`�Y���l����N�b{���2��9�4i����(�x�t�5�[�o�$��ں2�f���^��Aڎ+s�q)8���^$�)���E{�!u���=j|_�S�<S�3�7�rX��vy�A��=�۔W�g�H�7|;��y=�d�z寧���G(�or�+��Z2����z���	�>�5�H���k��=_~Λ����+=7�:\���.Ĭ���t�+ݬ����ڥ�|���eX�������9���UێK���]<�y��I·϶1��~� �81���)��<�N�G�Sy�3>�Tݙ{&mr�|#}�+�XU[[ǲӥ�_Gs�fg���!>w��)��yz{�>Rf�+m�J�V�k�]by���{e��S~}��DN僗<��)���^W�?��|�8Xy���mL�vw�=/�3���5��UY ��{^���/޾�8k�|�=��8s'��-=��	 o�U�ը%�}j����~PxVz1�V�nVh��s}�߷'1��>P7=~vr�s��y���Eo����rU�1}�p��rӗ�}9���8j��l{����qf������ߗ��X^�a>5l![ ��ne6Di���Q~�I���\�mc:�rՐ�&�u��u����C�x�U�"�&���vrKdw� �|�#f�x�o�r�O��-�{����n
γ������qɊ܇|��fW@����'{9�;)r0f��s_��������k��%�p����[^s�*�9���|t밽L����p׽�v�����seQ�8��L.sɧ6�{����t裭�Z�m�ssm�e�����w?e�8О�7�`�&vշ9��qn��]�υ�×�[���ۭ.�ۼ]ͯ�jZ}�y��ޓ7���yxws���V6�{,��B��w�`�MzȂ�������������p���s���}gn�OK�2������쬟{��!s:lΙ�y��l��:�\��9�Xoޛ�����b��`��d��+����.�zY�"�����Ӆo�{$��b�T�;'dT���讣~'Y�-�����P���I)��7����s�W]��h�r))����|�\xnh��=KΓ�[}o}���zd�4����]��v����n1`9�N�f�ߝp^۴h^ד��1�sॕ"���[m��k�j���W��	l�t�.
�M�s�9�f�����g^N}��6�%��������9<��ܒ�S���hNCy_`ڽ�!����VY�U�w�Gk+Cd�U�y�gg��<x��s���M�OuF�=�}��|>�{.�-�&�|�g�(yr�~��{=lf���41�6�=.�n2����9�n���>�y��Y���=w�{2�������*�|`\d��Ѥ������R���6��eT�~i�����Q~4.:������Uv߫�`�]{ح��T�U�_�'ϣ��=�=��G�nA�����q�������ҫV'h�}0��c�k�=f��az�_3 {ut�i���WR��6����s�q�}4�v=!����c�g�z�o]+����n�t�,%:��XO�����j���8���]FJ�+xh[1D�z������c�N�:ݥ�뫌����8�f󳝴�vۛ�>���7v'yu�D.����*r����~��H��{���O^tw[<������y�9�%������9\]^땧�\𭡊���|��q�?*����Ko3�+WJ~�g[8�u�a	����T��/�8�%�Mz;�Cq�|��ͫ�M���k<�:�.�S���i�z���tT73���C���l
�n�X�tm�nt����5)i{P;W(0��UUU������Y�J���^�?J�v5/p	%���w+vNgM.�]|���:�^��~�;�/�L㷻�fJ��E]�����KxK���7l��{[�Fݔ�\���/�`�w���܏�Tŀ�z-���;�UeK�x��l��{qo�K}��.���z��Yۛ^�۵��8�Z�~ʕ�]6���{wܥ=�ڵ�����;�s��|�ϣ���<�S����_���M������=Ϭo���0��s��m��q�v��bn�b���"U��UϟM��^K����2�˛]�2�yC�Q~�:�r�n)��;}�6�&��S%p�����zVAg#����n��t���Ÿ��ռqŞ|�^���z�pw����rӖ�ӽ�{듵��Խ�W9���'J}������u��_[��-�~r�Nt߇{�9�`m���ۗ-7�Tk8���ut:[��R�;�y �I�ۧí�S�J��oo����@�qMV;���G����왹.��<�&[�n����&Χ{5fT� �>\�n�^\��;���������]t1�����꫙�g����D��r�Ň�����Kb��-��懥��?'�jj�{��\���r�
ezi���������R����p�նa#yhX��Ξ�nLN	�k����p���b�N��9�o�r�m�s������vX?�w�{��{��&I�/�\�%�3����:��纓��ޯO�͠/OWݜ�ry�Vz�����d��:�=~Ѧeԗ&�y��ǧ��D��-}|�í��8�N��{%'�<39�L`{<�徏���O��z��t��y:]�;חX��������r���8+��^�kk�}��͊�x?+��G�ӥ�Q��U���b�-��z[���y��0cد��n�}���~9/�a}~�oMZ��ڮ��X���q������y�pӃ��t}�mzf��`������<�_��B]KGl�TG�!�ӕ,�R\�����w*NF�N�R�6�=x�/��A]�����D>�g���و5�(�P��ŚN���D�4�;�ۗ�v��GP���Sc���݃C]���X��k7s�+���Ș)���ђu���8R�S�*�Yb���t�����Դ̈́�E���l��n��R�f���io-����H�ki���m��=�e������C�6��=g�l�ٮ0��[q���4�0z���Jku�^u�w8�ݧ��t�[{��l]s��Pu*��W%�	`穥���a��q�me����X"�f=Q��ј�õ�Y���ɋ���zh�Q�D�咮�1z;�{��5�:�x�猈N�Ǐ%��(���N=e�+��3�Nm`����]�ǽ�ݎ����f�f%�s������T��{�;��x1���L��N�i�T��&G�
���)����|@��WMtl.�R�i �X3�<R�e���嗫*)kG��6���]d\�h��a��<c^9��U�1�v�N�WM[�3�Wl�Y����9hev�����N�@a��; �4�������?u��JgX6���ߣ��O�"�|7Y�h�F��遅%��
���ۗ��,���NTuj]���]�E!�ɂ���)�r;��S+h���������T�c��:2iH�;�b�V�NG�d��k���n��Xp�5S�N��GJ�WdV�S������n,S�^;�pG�^��x��;�v����OQ^M���y����N�M&ﵷ�U��)7�K8��k4f�S9�	A�۾�-�9��7��>��`�ojJr`}�[�>؅]��n#O+�� lnTV%k�Tr�e�
����R�#��R֬]�c��n *Ŵ���L.��Y��qw�U����eN;	]�Wk���,�D�t�ي�m�u�w6񫛈%�w�^<�+4n�Ⱥ���	�դR�R�Z��|u9��Sw{��-�Z���%6�f����^1�
@L�qEA����G�wf�i�� L<}/�I��*�W�������b��<d�[*�;�n!&�#���Q��9�Qt�ԕH�vz����ۂ������m�\N��ח�ڔuM'��R�<�.&��)��I��{����f�m�r�A�x%���;/:=�ԌME�e��Q}�����=N�x��[/a�����J�sS��¶x"����W�R�P�mm��v�G��@O<u%f�-K`���^�:�67ѲsЋqܸ��oU
c"�5�pzK,{٦,=xǜ�;rI�y�u-Su{O�L�ȝv�����Y���s-1�з�':�m�s�ɢ�pK7��-�r�E�k���lJ��'���.�w0�h�����r	p�-:���qM"(��g�^"�3'��U�j5��=i���oo}l66�ق*�*� �h��I"����"�����)��j���
"*����*a���`��H����J�¨����f�l�"c%�J)�(��%�k3��&&��������,�ʪ�̠*�Y�*)���)�"�(�"�"�hij�
�!�&�H���#3
ʆ���"j*,�!���21Zj!��*�"J�$����(H����)�����(����L$�"J����3���3�2H�
*���B��i�����H���
)�()��`��Z��s0���3�(�Zh�	$��?A �G�����g���;7�.0�_^�u��1�>ٝ��-'rv�X���d�O�8Du�A�Ev4y��r��D]LO�6���꯾�����<��������oE����O8=�g%�s�l�#~��u��s�y��K�d�<�e��c�Vz0�ކ���2���n����<������Nuw,���b�3�޻SƮJ��,w�ô�'/ѯ?��_^���ٍ�Z�I�E}��b}G�,'ƭ�[ ��+JPVU�^�}��Wӎu�Y��y�q�&���rz՝���k���[�%q�Р�UMG�r��i&�f��t��9��sl�݋�?�vc�E�y�j��֋�I�^��ԭ�����I7`�gm_��~�_9غģδ���޼��w�>�Sc{�6倄w˼>O��7=��.{��>��/v���l��m���L�uH���lQ�_��3�5=y]c���E]j��ֵK{l�fy��s�~���޸����.`���`N��?�ï�<��R�wFa>8�tn��2��bW���L�fe:���;�
��˽o��`������j���>�+��&��l��z��yK8�R(ʽ��XHjʑgY������ki�S�t��c����<����F���Y��9z���R(��}�}_}�u��&o/L���fc߫�_�\��;xJ�t�Nu'���k0��ꮂ�����*9�>N��#�"����nV\��Z�e��V��܁ӹީ��ɻ<�V�O��~؎��RSE�r�y��$�5��u�{���w4�.��SUY}�^�������bØ������]=�����1۳;��A5�K_8�ϓ�>�-�O�s����q��w�U��w?on;�.jSY���V����|��~��}Q��j���k���ٱ��ӯ�\��M�N��OlN��s�vfQ�/=��Kꑓy����d�]��o�k��'��+={y���/�uxG�Ǹ�9�^�0UC�acv�V�p�<t�=���!/�4���
d8�S���t���ơ��!�Q�%S�u��f��owAa)x��M_S$��-��iEb)�L.[��gZ%��Ej7۳8b{�s�r�#��N��TLX���R���ڔ�{ķ���SDY'���]�¶Bm[B�Ҳ�Xem���tz�V��i�[oy=�Qonp���(�.�G��Cp�Y=sy�����G:-GxT�(@w�Iu�!��5k�9��].�ȣ��I���W�}_#ɹ
�����D�OW�)՗����T^���7��A�j��zmd��^�hm��q��<��M�-�>��c�Qi(��`%�L�\^�i��OȹP��֌˘h�]��M��7}���͘7���֬>���wh�%�L�P���_Zer����t֋.^k�j��s8EꗌV{Ӓ�痢�,�L�	^$�,�y�I������-R^ȫZ�T�=��­�h�G�P��W�A�EB�`��.�=��ϥ�\8'�#])rG/���zy��ѢG�d���g��]Y�C蠗����iq^��%�\2;���qے���I��G����I�ᬱc�[`Ͻ�t��B��[�H�eY��~ӓ̽}�h�y�0o��i&l0���Dĸm2�.7���hYހ<���t���^��}�ai�DϽ&����]�r���l�M��_˗��OƝ�\z�^�]�4'��os�.���4����(���D��I��Ezfࣃ�}a�j�D�_���W_Ws��)�
טR��Q�Mpb���am��U��wӨ��赗]Ż��oCj���t�EsA�� �'��
�Fp�^��8ºƛ�]�=������΃S��)ϱ�(��>�lQ�`ŵ��\�t�¶��*�*+�%��waޑ������qt�M}�yX?b��)|�)E�@t��������t�踣�{=td�Uឦ9?=����}�N�!��۶�%3kM�۶�ivݎk9�7ҡh�o�<$/��E��,iz��%����y���E.�%�a��<����"v>0����ʱйoW�'����_�9R�;��^�X���t��H�3����w�X;AUa�$=����v?��:潵��Q�=�����s��8��`�<0Bଵ�Z�A������T6e���tҰz�)�=���w���%�G��j;a���g�q�r�z�� ��f�\.P�`��$T㕞̨��X�+ʌ���W/���3���_����}2��^��L��(��K4M|�����0̴�t{��8�1��o�(!���C���yF�Ƀڡ��~�1B.���P9���t�-�wu���қ��u���T�^.$#�Ƅ��:mbu�x;����Vr���18&Tō�}�}�J�Lk�6{X����Z�G��J��]��@����pO��3�q��	p��N���z�;��,q�r�ɰAj�(�����|jy%��V��߆{�c��y��2_���t�{=J��nt*�4��������ө�ֶ'|��'A(�n�4��u��81�^=;����殁,FnՑ�D"yͺ׉�����5��k��<�i����i+���I��pZI����V�q�U�:3��
YJ��E��bn?y�b8z}���r1O�ϔ0�TD.�Bx�V)v�s��x[�<Yv��LS���/�={�/i'<�zd��i�8)�Y��d��88����z�g�i$��r٤�1�z����({vf�^�4ֹ�Vk��{-�>Lt�t����8��׹ ��Í]Gº�-�C������`yL��C8f����i��K��N���J�A���k���B�8�[z�[$����h��T����R�˦^m[F�ZdE���$�#�<�2�ՒǙ�;��z>}6f�G�-õ�gqm+��q`&G�ԋ��e�=�Ę��z���|���\��w,��Z^���P�Gq�\P��s}GL��im�'C��A�+e@^�e����RV�<5�gsga�>v8��r��C���=�p���-���u?s����+�����Ny���:��F&�縋7�s�����z�6���U�|0�0����=�E
�L�Sr�rf�\Ճu�e����1b�]j�'�8a�ZRl��Nj��N:r8���̕i)Ϯg\��С�����Rr�wz�3�O�������ˋ���
뙛/ ��W=Ee�]�P���M<��.c�����3��~ >�o�uS�]V���US=�TDJq\C�yy���۳����A�����R;�J�ܛY�����7��t�D��g��	�c�x*�b;sj��?i�O_5�]�r����.���rs��k�}�C�H��KA��p�J�8��8�U�Gy���]��)�Pd��	�y�3���wZ���fq�}=o<�Ά�+�5��L�O�����8�����[x;��,f��7^�mfx�����0֣.����p� ��r8G�uʦ봋C�Wnw���Uӻ�Z�t�(؎� �"�|����B�/3>M#E�؄#�ѝ�Hq���gk.�z�L�oh�oK�IP�I��q�p��'MŖ��k;����z��:�Ͷ��>�@����ܪk���pm�g�}�抽pXRP`�r��K'{3�������p�hY�e���֍�M@^G�K�J�7�-3�}��}�4��0�"�VE���sS�o�V��Jns{�õ<�iJ�fτ��7�*ѐ�,U��R���喱\�O�l[�Z����gGwoQY���U�@j�c�M�EMoU��޷	k,W�.�s�ť�����d1U���n�׽τX+[}��>ݒ����f���=|�-a�,� �N{q=׽l�κ�f�Epkȹ+�v7j�l,�V�{����}�پ:��{����7�NVt����7Tk�xt���ݼ�K�(yw�a��ܭnsY'A{��+o����r�n��N�->.'�{�}��>�lI�[Wk�G����e��'�Ƥ�}�GR��B�P��ΣI���s2.��x�:��!�@���{��˥��/�x��y"��Ui��P�,��	6;ԋec�Q_�NB`.[��8�:����.�o�\��K���{�1��@�ID�%ʋEqn��yUFޚ�>�]���0u����۬��u��L��u<lTSKA���3�U��Ӵ�T��\�F��&��H"W~�=QgGu��w�M�3{<s·Z}�G�ݠEF�IsS>�C����̩�[w���s������jڟ)��^ʽ"Ny�fJx��q�%x��4M}Α&�_xw]T]En�p*�M�A�Jq�-g-�zT>lJ�j�P�Y��1vL�l��P�<i�5 F>�k���N}~V�^"R��ӹƃ���u{�g�1/&P�ߜ�kF ���2��t틳�Vb5�c4%2o�uѼ�¯7��(��{Ge�]O����X�ϻ^v�m/P2�b�vZ��]��|����]�$o$M�TW�*>4mM�ӎt�w�2��V�}β���WΗv����*�/GS��G���8�&ub�������4z.�)��?%d�ĉ�U��VO�;�΍Ne��	.��WF�}����o�O������H���_���<��P�	�(����,+k��7���hGs�5�e�ggk����&i��,(@�Q���{o*��lٮ�����r��:���9~���V�)�u�{�\�{�`N-+e@Q��"��Y9���J��%!6ź�^(O	=�cJ��5Oi�Sv�+��ݿ!n�3X�kD�rǢ��鿞�i`�l�h^4?��A���q�.C[���t�$:����-<��:���n�9�!�۱�e9�7ҡidu��ӵe��
�C������ٳ�8����d2�r�g�>��Ƿ�pm�39x�rޯ���#K/�hwq﷽=���Y��꨽�Eo�Z��Ey#�QJ�)�W��G�S��y�ŏ֑���)�}r�R�\T �jk�p��t�Zh3du'R�����t�u�������gw��l����5�.�i����q�r�޺=�6��΅��� V�+u���ݷ���5V����8��4MV�ya`��������%	���7!��G3Up;vE��V`X����1U�t:��>�f�}��mޤ�TŹ�������_��� �u%�]s�>��N�xEC�|x���/��ݒ�;s3A� >��a����ٌw�^���(g��،7=�,����y�L��(���A�\�����=�o�6��4`A;am �S��ϗSi��ڡ�=�7���cm0櫅�����^�{5�wG�^�g��D�
�-�#�ƃ�:z�P�uI~�8�Y��z�!di�{�{�U:�[e���O�۪u�Xy=hiI5���=~�KܮKN��{�yl�yP22f�=��M�3��o�ghOE�^6(O?ZHk+�Mq�U�Vjg;h�R��|�o���o1��nz���"�h�pS�p;r��o�Мb��m����{M�+3���.�r�o���oO�wW�7�
W��H���Z`��
z�J'��fM�4u�jZ��
ٞ{�'g^�l.��qhI�x�j�k7ʬ�pPS�0�g˥���{��H�zܢ���Q�:��s�E��m8T9�eCy�p�f����i5�cs�cK�z.JĖ�/oxʣ���Z�~�x����>��f���ט���AS�о,�"5Նt�dy�{CH|�5�5V�5��]���e����w4T�;� ]�uo���a{7}Ţ@�ǵˎ�Ɔ�Y�*�v*�Z��Ϫj�-�����e�)_sg2�}8����Ǒ�6�\��M�'��$K��:m��{�I$����+47��諸v�{ݘߪ��'ݑ��o�õ�ck}[K"�."���x����T�����X���t���Uѫ~7*va��=C=�չ*�=�|vq�՟R�B��ZZ��W6���''e���:��,a�t�r��:�<s�oWh�p��ؖ3��f��U�i�M�g�bBȕ�Cl��Y�Zk�qC�P�r��N4=ӳe׍3s��n&�?)�k�jd|��a^.$�/@��9'�xr)��l��<�,���{Ӎ�~iwoPs�'�b��[num��c\:z�Eau#��\dHf�/*�b�9��"e����Nv���	���ޓ�5捺�ؠ,�V'R"X�h�KA<�{B��2�R���.[:p�M��mUz`o׎;����V|d���~���H�`�kR��s]��3��TJ���u��/t��nUV/(#��%fx�*Z�5���}�����$���ZR..���<�2�nw����t�Jc4��K\���`�b:ȃ�������%vļ�0����J�n˨v�
�flN�k��Gx�|]e�6�6���nwZW�S�<���Sx��3���V�3��fkG�����:����8`%�?	-��L+u��2�7ˁ���0|�ٔ���p�I�t.�i�=�rg�Qn�t���m��WR��Ly��Θ8H���q���疌&���=]��l�<ʹ�Gk��\ay��C+T�dy�w9��
�vǖ��vj`܂�يSF�{��U{�����)ͥ���{�a�.>WVK��々7Ho#�W⮩�	�+=�Fg��;����t����v_#HO���g����3�o}��i�XFvka�Ã�Wre����l��#��u����@�B7-�Pe�t��B�$ӳ/EO0n*z���pǹ	�}Y}9�m�}&�TP�Hm
lRoE����'O^'�Qƨ�������J�;�
��Mo����I��;.��,�ժ���]>�3��m�m���.��޹�VZ�jq�G��!�Ջ��Iju�{V=�g(�6��m�7�E��?H���c��>�U�����Ԇ�;��5}^�����;]OC1ܫ�d����T��A6���7�Ew�
Ћ�����:H^�Kd��&�=��;�݈J11��@4y�wϖ���B�>�ST� ̾�5<H�f�H�E������*5s��]���o��շ�}���Ƒ�?@ev���0C�>�@0B�e3:���q��w"�$˭ �V���g���*��Ut�d��,jwWP�F4�oS]!���(n�Jt�)���)X��>7���QJ��=���C���N�#u�ڲ\���^\yw����)�|Vs��L�<*)ۂJh��ɽ[wK��P�E3x�r����D� z��k�%3��oe�y®��sF��K�h�Ju����_��Y��S;"C��Ʊ:�f���aVV^.n�S��F���y�E03�XJԇ7{���قk������/;7lF�z{�ewzu���b��Z��2>koˤ���ݹ��5W�n�|�� f��sCᘹd��gx �K2�Mmm�I鶨�P�2�P%E��_*c厏Z3Xur�5�}3�G~�i������#S��iY�X��|pm\�L�u������u�i��;Ei]Mk8�#����O.�@�V���(�wG"	������9c:�EO1�Kх���nnr>�zr�w1���8l�f�����L^D����|ؠu�6�i|���!'��$����9VR��w*V���f���mZŵo�k3-j�*�u��l��$�«�j:���<u{��w(��[�n�1����oWw�J��ZQ��_*��{�8һ�e�m���۾�W=��������Z�7��ol��
�k�ױ�<U�{�VQ�R�p�|�]���oT}����>��H�fǒ�D��S�dEf�Ue��@����1��
�
&��2Z&
fjf�*�"��2
X�����#�0��""20���j�*&�(��%� �2\���32�
k#,̠��+$��*s3*�*�21��"�(������̚h�+## Ȳ�,��"����*',�r���(��ʬ���2p�	��	�¬̜��30�r"�,2Ȥ̌��������,��r
�rr�l̫̆1��,�'�'&�&(�02��3
��,���(,�lĦ2��h(i2ɣ2��0�
30��"�j��#" �j�22k*�	�r�ʓ*#,,���0Jʊ2(j�,Ĉ����h���M~Ӳ��7)����&��݅f��*��3F��O=�1��>�p�/s�>n��x��� �i=��ޤ`���	�F��M)ir�-3�����b��0RW%B�l�-p�,���ԝ=^��!~��c�,y+(� S8l7)�	�pm�|1�	Y�h��R��쮡�����P����<�\u�<O��4�m�Į�l�j�<�\����O����cބ�Q.�����M����}[2 ++ݹ����g�e\jה8���ʖ8ᦼG�H�>�'u.��Ӌ�.�rs��U�����8����5y�6}�*y�p�+��O��x��%"���{�*۝��tEz����bc7-���b���z���#|���^�>�9�jϬMvu���.�y�^�^���J�� >�Z�)��N]ë��^1�u�&B7<W���Sl۝Οs/��R��i��\[,���I��ԋec�QC9	�-��en����{����Mx�(_�����-�r��\[.�Ϫ�H��M�Ήb�fb��)�2���Ѵ�r�k!�%��zxR�𕴑c�BӔӣ1��l�7���&���{-��*�^��STB4�W.oT����m�c�́�Oa{H�DW�bAxs���f�}�s�(b zquZ)��� ��������ќ��yȝq|�U�ho����;�7]6�-U(��n6�psќUYזV���*��x�:�'z�=��t����Ꝅw��0J�k���Ͻt{>wh_F�IsS(P�W���5�p��[}�#��=j�;G��עU�s�����zz���I��&��H��^y��|��hǏ�+��(>V3�k9n�].{*��8P�-��.�	��$Pf{{ݓ��>��S�|KKEj,WS��:�zu]��Y/&�ƜQ�����{:vi{��-��~���Q��c^VI��DG~�\��p�TX��-�0J�։uC�>�a�=�=�۽N�Oa�O�����
T=��������%0����nݳf�t��F}���ӱi�^�*�M�=����]���J��h�pS$�D�V+r� ��V�<|5���N��+�%d�6��e�����|�ZU�wF���p�M�=`S^׵cb+��a;ܥ���3|�5o�g�T�S�(�_E�!�_�5�a춖M�{�>:{�qG���3�� Uީ��.{��V'��۾��sn�9�!�v9��3�J��c#�{��B,��"�����o�c�ܱ�J&�խ'1����`|�ʁ�7>��fN�{��|36�:"�S9�d�a�wQ1OF��M��va�,S�}cE"w#$�ບ�S�^��v/{|���ݶ��jf������|����U��z���Q���EfuG�~ɳOyr���债��OW�D�z< ��5��t��7��4x�{g��|k׾�!"z�=/�S˯-2+��z�ʗ�X�`����G��,�f�dC����\y��v��]I�<'���xê�rM~�(l����"����oa����Ԕ�+��N�e�X��c>����l��mD��Y䕒�q���K���H�g��Lʛo8���Y��،7=�,�[�\�^}��9��`ZrG}�)b�����(��W#��A]��%�R���m=Z{T7=�7��B2���U�j(د;,�n���ۍw�����\���cYA2*��v:�M�	�3]o��zpҳ�[���;�����o�"↰{�ޟ^��?�a�8������S~f������f�G@��[�A���M�h�������tj�V ~�����%b�q���v��㱮>HnG��w��q{ۭ�V^J��p'�t;r�ȇ�4%��H�[qzm�Tz/8����Voâ�fT�~U�2���z�^q=�$�Wi�x+�iןvz���)
2��e�WXl�|�zz�{���M�;�w�J�V�Lo�.��-�A6��7�1�=�	tX���:1���Vс˶6'V_=!Fb�7Q�9L7%g�����+��2�Â���,���+0�G�����ܞJ�q��os�)��g��yP�d����v!�oK�k�¿��0a�ϖ��t��vޅ��Dm������͡LS�Bu@��,yL��C;6���H���s.f�������^��t�q�Թ�'�P��+��>�����>���޺'�c�
�b�Ȧ�E�rKizb,Wz;p��G1򸽫��ܴ����D�Z�Uw"�TX0uW�.����H���ҟL�3)�þ���3�Gq�nJ���j�Ǡ6��/gǮ��藉���s}�^��_<K�^��-06�2�;��]~�Ck�g3���{{�A��c������C��G��[m�U-��qBɘ�gQi�ql:�.W4���w��9χ
�a,�ɷp/V����=�g��I�>*i%�m��*�|��j�(�<���..k�=��WfE�Ӷ��:0����K���#��+��>�����C�Μ�p�i��-~���<K�!(����N���k�o�GYLi�����w3��޺,��mJV8.)Sj��-�2ۆ�;��עͧ+J��a�;qM���jw�6��L�qV����Hx��[�[�3q�ÆH'�g�*��-#h�U��K�u�h'+�Y�7أO�L�7�gx�*�x�W:����4����fnSJ^���.��T��|�\;T�ˡ^��f��Xt�?<�9��x�<���Ь%�;�gʗ��æ����z�QYϱa>��xa��e>U^��"�~���pL�w%�	g 8I]m"n���}ry�u�|�+��ՙ]|��2��0�Ü�F5q�+���8*��;r�txg�]��FNY7�vzu-��H��4��C�4ǞNI�*��9o|9��o�tyh���=W�c�6ge�>��@�a�c��F�M@T��ܪk������P�p�t��(-W5?eGmoYؤ^Q>�����U�z-���>ߥ��k����_��M<�!����y������-�w�/˦�qL��ne�����yدe,P�9�jP�+k�|�L���Ǡ��;R�Pc�,f��Vt�����ln�}i�5�@����v���v�G��I��Ok}Ճ��"�]�s��b�>ܶbu-x�x�y{��b���I$r�2�(k�j�:�>�91t�?t��-�.z�k�	t\�(K��F�˿qG�[}��F_5!����r�~�H7WF��:�i4���cN���-}�&��})�Ҍ��� T�p�1r��:o�w�Z'���1����<w���TO3G;R'�4L����c=ѩX�(U���E��S!�b�̇˥�^1�uﳍt������[�u�#<�p>�Y��$�z|��_S���}H�V|��P�Bk`�~�Y�:����6�r�:�u�2P�
�Z'Rؽ�uYh�/n]��Q�l����.}x-�uz��H6�6�D�ǽ�y(Nu��Ʒ���m�8H4-9�ڂ1�Ll�ш]��l#����I��j'�����FOm��f�x�C�p����g��(F�A.j96s�V{Ƈ;�k�c���q��~Y�r��x��N~�OK�Y�=l�׭ <=���?������<;#���$I�ap�7��q��r�-\�z%_���"��;���Z~���\���&zz��Ԑ��	d��P��ý������;KɁ�Ev4�����gNi���O2o���i���u�eW����D��Dm���RipЅ�T�tm'2��}�6%���f�jg�f%����葠�r���v&���6�~J.9���6k�L��͇����V�r��-��'.fq/�1������~�~6�иe6Ҹހ"�f�$J�;7�:�u���:w[�a�B��)�nYM����{Պ6yxt�,��S�#�/�����2���-g͕��"z��~�b�:KB]�A=��oL�4�,�	�h`�ӓ��1�ޝ�S���i��.�;҉����]���p�G/��?r���<;Ӻ�^)�o�l�qW�Z��ү�wFǜx�1=FV��J�2Rl[���_���[��=w���/t���:�e]�;���_E���P6�igޛl�mC��'7��j݊��=����9E��밡�p�<����p�V��m���s0o��'��B���^o_b~[;�>�g!��y�:͌Å�c�\�S�	������pm�2��=aǧI�ݮ���2��I�ʯ�eW����[l���^��+r�5}N$]P]m[�wr������e� �l�	��=�u&��ӍMu��U��<��f�I��΢�M����L�l(�����s��=�U�y��};��4�\��'�,�t{�,�\k��l�V˧��r����>H��[T'�;��晛�;����m���	�b�o����W�7��g	�I�0 �y �*_yb��y�B3��;^��~����m�v~�w..�ӑb��q%��{+�Ҏ��E�0�䔒�h��Y}�/W7Y^ڱ��e&�uz����cj���pE75�j]#�<~{�N4.��;]N�꼎�G�UG}G��x�e�Ɤ}�uo�����V{{[�TB��hf^R�ɒ����R����4ļ/[�څb���l�H)rWT�k(&E�A�P鵟'P�u�K��{��9o�2�&�s�������WbreLY/����@�H�^��B��=`z�.�/�����"J��&oCSn��{�G�חxEv�{�����P��X�)$=��\�k���v�Ö%�ȹ��&�.��v�{eёY���h�pS�p(a��ȇ>~&�����ց�I�77_���|%�Y����U-x�_I\F`�x)_�H��I���ORϺY;aLVa�C٦	n�~�+_>g�E�#���f�%�^���C�w�బy�`��agUo�45�^�û5�ی���B*=B`�g���7��}�{��x��������{no����Uޓ�R�J�ϩ�M���<>q-�r��k�LO���x� O&��!�֞k�#U�n���Te=·<S3�B���猫0Vgǅ#�����;JR��>�ٹno��p浥7-��S��c���N��Pd�_z�����Z.��4:o�q!��zpy#�n�c�﯆-�f�&�d���
��tY*�^��S-oMbL���wgUŢ���^'2�f{��h	]S�F�]�ڵP�U�N��}"��2���xWE��.�u�Rb�d����7�^<���g'%əF��@�&���_����_jB��C��Sn��L��l3.��P�Ա�zޮ߲\;�����U���7̽�J�ϝ����mr(2=PP��J��a�"͂�T8��kӍuD0���C/�}=��d�R����xȒ\c������\C�yv�0�yt�t�+O� [�������g���v+*�-N��`�.,��f\��D�a���}�Y���f��D�Λ^�Ս�������9��潋�j�R"JF����up�p���oǥ	��}�K����ۛ�����z%ޛkya����8短� A�֥t��P]W)׺�]8�N~�B��Z�7��˜���fx��������.�~�Y�p�0S�/�W�\{w/�Am����KyK�v;��i�{җ,�s:ȃ����p*::P�Eqʏz��^Q��=��6x�V�g������;.�Zg�{7<_��Ř7�
J�B�&c���g�?w/.�ڗ�0ʎ�C�Y��VQ� V8M+r�_ً4A��O��D��z�ʱ�F�q�	i��u�˸Z��F��_��\��v���v�u%�dCp��M����œl�\�Q�ja��-����Q��P�|Q��F����8x���i�H�>�Ӗ�AW�WuV���s��#G��a�6���m�1[n�I��9I�k(��GX֥�ҏ+���/�9�E�x�1�;^��W���{y��w;���#%2��%_��H��[ҽ�J�Y�Mx+7ּ�`�R����m^%ݹ�ռ������I�~ڳ�p�؟�gK���<���[yv��8sG��Ӿ�Yi�)��g_5^��h5Xd_U@|�A�rٙ�;���������#}r�wP�p�{�[9�?{c*l}o{��՟`������J��(_ ���Z�)��NfC�[��G@�u׻�_�s��l���������Y�I`|I:=�Y4/�lw�����Vki�\���;��]T�C�oW��i�k��JP-�l^�����qu*�J4��:��n�k��wj��B�G�X9z*��קZ>�kyd~VDq%���[EqaVYطm�-�ry^�c֮#�}��IW����&�%zf��V���\١Hpu�޷�]o���m�o�l({�/�C��<����zE�9��}=.yd�f�z���|���=�m�G�ᷯ��lN]a �����iǻ��T}{P�3¶5��Z�������$Ǐ-�x����bW�)O-�ڪ�%�a{�0Amz�ߟJ�%���_[8��(I{|��Ȼ�x���a���~W��p�4j�S+��@���a�a�W���y{�1�ox�+���W�]M�J~�uJ���}����|�Y+�r��q��8������k���8��Ã)V�����v4��Oy�m��9x���f.5^�V&�T�檸�s�3��$r���:!�0r��N�؞�������}�+s��(��d�g+>�.��o#�����;�L�aDOo��C�� �������a�q�6�?(X�Z�-�0]��eq�ʺ0���MIݙ�ҡ<{.��hl��|2=�VG��+��+���ة�#y��;�.�zb�W��Z:��rU3>̵� ]7MD�a��YNy��<�z��Y���u����`�*�y��kM]�%�=ǯb`���[d��xU����}��o=H�W��Y��>OLs�Z���f?�J㘔ƹ�ٝ�E&n�Ԫ]W#,�L�.S��}��g�<;�W�+��grj��� �8MkM"�%��<���R���^���vє<�|&{ؽJ�u`w�z����t�%ͬh��B�$T6�ٮWx�;{{U3Qv�s�)#})�kǛ�u_1�xL�aj�(��C�����ٺ��u@Ҷ8��Ͻ��>�GK��% Z�@���7�=�L��z/_�������*��s�.�no��oK�_F^��5�	��GmA���<�>��>��İ��ُOz���>n?{g���8ƐM�7W�e���M$Woٷ�m��a�7��x]&��IS�c8#�6rhu3�Fo�W���!�{�؃��`>��$bO�j����l�On��X�@�u�]�@��.���������l��q<-��>�++d/&�{mȟr��ZG4Ԯ���Ԫ�=����q��:M�'m��Kgv�������b{���=S�@��K��BӃ:��e� 
hAРF#H�$c�k�S�����4׈]�>YZx+m��uk���¥�K�)�M�q�(�������>hj�J���p�T|�Z��V���# ����9�@m�Z��̲��E9�F���N�A��e(c#U'o���J��R�5���[���	���-�x����v��}��kR1�f)s��F�{y�p�u=�OC���ZD�B�Ĥg$X�r�.3�n�	u���כA��������\
Ѷ�I����e����R�O��7����C�Kq�,��L{{�	?�Z�,���r%��Θ���CIn<H������=�1-�|{��D�-c��Y���*�'.��wQ#�Y":^�6 Tb�a���2[�\��,m^9|��.:��;c3Q��^��y�u��E�\��� ��$�3���F��%�
23#3�
*2���L��r*',���c�(��(�"�$���"i('#*�(,0L�)�,��,d��	��"�sr�3*"�,����)��0Ĭ�,�����(r�0ª����L���L�� �²""(�(2�0�h�
2r�),��&$�p�(�`�3,��I����0p�2�L�*��3,rr3�3
��*�"'
Ɯj3�0�2i�,��)(��0�+,�,"��"����!� ��!ʂ��,�1
�$����1+$��*�ʌ��
[1
L���ʌ�C'2���̃&"shƤ���+#)r2C3
�����"Ḅ"�	��)��0��J"�*��K3,��2'$��b�ʖ�,,��׾{t{���<��K���!\��X�:et��r��]:
�!t�M��hÉsv�.�{#GV�;�=�*�RO=�\��8��n�e�M"O���(8���A��[��p늳�7՟ISe�l�꽋A��x�cfI��m������y"�Y�$��^!���ý���� Ϣb^Lj�;��RܿN]&�.�A�c�u������$��#�YR��I�����Όio[P�d1��g_��Zn����+�|�F�a�>V���p���;J��\	����ݍ�U=�	�w�5��ð��h��g�����L���sׂ���� �-��놖�S�˛��v�4�/:���.���ye��tZV����q�9񘞥�,�C�7��/Y�^̗8��>f�l���[�4�7\�g�r:����~�'W�p�'[é���T9��ܴp��W�-�ҵ^)/%�/�Ǟ��m��יS��fRI��J_���%�]V�i>�=������cg/�IX�b债��T�{�_- <s�/�X2�[�w�H����>���z�q<7^�=o�,?p������Qut��ai�;���l{�$����@(,\�򱢹XØ}y�^�����姛DS�s��	�6:7����~W���}ϨR(���� B��}��;"{�%Y��X�x_aI_�p�< ��t���G�/'p�W��릝G�c`Rǁ�1l&6���B�-Ǉ/�8�#���Ϧ�"ӝ�{��M��8��^xù�e�B��A��'�_��J�O�|]7�ى��.�7�Q+b����FOP��o����E�&�لp�|4W���n�w�vNm���!ϒ"r�n�vS�J��L͝h���+{���[�]��7Z�r��:3��yGL�DНK��>!���A�]�˩����sǥx��\�=Ji&�����3�7C��C��NR䮩��PL��4��E�g�v�������7\�L�o����Vr𞩈Yɕ1d���hs�y+�uP���/��t��K�gi؆��Aַ���X���｛�"�Wl��2��eB,J�bc���k5�X�\e��<�Cf�+*<����W�+9qϢ����wFd�0����q�O����n]���4"�j�-�x�����M��MO���K˾,��ͿE�;�����ڲ�=�b�fP��/��҉Rםȳп\�k���?u��,�D��^S63%�^��ޖ5,�\��`z�C�5�'lD�'�m�`֯h&��B�~�VgHN���S�&d�7
[ER��I��t�x�3��j=�� U��:l8in>�z⫸C�N�9�a��hW+A��sE�T/U�1�=9w]�.{��nh�r�gA��}���T��B��P_��9֡���,��\&%���P�6B��>�|j��w�i�N��4<q�p�Ux����^�&Z�x|�+��ǧ��g5SFB�,�fu,�]{ztڽ;�d��%��wC���\^��E�Xߚ�g|W�`���U� y�R��N���u�yJ{j�=�4��2��;���gގ��ђ�}S�G�g�]������9����^��ٯt���EoS8&Z{a��NP�u,x���fg��} �l�վ�y��O\���}E8�ureA��%���M�=�Y�\� N_5��Pe�U`���{��©<�/
��!0�@����3.�����X��j��1q�F�<��{�q��������z���r�˵�Ӥx_�qqe��T^��������r�[9�����w!=U�91��=|ױ])�$�@�&��y2��3u�X�ʥ�mwl�#����^�mx����^�e&���B]K�<�չ����4�,���*��qJ-���k�ޫ�ܻq��W���/]�o�w�uw�A@gK��z�a���xCA�:�����Lf7�\%�����O��	TW�)�f�l�+}Ȇ�pG\샄/��~��k7��//C�������TDK�/�;���|��;z�Ju;:u�e~��+�O��a�~�����������.�%�	d�Ӎ���S�T®��X����DԡHƺ��NW�4͎�������F㬈?Ev�8e��x+�����g8��u��6ŏW�"+Ek$xg��g�����1f邒�Bx��9�y���zl�V�X[[�f��d�N��-C�Լ� V��4���U��DT|r��ѻ���v�k���Y�((#�����V�.��"	��Z��.�*�*�7�]\�.dy��Mޞ�y���|:��c\�U��$�e�+�+yg~�g/�:��W5�KE~#ZQ�	���}0���JV�B�h�/J��;������^yM��&�>U�U<v� 7�Vv���u����������V2�"���8��fw��bҾ����g�5�ĠZ�<�s~s��9�c�Q��c}Wkm߃'}F��3��}L��s2���.U�J7QyBVbG�x�>�g�)z3FTvp����$�z}O��x ��DwK�Yp�+���kU�u�RP�挾���=t@�y�-��)4�*���X��힜���^>{�w�ЛZ룸A&�wt�76��R�-(L��9ް�>~��J�H)k�����ȹ^AG�o�_u��)=�ɾ��yyT�.�Z�)��`�ݹ�R.��;�̯�3�x�B`��u-���e�*���e�Jᾼ{g�3��}���H���~Y�D���/�	μ}8���Qh$��l%�J�ZV���r{!u��)g�]k���*��֌�=��̽�Í��}�Ω��{�>���x�	cS
��}j�b.T>��7���}=.yd�f��]ԐF����^��wn2N�h���?B��!A�yƃ��������g�o�^�':k�6��\����ȼH��r�4z�T:'�#C�.J�S#�|��4o��W�K��z�}�_�B!�k0�avn��-f��r�pGF֌�����RK�#a����N���Ŏ��?{��絖�/����y�����V�B�`�H�l9G��sقy���	�_�yh�LK��rku�w�w��ǡ{� �S�tU�J����L����yf���aF����~9[��0��B�k_:���\}�V�߳h[U喦��iZ���ǈᘞ��,�}7q*M�)R�(vf
����i��t�)��!�Ю�O�W��p��&��߁����w�M����������s���)���!���8�|-o��"��P�[lO#,U��{ݪ�*1��]v�*�a�L����<�{&K�v��c_�ގ��?}��s'!x��/��<i�1��)��z�#����,�n�i�A;�/x�m�%��R�W��2�u�FRՖ=������P�ͨ�]ig�v9����v�A}wӥf�u�n��bW�Gp�-Ƿǽ���M�g>\�9����x��BzP�mL��1�D�w�� ��h�����z�"'��OK�޷�XdW��^��*=����F��-�=�{3t�^� �ԉdۄX	��<]I�<&���x���Q=4�8p�|�
�/la�^�׼drD��t���ᕽp�S:��:-}�7�/�5M9��	w��s/_�bj�a��˽=�v�T�Gy"9����y�|��晛�;��S��m�v�bI�����sތ�H;{r��K4M9K��Wl �au��dGL��̺��v��}(-�i'��s^��Z}�[���ji��9��@��R��cYA2*��w�:mMO���һ�{���)��H���={
�Yɕ1d�� |9�<�Ө]���߻��i�/���A�:����f.H5	�/n6zU�o��e�t�]ݐ����w�}EYޛj�p��C]4�����D1T;��g
������]#�i�f���,�ve�� ����<M�e���x�Q�=&��Vz�ҙ�2�\�O5��p)h��:+N�߽X�� Ƚ���j��Z�pL�E��b`~���f�&_1��Ǹ�]����kݝ�!o������D�9�����+/�U�K�=G���wdC�I�a8�7��̜
�V�s��x:���ouh�+7�"����DJL��OR?f��R�l�Ew퍞���=<5٨m���V����=y嶇}�,jY��,&�㾔�׹p�`S�E�7�*ڡ�tpg݀ ��lBP���Co�xK2��puS����P�xpY�hP���=둪ZD��������^0�^(1�?)�7����ߓ<z���4h��r���[NU�;���e����8	.��wC �s-+y`�ܴ��V�ȼ."�e��5C���w���d����R�|�d�0ڤK�2��;��=C���7���g���2==�M���]���Ǜ ���G��ց�"B7��p�
e����w9C�RǎM�z��k!y�l'�Y2:ٰw_Q�t���/V�x*E�:�1*�Ri���"͂�T1^]ݗ3�q�}P���wH�_q�7%��r	v���> {F5�1��A���g���'�dy�b����9�،�����O: ���}�b��*��R��d��<W�w�۱��������MV�-ǹܲc�S2��y�ՠ����?t��/���.���.Z����+��>��3>��:�S���8��U�oi�W:���ya��/�>�wF%��������d�\�H��+��(.ʭ���QɵÖ��n�~�y{׵|hr���c��91���qZP��7��DK�C�KA���}��ǯ+�s麕3����h�0�ꭸ)3���ٚl5���������a�K�#�fq�`G��P]5_��6��;IJ^je
��SJ��僜��ҳ<{���`U�ᐍ�۞/���V�q�����uk�p�p�:ZU�K����i�o�-r���0Q�dA�T�������+����{T©h��a�{7tx.��T8V���jS<5�W2X��u���$֡�VjTf8��q}��׊�W�|�k�9d鸲�/�7����a��Mۃ]��t�W��雹��Ն}9�%�
d��q[^K�C=�?-��r���Yg��y=�~J@��^�^�����aVz�O��y��i��a+Ρ$k�oJ��[�>�`�Z�ȬR��8�	��M�v�)�zI�2a�R��)�8;Iج,��m��>X�8�_�WY��ߓ���w@ܖK�쯝�.�����E�|��ոc7ҿK����'���M�zr�Y�{!�/�ǌ�;YO9�{���Y:�Ӏ�d��9���{�l���k��R,=�����ˊ���x�M���^;J�v�f��ڑΧ��|8������b�5nXdW��l �ؠϷ-���b���ϫ��G	'Gf.�;y�4)[�.�n,��=I[>'�	��T�z��9�Z�2A'�x16��V�W.zbn��_�L�j�Vs�����k@��3>�d�(I۾�z/ڤq����siR9eO:\���L�z�'gZ񞊽>J�0��:P�Eh�r����9���z����'j�!;	��Ӱ�ݏp\��^>�o(�P}�8�I��-hp�\u�{���;�=UfЖ��;�O�>N\#ө3צ�7��<�֯�޺<�����px<�Ҥ�Z@�"A/j��uԙu�<�.�x>~�b�ޜ�����:h1��9�<�-��wq�����`�|H__�Pq^q��r�-\�qVy��R*#��빝��3�^�r�[�{!Â_�ÓƑ�җ%b��ԯ�܆�T�C-rܞzCڇ̋`<���Z���\�4/�vs`�E[zܬ�+Q���j"�"��C�{���{��˲4�"���(��O�y]S�8��m�$��q^3�/����{΀���uy��Vl�4DP��3��ܢkk:�����+�S��f#��eK޸s�*z�`�j����Z09br�~	�H��ȍ�)yh��K���^ߡ�^޹�`�;�-�=�GU��wIYqB�Ev���4r���v&���,�<��=�ܞ4tї<zf����R~��੗qq��LY�.���a*�f4M��I�:Q>��*�{=2�y�>��k罆�_����>3�nxӘ��;W��ZU�wF�ǈ�3��WD�^�^Z�������`�鲐��n�H��<'���Wv���#��}C��1M�ѧ�ܽ���K/�>|��G|�7�A�=>�xdK�<|2�7���]Gm��?�%�_�1/{�U��IY|�8��^�����p<8Z�J�C,z�t��.`g��rY�9�����#�w\,��m�3)��=�rޯ�������m����\)Yt���<�g5�S^õݚ�V�S��WD�=5"Y�p�Nv	��=��Ʀ��xù�e�B�4#/r�˾K���¨<*��H��ϛ�q��0���v#,	�a����q���0k�vW�=J��;<zԳ�p��T��Axl8>�ws��r���
�U+��YB�뗰E�z��׈�'>H��\8$f�G5�F�h��L�[�_z�����~E
�}��zn�4�M�:[/��/8+�Y���ֵ=�XN6G=.;���������-����7:/��>�{�=�1�/!&ܜ����#�Z���}A�F�.'�'p!.N�<�iix�������p��h���M"�ؖt}9��)YG]���֘��.���bfg �yZ����d]GK�e|�e_p�n1���Q�n�bO� �格�Ѐ����:˾�ڂ��+�{��Rgز+���x��dQ�p5c�XfKyʖ�c2r�"�S�]���*�3��L�CKVq�#t���\6��u���-�v�ۿ��ؔ��s�6����_*��S6x)�[W\�sN�&G��Wyw3��2f��?Э�l(� �X�'.��{�<3.������9�kj��	��f�L����vu\�ff֭��CjS�����g�4���+���u�+T�B#5�L�E��!���kf{g -� &���@�[�i�����û1m�n��$m#,����˳��{�y�2ڙ�|�p�)nK�G��{i�H�&�r(���s=7�[g3g��^~��>�E��=3�Lȍ�*�3)e>e�[y������3Md��l���W����wah��u�d=����oT@��]�ب�-DE${�!�P�Lk<�����c�Η�z��v�6��u�7L���ɱ*��k���$�`���p]����V�Q���n<��$�=��B��vC�z\��:�D�MNl�����[����&'WvSx^T�y��O3��2�`٢��	�[�G�+W�Y�	Ww�yb�n�K��H�޶{K\�m5�9�Of&������r�N���@fr.?6^nJ�k�v�����m=���8�t:un�+���Ɉ�����y-�����RF$�m��,�����)�'�}�i��"��tK�m���^��5y��^զ��X	8���X���C��e���ݓ���Y������l�;Z�T��Q�l�ì�Y6P|K���p\�ö��x�r���YW�t[�����d	��b�RM�PA7p/�sR�k�������*��Z��tP����`.Q���;'h���A�Mc7ҋx�ǚ������D�/+^������i*���b��"7��� ��+r�s��<���No^*�u����P�]�m|��4���z�xr�o�e-pr��Ke٭t����eq�X�|�[�=l;}�MS���uo]�A���ގ�ٚ�cE(3g5�7״U������y�=-���4h>���o{^ĞF�uN4��8��`�}+�ʵ�.y�T�Ь�+b%xq���P��.��%tU�f������Oy���6`*�������]8��D&NDI�d�,Ffe��%e�VTA�aVK�T�&2��4RRY�Pę�T�DM��ف�TC1DFVaU�E46���%R�R�MPUDfaMTLPQA�MQFNJVNMff8�P�Y�EIfeKC2�YddRQM&Y�Yb�,E����UE4VffUfeEUfa�TUSQT�Dd�a���T�1�U#DESEA��a5�TEY`�FARULfeKAUI�e6b�5IF4�TD�ITDQQYQFa�DTe��8ac�f�4C�AAf.QUd�1QTIfLQ�1QQU�ea�$UPLED��9�Re�XD0A��ՖY��M6FQATS0�fST�U9�A1$�E5DIM%Y���2MdY�aeDT�T�QI F�� �>�B
b�q�-���5;�N�����Z�jD��\F�U��)���VsV�r,k�^����q%/�C� �y'��^ �M5����J���a�p6��"9�������V|�3};��圄'#0z�ٸ�b����j�bW�X޳�`� �/�ԃ�R���m=]��uݍi��?d�Ӕ�sXP�z�zׅG��Y��P�.�4��$�kh&E�A�V��^wR1����~�V:�'Z^�ߥ��������'�bp	�1J�A�~�t�%`S�]����Q�����ML�K�\����,w��3T���k�ϦT"+'�~�����}U�t�=]�P�j ����|<q�B�N\�������EV�.�>����/^A2hx����A�Z�`�����w��S|<�w�{�EI�oJE�Ox�R�����x�����V�)���,xN"�Cm4xm⿜\#�~=��粙3��n������NRf��>��6����`y�؅1Lu֡�3�Y��g6�v8-���X[^�w�~�n��堶����,ny�iz,�R�(1�?)��g��V^}}hzĭ~`�n����f:"��I�����$���ݖ�E]F
92��U������<9��e�v��U ��WB罬��ᝫ!�QꛇX�;-]X�ļ�(����]<��sĭ��&%k��v1��sw��1;��/��=�m��?/�n�Y�����%Q�<�2�z9�����ɍ�jݝ��R%l�|v�k�wi}8�F��EW{���f��S�`ܶf}Nf�v�����߲T/��u�fopꍷo{��z�YKm���[*�-?��2�;���u,x�����#^�2)=�w�Y��[��=�� �ű�j�m4P�=�1C�&bT;Ԛi��ԭd�*�o�w��$I�˻��N+�At�ע\8+B�L!�v����*+���,��'������=��MFqIc���쳟5�8�dX���d�\�'dO�������s�蜼q=^v�oE[��ج��XS�M�2��Nzz��b�]:����&�������Z�ۺ�ݼ��|�X��ZO8�Rgg#:�	��ܻv��^�"�^�x���|=<ްAW�#��@�L�(�:��r�(y�w�x�kL��Ry3�����/Ѿw������G��p��uϛ�����o���{Ґu�Sƻ;�m�W��M���IgF�Yޥ���׫�����+Ѡxǋ�3i���ח@����Rl��˗��)np�{�>o2��L��Y}���m�;{�:]���8���{ښ�x�"����i=������7ܧY��<Y��1���v��Ng�J������F�dv+��;.�����C�I��w��gsz����9������,��B�c�Z���"��N�l�}�
�Ƹ������ֻa��~z�{A�6���-pPRP�[��j^(�̣����Ϻ���z��ݫk/0x���H�YC������<P�,k�J�I]w�}+yw�NpI��zsWp��ˣ��__S�`��*X�`b���R�`�m�cݗ�ˊ�����M���zZ����f�Y9�~�g�}�4���𴱫�Rƫ��������N�-:�f�緧sØ#���k��E>����*�� ��V}��֦UC�dW ��E���}�3w�yP�j�;ٰ��LTG�K�Nz[��cP���2��a�=�RzV�jRKG�?0%���m�NP�e�==ܱQ&l�u��m(��ϋ��zq�u��B`��KRز������~�>��3ޒ����=llKx����-�.ߧx\Bs�.q���Xx��%g�|�6�R�����3u��Ǭ��Q�R��vN;��ܷP�:9W'6�ň��7���W#3�زλ��VŒ�Uk�;J[Q��V�ΥR�5�fuYvU�R���g79��:0$3�
ߥqȭ�� �:d���i�7�l��^8M��/g���A(�������Ƣ*I�e�R�� ��G�:і'�8��3{<q�ԂT��*^�\�ۥ����7G��!�4�)�B�;��L���<�'.qW��9��q��/VQ7��S�����;賆�޴ ��S��A�McܑBޒ�c��Vexfφv�E�Y�1OJ�wkQa���U<9L]�.=/����H��)rWT��Vgk!����D��ֵ,�=��׍ʭ���%:�	y0?Ev4�mhϜ�9`��p�I/|:R=�+��//�5���c����Pe���:���ˤ�/Wlr��(�[���m%�q��}���޽�ў�hRj
ڇҩ���P��1oJ��k�J����\ s�GiWgb��4=Z�z�D���2�!���%9�w�͡mW�Z��购uGC��Vj��eUa�?=��6r�3��o0)}}2Rl[�MB�H�OU�4۰��n&=�c�8����qtW�hJY7�>͝x�fv�ĳ�m��^4o��3����xdK�痃���
���H�Ç%<�
�LJ��Oo���%y�%ܯg! �
����̙]׬���)t˻�;yZw�^B��͚�跑ΰ�]循��t/#S�s��ʣ��SުO9����x�Z2`�+��^�1O^�|GYǩf���15b@�%��%l��s[zF	.�E��`ءi02;��hǯF�Y���^�X�e.X�H}���@�Dj�0���znQ7�<���0����N^	�\���DOW���=�~���!b���Q��$u��.�l�|U�p4/�Ď=5"^����{��=��Ʀ��>"��]{ٝ�6��U!l�I�*�����J��C6u����Nv2Au�e��7u�ަ��S{�G��v�6��O��Ջ�c�S�J�\xy���< X�=wּ�b赧��7)�T�3�?erY�\K��+�7�qvRJ�^;���4����<տF�g5��z��=�7���;5\8%����_�LƲ�d/L$U��)�Gst�����WI��>�>�VW��Vr��LB̵-J�A�R�t�$�sN��ŗ2K�Y�6�ۣ뙜"4<�J��P�f����*���\	��X,K�_��M5W��pk�|�$ �5��e��=~���j=u��tdVa|"�h���O�,�v�v���].��z��;7ZZ��}��ʻ����r�.�k��v���*�
��V��wZ�=S���M��v�;�_�w5���O*��N���m������djN���z���;8�4_^i�S���!�{�R���VP:������s/�clV	��\���h����a���~����fo<��$TD�=���J�|No//Em?S�;Cԝ_2w���}��k�F�uH���t����C��B�L7�.�N�������@5�aXs0�g�@�鱳ݔp#B0�@��v���֋� ��ю����Waɾ������^�,n9�,��t�,_�47-b=>?Kj��w}9��v�HOWz>�l��{/M���r�zdG����K�7<�2�}��>[���}�i͸߼�y��;7��"ޏ��Ҷ��Ȳ���܊��>>��X��g��v������+k�+��v�چuO^���}uE���:_^[�-�,)C��`�+e�s�p�ZͰ̺w9C���w%�n���%M�Եx�9��3=~�p����B�ۂ4jp�Ќ�ig$BY�vO	*d]�0���oǽ��N4=�;�e�^4��R�l�2,���TG���_ag��;�-no;weO���{e�O>�9�qs^�h2ӱX��]�V�xY\\W��X�����9�Gw�������^t{5�g��|5��}�Q%muA����e�b����}�(�W���v���J�B�=�Z	TmkW�ԗ��{{D��p1���:\��<��WNQsˣۓ����Udc}6(��uw9��]٩�Ǧ�Oo9RнS[)*�i��76�D4˞���e�/b�řjrDM������oY�6�D�S}ݥt=��f �z2�R�	�b��f�l:���6W,�$`Q䰯S@���H��2�A�f�$d]�P�z�P���Ι��Y�^RX����W�~8��ܛ˰�"e��U�Z �T��,��ͬ��S���aJ�{j���v/o�z�����:�+�Wo������C헙�=4�GbE��[i��Ֆ������z����׳�^�:H�\�o`��J�+�1���-p�哦��-C������H�_{��
�]�ՏPR:�N�fת-u��G^sD��Uw]JS�ad��لd�#�BB�TY̽��*{� �����lx*�}����:�ƹ����$Xe�+å�]B���������=�z��վ(�t��Nq�����:��E�q�?T[bq򡙯�Nׯ�r���u�6s�PE/��x���.�r�R���4g��d|<i:v�E��^�8CK��P���`��e��9���R�1u�/���k|��X�u�Ѵ��a�"�����O����ӛm�ʓ��s;o�b9�BF�����wJ�:-f�ht��y}O�����z�R-��dln��9���QU�u<��,r�u�V�Y��Ո�k�����tɶ�
��>^��~�	��/%Y��T:�����z�Y�vp�y���lye�^g��q�ә������xg]OO
�J��E����$�{B3֎.Aěq�Z�����y�򿢜���^�3�	��b��Է�v`���m㙞K�7�$7Ȯ)�f%GC�A�g���w��':���ky`���9%m�iM���t��B0$Ҁ�S��U�eӴ�
���9p�xN�}����F��L�pO�3�%c>�����]�EF�O5=�
�e��W)�S���zBΒ׳%e�/k��������2V޾�/��IU�`^� ��Db�醮��6�F�_]�6�[�y��ٺl�A�~���z�J��=�O;��+���:KK�j?p�voX�9�`Ȓ�ٴ{=��c�{��fZ_K�X%����Ӂ�6�c�')X*��>��":$���)-�_?S����ᎋ1���%U�K��>"�`�H�\G�v%���{מ�Q��twtl���8�T�8b��>��n(:�񿙺�n$4���Ah_طqm��ttk��&�WoU���*�vk8�ZȠ����������Ri���K��V'�eQ��r�V�A�����G�n���Mt&�^�ξ$�w�9u�f=���m�%f`S��:���ٳ^�g����7��W��0�&cD���L��?W�Й����g���ў��>��r��[6k�ie�K����sƜ�O���kO��,��Us��e������G�V��xm��e{���2RU٨^(O	�sƝLn�Gk!��w*]"�1�����1֠������M�{������Zur��Z��p�_�������=�{�W&��V�S!�۱�`�3�J��c#�{��V�3����u	A�~��p�����;=6zC�V�&��]��|a'�32����z��A��xOK��߲�e/,������M{��(�jR�O+����q#��?�.';G�J~��ꂘ�j��_��=ձ�-�l�����͂:�E�p8�K@��N�e��a�t�꧲Gᓜ�O/P��8-C��,M[2=s�19keY��fVTl�.i���ܘ�J�EO���v["ǩs���2��^e���E��NR�l�!ŞH7=��E^��!�>.mg��6��~S�$t�W'�#����@�1���3Ma��� ������(�����G=W���t"�h��̌�.�3F�꽾P>Ȥ���M
�]F+���Ź4�^��G7_�zp��vN��l=�4�*={]�]�Yur��^/����6ڀ)\�ՠ��g�߱p��F^	�;�U}.�4�.I&cT^�vxM����*���o����4:��C��|�C5։~�8_J�^���YϦT�+�u�C����ߦ�Y�[�O����+P{6� ���{��6��߻78E�1��P�\}2���n������dܵ�;2�B�5�Xk��T=�՚��G��{]ёY�����cu�q���9�7/��W,��L��]���*��im��i���o���Z*O�zR7�w���9��{���u�P�בּ����gå���fB_Q�U�g��3�>��x�Yo�+�KG'f�nv_��/jt��`��~s9�XY՝0�;&�)�c��Bt	f��^�Iu��<��k<`�v������8k���.��+�|Y>��6Ƶn�M��`���=�D�6�z>��w�Wö�np�ͫ����ȏ��%Q�<�2����{��[�a�ٲ�+����~��t�s�֙��R�5�\E�L�*�E���t�S�f��g�v���o������Lx[H�ޕ�;�7)���
-V��Ʋ����al��2A;
 ���%]]t��IjU�F�ų���!���@#�	�G�s��멤2�vH���ōN%��:��.m<��d��q��+ Х1Q3��U�;�s�[Kl�2�ɥ1E���fի)����D*�6!s�y��Ʋ��z�][ʎ[��E�`�֑nɤ��M�3�զ�#Q�<]L�ڞ�h���Y=���	8@�yїª��G� R���h�r�[���]#ٟ#�t{"�Z�A:��C5˻�3:v��_aȖ�^�s�5`/�%{_�����cFvɎ��{�o-�n�
K2���W���6u���(#��Q�خ�Q,��%%ֺrUO9��=}��d��/nY��&t��n3eE
	��+v��V���dŢTE�2�'�-�gw{<�������:��R�n�}Z]>�$ksU yov����\�H�C7�F&Ԯ)o�uŽ�6o]�\��V��5@0't���.�5�*�MոgG���U'o�����$'=o���{�˳9�N����Wv�R�B�sC����c(�&tW#��P�����mL������ú�!A�>���{�c�i:
�	V���,싳L�|��4�d�_W�6�_��Z-�֩�U��C-	%��w�gT�O���-Ș�=dM�Mi�(�G8��g����⢋�bMɜ{�s^��{���J���mT}��%Ꮛٝ�Rby�f��o�}��.i���gE�o� ���ކ靆i=� =�V,�y�<�w���6�r�axz�����G��3,U���Ƙu����)-ċ{�������sm��H;�t�'NA[�_Z�������C�:z;�D�t*�vY����fS*7K��LǊh�)-[\��ݓ�D��x��);��5*����L쳏.�{� T�T��њ{&����X���'Ea�n�W����8�6������q���d��c6��ڝ�����"o��c&���Y�)�[�~4U��`/,�1��\������ż���<�6�ݫ�ӱU�d�ιN��D�ڻ!��w:v����o�}6�E!u��Z�)�Ws�C�h���B4^.d�N?�žǇ���/^�0�C�v�}����>�y��y�аe�Pռ�7���ĝ�^��iB�n��⎞�RA�#�`OV��j
��	��{�|ǽn^�<�㱔s@�/i�ɃI*s^>�7w�8��|j��_9�J7�%��Ȗ�*�M[���cit��5s% �-zv�ִ�:����6�f��Y��E]è���u���A��F�+J�*��A�*e<�7�3`�^Z�䦽H�dE�����.�.�VW��L�#���9-2]�N����Rh�[�p��[C����@��()�N��C�O������\!�.�Lswǫ��iru�Y���O���|@UQMUM�i(�*�2"�(����'$���30ĉ"�,�Ț������H�1����,��,(ʲ"����"��ƫ1\���̢*���j��l��*&��) �����2��p��*������3
j������3,�̳
*��3(�������*��2f�h�#,(�b!��̚f���s�*��31(���3�����"h����23�)(#,h��̂�b"�(���a�&�j��
 �(��j��L�+#"��̱Ĉ�,�)ri�(�(�2$�"H�b�))�,̉��(�� 0�2���rŚ)*�ʠ*(�$���̱�3"*j'33��K31̈�,̤��,b�,̂ʜ*�h��ʢ)��*l��r���	��0��0��*�̉��Ȭ32"��(�2�0�*��bj��0i����ƒ$�m��)�=��[c�5�ܡ+=�spE�X���~S���L��L��x�͋�����62���a�:�(Cc͋������8�(��o_�EY�1��/ڲ��C��(0B��9��S-g�a�2��>'��sRlK��xPe�h�y��c�}�Z#E��%��EV�.�Z�M�Rw��Q��K���<�l:�����W��S~�K���|3�,�2���$�<����H�yz��N[���󊸇E5xl��>�9�qs^��a�bv+�K���t�wѝ�*C�u���q�~�P
ǯ:���v!as�6�}�.{��积��/]��1=b���|���l{��~@�-4�6��)���4eq6�����K;�ϋ�f�~K��sr�Y��o�+<ܷ(B��J�s\�g�*%�;\�w{)�^�I1S�V��=#ɾ��gu��Mj2eø%�	g>8I�ҰY���et8��Q{(����4���[w��.�Q�:�!��=\�<2P�n^f|��4Y��3��-3ՑD�������O5</��v��r;-foL��*��38�Z�Y:n,�򲏶�X���œ�g�w<����)LxHyvWKd�е���wuK�s7���J��Z�#1�5;
��i1�6���E�����@{S��X����"�ڄ�7�43�ޥ�y�w���W���U��F�㜢������OX��0w�#��i�3CiV��L7t��'B.S���_�Ś<��i��T�k��~r��K�:�l�m�{t�6����fK~���}:s(�+�_�ʥ�Lp_S��x_�1�"�U�c�J�P�s-�C6Μ~�#�7x��۵62�5����A����b�8��m}�[�{o�\T|lK�mR���d�O��l!M�H�(?O>U�+�ƭJ]�}v�v(�x�>�Ҵ[Y~׵R5[�r��-#�~Lz;�o����^����jϰUz��U�yC�X4�Z�$�-���-v��T!�b�̇˥�^5�}�!���;8{j��=1��L��M6�3��v��M�ě�E���(�)�L�z�'gZ�&
�Z��)����o�U����PV՘���v^}UF�zh?/4Ky7�Bs��{Q�����:�=��E��mD��ٍ`��!�ԴKZyJ��N�9R��'.
J�0�ey=��"��ǈ-���c�ѫw�O���;*�hwh� �5C���֙��X��u�o,���fEv�����V+�bҕ�GJ���K���d�\�t�������9	u�YO�R�n:�{�ϲ�/WRu_܍KV�CB�\/F9�+!�w�C9�+�Z�PǢ�vsW�[���J�_�ɭy��S"��777-�q�3ÝXzc��rG=
ȡ^������_�����xO[9�W�0ؘh�����*�4*��>��Ћ���qI�UR�Q=�u�~�(W��%L]�.=���'�#_t��_�L��;�<v�	�~\Z��#�|�]0}YT���e�,3�g��`~�Ev4�mh���>�.����t�-yAr��i��ۻ�i�]P������>2��ά>ުK��B�Ev�Ϝ�F�`9G�+7^�0�{;Iݸ}���ukltݴ�0�E�=�lի�S>�1`ޗEk�J߂f4L��v3��[��n��a&�O�G��Y�͚��˗�����u1S�>v�#<X3=ݶ�z�����>��f��!�G�r<������{V6 ����ES>���oٷa�245g+W��t�K/ۮm�j�,z(`>:�[K=6��P�1*z�#*����u�]�d�x�ӆS�ݿOU���3%�ִ��ݎ�9v=�J��y�ܴc���SV�V��y�kY��s6�/��Aa6xT����>u�^�32��9O��OW�L�;��3ծ����_kE]w�E6�����іSɳ��%�Ow /�t4+����Ume�����Z�K�Ȉ��~�������Kb���x�ޮX7O-t*���]��su����k�&^�}i����4N%��:�-^�M���C�����ۯ���b��������X�`��8��1R%�z\ ��'�=�^�����)u-�����=�Q�we�B֚�#�4P��饔����zi��AX�;�rr�*j�/$�r��<��^��;�tYbof�*��I��H�j�]��N�'=*�ֽ4�=�T��7;[�ˍ�x�7��<�-oe8W��(�(�}�+�$��?��O{��q��~�����Ȏ��?k~=��'�����B2�L�ر�WK�|�.I�\v�Gѳ;U��N��o��F�/�Z�V�!�����+���z�!g&TŒ�,=����>o��?7��2�#\�w�p���.�/�Ӈ��,w��3TΘe-��¹J��󏝻�" �P��$(o���9�~�L<&⡱^rC���o�۝r�4�_��w�����O}��!��M	�v/|)>[yv�6�o�w-"�N��uCO.��enk�*�)�6*9��=K>�d��88����;U�|�ee��Ʈ�u�MNǵëk[0��r�w��:�fh������Y���rs葐�h���X��*B���3�}ޒ��R�m]`�ޭJnDP�ތ,�j�8��u�GY�s�v3��u|�1��q�;��8�a����u�k�c_;�'���a�Ms罯t��.i�s��/�WF.��	^0p�+} �����Aεo�Nt��9�"�=��.`�}��c5�xy5{��θ�౸�ƖJ�\��^c�`WKx׭m�w:v��~ٞ�5S�:^V6U���O�V�{�v�c�K�7Σ(d�}��"<��*f�tۓڦ{սnv�&������M�
�ԋ�:��s��N%����NfQ�2��w[���0���������q�h�P�𹾣�>�j�gԶп����0El��ip�d�NN��N��8M}�T˞re�C}7����p�VZ<l-5�`��O �C�L!��e�B�׻j��r�s(��ޔ�5�ql:�ϓ��zq���'{̳�^4��xȘ;Cn�g?*&U���Y��{=��ܺ�6���U�BE5lF'<�,����{�N6�P�T�p.�яHT=3|�h\}��b���PP��v^}T;��ۛP���91���qZU�z�4�¼��et^�|�w��2e��KA���B���Sr��\��s��淖9n%�̚XU����4�Ks�y֭��y)��{F�B:}�$�vޤ5�u
��e¥�6�&�?6�bO�!s��Y�vg�n�rD���բ×��L��i��4QŢ[���2{��*�`��6�T�z'���R�Xի&���˷޶q�;P���(BjW�.k�L��D���k�r����ɍx]M�V�n���V��[kLC|�	����%� �$-t������ ����4ʵ��B���v�C������^^��cW}���g�	B�y�a~),TӖx?e�͗�c��HZn��&�e��3��gQ��ޘ)+��
K����ܲt�Yj~��'��0�ɼ�w���!���1:L�eY�L�poK��k���|��(���m�oz������p>��~���-��>�aJ�=���~R�7�U�{�x����D���B=~���MM�]{��u�vs�ְ��:��ʴd/��V��g���խA��,�ڧ�-�co��t�K=O��F�/,�ʯu�6��*�}9���_�����K��s��Y��y�M.��qіX�/��)�Ť8���w�\�����mT��-��a�>�u�z�v��5�M�B��Ԣk)��N]át��F��1�!�r��ԩ1��gl�:���Kݒ��1i�p�#1�`���[�.��=��^ݯ��T��G���y���١��HLr����d2�@T�����>���_�4S����響���o�;������Gq}Jǁ�e����ٷ�J{O�*e�s.E�	��������:n���'��2M������V"��S��8_�P��׭�{���'��-�5�q��
Q+K�e:��qx˲�4��.���gܽf��ӭ
�䏯ދq]2�[����b��Qh%�m-�"��N�9R��|��G�'Z0wF<�J�
���3w��۾�}�f���zP�V��G�;����h%�L�C���r����tR�����Op��"f�����/<Y>��r,$�,�u�I`�/�
(�v�1��ٳۉݹ��pd|�Q���J�j�P�Y%L]�.=/���'�#C�.K���n[wjW�'��wE�1JϾ�lQ5��Pׂ��f��Ev4���6�`X��_��~����|���;o��7ΒU��
�M/e������h��x�t���|�4��N8��n��y��\�}}rV_��I���Yk�E�\+w�1`ޗE^���y}j��{�<; K�������"g�S$Ɖ�2�W������/����۞4�������_'\l"�u�+�,�>�;��C�ɷNj��I��jr���G$�V��A�v��=��/���-H�{��.u�[ʇM�bs-�6���k�૤�%��$o�����l���.�u��s���t�KNߌ�͜&�ЋE�.o?y�Vk��t�8��6ȗqIx�3�AFlv�<�����=/l!{b�v�1<K��}���Sw3Qi�ҩ=���>̫e��.ܱ�5�u��į+���A����j��Y�bԐVá��NH�3=�`��]���3��-!�n�5��`�P��:�up�����-U���i�쥩g��~��T������>�ZU��M_T��w�v�15C��}�A��U{/oS#6�/�g��u��~{�a�+�+-g���\\�q#�ΤK=.\�Q���~�E��W��q�G�����h�R�5�-4�:�E����ƚXyq�&(\�_������x�@<�q���˜kܟeQ�wh�.5��K�d��z���>� �Yqn)�YOW�&է�ݰ�f�sUxeo�eWm�4rA��Rp��k�y�Ѧ/Ċu^���z���l	�y��'���fŀ9���t����H7�P�w��w��RIa栠�|hKC��|�C5։~�8_J�^�192�*��I��%D�d�s Y��,�@���'Yڍzj��/�9�M��Hp�c6ε��S�G.X1�-�5ۀ���R�ܒ��+�5�/�޼�����KE��ϸD7������#w��|�Bl �8+����6�|�OO��['�'Tm�eo��B�Y���~�~��9}��8'�xޞMp�	h�,t����*,�Q��x��i��>+H4xK$��8-%�Z<���k����p�ֶ�=S�]Z��=���)=5U�N�����ݑ|�M	�v/
O���h�P���T�,��9Y�/Z�w�o��{�)O�������,�t�v��fh���z��=��Ks�����^33����C7��K�,+s8"�ά0�7�ݔp#~��|V03��s���o�
�m��u᾽���눱��-��+�rPhC�܇8j������#'���]�Ǿ�^Ge�m:^V=mpvW��x���~3 ���;��V���٢��{�t|�l�ȏ�e�v�T,m5n���:)�¬����҇P�x{�̏��6]�����VT�l}W�}|����MC������\�Qӂq�Ճ�[hZt9]@Vˀ��O���c�Lތ�fN���S���=�޷��%ùYh�:V�J��b��G<:M�y&���Lo'�\;|��,��D�!��d�6�ya	\y�*A�&�N�tH ���˼��E�l��7�i\3�Xˈ��k�n��҅�>j�d��s�g9�\*���vk'Y�Q�7)k3?%\}��Jw�b�K'�r2�g��B(�7��w<�CM�K��(�Ǹ�6\�{'@~�+�.�|0�0�K`�i���1�o���\���{�,UN*�ձ��}�p���xN6;��r��:�c+w/������]*P'H�`�y�2�Qn�v!as�6�D4˞���^Y8�7���G���yNΌ֩���U pr�h6S/(S2�SG�-a��}gs�o=-��#�K���Ni�)0���c}坧hyQ�g��!��+R�>�L��2�P����,5��c�r��}�7�϶{�6��<}7���p�}/�K8p��ZU�N�Y�Ъt��|$ޙ1Q�y�,k����&
7dA�+����VxD!����<1dX�SK7�==kU����}5�F�u>��߳sǽ�f,ޖ).T!_�f0\E�哦�1���ym�S��5��myz}�$a����L�z����mC���-pPZ$���+Ԕ�>rKYw���{���BU�Ȅ�Z6}5 柶�ɬ�"����������g{@>��(�g����Km;KdY�`ݼ1�<o,Y}���Yb�#] w.qͣT�8�"&.<�ɢѢ���2^ ���ܼ�6<�t�l7�.�����\����V��=}EՈx�K�:��Vs��f��f�����E7��8Ge���=|�Ǐ�;�P����G�<&,��iznV(d�,yڷ 7;��K�l�ە�A?�d�<|-�M�ts�-����\����f�T��Pb��x'hL��e-Ͱ�K���,�r���ե����/_d�M����2ŋ��x;'j�J��m-��%��"ӄmEw�5�}].n�fWE��+,.�Fs{ʲٟ>�n���u�^�E�ZޔR����ʰ����	*�m�ok��Lk֡�lL�KD�w.w#�0+��xs��t�J������4�X߳������D��<^tוy ��Nx��`,ܤw�ĸu�x�S��ƽ��ڭ˜Χ�����Z����W�z��&��"�)9l��l�Z�n4*1�WW�8V0HQ�ћ�A���]vn�ai�jӭ�<�i&�n�m�ˎ�74	N�Xt�ވ�2�`j��G@�y�����3t�r��ύ���2��;�-���ZحY�����4Y�������A�Cf��u<{�j�b[��H٦����y,W�zi*����g�C[��γ0u�79�GW�M��ӝ�k?!�lQ$=�μ�Qd��I���E��Z� tp����
"��k��P�����c��'	��,��0Y`��4��IF��ܤ8�l-G$�Q�����e �Y�b�wx�+$�Ү�Q#B2�gӲ�ʛ _
�/z�I�M�����
d�\\�/���lX�XݽE�,��|(�ɑM��fʱZ�򕶺���w��&�R��'o���ڣ'<2�t[�z���Gh��>���E��\�4����)�(����ڒ�{$#p<α��P����g��VroH���ÊH����:7�v�vs���'��X���tU����b X�}ޚz�8�0�5E��[�:4�3�����`=�]u��"V�m�f�}G2F��V��c*+�ǚ�ht���Vt��ѝN��3�dV���CGs�;��g�
{��b��q0y�2��=�Y�OL�%��~v�+�NLK6PPA�a�D��VCu���m!ś�l��������nV�.�_i}�~ғ5vEQc�_CO��8�v�Eqb�:V1��^Cޱ���xXt<NRɑm��^�z��)�m����	��ޖ�y��n�4�������:
���ԵVR�c��|��6��=9.�y�[}�.�� �A����Y�� ��<��R~�m˂3ۧ�H�j}{$��\V�rN:z��Xos���f�l��Y��!ȝ����7��ټ�=ϒɕ��R����e[��ޞϕs���{�T5SD5VYU��RC,AD-E�f3T�5U0�SQC�a�dT41EFYD�M�DAESASQ���AAUT�QE4UUYd�A��UVFPQM1UU3QU�1R�UEYTT�3EY�dQIe�TYeS��AT�PMAfd�E�d�ՙfI٘Q�ERQIE5E�PM����LTEA$�QUM4�PT�XYL�MQTEQIa�U��4LTU4Uf9QAFFISTTQNf%LY�ESITMD0C0EFf�Q3Y�ADDTFV8M�E2DdaAD�d�EAfVE��LHD�YYPe�RFY98dafSKQ�Mc�fbfaNa�M�QM%�aAAAIM��VA�RDSRf94RS��TM%���T��T�UT��Ha98�DY���S��ԧ�Wp���:��c�s-���=W&�X����T�eHZ���fra�a��]V�d�!�u����m){�)o���~�79����]�po�yB��W���7�+k�%"ў��ǳT�����fL�o��x��K'׾�B��$]{��<�i�9�ʮ�ڿe3��u£�!ym�ރٞ&o�⒇�`�L`ܶfS��O�������+��>z'ۡ1r��|��{�Wu5�m�{��}6:Z�uQ�٢�\���z�Qe2I˸OJ�&cP��2�>�7�q��}�A�~t��ΩR�V�i%ۖM�ޤ[+>{J(g!8�oW�gZ��v=Z��>�s�d�ܳ��*���Q-� ��-��˲�4����~X��?N�������_�sz�h��q�k5��G�a��Qh$��m-�`�\^];L��-	˄yӞCu��\�NJ���w5Sm�cޙ�Ŀ���*�o��(F�_%�L�C���֙�~�=�k�=x�:��jڊm�ײ�O�����>��{��g0J�&�"N���;�nd#ˁSٻ(0�Oq�,,庱t�u�Y��*�>��.�Od8r_�Âx�3}W�/Ht�.׻4���B�<���{]9ѾGkkY8���N�'AV����\���L��mߚ�{^<����P��B����'sm!hd�E9�j\���-�[��l�H"�U���Vn�et�K�3����-~��Gx1c��O�;7tן�b�>�+K�����hg}\��Pg�:�c�WcN9F֌r��s��s��2�k'.~l{�k��h���fR墓����Ŏyla�^kD����U��P��)w�"Y��^ɟ���G�7G��˱5��G/�j�8VY|*#�1�e��f	G�)2<�5�>Rf� ��(@Ͻ�| ������J}�͚鴲�\�//��9�Y��z���-�^C�-$�N��
�ǼY[*���ρ�ORΖH��3pQ��]5�"\/ݥ�"o(gTd��ܞ�6�ǻ~Bd�ז���rǢƠ:m�%y_��1O\,Wc�q����])d���-|��Z��JgS7�w��imP溜��P��dwr߱�����b�o�Lz}N7���֙�Ek�V2K����"U����ƙ�N^	��Y�2\��u�����ǽ�t��>��z6�dX`���F�����S��8��1R%�z\#fi���l��%�pܥ��;��/ϭUx�����=��A�u't�l�w�c4�*�sM��LW�~P1�bޡOh���ۃE�:���e7��������V�E�"1Uu�tn ܽJ����zp��J�T�K��<��b�?p:�Ɇ����	��n���\l�i4���_4�������Uҧ�ቮ+��E�+a��z�j*}�w\�?ϴ���a��c3��]��]�v�6�o�`�ω8���Q�Х3B�E�5�ݙ|5ejCe�;����re�W���q��fQD�)r)��4��]%Ѫ�=��۽�A}���}�.��է�Cs��q{��e������{��e��o\c��רn�J�V����|h;��t�ϓ�f��/פ>�zg��M`��zw-�^z�cX��==Ǧ��u�Xx'�\�J�:��|.���G_�rƉ�Cח�}�["��� Iڗ��ٹ�r�:x����2$�&�I���r��>o�]�����Cb�~��2T�����]��Ն�SD���O��;r�ȇ�4%��)>[uL�țܓy��sp�9�藳�2T�f炕��*9�VX6৩`�d閨�ɴ'u�������8����e��ש��Ԛ�����o�a3;��9��:��N����3���W$�<��9��20��8����)jͻ�{}{���c\7�Ɨ�ȵ-���J��S"�ɺ���|k��ߩ��X1��+�!�2) �>Ш��²F���Ϸd���ї2A�jէ�o���8��N:���W�0A��^C9�{�zь�RL�&nr;���Uqw�Z!�,���i�Z���g"ߚG��~��r֨��뫂��m��<μ��z����aw�D}�e�̒����dN�܏5ݷ괵^s�ޅ���;^*�g<eY��
F�=���&{��"if\z8�kب�徝ڪF��m=�>��z�z;��FJ�����98���[hZt9]�P�����K�+sR�^�a�B:,5�f'S�<�c�&��]�.��F,[߮�GK�w�1&4=���Ț�'��Cmiiw�i���"͗:�.W4���^�p�tL�s���M�e�[|��a^.,T��.�����Y�⚶#�}�C���'�y���T��������q��[gŝDm0xȲ�fc�/@��_˝���7��m�2��e�Vk�{���k�v����ڹԈ��ť�w����̱�җ��x�˝�.���,�jKv=�l��q�wj��'�g���Y�K�P �CZ���
g�eD������=]>N�);ܒ�Ͼ�k�:����\W��~P�#�.�/�K8F����]i�w��ͱ��
x���v�˲�J�����R���'rkyF-_\��ԅ�ǵ�S����(�������jf3rܞم�+q)3w�w+%P�+�Yࣽ6c�.֮|��@�z�:�Z����%ң�We�,�V�i��2V��{B���G5N�Rϫx_/Y�_Kdu�|����τ�ʻ��H�돜ݵ�d{���	�)ir�>��_�s�wQ����%rT!X�1��Qk�,�>�C8���qL��;�n��8=Wh�� S�Y��Mۃ�>��t��pXV$����K��p�v�&y6���<O���?-�\���dq���p��~��V���*�H�w|��ݕyڻ�w^-%A�|I�?�{S5��^P�sU�c��VՂ=JE��+VRͻ5]ӹ���I��18����ɔ=�u��t���÷����/)y��Á�E�<"��V�͏l" �]�8aؘ�7-��K^:�����
k=�6}�ؒ��9�{���9w�j��]����9[*�!�PQZj$�qu9���oW�1�u�&C�ڮ�>��݆��t��|o��x�(*���rɯ��{���Ҋ✄S����<��u��&�����C����Զ,��/*��U�Q�m����.��vw��Fzo�`�W��(3�Z�)C�������a�	2�kP��G�y*:����wz6����Nخe")�#���)�r��X0f��9ܧZ����LYէU\:�<s0C�-x��fj0u��鶪h���Ed��S:]qRk}�h�`�V%��5�,O\^���>t5���Ӎo,�XxƂM-�[Eqz.��TO{�q�C�W��5����m���'j�0v'�7��StYbu١Hp�@	����t�\cוۊm>��{;g�qx�[�ïe^���'?{���,����+Ęe�NΑ$����n��y�R��cJ�v��q��,庱t�u�үڃ��P�Y%L]�.=/�ᰨ�뻗��{�8k�z�#�OQ�--��\1O\�ޝWz��şKɁ��Ɨ�ﳂ��s|�~���~��;=��.���VI��Y�\yIp�E������h�����i��}�G���
��E�t=U:��C=��=�'�m%����R��|.�-_��/�g�}^[��2?랫�`���@7�#Dۂ�&��D�̫�޵��9���'w�5��$r���G�v����ne��/��[�ZU�wF�ǈ�y=KK$P���Gx��χQ��|������A[��jV��~eMÊ�/�ո��ۖ=�:l=������=�P`���A�Rm��>i��p�.�V�Z|�tE9�M�� �(n`&;7nP�O�B�7��:�^v0,�C�ɹՐ�[kd��T��k2]F$�i��M�V��̖tv��I�cr�W
 JH��w;M<�`�=;���aq��|�m���,+�����gI��7�w����/�p�\�𘗨g��Hc6�sX)���uJ�����(�t��ՙR(��^��ܱ��1�1�e��X�e/,�����"U_= b<<{ו��-���OC닗�M��Zƚ���=^%��~�����u/Z�R��L�_S�b�I҅��a^x^��=;�;n�a=���{BqS�P�g��j妃6�N�*0��[��Hn�=���d�r��ԓд���FX���	��|'�,�t{�E�\k�vӻ���t���"��d̨]�:}3gZ0��yg �C{���^G��K4Iy��żNR]o$�4O6��R �f��˩	T��ς�m=Zj������B2���Ol��9�1�[�������^����k|`�@�K�JӠ��ﺇM�	�3]J���_J�.��{;���G�Oy-��\P�	�a�)V�F���K\�9�o�l�u��:p�^��r�*ޯg�1��O��U��-@s��X,L���B��䮝q��k�S�ؿ[�HL�e��R�ۥrOx�c;w���c�;\�Z��er�%2�ult���<=�2r��r/�{��n�=�?j ߙ��oY/�:���=�5V@�nK%��Ef���n�({[B�B�ͱ�9ץ
���)�N�kWr��FA��3�L�y涕��PN���W"XpS�s�;*��|��8.��I��:o8���c9*�us�,X�-�L��K���eZ�<�EG ��Â��҉���+0�G����W<��ߴ��w5�:GΨ/)�̗�{��؆oK�pXV<�0a�ϖ��t�ߙ~ۓo�>�n��hxAPc�B�Y�1�fW�@u�!�pX�sSn�k0�Y��sq�Թ�'�Pc)�ci�v}��VY⇷/���y�oՋ��SqgD�͜�ڧ�7�}���89ۅ�c�i�lee�Fx�:)�<*���x�����fU�MN�,:ěp�'L�}��VrҀL�3)�þ;P�Gq�nJ����-��>G���Z@�V.�Q�^���c�����g�-�c�߅Ր�2�����c�&��]r��x�+L����r;��s�{s��+��f�
ʶ(B�KýI��縋6\���N+�~{�A��g��5ݘB�Rs�Ӝ\%��F�PȒ\f��#���W��⚽��1X�}�p��� <3xUg��^�s� ���J����O&�A�qL{[����۵tNwPe���Y�&`T��.9e(�B�[�׆cO$~/�Z�\����G�{�)�9'�=T#��m���Ol�o��&]����{5Z3C� Ύ�s˕�ǘIxg��+ZC׈�ͼP���Hh�'�)�9I�<,�.,���1ݗ�U�,.v����L{ڻ°�Ū�w��m?d��d�[�ؼ�ڜ�e�����mu2�P�e�4�.#���{����/=͛�Яu�u��Ђ�7`�U�;N��5��СFx[$��<~���M�<�^��3m,;���[���J���T��V�p�Q��� (�#��y�ޙ���ɫ����,���fWC���"�0�;�(�u������<2P�n^fk��G	�}�M���|�F"bF�[��z���b�ޘ))!h�1��w�q�-������N=�=�'d6=^�l��@T
���h�������|&o�%�y��-	���[�3&���u�<��J�X������}��L��z��lpU������8����ϸ�9���5rܞ���]4�eU�̈��;�Ε�a����ʰ0����nu���{�훃)]�3���/�`	�gN|�ݤmR��l��[jy��Ú<��\uw}%09k�xP^���S�R��^�>��
���k�z���(R{qJ[��D�:�ڼ�=�+���*�`�.����e>סI��풣��,�� ����}�+�(�zF�O{�6��7����5͇#�&��AX|��sW��v�}�c���%˸�@��0
w1i�.'���#��㺼|�_���%�����=��BA�h�щX�(P����;Ԛ�2V)��|Kz�cP���f�VlѨ�y�V�A�����]ȳ��>1%�������	=�ew�iEE9	���u>�\n	s���;����/�zP�*�h�G<mjc�ȭ)��Ғ�`U�^�t�����ьK����1�x^	Bs�N5��?+ TGI����-�gս�Q�v��a�ɜ%�3���n�I��O���Ԍsۜl����9�C�[�]�v�Y%�E��sc2Э�������=}k���jr�ײ�O�$��a�*b�=l�	^$�ba�|U��?jC-S�;鋃���"LarС��8�vr�G�C��_���"��:{ ���-�^�i+t�gOTz������K��U�Vgk�ý������;	y0?�Ɣ"}Wy�$�=�;7n������|ݎ�_�ÓԒ��^+�^]�����΄��"�T�Xg�e�X��.U]e�����I�;��j�/�qELܙq����h���/5�+�����u�;��1��vr�EF!��IQv��LD�__c�Ǎ�H��";� \6[㫭��ޥ�G�O��{`#T�<�v%]ҫ3���+���Q�b֡�ئ�iF�v���#o��Wg;�%i̫�����f�W�~rY�e��L�ׁ�N�$}@C�|��N�cJ�#��!���%�G,��+{���EhG&�*9��YU/wW��]��,k:�nÖ�̺�m�w���cf��hؔ:�>�MV<�"^�u(!�2PF���5�>������۪����+û�GI7ة�Ư��:�����`m\Zj�������x_p�J�9�wQ�ǳ�ȥH�,A:�ҏ�g����s����`{�r>2a��ada�`F8w7��E��,�\Igǎ]�m]�}84<��@�1C���j����#ҜX9<��r����ݠ� ����6���+�5��[$Nk��8��A�7W����`w|o7�w���;�_K8!����u9��F���L�&�p/5A�Ɵ*��:[�N�O�x�i�X�^�	��D��FF(�M����|e$�B���(3@�+2e�r���c�ȪY������ݲV҈[ʯ�+d�t:��4��yb���d�Gi��<z�_)}5|p��v��. �-t.Jz�V���o���J��	�M�U3���*Z[B�n}�ͦ#�Wc�1�h�&s��/��t(���f�C�uѹ+�v 	��^Ūl�ᙐhO��\�x��k��լ��h$�Y���4q�SR���M��q��z�^�'�Gm'�#	F�l�Ŏ !�-#ft����Xv�Bc��j+���[�⼝,O���oS��|N'���n�s���K��;��.�`�(�D�t;���fOho-�$U�f��{���OC7J�x��ܬ�,Ve�x�_��L��HVe��ԫm-�̔�sE�,�\�xf�J[4z�����6	��|�{�;��0�6�?0Lx]}wocK�}��ٱ����_t��
��zZ&�/
������(\iep=�֭K�s.t�/gJx�)4�G�^���c4���5����o��%�x��w7����XS�y>o��<2�$�zH�ēȅ�o�}�!yw�MH���a�����}:��F!�p}y��Iw�+��+x�Թ�;�Ž{��k��uN��F�n�Y�A,������*�S.�s�*é�c�&�j���ZtG�Jc��SJ6��¤<�MЉ�u`KO��ީ�������o�tK:�;<O_���@k���1=���N��1��䥂E�øf�v��;�@�G��3��{pi��|x�}`)���0�5S�����Y,�ħT�f'i��*;�.֚={��PΩ��K���}���~i�u�D4�D�D�P��M59�AMSB�cFfSCLBMEESPTSTDDٙQACAAQ!I4U�PQQ�MQPUEE4%Q3MUT�T0T�1@TETE�dDQUQEDERDTMQM0Ifd�LY&EQTTU5e�RS@e�Vf2D�EQEUUfaM)M&MMPDddAU�d�UEAADSM%SICKMEL4�D�f	�ĥR�PRDe�EMT�UY�$D�5SHUDU�AUEDUSMU��9R�U5Y8MUCRR�TUED14�AAQ5UQ0f��E5EUDPD5AVb���ALL�4�Y�a5D�STdd�FVcA�DDMQ��QNFQA5QT3P�Td�S�d4�U-D1QES�d���!T%D�MDMd��UO�y��o��m͹,,^����{�<��-�v�~^�[ٷl���Ժ�q���L�V�Ǘ����L=�s��d��-��%�t��C�{�
t;�i�n`�=��6�~WR��|�"�_��`�����w��s���7帧ӝ�W�a*��6�I��9��Y޵�p��N����R�vgc�hn��=��&J_�ػˢү��(�{"&'�Q!���j��W_VU����N6;�2N��~�Ռ��T'(_�mǑ�]�������W��n_�j������}r���[ٷ������p�\��L���V����
s0kP��_R\�I�#�s�s����9�o<�#̱�3XZ�61���u9����e���������s������N�]c��[�qu���=o�,?p��6ϥ/=���8��UL��݋5������J>�E��`����hzq����;���L]pυK<A���}�M��ſ Қ��V��}�W%c�T3|'b2���0�:�s�{��=�ݢͮ5��SkO>��Ϋ��SǮ���$Fj�۱0
w�X>i���\�<��e�W�4�τ~�,����U𾱹U�)��3o��;!�F��tm�2�͂�Ñ������oR5��mo��d�R;�{�*ͻ�'�	��wm�7ݽS>�U|�:��͖9�H��J�:���<s��-_C��#F�k�7�_#�H e�=��j\�񩧵���_S����=Y�|Eq��A�/��&����s�¾�
�5�vx&#[��y�}�GԷU��K�9K��T�iȮ(>�6��_��[�,aa<팚=����Y7�63��9n-�,ϦTŀK����@�:G��u�p����\��I�G����W�ݓ{�GY���žg���92�%`�1��B���\e��<��wr]_�|Vm0�Ǯ����eg�]�J�Ϣ�h�pS�p;r�ȇ�4%��\یb*�{/Ƥ~v������`w1ޛ�Z*Lޔ�����CVX6�.�O�)��;���|K��p�ʓc�|�8�A�g��q����3�*������cR��
��0pE��A&ʯ^+*����#��S�� �<�n�f��pLo��1�>�N�+)��)��㹆��}�>�����4�< ���^�2G��Ki��cҮ[7�VѯV��NY�U��|�{Ҷ��Y���.��댡��c�+yC��to�id^��]���Μ��^}T�#f1%җ��o"�7� ��L��fϱ� ���br�����pY.�VE�\ӝn5և5����#wc��Դ蕏:�t��L����Æ��s� b�C��E��L��؇�܆�r�M9�.�<<��o�Q�1�Nm[m���b��=A����zU��;�v��z;��⇵�s}GN	ƯVR�B��`�Ui/�b��=S��jB����
���S-`���r�Υ�7�g3���{{�A+:�D��Պ�b5��S|�ٺ9 ��O)P�]AC�1.Ěi��Y��T8��xN5��hgf,8�d���>p��hcօ�eY���D����*�g��j��1X�����U*s}ݭ�Nr�<6���a�s�X�k���
���	���s�����;;��ƧsI�OWS����j|<��Nzz��b�ڱ:���h���mu2�3,e4���-HLف�ƣ/��������m���w��[��?<�9���ό�B\�A+���H�\�8U�-�Dj7��^���I���.r��bVg�y����j<>�p쬲Y�p�$V���D��m�t�j�����c�X�P���k���`�b:ȃ�]�^pU�%w|��z�z�_.JM-��[��|ز.��H]#�<�����Ku[�xɛ�H���Bɘ���2�fZ�Ǯo��V�FY#=[��ntTGt���{N2OEC�>�'�%;�ᷣ�sb"���W��G8 ��:��Q��x���BHV���]��nazٓ���Î�i�|��ɰ�Z2��5F�����[B�B �۽��1d�2=�\�uz���'L7J �K�gQ#g�z�Zcoʱ�	��V�3Q L���N~�Bf��cVגߺQ�`l�D'Z6}5x]_K(p�k���ˬ�6jĆjw&Z׼�$�kG.� ����H�2ޕ�ҷ�tׂ�}k�/j�T��3�����g�r����_��{�kS��T�C��{����.�i�t�~�bo�ϕA7��Q;�u�ZN�4�t:���Z��)�/��8x�P`ܶfS��O�q=Y���/�u7�{�}:�ו���͜�N	䭞�p�o �W�6;Ԛ�2WNfBzS��[�o��]�ݽ;;6كwӧ��)@�V�,��K�)%�������l��"|E+��J
i�_�%�{�bO�]��wo�{�ƙּg�	�U��-�uYx)WR����4���}�f�T��ݪwZ>�,����Vo��:�U�-�*��8�M-�[�J����~ܜ�Ev��Ov���ťb�P(��j#��ɡ�^��Ŀ�V��m���4)P�N��_S���M�/yv��`9X���6g=��*��oP�	�c����Q�s��L��'����S�L:K�����VM_p�z.�V�b���G;i^��Ge���u޾�t�9��,�YL*΍�n#�f4j9x��n��QDt`��O;6�����m�o�rf�m&`���\�|��O�$��a�*bɕ����L4�y�ݧ+��s��׬�e�D�#Ǹ�^�4���V.w��<�qP�Y��1vy)���{�S!'�5��}6�A^���XD*�GIuIp�E��x:��[Ӫ���Œ�`y:x���ٯ�WS_��}�.�`��ё؜�`�vz�Uґ���Rip��b�<�0�:j���/��^ڝ��*��/��"�`���q7=�'��J�����q���bb��<����p�~K�}�l0���;,��Ѝa�L�}(�9�b�z׍t���oØ�E�����>s��Hw��P��.,�W�?|�-+]@Qߞǈ�P�<ɞ�)�kڰ��ji��^�f��p���3v6z��fUC�z�!`f݆r�[��}�c�3�ײ�X=6��~mK�^wgY��5��+ag��S(;���_j�0�''���ߨ+8+�~�s�W_�d�����k�:S��w9����=��l8|��3��A�ھ�4����D���� .
n.�erf6f)V�̊�3�Aw}�o�
��>�����m�&��d�A�����w=M�p�Xnz��1���ye{����k�ͳ��)���ӭ�N��k[�H�,��Js�v����WL#�����$��Nλ���Ln%�F-L�ѴnwHg��mr��UW�w�a��=t�"�(W
V]#l�R��\]C��vG��ֈ;~��w���=�K=.a9�'�u��jk�}�;���Zh3�$���~�uxߌ��혘˗z��1P���F_��4�\�e��^�]���H�r�;~� {.,���n�P3�������wc��KO�fo����=����(oz�)�cyofN�j�랼C{�7ntC��
��� �g�!���A��/�����z����Zn_e��Ϣ:��S����3�v`x�=WK�9K�I���A2(_��^��W�k�5�{u&	�y�W�|^�g/	ꘅ�jZߥ�Xx��y�y/N�w�p��P%�8������:KL�{�K�g��gx���P�V>���B����u�Z��·&�3�kl7|���m�0y�/W]�{Ն�EV�.�Pö%ݑ�P��'��s�.�~��I�)kR�]�g׵�ouq��+�$Tp��N_��n�� ��9u@�TA�{�M$ښ+�h��1��f	�uvwΫ_d�,�����;�Y�QܰѠ_�����y�{�B�\���ݢqN�,�����oM��r�+3��d+����q�Ľ��o���f��e/.�Sr��^h�rVN�^�Tɨ�Վ�J֘���ٜx`�3Y�Cm4|6�]8�:�ב{��؆oK�k�¿��0n�z��젭���/�Է�uЅ��Z�����!A�P��<%��LK���ǐ���,#e:���f]�7�vN��89��%�ҽ�	^(1�?)��g��Yy�������*�Y�Z}��>��x�D{�e�̒�χ��P�G1�ܕ��E�ZwҸ��+�L�+�:��uJ��Y����z��՞{Ti=�f'.϶;U_�{q?�~�C����Gd�]�rV{�>�@�R����`�S-f�f'S�=�c�>���v�w�!�Jsӥ�Gλ��4b�\wV��P�=LP�	���&�Ϟ�,�:�.V�U�+]�ٗ��|�z�s��/��>KÂ�u!�:=�Z=>i
֗h.��񚽲�Pe�^��9��M�k���0����A���V;%��`'H�ǋ�h&e��켪�7�B"KS�ƽ�z��mV�ͨ\�<���z��b�\'R"J���к�x(S3��p��=�oy���V�IعU��R��sV����Ո�༴nĢ\V��������ꞵ�zfh�{=05n������ؤ̛�<��{�;������ME������\I|S��胡���
ʷ��j�j���,�W�6�4��n�3�.��e�鶺H�b%y��L�f�w���Xt�wzs�~��LH�p��y<	Xpx�r�S��Ӭ�+�B��\�6��9k����5Sa�G�\;����*�]���q���_����$A]Jb�k�.��~�L؋�aJw��{�x�x]�g��u�����p�<��t��ݎ>�o3�	����t-�R�ᮮd�׺ǌ�f�R%׼���@���	����3�}�-�x��ID��t�oԼ�u0�Ş��e}Mۃoʱ� ��o��I�Ź&w�S����aGA��V5�tGWl�e~�����������6�,��8!�u�Gn��ǘ��������.��0�~w	"ÙoJ�J�]<�W��(q��Xl�3���:l��3n{�)Z=P�?Y=��U�8v_�ςqYӞq�>�C�Z#�=�<�T�3q�7���;��/�]z,N������타�ؠ�7-���b���z�z;�m�
3����nlls��2��=��-�X{j�����J�P`�z�Qg��q'.���Ľy�=p;�y<ʑ��l�N<��]�#Ђ�"��8s�����.���Y3���װW�J����h�:����������Pr����X��Hse���U%m�y���;�{��Ry:�_y'9�$.B�tJ׾�n�D'���EOaB=��R,]��F�
{���|���f���=>K�I��~`=> ]m�;��6y0��A6=o�u�>E�]�;�ڼ�L�^zP��P-PKRؗ*/E��?69��U�b�Xw��v�O#.��wi6�>�H�~��x%	μ}8�����2���Z	;�}">����u���g��q��~X����h���&�<�\yV��m���4*��^v�UN��}ލ�@ϒƢGuԡZ�(�����s��̕1c��r�繮��-W�Ɨ��;�'�Dϻih��
+ƃ9�|�s�u��ڃ���ꙺ���=���ӓ;�����8����h�W��𞰈[�t��
�]
����[Ӫ�Up��!�� �7��ט�],���WcN}Z1�^�+���J��J�"6��yh��ᬰ�-����Zk ���L�<L���]$$P�j��4��>Neؚ��P�^/T�>ѩ!���r��U�[y���l�5�XdZf-�TWk�J��F��)p|@�޷)O�ٳ]u��Fʠ`W���R��j����;��i3�3tź�����
R�+�P{�~UXϣi�;^�UxJz���]��kV����bt_�����n*4�PO��:u��^�=�!I��~�,�y%�s^�OeJ�y#��_�\�"����2�o��{�Gi����>�k��'Ʋ�*|c�{�购uGC��y=K>�d���WX�{_MN��5��c�����Д93o"�v�~��ǆ�E�Js��>��+�֙�7wz9��y�4N:,`�o-:�����Uᒒᄹ���m����8m����Z�nE�ީ�m�LE��`�}����A�Pu���蕌�U.X��T�{�_M�8I�w�iص����^8I���N^���B]��K���u�2+��z�R��x^��R~����&%CՊ�	��% ��������8��P�s��r��  �Cc�g����$�Νƙ3�h7�|7�JiX��N�e��a�zo@u�]X��·؅�y�(:ok�h����du���ܻ�rZ�fo�b0؞�e���$�Q���=W�]�>nv�}ǰ���<s�f�q,��P��g� Zv2���i<��xr��������m���/b���cd����ف8Z[�ǸT#�6�cW�Z���+���Q�Q
���+�DTA_�"�
��ED�"* ���TA_�����"�
��Wb* �����* ��QȊ�+��TA_�"�
��W��������1AY&SYK�o x_�rYc��=�ݐ?���a��H�B�a�@d(�$h��@ ,� � Y�Ҁi�lk@@�Ei�-�PaP����&[f6،�mM���X�e��X[L�kLU�j���3b��mV�2�[Pլ�)mU
ۮ�m�4��3gy�*�Vҭ��mZ�֥&�ɒ�mi,���ĭ5m6�mEZٱ*�Y�U�Z�i��Tda1��-YD����U�V���  9�5��=k�D���qZ5�s�髲�p�t=f��عv�t�Y޼=���Ӹ��Z���Z��kίm*�\���3��j��h/  =�@5T��v��;wwb:����q�ʅ��9٠4��-[{j��{���^�{D{v�c��w;��Zg��Hݹ��C��g�p��S4�  �S� �(_��  P
 �U�E�
 �� z  �(�מ�Q@(P {�{���Z��]�ST���;���=���ֵ��څ�݄Ƭ��[��f+%�� w������U���K��{w�^ս��n�5��R)��U��mskX��m;w���X�Z^��c�;���Sjʳ-���tI�-�  m�@w2�\�UT=jy^�vx�z�ת��Z��뇵��x�cz��U[�OOE=]�v��G���3��Օ�wf	�l�v�ZV���^  �`�e[��v�ѧ�������;q�����A�N��+]-r� ����7�k�խ�"�hm�+fM/  �Z-6�ZC�k t�s��4�
��N���t��9v` 'v�V�dʳ2��f��x  ww� ��D�r�Jc������N���A%��;�T���.� �K:�܀٥M�61���1�  �킱� s�@v������ݎc�f��S�«Tܺp n〠L�Vf�Z��6�[<  '��Հ�j� s����%�ƀiӒ��3��A�S��    �T���!�   )�)QU &�     �{LF�R� �	�0 M4� F��%T���0   & J&���Hђh�jd�d��2A&�I�*UCL20�M2`#d��	Ǉ_�v�g�i)V�i\䆐�z�(Vi�L��YL�Z�-�("�ko�KOH ��~0h�tTU,*"*U�@R��~��?~�\?�����
@���("�pZ$
�V@s�("� us�E?+ݰN=�of��@EH/�Jލ?M�z�!�#�����B�$��6�Im��%i�bi�2�h�[�M��ǖi������su�R�-MX� Zz�jۈB�:ŰMlQgK)����*���ǣq�{�Qd�Lf�C1��ڳ�>+�)�m�
�W7�r�pM��s	Q����U�ä���v��e�&�Mc�:ݺ˸�-A�h� G5M zJ.f셲,�!t������N�ZW��X�/
�Wm+�-X�t��m��iê�$�pv�Y����;���ف^���u�h5�Z�K���� ˏ���F(����Z�v��Y��e�])5z3*5���
�gm��Z.�ހx���U�v�5
��/
��̭aͭ̊L!$�,Pc���lv��Os2�!��m43 Ů��f�n�C�Κ��ԯkse]��b��3�B�4���e$7�OK��8X9!n���c\C�Yem�*[��ԑ�,���Cv��9�M`(O[�,R��Ķ��까�_^����\����aV�4������4��s��.���R�AN���@-�{�QQn��m}ͼ�/mf�yA��v-" 2�f�+�.c���T9��i��.�C��h��Z!h��a���yƱu`��M�Y��H.�l�g��6�+_We}vۮC�	W3�I�i̊J+RЦ[)�i�Q
�ٿT�H�L�w@���J۹�.�^ұ�
ů�Q��F)L(r
�Չ�� �������藴�5�nU�b��䥝���]F}��h��&+R�u�f!
ˢ�H	w7XԹ<�l��
՛J�ƽ�P��J�1�J��3mebGNU�$ʓq���<��J(�(@*��@�XGh���:!���������N��A��ǖ���nT_ ��-W���5�e�����St��m�Q��t^a��f*��#>ل�h�sE3���vCt�w�ݠ�f*�YA��q�]��y�ר�����i�犉ql�o��e���A+m���=�u�TsCe;ED�BZ����Oq�[j�0(@�
�7t���o[�q�5h�T*�
ѕ����y����T�$s�Q����>ǫ0ݛ��K�����VU�}��*�ѫ�]��u�\q:b��ë*|uХO+�6hͲ��XLC���5Җ�r^TV^��W��͔t7�6]l&o��Z�IcTw;R֙��wx���۱n�X�غ����4 ĥa������ah'(�͉Y�QZ%7wy#D�r��7h���`�Y*�����J�i�i�C53Z�������̤-.�u#JQ�1��*9R��Ӎ-ۨ�;����Cr
z��k!b���ж7zXOC�v����v�=���ʞ"��t��1ĄN^���V��un�
W�X�Z��-p��ܬܬ+%*w�`�o5���Ќ1V�&0���$u1�]dI`�R��2��H�:y��[fݶ�5�V&���C���ΐ��q];q�ȷP9�e��M@�cU�09`��]�Y2�Z+p��ow+rT�m��H�j���?B4����xoE�:K�����$0�����@�#j˲Y�$�tVm��@�ى�V��0��U��Qm ����ߋõkMY���K4�*	caZ-$�-䯴�V�m'����s�XxE��	���.Í���aX�6y�X�+5�")4S���SwW����N��t.f�ز�2�F3.����p��5@8I����	u*I���ٌ��/�Iַ�I2V9Pѿ�yw�kl��`�1EW��f){��kVބ�]�˵w���4�J��{�޻Y�S�q%�G)�^5��a��Q��YP����Gd
�!xlj��\bɃ*i C��7�@TTa�n^��-^]$��E�)�0!�y�#f�G/R55�to-:����۷�����-�Q��Z{,fY��Ʈ�Y55G��T�ܹdmk�
�	�*tn A��rm�{.3��.;�,�[�+h�w��B�hb�ll�s"�XJ �e�uwFC%)�
Y���[��٦,r�U�ɹ�
w�ѤV�h9�-�O�̬:�mP��}��I� n+Չ�'�V-O�fw:ۥ�iG��RE&_1�+(ڥp}����#�r��m&���ҥ�����S�eƥ��2�E��b�w���,.��,0eh`�m$7f�� �CB�}A�	�7��D���a
�n���k,5�Z��Ƭ	�Bm`eR�OF��e����L�T�Ւb�J��jj�w���E恘U!��+]J���kĭE/k\�����j�c[p�/�F^��je"�ܽ])���&�7�	�F��t�bͤK5�Y�nV��)��=�-8w �(C\	1x�V��4�T���s>�֨��kJ�;R,+�V����׋�m=/PSD���+&��^KX�v��R���96#쑴r��w�����������i��m�GcX�=ˡ�8�jM{�m��X�0��.����R�R��2�J��FƆ4L���,�h&�\�4D��H�����V[�˭x� hhPPW1��̦�+Y�oX��c��&�q&�t.[J�ܭEЏ*��6n����v��e�a�y���)Z�CbN�Vr�ذ�A{u����Ϟ��U� �Or��隣�Uu
�y6��W�Y(���B��SC�H�(MɆ�Zb��+!�l*KMm<��%U��c�	�b|�5�^"F�`D��:��u�z֞�8Gv-T�v<eR�c��wԍ�4XJ�f]�5�[�#��M���)VCM*�k���F��]���]H������RAn��Xt�T��	j�ז�ain��Esv�-�4�UI��֙�+nK#��WX]�Ig̽�o��k2���ۣ�k�B'b���z�hJ����F$t�f@�P$v;/*���yj��6Nַԏs�\��aأ��_`�t�0�#m���wGnXT.�&�����1�u�a«d2f��x�`�*�@L���*V�s[*Ϊ�K�v��f$�a�3P�k֮�M]�;,�Zy�i`�;�{���ǳ5�^��Z�K3pni�� %n��Վ��м�.R��d�a�"�E^�c�d'{yC
�{�ʵ��en��˱�MX�]n�4�tK�9��Q���t��,���	�i��qɹ���k�vm�-T���Ԕ	�+YD�n)Y��
�����D��V��r�7wB�1�D���ge�5����ʐ�̣Ek���X2�-��(�y�HN;R�̖�17���ǎ�+��Vd�l��l�3��Y�4J��]^QO�Ou՚��F�>I.��,�Xo�{|��s�W�1M��l�@Q�3K0+��4�2�Ju5�4>��!������eݱ7��r�X��=�ha�2V��j�Q�Ԃ�NE�/��z�0J<�nƵAr��
 5يK(md[������uZ���|5��U��뼤Qv��ǉ��Z��:�
ʼ�`2n�V:�lW���[ۨ�ZY�-m8�^��+*��4֖�m^�&��a��^lcmщ賆Xf웑V������U�F�*P����-�t�g1�(�ʼͫ,���UD�.j$���׀��1��`S�,ɨ�CWF�:��]'r�J/���wRa��ו. �P�����u�0���[��[r�zLд�2uz��j��3iݺ��r^k��kV�qѬ��a!-�����5]�P'WX��T���yw�v.�2�^��m�2��3X�LP�=�1"�Z+sa'E������i��V��BҖ0AA��2���Rf��\`�[rR�1��D��1�7h�̐
���k�Oj"���wCk7�Q����&�:�4�)�W�#e��,�i@�v���;ȯ-����5��R�0F��2��ֵV2�Q���o7&��y��b�ֹ+%���i���FM�K�D�uh�0���n(]��6RYKM�WA��hd�\�[�AڤUL��Cj��C4�]#��6Rn$`�-d%{�f�[���$��ϘU�>��^v��M�vUw5G�4t�����QK�][�]��pV�W�r�^��F3-md4��&ѩ� ��Ǜ���K�	�R��`۹���K)ꔳ����S,�˔��Fjvw��Z���j����i��Q�5��j�qlO�ơ܏��f�)��su��H�o-ZAP��/[[�ێ�`܎<�^��
 ��M�ە���{MZV;�zl9v�K�&(7e����G,!/awr2lB6$�uj�Hp�mibj�m���u�u��lʘ�@�v/)n�Z[ܧHe���E�!Du��Ǆ�/�k�;�A��)���'.�TP�E�`�����A��܎��M����5��3 .�bזx>*����:B�����.�8�IU��D�7�Ӂ��Ks[t#���4ཤ!A��0�t5вNgf�a��g�v��t�>I�T>�#u��Ӳ(����Nj�)�
KU�qP��t�C����P�;j����P8���U�]w"�â�m#x�hbY`���u���'Տ�x]Zn�Ǹ��	 l�*=�
���CCXqV�M����?�TFc��m"��'t�#xaX啖����eGN���-iʀj��0n���[Y+!ݫ��)��4>/ �h�Ѝ w��O"/EX�/�gTui�]���<�w�d����T�j���Ӭ�f����r���tM�"�A��Q�r�U�EkGZ��%%{5����oM�h�)9�<��t�T����ջ�`�9[tp�=��8l5qH�n�� �Y9����eBM�)����f�v0i4Yy���L�l`�U�g���<$]oC�<�)b��TV6��O�Oln�ΏP�����2��+`�_N�t:L++��p����I�h�/m�-��-4�+���� �b��Ѷ��$ټ�öl��V�Yxt��t9s1�롹P\�`��eZ�b`w����[R��xe�����Z�L�f�ݒ��W�� 6�]��N%� r����N�\�Or�� R�0���P�F�hL*V��Ft��K��I��n5Yu���)�*�+M��R�uq��kz�:��B��ۂC�Fq���p�l��Z2�� �6�r����Qd��`Y�q	���\7+�#���U�u�4�b� E���ͷ����e�r�Ӡ�͝ڰ�9�sBi�d4mVa*Д1;וr�%�d���ܗ�����2�s�c��==��-��jCp7Lh�$<+�����[���/i$��hWʊ
��x�6Z�W�C��,%`4���`ޛ����TYk�V�V�P��u�VVvtU *��v��CG���e5���O^ЭPM�������mR�N�V!�*q�\���-�xX���Mcr؎e�۬�&_˵�58�9�p.S$䤬����@��38�X�^����1p֖*����9Bvq��R�����V�_ǧru�R7L�ܩ�݋)���yBA�K<ml&�.v�(�W�Cm��1׆oU��-2
�2݉�/�"�-�<k6��MLHI��3��<���L�+x��M�7Զ�}���(���>9�c��S�:��<��:{1%OcC2^Mܣ�+h`�el���yZ�ݐ���.bo���ђ�)�vr Ò�D����iZ����ہ1�r�x��#�T�V�8�/�_�+���9^�}�}�Wč��nmE����^�Xe��vm����|�݉K���4�ZݱP�t�^�f	���'���C8�.���dn��9c]ϓUú��ڰx�0*:���k�XqBhC"�c�6�����7��iV(�W@�2,���ľ<�[E'iX��Zr���ahJ��Ǫ4�&��Q�\��'(\��6p���ʼ4*��TKT&Uظ:��/1�6r�mL�6��*Xti|"�
�)��yϋf=g��!����w�e�b��r���hP���{M��y�ۺ����R����Ff/V���$h4��~�]�T�F�*M�+�G��*pܫ4��i�ͅ-�y�([�VA�םw%
;�j���F��%Έ=|VM%1���)M�G|�&o�:��*���1KpkIut�6�Zb���OA炮b	ωȆ^ͫйKiv���ڀ�һ�����x�o܃V��I6��ܣ���=[CwZ���_B��4����9��*e*�A x�mK\���M���*�B2D��rn7�a][Y.�v��A,���iŸ��4��5Z�b�z]�Xɝ-v���E���U�ũ���f�(��f+݅�b���e8��ڴ#��3��uwy&�IV����n,p���2��0��&̇�<ZBv��V%_��Mu��ڽ���ifb��Q��e��<���Ni�Y�������
x�����m��㠩�r'k`�No�܆kU�0�Qo3�U�����a[֖�P���MtG/���_v=!�,��QF�suVK*�NK���Y��\ulk���1�k�h_a�uh��u^m�B���	�fY�/Z�V���Fn.⹈�8��R��<]��Y��B������*����eb��݉Y[�6)��R�u�1\O �S�wv�y)��X��ڏCT9�׳�ə��Eغ"�	�kG�KἮ�k��wGe�ǧ��8rԺ��d	}>r��*΍��4U�3k^�b�M^婥��n�qfI}��|]�4�K7�WNX�ІM����Gz�*t�Ut���r:>�fE�v���.�`ͭ�|'b�ދ�Q��|�5�4�9�c�Ȼ{u�0Ta�t�ަ���1d{\�%g�K���ɖ�Z	�Գ��t��#�i[�w���A�P�cJ�;���\��r��@�fto6�@�i^��Fʂ�&�9r��*]���T�qKcTQn�!Y�{�s�L����F��_k��P���3T��uEX�aRM�-��X�Y��N��`�����-V��u���zN��Q+e3xQ;>VF��r��{����&-NU��I��S�6�R���J�P;��S���pZ\���`O�Z�y�I1֌Z��Y���dWSU��Q8?\��;�Yu��Nݤ�J�D�OE"�ٛvz���X\ٵ�U.S��r���h� Z$,/x�}������W;:t+=�ę���@!
���r���j�o=���V×�j{����+',V�\���z�92��'�pB���3���n e^�x�ӏ)�E,=\���E On�"<�3U�!�e�-WJ��Ґ�̤��Z���N��qw�kn�c���;V0����H�u�����꥕��,V�k&�d2i�Ǩ.Y{33,�{@�y9/s����ϻ����t�8B��k��Q}�fqy�������7U�gxg+���x�*��H�&XW�/�Wk��������VD����n�<М�r�+H�֙͆d���H kR�v��e������!�;��{��WV_'))(�*��n�/�u�4xH��euN\�
k�YNw<Y`1k �e�Ū�I���)8�<��4�t�NqaI�8���T��hwZź���c��o�����`���W6�.M�4�"��,R�U���Է(�:�Vj�ջ�^�'O��Rѽr������L�����d�7�@�eZ�"�b�Uɧّܘ�C�i ��c2�n��t&��fJ�I�c̝g�e��6�'���t wB��*�Wrq���3�bn�aK��{,:v7��o"TON�� M�:0��E�/L��s�2�B@.ܥa�r��3�k#X�2��W)�e+A��NXG����Ě�2m�P.),�C��Ҵgi���$���v�	���L��d
�uL�5	�Kיa��颴>�ct�D����]W�
��	QԲ�哰�Ţ73����SiS�Z�Z��,�M_V�
�u���u��zQ�v�S�ʚ֬��3�"!��^-A1�����8�z[�VHt$3UK(����@b-���g݌;Œ��L�K��-ݩwoL,5Y�v�K����P�o%y���F�t�	X8�I�)�f��� Xo���)>����挥Eq�)bk�j�=p�A� 6��(5u�7�b��F�ĵu��v�3"�(�j��wP�A� ݯ[Πt��rc���l璹Ւ�$�tۉ��Ұ����3�У�^����|'<��v��[gʲV!Õ�����]83ɣ�]�r�J;}@T4�_#Fn了��B��w��4WVk��7��7Vxf�>��Q8T�D<��Y��2���Vɒ���5ybA)ʩ[��7�]vFc��C�Z��PFm*r���˕��dW�����nm�1��I34��[һ^>>ǽ���J�[�b�d��U��{�4	�f�ŗ(��ŭ&݅\���� ,�[E��JK��4_
=���A��|�����0.��,u�M�6-��l�d�$.�A�;����w3*͛�5L7��sp�����a���@���#Y��ʘ�i�j��,�YN܀e�$w"8TY�˚��v�v�F�)eڮ^=6�.�#�FH�fa�����ƒ���K�I����y%s)a{3�G`ܨ{��7;�7��so�7��e^�si����x���
=]	r�ܬ-2�u+���o��j�(؁Pq��q��mj���ˤ5�+*K���	���UY:V��L��'7���e��y%%1af\�VW�M��a�(v���qqr�[2q7wo\�TY�B^��Av�"��ؑ���g��kr6�,��T�	�;
γ\7���0�-FW$�бۈ��w*M�)7V�ש��8^�<��)��j�����A�}!�� ����ӵ5]z��F�+կ�QÎ��G
�N�EM5.���l��4������ 9�cy9�gv|�Z�#�"�5(�$"&�쑹�7��im)a�1iV�<�֓0 ����=�"ݴ�����f�3#���r*�������Yѡ�JG�ʯ�����{Bu F6���:�;�<kd��WQKz�)�ьƯC�n��#�5����)%�p=�ݓ������m��d�ԈBK��w���4����7	9%z���쫼Mln &��8��3i�uw( Y�}h۫C����Ħ� ��[�Y�P�+�2�[�gt.stJ(��`$DP{x��['c�kT�+�HIЬ�hJ{����X]+o�2�z����r�Y��MC@�{3�S�C����n'�0��w�2�_ue ����u(�A�V{�a�oA�r�y+3T]3l'��	d6B5�c���Dm�!���J����:Ov ��@Mki=��hiZ����D��f'�;�X���ɂ Nɩ��V��J�m���	�93�hZ�����0�?�Ia�Z�G�"��
��]���'%��m+�w�Y@�O���Rfs@�R�Z��I��,�{cz( ���T�[�ES��ȸ�E���^h��tC�.+��\�����O�4��^�u��v+s�Ʋ�_.�e
�e/�K�g_Z6��=ie �nS�%�dR�z���|k���:CPjkP��*式v[(��%\���T�jm``�;���Z���2��#%x	ƥ�O����%�����!8er�sGsY��RKw:=Ev���:-H�uT릸�a�q����
{�h][*շ���둊҃X���<kSRg��mn�znU���hu�Vu���*Pλ�5z�$Ljڐ�!�0kS��L�%�#���P�f5�J�
�,�X;� �vP��,Q�*�6��NEwtX���ʛ�%���[x0=qe4\�{uU��BN��>O,�o�dȂ�M��By��3H֩�KQF�T�)d�0�C�B�����r��ͮ/U�Ur�rFR<)J�Y������/{��) �n��]b��R�P�x�[쁊��Ѹ����6���B����B�Y�L�:�5��֮Wc���:	ۼ�b�k�/��0��U�ww�d۴��R����&�r`YΤQpu���K3{rthZ�#���VE�$��\s2�)J�l%J�Ax�7>'Av����X)��� \�����v�$T�c3W+lH�d�]�ܦ��D���hfb*�d=+e�yf؜E/qg�z�jU��\MX;JQ�ݣyX�e-��xKْ����nm*�Z�P��{p�%��yW�;w�����j�Y�foB(����O}��G�s�<��F�N���H��}WvM����xFƣ�+�T���޺�.q�@�[��g��LkSk2�12�\�X��뛲�� E��VVǒ�ұn�P�|����jq�Nl���f�s!�z�\IU�ѳ�k�Bʸ�y���e��
Tv�����"�W���⳰���L���V��)����@�Kw�9�HΥ�-�W`ֻǹaǒe�6��TE�Ɖ-��6��A���W���Z�r���d�a��g ĵ2\#v6�7��^Bg*����Q�#�yR��a���̇ �5ܣ����i�,�0�7�݃����Y5��	UF_gta[3�_��?`���k��_�7lHl�s�����T:�3�hUDT�L���w�֬��6☹�zw�r�e=5��,�p�:�{b*���63�%e�s1�
%�ʖ�6b�G�\ ���'NF��y�+�Q�5��9"�.�\��˖^.�%�2X��^|�Wv��;����L���<@�}��!�5�`+�.mL�i�O�]�Sn�U��@E͵Dq �v$/����3��_;�r�z�=�!��KQ�Y;�W]ZC�We=9����Py���,�t�EN���n-�w���&�,�g�
.�����քܩ�f�����;�x
=t��޻�Z���O2����6�db��L����ڏIt�u�SyL���"��X�1Rx.���������kúmp�LD�Gs/EN\͜���X���B�H��U���%]i�5r����.uHm���hac#��{
��2���VSӫ���]�G���s��\�]��2�K m.љ��x��¾je^��4�8�%�8v}��ňWg7�y}t�ո��8���b�ۖI�8��wH%�������u����r5m ���t��)���\lE�!�.N�B�bJ\�롹�`��Gw>7u���.�7u�R�W4�]�i�����{�S�RN�-�t��}.�,��.�X7���(1��}c,L��K��]Q�53��;����w����(��7d�F�4�b�gQ��r8z�K��՗X�h��e��Nw_
��u�:�b�4�Ku�6r��Y�!��nhcR���(:�wX��u���oqΡSq[��1�dS�����������zf��}f*1�w_L�����Ģ\ A�]�K�"�HՄ���קۼViI`I���++�Nx.�e<�QJ���:Υ�&^���#,�ԩ��%e.���z�O{,2R�5�&�}G+;	�C����#�ܝ�J�|��[a��/3���%��zH�(�a��Ħ_]m&��,:05�zs9�<�5=�"�-gMU�@�R�oM!����߱\u*[]y�ꮢ^���[r����֌Z���4��me��,�U(֋뢥����)O�E9S9��C)0Yx��mp��D�d�w&m፾ �fM�jݥK�b��awEg��s�
�ޭgM!.�6L.�����f^i�EcϷ��C�n�-l�9[x�_
	
rD˺^�����Հ1F�h«�ܜS;.�칬�vX�/5r�AL�za��m��ۛO3�7�
A)@eeA��ن��1
궧�{��P��h���d��:�K,U��Z������
��02T��6��Ԗ�)t�^�ᘺ���L���On#��a��� L-�T5Q�5�&7N��vbȨI%�;���j��������ɮ�7������Ǖ�.H\{:8� �5�w�u5u���-B%�v�E�vV�S9^4+�ɂ^�F[6�ä�^��r�1X��|���ʳdp��N7Ɨ,�z�)|�Ķ"�D�u ����)���5kV��Vv��h����Q�0T���"��\��Y����؆����_fc�
ш�6u+���W;zWZ�C��}�:�C�O,����6;���bhb��(��I�Qu�7dv,�g��T`��k;#^X�����o>SR�[���+*����n��'a�Bä,%�|ia*f���u��r��
����K�AmԽ�7&�o�^f�6󍶵u�[Iլ4� �)V��'|7e�|���;`��הYX�] ���W�Z��{\� �=�],��V5�!�R�T�.���8�ڧE�!wR��0�_-������(�.�3N����T��NH��A���f�$�!�=U�$ �ʛA97�U��m�+�־��N�)��mf����m��_�pM��pռ\��8K�9i�$�f�s�����u���X�b8�BV��t2�cX�n��-R櫯�st�/��l7Q|^�Ȓi��f�4&e�M|.]@n�+k-:��fo��ۜl�F(�u��f�dēu�3:�#��'�Tr+�Xkm$�봕x{fY�H%Wʵ����w�ћ@�8�։6GON<��-7���B���2��Rb���$�l٨�;�OK�3�W�5�����:2a11� r�2N��|�&̵�K2Z��R�i=��}�&�rvXɮ�⛗zA+h;Jr�����rKBn���)rdr�k+��uL���߂��k�7�ɶ;%t���D�g���cU�#d7���kho�g��� M��L��Ce���0��*vőY�HK�V]�p��_S��ĳ>N�K����v��f	����i�X:6��2�l^��o�V�$+.�z��JH��Hw]C���8�,6,��:l��B�X�L�/�ld|R���
&ŷ��2�b������ԩ��[���1��7�FNj,�����l��L��g'�;e�C~̭2�7 a4T5KA/L��rƋ�Uث"���T��ɋ^�XR���©m��#�(U*��fu�'J�t+w���#�.��E�l4�V�[Mi[9*5���]���]�$E���v�����(9��>��sh�t]F���utz��(�"���Ӣ�*�������
�+��a����:�W�
���)�Sw���9>�mSZyV�!��Ǳ�5%�G�����N����Xw��U�W�7�"�6.���Pv`��r��I\�WҡǬ;Io#�k��w�>,�����r�WB4/�����%�L2��ங�I��:�SbTRir�J���0��rt�
�O��}�t��֫�V�fv-��w�,&�F���}����ݺ�X)�/�#D�U/F�� B�Yj�}�"���v���6٩��0+l�s���J^G�6���RS��L[�E�^��w-]�8q�՚�X�M*��
�=Xo��N�O�pR�v� ��2!��Nث��"T�e���v����l0�Y����)�����]Յ�U�h<���H��I��b]�-bW�cw�c��K���;L˫1c��_0e��gU���*�	�4�#��,�U��_U�(_B�sn��A].��m�U�OZ鵸���KXf�$���e�]�VOcXE�sq���к�qW��IK��:�=؁[)�R%}�u65a�Y��U��Q�yZ@�L`�
B�э�n�]�չ��u-�Й'-[R�k��r�rۋ�K�B19Q�NoX�Q˧�& ��0�S-�V����v�iT��t�vfP��3ۖ���5q�Y\�`�x���S3$�Y�[/N@e�t\��fZ��)���s�`a��a��z��8A��N�봳>TqQ�V��x>#���;�t��Dj���k��5�X4�.RQ�s�\��Z�0Y�����������3)1���n0h�fV��f܇�\��V&ʐ��1؈��&�N��bk�'��O)A���Ykt�u8c��H;E`GA��R�־tr�e]���J�ǚ�g8]��$,:d�3r�Elg���,�!2�8쥌�-gQzN�nҵ�c,Ge<4��P���G ��At�^v�#�-��[F�w2AJoZ��� �ܢr������[��lN����!p���ʆ�i�FL{N�J1ͤ�U�7�w�t��1�j�X��֛��ͷF��J����b�8:�"�v�+iT��c�˭�!�>�0�lV�j�Wf�a��Rp�*V&�K�z��D7�p\���Z�݊��Z.���ȳV�@l��Mmh��q	*@9-�"�-����BV1��P��(���7h�q	�@Ӆ2��ob���i��PTrٸ�T�D�Ӝ8j���4/5�9���I.׳˵K�9�MV�����Q�;T;B4t���ڱ�����5TUn5%ӊ�^��-�8r�����;��8�sw/��7���F9R��+F>�����S˝|j��K�mH�X�.�Zɣ586�F�Rs �"�K�[�Q��3��Y��bJ)�uҕ
�|5S�kf��*�xJ�a��4��+lgX
��gR�Pv��V���ed�|����Yuѓ��x�+ I=�J�3BL�W8%z�u�,:	�����Z��ޢ�Y����kt+q��Y��8�mJ1��[:�{�o�Q)��k����b���Pm��(�]��|�SS�����>�[gmW[JaN�Vc:(*�U�w��{�
�O��^Q�\9�Z[����Y�z���I;C��ҴH�$��=�t�G�fd]F���3Y��Uu�KVӔT��b��-t��ExU�����n�d���jޤ��\K���g�n=/qj��Gf�etw�1]���V��O��Av�� �Y��wl�����8	^�j�W$���I�"��5d�Z\�)H�*�@m����꼮U�f���[A�;�\�c/k�*ֹ�:X�uFQ�'*� v4p���>���l%]�� c-�5|��8�;5�гR�*��s6r�9���j�R�!�s�u���Ƞ�}Y�ث��/Tvb��d�+���d�q����i�脁s��}�w���]����"ƹR����*v��v�FnZnӚ�1�2�ƺ�7����QG�S�2���df�u�H�K�^��-��%��+	�r��6�|݇R���W'2��P�y�{�:�zn���%�Z=���.���;'@Q�����szҒ2������\:���!J�J�(SU��
;Y���i �B5����q��Ѹ�wW'�/]�b�U#ă8uX�Ȥ!2��n����ܓ5���`�����W��Ѭ�*�T��S+h_+/m�xGV���:ʁڇ���	�N�&�+=I+��"ށ��WZ�����&�RP�e�2�2v�Fc��v�-8����N�'/b�pt]p�yѰ�JD��Ŝ�S��U���Y�RN+�Owl�Mi/V�BR�;��[8ا���{]��I�*�9���6�>�JŬ���lT�aR����?]d<�.�.Ũg_^��Dup�p��(PY*�eO���{Eq�ۚ�;t���Q�;v�Ǚ	�o�V���ۂ�h�Rurk�iթ��aNNdP��$�-��C3��V��R�3V���襻�W�7���h�vF�k݉i�|�n�8S[@����:���b��V)� ]2�ov�n�f���yR�IV�7 �d�(c�@`�`��6��a���Z*�ܦ��Atlkq�ܱ��ً��o�:Q�3S.���h]�N�����.�@�2����P���Ҳ�i��T IOr �x~u
f|=ݫb��2w�3÷A���тn鬡I�]�Ÿkv��j�U�\�
l[zkb�ՆD��޲��@r�i�����'e��
�.�pυJۙ�q)N�1[�sH(��-�WwZO�T�wi�nG��+U����x�Ys��4��L	]$�in�0	x�J۫Q6E$t���b1;kA=�V��ۼݝNh�y^��m��r,�X*���V_�1˶��1v�2�[J,M&�AἻ�!��媕k5�4.�]�Y�m�.�A]�k�b]r���7؎I8b�]j{%)9gj��
R�q�f:�U��&�z9�Z	��b��  �K�y`�K+��b�f喤��A;4W:o��6�U�e�J��Vk�%n�����i��MCS6��\U��j."�_lR�V��������S�.|�:�g�LҬ�5�d�N"n򆘺�
��kUѐ�K�F��.���+(�Y2FȦa��ْ�Gc1]�
�33��ļ}��/�!t�N��X�6\��d`�.�c��&
W4h*\�~��fA��?����
�c�+r��A�Y�+.a�m���]jcS�+��l������Z�*kF"t�'[kT��+�PPvֵԬ[j��.!�V�SM(�%SZ(���*`�K�\��)r�ʸ��`�j,Wk�2�-2��CDSP�Y��M�&��1�����X�rܻ�ED�nj���q�f0Y�&Z5�h��1�0kPQ�U�f#�1��0JŶ���lF�v�p5(��)LED-L�er�.���Q��V�f�F-��LT�m֡��2-�;���U5�-�5*����R�¥E��]����a�i�O$���ϻμ��_oFuw�3T��+��9�N8o"�Ồ�b�ǃ-&�ev��)�z�b�����9��3�c��2�&��g�I3-~#��b�Ɓ5�.-��G��W�o~vIT�㎞�֏�]�w����I�6e����04� � к�%��B�a�9��.�z5�+��Ў@Ź]�oxQ�]R��*�YG,��.�¨��w���Y|P�����
s`l���ߒ5���P�ʈ��
�j�X����2��ޞlr����ڮ�c�����o�KW�|�@�֨*hK�)s�{^0���Te���t(�'"�|��P�Ҕ���]����g� ��z�)�J����7��Wj���>��^�K�\�����e�y��b�v��t.�<�����&y���M�l��g���vYS�ΎLŃR'�e����N֌B����[��<콢�8�e�n��i���<>wu�V�lZ��u��[������#�J^�/�q������7�pF�e^�ɕ��1s�Џ�?=� �����zN7� �q|B������J�\؏�#��w��4�6�^GI䇓<�� �
�x��[�q��ƚ9����Y�X����ja�q?v�I<����1 ���aϺ�W@��c#x�E}�	�0Z;�y�z�+�ٽYP���mJ�W Kn�g�46E+`Nʄd̨��+;#���W˓�&�D0��T��w�iyh��W�pVV�+B���Wz��y����Nl��6�
����*��+U*4r�"k�{UK�l�Z�����t$q�8��
���&;��.6� �t� ��V�@�ŵs8v�m�\�5�ޮj�ƺ��Pw�������G]Q����kf˭�z�G�u{#a���Z�]�@�9����`��HR���B;���+�|�Z���D)��#i�ce@�p4:���؆��D,Tl�Ԫ�;�!U�%�)E9�F�����>e��0Uo���9��ʽ��*��C�
;�GR��HX�dh�����q7���(���V�ۆ3����f8�e��ŋ��Ρ]6+���4��!X���j.�의�	I�)�E�'��w���Ty��-�!��ڸ�)�X
x�yA�L��ߺ�{ƨӋ<z-(��x{�SqW�x.4��՛Y�����Əz�z�j ��d_AТ`�Qv�S;��`�p	j9st��p����5�G�/��ʱ0��(L?E������[�d����\��vã]���)ݩAP�y}���&�p�u1�������{��8�����3���Y�?38�`�g��[]Rs���ۛZ[t�Z�j�`U���$��#�,����xL?L�h~G�U��ڔ!iC�JTc:Fj7Q t�8�MA1��bÒ��U����Jm����+���.Z0cjlF%	�G�@���� �a�����%	0|ܘ豓jC2;���a�1�\�ږ�LM($~�x�+W
��\�>��w5u�\����ve�1r+D@-
���x��(r�c�Mе�f�ݹ�:�PVr�]L�i�xև��:�@�:�����D]��+W2E^��G4��*d1R��o���bT��Î�R7�����BTiXQ�wY���;6�g�f����E�=��٬�u�L��SU/]��z�e�R�'/�������1�_<>T=����珮(%�gG��
X����Ye7t���c�b�#�����ݱ�2�\�E�_��:�<j�4TOdG\�t]�N�Q>�U�I��"��3뙅5�n�k�OE�[U�&�6G�0>7C�=���P?p]�|Wڠ|$޵}#Tgh��9�gK���٠�+K�2����P��[���>:xVDP�L��y��T���z��r���V�B7f���*}@�JnY�fa�<�B��^P$�ޛ#"���~'e�9좖U
��W��婵�p�\朱�D8qFE�T.f��b}FfR��O�z/��Up�Y�O�C�w.{owi��*>��+2����Y���[XB �%�3G0*�y�yP��+2#A ��5�j�d����;�&Wq�P˿�>D�{3�K�}�����t�1��s%i��xn��}��g^Q�n�,�p	(|��������X���}������Oz�S�pTA!���h
�u���%�]YJC�*U�Զ��W��:Z2-D�Һ}���M`¨����V�^��n�*j��6��˘�P��:<`��n�t�zV��d&�[��%uav5����i��zuLX:!تʏ`�F/�ՅSN{�����GFM�Y�~jP˭tr�?8-�Y�����{.x��>��_<)ǜ�Blj���P`��6�u��T��J�ÆwƎ��H��Z���ʠ��혽��O}=�Ct�M`�M�l��jVP�^7<ü{�B׻?wߛOƱ������h#>O��Θ�FoeE�^��ܨ����;r	�Q0�k����|��b�T9�5Boiǰ9
�T���_j����*�Z��Ⱥ���v �E C�:���_b&s�f����0�t�9��=[VCkq�òb��Jz.��A�ۗ8�ܐy��rF�{S�UeѧY.�:���v��	�Q���������΃��+��x�و�����R���O� WR��5�J���,q`l�gG�޼>�p���7)W�.��ٟ+_%�T����p�
ꁋ7nj��͇;��V5Ys�й��*��f6�y�گ`ʦ�⇶u�z]뭫�*z�+�׬.Ep����u�AR��GW�Izʞ��d0�@�d�#6B]�{��ኆT�9,*u�kie�Q�iTU�=r�Ų&�M���.\y6`�c#AU�Eu�`+:j#�3��j`�)�l5�^9T����.�:�Tk��4��T��8&�{Ֆr}��إ,�t�Wj���F��jS:+i�����Ш�{��M����éY:8*
�5<iݾ������xy�^�L�ӛ뛛��{�)��mK{N*try�oyN��)䧘y�9��e�_9���J���|��^��Y�������Q���X�t��ޜ���".L�.� Z�v]!��{�T̈BUs�����|�v��ʈ�nv�btoԒ��V��G�E�z=���կV-��W+�W+Kn{3IBI�ڑў��o�ux�)9*ME������_�¤�9��>$ݼ��&�`K��R��K�k.ãX���u!9��<BaF_f�����=Z������;O���~����n��7b�WlDÉ���jw����@n����� Zڊ��NI�����̎�]Ѡ������yK!���"�:�X����4*N��qx`,x��s`Ѡ�ϧ��v�K��T����ّDO�%Krnv{1X6�8�YS{כ����\>��^���UWG�����eJZ�|+5�*��-�Ԑ5�,907*�Ϣ���(m\l5'����V�QƦt=����m���5�<=J.�h����j�B��)A�j�W�R+Tfe�L��)�!�Qs�VT�z�cZ�TU=�S���Gq�^>7I:n��*���.٦�d��v'S�<�
��ae��p`�IrǕ^@��5����`��e���B��a¨����v���3̭�,��x�:�H�>6*;eҫ��j�ޚ�]�%"N� ����|h�uX�a�=�T�´:��<_B�n$n*��gI�J-�<�E�^�
�yB~��)R�H���_̬�~�9��<���:}�^}�Јwe�٘1�6TbP�v���UDEι���;�����"�}~���gH��R/�ьS�t�^Ę�P[�+�
y^X��ĮCO��#��OC�^���]M)I�q�jB�'yS~�L5z�V�◞��P�x��0G�_j�P$5T^Z�>U���Z�e�!�W����Kt�J3QA���oP�mxK�>���P>a��B5��#z{ws_ReE�N��	��b�#x�;K��T8�p�x��gjީ�SH��,Fz����땀ы�V�5�H��n��T�FΉc<�,G���z����҆���w���� W��^�1|$�X�kٔ|p���{��.>���񖽽u�b'�8Jܖ�ѕ�N�Y}XsenU`슢:�,�T	UطYݥZ���Pi�ݎ̕����
:*>�uf���SRʸ�#��4-K�U��B�lҺ&��6)~��]_/�qׅ'U���AZj�u��S���C\��(�7r�s�u��^{��vW�~�*U�`ܣ[��>z9t
���S��E�L��u�t+2�y�����[z��YBq���{/��9:�q*A�2�C��g*\Z�w���g�H��fmh��V����)�C���s�4����W ���>�ʗ�Է8.j��^�Ɵ4$�yF,e���Mv9k3�ꮕj��:|Cj��w���
C�{#���@.}y$��MX�`��%*ddN��}vx+�w%qid�:��u��t� �Jō������d$v1ʐ���v��̡��%77�QҢ���2J=B���XU4羐�{-v�}�g�{��42����X&,��&��� ��wx=�y�|N���=�����<��}/�o�E�[d4�S�eo��OCz��Ν��Z����B�ͫU eg���z1v)��Z�wޏth�t:�иq�#	W���)t՛���
�`�^[�H'�n�=Cٵ:)�
I����C��)~��]�j	y>�Bd��B��vlN�͈ؠa�Q�zE9Uێ�U㑃e��D�"��4�sRn�盽ޞ���Y�� K�.-���HnT_�Sӡ<$8C>�u{r_z��G�ϝBG�z*)��7��-���晓��f��ſ�dQO�!���iVG�C!䪛��5��-�u��5�
�ʊ��w��l�6T4	'D�z{&���
(@�n���Y��0k�Q}4�I��L�"\ }ʖ���T�p��Җx���,�8�]��bkc$k��_rqzs�mV�^qX_CP-�4�&P�#�t�Rm�fv��$u2X�FFlך[B�Y�A^*޸�{��]_*�S��$���l!n2r��G��u�2���_�޴��O��=�{g<�y�'��i�h*�(��?o\Ͽ�<'�z��ͻȶ�I5ߦ,��Gg���B�9�`�崲���Ľ�D���\0�e�yMtƪh
�mii��	�.�34Y9��>�:�j��m[ƭrxf۬6�]m7׫[�co$Ժ��Hr����n�r3�'�ٚB�l��]Ijn��a��.I�/]��Ʌ=�� ����['i��)t�_1MtJv�__K
�#V�a���-��HЌ�r�mv�3z���zÆ���Q�Y�h.A�"��[mr�}"*��z�Br�d��|��,�o����m-ɠa���E\�vz�a���;�9f���$t~���V�ImEKr��D��{[�SA(ck���Tzq�in�Ƒ)n<N�v*>(dSe�U�oc���f��̡�ퟒ�����ղ��Ke���GH ��X���ZP�g��I�h淹|uTL�C�v)�si�v";�y;�wz��ߵY�iE�[�����r���@�-p�|����kz���P�{�ޣ;ROs.{�<��8�DǄ�e�tR=e�����7��#��O �2�;:]��#�f��Jc��G���=��w���M��H��b��^ZQN�;R�����'����||����)������j�8j����H7:�k�Lj��e��۝wVi�U*$�� ްu��frN�,�J�h���k�C|�70�l]�sۦ1;Հ>�Zy��%�8�4,M�;LW@�6�t��Ƥ����4�640͹��H0Q��R�ϴ�)\�F�$R+�)��k�6��a�V��m�@aӱ]�������T��~�$��J�`վx���C��(ʱ)��Kp'kxt�������,���N*�b(R�Р��ʾ"ᔺ��x��=�� �&ژv��b�V��MHr���)�̵Յd-��G*����������Nǳ$=yLj���&��a&!�D��2�e���P�t��Oi�>Q&���]�h��Qz�� �,e&&k�m�$��!v�:]=��r7�L�Wj�Y�^��(�g��c���R��� �����õ���!Ɣ����2f�ɑ-�lL���`�#���Ƅ����{o�M���sK�\a�":��N&��W�ǆs�?s��_��_���ˑc�h��.#��nP�j�%�#�Yl*�fb�%Z���f`��3����rbj8YdD2�l)��&aTF1K�[r���6��l�j���1��)�7[w�@̨�P\ˆ-31p��7029Lʆ��S77ra[��MK�"�+�L-��)Wr��\u�Zʢb��1��\LA�����[�����L��e�
�����.��m&:�n��2��.Z�H��m1����D��%c�2b
��ֳr���mc���cALm�a�AV�S�r�M��st��ۻC�4�&���aiq���im*��ta�In�\��շX�֦$���++�*��`��n\@��IY����]MuSr�̡P�G5r
:�Uw,1�J�Z2�bf�\k[+bcq�-����o���*���ۿѳ;N�����9�x[(�,;��M����WS>����*W(7gw�m�W��]v�����~7�g���8H����*��tk���F��릢��ݩ�2�����P/���ri�L��{{�xm�;7�w�_S�^թ���ѿS��g�� ���~j���8���O�N
�< D#�o��6T�H�?Dez�u�S|iA�.tr[�R�`�A2�d�NF��ݜ��b��V҇�}!����;�Q�RaC�����LQ�g3C!R�w��Xʃ#�����:}a�9nn
D]�F�Ϭ%v�Br$m81���$��c�Q�nbW��5RC
��yh�+�?��zڭd�B�rd��k��*�C�^��@��4�Z~��x���W�~R�e�=�qP�ܣ� 6M_i2��P �����NC��0h^5ڕ`UC�?<+����Cxy#n�q�Q�����8t�<�LmI�$O�%Kr�s����XP�t�|9T�����{ND����Ԛ���CF�.�)`/��D�b;���+�	d����8Rc��ݼF�5!p��u�( dN�%�r�fT�E����5�om��dma[�*�_}�ٯ¬��7���.��z/�΁56:T]�]��i�S�h�����v���}V�
uB��ҕ��im���~�ZJ��>�7��E^{�~��H�{�rB3}�DP����#��܅�\���0��y�^A�����;F;2 ��QR�)X2p3��&2\��=��mg�Ϫ�o��Pt(��Z4������h��y���xgXr�����{�C�ѣA|�^��P��yBX�+U*Y��:�G�(��I͡N�rzub�n\bU�y���q�����@[���by
�G�@�d�͖s��'O!���߮9I��R�ci)ȥ<�^ԡ$VH�&�V��v�5�׆Ԃ��*\CK��n|�d:�^ڂ��x���]��zS�2��'a��1FT+�W�T�������_����5�Yw}��E���72�ޘ}��U��"gz�{�fQ��`��b�+J�8�p��-]�­��'���%&7(��QV�}m�zB��ܥlCR��
xl<6�o1D�ЁJ:�rR�Ѩ��Q
��8yHU~?������wٞ��ǨG�.,1;���5��|��IhGZ�����r�ݥXb/8�
g
����_�P�.VWT���m�Wr��y��3����wW�t�h�<
���� [�&C��*��[���m��f����(/���[��|T��;r^�^�ARzQ�Ԏ���a�j�L^Ό��ٕ.���xu!�*괉V-! �ӥ���,��ޓ����AZ:�����lӲ���^T��`ܣ����稳��#R�MAc���:jov2n��H�9�EXS*����c����[��C.
˺�$�0kc�_��st4FE)�S&S5�G�
G���A?y�S��z�YQdF7C���;�)X;y^t�dl)�#ـ�
*Է.ع}%@6��)1ݱ�'�#Pjl3^�=�gc�-fw��]ҭ�ؕ��(�Z
��?�*c	��y{�;|#aW�cQ�n԰��7���.2	�ה��;l5 b�;7�Ð�T��=;Q��G'|D��Me�v*��n��ªٌ�0V=|�k�����J�Q�c���^���S*���~vd.�*}A�-�;2���d�T��߻��\��lJ
͊�	��$9�P��ZV/�5�y>������~5v�I�n��ڭ��J���/��R9C]RU�^\>p���ϝu�O�dLL!���ݥ���jX��¬L%*��	��i�MOaPRf����������B��69J����hA���	jTR��"��;4Ә���D�̈́�(��jOH赔:Wn; *��͗ R�^"��,���;+�.�m�h����^��@�����{�E��!�BIH�������DU���"r��zƇAE��KxlUu1��)�넕��i���Pʰ�G����{~j�?���r�'��4��uF���7�WsN\���СCs��ɣn�T����3�`��[G/e��IY�HWj�2QZ.U�ES�����`��22�;r���xd]H+�_ѻX��aOst��U��B��=���V�w7����hZ�dў�w��>LerŖc�&���x��qL݋l�빊���#�i�?|:겈���ͦ����\ɏNZ����r��Cjkaa��I��=��Tz{�1u�Vk"������ף�]J5V��Z$[�{E��q�������X��'�U՚��x���ϕ�(��\̱^Po��Vi���(��.E	T��;^M�@�\�6�6`�c!���Bj��;�Ԛг�=�g�jKS�D��v		N���q���k�� 0�).t�(q�,uz���=Rܮ�^�Ź
�u�sѽZw��z\�S�A�4��� 섢A����4@�F>�F�u%k\Jc�0�ݓ糡PaÂF�;8�R2@�} Ѥ"�H������ �]O��1qJA�.v����݊B_��*B�/������4��j�^��uIM��U^�f��;��Z˰��%T���W}N����Q�D��XO�m��V"�WG�'b��Z�r���i�W�Ϻ�� Df��V��e�=IN�8{��s��{���0���P�N�ķ_Qm>��T�����Ũu��W��7�P�Vȑ�u�L���y$0�<Z)�+�?��z��u�Z�¬\�HwT��a���ڻ"3�W�PT�Ic:|j@rv�TX�v�1��'�m�ɝ>~���g��X(z�:c�q
�1�����l߼>���Mm�X9;��~�R�B�� *�}k$85��u�{�ЙRH�bm��,��ر
)�Șn{��Q�}�	���{��iv��l������[ߗ�]�������}�c^>B��+d���v�.�&1���b��:Py�`:u������j��c�(*�^�� �ʣ��sjX�a@�"��AUD�U�P�<�kZ�TU6g���Y��X�MD�r\z4��5����
t�9Eq"����RaZ"(^w�v[߻Ӏw���իC�F��h�{J�' �J�x�GP>�X�w�����q �O$s7o=��|�kg���9M��֜b�d�(�Sp�w�[7�i��Uq��ڰ�H6� ��|��8Ň8�����،��t�źSDU��mk��W�wtNz�}��+��MUF�/�����Jx���#:LO!^��t���1�"��"�����.Y�6mȽ4:���~n�b���K7�:��7Ɇ*�%	������;��㸷�b	=��7�S6��yMl}�}V��}�T���q �ò��U�!��~~z�>�KHZ��w�:�����tV��~G���b����UzC� =�*7(FFD4�i�l�n�K6Ώ5���U�W����B��ư�=uB�T�$4ř��)�0t��������⁺^uθ���+G!�h����noVl��!�F|��9�˳:�r�?_]����<ս�G͵8������w�s��rr��a���"FB���(&
�|���:d��l\�Vīq�%kK�69�(�,z���Ѯ�������lӲ���i�J�yr��<kw��`�X�*�I�hhˬ�ޙ��S�
_&���Bñ���5Nb٥N����dJ'k���2N��F�t+�	�8�aŵ֝��rI˥R���3���[s�B���|9��)�:��>���7�Xɺ�5�T��5[2�l�c�:�b�c�a����j1���	��#"�t�����#��#�
��[��rOQ�2ǼZB�e���Sθ��*��Co���%_�WVT�+J�p����>�� he���+�TϨc�[���|�Ѥ�a��9˕��Q9�ݺ�����ݔ��"��>~�A��Cۚ�>��L�hZ�`�<�rs{���鲻6�����P@�j�MS���>�O
�����훠�`����u&٫����%`���C	���G��_:�����Y���Oh0`���<�<�Y�"Ĉ�>�OJ�*�v&�ꃒ��m��r��H1�^etq���r/("�OL9������e��>\���D=�+Mh}j�y&�6r~�v\@)Q;��~��E�L�r#�3��+�حt���͊q�QڭŜSe�vnK��M_N5Ξ<��*����fo(��ʞV����Lu<���������lkJk�q͐_,�FFH;�Q�lrY� �����a
����e�/��>�=��g/��=��fe=r�ªb%�N"b��&�cs��#  �]KHq_H���?�W�puXB>�TI�V�n��=T�B��P�5��գ�k���c3�����:���RX�H,�^��ӈ�*�@9F���}sF��AE@�n���C1^ƽ��z�^��7��]����zlU*�w*R.��4��C�U)g�)@ר�����.�(w�޿Xʭs�!=t�� ě����e ��w2�ax�=cP�ReN�ߣ���b�DW�hr�ob���R�����G�B2�d��	v=��~��R���R�Z��t��К0�l�n�׋��uw���뢍���SA�����j~6����yԀ��Hp,���h�����fI�2�O&�DP:�1�h�VW@�TcO�՚�g�A���#���z���*%�tB
i���ه�l�I��h��=����[���Xq9H#�.M�����5�╗���W^9r�� T��N�����qd+�M������-�l
��:��tK�Π��� ᮺ����F�P�*P�Ģ�燹!�E�o����糾f�p���Mӎ��@:+)� l���|���R����,ی�ru��Y����ҡ��bUu:/jÈ�{{I�)Lc
��u�>��H���S�r��8��F�ϔ���[��}M���M4ir�U����H���`��NV/
u�<k���[kԺ�b�.N�����-�#<�z�H��� ;mEE�pٰ�'��VW��#_Ks�l��%
�B��c�T�@(��NKW`�(�?P�C�{�`+的]�y�.Ɗ�����0'�m��(3[��M�8��b���:t ^4����]P�p�+���@�:���=��m��}�^ f'�/^]������}�x:�\z|��$��� ]K�.%Q��`��E�yfWW��zR��]N�]���_[�a�&4q�vi�_߯��X�|��5W�))��q�XYW"��3:�F[M�v�����F�� �w��U�=��묖�Q��7:�������wi!��/A�rQ
=��i�Q�9[����姴CB$_j6F�RXA��]Y��gk�0�i9������F��m p�y6u"T575�h�ouj�]��__�©�n���.�UҚR��(J�B���Kжlխ��X,�۫�0E8�Eaȶeq[[�M%��#���+�;ɪ�Ar����B�)�I݋C�t�Տ|�[N��F���hF���p��3����1`)��ڳ��I�	<�i���W��r˧��u���^S:�t��]pa,�)F�!Ђ
���$�X����b8��Ӯyc��}<*R8��oW,'�S�xtGZQw#}9�׺6W�E��u����_Oi�D�����(<��W^d]ȷ[!�H�x_�W&�H�s2�y|�]�GCI��f*�:���E�QK)	v���#�z%�8�4XD��|w��ZJW�����: �db�k�]%Uy�mv�W=Y�r�3�%m��WP�Q��l���Ά�+�6��0�tyg��@0���� s5ϭj��ē���:Q5;kq`�}�]����F'Zy�l��Z�R���N��vظ�u����Zv��4e(��x�]�ʰ�&y�C���%���\���<o�FP�h[�h��Dv�"#;�1���:w�f\	�� 삌:k9����U���4�J���[�].��j�B�6�p�kֹ�����G�W �F�� ������4��(���7�ؼĬ��ʖki���pG�ٖP�\V�f|�uPz���
�A7���ٿtH)}�
����f[���Vo偁�'��}�ϖ��]­ܣ�j�iXڗ��<
��"���)
۹q�Jnu7�E�ɗ��N2"&N�o�^ͶI*oH��v�e�Qef�L�Nₚ\Ȁ+��V� �����Y�17B^�A�n9�)�v;�i	rf.L��渭��w��;��]�Pw,h\�#����xuWPrߜ�O��Oǟ%���f�S01EJ�2�mZ�!��2�7)fXT3�������T5����+�����J��1��QGsܙh�s0pLv�CP֌P͸�1Qf��R��r�r���̮��wt��m�9��nK�j�jW)f3)R�hkZֲ�]��fZ6�&1B��ˈ�U32n�`�2�S3t���
�wL+�m�i�SP.n)�LaU1�2��sq���kP����m��6�b)���[���[��ͨ��+�eu�2�(8�Aˎ0�M��wnb�d�n����e�ܵY����2�6�F�T���M��n]�K��mMTm��em��q�ۉn8mK53T�h��,̳�u5��+��n�n`7-�����-?�G�^Aۗ���&��9v��u�o1]��R���|�rUd���l������|U1��<���L���c�7
���:�g�5��c�l1��W�N�}�� �h���YR�;;�k*&���Y�z��0l�[�k���s��@���ɇI?!P�w�G��b,ׯ{�� �Xo.�:d�������{P���\WeW&�m8������q���U �L��}۸������ﰩ;gn }>�yHV3���H)��u��? (��s�N�v�C��;�X)�%b��醤8���~�b,5�O��k�<B�S����<������~�{~k
��Rc���:�٨
/�>�<@�:C�Oܠg��a�ζ�'�T�sg�8�MJ��aN2c��^!R���SXw��0:�7�;�z��sxy� q+;T��J�AN��	�8�d�/,��qyu ���S�x���h'��f���9���ra^�51�sܓY�J�v�����۟{���9�O>��R
t��$Ⲥ��P���LH,�:���(�?uq8�0ĜB��.�z�O�bAC�~f>�1~�� `zc!@�|�b���.��{�FP���l�&���0��f!��z���pU ���I�>q�0��+Y���:H)�1���
,��LMa�1S���� �d�����oww��|�����gI�H/�>�|�L��LC���Xk
��f��
��nZ(�T��?0+=N����J�q��3<�+;H���$x��X���_c����+�#���'I�.Ҥ�'�?r�>�R(u߸����~����%f+8���S�LI�*�&[>d�Lf$�Gٓ�J���%�?�Tr�g��{i�E�~��@0 ����C�O����5�W���6��񒾦0�h����'�ʁ��pߩ
�
�=�1 ���5E&wC����}����6D;�:>,�ߘ�6R��8��.�(�1����>cz�7OF=�L��z�"$�:]q���]�z7���D�8�p�<�lv(͌f�rCV�M.t��[̑W�B���U�W����w�O�ϒ��'����
�P��L|O�1�TP��������T+>d�>ÈÌ+5<���zïs@UR��i�I;f���,��!1�Q�S����_'�A|"��� 8�����e��X|�C�)��v��X�S���ԟ!Y��1=-"�aS��$�VO~��Xq��1�����w���ۜ�ߺ�������8���Xj~@�:N#���B��(t��<B���1��v�O�SH)���}�0_P�oS�'I����?yI����:�]>s�^���߸y��)*LB�ǿ`ힲc��r �g�c=d�
o3
������l�N�>s�ά5�l+�'}�R?2W���uE ���`��eI�<��w��y�~�~�Ϲ�+��R��>��AH.Z|ϐ�9�LOY�I���jA���E�0�>;����La����%u�f���g̞�׽�<aY�<�/~}�߻��>~���:g��5U@��1��8�����
��~g��AI���Y�=L@_yq ���bq�H=���,��}��Ϫ�1�s���_����:~ B,<aS��~h$�
��v�(����jA}`]�O5E�u�&��
�O�އ���~{�L?0�):B��y�Ԙ�=���AO�y�����?y�w��N������k����>���ꁈ��=�	�
,�՘�E%I�~� �g̘�}gjAa���x�P<��OY;q? ^�V<����ȧ>�"�j l�Z���;�0�q���$v���5��e�间qYP��>R�:�H,=��Y�����*q�a�<��H=Xz��gH��*C�wT<x����_��އI+�zɌ���j(v����}a�OP��?Q�a
Ì+��y���e�T�!S�
��p3���zC�z��P���<Ldd%���9����M�u�ʠ;��(�'�}���r%�|�$T����2X��e^�i�le�~�w�uo'/w����zƧlp��d���eE�J�����]�jwV�n��C\�1+�#DFDZ�2��W�UH�������� �L:O���S�1 �O����?'�1��!�?!Y������AaXs)|�bN!Y��3�(���Ԃ�ɿSY�%H.�s jq��A/�n���4��~p���$�tü������Y�N8���1 ���߹����}f}@�1��Aq �T�ÕT��Xa�'���1Q��
}�{��]�1K��9�'�F/�g4�i�LE�t�l  �d�.ނ�(�\�(�"�_J<I*��Nr���~��x��~����ïg�����fa8ϘbtmPԃՃ�"�XT���;I_��L�x�����"��+>f�B�֢R&qæʗ�"�Z	&�SX��*��{{���y矿{��>'��
�>�"�A偿]aY�Ă����1��Ă��o�5��1!��rJŚ����$�
ξ��Xt�X\z�D@�� T8R�3����g��l5 ��젳�J��V�*z�^���:�P�6�XVe'9C1'��!R
tvY>u���C��&Z�0��\�8�����v�����{5 �j}���RT�ͼ�*|�J��Z�$����L8¤m�����2T�����$�
��;;�:���5�z�̓�t�Y�������oIϼ��y����c��&2|}f%@�O�<q �B�]��CR<��|�P�OY�?3si=B�����Y�
�`��J��0��t�P���~>���~��>� ^P)u֫��Q)��-�ִC�yq��+Wa偉P*wN3פ��Nr�a�=L`p��ԂΘbbtr��5��,�;O��Nv�?}�����/wu}�><�s�%b���R
O�î��:H,:?nCSߨ����jA�
���Ă���d�~d�7�1��2o?gI?!̤���P#�cª@�ј��6��1�U��ٜ����k��#�'�{0#d��o�M;�i.�����&��0]�VKƋ�P,q���M��	S���}#㔣���Xu[�U�Ӱ��V�ӥ8�RK^o?� �\뮿s�z^������q'�QH30����*~�w@�1�W��1 �i���RT?ZAN"����v��,���P�l*��:d����gm�]ν��3�7�;E;d�S��jO��}����
��:��Y:LH)^�1��좆$���=|��5 �HQ�
�S���z�0��1����������U�o��9υ@�&�}����ȳ���s$�<I]N3����P�t��P1'hW��'[��c�f�}���g*�j�S�
�!�>u �A���y�����9ߟ�E���O��1 �X|���(���������1��܆�d�Y��}�:H)*�{�b�<2�O�P1'���ԃ�,���T��[����?��������v�����OX|wf����W��a�>�v~���Y�}�^�|�N}��'n0_P�{��P11���H,;2�1��J��]���w��}��$���Ol>CR�~�ɬ>aRy��$q&���(�̝���z�N'2���HVN��^2~L`}��|�^�7(�ր��#�2�=�e��{���DG����>�X|�T����Y����b)8��̇I8�@��3�Xb,�
�:�1�W����I��'���$�/���N�p�^t�y��]S���s�}����>����3���>�Rc8�YUH)���JϜH<�[@����m�$k�b�C�La�1��1��dϬ��:O_�� xD}����ˏ��[��!�	�Q�1E���0�<� 򞡉(��=��=aX{q�
�Y*m�Q|`T�bLIP�,�}f{HV0���O�8�;q'�Qa�}��&��q���'��=��"�x{�t��{a����SY�>���AJ�LI� ���Ma�<�Ă�3r����2g:�������t�ɯ����^��oN�%Y�V�ib���7k��$kiҮ�F���&�b��6���5�h�^�N��a[��9�r �-�7Q��<�$s#Hbvdx�J9D!l�����6R� ��������z?��׮�
���ǌ�&2v���_Y>�y9�AO(����y`��z�T=��Y���t�1����,5'�4�ua�H�8��|s��{�N.K��8 lL}{��& (��)1��I��ݚϙ?g��.��+5�짨����嘪�S�_2jOY�Ǽۤ+٩��%H,����ٻ�p��;��~{��E8����T�f!�~C����X���q����p+7�& /��>���l?!��)�Rk
²g,��f$�y� (�`Te�uRկ�����{ ������i
ä����
�ٙ������Qg�b~d���=B��~��}��$d�Y꤬�E ��"��{ 	��B�q�.��'��0���wg�La�+�lH,ǾRj�VwE������+'��HT�l�2~La�6��%}d�������0��*A�λ�k*'�~�y�����ϼ����_> ��jz����_�_���~B��H��1k��t�P�7�Z�2b�o�)1׈�FӴ5��~�rN��Xx�ǲ=��X���z`>8������Wa\�����:g�XjN3�<K�!Xq�&r4��YO9��������=���l�:O��`�l���QN�jAC��Y��1&%E�0L��y]s�8�}G'��;�� L�}�`����ǌ
�!�1E�����I��~�<�+���i<B�y�c=I�5*>�ﴆ�1�(�B�)=�����~;~�۾{�w���l9݆01����J��LE �iդĝ�Y?}f}g̘Èx�AH)���M@QOY�:� T��m��2|紅���+��S�ۿe�޳��������I�?2W���h��&�'jʐ~����Y�Y1 ��l���X���8�q
�;�3�Xb)���P�ٯ��& .w���{�}�s�߽?(v��2�z�:�&XJ֠�vMacz�Vc\'����}�����xNf�+�+��Ѐ��4�L�wr*��E�(\C�f�!�g
�V_גL`����   k"���ʀ.�8 ���!�<d��!ݰ�aY�o�;H,��Ow UR
x�E'�����B���~�$��T�'H
,�l����b��y>��r��g^�ߧǟ$�T���x����P韶Ɉ~������L���lԞ�X��@�8§�P1��Y�u����ɹE8�Rj|� �y��������/^���N!R|uC�OI�_�XbAN�=q��~B�P�������a�?w��t���:����IRq
����҈�W�'+�Ҿ�G���b����(%�gG���\�^����Ch|���V��<�5�����U��%�Q��6>��G����q_R���н5��,:��U�KP�4g���[�t��|]a�|l|G�� ֟P��X[ں��uAgS4�\��1^�T��Hq����0i{>Gƥ�<�x;)=պ���藽�L��r�LP�Z��	.�8Z��uw��4�Og�C�6o���g���!�7X��n}DӀ�� >��t��J�*%ߎ<l�!�M��S`�0õc�u>ɨns�cޙ�؂�TyZ���q
��җb�%j�w���Z7 W��g.F��V
�c��[k)����?^BD���I�R����b��E���S5�/ ���m�iw���赴�
�g-#oo��E�ûQ����f��iU��x�{e����]���WFB��AA���k/+�Τ�in��}S�;&*�g�ܸ�HH�pK3�5
�Mz�H��eRȧf�̨A��@�W�kJl��ǣYv�pH�
��Ѳ���j�9N}�L������}0D��x�T�:��"U����|�P@kML���W��gU�bM֭���͎y��#*v[�R��8�{ʟ��V_п��i����IW/%.�eg���P�åC����*���{�S�1a�y4�(DI���틘n�h֪f��P�X�p(\�P2��
9˹��lA�1R�"(��o�Nb+^�b�&B3thXRhS����1VV߳	���W�Π[�y��I^���=om��`w�t�׻��f1���
S���+�wh���<��NP��:,ׅh�׮��<T���q���(�5U�
A��u����]�U� y�S��[�i��W�7>�x <��U�3��<�6:����"��"����{+h�q�ŷ�d���Ю�Z/���.$1�i�GI�]�9P��%��� {�v�Nc�6l����C�T ��*��\�@kMu���fy8���ݸ�)����MR���D�(wRS��ɣj�!F�Co�������<�;Yi�qx:��E�
��̬t��=�X���H�#���+��XCQ���|�׻*���A��QXP�Zp���]�8�G/w63����Os�;L-���_�O}�[�.shr5�8T^̾s��(t���Q[���X�!�x�+�5��
��R�J����*���A�u����*�)}��Mpm#�)j~$AY_3�	���C�4��v��.9�.�dS��'�6��j�	8�B�W�D㞩����.0�o6;��A�`�ՙ�S������ 셊h�����}J�M'oZ�4Q�E�1� ���ٰ�(9.try�q�!���śu}��3+������J�y��y8�Tq�v��'Oi��
�� ҕ���[�!w��5aa%/����V�[A��kE��@e���R�F��{��������2��8��!���������u����������=��6�=��u��P���x�iv���/s���x:C�F5[tx��A$"�L hSt�}c�۩	ȑ�*QALB�>�%�x�o�墐�5Ê;̝���ޑu#T�'`��#��@�^�+��GT��^���.ڣ��C�:�6��^�/{+��������|c���#n��U'��6d\�P�ϯf��a�=�㰁��X��CD�3�����h1p1�
���t�ʜ�mP�qJE��7=1�D�.�^�'�$��V��=� R��'0��<�|��J�ʼC�ZF�|J�fPm�a^ޯ���A�r��?���ఌ<ŖH����9A���8�LMm��Db"�c��%{ΝCK�.��!��Z<�[X��]^��� ~�����#-5��kw�ͮ�.�*Ҥ9��T�Xu��U�5ify�\6�[��K����A�$�͡�����&�Ȇ��3�9]Y¹���Z��K�xxv]�☓.e(Q���yW�U���
ub*f��0�����k�[�<�+�_r�4`/�	iB�㤆�b�9��4�D��SP�]�S*��wq|j�}������:�Bo<�M1������t{`vU�*���ѓJE��A'}N��Y��h$+n�?�F)Ъ�e�P4kêB�raX�~���BP����ͭD�1�zm�������;G�i�*��|#��t$�ƾ{Ws����b60Tka�rz\Ts�}�]���W,A���9�u{���W��ch0�G��E��/"�Y�ty�?�r�����4/�N��8]��(�1�&�Nz=�J�����t����f�%gk$1��_���ϥe
C�haACzG�d��ǿ+W�u��_vU���;�+ ��:orv9��5F<��3���q�NN�.��=oM"�ɻyB޾�A��& ��>=�b�xh�iU����1O�۷m�03��Rr��&�P�rg,w:�GW]bY��V��u�O;���Q9���_֚�W�.D����R�2�t�GMSV�ԅj�e�4�<���w�m뼔,_{nYeX�e�9��Y��ܮ��Z��c\�x�uX{�:�t_����Y@�坕�)QOZ�h��H`6)�z�9ϴ�0��R<]ѓ�Lt7����4�>�\9#rrc�|4Ѩ� �աX�c]3�ɒ��`�k�J�W���'V�j�]ʯF�+,h����P��gVګ�Xr��)p�ޗ���o\�̫ �Hu�;N��ruu�T��!��d�6el����v����Pð.du�Oa.�l�8��`n�F��)�y�x�5������l��WW�>����s��K�+�`x�٩��F����j�`�P𗧺2]�G$���W+0�Q�|	%�4<ۚ[]oV���/��zֵƘ��(�>�1�MM����ǈ#�=[PC����^j*�5���>�H��y�:�,-��֙�yۆ��F��b}Pk�#H5�8��;6����3N �s��Z��*�+-`ɓ�G	"������.ަ'��vǫcqi�B��*Υ'V����Ajv^Ņ귕2N��3T��dS5*h�RA5�MA�?^un������z	!��z;�Ib�I��6���c6ݚ��V�xc���ӕ�f����J6ާ�c!�;M^I�Yr5�R�l��"�4]���ȯ#J�amC	�P3|	ǰ�;���9���X�L���j��kf���L�jvS�G%��tVX��(�'���6��uoZ�tI:���N���W���U�{���Q�Y�g$MnA��\Br�sW.��ziV2��Ӟ��t��P�ic��Q\ ���#������pDoN��&��-i�1�s�r&��1�enva����g!�S�KB� ՝W���ۓ:ܨ�F���2��5�"vV�n���z��x����9{�8�v�(S�j�p�	4%���.Ώ�j��:���aj�u()��V:�]�f3+�����ij��r�Zݰ�ia�!m��1��Ma��Y��+m����sk.��桪R�Ke"�I�`�3H
TP�Z���Ǝ��s]2c7G7u7R�]�����*��wGP�F���t�D˘6n�)Fe�ڷSn\�pk.�n�V��wSm�U��qL�ݺfۨcs3%��ܺ���QˎZ��u��wL�V�Ze�]���j�;L]��m�]st�\�\����3sm�f�2�8���S[�EUqnd�rܭ�r�ʈ��#����[��e�
.an��%����WE�r�ws"��n56َ���U��\̦[�F���s�n�#h�*n�kK[stݡ��v���˥ʤLs�ۮf\[iF.!r냛e�L�X�7f�ܳ]��-�2�.3[\�.9�ۃ���5��f�T�faGQ����i����3�˶ۻ] >��Or�n	fvRoG��I/6\��dWY�
�{Xo5��26�6T�:�].�\C���i�T�U��"�,�:|.�h�_<<9~_��8�>���n$��]���
���.��]ep�%��#�٦�1�F����vw�����ǫO�C���4��"�|�p�s0.+��5Y��;��lvo���m������(ظ�ѱb2(ȶh\�;��r๊�=ɭa} �`�|��,���d�j�W����+Ͻ��N������z�ooP6�����ᒧ^�=�ן��5�z�|�{�J=�6�\�Ǚ�.�^OCn���PF�TCO�xX�2�ü~�2��3��:�6Qe�2�v::eBS�U������k���x�� "k��/b�{�(����r^O��[���Xnr�����(��.�Y�����o��c���E�Ѡ�k������ݫ��y�{4�(DG�w�`�{����	���^\F�}���t�mX��
!s�+�v��A�L��^�^2d�+�b�n�o�ӵ'cV][��k"�y�92��.'&�`������0z��"��ZUZ~��I�I|����k`\�-���j�n�8��A���	�z��NI���*f����Cٺ�@���.�����n�r�u"�cK�	D�{fC��yK� ꎑ@��W��^^�|�Mħ�6j��\�+�ć�(����&C�b �t�ª��^�����ҬÝ��b0V�fO}%��UA�:gu�J��5�V]�h����|�&#��*yb�y���r��9ԫt���u|em*�O9åޥW���(8���^���N/����*�H"��u�}Ƒ'��v����Ē����)�L��b}v��2����_U��ʇq^h�b�ψb������c.�4�&m�C�t
��>��r��ꐁy ����ۑYY8�H9��n|�v�Ȯ�C+i1�B5tq{Ʈ��J��h�B�u�����7T���Z%f�Ϳ��� �SϮ�@ǅ�*�5ҤE#i�`n�}7@�/�Qu�}N�PU3Q����N!��|�5[��]�L��#�oY[ٱr����I1|��x�Y��"�T{W�߸ⱑ�-
]v����=��5���#��|�O��3�Ը�lWG��
ĎSNE`NͩQ�T	��DP��8�)�;�
�Ty����]Z ��V)S���G�B�R�4��pH�U3�ݴ܅�mR�*�APr%2����Wё�ܯ��V�����sM�}�Jw�Cì�<�z'�xS̞g��Ӟ��<�{҅�)
!ߺ���b�S�e�Cv��3y4`����*:K��iV����k&�<Y�Tɛ=Cw�8�w�\?>����Q@�>��,0=��3ri�� g`db��F��n�ULCs�^�+�c�}��h�ܘ�-���X���8O\�D'&��#��HE�hdɏD�'Nfn�X�ycpniMu�U�����^9������� ������g����z�SI�����GSH�aL�����י�<��j;���jDa���kZjT�,^����ʬ\Ê�X�=@�'J�s^qep�]h�W��i�(<����(�C��������owܹ�S�DO�f���2��o��G�9M��﷮�<�1OK9����0���������f7�E�K �~;g�T����:�Õ�����e��!�������7��*0l�̳��ͥ����z�ݣ���s�b�]@�U\�uS�=55�Z�?+���x���ot����+l[���f���9-}�D���s�x�/���.���^�%6��4I�	;�Q�;�c�|��;Vm�cf�o#u1DS��3�;��O�Ua���JH�*�O�UF��o��25��T��T���Z�.��S���˧����'l�����=�0�vk��dґ��f��+Z��:E�MȲ��)��XO]��J�?Vٮ�w��m�]*�[��Z��5��B��jF'WS��a��G��^�ﯖ�i�w���y�޽�)7k�$�U�r���4��
$��V�du��F�YM�����#Z�	�>d�cGj?)�g�b�]�F�<�}y�uܣte#�h�urE� Z�wIĢB�'Ck\��ꯪ�@ē��i�"��S:v��-}DS���Z�/`T�~�'�,L���fn��b�%���z�T[�r�у�Q��S�u�a��8�
��ຢ,ʊ��C��ShL��p�`�M�z=�J��w,Ɋ�Ata���d�Ԟ�Y����m*:V��7[�E5^S{.-NG��na�o
V�uݭ˓��˨c$W���_0m
�~�瀇�*�^��`N��	�K�|����案�B�Oq���x~<���<��B:$l?6�ղhٸC���M%8���8D�N<�����n��h����n���p��EX,(k��$mݜ
�f���6�!�q�<� �*d�����_s��*��Y�2��M��g��HU��b�#�D�}�8C�Y_1(]3[��W���n碌�)�J�2��2�x���j�f>D��]dCDfÙ1�E8�O��r婽{%��i��:b�}Gb��_Y�:��R�g~o���ӼYG3�0�����c�u!���-�������qN���Wi����Pt�UD4����J��9!�6E�{�����#0������U8jt*��<Ո�;�C��	z"��������	u�2���W��+j�s�uY�W��l�b3���s;*-�P�l*q��1����f���36;��X��zۧ�Ob�Fk��Gj�xRV�����
�4�U��!l���E�GY����@�k����kf��1ﷷ=����)����f<÷}���z;�qj|�wl��zm�ip�M�[�W�F�P�ǯ
y����}e9}{�U=����T+��Z�2��tQU逌�U����+® [���������P5&���%�#bj<�O� �=BX�b=Pa�#C&�Y��J���{���.�$���+"��9b�i���P���M������ek�;�e�tg��4�d�Z�#\�2�������g/@#���N]�1to?c�B"q��L���@��Q��V]9����S��P%�+�ǅ��N�}�;c6 ��dP�KzJ���� 3��K�:��~�{X���%��O�֛KH�Ȩ���R^��+�w�����Pv��W[},��=�_U�YP���N�'�|�;Eĕ]�+ɛ�#���0|�P��%]���!���������v0|��ꨊ��g�I����;`wX}����S3q����ٮ�9;7���~�qŃcJ��+���Qr(p�Qu�nj��ԕZ�O�Y�>0zGl�f��F����jT`�J��:|�;r�m��zx�<ƌ;.����R�B��-�plm� �)��AXic���:�s{��=}��Dd�aP�"t@�!�:-�E���������
9ҡbz���H%n�A@��7J���J����S�J�\kE�<;��Au��w��`ǥ�JA�SP���AJ��f�Oiϑ�������l��{ �"�HS��5�mj�P}����l��i��+W����{�U.�N�B�V�{l��l��;�Sg�br��f�cF�K.젥�H&%��G]��ݳ��������-1[pB��_x{�������FJ�1Q�}v�s䪝J�(��@ъ3`Vƈ�B�[l�PF�S���lj�01�݂���נR�G	�{
by�7s
󵧨a���0/|'�v"� ���i�h`����>Z'��w+W�ꕔ+��iV�=���>8<�M@/ ���iIMx��y�ͱv�u1�.�dI�����x.5`�x�iC��[�~�<p��\x:�
��7)`D�]>���
��/f7f�x��]����Ca���^�F���lFʉ���������K�'(;?/{)�=�=�����<K�g<��f��o��Z�[�{��6Y�SP7|�C�5V�pQ�L������lϔy��ۇzIú��B!�4��H�}�b�_�kb���^/�W��C��`y�6����x�O:xЭ)�;	mA�}9s�	���,q�t��΅����c��q,����l��Jp�k��Y;��2U��"��B���o��Ò�t���v�貣����s��J؜�3p>ҙ��'�B,T���
r\����Qn��q��L�e8B�T)��L	�ሾ��?n�V���\���d4�u�ű".�=�,FL셒EH���>��°�Sc�HT�^����t+�y�Ę�0�ߦ%�Rd3!bw�7�T�련�Pд�M2p�s:�@�)����bC��C���}�����7�>������W,�FUL&�>�����50箫� �Lw�뗞4`���C�w�*��^Gu��efĈaȉB�8F(q�
\}���.x�������Քmb-C48��=&�,ˉ�"�Mt�"�:B�57��_|�`�w��'0}�E�������N� �J��7���|^��%}�x
����7���J��0��/\�<x�.�?���v����?YLϹP�X�P=�������ъ��aXqǣv�UiJ|,X}�3��Ji�Lqt�|F[H�s�I�BK�ʜ�_��u�N����`Հ�
C�此*��3�$U�����������	�+�dY��|6��7X���
�W����su�v�;����u�1u!E���)�F�uZ��� xl/���`�Ok:����C�ލ��s�g��}s����uo��������y�����X�q������7y��8�����?1W��6����S2��x��@*Ae�t�%��X�%S����.��l#O�qW��*eW��� �ދ��z�{�!�V{VҴ��J��:T�h��b�t�T���k�e3�����lP�l^�t�zV�
ڰ��ȕ�o�^��c�ʄ6�Wz�.CG�9��&?��չ�3$w���r�iֺإW%ۇ�ON������/b���.v���Oz�3�_8{��9O�XxQ^���k�R������K;������L�c�;t�����亪4=ʃ��"��;���4�i{*�� b�%�,U�<���{��㯢[�|Y5�NQ��.�iu+H�;�r[����WRr��5��n�@8�x�u�aG�(�t�[J�^J��-�%���ۆ�
��i�w���@0��k9V�9�-q
	A�W�8c�-��l�[����c!ͩ�\�*#��ĥ�9l�C�Z�J�9h�ST�E�y�t��"Eج�(C&�<�R�TV��%��=�e^*R_t�8�r�C�3����%󊷎<Y��sE�.���C� ��(,�h�֬�s2w�J�kr l�ӫ4V]�f����z���a�U�]ok����-�]/Z��-)(��c�6��{-ј�]δQ��(��+�!�Rjɵ�5�/n��E�X���(-���,pܓ�C��z*�����A�w��Aڥ[�,�5�S0uv�Q���Y�I����X���'z�#G��9�P7.:,`t*�Xv��\���eќ�e-��k��V���%%g,��+Ԩ�W[!pK�=�W��V<u�O|��+�ݭ��h�1ZU1�`;g�btT��s3%�J
���#����⩠^,DCx��%xu&�"���=�r\\��p��t5T!\ў�Ejv����r��,��p��ӎ�[�σvt�tS�|z�R�;���e>�v��\9�2#��u��V��(�R�.�$�N�G�:�p���d��C,��`D�- X��&H�Ν(3f���X>Qf!��k^�=8�-�edv�W;j�}W��[��It�iY�=*ݒjl�-�c��ˡ�2-��[�n|����݀,[��r�aֆٛGO\濓0�=,ͬ䮤��i�'s��
f��>3��Ֆ�1,��ޡ�	'>���FT�Q*}R��(л;t5m��N�53o/h�AZ�f�&J�Wn��xU���ڟr��Ṽ�9��pə}W�q65[ú��dR��k8-��Yꝥe+Ѷ]5�ka�2��9��d�G8�j8��zwu0�S�Rۮ	�E��7]�qsz������)Cp�t]�p��|�p5��-��榫��[�u�ʻ��U'\1E�a�ܭF��2c�G��r�r\e;U%��ʂ�������}�w8�Q��k�����3������J�YW.)����-�m��QJ)��*��X�bas*�s0�#r��.nn�i�̳)l�5�L�Y����Db����.cq���,�ĶQ�\F䫻���Z�*�ۘfj�2�W0��-*,�Zh��mh�%r�u����MJ���2��f�v�Q(�s13-�S�j%n
Z	F��G6����p�r�+�&+q���1�jVT[J���we73-�\��.U-�Dn���m�[Z�L±B�R��.*ff\B�eJ�E,�L��һ�aEYm[[��K����70�#[1�[j��7wM���mTE�.-��[�Vd�,i�0�R����4��.�:1Q��㉔TĮ5��(�J8�-.S2���jV�Y��ܢ�e����������j>g�wu��%)^�ܴ%Ѹ��V�(Z����;H��U��˸��x{��Ә>��7{M[��<j�p��j*�4�$a^?%����f�m�V�|P����/�z-`7�!9U1:�8"_u~��1F��<�r��(oF	a�Q����Ʌ)��LG�!���c���R*��e+1r:��T�HLa��B�[�zb�B#P�c���c�;ӑ�h^TWk���ůsb�E��df*�YV��N@���b�P�<4z�Wp�
�=P}���@+�ʳ�X��~4�=ੌ��-eM;~�Ѱ='9ҠX�]Kh��'a։\+�T�9�F)�"ꐏk����f��M5��e�܍}W
=Q������j��[T�ȫc�(Z��=ix�C)(zKabF��R���7���A�lg�,�ͬ�y�Çf�=	RzT��|��&~��yV��HxQ������.g���{�W�5�� �Xs�������J��&�y��o�%��^�����{�H�L���V�v��XM^��ѽй���4���v�fVE]!�]7$���.*�}����EWCAq�ߞ���_^&S�!o�B����A���>Z �q@�@���Uν�~|4-�U�v�n��Le2t�F��)|MJ�D��?������U�{��fMQ%�6.��Yv�pN:�����.���k�H�[�J�\kD���x����n=%�wt_?;�X��(w5*������*�r��������ޞ��sJv3�=���c�_��u*č�Q�� 87s��bS�x�Ln\0�EߡW@Ce��r.�k���YWlF��)W�H�b�z����Q���P/5o�c�^��_}�)�e�4|��}���l�=֐CnA�n}�	4�AB���S����=5 �`�q�uf�W�[��X�]��2��EP�^ؓ.$1V�Θ�\i�YC�:���{�d�+̛�Dx{�Xx�2�B�<��e ��Ҭ��-b��v��p��o��gg	��؆�������9T�\KA+�0��] |��V ��2Ǣ�ʃ6�}10=��t� ���u0Ns"���3�r�|+��q��z��&f[Rw���9��I~{����Kx��ם~��5�=3��:yˏ}�|�͎~3��ؖDś��$�ޭ9{�i���V�=� ��-�dR�V�b����f͖�����b���R��ؼ���կ
�}N*��)W�N>���]HץţHo%DF����_r���A��;=�ܜz�mX�f���=�-��׶����y��=|�����a�fL��e��Z5��W)Qѕ<�a
�G�eQ^r[�s��>�uN�Zl��7!�5�3�.�jE���)5���
áM��*->�[����${x�/��.�1u�멧+���Z�x��N5B�P�@����M��o�r�:gɁ#�k�t뢡l�^����u/N���r�v�Z�ws�* ~~�*cgf}nT �L8�-xу�Q��׷�B��Z���wlL�8�vS�mq��e\�2�V����c�d��o8�U������|˺]Q��I��1ŧ�.%�Y'u���¸�Y:��R֫3��ӎ�����cO��W=�rx��?����<�雇o�3���%�_�Gۧ��W�Ss��V�w.���*�ձ�������g�_�{��p9[J����H⫝	�M��eB�ěb1\�#�_���WP��\@�*�@��A��F𷂻��7�M��XIB:3ҕ/ٶ�뻏������r�U�<M�W�ƪ9�qu9�����G�lӲ����z4l�!�삧��i)ƨ\�u�i���EDw�b[����]Ҍ��V;=���ظ�ѱ��+:67,��>nXˍ٩Ƒ=B����H�}m��~�iJx�E���S/a�GYG�8s���V��0mU��:�亳�^�uDe�c�"z�i�naƛx	���OEuP[;e<X}�B�G��_����1k>��9�b�87,ϲ9�@��6U(Ju%X��t�hj�V�����t�����t��:iq;2b��_43M��`��z��l�9�RF"+J۶��P�0[7"�m�ZEǃgn^Ժ���]��Æ��#��#g5����ꓯ�gb"��Z��{,H*�ﾯ4w�R�`9 �U���ܟR�e�
ڰ��ȕ��_�o�$m��һ3x��9H�#n�5?G�_�b�J���n{?(37���׫��Ց��&:���L��Tf���rY���O8�ӭ�n{N~�3�/=��i�h*z{7ܼ���%g�yQ
�y�WN^8rR�_i��~���a�����sE`f�&F�����p7�}��1\$u��d(�����q����1\��qk��HnAULCN�����@��˃h��z�c�d���ڮ�h���2aKx���#��F�M��[�ه��t�x���!9y��z� ���U��i����gR���5�p�[c;s;���D�PY��¾T����^;��R� u!�=bg�Μ�z�!�BXNɜ �2cӄV�	��k��7��i{��`�x�ir���d�D-����r����^��NS���Y�1����2	�[�\|�c�H]9Fyf\ܭ&�2P�z���8+5��DNӋA�Y��4bi��+�����<�g6���/�:ȭ��h゗�d��F�m-����&�����S��F��]Ϲ�Q\ 0�h���}ׁ}���Q�c��i1�B40��a�u������e@a�r8@�jp9�6w��mu�1^8���x+޾9$�%����pW|�
c�^�Z�ԅxҏ]Q��𽋅�`3I����Qj��z��7Ţ�Ӥ�S�8ׄu�*
S�!B����z��iKt��-�\�[úxR����i����3��Y<����"y�\�A�-ʅ˳���q�# t	H4i�L���O��	5KX[���&�q�$lTl$����)�
�E��*s�T4���>0%]������Ϯ'%EB�K��c�%T�yH��@ъbF�ދg�j:���uN(��utm(6uȺ��e�U1	��Wx�8�q_rc�I�Ţ�x�yٓ(x,[�ۭ�1��ˤ!<yCOE�1B��؍�����
��4���
�߇Җ���yLrw v�*48Z��йYN�܋0�n�ʄW����x}���b����(q�K�p3]8<'�v"�`C����'�^�v���.�ot�}�Ƈf��<�0����0�ټ�O�ܬQ�X�f"%�rԥI� *��a!�����������O���<h�Rz��U����:�;%�5X55��R?�:�
����82��>hߌE�&�aD*O�b:=�7k�g�a���k+ℇ�z?����ax[�J˘䖁�;3���PP7d� �:���s�.4�GB��� v��NH��P<|�3�M`n�:���Z�P.8!��~wF�+i9��!V�M���y�T���4��t�!,g��_r�-$��Ob}�6-(~�J�1�Fn?(KXjR�H��?Dʥ^3�V����tYB3@Y>/U�[��+D�t~˳�g�ӆN�Y�;����.���}�{�轃V�k�!�������7����|Ŏ�n)���Q�Gd�F�	���Hu�z�|]�6���v�Bmj�PwP�p�7��8@R�ge��Q�H�*Ǧ�o��2q�	Ҕ�?>�����N1&;�,ȼ�r,gPW�Ԇ�ũ>uZ갬:����;*.�D�(������po��ӿ]M)x�(�jE�WR@j�ġ"&]�م��Y�����A��*��ij�9yhC��!W�����q7ڇfh�y��1�}�%�D�Þ���&=P�L8�,�FNz�ì-���)s���g��4�޹�h�9F�d����<���nr=�J�&���Iy�u��:�]t�%�"�b̨��	��}s0��΄��α�/�o��Q�XLo(/���3�����8�����؞=�꽌Yz��L�_J���P��s�0��(@��IN1�eG����2s^Jy�ذ���.	~��Q�l�f���+�^�q[7t�=O��J^�M3�w5��sez��@���������P���q���j�5e�����Vv�hHbZ���x�AG+��A���[T��,i��r����cI{�;�̏vKё�q��ř��=b�뻎O�i�s,ؐ�5)�ə�hp(> @�28T�JOd]��w�x;���c�ϐ:k��T�r�j��B����~򬴠��
'"ӳe��0s�l:ȭ*��N�c���֥/�¯��m�9�_!�a��e�]�u~�
�$>4����L�e<XX�m
-����[��G){ҕt[sB�WO���/hl�P����b�:.Y5I��֋O��P�T����@��NG�o��mXnq�dJo?mw�#w����(���(*�Z��Ǫ��~*
���`��3c��uwWh���9D�ܱw[�Ύ�=B �=](EL��z@��!l���KH��
j�!��}�N�S�Syx����%/u��y��a��*���޹�&�=��7O��Z�7N9*�>� 5*�p���"{����<�d���=f 36ʋf�;!�U1v&�8f �����ռ�X�fb�𚲴D�N���������s�
�ٻ�A_�U](���1TˠRa��*tQ��܌��J[��#uedyЛc�9d#3N���(�ѱ�jX�j��23g�����o���੘S�T&����u�0��WS�a�hd���֧t���O�1d�b=c¶��j�_�/Z��b��= W��joc�u��[Fػ��=r���Hq��z���cR�ɧ; ruUP(�A����n�=]5xz
�1�g������yċ�~��nm�#�)�Q���Op�6��֫�U����.���
X��|A���{�^���oD�BLl�W�ܐ���R�\P��hf��x�6Μ�@�Pe�����S����FF�BG)~s�l���,�B�]��g5X�m[��+��<C�{Ԗ�������T��'ܣR
3UVajT#�t)�7�'�e�;��E�@��ADد>Z<+�n(>���mE{佥;��Qq�wK�&)��P5u�"��@[���O���ޯ�lu����p���+R�VE��w���clE)Wy�t�"Mql�E����pU�^�r�Z6��Yݔ�fU�c��t��Q�;���R�R�Xӑ��E�S�6�˶.��Ƀ��XQx.�+�T���e抾�����m��%�����Mb�'J�y|�S�
B��g�W@G�SMem�|���͎Z�3��Ŧ!�� O��ݫuh�]LU���<a�l��l�-�N�D��RX��f��y�-h�Bֻ6&]�#sr��
+,����B�NY1խ���.��"���;��k�3��ui���|d¹�Ht����C[5�{�iN����Kt�B3�Ȍ������ě�P��5��9���.���,踢�37$� s⬚���X4�nf[qsGBS'qy�0Y�	׶�ꤡ��p�k�`��Mn@�
ی��R7xp0�y�C��vb6�&t�[O�&m���y(��w���w�V�lxQ�}ΚQU����"pW%-6�Ga�6Fum�GD�ͱ;�[�H���ї��29z�����[i��F&)�{��ڷ1j������j���ɸ\ak%=tfb�@{́���j|d�q�-�%�<avΉ2rU�OeJ�[��ݝ@M
5�Ӻg��z���J��ك��R��Vq��]b�쾛�Gg*e4�t���
8c�w8�줻5�K���n��L��B '�Z�e�S���5���֥h�0U�W]�Ƣ\���0QGݚ�ai�N�'���tLYh� �|�4��$ܟZ��R.Av���r���c+sѶ��F�Y+E!�du��9���/y������c�nh�+�$y�,__LO :�g��V���s�9�j*	iP$��0Wj���犘�2R�Y:	`�N�
	c6&'ʻ�2D��'s��݇R�-���>���w���K��ӳ4���t�@U��o(�%ձR5ʻ����6��|V�Lu�{nWK"#�(�H��t՚��u������N��vb�;׏qb�ј�*%�����A[Zѳ-�@�;��6K�-�;]87�X�U��TY�9��@�'�����T[����s��<�]��;b���c�g�k-)�\���e�˗���R��ܢ��k�3.�2�9E�Ը�c�����jҹ��C-�S-���)A����c`Q֊�5�Pĭˉ����5kp���Lj��єu�j;w-�����&�Ƙ4E�S,(Ĵ̳v�]%W0�-QB�7�ˎ���$�� �r�F�w-r�i���2�Pr�n�ʨ僷.U�w.
�"6�qK�G]����mL��cSr��\�q0�V,�f4Q�MŎ�V���˶�70��ۻwv��9swfPXQ�v�nm��nM2�*�R�9��F����[�F35�S�1ۮZ[��]�b�ѩ�+����w3�m0Ʃ�F�F[3�-M��խbk��ݦ�nZ.�f�K.�t���������/[�b�Y���mk-r$TT���L������K>[���p)=Y�|^��9���2��"ʋxMW�]��3N��c깛S�������Vf��FǶ�����0�����ӎ��I i���ߪ|\�Z��M��ݯ�bCsFF����p5�n;���]O)QQ�dӀic��J<�d��nf���D�q��@j�=�ϯ�]��R*$W��mVsƞ �DÏ8ڪQNL]�����lk��#\�t4��"������zަ��@n��6|`������4��~�5¶�p�I�^�M)c���\"��ɓ�2%H&�(����FA��.��|���=<-���� 5[Zx\�E���4�����C�t��~�W������F����X@E��(z�@<��]!V��)`D�ˀ�Ê<x��4�5�,9�P�|��Eǐ�#d���MzY�Fh��L�g"�d�uF8�:c>G�/����R�@u�-���Q́}YחX���=�ql��x=��r�Ɖ��l3(��^D�8��}�m��L�=vr���M�z� l��b[R����C��A��p>ؑ�/�r�.Sb��bv�A�*�k�du��9gd����W�^�e�&ȏ�Eψ�٘u+��.���d��j�Cc��{iy7�.������m����^��(T�M)�T���]��y8����/>�����%��;�.������ؽu�(KXe,�h���_�ht���L���ӻE��FL��t����������$h�_���?n�V���zGRq}N-��s�}�$:E7�����B���
�����pXV1�S�(9�M��i�$81��״��X��)�Q�Ԅ1;ʜP���K������.�>A�"����3>9 �t�	y`�g��[5�.���vn-J�6����%R˫�'�'f�Ϝ��dÍrɣ%7�g���>-b�'}�vw�y��\��x���'��t�ys��Rܛ�X���=ۥ1����X;�2���E0\���1VP�1������nP�B�@R��W [Gl���>"���Y��Q���HP�B�ڴ39E�[I��������r3�˗p�k/-;Ô�.�wY
YʬN�D��@tड़�4������~W�URG��=Y��~�9t�{w����az���e�Ƃ1^��1C����r�B���)�`��p�~+UQ��������P��+t�S��Ğ�ث�1V���!NC��.��tn������h8بC����ٿ	����}H��AX=U�u��X)Y�M{2ݪgƵV�PC/�]b4���qK�r2�~ȗ#|���$u	���*\Z���iŌ�"0TS�ݔ�6Zr6k���("�n������k�O���1Ks���W���m!&+���(&k!u�_*ӡV�S��Q��X}YK)���@q�̾�ˢK�)�J����3��fB��箴/�.ǉ�9�aNe\Z��S+ �Q��:3�]4�%�=WԬbT-��-U�$�c(�`)qLw�mː�жr[짷�f?��������:2r��Bb>9,b�	�}��47�1�X����5�[E�w;��Ⱥ���0�DbkjJY{���{���څ�(�N���l@kir��qD�ЁJ:�rR���}�}��������+�%���^.�V󕦄����K�NAh�z���<6L��P�����6
��O��E�����t�=!+x���;�J�8B"U��X�L%Uk�cw�t����a��Q�ƥw5,h!�BC��5��Vݙ������0�eg.g
$!�a_�V]l�m�ۚ�Վ脞�k�u�zQ���Ws�&/�����+1U�U��^����Y�Z�9A�Q#��p����t���x�[��Q ��q��Ό��r5���i���4��:��W���zJѱ<�GԺ�-����(���ζ��1��3Ú�yԈ�h���q��ae�;I_l�,H/�\V�L�
2���E�Z�4Sx�<LӸ�I��<W/��{N�j��I|���4�A}���8�D� Y�
ǯ��Z��+? ��������E��go���-�<�q�ۥt�OD>͕�qK�%���J�9]s�q��a4��m��wٽW)cNX���Gg�bhv��h�2�?=-3\&5c>��-E'����i�[!��(��D�,�钎TፔU�G'u�֫�խu�q��Ȏ� �(O�&F�F۝Xot�/L��jwi[�8���ҹIx�4��X�m�z90&gѦ�7t��;Е��-�E�J���dm��T!�n�;!��{DcW���\7Fa�b����HU�ǠR;w�HoV^��g}����gp\�浺��*ܬ�LW���2�)[�E��Rd;��4���u��2zع{Z�]]�-�ghԙO�v%��Fh�oN��u�b�S�D墏5�*����:6�$���T+2i��i��u�UJ�P�6O^,8br9��º���i��*�J����MnS�ք/�G����W�Y4�r�|&]k��%E�u�c)��B��'��#��Q�fmp�̱ܰ�Π32�>�C)ѥMx�,�Nlۊ����1��Ne؜겶�R��$aU�ګY'�E1��}$]��0��Y@`�R�X��{\/��'�HE�ҭG2	�R\
T�cŎ>���A�M�YS�G)�F�-���Y-��鵹���f(X�5��'M���t�*5G(WBZ�9Υc��)�)�h��F��o���]��C�14Vo��ճ>ri��E�S��Q;�ឲ��Aa���I�;��I[]CZ��IW�αe
����h�y�<K-X�X����WӼ���>/7	�彵����)ٙ�Qf���ٱ)2a����o�m�]�*9d9Ό�mA�ӉZeۮhJ��u��e-+d����7�Ũc*L�����W��2��x�}�*�W��(��@1���@�>к�$3Aix�U��.8�H�B9u��[�N8u>��0�b����6����:V)/Ǫ��LJ��㖫(���:��r&/i�NJA��ؚ:�]+%�3��^F2hq����B�S���J�{'���F�{p:��%y#�(�R��go�dB�Ү*7�ӵ�ݪ}�X}���e#
�F�/�6����s,�۵�/3��y52��w.J`�7s�W�Q�fℭ9Y�i?{%7qz����x%Uy���6�Y�_V�Fz4!��q�x���0V*b�����5�jY���W��X��[\q�Hn4����Ү�P�K������O�3�Cy�1�R��c��*0����Guh�6��)�*�t6�������o�v�A3M��H�CY)�����iD�X�^-G��u�9N�uŶ���keP�В�)��gt��&�ӼI�a�v�#p}���J�����X���VT��vyv�.��fz(���~%YO`�:�sW��~k��Kd��_�{/=�}�LSս8���{|�sMDZ����.�9��-��W6���I�3��M��z�(C8���ְ[�}i[��$GD��
uɁe-}�j3q����|T7��b�Nmٚ���x���l���b[��`m�3#�3G�OK��]!W�z�����b�ٶ���6���:a���|�r��2��6��@߀U3ܖ�*3y/�T``��rQXkg+��B����v�y�FA��i^�Ŋsx����DL̄>����������Z�}Ȥ7.��:�b31C|�
$�~���;�ӗ$|u�=/���5���[�Vg(����MY��F�0�Z5E{��P�T��̷s5�orv���X��tz���R͹��4f���\K�3&���K���C���7��Y�h_Y��ts:�"jFɾ�TGHH%ss6,�C\�4�.��V@&�='�ՏNoh�:{B3k��T�/vܞا6'��<�1e�)�I�6$P�#L�~���]�t�fqS���hFki^�M���(���,3V��_oY���$�a�����Pֹ�m���A(_J�z}Y���u�f�
����V�}6{���${pe,K/5��T��E[5�6���^mn(��-J��ek�]!X���/J�xw��jk�;GaS��u�٩)8��閲ţ�T�y
:h�C��ʟ7ۼ�b��@R�;:�:R�g��g�]�����*2#x�z)kT�=!+s4�_$.�̺����!�apg�:����1��뻭s�E^-u��<K�:u�\,rP�çw�Bz���Ѵ\�&�v�2����کf��H�W�ā��Ô�ۓ4M�}�Ӕ[\�F�S��G���#�5z1F�����w36����~�W��Y�Y-��@�����R�ek�����Y������t32�m��4�6��$ʑ���t�eݳĄ+*�씍�fFj�y��P]7���0�����*zi�Ef	9�T�VU[ھX]��*�7�~�o���{;�Ӛ̼��*��7��й�=�ӏ2�Q�="&V 2��n��+D��m�)qT�r��N��t��0�^)}\�6�
��Uu����
M��n�T��R�v�5�&֊Qo�<YK�1�6ws\��ʅI-�]�2V�,3:�Nwmн���.ڬ�C"*�P�Ğ���5�8
�u���R�1�f	��M�j㊖����Y�ԊR:+H�m1��/"��\�C�]©�m�.`��P]��J���ѺZ �ީw+�Qq7��H�;]"��g%��:7b	jK�Mg��b*�a�rb����Uݜ�k�d]F\>���ݫH�*�;�,�},��<�	!˘ �RӾay��<˖�� L�>4{m`��A4����7��꼢��'yY�0����{�|��X�T���:��5��Z��
[g�[b�'�Y��#�Hp��e���):I
d]Վ�x�����B�ѽ,<4� ��q�y�WR��m$0�3�B5Z�D�R����TGs�1*j�M#+�g���/F��ͥ��E`0�꼆����[X�N�D�Xs�-�R#�M� ]�Y��vI9��}f�#4r��X�R�wX�Q��=h�b���A�Q&�3�e��I�3=>B�:ٽ�ov��m�o��#�8�bojKn"u�ּX�}�GV��e��N�w|/���Զ��(7��MZ�̠��v�*��k�'g^7�xML�Z���*ȃUs]�Ԩ-;?G��M蕘&Gsǎ��B��5��"��G]��#��cݼ7Kk��׎̤������٬rU�KZ��j��V�sw5�S���I��^�	L���{�Q-�V/`Z�R�]�qN�����*����\����6/8����0+���hU��GYR�wy[N�cq�n1�!A:1e�x�e`���'�oN�Z)�/Sԩ���ޭ)B.���	�b�&E��,4�疧\�;ܽ�2��!	_H�>�}�o�WqA}tl����-�}}����4R��h��[ˏs��i������ݷ��u.����eؽ�k�ɨ*�k��=���|�1�㼩�_@���ph"��m�J"r�����G+��¶�U�.�3ʙ�-��zgU���T�D8q�q�^����w��}�!F`���h�(��+7�˗,�9�&#��[K��q-
�%m�t���mk�c�E��L�`�̘"�eť�Q*�0�6�.4�����nỗ�̘�8��&d������BҪ�1�p�[Q��s��eE��3G)�c�3-��8�J5��aYs��mU�-pQaD��9�3(]�Աѕ�ݵ���e2���Ys����\��U��F,�1�)��m\�����e0�S�q��u��zl�m�ʙh*�Uj1
����[.a�hԹi��m�VTLp¦8˔�YX�ƳCnf��J�r����*b��bZfE-�)�[qm��e�q�-�jfnr�
m�"Z)��.�J�fUC��yw|��޼�W�~sʷC��	�W��R�k�
Ύ�"�S�3(z��q�y���&�O�����W-�Y�w���t��⺋f(gje��C��wboQC�ۙ��y�3�_wS�K�ʹb�=Q�te�ǟ!���9�n!��.��,s��{���Wf�!��lt�C�&YT,�w`�J��V�DR[�C6�S:���[:����t�]R\�4�����x���q�`ĥ�	Sx�'���ӌ���ɖ�Q�6��-�~sҬ��O�P�������#F�gkT��G����)g*Y�f{~k/Ϙ��NXU��W�����9�c(��b���KD6cX�eW���xe�:�V���a��+3��ک�m�J�#ځ�(^Va��t��v.���Kvh�Y�Nؐ��S�Ȗf�O7U�ߟ6��v�9���ی�*��z�맀I���[��BP$/�.+r<yQ�]MgzP�y|=�x_7�J�.�>	DJ5Dc��xREQ��^{��Z�k���~�b���Ҩ�H��v�ڻ����	Ľ�v"\GpaӬ�	��kQ��:F��L���߮�mD SM���$����H�'#�*tF�+9y�VWV|�p���=�S���<�+}B�HQH!���I���J�:�2��f�.���w'��艉,BHU׳7�\;{�}���
�(��W�
�߲,���j��GwQ��m9b�d�����bS�L�#�TM;�q�����66�Lj}cS�m켁 ��BD`mQ�˃��oZ(A��-�n���v�noؕͥ+�^Ӕy��������x�R7��m�l�#�(q}�f�q�Z.K<�&�QCćn�ag�}���W��V�f�q��㺢֬*�Q	���f�2�3z�S.�P��)���ȋ\�͕��#ךJc��31ٷ�M�u*}OI��'�[r(��$p�8��b��B�F5z鞝�Rſu"K�H�36�B
��	�X�X��o���\F�dEev�NP�c�9�;*��l�[sW�5��n�.���q��L�،BGqH�Ι�hJn��M�a�k��Q��U�Lp�1�N�Q^�TF��V�ӽ5�_;�{�~��{(go��.�=�4U��5�Y�RQ�#�9�Wμ.X��$g*r�о�U!�qt.����	���E|�Vվ�8Y��8�T�m�燨�+dc}Q�ôyU^g5|�/v���N����FmI�d����(�S�on>�[+� /�
ӥ0�K�� X���9|���<��7n���řҟ\���N�{CvgQ�%�:��ݎ��c7Ie���iG�y-��/�?�x��|[�7_=��'8������u2EN�-�t�J�洢6+�<�v;�E����(��7d���ˌ9E�Hu-�z���=�w6r�{/tG'u3�Q4�VG�ϐ��s�y}Ps��V��-�ʹ�h<t�w&�b�{��&F��nV�mɷ�wx�ˏ
y�*�\��wF_�5!<�x#S�M�Hƻۮ���2.21�s��*J�/kǩ����R��T�4���7���(�,�LE��\��UJ5j3�c�l�9K�C��cU8����d�ݫޥcD��uG�S��������a斤"��4/�Y�W�ݎ�(TH�Jш�͞�hP$\u�4Zʫm,�˝�:*^��\]���->�������)Ĭ����8v���Y���|͍/7gC����Lj�s��GnP�����]���[MA�_e����U};s;�m��9��V�V۽�+-
J����[���q�he�P��N�U9�鬹y�§�gqN�����ܧ5aD��B]+��{\/�H��C㨮��V_�ߎ�N1.���/%�*�)��#"鮣X)H�8�{�b�z�g'�A�6�������׈=�N�N��sN�'D^�s#�u�HΣ���<�)햌b.=ɒ��V�!mJM.�n��R�l�:��q1CM�z\��a�vKe`�5=�꤭�/�jh�f
���T���.�x�t�s�]I�8��ù����$��]|ŧ@�P��P	���1�츖$1o�C�SN5KC�e���]!�X���h���"��C��Y�d0�f��M۶Y�NKR�f�{�lŹخ�Ӑ'R�?9��+���.h飛o*4�R�o�G�G�)�͔�����URxI�1�5ϻ�qK|U;NC�h��Oh����
�p�����ѵ��]3��(W�Q@�yf� �tc�zp����C��X^륢�fy�a%{/;�Oo��V�A���Y��ջ�m�JQ��P��u�7�0h0�<�
��S�Mf��-5[/j�6b4�S(7��)31��5�euJ�oW\�x�seqv�\����x��n(�ѧ�S�;lgA�<�c��{�s�/��W��VX�yVuA����ˍ0����W$�z��Z��I!Hk%2�w]BZE?	CrcH՞��`O�'ׄ��]�ǖҳ�L�8�ح��3b��{���muoH�Y�1�ҧq.����{�� �B.ڙL�(�1�P�"7[�g������u�I�`6q��M����
��:��L��u�DA�>6))EҫL	��.�O��9����)����HP��<$>�\��2z����۰��|ڈ;v�e�s���E�·ƅ��t��=�=��\G���k���ի�����C��q��͘����9gx�7K|�{_^�o��uanq*�JB��#ײ���:����dnm���Yl��J݌N��*w+����P�C`�02[���k\�=U-��}u(ngW��J��F�;:b�wS~f�s�*I}~5�U}Ϸ�b�֫��iyg�XϼdF�[ܱa���o4ʸ�̎摋��ÂSwW�
D@��n�b:1�[V2�m�C�{Lw���TF��-�`�u�f����K���9��=� Ϛ��r�PU��ZV�m���u��*\����	�wS��o-�N%7osb%�D)l���+�U��B�l��e')w٤�K'�K"�C�2���q��d>ۛ�:q%�<!��U��VU\��E��,ؽU�^�U�>d�{�M1!���
Z�Vվ�:�z���G�re�6����I{��.xJ�9N�z�q��O��N���B,����ť�_I��ܑ� �����oFY��Rb�5�˿k�a�ܚ曓�e@��2��faJ��6;�+���Y���u�����6#]՗��6��^*��j��gm��Ϻ�*�̅p�͛��z{�!�&_�K�Y�]S#z�7b����a�-�E޴�!��˾�jEx� ���NϚ���w�����kD����>��h�T�AN]�9���"��7;��v�� R�
=wr��Oi##k����M��7�v�(��{��eٶ�n�un3q�̶S�!�����s6�D�M���r6�zZ*X֜8vgt��s�s��.N-�b6*��ch�讀�(#q\bxl,:i
3��6�[rl��t��%���P�4z.z84�>�l[�I�� [��o(^���U`e7}(P"5D�%%V-Qg{�c2!��IZN,Q"��x�+��v�.��]�M���GM�o*�A�3��4>�r�ސ�;]�2��e�\��T�����O��+WJ#˚���L
4�s��qE�cw��F�Y\�����NSe�[��r����e�&���4���鵸8����,m��bc4��J�4>����U�yo!����I-p8��׫lR2���H/0�P����a¹���y��u��)&hd�5��+w[r��
+��E�Cٵ���Λ{�名�]Q�b-\�\޳G���X-e������x����[�l�X��f��C���I榟W������R����m��&X��]	�����u	l�;S�2�DV�_�6��!��8UN�%r�@��}R]I��a�aJά�U��ڈ�e��R��G;s�@�L��C뜾�c���/52��8<�ݭwup�u-����p<:ı�"bbku�V���BJ��Ѳ�];=T%�P�����T>7]}ܔ1](�r:G8�Ĭt�h�����"�V_Zd�b�7�儧��u,�7��jh[��m��C�ˌ�ݞF��m�ǌ���ПY�a��[8ՁW���-5W�ٚ������퍿ksD�~j�����Ne���2�?�qf������s�+
��Q[
��N�͍���0"��R�,�xLwy���qK�Tk.��ҕ��q�U�W��:�X�1��君�o�H��Iù� �����&�)h<�TC"�RC�ы���et#��q�A�x�f6{GP��H��oc+v�P�;|]�E*���J�=v�V�Gp(��-㴪^�}�&�&|v������T|�U��n�KFI��z�_1��h�W�c�f�]E]�id��=J��5y�R�6:��[Ԋ�����{Vj.��J�y��Kg�w^<���*��05�O��2:�^����Pxڶ�^��o3B��èT!�ś��t�Fe�I�}+�m�����;��m�5�j6�����kE ��3����j��P����]Z�'�WBE�Lx�k��\�ǅ+�*�eF(���d]�7���*�-�0�g��s��*�:��/p�J֌!N�IɈ���]�܆Ю�i�-=6{;���{���=-r�+C,n�U�]E`n�PB���{z�"Ic�뛗`YjBA���+
��.�V;���s��]�n;�Kz*H��l�.�8+5�.p0f�Ipk�o�呌I3I�r�� ��[�x�3P��ܚs�0�e�i`�K��(��U����Jʢ9�
���o���=�n'����*�u
!a9n��}ih��2�x!��P�6�8�)�ٙ�լh�Q�b����@`�4�(�Q��,na;�F����)���5���j��.B��Zd���v�ً{,�+6����!rV�\�Z�Z�OI�6����w�yOS4�Zs6[%
Fӽ���o�%R���XR9{䎭���7i{�ֽX��5�pm]��i��CحlOj�b��Y�tK�֤8!��I֝��4���m$�����Ut� �(Im��7�C�S/���-���Z�,���p<���%3��Z��&2:Ks.��ֻ��e�Y�wNT=�!,?X�v^`�N��,=]Cr�7K�W�%M���@�dM�ffb�n�t��e�[e���I)b�)�Z�,A6��H�늸9(+����E�R�c�(�����΁��c#%c;�˝O� �*�{Vl��A��w�kǱ�rO�����V(U�-k�""���3m�d�T1%�J$Z��X�3�����e�J�(�bl��[`n[l\Lpq�Rʪe����h�[E�.5ƨUm�j�2�ZU[lkG75�f��W
�Uũm��"�e`㙖�1��5�k5�����Hc�T�P�l�8�4�����(��7)��������Tm�$�-j)�fҢ�&\qd�eAMaX[`�R�Q�vª
�)��5"Z]�3K&eX�(��b�;q�4G,j�B��P��.%V6�J�k(���Ȥ�*�+.SY��d��Fݶ72�J�Rڂ�1�hc-���[sҢ��m���Zcn��b�,�jn��W��,a���������O�oJ���-*ݼ#a8]�c^m��(��-*�[Y�7F��rt:s�nU�jߧ�;!͑�ϱ�מ�:ti=s�m��奓�0Mۭ�z��yȃ��V^+ʳ�%o><qB�u��ک��7�M���j�^+!��ۛ7	k/�7e�튾�e��#����sƮZ}d��[�7M�0��nO<{g�!>��BFm	�!���i^�"�iվ��dk{J��\.z(� `�V[z�<Yj�S���$���^�K��ؾ���y ����0�q��֢�u�s]�ii�֟wx�V��J���.����m�͇��FY�6}�ְ[�o��[7s���x�KA�����ý�MT'@�k\��Cղ��\OeY����T���x��􁣙KmgV���a�A\��*����^�ϥe�XeOvn	��)4A�J��WZ} �䝾�"����0�F�ЁJZ�r+��ZSw+�W�*RBq÷y	A؟V5cC���SJ�^M��s<6����+�����ԱN��T�d��!I��.#"��uX�.��j;��c&��Ò���i�X'���;��еN�^�\ i��&٨�8-�[S{��A�q[/E���n�H���zT��+����G���,�L1YP�rF�8��8�۫�2��Nr��4+f���,t�U�[���������W��+��Μ�w��TAζ6�vv��4'L�Tmy�sU3���"�#�\E�a��}��ig�[78H�S$d��x1���ɡط�M�8e`�T�m��� Y[U�"4�]:���>� ����+8�{:KD`�wkIt�
�b�	��t0)�*��7����>]�]�5a�\�T���C�%^�S��f=��9��p{��u.B���j%E(ӭ�R��Y�evC�j�Թ�}���v`�C�bv�����H'�؞7�R��VuG�V0�V���Ǐ�%n�Q�3�)��\ ���wKZ�d5=���@��}��6�l��I�=�֦�=Jo�6j���6�x�+���Z�<�TŴ�PB8t�ހ�c�]�&�|�=�KFΌ	;���taV�kh�tC-����K굱�b˚��c]-��#P�4z.u�x:E�(��l!xE?:�bo([Un�d�ç�J�����{w��V��Ӵ،�r�׳2�i��4e��`������AN��h.k��hz1p�ˌ[mm�����ܔ�m����&ԭ������j�Fo���:��E�	i�Ogʅk�F�*��559A��\1�ʹ�	��m��5S[˻�I;rAVsZ{�򬾻���z�gߋy�>~�|t�u���bN��3��㡷!7@�)�D��R�X�����2)��E����ec���Y��ڳ�)�D��7M_ob
֕�m��c&�s�ok9.:zzmo��͘�6�rXY��7PF� ���̂WghΣc��rI����067�w*C*̲�0{doT�)S����5����8,�;~���O>��⪳b� �+�q}�`K7�e�[�=�O51���~�������<}�ϪK�&\�L���V�t'���������*�D�P�����;��d�6�T���w\���n�8UU�ȱO-t)�֍��sHxk��z6Wk�b��}CՕ��n�gk;ge?r�GD,OxQ^N�Z�j�!>��!����)qKl��\n%���c��d��k��;&Rv퇇�� QuX6��wQ��E��P�<_��Ԣ���ô�i�O$�J�6u�ILȻ$��{*S[p������yD�Ƭk���dX��t��D�,�p���>�R�ymN���6�N'H����E)��b=�w�] �\��o��;WwJx��XMt�ռ�E��0�v��ڔ߉J��EM?ePH󫫲�4����OJ݉�[FKm(ճqDsq��z���-%�eI| #��r����>^�LÃe�l9:�rNP��B��1��*�pY/���;��(}�3Kr���s��kz(X!Q�{~	�^�[\�Vc��V=5�Q���%�S�=�hH��7'��Ժ�U�����|�F�79{/q�h��z氯)�]G;]KӢ>m�[���h�2�o-�b��gN��\�:o�q�l�&�9IN�����Z�`�����](C@`U�i�df�����8O ?�yb���-kwۆ�����.�o8���|~��w�տ}׫�{/�ܢ���}�or�4���b���}�M��e>Y��&�nR��HcNz�~~���z^Й9���k�o��n����s:s9�b���� dp���j�21��L16q�bj�M#*J�%��,�RpA�=!ώ��4p�{�I�WǴ�B0V�5#9FP���
����a7R���)=�|$��>���II�V�W:u�T�5"�G{C1W����)��#�Lw��s���'����:�������̗�C��t Y^����i<������M:r�e�?���D�j�R�B"����=�QW�d�F�H�y.m8k�ۋ5DO2����gSS=���u^��V��M2k�\��5��N�}�b�*����vN�SM��������8��k�+p�r����U��B���^�qď��h"�){���2��s9<��-I���s�mv�)
�[Z*�	���@��>y�ƫ���,WE0�Vr�94;gf��+��$npޛ������Rf�8V'�7�9Ҿ�M���(�W	؛�w&�B	��]r���f���ƺC�xs�*��[��c*L������t'�_T,�I'�}���m7�X٦5s|]�Kǟ)]Q�N�ȉ��2&��XQb9.܎���6Ԋ�2<�N�UU��ǒLF�6��w:�[*X�Ӏ����A�V�������OV�z9��täv�d�Ȯ1B.M+53B񰾹k�ʵJ.m���5�.ӵD�V�	1��e��K����4�N�mjˆ�ҳY��rA����b�/�l���C��.��\d�.f��m��k^�-��	�n���Y�d6��!�T�R������)����X�.�F�Ê;����򵄾l1�[� ��77�-��J�)�(Q����}��|��+��w���T��m$��yܭ^˔m�걭'�J`��74I��PФh������{��E�t9�e�"�m`y·Zk 9Ji�VV
5*�l���W���:ya��
��~{5��L˕��z-�4G��FWS^�v{�Xh:���&�CaNF����Y<6��ϕ��*Q
�πue��J=����&o{#��/xJ��<�ٲ�P@�	�$KR)��p��ME��ל��;M��q8�]�#�XeU��{�(��U�f����]OU;ћ*�����-S�#g
��ϔ&T���@5v�0�yS��*�{#�g�R���wQD]��%
.U���n����W#���,��b���S7:3KR]���a�%G�+��m+����Ϡ�͙ڗZ4���$�iZ��l�H��G:��61T
�#fOhh㇎��c��J�Gj����wZ�*���0^�j{���Pa�,t���B�v4m+�N��,��xU�C;ڕ!W��;���ހ�McW����_^�XI�,˓M���b�p=/2o-��w5|q��j�{���a���ܒ1�x�Q�m^gM7���_4#�R;Y)�]�I)�E���y�h\���Kҟ2�����w6���3��)j'�Ɔ�5t5�;�;�Cj���a�u#J�C�����<|�Dŝ{��f��t��/ٽ)^Z�]M+;�m8�U��إ� �]����{���r*�m�p\��%Y]��o�t��9I�;n�|�yWى%ܧ=�o����a��o�R;y+7v�L�y��"�170�\푂�S�����kL>��q���|U�Tf��ȹ�4��='C����T��Ǜ���Z��Kk��`hP�{��_Z���;��Ѭ6r_R�j�-㜅fz(��@Չ�nU��C��`Y_|����Ϸﻆ���oe��0�w���o�n�A{
�.}[�-9z���9�[��[OB!b��yCSҵy�}^��,�m���YoB�uS�Yշ̲Q�:z�V�)��X���P��j*2���N#������Qoj����a��oø�v��������(F�S`�`MY�`�)�����S�}
*�~V�:p*$��_�e��[l'����7K0��|��S�n8�=u��Vb�!�.J�F&��E��7#6浦mТ¾k]w�����z�|�sK"ە4��u�[V���]*]Nu|7o�J,y}��↍#�5E��@����PO��v�W
�%��f��c�*^ܰ�;q=m43�N�[z�o}{����X�G(.]���RoYl������{B�v��֚7rp���ڳ��"Y�x�*��l2B#F�Lk���s�k�Is'9zT\\��B.����Hch�(�ݲ����hQ`Ny`^�]��줍VC��J?iyv�1B�	Y)��tg��VQ�c���l�1�A
?ZB�r
{Ԭ}r�[�#��in�r9�Y��KZ�^�F�*J�D��pś�uc[jЩ|]�e,F�nK�tt6d��m��\<�=v���w>[9�Ib�J7����%�Vр_-e���o(��
�K��T��a�c�����&��4�og�1��饸����H�ڷ�[� ]��ܱ����;a�7|%J��`��>���D��"[�ı���kS>�И���w;*v@��*�uq�^ZG)�8�Y����St��bK�Ë���X7�7-�u�9X�fmJ�Pݫ����#��:����.���=E�{r�-t���Ձ������V����h�����D9*<�B�A�G�ͮ3wHћ�1�4�p�DN��m�rAĝ�
�8�Df���L����H�	-ƚ�W84�:�l���T����x���;�1c�Kgu��lR����|k��aW�C3-,���D���%%Ѿ��V�a�8Hܙ:��n%].;ڻ%�sU�N�E�gK�ѡ�E:ؼ]��&��%�����EL��:�;�c��́�J�e�6{vfE2�]F�صwt�إ�Xs{X��,1�v5�u�Y}oZ�V��if�4���)�v�:��u)xH6���r��&
y�^bڼflFb+������T�կڴ��c�5Ǩ��Hl&a�^I�b�r멁��/�U#,��NaeMY�<��2T�V�����q1�r�ֺs+RM��:�vo]����s���y�雷�H�CUK��K���ek�k..��B���XT�1�%��U\umK�QօMJ�2�@�cm��%jCnRcb�m�&1H�T1LI�(�\feeAVCT�CVbB�#P�MI]��b)1�)1\E���lXMʰ�DJ)�U��EI�Y��eUX�+)1&3Y�X�R9AH,Q��E-���B�*��ɛ��Y1�TAJ�CS2��Q��*���kEdU�kYm�8˴Rk���X�*�Tc2�*mQ+jTQ������t�+b�1�0`�e�*�Xb�cis2�}�?yә�EN��A�����@�맭`��AǱa�øHj��ڵ#�b,�W����xINS?�<5���鴨{)��e���S퉾��&2��� ����^f��Uc)���1>�&����������eB2����)M�̖��$e,g��`9{�Ac�候��)�t��Ͻ�JG�������u�?Z�\��[Y3�5vA��T;�w��ӫU��*7Bɖo^s)DY����mv�+��ފ�|!X���*y�2絶����]�&��e���6�q]' lP훂n7v��h9��"�k��l3����Ph��Nȸ�Y���������S�P�1�Y�gc>k�5��1gT����켎���'�Ư��g`��R�WZ�^��{�8�|�Z��/Q���[�Pݬͮ{���p;`��~����b5"ak�בK��쮾EG��%��2ve&�D���N�Hb��j�w�.���3�dk�dE��cI���܂%�h*��W6�� �R��F�v��fh����ˈ�e��K��%NymH�L�rvg����On������p��g1Q�u�n�TŀӀ�ڙ��0#�KX�0	+ֻ�6�l��'�PF�q)�Ħ�
g7��/a��S�pWH�����t�C�5��-�V�˻��4i��-L�v������*�����:�Ƙ�#S��VFT�F��ш�u^#&3�{��i��S6��5[����;87lVǵ��e�����q;ٹQ��p����$��tv��o\�ڠr�� ���F�+�O����Hv몬�C1b�l�j��^՝@��������u��"_�؂��a�:�jod+F^��U�l�@�h[�u�B�.���;fk^���	��D}��G�#g�x�%i�o��dҧ :�u�:S�[ڒZ{5no5%ک*ׇ�˰M��r���鵱�Kj�M�n�o%lVY��a����U��y�r��C6X�D�Z%�=��ͤa�#z����d�"�̎o�,FF�z�i]a����~��~�:����
m�U����(I������֨bw6ҹY��5/"���v���(q�%�2�@��V�:���*�K�2C��fz�<ay�����Zmkw��b�Է�U�ӣE���2^ql1��h)6D>&i7~CiX�N��귝Ȏ��F����cA���a�7�~���&Z��#�Is�pZ��_JJ�;ቅL,��{+}��(ע��>+S�!�)V#�k�vrC �-mo�:����Τ0Q��/͑��I�����髭�j��fcDEӲ��W�gY�7�s��]�#�O�R[,�EG�m�䔞H��g��ȩ=���E�ܕ�%Ux�T'u���'=M����o���uci��B�4��R���u(�/�	KX!�mg�>Eg��t�����v?�{�|r"�6��l27�]+��oE�co-9.a-��,�L��Z�]>�Va1����;de����w�g-��A�a���$���U��Q��9�	�*>��'�����?]�뇺�^b��(}��T�ڞ
�t��//���m�Ÿ�C'����J��o�+z(�'5���גu�y\'�����U���ݿ}ھ�m��Zv��uw��"�b��3�auJVT��O)�72�V�=]���3^�3[�е��n\�Lvu��śZ»"�����<,�Ws��k���Y70�]��y۩����6��;�5���B�`��hżD�aZ����B�8'P� �ZbV�!�̈́�{��;�fau6���T��%���sR�|m߱8	g�<:�c3b���<L���1+���`�T�ESqIĂ�ͺ��݈GJ���Cm-6h���+��q���=���{˹c\mӟYsB��Z!��rZ�d�اrEm�H1x������f*�J�e=�8o��B�	A�y�OYV�]cn������M^o�>�ᔭ���6Փ�q�~�}'����׃���7O�^6��z���9K��x�q�Z�i]vY���xV`��-em)��Գ����b��>�T�l���V�Y�b�B}�/;ˠ�=!���j���Tk��}�;]7X
 [04Iۻ�&D:�C2� )P�De4஝&g%y,Z�5d!^�[3Y�},��Z��뵪9�
חu�=;�<�.G�E�{������W:~��h)5۱io�~`���;����Z�3S(T�[@�oNX;�E��z�±�ZM�U+���2��-�}�c뮣��c�_v3�i�� �"K���Z�)켎���N8�L-�P�,�ީ�t��7kQLx�N��ͥ+�|Y���m]Kǻ�KB6t�{[���������W��A��d\��B�˜�}ͱ�L�[Dcv7]ν�ʖ5���#q<p��l��6�zC��^��6�6���h�����Em�M�ւ�Ȕ#e����^ڱ���|�l�ޙ���+�?_��6�:�;�}�LC�}z4z��(��ie�����xG^w�^Gw�ӧ%��2�|�0r��>֍�]~�,p����N$٨9�V�3��Y0�\#���RW_=\�y`�r�W7{1�^�\�(����=�!Qp�Ԋ�;A�;��b9M�FLf3���]LB�#�n�J"��F��Ԧ�3_{�����H�pˮ{����,#}Ht�{�~���7�WU��J�� ���k����6��99���bU9��{��*���^����<I#�5K�N^��u-�=F���8��^�lSI�&e��Z��V��F�'�h��G�r�tй�2�:f!u]��d��. �[�)햌p@�	����S욉D;��V�w�J.�?c.�8�\.���C��`��X���,�y�I�	�y噕M[]CZ�N��i\�a�K����s�yry�u�="�9{����ts�a�����Gk�
AE޻�w�t!��V�H�t�w���k��xEzv����*S|��v�K���(�M�5t�\�6��N���7j��������~�����/����.��/V@�c���:�!Pߡڜ���M�n�w]��R�3��n.�y�*�=�HѲ 9�&���\ss.70�y���*ؗ���E� Tp����N4���Ac�OU��q���<�&G|��f	�g4�m9Sݽͱ-��ֹ	X�̡II��s2�t�J�-�����+���̠/y��:m
�*IH���ޥ�4��MO�z�T�<1f�/R��rxm�E;r#��Ԫ��e�cy��~�N��L������T	�N[l�eNi\R!Nk���yV��y@����¨�#FE�[0�
���"ζ�$�I��{P���*��=i�쭼⬴�K�Jyo���e%�|���^��'�@�S���-P�;V��S;e�k7GyͰ�^;/#���t�ҽ��i�]�t�jV6���ґ�o:��E�Vc9k�r�P���C)M��n���W�����{��"G�B�
=u���,B:~1��5/�����}ZkĪ��]J��[-��=�Z�:Q�]�ξ�.BO#���[짷���߾���c"o2���m"y���2��^*��ޯ:ZkR{����kxW)cf_5Ӆ��Iz���;S!u���c=V���Ӽ؎F˷#�����pH:}%��;��F�p�b6)��ҳ�^�ʖ5�����Sۊ���3��Lp��z�T0&�����y�⽋4HΗ��u���$�d
�7�9�%�orHɞ�6(���e�̐gYwW�3z�*���l��תr��z0(�U�EJ����_I��!�8����d-P閸Y�u*�q;�V7�J��l𔠃{��b��%��4S�(E�̙�v�z&塃��r���\$���j�'���Y~�oT��3y��۵����*X�e�Mi�˘9J�Ƥ�f�n�1j�ӊ��H��i��n�Њ��^�:���3VtO�VV
���Ub6,����ıӫ�m���Nq��
��:���4��6�62f��8��4s��WU��]��C�b��+���osh����ܔ!6�;R1P
������9��J{�����¼�uɃ+f�1A00mxI�>�t�\M�ܪԴ�v�i2Ͷ�S�����xо�܌6È���̢\E��+[�_[�N�S�H^25+�'��z�{&;P������YnM�J��ڑD�`{�RǦ��Q�1�:c���Q*qfp�o嚌P!f�^U����7�i������E�F�ء)m�ᄭ�b��,б�J��	��yS"�G�B|+-U�!Q�kpg3.n���$a�ZͼĠ�/S�J�|�n��90Z��Q-4T	�sM�
efn3�t�.Y��<���[l�Z��}�'����u�1v��;)�r��(�:-�J1o0���6��VgZ��y𙵋s�2��\͈Tu{��5�������f^R�y����|���Y2����\���P�9�%���3P��ά/�%�����,׫���bT��δ���ݳA&�9�&��r�]����4_,���E�d��u�BWf�BjŸgC�,}�S�SD�D)�5Cou�����8���'���v��5(RP��j��� X��O���@4�%۽;�K毁�͹c79��$;�{˦lؐ���1�L=�O�л�(-�:u�®���y��LW�ڕ��-���"��!-v���H9��	N*����Љ�$�5�c6�G�/�]L��-"9.�7mݰ�3cj+-b�
j�dXwN�8��<F��$��u�71$��wׄ�C�֊ĝ�jpXnKֲ�\\�}�qX�j*���f`�l]�L@�҇�)Xܢ�2���OV� 3ܧ=R� �'�sUpwcX���U[F�	z��e��{x��I��E��q�n��L��s7"OF�3h-�8.D4�U���@��qCt'^��;���d�ᚘ̒kb]S�\�t�PwJ��_'�V�$UhAY��I��y�gk<߲@:�kP���/�M̷D�n��1��rpD�q�*JV���}iB.|�����Ŋ�:��'*R&�4-�>ul�;�u|z���w�'}[g~�z�윆�Y͙�%�K�`�m�p˛���]⻰�Y�������NTװ�gδƈ�	L3+y��^21���֜�$@ݦ7�f0F+����'rͧLi��J�Zy�Q(�u�Y���ٹ�@���6��{����Cfr����!<tZ�F(�*���Xi���q�P[P}F�K$.g�:wU]����䂗,���1TX���F*�*QX�d�Vk
%e��ErՊEAA`X�`��X�k3.�1(��V���+mX�6�6�TAq�-J�X�a��Ĩ,Pr��
ҋ�)m�s([ab*��(�����-eD�KB�*,ELu1\I�B�ED2�v؊.��k*
�UQ��6��"(��Gi�1Ab����X��B�EY�D�3��Ub�F(֋�,R�ZT�aZ�P�+��&��mF� ����˗m�Q��*\��Mk��ZҪZŢp�5Ԩb,QE+3+�U�+V�aQG.&e
�UE%m&0�B�hT�FM-�v��_����~�̺oC+%u�DT��M��"���N)��xk�X�7��kL�������u�.|��c�u8̷@�a�y�56�g'���R�Ԏ���zލ�v�ssx�2�^��HU�޸mG
��0�����NNﰾFsԾ<T�!N]=;�������*��t�KCx�ߪέ�(׋���ݞUDd�c8+m�w{x�w�hGF��^�Vv�:\M���F�4c�ގ���I��î{��N�R���8U{���9J��:rk5.jc���)Е]b���p��!i66�{�d�e��{��0�X"Td�0{�;ko��K{z��E6�͕��ͳ���S(T髙�/��[��f���Y�r��y_����=\B�o�w.����Q�tz��5��w{�ګ�fy�B�Ǿ�Ϣ����L�H��lGvq�=x����n�o�E�7�-�٫bv��6��<yΕi��!�s}|ҍ�-�@��I�Fh���|KLOG?6rr�c*��Ŏr�����ب�MA����iƙ���/��;k�kX�N�����=:��6����K�OekU��o���Gg#�
��P�W@o���4>��f�i���w]��m�8�T����������@�8uh�*�oBJ.%��FV��!=�VK�L1�EE���r�'�T��h����تa�V4KW�<��e#88�7Գ%I1�j��^r)�z�횳sCw҅ DC�-�+���]׹��$�)���feZJ�m:�B�iRJS|˱���	�ڨ���+~/�Y��k&�{N4�M��^�j��/'��G���=΁yQS��̨GVҘ�o8��WQ��WY0�l�^o����N��rr�h͵�,޶����J/\����̈t�-�Ee��u=��	�,{�7(��Nӝ���W��6;��F���x��jU+�V���5�;O`�V�.`�['J��+�:����EM�J�����p�>S��.�׫̓�CY)��T*�Te����׼/��R�a�.��h�ۛ)V�`hH���/6�X��.��|��nX�u��ܞ��V1*h���9�0�:I*��a�"BzC�V�~%���~��:.���27i.fP����)��G!0]	��N���I��w4���m�{8�Īy)���'jfav>����-�ew?=�9jM������<;�����g9YG��~�[=0<��k�|w=1��6#nx�Ѵݻ6����7^\����:��lqKe���2��U�	�Y�M�=5�`G *w}"� o��b[��HV	���4��)ʌO_�}��,�n��,4Ⓜ
���H[���C�R��f����3>�(w��!�8�K��+W�h�.}�V�M^����zDCbٜ�[rV��g�~S#��ފ����[�W����b��D7��Ĺ8s��u�1�Q3�wj�[�ӗ�z��(��GgI�η4F�4l��S���f��+4!��,I�~s�/ĺ����tO
��OjU8��5}��O[@����Uk�����W�z���p*���.�&Q�	�"�A	�=R�؝T.v��'\�݊HUZ�UHq���^����^��t��l�9��_1+�3�t�jam���(-��q���t��$��fQDYrz� r�JC���n������y�a��ܫ�^�i�7�^&��LX]�Md����Z�9v�2�ô0�x��)�4�Rd���%.�Ċ����ޞoؤ�ߊ1H��`�e�n�UB!�����-�##i����͛����A�P�N���2�:%twJBL(�t�o��N��W6���%���{0n�n�lq��#��Ԝ�h�6�|����"�3�\���'w7�0�0�ڕ,�zE�w]حu-�*��2�w��[�u��^�l@An���U�w�j�6���"z�Mb�����7�+�O�l3`J���V��G�	I4��S�tsޫ�J��F  q�~پ�N�,8Gp�B��2+i��},Q5D�$�F�TF�l�S� �ooJZ�y�ʳ������A�y횖6�'�f���඗_+JͶ�ޝ�(�v8N\�ˏr��i�:޼y"]�iV��;�ٱ�����Գ��1)q,�Y�5GXOH�K#WF%��ҹ�u�ñN��1�u��B��y-IC)Ԟ�m�����F�
��!�@�*��ٙOI�\yU�ع&���ڗJ�eP����s�I�E�Z��n�6����j����P���/��f7KcOQ����f��9M썛;�_Ql�$k��+Ӧ���K�|��'�����x;��$�rY�H��$���E<�\^�i����VI�_,E7�Ps���Ex���\�i�g�i���B���]RV�k[�N�R��=���b�hբ�B�� �C9&}\T��Z�^�9����Ј�$���.�Ι�Ӑ}T�UK������*��<\�T���c�ۼNäh��>f}I����9WZC�9YoOX��~���G�֮�`/��ئF��q"�5<�����*�m:�u�
���һ=%p��4�`�n,A@s	Z��	��[:���"fN
b��k;f�;n�*nt9��'*��/ydֲ��(W�Q@67����;{�&�tCl�Ԭh��g0L,�O0^M�uoj�浃E9�VT׬������E�;���E��ڎwWD�(1w��'��%zcY+v���9�o����2�V4�(# �U9�pS���2���>�|.�NTMf2Ü��V�:�n(���MQ��'�1)�\ nA�]s��]��kQ����Vb�� �+0����z�m��J���ғb��"��ޮ�CY%4*�m�ƻ/�/ex�׳<��Jr/���-�o���:b�)�쎓Ց�;�Y}|Yw-~���O�rK@���Z%M��t.�:����oH�p�ή�p�ս�M6 ��=*5	�+tS����TZ�OgyM��:���L����J�����c.�/uCw¦���"�:����"��e�%2̙�]E�@=�R�/�����aP�遃j\�ƭ�%��@��Vsk~�_��Fߊ�e�>����OV�:Zj'Ǻb,�=ݩ�1�Z�ӯ��%s`%!z�$�zd��ӆx�v�iLF�a�w���6�*}�NH���V��1�zx��k��o\�=P�L[N�3ÐX�m<H!	s��Ŋ���`m�`�)q����ۼCf�O�75�'���A�em�9Q�f��&X2L��$������yY��n�d��b{"K��Қs(6 b��q7�j9N���9k������E��s��[ڽjh����h�E��"Y0��6�{:���:��քh`F�&�W�[y���ah�r������g�P�w�`bX�랆��n픉�դ��*L��߉��-�K�&�#��Ac'{��Z����d����p�������S;V�Q��_k?z5��N�VѲ�=��>Wȭb�qe��mU�U� Yt�l�'�����P�.��:���S��!O�J����B�i>�%��;v���-�5(]]�-t�LM��L�S�KYg����9��w�Z)���m�E��(� f�	!��1z��m���.��Z�Ïk]͜���3��u}0���U˒b���§U�M&��L�<A��T���6"�է`ޚS|y�<ėBdi�MߩkX-ɷ��ͅ�!>�K:����*`�c����=�F5{��^�jVl��5[��
����
@���������hڬ��	���[����f]M'���TI��Xo�?
��"��+%-Ҿ�n6��������yxcmP��֘�����;�.��syӮW{ܒ�ˮ�n��5�]v(�;1tp@���@�y�bxF�0��7����x�G]��׼��ք'� �:�q��sC�}��h��f\�ى���b:1��j�t�E�Tw%�F"yQ��;H�.�SǛ�:oX�ʾN��C)ѥMf�7݃�_������]�u��2��Epۖ�54���V�ғr���4����J�YUoj�f���גb���a*�m�}Y\�B`�Q��ԛ���Iᴯ�c\�6����d��6�s�衏�k�2�N��>�bZX���P�w�	�,�I-p�W%5�(���"Mf��b�)�����p^kOjG���ʘ���8����;iHuP����BIT� @EJ�_ S��h�,>��/���{���Y_�r�����Za��e�@�V�D2��.PDD�$�Aؑ\�mds֊�,Zi@����DT�^Q$�3��o�Nw�}~��=!\�h*U�^�,J�P�h�r�3�(�k�Tƚɀސe�]�ܯ�l�A>����i��c��`�PS�tE?!�D���5��������jC��\5N?��\8��9x�����@�ơ��@��ƹy
���B�0U�ף`�Y���1X��P�;���������Sm���w��2� "���H�δ�cʮ9X0*zi`�&�-$��q�R��L��y�s �.�v�cS�T��q�I�����v�@�O�H�5v� o�M�������������z+<B�������:U��&�}K�|�u���7^Q�h����;�֟�Oxv`z�ߵy�����#y�*t'\`L�\�@�z�{<��I�Hz0��h*�P�a�T��_p��/��P(�*�<�m�{C2�A����PS��B3`jH�c�d "*F-�2 ��\fhh���)
0�P�Z�1C��JQ=�/l���\DT�T;���v u'R�1ܧ����?#�ڟf�;@��	��NQ�[Q�~�5�v!�^מ��<�=F����i�{�3  "��n��<�y�)�*r_;�dT�>K�4���1ڻ��P��o`��J��=�*��Q��N�p;;��������eCz��m�8�%[rM�=)+���r&p�Hn�7���!e/����. �z��&�E?�쯘=;���tur܊*r^X�0�˕{�Ẽ|�G����! ����PM�i�`���H�
X�� 