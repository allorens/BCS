BZh91AY&SY�60-��_�py����߰����  a9�|'�
)J�©l�@ -�mR�e�ْ �v�R�m���`   � � 4P   ����   ��@���� �D�� �       >�    ���  �R���vw`���:��-��ۣ׽�-�a�  y�<;��U;j�����m���ړ�k�����V�����.��C@�7jV�ݍ�Ƞ . �w��  �ވhtӭ.T�l�ZV�B룉.�Cm�$β��7-4k[bN�� �=���l1Jh�*y�wM2�[l��ݲ���tA���u��)�wm��  ��  8=�6����ӥ:��5݊:�GM4P̆�r�G�P��:�M�`�:�E ��s���Q�M�V 9� ��zh4��mN�rh�l�SR��rt��< U�1�t�1��S�CB�A��4P�6h4tx �  �0�  �M:�v���Bh3���h ��t��]x ��@P'��4V�)�t��\�1���B�Jj�                  �  ���Sɡ��R�H�L�h� � 1#O�EF�F&�C �F4��@&)�&A�2djl�O)��2mM6�5?"�	U(�0 &� LRMU&�ji��Ѥ � � $Dd�T�h�2i��  �2d��O�ј�)Ր�a�VZ�F�֢�U�7f��f�&�1�g���bb|�E�����������!T�@Q�@��G�Q�E@�T%D��_^p���,��EA��>�c@��@T �����E`fV'�~����\D���>��@���X"��O������o��������3�i��Q�N��$��a�z1��+��HRO'ę��*�
��¸P�B�h�p�� ���W
�X-B�p@��;�0�/����F�a9S��<�1�j��o��&:>Q��XVg#)u1�XA�$�p���ᇦ[�|�Wu�
Y��0��hw�q<.�*��7�XT ���\���C���h\8pt������9��ݼ�ݧ�,��]~�涒����9�o��zZ���i\>�^S�<d���x㤙/+x_L3t3����qD����&\,34�t���zI�����^u���I/s[ݩ^�]Ks�%��m#�ߗV���=�]޵���&f��5wn[֒�Z��R{��g�YM�-���b�2_�3��b�q�r�`s)�.Ot�������]=���ַ�Փ�]���[��]۶֤�u���kk���gv��zKn��%���u���~kr��-�ַ�q涖��]�\ktqلe��
/�x����kas�0}~�M�O�x��+F�)�ԗn��oO�(`�pQ,X�!!��ٱ���K�
�K/��%��BI�K�4��tO��q#V6tl�L!�H�*��^^�F���G��Çm���;��>�gN�?<1YM��paEga�z%cU����O��;I83q#��,�hТxr6(��������9��o3�,��xb�xً����H��v�;<se��+t����uG��Y�3fd���D�I�ຒyI>��i]ƫ��Ԯ�$������J��Jv��ic����$)$�$��}e(;�K;���i������{M�n&ɮEu��+��VqRL�I�'Y\3�[����62�+��IhPL�du4W�ݥpO�oJA�$!\���I
<,����3�$�Ё�!0]mk���,HZ׿���r��%��,o�8Nh���]�ފ�o�<z(we$t"Hx<���`�Y�NX��D���Q�+�B:.f�I�+�8{Ty{�VQ#����I�)vX����>���b�W �bD�Sd�BG	���[~��_�~U��KSf������X9�.&��o��*���Y��|O��R:�$i�hxō���o6�y�2�d���
�������'�\%�-�<6���4;�,:�O�n���KIbՙZ��Z���a�0��c~$�p���ф,�����äx�f)�c��0����̓�,�Z��n�ޭ^5�<��~K�N`�z� j̡�|oĎ	'85��2[�//'v�J���r���-nR<0åau��2�*��#/�<$�c����N���ǆhxa�Iqd�{r\�i-���yn��ܼ��E���v�{����լ��}[��Z]Nj��]�)w�Yym�_��).mi/<ZKX����Z��ՎZ��2�ݻ���I.���t��%�R]̼�?t���i{=���嗙y.X��?--��k��-wu9�_�Z^KI,�˻s���"�����ќJs������a�X�Õ��0�e��c�dcQ��1x�⇝Nχ]0���/!� ��-�a�0�`��3<�Y̶��Yc�VY����Kf"N�����a��xw�
0�(�t�F[�������ْ죖a��V>����w���K'zK�/8޿wy޼�ޕ�o82pP4a<���N��C��8�ʈxU���1Y�����B�C�B�#It<�y�GVU�x�.
���H��"�g��!-��^����ɾ�������-�]����i�c#���g�1����C�z25���o����eQ�r[���૑B�З�����3�D2�2�W���&�C]�u�+'��Ȏ��0u�<,,<�9��K+�p$�@�i< �rb2}+1�pC�ɾo]���O�r�z��'}oI3�Ñ�����ď�֌u;���]۷?$�-k�S�[�inִ���u&���]krw��'�..3+!�f[Xap7��to3�xb��o�3��|����d�c~;nZ�[��뻫��.�ZK'��R����<8k����	��W#�E�|���H��#C�]�Æ��"ňۜ���S�%�޼��ZYy{sM���p������ß#��8��&��ÜG�O�r>C�bG��̱h�pAU��Ñ��h��l:<���8���O� M"tS,8J0Tp����}��E�k!���H�S��<[})94xv,n��G���G�g�	�S4���m�/u���7�.��䢜�0�� �c'��W	0�C�1�L��T�@���P`d5���c��^CA'�Q�&�1GFh���:4Y:,s<
=��:���v��;�#
;��GB�:��0p��k�3�E&�Z�!�CYƳ�evv�v�<>v|��(��<y${<;�5ԍm�T	���G�D���^#T;u�Fƃc���H��{-�FQ��}���HZNZ*z�>�=mȋ�f�����������Q�wy�.�G��x�8�6��*�/B�7�F�|���
P�A�lЇ���C�}�X�=����u����'�YVs�f���p��at�dؐ������8$6M�1!�",u��Ո��ej�b8i)�yg���#���N$p<&�g\G���P�^;Na�W#h��P�xZ5f��xS88�vZ+	��&���	vz�=���G���tc6yG.G�ޙ��C�R}��	�	��AS�uO��Z=���=��#�Y�`�_u�xqKŐZ,�)���K�$�SæL�Y3ZZ�~�ɽ$��o�~K�:��y��W�R(A��+�U�o�KOu���k�w��K3^]I����2\a8e� �MR�q�gV'��q�L&�1d8�	�q�e5Ä�+��鈰���VÅ��Ob~:dۅ&,�I8�v��{!Z����"�p}
vxp�������;+��¸pxʡ�u�Ä�+���B�8�	�q�串Ob~;NL��{�>)���hX|I��H�]�p���!��ڒ�҅ӚxnK:B���S�ta��,���d����L��G��J�<��Wq��P�:6tl�����mf5���Øp����x$8nqT�;t�a����X�V�ļ�,Y���\�ח�5���kvY���%C��o=a�m�Xي��#��D��lQ<;N���I_$�����b~2�#��/����6;My�����b=�R�6��2�H�8�8�:�)�O�%���bAZA2�.��RO�'�V�5\�֥wI*�.�.�.���k�*�I������%i%�%ԓ�+��bWܔ�u�-&����;G0���Xh�F���=f����󡂅�Gq�%��k�|�
��NOC��g~ Z��r��<�#�k�[.'�߾����:1H��8���_	/�*����1��E�U��$�~�#�R$�=?g����ז�޽�"�[��Y�Om��z�QEc+>ya���xЈ�TI��ui�1ǖ7��5��y�㥯&��J�,R�����Wz���
�h-¨�U�dv|�4x�W�i�i ��͟{��0�vk	����&+(��n����'I h6p�G;�֦��C���	hE�z�L��j�*�]H�:VL{H�dK����a+׵��YN���Mk*�/[��<kl���Nǣ:K�"(��(�_VҶ2\4]
k�f4@�Ve��خ��B\�fꤴ�n�}n��}�4s��)�H4��dJ˔�G3k�6G���oe��U�L?rq�8[�+��_}�VH����tUGU�n#�-Sy��ن�^�,�I>�Od�}ec�Kо>cj��ˣ��Ƌ ��*�"�]��B�UP\$����%[�D�$�b�j��E�ī�rm��%%�>���TW��}We�͕�攽�f����O��a*9_85#b��<a��z�`*\d��M�^�8�Ϛ-c������m��h��ʹp��xq�jot��zˍ���|���p��i�#� &�b�ƅ�J�k�D�oT�x�ٸ�;s�N��c�ޔrYJN 0l��j�)�	m��O^,�f��GP�\N�F��k�ݲx�G�v$�dVt��w6��a�l#x��z�=SA����d�ᖖ���<OS��vnM�X��^ǥ8z������C�	<x��:��x�a��8�͖��Q�d�xj4t���X�"}�և���|9:{�)%�,��*a0�J$���ڑ�M�"����wn��ѣ��x�%�0�~h�g�x��#f�-�Ζ|s&�,�P,6m�"�d�I�n���:p�Q�sY,��d�35�I;�b�G�I⍖Q$�(����ӧ��0�I4��O;$��5v}�Ϩ�'t�d�n|x�0�e�}��O��Dgc�n��4F�x�ۣ�7 D"\`�����p��}(�#�����uaxQ[b@O�je.�ɿ���qE t6*"\F�|/m�;���E���C��=9�>O]( �E|���>E[jZ�9�O4l�����T��B�*,����H|����>�f�U�#��@��!�
�O�9~@�N�])�5��a��C�ӡ�ҵq�-�e��>h�+���1f������� fD�exq�+�6a�^��!bg�#&�|.6�0�:J�����}��� ���:{����'��:@����xaoh������l�}ݜ)p��&�e;z�Cs�����7�g�dd�dL�������̞Æ&���.��D������0�}��������&F��?PҚ��kX@H,H����8@�r[���:h��w����ڑ����%�a��YL��� P�φ�v�Z����OO��$�H�+��_��X/ 	��|8�vP�F���dl�r�޶%e8}FΛ>f�q��H�zT %�I���l
<��EH&}��:l�b�N�H�0����%����$~�'_NJcћh���)��ٱ04����d�G�QW��r��?�+�>�廘�)�|�*f�:Ufɑ��;r���l�X� �����'[.�D�� I�u�0�f|�٧�}Ϳ�:lç�<,��F����ia� Y���:t�����6R�k�F�?,j$��fΟC���|v$z��T�����[E8U���+0�E�z��R6YF���>{z��z�ъ$؊Η|ɢπFX�:��S��x�F����Mc2C�
��ᆍ$H��:qQp��뷄��TG3�$�F�c�� �W5���M_6x��s\0��pDt��+�P��,�=�m/y�h���[�8���<
��Uf�0����	���Zeޙb**����TY��X�����l���1f[�ORGG�@��F�?�����??��TY����e�x�tx��sD�K8�n�ځUC��:~�����(�MmeQ�����.zK<���}#:��_
�m@� ŬUI5�����j7*gz�o\ya9��#`����GG⩹�ۏ��uz�+YW#���? L<~*Ř�NX��<��f�eƃVM�s� �vma&͞�x^nԻ�����ٳ
�3%;n͚<o�����j�՜?ovZ�ڳҏ�t��K5�2~>ϐx�Ͷ{[�M,�%,鲉��䎚> ���=�,�;�vYRU�2х�����yΏ|��≳���y��w��D@����.�����/3|O�4UWe2N�*Ҫ��,��8p̎���h�$��>"�k��6�z����<���@����-�xt
t��xDz�����$�ٮ�(�W��<p�k��*F�<dŲ����>�lxh�v�ٹ�Q�u.��	�Y��'N�J�p��{�����g�p����[@���Jo?_'�$��N���R������1@�=)��(*�_7W��R(�ç�e�M� J:��4��]L�:]o)	�zQD�>Ιex6h���GN�-�F�Zن�n��Y\S:a�Ft��?��p��j��;�̯�7��5�&]���z{	I������M�'�#>�J4�k_�'��|`��=���E�%t٣���s�I�M�~9]yDѳf�<Q��IE#o&sⳫkU3��2t��:�f��'U�8l��(���p��5�%ֲQW�2�N0��`�Gv�V�1�>�&����Q��4~����� �U��@
��&ݸ���uV�6����w�f�>�4j�|z2�^�ei㤒l����Ň$��0��M�g�'UŽ~K��>��6���I�Y��5���,���|;�6a%цA�-�񕂳���|?�P���4~<�����?aK5�cG��d�*ɵ�s+^ے�de;���@��iSNy��V�iN!d*�=\�N2�M���r.��H�+�IF���l��a����u})�CWO�6� M��� ��cp�zri���l�Y�Gaڄ���>y�ԝ�yo�v�ϊ�l�+�� P�z�9�[˫:��iD
w��0�O�^�U���/9����tQy�����{m��(�GgL?�'!.�K�<h�͝�*04PH��=�4(���t��}�ӆs~�]vl���ƫZ$��B�ӌ�G�����I5Z�F��_o}�=��掚v�ƍ�I�Qa�I� �V�æ�S�M�������ǎ�� ��[�%��->t���h�E�5��:k1�Hu�Ժ�	#j�ս$Ç��ק�@�ꄶ�,vh��H�E<MkS� 8��<Ns��\����>\�6}���R���E�:���65R�T7uEXk`�ǎ2�S��]N�Q&�"��u���6|OТ���.���cJS�l���>�O����eq3"�l���qh�j3�rỸ<b	���� ��~�����Y��탚�;K˭ NKØ�Yc^f�e�ԁ��{�c��M�����/��*@ŵ���5��9NLrs9�:q$��L�v�Yd�F�<"&+���Y�c8��rD�눓�9��Mt�&2�2
�jق�^B��\��S���s�����ޝ��wQ�!�[�h%���ŏ9�޿O	��츖�r1�[=��z��आRqályoh]*�f�:1�A�<������bs�^�	�'n��F͵�����=םc���fbK]@�@�$J%�-m���	&���Z@���jBk"�x�ْ�����)F�!�<Yl��3Ɍ�DyNܡ<g�"KK^+�ח��;�����)_��OD��j�g��v�iebsy�rﶛ���B$~��aϗ�b��I�e�d����$	G�w%f��s�������ݞ�Yw,�<lf(�8^v寺!�t�Ц'����:��g-y�u*�:�k�Q��E�(���T���iñІ�[����LC��;zt��	�go;��kgt��p;�����	K�t�M!�hn�n7��)l���7I�LN��^Ya7+-�%"IAq͙�d�^�ײ��־��4{~����FM4�Ilo�l��n]���6ٚj{��V���W�.�B�y��^E��͠e��n�t�{{4���JG6�mkI��,3����s�&Ӳ�%�\͵��q�A7�A>��q�Hʎ5؄c@�|��!�),�bZG��뭅���_!z�.s�9'&.)��β���."��	pz� �9�M����@�z>��Ul<=�TK\�yY�fB�jQ�gZﭨ뫝mP�7��;.�b%��)y���9��G�d;���Rj�Z�+�{�ii{$�5�Z���2A�r�E9iCR��:Ю��"��*��r�!ԁC���=� �7�L�4氥�N�mbn
L��d�N�`L�R?��!�$�unCV@j/.�:��rF�Cۯ3v���������� ��~����.��*����Rc�);�������qL�|�c�l��+����ڿ�����^dffff^f����@<@xh ����=6bpl�� zlÀ�;��P�:٦��C�<�4~���P��2�3���(4�+M���",�#I@	��4�,����j�_��_�j�۝��@�   � � ƀ�a۰�t��0�  1���<4���c@� ��A��� 1�;��C�;�p�t���������E!Bu�@P�`K@��
��*d��5"�(K(P)B%"R�J�J�@d�2+u~�����w���C�<��:��� zlÂt��;�4 hÁ�@xhh����v6� Ɔ����=6�M��p��~����w�~��Z�CJI.C@��C@�-*�ԃJ�AB�1̯� "p��1h&*w���~��݇ �8�< �ta�p�@xh��x:��Ð8à<@���Á���l���@�;4�o{ 4� Ffff{fffut`6�Z�1��[YD���:�2iB5��+��խ�T� �N�%T�@��FAB&B�H�J@(d&�u)�
��5!�Jd	�*%	K��1\����ih�?��?��y@T ��!#��=];z 3 �b�A��������wR�����K�W򬖤�^I,Z�Ԥ��r^�Y%���]ܷ)Kv�)JRZ��\����互�K��{,�^�,���d��Y%Ԓ���wjInK�I,�w��-Kwr�Iw$�KW�]˫r价u.Z���d�]�$k^Z���ܒ�Yy%ԗ��\��w%��rܷ-ڟ���/-JRZ�wZ��V他�.佽��ww%�]ڔ�ܒ�K�,�InYyn��JR��)-W��ߓ����Ol��~��j��ZK<6%v�4�����2�2���u�tu�GFP�]q���R�th:�)*�YV���[.eڥ����ъm��B$�0g�hM�̹Mn�fJ� ۜ�M�LZ�r6XYe�Uvj+�sW7O�ݘ銟�g^�e6�S6�i*kt-�l����K���.'�X!��L.��Y��m-�0-,g2��<w-�Ƶ�����r4�{%B��؄���L��Rl�K��X��s����Ia���G8��-[e&҆�]�t(���6��:Z1v�xC@�`���a]�ͩVkHJ���:ykc�Yv�Mv!5tkE#���*������Wq��hlMv)��nm4�s��-n�l#
�����S,-�+6���Ѫ(A1L�v�:�n!�lk0UD��2RhAu�KU���)�/;u�
�Ԏ��5��+[���ek6��wa
�[�%Ʀ��Vi�J���]�M`�ˀ8BY��v��HH�Wp�&ŰԎ��l���16WnP���#V۬���6���WlBQ�	b]^m�Wkt�h��ib-�5�3�fҐ��Vw�t��t�!��eֹ.�k����m���jĪ�%rXSc\o;�w���h��*�5�4t�Ur�S+��Z�uټA Y�*��eL3r�ixjMm4ʫ��iK0GÂn]�-)i���ɥaŴ�:�^m�
Vd��!���r��q��&r:6�M��HĶ���w,%�N��i�ť#�^Q�j̸�Բ�;SaH[D���`�_��)���ǭBa0j���l�6v� �:�t����5�F�t�.s`M��6���;^Mi-��C�ł������鵶���p��@��ݹI-�.�Y�v��E�k�-+�6��m��A:XB3C�k�v���BR���մtЕrK2[ek��3ZA]���,&h��]CC�0���e�]����VR�K.���튵�~��W����`��O��9`����:vS�K���փ`ki�Ơ�d�y�֒�vf���b+)��in����ww���]tԵ�+e%r��E�y��ba�X��-��i���	u��m�W�}��HĲ��%����T�kh�)��X�Z�ˬ����.�SZn]�7�D���,�zس;��t��[e~nA�� �j��(I0	M�6�����Z����!�f0]�����m�ܨ͆�B	���T�A��Vl\څ]�j��\94Ksnܤ�5�cf�.m�V<N9ۛBZgi�\�bm��ء6�n�5��|G��M��]K
3[�KB�[������i�$m�qXv^���cU��ҩ���1������\���6��w�����Y^���ښ��s[���Y���B�YR��h3k]��"��Tlť�3b��q�Rˁ��m0ؠ�:�۠k����Y�6��\PĹ���S&i���"K�@�Zj�Rm���@��WX�.M��]�z;M�l%��t�.��]ǀ�Ԛ�#����e��2�]s�n�á��`��F��F�j(�i��on�m�+����%�r9�;&�hhִ6���	������+K+uЉ�4V�0����6�Kc�~M�M^�&��3-� �K��`%R�[*�w&�8��F�a��1���Rh]sK��b�XS2^P.'�۹�"�9�s^���:����an1�-JlKVZ���ņ��KRWU.��rl�mf	�%����]4Ѷv�l�X���s6m��.��:�W���d���AŷQn�ki����	��2kv�Y�e�� �FR��.�X�Msn�:cc�1�x`�ֱ�u���B�b�6�B�h�7j�R���3ﱠM���8���~���s��~�~�W�� zl�9��_�~��> 4s���_�U����|h�4�I4ᦘQ�x�If�a����2�'��$3�P8σ,vb�,�)��S����D�ؑ9����6q-�q��Wr�ˇK0:��mtHnj&5�2�+ �3�����w��b��+E�N¤��]L�:�d%o5лe��ں����#�tu]-R[�K��Z%a@��mI��$�[�v��5L!F�BXD�q��.˭	k5��6Ќ1��Ŗg�NK�,q�������!��"d�9��^]Mn6�h��b���RMϳ�Ӯ��ZVY|Ժ>K�Z3$����Yg�%]��2�KS����n����p�
洱�ʅ��+nm�aGl[�gngk�Ͳ��kv���A�!um����p]�R�e��/h)af���w���t�Hdۛ&6h\�f��ԭ���,�� �q�M��C���*Z�5�b��3��h-�K��z��h�r��/6]A�d�H��j��MK�uiеT�ݘ�tMVXy��5wfͽ���X���y�
�pBօ:հ^x�9��T�)8�����ox�0��a�F�D0j{g0gQ)����,����(#�9UR@�>�W�|���Z����R��K���t��8I�h�x3�t��7��_�v�>�)/���.7L+�Ju9�$��b�v�P_�8��s1�ݨ8�Gߑ�'Ft��I0����F`����F�0XcQ�
@����UG��f=��xj'�I��7E��]F�"L�Q��<t�I�ǦDyjgSFk(��Q�M�J��*�7�#Y��C�_��LF�c����Ŕ�ѫr����$`Ρ����E�g"!��<IP��WQG�)R�A��,8b3(:td�Id�p��
0�p�8h�FvF�Vա�� "M NS�C<@�^�� ��UaD�uR�|�2S�	x06���T���dF�,Xp�QD)D�����'��ƚ0���L\M��וQ����uZ-���i��)�/��r���ʨ}M��J�V5h�l�2"�x��]�L��qB�qP�t|�������svҌ#e�pۍ]��s��D[uчJ8�ݸ�"�td�2�Y%<xҌ0��<a4��Z��(���wI$�-"<�ui�s��g�
����<`����xs���3��RƬ��t���DI
H�����\6�GL9��.�_G�a�(�
U##���̧f8�5���#�K�QN2~ÿ,�'np�a�]�oG�;h�1OKpT=�7ўc-@I<p��(ᦚQ�xÇ�`�A,0�PH6�0ڽY���ů9(H�Z�
9����GW�M�����ysz�p���݅	$�=4��u��|0�Fmf�G1�07�-陳��g��k�NC�5ښ���׋]쒥���Uƞ��֭��|{oxo��5;ռ���#jɱ��ú,�47��������hx��y�S.3���q��l�%�QV���!PP�(�]1P�uwz)m�\)A{��d�B�T��z[�6��Y�S��D/,��(��)Q��4;E�+�ɶy�$����������%�J��F�L�j8wh��[nc��xw�x�P^�>��#����n��S�7�p�Oe�$��Y,���e�Z�������}R��l��U�D�I�s��V��ț*GӅ""n�"��˓��"
G�R�E(e�gF3G
 ��TQ�!���8R<�j��:�"��,�Dcf4ڌ5��R)V�ѳ-���×A۸��;��0��%3�1����!�E
IVa�XIȣk�ݜ����`�W�`X@�81��d��K%��Yj����V��B1�ћ� �b�`���O9:���K�zp�$K�����6��a����_�X�/f�N9�`w���3�N���"{�RDY� ����5��$�V.Ŧ�7T�Qʥ�x�C<qY!��YH�v�L��&�w�)q���C4�%�c~p�u,6M\:B�G��MwJ��L�9ѣ����m6�6�g�X���Tf�[��/n��nI}y$�Y/+ۆ�`��W���0�M	
�$=-��]�p�!1��f�"��g\T�?>�R�K�b���Ċ�����QIx�TQҟ��:tq�q��3�'�0��%v�����]#)b2����%C)��5��8q�m;;'7U뷆\֩� 5p�5S��" �J��A�_^�K�˗�K�%��y^�,�0Xae�ĥ���>���N�a��g�, �1g�7�o��e�	��;�0�ԬmJ�H���'uPPQ$�F�/Wu�4R�ʽle6���ι�+�0V+/���1�(���:{��/^�ð��gb%��yWZ��n�� ��u�ɭz��gK�>���qn;,=�YJ+):]-p��6���)a��c��c�}��J^h�h�N%��\{�xkkl��<�m��Ӧcm�N�#��n(,�5�N(\]L`ym�n`Lx1�x;�@~��,1�Ҙ���e�q�N�Ƨ���� �Ue�L�(jR�p�t������z���\����Id�^W��-^�V}�����Й���NC�� O#�J%,��J��<���#.���{x�G�"74��n&bU��`R=
����J��Q�=*��ۂS�T�EӃ��N��m�R��U�!iC|A�
���HEB��-��z������MYK{]#r1qB"$��G0�0��ň���f��T��p�FH�����<����gM��2��zF�F�G�ò4z=EHf���H�a�=���z<���J���f�C:9oHg��h�l6�p��h�=m3Fh�ǃ��d�!pz3Ftz3��h�kp�v=��HX=�(�0��8Za��i`��4p=G��٧I���zIi�F�G�����ɑ�֐�Rt��4z��њa=m�i����=��>����d���ĆK�4zY=6�@��H�H��idi�zF���g�"����� ��� |4�G#�a��O[��F6�F��ѱ�4���!�kF�}�@iD2�F�%h�?�P�tz<4�"�� ��$i��4����x=�i�
4�a�"�Q~�>>2>ʈ��~��������#Dab�K�Y��܇�t�If��a'v��7x�GK��m^7�����;��Q]>�^N�Q(P�����dPǛ�v=����sGJ�㇈�G�����=����|VA���E��^���/5�{B���wA�vP�[	�րBT��\몸�׻��\F�ѬI�Y݇�&d+24LݕB�r�i�h��J�@&�˱�r���"%| ����!��.?���y�~���/^���� 1����>�Z�~�Y������@h:뮾�U���fff}� 4u�O�~���f��������u�O�_��Ye�,����iFi�a���<x�Y<�B=b�X��$��8w������x���F�izS�@�/�'�c��,����bf`�1W-N�=3��&���Gq�!�bۍ�]$�e�= � v��i�����@�,z���1s���36�R�ѩ���L�ÃL�ن�}U����L��c�C�(,h�-$���	Dz�pt�s��}ۇd�e���c>CO�f��ˉ��l"p�_�����m��=�!)�&�/�:�8H�:Id�p��J<x�ƞ0��2�AÉ��r����b�X��$����c�g��1��h���٣Gɚ4�8i�~����11�sɪ�Ώ�ǆ�8Gd�"�����<���1�L���;�%L���RgJ!X!���ђ6�K�CfB�������
#It�A�ER�d/y4�0��=��IqI��l�W�rh6���
�a#��d&������_���Ҝ ĆO��q�F��vt�vJ�c�S�!��m8)t�y�1p:peId��%���d����������{OƆ�Tk�*W*��xE�%��I��
؎�]����ɦf<{|ʖx�{�P`�T���gm�5�l<L�z+�A$@ @��Ys�m%RF����p�ȿ-��'7�l기l$�ysA��H�,�^�5���7���eP�[(�(�|<��e��L�<�]P�@c$��:3xb�E���!�H}��F�q�1�i��Y?�~�< ���]$&�����м>��A��Ӈ�$I���;!�J� �Ϭ3I�D����TF��m�����w�$�H��WPtciJ� �:��=ݎ�Ꮇ&"d��=g	K�����Gi�(��i.��0��(z:�,���|�u�a�O�v&�L��ò(�@�(,a"�[<#��[M���$b3��`z����0�A�C���~�aϼ�3�0�hѝ�ğa�%�^I,�K��R�KV]^ں�Ӷ�6�l�DP�V+�Ȑq��=d;4`{�����8JY��
M��K����!?eEc�c����G��h퇇P^&�D��f��ٽɷ]���N/ivXy�:ұC����p�c	���Tf��r��,C�/�'�1&�^�v����#g�;��$Т>�TY�*7c��4�Qq�>^��jii�i�I����z�����0{.�LS����!#�h����!���]�1>#��_\0|�DCjD�C��@��j�@�I��>$�N�a�0�
,f4�X���6��m���&�~1X�VF�ߙR".�X0��H�|A�8
�u|Yi_H5�`�ǒ� �_a���LC����MXbĆ�JJh�A�3�7�}fVY�f�s�Ao9��u��$=x�羏8� �>`�%ϫviS�@���	bP��H����I�\i�W:vmh�j�)3�@��1&�чm�+�|vKa��Py0�!�|a�G��	�'��S;)3�H����I�F-p�y?S�xA����l4B�wp��	�9��u��3y�>i	<��q��܇�a���A�' �%vqB$aѢK�^Uď�g���$�M?O��Fa�0��a�O��%��6�`��4��[����}a��f�J�>$z�ă�7V}C��M��Pq�F�.��=H4�7�bdqه��޺�  D|N���E�lH|�)
��?�of���{٫8����b���,��&z�l��	9��2i��B=C�4WJG�V4�������LK��y��F���(��a�..���5c#Ĝ8y ��3��z�q�j���G���$���p����yzkq(9��CFCH�Q�R-Wm������!3"#�IC����9�
�̋��L���~�Xzl�&�H,J�C����ѣl�Cc���B9���C:i'�4����0��aE��ƘA�����d��j�y�H��<��xy�wE Ym�C"�����")�]d�U(K
P�ϓ�y��VfR�[������+7�k���+���N�����;�xϘ1�0�{Un
XIclܡ@ބ��y��T�����ă*�y��z��T�dab̘��Jו{������iۗ�!G��k"�{.+E�ߡ�mL̵�Όb_��:5#5�T�EB�����	m[���h`Q�@��TvQD"d�<#I6'�dr8D����(B���m<=GR�٦ə�=��ᒖ�`!�#��{��Rپ!��q����/sJ�y;Mq��3��̔��1J8����u�mJ(���"��U��͒M�l���E��%;���d���h	��?�O	6�Oࣨ�����52!|�JXtae�G���>dC�G*���r˅I3O�F�7�޺�v��Y�X������bxC��4�:p��?�t���x�Ɲ>>(�<a�X�<i�,��5ЋR�#�eUQ��5��$�H�����5���d#��L��Y��L$aL$+���F��0�`�	);&�n{i�N�i�k�������q��4�x����8�s�}:t�cn��QӪQ��\�Z�%	0�%p�0��Q*	D�1�3�Bw^�&!�L�J�mOŴ��C�8�
O�H<9o��G�-C�z����?�0��l 8���R(�G�2��qJ���0(�	�P��c��W=È����$}]h��:>,^D#���3M$�Ot���0�Qc0��H<Y'Vs���޵ٖ��i�mN>3�x�ﻷ�'k��da!�C���s!A2mr l�i�Bґ����d�ܣ�0�v�,�$��x�q)g�h��T�p�0�øR��Q�W��}Љ�,���Z��kF0�4��G��j���r~���Nx @�0�אL�3M�ugol�����1��&��:]�y�����Z6����嘊��`�<5�?Ϗ��oi:<#�F�C�W|!��}gSJ����JT7чȷP޸꾡��
TB-s�8�{ 0��ц���۶N�R�N���O�>4���Fa�,`���4`~:֦�$�IzO%1q,NϞ�X�VFG�����rI�J���:�U!�'�L>d�qۣ	rd�06A�ޚ�Z8���+��ߒ�Ra"����!]�qjӜG��go	�z� �F��+�@j� �83t��(�$��#Fή@th^8x��f.�8�E����I����s�������e�%�=��BI�p����5�0��Ak�E���>P�F4R��L~�x��=�����5�ë�uZd��0c�qW��P��va��o�F��b�x����혚|HքLl�̠谟H�`�M"�Q�|AF��5���5�0zL=#M��i�4z<��h٤h��e�:4���<�L>'������<'�����#毊���4��ьkFh�F�|4��!p����g Ѫ�����e�Fh��H4�0�L!h�=0�G��H҉'G��t~,�C�G��N�J#Fh�z<�DG�����| ��Í�idh�����(���C��z3�Hє3�Ӑ��٤h�ܚLF�Gf�/H��� z[�4ri=(�z����f����hz:�G����H�r=&8=8B�n:8���&=0��c4~n:�$pA63F�|��4eF�i�M7��dQ�4z<4�#F�#G��-��ti=2���zam�(�(gG#ѲH�g~j��~(��?�/���N�	����E��6�i�Tq�v714bU�X;�eJgN�#?!�Bt(lku�/U�fF�Tl�!*}���i��ºF�L��W�eU�Vc2�e�̻��1���4SoZݳ[U��)D�О;���v�?|{W]�ʳ^$�j�b�-:�l4�Vں�J*��4*�J�T�u��nw-E6� |���Hg����#�U��!s�yI�L�^�E���@5��l�9���*4nkʠ��U�tDr����C=)�=33��0����Ym�~�6��6�
�P��Y/�6Ӽ"R�tl���	�4j�Y�L���+.��޽��̧0h6L��֬�A(R}u�c�M�V�D��Xp`ꌭ��������%�#"i�_-/{p]uo.lM=sn�{��kyr`W�掬ˍ6.�c1�G�ݻ,�.WsJ��tz��!�w1�uK�+fC].��lN��c��<囬�,#M ��_�����P!����R���v�PWOL�w:����A�u^��f�٦��u�]>���ffg�g�k��቙�39�{ޏ{����u����{�ə���������{�����ffL��^�]Yue�w�גK$���ݖ_Hh�}a�@X���yD��b�$7��}�<�N�s���Vf������t�ɬt�v��2�S�l��ہ��K������B�痚k����a�������pLY����5q���#&(�B�[k(5&�6��gG��͛�hl����;�fC�1V'+f�[�י�:�^WmR�n�����EUo/m�f�>u�wh�`Ԙ����]W��>�vmz̺�W:c�/림���ސ;.��BfYO7y����ɽ�yz�He���]f��]��	�t�L�ѥ��c�l��Jj�����f� ��y��m+��4��X�ᡵ�4�&�]&��5���Wn-i3�*�'��c۱. �b�.׃����u�.��]F�]�G�� ���n|�W�)f����v�5M�3'>��	�j!Lv�aF�6Y����*���f�����ve#��*"e�M$G��b�8ә�do~���#P�X���?���m�N�u�'�Ԗ��� �uco�,W�(ŝ�����:0`���:g6����_�=X��Ў>�*8�7?�O��$�^my4PF��fY�<AH�v=ɴv^�+�ZX��!��%cL=�B('�H8�s��ta�+� �y�4�8>���x�J�	&<�r��*�F��}����J��+�u�tfq�bJ2��w�3~X�)GKC�u5~�&��j���F0���Pq`�|���QcP��씘xіi%�i���J0�a�a��ő�Ǟ�nG9��,��DDD��'?O��߽��Ge�h��F�k��a��Xۄ�߾"�=P�b.�9H��P��|zK���q�x����@C>?x��u(i�A�A�!@!�Q$�DR!D�80-ː5|Z��LK��Ӝ���Cf�u��l6IH�"F�,a�ݑ�Ȃ&g�t;S�jʎ-�6�+��@����D�B�vHp`P�#O���jV���(lp�+GJ	E�@�x���%.	CD#�!{˄�D"�+a!*$g$�&�t���0�Yf��ig}Tu�hÇV��)_v�[��L5~{��0���#	'�~���k��'�E��ͩE�X9'�1x�8�d���;���=1�ɰ6���I���v����?@H_]q>�̫<B!b��=Gx��!@��i4A��H�/��07����PL��Կ�G�U����|H���U0-��cI�:Yh�"�*��Vt"
�X���ɢץ�A�΋��9㇟]h0�A�N�4a�*3n���Aٍ'��M�>T�ECL=<��g_93��y��|���j-AI�7dDCpF�A��K:�΢��@P�*�׈\/B/�<ZdT..�ݒ�uT�a'i�Oa����0��ae�3ǆY�����%� �p����Ye�A�����_�0<�dDE��(�8V�P)x��]��k�}a��;sQ_���bS�А����c�ɻ����(�GQ�(5ѳ����50cH�T�����#�d;���<lm��ZI0a�A���A�l��gn'6&�ё�X��N�� kA�f�(��~���e}i�t�Q�%�}��#�%A`a�gWͳ?@���q��4���i��1{ �99�>b��z�H^�i�q�7���Hъ��^G��IE�(���ӧdO�v�l�Y�P3	�<I��M>(�<a�`�F�`�`�>�*�M!��*��쭲M�͕"Y�>��NN�]�X���C�K���7HR�)b��yV���XQ��o.�"��EQE _��^��z��bEjvy���gv����ܲ�c���[�����(����̓ffnc��V��ِg=�Xq���r�ۗK�~٣5Pg.ڥ�� z��(�:�8��#]�;>��q�bEM�UH���������L?~~:N��*���s�A�Ld2y�j\3f�I��ٚ֎<0%��i��I��	�k���Lon.�: ��8=5٢�3�gqI�&�(��Ç�&h�Ҏ�*���"""�r�G�1|#��NcJa��{6cF��\�6}/,�kBuO�5<ͦɄ�>0������^וkC뷉��N1��C/Du�=��W�Z=��'��gP҆Fw�_��²�U�[WI������	h�T4�����(��$L~�@�6�Pz`��B��|(�JL�G�(g��!9$D�[C�$�� �(�Ěi���0��ae�3ǆY��ۈx�M��I���NYe�A���~0ȥ�Y��)��5�����M��n!�j�>7��H=���Zֲ��[K85�MN��(d���K;xDJ)�������T�D
 $0�͠��?e�M��:d?g�1�������0��P3>=n�c1����w %40��ٙ��m��|��}��ذ����W`�/	F���-���e5�YĨd������2�5I�2�`�j8Y��cH��FM�U^V�Rn�}��T+Z���zPhé����N:����g��ahA�\aaD ��<I�N�i�0�,��<2�-��V��Z�oODDII>kvB����%Y��#:�9�qw���1�%��b�é0�X��� �8�DQ����$*K�1������):qqB�]r��>�(.�8U:�8h�z�i��f:6`p��|o�LHQ�� kS�[����@N��;�� �K�Q�!< ���IJ�4��>��4��4�ў[��7�i��$�����	�%t��|�QI�|�P�,��aԸ�V@�`t�V��R�w���@Y	i)�� 1����po�L�Og��9���<���J0�6� �QgW	D ���T��D���h[B4�x
�I ��$�M>(�<a�Y�<xe�s�v����w��,�u�l�|�����#	'��I�>n����No�m�=�$��F���3"ͧ�g=���%�y��f�N4k������б�Q-����B/���Ot�>r~�&.v|�ѱ���Clh��-zZu÷G���>���_:z�ơB����RY�@��&�h�B�x�Jf�ѪR��k�t�h@GeI$m�N9�����Ez�/&c^��,�#ᎎ��¸�Ȧ�C�ьF�p���; ���E��3�iӡ�ш�MZ�	\^�Y�v�H�XZ8��Р����۩#M�F�4a���L>:||Q�x�,�x��4�f3A*�ҕ���˱�GI�eN��z0ﶏo�j^��s=�,wFj�6�����ODDII�Ï>���kiM�p6S�G�.���ī���$y1D,u�[��v�X��Qw�����Wxm�ٗ��˪���(�':�1"��B�;�]�L+ֆP^�6�h�y3WZ���Q�K��)Kr9�;�=>�?#Ȉ����/?~�,|g����;>6r#f�GL>I��Z[�ba����M�D��>;�h���h�����`�.Ї
��/�����+F��!=�ߏ1���)-a��DT(���gXCL0�K�:���?�A�'s�i�^VI-�DCd�m|� �)J%1X�<��7�X���xgY(dB�WW�R�paC�ۙ�T��vG�(�"�M�Д���iIp�|�����b�/Q�ȓ�#%2`0bk!O����i;�ѣcۏ��Ѳd����<I��i�0�,��4��^䂌U׮�j�![f�1A��5R]]~���,�� �+�+���:�Z%hL�ĘǍ�I�1y���QKmRJ��X�0Ӊ��<�%b���:����<���a��]w�Mİ��8��ц�y�Pm��L�1���(�\}?R^ac%��$��ҷ����Ų��çQ��
r������84��U�
��ןx���&�o�d���ՅbЎ#FC��#��{"��8��ci�8h8O�I��kF�8F�B}߹�Ff�p�0ĵA+�����&�����L�юK�:,t��V���,����>�AF�P�?���L?�> dh�&���#���4zat��f���M'G��H���0z=0�m�(�(�
��o��4��֍��f��Fƴf�����8B�3�4g4ph�������`Ϗ��j �4�4x3G����A��h��|;�Hc��I�h��4z=����z8����4ri=����z3#Q������eJ"�њt���e��F��H�a��tv=:Di=&��ãIѱ��z=��ѝ(�J#�ќ4�OH�r=$���}:�z6ސ1��ѱ�4����ѱ��G���3GCц�<I���a�xF��ِ��0=4�6�N�GF�h��{��za�pQ�3���oa�h=n��(�F�h3F�h��@���X !����+�O�"���v��
n�]�C��e��,��ڭ��1��[�5��n�f��뮱3)/�o4�������z����L���77e�g;h�5���U��a`���}Y�=����.�*��6wQ��u�+B6�w�%�͎�e��ubɎ�)'(�މU�X��&�w)�����ʿ,����ޚ}��|���u�O��γ3>��@��4�ݙ��^��>���Y������wvfgo������k3#333/5����� �x��e�.Ye�������I{{-Yd'��>vԋ�<$a'����;�g���N�� ��	&G��!�ߕ�\R�$�C�D
�
�1���x��J���E��pσ�|!(�Q$#��rK;����#�o8T3�U�C��>̺7)CC)���&��ҍe���C�8rRAL��&��޿�4a�vN㧎e���Zw�#A)�Xb:���r^T���{���� �¨�l�O���f�?'Ha�����<Dm��4p���BM���$���.�3��L���I�s��,h�Û���eLٷ�q|����M�Xm�č��D������0�g<|t���M0�Yf��T�H�R԰��\��,��0�L��ϫ�خ�3�������{�Q �� Lg����	�L#���g����oH䄇9=��|�h}�[�+Z��7z�#�N]��J��-F�c�^�w+���3��P�,$0�(�q.��%ɂZ^ߞ�j%�:��Gm����4I�Ɇ�1$��d�чO�ѳk�#���]���a�3��^�TD�@�c ]tg]�A�a����r�{0I �����,�"t��81152�l^u���a���c	'U�q�ƆV��Q(�G=6��D�G��i2:I��8h��GA�TBG��
8a���|Q��x�,�x�������+�z��4�PS!����O��*eB�[`�$TDL��P�ah9u�Y�j@�, ғc�w�ߎQE��/²�҆��;�C�'ԯ��j.����������,�t��5������)[�@�*^n^(^,t9�.]٦�ҴaZpH�qP06HE�`y�punG��+��� ���~�4�va�N��'pl��c�nO��2h�B�"�M��n'�Hm��8�4tN�2j�$�{�l�'2G��9�����\(�Ì��R�W����-�F�HӉӧ���xonyᙽ%����G��~��{L��6Hh�A�d��{!�s�ɂ"�P6�b90FZ�C��\9!�`83˩Ď��.�L>|6i��cxw|l�n�T;&�3�&��M����to�nZ(tgL/��us� ��D�4��V�>BRE��#4���aG�Śi��0��0g��Ogd	� 9��D�����y'I��vl�c�8s ��ۇc���,�����ίD�㰃��RK	����%�h�v�'�		;�=��N�����p ��%��@���59I3f�Kl�����<�*u\,<�Rw�$�D�LJ�Y�b�\�:�yA~D�p�9�����q��d)����K����Jƛ���D"Y�G
 �HJ<B��y)�,�8��G�*A�C ix�D��n�\&P��< ����G����?�bi�N��O�8||Q�Śi��8p���4��{�&�M ���_w�DAD"Je��է���R"uXڲ����Fy��gI��w��9]pf��X�+]Gy=H��>N�ݦ�Ϗ�N��pv�'�p䝄������F��|TG�JG��qG��tX��y�؝�iv�h��}}=6��G(��n������MF9����!)�b;��XU"d�)�>]G& ���I ��?$JM��M��^.h���%�*,�;03P��[)�Ȓ�Ԍ>D��jI��)]D�@x��I�>4����4��ae�G��vy]Or֭I�h5-:��}aD���$
��M����˩�Sd|�à�'��fkf�ctb�I=�/>�||�^�1k�h��=&fEv�⓫��h�ES)G5�����Ry�"���
G��i���B%2U*���d�� 3�����cl������}?.!!��'�#M�`#���l�n���Ã�(jI�4J:q�H��h��HP�
P�Z�u�6b���n�+��02("Q:�'�>D�
19K���x���4>,�M<a�Y�<xe����c��%��[n����o�����q�Ҋ����㙆�թ^N���z�b�^F��,�p}�Y|�:O) �gdw$v�Vڱ�w�/)��Q�6Eݺ�-(�
��ECug,Kچټ5�^װ�'ve�Մ4����j���A�+h�tj���x/=<�$)��??�A��i�J-@X���T��8��T�a��(c;�ӊW��m�Xѵ�(�ŧ.0��C!�i��p���PB���եri$�l6��0n��i�&�2k�8R��@@�����"6��|�4m>�uE]	���)���]ň��D"X֢ʐ�.z���5�U��v�X��JI,!�M�#'�&]��ҷRB�j�\��俆�R8�$�N�����#�Q���"ab<A��G'��t��1��0f���|I��i�f�i�L0����,��{ޞ�Ir8��;x�Z��>1X�W��xs��3��IO��r�@g*BF�9���i�v��7����=2+���3c�,'F�SN��Ǭn�0��h�,ZB���hW$�(���V��D�D�x@1��
!��H��w`:2s�2�O`��}h�7q3��z�Ko��G�ϑ��M��i�zL�c"9<��C:��3U��D4Y�ە�QV�2@k�a��uZqJ�ЉD@Ht��a'ĝ>4����4�Ƙae�3ǆ{>��z��qB�>�53ҟ�X�V$�#�%�8�P��������#�����C[2QE�jΩ�Z�(�r�aᚵ�ÉY���]�'��H�(e��#5�9��z"J�(�uq�@�>}�|q�r7����m���*fJ�W�~�����O��B=����pg��pC��Qӈk�B�«i��o�Ȅ��VzCDq>O0٧��=O^&�)�gɤ�޲�(���G�htx��R����9P�~�>���0�"���32��Ǥ�x����铠�_&���i}'��]]�<TA���� �I0�������Y��x�,���<�g~��@B���:���ٌHH5Iw-��PI�Ix A01��$q(9�+y\p}R0cE���%i�^K�r�|�<:IT%���Hg&3���M�ɡ���UW���_���EzU��+�|D1<�e�82׃��ǈ��>nץq�t gPx�����Z��`�83���d2>m�$�{��Tup���P�\����b6�12it���^��T�YQ�t$f�+�E(GW������ã��(g ���Ѥ>�Ck��f����aƓ�������G!�G�/H4�=�l���H4�oO�ۊoH���F�P�f�٣cZѱ�G��V�>���\#��5�D���e�@x�Ӥ`�l�B����G�h�4�!�FL#òH���G��h�Q=4��C4lz3H#O�����K#��?��F��0eB���4���P�}g4r?&��n4zl= ��I��ztp� ��N�/H4�4z80�Gf�P�}.�C��g"[�$f�G����8�2�m��Dh�����c��h֌��|����N�$�סǉ��:<F��4�p��l�#N����f�z<4���zx�m�����z�f�56�3F� �f��FƸ2�|62G�w>�i�+�Tn��8!Oi^7|�ȅ�9d"c�U&)\�RGE�r����v���[O$#Nu4,bn���oNu�v+X�uj��C7˄���X��+΃z�飗�v�]#Zv�^�J���vg��L����>���ln����H�VXUr��#�M6SG
�f�NX
몼}Q#��=۝y��͞)˩E$g�U4#��J4a�B{VZ�u2�u�	��`���meJ�/+Vw]�G�����HX�q0!��Y�h6�ea��W�r<�a�6W)Q]�����̬G�m��	��V,��2���Qؽ��;?lg���|�=)GF�rm^%v�j�\��A����m1,𡀏e{gh��D�v�#�YB�Tɵ�`M�W�5�G�6�?��{bۜWmB��DT�lՄ�e��v�����)k�ߣzN�������v�zi��wκ�����f}�c`=4>����fg33������s�w����Ͼ�:�C�s���쬲�ݖ\<I�Ǌ4��4�Ƙae��2�BUe�g��^ �F�m`;m��L�ˡ%R]U5ia2��[�e�F�XA�vslS)�mm�����.�#�&��T͹kZ0�v��[�����e�W]�.%�J�J�ls0˵�me���Ͳ+e��.�\UD�6v�͊�n�XŔ�ڑ�2��˱����Ι6m�K��0�t�6յ�2۳uik��X$9���:iڍ��,J���֍�hcWP��g2kB��A��YK��6Ux��aVkK���nV0��.S:ظ��[�aZT2����j �ۡc�n.,&c���V��$n(� b�5-Ψ�B��u
���f�V�Pt.�R��M�<����1X�$� ��{�6��\����ۇ��!�4�Ar�"����h�X��-`�I=�`�ɐnT���DJ{{����NH-uk6��5��V�*�6!�BqPq�R
��������1�.sE�{�����6��^GWOTΣI �D��Z ��:Ag�K��+g�G.ȎFuC���c�q4�h��2E{�}����?��.��A�(�<�@F8ã�o��J,�$ e����:�Dl��Ҝ�AA�[�pѕ�Ѫ��D
$��Ԋ��o�>�m����ӄR���H�c��͛}����j	:��B�Aç�:||Q�Śi��0��,ec�N]r>�$~$,�3{�PН�9<���+���4:t��6���O�#�f�¨�}���9�E�lgȯZ<�F���y��P�^���Q#)z���1�-s��d�Eh��d���,���8�Y`�O�=���k�)w���	X��è|�V&qI+ȱPpd"�8ԣ��k"�����\-|�G�J�Y(�@�bT`�G�[t���|�:��0  �H4��ĝ0��M,�M<i��,,6�WE�I��
��جV+��\wĵ��~���y=�2vI8����OU��}�R���ϻQ�ϕ����7�@��e-My����p��T?x��K�h�XD�$���͘EB���U�$�2���J:�-a�RZt�P�B��]�t��<�NYg�nчR�A<�>9�иyD�@�*��QN�Q���#�v8�k�᪃��.!�/��Q�i ��9+���ɣ�X�^*����$�K8|I�Ɣ||Y��x�,���Q)6G�)��&:D�lv�3���+��0��ϓO���}TX�܅���z��G l�����lz|av3t�?LLk	��D7����\Xcó+e���g��>�RQ��ΝA8�R?/�E5�ΐ�m�1�({���Q���E�^c�!��V�$P��{UxP�y�)�
W!/0�m�����D`{I����a��l��t���l������:Yp5�.�$��,�J4��K4�L4Æ,��C]��;��ә��[V����,�+
���B��N����Og�|�ggiD֚8u���#��m}T�H$�K�-���[�>uv4��Y���b�VD�lS`��P�	u3��P�n�\{�s����� ��wJґ��8��6�P����H>���n$�Q��82��j�s��7'Ƈ��É����X�#�,�G����e/��#��It eՍ���m�J:j�6��r
,�Ae!��4�O��S
  f"O���ʊ%;�Q����8e��󬳴������5Q������h±�B��O����Vݞ��?t�r��%��r(5���G��IH��!GĐt�ᄖQ�F�i��i�XYc(��C�,!��&YL�����X����*�Q��Q�uU�r��%��A�䏍7�Ł�� ��((���OL|̛�����ӳϭq�
���PqC!0c �K��]<b���g��3��˙|,&��d��+GA�<I>�ϔOI����6}攔QQ:�8yt��@�,�Sq,pH��d"T�	$e>8x�㦔a��i�a��X�/�����l��*�8�?��b�X�#	�ۆ���ë��6�8(kT�>�a�;O��l�l���������tP3Qj�L��R)��y�S�H����ʶa�Yj;�²(7��G0��χ��tf%�Q��I"W����,�1�.�d�>Z� :2	��Dp�"H&xx�(��R:���'�޻�\�:��r<�'��8�@�0���ic���.a�~8x�#I����0��Z?�4�L>4`�0`"�i>���N!$n}
 ��")A��Ut�>�Gh�g1Y�-E�llg䙧?�����l�C����Ӕ�]�=�5������$�r��B�,�RI~�j��4�A���׭��pe�yR�=ȗ6��C��9cGEП�O��o�˵�u�c����]�"o��F7+#�x�X@ϗe�t�`��+��c>�g��"2&,����;�\3��},�@I��p��G>(����4�4� ���(�Qa�����<�u�]�&��bLT���������fs�@l�i}��{�XC��4e�v��^�{
ʧ���y#g}M���y��s�b���9Ҁl����X�e�Q�2��4��e����5�an���Ҹ���H��!k��GC��>����[|�v뙑�ǑH���Z>���FJ�(�!J(ב�#J|<u3�#�C������x���}\}��|�,���<�wb&d�D�4����簕e��D珑���#���^������odi�݁�8��g���.��A�(83��Ƣ9aQM�NdĜU>�(g���x�4���g	�j�I�q6��4�~�� ��Np��Ǌ>,��4�4�e�2�( ������Yèrt���{�i�����b�X�#���nC�c;=� '�o�0��`��]���d83��q�KD�V�N;^��=@���7�@����l(d�cRQޢב��S:d��:}_9*�8Y�+D���1Y�ӈ�i4��@ͷ�>dD�n0ځ���2I?F�B)�/�E�~#î1���e����ǈ��_p`s���jT���V�����%�;܆�ԩGôV%$A�	����e���yr��K�.���K۩[�Ԓ䗷�Y$����]ܷ)~R��)%�mir]]KR]�y/%콖K/eչd�^K%��}}.����W�����.���^�JKR]]Iww$��Ieܗ%Թ{.�K��wrԹ.I%엵Ԥ�0�Q��a&�if�i�Nx�n[�-Kv���ݩJYjW��jZ�nK��]�r�^�^�����{u)r[�\���K$��y�w.�[��+�������@�?����߈7��5��٬�4Q�8S��0��nh�c��m*�X-)}/Ӯ2w�d墹��ʻ%�au�/1nʈ��-V�)kT��]��rgh�s�ַ
O���xΘ����ۈ�Қ���+3`��.�"J�r:��We�cPCF�=�)ޥ��\�
 n�Fgb�glv��'Mh�F�um� 9x�f�2�mӧ�n�J��]u��v�Ϲ�}����f}�a����s�fffw�����l���s333�Ͼ�8��s�s��xg�<p���4��,�M0�OYc,���=�c���" ��"��fF�,T������c�C��k̃��%�y��H�82��;7�|�%�#V"����3����K#����^�dK!��9K]`�}o;��#2�
)���Ǒ�m������_A�P��v=^<ã8᣽Gutk��q3�<3�1r68m��æ�3��qnţ5B4�%�}H�yHt�� ���(��M,���4�4�e�2�(�N\"&3��t���8��L�JN~;�x��u0m?}��b�^Fr����-�>�؏l1�᦭�á# �<}��`�f?||K�-�Ҏ�MH>���M�$�B�*�Q2⿻�Í���<�Dh���e:u�8p���R*Q� pm���:u����f+Ӂçȟ|Q�2�i�̂Q�	�:O�#��.̰n!�S�I;E^��GB�t�<4�)q,��e�a�E]r�;M�'�s���#��L�
8t�G<aE�Y��a��Ye��
#G�Cr&c�P��Q���A%V؂�έ
�Y�t����������A)�˭�,C�\ �R/0&�g��+�� D�����z�W�Dy^Y�O�;��ӥ�D(O*�]�s���ۥ��Wt� ����d�+R��˱�CF�"k��C��x7tm�Ӎ���R���n��>H⥃��nڏ����;UI��#�����o)_�)(})yt���xb���R�N���%�����D�p�����$M(Ê�^���5D@4�0e(D#	Ym��X���C�k0���x���:iK����R!q� ��һ�pG���q������.rNW��!YC�����g�)E�5xD:��E��Ɔ,eagNp��,��M4�M0��dp��A�VDB}����ys�Ӆ����(T�,4��K��EQ��G��m�0��i=���M��<��k~)k�X2�߃�8Q���.C�F�JQK��J�V@Y��J8Y�kpq�C�����ߪ~ql��+�`!�0H����ł15�i�z䄰,�_I4��t0�M\9��t��U��a�\E ?��2Σ�Q!�8AE8x�g��,��M4�M0��d3bؘRr�'����.��'v���A$^K�(��l8��(��)=��z�2�D���o�����J�j+��h���'U���,,�����q3"Ip8��-o�0�h�J�|� գP��9,ds���;$s�@��A�x�]��R(aH�0����=W�rx��G �cm�%���|-E#���0��8��ZR$eYӧ8|x��>,�M0�L,��Y^�-�c0��Jm&�XA��" ��"}=�\X��}9,i6�_y/�#��("Af��a�ⓦ4��i�5a^��W���>�hI��E���G�����J�T�E�mPάF�A�I�8yA���z��Omk�}]�z)JThR
�p�g���>`1=���ќGVZ�ϳl �w����#J"G_1�@0�(�N��PB���(�AD��t�g4��>,�M0�L,��Y�Hc�S����"�R�R[���T�����b(����y�g�u�u�a��i^iT��Fݪ1��$�+��y�����k6f:������WJ�t݌�ݾ���sEV�u���ʪ��*B��H瑻����c:����
�y�+j�(
�'d��\U�Ѫ�ìoM�ד^�xh_X�ZN�噉a�Ï;O����e)���GO���|��>�θ���q[<���x�#�B8.,E�fP��q��<TE�"C�p�T�V#���>7�gF��-�e���|-t8Z8���媁�g���M�`�}��uG�߼�8�}g����Z��Z�8�/;��y�4Zh���u���~�MTqZ�x�nk�� ђA��N�p�O�(��M4�M0��dW��Q�-Z}���zI)��{zg��+����Դ�v�����kҎ�OS����Ն��׳s�>���ko�5wqGn�`O!lJ6|b�yuD���>����8h��y�8�OZ>^��ۇ��R��#d$pk3�n[)��W��[��40��)$���AH�h����"#�x(�.ǨjU�JRo�I8��n$`�ce�T�� �I:Y�M>,��4�L4�0�:8e�LQ�������LV+���<��,�m�Sm.���Ϊ8��ȵH��MmQK��)b'�6��G �3��4�����H彁��,�}�:��P�������<���~�>jt�
����깤���u��x��D��D�IΝl�>��cl�F�TOK�8B}"[oů������� 
�>8�Ԓk�6|-��OAՂ����2[Դ-M��A;��#�+$ex����>4����4�L4�,��AFk��h�����s4�Wf�L�:�b�^F}�g��`:\�>Pw�E��G�:�2�o�(h�(m����n[ǽ�}`CP4�%I%NĊ7t~wv���r����l�������<uy}����P������Q��Ͼ�a��g
%e3�+0��tp�,�G�B�i
�<t)����!�D@�,�jc�D.�;G;�GX������<V1ڒq�cD��]:�[�h�ӕgTuW,�J$�M9���\�}ujRKR�I%콷)-I.I+�,�K����չJV�)JRKv�%ԹIw%众��Y{/inY,�r�Y$�^�ۻw�Z�W��a��4�Ěh�4�8aT<0�\�˹.K�r\���~ܵ%.I%엵Ԥ�$�$���ud����u{u-�rܷ<mI���C	��I��pӆ�4Ӆ�t��4��A����.��y%�I{<�ܻ��(042e��v$;�hf���8�PHT|YD�Q���.�3	!�-Y� ��w�e�܏U�[��R��*Ve�ʿ�(f7�X]����H����װ�*:uUq�R��J��Z۪N"P�:�ca�J�sB�*X�b9U>�d��
5�d;�y�R���!a��0fIX$ݻ�[o,��ѓ㋶���[_1$`�Uh��p p�XLg�g9[��T��!0��tȪ���uvN���8���&mL'7쬫p2�j8�$$*EU��
�Gfq��HL��)Q��� �duU]Z3��*���A�&t���K��if�:-0��i�F]�m�%�CX�4�io],��u%���r�l��km� Vorn���&��Z�p͠��V-�%&�aC',!]i��5�����:�}�pcg9�9�Vffgy�}�p������fffg�����:s�wϺ����3��t�7���$�㇏Y��x�L4�
,��AD���h�9�930��uiE�n�`�H:��h��]��,+d�c`Q����2��`�����t�fl0�4V�JM�WDm1&#t�.H��\Dn]��X��.s/$�V٦Ia���`��Bv���H��]��F��Öe���j�ŷL<���`v�[c�lS 31%��[�B���w-av-���2mn�<�V�y��(j,ٖg6��pa�����K-	�V`F�n �צ&�!;nI�f&��m�m�斚��#��5)5I���n6pʮ� �Nh��dֻ���0��ۆ3l3-���ljknw6%�����u�p�����l�6v�;�ґ���y����M��\�::��k��Ҝ�&I2T�46�en�8I��V+��������δ8��k]���n���h���8>.�e�Ó/̃k���z���CK΄a�;sS����V�9_Q9�V�)�Cwnҽ�B7�[�2[�Ulꧺ�1�8z1�DL�WW�|�qvI�r�৅�����85┐����~m��\d}�B�J����XУ�2.0���H�������[*��g�Jk��C���AH�F���m��%#���^��ΣI]8���!�L�x�Qp��,�@�]���XPcV���ɦ"����`H֒vK#�t:X� Ӥ�4ᦟif�4�4,f,�n�����Ӭx�L��6�2yE@Kq��AD�-p���\�E$�_�)�����3��$fZ֭f�4�k��{&;�8#�<d�9�ކ��B�^q�ӡç|�Ge<~]�p�t���6��L��'��ncteD���� ��`��&8O�v�a���*�|�!���-��Μ����OǏ�uA��w~��q'�����K��|�m��QAE��$������ϋ4�i�Yc,���u���_�pfa��f&��U�O�=��x�8x��0����힬Q�W�m��IpB*I(���ZZ��v����e��6Y��7-����6��ٯ"3��0fl数X3��E���[�I����ߑ�H�jB�x�#�,!�ݝL$����=�ҌF���=���>bI��{�HTu�q���i�b�)J��	(g(�N�p�O�>,�ƚa��P���X,�7���IU*:uc�����b�^F~�}�o���+���Fb�p�<I�1���:�Gp��JK+��_�Ʊ�yuw;��Dޓ���m%S��E#�Б
�kI����B7��`oyУ��zr�����Lxh6d�&�gh(,�)-�gK$k���E����O�g�%;���L��~."���I�㇌4�K4�i�Yc,������#�9�+�T�5�]UCT�&*�g�a�o�=����7x�ڲ���^[�-9v85)�&-f?�,V+�co�ʾ]���]�Ƈ���S��x��1�N��!앫1#�}U����N5j�z�W��X:�s��,�)�B��2�:�_Z�U���Z���Ow(�\��u.��o�tʥQS�����*��xlo�QA�֜��:�tF�K�l�WTLǣ�)#�h����~E���Et��(3�
1�xs�}��i|�����!�Lc,�<8�����!�@^�`u\��$qA!%��I|t����gO"`�g����>�JmiA�����[��'���� ����o��� �Oj�=ƛ~G�՞�""��XQ�� ��K(�fY�x�L4�����ãs3"�)9&Z�D��;��V+�Ϝ���h��o#�O!Ks��X3����qO`d8co�J�����~�� b�؂,�ykl}ТĽ����KV8�7����Ģ�(G�O�34�v�s���c+:��G�����C����j(��j%�4�JV�p��7��z�P��8B�s�q���&5aW���������~m���j�ࣇ�0:X� ��J(�g�|Q��4�M0��dn��Al*Ԍ?1X�W�����kR�ʇ��3I"� ����A$�������]c�2�/E+���Q
�H�䃞��f����j\Lɞ�b/�<�I��{�{h��W�!�B�1t����Nx-�\���W�BQ�e���`|���D��7i�m�)�I
�Ux1w�>�C1�K�
Yn����X� ��0���4��<i�i�X� ���G�$tj�e���`>���ȈD����1�.��`�*l�I�۠���cM�m�an���JSw[]ݺ����*&�}�<۞h���t�h-z�fe��c�&��y��5����<��O/=k�4:4֢�$���%!-�mI�٣���dن�j��6�;:��&J���"W��B�P�t%*�c,��3���TJ���h�Q��{Z�Pψ(�M(�fY�x�L4�
,��AC��&j�H�u,�110�(ӔMe٫��E�J�.B�*g�ĜE,���}gC�ֆ�ڤ��0m�q�95�l�\����I��a��`�w���[��-OF|Ʋ�ƚ��kv��e��ʴ蕒���9�	ȯ�zg\[W�\�eA$�\󭤽�u>�ԅ���AQ�+�9�n�	\ZNz�^GE���*
�<bMTܦ��w*6ˉ��T3�=\����Q��GTQE��I�0}F�}V8���e'�(,�Aa��;h�m:0�̟>08w��0�-8|���)}+�]�Pv��>c(�aF������d�i�|� �������'����O��M�l��M*�h�x`!�q?�����y�l��x��Z��͘4ht��A�ĘQ��>,ҍ<i�i�X� �}� �,����-��V+�g��	_x}��Б�[��7���,�ݢfgS�d
^DGTD�����Ө�6�:�8Jd�PH��R���m���a)#��3M���7����	>X�yz°,�dx��ryKq�M��ʠf��-�;>��I(��?a�Ϡ���
��ȇ�uB�,8��C��%Rg�4��r�ܲ�]^^�ܲ��wԖ��$�Y-^ڔ���$��Y.�^K�˻�r��+�JRKv�.���]KR�K�zֽ���d�Z��Y.��I%����ܖ[���)/d���}___[�����������]�r]K��չ-Z���$��Y,�rݩ-I.Ie�K%�众r���Է-�v���]��R�+�ܥ�n�Z���K��˻4�L4���3M0��0�2I/n�ܻ��)JR��a��
�'�9�.v�+v돖S*�DO��������N�8�$��v�Zȕ
B�s�>J��Ӯt����L��#Վ�Aϝ3
�˶HM�F�?�}y�|+��a��Z*i���ih���<�楄��e������Et�vֲ1
�����S�)���E��]�a2�hJ�.���y�/�!m���&V�p�(p|Wҷ���v^�ϻ�������s�}�����>��;Ns�s��ffg����p:s���n������a���s�}��-Yo5�������K4ҏi��aG�dS~���b��^��}[u��u�( �����s��7(�����5G���j 6o�:#UD�'Ȳ\MR2 ��>�(�~�| ��H�RUf��n|�g���!���uR����GNM�����t����Ѽ�8�}Ah�7� �
���@@@S쌲�\�P�T��GWx�Y-��z��*G�m��WF6R��8b>Z���jB�<�I0��>4�M(�i�x��E7tp��Ɂ�KJ��}��DA��O��#��Ib���=(�����g���W�|��:7��#��1q�B���ޖ���b�~�@�0�p�,P�Z�%R���y|��O�hY���yc,�����jq�Ns��&t�)����G�#Z��b�u_|?.,��
���z<GW�Y*�ߺ�C��o	>$���|i��4�M0�Ō�)��e�'z���Z1a��1�o;���Q�z��k2f��|#�NK�xd�J�b�)�,t5#4&�&�a�X=t�H$�K��6�Q<�N;ۯ�����X�����z_e��ќ(K�U(r����˔�g�I/7�к�y�V7���P�ۻ�wL��RU��4��b7�j`�ŜB��b��ӳ|�1��������Vl�ܺv{=��S��t�`1���|�wdBa���,|'F�$�������qfm���EK������̓�h�;M�ʨ������+��,�o�.�\e���d��:���p�a	�f�P�Tp�V��_~1a/�������������ë��>d����P?.���ݒ|IFY��,�L4�<X�"���Dk#tª8|O�f}� �	A�i�_�q�Z`mNJ���>PI��r�6j4��u1b(��Q�╬:5���Ȑ}D�m���gIG��5,J�Š����?�	>o����s����4�} &!�(o�:�e���d������o`�'ȿ��qb-rC5�/�-L�q< ��)a���B$C,�7D�I��af�x�M0�L.|��{u��R^��ޱX�IxG�M�$�&L��4`��`�q��(�Y5�|x�w�Íє84򤼍<��D���C�lo�_v��EK�0Tp~��Ͷ�%����w�ч,�@��ᅣV�4�T���^5b��gQ��5.""!D��T-����n"!�\�B�@x���q��L�����a:G��&�ig��>4�F�a��Y��Y�s�X��(��v&�ND�,{��b�`��4B���o��(�������yq�ߏ'V���%�'�"a�7,�#��B�	u�yL�?s������|3���[��Q�,)B!p�PԅG�}\�k���lm�p�����>���Ў���(�<Z�(^r��Ö��\E<FA���,j�9��R�����0�^���2��tI�%�||Y��4�L4�<xe�M��4t�2��|�.�6��@�6][�z��Hm�x�F*E�f�׸���-R�2��o����A$^��e��_e����|ĭ�Ub��ʛ&:�we�ñ�E\r�Xi�
ؖ�on��A����7K�� ��z�<�^Vb>�J��6�]a|C�v��ۭ3)�w1dU��n�ѫI�����<b��T`�(!�:i���P�����}������"�GQ岎���DDC��������W���HP/�M���1���[>�9Lm7
�T#30�Ə�o�s�*f�XW#�r��,ɂ"U\�1,
�%xL��Մ�p3�u�a%�x��M<if�i�x��"��ۈ����<��{�lߞ�X�W������V{�9�~�!�����n��IF'���q#�`�na�=���a\08�֛y�+��tg�a��[����`K"`�,.��Aaa��b@�?�IZr���m566#6�r-�hh�����p;����.����2�(,;�Ll�D�A��H�"۲K$񇏋>4�a��0h�Fd�Ax��ǙP���^4"��Oʠ~�v��	 ���l��a-�7'���y|>a�my�
)}�-Ge�I_}l.G�-��~>L�Ȳ�R�7ϓ�!�%�&��!/؝S�N���L�?h=�C8�%�ч�d�i�ՇWQ>n��;��4��e���'b8&�"YL�I��(�|<K�m��68Z����p���'�4��OQ�i��<2ȡ�6Ȏ�� hQ���+��K�O�~E���	����'ҋ���~���L.W9Ɉs$)��|���0���h�G�݆p��Y�(���9_8���'I����� ��N�=�O�d8q�><�����_#�Y%|�X|(Y��]6�m���/lh�uB8��I�j;
FA�O�:;;wr˖��-I%ܒY/-�K�rK�%���$���^]]�[��)JR��[����互�ܗ��Y/e���,�<���Y%���{wnInK�\դ�Yn������������)I{.��r\�.��jԵ$�rId��)u-�w.��^�,����]˗WwRܷ-�v���/-J�V�w[��-�KR]��{r�����K�ynR��4ӆ�i��i�0�Ζtä۔�)JR�ի��y�|��:��oKX����d�V>�j��t�6���p���~#�|�����rR8Ѣ�S
خ�j9Ш��u'[�#�OI-����fm�-��HrIJ�J�Ѳ������4�N�k>���<W��AkՑ�s\h����̷�WUŭ�Χ|�?uT�#�6P�_/�3���m�A�7n�TA.q��4�)�]���b�Y%U=�on�8�K�����vV�)�kF�]z]�l+9&h�;|h6�Ak� t!:� ���uu[W`��<���UЭZСwp"D�����U[`�N����X��D��Y��� �!PEHeݑD�r�*-��|oq��+#J�]u��癔[nA,��^ȪѾ�Gj��.�?�+Y��<���{c,[��ڒ�r\��y���̑�f!�S:u[ql�%�Z��-�Rv�-�Z	/3L���n ʻ����]��e1�M(�9���u��f�����|ǋ/X��Yhۏ��I�'K�u�ޭ�uk��//;������ߞ�7�;��9�ڳ333=���ts���k3333߾�@�9�}��333=���ts���k�e����˫.Ye��i��(�4��e~[sP��\D�8�ݢ��2�����`a{.�CF��*�5e�պ\�.I�[��n��k��M�1��w6 �5+��lt u�۵��6XBP��Z�*�L:�E��	n6�m��I�0��M�KxR�.(�5���k�1���-����ZZ���`�m3�mXR�Q�!	o��d3�c�Z��Z�lBiC���jB�C�fS�U�X�Vb[��[��[�a��:3g\]aRg]�ky���k6Â�mn�t��a	��,�+	�d�3M�H[,�[�\R���1&yZf�V�K�[n�u��t/(My�3U��s�-"˜�2k�SB�.����bE�s$���4�iv���\X�������qcT��.����R4�?]��	 ����?�h�F��v�/Pճ��s��j���YVz5�y��h�	NE].̪ȴ!���ØU,�"9��)+���縡��4����j���,�˂�.�h�-
&`b�����
��'z����v^�"���O�B�E�O�n�%X��G/�8bt��}S���G��x�;�&�d7����p!�^'�N��%�ֲ�q���s�xP�{�~�2xX������y��k�-���i�{=�q�d-0>^�����ۅ(g�PB�X{�;���3V�FdG�&���>h��'q���GȮ�3��oǯP3iD�$��<igƞ4�L4�<xe�%�\LI�4J$��9���r�Y�rz8cch��O*	�8dp��)O�p�^S[
�:*Gtj���c��Q~\6/<�m�ۈ��w�=��IXJ���!x>CV���G�>:r�f8g6A193�m!\�V�T�b��~��S��<?z��h��q&I��OL�>!}���A$�x8���C1hwQ�9ӇJ	�m����������2Ft�&Y��Ǎ,�OQ�i��<2�$��DG�y̷����y#�br�9��*#����b�b�@��o��� N�����)a�}B�Q(��o|*�ȓ�1>OC�&�o��]��G
���g��	A8�Đp%w"�I�]ϲ�{����_���O�>E�|�������t}Z�>o��2��6��L�S��D} 5����Hq�"�b�<H�� �-�α�J�����{���g.g���t�'Ĕp���i��4�4���a�O�2��\�ث��2#P1ɍ�����#��� aU�4�~�=�Om��1Y�ڼ߲��af=p�j$�y4i�M"(�)�����_t�
A���<߳���w���f9.GWlEj�� ��DR:�|��A>(��A�Bi���h�(��g6�5R1��:?q��G��3�	>$��ƘY�4�4���'F>C�{�y3L���E�F�,C(�0���vI嘲����:Q��N?,w�Fؕ��!^{�� @��&j���R�+�����F���pܽ��WD�|Y��O`��h�f�<�1BJq`5E�{�嗜g.fѣ�:�]ElQ�K�UTy!��-	WB.��)�C���YA51(�?|`~����k���Ũ�t�.�v��\,)QU�!����8��~����,ʌ3�<7��I��?x����I�DPBK��N#ʗ�:������w�~�t���]f���X��jz�:|3�I��t�8��"Jm���:@�$�'�|a��x�J0����h���KV>� "��1F�=�5%7/1�����%>�RO\"�N�ƶ��>DB0��~q3ȝ8�P�T2�rm[v����l�|�|��
D�ūtl���U�����;��I'�Qh/s�|���LT��GZWP��M�H �W#nߺM>���ZSښ���Ӛ,C΃� �c�=�I����E1����5W=��u�V�L<fN�	<Ig<a��x�J0�L,��(�5�vadq�����D+�A �O����t�j)�w.������΃_`a�>��4�(�p���]/g���5��<j$���FL��}��8�ގ_ݞӆQɟCs.\�Ѣԝ���,��ʃa�I���a�q�Ԓ��=Ci�����Z��Mh�rb��`Ϗ(ng����\ͨG�����F����v�2M$�M8x�Ҍ>4�0�L,��(��m��po�ȇ.	����f}llm�"m�<ȇA��S�=��Z��6��:�p�D��!���7�%��$�ȷ/':�TD�˃�1�J��7�h}��
�H�W"FɄYc
%Q�|I$����`���_�zuI�/���Og�28k�ea��>���Lĩ4\7Q'���O5�Q��P;�i< ��##⺎/(�T>�mypg�$�%�0�i��4醚p��A,0G��IWR���v)��j��Wb�R)~W��EFWg|��D��Vy(���LF�h�1��	@��A �O��/�����_كW�%S�ק���՗7;+o��X�]K���6ީ��nQw�����A���d]Q�A����O�aq��id��Z � ��~�r��go;W��1��Q���ee�,H���A�b8Q�]�"�G��oIE�;�QO1PXx�X�J��IE���Q1%�����2w���4ů��bӣe�vcEޣz��Q�A���Q��.�!���>�D���o	ceB_��[�Ӽ���n���d�J:�����7k�m�[~o�D��D�I㆘|Q�ƞ4Ӧi��<3ãF����2¼�(���ͧƟ5��Ҏ#Q������E��>DZ�с���~O���S	��V�K�8hx9�����"`��M�*���,�����$����1��5(h�t={��nȎqG_e��%���G�d��?'�}t'q�J�W��J�z�����j�p�x�h���d��OtӇ��<Hσ�$�rId��)%�w%�^K$�^�˹wj�ԥ)JR��ܗ.]]5��u%ܹ/%�Z�e�K%��e켷,��Ie콻�$�%�$�,����-^˩%ܒ�-K����������W�V�}KRIw$�K�r�互�^�$��^æQ�L:I�L � f,m`aF�,�jWu�Krܝ�_�wr^��]���d��)%�%ܗ�__K���}e�����չJR��0f�<��c�9��d[y1��G;�ڕC;�Y�]��\�xB����wi�8hn��_�j�i�U�AX��P��^�\#���v�.�Nr&�N�x��,�;V�vǖ�-]��M�b���Ka3w�ZM"��F���4��a��T혪�P�a��ڻ�JQ�^ ��Q<eX�7�U���j��T���G�j��3�5nK+E��t{wu���� �ts���3333��@<��8��333>ϴ�s��~�����>����s�}Ye�ǉ<I㇏Q��x�Ni�x�#E�>�@=d	�A��[rH�N��|�8�(�A(�/
U��C@�J#H#�9ב��%���u����8�0�n���4QԻk�a��tIQ"�~q"�ƐM�����c�(~�61��V�*�WΜ8}I�-q|i�ߛ}G�/W|� �\9���ϸ�ޟ5t�w�r��̧�q/��M�^D�K�/#Y���cc ����hd.uH�$�M8x�i��4ᆚag��D��D`Do�m�/�|��i�!(���Dt���{ �r�O�jp���Q�N�S��)>�f!�E#R�>�����l�#��{ф�o�E������Z�Y����$��n"JX�Ź�����*�"��P|�>��9�2�����$4�Ϗi%�4���M4�iF�Y��<Y'gyU��w&��R.�(�����tq|eF�SM`�@��Zr�*�e*����l�wDm�8�ehjjn�)�p�[�˪I$�nn���:��}���׻����b��Ƀk.���}APT�^��맛껦c�6�W(]��r̼d*�t.�%��/�6�ⴒk����Wg@��E9"I!�(<���Z5y0�1bL�k��t�k�F��c<�>>>Y��Ɉ!���(4:����!'���i%&N��MP�x ��<C *��f'C��>z���_������i��v�È�e0���$���I�~��K�%��?�:�^������#̾���8`R�S���^��JFH�$�M8x���M4�iF�Y��<Y&
 ����A�f*+�|�Lk4�� $P���/$��	�Ђ�l}G|}	|�������=�;2'#J9
H Oy����]?W�wTE�ZN��4��V�3��a�ʦ�lvs>PgT���}S.&dpJi�R��^��Ϭ�@�������b�at��3�y&�k����h�x��B����+�'Q߼�!Z��pd�I�O><iF�i�M0ҍ0�ǆx�N� ��Kcʴ	aN��@ �~>+%6��b�r8Lxx�y����Y�����}!i�I��((��H�Ee��Nf&Yɞl1��_G�����=��5v����d}���tZZa*��	-�qj���p��pq^0KP>�H��kFyG��F�T�$��Ý����"Ƌ>�^�2v0e།O�$�I(�x4�ƚa��4��-|<�!�F?q$�HBQJ'�ZHY��û�h�D�$W��>��I��B��%o��!�N�&$Uxp���J�C�^���Ũ_Y�֮�F�g򜓈á&���q�����>��&�Dz�-�T������wt�C2`�04�R��m�]E��>!���y%�߈m�6����nCP[�k����dvl�Ėp�(�M<i�Q�oŌ��4U���5t}|�D(P�nb(�4�z�e�ʥ/�Ys2�,6YM؅��s���G�J�Kir1���	L�"}ĒIe��k4�4�^���mY	)�.�԰ou���Ъ�y3��b���8{�9"�-�<�z�4�����2>�uf�c��LC�el5���MD�q���yy?>֪R>��e�!����D�k{D(Ds�xYO�On�g��᨝p��9�,p�g��Q*��S\;JO������ӆ���g�Q��ӿ��7�i���=$	?��B�T�d�7��FM�UT��~����H���������>i�a:\�2�$�K8x��0�ƚa�Ox��y,��1&5�z�	�}�8�z��TZ�d�H<��u!�#�|�e�3:��)G�P7D*;a�>R#zG}��%�6vQ���\rc��Hg4�� ���L-���@!�ß:If�(�4��z����:l���}VR:�GwG�h�	�C�>gdY�i�4 ��p�I<p��J>0�4�I<i��YD��m��Ğ��lq�̈9�Vxc���� �$��J���֩�N$��}�$1E����
�WQ���w�xtLnC�cl���xh��}�H��K�W�G��������!7z�lD�i�2q�/�G�g�P�K���� ���n2�CK�%F��)�g�Y�6���+����_͐�DLFF-HN-M�}t��d�<�ۡ�h�FPI#4�O�<p�i�4�,�?O��'��b���X��t 	
���P�t�Ҁ�c�D.�=�g!���7��T�!(YK6��+���N�[��J�c�C" �X���>��z�m�y��Z�]�GWN���vXqp3ܲ�61���>Z>�әV��5����soᣐY�LC8t����f��h�?��?�?�P�W�UUTP0����������<6�������a�� �QW�#����4���4�b/D��(H�@���0L3L3Ǒ�D,�0QC0��10�!1LL3�00DL2CB�0�0DC�0��D�0� L�0�0���0�0LI��0L0�2A0���II�I�A$DD�B�DED�@�D�I���DD�B�D�1�A0DID�B�� DID�DI$D��L!AL�$,D�$DADL+ID�KDID�D$DD,�DD�$DDIB�DDIđ$A1,DDKDD���D�DD���D�DDD0�D�ID$D,D�$DKD���D�Iđ0�$ADDD�$A$DK�D�,IIDLK,DIđDI$DDKDDD$D,�ID�$AB�ADD�$A��D$DID�,�D�D�A1$,D�D����IC$0�D�@A$DLD1KD�DLDL,�LDLI�D��A$D,�I�$I$A�IA$D,�ID�D,İI�0A0�D,�A10�0DLDLD�D$D�I@D$DLLDL0DLD��@@ALDA$,D�D��L$��������� e`d����$2�H�� ``````d `CX�M@���
@0!"@��F��FXD�11 Hj� ��`aVD��9�jҤ�@ʐ0$	*@�2$�!��@ʐ2$��2�	��&�ʐ000��@0��2�&*��$�@°2��@��@�@��2� @°2,�(0$��02,�"���2�����,�@�00� �2,# ����� �@�H�(�@� �@��*�J��� ִQD���" �
	
B�0)C(���2)�C�ȰȄ)*CCʰ�0ʄ2��)
CC
� Ȑ��0�0��	���0$20�2������0$2�20$0�2��!	,2�����#��
H�������"C#	!!
@���"CC+!��
H�#�0��8C$0C��	����C�2��C$)�!��a�b!�b��Hb�a�bb�d�!��f!��"Hb!�!�e�!�RH`�Hba�ba�f�!�!�`�Hba�RHba��Xba�d� �Hb!�`��Xb��!�!�a��X��R!�d�!�d�d�d�"a��Xba�d�RHb�Xb`�$�$�"�X"	`�	`�$� I� &�`�$� � �$� � �H �$� ��H	 &�	��& �	�b	�$� &�`��$�$�$� &��+�0D@LL0D�I0$I$A$A0$IA@DA�A0A�D��A$@L��A0D0D�@1�A0D0A�A�A$�$�)@A�D@LL0D$�D��,$�A0�$�D�DD@L�D��0DI @P3 ��$�2@�d1�� d��HH �H $�ێ�$@I$�,�$ I$�2@�@�A0I�$�D�.b`@�$02@��� ���300$���� ���)0L3 L��0��I�0D�0�!10PDIB��L2��_�s�k#�g�e��`����2�� "�R�L��L$f��	��v�Waex����Kq�Z��"�fm��K����E��π`bfIa]��s���)YU�[���3���Uۅ%�Vp����B��������)�
�ê���s���z��EG� .^0�P�d����q�'C���x$ְ��k�w���6�b�^P��@T �@�',���" 5T�ȱ	�I_���>O�t!���2bv���LLO���������~=�X��?�鮯���x��Z���÷�z��0
 9�4hJ��@֢U�!�D@�P=\���@�P%@i M�p�"�\n��!3X���GA�����?��x?�C " ���(�@(�@��Q(�Q ���������Ƣ�J���sVjp.�V�	����S�����N*r�0* I52�5��]�W�[��WI��C��S�~]]I+u�ӥ�*`d��P<"B{���rc,]�&m��+<�d;���!�,��Aט�6�[iYi�K `8�*�A���f�Ь+�9��0"sv����Rx�)a�^b�+H�P�" �ǋ��Q�����@�� @���'G��8� ����3c�ba�&?��gA�>/N����:�f���7���y>	�a�T �RWcٟ����R�R����S�!�@1ș8�Ӧ�~�g��A��rvTM!f)��e9F��Ml�8���c�ԁMd���{GF"\�5����9A
��.���X:M�ʎ�,�����d?����?�q��]��P� f�s��f��F����]g�`����7��}sC3	3������ �3��!J��Rt�q�(	��Sq�G�`�o���C�?�����|O��Ŀ���a*@f����J�0�3"���aNY� ��k S����47����b�$���ߒ�k����dik�
Sߴ��D��&�
]zW�m��ܑN$+M�@