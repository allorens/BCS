BZh91AY&SYnx�L��_�`q���"� ����bF��    ����(��`Il�[-�%J�Ճfj�D��ٴִh2�lm�)-�Rm��U6m�F���Y�md�!J��bR�f����U�g�q�Z�ѥ
�Yi(�mXb�Y�V�Se2��ٴ,���ImkY����`�f���j��P�6��F-��֪lͭL�lIhR�[
�k�XU̬֭ęk6$V�U��jh�5MZڪ�Ke��4�[M-��kIV�5�ڴ`�eI���Z
m�������I����Kk#m��t���,�-�   ޽��Y�t퇣��t���v��m��W��
{iv�[Eڍ��3���w;�tj��4��^�Z�m�s����v�5��w�3;�pҭm6���U�����  ;流ٍ4�{���tҥJ�9�J�*{�6�ȺdDn��{��^ۭyᎪU-��U�Q�R�R���zTvV�/W��R�%n��o3�6����md�2�V�ZX͍jT�j��   >��U)RQ3�k���R�[z�;޷���O{ս�{۞���ͽ�T�B�J�{��S�jT�{���)�+�*��J����%�)U)y�n�h�T�{ʊ�V*ٍYfi��D��   ����U����IRU*S{ڻUS����N��PT�zR��%{��o^�����U�ު(R$��{�PSٕK{�ﾢ"u�}��J��ڊU)7���k6l�YfkZ!�ckm�  ��O�IR���}�Ғ�����;��U��Ż���IT��i�����R��>��(W�*��K�7�*T���s���F۵f��>��2��O>�ҕJ/gd���Y�-����l�m�  ���-�*wJܦڡ����R��V��y�j��${n������]��N�+�j��T%RTy�[��)kJR��ms���٫��޴�*�)v��*E/m�&ke�5��L�km�|   }�{�����\ޞ�yJ�Pm^y���'m�t��Z�:�R�wz^�*�N��nT�S��7��m�Gz��{�z �yn  �;��@�.��X-�Kb��m�ٶ�   ��})C^����U�U����Em��{x�J5Gy�����ꚩ�U�`�ޣ���U]ʳ�CG���S,J�m��m��@-l��  �>�ER��z� ����Poz�z��S��t��{� =��½Uump�:S�ǎz�ooa�JR����Qf��2&Ml+m�ʵ���   �}}j�g�� 
{�^��*��W=Uz�n�{ޅ {�x=z*�z��tz���@ 7��x( �r�M�|   �   ��RUP�2&�4 �F�O�1JRTMd���i�LA����)(4����&L��%J��2     5O�LJT3� �4a0�L���i�6����A��i��G�>�c�#�XQ�����EMZ�e�y�����W�#n��:w�{�� =�y�$� x�� �cl~��m�����;i��W������1��C�����l m��!�l��l�}w����������96���͐�o�pِ��8�d7�gm� �o�6�����g�M�d��� 2�@>gm�����d��q�d�v�ɾd�q�d�M�d흷̛|�7��>d=�2m�;o�6��o��|�7�;o����o�7d��&�3�� 2`����~3��;o���q�d��q�d�M�gm�;o� ���� ��ck&�86��Ym�;̘0|ɶ�p>d��Ƀ��`>g`����������2m������>d̆�}���q�3�������v�o�`��m���`>g�p>g��m�́����,�1�8���6>d��@�>d̀`��03� ��m��pl��&6� ��;��>d�`�������c�|� o��lv@ >g�8�c�pc2=�����|�0c�Lc2c`������}�����q��;c�C>g�����8����|��1�&������>g6��cc���|��`��1���l2�� �;co�6��@>d��87��l�>g�!g�p3������o�~r���o�s��vߜ�?9 �������87��2�!����8�|��L3�|���8�̆>d1� ~2m�&7̆��� Y �ɷ�L|�>���&;8��x?��3�*�$���:�-�[�w}(ԭ: �m*�6��1��-��]�TNUf�D���##v]lF��n��7*Z{ux�)Y(ٗ�^'�/f���h��S7XP�f���ݮL't�U�1���ռd�A�s8�����n�fV[�q�Y4Rs0�v5Q��o0�������gQ�#T�u�c���F��F�W��2�n��A;y� �ef�0L���}jB5�}V��]F���9����n��l��%ũ,{$x�ͧ&T-��h,�`4-�
�
�n:�a��%YVk��OmkZy����)�R������Kk[�d:*Zu���7��2�̄E��4G�,�7e@�n��Z)1�A	��=Q�����vN�-`��j�9�ԇP\;���,9�J�G(yU	ʗt0ca�M�N<�~܇Z��������aV�˽�z%�2��&2�ݠe	���c4s;��^�����[�6�+Jؼ�ۭұ$Τ�yGZlW���a�&��vh�%6�#c)Q������J�I��=r�{ 0��hV���n�+Ywz�f��˼j�	�J!J����d!s1�Ip*ӄ�Sv�il�*G � �-N���*�m��6��P`��k��ө��r�c{�!���ҽ:l��p�W�;rI�5;Z4�F�L�xu�ʊ���u2�]L�(d�Z�<�Cu�EbCMD8jm�oFY{{��W)=Ƞ	4�L��e�pji�%kz7�ec�旛@C����]fk�$'�V�pi��+]M` +u�[2:����=���`0P�-ٹ��1�.Q��:3;��q�MX�����,ŕ�j�N����jD7�#E�����.�ɎJ���#�B\{zp�&6��l�1�3YV),��	ռ	*�v�W�#�.,̳��<3mլ�V��E�wR�CE<n���3r=�X&ù�,c��5G[)�1j��[X�VQ1�����en��ϙt�<����O%�f�Uvf���u���(�k�h����̻�sAG�*G��� ���h �Dx�0�ĵ[Z�j��,-t�a�W�JL׮d�˭��m��1MՂn�0Sd�(e��,F�쌂fܣ��2�쭺Җ�����%��ɦ�[�����:���Uښ�,ke�(-/M4�Mj{���l%�tmh{���m�X�%z�v3��%0��Y�lcDP�si��B�u6����v�nb��[C ��xF
ǐ[�l֫J�����ݩ�v^��
��Ɲ֦wkeH�f�����1ZwM,�@�B��^�Sʰv����rj�B�nh�wu`׆\�8B�cC��A�Z���{���S'��@5g�:%:9�w���YJ���L,q�)����G ڒ!{x]މk2�H�0�� @T�X�U�p�ƙ���-ѵ��n��VQ������r�qh.�;qR�&$���ĘZ�/.�&]k��+/�m9Z��bt쇃^\�8Lu�AW-$t[A�7�����2]b��*xe���&���6��e*���`��^<� ��03��]�]�C�E��ƭ�q3Wsa��ʴZ���Sy�0�f�4����mkA�a��c2:��Kk�tW�96�]Z5����{����a;yR �9�O1mR��T53NVEv��n��U���Ќ��a��2�Y3��!��+Kf]�հ��*�͕�
Z1\�t���(MHՔ�i��v�U��Y)n	��|۪+��7[�IW;��q�2�+n�^U�+�O9�pd�In������{�����4����Cv�Ţ�­��b˻+.�Rmd�-5�{�c�1�sC�Au���Zb� �v��JQ�L��J��ә��Xq]H�&u���c�):YX+
�r8�7C�P��Ә\����fd���]�V�>����{YK���E�����7OSR�@�iF�zn�R��6�}i
F�����ͬ�VVC�Ռq�e,Y4>�D�N$dF�d���$�כ{��X��#���+2�M�uz�pW��b���d�z�����.�Qԉ:w�k	�S^��-�"��v2)v��;ж�(�a�Xt�z�#jn5��`ںD� YQ����+0�wtM�j�r��mR��M�]�Xb����ϕs7Z�u2�ۼ�J�#]Z����if"	9r���攔��a#��Ƿ�N�R�:�mΖ$�lE������<�D�]Մk(M�D�F�k/J2��X�E{����GU���!AѰ��*���h:Ұ�bݺ$��(=*��^6��H��I�W4#�8���Q�)k4��bnZn,��r�+F�T3S:�=�Yp�C�_E���H�*�V�w�
�0�f$�v�%��[i��y~ܖ���Z��nS{�S�q(l8i[�Ԗ�4��k։�C4V�A��[��}�8�C��Z�=;V�D��׷Zhm�
���r�� nbG(��V��C֋��6_�w
�X��͂�0����t�9���3U���MU��UIQln��9���8RY�ed���b�-0�	2�U���4���>7B�f�٦��g���j��emnn#i(ke[Z舃��*�#��ޝ��ĨeR.ՠ�jDw�ã�C�y2�UR��W��sv1R�VC�՛kT�GL���%Pbe��9�l��2�6�/=Pnc[CJT�BK����X�<6ۤ�Z��Ӵ��F����6�eq;�-	� �늘�ѱEo0��1FmZ����UZ�����w��C%8op�&d4�\TՃ�n`2�������:0�n2dƓ�W��:�2�ܲ�̩���W&�&�.E��Kz��t������śX�=$�⮝�^��P�,V�5�N*Tr7*�a�{��L�.��Zy��׶���k$�M�^�t	Mw�45[���sX�+
�Xo^�]:f���'�%�+Y��,�gm��in�̸K��V�74�.�Y��eM�U�c�GF'U�R���2C�������̵,�c JL�7yW��&
yM�S�m�g��v��"��Y|��V���`Żx�1�f�[;-6$�Y2��a�f��r�	�ڸ/q����KUM�@b2;'QZ��5KB656��͗�z-e-я^�vU�/-ۤ�P2;MF6XݫZ6<g]�O/j�S+W+��,,�Ͳ�ظq]}V8�YșzD�L,����m�M���m�fHq"�BJy-k-UwıLVVl� Me��;�93�YN4rɻ��Hkh9��ܖR��u��ּ�ųq˕�Z��#Z��@Z��b�E���)�p�u�j�<zn�#hU�vh�M&1�kVm-z�f�f�ب�[�,�x��"���T�<�m�<Wܗk�[���;--�w���^;J�-��F�d:��V�7 �QjW��{��e+)��`aW��%j���?��2l�,>��dP{�I������2�%4�w7y�x���.Ys�vm�����I%���i9�(m��HJ�͗���	V�X�BѴsthweL߮�-���rI���^����>wC���yI��-�%Y�Z�+�PP�Kc�i͵C6��\��˫�個����\�5�`��m�.9*�zb��-j��Z%{0ԗ!i^٫�·a�`���^b0�E�M����`&��I�.0 /��'��6	+5�����i�6���cLl�f��R:Z;�*��7{��f4�0 8h[�WkM�w(1d�L� na��[l[3r��
� kwY�J}�ܢ#W1��vo�5K�-����0�BJ2�P5���V�퉫i�0H�mb�ڲ�q�u���))7}�vd�0��eRc[z�^�Ƭ�ˮ��R�^!n����١��V8sTtv/-ڶ���0��b�
��n;*M�FV¾9AO�h����Ř��������LnÛ��	7@f�j�kU�i	��u�13M!Y��3s\�t�O6�M;n�Rf�P^��F]��+&	�+��G ��)N��j��L�]�q�I�ڏ���G*h�=#�ޒة����Y2�J��B�^Iʭ%m�㭇��ū��4�5��m4A��l�[�֦�G�텪]����� Ӷ(dXMͬ�u�h	jI��L�2^:3���m �F"���kd4���v¨��k[�)<��j:�i��0�թ�/wa�@��]��r�ʿ��cs	&�M�ѕ�$����;Ym��F�((�utP<�(��qv<��AnꕑnT�W
z�`i�(����+`�$�ݣ��YM����!��XY�F���V���l���2�>Ku^��Z�(CX�Q{w"�Mn�X���Z4��0"��w
�Vi��"
�iYz��O�ˬ�mGb��m]�h��S�ݚY�>�Zf�t�����V��2��4��QfɚyW]'��B�c��T�֥�))��뛥*2*�WO0ȝ�k�+#�n��YX7P�-
z��n��Y��9���z�x�V'�_Î�����uY4%Kkj�n(�d5i�鬶�p*w�
�0
y�Ҹ�\���D�#�LFѶ]B�%�r�4�b��AF�1k�Qֹ]����a�De�A}{�:p�hm���8��w.�O]��z�ƃ��G*γv�$9ouHY@Wā�Xƍf��`T_%>���uCsJժ,N����=�bq��f9�f�ِYZ�.91�&c�\r<v+v������GvC�t� ���F�IL��ef�0��IVc�;�:�],ԀO�t�`�uup�B�(T��gZ�*PY�I�^	`�������imV	ol��Gt�v�Wm��f���¤�������Wa}�Q��c뗯^-�#�H�cWX^�z����bOI9���ș�5�5���ˡSY�2� d�Z	����e���T��wfb�t3�!˛&�Sϩ��v�ə�̴cS1�;����-aҗ��^���p�"�G�,9��L�m���X1���-=�Y��¥A@�bc	��Z��t.��r��0��ut V�Ŏ��W��ى�R�M��Kd�R(om17�c�V=�����6�9u4�U`
<�m �s�vG`is��^%ʵ�:V�cie�`� ���.�.���Eb�ܽR)�,bs��k0Mܻ*T�sk�753��$�h[im
b�Bu9QՑMCov�i,�������1��sj��z]�;�*��Vg4�1�:�YF��柒2i�)�F�ɶ�X��x��e�{�������H�L�9r�e]e5z����bU/وѨ<mj^b�f�*��C��G[�͠���@����ћ0qnym��ř��J���[OfEcn�],5kGr�v�h,�ʹzj]Rq��j�xP�8�2�,c*��Ռe�����aR�/Dœ�Q#�D꼶����{.CGd��MN��Q��&�S%G�[lK�`(�-���l�{�ydb�+(^����/(S��.P�kN�&�\��/ul�j)�L�)���ۮ�*v�1L8�'��#v����f�T��T֨t��aܽ�jM&�1�+�����9�MY�nԃd��j�囲�n]���a�j0��9t\�NG�6��L��?]衒�)sh1Oe�X�����)��� V�e�sR �K�%ah��R�֕��M��ͱ[�3�D6�̧���.�e��j>�0e�\N�t�0�
��b%	�X�5d�����ye;Z�)���E��ˣY�[�9J��n��%I�L�m��٠�z�ٳ(��<0m`��[���Nd���@��*8�d����e�/%0�yif[����rfouL� 2GyL�sYUp�P���ִ���ǭb�[�Z�ڵI��{vX(4���}}f��u�-j��8�f݌&(e�>)XX��k;���$�Oj�K�S���8o �1��Dp�~+���U��p3enc�sΒ���-�b�M�8FڏV��{5%@��WMb�PH�I�ڼ�m{z�K�O̗�bM�,�Bn��m�dVb��X����͙['��]�X�6��d¯�b�,m��L��t���ֱ� )E�ш��H�oMl:���^^\n�.R,�ukeml2�Ś�1J��C����"�;�'��6J�@�n���҈���MҩZ�KQ3f%M�R��T;XA5t����9@4(��a,�܅�Pݻ�����pm���P��a�u�ާ���`��[ر�3&Q��A���Ul��k��Ռ�dQaKd8�@$�C@��<�x^�Ƃ�ۢ���2+a(%-8e��f����H%�d-���X�T�ou�0\�H1[L:�e�(�8����I-�E���y��QOh�{Kwu�jI�0H٘(@#�®���椲 1ظ��ha�
tl=��^`�Gh�>(�)Fݚ�Q���X���CS�#�1K��ə�Z�W��f��6oM�N���),a���|��/����e�)���b��Z&�#��Z������;˅Pi-��d"V�Vܫ)-Zt%�1��/f��a�G";u�*�"��G��X5��Z,�A�@�
u2&"��ݫ�M�Y��ܬ��[K1�J�!�f��Y̱�o�0=דP�SUf�n�����ʐ�OE0.V������. 6�h��9Z��BG-�[Y���+v�r�Zbb	�&-u���2��TR8�8�l�5֭��f��C�ˉ�]��/l�[ˑ�%��|B*j��y��7èy�9ը�2Ro�WЙ�`�؆�h�5����}S�g4��&E3&c�X�.NÜeu3L����:���u�=�͘�5����j��T-/--��Q ��Z�q�R���x2��N�=����fb�d��k[9��%�� � D�ǐ
�;㽶��ѷ+$�T���b�1���4�C˶F5�z\"N����]��!�S���Р+h�Z�csH�<��+8��uw�E�Z�&+�j��R��\���B[_��涫?��?{�P�-�����,/
�����?�����jì�m��D&39A]t[���nt^IZlڮ6�*���s3Oh7Z��	۸��
�+v9
����w�)����]���+�7K�9��j�]Fq��`ŻPL�D�Y����̭<��Τm�[@�׺�{�Uu0���ܻ��J�|��݃3pº��m"-땙rvs��Ӕ�����_"ki+(�
n�m�Cs8^Iʶp��tzk�ZJ4ħ��ic��6^��f-����LĬ�y2�2^^�j�����9��M*:�u�K�X�8�*�ȫ+�\���zrX.[�]s��X�>���3ve��E��5e,�i�, ���-�G��T��(�J�n�y�(���ـLVv)��51lx��V�GI;�w�⭑�5���7+�⮏�A�q۬���n� ��E=TR�	bnNc����N/	����x����ȁ�N[)�p��,���Wbj�z�(GGft��)s**�C��;��#��]�f�'�1�]��g|������7Gt[W��M�ARa�G��2���1Ό�T���]�e�7�%̂�[�	bi��ٷN}..
�B�=�a%t��Hޅ���v�.�R������w�=��։о-j����0vڗ�w�S�쫬�"�"�v�WC]�w��KV\��[#:�����������e��u�F���IKDtAr�Q�שq��l��ڗb� �Y�F�+k�[�%�Ags���&q���-�w`�o��n�y��)ʘ�r��9]��ۼ�Dg�]c���t��y��V��u{d�|%��Vr�|�1㮙�p-���O������v�����̜i���V��G�f[���Ψ-If�C/�nK{��CV��~X�k� d���e�S�+j�S,�L����*|"��M��\]uV�R%b�"�Y����������)�D!R�Օn�c6)��sⷫ�F�N�wݼ�şk��t+��Ŕi�J+��t�]��V�u�;�2��1q�@���!u�(�z9txA�
{"��6�N�`��������d�ܮ�����*�\�z�d5������J��+j�2�fU�qt�y��J�kU��mY4D���\N]EIS]�g�De��dg��*��o��߶�˫W����� t��[.�XRPh��푫�im0%!�u����S&�Ȣg�n{D`�.�񇢊w�uг��u� ��L��]{�7i�x7��C6�	J��y�P�Ԭ�v��(��V�s�ᝑ;Et�����u�+���+er�0/�͇<��p�U�y�g<���Is�ɂp�����g�8h��9���b]��̝vdN��M��z�<R�T�A���Ε��X���c'ʙ�/%�dZ��f�\PՌc��TU���k���|�q��:m^k�	j�6u���F�;s�I�|v�E�6r�AJ:���}p>|���Fb� ��p�kÎ�juxŗ]�a��}xQ�n4>/kB��T�r �
�A-p��a�[�?�F��$M/���[pk���¯7u.�������Wy�|�߹K�q�'�y��L2���Տ�.�Ǧ,4��l�٪��Nu��*�Y]H��ʾ�*$ 4���a3-�T�Eo�.�h[�W6^q*4�8��7FuD�=Fpm�D��[�'TЮ�8�#9���!��ERs���>ɽ�����K]W�E/Rh��=h��Uy������W�&��U�����DR[)���m]1]F�f�,9�d�/y��D-U�������	B\���]���:�J���ҧ{��9`ȟ��(7���y�
�����%�]��9����6�j�{ˤ�CNW\�g.��("�cC(WG�ҟ>2���ZI1@OV���3���yMecՒ>�wR[ճ,qV�Z3�8;n;�ڼy�WA���@�˜!�K~5O��J�Z�t�8���)|>���R�&j�r唩QjZ]\	yʺv�i��Z�Z]]p�[��Fw�,+vث��2
��7:7���&'�yK>�ծ��=�3b�;8���:p����# d:X�K�JR?lc-�X���U�e��v�+�}��|��ů7����Fbv)�=����[�_Z��o�י���� tP�9�����aR�SE��c�p�Y�Iד�����fWC�nPn�Z��������=V���d�X���'L��[���:�Ң�t��ͺaG8�T;sS�5cyL���-��G�|�m��򖷻��Ӥ�w�@4�(�]t;�;��:.����4��c���S0��f�o+BH;wJښ+���u(
K�gj|�7�J�J �4EN�V]w[�t�q{��&��	��)"��f��е
B�j4`�)�'ON�Fos�����b�����2�Wx��B�u�c�m�1�����{$R:�w|�����lb�f��X%>u*�7,�c7�����&Vh�t�(v6��.��s�$�35<���:��� ��O�Ʃ�.���n"���W:�QӨF�+�����6�7�o��h�\��p!�=efY����K8���T/:�3Z�����.ߤAOޘ���,
Ku��jkz��{p3���9���5vs���N����
�=.�[��K�����A��,�]����ǆ6�I�����]"���3��9%����\�,��k�w]lT�V�'��׷A�Ř�f��8�h+% !�31 F �w�L�%]�ڶV�]k�f���n�k��$w�-�XƋ�Xl[��
�|�˭��(�e��.&�p}�g��'.���:��Eb�o������^�Ui�
�.�b������Z���O�;�E��15�ި�	+�Xs��0Y�S�3&�pv�㏨�g:(h��4��J�_���9��{���u�#�Zи	M��V�e�\����������Rl�p�а�9�ḛlE�*v��;�9��-wl-��f�ʱΟk,GI"D�K]�Η��o.jN���cOT|���S��EZX�����ɑ��j�(4��_�Z�6%{�(b�m:&��V۔R��Y�#5��k���TvBBzn91\���񝇂;�q��s9%{h����ТoD��	��ׂ�ИZ�%1r"��*>B=<�A�(L�B#��=���� s�23�Hh��|$E�u�}��3�a�OS��+h�h��`�XwfGZ��ـI�/�9V� <Y5�&ZVE�Y�)?u'�����},'�.!�5>Xg<��wVN�-.7D�`�-�K{�	�&�3e�y��4+�ա���e�k��!����7����Tn^+�i
)�Luq:ʢ3l���,��=�m�A: �ә��U�)3�F�V�>.�����6p9y�)*頟'����grd��9>��-�/�+�`Q�lA�qҎ��彵�N�y��m�Rw�bZ�H�"�λ�˲kz�D'R� 
4��SW�4��l+QvB�X��	��1ֳ��*qxet�m����p;x�gZ��r�]kp"�p����XY�e��U�xjU�I�.1e_ ����_`��䲮̂��=�:ϰ�'�ߑ�D�ӊ�G����u�{RF�g<\7u�4��s�v�8��}ԗ��ʷ|L`�B�x/3��f&�9#\�ve`:$�F��aWqP�.���@�����{h�� ,wcnP��@ݼ	X��\��T#:���l�Dr+��nD�\@��IK�z��KZ���u��Q�EZ+�fi�u���;;m��wE����y�Gw���Tuk�O���m]wSe}��A��OvʴMۦ�*�5����G��û�:�+�@����(F�nL�&G����ɍ$)p2���<���)�
˕.��N�l]�����k�f�ReI
w�OךEzC@���k�x!�}����7#���1���\����ţ�V�ͨ+�W����f�Gx�rVe3���,5ֱ�K��U(v��f==��[R��� >6�w��Epq�Һ�k��;I���A
c�dI�ˮ.�_eY;���)�yH�چ�9�;��-b���&�ȏc��cgN�,�v�ӑ���[v��O8�=ٕ`�ɊG�Zޤ�ؾaH.t�8s0K���[H4�_2��<J�\��ɕ��f^}+5Kڅ�F�݄����� lӕ�;H�v�43q^f3Q��<.Nj�S���̵ �k��Tn`����ژ֋�n+�Z��y�}y/k����di���,§��YV��L��&�vج�� ��`���:2��w&XƵ>�.�W0g%���x���įf��q���:N�.]Sj��Ӝ�dk�Y�Y�m�����h�}�+z��7�i�"q�ʍ�u|J�IJ�P�$e��z����ՎV7I][g�E#���]�u*�=;&f�}Ev��\[���KN\�@�꓎�y@KQ�iM%|��\l�P��t(!ϸ#�Θ3�('w!Q�ox�Bf��*O#��N�or�%`
��J�l��亸�9��С@`1�[�F�g�ؙjփRD�U�v٢�a�x�eIi���8��/�_ZSt�uwn]��\,�b�Ց%u�*@,-W��h�$g��<J�u8�iWm1J��2%j�j8so��D�.nq*sR�>x����J90�X�N`
��ǝ��tٔ՞� ʄ�7ݤ�Y�� f���#��[���QTV��� �̎�4bgh�vC)ܬs�ۤ%r�GT	=�6�}a�ۄ�-�5`�8�z�#��z�o�*��s]/uK�{@�z�U���],ѭ(b�e,�f�)��d%Xt�C� �]��lq�V�֓Ӡ��w!oS�<�6=�pn�${l�w�k{z��.�ףc/�&d[�,��M!n]��z��EɊN(��8U�*:C:�fɮ�/�<�)��}E�����u>޸��tX���F�4\,�֞UF`���+x`�έ׵5A8a����{�S�%7wk��4g-��iTÖ�ư*|Z�/A�s��\V��kwgft����o�0n��1G@e�Lzɒ���qZ:����	�ԑ�K "��Y��L"Q��@���%�I�PQ��vV^B���l/%۔�V1�^b�hy��ˬY���>c��f�(,]���s-[X��Yr�)�Mh��͢S.�2^=� �yR��zMwm���΁F��a|bx���C����	p\s�M�J4���fq������&�z���XN'Q�NU��F �0����؛a�׽z�+�PA%��.��MU�$�#��G��/�٣L�)�`��B���q'@W6��Nd%D�XM��|����3����Ko8�Tt��mr齣i˥�j�l-��,�O�Z�ÙFɛ��Wʔ�:d��>ǜ�P���Jc�u�ަ�
�=���о�� \A�]2Pݹ	�ݴ /�ޮ���%.S���s�3�*06բ\[�Ԋc�ZWˈ��nT�C��s�!����*�b�L�<��}�b��bt|��۵�5$@��R�vP����o�j��ҳ�]�>��gc�s�j��G3;�s2S�Ϟ�H���M�W*�56��oLJ=��mN3��(e�uŶ��u��z�Qn��v�.d�02�/V��`�vU��IykJ�ګ�l���wm��rJZ���+m
ڝ�7Dx��ȻT�r�frؖ�����+{\z��v�(KW���p(+$y֭s#�듻5�+��
�cS7]lzR��i�4�w:,h�E�ܥ����F���d�0sl+e����y�Z���u�bY��	��ք�5ו��䩘�[��}%C�T-�=��/L�3�X��Wm�ʃ��>*�mC0Ւ24*Rcr���Iv�A|�u�=+S�kU;��,NBr���*Tcͭe�8�j`���3�I8��ǌ��t�,�o�����y����6���J���/9��l��\�������ܼ[���єӂ�c%��*V��@���@_l/��1)i��]u(�h�]][7���\�1;$��8��1��~Q���v�'�]kohB#���-� ,�ju�u��b	n	Jw-<Լ<4]DB��D	�ʬu\����;+�r�sm|�;�1ce⩢M��q:�Lo�]�[Jv�s.�F^r�U��Ŝ��7�-œ�.���#�@���c�"-��j�[n�PS��k���Z���<B�E�I1��[��$���n�ΤF�Z���Tys*�q�l���3j��oK��AAx��}�+bv�G)sY����z��9��ۦ�;w�h����w�DqaP��˼��b��6��$l,���ky����]s)���Uu۷�Q���K���y�¶z��\o'c���2�eh0 �"�Z�ܮ�� ���b�U(��U�Gw�TnsK+%-W/����fLgFX�����c�^vɺ��'8��T�/u*P��/�nv���sƸ��q���a����H6!�r}�U�[���z��,rJ�T��JY��Q+\�ֽ�N;k�wQp���):vc�0�M����zW*�7}t��+#f�{E0�؝����)�J��J�v�&�똪,�|�u��j�}�2��o@ۮ[pgn�@�shV��[�t;P��t�VyD�4��¤�)C+��۹AZ�|jl(�ی���xcW���M�h�&�H늇n,=6ȜD��oE�K��r���"w'���jj�۶�Ī'P�����A÷Wb��`w.zi�����'$�5IW|@�n��e �gԂ���t�"R�U6��R`��v��7"ucT�u�%Dt�
L�$��*��B�P,��L����+]EQD�])!R���F��Ͼ�WS�=�}{7>���vL��9B��a��
�S��0|�4�I�*Pm�p
R����Ң��@�T�D�e�U E�{��������q��������%�w�����~q���������������������o��W�	����.ޝD�L��2�Pm�}����PnS��Ok^`�l��\6��%����Ӓ1Im���\�6���ܘ%j5�P���ql�fk�_n��s��-��6&�
j��M4*�93j�G�s镺4���ĥ��:�r�Z�Ø�[2�lӨ`��L�*d�8�Օb���b[��X}�`�.VSNp��OV�pvV�W��I0QT�ǵYJ�W7*ܩ2��(�;"������:�Oe�1�cf p7�jqS9P���-�P͍��,�U�O>wԞ� ��[`+VgA�^��j�V�K	�^ɜ�Ӯ��w��'�a�}��j��ʍ:����D޽�\���]�h-���T9qk�)�rѦ�h8�l���_�T��һ:fT��������d�
	-�H�\l�F�.�CYsbr�Ks����'���	gZz�}zc�l��^��a�\�5��Э˚�ٚ�!��BZzZr�[W�lX�θ7{Kw��Q��
=�e�*�JP��Q�ͪ9��ܹ�z�S[�In��si&Wdl����� �zm�M��f,�pM�͖OI}%ɔ��쎖v�n�xt'4b���S�ݔ�ގ�R#C�7a��4������]7t|�V�P�}�؀F�t��/�&�oIs&x�B�m�*��6h�.^��ͷ���7@e�	y��M�gJ[X}�XJY
~j:�1�s���"ْ�D��YK���z����H�Gx���!�WB��;��U��;Aj� N_�Ц���q��[;�@)Hu�4���m+9���D����X/�Xͨb�g�:�5{�5�gT�(����-D1т�to�K��.�����n�Iw�u���B�]N�R[�i��Neű����Wu��� r���#H�X��r�%��wYLg��I��]Ħ`�<����1亶��[�uq�݋h��\��p'ų��N�]R�B	����1Ђ<5�͓_ucG �Ũo�ղ�D�t���9�A�2�HE�rg�h��pZ��@�Ji�v�v=�"�-
�&�B��v.5���0�vg����J��a�]t�FU�c���.���K����gS�}+v�m�B3mr t��`�0\�6q¯+9f��a�َ��^̮*Ƹ������C��km�q����e��H�0�irgh`��V��{f�M��`i��t])���)ʷ�Wx�t==��� ��h��.�l�#*�^2��[�e,l8Xq0`��p⹛���9�'Ss�P�)=�2�a���Jb�c&$��On���o.�O��tL����{��Q�k|��Wc`�×֟msZީ]�C�.R��*�h��<-S��#j�ҮY���}h����N�W<���M�v����Q��'��c��me<��:�+�]a�\02gujb[��R��+4n��C����:��R��k�F���z��=[I;�A�--۟k����Ή��j�V`�G��K�|#�n�;��V:VwD�Ol��.Y��ի�dx3+Cw����$��)̵�y.��A�a�w*E+�rTI�y��R���.�J��pd
��0�9�2�t��ebMW
n��:�5����+Ô��\A.�s%F�����kI�3j�X�KsV
X�n;-13Ev2�k���yz5��J�@^���z����;z�PT_l��2��Y�\���i����i��vB�q=t�;!���>��W��=��3&��'�rL�.���\M�i��YԶ����ˊ�h���*UHy.�� �՝B��o�4�k�u3��ř���c��@�
`ۛ��%e�gr�t�Ll]���]k-ܐ@u�]%-b��NV>յS$}ӫ���u����9j��>w�������p��ʀ��J�営�)|���J�X�8c��w �4"x����A<�����5�[���a��RBW-�p:"��l�8��}�ܟGի# �W}�8K�f^��h1*x+���Zۺ�ͧ�!���ně�&m[Vہ ٩�X��$͘�7hn�﹵+45�1��}J����)��ҥ��y�+3J��'-��O:h�Vj
f�i�Ԏ���\���`��
��Yl��4V�u����OI��lz�v���,��I��t-I�K e�[;)�th*���gp��я�5��V�]�wШ�e\��kY�6���OL���'��u�E�+�0ɵcz��fӉ#Oֹڃ����k����@E���8��49j�հЯ���s��F��x��Uۼ�����	�ϱ���9��eKыR�d��wJ�n�<�7t���N[��oKq�U��[Uw��	�u�S�2�s�+U��b�%c�)��Y���j���M䬐�sZ5W:íVf�1��k{y<ގUK\��"�4j���7F죕̧S	0��E����-��9�I���c����>X�9��66:-�;R��y�]�	#��˒��'4qW���P0i��=�=7YW ø���Q��E�T�A�#(^���U8�.eE���5p���/*]���x[�CZy����e�k:��8p�x��2��ή}��׽z�]LR{Fn2:�M�V��p���O���L= ����\��rK�s6n��[�@�뻛]H|G�[�>�ڇ�F,4ZA��L��P��&U�ʚAo"U���[�Qm�b΁�+�6[��� >�a����`�$���G�造�ʝ�LMS��sY�� �)Q̼�Qu��`:����}�ˤ��޳o�[jt2���-O����`��R��gs�(�z���:ܕ5[I�qբq��;���5��\� ��*��c}¸���u��|�:w�V��M�bI(z��&��&<t���s�2�+�37�b/9���x�GT��:
NݼR)�R@��u�x���{�ʹ��hn�kUɠy)�\�g=�W}�!tI�SX����x��Ԓ���r֪�K)��Ul&���U�{&�9U�Q��o�Z�iTA��V��mj\�����v�n���X���Gh��j�I���K�B�މ�*�`�s{P̝��Ṅan��*mLv�PQ iU.�rYE��F�Bx`=���t��>Ax�ӄH� ��̡�[f�K6\��o�c�Y��WNPB�(�×�����]�_Cϟl֦_L%���P�k����NZ��"�蔫�`[��٦Ф�3�QR�Vn�旛6&@\L���u��>��8J�l.}����ad��uɺcwB*���u�����R��:���>�َ�:��IG\�:��\ǯ3�Q)�5�խ��u�X��Ӱ�8���[�c�o��[Q�c�\�P��I�����C{�s(NS%��v���	��Y{;����Q�wR�F��#Qv�Ɣv�v���3.S�;=���5j}�5E�����Pt��!��(�J%��X��V���7oR�GKx���e6/VT�t�զ�ɩ�G�� ��^�����i�9[�#]�����*'/V�7�p��X*)k)hc;��V�
U{V�ї�M���ȫ���k���Q+�Id�E;�	5f�5���e����"�;��Y
Q���n�w��b�m��W�Xá��Q8�G_j�9Iv�P	.N+��z����1$j�w����')�����SC��ܝ��[�]*0��7:�7KR�QoRN�8������nY�b�
��ޅa��x��L�U��s�0�h�+����9bv,CC֑A��خ{�'*��:hc���Z��EjX�=�nWZÓ���B�؆�S3��A��s]�Okt*\�@���)ۜ�q�]ؾ2�L0q�ܫ��yAK�J$K�8u�n��$��٩*�nT�t/;Ρ��4��M=�T'(�2�v�5����Ϭ�o{�4B�x��s-O�Jj5n�=�8s�J�[���@�.�3�&���$��r���ܫc�7�tV��wl:������le��+�t�V�f�n��smt���7�{���r &Kw�)<51���^x���.�ym�uaʾ%AV�x�%� ��ڮWƏV�X�@3n�A�6v�t/�e�'�'΋P��Ky��՚�F�)�h�\�C��ӷ/������}v�"eX�#�
�YW͠1�9����onM���n���X�7=DmI�M�oV�`ٜk���Ù:���13�"<�=9�T�N$�9��Gv#O.SC8��ɽY��:`]H��m�j�bn�!Ck-�ksr�tn
!�ڱ,���ᵔ����7��Mm�˻�I�QX�N��n�9W�-��e��77�u�h��Υ96�j]S��#�N�*���tU�'�ZEY��aL���rkX����,��
 ���{L�jfV�^�JW4 �L�E+`��*þ)�(�z�r7[|�{0(%[ژ&Q�x�,�['˖֥Pe�ёqd����r�ofu� R5�Qx�n��K�\��b2��L�)*i۹n�V<����ުt�*9��Q��VU�N)i����������:Y/��W���R*�qù�mD�inX׋b���y]q!K�]i��V��@�JƬ�\W)�\���x�v���nc�]�Z��U(�2��7v��Z{(�Ks�����c���tٛ+�+���,�b0��6����-�ͽ��͢�fn ��ʂ�]���g[IX�Ƅ��1�m�����%�4N�Q�Zj �(:�-m�������İ1z�h��Ƙ���d��t�Ģy5��d<[��2N�x�e���j)��WNuQ�z��7�o��;t.�1�s�c��^� ;�/�0�;v�vFZ
^%Yz֎&�vj�`t�{��]��|����,�L�mnLH��Q��:o��������9��f9@,Je�Z�f��U�h�$^�`�e�@q���z)K���|o�6:h ��V�_o�5�@2��^�Q-=%Եgꪂ�v6�8"9�/D�;�y�
�-����8�.����Sѹ�Z�%�(\����!�d˘�P���\�WNWo$���D�x���WLvcw��\n�yJ�mo(+o�kX��A3Z�1�D�-�}� \�|��o��VL���k���BL�li�z�͡`k��YH��	9�<0�_e>jȮ��ަ�z����^I�0���u[z�8�rU�mua�T���RWv��{��SP������OFk������s�� .��.j���B���k�6�YҨjT�,��	efF__k1ή�{쬸t�}[�q3�.�E�n4Hy�����N�{`�N�j�;1Y�yKL����P�j:Uo�;��"f�ꏳkd�[�=��b����&�
���wk����-��!A����iK�Qt�)�[��;�	۷�6�g�a�YE�/�M�V�1q�\y��-���Ү��|�R�	go�:�R��W�J� v�Di�ï�n�1�T�Yr^f�:����|sJr�sWm<̜���A�״�\�2c.w̑����M��(y��Z2����
�NkF�tjL��^<������2�]ܷ.�W�g3���[%̣�]���\ӫ�̭M˂���v�Ir�[�*�%�1��R]��wC2b��Ԧ���s4(�l����Y:�;���3Z8o%�h����W5ۭn$��ՙo��]/�m֦t�KQ�ٳL�@����нh�� ���G��eܝ���)I2m4R��J�4FR��U4u�TB�vk-i��4��hܬ�Y-Bܺk��6�Vrl�SzZg(�]Jn��z�x��F�M.J��Ёt7��`��4�w̟��v(r����������c���8QU����-�k-aP<��+r��\1��;�1��B��'*�r�u:���DWQ��� ��š�֖�����<o��Z��)v�W�:�8��b ��E��6eL�26�ŀi�mҊ�^+��D�NR�\�Q�f�����m�9"2�#r�)�Z�}D����0b�Ԋu�Ǖ��F�P���GN��OR[�����e:;d-���u΀@����[��<���ۅ֑hunS�N<p�%ʓ�^`���,�����D��h�&�N�K5�<+St��β�ߐ�I-�/�&�Z.w���-���n��A�]|�Y�Pw2��l�[,>�m�v�M�g�i{X�D<�Z�Bʚ:V�i�HY+L�پ@0hV����Y�Z5�&-�R���l���έ���X;ug7�*�Ь^��C��I��ۆz��L]��oNa�{;m0̚�1��ս�wkv�4�bR_%�n��c+%O`���:��hJm�fQdS��f��p��$߷���!d������)�M��c�e.}F>N��33D\b9;�ok�D���+)�>f�W�N{�F�}te�n��"��)���³$|�銹x�{	U�kp�e'dK0A�+� ]ɛi�mtVnU�h[�qM{a\8(�ΰfk4p�"(�Ex�%+�T��d�I	Ӛk�.
��1=���7�����C֫ˤgL���8��AeG�����Ҕ�X���V�\\��D�M�3�pM�5����Z�T���Ƙ�̱m��t�[��9;fIrZ;��N�z`8%��x�V�a��(b�n�5jj�pH�]�k��)gb�1�.b�^Hq�(�a2u�3��M6�a�\��s�RR�QV��n��j�f�宧\_�h�ҔWڭ�TUP�r�c�� I�e"��R#`�!
Xb��ʤ�&(TaLN�f�uF���}��7�J�Wx��Z��BY(m�C$iH3��:�<h�8�R�¤ ��!}ٵ��)�!>@#Yf�m����:L=dEEL6l*Os�4k$��������ӂ���iv�:MwQv� �8�͔��Z���_���`������������o�-�����[��῎��[�����￞��:����XG��ؕ��w�w��B1)�ș�Z%{�\w��f*˥��Y������[�k9h�0mٕ�¯��Z�f<����m�۲ug7%��aH!V�e��l�C�oXi���FV�n��kya��M�u�h�Y{���5�6�:i��Ǖz�����p;�UƮ����Z��fN��^���+Y��Vo��bV,���h:���\��$F��j[�0��ɻQ*2���:vԢ�f����j�mW+�]�l)Qu��E����y���X���a�<��aTYe5e��v��f`|_3r�U{EVp�6)��Mr.��q�8�V��(9���z)!S̝������(��;�Xt����`�z�����:�-Y����ݬ�r�!v�`2�B^GH�����N���J�j��Lur�(�;�z芘+s)cLIJ'0�=�bB���dsu�iw>�9�G�I��&��ъ�AD�7+�9��r�N��f�uh�����;)��]}E�c��|ziHf
�TdvPŏ�; Պ�ƸFY��n�f��>Y4VnE�rQ�%"����l��M���2����L�)"���j"�����6�lV6�w2�r;W��8�K�#\�n��8�q��J�\ȣ=![�fD�twU9�u�Zy"֒��Yw�j���/����tnwGN��0�>�ұ��I�E�{�;�"������v^z��'��{�z~�������ÐV��!.���=JK��Ď��9�8�ru�bR��s7\=P�]ݹ�yЈ��i��s^��'�0��UE2�������UI�Y8l����5��Qq(�:d'N
�$����
��9G�jA�������8�p�E%�Qr<�ݓ��p�98������Gt�(�t�g9����h�IZ��:Z��*�F_2��hr%ih(�����C/u�j��*N��{��B����C�y��^��ܐ�H�����Qd���Y�i�"���Si�<����U.�T'3Ȱ��B<�Hy�b�&pI�K��N��1�Ȏ�@�·[����t�'.:�R���R�g��w+��G(՟=�%kV:�PTERv�:Iں8P{���n��MJs��^x氳=�{�	�e2>t*EjfW*^��N�[I9s�NuJW�S���\�DUw���r��c���}�?�ɯ�5�+��]��Ӂ�9�[q���8�FТ֍�'J�R;<u����j=�z!�6�l6�h_��fH%=�|���{��hW� �w@��U����5]t����cޞ���Μ�zAz;پ58m�E�w����.s���ӻg��#:.�cu>x�f��.$�K�&��'=��I\��-�z��%�N{�PD���1P}��<"��^��H���&gr���y9��6KH��Y�'\��ij��E��18�>l,�$���]O��z[��\���Sk;���F�����蜼��7,��<[�>^����챮2v�4�n�tf�l��t� �~Y�S���t<Y>G�P�Q��kj�LI#�T�W��S�o\��I���OO|w[��� �]�]<�ޑ�y�T^�.�w�o��ǹj�Rr���#�����]yR{�.�ng��QjIO>��@r$�WkĤS�^�^�}�v��B.0�ū�Z~�/>*ҟ����lLJcqGp�\���ux�iuE�V�H��ݜ���Lpc0��W$`�/Į5�7���b�w�'U��[ެ�Y���N.ͳ���o3���"�W�v6��f�_v��+\�p��$����b����7����V�po���T����ķ�Z���_w}�����X��1y�����LE���:��^4)��d1�Em
���(��(����B�5<���x�3ފ�מ�(�R#�m�W�>\>��C�w��y�Q�)�z�H�eU? �$]S��h?y}�e�������D���;�[�/����e�M��E�8�&�ۼY�Ǹ����,'���?��9b�>�0��_Q�f�o�3��Z�+�:�U�nF�K��A�:���b+��"��:=��I��^}F�J�N�^��ϤO�ۗ�s��ˣ=�y�d�g���/,[R%�|�+�*^�^J��V�J�[Cm��������#�c��׫�vg�{v���C�K�0nU��f�& �������s��Jޥ�y�<�柽�~g��Rs��M���b�zP��Z�v��Np`��mf�*Z�"�p�/4{�����M�E��9ȅ���!q��⥣a3W˨�Bk�RR��QPU�Yh!Kf��^KnL#n�&fl=9M�
ۃe�g�	z�s�Z�pUɱ(:��:!t���v�b�7,\kY��C��3�����l)�y�u����瑰OSq�Lg�,i$��zj�cD��*�_���1^n�}��⮠5��+X6��6F�3sg����.�Npfw����Z~%8���(P�.�JX��7��g�n���>�!��������Cr>��uu�[�Ƅ����O�WEQ�9�v�-������OX��_G[�|��^�-wl��o���Ǖ��Lmu"��^������v���*]��z���^m'r��ӝ�a�6ϻ�"���$�!���z�:��]G����/5��+C��\��e����kޱN���7rH�9v �3���=6.zi�������jk�VOvߡn�u{צ!қ�xO}�h����?gS�'���pG�S���P���g���G�uu� ��n�}�bS����qϯ�^|׼�w�œ��@�|3O1Q�����Gk�����z#7w������q}��D�E�Y�h��B�KR;��}�^$7+����+(}��s�\�Շ�y �cŇԄ����8\�w�
#���W�5BN�JݴBb�k*�N��IAnj��҃��<��q�X������@�~�[�d�6������kc(���{~c���xs��}<�6��{�,o�O��{NL��}�;mwՐ6�Ҵ��H�T�[�b����є1q�!���:rm���.dx�U������^>���xH�f�=���>в��@��,�kwhn��`��@Y��o1�
NZ�����,ܙ��"_�ψ���Z�G�/�y�o�'i�g�v��^�^˽�9����쓟�Q�c�ş�g�U�y���Wt�PoT��řԴ�rv��s�=�x6���|ȥkhyg�*��g[Ȩ��yݾ�{�M~���%�����M��jm��k3���VT�ꂲk�m�����%�Ϋ�|������y3��/������89�.�.�.�6�z|Q^��/]����E�>��ג��n��/OI�1MnT|R�ܗD��D���Z�(��9b�B��z^���r���8�yի��ny."~C��>�F�^�ۘ�P��(^]N��b�a��J,�@՛eoX\��u�{�,���/�u4���K/V:M���+��g���pg=���A���F�k���gwf���i��c��-y[����)q��b�BaO�Ԥ��������+������ηt�������.���AuNpKڱ=�G���o;��9�¸b������r�m_ո���8���ʭN�V\��Ь�����w\��n��>�u�`�M٣��/����O(f��[������	ّq��^^L�97��%��v�_����i���B���5��Oh}^L_d����bvA�9@^�/4{$�ɹ�OB}��}،�;����U���y!�E��M�}�^��Xހx��v�%^�5���c�3%y(������ �)�Ut�	>��Z���n�w_�V���G}��r*��y|W%*{^T��[Sܯ7�,��8���ҍ>�?l��s���_���`��C���߽���J���9�����k���]G)x8O֤��Pw<�J{���\oRۃ7���0�S\]��\�����d�>k+#b(�rU�Ɛ\��C�Mu�**��V5�W�	O/�����-�3x�>�Z9`; ����8�n��0�t��F{��q�VZΒ���#ck"�4WXPS�&�79ֈsi[An�h�=��$6�{N�i'4��6t7E��d<���������}}^�m���2y�I����/py�`_��4l~�XR�N�x���pS;�Rƛˀ-;).�w����#������!�l���������p��R�R�X���G2������?O)�y���%�Q����ѓ��ޭ�HƏ)�N�;��>��̵�[�i#;�o�օ���R걗����C6 ���Q�����#�讎�	��L95�u�w;Zȁ"�����ܑ�4��B>�`R���q{Taj��s5�\���;ڟgs!t�A��ΐmOg���ʧa<x��It��+��N�T\��P�7}�y�v�Z��f�/�z�׸u��`{Q~�����Ƒ��YC��F�ꄪA���O���5�������j`u������ؘ�J�î�X��3�[�3��s��Z�4Õ�u0�-�z+5���sfҺN��o�rK��dk��La��=Χ8��&���/����Ú`�N���
�^Y��o3�	�#��v�P��9Hյåe\٘uK��SC�'�'�K�Y�/�zM�<�=�By��k|����aO<�i������Q���ݣyq8�b��ݓ���2��x�W��7\�:�^��~����ĝ&���o�{���{˽�ڽ�yE�H��[��@�b|��3Y,��}Ο(���P�q�1�ze	~�{<��{W�S��E�랦/��K�'kO���;�!Q�܊!�5�4�{[�c=�`���nE���ӭk�ݓ�`�
�?�ʳG���U
פ7��z�����'~�/�J9K�[W{ն7}��ۧ�U!�W~s~��;�k��5Ԟ��O+%�vg�{Ϥ�=V7�%����v�.�:�㚝���o�f��Wt�M��2m��a�n�?�XBzw9.蕋�/8<n�{�6z<:�Lm���הs�d�������}�
��9\���㗃J����[Oo��V�YG������in�cl�Q�Jz�oR�n��q7'u���|N�Nn�>�+*{�I��خu��f�������R�>gz;65+���KR�(S�T�]�"g�]fPgy��,s�4]��fGS������}b�>������n` �A�Q8{)�)�0�4�s�My���������h���FUuݣ�(C�dݬ�~��d��^�V}A�zs�]=�].�W�})�C�c��˯z�.�z��lu+3�����`5�/ݿ{�R���V�3xf�ϫ��h�m�"6̭�6'Fh?x0.��d��b���=R=L���4Mc`"����w|�#f�Ϗ�;�3K��h��g�{e��=�[�u	M�r�S<������)=�b��^9GI���-� �c��<y1�k~ۜ~t�YW��sۃ���|�uY�#��o<�OG�Y�w����%�^Hq�\W��NG�gw��^j��E^�gؼ����}�{�mw�i�����0ں\�py�>sgK_U�j�ڤ�}m��g)]+i?zS>���}�$KZ\6�jz�#/[�Fjd�כ�}�����C)��u��!}��??eg`��L��s�3Ϫ���)��)�<�G"�8����n��X3uX�^�����.��K3�n	�o��B=�a٬u�[,�. �V��Ư��"<�=�K%P=���@�����ea��ۓ�KV�9�J'*�9�?bK�� ����I�~.�d�{ه;0w�C%.���7���$k�^����zw��'��wW�h���*#��<�����U����G��N��W�-���7���^�>�9�Q�ӽ����z��S�.��W4ˏ�+��v�Y�_Qr��$�U�;7�nW�=�gR�'�x��ʥ���iW�ς��Z�o�ߓzT�GfU��{�v�9��R��h{()`�7k�]ymk�/7�=�{:P�M=ֻ�A�y��S�W��{��aGG�*��Ω;�Ȭ��$v`����{������G�di q����6x��_	2�||y�0�O^�Vã���5���f��q~�Op=>�@/���؝��<[��9�{ړ�rP�qz�ynQ�|�O_g�%U��W���߾��}��Z5oeߪֳjx�ޯyu���L��+m��S8�7w�>٪eF��Z90�n��[g;(�|�woȯEo�h�Ea\5�K����;��&v��?7�ʵ{��)b���\��!Ҁ۳���|��7���P�B��l��<���.�)ڴwz�]��9�2����U���4��- _8��7���=��M~5�OOO4owŦ�:F�0�	)t�}�'R���t����fy�&L]���B�����~�[�ޯ�y�I�r�;��y])�ב��
��k��O��K�wc�`��==�L����M[�F�����[a�ޢ�x��[{\�K��q�#OM���͡2-�o'���i�1�`����
�����Wr ��z�u���[�J+>�wO��r7�)���p�״2�o'�M?y߶L����)�E׆i�Y�6�1��z�[�/G�̣5�&����4�HL��Ln��D��t�b����u���q����]mj�:"A~�!zn�~t�������OÄϧ�YG�࿂�ʺ}:��rs�ټ��_���M��yp͌)w�m����W���/�{����}�o�����}������y����@����)�K;��T&��M�2�����9:��$���DJ�W=:a�+Y����>�*�^|i_��\[`'b����yW��|������úI��$�^�Q�ok]Jڶ����/�[�4���e�����B�rim�%Yn����e\�4��OK4�|X�;s�D���3�9L݂&�;���GR���&oW:%�[��a�/8]J�Qr�D\]=�]����hr��i��>vhYҔ{�̆�e6�uv�f���-��ň�674hT�η�RS��(�q�lTy6_G����1������.�ݱҠ,Y���#��نA��I��)n��kjV�.4�:@\�w,��������z�o��ݧgT{�ARz��Y^���"�XA'e����v����j��+�������IH��$e(��*I�V*n���4/V\�ƶV7
	p�GB��D�(�6�v�n�@���*Z�bʮƜG]K���"<�f�zO�QJr�|��XH_Rmv�'yX9/O.��ڟ6�BNv�S�Ck��y�}۔�hn��6��i�)���D;��U����qc���F��:n�1;c�ز�~���u��T��٤k^�79�RY�q���j�v�L.�o'�޼��	�ޅE���ձ�՛�\�}�j_m]�4�U��f�Xku�o;��z�Kz&
_<�y�B��t��.ԷXҐ�^�ʳE5��R�N_N�bfu>���.��W}�+:��BUdc�2��C�b<���nSXk" ��)�}�w����;.��e����>��d�h>���W��%R>��F���%�Ҁ�>w�S.`���q#�\*�3�D�Df�����t��&��v�%���d�k�z��ɧUv`�k��n�ӻ����Wz��#�*�%�r8�ܳ�:��jM|odr��r��net��>�-^�U��tf㎦T�#�8q�C���4	���ȏ=���,�	E���X��5hk"�-`PT�&ɩ�ʖ�6�����y�	����f�乕�u���%�V����,�$�^=���\p*K����Τ�u�5�Zt�����dl�R��b�L
"�W7��f���c[�Y��)�\����Y,L����D�L'�
�wS����Z��q�ىT��`�[Xy)�>��h��:��5�FK�w�jW5/�ݚ�.�S�p
�C4�h.ʛ��1���9�Gl<����U�l.|�ͭ�`Ȁ��>��s�M}����>/by�m�������<12�⎵�v��هk�0��k�du�Q����.e���&�ǃ5�h(�J�I���9Ke��0d�{�y���գ[��ZY���E��%/�8�G�r�l>W��vL��yM�ޭ�f�ft�bt��c8��.�Z j���wH֮�������w۸� �x��M�u��Pe���m!���<�D���={H,�A��{"u�9��­b��s�#�J��k���+�jL�jQ���[��R�����"#R�	�G������xN�f�z��k���9�z#��){�gOk�]���N���׃��L�����-'x���lrЎ�D{�{�}7��N�(���q���{�V*W��9�r��ru�J�xutw]�{���#����=p�2��Sq#�z���鋗����Gr����yЫZ*@��r��ED�9/[���\#vd�y��{�*��}<u{�'r<�qr�=�R!�x|���z;��9=�[��_!��;�������{�����У{�Q^����C��~�dNi*�ʞn�.^�G��GT��RK��[��i	z;�(��x��i�����t�>��bs�9�J(�[��̏�r=};���׎8T{��?I8�$�L����%�B�TO���0<�Pd�T1�^ϟ}\"I�K�"<=w9k�8�}ݽ蕕$>���)$	̯_O
*#�H	\��}!r���՜��i���_��S΀rV����Y�A��s�rJ�RMQ�P�f��(�_O�>�Ĺ2}/ܦE�43
i]#Հ��j�^�Tť���v��T�BVfJ��epu�����w���l������>X��\����R7�E���g��~� Z��k$&͌=7���5V�n��v��t��Z	���B��D�폆]�F�ܣ���%�`��Ӈ�7N�ޱs�I�i�h�]���U1�%�g Rj�1���N�ת>��UI�7y���|X�E�j,�P��'-m]��',�zeh72l��U	ޅS�0�������+���H�٬�d}�~���\���B\؋���C��:I��)�)���~m��+/P��>r�<�dDKxn�<�Ԃ��#(�
ظz�o�1�����ӭP���4ɻ [ Km��]��~�KV�G����u���z,W���>m�������p�1�y`��5��oE\���I��)��Js��}j͇eT��)�Q=Q�bAlwO���o֑OJ�J����n����|g�P�R��eQ�¢ӀNT/h��5��\?���6F��ɑ,t�EO�����`�#��0>X�+�<&��F�%r���� ����s� x�w,��B�\��������/*�� ���/��'ئ��=�8(��b�d^�h�L��d������׸*.��6�<�F)��k@�-Q�4��#�<�ˈo�uTWwC��V��s+��G�/��ܽ��v�=�J
g����ޭ���ۗ��hѭ�~��o����X)�R���fu؜lU���3���>�EƢ;�s����:�ul.�6�Uэ��}���6oQ�%�&G9�(���f�~��;�[O��ʔ�eeB`k�ǡ��0��>0�Ze�ͱ���Q�}"}��Ӏ%�L~��_�Eo���T���ݯ��r0��N����$ST	���R!E� v��:�$�'����X`ah�em��i0�dhOV�}�ڣ�^+�6��E�0��mU�OI����It���d{q���%��n94S�oj0-��uT���'�d��, ��y�/#�HZG�����潋��u@��b沼;Ax�w&9�h34_���X�؝�)ieOV������R���'�6��mN,���K61�ݡ����}�x%��z�W�-#d�B�mE��# ��D⒱W؀���|��P�`8��"�㜽��$h�L�atʚ����˯.�!gv֍��?{Ҋ�r���k�.��P��Jxi��P�|��ֶ�ZևT!hj�'�f�0�to@�85N$��<� G�-R����	��=�7���<Dv���/t����·:W=�tZ���U�w\��� ���-o�qG�4oj=�?(2*��;e�k����1_l P�-tuƶ�ٽ���P҇�=\���;Ւ����� �7B/��\4�J������Ƥ�����E�v�Q�$5�sy��Z}T�ف5��Ie}������᎗#0s1 ��ݧ��֨͊���yż�l��i�,^߲��حlgߔs�_Bu���P*���M��|zׇ[�[��+���Y�_����u���Zj�w̢;��ݟ�����ѡ��ZO@X\_0	��V����ϼT�����WOٻٛwX�e�@-̡��NTZ�WH3T����΃�UA�lo9��͙n�m������E�f*�mk�c�zm��8��Y��� ��DP���vwƸt˞��n�p%=�뺩q
����Oo_;Fl���#I�#R���U%��� q��ք���iB��5#�AtrH\|�F���s�2�8v|~X1F��LE{pr��,X�y����ϭE��(����ٕA.�"�Ǒɭ�<!���j���lT{�����qT������'�Z�����_^���t��`�6�&DWx{}���x�M!b~�h�	�o�5m�ƽQL�6K{�[^�Rb�j9�%bM4k�t�N��^�V".:��^Y��^�A:`�k6�o��³���du*���9�)��|1�|���p؋Y��8��J�}�1�~Y� #��z�捧,��"./T�<���rO�{���v�uf����$���޵����ύb�̷uó�9�:)ϣ�?n�S�5�ۧn�9B�O�e�30�d�Uؒ1����
�f�������֠��܊���}��T�C6�M_SJ��;���fA{a��d�%(��qu�T���Q;���1^�d��5�F�H�*�
%��2��R���~��}~���[��x�(����D��k��gP�T�ݾ�xcz}��E��`��gO]0����D�撤Mi1w��Ċ���B� P��Y�|e��,��Z�Zp�0"�_!4�S�R���5��Vfo=ί#~�1e3|
�^3�qԽi��b$���&M4>.'�a�	]
�&t��Սt�z)��+�ᗇOEvqd�D���>��f����}+�J�CH�&��ùK'1�}��k���2�����j�aR��2���+j�@	I��� �z��07yr[ݟc����h�<�NI��#��v�a�d\��ڢ�ifV0�QS�0*�\Pwƍ7.�S	�=Ѧ��h0N�<ۭ�E)�]A�:Iv/	��In�*�#�Գa�^8D����%����W��K�GE�c��0z�}҆�=嫜��ذ����_;=�bQP�*�ɣ���\�t6�:�Cl3��D'-@OCk�Ց,��{ �%�g��*�{������7�h�c��n��n�7U�Mm�k>ZvC��܎��'fp�k7.v�:SG;���}�Z���KK$"^��>��������Y�"��7f�|¶�}F��͒�v+^C��,�N����"ifp�f��|=o*Y��F;�kiA�GM��R���ct>�'��M�[}����0K:��X��������n��v�Tq�F�b�:V:�i����ݝ��Ϫ�aB�i ��#r5�o &,�y��b�0�hU�y���f�f�����{�z�����8�{��a�ٚ3�k
�9?k �ضCc}@6�d3�M��d%^��p�ǜ���ZQ�^�R1�����+�uS�u�E<��a��#OΒP�")��,��J_��nL����a'1Gv���R�R�.�����l����NnH�#cg�#W�Dz�E��X�h���:�1�2P�4��6E�4Z��}�S�M�Xۺ�����cH�0(F�{�z͋�ZE>5H�zp��v���r�Z���I�ܙ�я�H���Gn�>��w�t��e�J��4lX͓ka�V�uv��
�������aJ_��i�CŇ眦%���rE�_D�W�$�b�{�te��amx^*u�^�Jڶ��a��.�qd����*��
�Pd�]?ɂ���Ϲ�"�f��\� �Q'^�L�3Ư��M�o\���"�f>�`�r|W���1���LS��yeB�ٯ[m]l�M�Х$�*��KIȕ�Z�[�"��Ke*�&�(�����>��ޡ��&}kwb�)�VTpe�;��(����[��(�X�ו��$��d�����ٛ�Q��'3p������,����O6���S��p=ܔ�S��$���w���=�;�El}N����� ��^��8�X;4W��tR~�R)��Js��ٟFk�:�[��7��{��a�^C�)����nE=�:0�\�PűӸ����#UՓl5�Z
N�%d��9�&�Ğ�p���JE����5W+	��E�Qk����(����fs�K[֜�y7�n��ˑ���� �=�[�6~���Z�g�_�B0�:YhН+&e���B�z��Unx��3��A�l�J�hbH"��� /1H�͙��ʸ�"E\�5;T�s�*������T� p�=_/oli�:��
���F������5yM�I㇉����95���}�[qi�9H��<�m��`!=Z�����D�?G�U�el.�3fb;}m���b�
�T��?B\���Ƈ[:�n�`+�:Dj��|�s~�5o|)��-�[_1�>un�D�$M���0��L�]Kf�հ2�n�wp2F������-����m3�)百��d<�k�P�~�H�	^�LGPF��S��z~��w�{�����͆���^i�v:��uߝR#=�[�V2�va����Y4-�i�}�G/�dS7��R�|Q��5!%B�m�qsJ��@,,�?feX&�=}?`�壶�[S�K��;�;�P�u&���â�Y�Ƕ��Isu�tdu�fˠNz~  ��w�u�Ԍ��]���v���䴭~+��P��A��ʶ�� 8~9�Ղ=\����$�-�F>�{ޜ.�%�;�\K���;�`ozQ]�R��6�D<�Ϟ̋�NIN�>�x���6Ws��Q1��y�2�{����{o)�Z���xk���5�
oP�V*}����c^C�����ωx��O�R���tC�y.�-�[�q��M�n[Nt����J/"&�u�n��R��fB�_�Ѐ�	L�{�*���8����2簶)?_�m��nv��F'��k����	V�5�HXۨDp�4s$��񈤡o yi.E��t�ק>[<v��ʍCG=uk����ո�+��w��ڛ�?R���y�[Щ3��X�[ �D�\^`ّ/lw���K�v�:�E�2�c���ܬ��jo"+��yHMц��&t�lM[֬q��ݦ���ޗd��K�ta�-l���=���]@�Ò;��|%�X���� &�,�]���93O_+nB`I�y�t�c��pn�����E��<sYL���H��5(o48����j|�/�D��<6��s�ɲ�h����XE��|��t���ʛ�@�߻^��n�b�e�{�-�'J�Q��t|嚸�QX|��e96�i��W�>�KV��gC���%eY��VJ�/�GcJ��GU������k�C:�>�����;�v�?f��eLB}j��iub���8��J�K6�=Y��a),6����vzuRĝY�(�/.�7���%�0f�9��zN{��{+����ꡖ��d%U��+��d��y��<.�ݵ}�fN��tW)��V��-a3m0����\�&4:�st�jKtճ9�=x(Ϝty�FWf�j~3N�h�cިh�k���D#��s�����`�١B��c$����ąpY���+5|<MoL񕾂�?���ml���c`EΏ1�`���������B����v8��`���@��M�iͳ���}t�U��T�fl9W��vY�b��m���0�{��*3��\�f>��:���j��0"���>Fgw)�lϻ)��r�_�����@^�&f�pG>i��.UM��D&�jAmѺ�	�[uQ���r����Ս~r�G=;�K�����(�@�����U���޿��2muqd��'-,3�8�����w^���fX����5ʒ�R�R���|c�W��o%��=9+,̻N�.M�גþ�X ����n\ɵ���VS��kU�I�!<պ+l0ν�U���4j�k�JZړ�7�v��,�WSz���'��[���蔼�]��ƚ�t��;]�|wh�K��{Pk�p�-�G���U}_a�Ğ�4ͬdW(��$�,�UL���m����T\˭�Vu����e�[����
�$�)��Rד�]�CN�Hy&�{~�N�XK���M7HW'@����z.&�a_Y����2ō�S��X}�y��<f8>n���ay�e�������b|9�:���E�+.3w2.���`��้�?�o�������}rޯa9B(���r_V��U�^3v�Uro:�+<�N{1����
��΍�'�m��[hl�xD��	�7�Z����N������ʶ�UE����޷A��u�B7?k�@LX,,�
<����rl���w#�sη����֧u,��4S��,qd��p#U�C4�#�5�p��Y��`(���YSSF*c&�j�}��z�C�>������ނgٌ�,��Mzxܴ9j����6M�J��|w���ỗ^�l��5�G�����Z�R4�33�7�b�K5,;#+�A���ރGy�Aڗ���3���tdΣ1�2m�zY��mF��+y�"kc��Q/`�� ����0'��ܡ�(1�����*/��z�1���g1�q��;�P�wQv�<s��^Ձ��}��I&����<���f��M�Н���z���jxR��{X��mŁ��v"�-�.�.�j���ܾ�h��(A���������8���V%c[���M�����?a`=��U��~.�m������e�nl���9�;�-Mk��5�ǻ��	�4��<`(���F)J�S�E�TĘp�К�uPl	�[��1Zd9��#��Q�����Җ/�mz\�e��E,�r��"g�>��?��1�T�����p�U�å�Wn3ʆ-���b��ڦ�	7����t�5�eс����I̔�����ӷ4�CTB�v���보����yN���ͧ9�%�~S��>_�ѨǬ8}�^�y0/��WΣ����/�ѫ���{6p�ϋ�eW¢��	�T/r����b�1�ugZhTÙW9/Kc�u�x���`�'��{�P��_%e���r�=��֌��{�R�X��Z�
i�P�A���#���ؼay!��Z��h8_���=�,��=�>������p��eV����_Vۗn�Oٽ~�bH"̅�dBy�D(�����➠��A5j��2�2�ӒT�k}Ra��О���\5}c��R=��F�[ ��a�=�{}~�o������~�W�x�x���w���o�C7����T�����x�ѻ������E��ؑ��1;��xj��y����ѵ��q���4$'uF�n�n�����V�<p����{��î��7��O[83i)0.�U#�)ɌtQB��Ǭ�qܓB���l�{g;�6���ǰe��b�F��V2�\��;�8���-�VS��&Z���I<��Sɗ�k��B��bĨhP�0���Œd��-��9�4Zu�2wŽ\�v�+.3��q�v/�g%ٔ����`D���/k��h^�
�%r��;8�te���ˡ:�Q�"D^H�УX��Τy���������I���<%e+{��i ��N�Mv�T$�9M>ki��n=8�O�~�����c��_m���e\����ҽbl/UӨ8=g �v*�85W>�"T�˘�wی���s�#zQЦ[��6^N�Eaa7�n�;%�i��G���L�e)�*SN.ȓA<�XRF�Ɋ�$v��unl�Nҭ)L�Q-k��M��Dru�a7�ڕ���T��9��z.C���>����:[��o���j�T9�%氛P����C2��`��Q�c���(S8o����7�\�@�f�|�]��L(N���>H+=Eh%�}�Q˗[HF���{)�z3�6��O�k����;�Ti�Ld\���U���!�
	�j3��4�����0��&Z�Y�Y�.L<~33
�iѺ��::�}.APnY�V�y��і�ӫ��\K�2rhu�-�'^m��el��s]��6��U��7X�N�C�:��u2�nƁ���N���@ײ���N�4�ÅV7���ِ-�ݤ�Vr�|>\��t�S~�Rhr텅Kr%ʰ)��f�s�}����!R8����Y���2��@q��B���o4�����,��Xh�X�=3-o�Q�$�Yn��Y1t�2�rwӕw)�r�����2;�D��i��m)KP�WW�su1:���6�s�7Èl�	�#�Q&I��}�I�ᑹܗ<��Ib=�l��W�B^P2��f�w�u2�c��
�׀:��4Z��r�MX���
,�Om`��C/yWLLr�\.+ƱgMf����+�$�+N�e-+��wm����A�ţr�oVk��vQ����[Cv��e-�27�n�ڄ�S5���B��̬�ڴr��X��ۼ�A�g�o!�K���{�rQ�)Ɔ/E'�c�X���,.���x��2���XV�w7^:C}4]���1��	��P�;%�]�&�^����<+n���(#S��iL��wd���nuM�KZ�]�3$�Q�Ab�G��sפ	���]J6+vmvM�+%��%S&b����;�W�1���vo���l���p��AxUt�.��e�\��I)}nx,9v��M��rG��|���S$P���W �e�V�u�3c�C �b�%��gK��\�1
�Ʌ��`P��r�͏M��S[6���,��[�t��۷�����ʴr�e��A�m����;t�QӠ����C$q�vP �&�*4�� �R��w���FP��9"z��}��E}\r��P�S�AEG꺝V��'׎�-���=Cֺ,8N���Veo��NQ�7g�#�H/�RB�]'2��	QDքM�E^j�E��ekԉ�.r��{��VɑD㋷�!(���Þc�@�4H�D9A�Q�(�� D{�dDp�W>��eU�Tz��Z�H8U
2Q�""��:D�QRy�	�3"��*�WT�*�,re%�H*T�HFl"A���]2�rCe�&r:j%r9TVhF�D^hn�E)ev�Y*Dg��B�L���0���t�wv�#��%̺�Dy��w �9r�ΐ�ʩP���
HH�+�Q\�*H�!�wm
�̮��"T���y�*
tA"�e�G!�DQ"��D�f�^F&l�^yϼvN'*�=vES�2��G9h��QUR�G�2��IVH�.�uu
t�"ݤh�7�<��ad���E�I"�$##�r4��Q��*РŰ�b*����"�}S9��09Zsb˧�k^޻j�V���a�Z��P�'���d}m�xM��� tDp,P�Uߜ~�������4" �����/8�c�=kɞ4.�I�����-l��FZ��5����K3������0M��녙<��o
���[(�ek��O(�#6GX�:��s�"؅�"6�UU�e�cA��Jƪ��{�lg����P�H4ySE?b���4L�X�2=�{U�`���:�\H�s���Ȼ�Du\��=��&��ޔI���BW��6�\�-��=Ht�d[�1�۵�ʣ$J�i�Ye-�q�윭��%�T�\3a ��q����R(J�Bb-@�v�dx??�K�76��ͺ�O3Ltk��Ԃ�5&n�pBF��mOitL�J*;c�t�6��yח�"�a;�&�n`���#��u/\�ڽwMᚖ��A�9Fm�k��k���K�~���W��}�2B�k׍��b��}�a���N�^�Tz���+^�t ��t�~�-�;\�S6Lr�����T��6dm	��Z=�Q�zW�8Jyo%`U�9�̯��5�<�2�eo�9pWD��z��)���e���vӰ�y˫�ޏi��>{���-�5�V��-}2h��K���&���^%�v�w�$��_!WATL�]8��/���~Â�ʥZ��>�д%����֊R.z���+���û�+�O�|,(�/nlEj����7��7�-�Ƹ��R��:���%/vR��;z�q.�*+h�呪�a9g]7Fp�������=��Y�Gw�����^�H^d�����F��r1��SK��/�B\��� �׀��R����O�g��wX��d�-T�����ǟy)� w��/aϛ��a�)M�G�b�{p85�H,-���<�֜�u��4��}ٯ!MJb�vS���c~�+T'�҅Nq_j&,��>7�4-�[w�}�Bvva�9�E(�*���k�C׺p� �%��3�%l=����殭���r6�=��v�\��Y�!�X@��'g��=ٜhVqT��n�����r^�o�Q�.�_��x���T�=.(����|�7�����	as�S�Vܹ=a�ky�|IX7iۭ��zUyV,��]�ʍO���}�[⽱+5��@N��PU�l|Bϲ\���M�l§�#�[{f7l�C�ͧ���=�ZV)��cI��`��L.�"��P�TT��ӖV��P�'���9m���$:�����S���Ƃ�AK���;��"��,��Jj����4����՝���� ��}��[6�U?���.���܌T��f����	4�b��,@����z�,�{qWH(�ͯ�'�j�.����Ȼ�/�J�3h�(���n@�wc�7h��I��5��uK��J
������węo���tg��upPwS+^�ERg)�'TC�|7����`J�@���8�kS�],���P�fԚ�d��6�&~��$��c��b�y~�"[��	�>v�1/�O�.�]�d��Wu�r�j>�1��>��0���)�+�ֱ��?|�d��J"1}��W��{� Bfzf��)����%6�#R�SUn6`j��d�y��� �Y��ᕴj�T�e}��Q�||X^��D<
}�k���������v���o/�J���c�/�7����Ww������%#���}fx�U��՗��ܚ{�s�m����g+�s�e�ULy�j�m��X������1Z����<��V�մu�>6'b���^�>��v��ҩ�9�N�XJ��w%V�rG�����ӝ�~gۤ�Bkʔ�c0NO	Q�d#�D`zri�=��=�E��iQO����X] swA����dbS˦m����g��,Z*�9A��yY�me}�c+���n��&�*���oЇ)g����:�wr+��R���;�:8g�X�lP���Cf0�1	��!�mIjj�5gm��3U3ѫ�z�"��kP�o5Y������e�t5�o
#�*j������]��)�V,�
�U9��/%�;+<n�ج�#r�9/�ov}r��~�c����>�����I�T
����xk������d��*��^�Kx�׳��vi�j漝�I��2_p�K\�V��k: %��@�*����u"�����:�������(���%���-���J��y*-�F���Ԅ�0�v�a��j��Aðb�6� �I5l���>�՝]��SJqc�3�W�O"�Uj����l8M�t#k_����.��C�J���򈽔�(fE,#�3���Z�c�:Tz�7���nk�w��4Hf�*�O���m	v�M�ɾ��1�#��F�Bd�����Q��/y���[l{�M������*�^(�*���vr��v.�P��G��|�.��qd�~%~����_~1Ń�~��7p��?mE�]����mKԣ��j��#ǀ��@���S�)J���B眦%��ۼK�n�Ӯc]'=,��/q�O	G3Ԯi��մ�'[n>�){T��R;�M�����BL��iv�"�P�^�`m�oB�k�t ɩdK&��+�۱l�Ux-�w��pܢ*S/��k��U��b�5xDN�5�@%��_?b{JE�]���s�<t	5A)�p,�WbBt�	׮̝��Yp%Ԛ�޶��K��)w��~��F�S�zla1�v�u�e��:���`�7��*�T�֛W�eJ�}c_o+.8Ө*���O��	���uu,'�nXp�|]@�O�-�qքW���ԅe
�GO��U%��H׍�;��knAZz���.��`�i�%�-R��7�S���3�w�4�O��[.�-�!���� ����*���;H�T�	�ι4�5#�!ҟ���2
tD=�@z�+��Q��dIF.���j���C�}Ցk{�eK����Ek��h�0u�xOD�F��OźCX+�P���&ɋ��lSNX���˴�k�vJ��e��Wq_^���wmHօ��dY=lg�w�a�]NWr.�/�B�}�*D��ٽB����r�4����Z�=�{���$��vv���@�ʲzqk"�y�K�~/b���t�kq�/[0^�}�hOB�Ϟщ��a���k_/j��Lhw��e�>W���� |t̸�1X��GOz��.;B2)�^�S1�,Y����2f���=����]�"I�*�#*�� @]Kf�ձ�}A�s'�*�굲�oiT�|�uƑr26|��	j�(I����U��ߤ:b��,�NF6n"m)�s�b���޻֩�����'%zT�T7a������r�P���Z5�7�ϴPy�Lv;���w*��O�$e��\����(f��iN�tLwzQ]�R꬏��ԥ������x�W�m���5lg�Z,�q��]ayY�����ď���p���4�+.�c�՞��3*�sw�,���"y�Qz:-�Л�ٺ��Q>�.�y9��w]�5&�.��W�k�T=�n����U.�7a������f����{�x,<�<��ȋ�LY��������;�͢��P��~?�fs���%ݱ���5�x�J5W
�mjޏ���K܆k��֫..��mAS�Jױ�2���I��[B����>�&����sԲֻ�K����M55��r'�E	\��ZQ��yEC����>�1��F��AK�d̅�gM���]�ZnEb��{���Ѿ��~b��"pB<���:Ŏsz����v��y8���W?aS�M��ץ��6��+e�c븦�db�_�8P���2����C�p��sfBC/�3O��I{fRu��S~ħ�_��/��E�[�����ʿG��]�2���v���B�k����G��a^&�1O��Idpy�y��R��B�-(W��{\LÚً��"c��W_�q���ЙS瘷��%�'�4��q�Ju��bW��06%!}d��٠Y�<Lr���ԭ��E���L7k�>巷>�ƅqR��qިOR�Rr�yU�jb�Gzo
�u�1u��j�_&,2��X\�����	rzFN���;�oB�0�f&�^m� mۯ��Δ�ܹ����o�-+xq����Gү܍l�`r!���%�f�]$�>;��yT���d!FA���%P�����T�P-�B��9oS�r����w�_�v�(co`�1�v��)�_}��7���{���gRHU�F!��Q�^�zzfM���i ��LG5�d�#־6]n�i�]N�v�!���	E��Z�����������+�a��9練 w�z�4m5��y^&bj�Il�jɾ}�;yL��lt�m�픋�Vd~��YCS�N�N�G��]�Ϯos�P��d���<Z����Z�E��I��ⴍ,omX;��<p��C+z<Aʫ��B����-Z�uaVr�d���敪����|��&%�i���������R7�~��R*��z�uKy�9F���i �^�Q�Ѯ��PV���"��_І�1}�����3_��s;��ξ9P^�-ڤQ��w�&����]�mP�dy�`�|`y�MFAS\���ş+�X몣�ߞ��l��e�e�ҫ�<e��[4ˬb�?\��U����׍%ح*�L�����1�bw|�^,���z�Ҟ��p>�0;<&�	�2˟���՗6�
�Ɂx�)�)��G].���f���_7��.e��z��G����:��z�T�ۘ��͉\�'T���d~a���ڡ�[2�P�^%k;Ҧ�;,1H��b�fˡ��7�RQ3B�K�K�3���l�0��<E:W+U�d��6���f�eY�����%Z�����jI��k4�;�N�K��O>�A�������|{�. �CY�gY�-���,l�8��1v�n;`_s| ���M� ���7k�;�By�k��-�í�l�����G��y3{�82�s�Qc�하Pƻ�S��p��6Җ�k����;s���l6�Y����N�GLG����<�g��}�j���lͮ��+v#ϊL��E��o����I�b�=hk+���~���˜��]�x�����p�2��j�Ǿ��d�)�s^�k���/$oP&���f@P<Ԣȗ��d��Ws�z�`�vB�e�4�|M뽟�t�aO�#�6g4�#����ض	����qO�~�"���O�$5ʹ{�w�Ǔ+~e�m~*W�|�;ޙE�7��-i^����I��uw~�cO�pl�op�H�8`T�^��ω�
���O0-aDbw�˨o���14Ǎe^ɩ�P���ѫ���Y��{�ʡ��0�:�����Mm���F/6�d;u�.Kk�Rn��,���C[\�0O��ˇ��?I�#%f>	3PW�3;��2"^1�'���Na��z�b�ɋ��o4�:���g���+����aF�R��C��{Y��-�@��=����eR�ʵ�B�<Sw��w���QV�<4T��bk95�Ѫ|�u��1���,T���C�k<��LE����y�9>��5�af*"�E��P}K�6dXP{�w+�u��;���*��6�,���b�k�赈�;R�d�f����a��"�]�D7��x|�x@m/l�>����%��G\��X��gS�xM/��D��DEs�o%�TUH�v}cf����Z�p��X��#$S]	���sRj�Z�΃&+"Y6��-�ⶵ��M�ϲ�_hWޙf�\�6UYXx�����u�ǡ"�ʿ��ξ�\���oyO.�]�yeg@�U��zY�obuvb�g�琺����_���^3Ѝռ�s��q��U.~���ɵ�E<osu��6������E���FS�c	��>������	Ϡ
�(�ޡkyW����6ȋ�ègPQn�l�v���YCl�Һ�y�1��/=�,CKa�6�	�Oܙ���ۧ�q�<��&�^��P�$�L��P�cq���6�nE�U�f\8X��q���
̬���R'�Ga�MW�L=�M)�0Yg����V�$n/(���q=��X�x��,4P+�KXG�э}
1v�{n/�����|U��c��е���3\b+�Y���:�Y�KL��|���G-*J�ZYZ��S�23dg�݋�/��m�e��əEϪ�\�fX�/-�o2{k�������E�V�gZ��Ժ�d�j9Sv2:`����3N�S{k��GIflʛ飭C1P��	�1�y�waGCV�3kyu��:p���Z<M�m�h8�����Q�Kg1u�&1�6t��ˮ��,ൌ�åq��W�U �x{�Sv��}�B6�'�����\��D-"i��0��L��m/���倳D���h��E.V�����뼸V�$�i�딯��DEm�a��S��y��بO�f,�̛;�L�Ԇ�^��T����({*]�7\�4���S������kX}�d<"��UaUb��l��ã|���`�v*�37ox�ǉ��;K�`�J+��]C�T^CQ�*6e6�f�3���EԙE�^�	5vP5w~�G��8���j�A���)$�%t���5���1mETF⎉!�<"Z�R����~�1^�N�IH���_\�*���C�)��ȣ�:A��b��U���7�P�W���l�3YPڌ���F�����	L��Q�]�p�+�ǩr�E�6k/��ؾ�\�oǢ��nH���B|�/ȉ���%����T�x�"ܳGo2m�����D]�B��|"��:�I�Q��je���㠷v��啲�֐�K�?�z'Zod�F<k��F�:
�eY�m�����/a�u`1���k��S�>�9ct��Dl?3���?�����z���_���>^>?������Gm>����^��%�ʀi�����ښ�t����-��)��R{A������x'f��Fs��j��c�~��S�M:�@4�x�|ZUy�:��Q��v�6/2�N�Ɔ��W�J����td��i��ڰ���*���!����R{����|gk(-ʲ�eu5&f|���G~�k]�T>�&������2V{O9ld٘b��qC�ɔ�v���*a�	d2C�0K��&��[<m�O.��5��	NJ)#ZtH�}e�N+T��<U7f���s�ul�"b�V�X��v	{c�kdݭ����g+��-+����b�R�@6�m_�V������P�a��p]��.�t��D05+S>0���s�B�WWN��Z]H�X�t�1e)(o/�К7�av�����)]�</y��Ā�yVq��&�AKu�V���l!.	��}����|Vo��m��[#h$��Kb�6��p맾*�z���/��&����Bf��ܭ�+����4nV�(wH$qڧ�V9*y�|�B�1�PXt��T�B-����ܓ�9�<�v
X)�63���5�F�$��z��u��*�#��wwz�M�|��m��l`���Z�Q�µ�to;HeE�p�'J��;;jJ�|*��.���^�"�w�^K<8�s+8�L�5�6��:�2���6U�1>2���u�i.�.��β�zA�KM,����5u���S|�Q��0�귮��OM��*�ǗkFmˬL�M�mՈ�Mu��][5�1�6�ճ8�C����cɞ��>z�v�3�sN&�X(��S��m��t��k�q'#�p[��I�7%�w�"YW�*}B�M�3 ��z,�._t�W�]]����:4�A�n�9*��
H�Xǹ�a�_�x]�Fا�`B;|P��ԭ:p�vf�\iS��p
q��ŝ\(���Z#k�E�l-(�u۰4fa��cw����L4u�7e�kI0�ݞ���M��}�Ν�t�s��יr�ּ�N�X�D�{�p���wr���](]����wD�:�J�H�[vVӧSo6Zμ�8����%�0�s|�=����70XX�Dv�qn-�0+�p���KO��+w�%�+��5������ɀ�h�j�0�)b��L��-9ly��ֵC�l�ޗF��Z��sD��aR9VǱ՚�YOYc��24L��-�n���)'���lvC�����w�b��MqI�=��&F':�z�������dD�s6��[j���h���k[}6l^�
綈)R��yq:�]0�Vu����/iY�=L�z�Lr�,�a�\�b��:��tr&�m���նYI��;kk�/�M��-���̃(�M���P�N,zE��r"�}5ҵk�ΙI�GX���B��wX�4J<�Y�7��]P�L2����?jL�� ��0�f��=��rH�Re�HQ �<t������ֽ��>�9Ȋ(� �A(�-�.帝�G��$+$�E�P��P<�s�U*""z��Q�h��u�B���]$��tp�ˑ�T��PDE�'�q�j��Tt���Tu�QތB.	$�A���,��9U2$��΅,��#7tu9&TQ��D��Q9��
e�YhQrֲ�D�(,�D�E�qH���+̹J��".)�I�(@����ݬ�i�,�E��ʼ���.��� �"ͤZe,�ΧT�J�u=f��i�A�Y8z��YVA�9Jh�*���*���EꅩT��b.�&J;�K�'�Ϊa\��+�͹f$$��RBW.F��"����	B?>$2�	=����q5gr>�{˴�]�U�<�O���_1s�0�F��,���q����F����o8+��0��K�����������{��VÇt���ݍ�|m��_��ϖ�=�^C��L,��=�� ����� �Z��GU�5�7�O�����ӗG�����R���}.4��kU��\�*��чiO0��y�F���D�=Vx��J�U��ۡ��Ԥ�<+YAQ��&�D>尾��l����ޞhlUS_%keov݌z��G:�Y�g�ti:όY����'+%��y�f59�QL��0�H�V��oq��ۅye��O֐�x��5�+�v˥԰���2n�[��՞D��\���'a�&�K-l���ޣ5+Z�5]�ĝm��`�k���_��}z5RY�CGk�`��Y�轊�pu{������LU�O+"A��.�l�66��({M|�P�c�4��}.�m�Cאc�Y�/X��>|�4���]�9]j��+Z6����[��oA��h�:fX�zF�3�Qh呲l�'�cq@�Z��=c���0���3Z�c�2e��^�cΤ�a�Nس�U���xh�,��.`EH̚H(�w҈Ƒ���NA[��C��,�.����<Nx-B�Bz���6T��������j�h����g����p�.��P0<H�;��>��Zǎ�e��Z�^�b��N�J5l�NR	�ޭ��㑉v/ik�z���������\�]�d�y+zl)�C?������hZ���ڃ��_}����� ON��,�\�߅�'�*ʠ[�X~U}F ��������񀳣ơ�S=��Q���]��x�^po^š����i�鶯wd�~[4˯ث[�@���uܦ���Iv)J�Jy��q�Kٹ�#+�_�Y�@������`�m���tĖ��ˊ�e��Vz����kXP?T1.�[p�u�Z�-�*��No9�	SG+�l�09�=n句�&C��*���9�:aA'�M�IU�J�eU&daY��<���#sr���:cƚ�C�`��Z6j0>9Hq������G�l��+���q<Ed��T��>B�}d3T�6�b�=,b* V�����k����u�[6���j�o<����U��n5o&��B�*�G���кb�;3�Ո�hP�����!����]Y>ն^�/��aT���jYaE���FL) �-k�kP&�@��z�e{=���V^�S�:m��[%嵳ѽ4�/yQNtt9K+��!�j[%ؿ��X71�8eH/K�>���{�yA�ڙ8�U�S��&F���O�L�q�����F���5kƙR��Nn�@��a�@��7Bu�Ȫ�Ֆ����
�,;�/U�]�Ur��g�Ͼ��5�dmQ�}�dq�4E��z33,��ES4�T9�G��{}�1}6�!]{G��&yԌ\�����[�g�V)�m�����Py��O��v����=�5��|#��r������*A��k�Gp��U3-��x ?0���Paոb��������`G�l������b@�εH�ilfgxo��g�y�#Q��b�Dx�>[��p��"f��~��1$oo�ɶ>,����"��P�þ��4p�`�:ɻb�wm�]�贱����6Ś�f���A-�\�%dI������yLK��}~Ύ�L���]�y���{TE2�@�l�~P�d��c���ar��R�(;^Ȩ8a��	�A����F���K	��M�Mc��k�j��Q�f���kƭ�a���#-��߈^���Wr|w��x�uR:�l�K[��njGW�����t4���M���n���͝���k�0�*�R�>�&d�������� 6��F���Nl�"禎>{�S�{lQ~z�T9�7���}J#� g���x��QD���9z�D[IP������O0�{�J���/r0�x�ƃr�=�f���j#n�J,�'�ۊa�|M̚���g�"��<��	B��������"���xt�N�vvAjT��@EE��/��P%����Ut��H�w��>e�^�>�]f�*?N��x��­;Dڣu�*_ۥaރ��ʸIo��[�<�|�p�
u0�xl�v�d�K�7�sV'm<����`봻 ��������K�;q�u��\!3�:�}��5n�Wx�W$e��nkQ=QPo�ۿ?�����^��_���D�l��c�{���oxM��b脜47��J� UyB0=y����;>�̠�9��<~l����&;�}a�e��L�;Cu�pϼ��L"���
�6�ؤSU�@��iN�����ZN��=�9۰_W��ܺ��P:�F�7����d@з^Z9�z��>:h_)��#ZK�[>{����l��s1v�0yw�u,!�?d��'����Bx��t9����`�y��K���=�~�%���Zr���O|/�W�Kõ���ă��h�?4|-�ߡu���wF�Ә>9M����d�mX�F'q����8�1E�c��juBW��\�/��b��1X��|�!D�b�;��F�v���Vm3i˷��?%V��3a{��V��~�	^�b-L?*�q�ҙ�k�dVhn\��8~=k���N���P��ڟ�K�`ozQQ�K�a$7��j�||�b����|Q�ֱ>�*;)��1�=8�������*eC��lx�Q)t�tm��{]Eӝk�%�uG�f��K���Ȫ��p2�G[ϯ��}�J׿gB���4�^����잼�lyx�膮y����K�%��td�=7Pǔ���M_>��;=������w\��(*,�^�>jg)��:�b@ƅZ3:ow{&N�U��+��)L��c_p�]uZm��x���7�p��Rڙ��Tٷ��y�i��oX��	vE+�@��W���� }_}T� �=�o =�k�E�46.�ϻWX���E0���^�x���_�@~��W0*�0�OBv��?!Վ'Q-�x�w'r�cK/b��υ�=�xj��U����.Q=M��~��2!o-����wv�7�\%C6�\���&�Xs2����|��+�Afe�s���!��^yJͺY2v�ӌ�E�Z��y3`���86Ӽ�S��IՆQLy�(��6�����/qa��`�c]��bζ˯�xa�=�D-1M(�ej��{6x�Ԧ)�U%������u<��L�Յ�u�;5��X	#��e,<�_M�^���z��.����8� 0����T�FVkN�˱5��k�X��Ja#��fqh�K<��n�D{�)�?���
�K�+A������h{�wK�#���wF�gЭN�-d64@g��F�,UE'7֯�=��m����������o,�H����G5�D3tꢵN�l&�l�R���%��ϱؚ�5}paY�D�99:�ډ��Lc[��}e���UIjlK�Ȭ�M�������]B^0}��5=�43.�"?L��P�@`��v]jUBVu3�^l�H$0�ӕ�˝��<]�LT��v筹�8ƽ���Q�XaQ��7@̇��@��@���/��ۖ�H����P�d�.xN
y��~}������c�M�M���(�~��J���!;�����;�B�g�
��7��!�VH�ǰ��b���3�.��DUC�w�޽g-�_��8*��������߬�Q5��Ѵ�^�fE�Աjr�^Tۮ�ݵWYl�p�����!C1���^Ǌ�5� &��+�S���	�칇�r��l ��W��O�C�gW�c-��j�P5�4���鿭�����	��S+yx�t��a�~}�W��C˛�[��1�T��ʩ�����mH&��&����f������2|Q�i~k�ik���r�N��鞎"�P-HȟsH�k��R��ؔ�j1���,ZڄՁ�I_%��`�F<|k��#�,٥�%&�|��>��4�94��	��J��sz�M�����L!h��r��ޙ�U�b�<��K%�V���h��_�9t���H���N�YU)��H}�0ܙ�ս��-���Sn��P�Hl�ѳq�����~P�g������`y���ܝ۝e�B5E�=�����Xz�U���� ���ŵ�̌F�y3�}�#�����#?LA�(��_Bq������Jڋ�jx��ӳz����
:M�޴f�u�X���-���7��R�RjZ&�y�6��yw!�l�<R���N�v��3�I[��a��vʇ��ٳZ���rf��A �o+gl��B��G�O�����_��G��⮒��1��SaM�S`�l�m�~?����ϯ��}~N�(o~V�ЊIW'�PK�Ҥv����V�`� ֆ�'�Eh?mܢ'���T���o����2�X�3�55�������Ýn�秬�F�k�Gɋ��4�yU�9a���1^j��yOŖl���|}yќ���~ީ��ٛ3�j��ý������E]���7����t�j�F>�Z�*yFE�'R����=v��L�=YIeZ�<�*��Yr��g���l�`���r�9֩�-��R2F��g
꺻$��"f0i����u�LdW�M��{"Č��S��D[h�HL�`���GTidV�D��^Tn�N���֎�dt�̩f�v��5�%��oG��ar�ңa&j>{BQ�yR�N��X�s�3�VM�.f+�G�`^eT��i�+��A���a����7N��]�hx�|dm�&���K�c.�rl~}B�E����{n����)�W�.��(�qn˃��(�'����iڜ���.hJ�잔��5x�+ȯ�z"�H�3�������yЃ&���m���6��R�Tá�>a1Ǯ�v�)ݟ,"ӜFU��<t�u�U��x@�"��(V��Y��Ccj��T�_n+7�|�����nx]�ZX�/T륳f��S��˒ئPۃ;gc\���3v�8���*]σI��%��
VEv�?T�]��q�v|��?O���|����%㟟vE��y��%���b�����t��i�;���ݸ�޵}��ꈮp��Cb�~EH��E��=�[E[R�C+�)x��܁O{:1�a��ҭ�C75`�yKu��T��PLU�l����Ǫ.\���C<c	SO�2}���{j�3{����C2 �N�ә�ܵ���:�/����V-�֪��H�_|{p�o����upU����x>(��G��3���;���>�c=��G,u�������Ѽwp�JهzLw�:FW�=��Vl_��T��Y���¼���d_��+wcO]��8�^9du�R������J�[���7`����5H���}�yﲸ��.�0��Ξ�Q9Q!Լ�~��:��ԝ�������5g��������9J�{��B�\ҞP23ddG����E�4T��f674t���ԨcRΑ=36�W�Z��l�O��H�ʺ4�z���Q�{�>�u��[�l�Q����,�.�`���3E�z^i���1N��	<3��NN^�.������'��{�w%%^��U��ӻ�/L��<u(�f�g��8[��X	 �AC��[dFk�tu��}�S̱�����0"�G��OvB�v��Vḻ�o*(Z�n���\H��}!���pb�R�哕����}?P���6��LC
�3�\�R)����n��÷s���1�o�'�H�?f�h�{��V��J�U�(�QP��j��t��U��㚨o�|DnU�f>�{�	�O��ivL�2����p�~�z�Y�K����W���nR��z'��0�ж�q���U/B�c@�A�꒤��̅�s�=��"��j^�8��m�}����\1R*�f�e���,(bR��u�^���]`�Vg��o<
S����=j�ۑ7��$�y��%��%Ѩ����%1�=��׈Z{��9ut�C+nr�Z���̹�<��V���;�*��q�+6��4[z<;��c׆أ��;��1���g{��߯�g<b2�����	�K6�kϕ����VV��]��^�é�۴�3�ך��]�Ga��#yJ.�!'Gͪm�s�Q��c��İ\1���zg��.�:�OW�[ውyOɺ(�|�<�yO#�LPze0&a7'��s�&�uC���vc��wTH���ڻM>V8�����te|:SU�w�{zr����*�ч�|~��D�.�\-����T5�-GM�T�٬���v����.>�3n'���ۖ�*�U�cQN0��uk$dF��e�X	{np�Y0��&p+C&'�-ÞI}�ӮY����Տ�8U�ܼ"�C��M��؛�(A����V�:�
������+ꪠ>aS.�vACl~�o����|���~�S�w�G��vDj0�mx�'VʡA��`�!�XdD=徿GكLz��nR�����e
^�ه�oO'���{ti:ϡ�� �Zb�a���"�8>�>�������ڻ�(b��ꨦR�&���rRc"�G4]*�mj���#Q4��V��5/l��n�խ���n�w�A�j�`�Y�sLX��9��V�ƷPdµ�8U��鵾�)�E�rq���w�9ρ>k�h�>��#b�H�yY<�G�]6dcb�,��0���Z��E��tԛ���8����_��R1�V�[��sDtV���6͡������K�Oe�c�L��zwn+[L\[-K؄�$�>͕�V�&j�="��$D���Q�8a3�1���Du�&��ܙ֮�E���y��z�ݦT�餂��J"25��`A�o/��,�1bxDvX����i���i�#US[g	�iH�4��M+�,E�+�[Q�R�/8�1�����9��]E�T�1�T��rC�j�K'KL�.;:��Y�v�۟T/xLy���g����z���_��{���>7��jOl���; Z����� pƳ�v���\�����]�ʐ�_8��F�� ���*�.�+�v�{�-	��,�jdSKY�)ٵ���^�Xs"�O'Y,1���jj�6���K{�%l��SYg�ٛ�Qڐ�\��t��m���B�%�oL�0Yvݧy\;)v�P��Rmmp{j��zl���e�΂�V�����<��8R���=ןKPvk�ɒ�2!��w�]D3�j���<���U�/|�J�uK;����jL�Ô�ڬ��緉��ݭM
\/�[T�b��x5��r�8�Q�0���WŹ���f`�/\w��KW�veD67�ݛ�ݪ��XE���O�}��
[̕WG$���*��gι*�|ڔnf�jN�}�GK�@�5��VS�d<t���)N�WE��x`�ǎ
�%���qŔ�`X&I�n��S��8ƽ�ۧ��,�#+Zv�(Wv&8��.䅉�l9x�ъ������ZT������Z�:�b^G�N��Y�D���� �q�#TIa�9��m���grx+]�೧X�]c�8Z��0��L�V2�ЩY'*�����Y�����Ր�T�ʦ���k$��m[~`�8m.�*�k_&��~6sM����R��V���V�"qC��S6TG 4�eqY\��K�^���^H56�s.I��/��󩏁s4�ݼ\[�}%�3-h ��p�$g9vsE�u�5�_��%ko7v�ă>M�4UmTF�V�ѹ[D���T�0�v��Y��QsG+��q�Na�ʵ5J&�����r�,�E�4,��wJ��Qɀ�H7yu*˛e�M�5�6����ж����Iभ���b�Ս�ҀWr���k(�Y�ee�|��vꇍmB�&�/���[g��YR�n:�M�SK��-���/^
D	���o�T�����Z�<X&Xc��m'p���\��� �ck�
ʸl�e�3�x(�gms�4#ک����Q�g�긛S9��f9b��l�2(U�{�Q�@p�R:�<Y�xH��+CԲ�*+x��)Ú����z�VLR�+F�y��P՗s�eym55]>1�0�p�#w.	O�ŵ����&M�-
��l�]��ށ�寐5��L���ưd�Q�w0r'2Z�FQ�n�딪�`.��q-�V��S�Ҧ�.�t���ˏ;��qs��'��v�n��yi`S��hr�m<Ckwj�5��a�z�j8i�4�'H=����,�Pe����a@��Qa��*�}�Y4���p&�Ep���MٵgM'��V�w�1m��]�4�Iv6:�G��*��^:k�p�*�*ω��R6�ҏ*T�j_<6"{�m���5ϵ�k�	M�B�HM]R��)��s#<��վ�yU����AlHb���b�.��y��=�өmȫ{<��tv�m@�2�K6��f�o 0����B=yuؚ׵���� �D�TI4h�]=7osI�Fwn��N������C��#�*��APjڋ.�H��:E$;�Z��e�d�(�G;�a	\�;�r**�R��UQ�T��2Ĉ����-՗.c;��3$����<�y����e%�R��Z��^NE+���HN�(��Y�!T�\�3���J�l�Ng�+�WJ�L�s�D�f'��NH�HUGrO"��(Q�y;�J�+�;�"�w�s "�t�!
�i2�C"���K��-��Y'#MC�E*2�e�%Vʠ����':9IS���ܪ�qR�E�w;���9�Qć�p��� ��qV9��J9��вNR����rJ���z�W�٩P 61e=�s��Og�(����ƪ�-���/��Z���=5�*�Q�z�[�JM��Gj@���vJ�ZOi���z�;e�j�.�e����?��M��ve2�Gl�L��p~�_�����~tW&�D�_,w�߮�BO��ٿ
��2��Ys�(�Ӧ�z�X_2��gs�Y����+�O�LwS�v[����fL˟��;0����H�xN���3^#��va"a��6j�[m��=��mx4�����3�Lq�/ĭڬ%�j�y�m��j�p�cK�>�j��;���a��cQP19?�ԗ+>�f�Q�t��釛�U٘����NԽ�T7���1b,���'h�(=uOَ��e"�p�m�jV�O�0���z��{���Dpm�����#�����J��dW�eE�ܶ0B��ֹv�0��Qn^��_�Ձ�V�oY^�Pq�)�b�0�فqy>>�<��Ah�W���f1����S��[�է��K<Ǭ�j1�d:��dp����>�j�)O(�# Y��"�>uCv}X�8H����9�L.�9�ODX���\����R�#6�d���]k�j�H����#�qz��r�_���{2�y�<1���f���u�Ȍ��d��2i�/K1�S�����h�D$�¡��˜]ʛ�#�)8�鵹p)[(-�*&��n^�-d��s�3������t���|�ܯ<�����N8��ﯝܡZ�d�Ʊ꼦���j<����Ʋ�p�Ѭ�r��[�^�n�k�j4��U��f�f ��Y�3]������ \�e�2�.���|GKZC�3e�%a�G4���-�I�B7�܂����F(J�$��L���mϛͥ�&H�X#�mr6�	���a^M��2��e�	F�n��ک�:5�R��y�5��<s5�k.���	�k��4��/Bj<����mtW�_c�bR���c�m�r�$Fbl~1Yӂ龷�7��]�0�yw�U(Y�= :�'�f��2�����p<s���k���닦Ŵnc+�5ͬkCVֵ߻�]3y����o�T��JG�1ŏ-�h蓏���w5;qp��p�i鎋�5�m�QE��H�Ĕ�=��ll<�c;~�_ƻ�Ɂ�/~Dk���}C�1bĠUiY�ۨDcul)TiŃ&W=��ӓ��^זV0֢nr^�ǲ�3�0r�=��B^��n��x��� =�R�������vv�oE��`"��E��S��Ox�GW�ȶ�pmK�P�x�T�����^C�	� ��\L��c�d�8�	�E�g�.�ؑ�qRTW\־��m�έ�5�י���d(g<�%�?�O<�)���&�r�4�HǸ���<��^Cém#	��
u�+/>=�fGAZ7��-N���,���+l�������q��oԭ,�}F��6��P�H�$orut>��-�]�K3)r��6�'oH�	��-�'����$
��m\��^�u���(��r���������|<`��<��<�dva�`P)�������ߏ��<�{��"��(lvo����#����y�E�n/���-"����v��vи�q�m_
n����:��7s��>{�����_Fmd��G�i����V����	�ݹ>�K\�����2S@��gS��H��Z`Fr��z�r��D-"i�U�F>UѦsW�i�Y�Ko�^���{|>1��w��oey�I�%?oF�|�r�7��J�B`ک��Z���\�'�,���.gP����-qܣ�~�������"_Tw��z� c{��꒹u����5f$r�ıʥЖ�|��P\�dC�㚽����7q��.&�v���.��r����vz�OQ]�J������E�^�����xjW"�uY�OD�=C�{�/2��l�&���ݬ�=;cC�}c�/��A��XIU�(M��͟a���?����J���s�z�4d⺵WEh���}���h;K���w\�����b��� @���
�Ph��_H%�&�~���_-���|o}o�r�tn�'����9�~Ô/m*�qn�)�o�cM{g�6�Ȯ��C�S�M%\��k/&+�Y`��U���߷��^����O/�)�ţ�VK���D8��0W]�~j@�޷�f2��rl���Ր�nK8���u�#u{e����k��m�ǡ�J�f˳׀bY��&U�Ltգ;�~�0.q��@6f���0�0f��䖩��S�-hc���o��6�k&��qF��$��)�&ά��
��^w�a' ��wa+<�{]K[Y=�=���T�Y"��^V�&/���btYE1���.������x��=s62K�9��"�#"��mz�����w���(fE�̃�o:��z&S�MJb�]�]Ef�ҽ�k�V׉ԓ��hO�
J���L���CsUk=Ɉ̍5M����8��gl�͗|EMb�p��U�-#%��3�%l=��V+E0��_"쁒
6������s��IӓK���u惓K���&�f��q�6��<�G��H��}
�� �Bb��� ��y{�-��=��S�0�s���Z��`��-�'��L�Z~g�UT�Ǟ��X�A�ĴlBI��s'��{Ak��b	�־��hJ��iL�8<c߫���~�G🅏�U������w�\��0MZ��6�݀�"�z�d@��G$WE���*�11ZT>��x׎.w��b��^�u¾�y��[�)l��
�����l�Z��{���m*�_|��#��y�3�ª�����'Ց&L%^��Q� @r�,<\�1��wfS)��y`!iCZC�B%���f7���>҇���X�����R�x?H�6��;�]��e���D091�<�S�#���-y��3ռ���o|�Lsa����+9ʠ�۬���*��L.2!�`<����l�\�Ҷ�ew���Dhm�xo9 �8���d5+�7��OH��y�/�O�'wZ7�t�s�k�� ����<nڛ[�C�$2E�E�w�ܢ1�v���[��/Ov�����h�d��9^�)�5�D��5M�y�Jh�Rm"����nȪ�,��^��Y,�d��=���a	�*le�qm0�p=�	h͚�j�B�j�Y?_��2�k{h�,Y��V�lhm�0��ouYX������|L�Q4����N���|�m���YM�xy������2�?T)m}�w�j�"d�Ro�nt\d
��:�����jD/��ؽ�zn��z3�ҏ�ѓ�&��.�GL۩�����m��$���]����P���V�F��	���[�u�Ws<͐V����9�ʗ8����(�5�������5�KgYG���?�%��VCթV㞻�W�����,5BjzF%��o\��	�D��^��Wm.���v:8g�X�fد�.�8���Xr�Z�EnZ�O����*e�qI`)�
U^N5�IQ��c-�T;kjL	�f�,5��uՇg�]���4˘�:�Q�w�����uw���`bZ�c����#�/(�/E���#��_
�R�[�yE�ܠ�|G}S�f&�S'���j�J��[u*�����+]��U]�)\���Joך��H�}��W���.2��Qp.2���GUb]�z�
�5���u2�qe�l�ޫg��1ނ��ez�����%�$ϩ�d����w���W�r~4C@��lYc�G���R!U�E)�eNHfFc�U:rF+$�.��咟��}6W���!������`e-����G�]kw
�]΂�c:$O=˟M�GwN��i��X��;��0p34^�E�ȋm�L�g��`�*x#ZO�}\
���}u��	��Nc�����vu1�����AS�J�5�Rf(+Ѥ�[�+����lZ�=���y�)�x�/'ɣיU-[�i�
�5vڕ��C}��u/"��\���exOm��M����G�@խ�)��i�[��Mz��O��mz	\�eӛg'1�ݫW��r��I�#�����M�$�O�T������>hf�D�YϦυc�x�1`�'���o�����~�aִ5mSj98ի�]ᭃj��=��p3<�b'��q�[3h�}�X:��&���Ļ[3%m:������s�T�m��s��n���O���� ��^07�6G�2~�~���J�shtW-@[��n�ňoF_,���B���G���ۺy���~�xp�61z�uk7/&���%#���<zʧ^˜%X�Dt�wz��ަ�<,>����
��#oTT.�(I�Mk���M�ر+���NTŴt�T����p��wY'[��G8�ѿϷ�(
(#�p. �y�3 � �T�墊B�ߒ�a#c��"��t���T/k֫kP'&0�O�eP7�����P�D{�"dM_�W��ߔ����;'װ�7�чB�;y���u]����gKv:'ųK3�Oޟr��W�-�"}�A�p�%3�o����CP���=��0�_�{yݩ��в��`1��1$��0�˲L'��r͹��W1'65�^�1���P��k��	ۓ�lt,k���"]zm���9-�=zD>}JD(�ڼ%W<��4-��Dkv�]:�]�}§qkZ�4��Z��5��>��Ҥ��`�ң���L�C+Y��'U�cوS����5#��d���P��Z]B�g@����R7]�;�5��~	���>�>��X���x�{���< *��:����e�f&��qx�w��y�׌����z�%z͝�M��;܎&7c�K��ER�^�黒o�|-���6i,5+�v�`�G(�b.7:|�U��C�+W�J�b-Gʺ�D5pw�2��3-!>��~��_�4����̧����e��J�+�����/�Lz�]�6�v%�:�����+����T�8]f4VԽ��P6[�1���O-r�a�2r���H�F�q��0�K�O��ѹA�l�*3���LHA�����u�	g�T��K��8Ek����-]��.3�π� ��?��@�3 �৹c8�4�2�o���;<�P�:��o�_YZQ�U//ߎ���K�W8n���!���<�l���ι�XïatN�
���IGly&`d�Kd7��>���<�|���x���E���{j�`y�,�'^�t��Ȥ��N�l�$�uCjKG�Atj
�/�W���yR]s����9>�\�U�#��'ƚ��˟�}�r+���avӰ��vԧ����Nf�����i[y�ӭ�8�,�6�k Z�L�-nfR~���x�	��H�Z��_�=�m�Ƭ4pbԄ��'꾅I�����
��	��T���$��(�<��8�UF�v��G^����������F�ʷs����*@Mр֞�΃��_,xh�r���^�o䧱����{��|Ą{w��n	�Ԅ��0�J��	�90��c�j�y���Q�tt]Gy���J�{.��R�ąv�XX�,�9oO0�-��}nmp@��$��f�xd~�jwz���XƩ��*<�u�,�T�q�Ki�՘�q^�" �>�jkYd\o�>Q�7��=�۹���
!�f�+���a���*eeL/&b��SGS:�/w�v�U뽆]_8�7x�F� f{9N�pF�wP??y�ݍ�Í��a��?[-ˮ��<��,i}Sc����Nv^�xwm[�.�ֻ{]������90j!<�~??�ߟ�^�{��? ���@�\ ��Q��Z��]��u�bE�b\�#�����N��I�����e��=�󍺒c��s%g,���w�t8��~TS(,$@}k��Lk�J��9;Z��&1��s����-�ru���ݴH���N4y��k��	G$]@%j�P��F���� B<���^9��f�66���򵭻�zV��x9HN���1�OU�7,���[-�lأ'�����6��N~�i��{B���մ������f#���4@�w��3��rƔ��2"K�XCaP2乛�k-��G4iڷQ9	>�Ws&��jw�s�`EM��A@;kȉ�h�H	��B�^9��G)�&k�<�ˌ����Z5���Lw��_�'z�4Q�[J�V=�Z�*��*!�1߽}��ʾ��yd�m�>�כj`i���R2'Ŵl�R�ͅ�L��{2�i�GMS�^kܮ��Xs�²�5T��D�/����g%��{��OX`D�K.!�eٳ)cpܥ�0f�k�)gi�Y���ӄN��C=E�$hŒAo�p��?R�X�ܐ��Дl�*�׬~��p����{V��%��Vsar�We[)QoCvz����(񋉷(P��-�v�H���5�%l�x�8�Wb�>&�zwK��J�
��Y1�+T:�f�ú�E��&q�m㺓�ٺ�=ͳ x��Wu�BE�/�:���X�=�a�� ?� ��-� f 3
鲇�i�)n�΢[ɹ�Y1�3���m+�Lx�ZD�	I�ބl�`|q�ퟞ�m(�m�_X���xA᝝���ҮO�s������JV�5���cfq����3dwK�_�Muܕ3�rV)�t�N@��g���"(�\��A.� �Gk�{nm�/��cEͮ��5J::7q�
�C&� �6�T�n�2Z���R�k�uE�����L,�+;$��j�r���B9��pLX-v@Pu��Y��P���}x����Z2_#�{0ni�4Un�}��k��Ö|���Y�lY9�!k�2q{VҖ9��y#�:���W�}��`���mO|+��n@W l��w�R�8��6��@j�X��j�:!�N�eE���!�ڄ�������3�9�^Ԭf�6"ujR#��5�^�hkXFi����umg̵��>���3�;�7h;G�z<vݸ0-w�H"J�Nمʆ(J�_{��}my�����?�u��埗�N�zJ��⪦%aV�z���T��޵,�@�m!� }��w����z�^�g���<���o����[d1-�����F�����c��*VM"N6�U�@^���֑)�C�gjL�[��n�F:S/y^Z��jf(��5ڨ�V�0м��Y07�H��C#��ɽr�C�c�S����Y�����9�Ԋ -fa�4Σ]���4H���u`��َ�0*$5�'�K���V`+dUF���ҭ&���u���T��[Cf��r�_:�*�vV�}Х�3\l2�O�Z\�è�XY�j8�2儓B��³�5�N�$��V���k^_q];v���	����]�{΃
u)�K��!0�:m�H	�m�s�ƌ��ڂ�к�ğ7)�ꭳ-��m��;dӷҳ��I���-x�����bhD��2!��ˮ��#����hzT׃��ș{�25�]6r룺x@م�9���*P/D��fK�.�i���$1����T�T��Z�rR�
Q[  (	����e=�}Ow�׳���Q�}�M�[m��[Q=�//2��R����[�.!�#�(ݗ��+�ܳ��=u��<�����hutT�vw�*48˗F�ǆ�C��N��5k�|4��m��D*�=w��u�qQP�9�uJ፳\��8D�HzT�w�m�b�k�^*���3֎0���
��C�s+�OK�/�vq��ѳo
�P��``���W(�2�wx��L]k*��S\���\���WZ_d�u�D�D*m;=]�w4�5��ɶ�8!%KS��(˫U8�<]���+�8�߾;�-ds�[�@�1Gr�,�spK°�w9]`��D6�ٍsyk��<�l�LY�rdw5�i�՘�ǜm$.�C��r��k;ڴM��FX.cXNci3����nL���&<)��H���*����c�mL��˝M�D�a�=ڴ&9�fv�/wF<t����^r��+&0��V��b6a�	�c�6�f��j]����� LX]�kӂ�ܶ�A˕-�n�P�Jj�4���M#�s_M�q�v��\%v2�w<t(+�+8<�]D��j��	��V+2�iq�������y�f���z J;�N�t����ƥ@�c�7��n:V.�Z���TL�i;��
c�ҧ)r:XE���Wmչ�V��%�ʄ�j����c֨���wel���:�Bg4Z�T	�C:�Й#us�5�]��6�LF�(n�B�H �t!�Yt���̳�$0�M���QJ��Q>���K����r��4,��Ƹ�'G�TqD��Fgn���������I�z���7�kK.��:5{�"���3��ޡx�,�h��$�kq��i�>���|�eB38*0IG�k�Cn�� ]�o�6^�7���I]H�n0����l�Ⱥ�z�!D�����'h̷�vr�HU�ݹ\V@�S}Q���!t�A�C����.TeVj�%Y�}H�"L��|�O=��D��s�.JBUY�S&�xl�á���-B��؜ry8s�
Ȉ.r*�7��I1�5C��juM�N��v^q�!'<�Dr;���pĔ��{��W
�0#$ �p�R��h�Y�m��9vS�
��z�컝ՉEQ�Μ(�q��{�NF���Yy��K�!�r�aP��>�������p'4�"UA9��:K�{�������r��r����F$�*�*Ud�U��17��+�_;τU_!�#̊��>���e�/���Q�C�o/�OT�Z���Gs�NdU:�R�Uʤ:�AA<�TWrH.Q@�$� ua����O�@�B��$P���}��'�i��y���=���j��G�R{1C(s�=��c�$	p�M;$L�	�}ԃ����>�~?|~$�N�TeaN֮0�W���>,��
��ŧt蠮U_��s�+`��N��=���Qw2�evRT���nQc�n)Kܤ5T���T!���j����]��f#���:�*$e-Y$f�ǟ�D6o��ֻ��i3 ��p����|�Po%#�C���wE���:�3�w�Ө��_�O�a^�O	�]��@����?{z5�]{6�����Ƀ��3�H��Rh?�r�_nu����E�}�q	�f��<��H�V�kP�v�^�ly���P�3X1VV�ٝds�1� ��W#ω��"���%e��*
z��~J�/@,[C�w��Lѹ�w��W:�)�v\�Y���Pډ�L�8d����#޼�3��Wxr^�Ú����z�fr�ڨ޲P��R���"���7�����l0�P]O�^���+K�t�*ڥYн��cW�=t����*�t�7�,.xD �橷)��T�őq�������_,z��)-T�m��4'�-l��؜3�k4W�	��̓VƳ�O�=%S�����S[>'v�lkM���B��Y��R��I�2-�]��;�r�jGq���PڃV�!�����ߣީ���,�g-Vû���SG��j�E�Ĺu�f'i@.)�l�tά&R�8�f;qR���xN8�]��v
5������$�P�Y��*����>���+12�N�z��s�y��C�Fu8�܆�G~���&��7]�N�I����[J���=7��	\bC�&%�@co����45�Nm����~1�3LD�5�C�[Q>�p�iyܾ��x'׫33ل�K��0qb(# j���X�7�g�/h���;S�B��0����T�u��2n5�"͏L��]��b-���ȟ���Y��_mU8g�pK8�i���3��;n���(��o�	��%�0g�{��v).��v�P�^��Խc�j��M�tr�a�(F���}=���е2���J�l�5M���f��ơ��z#� 1R)��G��+_��_Wڦ���ڳ��F)���:���y�����D߆t�dWT6�%��%Ѥ��z�h35��|��z)}�s��i娨vzG�q���Ǳz��,�uH�)V���.ɉ�*ͽ��Ҩ�!a3��i4kz9[N5z]q>�oAf�ju�VuQ�k1	GO��"o��Ev��e��#&�SD��,���}w��#*�:e����	�Ύ�u���}SW�������l��Y���u����zg�F٧s��>�W�{_QhEn"�Ҷ�mc-�zg��GD�Z�r�z50heZ�ʀhqܖx6��Ks�'5������R���l�a=f�5o�	������|�t镛���Ias�r�@&ɘ'͎�.;U5��Lz'��x ��7��7������W	�{��㼱�\�⺼���,u����x�3�~mلݞ���-1H���{�ᷝe=;��F�l����D����R��;�v���$wGZ�C�,��Z�nN2��C�j׸�F�	�$��V�ٯ�;*�Ӏ��<��}�a��S�9#%���":��Vdb6	
%�y��|a�P�
������;є=Y�������ҨUi]w�0;}]<����2�JK�£8t�sp��]PcN�����j�	�X3@{��S1�̼����-�ux]wl�RS��?t̛*��"�jҳzqB���P���]�|m�V}�px���{O��V�����8̒ٮi�{�+�s���>��. ��f��I^�h�k�v�S'�z���Ǩ�2u�߆�a4�Ϝc������ev�D�Dq��AK�x���w������}5�S��V��YEa�b�kdp��t�O��ƛޒ]��|D06��<W)�j�Kpn="1�<���?Os1�����h��p�wd^Tc-͙kk�����ia�o���a��Eꯕ���ۙɖS���pT���ۉ���>�:.Ź2m>!�y�ʘ���\�q���j�{�d��!J�o�8�@��(�JY��Y�}Qm� ��)tE�z����SW�L��ژa�%����3�YK�t����z������}���]�<C���1Ǧ�\��k�	�jf�j�mn�!6U��E]?���j֑[�4�yY7$�GE��ue�� �{�f�0c��^�b��{�m��2sAd�-k��	h��R�*��j=�m~���?fJ��[����"��o��gn.�j�@��d�,4�[�i�VU�r��'X�*����eV5��d�	��~�bG���&����#M=�����6F��S��u��X�ۗ�ɒ]:�N�X*�7v%V�^Y�y�=5���?⑳��+y�;��Q}�К��(k���א����Ң����ֺ0���X|:X�T,c=|���Y�թ]�}~�Ub�$T�{�y�k��3�i6=ja�����D���Q�9�R;^�F75����И���r$�-vu�P�MZ?����l׻-}:|k{���b�9�W<o�'K4��E��fz��G$k�@	���r�U�(��k3�o�?d�a�E���:�h�ش*�wZ�V7�ҁ��i�3�~�%��5Y�0���ڨ�Z���>����<F�g�<<��+7"D�"�C�������i	{���i̕�Wz�5�h3�xnt�J�3��nTb���ᒄ���3�S�(����.}�9S3(f0ɮ9 �;X��=���d���2TP�ّI6�ڼ�I��X�A��Oy�h�}�UYɞ�L���|L�~L��l�\>S^��gXgB6�>l�zD�����}yZ�����Xs!��7a���×5�2:K�����R��rE�ؙ�?k~�[h�MuG��[ETL�a�!Wig��z0�!]�i[�~��ܣ��ƚ���oG�"�k˒�Ƕ�n�oϝ�����JO��^�`G<�"%������fM�^s�w���GUF�lec���Wr�ןp��~�v��)^�Ɉ�S`?<��}��8�=}���<�B��u� T���Ð���p�@fyڇ�v�V�6�b���CUJ27�W���*~� ��ʺ�9�9(��b����v�}�ڥ��
}jg����@��I��h�"��	�HyeW�R2޹f�i�'�זE��d��F�����u�WE'��l�%9�vT�>�xfò�2`��Q���9<Q8}�WbRxG\#�WF��*�8�ҥs�*-99���Z�)���,+؎���>�?��|����_�x�+��kג�7�ѧ Z�o? ����T	v 0��h�m�8`�Ⱥ�R�9o�����s�I�+6�p��S�+�]���ŗY�(��l�]t4�2
g�a��t�t/���i��-U�ak�fj�+W`�z��Q���*#�4�]������71I�C�U䬏����:�d!�ܖ�ǁ�gm)V��d`M�� {d֋�ȶc?�����#ٙ!�b������<c=Z��}��9H�3T����86�J��v�뽇է��v߆��cL�"�.���T!G?��ؤS\ؽ���@��+'"�3y�9��9ģ.�Ws�%�#%��c*��$m+B�C皤Q���[�y\��[7kz�Oʤq׌�Cޫ�����)�K�Qg��`+������E�(D��A�d�H؍����/��ƥ1�Geq�$�'�$hcH���f����%�oY �]��ߣ/����?�i!Q�O?��<���.ݔ��]q��}�Ek�I�=_��C��RǾ��糱�� s�%����6��a��&�'~��VU�����*q!���՚9�_��Uߦo�r=!!}�+_�Ֆ�������PrtQ�㜼(/����g}�MoO�E_t�SUۅy�6�f�D�����vǒ���p�G���*7�C��yW��1��	��>�k�t)yU/W���)�|g1����T;c�3얚�����X�n��ڤN��ybD��k+Ω)R��q��T�+�:F��k�D��k7�1�;��ž�ܶ&�����xfO�&���6�G�PLyBi��Ǌ����wyJ��l�u��X����W�w�f厤��:�J:��J���/wN�e+��%�e'L*��u�U�x��`>�p*^��1L$wt�{�t y����+��~Λ"Mw�j�KV��x��X��7"�ۇj(ފ����w�НA3"�r�P�����>0�Ǳxb�O��YB����q��޻T���S={s��;��ܲ�K�'	tc��Pr��k+���ɭkfQ~§Ȝ��D�
��*��mU�AN�VepK��ױO��Z|�
���K�˫� ���!�F�_��id�nM�������U�Gy�2�bX;d��k����U7#򐛣�x-�����:��;��NY1ٴ���L)��>:�,�(4X�
:���e%NqOɺ8���W:��Gu�n��$CM�b��\	��FW�{������u����jJ�8�H�VW@�
yj�T�La>�<�᮳=�7k��`���g~�C�m�-��-Gs�JZ�����\��LlɶOo۲]�ݰɎ#���	�"!�-�E2�ӽe�d���䧢⼲9�X�	��h��G��0w��Z�D�LMf�Pm�³�=x���ᕻh ���j�V���-��O��*�,�w��W�d�n5!]>ٸ����G�8:����N3)����8d�ǉ����2�ŕ������j�祋�=��xō�Ո4�b^��O�N�e����d���$�k=��W-��v�hY|�in��V�������m)3*f��j��t~'��� ��j��x����_�U8U�ɘ�vCGk&���]�E�i���tS����>��I�y7��˖�R,�fF�}�3�L��L� ���j.�ʥ�������:�##�MMlm+�ߺ�,�ʏ5�KI�:��o�,Z����$`�6���ͳ���K���mr�(�c��f}���B]�5�G|�ձ#�G�u:>9�U2dص�Z������i�>�X�|�ӰQs9׳�v̑���/��G~�E1΁�6%,_��3���pt��T����%4W�H-��=�{�S�fjU��L�$΋��RڌR�|m�ћj㩞�(H͚�j�B�n��{h,2���zq�L��ػ��:��v���w)�J�[UJ���3�CE����Dn;�d�κ���ke�`��e1�*��s�T�u �+QQy0*��&����#S�1ǱeЉZw��7����Jj+�VF�~�yN�P*�7v �[j�8�Ʀ���-m�wК^��ޡ	K��
�&r]r8z(>9?dj�O!�q�\W�Ү/��͗����^�%G^���ȇg��(z���=W���87VK}Q��:�6��.	����k<��<�|�ܹ��^�>�`���t5�h
ZBw�+�2�k�h���wu�Jd̺�Zi�n�_9+�,f�̉�qW4�E7���ae</�ϥsu���C�����ۨ];^�>�3Ǯ}	��Ӱ��D���J�\KτI*�=�b	tqԎ��p�]�[~��Bo&|W�32I��u��5+ֆ�'�Co�� ���i�Aot�<�:�a�E�gDȌ� �	����J�_�
��F�+"l�c	��x�V�����Z�����C��w?~퇅_v�����j��Һg|�d�0���6,��`(6�T�!U�j��aP����v�e�Hȍԡ��^��f}���3�s�S�E=��~�A?v� �e�� �1���TA]zE��H����#V�����jY���D�Զ���wd(�^�i_T�������� �UI��"�@�R���¢�z�՞���d�qgפ@�|J��e[�uS�w�%;���K��P�V����
P�9�y��c�2}�y�2׻Ɲ���M]X{�[O�뼽������f�	���U=,���w�)���N��'�9���Oe`�Ȓ��{n/#�.���.�_\�"���b���CUY�)�<�[��\���j���	��f'珑K'���r�\�F��t�����*쏁�|:VIj�wp��2_>64ѕ�+6�����
8WW&�Nu�V�<�,�-n�x����lg`��rma�R��ANV�9����5iʎ���,>k��\��R�3��j�G��x��[kt��}U��3}��{ɘ��ax��tɨ�,�oPc�fnߒfH=�^>�w�+��9�:r뢹h�x��3�X��1b}嗎yw>.3iθ��	*���5�o!��YMg;G*�ټ�ʫ�X��G}�e?%f~��'��6�<B�\_�ʣπg���M���G�q��48����Kn]����#��������~�k3e�w��1�E�����xp6��Ou��Ӝܑ��Ӱ��|���/��.CsH���b�c׌t����O�4�ëV^Lǚ��ZW׸ժ>�ݷ�ē �"�.���U
9f���T=P��+�[B�@����j��z�`E��Ʋ򠶧�Q�cOY�����*�t�7�-s�#��5.���0�뉖�z�ǆ�����
�夺<�]����l-�hOV�|�^Fv���V�!�K��0?N'ݬ��4}o�,U`�t��~Ŧa�s�)����K{��'��[pY�#h�V�+��S�=�qKw|+e̷�$�@�$N���R٧�l���^{w#4�����7�����z}>�O����>>o7����9�V�<n��K�]����d��V��f���f��Iۄ<%8�/�^O�T��)�Ե-u^_0$ٍ�/�Gc��mV�uu	촊�7:A���K��l&���l#�H��
W�w9�jG|�w��d��IȬ�(��^��]G�N��se�GGn��הfE7�Tc��ظb��`���I�-�O�[$��S*}}�.8�]{����Գ@:3�ݳ�v���1Nʠ�0�m; =R\v��Fʲ�Ml{X(��c�/[B1U�g
ku�#�ʈp���;�����wm��C/v1;��������>�-,��I� }��)���űte��d�4��鋛:�=ɸ���B�~O�e���ʀj�魗-�����wo5kv���M�"�r���u�Ύ�eIJ�
�i4��M�(^�̈́������WoGk���֖�:��#�#t��ăٷ2F��u�J<:mb�k��1���u�ׂ�}�g�x:��i�m�
�ok�i�-)�P�U��+��&@Iuq[��꼽���w��豬�EV��Cx�h
c��׻6S�J�55���3X©�4§p��l��T����X��TӖD-b�d���*��^��`t>F���IN��C:挄�ҡ�n��6�YhS��'wjZ�������-�{,�)���t��M�����l��(nky]�A���U�2^�� ��iYm��,a���Q��G�i�����c�U{�ԗW3��/���/�V1�X�V|k7�\�'���M}a�C�֍f1�Zv�HQ�dk�*o������a{4��\���2Y��b!\�sN�+U	b�0/�S$5�	}�Ss�5�����0�E�R�)���*��3(�E��8��E`&곁�T_#�l�	]a��Z�w��Tα�����of�1�	9�Ṳի9��Zx֜;Q6շV^D�v�]ʐ��ӭ<�n�:��B,GTw�8�4�-!ڬ�����+�-an��ee���=�Z�Z4Q�d���ӷ���������'��X��yB�n��V�اٕ�c$c��|�Y���\�m�����>�ʊ��Ū��]��n�2�uӬ�E�)|R�b�f�@ZΕ�;7^����s�����gR�U��ed��qrMF��-ۉZ����!)[Sr�Q]v��2l��t����O^�-�
R\
��P[�a����i�k�6�q0��uڗ0�nk�w:d�mQ�o��ߢ�t�=�.��cT�{72����eN�����4�p��6T���F��뗰�k2��5���_`)n��˨�*�7���F�T�Ç)���XN��u���6�{o���ҕ5�+:)ť��m�G��oNj�x�Ded�UZ���r�,Xsc%�	�	���]О��nD�m��	�i+��M[@�꼺�:�84�F�QK����a���I[�/�Q*�w�KF5�ct�P�۫@�2|�p>d6��|��*��닢lW�eM����J!�h*d Т��R��ª�$~�����o��I\��8��nw��XI�ѻ����E�"�dTU�2J>���DvUr�X��/n:Q�'A"�*�;�r�V˓��9:����َ^	}(�����eʣ�.%뺓I!���TOF�����ʝ^p���=Ұ��O+�YE˕L�������B/���9}I��sʊN�#ן8�rH�/R:�T��+��⌣�y!r�LN�Y���.�n�q�L��;�c�U�:p��E���E�({�+�w���r�F*oA�p��B�� 'zPPP��뷽#�Qg<�����H�wM���z����>D���ʎ===�+y'�=�'{�	ů4��wQȌ̕bdUb��dy9�T�*��9V��ng�v���NY;��'U����strO
�N�����S�{w>��'��x��;���^�]{�=��!�_�?&D����<�U���5X��U����IiF��鱔���ۤx���Ư����-̫�\}V�g'<:u,]M�)�UW�0&,nV�� ��1R��Z��g���ֿ�*ױz�;�ހǵ���Ok&lh������?���rfFS���K��t��Ѥ꒹Wء+�LE�U��^9ʨ/�:��}]B��n��;ޭ�.�R����^�-� ��g��ۺ��j��!�ȹ�VQO�p����{�1���;V�c �=��¡k�9����t57�I(�'���|r�����¥r���KuF!n�u��z�M����z�es���u���3��� V��5�n����"ɤ�*���|�L��g�W ����	L��y��Zݞ����L&)�آ�����[�9�̡֛�϶i�^i�Un9.�v�Gs�����X#��҇�^��h��lɢ��)��u($�AU�����_Tۡ��@r�z�;3(m������o2�?���ǉru�C@�3��j�[��d ��x���qyֻ�<BNl2�c�q)�H��]O����j7h�~�ǨF[ne>*��Y�3��H�2^�˯jO!��u�5�;�y�m���<7;�ք���0*ߚ�£�}վ�g� �	������+���ǆ�!;C&;!Xl���Km0X�(��z���d�8����\n�1t.V�RY75ba��]$���룖V���Pol9�_��Y�F�p'��ڎs��=8��IP�@��W>)-�
��քa���/��U'�=��\A9�52Vbf�=�+����ݼ�����`["�1�^V�P�ƲQ�t��{�徜"@�|U�����c�n����>�#�'�����o�5zf99��u�G��6�ިOi��ZO�|b"�uD��eތO.��u"�+�C�H%
�#|���|�D��|N��I����:�'*E[uC�'l>�1wԭv�~����뢹g��A�(T����}k깦L�:�sD
���a�N���o��a{juƹ�^���'d4v��oT����j����c��;���㭸w5�![R�k[��fjb���Q1��x�q;�R�៟k�#��Dw"�tOПN5�Ֆ����(p��^�}h�UT#U����Mc�ka��$����\�!�]]�	��a���OkI}k���:!�a�t��U�,ͭ:֍�6~����;�9��t����|�UZ��qȎ��Ԅ������w�F�2�q���ߒN�$�jl�~fG9U��솣{�d�í��*n����N	�0@����+�tT�"|Zw�V7��2���<S]PRm^��?,�Q�V&����嗢��m>U�5�sj��u�2��8���b.����Yǲ5�����7V���m�Y=e���d�}���~k��R��-�Q��i�Ӭ��'`@ܦ���*��nRok�)]�x�b��7���;��+�<�=�MNFN|���䦛������J���.�Z���.�)U(JO�5�W���v��&Н4MUowx�j#��T�a`��m*�)�j�n��X¼T^L
��W��4�#Q�1�{�O�Q����v�{�>�g%GI��W'��%:aeT����^7X�����u��"�yˋӱ�kg��W�_.�p8f8<9"���\�?f�eO'��)?5�tsu%+_�k1"��f{��=�R�����r��L��1�̈�mdӃѕ�����R���#��=՝~�����ɢ�'l�[��鑤B,;��5�Xn
��Y����n����SVaJữ�BG�b��X�UK�Ж=;��|��\=ޠM�B���@=}��\�&�C��QWo����i�vi�����-K+��>F�u��[%ؗ`p�Ŗ�`(���Fͩ}K���Ej#�M�|,�?��|s�������g���=.>���)i��ԉ�9�>[�ΗA��/[k2Q������]�KT�:#��s"�ZǺ6w��Ǥh�3G=��*�5��>M�pU��� ��8�㬧��6�t���՘���X��z���,�jLh����E�t�&��3��IB���޷�h�T�w�n�J�{���[YX�p7�,߷,�,�p)�:��qr�X�{\�U�Wq����B��f܏�����'�	�����K��&MW�j��xf�l���'$�&�
���;i��1�4�c��� �R�/�ӱr]U]]���ku%áp�œ���?����c��o'��/*��x˶���w$]�ꜹ�[��i��h�G��d���R��iG���K��+˵8_dg�q�7C㾹7KRU���?V����w����3�x;�ϮQ\�ہ�R��j��'�:�'�V�X�F����1��u�ZL�T�ݚ��F�ɤ]Ĳl�v����ֻ�.�w��h{��^(z�}݊��>�T*ίp��9��6W��t������]���s�<3�mOt�N7K�4�ے�*S.��#9!}�g9K�c�����f�?cR��̪<��NNT/��7���\��)��i|TÙY9/^��=�N#G&/�򸗄�=q��ӧ�X����"��fsh�B�E>��,[C�O�"��c=I�Y��J}�ap:cɛ1~�n^�Y�,���
�C�f(e�W(��O��~��ݷ��$�VE��s7d��5�f0<�+呓�2:��%���p2��v���\�6T5��U囜���?��O�]Ў�+X^��̝˵��`9��5r2��Dw�5$S�Q�cX��"NdvCF��2�z/�ISҮu��wR������r�r���L�XtK�/��<�{k��6~�F�K~��0�r�4��d㡫�u)T�f���ȇ`�XB�+�׼ӛysx3��v�^q�{��~�2+8�D_�\a|��"�����'ֳE}6��]�������8�����9�xTL�� ��>�X�`e���]w3C�@}�����Υtϳp����{��u"���CF��_5)�iDX�g�kڨs1'k��Y��td��aj�n�de���
[3X�E����+�	�i��"�v�Ƀ�z�&���^��)gDmU�}}�ב������׀̈́l�|N�+�P��A��F�ϥN��"bۓ�]���DJY�9���p`�K�p��^� �J�̞�-�%]"�vǒ���h�S����-nn�>rr�o*.�xi����/Ե���o>��3�I4G���]�Rg�-R�N�ݳ$��$.{�����
`J#(��u/�̩�][�t ����YB����V��R����ҍ~�ً�v�fm��mv�G�*5_�_G˜%3�y(������c�ؼ+���>�����b�H����������s{�ι���i�6�YL�&�F`�5����y�z��V��BW'j,�z��\6��s+���u����v���z:�9o��B���R�e3�h�\�RB�7�֨u\SnC,[�:�z��\��:��E���Ƈ`�t�z��V�V/��z=5'�����4w$��|]�B*���KgL���z�-��{�sY��w�:.!az\�܍�V/^���`r��z�>��i{�T�=.|�8!��֧b:���e��gH�͗A�-R��`�SI�2�c���r�t7MM�E�͖�#}�s�OfV�^���2qh��*N:/)�7�C��J��7'��L�?O6ג��((xRP�ߔ����q|�B��{iM�Q�n���Ts��9�~�!�)'�	�fηv�S	,�3���>�m��su-��<���6�7Nc��E,�+�8DG?5zd�c~��@�gy�Z��zy=Z�����q��Wp�2.v��.��+w�GйH�BW����+����TS)�eu���uP��S��z����WfwZ,���GB��]���v)8�hOŷ�><Mo@P�">aY�H��'�vf߲�9>~�=��k//��S�ws��U+3eo�#��0M�Dڕ�ȝ�/yl�7���|m3�0����*���efjc�Vj&�ޙ�!o���dIMl����!�;ꍅ��鬦��i�ۡ�B���Ucޭz�RxvQ��Kf[�]}�3�,�p�b�&�n�w۟��yv|��^�B�w��)�+����}&�[�r��G�\�������^2�=P��5՟<;#
�7���k+5*kSWn�tu�[�G�؄�����h�UT#�楋R�׼D�L&�4�4ΟV�S͌v��\yS�T�q�P�&o��"U�Å����˫��}oN����,?]{8�7�n,���
&�����E�Zu��*��F�5��&9�����3�K�p�E벨���i�D2҅��E�wk:���D��0�����ؔ�>7?*�ND���"Z"f�Ҽl�ee�CR�.o�f�u�a�*�bݧ��[���h� p�<Op։����� ਷�Ё����#f'�wD[�*�E�{T��
#��(o:tǩ.�a*'�;�{�+:�$���x���CС��WO��'�ߢK���6	�m9ۣ����ܘ&�1HK�is�kR��w�<k�-ُ�R�9Gt���
�ō�Pgt�����(�5��n+�90FE��/���]NnR<�a�X���S�a��Z��������ئ���/B(���Ll:e�9�..��t.�ں�y�C���_?21jI�b��CYXE���y�1���>?}��XWd@�}T�
��@�Ka��4��<�a=,r��N�x�4%$R�%��SU��'�9�68��%�)���Էz�vp�3+;B�6���:�YF@��E�ꈳt�q0yޖ�>���2���mNu��scrXUma�s�Bi��KT5�'��0r��9t��".�Y�|�<s�ѧ{:p{��5#X'p�`�7����/%����qk���6���n޴�HȤ[t�W���������1��ŭ������5dv��U�$q���܈��x�gA�C����������˪����:�Z��C˾����.�,m���'Y͚�-);���n���v��	ޯ�B�gCdl-�,��%G�
�����f}
�c�<3�6�95�F��_A�Օ
�ņ���^O�t�; %���J��7Vz�vg�K-��g.�swM���3�6�����l��i����K�G��O�)�6r���́�/y\�{����q���:�!<�FO����,e���t��{�R��5�Mٵ�UZ�4A��s�VMm{�d�}@�0�BW&�̥�ϔ�V�<��2�M՚0��ƶC�
������΄����*m+���1�M�53s��2m��g�7-50�n��o` @.��p���*i��N���V��z�1;Z@�@֎�)�$~[��Ņ��pֳ�Hc�t5XR�YB���7Tm���"�*m�pofoH�a�3�Z�|���	p�{>�>���u���n_%�)ύ�P[�k�g0��@D�nf):p�C=�[l���ަ�I�=|�9Д��EQ�-v�'�`��{"gd�ͥ@�|�ܪ�@Ms�!l�|�������s�M_vLb=WSr��2���=ʍfx���]!�Lì�oM©���W8i��d>vt�:w�a��^Qޱιۉ�z!ݶvYiv�i��*���sõΎ���&�z�q/��u<wVX~K[,_36�����P���:�s�Vl�w�g��͍�En.e J�{���0�m㒆S<��5hB�;� V'�Q`O<�s�J�tqk�ynY<�gdg�'#uI�%�M�vdf��;h�&=Y�8{Wky���BvB��;�ՙ�b;2'����h�zd��!��y���p��B�I��Ô�"#o���N�ttoUjCW&�/z�KX��oʝ"���p�r�����n^Ǚ�M��?��M5:�N:�TxmM�L����ڰ>�d�A>&|MK�]�=�l�AF�\$�����_a�����|��LW�_:�@��L�獣u+;��W}���
��+(�8�Q�5-^d���\�v��3%�6#�-�(���u���nfC��-�!��Z�$ަe�����@N�`�V#xz���O�׳���h~��j�]ߌ�)�M��Ȍ<��ڭ���o|.�$#9��x)�;���tz��ש�ʮzo���-���yW'(/[���������u�̆�N���`rZ�*��Z�o�~}�t7J\�E���6�[���S��#$oo��5p�h^�F�l�Hd�!�֗x7-S�Y�n^7?e�\�!����?������+��^1��[�
l�!j�Q���`�ZX�����k3�|$�MCx��IXn��N�?��_�}|+c�e��$u~�����I�b3��[������֝�ռ�H�N�J����&֩�g�R��fb��<�luw������a5��ӊ���=B�N�﹐<E.Es��UL��&4KK_v��[�!��D$k�z;8�)>PY�H{G����{�>�O����{G�����[��\}|h��j�.K"
�9�h�J��ӑq�·wh5u*ԝ�Cn��Rar����a�N���:K{�X��+P�IQ�!�rԖ�↰��P���b.�6V�5���=�`ȱ��$E�p;�jf���n�ц�[�q!4����.7��V'cT�xe+�q/���b=�[�L�����,<�n�F��rG
݂������xs�� ���i����W'��N��˸�`�ke�f�����~��=�� �++�wsU��,��j�V`�3?7jH��W&��5Dv5��sP��p���p��ۂHFV��!��E$��r�Wqo'Z)gn����L��h�N�&�B	�^msDn���W1��	�Xqݐ�v.ʈ��^��uař8�o$�9�93����+7�
�%�y�M�ϲ���s�(.�y��T�>ɥ�]�ԩt�E-w[I��r��\���91�ӕ4�u1r����2C���V:��йDEB�M��1��5{�h�ms��v�GVj�>ͳN�N�_#���njmI���u��K��R�xr�=AR(���:Xy=ڲ�F�客	�#d뮲f��
r�K��3d���Z�+q����1&�U���Ɨ8r�XT37DT�V��	�(�/W�h�y�dC�[���ok�˴����
ė�8�M۠���i)�.m�w7i3�S���9���P��D���Mn�vPq�X콦nCÒJ�yzR���{���R�1P���/Dj��S)��DT)�G']={��B{vlQޔG
��(���3xЫ����OG+,EB�>�����b^��P'��I{�e�#�e���-%n�T�n��R[w{p������8R�lu9�vpT����A��"GR��ͩ��o��*G-X���1�ϸk��R�ԝ��Je/�gj�veK�t�g� n��©�Ǘ�J��Jٛ����>\�r�Lq�jEs�gH1�o]�4fH!j�eZ̥�����wMZ�]�co3�u�5�:�vlt7�I��Z���]4���*�W�T[�{G���NZ�|���t"t�vݧ|�&��, e,�
d�Vi;�]�2�� �P^uG��6�!)e�Z�C��\��P\0�\.4���7Eg+i9�/������W�s��Ň��W3��ʶa��s�.���h�V��+nJ�x�_R��R\v�U�5�fͧ&����E�A}մ��#�l�+
�{ԅx���a��;��G;�*�f�'X�a��WX�"��Y�'hb��'����d9mtyj
��=��Y�&��7��Z�)JU���dwQ�*���5��[r���:�<� �C�TK'����k; ����}Ҟ�*�=��Ҧ���L�/��V�^�W�h���ˎܮ���l��%9��ձ�W��c���t�L�X�T�7F�y��K�z�6�KD��;�u�b���t�q��[c/��Pvͨ3.X	��m��;n���o��GR���s2p�lIQMD�L�[��#0�g���s��A�A�
L�e8�)�0U�Q$������x�ց9m8�/��Y.�9���L�A=Ԝ����$ŒW�ȥ1y�T!�����o[��"��<#�gR��¹FִLBw�p��b'�
�Q�s�9W'Gt
z�̢>�ENd�D��Qe�TZ��}>��8db׻����ebc+Ot�>��� w���-�{�^�sԎdb�Dy�jki�ۺhҪ	҃s�,�'H��ê�K<��fC��{���De��;����u�j��r2D��'�y��z���DL(=���ܦ]n^8��qb��Ҥ�:�l/��纥�����rB�#=wRHNJ��3��DT�{��.iz4�M�j}hU�4�ش+B�B/��u'2�0��K3<��3R�!8h��aʳ�ꨤ�r�Iz���3��\�3���sxU���o/G����z�ݮ5U%� (�����ɾ!�ԭ��$��J�"��8QY�������{F�-L�ի�gR���>Kֶ��$L/!���2N�Y��8�/�K�1��{ٰ���[��F�V�i%Zj��mh�3��ǭ͵%va�����3��uI�{�w�5ۋJ���̥Ju;a�O]��!�����Ǳ�9���Ki��,���F���,����ƌ�oX���6;b�9kv5��(t�Ht6�Tkn�A�{���
T�fD0��16V
yb�/��NH�c�z<3��Hc���׽m�x=hL����.q�)���aSf��\fT�i1%�T�L�4�l�<f�ڽ0��h��,
�=�s�@;ޏ���"�٭Q�4��cS^�"v��va�ܜ���Oj�,2^F�i�n#M�{�nU!﩮�G�b���WY��:y�C�d����Aͳ�h�T���l�]�n���1c���~e���{�du��i���s�x'V)�7w^NU�k���ظE��{u3���o竱��$�&�Hen/�jz���ɽ�V��z�a"�'�N�%����#:w���r}~�)�q�n��q�j�z`���5:���3ky��eӝX8��^��'�ި�
r�Q����3�\naU�����纋��Θ��~�#nZ�KUb��y��.�p��b�$+�ח�-ٷ[w6k>�w��R��k����]�k�6q6�T�W���4����=�E���@;Ԛ'z��0:��X���G�9*���n�e��UG/&f�z�u�]aB�]]��3�tXfz}���h[Pkd�w��j��W>��	siB+t��k�M�#a��9�������؞i�ƽ��M����\�����5� m=H��jk���/�1����xj�'�53�1i��A�7&<65m�ŗ�z��s왝�l1�d�ɳ{6�ٹ+*s6mLz��c�]��4��b���N�'����o^����Z��������w�S�Rb5���"1�,��n�%<���+�� �����};��Υ�FX�)�lR0_=	3�+�<��K^�~��ɝ������h׾;��:mb��Vz�U$�y6=4��k�P��O	TS�c}S���"���)$k�Yg\ڎ]g�q��*5��~\��9#��f��)���I��jt���N��.obV-=�����4�P�/,��W��j�5�����f��Ŵ��7�j�ʦke#((�z/�2M-��^�X���|��8d+�.��������)����m��k�߸��;�u�ˇ������w����;\v�D�ĖW�P*�J��y�)n�ˆ�������=2��K�j���d�̀�P��|(����Ҳ��d��&�����{R��՝������Tx��[n�-4אST��:��"i�#�ާ8֗���u��/��6N���R~�ޞ�wj[1�k�!l��=nw��(t5����cV�"*��b�c+v��UהM'���<-�Gx�t���+\Y4�'�a׃�4�p�h�v���O�ty�Ԏ?�=65�!D#}���>�9�����œ>̝�Q�|KйJJ��o�o���e�;܅c��ps�l�E�9�K�_ #W;�9��;�����[Υnքo�|�~6D^���;s�{�  ��1�k��b�8��|y��)�
�N�,ik}"��)����c!����V"[����V�i�k�\�U�(ʸ2uv�]��V�a>�>�Sɧn"����v��V�w97�\@L�K�9�w�d8����h�E�������߫�^�Ѣ��t���J��9݊��w�.ŧ�V!2�D�c����}~|>����q�{ܘ`�^rؘ+����lh0��rr�{�Z��ŧ0�6P����rڽڴě����0$��}0���]	nl>MoH�f�{�Kg�u��v��:��O������.�omZڭB�v�ϟ��V��ή��Nj|���iM�R �XIP�u2��ΧH��bGY���D����M*���܈��r9p���j�c��Z�a~R��FD�C���~�k��mʥ���KD�ŬKoHX���{�=q���W�QyO`Ԗ����uH������8�����]��@}��.�쳸u�e��9+M����-�WS&���O��6�O���C�@P��tl�������9��a ����wr9U���.n�Y5_�����T��j�����)�e]f�vB�th�92�"��Y�3N"�����wgu��ɭѮ�t��ˊ�]Z�Gw3|h�՞tvt��A��X��-��6�ݛl�'��}Ws_��+��E�|��Y�J<um�C�9]:�ƶq�{�x2�3����4�?a +��n�+�g6�����I���*m�,]^G�{i�YP��5��v��J&QG��&o�����xѡ�Y�޿(��D�;$V�E�u�z�u��'��V�	T=�v�ʰEţq�7�"�
�,��XF�3���ȸ%Qۛ��)<V]C�cݕ-�0^U>�c�����j�����$n��y�z������/IJ���<�ϫ�gY�m%�V�J]!��c�q�>�n-���,.��l+�V�� .ɞ��.Mt�ܝl�!�9T�ĶI����-�~4�L���7;�y���-�e�k<w�U�jE�;�ps��_O� �@�l��Mɓ�Ӑs����v�>wABV���>�}su�I%��o4���3w����%m�6�=�]�Jw�Q��Ws���_&��Ru4U�G�P~��
?�e��fe�y��ړ�l-z�0Zw:��t���yD��A1�I���9��˴I���W�*���w��{]v:Z\\ݜs�,�9G�V��+X�tZ��it��ZuҼ
�<���`};iv��]6B�V�giv۹%�I��t��)퇙��=��]�����n<�{�Q�w��>f��R�\����;��Q���ܪ^����l������7��>��}n�`�I�[�͎��!O��v8'�Y�Kq�(-��Z�St��f7��3q��j��}�G������M�*��}Xb�g��2��>̊v�s�en����A7�	z��g
����=^n���T{�:U��[P�rcoU]�^͖y��uo Q`��!P�&���ݰ>9ת��p��Re�s��ݮ�'���;��k.�tG�S�I�h�F�
�lN��.n#�������x�};A�.IY�3?�vavޱ���Pݺ�.�J�I�mG��f�7������l�R�:�6_C��_����䔾������F���z҄����g%ro��OH�縵�_y����Ps�*Գ:V��j{F�t2�����5{��7z��	v �W��8e�D�J�]�n�8�%FP'��G<�J&V�����%��U����P�[��	��Bfq��{���"�����4���\��ھ�q0쉜�(��p�8�ٳ"��(ٳ��"�7�2��Z���|7(���Z}5?(^{1���s߀�9����XU�z�nX:�	�ݝ�M��z�߆!��~�����ٕ�<}xў^��6&���O�e��ڼ]��Dr*�1��K.ߢj�$GmM�ʮ�������}ή�O���;'�ٮ*���?���	_�][U�[լc�l�2���CJ#'HY%[4#L��2��z��L�nA��Ԑ�7_u��QYK��A<��)E��l����KYi�/��M�td�b����>{�p�<`�K*��d���}[cz��[�	���w^�9����;�g�$�v�������*�^r]yۢe�'\n���ӗ;�v�x�L�����s)1V�A�4�0SW
�Y�6 �����o�x��9����#�wW��H7kyU�̝�7eBv��خ��O-eY��P���_�*=z��O�g�=�����#���ܩ��L��o{�p.��6��[$]�i���͈�N�:mu?��7(��S\	�a��� ��e���im!�;�V�6���fl�g��`�f,��{c\�jٯ��&��U����7�vn}�E�m�ό��E��h�r9Ƭ����� �]ky��:W�zE�Hܿa�����J���W�ІnI�a�zn66ʪ�%��$T�.���Z�8�K�Br��s3��~r�ezl�6�k�ِ���_�M�*��uKv��ߞw�ŋ�wj�U�^�\�燎P-���y��!���8����:{p��4�|�hOo[L�Z�u�t��&ۤw�ǜ`�a���WH��Q3�!���ai�o���!�I��h�Ĩ�!�<0�vI�F_ ���z����ʺmltݥ��o�=��ɴj����>�v�,r6qy����]k�;�����s�R"mm���Q[ɺ|R��~P���՚�Ȉ��ͦe�5�czSG3��0���5�u�/��qy�FJϗϫ���ϿM�d���[��F��ӛ͛�b]� #$på+<�f�4%s�!?������=��N�®��|���^|�<N-`�vdd�*� �N�\�-rؓ��͝��%���5d�����ָ����M����t�13��x���]*Uts�K��V���h�C^σ��15/f�GL	�����>�� +\뽞,)��W��8��;2�3�m%�ܙ�s�x&;y���o#o7u�0��z[2�$����Vլª�ݲ��]>k�J1�6TU2��]Ҧ�,���MA�x��@b=�vFl�s���E�*�Ww<�c^�=�������i����I�n��c={�:�l���#!�%K:��\��0W���f�+e'�����ͣ6�u�j4�-uY��7��iq-4-܊��or��D�Tn`eGp��_�"�������}�Q��Q>�<�:V&�i힪�8ID���f�ޏ�Zw1��Q:�o䷲c �t�Gph=���Z�{���ǵ�g���ٵ]^��̛�mPF�א��X6�n������r+�������z��]��PgR��v:>�F|JkV�����]��uWer��󻴴�%���;�ܝÎR�c��.*�>S���k�ir�C�G��g~sE�>���ξQ�a\Q��y%��/�hfj�SR���3��Is��t���Ŧcޛ�wk���Vs����B�a0]�r��Yy�V𛣘���o�{�� n�Ӧ�Q��5b셗��;:�i]¢��s���A�[���Sbɑ��u����	�J��E��[o������ft�#��C4@gf��N�Pp؊*}b���7�=��m��cO�d���gө�Gz�Nc��~g��j�`������Ws0�l)�v��,�8{����Yн�F��׊W��#mr6[����1\�GuB	��}�̔�:�������_x����U?t���_{�:E�ʐ������!�m)�^3�.���(w ���{M��V+�����*��[���{F�o:;jp���Z.x��~؎=Ж��y�u�V��{M��9�Z*/~X�]�d�纖z��cR6Z��pQ�<#R���J�u�b�jdS�[N�\�FI&�tǩ�d�=�L��j��v��x8�����}>�O����{G������T���P|�����巽�.NB�V��x�-�p��E��Xw�y���16�t��r�=6�h\�iT�Ao٦�l`�pɹOuh�:d�N�}̩�]ά���������^Kg�e�bI�p�BJ7ZrpZ�L���)f���m��k
�"�+r[ي\����h�=�`��u�Y�t�QX��4B��&�ePP�-^k�Y��p`{*_�]�ԝJݩ�Z)m�NV��9G�lGx�����[�#8�2�����6�=͝�k��2��*뇞m�N93@,���Xͽn>��j�/�n�rY�!}�:�V�\��)�������S��B�X���w��Z�..�.[�w�EvJ�خ���Z�(��bY�tp��kN��|�'1���ţ+%I΀*��;/ p3�\hS+h���
m�G#SC)�s�V�F_Y於�s� 8b;N��o��S�r��A��V�e9��.H-�y��O5��G���Qz7��YZ��X�������P�Qx#z�i�8s �����Q`�aP9�ʝr�5)��W��ԟt��]��;��6��u���,�[AK���M�ed��ʎpy̳7<��HL�\��zSS��i��Zv`�7�ۄ!���f����;[p��.;��<ư�/�Y7So^%�[ص�W������L��{��,�\�J`顐CdDY�vj�������@�@�Y�����繵�FB�s����dG���w�U�V�F#4�f�_KvGVP(�9qm���o��� ��3�gb��k�fU��Dt` �>��B���Ε[WǺWf�4�J���v��ͭ��bÝQ"�K�J�&���;s��j�ˏ���=Fj�fE5��sH͙��	�Q��oD;!os7
e���{��:5�k`ze= I�r����7\�u���cx�R�I����U�Uԫ]�0�f-�����!�q�{�悌�*F�)��w�i��6���&�����@����
ucCj�MBg���j]���0���IA��F�m���ҠɓU�]4��{}�۸
5�	����j����%�0�
�j�,%z�_(튼�¯�!#\EBv�v%���v�:�v�)R��B�*wD���jV�*[��u�g`̉��Zr�y�e�����q=9-T_)��[�r�<�)�1|�Z������mW9[�5�b��K��z��4 ��-f� �s�s����U�}Q�KX�3w+h�BOô9�֚���t�j���!��3Q|���-���\���$�ظw3\˳=��Ƶ�9=.���ԩZ[7W$���Mu���}��5�ȡ�����mM�����	��w�/C�w��O(�q8 ������(0�*�[���Bt���G/��L�=Z޻
>kE2���C(g����7�;.��J\�].��aL@؇�J���=#�PS�Q�?^��E�G���~�aj%�~է��G��Ⲫ��L�D%����"(�w9�f}�]+�ʙ<=3۹�j�4��&y��[4B��&<��Ԓ#L���Je����A�A9�Hhk������7w]ݥ��˹��ϊ��z�f/^�{�a�NNS�����NN���D�eHW�	�-nM�=/�N�{��J��9��U
2Z*�V�{�xL�	�{��^n�q+�ZG��{��8%�IB�N�TZ����NfBFnIR��y��=-�c����u����y̷>w2��L%�7'<�s=>�z\�����U��`$x�*�f	:��y�\����N�8S�J�JeE���������r�*�L^�����r�'^K����i�����.mε{��;��[3�r��uu'w�J\���S�.IA��W�A�0y���]���-&�ܭy��v��������$�A?~��H��ɘ��0��ݸt_;OX��|�<y�1Kz;:�+������rq�زe��z�0�냤�YCkk�%��P���X�s��
��48쫪����/7��VOrJ���T��99{`5�<�����S
*"�Rf�V1��E��KvVx���Xh���T��:�}q��sU}�+��s9�`�{2+{�}֔*����uZ!���
��TKcDX���f&J��=f��V��{p�;V�����J�[��Ԃgg�[P�kk�aW�xl�ӭ�!�ML��GY��cN�w-�'�h�lEZ|1���a��ٸ�p30�/����>��A�����>Ű�q��":Pmq����ˈ����^�trj��d�B��s?�fU�˒2@*㞮�Mk�e<�S�0�:��״� ^�	kJ,i��a�HN��K�aR��Oɛ�Fz���7��x^n�֤�pi$�f�#L��(��bna�����7�[.���T8��}����\Bz�$��Oq�T˕;��Q�j����`_Uŕ�����~}\&�˂�큑Lm��E�����������^�uj�"]�]��o8���[�JEբ���[����b�ft�\&Qb���:�
�EMc��e^Ӱ�S"��F�a�M�#���C*h��}zC�୎�h���{�WBu@��+�S�9�J�X�i�w�Բw4K��Wy�4����57v�5�U 1�����Op��$K���������3z��sN�YD�U+s-��N��W�����*�NvB�n�����g"�l�ݘx��9X����W� �Զc�pB���Î����lyDT�H����d��C��a���!_f�ݫe�O�/��m��"�9w>m��:��^�R.1_;]o)�t�%�\T�F�
���D9W��*R��70��I��å A�"�cm*�|Kύ�TWq-���'�5Fa��є�:0M�L5��W�+��wlB �o/V�+V�U�m�{N6�f�d؜��N��~��{>:��=���� 2\���Uzzx���u^�(�����zZ��2����s쩝�m�;�.2�ۚ Wuyv򾟋m�L^Z���joMd�2qԔ넡ZK�
�4��9a��E;zc��U���1����yb�u��v�,T��P����G�����'Tp��pT�����nW&�8廧W��n��]����f�p��Y5b}ĉw+A|6�E���Z��` eZ������l�Β��v|�s+ǮZF��1'�;��� ��o����^NE��
�tA�F+9w�?q~�cC���'m+�����w�VݖM���j��-t�袦&�װd��h���RC;�lAT�3�lb30�_bU�&r��pN�>��T��]]^�w�%�DfތǊ�sp�]�+q*��2i�zk'��l������^�X�C����t��#P�k�4^[9�O1��ϻ�o��n��g�r�uxGS\�U�=���-EwzLE=ͱ-�����>\��Y�UM��2��]-~b�+�:��x�.�]��k�,�`����S��풀D�:���r���i9���u����e��MdAݑdm�&�H��T��[�	]>Vsm@h8���q��n��wF
|r�Ǚ��!v��.՛�Q4���N��n���rq��ˉ_`zt>�u�=k�P�݃mW�iôhn�ռ��5�*�Tĵ�g^�v�8���XN:[����c����287;4�h�L^R��K�5����34vZ9�!��'Q���Ǔ��N-ٔ엡��R�ڏIW�v���_�eJ���.���2Djޯ{vL�W|y�E�[�Ј�;<.�F�3���_��ιW_e��5A�׈�;��N��S_�ɹ��|i�W�^����s�x�}�ubG��2n4U�� o�����Dg���}�֎1��1E�V9j��\����s	��6�}Ŷ��j�g{��׳lnN�g�]�!�M)��:�-�m ��c�xfa��}z�C�[칢k4��N4jcgf}r�ӫc���zZ���x��D�Hd��eGmBo�{���Ph�}.��ĉK�'�]�o3x�J|�Rz,��4]_�YYDa�7���+m��g�EwT$�D٪�秡0�G^Z��NDf��>��r#4"��L�z�O�[>W�Ly뒙�n�"�o*�\�u���d��ٹ�VB�Q�K'(jƋ[q*i̊�����x`N����)պ`�W{��~&Y��7�W;��˟qٝ��Yf�tB��]�-3G:��r��ms�j��l�F�|*.��!���ؔo2}	���칼c�4�D�)@�j����O��O�jz���ʛP�������`
�n����.�JLi\&�r
!@��jřɼf�y����S�����27�e{�>W�'WXY�!e���v����G��6p����4{0+�����O�XuߎwJ]eJ�7 ���5Y~3�y��M\b&��"^�2=^�f����W#:�uy�-P֭�DMHm������%��YS�c��)���3pW:�s��H)�_�����[Z���L{�X�4�{]���PX�� �xW�u)���O��s���T�3�K��.�+�>���+:��n��I��/.jVa�}iޏ)��nt�"�*]��0�5�k�7NEˮȮ�C�3^�9��ҤL�{c:�y,-��x��Qz�+�.�W�|�0o�iu��(�Y��J|�twr�bx������b;׉�y�����ͽF?<��#6�)����q���}vcqi��Nh1�(0~
�f�jm�<���_q:������qA�+�eY�'��4��v3̡�x��ISh]���ꋻ�t\Ssy�U������z.����`�9��*����%�]���b�B���|�L���r�GbKr.~����9�����G�a
G����go#{�3w�5Pډ���>pqR@�Οm��9��[�H�e�ؙ�W?O5)p������=X��gU{�|�7��^d���y�!d�l�4�GU��O
�d�]h���S��y�*}�����J�m?G����
)��+e��{B��`�nun�t���3�j[.|��2�\il8���
+%i��K?Tn?!%��i�r����[<Lz|�q�5n��\�����f�2.Z���(��۽&*Emv��_*��Y�@�x�[-��ƚk�4z+�\�n<��q*L��9Gw��FE���\�/${�Y�����W�'v������w�;\���l�nh�=�no$U���~J=q�=S�<�feu�Ƕ����K��cNu���ӖC��5O��;]o)Ҹ`�(�m����d�i�c&"���2V鼱kqv�cu`��TT�}��4rKxִ�8�ؙTk�n�����׼nӀ::2X|�Ϳ�:&�JĞ�V�ӽ�R�<2�����8^��v\x�P��sF��5�KT�y`F��XN�����7):َ�v�_Y8�� �')�H��#������z_��뎏u�Y�K�r�[��Q}�7�q�6�ۗ���sMC}���3�08k���􈏑��W��XF�E9`ڋ��ܼ}�+/_I�W@%|u��3��6�����{V~9�ޡݣt�7�w9�3��d�a�'V���	���1��m��ՑP[}�;1�Fb�r��**�:�7t��y ��H�Ӵ�C�`d6c-8:a��͹���ob%�O�:��bޱ�[���x�b �T�9[��H3ҔF)\�R�Z��|#�L>�17ʆp.��4��R>�,C����y!N����Y�v7�{ ŝ�-�{=ʈ���Xkؼ3����}O~-��N�C��+2.�'R����� �zK�}��މ�/F���8�zj��l�nT���6>�nj�0�{�F9�Q�jn~������df$��q����3:aA�/7��k��$����3��j���$��хӜ��W��йن���;O6�-C��EG���)M ��B>�$�V6�_K��r; 4��1���ʌ��t{J�b��ù�9���Jnܐ���`�����MS�W�E��W-����*�[-�e��t,3=������q�A�S�zo�WDЎ��q�e]���\V�ONtH�M�Su��y�5P�e�͏z��ylQ6���)�K�i�t��e��L_��h�Eh�� �[����k�]���h��x�EL�T�F��@Mk����T�ȸ3Y��P)fQ���jC�@wX��� �����]X�'��m���DEݻ���^X�T���EP��^@j��%��Fc�t�K����V��Wc��
���IrZ��$gC�p�̓I/%P��s��9	o=��M�t���ξ��S��a�Ȩ�Y��򚑻+98�����p���LZ�����/7b�oM�����t��N��$��3����f�׳��F�����]���3YH�}Kg���k,|0y�:��Ӥ�u�P+���9Ұ��B)4�f,;b�����xk��eWcNr:3v��%5p�(�lA��c��㶸�*\s�)�Sx�#6��d��#X�ҹ�o�x-!�(���㽫UknWeoV+r��HL<>���q�)�\,�p&�$ ܟu8����N�u�{@�1����r���Xs�8T��77\z6����J�뵎�mI��쁘<l���1�ey�9��EH��wec�z��)�'b�06�h���Iu��Hl�Z�)�vh=L�<`Q�"�f)76N�-�]�@��"j�S*�{+PO�^�����,Ӽ)j//�VsNm�J׳��gD�Ʃ�eXԢ���Y܂�;+����Y�)Ʒ]�M���s�5���]���T*��YK=xb�g�:Y�IWZͫ��k1��x��:%��Z�S�~}�qL��+��}W�nr�o��vzå3���&�m��x���b��9 V��9U\��㙋�=0��,d�����9�`�)H���ޤ!�6�wt7vmٵ^'vA':���|:s�q���-mg/؋4�M��v�WЃ��Q����J ��1/o8v�����L*��r���ۻ��Y�ؿd@#~|�t��롋����!;;�1��"�=�*��,�彫�#7��>�Mauՙ�[��|L�����w��%�wY�<-+��7֪:��ʽ���tӸF��r�[�j+=St����x��z�s�'�;9�ͺ9�2���14�i�����}2)�s������ ���h���le�B��ƽ����q�DjU3���z��X;~s"��9ۏ��TW7p��xB�[^y�&���9�b���̮��ޮ�N�&�`�}J�m�E��6�M�2{_�-���Mz5'� �I�s�-���]o�NV���w��U�nTy& �]�YD��}g�&9�9�+�C�^�O� �wsJ���.�W�R�Psl���'�Bƙ�����'Yߺ�c.�ӵ�&��E �Bǡ�C����#3�FH�H(fFY<�Rc���q
"����K2�N��=>[���oWWg�s�F�	�$FHJ.\&��sY9~�ڌ��i���$���Gl髝1Q01%�z�V��)a��N���5�� �d���P�j�Sjk�cA�D�P-oxz��oO�������}>>^�?��>�ܓ�~9�W�;/�i���N���u��}��ʼ\���Rɴ��($1 g\5������N��3��d|n���{���G*�u��#�����&QŖy�J�ʌ���Ɂ��g\��¤��3d���~8�}���k�r��r�[D�4���M�yO�,���e
J���W5�C�[���p�a���uH�n+�˹�]�j���MZ�/r�Wc��{&P��E��YYUۄ��@�mIo���v�@��J�ӌʲO�h;�}y�ES��󨆓o)
/v�S4F�#�Qv�qը��QKAΫ�s%Hr��8v�����D��������Z�c<�gcVyc�y}����nN�Y\*l��h���X�Ϸ^P#6�,$�U���C�!<���a�VlO]�H���t�9[�S3�]������Z?*���4�yV2ӏj`b���<��{+��e-�;�EѾ�.gE�x*�*�j����یX��%�Y�������)��[ӕm�pC:�:���t0��#���΄�[���%н����W�N���4��"�f�j�N�fLׇc	R4#�Ig
U�T��%StA|h)��-:x|�f��-]�t�(Ȍ��*�:ZU�i�vD]l�"V���Jɂ�&��Vx���`1��4��2a$#PS�1Q�J�&�c;���7�8��Ֆ{uRi�a`��J>{�c���[Sy��Kw�ЊMn�
=�u#C�0���<ӱ3�f�r9*j����kr�ƿ �j�c�y4C�+�v��6���)��눚�[ա�j!7��t��G��	LT>%;��!w�#�/-d��[_E�dN����F{�+c�j���C2h���	Zf6�ou�8������xm]��
�x�^�c��v��j��sSۧ��V�#�����ZS�wڹ��n�61<�{)�ގ�wE�m���&��ӝ#����c����ؑ{b�B���Us"���I����j3g^&���H-MnH�r=ؕMo�<&� �S�rc�}��\��a�A��S�vH���ݖ��K�}W[�{Ǖ�{��f�_ȫ�\����A�&ݬ���bۭ}ӳX*X	e�{}��t/U��R{�
�u�q��7X�����nt�k��1N9bu5�XEfl�	��/^�Mn��P
*:L��Sd��z�1�7�����_��#1�gD��*���rٌV�/�ը� �����lM���έ�������2�_r�y$I�[*n詎��m&��FW\U+�,u�j��[N�s���ӎU�rH3��Z��+0�5��a�t�yn�Sc�E|�(�j Mr��.Z�^gS2����2��D뫯�\9cGo)ɓ����>iv9�Hr�l��5��M�2�ՠ���Φ�qo-�0���-���:.q�ml��L���Z�a�D�e�_c��Dc�����#dB��A�1��<���R}GqP�.��P�*GQκ�X��͸�[5��N�W�mԯT�Z&*fhYnnʰ���'e;41sr�mw]wtB.尽ѕyUy�8Q(�E;���Ԋ�0�n���TZ���
����uq���SCNx���^F��)��Owtډf�
�*TH��2�wWHr��P�^s���Z"#�ȏ��EZ�Hr��	�/\�#S�[]XM̽f�'�z)4.+��ϝ�g"�s�*.]0н����H"*��s��ĩ@׮�^�W���G�7'"���҂���{*+�E�䖚!Z���h�I���E��C�X�M�y�^�G�^��I��С�[�+hX���.���ww�]z����G�>�z�g��KW�k�V�fJ�IS�۳�e*h��E�
��k���fUG���xQ�K��A�縴7�C�θ�����y���zz9:^�O!zʕT��h�m��ܩ$*�B��Ms��5��}��瑃�ᦜ�����ŁqΠ�nK��ngqj*y)�F��g�z{SO�;���Hk?]4��~I�J�A�����n~Omx�Q۬a�<�}T
ǫe��.4�\�)�C�,�������S� ��O5��+��ٛ�۵����`5Na+�m�#�{��U�T� w|�.�^��ᚗo��((9�����4���w�=��5x=�����~+�.SW����=w���q�늷�ǝBYy��vlƇy^�2a�h]��n*VC[�����9�'�,�Wm��G<Mn�3;,�v�
�l��1�y��d�e��;W>��1��WU�ð�Nk[�^�qzՠ52(��}'Z�{����W?j;�7����b&��yn3�=g��i;�O+�vĩ��m�G{Lᷙ�S��D؜�e���\Y뵫�����0�ὄњ2ƃ�/;���2���ȭ'�C�5��T���
F@�1�q��{֟lr�����=S��Vg+�y�+����<����x���y����l�ջS�۝y$,լ|��:��ٛ�v��FB�����ƞ��	��,�ZÝ��=S�����NfYf��N�aj�=�¬�:��G�'*�Gncr����}����kO�f}|��2�0����R
W��fR�C�թԩw2i��3,1����ݩ��KCY�=�"&����p�4���W�1���3;�p�ng9�Ѽ��j�h�4��͹�b�^�?@���4LLޢi�c�T����	��f:�UGS���n���9Х篪�u��Oe�nb��_]�����䒰�sk�s%+�c��F�:�|��|�,y��i���z;p�˗>B�9����Z��e]��z��5��o�Ce���Z�f��
�σ��-��Δ�=�7bꝇh�<Ӷ��l���*Ks��igq/�d�֬.�o$ݷp��,�9ܛX��y����ۺA6�ۊ�s���	uC����s/�ط��np��No��ۛr�'��	,[��%m��k3��B�m�XW@�q~z4�����ʍ2>ѱE�� ��%f���7�-���U�<���^w�������3fj�,m��}aƂ�!�\��X���o3]�퍇���='f�Q�p�W֝����2��(� �ڱ-́�5{Rg9��wZ�yU��`O��9�Fa�4��$VyE�P7o���&s����3�ue��ykSl���^�d)����y{-R7�S\C�Ko�o��2@�Z��p���Lx���y>7��w~"��sC2�U��4�Cz����;����Eɏl,�۫	7-��c�:g)]�L�����vѽ!���e��� ቀ�f`+2,tk�P�����~�����n�Bnw~�������u,���wW�E�6.z��Dt@��2)��hGKms�`�B���v��c6�̇��SɵY�*�o�t���w�&�=w1r�!��\b�h��e l��#���UQU�T�[�=[e��͊��u�f���
Gi,��}E�t���ta͇���z4W�n�,А}��Mpj�Qq���f�
��Cv�ܚ���h�Dxt�{&-V:����g��ec�+>���E����Gc;��}&�]��-.�;3�(hQۦ��w��n��q�w��3�wה�w�J�+���a��Ҭ�����B b��u^��ns{��-�K��8*�H#˯cq1��+X���.�sf�J_�5�2�u�-Ev�rδ�܊b��M����޺l�V�?G�AW�7�*_7ƚ����]��'F�������f���ݟ1�����%Y*�'r|�7�y����|���Jj�v����R�9'h�&�ܸ��Vu)Ҿ� ��+�^T�h���M��m�z�Z�gH�*�+�]�'r
�>O�h?e����M��U�0ɸ�v���"��yQT��ީ���2+W<��
��Ya�F&~����wRniY��﫿�'�Q�]�|J#tlf����G%�f	���W�����=��~3�,x��r��̣������gyv~���7�pEd�5[��g*���Y�Da�zy��Y���}p˹�
�h�q�K�b�m̈́MM���=��u-�Z8� �<��vy�;&3�m����9ϻ�Gk1����-�H����N��4�%[ɦQ{,����[F���v�92�yzo���;��L����D��IJ�t�eV��Rt�m-K^N����z���&;���Y>f�_�9��}�;�W͹g¦+{���M�j��e���Ƙ�"�Z��pm��)ޫ�����ݧ5�dΦ�Ǥ���F+����^dč��W��h���b_4 c�Ul�U��ދ���H|dD�|���!d��0�sa鼌E�	�w�z�2*HζS���WS:�A�T��v=:i�_ؒά\.xd�Ñf�z6�ĵ�]ј�+cշ�0��)���`�3�g]G0�1�n���Ný9zC�7]���r��Y^fU%�x�'�K5��.�Z/��l��n\������lr5�0��w{�k$ݭ���$���j����l\4�8哧���w�e>�l�����m�1�P@A�Жǂ���O�ՂIzy������v'�9Y��؇m����Q���ܳ�W�O(����8 Y���[,�芖��{$:m�F���a�4.6�*�Y%�]
,i(^t�X�:��T��@'����jl�v38k�6D!�>r�wb���d��n�x={�A�Ib��
����QP_�^��G�x��i�IX�I����b�y���'Z�0�1GX��XQ�3M���4(��(���tt�-u!үI@�[�×���v��i���?o��������]�ݙ���V5��_
��������c{�H�n�7�ֶ���>{|WW�!2�5�e��˶Y�.���R������YV��Dm��n���q�t�;
���-�u=Q�v�������R;WP/w�{)���p��R�1�w,��8>�{V�DN�'�{>�T
�f#]�t���#���a�o�嵰�)��:g��C��|�+���}5��!Y�|�f]�|�-�Pn���,�X�Ոz��*ȱ'�X&�oSj�<lx5���S]U�=�x[�R���GD_N1'O0�"���Mj�[��l�i���zO���Q�+�eӌ}�����KeE��P�!<��&b�a�U�㥶 j�k��=-}��a�6��5ק�.��m�R��)PT��U�W�T{[�aS+!,��ǯo�*4�?�{�#kV��D�t.�ߒ'����Xc�ː���ͻ����^�A�:��(/�dv����I��
R3+#X��ц��2#�s�7��z�B�}�%�#mYKvs�*u�+�����d���ɝ�.�)H0�oI6�1�#W�䙷&6:B��pv��bo����r7��� ��k_�$;d4(v ��>�P$�X�!��{4MX,�<��ސ���͓�Kg��q��Z�#,a(B�Ck��L��{��I�FT+uN�g0��t�9��5o=ޡC�h�E��.��n"�9lM�?��$EfbZ�r��N�[�(�T�46����d�5l��l�O>��9Ļ���9V��0�Ix��9�뎩	w%l��m�����xю&b�S����˽�+`m��Rx�s on�H���6υ��G;DFE��cΓ�3�>����+�|�?��;�ⴵ멡.��:�3ٓ���v�(��e�lMz�>�XbYo��@ەރ�'VW��[��ׄ��Z�Boh����i73̠�oS9�jE�홀�Ϭ_F��}V����xM����E[����{��D䆾�?'��<��q���x�k��E�a���(�O17O�W}�[-!���C�d�ه���� lw&7"2
~e	�}���+s�9��f ��3tƷ
k2�_���v��5�ނy��Y���Tɝ�tG�7�-:���U���u�O,�_<��WZV��n��	���
eQ.y�)fW�TNuc���8��Xͣ+Oj�y9�GV�c�(ҏk(�|���C6M�p�6��ս�')�y-0����7�\#{;����YqWs31E!��|뤗�'�����7}F·�c���Oa���Q������^+'+V1˭���玸�Y'���LS�-�|�m ���W$���3��r	�*�x�i�t��C���7�s[M1&�Y�^����j��v�Z�$����q(�^k�E�貲{1��b�g2�=�b�n�y&�dH�eC�O%���U�4*�'RЮs=E:��M1��ʣ�|��]d�\���5�r��KF�c��뛪ł���Y�JFhx�9qgq�z��R�ו3\���[���ƛ[��$����"��?FR~�{��FA1�Y/�z��/���7�Ɠ����u�7��&ً����>� �P�ݼS��笨TWu�U�uP���b�$D�b[dp	���E1��Ȉ�b6���W���<yJn�6�-�Qδ�?�,wZR?v���u �9�r�s,_<Yc����Y���J�j�	��k�s��N�ݭ#;;6!9�#�ݖ��`ɯ��6��G:�f�kHnbCNLl9�r�A.�ݽ|­�S1+۷7�G a�iJ�nEn�R��RV�c���bo�ͮ���~������>���`���ؘ#�T�Q=
2ߢ�k�:���Kqua�s�3;$�c=�p���F#�p�[S~��{�"�w��{���o��{O�'����v���!�_�.���g|b�9 BK�`���8�#����3�R�4˚Y�������ޭr���"A�~/��8�i�s�+���y���D������K:�{��]��`��f ����ޗ��5�O���MԁRo�~ѷ�'�m��Oun��#E6�}#v�H&��t��zCTu_�Lz�y��H��嚵�Ϲw�p�ʂ�Z����Y2[<{S.vƣ��ҥ��~���3�u��^��A�g�J�7$в�+�fU%�l�C��:&+�û���_���7��m�>섖��i�	q'"�����a 4{��E�������}�͝uR�6���1�3��T�Jz�F>Z&��_:Z;�>^�U�]�ko�`��+.����Fh�������I����έ&�Z�*�o�Sr���2�(��@dy��\l�\k5%[R�FIB�[j
��<SlkTd���c-yֵϴ-��[|/�WKrE3R�Gb�"������3>�3H��j~[ִ^��S���tc����.Jf�G�p����4:��ݑ���SԚ�<,�tˮu�.:6Ѫ�5x��iSF�Lȣ>��T�~�F~��8:�c��U�QS	WFN��37�6��ot�R�޺�=U=�x:ύ�g��@˨=���_*�ڬJ^b���n��X�[:{Y<��k�eL�9�~�i�7�����2Jz��͉�5�����c�2�E$�%��z}��� ���ȁ~<<�����{�G��V=Z�su�lw9�����[���)ٳQ��川�wAȜ�� �L܀ڭ������!Y���X2�ː@�}ٲ"��L6�d���=5dX(��$xf�w]��R1	�9������������60���cco�����v�`6?�������>���;�u��cA�l�� gm�;l��d�l��d� ��8 �m��l�m��l	�6��0l	��v6D�2l &L 	���&p 	��o�}�xɀ2` �op�ۍ̀ ��� � :7q�5 � d� �o�h� � &q�� � &q�{;b2 L� 	�3���1�L��c ��0	�62m�8� � &v�d6 C;3� L� d�m�; gm�ɓ gm�ɓ gm��d0 �  L��3� L��3� &q�ɱ� d6C!�d6L�gm�!�gc&q��l� &Cd2 &Cd��&Cd�l��; ��;l���l� !�gm�!�d�L�d�&v�2l��[��}��G�����`˶�v0m�C��|���?O����>�7�?�?����g�������C�������?˵�>��� �ho�?�?�1��O�&0�ȁ������3���Go���C��Ճ�� �o���~����a����������1���������[��ll���� � � "` D q�� .  � 
 L� �� � &  d0 �& `L �m�� &  ��a[gm��l� �m�& �` @v &�l�� l��!�����^?��.0aC)�S l������������xx7��}����`m�?���w���;�c�}�� ?��d�_�c��o�� 6�������n���� �o݃ m���&��~�l`���C�������`-�����>���� ��������w���<�`m���?w�?�� 6����
��}�?�?�������~��P�8������� m����?�c m�����`�.?���� 0}���?���C{��~? �����`m���E���8��<�}�������c��o�1���B�}x60cm?���?�������PVI��]������6` ���������}EQR�R�R�D )��TH�T�=�RRARJ�����H)��)$�%U)UIB��T�JQD^�TAU �U)P��QU*�J*A��QB�P�A%'֤��"J)�(*��R)ET���QwH��
�(��JJ����T�P
��R��
��!AD�T��)(Q)QB��ED�%"	%$��W�R��[`��T{�  �\W�u�ږ��+����[k
wSJku������
��l*�+��6چ��)���]�}�m�0���]V�-w8tu]�ƓE[h����H*����)T|   ���
(P��B�.(P�B�
��(P�"��
�p�PP�B�r�*����붎Z�ݪ��v���7j;��I6���K`㲢�)Ѻ�)�]�v��ۻR�*PSlUR�M��"�   �����M]��ڷ]n��ֵf��;�waѭJ虣����*����[[Y�X5.���j4�N�S�m���Ri0j��)������IH����   _iCG�[r�ږڲ��4��Z�k���gkSKL�F��y�z�Ɖ���ڦE�Ҁ�J����S۸a@�JB��[jD!
�  ���Z(*� d�o���Uf� �e*�*�6(2��(k���L	d�h�Ke!A�5$B��D�R�����  �J֥�`�)Y�XU F(�ة��P;dH5�U�3a�j�!�6elUUeKe��4m��D�Au]r*��q7�  n<h��i�_]@[m��@Ov=��)L�� *�-�V�eFQF�٥a� �`(�w kA��R�BJ�E!�"�   �  5��v� l  Q��  m��  &�  р *�X ɀ( l� � YU"*J�I�"�^   Ӛ� `�  � hD޸  `� �r�  �`��Y� i`  3U`  l�EB��)k��	UT�|   �  Z0  
��  ZK@ _C  rV  ` (р 4,Q�: j�kP  x)���* d ��a%%) @����iR4z� )� ��z�  ��2T�   I���D  �������5�U�PU�,��W#�R�f_���mAq禯' ^�����}�O�=��I�o/��!$I>@$$���r@����$�	'���$���~x�߿���񖈔�T 5ř%���ͬ��2»�ŀ)�iюⲒגѪ����^�*������.��`X��sI�.s��,6���fA�2��+�¾���ń���]�̌'����f�O6�r޼hLwzff���Ӱ�4f*�R
=IJ�r2CЩ���n��Q���%�FL!W�osZd�1̬�ؤm��ws-7W X@��x��f�3�E����)l e�c�M;Xuh��D�v31਎
�y	�C!ɸb6����V�JAڡ�dm�Z��ج���v"%��mE�U�V�h�]��Z�+���!Z�R�m�Q"�iz�I5��S��下ۣ��7kOۖ���6��j�s�� g(�f5�K�@����t�{���Nd�>D��%�A�Bq��T���Ђ@�{�Q�j��۵��A�MX7O ����L��6C5wZ����"k�	͓�&)yW�i�h�YN�5{Pe��l͹Le�(2���(6��/QZ��'I؛���6��m�b��Y��:���m�"�U�j�Vz\�r���T/w%�`��٠���,�-k[������vV�����WӬ���ǐa������V���Q�mS��)iԡMn N��j`j�- �MYO&c�p��$ {w��PA�5�X�F�n*�[8$7qiC,b��$���x!���$��۷�^�ͻn�K)"!*Νٲ�
X��H�$n�3ק8j|���fى"�kE����N]3� �����MrL&`(��we���i��55���ͳ�V���ƚ�x�ws�Uhe�ש�̈to5m��$lm)�.y�"ΰ�$�i�ux+
���b��	�yL\�Gl؈��5ub��n���cA�f�:mVn)�c����SW���mEr���b�R�LE�*��:��/FF�5Ռ5�b��K4�p\�����d�����2�̀;)M�u �-��f�O-��S�O]��"m�t[̩� �`1oJ��ͭ�3)XKT�l![�wx��
�R��y��35+CE�Ii�Al��J�ܼ.ACr�Ukr�mI�[��$4���ʻ"�4��M6s1tr%C)C����l�B�mVȕ=YcI8e�3i�k���6*�Xp���	m-�͒1�YV%+�E�[3r�cw695Y��B1������`��[(��8j	WaŔ�9Tׂ]��-�%�X-���Yb�̀�w���hn���� y���T5N;�M�x)Ї-�QP�3* .#���E�gF�א�l�Of���tA#V�m��$���X	��`j�(��ʑ�G��X�-nb��Zw�Ɠi�6u�DYB�l�T��T�ʏ.�J�b�媻d3��T�%�[MR�YmLH �[$٘�7e�	`f��OU���T��70n��TI�{���Y-ڶHu�F$��Ƒɴ�XؕK��m�n����wATͼ�4�襉ޙ$d���I��[c�������ZwB��ʼ��:�X���y�p�L"G�Dz��DI��O?�n���[Q�Y�8����fP���a��0�R���{��fU�kt�n�r9r����	�-�x�09Y+�ӽ�>TC��0����r�J	[��f-'Z�azjd씝��3-ޫ��J��R�&5�a4�[�ú����	eE�$�l����̏&�E<@���M(]%WhLdm�2w.������Ոp����Ĵ��u���Z�Z���[vƫ�w{O)�E@��؈ln21�{��j[���~�j��4E�t+NA���Ĳ䦷5�]�hMkJڍ��ܸ�L��sr�9T!�b�}�Tm�ۈ8n'�6֡�̌�ux�Y�\n�V�K`�x\�R��LVU�t;� Y�H�^Btjb�&,�*�+k�/q`�o�h1���ٻ/b�
6��΂�4M�n#�l��֪� �	MMcs-�*�q���--8 �CJG%�6bfH�;�q<x�KnkjQ�z%� �1\���+�-�5ux���L�4��Vn��F�lhO/E���W��e��C
�ͽy��d�u+IN�A늶��K^����^�t�CN�"1C"ve�(�����>.�r�D,�x�����tX�su�s.��ܬ���K���|�t��h�U�V5�E�;E�ͨpY��D �kn�ٙ
� _9���9A@���%JXD0�ʫ����ҥ���1���:-G���ӷN�8ӕ�M��(��^�C�4���m�.&��S����ڎ�+T��N��Nc[t���P���������a����Q�OӔw)d�~Pӑݼ�V�y�Ai&��N�Ӻ��Od6�X7��ziF�7�h��KPjd6�l��2k&(;��I�k	vV�7,XU �"��F.ň��6]FYҰ�C7hڳ{%*j�Pjm�KT�ɅYF���x*^��tf��oZ�Y� ����
L�򡙔q����VfEX�/�n�����Q�S6��l���]��E$�r"�tZ�	]+N���XˆO)Rwh�h�
�Ǻ�l��n�*�
Ԯ�%�tac�-���5PTӅǁ�0���5�~�(���7,�%��vj�v��@�7\���qJ��2e���X�K���b��.�HEC���]�L�u�{I���HE@:V�n�u��4ֳ���Puw��S��/B�!��	YcTUW�:N#.3w$eP�&��[�7�JL��
��i8�W��뺿���󫲳n�el5�!5棑f�q��*�l��`j�ivj�4K�S�zf�R֠�������Q^
�	bl�����*i�i��5Yqn��݈Q�������6D��J0����d�Xs2��a!�5r����.�ƈ���͠���ժ,-�Mj6�z����Z$�f
��Q�a������E�Λ�khZ̸�)�U�Sj�y�`�h����T4J���{x���VD��Eъ����M! r�<�E��." ��z�!E�{�ڲ���9����"2�㻵DtS�c����ʅ�+i;��uux�Yѥƶ\_n����e희,"��i�Tw�鉬l0]������\!��4\2����ۤ�ϴԹ�L�Z0�˗N��1O�u��J����.�ԴD�JV��,�n���&�dm��c��h��l�O^���z��!*�n�6��J�R�P;�v^��%�Җb#E��݋���6�KPs�%���-�l�[F����)JК#\�R��x�u�a����1|�!mE��Z��2GB�u������@^��ei�k��X�9��i��c`1�⭌[a:SLvܧ�#��5�e_�]#��ݵL=�R�����6�Ew���`�?:G`�!�1�Yw(f�ѳVEfJEX���ʶ5MsK֣�Y�i/]��L:�{��f���S1����G�3([���B��OI5D᫙��eKq��@�-���Ig-Y��l�>'2�í�p*�ǿH�C�P���iD5��Ќ�9;�_mm�CB;�E���ެ�kUۗM5Vwu�E�T/ށz.�iF�!�N��w� -K��]���J����,�(�ޅ��Nj[P�w�u�eS�y�RZW�&کj�(F�p�V��;�:�:��ga�lV��C���9� �x8�k��u��B�H�y���;�! )	��X��*��I�To7]Ac&��-S�m�@GW��&&��A�-�)������:i�����{�5��*��j〵����6����Zda5���&�3�fd���ST�L��״%������ eb�5���K��<�E�2}��˦�u�(��luZ�-��؅h�����4�nQ	h�T�Yu��"�-�k����Ȏ����.l�{�ӹ@�%�u{�4�]f��qD�
�0�H3�-�Y�i(avoCW��)�
��]��[�Uf�MZ�����Q��V1b]^���M��Kf�v�M���5}�1eD,�2��t�Ŧ4�&� #w�����3J*�6�,�YF9V�e>RІ_V��i�n�],1cY�*�,�2�5��
2�(mhU/F[Fh�����u7.|�hP	f핊��*s	ҙ���
6Rsڛ[�����Rihd�W�V"a��B�2�6��D�����R��A�Y*�����Qm��� ��p�Q[6���23n�ݔK�B���3wx�A®YAv��Z�T����J�D�PY��V/��y�QF� ����j���Meiv:�'�n����	{/�Q�v�ڀ��^Ed9C`5��������a��{f5���K�Fwݐ��c ٌh�%��qCwYQ�M-�v�r!�z�]�5c�������9M����5Y�]P��`�#j�CP��)+�hKB�Y��9�U��1��{��5ժ�H_S���ѱ���E��������D��n*�OW.N�GJ�wME�!�MP�6-��	X�(��]2Q{���U����>�q�CVL�I=6t�cX�wz\�ndJ�� ��n�Gw���66���S�/c���Dh�� {��k4�	ɻNB7��A!S3�Ҧ�K��͚7@��D��9�h;�ʼ�{��ea��
��Br�S%�D��t����*LG�GP����	�Rm��[x�$Z&A��]�:�kM%Y��*�K[6�k7VJj�=�%Ռ�[��V9E|���!���{�z���r�h*�s%4�F�FB��e۷�z2ԧ�#A��)*n�F��ٗ���:�H�Ey�q�&���%�YxSr�&1"�5�J�;Q��a�9��Ӎ�x�(h[6���Wʓ�R���5t� ΍D�r���>x�srk�Wd�H� Vd�GĻ��x���=�vK���ަ�
��+YQ���4��;!�)�5C�\�!r�[�x��J4�Q�[���:a8�[In�Qd����Q
�Xԭϝ�]�' R1N0u3X�B����"�~��UX��J��E;����U)�@SЕ�zDF�ۏ-匡�N��TJ>���@�4F�<�^-D�,�<2��؄�]M-^U�j� ���r��@�Z�w.���ܥ�����:�����S;�H8r�si�d�L ��٩`�V�F �����#Ym���8);Ք�����i��u�W"E`�v:�rfU\��K4+S%O�J������q;�Aش��$�9��iɣ�%��>E��`��F�����Ac7iVIY���
�d���5Sj1�Kkr��H�t�����tn���I56q];��U� �h)�]�m�+f�Zr*3rJ��N�E�)�uP����M�]l�8��7.P���.��JJqQǁ��`"���5`�,F�Zx���,�2,u�%�:C3��T����S5`��[WxB�L5�|1��]f�7u��Û��t���7�.��x��V�^}���@����;n�� ���6v]e���V&�hLc,۴���.�B�����!8Lt��U�[��L�\�����]�I�)4�}�&bרۣF0�� �\n��]㲵P(�x�:Г�S/X��R�v�i#d�������͎��De��Ū�&"�1��[-�v]�eW%{q�A��g."ko/,Ђ����b��帖i�����B�Р#�]��^���4٠�*�r�e�P����7Sۢ���܊���j!/h0q8��cR�ՠ�^y�Mij=�n%w�j�
���9�U�U�U\XR ֍�����)O9y�H���o��b�q�����916�D++aVŻ�w V�p�J���{BiU��k����WR���kI��Mh�0+�<k��⎋ $6��)60[�gYYba���/N5�^I�,k�6�!=�����Z�ݵD��*��ѠWY�(����m�{�������â
�N�;ٯҘ��0�ba���ۼx6\ô���K47*����08�ML�rmQ%������]^֊[�LVE��n�V1��` Zbc&�A���k�P}2�ۖ��ѥ1�y��O�����\˭�/q�I%Hjv�Z�9���I��!ٙ�`��N^�:��4��At	�I��k��+u:Yx��
nV#w�<ۼ6�M*�. #�8Ч�D+ө3E��r�ⷊ�Dt�AP	kF]l�Cc�e]�M��;��dְ��v�+�
�v�ᖪ�hF���Y����i}*�7Wxͼ�ct@"6�]���]CQ�-=��$C*Ѽ�ժ��,��Ku6�]�JY���Y1�Ym�#. 45��Y{B�ԖxA�M*C/%8�G*^��ᙵ���y�ѵg^"H`pQ������(ܗQ9{n�+j��V\�ۙCSov[H��u��6���R�"WJ��b�\I�����T��w�R�V_�[� �����t�T$}p�*�=����3/^y�V3��X�7E[:��-���6k���{�*���(�,6�`A�I)F�R��>˃x3@[��e�Z�s�hV�����	��-�|bcveH�M#����/"(2��"����\F��Q���Y�kufd���%�p�91B�ۊ�e6��I ǚf�j�ޔ��ަD�}��O3E���E˹1�[ڐbî��
fL�X �K0
.��l�XyX!��r����b�B���1c/Ył��6�;GE#"4a[B����U��-O���Ym5�3q:���V��GR�졨���4v��5�sX�[��X���)(L�ghe&���Z�WY��H���uepY.�{\i���b�l����uϱ�Yy�#6�Հ�=�GM'{����A��[�p
�yj��-$���
��Q5���V�k��S�U�~�CvJ�:u�C���m�a��d�$�o[�oG!6�Kk3�<n���V�>]H��bu�1�!x���V���-�����[BK}/on`]�mA;-**��Q���s:�v���ݴB�B'�һ9��f�K���Ikɉ�u-D�v����T��na���r4P�:�a�F[�	��	NP�q�!c;T��0{�f�7�\3&�7:k,�uX�ɶMJ->{�g*Ov*�r��cg]��Gm�ST���Ȣ'3u',�WO0h�}��&��T�1�+&�AY��;���7��9�S�i�Ve9\t#.����ͣ�X�Wmn zE�UI�v�9����]M��#���IP%4��Fd7��R�O�bT�����]c�.��f�n�pr�-3�:�
�o��8���s-f�Q+0]�� ��D���zm�;k�)�ɗ�)�E)���o[��֘���Tq�k��g$P���f��R�H� �a���3lm��]�|y�u��3�D����8�P��[�'�$��u���9n[؄n �];���S��Ѭ�^#.�S#Ԛ��KU�� �:�nW<�e%�8�LY{]q� bq�ήA������g"�X9�`��/�C|�j����Ί,���;��*ڽ�����N����k�{]B���P�2�_٠�A3��0t��8M��e5c�:��C�++Z��@���S�iM�u�[�n�T����x�S��f��7Z�7kPN�xt���rrZ��1��ˉ8�%)u2�#��AG�.9ʙ�W�����֯�<�qΎNM���kx_n��VM��1�T�XK^r�+����F."��x�n�k��)53Y���3��}\n[����[��c�9u�sُg�s��u�u?�����M:�E#G2��WGoz;꜖ܲ$[�ٶ0P/w����������Er�W�]\�i�ʲA%L܇Wbmr��p��><�=F樫��ŷ��+tv<���ǳ�)�����s;h��.����I��8�-��
є��7��r����:�	�/p��iTt��&[�{�w����f�2i˗ N��
��V��v�!J_P�r�N�CK���4�u����Bw�i7��7\�4:-��������V�wV��^����*������g�eY	�R�WO�k�V��P�fA������CwO�F+�͏B��;��]���?5�u|	������IM���"H���9e��N�L��
�L�c�Y���oz3=vP�F���t{J�,���l*;Y���*ܭ�/F�+�n��r����
9\�	�W����c���[';�¨���5�.':�C��cq��U���f��D�ˑrG�T���y��1�)�h�aѽFÏ�I�t��\.ȭ�w#����.�9���9c��J��w%oG��[���is�nd.���!n�K�˷.s�i�����\�D�V�줇Z�:)ti5��Uܽ E�N�_*����Ǵ+Ւ��gx\橼&>u�m�8�xJ]	�57��ׂ\� �.�bT;)P��T�Ew���7&�H��ԫ�T��sK##l�ڷI�:��M��5SQ��eq,f諒�ݰ�B5�WJ�BpƝ�
�u^֞sr����Ζ�;�h�a��J{l�"��l�S��.�ʯWU�颳J�As?#�3����ۄ�i�ۜMB6YWq���K��2�E�gLh��ASS��_ ���h�b=��d4�*֥���f�4*�Lؾ����b��8(mY��X-�û�!�^�H�V3]=N��^��or��o��Y�fZ/HP��j�|��ys�m%�h�E�B:�wJ��7�˛5�eY�(D;�r�w˾�G���[=�2`)�w]]�Ir�N�ti���|��.&��3,	aV�_u;�df�E�t�ˡ�>�/�{�T����#����Z:�;����3p��9P��t�oA5�:3��.�lBr��N{b�5O��o9���ۅ��Fb4��V+�jSˡ���� �d� �r��˿�+�֪Ѧ�}4W�r��e��������W�y���
fpӱ#.�\e���L�{�̺`GC/�7:r�G]|s����� 8�|49־폳��|b�)}���:���bz��-��33vi��7Vh<I$`�E������[��I����\y��>n��1/,�w�3��`4m�#�+9f��m2�t"gL�P�N�Y���xRd��Є{�OP٧��,
|r<�:��z�\�J̬�z�s���d	nLz�%�"�[����;e����>�VjN�L�owl�Lt`� j�����Ǘ�g}�FTF�w,Y\�lӨ:-��S��(�y�f�{�ځ&�v��V���R&�\��hdk6^�[��F�����2���T���U�u�>�\���&�)���ܼi�P-B���lᴖ��ZS��q������w�4C��4oH�}J}u����Zv֝��/��*�%[5��xWC/�w���]79�dd�u�%�;�t=ǫ����2��8e<!�$�;����S�p��f�����yh�̚
b&xv,�uR����1�Lc�^n��,�j���v�gwJ�v毺�c�:��Q�_E۽W�/�jp\��\�¥����WE��]̚�3ݖ�a�[�,����.�#�W����`�9�Lx���L�����Wi0�f��&e����߽��WM�u��pȏm��5�S�/(:�)�W]�;��F����zBXY��'u��m�v�V���o�1r�����7�8�ٍ�]�7�g2w�w�w�vs���[�&TWfa�qω��g�k�Ēg��Y��5�qm�TYk�ef���[�r�`���~�R(�h�:��L��*�b3���u���ЃH�%���X�2��!�)0H�ݥ>�r�ݮ�����r��h�;\�j�:�c��� �s�ۧ�����ͫ�h�ɐ�	�{CPL�Ѱ;ò�L�.���M[��<�'j��қ�VU����gT�z� /��Y�ȥ��z�6��d�c��r5�6��뺜���lb�Nu����t���}��W[�)�7�h���*ܺ�J�誥B�^Pt�Ng0ödfe!Z�r��L�W)w��ڳ����������6�L��kB�;0VJ���o%�)�Q�YDh�׉����s#�I���sy�f�PrB���Z.������3��s6Q��ռ��6�k(9������`b�vK����Q�,���N]�-0Rg�C9���a���Iދ �v�F�:���`^*w���-��Por �}�^�Ig��^�^�|i�Ế��Y�ÿ��]gV,}A.��6��7�8�U�KG����(�/�0��æQJ�
��XwXtdi���H��\�A�0�[��ys���J����RYq̆�Ě�Yx�y�kq��u��6vT���&
I�CI��Թ�Â�,T���z;em9x%fP�N�4:ArQݼ�e�K`Q�Һj՗�t���¡�zwq�95䯸��n��J�d�\E��C�I�iT0_�6uC���4����Z�5���q}K.VH���X��D�YÍ����jb6��
�h�e˖6�^��q`;Ԋ�8�n6�
\(��}(;��u����)�K52Z�7<��V��[�̣��vE)R(��7���w����[ۘ�D�gTl��vp��q;ؠ�VЊ��=�Tӵ�7:�v�&p��Vb�a��e�JM��l$�)dD�gU��F���V�����nX~g���n�>�(�i##��^�c�!F�_4֏k(�4��T�9���.���̚�|HgK|��μ]W]�m�:�m��]��R�aң`���905w���UW3!}R U�]�eԦ؝�%]�d��ț��c�t����m��T��$>�7�o�\��V�A�T�b�iSS�<�Ѹ�'B.x�Ⲹ��+�Ͱs���4�Sϫ(礄�O~7%�K(帝��VJ�O |�:(����DE�j{"�L;�J
�؀��g�Co򾖴�!BVF��Z 3�Y4^� X��-&��,W{ӱ[�>�+�'`�x�˥;�:�s4 �vGArj�w��%sS�;^��[ʀV؀����k�ѫq���o*�ô%mXW�OÜ�&cв�P_C|����A�5� ȹ�X�t�;/*�]	�(��()V��iu�dxV�j� ��tA.0��6�riP�
��9x:�x�e|�Q��!���[}�`�V��rm:u����� �\�7΢��<�l�o7�o3%ۯ(����t�T,�Az9V5X-���[O���U����s�|�29|���R�G)e��e;ʻ��j�eNv	\�np���Fu��ٮ,YE�g#)�Va's��\�N�O
�va⦖B�%R]a���e��������IĚ�n�er y0^J�WP�k	gc҄�v�#�eMx3�Y{�V�.����ǽ�T-�I������B�N����D�G��FP�*����;�m��	c/�Z�2���f�K�J�s�G���=|d�]Z��2�|���iv�^��k;p@��9|8��]ג���3��Mzk��g5Tn�3L��Rj����&���Wm��v�nW_R�Y#����u�y���YsvӺ�I��a���W�>��'h����fr�4y�`�(֎���֒�={wr�Ê�T�<L앟
�g'�.��ByhV�M��#�]�f�71z9d�-�l"=b�uWN�5�G_e��+4�v-V'OL��M���*��w��b���^����r�c��f��A)S9�"9��oT���jY�Ԣ{�f�y�aQ-lr/��<�%B�*�ͮXtպ�z�j�t��3[��k.ăCkjX�]�!��"D��@rfjl]�e��p�w��;ۊH�]a��E�{;�T�5�*s��7f��kq]�Z��q�q�K�5�/��>������V��=��;���!\�ʌ�=lSx
I�gnuw}��Yu��Ĉq�xK{��m�s-�A�Նe/�v^0���|��u�5زĭV~ׂ�Ib�kۚ�Zd���&�+�j��5���s2�>���L���.��N��8�P9ʣn�����	>�H���Jn�ͦ�[!�Bѩ�n�e���ه���fm;�t�#�[������y��3�\�v���)�Iڞ�w$fo.�Y&H	��iN��B��ࡷ*hӽ�f..�$��أFୠ��8η`*�6��vk���$d4�k�'\��wWQ�����7��MPS�޻O_u
!�Z�P��T]%��lz@C^fw_v�Vb�ʏ�޽�a�}�X���1���eXZ��n�.�82��ز�w�Gƺ�8�9t��b���fiIaY�K��j4�gv�2��::n��D����h
��:���}����,��S�殮_t��Xq�3&�nu�$',��|ѪڬP�Ť�I�e��0��野�w��6P��㭦ޭ�(*�9>j���(�k��om�RT�
�J㼴�Ӎ��8��`en�>��RJ��b�)Z���G�r���B#��H흞JN@]7�Y�~sRܪ�n#�'@:��۝����������W���]"l��v���f�T��{;c\�=o%O��f�㾱K���}�2���J���p�����՘��ܬ��+�����gUEKM�41w�I��k��L��W�d$��}E r,���1�����X��N�X��*ѳXΚ}2�C'5}8T���ODU���KOHz`��������n���4��Q�o��.�{��Y�����7[Ʌ�خOvHӇ��;O��zj�� 9|*K�W	��Ӗ`l쾺��ۣ�%�ϻս���Ԉ����Ee�[���{9���]�ӊR[J��}�m�ĂzƁ����+�Q�6�Y־Ɣ�w��������W�v���|���ܩ�ý��.$ۙ���-��C�:���vj:��.�W�h��1��x�}�B��S��o���ԯS�uf,�#�E�as�!A�_P	^�-�Ih{��K�w�"��D^�σybZdX�1��:��8�٪��5��jh��	�ewV��'9���s&��'�]���Ô7*��S� �7ڛ��Zt��P�C��õ�\E�qٴBX�et�Ǹ�D1ӣ�_�j��W>�J�TYǳ:�+
yW�B �����>��`�s�X-�&�FWUp�B.e�;s'+�i�� � �h�P��i}����QVL8����wi9De�BVv2����t���Y��U+
{����s]�pm^�T��ѕ�'��'��"�Q̷X�<�f0�-G�P��]�Jn��[�`�^�ˊT#z��ݻ�Mn�b�zd���B��I�6j����+b`P�s���f����B_>S,�,kX8�t/E��3�d'q�m�H��F\�:�Cj'�ɢ��l�׺��t,SY�X�!*u��Pd�gKc(r8�\����ۏ\y�t��I�x漼Ԏl��cC���9��+�Y�����n�wP�۽���P�a��I�1��,�9$�e��i*q��0�a��"R��&55���j	��Q-M��kY��2Vk9yσA�tFU>:xF�c�i7��@��YO�yը�k��o**���C��m
/��t�W��vBE���)P�5[��Z�9�ckK""�`��<"����[/h��&:����+��F'W
�����.'����+x {Z��F�F��ju���5Ӻދ�w��RT]�[�D�a��nᥲ§bV�6��'k� x{������ﾈ�>��A�Kf���T=�ܻ�S��aJq�}E\��@�nf�9�ƉΓ�.u)��.bVxV��V���}[0��4��I�uo7kթ��إ��']�_w��_*m�f�X���î,\"��,�:�9P���M��r��5��6[��%eowsغVve��i���	����;����[�v�u��QQf��#�6������BF�������v<�F��*��t�s���k{{Pk��t����@k- ���Kr35)�e�[s�9Vs��u��1S�r��:W^��ޮ�-8��hV�����
4��L�Г׷�9wGmKk)p�l��e�I���S��& i�ln��!�̥m�9F��L��k��gׁ����Z���T5��Q���O��Su:�37{�Ø�l�S���w:�U�y���*��噓k/3���@�Z=��Q��\yk �wK�:Kog[׻n��*�$��R$�`��R�^h��o*ձ�]��qn^Yv�q�W�i���2!Ib,A{%�ͺ��\Qb��J)C�EƮ��8���+�Q�0D7�Y�J���v01ѺH�,��9-L�-��[L�b$s,�Oe���Q=(覎_�0���4��n��aS�O����dc��%NKd�Mld�'�NT.����jZ��WVk�4kAZ3��ѬЏn�S��	�ٸS꺂�m��'ԨGgV�B��L%ҹMJ�ڃv���a��,���lr��c-�XP��'���hgZ"qZpZ��5j�g-�>c�*���Ҳb˾�k�q��.V�UŎ�j�9p����#��'A���;8�S޺��p�=:-��v��]M��X�c��[s���q�Y��z���0{�7��P�5��;��n�V+���c�V���2����O^s��Q�{o;�Y����CY�W�H�V����"�ejȜ��[�v=��@��,��u�0nf �K]6Şvt�8��U��-}��>u�����jA�R�-�:���'����.��������ʭ�[ݝ-�;e�Xsh8*̫�|7iuMzoB(
����쥸��yHR�ו�VΥq���-E��+�nΓ�C:N�6G9NVuٹ�]o�W�آ��y�`�S�X�p�:�I������µ:vl7Bf�V� �o,a]&�qAQ����ʠ��\�i��9�ZSrV�|v�dLU���:/]�o�f�{�����u�V�k�������h���j`YY}�q�N]g_B8��=��6���3�R�n�/��})��F�v��OڜT����5�.���ɝ��<���a���=÷e6�b���RB�i�*�dUjep�Oؕ�2Pu&���yhѮN��y�eH����ܖ�e���p��+k*X�ǰ6;f���)�e���Y�vZyS(d����P�]� �^ꭕ6�p=������I9�S����3.�2hV5՚6k4��IX���Y���Ջ�,XS%+��G�R���B���Wn���e%-3 ']QPv�HnN��d�{�%�a�wu(e��$�V�gv���\�b�m[����6c}��W0��<����)�֎�E�v-�(�"�Mn�I=�2�LЄ�&�3��f�B����;�,e��ԑ�V��-mum�Ve���﷢��Z�jF).�&�8nɂS2��F9���C����˫$�:����9,�ui��*^�1uu"ԯ�K8;�3}J\��}�}�A]�|I�������j=�h���e�cv�O���mp��u7I[+�\O혾���݉��J`�7J۲���M��I!#|w�`�wZ�������S^H��i4(9���kY�����!�F�0>�̻V�[=,�+���[�wbɻt´b�|�Ӳ��E��yh�Ha4˻앉2i�b�n��I;�gV�6,뱆*l�˺�#,�Nb�>3��U�I](T�����EX�/�2d�eK��@�t�{����U���̵v7�SQ�]�K�̈́B��ީ41��:TQ�
}9�}ҵ�tV�9.j�7����j�W����z��P\8�'�aC��{��r���Ǆ��+km�Y3���䰦3|��nqY����(�6�����P}����Ql����VdK��ܳF.�v�eM�\7�W;})fN���8��H���s6�HS�X�n̤t�]��k;��Ӱ�W�)h������v��|�vM��:�I��=b�����]W�9엍��B�v����ڛ�u��7�F��@��{ +F�O(����u�1�[˜�xmjE��׶0��TV�Q����(np}u�2��/i�;P9��\�O$M�:��/m�Ʊ�G2��T��9R^�Sek#�/�c��y�g��㹳$��f��oKv�.�ҵf���5��k��g��V�jf�/�$�8�����κ����9�R��μ�is�Ҧ��;k���]٭NL�wL��0���j��+6(�삖��'E��F0��:B�X8)-v�-vV=oh�P�%û*\�/����t��4��3ֵ�v�]��X��o�� :�{y/��k&N���W�u�+d�S{^����ǺޛP�L�2ȫ�<�%vX!���u�q`y�W:�cQ���M��`�a��C9W#��t$���+�y|[p����9��;�Ӗ2��D+�c4���j3���oK�kM�]V/�A&�5�J���(�����?���G������W>M�S�����%��3�b��Y/(�,����i�붱�Ы�G5�J�#-i��U�8)v��,z�[<lG�:�� ���n�۳��7C��ig��v�o"s���5�
�\m��98�s�nJ��L}�5:�*�P�&�Ώ4�P*�f�W�lɭn��oOC]���u�b�[S�HW�r1k'K��ĂW|��E�B�� �Uք�Z����q�ͮW�8�����stCbi\��Eൃ-�li�Һ |4eݽ3��5�)z�P65���j�ٰ4*.Ժ�-RMfܬ9ږ���xS��њ�t&�B��n+Ø�sI�E��ѡxv���h©/����&`��n��໷��*4�լؠ�-�Ow����Nl��%�ݦQ7N��b<De��Q�N�,��M�Ey|m���/�GdC\�J��*�-�چm�z6T�̥�n�㩃��tu��H\�TZ�����I�C7����Ǻ��%��3�����[�m��or�RfX��n'P
�ʻ+w�u���9m��dꓮ�oX��˳���=;_tc/���6W��L�ӧ��ܜ����� [Wu��]en�v;�W:�u�S	*�m����)���W���-�Y�F�.(�W���:#3 �:KE4=/�XY*@��q��c*�H+D$�D%�����ԉ�����
��f���G���Ҷ	����p��
�)�hc�x#��%�	�6�����fwN��& wOS=cR�ap-����hU���y4�<����E��Bn2�-s��+nY�Ń"��7�Ή���Z�$�r��.�cX�q�Nd�%j4�>��׆,zu�=7nJ��k��)��r�/��]���v��vi��f (�F�a�v�G���e	�\����_)����PqS�����
K.@EwU���7��P�͋na|� /
7������qq��$(�F����rg���ϴb�x��c�$N���l�e�+k`��41/-�������V�"�nk�ǧ^ꋷ�
g�y�t�/��=�2vpb��>��'l�!)�Y��k�F��Җf
�*6��Z�U���9�w8:�ծVd���"@Ķ�܉ؚ�)+$���|Er�Ǌ6S�W;+���#��ܤ�wv8��a��pS�&rOXΧ���	"ڀ�V�F��Tm<�D�p��FR��I��Wj����:4s���3�F�G��b��n�9�j�9���|�@6��`�1����b�K��X����r͉��0WP�Ч!@WA��ϙ��z�O{C��U��[�,�4qφ�e}$1`T֔��yۈ������\0�K�;P���\BǦrɥ���
�5pG���Qv��XW=tC�[���_Kf)�������O ����RG���z��f$�w2mf��]m����=��a��N�U�`�P�s��ч_v��穹�&8e�2���#����	�GB7rV ��Au�lc�Z��pqBI�Jኻs��o��l��F���a����ʺeS����+nɭ?Iͺ���Ae*�}��{S��í�S���֮��;�vԖ7.,A!}�u��n�l�rS�sg26��^暚����n�;���0��-��:�x�5t�:�&���^���������+B,���YH�E�![{N�Ӻ���2��m+C�)��*�%vQ�xo��Y}�9̻T4`o1�(�Ð���=4n�j+�D��M�\)K�nˬ�]!2�N�D*���y�o��7�_*�K)ɔ,l�-*X�(r���\����0�,˖�o<�is ��wp��kgo1���r:׻ʎj_���[��+��}ݗ����5�v�eA�Sxuw1�أ �!�	��,�n��!&��K�#�%�n�5e]�t�4��[]���mF�Vۇ�$��=8�N���(Ĕ�wh�]��
�J=�Á	,t�l�^vLA{�ֿ�X����ZUz���T�\�D��]�{\��n#��ҭ���9�d�{k��];"��oU�,�o�B�i0$1ݍI�
��L���u��K6���,�.��o� 䳓�"]�?(9k)e�� ��v���J�I��au� ��'&�/��+����kD#{�Ψ��3�<��w�,�L;%\��T��{��3\�MKGh̥K�Р�n��ynN�;a�KZ��ʌ2���S��A.�vXS)���g2���̰e�%n7.v�a4QS�
�r�]ڂy�Cww�4(��C�#��xGit���z��	��<@�����2���%��&�V�5 ��c&��l����w��ѩ��c�墠f�Y��^6��'Vۓ�
��N�}I_l(o��,�(V�֍,��QJ�VU�̼b��C�wU��|�,�Ϸ�j]�ew֬U�.[��+e���^���Z��պ��eq�}�q��6NJH<�]ʛ�/;��i�D�K�`�f_>�&����l��j����um�d�`��Z]�ѳx{���r�^���鹸���'t�.�|#���,�R�V���GyRО��Ŗ���dtZ�m��7����T9K*���}�F<��Ub'��$�ޭV{O�Z��m��O�f�7��Jbá�X������AǾ�ᝍen3����+7�R)b�swN�].rz�nEr�v�gHp���]���x����`n꺄\�'ҍN�L��9V��Y7�[���c8f�W#�`����T�c��d�|5�-V�;�t���e���G<�f�(�v��\��y�_n2>�*����k;$�M��P{�Zi�����v���ï,V�H)��9�:��hLMӣ(xd���[{��6��D��E-�r ���`Y�ʠ� �׋�yE�l����1ڱI;Nts�n�:���C��<9W<�t��;�
y�E�Q�8zgr�P�|���ݡe���.Dw5�Ķ8�zvµ��ɴ�B�t�����F�ت���C'�$M܍Rٵ-�1^
��}f��p?"����mR��=��37AJQ��{�$�mḔ��\�;/y�o��"�؝ۈ�88ʘ�	�د	�c3h��{�+�ޢ��r>��&�i�s(��4v�閦2��Ic�3s��d�2�d�Vր��i�oz�BN<�!�U:ڕ,��j�R�n�;;l����+1*V+�lw�I��"����vb`kÊv�rﶒC��tV�n�ɉ)�ȍ�I	��z�i��H`r�F������ß;q`"�M��Z]=�GT�P�%b�{�����˵A�>�x��fO��9m�"�]���4��Wc!�m����ӂ�pN�	.�`��K�{�,����=�۵tO'e�TiJ�:��u7��%���
�8����|�#��k��l�����ϝ$��f�yN�vD.;ͣ(,��|.��R�a���p�w���Հ4� .�^�����; de���֛��Q��{k�v��e��"����}����O=�Z����^q�S�j�Sm�=�sT3���"���./�B��p՘���Y5{�9�I?Gbidɒ�1��s��L�=��Vk�T�;�6H���;M��ZBef��
��,&(If���>�0I���\M��X�k^_��m�I�G���/����z�Zv��֕��f>�]�@.���u�6DΝ�R�����o�Qҳ$���Ux���T�8�4h�D��y������\�f-�0(xp��U��#U��f�wWa��f��C��m�!�c#��}I�w>u�������ưPw�-��%�K��齗��s��雍�ݧr�;pIu�p0f���>r���w�u[c�.���}�|%Z�6m;d�2�s2�]j%pW-���s��o�:��v�����V\Ѯw�y�ZH2�ol�w�G�3�S��q��BT��sX�z�՝�{S�5{�/ I��w�u�1a$�Y�6�D���Jx�3����ɗً�U�|����/��x�Ӛ��־ ��N�F^89
vc�f�1��2@��*]M�΋iXF�[��蒡�t�ۺ.�f�d��vh���F�����+z;%�7)�Mť��ƒ�iT&��O���W=�u�;h=w@�v�ڕ��'��<ʫ�Ǘt�I���"��ta��X��^���v9���ݟ.a-�t�M�ڸU�U�f.̭�!؅�H �3���j�^�(r]gn��J ����Ҟ���P>�x{���}*��c��pr~��9U�x
ڸ{���L���;��W/�����$9x;��0l]wZ+f��T5>�ⷴ�u������@��A�S{\��A
�)^N|a�ȕ�i�����`��1��Un�Y(��;��f�V<u�ˤ���׫�˜�4�tl
9t4at%:ގ�wՔ����w;�����Gtf	�+;�J��s�������`$U�\HVN��n��f����K�(81��[����q�D*�C�	��j �"u�]@㡼wg<����[��$S�Q�8�\��tn��%����D>�u�@�^Fּ˻��yQ�qed~Ȋޗ\r��.��v�9:ަ@9��-�X��&��J2���U&�8�����.��uL�+6�lK�ݛI�ܧ��I%^4:劽-���d��n��1��*�U݇ž�s$aTq厶n-7�ٶ:�-69d	�4�b�Z4:_U(�9�Ļ4���C����J��U�Lr*���,�T�_e�&v�g�K��:�ءوи�S+��
��ʬ.�5��V�!�w:K�p����|�O�s��(oeno���v����)������&�M��٥���1XP�O���+�Uݼ�u�]WrĎJdk-��fs�m5��`y�d�.���l㌜��#R�Y�T�<��`�%���>Uϛ��4�T�N�s5�6�퉩��Q/.+;Y	�i-�E�A�����l�-,�si�2�R�Dh�Qm�ikEZ��-��eJѵ�laJ��kE�ںԪ�DTbZVU�UQ�YYS:��2�iU��4D�*E��V�-(���*�rb҈#j���[A��Xdh���h�0���Q*��G2��]�*6�ջVkUk+����.j�C���%V�+hm�%Ex�e���-Q�*�im*ʕ��Z(��+F�V۶L�m[KZ����LX��)Z�X5�jT��ͤ���-h�b#R�b���Th�E-��Up��ۙQ��+F�����V�j��+MK��S&�j-ce��"�J��QYD��&I�,�,��b��j�G*��T�Z"6�[��e��*���Q+e�A�W2�(�[E��Fխ���[K�D��h��&A�UG�`��+�b2�Z����U,�K�[�w���������2�[�X�}�Wot�qS��꺚9�5�v II`��[�V�ͻз���2���Mqn��Z*�u�H����А���ֶ����C��� U��=흻!����� ?W��"㜑 C�g�6�H�u�t-.�BS+�@��������KB2��:�ݤh�֨�:ۿ�,$�jY+Ab0e8l��g�_�v�aK���Eq�[��皵�e�p��ϱ9��TgN�����DD+5�-G%�_��/C�u�L,�.���$ASN��ٳ�^\�8Fs�ƞ�X��߹��$G�����>� �m���F���A.�� C�ܤ��p��>N�u��}��1(ή�r
9��Я;9� ��U#�sn����y�x}>��]��9d��c����X�������U�,*�OW�0����7�@Wٝh<:%�o���W����Eo��w����R�N���a����`�癎�p�������F�
�����3Һ}iq�	ث�V�s�K�ꊙ�OEb��+���岑ط1�
��`��$	�_N���5��Z��Y�U��Al3]�����Y�ڋ��5r&Ԩ��LV#ed���<x,�ev���d���|�z�{�pz���,���C�ʦ��z��&�����a����}�0�>����wu*|�j����u#]�ǧ����S]3��x+��t
��V�ZWC�8�U!_����}-q�)�a�g�ޭ��VJ�\�8���J���G�U�&+�{b��&��\9ܲ�9�K�N�Hi��F�����ݼ�2:q��t��
��{5+17;7�����ߙS��	
:��
�n毭����E<�5LI���9K�`�E�N�� 8Z��\@!��1	���V�Ä�wP���J�o�uP����0Н,��߰o�99������+ऩ�6&\(Aq�Tx˝Ù�/���v�ޤ�
><Nf(������,���y�Q��2NO*K���ܥ
sȎ�?D������u�1��y�[��\ey�y��r,wO�&��Q%����7T�h�I�����Q����[�˄H��M0���eqʬ�. 9
b�MP&*1���@��C�YJ�����;��a��N� �}�~��ąDaa�p��(_oK_�g9I��0��(�xt4m����vGnim�u��n���`���$�=� j����e+ߩ�ٽ�@
�h�S0���E;Y�bek�x�W�kXoz��/;�#w9
]7�ޥOT�ν�ѓ�T��r'��֟�8�n�9�O����((�Ẳ�v����vNVCS�I�k���Ww���̐WR���6��9'A�����\�U�.�3w&���O6�]����Mq׼7o�4j��nWq;��;��<���޶�3��(:�@X�rp�%��8\]�PK'���8ֹ���`to>x�L�a�o�֢Z1�����'�튳�F�{�Lf�������[�:�-���\�a��m9k�>wx��q����邱�eq��[�_ϱ�?1[�>������
0�)�������eT�9���W�QAX��ɂ��,.5=�p�ܳ��A�
��,:�[����A����z��q���5�t���A,���M4X���p{L&V
��!�5�7	�0/K���t��ًnC���xO�-�&�/v\y���vz�r%�ͧuE��Ȋ�{z�����F�G�#�������8�^_*�AuG:5O�_"A���mK������,ȯͬ�S�ø@�����=�n�W ��ɀ�ع�K��Y�^4�c��5��k����p5�Q.z��f�V��/5g��|��:L��mR�uu��4�(H\�4���iVG�1|a��s=Na�89̹1������N��8���wЉ~Y�D��^�w��<��F�ή|�Z*�_r��e�IZ�J���|;Z)gf��0��d�K �֙���U�=R���k�"\*������V�Ps*S�\�Ʈ{�Q�d\=ۆq��/����ݚ�2q[Kv�R�Q�6��=ܯ>��I��1"�c3D���������2�zP��	��Ê�U��N��ץ��.L��7C��+t���ɡ��s�����S5�@>����m)��f�a��>EH4z��@,Ў�uD�ܰf�q���{K�R6��y����v�fЮc+7�S�%�Q)���b0�W�ʸ\�/�>F�'�Ǯ+x��P�L�+.�5���Z�S�X��(�ܵc�:L�p��m����6�01��+|.�����s�E�m��Z��Դ���9Hޛ��@r�b%�������p�jȱB�����RP��vz�5���WQ�s�ϣi�<,��c@�����dj� 
x�����ۆ��vs۔c�a�bl�*/�["����Q3�@�(W�3��گ�l�B2��k��se�N�u}�.�}��]�pn��mB[��g���Ajh��S����κQ��ί���D*j�����͌��8�U<�e��Vi��$�[�z�`�5�ڮVȬ��Z�3�k��P�TY�U�(=M'���zo:��.#�,�^�δ�N����3��_N��:t�+awܱ�Q��v�w�fb�ki����|�Z���F�ۥ�r���&w�P9�����O�f�4ȧQ�3v�g�FH�Pc�GCr�4��X�Ж�WM9�'�N�o_Q�:K3�{��:Hĥ% �7�\���s	Rg5��.9��<팎����@i{>�w@"� ��J�v0]dˊuW���hV|t0�蔝w|�Rg>#��-����?")��ī�R�c�չ/��kHB੆-l���|[��x\7��K�t꺟.&������f���mF���e���uĉv;��h�q�.�p��LS�����L�j�M}s����X�� 8s�4ED�p���bbb�V��fp�BL֋�o��WC��s[
�js�`E���Ts�dU�DP��e}��F�爺��|�q�k=��X����ڞ]qO9Y����e��;	&~�咴#���Wו�fe䉪�]��1NƨN^j]�i�wJ<��c��F+���On���p�i�6H��tmp��:�~��m9���j��@��ΊQ�(��`ou��:�CR�w���3mw��)�^F3�����s�u�S��O^\!.'j4X�(p�8k��)Q��$\7���u�m���9awt�D��&�ve��Ը��>�����t$�v���M��Zc]��-��a��u���"�,T�qr�|;�b����t�ͥI4�M��1ر��0	����s,�������db������cR�V���Q�� v����9΋0����!۾��c��a#a�%���S�!��p;W���ӤM��q��
��;=K����zy�D�ܷ,}>�y-�C���~��|��t���65W��V�|��b;Bf@�����8�Qp��s�#t�o���֝��
���\�:�+�D�T���N��q�j�^C��e���jc�E\d�<N�!��ؼ�D����5���z��$����Rʩ�������8��n��M���@n�韺��n��R�tۤ��\���v��S7%�L0��<���U��葰�7�g�q��0�c�`�6�P��J���Z�HN}�ۥ�})�dQ]OB��{`��aA�uԑ��HF��N�biU)��nNA�dk�4c�� 6f��W���9�l��'�%>�M���T9�k0$�<Ժw��q�[��{� "�I�RT웙A�.:�Tx˝Ù��&Ì�VLhy7"&:��.��L��uC\�.N}+(�o�l�v�ㆥ�HY8�s}�����ﮬ4جթ��]\�u:[w�Iev1�\~��)�o;������3��ts�F�V"ź�OG*pf����n�nƬ�r�$O;-�u���HĪ�7��2�$̫|'tt�/��ɕ�y:t�J�m�wGBa���}]qu��EL���kZ��j�����+��ܸ��:��¨���H��9�Ì��(csƤwv�}��/��X����*\���Q\uR���;D�X����0uE�&�FDv���VK�S	�����¹ ��vI��]#Rp�ꏽ�wz��`L3K��5�k�r��N� _V�~�J�7X\�l oYZ��3�&��g�:�We���p�I{NJX�����X�)����@
�����0%�N�#̹,���h�h9�hl���vmT%�T�{X��bˬs�$XҾ�F�iU��Cw���I���kU�ms� y�.?��;���kM!N��pZ@�K��:<�vx`�Z4Ǻ����ޮࣞw,Jg�v��*��\�oi��2)���.?E�Utn�_ga�����E�uS�n߸��W�D��_շ\}�QAX�h�i�h��[v��1>�g�5l"Q�HỺ���B�GqSUL	����.��2�N�b�K.1ľ1p���P�su h슗��d�6��0�m)����Q?!)O�a�V��G	�����N�$ݚ�b�R�!�o�9���c���*��zS��^��{�/���dM�]AS��OkWd�+:����t��zA���4�*�Z��Z�1�x��8텰X��F��c���-�F�j��aw!ʅ,�t�J��nô��������;���[��^�h�riN�4Ro.����V��'�F*\�$x�\^��P10�]�R0�ilq��q�>���p./�pU��m�D�p	l��AY�'Ǘ�ձJ�f��x�'�����H=5{)ITK3�2�Ó��^<�*��G��F�c�J��{��j����.�X$��a�T�1q�3�;���9�=��f���T�uĲh��asm�U�f4�)su�U�&&)�D��,n�3���
Iղ��P�`0�v,��Z�cL�%'.��X��^��n��(��s�~߭�ɨݔ!�K69X�-)�@UsS>�����l��s�]�爛�7� )	<`6�͎f�3v�\Fm><#D˨L��0�v:������Y��6��4��s	��42f�ǽ0�\�Ɇ.�6\�l�W<��'o�^�纆Tˍ�Qێ��9�(��,4�:�l�n�����-�|-W��]5?.��U�+��~�s"������>�^gخ�f��:�o�kU�_�8���a(�b��藷�W��!m�j���JW��㽇������E�Z�:Za&2T��ȸ�fZ��	ٕ��mm?�ƛV73��q'-����W�m��r��*)��&eٌe��ܮ�]}��Y�����Ѫ�0�]r�5����1�M�K�J�E��ZU����;э�M1 _�]4bE��m�pty�VTN���L%`U͛��q�^���eR5 i#���Eœ���~v6C�2���W����^�⦫�o2���i�g�����ˎ��_�L�ߨc���8q���eK����k�}�V��kw�g'��x��t��t��(r��!Z�'���B)T1g�T&���-���8���3���u�'M�����{(EG���wZ���+�6�͔�CՌw;��ڼγt/;B�@}(6b����*v��p��3�4[,C�K�����R��1vV�]�%�b����KkE��D����C���ƇH�P������t��嘎�V���ʰ쬂�qʒFpV��"B�d����d�1��Pw��e���4"�4x�b�;1��Op<��G����y�B���PT'�䤀�.x*O��3xfM.�S��v��z��9V�r�Ȟ>�����uB��T7�ȯ�:" �:�c���S���|�*�ݡ")K�4y��ݼ�Q��6�ǵa+�s��V4�����6�o���X(u_��P�|T�W{�G+��f���ӣ.�ÐW�xm��~�[F���6��e.ꆁq�m�c٠�`d�����>��s6`�5����f����(��XY	�N���܀�Q��(9|��:^oQ��LMFj��a� Fb�f�|Ԁ��C�w��D�,��e��_
u^Wʳ����9���;�M�W\e�J��oK��Ϲ��cTt��P��8x@GbJ�]�{�P%��[5-�Cxv�pP�E�;�eB~޷��G:���B����5����㯛��M	�6��z��q&8aɎ;`��@C�����mm1��u�]��7g����]	��2��n
�}�wMė�,o� �]O<�� N�~g�\NjP����b����Kѫ�E^Oz#�p��+/��׏�":n|�8�S:<��O����;���(���'�Q-���r����|r4�.%�zk�r���^�ٲ��w>�@L^��(��62�_dT<�q�֔b��ޘ�o�Շ����'-��ߕh��Ծ�G�ʴ��b��N�&t:r��IŖӛ q�R^O!ḋ�m����:{�2�ҫw���3cm��/�ٛ���V6���H	L�9�M}g�[�j�"��}_=q=�q���渧:7���e"�hR��{q27(�����*^�]�0]m� �m����I��E��p���X۴.�
��<z��_�`�0�>]��N��*�{���.��J��oE��Q6���]����e�wX�۟K�����Apv�q�Z���0Zה�$���ȥ�+:��V�WJ�_*��[�\񬑚3'P�ی�s�R�@똶��X��bO4VѮ��w��V��M�|�
��Z���U�2aFt�+_u
/sO%+@�jEى:�����
$�;0���2�N���)<��ި�f��u��{g��2��H��e.�b[���1e]�t��-����һCV�����O�8B*J �\���gk�[x0O�jb�.U�K�������S�=#�Ri+�}�ZB��x��1)�#/~z�"����M�h�:6��K�'&T��V&������¯,�Sw*�@C~^5MX'�t��	u3 7�x��r�e�V9��it5�D��^����Ӯ�S$J5b�Ũ^��>���>�O92)��+�T/o���P�8u2T���,m���;nJ��N�Z'KE�]Y�Z���w2��S)e�la�_(,����̦aVS��;$�����{����q�0��S3`�{��9��i��jG��N�L��v�������>��3�R�f�̖;z��9h�|'�����鰊�g\¨"3�:�]\-�Ym&+;�a֮�$�F�=�N���&���썓 4��� �'s�v�t&��p���z�lٔ�D*����T��Jswb����:�����K������V{X�i�)ܱՔF�_q�*Qݫ���R�
}�u۠�)֥	\�y9lξ���I:���z+s�'LSb�m�5;���ڙ3|��ʪY�`n*XV.���0�Z�`^��g��FΊ*R��u�-�N�f\�\*���cV���)ܺ���c�#;��A5a9�u��ۊ�SYS��q�L��ֺ\�i��F��<�u
��i�y)#��#���s�)pF�^f�����k�ì�k$i��+J]*��;�P�b'	��c��0�l�kS����ޭ��B���{�Qq��Xq	�n+��,b2�N�U��X�L�yW[��]��
�.�9*B�4���K,NeE|�I�6e^̝��Wop9M�b��w:�}��N�R�ξ静�qd����i(8�(|�4�-��vk����]Gʂ��~��C�xot����;=&4�Ցc�@�_ ��s�i�g��pjҖ֧��������oG�)19r���,�!BwҬ�i]�V�_ms��GW���Ʉ��=�]�MǶ��ޣm�P�qh�uR�}G��'t�r�t@�P<+/�B��aV�䌾g%�wy;��-Pd�&hmS&��Ӛ�N�'�7hR�9�p�V��4�:�00�r����8)��v��WZ�zV�A�2Q�uɇ5m�]h�ھ6���]Y>Kn����yB�w�7v����� ��������6�����jV�m��v4����m)kJ]k�v�J�PX��ȕ�mX�"���TJ�,��Q,����cR�Z%�eKn��R�E�֖[F����[Į��o+q�eE�uɆ���Ռ�sf��hڈ�J��[U-S9�+��� �TEDDTaZ	iV5(�j����Km+)D����T�٫[c�Qep�Z�B�F�DQE`�eF*�5KiZfU�e֢֕�b�AT��kZT��YA��m�Md��[J�Q�۝�Ub�Z��F1���Ae+kbV�Ԋ�����l`���
"��䱙�̢*�Knh�QWm���&j*""ڥT��6�mF*֕���([�kUEFs�"-�R+9l`��ɄH�V�X�S�j�h*ԕR�¸n�Dm�����Km�b�iYm���-��+-A0� ��#�� Պc�l�S{8�GրV�Y����YrvVlz3AqsHP��[��+�oA*p]HL���x�Qj�>�q4H˸���;~m���>0�7����AT��'���9�g���x�:�L�I�ѩ�=C���d>����C�=C������������%"����>��1��"1:O��]�j�q����u��"8DH� Gރ����+>�^�}s�L�%g��C�=$x���Y�'���U���<L�uC�z`Vt���釬��'�C3�<fC�~g�ͺH*��W�9_���U�	��֜ɹ�Ҡn���F�P��t���fK���I�
��'~{�$��ed��=��:I��:�s�Ϝ�v�C3��8��W�J�Sh�d�!}��S�X�!��}��>�}*.���ђ��.\�ЄB��'��h�$��zyޞ�$a״��I�����ξ�=L�Og�ߺO��%eg��������!�=eVT��L�ƼH/��&�_��1� |�)t=~�8}\�ѫx����|fd�;}�)���+���8�a���g{I�=I_�y��H,���)�i3�8�_=����={fg�δ�~0*����L�2fS�7��DD�b#�D�w���н�mV$��*����9N�� �!�|�l�Y�%@�>j����&EP�|Iu�~�a�x�}d�n��\��z���a_^�;��'���Ru���0�@���0��9�Vթ���M.����t��̕�
�}ҡS�;g��|9I���!�>�����<N���>��2A|~hq���d:�=N$��L��ʓ�+
���ϨA��A��C�(���"��n��\�o��R���-�y���� �}�6� ��J��^����+:VοY��?$��9C�z÷$���8�Y�O�l=�IY��S�>�Rt}��z�C��?~� x����]w��������e�@\�r��ߨ!P��H������Vv��I����Ă��ɺ���d�S�6���+���&d��d�S$�
�d�3�t!�J�O�l:�c} |���������2�w�7��IR7�-��o����@�HC���P����x��z�&d�>�|ghd���}��� �����ϼ���^�����eg䕓���N!�W�}dړ�2]j}�$�
�R�O?u���ٿyt��.wf��.�}B[�K�ļ�Z����l����=���
e�9.��X��Câ*�{ŪWA�����T%pǼw�g9;����#����w��MtyR�V%�6'u�]��^<޹��#g�qo��;�7�p�y�߾���������t�(�^$����'Ĩfeg��g�q ���������@���!�d�'�χ�9�;C�d>����|H,�?w����ի��Agoi�}z�#�E��sӷ'��|DDp���zr���P�i'�>Xd�<�x�}�I?3�;����	�t_�񓴓����;g�}��!��:�c�$����v�YP�:��S^���DH��B?E2NШ)�N�3��}�ΐ<J�Yîi��&}a����@�x��aןw�>$�����p��Rd����ֳ�%gS�(q;d��?s�wv� ï{� -.j*�����P�"��x�ן�>�HT8��K�I�)Ă�ψ)�x�'�P�I��2��O����3�2�&gl��'���R�^u�P��Ă��î���G��B���kY~��� >��z���C���?0�<�d*�^����I=B��|��:�b�Z����*Vv�R��2�ya�H(p��<Lö�:�C��i�z���yIӥ6�>�)s�N�=���} ���=C���]��'��������� ��ě��� �ğP���~s�O�8�eO���t���:-3
¾yd��s�į���g*B����������疹)�Fi��K�T��}�}f~y�@����x}���� ��|���$������ ~J��*|����2?���> d��|�N���<I����v���:����\�r��h�mg�!� ����u�� ru�8�'�g�J������ݲ)<B�~���S��������iĂ��>�^�=x�!��&@QI����|H.@���}�p+$��ug���!�P���D�'��fx����>/�:H,?'G�9�&C$o�J�$����C��RW��?[$�
��:�b�HT�!^���u�������$镇���ژO��\թ /N�q�*Ϣ���T�x�K��)* ��{��*tö��RqP�3���t�Y������� �G�Y�?'�:�a�T�q�y���I��w�*�}}�U�hi�ۆ�.��˖u�ޛ+��0]�8�t�NJ�ל ���v[����}���1�t��I����B
u/��]���(|9T]�g���g6%���h���<���z����nI��kcV�u9�F��:�Wm��DR���whMUz��"'�y��L+
�ݓ��]}��|IP=J��t�E����sY;fVj'�_�O��^?�z��}��?'I�?X~x���3's�2�~J�$9�^��þ�h��	��Mh[�� ��1OO�c����a��q�g�ę��O��� �?$��ߝ��y~�d�T���Ȳv�|a�)Ğ!S�O�u��!^���C�����x#q�x�S7'�sh����E	}�b�~��/t��g�����D9��|}gĂ��������fx�&�y�q��!�����H*�G���:L��2úol2P����=J�!����-D�[�'�����H'�*���ukI��|�g�������i�'-���>�8�*T;~B���I�P>{���x�������}C��=�杧I�!�?s�|DD��">��ئ��C۬�3�3�}��rJʇ�����o)*;{s��:O��q:~�d�!_��a�}@�����
°��,>~���>$��O�n�Y*,����u퓱�>؋sP��D?|7���{F�3=�{��j��S��D��׳b>�D�
{��I^$����Xed��'�Yă���4;za�<JΏ�q���ę���Ht�U�!��a�0��iTx}�x���H��|��v���sf�����_!S�,>2��|�v�O̞�Ұ��A�y&N��
��3Y7t�'g,���I���r��U���C��:H/�|�3P�<C3�|�$x�P�����w��5�nll�h��b��p�E�#� c��"8D`��t3�����zu�:@�*�W��_xv��'�T>�ϼ�+I��8��y{@�^!�%ea���|ꁙ�%J���:T��U'��ϧ�{�W��T޾��w��`�#�c�=�l}P�&N���~N�<Oe���'�d���Rzʇ�����C5�Ag~���R|@�*O������2OS�i�Y*� W���0�+��9ϗ��Jf�[s�r�w����!��#�#�CS�����ʓ���O��z�+��$�^�_,����q�yO^�v��H>��Ȥ��'������Y>�a�~o� �2|��:C׌2�8��	&��]�_Ws\�������r+��a����
!"q�R�܅��`M~�rJ]]�����Wt���Qj;w+
�Y]E�yd����$W����7�B��Ƴ��X�oGNù��i<��%K�ܳ:���\�Xw ��L�/��G����o��E�@�˽�����{I���r�$giê���2SS=����Rg鬞'd������'I=B��>y��z�U����{̽�z��S��'�7��w�3��1���KΫ�	��|庍��2\�o߆�T���>��	�Y�A|E"�=O����b�H,�'��x�C$���=C���ɟ�V}N���T=aߞ��L��+�z��#��G� D��~�%W��h�����|��N!�����OOߴ��䕕�o�� �2T�78�+;d���a�x��a�>r�5�P�ɺ�4=eN$p����?'Hf'��=eC�~O�{$��}����x??u�{�akZ��$G�DG#�G/W����'�ox�aU퓯/x�J�^�o�z���2J�����QeC��'�^읥r��!S�|�ԝjB����Cפ����>w�����ð���35���������H������!���Vzy�H/�~���d�� |<��2VVz��?g�~�>!� �>_>�Rd2N{�>�d�P���@�*,���[�%I�;G�I���!׫{��,����߾�,�@�S�����'��p<I^�7)��;�fx�}��<�}~��AVO��1�%}fH=O��׈�'hf}����� ��{�&C���2�XT��D��ޑ�~�ܬ�Z����p�bY~�d�P����w����J�O���*�~���u�#�y�U��ur�PA���r�5��pϑ�պ�C�< ����y���:�;ȉ�������[�nܙ�������e�G�B�Y��k!�[�(W/���i _L��~9a�0uJT�I����6��X�aӻ���SY\4f�5��<J�3��r��q?i��2�x�f��!��z-�>22W;�t�v�i�c�C�}��p'��-�3W8��Ē'Vn�I��4K1[aӱ�,��3F�Q�^�":��j��s2�z�����˶�h�J�0�k �V�z�	p]������Nз�}�f��>��59��󫬁h����❾:�0���b1��r��ו<{#d	����R v�X���.D�e�sD���l��of7��À³М�R;nc�|��v�<vZi $��w d>\�g_X/�jy)7��Y3!�����t�p`�
WT��VHU8	8�\ɫ��t����T���\���L!��ej��Ru�CMW���ՙ��ư8�=x�W [ܵ��GN3\� l�T������ohN����L�Z2����<���j�S�IYp�R\7�#Dld7L�,�������]4* �� ��7k�S�̈́@��~Nwu��>LTe��4]�؝�+�yD
(#�IC�g�
���:�}�R����Nq���p��rf�����.q&�u�7ތ��ʆ�Ү�`��9��ND�}�N�|�"�d���n��Tc�ud�NxԄw&�pW$��gb:^�������VOa�#X1��U���卓ALv��Y,Xr�jA5<*�y�ۭ�~��eq��fr��9ʂ�n��{)�2��cE��x�^g��醴	��ؙ�o�%a��
Z���:;�\�q2�Ö{�4��f�ì�~B�Rp��<�^M[�T+78j�&i�4ಚͫ Qᩂ�v��DG�JӲ����j��� ��m��i�K�q]������g��� �����*�'������9;Ѯ�&�p�#��F�T��a���ᒒ�8qWC��?�����&_�R_?�4��m�`�{ր���H�{�wq�3���D�K��p��[aqŢ�P.�r�i/C$�po=UI�S�`�Q��p�c��yh��(h�I�lp6,ߦ�:�h�lj[������w�g\��*�����I�=���ct����E�B���ʔ�L�I}��ˮ�l�o��QV��W�W���u�oKok����g0���S����N�L��u�u��u��Q�����eT�M��T��FZ,?�K'�
F'(6����Qt�jF)�-z����ꁃ�d�9�*�־�w=&Y����l��X#�ۖ��O;��_�Z�c>��C�]�a�ˆ��@!) �g���	�r�h>y^�1P��/�6�h���/��~�R��7 G#o��D'��n��@�݊*<8������&�+7l'��X�d�Y��=�윮���qJͭ�y<Tʵd&8̩�@��ݕ1vY3E��Ӡ��5a�)ã[J��-f�
�.�ݬ�2uci��[��K�sR0�>xI�}�����V��,�־wRk�rS�js�z�jI�Ѯ�u�����/�B��4�,��M���l���� y]�����t�7Z��irj��;Nv&�a
q11�����=�/�,5���U9�Ns7�#�.�g�3#7`�v�l��#�u��nO3�7^���K�$V)cw�R�H���f}�U�`����ҍx5)���0Q�6:b�������g�:�V��yb.�
�g[�q��Fp���[�Q����v.0ot���� � 6��1D����&��|��Ê��jܮ�4�өXK+�y˷�s%�7��B����Gjp���p��C��I�.�j�Z�[1w�Ĺ�����9���qx>��و��w>nk�d��hF�Ϩwe6�2�/%^W��vͩ{���X�]�+�Qp�7�)��Pq�����#����*�ݤ�^c�$���!��dVRcy�p׸�v_��lU��;<'�ѯ|��z�X��L@�1��3�����L�Dt�NZ�Fz��s9%y�
6����G��J����t�U���v`�++:�f�8�����l67�v���v��ʼ�s�{Lõ{y�EoMKvtھh뭾V�G��֝��F��O�v|_�l���K*9�݋nU���}�$�)iz�o�:b�
�����&��q��o�r�;z�ۗ�.v\�ڬ�܋۞����}����S�3���Y����u�y�{����Ҵf�SG�r��Ե�,��ȧٛ��[����әr���K�k.
/������x癎�,`�Y���DU�܀Z�<��
�;�����]|Gm9����h��8ʸ(P<k�뇐��i��=�"��yC;&�Y�p�oj�2_T�o���װ~��Т�r�F1;�%<&�;H�C����`��]P�4�gI�ѧ:R7WRp�\���+��A<�a�*a�[,%�cW�s��x�KGU��jEYyv���ʣG(�ԥ��h�.�d�Q�������e�ғ�{J�~L�uٱ+�m&�,B�p�.��U��!�
�
��$as�S�X�a�ū�D�;��Ȗ��6E�c�k�p����U��[�#�LX��EE�D@�����d�F�LMy�8ړ�n�����k2���ćI>Ç=��#�ț��v�%2ʜ%��b��L9��e�R���!����5+I�Q�(;��3�s�j(鿓۸x��qlR��mRԤ�⨹�*L�$�H["z�McI�s--��x���|p��Lp"j�_�>�X��ճR$;j�CqP�4ݪ�O��ܚ�r�Vu#vū�=љ��;�f5c�Uw��|��[Ω��*���9�Q�x�n��y��u�O}��G�r&��E�x���7�*N�gW8(EF)`�mBb;��1��j�T��yOjT��1{���H��[Ύn�ţU�a��B{MɎ_NT!a�B 0��������S@k�����)P}3�z',P�s����C+�ñ>�0�G�����U-W9��G�׉��C/�]�zz�ϋex���Z"_<����:l��ʦty�I�Jfq�F�P=
6���!����g���I���ZX������^T�썑&$�8v��M+<�`ӷ3�S�y��76��&t�a3[N�,�'%���!_�K�
+�&�Go1�+�����2����&���Bəb9����h���i����r�)��֭ްR�J|��
�m.eѴl���&�i.��+sy`l豭5���MںD�g,[׼Xȝ���k�Yo!�<�}_6d�!��TD.�gI
:�킚Glf�nڨ/�lFmu&q>��{$`��L�n��Xf4D$r�hQ[O	W�K�f�^f\K�����o"u*�����'pRJ��̋���k-~�R�<m>Y?&��Vs�����v�t�.�s�vR��ۯxާ)؞o)�!M^�,b�F�⮑�?�!cz g>5�э\���V*�����%fj7;5�B;�H�mum.Qq2�����D}��j�N]�|һ=߸��W&�D�D�&CS��'z ��yDPRT��P��C�����x�)ni1?s���xỲS;�}ɚ���8��\��@��."��Tȝ�Q���qNk�*�.��t�(}&���9�F^��h�ʏ��g&1���R�0NL�7���I��w��I��a;���yI��ڋ
�'�!����A�r�%��9
c��aGR���i�ަ�ڶ��6��hz�:��ٔ�i�K�q]��j���gf� �'�)H�	�R6'3���
;����d��1�b�^�t�-�� j���P6��^��7Y�c=w������0��,�fӮ�Y_30���@Xu�4�'��+\-w��zT%=I��L���|�or�f��=V��> �`mWx�/��ek��w���(V+��1;&�D���u7a C��U�a�'zFK�D0�u�g���-�ӄW1��.?Eb9��kٺ���m���O�
��K�y@r}M�
*���%}�V�pY�QAF��ۦ�����v޵�sTu���"�%�u����h��˻����³��B�-�͒��Ҁ4I�k{2�ۤt���dP2�l�Ћ�܁�걥�����O37���rb�6��T
:G΃[O���e��q�y��W�,F�d��B���2����p�ܪf,W[˱4`��)�M�FV�lHs�p+c�m5��32oZis�=���3���3�.��O��]�N����S��x���܈���;%�v�4�Eq��L6�mҾJ��Hk;��٩g6-	Ⱥ�h�h��w.�mm��d�.�N��kx�3n�K����{X��p�����b�;�NIŮ7��-v;��I�BW����ml��/����:�C9�n�ؕ��]Hr�d��]��5#��_9jr��*�����HIgktŴ�i�)1-�����Y��x[� <8��hݷ�%t"��s:��B�L��M�g,�����r���Ç��mK<4��;f�)��@��F;�C��Ѭ�xS��Wj��x-B�4����,tڗ� �Zذ���r�jX��5h�η�&r�ԇ��;r�)�w`�3�gWP�R+�ӷ�y��x��{3m��f�%ʭ�u�II�1mc��uu��]�K�D�A���m�5J���5�j�te7�]J<�ʱz��n��`T��W����Y(I\iܮ0L���D�w��gE=b��d�e	���[h A@K���S7Ʊn�oR�g�t��أ��y�n�o����2+�R0�����4���^�즮��Q�|ͅպKx�[b��}�]��<0��pA���ܭ�#�H|vK�7YVnU�Q
񂦦������m]mbC\�>1��xz�gE]{uj,{9<�#X!Лr��55�W�p�:�򒼛L5\���Rط��������fPF�[��f�ԶF\��ZYޥ7+�<9x��S�����]�X{���e�$xve��
Vk}�;��s��]j�E�f��Վ��6�Kk�=C��C*4W\Y788*Ù:So�����Bkw�e]nF ���4���Ι]Lsaآ�	wţ�*[�Px��{n�f4�e\�9���Bj5�r�J��-��8�����ښ:���y��K2����m.T9�3~���M����NnS���$߻�X�N���B���:E*>ڼ*����76�
v��4��8��{�D��PuwtO�)��G��#�h��p�j�,�L�YY��h��v�}u�^�*�e�p�#���)�Bv�\$Ju8,Õw3��q�3�;9+#.Q��Y��O2��\L�����w{��.�d�EZ�2�Aњ�|k�s3_r��1��G/]Lw�T��S�	sXȥ����;�P3tj����ﯯ8�y��Z �$3�5 �S�}{��^���8yŢUЅ7�5X�뮺U�0�;���{��NS:-�F�b�=xv����v�W>�\�����������k訨�V�[�:=̑�;L�ݚzop����(�*��mb-��ͬl�e�E�L��֍�V��fJ��75mkEbR�2�63ĭ�b�QA��ʈ�A��-�6�a������J��J��YQ�6��(�Q��V�"&�4*�[m�����D�����
�Ѷ���_���n��1(�`��`�5��[�ֶ<��-��V
,E����E�mx�UU����.K�Ȍ�meѬ���V�DbEE���*�F��A�$�jZ�����\�na��������(����G�m7R����m�x�A��ujG�j*-J�����
��Eh�˨����^n:[bԣEykҪ�*"V�2T��"���U�WXѠW%\��*+%�����8� r"���<j�"�鸽&��
ֹ�FKv���ŊE&���T�Z�cmJ���E����mBڪ**�f�
�E�Ԫ��w,���yj��Z�bV��P�AU��DE�R��b��A^m��R(����4NY7�D[��w终M�����k!�Jf��&��n���o��o�u��%t�����_l�wEG�-�Ы�q��`=��]>̫?�ۘ��R��0�}�SB��H:�xCe�H|�o�z̤6}#�v�l���(zy�%�qm$c!�2�Uw�:c6!HU5� oT��"[�NB����5(A��I�N�j���q���1�Cs�Y)��bzd"���:0Y��\��8d�fLY���|�E�״���T5�)��I�r&l�V=27��G\@ ob��O*7Y��:��w��R�s�Bf���8ۨ�gJd3#�Brp��yd%m��t�]9�P7�z�*�9�N��<$���"Bu�Vb����c�1k�5��sT�s3��fp����+��w*�%�u�rQ=%i���u��O������֕�*��X�0��*toU{ڞWgqe*���:���z�/iȣ��o0���}u�@����n�jܘb-I:1c�z�m��fD1MH�9v,h� �:i��.QPo���wV�Ks\�玑4n�-v�{��� �e�4m-�c!��e��	��y�N�0���Y�{�5��ѷ!�"��h+X]������Ȟ��"�
n	���S�M��%m��t_��ҩ�Lz/q"�c�A�h�.gf�R�JD!c��%��ܮX��=���s�b���\��Ѻ�t�@���Gdn�!+�pi����>��ѓ1���Y��wM��;[:;'�f#��Cߩ��E���~ŵ�CyG�#�t�ʦw�R�$��
����qpve��+qp��¶yM����%'���iT~>zV��Ɵ�@�-
��U�(��үg8��O�iv���xa|Ÿ��,���sד��5Z;!>�r��W��R7&,F��!�
K�3��[w��t�qޛ˓۹YCb�[ЬƸI�㏝B.X�6��}
���Ajh��E}Qg�vp�)!F>��#O�g"���r��9H�e:cE¥�$bɡj@��:���m^r��Ur��N:��μ@�=�����2�
��x��i�����v�GNQE69N��}�s�/$|�����W�A�B\�ьD�+���\�6ab�f0E�ii�4�:�Eݵ����Q��r*_r�kY�J��#����yμW�F��8��Y�?c3��b���o�"*���d�~�Z:A�Y"c#��Z#,e�/�"J{�|�����I�T�q�W����zY��F۷�I�wqj�w:�M��'e�O�Q����m.����!I����h����^�H�{r�E�ո�{�o��jB�4;��	Zox��8�w����R�F�}]!�M��k�>�oDfg�|�5[���U}��}K3|���n��<=Ԫ�ܲP)́�>���2�p��W��@Zj-����!km�t].����式t`X��əca��g"tr1@��Yi�(��g�7��>��1�"��h�ڽYc�K��/F�L<�L����;O+o� j�W��n$p};�\�Ym��"C�B�m�Bt���cS;ë���\)AU��7	��;�J��b�q�(��[���Zp�����G��6�=]�qXb����z�C�8E�%+���"�x��'LW�ѭ7��2���⽂�eNT!_YzP��p� C؍�@ryq�*�g/Q��E.�bU�0\�%���s��s�e�bu��e#�}�|��b��<��\		�ĭ�����=�O�,}��&�9����W�M}Q":n%��$4{�+�|�_�K���ݦ�y���*#p�ʅ��!��u���
Ǖ:{6@�)d�uO#�ʲ�o]T��zB:��w
�&Q�.�&o�Շ�g�9l�ȧ1��i��Py���Uq�^��.bu�)
��8�NS��m��r/{��ॽ5�IR���ҳ�WR�ᙲ�1��s���uh�|���Cvk/8M �O#��]�uq���MA������NgT����Ax*kC7�"�uw+��>Z��J��{��ѕRNn���T�8o�
b%� <��@Q�rw'�Q��+w�_��yn��|B^R�s;v���Z���ۅ��\nc�� h��
%Q�*@ޙrp�C����N�#�:�#�4��-��/'[s�����Y k���U{ǰtb��~�G�3�tCwT���]OGk�������VA��!��H��*�F
�]RlT.3_���WM��
����[� �t�N.]9���-��'�94�&�T&C��{�� D�D]P�yj2�ᢀ */ؗ6�Vo�ԝ¡N ���KÙ�-�ӐXk�5�>j��32y)�yd�=�*��oV����u:�c(㈛�"���!a�s�uAq��"���c�}�伧���r*�ub�ݼ��
2䓜Q;g�#Z1��U���/E�M:���*�X��L}1�}���E-��6k�N���?���A��2��9)c��+�]>�^���I`��@��,�*e�]:�N�֖���Gʨ����1w�0C�u���#�JK��X�����������[;��$C}�uc#�U�jATҶe�Y>7}���G�ܺq�D�K�Գk-�[ۺ�m��G5IsJ�)���`�FV�^��+ղ��t��V�V�y���w����wK8�Y�y���&n�ky��,���r�D���`R
���-e�G��}'(���y�;NO�;����o*��Vt�e�����b�؍�tO	�*����	ɂ�����΍�ʍq��Έ�gcT�{��7b���w�
���(;1��w"��
�zzg�U�ٓ���zNó8]��!m:�F��f�)��V�h�5�1�2㑃j�1S�2�>o��7"�w�S`��"�xpq+�+�y��n���?/>����+���I���/�n�7jFX}�<}.�h_
��N��5�@p֍u[rV��ͮ�jb+"�E�U��Z��=<0bBWL�*zx!�aLm�k�b5���J���;N��8[��o9�u��_1?E'�>	�!�
����P��tX
n�/ �s@�ϵ��=P�bNJ�C��k�+�n���G���P��{���|�N�t�T,rC���5-T�n�1��	[.`�Us&��. B���޴�jb�F��As#��'
���|/os7T"�l_Q��A�� 4��y��!<�Dϩ��ȰJ�,"e'��o�������i<J[O�i�H��,Qv�Q36j���H��z��
W&��#��{�|��
�- �
U9�GH����.�Y��@e��toM�itX$=m��E�oAL�X%*����9�"��Sf���.�/6_3����ډ�5��݊�5+(�yX���磌ꯂȯ�<ѝ�hdK�kUZ��Qu9?#�������E�i>�H_���욖�p�J퍖{w����<�WF�HnlH�9�>i��z&_�õ��-l}�}����K}�,4�f:V-�o��)q�hhJ���Ȅ+�� �!N]�0��$�%��͎eޱ�37�Q��ozN�{���}�wA��Cf�R��6�2/������r��a�=�>u
_�Z��]_e�UXT_�cE�֫ó��ia��i��P�75Ȣv��D���T�kj^�SMƵ7Tl������h�f�	
���>��g��:�oˍz�h���, ��
�W��S�{�7�v���q�͓�8v{�,G���5����+
 b�O,s�I �W�iI�����q�b������f^�o�.5>���j
�IWx��������{D�g&�55_s�LX����F��ӆ�[�3���ebS��'�uE(��z�+��/7�G=�K�H?U%w	�T��p5����c��;�Yֆ[�L�v]�~C��P*��t�"��C��uи�V�p$�����FNܘK\��%���
]�Cƞi���	9��^K߁[�e���(NBc�����]ZY�)"�t���zdg,�v��G�H�&ɸ��p��F�2ӹ0f�l2�;&��K�+����ɯ'�TG�D}'#�m;�T�裀S�B3�<�H<v9>�p-��0�i�e�uoV!����i����x� #C= k�WB��B\�ы� p\tN��#�O2F��ȭP�T$�#+hE�K��T���ٯ|��U%qXseT1�XT��&t\j�ݰ9db���9�ѨջH��;�`�,�� ΐB�L�4v;��B]C�bz.����?�;a�t��\���N`/�t@�´P�o��\�U'�F���V�%W]Gp�qۄ"�LN����d7 F�)C 	��!2D0�t��(�P�^����{Du[����tu��@�_jvl�6��|��
�%�0�P�]P�i�"�	Z�3�0:h�-��Q_�v�aI�j��W��ϳ�D2/���J�fYeWq�G�^�rV�f3fP�@l/�{M:6�z|j��E�
��f�����ːy:�P���vu_l�t�=U�i�>�!�5=y4ܘ�&���0N� C�*(�7^� [�2ɬ�x�5�5�NFVX���Xk��{��n4��F˫��8�K��3���+�;3ْXl�CxB�>�z��:x1X*
7g���Pw=6y�ޓ-9gTQ��w;Y�!;5��*��T�QH��1��C4Ǝ���A1�R����s�iҤ��ꪪ�$�&��;}��تo��vN/�u��g�:��ĭ��	
�S?P�8!����bw�1��5n��nt� /������&�9�+��T�k��7�o%�Y�h<�����=|�wS��Z��j�qf1�����co�I��k�an}-��7�+�}SǕݼk^�k#�����{���� ��f�u�7�p�2eb�Z�7�9��NS)�s6�l��b'i��}*�)��u�c+�Xq�K=��gdU2���w�����W�*�;�n�w�����[�ì3|�S���P{�3�5ۋ��P�u��(�Di{j�I1�I�y���J��me���M��|�9+�ۿ�g,t��<�����8��gA:!��Q�����:��f�͞𦝴�M��H*q�����)S���R\=�0C�2�j9������m�s��z�:�X@h�t#_1KZ7p��2=���
Oѐ�r:��x�k���7�Tk��>2�񃣪����	���Xy3?l7�_��"䩹��M�0��j9Քyl�n�t����5oq�Ex��V���g�CQ��
�&�TC'x���^O3��T^`���kb���eɝQ��=?a��j���Y��gx��J��GH�ή\�!�t���CH.M�d겳��_W������92F ��3�.n���$*�TC����0`#��r�b��g�rM'7D�gl��C궥����ܼOa�F�cM�m����tp�B��p�I��e����-�]���c�l�rT$�8��P�d��-��9>X��7vZ�a�5�'�a��t�F����:����< ���3|��l���(`ws�}�C�g@�c��/F����kD]��o��$�_�L`������ Tr��&�U@i����6a���h�"]p��{b¢�e����xR��l�R�m����X�Gs�|��k;"�Lә�(Jos�K�^�{�d����Ȱ����:�.#iPF/e��$��[�r���F"����#�׏�E�Uun�K���E^.�]�cZ:V���%p]]VL�f&�$��5�IϏ����������WF�*�:�|������)ծ���S�S}ϰnF-=H 4�b���卸U��Q�j��U�k�Pr�勒�n��yiܸt v��fE���u�aMFe��N�n��s��,$�}����{k���ュ��⮌)Ec��+\X�MX�VK$<�\Z	��q�4�5��/z�}�<����!%(��.2]��}k�N�Zp�7m`�_`��Z�;���:?G�D}���ɽ��#���C�)��a:��9�+���{u%�Jn	*��Y�;A̵I`�0��''��\�/r5\j�q��K���5D਷j�5��qO*68��<��Zj��P nb�����*AQ��1u���L�6�%N�fํ�eGF���9[���^�_�2���ȁ>�\6�&9�]q4�1c ��1q�����"���BQG��2'�ݺ:<��i�{�j�]W�r����&��;*�c�����TH��,n���dك<�j3q�K�BeQ�-�x��R�! ��� �Zb�Y�����tXЪ�(,�dӭ�mHiE�sڒ��80GN�!��������H_�r�1�NZx�|J�a��B���M�Y����|��������5PF�3u	����e�:b0L5U
��Nz�O-��o62�lUȶ�����+��3�k����U�x�ؗڕ֚����CS\�'a9���x� Zkt��<:��/>�5�U�J��,����Ui����>�C<���6UgJ�U�c7�t�&Xg�/h3�U��FyJHF�1R̉Mڞ' c�j6���4&���T�2�r�{sQT[����ȴ%�)Ws�io���$�.� �6�G,��Yt�s��gF��Z��xN8ifN눃�Ւe��r��h�Q�X�	����Zo�t��� �`��&��=�jܮڀ�`�ă،K�u��{��a0\�swDui_Vj����Ɖ0�lO���eX�Y �Q��- �y�*`ǲw�j�n���ϻguV����3�ʛw6Hγ(VF�F���)�Wk��WS�����)ͭ��;�/�0a�ʳlXw0�����<��X=-�fNcX�*�+�GW����NWb;y���º^��+mm-z��0tt7��\o1Ռ�
/��3��YC�	���ܼ��ߧ�E/�U��,dLY`��~ nf%����az�.�;e�.�7�z9=�^�e��)��쩰�(k��HXr@S����dͭ)�X����6u�� ��z��w_�	�юtx�S�Y��M<��?vTޠp���;ܨj�r%[ٷ��hT�9ش���;o�gb!N�����Zg6mƎ���$64��ްc�K��r�G",q����D����;u�ހ�ޖ�ՙћ�]��I�
t����T��v�83NT4��(�*@��#���n.K/2�͡��X8cFԽ��h�rp�p�V��6Jui�����͢6����]rA�{[ƕ�N�h+�����<W�H��r�L��Y;��W)ѥ�V�.5��>�rm\b����Ѥ�\��f��ޥ������e����#E[C������jۤ^��	
n��7���v���ޘ�z�a�E�pj����M$<�з:I���ӥf5B�c�������=�7 ��x���K8��CtaV2�s9Z��SIg.' �c	X����;O#Wm��N�\ٹ:ম�&z>v���u)�\�YDt����dP�)�+d։M�s{���~�#��8(w��vn�A �s�����N,A�;������b[d*��	�����}M��v�J+�;�rΦ���;��F�y��y�m�x��%���c��S;ef��
tgo����/B��E-CTW�a��Y|�5]vA�[��5��z{��1wn�[�N�o!���[Z^ۘ��l;�'r�^��@r�,��Bä�X���&Xo���G/��5j[�]n�"�}���؄�$�wv�K�=�]])�hf�aV��(^�K�����Jzw.��^�4�U(��{۴W�����K�^��M�i7e^�uҍ�Jz/��E���ǃR�2�k[ڛ�ޭ��;��Q�*��tJ��/U�P��`��Z$%F�|��Wӵ�n����tzw}�1��͍*��rd�iX�E]��R%�C�fKo�5�R�H�mرZ�lR�E�6�3!�V�*��UV�+X�j#'3y��D+,���Qj�R�]j�UE�--QH��+��Knk���D�(�#mF�kkT��E�o6�Q+gM��"��ȉ��-��p��Z��\�(�k��[jV����Z��DUQ��ڼK�c����Q6Nsc�Tԫ��6�U�6�h�F�k��͌��ee�P��J/-Xks�ɩDVҨ�-��-teB��ZX-h֢Ǎy�\�sJ�8���\u��֝!^'�x�Qk�(�c�5���iU��UENRʔx�"�5,�]Ī��q�*`������"��f�(�+��C%�����v��ZZ�mƉ�Q�YX�<�����U�E�n9��o)UPX/9`�䠏8n<��o7�b
ZUU2�F�K�m+-��b��U��k�χ]�;<f m1Γ�p��U���+��䬔k��}k��ұ4���� � \k"W(GD�W��ǈ�;M�����"��(��y��Ӡ��[��Wg]@��Y����5��N�	V�xW�P��:q:���U�!��kW���wJ�-Jf.�����Ϲ��1�q�j
�IWx����8t}`�S�1�����wkB���W��e�ڭqϟ:�7"�1�
���'��v�<z$��И�;]v4����OGѽ��y⻄�B�����/Nk��vT��*��2[�N���]�Y�C�t�z��ޖ�t�����0�P�RS�����:l某�6�P�j�9�<�U	yD��C&o)��0@�$䁽.�g�J3%�2��E��%��Ȳjq��2���Ԕ.��'ֶ��0�f0W�\\n�J��3^ ��r��.*΂�p�[L$�N��S��թ�W�GL6z-��.y����NY!X�Z;`Hʞ9�R���F�S���#�~|^��r��zz�x��([��`�n�J�r�O��
Q=�eR@vFfU���	HX;��;�{P�����f�;5BL�o����jb�Q�'yAA��t�+���&n���r�,"�
�K������pCذР;W�� �T<�ތR��W��������ą)��^���ub<�	:��3"Yh%�#��b��kۊb$佽64����	�Ô���z��J��ᕀ���R0o�[�q��mn�44[y�O>�٣�Vo} ��Y��i
�V�}U�W�I"3v���mp���ѯ�l�s^"갭.�#7����'f͵ 6a��ԅ�g6d��Ďz����BȾ ������<5�s��S��)f���]�j{*�R�S�T{Kz��5:i�Q7Y��͘4PG������WeEa��R��ʄ	�����׬���fWTp��ۍۑƣ�ˆ�Θ�Y�F�[V������g;�y7ܫ���F�';;��ܦ���x@_o��������ñ��GC���W}ie�Ҝ$��O�!5��ojPVG4>Oy�2�h��/�&��^�>3A�^IG��
s�8pSmԞ��E�
(*�w�Y�f��3�'o�}�a���f��(h���u��&Tub��3F�c� H�%�n�z���0��-�L�N�_N[)�p�5����j���z��.�U��h��@W�%�Q�rw'�P��C���<׬ԍs\���
kk{M�/�¬w��+�^WR�_���5�	���"<~;��Xs8�řI��v2s�ٝb-�P?:�R�La�2kq7�c�-5��J�톧Q�������r�w�����9�����=�R��8��)s��^>����}�s�(��������c���̘�����<9*�{9N�4�=D}&��٫X�{5R/���gd�f ��n�C��LW��������މ֏h6jf��k���pL0��m��q���S���R&.!쑂���7L�,3�^��7�MЩ�	�8�`%��<8-�܄k�)4�&��Bf�<���� O�)����+�$��OKk��y��}S,h���8}q*w 9������;���k�G�p��|�
,��ٞB5��-һ��>�ـ8���J�o�Ш�˂�O�3����);����F�·���E�{��za�����묀���k��zL�j�W�2������X�=��o������V�q�>��q�W%��ۡ&*9�|�ಈ"��}u�~��HWn��zY��?`{Mgf��D}9p)�4 �W����͞�n����Θ!��?�g��%%�qWF��;� �p�zs|�u����cF���� Fu�#4��iHޙ	H&��қ}@*���=bSZ�iF �z�c�V�^+;�b�xoϳ�l���n0���ϓ��\G՝U!XoR�i���<X�ל�WR��N���钺��J���kv���e^)9
�� ��/�9:��w��&la�W-�fF���b����S��`<���͛�B���y�ǖ'
T�j��L3�������ѳհ���V�PVc������q;=>�myT��8Ӭ^\���uL>�Hb��Mr�rx��{HHכu��nQ�~.F���;2�]E^!7�Z�=뫽	Vݼp	y3�oE��KG�M�Gv�>0k�/ۖ~���$C��_U &*w�#�^@1�sЖ_�IR�&M?M�:��&u�Pv���ō��Y+i U��r�*�v�M�g0Y؊������v�H^��G	��ۇ��B�ġ�������1q0��ʽ|:���I]p�q3�����q�����5r��ϣU�F�d�~�NR7���V tmM"�j��0vn��u��利� ����K��C����I����ٝ)����Ջq��#s"��6w��*�R��Z1�J�o�Q�*�*��٩���j��fo �=�t�lv�d�W=S6��>��)^5[^�teq^D������4�U!�1
�@)� �+Ïͨ�����z'�8(P���gT��"�t@L4�p72�驅ž�Y<��}���&P����c!8�Q�-c��/�|b�4�1�d��w�\$������ú����^�l���y���æ\�)QG%wkO��ёaΡd�yW;7�c��9M��� )��֎�6J+[t�[]s�Vei��JQ���E�`t��9��ɥ��/zu-S3d/W1��[�W�_}�;�7!���Ə�}���Sx�9��cD%f���"��Xl9˰ġ��5���;Gpt�z��e�}�î�fǳv����oȍ�p��0�ƮmS�d�q)o@[nN��9s���դ:n5������J
��]~�� �cc���3^�mC�������]���<�O<7��W�M��8����Ն<4Y��]Zb��E����3�X�^�4*��\�5�:�.�K�����,;���?{���Xb�ݢ`�AHV\�0�c/�9�k^YX��{X ��;^X��J� ����M���x�밻�F��t�w��.��x�<:�� ������&y��?v��Q��t����Cr�1�
���i���w���BTP%�[V�чrgç]`	�q��9
���k+s��j�,h��R�-��7�s�7�z�Rg�sC������5M�@R�b3���V��k��	�eƟ��<%*l����U��+�+��Sg�U�Ǯ��*8�͟?F���{�_7h��	h죳�l��Ģ�{m7���izN�W����@;����J���_w����6���(���ýf���F�p��(��%����
��]Jr�3�~�A�K������9�-��[E��mI#Z�rV,���f��&�Ǹ�8n��0N��������Ƽ΅���B��P�3�3�4TYB3�� $z�vM��!�^�yU�K^T��]�V�R�К�>�S��ok����F����Mą��Z:A��L�pF��%V_\:����S�ڜ��ٌ�FXw�t�Aʚ���z�;��܂,c�i+���Q&gH+6�)=�*�z&&��ѿ���&�ԙ����mH� ��Q���*�����z�2� D{�����G�,G>��|̭�X7�Z�)�@4Z�٨T;�4e:!9���ɵ��e�L�t�{p���PC�/+�W���d��gx��=���i֨��,��_NTi�ar˕FϺ*x�3��8cD ��D��*JFY[8(F"��5#���2�\K���#@'}��}ݰԺ�į5��׼�b���`�kqmu��:��qN�R/\I�뵃�K�]1h�T��D�ol�u���ݓ���N鸒��\�v.&��6l͇�����������ϩ _�t���O/��BW�+�k+��צ��ֳ mz����5�;��r�-f�zi�r��4�oz��V�=�G�˨��9�oV*;���m�˒g����:/�>��W5�6��G;���^o>��ǲI�f+�Ţ�u�x�=�+k��Q���C�G��+DbM�>�X1չ�k�tp�����ꯂ��t������/�%��â_����n��;���T�**��>G���8���2]6���=�q�с��Ef�&	C�۪@M�XJ0�Bل��:��aay��d�4[�^�u��r��>�8B�Kt|�:��1W�T,��'��̓r9᷶�r�q$�>שvCy?)�n(vo��Q�_Hr;�e2=���z�{4�t׾�~���M+�qݯE���w��_%	nښ���1�����e���'�@V���y���K��B��m>A�̯��3�={T�0~&�w�]�}ˢU��t�`=wpf\qN�4�|�S����� `7��`hUζ��&8Q}���Jܼ	�_�ǖ�cg���a1��7�Mok���󜝳�\s�r&&
ݨ5�Ql*�9����EK{J�T6��Y�\Fr\�>�Sp��	i��Gی��R藺��'�k�HjYVuNy�d��zG]+�o�{���d�'R1���슺�Kd[��嗗�q�YK��܍�Z��j	V[�#9˰��g��w$j'�2��+��}VԲ*`Z���@�{��^�|�y��}��*jv2y���n��a�2:[�+��а	��tV�|s�u:=lV����ݵ��_?�-���f2�Ou��_;��O+�to�Z~����Q~9��<������]����1��X����]P�WU	�;_uQ��'oZ̙�U�3��ST1±�Gm�U�E�u��QmF�Y���ď��`�v����[7�Q���Cih�=�qq��K:�1��Bj�xg)u�Yb�^mu�]ݹ:C^\����&��m�Vu
���!w��
���Uə�=Vj�}�z�bX�}�)�F���# ���J��k
��z���Y�m���z�a��+��|�kyx�o��ҕ����O\<��j��N��R�td���m�K/�Q�i��q�n��4�n��/�r�d��5Fk�.���a<�s?�U�yb�Ϸ�]����T�v��\j\��&$���F�7��]{����ax�� ��F��ܒ��������)8�]����i�n]��y^lɻ��Hm���Z���3	��I��w'G�w�V�Еm`���H��ϵws�:�͹G������cjK�f����u����*����D}yL�ok���/.Q�к\���
���ބ�DMG����s��l�oe�e}=[�7tҐ�X����	LS�1K ���y}�󟊿D��}6H�e�y��ns�m������Û���E&8i]�im[Y<J��Ԗt��ګ�^����a**�RwW�CWn�-�8T�=iV��Ns2W�u]X�@ˈ[�V�����.{Q	Qu�B���>F���F���p�j)ə	�se�/-��U��*���c5:Ֆ�8�hajឃm�{�]zk�=����.�jX<�~8���/'+�^�_n(��-�J���+������{��պ5F�[{5�Z��kj��ڠ���7��K������|�����n��/����ja�X9�j)�m��ih��;Q���E+[�^�>�ȭ��|��{9�yW^&�E��r)fＣ/�M&��|��/u^�o�%�;�^�F�������
��j�.V&"��Z��Ⱦ���܍
m�E"xT�RԂx�K������
U��ukM$�9�*�l�#Tό�R���w4!�7!��<l�evi׸Y��&q�l���e]��ق��p"ݎ�-�R3f�^��W�}U�j�կ9{���,��%����d�r�c��?zh��xw�:���9PA;��;��m�.g��pbw�Y�'��}oK�)�}��]hq0�5�-EOm�����,jL�U��LU�T�\�����_p{6���3S~�˥9�4�nR�%��}�!)
7�%��K�Zk/ud+�S�u���)3��<JK�I;�����r��6ʿ�BS�]29��2�����7x��*ﭶ��^��cl�]Q�
��T���)G�B��W��$+���C����w�SM-�=N��i�*��	�,�=n7+k*f-�Y��R�����ɬOv���I��|ռ�(}PR�ܸpU�1��ݍ�5|�#���h�"��_s+|�|�{5�{;l���X�Ck��ctkS�xN8���첹�ޅtW�}K���;���Y�u�{{t�Yu ����0\�k�r�֪d@�#y�yz���(�P�E�f��I��dE"ZT�s��^�S[k�9RܙW�>�h�����Ǽ�4'Qm��L����:��QV-���N��w�Y�l�H�)*ܚ�
��.T'Oi.��<�5�k	ڔ�Jt�s�<(��{�}�0J� ˢ�M.�kl�`��$�en�{���H���Ml�4V*��e@�1�8z`s��kp<Z�ُnmNV���O4ckA��X�-n����z
KA�u��!y�d�4t)I����Lr�<�'����Wk>��1}[G�����M�c�Ͷ�ˋ����p�.;�)�dS�*����1Ђ���L8먩�nik�[$<�W.��� w}:s�.���1�Nk��=�{}�%�<��M���o�Ц�� z�"V�9B��1�]��]�[�p�M�'R�] �E(��l�[L���;�\��(��S��]1�je��+&��퍣ڙ8(��>����c�w���;p���y����@y�0��K�5a<��1H{�%t:v�L6)Tw(�B�"a��}i�Fs��:](��G�M��k2�X� t����ɠ#�[M�����M河�)]�@S�2Aq+@�V+�0c���}h�3xN�ت��	\k�Z�5>:�z��K~t�ԕѮc];���z��]�r'5}MJV_ܬd��]B��5�[�Y�q�"�h� �A|��u%�V��;U "��v�x��:�Ƹ���<u5hJ�Z�(�:��sV �@�˨��7��	������7*� Iur�ò,��f��P}��1S���3#a��h�s�V㋙���\j���=�jt���E�� �Ŀ&����P�vX8brz���8wAsyM��zd��Z���j�5u�ko�.���:���u��NC�,(p|L�9w�:�W;�AӺNeE.Q�KL��	�}A���S{�Σ]�X�B�, ���|��]l�#��2W_m��uΠ2���2��5[���ʼ�ZX�h��v�(�ݡѼ�������`�}2��ť�Y]գ�lXk���Q�2�54��ͩX�3y�N���]��lѰz��)q�b֘���'X��+w�s��#�w�>y������!�"V�P>Cfպ�ܻ���*�¦����2���U�iE�I9ܵ^�d�P^G;D���!I�(G�4��sy$j:o�:mp���xq-�f�,Z�p�a����Bx(�l�ܼ��sǠ���.�؏_C��[��e�Q�W�j>���6r�,i��JE��s���{�]Z̫��3{�"ݍ|/ �6:`�`��dˡQf��' �1ϑ�N/��b�	.�}8ܼ���39�����\��t����zLF��1��e�;��9�L���0�
��o��Pm���Of㴞�4}�o��G�C����)g�Y<�R���Z���ĳ�x��
#�>��1T���eQ�UH�S��QQ�X)�)�1PU�b�"��u��[5�ڙ�(f�mX���(6֍�Ua�V��R���+��8�sP3W���رB�j+�J����F��1eUQ�(�Ė*�Ԣ0cY+�-cl֪�f��YU[������	�T�V*%֦�+*[���kl�(�-�P�R�b���"kTx�yͮ�+��KciKTTF�nJ"35�CR��Je��g���EDPMhր�mU�U�X��^$�����Tx%AB��Ҩ���-X�cmw.�L���\Z���9�]n�$--hź�Mv�]u��Ejd����Qձu�QX"��ÏYX���k3���;V���(�K�&U��li��"�R(�̥�R�TDV�J�"�T+8��b��ZQA�X�'-cdŲ1#,V�"o�����{/��e7c/�u=/��K�/��g��:�jb����d�+�I�q��0���������ib�4��菾�&U��[���ܤv.Pw�������=����K�r��
�ՙ���5���rҰK�Pc���q���>gs}�i��c����/i�}u����5-��~�,[�^��G�f���.#�m9��y��3
�a�s�h,��;���VqË�F=�]K�>�[�%�$����c�t�V�Ol�x��zy�����}:��_M}�"�oL\�w7����������J�0���vm��y��U��>Ρ��v�;ƫ����<�쇰�ʅWBE������ޱ{ڒIk�����º��y��1;�T_%�)�825��ת�N8�i���e�/T���+���~�\����8� ��T~`�;]uV�ִU��gk[��I�e>��6ۇ����#���9^�יє3H���ӵ)<��s�0Was��1K�����ތ�t�	*e����Nfsh*�Ar+k����tM���辣ر?��L�����.��F�<ψ��3N�T������7<��fXfJ*:k��qxVʁb�wU�0�!���k�aWe7�v��v�_'����T�ۏ��7y���"m����sBv+(z#��	�t}-����ݙ�1�b+�B�wve����OS��?S���s���U���Jjb^��EWuA��[�p�௓8�a3�9ga���V��������uCy��vQ���؊�8��͸C��R؛�{���Mr��	1T��n�&��)��f��ז���h����q��.��_|��k�����mA���S�`d>�-���E��}T�NH��/��7���E��z�����Ap�ƴj�k�Ɗ�e��<�����h(L}
Ļ�6���=[S�v_R�U��]��K)f�顪-����*y�����[꯷Tk��7͉}�˂`R��iT��)�^i]�N�����IioÍ��죋���:�3xPTq��Q.w���M
�����ߛŷ�u}v;�
���ֵy�����,���`���9���>��l#7�Ѱme&�;6`ۨ�mt9����|��{�-�O.��'̈�Kri��%�رa���t��&K�Ɍ{�н�'I���z�l�a�9��o�z'£F�Z����P��o�޶H�����_}W��-��sB��Nw�z����e|�kr�ڎ�\�y/C�*>�kҪǅ��9��\Ȇ�Eb[�\��q��c���қ�q���S2n�i�BݓK[�)��J�%���T_5��:i=w�o7m�ї�@A)Ȟ�d��s�%	g��`%­s�Q���G�_u�j�ˆ\�ۚX��Y��u2�r�%�Ȯ���C���q�cn���vB�Y.`n{{����]p9o��E�JQ���h�y\%k��bw�������n�am,a��7��s���2�F�aҖx٦�ը{u�w�s4�$+s�z��o��}���qyIQ�IӸC�R��.���{�L�y#�:{�;���ޅtc��bk��*.��ۇ���»|:2����T�.�jr@�S=�F����Qx�V��;�z���Z�*��=��s����o��$�Cۣ]��ȷpf嚴��Ny����c
T��W$���NB��!vT�[�o9�
��i\x���:�˛��&�V�w�y
5kE+��=u�ou��wu��j���Y��̭���x�N��������}���}_}�V2�0{ݵ��:�U����Ϗ�W������5���|�@��Y򵽽���)��;T��٦�gxdʣ��+����.�T�Ϫߞ
Ŏk17�^�Q���w�.ͧ���vX�[������:D2�:�]�1�5�)�IU�F�[�͇�c��m��t[��~�nB8�J�쿺��
���T�2���7/��N�=���q�K&�Q�m�����7���!\�r�]��#���Bn��cPz`��Tk��%x��s�CZˌi6��s����
GQ��S��j&��p4-�d�k���|�,�ܟ1�QQA�bj�f��9����Gv�յm������	H�ީs?�TZk6�������*�r�.�6�w��ƵA��S�j!�P#��K���A��orҩ��-�����Zմ�}uu�{�[ъ�噊R�_�m��������R	��F�hܧr�����vOM�Ӱo��<�M-���y
�GF#.������B�N�X��S�f�@B�A�|f�����f����h�%
�J='MۀNK_Y��*�K���_��c�{��ö�O��~���"&3*/d��ȩ��g�ˀ�2��I���+y�z���Mbiȭ3��y8��!�/R��P���4W�}�c9��'��ZL����a�}[ZC&@t�:j�9Y�r[���p
�8���kSAU��8��}ݾ�g��.\������U!��	d9�+@i��+��4���v�ዕ���ZO��o;9eߚ��3�(Ε���vз[��P������f�9$
+7;��]n+��D�p8d��MJߡ���{�U=S=�>)m?[[�膗�/೸l��	_=���u}y9X�}�;)1���|�k���Kpd$�цYW�z�r���xqpMG��?�R�jr���UۉbV$b�LX�/���Xal^����&�߇b{ft���z�1ٚ����/p� E)���}��3��7�ڜ��~BC�*(t��կݷ;�d�#M������i�}�a���
���$�Ld.��x�)���k�D$p��(٣M!W���Kh|a@�-�ylC�)������F��ݙ|~��eY�y	��;��%nW8u������<�d�ٔ*Χ}đ��Z�/{��l�L~���Q��e=�w�Vw�5��}�kSݚ�-��cYQ�D�1cv(F�YH��u������t㯹>w���wm�oiM�|l-�
f��A�)Ru��s���[��w��</=�(��'��i\k����9�uǙW��o*��Z}<��D�67�7����� �4Z�O���
ތ�Df-��������1ip!��	W]�ٗ�:�4�:�0��q=gm���}�59��^��Sh�W���%��+�g�,g4���5PrJ����l���y}���s��JI�Sq��OԘ�QvWƖ���͈k2�۷��&�G:D׫Ö�S�$����Sp�+a�;,�������I��&+'�=�OV�ֹŀ����rV]�Vۃ��R�+~z��jV��Ko��;�ݴ���s<�R��\ߝ���u�|�.�5;��mFʸ�yY���tФ��Xv���>�9̗(?�R(��G�#������,b䔨]I�J"��@~��hĭ��,��5VVV;�4l��������JChQ��\�����q�+k)b�E���)�|풆$�u�[���K�J���b�������/U�n{�i����Бh^;GϷ�o�w�4��C�O��eM�=�=�q~-Of�$��t���[C��v�8������R��R�������xI�=�I~�-�9��)�T����K~m���Ī,�U5i�w`MvOR-�ם�/"�Χ}��i<�v�\9���6��wQV6�G�s]q�ut��w�>�.0�W9\�eR��_Ͷ�)���M�\'��@�^a��ۡd�pB�k2Ou����-�]��͗�7Z���K���b��ǻڕ�FS��t�Q�R���qgi)��J\*���Q�I밚W�v��.[��Z��b�5b��r�A.�	F�E�����曙� ��؜>"��8��l��9����ܘ��QL��9mJ��}]v]���k��%�k��ى�&iN��:�Lb�B2��(�9��3}��Mv	J��,-��gnr%�>�������w<�b�v���8~����5���NT#�a�YS���%�Fҗhd}��>�`��B�f*s�W���N�L�Y7��yͬ7�F5����JWga�o-u�-��D,gREWG}��=����@ř|ym���v^���j��b�5fWR�X��{E'�e�<ud�y��I��)����A�ݣ=%fTl�q�V�s+fT[yomi�X�=����̅0چʹN�\�NʮzǳV�,�]�Pk�^b����c)��G�^��t�zJ���'Dk��B�m+�q�_��k(�����'+��s+���/�,��͒Vv�-�r��S�GC�x�s��e}���Pq]E�u|�"5�u:pLvB�֐�y���s���\>1�����)��5o~�Ҿ�L����p��^���$ֹɿWa���iOF;��6[o�"�޷�����V��jpݫo[Rpv��뾕B������9Qږ����S{,L�븡pu�[�2��ư�� ���J���j��%b���`�=F�jٲ�9\�!o]�kG3�;�s3����mj�U�J���b��{��L�s欅)E���f��oOC�B]&�u�9V��P@���w׆ԇ0ʶu���(,:ЇtL�}oTU��u�s�>�`�.��Ꝋ����t�_��WՓ�\���ÍO�9�ݜ��s�U�_[�%�%�����TN,���"��xC".��;e��UNw;p�)�mC�L�P�7]�����^8c�S�M*i�I�����.ғI}�;���dӤ��eX��J�oGL�댚�2��%'_�[��7wZ�։��rL^���)�vg�KOvt�RHJ ѕ^��E=}�Tz�R%�ˀ�3�i�j;*�֞BE�]�h�9%�S����z��02�(�٦%nN^'ݟs�L����w�MkY�r.{fߟ�f�'�OK�_gxh��T[Qx:�Ŏkynu�
헝z3Vr��/�hUrP��L���	��첻h���W�ö��<�ҳ[倽/�g3��M���}��IT����m����h�-�W�a��ez��j}c>���m�9��#�t���oV���%Ty�9_�աHejXѻp��A��ֆ�	�^�=Z���g��:r97^ɣs�Xw5[�k�x���S������f�'�׵�#�*�Y7t宩K��rw.���'��^����]G:���]*���|ȷ����Ӷ�7�ڜ��U����������g���o�b]E����Lb|�\u���Ω�4�g|m�[#��>�i[�GU�H\���T��m>ŵE�^���:��k��w/Bz+��F�?S�M�n+��Y<fq y�qʣeVh��̺�e1W9�7�Z��2����Y_cý�8-�D��k>���ΐ4���u.^�%�v��%WXĲ�mvS}_)�ɸ��# ��r5�OT"z(�w�����ͦ}Ϸ���Ա\������q�m��Lm|���j�c�t�ty��D֥�w@�N֫yђC�_GrYx���OM4����[R�O�q��,l�9�Fk�.��f�:����.wq�:~�I��Z9,��̜:��PSn�S^�'�1����yt������`-wٗ�:�4�]���<�
��kji-��o!W��M)G���Pa9��+r�'��#@�7^ښ��o6��v�[hJЕ	��jk��MX�\PwM�1���m��3�膐%���;e!��Rq�H�#��[�ȳ**�{)Z9�8,[��q.w��l��,b̊ӆ�)+_u�샆m�M<�s�z6��%����tY�ە��U�.p�5,9�Y�;6�A�����m-��|��4peU�L�yr���1� �H���L\�.�Q��r�U���{�P�-�vt�vSee�o-H:��r����)1X�� %��mڻz �?�_X�u���8ݵ;幌W'{� R�öjȚ�F�������6��ޖy���e!F��;��q撃��7��l�wZ��zo+���R�=���R��}�e����u�z�Ѓ�$��!�e�B�~ȢJ_m���9^2*mbiQ�6�'u��gL)�Y}���Dq\��{}$�J��m�ݐ���>�0wߍA�sJ�L˵��vF�8m���/��1�#+����G7�{%���ɭ#2�kjܧZG8��a�f���(��-��z;i�o*�\u�Ԧa�1�7y�&mfX<� �\[x�m�fm:T���|KG���zu���r�6�63��%�x#���8�']�����;Wb�}���;��f&�e�\F����p�yR��΀�!��L#���+��҂F}�I٨���K{��y���5!�c�s{�pWB��{@#62��:�j����Y���һv�Qwe��B�R��^�fb��s��n�lNc�Z�cR���7N��'D��1���3�Jٮ�2�w9�e,s9oP����C��1-rN澳�U�%��)�{[�ӻ�VdǳB\%Y�����sqI/�}`�`�^?�sv���֐��;q�ө�nDM*]ĸ�%k�v���T1R��vAK{��lת��ͼ��:�{�Y|��ؒ��"�v)6� ��*�ƪ�=�5��-?�1=�N���I��>��]�7�3��F�#�S�Vq�"�Qo6X���3@��� V�t�)��9M�Ө�f�:��`���	��1Z(���Vy�I���6�+���nrp�۽��Y�iD������FH:ׂ�o<�ݢ����X1E�z�m�n	YL������o.Y�mB�]4Hs'6u_�V-��]�����8SWè���Ӵ���FG���g#8&�Y���M��o�'�1h�[7`J0�C+d<۝�u���;;�9��ͷR�y7�����o8'�3��G.	:*V�!� �
�&�:����	����R[������0�P�Jne��w#%���2�qN�,<��%%�yZ�<��p�Nv�vOP���K��u��c\E���8�?����u�=�R�\](;P%%sZ����d
�Od7c2n-ѽ�J�crNn����͔��qơݛ����^<�v� T�)q׃s�:t	��+�؃ttU;��U���ـ�Ft��e�5/x����]vڛ�W'�*8���䄗à�����9�c�s��U���Z���l_ԼF�1���c�.Ki�6�"�]p��9+U����m�<f�)�Z��S:s"�VUb��l�EY�K��V��j#E�X��ƚr�ڜj�b�TU�*������e9J�n�Q8؊��R�
ʅ��V��""��b18%[j��AT�scEb*��eQ��*�ʕ�#dG�q��Z1F�yv�+km��TUV6�8�!���`�,^%�P^Z�f)���US���(�Z�*Yh�5�Z�H�e��#YU��EX�Z�EU�U�`�ͣ��ӎ��"*[yIKi��Asg�)�q��E�f�V��"���g*����Z��D�AE��(�P�R����3F(�DTfe��5e̢�b��Sj�dY5�V
"�e��r6�TmɄL�L�X�5�Dmm�(�lZ��]u��Z�GƯ9�NY}�qգ@���R��35����]N�и�}�!��0��M9T���p̷(��'Pޭ���������I����;_>j�LҕP�E&8l�F����3Ƞ�X���K{t1jj����q��%G*b�P���:
���쿠�۳��`Vh�⌓t;p�V�q��-�ŀ�r|�>dj��Q=p�]�s��Ě�q����Wo㚫��ux���_b��u7��������Y����C�.'�D&Ͼ�����j�����iw�ֺ�ާ��Ś9�7(����=�Z�����ĕ���1j��:��V(��n}�p��pTP0v��Z�[�LUެ��]P�t�4�6���lO/�.�=Z3Y��T{^�$7^Nƫ�6Um�ا���Rݦ�l�m�H7Y�2�E�h}���&�g;8��NW;�T�n���{)�9���[�hն6���b����;���=.�;�5���\��q��c��7�&��Kf�z�����OI�M��(魰jש۸���2�̔�Hy��M;��%�B)Nӣ�b˼ȥӅ��"�|i,^��k��.�kŗ�vh/i �Ϻ�f-j�������μ�6[[�Zڗ[|�MX]��ز*ٙ��6�{I��r�*��U�S�$�,.���?��=��9�����Pc�K�}��nF�M'��%4�W@����M1ݽs}����ns��ݨ�-��G)�	TK�	p���/�Q�<1�]v3�%u_kLg;�E��'p�w+��%�)���*���Jb�2��j�����L�&E��}JF�9�z�@o4,lk��WH�K��s�U��v�ȕ����7o5;���ˀ�e����v[9�sq��x&�����~�K��]��qT�3jT�5�Ql}���lqY�Q�Ne���Ȕuv�뫃=���.��V4�ύ=��귦qc��s���̅#k�@�u{���i5l9슉�<:���w�w5kF�iK��=�Z�i�bk�@���y7�GD��y���P迓/�GP��ϖ�~8���V,2��镸8��%ǟ����{���m�s��s����P���cp>���@��Q�Z����A��v��~�̪5r�m��ZWViI%�]�찓yn��-��h��y��G�Qۃ��{�\Hn�������U�l]���VvR�P=�"J�%�4�����Wy0^�@�>�`�n�5:������ɢ�����b s�c&uO���z��}����SR���\��N����9�T�*I�[�N`�ߣ\l��b�ս	�m�֩��F��UOK��T�&�x�lm7yҜJ�9�-��*1js�����e^ky��f+v����AV��hOq�6�x��3{h��@ㅽ����Ğ��T忏�:��=�ri��c���RBg������TD�5K��~���5#��ޚys=�ϳ�8M���S|�r�em�v5Ԩ1)1|��/�Ӻ�����O%]��`Ҝg&�$�Ϸm�մ�ۛ���(���:�ƞ{�in��94���U�ɼ��1K���Z�=��+f�_%O��M �`��U׵8�F�ِڻ����֪�F������<��P�����Ȇ$�w�)Rq���_�1\�y�vg|���Þ��:��QU�����Wn��Wu���r�+�B�cbV��'�|VRL릲���h�j.�ݾ�c�٫{�٘��5㲥(
��n11I8��V^�b�늆��	�l�8����Q�Ȝ��F���ga�K;��K��2ng�d꒰�7*W>z�����\�-]���}�����׋�秷Wo�n�u��d+�剤�
/��4��v�S�1����k/�B/�7��kU�ܓm<���>��˅@[LvY]��W֗[��=��Ԡ���y�=J;�}Ӯ��s���j�ByN��u��:�͑�F�G��>���
�o,�nμ7�c`��j&6��ny���/n�����#�n�H��6�uYSϺ��z���
1��R�^ߚ�ȏz�{ϥ��xL�� ���7Q�`{��vw.|�R��.ߧ�����=��U��V�fw�7�ޥj�R�������5��tZ���n-m�s����E�ur��9%��ӊM�]X��mm�ml��wَ���<*'�k1���Qm��sAuf�㜸ƭ=��:���\?WK馃�)���8�$R
a��mH��A��u(�o���f8��҃{�P�y�;۾�׃;4w��7�:�V�i��|�9'Jb�s�uv�wh'�m?3<#��Fw70��l1��������֯���k���"=�Iܡ�U��{\�3S��=��E*�UZ��\9�����[P����۔��Ԍr(��k�s����W�bv&�&�D�@�J�I����5��:~�O�M'���Q0��9�E���I�9C�BS��J������x������7 �uZ���yغ��:�V`�]L�\��mJ~��]�ٜ}Vܚ�uN��c7�r��ݮK�
ۅ?Qv��Wp��+��[�
�w�O�&��ݛ=�zC��SS��������7P�D�c�]xin��ŏ��}6Q�̾OH���/���))&%Cơ�spV�p��j&���mlu�>]..��U���xg'�C߹��mA�w.*���|2vC�U\�y�Hn�nQƪ/1W׏k^�1��+�����Bq�ңJΎ�g�덩�0�tz�Ki����~��|�~+��Mue��o<k���x��y,��J��,�̼��kj����q���~8��}4W���i���x�wB#�y(��4���V�u���/���#.V�tg̜twiM��v�I�N^Z�k�Ԥ*s�/v��Jn���{'��#U�A�(,S��L�Z���vx��Y�����w1����+�Ior��˔i�ݑM���_���^�ԯ�{���_�X�j0�b��nZz�ΚǇj#�fCr'�C��9���ېjE5���㎺����[p�a�{��-��f��t;�t��
��ݨ}�MOTr��J�\���g'�l�Q�_}͖�>��	����8`5�9��١V�= ��c�K�U,�����y^��ݹ�ӯ��r�[�`6�T�k&��6�
"�lk*
\+_]�j�OY���:]o*��Ew�u�+�WuH���=�ݔù�uHk;2�w�NN-�p��K�C H���S\3(��+�uCq���ɇt�+��U�0���&�Z��4s�fk6�o2;��е�is���:��݉�r�+�]�ne淕�yɫ����k,>��b7�k!ʩ����)Z��m25=�ԫg�\���w���ݣOj�2�'���)7�	:p���ZtS�C*l�殯v�m�q�z�8�>B�Z���Y[	�7��.��ء�9]6��B��,>�ȹ��;9v+߭��;��P�s���fj-n܋	�J³���ʿ�2�,:��P]N��I����1 �=�R�v��G�+���le�ʇ^q�RU�jՃ:7Ү���(c�v�0����%;9���Q�'U$�7=�P�6��Lp����"�:���qc�\��䬸L��E'U����j�o3{|����)u�V@u�����o�y��`�f��.x�{��=G�n�����?s�W��Q���Z������kou%�ֺt��lS�M���o��?u�v�W45V�D7�4�\��fUrT)����ư��fs��^����V8Ǹ�7���[��p�mD>Ε�6�Ñfn�_�@��*%[�\�
��똹�Vq�Qk`�w��i<����kq�m8U��rWA�J�&��Uv;Y�1����7ΌY��ֻ����xy���I*����[ī��ݏ�Snw���(t�~ά~�DN��޺%Y瞤�k���kԷ��s[����I�Ц�V|,v���]D�2���k=@l����٪����E�ܟ8�����f��Ar�	F��/"a��X�&��>g�b͈�W��h�W~y�)���ݓNg�:B��iq왞+'z��:��*^4X����}�ka2p��ޘ%�&ћӦ����.֌��q�j�.�l).qWv�H���^>�C�>�r�Rb�I�O����{6��W�Z1�^������boѻ��.�Q	4�S��V���wo��Cxx�n`��,����y�Θ�29u��KR�.��oxt��/��]�3���P(K�e�-c�C�1�k��w�ٗǓ�����<{�^����1{��}�X�Tj����%��m
��g5����9=��ק|c�����~�;a��B8�����Lpߋ��/O����Sە1]�Fμ�]ڥ��ڋ�g.-�7je�V�4�e�]��(M	�ۅ�m/�.�_7¹j>�1��,�q�B�Ơjw/X��ʹۀ���x�r眾�z7�t������r�-F�6��j�pq|�T�2`��ކ֍Y�Ԫ����ʃ���輜���oe�-�\�WN9��]D�ɺ�<w���jfƭM�U>��|qv��ݥԻi�&�{ʼ���S�S���'@���{�g���7���o\�s�Ʋ�io,��nN��HR>�"�si��V���o&��P��J�����Ӯ���D5�ժ�]�XP��!A����.����t��Us�]g����}����<8��H{�[s�r��=�z	�qh�ok'���o��f[O��oj��*�N�o}"�	ƩڎM�4�Sͯ���v{n��J��D�S&cU��Jŏyt�x^���N�];�cYi��)���+�ݘ���=��R�Վ�̀-���Q����.�+��R�g�ˇؚ���oR��-X��Њ�oT`�v���qdlk"�v�\�^(�OMCM+�qݵ;=�~7��%�ۋB�X�)��6ʿ�BS��J��D�5��Tϵt �l�I�zkν�ѭwm�<������1.��NT��mU
�϶f_?};����<��>l�9��ގ��E�4��_�뼪�_�����is.�=���Q+��p�e�6���z��7
�D�4d��+�}���,ـfNW���B=K���Y_%G+䘪mC�7����$�Y�^�2J�dqPj-���[0s���zmWt�a��_i���M�n㥤�r�ٻ�L����^e��J��]���Jffqn��UǫW���.c ���8e��
n���kT��Z��2fǉP��j�w���nPn�|d��7���V�	�7&N��d��}B �sz�Ǭv~��f:/���QoL�,c;JK�o�N'��(���N�I���}�Oz�%{�ۇhsV���h�=����z��>�[U犴��l�����6��Q�T�kTk�o����f]���iQ��z���5��NO9��e)F�>v~fgtSO�l�v��������)^��kƑ^��o�R�s�������S5y6�T8��s�b�T�X������}�n�$��:9�sk����܆���W��8��3
�fX��y�+�orޣ�c�pkyU�N�r�^ʥp1���[�ި�5���3pi�.�2��ư�� �[�%A�w�k{���+o�|5�/d�0���Ǚ��n��[��MO}S���%8�ж�)�
5�Ҡ�)p��k1GU�r�D��u�U�9O0����p�d�t��	X��l$Y�	pF�-o#
t.β�㷶�I\�g����(iBs��̱V�g<1\D5��n�Et6!Uµak^oʊ�!�r�N+�����%�e���2��ysytގ�X�e�S��:8Q�.f\Ђ�������\��,`�=|;�Xc8ԠM0�q/��A�{-T�t-yi$�"��e�\���"\��4n$����06Wi�fd�s��X6��n�
�	���Զ!ώ�AkX�Q޷vݷ;R��g`�׆��
YAH0-3��+{�s�JWk��]�kzs�Sx\�P���^��8�d�X��W=��l�x�njX�w$����&���,͠�;7�MtTt�Ys�E����*<*k��k=������j'�h�s7��g]v�Z�2����`�Ftب�֔X�hDʛ�^b�o����v񗳚A�kA���<e����\��fvJ�:�Y��JƷ��/������7�i,��:{HF��52��K=ZGB�^`ȷ��;�g,�E�����b�t&�9��l�����V-�SR�uK�:{���0�-<7B�V����v=�C�2��"ܺ�����G؁yh�\k�p=Ûg\�����J�N��'��Ň��fE�:a�TE>5��M�8MF�9�������s��x�U9���W����j���B2W	7�v>��I�7�,�]�{��0e���U�
��ɘ;ʹ��-
/ׇ��)"�_ݼZ������6[�qo2I�:���6耹X�Z{��&��W�l�*�o)'�3����>��P�n���3����[�D-f���u����h�a������9\��*�aԑ��]�sr��Y���lT� }R�㩤e�e-�uUf��r�%L�{��c:-˫�ť0�PI[x���J�s�zͷ�R��'��r�o���#8b�76�+e&�Z9u���c��@[�ڰ�:3i�QG�Y�dز�,XM�T5�|*މ�B���)�7�w��KnZ�S	���&��m�U�k&������9HA\�r���\['q�}���VԦ�0o�^�8e�&�n�f�;IN��� �z,Jј,�mr��;-�!۵9�x�a֝�ޔ�[��f���uҁR���
�����C\�}-=���o�m@���"��N���z���J�$ERL4�=���xa�*�$��ٰ'��G��|%c.�������q fg;zM5�������Ko���7>�!�6Ť&��ʮ���������$�Ot�%����0���7*�tm���S
vT�$�Ilxܭ��^C���<^j[�i��}ewH�ϑ�W�F�.���-�G � |�wv/콂�,K���8���D�i���`g��髍�(����fO�<��ۓ(�Iګ"N���s��F��>��ڝ�L}��2�#�i��,$7�g�0l*&�F��:���E���.��1�C��q4%�Gy�%^U�䯝ږ�5pһ�*�Ǧ��rZ���V��$c��b���}]��Bc5g"k^=���L�ΗkPe]^[�oS)&��>�1=��jE��]�U�˓&U��6�!F33k"���4�S4f�Ҫ0X�DV��j���;����Y5P�:mEֈjJ"�Җ��rV��PX"�KK�X��R�M��^3&J�<�����̷VMl	u�Q"��X���c�����L�Z��EET�E3VW0�U��V�B��5�Jʨ����VG!`�L�Ȗʉ�(���4�kZʨ����GJ�H��b��1��T%U�)RV�X���3X��J봱EEB�ef�*樊d�«A�%��l�Ʋ�r��Qcl�J�h�0���k\�h��k5)m�����TkI�\&J��!T�P�ԺŶ��k��F	R�"���%D�Z[[lFĈ�k-(.f��H
>$f�zx�ݚ�j��e��v��.%�ݏ.�V��'� l󱹱B]�V������5݂N�iӷy*�����o<�rur��c<����3���=i#A}�ƴ�^úR�r��	h��y��/���f�K������Lr˸�N�G��w掿��O@��.U�qh��4�]��k%�t�*�ޚb^���/�ʎMu�T���j��ԑSsد3heca��C��h���eA��l]�Q���W�%G*�tV�
*S��L��og���Y"����c�A}�imE�uE�3��.z�<��v*u�H�û�/�=R6��䡡%�\��tV�|k�D^b��z�2�UM1�A��f(B�+�<6��G����9]��!�8��t�`���KV-�T3�iW���۳���'��O��S�5�6۝\29�K]�V�2��csc:o���.I�K���g��*���+�q����g�;�u���?C0��wz���w��E�=�o�c�Y�9=������V����ب��m�A��sB��VW8���ҝ������B��ރ[�{f����|���h\P�\�_5Sx:l�R���f��}<�{t��RqL���H�ّn�7�rdi�ݡ��Nʲ��:7W'���\��wz3�4�F�
���J��_����ːF������ӈM�nMm�w���W��z�'�&�7�y��o%7��Cm�����j}ej��ŤhK��)��B,)'3ki�j\.��M_�[ǩv��ox��Gc����g���8��8�/ie6�d�q�Z���O���,Nm�գ��Aj��&Z��X�Q�uAʥֳ�$�a�*-������Ri-qܞ�ߩ�GoMAG�oIT�nغ��v1�L�9���s�Z����2���e�C��ʀ�ޡ�v�e.�9���QU!w��ĭyave�N�K�e��N������jJi-�ἅQoҖx\�!l�V\�؞�T�z�bN�c��J��z��O���[j��7�9y
�����4��a�����ڮQQ��n������Q��)7�jb�P��V�LvY]��Q]8B�A����sɿU�oCZ�V���a��Z@Ss츒��shP=s �k8zQ��l*����t�����cs��
�Sx�t�hB��:@����#nW[��h�z��V�խ�l[W59���;�쩡�6�boB�|�m^q�X�'Q���S��pz��A<9.{z[CZr����z�k~	�h��V%ް����~�c�j����ӘE"i�%��;��N{���%��E����TaQ��5G\�&nV�G���n�7�ZV�5+���N}�ި�-}qË���b�U#p��T>7d��}�j�˥�-����/����q����s���pԀ^mJ�y��r��Ou��x���|�QM'�K5���3�;��lW+�4ۺ�[n*��bD�Z�E�����R��ZM�q-�t�������b�U@& �/n�W%��Ԫ\�y
�J�e:�����or7;��za��	A<��Xn���1Ӆ�qЦFF��{�>j�F�Oi���&���n'���g�^7���jzKS��p�u&Z�7��e\�ڣ��������+lVhOs��6R�z�Vi*)4�Di������o��6�e�S�^��K+}��|�L
�qgB�^N�\ȭ�bf�8��^¨n@ռ�F�I���p���t�}�m�WX�p`�Ů�ק��{���	[x��#�[ra���R�˹fֆ�5W���X��D}fj{w[İ�6y;��On�)�4��W;$�t�[1��K��w#�]��uUUvfZ�aM'	��>�P�[�z;��_[�4�v�u���t"T�7��!��ˁ�3���Oj!��a�2ʸ\��c�z�6����q����[����3��Yк��'2ۇ�j�yS���:�T(L�Nl;j�@o0mUȴo��Ji�H�e)ޝ��=�*a�ٕ�,=Y�fyv�t���y��`[y��ڨ�{�AܶU���s�E��l�n�ZS�le�w`�e�����+:�p�P趂�}٣E)�]���)ޞ�P��yudG��V�SϹ��]���R��~Q�|�e���=t̙��[B��=�Q��R�N��<�w�7���=���V���@�W�8�{�0w�v|q3k�ur��m&�}�ȥ����9nf�j���ݲ��K.�`���Y�Q�z���gY�bԨFc�#so���5�d���&�O\�� �`W��p����B�l�X�Ɣ�Ӝ�C���!'Q����o���b��X	ˬT�o:�T#i�ʤN��a�3G���pt7"Q�j��'Nu�z�V5��6��6o6��ޣ��bng���ȟC��բ=���&ų����Y�*�tT��r�s��M>�ޡ������/md�Y'�L�j�=%^wT�9o����p�f�-��u�О�Cv�k�wܲGL&X]��d�ISZ��p��yx��pI��[ђ�'�U�K[�ڎ}{�3@���*��K"彙���v��ME��|��7���S�9�\�Sl�͓�t�*���%�ͣ���ek�ڬ�4�Mu��w��r�+k���6���辧wQ.���,�h��`�ܚ����Ws)+#�r�پ̨u�6u����J�7@�i�Z���2�x�G���Ɛ �Y��N�����Cj#R�� �j:� ��5΢�;����ӬX|�Dv��6�W�$�J*�<�����>�]`�5o��cQ@����	�v�Lf���X;1�e7�n"6c(:W(�0�q�kjS$k��&���.W�$loB2�����9��Yjw,��}����}��r��x���D�����r��" 3�-\��H��֕�߹���=�-E�~}P��X+�<�hmi��9�����}��<���r�19j'z۸nup�q�l��؉-������Jx:���;��Y�r��T�㨵9_b�u�791��'ky�݄����e�W�,^�X_k?��d�볗�Qkas��M�sbJ�{)����7��z���Qq^���??!6��T9�t���]C~7�e*־�Ë��{���Mm�|Z�{���<=אzJ�?"q��]E5��WG8p��HyΑ�n򭖫�ݦ�����S}K��P;Nƶ��8v*2����S�a���p�B���vQu�����T[��\�s����J��ح�7.�T�oy�O1��Y��U����z�SIF8ݯ�yJX�Z䫷�{����%�(Vj��Ô:�BR���� .v����w��/��u,�Vl��R�l:]�+`k�%�ZІ��2��!],�m���U�[X�qR�`�|uT�Lr-��W�:M�\�>�OP�6�Xt���BХ��C�D�p37���8n�4��d�
�ȫ8���}�3a;M�V:����G�s�V�.땽#��]q|�rЂ����g6���UC�"�l@��#�DWZ�]��S��hqH���6�o*��at��rwm�C�T#[B���~�it�YRϳ��3�U�Ɨ�ɝ���.N૎��	�Lp���=�"P9��+�4�s�5�fqc�w�u��.{w�P� .C�kW�{����P=��N��f��yXU��Dr�Q�GWɨI�62�ݞ��mت��	��!06�m�k�/2b*�TaLMF(ޖ�r�����*�a�{09T��k�}.�ul����l]�͖e���3����c������K��Y����%����2�j����m+��۠�|�������`m�bw��9���7:�K>����o�Ҷ���k��<u߉�K��/&��~��p^��ŵ���jM�onU��mƼ=Q˪:9�2�W�ή��Z���J�a���&'�1����Z]��B��r�qn�R�oi3�����wn��0'̩b�^�o#ۃu�[�9
�����-hP��W��D���Syf}�����eܢ0��4�9H���'n¨d��`�ٱ��W��s;�M��5�
=���W/���k�TE�벹_�*��ַ>|۹Nz]�s����J��xK�쭔�S����RP�]Sb���8-=��\/W���=�^���X����̒���U+K<����xMPt��<��:�'�]�I�����z������x��<�3�$�S�U�8�e�,>m�a��/���S�G\9M|N���W��^�7G�y��N�"w4�Vf033�5:�@g5:��ZG=�A3��:/��@�~�IwLE�P�s�"��2V�qy����<>|��9��7���Q���|߫��4�h�s.T�CEFgL{�vl��E��}Gӭ�z'ޝ&b)O�ч��;�#,m�~����_�2���r#�9{�P3��o��b�6���{Q���'��>+ȖO��;q7QLMt��,{��3�9��<����T=���L�=�����P��EoxRO�ۛ�}��aw���5���[	П
�OJ�%�P�V�Bj�x�窀�o.ǆ����Q˙c����2��ϴ�q|L��&DLT{�ݪ��?v����{2���M�F��Uv�v)x�q������˴yf�!�0H��
�c������fټ.��r�h��Zt�]�gh:�r���I�˾�R�+wVs�;��l���ݭ�}�e;F4@)fR��мs�r+&t��Y��
&h�u%����V�}MݖQ��@�/��<�M����p���2��T<�ٕ�-�ϦMY4�%�>�:L�ݲ�[~�l�%G9i�u�[{gM�4௢%�=�'���S�Q\8�����;�9�=y>3�_�~�,�O<�z��9�ٳ�\�k}��σ���}��lwL�{�ZX����t]���u�H�}����r���k}W^�9�F���X�W�ߪ�}���Իt�z��Mׂ�o��ɝg�[w	�M;1o}ON���"�xo{�y܁sjcR麟n��1��[:�^:�V�����Q:�����7�od��2���>1��Q+<�����^����8�o�~�8)�^�(�̀``��(	������ϭ�g]e�z��xw�.�4���������9���_�áNQe� 6h�~绎.��e<SJ���'��D����k��W���c#ӝ|�ǈ�1�p����i�y#����D���^�������Uu�4Kfʞ�̈]Lz��;bo�\�_���9�F�&��_��ʍ�;^���*�&m��c�Z3}�^d)�6L�FOa{2n� �����'XgC����®�Ҥ����31�|c�|��#6��-��6`�4f���3D#Vx6A�z�]˔�֌�qM�&f��Z��t�T���	��F�.}���!�s~��N���}�vg��	C�ϑ�O��,�_|��VKy����鱼�'��k W�WS��w��\�>5~���~��}��wp��;8~ǈ��ʙ;Ӝ^��5���n��Ϝ� *=�G���zg�h4�څQ~��y4��#j%��d����o���=�+���QKӌ��o�G!���g��ZK *�,w��=�ڷY5�J7w������LhcL��)c���G��K�����wI���zs�+�(?�+&�s;�z���"v�u�K��'Ei����w%�ڳ���������}XP�y�*kv<�ώ�L��Gx�X�8���������~��<�~$w�����֭��y0:����Y;�e~�c[/o������x��G���\��{I~���@���Y�AQ����՚�{�Onֺי>\���`�t���i��Q�%�;2���w	�O���w��9s�/�����Ͼ���fG/[�{��/��q��{��(��d	UX�je��E.�t�-����fcl�L$�Z6�F�EH��9��(S�V��qupU)�o"���S��ʗ#����6\�TR���*г�8�b�\d9�3�����	�/U^tS�����\�H�������D�e�eXA.�y�#V^���Q8������4�L}�0�v��n�0;�]�]7�>��o���:��Ô�\uy���ƟS�F��]��s�|������Z�[��GǺ��^��V�.T��N��v,�	L�F۶�i��H��זmfJ	�
������כ�b��2���կD"AJ�pL�faŗE9��`����Ȇp���ސU�c�β�rR�ݮ�� J~�߫�{@"��fЩlhH7�Ĭ����� ]h�+����"e�Ub�sۡ��W��Y�^T�ŉ��������!
dt�6���82@�ȱ$��F^Wv��'�y��Qd�\��臷L}��1��t��a����X�m�Q�g�eMG�]-�4U���V�
���Z�K[�|�B�jA9�%}}������ו����F��n,Dv��ު�=��;�l�#x��JW,آ鵛7��ה�1�.�v 3���k8�<��ܣHǘ�V���-��Dŷ�V���o���+@:�:�(������^�$�{��B�.�:�d��׊*
���t�`e��v���ܮ�)jp�u�c�B�ҍ����I�w�L�P;���*&E>4��p�w�.�R��e+	�Jb�8f��ˏF�:�v��=<�F��xf�0˺Qw,v�5#*IO��0%��\���./C���6��ҍe���5��)<�����(�!(�I��,O��$Q7f��pi^�cښ�&��P��]�82��T�k$Љ��b��G��y{|�]�t�M�\e6o*�pV1M8�ٸ�
3��5���
��9����.�f�X�Cy�����\����>��on`��/J��Ň'�h�,G0�\���B�`7�TҶ�w�	[ۨ���A� \���Aa��¼�B�Y�V�	�XY�ih; 8��K,�e����i���P��n��ew�G����{��yWf�@��ǚ�r�\��w��D�A�ondwK��D(tz(m�� v�Բ(�k�;�Ɲ_գo����v��� ]ٸ��{'b[Lb�]����@a��:��:�gv�sչ�&�[[:���T�ۗoD�Ӻ94�Xi��lK��X�y����e�b�;�u�1��4 �@e�8�ޥ�r��`Դ�V�����f�12,&�I����n���hõ��� e���Ӧ�o 2�]N2����jXPmή��G:�6����s-P�t��̸Wk�_N�������F�w����+4ww2����F��Ɖ��x���&+'#�8	{Yj̥�i�Lb�����7P�͊���ϲ��jtf��<�M=�6�\�^���[��i  �>�J�ys�"�ҫ.)Y�b�3�V�ԥ���E�5ED���ʭy���Z�P���J֢��m���-�n��m�օ�&@L��6����U4s�V�7�%��1URմm�iJ#i��-��d��҅�)u+W��	�Z٭QE�m�ضݩ��̶��Ү�YV�m���e�jĮJ�X��KR��-Ca�V��0�J��[[A--x�U�숢[m���j��m�ڻh�l�ֲ�����-���cP�;6��U�J���K��U��*�1
����ul�����JZԣV���Z2�V�8�Y[Rʖ��QQ��s�V]N8Q�j���Us-�
���m��n�N^<�F�J�lg*#mu�J��3���s0�V��-�
̜�31Cj��a��-�l���m���£8�p�i���V�R��Ӗd�+�볮֨��UTyeg-�\�
lk���-�k(���pm���kc�l]j]��η
�DQJ�K(����mLlmh▉Y�IC�(��RD�QG�)S���]bHk�����j��)1��	�\E�vjXw
C;��(�voU�y��|�	�e&vww֜�ms�;��)����<��c�����^-�����P��u���CꜧB֖v����ڙ�$�'�<6��G��!������*�8�/����(7JWbN�"��Uz����(-���ޗR2	l�px+�VWb�!#�1{������n�4O��N.��Ԓ�E{:�C
s���=�0�C�F��:KGُ��H�����Sh���I>��ok_9��gϺ�>�Q;�u"�雅 5;�2�S�}gIh��a���9���xo/�n/-kk�Φ�=T����
�~� �{l�Qn�Q2�a����"�D.��RR����'��|71��{Q�gt��e�Oƣ��W~9����s�y@/z蓱���Rnf8g��x
u�l��59�>�^�E��"��^	K��؆���=�t<�ɏL�Iú���j*;}��d�>�=ǍLv^Vq�Ǥ�s�n#��W�Տr=Q������>bp\���ϪOz��B��W�x��}�%,uߧ��Wד�:ρ�ܶ �Y���S������]�SE���d<��j�&T�=�x��g���G��1��uck1!�]A`��� ���l����r�+�>|
��H��`8Uds���	&A.�̢lH�eJ�:>,҇oF�걓.6-�V.�[���{��b��[����O���<�@����j{�,g�ͭޓƉh���
�2��Ou������j�n�Fa�c;�]�ioy�7o���uo��=��Ca{Eh�Y'N�L��'K���-�)ڥ�4j���&w��q�5�"��j������=�������SǢIӢ��)�:�U�C�#�NvzZ�U��?����Ҡ�=>�̿_���W�_�:Ͻj��w��L�E'3���j�tKD�ve�Gx��g_�>��A�S� l��ޟ#��|LG�Bo�k����ᕾ��}�c��L�R_3,��|M��e��?(s^��L��hܾ�wu>���Cy�v��(o�U �6CR�؉�bb)�D��W���pY��v�ՕoПI�s'��)�w�7O�7�,.��Y+�z�~�(���|O ����_����=�;:<��S�~�Izh��r�,�g!Q��I��>�Ǚ�xN��z�o�\�_��ۛ���Q�.Sœ�[�F�^�^��=�<s"A����\g����W[�9Ģ��N�g�ȫuNJ&��yV��z��O��TvP�d�	��\f�Z���V��S��'cO��А�fN�G..E负�X6�*|fj�AC�!���8�'d���+b�"o�D�����1�V".��)A�SAh˞(	9�Vv��z��"A/|�b� %>���0U-.�v�tb�=;�������Uu�f+��:�Ý��|���瞧��ǜ�L��ր�=�^���D�^�����}R;q7QMVѸ�>��1��I�������g|���4�7����uN��d_7�H�g���u�+t¼�t��/O��xh�|��z���
G�R���<ӻ(�z@:���M�p�J9L���y��6��WT*�BK}��J��˼������Or�2!z���w�~˸�<�g{�Qˉ����1�����gi�4��y`�{j��l��9|��d{�wǉJ��n=�WmQ�H�������')�~.��e��3�W���2�2kK��b��k������N���:�����j������M��q@:�\dҪ�<c��N�+�Uxf���L�ː1�~���Ċ�c��ԭx�h��K���P=�}�y���Y|7�kQ�����𞿪���خ��_�gV��ރ=�����S�[N�`#��R������K;ɟ}�:l����:�u���~�H- ��K	M��0&+�p��ˆԟ9�xl1��o�˞9�:�������,���+��9N�Y��z_����,x��":�1K�U�O�ˡ�6$[��:j��WYA9�{5
�J���bV�:8���z�o�t�aw�+-�_YW*�o���ne�p}�\�T��W.��Dd��fiN.�Fz1�}��p�^�q�-���c���+b�Uz�r�t��Q`B�g���VV��>7rb窧����4
<��ǲ�6r7�\}��^���b��ˀe-�9�i����{8N)��:��B��}�o%�3���V�p�o�ٌ��v�w���S�qU�x:v�j:_���U0_0az�Hx��.���t�:��&��w���ԋ���~TvۡR�s=f\ӻ�^�̂K���G�鉅�D��>�i�%���e�_���@����+�Un)d\[�C�N�k>;���#���{#v�E[�@�L�z�dƾ�	��մo�/ǹ�n��d���ى�5�g/G3��5���^6}�ݐ�� ��Y�%�>l͆:�h��>���}��i�ѻ�J���4�*��>�iب����ٸ���r!�]ǰ=�MG���ܙ�\^�>���+���<�>c}�Z:�'Q������X�F'۱������u�~۸�D�p�Ucڼ��T���k�����?��;s��������Zu���]07���z��az�6����ߟ�e�'z�*zAe��ʼlT��|�2�.�������_���*���%p.j��V6'g�mR3��9х�,�gv�ݸ=�W|�rbB�h�4�E���b����NtǄ%qǙ���7w���s�˧����f��`l�n�෪p�x#�^���Q�����|���ws�,^£\����b���#���;s3T˟O�5���>�H+�T�}��Z�;�����dUC�_emC��u��@�y��>�TF]0O��9>�:1��"}����߼���CGG{M!y�QۙcM�=Q����>����6<�xȧ	��{��΂���F�C~�q��*~>]��p���2#��Vo�X`���Vۋ��LY�]-�Ϥ4�=d�9c]?�^�ȁ������qw��7�\kYR�Fҋ�Y S��(67�S8�w�|}= 7u^b���y(6n�H�/zس��pz=
V�~��n;Ӿ��0}'�D���T�&��1�I����W���D�^/�TE�_	��lKZkjoM�\�q9�'x^�ޟ�v�䨍���
s����'�s*LdA^��	h�T��drK����m�9�O���ԙ�����P�_��ǥ��X#�]̀٨�4* ��a��"�Y��U�K�}�׮�w��{����Q��~#�<
P�z w�*�S�'"e���c��~��`�d��?�^�ѵ�ԓz>u��G�5]��	�X^�C�&�FZz��/����7t��9�E���j!9Mwb�>�6��ZP]�2!mr�J�@. ��fw5�r�Ƒ�y�S'B]�h�dx���=������V�a�X����]a�3�5���l��}�9�e�����j=q�+���g�v=[@?)$�>'Me�P;��{lx���(׾��:��C���EF���e�n�F�7^71~��8�pz�s��ȫ�v���g�,�\������I�9Z=su^V�w���j5΃5�q�d9�|*�+��{�F�דꨨ�S��&���׵c�W.!X����6v�{'pü�i]��f�r�;G������F�fy{2��z���s���eءy��w���Z9�N�<7�{�l���o����ɜ��g˗{����;o�
�Z���x�(�Gz�3ފ�k$�ۙc<n'e��S~��	���S�4lMM��hW�zR����z9χ\j�����N#ݿ?\r7z�*��s��I��=�����V^z�����U �2kO^L�6\��uz�v7��/}S��T3�j#�n㯫�~Q�r��܋7��f�����}>��X{Ņ�U/ӲPj:��x6}�!���z}����7��94�^z��:�����,��ؙF��7T����|Nܨ{u�ϑ�GNmz�ג��Uj�/u���e$"7�h��X��5Z��| ����ʱ�x!y,�fQ�+,5O��d>�{n#2V��V��(�=6�颯:���=nS��T��Gi�T
�s�L06�&-��5x�d�j���!��]�R���+E�՗[b4���0�3q��z%#���#�!� ������rM�w�&����q�x�����~�č$����Խ���3�m�cw��4W�����Pe�!���t��+�Cә��'��<+l�U�֖���Ų���5m+�s�H��q�}�:*�n�[�W����^8Jh��X)A��D�^������[7��ә����{���~����_�½�.}�;ŬѾ׮[���h�z��$=;鉄�-YN{�FJӸ��������~���霤�lN���1W�5γZ�]���D{� ����(��-50�r�LO��m�\��dB2��6�(��p0ו}o�*v��ʊi����z�+�73�v�n���n�W��:�V�&�����UTMz%G>{�W�1���~uE�����/EQ�0pF�=q�������!��
�͌���G�G�2�5q�f����Ϛwu�Χq�����[�8j;�Qˉ���c̾�Whd�X��=�!~�ޭ�g'b4���X/���\�'!q�_TW�Q��U�3�[(!�S�M��G�!0vceo�����Y �%��m�Q3B�:Ƌ���[!��s��
.�[��}��;*�Ot���W�^�3�W��k�¶���A�������W\hz����w#�N�_n�A����P����a��L�(��Εܶ���4�u��
���4�}q��FBl��j^�Z%rt_�ɭ>��X�7��鸉�$�����,O��J�fąѾ�6&�c;�#��3�<�f.!���q'�|�X�3��ɝ��t������u�b��i�C�=��xj{���3��ԧF�=�;;�r�e���,���~5��ɝg��m�'ϕ���w����P���o{�w���|v;ޯx�<�׳����A\d��!��~���w�GǫHwS��E�ݾ�漙���}�+�d@�W��es�_�6��S�Y�r�3�w��g>��뺊�g�*z�S�=�ܿ�=���F�O����ٽ~����)��W����Q^m���OO�I����ώ����_-y,y���@*�ھp߭��S̿t��D?�Cؘ��뙬��;���R�\����<!��ڥ]�=e��0B���Z���P�uZ��zy���߹�O�7.?~U#����42��򉉅���11O��@h�w������>6.h�����zP�ʝZ8^�dC��=�m��L�x���}[GӴ�޹?� � �ǉ��3J������5�-�w ��� ���f�)�&�� V���V�
G�dWM����Z��ٓ�����IY���e�_[�n���\�l�:����h��()���}p2j��o.kK�ه������)�>T��� ���dU�QD�L�-�3a���T��G���>94n���\<G{�^�_i��Q�J_N�F��=�:ȹ����I�9�/{���t�]�̾��{�������Я'Y�>fw�R�m=ˏd+��sd���w����9뺋��|��>�}���D�3�g���;�ד���k���}�l
��{#�"�� aq�>���vO^s�3�,�z?SkM��Cg���ğ#�f�W��f�i�@�wm�js֜{�NU�2�+���,�=���D�������HH����N鸉/��;;��==GX�L�I���<�ל��`Z��Ѝ����8������W{hpϻ�i�Q͉�0���P�J�\������5�G�~�+��%��u;���^��-���7O�z��a�yl�(UL4�{j�u{j�_�����=�¼�^��/ŷ~��>���G��_�zyV+��ǩx�c��R{�%s^�9� J5�;�`MO/I��A���G��h{�3�#}
���'�n�v)�uu�߫Cu��庇�T����#ԣ[��&c�n�5��;N��j�]��.*�o
�ږ���Pq0~��D�|y�z�I�{׫a̵�xY���S�G~��y�;�[�5S���Djms��nm���enQAu8(�]D������ox��G�X�#�Y�ϜK�G�WU� 6Q;�y��^�Z<�yLol�Rqb��G�T��|�+��2c޿dxq�j<�75�n���K��u�V�lZ}t������/��<$Z�RG>���/>�Y*=���.�<�nd�Z���Gj���@w�'7�����g�=����?%q7�'k=g�e�Ӏ�&B~o�Q��=�d�~�b*��[Ŀs�t+�{h������Ӑ�^��f7�=�w�Ӭ�NK�\{�d�� ���^Ϸ��e�֊��ό�i�S����U��"��s�=�S�Y��s��y��R=/��51;c�5}��x}a�fV#�V��U�7P��en�q���j5΃5��c�	Փ�n�N���=�>6��ةӝ��U!��} ��ڱ�(�+� %a!�͉څ���0�g�w�A���`Ǳh�Oydʚ$�v�-�0�gZ	���:pw�{ۘ(d<���t�-�90��F{��O��~��
!�X���(�KG��m *1g���:�8�p8�{����ފ�j�Ò���USy���yԼw&�~�`��TOOuH3�;T<%v��j����!�ֺ����j�{�����	(˵�C2��������F|�Nզ�[v��N��L#B���̠a��靨Z�O������4Bx�{��.m�C4�)�#�m���N���]W�����n)A+�Ǻ��^�y��6I���a��;����yt�m�Fq�M���ؠa���\ؘP�y(��l82%[C+�qh�hKSv�]7�ZIJ{���S����)8;�;'G�]	�1��x���é�pP㳚��J�ެ�eB��m�Sn�-�p�N���t��'�
��#\,1�Ck�"����7x�Z�76�V�a}�Gp��$7��b��"���#e�i�i6�g �3��EZ8U�7������#r��QƚdfG����4B<�ۖ�5�n��2u�� u{�ѽQӫ���l�v�	��XWί�7��9�|-�E#�qR�����XDk�JY�'*"ؼ��8P��wT�wgÑ}ߦT�]���/NM0�FL��4��F�����p�+�� ����-��V˅R{����սEhÝ�o5�2J������F�֨U������@�G6V�#B
^`��s3&m1K+����U���yRNU�j*	L�6p�`i�+ّe�>�����_���&,;Q��7Zh���PX���Wb�[�u�C+��X��Qu�#8��I쇒�Tzۛx�^],����Ba��#b���n]����-ł*��,������z�D����v��e�.�a�U�����5q�#J�b�1�񰮣R6�^s��RA��3���Dr���w1������SI����f�ck�'��[�� &���G�v"��0�+//t�/� �F�G����JE�ɪ�,�7�K*��7wB��ZiÙB������V�0���4��xw���e��F��5f��d='5����m&����j5��6�7n�|�l3�K�n��뾤�5I�WC4��}} r�T�r�WP}B��q-���FM虂�}C9�����"� �8��M�5j��³av�ԃ��Ջ��l<�˙��f6 ���?����\�b���x�:.VJ"gl�"�}+Q�i�Lke�7Q26�fEJ�l���ꚲ�#<�9��3;\{��s�^�m��j�iqn�r{�%:�z̭A��]�L�@������]p���hL������c�Kj0C�{����ػ�۾���XiԮF��.h� ��k�'Uvݫ)-�%(\�U���Ɣ�yۇ.3��3k;DTitX�c�=7.I�c����Y�ͳ!��\�{�;>[ȓ}�C��v��9�1�z�N������J� ��FЧW�����
Y[R�p��v�qH�ԢSSRdF۞3:��p�Lܪ�R��ej�kZ[]J�&j�Zڊ�ڂ�m�.qh��RZչ
"�Dq.�3(��j��թ��v��Tn�ZQ��֖�j5kj*�R�J��h��b����V҉X���sLZ�)L5R҉Fڧ5m���5�)F�De�u��9F̔�-�-mh�eV)Z��J����´U��X�R�,)j��gP�����j�X#���򗖣�9���E�-*�UU-�u.Z�\T�)fk%I��`�k�eiF��)K����ȕ�)�DMKsfM������cj[X�fMZ��r���c��e*UQ[VZ��s�s:�LѼ�+/6D�+k���r�V�3�D��jaF:�#��,��U�mD��0�&�3QDM-s6��j[h��u���b���^cL�X��E��K�!��Z�b֥KJm6�lX��Q���L6�KR�j4o��Zʎ��-��^Z�)e�Mu���*��[�5���7���+kw6��Nl�R�u�m�9%�է�Q<�R�՛n'{W���C��)z��r�IӔ5m��9��s���q�Y���K��7�|:�W����V��}����:��s�2c�r�#��^{L�{�G�>?�Z������ZY�T�~c�����߯��g��+�Ź�*��ޘ�\��'���ӥU��z��?W~���A��.p���{ōɝ~���e���uA���:.�r�W��/�gc����cM���*<}��;<��¸ș�G�S�U0(�>'~oj��s�֙��l�#v�S�󢇾<��ȍq)ϟ��m�R#a�oC��@�;�P��t�pŁ��$ś��
q��kRj�ߟ\�X��/!��7�g��#E{����9E������7?\���W�����II�/+��d�nF���D[J�o�^���B<ˏp��u#_��E���p*������1yO���`h�}n�#pXmB�~9��'�]k�������C��6Ubf�a�> y�d�o�>Gnba:��4�tdA��;�#,m��adz�_�+r�{�,����Ⱥ���Nj}�3��/e��>'�QZ;q7P��+���5[F�χv#Lky~�vMt	��b�y�GԖ+��7^C�)㊸�p�l�=.�\ЫG8Ћb]�qB���5[��I$]s���M����< �Yn��+�-U�]՛y�嚝��Q��:�Z�L��lI�ݦ�%F4��Q����ø�q��8�g;�6s/D�b��f������;���h{|���:ݏ9ؓ`z�{��<�%�3�v�n���V�g������6�NaS�6�RK�J��0y;�|ꏏ��rs�c��DTG���_�L��fl/od�=1�u,ؽ7�j��_���>7���n\?��/�#ΪZ���ơ��2=�gp�w���R����ڭ�̯{�{��g�_ثC��v�tx{f{��p+�z���E��#ǻ:�}��fKR��0*]�$��O����ҥ���2�&��>�c\���l�:�S�y��xFH�ei3}����'W���|�U�jʞ1�/�U1�5������t��찵w���yb�����~l��m�g�.t*�{/���m�1f	H�D����Uƾ�t��L�>Ŭ�����yg���F?FϮ�nB�[���y���xuì�6��(r������nj�Nl�șO��生G{�w��~*{���Ty�j{},p=����^C�%F
'�>���㴺�y�2,W�l)�nh<���z�9��C+�G�_��g����g]�GE��=�C<o����
�[]ob�5������v:���f�Ŗ��Ҏ�Y��6-�����z�U��UbÖ��u��èU��6��M6�cέ�d�s��E�ag�˱>���Q�7�"�qw\����c�����:/#�.�x���Pz@�\E;�_-d��w#[��r�;!��1q���ȏVy��Rw��Zeͷ��i��n�B�.K���&&�Rr	^++�2W����ؘqk���f?�;'��s��F�n�>�I��pF���(蘘^��LS���	h��6H�:�~������{C��������]��P*�gנ<��p@���|̶t�����3���(	�kwe�_���>����(F���k����Q�<�� /{���&���[ַƭ�T��5
��yOd��9'ѧ�}F�J_N�F�?Y���� x�7U���$�I�~g���^x��%����sr��ͭ����cL�j�=p��G�����9:k����M;���0�Q\�̬����/@ݣ��^/
�>gn"v�?a�>���e��ke����`a�⎆�׹y*��h>��(��8���f��0�}�厽r��>�=7�@�k��U�9n>Q�����Տ�F'��8�Z:�<�С>�Z.	�$;>]UDemCZ�huH�V�5ч�(
�V��Enr!
;b�:�Z�l�Qs��=�|�2(�C�`*%�;��s3*F��%f�T�|��e	M�uVCFэ�V�&K� �n����0%���$����SG*w��\����5���y!�����5��ٍP�^&��N3��;��;�C��%�P�X����Z�����w%�T�q�!����ɝss�����wq�߯�s�t���߮;��:���Ez0��!{��=���\҆^3Á��|��L�>����C�wz��x�5��TT�.�q'&��xd�+U{� J5; s���yzN�d��{S#�޴=����;W���|����o�|��6�=q�r�1��]= r���%���+��F�K�V�J��ưzEA�~�����=����~�l�9����ǆ)�����'�wT��A^���Е������6�z��z!Ts�v��p�ԑϽ�ϣ�dh�S����&󞸙���d� P5�������xs�S;��5��~n�o���p�k�Y�8��v�T[�r�ĴH���g��o���{J+q�^���`�U~�'�����_���R��Ϛ�W���s��rVP	Ē=};�^g���:ն9#�4p�>�3������Q��i����,m�vn2ۯ�þܐ=f��񁓻*aB�8�g��ʝ��j�u���X$Ր1��UK(p�*�%�ӆ�16���w{�먖�M�v��D�`� ���N�׮}s@��ר�Ը]�Tȩ�/2�B�u�6t1g�;��{�z��gO�Ո�{ڛ�^s�C�4�̜�*�ZK;Ӕ�n�hM9�������̝�cej���I�=M�5q��^�Ѯt��l{�=D�����Α�3ux�y��P��S�=��rA@J�C��ו�a�ٵ�3��}���,���X�jz�R y,��g�T���ޠ:��<�N���8KG6v����~ݫ��0�Mc�����zy����� ��v��;^�jNC�@�[�Z.�V���t�]�b=�����yoF�X�:>�zP��ۇd�sq�������u������N#ݯ�������`{&��߳��]�-L��y$n����=u^�kK�w�:�/�49�W�Y����ǝQ�"m��6�xI�>>�;����k��%�~���]"�|=N��u�H<��wa�b�SS�7�9��z3;ϳ�R��E�����q����lL�R|���`O�S���{f�&�x�Kޯk��7ѯ���O{ף�8�1��G�LM�N��Γ�w�jO{A�
���a��>ƞ�i(c+=�5�������KG��u�ޯW�B��ˀ�~�1����R]G�3��s�X�'�ӫSH=�S��x��ϝs���u��2�=k�/��;D��3��v�m�7�;��[qaK��f�Η[W��!�S!�N��0���5����%%�L�wK�-������2�[ �6��"vpϢ����a�C��-1�\����WM
>�0o얏�5�j�Wp��;��S;�8&+��evU���>����P�G�+�'} ����
��P���#� ���.��g���OS�GӼJ94T{�N$K�U�Ҫ�
�mB���^]�EE��%CGL^qt���=�#gԸ���R~�="�'�W�W:N9��y����^�Ngc�8�;�:�<M�%��7P��LM5[F�\�wJ�:ǵ�;�z�J'"������urt_�z���)rlG��!y�R�|���C���0�XKc\m��o%mI����.�1П
^�(����,��s��wY�J9s,v��9��0X��c$o�L���x�{���3iq�����ܸ��{���U,��޸j��=���ᚋ>�<r�J��מP|Y�DL���졗��<;9;��t��`Ov�l{b=<��!�������ٝ���+}�v���'����Cn'i��ɭ*���:��Ov��S�����31��p�s{�:+�}zts��*�Ǖ:aB�;��>YLed֖/����@k���w(�shMO��o&�7ٓ|��Y�:�v��� ���U����,�R����/���~j�	ZF̎{-(����n����s7��Al�q�]��A*mH%9�l����l�I#P��n\62�Y����[�ѓV��gWno5� �	���.\��g)h���|w��{ΐ����(��`���툪�㊥���8�^���l�W��[�}<sfcW�iٍϟz��=ޯ3����u����2�(ؙF����ߎqI��N�Kg�@���e�|���:���{N��WR����1jz�=�ѹC�fn$�q�n�����=���+���^7V%���=�=)�����(ψm�(W���P�L�Ez#�C�\f�; r��]
.Z&�X�;��V���M��G���um��ŏ����Y�wI�Q/���Q��A�(�;��ѠK�^��g����t:D�;2���*��G���i/h�F�&|=⋟a8{��.$W���,��10�r�����>Ɇ�������5{��yz������6P�R���>�@����� ��^6�ɖ�\L����rD�+��h��,��=�-�Q��wP�x_ϟ���7W�|��
�W��,���,�����2�qS����lYW��y�^�6W�m��l��K��6��)И���6}� {�u�q��y|�[��V����y�?w_oV���Qt\�[�H� ��{�D<�uS��e$j,bޕ�!�q.>|��
�#+��ۦ��/j�9ՙc;��m)�u`6}�)���3Wo6���L�����̎JrG�L�;�����ς��kC����c��G=_'���n�}1惟}��T)����umw�W�֚�v�+���/NI�;Nׇ댝����Zn5��f�-�x~G�ʮ��fo�d��S�|���{��U��gL\w����KGnv���W��f�i\�:n�zE�����%���p���H�l�K^�Q+-6�_�/�ET<2�{�7���zK$��m�/����VN�5~���~&��N{��θ+���C�w���%Us8"c}��r�R]%~!28+UQ�ɝ����&s�w�ϯ�{��/}Q��{����Lw�qڎ�Y�-�!h�{��`��>����S����|��c�}ON?O�Z%ӏ)�po�0v��tU�1՟ub��,�g���DOH늦�O/I�ݤ;'��hz8GW��V��t��{ʼ�����;����Z9E�n�4��g�Y-�M�a^/yf�Ɏӷ��˟v.�5�����v�Gz%#��#;޿dz�B�
�`����Jo����վ��ҍx@����v����wx��wY�V�d'9ؒ�Kg(���nyʮ�]�wEm�X��p;&a�\���`O:�}v�Q ��PTڦP�܇@[$�Ev@�d�6t�?+�!*�5�i�����TԞ��tQIt�G
:fi,�H_��	���ȗe$t\:�$}�q�,��=^���p��׳3QU��"�������M
)��{ơ���Q>�����g�נ�� �/>��T-;.��}�����I�χq��>��Q�9�;���L�7�����Q������WWG�w�jT�Mπ�{��5jY(����M�q�!���#Y��FX���g�������$y(�n��j>���#�>�u8=䓞s�V���x��W9��O�I��s��`w���p��zo.Z���}VO��vG�'��ՏC� �� %a!��^_en�~�^]���wh�����u=>�>��<��BY���:�jOz@���˱B��Eh���9D�G{�s�^�����y�������i������`
�;�8�:�9ِt�G��EChV�!�S��y,]>(󉘽'����vWT������Ι5jq��N�x�y��]��������W��r���#tܹ�zeY�/�&w�N�s�uz�v7��+wo=!E犟�2x"m�=O��{q��+,�G��*`�]�u��y\�!�������Ж�k;��u����f���B�K�|�lt���2r��NL�t�Nt���� 
���OJ�q�Υ����#�vz��M��t�d���C����vN$�B������k������^Gl{kQ�Ä�n"\�=2���,Y8�>��������'nk�Cb��+�O��5W��{��w"�O��
�\n?m�Y(ԟ"�⩁G��3z�~�({|\��{�|���F��^�5�|{Ձ}��H�D?W�9�A�S��v8�F��;ȉK�� ���OK����G��W��=��#]�F�y\z���r���a��Li�<^�s��a���7]��X� h��M
��H-b�]�F��q7�֑���"��p�	:#g�'����gܡ���\��{70Xu��|\��2��_��%q6ݬ�u�q�ћ�P�g����ҕg�D�s~��DM:�=$d��\���WH�g�pi��:�c���~Z3����F�:��zS�0J���N@^�Ts�x�Z;q7P�'���MV���A�����u�EW,|����V�cUrx?�����!ztG���DϑW7P��9��ǳ�i��W.��{��j4�O���~-;�B�QF��@y3uCþ/EQ�$��e=���Yȧ�Ko6BX�0<>4-.�A=���;�������ŌF�]3\4�󲓭�Vt�]Er�Gg,$)��)�_b��l�b����`��m�mr�i\��ֳG��t�Q�G)ٍ*G`��cI]���0�vY�c����"m��n�u��q�[�x�Q}t)���\�o%qQ��va�t%��gdx9KV�U��3��cz�Z`&c�@��E,|5,V�oA�l�	�J*����E����]87z;!�ם�œ�t�Po֌3<��6�;i���:*�~ɮ��=}]�S��(]�n����Gm�ol��U�LY1�زU��-��㭲1�ʘ��<��n�[ΡS.$,���WV8_�y�w�;���s[a��e�1v�����q��l�N��R���6�������$b� �栭�4����߆b�p�E//�d�C)�-L�R������V���q��q�gP�KH�{�Mӥ1�h1yϴMm�c���G�ոG��]�b��fʏ���<�]�}����b΋.v�:�Wa��jB�ʶ�*b��q�4�Ԕ�.c��fT瀼Ûڦ�j:V|u��{w������J���+���/�=xxU��ĤY:��h�]Zlb޸��烰 �9�����sX�g5Tu8�Z�V�9s�̂�7YA3i�ַ�3w�݃���㚭�6,���[�S�}�L|���/dX���U�Q��5���\�k�z��ncɒ�̾	3���w�榨�[/U�HN�o���&Ҙ�@���0ť:f�I�_�]N�r;��l-�&��4^ʃqV�!�]N�5��9JDF�֫�Ф�c�;꼳��)m�ܼ�#e/7�udT8����(�)����7�W��fg	�X��o��m�����X싮��VR�ĭ8���Ց���H&p"Ҩ�Ac��=[#B9a���u�hY�30�A�1��u�G�B�hW��C{� �s��[Foǆ^�9�Y=W��ľ��P�nE�����A8�y��U��d�B��y�y�1:�r����^��q^��x:�X�N��֪Q�J4�z��6�պ�`Q҄7����qQ��:�,s)1����<��ET�Y��熥%ݯ���][Î�.�Ljm�rW7�K��Ŗk�	J�X��j����T��jF�H�8�g"��SV�;�Z�+Qwc��M��A�[ [Qw[��8����v��w�����s���]�60�c���͌Qv�U����8�P�79h��!���+>��Ɣ����ӕ:����Kn���f�AV���2%�h��]*9Qz¾X���X��q��'pss���Y�XMJF��qS����k�3 �}�qS4�M�-�!9���Yj۱u�.����N�<�a��,��4,�u���`�Im������]-�BP\3:��ʼ�k�X싮���8V�߮�ۏ�2��NA�ppu��#Mv9��V,O_�}�qM���9,�t�t�;�7��|�I��*Rʈ�)��%E��<��a��b�K�ԶZƪ[e��R�����)h�F��3U&�-[T�]��[Z�y�5���R�R�1�e��nZ�-[c�%mJT�ʹ�����,��F��ı(Q�MvF�D-ظ�ۜ���Z7�3i�-�k���qm�G4u*��S�b�aM�J�e-��DN`ج���ԭh�sg]��aʶ��NUZ5�5Yo5e�ڵ��ͣ��i�E�6��R�.�Ա��&L��[r��*��eL+)Ym9�ǖq�R�R�L�qJs�Z���ZUej"��թ���H��%�+Fjmh��G4V3*���#J
5R�i�MmE�숗&r(*9��T��92�m�բ��F�┥+�]�k+�m��kT��.f��e�V�0�KMs�S[J�YmR��)W�g)�����U*aJ��l�TeR�Q��S��R�V���Ѳڢ�F�9�uYmKo9Ex�&�rV)�V]�W;��Ʊ��Vؔ�jW9F��]kFڍ�UE����.�h5/,��6�K*U�5- ���@��-@�B��SHŖb�g�T���Z�'v�7K�[�|$�K7��lj�����2pvϷҬ8��.��ޅ֐��R�'yk�� �����B�ͧ����&j7.��}���T���Q��~�ȥ<�U%�T1�ȋ�6���G�y�O��M����������Ǻg��_�=�z��OVn�����5����*1��O��ڊ�=���ǆ(��c0Ε�>���r7��X0��^^��7Dw��﹮m_y�s�E��j7�Tuƽ��
��;^)�/c&��y3�;�_f�]Qcm��K3�mg���]찲>�^�"���#��F��\5������n"K�z����ޠ�o����gw�P�̯�Z� ���F5���^�^g�ޠ5?m���9}�'�Q��c�� �*��Y�o����'X��p��˷�p�s�u�q�����Ke��_��u������՝�1�V��P<9���n��]����Eb�6n7�\r.��s��"�=�OW�����ה�e�@l�A��׮�-y,y��t�����k�qU�f�fxTXW�;;�}�f<�*^>�p�{-�<���E��0[=s�EңD��2�n=7���/�|���0���
��1��'���v���4��g���J�uyo�Fdg,}gϥ�fFyn��ʝ�'}�WR�U�����@:�چ����� \�����X�7�]�kv��wОޮtQ,)Ks���Q�7h���Tʡ13@ݼ�Ի=���~p��e��J.o�$y߷2&C�j�Gn&&��g��L?zF�V����~�>'���3^��l���U~8}��X�z��nA���D�G�֫�|�f������I_��>���Nv��i��rC~5���W�w����3`Q����ʺ޲.��9��9
��֊�O�gF�4<;c6��[��Q����B/M'b���>�=�w��_M�x&�� �-��7$��Y+=|��a^mhw��:X�3���\'����7ԫmC��n�ջΨy���>���[������7��^���v�v�?\d�_�:+Mƹ����G�ё�p��/i%7��Oy���Ր�|�U�s�C�}�ʱO�GoxOi�-;0�r�ō��D����ѝ���ސ5�Gm�+g�${�/�Kգ������Eh��	�7%���:v�
$w�(�l�[�Gq�β�_���'T����c�4�_������O�,�g{M ��r��:��EX0�(��+�4|Y�L���tx<UP�2g}7����uQ����=�����:*�'�O�*W7v4��W���A�}P��ச5(�1����9���=�޴�'�t�j4A�&�jզ�v}��SF�su���OӮ̯SZV���(d�:V=�μk$r�`���
��:^͚��D�HN��,h��hY�S��5�Ƒ;�V�76�9WB[����,��UA�=2�Ⱦ�øݪN|7�~7�W�Åν��=���_�����=޳��Q�+��R�Ʋ���d	D���T���^���{u#���L!]n��+�.ѽ�圝�
R:5Ҿ~�q�Y�dB9E�����9O�F|Ke����ɶi�zj�-k��Z��;ևy���u9=�dxa�j=qf�%��-Q�G.���<v���^�mϥ���9�+�ُ�
�v��|�ԑ�{���F�[��x�<���qwJcP���u3W�˼%�zdF��B�����gB5�����>�^���W�� �.2[P%��]��fיu> %,��}3��������"��9��Ӑ�^��?����ߋ��~��G�9S�<k�`�t��I���@+^�$�[�&������1��!���"�^ׇb2��fxޟf=��U��Σ�}�V�Lc��7�,z�{�d�gļ7'ȣS^Vѓ��MG�}���of�3>�)f���}�hzӫ'�zB��~tO�Mt�A@g~���م�g��u1�Vɣ��âv�����Ŧ�����9*[�es�S]��I�����k�5��p3�.�Z��Z�5�a��,̥��\cQ<<ރ�#�;�&���D�y4v�f\N��"�Lco��+q��LC�&W<��=MZ�D�D��N�&��b6�(��KXnK���6k�~��2�W=��
�+��cUS�'��O�v$_��N
��'N)�y�B�;GF�zqY�[
޳^����8�a�ڭ7��=7�l��x�~�e^�j=��Bq�e{�wh�Wx�Gh=d��}3�:X��ۅd�\�`g��k��k���̋�MnK�L�n�� �㾦��폕�-p�`a��b��������L\m:	�uz�r����r*<#_
���ǚ��T�����{]�g{nQ�8JF��s���Sn{Ō'_�s=3��nx�{y�7�	����l�����~��n�\m{�<c���5'�T�EShf�W
ے�}�������}������>��z�o��:���:�u�����rLϔ��	�$�eL�2���;�Q�������2�F���[�\{ ?Sg7���N�z����.����'0k�^�.�x��MA<��W��nP;���luG#Qm+��^���B<��|�^g]FٕouMR��;��"᪯Qp og��,:�UB��#�Xo�S��7Q=���"�x>?{6�F�Ti������F�U�P-Aܣu|�j�ؒYۋ	削�sK��%�SɶI�FKz�)�5��
����k�w�=�+w�Ɛ���+���J	��ts�^<&��]L����5�®R&�d���7��@�E��y����5�ݻGy�|����㳨���OmN�uNJ'$�z�&&��4�t�&�#"n5xӆ%D���>k��ϡ�Qǧ�}��L�pq�nA��׉D�D���M�>���0*-nyP����Lm���%v�Gt�݈׆�5'���>t<�#�S�z�����?
@�ϑ۔�|^�W�$�َ��8�Xx���My��
�=]&��O���p����g��E�2�����´Q���\b���Cb�wo�,�g�49��ڏ_ٵ�7��3Q�p�[˯�ΪYG>����π��c�jY|�gM_�{N��H�o���Zn'e��NQyU����e�K�}��p�ſ?z�8������e*�:Nq}���Qð���7�Cnv��3�Y�+\����x�y�߄[U��1kyj���x��V#���ռo�U�\k۞0�ñ^)�/rkK���gb�0�k<��C���w_X�u�H���;�*����m���E��)��^���w]��wWOg-A�Q������v��GM;1�������{o����4?a�;w���÷6)�Ny< ���j�uZ/N��]G/�ᡃ����[�n��J��րЇ�W�3#u`Zg��;*m��m@u�Φz�dH�G$=���c�Gh#}i�D	�q����e(�������;�Z'\�u0�F>�R�ݜʾV�I��O�韫
	ɘ�ʣ�%2�!��?���Oz��#Ų�7=�!��kS�N^8S������,��H�e��C�%�s���b��y)��h{���=�z�5	cC�⨹�9r�ڞ��u|��7���)�,��@l� r����N��w5�
R>�p:�Y]��I����c�ur>�f=~�d{F˓� 6_LL7V��A+�ayu��a�]/����ݫM���~�U���;b}3̠����s�{��w�̉��sp�h��L/�O����f�3.6�Ӳ6�9�tL{ݕ�9�̧���,z���>��U��A^�`����PC�^7��,�%jR�DL��IFl�5�f�2F�e{�hޗ�ݐ�C�ߌ���k��|�,sX W���۳��2v��J�����x��'I�L������͢�vN�����Z��������f�B��R�����M�G;��[�}\M�>.r���H�ܰ�6�;�����zL��,x�ێ���g�2@Ȝ�<�/}НQS���p��q�y&������"O�۝�כZ=q�������>����vd՚���s.�4��K\UH�g�l�ĴEswHA�4}bRv�݊/e����K��4�m���]��w^qORP2z�Դ���X&�p]u���'R=��-�����:n�hiWK\Y��p�3E����ul{]sǻ}W����Er��}mP�k���O;�r;��\Ь�{l���'���Z;N�<��?!L��TI~I��{f�� b������H��_ޜ���B���Z-`��3�{mόj{f�{ʽ���T,5�V�z�WY��P���c�5��M��o�]�uy;C��g;���}}R}AV=<�h�<��n&|0��Q�x���Lϧ������w�z��=����wzv�r.�z缶	Z�=�л}|9d�<�D�S>��`_z���2��>�~-W�Ǣ��L�l��ʯv���g%��L�R+�''����CJ啛 J5�z�S��n2Pl�<s	��=�-�18��%[��`����w��y��w~�qs~��t)��[+Լ�8�ޔ��owp�Yl��b1Vk��3g	������`+~�:<����}�FyӸc�
s������\_�1>�뎖 �c'jw��c��U�`{���-cꂔ,xّ��M����=�F�yj�X��Z�}���Me齖�T�F��5jh�� 4s#P�m����W[��>��T�^�2�\Z�$��ƅ�ZOzX̀�!(<�_=܀�5�*@r�rweMRR�+�u��t,�JiKyۀ����iY�X�fl�7���|�F�-ʼwxU-�뇜�YN]A2"�gR�u6��<����^NK%Z8�ߖq��ƹ�Y�qR���+˶ȫ�S�'&X\n`��TD�N{N�~9��L�+����y��7O���͕ʊ��4晓�Q�e�j���l�4v�鎼��.V��|y��y�&�c=�ئ'#��mw��G+5���Ǽ�{�Χ�<�O��+	�&��������k["t��^�'�x��7�W��N����{#>�:�!���\5D�Vr$�;(<���8�r�M��s{����{Lz�6���O5�lQ�Y���󪖤�z��{.���ZRQ;�n�r�}�Ə�:J�&:Ϣ1uC�ڭ7����p{m�/V;�9㈳5���=�<�����]dv�����<�kE��:v�g����2�2��_��Vn4�7�q�|:�5z�I ��.7��n<m*_���O��u���ޫ���m��Z#0ϗ���p��i�����X��yW���]�ϼ��7�cN�>�W�_���{�ב�[E�<JF���T����*b���#�����\y��>hz����\GS�ϙџ?z��l_��۬W����5ה�H������""��
4k)�����l�A��-���y7�;zn���6�g���s0O*�z��(�vN�����ԍ�^m.΂�z�-�����'0��,w\ L�vOeۼ��Ӽp�,�4,�]�l�9��no�� +�9]ײ������̓�3�z�Aj�x	��;?���1����9S���3�<�z3|�6V��îU �6C^��^\H�u@ЩY'�_xS��'q5�"n0����#V������Ac�{��3�}C�3�`8�gt-5T�W��C�X!��t���B�t���h�r5���%1��֑O�v]�Tׅ�i�>�f�c�V��Ϥ����aժ��7��ә���V��6�L\� ��8t��;=I���%��t��̳/��K'=�<ʹ���VDӞ�љ[��y�z(�������)�[^�_���m�/{<*}0<��3��N ��{r}n�J&�KGn&�[q��=�['���]�I/Q1�vңj�ǐ>�Ԝ	zi�}·���=@�Yy�Jm��tӲ�2P�y��.5麄�wz�앥��s��v+�����y��]P�w���&���J���P��$x��:l���h�d��m{��|L����o.�;�:�e��F�b��;�ti��W��Sh�j��~����|�Ǟ�fQs��q������`������=�ap~j�+�?���bu�v@С��O,X�y�|`�H
�a��ȝ��X��M]S앏�T��9�f�nrt���N$�������7�7�Tר:���9�hf�9��(TKb�5��/d|9o)Cz=9m,�Ѽ�d3�G���ԁȼ�Wg}�Uüs���uD�G���W���.)c������
��������>�6����>G�uDby�og��ռ|�TW}�nx���;��>Y�S�ĨQ[a�f���h�1�$ΛN��@k���]{ċ�o���ź���e���F/0JG]�L9�c�1>Q���2����_��3X���em�'�iٍMz��7��w/��_ʲ���
�8a���TL��m�9�>C=D�������P�����
�����ʣ�z��#}-��r�{70d�ǻ�7K�l����[������b���c�%T�;�!��M߁j1Ղ����dz(M(�9�ܱ�r�YI�>�&���ת��dt�}�������] �D�d��v�:p��7ۋg�J[�ֆ���v��/z�1��T���I�Q�p���X�0[;q10�EҢ��HN���W~�i3���#g��wc�����hM�'v�X��}#NN�Q^�n; 5�F߽e{�Fӟ��t��C�&'��KNA)�&Bt�Ꭶ�����{������>��!$��	 BI���!$�Y	 BId$�	'���$�Ԅ�!$��	 BI��$�	'��$��!$I?�BH�Y	 BI䄐!$�@���!$I?���!$��@���HIO�!$I?���!$�r@���I '�d$��b��L������ �h� � ���{ϻ ����r>�PEUJ�Z{j���F�2�$Ew��w�*'�5�ܻ�;���V�յ{���ޝk͔�����ֺ폤UQx;�x��^���4��eW�½uz��]�����:+^��gR{ơ�Ģ9w6l֭mS�    ���*�     �B*���F�  �  ���M       ��@�J��� &�L0	�	��ET�(`�� ��  D�A�L�4i�oT�h�jf����][* ��%�!UD��4#pAB()e?""�%������g�?���~����ED�@�ƀ@S�F� �Dd�P3��=U�.������J3b��k�cwIP;��ߐ��4Q	46>�<��[�֘�Z��K�5�B}��������_v�S1��$�x�:��w����m������+�T.,ԣ�Xkahk�yf�5V��[�t#�Y��0����x$��B�0K���ۢ��{r^:��.��bO�L�f�51;ش;��Ce�T�����D]���Ma�10��ϱ�YQ9Gr\;�Yœ���\v����X�x�g���NF��c
]Xԙ.�Rf�wT�Cj���I��M�T�Ż��nZ5(��%E�B.P�5��32�U�P�����]��f�,��᭤��Y��ڇ���7NΌt3H`�1
�W+�j*;���ų[v\H�׌�U1�X9ҙX�TզV46����E��R�$�޴�,6���{����T���{�ND�UKTTx�K�.�)،=�r����t��,�X)�&�7�]8*�[%ˀ�ChU���R�vV�ѕR�I�^+����,^�5@�`�3�>Fn</,d��H�q�$�L������AR��;�
�T�ݤ��h놆�Y��wt�L�D�2��K�ci����5�,��p,��]2M֠m^3�B�-�X��	�¶��Ʉ�ʡM?��Ie��
�e�wT�
�8z���;���5�H0�i6�H2�GO�������C+/��Uv"h�|���uuM�ܮyZ���$|ݹ/���o���I��=�f�W$�+�Q�wl���*�*ӜMZDt�|�J�JfL���͝eJ2I�GI�/�v��܁��l�2��Yk(}�Rڜ`8�Ng�̋Q��@�}�(j[;��-���p�ݽ�{}ۈ$6j���2�.��Q�օL*�#���k�����-t����N䲊<Vꙫ�V�\�H*j�m<�ԦD�*}WD�c;(�Pv�#}N���x y��nQ�P��,XR"k�ٜ���dv��x��T�t��f�vB���$����F���y�I�Ǚ"�t�ÆgYj�>%�i��&d໲�Q�OZ}|��p5��v�bp�T���f[� �];�55��͙���nti::2j�Rꡤy��T�s�ovv�õ�yNw-����o̵
��.�v�l�0#b3�TC�;sf�5��)nP�"�u5���_L�]S�iFF���ME�f�w�;�$X���-���޲�btV���!��Ny�՜E���@rkJ����#�x�N�ǡ�����Z'�g(��;��h<��x�՜8���;��v�3w�Kl�;����ܮ�z�yJ�jXo_ήJ�3
J�\��'`���}߫����yhm��+�:>b��r�!�-�S�md@�M3K �'a�#����~����/�� g�[��C�/DV�x++n�-�:�g8�
�]�Wl���r��)&qVڎ+�7�̖�)�TF��m�v�Sg=}E��X��wF�`(�]x4���v��Z91��b�NA�R�ydN3@԰��@E���J�]���ҏ�o\{��N��]�+^�RO�T=�<2������^���$ �Akjgp��#X{�Y�k\%^Q�Am�zq�k)jدKj0Յ�w�&�-.��"J���fv���[p)k����M6��n�G��XЩ��Q!�UH��s��;Dvތ�z�R>W��/�MpG�{��EBe��dn��D��N�f\��u܎�A�]�HP��غq��\��X��'�2@�*�ͤ��к��(�|w']��E
כ�ه����r ����e���ր�q�\W�i��<�G!%.s8W*pwV&�4�bbh̸�����c&��@�B�)J�˺�
h���̣x�T�Ӂ]�c�8�EI�bi#(1���ړW:gM�SOy����������3\���){R��dv�e�g��K�xH�;2ҽ�i���thB��y�4vdr��d�vѨ�rs��W�;dٛK��Z q��ukU_ձ�b��%�lm�z$I>h3��w9��q��O|Ue�Y�t���m��,"h��I�I	̋��eH\��J�p.�ն%����y�cʆ�X�{��J�����x��&Q%�P2~tT$��7#+�ᱥ|c"� ��[!��Ia ��$�	r ���1��,�v+������ŉ�$z$[آ��fiC�׳+%�61��l��}W,��}�gO�2�/����s/�(WТv��7��[r�k��̿n㰌PMw�̣�4��v��:Y�4R&{��++�R��6,Tq��DE��v`O)�w���BV�
�Wd�&���(��Gx�ǲ�f����))g���V����� 잶�/&�p�ң��u�{�W���/9\��xu*�y�z/�v�[�MNa�ρݛ��A�(郐�ϭiF{GA���5��*�]z��*]��K�����Ve؍�*ۮ��.��� Qy΁j�DNΛ(4���F^�Z��a#f&o��ۭж��Y��b����4wZ��Xl�OԼ�Ռ0�Q��v���=U��U^�$m�P F�睇�^�{`��0�=lu����s���K�]Ϫ�e*D�s(�	Eˋ�2�}��������9���L��=�� ��[R-��\�X ���e����G1
Zǟ29~��o2�E}uA+��z�v7�0m#+��Ղa#���fQ:�E�SW�c�_����v�������n0����Ț�Fs(�'z@��#���}��sG'�{�`�73o�.3gju)yZhV�z"�!�{�J-�<<[�N$�]���Y̘ː	�(�&b�I7I�0j�D��N�˿.�A�,�%eǋ@�T�ԥb�R��N�����HH��� C1)NB<Ȝ��9��!3�h[��A3Z�)�{TY��xY��)�I��i�i���G����sX����"9��ۛ�EV��f\�=��{�Ը�Dm�H� γ�<kw5,Ty�Kͯ:�6�{^����5͵���e]/Co�f5>z}�֕�^~����צ�냬���D�v_�g	�*��]�������Eᮒ8@� Lٜ�ROWj4��y�䖬O�.�����=��q�m�M�P�s&n�F�A�f�fa���-�����@J�"�`�#��/�mB�b k�d@b���{����ѕ����P|H Ā����o[�D����JQ܀�K�0y1υ�	.���s)�	2��`�������܍�az������F?0!b�R�,��k��`��<Q��v��=}����w��Nӻ�Wׁ=y{�f+"��F2����gvr���F�-F��n|�xc�\�I�	dYLg{�n9�����iF{h���&���r��O�*��j42��^�V�~q<��S��VzWН�;�G�_L����I牧�9���m��Nxa�h���&h��/�A>�u�AS�v������5�D:$D����@�=���De��S��χa��-�W�g�|._�X��>�+�`����X�Dr�5� �Lp�=�=�kNIG���]J+�+�__b���05��VJ�7�LP&���%�L�K���겮0�Ky�[;�O�콪�a����1NQ�P92��)U��	4��f�r!�I��
��P2�#��5F�k
��ӞO�@��C��)�*�1�+͔6�
�+
�e8�׬V�6! �^-�q���˜8�$��.�=3?u�+�K?��a�>�GТ0�}��_e\����k#�k��}����J��)M�w �ۅg�Q�W=��q,_h�<iݜ��O�Ǣ=!��S�e>(���"�(f��B���{�Ē����b�7�}\b�'��;U�w@ܽ$Ѿϥ`g����"�:4����)������K�fC���S���(ϲ&���8O¦(�t�!��K,mH���T�]ٷ��9�y[��>��_>i�+��]�m����\�-v@�K�Au��^#�.,�]����s��c����K��jߑ
c��1�6M��ж����;&!/��β�5t]R��e�.v7suj��f�7�ol�=��i�� �����e�:(��sp'ኙQ���{�T��ɕ��y�TI�|���A��oGەﺧ_:�6��\T�U�zgk"[�ģ9= _��aћ������闼��[x����ǽz'MF�ת?efӝ�.��ovnv�����)�r�<c���4*�Mw�k���<�����rL�?�vsI>�����{sD[�[͜�lhO-�y.a���4o8�K�\�m�U7�9Å��8ˢ��!��&�ne�StĦ��}��O���z�t5$]ʶ�}&�� ��bJ+ �
���ut�-"l�ȫQx:��I��P�9*Ke�x���[Y��n�Ū���CK6uNfle�n�$�.2��$Q�MB���ߎ޼�_�Ei��U"!\{���%�juM��D�oJ���5��\#l+}���Uҏ'z��r�(>l�> 4e{T�ӛu����1:���<�@��1�̟4E�8�����Ѓ�>���l���/MmM���`�g��wZ˘x^�U��ֲ��ꢮĞ3�/�7�w�0f�	�Z5ѐ���=q�&nj	K�G��<�y9�{������ԭ��Z�b�3��dN���^HB2}���g�F�(���3�B��k�a��ܥ��������g��fq�N:��n�.j�=^�׭=r���R�ӓ��8Ż�RFAX�R�����?��k@�$�1-39��s��$5����q/XZPq�-�o�n"O��� O;��庉{ZDM�����[��
���!�n��đL��v�#�1-*,�mn^!��;A�쮳�+�Y��/�i*��@�) �N�7�Ҷ��T4���Q|�ȋ�����ff�a����pF�do�H�S�[����d�8����O, ��X�L��A�� �DIAQ�6��		Xf,���K�L_k�Dl�,B�yl�@Q\�s��|�/0f��k36��)X�6�D�C�����
�[8������6��3��w1��CHH�����K�1@�xf)h��a�,p`
,4�r/��N3���R�{���3f���c��؊"�d��m�4�(��N����J�k���z�G �X;�u��]��A�z�G:\�c��}1fǙy������=��fn�wO"ނ�G�16��S�3��ۨ�3�k��U7�Lh�dA#s�l�Gm��	��e��]v�Ź�e�8l�ŮiyS�wkm,_30qa�fYu�H�,� Td��i 7 kne���9�`Җ�KQ�m6���$M��@@�;D4�Z:��!���U�nP!�8 ,j���n2R����V���7����4ȇNb-�&c���
!@� (����8����{,1R�"c:�t-!�
���F��ȆdY��Ŏf�����]4���[��qo� �[ x�bA#v��#��`:\70�oC�AaIق��`���2js׾�O���-L�ה�����L��ˌ}k��	�?�dL��xu9�{&w�纊�I�����2�_��B���8�;��ĳ|��+�|�4��۱s�=/��N�d��y��
(�$��ϹR���>��H[[�v��/�>��lr݃�4�FO��n��b�:z�d���B.��,�%⯷��m/3����D;τl���]�>��*Y�:`��p$��Xl��9sY{���|�	��B�݊�>uh�Q,�}HE��gr�>��-*�:�]ڕ�K�0|!�TǕ����n0�\_������\���������30(��wf�V��]z;g�h��U~ˮ��,�s��:`��b[�V�wq�={3��\�E��8����8�IR[̼��R�m[�5��{د�*㦹Qօ�1><qb�;�����s���1I#:�j�9v��;6��#LZ�l�{��F%��>i�n�Ʈ&�D���U�PӮ���f�jv�9gU��iX��"�%��e�i��*2P��Uz��E���!ɀ]�$�"�{����~�_�C��C��R��\��4�%憐+~�����j��sҫT��^����x��{�Lf���YM�<&�V�ǖ��.�-�?!i��`,�;z�)׳�G�6Vz�N|�xB>ξ��<��7E%���
�"������P�σ0*�s7yE��#Ux\t���E�k��҂|�h���W���ʓ���}��b�`�;}3����kӄl]��W��5<��O(��d'���.H�;��]gf��� �c}t쿶G`�k�']ʋT!�=���
׾�j�f�P9�kJ��}}G#'7x��fh��窐��]�fBB�B��/w�lD�ήy�������Vgu�������4�11y'�2h�7~�N,�`s�7{*.�=��Yd[�M,V��  >��z�:?�rcr�c�"����1��c�nGrh�}]>�Uy�{{�`G�\���c�c6��?�8�u-�w��ܢO����x9:Vh못��,�I�����9���>�O��A��W0��F�s�g�ؓ���sfr};��E��ce
��ě#ٰ�&QvP��:JV-z��`Ċ̩��P"�-�F�8��G>��RqF��b��)`"��D�$$�$&d��l/��{d�&]e딧�U�`�c뻑�q��VN?����?č_kg����A|n٣ԾX�1��9�������cg˟�o��K�9���
�.��-�rwj���]��wH���ŉf��`"���(�
�yװ��\�Wl��p�>.��t�>����%�o��t���׻Z�R�����>x�l�(x�>[�lz::��=8�s�=q�_eՍS&�}X_�PI�f3S�)�z�inoWm/33G��'S�P�\"1��1-��(p�,�es؉������=Yᐉ���Nq�s*�!Ҵ���}~c��"oB7�A����T�"9=,�q"U�����g���а���j=�h���S�릻\>�L����a�\�Ѹ[Fz&�
y�mnQ���&���f���"	�rA6����¼����C*'gj����a~X������~���P�0�z��dZ���d������G��4=��K�2�'j{�U���p�O�+��iB��
n�O:��m�Ӕ��ܔ<��T�\��7���b���骝��gS~X��a�xb��P��BI�#0L�;�N0��v�c��0��cU$����}g�|_S�$Z��Ass�N��3u��OL��u��v��2�ռ2�h�"�3*�X�E�P�3S,T��m�Z�0+/.Lf�,u+��(��y��I0Y���d[-���u�L�%�^A;^���]w1N|��w�D�o��Z��b��D�޶�5�a%�=[��������!@e.�eM����y��@|_'��>���{'y	�]��O�8��y!�i��Q	����j��
:��������L�j?l/����Q�I�}$���th0������7��Oi���v'������wgC�*p`���\�rb��M7��*LlY�ƕ��`�y�,D�&E�w{G�!S�ef����} WbW��ڕ#�V��{�0z��
kIHcP��|�Fn����B֋3ض�䴧�t�מ�B�<����4ҍ|z�sb���S!�j��f�t�8��/u���hY��3*��I4�]B�
i���v��]+^LOv���+3������J=��7�sUe��7܅vf��-��P��0V�W�6<�)^p�;m��x�������շO{1Ȑk�q[dE<��◚����dAZM)�ᣨtQ����.���^ծ�ǖ҇Du��5�)X�G7;�i4���)iz嫪5K��y�k�!��Zk9ƨ+L!^��5����5����F' p�,U��P87�݅�h��Sgm�ϒ�yb���;3U9�5�Ȯ��S��ed
�pS�fa�ǲ��t�gJl�5���ʻW@��tк�4�"�A��.�]�xx.�L	Ӕ�a��XB����d�~`�҄@KK�X6�*�#N-��'W�����]�{/V�[�'��y&�`[0�A�M�Q�u��d�	ĖHvK�g����Q:�')�Go�^^���;8a��6���{tq��R���E��n�k���\q,&����L`������˒�1k�E�9y-\�ƻcJ�N7�d�8���}�(�+{��v���ݛ��fy�ko@����p;�_{��gl�}M�l3��r�ҭ1;�[�ht��u>�߬�<���|�<���k;,���k���KH��{�(���@�������P.��Hkn��ƝR�N�e�n�i,�V�%+��<���<��i��Lw��T����T�?�||/�7.�g��
|�Ct���{>�穹��ҧ���|f��.'��臣@�鬕#ov;ץ�OB�L�%I��ʉ���	��t=��z�#���D�Ϣ�g����U���έ���*ז�%�b�ϵxP�H>�7�@WSR�Q�I]K*FyRD+�h�R���^�<]Vm[�1�P��;��D����C=�v*���Cjڽ]����;ʨEsK���FU+�s/�v��j"@U��y��H��Lњi���e���
��X�w)�)M��[�ox�N���͍��J����c�"�ɷyz,�}�b��_��U��B6�O�]�����f�Cmn������B�$�~e��I|�	�,�-�Rbd�I�."�99;/v�''&���t����2$�eF��}[����o��({u����C�0[N �������~�t��u|0/�!zmOV�	L��=�}���-�ZK�i,qڭ�P�o$(��+C�ۼ�e�����qG�l	��$;j����b���*ٵ$��5 �fqY^l&���C'��'�D�ɋG^ ��W���&�8u�DԼy�~#]*�#u7Re!�wu��e��,���xx�[O����\��[C����+^h�:Ohi$3�u���m�%m3�'g��Q-A�6mF�ݺ�γ��'>}m�חS�_M#:^ |��P�:il�`��e���d_9��A0�%�.�-��o��p�yw��� ���:�=�y�ع�mP�C�,0j$���ތ8�,~�fe�n�v{��q�=;H����]����P�Vg��=/��,�!0��.#s��Kj�fm��9P}��t��)�ORD���ʸ�$X|8���+�޲�SƄ�H�K�*wp����~����i�1� ^E��5�\G$W>:O؋��]��̾t�	�oc\��=�Y�HuQR��I$�%P��ZQ��
*'�ܔ�(������~%S�Mi\u(�g�E�K��}�k U�pŋ�X�a�����!�Jx���drikz�:e�"�{H2q�@�t�z�?^T�M�xn���c��ֱ������Pi��c;p�PӘR��tƍ��QQ?�o���߷����آ���AȞqQ?�v#"R��8����;(;�W�dj}�Q������=f�O����(����|����� �����l	����-���L	6O�V-��{�W���q��y��s<�Y��V|r�5o"��rXQQ&؛��֮����	�ED����l��"�`h�X�ZE�[����uN\�s��TN.C0J�3��uE�����t���4�_�/�˚��r��������i�������#B�����^a�NY�O�wx�G�c%�����:����Ͼ��^F{<�L'5����������g���>N�I䈨����_��d~��]\:ؐ�ҍ��>�@ )�Y�TO������8�4T��a������h`(����?�� S!���HF�l؝4�5SDP�\84 �GXd07�l[}�f�*��M0�C9���J��C/����.���6���l/Ru�*$���ՂN�Ǡ��c��?Á�3�Cs�?�@�Kyw��>�l X��������>	���)o�W@���
DTN��玓��'�*�W����=h��K��g���?O�}���?k���:������3�ЎE�Q���!�i�^\���>^�3��}�˪O���5������/���u���N����]�2���hC�g�07{!�G�z�]Z��A�L��:`�EQ?��t��OG��t:u��(�'�z���H��v������R!�-�g�����B@{BB������rE8P�����