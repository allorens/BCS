BZh91AY&SY�4:8ta_�py����߰����  `�~�  
�U
 ��y�hh *�'�B��x      �P (   =(    ���P;��;�A@P ���ҹ�����=��m����q���跛������vl��;�{��m�}��>�{��;o{��zݾv������n�|>��֪����>گ{�������t�[|   ��>������������^�s�W����K�ܾ�z%v{�ܽ���n�j��z=�mm�z�}���T`v�k�v�X�T�Z9O�N�Um�2�����+�g�  ����4���Sm����C�}N���oMWn����gV�3�{���>����ח�t�î��罗[�p�VC�]������׻G�   'a�s:.�����p�n��Ӿ���sm�Ƭ�у[�e�v� 8���{}�&|��u����o��|��ﾾ�om�wo}�� <   "�}��m�s{��������]���w��޽�r��u�{i0�R��������]��V�}��w�ޫ��o^���v��      
          �      %S��=J�R #  4��   j~�D��!�0�� L�	M��jUH b`	�2a i"�R�L��h104i����$�ELMM1'��O�����zb�����T0 &L � !�M�x�y��*zQ
�H����ق� ;�� U� (������􌠢�p�ҩE�������B� x� ,aH�TU$(����[ 5U�ɠ�	�"�`��%�H#�A�AA5�C�|��}�o�����3bɭ};3��4����Q$�
0eaxs���{�|Y���p=�t�D7<8{�n:vg�0�η8VSw��v۵6��eA/"�"- �"-=,G�'��{����D�7�+�ݲ�K��6�<�0���%��Aq���0;��	��-/�#�Dt��Kb8'8���x}?{"-"Q�����y8�q ϓ�<���9��H��D�؈L�H�8�C�$`�f����%�FbbaC�#�e��y�(Hn!ȉl�9��� �����#�*3�	c~"D�H��=#�aD�8B"%؉�H+�|��}HN���1#
)�#B$s�M������dtNDN�#�DOq!�ď��=BbY%d�C�>K����L"�,D��0�,��D�"{�	Ή�H���(��|�ap�$"O�;�Y#�	����Ds�<p~�"_��D��VP���G�HN��$|�E�`����B"_D���Ύ�R�H��aXa�P���vpi��F �?�Np�Q;I		�E�����z�%�w jբ��D�RĊ:�Bx�H��&�vb�ʈH�B9s"_"�J�H������g0�d���8�ô>��0�:Kd�ga��X�,N���v{���(�~�k���d<"���9���>F���DX��e�Ra��rb��=���ü�_Q])<���'��p��I�	h�����/�,��G�0�Y9�8��bx�%��s��C�Fb̳����v��q�7ݘ�Gtr8{�G��S�Ӑ�s�I��C������nL�"D}s>f�p�D�k�Ԩ��G��%���C�L"7X�<s����DXJ8��5G�X�G��1�E�(�@�L�#ژDX�*.c���L�#�0�1	��1d��E��x�a�L"K	�&$Ntj"��@�L�"_�N,ĉ�f:@�>DX�:$ؖOF!,�f>F�(zD">"��"@��ι1"{��?dU�$b�T�#˘D�� ~�D��"P�xf0D�ǎ��F&b<O*a�L"t`Ɋ8s�B$����α&\x���� �'I��H��D�D?D"@�(X�<3a�����1am�|8A僳%��)��	뎱�JaV�x����{��º@�'x �>���$BX��<k���a�p\Ze@�L�ណ�ߦ�|"���I����"7�xFna�F�/��*�������1�����(02Z�-��H��[c^m`d�������cL�čra������#�\G�Dxf��X����f<r�<w�y%.<a�tuQ����C���k)�3^�w��}|c�'!u��R����ϼs��94KR��_cg�3���|���,��=��@b�>��Zί����gؓc��E	،;�LD��yS	C��u�wS������S�T	��A��@�X�P�&v�=�Lq�	��a��,,x�G��Q<���N��M%��'�^��˾��/S;�7J��ZZ^<�S.���e�
R�Q+%�9�U��x�R�&�@����+>��^gt�wK�aUg��}��{��u�β5��(|���ߘ�}����ǡ��3��k>��_۬�M�3X�3�̺=����9����� 2����U��J�����3Y"��+)�.��������/ ]@T��r�}��XϺ}�}��[
2j�o���b8���~ʈ�D�K�?a�	^8w��1�o����,�I�1"Q�<�YY��0r����ɣ�ȏ1ab/fp�rH`��0f-�J"'����'�B@��J%�P��%0y�??[G��<�B%�Dt��D}��>�	C�D��BI��L�Gމ���"s��D}��O��1=�bQ<�%{��!����16p��L�(���C�"tN"7	"g�X3��J'��G&0O�p~r%��(N����p�H=�I�Oǉ1��ˉ��bh���I�<5D���`3�5��9	�+�"$\"v�Bt}�K$��aD�0����1a2�e5����85!��"�$��τ�bd~��	3+Qnm�X購vSrt���Ra8I��˶'�AEy��Q���K���B6��+��T6y��xu��������3���B5P�ˉE�1����#�Ta�v1##�EDaG��G�=�Ec�S���Ʈe86D%�L�`�DY� ~���{c�D#1eD#��rٙ�3%��BH�Ft{��/�+/1Y6ٖ�+�̤�㪗�..�r��G�ߑ�a�a�|n��a�=Q��n7_����ϱ������չ��u����m�}C�]��/��S���Wj��!������V��߾og���� ai�ý>����2�_3�;���Ƭ_|m
j`#9�>�_i�߱��|߾5w~ohlm��>c�T_a������9�rxmN�c;s>��8���}�\�9��&�¹$gb$�BR�JG���0���!.����12؋(��	OH���{�{��.� pɲ(�'�<&	)t��f$X���s�0N8F`�^@�H.Q(����~R��p��J���8P`��ϲ�����OH�����0������A�k�T������#�����c����;'��uK�yO�o.�,�:wn��;'r�������N�;0��N�ڙ�`M�����>�����L;k�4yG����P�Y;y�b�;�ݦ��~���S�^?-9�H7�9;}����'>̔��o�[ߋ�n��ȝ�_];��`���hM�t.��}~#������#����_�d���ux�7 ����O��a�A�/��v�;�ov��T�^L��}��y|l�~��`}�3s;'M����nMU���n���ҙ�h�=�=��������F3C�����+�֏'o٪�7�w�m�OO�D׋;:q������Ň��-�����s�H��l�~��0������s^f?���������5|⿞c_�dהUF/�M��������A}߫���%�nS��'�}�R��Q��C*�<7�iv;��M�U�a:un
��gd�G�}����={y;�5��RY��Їs.r.�[�Z�������h;��ɏ/g�oӤvyCs�}�/S���χ��3*�l�a��m��f{]�b�v�k}�}ݟ{ކ_�����״v���̃�.�O�l����?����_����1}9�>���_��@=�`���d��;��� ���8cOZ<v]�aM~���z�t�W�s3�o��9��r�&�.����~|����w���uv�0�{������t��;M3lҴ�FF��0�86���\����g�z�f���ǻd�2�j˟.�Y:ø0�W�Zj+�2�}�x߱Я�V���Y����~��b�`\��n�Yߨ-]{�dNF�r-�|N���{O=)��fs���n��m�MƲ�>�:sI�[&��30�e���:$�0�Ј����~z���D�P �@>�?{ǀٛ�n:wi��fwe)뾝�dk�T��Jfߧ*ou`�s�q[��o{{h���F5B�)���^�^vV9얘�6Ք�M�9���Go�6��Z��w+	�㳅����Q����ǰ{��kYܲ6&n��~�<.�ʈ����s�����4�Mk��:=�ǉ��X�}(.��s�̸����y3�0L�c8�9}�w���v��e�#��&�c*�Pa�ßt�Ebג�{`"H�[��U��՝�.vi��ǻ_e&}�.���o��x���Ƚ�#�z������Z�}/�*��Oo�KG'U����>ض��TX��ݽlix䟋�Y�m�g��~<Ao��b����>�sS덩�3�7��"��a�ʜ�{ɭ�gw?f��=��c��}�̦N���+���ZwO��{���s��� �b�uw�������Nr��,wv�f�)�nC�ܙ�f?v��M�^��]�g�=V�br�2�p�c|�2s���ݼ�]/{����� xs�gOz�}�ۉ��OH����N���v^��p��u�n�}�m��o�?�$�}]ƻ�g�۽z�;!�V��^�����3{Ng�*�\9>���o9�GW"ႈr���$�^�TDT����ϯ=��~�c9�-�(��/9�q��ឣ>����Tϻ���I��zo�g��w���Q9�u�����cO{���l���:�)�7ݾ��c��{������u�p�da�u��{fC�{�c�청��(��r����珼=��$�3:�c5k����i���!<fg2h���)��G{ғ��c�O��������������Ww�Y�������Py�L���0؜���},�d������X����͙��703�w�@��/Ok�y�|�?{�/��g�6�U�zL��R$$s����ڱ�y������<�Q���{�۞��.T��B�lO�3�E~�J^�Bk�$�U�s>�s䝀�n�!��7�����d�Zs����$�OcY��!��{wC؇w�$+��c��]��q�[-�0w�7wy�z��{�=߲�d��<h�?�Ӫ�~n�$�m����9r������O>�oW�ݞ�;��0�.���.Ѵ����{s�t�SV��r0����̕�;�t�~�*�G{�N�{����v|�vw�>V���]��c���{�t2CO�&��&�ˁ����ӴxV�b��wsy�VkS����&��e�-�l���gz��������.7�M���ׁ�����vcs�k+��;�#�nvl���*��.��Q�K>L�.�����Y�]��w?I���쓓�S�T�}tf��T�����c���\¼����^od3'�;^��,��>�b��v�N>w���}3sX�)���r��ڏk��.>�������Z���vf��H
�ǍYu�x������N��Y$��Cf9 tf}d<�Ж�LV�t����`���[w�"�5j��O�M��10�s�����v\��6>�ߞ����ۓ�F[���5��2:����!����a��_��{��)��}�$Vo������]-_H�����]���;!֞>�h^���ѽ�[v�a0�Y�k�Ɲ�2b����噰#rf�Х_K�I����bMr�7���`L/�;�";u|��=ӛ�o=o2%�50[���{��VGo�N3��&�k��C��a�ө�zl]���^����b�<�=���;��Q9#�R����=;�9�Ȭ�gw/s���~���ՋUwVZ`�}�������^g{z��}�wg��&������g�z�$��K:�O�ɯL�*���^��˥��z�$����&Yf��.���5�OK�3���ݎ{�״���̆�ۻ�K�d��{�I����a�ϳɻ�|u^oڟnn����3;�:<:O��ݒT��>�~�;��1��$���h�n:#&�©�'�<��|/�{�^�)�������wt����7���	�ɛ���R�W�_���K[<�����%T>��B�����==^�ߏ'@����2�����	���$��bx���b�|����Q�X�j5�1�ny���!�J�"�R�Q Qȩp�*����"��vd���q�Q�2U9S���Ej-�C��-Q�Q���W�Ȣu���n\�n�X�4U��YJ��e��E#�j�S.#���Ō��j�[dlE�r�J�?�El�>�1w)`0n6Ue+�#�ڰN�1�mi�u4iY/2Ե�ۘ�.�TU����!�\Xک��Ӯ�d��
�r���v�.T&A�u��Ö1�l���d���
��KWNL�&Q��hR��FP}0��4g��	�q�]Z��Wް�yT%י�H)�f,ʛQ����q��ł�$��³Q+��R4أ�8&؋U)Zl�:l�T�ckꃖ'"Z�:�L+%�"85�gU[�w���U�FT�V���-�F�A?�9[mbnȨ�U8�h�	*�r
+�@�㙕��X��&�pV�E$�%������abm�`�K,i/!ܢ"p�'����)DU�X�kB�� �&�j���0�*��!G$t#����Q1�UѶr�&ډ�����2�Z��9Jڒ�0���6E
R�r�h�(7_�T>7[�"�%�ʉ���ʱ��H����Z9��U��R���ELU�Rd�I�z�oB6����7����d�FB�y��ǽ[f�b����{�3��Î ���|}wڱǈ�f�d��@�c�-�����j�&����������َ�ݢ��(��'[l��9���'.4��nA<w�Mj��U��'h�i�Zm;<���hN�W��]��ӣ1�Ty�9}M����c��h9I�;%+�2v�L���	g(��Q,|�1�Y�U��e/%,��U�!���b�x�U���i��e�8&DXEz�f͡eƈ�Ƀ�q�Ir�a�{f�>�5^I��T���\��\�u$��*qZ&(�;���'�IdU��STQZ�qGm���P(�6L�w�}�F�c�t�bho'D��xˣ'��b$�IQ���l�� g��ֹ͙	� ��d=��-]k ������-�-"��?���nIR�!�a1�>G�?���쌈?$d�"#�#����/�?��o��UUEUUEUUEUWUU��UWUUTUUq�UWUUq�U��үUx��VUU��{�qQUUQUUVUqYUV�UqaUWUqa��"H�(���!����"����"�(�
�$�@ؒ�I�Ǚ��7�����򲪭�*�Ŭ*������������
�����������0��k*��G��UZU��������ʪ���U�W��*�U|��U�V��9�s�(IR��� �H�"�"!QGQ��R�F�(]�"�M�&ě�2sٙ����fc�W��*�UiU�Jʪ���x�j�U_*�U|��U�W�ʪ�������0������U=Uz�ҪүUUmeUV�UU�UU��\̜��cHc m lCchc�|i}��������ʪ�����ʪ�W��J�UZUꪾW��J�q�_+�U|�^�����k
�������{��2��k*��0���������������|Q
�d ���2H���H) ����h�	PV���ݒbAbV� �?!�>>��@`BDa'��ϯ����܁�������z�2{L���Q�2h��g�6pИ""ag��D��"""Ad�$���HD�(N�tN��$�""%�&	�DDD�0L0�(�(Nb���$����0�8A�Ab!:& �ŉD8'0�� DDO��Q"�""P�b&�%�%$�8 � �Y'���pL<b����~�c�_[�G8F�'�e�)\�;x�u�b�mQ�M�n�$��Pe�e[n$��ȥi�Z�V�'eJ0����<�	��b�@R�8�c�?��ry�Z691�\i�)����ܴR��Qi~��<�����^%U��0����i1F�	�9e���B9n$���ձ�Fq��´�h��O��<��W"$��NV�A� 2E��]��m�6�
d�`%�G���$$D�RB��n~��O��g$�<�)0�b�>�1�ƈWe�%b����\{��(�k)+V@+��lV+`�$ ���i��4b]��p���r�\Ņ���[UR4�11QWk�-�a�'����Ò���Ą��`��b��[�Z���I��ʔi�*�NJ�I6-�88���+!�cP��Q����,���e�Q*����BƉy-�;Z�
;-�VƜx��}��Q�\�W2�uV���SC�>������QUj���ߏ��>#wwwwTUZ���w��7wwwuEU���W~�������Q�i�`�&Ag�����[�霊�7[t���[�1B8댨lW��\n;*j9"��V�0���J&�\2#bz��3�"Ь-Q��+�m�9SR%���V�K�q\""ڍ��F���D:'���T����m���'��5�2��BJ���$.ۉ�x��GoRK�:N���'PG&�E&4��m�թI�Z�h��y8䍶�"a$c��5j�3��� �B�GV�K��Vxhg|�l�u|A�Yf|Y��Q��yy�TZ�j�b��y����:`�vG+���T8��	a�F�wYF�}j�L9,���MЛ��sl�����j���=R���O���n���o �2&�*o���3�	~∥e���Ax4�ͲDr8��b��Ԇ^��l����_ВC+ǖD�xӧ�,�	�`�&Ag��פ�!M�k�
��=��;eW|*�q#ѯR8t)�0cL,�[8O�)�N��,���a�ެ[��H)wr˻���$L��v��g��rA	@�r�q'�R��,��CG�@�|��Ÿ��vtdٽ�FN1&k'��0�㦘iFY��Q���2�8J��B����m��������#�u��w�5{�E��&bъG�N�Q��l#���Q yt7��"�t�t������Q�H�7�
!��N#�N�4G��Q)�-��B�q�@E<mI�t�o�R�'�p�|Y&p҉4��0L���,����;wS=����/3���fQ
�m<�v�j���&5�mxa	\<�^<��a�#{�eӓL��Y�1a��0E19�Kj,V�T����K
���㢜�4�Ա,��LV�r@�vKU!h��ڢ����U���g�����Ņ<���erICDq��8/e&^�Vm1Z����7oF�5��D��5��])��Q��drT��Dq]⋱}O�k���HKa�x#�H��E�DI�s��L�������A�c�J���I:Q$�Y��Y�XYc(�����p�l!�@ɦ�mJѨ��c}<Ԫ��iq�'8�M� ��W��]���o�V�O����
>I��כ���z+x�	bD{	�3.dķ)l�t������AJք�x�\���.t�t�u63O1��E&{��b�!!t�	$�,��,,,�V��Z8����'S�+���,��
%�cA������<}�1컗,�ugL,�e�Ч�*�ߓ["�lU�H�;HL�Y����fC��X��s@xY��f�t��d#����£�QD�A
t�G�Y����o�O-]2��ۤ�4�I4��,��(���D�$�T�$�UN��� �6�0�� |�z8&Jh�j{�W��qTՊY������T�sx�E�U#�K�X�F��~,��"�_%��DlX���N0�C1���D�q[:��Q�kp��CX��IgL(�,��(���D�$ˏq@��/7��f<V� T}n��D7��# ��5Sp�Ʌq�u�9�)�x㉘�qy2��7	w0��u�"�M�B:�9jHӊ:+�[֪#k0^ ;E��UR*�J����:V�h�F�He%wG�2��\-`��u]h��yu�6; �����`�}@US��ϧ�v7}v0��^+�Ml��׶�ia�nxGr�="��6l��=w{��/�m��B���jv6��7�qK@Q5<��;�6+Z=K&�><,��,L0��<T�%�ƾ{��L�C��*p��z< mb8�H8U��]�Ȏrpf#C��w�*m̐��;���-�#҆�x��I�%R<b8<ޗO���c�:�7bBl8�~Ng��6d�#�����K&�M�)2�9Ѩ���>D8a�	�!c��1������x=0�G��I��R0�4��F��i�t�t运�x'����xR�0�����z=�$h�kL#Fh�,���|^c���Дx�}ŸI�4zY9�F�D�z=4�>'������|OO1��GrxtOc��)���_-���?V���?
����>O��� њ9�$�֔A�VYFH�h�y�	I>���������t�~!�|xv,����x���xvx|K6ј=�A��ri3��oFͬO�6}��C�>�Q�bv&�I<C��0kx���xO����Č/�O����7��L@�~���C������}wpXnz�c�y�����o����ٛ��﻾����/���nuTׇ���3gǶ���fz���=/h`���22�j�_~�����s�>�ם����7�8w�Y���!ǳ&�~�^���4���[������{ު���;��{�����w�ꮟ;��������w���x��,�4�0K���L8a��zD��Ui����p@7@�s��L˫���˒��E�1t���؁А�C�̝2�!��aNq���HuĲ��!ww\a)(�kL�F"	�y�D���~S{�h��Dâf��p�jd8H�Ob�9P��
0��$�6Cy�W��}���GR���FI�ϖ�`�`|��hC"�᫢Z�5��$@�!ĉ����Hl��ۍsG|!���O`�&�Q��8i�ύ>0ҋ(�K44���K8a�jBI�jmUU�D
H���HD6@�#�	����>���Ԣ�F��G#�nK�!,�*�帹���qo/qK�v�{�� r	�b��u%	G~�(:}�|7r���4j�?ధI�R��J8 ��tf �0!â��N$
!ĔC�9K��ȏlZHb�F����	�$KPt�]bJ�ov�J%(��O�^� ��gBC�jpMA$�ֆ�6nz��1�������?��0?�a�Ζp��&�Ƚ91�ǔk��= ���֛���V3\��ˎ�.�5�MrM�[�Ud����#�g29��b��ν�bo��`9)�q�Tv�Gah��`T���Gc!'~Ң��f���ə.�`�uM�&ݱ���6n���O"pN�P�|���:�c ø��QJ�P�6���6LpM	���98hq%(�c#�*��0z,R��P��K����!���U��'��l��`q!����b��@< D�{�L�I�
(�=,�e���C�C��d�t`}�d��42"�$�� �4!�_��}ւ�qG�	U��J�.^��9�@�&�B�Q�X�<0�Z���H�\��zl�:�4&��$ٳ��4�h���00�$Å�,�5ۻe7g�9��*���}(> a�r!ج2��%�$�`}�wF�:"X�������rB�;BL�u��&����s-s3D�2L�2J0�@���T�X6����s,���wh�5A���/��V%��*�D��<�@��'\F��0#6Y&�������fa���4�8P�&� ��z�*
��9Μ^HVm������%�0�-<�d�����#���e���h����A�؊��#șHi�!
�`u�,��D�ǮN�� �R�q�Q||ad�a�faFY�Që2ƎG9CM�k#޿��UU��W�U]q�% cJs�\�؇�C�
I;��)�.A:{izM	F�8r4�H��&#��L�5�Z��+rÀy�5"hI�*��b�E�І���7�iX�j��79&.L��X���$^0�0"E=hB�b_��5&�')��4è��(��R��aI�a�
"��*J���!4ꆬ�p��A2�](P�jMu�P�$&f���C��0�S�#,ᓡ-Rv��!�r���'�g4aae�YGN��(�6���둌82�1�H$)�fs8����Ҵ��t������h��!�%�h��z��hR���H��7�nX5��!N�c[��E^�����'�+�H^bD���H���D��d���b{2;V4�0�<�Κ�	�NI�F|R�`0@j`��nɉ���j�j	D&�t!�!�0,�A��t0NJdI���lA4Ġ�!�!�"�7 X��5�<��4��W	_a�I�~0DK4�:t��&=0C!�"tdB"h�Pjѫ,R(�Zr�84�p��� Õ�c9��4��G��(�ҊXd|�&�*d�+!`�YiQ[� и�Զe�9�UUQַ�$��b�Q��]�P8��l�)�E�[��D6�i�a��4��<�XӸ0>���)�p.�]+L�Q�.�d[�(&�ܠL�	��b�(�ç��Dl�a�D���0Craz0������8a�J���:2R�"� 9![�B�N�$e uD;:�N�}|���j�֩�'Iqvؠ��6 F
�-,���o�=x����י�l�z��7��9T�Y	��ipv5
<�����<���� ���È�X�W[�䚥��|i��i��,L0�L,��I{̜���tl�r�˚։��UUT@�߾6�D;�$�^����Pe��{��I.e�b�-A��%�vEȇ����CQ���6�q-������X�kRt$-��0��a��#}%����Hf��{F��S�I�2hC�M��FA5�%<��h���u�� �Bd�(�mbQ^Z�.$d�ڋZ��c!���H&��s*��C'%��5�2���Z�ba����.������u�A��bSz�}��e�Z�KS�0!�����p�L;:,�Oa��,L0�L,���!"n*��!Z Q���*��n��R�r$�
0�$O����'BI����>�'�y~ϱJed؉��O� ��Q����:S�S�v!|ߛ浳o4�nl�/��jQh��^�>%9��(1:�I�R�a&�<�zp�W)�nA�v{�r!Ї�v��V�����4Eq�	$j���hH��G�,%�f��G
nA�@�wlV���3(p���<i���ŉ��"%���iӆ��Z��eW�9y���,�"��Ϊ����ՃD���č�i\0��p[.�	�� ���%��t{4|�0a��~���W���N�n�6ˣS�d�4!=5�`�)C�d�oj(�wC!�Ԣ2DFDa��76y��J��j%;���`}�����1�i�8(��fR����|CZi: "\�v���'a"��a�J;�5��)b'c��etFQ��y�l'd�!�e8N��G�p�i�ag��H<<�#G�����:iz=�4�I��<O��8)<D��<B��k�8���(���HX94�����M���t?��^
p�p���?�"ψ�`�� zM#Fp�4zIi<�G�/[�&����х�u�����eS�3�b<~)�8b(�
'������z65f�Cѫ<Bђ@�&�0�>��='�g�Ǚ����|M�Ʈ"x����,������i�<��4�	4���z6=O��>���S�G�DؘA'�^&�XxO�O��x�!��%�#�br''E���72�X�I�<{ni����K>�q���d�ϕ�]����o�Z�ٗ�*x�󊏹dy6,Qߞ�f.�A���٘�䅱�q�O���k��OL�a���R�e[l��MzaA�:ԫ2�%/��H&����bv6e �����K��ߺ�	��D#Uk�_E�\
���L��r� � �||��S�y@�+lJ9���ɒ�{��I4�G��Kd5jr��ս.b�dʜ������w��b��[�Y�9Z�,������7T2��Uܸ!9��׸\���"�$W-��r�,܁wtY0��V��A�QL����9/����T|�6�k�1a$�|U�"؝~������L��
<��ǘ���|sN���u�_*=�Gߏ����s�ਬӧ�&?��������ѯ{375���TK=/W�o䘤��Mv��
I%jKI�Pꃑ�*��R��� ��u�b���("���:��DTcx
GN>�a\�A��$���X�j�i\�c�Ҥ����"��H�8��o*�FT!���ME��ӯ���TR���9X��*��dn!<Dq�T"M���EF�`�;B�pD��ᑹ=��3*R����#��,X�Y[�>ϒ���Z���w�������wwM�n���.������B7gwwwmYW}����UU�e]���wp
 �ǋ,��4�D�00�4����}�'�#��9�k�ɐ�D���i���j|l��1ҷJ�x:�$m�嬊��3qI�u�U��$F��@�B;��\
�QX227c�|��m�%���Z`�Tt���8��Ub�It���d.�')6�0�tYX0[$��yF��A0���]�K'/H`�vS�+�p:�S�e�����=�d��ϸ�����d�2øm"���a����G<��{�T�cd
@#�+C���w=B�a��3MyM�L7YGtQ����~��̬�A�눁��G�o����J ������iéV��Qg�P��JvI�
?�?h�b`a�igNu_�����⪪�;R�����Xh�8m�CQqZ��Ϭ�M^����n%%(�i/"&��GQ��a���8AgQ��8i�����jp�I�ah��+��@D��̥&0Г�Z���Qd�/F�0�.�sQƪ浰ԸZٓ��q�r2}:,��M�qI����^�iR�q1���9N7�!�`xC��8=�D���MD(�5�l�Y�Y/~`'�O�~L4D�00�4��R\�t$��FK���⪪�����q��id� ���	2�� C���%��K-���'�YD�5��ٸR(H�����yQd�N���"t�ۤq�M�)s��Y���}:���8����$1����Q���l=_��S9�pIV���W�p��H0O���jg��������[eo{���̓�]	��hd4=X�'�P�F�	�ʆek	r��Pv� 9��������?xO��Ɩ&��4D�00�4�y�U<ݤZ7�ʪ�������!�]��,k�znC��gs
���P;���'�O��̚����+$cNIw�_*�<�����a:K4�����F-$6]N$MJH�v[��l��B�
v��.����h��$ �@hH�ïj��z��0Ϲ���U����]̗Ű�a�ξ�ҵ��Ä����gKIE8K��.I�����2h�>=½Z�3NL%&�6�)��4�r�w�&��'���h�b`a�<pú5}�Cˌ�/Kx]av�\��AUt������qڈGk���7��yH�M�>T�B
�D9$-���c���1c�Ɏ�����O�ҷi9	r:�V���UQU_�j�����UU a���A�%BcVIX��vF��ɢ���(]�\�Qx�Ś2��ƧuU¦�	�d����8�N����Uӫ�C/ؼ��jm���cG����gE����~�{����"�oF�'t��Yu���xpق�͝�[��#y�ivJ�B��Up��U�4|8r�4qQT�%Km�(�{��җ��MFh�jx��18l�A�yM^9Sbâ�
�k���~���?%��&�%���Y��������a��3�UURwM+!��Ci�Eَ�U&}�ª�4��M���gF�vD25u���ƫ��cp���3�(�q,�[���F��t:qUR���`����U�&S�X�;�|p���8rE�X�3,�S��@d��k�6أ�tBdf�V��Z�AEy����e|���*Q���㬣�ϏaE�|a��Q����6Y��g̈́��mUUH��p�^wyQ��y�����!.��`/.�(������4�Ad�l�Jd����G����qD��0:o��e�����e����$m�s�#��sD�5WMu��ӡд�j��o,��DEZ�J,>�a�U�H`� ��Be.��7&%e2\,��Y(�Ԑ��<-u{�Q$�>+����(����M>0�M(���D�4fߴ���&&&f�3&3iSA5)-٭nm�UU �s�ѹvr�W|$���Q��J|�	�4�n���M�*���2��D����l�&+���C�a��dJ�c��1̕3���:p�'J'����BҠ�4�N7Fb$��o�5o���dN��a:>0����"T(�N�F���������Yg�3�p��|I�G���x���C�Hp�g���i��^Ifd�E0
}Z�G���XK�s!f6��:s�*w-d`�U[Rɗ)rI����,*b�W�����f>�iDP�18>YF�| ��ڥ#AU%�jX�Tay(1HS���X��߶���w��i���^�F�����U�<?G��m,X��bl�$�Q�"�U=����M��k���`c7��gF����CP=5�����Ɂ4��\%Ӗ(����&�p�q�.��`�R�?#���Ջ�����c�n�#vBT䐁�n@���b]�7濫R"
��4O��,�4M4��::C��<_�6�0�3�$2�Efe�HH뗵UU ~=�u���IՈ�!�N���;�f�Y'�G
���ae�4ehh�F��nO�W��,>PJ��"�sx��>�Z���P:�$Sk�|nW(�2T�V�R�#�ܐ�A}�8�[�R�QN���C�o8mS'Rh�750�#�Ys�G�()�9�|�3wz2�C��4�|<�-0 �'HH4��R"M$M'HM�:M!�Fi�p�4zI=�L �z=Fi�<i9�њa=m�cl��֎[�<A���CD�O̏���<g�/����>/���Æ|<������zDKzA��$u�$���3�;0|L!�ƺ[ �D�<I'DL/?
3�D�S�|'�<��Lz9�F2�4jG��	��h����}/c�~���{_-0|Hx|y����l���>g��z=0�i�Ri3���7��4�
'��
{W���0L��4}Ӥ.�A�<=�����m����6g�M6����4ޢ&8y�C���?��^�on_��'�n���I��l���s�����o{��,ɞ�G��ޮ�ų3ѷ�����}���۱�̝a��dG���ǷY�sQ蘉�����G�M�r�����*��UV����U�o��wwu��YV��U����U|�ŭ���w��x�e�x�M<|x�㇎�N��ǒ��5��Um��I�͟��Gr���u�V�����,�d�F?}#��t>��$��������w��qLs%)Tն�%��r��-nۭ��y����/��ެ��7O"��JK�M��:h�[=��֒�g:0��)M�46�78''sɳ�m�"%q����g���:t�>>$�O��4�J4���Q'9�������3��|�K93ʪ�@i>�N�Z�����C�钭0��^����Q&��'2d���S\�H�",!A_h�L��Y�x*P�AԊTߋZ�ϽV=���u:�9���Su��2�8�WN�B�Ӳ��N��\q2vlCZ�ND��J�^:��o�0f,R��Q)u�������a�'��Y��i��iae��N��<2N��/���¦�m��sr���Y\̐�<t�)�0�?��[oxH5�zJ,nB*HO��Y^f�cp��L�2����$P�|���.W������Z��D�R����I-�J��t*c"���ʂ`�__�UU l�M����!�0���Nw���#�nL��GS<z���I��[�~E��M�(=�����g�!q|�cm��,:2��mÈ�>p��\#e��Ę�0�j�G�XttjB��	`�O<_��4t��!���cі���Vҿ`p�@����g!�������c�k��4��Z�33+fQ�ĩ*c��[��{���s������w���^��ڋ�(�bζ����E�QGŔa��a��Y�2�8O�o��9�.������,��!�?p��=47f�{12vn:(�Өvr���]H�m��k�CJ'�F.��9J&������Ǥ*�hQ}��W��C�ɒs�z�������&e�9-b�#x�2��e}F��(�xM���d�b�ò��C�"�T�}%R���k�q��8�>/��g��E����$�K>4�>,�M4�L0e�pжV�)��c�$k�.\	B�2������gk��̸"C�c�x�f6�j�+��O�\=u̶� ��Ѵ�~4~,g8p1f����DW:t���2 I*Ԓ���sB�d�c	�����q��`&u,1�1��8"et��	�F���V�Ҹ+�z�ڔ�X(�.˞<)�>�r�����!�s�èQ ��_(�I���Ř&�i��a���ч�1r�;T1>d�E�1���UU C���$��>?r�Q������� Ô�a��)�/XW5V���f����f��S��Jw8d,<�QώmCH{�/Ga��h�g�fGQ��@a����p$��c�����X�bg��a��Ç ј8�6>��1���@����ȵ	���QRI��ƘiF�|a��if�`�$ᬁ��DS��j	Ĭ�:�mN2`�p�^U[�tÙ���1Mtcn!�>��U��"Yܘ�d	YM��BX�v),�
���ڞA�NBV���]�<���&�V��R�ح-�R�ҾE<T�����4Xu-!u5x��
v�G��ˎqaA�
�a�\<�P:L�â�,kNW�k:eg17gD��=�CA��:ѣ5L,��6hC�O�|��7��i_����J�D%�Vݎ�;��^2e�w�J��������ւ�@|��������I��(��4�M,�d�0�1���j�ۄ�>UURyFY���,$�P��p�Dm�i�4�JE��"Ϥ��_o���y�WH�|Y(h�h���te$H�L�_[m�8E�R��!j��X��^��W�~�Q��#��I�2�P\[�jkظ[�d�t��6�nB��;j�,`��o�F5�|�駃
E|ܞ���uq���~>0�N�aE�a��x������M�R@�"e�#Q�|UUi!�.���*�[�^�����\�U|J!����j:���e�����:2&Ĵgg�0��92Fz}UEim*ffQ2��Sbjt`"u�s6n�-��qn3&��~���4a��ٰD׃��^<���T�I<3��.q��Q���.Ci�Õӄ��C��ɳ'�Gg��a��ie��2�8i<�{�y�$B�U �e�Ld�'�y^]ڪp���lDq�3��K�(�F�q���k�M�8��-a#���&�pEBT�@�$������c��Գ����jy�}��a���=��3��f�)����
`���*a５����l�eSvQmx��0�|>l7mP>!�;���0OHb��̆ĔH.G4��(���>��g�a��F�:BA�&��i	��F�a�0����ti>h���$h��4v9��F��4z>�G����4kL#�јi2M!h�oH:i��h�O ���/����x�<=<>!�<hSG�����<;<;<:=m��f�F�A-�4��xK<=4>& ͱ!�!<BI�D~4Z'�JY�|���x:�=��8R�'৅83��؛>��م�S��<3���8?��tp��x��<>4>'��p��<<4�M���(�oH����f�>�+>O�>~�����p�ˢ���k��l~�τ�^��O��ڴZm�n�*�k�`Q{���w���3���!���a���jdM2�D6�����U�D��K_���_q��{1O��ɢ,�E;�~�����7����r.��>�{�5'�L��r,�t��;6d^�9��Co�;p�)]D�B��1�Y�b�
�ݬ�3*�D�fO��w�����(��F�7�}��zbMꭽ��I�V��v�#�7����e�hl�6`��:����$D�`����&�o��d)wf���5�yo����]ɱ�n+��)�]�lK��D�ۿ<�g�g��1����[W���(�^�����~�0��%η�G�����n���7�U۪�q^��}^ы��[�z6a�IDצ3�����t�E�ń�̽��N��v�f8.Ʒr=[����{��3�-�)��̾;�Y�gq���x�s2x�gy_N�������u�Ic��E�U`�k�F�����Rdj2��v�c�>Yy%�BڤF�	S��v+ϞD�S�NfC�6�rFY%Q�5AK#�UF� �6�C(�Q�̫%b��݁%R7d���RG�K%@
��]�02)S#�"��V���ܔ#8 ��q8W_�E�f]X��PhN"�V��R���Z��ڿ�ʼZ��Un��UZU��o��wwu�J�Z��V���UiU�U��n勉ǎ�Ye�i�i�i�B���_��Wd�/m`�Дib"����r[#@�W�Ufeo#8�Q�9d��i���	8Ӣh���,�-r1�)a�UP�1��&�-p����N*�@7-�LH���m��зu7��T:ء�Ls<n��?���C+��xa(��N3��t����t�\v�[j�T}ppd-D)5x���C�S�ٓ�VAN8`�z��e��>4������:tgq��TJ5E�>��u�Vb�Ė��d�<��U
�2�d��!��9inDC ��$�Z$<2���r8��(�B:t�M0�
0�L4�O���!�e�>5>�l��UUi�,�T����Iх�-��q)�"���<X�"�E�4=��>��35s5��ON�O�uo���9w��K�ƷG��N�����S��fÕ�,������S��q����AJ��G>⫚��$���gFP)(:�Ty|��|��:0CÓ�w,)�7�S'ZT�:|�0�,��L4�M4���!�e�h�P�(����Ul�X'�Қ<��0D�0�ϼSA�4�J����ե����sPá�3��(d��N���@ϡ�a�S�����{�^;��]Sj�S���k<�wN3*�cl}i�I��iE� g�f�gB��P�:�,�3BCF�e5E��rSӵ׊��(��>�0��ň����aF�|Q���i�XY�6Y�zPMG֖[p�Y�UVQ3��<9�::����rjy�N�䜛�6ytS�0M{�ESí�#cRRB����緞^☗����0NH{�gsf΍����by�)�r]{�7Xl��=�ˣ{!}�,�P�P{����>�ȱ�2>�|XmD*�}DF{
��p������X�@&2��~?&�h�`a�x��4���H�v)tB�'�#�Aٽ5��фS3N��]8�	�d���n跙"�A2;��h�u�3�gGX[ʇ"�LuX�U�!4p���9��n*��x��,����m�[�9����ۍ������� �V���������F��~%�vu&��C*�,�K<{��Jp�B�x��G�}���r�.})��M�=	��x������]�0�Ǽ!o6[aD�	��U�9��n }A:�s��5�E=>߫���]Q�a��d��iUL��M���L��<)J'ZA��J((�D	���M�pደ�Y��O���>>0�M0���D�Y,�:q�P�x�J��$%�����s4BR'N�-j�&�ݏGџB��E�O�E��fD�:0��nP��&�V$�lѮ�4'Ӣ�Z��{1D.��أx7�$#�
&�)#���e�<a����-����К4v"'q������[�2ސ�͐��M�l�!���;,��������G�?h�Y�h�i�`a�x���{���iK�������C9W��ó`���A)�;qԚ=�j<���-G��-}���w'�ð�G)�l�8-��%��r�fLűT�)u��%֮�L����9F�	�����L ���~��V0�4�;%(�#�\5�7O|j*t���_��$!�9^�EY�Ό�qQu<�y��=@�z�K,D�4�0� ��	�M�x����B�⪫I�?}R�HU#�>EYëR�Ã;�x ~q�J?����F�r"�-��#E�it����C(���Q���8$!TJ=\;FB��vùx^d6z&	�$��ML�j�ڷ��S��LD#�����C(e����(uĉ<�Ppg!��A�a�Ęi��|p����6Y���i'l����l�!&?�C0��z�I����v�x\�-�tʰ!�&ř͒D>�t��F1v�,�k�TA:�S�v�**n<N��mX�ԇ$Qƕ��n���UV��on2^a�.D!�TVH;yF�IS�7$P7��_<m�Af�V`}6ie��d/�M�).S���莐�Q�H�R\�(������т'Z8d8u92�x�^x:3(�>��!��>�QNB�P�63G��=�D%����g��[�H6�I�
�u�b������S�E���>�p�u?�QI�r3	,��M0��<|p�Ӥ:'�:��� dg�az�!�U��5����i�s�i˗���m�N�,��e4Q=��:<&u:52	�jGS|�󙙘a�B&�l��X�I�;3$.��)�|���ŋ��k�òA�!��|B���,����$c"(��h�D�Q���|�Ѧ�ޡ�&�X���b�r�UhSnVԖ��ra��a�a��0L�	�`�f�&x����<��g D����DX�(D��t�� D�:""X�g K(����<�P���"H�`�,�t�@�"H�tD�&X� �t��K4馚i��Y�AD舞0�
<P�t�AC�$%�N��:"P��M�������[�V{r��v�}�����)�O������������~1����߻���ٸ�ˮ��d�N�xLg�_�ϯ��+ѩΰ�b�Sq�x������5�#����'�t���[���Ɯ%��O} ��On-Ɋ-'`n�L)�׿W�U��T���_���fn̷��vr�����t�������ﺘ����gr�iU�U[�����iW��Z��V�����n��U�U[�����iW��Z��V����(�Ǎ0�D�D�N��6Y�'RHk���$'�|?�]5C|�ȯ�Cf��f��Q���=��ߖ�[Lѱ53�����%�2��|aӤ!����Z���9Tt) J+(�䲨�ء H��<t�fS5P.d�i��\�����H�'i���R�ј�U��m7nNJs�ML3���!gGC(� co�I$��I(�O�4��gN�!�8l��Ԫ�ڽL����fk����UUi!���ô,8�4��$�
��l��2������R��B�E�x����>>�I��6#��Ƽ�J�v'3�K$a�=�O�W�/�H0��Ԯw���3� ��͘J?	uEg��"��<3@d��>,T�\G���� �p)��HH�i��](��E�#	K�O�<`�OƉ����aY�����b��Z��<����i�\Q�\������1����h�kV���̍X�-�&:
'(XYl�;+R�ddM��i��HG���x�Ro���$7�f�

)H(����.񯀩L�1�6B�d��酘��`�؊�fvQN��p����;(������ɲ�h�MNaf�K��Y˧)���e�q� \���~��e��Dy�Lc���@�4�� ��{�WNt��pZ;�q�9jFA�EQ��a��Y%�2�8l��ȣ�1�N�����J<��c����V������M�)Fi�ڊ���j[	G���@p���d,�|�!�%2�HA�W׾oz|Q=�6姙��&f������)U,�I�yӄB�sx�R�r����L����gp0D,`Ġe^�k"ԔH��Y��a�?	����0�	,�����%��c��ޗWf�.e�M��UU�K9��g]�ób�R�KI�Gb&�S��F�AO!�f�M�zY��A�u��|�LqT�bfX�r������6�����_Oa�HC��G+t]<���k��+���=��Fr��������C!�7�RJ(�7�>'Č���?����tX�%�ko��(g{`س<|i��4�O�4�$��Ypӌ0i�Gb��Ծ��UV����õҏ�a������q�0�2����MR�{U����0�2LEl���L�fL5U��|z:�I]:�z5� �ќ=�[}C/��x�˵,��
��1�_x��(x:JR���J!��6��P}����r��B�t�0��(�MM
0�$��E�S�y�����(܍r��x�U�����q���[�X���H���V�l6�d��r�-q��j�6��Yܸ�s�T����԰��[��W��BjHGGF'�	�� v�8����m�ƅy�z�)%�NV9@�r'X��T4�c��5j�c���TM�V-�����G���*�A��KmZ,��OXa#(�Bl����>�:@�%�G�[F|a>E����#��d<ln���K0�'~g?Bb7s0���p�`�`�r�C�=�N�΢��.�`����$�ǋ4�D�D0�	,���5�&� s�UUi!�ܢ�!�?Uђ�ι��
�{�4#=n͈4���:21�S~Rs��/��pcG(�t�]|��d����5�Db��`�u2'!ɐMK�ʦe�a���G�g�_�R��B:w5"�+�1�,f�tf��-��J(�Oh�&�&a�Ig�.�d�k[UUi!+���U�~��\^,d���å��d/��ń�H�1A�Fʒ�pe���j<�q��jfYq��in���t�����Օ�1�@a��Ya��ժ�^=}*F�C��֢��76��V{��.�1�k�����a��i��ag�,e�Q'
16xa���Y �S)r0��UV��Z=cknA�PybR2��u�����.��5r!f� X��IL�ɤ�	G2*�KG�ay4|x`�u�1qn7!��%�8��Ã)E�=��GBY�2����qb�!�Ol3���ԝ��L�����r�7>�}�'���Ord}3ㄚQ���4��,K�$D�:"'�� D���,DI
:'�gN	�b!:""X�g DN�"xD�<%	Bt��D�$I�8@��D�<tD�bYRE	GM4��i�M4D�M0ᡦ�i��4D���xDL;�(J8H� � ��H�'N�BP�BI���LL�1ɘ�;>�8y��Y�؟%�d�ȭW�PɊ���ܼ2�/M3q���j����ӛ���M�;!]ɯ>o��7�������N3�>N��j���z.�]��5oqE�$��l�N�[�-�"��1�Lx��Uu�ӥ`����_����A|�Z�mU�B�F��v>�fDZ�i��iy�@�L���Ց�j�j��ʠ��Y���Om>��a��3m�VwV�"����m��$p�tZ�ROj�w׽{�ߥ[�6��)|���Nb����>������Uv�M�}�77m�U�x@���5���O���p2��e��Xafi�=����7S[s��Z���
K>z,�ɚ�}�h J�q�(�u����⼨�����F0�R���8�g+uI)���V�����ņY
�i��AJ�y,�b!^B�>���+��z��E#�6���7*	dp�Q1��e�I:벑�r���ѺZ�I;/��d@�g��̐��%HD6��jGdh#n�*�
��d��Z�;P3H�ۃ��N']⬭�cj�Im���'�nw;���}��UU[�����|�V���ۻ����^*�UUo�wwwu�UZ���n�h�I$��4�K4�L,�e��
$��~#E�r���[FX��3B3VcTTE�ٕ�	�E�S��KT�8�1�GrUڄ�-��e���Q��Y JSuUU��j���bՐ�G㫧33,���S�7�O��8���B����0�m좨�.�0F �`{�lU9C}�DNu
x4i�&��# U7��J g�j195u56"zaa�2�^�͉w=>�+���1��VKk r�",NW+�!	�߁"�G����8PǍ��j}B⃥�||Q&Sa��Q��dI�;�k���q�0�z���B��ՙ�'�'(��5ް�t��@�H	�m���}Hf�X�1��h�җT�O��4�ل63�>1qр�-�l�-i5�:�z��k--#��1��ۄ0T�,50ٹ�`h�=A��	�\x��ܖ&�r�Ep6�"@��\��BPY�IBh�ibi�i�Y� �6Y���;�uUU�>�M�#虁�5XJѓ_ͧ��$�DCG�������;����tz��}�/m�^6Z9��ִ��]����y���c��BO�?���x!L;����|:�K�����FK��������.,���I���|ifaE�:C�p�g�=�|/z���Vf��UUZG�ytϲ�2�h�p�*ƽ�'�J=F�3�^��[����KLɐ�vb���=FW(پT����8e�`f$��l�/C��[c�"�^Bl�yJ8I�U���I����ܹ��чۮ�t��o7$\��� A�cӷ��2��&�~�3a�g$*^�77,8ɼ���O&�~,�M0OƉg0�	,��|� �>�V���#�i�L.p�ۘ�V�b�Q@���o660�F�	b� c�)��l��q5Z�uZ�b�+D�D�VN
I$������1$K�X���UV��a:IQ����չn�vUi8�14GF��,,�L��񳜉�S��5���d*��kmZ[>�&�ORl�t�j�@�P���+<Z<bJZą�C�缊���������l���2�T�*���訡��V4�� ��MN� ~`*2�L�Y\�MM�vy4n�Ӱ¨����}e�Q��ibi�i�Y� �K5Dr.�DlUR(�����km��'su���M�{M`A�]d����=������A5�ь�H)�ܘX!�g�G�^JdC�ٯ���K���H�,HE�1�����c���m�K5D�>������o�n%�u��$��2"4�h-z�ϱ� ��,���aG�a��ㅝ:C�p�e�׮c��i�����ʪ�	�{��H1�>�Ul>�����r�@��띛�^�>T���gAL-�	���2[J�\2���Y�Z�J-���P4��>�V��1`�	����a�P3�|)�|�L���S ��0�jz����f	oV�|� �|QE�Y�Ǐ�t���e�u,^K�^:�DѾ*��'j�^�'�����eS^�}��s��5���!T�Íx�2�l(:tAD#�.��>�ox�Pl3C�Q���.	�L����X�5�$#CGܦ��Fx������qZ$�K���8O�z��Æ���a����3U�f�4����,��>4X� �N��69��k\�G^�`cL���q�,.e������ ����ۗ$G�}���T�X�,�ޝ�uӤ��X�T�f2cPCj�B*7Ex�U!�l�A�HP��Zڲ�.�X4��Fͥ��wʪ�	ric$���a�"|�4�A	�U|�pm�W��o��֯�=F��A�:�rh7="��Y��\�Hxly��z����t:i��Y9�9Θ��%�������R<|qQ�
9�<[��ۘ�̮
��L0˕9QY�w�=O�L�u��n���d$�ŖQgŘi�YӤ:'�m��m����c&�uUU�;M����$4	���]�V�4f����{��<�9>[|6	���sT7y:���Ϗ���E����i�\@+%���Po?n	�rnÇ��h����N�n����c���K�-Hs�X�){�A�p2T&#�i��_��ʖ��0��0L�0DD�Ĳ� ���K8@�"H�(L�DLǄ�(N�t�� D�:""9�H�$��<'D�1���	�:q��"H�@�d�G�!�A�pDI�DO%�QBQ�N�&�t�M0K$A�M(�M,�L4D�0���� � ��$��!8tN�,~�UϢc����=>˗�S؞k/8>�s�{.J�+�}~����_�Fş|u[�/M0�����>Zh+z/��^ݐ�Z���ۛr݇E;��ʙ{�2\�}v0Z�gU��,��轎�O�~s�2z�z�_9������*�	�K��57Rǽ����0NO���ڒbb�=	z^ܙ����UC�Ko�:�߻%���ۗ�w��UUU���������UUV������UU[������ʪ�UUn��(�ǏY��i�i�Y�!��,������}Eַ��BI�p2\:J,�����EQ�g�b�C�NCFü��s*9k��(WTSN��7���>�.��&��m:�v�f���pͭhu4S6>ò22N,_#��J����E�c�0�������`�h�p�0���ùE�����BaΪ��Y�û���!�������!��F���J��F�:�!m���	�M�����.�[Sgc	�s�&����d���Q����<�~��th棈����ZQ����!�0�7�R��j�$��M+�
k�rcR)Jū�ϣ����D��.if�Q�EY�ƘQ��dSrp�u�Q}�Ae�ʠ6
��9Yi�b�)�2�K����c�'��|��&\F<̷Ne��e�1�-RK[���ಔ��d����UT�t���^Zj��z��ѽ��]��!K���L�c��,Mѩa�zozx�6���E�p�0�JKGxq(�C����a�v;�Q�U�M^-����[������:t��������]��Y���Ɖ΄��+�g�1;��}�(��Y�9
��Ӷ��ʛJV�l��\��DL���x���g���'
��Q�����K?	�&YA��6�Gg��>�UZ<6|B�̦�4���q�q���GV�|W<V�@��R|ф�!���9�7�Q��Gĝ>D�E}�}��3+-n�fcy.C�_NB��Z�;4�ӹ�L^�����7<��v	[����.���EԻ=�agƉ,�O�,��0�ϊe��)�\r�G�`����5����F�<����b[��SgA���{!�m�o�
�ã #�զP�M���E��*����y���=;�UYY.���Ӛ���J���V��O!��4�S~%��s�۸Rq�a��l��������+�R<���F�x4����
�<%�Ɩh�'�O!Ӥ:<�fWӧ�3v.z�kM�*��&V�BBUOr��T��|0Wa�ܒ�����m|�;�R�v^&J��s(�Ҵf���������"��E�Q���F�`h��e�	�ǆZB�=�~^>]Z�!�2Q��3�j���a}&eJhC(k��poxDD�Y��?x�,D���//!y>���|�X{ZEp䭢�V<q�A��p-D�m��
ܙm.KJG��b�Ikj8雷�M����C��-�����w��C���`�#nӂDV�2*ڌE�D��b�J,#qo%��$�UUZ0ɉ���"�F�f\�T\�/X[-��x^��Q'�i�i�V�uZu==x��T��ɳ	��\;Jo�n���s����I`����bJz#$r8w���|Y$I��PB8���o�	����/6�a-rU�#0��+�JAj��uG�iH�,��D߉�Qf�b&�idaq3�&3̿].,��uUU��CE	�spÝ�'a���x��A��~��6I��uu*�1p�Dў�M^.�#W�2BM�{����a�ق3 �m�P�$n5���L
�{.���v�z�W�3�Z0i�t(�E�p8�+�6ݘx��4�񥈘"a��a�M�����}�Գw�*��j��jI>^:}ՙ�0%c�LG�	
 ������}��V����f;�:�f��w�^�^5���٥�n*�����}4h2B�ϩvŕ�)�J]IumU�x'���A*<t��8�HYΌm�"C�(�:��Δx�4��L4�0�	�<G�aBQ��{���ei(�&v���GV�>���B��:E]�(�Q�^IQ2�J2wc������������������+;9Գ�=Ȑ��C��OW�e�\ʍ̞&q��<4��Ql���s��4����I��b%*9�`�8x�4�񅈘&	�X�""abYD��$��D:'舞,K,O	�:'D�D��DD�<H�$��<"`�`�p�:'N	�"D�$� b#�� �	�:tD�bYtN��4 M4ҍ4D�<H�$����4�M,�B�(�&�� �"$�Â'D���	�����{�I�4AH����r������������!7�x�fW�eB��ve�)i	��9g���S�Zܩ�z�����ᖿ,��:ϫ��&o^���U��Vv�}Y=�����v��s��n�˷^ʵ`0�F:>}7v?Gqۦ
*�(��J�M��7�2l��=[�f\��a���
8B+deZU*���VZ�" �#�	����R<WXNYc�_����;�E�I�]��m�Ejg�]����lx�B�8="�G�Ga��QWU���&L��֋}ܫ��{|$�6C;'G����	'���c2��O!]	mFJ���݊�=FJ�@Zg�w�5���H�&=3ڢd�������qaeg��Pgu�gZu�}�5�hJ�	>��@��/;S����T�Ȣ�����1���Wk���4ℊ�n��8ݱ��F��J��Ȥ��@�9E"�hC��r��fC����)�(���Ul�x��X���ӊ��h�M9*���n�>&���bb��&�lO��2VY
��-cl�ݬr&&�m"��9	,RI\�����/dPF<u�F����[QJD6��"��Q������o��UZ����7wwww\aUj��������q�U���wwwwwu�V�����<ae�0�K4L0��0�.���}�&k�u��12e�t��m0lR!2I[�u�2��)pY��	�Тy�\rD7�n[ʤl��V�D:�5x��R�]���ɓ	�5Q�R\&��w*��e�q�I���.��.�2E%ݍ��z����4#��c7�Z��L�MX̒d�;T(z��Ov��Vүt�Ð��r8�p8j�ј@�<���/�yt�> 2_V��|�Hw�de�T��Hd��1f]�ԁ�=\<a�K��\�[�:TI�O�|iF�Y�|P�,e�p���¶�k���˻�)/�Y$���ƪ��DGu���� �o�&V�5D����Q��98uf�à��0�Ƕ�qΆh�{�!�R�y=�pu��MAIeI��������Ui��8]Z�L>��c5ʆ�f�>%C�ɤ�t��~�jd;9ϛSIT���G�L��,��E�|YF��&YA��<Yn����k��m��Wa.�����IF��e�o�*-)4x�Y�a��ep�Bg��5�YA@-z_
F�'[]:�)���� �C�ۓ�n8�2���Q:a���P���p��[��Ŗ��;9(\��0{�*��a��vh�0��@:�7�*��|�A�#~ �����$�YF`���A�ag������UWy6�]��:���qs�Cp�<h�`}�o�r�e�/-����d�k����Wju�TEh���_*�����.=�$���ѐ�?O�o���,*���J</5��`�f�{4PwV��Zu�2s�B�����f3c �|�,6P(��ƨ��j_$���0��0��(e�3˪-R�|�0�~��,�#�؞1��L���fY-�3.JJ�[3�і����9��!�i��ݙ1�x2�RK�QB�6��NF�,�88UVf^� ��B�QF�
됖F�:r��� !2M($�G�6�_R^,��0�Ѡ��rPG-��n�p�K���p���l]
[m�!�)b� �ӛ���CGMQ������~o	�LFT���[���^����;D�!�,����x��K4�4L0��0�8Y��i����/V6�;$�Q	�&ف�G�wc���s�錅���.�㳁�S�����gk�+R>Z���|u�9�%��ĭ$���9�Ԉ���Z�J���_%�A��T ��k��KQ���G��~(�|xa���"mM��0�ojᤐ g���G��9,�ό,�,D�ap��&��uKz ]�S�O���_-K~����]6�=����\V.9��y���nl��C���6���G�s"Tk�����۬m3'��v�4p�<h7*�'�.�.��R+�<Q�u���lիŪ�b���\*V�ƅ:��.���ִx�"���x��4K0D�Ƈ�����ը9�\O����|��j�|��%˞��y)�PՎ��6&Q�7WY���g��Q-˳f3�.�i	��T}]a�Z��+s���l�tm�l�<�j)�J%!}*$�7���Xb�98��۰�5�qu�.�HA�nX|��K:'�ıL<~0�"�Ԣ��qݘ\��O3�̙'l�Mq�Pr�.�X=6��^4kV��69��
�vZ냳n���-QZ�p�NNcr'��c�j8XW+̅2'�H4(�_uڋ�| [�q굗�H:�R���GP:��te�C�i����3��*zH��W:��r�i�1%,D�;5�T��7>�MG��ߔDZ�F�Ҏ��W*�+F�}���e�k,�WI��Q�V�j}����s~���>B��D�.S~),:x��?if��&40�,��U O�C��E�\��g�*��9����a��e��.g�69*�����{l��h�il�8�����9窿�����y��<��7�n#�ga��u�ĩ��|p8x�P-^�6��+�:�}pC��KʌE���&TG�L4�	�`�&	�`����e"$��:"""Yd"@���"&�bP��t��H(DD�<H�#1��LK �:'N	ĉ�I���$pA���Q5�,J ��8i"a�i�h��x�D�(D�L�<i�I<A&�����"@��8q�N��<'��ܿe�LG�jƺ'cP�e{Ԙ���oz��>�>���ow鶱�Rb7}��~כ�2;�w����g~���+���v���_�{/e��|�6w=7��-����f
��07*��_>�ϫ���{�V&=���i�;c�����t'}ߺ���);�l����}ȏ{�ۚ�짓s���98\u'��
�4�Ϭﲫ�F��}�7Ո��į���+5&�����:w_}��.ܯ,�[����{>�vz���s�2�	�����=����;�z��]��wM�ێ����UUK������*�UUR������UUK������*�UUR���,��4�L,�$в�YG	5z[m�R��!8��>��W,8�����y�Q�������x;!�u�58���6���\����r�a����t�I�pܮ��2���'ƶ�+J��޶�����R5A*B�m�K��J+�m�X�D�Q0�b���g�$�K(���0�M,e�p���}��\���j���ɩ�pMɭ��s��|[���f"cjэ�ѡ��E7MΒ�0��7Z��֊
A Jk�����k��4���.|��^F����ZS*e�ce6:#d�e�qi9w�氾�r��A!����i��Y�a�&40�,��zF�Oy��w���	��!��l�߅�#m\��v�G*�l3e1ǉ��b�Z�w�u\1�ZIk1b���إ[#i�t�U"
��LƘ��s�7k�9b)@�#��qZ܍���Q����<_ Jn3��ZY$!Q�J�uĤq#���[��b)|t��M�j�I��2Q��2�������6x7�?�����N��pɳ���:��f�]��q����?e;A��$9��k7fK�le Q�J+� -�7�$%�A���")���gO�>$�0�:l�t��,��eJ�Y�屆B^�m�W�Q��(:��0i�U;t,�4��*	�u�t|uЯV�E��z�=;Պ2=5U��'�~ �5-�y<<��9��٠���dk7v�-�X�`�Q��m�.�1kT�&�����\2[K1x@�\�]dA�*�G�Gcl�L4�%Q�a��hYc,����\�L�J��:�I�l���e.�L��dV�g�^�׎�����i�(�G��G�T[�%��r�M�f�?Q���:rB�D�o��m���H�����cc�I�6R��|A�:~0�L?%�&�x��<���o�sM��r�U�j� �ӘiP�-�EyF66��}�B��՟�S�?;�1~���l�]
	��fm�sW��Vp�/ʪ�n�A$t]��$�)�\�A$�̪�q�l�ɳp��ݹs�}�ܙ7:��Eb�M��Qtp�.N����S���4���(���+�,��I�O/��(�Sdncڵ��b4[0*m��"e-�H���+�U�Ё�6vClX��Uq�Cr���AR��9[��W["!q��l*r��� 2��ŭ7A��'��W
X�gL=	���4`h�K���J^p�^��l��'lk�U �U�}�9G`���$%�Z��U}�X��o��Vc��Uʈ����y�O<%U�Sr��5��٦g���OP��>Ew[�~68|i�~aF�YBvta��6ȢAP����(�9i���tդ�B��uH�o��9�YW����pl�NP��/�4�9Un�,�n�r賻�_t|�Rxl��4}��V�Jr�ct�3&�֔)�h�R��S��+=�FxQ�^Mp����^�6hTL���&�4'�ָ����t�N���E�(�ŉg�0K�adx��|����V1�e�[,��I%J��Tg�a�����h���6>�0��
�k���E*xX�'�p���}�=����Rc�14(Kc���"���ᙍgݞ�|z<!��E��8�F"�0���#���DϺ;V������5������l�Q�jT��æi��i��p��t�,�a�g��&j쉧Z� ��UJ�{� ��ķ� x�}G�}��w�Be4r��b�7�o(Ԓ�9]N:�R� �m��C�G�#�k��DDIz�H�NM��eh��K�U(��1dNҍ,��(k�y�6�6[!�g�jH_~,�WUq\�n��m��;�G�E"���O?h��?�{a!O�H�I �U���������鰸�g�ia�ňp(((� �.�(P@�LW���)�}mq@�)"�P���	5�A�Db1��(���A� �b0B1F1�F"#���`�D$b"0B11 đ�F�! � �!��bF�@)`�0A�#`��D�A���F�0D� ��Db"1�$��DF#`��D0D�"1F	F�1���F#���D�"DA��Ă���`�!�I2�0DF"#��	 �"#"#��0DF"!�#A"�$���""2$�"#""2$#" ��"	�(�Ȉ����� �0D�"2#`�����Ȉ��"20��F"�A��ĂȈ�`�#A#""2"�F�0H2#H�`�#DdH"2"""A1 �D����"2$�0D�"0H"1A""�!"#"""2"#�"1"���%��DF"#""0H"�"0F1ČDF �� ��A��DA�"A���� �bAb"1" �D����F��F$��b"1 �D`�b ��F �1��DB���Q`����Ă#���D`�##�"1�
0DDF"#"DH1"#b"1 �"�Db"1 �Db"1����"0F� �#bA�1���1Kb1 �	F0D�"0A�F��""���DF ���H"0A�0DF"##��Db"0A���"#`���DF0DF��D�AE ����B�( ���@�	 ��(�D
�H�J@�B !�� D!�@a"BY $���@BA��@BH���!�O�f"� !�Ma	@d��H����� $�!ABP�$A 	 ����@BD��K$�� $�H��� ��*���@`�@@�����	$ �� ����h�P,�T% @`��@b 0`F "@b 0@D!D!`��@`��@d@DD(��`�1A�	`�� �(@P`�d�B0A`�FDA� �b ��D �2 � Ȃ2 �F �"DDDA�AH�0A ���DA�AdB"D �A �DA`�1A�AdB"A{B�A� �#"DDA� ��b,� � �A�DA�A�2 �ADdA �dAdA#"�"�"�"�2 ��" �DA� ȃ"dAdAA$A���1�0A�`� �� �D �A�bA�����Ab1�I� �A��D�FD� �"�`��F1b�D�! �1`��D �F �Ȃ �`� ��D�0Ab ���B("@A�"Ab ��1A�"A�A#@dA`�0Aj�!�D`� � "A��"A� �  �� 1A�D �  �@D�D��1@b���� "���b �"�b`�����0@`����
��h� �� �� ��� ��F!���A� � ��1�`���5,�!��! 1�F @bb.�C"! A`��#�A�B1A�"��� � b� 	���#D!�b������"�@`� 0A�1��$��"�@b �F 0@b �$@b! �F �	�AA�`���b�B0A�0DF �ČDF1#�F1���8�P��A��.l&^�V��R���8�iA�EQH�X�1�h�5�����9��o\���ȞA���w�z���\P~����>_w�6B��'A��>�`\��o�
Q ~����z<
�~�_�W�]���P�0�"�������C��������`d�QU� �}�}�����������DO�0v���P�����s�G�?d�_p��=��hx1(�_�	����!P{����|��<BB)��
��;R?���`�a��4�a��n���3��!�K�%��*Oc8��D����g�/
hZ�s�C!�h?��$�_o��a/-!! ����<�����ҐDP���(U�U�Y��E�U�+h(� 
0�����A�����@�xnV
l��X.%a�_�~Scq�~ "@�! S$� ����"�jQ@���

����Ǩ�oއ���2m�C:��*�#�f�{�C����Xx���������!�����K�>�j��*�4�(�3e��~�~�'�O�����> h���0�;�&˃�� {����d�}�q�`�~�"�<o�?Xyx���Xu�O�����ꊠ>h{b�g����;+������pP@>��hG�}1J�0!���*������T���}�?;�J	k)�v}�A�7W��`�\C�@�)QL8F�D	<�,�]X<�a},h�7��"�_� �c�>j:���������E҇@�k-;�h8,��t�,A6��؟��T��<=���=��}��EPP[�0��B >)���x�����������"���|Sе���=��? {�>��� �~T�|���G�����*�>E'�)���Q��+�� ������۳��C�����O�0���D��t� 4�(��a�ן`��0� ��?;`��@-�!t�{�n���:�B����sX>S=�q��n�ν��EP$�q=<�<r^QLeD�bΏ |���0����z��۴�]����F�\L"�<��}K�_� �Q�A�+��~pl�;9@?_ߡ�|��j �v>A���C��vO!�g3A@��hk�	��%?2H��J
Q��`�G���������)����