BZh91AY&SY�$�
ۇ߀`q���&� ����bF��          ��(R�	P� ����(��ER��B*IBAUP��@��J**�JDUT�TH�JT�)R��(�#ѕPP�H�TT���(��!P��@J�JQPE�$�J�D�%J��$UI(AD  �T��I)\�J��¤��"`4�U�JD���T�*���� H�EJJ�!UJBJ�HB�*A*(�{*T)TU�   ���j���1�۸�ڴm�]�I+]pӛ�H�Z��K��E�wc�ݴ�uS�vm�0�֭���K\�v�J%*Q�kR��RQJUT��  m�(D��&:H
�r��*�=��B�*��<YҮ�� ��I��aK��"�U�T�
�l��R���j�G+�t�P�U(UU*��$��*�x  -g ���5{���JR��^q�GlD%Ls��օ"�������֌��=.ڪ*��{�UJ��y�!C��X��$������) T�p%DU Q<  3ު���G�:�V���yWL��{���B�U='��J��P���צ��xu{�R��Wz�8y
�*�{z<Ul*[����z R�D�PT�%(x  -x�R���gW���s#l�[��� *���*�U�'�綕���M�o{�J����%*�Vy0t��K��'��@�l�y���	J��f��D)$H��TE�  ��RT*�q�J�*��E{�U $W��m�R�=�v������q;��44�t��U*����r�QD��r��X��u9�B���������U�<   Zs�)	*�+B$��+
��p:hh�quJ�;�U�\�uʵTL:�� ��]WK���[�J�
��@R����x  u��T NL�4�\
���U���V:)��nWTЦ�wQ 6��iҚ@f�l���b�����*�D���U$ �  ��)F�Xt
�]�wTU�LEU0�@Y�.uk@s& En�P&�(	%��@��DB�!�`��UU�  l�(�[���E9��*@ұ�EP�Ӈ@U-��]4� ��K�QU�N�UR��{<�ll�   J  
 L�)R �L�10L&�b)�IJ��0 44�� $���&�)�����A�OP4"x ��H@     5<�%A=M4`C � i� B��I$��&�=!� �	�o���1_o���UM7�w���feE�,����|��7~s�@~���������*����@U�����������T��� ����4Q U���%O�� */��_�������2�!�������:ɬ:ì:��í�̚ɬ����ìɬ�α2k&�k���k�ck&2k�k�k�k.�cˌ�ì:��:ɬ���k&�k�k&�k�kL��ɬɬìɬ�Ʊ2k�����k�k:�ɬ:������ì����.�k&�k�k&�M�ì��:���ɬ�������ɬ�ì:ˬ��k�k�k��&��L�ɬ�ìì�ΰ��ɬ:ìì�ɬ���ɬ���:ɬ�ɬ�����ɬ��k&�k�k�hɬìɬ�ΰ�&:�kk2k��&�k&�0k�k&�k&�k&�k&���ììɬ���:0k��&�k�k.�δ���ɬ���:��:���ɬ�Ì:�k��� � :����&��2��� �������*�3���#��Ȏ����k":Ȧ���2#��k :������:�&���&�� �*:Ȧ�)�*k(:��k� �&2�(�:�.���"k :�����	0#�
k:����� :�����"3"��.�)��k:�������������*���������ʎ��2k �Ȧ����k:ʦ����k �����)��k*���)��k :Ȧ��������k :®� k:¦����L�:����
k(:����(� :ʄ�k :��)��:Ȧ�)��� :*�:®�#�*k(:ʎ� k����2��*k*����� �:Ȏ����)���(:�.��� �.���0���	�(��	�(��k*�0k ��.��"�8�Ȯ0����(�ʮ��k"�������
�k(��.��Ȇ��� ʁ���(�k �����k*��*k(��!��2+�"�(����"�*:���+� �k ����� ��.�����.�3�:ɬ:ì�ɬ�Ɍk.0�k.��M�:ì�ì�ɬ��3�8ɬ&����&��̺�k.�k.�k�L�&��&�����&3�0��k����2���&�ì:ɬ8�c��ˬ��c�c��&���:ì��ì8�k.����.��0k����&�ɬ��k$Ʋ�k���ˬ:ˬ:ˬ����ˬ:�1��ɬ��ΰ��k3.��ì���k3&����.��.�L�k��Ɔ�菪k�&͆���PΉA�tD&�Q�?�FJ^k�5��g*ޔc3�LC���Ӱ�V��z�#�;R��Y��]�Q&	P�Z�K-�զ��h����jM֨0i�Xrf���^ꙙ�������5����x�Y�K)e�x[k.����"�-����ww�WX��.�Jdɑ�N��ɬ���e
�f;�*����y$*k�:�D�M�Lՙ�8��!"����\��*�H�U�5Lڏ�r+/�+Zm�R�e�K����2<N��)����6e���Qh�f��7n�T��i�lLcC/2�N��f���mcK�A���勸�s.�Lಚkelbʚ�Pm��6�n��i
&~��zu��f��uRm���ŭ�Au�v� їCm�t����j��Pjīz�SMi�%ԡ�Ҷ#͜��x��Z3T�ALI^U<�^I�ƪ8*��[�X��5l0�bS4m�3�qE��b��;�d���[��T�ǕZ�p �-"����aU��Qf݋lԈ1B��F��N)�Bn��ۍ]�c�0#m����ХA�4�"^�HԕSv�@���	�r��֑K3*��*�w`hI� PH�*�P�qS���ܡ�6�(�˛���w�
�c��Jal,����ᲯK�ZT�[[������×�t����U���J�V8f�{���Cv(n�VMڹ-V��֓�)I��f���jSK)�&c�;[��THZ��B�cX��2�ub���ax��E,W���Ff��&���*5vʽ�5t�֌�p�s%j�e���h��c��!y�gvʬ�ףCm{QiV�>4¼-hw�1ѫ��.�&֫�>����s¢��۬�+h����
�O�Bi�J���'lϵ�ܰn�i;PTt�мv"�Ni�[C��"�:D)(��Wcs"/u�[SFTy�Fu��Ԥ�IR �T5�v2��֟�*8����wW�tuJ8H�Ii۳
�>Q�*L�su/=�bm�	�è�F�8��t/�v�Z��fb�����W�(�BeD��5]я�{O0���ô`%Rp�8�jк��NP�6;xp��m���!n�)Z��]���t���/.��+%Zb��M0�{7Ս��2hj�HL
�/(r�cwr^�9*�н��9��a��J*ݲ@4 z�ɠ�Ia ���ւ�3B!]l�zFՂ֤�ɹ������Ȗ|o"�L�[Z�"L:9^�"���I��׆�[c�W��pm7t�/i�3hӭ���1��A�X���l{mWYD�8ٹN`��mK��N�ifa��7wÒ��أi�V�U��÷�h�ւ���Ŕ�Q���bnSw�T��	i�KM2��z%��:pÉ��TJ�M�)�Ӹ�	�k�.]�x��cZ��t�,�(�7GN�Vk(LT6K�2����
,ক���"++NX�Ŝ���=���N�77^A��%�����w)��~�P�xr�M�ܣ�ûjRd�é)ӵY4�1Ƥ�<ߝd�u�j�3)��. Ȥ��n��������7hS�%�&n�L���%��"��b��-*7V4���NZ�d �`���R!��dV��������5HP��J���F���2a�n1���mTH��!.�N�2�x6zj�r2�����)���v�W��ZmQ+f���`� $&�r��b���H�R�M�Ym��`ײ��N���Q�E6ȭ:�ҵc�QTvY�SV!2<V���ݰ�{�L��7tU�2L���L2MĶ�S@�3���=*іkH��D2�m��nH�Y��R�I��re�+ef��%��e[�6-Eki��4�c37v���ut��Q��M�T�w��1��mX��%����Ga�x�eє��؁�me�ն4�EDV�v��(i�VN�L�Z��*�+f�Cpm���.M@��Qr�G�Bj�Lwqʘ����La�D%������f�U��p��C��(�o]�Unk��F��b�i�0��S�DjL&څ�M��~yN�h�-�L��t�,����L��������/*m:!�;67)��^�eк�*ú��kyqnU֍��a��n���5yX�ٷV.Sѱ������nL2��b��b�M,�t�}��j�J�:Sb�%x24�N�a�A�H���Wg^nQ�����h�V$�"Ҙb�1��S��U��%�Q���m�q�N��ҥ��, �R���L�L�U�o@�������D[��5Q5qa��[:�b *�JU�.8�̀�(nU�Z�����`^^Juf�q�,��t�,LR=�9o5lfT[�,�2��"	Yf�lX�lm�,+��� ѻ4���%	�Jx)�W�X�
Rƴ'{�ZѹA�tB����$r(qV����/�2���;'5	�[��n	)�KV�LˎѬ�Z�j�b�L�p�@*y� �3������+�լ7��Ѽ��`!�iݢ�*D�ԛkPZ�̕`��·(��f���*fV��%�$�ݺ{.�z[���6Kњ�nN+.��Z�R������`Q�y�&hʿ��ג����SmF鷗2�5l�\2媉�Q&ֈʫ�(k�Mb;��V�Z���@��c��Sz+ML�����G �J$�"�{�(�]��X.�߭�����n�l ��p��"�=0s+cX�Zʙ��]ẒQ�`��0��׈��ǵz��{W��K��I��b�˂�2Y�[��TZ��]�!����u	TS#k�n�`q����0�f�S�[�C3EcZ�:�ޛ��8��+V�okC��Z&�y�.��^5u OPuh���Nl�T�Y�EV���ג�cTvV�SͶ�S�-;N�Su�6����Ʌђ�����kY��ͤ��V!�J�TA�07�Y��J�K)���w��� "A�����wZkXZ�yOkR����&��L��k^���Ne�F�v#����oE�L���V�mdz���Ǝ�5�=�MY�x/�*�ʺ�]��2ܷ�qo�KCF)��)nO��I%���vC6ҡ��CA%���V0��j�̭��V'������%�Ŕ��s�e�2����mP�p����	��մ��ش����<ʊ�)�JɓHE��*�dx�*�e���a�W3�B���#/h��,�F�J[���wsl�WY���G͆6˩r�׆�MyN1�\Gn��g�a7l�i�2w$
Hf�5;�J�^'�⩉��f�hY�������;�Z,7W��+�(m��I�kT�L�n!Q��ֲhL\͔]��/F�f1���$CK4�!T��s�k6���jk�GU:.l��a��*�];x2��]<��>�ȫwN�G(0-Z�t��e=	T�V)�-LI�oU�Q�7���)l���L�d�;���i�A�Չ�`��54����	Ƅ�����j��Ӵ� ��j@�Mu���։�e8u]E��"�Q�Si,.^#D��R�n�������3h���үje��f�Zh�����V������v�Ï
r��=6N+�׭�(�X/��� 
G&�Tr:�a��e���"�0��a�e�
��fVf�tԬEX3 ي��3ql�P+fk^2"�Z���i�YRMT�7�'w.��b�KEm;�����v\ ��m,���@R1�A�C�6ֆ���2�
�i��2D���ޙ����ұ~~��P���L��X�Ko��ț��`�a  {�g�%���-��f��d����ZMA��-A�9Xz�
���V���+v��J��d��;���K�4F|k�c1UZ۫��UYK$řS@���Q��`�Bʚ���j���#F��Z�y��^����-jHd��N��f��$���r��h7J�%f�������-�4ͲtӐ;�3(�i�+Efo�Ջ�x��jF��s-�&��v���KY�����v����Y�	sp�U������K�ښ�<Ъȗ{&�b���&���Z[�,e�)�h:��	Z�3*����ŷ@c�Ne�@�r�+�nA-�S��d�aC4��7�B�jH5�s`z.�T�JY$�kU��M���^yjgu�IX�����]�JU1�N��[�r��#H�� �X\bVnR4D�F�0^�k�_8j-�$m��Pأ6�'�˴�Y�&��#!��X��楛�V�g�f%XɁBoP��3M#�\I^]�C\�V�Ue�h�=u��X�-�0���1�ti�R\YQ�9@;+�\�kr�1X�zj^)V�n�i:�i�2���6+0-10��EZI�`LKb�\�K[�C6Xv��3�#�N�U��ԕ�I,�Pa��LXv�IM&��7y)b�wE,W�/�3�A���`�Z"�R�lJ�fR<²A[��X�W[�Ҁ�qX�jX�9z��n�p�X;Px�l�"7��t�W����Dضe��<�-<,�Je�o5���]�,�n����J��K��5z��W-h��YYS�n^��ele;"��mYV���Vmk�Ʀ�Wx.�fd%�*���F�:�m5v�ekF�f�������F%Cwq�ɕ$dd8�P�E:/t
��(^l"�W�e����qY[[x�O&�~9��@�654lэ8�R���;fj�k*��q�9B�����5�ih8�+:���/#GN5N��k*IHɺS�N�j�)�K^�c)nk#*ʠ�)h�拙@�:Wk*��)kk.#
�v^\$YAK�r'Q��u�,7�b{����\���t��j�j�wI�t�z�9��4��p�ك.���(ګ+���
�=�A���Q��C� W�=���Y���7�j`V7��D�BZ��B6��ɂe҅�sF������p[>�,nfN��f��ښ��Gn�Gjh%6�t1P2�5xb��z���r΍��%e&R��%D\���kn@�R��Q�n���`���gvS��D"�\���-qn�q��	��'IB��2i�@G���9Qڛr9�i7�Z{�y(�Zٙ�\� 7F�w�d��o(άv�嵢PYtQBL���Yw���yx�[�6��E�sT�Tֈ�L=�Zr�ɵ �&]&�8C�$��g2`)<d ���o`4N�U�g����b�+����KU���2fj���6xj�7�KR]CGS�Ǖh�����rPͺ4�Cne�@�*dT�3rζi<cj�r+uOAR����,<TF��r�ǋP��V�Bdі�R߫1)Z7&���CiB�wv�L!�w��y��6Rz(PJA@-�Q�sz�du���"���BXu.Q��Uy{G‍�J1������y��Y��Y-`Jts�B�Ń=v��m��ìZ�95�U���.ZYe���&[��.����M���i�E���*歚�FXTUw'a9)������6�Y�2�6MEh���m�4��h��	��#�n��C�1,�^�I�����*�eշ�R�	HG,�b�,��ll��hZ{/km�MK6u��{{@=L��@h��L���z�T�;1d����
uy�(�FZ�dǒ9�p�2AF.�FC��Ӭ:e[ݢ�[IKˋˬ��ZB��LE���^��1�)���Y`]�i,!�'dX�O�*��x�TSa�2��sv��k�W�kY	wF�R[��,� Z-hh�,R`n�p���̊�KQ9�(=�w+e(���N#���Ǎ)OE0f--�I��Ր[n��V-C1�^�\��i��B��8U-���݅�9��K$����ċ�`�ܷ7^�G�⽣����Ҝ÷KSyj�f�DE
�Ʀ�LHejh���n����N#mD�C7���qGAÙ6b�R�ϳf�ʻ�ȠL�m(�C��:�R�"֑Yz/0���؝3�ƽ��BE[�	7Щ.Q��3[�v�M�ݬ�L�:V���[�*�M����-�@�h�����,��v�pnG�y�ڰ�����#��.��y*Ż�Y�7ͅBU�6�������l����Mm���L�]Y���V'�^]� )8�zm\Ɖ�g3��D��L��l-�n_[�IQ}B��#rX��`��s�R�ށ�;@����v
a���I��
��Z��r���&J�J�k�ЇFS�r����xK˥���á���Z������C^���U�T>s'|�x����İ��Y{}��%��&I� է�0��U�|�)��E���(���{B�I�XQ�c��&� ����������!��a^��4�p��K���ڥw�2R�jW����h�O��T��4E_Q$u�a��EX� �V�C�A���3�����\��B�avK
�}ä�8	y�XM��n�tZC %Щ�J��/5��ˮ��M��=���W0��&S%�D�Vm��j���ٛ%p�a/M��Z,�
��]��IZA�j4��'%gܹuR��V��V0J�4�2(N&��AN�n���3�i���̍���\6�9���6y�d@q�)�,��Y(��uq�(�0��ݡ�IT�3�%��
̜z�����V<�-�զ�����P�����1�Q��ή8y��l�E8V�g��a�u�� ����Ɠ�}/�>�6�Eg���`��m���] j¨m�Y��Rn^ 2��+4��g���)ԅ!Q�ܾ�aз%�2A�g�]Պ)
�cAR���v�(fl�r�e�F��Q�7WGh]f%��T��JY�5� d˼*Y�r�g��5�h�NMf��⭈,�qYO��5t[6[ Qe���oU���A<� 5G�g�<�p�9�`Q�\ܘ�\�nx�^��z*���=?��`��WVϊѕ��MK�n���N�5v���?ُn�3���C(�/���-��k��1��e�f_WL�9���	:�ʂ�5M^X��R�#9�V�WI��e�k͘��+Vu����z�@a��q��S�8J�:��d��R>��;`�-�|�gvk������XpH��\���Hxs��h=�\�D�S빢��T���Zx�ۘt�tyn3Xs\f����z�N�����!��K鴏R�C� � n��\���0Z�(3���=t���ӭ�����P{F�<��2V%�L�i`��_.��'B%NX1.Zڤ��5�E�;�Q�`^�imڎ1���ֆ�t'^IP]����U�(*vZ%vs�b��&h��Ft�$L^�s���uen��V����^<���2p�N$7e�"�����ڇcڒƛ��5KEeLo7&&��� ��f��[��������;�|��+��.V[��a��7��o΃S���ш���7�B���%^v�7 ��/�f��n�ЂSV�J���m�����сr�N���gW>����e�֎>�[��g:%����*Wn���وv��vr���v��� 3)���AfK\B�|�k�wbRZ&ef檒�5sk�jJ.�:����VRm���rƍ�3}&�;�VQ�nc���\�+�kQ��{���Ք���ji�waf�q���c}
u�ޔ����6�P�U����e���,
KZD���B�Y*��iZjTu�vR���8M�{����n���K���|�^�y�Ջ��jF�\Ou['�H-�#0Vsl����Uň�79�,�\��rٹa�����a�ggqe[�Ă�{P{��W>�}v���Xףo�#)�*�>Z��c؞�#υǿfK8��?c�J�8l�9G_]����D�c��ML��/p�j8:������[�}}ylڈ��űn�_m<8'=�{�q��\��߹^Ȩ;�]I�-�h��Tە1ۧe�d��	p5�DQ8����iD[
<�u� R�P��
&��<��B�V	�u��#x�`sۂ����eCK#��4��?���P����H$�?}Y�oVI�.��a��u�ˋH�*��KX�YӬ�};���}Z��I]L�C��7.�z-�1kj9ғ�[Y�Rצ�$�O�Ng��·[R�Q۳�N�L
��� ��+2�u����,x�ٯ\ո���.e�Y��r�,ܤ� \�v��V�b�m����)�>ܲj��yv��Pr.���(�X&S&�c�賊'ICQ�2��;��cW���Qs�.@�c%�H�`��d"c���v�e���bGEv�#/�n�)��1�_s�',�t	�p���e�E���Fo@�s�=��5��J1�Y��p萣�qR�]�]1C����j9R��zE��[Xh�t���\���/Q�bБ��2��,I0��+X��-3'P����sGj1ֆ�N����8��/(�*� ]z��N�V)wc-D%��ݎ�N�r����Q�Y��Rws��OVl4 ?n8�67�'C�	�����F�^�wP��C��mԊ`�cB�m���Kz���sh;5��T��N<6��jP��b���f�Y�M��/��oI��)�W4D��s䁋r����K������i��4u�6�w�
�6�TZt�tۛ��֋V�8릁�dGe�b�s)�_-���,.��LTtC�1U�El���zZs6����֒�j��3�d����R�q8m+��bPa���Po6�N���q�
�P�tm�\_�b�c5�ހ�U�g�*�ڶ�<=����>@*{�m����f��U��3�	CĲ؀��)Ǌ��Z��\*C���8��:��[� b���s;��R�c-ɍ�a�B���#FV~���y)����7�.���g0hZ{�t��)VF�{�,�ܾ�����\�U��	��);��M�^�1�@u��MO,��"I�p�f��U��v4;����N:FA��/�.�Ot/�M��ѰF�t��PKw�󻅞r5lr�f(�}8*�p��1�®�7��0`.Y����G�/�b}�j�GC}:,�������{��Ӻ�:8�-+�U��Ϡ�u��X9��w�t�J�H�t��lER��B%��VVnLy��5�w;e-��rӥ�b5�D���g��KHhP�ej��B�2��}�#1�X�Z�����{���Âݽ�Z��7��2�y�vk�{�#GWL7��k� �ܟp��ef��h��\jMTU]^�=�kA\>���֕�����n��T����e��!���M�����̰zH�Ph���g`΋q���K��:�8Y����\*��Tf�8�K2�:�=	W�;-�b���5����M��j�B�b�"yu�mwT���f��t+vpRrw�Cw8��r�����9�YV)�5s�}�:�D*G�Ƕ�zH�)/ck�_ut��+�Ɋ�j�n�"����iq���앇�XW\���@R�G8��YRn�8�RL��I�i�:��'s!���D���64�[m�������W&\큌>��[vk�	��>C���Y&2�w;�{8SR��8V���Q�\Z��=z�;�w6{�[���X���j)@q�2��#���Ln���\��D�V��j�f
���Y/�:�d���,>���CC���[irn�+K+/r�}.�4Q�p����Uk��'=���wFi,�rXv�� En�6[v�v��rR\+5,((�{�6���V��s�sǦP�;�=%�" i�a��s�e�z�;�ԤE�ݨ����ھ0�<7��B�Ur���뮾��j����bt�Y�;+�k���Z���s4�����md�x�Λ��y��:�#���4c�qB��D��^GS����a�I<�=Q���5o 5sԫ-����]�s4R���f�ۼ/���s�z+u��Y���F��/7������^�����\z�NY��mm�4Ti��AHiu{8֎בiz��I�2���4����i�=t�����yة���5q�߉C�oY�:RJb���jh ��cZu���V��i��1�b�	ث�A%�� ���6���)�%��1jΜ2�#
�2�� �������ћs[�fc��9)�*Ɏ��m��"w���iwW�>�����.ĿM;[��yq4��wfA�9��Ò�Y�t&�q-��N�L�����uʒ��Nm��lin`�S���
�6�=1�l�.�������݇�ֽ�<V�܂Z.�Q�[+�z�cP�8_Ww:H�-bЖ�L��fm�:�J�[���<�Ǎ`�uc��(��,{��n5���f>�.��*Y�ύ*A�=�1[��#5�.�1���Wg��y�g7�� ����[L�'}�O̷ƞ_n�Aӌ8Mp޹j��>��ej�g�;ن�sW��U�����LYh;=0���I��㣪�6���M��խ"ή)5�`��W����u�e3vUGH#+U_{��T�*9��au�NM ��؛U��6���'u�S�/@u�����r+=T2�0��T�y�z�����K�~�}\td����o(�*q�eXe�9l������r;��
=fdɷ� 5yF��.̿4�wn0�*��W'��X��%�__ow1ދ2 4�V�Y:]omwf!��M�5Κ �F�4f���K�Ҏ�ı-k�%��ΘȤ
U���Q�j��%.ݢ�i!�Q�4���ߺ���hC�2�Q�X�Y���EX�Wۦ�f]�SI�=���j�f���>ԃ���r�\-S�9�zV%7�b|$�HP��˾�OG+Xs
lP��t*|�@(�e��3�W�t.��EHJW�rX�sig;~[�J����S:X��h�B���.�t�b�*Ч�S�7�K@��G 8aY{� �3^r����1��F�RP�u���:#S{�ߐ�L.ܶ�� x���Y��Y����X�??�=���Q\�b�&�bnKVb�Q����ȫ�(�"�
�uE��<����ofƢ���B��q��a]rY´R��/��Ϣ�mX����7Wm�L��=�d��W��R(��7� [����#�6ܩ���}�Kz�*���f���Җ�gk%ԭ�ky�c��s���ĺ�sC�8=v-b�%��ֺN�q�hԒ��U��2��� �Zt],��xW;~�`�3�1��+� @U�'C�!��b��2�&����h-�鼕ҁ�y����/�64VR����.zT���N���;�l��t-ݑn���	��*]����Pm�V9�7i�,L��*�� �R��]םf���*���u��l��iWu���;W�1�cw`��Bm��Ĺ<-\cl�4����{Ӓ���m^kO� y�8�%(���y��Ou���-6���u��V��X�V�O����s"y�29IuᎴr���g�砬��*ݗM���nUI6�Y�ט�.�E�� *�8D�w<��w[�cz2�����>� *�n�tV���2��j�K�{�҅,]������Ϗq��YV	Bd�o&Y�>������R' ﴬ=k��� ���+�C��QKz�ը/�Y���:G��R.<��1�ݗ��'|rV��}QN��,ۥ��olĘ���&%��`v�IM{q�8�S��q��Ý�AT+	''�5*�ʀ�cP�<r#ǉ�PS;��M�ʻ���NL5��b�-h5�:2��g/tӾ�t��X��J�	���4,�X������svt�ى���AW��C5̮7���F��ns���pY$�E�a��˟v�,��5��qw���ݎ�qq��a�Od~;�<Y{s�}-�r�4ڸ���Wn!)dn�`���	���Qu}s��tHKq]�)< �VX�N�yڪ��Z�Z�϶�e$A�bP����X@윍'�q��ʹ��u�Q�ހ�a��`}�7Pm�N���I�_%g�E�/&D:��]	Uss	E�����sm������C�OzU��Vl�]K������q��p���_�	%��jb��"���;�>�6ٷ>�X8U��%J[_r��e1W/��E1�][�N��|#�OVս/X�N;�CI��z� ��%��t,P�2����ea�������Ĭd��}�8齎o-��[�҅f� ����7`�owYB�Q��Ⱥ�me[�M��0+��m�ˆݣw\]��$ZV��4�s&�,���>f�qS��&�K  .��W!u)	�{ԛ��U:.a	K�Z�G-�7oos�U��`Ǐ��]�PA�MڏB�k�߬�yA
��9ѫ�����'�Z�����#�ۗg��8:@����^�S�wb���y���U�[t��^ӝ܁��)�]( ����z�a���D6wCʞ:�l�dW��\[�,[��%^X�9�i��Y�J��$���θI=���kV#jd3e�[�u��"SU@����ї�Ж�V��x�R�i���zL�Hwe��;�/�C=��V؝�-0q�Y\E.�J�>�y�o������	R�C�\9�B�O]&�v�����}�t=|SL�.*�-[�3��qf[�1���^�:�5���MǼ�͝sXL�Yj�&��MbUΚ�N�������>�yjM�ڸ"���&mh�+ǥc)��s�,W�����	��m
Z�i�f��3)v�i� /Ta66�2r���*��m��ŭ��}|�e��t�����,�E]G%�t/�D̢�8����ng^��CZݫ�t`X�m�=aS���k�L��V�X��nQ��r�[ÏK�-�vy_a�~��aS��hRJX�l�
��\خ�\�K����v^��+��o��Lw�16�c�����f�,��Գ;_KZkXumcԗ$�޻��Z�ɒ��<�l6��H�R��Fu5hjqf�V��U��,V�c�&ٲ��à�@�kN<�E�g�9�}�RW�m.!��q�6�B�if��x=敜,�\��F�<�Y�[���ܷ8��7¢=���/���qE�c��9�l�y�n�0K�o3�V�*����+K���` ,u)>����ќM�|+����t�Qm�_*����<�p����f�]V.�Ba�T�>�xm	��tY�K6�q����WϨv��e=�w]k��rT=fo�L�]��qS�'[�1���N� �.�����d)�*i&e��"�G�D�!Z��`�Ǌ�m����=jT�t�$-t�H��� Jr�!��B{HD�Imv����Cȸi��
���)F�ai��'ҹ����R n�9��4%<�V��!��q'�����*]MXT��h�]hL4�+F��)�I`��c��*_�	��P�t)��]�PJ���
�hCTZ�PD&�܁���
N�%�f(STh-: �u9aVY R��)�yۻM��Xd�x��j3pQ6)��л��wr�%ln�Y� �i@<�H�'��P�[�`t� Q:�\�(� G��2b����*K���t"��"%@��^[tr$��WWJR�.�<������r��) �K��DaM�Q�)F�v��	�{bn�Y�foe�B4�EQW�)�t��!�%�y�:Vn��:"�e��) �=��kL��Q�g�R)R�C�:p�RN�&��t�R&�4�ctITt0�
7q(E!A�m�9�Van�'V��V��d}ה�6��3�B��J����w����UAD?_�߱�����O��P@��>W�.I��b)$|��$otN�6��Wk]�(�h��k<w~	@�]��AGU���g8����`�hTp-�H�ý:�ji2���8���	T�	�Υ�ѹ����ڇn���s.r9F��E.��[��kSd���{�I�W���`!���3����T�z�݅K7z�o[nD�ui�Qej�-�Y�&J�-������v16�=����X��F��]�g�������e�t�KUe��S�1��w)��|q�#L��Jݴ�T#L;���]����+8�QC\��x���3����Q�^��k!��%ۆ�J�W�[O%��̽w.f2��L�v��g�;����*E~��<��c�'�<���zJo���y�_��޵��rT�}(�7�CT����˂�=F�內�c��ܽ�XOl�uJ�|vR�l�a�\�&>�=�w�ܵڏlwb{ �j���|.��A2���&E���ɜ�ܱMgk흳��f��R��M2���1�غ��=�{�딶��ٷY����(2�̡b�ʕ�C\�	�����ĵ�u.f" "$�'+(�����[���@F�A�"�VF��I/oe�Չk�P�ӭʘ� sB�F՚�\��捽x���ǏO��ޞ���Ǐ<x���<x��Ǐ�<u�Ǐ<{x��ǧ�<u�Ǐ<|x���^<x���ǃǏ<x��Ǐ��Ǐ<x���<x��Ǐ?^<x��Ǐ<<x��Ǐ?^3Ǐ<x���ǎ�x�Ǐ<x����x��Ǐo<x���<x��Ǐ<x�<x������u��~�_��<x���Ƿ<x�����Q��,��%���T�k�1-�2� [��N���x�N��E����KL�:�g,mp��F]�����+r��y�i�];���6�DΘ�R�]3�{Q$��Q'΃���; kY<���wb����626��p=-�`�K=R�t��S�t=[J��uI9h����s��Wt�����ց����4�X��a׭�\{r��y�e�u�%����=�a{�^ZP�r�f֏'b4{��ռ��Z�@-\]�HI��u��g%��8��q�zxӭ<����d#w����pgLa�Թ��x+q��bn&�0�:�ӎ��x�an��e_J��=[�8j�k�R.6R�հ��47l�P<�b��U�LjWM\e.��_2v�5u�R����;�9f˛���H��ytJ�:�ZNe�3{);
[��C�������Q�w[�5���YN�K�BY/��ȃ�r5¦���f�h驺�RȺ�k��ܷe�����	J|�:J?��1+[�{W�(��z���`8����dm��iW6	����:��l͆�s���VP�	/8�5�}˺���9��/iZ���8��ٍqS�R�I�ͷ�_=��wP�%T��YJ���DE�B��[�UW�Ç������_�ޞ�?8��Ǐ<~<?^3Ǐ<x����Ǐ<x�x�Ǐ<x���Ǐx��Ǐ�<x���Ǐ=<x��Ƿ��<x����^<x���Ǐ<{x���^<x���Ǐ8��Ǐ<~<x�<x��Ǐ3Ǐ<zx��Ǐo�Ǐ<x����<x�Ǐ<x��x��Ǐ����~�_���Ǐ?^3Ǐ:��Ǐ��;��ݧ�k��o��1�6�f9bܺ=2�R�Du�A�7\κU�Q�O)	۩�����ߕ�f�9�adn=����S���&Q�7I��qww+�XžIm�^��1�r�ec�u�����	u����N��z��j��k٩f�lQUw0�u����}�[���C�R6��'�M���\�"�[~5�9�
]���n8�z��^8Y<W6�Fl[e[u#�4r�!�5 \&��5��{[�2�[S�o�ʺX�����M��P|���;sd���Hѣήh�VgZx8K������o�J6f��p	��ء!I�3Y����0!C\��!-���{fu�1J��K���ͻlխz ,��cf'uk� ��zݣ}�t�F��!�9���͉%�O�楹���vwEѝ�@qw���#���{uv���,�`��/\�TD�(�d2�[����M�\{ڻ�3�Q�*��{������j���\4ө�ԓ�!5M��XK&���Oug�\M'V�[5]�롃�/;�{j��t�%3 7R�X���D�2r�є�C���&jwِ$�O��Geq���n��Y��7�*d��)��]�hB(�A�R�F�xo�7������~=��]x�x��Ƿ�<zx���^<x���Ǐ8��Ǐ<~<<x��Ǐ<x<x��Ǐ�<x��<x���Ǐ:��3Ǐ<~�g�<x����ǎ<x��Ǐ<x�Ǐ<x���ǏO<x�Ǐ<x��x��Ǐ<~<x����<x��ǏǃǏ<x���ǎ�q�ǏO<~?^߯������Ǐ��<x�����˛�:����ֹ�rt{�z��)�`Rީx���x֫�K����˦�9:�yÇ%�&1�ɑ�]�%e]& /3�Auep���S�.�jw�]YWΒ��ue��;�`ns�,YWX�W+���o�y>F��m�(f��+h_Z[}[V��C%�(إL�e�w x���L�:���ʙJ�_17E���et��\�%�XO!�d�< =���S���Ռ��d}K4���try�S\2s�Z�d=Ӊ �%�)�=u��iz��vP;}z3'u��'�M�e���[wԋ]*��ʮ����l���),�z�0�]��qe���N4��BU�8�fe.���v%'y��ȁ/��6"���Bi-c6�ޱ�^SH��6`"�n�"9�d����~�6d�LƩl]J�e�^�,���Bf��Va��Z��*HyLI�;��(qնV�d��4:��]Z=']�R�[C���+�\ŗ]$�2��z��EEt&o�ѯ�Q�Q:��ïS�6λ��O�,�nR7J�<�'$�k���h�|�v	�~7Ru7�����lV��y�|.�hZ�u.ܲ �����G�K=/�4 *ː�����̇BP���T��(��|l������,�[`f��?a���β��_c�ճA"Re�i_>]*gv/v���z�L���[k�5EL����V�W�E�̷9�M�n4�Ju�3�����bRW��8EUU�͠&tR�[1-6/s:���e�I͇3��J�#Y��^ ��]hU�(���B�е�.)��-4����C0,Z/Z[�\S�]���r���_J�e���h��|��@��Y�'���J����xX��*�����%Z'Y�u�&��-
�Q�D�8n&�Ջy��v3��x�^�0��I�<Usj�=�ۚoz���9���S��HLK{�����='��4��Y�H.�[6b�f{m��ބ(j�������(��#��H>��A�2E�<�Y��ns�+�JZҹK��@@�%{yGH��wAh��ש�*�_1�����m��SV�^�푢xT��؝�9Y�����m��;�����Q�
�(�)J���YZ�.]��l��U�zJ�u��W��k���Q��;�w��y8y��m��/-�:����9���v���a&otȤ֘;��>��� ��= `��I�
�bp�"���
�S�N�\:��{/P���6�Yu�b�t�շ���A�X�BX5�R�������)0Q�(�knX-��
��P�,�p"�V��kԙ�{�Hn��1b�ӊ�h���u�Go`n�Z��W�[ `����uw���<T'�5(hK.��t1]�U�j�X�9�ʇ���:�z��Ԯ��P�K��:�u�����a�� ���YyB2j�7{���Tk��7�Ǘ��g
�15�l�7�jp��Vv+�_=ƈ�H#OK�����.+��gQ����3X����q^+JmYf��/�0����Ħ�s/�E�h.��yH�7�n����zhn��;Z$�&�Q{�Dք=���]� 2��{�%��v}��8fT�<�k�}4J�@��䈙_ ���S����`C[�m�a�Z�U��|�Ҫ�Ga&C�V�xν߾�L�Hѧ3����TA�:w��֨�ApӉ��F���P� �N,�/� Mּ�x���!Ӽ�X�)��fv(i}Uq�5�;-�2��z�3�E[��s%��b���r�!ʣ�j2�[��z:���sxλ�p�1t���N��̼�
���+Σ���eg!�@��w_}�*p�ʆ��Y�Roa_Q����D�եpY�Z8*z]l��U� �ʬQZ����Y�X3��9:����x{�Җ~_�U���Ӱ�Ub�xn���/>��l`�l�43��^�ْgp�H�Ֆ��Q�А/N6B���f�.����8)�z�F�orΖ����`�x�ʝi�O�U�Y-֎	,�G&V���U{k���z��HXnd4n�"�"$��l$�q�F��2w�u������6�����Vv�L+��Sby֥��nbt���V}.L�a_N�z1(��t�;'5ۂ��+0IM�66��S�̢2�t�ꩊ*�LT�o��jP���tDdi����t�р���F�U,��h��T�Jۻf�i[v��Չ���Lں}��&j�18�6Ƞ\�+Wۄm��ԝ�	��Ɯ�,*:(_Z/���ѽS]��F���&��m��m�>Z�Va��+�=�u�=��f.�V@�s�e����-") �wC%#�-�x|��!wQo��o�5�iL �G5���R?��f�llЄ�J�[X�j2�}��f/��ӍЙ��Z�mz>WJ��
�����6%<��P�6�s����(�U��a�5�ֺ۶��c�J�/+at�ZZ����+���툴)�r�^Y�"�m�}J�vi��tWu�R�xo�u.��s.!�w|*�<<��]A_Ph;��:������.`�G=N�s��R��gN��L�f�N�JΘ�7] �)ĴU&�c�F�Zl�;8k�y�@dا5!�rЧ�f�S���y��ok�s�(�dp�ʍY�N]���`���ŝf�2d�Ǿ�O�*��w��u���}W"�#Mp�r�}�oVegB����`�"u8�H�=��2�z�×�43v9���>�`�	){�y�B�C<�35�z�d��Y(�8[|�����D�j�u(S B��iv�q�G�ӫ.�����o��<��1Jz�� ��j{�me��3�*��+;u2�E���a��Yֲ�4w9P��QmVSc��l��>���;Zʭ�VDy:ms��,�����o��Y����v�q���'t�$nEփ�avչ�FsV��G\^��f�c�\��0ㆆN�{��%p�|��a���2!W��FB�$U���U�/@��m5fժb,�8ӦCa�;�mZ��n�W+)�x������N���\(+L�J!�5=�)Z�ձ&��o�b�Uo-N��(���y4��fl�(>t�ri��!�]֫�ё�f�``���I�^�N��h��%9w�j�W��ԧ0�kugVj�A*�,Q�䕵�T֙�v�ht�Ҳ���y��mIOr7����'_]�
���1�E�z��u�(�t�R�����Ef���f�۲	��/mo�`��#��b��]��mFAn��b�:m@0p�N�g��͔�ͭ��W�R���E�m
��V�Bu۵*�n��k����ML�Ռ]�'��(���u�:��\ɺYc&�,ڷz�N���\r:�e #�Q�.�6C�*S�y�k��ü���r��i�ts�B�n3BiUa�1���l�w6��7���{����;U�	w[�'�,���1-��dR�U�h8�#�D�tI饁�O�9���P;T��0rΞ�]Fk�G�D�h�|�;�e<�@B�O�}���tϮ͌�(����Z��O:m��+ i	�ѽ�{t ��z��}��o:喌�;��U��3/`��e8$�Y̞�4(@��]�Q»8�r��e���Zq�mN��rM�Di�����o���+ll
���!c��vFl�^�1��qZ掭����*���Q춺M������Pu�5L�Y@�F����U�v�ܣ�@�l�Z��k{r��s[]J�Ur�Ѷg+���s��Z[�����B�[��Z�A�_]ِj!x��LZ��i��C��y��*E����&�Pj���w-b�In��n�֫E̷W�)U���8�Q�h*��Ea�S� ���͒����>i�}�r��3J��[��M���57�:�a�x�v�K`cv;࠽�j�+"�8s:��.����H4S�K`q�z���Mu�P�v��%���x�b�S:�:��#y�u���q�2�Y�r��8Way����ю�1��]��cL��+oo��X:� �����,(E4���s'����ͤB��Oo5��̪���"J�_e��ރ ��������E���ّ�[���{j�YX;T�Q�y���E�^�TȮ쎴��r�+����`)r��;��ĵ�'{��]k,����kq�ve;�q\y������GE����4ԕ�gm���1:V]�h*f�[avS���:m,
i�^䫸��+�r��d�	���m�c=lT���N�%�f�ΥǱ\�4�q�X���ڰ���:��G��"{��-�S.
aW<�E�Ik�$�o��	��<���5�X���T�B�;�v���kjj�;��RTD�+��u4h�������е�'_G��tՖ;�|^�9��+�9X
�CS��]+��|OV]b4^���]Yb��̂��gnd+�1���yO���T��9.XʺfeJ�r'���Pv��t��Y��Ω�l*u+�=�B���5��UR+2�]�3�X�q����]6���j�j��bm�!���9�Ό�"����`�*�l�ȭev�Mv�D�{�Q��鸝���1�\�2,��0om)�@7)���n�w��l-�ڼ���Y��lF��u���.���SX.|�˲��j�|��u�V��h��<�m;�wԅ���1p����7�P'w	 �N���ϳxj\Y��wtŠJ����17��z�N�l�����í���3��E�Y��8�������1L@xxW�E)T��՜@�J��g~ڴբ[�ʺ+S����ٽ�8A��,I�@wI����/ ��E �$PhD�Iׁa]���V����`��)�Q�}�^5�͜U4������c�xe�<�%o�Ҽ�l��Gr�u�U)�����N
ֱ�+������U򪾧�q�u�/��*����0��Ã����q�]-Pr�l�e�	������pkF�8�v�0�.�8,���pѼa�oy�3Z+o�a-Tܨ�Y�A��5�:�s��c3��rd:�U�{{s�e��S��{U�%=ƥ�vM����C�6�:��"O5.ŝ�(�T��f����gb���8�8����zir@�ʓ��u�v��Y��	��oqp��m˧S��r=�`��ޢ�*:"�3oE�OH�0��t�G�k��##�i�vu={]��IQW���}.\i�_P�*G5n�θ+�'�����ޭ���:�Z��fW>���W*ɘQm��"��Y|v���9sЗ�9�w{�fV'ʩV��P6-u�eu�y3X��`�h�5&zq�[ �dTj����c/B�wE�q �}0�c �i��2�$��k���wayҎ�:��5�F�&��ouc��i�@<H�%�:��=FTzWS�4�Dv:6nwP�sjv��*�+�x��^�
���v⛑����C��B{�q7ĉӹS3Z(�YXa	�%�'����S�� *HR)Z�T�%Q�:l�'�3<��E��K Rf��� �Z�@�
��U:�O�� K�"��N���S.�E���^u�}�g�vZ�vrM��%2���c���d�=AY��Q�u�n`�%f/�\g^��=�===?G�ǌ�?O��1#��5HRP�f�TPd�a�n�M�� 2�`�z��3����zz{x������~<x���y�'�d$Ml%!�T��y��]O�lѰ��f��{q���������~>�����5�Ù��9��+��ԧ^hR�}��Z��)!-��t��uU]f[A���fe[���Q1A�afd�AP@�3�H��b��v
��*#l����*�e�"*$h&h�q����Ȃ"
V�#";���H���"���M��̐�,�w�:�s(J���q��s*2�c:�*�Ic���Ă:̈�n�f ##*)��2���&����)�ʢ�:� �����ܢ�u-�s̌��1��u2(��B�0�*�0 ��L6�-��j,����2h���6�2�0#c3)�(��g���Q��2�r����w<��H!�����Q�F&�lc�VM9U	��[�uu˒���[�F��YVa�n��wJr�L��̞��3LL�wcgc˨M�%�è�0�M��H2�blUw������M���"�;���Ɔ���;�e�dV��f�桱��;-��bu�Ӳd�n9��eY#Ef/���i��p��d6�s����}G<������ju�s)�c(8g	�-�8�+�1C���	K���u�g!�;�+������yz�������م=Yk��1�?�$��̍�k�]�CU���0�%�/>����3۽ ��^�����Q�w����޸���������U�Ou�_7�d�(�vn�w��+�E;�.^(��=�g�_��c�-��&�ɣ���Pv|�{���8'Fӭ��,=���'�򳽾�D��6���ڴ�=髂"U�w.��D�h|�d�E�r��g7�~>�$'�J�y��Y�-5�r��٦�5��v��F�JǕN>֜��&we��pڛ��y�$𮆽�P�`�]C������s�3�����J}U��(�
��㦘���h��׭�k=1��H�8��"sڦ�kb���=�D�]�tw�
�c$�/�D[EZ�f��.�u�y�41���#o���ۺ��~�et��eJ��j�q���V�)c��1گiѦJ�)GF��1Dwg�})�`l��2U��J�gT�n���:3�}Y�:]�ٯu�sJy�E���k6GWq�|Uܕ���ó�Wp�}9�U{�n)@(1Z��6�����L1έ�W����ݖ�;���)��\�ϭ��*.Y�A�!O,[�ٻ���>�\�>�E�ͧ���O��������]�6qĉ݂UK且�2�A�ͥ�^�cj��>4c‘R3���ג	dᶲJ��^��w���M������ƌ�y�i�xP�\��,g�>��7����BB�p�ky����~Rs�\�)��s�xk��P��~���Y����^"`��z2K�kw�]�옹>q�8������5�D؟nLe�No�A[ݙ�گ��MjI ,
���^�'3v�wJ�Tm�����9�?GS��S_K�f��w��jm�=>��y;�����Xچ�&�V��w�x||�޶�*mf�s��m�|\���v����率�6pw�/�X1�G�k䲳��qbrzE��[���'8�5�n޾�=�Z>�1
�7~�} ����y�v���Mq��f����0bn6ؒre�}��~~�Y��$PīZ����2o��\��t�"��r�e΢h�&�JV6J��:�[�g�fEƯ:$"ή�dY.�;�&��ݣ���+��>���nkrg$���޳W�D�P��>����w{:�瓘I:Gc�޸� >db��\�Ϯ.y���=��L��][�{>�/��w�o��5G��u��<ߗ�?"5s���=O�w�M�V��_���_Q�_��S������pb�L
�@�U�[x��#��k*Huu����r9�+�Ww������@�'�l�ǩ�ؾ�d�����������NF�s�3���,H���y��<e�|z�����g�H��n��f����f���vG�ܳ�ެ�ʷ������gw���-�TO�8�_�y�']Y~�[�5Y^��T��7�\�]�NyÓ�хj��s{��Y�;���߆:\s�g�R�M��̻�uoz��!2L�G݂?��C��lӯ�tU����V*�::���r��S�ӏ�e-9��w���ShQ��%��]��*��Fr���D�%J޾ǔs�a����R���m:9Ƅ�q�Ka;K�D�I��Oks�O�����O�`�{�4ĭ�=³����V{ ��ux�M��fd\u���i��t뻠�E]U�֩�O��b�^{scEl7�������ol"���_�����g����!/+>�>/�U|9�Ԟ�rr��ώ[<h�d]� �s�"+%��%�f��4���� ur`�g��(��~�4������/z(����\���������{���y���|z�o�;����z:�9\W��$��|��x�c�I3�}z%��\7֞��#�o�zp{=��؍=��9�9O���9��{�����<�b���T�w�Yރ�8�Ǻ���{@�ϱH��,�Ꜹ| �]��?�v��@T��M�e�����YT�s��U�û��"�}�Ӧ@����:N�i����9#q�� >�~G�u��Ʒ��S�߇}�)���X���������Pxך��ܽL�}(�jA*v?S�6��.�ƌ�y���^9�����Y��[ʷs���/�,]}�j@r굵�V�fݯ'���s�*���	uȺR�̧k2�E�gXYM:��v�+a�\�;볻�)�6Gyo\��q�J�l
�M����H��OQ%��Dcu�e��' �@�����G�0��en�ٵ�_X�o�(�Sge��˺i��]����؀65踓�x�y�٣��" 	d��2)�%�b �EF3\�V^X�%���� ��
�j5�\s?b��Ҟ�{�:=��ڋҟ�����d�]�oҟ��:����΀�(��>:]-���F����秪q��QV9��*��M��_1o�T���4�;��������3��=���E��(@&�t����d<d ����,_g˗����>}o�_h�}��r8~�����X��J<��_tٸj%؂2T�3�X~�ȯ������w�_q��Ku:Jb����y���8�|K����Cj|����|�}[��=�sg\w����KU�,�<��5V)���ӕ}V6wr��t�,��4�f�V>�3�׺�o���Y��Qt|;~"}� B
���&%�7ض�o����u�7�n)�f\nħ�I}+"\�F��#(%֊f4 �Wu�L��y��7�	�7׻���p���|g��v��r�૳�ȵ��v^�����ܺeLC�4��J\�����wSh
:X35��5g=2��ɭ��#�p�2�,
W��U���4\y/f5�n$��f�/;�$�s�3�i0JV���ξ������������-H�w���tWI'sh
��k2#y�'j�|6}���Yj��is[���66�u]��Ԛ:���'�MT��GF�{�7b�y�o �y�I�?*���k�:u	��	�
�{��}�<��*<2a��O�w��I�3�N;9>�!���:/f�lohD��c�dc5�Wji�ӹ���9�Z=�^���Y���d/�w��������6`E���I�@�2.s�"74���̒;M��9}���ĉ��>���w�~�>�5�Ӿ���-��w\Eln
$���BIZ�.�()�*�~g��5a:���t:瑩W�1k��R~�ݔsnldӴI��֘��ԧ�-E�>a��{o~�t���>߼�ܼڜ�G膱��wYo�e���.�K!��u��5��z/d��rBif�"��3Mw�+�v7v�<t2#q\�Z����WûԳ���zjO��)�)�7�����L�.wY�ԛG �q�a}A��uݬ�t�����gRy}��	b�%s��7l���oq=oz����{O�^;kHT��2t�}�����I�&Bm>ط��c�U^b��b�)k������%}���D�����fyvVǷ��9�U��~S��gW:��Q�z���d���]+v�KN׽�iz�m���C�Vy�"��쑷$흝=o���#�+'~5��^*���F���;{����K�	.�i���sx� �����R������+6��j���[7զ�mwf`�'.r�N�Y8|����n�� ���q�ݑ�A���8y��!��Ŀ��'��0Z;N}F"�й��ެ�����9/���ǰ��;�~ʔ��|�e��=̍���.V��4�g"[39��^��v�y$�'[=$(����m�������z_��XUb���扞2
��o�o+��&�L��gɠ�r���{�w�9�k۾��m��<�*I������oq���:���@&�u�x �/�~p,d*�k��W[WaҦ_�{0C�u�ڠ^Wd�]\ZlbU����M�m�|hU�"p���T�H4�kw㤌���	j�cKy�5��;�oU�+D�yfED:�b��r8Ү�\:�>�BB�r�b�g�8!'���a��-�Iu"��k��ȄE��tb��^OkR���2�rf�q��_g*�&n�O<�7�^�T���=�=�E}:� ��fkȜi�������Numn�d�=p.�q�I9�N�B�U�Z<�à�x���\]}bM�V�~9w�CQl6sS+�6oA��
��Z -�'���[�ρ]��|���'wݿz�t�*P��w����zu1�')�T�}`*��*���U4��E��rɄ׻)�|V��k��3EuxJ�g�s��Pڒ��܃2�HӧE����9��w�f#������֯��wk�$�Y�g�6K�
��� �Ou{4k������޾}k~���}5�r���zq��"��2 ����<����|4����L:->0�2_������;��^� ݤ[{���()��}֋nz���ڕd*�6�e�@T�n�z�f%3�������E}�1�����)eV��*!�iXZNn�0�+.lv���w1a��HV��L+�]���2�5/]�ƛ�g��<��(�X�
+^n�|9����R<�d����ڝ1��`�jo�j�=R��,�|�����+�I"#����h`65MSTإD�����Xϔk�QB�(��;[;[#!��ͯ����Œ��h�����K�[���^q�Å���L������&=ݧ�����p�|tPn�iͦt�����x�āV�����c�?o�_�#�Ϯ�|OE�Y;�ځ1$N]���x���[k�i�-|���S#�<�g}�]�n�h������1q����u1�RZ����dP�#��+dT��}�]�s�M��|z���z"�g�ǵ*�=��WS�|)�P�U�{k+����<W��\�y *�N�~᛽���q�Ο�O�g�ԥ�D/�Ů�]����X��o�r����y��Nu��^��7�_�=�%7���b09��`�Nw�|>���mPA+��H�3�V�;{��ugk�Ͻ��eϟ<{m��Z\s���������k=����5:���6�����yɛ�/4�0��,��d�gZ����i�x�9F�6�J�����`�Xpѓ+�*ms�W����g^ʸ�غ^��FW�W�1^A�8�u�Q;Oa���y��O]���7��p�gjy���7R[��]6��H��T���N�Y���}˚v��%?A<3�99���T�x�W9U�}�>d�`�B�.@��y�{{g[z�4�n�@aW&�Y�^U��+�>���c^�r�cI��?�xq)ӷ�<>�3|<P�]զ�v�|V�zj�,����K�M�t=�'m��t���ھ늽��˚�-��k���F?[ϑ/.��*D��v�M���ۉ�p�m�D6Uͬ�nH��|��#%�JaxaÃo�����|˞)�?�\�}Y����T}�zp�w}�W��|��c��|�U�wEm�uw�Q��'�����pBYWؽ>���z{�|��ٗØ�i�R*=���Ne��hB"�P�efRU���,����0J龽y��z,���˷k��׹]OY��u�p���M��=D��I��}��'C[�}^g�ƭ�j�{$#~������N_����@K�|M����)~��e#���J#�5n�T�1�������k{�ԟf���X�nV���t���-��06�c�tR%Nז"���%���ow+WW%��%�H�tG2�9�M`\����6��9X����M;J`�K�w�ښ���+ZO�]�e��O~�b�%F<�F�oG]=����W��Ӹwj1�.ok���ӡy�������o�#�R�� ׷&�H�=��V���
�w�¹��=k��G��VF�m�2���n�)��)�g�)� u��4�J΃��ɺ;p�����lVbn(�fs�N�F[����TZt:�4�2Ȼڂ��$�X�0��٥CD-A���3H(��U����.�Fp�\f�Q����:_)��E����٘�n�c����7�l�c���]\ؾ[��u�q,�_LۃV=�(�n�I�Y/���w5�z�!�hI�=��#/�c����)���i��T��y��y�l6ŏ�u-��mq\W:���Ҵ��%�x�0c7VC����'LZ��H����\ӟE&w	����Ruު������������O��oeZ�YI�o�m]�� <[���������oPW9�/��o��J ���W���� %]IWXvn��x���v"���[��V���ҐTF����tN5�U0,ٌ�t�²���;�����x��&�i��$��0ν���8�;}�u���X�k����z�e�|v�{CN����C�\�.u˻Y���A�3oAbWQ
��XӅ9�/{"-V��t�]�)@��ݶ^m�ulM6�)4�T�b_.��v5@�V���Co�]�As��,PrG����0�v�X�Ƨ3�2��HC��nٹ(��Ae�V��X^�4J����]ۃk���}xh[ܾ�ʑ[�r�
v6�=O;���T<�Q�[B�L��|��%�ᚢ.�_k����$�EDM����Z�r�Gq4��,=�<��{H\�κR�-0�]�[��	*�2���hI�w�^Μ��1q�3�2o�FQ���ɥG%���.��ח�5�,%���헼f��c�듇0@�0�d1v�r�\p��¬Ն�Nv����,꜈�_u�sw�̨&����T׷4A[E��6�a�v۳�v���h53Vo:�©Az��Kj[т�*7[��K.��� ��Wz�q��M�|��S�>.|c�\�����9�N��e1�,a�E��X�8�dğEխ�y��{k���D*��Y�Ej�X{��ޓ;����RH��zр^G����+�z�U�Q�t�U��U�%��v�B�v���Z��qt�Z�>�8�3�˽b6^�� uM��`jQ���
�o�߽�߽��%E-)�SA��)��dU��I�����	����de�v�u��Ƿ�׷����������Ñ���22(l�)��ɳ�7�4�v�����+;ݓ�2è�#$�,�ZhȮ��^�||}{{zzz}^>��<�ry�&FFK�4eEY6a�VC�fKC;Q�����_�zq����������>�}q�~�`���>˶�Y5FCvᱰdP�%2vs/Mr����*�����ѽb�P���NIffaGvn.CM��d��Yd�R�le�ٮ�$��i�����nu��F�d1Sw�YVBS�@w�lFBPc���``�@P�e	Y&E.HUfde�C�S��le���[Yed��`dd��w[�t��2"���1�(��,
�]�����w�{��(�3�6ZM���2���r湥d�%9!^�lً��aY? Ȩ�
�n4?c��;�d�2�6ss*\��'c3 ɦ��2\ �5@W�yc������r�^`���7�J�e�n�92{ =ݗ�����ݠv��:h�����,�!:j=f~����u�����z������`[cW�c��1�a�����D�����!����&��3O1U����V�-��l��
�h�MuS��@H�5Cm�m�q,JSeù�t��ן6�TԵ���w��)-<��&3����Ƞ����2e���tZ���p75�f��5�:���M�e����$=��*P�>F���S 8il�xod����Ԃ�`|@{��.g�B�^�BɄkh�������7 <`�+���f�1�ҙ�T$�2�8[�������5/K�Ɗc�h쭦��\�5�8�@�X|�5P8xv[��P�w5��:f@�{I���(�n1n��,�|2�FӋ���5��](� ���U��q�ό�*�>���p3���W7��@���*4o=2�z����b�[��Q�=��FM��fZl���d��g[�}J8�tI��OI���^�啌5����X�Y��e��qި^m
��?[��a'�m�*_	g��/z�KP�����Ǆ�~�S���Yg���O��ʌ��c�P��9 �u��	d
��V�gèBl��ؠJc�sjo�Kn�j���<M����K��#Z"$�PF;����^���Of�}Y�z�k�)�����ډ�fU�w�%�(�V]�Ǿ"��#~�u���Yʹ�{XC����+�r���d9�滽��Ԝ�� �3����)�A��]�;5�O�5W��� Ee��N�ۡ���<�[�q�ܳ^��q�Z@2b����X���:s�9���ڧ�A�x'ʴ����*���t�)��Btӗ;���M�И�/�$Qs�_�Z�p�׈�֝_3�1I�bQ3����F�ऄڀ�Ft	�v�|*=6�Y\��V������kC�	��O��4m��|�u:5�*��}�:|��{�/���	<!�Á-q��&�I}������j�����P�6��Y��nW�`����ێ��I�*!{Ⱥ�|,����ĶB�8�P�cXO�>k�3e�!u�U\��^�j�P�hx
��5:@U�L�\��(������4����ŅkI��Բ��Ï�m��a������A����0�����͝)�� �0i����vv��^j�P[��X7�q�u�;Y�n��p��Y�p�I�#�����(��)v!�|�=�)�����	 '�C��:�Pĵ3���:3�Ax[	Hڷ �����c�|����&22|��f1R)�v�9l����Zc��y1ot!\!�S��Hx��Q+�mF�G+��p"�gE�0/��)=[,��.�K�q�ư�^|8��ҿG����(ܝ,?���(�|��`*�>���J�8<�d5�!�kc�4���*���lԠ���=�X�ޔ޴x��]���u\=�Ō=�J3� �*�L�������x�\��اlσ̃m3+c#m�l�q�Hds����f�dV1�Q�x��\
�C�����O�� [��N3�8��ֺ�������qB���px��nni\�u�x������w2=pX	2H./i��.>�	S��G�(����|�3����W��M�E�.OR�����/zX/T�� �ۗ�v#�\xZ���\
^�y�����A�8���3��)���r:;}Ť�[56���d%���>y�,�XŪ�߱mxu]'���0N�m��\�֢B�T@n@DĨ�@��9�,�ٶk{��w`���۶���oA��Ac���n�!���1���%ԁ,���$.4��FA�~j bЀ���ȳ�*���
mW0H�e������
<1i"(���rq��_i�gh��I����T�k�P��su�r�	����������r�Y�N�Hq\%��P���/�L=uN܌�{�jt��2�	a�^O��/V����������ENk��Z'[�#>�#K�5U7}(g�����H7��i+�@s�&oh�7�bE�W��5�/������ԃ^����;x�׼��<�s\1��O���!ѻ��dm2����ڵG��6C�R{H���S$M-�����3�J�|�l�{�V!o
�������VyBz�ױUݚta|���]��FҥC.���P,Ԅ|�y���WJr���]	��>�Wq��fVu�N8w�w
c��U�s���uۺ��&_3��<w�a�`|��s���==9�=����مr���/T��E���{Z�@W�K ��G�a��J�."y�a��c(�;@p"] ����5����1��Z�j�48���A�5���M�	�"���0.cZ�{����g�~׳� �F&[<@薨��R�k�g��i�@v��48���<��$n]���?����^꣑(��Ǚ�$�`(0y���0�CA���wE0�Ѡ�	� �W�c�T|���v�f.��Su��m����ץ�	Q^���vĐ%�s/��-�:��s`M�Q��99����e���&[H	�U�a�O�O�<"�C2�|��=&|�.n '���Dkɘ۱O�{a�b�x^��B3��zu����,v�� �)��	7�/'ùD�L�XE5>�-tE�3+��]r���M���=�2|Nݰ�+1�`W>T����*��+\V�iNC�Rqa��g������	j�DbP�&��ntQ�^�� �e�Mİ�Ә�=�?2���@@���,�+�n mkt�-�"��)@(K�dw#��w���@�����b �r}f�:��^C��Έ��	����u��ϑ�vvگ��&�y����`:��(V�i�!���단�3%o1���;�6��Y}.Y%��݈� �0nw�YȠ��<ia"��+^�]��o��ʷ(=�V�rPyG������FgAڋ]dZ���O���N�����kPh5u3�ok*�__�__����ёhn��gRd��x6��u����;�s^d(�����B�'����	���;��B��"�8N�.<��Lb%��Ӂ�Tz������W���p�٪ t���Зy5�!��ʸZ���N�@V?4y�(,�M����=�Q��.��|��p��d�0Pu�W�B_��9�
���y�L\{���߭�eq�ϱ�)�����M*H�`0�}�i�˗P���Y�f��,�;b�1��X�=5�V������(VϨ������J=�AO��6�bNړ�$��np���[������Q�� Ud�f_�X��M��mU�a�����C�<�><�J,�%\e��_>��V.��Qp�h�ű���Nuw�{N
�v9��Q���i_S�����wJ�
��w��x;"|$��P�!�mU��%s����@EX�|`�[�	���h>��J�Mu�,,���-m��3h[�O�o?(;�H�z#�Bf�V7�)V��*,��DK�8�,�������ޑ��i*nph����[��?�Rc��wݐ�$W\
���zI��^83�w�Ny������nd�{�O���YPE��y��-���MB7��	L�~�t���'kWs6�Gi� �_u���J1�P�Y.���;a�kjW��$�v��	N�pek�K��{^��U�5����Z��⑹��޳�1����v����J�^���G�?��T^vLB��;�s���GW�<z����)�C�ؤ�x�Se ��=���y����-�1��d�#8���P4z���%o24�C`.'Z�����*�ɟP���P��ڮ�X8潘a����x��3�Vv֗��C��oC�j#��i<�尘��~�֧��Y���n�\k�����N�P��(tuL0;�da�5�NO�sة!�1I��f�/;�U)��nCދ�ڥ-y��U��+�v�������DZH�OK���P����	Ք���oIm��Mv��׊Ut�o!hsñ��u�Tq�B;_Oi��'�@�RH�T	�D.W��x@�/*a4�꭬h��]D����8���&���\����u�~�����A=)-�|
�|V��/��A��<TB����R�Nׯ���y@��j��~h���|L[9~ͺ>��������� �$��UZE�]���Y��qv�k
���2�D���57�1ש5h������bo%}	��X"����8�&N]������%ݧ�Da�ں�V�Ų�z+��}!ߧH�Y����Į��D�U��/�݆�H�W[����R�ce1c�Lȇ>ق��`��PU���N��'E���_.��W(u6qL&���p��=�wN����D�-�;����ٮ�P�@0�I��ʙJ&�T��8h H-���xU
��U�ܗ$�n�H�r��]�ջ�	E�]����:��U�����&��C���Nr�	�A�|z��oUݵdn7A^J�Z���O�'z�yK�t�DǙahd���KytE��-)LM���2/�<�����d�ٟo�/]1����x6�0c7���q��q�����o\�]z9�o1�]y�'&1ϸJQ0Ýl'P�C�(R��1���KѸLi,�Y�q�����07,��G;�#�kf>=^���/��X�]1~��R�e�����t�h��ח�r�����`G�fsW���0��uC�L�d��%�g!|��XzT��03zU&� '1��k��T�AY����g�W���z3(W�79/m�6zP.��sц���l4�7�Gwd�/�[[��T��-u*\U�94Ž��Ν���.Ջ�a+˃�z��K��&�O6�����2� $���*��}��W��T���qR�B���JV�u���^nc��2$�Nj�������}��L���}��MЮ~.8�=�~����a<�@�1�^NE!��
t�|�5����53g&���R��1Lk|Qxb�vf果��Z�`ͫ�٬�B�4�K��1�X��K��A����]���؃� n)۷�e�2�'����Pr|fl�[�U��>.�wV��[;c��NHX���ʠ����S�����i�y�k�1�aw�Ȇ���{f��P��A�N�B1��͹
K{��U�6_"�܌]m�Or&��1,9\A-�~�R���Ny�'�؊�t8ξG
�F��.�"{[zy^Y~�jo�f����+dpN�	�q���@x<]�����t3z��JD��R�p��k^�����f�vC�%�1�7����e��� =�jby[�)稸�[T]��v�˰ZԆ�Ƒl�w��ؘW-��{��ﵡ�)��2��<5�\��jzd���1f�<泀��j�R4���#T�������!��H;�r�c����e��[�9lna]Gx�Y�c
�f�,K�n��e!A��	o6�X���#�ڄI��ާ�uu4{Y�Dp��
g�܉v�.�ȗ�i��rQ'����M�1NS��v����+6�F�B�:��ZC�o"g�'b���1?�]�=o��)�N���n�#lm��=g�,&�a�I��@#���į�ܕ�
���}��{���S(�&L�z�ÏwG-�����VWk�?��2�I7�l���#�n�(� �dH�f��W+�	��7t�l�}Hk�6D�ihO�'�7[3��`_��P]�q�*{`��-�J>��Ǔ�y����h����Y�_9�0F�n�y�W���U6��G���$�}D�n�7
�!2m�oL��2�_��6�k&�HJ/�^C��	��{.)S�WQq�|yN{��HA�Z� ��0�Տ
5V��`{�R�o3�Η�P7M:�G;dY]lr�]]����V�-ȅ�a��Ych=uJ΁o�M���N���Ϲ�}������R��˞���a ����k�P��כxc4����*���]��Zn�R��K�q��.i���t�h�=�W���@������M%�o\lk�R%�ls\&1��2oc�!T��N�tT�Q��l`S|��\�����44D0ˁ���N[�n���/m�����jvļ+e�FS�25����i�	�;��g!�Y9LnokF��5]���虼�m\�w(�^��(��3Ԕ�n{>~~�5�󣓤��t`��ԍ&	T����l���ԣ�7؏A{l '��iQ��cb�c&¸�1`�4�V�a���S=�\�,�|�y��v�&8��n���wc]"h�̯nّ����.��蹫A�_��'ON �1�@(��p��j���S�����;Á�儽�.J#  �\Wh��C���Y�1}&�Vj�_eP����]��Ŋ��E*�x�H�Au��g�q�!jB j��M����N��.#��ojK�c�k��⾺�G����|	�:/{+�7���#��v�SF'J�1�S%>�.[�e'9�韺񼿀ȧy��O�r�
�4�H�Ś:�.�c�(�A`�۳�b&������E�j=3�aݗ�aT-�Lk"�gWv�������PU�M��-M��M�޿<��P�~֔�xB�U�Rܐ����=�h�rԭl�!?~4٣���B-���u,���s�g����/@�oI1|@�0S+=VИ�t����k/�Is|�v��U�Ɓw�AXgV�Ι7������~��%��%U�veV4�Dfg�*�׻�B�ka�)������kQ9f!�����7ٮ�'��չN�3�����2J�%�v��ʒ·_ε�+�l%�r7tP=ѬC��c���V�BW�4si[�������5O,Ķ�DD�ϙ�ֽ:�l��1��3B�J��`W?�M�E���^S	:�g�<������m���P��bH�B�.��1@u�v�#��u.#^�| �˺�R�Q��J�>A�yj��!��y@���[D[y��A��pH� �ਃ�7���<���2Έ�?�*xj�=JK���ƥ��֔��*T�cI�yu�o�	Y�U)ns��S�(��I�Ҵi9P�e���#!��!F���W�:��/6kK��JpE�V���K�p��/OӗƎ�ù$��m���6��z�o�M5!�2��8**m��Pv�oy�s���fﺏ2��a�A�Ūꡍ�E.'%��[�J��a����n�UgPG(<J��R��r�d��j\6'I�'Iq.l?]��'S!ڼT�vlۃ��f�ioSw�I��j�}L�x�������45���=��ݗ4�
f)���h�r�WA��z���げU���=�|�B����s�눃�-ܸ�u3�h,��*�S\r���U�+�\&�Zћ�H��+\��>7����� ��b�Xq"E��of�6:��9.�-+�l�·u0�;���s5jT���ج��֧;�P����a"����e�����L����#[���)X��h�eֱ�`�ɱ�7,�U�����cT�5�K}|x��y��,�CU�3WT2�R0�GO��:+v�Ck�:wƊ���-7)�+�\�/0�>��^c��}�]a�˓��WK.;��2��(���C&tL�+V����l.uƕ���a-	�eI/[�y�ro�{N$��S�㊞��l�����Cɋ�A�i)����e��N�v�*Ƌ�L֥5-{��:�=
آf��z{b�
9�7�E�K���K��4E_\�8Z�t+y�o'3֫�%�Z��`?
e��	R;�ũ��y�r
hK{�^ +��n�}և�nZAO�/��Z��6�^��\x_wč\�eڃ�6򺬴M��P��+����Ǫ�s�ǌ��Z���0P�B�<��Nb ���ז*i���w��*�.�j�Xd(l��'�nM0�롵���S.�[�z��P��P�k�rˢ������:`�ܻjb��֭�%�1K*���v���o߆]���I��(��j���Xh���r%�c�L���թ@��wj�}͛�<�:���Ňz�m���3�{I�df ��VR��k�b���7�:�s�>{Νe�(��V�Gۙ���L�;p�ЭRi����ij�<Tg����6T�5Xϐ[N���Cy�^]�]�K�Q���q̶�2D�J=ٻ�'��zHN§�M���h��ָnJ�(d]�z���T��G��u��ن��z@+ ���MW5��޺�v�Ӿ�a]�� <�]�}h�����n�߇(�#���X"P��(��umM���v���Q�]�K;B��8����$�b��w��҇a��Me�F�N�!��jb�ƴ)�po�|���+8�g���W�V��ogrL�R���Ww3F%P�����'�%�T���J~����b��j<d;KK��'�f����
�s9�k:�e7����YK�N�3�+��{2�����(5	J��B��S��6���!��*R�@:T�p8�����y B��E2RE[B�0�m
.�g���n��2q_g0�"�2�6���b]a��&MINI�dx�{u���׏���Ƿ���������`m�l������d9Y�[wuRUm��MΕg��:������������}}}q�>�,�}δz�#$2W$������h�3����i={uק�___����oo����q��)���$��2� i���[�y�u)F�d4�Q&Y?%�L���R��r����0r3
�	�a��0޶�jM��Ǭ�Ȣ�ɾgr@uCI�ReE.Gv��d�P�MS�FH4��6XylR7x�m��Fn�Ԧ�!Mdm��S�dgX? ����.�7s3��,�J3$��ri2�*(�66+p�+&�b"9oY�m�A�QEpe[d�0y�G�:ӝ�uэ���nƨ���]E��r�)n{W{�|0�՝,�&��U�Q������f��X��V�5�ӝ��u�O��]mloGV���X]w����[���)�2��-
��^��;���>t_���E=�������τ\N>�տ�7_��2�`�V�]�O$��ѫ�;��0��<��u>;��-G'l���H�u�u�܁Fw*��q��rB�˩u:��k��*D-�L��y#5�]+"[ݯ]��^�Ű�aL��5��z;���/�{�Б�1z遴�s�8b�@4��ǜK򓐣׵&u4[�{�=� s-��j�)�;�����l5�kI\��zP�*��g�sQ
T��:�Z-��52�kqJg9����J�e�'�6��ͅO������̼o��cXV�Y�E���m�Wq9�����)	12���5d"�mǙE�?��`��Y�).愆xs���17"i�rR;r��0��*�T���a!�:B��r�R&�A�F���>4D���(�ԍ������Уݵ� �7d`I�J���F[�M�P6����uW%c)��n0�UZ㶶��d��9��N�tqd4��SHZ�l�!2*����#�-'�
H�Y�q�dJ�b�6:D=��9G
���7�"�D���k�>�4��a�q�*�7Hk�ɷ�8�ks2�ӤC5V�v[��ݹ��5��|p7��
���N�ʝV�]�IG����3�=�2�;ܸ�{��~�mr�����O|������y�9�^n��m~����%`��2�H5! ҋH��f�f�S����v�ج^=yfe7�t4��T���X0�碏r�`)ƃ1:^a��G5>�^6�kA���K��E���]���O!�杰�tLu�k����h�{ew3T�����r��[!�Oz�
&�ی�|k%1��[HP��+,U'Ĩ�f�/�z�v�\n�]>p�!�B`&%�zёe���6��$`��O0�QQ��Ǥɹ��m�f�6�wSb"V���b��NL7�xț�<_�]/���A/��M}3A�^)ļ�산�vdM !���Rk�ڤ<>M�y=i=�j|>�������?~���(�sO����A�0��a���fC���PV��9��Y9�m� g֫,S��3d����J���,�����Y<AN(�&�Fy�^�T����	�Hjk�mZ�I�M$\*x�z�;s�t��h8s��,�/$Ք+U�Nn�i�hr�Ŧ*���؊<��������uy�|��n���������5K9Y��NH�q!��Nx�f�m���N�G�C@ˁ�}��7^��gf��(��;�t�jWWbm��z���,(WLj��n���  �LWA���ѱ��7<���v��	muD;�k���"������$Ot^P���?�e>���c�+M>�|�86��]�{61C�)z�����9���#��x�y<}�x#�� �����疯�1�6�B;����q5�1L�JA*���!���l&_F&���$H-۳�ko�GQ�Lj�z�JAu��!���	�ӕ�
���Άq�v�#Cq��%��{���Yt��c�-�ڻ��XB�U�DͿx�Pt�oʪ����P_ƾʨ�~����2.j%AKi��?@��: SO	�L���oUH��uC2q(���L�J��T��S���Kw�^?c�-�l�[3�W�JU�㜧P������zm*�M�����V0�
m��E���g����.�]6e�#��	Ƚ�r}7�BF�%˼L4YN.�t���M5}כ��UKM��`��~��MDhs�
�������n%���oa	o��l՚��Ϸ��仛���4�_׆C?m�<����@��(3�X���b���*9�������*�9��#ZLJ����-ݎ���}���{nm�$F���&�@w�L6��;4��I �W8�y��j�K e����,c��C���v5�vA�T�����X,9��x��PX����D:5��x}�.oԞ���_w�6ݼ�н��Ca�>F����;T�:�z�qP�W��2��V_ؘ�:ܛ���gL���,�#�6���ӵ#a��*:z9B������dv�k�>J�i�nkf��'+��(��]V;߿~�����d���}��O�)�����P��ۆx�Fj�O�'u��dg�8fM��^v�(���ˬ�S���+�a�QJ5;[�N6rd�I�AN;���@�k��lnDtN&'{@!�������A*�tR�9��s}j�D
=�³��Sc6�q~='�f������"��m�����n�X��dga14ǘ"�[��1�ʖ���
�� �66S�P,�j�.��V{L�����y��,U�Ҳ�&4�N&-ˌ����oa�Hb�f�u=�\a��
��N�.��L�;�X)�\�>�1��p�=�R��Ǌ��O���\��֣�E��T2���F(J�#T1xF1}ĵ�v�[�O=tFu���&E-��G2�WRX��Vr�}�ΆT'��n�BZ�D�m[�=�K[��hI��9�:j四J7�ۘ�yz�)cn�k�.9�Xdd���^7�=m�|+�A��z��1�o�]�5��d�3���r�#����5I�M<踕����Q\وbh�G2�\o"��� �f�ge;f���K	ը�ΰR�+=�W23\s�/	�;6(mT�]�E�-M -�t�7���qKWT��{��4| VU���$u[��Z�����O:�N�2U�sլ���t�)����Z�6wi�H%wZŲ�n�`�c�X
���Q�64�y��X哽u���u���B�����!�\��P���y�:,�ݞ�p��"!�<[�oන�̚�m;Z�^j��C�s�ֱ�q-��0&"�T�����C�j����K�n9b&1_u)ܬ��R��gt�h��P��δ/+|���U3s�+94��ט�;/.2$R����\tkbG(l8�LQ_˩��+�:pK��|z�S���5RR'��U��j̍�۔ɯ�,��X��[RH���L�B.8�!�����\̃��=9�R򜗿S�@�3Z��Ʋ�nտ�����S�=E� �7&a�zݍ_"j��j�q��9<i����h�rv�q����^Yx�[���[�T��,��7o����M��ow�����A��"i��H��p�1�VB�l�@[���X5���1�p�ԗ�vcY�g�y;����S��%c�kL0E��ӊ.<�X��yv�u�%�1 ~Ԟf��CWpMi�4�����dbi�����}�)�kQ\�ߙ�d<h�ߨM
SL7S�x�no�ȱ���1�[�(xv/�Ku�ci4��4����H05�R��⹜P��[#!���<Y��� �U0���2!���5k,xZ}�K=y�ǣ(q���
�<u���Jmu�&!z�ȑ�.9,[�v��gT�7w^�5�f��yoy���"U:��\�#��nj�;����'��z����)\D�D�ia�3{�  ��(1�x����ǯKո��q�_K�
��0��x�����Qy�3ƻ6�wR(�d��h��2*�jt�C:<%D_x�c/���-B��rC�9	�������ٕ��������������N̜e˱hRV.K�X�,�ޖ�����X�sM?��*�~ӷ,��I�q>)�L�����7�]��ŕ�jȀ+Я���u��u��������~xޡ�b�nLl��!3���yoZ�V�ʪ�@Η�Ri �58~��\��n�6�M�G�V�c�
�������3�0�)�Ŭ�;���;R._^Z�t�>%����TU�3I��f�L�fnE���2/[�)�ڲC��)��R[�ኔ��g�Ͷ��qB�$J���̓�����"M�C�J}S�®��Z�f�w��XH�dp��?�#�ےb*y�q9�[���5�p�Y,5���փû�~ʏdF�V���v]=mZ�P�n��D�w�/�(L�a��b�%xPqa�\ש�_&,z�S��>&��~�����L��iR��啪=޴N��7n��x�,�=<q���^T��c_w�}���{P�; n��W>��j�c�7/:pդ�y]-X��#⫃���7)h�t��^���w�Mo����̞�c�9	�/kj%�1f.�?dC�!B��G!(T�0aS%\r@F��Ϟo����Yz��.�|��zԆ�25���r�]�^?�,�\'ۏ��
���l����疚�Ɨ[���
����#ٯ��@�w�!���ޤM�]�'a�fSUTqȴQ-z�yE���L'�h�U}8_����l�L/U�M{6cL���	׆|s4v�W�>���F�_��������=6�F��J���Xi9m�"G��27{Ӣ&T뚜��ͮ�ΧrUC��_vR��g6%q���Q}�㎋���0��}ĎƠr���F��TyY�w#6��=�#\S[��{��}d�ay���n��L6������NW_й�# ��r�w��c�~�]2>��I���%��y08��]"N_�d\eL���}�E�y�{��Ĳ�2��,�e��k{k�fX����{y���H�4o�PWf�{����ɧ����P2|�Gdw3�8̦[�U0��^����OW3ל�i�c�];�$�M[^��Anc�hL�^��11�o�Z����.�X*�6�%V�C��qӜ6{����`�Qm�s�`�{�����W6�ۮ��_U�Ki:���Ճ� œ�ʔ�݋c�q�u:ʥ@¶���jR k�ur<^��M����8�s/8�굹㜲�
g4b��.���	P�bʻ��v��Ͽ|?J��U!��Q�F�ZB@� �����ι��!|�KG�c�-��L��z�K��^�E'�Uf�7�5U�=�K��SR&{��@��.����6�Jc���}Y��Č5ٲ�Bq֭:�x�z��y&�}Es��;�
�ܠ��7Y$ZZ���t�B.7���MB׌
3�&��g=dá-��\0�1��c<�Z#*3]��cm	���u8p�٨��e��[S��Sxkt�Eu�����v���ǒ����m�a�O�^�k���#�2�+�	��[Q��i�NF��X�:�\���j�?]��r�;]�'���S��e��D�\u�N8�+��U�2���Z�E (�s�m��0��T{wUˆ�S�Wd�Ѫ[)^�QM�zf hU��6[e�����Dָ��5�T��W[qR��(/��]��Sr�q�P�\g1��eʅ 42b�1�Ng��2GtxCCYܑ~��2�9W��f�,����2r93 5nӵ��p~�&Y�����FˮN1\��!��HB�彼���Q��DeI����[���1/��}��|^}�@�|lf�4�%}_	�a�l@"�i��I��FPa��&��h��(i*�Wt���k���|�"M�Zu8s�7Ob��iɎ�i�l�/nЊ��]��;��8�Q�N��m�V]n�ٝgFgV���2"l	N�� � ���H x�	����9-2��7��zFD�C���S�����ZLx����1����M���	�_T"�/�Ι��:S�*�����ԣ4^Z��4v��"�� v�z�%
�=~Ǆ��d�`%�M�VШ�[�LZ󔰫�4�UB�S͝&�֮~}7 �� �/	s-2Gd��D�=oBeε�>p�J�nMw�{�@ݱh��6�U/��Y0�w�m��G��;+%���y���P��k�%�2�c�Oԟ�-���u�e��ꘒ(濡���d����Q�p�c��M�|���{�5[�a��'�|T��e�w�Ӳ�h�9q	���	P�Թ�\(vF�C
1��;�xI�-�</Z� ���軘�]Ul���1�r��jYo���M]N0Q�5͐��.o�'����~d��f��]�W�)�$`���}�Sf�;�<l��TZ�����[uO7}&������xl�M����ϱ�T57�"�F�IG�x�s�
�Ln��S�.�E7IS5��}X���ec�j%�y��+yq��eh��5답�����H'8���b!ee�F���BY�G[CƲe��2"U!(�Y��8�c4�K�*i�y��5�䩕�[�q^��.m I�(DSh��O�3�c���Y��'׆ڣ��Q��_g�a�}�:'�(�7���߮S����b��"^Z������ {������� !��@����LW��֝A��Z�\
g�(�j �e��6�N�Ms�вķ����j�ۓX�[���]��^�*q���٭�T{]�P��!�b&���´y`55b`x�~T�u���H�7��.x�-�y)�nڡ��i�`Xc�V�5�E�'��^�1�a^�,ݻ3���Zܚ�V�Z�r;��fuH���C#Q-����u爂�%]�LۺoW��ڢH�Y�3 �m�L��M>P]>T��\�%��SD�ȧ0�Si�Q���ns�3��%L^�7b��P�*�9W��C>�C��R��7��7�!)�aN�+��UZ2}��6;+J�s�վLOJ{ǘ$�/<6;:,������H�c�UmzV3Ǒ��l�>�>;*��.�Ӫ���3}�'���*�y��6��vF�ytT�3殩b"����d��>���@F�g�zv,8x��5^?��N�7�%����\}�e'XT�0EmP�}���9\�nA�F�ಲ�~�i����Q�6󌩝b���'3�	q�h���S�ocqJ}����߶���\8j|�xx���oG;����F5ATCH��P��^�������w9����&���;Ss��^�K.�ˑ���%�P�:�%��E/*�5Xe��>\�*j䮥E���eѨ�곡ԾR�s*�^�`pm�ڗ}5�jɅ��\1
���Q#.w�@�������,;�$�ͼ��n��o%5�z����WM�l�Rܝ�5Fl�K�/+��'��V�; �f�w��	I�Zʾ��l!i�O��o14�&��gY^��+��%aZͨ��V��*��=�͂���JɅ����Ѱ뱌j<���ir��8����#zpf��6��y0��+�à�ٛ�ƕ\��8r��9y5P�hW]o�t��#�5�rMGK�Y�AS�U��hJŲع)/�ЮݘQz�����f����v�޶�/Zɘ%<h]�G:;�x��8PoY��y[*�L��><��:�Q��,J�N�̈́�E�F٪n�G}bSz����tr��H�T)�����joe�Ӭ�fl�|DD��*��Vs�F�WZ6��L%[������Y�.�YK^�,]e�Z�yV�I�hm�������n*���Y̳�<|��r�s]�CW���4ö�ы�55��ea���[X�.�&�[Y�U�Y� �V�c_[W�"B��V�I�BW���5^2kf�)�اE���O�-m�����dy[nĔ�a��Zڷʮ�JYZ�	O����F�sۡ2�c(�ғ��M��n�NWTJ�u6�wmv�K��Xv�RŊ�K�`x���KC������cGe�E�ۓ��h�tR��)(Vj��4�jf�&b�}�G�E�f�G���&�l�4��a���gh�86\��b�lt�0<��P΂�[Y�-7��R�����|~�Ntre��{�3��֯���+p(���dA��Ұ�&�wr� P/���2	W�oQz/;�B�]�˻������i*�B�S
�;��s$_<r�[��x��@�Ǖ!O
.��6ꃖw;�(q����[|�Z�g*h뾨���̺ܶ���i���g[����*�nIL$-<��Kz� 2�b�ф���#��]٠Y9��\i>U��2<%�+�6�W�ifU���8jGb�Z�,��Cb3Qd�x��N��}Fs�7�yhU?&�4ڕ=-k&��%���$�"�JC�;�[�ZN�;Z���*�U"��=��b6��ORC���q�� �
�s��������g]�,f�\w7�:����}�� ��[���z�d�� � ]JK8O�k��뼽�F�5���t�5��yJ��sQ�b3��{x�_�l�UB��A�6v���
����!�ȉ.�ʫ<��޳Ƿ�^��=>���_\q��X�]�#��20i22��r,2��6�Y�ק�ק׷����������{�R��J���"�aY���9��feU��>���������������}}g�{G2����r��(<�z�����������<�qH�rȷt3r�9uY�6Q�9�VI�QRRnnf�E�;Run�A�6�PLic�d��Y`Yfa���B�NE�i�����GDF�e�Yd��D�4��C�N�A�aHlf8YcILU��fd�Q��[�DY�-�n`[���dDQ��UPf�n瑳�UT�3f{�HD5f5U��e���\3(٥���ǐ�#T�o�9�m۔N�}wb��j��ᩅ+�]��Q��Π�H��s4��(�瘸<$lWk����*Pw�����|?dD?C*���
��A�TiR�@�`I����{�r7rj������=/�>t�)i`'u��$���#�I�]���a���*o:���p��w���w�*Qf=�Ɖ�2d2�ɰ�{��O����/���S�(�y����vd�K���yjd�f�Ƶ�ԁ&�5�p���O��$�b���F�V���,��l}n���؍�u��P���'D4��b'!�!��"�����PʹP���EUZ��U��xِD�]g/)�](^)�t	9mf���
�N�0�6ǔ>�J�Q-·����?Ni2��|��88]zkkwL�U�kS�{��b�1�>A��L �ޠT}z��"B6%۫���ԉ�
36�;&�O�T�c��r1�����d<�ޕ�<�\f:(��aZ�۬(���ja�S��L���u�<槛�+Upޖ�n���_0���P)A�� �z���X�o40�A��:Y���T�E�n�璩[%j�Li�*}"�.Ӽ��USQa���9���u�ͺ�2e�v���k�Nua�mȹ�H'ݘD8�dkc�0i�\`��O8cΆq廧��4kJj�({q�3ئ�>��!��-}q��B�[����8��C��{�Z�� ����Wfr��u��y*��!��=R8���,��)3<�zފ���1���l�w�q�[;j�L˭e�|pb�Ӵ՝�2�gϥ���Va�D��T)R�Q�������o~~u����Ʋ�@��r�ۇ�������'�	I&L�Y�&0���-�7���l/7�m�+_�O{_�Z�x3|��,�h=S�}p;��Mt�2�C#ء*�WN��9߿w�]a��&���v��[��	T�r{���eV�/0���iz�nT˟�^���)x�mcC?>�rqyi��7��*�t=9�_�Q���<�{�K�L&�Ji��Rx�d�e�ŕ��Nw��M:��o�L��kG����y���X�?�����f��HQ�i�l�T��۠o�ڣ�6^0�݂��r���@맏����E�1�)O7��tLk)���u�3���oOR����u�ar�w5�)��+^ ��5��%���5�[,޷]�5b��V���#5榡��^��]Fz���v&��qV��+�	��v �>_0g?���3�;�U.������e�93>���r)��m?�s�ݟ=���%q�J�b��MU��o� �Ry�)�w5z���ð�ig#����R�`�����1����n|Ԅ�Hw#ȵ3\�&�_��A�������ڳN���}������m�����5�T��h�Ћ��]vn�ie��LZ�Q��*��_�����2���qȣ��#t��Y7.٧�L�kW-Oh5�w�����$�m�r��k霋��9fh�n&�&�U�[�{���>�_�F�DL�0eD2T%����| ��tz..c^��;��,g�R~�#H�hr�%�^��`+TxR���.��h�Y�Q��_�V�3�k������� [4��8�dkJ&����
��S�p�۱�Dh��[�4���֭�O�(7l�n�H�!)�îQ����ǒsN
�L[�gi9�5�4ƔBm�;�H62OM����H6�f�#o�7����P�@�Nc�հZ���{���(�uF!�I^�J~�P�ފ��2�6��GTW��8�P;��@̧D?^�'h�Sj�ʆ��r�Ţ�.�/kYU#�F�0���\WR�����n%�`�ľhJ�T���r�1�����a�U����cÐ=LL��������jz��c��~� b�أ�������d\��j%��7sv�kG�1�M?� @�j:���_�A�m���h,��C��̽���͜V�;��lك�i�|�{T&�gU��6�Yz�^=le��T��&�ޏ@CX��ZK^���(���L��nC2���i�9�e4'y/����c�[p15�y^Z�
i��/Шx^�%=�h*�/��[��Y�.�Eʚ}�U���İ�8��Z���� \����!<B�y߽Z���jf#;�u 4 �{�{j����K�&q;*+ז�w
����x��`���ֶi5)֢�:qT0pC��>�����z�?C����"d�-P�)@�J=|߿}���?3~?&8^;���ض���ݬ�Y�	�P�]�cJ��J���b�Zb뽋���/ڏ��9��S�s��8�m���&��z�"��B)�n�cͶ�G1�&n�7" 	�H"��-�>����ڪ��ָ��|"���k=�^ ��\7�ɞ���wq�Kz,#Iy���^T���Vt6��V��`}T٨L���4�r�k��[Q�k%�dx�a�P�$6�4��ԡ@j��u,�o$Tk�v�K	5&��g� �wJ�oH���x�5@f�������\��S�-긾}�w:�i���eF��	�&h�pS0~���]����z'׍:�u�����c��%�G�:WИg�֞�45V
3'��BrK�5.w/�V�O���r�PΤ�Khi'z$5�Z��!D��eU��X"#>+����O	�WN�� �%	1��;�QKN�q��G��9�5Z����,����$q�����
��~���8���w\D3NK���TM6�̕�Ok	V݊fT�P��,�X�U�"ڕ9L6���%cIq�y^��L���{�+�W�Aѽ��;����2�cd���I,6u-��P��x��3uHg9����v�t�Wl��Y���7M�y�Г[35�aV+y��,J�l:��Y��%��wWrq� ���A�	�0d)B���JP���4���- (~z6n2e$SWٌv��t�	i�u�z,�w��J�����&��o��hky�{^;OU�tQ�3���m�@�Ӹ��m�ϫ�E�4�U��"=�E�Ш�A�[�f�Ϛ��'�q[�7i����ڌ�-=D�L����؜��	�.�v���>�h�N�I��/,"CN�ު�s�E����2�,��H!�Y���L���Qpb�g�9(����6����֣�8(��1���ɮ�0n�\����=j�qG�qi�p�[��X��5�ծ��$v>݌ĺPYԦj*�iM�H+RX�sE�HcM���q���z/8��o��Ŏ8�����5\�r�rc
D��ڭ��F�֡Ϯ��}hǏ5��f�2��!�gǨ�dTd=�<�yN����hۄ�uC�����'�5�ek$��sqz1�����s�ne[a�%�xyP�W`CF �����n���I6�ae��p��e+f�O�� ��뱸��9��
�l��4q�qK8��m1 f�j67�`:9�	Z������{(����u�=6�ZN�=�Q��b�v;z��T�xRa[����d[O��Ć�ͥ|�3�!hДah%��@ڎ����������>	�6���� '\m�\b�������y
?�"d�`�䔍*`��d�B�"� �^������b��p�-��:8�����ڧ !�ݦ��xQ/�ٍ0��1<�L�C��ޥƼͅ*����=n��֡��mA�Y9��,m50�/�aF���k]	�;���K���n8?=�_Տ%���2�NSz[`�w��m+��˅^YKy��'������V�n�� ��mD@���*�p�j]�ã;x�<�����T����p�Ǎ>E2��QtO���X�~ޮ?O�t����\xv��p7jR��.�]���c2^�0cҘ�ij5fh)K4�j˹l��#	@�q�ki��K8��QiF7��#�x[�3'��W �����`�Z�{�f�eӽ�4â�� �] �r�<7�S-�US.{��)���`Q,���4VT�,놕�[ Bȱ�m�[��i�OK���mf3>�"w����َ|1�A��B�x��"����l�j��߱���a�oc�6+u®k�^��k��*&�M�-��z��Ȋ��{[��ְϟ�"�q�d��t,��#aA uVFwC˗�M���#dӫ�1�Cs4�̈́by
3��yx�왇��
ݽ;��.���7_8�XEU�:��s��(�s��k��ivҭ���uL�����] �:�Z���&_9��;I�]>K�qu\]ǲ):�h��2�t}�<e�y&�fߜ���MCWW�Ja*��b�˹Y��8����m���W�2�)H2�Ҹ2�� }�	��Y�|nΛA�x�>4zDi�U��Q̶ÕC��Q�%��y��8u��V���`�z"B4b��ty�Fuy[>*�cj5�ol�W�����sm�����8�@�C�4���g���������ŵa�Nl�tK^(M�/�Y���m�����BB�6���ke�t�M�U@�^Ai�fX+�	���Pa�Q�*90kj�%¦�S���M�[�bsJTӛ�9}0�;ٮ�,e��I4�6�C�W��sV�����"@8���si;�8^g\�u�nh\3m�@�yթ@,D�fF�<����pܥ��j$�������E��ry�j��9�5y�6��$!)���r��Q�$Ɯ��Ź7�sˍ��r�x��[�	lO'!<�y�g��i�֑ܬ��&��o"n� �@�M�A�]��K���d�<,AQ�9���Ҕ�	g<�ظ������zZH��OG����=�u@�g3}.��֔�R���a
�6Q�1�ֻ�wj��U"��`iO0��G?R�U��)1�]��i�=�p?�l�N����0&������t�t�Ȩ@���-7�We��a�\칋	��$+�.' m���Zhj��i��j+�_y`�x�n^J�Z�{��4jɩg�����ND;�V��@D���Qޠ�kp��S�N��:B��g�����~����a�r�@�P)	QiOϼ˺�]/���Lp��҈Rf�z�8v!�hã���q����z}��{-6�Hs[9T���e٥vҞ�q��eAޖc�L�t-��AJ�aBV�o]|��'ܬ��=O
��b�}�2j�.�4u�t��kf���ժ�%��z���©�'z=Any�+�Qs�����w�����7�|I��r}�;[R~W]�(��ځg�e؇�'/�����8�Ǽ��]s����yZ�:�x���Qz��0P;�� n'���o���oP���lub�~�-m5*p�ĵ0�+-s�9���<�r�Sso<�Bd�ș,�x9�giQ���-��KOf��)1y|��������!�3�^*t��T�Q��ob�j��r&1��X�5`��:$5\��D�j̇]詷cޞc+�6�WHL[
NZ��#�I�4�:��6��~��Cou�ǚ׳Uj�C�U� ���F���I4,�� eW8v�bw�݌I�����rrc	�u��g;�f�aG�[H�� j<�C�P+����W�����9k%�\�L���檎��k-��{5έ�K�����A�O#���W��/���]��˝���%C1v�o�ʏ����V�M��]�YdBz�nd����Kpuj8Ӗ�	5v�]��>�ԣW}J���ܗ����}®z�_D�n��w|:o�~�{�0��C	W%��(���fYO��)����n+��n�6}�э��e�&��KW�E�'�`�
%E���G6-<"�,���K�Wj@�G1U�hbUK^!�m&���K��������l�FDҹ9Q��l������hd�5� {���BL�S��b���7Ni�A���-+�45��i��UQ��zp30�͛Hk .�-��"E��^��y���4�(X�zX�v�8���1�U����uL࠭�S.�m7�W�D9��vd���Re�6����9o'&�_l�P�j���v��8gM��}	�8�)>��0v;�+z�Xg�"?}(+U����� �?�ؑ��NS��l��7�lA%a�np�̚M��ב["i�]�xW���{��XV��di�l��nGNdCy��� :e� ��f4b��^<��q�e�tb�W��t6F�t	I��vg	�h��,�%�K�r	Ғΰݨu��m��[!qk���K	���t��Т�zs�D��QV[K�U���;�Y���t�y�� ��-~8�q�vsTz��y���>��f���c�/�&>350����j�ǋ툡�8�w@�x�S�����׷��5��W@�0���j��x"��&������udNZ
���*�n�K8m�I�wewm�6ڜ���Q(��l�4Vp�+��^˵� է�����)ǳ���>vf�y�>�s��o{��SdO�`dl�ZRFU�J���Ͼ�{��3��T���|��(�֬�μ�5�w�Q�D�'�U<����}�(rϸ�՚�_H�Şlo9�I@����䣺M7��H_	|1�2+�L,1O�@��֬U���
l���i;�v�m\�����K<�/L���U�3ϑB������:`5�mf�A�p��Ͱc�5ι[W_[��'��i���Fv%��73RASg!+1���j����X�a09����jM�]L�w���|	�\L�[�[��C���y
NO5�%Ǖ+L'��vҋ�P3��=;x1�S��]R�!1k]l޶ ߷�<>��^0�z���E��H�T��㗶�N�9��jy��չ9���[�`qA�H.7^J��ei�cNe��e��~=K[{����յ�3�S33���m�p'�Z�����n3C�{甂~لC۲ ��g5�����Ki4������m��9�1��8��I�6� F�{t:h�d&4NP�{��l P��.d�%%�Rd��b͓�y�*h����\[����o���\�_/Yէ�ڶ]�N��|��b1e�:��kF-�?�T,e���'_�t�i�:�b��RL{�A�dw�E�Ʈ�"F:9�[��e�3��Âp�yF:d̂�un�C�����Lc�!�=�T�:���]�}��9|��i��*]]���n�<�'V��$���=�0 �mB�&�p��F��񉀺�3!3.Q0o)�>X�#xZ�y��O#���WiƗ+���&6J�)
��(�2��W&ۮΨ���MowZO1󭕖�C���%[��{�� ��En<{/,��z���k�Q��V�_+�D q۠��t|i�t���U�N�9[�����3(�����˫�c�g�Χn-�K�wV��ڲZ U���g'E�v*���/���o�'Q��"<�Ĕ����v_C���x�۬�"C�N��
��@����}@70���m�.�V�t��qD�9b�u-�̚y.cC&i�M)g,>ɔ%#Pf�\T�����S��w�#�QMG�^Ol��.�U����,2�P���F�rpȍ]n�B�)^�.L���Ղm���=�<.f�B��/EQ�"�#Fch��q�+�;�%G���h��W�h)���ӝz;9w*\���OfV<�g &����9��S9DGO	��u�VDb�HVp0G|搤:Bնб{�E&��z7�b8*6:�oyVGx����D� ����g+��N(�F�n���5��6��,�;d�n���2*�aTo��� �5��Y� e�5�P�C!䖫Vt��i����D
���|.�9F���L��]JA*�ë���mk��j��O�ZCDv�`�V��u�\�ƂB��2v�7+��l92�*`� ֕#�3��$gWW.��Ȯ�/
`���\�{���/�_'g�!L�.�������R�#;���O�2�Er�Y��h5i�P�@v�t�˔���c_2��e=�Yº�_+�`��L�G{��b���CG0���ڸY�}�hN����R��X�熯dPX!�|�IA�{#-
�s�P ��H슱W7����vN��רw_B��\ m�)�!M�M�d�r]$H�n���U����s��(s;�waltR견9�f���l�;>��i<i���:�*�Y�v�H�kk�����.�g�E����!�w�����.������~]bn��c�Rޣ�9)5�����y�u��;�6k +XT[�u�>�.p8��u9�9��ӧ��3�PM�����.Y�\��..�ۛ=��SBvZ�nS�0t�O��;7�8*ż&�&���Y�����c�ζ�U�w�  V���N�a���1����γ�H��#M�槹<F���,Ɋ���K��:���úe!�:D����S)��ݮ;�rl@N�L��K��K8-�%d�s6�Z�G��e�C�K&�\��(*�(���_f�t�<Z��}��o |m���Х�H��cƙ4�EFCl���MG,A"K�{�T��]�i�m�uQo�v�@���j(�5H�)�-
�Q�X��Ѧ��d&o�rN���"�L`�3*���^?��o�����������x�Ϯ<=�NO�XQCMdQ�4�wpȮ�'k1(�&�'3#01�Y�^���ooo��������\y�=���4�L�FE�8Ff�����Yf�8Y��o��oo��ooo�����������*�a���7t���lR��N�a��xa��0D9�f`PUfg�DCDU2�A��9e�c�cc��z�fe���6�eLEUiD��b?-��"��#*�,�12�̗c�&&���"�K 0�������/�l.A�UV�STU��v���0j�z�����0�����p��F��S�JVYu���$���AnY���Y��I�>��dU��2�TM
�j�I%6,�)|r�mwV�� �"�Av��ܳ�L���'U�U�Otf;�ᴨ����KyC�A�#�T���{�҂N�E��~��ʢ�ѠRh�/�?T��?%)U>}���lTv� s@W��@�^�����Y ��ZE�7���A�R+�NBh��\�ޮ�]\�:��f&�]�(�b$6K���x��֩y`5�p'�ꐓj�3ylE��G%�WtF��z�6r�V�G�����,�&������7�8��a4�x]m[g�+,n&�jn"\1|��i�G*2;[�o Э`ߡ�,^��d�h�&!>�zL6��gr2E��ޥƣ�i;S���zE�b,<���[�� f)�j8oQJ��c3��m�P�¨�Y.�2���DkޱS�龁-Kc�o�'QA(�尡��ЙB���h����L�3y|.xh<S����:}p m(:seV0ZEs�/�Y�x�yڤ�֘����B�vl�|�h��,#���A�Z��ݞ6�h]a�P_���sʛ9L�8�G���WQ[��/�.����(ߩ���yy�&
Vg6�&���"YWk�U��1�R7�����6�v6z�&�k^|lŻ�&��W��(��fc:ȉ��47ѭ"_=^y¦�'�ˍ�=Ў���4��7h���SS)�N�t��۶�{�u�����*u*��\e�/�'="��׻�S�6��6KM�G�uC�{��9��|:�kvr�^�3+��5�lu����K���ŋW2�s�g^s��眯�3�s���҇�dHe<�����JZ)�ￜ������tͺL���	�t�B�0P��S%^2�.�@�+.c@� ܙ�Ī�ם���5;�(�w���ܓ�#�o�yMc��UL�Ze�1p�ثh<_��t�]����)�2�eB+w	{�4�j��Е�����uQA_t����c���c��AiYJ�a22_�	�-ɢ2J.�u����g�)3p�	W���e$�@�.E5����.�@	B��^BX��&���i
�v�|��(�<�؆��T2ޒc�Ƥ��L@�aIk��/=o�I���-\��5�Xˢ�U�$���O��|\	3��T��$s�,�d��ĥ��O�z�w��9�^P�]�g��<D��	,��d�ײ�17��Q�E����my�)>
����?C<��<FFՌ���!t���g����(����F,�5C�����nE�k�0��]�+�(�V�S��S�.2Q��/�a��ֳF�Ǒ�:#Y��;cv���2�����r0��1#��D^�w ��i��ͥ>��^�@��1��.v	<�e�Vֵ���6���Kʔ���®�,�t��nOݾU�N��)�.�	q"��J]	ś������>Q�}��k�&�Ò஻"��:�VS�*U�8 3�#�	B���{�򑉇"�N�����<
���Z/��)JR�k �t���]����gR%B�oxnV��Ś�W��A�{���6�>�0�GѼ�/?:/b���>�a��������leAh�wV�V�mNj�<˚)�K_�5>�ez,o�Z��0K`X��e�%�X��X��#Z�e(�ڬ��u���= �AN2����=!�V���2�>d�	�<U�1)R����O;����5�s��dgP�m9#7����*<5�5A+d:q�ca&�ymr����h��̼8��&s���$�7�9��մ�8Vq��=��Wz�@����0�D���C�ys*-*tf��k��o'[8�Io+��~w!2�����e�����C�K4,'<���*�r����L�_<�Q�a^*�ݖ'U�+�N�@^b^\=μ����i3wF�ۚ,�C��.�����p�cُI'�yH?��ٖ�T������X��
�u�±5�GD�Fk}��'�g:��+�������� ���,���fX�`��9U��8�=�<O�𪕠��=��u2�%�5�3k�Z�Oʯշ�=gy�%��շC�1��5S]�}�3�ߑM�c3V���:�s��CH>]~T�
�#|\��Oi�3�-��C�$�uT�j�M��G�Mkp-+��-Xol��Ҕ��-���h��n�N PZ�	4�X��*ܾ��{.�s�}��}����;��~���C����� RR�;Ͻ~{�����y�?>߭Δ$�2��@^�XC9 �w�WY��|��ޣ�V��\?�e�+�ϥ1�VWp��Hq�lV��Gue�uIW1נ�3��S-�C�K��<�o;�hE�m[5�]����N�x�ځS��1��$�ituМ�<�,'5¼n"�eIn1�h�Ca��R�5�$��Ջ[c��~�)����"�'��%��dɏ<�yO"�Ȏ�tU�3�y+�˜��"-t�F� �_�2iрby��6pڠ�E܋Q�(�bB��	R#&�윽�O�}�L�C:x�y��v]W���{�2�J�sq��aH�:f6�!�����W|�s�����|��	��LX䆧��ށS�ό�CΤT6lA�v���ߋ�n4Kh�i(Tò�WW��熞�p���;_��藃��Ψ���Xn�<a��Zq���ir}�d��&nc^�����R����ᑴ{�G�ڵG�TC�Rq瞋�ل�*��b`��ڢ�7
�zY��D��������RyLU,���o����Wxȋn��̩��Q%�b��Q�zͬ���#%�Z�<����b���t�|M�_AIg��=�4�!�I��Ьg|}�Q��_'��u;7��@R�+,���i�}���+3�N�`硵�[ݮ���6�*t���Q���'*��w���F4.��,�R^10ы�,4��Ubη7�޷;�����h!��Z�.D-~՛o�z-"H%M�b��sq����C���A-i�ܱ��)3*@�a���n&�8M/�c��I�;9t=���5]���Gz+�D Ƽ8�m��4]/��B��Gέ1����85�4�˸Z����[;!q���p!���Mb��ɐ�h���z�۲�<=�P��,�/��L����j�U�ҺN����b��7������ӗ�e@L��g�k{k�f_��1��e؞�y�C�''��e���y(��	���u�<9���[��>��H4/���[V�{h���1�g����W����V�a�!{]���V���&���z%:����z!A�X���N�y��Ji��N2�\L��z�r�����>*�w�Y����R��c��ͽ[1C+`��e ��7�J�Y'��JalsL� 9�G�W�ۃ�ކc�Z�?�<b�[�Y��v�i�z�T�E�└{���x��[�7�����Rڄ_�K�I8�V$��5��A��M7�.���5y��Sy�a	.9�!����/��l�\���omy�P�8j�� lgTۋz-pUɌ���n�"0�+�\�[R�;��k�Y�n,γ��IԨ��[';#'f˵Lݺ��b`e��O���2�4�T�)��@u���S�Ü��Jo��[����s�{j���H��m�b���ߟ~�~��0�)x�#CA^4�A7U|����a��H��=K�NzQ��5c���qX)��@ځ^2�^Pt֡]	]5��v�D�bE@^����(��p���r�Zn�z�rv�p��K9_rΚ�U#�I>?5rʮ;q��Îς���y�!�X`N<�3�6��iʻZ=�OA��E%K�d�Ga�zs�u���L��mi{��\�FQ���,��,Dz�3҉�<��/7K�z�Ψ;ٙ�X3ۜ�!d�=Tf<�^_�Tz����kp0�C��@BîQ�Ƅ��'*������5�d�;qQi�4��s�ܴFe#Ux�{�9VٮH��q;��B�e˯:�6Ӈ�|tK=>R��J� H�#����=�h9R��7�y�=C�pL��_D�x��6�x�^�Ǒ�d��~~���נ��Ȏ�iL�*#�`k���e��#	$��W(P��M���P�64FZ:�ݳKsB�2g�5���n#�|�ޒcx��g�&[�9.��#���kq��o��K��f3wM��
yosy[�o�l�w=R����b�L�v0��g�FK׎��%�{�RO��ʴCY5b⒀y�#i��<��2���ް���RR�yٙ�$M\X����Z��q�(V�΢(�L�X[}�jlWt@HaT��.J�ޜ2�;cK��{)V6
�y�v�=\8�A0�bם�)P"�	�^��>�y�y����o3z��$y�F+�Ｇ�D�w8�}4ms�P[������ܪ"�$�>���=0�&��r��m�k\L�Y�ࡏ+���7�3�Q�lå.��7R��4�Y�j6T���Г��b{v3wK��0��h�M'��74
g�M�.ݜ�i5(���<��0ױ�K*�d�3�X�]n1�xs!)0e�Y=L2�6�3�9�N�y���kŕ�6��\�4�m�5i��0m������}����q����@P,��nk�ŵv���޳��|�j��}5Q4lc��m�Jg.�c�Lk0���o46�W��VBL5ޅ��ek:%��
��N������H����8`�}�J�N�
mw�Cu��P5l�H��Q���1u�I��#v7ܩ�H�n�^0�CUxsH~YB��+xc�[��pƄ`cAvn�ü��MtC�G�L�k��f (`�77cy��.9(�ն=M���Q�)�Z�'5�z��)E�,C)��$��l�����	ϪfgK@�m���=��GiH���C#R�#�0���N.�*�º��r�yC'�5�}� ��B�N.�]) gvi�VV�K����Ix�I2�rG�q�D��X���0P��h�y*� ���7��,��V�K�<��&E۽��~���i��ι!DE����u��"�̂��U���8UX�̪�7�����D��g�󇏁 ��ĀA ��ʼcXw��t�N�/G�G���L��7�s8S�`�_��Rm�΢P�,-N�%�ڜ�~�̛�ƞ�s���l��f��%C��''�Ј�<�*�X��p*@~�Y%cT�vWa�u�Fn1IAS,���,e�M������ ���fO�F����j���%���NV'���RԽѩ!����\v��r�#/��H���Mt�x=�Fo����g�x&��-S�O���}�-��w �~m%��ٓjq��BO�
�.61[5�����3r�p��i�/8�V�V�&E�H*`�y0in�)Ƃ�u�$���a5�c�!��{em�[G�:��T�/ݛ�;&-�b��4��=i�ԳԸ���>���
��i�(6Q�|W+��֢�+��9\�G�T��B9�ر�����3r�vo��7�m����H��-�T�6��q<mV��"d�9f\W0���X�0��&ɞ:��h�ջ�U�f�
�AW�m�y�9M=�*=�.ʱ`��v�r�WV»[J�\%��"VS.�OB׾���T9=��:$F�5nn�x�H�eq�I+��S2����ܨ3����)^g��×�,�/�\�����L��� ���a5	��a`^�{9jӯ����}V���W�\��.�r�Q�}V�y&IvikuӔ��M��V'ZKlN�q�:5�K@}}C2�������Unfu���x�Ï�j�{]�3�{���[z�7�v����Rx����yb����x������
�h -O�׺p�K�&b��2{*o�8�'���l!�fr%� �@�`�Y�Aa����j�3Ͱ�v�eF]Ҭrf{!��^�B]���W��=yI��X6-��:<���'y��BM9�#��8K��[�y�R͡�p�aD��Ƙ[镔U-U���أ�:����D�r��>0��[}�Ց�����V+2���ha��H�-^
�hNɭ��e��)(�#ǧ�E�O��׊`P۪��A~r<��,q�p�7d����_�+���9� �6a��l ��/u���O�[�b��ǔU|�J,���u"���4@wW���	M`&�'(V=�V���L���`z�a*!�����KO��u�^O��a���he�9���8��,�ҭomW<%��M�l�g���Yi�I<�pξ�L����(��(2Q��j�4���hx,'ze2�6���u�9gl�d�|�o�n�Ne�t������O�ء�Fˊ����/�mX�]��=���t�h3���yb�+	�3Upٔ�n�*�mT)��ZS��e���Ȇ*n�AwV��y�� �yUG�&@�f�ܥ5�e��}'p�y*ES.&vx��ȡ2���g���1&S��v_��q�U&w�p�>����!��B	���Ϟ���j�r�����7SM��m�Q鶧o4j
T�P_y�+<�m]�:�ۦ��Y΅y���r��{�S�/`�R}d�����)\�z��]���Et
:���.멋baBc�������h�oY&Do\�è�[a̍ׯZN'[��}H�肹E��M26+���vU#�Az\yy�i��|7�.����`�&z�L�C�S	�ZRX�Fz�i��5�w�"��ۭz�CH��K�X�0�[�ۇw#\�!�����v�x0+�q��{+�'�tC�Q���Em˽g(�^P�W���>HZ�6q!F�p�|u���;a�P)G%;�_�S�FQe~����7��X�?ӕ���Le�SY��b���&H�`��,$C�HQ�u/��{���y��c�=|�i"�m��@ƳK]�Tx?�ӺT��D�U!� 'um����X��Gj?���2��@}�!�c2}��(o3��>$N-�~���}���>�S��e�mm�]��z��*i1i ��Px���W�����ۤЯ%�9�_zK���	�=��0��T��$C-�s�=�܅�ǂ��hyt�vS�C�T5P��'@⬫s8����/1nJb���Ya&f��r��t5���9��{.^�ʟ�T�ԟ]�o*���b��[h��qp�X^�x�b��kF%�﫻��}��
�܌n�C�d�r|񎒎�������*�-�s�-Ѵm�WK*�m��y�>��t6�m3󭬅^�.�.��[��m;�7Bq�G���� wy�zq���ڍN��2��R�|`�?.��o��O*��{>�=]�ع�������k��5���'��DT�}�"�/�Uok������]BU�T��fz����5Z����Vz�V�
�}������Ԧn�Vsb��:'i�cV��d�]�a]j��),/8�(hR6j��e���=+v�uH��EL�*�=֠��uj����(�6N�V��څ���%���ew(	������Je�k #�s�hp<Ot�&
�kP1�y�;ѡ^_n��PI���܈;R�;��D�l�4-�α�h�	Ա5bZ�fp��o�]z�;3�-�g1idA��+�˦^�87[&���E��i�=*6�����C@'Sj�Z9�([8Jk;iҝ÷Qaμ���t�jƼ�K:*��{�ݡ�@ꍺ.
��o��9B�1�E�˂^9z��*5����ݻ�wb�H)�Ξ���Gm�D��^N��y��g\���}��e��N������پ3ҕ��oݷ������Nd̨��̏{�!�Ks�<E\�x�ھѦ<�Ls7ϒْ�ݸ.�j�$)nc�XWd�7k%	�E)��O�˥X�J�k���;)�^�L�x�ֵ[�٭�:+�[7��h��/�a���V�
z����M�,��/zp�8o\%<#�e�Y�ݜ�;:����a��%u�m.�Q�,��fu-�F]�Yl��g.�	*���N��ᒲD�Sw��K�S;r���9���>�'`cc���h�a�Pae�e�pb��\ws5�|M'Φ|�꒶��yZ�R�t������L�,T��gD���a��{��I�zV��v���� UfN5���B��RU�f��0�ɆV�ݝ�J9y㻩)���=��&�f+�<t�Ԑ]��㯀�cy��C5�eh,�w�ԻW:ڊ�Ni����h���pb��]��h�3�U��r��<�Nf�HO�k�u9�,M��կ�7��s/=�i��f��Mg����1�����3�y}z�'+!���wI�yU�'R[�{0r���a�g��x��,
ޥV��{�]3�!WL *� E��¡����YD��;Q��4�a��l�?�u׷��׷�������x�����$YdQ}�Ē�Y��0��3
�2���"�ɡ��L����Y�^��_^���ߏ�����3��`��9�f:E�f�dffnn�9����F�fTT�T޽��������������}}f}}=h"���2�3""��ȓ�ɠ���"�0���&>��Na�FA�,�7;�jL�
�2&���J/�U�w�fbQTS���������̘���#'0£11�(�c ��6�2r�0���Fq�0�%��,��l*��2
J(�����Ȃ":̢���.���#(�1����Xl��bw��DU4��X�u6��Q��Qf��lQ�d�E�fXm�f�a%��y��SQ-Wq�]XEfFw���]]AT�4LA7v'xcD1IM9f㳤M�d�H ��G��x
����
*]b� r����l���_K.��捰
��4���a���j-���_�~���b��x��=��{�O6�}����Z2e�>/^Q)�QL6a������0���ܦ�I�L����n�7��g���B�3>(Jy#&Vs��58�,�����R��.�ۨ�`�kH�>�zUٙN���ó����3�oT�#{II���)26X��X�Ds9�Xd-iuܴ(�j���n����ɜ��\&I�lR}��B�dv�]��i(��K#���kE�Q��Y�fU��	H�����X�B"�|��UW8���8�<)I��/ب^PYX�Z�'+e�ѱ�9ݑ���U�4�6%NT?�.fZ�+	�8����Ϻ&�M����\>��s*둃X��Cp�0���M������C>�bc��)���E�3�;v-�����sNBG-̴��U���v~�;r�@
���Ī!)�9K��:��i��`�����{��3O���Z�T�K_��9�Ԑ����5���G�9t^�ߜ�|0���ɩFՓSz�P�#���.k_y��eO�=W�ד��2��R�n)��5�-0WjU����V|�jB{u�Y,-m@�v���soW��臉��qX���1��꫏;ߓ���K.��g��B�'+��hy�c3���击�V���M�L�Wu�J;�g�9H2f��FAsչY�=���HY�]�a�5�'����<@#��<�ի��)B�~��=cϦ{�V�qqR.wY��h\˅Z�`�j�Exe���55�dKC춪殺��m#�fH�����h�CY��ރoC�s�3E�6%��"���-���G���a��|L)E{ܧ���㲉��'�����|��r���gK�S�G��b�:�s4����cBW�	&��X~z!�9�u����D25*�xmٶ�3x'�2��^�U�yK5�I/�0�B]�ƹ�����s
	��y�%�����u���֝��+�&�O+t�gH}5^��RN=��k����Lw�D4Y�,Na��k����ҩ�h���S�z`0�Ǭ�A�P��})�����U� 4�B��L����5!�Q�Y�P1J�q�7.����������(𚚀�n;�F���uÛ]�hU�D5L���;5ws-��m��iy�����`2�A��K��[i��`8˹\���	T+(ut��O���j���3S÷��H
�^X�aY�Fq��R$����G[����_[Q=�/�K��k�<��:���_^�(���N��ٹ]sT	���9%����cUr�)\�`�9WE��\�0��̾��lr�#�ź�o��o���V�*_}�x����\�^.���mp�ͼ�Au�=ΌfL$��d;+a���fr%��Aj�+{�we� H�NQ�����~�^�kl�
<�w�=���o�`@�I+�Ga�[����snF2�f��=����֨:�ˏ����)�p��GX��#�֦��j;Lr�)$��8���>���t�k��qK\G�T�CP�#}�X��gM�`;7�8�lgYp�d=���U:GRz}ހ���jq�\��v��j�js�A�sA�R��
%����4�A�9'�Gs5e2���_۞�hU�.͍O	Gs�J5�&���ȝ�I]�WH���=�˃1���� �
[�C�n*r����__@���T�h����S��ۮm���h���%B�D�L,���Pm����g<m���:��B3L��ԶOH���M9q�_p�\*7��	ǧ|��G���[V��*!Ĺi9ʍ�*�q�WL��mO�.u�#5�f&d�:�Z=)�]TG�L��S�ח���]���!�'z�7�.U7Q��h��s���:���yH�m-�`�����1�Zp��s�K;fg�G�m�����!���Bj/2.r�r-����̣7Cf�bT�F��AO���$EC�l��K�/_c���3^t��`L����̽�$5���J���t��ޱ���a��,�m�g���H�ʦ���PG�m2 ����ٗ�����Lx�6)t�̓�Mh��Y釱,�v��Q���QS�h�'�Ss��| ��� W)��UʌZ���M�"5N�	p�g���ʆ0��Lټ���cV��d'��}9.�h��e�t������;�	�Ѣs���a������m��ɸ�X�z}�j��g"P7P�?�WF�!"#�}���U�V.~	W�T��o>��g�iʋ3/O�����8������c�`g)��qM�`�(���f�o��R:�L븳гִw3CX�aT=p�E�\-��v�0�׌D㿹	ޗ~W���$刬�9#ZM2v�ceٚKw����\�gva2GY�� ������<���I���@ڔ,|8�"ی2^�)�Z]���7�[U��-Ù�Y��4�Jb?��z��O'd�����zI���G�Qg}�sn�k9��.laR�2�B��<"t�L�Z�b��5z�<�I���oR�x�h{L֬��d�׉Ayp����ly3��p�͛^i��>h9j]���.2��i|֭We虭w�sm�iv=��]�q'�C	�A�o�aE�W�л�(Z�%�9P���3&YG���9_VL)]�v�T����v���P�H�7���{:?d�����䍽cU\F�R%�*�5n�U�䞨9ƣ��ryV��}����a�Ҷ�<�Un���zX�����G�����%�Ցn4{p�p�WN�qi���y�60<���w�
�P���{�U���~�
�K'I��:.���� 1��a�Rpl7�)wc��}>�����di��`[cW�`��zF�,]�"�Ft�gb�yG��6�<1[�NpG�ٯf�j$�X�#	��6�e�09��C��b|TŘܺ|6\5j#�ټ��o^����t��Q~ ����j�G��'6E?����:/��w$v��3\�'�jm�s9��x���3�d��.~�V��{~LӅ,J�L��0�E��k�+�ji5؁�{�$u�`=3��;3���YK�&�$UA��͈T�0��N&N�����q�M5��v:L�c{O,�h����[B��3�J��ܙ6-���OD�����8E�[Y�2̷+q���-����ox����h�u�G���i��,�J)m�]�<����c��8�vD_�����O�V�=]�}�����]JV���27���
f���s-��˹JaF�ɭ���V�»�Q՞���oN8%�%:ձ��/I�m*�<4�V�!U��p+Nl�Ն@u�~o�~�T�z��WIV��X��N����~��X�ړK?���}��/.��L;�ۥ�,P��c���tW{$&�aa��r����K��۫�3h�d�L���hw-�� aٳڌ+�mu*d�qT���<|G�x��U��]�'7ǥ\�o�9��a�Xp� �O���=N[���}��H�\�\�	1{��m�܈��X�D��SsCq��ۑ��̨���S���&�O��lrbIf�w4��ɭ&�M���lȍ�]��B������K\13����-� �뚈\�ς^K��2�B6�E����N2r�X�Ef�d1Φ=M�>��|/�h \��me�eh��Mv�LB����=�������az3�+�s��-��zC�����)i�Z���4�:��\X��]�ݙ*�x�N�:>@7�Ӳ%�7-�-{�uY���53WC�tU�6����S��ŧڨ���y�w 	�p�\B*��T�i����J٧���q�������nݕV��_u����IAk]�Y�yd�M�����MʆXo4�"��ý70J2J�M`�Q�F9�^�l_ټ�H0;���^7�`2{O�:�ڛy1yBL�a+=��Z���'u���&P���/z���@칈sY(wc5��_d�.� �].�j*Kgm�= ��&��P�"��:�݊Y�������mo��р��ww`uwKWX� ���<��Q�*B���Y�V�I�3�*黄*C�X1�w;���T�ͨ�	�l��V�=�f]�z�ī���vu��6C��Pm�m�u����O��C�@���T�xVʽ�B�hTy����Q*�Y
)p:��q��R/�ȃ�bz���Oo ��8�U�kX����ޥ�
�A��lp�F3�u��XD��^��ǟ<z)?_�m��1���)ͤ�u�{׊���9���ȁ�������e�?�i=r���/���Q�q��b7K�ju�2���$Z��G��T�����{�F<ˏe0�cP&�sm�kC�l��Qڅ$d��\��O���O�N��ךv�!��e�g�����8W��R�rкX֮T�t�T��~��a�M���bW�ݻ�P+[��8r��ʱ��h
���HNV��[�cE��l�j�HKT�	�m_�������}=��a<�h���0l�h��p�����1
�Y��g2�Y:2T�32�����B�j�.+�v]=%�0�,0
��M��j/k��jl�0EHi����ʛ��L�x��f���l��T���ye"2x��CT�~�<��f;��O
daj���]^mT)"y(�r�1o\&Yf�Nm��� ����^�sQM����i����P�	���ɾ��WW�ǒ~�{��~;����b��*Wɜ�&��#�B��lє(\������o��ʹ5�uʿ]��w]��[s�w��6E����evp`�8ڼ�o3n���v=E�1��c������<�0��*#{��-�nc?^�{*�:�jH0�$coS���e����թ��D@0{G-D��lZcN��"�Q ��]�w��3N�Kv@'���b��3{��[��
�%@��vA�b��*,X��h�:�u����Tx,n748���$�t��T>�3��eE��$!v�Q��2�&C݁�*j/�,p��+�}�X��0�E
C�m�=�y��Ӱ��ܥ�;b1)��;)N]J��s��R|�i��-��'}������z��M�d&�nD��Lo2ƾ�F�1�2b��d˭BRO��I��q��k�oa�nx0.�΢�#��B�=����X�3%��`H�V��/�Ϯ3j�L���2�M�S(	A���Ì���u*����Үe�m�L�v�2�\�l*�t�z���]����3eL�W�D�C��3=jwq^��%����$��T�H�Ξ���S	�PJ���������Qqm-�w�[K6D6.��/w�+�ݹyy�Am���&.&�`(��A�k�)�w�Xhr�]ͳ�l9��j�XJ�
l�j'�f	ʏ+AݹAR[�uwtk��]=#����skӅ������}���;�~Bx����\/OY�_ �������bu=s���J�-QZ���|�Ք�:�l�gabv,�[yH��qޡO�ξ��y����W����0�+�]���9#�:r���'MS���og�*��\���*�=�1̵���u��8AU�J�k���2xr��77��]k|Lv|"���ù��p�":��˛zN��� Y⛫����[�|���L��Ϸ�I0�-�����6h4c�1X17^��\����[�Cgu
z�Z��gO;HO��f>w��5l�B�`c�N�������.:�:;7#�/����������S9��.#-�4{"=��R�3��MI�a�����q{-q9��w|fъ����_���N�-�-���
rk�������e*�)^G>��J�r��罵݁��SThjSR����'@��މqt0�p3C��ފt(dIe��~��ܦ�Yn�	Qz̆bbL�㔘��ż��w�S�ze���q^�n���$% �q�"�n]3
ef�o���x� o�ih�6��w�T�>�Y4�Q�O43+�:�{�;��� ��6�ݬ�b�T1�ҙ�b��Ty��������!z��T�T�Ľчn�S�,TN��M>ͩ������)]eoW[J4��F=�Ռ���3�8�N����� ��)�uS�G�*�I��F��A��D��R��w:�^n�&x+ދ�b�Gn.yWI���z�������J��Ṵ�Ṏ;�z��1���>v`���a�"i3�4�$���/!-K"Y6�	8��jɷxi�=��&_�e���9��`�gwnD*�2�QLZ|/�Gg�3����˞�=6�~�Ԋ�絪kӑ-r�e���A��S�E�+��(B��^�,�@�nCE(��u�+âU-| �)��z���1��R^y�R�"�!�mo9���0�%� �/�W���mc�#��KN8%���ų�i��\9(���2���]��ɴ���Ґ�ˁ���F�&/j!�[�C��c��1�y�q�oX��Q�ݷ�e�E��r�O�b�[($v�q���|a���C��C�9�N��l`צS8MP���:eЖX�@]ތp�5]<Ǫ�?0�\�F=������E�>mi�vs`�F�1MNS)g�1�;D��fs�<޾Q8�W(�ڷ������^�͏�#�a�!֙�*��F��2��t;y���!.Ga!�t!6/7dY��
ob,� -P�6�延[F�]u��q����#VB�2������,�a����`(:���l,դMx ��d������y�� ��\IlUnlL�u!��9I�Q�lW��"	hh��ǋ!����Dؙ�Ю�f_R�W)�v��+�wO� ._Z�5AZ�bU�����K.FO��r�̔�� []t��˫�y�q��b��WN%�+1�5k���ι8&��#��l��qJ�{�6��k��P��՝�$�@+��.���'r�Յ�S\���7և��T�S{;R����j=�v��G�����J㸴-���t���g���}R ^�y��.i��q�w/�p�"��☘i����(�����fc��f��b��G��	X��+����ժ��K7i�����e��09�2E��ۡ9ڼ�R�Fk&m���qRW�:���xwou�Yҭ]+�p�U�bO)��,Zk�T̮�W	�:��	u��ŘL�g>-�FxE�&�fޓ���7tm^;c�ͭ@qXw�
ͥA
�3Gj�k۷}�s:F���܃��34򡭑0�T`!`��e�7�;ޣP��f�ɵMS�v���J�3Ѡ7�b�(v&j��1Qص3E(s�5yi�������aa���2��r,���,ݾ�
�]��03��T�)me
N#��Jཛྷ3�$s*�;'V�q�ƪl���W/*�\t�Xk��7���و���kʹ0m��`*��sa�<��)ծ{�Ƕ��o��v5t7D���CͤH(#��hyx����݂�2����JY�Es�u	��Y0Ve�%ֈ�$_)(-�#��`�ԝ\G"�7�s��,���>��ۛ��%���;V:G)l�G��(h����9-�2Jz�Բ�@Y�	*uvAU��M�է�F�H'�9�x��juuc4JB �^	\���7�Ǵ�
qy�Í��*�u[��Y�.���*�蕖^��p�`wO:���h>�v�y5,��r��M����:��9������_E��k����F�)�J���(T��lxsl�I��@��<�=-#8��i���A�W��J`}�!Le�5j%ԩ�`*!�/�_'��Ko���/�ͥ���N߼{i�^���t�uV���
�h�vh��2B�8vl?4�t���ϭ��0�f�m"����˾��C;:�%�C��v�
�{��"�2����7흔�z��/r����Av�d
�&�5���`Hu��'@0���	-�Z��.���-��v�|np����s���Y���u���}����yD7 K��Sw}�홵�ιI��0h�؛��I���j<��޼8���z�����:�`mG���Rǂ��p�z]f�49�Tle�S�p��mT�\�i����n��zGu�zQC��f�P��^M�N�M:�x�7i��v8L=�.�V�|�oZ��'d�nW���,��X��� 4���a���E"j�l1��Ӕ�lQ�\�y .`h�4^BTF�,?]%R��ٺ������P�QSa�E��	U�[e%E*D��ځ��>��L�SM��8Ve�8�|�ȪX�!ɳ2gp��z�3�:L������������������ ��UL��deUwzuхY�de-T�T�3E�1{�$OO��Oo�OOOOO������ׇ�c�M5eaͰʃ7M��(=�#s��*K2r�<�&���(��j��3��>>�====>?_G��g�"��\�R��"��7Cm*��;�gs��̦���7��2p"�31�*,�"��)�w2a���!�i"}��n�
#q�b��**j����2��))��c#��w�6a��'�GV4Y��UE5�p��fEEv�FfEER�%UD��f�2��2Ȫ&�����
�H��%����(�")���eTfeQQeQE�U%ADUSS1��E4�Ģi�������+���s-̊�*:�c�Ƃ�
��"J>FDDo��M$����SՅT1d�MQDQSTP�dd��> Uc'�k0�G��]�i�U�i��j�26z���6�[r��+U.x�,�F'y��
�=�y�t�.��vH�l"�
�  7J�%Y;�d�^��D#�nKه����C�|��oJ����,�ӊ<�|�n��mO���kg�ܹ���0��h-<2�.��.�c0�_ʵ�Kr��Ү+�̅Z�?=ᝤϳ���/>N�	���˫r����:R���C1i4�al�U�i&m�P��j���v��d��O�q5���X�)]8�A\�)Δl��vB���`�(_=$�Ze�c 9��fm�"��,x
�Ow˭�]O!J"��C{W�S�|�[��\��m�,���DA�Y��1���m�x� $y����j6����Xe�*�y�3��m��i�� �Kŷ� m�r��⮘Vr�PD;d<m�%;��_{��!������[O�?'M^�a��N�n�2$ˠ�`��v;O�;+���-�[}B��UT�1L��Jb$��磬��]8�[�u�:��t*���4I��ʱ�`Afhˈ��gy.�QM��<��UǍ��-협�D�cǭG��S���:��)<Y�nR�Ar��fK�M���Z�ˆ�?~J����(�5+qZ-y�v{��d�(;�[�1W��L�"ù�W��̘�dN�$�ۖg�$߆�W�Du�ܥS�;!v�ϣ�+Z]#ěW7� ����j$���-�G�w����}Ɖ���1G�xt��L������@����`OJ�z�c�������ն��s���Ŀ�<�^E�yP�L�q����x��FA��aA<���}w���<����_b6�F�'���=Aw�[�]z�{`Uj�.*�˧�J{�m�<�z;&D�TTPfl���r���g������#�(�;��ōhi|>Wo@�֌d��{ǧ�=o�_W�~�}$�{��6=�CS��p�S�1���	~e��ju7Qm|�6S��D��X��6I�s�l�Ka���T�hs���l�B�i8�j�la�|M�+��e�v�
 �.�-hκ�`{USs��.S���rid���"�
k w���UY�/�E�I�qje#��=�XC�=�Lw�5��8��S���߯==6qœ4�T������ 4���}ɼM:���oX�[#V��9!�C�2 �h�
9�5�!<���2.�:�=�`��'��V��,h����=�O�������{�g��V�$��_�k]X5���7�#�~ꤱ�f��=����e}N#���Բ�O0>�T�u/U�Sփ���ڏ�f��k���}�P;���"ɕ;n�S�� ��Z
]��k�u"�2	�5�����a��g�vwl0هu\u���PN���:��Jǘ�k��g�A%�w����U�r0�s�%��)M�۷��m���20��t���-��T*�3�}�;����$V�U�n�]�2��K3�Hg��ė��Q<�c����*F�rVR���%Y޽�����v��*=O]/�eGf�'1פ�XC��o@�恩t�]��4+Z�l��u˦�ޠ�	����R�d ���=o��Ng��{1�E�֕�}h�q\�̶�wuv3nl<�T��\<ܒ���7s��L���B����Z���݉��t�N��ǻӂ�M �%����Rx�sC��˩�Sr�{U�a=�/M��;�kN՞}��g�ޢ+�����'`�Q����6���)1Z� R�ͫ\�+�k�tY��o�q�_�����^Ӎ� ��H$�g�� �k�SR�h��P����l�iJ4��ΟEڟ,v͉�T����5�e���Ɯ�3�8u�gfթ������r�ݹ��p��t;2�$a�:�At�Z���\������VW+!f��O��|���s:��{�e>�F tY���S�i�5֞��J�޶ַ��U1/��#4F�sK���V~��p��{�O���];Sp��P�[��c$3H�ٯ>�����Ya����"a&�y�<�'{�V�f�cMs�ؙ���S=r����WP7���A��t�=F�79lLud?���$�вFq�i4(���F�E�#�6�WqNC2��w39{���`ڑW��Sϫ���)���S��x�;��"I���v����D��i�.�h�K��?��+��YId��D�b�g�J0` ^>C�/�R�C�o札[��}����?'����{�d�%�%e)�Ug,�!0�:3\�*zot���M2-��;���L
���^/
���oX�X�%��k�m&��9��x�ǐ���Śd:� �"�zY��u+��3׬ܚr�Hؽ>6p��LVD�0owD�?�-�#L�������y�j�ކ�������s�H��x����E��sY�{h�ó_����[*j��Y6۔��QT6�Qy����#�ջ�*f��;��:.!aԥX�0捫�G���SA��],#X Hu��EJB��;��ŬO���7���˸Gi�ɹ������vɒuv,x×�}�_���=˹Wv�O� �w�7�Z�eS����3����_=�97ks6�\i��"��Jgջ��IR]�l7+Br�c���@I�S���Q2:���(�qr�%�D۸ë/��s������+'��oB����ܱA����&̶�w����`�<��C��*��Ӗz<� �St��:jsZ�駽I<��$�M�U�\��ߛNoo{�T�컌��x�ە�*uR&�[h|�)����q��s�ۂ"e�y�k)�ܖ���=���g
�W�Cj���Yp"�7�*Yߕ�ٗ��/��"7�u�p�$ќ�Q�QN�x`Od{�|�Mbt��/%�G)5M�ȇ��^�SYk/3�g2�z�S�r:0�y��h��	���֥�cHܱ�٦�Y;ox-٘0�,�Ӓ ���*��o(��	��6�8T
Ě���-ս�qI[�oO�މ�^�qRB�-t=�K��ec�c�i����\�v�j�s7`g���;�1P�b��L$q(F�Nat{�X��voMRϤ���ٜ�#���:>F�YE�h'KM�/^&��Zz�u�*�@��.��b��O�LS�;��T��:/ih�T�U�h�9(��T�Y���6�k>;�~�/�>��3x���q�m��+�C��\���2���c���3"�I(�x�$+���[�[~�����y�}��M�8�~�~��{��i��É>��VP�;�J�
�m5q<���>�Uf湱Af>M^rl{����B�6�Y�G�������Kj��x+�5e���ij�1��7lL6��pݹ���l�kT��GU��F����Wɘc>���Zf���#_�s��'�y.3�h���q������0�6�;	��a����e<E��{|�B��80]�
�ٔӝ��ڞ\0��Q�OF�s������if�d"m�xa�t,]��)������t�N�P��8]���n��������4� ˹���[�K�";
�y0����h9ہ�������ןQ�wVh��������f�������e��d� �G��S��3t�z��B�bwTt�F��.�=J�[0�R�7u=�e��X�.dW;�+mt�U�>`�*ț�d�u��xe�+zt@�N�n�|^2�w1���Ƕ�e"5����&z��`Ƴ3j�k��Z"�1�ɜ��=ҢɑzŪ�����8�n"�(��6���`� �(��{���8w�O;n�yۡ}Tӗ���3�C��|�9���x���~�����_i��֗�gq�����TG��)YkbE�pQ�wj�t�d�
�_\�݁�@9L��:��d1ڟ�W�좗ܿ(��:i�*oپ8���گێ���A��Ad���v��wf^IMǭå��e�k՝��.b�c+V����ï�w������Ss��W�V�7G������y����=-{����Vz�=��Ἔx�@1Vt��7y:�FQ��+�ܝ�9O�OY�*�7>��������6/����N�yX��|�gfd*�<^��d/Lu��uʺZ̲��`S�[��Ñz�_�$S���wj6d��۸��׹��R�4�#vïQ�K���l#�0mL9s���*u�OJ��U�V�&>n�>"��;,�i�p�'ڳ�q�����G��%cݯr�$�=��y&wt�guʺ��ᐹ���]�/���4�hU-��q�WmWP�Bh�y̗Ҁ�h��s�K �@Q"�m�
���5�S��;j&�Yv@N�gﾠs��#q}}�t�%^��,*q6���e�q��e���6)����dZ8\m��t��u��z�A:H��A�i����Z����H�p��twsN�6���n%��P�ػ��FY��=6d�;�P]SO�O���\�$]xh�DE�����S��l6����<I��Vh���7�n��T`t �_Hq�ɘ�?"�`�w[����r�90�χ���3�1��m���z�lt/=����Єb�T�,�nc\���&"�j�WI�1фf�f �o+J=0��m��6)�d���}��9<��f���LQ�4�D���(d�>�U��[�m��Y���6���)��jU�ټ�Y�r3��_�Ы/=�e+�W������K�Ѵ�5�s�"�W��a�?NN�l�UxJ�9',��ߒޟ��^p�Mu�t9BtN�Ou-�1ɍ����ggms[[�NW����7TB�,4Ԏ�(�⸓��Q�{Wn�b����{WL�@oSo��5(R�R�o�'Y׼�R�7�#��MA����y�NA�ܖ�������Xt�DLO}%f���]G.��@yP6i���)b�T,
PB�f<p�k&����;�1�C�9��eK�n��G������>�K),\�"��쌹�}�k��8�yz��ƚ��v|/
�؅�,U�,����ۏ<u��8�(�<�i�l��э�5�\�.F�\"f������U�lfF��M�{��w��-7��ɤ��<�ge��n��~�֊���GM�I�1�Q�
�Вt+B2�y��b���c~8������}��~��D��V�&���'Y�����u�Wz���]�;שE�S���c���r�����%Y�}�u�=��7֯%3gX%9��f!U��}���J�Tz��ٻ 6�b�Gm��]�a��9�r��)ף@̾�g�`|�`I�F_H��z}b�ܘ�ǎ���Ԍ��}�A��,�-���|)��*�ӣ�o���H��aӦ�-��~j:c0�]��c4=�:���Vі��@[{����-d�Fo
�tw��-/r��H+&@�A�͍^n�ͭ���j�,R�W�W���_L���XB85kB��F��p���orͮ�!Z�g��b�T�x<��y�����s���|ۦ��M B�i�+�8��A�e:�T��=1|��8�1&걳7Te�O�1J*��o�=ck1ᘙ�c�KbQ]���j�����D�=w�YZq�[��Wy��n:f6�W7�ύ��Q㵵9q<g*�9�M��57��䕻�6ך���V
�o�G:�a��u��i�V��u���c���s8�������6G.����-����v>j�}����d�^�>e��"�o�Ъ���c8ל�å�1g�����m7U�rY�HHw�p�r&�F�Di��d����נ�܎�����9�UW���Ma���[�@\��-���G��>��<㳂���.x���0
�w{�v��%V g�������D���Ѫ]g��J�^J=��hPw7���F�Tm�5=q,�9��gI=A�V8ed����FgW��������g3;p�z#n4hɽ�v���(!�����!��,�:�N[F��Wqra��u+�̜5���Ya�*�k�=[mdUi����c�sX�Wu'ݚ�+Њe���+�:�@��kvY8��Z���z,]��>Z<��j����3�#��m��-�*�)]�qW�a�;2k�[�ͮ�"���}�W+�Zm��Z�nsS
��\���^�p� ��N$6,h(Ί�W$7t��;�Ѐ⁇��gL���K�q��so��V��9����lU�)�cq�X��lǊ2%��������J:G�.�o'�I�˺Ԥ5����]�Y'��i�q5w}�JP֪�a�]W��i��8܇�(��YS=Z),�ѯW���ml��ӣC�5n�ʶ�n��A�ܳF���[�en7�HÎZ}�ћ�.�@iwV�\�h�҈��+��>]kD����z�Z��ج���ڴm��;ή4��upWb���
��h�Uo�f�@�@-��h9R]�O�Wc��Tp�gn��	#]k��*Ȇ��FOPU���@mf*Ǌ�r��1U��������[�e�D�ٳ�&�Q�����sn��D�f�`)��NJ)	�K�E�TQ�Z�)��9׸r.OR��O�&K�?�
c�Z���z��S�]�^R���wvX��9�qc��A�ʠ� y�d����l��B����AP۩���VPb���(Rv�l M;\WL�Z�u~�}�<��7~��۝r�5wTI�qf(V�FY��e�;��9ߕ��7��U,n��"��h\G^�su��zz�&��Ҳ�볌E<��D���|-��Y�������ㄧݛo�J�^�ln�z$Z��x�_!9Ȼh�+	�i�hH0��w7~u�*=hpj_�s�\���� ۶C�1]_�K.:c/m���Vy�����g U������s7dΫia��WVr۲X��d\cڌ:+y�s�{Go�A	9��hVe�W�����6�yeG	������x^���Z�缌��Nz�u�5��1��_P\it��9ѳu�2�)�m�Ms��ӄ�.��@J�`5�%�I��^�'u_ �Guw]�y	�(N�Up@���+WKodw}�n�Q��;��GEq^fU�ug(��{O�p}w�nY}Ò�ݸ��4Ð.�o��ZG��v���>���.%Ok�9X�EҊ�x��l����{1���WP2p�����B3U�r��!|�^�@�E��(n���P ��WS�������X����mζ�^��v1��C5�&��e��u�J����YPZ+KX\��눻eԇ��\)ouq�([/;_ַo�K0�\�U�[��tC�w��leA�rM��|��&�r��5|�cr��5e�a��I��OM-]��O��2*�Z
"
	�C0�0�j�c�b,��������=====>>�>�<9�Ƃ���j2�(����1��ܓe�p�z�J	��"�(������=��====>?_G��g��������j"
 ���2f��.�
,��*)�L����k���oo�OOOOO����������YO ʊ���� ���1��sq��"�*"f���Z)(��w�,��0�/R0���
��"*J�����taKIIf�aUT5n뤕DRLДP㛫�"R���c���a�U�[:�ʊ�2ZF�"3	��nc�PPS}����#�bJ���2���!��*z�(
h
h�8)N�QD�ܘ���d�Ù��Rfa�f�4�CCTQ��GQ[4,��h�������&Y��s�5�
B��u��f����J��O=;0sЕ����9*Xĺ�5��9��A�wZ�3s�{M"�uf���.Kw��7_5�>�|
9�b'dp̀���-.��a*_	���Tr��-�i�{�M��_5u4�;��������;�w?�\��8S��tZ�m��G��^P�v���j`���0��-�@�)
�췯��Ĥ43'F�y>���� Q8��X��}�7#sm����l���-y"�V����P�� �{�Q���SV��.m�ع��fq��$q�{���ꄼu�)}�aT�O?8�A������H�Jbl� �â�^}zg�tPY3��7��XD�9-��&tK1��t����*c0�H��ꐮ���Eq����請�u�����ro��L./U�-�h��3�=��R�5 .0ء�dN�ч�u�n���L�A��R8��Y����,�NC�5�����å%g�j��|�� �V�����
|���u3`����������)@�㭺��>��]�x�����\���m��[=;*{D�`�s�h	bR�Xs_o%sF�b�P�}D����9V@̮���<�mܖ�b��{:
���R̆�a}�ؕ;E�J�}Y+��i�S����_V�e���y��#�A%�3��ol�;���**�+J�U�Z��oC>���}�>*�|��p9[|���=�6�tv,[XK9�<�����Q�f�z=ݛ[<�w�� �=�j��b�����_��'6��s�1W$�lq/����x��<���a��1zy�y�.q��1u��]^�~��Ӌ�f�K�e�OHMz�6ξ�s��|M7�&��i�=49�)�2= tNoT��u�=��Vw|��{��9!~QN3�ۨ�>�|�C(��Xl�t;����x��SN8	J�-�U���}V����{^�9ݱJ��g�j,Ŭ��\�����H�\է�OUbk1c�օ/����[�����9����cs Fɺ-S}�ܳ��7���p_6�tb�Cg�b{��,��QcX驼g7s&^��u�^��3�3�V�h������h���7[v�ѹY���r���݋��|�ػ�X*j3���h���+��Em����7^V��W;�K��!�U��K�S�;~�#n�Fʺ�˖���^�r�ļ������V[��J����X3]�k ������!�.��2Z�i�`]�+k)4	4�`�@�?W��[{��߹�(w�}��;���M�*���X[�+�x�JT�M�e��
:�Z�5{�u��P�^oՉ�:�q��y�s�y-:��8����8�Q��ySHOl
�	*�C����Y e��e�`��v�n�g�2�fxZl��p�PbdR�>��=�������ү��'V|[un$FS�į�jWra�^W��*���r��y��0�=}�]_jpݘ-�5�Dt��7�.�ω��wh]aQl�-�|W��lMo3gev�GI���]"�B�Jϕ_��u(��6g�R�Gc�6E\��i���<D���=϶�N���݃���.W��č��*޽I�������:���{'c�5��g���Q��u��YU�x��R��}
Ќ��Ѵ�:�/f���?+m�4��I��38��/����'h,-�J��6g˨�o(��� -e���^��Z��:]>J�g~���s��:ֲC��J����	���V�����s�>�Cۀ��v%�ȇ��q:�]�@�Ν�A�@2וaֶ��v��{��i헟��ӳ"�A,����4>��7�Rz�B��`f���ә�P&�=;�N��b�i"&�c�@�'s��U����7�����X|m5�_%���n0�<	����j�v�7-i
@� ����<à�V:��U9��ۛl��]����@G�s�]-���9��\�Q1!UD��[��zz'o�L�3=˨�2F�U��e�L�::�u>�j]���D�����UݹmH� ���mG��` �9�*i��vo��;��P&�����6\�X9KZ��t��a[!Z�.�j�;)G�m�IN�ad���N'7��?Ĺ�u��q)�Iθ�#"`ts�)s��|�<��5�L��4���8�ܮ9�]�ѷWG�����4�5X �y�0�z����z��I�v������r������]U�V���H��^񝚍�f�g&2~/*�~�+�/UnG����o%hkjPc��۫2�r�R���l�D��1�d�q��w������1ѡUc�Z*�R~Iw^ӝ[��!2��k�Y☭����x[�Y;c�]{�sxi�.A�Ω�;C� ���9��p��>�Ӊu'ǆ}�|CԖ<������Y����g6�x.*�/|�ճF�m�g���3f���<UoT!�/d�jY�G�h�-�ݩ+�e��XB��ԕe<����k���J'U
ت ����XR��v���-V'��������:gv"'w���#=�+� ���	���^wHГ��WV{��2��TEue�B݆cёR�!�mxIs�$c������^�뀯�2�r�LJH�o]����tz�� �/u�;����W�L-���46����;�[��et6�� ���܇һ�ưq-��`6���d$��y)�5����s5:9�;��e�1l������!2�C6۶r�f���W�g&��,��m��#�r��ݿy��ݳ�֟�-�M.�Ϙ��1�d�6��j�A*DM���T�zL81U���Y�� �M����2�.uy�:�fN�����چّ�8U�e�}�5��j�`�	1�bLİ[�dw~�}Y)���en.���f�W]u�=o����zz��Zj����5��a�PY@�m��.���dp,	l,���O�E�~躟Q�_Z6����g�p��]�k='B�xYL�6Z��L�g<)xwј�ܺe�-��-UXIb���0vf�<���bux	Ŵ̥�Wʿq�[��7}�Zaꏒ���G�D�/4��.�UЖ�R�z�܎7j�I�}�A=�����Ďu&��z��|�.��Gk�#^9+�T��*�9577J��0Gci�@i�ƪ�W�n&�t�����%���s�u݃��3�z���ۢ綸=�c��r8=�m���eV�sOTކ�Zٝ-H�Η:N`��~ːAY�y�>�2��~�{��e;f���5ѷ��+i������͠1-T
����p� �XG�1;���;��j��Fb�o?F��xadL�*��C�u%1�ˀG�%А��l�-�瞑[����rUn���7�^��F��P�
�	��2(�q^����k��{� ����W��Z�FҾ�Obh4%-=i���d*?�9������M��	6�p�׿N�+ �ӳ�������7�,*]քԓ�a��;�}F��%�o�E �$ŝ�e�� �ReW��,�H����b�oh�:�e�5d�ݲ��i�=+�$Y�zx�ˊ{ސZGyG�4��%���g�)�p���y"���P�1�j/c%���l��EEd��Aԋ�g�v��0VhA��a۽)�Z/
T������T�`z��f���OZ�J#z#N���u|@W>�.��h��0��L+��TЈF�R�M^�V��3x*�m��)�b���@آK�h�d_�_dt����*��/=�#g"���b�b�R�����iO�|n�gwns��jd>J�a��˓J�V I�X�ŐVJ������x"��E�8zm���d����O���e�G:��Jy�{�٢k��ӥ�/���[ )H����q��O]��'|�J��5,��ݵ�=�2��G&�����f�A�[AǐwjZ�&�!l�ڙ��|xq���.�v�-�Si$�VZ�5e�˽�X8�Х��|��>�֣g��c�o]�i6�y�����O3T��.����k��A^��.�+�2PЮ�u^��%�������f��r�`q��N�g6=]Ƶ��si<��d����7oPs�"�;ی��I�o\yڹ�bV�O�Kh�&���;��74�m{�}T����=�+z�T�ۀ���r���̭��!uuV�n(������o�ɔ}��m]ժ��Rԫ��v
��Ɩ�SF�o"�1Z��Y���;�c��pū(�e~�:���'/.�����g�6	�@�G��m�A�;xp^�B�=������aWm�s�DZ)-l�:�7X�a�R8Bj�����$�hd��lM�W^iE 7�T�-Uۈ���6���쓾_/ ��|�_4M��K,��2��Ûb]{��=��pZ~Rw���[����b�LM�`�3�v�/VJ�0�E��*<z�D@�:_�����|9�>�ǐ|5���4�F5������N�����W<�H��"�\������o"3(��H3����	�>v�B+.�Xǻ5^���o�%JLS)rN��y�Pd�1�m'��lV)w�D#�����ŪxwZ�V�'1��/&�����L�y^[�MS;h�b�ӹQ���Ԛ�-�k���⪝0�.�k����Ӹ]L� g^�����Gy�!C�ʍ�i B���24��N�����m%�^V"'�;J׏gŧ%vD�V�f�[X~�mU}d����V�Z|���Y�Z/p�٦�U��*�"c�R��b�Y�����(�61_�+�3%y�k�+E�NY?t�h��^>���ٽ&	J��e���1��m��tMlvg+�]y@ɼ��qxx5s��Q]����(�V��h]>��h��9(�w�s��[��Lcb����˦;5��{�e���}�.fc��z�A��f������yWp]632E�P���9^�6O	�g@��􈂍	vM�=ձ���U���j����#k:���	�Y|Lb��6����FP`ڢ��R��l�ᣏG� 7g'#7���/^�R9?�IY�� ۉ���[�Z�g�-����Z�9���IR�k�!�*�P��Y�G}Z޿�J�|�ߣq��/��{,����2�wwH�:��=��ؼZ�\���D,o |�����8f��Q����HRl�e\�#9۶�#��2�u6+z���j��x�9m��锊{���_���m�"�ّ^�*�"����n�	�q��3�����M��"�ڹ�I.�"���b�\/F!�����6������?VW���7��O�_����Ϊ6��(�Wd�8���XXs�ٳp���ɂ�RT�)+nz;�7�i>"�m��w����k7&8�ppF�Ϙ�̑�Ϸ��vh_c]��EG@Qj��[���dp�[ВCI~�Lǥ����@d&r��a]�B"�h\^/�yP��'��ҖNd��)���u2��s���"�4t�t��rK�V�c�^��;�+M��$�]�]�lmx`��oS�k3vJ���9}X�e�C�iJ����F����K�dTq�T8�0f�bj(��ؐ���ƥ�!�W������#����G^z�<����x�vo��i�Fsξe=�+�k���,���T�sE��ϴç{�W,��`�vh��ܮ�qӷF��]�;c��ݜ�*���|�}�ic��Gx�����+z��w��c�Z�t&�9^��>k���#���)&T{�Z�h�<�_ �dϯ���\�;̻�˝هy�1!���A�u:p��q(_�#��,u���!��[�N��E�lu�.�r���O��i�]ݧ���}�&K]�1�[��z�7�>�Y\k�=zӲ�C���>��ҋu���`�V����4Zٍ1OZ���Ix����Ǆ�Q�S���{��B�H�Ώ��i���uR%y,�W.쵑Zs��S���)�j�L!��cj��+�N1��tz�[�Ų�'�jX��r��t�o��m�^V��qs˹��mk�5}���s�hP�:���bR����;+5�lLQ�m�e�[Z��i��{7���3�F'�7�Ն���%ȋ[b�n��7�L��i�kng'�r]G�,B��$�ď�J
�|LWY��γ�q����r��a�c����B�ڛ��)�'Q�Dq)��z�J�Cj����ř��Y�@�"l�7�����rJ�ޫ梺H��t��q̘E�GG�������ddT����4͘�x#�W[|EJ�7!�vY����bN��V���NF�;���O:�3� t�}G�����8�V`�d�w+�7�ա��G�ͱ�bں\��>�jI��n6�޲M_\�=rL���2�`���j���:�^0����C�9�g���g���ûN��51��*�r�ª�
�]�\��<9Y�Ufa��<��c��ݙS�֋�f,+�[�T�r�۹���X��BJU���=L��ۼ�,���J�";|A95\�5�d'����@&.�����l�U��4X��;�4@ą�"q�Nwfc�S�}���a����>�ow�}�����R�s�i��С��m��o<!:���̼�z�Z;�>��04�wp�U�s���v�)�B�na��&�tݎ��wKX�K���!�r��7��\���`M�_�o:�Շ�il�JK"\�wi����S9^C��v
�{�NeI3�Lµ���P�RWVw��̳;CUe��b�zi��%���Q�&�(�WP{�{X/��!���G�P�����x�>�)�gÕN(V��2�Ю���Ȧ�BI�v�Kx���z5X\����5����j���9jWvf"z��]vx�����*b�w�k�t�^�0Y��r���c�q��oF� �'��۱�%qH�����+Q�'y�z%���ε���C-wi�d�"9ڨ��홎�u/_v��m��T�� g<WE=�wLe�9݆����K�ݷ�f�.ި���NZ��vB�4>�MT�4`�������L��ѻƣ2��,��jq��Y��p�{�vG%>��8l�� �*L

��@@R��G��.H|�4k� ��,@�������l&��R�m2�4���yT\����〆i�6�V�d|J�@
�IL ¦"�yu�9�ϲ��=B�0�=�b{�%��(���l�+�0�h�$��/��8���ǧ��������}fyȪ��QQ)AKE'-�$�r2��[,)��8������������}}fy���#��pr2��L��)c�:�2�rr���)����oo�OOOOO�����3�����=�*%��K�3r��=� ))�̡��a�w3c+�,�>��6(�s�2��!�C#"��mQ�1)*��"��ȳ
��A�l�&]YHm�SO��f4�4Y�ff|��I��b('�`��6���h�r���ɂ)"
B�C#{�\�&
�#�ɠ���r�"�J��2z� ��s�3�2����H��ZfC� )+�� ���6�)�������a�d�uX�JWvP;�9-R�MRSCU@Q �;�	�	�I�o1wd��)���,{�in�Cn]�����k�	j�g�8I�Κ	�DR�`����S�F��o�ciS�F`�N���t�3�D�@Qa�E6�)R-0���e����'��i�E�t��8�C��t���	,�^Y��m0%�t6�:Ƈ��S�sl�4lf���Cz+�z�i��%Q�C���< ��G4���.º�+0�p��4�6=]~���Z��K�c#�a
���ޟ>�)�[AkigfO���Y#%��U3���8U��-�/R; *���n��;w�}U~�У�/�VX��GY��|9-���q�WۯÜ��HV��d���=�
��>�c�0����F`-2ǬȵG���[���
��W2�/�sN�}:j����o�
Xя�^�U�6׬;uu�7�wZ߹�ٽ���@�%�2��l`�D�5��%w�,��Y���eMo6&��&�AyK�h�u���";x*�l�M2��<fU��7T�Pc���\_,B.�DMѺ����m!>WjI�*d�3�.wj�Uѡ�*"�?e7h@Y�a,�Fs�kZ�gh��1eΗ�7`����.�Me�Cu��Q�������J���`*[�bY�]�/R���O�Öw���:��H]w{�d�������T��D 5�P]��Hr���c�WՈ������n�о�J�7�]?�%޻�@֘@u(��h�hb�j�����j�+O��< y��A6� l����jW(�Zޯ[���,nY$����,�tE�Y\�=R�$H�L�r��sb�T�{Ӏ?3��`�Q~{a;�໳B<��k3��ϻ��'MY��n֣V�2w�{�VK�[��pv��-�."B�Ѵ ���3$Ma��b��]yY=6�����v����UFg`]j���,Y��Ux����ށ�{����p� �{"�K�C�<\	�٩��US�A!v᜾e�)���	E�WoHt�I.���­n�����9�u
�g1a�uH�C�3eb1��3�Zr������~�&�6#A���a0[��Z��x8�b�Vdq"��Py*=�M�l��ePl���t��p���Q�B@�-���1��ţq����"���v�Ք���V&;Yk���BX/�?��΅�Y�܃y-��O�(8�U�7��{�GHV�^����̮�Z��kmV�Ȓ5E9�n���m���ht��}L=���f�>����8{g:�"��Vq�rF������"�*�q9g��j���^��](�_VF�>di��-%��{Lv���f��5�+ `�d-%ء�ZJ
:�/ra���ka����Z�t��m� �p9Os*�\���G\h����sy����DNh/I�YOݞ����#�.�4�9�U��d;_VhSM�`��ՑX�ɯx�kP�S�uU�߷]a/(���,��L��3wl�_�]�{��ay����U5�~��Τ������*x?��~�{n;i��`@�@.d���r�7!�z|�4���ɮ�B��[<�KW�ٍ�K�udIB�d�wUf�H��]���a��줅�wi�|���L9����K,qK��W�w���7,7E	Ɯ~�³���9��z�C��c��&�`�p6�-0�4���٪�������_�4T<GL��.ݡM�%����G��������k?}{/��K-�ھ��u)U�+r.��-wp��fR49����K�W(�Q��µ�ޠ#���;�B�ιYR՜|�;;WQ%�f���5��[�/P<�K��p���5"�Űue�]��1{�1��.�
c�����60��w�c%�U�>m����: �]"9q��L���&il�{�N��Y���vImG0�b��f��i�~�;���;	��i+A�r;y�0��6�;�h�M���2N���F!;<3a���,��HxB�T�[�lI���%�������eǶK���A���ioG�׍�t᭡�<��wU��N[�S� �{��W���wi�<�O@l��r�BX	��&��&2��7{5�I�zB�#%���q�yl/��x�#�<7gd�4��/����^h2��5��p��-���Df(��'ع��W:e;��7Y	�/t�d�2��4e��y��V�wH����=w�'5Tڇ��&��n;%�0��\�^�5�KD.{sZU@=��ç	�Փ.�=y�����X,%[l�
AT��NNR�}�z�F4M�9��8�u��H�3�9��~\����T�B[��(��;�eSM�m�9Aj�8���K>wQ��+��i�ߌ�8^��Dzɱ�NtV�[8�}�B��廋%�+�����e�݃�1{�Z9��WRٹ�A��}��5̽�C�4�UY�g$����!#�{�&!к�B��F/C�����ysy�+-�'U#p�m��]b������qN
!�<A=W�Y�lNh9D�����=�v}�0��pZ�}���E�/N�k�GCԤU�ȸǯl�0�k�0��ш���%a�vҀ��Љ͆�Qs�>ޭ��y#��'�ܽ�����ej��<�f����o��ms?I���49�Ⱇl�#��K������l��k��衯�;�#f�׮ަ��|K��w���D��GKn�*#2��.k��vK��\��&�:tG�fϫy:�R]�oΖ�rf�oYw�n뜷/8{YST����E��8�t>R�z�1tz �.��>�+>��X�[����֊A"���bS> ��e�����;��u���mHl�uݷ����"��� �V�ZH2��h2^�k�����f�a���1��j|�=%H�~��_����5���0ʟ;�XU�Y�̬k��H/��Ӵ����r�d��s������j�N���'p����L)��wf��)�?q��i��{m�w�=CS��]lӔ-s�`:iU�w}�/&�r_<ʒ��Nʭ+d�<DL�y�$C�_�{��h��,v1�"��
�������it�R��\��3�0�"���r[Q4H�X��p.zq�c��3��ƹ�P���5U�tfoA��WP�c�m��R�;�C�m���I�>�2�GZ֍�Ƨz��/W�%G��q�U99|$/K�c=9���+��~��e�Y���i�?s�F���e��Q!j��4E6R޵�i񃡘�۳USm+r$�.ȒrtWl�Ͷ}Lx_��7n���
v�������6�GE*̥Ͽg),Iq4ig:�ꬠ�eO�l�@b�M\�*+�]��-��ޞ��fk���:%+����`7kP,*�ݩk|*��z����VE�L�.3{O��C9l��"Z�VB����Q#���cʟ��!SM�y���]eY^��>�,=]��!f���E�@�	����e�=��04��;��$�nW�y����n!�N!@htlXV( �r�5��&,�X�E+��w�K�2(oQX4��vh��Y�/i����T/��Ty�zLY�h�x���9uu�x��c��r<������V��Oc�D���9��p������NN�{%��Զ�~��n��E�w��	j[��Kl�D�:����Y��^O��T���Xv�ُ��#�j����{�֊ɭ�YT"/���Z��L��]���|{l���|������q�G�.ؗ�g:`������]ϛ� w��U�l�;�~��p����ڳ�$KF���ŝ��73.�,ȵH;3�!� ���_Us`�q��S��;@�cA�o�Ƈ"rSQ/�/kO(@G�L��,Z�D��͡���^�b.��9[�,^��U4rvl����M&2cȃJ}|k�1�S>_vP��E9x32n�+/Z�CC���'ٚ�<��`OS��&﮼.��O1��~v�eNq������/N<�`�\нٕ�I�`��;G�WO���DND	���q.{��7��j3�nٹ<ps�6r|M�����Kkz�<Ӎ�z�ܹ��aw30)��ry��v.��M�ܵ����ypDYA����,}�ܟZ}G~�n�ufZ�z�R��et&V�c�;fV]�x�t�����0NTX��)�)��&�Z�������w���<�J��^�n�N��.pfZo��>�H��.qM���+��x�}��5�����{Wp�\7i\�bmd����V�^l%��.61VO���/
+?fM�ap��v�ՉE�}D���V%�c�M�u���Y+�G�v�lr�afi%s������F�#3��7�!WD�L5/D�-�H{`�Q-�)�Ŧ(ɬgʞ�zrw����~YvA7���9�x	X �=k;6W>b�qb�E_.ʨL_ȑ5t�N$"Q�`��[<Y������`1��?-�f˴���Fe��"&lf/��ʽW�3��]�raI�b�+�F�= �0(C>� 6�Qy�2R���^�:��ݮco���F�׫W��D�Lwf�8}�������3�헣[��\"+��!���>�>�O��|��Ɖ�8�ы����3�Ӥ�E��FW���׏s+�C�+�''�������5u��8�p����䪙P,��`�!����@����&-�h �T8��\��\��<��O;�ݎ����Y7	p�Go�vCb�*�����!WR����h�7.�u�bֻ䛮�f��dSZ��V�X��!;�K$ �pX���%Hz�u����� _	/���CDa+T�ë-ݺ�誋3zz�4����g5S��؅��F�!�;.��; ���}�;���a�����fcla~��U/ܟ2�ؓ{� ���L��i��cl4"��V��g�V��ew�/�Y���$h�Q%�1P��EF*f���	�l,�pS���2E7<E�b�j'{$���z�<ՠ���5����g����]m����U1!Y�WêO�MN����%�H��s�!f�����]�fD�w��y�5���)��p�*��� � V܎5(J�nk4^�v̘����b1�e��d)�4u�$�Z��@`��Do�8]�&��̙��,�z�nY&���8��Us�ב@И�S�Q��kV���
ʋ���rP�n� d��pU�yWe��n�n���[��ǝJ�106k��CM\����s���%���=�����Wi��g��p֟�~k2Mrx��x�)��e��k]��M 3wƗ�� �>30�_r:���]���
�ژ���=�z���w~~��|â8�q��	eU����'�70-�r���+rR�٦��)��b���
��fb�3I�;�[��s�0�8�Ț��}[�"������~�1n����syw�T&����sHC�챷��i�ɂ�9Ft��+�BY�� �w䐙��
�������Z�b�.�ݳ�^�a�N��5oEx�	‱��f��_��@�����kD�J���4D���˄�={f��{r�=y�)я��Vz�ؒ��WQ5u�-M�ͨ�y���]>��=^������=��D+8��x��r��8nB��DwU;b�o-$P¨��a��\퉞��N�Or3Ji��+�����3���l�s���N�W>*٠�d�3g^A���5���7�NdJO�3r��~+���U�fw�}Y|�����Ed��5EZ���۶G��?CY��df^��3��1�d�5ZVe�*.�Oj����@��r.I/�mE6�{�h7E�P-o_��#k���Ľ]�>m�Um];n�+�e��Ҳ��Ew��I���ĳ��!W�~���]���q͏�;������=�zxtj!����7HX��Z;(W9j���}}IZ=.�-<HV#~�r�xw��<5�Iٹ^���U��U�;����zŔn��뭌������������-%qb�v�M�,P5�3�*�����n��NC9�Բ`ڄ8j�f���^u�̙bv>�v�Y��L���U��˰8, 5�4n�ۃ�'� f�x�A��{*���q�$��۫yٽ�J�]xT*R�u�+_e���m�����˟^���G�9����j�:8h�2��n�}�E�oC��I!����4V�@�ʑ��U��!G�r�eQ�]ճE1*���R�Wv*p�t��X��TE؜�%��1ಟffM�"|S�
+�.�Cr�0;��*U�n�AR]c�4�c�S]D�ud+C�ٹ�y��/�x��3������V�6rrInZ�]u�y���GFS�h]��7v�%m�����Uଅp��R:Ȇ 
�m\��q��Ew �uK������K�_�(v2ծ�g!�xr�#�8s�����G�rR#��B�r�*Y3�k��][c[���9�i{k�����!�6�9�\�9t�k�!��A9d6�V��2=YBC`si����93��(�1��իb]k���2ӗdzP�f3P.�+I
�W$?qQ������ph���,��7E�W��+�B�,��!}�`Է��Pb9=v^2�Ԗ���gf:�2h�z�>�#U��ZV��B��Y��\��y�>��K�t�w6�2ՇRʞ^�;���7Xj}�7��^�����탱��-Ă<z�N�(El
�N"_J�X��8C�-�8�j�p�gj�k|��v�e���rw��!fޭh9����Ub��J�<Z7]��[.�=�g+�eK4b}�]�q���Z���[s��t�#��.��������a͆^�I��+%I�������en-�< �n�z��2�p����9��>=+;�o�yL�G�l@f�Z�q</g�٤�`E�җq��]
Q�i�z�*�XV��)��������Mԥ��K��n�>�J�.P�K�7^��E�n�^+RA�T�!W`ȣ��33)skU�C8���v�
Lju���㻺c���4�~r��X��9ָ.�%�.4;���1��լ���T��z��[s�yӥ�Z(��%=�k�N�����b��U��e�Eg�]1%]���,w�6����ؒ˫�}h��nV��\hx�
��"�=G4�G:q5hP Z�t������i���J��3�����S̰	oUٍ�av>�0�c���Y��p.����y�Z&�ohCC�����K9���]Ǝn�=�8�s�����]܄�:C�� N]G��5�NL�X���,�>�uT.�ƭ�hj��&Z(�g$bP����%5U���zz{}zzzzz~?�3����+ؠ}�j�*��+}�a��&�|�7
22*����2��G~?�����__�8�}x����2��ZJ������r�v(&�2ZZvW�8ν=���===>�������rV�Z_}���((6�-�,��&H^fA�dPr�
�����	��X�w�Q�z��`)iiF��-M&�
���C �iJX�:���gXui9]���EE% P�E�9A�KM&A�FN!T4��@��9�e�E�h9HRncKAu��R9u��F���d�Y5^c�J�q��)����qԙ��r4�[u�m�l�CN�HS���re�r��2
B����MPHQ�ُ�Wo9�����±Sz9�9ۙ�n��J)l��X޹b������S�ғ�Z�
n��v�@����!c��B���j_v��=�_ۘ�����V��[>b�M[���̫����rnE�J^��9��[��~�ڮ��3^�`��+ �R�����p��HE��/��W&��w��<ҽ��<��*:�ev.����������}3�b2#�������aoa���,��@��W�i���o'"B)/8�EּSra���\i�i)��}@u�]��}�~��p�i������Qh=8�()�ۆu�[�a�*��]�E�M]�9ï�������xY��<Ͱ=�(؊�j2׮���i�Z�k�8vư���gO0ӛ}��/{`�-�;٬��y��hΦǗjB������ux�㉐)8v1��z���27��4]��0>�4�vr��y��w�̹*�o���^����C��{E���b5�1vv�����bY���i
�Ksꕈ82�^�Ǘq�$��e|���I�́�=q���I|�\\t���C�(#1ڼ+k!�=����*��^ues�M��=�b�V��r���_nR���B!yc�kɱ�y�<��z�i��T9�V��W�'���w�祷�1�uh:��0P5��`4�u
��Sݒo�-�YT�׶�U��R��|<��0$\�V+7��H����]WskǼ�׺R?~��x��g|�`c��ѵ�.F�f�i����>������|T��oUF�N�z�y���v�������J�#1�mO��D�lyVNo���&��_3�bEוB�|g���7�|tǳ:=.fq�㒶���e�*��U��t7h�ub�C���e�}y g� ��ѹ�(�[�k�Y\R�؜M���2�r���M=tgcf5(C�`׺`B����d8����n���CL�/�*:m�'P�����
Wv�P�������vZp+�gw��LW^�:���جʴM@k��2RIcC�ce֍ڎ��V��\T>��^���y9�0����T�֘l�'{w��H��wb��֏E�8��3��?<)y�\�>����c�h�.�bX9�vtqږ��J�gj��%�R��jN����楅w�B(��VtWU�.�.Ů��tDI�]��@gWvs���Z��,�=O�
��7�@�;&�S�:��$�:t2J.�@�ְU��$,�b�U�yf���M�E��~�_2�2�m�
���p~�T���4F2�N����\��m	S=00rK�Y�����vB2"���"��k>����#x�0�QR�׮ndTM��)���B���\�ܘub�=�k�=�����T��f����T�v��Mi�}!Gi���aӮ&<gW[R��W8_0���u�ք�@�b;����-���+x��tK�V��SY�m��������NSf����be�t6�=�]�"�T�>���q��ݞ޻���Tϖ��'x��T� �2�l�x�1/P�x��>7��r�u��I5����P+<B�	��	�����Xf_V��ʙ�Sӻ[��5���nKΰq�{��Ư�d(��ˮ>Ӌv�&۴�Mۓ���w9� >�l����pU�}W)8�[��0oJ[�o%���J'�~��Gk���9FU����Y.A������ūq��BE�����������J߯{��r��J���y�|�q�إ	��1�1��|:ե|z�V��F5�0�δ�Vɛ���mk�y*�F�ا�������S����wut�3�����m� ��hY��i�iK788���)���]Y���<o����cJqk���Wy wT���Ѧ���R�h6B�a&�T<q��[��hɠa���s��a.�%�B�'��X�Y�Z����f�ꛞ~{�K۸f7ݺ79+��g�-�D�ӸW
�9OJ�������®�i{�T	y�T��S-5��ky:Kt�u�M�+2��wn�s�^�->��G��U鞇�3�F-�[�������w �2��fܑSlJd�ى�̹����]���I���r�χ���k�f#�y�����6��F�i�pn��4�H��HϪXn��m����4�-�c�����ܽz������K7�>ga���m�<�mֽ;e�x�ے�΃q�Q�}�C/o�x��\�W�s���\c��
�v=����2�Ha��*�T�5I��1���j֗�[��v��=��-�pZ���T�TĶ�Vg+�QwZ��R�WF��sO�u;�(�s�:�qÖ�j��M*r9�*?�W���:��Ǜ�N�G��\��8��"���{·��$M����DM��Z�Se��yB(\�Οf)�L�t�6�w3g���ւ�����ј����G$_r(d�,�P�MM�3��.�,�2W8�r�].g�Y�a������e�����i��f6Ƥ���Emmέ�]��}M�� eP�><��t-$6�Ռ��CIh�}�DA��f�����7�Ue�(�~��k(���Z�;���ю7��M�1��|x8��T6O<%�,ۋ0�d���J��,�z'bq#2���e�����); v�ed�D�+�KdUM3`-I�5�5P���xU����٧.����<F��Q]�Z��M�I{��uM���K��t��x���A~ܺuƛ���gOK%�[q�Z���v�ӽQ1ۊ��ʋ4�u�ϔx�z�B�Z�n5��^�p�u���Ց+��]�8:�SMhp�9�6���x����f>�+z��X���|5�W��|:��X�@�և���7�hT�綕Y�Ƣם�uC.xI��^(��a7ι���}ׄ��qT���K�K�]��`��oJ�}�(�
�pfhl����ɢ�*�>.Ko2��v�$�B�pw��>�k�$l��U��j�ᚢ�L+eɍ�W^�ӕg�'�W�R^�T�����9��c���l�Ŝ�wx�b�m�]t��-i�u ܶs�N��1��~Us��.Dl\���;��T>_�i�A�"ֳ�F��n$л�10��0��lOV�kB-v�F����Ϣo�ʦ|���q�7�nJ.���zoE����u6��ӳ�>|J���.q�eJ�Bb��=��>�}Xj�(f���:����_�GKac�.��1X�|=���LWO	�{������K�.��'�k$su�V,w>�M��qW7 �jl������:��ܭ��W��q�J���m�*�e�W�M�n�+��V+�5&3�Ψ�
�_ô �FF�{����K,qK�⬠��\�N�����SJ�q�c`cӘXT5�A�u!6��J���ۜ.�����x*��7���P.���Kߘ̜�+D� ��t�[���K6�L����G�3�A��J�-c�yi�c��%��׻J�TFw�|\ *�o��V�4��i��Nw�2�H�t4Q���4e���]���x<L��4}�W��e'%��"�y�O<��u�4h�ә�e�������sW��D�`WEz�j�k��i��𺺷�I�{䊤U����-ܔN*�������&5o.��`OVQ����MF����ޏ]�s���w%`2��I e��y�K24��>0rr�1��`_A��R�=vM.0i��V{��_؋I���kw>�ev��~�4 �T�v�GC��Q*�qֹ���f���i{3|Lv��]���g̑��j�6�}r���/��5��kh����e��Cld���.}4�׾+��6�Gl^ڿe��.�t3DmnpOݯ(fd�L�wP!����<7.C�͢}w;eȸa���D�X_
Yn�MI�nq�Xc�f�kt�Ēgp�oxuF���'����p(���*�q7^?��\/GZN�m;MV���NJ-e,;��1�Y�b�k�nsu;�\	Yx��X\;Y�?ǝ�wgL-f'>,כw��g"Y]�bi�"{��b�Z9��u����0���˝˶��-��2��uV�����ʸ3���w����d(7wW�T�2�0��Eb�j=L�e�;u����=�ͻ�����-��]MJ*(�縭��'+˰i/��9�c���|߻�2��m��[����5\��Ӫ�Ѭ5W
�5gd�P����}M�7Fq�+�
�����pfA����뤩i�rne�VĆ������n���1����q�>Ń�8ޝ�S���I[9�Qe���tx;7P������k�*ʥ�|��]d{��7�8��lq�)��+q�j��Y��}{����*�`�{c֋F���q��ҳP�#[�:��]�(���9C�FSWW��^R�~3*�v��"�O�T�4��TY.v���J�����SU�Z�6tnƳ�� �P��OR�f������Y��p����yyv���a�`lH�k�B��e��F�B@��D0άJ� s���mL��D4Yͭw���Xo�Z�y2vk:��x�}�l��"�<6�R��?J��뾸7��nk�O�ތvu6U��]6����+�x�5O�T���9�&�#� �������;�3���h(�΢UW����m>_We�5=�n��"ye1�-㽬����ۮ��_i�c3q�+�okEk����Oct��^�l1�Fy�c�St/Մ�G5]Ts	ɡ�/>��Տ�m�.���^So�˚���v��s�gˮg5��w��vD,&�x�����M�1:K���i�N��m@�`+c�.�l�ě	I$K;����xTf���n���]G;��l�&���:�h�rwӰe�
�MM�c��Ns�@�����@��LuLO)j���ر�{ض��Lv���E%3��a���~���V��l��]��F�]W�x��K%m�r�V_���g���Hk�j<��;4�Ow��gm�k��Epܬ$���0��Բ|�4,��	fg��ek�k,�_L:gaӪ}�����"/��yg�P݉P]�G<$��rn<j�PD��	���~΃�f;�C�䴝�"�k�����5���Ύs������v� ��AA���\��M��x��"�5w�;A����d����fXF}��F�h&duӎ� E�	�u�����RӼ�7��Y�5nԧ�"�j����Kȩi�!�
�&T��ʗ���q��fV�}�KѴ�.���1H�:;#�܍�yW�*����u���Ѯ�c�D7^���ډ/�͐V���o�E���{���2���Z
���O?Q�~��H'�;+mwwU-�4�&���e���%��f�Q\���YjA�β6I�'w�B�-	͟c��
�yf�g�k�T�o�Ut�m'޲t̵��X�e ����Ed���=;ᐧ+.���{�7�a6�>na4�x�u�D�ߨ�n����dѺ���#,�"�qi�h8�4�]��L�a�jz��U������Kw�'��خg��k4�~S>�ٕ��F���U'~�[5��$|�܄i�����6y�k���ՠgS7N�=�⩻�:�h�N��z��5tTu
�Dqђ
dV�y��e��x���"�շ�O�?��[�_�~f#�\��Q�'���� ��((#�ݡ�� �O�YP7x+�ʄ! ��2�B$4 ��C(0��¤!"2!"P¤�C ��Ȍ4�,�"�L��!"���B��l�D��!�
��'R���B��!��� ����t�B���� �H���B���B���@b!���
@�
B��"B��
H����!(�B(!"�C@��B ��J ��!�@�� �"H ��@���J �J �h! ,!"��C@Ȅ!
��B	B�4�f"�@��$!
�(B�B���M�HB$!(!(���B�@$! ���C@�$!"��B!
�ʄ!"�3"C@�$! ��"B�@"C@�'�;���w�<�_�*(� �
�0��v����$��^k��l5Ҧռ0csLX�;w�y�������������TQ��( 
���������?�?�/����8� $��B�����B��-W��	��3��HE�g�pDT�	VaB D�!�I`(�$ RQ!`R eB!$IP�D�D!�D��IYP�$�!A ID��H$R �H	D� Q�Hd�I	�%%�H%T�B@�H�E)VF�a�d�fA�a$�b�@J�Z �䐂��J�� � �*H��R!H��B�B�ʅB�H�@$Ȅ�A
@$��0�2	"@$�!$�@@$!�L�a��X?�����I�j���P� �4��_���������?���@��><� 
��*��LQ���w� o�1vt@ƧH^�C���z��O�� ���_�C�����������#��*�?����C�оh``�����:w>���( 
���w�B� ����P/9���y�ï������~�����C��" ������W����)?���)�����߁����.��=O�BO���W��`����� 0��������9��Ȫ�/��0?O}�(������o�_���O��PVI��t�p�@��` �����������U�T(��ب))�(E@Im�H
�RT�$���EPI*�)J*�����
���RɊ$�DM6�l�[T̂�2�ĥ�Y�ڒd[5���5�l��S-�Ř
Kk4JڃF���X�[E�6aV�U�֥��i�V�C6e�)kcVJ��Z�پƝ+m�JU���lj��fR�6��l���JK6��ښ�D%�1��b����b�i��UU��Z�ɛ[e��E4�U[f��i10�veUS��H�p  -ה�T�N�u7:҆���+�ɮ��X�ۺ���`�)]�ۣN�V�]�9
��jj�]��n�]�Nja�ηWmv���p�]����wA�F��4�[5%����l�� sB��С@(w���)B�
(���z 
(4<�ۏ;�
{mn�s8i3]���tVWl�m]�[�)�C��Z��i��uаw��@ݶs�����.$ن6̘�fk&��o  �էC�Cv9����N�Y�ӧi[������we˴�u�c.�ӮΚ�n�t��WwP��n۸;�+GCL�k�۶�'V���Z�>���H6Ʃ�M��"�  ׅ�h+Q���k�j�,��0�:��v*A�[q v���\�M[��Lt[���n�jOa���֛�p:յ�F�E��+k[l��  x���N�p�۪�ح�S@;uW53
���sN���ۆwt���n���w�k�-î�E���C����u��[�UU���)%J�ҶfW� �4�E��t�N�\��)��-�T4wu�T�[UJ��*�[��*�u�u�i������SZ(��vMw1].�aR�dU
4�F�hd���  c�{6�K\�WT}�7T(�w�j��U
��tP��ކ������P��4��\��))*a���
IWr�QT�{m��U�U��m�6�R%�  u�>�Hi�w��R����3�T�*ާt*P^�={�i����T���z&:�$Dm�yTBVƽv8tR�T�w��Pwz4�%d��1��mU�  3�|��)+�Sמ���U[�o���{׏TP)�{�T��ާ��@��y�z��$+�X8����={�JAm�WsҔ�T��喊6��ƭ���*E���  9��٥�=��B�y�=�	"(^���Vq��'w�ׇ��EW��7(�E(�ך�U���׮yUJUI�{��BR�)�S�)JT � Oh�JJ�2�E?&�mT���@�O��E  5O�4Ԫ(� 	4�h5U2 j~�����"?��7.�?���(�Q~���5�lw��=����5���^\o[ͣ�!I7����!I6HI$�����$���BI��!I�B~����D=���?A���"�YUv�l�U��Z ���Gr*ݷey�70T��O��)/hR˕�)B�lGM�Y0]ն��y)�lR����wu� l �i+dS�.�^\Iۆ���)%��n�Z�rL����V$mn2T���xU��KLug<��Z��f�v8K�7!Cv�����V ˻���z�/�p@>qfb���l����Kȋw���/fj��6�lj�1��[Filnn��z�Ј�%��JU�]�6�e�$5������z�ʄy��N�dt�[n[�ZP�"�Y��C6Z�#��0�r��OU̲m�3*��,R�B�.��kMXZh��wi^�����ţ��B��tv-��e���X�k�+
��3������QCh=`a"͍�@A=�fc[p՟��ZV$�!�
Z�Z�aRR������'��>٪
�&<T�]̍PG^���seS�2�k�[��Z4(��ftK���)MR+��٫����Fr�N�F��]�T�ncU�n ���pnc��	f�Ø��r�r8�Kˠ-��oa7� �|+"�b�{SK�u�l�B��V�9YJ��A�u72���h����0�Y)�[J�ƒЩ�s(�8�Q��͡Rnf�!�urc�ƭh2��V�`䠎|�V�5�dR��YD���Ҙ`r�`9��E*���*\ܥ� Պ� a�Z�ìn�m6���Y �B �PVNA[�Q�Wj`^����f��.Lʓ4��)P�Me��#)�YA��!:r�B���me˻�w۪�VF�a�pl�:� �ͻY�t���tLu�wu�2�$2��X��b�W����1̊�d'�MK/2�;>�Bun���U<�kba�[aP���׍f��E��Jc0PbPFԬ�a�NH���]��
D��c�!�Zf�Դ����B�1�x��j�Y��,R۩�u��ȗ{�s1ӥ���K�N�5�S,�9R�A���;��5�Pm�$J�,�/6�Sw��L!�6��z�Ut���b?G�i<m3w��Y�����ո��ԃ��1�a1b�lb��j:��4�ͩ���CEU��K����X�.dv3pec&U�����!��P:�bҥAa3%7�*�ll��4سB�S��l�3j��U#N��DĪ[77卩�r�/HS7]f� �5���ՒlN���
�e+�j�X�۹�jC&�tY��/Y��P��l��o`�A�����Vof��!p���XӑL����*yY!��e�4nT���F�۠UiE�;>�
�9��ˊ��Y�J�V�ݸ1s\�MelRi���JY��6�U*�.��v�(��BƘnՉ�6��N�;�Y�1�͡�/X�֪��**���;�'���{4ҳ�h�wC	�@i�`W��=ؠt.|���$kn!RȒ�n ��LN��h�W5�(kf�a��Jٳ� �0��fS��`���;Ku*u���%�i�A�=���bbu�]eŬk�i!4�����ˤ]�+TJ����xsw�л�1:;�mnڻF�cf��T/C��̘;Q�L���Y�cnU�lc1)��t�@��5ұ�p��o�A����i��6�lp�@@�Vo,!�D2���Al�xr������t�P��@av�+�KA7e�ϣ5�%:7GC2
,���#�u^���d-�(�V�`�4�(�����e����r�f�$��j�A�VbMJZ�Ҭ�Zd�ig�ܰ�]�Ų��}���$zے��Bf%QL�B���l�E-�NF� fDhJ���'�\hʿ�i��U�ӻ�A��m3���N�&��@��ܻ
�Tm�����2�jfQ7�,`aM6��hLt�VM̅�m�8����Y ѮJN��T�*�a��L���aB���yXD��6!G{-�Z���jmXC3s.�6):V�%f�Rn�y�+/T+�Jff�k����l��۴���J�ܻ[-mmè��A�)5h%@Q��(-��mn�U��&�7�Z+&`۽V滭�#4�l3�6�3S�
s
o1�n	z���2�H�12nмM��"Gb�w�E8�&��U�J�1��-�-\ܱn����2���A]���t
�P�F�X
{JbR;��f�Y�z�M�t@<9X�X��[��<%�F*'���Y�HW�e��t�SM�se�m�6��\9p��锵�lf[F���2�e�r���("LUCD�f��'.�-ρN� қ$`��B�.����[�p�W{1X@,��ckmأ���i�:�Pz�73st] �UK�RE1��)B[pfL��=��G����H���#�����{A�6���;�7�jX�[Cb�j���4�H�Z�.��KR�����a+�F̨,X�OF^۶�ł�6��h����GN`ˀ+���$�6���!+��S�V�Dnd6R� i⸨��*��*����S6EK2��[�
�dq�Grчe��*s!a�)VFVZU&f����n��-��4����BQ��0�.��]b
�P�G 8���ʘҳd��$X�c2��$e5f%F�7f�qO���!��Z]H��XA���Ss/J���(
��eD�)һ��+��b�v>��Ad �r�+�Sց94 С�L�p�wF�ɹX*�!�v�4wB��/>�Qi�.�JޥJ���h�z�f3����Y�GF3N�:P����ڌ@��t�)=�&�H3�ie�ܭ�����j]����b�(6�V9�SN���/f'{x�4��{�5T�a(�݀���p�����%ǫ6�T.�*3��ܶ��Cwp2Dj����4,̉�,�v�!���r��.���i�[����ޢ�u,�[Q�{�YҬ�5�mF�(�J`W{vrR$�N��F���-7ic;B;����$��j;[�2��@e9q[1[���ң�r"mL�Ri3ͽ \��M����a�U�iT�07&K��G&U��k
%��)����V^��֫��L��mēT���܀��t�Xf��-S��26�ln�RwAR1Vkn�kCD;o^��śG9�V��Z����qy9�(�K��֞S�MjyCSf6,A�.�.�s\�`�Br�M#eܫ��<�sE+���ѵ��:4���5(f���OE�� 06 %��xl�L��VkR]nR�)�8b�CDH:
�d5pєE��R[9$��i�F��$Չ��&�Ȉ�j�M8ki:�\Pf�p���JX��"ѱf�аr��	��Ќ��X�#���Q���ul�nJ!3�X�&^"v�>�Ԡ3R�z@X@����*[ESI�f�yv��6
N�����fU���])�c�)�7Ra��nL�b�ǣ�
Y��H��!V�r�J��u�sf�V4l��Z�T[@���J�h�5�8q����j��eb�oi5��kC���Xïv5�7�f��X��,�����ќF�5�@��0���d���HѰ��i$�n��DR�Vm2�37f�K�luՂ�J���ۡaK��c��[Rh��%Ql�*�K������f��.�*2'��W����1�M�4 �f�o��3	�^�j��*d��I0(⢝ձ=�46��ڽѶ�M�p�%ynʽ�����vh��o�hA�d+�Vd���S�
J��2��el�H�E�Y��	g!OhM ީ� ��5J�{�)ȍf^]ȫ]h) �Si��uh5tohڤw^U�L��x�1�G/3�[�zUc�5�[���>��,����f�j�	�Of\%�
�.i�q	vr�X�\T#�-'�a��p����(򆽭��8���[J��sRY#`�V`���Ӛ�У��:��h��x����f����Z���q�KN���*Ε	(S��M����J6~D�A� k5�vޝ��:�7v��m���B5�L��ɮ�;ut��@i*�ۘɲ�k�����K��x���ִ��,�XWZ��-���@��-9�:N5�n�{�Q���ؤ�������˭�r�Y.cK
+IH������+1�Yn�f��4��D��R���v.P���3�wM����$p�}�̰��J{!i�o!� �:SSڰ��ۗ�n�
�h�.��nљZiX��M�p+�)CFE,��ε>⻻4E;�B�7� �&��Z�U�[XS-f�{�Zv�h�u����@aUwv�X�E&����ATwt���A����D�l�lzH�f$��`��&�E�-R�Ƣ��:�iņ�@N$�MP�X�J��
g1��Y�E��v�@�+9G/B[���Th��6�@���Yw��W���*����bc�1�z0]�]��e�u8o;�]:Y�Q��oK���
8�B��t隻?ekt�1�r��`�l��j�fXh�4m,��JD*�v��Z��Qf�Z�� �.��Ѭ؁�R���lf�eY�&GM�t&	bWZ���D� \���KG"���#q<�4^
�M卥��M�.#������[�Y��\.�!J� �H�%dtQ�Wڏ2m#�Oflv�v)BCW��U�ղ���"�@v0�WEbu���5w���V�*$6�2�ɌVJv�1��s.�0�Hn�U+PصPqY�\Lǚ��rk��$L�^LDX/0�Y�mM�1�A3��ݳ�P,y��;j��,�{#��&�n���.��A���Bȣqn����{n�)ϖ�A�`j����f�@��r戨Mʴ0�v�Խ������JdQ5��,0-�X��;�ce;�Ԇ6��%[jC/�UL��W��Y��Q,��6��f$wGP
ٕ��R Xd�ʆ�2���Kh;{B�i���Nz�^i��9���%�В�L4�5e����"�.�l֝ӎ��kZ�M���������=D��%�W1j���Q11˨�b)��q�r��y��m&k7�N�z�<b��EH����t��&�1z2�3��J?MKng���"4��)k��wGlHp��hV��{����6�y,3�����Y�<90��
��r�+@ݭ�9��d�TfF�
�M�!�h��30؁���Hh8�n�R�,6]ژr���5D����G[5bt���v�\�mS�b�b��˨�\wE����ؗB���q[*&�X��p3[XS�L�n��1n�HyX(K��*Y-莬%��V3�J��cͼRn�e8���g�A�36R��)b�u�v���4��D�+q�WGE���N��M�vZ;s!��;�67�5i�c��k%E�hhVӣ��K/�%n�M�L{+!q�m��oE�M��^���m+2©�k��w35pq`�R�8R��:�p �:jA��0�{��7VlPxأ�(�7teB2#A�&��A��K%�̰���-�s�.��l�imK�b���ı�ҽ�ğ�a��ɬ	v(� $��'s�Ø#t(����@�i�|��ߖ�[r�W���f��U��\ʕ�k,���2�3L?��H}�sQ�uiUգh����R�UˠC�),Q�`*je\R6�*
4�P��B�o m��8�5�p�)��ַ*T4�2�20<da1|mSƵ�!fd��l���$�a�T�
w+�Ճ1S.�K[�XCV����$qJ�Ћ3m�[����
Ha�V�B�m�κ�5��W����r�̚��(#,�V6�A���p1�DGE^��m֧�����{z���
si��ݕ�x5aQf=��a�����5A�����O3t4Ӭ��+�"Ô
s	�3)�p��,�_ej��r˧L�y�IE�jhjm�W��X������̛30�(K��!�p�TV�bu�l	����y*ΧR��ʤi㣖ѨB`�Qխ�dn��m��Eo�J�C3:�,H�"�"�C����0B��K("#�����[���CE��8��)�V6?�`���y�!WD�Rd�a��ز�̼z�����[a%���;W�v��LV�M����
��ϑv+"�{��Ж𕵫n�%�-q}�;���z��歋~���5���j��k�U%=�*�	��=�9[Y�M��J��˨�)G�1�u�i,u�p��2��G4�M��-�+(�5�٢�-K1Sc2؊5On�%{M#W��+�ᛃV�:���a4�Rr5zr^��@7��2E����,ְE�,:�"�����E�C�1k��qn��$bT�зr Ӹtu
��-I�L6֡t�HG� z�U�JW6�(�eA����=B��WW����u�V�Y`*iU�N�����[��e��:s��Ye3�#Gt(��^��QE��d�m���P��{Ck�62ɴ�1��z��Z��7M��	5�1mԘ�q[r����ˌ%BV�����-X�v���u�c�JUˑإ�X1�+7U�.�@栯3C�Z̛�����/
i��@�8���CY�h배"5�,}�r�B�Y���"�VƦ�[����j���W+C[y.�6%�mF+MʵGI�4 퍦��ʰP�8/`�p������(� ��:�]=h ��7v�8pȞɱ�k.��+ 'u�ܬ��؝�[�#�Ur��)ޥ v-J6� �47V<�V�K�A)n�7�;b|�ɭ *����//��B�8� ���l�y"�0�ik����u���R��]")]J�N�[C-	�^�yqV�$0�(e4H=�j��)}���>����ECi�
�g麤�yH�1�oiIQ���	)�4���⼡�����?�ԏXU�cu\�I����S"л�i�K��p�8��7������܀R��R,:& ����0�N�e�Թ�;)`��֐�_=n��s�)��>�R�k�T�ؓm�쪺�Uԓm��s��\�e��S���ٮw�۱nZ���`�f�x4�.�ѱ_3n��=�_+�-ۇ���9�-#�#�_\ײ��x:ROh�!��S6q�卺���e���p	��âԂMw0<K?*Y�-�^�X��vn�����=�@�mq�½�&�aVI�z��y���1){��,�Ι��ݽ��g��v�.�^{��E�һ��r��JKrw�h�D�]���q&�=cn�euk$����V;o Kҝp�L�x�1���T�6�0����{���i��9wn�egv]��qXB1���W|�2P��l�����^@9LD=�����@m�76�5.0uw'28oU�,T�2�)6�J�mm�yxԬ�����v��Lulݭa��+��@�W�1��*����(]����zP���8,.=N�r}�VѰ�;���Xw�"W��h+���gf>�F�rf�e��1'k��ˏw�BEEڊ��/�=\��M�yRb�mݬ���Kq�J21�q������a���Z#.���aϴt��rk
��v(ǵ�e8�Eۯ�Zϴv3f��O{��TLnQ<v��8��>�R�s�a���2=�rA��6�\;`EF���PګoH���ʙ�\�;g)[ud�49.�Th,�$��m�Q��6�N�Y�r�1�e3J��\�t�'�F�s{�;�y�hi����#���Ȯ���Iȣ����+�_
?��	w9�J�Ol&"�����o�}��e=�]��7��2՘�6 �]��E�A	�(w3�� �����N]��m�{A�|�`S��V=��K��7����swV�$�W3�A��	�����n	S(�V���>�����MQ���wR��M��db&�N����sѴ��X�A�wv�{������N���]�R=9+B��&�[�[oi{p��Z��3�%ݝӐ8�[ݼ�F<�@� #��I�A��;H����79؁X�!s��~u7L�Q*�W�`�w�\v�E�Jpu�=m#��ys���,髒�UjVz9���Cɶ_0id�.%ְks�;c<w4��!����IG�
�c��jB4!T�rr�Z�/�����" �'rG��"R9�-�J��k��o9�S�㈿��
�
SR���^���Ҧ!�c�P��7�V���[�Mp)=�k3�+����tu��Pq�:R�M��j�
�K	JK�6O������K��x�5���>f�Z�#����dWӤϙz��l�8zm�&4��2*Hjr�y��dZW�d�z�6>$4�-Ɗ�~᪲}�FK�$�Fь����>iK�ըˡ�t�uN�qD���Y�ׄȵ�'VwU���V�\2u坉�VA���Dᗂ�8Ӊ��'�����k�Q��ܷD����b��[v��ͫ9:�����5n��[ւ]�g���k+8u`er��c���M��.;ù�{��E�k��Sр"�I����@���EVȱ����^�_u���5g�7x�,샺v��&�)�/�ᶷ�`�3iS�ݵ��P�J�()�\Q����ݝW�{�?�Zi�������h9�TU�Xz^doR��]�٧Y�˨m��q�׽ �f�Σ&�&NFڥN�C�Ev9(H9�K1���iD:9�j����n���,ÐC ���oΈ�R�2�˓Mb2��܌O�f�be��.���'5{0�AD�z�]���39h@�훂�Y�e�}|\lN�\Z���Е��/5�nk����qaͽ����K��į�W\G�
ɠl�p��eq�V��j��µ�Ch���LL؂�U��pl������l�����H��M=�����8)K�K��
��`�!�_^�<4U
��G-=���Б������^�ccc%�-�`te��5�3L.����u����kX�jc��B+��E��l���ũ���k
�t)�k�.�ȸ*c�̾,��qu3vQM�z�p�[u��s���p��o@!,Y����̱QR�n�;�c3U*o,	����k��	ک�.�����N]`/��[�2���T]�:��%�1�y�	2n�H%3\�sr�h�e<}���<Tb�}r-�ՎN��('u0>�!V�pc�C�V�Z�5�[��r2p�N���F9³	"���SN��GY�[���Fv�O�^�b�ΰ��G9�ay;(�4��:Gټo׾��V����?�����Ą[�f��μ��{C�/�ش�k�t����C��ᯞ��M "[���1�ք+�;G���zE� ��J�#�+yMe���x��ʷ�#U^�3{�d}�9Eh1[O0�}\�H.��ؓ��#�����A�b�չs�ЙCX���a;��ڧN�F12�]�؛*Alz[(�O�W���3�r�� c뽎Y��
�n�T���6��K��]��:׶[Iq�Gr���H��lv_6�
���T=���5��d��9׼��ZS��r��A]�Qi�}��vuΜ�˔Ǧ��p�߷:]��cL�*g#�ć	W�o��4F^��m�[����:� p�U� A���N�T���D�Cq�i"��V+E�\>p�E50Y������O+��q�兽�-��/�Y@�%͈�ߑ�֫�e�Hй��m�c�����]����d�#n�*�k}�vj�:*z/,Eoj6쬷�#�	����Y�B��5~>�.�1Ѐ�yJsc��G��%�ȡ�2��8~骲���ʽ���9K1l߲���!3E�-�#��
��)���+-�&����f$��82B��ՖEW�}2[[�dn:���0^'QsZrv��Go.�i�oC���ۧ�ɺ�\swN.�ESo6m�*Oq4�������߄�{1�\#�h#����)�+]yR�$�=;%�	����7%�u`$4�l��(u��1��dҤT�$3t�s]J5�%)���es��I��W҂�r#����$n1�<S8U83���CJ�ք,���k�r*�Ȅ�d��Ͷ�m��ڪ˝V�5[O;N;t0��F�!���/rr�:��{W�6�8��)n�Ó,����v�"��i�Q��]�"l���*�p�z)r�~�}0�E�ҶgV˦,�v5L�o�P|��0`9}�V驼2^�M}�8�=�2�.J����]^����]7H��������{r��W�1�th�
߽���Ud��#Z��A1z���!�=�WB�(�*����otn�%D L��;��׮�\V�!�9��c�s<��6hIQ;LC�lwN�pR��譾��h2���B�_�wV�������<���yצ�|��0sp�V�N)Y�i��f*�Df����:V��;)���n.�s�ҫ[�؜�x�)�M^8uka4ޝV�q��z˂Q��گx��3���;+8�b��w�f��Ge��O��Ѯ��"�.�:۵ݳ���v�s�o�:�լʾ�#��@C�b	Y�][�9f�Ц,PBu�m�D����m7�|'ךU^9'LMdV�xkJ"�D�e�y��ب[�D0'@��ʒ�=F��+{�f�;r_A�=��jN�B��JU�ݨ�Wt���"�j�.��X���j9}���X��F��p��6���T�De�H��.�339-�[�^n�ۯ���ru���o�����%��tu}��KWU�և#kr��AᇮsY�	�]U��#ܸyu'0��JP�]�3]o3Ȭ�ݐ��������Xt�iT�Lm�b�n�;�;q�����dT3NS�K®t���w�E�&Ǒi2�A�ۢQB\|�RH��3�y��Y�JA.���9o(3���IԳ��-�#m�;�H�h�_l9^���Z��Fz$�1�Yk���X~�su[����ָ���*N_V��7k)P�y��0�b7J�܏���)���7c!��6���{YWl=�/�Z�'�B�G��9�Mu���C��U�k���݌Q�85d��\G��o%K�9ĉF,�7lR�h|���!�����B'��8�wu��{%]�`�%����d��R��3�e�w�=e�!@�*�W<��AZ���3W ֊+��o�	����%���f;\ȞqY,���e�85���,ӏ/�U_3�L0��nM�[���ܦt���-�+l�Kꋶ�0E*��47Zt�\z�^I�wO�X�;��X�"h�;"!ͤo�(��fu���b�R���gma�uu�N�څ4d����"7;8�|��m��vτc��$�WM�xƂ5;n��JG+	�iJ�\�9yU.^'��!|t 73�P�b�����t�i�ʻ�ԩ{�d1h�U�`9�K��k����kY�MV=�Jky-gS�留��L�WVWk��*V�X(M����y2�s�����vL�\X:m�G�{�@�Euz����E�}B�!�7�v��$[�Q��1��";څ��K�ۗ���'T�`�C��7%e,�o��:Oe�w1�"o�\j����,_�@��@�`�oP�C.��6
��0��17j!�8��̾e���}K�w�J����eB�FM�Y��Ђ��]�v��3s�S��J͹����[̂��ZW��*�s�&��+\{c=�r9��ƌ���T=VȖ`���0ȕ0��䮮b>�b�[[|��f�K�P����s!��Yz�w�7���\qX��Fr�k�z����gs��9L$l��aҖ��\�$r��2�����F:v�N��v��l:ƈ9f�n��]����a��&������j�5'S��:��qi�'�	Z�ì��"�����򂤮�`*�>��p��'�H�P@rn��*�[�x7Q�=����ک�8AW�;�F�c���ê�*�pě=[�s5�̾�Bђ5��B��2DR�%8����T{�`&5�h��Ln�jJ?P*�$D�>����a�JM}R�Ķ�2�7�C��1uK4d��lݚV/���n�o����2&N��8�̨�jx��2�A���VE\����חf�-��y;�Jz�+c���c��>;�¸�h�t���ѝ����iѶ	������}���6ӒRAn�=��b�6�٤m�8k��/$��GL������R�kQoM�PTF��v��B���v��4$h�x�.��47h5�}	n�Ͱt��ʢ.���2���N"쐮���;���]��YᲵpW׹Zɶ9��;�B��F́��c�G��p���Kh0�XQ����5��/]�n���KB��<DPYyI���O��L�*e��x�s�BtC2]��^Bi�WM\h�θ�y,��y���
��ɚ�.[5�6�!�^�&�H���Uq��3��b��毕�yZ�]���U�P]t�^�LÊN���!����>�����R:�歾�)v(SŔ��?N�Y��a��T���GQ��_]��sF,��R��1�r�N^�����LIɖ�H�b2A��<�����B�/{):�l�S10޲�p%��x�0h/��<�����͘��7l�ɯ.��R�p�_CMvt)��"n�(��!���b�[�Wk��/UZ���-����ݨ��9��m��r6��X:� �e&��|���6�rܼ�Wi:��8����v;s�ufMGF�NS��g�.�R����f�jCB�Pi���*��awvK�sJ�@Es���Yv���[d]ç0r-�z���sX�	a��Р��V�1��ޫ�d��ʂ3:Qb��G3hD	��En��HP��%r߯��5No}3"���Du��+̂HH.�)r�3�b>�}`f�̨Žwty!]���R����F޹���W������x�������ݶC����p?mE�C�6�=
K�Q���+��7�$�C!����s{���\,=L�Jf��i���[y����+��2;��A�q��s��n<��ǒStU���Sڭt0��A#�"��0�7|�lO�_CQg ��}�;���J�]u�|�`��w�qSu�S(A�Ha���t�<����4��T��_&֛2|�>��u�]�t��b�!����ѭiM�N����&[6�C��b�C��lo���'��rN�p�mHR��:�]]�wf2&�.ܫ��@�03w&gA(�iǏ�$��|���a97� ZK���x�X� �8���;�$�%�B���q:��cT��Og�~���RĬE�n����z^t���y��:`h��+�f�#E��<3cQ�Kn#��]�jU{�^0�o�Ƞ2SK&>���0㶹�7z{>Z]f�b�mx���#۶�kW����[�C���}��w����l��W��~oN�+raﻣ��Ԩ1�&�Y�k+�ܗ�c�<5�E=3�|>�{%�)Q��l��j]SVe=]K2�����hm�p�o��\v��I�0�Z4�f���*}Ȼ��y�2�N軩�B�э�]��
���Q�WC�&3>;��Yqة� 5�2���k0�;��N�Ŏ� Z;'+�Z�`g���q.O��8���\�j�[*^[�ۥVbv�y��-��9VgH.��R#�<
��,�f��&����me�K��+�I�>'�H��tj����z�&s!��Qn^9�2 �j�������*>P���7��bA��Y�%R9n})�������i�V�49�n���m�C���MG\�t�.�Eŗ��]P����S�����t-P�:�Ef�ئ�FlڗL�j�����}���?(!	&s���<�9����3��nӭ��M+���	Z����f��-7F<b�8nn���]Hi�њ�SX��8ep}��p����:���J�r�}`�[�r�'Р&�(%Z&���|
��w��d6)+��|P���u���\�n�d+��Q\�Y*p����E�[�sp)���%�_7��_'�{��R]�����%Nw���wjL�{�Q�Bl�rٮ�/�\��Ms��U��e0�nsΘx��a�Mx��5�%Dʽ<mu#������_*[�XuWc7c�
�h��e徱��dZ߱Z��[PM�v�wG���Mt9=U0ؾ�9k�;J\]p�Ag'(��]�1q
�{+-�\IL<q ��E˽ٛ�����Y/1r�� ��۽'���<�
�]�,y[�ɬj�WLs���aU];vkJ�f́�++�͍�徤0�Na�c�0o�����Li]�h�����9���͝l���G+�16��{}+��Ol��FT��=Yl�Ūp2����@N�vm���Rq�S�0ݙ�	R_d��3���˸�ȃt؆��#G.6�I��N���]rD�ޘ�eLL,JE�ۚi��k�ဓ��*;o2���wV�C�2�w7��IѲ���d�N��1ag'ݺb��2��B.��7:�<>9�"ޙ�b�Ƌ�����'���y����+	m1��bA���Dt�c��p�ǇP~�*kxK��T�;j���0r�"#t�����|"���
�9ik�p����:�ѺT�w \N����Q�@�Y[�ߞ@��/5V���w���H-O�/1[�y���Q��0gA)L��������٬�la�F���\m����\{��Նbm,i�_X��)��#u�yZȵ�7��;���Թ^�
�`�nP�+wk�{zNdvP�\B���ܱ�X��r�6V�*�,e_D�U����[.,C�d�K�C8�	j�T;5ے�����[��T�W5PW�:8�6ޫ�F(��P�;�� �w��.:�j�ے3r�2���7]nY��k9�(�J]q��xEk��C.�V\��1�D�dEm�,�\��Ŷ�Ԏ�F�k�q�+V��o-X�!�Q��7,���>�܅���U�jò�TO����Z��mຘ�6©����f��^ ��\49�P���Nu�1k���vn�{�@�,0v�.�/�:�����
��w�8�=�-�Q�U�/�JR���5�m�Cp�Wg����-����-�j[��9���b���7�g*[��k��+�Y(��@��%B<�-���W���"�b���<��J�7]��;ٝK��"����#Y&�ݬ��}��;$NW�G	�K\�궥.\;2�B�"��^$���E� ��F��[��-�쌚[�!b���J��˔ƌ�S�و>�dS}XeE�pϨ ��X��Mݩ�q%�sF�攺�����ׅ*�u��lC�P��2�#wlh^�M>�pH�YF��厐JMD�oHk�ѰMB�OK&�V昊��Z�ʄ]Y%�c��s��]�|����H�"_k�Ɍ���i�S������k@k���L����h�vt]Βhu��$�s5Ǉ�`����01[�Ù�ݔs.1Ru�"����z�"�|�`���A�[������q�:y�eevL4�]�w#r�&^�՜�WY\=|tɫ�t�2,�N� U��G>
�����7g�%K.�͇�Y��Z�n���*���iYE��ŵ}ڈG� 9��S�v�*�y]Xi1��2!�V�^ܔ��+%{�a�3n`�Wi.+t��<�-'W�:�ЎO+R{�n��3O'"��y3Wu�6:d�zxƾm�H�2�eifܘ�@b}N� ��D�fF`t��wn�З3��&�5�ڵ�@�B/�r*ʰLɜ��a�N���9��u�n���͌�7�0�V[9�N�:�77f2oX�'��/wd���)���F�N�T���֧��|�L�S��Ŗ/0��Cw	5}�9I��ө��*֒.�H��yA��e�7t��N)��G�, VqѶc�<bǙ�K�]�n@�T���
]JWD�-�n�����îr�r��e$��`^�F�i)n
���j�����p#N�֒���U�siY�/r���[�bA�wx�\;b�R�*ޅp�B�yK79%w�y�]���R�=�̈�����C��HU�K9
7����.^1�:4a��(<]yr.Sv�c��#�i\kK����07p��%��θ9�䲦V�ɹ�Vj���Q��Y����s��N�yz�"�e_B9�g�o����� ֕�Lԕ�<��!���С�+;�z^�
�B�iw1+98�c9��a�*�6�7�w����FiAܶ����'=.�so�)��)+�N����J,��.d'��յQ�h���>�+gc�j�PJs�iUb���Ŝe�\��W�� Gf֡/q�]�1]�w�����Rq��N�0���OEi����[f�����b��1LiߔWΠ2�&��NE.�{���7�wV���I.v�+s�#�̝�@k�iP �]��~��46��Y"M�H��iz�=���F&��(�[7�4Tۭ.�抲$\;��0a��S*��Ae�B���h���fS�7�9�wid�@FeҼ/e�1�.������ ��踖��}u��E��>��it�L�*����M��	�j^h*L�n+�+DΥ��\M*�ŋo�殮�K�|��o8]�w2�)5M���d�Z����DF|���ȶ��"�1v�V,�iY|V�i{9EWA�1j���@3bM{�ro*r��Fjc��I���lZ����>w�X�Ln��Mm�`���=4�dY��vD�%�ù�x������5��W4ȯD* ��1#��Ija��s3h��O(����FlΤ��Թ�P4Rg1S��W4��Z�Թz�Y�{�Cn�����O�u�Z+h۶�^pbf�q���u�n����:B��3�GW��f��:FmU]&85Ϯ�N���7�6S��	O"�<y6�Æ_э\�.��mbz[=���m�NЪ�+Q�`�n*K��Bē�$@���t��X��j�U̇�\�ص�܇��xݔ���[�7�?Z�f������k�N���'+�]q�6�w,�\Լ�iem�S�8jh,ִ�R�]l3��Q;N����n�ς{��`�ŢF�)�2�����V�eK�Kޑ��R�d��j������0j�+^�IC�L�&���Wj_A7�a#K�eެ���**��%�X��t��i��ٸ�vk͜Vtmq���5�ח-
�"Fq t�2�ك
�,++���������8����KҖQ�]s�a�M6Fve��X��k�c-ء�TM�1����w�1��Qy�C�i:j=Kko)��I�zPKW8;�!P�pv�f��X^�H�&	vN6�.��X���m.X/�k囂�G����h���[Wjt���e^�}��W7*e]�n�5���l�����6B�^S���<��Ugs˝t���sЫ�L��	Y���P�^�-�;_Rd(�E,���4�����Vi�G���6�Y��w�8E�b��):�!� ;*�u�z�
�����sx�������4H�Kh�&�']���1��z�dJ�Fr� �f]㾚.�ix�= .�wW�].���pBw���ю�ܬ69Ja�d��`��)���&�O�+�%��ٙa�7;a�j����Mt#�{�/j��}�N�ס.9Y�ҳ_r j��0mLim������z�S ����D��tjqs&�/xۻLb�V!O�6�A�%h�ЎA@��)ł���m�J\�XH�*J `op,9��6,��@����\-���a�Nѣ��X�λ�%ҔYO�IkOPJ[�Oe1�^X�]WR��b��Ng4Dᝮ�l�gT��P���m.L��Wo�Ÿp��[�F)�H��f��V[6�ګ9���ڱ�0 �4j!��8�m�B���(%&hǻ�M۩r�I�x���dن��׍��X�_]�l�tWk*^k{�OvlV�%a�@�
"�E��[W�@�ж���o��{�-Դ�����t*u��pJ���+�(UCzV�����K���q��2�{U�/����!Q�ic���!��']�;ͻ�l�4:��a�/�x���.�R:ޫ���zdյ���v�p�p.��J�K����ZY������$�e���|nf��d�cڃ���PҾ����W�\����fHH�-����fN�w0����������+#���;`�
6fʰ��t�A':2�$M����u��:��O�Ļ��Gv����(�H�DBxq�b�L�%�	jq̩��v#���L1@v��F�:�C&�MJ(Q�1��i �u��g��/����z�&�xEn�]���It���t���9���I!�G6����څ-���(,��ʥC����8��TY�ť�n����Jm�b�t��ϊe>:��}Z����r��i���E����U�j�*��Y���ڛv�MV�SX�.�L帲���\�)t��6dx��H� ևͨ*X�6,ZM[0rZLhbW�К�i��l��.ʽ@2�,Ͳ��1��n5�S���νv(n��^R��sq17)�Gg:�x��ãөBԴ�{���H{F��hƸ��y�3�-	�먁6�5:�.7f4�����6��٠�ypR���o6<�쑔t6�*h-.�ڵ^TI��ka�{]�ָ���K�|�.�*fm�z�F�t&���&��vK�e�[P�<X�t���*�q�ݝGPFJ{N�-iS0�݃�lO~�����:�P��,��V�H����O
[�5m++��iJ�|U���]e������8K"mj⁝p#���WWٴ�-�6�9MM�x�Uw.�b��K�J���]���}��ob4��-��I^���^�����ל5��s�k,t����� Q�/oH嚤´,R����S�h�V�N.��+^t֎f�M�������r�1	QI�z�hv�xe>k�Q�������*�&A�e�S�Fv�������w�:���ϔ�����j�U�2��E7���<����4�C+!�Ǻ�܂]���r/�eGe��BŴ+k���)))�uw�tVw{��V���Y؎��mG�k:�v�e9��YI#;�V�F>u֓�Z����V7&V'r�f����-������\�Ss���u�6�1ڹk�;�V�]��] �.�rч�j��!�X�1���1X�7�w��]1� �ѕ[ǹ	�zK�fe��iؒ��o��n�xV��y/a^A&�y0I�U�ۺ�	��B�ɓ/B`�(Q�P�kS�{.�e��".�o"�Z 7�>;�7h�*P(�l9�]��㏭q��R�2q��*㿘;E�V�Z�t&صO9��]�͙ד�Dˤ����5������aP)=-�z���E9�U�`��HBx���ȅ%2\c;��3�/m�f�+��B�-�{f���va�j��r�b�N�:9�+��Ѝ��r���,v3��C�55���,��b���;{�2ƝΧP��]�h�뻜ʭtP'֔A�	n�=q�-j�ǩw}�'�W�L���(��	�U(��B�a�d�����=�V�}�$7�_�l��Ya6ʊ�e�WB��0�y&���pG�s�VV�q@Nwս:�ٙK����"%�]�y���+w��v��rt<>O��WYl��n�{����VwMRR��|��B�+pj�3OLۚ�C�E�Z5�� ^Q6�V)�7.F�����[f�`*��ݰmusB��z${J��<�����.��y+(�P�7 �YM���,ղ�dɏh����z��c燑ʚ���+0g1�STs/�jno;�jY�%��@�wy4�2���#�nļ�Z�"n��@t��'*����-+���v�%��ѿc'�Ak�m���Ɏ���:�[��ӴKw��� �5��z�a��q�iݽ¤�`�+L��p�i������TC��8>;.vg-}�Rym.�6	i�3���P^hs�+��Z��m��k%�ut�w0t<�Z]M_7�V$ج��T�$:�͠���GE��l�QA�-V�>:+��>�7��C8Ɨ�n�V��P\���G�qn�7�������q�����[�*�e@T�⎸ƥ�\ApF�����2}������gNl�f5yn��G����5-�x�_V����o����|ݢ	�v1�V��#�+N�+U5�Uj)��o�K�2�tSX[����)�V�?Sq_���N&��أY{a^����WIW�.�]Y�i�7{�뒊�E�{�Ou�ٵ�kn�Eַ;��x��t�[HS�ag�`0#��G RwG܈�VB`����UEY��6����pP�Z�8U�%'Y�����/+0�s�=�O#,gॣU��v�
�Ҥ.Pt�rg
8,�C�+���t)�l��;�d�Qm\�4���:+��i�˨��;]�x}�����n*c�DV	Vp6��n;�������*�&���h$�x�5�)������4S)�9/.��B6�Ƹ�fTr3���{%3v�g����Λ��N|ʕ���X`t-�Z"�mݺ�&媖�aީ���S�t�%��6����d2���t�C����Y{M���.�9G��;�����M%�T�u{t���]<\9\����
]<!��1:�B�h�׮�-g6�^V�"[t�h#v/hV�U�L�KyL�i�I{Ў k{�(�k=�.����{��n���!I=�������V�k$y��Hڧ@��B�4�,K,��f>�(�[��U,s�6���u���j�U�[��2n��m���!�8ꕊ�S+�Z+��mV�
-�K)�-X�*K4p{��,Fh��GnE�Fk�;A���V�9^�I�Y.�uGsL޹�
Fx�
���J�)�"E�O���,WO[��4㎥M���kM��nh+����K�t>|�"���C6MЭZ���le�T����ܹ<f�.4�R��ʖ����6M,�ox*���{���,�]�݁^�S�m8�"G{�-��-������v�Y_�٣�6�I�	R ��C�,��:
[�rη��o/�x@VWLgЦ)���T�õ�-n��[9�c���4Q�Ꙩ��YxE�43�\v��^�₮�N*nS�5;��}/���T���E�f��Wki�XB<h��hQ�.��s��θ���#�X��Q$��U���S�\X�����+���:Fu3���{ІT�y5%�u����ѧ8�>��y����Z�N�53�,Z�ޢ�:J}x��P�>���xt,���� �.�L�̙2!"�������ޣM�٘)b'.H%3�O\z�>�0l�����I[ �q�sI�}��ū���g/-�-��$b��8�`DfW��e:﮼�����QAulX��TY_D�eb��Hc(��Y�Y*T�
�VږЩX(�-P���2�J��m� �� ��e��R#EH�ԕ�²
�T)��E$Y�LV!W(fX�,�f\���Lh�cIR,*bJȶՐ��Yam������kT�Da�&2��,�1�Ԩ�3(\���AA`���(E��T�Ud�V-aY(��R�%Ɔ1a1f �R)�TY
ʁPR�VT����\d�+�**�&0���0��dYX�m�XW��� ����A@QH)��,RDf51(��1�
h
�PPU�̷��Y*�m�($P�I�{{�ܦvx���b� HҸWWp���kC�ᚸ9��gmÔ���0�[�L�j�龓@���|�M���%��L��v{����"~�S��`	5_܂�����!�cMG��*7���h��iC�"_OXW��f���%��� 1�����*�_�9������J�j5�Y�i�H�9e�}9��'/��M�쓅�v�"\��F��Ӓ� �1,Xc*-oݴqxblfZ2�[�i��*G�3|]��ϳ��f+�Q8+�m�ǔl�&j�^�^<��.~�{uz�o�{'��u���5��LwZ�c!���E��n��y�hgބ�4py!����Fsj�Ӭ��{*,!�Pc�r:�e�%/k����U}��>v]���ǎ��}�c�MΝrp=���0B�9F�IC��@W�P�v�;����A�w��4K74��ot;p��=�o��m�Ok��]Ta�6f}qf1��ˁ�B��Nޛ�&��[�%�)4���7,h�ޓ�oUp�pM��<�괸�{|�oP�YxM@�U�ճ��U
e�R�H�1��F����g��qJ�H�*���|�W����=��}�}�-��㫜�{K�4���������0v��C�&ak�م�Ņ��G/!��^m��=���$N�mќ�{��׹���i���j�%gq�/�ǖ���d�qN�|����Z\�S�U׿�J]�4+�n��h2�Ԯ
s�Uc1�Ӽ��lUx��ا5Z�Tx8�s��
�a|�g��r��4���uF�*O|�P�A|�H��Td�c;^kS�tw�*�x�ܞ�S�_6��|'�� Ʉ��1����'h�4��J���č���]�f�, G]P���4!��$S�@�d:r��]�KS����޹Qz�d�6'�t���@sj�ͨ�ډ�n�{va)�l���2v�e����o���6�ހ"�RF%I�P�0X����Q�73�@VY$ޭzg$;����ooi���/���'~��:�5`W���P�'�>�tkl��gK�J뢋�W�oB�XWp�A���x�S�_{L\�J���mEZ2#�ˡ���n����r�l��j�z(#Z�:M0��(=�PФ9��mP��W��U`"�|��A�[VcbjgX�v�sGn�N"]}�r�v��N���L gKq6�f8�n�H��j���c�_�ξ��?^ق�׬ʿk�ԵVY�S ���U��C�ٮ�����#����@�����0�)mr|x���;�v��c�Fb>��7پhٵښ��ݽH���h��u�3#��"�W�lFiA���<
"���2�&�-l��e.�ҢL�\����Y�n�r����%]���}lY��dȜ�,e�޺�Ch��'#�J��uuJ��J����4��^.���l�G�	f|�p������.��7��^m*��a���5���qC�s���ۉ�8#Es�#t�Z�F#�?�'g���U�	S3FR�8�yY�)s��&4|��O/e3�P��w��������+��s��n�����ǎ����*Z�Uvb`��A�S0*Ӵ��9�|s!�>'�b����?\c(��nG
�Sݫ"�.���F�r��W�S�x?�\7׏�𚗅�`>��r��S�[��db�љ�_Kq9#'H�=B{�%�ed�<��*K&��̪ͯ�e��]�S(���,�f�_m��N�K��b�.��.�e�0'^K�x����=�AE�}��:�.n����%���t�{Y�oT��.�6��o-]�`�H\T<��L�*_�v��n��[��5|�a�ٔ\��)�ty��r,��t@�O-��P�^

��.{���oP�3���W</��B��ňb����[�Ȃlw��ʫ_�%9?"�q��v^K�ܝ�\�AV��No�}�3}�w{z����2�^k\���G�|V�KN���j��-y��њ���v��,F�� Q��qw��5�r\fwnr�ލ�����T�Y�xwhNE��� ��Ql�}�e���!��袋o�IW'����*�Q���ރP펡d!˝[)ˡ=6#�i��K�ݖ��i� ߦ���"�Ro<vպ�Z�??Gc
�i��)�2!�Ԁ����]n������������|�.B��^<�*��[�3]��r�ChO+�M�b��4&6���[����Ӥ2�B8\7U�mu5	�T1��VH�+�6\�n;���r.Ն�u+M�>�.�eP̕�}5��ә҆�O��T�h�b�8/�r��2#�������ǆ�Z�凂����'��tuK�(��#p��ȼ�΍��K F��l��*����Y'�Vp\d�!_b�1��~� ��*zc΍�O/�g�u�`�^t�ͮ֝rp�ٌ�£���_E��72�+ِ��ڥ�ӱ�pˊu���;M-O %�|�LşLPў�t_(��RQY�]	��K���E����%/!hY��i&G7;}��j�[�t�5ԇ)�"6Ӣ)\H���`�Tg�ˬ���ECW[��c�z���8�V��EѮ�fY">/p���)C~5��o���hV��F}�:[��Y첩
՛��*${以�}\Z�.ѼӶ�,��S	u�AU�
�S�tP�A5L�3��;��7@p�H���������Ւ�ܣ���\w�_��r-���iB&N��QK�2 ʐlUH��U �N��w��r���z�fq�Pt`U��c>h*�r4��i����%�3R,(F��gU��%5{����	̮=�3WDd�׳��1��O'����9�e�D�)D�Z���oZ�_y�|�>Dw|�$,�1o�NC@A��܆�e��� ��y�{$x�3پA�� z�`�G�{U���V3ƅΧi�<[Bx׏GWh���8����͠�Ss�E(������者��_p���G?��"��3�r}H����L�眺zf�D��'L6Z 6W��E����Ӓ�>7LF��kJ߸��
A��d^��d�甡�e�_G<��Q��<������ ��c~;,lH3Ab�R�z��ʱ�!ZtH���5����yT�� ��'Y��Yx'�&�z\�I��dƧI�777g���s�XZX�p�ؤu������@�yL���_��|B>�g���3c�ɣ�X/V
2-���q�%(ALL�_x��g��W����y�W�N���.�C���`i'^�nIǣi����Ԉ���-h��P�fG��2�*\o:V-���l_d6��vm�K��B��ˇ�L�7mI7�~f��j!g:����<�8|���Δ5����#BV��At���!Ƭ�3A�_q|2�y�ésl5~.P�ngd�S2����yV��l ����"AR�����KW��z ��h����0��M�
g�t�K�ص�u��U�;���g;ع�q���Y�^�e2��ʍ-5{�<}bq|�
�I@�oQ����+)D#�x<��Y��T@��pb!��m��j���"8E�s��[vkF�";���-{C���Na9<.���C�4.WyK�p���ZC�&}x���r0�Rx�������Ԫ��N��I��8#Y�T�U!
�t�����ʅ�u�T��'(!a��.��S�o��Θ�Y2)�Sp�l���޹�ud��ؚR'���5�7b1Rh�2�q\����c��)�V�u"���!��$\t�X�:~:>1ӌ��a��w�B�al'`\5�s��o:���_S]Pŗ6���K�����j-� &:b�G�����锱,`!MJ�L��l�挲�mc�_�b8#"1����܊��t[C{l�P\�[V���t�ZеA{O�@�f��GV��OH�MԋP��Z0�.�[|2���Vܽ�:7;��y�
�9�A!Xx���j�E�BN�g-��a�V��n�dA�ï-����*D��b���SX8�g�3Ir�ޒ��АC*:�B��ًn~|n'�d����|�	E����jJ�v�^A7�c���pl�v4�ʅҲ0�֨}a��P�Hs�1A���H ��˫��8�$����Rq?}U���Bn��N&U?��;�XcaL�E9�Oe���U{F���riu0�Ov�ugy�+���Q�o�g�u�~_'@��R��P���ۿ&:�Z���ҫM!|�4�!:l<�A׼���܆t|��2��*�J�>A�G�jjGE�yC}4a^�)>�'�5޻��8�k��N5�͈�����c)�5�q1[cn9w�z���} F�^s�
�L���N�쇹�����<�X��X�Lo��!�j�}��<%YĶ'�S��"��^�� mS���a�\c)��>����{�yt��N���u�@ؐ�Ų��
:�R0�\��U�L����1m�R:��g��/b�h�E/�?y�km�꼯
{�e��Um����Pyo�_ؾо�[�����{;�9I�D��-ZxR�b�+p݀!�j>#Ȍ�r\\�׃�#y���J@t�w���l�Ԋ��D���s����C��a�'$J�'��U��5e���F��*�+��U�:�#�8��l;]��mއ8bA��8�.�0oj�K�g
�0�2D�	ѵf�CU+�\H�ɤV|��s< ���Gt�.-��_����2��٘Z���h_|�X�#��	������{h#$g"��4�Bٞ��^ݷ�Ou�k'�K(OT���&�����4G��aW�<�*U*1i��H<f.��͉ӵ�<�W�mļ�0Y.�G����s
��w,��b:a��5���5�]�br�Z�io.���R_Z��&�>�H:���̰�a������<n���j�j Jw�jU}��r�OLO`��ߊϪ�=���?;�Z.��6O5xW��C�0������l��	��N�Y�d�%BǪ�y�gڞ�bf�����<�/Na�F��Sv����6��ee��)�QF4!5��ʛ7�a�UB�D1y��.r�s�a_t�}�oc�CIq�++�B3����:^���M��d��0O}J�K�y9�e�e��y��.-����O
�q�F�����1�.��;�F��qCl�H�j�1VM�m�7����U;ڭ�HS~I�WAx��E!�i��{i�Z)Q�={|+�$��.<�����(4�V��qg����Z]NT���m�w��5�QɍN#zb5{�<���gj��=w]���D���yW����Ƈ�n)���1�͎���8:wp�^ۃ}l�<w'JsA?dҸx�b��U�_����_���
�d!��jv��ѭ�p٩�V���y%�C���;w>ӝ�7Ǵ8n�D1�������@�"^�u����)���u���s�Ш���(�>�8م��B���\�>y[0�UH{5l�+ד2��a^#��-�a�R�^�\~����cp�7(ENؼ���)g�_'[�h����6�l�"�o:%���lC�aC�_Od�zL�6W�lOW��kԡ��g��H.���1���[Y����&u�
�b�&6b�����Ok���#��ˤZ��r9�I��!�
qx �Ǘp��ϱ9QX�����(����X�_�)�f$^I��U���ِE��t�o��bbb�V��f_�a��b�w�=t�m��t�֖�3W��(F�b�K� s��(�Yn���G<��S�xy�L!V7����}��`3);=��xc�� [�M��)�ܕ�q4��i���.T���XT���իH�'ؤ�p�I}Ë�w~�����[��P>PIh����;�3#�+8�yD�	�»����[�m�%�51.����*���t�D�h�����t>o�o�J�R���9�KX���AWe��,�����!n�f����\��4 >��veD�+�1Q|��{���ߩ���%gvuO5|��A��\����0���T��<(� �P�_R"l��9��8�o�Jǳ���h�b+�R���@Lw[�c�����)�Ϟ�	mQ�GNb�Ii�x�\�&��D1f�����0N�,CҀ������5Q��F�:����x�a�͍���rñ7�鿗!g"_0�����n�͎ c�چ"cqPe��l�uMg�,�'�=q����{8�t�V�8�pN��퉙}e�߳E}V�Z�}�tf��i*�41�f�b�0��}�k���Ep�RB�l {"*�	��p�Zs��y��åz@��u��*)�vm���^��2�|�cEq�1�Lw�{@>2������O/j�E���O:>�� �9 �@W�(~��Ok��*�^��U��hF����j��Tm�{طW�����1y0��̪�B:���Ժ�ZÜX�:�e�aG���o�e �%���v:Z���7.�m�]��������{���o:2�Z`������1;Y��Ҋ�6�u�Ɲ�3C$���[~�&z{d�>Go=��.�q�9��ӗ�ӫ]tHzY�9��B7M��(k�V7LlZO;rt��G9��5�� w�N���-ė"�]��e���	-�ͭ,�rJݩ�,qgo���B��30h�x�V��q��k�1v�_>{�:���!}��DP��VA��}�os���$��dWM{B�ho��}j��~�2J�$)�]��T/���ۇ�x���^!��U�r[
�hw j����e�A^,զQ[qh���yo�l�\7�4Uu\ RN�tn>���-�{�^��PZ��|�}��9>g�A���4�g9&͇(%��F��(���c��^�M+I�ѻb�8�9��Wt�<'E��)���mp��۶�jOi���+}tZ��cka�/n�3�t���j��&�r��ɹ�)���ڸ���X��26�&��B���x�I�N�ûv'�䭁F��me�] �7J������6�)��1s]dwz`��_l�f��E�Gh=�nQg4AAP��'�y��qPK��R�,lm�k���ݹ�ݒ����J�Q12�V�իN�&J�.��7*3��Ѽ;c��l{F�.�m4ղ{ ��	��g!�J�B����b�hХf�Pb�!���I:W�G�I,��8��R�Fs�9��H��Q)�B�<���iضp���:��A1v��307�[i5���y�anC�=�-�5{uh�r�Vg�CQ�u��m4�z��W��Ic�V�_f�R�7;q+� ޥ��q�a�l��uاlݤ�.pr`�{�$����y����g9�*dZ�n_J(X�(t��fXu���@̟:Ttވ�\�:�L�ML��U�njWó��'�"�p<���5�t����	c�)�B�E;���O#���vt�����f\̽�Ñ�qe9�g��������(kzV^>F�zJV�dV�5�Q�7b�mp�7���ϔ����oQ}�9��y#fg'��ky9���n`�vx�1��x��u`C�c�*��w�*n;z/g�]���;���Rv��v��o$�#�.����y o23t�WoS3wq��8^�R"U��ˤ���3@�Lzl�P^�{fT:��D��g�����qRE�,L�� ��W�2��U�T��ӻ19S,na��O�t���#�!�6Y*�#5�ԭ�Wf�o�"�6�����;�� ����^[[3)|��v�%)�o��[طH��4AU����&�s���n8-�iۡˌ�W���kVR����+)�M<"��C�c?f��H��V�6�Y������-���|�Ι�7���uᜒz����fO.����H@��k5̌���d���46��(^]���E���N�� N�݅����]��j���S��D��ǉf��6u���/N�)�r��dѧ�U�Gu=���@H�aX1���2�PVДdXE"�J�ԩr�3��AjJ��Kl��Jֳr�C�E%T
ȰE��"!U��#JK�,	P1�,�,�VAAdRKm���(�$� X
�B��$P�leF�TJ�)X"���Lf2,Qj��&e�c1"�dZ�X�6�����V�*�bLT
�
0PX �P�Y	��(��"���%W�R)(��11��Z��Z��%eb��T�Ь+YR,
��*��b�l�e�b�cU��1&+�L@r�&%jF�eh��TR �J���e�k*T*���Ŋ�S;�]��w�D�`�Sv5Gd�}�r�J���jm����.p{�e.Һ��4���>��|�Ԅ��r�%�|�)SY�&�o�w�z��R<a���{֤Y�������>}f$��X|@Z���w�:@�Vmz�=g�>@�o�LT=aS�o}�t�~���zVx��|�>��<#�C}""z������幆'��o_}�{�v���b���Ȥ���^�:�3L��s�jt� ������c%TZ*�_z�M=N�x�OL
Ό�����bN̡����p�28Џ� #�����l���EZ1�5�o^rv�Că�w� �׉1�fs;N�x�L}I�^�;d��ΰ$�+���1�V!Y���:B�����,� �f�0��Xa�����H��٘���s��!I��m=����6�NӴǼ�1�$��rs'� ��OI8�`{�f�@�bt�9̓�钲��w��:H,�s̚VbJ��S�b�I_��L���ϨDCD�e�'3�o�C~����z!��d�����I����1�9-��J��Y�N�1 ��}�\�m��]��q�����N����y�H+�}�t�3Hb|�A'�vЕO���6��ivDE��>N��� ���l�Ε���&��+�i��@P�K��jwa�>B�d��^軸��>Iw�ڝ0��l9�I���Rk�惥`#G�B<gqG����:�Z9#<bg�{}�^��1����[�%B��|���1���b&�T4�U'�����mH/��t4��yd�:�ɤ�!S!ѫ�Ì.��<@�8�M�{��:偈W�y�5Nݾq~�~}���:C�p�:gL� �ε%f������*���l6s�������k�:H,�'n;�Èi �4uCi��B���~a�11����|Do��Ʒ�|ӣ�-&�
��58ͫ=IRW�s'I8�t�2a��bҧg��]IZ�+�T��8���ĕ
���c����%{M��u�6�Y�;C9d�1�-�tzu�{c��8�_{@@�:}f<7`c��;�q�*VO.���m�C�N�9�$C�:�sz�At�3y
��%d�s��:CW��;�4CHv��jc%I�TG�Q���x�ٌ������X�[��cQ4��/axv@�M�V���:�P`tw-$G�����'�/z��}s����8���J��t���� �ӊ�L�Q�'}�/�����n��D�(�גp�i7w�,�S�ywE&B	/!�WDo��*����-�$�:�Y�7.��K-�����D��f*�Dpn���8ɤ��Y�wdĂ����l>a\@�y�!�LORz��~�P1���1��&�'���Hbx�0:=�j�0�,��&#w֩�>x�"�����*t�T�}h��#�,C�@��x�z�ά1&��6ԇ�x�P��OM��̟$�}�C�>d�a���1�!��51���V��É��ޝ����y�1����rE4��*{�E�'���4�:���d��Z���LH)ѻ3H|�����I��8ó�p��<I�%߸c'��+:�t�����$GۻNKxp-�����)*θ����<�z7�!P�J����� �׾PSL�eI�u���$��1R����=CH*��z�!�Y<f$������ 1I8>��:�0���N%��}c�@�JÇ�䩤>I_S��9��
$�s}�'��{��'Y��>N˘+�� tsXi�2T��^��$�T�=La�
����=ađ�x}òw�S�o��]�����H9�0$5߼���C��d��� ��䙾���NЩ�;޾d�AgI�s!�T
������c
������&!�&>&��i�d�9��^?#w}�T��/�3z������}�$�!|�q��gyH|Î!��=M$|��kI�+����T��SӜ�4�N���|�P�%d�����=$ă���+4��+7����zﯓ��vb����k��#�"�E���$�u�E��gl�ٖ'��q�"��+����o�
�$�]?2u�i ����>�c1�Rb���*�} H��N�?3(mw{�mQݽ�{�}��m4� T��zϐ�񜚰�Aa�h��}I�bA�Y�0�Y����|�C�+�x��$6��5��B��
�O~Ì�n���g�:ea��I9��zi��Z�y������}w�g��+'7֔��]y��&&�z¸��u����1��ޯi�Ag�x�����%H)��Ì��������4�G���;B��5�I�Fm������N�uuo�=��͔�-�k�[�=彣0�v��aQÞ2��}HsU�͜ڐB��Cl�iY��fQ�u�'v�b�y;n0�;�I�gM����u��A�̌� 駱�)�FUn��H53���͒����t�I(?~����T4���&<�o i����ϰ��OY�ã���N!}�x��];`T8��}��<N�>w;���'��2�'iRb�W�w�	�﯇����5��� �0�O��ݰ�Ԭ9>���x�& n��d�*�ė��h�!�NЯ뼆&��%I�(�"��Y��4�S�M���!F�0�xE�D�kq�O����hz��^w�}����1��n3�K���הV!�����6�^$��c�;N!�/��P8��3�17�bAT;>���Hm@�̰�1P�K�<��z�����]��:�Ѯ����{�x��z�LH(|�!������7t�Y/W�;��&�ǎ��%g̕+{�j�U�n<a��i��+��(C�>La��{��6�Y��;��1%H>������懾��|���w��>IYP�>Cެ����{y��Rm6��{dĂ�n��4�+:�ϐ�
½�a����J����ed�_w�5�'l�?�D}� ���0(G�����=�w��޾�?0*0��{����bAM���Lq'�V���%I�ެ�A���΁���@�+:�4�L��La��1���ϐ�SI4�I��g�{q�����}#�_�;�c��ELR�Y�n{�B��a�+>g>�� ���}�t�&ЯG��RT��P����'N2u�4ɲk2,�%�ɉ\H*�D�;x�$�<�C��������G�!��D��{�D�6�e��:�O$�� bAT�Ì*q��9�}C�1Y�C�ä%Cԕ��oG��H(l���:V����L�K��s>ΐ�%ea���gL�+>� G� ����L�9��3��|<��OX|�&�vÆL
��|��ug�t�Y�zZ|�!�J���w��N2��x�vsD4�
��u��6��T���I����Ѿa�VJ����C��~�˽����_75�^yǦ�b�-�������~-F? ��'F�,>a��n��=B�C��q��P��{�v���1 �s�J�礞�Sgy�*ɴ�5�3�:H/̏7����@�.�^���s<��:���4r� �=�����b8��F�L�]��t�f�j��#Y˃�A����\>Mv^"�V�kh�E^����P��[��v ��4aO$��(�Y�������x&A�C�6��駷�!׫n.���#�sZF%����z��}��������Lg2Ɍ�eVv�MP�M!Rx����d�hm&5���Y8�t�&/oΧ�Ӝ����|ώ:m��u�L�R�D��e(*���k���F��F*	�쀸��(;��
�~"����oQs̴r����7'bl/H]�?.J���*�����U泊:�Q#�2|hB.u�Yk{eN.iő�-J�p����;�2��(�Cz���U�!�N��Ȯ}�x���������Ұ�b����aT$�ٿ�TG%�Hںrz��b4_w��I�Z$ȗY������wN��Kfk�>�V/��T�f5Z�z���i!�3���^oQo2^�V�rGU����c0�\�b5�nP�o!���GC�S�m�X��5�x�.��ֻ��}�驠��A
�m[�5|t֫�^!ZfC��%���K�b$��ټ�5�j/L���}���2`�����,���R�k�y�3��u�� Ge�s����C��Y`8j��D�q�\l����tۦ��+�퉊�u�Z��TE/L�b�E,�Fܭ��.�c�X������5v����]��'oAWMJ�78�u^M�
#����ծʊtU��ε�G�ݵ�|��mJܠA�{���0�De��%���*z���J�Y@!4e�{>�ow\�eV�<C�i��N�6��sIAk}�>y�f>�X5��|r��v��f�s�������]t���V���Xt�z�(FP����kOTc�3��0���
��Yxm�L�:�c�#\c��|���R	�P��[+_3�'o,��(��Hq.,^L�w��Ue3���q�e�T��A\��˥,�j���36��p��3�P���k��|y�c�J���Wl�v�9̼z>.�ώH󯞷_�U�_����O�"r��P=����%İj}�Bw��4�S�WH]�����8R���(!x��Vw���`���̩}Vl)��Z�4p����g��Z�v����<6���a�P]��݁�*-�*
�ԆP����LX����*Z�ץ��ҟ��;� ���j�����.m'"}l�]�:�n��P�=Wz/H�R�u�l鴸.���<?Tbu�rC*���qʝ�ų�f�%M�w�w@%Q	�z�vǛ���=!��.�IRߔu�V��8�1T8X�x|-�OD9�mPfd��ܣ*&N:u���[�z�z��3 A�:n�;.p*a��5m��S�8|v�?ʋ^�a���;1>ՠK�'���O5�;��6�B��{��`��RO��`޾6�$CSS9]��s�o{���X���8q�Et݌NY��{���39�[�|�zJ]!�n}�`��{S�y>��7>*�$+�L=5�t������0�Y�����u�i��i��wHqʑ=9��AV+砞��聇��?���P6���:ϑ:��2�k{����2 ���!��`[��a�]�������N��f+\ǵz�k(��e����'��
�Ʊ�39���x˯�rw�4F�MQӣ"\N$��8�J5Μ��{!1�O�?P��-k�kِ���M�gp�O:��}�x�Z*��<v�����Z��k����߅�;�Q�FUlY�^�6J���M���fӜ�W���2aR�6Sw��{Z:�;:/�0�|�e�B�YC	�6.e{*��X�"��(s]�ރ+�d܂UU�+�eL�0�i�OZ�R�X��*K&��WE4;���<�oi�f�k��I��[�k�Pf��ߝ!���yp�A�<]�3��%��n��	b"Z���S�gQ�E��mOj7�?jN�8�H�F��৖��,tGAh��㖪m%=S�t������S�Y�9iP�����u�iR�X�����l[=�%���$�9��P�ݡ�"�N�a}�kc(��nm�M����]�
bUr r%%��)�.[��R<nP<�M����^���,�X�bL����)���>���<�)s�W����Hf�1�<T=���1����%��@�|[Sq�ټ+��]�(9}w[�H��(1X��s�Abş|��n}w��BOa��Bfa.�"]+s�G�ۘ��,�ɾ�6��n���YZ�$!z-`P��גqأ{+Ž\/ C�����)s�.�o��$gZUs�n\���Oѐ���L���9P��+I��X!�^ǝf���P/\T߳��=�JdV���B��@>ϊ��
 cN�1`]W�=
���{Bv��/"ʲ~[A��E�sX���8��5����ʥ�ga��<�,�e80����I�8�6O:��0)��ћ��H��U����Έ��u��2i�񍹟���=��V����9�31�}pO�X�\�\+΢�����*��
�IT�g���Ң5qT�~7�x�:Tj.�g��J!���5�u�#{(C��z�K����d���]v����fY��^/���ˑ�Wt#�A�O�A��t5��W�/�
�X��a=�����+��^ŀ�!����t�ZH�2A�{Ǐ!��/y��r����{���t�{j�DI{�p�gvZYz�y��ֻ��b�{s0�շ����,�<�bŦ+A\)��]B;_%����+rԂ���s����j'cߋ�9�¥<5�[�=�/�2_����oeKaWj��ў�������_C�7ǜ�R�y8*��BhH�[^[�R�{-��(��֩�z\'U�F�nS1���4J�6`wU���u~d>���ڮ���[�ʦTIkOb�N�bL�ѫj�T��@�v�nX����Q�uqv�d�49���~���fk.��\�N�FT� +��gC�N�1�8�zn#�&Uۓ�9WR��5%�+O��a6���G*]$���ǰ�S]�J_^�ʡL><.!=�*[ȓ��[{��b�j2�d�6b��$LMz,Aq�ܴ,$ϱ`Jr�B�d�Y#����G�s��Y:k8Ce�� ��d_E���N�� =4e�eoMl*�i�d^��Sk�0����gi��8Ru[9�yLA�� �޸N� ?�6�����dzy�(��'VV�4�WIl�/�|LXރ'�C�@6rN "{d	����E�1&e�u�U'�T],���z���E��5�K�d֔*�F���6�g}�o�z�$��!���+3��r���E�{��,s�� �ȣ���{1�5��U���N865�-ἁaF��;��-�۹�-�M��K�問9Ն��B���ȏ0��)Ec��b�$8cVކd����m����e�C~�=ʰodB$!>֥�J,<AS*���rX(kD`�*����f,챶p`Vp1�t��@wS�a��ϩ�Kňt7F3I�X����woy��Ŭ�o0׫�ف
�n������V,��.��$�����cݮ�9/2��5���mQ����69��O���?�KU�y�3���v2za@֬��3��m�ש����>��	�!ֈm]p���~�ۺ��3�L����o�I�!��[!��\G�"U�(/S�K�sn����r����G��-�F-L��yMk������P�Zٖ�{n:�ɝ?XC���4�,�7�K+�3ø��6�-�xou�d�@v˗j��g�)�$��N�,�(Y:t�ч���d3�m�|b�Gؑ'�W�3���ߥ���	tv� �*�
0�]<ʬ�i�s�+��pk�h�~D�f�w�ͅVm�D�N�<}L����.˪���*D����ʅ����yJ�(Q�]{r��D�.���CbPB��!ʙ�t��`�(�|"9d�{!^x�M3���&��nW��A�N9���y�q>�w�U��Q0�U��k�����F��B�:=p�;K��9u����.jN*��o���dS�C[��W��m����/0 �7�>5�weLwN$��<��VAvPdf+� 5� �]D���@f�J�{�-�v�ݨ��0٢�h<��:-�_@N��
C(Q���+f�%V�FSǱh^!v����]��%c�
�Xi&��/���.m'%��	�Ȩ�uP@��6���:�3���q�3�q��g$t�ھ���4�5X��.N�c��~|J=�l�1��U�MJyF��sy }����I��e����Վu�"�p���_ٮ¸�*o�K�E,?@%���Pa�|q}2W!���2���me�����Bj�ÔʫP��)��/"�C�����1H�Ҫ<E��Ry��+�}Q��7n��۝�Xo�{_o�b���4k{%|���<�����F�ä �JP�UP��Ԅ��&E7 `h�4���(X]�x��\�>��qm��3���j4�Y���f�ð��µ��w1�~k(�Ӗr���:�)d��f��G� ~���ig�L�0V�W�o�X+'��Uf��P��o���T4�/[\�.#L`�����{>o�ݪc����i{O^�1�g?x�/������ќ���o/x'���$��T�1v��(n<yGV���4r�'���b�v[��y��uI��c��b�R͈��b�F��8qtY<o��e@%��ad�n�lujl�fM�����md��[>��N��7q�e�.�{R���gl7�<Ԧ��^0[�	_�]��7G��4MUqk�	7k�{�z^b��`�έ�Kc�+Sl�&A� �3f�Ѓi�sG�@��n��V�Z���:C۔�̎�i�����y�G.���4�E��q�U��S�k$P�45G����mZ��Hc�A:�d���J�s1���))ס='�N�a��Am[�-Pk�bi�o:��|�\S~�\:�)�څY7Au�W$y�ܘ��C�t91x��n�d�Wcf�c����!��������ި��y�|�!k�B�ͦ"Vm�U�*IHaYq5�ldW����uQ�ӑ��n!��(ɍ�.㒓ΤZ]]s-�{� <0d��I�8I}�7���eF�r�!�hofH�v3(Qá۾9��� �:ݺ.w��A�j�R�����s��[��Җs	����kmz.����o�n�t�B��-AQ���۫R��#cjM�R�q�)pM,NP[O�--h��w��Ź��%�M�7�8�@����f�T���{8��k�&cд�Y�f����է*�=���)r۬�থ��-���Hm
�u�m��J��n:;�C5�ة���4���aT������P�FV��2;�2�������v��c�.�£-��#;&20>�Va|�#B�a�&bʚ�׬�y�
ZrrC���NM�*c�˃#T���b��V���v1�J�*�'$;E�nwX�U��F �gt���{�2��b��e�iT]���� ���g$<��v#�T]�B,벏
�a����l[�e[Ӵ^�Ԍ������Ws�5�-z�G�חY���ݜ��w��;�GS� �3lq<o�f[4^�-dm�������q���tZ�u�����JC�)�)]�K����vp2�q-n�kd?�b��T[�j����ϵg)�'��l�=����{����e�pDX�Fl=t���ٰҭ� �*�ZP�,����+T"���d.�;`u��f�|�y��Ug|�	���r>7H�g{���\��`�F�*܄��R��Y�d9x$�z��5�gF'�j� �2��ٻ�k4�V��F�=Ln$+k�4��m�$�y�'.�C��s"3f'b}ն���N����=Yx�{$RI8f�um�L+���ޕ��"q_u�F�^P����ʱ�̔[T���g����.����'7,�B���Ow2����Dzѱ|QEFP��P�CI^��R5�u�����t£ �]�F3f)4RcItovTY�l32q�^�oK+7�����B��7]��8#�@$�kR�U"�,J���
b,�
ш��VT��@̲�(*�ˎ$1̥�EPUE���1�YX",�Pm�bV�W�%Ld��J�YS��Kek&e�,�R�-��lB��V
U��m(B�iB"�QB��ŕ*
E
����ʘ�
e��+RQ�RF��,B���VKmC�@F�QVC2�,�R�pH�3,�Z����Kl�E�9i�E�e�R"�`��Qd�s(DL`��2��2ذ�1A�Q�k�����J��+*������1e�b�(�(
EF(��*�kAe)[*T�3�jc'�{�[ص�oj-u=�˧�3��вv��\���5�c=Q��d�*j�Z�-��*V�����wWeF�得� ���}Iz�BT1�VO�	��ˈ�x�q�؈dR���O�ڡ%{jb���܍��Ξ��
7jа�s��$ ���`�`��Y;̾S�j��R�P+��<yb`�R�=��;1�Ӭ[���T+�8\-�nk�8_�鐊�`%���w��#�����=It�H+���1�kr~)N�:ܑ	����
zX��A
�I��L�̍�n�4g��nru>��)��S1�!f�%���gK�َ��#
�ǖ@CjR�^/�cj;���d�B ���}��)�0_�Oa��L �\�p��YS��5��+ x�Nd5�L�lW�~����V"���ҥ����J�c��^�ρC+��!���}SݙL�].\�*w���A��D��9:�2��|	�|w�r�m�V��Ӝ�Q�rp6�q�v�Ń�ؤl�
��w[�K@8IRxڈ`KǙV}��v%���wa�
(7��*�����I�=HW]	Ʉ���1���60KuL<�,�e��L�,0�����k}�V��`݂i�V����VG+v`n�U��y�Qz��g��ߐ���Y��X_,��h�oT��Fv ��QS�ޫ����f�d��{�%����[���Q�����B�q�N�keXSu���m�ݥ�s�R����?�_v�G��W��}�[��F�ݬ�Nɒ���.��R�d����U�Bon���æCy$�T�i��>�&81�ʜ�3��؛=�F����&-]�ToK�<�T���}����4d���r?����R�-��m`�DU�����|���cC�7" (j��n���5p�j���[�y\{@�y���C�U�C�T'+=k��%~2�����\���=4��홝���5�뷧#[��N�m�=��>�<-\��0��_�[���z܋�#x3���	��to��~�R��r��u,h�W�8'��9l�()@r�m���p��֗_�޾`z>��������t'��#ǚ�=����<w�e�ـY�ӛ����[�:����r�FTJ�E��^:�DsO1�˶@�c�v	�v�;z�ۘ���m��������	eH�u5${*�˰�0��J{?$a�Ѡ"�ghșoE�s���T휗	�fY��nY0� �E��<r�%�Zԧ!�
�� .J��Q9�c����nnk\�ׂ�lύ5����զ���g2^��R�˫\�9���o�b�ʻ2����4ۧ�Y�H����X&�����Wܪ:���K(�-mSz���%m ��WK��U"E]�M��G+n5u� � ���0��������Gβ�&���ՔpzqR5s���@Umd`��CR�ɐ��c>�Ղ�Un�v�`Աf�*͖�F�1�kb����s���OOe�>ɾ�'ʌ<�*���ۘ�J�P������}&<�r~�hk�G_K�I�L墦�"��J�$����7���/\O�Τ�{�Qb8��E�U�Rɋ�ewB�zjx����tץV�3X�>vv���+q�=�/&b��]�����b���2�j��o!���E��
F���gY�����p9��pԯp

�Z%ҷ\>���Kke�=��B���ϴ;��,� 4�[:t*�yM�`�Ӿh��K�8lV���h�m�Ǚ3�ds�.:�U}��� Cx�
�,c.��dp�|l�l��M�i�z�k�kGZ����Ƈjsω}�i��PRci���eF�x�ȍ?1�p���2����M`��>�
�)�'�Xt{��w��/�øɝ?U�|��M/�O&t_�3|����okҹ�گ��K���D�����*�DC�ܼ���C0%��2S��AXZ�ڌ�e:����]u��(!4���JnUc(�nr{�gnq5��Ϊ��R-��fa�wAu
�w��	�����9�Z����ֽqK��E�Y�M����ۣ��n������菾�>���T\+:@�?�VRn"f���E�'C����)��gt�ta�M�n\������/�eV
��~�Uj���5\ T�sSY��M9���Ǫy*���˻1�[ �w�	Zw bt��W�`��9��ET�)R&�0��<�H�Ns�Є�w%˔��}�pr�"�W�X��~2�AiP����z�p�+7��{^�뮊�w'��4���ݨW�͗���Cv��wDPRT�P�PN��y�ぺ���٥�O_E`N���f��_ӐJ�I5�C�Fd�} t'u!V�sp�;7��S=/��� ?�`Gnn��D��!�~��/N��T�aRT��g��ώ�gG8�L��X����@�6�
�wJJ$Ɏ�u2b¢�I��Tic7��B�<�M���[%G7��%�U��z������"S`R�CG:n��9f�xz5N������Wd�м��j�V=N(0J�:,�s���U���'�oΨ�ӳ�K�~
T����f��]��Eݰ�2D::�F�-p��[������r��e]�piou�����[2:�-���v��o�V�2��X6���GdX3��	 ;,�S�4��D15�I^��_u&�!��n{{��Uv'd�{�}������X���Q#�|�Gdl��Qb��U}LN���ݔ%w����C����5���y����q�Y���fԷL��M��� �l�:q���k���s�4BvS鎮����k�ni�t�v/}LV�r��XʽSR~��QhX}�6���5���Qk0q�D��h�ލ��4]��kh�l��9�`��1�1A'ܙ|VDve�}����];[�ŗ�X3/��ӊ�y��<���������0�#�Q���ǅ�\<3�挽�z���ْ�V6g�[�O�d2��ʺ�!��2���W+>�@G���P�,�|�z��s���O�y��u��U��b&8r�,v�C�˺�8ܔW|��̠��ٛq�h^旷Z�Cp�/�מ�+���������g�<-�ۏ��-tG1�S.��iq̏���qDf�C�ߩ��W�Ԫ�|d��.�huҾ8=��ʰW	~B�;��z��g��5����U��e	�+�B�����S`�*{B~K��.U9�C���*����}`�U-K�����ܛ],	!-3��ꅮ�n�a���R��BW�DI>�F�-޼�Ú�>�nv�O��H��H���e e4;�lu,;}��͇�wG�<P��`n�X�jse�n�r���>t0���QJ��m� ���*�k��}��n\��?T!��}�UZ�IE�9?"�{�m*_Z��M'�����̰�Y���`^+�%X9o%sW�+bD`kUro�ܚ�k�O�|�x��7�;|��d����V�~k/�u���I��<�]q����"BMP� �����4�K��xO@\'s�d���֣����&F��hO+o��\�~C�D�/�2ð�����L1�8X��N<6�d)��|�ڰ�ra����'kf�4�����P�|k���W�ېks�I$�[��͜����I[(�rI�տ��+�V�U|�yJ��*�$Ef�=r����fq�w�v%s�,��-զa���O|��2��{)W	
����*a�|���G�чu�JW�x}�s}�8�����H�1K�����n{�(�Z�kz���T&+=jK|�"�[��Tv*sy73�$�����1���:�1k-�]��'a���*zLh�����8`��z�z�D�Ce�V�L�z{#\7�E̱���ʫ�(<-��j�t�����Gh����nW�X�߫օ��G���~�oS�]*!���)}���7�����������.Q҃@�D�0ܝ�e��pRs֨�"G�q���WX�����V��ǭk���A��f�tW˥��Ex.-��,s�[W�/6hM�wGl��9c�̹�˻�D��5�n����}�����_kW�y���Ƞ=�4W9Y$&j5mB�҂Ҹ��D2�O�*� .��#3�_\ۄ�p��&=����xo�0��7�`J�}s���:�sv��h*�6OK+��������Մw��ܥ����<��i!��-��7G�xI���E��emח5/#�7ֽ�;����s�eΞ�pe�n�Ɏ��_2��;*߈4AJ<�9�:�بa��[]�r��ٲ�����>tt�n�����Hjw&@zo��͊�4����d�yO%���Ȳc�f��#�,4����X�Ǒ����
�!���QXA�x�o[�3�2m#=�ܚ�4�/�|LX��z@�I;6m�@4r{l�Ed�����޳�+4Ox�u:��X c�寻"�g�����V�>A�=�.�֏�Y�շ��9�˒�in�h�;(�H� ,7%�9,h������O���S�� �g��-coo)�>K���Z
��=���{�Z�=�Ĉ�&����R���zK�j(�{3�6n�9VG=����e立k��&v܅OF^�ߝ�Ǥ�;8Z�OW&�l����Q;%gv<�Z+%���ڲњ	V�A��w#�Mr:k$K/.�2�㮀,���"8���}չ1������)	��D[����OCo�2M�
妊f\�}�}�}�ݾ�s������s�`x�6{g�?zñ=�鿼ѳ���:GUl�lbӪ>�ߝ?l|�!��~�7���gk�_5u���G,5�r%֍=*���*\���2�'\��&Bp�/���b8f b�jvɼsn�;�x�(`��G�(p�G�b�9�/پ�;$0{�`��7`)�+����E�|��MpK/�r�\v��	uTb�(b�ζ�9ֶj����z���v�Q��SY�C�<7�KG�*�T����2 \�9$�S���׾�]�z�/���<k֢�'�� ��a '���Ug�HF�[���Qz�ĥ�:��HZB��]������\1���H�T�$X�J��^�"�V���X��R�9�ҵ��s�N��&%.1�*�2�ja(��sn����rx7;TS�x��/�y̍����5
�����t��"~�tD"zH��ع�(Z�l�_y�g�����l|���qf��ɵ����}��i'��ψ�ܽK�u� �z��*wk�N��a�8fm �5N���"�P�E��]��B�m<)�\�7D�;Ԋe���t)�\���î��g���V�x��la ���Y����f��F��+z�T)���Y^����>���Q�ܚ�dF*�Ø�˛�"���?V)zwC*P0��J�\�eǻ\�+�i��\;���m�O�F��	oh	��t�[�]-]	��4�^.�0��vm3���csJ�*��}���p6GL&�3��ЍԂ+�h	�7�Z=�u�THWY^a}��W�ݠ׹&���X�ȱ����L�#��'z!�Pb����b<d�6t�X묆{xI����f��2--S=�S;7�� L�,_*�`[�Bt�y�"�9#4$�8��W�D3:�k�����J�$�@�\��̝�}.�o�1΅;�,c<r}���*b����=T�y�-T��
���ߢӊՌ�xGQ;=*��*��6>�ֹu�y��ee�s
'<ͻ��:d^�&�� ��r�!�H�W���K�CHpߢW�Z^���jC	�u��l�Ƹ�:�[%Fɴ~m��u�4k�=��Q|���tR�]�4.��9��BcP���Q�[�pf�N�1q�,`��O�g�县�]�Ts�0�9�U)�ty�}������ϼ߸D�������PN�`�3GQ}<�F+��ߝ���|(ԕq�ʗzhKd6�p�Kb�cSC)u���*6��o�u12XŪ�֞2_3y3�v���#?��ia�6r6�3�������j�GT0���W��YQf�0uܝ����a+JY��}_UW�To����>ݐ?%<��گ�W���X�Q��h��s��dp�Ǖ%���F�f�e+���­�s��+�`�e���;+���$�Ƚ��|+M�nL�3�Sy��������[�u	�P�7�iu{MJ�|d��.��UҖ?q��8B�����O79�]���d�ݷD;�v䱰`������S`#�!F����6_������AY��&M�Ԟ�ه�G�3��A�2����:h�-�O�R|�3=m.�w8Y�+]�yw�ȭ�n������I^2t�d�>����7�`��r{�m���'�7}PL�x�B�Ir'�U�\3��c>ޱH\qb(Rj�}�T5�����K�/	�Q�ժb��N��"�o���m9:#�&5��hdr�,�D�P�XvQ�V���[\9R����?�E
ZZ�L1��a�\�l��P��~�p���Z�ө�˃�NR2k�KU������i�&,1�4[�o��^΢����3�V�Q�j�չPp�(+�{���JM�˓��⸻m� /V,�"����������W%���LsE�r!}��Q�L���R�Mg��^��U���y�˫�&�I��}&p3���͙!�}d�S��X��ܚ��A���.Co�en����Z���e3@z��o&�Ҧ6P��Hf7<�9)Zݫ���/Q�7J�]�ϗcp+Hp��`ј��&�(PybJ���Ve+�P�Gm�GjĊ︓��X�Jn־BW����	�{J7)�k@s��L�cm�Wgr����r�T���]x�g
�����k���2���m���3���:�p�ue�@�{{�a���3H�xw����a!�Je0[���n��lid�݄�>P)��t�k�x��:�9 �3zﳻ�2�]F�.�waWp�5��n�q�ʮaސ�<���J�͈�Y�{�ܬ�|�U�oD]�T���]�y���QAN�ь�WӮJ�hf�!���{�%fNJ�*��`)���Y$s#�9w��	ė��];z�w+0۝3 ���5�J��o��A�G}�L�".vk81�R�cލ���u��Pj��C��Ԏa����+ݬ��O��I6�m.�,.��`��N;pd�F�җY��)ڕ��J���j��\��}�A����.��tlӸlKz�P2g<��U�r��v���q�_m��&��KB��z$��m*��M7G���7�\���m�3�S㕷���A�3R�b���EN1 ��`��@�"�(4��#rZl��t��%�Ź��P��][;�ͶYW,D���Y^-:6�޳�Ƀh�:�["Yr���cC�\����gPY}n�i�����D���0Ȗ4��*0���]��ht�i^$\�:�6�wWiB3i\����a�"8 y�����g���W�e]��"���p���:-Kam1X/�nɦ;{^�ТWf�D�T$�׮�0ec7W��X��*�NܖtUe���}��9u��bIfrg*cZ�][W�9A��Y�@�j�H�ԍ]�ʉe��:�Fwp�Sr�q͌���N�G��WSI6����<���#��̎
��Ӣ� ]��JΊ�\� ��i�wjRA�Ks���Ʒ�Ě�Q�8����4�����n�Օ��g�$�)ExN��o�-���;���˕�6�9�%nч�K�M!��qH)o�P���g�.#��S�fq-T�}�R�O�.9ARr��\6_��[YJ�̥t�].��\��)�MXydj�`��4*'���%C�vm�*_qQ�ҡ����`.��8�5:f;�_k4����S��"���/�"3�B�*Z���Qn�'dma�L�Dd��A�"n��{��Ǿ$Kz����A�y�����ޭ�J����4A�%`�XAq��`�F[`��Q-�P�j(��J�Sb̥`�*����Uj*�i���֑f%AB�d�b�"-H(VDTR1E�J���6ƅ�e��1�U�Ƞ�J#W(fQ����aZ�
���E����k".%�Ŋ�ki`�X�Um�*�j��Z�і�*��E@������Q!QJ�Jȱc�(���1��1F*��E��[e-��J��J��iQ
��)RTZҫ-,YP�Զ�dX��6��EUU �dQ��"�)Q�5�QU"��Jʢ*$YRTTF*�EEU��_���re�-M���`rtw��ֆvR�0���
i�ƶ/.�k�/-F»T�h�;{:J�[V�U�0��a� W����>��t�m��R��'I�x�+>83SR鿝I�q0���sXP�s+��(�V��޶�����/_ڭ�*.������v5�E0k��R��WhW4u��m��!޻
�7���YU�r+�] GTl�c/S��[�ђ��8����}��vjH�I��GczohZ3�n����RW�CM�d���t���k��O�yJZ��C#���c�Asv��k:�#m����6�TD��V|bBgV�.���֖G�5�{��8X��"ӈ��}:�o]�q���$Q���x)e ����Q��s��ۼq�.��v��E��N�	�o�Qo~�l��`�P:���Bj�x�������<@<)ԓ�F<�u�{�^8يt�7,���凍�k�2�nQݻ�j��8�ޕP����hX�èWH�n+�9��	v1yvry�]�̰�~�a�'��;L�WI�LR�~s��P�/ ��*�/�ٲ�W@>2Y��#�Gi��:]�؂�!N&;zeէ�o���]�ē��*꽏t��϶аL9%I��������\�ڋ���|
��7��jkRE��h��4����u����sOAܼ�r�).��oܵ�Vj&��[�����}B�{Y��5&[���ش˙U����Rp�N���Cu��}�]�:f+��TLwk�P:�C?�>��OF,c���*��!�)v��ɜ׍��{���V��������7e���2��}���qKZ�wmm#�����q	��NSoF�ly�To������s����u(��u�nv-��]��\BPb)Ҋ�X���8=�^Ho��m{���zUP\{ &��[aG廞�/.���/R��Rƺ�^x��!��f������d�+O��sp���oz_r������Qgb�U^jltE��r!�jt�i�}u�n;N���U��k����թ�j.+Z����wr��o)��Ҿ;�7�����%9B���{�D��7�+�YX)��~�x�{)�⼕s3Do�RD��w����{b����/�r�	����U����Ӷ{$!NX�>zb�N�#�/^�4�#Wu��� �+x���kB`����w��T�f��)�=�b����E_vK�r�2Gt0��:T�.��&���Z�j@Xr�W���O`Zmt��6;��n��{&�fkU�K��Hބ��I߾�����='�:��8��N�$�ϛ?R�,�麸鄩��á�}'Vf����T�z9�]���痋�uj�ܘ�KdӤi�eF��a��agZ�Z�N��ڜJ��rw�w��n�u�}�9��a5��{��S�{ �Y��a�O*�����+]�}�a\�w>v_S��*,ɒ�1O��.3Jt�TY��d�/џ��U�~��5��*��
TK�T ��Sd蚰���Z�����	�^7�=��Y���)^E�*��c9�-��N�dn�5�n7q��_q�M8}pT۸F�h��/��<���vVX�EC5�4���Z�R��g�J�ީ)�;P�㰬U>��}����� ɉ�'oL���~+�7��A��o9O8Ջ�a�OYo��ik�܋�f�Ff�c��\�Cʃ�������˩{~}K�ʇ��׽$��ms�
�'��Sd�4�{φ�=k�����	\/u%N�N�z�T��u�b����i��H7VG��pW[=2�Sj��H{2�fE% �V�F�#������9�Ӆh����}�-Z����b��}}Gٷ��Z�tt��tW��y[g��*�\my����So�Gaq;o�h�F���5��{Ϫ����f��r�o�Xű_!��z��6N����=u���r{nҷ�>�~qS��i�ϣ.VH�V)��ǫʪ��?I�� 3]��g�>};�L(W^���{t5��{(R�x��w�An��x����b���mN��,;�>yэhr��	[#wf��t qvb��=���\-��6�i���t�Wv�/��guYQ�zU�i��n2����\�����%�X����v`3��7�Bۗ�S���y�����~]�dȧ�8�W�JQ��_r���v��.x����*��57�wZ�Ocۜ�I��&�uaj���u�����j��[�L�I�[m��[e�[�½l4�[C�*�;��>��FhKk|�܎�U�#�V���X�])��{�On���]�me�B4y. Vb�ag9����:)�%���S���#$�p�7{����\3�c\�/�Hٷzz81\��f}1�4u�����T�
�G�n�r]1��\M�#Ƀ��Aw�Zy���Z:��d`OofN��-��2�-��}��G�/Pn���!�K����F��ޠ�51I���]�k��'����Kq,�1ˇ���;�l�|7����\+	w��	��/�T���Y�zpC�b��֪⳩vZ	���e�彳���{y9Q���ꉎ���ӎ�u��%
v7)��2q�>�p�M�m���.'ϡX�Q���c��aL	u��W[�+a���pkw��`߼խ�r��{,�s�Q���:����Z�^�,����fN���[U垭�ǳp�����}c�<���:�W�����ʃo�==��m}㞅y����}�O6����;z1	C�k¢˵]�M�䶵3��E�ue��*�Jx�����=�{)�8�4FUc���Q��8Կ��5C>�¯�&��q�.Dyߣpoz�B���c�Ò������T2�mɹ)D�sSb�x����؞�떂�4{��ʷ��H���ȣ�����;ޅVY����o����91-�5�������aho�5J���U�ԥM%�и��vF�;�J%"��M����Ŏt\Ov��Ǻ˱�2�!c� ��5S�u0���QDd��P�Ÿ�ޅ�n�s��r�GeF� t,��ßV@\��Y��7���Św��n��K���d�Fl(�ֈՇ�3�I������ܥr�v�`\��ِ��n�����G7p�О<a5pq�>nHv'v�ˣ9�[̰�e�s��;��ɞ��:�;��s	eQ���:JR�2cHՌ�ʴ�a��cۀ�w�*I���P��v9ϲ'��uo+��5+}Lme?�FF��)v�|«�_yVn�ͯwVi�/g[���{=����Py��+~z�r�n����x��T
����&B���r�5]��>�➣���5�+��m��Ge|q]E�YP���5.S�k�ާ���;���ң7�8g�jwg_��n�9�A�����A��Q^�s��v�7WR���T�Zǳ��u5}4��ų�n;ȸ1S���22Lfͧ�8�n2��*���5��u�6}ch�X��i��$��-��srA���������3��5���չp�$��u�ֽ�{�d8lӸ��Ϧm�eJ�㰱��x�D��"Y!xP2��*;j�0�V�V�l�k�ʖ7���/Tɑ��ꪪ�����'�Z:��\K���UgF(�[����i��ogGu�J�Vp�l�K�5��rw�ޜ���d�*i�b��[,a|��[�u׹.,�1�z�M�Y���s}���`�SiPw�^�esȜ�Y��Q�\��s�c���d7�S1���x�0�6�1R�B}r���P�q�o.Sw.9)������tc��N��8���P�5���/�Ќ��w��N����y�t���~��&Rz2��-�9Z$=��V,�ˮ��\�����yS�?��.���1(S�ý�_��
]x���*�[�"�w�"c\5��<
�j ≯Ҳ��������?_e�tUuy��#P�	�P�e����g���x��vՁ���3$y����,i�eOq]L[�s|o�\p���j��f_m�me孷�rRh�xge�Y9^)�mmݖ���v�;)wk�h�.���
e"�h/��Q��p��܇��!~�`z�v;/�W��
]cW�GCZ�ͥ%b��f�S�&��D�G8|��E�"�;�}G٘���9�yz��v����$o��T۸Fȟ�`,��(��%`��|�Tu�{zj��ON�z�s	]��!�C�v���@V*����] �VMl�t��)Г:���:��sñ��]7ҧsC&�a(�Ȍ�e奒�^��S����쯎+��L�}�oR�:��||���'QWC�.��fc�[��<XߣV����hz���8���B�Ꝙ}s1��B��[L��M�K�M�d�6��C^���\�䯸��Wg���.�7{}q^�c7��ɋ�y��{���>܇o�MvKq��bU|������#����O�ߦtc�ۣw�e��j�����y�dC���Z=Ef�bU��=&<��u�+��1�r.�"��>��k
��}5���>��kh�N�7������mh#�4rh�[rl%�>��^.�ſ$Ҹ|;�u�L�����!Wj㵯֊��`�ba����Ë ��l 	{��k_4��f��1��s�����׵�Bɟ
,�瀺�Γ�`�V�f@��<�]��ƴ��i��@�k��'N�F��.>�y�s�r�_C�݈�7Q>r)�S���舏��ĔVSژ�nV6)�U9a}ws�}�VhV������cmmps��zq�p�:�)⡆�G,������.�ϯ���q�k�U���v%J��+i¦;�o!T[�I����+�b��U��uy�-��ݿ����MT�=P�༅_>����Q^���}�#��)o���`7rN=5��sUl�S����`9�v'��`<�ҫ����P��x\��H��T��.���;��N���p��=N'���ٞ��4���S���{��H�=;�v��}�q����Uͫ�b����u�Ք�w#�Wڝ���|u���x2��T=Qh\v��o�b�Խ5FoeZ�'�ٻ���É����C#�bw�cp\�Б|	P��r�.뮞!_��Q�y����w�)M�9k^��yy���^��W*�����$����ʦ�����b$�P\մ�8@��tJ�rsc�ʫ����5皽Z�A"gh;45֍W��WBzƙ`��)���)�k­��(��MZUϥ�x���9�g{R'T]Ȧ̵ow�>S���%ǅ��3o9�g �c�����Y�������!cR���켕���E�U��F�����^�׽P�ʇ�O+��WtT�R�'Ss����^[�<�g��],b|�#T��)嶟vD;|����K���?G[���#�b��8F�g��P�t���F�U�]�\�I;�5#&���5	�kxm}nۿ����øp�bN�J&6Ov��h@o��m�/�^��%ܯ�|;v�d�t��q�	T��u�'������|h�<�zA�YܡQ�9���e�TBo����n�����r�^�R�`N��ycn�N��|72J�/���n���n�;���y
��(�H3u�!����Y6s�.R}�Qg�,g5�̅Y�è�ҷ��5tr�e*\�̲Ud.Vr�kDLC��/�4�*{e__�|:,�9�wx4;��o�]�i��ҭ~�;�BL��������-�X�&� �N�=��i^)���6��F��E�0�SkxT��&�����ݢ�tXW���n���.��o���mGƱ��D�R�j;�{��mu�=bR:�#3k�夤�Y�C.WN����2ff����s��@3�/a�m��ۑ�}k{���oNT;�*]�u�Z�)Í�ں,�G��Aʁ�]��qZ=zB�U��Ŋ�鼨$�{&�&��v��d,���،5x2��}�� �GI�q�\Y+�I	YS����ն��^T/�i]�^��޵M�U?�x6�b�o��j8qUf�gc�ml.�&��6�2%��)<���6sR�T�6U��{6&5��eZ�}�!�](.u�5�
V�/2��ha|x�����[BW�dҳGF���<��-�WD�^����1����)R�|��LIc��t�{m�S�\R�ҙ}�X�s�7EqsO-���n,Hy4@���<�[7O�����D���Qr7S2�Qqc鼂�dsn�\��;��6��]�$��e�u�����t���ͼi��d���u�i����)�]j�]w]�*Bi��g
�O�����gI'��M!P�g�Ħ<cT���g���-�yI���*Ah��\H�(e-��W)�ӝ���J�KU��n
�V�J�!P��k"����^���[-}YC6(t�^�l��4k�r�������[��ZV;-Yɪ�;���ʙ<(ۓ��L��F�tCZ3)�ps�Uc�u��B�9�=�t"��V�e�S����"BwXP��43�U����b�����7O�s~��:l���BJD�3<]�il¹�̎9weMVsU�mX2qZB�C4�n��.y�P�˰�>f��0�xtd��$��ũ:�0	]IE��`�GK�*�F��z�|�)�����q�B>���G���^k(pޅ[w9n^�p�Cvʄ A�ۂ��1�a�P-QFS�`��D��ev;�'[
�1��Q*z�G�F�̜̼�,6"�
2��j�R�4H�K4^��C	��=�yn%Pr�^W-��̈��v�]r�)�{yzn��4�j^08���K�҃�ʆ�0Y��v\.�-�+I�.���t.���.Lօ��/a�V�r���@N�/��~��"��t�}B�of�$�:���jK���c�Wnp�d�=�#�Һ<2�*1���Pd����ɼ#u���v�{�#���#��뙇,�혛��Wy���IR��P&'T��vo�Jn�Ѽ�]�,�Jda&�b����[om��Ե�C3��p�D�˹b�ZOI�s��r��)�}4��;��]�۷LȲ�9���՝3�*{�tzSP���{p��ǹ���c�O04�-p�Ԇ�]]��bso�Y��f==l�wA%���[`t�ڶ4����U�dxkr�ax�.p*H���r���Г+Nt��$ap�T�6p�s�L�zu��\9�t���pM?�lٺ$Y�A ��?E�[jĊ0T{h���U�X*�b�"*��J�TE��+���KE����"����1Q�YiUTU���EEV%JZQTV�@�Jb��b�ԩm1(8Z�b�X*��ы[�,"
J�b� ��V���1*"�-�b�Rڊ*���lH�m�6������FT-�(��""�EVQ��ib"��"�TEQ��Ո���"TkDF*�Ec��*"+kJ���j1eJ�����+YTR�(�c��E�QQVĈ�*����(��**�
����EDq�%QQ�A�J�Qb��"�)l����^[��}�����N��8B��	;��5��v���W�h�8����n�gZ0�¯K��Mޞ����r]vq=��}UU_y�F�WX�7�v��X�O\3n���/��:��1W׏s�Q����OE�nTvsՠ����V�K�z��7�5`��#��m�}$�\�L,n5FO6p��m�̿����w��\�Q���>E��7��-�r�ޫ�PM<U��\�'�gN.��W����[M�f��a�5����3�NL�	x���K�kp��ك�%\��*���G*�K��Sb����w�VT*�S痢��y�=��'3�2j�,�ΰ+~�vY�ʘi;�髥����U���ki_j]��Fucx[ؔ�$MF��LS��T.�=�d,K�N�l�8�k������}0����Zj����]'�^�o�!����LS�Q�WvD$n<͈r����(X�:L/�Ʈ����s^8m���5L�b�;��+uR��&;����|���9x:��5��^WA���)t�|r�Ng-����u�(�0�
v���.�׵״j��[�-�U:h⥄9���l�=�:�Qs�@��^о	�ԫ���'̘KBn����@�Q_\��<�d.*���fi�gD*5��J�p|�Rem�>�舛mq�ri;铞9ЎYS�	�B���ҵkp��F���3T�=�C��m�s����э��}��T���-�b����D��O?02��;o7�t�����7�u7bb��B��K*�1K�Ӫ��c8��8omL�����.�^�W�n���n�����PN
/m�}���dt�{Q���j�����r/��VLoPu�C�mC낦ݣdO��N_mN�0���s
�q;m���*�ǵ��J���J���69��7��6�n�)1@�:Îq��=�R��:Ⱦ�W��bzk�Pz�Gs�u���a�G=w���;4�Y��գ�-���P����Q_�f�oH��6FfT2�^w#���q)�'H�g�}�	��g������x���n��z��c\J�Z�3��{�����ܳV^`��TU���El(�@`C��9���Nl �w��O���=�X�c��}9!+2]d���߫�}�^gǢ���f@}�\�g�9%��U�v���l�K�\@O�p�I����\�U��
��c�V:)Գ��Vb�XI�m�����f����Cq'B�?}Q��5��J3���]�V��K�n��7����Iy�Mr0dO�/]F�/u�o��5��?�n՝Ues��j�Jyoy�:{�)�Wl-='���bj��[�k�Ļ������S½�b��_I5��Ʋ�+�3��V�TN����,�me0�{�"g�Ϗ	��'AI��OM������&���p��ke�u���4髆m����O}P�Ҍ}7q6&.i\�쑝�z�'�]��9$5^��_�3��݉�(��j�rʉ�+]в�v��TM�V��.[�x�Jy���s���
�W[m�+t2��!v�W4N.�|�ٴ�*��ݹ����엉��s��O��j�Y
�A�X��;�X�&z����7V������E�t��c�5����y�W7�6�MF�MscV����w-u]��Z�ƻ�R��[�K�W�
��,�:g!� y�-�/��S��1l�[\�2WP�[O�K[��8�,�s��7rWk�&�ߠF��|z��5>v�3�Z�Q�w�sp�2��uky����k��;��\5S��;����*	2�ʲ�:���gE\!.��6�*h�Mћ�(@>�菢����mP�7�ݜۀ�U/�,�O���m}y��'*1x��|�n�%�)� �l�
W�����nm{���{�q�G�[�W���X\�mV4r�6|��Y=G�o�V���j��mS�k�Z�iײʆ���G�����yK��� �7���n�?:���Nw��ɪ7�=�t��]���MX�R�z�D���+��r�ҳSwэ>܊y��h|�H;ђ��X�r�7�G&�J�*�눚�֨r�/��ZSˈ��J�$��A��lSU����a�۵���{O"z�]yV�¯�&��ν�_�z���ۭ�oSZ;��7�Sw�یQ.���>��A���A�o���߻s�)J�wWs�-+���Ӎ�r���4ʲ:Qbu���k}4���eNm���un�R���
���:F��U�>� v]��L^=�\��ˇ�$l��+�2�ꜞ�Mr󮓵nץ߉�S	?g�߫3�F�Y�i�=���]Sw��ӶU%щ=Y��ZAq�X��;�T�WY���#�ds���!p,�qj����-ڋVB�Z�YS��Q(�u�l��T��nv~���!k[2����Gj�OL�N�.̸	�ݺ����@w�\7
`S�i���W?B=[[;*u��H{����;Ϣ��ne��,+�a�}N�;L�7��^�涱��;�觹q1Nю!�m+_?*{e__�|:*�c�|Ƃߑ���y��3$^�P���'�a�d�ٰiu^b�zf1`=U4�s�u�SJz1�ݗ�ye۔jNo�ճ>=��'�G5k�vza��KV�l�s�3��s@�۽SϗIqP��������v��/,Q�_m9�.{��n��?:���]D^NV'��A���žGqݜoh��|vf�#Y�b|�1=�y_w_\�}U�k��*29cٶ�S��U��g�*[�F�f6n{�{�$T��gEQ_A~���u�������-TՔ��zە���^6�k��Z7c�&�ߦ�[,b�E������h�wĄsR��UZ�:8{��1�3���&ԱOw�}��^�*T��L�X5|��-m>:|��2��ĥ*���ɛ��I9a�u�O>��R%9bȫ���wH� ���3%a��N�rI6��n�1�v�ua�9�n�]������)f�D���}e��H�܆�T�e��݃�T��LV)����w^o�%�\c#���>Sώ�\k�QS���}��ڈ*�_n�!q���G!�B�e�R{���Ϝ�b���+ί��e�ִ=���[���K!G�Գ�uec��.�I�φZ��~�ЩzN��ҩz�R��y�)w��`Ҍ��Fn�P0%���韂}ve�bu����'���)��8�#���{T١|���~�4�j�U��~�Z��>̅W$e��:z��}��n䍚��T��&k�.�{�j�y�3�ss�ENڤ�
rG�b��t�������TN_|���W������e����WC�3��Q٥&�w��y��g9�{�Af�o����zG�=��<�-�p9p=��]�yH��K_^3�ߊ���=�7|�
C�v���48UD��B-�4pr�'����"�X��R�l˞����.��Qnx=�0�}ѽgf��嚐�U���{�0K��A��X�u��Ι�G-�����: o�'j��+I��M�w�9LB�or�*�p6�q�s�═Dcܸq���>^A�)����F �H�8����ʌOMj�t��*����5�J���Ұ&y�n�|.c�̯�����us�`g�o`�Xpi����t������p��\[�]�5���^j���V���]E}����!�� �I>�|���eV���aD_7���kq5��a.����j-U4mEJ���2����z{����e󿴭��M�4����^|��@�u�ՓkmnL��͇I�s����19ʬ�+�ƫUҞ�.O�>��4A�Oh2��0��/��1��<&�0�H+��I�w|��s��>�+٭�۬�TN���6�3���eBۉ6ᖚˈ��[��1n�wP�����m�8M�i�e-fm���rU���=	���X�ml��=6yy0������:u��{�^8�Qn�M$:�}��	B%�����vێ��
\�c��d�V2\�Ŭ�h���v�Z�����ڃ	ᲽS���P�v}ՒPঌQA�C��V�yhh�EM���y�=�8Z�4��-{)�Te�a��$\7����E;��;]]ֺs7��G�v$
}xݗ�ڽ��̸	�ݺ�
�W[COa��j�f3�s5|��:%���Dms��ރ�����6 +��a�}N�P��*㓨�o����ck"�L��=�}qAUI� ����=�3L�j�nqZ��	0u5ٯ���mH[y4wk��ĊC�d� ;/�1��E.ߊ��K�Nw���y[a�B�$R�܋���m����'8�+O�K.=>z7ٱy�����^�SK��I��l���p]0���[r���41�n���7)�죊���_k������$~[9��t���WJ��oB�k��]�{���ȫ܉�^�WC��!�YQ���x{~-����ֺ�����*����&V�3��Mè����<��Üs�7�賎��r�ҳSw����y���]^l.��{�{���[]^�N�6�_T�Ug�Y|�5J�Ҟ
�nY,vwcދ;4�d�#x)��wq�2�ҢśYȳ�˅���,���{{}P�d�x��w��Nլؖ��d�x�F�̰�wZ#���ȳU��+�a�S�;�Žݝ�"���3P��Cm͖:���[�����&�}������Sp���D;]_r�[�׫��K���I�ͩO��-w�>�Ax8�ɛR��Q�c�K�k>�m�D����(UPʅ����)F����ݾ��}��;Ӓ�]�+R��������I����?'M�e_�U��Y�!T+�㫣b���α��9;�]?Ef����;М-�]#QJ.����gq\n�r��9�}ˆ���<ʉ٘U�]�p��TV�aގ��VG֋v���ev.�B԰D놶�<��~���̿���c���8o>[�<�i6�VޜP�=A�u�ʦb�٥��خËo�]��au��J,�v�UBj\p��������}��TE�*����7LԸ��'z�h����;z�QUm�N%Ƴ�ۦ�vfX�{� ����>������ki�爮��X���n�IqOQ�o*i�Q�یJ�t'gF��[�W��9��RQ+O:�]B���W�D�촬�`�+kc*[|hn����&��/��K,Z�6��ͥ��L�\�r���d4�5�����r��9�1�g#Ў�/��{\F�V�x�;}/Q�fh��;^�Ԗ�' �B���z#ﻹ8<��MO�U��ד��7�Tdu���5b���}4(����r7��g��@Y�v]��뿆������3�[�4a�sN\�$��{�\�ͪ�[ک�6G��;Q��B��,���g�r�v�_)�ّ�l��UZ���o5�b����a.��M��j��'e��u�B���2���N4�Kym��-�5�*���%#\���|�9R표��W�b���oW�_=T���C�l�DZ�W*-0�N�;z��~�45t
�
�B�=s���t�<\w-w^�t�.\��s��6�;\	�*�A.k�\gM�t�k�o�ח��y�4R8�I�Vk��ޫ���4�(�_��_��3�
�f���"cP?"�$I3}�>�,o[�������1�CU��YS���u��W� ��ōj#��L0H�ii/�������9�g]�&}W3d�ʸ�/�4�
�MW^6�d��5��ØgU�����]�V%��5��n;��P�qR�����A�R��7Ol=ʺ;L���b.0_
׹�]�H{#�8i�\�kr�Q�c��V�r�p�.����d,��CW�ûHQ������J���]�ԃ���,��E-n�c۬�']�O-#�סSx�C���wf�",�Z�/ ֋��hgc�k��j���'u˧.ɶh�,?�a�!�5���X�@�ʎ�t����`C�-Wb,Xj�i
��n� 1D��e`�E���p��ØȞKWq�&�qEv�0��W��od�v���gn�q�=����vd�P0n��
]���t�'����:�Vs}�����8)n�٢w�K�-en�� �jn���@]�l��f�w����ۺb��=���硚��&���k�F�[n� s���\����D��預��i������U�kT/�\�;CRY�Ԕ��32��������E��uP�<Ѫ�Q߸3�R�f���[˱�q��[�L,��ox#�������)��b+��m�31v�b\�s2&��yl�WRK|����"���ճb��)>ھ�;��S�
�X����y��U�Gjˊ3�������������Y�kÏ��p)�w:*���Ť͸.y�}�r�����m��\h�;p�I0]��(���ԁ�t��U�D��ns�y��y���<���ھX]nZ.��,J�:��60��m㶲-ɦg<���]>�t��b#���؅\���N0�^iw�Pj��f4r'6�Nhm�|��B�J�:\����G ���ӲgHޕgZ/q���,�*��5��,��-k���Ma�Ɏ���̇_z֌�,6�̖4i��踴�f+_vA�1d�[]XU��orN�km-�����r�fT�D�\���v%�J�WX�{#އ��H��-a�d����rZ�v�ץr��H2���:�X�p�^�mԚr��z�k/z�e��
��˩[����Y!��NJ�Y8�V莺�ʸ&�8��9��۾6���Y��*6�b�
���1�[g<���[�ҊfT��rFky�n`�]<�V��-�.����+�D��e���ˣ�dᇁXp��3���v]w:��vlj�RT�YU�F�<M�3����R��ٮ��N��M�p!Ie�b���M���/�)�R`�zz��כ�p�i_h�4�+KM�qu�.���W��J�ɢvwX3���v�0��Pg��M�RX�{����Ƿ�G�)&�˃�������'.L.Ṫ�����Mm�G_'�i8��P�6ܘ%|�`��^���C��]�Tef8,�Wj���
K/[�,Vw(�t�1�)o'q����nY�N��Nl۰~$�F{h[DT��UdEE�0F�6��UF"����%Q"�@F�cڪ��YUm�TjTDEU*��ZP[lb+%��J���D����QTTE��UE�#�T��"��D�"��U`��
0`��UTkV,QX1cձ\�� �5Q+Q���*��j"DUX�rʌJʪ��A�QQ�����V��E[h��6��+t�����Z�EH���*�
j�TL��Q)��,AeQ��U-��F�U(*��1Tc#��mm�PTE�mU��)iYiDPE-���ʂ**�e�#1�TQ�j� �0pΚuw|06/�����7yt$QA�xﳅ%Ck�cs���'`��2�e��}��n-!�8V>+�TPR�N-4F	������n^�����nभ�&{��:�������4���)�U�:�.b�I�𓗣�{��Q��;�P�ʸtD�L�/�ڋ������V���vUn���u���;�'��
�Hu�z��&�|��C�N5��BЍ�=m����w:���ʈ��W�j5h3��WoQ;��w]��`1�|������UB`uӑ�_WQ���]�5���l�^���t�;�c��@���R��]�����N)��Tb�nCz��F�^e��sV�T*b�1ŷ顿6�����5���^������z��G�͕=�q�����)Mc�n4)b{��v�;���Ya./0q��g�H��d��z�׿����s�}�y�>��6���otn���cl��g��Jn�h/�l��pbu��ʬ�w�ք�~{Ϲ��1A�υZqnnȎ��1��DɷV���|z�"��,��fI�Y�Hc�̎�ofi���;ʳ;��}�ݼއz�v$��4��Ǫ`�N)q��b�݌Ǚw9S*��Z���x����@����u��Vs����v�wK�o��g�X�3������u�ʹ�gd��[PД�B͛��LDS�2WV�U��]ŗV�9�(���먍��H�w��̌���],�\*-5��l�OVs��z�Jsx��J����+�ù\F8ɧI[6ʌ	w�9`�hOC���B�����md�O}��VhT��'9�g��:�5t�5�!,W��&3���skp��X�p�װVҿ��:��Un�"�'
���{S�>��oyΐZ}t�;���b���]��;��F�j��y	�oq
�0��V�n-%gT�]᥵�LE<+���ΗY�vw�
��%~�M��/b�5�4S>>����a��|W�.ڼfc8��|��Wͮ���y�J�
�pv�e:��_<�O���m�:��P��v�g�aO3"uG<�X�IC���N8�ֆ����_C�7)��8����î��T�$���ʬ�mfU]���s��O�[��˪,ت�K{Ir;���Q�^��i��-��[����J��Y��wD�H4&�v��y�e�|��:0��$,a���P�o���a���k&�W��r�A�ά<��&�R��#�*<E99���6[Л�0��]���ﳗO_��Q����7���\�����Ȗ��;G8V|�C��u�R���P�'X�_ZT�r�㋴���<��S]Y/<]�7�c4�t!���͸d.�ip��n���l���V1��_Gt��������&$��iy���td��zM)AN��MA�j��ʢ�稭�V���R���T�Jrdڮ�ۮ��S]���P]�aD�E>Km}�+QdX���Ϝ���[�o%�Os�{QSu}0���wq�e}'qXs����j0j�C8��X�v%��.�m�6���q�2S��2��'72�K\��{�\jq%N�s���V�}�	>A�ۛ4��,��)�M�qs3lp�P#�T���� .̸	�v�[��Gk�XU;�2�f]�t�>����(����C�W�
�tOI�:*��WYN7��nZ��R�k*V��u�ȱԊ�~K%�Q�oc�T�*�5f+7/��{��gV��a�c;m1���k`<Z�ܕ��ያ��%���ǱC��ٓ������ޗN�1��tZ8��컊���D�>��S�S[4f��ZF�<�:�+����,���s�vŏod��@�ήїͰ'T�#Q�.5�u�*�����XU��ق���\��7f�`��X���ފ�z�e���^5;�}�:������/�믜��ʨiKmE^��{8�=�W�k^�1��齎RTbΨnL�V8k��:OUv�2���ހ�R�C�8�֪�}���T������pu�<��9���2��j��"l���~�YZ�<��{_�cO�ۦ��luLꎭνJ��s9�s���ݒ��Wt^fۜ�g���G^t��u�)nh��H���ҳ:�3���y�����hꅘ������ִW^��oPz'1�乢�^�����1��lE8نi�OWM�k)��_=�c���v�<��s ��([r�N�2_��n2�n{_\�����H�ʔ���ņ����piE� �� �\�� L��R62w�C9/"\3Q[9]#Z"eq��:g3s��KG�OwZڛ-�&j��f�ZH7f��]H�ZD������=r��-ᑓr&��BX�����h�yY`�m��؉������%���/}\=��?Jq5����z`�'���z��]��<{N�!dl{��\�����g���s.��.����q��J�z{D��<���m��>�L�rʸ���D�=w��w�AC�����)��~�bْw������"��P��᪈���Tb�]d�R*V$��D��-b���c[�e�;��3e�u|݉���B��4�65.�{*{vJ�)r]5�'�a���I:q�C��ཆ��m�\��:38����i�{��ޡ��I��2���~~Y�}��:���4�K�j��央�F�:=w�$do-��o�y�v�7�������,'V���s���eYnz�|׵�W�P�;^ˊ�j>\P+��c~}Z*x����v26�o�v�+O��C�s��y��Õ�@nS��_WW9�np��!v�"�r�0� ���E{���S�ە ^��**�s�hܼC���T��r�9]OVд�kdU��^�K.qw7#�K3ޓ-@����&��*�ޤkrXR�6�|F�]ڻ�8��E=t�Ɔ��uh��a���2�)*��j��7uT�c4�e/꩜��>��zGY?�R��ˊ�oE�ޭu�^������U_l��"F<�fR�˖����
v_�z���-�qD�_<n��Ǹ5������ɐ�u��3m��;�A�C�x��c8f��V_+Ҷ�7�����L)��q^�k�V�-��X��q�1*��D�\�V9lY]�O�;��= v�-4��5�<��v��?�k]�6�И�_�m�A�R����7����|e���+h�핔񦭽�ޅ�HΞ�t�8v�+��*�tJ-���Q�G���G$}�QY�7��w��wF8ɧIM��_	TՕ'��n�VJ�5�=���\=���w5�\���m˔����3|��*.>�XZc��>���^��؜�3��.�М�w;S�5��:��V�wF�)<q� ���Iz[�
��y�C�W
Ս�o>*�7�u	�;Cؖ��Fo-�T�Ӑ��Hjﱼ�2��S$���MWU#A�œ/$�.c9�((�A8x�#Rꕶ$�}���92��ć:94ɓ��iU�ܳ�����\��EowjR����Ѥ���o�҂�e��i���y�g�#��sT؇\���7k,F�|\�g�#/�:+��N�:�<&���j�����o��z�b{�Q�N�ikz��.��!���j��#}�|����Exe.V��RҞ�>ַi�]����;M�8T'>��~�����N�^i:bNc�f�����>���`�o'91uz�tg�{�����rb������b�K%�ճI��]^NTb�z�zTf�p�n��c�^ظ�KӉ�v[�*w[�c�:�z�YL�x��q���Q��켽�J۔���<&�ٶ����RP9���w�O�%~W�n��J,㨷�J���a��:�-^^۷Ϊ�J�Nju$�b�R�9_b���_�6'F����}��y�;���r�^�ˈ��njMvE74��*:1�|`���>��;S[wT�1!�>�I�R��@�ش=Ά���Sw���`����j'��C\��}tn_ڕ�;�\5�Psqn���l���VU߽ʷc�wٮzM3���$�{ʳ�a��rtK��XδMZ0��eu���Ú��"{X�B�r�t�[N*kq�4r���p��'9Ǉ��ER��B�J5�B���ov���)YK��~�ͩΑ[�����W�$�{u�9~=�5���.������4v�Έr�Dq�r���<��7w�h�:t��ui���_OK�V��]���{�c��}J/v�])����Qx�����`j�j���-wpfXN{u��O^m�����v9V��sG��Q
��:���y<�U.]����SI�wc���(�1������3e\u'q4����;p.�<<�٭XNz��`�WS~��g�U�����v�&&[�nેP�D�o	��~4�l�$��Nn	v���K�<#=��z��C��������=.�7'����rrEc& ��z�vB{����
�?;T��T��Κ\41�z��]�BXڨ�8��*���T��	 �ב�[�Qy9����pX}��rY���ӕG('���'�ZA��]��>�+B��>��K�y��k����	��s�CB�2oh$U��p��&�1��m�W���k<���x�v��¦�Il�¹k��WlS���Q%���p�q+;j���ڗ��BÓ��G\[�d5�&vSs�XzB6�mq`=������w��W�G9s�|ɬ�F����V��q��h��v�/0qU�\⯬�cL�B���\r��E>��jR�݉�
�M�i�w��j����ruv%p����<�+k��\��e����x���i�-;m>�Oz��x�C�Y�;%:R=V��z{�ӜQK��es��哥;p��Coh�sUK��]Ɛ̘�Mh#�H:�EB��lT�/�Ұl��N�3�|C�Է>�����k���p���&<#_ú^�zy�>�．�%�=H�zTr�J:�:�5���K�Z(��`J�������'�4���B�L�O�'_؞�N��:��V�E$#!�k�W�.���0{��q��쌩�z8���]��|�KWV�!�'���8�	m��0:j\Vrq�N���Sz��X���W�!dBN����Uï���梔LԳ֩C/�aܸ��Q�jI������<�sEց�"烘��AT<=�׏�_�y~����� ��
}���52ӻ����0���؝�uOk��^*�J��,ɸg2��c��701�]���`����==�u��!��4蹮��[� ���c�!𿈨Hܕ3�&0u-��5�.�=�Щpp[A������P��A�җi��{�nm��}����Zx��q�T�ޕ� Q�U�X�>�r�D�ȼ�x�~ՠ�&�S��=u�<w����!��	�8T'!��=G��[2�{e���<�$a���{/Zjvo���M]���:��j��tߠ������to��+�"z�nj��v�\_�NS��Ηk�YTgT>�+u�H��?5o}��#�T��Z�q޽13\���p��⯣c�����Q1݁�����i���Z��p˘s����n;9�����V_R������^����������vd}�w�+��ޛ�&IQ�BU|��Pu����犹}�<�3B�5��N�wo_��^g������ ,ͯ�1]pT,���2�M>J�%rƥ��3D�z�tS�Ɋ��C�ƶ�.�����/��
Y_)����}�sY�u��i�uD^Վ���ٶ�s,&�|U�:v�B��3�U��
�@����mj�����`ׇ��2�|�n�p{t�[�.����n54���@�9�C^{Wi8�Of��J�?:`Yb6i�nk�2�1�}O�WH!��hWwN�F�]2#���l[C��VV7N����8�3\{O���v���ft��Q�0���Ɖ��l�b��4�".X�ﻂj��Ձ�(��8���c����c��4����:��g�<iZ��V����i�Olow����諱���4ts$.�����1�s�E�m�~";�PN�[Z٧@���N���,%�n�Y��v��jV�j�Xx�ԝD�DݧW׊��x��T�mK���L&�i�3�Οm��m<T�c2ಱM80#��Ϣ�hΤx�jt��N��ۛu%zFKIt���(��.���¥%�q�O8_i��(�P>�cD�
ۑ&���U��W{i�.�c����S3q�b��Ke�Kakn����2�|1B�+폚�рo�왨j��S+����v(�17/�Ӳ��&b�RC�JmK��]t,��J��wO&�Z��S�6MM8*�W*��
�k>�W�)�ۧ��6�o'��@�i��^wQ�,�\�ٜdfP����=$U�� :�.t{���W����7�]� V��	V����Ci�)�p�� N �삥��[?&4�G'�]fޱh;1���I�Nj��p0�C5�
��c)ܥ�6��n�ɩ�9��_�g�L�O]�<,��MF��_^K�򠘳6�vf����OBf��B�(��۶Z1vp�������Wt1���VEu3Ưo�^p�������'���]+:�[Y97Q��Ŧtbu�Q��}K]���TZ��h\nލt�G �.�7� ����������'��������uY�u��J�i��#�aCjN�lh�z�$��1��������w1*z���4�g1�Y��۱�v��O�"�b�=�ه���-�6���B�Ouaz,̧j��<�HJ��� I�у`���]4@բk���";�[�y�����eޙ�ݷ,�>H�$������)j���7�^�ԛ�;j���#4����W+��Y}E�oU�p�r�KV��z
n�v��}�vr�3nk|c`7CR��Uv�Ah�\�&��Å�q�E+��Ѐ�6+\X+�1n^p6]�:�m�չA� ծ�p�k�X|�p��Qd�����	�8�߳��!�=��&��[�G�9��`�[��cJ���ݨ�l���u��b�-gLnl�*�ceu��Eq$n��0^v�F�V���]�;4���W��g*�.���Ԇ��Ɠ�BS7|��9����Os!�Wu.�no�������'; ��Y|s2NN��f�1[Qt���ԭ����S�N�g+.�*�K	L�3�&�t)q���CU�du~��r��N^܍όy�@���qc9�/J�p�{®6��#y�"l@o���WzP���߻�PU�ְX��[*Ŋb�,QU(*�B������c�ֈ�mE`�WhV-B�h��jc��*�b��T\ˑY��U@�UPAV��((�J�*�[k�����V��� �[0QfZ��DU��q
���QA����E��ˬ2*(�0X(�,b���QR"(*#��DdF*�Q��dDƈ�@PX�b�m�E`�-J�m�Z(�,Y���+iUU&0���k*()X�R��d�����@�1X��j�$ƱH��)iX#���R,1�D"�@F
V������)
���DP1���6�X�D�QF
(�D�RT�)(��
(��r����X�@| y15�<��%�e���f�2VH��o��UZ�sX[g�X��:��(.��*:C+��DgA����T���v��wjO��ѩ^8ɧI[3nW�}�������)P<�떣c����o0=������~�r���>ߨ��og�H$�秼�,1$�r�M��2�Wn'A��.��	�ݺ������P��+��o\�`���c_Ay��A�݄{���j��7�e=~߻�|��8�n��F�����r�ܨ���*f8��6���)��9�Yvtj�d�qvOrW�F���Uꆲ	�H�5L��4�o�o*/1T^3ٶj^%BVFM��X�lq��Zx�uݫ�T�_=Pv�nq�b��Y~�=����7�b�M��~��Y0�K��o�O���/Q��n�t㋍hm}v�:�ϟ�Lkf����)��ͧo]E��b�cTgݔ�g��~�~\|.6B7�����D/����g���<G7��b�~�{�ǖ�Ր���'��6������7D:Jg����.�Gv�S������X�����h�~y��ڸ�F�Թ�e*V���b�����V]]�:�㰳�6�V7������zf�Z/o+m�{��T����("���ƒ��>�Щ�).�h��Eԣ��P4r�(��4�M��u�g��T[C��������/T�Lr�#��<�������T^�-���nmnU����ǹ��N
d=�a[�����"�ljObk���Iu�N{Cv�=�Kx�ܽP��,)�<�Ob͙�_��H��fu���.=b��L��O�P:�����Z}���Ju�G(�	�ENqߟ���ɞ��3�Į����R0�D�ܯY�yE5��7ˇ?	���haQ��06nx�7~�u�ɭI`�.7���M�*ْ+Ҭ��h�6a���Xoґ�\r]>݅~}�u]�ݨˮ�h���ё�F���>spH��Ԧ�|_W�����0�Wt�܊��y�i2\�X;;'o�I3�+�y�� �=�E��$o�t<X�0|2�j���=�r~9��hɼ"]{z����:k���m�T�=�����[��\�G��K����;8�w�E;w\Un*�q^��)4��G���@b��������G��yN}� y��3�+�U��w�`6�b]��N�7=��'3�ry�?WO�C���;�֭�Q�v&�]ґ�<G%��Z;wg
�h����Z:�Z���$9�8I@Ν$�s;�vv�Σ�>սa����/��v4�0�ʫ_N,�����T�Z=��z}d�t���g>����*'���u��|g���Sn(mV]�61��x��Ԝ�uGmZ�1���zj5΃*1pcާL\CUS�.=���={�����Ư.{9k��Hq�ap���:n��|r�u��-�f�i���zo��&ջ��k����cJ�{�5��u�i�y�"��ب��좷���e��څѓ�szX�k�K´�����M@�X��ճ���ϯ�
�{��W��R7M�ŀ�g�g�+/\��EQ�z��kc�}�0ߤo������L�5�^�F��'}q��j�9�Il�:u����|�z��E�W��jۧo�q;�EG�3�k蹞�w�̏(�/��|���;OǥyE�h���Z}^5R��{�j��qW�!�.-M���V5<�nS7�L���G;��)��.�~;q�6='z��K�$�gm�V��>U����J��G@����^.�mCF��mC��t�7~y�˻�����'���<������,�6Ks�X����� l�}�0���[V���>��i��z,��d��;	^�K�l�n��'��wZlR[9&��ݨ]������ͷ-�籑��C�(؏-pz���]�s��QX����,�1�*��m�ΏU��ub��O�^q���eMw��Յ�yɅ1կ9�k��Vlx�tgu�W~��OxߛG�3��8:�M�����#�у�9JdI�z_{:�w�\R�ͩǵ~q��yo��+�_��L>��_�G�q(���]���"��9 y��* �A�������r��ߙ/�i�xs��%�C��%�S��.�9��5�sJ++�9 T�fkŕ[��9#^���!�1����aw��r���\2�ʉ�Q�S5���(�H���٦��3�G�ae_/@'�E����K�9sjU��Qml�{U^+��c���&��6/׻��K�lȬ-͠�'�*!�Ƕ��xj/1GW׉�=��Ls8���	J{M�p|'̭��K�'�o��?�H���8�i`q�%�~|n�D{D������rnqj� 1�e��w�� �g�2���[�i���g}�*&��NN��hO�TN.�-�TյפM��UK����6����c��kK/��cq<s�rOƣ{�2��1_>��I�� h�.l�Z~���z�q꙱Tfσ���j3���!�F��>���o�ht�/?f�+��Wh���H �2q[��U�Ѭ����:1��7{807�.�K��om�\C�8q�dM����)�H��ܺپͻ�q�fGq�ϸ"/h�Z9��֔ҙ]�rW
�у��Թ����W`�5j��wcG�M[Rh��s������]T����A:��Y�ע�����%eT{F+�/�ɝf�g�<��C���;�U�{0r��3ެB�	���g���^��_���:��EI����XZ��3�53�������5~�b޵��*�(ɶ������u��C�V�)�,�|�DS���r(�����'.\
��"�~z��g��ξr��b>�~w
�u{���}���O��]���ԫ�X &j=*�o*�d���S[���v�
����o�C���,*���7�l�G�T������G�9^��|tKfsOO:�s�7Y�ü�<�?UHd�>��\�϶X�գ��y����C<���G����; �{��obI�tX:ό�R&&�W���KGvGt�7]V�A{^yj��i^������[�;�wfA~�nQ>GI�W�1?E>��q���g�a�^�"�}8��F�Ֆ�{�}2�K�-�� ��~�1s�RG���3C���#���IX{F��t�U�Ì�9���[AGTk�4j9��������%|�2z��c�M/"/���$Ćp��P��Uo��N`x#{9�s�y�[�����ԕ��7�_('��i�A:΋�u^4X��b�BKh�n��xiW�'s��P��b��}`gE'e�o:]@�	�s��΅��p@gq=���㮘��y���h���]L�JYnc�$v� �nv!7��WZ^Lϡσ35��UU��T\�=p�M=uZk,��|{��?��������jΛB�����=C�9�.�p,5������ww��@�>9<�M�1Q6t��'��f߳��gFĝ<tz^),�ɇYZzX����8�oup���d� ��Z]̎J���'�g/5/^m�	�'��H�I�:����Qmm�ΐ3�T�2���}��xtcH��^Gy5�5�~����#�E!�&YޟV�*r(�����L���&h߭]F��7�׬z������c��]�����v��xכw�#˅ �5���\%@LV���[�DL��/���c���ε��lÏL��o��C��<�ny�x���7�\nG=���uLۧ@>��+��~��^ޟ����G���y2��U�;�KGC���*#��x�C�Tz���ts��
���9��.�6\���UHʙ~ Z+�ҍ�竇���t����{5�����s~w[�(�yA*��K��Y��(�Z8�{�`���IH�S�f����>چ�븱n�I��Vn<�.�B�Hi�ߋ�h�s�]*�Y��S"�3�z0B��^�eF��xr�Ɗ+:�_`e]��98r�ZE����6������N��#�KtvZL�¤.WJ�N�-F�v�n�ፙ���N��2�`W]��͂()���Ü�����`p��n�?O���'�l�ٿ�M
���a���a����'o�i;�Vg�&&�Ƹk��|tz!���]�꜑~t<X�0|1�#")�i������66�c�����=g[c�S6\��Iȗ�~�b�W��2CGzn�މdozB���$���%V.^!�=-���@>Q˰�6��s
!��%K{���+�+�]+L��w�"K�s�픴[�<���ʵ�v�xl��8��\�Q<3yQP�!;/��q}q�>��\M���O��/G���6�R=������W�騍s����	�����d��x��T/z�� 5�:7Ra�8��G��[���՛�3]�L��� Ў~�6����OۛSU��L�k<E���:qݩ����#�\�g"rx]DZʏT\�T���B6b�}⛅��zzN�=t�6�'Ρ��*�F[�G!��n<�AS,]�K��_C��gU=TWp���8��9銈�#�j>�!����gt�7�c��F�����6OqҸ)��q�%<�b�g����\�̒@v�"��bY��.�r˛�ķ�+���`���ujXV�\���JE�c����L*��xC�/k��� �A���1	gG��.�/�0�)�Ż�Q��wۗo�$8닛�����OM���X�kf(�P�}��p���/�X}��.g��~=q2<��|X���qԶSu~�}K�ِ�w��P~�ї��鎻�KK�l���h
w���j�X^��xX�<�z2=�|�o]�]kYV{\o���i���v�CӁ�m�	Ѩ�욌�4�V�x�ͨh�_������pЬ���P:�G�5�^oz�p��W����\ ����ޜ�#+�n�7=��"��R���]�a�k����ڍ�]i~��g}_�܁q�W�q��ȁ�⩑9�Nm���\�[5,���{��|=��'�U���u6|\��p����SC:g����K���n�}S��6������K��k�Uq3J_����Zwc+�u�˟'1��s���7�҂f��m�U/�Y�({��$z�}���B|���G�%��m�\�wAb��^�?Mx�9�ވ�L
��ٴ�aK��@W�mT ���7���ډ��9f;m����꾯�+�1b�>�gϭ(�1���TR���2��.;�޲���t�>|q̱��3Aᨼ�y/����!�u~}k?T���^�1��f��0�A�*�R�X_>y�����#�Ջ�;4�� 5���q�s����S�#�3wY�dl�q�W����{n���q��W��Fוyb<�WtN�XU�T��Y|�e��6.�̭3D�GlN�o��ɻ�I/j"s:��ts9������E�:�ȷ<������S��u"=��rx][X:G�%8�:�g.���e,�F�&�N���8�&ռ�&f����)�X�*&�9�N�ŝ�A�ϔ��?%��^xK�]^��5���(V��#}7��wae{=<�^��s�Z����<c����6���9)��螑�{"��+&����}�@�uH��� *�v[�kF�J)��p�O�����"��Kh�����O�t��ET{b�c	�z2g�<��u���L�v�h��!����Ɩ�l�Gex+t��ݤC���N�"j0	�����o&X^>��[+��d��Uyg�8��	�'Og��Lh�ʭ_�7%�~�%?����6����SU4�����n���~[<�(w}0�t�ϟI�\r7���O����Ie�>*@[Z_�nٵ>�Ts�n����k:߇8�-EO˸���Y����6`e��.f������,Y��/Gt�Nύ����j#܈��g���įg`�L�<�pw�q�9���� om}Ó蕃*�s���@���B���
����Ew����~��/ܰ���ڶ�f���/��5�Қ��*ӝ؜��&ȵ=�<���0IۭmkY�c̮<��>�(.@�/t����Σr��t)�׽�V:N�ǝd������0/�L?@B|ȁ���T��}>ÿA-�ǩOq�N�]�t�z��9�]��od��(�z�X;�*�:��"������d�MG��14����a�w`�Q�T+h�\��r�{'<��Ѥ{G���W�<�hs`o�`T[�\�^I�m��2����57Yt�v/;n�b��Ϸ���Ȼ�tu}沍F��x��Z�h����4����3*������*��9��&�g�Lʌ<����\o$\�=�S���~��F���%�����?�T����r=4��h�<�ˆ��9���6r1�Tb�=�p�����q=�5��aM�w�T3�i�XZH/cћ�)��9�N�{2}ŋ�8TF�}}L	�V��������=�;X}�guW�x+�?B����-�mI��������e��j3�ꎩ�KPk�Jp��,ox���^�eW�\;�����>6�n�gn}HiS�}kiq5�����N��0�=�q��+��~ǰ&Γ�����3��u����h���$K�.� T� �벵�;�fw��jN�#��4,j��z%�=�O���N�@�,�C��A:w}/��A�cU��^6{|"W|�a	*�:�:"Zn)uv��o'�X�4���vb���6���[����Y�WQT�~�t��	E�}J��f�KU9�ٜ&ni�1��(&�.���Bt�{�ui�aP�2fE�U�B(Q����5�i����q��@m�m��������w���I\���6���U��|����%�Ŭ�6�[D�7S:��c\�Z��	Ik�i�gq�B�E�x�zn5Z��u��k#Y�{eɂ�V���,_!��	�$7���rby�ը�UĬ���q�W{�1�Z��|k�jf3�0���apq�K���8���qS���Y�>���������9Z/��k1���\pZ��˧*mKsuvN|��������]|댌+ @|y�L��2��&C�Iv�
����,U�e*�R��W0���
�T��;�&���wz*�qPf�Ӆ�Db˱�^'�����_h�뵶3C�v���-c��G'�v���;tC},��o&����ε�jwR\߁��/�N�Bo@ O%]*�΀��p<ډ�)��R�s��<���}�Zr��;[��\�٨0��̓DX퇽��{�\�O�)à̎��T{}	{�wL���j��Ʋ���hWnì���ޕ�7V+����E�Uͺ����N;:�r+�$Q���v*�J��w��tM��5t)u y����]�Т��pE����VI�{�*ܥ%�
[3Xt��[�%iD���&����]�]3Fd�phX5^`� L*���̤ɽ��u̽]�+B�BT�C4�	��w���`@��έ��/m̳���4�R��/�&'F�g]`��2*!�k�e�쫧6�U��ŴՔ���aU�_�,���]㏬��_`��������aQ#ݽ�N�^��X����ԬT�Ƽ�@����w
���
]f��a��x�k(C8L׍o��`u�9X��̟�����3!i���[J�˽+&�mb��4�ݔ�{�����ڳ�HyI*��h�_i�,|�yf��ƀ9YQF��,��a5�I�pa�+v�6g;B0J�_����4Quk������;�o��QW��	��j�d�i�\K)ƹ9�Ři+:S��M��=���l����B�	������]��a�2:\戧�e���n���죎��SW�巇���d2�^��4�I�5��CwO*���d�ﳣ+Z�|�5溹�ݤ]�Zoz� 'K"��kU-a�'fpj�)��}/��+"�q<j�ffk%Ҳ_g
0>	�v���l�cB펊=u���%�C�˹�R�K�;دC�*��aM�����I�]'�6"K�h���y�lMH{3��ȁ�h���)�s3s�b�tXz����� 1�P<�CTPD����OR�("�Qb5TQV\����2ЬAYX8XTXKm"!iJ�Y���LaQT*X*��E�VF���DQ�%�J�U"ň���Q@Qj0J�j*2,m%�-�VGM�Qb1AA�-L`����0P�& �&6څf0�f:�$R(�f���P�U�
��Ym��*��M[V�Q��`
)P�#�EE"��AQATY���H(�X�"`����%T�RQ��%�Uk%eeA�X,Ыm]a���H��P�Ab��CV��8Ɍ
��2�*�-����E"#1��)��b"ŌE"�LerҲ�"�V���1L
�����[lP���1�au\���ܦ*
�L�H*1U*CN!
��(E~��f��|�3�7�26�����:^(l8ut���̑G�kj����J����/f�5��i}�JIb]d�vvfP�EN������Ϝ�SO��Y��)�{��R;�PF�+�ƨ���)��G���Gq�-s��)����ED\�|0�=�����h�ϟR��iQ��t�~�<�h�}k��9	z�a��7] �"�FW�-�*-J�u��«^�Θ�p�g�J�Ϊ�u�v]o�MS�e��+�v=�A*w�T�+�^��	h�26����ƥ���{�<���=[��-h^z|�S�o��u!�}5
0�)�Ā�̣ >�YD�wy���M^�۫Z*q(���:��x��U����=�@�,��#��~� Dcٷ�G�
�SU���Y]��_x�_�a����P�9����3�%܁��,
����"�QZb����z�3ׁb��䇐}�B���"�^&6��}B����1��P}9����l��]�}ۙg;�7s7\)jN���;sJ^+E�����g'���xTo �*!�BvY��ݽ�[�fe��)��ڳ#�[��D��>�MK�۝P��f����k�Wظ1�:c�)�ο`���Юٶ����	9xs뺾za��J���^s�:�4�������"^c�cmV[̨r�`�|�Y��ذ�l62�8��e��l���˓�d�s�
�ӷ�tO��j��3�-��PWr������	��T�M�W�N�t,X��zQ�u�z�}�B��^R@�5�4��Wӊ:�[�W�a�<��]yA�7�`(��:w���݁'9�-�bt�R29�X*b:v�D^��em���|����9wiw�˜���>���e�@dz�[:�Q�}��
��Q�P����>��U�핳}��?WK:���n.g:b�:G�֙*7���ֹ�iȣ~*9ߪ:߶���S�4�νm�y^�K_8�=�OY���{�U�LE�2��L����׳#��,[|������&}�U��p+�Z�:�M\�U�nǌ+��Tͺ�E�}XD�Jf�e��e�W;��uf����
�g���YW���=Xm)��U!�p��Y�}r�`=3����+���4wQ���v�n��3_�y��V�EzwO���}Ν1�v�/�nn=2��NQ��-�.�Z1{��?/\�Lu�4�c��:���VhQ��5�<�Ӽ[äՇ�L��_�7����^4�/O���Cǳ�<�99����<7d�*�Tur�l�9���7#[�F}\�I w����؉��v2x2κn�ϒ�n����2��n��im�v��C��GlJu)�6��Zf�3��H�
��׌K�t�L�'w^y6SU:c�X.��`rRu������6��]ݜ���Uh��A��I���h�[s�g��c��ou�i��d�ǆ-��1-k��9��~L~�C��~��g�s����Zw �R�1��u1�_�TK�h�|����]�^tz�L�M�9��}D�C��ʚP���ɉ��X�gK�xZ�*'�GsTʻ�F�ۮuѸ&��3x�jXʗ>�k�j��ex�R~;sj;.r�u9�>�=���L`��(oZ���{����ܯ&�:4�p}�G��h	��#����I>7��c�������ͯqĀR�zLݚ�=��筢eǔg��w\."7�,��������vQ�q�$���!a��c;�¬�T��f�viym��*-�^���*�:����
/���Ͳ�y=7�=ʉ��l��jI�+��ku�H
��^�ź���8���ur���兆���5x__��z�Ӝ�{��b���Y��@tǈ�N�5G9C<tǵh��"T�:��2�ɭ,^L���@��܎� W��}�~ގ��������짙õ5i���ٸ�K�VET{}��'Y��O��6:���Ț5S���ɧ�\v��;�M1�W^2=��}"\�u8���b����)����gT�mرӃi��U�����Aӯ�4{�!��ϵa˜K
s�<�s�v��\�ξܚ���u�7�M������`�q`AYء<1�uatx��5nn��86w+o��,����/�<�t/2�h�W<��ݩ�حFJ䷽�x����r�_��i�;��+�z�+�$8�g:"�̠��G���1V����N�T.���#WT��ށ���2+���s���|{J�}/��O���v�/"4���ى�b���;>�;�)���K�?ET���@W�(4}����C��m��y�o�x��N�����i�YSZ���^����l�A��U!�U���x�}����;��w��H�>ڕ��v��g.�J2��Ex^�,�"��������0P{U"b~���9�-l�ǩOq�ojQ���ʝ��{�%?Q�����w�;ʨ���^7�Pj{&@zj�&'�}[GC��Y�����=a�D�Ώ
�����g�Gl�h�@=���X��W4@�y&�A�m��D4�o"p�{�$��-��Ѩ�=�Do�(��yѣQϐ����T���9�W��c�D��݊hZ������9�`�ߖW8��xL��<�ffGg�"�+:'<i��8꒍���JU�
.1��'�����S��N�ᷓ����}�;,����d��x��^��G���]�����Cf~�$��Y�ю�+3��٪�X��� :d�&��7�#sO^���ŗi�-6*EVz.��̊�)&E�d�'��Q]����#�9�F�l'�\4f����#���:l�on��a����i������9'9��~��ϙ8c�l�)>9Q8�����¢�V�:@�t�7�[x�C�=��o�+ef�ȓ�6�c9/p����Sტ=�+EǞ��.I�~�J:ʋX��"��5�u�9�o�(D�y~�=NB��t���~����>�-��cږ{'գJ�Z=kj�^����Z��W�~��3���͹�*#}3��^£���Zｗ����~����VU``��]�+�n�"n��d����>ݨڋ�ޘ����n7����Ί�g�9���*�F_���)��;�M��^���L�k:�o��>�+��>��(�#>�h�y2���_�t�����j4�IW2|�>�9��l����+Iq�7�g�t�Oq��>g����s���}\3���Q3�F�7}��(5F�6���yӸb�ӌ�u�2Ot�*ۊ�T�RÄ�}�0�F�b���9���|�Խ�x{���H��<&���Pe��/�I�$�e��ȯ�;9�v�g=*�we,kﾁ0�k�wTuOm6n�����W��U�t�P�xW�|��f�'Nd!	���S�흅�(����_"�L�KGaJU����TG��~��w���6ރN���0�kwڸ���+��m�AHA�J��8ջޝW��Lg
%C�յ6uʑ���x�>�ȈC3���j�oX�due�M�9�0әڹ.�)Y�K��r����r	xR�|�&\k8�%ԁއ��H��'4�tV>�#�}K�Z}˻�j,����G�O��Q�q���r#}AGWrf���t���@����t���=�E�2�m箕��.�i.��)���҇�k0��:O}�t��c֦�b��\��H�/{�� yv9�hW���C{�_.	����~;q:��}�u^'��΃*1p�F���sWO�'�B�/�}3:Cz�N�i	
X^�$麆��ÓG>��:�f�:^�����UK����q�ƥ�ˀ���ȏt�"��Ʊ�T��M�m�g�6/NOSyo�n��z����֔O����q{����֗�Pߎ�G�p����W~��<��v)��S۩�o�P�[�R]]�L�d�=W3�b�:G�k�2�V��A���sJ��Q�b��7�4n�u�ş��'��:��VEV7=���dγy3�^GL�(�/��|���n�ۅ���}��J���ۓ7�s���*3��f7�a.5����VG�"�)�%����E��`��õw�:���XE�t����(���D�F����R����V��:���3im�V��M�GUp�Y�v�@������9F�B��*�=���nNܻ���;�ʹ@3�mq
�����fېjhRb'V��i�M���\�N��.\]��o��C�zv����)��r:�� ����������m̰g�Q�)�"ԯX�9(Mp���u��#�zc��)��n�o�
!�t�\G�z�d��3�������1�e�5���cֵ���h(�/2aiV��k�>�r|}��N�ECj�%ƒ>���͉Z��S)#������L����`,-9���ibWʯQ^/�G�#�=�EZ��t�=���9u��w���z��}Q�ۥdO��tYs�9�g����K^�1Av���z4��K������z<۸*��I��K�웨{q^&)��8ϴ��2��^��<2�Ô�}�}Թ�����*��� ;~f� _>�k���'�6���-f����+�=���(Ϊ�Փުp<��ǃ�'�ik�|�~�<��o�@/1%��U�ñ�P�)!�뚃�@��⮶��>��2f�����xjN���J�H�U�Z�G���2Gaۼ�nez������OP��`u8�ps9'b4��z�ÿt�d���5�2�k�yS���y2\)��	��n���2��Ǫ�
��*�H^_��7t�ak-�}SE7��t*��1�!6`}�W*��/T���d����AX��U�#��nm��N�*(I�CK�\T�� �gk��F�ޛ �X�:,��T�G���W؄�I,���h`H����I�u��t�ٽ]���b��x�h����/�d֗q���nvvx���p�.��6���6�l'�~�I\އ����������;l�E��T�VMib�ɝ�� k���{{i�.��gK�Ue�,���Mϭh�o-�.��_�tSg>�N���=�K�9Ƣ�X�h���S�����O�ȡ���u�r7�>;�,4�]�0��fѯMě�Q*4�Gy�Iq�����7�Y�cXӏyr�q��g�#޹�����r#�+�-�_��[�(���D�����
�Ǧ��y���᪯V6���T\�z^l�h�{�󤍦���w���5�1_zU����3Q��dB�s  �7*���k��3���r����Sɀ�.X�>�­����1��/} l}�/�1G��1ROM'�+S��8ņp�`�񣃮U6��K|`�G���>�šR��xe�{H�*}ӿ�/߶�Y��B���O"4��r�B�����0X{qT������8KGw����[�j>��o9پ�h�E�*f�/���n�Qn�nR�$��?��m�vOt0��#A
�}�F���Y��rku�+Ѥ�eqy�5�@�V����YiFb�!�@k��XL�VvX���������j�~�tn$��v�z�mU�b7.t�3��)��s�)�q�W8�X�kX��kGǧ+սס��sQE������G��:��lS�)���@7g��=_s�DW< W��c�_��m�	��'4ڿE�`��S1�|��ܽ%a�-�/
�PQ��v9���O%���m �Zry_�1���
�ڗ>x���kQ��5�g���X:�q���eFe}���녽T\ž�8Sip~��v�'G��K������3��?IeΌO�t���s�]E����s��`g�_�<1��db/�su��2�ڙ��Z�\�N]�	Ƽ��;���I�ʉ�ui��xf�gH�W �~���y�/��3�DGw��/գn&$'�|��.I�~����X��Σ���B7�s�s~7�[\kʐ����`T,�o�V��h/;�4tG��B�ǵ,�D��iS!�)�1;DB2),�o�N���9�V\3���O3��t;��5/��F<����r!v֬��x��)tb���� ��p���&_�߽ʂ���zn�{M����ʽQ��R\�k��zQ�=����t3n� �>��'�DUϑc	Cݪ�����}��i54�[��lɊ��Y�"Fx�kg=��Mܥn���F�լ��
�)�ڂZR���ל���
u����ҩ�f���4�yx��׽�R�ww�cq<*ü<���ܺ�t��c{���o|��y��QV��V%�վ�&�\\u�_�.k���x�IufD
Rw{Gp�U7�G�׷�gh��>���k��Q2��J�͖�Z���{��Sl��ћ�N�z�^Ӭ�Z�;�9ơ���4O�vL��^�e��5��fMD�`D]����ӽޟF���Ã�)�H�o��@���GP�/���7�g�G&OF�f
�L�5X\��>%#��&�.�p����<�V����N���yPe����ͮS���=^{G8z�^/��nϠ����aC�~�f˛����ր�s���VbՐ���9�=�ܽ	5$5TB�웯��Dz��#b5���F�cV�����LTk�Azk�����ad��Ol�x��zXR���-�=��4���-f��卒�����Q�D��o�U�@�QJ�댫����'f�9��u�? }G��:��E��Qx���s��A�9!�y��7���g �W~���E�Y=����+�O���9�8Ν�vw=�h��W�>]�Ը��c���G̶zn:�~Yn������˄�y�"���Wϱ;p�"��G��.Tȹˣa�4ό�T0ϲaEY�*k�!^je�[���M`�*�gWl0eQv%��˟Q�n+F�;lӫӄ��K�V�����rtΆs��:�! Ƶi��XW��[�*�j&79R�eڝ��+65;�صq譾Ϊ�YGvG�$,Ѻ� XpY���&�G��Ɣ1��I�ḋC/f�w���'-�0�#�Dpٽ�����A��wM��e^ν+�;��*�|+q]�`ƉU'u��¶�˙� j�⑧[�ky�m��੮�V����Z���pTe���jf�V�KK�˨Zc)�SE�7�g+�-�,ܥ/&��qX���7q1�<�����եq�:�BrG:j7��#�%(�RU��3��
+K�Q�7s�;��b���{j^�m���3@{p	e�f���w�i�vm]�%�ݮՉm�dt�R�����ܙ�<<F�t�v��s�����%=�װ_p�@h�;���\��[9��u-�z	N����χ�Y����:���(�_S�L4W�=ϊ�ǆm`������];�;�G���c��Fc���u7��2'*��w)lK��n�ryq�0Qcks6�s��D�̑
Tm�koo+X.�ha�`�W2Ly�K8+�f[N�`�f:V'kr`��U��]��t�NUj64��s\;w)Ke� O`��t�/�W5it��t��n�sM8|itٔ����4背���ȏ=�g
Fb}����>V �G%e�u}�9T1܆��O��xj��?K�<N�Y,闚��Q�U���Z+�p��w����\�x�z���]6�����#���:w�:˨oP���,�Ӯ�'�C2ʓz�"��޹)>�,��_D��>�3p%�S��&0rKՖ2�h,E����!��bR��b�L�@�u2��[!���\�OI�shm�7*��8j*_��vt��{�X7�Q��xo�:ct���8�TuQ9ĝ4US&�%X�v��z�}'@P"r���nڪj���6ֱ�҅�;Ǔ�dcITqTKL{�a�v�lr\`��.��l����T|��x�抖o1��v����R����T�8-k/M�B(riحl��	�/_.Um�����rZUխ�hn���z�x..�b��uw��ҋ�o�\zdV�T�C���S65B�ϭ�\�����:���FQXh�P�P�5��Α�:xD��#�p{6R={�4^]����kbH&�tfb�kp�����x�!ӏ����S�wN��'C&#��i���-��k��9��`̔bc5�腋�������Z5�g@�Y����>E ����{�!���;�%]�����}�횗���]Q%�����ݜ*�tٷ�ܨ��*E��C-�V�R��TQb�!P�QA`��((-J�&Z頱W-�ա��E+*1�+"�VAƊ��I��#�*�B�ZE����:�8�ʨV"�A`���"��1̠��ۉ1����dU�kAAAAb��*�It�B�*b� �4�D"�5A&�k)�D��b���V����4�f�X*�����R"�c
�B�Eq-�X(��i`(,X4E�LAjT���V*� �Y@R"�,�*"(*�R*��0��4�F(J�Y4�
VV��\�0�Yt�*E�
)�R��.$���X�P��AAVL�\�X��1RE"�$Y��] `ŋ`(:�i1R!Y1�A`�����"1I,1�Rb(DE��w��wߝwu���ɸz�B� K+��k��9˪�}���]��V����*}���'T*eR����޷pHum~��G�n�sq������_Fs�+�Z�|Ut{�	��{^�����y{�!�N,q"�.��9�}�do�64��r����cc:G�kL��Θ>���wK��t�=К�v�]y���pG>�|j�м�Yf�Β��[Z
Ȫ�&"�X�u�'�[��B�|σ���q>[��U{1s=�������\�6!�ci抯�M��\D
�L�,w�g���>�Fnk�'�����`���v�OMOR��t;���>�d���d	����R����@�����z��t�G��Ez����,{n#��i�������#�Y<r�fL���c^[������k0{�}���\�/.#w���Q��׼o��q���S���NOuo�������Gk{�c��"G$��._g����⯺��?W���Ni>4܆z�cG�7i�u���i��́�7$�_�GeB^&~N{�@�Xs�c�!�>�~���-�sc���Lnl.S���>���:�<�*+�9 W�B{�niGeE�L.��7Ō��366$�뾮s�$]�J���q��x/g�?Nͩ��9����N͡�ı1�� �b%z�i��lr�W��^N&`[��_���ר0]p*�̏�kT��6��2u�2��v~�-�u|�sz���ᑗ4�9.�Yyt۲�|nf�f�϶�L�xr��6��s�f��uì���8��z����A�~�L���NDI��v����7���Su7f;b��>�J_���Z#�\y�W��ᢹد�uG��9��tȶw��
	>9M&=�f��ո�Y.��Z����>������&j5G2���H�)��:j�V��.n��	(�O����'�#'��#��ϧg��_,��M}���5���?m��;�3��_=jt�<ʉ��pV���2�Եy�{wڣ��}ޒO�ܸ�6���3�V|'
�#}7Ł�]��Y^�O��r%+B ��~�|�i�}{Q>�GLsz+��O�aՕLeFMib�ɝ�� k�#ه���O��Fo��jހ=���틝
�~����.��=�-���wIYU��ԸU����j�k�X����PY���l�����q�?ϩ�=\��1z
�P�6�p'95x]��ŝӛ�������'�]<;�7��g|j.e�x󹇢]{�N�=���J|�,���p��/b�VӍ9љ��O�����1��Yk���|w�0��$q�������N�Q=ԭ��uTn��&�+}R�C�i�52��=8;#���EUni����c3)��6U�FI�4�ރB�I'[[��m[�i�Tk;:� b����̮Z3)�y6�#T��Ajvs��9�`��M��Ɣ5�ҎE��_`̺�S�.}jkLp�Ҏ���&f�%���z��.@{2E�,rǑ�l��/z�<~��_��:�B�u�雇w�E�{D�q�W��Ҥ��y�RL����>
���<���/�v�X����zv΅�(���@w(�\j=p�ƌ�K���g	��]��>P�*SֵҞ�ܚw�S\5�H���`�������:�=儁�/�51=�A��)�m��}���\2�wlL;*7�&*9�S6_ �V �s����=2����$!2�{hM�FMﳈ��稆���Ta�-��To�(���f�7 N�t�Q�r�|=m��7s�.�G�
��'���㓒��mhw;�5�ƙ�{yfd>s'��⧏�1��>�^�ť�L���.���@�f���O���~������m���.p,5�t�TF.�N��UQG��9N�����2�3�?��t���B^ɣ	��]�"N3���C��+�X�͚�k�1��ӵS�-4(������*��i��~Z6��*�X)��n�g=iGYQkv��t��euTQ$*{��	� ɼ��U��Z�'�ɯ`6{�Sʲ��)U���h'�W\d7Lb3n!3]��nU؞j������y�X��gu����X�Е�,�Yi��{�#���p-�tm�*��f:��S�b��wZ��ݬKW�>�)U��oz@�n��կւ���C���3tK}(aR��Mz&�XT�3��4xk�!��F;�Λ��6g�o4��>gq��4מ;�]Eu�\�l�W�NRq�`�Ƚq��0}p��5�Q�s>���_�޹��w�;��W��>��7n���m�'��U��^nǊ��d�ɝ�yW>E�%v��w:Z:=���hw8�&\������'�\vϴ�K�P�<v�1τ�+���$^L�@��R�]l��y�%z ��Vۉ��ޗ*^�R�+�{���^��G<j%��%@{qR�^��T��աmׯ`�x�.}��߻���S�P�:�$_�P-����ȸ~�M��'�@<���NA&����/?^.�q���Ϸf;g��9��W���g =��Z+�uNH[����E͠�i�^[�Gxa� h�yQ�p��g0��3�k��
ٖGe�s�@y��'<|�_n7��Ѻ�\_-$(i�r�i1�m�O��Q�8�������/Ū��V�r�9��T%8n~�7�Q�Qm�M5/YR�ޙD���W�'�x@QIPa�ZrM���g�����y���1jN�����A�y�R�12����7�ܻ���|�B�w�74��H4�_[�?ת�m:���q�J�C�HGl5�myվ#���&�A�'JV,�;2e��W[ܦ��?�%N@����
o+�U��t�ÿZ�=e����8��}�ni{X��6�w7��/}D���Pw�#\����'�'�j���ꇵ�u�3p��\N(���v�ʎ�\�>T��U����Rȧ���Ci	
>}axT?	:n��|r��Q�n���t��ƻ'����O�<�V���zz| ���+վ#>�5�t�z�
�`�}���IFʓ�g�-`۸9�-n��qq;>_ZʇW/�5X���b���_M3�a��xם��c��IN�[6m�Z�Fw�Pxn)�J��T�fp�'=1��R��������~)�b�o�9��}����q>l�{��TQ����l�C��dU`��x�s�����ّ���3C��Y5T��{H�\��A���;���Uꌸo(���f�N2�*�	��D
��)�ہ��K�w��;b�{}��f�s�Tj�X.�1�U�Q�:unCR�g�w\MF@��\��\J�at�Z^.��	E׶��__����#�����P*!��~
v�/"�n\��ȶG��WC��Q)C�:{ʱ��Z�:f]]�]F��t�I��Z{�~�s�i�����5����w�v��-� ��m��z�::�����&-!f�y�YG4\�
�i�h��`Svq��,vWm��"'�A;��T�����k�����;]�`ԫ|��2�}<���KG۳��T>u�l����L���w��H�=A�����51[s��\ɶ.H�k���(��.���7q�̨��_r�l�s�O��t��󧎏�=���J`��bϟٷD(v�"G�K�F�e%�et�8.��rc+�h{��w�d»���Z\�/��<��q��:����L�+`���iGmZd��N#��,n�N��f����
��z�Ÿ�TO
��T͗�=����5P$��0�D��r��Q�Qk0�cޜf���Ĥk3��{��[>�j���+�K��5m �gz�k8]�:IElz��w�gBȑ웊;
�Ќ�j�Fqq{��;��2���.#y"ȯ������;����)��̎*5%�$�z3a��N-"��b��a��8�k�1�Z���yg��)�.�Y�#Q�W�ĸ]��G��s���IZWӒ���.��]>�Y��,�����{;�_@�s��Hzt�)�[�����[��u�������n"\�8����ɭ,_�3�7�@�pn���xH����9��w拷7�aV��N�U�Tk��Ԇ[fi#,4�h��v_������ݍ�_m�x�Gc)�}��R��]8�r��X���9o{eE�{*Tzpql`1X�.�K�S:zxu���%2V�\����T����<���Gm�_5���lzxs�7���1p�E6r'ӺJ��Y�R��SP�tǱ�)㷡%ɽ>�ɔ7��j���4��1�~;�M1���׆���ϟES7�p70�w
�f� �+w[��eGU��'��Ω�v�OǺW�[�n��,r���U>"s��VEq>��4__z�����ͦٴh	�\�\�9zd4T}��y�)����O����%��)A��o-�Nr�<�#�����G�P�*�ar�ȹc��K	Ej��λ�I�Ǧ�M,����Ѽ��R��Y7#
�N���rx�x���U!TL����>۽$��N-�7�o�w��M�3�Qsg�iW�.��ˍG������줼LJ�O7����>��e_f;~�����9�,W�ګ�w>{Հ/g� �s�P
�|uG� =;(_Nlg�����8y��Cn��v;*#9x_�G����K�'���{,
��z��ȵ�F�b*_�UKk�wP�83cF^I�\�J�/F������#��ٸ~t�ϥ�h��M'�sk�Fh�B��&ە�zh`c"ܐ;�.�4%�$���X�Hj>U{��wԃ�ʐ��2��gAy̫���	�L�Vf37
ar�r�fa��<(�[�F�h�	�����ˆ� �g�y�J��.Kjj0�(V�]v/>�\O���DNKq�Z����,i���ǫ�fCĝ������l{���wbs�;7��1�û3�|�/�,�=���=�=_�_�;���N��k���F� ǹW�[W��^�X�ߓ��Y�z����*
�o(ኇ�'p�R|r�qG]ZzxT^J��{�NKݥ��b�5�ncy�� �����'��.=��YY~1���c�=���>��u>��w��IW��jg!߯�ŸJ������v��c��M?O^yhpȏ-��ږz�K�.�������h3s�<2��;�2g}7��72�֞t������Ԣ��o:�kc!�3Y,������غȴ�*�	�uQs>銹��7�(ui���7<ϼ{���+�5�QJ�9�諢�x��[Q�yE�[��Qː�	X�˟"����U��1�� P��n�@^�lzx�h���^��#Yr�-q.�z] �}U#*e�Z���hp}%���׹z����R�`�/R_��lg��ǲ7�/�Ӹtn#ɅOt�;����B��`��~��:�u�JL:m����)	����:�{s�-3~��c�oh�[~���5s�u��{w�^�ֻJwwX�'���nu��9k��czgJ�:,��ngH��g��Y۲�.�U���[լ�ն�eb�ނCvm:�4rֳ���җ}���΍�N�w�>چ�{��I~�@��~��W�|�B侞���{:gh߻-^������t�҂>��«�2�q���͗kA��u���tD�ލ�<3�Hs�h��IJ��0|2�j��s�wl�:�{|�C�~I��}���L�~�g�'nm^fnz�ְm S�$x��s~�\6�����dgg p��tTm����"GP�^�8u�~��*�Y�~�H�ӓ�n)K�ۉ���V�w���k�s�νU�>�����3�НyQ:+��T�����҇;�7R~ ��5,e{T=���c��>�d�Cq��7�t�����ki %+��53>!{WI��D��'G��I�u�H��cbu�e�ɻ�վ��'��������Xk3����e�������V�q�������#�B2�Cc}훋�������f/	��}s����������ej�&#�V39�w[�����m%vM��7�o>���D�-�Ϳm�r}����c+앇�.g�gH�MDi��7��Of�^�wc���m<����hQ��_C�;.HWT)��k�<�����Xm�̽"�Vm� �챸�u/i�
rգ�F+)G�P��ɉ>}ҷ�D�u��:�:�	|[�-k�b��WCF��#����}��Һ�v�V�6��úV]j�'y�3��BM�w��Bm%8�-8�ｓ�n#��y��F���-�98
練	���/��n2gȵl{�[Es��}�%�'���_�i�Uj�r�ό,�
�\�e�EV5<������]=�;�W���ԏ��Y����X�z%���i����Q��+�o�2�|�V<���9젹 ��Vz}��}}=��#j5�뇁:l��������n�p��G����x�-ﶋK2�,{���)�X��22�z�7�����4j���:��r���Ϸ�:.�����n�n��䛋x{��ɠf�%��73�2& ��@aa����}�:���Os}}xL�3>)T~=�?.����.�÷�?u%ȁZĶh��쨊�L�9�Ҵ�-�%��<^L߱vi^�F&�9��s���D��n��5� _ʄ�{"n��O��jr�:��~^���Um��aޭ��
��r���3Q��Al���C5P��WR���ʇ�P�|�a��[�{��wIV�>��ғQ���_W��T%�s'�yH_ǒ���C�'�3�[�(s�[4�����'�\�Є���(]�8sx�����5�n���;��^ՙrG��S��Ěz�Q�AQT��v]�:b���=AC�VCH�E����S]��Z镓����v�А=�w��!�z�g1��9!���������9��03rekCG^�Vt�C �{Ә:��ġ��1��4\
2)�9r?j=���X�0�n�r����:'&�ב��\�P�P[�V4g[�{9Q���J�z��;�F0�RK��X���N�0��fRW	���8�hx)��9;�M�����-+��m��L�S\�m�C,�Z��<�ݾf-�w	eǘT`�cf[�V�hYN;'l��d^\������w�����
vs��(]���8L�qc���Laiѭj�����#�i�C�d�ڡ��T���Z͔��db�A;�4�yB��g%\���s��!���RB�Tw{�=�*oW�t�%�� f��eA*ɧW�[�V^Tb	Q�t�jG�]u���p�L�fsGfH�u����#n^n46UG3�
�̀�f��2=�^���to�0p��ˋ�U���4\��9f�=Wn��6ԕn�a����7ϫ%���E��z5����4�w
��7���ID�yQ�ݖ��ݛ��ŭ��up�1r���G���oMyg�j�Ţ*�[�^v%���o�<�2P(*F��酓9ܚ�����	oor9T�+�3�qֈsc��B�I�cD�<	|�o�]����p�i�.�]���ʻ�l3cer&���73�w�Q��5���n���I,uz:w0gH%g`O��e E�+z�Nde�<B�6�-�,�ȶ�c.�qC��k���qK��9Z�\q��ǭ+����b���1�7��&�˫�@^��AY:�VթH�gS��:-�T3����v�M��9hU�����tt���=�Jp����lŸ⨑���J�!>➽�Wp%f^[�e�f�j,�Ү���Φ�]sٿ
�d�]n�T��o6>C:e5>C��Mv�b�-�u��ˎ��=�v��	7�1E)0*L�q)�V lҕ[��pt�S*v���dbw�=��0+/��u�z��ϳfl��N�vV����v�A=ϻ/Pʋs#A.y����$[hE�[��yX��=E�-�vuN]�W!-�Zqpɸ/L\q��4pp�YB�xW�&�z2���;(���<'Zp*���AXA��N�f�y݆�$���c^����*�.�d��+Y�����6mCa��SÁ����Y�;{!���uD���eM&����S�ұ)��r�"�oL�4��_л�$�9Ryn���k-�WJ�֫�1���w�,jC	y��Kjh(d6���V�;Np�b�w��ݔ��M�
KGU�c��SBeɶ����VT�!2W�<�3T6:lF�"�U�w�Uj�,y-�R�����N��~m�v�_m+�l�yڹ*���K�5��`��:��Q���T��|fٖF)��K�xp��K����R�[5K����ᶤ��`�1T�*Kl�Y�}�b)%�%u�b �-(�*�dQDVMZ*1q���U"�UF"��F* 1nd�d���l��Q1P�Kj5���CD���+-%�f2T1��5l+������&5���#Fb��������`��md2��i1���QDdT�@QdQ@�C1�AV"�T���E�q0H��J�C��H�\@�LeH�Y"��pH�0��
Ȋ*VJ$Ē��1R,Y`�(,PRB�b�r�TT�V ��E"�R�X�b��* T*R�-���R,PZ!UbJ�I1�
�XT�$X�Z�� ��"#�Sغi�j1U��yn�vXr����[��N���bl~�mEڜ_Tt_�Ʈ�^�tJ���]���,YE�o������_����7�
oj�i����荨~4�����Q��Ƴm��������Ғ�p�x��}{]���qx�<r�f��Q9,]9��nvs�<���X���Nk|@�УvU���u������4˝.=��
��*p�>�vpJ_�p����r�<=*������M>}{3��6�����Kҳ=��V����h�S�v��!��|E������kO
��q�ͻD��Ǯ���^[���+vHYｷ��/���u��Z�]e�{��9��%dUG��V�� D�'ׅvx4����X�R8mo:xn1�~=�~����{m�BP���Y�9;�c0vs�@F���,;\��uϢ&����W��ɖ�}�*�^ӑ�◮�8/�Z�.:����[����@R�^�{����E;���r(��@˟'/L���/+����F����ܣ�^�V+�n���5�����mb�{"����9�/>�L
��#��aU�h{�&�>ٖn��1(��N4�y��3��j/��G�W���tKf��A��T�Q)�Y�=>f��Z$�*�YG%F�UP.]\���n�kN��^�ɽ�^ynP�jM�{��޼���|��j��b�*��w�^}t��0C�(Ip�p���ɮ�O������vQ�� �S8'n�f�;��QB�kq�Z�@�w�qթI�j6Ea�!��
���F��ݼ��E����j�í+����:�]�X�l���= y�{2
�lT(�>g�n�pFn��jѓ�d��[d{{}�4��_�e�'�_zwK=����`��`y�[��W&jD����B��\��br���8��bay�F�0�;��	����&*;ʯ�{��pg 
�����c��Vƛ֚�Lː����͆2�H�J�=��Q����PQռ�Ѯ|�~9;Z9���wW�iBZ{s|�{�9@W��^��>4���E�Ϣ�`�LJ��eF}���q�v��D�9}W��m�;1��)���`qF���'�a����;s��ڹ�.���Q�?���`�/�5Qrc�vd�g�n��րt��x\zq�
ƙ�{r��hُ?;�����:����q�}5�/<z|�mw�����w�Sb�[ To�S��h���)���`[��\�:�Uo�M���
�y��q,���ﳫ�� g��G��l����Uoޭ���1�P���J�����S�Ϳ1{~s��ӫM�ū�TuE�㚲�{�F��ʍ�O3��:Qxl�\�ѼN``�b�~yP9�_u�4`�]\��[����b ަ�fQi�����ڗ[8u5�Q[��HW'FT�o#�Z�ye��T2�q���+sU���v_@N��9P��a��ge�ٸ�&�>�V��ܹG��%�[�����ָ�O�]�Q�k�)�6+R�+Z�˙�LT\���#�w������Z�D�3e,���Q�7�\��q��,�t�,�t��X��"���<*�|^Df�F�-���=��N���q������<���rx�wh]F�� ;n!)�{�6��9�Uqnq���}��f�N�<�Z��p���t�|��~�d1�������x�+!g���^ܣ��nV�<����@~>��WַO
�M{����=x�
"�uH����r�n��c�غ�v��^���ig=/�$n��tУ�a����I\<�+���xc޽ 5�]w�'(�tP3��u/��k�^+�E�G��A���I�a��y��d���{�(|��(������c$!��7&�:�����j�Eu�$zd��͈�\2���k�a���1��k�B��ɹ��ʖ�qގ�[����ПM}zL��*9K���MK���mGeE�`�cd늳0�;7�(�8�Y݌��w��eǖ-j��_w�u��_>�1�q��B~}f��~;q:���X^���df�]DR쭞�ʹ�DL���-��y�w�9�����JR�S@�k���r��9�ã�r���F`�;��Om�����ǜt�fIC���H�±ۦ��uS�su\��O��t:��[ĕ�N_+.ċ����1Zx�"�vi<o�{�+��0�s�ʌL1�S�/������6��PД*���lgN��e�E=�
ww�����Q�:���_j�Qx��gf�pV[�/���G��:V�v�q��A��z:��>�Q|����={E��ti:X��+n*����M�O�m�&��Kщ�n��o/ם�o���;�Ȭ�������O�h+>�c0Ηd�1��\q��%G���4�+˥�	I����-��d���w�G�YF�����Kɰ}�Pu�s9�e��ՕFݷ��+��F�zdj�ë����7��f��z��A��c��roǦ�K@��t����U�f���7�\� z9O#y3��찠�:�p�K��m1��^.=8:�o�h��~͕!moD�U7��|s�V�l�J6��~ه����g�s��)�t��������`x�Wm�R�{�>=�
K��9��r�����@�KGۑ��}�i~��g�����@�ɑ3W��U�b0�?�k)
��]'��Gq9�2&�q�@,-9�/Ư����A8�/ʦ̑3/�-�B$�G��D�#`KS핂�C�*����WΏ3ߏ�hRW�a�j*ha73ι��<�ɤ2L�rM@'2�o�58l��t�*ѓ�]ݔ/��R�z�ĝeZ2���{UvJ���7h���j�kj2��h���ܵm������Y(�7�}�u��ˢ��'���
fQ9N{���~�a�\�����joH_�a���9ꦼ\>�!��s��M��K�����ɒ�!=�4���-2a�q:�i��d���)o5G�������VK�mS6_ �O���@���x�R~;���@����]N�Y�w`q�����l����Q�����o�"�?H�2/�~S�{���'�����q=��� ͚v���f�a��1GU�ztv�71���I���dS��t���z�Q=�1�������E�SG�'ƶ>i�'
�sc�ZZk�5����e��ci�D-J8^��N��Un��>��ܧNz�/>��D>�N�q>S������aa���/ޮ�q}6��r��t�hqW�D;N��8���}��Q4�(銇��>"�.�c0Ζ� }�NUyk�Kwq{��>�9U�H{Gm�K�_���yHu�e���E�x�6s��{$�2"����&��ֶ��и���Z+��5�����#�g4쿱�~:����u����rG������zr�em��M�|l�-��3�����f��;U���٣2fa����ݷ5Sg��st�go�"Fmf6^5�s�= i�-�:F���;
�Z�gVBe��nE.��5�!#m������Ě�fC[jʨ��^��&c#�E���y�j��!I�ړ��rf(}]�q�S7�,/�TR�w�9+���/Æ'W���@��3��v�{Y�������.��s�l	��}~��ϣf�F��P㜤fe]��"����aR���|3YG(�������,��@l���ET�.Xs����'��gs9��5����lAX����~w��C�.O��ѳ�eBR<�g���ܗ�h���W�oi˭̹�^������իGTrZυ���Ӿ k_g� �r�B��n��SD���Sr���w�N��V��%{grc����l���؁��:����P���J�!jǛ+ۼ6��p�˵b5���p&:��0�����3e����`={��>Z��k�.8v����>�z��g��f�9SY'ah�^�i��!1�yѢ�r��>/޳rq�Z{G�vD�w�o�� ��\���Lo���W�W�8̨��%X|?^�DcʮU���x���^�~��̟L7�
t�6�c�4�I��I��z�������ZA��h��e�s��zob�Mk�1]��m�&����+/���:�*ָk�BW.!3:�:����3a��"��#A��oIT�agB��-U��Ob��8�8J�iՍp��7g+�a��H��A|��H�'(ɻ��u�킴��Z�X��Iph�F�~�f-�6!�:��x��縨*����+� ���񼏧u���)���%�%�O�cѽ5�|@��ux	YV�����p�wLH��
����.3��uŮW}�}N�eZ����5� gTj��nr=|��O�kF��[X���C1��o����p��{��S��*�iS�E�W��'�Yp=ƶg�W�Ξg���|����(�`��GhW�㸻���}�ϵѢ�V
Ȫ�&���e9��k��oJ��Ɩ��c�X
v\�i����O�H���j�o���ȏuLۧ@>Ϫ�	��EEϑ`E�h��z���uU�еj���)��h෣�t�>�����P��҇����9��"�Frˏi�
ruxߪ�(�ec�w=�gՑ�«�h��;c<��=�o�\��1~�f���{�%`���f�g�3�K����U!��u�8KGٟmCV�"ßJG��(y�E[�r5纉2(���t�ѓ3��}d�M�{7��}.�D�9�&9���Q=�ٸ.փ�1�:����%�
>�܆ˬ�iLU��Ɏ+Z���6k�����48U��;Ԙ��xxlW��2 ���#"��0��,�6�8�Iݤi+RG���|;T쮤�Zk��V3���ȡ�Øb�N)��Ww�Q�l���)��I]��N�Յ�L�+��?����D:it�]�3 �b�w��wX/�t���b^j)���Wv�����F������*M?HM� ��9"�"9Ϣn�����ZdV������ľw�����n�N�{�ݗ[AGTk\jb��A��s�=t���Ĭ97>G�蜨{y[����%�vMH��.D���r}�Kj6�uʬ�M��F}�t�~�VՐD�y+��#��M����C��vk^��1�x���s��O =��ٙd7���Ci		�������'GG��88�N�,�N(vj�TuE�Xj0�;7��`
�V��~#��W�H��s�Jr�Ź�Bo�Ю����A�~7۵��w'Nܺ:X���]��gC=:=/]G(�I*��9�]��\������<�7��+����g��{Dw�tESQ�Z]�L�/\��\]\#N�5f��s�}���_�iqg���#ڶ�56����ӳ���.{ŋ�xW:p����+��>|��D�+I�2�����8�{K�Uꌸo(������r��Ӿ[F��h�ɏu� a��n+S��-�����g�;���/Gm�IA.�/gjF�.*�:�V���a�&>��e�ž^���n��F�S)���ئ;{c�Y��WB���[��L�7�/lHf�7-ަ�l��V�o��Z����[$��2�o�\�I5����9\@�����ɖ���c��`��#^Eo�xuʯ�;��>Z�cT�U#3n������X���̰ܨ���|�+��.���	�G	�]��E�N���l�[;����㋬S��\a/�b��9�[�����CF�/��ۯZ�+�ز��1B*iJ�y���(�.�W�߯FDzg�]��"g6�D�r���x{��qcթi�q�>�^�V�I���Z�y�.sI�nF���_<�t@�^�l�A�Ҳ&����z�9��>s���{;+�w�_Q����w��ϓ��/�9������*�U2@��G�n��O�uw}+�X�T�y��)��&w���F9zv��X��TO
���S!�l��8�*���<mk�'����{מ��Zy�ڏe}k0��N��/U�ᢣ��cy�� {��ůR���{vx�o]Wb��,�L������ט��%��=����uRc>�H�;<�Z\zm;�Md
���C�M��`�"L�{�<nW���1b��X��+z�3�j#O�ޠ%6}�H�V�]�7Qn�Ӝ���lE>1vq�LE��;�\z�*�ߪ�����0�u����:��;�M��ԧ:ɠ�ʶ��v��̩+Q�N�&�m�(��jv}b��օ�X�^ܙ�C�d1�U-������Q�a�w��Ãp.Q�{�Vˏ8�J�ſWR�<����7$��s�4�{U�_�>���^b �jf�Mv�绌/K��2ۨ�]nt�׼j��	�5��o�r,��oz3���{Y�U�*sE�~��Ǧsƣ����!�}�\ ^�'�㵣k������\�[�ٕ�=��~3����5���&NL���b�b�g|n2g�<����i���Kg.�cj<��0n\S��5C��Ǳ5�� �H�>�s��ɨ�&+�p��QnX^<�a�s�/O3��`>ٺ���d���#Um1q�h���k���dP����'/6h4o��p�=�f��6 ��U�W���	�wO����w�ӴQ�}�@l���UHʞ\���cN�����n[��.�v5ǚ��Cn��?Nq��#5�9k���qD�l����*�.�<�a�����TE�w�\�}Ǒy��ѳ�>��ữ3�!�..l���rPD��<��.�ʡ6�;FM{H��{�)�&'zV;�dZs
��R��ށn��D}��!	'�@!I?����!I?BO� �!$��$��!	'��B��!	'� B�~�BO��$��BI�BI��!I?BOԁBI�!I?BO�BI��������)���7� �,/�),����������0TO�UAD�)@��((Q��Ғ��D���H���)D�Q!R���$��)w���m���JCaT�Qe[m�5U
��f4��  � ��,k2lͦU"��9Ӑ��-��Ѭ���-,m6��ER\'�UD��r���i˔N�Zwd�s����K�)��w[��[m۹��;L��ųvҫ;������(��R�e5��j�$`�&�fѠ� 78���e�[Ḓ�%����6ʕ@� ۔�(�Kf�ciY�U5Yd�J���Y�mm���l͓*�k[6�f �
��n֭��f��5j��,�[lw��H@ 56�ʔ��M 4i��d��$�R��      �&d`bba0�!�&�O��T�       �D�LF�LBcQz��4�5R	4�BU( �ML�  �i6j�f�{e��Sm"�nҀ���	C��������*�@D	��!PAbĲ�?я���~���â�h����.�!!�bB1Y
��Һ�(X��~|��p ���̔�&Za����<{daP�l�Q�@uo����0��x�+-�R�-*�p�S����^|r�e�6�R�����V�C89e �w��fdJ�h2�}�,
EJ;fS�����#,1�5��W1L���+�ܻ"�c�^by�7v���!vB��`�7Pb�.`*�;dC(Py�+�1�Th�Mn&�[[�H���ʳ�u�f��9+��fZ�'r5��t� *l����^��HՊ�b��Z�l��&�,{D7�P����=4U�X��a�ұf�1M�tH��� %7��sTq��ʴ�3%f5�����c�x3a�R	�6���)nL:����3.n�KU���+s1hk^SGR������"�*t���t��f@�������ۉ�[�h��eː�Q� �ޝ這8������@��*�eb9�ndI�̥��R�.V���m����-�; .���Ե��Yy�u	v��rF.,Ӡ�S�AJ^��.��:�8�D����s`�D�hm[ǵ�B�H%mԦp7YcnJ�;�Wjf�gw��e�(�PS4�� �������ya^����ȐK�v3KB���W�LAtve��!vF8�#*5�{�nK�`�'*�����d5z̖�=���mGX1;H�!a��X�^����+�dN\ܥi*��HQ��b�@��ܩRPJ�Y����cf"]]�f�9r�h!����R��VP�0���w�!f�i#Fn�GB�i��)���@�f�b�ڽ:��m]kp��ۢ�1"v�XYp,{r1Co ��S2^�Bۻq��Kf�M�W��o)e9t�3fU�S[�h)�V�-|�2E�D��*R�h���B`B�u�d�t�B�n���J���%-UX��y��^%���EVm�T�d�J��K51G�K^�j�k3:�3K��(6���ɲ騐��Ja��1)Z)�neՁZ���b�`iS̷xQe�c	*�r ����V�B� ��Y���wDd
&Y��I[�:��-]<
��hk5�k��B�-��,�r�S����5��V��$`�w�lx2�E�˂��k6���.�ݖ��xs�	͒��^�ז③�ި�{,�e���n�m:������VK�����!��Z>J�-m��Su`��de
��K*c�J�MJl���)C�����tM�6�B�BX#	���6�fl���[	&�՜�l��CA�����b�bb 3��.�bTc,�;M]�R�ǹ�u��d�7ZB�<ʒ�L�y[�y��3`h��e�TD �ݼ�/^��ё����r`B� v����ԭ�ظ*�̏�le9�����JM�B��T)^��LY�@�R�71X�>ƀNY��5e�'*��7j�Z��Z��^X���[��˷2���f�������8K��ϵ��Ť�-[�����ط[W�z+c�dSL2�kf�	�n����P�0޸\L0+�h����Րo�b�=08�E�t�:N�<Wl r�)�X���ё��r*ܥYBY�iö����=�O`!V9zwkKЁܬ�VƵkٲ�t^���ƫ�/ZJ�k nõ��Dhڨ�z]d�Z�@X��v���IOD�Yy����ɳhil�{W�`��;�"L�E|-&�(#��m��F�Y��6����.�x� ����V�EC���,QKy
-5.�X��-�ٱF�cڔ�Ć��FpVH�׌�&X���'���e��F�z����i[���,���SvRwt���i�(�	Ifj�L�3U�qU��&�t���8�0���$�*�hI`�y�q
͚Em�)*V1�	��1��U�V`b��5�.��MLĪ,�2͛�U%Ԣ(5tРs�c��m�.�x䇁�R��N�J�&����C��B�H�ܫXp �'+��5��ъ��Z��	�z���j�#$+U��k����M���:�H���JF����1'�n�2S�!�Ï;��յ�4`���3��'Ӻ^�ֵ:����U��[�o&ɶ�R5�K��ʗ0��
���mub�<7��W��|%m/�dA�sd�2 yZ˫�{�u�n�ԟb'ju��g��㗮��/x]N�J�(�Sa謝
p�:�+v;�W��%h����D|�p:�_w�Y�]�W�NY���S*a�ϟ$B]y�r�ӻ��N̺�Y!j��OهgK�y�.��z��f,F������x����Y�+4�Gݯ��w٩�!ø��Σ��;�L���0h�
�6��3�/9!-�1�r���s+���U�Ѝ�CME�f�>$F��iX {F����J,ɓv��$�M�&�^صE4s�t���o#��t���Q�I-v.h���k��V����5xj��+��ֳ�J��6� N��#�:��鎐�_���J�k�q�g��f�A�"{��_Cт����=�,�IU���
����D�]��݊l2���'�cߤ����+�;i�(é���͝���\Oe:�iʔ26�gn�w�ń5+#V(�����c*��F�:�Vu\�q�N�;��G���4�.�t�M":���P� �{\���[�4*1{4�r؃����*�TZ��-vc���r�Z���-�r3Ao
W�ʊWvL�}z��U�+.��8�S��[�X�X��C2g#�j4���xoG^�#���P�xEgt�OkF%Xw���ں��Y�'n��#�p�K:\5v�)��'���vo8�߱[�S̻�ݾ�;-C�ӊS�֨+���_G�m����#���B�6x9ܖvt-��t,���o�`m�o��0��C{:�w	�&�j�k��2��p�J�����v����u�3���U:Ԍͧ]ņ;KFԄR����#v��)'�I�n f뫂^���g'+V���n�L��F���Ύ���v� �m�g��Վ�?&��*���6ы7;;�gej�tu+.��߹��	�k�.W6[un�`^nҸԽ�\g��ӯ�n�b��-vг:�b�U8a�5���)My���1�
il��<�P>C�/r�5�<�Y������7�eS���j2Ҽ�֪ȶ�sH �Z%*��s&�G�a��
U��8�PB���T�G��(��Ϲ1�]�`��U1���`Ert�yY.����TS&�9�.m�Й��\f�e$�;�z�<p���y)K�u{�Bq��^�q0�i6�X�M�K�yӇv��ԥ=�@m���x#}��˥eҏ���;�i{j�	Z9���:Nޡ�.�$d�Y���d�Q�C$�=�"��̍��go�_+{O�G�e�gw�캼t��9�0F���.��#�1e]NY�rY.tLgfm����p&�(����B1���8#��
��}�%K/�7(�R�s�u�Ό�v��A��Ջ��ԓU
W$��;�C��3&Xu������d��b�\޺ceW ��<�Zn�z�f�q�\y�W��j��\�_#�󕠶#�e��= r�����\�+{�h傮�(���ya�[�T��{&��ZH�i���f멮΅xҝ�@����8}��oE���>`7�]��SW��W]Z�no6Ș��.�V㌦b��S2g=�^>j�S]9&�|��pI�48fXc;CeqRoݻ]�Z�خ����3�'�<v]͌��9h�	%��8�ZZ`�7o^'re2����w����H�5�	������yX�`m���V����vG5�������Csu oz�����O���ݥ:��+]M�"�9�s��˗rbK���u�$�����Ix "S��l��a<���[�k��7�,=u�j�K��W!����_e���Rp�&�whn��x����ԥ���ʋ.O��0C����ꓮ	��^ޝ��e�EL|쉘3���l1�JR�U�Zk��^t�٨�i~�2���E}� �Z	�;� ��n� nK���P@�v��l��4?�C�/��#�r�qkX�Z7p�/#Ϳ��ԝJ�|)}Ո���K]�"�׍�p����7�i���{�{kn��+r���f��l�"�ժ�h���+�SC�R��: ���Q-�o9/V��7Ws�u��y�P�>@;ɳ�9���U2����~�v��u�%��<[ �E�����X��(�H�Q��M{nJ]��'�w�{���0(�ɤ^Z�[����y�ls4�|�1e�V�x�ۓ��HP��m��Æ�X�6������	�_^�`o�Z*+��1K��ɻ�5����.:n� �1v�@�r��~�9��:>�n7w5�j�̳�a�2��o.���l�7�	��N�
��ʒ�Ȩ�#�ڻ!t!x/"��vR��s�h�Q��5X��+z��Nu{�m�[�|2p��i������7M�[1(]�\�Uj��2gI�Yt]h�Mm#9�ŭe��R�>(�[�^����Zq��J5u�U�i�s��yUq���n�z�λS��a䴢�6K�n+�ݫ�q�`�|����q�U�c7/r����5�D��u��s6�cWo��n�(n�t�x}Փ��R���fꘙ.J]��fs跄xkyv�;i��y�b�^��u�ڑ��}y���e �9�w4�gX�3Hќ:���W�4�_nFS\ﮛ��a�S�u�����nŝJ�&�e�[� ѧA��e���o{���	۠���p
h��c辱}��Z����'��S�Ĩ�	�W�.qVA0�J��r��l}�R���p��(�S��kx���l��b��,��:�\��Gi��g�Y9��u����3��p�bQ���7]��AT�q���KY��>�ʃ2'�|���W�������9'�gRܤE�i��UҴ�5N 2��<w���
���.�t���tMC�m	�4�C�Bt�u[�h��=���f���Ű��b�y�f��#ɭKp�@�67�e�M`G�$S�T�R�!�2d��&���"��jD.\Nݠ�y2��i���y�c��n�����wU��I����0��Ys[	�}v�r��^%�]=!\��VZ�X��F�φ �Ӭ�5ɴ ��7mr�WH�|*�S1��>]\m�/���=rY�s+H��B���\� 8E��+��ܶh�`c��>����%n9[��Q�(P��-8V�d�1e�M���߂�v�I���!\s"V�ioc������J�a�	xsK]���l�V����VN�ƖwL�^�CD�4tr�� n��L8u�8��w"�C�Ұ�L��@�K8���=[K7%��%B���3��v]�41����U��h׷uc��}_X�{��4�ޘ"����+Mwn�T����ݶ���M ��Z	��,_0���GL�P�&�=}�0������oJ�7Qj�2�!��bRV�F�sN��St�,n�5a��f"�u�l��"�#������{u�4pm^2fc�L�ǽs��g�L�bL�F��v�2Ш]��6�%Pu�p	�k`C��&PW�: ��Vn�AX��Ѵ��7im`�Y�/.Zo�� �t7����y|kL�m��uog�Ɏ�������n���p��쮶s�K���I�N�6pH��\٦bm�k( ��3����]mM6�RN�n_Ӳ�3��]���{E���e��r��a���Q���ؾL���yQb��kL���!Sa�,��#�U���p���Y��sn�����1�F+�R_ZW��f�K��v�C����c�T��V�^^Lb�a+v���2�t�����#�Vpk�N�8�M[kn�V�[l71>��bΧ2�{5i9�Px1(�dB�c�Ɨt����v@���U����1$�!e���sE���o�}F���I���Z��x,<>ˌ�k�s78NBX���HKƸu�������� �`���� ���}ڌ
o�7�?o���%}�U[��yt�P"L�9����s[r��=���fP(��'��t�Di+���;��1��f��*#ys'�H�W��$�u��%K��6�Z�Ƅ���c\��^Ι7)��$���0��|e��$��lfSŒ���aŪ��W{($.�)��;��Ւv3[��fڗ:VRᲜvBbV��ݧw����.��c����.C��^����٭í�櫁�9޽����},���FEzQ��ֈ�&�S.�nP�t��6d޵�Z��f�Q̸۬���fT\�m.!ij�jZ�+Z���l�Z%]��5�d����̥�kkZT���:�9�b�Q��i-u�R�ܷbeR� f�� �uVW��/'{z�y��h�.�;��;w7z,�\v��?�\ڠ $���^~���4ȶ�- �,���ǵ=Ѥ�����}���?dٮ�t)M��T-Ｘד\k�h؃�ʤ|fZ��OwW�}�b������F��B#��_��n$ٿ�]z��[L��.L�i��A�ǆp7 /�u|:���t�w��q�����m�����E��V.!*�q�G���5MA�[7��ޚ]u8Y��`R�;�;W��h�m�:ܥ��E�}�8䔴爔;�,�o�n��2���2o9��N;F��N�2�z|�=Su����Gdd�gq�2�"�Y���ϸ�<7K\o��gWW�V�J���(��cw��]���|�K˵�ި	�W�1��7�,��W?j�˞�*��uɎ��L�|����;���<(��sO��uc܆�+]�u�=�|���ܦ��� *Py���[|�3ǲ#Fn'7�]t�=�˲��CO)����L�Hs�*:�����wܮ(�kj��Xx�P�J��^�aط'Vj2�r�̫��uX�G-����y(zt|_3�U%�J����F�V��Hhݨͣ��/[au�jn/�W�*N�z�E�'FU�x��v�[]=U��۱(�������^E�O^���7�E)[�s�����::���o&��$�Q��u��f:�^'�#����h9s��.ꩣ3��vR�j��P��ꋩ������ҹ�
�z���5��P��u�����Hm6z���ީ��n:<cŔL���<��^��is��o��\�4�V\U�֋n�5暮F��H�rc���>5y~�_h�tF�Q�:?M�.ï����z|�n3Kj��D��o_g�����e�G�b<��Bۢ�܃�Y��-M�q�.���u��L�vw5�����v��d�QF:��ُ���`��v��vk��b��.t���n�f[�;�޴)��mu_�r!�����j�����)�CI
(��+�XG6����x�� mы6I��5'f���両�Q�Ф�Zx�Tu����L��NF�Zv~��{e!�̭�|)WTltzP��e��\�U���Oj��!]��uf��I;�Wng�z�.�ھA�<�/T�V��-e\L�u����i�[��&�x���w+���w
'\���Ck�"�B�>��.OE2��~'�ٺ�]����\���ۅ���h��g"�*��j�י+�O���Y��zj�j�>�5��[�5���ý۹�-��MSvwf����Y��;�>F3���k���^(�w&����i��oMY�k}�i��cUnCJ��{m��#���T��3ꋣN"L2�����Gm���ow@󜋤�zua�ny(hL�K'OV䔹��T���a2�gh����0���q�3�}�͏_e�t�^�ߣt��Sj����J��'�bu7����6�f+�j�	��8��[�]�΃����:����Bg�N�cEi)
���ݹgS~�[B�@%Hoc��A��.O@�
�P��'ߑ�������_�)c�:s(vY��ӓ�l�g�n%F������2�f(��o�{�έ̷/��Ӻ��N�7n�pfC)��t4�=�-X���?�k��I�c�o����m�v�r;�gpg<�pK�f��0�v��z�%{G�l���S�qU4�WeC/"�ob맯��U&և)s� �\�L�r-ѽ㔸;j���u�]dn�8�N�y�7��l�
��k�R*	�ps���_�>�������f;�;t7�'�
������j<0S�YY��5 �,P����6�2�3���6�!r�7S�ܥM�{h��*�%iV��;t�5V��TIZ���Y�Nٰ/2�i�o,�JW����Idiی�Z�eAb?�Hc�2�?��13.��BQ�j,����yQ}#�t��)�830"�Q1R�]�`�h#���J�faZ�!�m.�e�ʕƦ���R��EVZ�1�ն�0��s2���ihԵE+V�+��2�T[uq���b�(�-�3QF�PKKJڦ�q+SYU]k4�L�����:�KQr�V��j"R�Z�Ѭ6��0�b���_�b`�V�j*+8-��֒gR�������;���D�ʻʏzl���%���F_�'�*а1V���w����YU�ϫD|�ڶ�r����:�rC��۫�h�DL���J�t�B�U��|���ֳ��v���3z��w�v��`�#���y�P�,�M�x/]g�EC��w02��ʅ�^*���J4�٨�>u"���pv�'[U}7u�f�/�;C6�1����M)�/O�kj��!VK�g D.���[v�:oE�X�xZӻI����OC|=SRE���]d�pN�\���4��nҞ����Ko���c=���Nͩ���NѲkxr��l�kCs|�]֡lע�Z����:ivj n#���o������kޤ�KW93J��B���z9̻2��ϵ���wzoQ�ua]L��Oq�"��1S¨U�� �������P����:���x�F�p��"�Q��<�
 ̞�G:�vTp�����e�ƨ5ה�>�1�  .�I�Hz�\���~;�~Ha8��	�m��L�i!�&��d�=�a
����ܓ��O��&���!��$)�d'�C���������E�B0<@=O�LՒ�q �H}����v@��06ȲVIĒ_,:�? g�d�$�@��|oڷ�$�����mz>�i$��&� � �s�Y'C��=Ha� ���iu!��2����oxH
I=a<`w��!�@��P��qx��I>d����7��b@>`cLOև́�Cl��2x��S��Jk����� m�1 pd��B����R9b��!�@�����;��A��D�kk�v`ܻ��E�K�]L�Y�����ֶ�/?i$7� 
C� 4��$���Hi��É��9���d?204��d�����m	+$�J���M3���l8�;��B|�?!�H�=HY �CI? ����t���y���>gY>a9�!���4�HNy_������C�M2J��XI�m��<��@�$��$:�T�ׇ̐���ށ=a����I�!���﹒I������:��~��5�C�@�@1��2(C���6��$�M�d�Ԑ�=�^���!����$�I6Ȥ��I'�I̆ćK�k�}���{$.�!����3�q$�a z�O�<`2m ��	߹��� ��<@��}I
r�>� �� {���n~|�������9��ڊ�$���d <G�.ё�S}��7���_���9�Ѫ��(��E��'����1��(.�c������FRB�c�%!�8]p��N��Ͱ��-�A��ֳ�+�4罺�&�:Od�4��u7�+�LJ�l��	�s(My[�b������v��a��żʿ�2���1�����s%p�w�-���%g?z�*���h���"�߳uö�̺�E�r]i�s�J�X�(������%��^ӔSkС����<p\�ǰ�0 C��rĦxd�Z9�T���B�IKR-�t�Gk�}�8@�Zu��yt���Cf�Y�5j��:��\,.��+��Z���M���qF?ʽ1N�؆�Ws�Sn���*6�1WÔ�n�Eô��Z�|,��Ϯ�~`�x���{�-I���Ln�V_�4x>4t�ds�,P犴zH�ۻ�������\ξ4���|0>5t�~���j{��-�V����y�Wl�oxs�;6N�&����_�+�t�o��g;���?]���v)���҇�S״s���*�9l	��j�K/W��[�Q$�X�]c�g&4�E��D������t�e�뢼��y쨲D�	����O���u��A\�:�ۙ�運x��j5����,?�]��ǫw�:Vgg\Wu�KV���.{rf#�B5�5y��Q[6Z�JdP�^��:�W}��W������Jߣ�i1zJ���R��g6�R����@{}3�|�����
5{ֻ�_��}~n���K����A��.�ohwXů6��1Τjx�����t����H���ou����l} +{x%G�H�V�Y�p�c �&7v�
$�<�1A�S�M#\�&��k�`wx���ׅ����{�/,D7��O�����C0�����=Lv�F�Vt�~ͳB�sQ�v���2Ŗ��[*��l2Sհ�(�q�T���Z=uaaH�/��q��7��v�B.�,]�+����N�~���O*�3��T�b�DDfF4��Qd�T�&h�*�VK4�e�B�Ŗ٥D� *?�
�	d�0�zʱL$`F���$�mS���G0d?A��MX5	QK��X�`"��G���9��Pw���
�,��й�j[�R��P"���;���[��dMi!�y�-U�g1S��
�8��o���o��=����w���X�.\(�Lq��գ�\<˕eDcYR����m�m�-�Z�hU�+aDP�1���V��J��c����J�����B�V�T�mn����VZ��,*fc�W2�YX(��[RȢ6ذDZ�YU��1E �A!�������M.���+U,�����W� ��зBm�<#� ��������^��� ��U�Y��mkV��r��Ѽ�r�ʣ�+�����>�}�i]��ʻ�Y�*�'(��L�.�
G�,4�v�t�ٝ}z��� ����/{8G�i/<�<�G���y99�*T����z�R�t����3�;���,�� ��S��\�s�5�e	߯v����J͚V��2�P��\�ycm��9*�h���u��|8�+ie����M�� ���>��AW[y�yA�Z�<�_)���R���U��#�xJ���總�i��7��T$�hbp�d"�7;+�-`�r"d"�i=&��I�k�w�<�J֣�S�tc"g��=����U��d�:{ח���?%[��v��xX�F��K���=�y��m����Vr�D�h�p���2$�۱w{B��\����֊S �n	��d�]���\N��t�qdO����⊬���>�|n��[���o�=�z�3��I�'ﾯ���ђ�R�����Ak�W�U�U�]Ha�S���G�Z���RN��k�T�:����^�FUF�>T+�׃�	�NT��s����ã%�jO�K���\�k6����J>�9�f#b`D�R�-��e�Vu*��2�[��RG�2��K��箔:2�w�-�R����[�ٹ}I$���{��
Z�_d�u��2����P��g����>U�KE��29v���	�ٗ�7��[o��鼗AR�{ǚ@���ovr�����.kSsݕ�Q)C��;����h%�Q��@�o��7�-Z{��߶�	��$�{ �_�h�0ǩ��	��t���,�j�ڶ��C�)_�zŋ��SG�#a�Z��nNew�Z�ixl)e�Y����o��P��v�?h۩fs����t��Xlv=Q/zD%ٰ�4�G
\�e�C�&�v��{F4d5�B�c�Sי5(��ڥ���ɫ�ٸw9���"u�9�f敏�cz�9k���k��U�N`ڝU͵���]�f|���(t��ܹ��\}P+��QO�O�9�Z �����V�7.�z���_���/�v����t�ddu���yʪ�P��Wc��Bn������xgb�¾�l�;+��{`8w{ٱoG�<c���#�n�)�.����'ǝ�X�o/�,0�Y��V������s�L�|����Ti�,]�"]�w������< �>�� 
�H{h�����[�3Ya�����)uӚ���כczJ=mK|�؊[��G9�V4�n�҇%,��{^Frz�o_�;۱�ә:�P�;�wރ�Ed͊Q�/��0U$�=�3B8��{M�xh�ʅ�Y˞�V�L!�����
�]�{O��Q��VP���#&k^��E}&�9���Yix�oo�J�6���g���#��
�}.�v�L�|���o��Z��R�s38?5���N�np����D+�ܔ�M�z�TձW��{1�'\([��->�K��:w�0�/�V6:�r\a+i����mm���7=�bP�Y��V���Ԓ'��L�|ߑ^9�kiߍ���D���t�Q�:�vz����3�^�~#�������IFp����e�M�M�sE	�m��yM�y��7��mQ}�*��Z�½��˅��v4v���/J�2��	Z���o��N�7�̢X��BGPM�/ �jHZ{���nҝY��8��V�v`�a�Q�7M�;~�I1ŃWo	��.����v���}���q�2����)�h�X����E��\J��{F1�r5M�ew�Ԯ��R�V����G{o����>=6�K����3Z�`��9��:铍9cn�i�m�lt{q�%�1nΪԞ����^���Eh�_ً�l���^7EVi��L��&ݭF�V#��Ul�ڒ�BBے�xm�#�g0:l�wjf3&^92x� ҧ`$K�,��a�Ӷt,�l�6�ޒ�U�n��Z�+�ʻ8����h*�1�����:��vZ�WFL���&�2�;;�����(�T�$QV"6��V�*��E�
����PF#-�TT���L���کjV%ZQ"��*��������FQQ���+ZZ"Eb1s.��6��4��Fʪ�E)2�1o+�����4�}:��q[+�<<��{�p~j�w��^c���m�Q��N��u@����q��)�I˛3��s�}#R���42���}*�1LP�T�u�.9�<��x'���s�^�ͧ{q�����,=����L՞c�s�j��EHR�p�<*��A��������	�>0|�@p�/O�w۰�g���H�^��]�p�h��;�]غ����Ae.{��_���a�U�K��o_���g磌���v��A_���7f�~g���]�>���˷i�ǽ��a�����߼=b����z���z�|�l�t�{�M'>�8�*�W�h���@��K�����*
���x��秛����o|��l���6��j��-�4�}������� ���l4�
�HJ��K��� `Zk��b�8S:
��� ��DX�j�8P�}��$�Ǣhg���^r�9��[�;���,�b��a��}_W����V�C���|M���<N`��w��9����4l��1��wnn}0�V��Z���=��w~>j������:�q���k�7>�>&��Ӝ��=����}��v|�߶i�Vyn�	�}�Q�Jx�9�����*���Ѿ5~>Cm��*7h
L��H}���7����0��5�>x�D���W�0*�FÎ����ΟT\||@ĸ��nĐ�p���՗,����F��L�|'eWuL�Բ��j��~����7����rf��ϩ�<^X�����n���'P�Y��ut���=N_u����J���M���T.�;�g'��Z�1DFߓ
���g���Y�+,�#U }HQ�LhH��+΅�r�Z����kEV
`�=Ons8mO�|v�f��=N��<g(�틞�uYB��xpB��^�5�������r��<*�����OM@�*þ5��A��c�
�0|Es[���0�ǥ�+a��wK.���#\��˴�����N�WW[Ǧ�.��{�3��E~��y}b��S�}�����^_�V)�O;f�Vy�:�;���;}�:���FK������
:D���
��I�m�S���|���^��b���L�����F(�v�0!��U!_��/�=}���������t�?3߱�r���}��f����d+�8=�Eɸ�"cɐDd��hܗ��U�+�F�`�5��Vi��U;3�<�M8�ƍ�$�ތ���\�:E�]�;�/p�GF�%��#�B�1;8��i�a9�G)�ﾯ���}���~�����o��|��r������:��g�m���7c��/��9���OR�Lz�~N;g��ȡ�I��b���@�k4.+Z�>��-��Ui��١����|�>3������(���Vf霳g���Η�q<�&yOS~������륜M<b���<�O���������
�����򗯻�y�c�zΎ�k���!Y���1n�����<�9��O�<<Ϳ0�>yʈ��_z��~1Yg<j�Tbi� ����O9��+U�������\>� {��nf*Ⴈ�c�
t>���,X���&{eA^���c�1?V'n����*���i����m�;���ok�էO,7�<k.�I��9� �Ռ�\j+�e)�P�u�q����0�F��*�����ٮDD!����W��eY�<R�:��x�ї�(���|p����Z�]]���6J##o�E������G�U<vΧ1I�S���}y��s�0�s������b�e�?Q�e1�+|mi�HK(W�n+���X����w*c>�6�o��Ϭ�x�g��.�S�~_��9ϵ�ޤ���{��wVu.���:�c�Tm+�8|�Wh�ۯ��\ p���Ǉ�*
g-�G,�o�{CJ���=���̼��;�uם��2�Կ���7���*8)D�yku�C#}$v�>�3[�;�<����,kYkidv\-䧿 ��#%��1�����خE����'��b�sÓ����e��qX���������Sb���0�\*ÎG������0�ã�a���������)�,ֈ)�*�A�$���ϝ���+=G˧��s�f3�m}������
0�ł+�5��R��H��v��2��1n��'�<�׽�~�:~J¸�'9O��׃���f/i��4�x�q���f�뛿r����7�++����&��q99�'q���r���!�y"�B��@�+�*�<q�ˣ��5KO�>�~�j����㫻�DS>xj#
7���+������ ���
�?p"�R��ݕ��>T>���N�.�Yg�)����h�	��6��]���s�s�y���e1=J�B����Xaf��v�,?A����1 ����}��h�Q��Ӣ~�E63�=+��}�4�612��=x��L9C�UDw{����V�+.����;����W���8u�o
��@�I��WƵ�Vv��cBN����:lV�1��;tkwv�^���K�5|�б&z�U�}:����9��� ��m��x� ͅ��5����wy�N��"���fp��WY�1�j(w}��C�)�Γ{�1�qS6�'^�A�꒹�8ge������I��䍈���mo4h���1���[���N�;m�c���7�D�j����s�wzs%��0���n|^��*h����O�Vg,���N<h5��Iw�+�+�m�=��h�ŕ��tM�75$l���9ө�[i�S�bҜ�ǽ�72�i��g'�O[��n�MBA�-ByԱ_l�7�����C{��Gյ�;��)`���zs|��;��������;���iY�K1�����+"�Uێee�EU�����m�,DV*�-��Q�F�3�(���%V1�[EEX���"�Q���X��2ш#Qj�7�߾���{����z����oE+Z�����=�+ߐTz 
R
��W���N�v�+Cb(_!��$R���^�FO�V�c�"�Q�j�'U>G҆���xn���U�Lo�j�10�:�m�����a��p���W�ơ4��~Z)*���8x����W5����L�5�ǝ����yޯ��iW�C��9�����>{��A�/� p�a��F��'�m
!��c� XD\8�H_g<�j�<���y�?_��e�Uu�iC�7����\������:iO��q��_}��#��wB�o'�T���ɱƦ&~�/*����Ħ \h�Cc�|���C]��'���g�`�dW�����Pi_v7~�g�<(��(p�^����>p��]��*
�Ǣ�]w�_p������.%����|֙Y�{����OyC[�O��mֿ5�U��V���4x`�<�W��+׸��:�L8���t8��kutRT�1�'wVu=��^c����:{~�U-�f���*ݶ+�֣�|7��T�{*{���Io_� x�C�B���4!L�G��qYg�~�������~g���[=�毾�Ǐ�PҤ����y�a�L�S��~O^��6�{vS�E[ V ࡯��X.��;�r~0v��Q��e
�Ɠ��U8X�U�?1�i}"'b=uI㉉���9���sϽ��-�M�Q��b��c���ڹ6��°P>4*��SC�>��.�Y��)kŻ�ĝ�wn�#� ǻy��	:�>��8]��Ӵ;W%_ �y��:=�{�h���������|��߷����Q1����/������}ޟn�:b���������Ϫ�v�]��R��X����q�CV�Ш �^�*�>�G�߹^en!�/�5l�A�:*���*��VU+W�-ڿ��wA����"*��8����V�AG3�O-�mH~��`�>�j�4 x�L�>b�1��i����of�0��H<�S���Z�Q^Dm���#g�[�udm��ĳ>Þ?\d�H�d\�`�
<�~��;����@�#�MFEx1�����!�o�����Dp(�n/�a����kFw�
��Z4xR�j��5���t����ϓ��N3���֝���X��x|�x1�&��C���h����׸ֈ+�*������AV0N5�i�.A��5�1Y�>t�s�s���w'��y�s�L�ueO��y���4�|4�E21�,ז�;�AjG_���U�#�{u.2��x�ɝ'D�n�ui�iZ� zkS��G�<�TD	�80�L�U�>�T��*٫}��Y�x_/NS�OS���>�}M�����s���2���M�ɧޞ���g�����>�q����5��_���x���p��c��}a鯌/�m�O>�8��@6A�3�;a�D��@��xFƘ�F�o�_�����6�n�<g��LS�7뼙h����g�_;�i5��0d��v�Gr�J�����uȴ��ӛ)7ʟM�:���fΏ�����ϳQ|a��g�N~�p��o�I�.ҤuR��
�U��ۊH>�I���x���Ξy��ͯ)�Rb,�}���<�x|�;t���m%}fs��9P`�*a�����AT��
~+ϵ�Χ��۷�PҰ��S�;��4�i��!���<��0W�w$<��>b�SMt��}�����Q�����4�|s,e
UrM
�C��{�bڊ��n����
"9�$'�Ϝ2�t�hq�&:37�r��� ����>�}����ͳ�-2��]#\)qb����
�`���&�+�����Xۢ"��u�RX�g�1t)�
w5��&��XC�b�|ǁ��X9�����t���N���(�t���sn�v/ω�)��)*�^���1����]�g��M��5���N<�~|O���ę�|��<�w���ohu \\ǥBg�i�O���1Kj��������aUS��m��Bw�X�\qu/��M���\)�C󜩣c�����j�*�V�
`
����}��~x+�z�h���+���VL�%��T���N?@G�����f��YB�S�CX(�"�xk|�.����+!���+�޳L��N}M�&��q����T۝�8/�%�}��*���=Q��~��f��՘�
�'��������v�![�B����=��t�wV�h�:��*�p鬃#�<���)9�Y[h��Y��GMj�Ͻ���F���'��OwO��^0���w����>lF���8�}Q��-;�����I����x�������W��>���B�ѦZ�4���o�t�_ATG�(��4�IRd��OS�h�_|)�>�8ي��#Y��� �>?xR=��w���ޏ� ��k�&�{�������0H~s#� ����3�YW��V\�{J�G��@o{�E
�T2����=�]�1�]k\t�N��YSi8�9u�K��� .�
��)z�u�sS6��dj�8��2
�<��;v9˝3Oan���L��z�8PαQ@������ww�6�
Uw�Q�����ö[���)롻X�u�W�.�s��`ta���4��S]H�be �eh6Gj�a|y�t�e���d�w�`���Kޣ��?�#�1�����iP`��6��A`�ֺi�fri�n�����5
Ds�zp�ŉ/B����YmIλ5�	ڂ��Z8Z�vo s�zL��f��Z��r�f�h�/fgU���t�0E��q=S;��oPy>�DT�J��d]�%�w>�c\6B�dR�!u�5��P��85Bڇ�}��з!yF�ᳶ��PT,��ް�y4l\��ʼ�Ğ�YIs��������{GV�;h´D�(b���R�PRҊ1\eQE`�� �dTWm�E2أh�����E�F�V�J�eT��([Q�̡��l���J��AH)��F(�\a��q�`�a��ֳ����+k���Κ����R����k��I#�o�p(9Q�����m	T�!)Û���Z/xy��Ѫ�\�z���נ��,'Q��Q�|'��$o^l�%!��hf����A7*���z�n;�O&����r��^R9\re��;�ӝ^}�nV��7�W[�4�,�W3���Fo��c��L���g? �b���3�sx��4����������%|�m���QQ׻&Z��_ &��^O����S|�$�M܉�>Xjo�_9�W���vd�4�����r�u�zw����񊁬 �ώ�b�Y��vzF{"sU�x�{2���塛Ej��'����r��d�����P�;*�l��(���]B_=o{KV��~�GU�<V���۵�*3�j���c5ߤO��\�o�w7�e�8E�L��=�A���F"���Y�Nٝ8xd�V�|"�ݵVN�����2�Q!��9ժ��MFJ��*{9�³R��U̚��YG_�ZT�Ul}�9]��jͪ��}qT�Y�u�#Hiس(��S7�ް=2i��wEE�͵n�F��Q)��ą�n�"�BQ7�$������6�!�oy���F�k}N�[Ӟ�'�$k�&Beu������� ˽���{��O��w=����;d�E���l����՗�xEs���6�t�[v�.��Kp)�Ȝ��a�X�fk��+���'/xU��\�<���ܚN��d���Bמ@��__�԰��#�/�#��b�Vom�s�xub>�O���ov��-VK��C�{��˛��}�^Ci��x���2���S��rYc��N�����16{�翾�����]���Ԋy|,��8�wJ�ެί�����S�KAWi�E�v��m�����Q;.��@�Xu�.w&��w��z�>�*�^>����QdЇ�nؗk7OM��nU͞�,�Zl� �p�c�)��Wy]+�h��1���E��Y�w�ם�c*wp�Ϯ�8�a�>��Owg짐��G{o���D��FT��ۡɽ_�@��/6q��@��\j�\�����2Xr-��Y�{�k:���kr��Jc)z��]g
{Ew9����؆�G�"��-���~�������O=��Zx�bu�^{���A��@{��Šz����W��o��j_�G���i�2�1�m�-�i>K ��|�ɖ�o�G��{�B�k���1lq4c9����)ּ ����Y�^z�}�JH�WvF_:Z��6�D[+���]��׶̐�l�GK�۪��K4zY�3=[����vI�.�o�,c�œ���8J�j֫� Ok��(���/�oս�fd�wV����%8ᜎw��Oh�����E���y�����2Y��-���e�����Bp%���W��ۖ���}�����L`um��Z�{��ǓE�����n�X�]��؞�u��z����&��6������*�zj��gFC�̈́;���1���=�kË������*�a ș���-/Z��l�����g���4�����O���=�8���|Q��j\�ezuQnW,mw�5
��\�V�J��pN�O6���9og0�7Lis���'i�@hCg���*�l��[����1md��j�TB��q͂ �7��A����*���v�O'iuu������dܮT�$�j:)�3�O#Ԩ_QW¤�k�=�Dh��a�^й\�-�K;&?�WIٓ�w^�Qp��ޚ�޶����{a�F)\��ԔW����,���#n��՗�3y��7����J�5f���SQ,�]rZ��Y���Rc��Sᖱ]���(!iWvG1�>D�/,#�]��V>���j�mn�]iZ2ğfFA������*�m����AS�>���Ur� �b�2J]`��V~7r�$���!J�+̄�RT2e��t�(��2V[F�c3v���,�� $�!�2�cM7iՈ̴J��[Į�VVd�Kp[�"`���y��e�w��ь|�E+
�F#Z�m�5*��2�,7.
V�(���
T��T�U̆"��\����[*V�+-(�4*��RS)QE�S��D11U���Z��[l+1"±V�pB��
��J�`��QJ�����ڲ�"�1�"�1��\�\e�++���m����k{�J� ݺO{�^_)���:��S�5v��6etj�`�~{� �ݟ�N\������+��ʹ�ą�Z���p�B���[�A����Ҵ"[+�%�����[kā���x#=}����G_�
��E��zJ�Cܽ�-.��X��@������fΗ�_1�?E��4�נ�+-m=�]��2��!3�4@:"������t'Bj����yg+�B�MBD[׽�/v5�p��4��s�欝j��YK�*��ͼ�K>�5���^)����W���6��5�.������/.!R�z��E_F�^��4׎�ɝ]����q�F@�eU�_�2��ֻ'�]4.=��7ճ�%���v??�|{�
[����t�}|�Y�G��[��=��MU�������n�ci����s�+r�c}����/��b]ҷ�v5�O�w��.��h.:H�#e�>��L�J����ww����;��4e��J���f9]hl�NŠ́t�6��q� |{�ݵ���户�pP�!�hwʼ����{Jw�"�>�:&]s�k���+�ى���~�?8�_R����%n� ֬˕솽�6������+�ED��.�ud���$,SqA�Y��O;E�bFED����t~����M�z9]:�Ms��Sf>������7����^L�E����fjY�W�-�ӌ�f̏o���9MX�,��V�ut�T�ݟs"�C5�m�)^�ILe�aWw�+\v�uĦ׏���m����)R������	�/[�s���ݑ�B����
7���;=��Q���c��;܎}��q����㽃S��!�m+^7��_��i-�4�>5���q���룔7�bwU�b�����zQ�X^�B�>TIo[�Ǩ����zr�����a�#�c8�R7R�3<s6��[=����ܷ��{m�r�h[��j
��:؊�*qq�]�Nd\a1��^˖�WM`�T��Q���T� �1���O�k� �+��>cxѿ��?k5����<����h��R[��<�J<�Eo��gy�7V���b��UMku����vk{K��k{!{NP�6֣���ӹ�p��D�T�x:�Of*��R��~�<��y`����y9��ӓ��:�<����>�6.�S�ޣ��!�lF�׵���s͗\r���-E����=�R>ӹ�Cpj��p=~w�G��;�)��^/�&���S%iy������t|�R��q�Fr���}�����n:���;�T���}���_B`�@�ֆ̥�6��'u�s��'s8�D&c�����Jv��9�˸SZ�US�$�<3��t;yW��ߜ��+�L��t����bJ\ڽ��af�)���lhC�r$�x���ɾ>���\e$���k&%�ǒ>Z4��]L�;N݈3�<�e��hsٝ��	w)�#����2{fjO�����%79u,�;:����Á���Ѩ���1�>n�qOpK�۞z�uimk;�㊲8z�%۱�����Ӈ�'n�3�,[/�'�.�D�<��=�`kv���izd�U8��� {I�z��ɜr�2j{T;W�o�|x=u�۩����F��o ~S�{��eO^�&u�Gϡ��%h�uH뷈(�wj��	e;Z�[e&�P�푫j�dB\�Q�*^t�[1��C!��+*[Csg(�iG��A�M�y��vT�)oWz��gL�lK̜Kwx�,`!X���ܨ�;(�Q�NB\��I�r��]���Q{��9�8h�j�g�EM�G5[,�����"��<��m�3J�Y��9tB4.����]@Z��R'+3%%jd�0e�P��a4A+,��n�1�r�����F�Ph]]@�9r}���Eܔ�e3�A����d�C�v�`��w��Q��+���u��B���ņ:F�q�@�l`h]� �!�i�a�cV�K)�"6�0��5�`������K �N7�:-��((+�**+V&�)�h��(5�QQA�Z��F�QD�-��0VY�&Z�D�ニ��Vm[(��"�4�P2�b�����ԣ��&P�q�
��X6�X,+(�T�T���-*�3*�,UU�Lm)2��T-m@U�«
¤QR����G�\�*�v�HN���_frsl���]�'�q��<���i�
�l%z���N-����.��qq��t[����ٕD�:g��W�d�܊[K�;��U������xV7 9Y �ˡ�1�x���CWճy.��y��#Uʃ�����8�:Ն����S�Mc�Wf�r�f���睢�uՎ��ȕ�o¶��yf{q��κ��p��;ىb��٣+��ʁ�ǻ{[��e'����s�N��.^����ț��`�s�x%�jr�;|���@�r[�m%X1�Ʈk���.�����ʃa�Iz:��^'ᅦB��]fmX��E��o��\��q�HK���1�=[w��gV���}���Y8yG~*�����,8-0��g��ɉ�/�4*���Y��P�oq�Vqu|l�YEW5c����O�[V/^�����I���=(�@n�jYʜ�wk6�M�ֶ�a�ncp�I࣮�I����6-AJ�n����͋J&�Wۣ�W@!I��Cv{�o���y�>�#��{K���Zr���=�p�0x*�Z��s(^츳I��Cs�[�j�N<�ib��U� ��*B��:�~���vȨ�j��kx�{˴�մ�|K<�G�n�i
lL�;�����Ҏ�צ��T^�w�_�!V����<��eڒ�w��`��A���r�e�+H�G�J�Mz�g���L��]ꍎ��'��Km���ʏmP����^[�tڱ%OQ0�n�b�ę�*��xr�M��gae���If��eI�Ӂ�>P��ɫ0�EλC]��"T]Ҽ� {�DA�L魗�3+���f�-��@�;\�&	9�G�`��돻m���=��]y�"��,St����ݻ����Y/�E����仵�t�=�{��饳y��\�v�2���P�XPݕ�κ�fm��k�^��oNu�f��}:W����:y�yfV�}���Uw�A�î��?#g��M�{V���)V�)W\�4�^���ھ���j��F|`�6��z��U�4z
�<gJQ{5v�7�r�'"���f߽��/���H}�*��G5�$���,S����J/v�"<�[��UUڶ��FC���>�Z���dJ�[ΧAևY�E�V"oN�^M��{��Z�B�-�φE2�:�d�9���A�&���ݪ�jp3gdu��,	D��i�<��u�l�[��E/}&m[N�V��e�eq��G|�;�Kq��'F�|�c�]�[7������k%��,4!t���qH���6����Se�V�:��,��z�Q��ʾ�n�fCL��}��n�:�\��T��2����<GVrv�E����n�0�L��pMm��æ��_[{�jR��\�1������חuQp�:S�v�t���OB; ���[+=�B���m|n�<�<��].��د}q[I�Jn3*����}�ꝸ��~�R��]����39C8�K1��!͕�#��g%<!e�.���u��Ls���3�<������T:<p�<]i�}�<�y�h�z�������Z�t<ڙ9g���ګ����:�D��K�Y��]Y���Cͺղ$�lOcEb�}3�ɗ�v"5�|>W�ma���H��;���Zt����UbM���-�B�=V��̓6��d7���k`j:�':���Ӷ�/WW%�d����L��m�>ػ��~�3k6<5�hw;Sr�ʡ�(��e�����:3tN��m��X.�c3e#3��EN�$��8��q����5�@�,/h@[ɌPTbxk�`��7d+ �j��j�)����sfu�f�%^Ys
wv�&���X��LL�,+�R�A&e�ˊ�L�yF�����X�I�1���eYIf[����@&��-�e1K)�,��n�Q��ĀH�h��@%��HE'���wz��y3`L,b�x�0�7Q:#%��9c�R��h�]dDʌd˭��U�%`U`��e-T��lXT'r���F-IQer�T.\dY��b�Ee`V�UkDdX�Y*J�fe1��e�J�,Db�UPU�4�l�`�*�P+	P[h�)�+����~������Ï��7ِ��ft���_��P��{yq�[����D�S�C���F�y*�����<[�f>�s� ʍ#0y�1�8��ͬw�!Zuh�KƖq���"�-=�5�� e:�2�xd��x�n�) �	��>�|A���*���B�jV^��7+۩cK��ޤ��"���!y���x��o�o���������=�V�<;���1�T�5r�u����U_[�3�\����T�q�5���1�{bV�͇}#4r�̺��4�u�3�-b�_m8��Ӽb��q�ʖ��c^o$���<ȝ��p�YHv����9d��v�H��9K��k���g�H���:�r�9g��"����;4�뛌����9��^w;ݻI$����Gp��b��%Z�0x��,!sZ@��7+.��G*r��Y}�F�l�c�1|��nT@����ܟ��T֚�nZn���kd�_%�n�{�v��o��T��i%���T�71Kf�J��b�C�Z��tv�S0*f?w';0�Z�5�;���U���f�z[�H�6�WF�'�]�d]��~����+y^�%��c>�M��}�7r
l�{eF���xcwY�V�01̔��b���֞��{c;�rT��sPy!���c"N���uu��Y�ʆ�؎�7]�J�Z&z&y�Ҩ��a�. ���}�fN}��.s���eL8�(�4���]u��v�5���R2���Ә�dL�^��:w}ޭ�\����VT�EU7�S�cj3<�.���*Pu�kl���%���ԯ[��#��|���S�v�SkN�K���|
#\�]�c�of���}��668H�C�����}3D��E�t�U/V�\;��i�՛���Z����PT>�N���8�ж�(~�:L}yI+ν�-{ P>o�������pL���}�gFM/���nɣ�����V^6ι��>��������%��T.M�mI�j���.c��
�kB��aQ�a<6��5p�qb�/� kjle���d\��y�"�j���l7q-��砛uϖ׃5��s�g�)�%9�y+Gdj�T�Tv��V�6��y��n�Gc|À�>���_�˺�O�v����ά��nT��6�.��`���=��ĩ]�ӸgW6�jt�;�1wV��y��N���pq�K������á�����r�p�1���3�܎r��
"�ϯᏋ���N"ҫ�{-�咰�'���OV5�+�^����hJ�~q�Oj�"��F���9j�{n�]��!N��ݮi΍���C��W]vH<����wM֖7�|���t�Hv*��	��ŭ�n{ff��������z��x��/�Ҟ��A�s?��+���ע���nr�X�������8�w�7�r�.�̮�k��G���\��q��y��nF�s�Cж�,ڭ:�¼R�v��'�5+E�8�*�+���2T;;��VsO�zi#��Ÿ�m;��:�޼as�G��"&��l�;2����C�5�R�{�<�m���Pz��nQꎥu]�h�/%T}�u��/�;��[���2Zx�Z�Q}wq�_Ri��}��z���3W(J�T�dW\�^#����!tñ�u�� ���r�\8�e�j�/��]G��8��[�3]A77",���t\�s�o=�tݐ(�N�^'����ā����6�6[u�W<����o3Ft��d	�7yN'�Wt�۝>Kn�"�V>�Mt����5_F;
�{%��|����'X�4�a^�Bd�y9L�j�)]/}�YݣC�Q���֝�'p�b�,��ظ����s��N�؏:��%�M�<U��[���Y�+Ryq�̭�ʉ�=�L�ҟ��t�~��α��U�93�5eu6�pl��v�}��쑬�"�w+k�u�(3�Χ���v+�m9ӰR����YJ�"��Y�r7��N��@nG�f�u0q����&+]v��n-86XC]�wQ��P�V���g��qp���aث�����MK���k3��t> 
}h��J��Y�#Z�V�eE���m���q�Th�X�d�
�!1B��8���bJ�JDJ�ذP�U�P�YmĨ�
���"�*��2��q��Yf�GE.���kK��PT���e��b,_U�'X�gz\�|ҷ����^�qP���1���7L·L����`�ڼGD����":�G_��ںr�ۭ�;�i7υ���:��NEҽY ���8������O���{0?"�0<5u�%v�v�f�iߝs�T=��]/w(��YN��W6B`0�}t���(gwrܝ|��6+��{�k�;0{՞�������w�jC]���%W��0�f�.:�=#t<��ܕ�,��+�u���9�U��u�Y�5�*�:U՝8�ys\�w��T�M!<�ő1u�ya�V�t��{�*v��3gHUΰP�M��z�@&8���X�Ϻ�:�>a�7�w4���&gu���J�K���k|�wӆWM(�odÞl藾ʌ�#ϥ�������C�)�G��*�M�OSG������n��J�rv��*I�f�\���+�/�-T��e�D�!���P��}��*2���i旸�ܞ�.s���[���kN����}�2���w7LZ�����d���Oޅ������g�u��yjϺk���8�]"�s���6�c"�K'�V��\���Z�
ߒ�㒢��ɇ����n���_�_��W�X�5^.���|#4(�)��b��'�8��(����c'�N�i��ޥ]놷e��xD�Z�I!���*�xԝ{�QY�1���Gi�� �S�Tm.U��Y���$��T;��v� ��x2�]��j���T=V�ul���U�((}��܌��Η�*��\��I#�#�]������[� �jfL�|���{]��Oc�Ⱥ��S-�����^��K�S4�,�]]�g�]<9�D�!R�{��]bO�g"C������KW4�D1�v�3K�sʲ�·C��/b�����w�sC�f�\�A�7L�i`v�r�	u'p[}w�U���2f�g$��y���xS����O��7ϡ� y}Py-$�ؾ�F���l���:2u����r�ҷiG�1�{[�s�@]�^�F�~n7R�;�ڽ���Q��w���9�ۆ����9��sU4�obD=��۹����g�����8j6��*���P�(meO��z����a�<͍���&-k��_9�%r5��>[��D�+k��JW��G���\�J[{�[�B��f�⋣�5��E�--w^Z��kĴ��S�x3�#�����b�ۧ�>z��U��R����m��=iٝ���󞜦!�N�c)�ϵ{��+w�\8�q�-��p
�؝�8l|!]�5�;"��:�b2q�(��Q�N	��{��bc����}�w,��o���+�Y꺃.�>�1����8���EC�kO9a�s�����Arܚ���뜩��������t�\�l�4�;}MA�u�6��P�LWH]�]�O�2st�ǽڑɵ��2���\"9rY�W(���c�Z���7kPc�y[���sU�<�fw�{��B��pc�;]w�#UW��o.�RI~*��g�>�5�*K��"{��Z�zF�W�-o���ޛ�7�{򃊋�Yo+��,��)���������*V������q#�� A�ؒo @��G���-��,����������7�_!�  @0��n�JkQh�S]� x��`u�N0�L����WH=�'
��F1l�3��S釢`����������R35g����<(w��y0翗���B����AF�Z�m��h��W�f�}@��A�@�N������bKa�c�ŝ��A�?��5�=hH��;�ɇC���'�H��  �w�l��v�"
���)��W�"�8�5@H�>�T�/�e�)vN�CMZΐ9�b.���7�X+)� �� @�>��{��?�8#�S�_��4@�;U����νd�����gCYD� ���� @Ũ���½6��e����Đ}��ܖ_\Yy�j�Z:��du����5�dc�!� �;:$��0��U���Ði�L�d��5�St,��h>�2鿙]��"�����t�̧�
�q�=������y]��p�>�&4K�h�2 ��F��q�B
bo s���g���D�9���aո��H��T��� �P��q0>ћ25H#�\9E��BАд�u��Bk�����y��`����29O�b��_iJ]0�|/f�Gu��M��gS��	^Z@�	�|1�Ff y�a�i�`���l�f� &Fg݇�	�"椟��KBϿ�IUi�Κ��4���+Ͽ�$v�� I}h�b�g�ꞥ��}o?-	�1sfA�ߡ+D����$x��aY�	s��ϻ��=����g��e��2�v9QU��a@��[�bD�
��ք�4���j!�E��-w�y%��5@�� ��0/Q�R����4��ߒ ���pMIP������d��-�I��:L�"�y����m��rE8P�ĞЎ