BZh91AY&SY]��j�l_�`qg�����*����b@           p                                �(Tٵ�d�R-�S� �                       A@�           ��U*��(�B����
�EIPU"�*R$�(�QIR��R���T��H�	IB*TJ�T
���R  �(�P�$�*H� ��:�ݸHNcG֗��T=��J��"r�@wn�@z:;h�s�m���sԥr�*� ԇwu�   ���G�AO۾��[މW��R�����������z'J�0���=+y��GA��34��՛A��@<�\����`   0σ�*�����{o�J;�=�@eօ�G3���Z�U#�s�*d�ל��t�`9ڂ�ѻ4'9�Ivy�P�j��4�i�   `|�t����� <k�H3x�C/M*�����E
+� b�9�p�# $��!
d����E    zxz�UR�B�R�H���mQW�s�l!�u��t��w
���Pf��f"��p �ΕD����@G�=�s���9�4��p   ��U��
`{>��f��
^���N91�Ч{:R��I������!:p4#/Y��
:t�י�:`   ��ﾕ >UDT�BJ�$@����C@)�J�iQ}��h��x��s��=��z��vr r���m��[(:   ��J@x<��FA�L���1��s��9R�v�.`�UӀ��� �� p   �)( ��%RB)J�R��)�)��� �����Pu��3>��#S������BMȎm�si��`�   o�J( ���c�Gv�������Jh1���}��뼪� ht��1�@9V��|  
�P�  �"`R�Q���  �  ����J�  i�     �ѪRS��      ��Q�J0       ��*j��      )���&LF�L�<�O�<P��h����~��$���_�Ȋ6�����I'0�N�&����

�_�"�
� �"��"�*������ *��C�O�w�w�_������[��6����Z�[m�����^@D_���6R�􊊢/0�ݟճ�`� �X6�`�%�m�lb[ؖ��0�L[`�ؖŶ%�m�l��i�l[`�-�l��1m�l[`��-�`�*B%�
`�ضƘ��6���l[b��6Ŷ-�m�l-�6Ŷ-�m�l`��5!b�ضŶ�m�l`��[��Ŷ-�m�l[b��ض��-�m�l�6Ŷ-�#b���m�l[b��6��m�l�6��l[b��ii�l[b����m�l�ض��-�m�lضŶ��-�l[`�ضŶ-�m��Kb�ض�-�l[b��lZ`� �-�m�l`܉ �l`�ض����[�����-�lK`��6�bF-�-�lK`��6��S�0-�lK`��6Ķ�m���b��6���m�lKb[#ؖ����`� �����6��%�m�l[b[�6�C�Ķ�-�l[b��hm�LK`��6��laŶ�m�lb��6Ķ�lKb��6��l`�`F�m�l[`�ض��2ؔŶ%�m�l[b[ؖ��%���%�-�l[b[ؖ��%�-�L�0-�l`��6Ķ�-�l`I	lK`FĶ�-�lK`�ض��-�-�c�6���m�l[b[ؖ1m�l[`���-�lKb�H@�-�m�l�6Ŷ%�m�l�-�lKb�ض��-�m��#�6��-�m�l[`��\���-�m�lb�ض��6Ŧl[`��6Ŷl�b��6ŶlH�ض���1m�l�6Ŷlb��� �!l��m�[�l�-�[إ�KbŶ-1m�l[b�ض�-��[��`����� -��� -��-��
�[b�l@b�r�5!�"�LUm����(��Vآ�B��F�܄Qc��[`�\�Qm�-�U��
��-�E�"��� �lEnB(� -���Dd�nB
��F؊�[`rE���V�+l #[��-��(��F��`�lQ)�[`#lDnB"6�ؠ�`lAm���DF؃+l@nB"6�F؀� [`�lTnB
6�F�܄� �b�lAm���E�"6�F�"�lTm��H@Kb�S [b�lQm�-�U���V�"�lm���Vت�[��lDb�[b	*��"�lTm�-���� [b�lU.B,���AV؈܄Um�-��*�!blm����� � [b+lTnB(��Vب����b�[`rQ��� ؂�[`�lm�����E� ��V؀�V؊܄nB�R�F��V� �ؖŶ-�m�L�-0-�l`�ض��-�)��)�lK`��%�m�l��6Ŷ%�`�ض����m�lK`��6Ŷ%�m�lH�ؖŶ%�m�l[`� ���K`���m�l`��Ħ-�#`�ضŶ�m�!b��6Ķ�m�l`�)�l`��6���-�l�`�ؖĶ�-�l`��R�%1-�lK`�ؖĶ�-�l#�6Ķ�-�l`��6��5!`�ؖŶ�-�lK� �ضĶ-�-�0?�EI?�=d����+�Y|����yJ$�e�&$sL�]T����Gu����^�62�&�<�k�t�W�"��5)�T/ଷ�C[�y2�,��
�]ݼ�MJ���d&,X��[�o��{���34i��<(�\R��	�܊f�c�KFE%���op-�[����Q&
~E<��\��u�ǗZӥ���ͼ���4v�&��w{��w���peL��=��8��WWU�R꩸m��ktT��Z�L:L��r���<�X�{X�j�Ո�eì�*6�կ*�a
ެt������͵�����YWe��Y�5�D� �bUش1\w�cqe�j�1,��0�a	�2��qLB�V&��܂�Ռd�I���q�2���5��&n�f��]Ú��μZ��=���B�i�匉��!�B����$hv�j��:Bh�-��:�f%Y��[���rG7^(�����-Խ�)��e�nY�Z�$��66	�F[���)I�:��h�����hs�\��UmU%�r��;(X��s%��qE0�S-@����f��є�ᅷ{/�5N�	�u��kƑ�6�L����)f�k.�*���,أ����Hs��2	D@����:o�hc��/c���[V�\�#r�b���C��
�S�[Ij�-<�~4���Ib���бV�N��	���Yەot<�Sոp�[���̳��r�jI7�؇qZ*��
@�e	�%���WB���yVQ;�r�L��j�a�Ŵr֧R����GH-�(Z�R�k[��*݃0mnm���(U��q�4aBmԮPnPZHKwU�=UY�� )�o7�%f)�KnѶ*��c�ڧJPD��;�w�Q�=�,'��ÇF��n%c
4#U�����&^�t6V�:,�D�袶�XV�CE<^(�!ʫ�J���a+q�vb�#�x����)N�dXv`h]�����;۫�7�%Ե����A2&em��Ӧ�^R�+ ��;�]�J�ù����[Tq�����y�V�t��T��b�#ܳ�oF���7[bk�ܥ��э,�L��˕ou�[��u��΢�p*Ww�d	�ZWj������/�c�1i��V�9t]�n���.�ah��bV�K���=pԞ�"ָV���L���Z&ɒ�V���k9��sJ��[ێ]�ֈ�Lr���cK�jC�l��nV-́m�S)��
)�앵��;(\oY�oeSx��Y �.J��n�8�n��J�r�lb�ae^=�3C�J̣`���m6Z�����qd��WVY���țwgjU��@�Y%�{�9,4�2]S��nͷ!ڪ�L����&U���^�.���K���ne�1�n���v�X2�L7
"Y�	���n�'�N�Pɐ]�U�+C1eT�Zi�u��v��T�;B�D��H�o:eUav�f��$�������-d6[�r�U
c�7�j�*l�9�d�x֌w���b��x�*����̝�n��[+���8��W0���{�JR�*ȴ�i���\p�P���/�3]�W�T���V,����Kj�įN@�k�s6�fZ��d�uP�V1���+B��*�BU"(�Am`��
��b������x�m�uyL�6���&�b�4��b��!+mZ�������t������L`uU��/�;~���h�6Rʔ�!P)�Sɵ���se�h+j�"�.��J^���!�G�l-�QlUi����+5��m�r��T��X������H^�u��DA�mGGv0�b�rR�wm�4f�pݚq�m�1���jCW��W��ͭpI�Y�7)n�7.Lr�P�xC�܉+!�2^Y[�.�ѽ��#v��-�mc66��fB�n�w��D��,V6"gSc.��`��(]�'(�m�5�V\��"H+,UY��]:��t�]Bp�[�ZMG�JV9WG$�����K��V��/gJ�3�û��PB���-��<�KK�J�CM4ꮊS�u� �F�Vb7{�!��v�`Q]\˺Zݼ�PB�,�5k�pf���d����M�b6����h���۬�D�\z䷴�k�&r��֪.]e�:%K������ɉ1
�hA&��-�*�m�P�.��3��r�U�O"Nl��@�޻w���6�t�aYyZM�B�d���׺&L�/`#��R�M��t������V+[���#��Ɛ�GA��CR9�nX�Y�]�!�r���s̱Z�eĪ�������e̴E��m�j�;7��yz؃D�F�����;d5��e���t��*�'�Yױ��x��ٷI^�i��n+t�Z˪�F��KKjn���3�grX�e��b��{�Xݛ� V=��ݑw��so<�a6��ǵ�U�*�ѱ�7n��N��ټ�����Bnb��c���$��c�snav�ө?8��٦�ئ)�m�Tōd.�+a|��Q�#T�I	�̳t�{�V-&ٞ�Qbw	Komf�b�!���7B���n�{KI��j�U�ٻ��U�.�]������t't�H���p=̪��p�F\F�7� �VH�X�˳�Vb�jY�P�N�Uma�-�2��M�z�_���-y��N�ͼʖiX�Jٙ�T�/n�"�0��a=�"�ì��Ì`i��ͭ۲�X��U�F�Q�6�Z4l���k5BC��4�Tr�F��V��)-�2���s[t����禋��C`�ۻe�%K�D�����*Hkv073j�Vǌh�P�Ǧ�\�囸k}e��y����n��f��uA)Z�ј���+���Ӏ�v�,��w�Y��;9��j�<h(n��+˫*�YǠaS�E�巶7S��cM���GAr��kfڪ`�5v�ޥ���z��{i)�4K�2���uiں�L�JH����v��370SjyЫ��چ�M�Y4Ҋd�
lD�+S��Z�/�ȝjZ�z�n�U7&�۶����Tj`��x�H��[`�Ғ�^�^b�/M�ɛ�1-A�J�,��XqI�`rH�@*-ʗCL�Z�Y���(/��ctn�苛
Z�I�d7nƚ�����d���LØ3w$��6�Y�.�F[Y�7�bu���V�/*�X����7{H<�����l^��ṇWG"xc��B��9��P&rW-��B�%�	V�UCf�ǲ�B����S{Z�"��v��LU��ùh���Y��6��=�אccF
7w5V3m���]��kI9�Tq;lZ=8��9��"�˵"���X�r��]�U籨�ΫO&�8�M��n�7�
YH^l��!�={����-^ѣ�\Փ,L��ͼ�fbT��V�G.��&L��v�-�l�z��������6��^o/*����$�P#`@�˪F5@����P��t��b���N�x�ѻmX&�ŝK2�y��-����&V҅�p���[X�%�*𓸘���e�(!���%S�UB$�2�Ci��W�]���%nɾ�u\�q0e;�̀�*�q�u�W�[S�nJ-���BMq��Z�ur�n6kL���ܭ�s�lze�2��P�*�MM
�6�ՕV֛�4���u[����e�B
n���AKǎ�˨��o��S��j�Z*�5Ktne^;:�FZ�æ^f\Iۻ9��UZ�A����r�f���nP�ǋ0e3�^�{�q2�m�R��w7w�-(m�����l`4���Mʡ��@��ڸ��۽��'��܌�b�ۅm���&�������ePU^J)VGS�)�)
�[����ۺG{�nM9�(�"Ģ1w�u��w�i�9����el��ًuGq:9�K�Y��k2��ګ"��;���X�de^A�1<ķ����pY�*�<lܧ��
�v�#.���&���m���jˁ��SM�`2�t��6�m
�6;AU�ߍ����y�6�������{���;�9\�n�U�mn$l�
�w]"60Q��B�v-%�(�ɧv�Ee:��.L�8��:�c�/�w-؀�+D��;6^U��'+wΔ�-ܡD3cݒ�#���M�͉�uz]�f<�Udq��܎Xǖ�nͅ�tn�
"��h�.�6�[X�e�;�Tr,�z	�L���X*i-�{��S��"֤-Q2\Z&/c�j���H��w,ݚ���l;up����+=���4hB�Cm;z��v�Uݽ4}��ʱ�+0JǱa���ڳ�T��`���f�k|^f8e"�CZSX��z��Y�Bu`��
�\��o!��^ѵ�0[f̱zki�y��G�H��rn��F*fi��Y%:z�5nYa/4�9��(�`!�r�ռ��[L���AͰMe� ���R�Ʌ�6�mhw�H�Z�[��^�b�V�,�6y����	O6l�{I=l�E��u��(̹s[�mlL�
�W����w�'h:!B&2(�Ǹ���mԆ�n�m�el�����.�MZ�v��ca��6CN�편��d�kb/%�t,�A+���a��]ʤ�Y~�¢�Sq��۱U�7B�@������F��
��:l)�F*͛6��n֣��5wI��ى�ʕiUU�Ԫ���k�DV�e=H�˷a�oXnK݊���Iڗ�b�X�K�%ܭ�b��h�Eʪ��)Vښ4�K��B��n$ⷴ�؎e��H20ڿHn��Q�Bc[y�a�L��V�x��5���+I;b�S�����[��W������G���l�����Je-ӈ�j�B0���wlf
򴱇R��O��2\ӹmĖ��w�[v7j��;�F�f5v3eMb���f1u�t�(ƥn�e�Y�U%x�ܳ�W�WA4kwmkhJ$K�s2��WǒL��ojvl�&kڃNۊ��b�j��v�n�7X�.�6�U�0�*��FHve˫Ũ��UhjיĞ��KY���Q�
G�w]�p�s#�f���)�i��-1dX2�q4/6���VaUj[Q�JY��8�����/}c;
i�b��%L�u���I�F�J�lX�p]�ה����"�Q�nc����T�B��mJ�\�U.
]Ao�Y����������(�
%Tw6�e��Š�ٹ-L+g#AfeL����he
����T�X��z����q�Y�����Z����n�Uɰ4�һ�s2��t��[�J�(�(��C(�Xt�%E-�n��Цn�i���C�%�q�V
���w`�����'�,@��lU�B漇�l��n�-�Xy��-�e�U@�7j�`Ӓ���1TX]e����8�ecde�p������ň�۪�ۭ����!���\XVm@��n�������l��ڧ+��M��O���Sv`�=uC<�Ud�ֵ���ic���d9W�or��YZԿ'%R���cuѼ�9RftEf��3q~�ZE)�փ�U��ܓ$�sq�k��we���יW��R��,�X2�-�YWvVn�ٲWhT#"dx�+m����ؒȕ���ʀƓݦ�x`��fLͅ]i�c�:�4(&<4*ЀW��4ǠK���uػ��u�:��]�Xʛw�CA��2���'�(�3�.�^��*���*�'uY��ڍV�F��,��W^��\��`�ǵO�M��m����3+�C�P�M<�w��CŻ�R$��yB����0�᪼*��סг�"�Y(���T%�5krJL\іp�Ɲ&�X^jb�8p��H�Lw��H����cu���L�^Z��Ɔ�N��Yf�bH+f]�;j�؝**�V'32Vi7�W%���hL�i� i�X�!���6��^�C+0�Ѵ����Y�O$�rez�)�{/R�*���!��~}GA�P�q�ٰo�E�7��آpYx��m�)+�l�+n��lX�����k2ތhDwr����e�����N�;r�G��(��d&��V/sR�uH�ըZU��r�U�y�t]���]5N�Qu_C����e�z���C�䭄��	B�U+%U�73)bN�%x���$�/%ibP�)��Ⱥ��'�%*el��lɁ���O1�ϒ�S�%V3�ay'���%Ib�X�'Kt�))Yy=�)W
e?����ZR�I%�|�������(�6��\��(J��D%*i@&��x>�>/R�M�Y�)|C�0�߆�>���^R���DK�Ҡ�G��������fK���</��|�쯓ؠ�zC�`�|�ɾg���V�(�󭜳&OUu]V��Sk2�*�+J�����J�IRT����Y�e���T����,I#�|�R��L)�7p��2�ç�~�0 z��K~�|)Rꮪ�ʧ;%�;M�����T�T}���z�����'���l !i�Y})\���)F��Q	Z�O	J}?%@�ޘ�]��[�R�z�ؑAIZ@�H^>��^z�)JW����WZ�nZ�𾻣�u�uJ��/�O=���~z!��0T�Ɩ����������>��)�Q��JR�n􇕒�p��h��]�S�uWDT�6�+UwQ��N�+�E҇�����<��������M� �~|6�m�7y� 7�{�ψ�����|��{�-]��C�R^Kĥ'J�N�+�J�H��(�V�%K)G�����> A�|0����$��3(�x���'��/$A�1�����K  <,��eC�� 	��? <����x}�oL��$�BK�1F�{xj�E$	ˊ���<z0L/bUIRIy'`��R�Q��0˫X��P�$��E(ta o����	��`�����!r�����ߥ�U}Y�}��*J���N�JRuI<%Y7�J^R/E�R@�'�0x ������z���o@O���*����ކ �},�Rʾ��d�ʥU�Tru�b7u��U������y��� �'���oа�X&�U�:�(����Y�R�+*�j��j+s/jd9�6r���f=��{��*^���ĥ$��Y�ʋ��y=��i,R�]ҩ��&RIBV����RA�2��V���V�%�C�|�V��-�}���|�����>ϟ���>�����ڣm���������j�V�-cmڱ��m��m����F�hֶ5�֣m�֨�m�ƫZ*����TmV�-����Q�TX�k�-h���b�ū��X��Ub�5�F�TmkE��E[�m�ձ�j�h�h���Z*�6�Qm�[j�[TmF����m�Vգ[Z*��mEm����cm��hڵ�ذ�"�*� ���"H���b�m�[E�F��kEZ�Z�������@�UdAK�|�}E<�_��7�vr��(�C6V�ޯ%�MU˴��fx��ї癫U�h��G���m �\�C�(HT{<��j� �!ءu@���w��MÐ ��@���̤{���W�$���s�<���^P�/˵̾�;*d*����K���I�pV�W�<��FrQ��)�+]�NM���k�=�_|��{~�!�"�+�I{�`���r�s�B�\ �DI�sv#�	�ۤR��AU��?��x*�*���>�v�?����?Ȳ������?��C�?/��~u֫��n���W�p��_fљwU��ٍ��dH$�K�5T��0muf\��{��gZ޼����Mi{�R�Ob�W�Y䪩ͺX]u*�*S�N�H�����%�\m�u�Y*�����b�&�������*H+e�V㠔n����d���a���<�ɼWy�*V�egz��u���}ь�ñ)K�U�>��͗2�[��Vƨ]�u�qOy߽1��u�;��qG�eP��Vm��m]m�]�u�bָQ��)�t���L��9�fm
'�(]GYZ b��`���Ǣ��\���7�՜��A#Cdy�*�w4���]J�����3s^fm���ڻ���^.�
I��f(�j�ұS�aWV��N�ӵ�΋�q��ͭ��P��r���,4�t�mZ��+{�Nj�%�l*��Z�ݍ�y���pv'rk̫<�!��__f�tB[h��ef��c&��{y�Â�Yi<�tY\/ݮe^dğ
���wwf�bv�+	C`YMGn�M�{�����2��<���`�%��*�1�i	�7�I�c����YB��곷�CE:�U�۬2w�:f>-�&	M��[�kiX$i=%D���[�Wp�+i;ේө��:����̍��(�o QB��WO���њ�V����U�|z�ǎ8�q�t�8��8��8㎜q�q�q�n8�q�q�c�8�8��i�q��qێ8۷q�8�>8�6�8��q�qӎ8��8�:q�|q�m�q���q�q�q�8�<qƜq�qӎ8��8�n8�8��q�q�|||qӧ���8��q��q�|q�qӎ8�n8�8���8�8�=pq�qǽ��w�{�����,5[u.��C+繠���Xsm����l��U�L��U��π ����sm�G�Bw�)]���Q�ZHs�=g�ىM���1�c$����b�\ٝu�mQ�{�*�vw�H�I�np���,=��V�V�ְ��k�;������B���kYSc��xpU�.��ފc*΄���b��z�����z*�sò���!y[$$�]�g�%:鞾�vy�S���Ļ
�u�;�k����{Z�v���cY�;�٧��Z�"�;+�a�z	�Q��\�z�ݏw��VU\'f��r�'r2s��X+���=�O+5�i�e�S{SA�T�o]'۽dq�y*�U,��4؆�Ԗv������a�GYr�Η��k;���Y΢�Q��zh��`ݲs�*��aʻns@�8fa�ږ�G�[̔�ꚺ;�n���soj���3�W��ݛhP��0W`㰩r�y�r�oM���Ff^�Ԯ���U���4�֤Z��$ڷ�V�S.�!��s�|�,Z��s�����t�&��{�ѽ�y����"�}���h�/]���&4�'{SP������Ue�y��.2�]��9��IUМ1p�y2�5˻�m<t��ׯq�z�q�q�q�x�8�8�q��q��q�qێ1�q�q냎8�8�88�8�<qƜq�q�8�N8�;q�q��q�qǮ1�q�v�6�8��8㎜q�q�q�q���q�qǎ8ӎ8�8��t����Ӄ�8�8�\c�8�8��i�q�8�>8�8��8�q��q�qێ<��ŕ�\U�����v��BoF.���S�"���K��x�	E��,�ڵYl!�z�\5Z�9T���@��:vt}}��������Ct1����7i�2n�k�Wr��\�2�9.:f��AREU�o ���t�|9T��f�p�_I��mKܵX�{3jʷ����,���7m��1���z+��uly�ٽ��G�}Zڮ�[*�X8��CV`S+ۺ�����,P7�u���a,�n��g�ųw�z֋��h��dWV[�Tt�j�m��))��p��'yt��esh,�A��|4:��ܠ.����6�wUT�
h^�fX�z�N��dܮ�2����gc�W*�y�C�:n�A���4غk���VU���Um���w���YB�������5:��Ï�5TUY����#g!}(�k��G���^��C�b�VK�Q[c8��0�9ngV]����볆���A�^V^���&&�x���J���Pp�'N�Gv� �[7�ֳWK��M�H*���]f�]��5�7/13�os���aج��<:m�&���wD�c&��$2����j�g�rѬf7xu]S4��yg^��96��"�ROe���XN\��:ܒ6���N<z��8ێ8�;q�8�8�=pq�q�mǮ1�v�;q�q�q��q�N8㍸�8�q�q�qノ8�8�88�8�8�1�q�q냎8�8�88��q��n8�n8�M4�8�N8�8��q�q�pq�q�q뎝:t���q�q�v�q�q�z��8�8���8�8��q�q�x�8����xl�L�m�U{���݄�]w�v����_w��૽q9���T�W*��΀&qV����=��KVW셩��X��f�ƥ���Gp7�R��o	t�8OF���/�u\�-�u卝�G)Q��J�-s���5�<�=�k/�wk��|ɖy��a�9(�>ι�6����wb�U�{�v��Xj�M
���%PAYe����)�&��05��m]6ۗW����s۪G��f�m�e��ȹg'S�5՜�ws��Embޮ��^
,�ޥ�q��2���xZ��V��&�����u��ʳ��ݮ�ԯ��Ѿ�E�| �d�
��c�}77D�W^�3�c�u�_e�JY���}�Lh9Oc�,d�6]־��զγ�מ�ss*+u�l�\��:���YwTo�u�2sW>��Q��^��cs.�RS��!N;�cQ��A�գM����֖Dc���yfO{�l-��X�4\����lʻ��ޫ�m�h(uң��ꮭ[����T�F��ŷ���w`'<nh��=�;n2z*e�i�t�7��^�F^U���7��)��Z܏�,�G'gpԱ�m��fʾ�Y:����X�*1;.�v����w�bf�C�%=ȅ��/w>\}�X�鳘��7��t6��Z��}�[z6�^�&R#���64bLr�ч��iܼ㪆M�uӳG%Em�����u�sܼDq��*��c���:�^�S!���{�"ڒ�W��&UUi������pS�� �!u�0On1Z�64�Z�a��'�#�,�&B/����Mdh+�t���o]��e^T"ƍ�n�42ɉ.;�U���Kz�܁��ؽ��-��IUu���b�R��*�z7�̒]�2����;���L�Gf�/u��	=Z<��ҷ7ye��όb귒�"�C����D�=6̻��Yy�ƬL��[��fN��,���a\j�bŋ�Lڅ]rc�mbM;ݠ�X�D�βDJW;EUĮ�Q�v��-Z6xWnc��q�a�7N�or��M�˱8��h�"����S����,���^���ΰ�aU�`ګ{��ww�3^ͩ���R��S/��Biuڣ%{V���<¹;U�X7�wc�G*���,�s:�Z��.�=yt�8�/O(�7ʝS�o������'��Vۛ���T���̴̼������eVnu-%Ub��U����/5ӻ�6f˪�hX&�b^ Y8i�uEo^o;$�f�w#n��f���ؿgKx���=Vե�M�̖��Xy���1��X���B2�W8rk7���J�|��5U�#l-8*�1- �f���
�s��YV��~$���b�ʶ�8���nțP�2��]��Ȥ7����u�����,��`<���z<=�˕!��M=�´-{j� ��\�z�^�=�)�r��/Wn�@����|�x�K��*ҷWP�=z�0<-XV���	ߴ�s���n2�Rw�l̇r�r����(B��o��/���xy�<��v��sQ���[�QJQuѣ`��vؒu��r��y�7K"�F�u~�@����#��|���:�/:�x���3\���W�h�-��m�%�K�c.h[%J��콿E�)�J�`���tY�:�����	��R��{�p�`Gy�vr�bJ��o���V3�+Sj|Ա���͒��K�\���>���v�ÛT�duUDȫ���ܯ!=oRׁ��Vi� w]»�MjU�y�Օ9S̼ͭʰm#	kVk����W뗹]����]B�r�+lM�y�H�x
��]K�!h�n=�����xh w(��\�Vn��qa7�B�Ç��S�j|�U�m��_u[oj�P�b��t�.B�2��6;�.�Lڔ�D�}�]�f�{-x�#��؁�%��沷YAl��6Y9��tuV����Jʭ��[�)��������t�;ّ�cu��j������k�j����d�fE��Iw��T��k0��\fe�]�wY�u�y5��8�5y���[ՋU�L�$���PV-�ܪ�B��F�N����X�i����Dܻ�Żv�uU�J��t<< Wc($j�g3���т�9�]3�nP8�fh������e��6�v�=��`E h93��|V���,��f��^�lm��S��_�`�WAf{�{�v��G+r�N�m+n��ZipFvtmcڽ ����'n�6�A�x)��i��_V;�;HEh ]�f�4�����vk�jh��{f�ǂ��]i�Vhڑ3G,l���&�T�a�PW7J0%�	Eд�W������-A�[�Z-��m�sj�d�(׼-Ә��#��-_8\��2���a:����^�ţ��8�/2�8Uou�A��Wm�Y��,��ݦ|=�`����z�!M�[}S�A�(!���G���K�����N��#F�G�a�Ý�G%�6���Q�,˾��1:Ѓ7 �a²�Ok��Q��'�SW5\37A�	[�(��R�AY��µQE5�ۭ�y�Gq���<���	3y��+jM�N]]��9-��y�t7�i9B����&�nQ���yi#tX'��~�=��&�i��N��tg^PW��g:�t���\!�Z����5���'�meU�h:�x��vq���e�����V�eU������*P��es��+�wZ��E�����[�^,����%-��Gס�|5�6��ں�g;�=�[�:r�c[������(���б�=D�kUb�{zi���O�ν[颰T��-���/9S�d)�o7V�tP%��CP���N�:��~W|����ܠۙ�������[����6�Bn�ql6WS�����k�sΙRW^���(�h�,�.�UֆrhɩgH������U�s%�B
�!�-_/$(��-��}���zs�l��ˬ��O���
N�n&jV>�N��ѭ�S��v�M�+���6�%�E���/)$��N��wu^eʾXl#��c!,u�c<R��WKR�(V���Xzû�e��i7�yFM�=f�o�L�˥d�����^�j��r���wa�Z3.S��s���]��U]2�яxܵ`��1��uX���\�^�WJ�j��*f^����h�f����c*u��M=7�G%K�s��J�r���6��yTI��Oz�nT�ӫ����Y%�NL[��WWev3Y�zuFb�ו���W^�]ӝ>����y��3�떉�[�<-F�L�њ��6�38�{��)ǈ�-gv���#vK��GL�z�Ҥ7�e�-g
��^�k�>ھb��n�j�q�mcB�6�Y)T�뺩���]��*L�p>D�BG{%k�*��ɔ�k�X˛*匳i�J�P*p��W3�b���i�X�c�.�7e��˹�&G;M*��q,W�XF��&��,N�����-�,6�,�� �wN�o�]�z��0���{s���`��2��_.'��A�=���PK��Ρ`��s�r�ힽ�Uf�Q��.�f�w&b��-�U��7�2�Ȕ����N�� ��[nb�뷰��V�!��׎�GV���^���t�NBf�9%w<y�6���kA)r�����QD!�t�=�N�ڥz���=�z���u��:��X|eH�*����m�er<�*#*���Jig��{��^Q�/���ֳm\jg]���8�&yY8�;jR�f޳ݻ�Ȝ����][mY��Wy�Z��DX�mub>'�yf��n�Y�Og��\Ѧ�,�Pf�!�V����v���{!�2lΗ�*�%Y�����5b��:Wu�g]��LW�Z�z�+���	riB��cCv���՝o{*�]4�^WQʫ��٠��ˊ���ba/i� A�w��<�r�愙�Wn�`N;��ǎ��T�&��9#�-��Йyc��Z���S7g���� �3iC��+]h�/on�*,D�K#n�6bH}�Y�m� �d�n�q+���=u�庅��v��T �=�ȳR��u{��^�.u����'�8�!�������;r7yr�nS)�����ګ���H�Ь���GJw���i�Y��'{���;U��z]�*�kFu+=֮2�om��9z��؊�vB��C3��`��'f4�x�w��!b�e�[�F5㎁�JZ^mm>�H�jþ�$B��Uw+����;�.��r�NZ9���B�5`꣓���A*���;O���j�b<M#�دI�9A4v7U�tyw�n6ѥ4�l�Cʮ�Y2�B�C�N�,�A����Ly��a��0)�/��,5�Q
Q�۳��EE|���v�i��E�d���(>ͬ��k4Ra����)X,�c6CX:�%��Z3S�y��U�s]m�lK�)$�/�5��M���頷gki^+��Bh��m�ۺ�m�삦��v�zk���z�za�!�ۅ� ��ٖ�ɄJ4n�ؤh�Y=���rѽ���78*UF��q�Lh�G����#Z�F��P�CY�:�_�UR��qRDE�M��7��!*�5i���[ݒ��S��3h`P����E��W���u�<��~��@U�Y�����?��%�@������]G������]����(OD�����Cl�,
_�_x�k�<��"B4�jԬ��vB�݈	b�,Q���f�A����l<��7�}�����q3��fv���.v����nL��-�U���)5���fS;M�t2b�;;�.'��K�61[r��,�l �15���um���m�	�����{Kt3�Yo���5,Դ1��&�\�
cZ�k*W�X�{L�1��d�L�یr%��kq@�f��[�n�������fh��6n-bY�q�����#�ң6*�v��^� XJ���fQz�=ib�3.��q)I������&����&�k�J��*���$a1���Ԑ�t�c�pՓ)G1��h�4LK��7�
i�L;�9���rk �v�W�x��⦳jA�1� K�1@��Rh6Ū�]X�7l�54��J0�-�,�!�qyЌ�S���nĺmq^n.Z�����j�U�c&m��#kh�vW�+f�U9�&�L�	��͑٦�cRW3W�n��j�3�K1SQ��1�c#�B�&l̶cbn,�R��nnu%u�c)��rmA�2d��K��p�U�4"�ز�#e�&��ƃ0E�L�m%��i�S b\�@��#6��m�� �-c�CkmV,�f&�i��E�&6͙��J��c�̫jD�:��fc2n��WZ.�^۝��K�rL[�����o5��g���LdZ3l�6�ҭz�l���e�X京ư�nmB�B�`�h�"
��t0�.��1A�i���aţ��v�!��؎�0ح��a�\P����V�8֫��YA\�'�9��5h���h۔jB�����Л:�ocf	�]nH@����c�ţ�(
+�e#+s�k����i��B݆6nn�H6�.8G��4�ɦ����@��v��m&���H́Y[���%�8�(\�.�R�&�npKu�pK`,\�S6VĘË���P�Wl5��J2�Ѕ�)�4XR���TH.���לL^�#�.�1�mfóh��vt�,P؃r``V-����U��J:K�4��l�\B�P�.4&�WJ�uא��^܈4m�V�cC;��n�16��]���(�*�^٪af��J��f᤯7�{X���y�Rn2�܊��&�ÓLA��]�%hL��m�$[i%À���f�֎�IvLF��jB�p�ՙ�i%P���v����ԚR��G4���D��:�B�m`ZE�Й�U�(��6V�b �e��4����f�gQvҺ��`����Κn�<�1(�ҙ�.K%�&
fښ��50Z����:ǵ�Z��!Q�#�K�fـ�b��f����.��f��6���x���غ
�vQ7�4��GmɃM*b&�b���	���U��Jd���ZY2͝k*4t�\85��q�Ћ�3��L����5elH�J9�J��n�B)*cÀ.�J�1WD����o�ޥf2�5�sU�R������^tR��oD��[��at6�0�Q���	��5�n��1P���JK6���b��h�����Z-V�����H2��H��L����r�7l]�U�&$e��CVf��V���CisA�����%��������\*̶ِZ�6�4�F�(�n��G �[��a�-���Һkm���8˅% �VV�{2�YR�{(XJ�]��ʉAM�hsM�V�7�^�]��P�-���fUЈcL�ݛ!lp������:l�5L�D	��6kݻ쐲���B�,q������^�m�u�R��s���jǉX��n��n&�u���6��ڌtK��J�W62����v-�R`aUYa��kZ�eQT\@��J�lM��җ& :-�M#��`���é��B�LR�6���v��	)7b�L������b��E��Ř�lU��1��c!�����^�Y�e�H�D�vݪ�iL�1E�����5�z�J�s�!��:h%�&�0�.©��6�bc4�p�#
=ZGV�.�gM���72�ٛ���ǘ[��6�����
)1�l]3�-!�,oQndYJ�0���1��4���GTw`�h�DC�'�x��j1JE�V��X<�b:Zq.��-!�LۑʩXhB�a�1��	i�/,���i޹�%�M�6�L4�tHn-�
�Fq�F\�m�n\XFhи��R죑j˚@6!k����cE��e�ie��F��pƤ��N�����5��΁�7JLW6RFYjhƼ���tBV;h2�vq1F�u���f���5�;�*�Le-��y�0�-�"��)7i�VF[�m�6\Q"ًu�k(�V�%�*-q1������a�!l�`6�k�T�Zm��B���7l�kc�dp`.b��R:���� ���iu�@��u��*]�h�@m&��v��!K���̦b3K��f����i�`ZK(�Ý3�����%�!lpuB�Fےpbʨi��Y�vaqu׮��;f��e�r"��Y]�C=fq)aHā�I�m�����(^J ��˝p�R�B�-�!	i�0Ѕ��ķvф���[��l�JVkl��.�ї.��0%�2.(�m�Kn���!h�1]���k��D5��$Mz��-,)xf���k��╘M�15"���GRP���L_��{��%��c�&�S�M[,�XuE�6ܷ$��jڱ�L��mr9�]j|p����sn�[fIV�RWk���tV��9���P��Zn�������+�%&�k*���R����y��u�����j8�*حV�.{_�`e��ka&.�Z������6�&�Va�.]�<�ږ*���h,��&�4�t5�4�����-���V�iJX�`Q�K�e�dD1"���j����9�%�^,ٸ3ê�tؗLƍԆTp�AЮ�5,�d�ZY
*�%Ѳ��](�ַ����\r]l7ko��&In�ϼ��7Hͬ�HR8��Ɩf:�6���k<y�-j\M������	n4��\`�haZ.��qI�.aͰZ�p�K����"�53�c�Gu��kyISr*�B&�-w���V���s
b�,�Qа$�vͲ�bׂfS+D�b�ĀWM���ĺ��14݉�{$C��Y�����u��[���f30 �.�"�#�kj���ʄ(���q�Fb�\��)��ܶ]++��re[]V���M��Q̰���M.!��YP�r�v6���\�!k�-Ձ�,k��f���"�%z�6+D�;-r�ݸbWSXҰ�H<�d�1V7dp�ٱ 2ͥ�Y�L�ڳ9��3�X&��1lq������b\͔��ư� 1K]��e�r�iME��7X�1�49�)n�K��Ħ�%K0����04K�76^F�Y�*WnL�ي������Д�[l�Ya*���T�j�қMe�4�+��	!�[G$���l��]6Ԧ��kg-Y�K��u��A�b�%�P{e�]�5
�+�]-����M+��!����8�٨�LG9���R�X8!�V3�$,i�Q���!,ԛ+���uj�0]����f������ţB�VY�R7Zln�n@lr:�kJ�e0Y�6eΰ����R�)3rs�Z8&��u\R�b�U�B����v�&k%-.��^����ˆ53�C����������kX�lr؋���M�Vʭ
���,tMl7���D14�6.,��̻icU6��ؑG�BSb�隖\FeB���J��j��̀�&Mr�.h�[Q�Uu�h�"��X �4U�6�ф-�˩m��E�������taqC�E�48���:\67�KKLKi��\�98%�7��v�6ʮ�#�`��l!��&Ee�g.J̈���ֻ]��ɍ�PYZ����@�;X�1�7HXhZ�e�i��uV۪:P�6ie�Vr�\�<���*Q��͘��w
 ���� X�c%@�!f�t�Mt�g0��ل2�p#{qtUƄ�����r�!�i4V��� vm��u�f�h��.E�Z�q�]�YX���l3�F-�
�#H^a,[f�q�Tfţ1�T/=�[1@,�����v�ަ�f�-!�*!�J�.t�C2⺊�
��h�e�����kK(��,��q�)B��ȴ���Ĺ��y�}�T�1���!�pF�[ �2�cmA��mT+)(F�Kql���G$f���X�Mt�Rݐ	�W����{�ˢ��V��i�`�Sla�ekD��5-X�(��޹��A�V՘�%\H�.r4v����J�wU�d1��9���˵�H��ܲ�:*�8�!W6;�
@��F-�a�2�M+e�#	�6�WCG8�p�2�.e,�k���alԈ@�HT6`ʘ��ڄu����.ؤ$%�o*k)
#��MtZsé�3�Օ���3�
����UUUUUU
�-]�B5�5��,3�21b%s�%�[hK-������!�m=�k�%��2�#.�^���b^H�m<7�Lx����Hԥ�w���0�A٥�%�0���@땅ш��й׵5�CBYY�&2l�j�TT��R�M-��b�X:��G[[K�m��b�eU��2����=I����<�5_bu؆������Fh]6��3�.�i�A��)L��k����q��|��i�1͘%�136%M�l��B仐�v�!1� �hPM+i6�fȗF �X�]yMsWgR�.����	�m�h�m
\�E�2؏�����:��u�׉X`ʗ�����e� ���ٮ�E���<�@���u9��8�)��9���)^�Ȳ�����
���y<��,|�]{SX5Ƙ�(u�R兮��;6�T�Xk���FLjQ9�[�@��'���B�'����tX �:�sH��j�)v-q�4%��MH��B��9Yn��n��W@��kc�͛q�G[f�`�p;  5|6��=:Ź��b����d������v�v��q�z����4�ӧZ� �YA#}+�1�$��(����t�8�8�=z���M:޷��֊6Ɛ�DhS"�!5K�%�qӷN��8�8�ׯ_tӧN�jH�H�H��
�b���]���s�+s&�Ӵ��ź��T9rN�C�wwurf���uӸ��\��h��˻[rH�u�ŴHVЈ"��D�$�R�s���mQ�	mR��wm��;�m��+Ǟݹ���a��╳9F�����mMp�T��Z��.�;��B�l�}��<MrUݓw6�/���≮]���o8�wg!͍�^&ܨۥ�Z��ou�k��7M�ʹlkDm��Rܢ�`-�r���jꭾ>|5���Q1n��L���^�������c���[�M��؏��|~_���
1�
�kw�:_zx���w���ыƘ��M+�$��Bd��`K����2�nq-#D�h[�Mr�(V�eu�J����q���a�5N���� �Z˭�f6���B0�u����������b���/37ZX��*����涚k
��� �m�I�4Ա�e\D��]��0�]���ً�L�֓ 6����hIK��v2�H�ĨV�J].��l6��瘱��u�WdjXi`L�
M�m��niq+�.�o1�%-48��YsɡŹu�!`n�HiF9�bܘ�9
kx��H�٢�"L5J�yr���|��-�+84+1�s-�"�p�-0Qe�Wk\�.�n@@H���[ni��#B*�)vm��0%��1�q�'U �!3�B�:��
V"]�Ҥ%���b�cP��Zffd25-�HЋ1n�	JCZ�#vu�]�B�sC �hPm��5	��Y[S���1�a�P��T%�90�"�՘��W,���]�x����A0TqSjї0��]n��ku�[��/ ,
.\-�#�r��m��|g�ɖ��X��m�Dv�F[0�!�,�+�ԯ��d��;h�*����k��4�u�d;E�[3�H���Pݴ4
�5\ۭi�r�d4&Г4�ʻ9n,lM��츶(踫��hk��L�x��aȀ��0�[4ca���l4���`l���ADn�D�\�8���8m�G8����+��2;$�x�����^��!�5��{s�2(�q+��!�6K�ؙf�$5�B��k�R�i��3BE��E�h$b��,��tJ�BP��h�h��*����ue�3U�f�yYe	K\:�������r][�n��	IKX�Z��Jc:��Zd:���!�ٶ�����KB\h�1F�%�V�\k�A���$�h
���]3,@,Y� 3t������=�#+ޅ5;�g�*�y�*�i��,(�qԱ��ǘZJ�YAy��`�b�$K��`JaP��匤lahJ��
Z�- � �RX�Yb��[C���ZJ�QV��-Vk�	������A��F ��N
�k���eQ��Q��4�,��\h#�%%@_|���}��Ϛk~~lF��LP�� ����c ���U��u��sY��F�}��c�I��S�N��O_p�y�MMm� 3f�w�ken��y��	(7A����gt/ۻC2�[&Y7[8�k٧"bNbj}|N�N�bǓ�\C=x���$���߻�~Y��)v<�l���X1\{r*��%��h�x�8�MT��Be ���O�fc]���lL���VM���MVݡm ̵6<�M3���J����̯��C%�Y������K�R��Lg�"ҪL&FP/r}��~�>~�m�Ŷ�Kv�9F*�tf]��r��n��̈O��!��2���R�l�V�,��;��,9����^Z��g��N�"At�oǢ�t�>�/(����D�M�ڸg�K6g����%@�γc���Ϊͤ���e�����
*�:�G,�oFn#T�)I��T�����b<�ŋfbŐb!��U�/Nc�^M��^NV�ݿ��&���)SN%+�$��W����)�!�	;/>?}3�m�tK~}��$���+ b}�]��������N�t��0������C���)�U!2���{�cP.l��|�X+�tR�s�:.��I�U����|������p�W��{4|�#e<pÒ/\��wXE�m`��]/]�К��Tn��l'T�j=�7�n��h}3���{�y���|8�����6y�n�y��+g��x�������������'t����P�v#a93��|�V}�����gϨ'^m<�W�6�� �#b�3Uu������珵���"+���α�Z5��͉�_T���â
����l������M�nsf{8�1�`���]ܤ�f��}��Qᝨs�T�v;n���ګJ�.�_�>��� +�f����g�s�{s�g�;�'��%'�pޠ�y���z}�o��mj�ߵ����}���`B�L�3P��L�m*�P]�DAw	-̦��M3.M�J�&,�u4F�ʫz��XW#|}����V�5H L�}�J���H��Yl����u�� "�y���h'@1//χ�\�qBc+ג�3u)��N*�#iəW��O���� 7`�� U!%I�`�����I_Dw>��9���v��}��L��0Ϸ{�|�9�z��(�'Վ��Jg>���,}��������ｃ �q��Ĳ�I�m����Ѧ�Ui��g�݃ADmM7�-/b��z�\;��g�܈kջ� 8�@O����S��05�w�M�a��m&ּz=v��1��*��7N��FN*��֠�U&���c_e��j��_Ly� 5�3M�B�cK��Zh8�P�I��s��X&-պ�w��L���[i�^mQ���[~��]�րEQ���a}{��U-FeӴN/@����!��}�&�����av��	�O�ժ]��1'���!2�^��a��\9_x�����7��D��&�Bej�}���{u���{P�W���^��]�ֆ8��Rڃ~9����2��X��fwge�KB�g����FG��o�fNݩl�N�W{�z"�S�eޯ{�:�j&�)ef}�����w��n�qՄ��݇bvlT�u$�����k��(��Ys2[�vQs�9�#�jŇ�L�ĘE�ɋ �z�8�ɿ;�a���ey4��
��j1�rL��B
FX�d��
���uֵ���܈��3<9biL���]� W�t,� �3[�1�LD�3r@qLjK��q[����ʘ)�.�� ����1̛U0��j鶆n��%��L���Pp�:�J0�jb`��Q�vI�1khmyƲͣV�ݣ�ς�	<���<�}ڰ%�v�]rW31�h��Բ�����U~4u�hYt��+a�����-��F!<DA
��x����@U!2��ʟ7���|^.��E�E�߸.�X^�#��S�M��W�3�C`f��v��{�ѹ�N��>�ـ���ߛ�nٯ��b��ye���7^yA��g3�s��a �c��`終����;��؞�zJ�͍���ݦ��;/����s��_|����w�ީ����@]c喙׼�^.X�R8�t��OF2��ۏ��fGכ}����u�oI���\�	�������/e����ku��nc���f���S�4�z�JV>�>�x�<�T����y�p�Ӟr�fd��W����etm�Z@L�ĺ:���&V�D���������s{'ת�|c�z1�M�U{�W3ll����2�U>�.�a����]s*>� ��+�|��+=�3~{�==��s��eWx�Ssh�w5e_�fL���4�/�}�)��y�Q�UB��os���޽�w���*��6��Y�mXܣSw�]Si������X�ت����E���&���h5���&��``��r��ϧ%����G����}~ ��M׃d|����?U-H7t	P)n� ��[�0\͘��n��՚���
�[��=$�����92}�}�ܶ5��r�K���������6݆����d��R������[������FRb�[u��l�U�������eCI�U����v���)�ժ jc>�V���w{�2�����L�i�����f�B��5-�CB�^<{�lڞ_m�����潲ӬČ<�ݏlnM�?��)=�Be0�A65TVH*���
T��x�T)��3rw�}|��ELsC]�NtMG��˴��Y�6����pe	�0����Z���U듵�C�{5�P�@L��${�x�S��cD�65���,�oe�z��\�]D5�0��
ABe�_|��5�;�����w��or}��I�y��ξ�:|�mV}Y��K~@���E��ō��Uh[K2����T^���֙@`�*P����f�ն6�7��.�����eY�n��B�6�Z(Q���yr^v��~�f�̐'[�H&�uJ��۪�9Of8P�u/o�o~���+����;p|8ťC�f�X��ţU�6,����s]q�ba�ѽu���>���	��J���t̺����m��y����L��n�����{�{�7��s�
'a�"}rf���5e��=(���$�����f�#��}E!~�8ڵ]�4�.�e����ƶG��������;A<��޳�P	�bg�c&��4_��P���yҏ
��o�-���e0��)�Z׽i���g�n��Z&%e�b�+ M2��G�͵�C��>��5R�@������ζ��>}s�VY�ڇ���מכ��ϐCk:�*O�� '�	�;Q��LʵsZ�<�.stE�x�@O����;(gPm���t��n8K�^��>�ٯ��倩��׳����}�9�)����e�zB�y�zzF�x�utA Š�gim���n��'c�oh��\�n+N#9\�Y���h���D�T�B0#���XI��o޿/��-�ܣ>ߪJ��p%��.i���P	H�K��� L-��oV��͎e�9ut��Q5Jn��4S�9���#�10m�v�M���L�B!l蹥H���+.ٺ�\lS�
�Ae+.��K�]a��y�)�����uk�^�i��`d[u�8�XU�RnP�abY�W/^�t�Z��x��VY���W<�Wv��`�EA�Y�?91$���&��iaX)f�H�f+[\T�EM�*�J�Q���UY?gխ���jgצ�ړ�%�E���Z��Je7���mϜ���&����\?YO���K�z����<�)9�Y��_��L���(4���cn�W��$�ۍ����7w�§�M���>n���G����%m��%{P�U�b�7ٖT�r�>��:�'���ܺ���g���{��;�1�343)�fr�E1�Ȇ���C(��7p�9@�K�tQ�4�te�Ჵ�T��ˊݦ5���r,v��&9�m�߫��7B�g�;n��wz�y�ٸU�wҽ2�Su��|D����ϯp��;�sr��Y��-fm�I��TV�2P��lh�x�ݸ�2�Rh*wS��ՉX�W�/����2���-���� ��X�0X��.E�Q��:��EI4zPj�z\�ǟnW��$��+�&�v�x0mL��Zf�D�u5�mNxY�/Ɇbff$	p��s�}�bzՂ$ى�@}�B�tsm|>wn󯤠�>�9O}����u��oyڒع`�d�� ��¦Ms>��]���m�$����;���@�լ�Qʉ|����6�7m�h\�T�������h͉��c���\[ڛ!L����+DK�����ѷ"7LV\��]��%hf�q�F��Ru�g�����s�Fe^K�HcYdfŪ��$N�w��c�s�y�(A�k���B����Ą#f}�GRP�U�ǁe��peǖ����)aV�Q
�֓P���t0�ܺ�s��U�V���A��t;��xfTa��5yR��>S�ٌW��m*��x]�Ӄ��s������ޗ5��f��f����F`���u�pi�Kv���f�5�N��M�'UBMJ�^�7's<9Sa�2j�LW}QvB�N��{���j*�h����B����\�s�]��N��\��uQF�G&뙹/[��F��n�)Q��*ٹio]u���V�s�o�a��G��}��geF\��k.�Y|�k5x�fѐ��"�7�>�禰*��"�� ʾ�n�P��/]��yy����e��v�Xvh�t���.���kdP<�ަ΂U�[�b��v+��W�GH��{{��ɹ�E������eƬP�N�uwX{n^V��Nb�Y}qg�"�t3e��ެuO_V ���BlX�SØt�US��"��	e�Ws�N�aq^����I��s�i�;ޝr-'"/�iw|gN���|��3���V$v�YՄ���'pZz�剹�F\iW��b�jܿv���gY�̺2�3IS���XDӋf)��X�`�F�̽�͉_j�7F�&aY[�s��Z��E�L���v<C���wz�{)Q
�UGX�xl$�p�G��dVW�����%W��YP-P�#�����P��b����]
u^��B.�Xu��"-"u-]�?�>����r]Q*��<��ʊH�@
��##!# 2H��ӷ�N����8�׏>���m��m;�)U�ʧw5�����Aj6$!���׎�1�����z������n�v�����2! �I H�eI�d���O�;x��������ׯ>���v۷n�@�Z+5DZ������5�+F�b+Ƃث�nZ��k��Eo��TF�l[_k\��1��lTV�j��4Zѭ"�#�n7	cME|��-���M44��Oo��wWVg=+wS��x�^��#WA�&g�ÃT��
��32�t����n1�aI	2�z��c��᪓8{���b_G��/ge��,�������x57;����"O2�6�w��Fw�Y}��9G�y�B�6|u�0�7T�'�=�}���ʼ��`.�p7�Ro�h�^$�����"3C
�h���0РY�g1 �	�G<����	�Xkh��
�Õxi�7
�{^g�`yYo�3����Nc����� A�B�w�*{~�x
j���2�Oe�s�aU�pA�D��ѵ�g�i�3�Xe��!kHp����D�w^�n-q&YJ5Qj�O�I�fa�U��Ӥ7�u�E��9�E��4awˤ�Ր�  ��78$���c��23*�d�5G���'���il9�l�'#�P��G����� hb�HV�� ��I¼��/������ l��~|�o����s+;qܫ��(I��i���ݼ�%����U��v��=y|zȉ���N�p���d{�D�(1�#�DyA��d&r��	���C��}7��ff����X��u��O�ctZ�t�-���+ �t�n���Y��(������n�m��#^��5�#2\#H<:��V�i@&�׈���]ނo��H( A�nز�+��ݻ�{��y���Fe^rTppko���K��@�5��h�'��c��K��*��&�9aB.�w��������:r����wZ=7��/���2`Xܠ��zṭY���,�H��f�\8#�ð ���T��]�q��0��s���R�� gp�]���T<�a�e>�h;��4�}��|����z�Y�nk���9��0v����Ʊ��	 ݸvf��;u�Fg�9�j4x�voeb�>B�p�h� �&rRlkVC]�Ò�Wj�����R�q^�zkxo�/��sY C�1Z�͖�v�������
{�n	��P��)��Fy�5#ׄѥ�[�p��{�{]�$T��¤���ߢ�۞��;�U����:`e�����c ���s7�k�yZ���'�ֿf�'�����][�q{muƃ#���4�̺�!���c2�J�Z3EA�Ѭ
���!��k,y��*-r��6�4�\(�S�D�(٫f���L�R�XJ�Ԛ��Vˍ��� uؖ
d�g0�K�fj� ��a0��U,%�*��:�]vtl����.�Bd��)Y*�J���Z�#�����ox�LZ�[�c��[�s^lu�X�?���mj�� ��.e�F ���s�]mKu˂��*��k�>�ό!y$�;��v����K���x�>��1ى{���0�z-#�/�qP���VB�ڲ\��Rq�sT�f�6�^�����&�%�����[�(dfgc�s,8@�g8r]�Z×�y����x�Z���gj�gh^���',5J|,j�DZ�`6�Ђ$��kz{�|���@�9�Lϭ��ْ�v�����V!U��m0�����(MG��������W+������2����v%ݔ�	� ���'��:}6���7jτ1
����P��=u�b��, vL�8z{��<���������f�^�j�4�#c�O�<�{��炷l�%5�M�v�oe�mAf���Y��	�,�
�ٵh"����[\G����������Uy㻱:��[>W�UH�s��v���艠u�0���q ���i�D���*����.��9�\f5���
Ǯ��5s�,*�%O��bp�lm�q�rέ�>����K�P����c?����ú�9�/n�>���ģ;-p ��c�9��@�T=Si(�	h�f�N�6۸'v��%�ő% �#�c�DËo��լ/L�w��"��=+�ֹ̼L8�����*vp©<�n
ۑc�ϖ����|�;��X�t ������*�9�8;m��(?
��!j׾��9�^sVB�\Nr��=숼�3��ڱ�����ģ;-s;&v���(y��am��A1�R��H*�|���y�����( �K�\�
��F��j�F�e�LVWQ�ղ��Z>��:~�ߤA�˖ 8"��ک�8Q�fx�A|���FRS�:z���5j���A��v�7hA�9�8@����i7�,0�A�V�������ۇ�F�J�lt%b[�M*�dK��3
��|��/<�-80��v�ńy�ص*"�z�@��S��r���6���/i�v�:w�P�Y�UY�;��r��1�ai=�Ǌ�ʼxS5/��&}Ts�m	�,C,X�#�L����hQ�߱(��|�Ovq!�����;uq>1��Ogt�O��k��A~��fh8�Al�<t�K]��^��ǰD���X()�`@6|\c�3wq�����:L4��gLi�!��1l�(Y�!�Š7ƌ�X�t���iUGtv9�N���z 9� �"ŀv�p�j�5R	2(�9��}�&�J�Gq[����i]\Q%.��7P�R�j�5Z#�`�a�z�pA���k�gcv�{2֭=]�^�. ���lW�ь��t ��{� �&J^>R��C���̭3|sC�L����B����#��y�E���d���+��؊���;/?N��@�� ����@����A��dz���؉����P)yO��cg���i�>.b��-�᪐��`�ER�&��`�����cz��v+ѣ+�����-m�pؠz�b*��a�k�L)��lg����1��:�F�ݿ��@2��z��z��q�Z�d�Mel�U�v*���*�X�Y]��)�9!�$�>�cQ�5P���E$BE���=�g���!󴜜��Bd��!������{uL��4��x`~��՝��1z�6A�&y�ܠ��A_��"x�8���C3I�����>���%(���i�
B� ��-���2�Zb��o�6�jpXn&sT��'��;Q��"���WM�nέ�����sU��{��Â©�g	�RX=D��W���6�� ���I�����;�h���^�p��Łn�J��h���bi�YwOL�n� �~L�*�5Rhc�a9]�}b�
�I�հ�=ܝF/U�y��� x[�SB��P9�=fٮ����J�U֒��m��r	�@;����kP���,\Xr�9U,�a�o�9aU�"�\,A����ۇ"�6��;�޶X���vq��s��Ay����q�)���m����CU.ٌ��Q��ބ�O$Z��j�X����a�u��v<��vo�dZ�m�[��+,t)&(���tS�vԤ��Z�(4��v9` � {�i�TT��4�BD)�4%�1  ���9Nc2Tǽ/݂��QO~��}�y���� F[,�%�����[A�j����K�\�6��cuv�m�m�!bڐ]͵k3�\���7��O��<�5��D�vs�+J�%k�ʀ0a�U[,V4͕d�q�ʄ�����V8��o�wi�B��!�,��ښb��K�j��QI��i5R��]n� i)�
.�'t�D�^@����fo]��j�̾�z�;R�W܊6�V���A(��y	8�X�iR4E��J����a��ݡiP8�[.�B璪�In��_`�f��G�Yi�����u.���^1�o;���s8��TO�X4<ðv�PZ����7h�A��J�^$�����(	��4�b����z�b�9i��c����Q�g9�7�)os�F�H80Ʃ 9�c;]�c{ef�=�O�=�k ��a��Q�Pq<.��K��X��|�[U���T� ��@9�(U.�E�/��Π�D��GL(��U)c�=���;�Q�3y͑��FˑK��B��\uV��a�E�;CQ��H7��'�Y�d���{��h�!�n��d}䣬m��:�F�^�s�0 �c Fc�yVl�,"�=J���e�G�{��blY����2�j��dms��.���F��]Q!T&�)�+v6\C �jІl�B�1Ņ����<���q����o��֓�;�m�2�ٚ���<��I'9@z��H���<1��oس_]i���������"4D�/�Gy�bJ�n�CGb�$U��������t�ںܯC~&��"?M1�Z��H��Uj Ȩ�X
%!wI�J��A��t����;�wʉ�����	�e�"����U{�sޝ���Y�ce� @� L���|J^>����N�����f.V��b7��#�l��m�a ٲ�E۰�"�]�ުV�ї*�(�"-md�S�)Q`�c�V�"xM����s ��@9`������� ����@y��N�
��T�4mo� �����c0-�����*�/{�YY͏�	N �;"�ݨ�a�z���J޻z�#��|�����W-�����n�;U�.8��r�ihj;r� #SD��X%6Ӂa��U&pRvh��>��
�^�s�w��C���k9iהu��r�!�p�m.rﬨ��C/�y�3)u��=���d�+sA�]e�ub�X�L�Xy�A	�� �f��,n�3q;4� �&"��:eF�S���{��o�ݵWl�T� ГM������0�osʗ��n�d_�l�Q��@����p>:i�VГ����p̪4�e��$��U_@/ӌhQ�1���4ƑU*"$��*!�I'�����)�"k5��g�FːZ-�9N��P�J�J��dt<���x�D�y��t�>�W���9��A�����_���L!�-Á���`A�d44]��,.n}C����x"���b<Y`�/�8�]7O\��n|��9�찀nӐ�k�1��&�g4��
t�
%�Hi��M��gC;.�X̛gk�d��Mza�A��8 C�j�k2@��;ط*���1�5�	���af���l)=��y9�9��N�M�Þ������ѩ�1k����Յ�=����v�>�W��;�q��N&g�v�d
��m8��\�߱�UyÖ���x�qT�ذ�wcJ���ȩ�]uS�Xh���ꢸ>�����|TAgL�IĲ�.ơ �E!.�d�c�X� �]���E� U;�6�S�įC��l�288 �fˑ}��gqml�1#��=5F�P�M�߾u���{��ќ�R�ܑvot��+]l�}��q�[ck7�|ֵ�:y����6Ɣ��+mۭ�tը�j,�Mj�dQP)����7l�_TP�/1T��2��pj���g>𽣬1�a3=���y���(��b�8 �Y@!�2=*�����Ý�Þ/����Ji��$��0��Ъ��6(�f��Q�L8��u���$�&�,�<�Ap̢�s�[	�Q{,���=ou��pK��5*�u�0t��5�� ]� ������j�aױ�L.�L3�4��NAm�`��o�{������vj��3��V�Co&�
{)��s؃�K�\���N��<�uT���]�<�A�tR~]^}�z.Ɔ{�kS3����2D��"Hf��;�)�����9a{�Dv�����޻��	�2�M� ��=�rλ�y�[�'W�T������ �@m �\���vف�ȗ����y�{����L8����h�m��ld�(��R�y��kN�a����s6��Bz�\��yG���Ŝ����v�6�GK����锫\�n����y�8r��M��������+!Ƅ꾊�v`��&��B
\�����+�sK�:TC���cvu�Iֶ�z�M㴍��[jK��^�d���30���YX��r��[�wW�6�]��y����%[n��]n�8��ů��md�j�f�ƒ�G��������V�V��E�B�����鵵�\���-��z������ъiz9���w�W`��u���R] ��&�T�������y�hP��ܦsR=�𫗗�cz�T��h۽ً-4G-�#�fg%����[-V��V[}�ɛ���sg�;9�����M̌�7{{��L���s4���4���us�5��їu{�/.���W�Ӥhavw=�R�ua���2ҥi�ոh�K.C�c�7�9S
wt���3���m$JTyKhwf�p�:�]i�ؠ�t�VPH;�{ L���f�C\�1�+3F�r���&{Lt*�T����2����a�����9ʕ��n��]����2����}Y�Ζ�o��9xi�,7�N�1F�:C�ʽ�֫:��m�a畛��s����q��#���8eҮ��f[w�f�+�|�!�EH�Y�d�Դ+��em�ʷM���ǆ���p����w{qPRޭxy��]��U%U����8����!�ˏ/6�We��,�@�� 8̡d%D�
Z�<����|��Т���������H2) �m�];x�n>��������_]�v��Ө�����"�Ƣ�U����ӧn4㏯����8�����nݾ;t��"H�2�����;q��q�_\qǮ�_]�v��҆��v5B@����)"a�B��@*\U�j
v�`�ME��nyZכY��r�嶊�(��U��������*�j�����)S^�ײ<gW���҆�g�ս�<Cv�[mFi��i�ɸ��Ch�����v� �����V7�"��e`e�)I��\b�����c�]/.Fb#4d�L�4�\(L�IVg00YA0�ccZ�׭�s�G�C�.J3�J�r����lŖhѢ�l­L.�i�7&�ˑ���K�F�f���� ��swVX7$�rY�p;)aM;E�.�����w9V	��APٔ��X�E���.���Ox���gjl�6t+(�qq*B[Џg#4ZADr����֊[�nme�H��;9����}��.s��L��9,�WlX�.K4�U�7�"��-�hRTu��jK-Ъ��.Z��7d�,�4����3�E`�L%T�[���=�1]�Ye/ie�ˡ.sψ>M��X��j0Kr+y��2��X����tID��4)����&R��.�+�`pM,�"R��m@���lj`��c�l�G�� 1�u��Y��e��V��(/m�4(���3��D֚mi�4�AF�v�r��"G`��X�7b�f�	t�°܍�s4��	Q�ZF��a�[���4��iwc ��*hU�&������
��"��i�h-���b�к�u/�T���hֲ�ۮHGl`$.wW7M�Pl%��l.�b��4�f�d��(M6�n�:�Shg[5{7$yb;��h\L"땔08P��4w2�i���̈́n+��qYK5Q6�,LC#�./]46#�*�V҄��Ʋ�Q٩f⍚�+n��H�䆺W Þ����}��p!�I��L6�����@T$�vfe���LV.�fiJ��.̶�Y��P1����{]�CK�kc	�v� 0��XX��<ڦ��	�й��1�R�Klb��������0��[���c�]�Px���\)Z�-�RL��<��k��ݥ��	z�	u�K6c�R�E��SmD)&�����	�T Vk�X�їL�%X�#�L`j�.���U�p�����D���B�j�(�*����׷�7����D�����_� ����z��Nn����	Kr�ܙ�v�ʥ�PS�cn����i��1�xיp@��fqoYb次6�+���u6LX�����4D���.X)75�!s5 �meJ�ji���A�slme��0m�ٳ�9��%��x;bR���LGL�5e���nl��c��X�إ˾�}|7���~~O��WM�(�ӟ��f��A�(bʩ��i7!�V��f�ۭ�&Y]�c.%��=���=xte^Pn��K��Ro1����u/��/��*�`kX�Au�HP0��0�.� ������P�����x�;Ja88�-ܥ�=���+�'@�\Ac~L�HsJ�R�A\D>U�f �j8[�Aq3U&�Rʀ s�⦖v���e�����I"	]q:�9�����z��|������Ռ9\�d�*����4B@YJ�8�r	�O}<+�}/�|/��F�obX+�TtdC"-���M�K"G5e�r�$��SS�pEUj���D������b�W.�*t���y �&X�C���uhf �v��I��1l����9П���	���Ђ83���k@�%l�a`v��¶|�=�K=��r��A����RyՋ������.�����S���Y�ʲ§PqX-L�� �KŪ��!�n�+O��$��ae5�����Fz�ayP>�h���y]�����L7���K�[�mqv{:K[n�y[��F��^P�
5?CB#M#B1cCH�Q A
C���>���=k����}���i��&� �䘹`v�8U-�/�:rl�B2����ES�,*���B#�B7@�`ŗC��񱒮��'��\�s� �}ARP �^����?:S쿗s��6$vm��S�/�Z;ox�?���g�A�p!Rl�S+k��a�d�v �j��eR@9��� ������#9�u6i8s�͙���N��V����͆k��7+s�'h+�}����B�!����6�̺�2����6�aRa5#IQ��˟���0��a� �Q��*!ڣs-t��	7u�C�.L�S3�wʁ`uYR�{Y0�p]�c ���]�t�]_���A`Z�ۭ���W��͠FB,@�l�pA�vEݦ�3���[Õƭ9�',(�j���C�i˕�NH�'�zCݪ�o�[[8m��"���v,�L��l�n﮷����찋���7�Ze-�����򞈌����@?  Y�@c�4�44 ��Ң�C33�9O|=��g�_�
��O҂>yd���������ay +k*$�6�3\��XR��ES�c{�[��.��l�1��r<�6�L#g�֮���LA3��)�&H@��.�=��(r�=�5w�f�.�>�U�*�:	�	1
��t������w�����v��n�9Y]��[d�k-%1�įm��P��8X�N�.b	�' ���k<�5I؂j�������>�</���d?�2�v �k��bS��B�7h
̺Z��
v��oF;:��'w�����C�a��LuӐF۳����ڮ*�ѷ��MX��R�ک1���f��٬�u�7H�X�̨��gފ��/�d	�ѷ½ew,�f[��2�<Ɓ����Y���SP31h"=9�ɝN��`
�ulp�͝�g��T��c��#<�g��DP������)�=�ZVݵ������j����e��H��3�|k9���p/����]u�zP�V�RO�]�D�@��Њ�����5VDQd ~N>9h8 ��K!I� 骠@"�|��|c�a�ԛ��lb�*��_��p9(3�� T/ Z�V�#�;�nlʿ ,�C`cSb��J�Bk�t^J��6���Q�ԕ�,' ���G2e��pEr��@N�;��z#�Ͻ����h��r�6n��)\X�@`�p7e��S�?2�P]�Q��x��}2ޝi5%�g3����ћ;E���7��{��C�[�0.A3�@��D�'�;��vɠx�+)���Y�[�D�T�����A�q&�' ���!v����Ӂ��]���n���8y��u�1æW�3��fPr�s3\�e����a��l;��9ʶS(�\�y�u9��ADH ̪ޫ��ٜ�f�k��	����\�8 H�{�g���'.�㉏ݓ9�v*�6�
�l��A/^�k$G����U��-NJ�en�}ى�Q���r�R���<�L$~`���P���(�� �Р�f�f��F+��5!-�Q2�e��ᵆ�5�A.Y���
�RVa�]A�̓jl�](�A�[B�+{���l4�-���-z�b,���	JmD6&�8�SPf�\��u-uLM�:@.��fƭ.yfV2����p�Ԛ.ȶ��u�(6i�-vM�4����m,����7g`\�S�WMr���UB�º�Uw���bī����r��L�3Y�G&�$9X����dѺ��̸��Z��(T�IYB��B�l��at��4�K�>���|t�rU;�b�9ãd�{�u7�2�6��BixɎ�(x���G."ͧ�锈�!@�d�������]z�9�i�hxzv�oDw�p���m~pA�%�����p�_�|E8�"��<�����r�vsT�y5R���=3�	�?Y�V|�����gv>
���>W�G{���h��{� |��H�?��z�` ����E�6�����~�=�1��i�RiR�ƒ�24=)��H �'IH��%A�zJ����ǟ�j��b��׭{�5�G��_38������������oMb�����K��x,4>����-��Y��k��˲�n�.��5�Ԛ,"����'�� ϓ�����;�O�Ef��mN���8�u�WDx/k���#�A%�!�U��&_�^��_߷��[��Gqq�|�G������/��L��D���D#�'R.f6���ݧ��gI�5�&��i��yeJwB�j�]I�!�̬��u^P9�ۡ�����UKF�c�W���6B�l�y���}�q�~E~m���Ɔ�tUeւаU�H�@��B�N����v��!]6O�Q���Q���
�����q�t��Y
I��xl}&�˾�"{�鎛\A�)4]8Il���HW��5�X��wK�K�i�������6=�o�yw�H�|���ճ1�����P7H;Z�ñn1�q`�&���g��g���U'�von���9����o=N�O;M�����#u�w��>	DI��M�S�/�:�E/U���u1ђ�6���bed8 ��MMJ�N�Nj��q��~qZM�p�� %J�l:��������Z��1ց]��ݶ[��/���*͗V������^��~])�>��m~!�^]���:[���C�T!)IH�o���������V�C����ܩ�~�#�����҃�,b����X�)��
�$+\8$m'qD�P�J���}��'�v�0��ڂ�7��ɸ?r�z�v]���D�?A��fs�z��z�ϴ̫ܟb�w`��z���҈��EJhh)��@B 33� sT�(�EL?���DLt{��K�7��=1/MRr�NZ�N�!�Kf@���ڛ�ޅң�9yͯΘ��4v�����n	_�8;i������� ݦ�X�q2��5�ǧ�w�ggE�9�M��p���鐪@�{owU.��(:"V2��W\k����Mfr]
��a,%f�@��<�6��})j�H��2U��o혳wQ���.<���ubӧ�2��"	����J�@W�}{k�L ���AI�"�È|����ֽ9yͯ�	)˱W��U!]����Ͷ�9�L���;�%���bvs���2�!؝��:'ZrT�,��1�`�u�3ԃ� ��I�������>�0���!���#=�w�w(!{�ų�DD�{�������K�DDg����I)�16�ЅS��z����iM��}TV�JM�`f��0�ڠ�]ϣ�." ��B.����f`|�d4����(5�RD:�q	c|� �j ���p�T��+b�i�/d=��q*m����_�^�=k����a'�y� �3�����~>1P��>��j���F�I�mƥ)/65���p(�����;����sl��X�'b9�X��LZҿV���}����k�o;�̡��<F:
�C��|$A"@�%y�L�T�KI���'�Áڃ�;�X���G��q��b� ���ŮГ�n9}���9U�����n������ÑT�&AU8w�eVyԭE������-LFU�6�LP#i8�8"�3�������o�)����Sn�	�O�]���}�sM�@GO�lLsoh�B�4^��$	P� �t"�c�.�x��S�u<�,�u��X��\�����̪��1jH ݮ^nq�/$yj�!e�Q_�Ҳ�Ju�8��]��]\ͻ�ҤY�tp����4�����u��wZ�7�d��=��s�H����@���hhAJ��}h�{��a�|������'����U	�е�6ƚ��Sc���C0Gj�!r��t6�Y� b���{Vy4Ye-WX6Ii�u���i���\l�[[��m��nL�1� ��D4ʹ��J�ᄴb\�v�^W��"�޵��2�[����
�Z�Lh57:W:��Ɓ���<�6��lsH/�$�f�:�v]s�]��=������ꙟ{^�;��^T�U���F�����	�!��u���aqͱfm+�b�Pe�Mj�%�����z�v �8v"�8 ��Y������2�9������{���NF5[�#��x��A%"	��@S�j��+%me���y?�w'�;��b9R�̵3��M͍�Ñv��ullV�!���
�P��d~��� � �|d����wP{z'VW��y�~�.���`���D�@I�og�>/}����p�����T���w�4w[�F]�y�����>W6!���R�`�[I�U��jzL���Ʃ9ʩ
��h�t�
�=�ܬʖ���jt��Z�^"J@�$C>֡_�[ί?>���O��ft��Ў�iui�P����*�2�Y���n�5b<��w���
�?�G~�A��*���Cv-P��A��X��\�#�*v��u`���A d���>�v��7h	1g����:�e��{3ur*\�==r}���3��1i4蝽�����3���42�A�^Ǣ�uU"�	�{�OP�z_� �b@� ��ңM T@F@�8�:���1�x��ѵ󚌻�@�\��4\�|�Ul�A�|2���D�P���^H'|���E��� �,δ�g�D�ё ΂��Dg�<پ���$�a���鐬B,�T�ȪC#�ݗί{�F���M�r;�;Q��\���I㦭�ֻ
�<Sa/�&�K�Ng��z�U�	�ӧ�PW�0�||F���#uÍz��}�\�Ee�4� �Oͥ"��
TF��2z3�fA:�z�Ж�!E�I���6MKj\�Q!b��Y��|Nw��N�I��I�j��w��������1���Ѹ�����"p�2P�@��W��^0���~y`�pr.�;I�;M����wٚ�����%RpFp$��<sY���8��O:r��,)�{G�+���i����8����{�߿<гP�ºvd�����)^m�w��8���k�Y�H3H1*޵(�*�Wb���2&�k'Wk�ʌ��qNĶeTUԒ��V���O*��-e�x�YW�uH1֜��n�K���ܾ�*��N<۫K��XO7vtڌ<b���0�S����;���>r�f�h��At�q�7�f.�cj���<ˊ��+j������̦�煇��y#sFICko�|w\)�v5����/��v)��w��<4{��bu<m^<yz����8��l��֪f�y;��%�јE<-I�S��hй���l��M.��xmn�<#l�Xj����uAT��z��wvwm]%��ҁ���ۺܣ�vwp�Ý;*��iY��2��C�D���ާ����_n����X̦���ZWY!�%(�[��u����]�'V�L��r��щ�ط��.�^����n��\��WA֪���t|ume=K��o<�d3*�^�1(1�a;0sO��b��jpג�u���nS��T��h�uK*��Qg]�a]���&.�)V6�l+�y���vĲ�i�0@�]h���
̭�/8��6�t���宐�zfKxs�i���Q���Y2)�+�����]���v�-`��4c���8V��f��z��Cq�U��δ$�P����K|�&��I�]�����]�pV���&�I�wbrfѺ�U�H*��B'^��F��<�>�� F]y4�q\��󇈊��)	ҐhK&���L��|"����J�Qk� �ʃ5*ԐT$�}||t�o�6��8��=|}}v���H:�E�MD �@��>�|t��q�q��z����۷o�r��"+ ȣ ;���|v��|q�z��6���۷o�yd�2&��TV����j�ok��ڢ�k���Үj��[cEck��cb������V�V�ޖ��V��\բ���U��Ƶ-h+Q� �j)QV��n?@߃J��Х44 5<�I���V�*��/9��#ڀr�ށ�^b�hH1I��h�d����T��)9j��w�;���Q���-�R����׎�Ӹ��~A$H	)ES�p^�]�Y�^��{1�j��f�W
��z�އz��r�Z��v�te<�Qޮ1�#}�_���2t�
���l��� 9 ��0[J���,If�-<�S����~xH�[�-����ۻ�
^��_��n<����<�������? ���� �' �j��꛹�lnkFF��m,�-v�k��,��~���((/g ����H;��;ŝ�U�wP@�ԼF֑C{�U;�����y���1��ǻ�Q��_[����^ �*j�85I�Q��a��$s���8"�����|��݅^��Yyͯ��փ�쁌ŵ*f&Wq�|�"�Ɗ�T���et��C�b.�t8m'�1�i7QY���j9����ph;��R�y��Kz�^)�;��0mn� "��i�����C�鿬���W�1�M7n౴��|��|��o�r�w���8bA�� �X��RAN�(����>��K�ƹPp�xrӾ���76�F5YI���������؈�iC���ru,�A�p��]õ�i�u���$��Ҹ��7��qԺ~;�l�i��UÜ��s���s����}�=�2���p�1���	둪��o��&vz�>����u� ��/I��1� u�?��7����^��_ǋ�|z��y�P��`��wS#���݈9�K���T�Uy�nBܸ�X�8���Ʃ�۸�Ln����߹����CP�7��V]FǛ�k�G[c��L�z��T��� �Aj����	�m�ر]�Ӭ�p��wv�������Z��m��؋�ڥy����'��%�+ܔR���cN��	��E9C�fw�z���o���f�W}��y�%�;�gv-Ӎ"�J�SU��5r��__������A�w��VW�̹W�%+3�$B���TQ��.a��Lk
B�e�hѷLV����� �[j:�kj��k.��.�0l[s�2��.��Yn�e�`�a{ǥ%%t����1{qLK��0�Lb�ڈ� صIZ1��V�\$a!��83����X˸чl�5��١4	�$�&����fMf��"m6�A�4B�`� �0���1
w�V�Җ�r��3fV�j�7hX��iV�Y�T�6��]va�Z�����xx/�W�r�D7T4�p,j��Vr��1���pp�M�'&��W��p8o�9�AȪL�!T�T�3yoܽ}�t�\�wc\����c7yrqv&�ˈ �' ��g�I�݃��n�GZpA� �N�H;y
�/׻Q|$��H=��/�=hW9��pbJ>��	x��^E�@��Ǝ��WE����,��.R �){��u�|�;Εp�M�z�v"*N����Wz�ֶ�c�o���.�t��hdۇ"�1��w:vm�҈,�Euڍ����\��� &Wd�vsv�Xݬ���S��٧킐��P�7<a��T:����dm�3h]uK����� �-���C3���2H@}�������3��a�t*�#9��=�P�E5g�p�nݼ��KS ����:I�ۧ�e�%��-\)�>/Q5O�{F��pot����t>U�9d�F�.A�$M��q��ږNֳT�.Q>�)d]{ݴy�+E�DQ�ߞC���M44R�C}�=�}OZ��U������*���q��U ��qޟ�P���A�9�9n�$����v�ٚKu�ѠG��o��
�*��\�v���L���Y!P��H!ه�H��`H�� �A a���~�ٿ�������p�P�S��8(��;@�p"���4��A�y%-������x�H&��w��x�\p�Ԅ1`Dc�:ُ,|A�q����4a�e�+Jk�wwPR�3F�&��uҲ���z���Eæ�~��Y�=�f�����la��L���i�u={[������Fߗ�G{nԧZ[i7��+b,ܦ�@{�Lî�aw�cY�@�"�È���f��r�9����fL4�"�~�4gY���qd)�N�"z(|�g�xѻ^s��#|���/E�̮�%TQr��Z�m��{#�KW��Z���sk�mWr:6��]�gG;�w[ƪ.����T|-�2L�&L�&h���"!���跏Lf����J�c�,
����,� ����`^>�v:��[/�Mښ���%҂5I��x�96\�kS89��2n�5��|h�x�yš��[�����1���^�Z���!��;p �.\c��]���dz����>9`���ĘN��+.��k�r̺\2� �Ä���!̶>+}���C&�R ד����F�zc�t8A�1f�-? z�절 ?=�~0�@�7PPΫ6@�9MS�^�OV���[���M��:}��=��=E���5)��Qj�GVg��S���}�YЃ�z�r �>��?nw�˨q���f+�TE2=>�^�Fs9��4d���ށ]�v6�ɃN��'���^}�U�U�8t� ��J�����`J�h��q�A�ǟ!�c��k(�|������l�Zќ���(nð�/���U}��X�k8�zhЧx{�%FϞ<�/H��&A��&3��?;/���<�]@g�yY�E�`�E�zez�D������8}Q՗�i����� �H�+��O�Y���˫Ώe�F���n�� "��	����^�B��66�V���+e!��=����'����G��KA�R�A�=���l���g3��ȋ�*;��͙� or�8ݐ p᪓85I� �&�9�o\���.�sԜn��q]ѱ�Ol��C��G��nЌ��2�\��O��p���pX� �CU8	�� �쭮�3��w�q]F�O^��R���'`A�p6��elA�Y2i�s����Y��z��C���yc35ד�S��g5�L����9��=f�=�����źݞU&�^N����Q��[��c��p�W'.�w�ޏN�2/��|��M2�S��g���}y9=��Tفqꈪf	sГ3qh�{�k2���+-/p����C�G@��v~�v�����u�AI77��ňjYʃ�g��4zh:p����=eЋ��۶�氄\�u[�tkU,jٱJ���F�[��� 4�!��]��d�Sb����tpflm	�Ю8��+�qnQ�b��),c�],pB�:�Z*��l�f��It�D�mКl�&��b
��1��C "�\���M�n�� ��T�/8�#��(�J�a6֞՝x'k�ݒ��,�YIS6V]����ti����yɷQ�Q���O�E!��A����;1hl�g���lL𩧯_z�UY�*Mَ��*��!T�� 昡>F׻ � �x���3כ3bk���1Q��(8���Ȫ�A�bA�Q$f2�7s����vsT��j�^ǁj�<���|+X>. �ҩ�K.r�LR��Z�¦6���ϹC����=>m:�\9�/d�4/�����"��9^�c�C�o(��Xb�Χ	��PBb�ERj���y�����0O�;	�{��}�k�����R����נ;T�r/ض�?���y��C��� ��+4vC ����"7R	�
J$�r�K7��ڝ�/��,�L��'-4�W��Z�u���`R.L�%�V����3��sPr�p*��5K�v4q��tm�&y��M:9�5�̘�2eqz��v�5y��m�B��9��;S[}{��ԍ�G�
�3�[Oϳ�����znX�,C|���"����ώz���bg��={:��T��"��ݪ����=}x�c
��{�CHy�T��$ɤ����w���H��˟l���9����P׮*�8�p*��5�;��jwj�Q�A6�4�pAcvY;@���lmr0+���A>��7�?]Ra��PlA"% �@I�?M��)VX�gȁDwx�v��;5��<=UY�I��' ��g�8 �T�<cIz�@�9��Eᜨ�u�R�̑&�(e�0U��흻��*~������y���R �~o���5�����"��C:Ν��Ŧ� ����M��nԐM�v!v�҅{�j��i�uް�֔
�c�����i_W�>�p��}�^5���qD�/I^��ʙ|���ڍ�Os� 陇&���vu�*�\/��w�^"z�k�x��'Qn��Y���}ŢS����`�O�,C!��)����y�UQY�+�]L�i٪���NER{|w$���|���8x���Ȍ��n�렯+Z���E�!�EJ�{�ݏ��A��DF&��`7��销 �*��%*M,��n��8*Gf�[���p�or�u��U!��f�_���q@����+���st�&.�ɴsc4H��rE������?:�_k�̆�w�b-YE�9��׉<=T��2��įs���� ����tړ��KBl�c�BH���g�~nX��\.+Z�w��܎�;r�ek=s��� ޸r"���2;=�j��e�8:��Q+VC�.�kȾ=%~�4��_���WC>�O :�&�E���E[�-|y`�׬��/̠����J�/v��g���U=c��\Ac������eF���{ϑrq[�/����ç���к˥![�&T	~�3�#B3��gxw���Y��nk;�wRm�1�6�?�K������8�0}���S�v��K�����J��;\�d���U;�"$\�Jʳ���߂��)6Q�	u��Gf�Nf]e1i�4.ѫ3}}�-�����	� �1Yj��MR���nGc��pC��!/�u=(8 �]��GO��PDH�aEx�?���'�d�-�����VC͏vv�y�T�~���Ne�	Q��-��顦���Y�6��A�.��N;�n*�?���5$��WӲ�os�^�>�zBh>-��p[�n�w&Zv!�իx:�;�Rj��9�BX��^�|zx�|�J��t��X�v���.�ݗ�ŔA��+�H(M�N45 �^W�\f���͍���#'4�s�p����&WA�M�Jȓv��� Ub�;����
����;o��kY�O7X4NM�ʽ#v����Crɭ׊�^����ǵ.c]u{jd��m�Ȳy��A���32���w燫2wl���F���о7A�e��Wb�V'�h�	�bMh./y�kf�˦k->��]�^ y7W�L�v�VM�][.G��I�ܳu]�2�w5i��̲v��uc�ꪶC͸����z.�t�L�}���Ħii7��֞>�i�op�=̖�X����6�r-�+oC�R�.��Zx�=����x��nC������}2�Yҍ�Ω\h,�LK;n���\;g�u�XM໌��s�k9q���2�<N�r���b�K3����аQU޾�;w��[Q��!�j�e>ʫ�;z��쫝��ؙ]7� :��=�ԶU&ŊWt����wp�%��櫍�w,�gSg�8�cW2�}�"�7����
���Ǘ��%Ɠrg<`3MP=��FVU�u�W9_w��*�u.f�d�����E�KoJ����w9Oo3�X���%��Ϻe1T���V�9m�K�&�.�ŔI/o8��KG-Hu�C���R��]S*������fk�}�X6V����U�k��wme���f�
�tbIڴ��+H+����w.
h�&��Uӹ���Z�Ѧ�^�+��5յ�[CX]����Gݼ�co6(j\�E��b���ib�	)���z:��m�հ ���P��$
"�h�$�U2�*�5cn>y
E+�x��K�C�xl�J��m���o������qǯ�q���nݻ|A��Q}x����N�q��qǯ�8�o��ݻv��@� H⇐�	*5��O�t��8��z���}q۷n��	"*�EJ�EW�(\�"� ���"�P� 2"Dn ���A.�w�A��47#l���h��؆����FkF����UY5X��k��41f�~��{���=�Y�,�f+�u���1l��.4̓nI�-��PBF�괍M�T/U�Uv��;�ѹ��iZTε�[m�r���5E�%�ʌΗLGD���6��f4�kfe���u)
�4�,��A��U,���f��[��R��im���&jh��b�lM͘8�Zv�jYq��4��a{SdEv�iYDYsٹ.+�0�f�J����U�WF-��J�X�Tl)�;1`@CF�� gb�`���CX	�]f��M�D��eMWi[2��Jn�٥��ҁWq�!��̳V2����2�YF��02�5�Pn���f��{V)L���v�ib�y����*r��m㴕��ns͹���&��c����I�0T#F�ճԧ1�efe�ZD�b�9i`��H�B]L�e%�ͳ����s�Gi�J�鰻3FWV4���u ���I�������UE7W-2)HTp�0Խ]J�A�G\�Ҍ@�k��c.�Y���)N5��K�6eb˵�-`��P�v4�	P�bS5�j�et4#��ny���G��۩�I��^Ö@Ki����+6&�/f[f�"��M6�4��"ո��4v��Jv7b��Sq]�e�����+��n�a.Qæ�l&.F���R�4�ʖ��k�Ö 	���V!R��d��Q�;[	]"�m�e�t�C;�2mŁA�Х
R���).�Mk2p��Zd��j7;E+#
�%��^
�.J�Ka�d�el��M&���n��8���(��.V�.�bd��T�Y�h6�0�%� �n^b�k�٢&R)������p0"�k2�\��-5�m��XY�)G\Y��,��*��CL��p��ܺZ�Ѹ�dq���J�v�&�9�k���,��4����8,{0���b���ͶX"a�"�\5���q�������lTf3�p9�k�;��1X��{6x�G����o`��H��	;/[kuM(�"SS`�jQ(E�I�u�4f�*����l�T琗.桰�D��#��!pQn1�m3�ҥv��2�����ch�0!U ;U ����Jn��]�#F�V���%�՛$H1��,���v1���ɶ9ķVi[c.�l�a1��F��`b�t��@�։�q�mRIR��tڔK��Z$�ΪXZ����)�Y�,*��uԂ��Ѣ��!Nԗ&�hփSJ�ka[Ku��4ŅT�}hS��G�y`Sv8�k�cF�!�E�y�>��V�ru��Ƿ��g���r�-�|Z��́ �佧H^2P�2R(�_��ˠ}���ZŪ�f,\V�u�4d.-�@;p�9Fk��=�۳L9�7�0��X\�`�{��mc۽M�V�@�����>��=_zWi8 �ӳ��R�A)5R�8�LV���@Us�c|��*��F�}�䕩��z�����fgVj��la�A��4��9�g��^E*���^��t�l�kul'(��寱�_�8a��38�p�Ѣ�T�;n8���,��qK�IK�5Ĵ�7b��n���`���HC[o��>:\�׮W���Dc=W�����*)��Ҹ#T�e(阕ءax�;�� �N�Q�@��襙�zD�b���1k��Y�����n\G�W*�n]M7��l͡B9�"���\ӳSMt�I:���N����{;�7,C!���.똸
���)���+YS̫�|d�ָr�hzߔ]���)p��2�M���Z��]�n�D˽Ϟ,f���9�0�%g>z�xg>-l�k��>��0E��o�w�0��̚G�k�F�v�
���~��.���A�u�A ֧ ��{/E�e�t!���}�^Ӥg��T���E�ҽGܺ;��h;&�
~��J��y���2d��;T������y�X��(��ʤ-��%*���2���1�8͢��l0���!Yi������x�������N,5aj���R�Y�y�~�S�0���˚sz�i���B�:���E؊������F����4z->訊����MT�����/���E_L =��J��K�A��M�zli�O�	.0��@�k�p�Bl�E�Y� ��;+�g;;,�Y��_}H�{i�8��:����.�m�W���uS��x�Km��Yb��������N��љJfeeq9�ڧ]��{���RA�-��W$g��߃1�賈���Roʻ�k��~^,�A�9�~"���P�Ӭ�9��;r�L� ����-A���Gz�z5uR�#�<����r�ǻ�40+S�-���,i �T�4�n�Q9&Կ��ic΃�#k%r���FX0�Y�N( �3I�i9� �p����/�����@�?q
2�L����Y�u�
�����Ă�7g]]��,]�T ;(� �R�W�;�ح��<A�㲩{�^�!�)xDہT��B��Wj��r=��<��4u3��r��}���?i�5C������ԃ��$� 򪼭��x!S�غ��@��H��$�$�zj�a0�|Rr��+m�ez�.*2�t�q���ƭ5R�-T�K&��*��SáŪ� ��u�S�o\dڌ��1���O����&���QS��hJ�3�?%�wt�u��
�U��J���l7_l�����oVuGx�������wT\�g�PwUx�n��e>{�X�,C] &9�����T���AY���9-�z��Q��6���j�{$ke�4�A�Mx��@8 �������|�S�t5h��<D(� ���@���vh��f��^D�f�J��cOg�Ϭ���3�pES������:�G.�&2Ȧ���|��O�ݼ�}� $� �5v( ��<�n����痞�4?��Ɗ,+�o�8��](������j�	)��(f8pGzЕ����%��9h8M���ͬ�+i��x*��A<���^���ݜj���ת��5_�� �]�b.ӂۇU;���Y���S�]�O��o\9��E*!�ɵ�ˤr�2c/���� ���F�6�q��N��I�$�%;S �;�ȳn ��ʝ��F��<�	���F��4w�=:�T?x�e}܂� �D�E��i��X��|lY�J��>7U��Tr�'�˻V+!g��1�n���[���a�t���>5�-,�zn%ŷ,C|���X�K\s>��o"��_�R�}j��5��7�:�9؎�.)Fa�B�K1���f��P�7*:d�&�0h�.J8 �,�\�n��V�j�m��%ce���\�;6��ٵ�bXji�� 2�ob-e�KaHB�@�D��d�16��m�#iJ��Dycf�u�u��2K�c�7�CU�WAmL����+�DtŮ���3}���>�U��36����l�wd�=��ʡ@���	T,-R���;�;iE\]�v�\ "�u�^%u%� ���&v7I��x�.�՝��b�VkEp'w�z�F���)U/ժX�����q�E��4<�)zl��#<����M�ֿH��(F_L.`[)8-4��n�Ū�@�S�4X/
�8 � ���
��"�	3q=_�x�;�U�uڸ�3�B�I؋������P����'^��p6c�k|��A�bv �T��oVvw���{�̴���j�֩�@��`�Q�" ���n��O���� �q|��r1m���	��|F�z���d���u5�&B�.�����MJ~�c<��1��C[�S;YsFmY�⡨ʈV�4��-�,_�ߜw��2Yg�׻�2�3�ܜw�<�_aȞg�pV��\D�-=���g����Z�8"��~U�O��t����fVٽ���~���ʐ��s6�nl}|�DV.:�����3y�f}#����lY�"�W��Ĝv�ňb�1�z��vS�n_r���U��M�k�	�A�y���I�mV\��{���{�;��,��p���@3~13�S���9 ���UQ��.�^��2��Ų��K*!�RpZ�9iHw�u]��%�e�`�QLAi��㏔5h��q:�\ɜ"<P!�"��5L[~��% }%#�|�m��h��p�cz���r���QGޛ�k���c�f��� ��e���ym�tj~�F����e@�К�qf\Y�t���Jv���	t�D'���GA%ÀD˻e$8�3����Ց(F[��MVp�|��tE�����=I؂�Nť	�@j�+Tмs��	,����*����*=�Q��GX�Z�UX���KX[!h;���A��N�y���՞���;�"��G��|��7���^�r���V�8u=)^��[eE�GK�&�O��BB��,����M$ c�(&�ňb�6� �~����1F=7�D�@�s�pA�$[j��]˰�d֝��#f��>�dO�;DB�������!�6)sLbr3_�'v<���p���Px ��N<�#K��X����+|v��a(�B��0:����sx�ǯsS�vo^�BT�r���5 ���i�;,��]�TomwSG�*��n&j����a��ѭ�<7is&Ĝ��3)�-2�s��fwQ�^�Vw����e���z� F�! ��#��H�!@�h��?�,�Do�[N����!2��tk���I��;��؂k�!2�0滊۱��G�b@��"hl[B�4��g��B�q�J��op�ǯsS��G�bP@��C����T�=����o��X��9���"i@�ڻ9��IE{/9���������هJL��I�dT^PUo\���S��&JW�Ċ;��ν�L6�����L0��U��FJ���W]�R�	��j�����3|=� �?0cUG~��7�.HK.� A$�Ў�/��[�{���ڨ��m.���-�1�%i�����rC)�N|���0yx`�H?���5��Lc$e�F�]�H��&u]�[{��,YbA�	���0"J ���V�d�Ï^�=�5鮓.":lI�K�g���n��t�@¯�Z4F��b1�[9��=�r��=={/5��� ���6���۟P�Z�x����"K��L׏b����&�����SU3|����n�X�'2B L�s2�b)�6\���sɴ�m�#�b=)��hY����8��e|G�"��lw����3���3)����L���e�ڣ�vji~�� ���7�f����W���&�A�y�� Dˊ�Z|�gp�qUFm��2�U1Y���ӱ���6�j�u�Q��B����Sn�.:�HmT�ag ~���F�Ϸ�j�`�[�|�H��]י9}�C��ި�����0c����}�S�����=��}S�p�#f׍�]���Ț�yJM�R��\ن�ꂧ"[s���L�,E�sK3qjB�oT��*3mA`��.� �v��A�͕���]�Y�A+iyU�H�	����v�[K*� ]�0�
�f0�A��"f!�h�����F��lX�����-�Љ@�M٠j�.&�.�8ᆥE�/l@�Tw2�]�1]��r���5�˘�ת�E�vB�	
�DQ�ey&�]���m�� ���G�(?1�\AN���ܸ��l�S��u�C�p��NwN�j�zױ���	9ʸ�#7�,�fz����@�Je�C�E1q���
p_���o��ıDN�M�"��%^�x!e�P΂5X���B�@ �[�v)��<]�>y7/
�BN��-u�Y��\e�5��.��1N���-2��2I�o���o`&H/.5��<��5��('Λ��n�:��g[��s�F\{V���/��v�#[�t��[�>���"dAx��@����:���Ë�����ى�\ֹ��[.l��@p,�W���mȨH��_� ּR��� ̠�l��f��h�P�j������Aڙ��j��O�ەh��B�2���ǽ��y&��B��9I�5NC!U�PB�b��c����qaw���85d����ް�k�j�vQ��H��3����2v�wwE^ʢY4k�;�a��U�Oݾ�`��{a�|m��-VtW{��\�E��k���L�Z8w�X��F�`>��{6��$���J ̸��y�o�m�������s8,MJa��{����W\o2�����ͯgnͪ�sR�Lʮ��������-�|ȔwP�����6�0#Mx�'�~D�hH� �k�@7�zy�CK#e�io.���.R������s��A�5I˱F�,#�f{>�y�N��7)6u���e��g�!�%B:!e)�kl��58'ԑg�p�D�H���:5�<��c���6"l���	`�$N��Dۻ$#2�ZYN!0<�[c�,�Fm!�b}��q����� n��,��8pD���]a��8r6]����t# ���]k�~�j}���F�:�a˾����P�ΰ�vT7c�e�<�Pݮ��^�fV����U�r���U�R:�;9V��E��_o$z�]�"���~=z3�81�T2
��78�S��'��ov�J��
��6�� �-�R�^��Z�I���+֎���JNfQQT`��&͝m�A�\��}ON�v�u��^U,Dm纻sM�մ���9op��OI�3��_C�s7�[\n����X��U�n��za$D0�Z5Z-���+���&e*}f�����=G��V�emK�+��r�(�ٞ)挾'���y<]#ܼJ��]ٹ���GpS:���9�����})]>���]!�:�ty�q]���u��	2��m�[Oa�a�������}d�J��U�Zݎ�:�L[8Wv󵰪4��d�p�x\õ��3�[c*�(�ۼ;�W6+0ou��U�*���c�8�����]�1�N�9�se��s8bظ��kqd���{G��]@�ք��ɇ�K�1��f��𦲻��9ݜ���^�nV��D��ɒ�l׬ɴԋ�*��D{�i��ji��}gIH�Y;����ޛe\콝yخ�7�Pٗy�,��B�f�v==�;'j����-�m�x�vF
i(
�4!�)4�z�|�I�L'�JJJ6�p���֢��O=�thLI]F���D�	{J���t >8  �v.�k<QKT.�7��\B��qu�e[���g���vt���GJ��}���������eEC%y���|	��$_i%�i|�-�6��8��p �J���!��y���H��g�}a��|��o���$��OEit`�v=1�茸�#��*���K0 n]-E�F����Ǯ�v���:q��}qƟ\v��j� �"��dBBE:�����n�8�:q��}qƟ\v��fv��"n T0X�.y.$�p�)"5]>;vӷq�v�^�}q��]�v� yȋ�Y	��&�^>.�h��^V�-�!�*��D&�N�t�d6�A|i�<+sk��jwh�(�d����[��	��؅AG��v��yxI�m�\��,cU�c^��6kJ�ҫ���x�$v�ňb�6�wyu�����ٻ��A7���BQj��G��8�M�e,@�̩/�zו���-���,d�e�!��D�{�e�[ُ�W�m �,����ף����Ec�H�$"�3 I �ό�� Тe$ӱ�z�a?�jEF��i�2�������I�e�\��<��>l�\�Μ�A{M5.�+�vR+���qP��
Y�޻6~o�=*�ѡ�.����8$����?>�W'��^��v!�Z�7r"��3����g�M��� x��o|�o�)5N���A%�7dm����=sZ�D9n����~�"�$�|��̼e� L�-����ڤ�BMf�5ؐI�U!淒4��Z���u�
\8�T2��p�Ey�Ƿ�h���yve�+��Ō�3��ǽ���O��Ł9��in�tk���)����2f=��Zg��F�5Ze
S@�f8����ldK���]gJO��w���.��<�{�����c0|g!�/Ulԧb҂��	$	�2o�zN����O�7��u66��<�sZ��۫<l�^f��>���]�C�����lݵCs��JC]4*�ɱd@�a4�i��'����Ē�"+���)Oz����z�+yc��e@�֓cCjD���]�y�-��0��OZ�M�-�*}�z�J̙�
�,D˸$�L�kv_r2��ܽO�����s!�@�Ɍ���ٔ�{�g��\4�&�0 ��AȪND��(l����CE�$�x�w�q��ɋ3��e�Fʞ@�����lwEI�H�^nx�OP.�;@�����qWS�^�;�G2넞�փ��y�z=o���s9Aj�I�p�2B �2�L�l�~C}�7����i�E����������G�'13�MCA�L��:��`<�.����x�4��d�*r�����/er	��a;��]B�_|��|�_�H���e��N�2Λ�r`�yAp���J!ۃ!��]��8��*�|��R{�ﴏ����.�]U2�bS���L����vQ���3��е���6ـ�@��`���Z�Dc0���T%���),�N����`����m����X��,q�@*�����)v�ٮ2et��G%1���-W�3��^���Asr�s M�\���n���&�1c)��(���Ŕ��4��v����>���xm.Sg���e�"����Ip���:i�����Fj�ˬLG�)���Xn�&��W0M`3:�a�!ۘa����p�HLA.�w��3Mw��;L��C="�^����>�kn��ځ]8v"�"f]���oui޹�N�e�ZL�r=I��Nk��O#��xI�=I��$���ZUom*���>��O���A_P@�!��6l�C���v�w�:4�<RLü�:s�O��u��k�Jd�v �2����[nU�>�Zw��@`H;�L!�-�v� �5��E���Q�K��|u��pA�1�!�zk��ۥlV�j$*L� |ϩ|[�2u�?`;�bࣝS������<[�0pAƝ�y�� ���9�V�77��6g} �B	Jt^� �e��[a�y�$&�eE�bŉ�`R_C�>~��ϫa��6k�T[�:b$A�1�������D�������BiyL������Ze4�"�[�dN;��5Z>c-ڬD�.+@���d{��oOW�+8��`��G�Zɻ��y�]$�&�pi���]��m��f�ud��c0e�|'��_8v��c�gRΉ�h����bɨ
p�L�����q��}��ƦM�mA�H^�ȷS�~B���c�ﾐϿl�(�x���Nкz�x1*��b$�N��)�`�HDL�&|�+�D^�ڍOc<E��p�hmÒ��WF>��3�����	��y9Lm_��}�z�eP�����H�@���$E?�A):R$M�x���{s-tNsFإ�����{C���pI�!��> }Kv���(�bP�ְ�Z;^�&�3���,l��&i�L�'�QZl"O��yx ��vc��s��iML�x�����,�B-���A���B$A"��ݬ{�L�>�d_�؊M�����}=�ǝ�\ �'�C�F2�G����1�O���� �'qd����Ƙ!Mۊ���IԍV�^S1g�b|�qA��Rt��UkP��ܮQ(�o\�Ȳ4$���`�Y��c|�n�Jb�$��Rv�˫�1 KA2B,�8^R-��ňgg��}�Σ�9���l"�D�x���Fvn��T �Uh?���FE��֕S�7�y�c���,nnx��Uk��_�G��2o�_��$HIf�-��mo�\1\i�W��w܌�1��y�ԇ�؝�&^-��� ���w|'/�$]��M$i'�Qr��1�����:;X�+��u4؛ )+�.O!�h��h8�p��0�8�q��^���+��Ϻ�����@�ɯ� r����U( ����ự�!8�b�1;p|���z�z���A� ���p�I182vS����������)���-2��c3�F�DO�Ȱ��-�'���vcٓ��\A%;��E�3�2��ȮE�c�J�B����@�q���LT�Q[��}�6�����gz���K�Q��U���`&�*�̉x�x��x}7���mp�SM���8+7�����:c�.��7�Eh�|���,�a��Rj�e�c!%��ޤ��c0v��>C���������[	�	/D@5���/��Mc�v��#^B��ڗk4|?"�YAx���3D�-�~|���|_O?�_�!����bh����71��]�0�7
�e�����'�e���e��ע�L���Hp4?{�u̼�:h���qޡ:v�d5����n��d�e �����Bȉ��l`s F�do�*vt.�i�)!��>."�܆��6���z{� ������&-|�A��c�ɏ��z�zd�|��IP�}&x��媈�DN�0#%"JbL�t�L��ni��:[]�����wbh�-�^.��}�㉸�&�5�j�Oxo��М��tɤ�3(;DˢNA#�-�!�,����ݭ��
��H|CE?�vNER	3��4�,�������,ڜ��7�y���vmp��ϩ�#0�#\Z��+�8�=M��W:(B�T�f澦j���+��M���b��Uf.�}�����X�i�x���2����2��a�b��\f違V;ak3Qm�����MZ�ut6��2Q�H�nк�(2�R�s]���v�";JCWm�4���m�v��Q,�,tbr3QK))5���b.��ԠX[�jV��l�kl|�/��u�]#q�f�cf\j��$�ֵ�s��	�
R�%j��o˷C-w��n��&M���9�/���Օ1`,ݠ�Fn�����k������`��b%��q�WƗ�n�rq�-��D��Rv������T��Ù�!�;JPf���`�����U8r&]�D�A��	��_���s�d�%�����q噃��:ew-w`�d�:�LQ�ʩnAj'ēd�W�2����� ���Am ϯͤ^1O��p{��}9�̿a;=�>h��☂*�;1����Hv@L�b0{c��!�ԮIa�i����j��Rv�����ޤ���bG�NKb��׽R:���D	5�=�HCS Jt*��'��ٌ�LB:q���<�,j�ǺN��q��ed9�NA3+=s1[�$�GzyX#��,��f�W:غb�j���Vl�D��AJ&�)�q�w�%�8�Q�".�v��Nx�q>�Vowq>wc�&�g@�8L�u8p(��42�r7j3vF���f檵kh�o?2g��+f�嗛u,��@e<�&C����}vDX��8�ְ��	��IY�Og9j!������ϒIRj����9w:�en�F{n���q���a �r$��ra�`~؂n$5�Ctח�d~��D}�.��I"����5�a�ko>gc�&��dL1pfS��O�M.�!u^����U�.9�Ÿ�ˇ����g�aY��8(�=������+<A2O/X�'n����Xb�>���;��Gh��}���W(;y�^� D�1�T�H��868�����-�w�4֖�AGCcc�е�HG'��|����b�p�L�$�q�onڇ��I#�� F�:�O�Eסǘ��-/̑�$�feXN��h�e����y�+���jV�V �����<�,�}́�hDh�A�=~8Ey_���5i��x��XT����"t.�)}���q�+uj�JT���^\S;u�k��V�e�rz�wØ�o�B�S����6���1b�f���E �OCvZ�4i��r�r:�r��r�p&|_ti��;��)���N��k݇[ל����{R�H�M�s�7��2������Hw��W���4�:�Va������b�ÉY�M�]Ζ����U8r*�ؙ �����1�7TQ�Ƅɜ�r�<$���܍����Ζ�2:6T'.%������M�o�����v,	�O�)N��/4�b�4�a�ܟ&X��������kAo�\7�	Q6���^OY#\�U�����v'�����9z���@ի��j�D1�V�]�f�h~���I�1L�3�<(jeI0�(��遚��m'�&7L�j��182��,9�����Ae�p�3��(����D��,�L33gJv ���L�fS���u:�f�\��;���4)H@8��7z"7�}�N�����4!����Z]ը�	w�J��f��r}&�iZke�
�umQ�#���T1�����ܐ�}����B��%3���D7A�h��_e������	�Qc猽�{���W	�Nd!�*��J���������'mR�K����k]��n�ݦP�ck�z�t|����@��@d�`�D��S.�?{�����t��.gE���F����`Ҁ �P@��Y[� g�� �ܑ�p�8��8�� ��;�.�wW������ipM:4�P �4s�6�9?cH8�!}	'�U!�NA4Q��1�z�qǿ^e��	�}A��ZpAˋf/MS�-)�U��Q�5��41�C�iDL���7l�ѵ��f�$È�����=�:!�#Axx�f��lfB�k[�oUe�Q6Bec���|(ţc�����u�^�� X��pFJrA&JL�ǘ[s}�ҩ�|�A��R�*������㔩�egj���9���6�t�J�Q�c�l�spǽ[z��+�1[Yis{��]�u�oV�ut�O��	�=Lv��Ufֻ��Y�_����=[���\R�^@�c��\�j���y'�7���q�ɢ�+`�]�q����zƹ~�v�y��x�V)�Ԭ�*[WUr����(�7Q�wN��
��R�s8Ws��ؾ�fbh�*{���f�;����2�E��UGc9���.Y�۷}Sh!���i=V��^e.�L�ʖ)y��.�y{\��x<o�]���9ۙ�澙���H��k0�������,˜ua��Y@�ٲ�Y�Z�*��]r���p�6qR�٢4y�5�U�v#*��:��Nvk4�=8w�t"��켮�sy���Q�er�1\�w�5,��b���Ր���먃��,���mR,j�\���K��S�N�{����WY�Ϭ�*r������ݷ)��iұ�I�&��\,fw;%Iv
u��^��ٱ�x�U�rœ���ǳ��iUꕱ���>�ߣ�Y��Y��	��^N�ע
�k���.��e��=K��ٻm�pܗ�v��gC�tvVLu�Xbn�އ;e�ڒP���o�]�f���Ǯn^μ�6���hU�*��y����4Wm�g;n�4pB�I��O'"Eۈ/����-�3�O�����M��D����� D@XbPEyS����Gm5��e�M�}��S���|}��&��O>��/�kh[a��{Ϗb��jz�QGT�B4�Y�3*�� �T�+1�DzO�'@D����=�5t����捋a4ɩ[z�ۧ�;x���v�^�~��z޷���fd���,_t���fE��������q�qێ=z��}x�Ӧ�! DE-_ģ1;�(�B!����lv�8��q�ׯ���N�>xH�H�T��$]��*��3k�R�/(��QAEh�A�b#��U�],�,���Pi�:�u͹Ҩ�&��wt���-������DQ�.o�x��(�a��E�0{����I����߈_z��҃��z��jz%5ҡsGhb��"�]vW��^A�mst&V.n�B��L�s)Ð��Fa�-3&�n6&n2!�Y�Uͬ�1Q+�R�`�bv�*!3��H�,T.��B,HM��`ta3T��eИh�=H��.���霦�c0h�F���j�iJ�4�\�KM&Z0��Fݝ��X��c��F���l����L�R�b�bZBWYI�&,,�cK�\S6��P�0b�Ջf33�R�8��ж;6ӛ��V���"F���i
m�$��gѺ��� �k0��3Vb�h喼�EM,lٵtZI��U3`��r$��lU��c�ŮAѩL�44�К���,�Ͱ���g0u4��]F3X�³k3�,�X�m�W��)�@VY�M1IA3�J�Zjfr���3M�.����'�v�1T���,��rGj��j]��9H1�(����>��޳a���{]v�ʫl����R���7[���4���u`��NP���{jܳge�6Ma	���BT�i�[�Rfl:�\�ޡ
"mf�Ө�;�9��5�e&���: XЉ\SD�F�ѯ�0�M�l�4�	�@�l�����l��MTm��V�\l��ͦ&�Lݖ�q	k����b m5��,�������nS�%��3D]`�bii56s�b����q�( ͮ�L�A�u��d�K�i`��*2ئmƊl]t�9�Bd��5�.Tk�����ZKM���X(лXF�^,(�c�M�W[
�L���@�ch8���a�b]����Y�Gl[0�/Lh.SRR��f��SkB�cs0�2`�%���4�Q0��k+�b�X�Bh��A�8�&k	��..5�b;V��4�$`Kl)jjd]��x�PCkG^�0�C"��U\�3n�4�.��=�۴�oh����ņ�.���R�q����=���/�ہ�MnV�1���1��ّv�/�����31e�fL��MS�����F��+{�!����y/�P�,��_�Y��I���If�Fb�^@
����.�)i�eIvE��ړ5+��bljcjWB^[u��Ď�L���cVPX�(U�l�P��.�l����6�4��YL�#����o[��DЮ!�Uh3dA[aV$ �u��t�c�愩rR�f�,� �K�X[GZ&()��e�(�n����[�E�x3;�]��&`�nڹ���7���Z/�̠�������*��6�,ѻ\K�������$G&cm��w���aL�qg���*�ر�T��=vWUO�p�Z��wT�(:�K�>w �x�v�9�N��k�7h�cMP�!��x�> �8'�u��]α�h��x��.'��y�:���lb����"��^>2W�!IL�e<RS/|E��~�tVQF0�H����Q��{/�B��.�����F�A�h CtB9����P�d��!e')�4A��P�}]7/+�H݅�ɮ�1ry'��ɺ�#�O)�'ɥ���Ŵ�49��ܷ���z.�o���>���Q��u�3G�0p � Z�ÂH)��%���B~�#�DH�z�6kn(�.,W[G��,#,��a����#az$�?�M���1F�8 �-#��)4�h�����{vy���NLdfmm�Ȥ�N�2��Dˇ�!%�������GV/!�9W�"�0�X���b.�ű�F��iR�8ps9�e�\ٺP�0��+u4`4�k��&nX�,C-C��ؐ$��4W�k�jz��n�M�h�r�-!�JS�'[��`�nӻ&�@�e����p(�j�?FN=o�� (�n}��}B��]c��|YAD*\8BRH� U&���c�cW�,t��pA3)���>,�;�j$pLg����ܺ�{҄v�8y�A�p�/ |D4!��^#d��l��χ�9�m $E�Y>'7�8t�'��@p �2�����A�[�Y{�E���{�=�O����͗D��ak���̨0�E��E��:���a�S"���=��Ώ2`�Pr��QKW����1ǻ}�&��������v�|lC�P ǜp�jgc$#2��&e �gP�';��m�o�9�'lz��.7�J'��@ A�A}�fa���A�9#�䀆�	�D˸�(�
���H�Yw!��\k�I;����Ţ����1K�������M�ˢ�}k�Sa�]��dE��W!b�v/��I��ňb�7���#�s֎��z�� ����e���,3)�J@׳�%{���Gt�=!�����x��.o'�\:M^�9�A\�P"���ѹQ7�\����� Ze8 �d�	�w���!z=�c�+��B8gr퓳����`A�A�4�P �(�T�P�����@�AB��K��WQ)(jٝn*Ph�+qA�3[ mg���~u}�<��V@�&}�'��򁫽~�S.��6P~b3�0nE��A���B 6�Vy�GKL(fS��"\ Ay@n��~�Ԕ_>3qj�p��>��&k{u,��4y�F�B�!{���l�ͦ*=��b
X��&pjӂ!�{!�yNL��b��(I"�m
��?xJ�j�����J��[AA����/�t��8���wHYy����X��������Oz��e��#-۴o:����T���ػ4�{+���hý���m\u-���好a��6�a�.��� IK����G_�1�r��XcE39W����@��A��I���i�͆�Z��Ii��՚V�jǁ�<���Dgd���d/a�l���?o�e'��~�<�q5&+ս��x�vh��3[�^�m��]�%�*�&��BdʀZe8�8]����D�������2���c�҆,���n�f���o�A�(��":%�y2{���W9��\A�;N�S/���r����2lt��2��A.7GVMx!� �骛��f�wN�����IAx��%�E�@���!�cV
b���* �A $��և���+�9�C�ZxH�A،齳��g�ehpe8P ̸r&`p5z���|GuX9�����FV�W0,	�9HFaKe���Z��{���G���=�\@Y���ʘ�o��[
��Fm*����@�+�jʝ�}�ɽ�)�J^�[�l5���nX�,C��A����v��.$��v��[�į�aF�͎2��R��M�˗Q�`��U�ɕԗ�Ż�-8��#RQ���C�^gm�<cv�����vdѵc��1��WY�U�]����k���P�ŴD.%P�iJ��"��鳰[yZca�;:Պ�ҪZJ���8���]�*l12�I�6�r�6T��J�$eę{>?eTL�z�<Z�k"������RaU�
���s�la3��amT����꣛<��!����G�C���@�T�6"+�ʬ�ӯ4y �X�j8��-(��p��jH�fS�A�DE\��M�&�� }�
_p�����!��sO �iS�e�q�p�tmϫ���	ZeL��Hͅ2-�>��lD�����*�>���+��'-� fS�D�f����Wwýfe�&`C>�g��5�+.;���\:{�m�Q�#f��Ѳ�<�(	����4�#l����2Ȯ}琟�9<����T�4��WQ29���"�D��Ɋ���b%��ۀ�n6�Ri� ��U�`�b[�C�M9���oZ�([U�|M\�*�8�N��`�Y�e��������7W���E����V=*��dz�j��F%J�I]Qq�F��Ɍ����𮢞�l��lV��c.��J�/��V蝦���0c��}xF�=����gٝG}8ak�mmȻ$,�^��15�����u��ތF���'�J�[������g�2S3l�U,�XӠ��_{�/c[����U ;o)+��]�2���eJ�j  GO��hת����;2�T�4��-0�9��w�{�Σ����B@�5�/
���׻�~B^A	�W	�7V]���m2!Y.a1�eУk,fZ��{j�{Y�
��HX��R�����<t�t�x�����!�j�U )� �cz�������ɴ�cmmvB��]�e>kL�ݫ�F�����3��l��4��J��1U��o���?V����XV�%:*�DU$2��}mh�`�oy[9�-��'_`��ߥϵ7�(^��T�wF,�Uu���z(��Û��29T��|'���{e�)IIY2~��w~��pw��L���L�g:�EN��l5_��P��R�b���<t�4��k"EW;uf�j�j�ٻM�YH@7�z^9����8����ٰ�=k����|ٕ�3<�/6(ďo_�����߰`�-�&�J�U��`�,���]]r�n�^��2	���@L�T+�Vf��_i����ם����z�T��BZ�ija�R�+��v����O�1j$��t'=�I�gCN���1���=A��$I 3�r��b&Tʙ��Y��0=��3�űJǱ6F���I�^e7��G\��=3�ֆb�@�r_��m�⧂g�ézkVz#�X�����LUx�x��ݳC'|m��;��W�����.�soA����w���ڽ^�����=��[�Ƙ�1��y����&�t�*���T�*+��_d9��VO���}�:xe ������H���r�Q�GKf��"�E�m)���)��c���.�E#=	�����/M2�e�ul��F�fF�Z�g�M�ҭ.�ը7������c�'��#��۴R���ܕ�|6�z�c�y ��Lqǆ�vX�H#wu4m�&&`L��(ȩ=�`��L�(P�&`���;����9��Ų��2��c{8���Y4y�Ƀ����o<_pr�72=)�5H�+�÷��X����1�MQ2�ݭ�V�y�k��M��{xm��O�}�ܲյUUy��}	W)���"�蔔N^h4-q]z���>f�v�M��1��ߙ�77��u�.�Ժq@�d�����Qo�B�Ѷ�,X�e�:�Z�uܻ͍n�
�E�UUEYB�B�0�Ju��kp+�pb*3dlRX�#��7�ZL�ss�R�ZѢ��1����������[�!T���Q�b-�m��걚%�������2�,6e��,�n�#Vk���#���4[X�B^c�V^
m�TV�f�P�օ��v,�U��ԍ�,��
k��f��f��|���_ĸgn����n�c�F�ƽ��jJ�)h6:_
j�\s��"�\�J���M�=f	�ەE� x	<�h	k�j��J�I>��f;����恕���M�/7;��S(L��ѪhM�C�Bos�/�Oes��	�&��
����Q�T���t)�dm�v�ʙ̧\�w��uu�A�w���[�ӷ�;.7ҿs�u_�(	t�eb�U�?�=�q)4�3�C|O��Q��}�#�՝wW:��	8���[v�6�`ufV�Ys�;����7��|�>U�g��ѽ�?�+8�P�B	d���@��d�������ɦ�5#G�pK�At���X�����̩�[���9���;��>
�̍��aU�3��C=,m��.�%�R|w^��N8mÑ�p Oق���2,?q��P���Zy�f6�1�V�,�_(cYf}��6,�;,X����D��c|L�#,��#>�wV9�r7�=��Dn��������3皧AσɀM϶Z���#˾�Y3W!2�.�>���r݉;D\&���e�c2V����~��y�<�FK�[�Ǥ�V�)�b�.&L���u���<pj8�'2��.����p�
l�h����1p�Fd���aB�J�"!'w76նi�c�KK���6"w�rQ��"aDF@v �h�B�L�)�w[�A�#4f��¡y���w&j�Ŧ\L�F���EW]OD���_?e�����R7#Gm�N��{�LծŜ��S��~���W!�v���ww�A\�r ֫�\�� �����|�����s�5�^�^!wْ�:=�GI�w��h^!����4O>��j�Nj��9�t�*�V��;��S��S1?sɕ/��Ȳ�r����Z����j��-���N�A+/L9�+��η�Ρ�7dCɪ��Р�;{��m{7k�cuJ��%[���к���Ư������x^Ѥ��p��hft�1������۲tΜn\Vlx�m�Ǖ9��4^�,�;m��Z:�]�w����]�IU�[��:����kڋ5��ݳtѺծ���o�M� �&�/�sy��^�ɇ+7N_x��,�[���d���t7�n��lc�Z/��4���󘞔�h�9n���n��gOm�z�vM�]�]q�i�M^t�&�pNe,ך�@ؗ�v��SK�ӤZ�>4F1H_WY��gU�Y�۝$��tx�;f�jwwV��d)!&�f.�t+.wu��`���J��ʕ_V�({t"����UcyU����7���	��*�[�3�	7Zon>[��*���1�ص֪��VW�t!Q"�5Y��f�Mtջ��Y���O���M[�Ϋ�u �W�TL�ެ�����^noHv�c��$��UuZ��/2[��#�4^y]�X�ܥ|�S37�9]-G�ؗ�����m�v�N����}���U��^�ŪJ�'�n4)EҢA	U�e�ea�HP�Y'޻�R����Oǒ����(�/"z�K������T�M�|!���؋�Rf��
!!$IR�*�_]�;c�}q�x�ׯ_G�n�:|<YBBLP,�4���##!��!!�___]�c�q�q�^�}]�t�$�BH1o�"�=�4ǅ��M!$�����t��q�qǎ=z��}v�ӧ�	E�a	�"ŉM��W��de"S �d4�$Qdɦ$j��ƈ�4i�2l��&��Ȟ;\�ٺY,aD�,��H@���F2b��%��(�ā%##cBdă@�����H�#ñ�&BH�a$�&����0�%s��C)RF!��9EHB'�1�c���u,�.��aV��9C�1���2�Bg�a4̥�۳�/��h8�  Ne��8�u�,��i݋��A[覮Ȥ�V�^I��	����5<Y��v�q�Z��_�m�N���s�&!2�L�hWJ���m3�[,��YvWT!��))H�v�Bn�m�%��%��Щ����5�NS�d����X7Ǫ��s���������b�M�風l�|��BD�-3�(�ȏ6dG���V���_0���!��p�!^�#����OT�ړ�j�U^j����~�Nد�Ӿwf??i�9���w�? �����&P��Ϲ�Ol7�k�Ͷ�j�E�+���t���t�1�A�<<�`y��]\��҉WF].����z^t��~9��$���=���73���x���Pok��p<����6�n��.�Q���bž�����e�a0�Bg���;ȏI�U5����/��\�E�޴��Lǘ�G6O����Ub�r<C�PC�K3���RR˸�4���V.˻)���?o��C?�3�+�'y��4��z~�x�V||z���)"�/2��e�r�z"��Z-qC6MN��|f/�t��;e����ֿ�F��k�m�j�uP�0��l[�]�J(�����w˅�U�����LQ�k����B:�V��+��7^��:�=�r��V�;�54�T����N��Bo��U �)	�(U���z�aɾ^��<�{���l��a�͛�o�;%WRF1���/�1<�g�?�4��_I5��ga�#M�s�8j�V�W�L�v��=��y�'����y��,@��S��rj�A��/y䳫�B;
I@DFrJ���0�pԴh�Y�c�9��HB��i@�e�֙E]e&�%/�yht��j%p$\j��3R*�*�Rg�.8l&�VW.�d���-6�e����.�v�T+�v[tmm,T�4]j�ʮme�ȃmZ�&tԭl/&/5��V� 5�6�H;���hx��%�;W�v�V!%ݷ�ͧJ���ZdM���gN�[����41�l��m�YSlU���SD�u�HG��]�ڧ��Mv�SL���^w�;���*��3l��J�Cu	�"�� zXw<��؈@n�ij�m~���=�lS�����H�ʥ�M��g��g��/Ҧd��}}z��#}�"T��7U�׳��{���`[2f@y�8���h퇯G��fy�M�=5�7Tc�9޸Fa����J�i?}�6݆ۚp�i���7�+sD�Ok��v��ɪ��S3�8o����|����Ա��6����+����4LF���SR�F�(6j���1u�m��1��=�Վ��߽��k�K~J��s�j虜��`�7���'ա�2��$��N�&�r���W��h��Ȭ#(ӳ��бN�=y�6��u���Y��M��W^�0V��]��q�|����|�1b�y���7��{:���`̍k�9L�ܼ��.ϭ���U���UTUk��Y�	1]۪����?Q�\p�M)��7�!��w>xil,/ڛbg{��9]{���h=@��w�]����}I�[�T���"��=`xF>���8/�S��ћ�5������.�~x��6������Y֗�3����he�I�-ƹ��0F��If\ye�Y�l�hzP+:�^�S}Q�w�f��������=�׀cn�tL�L���O�n�҃�M�F=��g右3߳�x�׹�۪�~5\^�ម����H_��'�`ƫ��99�O����S�K�c^�G�ݛ��x�f>�w]��s�/&��]��mg��Q�C�EVz��T��ŋ-�V��]rrV�
�A��>_5��>y+�W�����v�J������{-y��_-��z5].�pظ�vpE�^/F�zV���u�����y��	YWY���~���Oڧ=�����8�rX��<ɡ�eVhA�������`k���QJ�Vl�U�XU�$-V��uE[Q����w��t�J�Bf�ҽ�âm��9��[ڟd�=I��Ƭv�B�4ʳ��[�3�3��R�V�]�k4�z���ƺ�f�<W�.Q;�4@L�j��@U^��{�Ժo!�$R^z�6�=�|�B�~�n�撃�i([o]i��|&��@L���V`��tV9����Z�{+�ҍ��j��,,Ml��@�~��o�]��}��c>�ΰw/+'��|k���N�:ڱ��6�:�a������֜�jW��:&R�ĤX"�����S{�و��zI9�a��AU�|a�D?D""?����\vX9��,[�?ɶ\e!��qT�PU(���E8�s�1�T��j���oݬm;8��`��v���G�uiZ)"olZi��/h������V�VYSU��y�����	�f|=)���v���>TB�>��''&��v�MT�W��M-�y�фn�JE��������~��r���^�c�#�s����B9�Bfg�%�y���ZϺF��T����cY�ƪqT��v�qcFX��ڶQW�vfwQz��|�s�D.�� �1�ڽ^퉇���jl��[E���j�&j��ej@HZ���j�������,ֹLoC@(	���G�i����=G �~�뉠�k�n�Z���e��`Ğ��|7y��)ak.	9��5�mL@�H�Xٲ�<��f��%�!�(� ,[�?|�ca/{b_&��\��!������t�"�RYF��Ml���a�J�Z�9��d͌�B��ֻ��Ǩ!4�Q�X�ԥ��+.���-���e�2宖�K��1z�%t��ay��m�ٖ���i0� +���k0�/�ѳj�9ڕ��\�U	���Ѱ�h��s�+��Z:/Q�ɫFuݨZ�v.���_�.[	���]P��iw��7��&��K���^����f�#D]f�0��k���e�P�w0bx���{�vsݠX�+}�W�ƣU�N��eu�B�pmG��v���+��p<��'_���t.�K�vK�{�TG?��{-��U]]_�����+k��UJe��M=Y�yx|���J�圞��ɛs^|ѹHq�2���N����LU3�&�v L���*�o�ޫ����˾+ț��i��U8�T@�B���`��C�m�{����k�":8F!v�P>k�s޹�%��i�#QF!@�[��S2�tU�GK�SM�6��j�xf�+h}?'���vzMT��zgw�{��זo3���!~���A����,�e71j��K^Ty����}���Hr�vAC���pj����>j*��T�l\�3F�+�<#Ԗ^����D�)�'$���b_C��bŋ~&	'#���e��/va*���5<[q�^]����o�j����M]��Y�	7.e9�������ݟO��.�3�{֢�l���?�"p���vfgޒ����H�-���^�����7N�f���������zө�>r�-|�j�(����~���E���3�Wxu�/C�Wq;U��㷥	i38�w����ċ�(�P��t�[�GL�V��tj]S@�4lm�:{Ғ�6'vٗv0&SV����N<s�=O���>m2�Z���Ri)�S��U:�6S�7����=y��R�8d.�2�$���"��Tf&2��n�C��'�}__�趮�7,1B�R�Bͻy���˱EV�K�n����._dGm��dW��v�Y7p����u��������}�ϊwN��þ"*�Iٯ�q�4�UI�e�产�C���;?,cT���S}z�7��GG�v-t���m��(L��ɦP�ݕ@�[���o���w9�!�L��c����	Y0rxd���;GXT�r�F�h��-�κ!5x�_C��O��gl��M2���a�k�W����1/�wɈ��$	Jeb*�L�éU��U!�����x�{=#5��
�~�z��﹞���3�k�&HU����$��~�n���N�)��LfP-3���S��qe��c����'ٮ5�k~a��=w�5�s1�����AYF�/6���N���U��]�Oq�@�2�//"��遛,�������5)J(:��Z�4�bŋ}]q�ɦSL��-&U�dk�⺧~^w�R�z��Q��z:84b5�-3�����+�tT��uo�g���|O�G��ܘ�E�5�#E��8�\��c��,J��D�x(�r�ę����V�4kn߮�ǻs���}T����j�%Č��Ht�v��,���L�:*rs��+;Fޓ	�k����Z��5S�-+S�)�S~}�>$��@]�&T11����#�چ-�0���U�|���c��ńz�*��-�����`B��m��p5k=R��o�9��4�� �G��x|�jn���h[U8��AW��U ��咢5������(��v�5��S2&q���3��DQ�L%H9��Mݩ�V=S�̷��w��oX�<��ot���\jP�>\�j��kyu���pU�"x��94�@��j����R�a+ST�I�+�*QՋR�ҫ5�����Nܜ�wc+c+��!�^�]d�����|a�xd:�$�-a�n��WiM�{1�m��{��>�=��c��1�9�)Nˬʊmp��=y2�CEdު۾vV��S���q`$[
��F�;.���\*��A��gH�f$Lv ��,冪�oI�I���z6�N҇���9���f@�bv9f0���}D]�	�Jf|nQ�w��7�� *�:�)Jn���0�zZ�x���)0t�s�Z�V�>9��fZ�e��a��f�ήYٺk.�������&����G6���׷�+7kr��w����a�#{�!rI`�������/M��}��vWU�����A''^ѫI^>�ӚB�X�S�`��z$c��z�iś��g^Fv�.���W�7Kof	/��ymJ|#�{�_Wvn��79�MfPY!fd���{����z:�2Z�"X�=x+�b��-�ķ�n�ˤr����v�	�&���/1r�z��Kf����9[�r��/'pB���v^����D���ԩn����݅��_nޝ}+7�P�#�	��{y\��8�oVv��<�u�uK�F�R���z*�K� �C�����[ʕa$�>��"��U]�ae>��akm^�B#��!B���	y�8�3� �ׯ^���o����^�sb%	�O}v��@!�Fx��C����8�z���}v�Ӧ���&�
h!
D�0n��E�FI��$�d�	����c�q�qǯ^�}]:t����!!�P�1����@II2���{�����8�=z����:t���I4�&d0���pّ5u� �s�(C �E�wa�$�z딄 SMDQ�&�&Q�f�bɨȐ�RI) ����A�B2��5롐����2IA2�d!���"1d�Wq���Te�,D���/-�)kˤH�Ʉ�&��#�رJ!CM��H��Ҍ6�DEF)1�/OW�חu��&�+ac��Dڵh*�&&X�ֻ�=cN�ך4�v�kZ"`M��N��͈����u�Y��r�um�lj엕�2eWFɱ(�L��5��K*�h�̯a��F���������L��R�̣(b���%HYM�bU1&J��2�T�b�:��uv�Z������еbX�ˮ���Ʀƫe�6��F9H`���L�,"gX:����4Źf��K*R��E1��s(b4�:GZ)Zl���f*����K7Q^�r�������Qs���T(��P��uDn3����EjLlЄ&ڲ-+��n����L�l�s�����Ypԩ�K�;K�3��.�#�`��"q`sZm,��^�t0�B��*G%��i�j�9��6�3�AYR����PM(�;�Y�������6Ռ5�25Gjˈ&��ls��7Е�KY�9�i��2�`�k �J\MRl�\1�5U�K�e��t���6]�dG&�f��u�UI���aup�<����\[F�EyB½�:j5!�m�X� �hp�[��]̘u��b��ق��HKm."`�A)3�Э�b*j\Zh��ķil�ńbe{Mr���S0X�X�ku*Z�Lu���cMMaA�an[�k��-�\���6Hܼ����s4.����+j�Z�ҳnv�ə�u2!����g�RVha��a7++�p��E,�[�f��B� E�Y�e�+��e�r172݃0il�������YBL�٨3VYQ��@��b�h��ka�kS$�t��<�����Y�1�2�Fk��"�]ےs,���Z����+�zzkbDn�`� X"�V-+a�F�f�6�YvZ�w.��F��&nm�Z�i���]���������[����ج�������j�.�a�nft*�����[8����]t]�5�H��n����/U-���7J;��|<{�e��ؼ�1
�Vi�0C�-�p�� .�Kt.�m�Af�sS1ET�3��!�,4���V�6Z��@,X�ѵ'����?�)⨞'�w��M1�5��fn��/TrŶf4	�e��X��2FiNt+sf3yvl���Al�8q�i\{ ]�*ٵ��+���ƙֶLe�˖�.ٖMձ/\u�.R�������D(]z�,��X��61؀��n�5ΆNn���5m6�� (�5t#�tq�6�v�b�9����y���Gur��YX��S���$�|��~-@u�e�S\�L8���*�3XKla���me�b�D�����7̳҄�Q���^*���{&,w����42s�@���+�ϙ��	4�
�:lم��>Șm��j
���=���}��T�N������l�;�l͆�W�����r�KU�)�O��:��᪰�M�z��3U	�Es�Z}A����Ɍ���[/xe����Mb�h�nP����O��m7Oĵ��{x.${�O�m�2K���=��*j��UL����x���S�@0\��B���PhFY��ة���4��	�wu�x���N&�;O/J2+=����<'o��g��Ny+���v�����/5y� &fh�=���R�V�Z�V�VN	
1�sw^,�E��/��=�O9Dmӫ&�����d�=�F�6)�]��K��<[���bžO��P�M��K�x��/�{&=���^�&e���Ϙ���᪐
fX��qKxlO��)=�#SϏx�Uų	��=33�KVwFB���zm��=���{��	��9yōbq+�U�w[��jhڨ+��j�4�!_p�}����^+5K�{":8o�e���Äf�E.тͪP@.��h�เ�Z̆"��1aʬ�i�+��@׈L�(L:>��~��$�Ճ��3��?{�wP��W�q\D�g�4�e�c���߶�]��N�j�gl����	����=>����Ԇ4SJ�	���}�O51���b����K��0�e2�R4��*�rc���E��o7�ݠ�C��jζ�����������,X�bY:PH"Q��V�j�~�C�|�}M� �����վ��*�gΑ��׮}SU��G�b�\�:�-3�BD��fX���UL�?�6�T{n�'Q#��m��o4�(�ڕA?�y(�d�\'��
�
��e��CPs���e��
��\٢[�0em��o��Pt��C�L��(>nn*Qxr�z2��j����!�ś�5S�!R��)32!�7�>	�Wq�5QN��p!�Zo8ֿ/N�}1���j�[��ܚfe4ϗ��e��Qi�ً����ͼ�ct�{vy��;L��O��K���F�n��c)5^u�U�ק��C�so�[��������^`4�l����Y9	pc��cZ{>��4ù6 �^����_��D�ηKU�s�1݌��Vi�!猩,l�r���&LX�B���ș�v]���]�\��G�+��P}��Y�_o%5^�9�=�.�>��ͪO=�{�Pvzh����F�I�k��sRgR*������`:g�*��Ju��p����©1Wس����s��pY�Ob<n��py怜bk��	�ge'�����L�>ovy�o2��^2sǯ���=(6�Y��WX����-ҚffL�FO;�z1�)��巡MO�֏G1g]g���ֱ>{�}|�^��n��U��s4�u����i���q'�^��2�ަ�m &P�@��-2ۨ���HX�3�^6sǯ��;���Й@K':����_u߱Ƃ՝p;�:��Eͫ�r�]�;.���rJ˔�T۲��մ4�R��l�{}��_/�N�EH%ͬX�o�&H����,�Cr����h�]��ñw0H�S��j�5ۊ�x	��l�4��am+���3����(^ �H5߾�`��Ύ��͡�X�ؒ˦�����e�j*42m�!a� ˮ�dr+���V֒���P1�@�3
7)�c-7\�L���4��X@�6���뮐��̪��\�c6ke�/l�31(m��h�U�^>�~}O6��v�|���j��Ȱꚨm�X�#%�x��
������6u5��B�L�v�˿�oeE���c�E��U)�f�w��q3굱QZjhx�H}==���}պ}�ۡY�9�{޾���(W*w��;�a�2߶4�b؋�g�]բ��ӈsCca@V �j�������vR���s��^�|��dA�2�@L���S��~���kz����O	{w���	z���&f`�w;N0�4���Bf�y��.��j����sz��ާ}i����U�'��~�ھT����ϝ��<�?m~V6�2�m+��J�vc�ču�!vz��v],�*f�(��~|��m��Ԁ,D���&��=g�+��N�묈~�{���p���	��**�o�o�+FW��B��ZQݎ��G�a���E`ט�{�9�6ƜV&�\���.��,��>�Z
i����_X6y�����w��|%UI��-��f6:��I���վ� V)��i�m/��ȏo!װ'H"��љ�O1����r�ʡ����_�ִ7��/i{Hɔ����y&��=qu�=�k�!�W$8;;�]q�=���r&㭓&B�f&SCL���K�}������!f߳>_~�zx�X��&�v��ݗ�"���K�e�q�#\M�X5Aɷ;J^���ˣ����%��6:.�y$�}�ϗ�2��0��s;��o�w�=!t�����y�ڼ�/ؚ��8�@;��
j������wQ׌�]7���^ۦ��ܽ1��P>�C6�k�ͻ�����iO3�j���G����˔�'���|_;�z�y�^M����#vЫ���b���MϾ�f�jR��j�"}ݫ�'4�B�A
�Q+��c��c��w���#��U���@&=.�>��7�����[��z���Є_�M��ޢ��v ]���<�����;5����kv���7ºV,^��~����z�o�s>&v���3�h��u��8,Q���	s-��]T�H�(lLU�����h���
�� ��m��J�M2�!wQK==�Ȗ̳�1���_5;�Yh7�sU8�M˸x{
8�7Py�0���#����ۑ��VُT$�WGt�e�41�L��e3ʄo*=�|~ ��y�k^2o������sf��ݦ�+�iW���W:�*�7�z�=���s>�VhޚA5�n��|��.�
�5mΨm�=�u����fw����V��Y�/�޺�y��j�xC���;�\4��Br�p�������ś:��d��L���8���S��)����Y򟾸�d�t�+�E������￞��B7�1��K�S)ILv�g\��΅���0��Ð���!<LN��0ʡ�<���Ա�&��x���>�k���;r37g�3ؚe�gZ��2�l̑�.ed>Wt�s6y�7s��~^�>NZ��I��,< 1��H2/X��Qw��\ng��>��ۅ��\Ϫ~�۞��:�nۯ��Y7��F�v� JAfVu-xً�O��m����� Bc4�;�ک�i��HE�j�"���F���m���쒯��y �� �P�fa���E\χ�l�u�R�I�);6��ά��߳�+�w�6�f��N���𯺲o��P��������݁~TAX��,X�b�Gn�>k֦F]�ez��t�ܨ�	[�MDW��6�C:�6V�i���[]R��)K���+v P�$&-۩�#��L�A�R�Y��؈�1���=���΍����lh��7cX�R��I`]�'��Υ0�5�/c�2�ӂ�+r�p�&���r;V����T�T�c2�d�^���fY�ořUP��ʵEb��UX�����b�fA�����QLP��8J��~�|�}i=ߞ�o���4������U�z�ƹ�s�l��~о������~��^�����]���[s�Z��_=�v7�glHUv�^���g�&�n�I���Rbҹ�VO.Q}�6A�S�%_�΍c�sA��	�Ze�j�չ.f��,ۯ�2�6N�l��]]�3�S陻gK�4��\}�/�1.����_��:�''��ş}��D�tZ%��Bg ��f��=di���x�o<1#Q�����0`�%�1�*6Q��{x=��w�����Pl
5���w�*^	�s�\U�z�����֪v���.O�.!�k�"6d��7+/�8�mV��8P9�z,J|e�M�\�ҷU�1�n�n�1=�U�u��@��>:c�k��g<�[g��1u�ڦy�P�M2O���cn��z��GQ��a��]N���+����S��ٖ�OsE�w3e	��1Sdm	{X��-Ce=B�Tk#��zE�V4IY�.��]���f[U=R����w����F�y�Tf�ً���j��\�m�KE$*;�Vw�.e��Z�-��f_�|?�O�srle��5�p���Tj�i�*���m�q*
 �Lb���v���}j����?d�o��ݢ�/�w]��S�ݲ !���cT�&y�2�K���\gg_�a�3	�u��I���TVX;�S2/EBm�3�&0�.�1o<�Ce�j��M�hh��k���}�^�����&�p�[Nt�-SMZ5C&w�𙋥���y�Qk�V��I������~��h>�^��F�uTzu��iq���72���eQ���r�w��9���k#�t���Y�i!Y8��.����A�i=�kw9�ѳ9*�:�9H��B��EG!緧��9i��u�t�m���vu��j����]�[us�{!qRSN�h�
��t�6Е�j�����y�>����h��)��8ni�~g�;|˫v�s9I6�0��.S�\�;�hQ���57*��#�ſ{�Y�N�V/wc̤5�=��O�[6�ն�Ѕ ��������&�P�R���#uCh��)��t:'�Y�K�&򫃪�Uw�%�R7�Q��������k�o��r�a�:�e��xּ��}`�=��-�V��!s�c��[���_;�j�:���ڦ/z�z�ﭴ뷌��f�v��Yj��s0$2���U1�t�
)�F/GL�JX򱵡m�9��.����Ҹ�Ś���]yw�� �2��կw��
�_{�ž���W���Iܩ����t	N���pCN��6V�뢰=��8ՇQ�ZW50�]n,T��T��*=�g�vq���}s��k�xCi����'M{�ب��H-4J&R�*�"����ڢp� I�n�����~?wѾ���/���N!	�a� ��lD���&�$����������8�8��ׯ��t�ӧG��^l2� ,%�%g�k��D4�hЁ���n�n8�8�^�z������o[�yl1
(�c36D�&"",TD l����^����ۡێ8�8�ׯ^���iӧO��"h�1|7M)*_=�E��фe����6�L5D�b(�Ԓ%!��ccb#���'� �h�b���M����j0"��sk�� �m��@Wwb6��Qb,�F�1A�dF�	Bi61M���b����c�*J̒�q	Q�K�r̋ys,�(�m��k"�gY�ATX!|�̂H�,�$AcFw������S3*�����;�J�,��L]G�7T�4���,�f@��2�g�׶��Ң�]���&�2vvO��E�?�_sz���Oϕ��+zn������Pg����y�9��٧�\��
��|�fH7�\ Zz�L�T6y����{/����jF��ٖ؍&�YF��J-j���4t��h�.� �����f �B���׺>���<(�>�Bܱ;�2�T�ﺲ�n7�[b�g�:+�նogp�A��n'=&L���l��g�]���3�8��H�>��/&�L����s���U �ep�;�w��`9��!���lJ~�kڨ|ᾞoJkh���!��<َ���0_Y��t�\#��xA���}�]*��i�:vCw��*L(��2��2��/��b�2c	P�L�t9���,ū8t&�)�%��khj��#�`����Vq��۵��{ּ�en��a30a`���{���学�������H�]Pj ;%����L�.	C��s�å?b	�&yKPٱ�b;o���^�h�sU{eVz��ڽ*e2�e]�zǼ`���N�f�.<c}�����\�H����������DcPƩ�?;�x��~Â������J��٣^����n�h�o1�z�e3�U{^|����&�S+�����Ƶ�E@��
�l���Ƕ��az�Pv��C	�y����z���W��ش]�����Ø�)j(Uw���AC����c�pS�{��Yuv�Q�����hL���wE�CL��9z��v��bk�tK�Wj_���	$�g�y�,X�=چⸯV��z�+���[R��Z�`��vn�B�+%�ܸ��M�6W67S$[T�l,�lĚ:�����͚�KU���h�eXvъ��Dt��%�4X�ƅn���fل�%6��E��FJGJH�խ���$5y�t�[f����IV. tRb�XQ	lp��e6�i��7�����B�I_nU����u��j{���֎�g���z+8@�C�!~F�4�����g�0�h�[cZ��B�ľkw����7�������jg�^��߆d�j�EX�v(=!r��S0�2���u�j3�*!E�&�b49=�-~P/u�]����6��`��Tthv�}�ɇ�j���HUV�Z�ٖ�\͟O�p���7�ޘg/12�%�O3��@�4�f̱g�;��oӗP3;{Zuŭ/1ԡ���	�3�yHL�;�+E�k�m`ǌ�Z��^痛��RaU,���k�y�.qQBt��<p�j���garYB5RWBWU�Ĺ��-ro=����}�?~�m^�0��z�yGp�wxo����.X���e4�f�O2��1�n5�[��y����UV��c�Wl��WĢ�ݮgq�μ������cTt�7�*t�k7���Og9�^ݢP�,���ŋ,@~�&ܤ)�����8[�e��ؾ�R9���G�<���q��^��%	1�?�s��W�J�YY|������úf9��Z���Q�|#��BznT�<�O�cE��[�}=2��n�J~�Q�x���u��	(H&{t��m!ם����cgs{m�2�L�svrz�<:��B	��E@0��D"���dM\�.V��q@K�q��a����BqL��1�i������y�z'af㍈�K|����v,���S6p�6&2�)��.iz��e�h��~��[��+�Y���A=~���N���c3ċ��xJ�y踷p�K���Bnh�W�C���Y�L�v^K��my�t]�[Y�{��J�sk���]NZ0�R\�~>>>>;��n���+�	C�mU�[YU2�zX�-�2�L��W�:��e���6�9��nWg��0��6Jw�;(m��S�/���@�m��n��lG/�/�?Q���m4��=g����<�J�S(�=�vIS-��?>_-���s�-�Q+0�u��u�l�$���\ͭZ�� Ҡ܋
V����e�Pmy���S�}�Ye�r�c�=}7�ǅ/fL̴�eq����d�����ȷv�r��=�8�|��%��UWT�xj�1sT��w@7κ�����p��<�-|�.o_�D�(�&Qi�|;��l�v6f�3#�v��,��*�fu��,����x�૶��ۼ�����W9��C�*�s#Tr�y�*X�Mx�S�����*��[3�;;�A#�-Q��12¼~&�{zc��y(���7�>'/�z��1�j��+�gtG1�sF�!bg�Ri�����=�n�n��gYlؕ��P�y�.^��������IY�m,G�������)
"? �G���yU.cT���O�p�skxf�S���������ꪙ�3,��,z{�< ��]�q�n�{�k��ӌξ�4�E�W(����V]:��;�R�S<�ݮ��i��m�n�N>�I!�`�Ø�A��NX���v�sĜ����YS���2i�����M�,�#҇&-�݌��r���W.�?�_U3�N�&�+v�.�L^�Nt]��͏>�ӌήl�ۓ3�gJ�>ko[Ǯ'�4�˯A'�5+z�>���N����ח;RU{c{p�ӂȿI(�`U�]x�O�,�U�����h�>�u*)�ρ�1�b��{K��V;���~���tl����u#@^�W.�:�Gb����ݡ���"�-Z�Jk�R�*��Y�؄t2˄t��cFZ�����eЙ��ul�@.F+I� ��i�M�«
Kybc!@DKL�%���s���B�A�V���5̦8�b��@Mn�ܬ����;U�^�d͆k��k�*��������.���&*ηQ`��װ����
�/�}�[��^�`5�,�0N����.љ[�Zd��B�<CÃ�S���. �M2��Sw�D&�b�CW�y]�P�I�ܽ���������fi�`��/*�u6h~��F��n�oa��T�Q	�ƺ������#5�	�S	�2�4�{��c=�Hͮ��N?dӌ�x{qL�2��˻�w��}�u	�&Wl�Y�nx��l�cU��i�Jn��M�Y4�M2�j����)�Sz�c�GQ���wa�k�qS)�2IXj���I�%BgN�@N�1��V]v�a�Yc*sRPC�/	C���lɘʧ�����4�3�v�׽g��b/��cT�RHwj�1�����j���	TC/^��A�j��C�J��m�I�{s��=���_C�=$�\3&�Ԏ�:]�}7�ŋ� fd`oM{����_^�3�3�CF�O_���(o:ُ����y���_��X�Ao�K��յ>�9��\�Տ�TϽ��L�lv��$���%�����]>��[�N3=�z�
ܨ�]�q:ާl���7����@U!3o��� �����o��ƌU�|��;�L�D���tz�%k��w�H�0�8t*�vV�A�K���#�m6�P3�J1����N�����m޻�j�����#���U�14�1����<Y�aN &}0Ŧ\����k��i���;�����T�3����>��F��)�j.���MӰ��1�N�H
������V�k��˖��E����b�e��ҴЙa?IIwl5�Z��&^(��aS�͔���ojf����}����%��[��}t�1�P�p�U]��C�zv�yb��[n�j��B��U39׶S�.g�r@�5H�yK_�+�5[k)�\[BW͒�e4�i�g9l��+g�+�s��{T�an��	�;U!3U[ldߙ�4=%�/D	��q��6�m*��,`i{fZk
J��]e��	���J3��D��1�S⇥�	ʍ���;|��W���Ex%n|��e�%�\e�*�SU8�>�x�ɸ�}��<��
��Ws��pI�a�eR���&���>B�v�-��~^�B��*��8u�z���x���B\��^s��I�|�Y�1!v��n���{��{��{+�ژ�Cjsϫ�9��b���<&\�xw��X����=�W��
�<��fc��&�fx��i�FJy�]���:�_��� IU>���,F���M�M�n��BAO8�+2��Z��,��np�|Ջ�7���T�p�=��@�Η;[�z��`[.4��z�]c�)A��b�\H�!�S�\U@��qy�����o�(fWpz�Ӱu�[j=�32�}��	�h葶�<��ceWS��s�П�3y�u�eUo���)7�3�5Ri�g�̈M��"Q�>����E���w\�I�P�L��A����9��>R�q}���~�{.3+��څZ�q��✱�32��K8�Ч]wؾ�>��ś��+U�w�>�C��7�������S�i�T��( *��
*?�������(,����u�MP� ����2�e�5-��2�K�K5�+i�����fڙ��ͭ1��R�X�Tʩe�2YZ�,���ZejXͭ�2fژ�mT��TŚ�6�Z�Z̵�����MKk,f�55����R�55�������jm������jmi�����ԭMJ����ԵMM�jmSR�jrڻR�jmSSj��T�����SR�5-���MM�jm��U55��mM��MKjjV���56٩Z����ڦ�ښ�Sk6��mMM�jmSR�5+SR�56��mMKjmejjmSR�56��Z�����SR�jkSR�6�j���Ԫ����ڦ�TԶ���5+SR�o{O�P" �E$�MM�jm�Sj����(F��B ��D$�hB
+<�hB� �B(+"��B +t�R��B"+ ��B(+ "�B
+ "�B+""�B
+w`���"��B �"��B+"��B+"��B(�"�H�
+ �B l����
����
��������]������ �m��ԵT�-��Z��TԵMJ��[u�5*��jjU���56��6���"�����j�����R��jX͵5*�R֚�Zjj�u���՘�֚��Զ�-,�Le�5��ke�6�B ��`���P�������QU$AAQ�  �O��W���O��߸����#�������C���(�@~k�����?�������~��?�������?����DTE����������4x p�i�"����>��C��_��C��P��촋_�ޜ��P��N�~�?@��C�JEv�ڛlڦ�Z�T�E�Z��6�UJ�Tեjm�U)��Զ��V��ԭ��jͪT�M�V�*�m-�����Ԧ�6Ҫf�+M�Vj�m�6�i�F�)����M6�$(*"�
,��)��+j�j��Zդ����%Z��I�ImJV�j�5�f�4�RͪZZҦ�%�j���ڥSj���"� � j��!(?��l�S��@P E$�����/�����>��>W��~����H( *�U���y����ҋ��٤����a�������p??T��0��9D_�����(~$?�>��t�QQ_p~C~�Ap?��%�x������+�I���&������4�Y��c��~(���� *�A�~P�?3�>�~�����~!���O���� �Р����?@�?� ���<�x~͡��?��N~ K������g���>'z�Rw�� ������VI#��IH�<���q~?I��ޢ*"�C���[4"*"���6՟[��!����(+$�k#��� �CK0
 ��d��A���                  @              @   � �DU@I@Q@�)D� QQ( P
�P$  U� H AB*P*�� *�UIE%EU}� �(IJ�����P�	)JT��H�*��%TP�*�J�!HQ�B��**�  �"DR �D�H��V���j�N���;tW�����9�
�tN�u�M
x�����J���R�=9�T�z {�罃m���J�J�� o� S�A���AA^#O�zt ����x@}V�q|�=h)��Bzҭ����yi�ԪU�#^���.�Jq@����YV���P
� /�(B�"�EU$DHT����eN�U��];��P���R�N<�8���չ�S�\M ��v�J�nЛ�=i��t{`s��{�((D��+���űɥ�}�I�QJ7gAW�o{Ήz��P=��`:���%R��ꕹ��үz�אӜ�U2�继�J�* o�{�
J�%EU ����C�1�w�-�R�aң��Jn�S���p����n�;�*' 6΀��UU I/| .@<G��$� 2f������. ZΨA�[�T��I! U(| ުQUUTTJ���EQx ��v���݀���S � }��7� f `r*� -�T ��p@��  ��{ =B�� �t d@��C  39DC�l9 7`q݀C� �@$)U�   ��UH�ED��EURG�f ف���� nR�W �t d b 47` �H @@`	PR�$x   � 6 �U� �=H�`:�C� 1�QU\ Ðu��u��y�|�O@d��F�di�M��bJJ�z�24 4�j�	*P��R%#M`��)B~�@  3PI���R� ��?��������rI&����G;a�(���QYF�>�����!$���$���m���v�խ���[V�ߖ�ڡ$aHHw����Jm���_�p�m����ǅG�ι��[g$:�p�p^�ᡬ�y@�����ʒ�ۏ_[���%O^�R�I�����,�� A>��K����od<<yu�!��.���. �S��b����&E3[�.$Q��命�˵cXr���ov䲇��1I�Q�^�7^�v�7���.qނ��t�hq�ɢ����+��Ǐ�wɭ+�٢��9F�fӻ���"�4w^�8��ڳx��-�m�I��j8���6n[�'�]h��bˋ(=g.&�v�3���Mע^熠T��5�p�8�7�R�C�Cv��E�q>Z��@�l���f��<���7&�vSg�y��,��p�Oo-7N���!θ�4�6I��Tr�ٳw4��9��	���qb�]��f�#=2j(w�4��	��h��A��ۑ�1rP��rv/�%��&��ܨypӦ���l9��M��/I'],-��]��Z'(�AK8��T�xC�i�Jۨ�\4t���|�IR��ז�wi<�q��e��v��ˎ"PJ����^���G@�2r�	�����P�<7������ĳ�IB9�^wL}��73�\��h���So���|V�E����e���\�*�=���ٳ���{4G���������c�%<m&�,I�i�uv�7om5�;�����.#��`�:t�ظ��[֜[4����X˧���)n�ۆ�X��7`��%[!�뷾�f���u�'�J9���ځ��^�v��=<�Ӓp}�s�+�>z���gL��'�Lyb�/<��������7�2D.�3�H2�������$���"j�[�`hLfD�:�UѯOoQvd;�Yu���t+Q.=�<ν�H�B�e}O$�1�2lm`�*>�<�?�c�pZ)#F^i}���ns[�L5���%�`�>�c���F�yú�e ��΄n&X�rWue���w�XX�_��]��V��9�^�`N�"��p�F)�������y�Fޓ�/���8���\�x��]��&��]�����ˬ�����|��W!˒1�;���x53r)�+����^��_$�����je9װnIک�R26��k�\�fl�IɷJ�R\N����}��bp���ni}pI�-��z;���I˚�^�:w+�̪X�EG\g��/:�l�/P8��׫N���X/M�,�9��Һob�f���qs����� �[��w�"wAT��^h=����˒vRE�ZI�#ӹrC��W_6��m���MM���N� ���b�S�Bu`�&�mln�Eil�_P�Qp����+"`>�,q޸������/;
�"����v����~��I��v��z��nq|�)��s��/�o��<��::؜�+b�ɸ�4���K*�Q3;+{_e�tS��Hy��M�;pɚ)��c0:�롶�3L����-GVcpt�wwi��U�:r�=;�#��H���v��[�e�x�<�tLlM���^��65�@�&M�9n�u��њՀk
���$͸:��$%ig��T��9���\ط�p{�s�	��{v��q�� ��H�~D��BQ��K�1n`�2Zś���b���Ӈͳ��:�n�Z��Y�BuK��d�{ �0��M6^�tӺ(G���B��XI[�������L��R��p�xnn,X�j�x]ɐ�E)�6ݮA�M�x�sO�����Y�=�����f�1Ge7��X�c�$,O�N,�ɍI�an�=�^� `��ɗ���;��0��r����2X �xLO�onJH}�U�:ۣ6�����c	U�Ԅʹ��k�'7û##����Һ.{��!�R�8#v<�v �\�T�CBP�sSЯ���I��&C�������j;�~�:�C�s��T������Ds�K��5��ӏM-?�#,�1�-T��qܑ)���Y�~�����$���#Vi�ƾ�6i�;�v���XSFDƻ�LC ��ww`��8tQ�sMFS��̀�/{h�{�*a��vt��5Cu=Bs�*��X�!���R]ͯzh����rs�ߗ\=����٫����e���	�ʴۮҔ�+,7�q]�1q#�#��L�E�I��V^�9��'���qL�ս�eY�!���f�ʪ���yj�ޟv!��r|�}Յ�c�Vp� �h��î��1��o!&��әtd��N�]��j:Lӭ�5x&8:����*Ɛ{�ᓾټ
�
ït����1D�λ���;]*ѯE�%}�gFYӺ#�k=8ao7N��=�����w��-[ ��M���a�wQ��䋔n1��#4J$�k�!�Hc�f-��mCP��vi��ٺ�Z�y� n�u���Oa�M�j\`:��F���;&���5S���⛼�{�3�4B��,T��ӊ��,yY�^)&�9�4��B�\��3�v���n&h,��ݟ'\��Ή��"{j���ط+/�k�A���!�L���!��c��]�*|��aZB�f�ܯSTn�vd�c�A}�h�,�Gti;Vr �]Z��x��ܡ��M�� )���ZR�nT(�f3�1�:��4�2h/b)��[B�^�Ч�-�.N�Z��0��7&vޏ5���>��p�ce��7 :�Ҡ�9`���Hݤr��r��Fw���ɂsٻ�q���&Efwm�� g���ж�"��}����w�f�k��g���������W��]��!��Ml��ނ	�sp!�
٣!��{Rb����&;���u3&����I���6_N��tz����Օm�{�r��Ov������^��䤈!9�y��^�ߣ�N�2�p�����wP`��S�7K����g�����S��4�JNb@59^���� �3�b=E�V��
3S��13�ɨQ<�ː���MDFC��8[�������<jŨ�t�MFGĽ7O1��ٔ#��Հ6��c,#�qU,+t��6%�Hp�G�w��nё�ٽIz5*�}���>&��<P5L M��ah��}5��{�iكJʺ�}8�Ծ� $_qK�0B5M!�H�{�I9�e#凁�v����/����E���{7cx �83�N#�`�-�N���$�r�� &Ħ����0i��槖"8�G��WF�-Ӷ\7�Io<�S����w�@�A�"�VE.[�J�ݲ��T�EU+���v-e�B���T���`���z�ef�0�DK�1�/Xx�uA�s��yFu��u%gB�n:�oNI9�$��؊�8��'���j���Ŕ�8�;�K3���B��V�9L��5~K_�ݝ��i<(��1ّ��v�l�M�9`[�g�>�;"��K&.�y��ta��7�_��^85�E<2�ޝz�����0�ս�rv�L��v��R'J=���-��eVlS�;�}�aQ�i�G(ޥ��t8$�LE��h��Äi�����\ِ����s�A��
�gqA������_=��;��^H�I��t	;�gov�u	\k��D<ףz+��|�Jϗ�&^{U���_���Yn���p���kŸ{��pr�w7����ɍ��*ݻOC�r��P{��'����,(��pC&�e��[7:�d�{h� ���iD��⹼[��� �.v�։2�	I����ﷵiA�]��*9x�З9���ʴA1qƶ7�wu���N@��8�3q���{4j�5�m	�R�Ã�����������f�����.St��[ݕ$�? ){���6��k�NLs�u�.X.�7a�'���\�����0������뛴F{������ǵo Ċ\�����gsK&V4������5�m���R=Fv�j����{�D[2�&��6�''Mh"[��L6�P�)��"<x	�RH�˹����}U����9ôo4���	�3r��6w*��j&�ͥ(���:�Ϙ��,JQ���Z�+�1����9oɀ�:�՜�,�ÂǊ�=���W*��58:vu�7Vn�on���ǝG#}ݯu����{�k3�]�33Gwa��Ýw��9��o#�}�"V�=6�{���=��N�>/��=�3�ܡ\bu����wwL�?$|�s�r0e�ñ%�R��^�@��90z��X�T`8U�;��f�%�Z��!�:�3����.��A��Ժ�)ڨ�^��6�.n�:v���f=L���]���F(�<�"��ԫis��W8gs��Ґ�ƈ<ð�ø:M6n���Ʃ��}� FvJK���)y�ɚtfÄ��s����-��������t������-qn�aƠ�q˼c��AA�9۪����_*�Cf����k(��U����]�������+��M��㺻`U�
=�$���>ղ�'�i±��nwd�{9]�Z]n�vI����а�-�o�ɮ�q peQ�ٹrf]��g��y��=����J���l�w0��\�����;zU�n�ZL؂�:,��x��ٹ�$���[�ν��!C���r۱�[6v�!̋v�d��d������,��i�h��h��Q�C���Em������-k�݆���l��ӗ��[����]y�������(���#��b���d�.����w+���#��Ős��c��#]�r>��������˨W.温��At�f�ks�9�O`9)�O�9I1��g,p��fT�v.Ӛ���ؘY����%���{��S�e�ݮ6G��uȔ:�T�Y��:ou�s���^F����+�2p�`�4v5������p@�*o`��T�Ƭ��v��@l��pMEH�+�5�y�d�+�Ѻ�q�T){;��uCѹ��n��aBB��ܫ��yq�����Cw��TO��Xv���F�+y�h)�*ٝڅ�KG7��aLVN��x�]ڞ���8����=�-ǋ�|^\L��)s����fc���{.t�tݻG:�nݒ�ru����X6��|;wH�ɱ��.!-�x�a\fGPQU�]M=�:�'�CָƧl�A��5�l�:*��9�h�Z��vtF�z;���g$�;� b�u:.V<>K9vL���f�$û�w0we��X�l+H�sj�zٝ��P?��Q���&,��7�h.����g%e\u�t c|�\���N��v�N�Ń��G!����YF�;<u��b�D�W;FX�RRh|$w�8M�����1���ٷ�¤�쳻b+���ZvӲ;��6������!����Zl٠g}���ȇws�X��1b����2J��#I�M�W��,[_e��;5�Z=5��;UX�j�v�m���:	���%뼀o��������{�CPM� 9sO>c���v�v%���ݧ�����z ��R�T��'vU�!,<�`��/@�k�>���]Z¦��Y�_�*�Zo�qN����ݑ��>��QA-3�cD�=æ2�J�h:��]�/V�O
���j��Ω!�z���OrA� a����O�~m*����p8�F�:�+�|n}���{�����
qf��=pLR�a�oq׋�o�oU-p7	��,�]E�L��ٔ�����㒼.8��8qSi8�:n�V�R�;������.�֘��z���]�j3����nH�����a�h�ۼ;����&��w�h���K���Z�!]�3����p2��`av���{�Ib`�õYAxU�2��{���ZVF�2��f���݉��N��՜I�w&���)lL�K2�x��1	2a��)�ݻ>�@I���H}΢�u.�5l2"Z�yɻ�^��ko�ߓdl30�3��1�s���4~$�4n��̖_�3*`FZ�P��|���=`�T��#B�Ѕ�
IN��EpY���ڊ8vQ��Ś���t�܌�z��FAI."�F��of�/6h��9o[��ߗ>'qpd߬��92�%=j�Èr�!x��owb�&}�}���ݔ�֬��R���7pG�B.������LgcU+19�4��ǲ���d����y��6�=q,q��ë́����
�}��h��㨅��Xh������רm��D�ױE���f�'t;.���HPeǋ� ���|��nv�>�k3��@�WZ6�3͚:��5.'��×4#�2n^�͌�xRň�/��M�0�lQb9>`;��}�%�qt���G.�ڌb�0ܡ��Be�(�Xfn���=���AÆe�g3�7"�c�.��i֮�څ�n��wf�?L���p��d3oiԪ�WGw*���F'sN����>��bT�)��kT�ŹZE���J�yJ�#��ʶ�hNƭ��n����3z�R2�9{IvB��&P�;�!gGn�x�R�#s�I7���*���t�������xm�uV���ޝ3L�;���*�n8�L���q���斀��fB���c1��h��wzG[dj��0y��3�0p=	T�m�*wN���'��[��&.���٫�.�]��y�L��YAÛ��qڑ�_M�{v#���Rq�5���ڦ�N-
�E��HX��Z.K�h�q�����u�)�� �F7sGLZ>M]���! P$"�B+k����ѫh�����TUF����5�lZ�h�F��Ūŭh5��[cUcV�U����E�kF�UE�U�j��U��[حQV�[EV�U�jգ[mQQj�lm��ըګF��V�[lV����6�QUX���T��[Q�RkEmlm�m�5[F�U�[�6�bբ�X��ƪ�Z-F��k�V�ڭE�lmj�V�*�%mE��6�lV��cTmX�5�Q��V�mb�ՋcZ�4T[U��V�b�[j*�V���QkW�֭m��������������_߄��zz`���c*�j��寡�f&�����	�1�E�b�~OPܣ�3q��~[�W�~7U�~f����5v{4{{�R-+z�(����8TXy3KʦY�Z���d�&��f�c/=������G��q#���簾I��[�7=��lf�";寱��� ^�ꁼT��^e%�7��~so����͠�ݕ�|GVz���d�i���@����u��.��<Ҿ���3��=�ݪ�y&d6�G�V��wT�cUM��Z��F��:Fl�����X�c3F.��&�q�)��ܬ{��=�ڽM��w5�A�����4u#�7@�M����r�ӊ�W�3Jp�n�8�u�\Մ�MF8��H6%ʙ�H]K�Qyne1;��К̀��X�'d�AT�9:�2k=�j�K�fN��<�s�˯8Bn`����Y����5�Mtڈ7`�b��0\�"��Ӝ�&z�{�� ��U���:^�ɤ�N-�[���G�.`��z/K�p�Ӻ��smH�"��� 9[��y��"�z�i��/ y{|�nD�3�gr�ܙ�Ri��:�p������h&�o���d�5?	$�K����x��W#btbd%�/��a{��$T�u��p���ȷrn
�[��ә�Z��ٛ�s���(��v[�º�T)�X��~��J�`Nz�8�ː�VM��~�t�Z��]�a����v��!�6��]�l�]�[f�2���i_Ob�`����e艼�qYvK�4 *�Q�I����ZcRd%m~~HJ�<��/&s�3�-�.�w�s�m�X5k�8^�wt	n���p���G�P�=O��+�����K^������ٸL��΀(랆�}�j���e<d�nNX��"Y�p=p���M�0�N�[�I��6��2(�,}W���j-2�K7QQ�;��1*�H#*��=�NG��Co�����O�.�=���t4v4Ь�47�}�����d��i���7{t{�bc��֦�Ր�^j����`��V�U5x�!
�܎��<'n�����|�S�ͼjo��//xt�z{��ݪuH���iHc�G�'��ۀ{Uےf�wH��Ǻ�������ǻ�����ܹ�W�;�F������t���jF�d�,�7n��j����f�G�D3��,���Q� ��ut�PgU���H\����ɗӌ�M�9��ַ}�I�ʶ]�,ټ8}�*��$�`�*����-�|��c�^�Pʡ�&{�2ų�cjg������L�#o�
�5k|w�{nk�wX��{��H�M�����ؚZ�cz�f���+5,�š��*U�67�pP��׾�3�0��fqX|��k\9{a��p��`�U��{8v���U:�P��m �+�h8z���j�Q��&�j�+�U��xyvt=�S���m�!�*����]�g�& ��-���|@�9Vn�Na���@��X']��T�[v#m;3����*����ad{n�Dh9{&x]Z���yV��~άh�9���4�L��8��wX�7>��:sZ�n(Sޝ�KӶ��o��b¯/�>�y���nn)��Z'�l�'���";O����Xm�-�/Z��lc�ܩ�ۼz�KG�,^�d[0#ᗖ�d���X�(�2��R����a����(����仳�4���>#7aJlɣ��#_]�W�"CVn��8�n;��v�Q �=����/m�.ow�G��|5����UjW�}������!�b���p��*��A � ^�tr3n��i�>�E�� >K/D0o窈)��)�ڶj��+3t�J�Da��1g�=臌ò-ڻ�Ȏu]����o��	�]h�\�]�oWn���ܞK�W�do�g`�t����umP���i�*��/�vr[6��w���g�e�W�����k���	��4�V�P�v�ilk^S)�P��t&ē�[lm�n˺��9t�huj��T�D[zӚ�����C1*��=�4ƃ��J�t,�_^x��nw���Y���{t:ܽ�{��c'��,������<� �|"��p��4h�4�3у��93{���i'|��| �0��0B]��[�P�=Z��"r���k1M��%2K�"`Z�wp�@�;F&wa��ũ�5@���td+p)��w)�v�Y��_�z�>	�p[jp�ݡj�Ջ�v��nJ��M���q��i�s���N��ݸ��`<���R]��j�'���}�D������=�D�����`��[����e�y��eS/ D�W�<#��-�oV���;���1�- ��%�8�����T ^��<i�׊���{pҥ�x����&�� �sq=��"s���A)T�O���;�x��=0̙�[��ܦ�Xp^JƄ�1���Z�g���*�M�'�&���4���ަ��<���:v���R��ios{��}�JD�5{=篱�96<���-�T:і������ۛ�ڪ�L�0��K�S�U�{��zc{�0�tǗ������Q�f[㞰��JMػT>�����8���f9%��Rw6��N�՗g�Y�;��=}��ua�&���x�7-�/_ ���5��0����1S������`N���!��Ľ&,����]#����Rt笮G�={AG9K[M\��x�P��e��n��j�}��I�q �Un��^{ɮ��p�bc/ӈo&{����s���e[����)���?�ۅ������{ѿ�K�4ʊ�n��*�c}G��^z��a�=;��}Q!I� {�7=`Ϋ"e��6�8Iz�&!��'� �����V,d�Ys#u&���S՗5�b�f]�@��3�i��Z�X���f�h��ZQO�g���}7$��*_r��E���Q�� ǽ��*kd�j�_�zwv��=ݞz/���܏˵(}��3�2qzy����j�A�ݽ�ߧ����$�|蝯mH#;�yf����\!^����O^��&�CV?q���6?$�{˕��ܡL���%��n�$�;���:o������i�P�ؗ-�XJj tm��{~�thG6�ѩ86�)]U+^r��d�ĜV."�*	��ÛI�<,�4�����f�w�����i<�w�>�ż�@~*��n�i~��(��R��X����v�z��R��:/*�4�!�Bz�3A&���P�KΘ�W����+��@���ݑ{珦���f��^G���w�
��2D�^z�\sO-������8n�;w�nfK����Z٠q�}�}��;to3��Yi���~��54�ۖm��xQ,S;L/�(�H����)s.�wB�-]K�,Ø���'*]pb\�XTm_�i'j�8�EA�!ik�{�u�;o[�{��AH�!n��&>{s�����h��hʯ������|{�ȗ�O�/A:���&���)��2v>�d���6�uyGf�d�-/=��|�{�o'Nn��Q�ta/��L���JZ��Q��Ļ�z�l>�r{�gN�\Y�7�hT'����ocG4xx���|_$|k���n���;��sB��=f�Mi�ة�X'v��m�%^��jꇹAqv"�S��E.T#���f�=�"Z���aB�<z��i
swt��MG;�o_՘D��nz;�!�xp�)���_"w�f�y�:��	��[�9޹�zxj���^�u�ۈ��õb�}2_[T/G=F罭eޥr��B��F��a���͑}FW�;�=iXzw^�����՞�5?,4n�ߥC�W��Y[�/�y<g`��q�|�<R�*;N��o����ޯnӠV�m�Z�v"q�n�J]ӹI�L5{f��r�{��/��G�a�k���ۗP�A�#�e)�_a�����ŝ�,�(y��eM��~'#�Tw5
���Pb��E�̬!�b�JZ�8LE$����נ�"I\��YY[�E]<uC/1Ju�b�*��
	4bQĦ^ٸ9�]Q]�<��e���T�gb��n�N�Ks܎n�"Q���4"��� ֍{�w .��y��ةzV�a���.t�	p�]S�٬�J�]MeE�c�^���5y���O����3���B̈́a�L%�o ���P!(L��qwQT�Xe˛u��2Ҙ�2�Z� јC}�x�T\@d7$K��2�~���U��O�Z�E�p�y�E�||�af��j���c�
ˑ�结�w>^1�`���ۯj3ޛ�r�E�>ً�Cjc2؈�УO�n� ��Gh��B��6��&������<�Pp���+ױjB�jf͠������VsXY��==�f!37�+7E����	�&�c�t�d=��W-o�K�d�>���Ս�d>�܆q�_q�&�~սbț1l>G���T�=��b���|�-�Lk�ʰ�eX����u�,X��>�ɷ���wQ9�hd�(R/�XMx��V�x^���I�G/a���"=�<w;�� �ݺ�X�FN��� �ӑ���,��{�����WA���@4��O��Ҙפ�q<'ļ�,�$��7n�s�Cj����߼��Y��B4˔�zҪo��4X���������C��\�ws��.��Dqo�G�cI�ȯx��c6y���ox7�7�]�Z=�J��t���@9j@f�w�G�hOn/8�t�<w�����nV3p.z���֍�c��M����>�5{�0��s�����j �^)kl|�o	1�m�*wt�4p6��[�`壜`��~L��*�>����5P�h��F��"�&�zŔ}�wӱ:;hr夫�o9hy�L�k3j܂*��E8�d)3�5G�5x=������g5s|+!��u�0�у`�θ�4�!�����m���y�����A6w����v� [����tn�0�%�R������޾�k���x-�͡]RqIU�Н)����dL��Z���R7�3S�,�Z<��\�s�E�/�l����z����ҷf�[�4w�x�<��܏sހ�#�O���+���7G�D���;5�m��W��6W���R�4���W*'6b�y!�B�t��Z��ژ���3�MZ���gi�Shc��
��F�×�D��[��gn��n�<���O�P�*z��\;U��wI��X��tT���k.4�s�صS��#�����Ų5�X��^�����q�Lo�Y��T=1L$��4̞�����u�}^������	�G>��=wqf-�+Y��8a��66�^�u�����{�5���Cpc?K�`����O޻��N�۪�Ԩa(f`S3�̷.�����4w��Uj�1z����!��]�[���jX���#U�z�דBC���Z�������ۓ7ݐ�����,��{�8�x�� =�A����,�
�W6/#^X(���l�
�f�6!V�9����D��=~��>\�ȖN�MU��|��ˍI�U�y�����=���7ӽ�g,��Dhî���@�l��#)-Q��װ� 0�k�'�����ᵩ�yJg�gj�vf�Ԙ��c$������c/0bq�v���v��At�j�u�Q4d��q*�!�O�ׯ�8�|��^
R�3�7�G��O9�ܧB+�<�v�Bz�y�;sm�v�
E�/;7���~��	�4Ǖ��+@��g7�N�~��B�t����g�L�'��/��m��!ٯ4r� ���|�%��K6{}r.�,�Nԃ�P��Q���%�(f���q�N�H��װ���w�!�W�E��$Ŵ���t���3�е��+aB����#5l��a�j�K6�vc�v=]��<\jas���z��?g�����qo�~}���S����l	�o\�}��	�ٱ��x䂑4�kFn�	�m�M�6*�͸I~��ph �F{��{c5U�j_o�a�׹*g_cظ��1R�9�&^o�n��
z$�`�W��k���>��� �LK����-��u���Lo���ly	�gx[>S�S���=�R��A��������Ti��慧��b6���RE��in�F�uY�w*[��i�H��3ֲ�;��C{$VؚY��*���-����a��{9�ⶅ3}\��p��vx#��2u�ѵ�d�ƨ�tD��-�$��` ^2��������Ѻ�u�y@�B8�OK��`8�ٱr�η:����v+��'/i�e@q�u���۽2�x����}�t�o��g�����E��1>�����TSHK9��tk�E��[�yyx瞳�5]�]��n�S4�br��,�EF����Y`Q��ŗ��T3k�U�y�{۩�	T�̹W[��M@%v��PP/�s�"�ӂ�ל�Cɸ1>�>IdncLYSwqs�ޙ-���8�t�%�^J��Y�"�D�6�4�U��Z��|��|1��k�}�<�A�SZ���� ��z��s�j���6�$n7F�dV�N��Î��Z����'t���Z�iB�\yzK=������.�,�Gz�`Zs�@����'�:B�uh�!{���<ڬb�&�6�3T�����T&�1}��/"�C�b{�Ҝ���t����Y�x�k֓�Pp����r�1D�Y��=�*)z�{0�܉%[��F�qjZ�<Z�q��Y��}�3/MXd���yS�^F݋קZ��L�"(�Q+Z*j��NM�����4���+D˾`h�Ը��#���囸���S�����Yݳzj��1���ӊ��f=j�	�0R+s�.@�.wȥ���؅5吡��\�s��v� EW�҉�#w(����|�W�������P�h\Ӹf�26�ޜw"��tw�}G�%^�LgN=�^�j�-�Ȋ�jkԒ�i,�ǮY�����;(�P�3���>����ϳ��N�I�����M�9Mb(`%�2`�F1j��Pe��k�1
5l#j��2����y�/��Z���Q���d&��6kK#���j���L�Q+��[7\9+#5؀��Û�m� �*ǆ���m�1B�.%��c6`7�R�f��y¤V�P�-w`�V̸��XGA8�5�%�mU�A��#s55���4m���3&���o/5�g����ƭ��bm(����5���^�ئ���S[vbr��V�J8���s�3L+.���%�H�;���@��X8t��m���>6�-[��#���R�U $"���ۋ.k.`�eB�޼j]	���RjWm�i��sR��l;
6��؃�kYf�j�Z�I�.S���t)Q�T٬��7n,��m�mlX��X�2�l���JZF�J)t� �]M�V��`���J�*�n��!���ѨDt��@J7Gc��l�u&�F`Fh: ��0��%e�ȑ������#+���í�F�!�K������vȳ]�F�#��R��-p��X��W�p� �l6SPIa1��H����3j�-���AFef�����`�+l4)eы�j�8"����٢Rڬ*ˍ]pQ�EGnԴ���f�o	�`W-�%�IFx.ԣ4f�F�V�]ůl)"J�serǈ@����M.u����H�e�J��V��TmWm�1�Shm`a�gZd��I��k�5�a-��@�\�k��{k��S9끱���t��.�D��b�[�j,��c]3�n�&6X!��)�M�*2�ٚ� �@�ԁ�nȄ�Qͮ*`�	����	�4l�qAs3̸�j�$ZY[m�$i-h��4�����č͖�����bD��N�.a�g%�ѕ,M�������Њ��5�t���e0�[��j�)�ct�G��������.)���R���h:$�c��:
�r�U�m�XF]�M�,�E֑�����X@c[-%s�Q�� �p,%�i�ۀv���2fb^[h�i��.�η6��L�������p�Ma��a)�j̅�slKX��ٴ5�A��a�
��J�-HaER:�u�LU�(т$*6SM��%��
1 �G�u˒�.t�X�,�"B�HWb�t�˙DE;m�:Q��8H�q
�4m4������s�L�u�{Fgguv��Iv��Fx��Zy`�r�w7G�ۋ���������͈K)ܩ�v�gB�t�/mhgB&��KXҹ���O	�]K�35�t�-� �K˛��ih�m��ea�Tե�Sp([e�@.�v50d���]�q�X`�1i�.�5�ԗ�-YyCѵ��3n�&�Hq&�LA�$��� JiG����<��6�Ű���1b�Fb؎�t��eҭ2��
��0�m�cR��pWZ洚��P����Rh]F�α.fԳJ-�{&�4�P{^J�!�����V���sYH�ңAL	Ե%`.8�P-���Ј��e�]*ۢel�q���f�q6;�%�b�bb�,��5�Л�m�4��X�0����a4���hvƴ#��`�"�Ċ[yVX��F4�3t˻L�=O�H�(���J�K-F�&s�Í�l#2�7`���mv%WGc&�q�%�E��H�ŭ�ڻU��+U���ۊ`ril*�X� ��JP�Iuv��s3"tܙ^��/4K3a�R���5�c��,fĎu�0<�"K�M��#e�E1�2�@R���L�VQ(����4�pK*f�)\�c@��Z�!ե#��s)���&�neƴ�1���@��2��`�ۭl������GII�ʑ�7hkΩ�k��z�Js2�D��0�D���v$�Es�Sf](mp��4��F[GB���L�:"6\7%X�bX�*�[I��lenJĶ7m3�n�-��I��!u�v��Ł`Ѹ��[�W�n�a6gq�ƶ�$�څ�e�4��3�ĵ��q�p�MZ��j�j�Ml���-/S6��桌\�Ívp8/X��Z�� �8cZx�<����
�E���rj�qv"��KJ	�4�9Єp���ff�ĄGR�U�К:kD%�Q��n&�a���m�LrX�f�1�T"\n�\ ���2�Hn!�$p[Hb�S,�Y�Ge\�Z��f�g`�b0pdQ���[��V�����������.51Hݰ��d CdىV�5e�����]fȡ)Wa���`�*9�ֱ���pS�6b����H�$�l!5\�&�Q���s�)c1�ٔme��m��̸������!��vqr���u,*.�`mA�<3�1���K�K6��`(�-�ҙ�)��W�5����QU�,"@v�i1�/n�1�[��(عm��ɕ,�v)[�5pɂ����	u�A���y��	Hy4�st�^;6�a�ƀQ
1����YW�.)�λ:�Tփez��Qmi��bY�c�����M.�t6��CX��\M�R��ZZL�d;b��%�-��a���Vb�tA �r:�H=����x��A�K-��]m�F25��MJ�P���e#h�.��0m57mn��]Q\6�n͸�	nx	\�`�����6��Vb�YX�n�lg����
�uw\�X��ڜlS����X�F���X:�X�
;4����Q*�n�%�Kc���*�˛�¸�[HQ�f�[�3��ZL�&�#�����femK07#�.tд�kUFZ �S��
l����3��*9�ݐ��4�E���7M��-#n�i[6���Tʒ��uP�f�1����)�i�lD&-�n!����˦�K�-��5�h��B0����z�[��������剮���[����b,�+�ٙrb�$�4i�Vf��lkcZ,��64,B:���TL&�u!���f�I��kn���Bd�V�6�Lki�Ku�,��2b�!.��tr�6�,z�D.���&�l�#L��<7�M��p[�G.���tx��t��qe��$c)W�C��ɘL�mZ�X&ڱlƍm�5^���elZ��t�YF�T�L���"+I+�te�[�ZM��-ҭ��(�i�0G��`ks�����M����2�\\i�d̶ajd��B�X�͍��4��\k/c!��;3xҴ#��WT�,nd���]����H��D�Hv�r,�[��[-�X�Z�Q��b��c�C1�3,�ز�\�C-f��6+��1��ԫ��΄p�C4m���t.4�>>G�x���n��R�k����,��B��¹C"�ݸ%�،vq.&e� eт�(�f�J��L[-WR�WV� XəlX������ـ���U�U
��K)R,�*m�J��A�ֺ�j]w.�Fd#���-e(��w1�L̰`.�,�2�R�H�]��3#[�L��j��bk٪T�ݵ4h7Ec�Ce������47�\Ə���S,J����`̍��/;ΰ���3u�!Y����n�K��,4ѴVZ�cR3�(��Ո/K�.5c�M5����.����5�U"7!tf�fѷ-��qm	�D� SM�
�ݘJ1(
bh��2k�%Uvb��n�t��wP��L�L:k+t�ƶX�X-��[�j��
U��U��+ZѬ��ک��VZ&*��Vh��u(ڴ8���.pF۸��M`:�N]n���`��i��1����+����+���P�ɳJ]��g�!�p,ҫ�)lR�h�ea���R1�2ʺ2�l�6:�2�)��u&u��0SFwcvnsM=���#����f�%0i�b�5a-K�j�	�˵��v�� P�"�qb�Ӏ�e���-a��]ZqE&��Ue�!��u���d�,�hYf��%�B��
X��1��i*n��*ˡ��R�-�IY6ƺ��&�Pt� ˫��u1Z�A�ی�K�׈�&��K%c[!�t-�9{vX�uc�m�	����Zl�՗#Yy���W�L�^Ժ��P�C���%�0��,66�6�����L�)�Τ�1
�hZ�b���ch���Jg���Mr�gDh�F��Ջn���Z�5��p��mbpYo*$ڎ���SBٖ���� � �I�%4VRlL����!��u�](�;�ukmĩ��*b �K]P��]T��c.��Mh��\!�\h�
�K����n�������h�!�d&k��+�%�04I���!Q{]�@�s0أR�n�6��!)�#�KaI�B�Õ��6�1�����-�tRX���@�\��s+���%�J5��o� 5e�H�$5�9�t��G�qf^b�Z��J��3+	q���k��/mu��Ʀ�,`�Y`���v�&��p.�H[cKD�E�V���K�V�y�d�z��Y[kjv�T�ي��Z���K�le�n��9+�3���R9�J�`�)n�0HVV�k�ݡuCjC�؃1-
���1��mX�#�1�3�;6�۝�DLSP�X&-�6&�8;LU��p�CTt�֖�e��d�����!{`�B�f�2��R�h�n���k��Qh륔!�M��Dte�3.%�n�X�i��+�24�b��c���-�QɡF������8#{j�Bi��+��#/�����M�aJ�S����0���S1�G�m�a�m	R�Az*]�2�1���eZ6=�*�<�Z��hLZ7#՛A^%t�ٺ�3���P��3as5�H�+xJᰛ7^l͍1,��6�m�uSF\^5��ȥe�A���Hl���s#t�4(!��S=Jї��1M���pi�bZa3)Πi�m�pg��kxfF�in�G`�2l�WAv�4/$�٠0��
uѷ���@��"Z��.b$����:�3��m3	p���n�G�JX���L�Yi�[�8��W.meF�����q�vf&�m�+��,vƣƥ��5�������Ŕ4mՅv%K���lMS%��([.�s�-�E�p�X[U��7\̪խZ�b�\��sY>qN D�Bde��&�3#$�(BCI��A�a���0�(�e%����""�I@0�h!��b1��IBF	Ldc$�E&I�)&0"�04ƒŌ��ѐ�d�5�S,�0d#T��d��v���2�M3E��)	�4A� �HI�\�CM"$��)1�(62j1�J��B4�I���4%�5&F1Bj*.W����d� �آJT@X,���&�PA��\Ɖ�ȔE-�dƂ(���@cDBd�ch"�B<�$�v��X��\&�1�c73&X�V��7t��`9΅����B�er�+���"����%�*�m֒��d�4��4�A���؎P0����[���S;LF;Z��I�,�L�b�K�4��k\%:�f:��a-�����V/g=�Mk]PJ����vFˆ݉v.��#p�I��"i[�	nk�]n�[�F�R��2�-�+�Tv�\���5+�d��a�{h���Yq����`k�0*k�����Y�S1+H��b�����n��j��]M�X�`rV�l�S�ʆл�3D��RM�Sɱj��b&�Ki�T�]b\£]�,m�v��ʶ`sL�%�in��k3�+��#��m��봦��F�]��;i����
XU���b	r����5� 6h�l� �l2�m��t"��q���*��D�.���HF"V:�#,��NG)WD�ڔ�Nk�ʒ�)e.����ai�`��Q�Z��#u��+ ��b%ͩIpV�a�Q�Nf���lGf�m��k14³R�`\�u.�vKM3��Ǒ���<��d8uIYV0�gSXSZ:��ņ��1E%���K���t�KZ���6���5�շaA��jUv�q`clRj����u�m���B�h�p���f1m�K1���Hr�b<9n���uz�+ti�ڐfQ��֮%E��4ľu�3�γS59kth�-:�c1s�!8 òպ5�ݦ��˓Z�R��7.��ts��I�s0�KFкl5YC.�Y�Bk��S܊��2�1qf��]d4=r�腡��F��$�hl�F6)�	���B�v�t�4�]���Z����B6�V0�[[HX!�'b4k�D�Jbʎ� ���Q0׀�TC]Ya�XY�4m��HJ�س#�	��W)�0*:�va�M@lFڬ�]�X4��IGUN�s�ⅸ�]&�L]��sgI$3�Y�	dh�G�[(A%�#c�B����HZ4Ё-<34%,RlN��T���o-V5l,�ʑ��
��Z�z���J�e�)�eeAe����"Z��a�b
P��bR�U����C�=j�%�l-,k �o2�Zš�ʹ�lk,�3��GK%���?��~4l%dfhM�(�՚�[��5�"�f��.�56���d��"�_�!�C�Ả#2�eZҞF^M줂/�����۽�P�P��x�wdQ݉��A���aTtI{]�rC�$�
"�iU�:�V�U(SR;��A�Nf]k~�g/N�5�D�XqЋ�٢7`O���n���6�,�"sKP橻�Y��A���� �F�ר*�����p����x�@�3MoCΌ͝�m��x�i�v�s��ߨ8�s��@�U��%#��4;�4���Q� ��	+�]X��J�
|���h��C�����]�ߟ������KcI�<mu�/]A�l���P���Aҍ��FەͲ��֭5[4��ס�1�����/N��N��An8�E��"P�����ߐ�����Rff��̢�g&�̈́�H�5�$�)Q������Md�f��b��̈́��ywqv��{����.z��}�_(��� �RPj�������59g��� ��D�V�tr���ۖ�� �Jk��KLo^���eW.s+��s3F�ؒO����=�g�j���K���9������{E�r�f^�9�>z���;�wɯ�2�n�N��'��:�9��A� ���{W�}�ݿa�{ڴ^%&fkB�Qqʐ��n�ux���E^H����memm�m�x:S��"A`�����?��|���_L�,�a�uk#�f��s�Y�Մ�dy�U���]7����O����=�Ht�sp���]X�Vj���ǭt�Ε��ڀ�A�@+��nȟ��vh�и�Z$������!>+]
W�O"���AN;�DOhhs+Oz���W�����JL׵��E�6=wf�vA��)���ލ��[�0]���8������|��X9s.(V�$Ov�SΕ�N>�L�f�"N����Z�ٕݙ�U@��8q���8z�+on[l3�:S��I`��whW��O�����GF��\�!
�^=�> �t���yo,�/B��)k�@��S��Ms�֦߾��#;�-1�̽DL������^�b�/�TS��"sȺ�98�D@ ������# �O�g�����:��L`�ꆓ]��!a��ʎ+\A#5F@۲�c �g��~aǿ�hC�� ���n���M��������>kz�eW�>�sׂ;���}�4�U�t��i��k�8�S[J��z�8�
!��C]�7�Ƅ�	C5���	 �����l�D[�MH�C0�:��\�C34{�x��u�wu��ݞ�৑ur
p�6��28	�#[wp�{��H�=/����ޫH#vGlt��Ż��{n�A���k�^���o0G]�Y^j�m]��%�W�����4Z�a�Le�,�w�����Ln�{<�z�t^X,���?S����Q�����a@����0|F�n�xDq(G34i̯e���O���U�ia�Ր�����BB��r8�O�!G��V��N>9)��I�Υ�w ٲ��pAp:��3T���mkm7����aĢ�Ͷ�9R� vd��H#H7v�zko�@B>�aNAN8w�[3�١�,�#����Q�:D��(�|AMm�Y���w.hZ�!칷ϏS�[Z��A��n}]�$�+\k���eРVD�Ad�ۿZ`��<f~"p�_!���jj�m��/5�P�}^J � n�� ��M3�3a�ڬ��3S��"H��ȱ5�5{��)�)�x�h�e8rkj^iN�^�I� �ݡ@��H#`ݛ���QU���p���6����u����	{�^#��� n�
wN�N�9:�M>�����_6nrzV�6�L��̾�B[�"�V8�SS^�b"،����{��k׹�6���寊-b��%�V�!f��5K����(D��5�9��v"JY�Ț�Wn-��P��7GB�@�ivu&�5���q�JT���R5Zʑ�+-����[Ɨ���%�nH�:ʔe��^�Ju"��V��ShB��J-��˸L@5`k. ���eIA�L��nI����l����٣���ג�d�0�Pr���c����O�q��-��ЩA��ijM6ۆ!�3���e V;eܩGA����q��u
v$�t����k�1�z��>�>�x��ڞ� � �� ��F�%�Gއ����u��<��0�^�UX3Z�N>!NAN8�h�N�x��
��3�!�=�{T	�����^#v�j�TS$L\�rq�ڭxޠϸy>�� i�ݡGv=�Pw�F���뾡Gz$��Gb��]�ݱv��(Zr8� &�S�ў���j�~���:F9�z��X���非���Α©��'��N8�"ӡGv$i�6{ˈ���`��N�n�Cibh��:���+D�m�.���)@�lފ��5t_o��E��Q�˚̳�5�å�[U����%�Z����3J��2���'�c��49�b.%@d}<�%�C�zE.�B_���Ct()ʩ�7��y���ȹq�5�ߗ46�Q�
�� ~�Ա3��}+yD�Adv)��ۜ���F�J�G�	�(���s� r6v�J��%:�#���L�-1���f^_�*�~��W�67y�<'
f0'�� �N�ؐA �F��������<�7d��m)�Aݑ vOM�ttru;:��A�%\�"p���X��v�D�'P���s*�AĤ��4�W/h٠лo��A�"�����p�ѫ����P$��6;�2+@���<��^�Q���2�cb��ǒb����1�;X�J5��gTB��8��� {��$;��7�$ݡUX3u��|)���8����{}ߓ9��Q�U�bRff�.e�A6�z�`�ɢ
R'�zo{��S������y5�l�i�:�)j^�n�G�U�������_"�/]�W/�ޟ>��-��%�r�4{�֞.!���|�+*dI�C	��]͉�#�*������̣8鹽
�NU*y*��*�z�2��Kvv��t��n���}@��Qh�����G2�ܤ��:��\�����5�5"!	�����q�%	�랻r�Y���0}V�Ԥ����iŃ?m[꯱��g������l�o1�{���hGl��`�[w6�q��!�nZ����H	�.�� .��@6�2b���vvŰ���0��q��T���U���"s3F��V3��k��=�8u5�ܘѸ�P�v)Ք� s����X��32�������<r�]��"�.�5���*3��S385�G�:wcl�gELu� ��/9�B�h�r�f^�L�5�y��lI��Ĕw+�[��a� �y4g��LB�fh�9�bw�V��7��� �N]y8Hכ\�v���֚s�q�AJ�*\��di�M����ww�j��Y�]dUx�pjZ���z[x�M
��*�b0WP�j��[��l��c�W�.}ǻg�;�ZcH�f^�32�Lu����1j��I��}B���J�����13�\{�� x�P;� A�Cex]��ؾW^�]�LZ����Ɇ8
�5z�nڍ%C�B0�V�K�i5�]i��gM稸�C3/hF�f����p��o1�x�5�a���L���ff�e|"�P1�|�﷪.6:� _D�A �#�k�.��g���b0n>�|R�%G�ݑ����AF��]��m#���e��̠����a��{q����M�13�{^F:JD;�ths*�q(L��h�K�Ȟ��&����8P�z���|�c�_FwoN��G�|�&�{��P���՜)�#�7�Q݉ ��AwhQ݇Q]R+ő�VN���g���b0n>�%|A
 �ٰA��I�����#�i�?%������0,_f��F4��G�ꉳ�f�X1Qe�tƶiM�V���A����������~ͯ�M>4H�6�ªє�ZQD,ݴ�i���k��=y �q�Q,.5nu�6²��BY�M6Ԇ��aH��q�c��URm��L!VZ������.����[�pSLQ�g$R7;��6�Ў�n�,��+0:�h��J��
,,��$8�R����xdR+����1e�ȷ�Aś�/Sܩb�������l�F��飮�SiM)D&����T%��{Zyn�6!u�TF~?������O���whPY�	+�s*bg��f����ݦ^&#���Q�U�J���@�� �5y{W��hG9ي�g���1���>��f�����i.��4� 3���3�"n�
v$:G9Ȋ/�����ל�y=pvWh:�#��l	!7vl��Mx�9yv���k��x�� �0���СT��b#q�13�\$p"m��e:��R���� ��7v�^݁$������c�u`�YYrY:dKɊI��ļQz����>�� i���."gi{ߢ��Js�WF� 7J8� ��,�t��6�`GL�a�T�6G,u6v�����OD�!��
;��H�ͧ)w(���v��q�WtwfDL��"���Ϩ���"9�z=Z��wfv��1��x�Ǎ����ŧ��hΑ�����q����Wva��S��mV��3�͹�*1��|GaӜ!Ru�5Y0��ֈ��`_l���Ú��|�NI�}D�}�\�lC�Mr��l�G��ϫ�vG#�����_o���Qz�Ϻq�E��zD�Yq1��fh�9�,�ߜ���.���{�|0
0��܌)�s���X�ې8����e��9���^�C9e�4����̢���p�u�qr,MbÍ؉�|ʑ9'\w�&��A��۱�H�	�X-!Ϋ$l�4��Yb��]q�3HKuI��.�U��f��XM[eժ��_�(��jS���L�;"'E��^��n��*�b�Ms�_"3�e�3353+�bP�w2�k�s7�{�|Qb��܌B�G�,X���l!@� �"z�G{�{��u��{z�9��fP��]2�Q�Y�el(*#pv����Ig�Ӟ:s���jz�����]Fh潊�����-�<]2'w�S��nќ���9�#b@��m��jn��>~����`����oY�,���]�4y��?\}�|=� @����ȧ��Uw� k<{����z^��Y�=��N.�l9j�mCs����_xPPź�=�t��O9�Ѽ3}�n�u���E��:+7�ݞR����N�4Kx�v�[��2&ë��{� ߞ_a��'�s�ٚGLZa��o��ġ�wq�A�5M�*6�!� ��p�U+�Z���ܼ���V�1������V�/{�u�d���z`��B�SDE᳦!k�a�3��eNA���-�>�B��������%�̈́]�<�E����/���B�:X�`/��0���u	p��-�,<�4(�.����`���� e�C�ӑ����a��M!��0T�}^k���F�T��1�G���b����ͻEr@Y����U���k-�@��fIys�.t_[�%O\�B4��`z������V.��E��	��3���[[������*��{y{ne�{��	���z;^���9M�QIH�ȇ��*����-?d�}���ȱb�*!�^Ѥ�sC��<�v�M�VsY�^)R�r�H�vq����4<;�WmΫQ�gKlX�����zS��v�_�k24g�{;Y�k<r'�sx�� �-X��I����SV3Hi���.ӟ[��M�/~�9�O�bȈ,/����i����эAd�Ad(�4!0Ƌ�T�D�4b�EE,h���Ww`M�q�i�B�EIl�4j#PX��2��`ؐ�#s�h�d�M6("-��ĉ��b(�!��F�`Kb4f���"��"�����F,i(�j1`̴cDh��E��(����m���E��E$2ɹ�%��-j5�ѴjJ
�eE`���E�E�ZaIA{�w}�����w�ye}� s�Z~) ��JwUB�JH,>��H)���`�Z-�j*�.Z5�����!�y�����������y
!I��� ��Þ��L��I� ��
#��ي�k���*�T�Òڠ�
J��nd�) �k�����n���O$ᤂ�T� ��w�nH)���9h�M��v��hמ��ƾV�n0�r�I[釿y��~/�� �S)�T�|�^�����ֱ�/��������v�RU�QiTB�]����Ü��L�d����Qi�o���۟w��?t�Wz�ƭ]5ut���&�R� �A�wM�H�J
 �X�6:\�o��T��RTB�s��i�l���S��I���ʨURW�J|,�n��ۡ5��FO����
Ag��ֹ���W��uUCRAaS[��c
@����K���7=��Z-��|���(����
AH/ky�Ûv��]���`)4�L7�\4�R
Cz�O����g��z�cV���<	�P~RAI@�0��p�&�I�ܳI���������Z�ϵ����~�i �
@��ZAH,�d��T�) ���桴��c
@�(�����L��P
��d}��`��{E��W1T7�:>G�>�X~����QiR�RAh�� ��Ss�3`�I
�s�i ��
H/*�)#�֫߳�ۻ����?0��p�&2�
fY����i ���YTAH,9�\4�]����v*~��t�d�� �@�> #]�@P�%$��ݵ������(��)f�_�o���m�n��~_�$���@k�|�}�|�<Fp��x�eZ�F?R�C"�p��CA���V_�i ���R
Aq�H���Ü��I!�T9E�B�G*���s��i��;-�+����^Ǽ����'s6qs\�����>˄,Bc��fe�{�Wq�����-i�ۚ<�V� Ar��uK��ڥeTݣ3���Q�l��E� f贂�Y��O��R�9�m ��
@�(���RAd���H�p�=�?n���<y ��ް�� �=��yZ�u�pߨ����RAh�@��� Sw��L�%&��{�_F���y��h%Ss�$�����kןzo��7� �L]RJ�{���6�t����Ö�&~�@�I
H,�Jv��-%$��H)���=����ᣁĂ�]�) ��,1�AHQT�E�Q
H-��Rs�3ᒒ
!�Q�����m�Lu�kǫ��ocD��8�/�8�Q��$x ���p�&���P+�,�A`hi �`YtAH,9�\4�]� s�Zh@����?W������\��i�Hz$��ý�p�Aa�?v�I�
H,��x��?_8w����޷��x~<�Xw�\4�R
2�H?������~k;�6 S���L�%$(C9F�
AH/�H)(B�s��i�`�H(9�4�XH/�u_���k�W�T{��H�'�j��'�IT��~s����Z}E���)���) �=��6�R
9E������� �5m���3�g�����Ȍʁ���d+�؞�&�"�P7�Y)q�u���/0��m�ǆ�	Ɍ��!������=[���{w��tlc	QYPR���q�����m��L����h=��F�As��
ʘ�j�\SK���r]��1�`��lkCL��t��,�x`Y[aK3*���t׎+�/�-�6�ښ�)��.�8�b�����B�)-��GXa�����m�6�)v�`Tln�5]��+���v �6�KBj�6u)p�,[!S*�i�K�39Ͽ��������I.x�Xh.��c@X�vz��m�!�v�����ֆ���H,>�.H)������!I���R
Aa�r�}) �s�ZAa���s��w�g>�y��$�A��$��=���ɯ�<��놙82�
�f�M$�P,*�)��.H.�\��z�|e\�nmǽ���[�޷��^������o]�>H,20��E���Y)����g��:럽��k{?qۇ���~���v�R
{E�B�UہI ��9p�7���߿o�.9�<�P�3�H,4
���RZÝ��L�e$
r�$�IyP.肐0#�%>G�*�ވ{��X������ֽ�;�-?�*2R�RAH,.{;�m ��9�-&����L��P��Ü�ݤ��f�=޽�u�3tZA�(�$�]�R
X�L;��i����P@ %��'¼�+�a?���K)�ϼ9 ���
J���2le�H�Zz,՚��_o�.��3o��DAH)�T ��\4�_̮U�x�r�h��Q^-�K
�9�m �r�I�es��k�զ#��z���	 N�d������,����ÿz�󴂐��;�- �RAk�p���L9�\4��JH(R�H,=��~���}��MRo��b��!-�(V-%!@��sR-�`]�P¬1y�m�U��D��~:Rt	Ԓ�?�ˆ�6�H(�٤���H/*�\� �
�9ˆ����s]����������~�h���$Q����׷\�o��(v$����Ci�����ZM�Y(e<����Ü��I!�P��u(��O|3��Wkg�_E�T}hVI�������$�}ý��y)P��G�H'w��y͝���o��Q�?|���	iҬ��eW���L���S��L9��$�@���O�	�z#W��oR�ks����R~���2le$
?r�$�I�T���7�|o)⡼�ᴂ�`Rܢ�E���v��V�^���Z((��R
AyU@�~��w](�R�������G�>:@�"
A@�h���!I���R
X�L9�\4͌��P�r�$aI�P[
H)>��>���߷����ˆ�:�H({,�A`hi ���]Q �C���i���v���{��Mw�w^�@���O��YL�n#���#���~�s�Vg��n�C���
@��-&�) �S)�TȔ�Xs��۴���T9E����9wH)hÜ��L���{]�u��ZACר�A`�X���9��/R�Ks�#���	'�)�}놙6�H(~�H,$�P.���h�s��m ��~���>��z�����YG�i^�k�1p�6x�Vԩ��3l\���6�`���̴��}$�|��@
H,��O*�) �����m$k�U�x�¹h�{ݨ�����w����?g�}F�ǒ�높
C��}�߹����9��p��Z?]�R
X�L=�\4ͲRA@�(��h�{�_-r�nW5���� �j���t{�k��Ϯ�m �1����ʢ
A�P���i��v��w��i�M��$�@�>� A�#%;���i) ���u�aH�������vs����AH/�P��X^��봂�P;�- ��Z�����/��������>�?h�2�w��0ED஋Ju*s"�.c���uN�:d�,jQj���S�;�9��.b�7�٣۰ K޺˺���۪�^�$����x{�z_���o���LDc��sG��a��5ؐF��r�dv�q� ;Y^N3��G��Ӫ��d�+}^j�Bn+hמ:������e�4��^�9�$h�t	�;B��������Q�����]�xDM�NeX���h��G=��+ӳ�j$#���A,J�lLF�Mf�+��h��j1��6�n��lY�-�k�0={�'̈;�4Aݑ�vutm8�J�c�������o���s3�X�Ԩ���@�T�@� S��nMȰqD�|B<�\%�*Ia<���%wf;a���f��w(��J�/B32�*&fP�)�~��7tL^S�r�˓��ʹn���Qs53+�1���h��h���J �Ǡ���nȐ�mkji�E�V�]���{5��J�[�œd�n��6{g� !��Y�S,��c����������?o��>�Ę/5~&�h�}ٝ�m]]J�;M�mIQqs�� �?���4j9�`�8�33F�v;���L�"0Ev$5����H�u��Q�wf�>ݑȅ�r�aQqR�#���/9jl֦��й���l�ƚ
�L#sw�V�hMWM�����#��i���-^*W<�:N&�*��/5��5ZC�9�N�|"�TL�ֆ9�Z{>�۹�/g#+�M�� �;�HG+[SLO]�O][�x�٢3�O��4[��TB��}V�z�ff�9�pDq+���um��<X�F�}y��j�-ǥzw}��(��ʕ̹��,Li����L�ڟ/s� �0|wv�J�Ss���n�S� �DAP�\�Y���A�*[�33f�9�Z9R����p�T6���u�}Y#$�g����Fy�}zD��ZcC��2������7Q�� T�̬��sxs`�`Ǩl�Y��n�(=ƟE�(Kʊ�u�ǅ�Jʕp�qe]�Z:���B���t�䚈�g�;�w������/*Y�mu*isEwbXBgۑ3��4�gK�Z`2�M�dR��+tX���S�T종�mq��)���ek�R�!+�:�a�W+WD�TN�L����K�T�U�p��F�[��8���p�]�6r�(f�k����J�i�GX�hбűma-��ט f�)
���[�2�ֱ���	*��e&E���	]�˾��~��?Mh�NԺf�����8��Xijl�\��A�Y����B�|'�!�z��;�$"R�O��:�,;|(aWh�O��m��G7\� ��h�wf�wtdY-���shT%k���Y�q7YW)�4D�Gv$�u����3^k���!���n�㘲������da�p�9�t;|��귉�s�3���}z>�����Ѩ�U�p���܊��绻p�]�(�O��!�)���Px�������AX���y2��V���O�@�4� ;�4A�$�7i�Qf�cW��*�X���u�'u�r�q��F�@�Ă��M�����K��17@��4&bMzMThk�cr`�͏(��R�4t��ZiG:륌d���|���
�O�G����]\k֝�U]��9��C�@��ԉ��9�AΑ �`���
v$�H�#�D�2/�yt����®����I�V����o�6�QHԭV�-�.0�k*��Sl�ܳ�UV�ieü�S8�5�Lf�O���s��;�"��J��LU��%����I���3]W:��j�;e���_�뙔|��c��5ܭ�َ�L��f��g	��dܷA���w7�i_�#-���A䔎Q<|A���
�G�m��;�'�#y������g�]���MEwr����G"�P�wbH'H�F�Я��Ԧ�lN.Q^���CA�"B�\�8]���,7�@��IG�ݟV�s�r�y�=����N��6�7e�y�h��h�/��V�mf@ʡe�ц\A���M?�{��}�f�����whW�V����Σ��˩n;�t���\rӂ;�����#�ff�.e'�W9/����8�Hs�������i޹��x�SD�F�r��C�����v��Oe|"<B�3F��R�GO|���9�Ms$�p�'�.��wٹ�ɭ��m��^��<�a�^�V�x�U�0���yu�l�z�zou�G>��]O���z���#|.�b�!���C�N2�3/H��,LhJ�W���Q���JQ�H#H��)�o6�^NsY)�\�q�l�n.�V���u�G��j�:�&fkB�Qh̩C���k:e	t�I}5AmH�T�+�y]Y{��SH3���� �vȒ4Ǐ���K��SY�A�OKp<�A�e���t�d٣,�f�0�*� ٜDc��4�f�}����XC�{��v$��pQɳt��Жޡ��"�eq~�V� n [���F� ���2�v[����\%�sãA`��:����ɾ{���L����!=�@��(�Q�FL��݊�p$}Ne�<��-Yp�e��
�մ��g�][[��SH3�j}^� � @����a{7�pAC�$Yz��c �(䘺�
��K	�
�A��V���3}��;SX���We%F��� `���Q���BU:Hd�dґ�=��p�r��ut�ʃ�n��ε�{|���N���L��w���Q�@�ٲ���_�#]���<�|�ƻ��x��T�q� �"<C�>ݏ`:|�\7�vS�y1�1Td� ��1 ��$�޹�#5.�Z���R�J���[�&�Kl7�z���\��`���{���};m�SH3�gVR�U��4�يD��㻴(ؒ	� ���};�/��x��
wy��/�aȆ>�Kp$
�@;�s�yyw�0���ӭ�y�4fYc���%������H?xe�m�o��������{^]���͎e\F8���@P�=	�Ʊ,DR9�
�G�j���%�����ݧ�қA�ud׈9���{ʿzڼ���<�Ϲ뙕�F8�A�B�;��r�W�e����Ol���}��Z<�Nf^���Pm��	}��G����v���cB~����{���f���G���4��{�_U;I��p���>�����t;��f��4��a��>��1i\�ڀx���v��2&��e+,��Ԁ��g�,����[4�dNL!h�TD���M���:Ѻ�HE���U:�&���h��L�8�Q��A��'d��k>�|���ػ��5B��u$�x{�K�d�Z�'v7��b<�5S���r/	�1[�4S����oe� j��ʘq����	�-������|\�Qc`���M�&n��V���$�	��"��qv��;�e��Jb�{�c���"	f�1�m�:���~�lS�Ѿ5r�ٚARV[Rۘ�/CV��3.�7��Q�0u��1��T�ꝶ�ٻ۽���q�M��ݻ<3qﯛHp�E�ߏD��0@���y��<e{��&�Փ�jqI����AֻU��-;�,ڱ�̧����{���aw��5��}�'�C��\����y���o�֧{!}�[+��������ɟ��u��Zfmǽ����Ŧ��ϟ"�g���x�{�0G{��شF=ʪ���`[�����7Z�7wԫ�g��Ֆ���V/���%@�����u�ٸz+��Dx'�ȟ%=��+�V@�)I��C/G([��+�����kݞ��8{7L�B��C�U��0{@y�����Dd��GV���*g�z.C�쵳1M�j�7��$��Jv��Q�=ѳ- �9��Ǝ碴�ч{+{��[����Ȉ

����-H�5cX�V(��آޫ�IF�&�Qb#ʮQF�ɩ�Ehшƴmwv�E\���U��cQ�[DF�"�b�r�sBm\�r�AQlj�\�
-��v��Z���lQ�F��1�m�h���b�%s]5h��R *�Yad_��Wt����8 �޷X�)i*�h8�%6�u%�:�jh#,s����
j0�ج0q�+�6Wk.����䙮�vH%���YX8h���J)�:���\[M�]�;C�^5|���<.୛B��R�8´n�l�6��@Ÿ�HQ6�Sbnm�����u�,!�){()��Da�,.����1�v�c��16�́C4hRk�`�a�	f���K).�f��)jEզ�(��0��0�j�]B\B�����P����.!]���m��s�v�j���&Mv,��%��V��v��6�Ffµ��l-u��Z�Z��B���Ñ���Zk[,�GQ�h��7�Ű����㩄Ke&�mU9ژMJʒ��h]�Wk1u�J��)�����n�s��AB[]��T).���Iu��t�DF�GV�1;6�[��2��P�(���iu�!M��YE�%6��.�\��j�٣m�LB7���Uf��t�G��F����[&f�)Ic���%ʆ	@Q��5��c[f��m�j7am�T G1�41���Rh6�������V��\�3��n44�2�{Bf*���Cnf�,�ʭ��-U�ѷs�����d�ҳE؄��7��b(kˬ��ZL6�n�z#5�΍B̑:�1��Y�f񝉚�FP4 ������<5��y�\�t4����=u�S��hГlMB�KA+��UqFh-�1FM,����+J����k�ܐ�
Ȍ&�UrKBfU�U.,��	�&`h��r���f\ǲ��K���X:k�C�[](�l��6X��6��Ki+��^De�ד�IcXLT�T:�h^���e�ک� ��)Kv�����p5��e�afB�i�+�Za`�鹥�;9eBeu��j:^]�"�LV�a�Mr��Q�Ժ�whFa�jd��ŇYcs�V�X�c0���U�f��m�\Vfq�2���m��.��m`��Y�)]�B�I.�fian���dbЦ]��cs�'wI%���het��<�"�y��c�v�\�����*��3R��٥]-�5bx�+)��t�(1b�Yn�0K1lAiX��6�.�Yo̬m�֢d�6�q�Q"il��js�6��` �W ;��^SE���ua
� ���)Z�(܆�]�&zd���W5�&r���r�K�b��k��T�l��J8!��������b�����.�	�5(��GE��ź�Glki��-.53���D������h�p$�0|}��)�f�{]��[t�*e��Dy�C�Ut�d��qǧ�H�t��	"6��j���lyx�S�]�.5��l�x�Z� ��٢���[�d���@�ī��H�� "(��ݡ^9�$t���l�'�p\��zݜ���ۧ���hc��qʔf\�bŃ(��k*��]��ޒ�2rŃ( ����+�1$q�����\θ��".G^��)�]Tc��l#�"�"�݁>#O�ݞ��,��g�p^ND�K����6�8T�< �ٯF9c�|-��_v�'�ɛ�d^h�_G Y+CMG[(؎.f�W��XTٕeb�iZB�	{f�&eB>��B��xi���-��(v>��!�O�O�҇�0_c��	4}����O�Fh���/�O��=z��y�2>��Ԕ)���sO��k�,[�v�үXS�q+� �\���AѲ���n�׍7��obS���;�=��R�p3����� u�}��T+��j�./�n]e��w����
v"�Ԃ��5��%�'��4���%������,/�<���+��B}��Wߡ�{�v��N��9̽"}�,fUL̳Q̩��/s6�ȃ� ��P�R� �����1#��\�->�AN��!������O���^�=�,Li��^�2�`�9�m���Uv��qW=m˫��q��*#7��әV"�u篟�w����?Ob۳�Z��l�$�G�t1��H[WX�G]��Y�;1���{����~Y�>a�߽^ ���M����d[X[��巫3�=�f�	��by�9��C�V��}�oRS��-�c�b�8�	dC���p���H.C�P>8�A���¢ݷ�9� �@[�$�0���FfYq1��fh�+ޮV��Sz��м����[c���E��N���x6�� �g��aw��e{r����4�Bg|%�eA(��Ԭ�����_�e�Kuq�Ẹ��M j�����#wj�8cjj7��u 3��\�A��T�V����6���x�%4C\��'�s�BH�ǖP�� �0`�o�U�{.�S����w:G�S�{;�@r����:�I`ݟ^l��.6��.��Q�=v �>7�S*���Ԅ`Ɠ%�Z*�a2�j�&�^V�.�R0`iVcB���z��Yq1������_}��v~����Q���49V�f�G��l��b"cBff�#�A��|�i�����ϓ��<�'�n�i�ek��|�M@{"Hӗ!�*wns^�7Z5�V"8���s2�\M뎯ܿ�C��KPڭ�w�a�=��6 ����i�}j55��Nh�;$I@�ݡO*�V#=g���⥨�	� ����#H����v+fyH���:�ag�t��t�٭x��y��������,�M��g���v��F�ܭͥ
�{��T���I�ff��E�fT��e�����_��ߚ���{O����7�F�A�>Y�D3�e�Ƙ������>�}�;���i�$��%���9��7h�ƷQ4L�tf�͠����]U{\��8�{��̯�c�G�s�OH=������6�CC�[ͻ�9=R�g�B&e���.f^��>��[ތ�!�8,���E,��C����qqR�p �"!�Gv"�ۗ���6�	�ލ�(�r�3/q�)���]*��b�BX��q�Pg� ���e�c�f�e}�}|�U�y5�?���+ǔI�@�XU0�G�D2�7#�(�MT>8�y�4G��Ds2�̲ٗ���Y��7�׶��{�
	�ZVo:��⥨�@�mP�wbA�Z
:j���͗����l�~� ��|��� �����n�ϴ��6�yԶ^.�'�I�ޖ�A5w��	Fo��;�,�N�
����g�wIY��{x2l*�v�5ZF�PQa0ͻ$��.��A,��n�c�R��i.&��Ǝդ3c��n5�s(��Wu��j<7b��c��C)	n�d�պ�Z(��nih%��+4k�K��	Cc4�]`�-��^Lh��l�a*A#��gHv:��۶b,���fSR���l&#���t̽J�	H�u&8Mk��ְ�)��ͦm@3��߷�o"����Rk2(Lp��΅.� ��f��)���k��Lٯ����ٸ����͐wdO��Uϲ؞[���}��&��ýXC� �j|��B�݉ ��4� �(=��s$��܌tH ��yAQ��A�����H���vx]eu�Cσ� �iϫ۳�ջ�&�O�Bۊ9Svw�g6�LT�A"����IL���@�Q�킯i�Zׅ
�M�qO�nȞ�˭�[�6�[ey��7�4�򱣰��H���2��ѡ̫��f��^�EVx��} &{Pb�a�A��P/yE���fe��c�׭u�{��*�ޗ��߻��7f�/K��@m2hAȮ[AC�i�Y�E��\08��=w�,!����Bz����㻴)ej�+����RjZ�"X��ho]�3y��Ӝ�c�33SC�,;��r:#��ʚ7����fT���u͓n,a� LKP��N�S���*����m-�8I�,򝩫�H@Y���{�^0^��&
���0���� �G��ٯ�	�K��ٌO���+τ��:�_�)H���n����(�?,���"�wc��bR��Z�_:MZ����t�{�h^�f%G3.k2�f$��#���$-vX�`��?n�鷆���f�r�8�E##;��I��}�V"�*	��9�\D6= ���bSsq�W��Gb�7<���<o�3xo�xu�����e�	�33`�Q��)-�C
��� O�N�V�����3*�Q��XY��f�.X�Ɩf�.��|o�}%A}�ʱ���6sN�����C	��)fU��V^��蝽�D�5>��F�G���x�U�Q��p�-��Z����˅&��q"-m
;�W���"6:�RU�,�Mѡ}�2����L�7�T�}���Y=ں��	�Y��K���*#��dlcfU���R�6�H&��IF.j��gD���|`�`��=�3b�d���x	��]��yܹl��y>��d P����`"s���tfm�� �<�Qމt��b�!V�R��rM���@�'	3�:� ��� �H�F�>����Ոev=�p�~G����s�ՁF�f�£r�8���Яؒ	�O����)��\���M��P�@lp�Cl��JW6m��6�{F�=O^|���훈���wf�nȟ9��}����ɖ����ip��k��|��#Lx��wk�L�`�F&_2kCʹܿz>{�(B}�܎�c[�@���Ǡݗ�l3E��zD�0���쁦�|@��]]Ċ��k:�:y�]�cW#r�ѹ{A �Am{v0:D��A��9�ܢ 0A��x��#vD�������ow&[(3�{�@�T$�7n3o����M�kU.�U��)�:�]�9}��3�SS��\oT�:����X3ݵs�������������s�|�tw+����I }V~M�3;�fഡ�p`�n�JZ��D_���@	f�����3x3a�
��;�wvh�7dJ�|2�d��2Ȉ�.�v�[q��G2�°3֚�r��8_�|�-
�`��)�	zl��>��>�Џye��32E��⥁F��p�]\K��)�<���}_u4��١�U�1)33A��.'-�\ܬR�w��S�zD���}���E��-��A7�4{|�Yu�l��F:^@� �whW���n�]B�22���{Lãz���a�P ��q�Oٗ��,Li>Ӯ{�_}���W�3�;�O���whr�j��wjɨ�f^�6D��"�mFb����x��b1�33f�s(���̽�_o�r�{:���!OjV��(Sid:p�<p`������(#�j¯����'X�������-Tj�Fe��@l+�&Bfe	_��e
{�uL�5x�U��)��]w��w1�_|��b��6}z��!>>u}��.���]5J�Ɔ��U���uW[ue�k;g\ �Zem��j��4,qaWfi�֫z,&���úĶ�ssI�G��F��6�.��A&�JL�&���&��ΫB%��Q�BZY���	@V�D�ca+��Q�3�4�-����!䩪S�&�R�k ۜB�	�ַ<q#s�̖�4&�pv�H��L���G�6:Ҵ"9Y��}�	M��[��ѡ��tn�.��уSE��%5�7���O��P#=�hәV��fg��/U���P9�ao�C{"��٪� �:= �s��̲�cH�f^��.���w�Q�+ܩb�EFwj��=��@��wcfӹ�⌊#�y�Od��}H��͐F��a��"�0\%��]��Z�]8A� �ݚ�vȐ� �v��0g�.#ė���a�����i7v�J����h�"ƍnG�$��u*��������/Q��LhE��ЄnȐF���ݕј�M���t*��*�VK�EC�G��Ȃ���:q�%��=��x#g=�Oڵn��K
�ek��2Q�����E.���m�@)1^f����$�����Dn��ڶ�Uj�T�C>�)�QՂ/w��1@���ݑ@�Ă	� u4�<ڒ���Xj͡��/���z�F��Q��7=������n�
��͜���K�^���S�f����h�a�����MZ�$J#wz����̋5��Dʔ�e��o��0�Չ�2�O4#�FV!����`�ܽ=��ׯf�'�Y ӣ-GA� [���a�A�@P�;n�uB�j�@|����������Y+N�N�x�V��!dL��p��;v4� @����` �"���G^�Q#������ê��A�ȱ�[�P>/`	�sw2B������z��o���v�U#�q���)�5��T�ֻ�l8���2�t%�=����Ը�hC���wd-�[W�ns�F�u�:�D-H�,��D�@��E1�32�e�������}瘛�ۚ �/��9ܶ���N���f�gH������o.6�7Rn$�1��s2�C�_5^9�O��V��j]���x^��w��7# �G7lq��<�[���p%��jx�l�C[,�r��[d��uR��"�CKbVFؕ�6�6�uS�yPpEc����Ad(��z&�~�XX{�܄��~~���{�f���cיgv\>v��)�!�/c0ະ/yzmR�`�����x���w_�����P�z�Ϫ�&�T��F�Qzl�4n�0���T�:l�4�q^�[�I�'EOIQ�����UQS���u�L���EYo/����"�(y��:*q�Qp7[m�@��f�O:�/�xP!�m�[�}�L�i�Z�{�Ϟ0�g��0zf�Sv�D�U��3Rن�M70h�F62N`@�1Ȳd�Um<�e���Y�/z�kE~���?w�NaX�^Ǭ�y����k甗���}�.�|��5U�_�B�[��P�D���t��!�l�&e�9���'�~(y�W��t��8�\�M-,��4^'�\쩺�|b�[PV�z�'�;Anʾ�X�<`j���������|�I�%��C�{d���m8U���|ߜ~T�(w�L����tzy��dv'+(D�a��8�1{s�j-���yWnH6v�ґ.�(�q��k��+'6s����*��V�""��0F�oE0���c�����[�>ع��iL���V�'\��C:���y�9���w{	�M޽�w�z�ͤ�o��s;60��[��/g���=�w��^�x��So�"�\=���>⯱��c�ܔ���
dk���
��!�i�?.=OK���h5�nQU�G+wqT\�ͪf�DFѨ�b��cV,Q�!�jɫF�Qj)�F�h6��E5���4j5E�,X֣mb��F5cE��m��[F��lj-�TZ�h�(�ɍDo��h�5�[�5�njJJ*���h�-�Z-�rr�Eb�1��ڭWc�����L�d`����	 �t����&�8�=�ˏ��R�� �ȓ� G�����*�U�p��q57����I�3y����7��`�j	��j9�\J3/~;�ٜ���tw^Z͇���U�T��28[>��"A�QQ33Fo^�׼3>m�i�)��-,��"\gʋ����Z1�\g�G��Vb�_@�Gvl�v<4���Ȫ�{�0#��l���S�s9txDq(s�ޑ3.����"���GlT���`�ǣ׮Gl�Uct��[��jgp Y�AOhQ݌l�k��R����W:�	 �ڴe����䧽��i�[����Om��T��z>��3Y��Q̩�h�o��x�=�e��noéC�(3�yST�oM@]�|(�A:)��,)����*db�lq(TΊ���B�8�M���ⷘ�t��Q<$L`�TsO�f5 �F:s��Z=��;ۚ׋��?k>��v��!!�O��ݽDy�,fU����$hpNa�n����-V%V5�Mo��jg{�`B{^݌�#k19!U_.N��h�M
��6��[K(�0�@Y���sڵ3�Q�6���ue�)V�
���P$ADA�ٯ�dOgc����Xԥ5�}"�qvt�s�:A�"`̢������11����Ώof�xq�$3���w[�7w�h��q΁ @:D��t�F�x���Dw�FH�n�c߻zF�[1�33E�[(ν��ua�|�k�uQ� �>���x�ĐH� �ݡBqn����8�k��"B׏\7��Mc��V��
Y5�}�o3�z��W5��=R����e}���p��6�`tuOu(�t���.��
�N� ����:�NY}rY�z��~���>g���$曻�;QS�svq�V�r;�"}��b��Y��A��y~uI�5#��p`�>y�N�/�����gٙ���[�l���JZ�vЄl݋5͠Z��v��6K��-, 4��!{Ћ�
�Y��	�6�a.ã�����-�l�^!����cB�F[H:3B�G!�R��](�A�G�P`hͳ�j�(С����71�´Dh녗.�n ؃�m&���BUm�;��L͈��+`�p
�	����=b�Si��w���!��X\T�%.��s(n�C�g��fj@�kH��EQtܹ��B�z���.3*�feڤ��h��7舖8�Ts7�Eş��D;��}��hL�ѡs(;}4��X���S�~ �"|�����[XZ͉�>�Y4AΑ'�/"��]
�J$HF����` �4���g)�T�����q�g������,F8�9�z#v|6��,Z]<ډQ���� �b<wv�v�ն5
�Q�LJq�1�$�ί�o�՟GyV��i33F�9�Z1�A�٧R����;J¸1�v��o��ïvg|�)d� ��"O��7v��N�U�[�le!H"l�4A"h� �r�c&�GMa�i�X���ڷ$!.Xֽ���/��� 4�W��IL{��uWKzN��Aѩ�
1=f�.��N�Y��Ӛ̲ىC����7�w���//u�����N�)Ӎ�V�=$�32v��x/afcp'��Y'���˭�ͺ��4�}��%��+���+ic�:�c����� .�����'B��:�ơ[�w�bP8�$a�7�(���	*&�N��f�^4/ޢ�G�̽#3,�ݲl��XR޶��ǳ��	K'��|3��ls*�}��٢��e�x��C�C ��ʧ�S�C%�&^�,m��u!��E��]�x��I��	�٠A�������ǅZĽj�u�k,}���s�W�����(G��2��F+�'�������wVhŹ���(�M�i��؉�l��6����E�Љ�uЄ͇��1��B�@;�4vD�v��O��܌{Q��%���u�Oo�*��H���w7�i�`�ͧ{!�]s��}�S����[���
��9�$�ݜtb�����9R$�J�4A�'��0|@��z0��b�t�\#q|�Rȴ��c������:�W�{.�z[=��.�[�l���a���k*50nm=������{ànmL����-^ݯ���R=�h�9�b.� ��&��خ����P�z�sDn����jq�y��j43� �R�����}�o7��Baf��"��I��A����g���� *��h���0�� ���s�I} ����0��/��׿�w͋?]����8���R-̺�U#������`�ٛbX�`	�6{���zh��4����Ej�:6���1��[���cV1\��"�(P=�lĤ��4�Qh�U��_Y]��s���>Jv�������ڍ��)d��z���o��Y�]횎r��{whQݏI��#���wn%��G5W�X�e���S��P>8�Ilz�� Aݐ4�!	b�U�8rqϖ@di�}����W's�j���qǸ�� �lUlNt��jɝ����k��q*�v�v�vpV�+�*(��a�Z����jY����dF?/t�7�߂B�|??�WĠL�֦e�^�wvcLX�u_`��,�cT��f;�ǵ�%�^ ��"|F�#wk�S�����翓�����J߰�4!f��˰��*�V�g�h;6h�˦��+��bݶ�HC���-m
�ݏI� ,��z�-oz�� ����d,�Of�B�Oj�A���hݑ>#O��wf�E��(E�{��@a~>y�+�Flڄ"�p�3B1�6D|�׷b�r�簾W��w�#�Р@8�	�wf�#vEc�<�^-����{���f�hg�A�Փ^#:��(��L��&���UǶi�l���h��%*޸�[޴�,jr8p$�X�~���ڭξ��Qe�&4"9�z�H�[�&#}Q�5E��1R�R�jmBm�Ң��� �d�
�݉ �t�Bu����xyk�X6���7���]�JX?��]@q#_���O���#d��;�2M� �:�(ښ�D{�������o�4�o�gاԈO�
1�m؅ `�K,F����U���Tn`�,�jP��7Z�JQ�W�34#�kj����R���L١2e��514�YF֊�����j1湍Y,& �GZX���[u����	�60Ci�^��0�a��$��nHӱ�@�vJ�c)X�-Ս��u��+�A!G*�TJ�v��\Fu3"C
ͤ�����,�������u]�մ�XV��1I�Fa�cH84ܥ��V��f5��|���>��B|:��߼��'ݽ���{��Of�hg��7\}/ߵ�A�Ջp8>���0}Fg?]�{�5c�+V'��8�� �D��KC1r!v��XI�{	 ���a?gI��k����Ɔ{�^�32�Lj1��Bc�Voc�FM�`���EE	����(G��s*�J349��F��\�����'ݝ���y��/f�hg�'^M C
�b�+�Wu���@�y�L�L���i̧ǹ�����ָ?"2�eN���sK(�������?����y���ճ�e,,��)`3Js
3)��B����O��:��˕�`hmR%y���-����O�=�x��
�iQ���`(��8�*�Kt( �$l�鹸%(`awdP;��f�9��_M�Y%�Ĥ�9�Q��|�/p���w\gT���W7R�{��\]a�J�>�[P.�K2p�|�F3X�"v�&d%�����)l����#��Ǳ���+^��G�u���$�!=㢂��گ!��(�D��H7v��AHḷ�9�[��/s�Z�:��Ns�x~�-�@�e�L�,Li%��"�=����(}{"|C1���ݠ�\mb���Ε'Dq�5�Q�}��ts*�|�����Qb&T�3'crz�7;7@��շ�2��V��kxq�"������\LhffY��w�|��)}��|��{��5� �p���c�4)�c�Κݭ᫲ۦ��p��L��}y~ý���Ex�Đ@:Fr�=+�e-�o"M�.��Qqю �����AvD��ݛv����-��g@>:��ё���;��B���8�l�
;�){�nr�u���RwhЏyE�R�͚n��d��o:kiF�<�+&��$\A�/E�nv?���QT�I�z�
�o�1��',I�v%�vf�GLkt�MGT�,�0>���ߤ���酎�U�G�x��ti��7v����r��k�ԋ�$|t��)�Y��o\9̈a7#�́'��=���p|��!ܲ�G3/B$̲��|�k�鮡B��w�N:����=�ȀB�>݌��3u���@�*l��g3@v�	f��F��&����`]���v)�BMZ������\�C��[W�jśޞ7/o�~\���˜>D��.�����Oמ���,1���Lʟ8���=�|�FDҾw��x(������@ƕ�Y����y�}@�� H��ݝ�:N���������Y`��gy��L�-1�;�Br��z�
��{e��hS�&���]�<��49�h��fl�Ҿ߬�:�=P$�*=�O�۲&�d=���S��VhG�r��8�9X���
Qc{�{�?@7υ��[�����?53��Ӆ�+���<9�8��㜻h�B���v�s��D�4C��v)�'2썻xgߏ�8�9�٧2�Ĥ��49���dW#I!��{�UvR�\�!�Thm��	N!�E�o�Z�l�ʞ�ؿm�xY�����	�7���Y�X����b;�a�������0M��od�/��,��7��x�ݠ�\u�vz��
ʃZ�E�ir��3�q�0u��O�e[wp`ͱ�R�};S���D�K�1�sR��No�@ ֹ�s�H>�q���y������Nr��B9��C�V"���U�ݍ����^m�V���hM��ٰ$�H�wvhwdI���b�*
��y���墜�n��y"VT}�?(S_����a�Sm_Z~�M�w��_¶���ӗq{f���#�*��f��5#�۴�D��0b���c���q)OR�;�x�Q�W��<U��|eD��W���4)�f��u�cv��n?gy�@Aۀ��af�o�0�2֪è�rx��l<�7�	�)����(]20�C���Y�$e�n�iU�r�,d�|}�6$;ޯ��|T^�m��v�	�=��1{�[T�p[�K��eq?N�<�� x���)O�_մp�{�(�Q��� ��Ph��|DY�½�n2-W�lb�x{.>���2ⲬFtk�˂�,��){�1T���b43kش�dj�ח��:N��;����¥�?�l����x�}qԐ�-�?���X��k��<f�Wa�zn���4#������10UQ�Ѫ�[bܣ
����Ӟ�;ț{(��98��Q%[��B_T��DLTF�Ќ���<'e�⳧��E��r�8j,'06HlTՠUu
�%E�2`֒k$�EV0p���F��w��;��l��3^����r#oxI_��4���xy/�x����|Ϫ>P��i�[��~L�������P�����t�j�{��;�8Ñ�7�;v����{{D��N����PC�W��s��y��)���$츱���W����A��H��
$�Χ���[���3�a�`t�o"���-^C G�1�/l�����}�#���Vx�>��b�g����/={N�O;G��d�d�N���5�&}>�Ǘ��\3�G���L7�!]ެY��A����@(j��w�__ի�IϮ����I�B) ���Z�+�KQ�͵�cZ)5b�h�ݭQ����ʨ�QQF����ʍnUE�\�VܶƵ���Esn[�����Z��h�ܪ��ƮX�[��k��Q�6�V(����s[��y�{��;�,W!�b튰a�[�X�m�+,G�ݍ�7:�[TpKcZs�$�t�q\�kX�4�@�U�L΂顲so[F1�\������$o�-��(Q�����Ԛ��#X�6��h� �B�jV˴R��L���[/�)���%
Ѹ�,5��\�,ѣ�%(4M)J�٬�)FgKL�ӌ̱֖�)od*��A�쮋e��އ#�2������[�]���*��Vm�h��k_/���ɡ��CVTB���b��
XZK3.��#Y03`.�(F�"d�md(�6��l�s(0&�0��(��vqf�v�u1�!+(�U�cE���S�e"��LhkcE.M�c<gX��F5�ah������͊��9���-x&cR,	Ef�1���v
îXKP�5ۉun%m��
A��GE�ٖ�� 4²�����ݬ�n�-���Q�{\V�(R`��7n�PHR���sL��]�R4�h�Wv�5tMq]j��4��
���Z��-�]�ʚ�`D5u5+Sp�w&�(�Z�$�D�*�L�0���hh&�݇;��cS94�.&�޴ұ�G���La�nol�tC��am��:Bii��]f���w9��\mҐ��,7l��q��T2	�SK �5LF�L+2��p*T��` ��c�\CJ4!���V�\C].S78��c(Wm,�if�){Jզ�D��Em��`��4�Z4fqm��tv6�e�]`@��A�[`�uxm+\SЌ7���%������D����2,q����"[is��nMX�NJ�*Z؉vw;U�80��V�p�3PP	kIi�uQ��6�9(.��ձI������qn]�4ƫ ���w.D���f��B�q��*�)u9���])�L�il�2��3aJ��],&�"�cM5�Z�B!Մ��&5�Uf��ffԂXK�T�F���7���,&�sh��8ojv�x��-o���MpW�4:�J--��
��˥,Ɔȱ�vb�����͏6�yU�����%�1�,��t`r�e���j�V��/-� ��,�s���1e%�z#�n6�,'�t��6��(�P��PlXktU���W9��vR�`�ccpB��ba5��ݱL����f�xl#\'��ݗ��m�eC,�5�Q4��M��.�;��
�"-�s4��\�W,�U��B$q��B�� aYkU��L��}?k�M��L[H.K��,ҩPY���N�T3��1���ĀCR��7JF��:~����ޛ�W߹��㺕��y{����eF���Q�#v7`n�s���KW)3} n��Sm��۩� ����uEM3n��[~�x�ڭ����*rΡ�7�{��ZÉp��gG�cۻ#v=4n		,���P7c�ܜFީ|���9���ב�]1��E��l�ީ�q�������\Uؾ��N7��ЪsR���H��_z�=�m?[���?C��_w"�~�	\F��	�=�����X��f�]���2��n�aˇl�4v�yl�7v|7b��av§hf�R,N�0��twG�������ku@�s��խńȋ޴�;�e�(r�W:���!wFB�2�_�o��7k���y�_b����>��->_;'m��H���h"�;���U|�E������˽�9V�z�<3�ww��#z�|c�����v��YR�n�xF�SJa���n�}Y	�큻wdYn*��b{�;�ֹφ�}QnXR�΅R���j��Ԅ���$f���H��݀7`ݑ���n�w�ؚ�ٶ�<˵���{�c�>�����Z�o�Y��L����XMۘ%�W�pM�*���.2��MIg��]L@�A�`ϝw���7cwd�;̶���E](:�ФH9.�m����>��{wgv"(_t<���N�T�����QnXR�΅R���������������[W�i���s�qa�=���z]=�0,��b�Ѥi���o\h��}��ǎX�)�2W}S9����t�7�*�S<�Vy]�����ߧ�g�>����e�W9V�_�ۻcv7c�<q]X*��}��C��N���wJN�nD��DCYӀr�� n�������b{^��lf��7Ώ:Q����;�}��d�r��[J g�uq2��a]<�,��ֆ�˩,��.�m0�+	H��n�\���P��� Ѡe�x=��}����+�kU�U�ž��k+57���{~���ݐ�����k�vB}+D�e�n�tUғ��[	��ߥ�u�_L���� ݍݝ��Z�u�$m.6��r�����-��7cۻ��Ò/\D�f��ۿn������Z�q�m���u/G��o��#��c��7#��(9NBz��+�n��9���;�P:X�|��Q���ڼn�ϫ��{�}��-��9i��M�ǒ�7�՘}�Ԝ̴���٦���|l'����D�<�|�������b�e� 
��;hǩ]WW2�0�ksé�r,�ٍ��[L�o�޿Y��~��v=j]��/^޳M��ح��}WJ�7�|;#ٻ�����Q�9H����9ǻ��/%=C��G31>��gG�v�)��+�.�� cSỻ^���#QNRK5B��vP���N��/�}��t��O�cw_z�&kg۝��wx5��v�w�]�vw+�7�W*���$Saun�	�]�>�����B5��']�=W�}�^z��b}� g@����z��W.辬����W��� ���InR����ؒ԰h^��������{�ϓ�Cǖ�q�rL+IE\�����OD�U|���������%�`��2��eAu�&x�c�Qţfe�&k���Ԧ2�Y^�a�,�%��]�MW�C����L���a��q2K)�͌����c��,�k���u�
0Z�m4]�d[V]����iJK
e26^#�6�HXL�&孵��Ѕ���l�v��PŠŉYT�����	v��1e�;��(-�\5��bge�k��'��vWGR�1�*2�7Aԍ�l%�iX��Է
ѫ�4�������߫����4W^���㓯��qfv�C[�9�}�~��VZsq�#vT��}��էY���gv�\<�dg@�
��ev�c�WG��wd�u��S�"�͒+E���������5�ޔ��m��s;��ʢ�s�7�ۺ�E;Ohû�:��fs9��c�R�W�����me���$�ќɵ)�f7�����v�\l�gt�$���"٭e�L��"\�6������(ʹ������V�`ˬsv�S�Jī�a��3\���Fֲ�V6z1�Y;y���n��(�d��ƶ��|�$��{)�Fl��S�w�d��jq�P�ŎdF�RZ�]R��S2�X:��$v庑�+?tE��,{λ��5�.V�U.9��V�
�s���4WZ��v�k���� -rF���3�nZ��Ԁ�$�$��WG17|�!
��털*����R���ȵ���v��Q��^�mGe=K'oq>�1\���@��kJ֩IJ[{�b�u��۸B�w�LuY��'i��5))�@�g���Ͼ�|����TsոSLR��;�̥,�Z�1f�B�4&�6٦u��Ͻ?|��ϧD�KT�e�8�Ҽ�t��ވ�\ʘ�z�³�5%!%>	Ff�[���'(v��[>ޏm�8�M��OZ�W��f)y$[��+���&�%�>݀��X�K�i��A�M��·���M��|y<w��O�
��U¹B}Z�K����������ߘ9O�e��$Q�z���?*r�k'%��v����z�yk���y$����p�jˋ����>	)��q��%]g�ƮU�/�x�����))	G�I$�B�จ�z�U6Wf<j�f�}�x�oBJ|9ǎ�j��h���ƴ6�B�ś�YbƂL@v�����&�+���Sw�n��~���)�t]�.�{M�:���E�)uK�u��s�%>	)�F]
O��Q������|"3:1��%]g{-1�����O�yr�+#h�[!fH�IHIHIk�������ʮȷZ�<{�Nnn'ي}�	)IJQ)�`�v�u�\&��ݐ� ��Ӣ����s�k��>?X���um�վ���k��M�������\g;���h��*�o��Kc������n�6oL�ۅ�-){M�ʆ�z��wF�>	)	F�kB옳h�3
�f��%]o{-1���g_JP�7:s�vH��[kA��`� Ԃ	4a�f�"�5\T�V��DF��X-�lm�`�l��}����K��7s�Ҧ�v�Ƨ77��غ�y��j@���$��@	+T���o.:|�'�7�C�u��bm�i��O��@Z�-��m��3	u��5�I%a%���^*9���9;�������Ʈ
�Z�	@	)	)�Z�ܞ���ؔ�o\�t�^cs�7��#��,�\�L��͟j�J IO�JRә�2+�09\��+����ؗ�O��Z�$��"�V-͓��}Yq��j+2�b��Ǆ:u�r�{��Fs�ؽ���Z��8ǅXs��/c�����}\����v3����L�O���I��N�����$��vH�bJ�✴̔����u9S��+�V᭿ń�)l�� %#L.��������V��mak#�`�lkL&#��V1��'���΃-1�͐ڽf#�"��ƥ�8]�#cuZ���s2]c1�3+����8rfֻB�ÉK�H�ZS@�iN��K�:���F��@kk���D-H��&��x���x�6��v�����EIb�P�җj�iK�2�̨�1��33X��eX���%�2`4'~����% $�Lft�11+{�-������/i��3T�IO�IX:��jj�ͭ[�Xc�t�77y8X�jμn)-��� oBJ1��6��qn�ɹ	)J<����.ra�[�2]�u�ۑ.�'_^ǂ�!%)BKC�<�lq��`
��~	)����&eo{8[�
�z�Mw;�qr���	)J<R�ګ�H���`+k�67eg7yW���+T������2U��:cLE�����K	`]`��6�{4@���ЛSbW31ÖˀU�;��>	�JR�EN�E�fd۸��ޚ힥�0'5u)���$����B~����@��>���Ieu���X���3ª0���[�"c4����ح�+j�I�cff�vE�C���M�J�oO��w38��e��
�F����و�9���\����!{=vr�GXu�F�vsw�{��m�z IJJ|�q��r��8Y��@o)�I8�3��{�s*��m>���X���99`<r=�R���$�b&p�\.A����}��\��[#_%a$To;���.��GI�2`�xLF�6�tW�-3\�s0l��a*M�;2�E��Q�h�=��RQ���U��j��2os_C�X}f�3K��] $�%	)�HŸ��1iޗ�f~W5OƯ߇�d�捧װ�	*o*��Ɏ�W�@���@I%a$�1�7f���ōM��,UkkfC3���3�iS��8�)�t������d�3����ڱa+Iᾖ�~��3�؇�������͍��VEm���n��i�F�Qyge���3�9k������d>���1=9f�;�$V'�9l%%�~sI^ɛ�U�<|
�x��"O��:]M{�Ր��,��d�:y$����i����^�]>byt��iWZ�����C�N<�^(�@�=�\¸p١��i}�ϒ��c�|� ASˣ���|���P�~��p@)���0f;�Ӝ.�lV���7�ڟbj�{u=�s~�Z��O*���-[�N&B��۝n���!� ���;���S��[��zݻ8;\�ZF-�j �c������ղ���j:'n{}�����W?O."5���9݅�1|y,qs�z��iE�f��Z�.��7�#��������NOoh�
U�]��u�"�W��w'�/� ��<�x�ɠ!_��ޯ�b�T�߽���	'||{����.ڱ����K;���^/�b;S�0�Ç�T-"��;��+��=�df�]����T5$u�g��>ݝP���j�t�ъ�pkCpUT5T.����eX04�FcV��RV�����Ƕhޑ}MzX��VN[�Ӎx� O�<��{;{÷w_n�+�I����Dԓ7UNF��8woS���1�C�2*'BŅ��lee�Z������� 2���cڷ�i��˨8h����;Ӯk��y��s䵺�|ɴ��(��Q�+`-�W�j1�V�\�r�b�*��Z��6����ڋ���lj�wX��4F5sq�F5cV�r��"�ƹr��V�sj"�h�m�j��[r,Tj�hѮ\ѹA�Q�Tb1\�*B�.�wqh�r�%�1�h�\��csc\)51cW,t�#Q�r�gurRA`���ϻ��wo^�������_HJ<����v^�2OW�rI�J=���S��
K���� m��/�P�\3E���r������%mT�'�K<P��6�/Lm>��-rS�%
,R{��ף���WԻi*:�)��:�`lיfo:l[��rPFj��"(����5U*h���8IH	)(��;�d'�J��cM�����w�t��$�%>Jv3�WU9�:����W������x��S�[��
�>�%M�e��ҭF�s��|S��$���BӃf�^�3�Fw8�ܼw1:�� z�$��%]EiI74��!j5��JA�9c�&N����Y�ζ|gF��J�}����^H�ֽa�7;��w���gl^�	�g�3�|��L���&��:�y0�o���C�����Il4��΋WYS�3����%>	@IJK�U�[%Ҭ���4�r�]h�V��j��JBK�nP�w;d�$��n`C�A1E�`4�%JmK�u���U��g���s�h�=���#��V<��}:+�h��'73�N���D�';f����PS�JD_���ӝG�J��ͨ]�<�A�U��&WNŕ��܅���Q:"]�FOP3�ا��䔄��%�ٍ��XO
�y��}i7�2kw_m�]	)�IJPe��Z���ڳ�^Hj�R�5էc�e��cٌ�޽�V��4��(:z���IHIHJ<���Ys���B��Z}��U�����K�%~I�ۃ�cW��Pے:�bN�z��iȍZuxd�|�%]�o�7TEnFV^q,:���Vx���M;f[4��WQ=f�1�f6�"I��Q�3�p�ж%i#p	Z��[MJ��A��Gf����HR��&r���%�ٵ5�6��QB�%!l��	chv%BR2����*�f4������l�Y��u%��L���Z7P�"ڒ��U#�%�ĺ5�I�J���n�-���L3.V뭄�h2��UB�ky�c�l��c��$�F��[q�i�4����� �����`[ZFY���7D%��T[�`�ZA��"K�a�KΣ��tw9�J|��V��ʷisܜ����LFuX���a�q�ϒR� ��*���uN�~�غ|;h�V��W�{yof2��됒�Bkw#�r#����>JRK8�	�c7o&��s3�	[��:�}�JR��g*��-y�j�ë�<۷k�ܩͬ����
��WN٪��fC둛�XIH	)K��w>��+��i��Nnz��le>��ϒS�o�������&��
�34$��}6�]H"l�t��*��˙�9���cUr�L�[	�}�޾��4��$��t��s3W����K�و�V������<�����e��-�M�h��]���q1�f<�X��"�,�qQR`ky)i���N�[n�<ހ��q�	�R�9�6{Wxv{,���'{{ף�����C5ϹFF���n���^dl��>�K�g<�DN��7ٝƧ�)	G�J#E-��3�z�f�4�g����{6�	)�I+D�j����(	)IN	��
��35{4�;�e����9�+;K۪˝n�))�Q���$�P�%&��ɸȻ�}�Uֺ�9N�������gw.���4�3�u����g���M��I[�Xݨ�[4&�=J�{[v�b�MLA�TEUz Nhԏ=iX	)�Tk�j�g��1�l�>�
r�VP���<�y%!%����&�D�
�!7>�Yvʕ��M�U&� �'HJ���B�Y�y}�y��ϩkVRS䉒�3�=��7�vR���s>�7�כ7�Rn�.�^�A�n������Ⴂ����f��Ovf��=��X�;��n7D�ڭ�oj�'i�elޮ��O��VR���Q�]��=��Y#�<R��:��vzl,w9O��3
�ye�Ȋ6�֔��	)�JR�$�^tK��:�}³�������L��H��I%#$�������z�����zU�-�3GM+�j��K��Xʉ��l`v�V:T�k篳�w�Y��J�5[V����X�kn�p�@���{�����r���$��U��m�e���kU�4�gUOP�n�U�N�fq��됒�z�]�>��}�O��$�$����È������*wg)0w8Y�ؔ �If�1��PS���!,:����w����ۭ]�ܗ�8�:��syV1?8��4x�K�:��~�cn�ᇘ�����Љ�ժ��wdR��݆����N)�[{׉��#�<�ӗ#���y%)$����+g�mH��P]��U�n�fq���ZK<"�v�P���(�`�PbE	W�IT5k7bb��LۀfJ�̺+],d������ꐚJ���U����/fu0w;�þ'3�+w]���$�Y��0�]�,DDTˑ���#U�oj�n���Wxܑ���_���rm��z��ܜ�%)@	*w��puOP}��Ջt�bq��(ZK����]��G����w� $��֮\{][������[>��wyǱ��'��y7�t����y%)-j���q蝐.+ov�v;����{w���r}�%>I,O-�n(�]�f�`\n�"]�� Wz-�=�ވ�c:�r�Za�x�o��X�����Ӝ{|/p��]o�t��h����]�M�B+�{��z��� �k*�l��8�[����A����R������jJաc4��1��
*�M��ʘŏZsZ �]�;���l����J�1M�ؤW8��c��)j�;Z�H��ME�0\Wiy��ːΙ]A-�5�-���1
K`(��9�:p���[Ƅ�	uf�K��h�B8�u,&#�&;[�$Y��e��΄�=MT���j�P�����!�m{�e�����A�j\�2�6oվu<���PLQ �A�BdP�^��ןH���J ���L_P�n�źS�8�Op�uWa��#���)JRR,T�J7/#����J���ky�榱��R`�p����J[K#u��7ϥ��v���d%	)ԥ%�+�:��wn3��m��f�ھ�䔤��tۭ�PmDD��x�_����8�����źS���b��bP�mU��%>�J@JR���2{��E��|���y��+;��9�!(IW�����ޥ���=S�	�.��4�f3k3��dp�Ȏ�BU�Si��0�f�0�}��'��P�������1��m=۬�F��ّ2��l7�))I%~�qd'MF�����٭tӫY�6Z?G�֩��^�Bx��6���n2���(�;����5Y�����ͭN7��_��)�辑����ͻS���{IgEE�E������܀�y%)&�N;�����*y�.P�[����Y��#7������vX ��O�ܼ}�,P��F=��]�Vn.�3Y�J����32|�%`$�������A�(�H��w]�S�;O�(z�%>�I����q�`�vp4�����1�n��j��\���nX�L�宓Q&M
��DЖ���$�jR09�O�]��m�6K� ���ފ��%))J".��c�\���[��O��fʾ���m빼��\,�В����+y����7S�wF�R�y$�&9���D���[��n�V?0s�w>Γ�|VM��d��0>35fF�{`�Fp1�������m����j�;��y�{�ι�\S����j z�%>JJ|#�v����osU��`s\�2���W.��:�t�U�����!%!(�JBJT�FSn�nRͅQ�qj�y�dw����ǻ�gwz�˪���	�Faג��6vf	�j��f.��@շ$����0R(1QU�=�	)���W�]t�o�MS����]՛�7Ƅ��Y�� ���9�ƬI�[��7.G�sa�s|ʾ�n\�/8Ol���"�LkE�r��w�;�y%#R��Tmv��6s�Z���w'/mw��@]	)�I"29f�x�m�{ۻ-G���zz�k�T�mF���pK;�Sv�_�y��8A��G��x��C�Lֿc���� ���+٦h#�rۥ�p9Aiڼp!DN̅YM����Kw'�91��þ�#�_�}W��IXIHJQ�9�n�h��ҵ5
�([r��y�[��(�I<�[�.4dN��ho��j��MWJ�1̭J.�\�3	hb��A�&����D�4ET�����|S�6U�G�,��pr�W��51m@R�}�KQ�eNWG7��}��a=�g��N�m���[��BI�VahD��>\�%%)-��1f�L'P+��{���Wm�C�[>�i_�RRw:�s'�EgH�R�fʸh�>�Z^u����$R�BLs�nh����jIX	)	)�V�Ukg}rX7����o��;�[Q��[Z���^��Q���Y���[c2�8̔�9qNQc���1�:��Vs���;�0�~Ge-��_֘����	��f�[����z�_k�-ʄ4�GrL����J�gwi�nX�������O�=ΌV ���Lڲr�D��R;�	�v�x"�輳�a���Z�������j)�l��CY���-Z���X8{�����RoA�#+/�v�Ǡ�Q�2�����Q�ҵ�'aXN��#N��O�WO��$B�*��j��\������cٻX.�6K<��:�&^�oZ�C5�ʨ�V�U�O�]W�'V
�ӛ�7�.��,C�A��rS�����zs׳u
LΓ��;��J��L��=ۚ�Y�w?jL6����>��]���׫��-���總�2-=//j���G>{�=��G�7���e"q-ښ0�Z�UҔ�L��֪�����&�S�R�1���HN�ZZW�qA���[d\߼�@Wb|��yw/$�G��*��~X�o @��m�靾ر��9�b�G�MƆ�=���\�t����5^S�b�Q� %k�w�������$�ۗ��xHJs�����ܱ�l�Lp��vz�Su�صQU�!e��A�)U-8rO�鸁[��}uWu�����^�wۑ���WTY�ᔖ����.��EyNE��=�T[�� m)�����|Lv�A�f�л�S�u�{ܓ��
����5U�S5���*�5:�2� ��ާ@�c�;��W|W�r��x.�.�b��G=4h���L��^��{7����)�}^��G
)���� l�pa�;�ym�ޛ7]}yݷ�v����E��*��-t#DZ�h�����(����`�J61��hۻ�Q�5\�X��i+
��A�)#E�l�71�r��1BX�A�*Ʊ����cQX��Q����\�A��LL;��6�.n��Ɗ�b��QbŴ��� ڄ��]9�h���jK@j9��QBQ��7"�I��j��l$����ϯS�Þx�T��R��6�e���L�V�q\[�Q���@Cf؝Mq�M���6i����ňU	x��������K���F�ٮ�/�y<v���.��G�&5
;Y�h����^�rؕG%��n�)���݋�IDy�C���
ۖ�Q��kFa�z#�����؛��sm��!��J�l�3(,t�h8iR=��[+��KI@�m]���H�X����cMe�z�-E
�lu ���-�G.��P&� `�cT��f�M�[�*ō4hb�iIa�%����^��1cF��C�C0�f�`CD������]�c����!6*�Z�n��T"�m��Y�.m��ݻ��3lvi*�d�p[�E�-��m2՚�0��s�ci��4D�a�����K6!��]7$�+����F:�[�l�0.siel��lK�H�t���V��k�C��[G$fĴ,Xs,-˴5ñ/gQBʶ,uX2f�L�Xm�;@u��(�j6J��b�YP�y���!_1�:��.�]�x+�����Իv���v��R�45",ڈ̛�	���s+�Y`U��� .���+t�C�<ֽe��ǖ&KBR��CI�R�Akؽ�R��͢��1U��m���DH�[���h�-�λf�(�+����kMuk�)�Z�a�d�YD��e�s���kB�{m��8�`�+�#F�=en�]��C��Wf�E�ٍ8n���Ѝ�Wf���Y]ֻK[�J��\ש�� �$��Y�kp��j\k���䡶�`Y�S6�%���]���6�f,SJvI�v���!�j��6)��5X�M,�&�e5����y�e�t.��VŤ6P�.3))��s7-惋E�0R��jK��Ԗ�pK�Ļ$kK.[��P�L�"1��e�H����i�\B�ҥ���,�Z�:���Q ���B7]m��p( bL-�Kٖ.�8q��[u��,�R\W�k��h�e!�FK��h� �sf����[rk0m�F���1�]XU��k-u����6� �����]�	�l[�%ʕ�a�umM���3�m)����5��8AYh�v��1�V�k8���(��e�e�#6�PZ��͆���Wh؄�0��vc������i�m��Gbb]��#�-#S�h����)s蕃K��R��nɶ㊬�5�j�Z���f���ۆ���~~��p�hMl]�fkE�)�3h�:����� T�4"f�P�����QQn����W�	�o�yW���Fw�C�c�9[W�+�$�Y���T��&�P3Q;��vl*�+1�j�Xʭ]ᷲ�L�Yu1�Wy�\����y%!(	.����<3(�b�Vp�}b�խ��}�q�|������>�*'de�xs�]#�)�]M�gq�R�X�����:���Ti��3��s�\���y$�5�B�5�8��c�t��;��$u���Z�od�RK�و�UDi�F����I���<���v�ș�_9�ae��hM����
=�����{�(	,'�4v[�a�U�t�D]gJ��������%	)�K��������i�wTb���G\n��3�V���Ȣ��-����_��W��?-�kC��zɬF�w�CTg��O'Ϝ�I��}
R�X���9ٮBT{��%=�f��f�.��>�$�$����D�U�v�{�9kJ^u����]	)%)BH��q��mΕ��$��ƶ%�x�^*6�ǱS�Gj�W�v{�9�I_�S�������9{�v��u��C��T�*�&p[>ƥ(�I��#��0@��`��4&H5�n���;V�T��c�M�WJ9�-��m���ۇ��'���s����Q�\�6�>R�<S��1+���7{�oX�JBPR)΋�Q�w�)����2[����l����Z�%��d�fz��� v�����$��%�){XC���e�L�f"'�a~�΄kC��0s�)㮬EJ+����6*��.!T0�E����*�[wR�%z��ɼ������V@�OVi���wV��tf�ղ<�%~I$�r�L�T���ǦCZ���G�z�f�b�����w:�{7$'w:��Ǜ���(�IHIJ[C.���<ճ�JxC�1��
�s6ˬ�-���S䦣Q����u�dmPA���	J5�裘���W[�3fq4�ݓ
ڐDU2H���yO4��JpE�z�Bժ�y�dNeN�D��>NS䔀�{kb�Uv�����Y��ˬŏz���W:�z�d{� �0�B*e��7ss��zs������������C�T�v�^pyۮ|����%#7.��=���R��.��v�J�j���ul��7��u5y��n76��9;P��ڽ�Ş����=V4��u�[��x.�k�Q�q�26�q̐���򾋇��Խ��M�Խ9n�MvN���~��Z��@	$�@��y�9v�ݺ��[��J	���7g��%>IGijY�>}O����cܳ�F��iI��Q��l����I��1&M
���b���sX��V�8';�،ե�O-)�O*�N\.����S�%))��_�w6�/#;zG%8&�c���[Ko1閸ul��*ؙe���ϛ��p<�����I����\�9�Y�q�v��]��n��.�$�y$��;�:Y�WgN��ԁ� IH�8k���Fj�۫w޵���&ј��f���R IH	BK��0:�#z�t���,x�eU�0�xul�)JH�Q!�R9Cvr/�É��0�{DM29�F���읂ׇ���H6��̿����	)��,H����3�ʾ�j��DQ�_�=�.Z��:�ҭZm��M�L�s���1�1
<�©�k�%�ꑫ��%ڛJ��clq�Hى��F!�5�$�Kc��ڊ���Íb%�me����͜ڄ�Bm3JM���BB1�Ջ�e�vܢ�pַ�+ƙ���d�h`����5�ѦM)�3&�q����Q����ѱ%��ZE��`���	[-;ZaH�pa�l��~���t��ړ8e.�ZZe5��3�!.�f��&����F���DULM��l{7�X������u��X��}K�6.�o(T�$��y$b��S[I
���R�|N����f�-��}�j=��]a�$�s6/:�iO�S�$�����u�g+T�j�t����k��@�R��>-��uC�Z7��f�y����^�}4 7"G'y��}���+uf/ዾ))�w٘P�����Yj�ɹq$ۚ ��
���}�4#�LO�}??��f�-��ggޠG�8.�6�A7!F��$���rA����PTl^�Jk�kbJ:�$6�$)�@�e���4�ar�3P���Ǔ�>�$6�[t+Fc��k���]��qs���-��QuY&���W��x�m�ۑ^-�ߴ�ñ|��6��ٝ��Y�������W�W�(����df������2����Uz�N�)9g�\�t#}1�+�a��3��_�����D���o��#�V��_�o|RS@��$��ELO`�����r����9�!�B�[�ۘ��R����
6~�u�5{���W���5t��4!��uB��wz�>+z>���y"A�W��6�W�c�=6��S���2��p�������}e����H ���!�T�p$ۑ@��]*��q+#jFj���������Y����>))��D���W��t���4�������Սr�%֨h���Ԛ�G��燉�)������0���6Kc���_��׷4A_��@�|A�-��'�s??��j�rU�3��Eq��ᥘ�fРS�A�r$�܊�m����pG��TOF_�+�s�CFS���\*�7	�T� ��Р[��ᆲz*2�@3�h�}"���mכs�7��R?{��̫�W_
O2oE+' ?dK�l,�#@�Z�P��p��#M�(�w4��z+��`���������&/�o��'�5,Y�6g���Tܞ�W7�I������;��|��?�O�mЯu����]L>�Y0�6Q.��q�͹��������f��1_�:�\ �������������/�H!�T	m�[�y�-"wc����)9��]/��T�s�����~�5���B�-ğ6�9B?�w�~�|>|<����
5`Ǧp�%u0U��K.��R
37$ծe�h,J�F������awP�ۚ7�2��o2���6k�w}��z��v��eϒ�D���}M�n=%�>�އ1>�T�׮�<A;���y�v#u�2�[�>�H9���E�wXU/�~�"H�u�nh��I��t��Z~����sU8�J��a7��>SD7�B�n'�͹�u�Wq�闽3�������h[���̾�����a����
湢0M\/�9&���F�5�*��V.:\�m�8͝�X���y�l�a3:�ь�X��nҌ�a-� ��n)ź��䯇��J���%�(�H%�>�ۯ7�����8/w1����hd�A���g��ޜ���P>)��#WP���7!�ق���Ǵ}6,��s~:�#p�� �r���[eاg9h�l
]�ƹZⰡe���~0�{�A��"A��6�ds�?i�����DZh�էr�}o�G� m�t([�$W����=�~�_��S^ ��v.̾�����aɮ�G�uO��"Hm���C�n;�N}�A����B�q$��э3���(3#��ǌ���W���
p'�j�n}MȒuB>�����˚y�}>�vH�C]U�܈��r����
~�RsQ���|3=L��q�uܮ^@�Nx��P � HmТۛ������QƲ�p��������̜�����v��@��4A�mϫͺ�	=�Z>3c6܏�늈��u*K�ZY��ѭW��UE�KF�R9��z+x�L#�T�F�q��Մ�n]̑�=���n�|]��ݓqv�h����l�bĖf_���[	�0�2݃�;4k�6�WQe�SE��zUt&��F�0��Cdv�.��x�T��Krܨ�\�cB3Dqz�J���a]���f�Y��U�s9�K�M���˜�D��ŋ�y��l�j��W-���n�6&`f�eȆɲ�8SD�
v��5tͨM�!�aR���*�f]���<�J�n�91m��ef5�bCPK�����a)��؄Q��vK�Hj&��l�J�&��kp����4�s������?}��~����A���������g3Nb��O}CQI�@����Cف� ���� ��
���l���U�\Qc��گ��S�!��#��T��|�{�9�u}B�[��;��}/_dc�+xW�}�D'�(�	 ��W�n}A�kQX�V���577u��9���<���v���^)�y�"A��y�B�n$��[��1+�Y�hW��$KnT�._}y���|3�G�t	#���9�灂�������m�[s����M���/U�P�ѐ�B__�W���G��o�>_9��O� ����O��뙎ph�F��\���&��Ʊ�۴��tWl�ZuHhl�RviZ��B&�T�p���?(AK�͹�r+�FgWN\��"�*s�k��*�G�WgD�U��3@���Gs�W�n�x�|A-��E��m��vd�a�p�b̄*�F�+�;����}2g�ٲ2��>�ԻHw�B:�L��9�O��n�|ңJ���5]瞷���.A8g/��^򚝆�~�t{���)=�=��}�n�����+�]#nP��L}�}q�2��$w9{��܉6�W��t"�ƨ<�H��_\���5��G�>��� ��
-Đ|[s^!�@P�T���ό��pp�M�d;��]4-ț��n����|�<���v���Nb�!mG�fqȎ�41uW�'B�[�[s��^n:3�ϕ�����u�׬K���Wۡf��W��yt	��Qm�r�>�{�/Z������j��#l5G�U�\M����ڕ�������Q�}@�����Cn�x��T���ݟ��^U�(�Ѹb���g<<�
=�$ۚ6�P-��8��4��/�L��ų�}"o�q��ӗ�I�fWõ�(s��"A������e��6�W�tH ���hۑ@��nd�}�Ol��G�ss�򲲼3���.y�:�eO�7ik#V��w����5q�y%w�wDCh�|�μ��kٶ 7�;�m���9O��y\M�����C#�y;�b%hZ��P�o%�����{a��>�鿺��݇�R-Ƿ߷��^tޓz�ܰ�w7H���zmɾ�5��1�֌�z�y���ʷulg$�U����%��j�l�^�S�@(�+�{�./=��h����b\U�۬܁�ảtя]� ������������S�9��H�k�\r2�o��zEw(��ڄ������¼��F�#2��� w�rø�����3�L�kGǙӛ��^��V��}���m�	gUR=���I/K�<��v�3�ffݭO��bw������|�w���/y�:^ƶ���+�u�P�wN,���g��؟X^���Zλ����ߎk�l�6f��T:ۻ�x�A����0��8�g9�<[.2�gт������k�����Nr�|Jӈ�2�G�؆pЪ�4���9}��'Ýۖ)������;��&�o���H�/�Џ'�u+�X����g�i�#��X9��Y�"�Qt%�ηU�L<0ᇮ���������퇗{��;l�(>W>�J��⩢k�]ʜ�O�fnv�����6���an8&�����Q��*��,ɣt���تCA��^В잯�F�	��A�5:iݡoNn-j�����ըf�m�e�<j�v��e}���N�p�����H�,�9��$��6�;��fQ�Rh1��!&�i-"4Y,�,%Q�"I�*B1Q�dĉb"�@��r�QcD&�I���I*M%2��IFC1$I��i5mX��I�$�M̑fjLA���4�)%&�Ԕad����PS#�1IH��$S#d�C&PY�aA���A�!Nnŋ0�0F�jdB� D@I	dЛ%�h�Eѩ $,&,�M��f2�D�w]�"#D��T�2&b����@���̱I4-�1�F̋+&�BN릙���h$BA$� �x�-NiI�Z![:��]A.�@��!��!H������۳��R$>�W�mС9��嘆��W�A��|&�٢6b���ع�.I��Ϡ�ӄ6�P-��Cn|ۚ��t���`�h�� _.��Nr���N�.����9�A��u^!�B��~��������
|�m�D-����20�m�u��ψ;��@�ɴư���̹���������C����x�|A-��4uj�}��Ծ=��|��ݖ>I@`@��wM AȐCn���!�^�}�xW�n���`�U{~r+ӝ��|%��
����(���ٯ����u�r�ن8ښ����� 6�`�5���^J�}Nn���g58��]|;\��c�!�|Cn�^!�B�q �n;�jg=ʅ�������jO���t-@ޥ�������ݣ�E�97��jã����'�j&wb[0w�0�;�5w}��ġ���-�'�C�0d^G�;�]�jV�b���k2���|ڦ���!�@P �����u�����k�F���!>�7��-�*��R5M��D�Qn= ���8�b.�������b%
�t�x,Y2[GGe2�"�KLe��M�5A��-���x���hG?Qb?�{F����Fuȑ�.�����Nk����k�
�Aߝ���'����!/��Cn��I���L�Bf�E����s�:�.�}�N��Ծ=#��]B�nj��0nM��Gs���PnD�۪�M�5=��~���������aU7P��� �o��r���H%�4Cn�B{ ��w�[0}�P��9�r$_��lwVv|�5��Wõ϶���v�8��T�^#��x���q�-��Cn� [���o����~���
�'��~�GQ8��D�:�I5�+ŷ4n�q+�s=�sdnm!�Ƽ��!�K�MD���cnl%����{�!�*�R�n���\�wZ��'p��d����]��m�"����6��X�B-8�9�AX������;�4�Թ�Z�f#I��ո�Q�	��:p&Hf�n�j��ClʱE��E�8�1e#��q�75fG.oZ]i1���e�=�ib�;)"lI���p%*����sGn��m��3e� Z�m4D"]��-cDs�qw6:�6K2�+��i�K]�u2��)\e��;vv�к�)4fH�%� ,`�c�w6����~ė3�2�!\�.�n�X��K�&f�Y� �xE��%��$&�}F��s�� ��W�n�Ng}?\9a�7�4_������sX�p�}�J �t(�npۡ@��Hj����q׭��~�O���7�<3{�:���fr�����k���$6��|~�.�݊��$~nk��
��Am�mƣ;J�#S�����u�g�'�ؠ|-}B�[s@�rnD	��w{1W7ksgA6D�tx��W�3���}�yR���|�}�7��M<��q��9��$)}4Cn�[�$6�W�n{;u٢�ԇ�/>s����'.�v���ϫ��"A��[t
�m�T����z��XJz�~p�+LX%[����cn6�ee�-љ�K4��K��3��������<O��Qn'�ۚG�V���W_F�1,�D�>��_tw^�װywP�ZsD��
�����QW</e�����)����GVJɖ�'����F�G8��K`�	���$���m�W��"�1��ͯ_q�-�(��|d��#w��u}B�3�?���R��:��q���4G/�Qn:��O��p�;4�Ǿ�$�
-���jEp[v>��.����$fk�����S���	I�
�D�۪��[��D�8��Pmh���J'�(�A�m���_���Q+V|"��W���B^��� �g�/�4!�Cn�y�>�܀�,����o�B󏾡B~|��
�����/��+�~�ܾ�7��3��z�5>��H�4"j� �K؊&22�p��\��rR`�Y��0k���h�\�m~G���	 ��y�: 7"E��ӕ�o�tf������<#��l\�x��P!�Hߺ}A�^n=��5�-����t� � ��:6�O~\��J�|"��P>:�I5�
-���]���4vH�״(S�nD�ۡ^m�0����\|���ڈˌ�X+c+{��n7^`��Wf�{F���Ӱ2�����Z�"��0��x�l�`*�B)ue5���.�{�|�}�	�����4�A����	ߗ�	}��ԠW#|~Nh�܉��|9v���}�L�|;{�+����WG
�r���������@�O�sD6�P-�46w��^���M����5]	�g���\ 5�
�<��������� {��\�vKf�غ`�R�Gy�f��J�԰�F�7/���q�~����_����W�mС9k~�/��~{�~N>"�>ˎ�C���C�H���� ��mРAn�DF���D�g���<,Jh��D��M���s�p�Q3����n}A}"A��m}&�|�c��P�{�A�?��A�n��g�>-��(o�Tu�����:&��"V��Ew�� O���۝ ��I��ޝ������y�>�D�9��ۡ^��x��b��=�q�k��})���ep����fT�-˼����W�+7x��(�$�C:b�ї�a�h�m�G��LS<���썦��tsdҩ�!6��^9ݟ��\zA��͹[� �ۡE�5�����H�L=�ng~~�����@6���Cn�x��k��`]5Q�<H�DU��m�]�I�굤�I��ך1DJ	��4	��sN���(��ۚ��Է��蚯��Q�>}"l/�!�d�]�0G۔(��k��$6��-����IY�S��Ƒ��x���	�[!����OnTo���������-��ݹ4B�sDvt� ��$6�͹�nB�y��o���ҡ�'�<݋�෠��÷�|���+��>��
-Ă/^''J�rv��j��T(�D��[s[gV/����*5o�/�	�Aw.����j)����m�[s�Ȓb8�wX��p~�P�'���	}�>v�ܕ�8�M��� �_P��O�>-��|g���ŝP��TiR�shb��Iѧf	E�f���;�[/nr�s~f�ȷ�W�{Qž��vxN�٤�vћ��U��ӸÝ���!�����b�b�6HE�4����1-sM4ι�tX��eL;0Ɩ�D�)v�77GY��٥�ɜ�&X�Y����,K�9ʖ]kØGB��rZlg5��tD���*�li#k�K�����v�W�Iff���Lc	��i���;"�)�uv*h˔kK�Vm�r���V*�74�c��R7^";JhK�,�,��=]b썄3���B���ıͶ���M�<E�F5��A4����d�f�Ͷ�tn%���F�Y��~���~��A�r'~�9v�f�[����v�ӵ�V���g�'�.����
��Knk�0��348��)s�'xW�dI����_3��˅���
��C_H�[s�W{$���:�ا�ђ$[��sD�I��x���\F_d��F��}��[��~�x��)�G/�P��A-��ې{_L�P��ʿ��� E-�@��� �"F�Gxov�n��L��;{�J|ҁ��_]AcHm�{{�P-ĀA-��r(�oq?�D.����K�˕���}nZ�ſ���\	 ���E�5���n�Ϳ����M��y)����VS\;�#-��p�M��#Y`$ѷDTEA���Tf�@���wH��t#)l����[ƳeF�8���̣0�1�u�˹w�s`���У�A�4m�p$��ܻ'숭����_L\�w�GaǼϥ�r#���hʼ�����w�=۹F{�/E��LuW@ۨ�)Ƶ���O� ��;<9lwmF���"�w���
�Қ/�H!�n�I����sbA��Pmכ�g�n~�1;����"������j#����(���(�׈!��t(&�:ڳyuS��5���6�W��l���7�6�/������^ �SϪ�N��h8���ϛz(S� �ۡ@���Xfa��"|��v�zj����w)�M~r$ۯW����{�Q8 ���%ڬ�͋ى�R�s��"K[��њ��b8��Lר?�> ����B�"�[� ����C�{>�韚�������Q����mn���ϵ)�P!)�$����+���>���|�
�]�����&�Y��~[A��h}�}^n
����{c��;5�F.���>mР[s@�܎�j�����_m���M�3*\ɀvPK,��Qླྀ��b�ؙ�˝�Us�a|WQݻ9�oy<}S�r����|S�<2N�dӑ��wM�M��������4�"|Cn�x��
�n<T����N������t(�O�Nhm�K�{>��r�5��K���Ț��>1�x�)�wH�t+͹�A��B~d^|�?|�C��Cw��m꽥�c���O���� ����iͣ>2Eج���5&��i�͍�V��um��X��I�dׇ��k�]��T1��	ߠI������N�}]����w�����=�4����W:A��H�B��x��B�[� �ۚ �RZL,��G���uD�Ak��m�w8�����LLb�lw/`I��W�m�����#�J���D����?'>�܉6��t>�Θu��7о��]<�����+�;����o~����(�H>�4Bn�B~���.�~��^?w��nD�J�8�����Nl��;���SDo�3�}�;une�fu�
��N���f���w���x���Z��J�N�~U� �":�ۂ�c><��׮/!/I���:�cf�e�co����}�C��>�7�����
�n;������;��9��U�
������_דI��_��<�'���(����l��8D�M������<��ۋ�J�,��*�����&]�]`�CK�r��f����z*�z��� ��D�۟SN��{A����cJ�N���~]�Q��*x���^)ĐAm�ۡ@��I3����g��Ϧ�A_H�]}��~�_;�q���߅{5M�@m�����k�;*��A�O�r4�Aܟ�wӕ��v��*-��V�&��2��ޠK�A�E�5�
r$ۡA�v��~��{���"@!��^-�skh4�V�1�K'~͏��>�VL_��4��%�4Cn�@��H ��B�[s�M��V<�AT7-F��?^�������߅j�/���t�=�W���:*"[�!��٧�ںy��97u�l�{8 ��r_zm��<.��u�9��_>����W�� y�^w�H/XvN��{#p�ҋGf�mN��������J�BY��S�?vmM���`�4�7��ə�t��7�7;n�e��/7�䏬�{@�\��C��0�-��Ǌ���G_Y���������WN^���m�~�0�h�۞>8�
�W��=��O�=��M�k�t�D���U��vb�盎-�ou�p�bZ-�Q��Z�O�'Ϣ�x���{����n�NL@�VZ��y$*^٬������-�p�\{=v.�<��:a�#a�����4���Y�,����hk�o�5��¼��� �;�y����,x�ne�n4�}缟����n��u^�pLC=@���揠�a�?j����!�=C+����gvu?V/G��}�XX�O�Jq���[�Ƒ�Ƞ{��Cq�����Y$#Q�Ş~<u��v��t6�A�a�F72%S��(���4c��Z�J���E�4�Ejh���O�bR-Wq��N���	�H�N�I�z�<u�#���<��::�~7�N`�ͼ���L��0�i��rOt�_I9m���N�$����4��3�*阂a,��w�m��S�N�㻒����!$to�q4n�1炥Oj���C���U�9��M���X�0gEA,��:187�H��/�'�˝ۊ�O%�ln���pic�I��/c�7s�d�S{B'���ڽs{A��ғ�$����e���Ch �4�����FL��i��IE ���H,���a��! ,D���&
3,RJP�dB�$��&)�))��HF̥��"�$HKD�S@��) �J�&� �!�"@ !"0QR	�K�B!�0�K��@�0A`�RD��1� ��(��"�)(�jL& HS�rchf�d�HR`��(�5%�!�':������d1&Q`ĠɘњE2fC�")�]�i�	�	-`�"��@�&$% $��ŉ3ĉ�bBM(����"B`�d2�$JM$@�A��1DF� �rI�@��绽sZCh��1��K��۠�	A�+�F�Z����.�+���1�[�dF�e���a-�v�JK��W<�ٔ��tl\M�HԎ��l��xH+\h��2
�.�6����4���[��q����b'[Ç�h���؅��
�bŹ��$��b(;�k�솭&�\Z������+̬2jA�hݹLMp���M���h�̈́e��6.Ԏ�SLP� �T��Vͥ4]�V�n�0��\�VY�Ґ5�EIWj����un e"�-��˧����q5,��Ų�/������p%��Ti.��32�*``lSRV�-�S\8�i��"��HA����0f��r[E	x�+��0�e8�W@qS1�%[J�H��I�v�1��M,����h�!�����5u�Wah��&�� ����b�[P\a�&թ�.�Yv5��#�ն�AZD�JK�o9m˥fҭ��:��4ibb�����`l�m�ݕ��5�Tչ̢�m�4�h�f�j�pR0��jGݦi�W0v(n
Ff\���Uf/1��ٰ���0, ����4�L�K�v�KTl����JM�i�A��Z�aX�kJ��°�,q������X �̡��_����B��"�Wi�����Ňc�)]A��v\X�4ce���)-3�����#�0�l�Lgj�36[JpY�*mm[P��.o$vܰJ���=V�qb2�-�=�2�*�ѵU�P�!����djG5�Bکu�s`�]<l�!����3L�e�@�n�[�SL��a���.��׳��Ƽ�t�XHK.5�vex�S&z޼],�(1s4*l�r��pĴ0<n	j��4u��:��i�n�^6A�0�a�ѳ]�rXLmѶŅeJ�.�f4	��ir�&� j��H��f�,3@���n���Z�6����i��p�9tƮ�GK�4Kإ�D�F�W^��)�v&xL�h��JchY�ͮd�#[)��SD���U��\���v˓Rk)�)v�c�3n����f�emlZ�8���Em���RWJ�ƒ��[*���"#r͛!�x�v�l�g�ō�;��º�u��`��le��3��mƂ���֕.aw$ՙF��m�@ �WSB��Q�.M36�eH���k�KV`�k�h$M	r�1������M4b[�:�����<�k�n�`�Ζ�r��>B~�ɉ2�B��.�t���0����j���م�lV�2�^�
c�x���/ߨP-ĐKnj��o�����%]���ޡzkA�����DAW�
��寮A�m�nh�Ň}6�B6�W���[A�ڷ�-)Y;�l}�����|�P�S��Wj��dף�P2��Z��� g�t(���PiU@]_5=q��aT���N�û~�j� ������nE�I�[�������o�j}]�B��H%�4)fF�;��.[�yH��$�k&�<�}_Y�k��>�m��ۚ�H!�3�]^�|�{��7B�m������V���7�Mx�>�Т�O��s�ʆ=�`��y��?������:�c)l3H������4�a���\�ڷc$ ���_�!�嘇~��^mΐ[�>���ގϢ��[y[����,7���̑k�r�:�Iw�^-�q |n}�u�2�}W�rn�&Փ_X�Yw8%jZ��-4)�'s-�3�hk�)J�65��-��l(;Y�@�Nq0f�ow���*�^nj̇�]����镆��u}ٗ��W��^j ��P�۟��f
ٖ�{:@w�(ۚ ��H!�U�t>���5�~J�g%�l5��w����l��
-���[sD6��=��8:��Ar��N���3�Y���m|ͷ���������#��(��h@��@W��:n=%�>m��[���N'���ֆ4�\�_����˘B�+�y}��	O��nt[�����]��[8^�r��Q҆��Xe�nXh�H�GK�́j�ttכb	��Z�������~�����Cn�{^�+��o����߷c����v���3@�-*�zKn|��P �A
�겛7�� Rs@����/��s�Y�6���ó��j���!�W���1W�����#�H ����nF��O�s����G�j�l^�C�<3�"-���W��L7'��&�GN��i+)s���z�圄n�*M����8�Jp�O%��7hjT�.T�`�����'�
 �����	w��S������4>]"A	���t1]m3������������f��CA��]?H[;��Ȓ?|���An�|ۡE�/j��9]B���,W�$F�x�wl,�n�s����͟���Cn�x��(߯��!����}����X�۫��E���d64�be�kXg'Z�j�\SU1�"+�:�>>_)�|�
��[s^��p}�}y��q����:��$Xw1[��@@E��Q���nD�ۡ^m�#�������eW��}B�f�3�/;�-����l}���f�#���R�q�1�u�VT�#yȠ{�I6�W�nk��Z�ٌ���2s>SUN���O)OTcw[�Α�9�h��� ۟PmТ�O�����JP�ߧ�>ݯ>�>m�R��?}_V��Ƶ�_P'T	 ��ᣭ������?�ğ7�^>�v�Y���]��^��3P���v�g�*��WjO�y���xf�O��ا���cS�#a%����A���^m�[�$6�d�H�gJ0`/H�T+s7)yy�YM]߷c�	϶h>�Ȣ�I��ޝʧ�ۧ���&�L���H�	Q�L�� KZ�ؓ���c�P"�W8SlZ���}����)}B�n}Mȝ���}IOȭNk3���
3w*>4v�t�G�}MH�x��
��-��NCv��q ��5Hf�3���nmױ	���	P�nfz�"宭���D	|�@������Cn�x�ۡ���|.�.�ګ;�x��-E�߷c��l�}�E��-��ۡB��jOٿl ��u���Hn���g/����RN�3�˾��M��l���1�Q��'��s��w�q>͹�-�q�4��S��s��
�ۏ�����1�b>��^J��5�B�nh���/:4�AF�<3�2!J+s��?��
�y'.�O}6ľۣ{rF��)��K�����v~��+/:�.3���̺�ǌgyE4 ��}ۉ������p肤���n!�E6��.�e��+X��K-�;A�13����l�RuɢMX�uh�΂ոL���l�]ZJ�ՔW#e%�\\��3(�2$���;D�bJ�nZ̄#�Ί�ZG�rpaF�&ҷp��U0r�
V�a)]��1���-%HS�͕cXY�R� �5Yuaٴtl�6ݶĵ+��Kl��R�`����2l#6�*����6�1ȅuŨmr��	��Pft
�g��O=�=����G���W��t(b͜K�϶���Fo�c�;Y1����|7�B�<�A��Cn�@��	"�7�ugnC�>�Bp'��_j�~E|5jw�]�zҟR�D�ۼ'�}�r�b~ܾ�^+�H%� �܊-ğ6��s�?�q�$�H�o�4ʭ���k�	�#�R�> ��y�:n�Cn�����sw��9�鉟7 o}�6�V,�|����:s7�� ��f�载���KB��I��!�T-��A�nU��,�ҍ*dH
_5��c�e�y���
�SD/�H!�U�܉��W��<<{��X����U2�3�v���n����pv��:�؎�����~B�_�������zAm�z�����]Y���m1	��bm1�^@`���@��[� �܊-�����Y}{s$n��������Q����ZEé�:
G3b�.6�
���:5V�0�p:=�8�"�B���hB���S�R����rU^:�
ś/����m|�	����N}���
����C~���|��G�O�V� ��mכs�nFI_^���~�Q�������[-�χ.�P>6��!}A��6�P-Ă(P��2�#K��F�Т�H ���
�_|o�2����#�<�|R�>"�����?��p�����I�nh�܉��H�g�5.��G��(P�*jfv������A ��4}�^��-��El���5�˞7�z�"&��5@�U71�g��3)5��:덡��enr fٴt@
��_
P$���[s^!���S�G�[?Q��χ.��o�0d\���������q�nh����<\8�>)}2��_|ri���YL_	�#�R�%?�P-��3������-*��4>n@m�ۡ�W?`����i�zx[1wl'��ǺU�-8B�e�.�P��)Zϼ���M�w���Ϙ�C��dZ������)�[W���f�;�a��J*A���/z���w�q���>��}�7 6��&�옪�k��,� ��У��Mx���.���~Ϭ�L�p�P>7�k��'؊�Iↂ1e
��P��H ����t(�ҭ1x#�|����{��5}y�VK�r>\ ���ۚ�7gc��}�����߯=V�d��uխfuJ.�����݌�,�ŷ*6iҤqZ�J�W�>���C�����>!�B�[t(��YN���~�|�|����vY���ϰ^�
�I��mר�	GLP����j>���7"B�;�]�}gZw��P>7�>��6о�g�e{ ���x��zKM|ۡ@�A-��YnL���lG4�ѱw��:���y��p'�/����7 6�PUp~3��ߟ
�]��l�o9��
��q�ܹ�d/�ϓ�|s>�"�x���2>����]�2�>�u�F�R0'�0GH�d��sbt���k��:�a�Wo��׊p�Ł̒.�5�j'2]�u\��B���G�H>�t�!�T	N�۟6��7��q��z�D���9|�~�r1ŧq�����ϫ�"Hm�x����k�|���cٵ5XcIA�h��KZ�5��a\��[M]A&U�1�.�4f(/�> �V�׈>�:��zAm�*�K��Em�}3���K� ��*������{B�??��!���-��V3��X?&(���+�}�(<������%| �|�|A9�Mx�>_P��:ʼ�U�hX?}sD_�O��>mР[s�ș��8��
$���gO��mE'q���@�Κ �>r$۪�mТ�O��:�{֍�S� �T(� ��涮��+n�>���_}@��H"���ӕ�Ti��@�h[�y@����I��[�B��}�=�+�ٱ�,�w�(���8�Ng�@�����H ����	Ss��ݳ?�0y_���z�C���ʄvOQ/�1_x,�xO�*�!�s��f���N
[x.n��r����н�,�dLG߿;�ϵ�J�)�V��G�.��M�K.pg�K����Wm4ۭ��Z�0�,.-���iIC.3e����e�
jZ�uڭ�5�9Ơp��K������,��(7Mإ ��:�.U��2��,n���Da��p0�,�i��)��u%w+���6��s5&H���W�v����Fbb�V�Z#ak��5�\������m3�(5�6�5S^ʲ�-J��	�)�ZY�1���1SF�p�_
��B�Ȣۚ ��s.��Q��]I�g��PY��o`���>��~��n|�0A-����\*����>s��6�q�����2_	}���	 ���[r�X��ۡbX5�񱣪D�1:�|_9�A����Cn�o�'�u�c(5����l}
/~s>}Ng�^ ���@���n|��y��}�&v��
 �YB����܉��7�{�"~%'y?�#��D��_S���|�P-Ă�n}A�B�nW�>����h���{���ì���}	����j��t��5�r�=�~=�T-�pX��ʋkl�ѭRF�skF�![,bKX[j�o��������A	*��
W�>�H�yg3�T�_gJ2"�w�>^K��8�A-���u@��	"��p(�<�>=�kɦ��;�CWJ��D޵�r�:��@���ȣy|r��ܴlC�D՛'�ۺ��l��g����h~r'�v绢�|Jי?����D/�O�m�΋��U7���=� ��O�ͺpnS�v���_���h�7�a��H�%�½� �7�6�H>nD�۪��M��}N9w4A���C]U�ۡ@+�&>�o�W�
9�>��A9�M��p�YG�DB�;�$��MۑE���t(��h��T�>�������g+���O|Jי<oޠA��� ��y^!�B���كq����)����s�Hm)5]��������1|�c(�&�X�K7[�@��1U"��O���[�[s[��ô�U���$~���Y-Zi�~��3�<��x��>�܉!�B�ۚ#�P0���v��B�AV11}|b}���wG�Ϧ�A/�W�qO<�|�I7�v戽��p$ۑ@��7# ����g��n&)V\��o[	N�n��M����0�{� �z�mh���E�W��o'�}�����A�f(���-�_��ۛSv���{=�T�Z�0nk��{	²r�]�˄��&.�e�����Mỷ�3=<���5���|�Lͺ�I���+{=wգ�ĳ�צ_go�z[�w<�&��x�ێ�/��gd���`9�p�� ө(�����ܧ������f!�{OR����Jܞ"3�Pʝ�eɡ;:�M+[*��9��hӚ��w��DS��;�����og���B3Q�*��p�sJ]y�����8Z�@�k��gDᷡ��I�Ԉ��TWm:a�=#U)y��嶿G�[�4T �n-�nB��-`J�,⽥�}�����X3��H�������������wv�iR3��ڑd��ݡ!�)\��60�pvÏ�{|!��%䐻�R-�k��Y�c��/��1��h�����T��ZU��T"�K�fLP)d�+���|�����'�����n6�C髗�\����l��T�;��7eZ�u�S��!���<S������C�|p��>3P{����u�����羉)n�����Gw�������k�3�r�ߏ�{[�"þ�ע�K�w�p������yE��$������Ov�/,[ɐߴb�KLo��ݫ�J�L��)����)�<z��xf���D�i�V
o@7U��}|��-�����[��j�}�B����/c{�d�G�ӌ��Re^~����(<����z������434���	(I�fHbH�I��
	
Qba�Ȕ&0������	-3%$�[�fRfHƆ1���)�HD��H�"(F@цĔ�JBM�#�*I,�$�$13�̑ �1���� �fS II44�	!
Ld�!;�B�e��ab �e�E#2"RH�M4FE��I�Sc�d�)���h�#$�4�*B4�с���#)QJI-���1%52F�HFI$F%CFhD�fB��,ӗ1�I&B!&��%BHL��I���24�Ĳ
2dL%0��JP�X�c$�X.�fJD�H���ۧ��9I�|g�+׈+��>m�e����;���~��&f���G�H �潼^��u�����!i�K������@X.;;�����}@w�$�܊�4-��>����|*����(��0��"�>}x�w>� ����x� ����B�N:��3x�[a	��,�q�0����X:��@@6�f� �!�,P>)@���y�:!��/[��8�O�u��B�T�:nz_�>��H#����mТ�H>m�-5w������C��]c�B���P � N��(��(E|��0)�+�>9�Ȓt+͹��=��e�&.��4������> ���׈?/�W�q �[sD6�����3�Q�� q_�W����?2���꾳����~��Ǳ��G������p�y�&�r%
>��z�ҹ(dG�چ�j��up��}��K�u�h�p�-�7NT�LL�>#Z�W/�W�q ��4 6�P���=/�1�u5�'��U�2�����/�}��#~�[s@�܈��4����&�x�]
dl�	.�x�@0cKͅr�&�ui6X�e�!�M�g���������ߵ�^mȧof>�_OI�_i�y�t|{f�"�f�}>��hW�D�Knh۪�I�x�Ui�&
�����H��x��u_a�L�y��A�s�9Co{o轜��&U{z0����>mכ� ���a�n�L��f3��2�ᑺxK��@�;�P�[s@��>6��5M��P���_�Ӥ� ��������)}3�Z��b������s>���_�{镻���P�~�$��W�h��(�I6�P-����F�1N~J%����_�]W�~�-�ς��W��� ��O�m�y�"uom��f���[;H��W=ʨ�0d~>��:�K��ٝ����b���%��š�Pw�9�^���mjg�2��L����1�V��	O�E��[�],�f�0�NӘM��彲�.;Dy-mS���98���a�Mj����T��n��2�$�6l-@��0s˙�aک[���H�,].�:4�E!�p��)��k[��YN�VL^�ܖm�\�["��T���V�6Ǵ��`z���ve�f��̔M��,-�3[X ���ոj�����sNnH���nLM4H�k���|�!	��r�ŉ�kL]h������XF��΅�4�Z�ͩ�SmZ5zj�~��Dg�B'��F��jZۚ��}Y��}���	}��`�_i��y;ˠw�@`Eg�(��h�܉!�B�ۚ"���5N�v��0���^#_P�;����>��~'g��� �Ϧ�w΅�.�S�W�Ha�sD|��@��� �܊ ��>nC���xN���#N�}��^9�t�ς��W�)��ȐCn�y�"�[�g?�r����E+�� ��
?}�ny�]X����Fh�/���	O��_��|>�Cn�Ss�Ȓw��u�Q�2�W���-㦷��tU���Ϧ�F��(�A�m��{�i����ϟ��p���Mt)�l&���5�L6�ꃸe�Y�h:�<�0�f5��?z�=��'��ǒS<���:/�>�s��.����A�'�2�|�H!��W�r(�N�y|�~���G1��z�,���\MK�K���1W�O;��GjSW�
~����\��^�I��ɯo�Cçu�s�f��E	>>Jw��D����W�Ώ���!�8�՜.�����u�>�Aߺ�x���ړ��D���B�-��!�Cn�ŷ@���7�Q�w�_���4ƨqI�s�����|s>�W��B�q �[sD6���|]tp������B�K�nD�/v�y��ݲ����<��#`R�g��N0�w���s�E��A�4A:�p�F�=�wR��O���n������
�H#~��nt�܍�� ���_�5>{�������nu�%�{a�d\&�Z	^�5����-�vt�|����q��ܐ�����[�Sn�{�:69�O�>�E_����s՟�*N�b�@�A ���u@��I�S��>����[?�}̼|��3n^k>�G��s^>rn�b���>��@��S�A���Iŷ9%G�<���Я_�;'o6e�LI;�T&׊�N�p�&��nNاK�.���_�����-yk���P�w�Z��*E�>*�����VD^�lܩᓺ~���I{�͹�AȟuC��qYunl�]X��s� �6D����[t+�ΎR�'�T�_���Οv^0:U��G�ﾏq|�mРKp$�ۯ6�k�#qvONep"����^|�8�7"�ֳ���}���|�I��6�nS������^�� � �$��9�E[���<�_.�҄jd�fzV�8*�Q�[?���!}�@���
-Ǥ��.����39�|2v��_H�5�֮E�=�C�"�nh���P>)�������b�,����}��;-~W�uLU�t|A3��{�[�� �'����7>���@��I�B�[sD7 ��:F3O�x�*���y�nE�g���@����|�O�m׫͹[�#n��������^ ��P�WG������)�i�okᙶ~��@�Z��8�o�1#�zћ��*m������e��*��+�iCJ��r���{uw��UC�,p�[	̊�Ȫ+n*o��?/���D�ۡ@�۟Sr$۷`�B3?G�����B��<�<��ꘫ�� ��ｽ�
�����?����߿?��O��Lє�h�HB/W���Q+Q�Q��T�uHך�s=fߦ����������m�x�܉����1����!kY�y�
	�j�g�N���*� �H�G'U�ۡ@�H ��#��?V���������{Ǿ�W�~��ᙴx:���ᯨP-���|����4`����W�}>n۪�nDd��Ί\f}/�ʎ�Boa�1W�t|A9�4��E���	�3��4�@@��EwM�	�^=����wL��g���(��^#��::p��F.�P�7�W��y��-��AmТ�o[�;�o'��_qW��N�#y�xK��	 ���������L�Ut��w�)V��İ�6�{����]ཧYi��6�Bpg}�C듟���B���%{�x�4S��0]�5�߮�-����O�|��� `#p|&�֍���bX���qL-��Ȃ�n��{6�F���ѧ��S%�5��^��۶�CCB:��m��ʑ���-���XEcw\���I���� G\�4�Ds��.)�i3]09i��
3k��f��X����*�M�5-1�Sۘ��ANΊ��X��9�ջ:ky[a�QaK-ΰ0j=Un�F�fv%<�������4�lk��>�336i�
��	5v�`�e5 Mf�Lr�gVhg���K�����N�S�D�۟Pm���vT4�̪b����GP�)�С��r�x��E�H �����An���}�	}Á����'���k���![Y�}�>=�h�D�f��W{����߯��P��$|Z��x6�Qn$Knw*�83���N!zv�fW��m����<�Iou
�4>nD�ۑ���g_q�N�Ր0��B�ۑ\�yL6I�̪b�����r�}6&��"Ov�6���9�I�����7H-��nX�{�d�u��r&�ؼ��p��͘.�σ���S@��$6�|t4O^i}�߾�f���#J汤��fɬ�w���r2ہPLԑB"GʡA�zk�>n��H[�]�}�O��_#kj8K�����o>����~���A�"|����$%|RS@���t�5��EEf^X�1)=�-M�gt�K�k�<5���vA��9SPY&��z�������K�B���'=�7�0�x�G ��'�˺�=z�����bU1w�t|A ���V�^J�݊�V��4v��=���-@	G�S䔃�}�|�M�11�+�-�lɦ�p}�Ov��$%"|B�B�)D���3��W}q�?/����
;�H �R��W�T�M/���	���@�CO��/�'I�Z�D�%2	IMBR$��;,ţ���܌���څ�=�LU��AˏH\�P)D�JP�g�T�z��}�3��Atye]+��D��e��dų9h�J���r�٪S����?q�����%4>JD���[�u��y�&�Y�}���.��-N�|� ���J��H%(�w#�]�r.�}}�{�@���9:��*�F��|'�����w��J{ᦺ�2�o��&�+�j}IH�BQ�IP�՟����+ �1E�p�}��'^��ݝ������8ۚH��f>��;�M�:���=$e\���ʻ�a��\��f{��K�{��k�S�wG��$��P��I�BJFP�qTb���������1ȟN}IH�wk��wٙZf�Y�}���^t��0ʖU������"�g�WP�R���Q>!%>JW������2$Er���y��(ŵ	���?(�ߤH))�A	H���ϟw�t�F���ܸ���k�P�W��)��h��G[X�k�5Ҳ�36�UW	�{��C���f�	%3⒡^�Y	����R�F���^���=����k��3F��j�s�qU�� E_�_F��ׁ)���ճ�ޑ/�����̭3m��>�	�� ����l|����זG���$$��FAJ,L����D�F�g�k�z�U�Tp��y@�A��%8BP$���+*f>�Ϥu��'|A�$��}>)*악}���U*uq�t|A�'� 3�`��������"�}m�]������;���㑦�Yr �5��4�ժ/�
*.��&k_����~��`����V���t|%8�K(�	 ��IIMЛsbCr$}�[��_ӛM��>�H>*�hG�RV'�%C>��T,�����oP��<n�e��J�M2���k��ۇb�:"LŒ��+NsJ5�g���q������b|�zJQ>���y:�_]�Z�T�'��ۭ%aߦ����Y.D��MR� ��H ���}��ת���1��O��ШŊ����R�ӫ����Uǥ�%>�ם�yU�G���#�׫��H �"JJ}A)7�6`��|�֞Vl]�o�� ���@�H���	*R��=�a��n�8���O������u/��Z���'�-��"/���w�F���|{�@��"|BQ��)$S;�þ�wH�\����4��sq�j���X�U�2��B@���$��	'�BB����[n�[V�ߍ��km��[o󶶭m�kj���m��O��$��$$I?�$$I=$��m�mmZ�}[kj��򶶭m�kj����[V�ߞ�ڵ��V� IIO�$$I2HH���e5��P��`�=� ?�s2}p ���                   :       (         � ����I( �
)% �@PP�(JD� �@� ��(( R�$ }��I@T�)"�JQPP$��U)RPA@
)T��R��J��R��I(�"�"�
 �>    aEU$*�$U  <� r�E�2��݀�蠧�=R�!�
���EZR7� ܠE�@1��w`
$�@�  ������I͠<r� P
݃�k ��=��  ]�R��
���`�� ��� ���P�Q� �Q*�P%%B��� ���g�Ԡ2А^����J�=uK��9�����U��s�Kw:z5^mB� (� 1���RW��nP+�z�"����XZ%����T2 iIU�QZ�*�6�U]��Rwc��* H�� ��
���$����_e�nZ�M���JT��zhּ�]�Tp򒛪P�l/f�]��)T���*��J��RR�R���=�/H	�w�W�{�������y�J�΁,A����s�iT��w��+��T��J�B�-T�Ӌ�U{�Ǫ����
 *�$P�|  q� ��R�U	I! %�HTͩ
�fe)U8��4��[����[���P���(�k���[��x�O�*�I냩Hn�O`  �T��  MW�wQQͪU
q�%[�2jR�9�UW&�@�c��֩��Es��ݺ�)F�t�In�*��:Ԓ��IJ@��   ��T�J��P	(P+�R�Y����wIB�v r\ƅ�)H��ݺ(�.��P����t��^�HU�U#-*E�{�
��+�   �+{��Y�
ܢ�[��g�	
���l��j�.�{�=�U{��*�" rА��4n��~�LiR�@j��4��A� hb'�JT�MM ��A��%P5*Pd ѡ���*L����	���H�3�L�� h������+����A$�$t����?��Z�{÷�$$ IR�g����	/�� ���%��[o��[Z�ߥ[kV�mZ����y�O�O�~��L���ʺ�$��{G\���f��6��d��2�,9�Qێ ��33\�&��᎕^G+6ƅ���i��u�����c��yB[�K	X�`eSPغ������oe��A��Tl�Vj�`�^�]�C"�ںyv#9D�e�33Y���$�m���Y/Jٗ�pff�J�׊�M��'VC�l/UZq�!q���1mM�Z-��ȚMhۆ�aN(nUW{�e�9��㷱ь��I7�=����m�6��[��ܵ�U'�b�e��e�a<oj]-���NӼ�C%��[��]*r��F����V'��fR�R�l���9l�o[�̚�BTGj�Ee\�ua������of���m��V�_7���aUe;۹h*ۖʖ*��{�m:+,�D�/����b\(�ͨև���a*��m�D��H�-U۪i�=8���ڥ�YDgͬ�0�(:f��*Gz�{�����b��x� �GJ�JM���چ�N�[��<�����_Hm�Rٺ�[�ΕWj��yy��w'h/u3���a7U���.�z�aT��:73v@�[�r�؎�������dU$���ձy�G4DLR�!ij��ŭ#�MSV��/o�p7�ՖVm_�#�)R߲�X6���"�"k�q��*��L˄*�_k��k^�l��M�.�]�7��ɩ�e�rH������xEbZ���خV��-K*���\�r����Bc��D���U(��SQj@`��ݬ��5�X�Zȍ1����+mX�5�T��mV,[{U����W����Ul^<��u�Ϭj��6�TMC���;Q]؁1,C^�ͭ8�i6�īj�'GV�I0v�U��`j��t��+\�msMVcrf^չb���J��;���e�5eem����X�c/kqV�Ah�)���S&�������o�4ٺY��%r�3M���-eCF���L�*�d�L�JCwq:{[-`�5
ݬ�}+wU+@��W"z[F������6�i�u��6�
gT��xZˁ�J.���z*�#R�X^AUX�*��N�^���[O}q�x�2c+w2+aK+��N�h�Hv�i�[�m��۔�������+�v���r��(2��n̄�3��T�G^��fE�e;�Xc�L�:8�j�lиF9�Ә�-�����˵)�Yh��:QB��/�WM勱��D��J�㡑�ʊ�ʃr�%�VM9LUd3݁m��b���f����5ZrK�YGmɢ��U�V�L��ip^��Z
8�@���y(�*C#��zm:qV)5�^n�M��"�:�y���b
i
jЪ���(�l���'�t��U��[L�:��K��ʣ��[�w�.d�1��x�Z����M���"HF<��j�ʸ���wLXr�re&t��6�@�Uef�&-��i�e3���j�H�^��1b2�6i�&�g�1��#�O�{�N��3B�A(��2���sF+�5,�KCmS�C�B��y��suY4��eK�sF�1�J]����e�Ut~�ܬR�fe�)fA��V��tì�J��B�C�����V6���M���k�s+Nb��*{�˩��I��0���#�yUޫ&ױ����ғ��7�L�>/,��B�G-m��x!�3*j�����u�R�N�=z�{�ɒJ*���)c7P���D��ٺ;ӽt���Y70��d]lu6a졆��e����A-��)��Q�Dn<An`o2��j�ڻ� [�+'FM�P�Vk];Q��:�6�5��f�ݻs*���F�ӳl�9R���J��ߒU��eMIOE��ϒ�+�v�۬L�~Cv��L?P�9��љ(�RR��m���jɒ�D\X�V�\����U�(�����4q�[����O-aǈ��mi&!��.�)
���u����Y/[M�\C�-.�7����j�]�ə�K4\�2'J��יu{�n�Rni`�UU��b��j��T�Ɣ7ww��Qz.d��-b�0�x�9p�������ڬd亯�E�ct^���Q��N�4˷(i�X�ګQ�p[�VV��ZW��ݬu)Vf�NLTrk�u!�����z�d<T&'I]"�VF�˫�H�҂[�=kE�4N!��\;1Z��-��s!����ĥn%�"-�#�㽱aR�����Qc�n�AdFme���\��5�����w���(ea���a�$Y�+H��:�J��[�*�ժi�{{kp�9�/h�#Z�N�c.��՗������0�;��)�[Z��c�)�9��V]X�G6�ICMdѶ���&�Q7Ct�ؕ(aӵ�X�WDb�oq]�ŵL�9����TR[J��[�.(����,c;cID��֙gdE���ޅX�.�/�,;��U�(jȷ]�4Q
�����5��UJ��h9�T\P[H��t)�=R<;��B�nf24f��]ju�(�6j]��hd6�ɘ]X��wj�9��ۏ[ˬ��^M������ͺ��(a�wVj����H�L��߅ �v��k`2��j�n˪!H�P���¼�Ɐn�<pf�bo�i�v�5�d��i��Wb�\{tj'{{F�T�E^M�뙫~�n�ݹ�v���V#e�U��7.�yFSi��`���V��A��%{�mҖ.��.�-�K�GY��r�d��[���ܸ%��&�wsa���ɂ��B�"�i��Y��4�5/U8�bv��C�Dge�Iu7�*�e����S�5B���աpȫF�:�9N�l�o	��N�뱑����eM��t���y+؟p�݄kv��;Z�����&EdǦ�+�,�-Ml��l�S7!ܸq�yF�Ǘe�kk~!V���6�mAg�����8%4�U�Ĭ�w�,WPզ��3"<�d���yz�˭�k�l��I��ֳ.�b�[��:;kN��3�m�j�j	j��*�+�׸(���ݩYYCA�,�״v�U��IJ��Ɠ��5h�7��!/N1T�`Dފ0ݜ�cK�7U]Gf��vV����V�wx(�ܲ�q�(c�Z��0T�-�3G5ŊR��ܦ���є��b�;�ē[�u3Aj�.Zu��J��;n���v�0��U팬ϝ�t�%2d�"�
�(��,R�sv�^-(V�j��5��t�ղ�fo����7���t��U�j�M՗�d���7kS+F��^#d+�O��(Q�wQT��j�[�h�Ovk�W�^�쿲<����{�[[*������f������r̔�eKp;��2�5y��)LԐ�6��w����-���M�M�(SS+���Vb$�J#N3Z�kŴ��T��%k���̽�Y�E��h_m�_bܽ[�N����-�"&��;�pe�w�5��f�Q�y�+	�M��Z��f(��17Ime�
�m���9�Ik���0�6lQ�Nݦ#�h��Z%���0c�i`��n�u��&��n�/5�*��@�j񚴡Uv�ˤ6hƯ7@��ɛ�20��p�r�Q#&P����vɬחL�&�i�O)�ؑ�S��5[���Q�܀�֨62�^IV�yn���n�*����;f�9u��P���3b�����j4sa�K�k//97���uZ�3oKkc�AR��EH��c���^�����ښɨj��L�m̩Wu[tͬ-�/;[~�eo��XݏV��R����T�d�t("�)J��]��
y%k���P2��m!���E��݌˺�(P"�:ڪ�Y��O~�)�,z��Be��������5R�o,@�D�V�m�j�fRA��K��7v�Q�����X�Y�%�2%M����#U��r��H:t�0n;)n�� �q���˵��]���q6ћ�\��h�Դ�ܠ[��l���f��FtԊ<�{)k4Q1�E:�3^#WQZ;wd03�oM
�tŪ���YE�LV�#�B�V���6,f�YB��b�
�٭a�V��6�=�`͂C5�.�=�65���Y�B���Q����:��̥[7l�x��t�l�0ӣqn�Г��v+�%d��D�M���˽'�k'h��,�#utp��J�0]5�4͆�$��^GTp��4L
��5E��NF��i	��[��`�0��f�2�rl�T��զ� ���ub���a������D��V$�Y4me�j����Ib|�ޑ"͸��Qڗ1�gN1UU����o�ʩ��ލ��1�ܼ��r�ĵC[B�ܪ$������f�LAnF]Ղԥ{��&�
�F��NVI���n�m�X�&�5%[x���T�%6�K����r�"�QIh&p�iyb]Y׮��r&0���Kją>��_$)J�L�3в"���L��N��N��w#ә�Y���٘�+�v��^ô��Ŧ�IF��۱3�6<3+,���a���bY6����������z�X������F�"L�ؓv�Q�ׂ���컔�G�謿�0-�ؓ��1��]V�w���h��ʽ2�+Z�˭1���kA���)E1*�h�v-��u��%
m#���d���Q�R67"v���X�P�N�&ٗ&j�hk�������w`�Q�wW�	[	2SyjJTK�x1[7Q�ܔr�r�U��w�޼�$ԭ��V����fe;�����*��`�X�uZ������z~�j�ab��lZ�p�+sF"(Y�T�B���U9�"Va�w� v��Ć����M��;u��0�ԁF�k^n\D�]=�WJ�̚��i����*csS;wE!o,��I��6�fmը��i��),��B2%�[)f�H�Z"��MVq�J���,�i��Y�R?h2��槻�[�t��B�Vs+Z���^i�̚C��8���a+_Q�m|Y�x/��#�C��Z��f�a�f��fG�DZ�Ŵ��؁w�qX�GQ�T�y+v��v^<)a&�����aٕ�mӇfVS32��1m�ɱ2f�NQ"�E��5Ph�ɤ,���V�%f�*0�7{[�$ov�>��i`���Eɚ0��b�CI��NVP-��1kq�beUm�'�z�gPf���ji��y�2�&�Q�T�Л��"���h��9obD��U���5����[n��UcutSF!Z�ˢ�x���ҧz�^b�e����WXl�ә�H��ն]V��e����ּo��v�c�u�<k�R�i�ts jAR��-�-��ˁ�KY�p�n�L��f8Y�_��Uպ��uw�����?�n�Yr^jq��A�ڊ�5��[T5,����h[�2Ƽ���Cv���bӺ�D�j��z����eT��Ph��j0�X���j����z�T/va�.^۸��˨r��:ۈ�[�F�I^At6)Ey[/.�Rl��.����8�F�\�W�`1ز¡3B	n,��e�Xu)R}��{�͹fɹy�۰�*������8T���M�c 7WO+qi��A�o�K�A\��-ֽ^hB�;����R��Z3�FHɫ;�Dj�˴e�B=�n�r^R��Vcc!_nۼQ���&�z~V�%&١�#)�[T�=/Y��la�8�ԎF�[ͺ�l������Kuh�T��;�N��x6���[mL.lVV������MV���Ɍ���#������+f�#/kP��x��Ƀvr��6�0�̶�:T@�Wt�͍�w�[���}���v�x���7w�A:;�eM�A���5dó�`�5�ۚh�6����:��T��-�m��<��D�wgM�[{�5:)�
�e��^��𺧅���R0�ȿ��z��u^ʙ.��[k+'Ղ�55=���ĻM�9x֧��F��#N95��ct�lɔ� st:�p�̍ЙZ��iR�q![�'��h��V��&�Nh��(麺̷���˛Y3e�lW�嬁����eV��s/s>Ǒ=5�.��y��Yx������`���Wimm�]�@�2��4f�:ne�E'J�C�l��굇�^e�<+t]���w.=2�
;v�Mj{۟h��ۊ����
�ec�bt�Y+K��G�L7��Bʘ��DSѶ�[Q�r`��	���Xy�,�+*�w)ØK�	�b�!oo,�Z��͖�@�ǵ���SV!��T�]�ոv�5�4�iҖa��KB��sb�0*7�v�ie�Z��!�V�ڬ��	c���Xj��#.��n�:
f�rV�k�e ����9�%�Z�cd�ܳR��O�
B��{X���ڣ�n\ӹx2�˷3-��-�������p��h�2G٩yN���S���U$��%@�h$�.�֋�Cn��Y��V\��Yn�љ���f�%�uUL�z��n�*ܧb�s�nO��
���W�p���L�4]����/j�i]��Sw���R�@�fn�tUvĨ���N�e��U�Ȓ�̭ԋ�U������L�۱2Y7uB�/u��F4�Pڼ�@��mV��f���-�=I"]BsFn\x�0�ڙU�;��%�ͫ�;����ɴ�Y��X�r���x��%f[�VKxu抿�d�,��jZƍ�y-���Nf�.��'nj���SUL�;��n�c�(ڛyD��+�9�wMRc4�B�	淓2rXߩ�r�n�b;�ƉM�?`WB��'%eE�N1�ڥ����[����Wn\	\1������?k{a¹e�6���[x�4��;Zj�m�wE��7[u��ӵAv4)ˋE��!
�y]H�.(���ӕ���b��y��Խ��p���ov��!�\b:�b���ia(Ǔc,d��q\��%I������:�];�M�d�7-��n��B;n�r��4���"�/�IMdB�e�vr�J��`��ʾM���K{�d��Uւ�{�B�uD��R��M˪������N%2��q���ѪoFҫ7�SՑ��ŋ��nbMT�Y�������2��P�M���r9��O����;1�p�����-hHM��ڋZ��E�����U�-[Fը�j-Am�cm�m���ŭ�Z5�U�Ƶ����*�[F��5Xը�تƪ�*�mlj�[m��[TU�ڍ��*�ElZ�m�6�m�Z�V��Z���Xִ[jŵhՍVƋV�mj6�Q��-�h�j�j6��QE��k�mQV�V�m��ڱj��U���ڶ�U���Q�m�klmh��j�-�X��F��UX�ŵ�mh�V+Z�ձ�ch��X�F��նѭ�5�ckmEd���H		�IQ�}�~����^�������5x;�k�;괅Ҭ���z�[T���1\��g[�	B7 �VR]T!��#��PάR�*͋��3{�	���Wa�Xm����0,�4��q-w��Y"νW`�Uw]D��$.�S���жg�{U����{f�崪ý�p�ǿX�bWU�[���د�>�=^����VE�wCSr�2ٕ;���K��,�[nՕ��}esM��$7�L*�%y����_�fm��6�پ8�
��D�M}����o��;�q�v&M���wd��v�&�h����UÌ�pQj�,�2��͹�0���+)��F�Q���^�����i	�z��jh�.�*�����8��v-o>��W6�EuT�ݛJ훬��orکV(v�š�%��U[�R9~חhQZL�J�����N�mQ�NI嬕���n�u�i_aI�k��˽�Gg\Ɩ�Ǚ0Z99�-�w-=˼����D���������۔"Eֱ�u���� ��X�Ţ�sk �;��8֎[�U&���+o�Vk�0fu���k�̼˗؝�\2���8w�,Wt��V����DM�$F�un�-��X��i��Ǭ�s%<n�{�{��)ވQ��l]�cI������$.5�X�Q��'v���#�t/����e�6c�\������ �]�ɋLj��i�"(�]/+�WR�2���x���n8��t���f����]�+ރ0oGa>ÌU����*��f�� �^C��2b�Z�z�"��E��r v�����w0��h��u��N��!��b�^5��=]�o3D��,���.��%�|r��s]-����tR6������t�\Ż�b���6���r3�:Sx4Y��	d�c���RK����+q�o��R}['E}&֔�^|M�*ﱠ�ѝW�u}1۴�V���w��`���*]�U��{_v�ѵu�Ys�N����g8�R���JBN��M�S�y�s2HE���L�^[�)fs�G���Bu��\��-�`ʞ��R�c1TY�u<���:���D�l�L;�qon+�"��ݼ��}���$*�����s,er���
��bn�v�^�벑��*���{�n�6}M*��Փ�~t�Q�1��/*��Z���3!�cv�]�S�T�sq�.m9P�;$�UjL)�-�A��8����o,·����TZj��e�/&ḛ�74:��g��җ5>�Ef�U���+5����=���J�☾��ݕ�r�fY�n�����0��EG�KM��u��KˮN�e������d4Aa;U6g���i{jU��yN&���e](F^����r�kv���A����A�j��F���)T�ض��ξ���.�a�T�63I�(�� ���O������ev��*�h��!�Ah�y����3���p�y��J�P{z9Y�(V���U��svm���kR˺��'�Z���A�4���^<�y�pB'�Y" �ϑ�2�>�D��JVi:M�7�Y6D�\^r��}��/ض�v�M�beV᪳�UY�w{m���Z�u��ks`�JG���!�����qW��igR��+���ԪTJcn�5B�9�횊o�N|�_q���Xk�ŉ������̽��-��{OLS���ڍJ�R�n?��p-.�%�ΐ˅.���Cc�[���F�Ĥ�.�V黽쭱}t��N��IF�Lj���F�v4�t�o-m�r��;����lf���=���l��m��2��ZD�0dzs�
+�3�y�+�.��nS��!V���V���[eJ�)N*�K���|�Z櫴��渤�9�J�.n5����t7a�	nlV	Җc��;ps�8�I�Y����w������q��ɖ��옞�|�'�s��]Ʒ��#Xհ���7��L����f`/V�L���*�A�g +��P4&�*!ڷ�V���׉\�*���׼�qb*��N����	���+�.r����ˣ��SR��͢�W��Y�l:�����\�����X�Y�I�6�K���*&�`�[u.ᕥ��E��J�4�]nw�mY�������v�2E�f:Wk��n!�U�ǅ�[u����?BJM��T��uL�'�m�ݸ��.��6����Ơ�u���FU��	�3z�,��9b��XN\���pU\{���<��˟=��i�j���h�?=�ݯC5�~�ǃ��N��X�KY7W�\st"Ϛ����\��%c����|�6S��Vf��ۙݹ7�{1'��u�j���L_�b���3�1d�w�A�]f��s�^��o�5{N�X�5$�ⱽ���]ujA�`ӣ�<��/��	1,�9��DU��twz�b?_�ټT��$��v���3�*m��ǔ���JK������*���ګ��Xn����������fc���v�ε�uu�srd}��#��.��.�rC!b^oW�A�Jem�YY��U0��+,�®���^��nٻ����%�l�Έӵ����M�Ü����.������!�gs8,82�1.��Ywչ�A��V��2^
ûN]�f��t-�W�]2;~�hZj]^�k�C�=uW���\
�0mwf5��~�L�����mn�T*���Z�{��=5���sv��A�Ӷ�
��]^m#��%����ѡ�S��jԵkR��_pY�*�Q�R�]��{w���{6]�}���HS��������Op�t����t���M�HnY�N�M^D�&�b��z�k��[�l��gT��{��mS��'�;��8��$<ߌmFC�,n-i�Ѕ��y���#�򷎕����K�����Ge
�1�Fﺫ���*!���B�ЖUR!���a�0f�7s�Y��y��UҾ����=]c4�����ZT�#�V��m�ifowpN�?+�)�-��Ȱ�w�5�껗!_%ϧM���;���Ҧ2ʌ��{�f�GQ.�(wMEJ���cuqv+�x{��ff�fn=S����Y�L��hr]jG���z��&j��Աf�[�3���{(�r�,ý�����Ht�C:,6a�a�ʢ[�{�_�
�N���~���`[VØ��ՊYe�h:�l���u)Z&s�%$;���Z��٣T�̓!Ɇ(v̐i]���'S޺[�ܢm*�Dޘ�U}Q�q�so�_���*�Y�fy\n��zld�Ƽ*�9D��ZOG`'6�Z��n<���ƍ�'Tֳ�����,�GStt�Y�܇`z+vC�m���~��P����m�j�^��Z/n��VU��:n��Y�Y�ٽ66,�J.�g%�{a������U�g;U���.�:C���+ޫm��r���0s7�]VӰ�5s[sf����Z6ѝ�'x�="h³(�qc,]��{E��b�3vͫ�p��xom�B��SN�v������	6�fi����5�r��[��"�A�-�=z2E�1�Yo%����HV`yKv��Qv��u��5��ݾ	�+��N7_mCu3:�ѝ�i�op�d���,o0�k��{V��瘳N��k(+.-c"����8(��	��ܣ\�&��YC7Q�epښ3(gZ����ݥKLS�t����rwۓ/C���ۈ&�	<]ӭ��`�8��j��P�zt-\Qܪ�hHQ�qou��PǷ�w-��%�Y*j�<��1PP�C�ݠķ��'\幇9�$1��޼CNM�٬	*�UA�5���]�ϯ��g�3:����"�mǌ���n�/a�������-��3�gT[��.HL���4�K<��W1ZU��Tmћ�b׷MP�=x!�Y�t�j�z��;��eb�؏u�e1�i�5���[�=���ȧu[g�+b�K�jeQ��r���f�{�5ES�3��C�s06�J���Q�%�/����w�%mk��e��K+mGVFK�w��1Y];�G/3s��%�j��7&��]k�[d��#��_5*��e}�7#5�g8���L�����pٻ�i�^I!˒�܎�������c��U�R�����2��e2�멈�[��q۩��1��G�b5���[�R��Z�%��7��h���~�f���w�w�1AmǑm�k�,��ƋV))���6��Õnݼb�c�t�+���B���	�.�8�mފWt�
����iX��ג[�]��wd�Wdr��Kt6�ݤ�˦t0�[f�S�kf��Ӫ�Ke��C�e�)r�*>���.��n��.�S��ۥ4��9��ژ%����V�m�ʂ���%p�!u|xYe�3v�^�6��e2s/m��Y��I�&f�tD����X�d_u{
��i�b�۫�M��f)�7�	��k�ͧ��+2Y�`Ռ�;\7��uC&nV�'�������Z�r��9���g.WZc��b�q=�^���f��P����VVZf���4�;컹Y�w3~Z�r�˺��r��E�]�u��pZ�Ј����{}��2�N���\�s��O;F��^̼����2�GrYGG]�\=ϖ*�׻skl�C�m��/J�JPM�h�U�{�(���p՚�P�W,��>.�x�ܣ&l��O;%XA�v^-v���/����,���w�b_u��iӌ\�}�7(H��r����띜έ��1����{$���;�6��L3�;����/l�wy�[�V�j��ijvֶ�U�F�::)�N�Zw�2�eR��0ne�T�
�or�w�45�mM��Mq,a鷞�uc�ژ��wI�I���%�Mt����o����l�O�&h����m��s2���4���k`���0:���X�Onf7�Q{�Sz�3:�×jQ��t(���W\�P�Ǯ�JeqsC՗3�d6~Ôm���P�T2��[�5}k�<��j������j�ޗw�0�X��J݁$�;���ͻ����]BG�swn�Fq��*`��pL��xm��5�^���庇j��:�-˶U%e�Ep�KQ#1�d%���s��՚�Yo�oZ��x3VQj�]��H���݉.w��uyUI��l�ܼ�c�&��D�[wJ�39��&����r�ɻB�Ty���c�`��R�Q�G5K���qT�b^�۷�V|�wi�˷]&�w��e���W�hV-e���!�/�]�6�j��}��VgZ�ob|R�����M�ޮ�c3&.�(������7��#-&:+j�UU��tG�w��8|��ɦW\|�_�|����ڂ�u�+���ܒ7�jʭ�X1VE]w��Ҧ�o*ֵZ�&0��R'u�#��%ۼ>�8d�.uL��+$��ַƧJ9�&���������e�k�aë���y��׳�&�7Ws<b�d��c�S�۽�W�r�!��s4%���V���X{�KQ�Zo��R�����R_-�gR%gg_MZ�/%ػ�D�÷��//ػ�UÝ:�틉^X�Q��u�#쩍}�hh�͖�ï]��Ɍ�k,�����H�(g3L��v�j�	%١	zE�6�t�m��KU+�n\W��|6�b�sqB�C`yb��n<�O�w�m{~%<~�nx�X��T4o^Wۦc�Yz���z�n-	нP�=HrS2\�.�&�j5�������C���'�Y�qJ�){��s��7PZA�Fƒ(n'���w'Uaɦ���5���*�N[�b��{I��y��j�u։�����C7�lʷ��ak�L���-{*��\��~�։�i�s�u��}L��V����hW6y��C5�R*:�̛�s��A�p����|�Vbj�V3Z՚�%�v��]|��a3��i<r��.k��W�u^��2V���b�9z�Tn�N��Xݍjĺ����/KS�n�T�vG}r��r�	Zwy83Ҍ�8վ�[R�Q�"e�8��:+�X�yPX�˪�y�[�^7�c��U�Z��P�3��ڼN���N�,��UY��8Žt�#�����Z��=�kB��w���t���B�-�z���m�he�{A��u��󖚍ݝ�|ѥ�A٫��䴷1�7l%�N�c9�De�,Ͷ�M�P`�o��r����i�>Xo>�dfU���qb�$e�gt|� �h��+�ҬT�;{�	+�)�+��y�.�ٹv&F�J�O���ΈV6(����l�����|t�M�>Vl#�#.b^ٓ��U�7d�v��L�y4B����WϪm���e[Ϊrt�ʽr>�G��9����Q���{m{]d��ʟ���^f>ᠺ�o�e����2TFl��Hv��5	��c^�Ό�O����Gg�|Z��d�;��^����}ڏD���=qe�ahjڱ/�ͧ�����=s��W�{�B���+����������ھ���$�&�Et�0�e�=ʼ�J����<H� �u. �ъwK��qvl�o��[�i�Ӛ�7���-V��~奐�Xa�x���h�FmS䶄ч��z��2IT�������?9U�n+TM�W�8+��n�Y�rٌ�1]�	�f�����=��\�yf�(�j�~Ti�7غ�����F]Լlec�j7�rF��0�TQ8�w`ևM���`��_v�p�*��i���X�K�S��Ė�Y��d}uW7LX<����:_Q�J}Y���Q��#gV龍=��xwDv�5wv�����!���d��X��^�x�432
��ctfnK�&\j�
�)3f�Œ��͵|��n]���j�OY4wa_A�TY[�gC����6�%��x�`Ɛ�+{�+�Ъ
�_m�4܍��s4��]�eh�[T���ࣗJ�nӕ����Kl��:׍�d���i��̫�lئ��_S��ƾ����ì�����L��n.�!���'S�g�8`eػ�1�\�՗Z�*œ%aqM�8�A�{�.�]$�k�9��m	/*���uĞά?q0���D�u}w�$n�t��t��r��s��#�=�?�	�RBB�	$����j�i���a��l.���y��,/F�`��ܩ7�u�*�7lOT��{�mݥ�4C��d͜�%qϑ�ِG�	ɶ�Z-m1{%q���.�a�1�m.ip��
\YG���`��w�pUt<�V�ι:�ώ���WS��Ʃ#r����ë��uƌ
�4àc`�:䎚��&�Š��6����P�Ò�O[��(W����9�.
�K�v�!�u�W̔t�-�J��5]XWLT��1pon{h�� g��8��1����}���v&ݮD�EC��L�9֩�j8�\g`��up�twC�m�κ8���s��̧aWEH6�Y5�{���`�˭�N�m�7\k����m�m^�{XLJ5���JWk��fb�<���๮9���X%��ɥ���u`2�e�6�mtĄ�β��"��Y��h �3W��=�b@�=�<;,C
�v��s.\Ѻ����c
We��B�Ն�.�muu���^��������Z>8�v�i�瞛
�[wbq��@��ľ����չ�k;���YZf͡�`6DGWB.mV��-�uq��y��R�5n)�`��rX�R8F\mH����2�R�t�0�4in���eb834�ײ#�{mї�*񨲯*i</�Οd�d^О��S
��yZ#�c���7)�f
KM،ر�(�n�pS\�]\p�dPv������c��JjU�I�vUv��эҎ�8b^[�l]vҤ�:�6�U�ٕ	��:��P�t4dƖ	�u�-ѵJM��-��U�͍���"���v5��rf�Z�.�Lhu���sb�ru/:��O�6Q��Zhƣ+�Q�5Ͱ#&�j'`��݉:�C��q�j�՜ڞ��u�l=4�Fɛ�y�i�R���P��g�3�p��U�禳�,�[+	��jhS]U����q�^��Ẃ7[f�h8҅�Ƽ�bY]Z.y�X�h�kL���Z�R�mkF�J.�c0�3n��B��h�I�e�{A���@J8��Ki���jD�-6{�Zm��h��n��Q�k!.	rV�,c`�͐�����=a�,�����6�m�ezx3\>���;:�N�|���j�k��ʹޙ��8)���s�{��q��m2V�cw�9U�R��T��KP
���H��Z��b멼���à\z���4�`��u��n\o������s�]���3=�_k'� ��N.Ѷ����^��
�q>Ձ����yM|}��ﳺ;p�M����n��6��$6��&K��0�9��-L��R$a�J1r6WZ�sC/0���OG&��y�6��H&�n���;j�BbM�4��!mA�b��Q�5��l���]a,����[U�7�*N����|QݽQ���L�a�Z �9m2���h�.R�����;,�� �=.X���gD�\h犃�;��d�mq���'�Ly��w��X��H�F&
�k,,�n:��KwOb;.�]j��i%:�z�����)�h�qh�f]4ͽRzŬbLWFY���||B�Ls�1½<��i��pf49�HMf�2�T.0�v{)Ɠ�G�O8����wY[s��{B��S�t�P89���z�5ِ�ܺ]��;3�\�
������ƀYe#���гP�i�-۰�����l�n���ž����zf����O�W^:��=A�[:�w@�9����c��M�3K1s��ibU�1%��v/Bv�����Kn��͂���2ݝ�f��8i�:ͮ�9,�6JM@�a�l7$�\��7m�b�L5�l<4��������G
[�.�6z�ih����Sz��������t��L�fέ�	qq�!���7cq��q��\4��x��)f��Qs0MD����ܷg�5ڱ�l����	�ŘQe�fS�ؚʹł��mU��cuzq�G=:�u��{@���&�6����,��P!7`؈-��Y2ֳ�Ѷ����,�q�颅�7n8����muH�Bme#e�Q"#.!�t4n�%m��'q�8v�4=��=��͢���&�{l��:No���-�7���nA���ϔ��u�/��1��W�����Mvfۅ�(����7u�:�Tj��n�V��nE��Q+06�Wb�k�]g�8�ܓJz�vx����ܦZ�A�����v�T�i�1�	;��v|�F;<,�i7R[���J�ݣ,�km�B-�؉ց�:#e�żQ��8�r�@�.�m�6ʖ�%`%&bi�P��앁\=�']���g��//���z@�d����X!n����M��	p\�M�Z��ɥ�-��}w��Ӄ=
�����5t�k�ܦ��-U��ն5�
�G��E���}���#&��susk��=J�D;a�plp���Ksv�;K�*¦�f	b2�c1��^�)v�gq��S6�ޮ��{6�&����N���2��{pg.�勄]��t�����̐ƺ;��w.��t��n��m.�o]���M�n��ڶ�[� �Mn�O8�ZՅb7\'�^M��X4n�����z��m���n=�����&J���ۭ�n���)��ma-�a��Ji&�=��<'�!���x�����K0��&8F;=�i 8Ƭv����`X�P����FX�^�;d�{3�cJ���TR8��b�9c�S�3�[rOTBָ��,հ[�kie �r�ߟ`:�`}���l�v�{r�ut��6ĥ����kC�:�ق�Hz7���>B�+� `YCP�M���GX���n9ʬv^����z���N�U�����Ʃsy���ՋxZ�&��!ahH[���Wns��dC���r@��aFں�:�#B���s��v�mq�؞�%M�n�͸v\Zِ#��BFPe�Z�fl�[,��Fe.�G��C!.3�rA�{][�]l¦��`�[�A���W1���3ZF���Bҵ�.�����c�O��H-=�Y�{#�K���:�n�����9a��n#b�e&5�Ƒ��q�t^��p��Tvձ���l�"rA6�j0\�w\��݆U����'Np�t��+�u��
8�'c!� G#��u�=���+�M3�28�	�J��<mFe�2�[��בs�S�r�7m�M�G���ɴ[O�����V��s��ֺ�3ڥ��A�����w��>rn�s�E���0ƴ�r��&�XL]�׌oGA�{tvͯd+��7��e�"U����0F�s؅܏=�]��e��$��K�HbYaWmuvc4�c%!X�h�[�I7XF+�u0����[�l���Du�X�ڒ�5�fÉC�:�QZ��s���m��?u�,j��>q��9�9w���4Z�IٖRA��p�L��M��ۀ�u�Y;[$��t7.�F���fp�k���77{���"T,I�r�l�f5�̼�v%��<��`v���ѱ�����GLK�4�Q��=��ɇ��޹���Ѻ�9�\\���3at(��a��6)nѣH����.4�����fY׍�bW;W��1KVV�H�l�@�����E�g.ҹ�8�X���������n�3��e|n�\ �+�X�h�n-��(ZJZن9��V.��A����M^�6&�0�۷���ܢx<�[`.ձ��������5ļ@۫I�F�m�����[�$ S��l�ڂ5�1v�3�ڗ�4xꡳ,�k4�{a�K��ƣi��>~�����ڀ*{�w6#�^YA�;��]ct�lMh�D5��k���k)c1-\�m�V𘵸�픻7�̼�-�]��x3������s���u��L�m�[u({	�M�'D���m�k��3��8y���ldHa9%�&�S�bb�[ 6*c��k�.9����'lf��:��K�����|vu����),	�֛���4�h\L$x)գ���bV0�ʑki����@K	�`5��5TR�(�6�{T�h�ƶ1,�#CF���Z�l	�݄x'��<�;��]�.r��H�c�cK��Q��/]�����*E*��S6D��2�6�X�<�Y������ƻh"���͉�hW&�)����.��:'�ۃ�m��F�s1u��!�X�[O[l6-�n5�Ma��݃�E	�88s�������e1���|\q�O����ie��G�m�3K�	�F	�m�M��A��݆y�g�c�,���*��h���*�Ƴx��N��ȫ��[��ޞ��kB1�qp�#�`ׁ�Òh�X&�Z�B�m����LD���d�Y��7S�kEVzK�wo��ZnâwWV���񻈰\�s�,Lϔ7Fӻn:X�Bi�I��G6�sc���{Xn��͝�����"鹡�u�[UE�l�ˮ6F�
Lh#����F�X��հk���SI{6L�s�pe�vz���{SXТ(�9�7Wh�rDl�{G퍤�.tj�n7�^�,����u[�x���HM��5���`(	�l�rk��� �h�X�"G��{j[�t��rΣs���	���c)m`C=�Ssa�d6�=n[������b�su��BC��
��Asm���L
��Q+�&�ڋ�n�刜u�Þ9�f�v7nh���k�;m����}i��Oi����ӺM��H�wR��+r��vѶ6#�p��2&�DST�ZIu;'�y����m�\����w!��l7��wf�3�瞃��d�sۥ�
�U�����*e����'�]#�3X�`�5#k\�f�����x��鵗�rK���#��\�n9\���U]t�tr��\\�Nڗ�y���-u�@�KiAa��Z��kARb];�R:�]p'Dj��X�������sۨخ��\����+�k@u�s��36��U�v���u�r�T�uULUU]U֮�����H��dFP�D@h�ؤH�cgv��hѐ��AT�F ��2RD%%�b��$��I�����N�&#��b�E6#��1��X�d�(K&c)7wR�3&4�6H��a4�ٔQD��)`ѓ�I1�.��ب�Ɲې��3`0ll�4h���I��f��Fň���Td&�Lh��cF�4[3"�*(̰D�F�-��5�nT�6(�EEF������5�� ",`�-��cBmbM��#����$T��E#ݴQ��%�F�HRm!���UWǯ�ǝ'J�le�6�u��{p0�F�5dnx<lF6(��޽��Gk�]qc	�x�g��AJX�A�.�����[�wzs6
�P�l�$\u��s�Ws����b.pe3�bhZ�f�Nm u��qH`�/VM�B���J(�ku,���݊0Ҵ쮔+ �a��]Z{���ݷ3ۉ"�u�@��4m�ۤ���n�ۡ5{\p$����Z��ո8&%���ɹDۑ�ui:��=Vy.z�pI(�@����n�]���)�sf�4���f2���-����f{JgP�704A2)���ttX�Dx��[P�F-�k��Ї=�=���6������q�/�hܛ��s������[u
aa�k*�������\����<�z��0��0#-oa�Ս�^�j+�<Gld�̜���^V.�s*�`��W�����L��C���V�'�zt�#��0��b^���@eЌ�]���ь�E+�7[��b�y6�z�J�l��Y�n����vY���n=�s�8d9<E	p�iy!^�ܞ�h�5�I�esnYp��r�n�Ci��e��f,�A���q�	�P"��6{��Tt��
���;}�c	p,��Ž8흸���{E��u�M(����Â�M�\����PnG:���=�l�.1�z�

��&`��8�tv;[P`7-�G��nJbpS�6����hMt��zI;i^�5��i�e��1� B��1V8IY�,�u�j鬃���P�͗ƪN�:�sxy.%z��k�.{u�b�Ýs�\�卐a�K�֬�]�0K��Y�FK�e.t��=�F!m���"�%�F�ai�SF�ʹЃg�{t���a�����v�cn�;g�H�-�%s�Y�"f�ݤE�iA�7�;k�A���iY�%�ͣ�-õ�e�{CE��7=�4�s��顶�gI$��U�NF�)Km��l:��,�T�հiQXF=hE���,-d#X6YAR�60�W�T��Rym hֱX@-�:�RF��mb�x�*X�`��xeX�	h� 6��Z�RT����<4`[ YJ%�e,a`�-�^�x�XR6�X�-	j6�YB������	������W�sZ�4r���2�&*	�s6h�֌c��n���J���C�H���?���L�ԧ:jy��>؅"7x1~�u߯���A�a����D� D��	�&�p������o�;��_j��4�Y�z�S�\?�LrF��&�-���� z�2;��	ޠ�F�&D��ͫ�
]��o�ko;T�U	��Dѳ�v�w�_$`?���d�FY#��EdZ�����J_~2D�jN�K���w�!�#wx0A�A�+��6�M��f�`D����d��A�D��}^��Q^����P�{s��M�z������m��)|?�%��� `�
��E:�#aϭ���ݶ��,۪:�i�֛�s�w7<�/�G%?�oF�H� �@�f�u{܊&�{D��sn�7&R[�_^P���d�0d�&H��y�	�sϩmr�s�I�ml9$��݇�j	��Ju���uŦ�
}������Q�]U���7~�v�[w"[�%!g�ǽ�P�z�c�3���'��iv�y׷����;( A�"�^r�$S>U�4W�DO[`��/��D���3���5HV��Zx�.�=���%E8"��q����FH�J@�d��$B篷7��؝�Z�-�a�rD�"J��哺Q��fꥃrs�������`��N���o�Ә`�@I�D��d�}�_�ڰ��ӉM鴹j��ɬy��q�� �?��0D�.��s�nfrW�}Z{�#Cm�a�P��6��j�ed2�.���QYy&)F���0Ke�V`{ɂ�A$a�d�?�����Ʈ��������}������Y�w]�A�ٯ�����&�?��As�P�30C~�f�'� ��/yL�`��fj��rs����"$�U�,��{-/�v��R���"�"ĝs�)vne�5� ��X�b��$p��3T��MU銷���oi�������G�������R�0l>&	�u��o_���ՙ$�~>����J� �2D� H��[���{t��O��A���f�vs��~����E��q��?�xo�y�i!�� ��0� ̔ ��c=��޻����q�اw�x!2L�K��	ۉ�w�@�"����Dz��rE�u
�i@(�4�	��t\��8�Rf�b�:�lb54���-s��e2]�/Ӽ��ﷰ�)A�)-[�M������S�=y���f�*����`�rd$A|�0 � �{�V{�J>��~#݌?���`�wg�~w5��W�\t��(�S<��j݂z�2:F��Π�2F�&A�D+B�=*��oU�ޞ��1��)=s;q0A�	%���F�J@�{���J�▯�I�0vR �"�s�Wj���bЛ<(9�s,��>X����:��b�ܛ�^��ݪ11��Oߎu�"�In?žv&��H��,�����n�Z7�fK��`]��e�Vʋ�5}�DIfH��@�%v_���/�3�A���+_<n�[T^nW��=�_?�F2R �$S��|��:���}|}�I�E*��Z�0s3��Cb�/'<�]�4i��Oʘ-� ��A��`� Ⱦy{]:J��3],����Q�T��XA�#��������� � ��V%^��|��N�"	�����ku���K������� ��0��&��E+�3_ː@��lw�|�A$_?��LR������oO�ō��M���{ڙ��%}fH�G��^깇����>�����@��~��:uAj̙���vs���т���ۜ�C����Ό1�$L�$�?���c�w#�P �4��u���K������("��H� ��y�z��/��W�����_�C�v�{ۺ%���r����QUc"�}.@����x�;Ҍ8��
�������Z�i��n
�[[��Zy�����E��*�;�ȗ`r8�(�qJM1/CAE�/���ۃ�d����ټ4f'8+$�=��/[z"C�msq��w�+q�3�]L�����0�%a� �\�$�1��u��\�̀�W[c�:8N�S�n��؇���U�z�[;u�Z�)��z����=�7P;��}�(�sÜI�nR(����TÎ��l�w�L��vt-0p�j;�]��߿���n�VY7���{D�P�N�n٫]��
q���B�.H�*������8���Ry�J��w�n,4=�����m�VZ����0� �DȒ0���!s��z����(,����"z��{�v���햜s�n?}�0���%��G�J�;�?�"H���H�$F-��WyH�eͺZ�t�X-	��P'� l�3$LG� �"H��<�^/_- � �����I��g_b��^�(^�_x\t�AH.����`���:���tL$��IfH��t�
~Iu���N��Yٛ�Z7g	ۉ�A�I���==�~�L~�g�W���J8]����mѦm&+˨�i�kF1�ƘD&�T�2��+H?�L�w0���FH�����犧M��������o+�P�u�sbd@I-��2D��V%e�v�Ƃ�YlU��R摧��Ua[�k2'��"�z@.���o%��NŷY_qE�n#�t��̌�K�C����#:0�gw2���m�xh{3h�w��F���޿j[tho��/�� �;( AF2E��=�����v*���&��^��KF��	ۉ�GDE�F��?I~u��e۞km|�da�vR �"bN�^w�:�6G��������U�Ϗv��O�A�A$a�$Ld@I^�^��<v}o����4�v̯^�ow����d�G����d�L��T��iM#U,�MNV�AP�����]�ap�GY녦�<��)ݳ��+�	i��2���;�� �"w�{��[:JN	;+��'��|���1��!��&�̢�d)y�4����gY�W� �_#���}۝o%_l��6���@��� ����<]�Rݨ;�!k���2r%�0�"H�����Q\�o�����Գ|]��BD���t�YƊQ��ć�[$d��-�8˽��sfbp,\�5u���a�J��<�V�ş]��f��U<�S7�Ud��=�L��?���"`�#`U���9�۷�6�9h0vE�D=��{;{�/f�kFlC���D?�ͪ�6���bc�9�BH�J_~2D�E����e�L�
��O賦M���7$y��P����rP@�6G��}�D/������h�4�T�
{��֎2�����M
��BLY�p����)5�
�Wc�rz �I�I`��y��ڦ�^�[�x��˓�צkG�$4�޻��#�� �"�I�%D�m,�������`��d��nޝ�[�t��6s�ӨY!�����br�=��� ��LD��d��H��]�ݢ�_���nM�H���P��8�� �fH�@�#���\�t~swmv��[5h#v���ѿ��?�$�/;+N^��4�ep�L����Ѵ����s�&w�lfnk�����_5�yC�|X��wL1��#-�oof�;��٣��/��#o}�ή6׏/aݟ:�Y1��������	���D��A��I�Dv�{�1s��.Lr�d�����֍���v�`�r$`?��b����kM>~����Ym�Bi�[� �1�I��]k�\���S�1�uStJ�A�Ī��KO�;b�%/� ���oo���H�~�P��6Y=�:v=\ϼ�����A�"`�$@I��2�����r�A|�cM�1u�:�������K.P
b�AΌ?��C�s.��y��L7#`��"H�2D�2 �!(�w��^8u��g`�Ǧ��n�8���dI��"),]Y��R}��6�����3�H�$N.齯���f�z�N�M�	�A,U��#�u���ɢ n�0AyD�d��D�/��V�X��f|�ˌ?�Y;���FL���ep�S#: ���?I��}�ܳHyy]��z���<��wMC����6_���qV({�ϼ��{,�6�*oj�����fz�Y��+Kg���}���-!n,�Q�l�\gY�v��L�����q�+۩Cx먮v���G\��>�sa�Mm��U��!Mu�h�A�=�:�t�u�c�-��흷Ձ���DF!^��9��Vü�f<ήt�'	����l��f�a��E�<;{E;	Pu:�@�5b^�${,m�뫫,�if���3\�b�Ek�����X��q)]��|���N*3*�F�֢�ٻkw�����UJ�eA�d��gA���t ��2D�P^�Fgt�����ލ��0vW��ˈK��$ݯ�;�����#�H�{���c���>�=	=S%�ަ�ݹ�.��+r{���ټ㒂��"�H��*���[b��D9N���,�#I�Au�Պ��is�&0�̮ ���FtA�)A�/��K�x�Ct}�'��_k�L%�޳y��h9����� ��ڮy���I����"`�$a�*uL��y<<��1�`Wt�m__=��Z�Cf�`��#dA�$O�'!{�3�d~��]�Ԩ��EҠ�$U+��I�\��2#, i��v�4���rP%�'Ϗ�)���("$��0�ʝ;���=�c	^�p?T��՞�2{_��s9�w����&0A��!<����]�	ɦ�\���t������ ��UpdE�(�e׻��7T+��I���w
�R��o
!��.N]csk7�쾽և3S�m֏fΘ#B{7Jz3g0~;q2�"Hf�n���36�쉐D����2E׵�e-j+�Ž��ީ�s�'F<��>��3$O��D��UY�jU{�{�@������F����o]��f ��W�{S"�� �::����i���F�J$�?��sզU6���9�o^�wvЗrz3g;q2�"H�#�����iz�N?�]��'��h��nP�eX71f�ѫʶV�����&[~ʭ ��L���% AdLT�ίJg=���.��C���1��}m��3(��� ȂIfH��g����c}��=��bw0x�z�r�����%���Ό0d�l_tmCZ�onX���{c`��H�2D�2! �nx�r�{U�ęw���Q}Y���X�ע���߭��	Ըr�k���\���.���2���˦D�ڤk�;����e��=̄�]^�H���͗�o핳���i��ɮj�"�l5�ohڣx�j]S'm%T\�͌��&�o�lӛ�'��q�kiwE��`[��-];��Z�G`���x�X�+>�O<���!-�d�ͱ����]�L��{�vQ���5Zjc�a��t��v��nҩUo�M��5v��CX�����j�&8iVz/��������i��)lYfm����S硉$�������o�O/!g�O:Ib�昩vh�k�8�<��>��6�]�MgU
��+W����g[��{ˈ��s�Ѹ�i�t�+����RV0��+n�O��{�%�ͼ��[Çm:	@��]x���2�����I}�[VvH��gi��J.qu�c&	I�<�v:ĽUw�g&��W/7H�9ZQz)�H}MSҥGY^®�8.�z�,����y�s��.���on�V���n��Aj+s�T�#�==g,j�D��f�07���O����U��+��.Xs+�Oi�����Yl�S5�OUD䫝Y#KPz�ڵy�g���̇Qw��/=$
�u[��tt�;w�w�]#�b��=��d]*��{|�NJ�j�*�̹q^�ݹ{3�K�*5�ԓd�h%
ꠜ�K��8�H+���f��'EWe��}r�����.fUa:�&��0)�K����i�E@kX���������(��i�IJ1��fDb�ё1)	h����D�'��+F �QF�&�h�2!�Q��0b�ٚMB&4Qb*,A�P�6��&؈ƍF�Q�!�(R�5��ld���݂�&ō&řI�V��fFɢ�50h����b�DR!TZ�r��
�n�,Z�kE�DjH�cX�jHM��KD��Dk��X+mDEE�DQ'�Nʽ��nЗr
z7g0Aۋ�' �G���$a�)|�}�n��ܬ����$��N�;�mL�l��Qt6o �9(#�5����
���� D���2D�D�I8:�C8ۛ#ԥ���
��\��׺ ��_xv�> �F2R �d��(I6������y����� �֚�Y��4Q-���H�Q:��GA���,t��4�:��%��e�~��"dBݺ�}*4=&@V���Z]Cj��ԹiuGH�rG��d$O�*�4{�e�N�p3r���'�N�=�L��y��ٽ�`�rP_$A�"f����`[�6D!�6	�'�	_$o��������n_��v�/.�X�J�n�O�S#: ̔��$M33((q1.s�i��81����ʤ$AJ�ܭ�ǡg�&��n�`�v�`�Wz#��2�6��Ӯ�m
�߲�듈�	��nj���@��
�-�<��H+T{7��u��� ��WL�,r�A�g�[�c�y����Na�(	"��"H�����B��^���fn6�e���@��"F2GD#�q��-ɛ��)T�+���-�)�$�@&���V��*HX	�M.�m%ҫ5W��|��&�:'���$��$Ct��^Sk� ��^!���xrn5��d�W��� ��}$��J�;�~��U��4��|��7+v�\ꐳ�&�Z3g0~;q0A��"H<�����}Y�W�#ͥ��6&AG��`�$Z�/b��+�ˊ��3�d���x0A͠�#da�$L�$��L��VY�H T3� �3�9}bH�9��8_�n&�J�%q��S�����Q���ua�lL$����"H�H�i{2�n��ٳ���ղ�N��Y��h��n&Gu$��F�J���7�t��0��L�l��CLk�Y�3x���z������:��B���w1i.w\��d��{��~�B�Q�W���!x���gm�U�'��/����u���a Ǹ;����\{��=���9%�e64�6BX'm�kM��d�&��������
�����x�XC/h���Ы�&l.�;	)Z�Ҙ���^^�b�T��ay��Ӊ�㬋��s뛜������%��MJ������ �%��jÒU&4,�-��2U�+m"��-e��&�M�}���_6^��Y��#l���&Q���b�u��Tq�B�m�*�A޴�鱆d���&*Iܖ�mλ�<l:7��`�K�}��k��7��7���("$�0~2D��Es�wݡ����3��gvN睊�IB�d�z�0#:0�����_�V�g�&G_0� �P@�$IdB�#�V�C��-�]�ީ �Z/g �;|�}�	%������Q�Y-�鷋U�2�}:�	�&M�Դ{n{�LfǨl�`��w[ɕ��4����I��"`�("$�c�i^6�_ �=�ɓ'��IB��+��ש��fJ�"��WRz�;��V���7m�"�)��^�5�+�avf2�#�F�	"� [>$�����E��(^j�5��o�zH0V�l��:4������������|��*��DȮ��g�أ~�k�Yvmu�u�䕓��d���ڢe���)F`���s=�3q�So0zLw�+�hV����ړj�vfN�aWu.���%���w���$ ������S���1���P��� ��"�y�=�]jA/���ɂ��"H�rFz���{�[٢��aOd"��+�?�L�3�)���$`0��h�*�������-zD�"J�{t�.��d���zN`��O���/q��0x/#��J�|d�����d����^`�S,��>v�c�O)��W{��U�btc���l�3$L%��g���7%z�vK��iB�s0�{��G���lk�\���xcu��j�LS���0A��� ���/���������󰧽�fJ�<��~���LV#w�)A�&D�����A|�����],Gۘ7�X�y��9/5��ػ��=�V
����\3�DI���N��-HN�<�){{+3$�Rm�KKSP�6�n�M�s���ת�~O�R��s.h5{m���{L�M�YR;��k#�t��\�B�Y���m���^�&�ó�"��ʫ��ʙYϗ�A�A=�����7���Ε���bFnH~�Cb"!�K؆�6f�LCk�(h��E1�l>h݊b؆�ݐ���!��>e�q��9�n�h�����!��LCh)8b/} }�lCp0��G�Cg��������#��g��-�̉kɥCb>�H��(bGrkxz돇��LCb�az%�MC��{6@�!��wd-��6""nı��C�wh����҆�ݔo#��ϲ<X#�h�}�{s^���;���>@_6C�i�|�B��<�Hг2@��6�(��9��/o��_|@���X��HI����"�I�X��%���DkR�P�:�RT��:��D�c�܂��5��!г!	K̔.�f�O>�r���t��� f䇚�̷�G}0�B��HEwe	Rh̄����"-�������o�X�Ыr@��6���ם�����"��g��n/}r
���HE2 ��0�/�E�+�J �vC�BAy ��3)�`�2PR`��J x*��T��������{.���쇆�6�e
���Hг2@��0���CB9tg�ldM���E�AbhF�����%4!�̔.�f��>�r���t��� f䇆�44p
Z��9�_l�/�y�oR�0���=+Ə���~o�Qm=�QJ�{��0��7�8aK��Zo�!u�oM��]c5���p�|����?�����/��#@fd�i����Mfd�%�fd���|s���TT��ځFd�1}����w��{����>�����07�T4!�ܤ"�d-c̔/_s���ן8���X�:Z]�0��]��Z�����u�w		�(���U6�k@=S!�hC�)��(E0Y�()�Fd O;��ڬ߽�g~��9�������n��G���rD�hY��)4!�32P�2SB3% w>,ڽ����j�hYp�i�ߥGg3�����W���#�^ ��1%܄"��@�(>�����3 4_d(hC`e�PІ�������a���_;W����ۇ����ͻ�{���V� ������hC`o� ��ܤ"�B̀%��fJ ���"e�_Q��<AU ��{)��o�((`�љ w��s�n׼K�ל�>@}�!�`_6P�����mn����pM
����m�(h�	��My�HE2 �빓��Q\@�jP�{�履V����W�3rC�B�s �B�RC����i�2 9�o�޷����3K��"�n���nc��Z=���'qz��W��]�&Eҙ�6z7��m�]�Zr�s�̩��k94�|}��x��r���I03k�$��ix#�P�D��#��XN�[X�˰6�M
��/*m�6���C�k��/IG${�n^.����hj�`-�*�x�W��v��6b�G!q�A��jE B0a�f�̍�X��d�0lu���@��ќCY�� ���9�79�4myʈ��*W�f����-�X�I1R�2.�������b��V]��i�����b�E�E6�vV[*5�C�
;M-�]�0+[��&.��t����C����hC7$ г2@��a�����ss}�����O��O�@]�y�2s3�9�#�G|hs$�Ї���� phCL32P0̔
��#B;<��>�{���U}=��~젤��2 '��e���^�=��9� >ݐ�hCL�Ȁ�� �fHwm�뮽&І�vvP�\ R�y �hCY�HE2 ��4�$_ (L̥oL��7��V'1�yiM��۪��Hy�h9��$��B)0Y�((hd H4fHRhEFnw/���{�W'�y�B�����{�BT�3%�߷7��ܭ���\���.�<����
��G+3���'y�\�}:�u�r�	h�J������)��(EfJ��3�]��|;��@��E����ⲽ��V�>ݔ߲P�І�d-3%	QH� M˰C¿/߽��C�%�N�"�k/F��q�;	x�\�t��|f�lt�u�X�D�V�#�4!��� ���B)4,�Z�̔vs=ٜ�{�>�{��W�7nP(�\��Y���_b��B ��B)0^̔�3 Z3$(hC�(T���ˏ9���E�T�R�=�����R�."3y=5Rh��ׄ�%$l�D8!3v<x�fX7v�����:���������u�G����D�ME��A���4/n�І�~��@W�w{���_z������ .�<4!��$4#���SB̀/�a����z�(&yr4!��@�2��,̔%M�s��П�ea�U~*d/M_��k%��| ��@�0/�(T4!������i�fJ�2Z=�+ӽ���}� ���B(�-l32P��rg�r+��먊�ې�4!�Ay���'7ӈF���zPP�4f@�fHSBY�"�$-3$	�{q��	�%��_}^�k�}�W�ȷ?yw愷�TЇ��B(hY��!���@W��3�z�������A�Ѱ`��y:F��K�f])�h�	cUCl�:��̐�hC�y �My�HE0Y�((`�4f@���e�ۻ^��N_)ǐݔ��n{L�zN����[B���������� �hG.�c}�����hW�Z�_�(����r+��먊�ې�B�^@)hCW�H3%w�K�&��H�ɀ	M��
hCy"��@� q��$_ ={an/�X���]~�/ӎ�z	���8*��Cn�z���o�D���Ǣ30�a\�YI'B�!�\�7�G*3�_.�a�]A�r��$$���og��s{�չȷ~@v�?4!��$Bw)��� K@�2P�32B����Ɲ�L 
7v��`��(J�3 N��2��ݯD�s/���n� ��(^M��}��Aз�(hCaw����̀���2ASB���RhY��n��c
=��#�/ݔ�|�}���>���u^ ݹI^@)hC/r��`�2PP��2�E��Uⴾo1W���T��i�������]v�Q�q���^��k8-�c�r�]5�ٔɁ��P4!�-3$
hCfd�+�{;�^�9��}�|������y���;[���~�*�A|4#�r�SB݀%4!�̔��hC�2KB'���+�j �ܠ��/d On�2/����5�����hCL��4!��"ZfHE��ϡ��!0�d�)�/`$hKג
��<̤"�d-��@=����.�2�<���ˇs��gA� ���-e�)�����ƀ��
��>�x}��+��s*P�4!��@� q4!�/2P}�f�����~����� 9phK~�M��3�� �������W8糏24�>��i��K�3��ջu��ń���I4�tlm+n�[ҩ�P��E3��O�����b��A��w�����Bw��@_�	~a�������Rh3 ���B(`�2P?��e�M|u{ ww��^�վs�s3���n�y�+��&�f�"F���i�fJ�L��y�Uنy�rk9�9�s��
� J�<����ͷ����\��������Ȅ
���M}ͤ"�B̀%��fJ����՟y���l���v�<4#���\QOӿ;A_@.�!��"�
�҄��2 $h̔
��(TЍ̿��w#����4�A4,��4!�=�J��wb���{���;���0`o� �hC�m!4,�fs���I��"Xz�P�9�HP1%�@)hC��B)��E���P W�����-EW׎~+���!ǐݐ�І0/{(T4!��"SB����6�(
C@f@JhG>���]?t
ߤ&�0��B(hY��32P��6�g�}篞������xhC�-��&>�*k���
�@��0Ch̄��hCL̑� �3$
�~7���P�0�jP��碷��{���m�������
���B(hY���9� �Z4���\�Z�$5�%�ݗM���ʫ[dn�&Jԇf	
W������޷}�����CV��gӰ�{���d���4>.5��}4�\-�	�E���r��ma�w�{����O�4�4�ߊ5��}�oo>x�ތһ���uEVK��nV*�N��%+[�1!���f��G)`k�����e뱰��
w�r��]��IYuY��Hn�ԷYA]�K�K���ڄ����M�KJ�{egv(q��6�+s�Ɔ)�b<����Q�wB����5e⿺�P<���o/�5�N���u���
���{MH���ǯAhV������<;U���U���w3��2g��j-��嶣#<lR���7�$�s�1N�g7�j��_;�*�Q�GGhBhdm@��e�yݖ�QD�w�LR?;|<�o����Mң++n�N�;��5M&����F�X���ر�o`2����e]�����*������FƳk4�$M����PRAd�ư�'^-.<�b��o�����Qj�d����7I�eZ�F���=.ÕH��ʥgi�9P�Hb#�Yfcs%�]m
��R��A��	=��[�UT���sfo%�W9Dk��i%�a}F+�UF�nwKʸj�فR�V닐�V!�PUټәA��F�#���%��f�;d1��bʻ�{�M���
p㷼w�^���,��ǲ�ܱ=�V9�&m���j�ΤONJ���nﲟ������L�TU�PB�I�u]��w�rnf�F��,�г��=-%�:�8�gE��Kg��?]��/4&�6�4�j"�QI�	���i"��,EA�+�F�`�J�6���тŊ�E�J���,k	��T��1h�lm�r(��#	�D��IV5F�Z+i,�Ũ��k�\�X�b؍F#��RQZ,��� �rܠ��d��b��F�@mFƆ&#X�EEcbJL�ܮ�,X� Y�e��z��oz���=��E��Su��^x�j�\o&kr݇�,+�,��v�:���9�l�<�6"�]��lq���g���6��?X<v箩є[uv��q�a�i9<n��tGmi�ɹ�k�;\�q��[u��������dl'*�H]���A+�VŸݧ@[��L�eE�㖵��Q�H��f�n�m�L��{m]�r:9[�1�V��.�&��"򜝎)K�.�R���m�"h��6f�.��m�	�	4���ՃQ���Z�=ڼ�����J@�v�Zk�6 �A��p�؟��J����otE�;nҠí�C���f1wV��2�0��np8[nf�-)�tn���{{�𚙎z��z��]u��xgl��?o�>՝6ۮ��\��{��� }�E�V�ڔ,�n�mY�E��d�bpG��LM�i�r\&�3�"�#�l!�@Y-9�tfN��/��HS[^����޺���-�gP�%���(<n�����%���ln .mpo��	��v��C�Z���<ģ�	]�v8�H�XL��
�C,v�]e��Y�-���^4Q�Bݜ5� z� ��:�X�)kv�c`�a-�a	��d&�Mu����$�����Ҏ#^܋���p݁m�v�>y�q�J�NP{)Ÿ����GI�����+k[*v,n�U����DJ��n�:�Xܸ#`b�n@��8x������f]�:�V�!y�1jgmT�6bZ�u���͖���҈��3j������ݑ��)Ѯ��fɬ �Gr�q��;B��p�7����7]�*-�(6�.i:�m/%HV���Vz+U�ǟt��m��ژ�ijҲ�k�D���w�N��S�e�2��%�����"���z���9�d�3�Hp�<ts����{���m�U�c�!����]�y��0��/�J5�tg����Kh�L�M۱��ٺ[t�GG�=ל�r!��~��v��܎��na�'�]��ۋ�`*����w���瞾7�Lr��YcM �r��[��+�a���ZH���I�(�㋌�p�lF�q]�B��<��P�l��B����wo=�^��Q�z����0����n-�W]�lYl��x���g\bar���w`D0��es˭A����K5�q��c��r8u��Ī5�15Q.�۴� �9�B)��n5�]3�B��nr��������@�7S;,������vᬺ��.�,��B`Ri��ӡ����R�ė�KBfz��,̔42 .�/{ͬ�E��9�3d<Џ�������*#�a~c��Ƅ3� �h[��%L32P4d R���M�Ov�55W��G��|г 	hCa��@R�������k��������y1%�K�RC���'�9�;Ù��ѹ��B���B��2A4,̐)4!�̔�l�.�=�~}���{9����m�����䂤Ї��B(hY��l32P�32P-9>�}��j9���	��hC����.�e	SFd M�=�{=�:�g~ȉ���hJ���@Ћ﹚vHϜ�>��������wrP��І032APЌ̔"�B̀����&v{hGwܔoΰ�{��^���l���6��HЇw�B)0Y�()�Fd z_[�˞kn�,rDu�!�69��{z�u���������.d��vn[=v��vd:І���*hC�@y(K�32Pw}�l�{��Zc����ЎfFm��nt�e {}(F���B�a��������1��@|���r��E�߱e4FT�)+��0d�*�5�am�B���o����grҰZE�b���"��p��=�7��4��7ܛ�|�����?�g䄐����G�
�l���ѿ��ʍؼ���#��&'Pܔ���&�n�"ZfH���%vd�P�a��P4� R�� ������1�H� _=��w��l����$�� K�cAy ��/�HE����!��2 %4fHPЌ���;N�ɀr�Doe v�@�Ba������{�Y>�{U�2����4��\�������ߨ��#�
� J`���w?�t�����C\��e$]��7�Ϗt�W��;����܄��$�U�ן~}��aྱ������X���1�I���ʲP$1$�"�_0��j�~��;b�����
���W���l�1cÊ��twL����"�1$�V�����e�������������;}=�\��ס�[*�p���cbG$I����>+J�z��$f��O.��|6��;������3�Y���ek��)�}|olrvs;�E��w���
����(-���ZF���Yao�>���������_g4��6��)#�l��y�|��s"j�`�Ǳ	#�|��4��\�����bnp~��}��T�#�BH�F�Ip�-dv 35����U���O�wHf{�׬d��	#��Ή6h���<���2F��ܴ����Z���V6ƌ0 �Sh���DPA�Q �i�TGg��)<�	ݾ�#��?r�Rsx%�9��5�;�z��9�0�t�\$�ol�?J�gޫ����R����$@oF$�{m��c��fx6����0$RG$W�=�k�d���ʯ;�m>��C3�u���d�I��G��K=��=P�]ܾ���k�����qRs{얇oM[v��p���U������:9��i��8�wn�"IՇ�`��IMT��������1AKޤ�!��WW�����]�3t�U�����~���s�$I��������?�u�뫚��%us;�l_t�HĖ�=1�;�A*���I�J-"�{ =���g:�qng�t��4�_:�[��E
h�J�:��[����~�ٍ��k��t�x��R�U�L��t�����$�8(�u�Y���;"ٞ���:)��GI��2[������^��������l�$�ՏD�V}^akɘ->�Ϸ���ޑ|�	$�$c���{�7�^Ǣ��E��s�cq>�k��t��sB�,�
�/��~��rF�癩I�]^��2Ow���nw=�g)�����o�Z�H;"���[��m=�����3�Ry鹓����看�M��2,5���Ҷ��{Jm��ε�`��7|n�ݴK�e��=��:b�}�| +I�q
HҢe@�k�SCXr�8�m��"�� N1�5�h+w.���w=�y�,�\ٺ���6�V�Q��թL��W/�q�����h7�pXx6�ۄ�nC���n:�{;qz�۵u�jL�+D®д@��dq�ĭc5͔�Ԋ�6����r����r����YV7U�7�K'�]��1���]�#.� ���x�qbm����5?��1nGF�z�)�`�m�[�p��e��b\Kf���N���@^�ݡ��{;;�kr�u��f�;�_B�q�i�<�����1"G&����:c��/��{����Ln'׍w���Wk��L/��r�_1ܤ�v���o��$	���N[���Ӟ���)#�HĈ�;�^��&Ȅ�7uOggenW.��4}.p��m��y��~����$rG"�9�v{jvՉ"���G޼O��6�{�1nM�}����X��w(��%T�"�a�� &��Mi,��ȍ��\�zӁ���=s���O��~�ϲ1�J���}�rP����m���.���������F��#5s�ܲ����ܶؖ���s5�m�X\ɻ�[9�M���z���r�Uضc�j�{F]{uo�$�GN4EG���:��k�uO� 27ܽ��+ݿ;�q|����꟣��|6/�c�jQJ&���K�H��}$cwbә^���?(��N}rj��1{��#M��IJ�$�606)w����Ļ�IǜK_z��B�krX�K߇w9F$�M�TW�oOem����'YP�W�v�vw�����0$f��*#���G#�G��hJE4A��D�nl]n���y	��7[�D�KL�T�a��b�:��Ν��$���k�{)oY;^�z_�׈M���Z3w��$rG��*ͬ�ic���쓥�.��{�ys����ﳱ��HsH�%`�lw/�zI�/��g���A�d�M��ֲ���=�*ő�i�k(T9����ޮXpec���Xi�j�m:���=��!,�ћfQ��I3�gF�O� ��g����
�z>�}��������-��w��ɡ+]����;��_�޵QN�����k7��������ej�V����$`H��1$����7U�Ľ�_^��r�\��ñ������$�;�U�c۱J2���tE
�C.���eR�!�meV���ȩN�����ܮї1�Ɵ������n��~���r%�×=��8;�{��r�n{��H�z�݇���;}�d�����xc��d�r{���L�J���;����@I$�$��O�پ���<��������I,I�}Xh��7b>���ھ����n����d�{�s���gx�T'{�����SP�{b�"� �F�v�����6�n�'-<��u��*×��u�Up*�M��iw�uXś:J2�[u��i�l���f�{��HB�y�f��E��wr]�ܢ����~�l��bI�
^��9�#7���׌d�"Hs����>l�K͐�R��!vݜ�Pڧ�ϱhˁ��m^��˷]���v$(���V�!���מx�J�!%���_|t�r��I{�2����$bD��{|+��5~�d�=�N_^��}̗;��������_j�n��/�-�d�u�t���D$��!9_<t����gף������=׌d�$RG$a���:]�/<�H�ݠ{Ւ����j���؎{�Z��y����I�G#w׾2m'�y���t^��{�{�\��}�I��X�t��>����>ov壝GZ��C�eI3xV�2�ϥ�I���-��oz��#�
�&��]��M��\:�W>;ȧ]�H��p�"(����ykA�B[�"�<x��ar�6R�F���������E����5������!lٴe)j��hh]�hĶ[����jn�d��u8�����;v���XKQ��oP�)a����b�F�E�L�l�q�X�^�Ռ�֭[�p���[�b�6Tv�80&S@��jGB[`���[Xhi[�,F��w:��~�~�E<*&BX��.�XJ��T"�*gn��#G����+Ͷ�f�W���1�BHē/}��?d]��Ԟ�v�5S���;��dbH��.���5��X�޿jf��W�اW	���j���-}%}��nyv5�b��V|���I>�3���kr�l��R5��9.��gx	��đȾ�0g���A��}��n����pX#���l�����նĮɘ�V���d�H��l�!dfڹ��o�Q�>��^v���v0;�����nV�	i�ZF�%��TX��(�u�f2Uo�=�9��bb�,�A��g���緽���"�I�6��Sk�ز]ݾ������q�u�C�c:?�BI$�ބ���4)�OF�u̼�īٛ~���H�5nd�(��WU��*�/)貱z홳����I�-v�k5Q��cծV%�$VA�v{x[���쓞������g�+3�������j8��z��]�o $�I�`�ռ��yj���/v��/i㝚����oc�F$��NR�y�M�?��_!6�u^�z��JN��wv�;�ꋣ3����!$c�#�}��$y��Ś��3����t��<����:KN���WT�x��&�mӪ$=��њ��\�7:H�����b;o���s�z��Ձy[��Nߤu'.��ȫ�u9�\��Ue��sH�_��~���n�����^�z繥;��m�'�_ɲQS�d&n\O5���H��I=�=˫��-W~qݕz��u��Y��!�ڡ�pv���`��Jt�w�!/BID=���X&>�.�ik%�x�Īi���2��z�i�uwx���7{z5�M�e��vuЫ��ff�.\���W[n�S�*�����^�wZ�Ԫjvi����J�:�R����8X�}�۲�ӭ1��ˎ���k�Cu�RA-�w}6��2�p���a��$����dNt�	�f����e�駈/bPś3oo[�(�Zo��[�u�f�7�� ��FgۉmcX�ɥ:���1�^W9TE�d�E�e��:3�_X�璑�vT���w�vM���Eq+�{���U4��vS�s�JF�_^ˬ�]&��m�]A\:�1BP%ؕ�����}	z��X���˙ǝs�ku��`��B�3�z]��8��c0P���I���FqzoJ$�E�n1�3m��{��R���-�W�z�M@fEx'�2ަ���͇}�+���et	YtU�:���J���Re	"�k9u�M�BL������pԺ��^��\s7��d�p��9<T��n�bs[C6>�C]�E�^-;y�����������ײ������j��fۘJ贞m���j:��$�:bKT<!�8V�����) �gZ�������D�6ђ�w�8/$�[8���)R]��Y�i���t.��U�|v�:̻�%uJ괓$��^���ݜ9چ�����B[X2�t�mK��:%�(n�y�z�����zpa�f٩�gh��3}w������}}������&��cF�Z,��#ۛ�bآ���n�-&-66*(*E�b*�[�
MlbѴQh��}�Q6-�lb5����#y�Bm	o:]ݍ����h+Ovܼ�*L�b�˔F[5r������QPZ-���F�\��E�ڌA����,���b��E���QY1a5=�
61�X�Z1FJ�r�6*
L���[}��b��W�����3��'�%�&����C�~�{��z-�
����8Crmh���耺�z%R�;�l�v��?��I��;��ά���2W��>����RN�f�ל������Ք<y�#>X�J>R&,kl�n�;;��b<��:6m�\�C�*L�n��9v��\�E�|���j�ˬ�3����;��bHđ�������wj�+/=� ]��'ga��iѯӀ�D��wE1j�]�Io}�r�cկm	��$bE$�f-��Z��[�[K�x�m�'}�_�[���}���Iy�e5���{C���wU�w{����Vd���ݘ��<o4߳��%g��w8r��^�sdZ��z���U��w�|�[Y��Z��y7��j>ޞ���x?;�s �w+C�%���y!$}Y�@_�Qwr]�wr]ߥ��"Z0]��x6��o�����*��m������{�V[�]�# ȋ)P*�K�@��n��:安�k�A���<�f��m�TL�a�4���E��v���wy���g}m�'OZ�ϥ{Ǫ�p��z1"�?���c6��tW�wd�v��t���ҧ�Vf���.��_n��ws(��s=U.���.H��]2ZѹUۜ��%o���������$�	#�
Ʉ���Z<�}y��dF>��<��ڧӼ>�U�$ӂ�{GH�ؤ�	#I$~'�{2�g����羚>�^���6�;���d�,}$�~��0�F4���b�=��y�pT%�x_���ATk|:|��u���;:�.n�J�E�{�7v��ϣ'�29>:�$!,��DDD��*7v��98�ק�	�:0g�L�`8׷!عɮؙ���d⬎f ��8/7�����<�v\�eY��%6�3c�bl���e�������uq���qjAӰĵ�����A�n��i�[6�:�#�c.d6�0@ڐ��k5���`��wE=>�8S���k}�y)rj�Vv���F[LB܎��mٌl4��4t���y|�L�ݮ��R�bjd�FYLh��l��&�ٮ�\��%�B����]��d�w~�.;�:\��Ի��Lz��ނH�_I6�P�-��V����Ӹ	9^���w:�^+�Ӽ6/�o��Izx(x�κksv���wsE���$�#���zּ����6�;�vc��D>�1$b�8��_�]��'�	߸E�;�&��87}8gY����c��cv1"F$�Ox��k0�Y�LatՌ��kudΕi<V���d_f�I�Hv�6{3��i��a�H9M�l�=��쑹L��Dhh�n�ڏY�6_7:����r�H���r���7��2��Ց՜~�5�� �BHđ�=��jy���N0���e�1jw=� ���:ed�G�!�}����a����e*����[{���y�+s���pMk�m�v��		���}���=�6yg�C$63}8�Cen�e\�cF�zN�����F$@I6��[�a�Y��S�(�w�3z��$����p!��5��ֆH��H�͇wz�uv�����3ዽ����qn�݃�w���I3�"Hē9�O�Z�s�/��[��Z{���o�	�H�*�X�h��ˍ���f��`n��Z9�[���鬸� b�0%�B֍�'Ti�i==�Ly�%�$j�\��J��d�
���ⲘS�M��Cd	 F���)��t:c�l��=�o�w�ڔ2�xvc;��]\W�]�%���+�1'���$�`ܯ=v��w����&�ێǧ
��j�'���I���U/i���J�>�ҫJ3]�����x���J���3�ɋ�u�	׹� =��~��{��;��o��w�^E��\�X��Ul�TB��q���H�٩N1OA��<�;���;{5�r���=��`�_I�F�N����n���ߴ�=�1.�w��c�gt��M�C+O�n��Љzz�n��j�3I
hK�9��b��ڍ�T�D�H6�/>�>b����������wn;G6�a�w�3�F����c�I/f_o���ӧ)������3B�[�<��d�|6 3y�&��0��me��9��"��E{0��I�V��k<==�1.�w���9ȾG$����=��_%>���[��^��T��;�kQٝ�좲n{�!Ѵ/]ZN�Q�L���OK�������&^#m)x�ŽY�MB�t2��U!s6��;��J9nJ���}������NbE��G$I���4��.��T���4����/&��w�ټ�IwyA9:�"��KČ����])a�X�;m�J\���X�a�mY��S%��2ꖯ}{��I%�$c:QΆ��}�q黩���P��sȽ��~�	#�H�W=+���~Y��1胻�8w���Z�K���:I~��%�=��g���{���$_	"�:�ק�r�.K�nU�^msx6w�؇ٽ$�$�X^׈]��fݡ�G�t��%�����wS���������4|���{����_	##�DX�)�T��������=�R��g�:ĒH'�/�B��f�ɐ۱YF�f����iK�(�0<\��Pںi�����]��@](����b��.T��X��rr����hg���~|>\~�E����v�^"���m��q� ]ŝ�#��m�Å퍬���H౺,��f	[2��ʽ�x۩�/G]���D��S�]P�r����IH���b��ݵ�m��=ceۂ�v����T6e�;����V6���r��h�m�bΚ0���6,��16�.����X^��"�n��^Lp�;�<����1��(f�nn��#��_?�?���9�=J�0�:���ł1�M����X]�Q�e�7����o�K�9�Or������d�}8:����vȀݭ�CwS	ʯhV8���	�}ٶ}����z������7��ר��h�]قr�9����&IM�q�6-y�sFL�S��=Of���$`I��#H�<.������wI/�ǰy^��y���	�ﾑk�q{s���KF�I]��ͫ�f:�qΔ�Y�y8}�h^E�Cw|N@�0�S�f�~��/�-�l���
 �t��5�hK"��l*�t�*A�H�H0AJ��Ht�Z�{��1%���vq���W�;��y�a3<�;=z��LRsHċ�"��
Ľ��;�H�h�cїĩU���D���1��S7�;�
=\u��&��dT5��q�k��u��z�,�Ưa��� }�������f�ն��rJ4�l�>ͯ��@I(0��r�MWs���I�C�k'�+��͖"��s'R�g���օ�[�H����y��V�[�oپ�"Wb	8�oG[�{��w�ھ��馧;ٷ��X�yȾ�1$bG��,T�!{����g.�Ք�NiF���n�ّn��w���s|����+<��b���q���27S���tc��e�ʘaRl�5�J�t3|&F>��_�H��Z"�V�wR�g���+.c�+��P��k�/��H��Vr�O��������������=ԤW,���F'/���Z���W��t�	$������gs<P�z�m��tc����ə�u�S/l�Ar;"�2$��&�H:���N��߶�����j���[�S#�6�^�!k�1����}�^I�vw6�YFt���/�y�#E���7���ۼ;���7u	�D]�[3��Y�o'�h/E�)X*�w��ޒ`���H=%v���s���4w���ͯo�zwv���u	 vq�fyv�?{�Vy�	�$2�0\Y������jn��Vl��[.������R��}����{��!$c5�i{�{.���N��!���e���E��w��>I/奈M�q��k3�"�nj�D\<�gu*w�����й���Z��;Н��!~���wP����׵n�s���c`�7���i�o{�o�����$r/�pR� "�|��&��Iٯc�K���]v]R�= ��k׉�w���o8d�lnQ��wD������d��.I�7��zs<2z�=�[�S��z�Fj�t��Ո���j���z�	�c�)#�9����7ke�����A�;��~M���B�-������f��y�{:�y�N�b�iK��ek��m��*�&��LMC��˦�%���z?w��ٱn�����l�ܶ7�O|^N��X�}:ᕓ�Bo-�[��ru���Pھ�Y���}��9��ٽ�ݡ�۲���T����F�I��ʞq��9�<�ǜΔ|�ɻ�f+Ȇ����%AV����߈=̉Ҿ���W��:�v�S"[�2�q�LYt:�|�)�(3|���d��"D�|Ȓ1@ȕ��twv������׋"�>y�ީ���ټ�2W�f����|D�X��h��kj�;�ОhIU�׶�RȎ{�cڵ:��sҼq��6�̉��SU�=�	��mڱ���oge�j���:dt�v7h��m߃~��GL5/nk�	��-��g�i��H�����`��D�V������1���PN�;����ޚ=
�Gw!ψ�ǭ+�-	�z樗9�4Ш���y�kfn��Y��[7;��<{��N��fN�V���S1c����$r�R�5T����Ȣn��o �G)ފ�2ʨ��k��:K��sөKo�
N��Mr�@uU�v��[�����9�j
�1^�7v�u�����{z�@ĵ��NV���|�~2� ���ͻ�gp��*�״����a�z�陳.�Z=~�n�<�^.�ژ2���X�vf���'9�dj�Y)2�[���/����m�XP����v�U�A�T�a�Ve�od�¥��cy�n驨SiZ/cYi⪭\�u�M6E�.�B��UکCw$��菰fm��m��ݫ�9��AI���g՗��|�ٜ���L\MՌ>�/�Y��q������3j���P�c�u�R�,$̭�3o�ƊbC[Y[S
�ޫ�n��N����eK�4���֪߄1������T)����#���۷��8�U\����v��j��z)���D�bh���h&��ط$7����3l��R�������M�/:��!�u�lb�1�T,�Gz�ә��n^�L
4WJ�p�1��P�iX�D��A���=cs�g�b�x���{�___wƾ�ƣQQR!�>]6,j��FkF,U/-�t�QEr���V(���[r��A�nW5b���O;;��U�j�{�{��wu�scr��(�#FأTW�r��o7A�Ŷ�r���y��Pk���ɱ��LTO;d���,V("�5�e�m{���j6-��ܣ@r�\�[��ݣo��ǹ~~1锣4�+%�M�Z���);��ͧw=��E�Yn5�V^���^�%Ð޶
��%'�@�����ol��I�"E�vǛ�����+�3S��]b��Tv�ë��on!���p�@�-��D�Py�͐v�������6H���ŰX"95�T����]�#Q�3�n����X�vҹ�9b��a��c����3�X�]��/U爹�!m�E��˹� `'l�sƇg����]�bS�lYf� 1�l���[Ohe�5��12����nd9�Ѵ�ǂ��m�<�)���e.;t���B����0����zz��s Q��f�h�&�챲�4b���Mu��q�>��h�$B0�s�J̷EH�Z�*7�v&���,�h��"�c-�)K5]m�e]9�6;i���jU7�#k���Q�nɱ�չ+)Ka��f���qa�6�(�V�R���n�vkI���� �[K�+4y�賸5úC5�� P��H�-���c=���`5j���X4O�m6.�Уy�q�Z�C\�������q۠�n��m��̫�"�;���X^9��O0��>��]�wb��V���6E9
��֮��Gnl]�í����t�j�8��k�t���b���5�x����h����Ch�[e�Rt[c4�D��W���G=F��q]����<7�ml���I��N0���Sd�F�y&�j�3������!.m!����4@�ۍ�4#��	n���>�9�z��C�vq���t�\b�4�5��Fش��!S\��ٰ���w\��d��t���>��m��q������[�ƴE�9�����`�Rj]��iR¹i��z�@�e�J�+�YѪ�g���ƹ�3]l�0�utB:�`JK��-tH��,��)!4.�+.�.���7C��GH]G��At�����W�-���..c������3����Z� ��㪫W���>��;U�U�b�M�5jN�ljs�l ��J1�ah�#������V7[l^G�7�W�m��7tF@����;���v��qv�h�����2��^1�Z�O�Ny'�cqu���=s�V�f��X��kY�$�)t㙉}G�[�7j�%ú.v󄆮�d[����'�vI����f��Q�Y�ipb��bPj��M�ű&{�M�G�<��e���]����uF�t(���T;b�a��H�bJ�UC�Ee��Ƿ$��%1���mA��z�}�n�]S�4�H�ݼ��KF4wn�\).�w�J�$e���>�w�UW{����?lA~����waj�0���G@�9���lʫ�[�{��n���_$�("E�TM���ݹ���t�MmՍ��%|�R.�+�$wp���w�˿���$��A;��c�6��S;����h\�ݕ��/w��:�7��e'�Ħ=�E��P��"�_ ��\:Uq���Rv�h�'e5rz��ˡ��ݩ�~؂;��ݎT����4�q��B����F:M�	�Qk�����	��BSζ�@(h�=�������`�1|�=�B�2'�	٫b�]z�d�EV6j�=��nѬ�W�;���U}"�D�$tEW��W�Z��*���V��ՙ�cr�َ�q�z]�o-�u��-:ʧ�Q��o	������G\e�=C��uIԸV��T3|s����]���g�-�]�}�z�]S��ھ~���DǠ�㝂n�*A��QJ�%���]�)2�E�[�Fs��m�H�͒rū���4\v����x��>�:��AH艨 e���E���ֈؗ_aOs�R ���C1aޞ]�z�ңk�C�����o��'��ߑU�R܅w���i1�o�!`�8���G��B�w�W����z��U�`��_2�+�"`���Sݙ��#��f�\K��d���������oE�5�lk�S�g�4،�3Mpχ��K,��	�7u��#ungx��o�Ԃ�=�D�E+�o�ֻk�w�2	�:H�2/��ح�G���1|����q�<��q��F���d�F�� �&e���e?o�[�1 ��y���a�d${G�z�:��Yw����`�R��Oa���)K��<}��T�m�2���gK~2V-u;Ě�:�`�8�|�pG�tem���Uu�%�����}ީ����{� Nu|�"f��k  ���D��d�2����F��"f���/fgY;}��d==�&��?v�W��~�V��.���ȟ�n�� ȾM�(]�a���~�g��<��]3u��F���`�) Af��#d��D6Ꝋ��
�����Gh��n�s·���s�3��[�� :B�&uuu�%H�������a�"�2G�.����jy��R��jkÀ�Y��~����Ld0D���L���.��8�
���_��?�j�}�+o���̃E�Z��GD��"�m;w�X���.U�$c̅,awtS��w-�Wۙ�#{���I~�]T�ww�r�E��$�_����ؼ=x�%nV.�K�9��Lw)�;}�j#����dd�g��m��z��.�fV޳V�ùv�u�-��F��{�T��ԫ�忢]W
�j�dtI����v+t�u��|�̾�'�ѹ �e��A0�Gu��;?fp-���{�K�'���A����;ڟ�o�`Ș �$}�g������j	��t��3��\q�[�k���^�����)���0-֪�SF�!��@9��FD� ��a����}�{��ڍ�N>��ϥ�~�mx�~a��(W� ̉�~2G@��v�"��O����{S�r��ڡ�6�1{���"oP�"�݈m'���,ڒS7v�,Ȕ�w$�]����4��o�:��M�3 �S�_w�{W����|̑�6.�؋5`�h2&c�E�;/���4��	"�@�;��9\�R��t_n׾ �wu0A�A�PvU�I�����NE��5C�|Z�(^�0NyA�M��E�#}������B�z����!���/�֑Dl轹���=e��Rɒe��J��-F�(��mGJ��v�glv�4�+a�E���>��"�j��B��Z�ez!�NN_ms]��q�]u�Z#]�1n��e��:��Ͱg��I�\)�d1p�F2 �k�m�[ �]JJu7
`(M+�5�%��D�. )),t)�=Ȉf��&� �8��M�� �B����R��*�,�R<7K�������kX��L���v�QAj��ݵ�-��q9�;���++=�!V\ix�tn,]�����M6��q�����SVD�=�l-��ӱcY'��<UUb�c�;��YJ��F�3� �݆d�b������w7�X�ĎJ����������d��"F�D���)>Bf�`���lA���}�{��iQ�����|���$[�sh��SNO�_0�j`������?Ib�ݕv�/5�. ڰݾ�"�/q}r���.0����#u�s����{�ę��d��|da�Θç�����]x�A��GD]��
��y�"`�z:"F `��	#�D�"h���o�8v�xl��^o�Ш։'?��7P_�U|db�٣�nWj�{��Ik�a7��9�h7k��sPءF�魔�2%H�L�uP�ަ=� �|�n�')��}�/{���-���*p��̤V��|g/��2$�_H�	�
9J><=�*B�i������G��`Ǧ��Yx��ظ0kӗw�,�ۨ�WS�S�I�P��^�ɒ$ɤ�kSQCȚv�6��O27���?$������O6N_6�#�gs��އ���=��7�3"􊾬�Ta|^���>`��2�P�"d#g��W��݋�w�����TkF��	�H�$����2/�ή=�[=��eͪ�ZA�A|d�A���w)��}*��[��|�<�{�/�Q�2�����L�����%P&D� �`�%�Sԅ^=��d���Ae������2i�R�x�y�[��ș�d����4׻l���!���X���s������m��ג��qe6�jac:Q	QE����N��XA��ٳ�Os����TkF��eTU������W�H�D�?#��Z�>��X�����wVGN�jҫ�W��/|'<�`gu
2-���r��n�}@�90A0�"IB� H���+�J����Z��0��u���y��52L�f��Ъ7�<:vE����/��]it]a'o:�$�1�u�����S|����ve����s&�UO]~.:7�0d_3$t�����lϩ���!ݰ�ݤ?n�����8����JPn���@=�76�J���^��2z������� ��%~92���Ѭ�L�'ӧ�y�RR��^R�e�y?gu
�Ș �ö#����v]�b�2�ɭ�x����ke�/br�!r=�<A�@�t%:TYt���?����A|F�	y7�49�&z�zXK��"��U}��-xw�*�����ؘ �#�$A�dA��n�5CBۦOs�>7 �0�gXs����jZ�w���L�#$�8����sO|'���j�A;<�"Șd�'vj���U]޿y5<��"7< ��gs�}"�"H�aW~�]����a�2z���C&��J��9��j�����\__6ru.D#����v�J����[��w--sn��d#}�s�oZ��d�:��s7�^���<r��ͧC���w�����;�K�ȓ��}�W���{c�L`�"d�(�C1�7s�*C@I�໕�7����xP �&A0ȒP�%ܕf>k�FGJa�M��袃@+f����@��JD�tk.��Y��_��Y~���g��D��{|�n�����3}H���i�>���P���J@���n��wi;u�����r��#/�Ϣ�/کa�|�F6�w\��Gj�^����U��?���	�@9%
 șP>�����g��>�s��5��љ9�z&"F"IB��}"�E,������Y��>z0�;���:���n��Dq�>��/(w��Ǽ.e��	�����L� &���2/����K�TY,�ˑ���� ���T�θ�KF<^�~3������$y6���^̥��̦��*u��k����W��8�u|����ue]�D�1�49j���~�Vo\���*^�3n����!���Ok\ʒ�6M�I�� X�}��̼��2Ͷ�)��)�%=f�]8����^����
[����B���a�[��Җ�
4F[��Ի0r	��%��X��[���h��J^�'gO'��z�R�:!t�qn,4dn��-�����z����\���-��{Dv�1�QX}���ll$�\��6V]K2X�M2�w��`�~�;\\��t<m&{-�Z���"l�ZMj`�1Y�������e�~>�~�FE���'��Ϊ����Wֺ]t��;��T�O?�G��&H�~Â���W�A�@wG���w�w��}M_Z#7�s�d�_H�^�lX��0Gl�_NLD�?��?�H��+��f�1���Id����6X�1�}���D��"dd��0ī�����x�ˡ��g:��2m(vj�Fe���FL��m"
��@ݱ�U��Պ�^
#��}_F�D�#�$_H���^N��@#��������Z/��8��_\C�FN�FD�Fѝ��?{v�,��͢������܄�vv�;:.�i<��m���! �f�ᖱ�wi�@n��+��<�ۊ&'�xl��V/��m�꽌f�D���`�d��"F�2 �P�^{����孮	4;��z����Vxw�_�����t�{K��sGv��FU������K6J��qT��g��A�.�6^W{�J�=C&�*H���\^ۭ1% A�u����5g2�n�iiw$�ȑ�;��1��% �#[y�4����^��g�n��<][�C3�@�r�W#�� ������>R��-�_g�Fg7��A_�e��t[�v`�1��N�LdT�Sku��x��,��?w��"F?d�(ȷ̮O�X��`q�����E��ˋ�u�&p`��� ��}~�g�)�y��O��̬@����Z�e&M�!]��iuۺ�uܖ���D�tƟ�����?g/�k�A����F���/N"�W$7|l����|{cv�nJ�E���$�@�"dS:S^��XN7�q!�ݫ�.��[:���f��=���&&?v���{k:��0�'�h	�A�$b���D�!�s���]h�z3�ۼz�}��S�3-�wt��/���e�r޾�'\��UKY=뢆!��h<_]�4^�f%S�*����;��0�'9wnX����7����8���)�Q���#��j�L�s6���M�Y^,��Tr�M4���|w)��'Z�	-��O;�v$�<�;�f���v�	y�1/Q�v!b�z����J/�EV�;[��������)Nܖ.w�˫�ct4G���95U/�a���Cz�n��\VX��U%wkr9)��f�.��ϡ�AٙF�n����n=o�h�fEsԟ��eg�j�k_J��ҧ=����k�̻������q�PF�T|��";o&C:�9�͚����V���O������+8���\s�F�
�׺]���Ł�J��]��1n�NL���i��o�3��07��Q�5m�Ea>�m�󻞘�]fj�����BT�!����VB^D����]�lru��`A�x*neJUn�s��l�KÆ��n�u�z�����*��)�UۊO�%-;�{�0N����֥M�z�l�&�2�6)��D����ǒ��A�;꼾�A]fݷ��P2��I�q˵������h����^�BA*�a�*��M<<83E��M�w[e�D����qU��b��=Ŗ�����5�]B�wG���O��r�\�6=�����W֚�d�}�杮:U�y2����<��D%d�ޥ��ӥ�Wfc�����7N�7�κ��F��[W�vrvÇS��?Wn��|�1�C11�66�Am��,%���r6,[EX�Xڞ�n[��Q�j�����b�W9b���u��\�ks���Q�h�Z+���]5QV6��[�Q��\+slnkE��X��\�lE�w�r�+��\�s�(�ȫ���,E����r6�u�j��w��0F���9��KE\���1PZ#}�$~G��RN��w9����P'y|�0ȒP���0dL3�}9$xs�����"`�$u�<�g�����R���|� ̠�"na�<���h9��(0D��v/�BȒ����u����+�����^�vh�Sޯ����ڂ;��	�9/޻-
��\QOS��L:$��<vb��ύ�:��#���y��Q�ͳ���_�	�����|d_1#})�99���6�FL�q���H��UP��$��T�w$�w
]��2�98N� �f8���Z`A�λ����b۾�mrC7��js���e^�N�Uf��.��u�P �/��0$�_�Ed�&�	^����5$�4xT~��j�#�d_3$t��բ�3��;�f������D��&��^���LPoo���?n.�-��Xk��E���mJc��٩��9��b��K(�wܫ�+��ߵ�ƫn69�ȩڽv՜���F�*'�C)4D���m���x���r �$t2?�^��܈���M1�ǅ�y�w|�ܪ��e9�B�2'�F�K6*�xH˭o1�W��Bf2Ĺ�u�7O�9�s���:���t�WԘ=ҁ �_NB�G�	g�峼�S�T��Q�p#k�̗��ko����n�3g|�?I#H�>�����L�1���H�ڂ�z{eo�G��FL�'% A5�݈3-byR��d��D���41��Wq���W��g{�o[<x=33<���r�f��z 2s�2���U���{�]ܗ��������.���T��G������wm_���~�W�w�`����$�(Z>�8-���oWm�����=�Z2�J�6����������wr�j��w��Ǧ4�q�'���L~Íz�~��X5e����e���C=WZOqj5��o3=��.�о~}}�譟=M�M��XڨK+(�,rs�@)c�k6��"2xdT��mo���i��i��H:�Z��^�ur���G���6�+��jy�qZ���@�5�{�&Ӷ�,��q�Z�����7j8ݺ�{mAo�y�����a��õu�y�9�U�:�&�)����H0!�S�sv�s��rU��֨/$�B+���J�Gm�}��/�|�k]�u�����HP79�2f�R�(�*���v�h��C��}���3"d$s��{NMۯw��rCg�x���o�1��(辑"H�?�@�2�<rӭnP�G�7�ȇI2��mX�q����N�tta�dY�u���7P^�4����	�A��P�dO��Rk�\�yvK�bNu*v(7;y2��}"ȟ�[�f.�G3�1�ܬL���=�5�V߽�Hl�`��?�-�4�A����� ���;��uF����y�f_��O�d�����ã�"dd�������������܈�1�4��i�����0�S4�� F���m�1��霹0f_^�z�������
2'�H��ڛ{�7޵n9ؠ��~�_%��+���n��D0 �$u��Ҝ���RO=��{e�v�f�r��vk�v���(wy��c��ܢ�����6t5�l���V����X��g�����C1{�q�8�R ���f���^{���ʡ��f�_{۴����E���� ����� �`�%|+�>����s����˿U�[a�ǻ/��'n:��"�	�:"Fio�4#�yOr9�B���A�A�72�y]�x挹�?�R�����A�>3~/(�;̠���K��D$tA�F�#^�,��lϜǲo.S9m�����0A� ��_H�����ųr�׶WtϏ+T(��ؤ�[����&�6N�r�������.4ݫ�[��m�%2��R��Q������~#M��×����=j�N�<eۄ1��X?I#"dx�[��OzK�O���"
�u�_��u�9'��ˈp�"S��F]هٵU\㎪��S݉?f󯈑}"�� #�|�^�c}����a�5uE���S���W������F�l{t������k���.�ᕜˬ��B�S�t�S%��v�on���1�C���~r�f������3��r0�J6�<�Š���� ��"$��7P_v��v�X+���ە��n:_�c���V���Ϲ|�>�H�"$b�2,g�:��\����.��z�z�a��pfN`����5F��m�X�3*%��A�I"�I�:�\W���Az��z��x�9�\b�I����P���� ����2G[�<�U�3ӈ/�U�̓��?TW��ޡ�1�v�O2%���S.�JN�$g.���+.D�{�/�͵~'g���ٵ�A;q����m��%k����ܨ�dtD�2 �P�"d#�#Wiuo���ɮ����༜ �L�60ȒW¾�dL��Bk4qq�7���7��+d�g���܃fyW\����=�2�sL�~��[��µCr��2`�e�Tk +L}�Rn4W�M��&���/z�wW.)�wq]Ty�"�[���[؏mKc��&A�`I3��	dI.��Q����)>��\��~'���G��+�'= �A��d�J��yvo7�����uI�ke�����u��,4Gr�oN��ö���e]g{16np ~=����W�u/˯q�w�fW�pɃ7��&�.E$w�"�_n�d�����ȟ�$c������=��=9?�f���/���*�o|�3�`���Q�h��"<o*�y������|�P�F^7��_o����/��J�}�d�OJ��ᱍ��J�~�k�dO�	�:��c�n���;Uh2{����y9z�]��	����	�_,�L�K�~\�?�P�2/��: ��+�+���~�^yC��y�8��l�"k*$6!����(��ઍ���d�݊2&ea�t�v�wb�AYIV�����[#�{t�=���Y/P2�T�ԬF�^���ه2�-�PP��`ѕ�u�wL�A�q%0j����`p@��SH���0��&.gP^1����v�;��g�ޜv��SXz}g�#R�`�X�]-�в�3$^{E��Ek�Tz��g��Dт�i��*���(fb����,�̲�¶� ���۹��8|q�F��^K4Z��AH`c�����3/]�&�
�� [k4a�cPiE3�1DbR6�K��|�l�?́e���ǧv������1�C�x��vj��N�O����]/�H�n������L��'����_5~�m�f�����2GDH��"�R�/��u��`��/���[�׻�\$����)�A�$�<:�^��߳�����g������AH߫�U���Y�a�g��܃z�������3�9�E�_�I*����bz�k~ �a�Fί��#���Ƀ��!��e}�ߢ`��KZ�����;i�A��DH�&D���(�Nz��W/`У�Yo��o�����<+�ɀA0ȒP������ƸO��p�B�4ªE�L����6�#M)�la�D��Ew1-ɻݱtw�a�K-��륗�0��?�&H�d��.��Ҽ�˭hl��y*��]{{e�GH�9)|A�A$��"df�1�+��v#w�u}�`�ޞ���/]��Z��� �J��V����S�������أK4��3�e����iD&h�yc�#�D���Alv����p �o�2�۵w���A	�8��##`�dA���"`�#@�)���[�<�+^pu����3���L�#�%W�F�D�
���wumk]��4��&H�l��ۜ9�3��i�����:���l�J��L{�Je�ҡ�w�]�,I'��u�{t/K��L1s�^��P��&'3���r��[�0d_3$f�����|��4����T�\�[n��"M)�,ݛI��V�4\���d5srD���z��0A�gP�dL�0�˺�^���et70ع��Jv����~�W�& ���+�`ș�$vz�5�s�u*xe�;�_M�O7g:�.�*�~ƆJ�uᓨQ�ZO�_�es|�0*�}�FJ���}ز��}v����mޞ����ݘw^��&n��r����!y���r=j�},<����y����n�g��T\��&̰��}՘��d�!�[KfW��&9۵�A�#�LbӶ���6�*��!��;%
 �_H����ς��y�s8XΞ��3�;'GcR�2Z��A�H~;��H�2-��C�ھ=y�j� ԷBoyuJ˂�J�k������wi6/�\�������u�t���I�f�,g�3f��kkn��֜�9\A��\k�������J�r%�w$�˻�Reܒ}���zN��9(��^�k��n�T���t?{X`�/��: �dA����}Qл��A�L�'1�߯ς�Y��x��ɽ�`��� M@nꃙΓ>��Zd��D�a�d_3$uv��� ا�u�3V�]!�j񱓂�J}{fD�F�I~P�X�ߡ�Ȭ��7%���}���
bt5�KnW�s�?���Fm+����K����~��P�l����W�U��l������gc�"ֱK���S[���l�9Z�}��8~�7����>����?�2JdO|����e1ϲ��.��ڂ�M� ܥ�"��?��ο/�~����Q��b�M�km0��Ap��:Z][:N;k���p�E�����׽y��y��v�?n�y�]�b�t5�^62r�kt�>������P>��da�$��G����8��;2pd_k�r݆Uةe��uQ[���s�0A�""æ&�nOf�:"�"d�(ș!����e��{�Ӯ~��`ޞ=��A�a�$�_H�2'���+�j�_��?xO��r�� �$Owk�ɮ�wCX��bo�J�������Iϟ}X���2$�_H���$a�D���VU�������]���h���'o�~��D�?#��*O?%=wsBh!wHvQqRu�w�^A���X��e�*t���ޭ��B=g����i���웦�V�U�w�&yǩeJ�[�ʸd����ưk-��R-�:��cm6:JF����V���t-�X&1�S�ֱo��W�kY�'t�T�U�m��IF��μ�AQ��u��9��v�sC!
�VorW��XU#1���{���i�ۑ�\�*�vl��r�V^����~ʠbʲ߶{%k�V���R�t�u��e�,nx�b�.k��%��������-qiS�,�,�͉
����~��Ǝ˵���z��we�.�6%1�"��a�5�&�j�:6�:�WȬ����GY�X[/n�v2S���.�o��˩��і]t�R̵��z�wUZ��㛽�w&4���sY��w��nMurYsmM��=�5E+�T�=Z�,lɰ���ѻ��a�[��emc�����ΫW�^�`ۜ�+&���n��w7]qbT�F0庇�1��7�ʋ�]X���]3��M�����o6!V^G���1)�8f��};k4��*��*�S�"S�5�6�ӫ ��T��ɷuIg.̔��K��z�!��ζ��r�Xq��[W�~߹u�Rά+*��(3�Nh۬J���c��y�yY���u�<��B��-#c�\�3r������`�M�7ή��ȳ0�Zz�7t�k�J��oe�Uy����^d�18p���m�����M�t��QW%�����2,���+�r�S��u��E��X,�-�Wu�"�<���āԅ��fS��\;�?i��ܹ�u�r�����9ΛE2e�w�EA\ѷ6��"4$$E\у�5�\������nQ�E�]�\��9����؍�N�ʊ��۔k�4�u޺�6$�7]�{�y�-F���jSst�E�+�2��-
h���'v�ǜCA�,U���:�˩�2b+�h��HL�1���Js��b��h�FcM*7:lC#A�Q��L���A&�pƮ����Dlci/5s,!ns�&��|���[��4u��(��r^-�1
IR�QKv�����c�l-�ÓXµaM���X�;u�(���Kdv��ϑ�fA6tLu'W�0o�Ӳ�&��e�&u���$�[�N<�`�nY�ù����3秹2�,v1�����;�:�<�Qna�7;��#C��j}tanЇ9,�s�(vX'A��,�N��9n���º��Rsm��`7b^�1��z���]�YMٱ�7U7�f��r��o�f�F�P%�
���H��%)(ön�k��Ƈ�fP�C����<ޖx�@-�q[[N��{v�����e����Bok�\�pf�[nj:��q{���+h3��!�zR��u#q�Y�nk��MgX�f�����M� �]���v�vb�z�]��VK�)F��3qL8	(��1ƻn���	-L�Y��fj0��s���{�E�ju.�@	�����v�v2R�-lHG4�k��GK&�'n���x�[��� �ΓH�V�kD`2����֚iK0JZ,e렶wB��@N�sgD�Lk%d5�c�;n��G���><���s�ʡ�X�HOG-��S�5�a�Wgs۫nď��L��k�5{���,v��3
	F�X�.��7Yǧ�P�H�>h�T�ZCXS�.�B�n��1�b.]�v#��V�unq�Azɹ趩�rFv�@���S��l���81������ԅ��&)	��m�ٽYili�4����Mc��׃�[������'n���*vK�Q�հ��"����S:hb�ȡ-i)����sc)�a.ۤ�q�鶶��O==p�F3�<]<zդ�oC�2�P�WBXYY�1�!�
�Q���BYUc+��p''v��;C�.s��s�j9|q��\;�y�d�S7d�ae
�ϲ��������CǴwne� � �g[vWK�rf���g;%��mcK�B�ufҩ F6�KF��6�뮊�c��d89n۬�9��%�g���!���yɐ�Ν'9�эV�N�&F%�h�m]���j:�g����cq����{n���G6�d�vpEq�q#˟Fء�e+.�ѐX�h�A�4Yqta����E���o�ܶtmf�N��&����l:�h�m�L^fVhq��s33�D�f��xM���l�#)�T��6���� ~�i�ZK-ef�� z��\��f�q�D�)&Xm�� A���f��j� n����J�^�n7�a�;f�M�z* ����_�+��d��#3}�;��MN��R��wk����!X��bo|�J@��0��6�(C.��~M���E�FJ��g��Roy�#�8Ha���l7�������?�/��d��!��X��*�b�;(P;ɂ$A����o�=�ۂ�M�;��"��5�j�f���_�?�VA2GD#ȭae�}K�����l�㛔�cY��� 적������n�j{y�e�s$.��'&��b�W�Iy�3��Q�S<O�v8���bl��IӤY�k��/�s�$�_�az�x����H*ٵ�o�#~]�
g[�H��L�$tD���0�Ž'��o���8;�Q>�Upܵ�`kv��iZ��Ĭ^����1/#���xЉ��RY}Y5E���
н�1�Ӛ��(3�q�l���#}�<�w�s�&>7����D,�&�3��^�����\a��� �ӝ$A�?n�u��u�鴸�)�>�cY�����A�A:��a ȒP������P�' ����wP@z�eU�Sŉ�$n���Έ�����<&Zdg��$a�d@1$�@��ԩ����M�3© �]�ڕ���"�����jF��%
����2�(~:��7��G\�b�&�;�GH
Y�K���v͌+���ۥ��6N�	����n��H������wu07v�mMO9�+�lM����:�K�Ll�!D^�{ɐ~��D��DȔ��Bg7aeA���؃���ʽ.x�:D���_qˉ�&�@�^Ѫ/Z�d˲���n��0��� �?I(P2& �O:勥N��r����Z��k����3�mG��nݽ��9+k*��Z|�����B��9D{��_rշZX�̧ڛ�������W��U�,d�`�2�( �����+#9Y�qh����9�rA�՛�:�q<�!X�cc%2PD?U�^�&����X� ��0D��2%�u�����p��\�ɼv��&�ܕ�|L_?� ��"	��/{y̔޽xD���y�
�.��5��H����a�A�Y�VRg�e�Tt�m�0ؘ������DA��ݤ#u>�t��������*45ܬ��A��P���?��#��],q���C�r� ��n�����B����J�6�oc�Խ�{�C�s�
go��cۉCw$�$����@�^#��zћ�4�����ĩھ�;�u�y�"���:"FK��^}��YA~��9���A]z{��=��ݘ_���'�cd�ڎ8lN����<n�띋�WY�\+'���mκ��Y^���Xt�B)�B��W�U�¿v�,+ؾ�k��Xڳ�6��������d_0�� �"�G���x8���,i����ޗ����R�o;�	�AnG��_��>�e�>M~`�Z�X�m��	�/g9ͼQO]^�5m�n�!u٬6Įu"��{����/����2 ����n��w��b�ũڼ~hN�����}"�~�:"F do����]��ɶ0�ɐg����Vu�ΗeA�.sr���A�����W0 �?����F2& #Ͱ�4�`�87�~%-�d�U�]��x���,`�%
,N�5*�GR�A���ޡ_H�_����]А�qJo/�w���$*�u�؇bdf�$0L�$��N�FfEd��F��t����K����씁f��#w[�����JZ��K؏�e���kN�u]���!��
��4VͮZ6�긙י�F��yh���~8:랞C�#\S1���B�������*goA���V�M|~�N�1J�DV�+v�� �.�M��R�{�=��Y��e�������r��j�l�!�ܦ�0�3.T�Bۮw]�b�jl��ͳ4��V�#ٶ�UF�lo8�v+��6˵��v�Ԝ#�0;��j�v�mnuQ4��u����UB\��Ux���ŷgn�XʰK�0���Ln25�iM!D��W=M3���­�f�d����!��T3n'pA�k�-�f���i��.�,���嗭O:���	�:�a�ygK==�]�V���+`M��҄Aޡ�@~���r0Ȓ1@ș-5l����"H���A�;5��&�j�%w��w�`ฏ�����n��'�A�W�/�H��7��ќevAkoժ{1.3;y0F�G�	�+u-�B���q���JV����0�耒<;�{:��~�WX����w �M����Az�������%}@�"`��	!x�{G�E�ܟ{[9��9�ט��eUnJ�':� �2 ��0&H�eV����[˜%&��\�Yn�]J$!IvC2��;���r�h�lp(�v�����{����Jc[�E'w�˹:��A��o���T.���zh]l����>�%3{�Rj�U�|1�����w����TNS[թ:��|S�K2X�,����y�&Z�x�wn�觲m�ȗ�V]A6��/6&�X�Ur�]X��lSw[���p�t�U`_f�p˚�zՎ�����{���9uǢm�a�c' ��FNb���v>���U$3PKw��z'��L������j�҆�8��Ђp��^ ��:���ȟ��#����4>%���L3A��0f������t�[~��t`�s9�J�'*��ύ�V־�B�D�&H�D�0��e-����1��{�=��j�y��'eA#���&ل`�H�+Pn��@��P�ta+�nMv���05�(L2�g/f�r�-���"�����n�w��g�p�Ƚ�
̿�����5������&	�B�gٗ��u���z�H2 ��s����p��u� z&D�2$��u6ڞ_/c�_0g��"D2& ���Gk�~�AiO�x��k�����v��!u�i����3�Zr���=�=6���.,Í�d�d
U�^^��L��M�E�R�np�s6���8�u����3���Q�2���P��xͷr���.�FJd���/Lu��8��Gn�F4�+��{����~�8�q#s��62 �P�d]�V<�q��q�}<Vg��^���_nW|A�A�$��E���W,!̟�x*��IQN��]��,�WS[�E��
��&.v�6��ޯ�� ��S��$A�_A����s=�<�i�u<��C�q�����.������X �#�$�@�"d!�d8�q�x7�/����� ��e,�U@���\A9|��_n�2����H݂=͂dAF��;��#u�͜K��5�u���y���w �/���$���b�쬳�G���`�O����M=���`x�}X�y��%D]�]K�Zʛ=��w|�m�
��z���
�Z?�E��z��qK���3�j3���\�h[鰔��^Gv_k�E�s+�����s�$��}"dM����3����1^f����uN/g�OT�x�z: ����Y$w}�}�s�)��Zk����Xj\�Tk�I�]��N����L��-t�b&kbb{>F[��A�3�H~�A:�!/ݧ�����ǯ�Q�Tn��wp����ߤ��weQw$�v�@��dc<���^�o���.�ϞOf�k�ՎW���}�� ��_۴�d|�3:�P����������%
��­�S^�[�v��E�3�*H�A�|A�2&A��#a;9�u�r����(��db�rx׻:������np`�}H�͗Nr��"L0[F�g�]�����0dL�d��?H��M��Y������B�z㞹��[��lgx	�A�����D�!ǽݻ��.t�����e��b�o���5���#1pr#5�g���?_�e=�-����Y���j�:�p�����9ڸw�j%	�Y�I�
�%�D{����Պ�f��i�ܹ�.���y�r\�l�κ�	]���<�hG�����Xfj]�n�j���68ۂ�y�@�ڤ��g�k���:���;hb�r��qvݶJ���v��`U	T^�q[e�Eb�+��1�&��M̯Tϖp��6��k�����N�;�q>=��A�l�zr�4ϯ� ���n�³[��܉i�w��6����0v�f������io�~~a�$�_b�g(+�o�/T�x�(�]}�}t�z o���A �#`����=����n��JV�rR �ξ�����e�ǯy�y2��ۖ�C�i��O�O���GDH� ȟ�d�ۇ�<�q����n#}�k\�!s�͠̌3�HwP@��橈��-�RSqFMu�7�`�߶s$��x����@�qx��;Ֆ ;��>�:���DF(�==�!X����og��]�r��?�)r ����n�o�U��>oo��6~}���+�r����½a�<Wk��l؋�&a�+LgR�W�̡��w��a�ц�3���	�����q�ʘ���b�#�s��:� �oP�g��F�dO�6�������,���`��S�������ٱg��mA�譤�u������evX�T$Z�^鮇�w���i�x�&���<璓���<�5~�ʁ���d�6/��: ���v�ݣyd`F�/�X_l��;��v�������e���G&J�'ݣ�uY�v7{��F�I����}v�f/� �k��zR?n��w��Ύ���R�9}6�#8_�ku�w�	WӦu�y0A�F(ȟ��dI=֣�u��t��y��@^T�>���F�'2K�� �������k��xup6ՠX��]T%�Ĩb�׈1y.q�iF@��;�m�ַ\dK����|~k�@?t�@Ș"D������xuY��^��c;��C���� ��|D�3"g�#�=��2�O���PFu";ڟ�7�9�]{^�M�'%7��wi��Vtm����ܺ)^D�w$���&rq�l�G2����h4�3i��W\�߯�M�*o|��AΚD�M����Z�Z�o8��݁[�]G_�gS9]�{���m��5n�cr��˿��G~@�tK��Χ�7Z��2}��p+��8r噂��M6��ixF�OD'���,�%��TCw����oi��Y����r���u*�����G0<2�A�i�[5j�J����meVk��d.\���$�U�YMb=�9]�j��w3Fou����̍^	�j�S��M��w�h�5����e�|KJeT�M��yu��So6���ut��/�6���
�*���2�Uǚ��V-r��u���R�<f9Ki�f�\�U�Y�j�� �M�dn��i��#�ţ7��N�D�n���q#���0�&�b�t��J�����h���������]SF��ܙ��X��s��xp�I��Ivb'�v�=�e��c�r��ٷ��tE��uoK��È�[2�-�w����ofER�z�r�J�)�Y��,�̗*�u	k4]Ŋ�^�ȭ�|Wy�o�Dp��7��VuM���y�\�Ò�bN�uś�q�yQt�#��-�5³�#���$�,��N
�0�p��8�
T��AyOp�2�nʽ��r�����2�� ���\��ycT�� �
�{�7�!�m_@�+{����	��st���)B��]��t%?2<kِ���ݹ��P�"t�i����b�����IԻM�r��e�ށ�{�;y�}����7:���\�(U����\n�9v3u��z]������(�*��r�v���I,H�:�wffcl���gwZ�4F�4F��)�(���H��&JXfI-&���SAhƌjJ.�W�v���!"�(�f�r��$Q  �$%��ȍH�nW0��L!DH�%D�4b��(�22�c"�#�2!�&��ↄ��)Ca��dhѥ�P��"k�qw\�))��1�!1�hEN�c�]�ɤ4(�S&%e$��RƊ��Ȉ���@2�L�"bRE��B��4�]w\�C\�D� cFG�����/�����$�rE��~W��0dL�$I�Y{�y]��r��`�*� {��!ڭ�A8OY��^7�����Ko+7�����;�0d_0d���.<��{���/�%�N���g�Y��R��o �t�(#��4�}U������a��o
@�rD�V�.�;v�`.���x�6ؠi"Q&�S��/���"7e
�DG���\k�/�x�V[;R����Ǿ���g�2	�:"F ȃ#z��&Uٽs0h=��=�?��[g٢��lI�?�D5�4߮_�w���w��C��L��Έ��?���G������p���r>M�� � � ��Q�0D�0D����vQ^�Ù�� �܂#�������;����{b�!l�� ���#Y8O\��(���f{8�"���v�i%bn����Z��]�:�����B�<�o�U��v�w[�oT˦r3��-�	� oɂ�g:"F?dn��v��|�.�lN�/Y��ʮ%���ؓx;��� Fۨ9������'� Q�He �a��L��h\̲Ѻ���4���Ҏ���Cc5�o���,�?}T�Ⱦ#��=����n��M���<y�3������H~��JD�"X����<j
!�o�����:�.��Q�+�'=���0ț�v�]�{��U���`�r�%
2/����H��87U�N�́xzɛ�ѱ�8�r��5F���A|dL��mm=�o���{���� ����6�����#�n�J��@���7r�ᜍ�ԩ.oS�2$�_H�bFM}�T�.4��B�퓪��x|6x2�j�����D��D���;AV���|�s˭��
*�����"�A�˼���1J8g��I�UIR>0<z3]{��dA�nY�7dV#�^8�1)�c�:�A�4�������)���
&�c�c����1�=��σc۰��B����^�9����Gs�N-�b�!6t�O羾{|������ɹ���y�1��vx�v�䚕3LH3Wh(��gE.��d�%�,%+�Yk�j�G=Yi6h�-be�R�9m��f�i�{c�����wmXx-Cm��R��cWkk�s������ʲ�lz�km�;=M�i�����ݱ5k��Y\����s�ڃ�P�dO�$A����a�>̎6$�=N��5�[��9����v�2'� �$t�+D�S����u_��R߈ �jpm�����E�dEP���A�n���.kXˡdL��)�0D�����1�#7h����V�7��S�x�ߝF���"
y���!��y}�F9xo;�ޣ�/.(ؓ80~;����������>#���#���E�H���'��;>|O�m����������8u��I�9�Π�"��ݤ;�5��fo�%���W��%M�MF��]���n�:3h�l&H4݌U6~I
i$ݎ�����W�(x��o㺂>�H��hv��zW6��{=�0]�y�A�w��	�:"F ȃ�����aG��by���ޝ��KsA̕}9D+��ZC+������{F�Jwkqf$2�����Y�o�;ޕ����̕��e"E���oQbM�}T;��|f���a�$��4-�D��sa����Έ20��22Gw��o��31�x{x.�T.p@��_J�2�0ȒU�f�a�{�B�a�F�v�^����s�F�Ҿ�s�0C*fT�EZ�8�R��{�dH�ȃ �$�FE�}��{�^�·�Fl�Y�tt�o�(����r�d@n���CBd���YgZm0�RtY�f9�w�X�����.�
��vɢ�r�ڠuqף��H������d����Onw"���b�j'�!����a��@������a��ݤE��m�,��V�����_lA�d��ĭC�}92��x����@w�`ȵw��=]��_7����r����"`��oo���\i�T���fl���n�.��p��u��ϑ��̖/��bdJWvџ[ַ�޽w��k�P��;N�E{7GR�ɪ�O%Y�آbL��r� ��F��?���~��ě���׳��6��h#җ���O��}{7<��32J5B� A�@/vPۿ'��=��!dI�d�A�A����y����4����.i��ɕ�����Έ�A�dL�$m�m��a؁�h��e�,�A�%Uv5-F<���D�qH�ja]JM����˲g�|���Fɑ�|���.�n���%��LI�ԧu+O�'�Q]m�@A�<�gu
���2&AH�ӫ\v0���&�3��ɹ�wfd�j���"��ݥ���"�g<�F^ ��_n����cu
���w�v�o_:S�=ܙy|�'o����Ⱦ`�$`!=خ��o�ʞP��c��ݠ������*�OH�1&pnR+��މ0�V�zť[���L�ˏV��r����5��.Yа�Y�	\ԥ��ӷF�`��N�j��̝�6��j��pm�E�s�#w�+�=`ș#��a�d]*��x���<��pd��}�yl�E!���j��P�dL�#b���=�����O�T�5�dف��ˢ��%�{s ���X�ZK5��}�gY~��#��a�M�+��G���e���!z��9�-�d���7�3�O�	�:"F ȃJ���N�Mnw��������л:�="�Ě��@��.��1ˮL�Rڃ�čfl�.�]��#��՟N�%����'s)�`�� ��P����#H�(;���ʧe���=_��?�h/���49����R*���@9�L��ު&�h�}��nU��;�	��);��@���7��d��+��鴮�F1:1�10A�2$�+��>{9�PS�U�,^1R�g����I[�����3�ٛq��\�"�������1�)�r��1��o��1����j#�g���=��	�p��"�������km����%��ص��N[T���^e]=��%1����w\u��;g�q6�=�8�tu�Bqv��:c���U�fڢ�Qklx�#$�l]rܜ��h�ѷ\ר�]��t��`ԃ��7C;�r�Hᴄ���j|lY��9n-hv@�ۥ��d!��jf�����Y���	AB��ϟe��/��K.K��1uv�
\X�E�<�0Z�F����#G&k�|,�Ͽ]e����L���o��'��'s)����g^n�zޤ!;�Wǹ2�0D��	ݤ���{�E�߷��u}�+!�Oc�L�U��~9�LFDݡLV�V�g�F(B�Wݖ&u I(P2&21�=�<��nn���J~�r#�x�� �A F�u�d_^Y����UY������#���unO�t�Z<'9R�p�y��&��8i��bsI���2�2$�r��^�;�hy}�PG7���>�;K�^L^ ��: ����}`��3��q[�j؇Ϝ�J���FKv��x�$���=��R���P��t)|�!�B-`��A�vz��n���g{�b~��#�y��^�#��]9]-}c��_#�E��d��	(�T�2��Y��,]�}m2���fF]L��F�]h���dj>x���*Z�c�jn�I�+=CjbA�'u�z�R�n,�c��D$Ld�޸�'��zs-�x���#$b�2*��k�Q���� ȒP��1���a_*��;���<�>9].�W����}��2/�2G���[�pVWxzz�#r?���1/�7T������l�`��"��&\��=�_p�a�dLL���H�2$&�y�/0�k��*��7��:s-�0~9�2IB����20�ѐ�,;�m�D��h��rݬL�nQѮ��qn+�Ͷhu:͋�[p�bj2����	�HȂn�����1J�;��WOR*����R���L����㚘 ����0N���^�K��or|,�_~�A���Ž�=�":�ȇ|v�~��#wu���'`X�a�k� ���R0��0 �{��z�Կ7�#�|��y��Zأ� �hf,���>�x�Vhb��W2����=L������{���t�yv�^������x͏���h��$��6#t���`�����"d#M�ݨ�훫^��A�A60�;� zf%W��U�Ԋ���A�rd7�ڗW�zw۸�yy�2	Ώ��dA�$H���5���!��#w\���{���2Du����u��n�㺇,�?}���|�B��Ҹ��G].���6f#���9ٝ����H:�۬.��z����#��|�;��ɇ��'���A#7���Ė�w�4�;�B�3ɂ�?��U��DZ���<&�G�,/��_n��LĪc6�3��*�W|A �|��a��V���_�|GF �F,�@����;�w6�g+���מ�H�s$GX�8?���<F��� wk���S�^%�i�Gr�{����WCRl1"/8/�("��T��!Y<��OX=׮j�{	O��׏�[:w�*�[��iJ�[�J>�)�Ȱ���]�0T�v�Î��/^��Vd+�,e��C�K;pH2���n�s�ӷ/��r�w�j�U�*����������E��$n��ͦ�}X��IۤK�Ǒ��5���ϞBf��u�`z�[\lQ�$6�j��z	�PL��ڲۨ ������v]ܒ���pc},���~��Z���#�W����L��+Ă���V�@���f���͎��Rl1"39}.�\��v���P�։m��i�Če܅��⻒��]���j:��J�%���ܙlA"d$tD�c�Ci���J��J�z�wPO[������w$�ld��n�C��gE(��(w����� A�F�]��g՝�}��}3El�ʳ�Rl1"382�.k�D�}���:��u�h�U�3uaܼ���85�{�1��I��iQ��Y:��ƞ��g|¡�k��0ڛ�{Z8�׶/"��y�c�m���Oj��Æ����.�C+X��w��9S���V����;/OP��F�x+�cR���g��x�~ʺ��K�tUU?bax�s����*Vr���c��x��{�P,W�坜nf�a�۪��;#��6ݣ0 �#=�/7B�Y�~c=�[x��uA.�c�z�8��ơ����*��C�N]8c���$�hC&����*��s�*����:�a�>��n<�Úݗ&❒�:���_VS�S�Vjy�*�m��\��@S���2�*�#�|�fү�کVE�k/�)���`t-3�U��ko���"Ŋ�1��{X���-*Y%E����rǤ^�I�ʇ�=#c�^�9rdH�#1r����av�����{U��a���9N���%_=�ߘ�Oi����{f�^T�1݂��9��F��n-P�l�1{Dj�� ��j8���ٵ�e����y�z�^i��y,�3p�|sSe�:%y����Jk%�L��I4Y�(�סEr���	P�`9�S�Es����s��*ҹ��p�R���hT:��C���	W�x.�b�Q�Co�.���\�u��U#RUm�\X�*�J�mi����{ιH��i&��;��/�� �; Oe^uu����A�i�|��`�����Ѽ�W���)��}g6��=G��u�Msh�3���C��:��(̪��>���ꕽ���a��0�{҅ݪ��$	 ��14A"�0G�re$��	2fI	4bR̂)#$�wWd���R�� �@��I
 �$�QC�BY@a (&̤)�$E
sn1�ef�  hH!��PX�L���
bE�3("�Jc �Ɉ�9t�� h���$��)"i1#0E"$.�	��0�$ĩS�)�d�(��v�#I��!fF"���`R"`�F�L��!D�0D�E��t˜��AF�(Ȑ��1M"Hf̆�hL������ �1%)�� ���2RfIF��e0���d�!��D��34��8�<qߟ����;�������t�Q݇���=��pGM�ˑ�f�XX�h.���`���`:@���'B�ը�=r��ɸޡeu��0m���R��Cn���!X9��pq�u�l�,�/c=��+�
���y�����=m�]:����lx���ۭ����d�I�������7^J�m�+ט݇Ǌs��b�WS��^|Q�>-N���i8tcKӐ����f{DB��Y�۫�����P"%K�1n���m4�
zz���u%뮒��g��Il������Y:�i���MM�HZ��
D L��!�jۓ��6����\9i��0ؚQ�j'����aM��-�݃�J�p�g{=Jr1�hz��9��4�q���l�:��3*;J�͋Ќ��-	.�+Ψȸ��Q����[Eո87a��a�q��q��;��l)D�!�h�إ��ŲXeL�v����+k���]X�B9&!��l]�\��m,�FdN��j���#Ɣ%��K�ai���]s��決��qm�n�p�j!�V$���X�ܜ��Ӻ< � ��c9�a��>sQ�k];%�\Pv�q��N���>w���;���9�:�{;z��)�3�۳x���C����׭��L�M/0�kh�Y��Z�6��sw�#۲����]�k�:F:�W���k[�\T*���Z=�;�t����<$�9Gi-�)O[v�nݬ&��Hg�rZ !�5��7WA����*0�fV�#���t�����.٢��
�n���y���%bFTz�Ѯ��p$��r6ln�f�m�N۲�tF��	��dȑ�r��,X���}�!K�Bt�[%�s�]�����m�vp+'J����eT��F%n�ڎ����������zւ&�w�u�ܗE-����b�u=�z����0��������m kv%���݀��b����x���*����,#���0�[)R�և���8۵[���誽� �m�7g��!��:�j�
1�n��i��7>;a�\4W8����#�����l[¢���Mv6ؽ�Z�8Y�6�ug���0��\�7h��UE���BB��%�����^#��N�%㨱u�����42�66�u݈��k)�.ɠo�����YD�m)���-���U[x�ƨ��]rOnc��K����	�f_���/�Y{� ���n��9f�AX����PK�+��z^_q��R�S�G�d��$0L�2����7k=��u�;�A�}���w$��2D;㸾��'x���+P�@W��2	��DfD�#�"��C���L䳄Rl1"38 @2��a�"d`I2�����w��.��=l"&���7К�l��AW�W�{�>���׷�����&N_n�@���$�@�b�!U�ܪ���výo�t�,��IG�\�0N�"3�"$�_�a�}m�1,I|PB���RZq��Hf�F�����t�.��ݬX��G{�>�ǷS�;����c3��݉g��bDfr^�]��W%u�A�ދ�$@I2�2&Bae�p�tcz�~���<ص�w6p�ӥd��7��ŋ�5Y�b�,�/C����fes���N�7xd����_�A��p��cp�_p���ro��>��Q5s�� ���D�0̊�ށ�cG o���/[�|���$�@Ș ���뗣r���U^�=F_d�F�gw��L���0ȒU|D���B�\�`���_s��0��L��Vg#w�)g�l�����A�t{��U]�Y�!�0A��$b��0D�������y������՛�Յu8��j�/��胼�2& �v�{^���+O>�m�٠���.�C�Qr�p�7�����R�"�ml��䞟l�����|�����PA�w};ݎ�{�l%1�pc�sW���o��X;���D2&㻩�G'8߰8�����''�ȷgB��Y7e*#3�&e> �s_۵��pət;\�~��y+��&A���P�fg��4�r˔��:��I�Y{���W�B9B����Xw��o�5D�*u�띕K),;{}���:�Y����?fc	�x��{ד�V*�W{K2YP,[ǂ����������3���0�ۓ����7y
"�1Fz� ���[����/W��a4�l�&b`���
ʼZ�v��"gW���a��#�$A���[g^V!y�@z�g~�Iɢ7<�=����	G=��ba�JlÁ�H��C0,\��㣌��7��%�F��]���A�����K:�L�:0�J��FƷk�б{��F��^v�;���먳��a�{�?I#��
�Z��a��T�Y���d��2�=���-�͜��'z�3��,$�ΐ�*yyџ`���+�����F�|�2G���G���j��~�l���`�ڀc:P�"`da�$�;ɣ<>i�A�{�+�#c[��n4;��F�N@es�#<����W�CD['��_,\�+J����F�* ����Ss��)#��pZW�K��Z���~��*�8������H�DI(P2$k*�u0�(�M˼�w�6���8�c�z�3�����V{$3���yv�e���`�͛���u�\��l���rX�9y�C%�KuH������@辑$s���F�l�ͤ7<�ԣ��*��&F+㼘 ��I�dO�8F���_wP����ڡ�AU������s�F�ql���D�a��艬?�@9%
�Ⱦr0�v�{}2����u}'�t�
�bd�$�_#Ș#rK�L���?���0z'��H��R���*f�Ī�_	�@_w�������9���,$�_H��Dhl/�L1q�����w�JKFN^�:��|��<��j�K��2�{=/q6ѓc�fо�=�:6�;�T�G���Q�PUY�V��]Q{��=7�{g���5�a���ÊQ��]��g�j�޸	L��Z6������v�I����ˮ�ɹ97Cv�k*�c�=���֒�ۇ�vx��`[���ó�B�44����-�c�M�ki.�Es�]�R�Z����]�q��7��*M�nIs���y����M̝:�i���61�X�|�9���v�vA�S	ں�#����ʌ&v%��	t�
CV&�kZ��� ������hЦ��uIz���f�釞j�g/C�i�f0೦h0K,��u`� Oz� ���;�������_;���V	��v���˳��=_W�F�ș�H�I���u;U���~�|6���+��I'4����ڃ�B�DΆ�qz�t�"��_P'�0A���J�1����~������H����;~u�y���A�:H�����ͻ��å�$�z�ɂ��w��}�꽧w�GGo1�10ExL;k�������@W�tH��	�:fEb�f��lw�v'����ޕ]�dݕCo�����B�2&21��Ö_�~Os�|�t�����&vc�	��'�t븂��i�X�蟩���	SZǏj��<�I�PC5]x����C�\����,9N]8=�?�r`A�:"F� Ȁ�A�����	��x%�W�L��Kn�չK�[���w��uV���Tw�/�1x�0�u���B���h�Qw�	�e�9Y�3�Ӑ��{���\�w�GFw{�1?�;�"I9=�ݣï����9����H��Y�MM��r=���s����UL+&l�*�{��ڃ�(Q�|�`I�Ĭa�^�ҀoXdI*����mw�}�HX�+� ���=[/��r;�VO��A>���"�AJ�z��S|�X��19��=�w��#�;��m����#wW�n�w�U���D!�O��P�6e�������]{�b�"� ]���u����U6�LJA�|F��b�� �gx��l\�L�PU�!o�7�9;�|�F5����)��F]�P�w�^_+��w�^vЀ�-��y�Á�������b�W|A.�2DݯV�fU<�ne��_nг%A��2&�
�8nKswٗYw[^w����bhj��ӷ4fU�cA!�wԂ��VO�y���n��&xr��s7{�W��
�:L�Aә�[���S�z�vqۉ��ѝ�3 ��I��20�2/���0j�ѽ#�$_tW�${�̞�=X��g.	�<{P`�A�-u�v#K���Ȝ���#dLD�?��t��*��4/{��ܷF�~�0x���A��� �0̉�	�:��Nw�����v��lF���;�-�2L5#���.f���C[�n�׮���|�����|dL�$a����w���{&��l�8��ךsz��exG���+�# �#�!~T��SF�=����&��Fw7�NwY~�Co����A�$b�2,ګ哶Pߪ�dU�D�?H�"I_
����Y�W�k�o�`�(K@�����������&H�<��GϚ��(P3���#�[�����ރ��s����Oخ�L_��Џ���+|�:��-ͫ�E˘������\�C&1J�j�(�=�ifo��n�O�:R��ʇ`���^��D� �d��2?�Z�F|'�<ߜח�f�.���t������ ͔("D6����9��U⎆�e&�L�&�
�֗�X�{����v���xf��hݨ�i�������h耒`�:=�����;9�}�1%�U*��"��w� �#�D��dA�G+J׻Ŷ���_?��Y̽��Cq���9���(1|��0Ȓ#[�-���5��3����@�$a� ����Mk1W���K������lpR~{Pd���` �#I����hG���m|Č0GoU|~������V���:�������r`�,mסYJ�݆�}ظ~;��#`�dA����[�E��(g����Wno{ޖ�U{�d���҆��%����+�:����;51L�J�+��dK�����Wٙ53�ZnCk��ڛK҇�U�G��A����8'���}��t��Ab�ܼ�������,o����qh�$��u��-�.������(��e�6Qi�G:WQ�0�.^N��=����[�}��E/n:��,��,�[)M[x�G���\)��ٍ]��i��	S�d�4S@-���u#�R�6B�W���;m�Z�+\���m�*ص�n*>��ѻ�Kl@����ΝɱD�a9�0T�<�g��!͎�C7cgQ���_!��:�1��k�$D&�n����v�qB[��d�j�l\�_��^�|u�}#����?$u�I�W����N�	���^W0�ƭ 4]���`H��`��O���˸�<�T������L��*�s�������0A_ھ��Ҿ��7X`�y> �(Q�?�"F<��
N�`����'��~ɢ#�L���/�#|���%
��fD��h̻��]�Y��W���J@�wu>ۯoN|��͎
��ྙA�ǖE�=}��wU�`�<�I*�2&20�"Hs�ԭ��A�0�G�෯G��|�N@v[�"�Ș���|��Ν�I�U�0~z�ǀe�yJ�x��T@ie����a%����/�}|�� -�B����
�m����M�61NQ���o���	�o㺂;��#�Fׯկ��9�V2|6���	�9oM��7�#��[���|q��y�z&�з6�M�?+�w��x�+3_��k����jR��1�j&���W��>~w���P�r�2�Y����Ћ�����7%z��"n� y?��D������o��{:�{
�[��|��z��W�d��~9�t؃ Ș �6:H�p�1�%~�Eo���u"�z�w�ݝG�̆#�\�	ۉL��g�{{��ݠ�唷`�;���#��"G��v���{�fb��y���\��U�3( A���v�[^�Nzҳ�-}+]
�a�COt����b����.��q�5qMu�̥҄�aen��|��>�� ��0�U}"k�������_5�/oݼ��WOH#5�dLL��"F `�����o�`��$A��Ν�5���<Ύ���	�� �7�`�%T��/��~Q�2	��$a�"d���ͩ�Y����uv��]�]U��VK?9��V���(�ٗ&J�z{�b��Y��������I�X�,l1�B�*M��CpW�s����U/+�V��(�^�V�1us�u��ΛyJ�aB����D֊�y�G�D������wH�f�固~;+�u[��Q�Ӫ������wwۓ�}��=���UW�>C���qA[U�or5�^�WG����t���m�K�vi��ٻ�I5�����UOy�l�NC��$^�͞�5��)�ka�S2	v�yk9/|�.�Se۳ {
������3Y�����hE.��-�3(Z�%|�c)�5�&�U8��h����K��m��ڶ�X\j��v���a�jWw���M�{T����L���|M������F�_�e�cFKMcķ�Su&�ڒ��{O���y���Ĕ��#��0T�f�ɔԛ�H�&� �<�ҏf�Zغ΂>�&���x��|ws(�u�y�n.��teՠ��v�W/o4��e0� ����lvU߾w�t��C�w�5��b������x֜u=ڧk+N��.:ÙWϪ(��h3�^�UC:��{��i�۞�sZ6��>G5�%d;ϪF�fvfu���x*�f�鸴�%)�]�B�+rݤ�e�V�V��ngb�x*��i��5�<[��YwGA�#�ʾ7�zu3Gv�V��/��]ޚR��Q�7"���k^�]า�̎�\����y�u~)��C+/�ƽ4���o05c3�U��2��_y+~l�I9�`�vq��űt�w0�J��ٮ���[o��.�/��(AL�X"P�ۑ1\�H�0�"C&H�I����I����ɦ��A�qH�� �	��!1($Į�B�"1�!����f�)d�4���%�RB0�I �t�D�1���(�IH�F%2R2)��$�ᄤ3��Be&�I#`��D$L�!N]fL�0i�K,V&��i&��$�4B�K)2JF2E �$��0h� *D�� �ݹ�IDȔ�&T�d���q(̋(ɐ�"�LRHI	RIHI��� �h�#"DbFARe,n;�	�t4b���,EL�,�d��i�wm�A�H�$54̑�Hл���+�\��&�i���������'"�UY��'<	�|��A�%
2&A0���ǜ5��}��^P@��_1����f*W:�9����q�}i�U:�s�� ��>��'�:"G��d@1$�Gv��f���m�\ۜxc���QvW~��쒙wtReܫ��������t�k4��&�b*fX�Q�v�]��<ppt�\8{A�_I��[��Iױ(A�͎�|��_�~2Gꊧ��U]���XhrM�RC�k����$a�$�@��Jו9�f�^��e�W�{�}�gko=���7{���u���G�t�t����{�?�2J��A��c�	p�Ov��ӳ��ʻ���&s�1|��0D�B�"F2&B����"{)?y8� 堌�Dwu?���gn�վ��Co�ڀ�/n�pC�ZGc���Mn�۱j��N��2�d5�V��}EA����Bw�Mz�M���(�G����J��#u�c�1�=�V?^j{W� �J�Dȑ$���z���|�=R�bJ��s��Kٵ�w�@��0d_0�٭���j�r�l�dڗ{
[m�u����Z����ţ�s�n]��kv@������� �s���u��ٝ\V]��GD��1[�Dʏ2����B��#��W�/�W��$u���ı����<��,���:����T~`�ڃ ���q��kqs��l27q��`��2$�+�����X[�����so����b���@���22GDH�b�u��.C/|�U ��b����f��'o��9��3�^����s���@����X�/���d��"F�E���+r�w���/?e�g��[��o*	� ��A�+�$Cً�m{M�\��yVb���ʷ&��D;;ު�h&�Ɠc����2 �N;/Z; ~�<~ǣ�ZNt4�۲���]y�z���C��O��Zͭ��p�7\�`M�/�(86^����y�] t�u�1����ږ��Q��!�q[�4��+���Q�֏��
��q�m����h:d_oX���5��F ۣKۢ�vD9z�M����%���p��IF��O��Iu��nwQ�8�I�N�Z��`������\0��d���n���AN3'D(�&ہ���ϯ�,?D���ld���L�]�;ۂ�����YT2���QL�4�h��E��AȾ}&���+/f+�u���mF��\Dn��]+��aߕfF�����wS#u A�@:$�-E�w�CG��0A�����7�˃9��3dm�F���o����W�/Xf�2>�tA���|��44���}�6�uyg��[���P��y�%1�]�I�ı�rK.�>4��}��w+Գ�A�td�1�f���cɷ�u�;ȼA�������{�=����3c�Ld@9%
2'�>Sk-�����훜�"�,n�tK����H����纇C%�nq�����_*�ZX;�I���9�6�h`���і��݉���&u�	�r�|;�]玖^����~� ��O�7���Uy��Xc����vdX�B|A�e
 �/��0D��"dE���ɿn?R���k*�YԵ��-t�4�w�Ӧ�Q�V��o=����x6��Y���#����YO*�A��Q�f��.�۵��<��x����sPR�ve\�W��N(ׯk� �o����dPP߯^��t��?�2�J��$_t�QK�l�\͝܆q0N�<f'�#�$�_#ș�G(뛷�v����NA��6<��vN�mN��4/� ܠ���ז���E��A��"IB� Ș ��n�z؝�~=� -��]��3��Q�n�	��7�`ȟ����6F���������QJ�VX�%;5�=���&�������N���,��eׁ���nsșF5~��z�F��C8�&w�v���7z�1�$�s.�5w*�>M]ܨ~��O�f���=� ������:��;V��P�����{%
2*���{<o��^��*��&D�2$�_#^��� ޜ'W]ĭ��9�L8�oM��l��}ɻe������;ՙo�-�TR׏um�f���(�
����wbûɘ����bZ���^}z�F���$u�!Hா'���(W�rdH���vw��hn�3��\�;t�?Z�3�ˉ_w{�cHw��v0��0AH�"�"U�\�v�S�v0�i�+&��:��>׆0h_�/�Pd3e}"��9���+�]��>����_�Ѡ\5��k��d�ca�(FArZ�C]��AЙ�	�RĘ�%��ɥ�σ,���<�P��A�_wns^�ݯ(�'y��m���s�/nMQ�{�`D�?$H�� D]~xF�:�^�N^���a�W�$�|�C2��'D���ۤ9D�ӷ�ͱ滕��W�1��9ɟ��纂v���9�&?	��{�(�����ߘ'� �I_H��dI*�Y�Bz��A2�ߑ�H� �����a�ڦOdk����iJWy\>?_�26�3Dx����,d:Ve�|�%���ٛ�-[��;���:�R�U��Ln��dHs2�Ӕ��]tt���ӥ�M-�kH����9�H�?`�$�(�3��-x�U�U��wd�<���pK���#ݒD˻��.�8�ߞU�y�Y��ń�M-X1�+(����˓x+�ʇA�M�P$UH�ꚤ�/�d�� �fD�'wSy8�oo����!�J^�OL��D�Gy?�FJ��2'�m^��&&��@��P�0��2{#]�|���w��}i�AȂ���x��l�ӳ�J&Fu�AFj� ��;��z����K�̑��{2/�ݡ�|�Lk�$���R��S��G���A���;��ãȘ �#y�:����So
���w�2�<�*Ե��O��_=�"IB��|���D���������?.�g;��򫴩Ko�����o0��3���܂���s�.x�ŉe�̺�*����鯽[v:MV]�v�d��y7v���i�D���{<��5�5����~�e�Y���1wh$�V��T�@v�X�ڞ�%p�糇;�;�s���n��X����&z�I��X�`�@D@{`�>d����9vrx��P��ٱ=�l\O�(�⚶�t�ΝGW9����:j,nvP�N��ƞ}�AH:ո����9G�9�^:��ūI�+	L���:��d1/gbKKu6�y6W�����aJݠNy��k�������D3!5�vŏ61Ita��v�#C��@1��( �f�zt�7Cs8�'Gv�P��l&�;W�3����0��2�H�1���_�	/�� ?{��V��g���B��6�ݨ2�f�
2-����ф0�Y�_H�bF�I*�?H���j#==�%9=�W~�KоO�W� �r�胼�2&A �$_ji��E*�`���C  ��a�{k������2qi��Ӱ�s��_x��C��Cٺ8s[��?�V #�A0̈=7�Q�URa�_i�p���hAC}�����(PD� ����6���=�+)hI%��l�4��wGm�,�Km�K�0�R�b']��&�ӱ�ӑ2: 6L�����9������a�J^W�Ŏ�n��񾭘���_N�����$��d��l��{�Tذ���٢��N��~�%�7���޵e��h�+u�C�̓۽Do��*=��2�g �k�j���\��|�㽩�� }wrn@�1���'�p`��� ���I2n�zz�"/7�����0AF�J@��/��&NU��l�P.�;j�7��0L�M�0�2�D��󨭮S����A�A3���2Fg0���s�k�ԥ/+� ���i���۽Q��7��?ؙF�J��0̑p�{�8�:
��;���5.L]��	�.!�.&;�"&��	#C=~�:((�tj��}������Pn���:�`n�"&�W
��M�տ�D�=��%_�$M��ޢ��5��Q��^x
ۗ!r�T$<@?�цd���"$��d��oeUi�Җyxx���H�[ԧtM�r�*�S�_q���#$IZ�����'QM�CO/�v0Ou ��?��0A�D(=���d�����,�;GB|홲��<�j�7�����؅MD�'D�'J��@��C,�!�:Y�J[���#�یOOm�5�B�^�L��H�~ 8$�`������#$��*�"(Iɴ���O������;�x%��Y�
<�����Nʠ�f���~NA$�?��0D�G7b>�~�ݰ�=6�Ε�R����������rG��dd�t��Ǹf`��ΛT���G�L��	�1f��3�[��bg\�K��_<���A;�d��d_yz�N���c$��1��]B������;��$��*�?I ����ܦmu��g���ɀ����4�y�h�C}|&m?n�2Es�`�U��e[A�����A�DF�HǷ�t^���mefx�~[�ܐ}z��>��d�0���D�D.�r�u���m��A��aH��ٛ�]��c$��9q}C�㚅�
oX���R���]_��o�mo��'��]�#�M�*��8��^6S��a�N�s�Z���7k�
�5��S�+N 3s�d�3% A2E�0�2Wy��w����KL*��ڽ��U�i�Q�����`� �U��,ۣ%�xO�__����X2��:hi\s.�u��
��^g&�������iq?����Ͽ��G���g�uw���+qt�
{+���3)�&Q�洃��3:��+"H�&J�����کL=|� �A�{7{�@�nX�F��	ˉ���$�/=����R?gD�H� �HL�Kc+-W����IO�Q���Dm�|&m �c�d��$A$�-W{��s���ZG��������`����Zr�WJ�����m0F�)x����ܯ�9�0D���H��(���{l_��޻�y#����o�`>\.�2��Uܓ䐐�%���֭����Z���mmj�v��ն�j�Z��ꭵ�m��kkV���mj���֭��m��[o�V�����!!KRBB�$��	.m�[o��m��[o�mmj�~�kkK� �$����%���$�-��m��PVI��P��@�W��X���y�d�������     p hH
�% ����(�� àh �|O���]�:SM����=�  Zγ� >\ �٠����+�6�$�5W��➀	��ǀB�
`�<}���h ���x��	�xA�`��@    ���
RJ���� 2���IUP       ت�Od�  & ���&L Oh�2R�G�`C 	�р	ODT�ʀ�4 �@  �$�bi�Ѥ�ɠ4���I����>����@��G؊���a�.���>eP2��!TP2������?���y���tDE1�A�\$IZ�PT�����Zg�A|~�>;�"��w�/nO��!��ؓ��P�s�y�@��>?���S��}SsB����Vqڙ��R$�N$s���9��FЏQ�	Ҏ�x�EN'͌5��"�w"�$��'�):v�n�D�(�$&�ۂ�mRA�K�(�e���_	�e·�p@,�]�p81[@��I�V�	�cX�H�Ro@��N#OQd�&D��5���r��v�=wL|7 �Hܦ+��u0i�;&�'8��D��2�82&�Kν�d0R��$E9��'���F�)8��D7�գoUpHPPcFD����0�-�Nb����2�N�k�Lu=���kL�@�勒H2lµf��Յ�˳DU�m��m�v�;"��f��u5�B#`��G����d��C����;(<~�<��㦴��}D<�d�2�r됏���up�k쨋���^��+��c�qJ���H�7q�9D��'Ӹej#�.Lh�2Z��v�A����H�M����.�'_�U�M�^����w��� S������67�;�c�7^���3q�`T��f�*�&i]��GԞ��cL��U����'l�ʻ�J�b��g����׶jD��w\�F�(gqD�Sp��k�a]1���R�U�˦���:`��d���V>���5t2�t�ǆd��LZ��:��N���Y�9e�r�����|��3���I.�T|�.��Fr�ڨ}�����1����A%��`wqs_I�I��熮��x������8��Oe��<@�zjJ�Ҙ�v&2��u��� �8��n��hCf��F��V�5����J�Ӷ-��M��p���A}��������;R�PH�p��G����+}�>W#8yX���{�'����uh�<4���oWL�T�6���K�w�}��փ98W�O�M3���e3�{c�AI7&Bkl�q�|�Z�l�vVVk[��M�d15L�(�@���F�s��,�*���N:_%�~����s�#M�Nqǜ�ې-1������48<� _<��(��(#H@
PЩB�ЂҢ� ��*�J�R����x�]�g�}�~�E��t�:�(!�n2
u��&@Q@�&����m��_tcqC�P�����0�������"��j�&��cN�]D��_7=�.��'�ԛ�s�9G����![ |+\�mD��I��p�V�Z�"�oU~��L�8
s��aY��$qUqu$�-�a�K�e^����<�{�{������Е;X��j
��.��r�/)������/,і��x8W����c�����G� |W���%�6P�����G��]���{�@�;�'�zW�G	j�U9���>ӳ�y�
;)���en�e�Ǖ �?P�4�7E������Tk;\C�͍����4Aw0ӺK'{��
V��P}۳��a����������;������u)�NW{y�~q�ɆX؅{;Y���]�o���۲�c�]�;��w7���-��i=�6��ظ/$���t�W5��}���Z��3���j��K�_��[�[�>�z��Vn�%=�:3L�X�(���Z����k�z䜅�{��y4�O>�S�w��l�[ ���fV�2��ܙZu��a����Wا��_)�o�؈%$yX$'ȟ.̜��<��<�63E�z�/��LiY���A����8�&��Ft��_E>h�a��aDI�� �-f����Z7cb"V�Yѕ�M���*VA������Ym��R�8��nn�ǯ=��{<���QD!���Ӽ�Vs�X}�w�5ޱ�{砅=�}��w
��T֌am��"6˽�:2M1I����^�<���U�z���]�+�Nʟ�~,�5������x�
�!����K�/��C�#N��k�[7�R��3p�50ZC�S���X�S���3�s��ݽ�	e��S�#��^-������%��Gs����չ&G!�k�u��	��ϺC�Z���w�`$)�k�r�4��F�Y� �D'U�`Ԙ۷�F�Q1�ovs9�iB�%���<'">��;[3���&񴟪����/�8['n�Sp1�95�kj�wp�
�mB8:�oΛm�]��;隸���Ν��"(T��`{fa�b��gx�c���6]��f�7m��3;]1���e�|wW&���f%�g�;�Iv]@O�k����q;��5�nM�\\cu�X�e;S��'�܍��'����
ۮk�4�n�N��5����z�t�]�m��n��;Vu���W,ruی��l��٬���Z�nF�3�+��7eM��V�E:y�V�j����k�:F�FU�9p\�ۍ����e���r�-���u-���SA���N�-S�q�]�3땹e�ȷ=��[69�e!�Nx�ngT���&�.\�l&��v^�M�:/㍭R�g�l�ӣO-�i�iM���I{a3mVRvٹ��؁ �C	�#��]&�Y�7W�s�Gv5������n����`�髤,sFT���U7!)�к��Ԯ�����ݹì�����R�������u	ո;8�G6ȇ.M�t��n��~ ��c�\�et&�D�Zl��qEq�՞�����-�4>��-��;iwV�ŉ�-�&���);-ne�*��<�b;'VA��"�ju�p'��umi	V�t�[sr�E���v�V�ӛ�7��`��lUUUUUU*�UUUUUUUUUUUUUUUUUU5MUUUUUUUU)-�:ێ��U]H\���5UM�����9���|q5��m�k���Tau���:eۊӶ���ዖ��uV9�.sڤy�v��"�Gn���.Y�qs[n;a�xvmbP�m��a��M&�Y>��5#���R8D"2!�5��gU��Y�r1�"�H�Q3�9'2OaDP\5-�s&*#��!�ʱ�#E��IY9�:Aq}30���^�/��{c�xϩs�ѫ9ѕ�sֵ����sq��t�4d��͡�<�	�ruWDm'[������|u���ݧ���>Knǈ��:{lZvv:1��;�OB��.:c�WW^�鉩V�����FF�	H2�N��Tݖㆠn��"�;����>v���gg!�^T��?[w.�A�z��z
��B��Ftrf�߶�0�:4��KR�J.�01��uJpB#�U����,�
&:+x�Ҟ� Oz�kB]$nzV��{��W^f���,�9��nsS˴�"	9������W֘p�s� �j�Z|�fnL��$�&����7t|���c�#�z�����ճ�tü��᪥{�+r�1��P�4���;&p�7XK�&h���NSoĥ|fH�\n3�.T�F�C���d�i��E�$��kv�^L´�Aŭ�-Sa��i�_��Ԥ���-L�n#[�8`���L�q �5
&���s������Vy\�3�9N*Lj�3�����2FE�'U뤈����Kǎ-�JԂ��"�nP���r�JNr~f��cGolE	=�{����Ð*�*{���}���^�['(�b�1֝�xؘ\�b�'�!s���n+��^��u2���tȗ����0���z:����&����wv�U�Wl���K`��S�:�n�W�4�;��i����ͷd��vۈJ�g�h��L�Uf�o���|�C��+��гFH�N�n uj��P��2m����-�D5)(o<~Z����S�Ք٭�P���Qtʍ�'oP�	\Ӄ����9�H�p�Ú�<���y�z�x�ᚤ���������6.D5���\ܟ9����8����������E����R�)g{">��N�(|�����G:����^5��_����S;`�U��в��j�45��l�rf��5���>��]zɸ����b��g��*t�`UDQ�$m��fDz\+���`��\��W�Fu�BN�6�`O	��csi���_(�O;ټ:�F}>|�0HRE����B �՗P	��婫�o�D����\}�>��+ꞷ�7g�����?W��j"`���A)QL��rB�}�+���'Ļ�SS�2`L���i�_۾ql��6�vF;O��}j�Gmi�������l��1{5�`�����g���˰��i�H�d�v&Rz`jԄ&!Cug��s@�s���M��#�5���ҀpMk;��#옮�V����eV"��<���,���ʹ���N;�1u36��������0p���'q��HG�"FQ�1�4ƖL��gx������c�2����c�r����J�9�8�UL�i���� ���p:;놻���O�~�<=�������=G��0�ሥM�j�|�����Hi��C�{�\�M�()(�9���a��K���ɴ���`"1��	�G���u�	���^��_KG���cqZ(SJյØ�ѝW%�ĽJUUGeﾯ}L��	�a|4����
���I�y�CX���R묚@�%=u�\����뮺�u$���ɍ����^��z;�w���>�>�wF��m�t�n��N��\)�x�9�羝�T�M�:��CHw�0RR�m���\���!	�P܀(��>\���5(q�ad]Ie7�~���K<gL�G1�[o���`S����

JJ�\T�S���x�"G��a,�����e3$-X���k�e�(q��k��QK�t�}5v"���i�=��;AM&��I𲏀��`�j�VN9�US����s'<�X�/;u[��M��뼥�;��5��Ӯ���K�w��K��0�E��F�ۮ�T�0<M��hi;��CHCY�uu9���˃N[\��LǏn�.ܐ[C��t�3���eď��d==I��Z�54�m��<�ܟi�{����3�ּ���_Hw
S�r���|w�8�-��ʕ������董	?#�y��@�I.�)aē'�1�m�#��,UY2c�T���E�s[ r61!b�K&D[�	�s\\�t�U"DȆ ����@/_s%)�U�mH�[l�n��%�u��<M[�w�m�&�R5�;�	�WbtH��ZN�ڣ'=��;�۰�z���=�݅����X�x6���M��ToZ���<&�vn4��حƬ��UUUUUUKQ5N� Dܸ���򳖘f���>��n�h��\^��*�w&b�D���4�i���)sp�@����N?y6 �1/=i������5�Nڊs��Z�:�;�3	AI�H9�L� ������x[wwl���a��B�>��ѹ��E̺������i���:k�iK���AR���v�u�^�	BP�%	BRBP�%	BS�����|a)
�)9۷mXJ��(J��*��(J��(J�u�m���c:���i!T%	BP�%	BP�%!T%	BP��;u�!)�!(N{g(U	BP�%	N����)
�(J��(J��)c%	BP�%	BP�i� ̅P�%	BP�%	BP�$*�l��%��%	BP�%	HU	BP�%	BP�%	HU	Iv������m�m�}��+����o	BP�%	BP�%	BP�%	BWiBP�%	BPg�z�u��(J��(J]��%	Hw��:BP�%	BP�%	D	�;h*�"P�H�*�^l�BP�%� f�e�%	BP�%	BP�%	BP�%!�81�c���LgCƚo�%	BP�%	BP�%	BP�%	BP�����Ma(J��(c�at��k�H�1�2�%���#ā�����`�eC[NO]��wyG�����RP��:�g~�e{q���|�f�f�����������o���)��R�q�ր�-�@��^�=�$J���xy
�E�.f�X�xg���"�,���$	�*��h��]�	US��p�_���x���hܽ�mZ�N��H�:��iN�5��K@�"��t]����F�ﾉ�^w
���{��(��veC�LQ ��l ���H$!�3ceiv���_/{�M{Ê�3���޿�U���(4�j!U�C�_N��7B$�:"Y����?{����C�Ԕ}�	��	9�"wH0��SVLu�Ѣu!�l��\eX'���b��A
F�Mmj��<�õ�(�U!�� ����V��ۛ�ϔ�I���@�z\���D��RF����#����=������:vlr�4s%W8.յ-t�]�UUKJ�?����#IC�Iԕ��hD��2`���q��i��޷BF_�r!kA�y�m[no�p��S� <��@p�e�|��J���$���oR%�Ό%�����n��s�I�M�O㯍V�[ê!�B��}�ط����N��p2N�BjÁ�ŷ���Cw#�s�q2hKM[T��A�wo�WEV���/��]��wݞ+5��.,��k8�f��ea�"k7q銮�GW4`B��U}6�$�!�"%���GnPJI۹��Q^E�	�R않2F, �Ҏ�y�"�a	a�"�T�r���⨉RH��=᩟�J��?����>4r���;)=�B�m���ƻQ0DBΚ��d���}�߁ ���r��;���?��{͓��7~��,.��
E5@�͘7Pg�Ȣ:��*�s�s׵3W�rEbl��;�Rg4+�=X�1�i�ׄm��2�q����Ayڽ��h�t��M��p�)=χ|�	1
��	��.���|��K�#��$���̒A3k:�.ӛ�p����)�!n�Gme\��GzD?�/lЏ��/�m�H6W.wd��l��S�[r����I���j-�F�=�&A �⍑ ʓ}��AV��Tw�{���g�I6�v�ݺ�%Oԡ�h�މ��RV�j��Ϭ���f�H�+�$u�u���t��S*x�4G�x>/��s�;Bm��QL�s�OճBp���R$��7��%DF��$��	�M֛	���Å��	/�Y7Yx��F{sg�A���UUEY��������9�ð�8�$�ErA1��j�f�t�L�>�z�$P4�`Z��LB����`� ��p���#"������B�$�Ј[ ��S��F;��;����D�P����OE?}�$���Gk u�<]v��c��d�N���s�V����m�(�Ů�|��L�뮂g;ܩ�wt�m`����U�P��Q�*(ڑ�a&�J��m���+��#����,�ԏs�PBhC��9��b�&#1\�T���e�Xh�-\�mܰ���<�G���r^n{��Vt,+�
}�"�4'� �=��:��
�]�\{�c�I��q-��5rg<&_]���A�C��ނo�V��݈-}����T�ȍ�`B6'�f��{�
j��$�ؗ�У��e�j��,ӃZ���=[�+ 1��j�T�^+nY6"A�+�h&�Vf��М"�|�n[JR�J��Ex������qX�q��޴N�rVؗXM4�h]I��[�!E���f���һ\�XA�n��k=����=�M��y,�,!��^�ss����.o"t�&![�R�MUUUUUUR�C��)�6��v�!1�a��L{�^u�v�ٲ�Q.��Qn����œr�UZ���}���}��q�f#JڤZ��ڑ;8�Ol�&ȃ�\��������mH)vΥL�"�j�G;&��۷��p;0�d�#�'�R��P������H$�(npG=���Fgfd�ݙ'dЀ�w)��Nw�W��$Mg}b�_�>T�[��Q�D��J�?(�<F��BI$���ҨY�uݹY��{:����gQ�6>����ĽM�J0�A��Ϲ����hb�!���ɼ�z��2���RE��9V��Wt)0b�P�7��Ը|޺�9��
i�m(M���APj��{8�j�g��\����\��/w�ђv�!=�$��gOT \��N�J0hDAD��d��S�K�.`�l��ꚋ�,���8���.��I���+k,Od��uO��|=]��~�$�/��h��un�����R&w��d�F�W̹��ٖ��x�`-�i��s���Z[�ֽK��� M���s����F��dRTB�����]�����]2�+�!l'�b:;��̪�e=5k�r�6z##s쫨7�O�8ؕ�-���Yɸ\��6ZV�{��X����t��4G�zg'n��r���h�� зwW������S1	�!=�q�p۬N�y�⸸c�-�ڬ�;.w������>�Ϗ���$s{�.����oM-/*Xўw��f��iޑV3>y�td��EՈK�6*�D<88�̿p�FP�#�.{5�;��jG���P�1���-�^�]wwG7r�:�7	�%�b,#�G����}�A��W����`È��t+(ܯ�ۋ�;�9{{>[��9���U`��񋠜DZV+u`��<�H�R�6K��/3���t�bZd�{���M��"x��M�ƾ@�<*��b k�]�l*i�s���oM���	�n�Yzy���ޝڴ��"�/wf]��+�"��M�E�)R:;�H4!�!��k|�u�4zbG����z�Z�����C�+j�)B"ڪ����wb"�H���$���\��������sPvw�r�<ȝ�?x��[�UC��dRTB�o@��b�o�4��׌mNGC�=|��a>ޙ,G���V�{��xJ���d&(0H"$�|*>�5�X��▪�i�vw菾0�:�&��r�'>(�I�����w�{�L�a%�ɜ7zM�i��aT�z��em�%��:e�1�=�9�=H�_oʎ�"�~s�NK�v�����X�J`��� �J���Ni��½��#V���uD���WŨ�ʄ���}S{�\0i8M&a�:�	�Dv�{PD̸�TA �;9;�뜩�7|و��k���`�C'����0�we.踗�X+c�z��&d?0�U��Ċ�Agd�&i<qJ�>{�|��m���m��pnؕ9(Z��qn�KUVj��~;���IQt���]y�\�6���Ω�q�EtP"ySG)e��c��`�%Ԝ���`��qϯ��~91��^���W}-bD�������D�K�Y 滥B��i�H+�Tw{}w����V���6��w'x�e{�r.rllD%���Y=Pnƒ��O�u�i�R��H���U�Y
6"]�ng����|�פ���i��,���r� �������$\��>V	����&^��XH|2�9���w��Jf��i?m�կ�_t�oR+�pxߗw�y�C
Yb��4���דA��gE;�<�V���P]^���/tt�r��\J�l-E5�xK9�2��;u�m���u-*UT#3�S��/B8XEUAp^�3�\'�R9�����rB*��/��x��Z4��Y�1u�[66�����ܻ����{$Z��m�t�n�Νgk���n�g����"�u�����iw��fk���!`�o��fwA���\�+[+�{]�e8��E15UUUUUUST��p�r�v��z��i�����_b���O[6�9�ۍ�kW-�,x�������������:��Y���1�����;����$��&gĹ���[gV�Rb<�Ю�*���r�f;�_�7;�&�����K#�Ac��!^���&���[d��丧�.<c�5���o"\Ͽ�﻽���@��}�آr�~q�Xլ�=n�TNE�WJg#
'9uD�I<��Q��x�Ow��D�l�!,D%
��}q5[�o��9�h�=2}UuDL.�%O���@]�j�B3���+�-g�FҵD�b)cR�[QـC�RUU��-�|�i,-u�燷�f9Ҹ!��q�ad+�bַD��+��tDn�P��vL.�S$��j=����y�I H�Y� ��z~�ڏv4%���(n���Q'�fD��C��3]9�n!�"b�����GE�P�	�����&���\�Ad��^{6�^_���75��h�zGsz�Q�`�^J�F,W��WP;�MJQ�F|z��P�M��^�'+\�
�.��6Fw*4�#q���������2 �Ty#�`�^)�L�Ut^��U��m��;/{��$�jBs���0I����z8� �����T�F9��q.�e2�,���] ������5͕ů���Ƥ�Ԅ���话&�C\i�/Hce�ބ�2Qn��a^��Jy�O;~�*$�J���j$}H�z���+V�>���n�8�������ｫ������-�z2�,�3���qc�/�O�WV�����z/�Ɲ۪�90�E��W��\ر���c�+Y�ͪ�F�T A� ��>�%�
��* ��!�����਩&v���u���)v�9�k���(�H�Y�L�P�M7��U�=��Թ�߶s�ks�i�Sf7>���-���	���MKKEh�ķ��Mۘ�xJ�����̏���#vb�P�_���Bִ��D��ꌑg�hxB�ﺸ�'9���]��+ �� �V`)�
Ai��Tf�]1�Y�
$�m�i�	����K�Cf�����v *�(�2�=/�������Y�z"�BP�㕛���� r�NT�����K3�}��i哏گAͽdm�o{�0Tvl�����'1s�	3�-��I��2�U�����)��#��aB�}�f&`u�I&J-��]ϧ��A1ܘ �N�J2x\�n��l�@����W2���o>��~�쵭��{ꌵB~Q�N�{�[�36�&'ŉ�$b��i3����;.�H�S���b>����Ҳ"�,�P�����^��5-u\<�*���ۿ�7�"L(�W@��k"�T#츚�B�SM"
�[ц���$��FA�w8h�osf�v[����Ka��KQ�Q&W;3�H��"��W6@;d�D%A�Q�j ��n��O �Y7]1�!�ܪn��T�"�qc DG>�Ozj�4��e�b�j�.ť��R��t�3�=��6*^�cf�R��T��T�G%��$�E�7BxĎgfY�	�gRf���
��#w� ���ʇ��]�d&h�O�W<]����/^�q���c�Վ\�>��/=z^蟪���n�:h��^ö�/�c�3y�ϻ(���5�Q��\E��H,Z�q&�1��T�kD�1��Ǌ��\Low ��`��9$X�-뻎� �S�lX1�,�����$V�\$��#�$����]R�y5.1����yJ7qeETM�5G��VH��tG�[2'k�I!��|�ջg��×��=�x�ZtY�����qn��fꭳ���W�9��&��a\U���,��&�؂ɺ�9�<�=q�擲��y5	Zj�������i*(�3�;�q�A'u��7^��{o�~5�W��^�I�աf�X]�UUCB�__�~�8�%����q`�u�L��E*�SAw(!֗q I׽"H�_~�&&!wd��C]mL�?�퉙;K�3�Ï#�r�Р`+N��`����,�Ni�JQe�*�Gc�T2�w�W4�A3�s�0_A"`�D3���p,��b�����R�VcU�r4�+��ÄK��Gl"y�/����co�{I��'�}�2!�I��"��}������i�A�_WL�#L�A�Hl��7*5PN�GB�v�fU�0�ax�
eG�.��=�Z�h��>R��)���<�l[�&a��d���S5P�&��@�0	��}���ը�I�(ny-4�*�U��5M����X^���mv̍#9t�N.P��HV�кD�l|Fl�("��0]�T|��)K�>c(�`�.�����vm�ְ����=W\�\B4[�S�1�gr�Q�!�n�3�\�=+�$����Us�����,I�k�I��P��Q�C�Jyr'+��J�W��`�+-���D-�@#:k	�p/�%S��臺�Qp�糷6�N��j���O����澾w�����O�؈����/��Ń �9+�������y�]�f�2b��4��I!	L��dg�޾�5��0��y�HB�
�2	hl�r�� e�)����&�C}G��B���sz�bD�;��`���eBjE7=�ˊ��r;WEn�L��$ڗUo����s�t��}޹їr��A�o!'�WU��]-X,n����܍[����Y��O�ݞg�q9F�{�6�2����$��<@�Gш��'t�)&@�+��k���/R��.̈�`�fLS����	VI�Qn3"b��\-Qa��!E\z[W�����r�Id�d����'6"3���"PE;>W{�\YO�O��*Em|��=��nP��N�\H�m��v��v�����*�N۴��[���܃7<G������tOb�B2����t����ԝu��僆��6ԯ4�s�[W&�*��7M�����L&ڄ�p�;p�%�P#+i�h����I�*;!��Z+�]H�pi&!��5D���=�Dm�F��țU�a�	�tɓw��Ds{0N���m0k���F��򏉅�
d�ڑ,ګc:{"`�r$Cy+AɄN�N�z�� ��Q	�P�x��qA��v� ����H���J�f��>��O��V�&����W�-�S�$|��n�W����O�#��hW�����(r�@�k^�P%��Ubiz\�cT�!�`�wn*����#AŷLb�ܨm��i�=�-N�G�뵫�B����d����P)���O��щ�ƙ��P�)��d��a�9[1��M����J'��� �]�L��r��oW��m�l��F�c9�I�A͡YHO���{��\���rzf^�'r��ej#{S'OP�2�&
���0�/MY ���5-M�T@2��n��3��'��x�<���GEX�I��������tε�D��Ċ0{���m�!��9k�/�_"��|�O�_�!�6۪��@̓��E��.Q0PO���>�<�@��o,�����)��x��S���"(���a:Hs�X���W@�0�����""���a+��<�o��;xm���d��ې���d�_>��ЄA�W�����v�2m�j�<�C��ѫ���oʢ(�}�i�O����������	yE�'�H�ar}'o������}��j�Z���v�OG�=������DP7�@������*�;|��=q�62���ߡu[���0�i��=y�`���>�#�5o��NCP���C�'��"(\ɧǆ��.�Q@����4D�-j��a������}��nY���?��c�E���	�#oh��G��w���<��×���rx=���_�=��}����{�X��	��(�x�v�N���3�����5��8��W��z�C�O�y��=a����}���_���'�2z����4o���8C�������E@�^��
"��>��<����a|�NO����985L���6�� �;9�&��(<~g�n�*ˮSr �C�j���k�,F��(s�.Wm�}a9�O�憺q��r��Q����{�� }	�DEO�{��x��0�#��O��˸�����O:�G��y=��z?q9�=hz;}/���O�'�x�w��p����""��=ƞo2�}�>�ҟR"(���������!��|ݏ��=ף���u��6�Ul����dsy���@{���w�;}�s��|�����9^�z�Q@�F]=)���{�Ӷ��G�w��x�����:ƾ�q��j+��&����"��a~Y�����@<��|�1����EҾs�>bM�N��Ӂ�5Զ/:�>�i��"��?y�zS�1����H�
��x�