BZh91AY&SYy���_�py����߰����  a6�}  �    D�        �T�0 >�                  }͵R�����*��&��X� �	�� 7��}d�$(�m���O���޵�ܾ�o�ù�=O}�}�⹳��^������;�y}�(��|;��t5�����Ͼz=�gۉ�=ۧ{�g���;Zi�����{���Kg��/Z��@y � ��b�T|z� ��_m���_c�����x��m�{��{�}�۬w��F�{ǟ>u���$�2.㢘��c\�w�gG�||}_��ТVUw�ǶW��wφ�I�O����Hwn� ��E/��ք(oxy�6��}�{�!��M��s{�p�3ݺ�1<۶p���M��i'΅�C{����"�۾�����#��̻4�J�y����e�=���w� �{�(�8�� ������͒K6�S=���[yٶv�{�� +k���w�^���f�q��P�S��u=����>��w�}�fQﳒwۤK����0�3����]�K���(�mn�S��4��mWZ��{���}c��:�'m!�xz^]<�g> <!�W�}��z�z�μ���S���b���ޏ.��e_Z_Y�>�����      AT         Q 
  U?H3�)T�zL F	���	�� L5<R�5# `  4�)H�U	�M0 L   ��IU$`i�  �M0��$�"h@ �x=M'���4xS��@TP��J F��i� F��&�3��d��D	$RF@�O��P�۟z�5��* mKD$�T�6����� ��9$�G����������
����K^����{�w?������/����4|h~`�~�c#	
����9)Z�(�����*�"/F"�Da�A�S�Qs�C�?�P������?/��ꕓ%��]2\��S���8i�H���4`��w+���F��'J�J�C����R�4�R'_�"�VvW���L����J����L6�������w)M�D�2��F?L5١��.�Z'���NSL�5�㒒��*��r���Y���f�Y�4p��y�Ts�npL�U'K�Ue��+�N������]�9:k"m�*V���I%A�������}����>��lM�)�Fc+���Xs&�bL��RW$Dnu��gd��N�{Ubcʮ�oq�T�&UR`�β�q�J���Ӳ%�2&�������"P�L��	������s��|�H7���}�d�}�+W�ߎ|s����М�\�xӠ��X�L���)��J�>���]Ӄ2��IlIz$��Q��)7�)(t-I,I/$��O�W���Z��FIrn;�&r]�#��9#���2��!
�|a�Ț���z=��}����w�K�S��&G!r�HH��xMp�NaA>�fCG����զI�9�'h�r������s�3��W>ÂN�Խ�Nj}��s��9F��m%�KL�Ժ�'>։ ��WJ:���,�r}�r��hH�;GPLF͓D�����&�hѿ��r2}h��Iz!p����;��2P���ޚ:�����h��6J�q�ԡ0H���ko�I�
8��������Æ�%�&DK{)��lM��+dD�&�?,��N-���J���\4:��d��I6A�D{8��k�~��֥|�D�O�0j"=쯑�]ԤG�����ԭ��r�:�Rk�^J٢�#r�9l�4[�Do%p�0�D~��F�JDr%ߧ��R�4�Rk�G��R��벾~nR&�R�&��Dر:h�(���D��D�2�h��;GG���8QC�	�R�1ܤ����|ԤM;����u+��+���#�/s�i�nJN��+��ܤM7)�ʳF?L9١��,�h��K���+RDM��r��_T?`����Y�,Kd�֥������7�=��U'K�Ue��+�$��٩����Drt�D�2�O�:Hp�A*��J15*��}�UL�#ɱ6ܤY�f2�kq̕�2J5sd�W$D�Σ��a�(jpN���1�WL]S�$L����%�f�h~�l�S�$F�NI���յT��U�:�9 �},n���G�-�A�Hk��䃯�ܻ���5+2f�%ð�����0��N�.����(�]H-H&W�ړ�I���ҽ��0���,ʒ�$=	�I{�{R��O�I�����bAy$��<½��RŪ�U�d���ɜ�q����I�5'��[��w�}l��C��Hs�q���Is�-��j]�����$I��	C�H�>4�o=Ҽ�M��A1BBy��SUGbvϯ���h�9�f�"j�u1p��Be�p�'p�&'LK8o}�8�� ����	�8�`��'I��5Z*$H��KLĖ=)�5�p�	�	�1�=(����>�$�sd�:�:���L����Ze$�N���9	����NC�uB��ݗÆ��5���&����[rb`�I0�WrI��܉-�ZB�'S���	,��Q|�N���3�i�!}5���ƃd��C�%ĉC]��7'��i���)!hu�p�4h�%i�BkI0�e�#�rK�>�"?tH���'p�!_'Q-6&m����obl�H���
rG�I�a0I�La3��-������:Iѳ��J:��7#�S���e�t~Ä�t٧����fD�c}%	�I�LvO�3d��I;Ԝ�D��Qߝ�K�D��0��	ٲ|��D��8���wbjh����A8Q���H��J�''d�C��:'�q"hw��Wh��ğaҘO���7���Ԏ2Q�0N�N�-�>Fa8h+I+�)I�E}N��"q3?&�����c}%��8"btSe}BD�$�ȓ��p�$âDD�l��L�RQ�$L�����xO��h�E0���7Ԙu,��FB?_�9��
4�Τ�&	0~æ�NsBv	�1�/F��}���N�/�����pI�0�0E05R�g$IBs�Q*t�N�:�+S�;:ĺ;�?Q�ڝFɻ��Y����%�<�D�Ա7��L7�gw8m&�M��C�N�F�p�HX��Z�*���&��E�lJ��67���,Y��,���5Z���7��l�u%����/�+��%u����9�ȝ'L���"&w�0��q)%��kD3E�MD��7ڈ�����O�z'2��]N����<9,�M�ڜ�Nu�Ϩ�'N�d�����pk�pG�Q�\�ٲȔHԯ�]������o纩f˓�N��#s�Y�h�DG����f��
��ʨ�6�pNDE�Y�}eTDM�D� ��S�#�TD��M��A��uQ:oq�I;�)��Y��`�"'Jd�Q��D�Ԣ�'cS�O����T��<ʉe]��I�d���H�"'K8V�`�U�&֥	ĳ�O���T�ʛ�N����f�ڔA��GZ���R�fTD�ڜ �|�ʩ�|��>n�"e��kS�G����S�aũG���O���T�ʂ�*"oMJ ��#�TDΉGG�"%��g���&�魚:jDy��"�4%�tMm�l����y49>�܏�}��G4t�ܣ� �����ᠭϠ_�A����h��Q�&}h�w�h�y6&��WD[��Y�¬���E��%�����f�az�Ӝjl�^�>��K��Q��־���pH�����!>�$�g�9>C�>�S>��C�TF���Q�'$�����K���i�Ĥûjt��t�R����'��_�9%G�������,�o�Q����[.>	=O=�����t���������H�4}>֏�����^�.�d>�H��#��}�G��|:N��K��N�u������n�/jt�ڕ�e���G����M��?^Tn_Z�r��U;MK��";j`��|{��0hI�CIx"/���4d�]�N%�h�`�;N��G��d�Ա����г2�s꿤��.G���:4���>���D�����[}�Ǔ��I5;'�܉�Ա�cq�Q�w��#���(Vi�$\4L�!�s��>��4�B��G�$�O�npK��*a���K�Sw1�eT2=�ar}.O�(�IR�;$u���Q�v�#S�/[���|6$��l&5�H:	b&�4{">��C�We,��NT��nO��'"Y|�"_F�� �'��+��~��֥|�D�O�0j"=쯑�]ԤNr2",H_�R�&��D�H��]4V�$nR'-�f�~���F(��n�"]D��$�>jRa�r�:�".�a��e|�ܤM^�pN�����:0Z�d��a�Q�#Aspg����#�S��r.+�c���1�V�	K�[?�{��BM
7,	I�,{OGX�4!2����f��I]]��j��h���pf����w�G�gXkaM�F��V�	q���t���]a���4�V�����7	Y
�-h�#��U���R�N�ş�cZB?/�;Y(/>��6c��+p�DlP�����7�hٕ�d"��a�$�M}'a{�a]"23��	k J��a�Ne7��Ӌ��p����X��rV�xڈ�m��Ng�͕hP�ƅ�4T�n�E#��lAi�B�r�>=8`���Ǚ�!�h�
�iW\M�H�i�*øm���+�w]?�a��7������1�+�.��ݲ��^�Y�['���)'ޯI�U�N��QWc6��񮾱�R��z��VX�[mi���mds�=6W��K4���vOg�:1a�)zI�N�P�2TS��:Qp���-�U,%J�l�*�2c�h��t���?^��=4�K�Ôk�	^(��N���ѻ괝�e-�#::��l��Ԋ���No�W\*�F�/�iD����GY��.?eC��������XQ4�N�;5̅툑�1¬�w�?=0�=8p�5u �I�����5���܍������<p,D�MǜE���'\��O��37_ĕr�҄Sgٰ|t���Ǣ#���zq���c��ۏ����O�'����7��d�(�-udE�xY�Y��F��/
�뛍����ZM����ʍ��)��r\�{�N-M�Jxy?�֕#�M?Lx��U'�Lj�O��'r
H%��֯��7�۩7:r}�`�қ2��0�3�
ms�9U�56���<p�&HK*�qd?j�Kj��r;�p䲓o���9��N�����nB>��B#$Q�x������s
6����e�Ϥn��[�,,ef���*�.�������n��0�(�T~q��6Ui' T�l*����������oM�9|<I,�Fn`,�q}�~�ҏ����~X0�s33=�9�wN�xm~��n�y��w���6S;��
�co���ҙM�&	`.��s
��%;�z�5[�FU��cYr�2�
�b��j��sq��M͌-5ib�2�l��.R�-���\�73O����l�s�2TYS���Y����]��x������y���_b���\��et�OM==�o^�������O�4椆G��5-c�)k�lå�w���0�;��IG�Uȵk���CCmE4b'��72��4i���9]����oZ�^(�=�>�۫[	k
$1���A"�]�l�d���l�Z��^,�r!�"K��FfL�.L��/t(�ՕbO���6�a�.�.?oy;���ٍ,��I*�)z{�0�<�B��s��0ll�����'R������⨬�<�6���zwz�]	/|;p�s6g�������M�����W��$3�Pj�;�4~��zq4Q;0�P�p,�,vc�ixr�E]=7��=ƻ,�;�B�ב���ˀ��KM#�}90���!���I7{m6�}5�?<����s��F�a_wf|}q)к�RvW�XH�N�X㌧�Ys%�L��1���a'	QQo�1<���=��r>��C�[��o�㸉2�/�1��L������ZW3	����醵��Vuf�6��^�x��Ӳ�{�b�;�0�OF�xED�v��2�ܸwN��}�8k�qn�}(���d��x@%݁#�pDK�@�Y��GȦb��az���]dw#��i%ܭi�ޘw�#S;��x�_{F�����s�fc~A�O}���;)��m{��f��d��̊���sB80lDo�Դ�X�N�r�O鹭_�ᕐ�$�]���:�J0�㬭YBʙW#���K
J�un��10�,83�6�7N���A��Km!�Ͼ]�õTsv�4��4�6M�_<���=8ott����8VW1�+�a�u�����n2w[scC �^�F����Æm��d&tw�릚zT0�����6ۍa�Y����ӓ�2l�de�הB7�+U��E���_���rV����NJ�81��\�$|Vr�����$$��a�߂�;�h��ۨ�g��k�HWpَ<�%,q�V�Գ.�����)�a�o���ގ�ŭ�Ī��fo���RK��sk���O���J(�����j��c8����h�O��+������N����4���No���������2Ǉ
�ffS���D���5��)�&|�����a�*�e�=���w��1��o^J5g���I�2*k�#6��n�5z��
.�9�Ȼ׆��_|�}�>��5�ѧ�MU�z`�^��Ҋ)<�����m$��G�F%1��q	���������M�a��ږ=�s&<���yfaJS��ט�2�ͨ�6��VU7n�ç O�2Y���\���ա�Ռ��������A+_�޽˃�p�f1���4Z�NL��#fc�QQFJ�,�;���s���1�Ӎ"��cα'�g����d��>P]��V~�fW߻vfnH�ܮ�yQ���Ǆ�9�e��V��� ��}������F�c��J6V����ٮ5��[�M��S-���z��Ɉ���,+.�9��3�����3�v爆?h�M�re�©���4�g���2�ڧz5$���N��vRw����ˬ�ݔɇ�=�i�X���IE9�c8�f��n��:(V�B���3�2�������ң}{̈2����&Ǖ�5_���>�u,���?^���+���l�a�xd뻸���|eaӄ��z��}{pbE��P�WFFǷ�S�������[�������+Y���w���t�_j}'�e����.�i�F��ܥ4~�p*�,��A�?z0���nu�R�+��Q��l-��x�"�R�Z@�`MdȬ�;���I����^n��(����ե?�'��/^x�l9f�aI���F�?�OB2�6�w���wi饳O��&������"��zE�V����d8]g���&>���p���D���+Y8.�2˗2R��2fa���¦��:}��N���b�uo���=}}iT��d��o��2�n|g~�����y����f�ꞝ����e�̟~x���Cs<Q�Ņ���Ɲ¨��������,�����_��珽p�wӷOU�Ӈ�0j��W?V�35��)�$[5Z�����u�*�k���*w��p��I�z��Y�"z���rʹ��(K�4�?tPC��=2Dz��該
����_8z�����xޭ6n|��m{�ӿu�Ւ���S��h!V3,gԪ�B���t�uH�xك����z��φ����t�R{���Ep�0ׅ>�9��:�~37;[���H�;�������q�J}(��?N��}����_���{q��{��������Q��,p�?�o �+O~���ǹ�NL%�Ʃ�M+W�T+
k�Bѭ�������>Z�u��xw����m�1����Y=>��w#Y��t�t�pf��ė[��?�<#�p��&2IΒ�y22e�j.�C�O����C�c2f8K9E�ᰌ�a5�3"5�q�ڸ�s+D�V-U��fŚi;����p�.c�]�d��ӛ��'��jd^�ϖG��޾����k�sJlR�,BJ���N�&�m7r�W8�{2y��%��[�鐦v5��ͫ1�u�%��[��w��y�0z��� nw"At��Q�6Z?}���y���pd�^�6��=���C}%��:��*�@̿nc\�g���?���~�Tm�����/�u�l��䁔�O��m������,}�BO�>�J�A��?��0�A��'�������A%+���t!��ף��j�``RZR������6�)&�����:K:"X��cwL��9ӝ#��]fᫌe2ڑD[ �A&}��E[���Ⱥn��[f�jb5��~&7�V}�^2Օ^XY'za뫋���=������w������յ�E��	tؐ�s\��ux��"or_w����H3��!�f�rZ�%�q��HB��5\����,L+��k�1z�88�W����ڭ�5a�R�4�(�l���z�M[��:�-�[�K��e�D���6�Ń9�݅�9��E�ՑA#��toG]��lbm����g2��(S��<�"�\��ˈ�_9�6���>c���8KE:�-9:q��h���5>�x�F'u�6i	��w���م�;@������`�����4������8��К�n$6��f��aڽ���cD�^���B	�a<g��2�[$��f �Xa�D..�Qqn����7Vk�(d\��v�#��ذ���W@϶�c�f�� �㇍�,ā��XYDK��kR��п&En��GI%��]tJ��] �d��������޶b��K�HH�K|����Ց�c2����P���T�vCjjj�\�c���w�Ͱj�װ66�Lb4���y�-���&��zAg'5 ��䝆���okl#���i�t��5*�ڨ^;u�LRX;K7��(G)��������BE�)G ����j����+��0#��A-(�jF�E=>�4i�ё�T����ְ�HJ�C���z�o;�3W�X[C�|�?g��^/���m���<p�'�*�q�ȁ"J�6E�t�#*2I2sF�twH�҉m�N"���u�==�ml􆉪
7<(��J:4�w�����T��E����Hn�hHj�H!G���Ά���K���	�Z�Б(��x$f�NoH<[�	�0H� �J(�ĉ�ļ���["g~A9�`��[��I[��|>�0��������|m���Kc�3�>�|UWH��E�h�G����:^���t]�[6��M�p���I�[Y-8`q��lk�?Q���}=�㍇L��,��	����h�ּGO�A�n�T^z�VJ�
*�쵟,P�ǵfgзЕbH_�
fL���mOr���H��l�Pɤ[u�\#�Mα4S7���
��0ZO�'iOZ��@��;o-�����g����(\bV�fQ�δ�#5�fWW@�B	��
�M�d��Y�a����淳5��J���}�}|�  �-���>_��!���̄�!P�h|r���_������@�#'�Tȓ�TO���������k�?�mi\b���*��t��Uҫ�W���^*�Ux��Uڪ�WJ��Z��[W]��V�U�����UWUU�*��Ҫ�WjҪ���]�1U^��Wj��Umb���U��t��EUW��Uҵ�i^+�!�>���$$�ԶYdE,B�-DX�MI
��6��A�$VE�dF$AP��XE$�n��j-H�$[�-~8��.�UUQUUQUiU�W��UҪ�WJ������U\b���*�Uz��U�w�W��U^��Uz�*�h�����kJ��^+J��*���Uz�v���V�U�UW��Ux��iU[EUW�U6��>>9��$��ꈶj�HZ[V-��%�E�"E*
f	h(ZTH��T���ն���z�&�J%��b��ȩQI�~	>>�}>�$�����ZUVեUmb��,UU�U�UKUUQUUQUUV*���U\EU��U\b���*��t��گ��W��U^�UU�UW��Uګ�iU[EUW��kJ��^+K�W:*��ҫ�W�Ҫ���R���@	Es�#5dV�$�H�0���;�VBO�� ���h��h�w��{��v��Uګ�W��U^�J���U\V�U��ګ�Uv��WJ��UUq���������1UV֕U�U^1]*�Uz�UUb��WJ��]�J��*��*��t��U��U\EU��:Uv��b�Uw��Y$A�$RA	��%EJ�p��hTD$Q5h��e�vA��ZAjIAY�ؠ�*�*�+���ya#t��5N���	"-�TE}�>X��	 )UmKj�����s������	�}��Q��>��}����͜8l�!@� � �	��؜:tN�D�DDN���8AD�8"X��&	e��
� �AHpM	�BhH&�N��X�&L,D�,L��:'lDB�M�0K ��М:"p����4%����eHlDN����B"P��Y8hL:'D�f�6h�BP�A���B�M�"�BpM	�Ĳ�:Y�q_�;X����l�x�u�{���:�W�bݴ��Y�y��Ժ�4,�BM�c6�A-���o���"����Jg�Tv6I;��D�K\?	�`_a`]uI�4�͆�e�s��,sԗf�*lYf�A0ۦ����k�p���Mkd\+�fQ\m2۹9�a���DI�����ZjJ7!tś�%���P�,6�3�/5(�>җ�Z�VS��5���,]H�hh
m����x���e��~/�a*�P��`���@�R��&PP�S6|T����lb$��1����$.��e�Zfl�H��u�����|�z0�ִ�j�MQ�XM��@���E(ޛ���k�|�q�v�,IHy�g���l���ș���KتH�Pq�;M@��E�B/�a��|��#-**C��	����Ox��$<��B�{ޒ�'��u]�H���d�f��H�u�jQ5��:���I��[6"i������,�$�>�����j���:nu��W���|Jx>�5�\��Vi	)]~��	s��`�إP�)g��m�jz��N���ύ��g��%�`�@�dK�V~}���Z�����ZdG-FK.k�v�B;q��ϛY���WW��묏TY]l�¤�h��nB
�Eee�B�Ď�B�0%�0�ग़��������ͱ,�	R�?{��#�..�W�k��x��Ж[��#Lk\뢲٠�Ql<Mp4�!Y�K4�s� �m��-�v�^MR��r�R�n�)���<l\j4������(�6cޯ�[5�D�J6�ӳSj����nD6e�fj�I��V��r�B95����i��Bi �b�6_[ɱ�x�:��͒
�Pė�*,㾴�$��`qg�]�7��j�U��]n�ؗm(�OiyÅ5ifM�C���$W�2��L�m��'S�!��]����6T���$[a�J�$e##.��2�,*�d$jbF�|����>s33�*���W~�����sȮffyEUW���}��s��\��򊪮1U߃����<�s33؊��1U߀ �ﾳ�hCeٳBhM��:"&	������s���Z�e�i��]�]K��f �A`F�kbk��-�{%��̉�B�R��anG⎲d2���X&R�f���`Y��j\�tghH[��6�jQ{93C7,bĩ6��#I�R��n�M�la�ux�-.o.�g9���G�9u�) �������	�c2ph��R�	A Na-�$b�����BKe���`w���x9
~0��5W�~�N��؟d4�4�L%�;��f2Z�
�$)7�'MM'$�QR�!ı[J�v���=*#�"ń������Noh��>�X$wڤ8c�n�J��h�]�Y�y�0��OG�8,C}p�;0�}ӆN�4(�͚0�f��x舘&��	��\�M�I$��C�0�����4l���\���x�F�2q�yz�d1�+ub�FfSi*e5�!%�,)��	��F0�8|c��zP����,����\C]�`�+mM˭�u�]iK	ljEU��ؗ2�JM�C������r�%U��`)�U|a���u���HIeG�p~��tM�Cf�hM�xN���l�(�0��r�MWUK�Ni�圃I�b����Æ��p�4���-�IgD�d�[��8tU�����>;�3�þ}�#l�l�8M4�,],�w$�t!i����'��ᴫuYuBVϊ�cRR���40R=�����O>��ҫE̻�%���ɸF0�XóM������(����4�z�>Ե�&H�Ɉi(/̡I��]�1%U����v���{4���xq�q��6M�`�قQb`;�U!5$�I�NT��̆�d2q/�&5�i�D�����0��&RN|�N*�6d5��&|C;�\;�܇��i���1
�E$XL0�zK�;��!TMc2e���+î���[%����v������Eك���Jo9�QE�
�ikQt��].� I�Oʎ��B(�͚0ц�ǏA�����ޒ���D�� ��TB��C2��=w!�5�)H���$��3%_��/�t��x��*�1l��;i5��݁�5g#E#w�_���=�e��إ�*�1jMV鋓g�ݣ�u ��g��S��{UT��gf�tJ�e��d��)e���Cms\:أ�ԛD�Sf�d!�{�
k�����:;.N��j�^���E=���#3	
x��K˂�)��Y�V�[UWSٟG^��:iϖ�i�:��� �gY���$!z&�x��2<Vo����IO0�.1{��bn����9�p�������d�! �8�d���=)�i�M	�6"'DD�0N���WUr��m��u<8�i�ƞ>�8jq�J;�����I*��x�F�9��H}ɝ�
,���i��΂��$�.{��70م8[#�u�����H4�ƹ����L�)��R�إ��ƛ&�;F�B�̎'Ls�	���v$_'��m_ôߍ7N|p�f�(�͚8h�e��"`�'B�Ô���u���7�k��$�r��Kh˩ H#cAĳ�J��<��sI'0��d�Ǣ�3I���'U�fD�S�;�����F���+����뮥n(�\�7+�cQ_<xǓ��̊�]�I����Ṑì��C�s�|I'��,6$T�R�l!\�CZ�`%��e��ٶ�b�r��,4��uԂ��q#�k]��nԽ3�y�0�i8�̷�:g�ͶVn��'g�%�o�`���gx8C�7Ӈ�gP�)��f�	�6a�tDL�X�M�k!'5US�7��s����U�`�I�nS;rq{b�9���K	�bת�w5�*���nu+a��ͦ�6�p8�0�X��F����=Jt�e��%(�E&���hLv;�ֵ��m��yg}�:�{�k!�%8�I�i&�j�U�88S6�&�QL60��r��\��޷O7:��'_;t�ݜi\q�m�q�	�0L�ba_���H�2�����k���+6��7h�ͬG[\��6,��4|C{L�鎾��J��1g�ϩ�5�H�����*�T[���3,���2ԅ@,t�.�f	V��nᬭ�`�+f�f�-,��mXNI$���u2�T.�R&^�H�õ���
T�iBDFHdf��=;c�X����G���)�9\$d�%D�CI���>�¶��ϡ��|�|�eF�)7<$`ѹ��b�(37(���R�dm[0��CIs�GM�ǚ�HCA��F���#��kvI	$0Xu$���y߈�X�ѰV�j�<u�!���(g�G�j�fw���kO�ʴ�ϧy5��cm�8Ҹ٣6x�:"&	�t,L5$�)z\_
8ON�{�{�pzgRYh�Fq6h�.�\���07�H[P��o����)Ik�oe�rd�,��ϳN�sFyiK�g���w��r��Dl����V�z}J8&:Ic��2DѼ_2t�Q��	c�k2G2HRB�G����w.`�	��h�Md�]&�ԝ_���c�[�v��v�[i���qk5j�%��/�-W�e~W�쭩[j?4Ӌ�g�_���Oǃ��d�z?G�t%����'���5|cx��1���ƫ�cmc5q���/�ո�..>jc�[��]>&��K�O����'G�W-���i]+���cS����b���L_�z�W���1�\_qu1�L^�4��q~cL_������M�q{cXⵋ�۶�qqqqq�Z\Y�5���Ӎb��Yomb�|�,�xƦ/v�4O��~�����N��~U���\x�.+5�;ok���5�5���b�5~k.j���]yo��׋��]�a�х�e_��?�[�\[oLmU�W�Ūū;sV��M1����\W�1g��JvM�f�l�n���ҲJ:Q�(���/�X�f;��S�?+�4(�J��&0���/�|]]��D�ޜc}���z7�Q��e�����z���3p��A��C���K���Dݸw���{��σ�����33���UUTU�����9���333�Ŋ��������o&Vffg��Uqu������ef�3=����U�U׾�(��G�+�M�m�c�|�>c��a�������Kn�:l�y	!$$�07<U!���a���UC{�I	u.@�0�I���dN)zQ@t��$8�R��s7V�,ܠ�Q�]��� @��G�G#}���~�N>�2����t�Y3���/i���&HK
�١'�Ĩ��Q�u��	��e�<(�'�ZSH�r�+�~��OpLs����V4�aN���፼{e��,~�}�߹�wߍ�4{OV%f��ٮr6�Y�*�ڟT���t��%*�Xߪ����a�F����rb��<�����8b���Xْ��WN�z������׏^=c�7��)�6�-�	 �	  N��d�.\�d�c��j](�6��E��<�4��@�D8@ο|'�ѫu��uP�j�3��h�J��C����q���)�>[��J|��R���&�Q�m�)���p��A���2�gbw������Q^��m04D6�I@y�� Sd �^5#��U���]R�͛�N�f��t����L.���Pd�%�(3}�~E;4q?^�ÆSjdTY�M�MCȬ�ȧ���n1��n;SÎ�Ӧ�6��~:"&	�t��Fi3*��M��W�Y�YPA���;�$ћ#)bP~��PM��	�<P�F)&,L\��fQ��QK���c&�x�"V�M�)�Kr�[U$�X����2�����L��f�i���NX�ܔ���G�߲ �HK%}~G�sJ�j-��3�)���b���N�ٝ(K�:��f�}8�}Q��Ӎ�Ѩ���X�rTj,��,A6ݡ���>ar�j��U	D,�a��@��8�$.y(|#�{��h�Q���/��[]G�d�^J���#j���Q�q�s�O)QY#M<���p���|����`!� p�HXT:�	 (�th|	��H��JX�)KC<�(0��C�3�	����ѭ��H]�+�-����wo� ��07�������f��2S��D�ꪘm��&�2�z����x�G+�h���0L��O��SӍh�RRBHI}�g�|�) ��ɒjJ��g[!Ij,8�.����NR�m�vh��ER���+Uj�z���t�!z�v��-Ȩ�t�,���Id��B$uv�b�o5�َǙ�;�%���֋'Xy�^���-s#�;�@�^�
Hl�ADJG\�UHJ�a������-ۆH� g~�Zj�7һ�4�x��]J����;R�;YK���,e�f1yz�	���|^�J�\��9 vp4H8����D�pN���Qe���yJCD�h�_%�g��ƚY�M�0=�(�� gRLJ�т�Tw��,:x�ۥ:8�]:m��~8x��0DN�A0��O��;�ۼ���֝�I	!$&	��U�j��e���)<�2+����Bɗ%����u�,1��ܖ��nA���0�N���;�3��Ңӿfb�b�X�ȴ�XݡoR�[{�blY6$��$��8f��bN�7�?���v�~m�JqP�q�K'�Y+��O1#���8~��p>��o�SW�#�j�,6n�u k�K�M���*OQNtd�R%��V�A�X:�Ӆ��ٙ�RjFq��!e!�%�x4�]"��k��p����pX�p��B�8�h�D�䁂a��F�8\v8C�h���?��0DN�A<��d��ȟ"A�$�����C�8Q=��UdRHG��ئ�є��P<��E�3�'�"�$�p�;�^H��ݕ\��iYǣ6b�*j�w#�Z�ӥe���F�~��l��,%�K�=%Q�%Ͱ5*b���+]�eF��s]��!Ў&CnS�<���4�/Y�����kcr�,<Wӯ����>�i��{�Iən�����ۣ�M(��"А�{�*�q��Q�����O���[�=�J������,��ѥV�?6�t��6��=tO�DD�:Y�П�aTI�8yH��M?4Ɲ��C�l����̔�A��)��8�a�iaU	- �J��0q�(���hbH�EM�.ǘcx�g0�(�hU�qe��07����JC5��miRXKv+M�ح�u��&[=���ϓ���@ �g���,ҭ~nn�kId�ݭB�p���,!c2�p�ÇXV���*ů{]>US?[l�&�C%%拐�&誔Kzn���!�x�� ���z�C��nn�ֵ�y����E�KPy��%�X�������S���5��*٭4����喧j*�M�dԮjqcl4���0���x��U.���=Vg~��kv�I��|۷�F�Px�ć7�7! �
={-b�L ��!KV�C!�O1��1�P�4GgF$��2+��z��A��R�p�_-�R�v+Fȝ�7:d��Xf�
��!U+)��G�^�0QgMXl�4a����0D������{����:N��nfJ=�AUT4A���y������Y�SI�I0�H?�uݍ��<U��*���!�y�燇?~Rd}(�%�L��؛�}��h]��������M&z[G��M���5���<8L�>!Y�C�k�׍�M�յL=�<Fr�Ԧ�^MݗJ]D��%$)F��>���8�0��q
C�4�|y�R�UATh�l��|hpA�t�K���.D�[����dx�ks�lm�����8C�4'���DD�,�L?f��	!$$�A19�0�Jt;�8��=.q7C�n\GitŨh�;
B��%J�7��F�%Y�����'��κ�	�HY���,U�rԂ�@�wq��	ѫ�j��A&�q�����������ڎ��L�)��uD��=3���:�LL⭨�^��K�(a��ۚ�/�����Ւ�a�w���	�����t/�Y8tܩP��$�􅘅�: ��oɶ�I��M�?4}a��8pК0�pO�DD���ӳ��<�^��esw��%'!$$���&h��:�vO���zI�WfҘ4A�fM�K�w���_�̈~bV �L�_I��M�p����ۈBAM/̽w���Hxm{6Ӡωa�G;�*��|hִ�=wmjK<��6�\�`4�e���Oj����u;�U����9h.�sfa�i<=6�zA��d�R!v�GK�Kz��q���8z�cӅ7L�Lʪ(�a�i,��$ÜL��g���O��O=i�W���b�}�X�..>i�vƻWJ���²[q����XV-V$#�!��Z�OS�6!�!s�7<p���9&̕�%���d���5���X��\_��wMb�5���wb�Ʊq����qq�Lx��v���ū�̖�~]Z��g�-_�U�_�������_�h�bΗi�4�w����xƞ�垱�>i���q�LW4��q~cX�1���Ƹƪ���loo�ޝ��������Z\\]+�5���]b�cLzk��Ɵ+��χ����8?I��x$cL^6��qq|cXƾ\^�m��W�.��.;k�5��qr�k���<c]������K�Ӎnۋ���>)3�~X#��~G�D�Q>]�@`�4~9���9�5��cOX�v�ׯu|i�ֱq~
��>�Ef/�cTO�S8x�k���M�/��7#�����h��9(����V�G"c	`Й<a.[M�y��v�l���fZ�d���)@Cs�7����Z�1�Ia�Z���q���y��f6ڄ���*ZEab��`'�c'�15)��Ӊ���A�0NȡS�i(�d��s���+\���dm�Љ�嘼��+��KQ��'�G͙�(9s	��d�\AA�x���/Z��:�7Pq�ֆ����l���L�a��i�X��QkXq$�H۹	t&x�V%G,�D�p$�E�cqc�.AY�YY(�@\G�w� �����v���t��e��)��?3�y�&��eҍK.tb�x�2&���Ic��·}�缯�s�:�I����}�#��$GH��Ǒ��سKfb218Ȇ �1d�zhݱ"d嵘��-�L*R��6&pz�N��������b�F�s�jޓ��;�l��uh�ۈ�Yp_ѷ���4u���X��4�d&0�)6���zt�rH���b�n�Ѳ��B�݋���+J$��@�݀_�Z�e
Ȍ��"!��,)I#�[t�6�X�5���0>��x���y�:�(ݤ��( ��!PFj��O�9S�U�r�q��a:�x�l���P�#�/����n�5�32�߳ޞ������}��������>�{��{�[E]x�����fk33���{^���z�W^�{߷�����{�׽�{ٞ�>���N��۶�Î�Ӧ�6�<tDL�V�$�2�U�b�1��N�����t-�bm6�ŗ�;XrM��I�j5�gj�۱m/7b�Z�X��0�k��S�A�m�݈��vl�9%���dV�ۮ�b��d�ʵ��{z��x�a��*�#�m\��2[	���k�r�ն[#�iu�CAo%�.2�M�ml��.�LIe���+��M(�4F�a�p�:��)JR���c��{��n1O���=�,	Io��j:���<a�'��f,	d7�,�NBc�*/3�>ϰއ���cl0�v�wUTW���a˂�N�$�Vܒd�M˜(��L�L%�d4��1Vbԣ�<�Nm���B�r Jm�%޴�ۓZOuc���A��`���d�m�������I�7;�-<9��!		 ���L��p�K��>gR�J��n���'ؼ�?ē�~����h�����P���B������/>�"(�Io)D��V]�N���66{�j�=���qS���Ӧ�6�����"`��X��[z�m�5swp�u7Jߦ����_�1�L�g�i�c�l�n��FC�を�D4q8�,�����v��@L�%4q6i<�M���Imw�e�bz�U���xǦ8\nC�^��*�-Uh�J.q��嶅�6M��x����tg��x�Ֆ�nt^r魛�_SJ�h��9~H�m�lP��n{Ȇ�b�sGG�&��s�6�zC�)���Sgi`�х�	�ܗ���Y��Biɴ�s��8�x�LUqҺt��ߟ�>c�0DK,Ha���U^��k_��W7S�c�&A2&y����'�4�R�%�!�ܺ[%�:L�H:#�6f�HHE�+Od��|Rl���w	�$�/ �O��ʄ�ѡN�Koio�'��n�a4C���G���Iy!t���iN;�y�&�	le(lD,珪M��v�KZSkR�^�,u6p�GSɫ��D��	G��*HI�$�cI�Ӄ���4p+p��!�~��šUNM�M_9��-;+F%�y4���ō�2��0X�G����㧄L�VI�ژ��*T�R����&7���a�6\lAɂ��N.�<w B�����tŸ��6�58���W�X�9�QH��C9���s���>4�xA���'8�i0쒦
�cC��!����X�eB�X�V<��a�$ɳ&��9��!���rLW��UO3����m��q�ò&y6�J�IU�'N8���a�n>*�8��r��8QÆ�4'�����&�e���}�u�(�	A�Q+NP��N<È�
A��yv�>}�{�&��L=/乚�8Y>@쌃DJ̨41��q���yS�鏨Q>oRNI�һ�+���H��(F����y9\��(����0��JR�%�z|>CL���4�q�?fl&z���{ǧ���{ϱ�%OR�u��yh��j���~���̎2���[n�۴ɶ�,f�Q�	����$���:XI���ICDN;�(�H�F��,�S� x[������t_ww,�e,�):C���,;n��\!�`]-E��O�~TS�������P��!�Ί'�ؒB�i�iw��Q�F~_'����і�A+R1 �D����!�&R�a.l�d�e�v���ŃɌ'�F�K!��|S���C�ӆ�8p��F	��㧄L�>�g|���Y�g�٠�a�EQR��X�����X��6K�Ļ4� �4Ɯa�I�L�`!��.�5f��5r�m�9�m��$�`���scx���j1��rq�RY�!!L�c���9�VLa&��'-�oԒ�Mq8�a@��}�g���.L���i�:�7�Æ��F�nхo�v�<Kg/L���^�CGy۽{bx�X�h,',qZ�s9��K� �8�c8K�t���:h���4��~6�m8�Ǎ�c��;c���e�?/ٳ�+��d�R�J��{�ɉ3;:�Ix��\t���Ӊ��R8t���X�<��tX�
ov.��`
0�L��.��\��e;�����B��*�KUT�� ��S!5l{{���Q����,�J<���١9�O�Y���t�GM�ǭ�����i9�G�5RJ�^��c����r	����J��n�]<;��]�t٪k·�,���І�5�F���$֍���l��ɉ��Eв;/�bք$j�r�y�9$$��v��cN�_F �ƀ��6�mccԤ�t�`xY��j��)%��=�ֿ:~m8m�m�n;m��O���xL�zˇ{Rk��ɪ*J�:ԮIΚ�1�b=�g����dnJ6X��$�i��V��׾�;�GE���� Og ���>+�=�d��J���t�a��@��D��w����}d�mO5I��+��V��a)#r�B�A(�K�]�G��&�F� 0j6_0�p9c�%.��Ίa����Q�I��}�O�Z\���%�W��ڤ��.��%���i6�x:M&��0��7C�����QUXt�](�M�}
�.Y�Y5�Rj�Sǌm=6��8����t��0DK,Ha�;���o\�Z޹�oޓ�D�I�;k��qq��X`�y�N2�9���r�Y��!��*n�r�!�M�bB$�`����'J�'|-�$��U���Վ�32;�,9��d|c�1��c�3]���׶�1��Sv�K�V�M�p��.�o~��O��i䥄er�����HX���s��JJ-c+�n˛"�m�Θ)!�m�%;N.mѓ�H���)r
7����p�9�Hg�N�,�wIKt��6���RT�krK�B�I�v]����m`Y#h%L&d�L�H�5$=RF��H� �!֜_7�$���(9�ydM�-���QbO��aH�ʚ�
�e@��>�9+wmپ'|+p���<,^9H'Mؤ�s/��:]4w����oVy��c��ͧf�W|�c���㧏	�"YbC�H�B��:��1��	��>!�(��Z��$M=
\LT��)�)�B� ��ܼnV���],�:�n�R��{�%Qa!�6�O��TRJ�HC4�2S�RX�A6kD,���I!��mk[I��sm�$F�ip�i�����Ni6��J[�Nt�L�6Q�nJ�[,�t���	��M������ѣ)G��5L(�&HWn�HwG�Ub�Uf���(�6��v��%g�MQ���s&�7=������#����q4�ߚ8D㦍�h҈1s'���:[��2t���ڹ�~V.>i�[�lk�t�\[nj��嶫�վ.�W���	�Q���a�`��Ú~!��g�8~!��?�c��p~,~f�5��ZxƱ�_�����Z����]�7�/o�b���jߗ4�-Ӷ5�Ηk��Ֆ�-��Z�,ū�U��iqX�Y�58Ƙ���Ә�b�|V/��zƞ��zp��ҡ<t���<J'��/�i������|W�\\c[c[cX�m�\V./ޮ����~Y�5�����~|�.��_1���cF/v�Ltӥ��]>kj֗k�7n�Ƹ�����������./cx��cX���x��.+-ƽ�ׅ�~'C��^�Jp~Ք~'� |X��ftB|*�A�����Z�ۍJ�\]�.Ջ�b�vWI���a�&��`�bW���:`�'O]�0'��j'��A�P(��T����%��G֤{��L@��i��+h�ԇ5M��랯!���:�P�QB8w��p�FE�*&�Bh�I	jD��`B-�F��5�K@�[�3�C<�[�
���K�p9�K��9�V�+�a�3X�=�g�.��	C�Bj��w1�C0�����ə��d�:r����I>C��8�}�ff{�U�}�{�������~�ff�3=�J��g�{�՛������f{�UҪ�����kZ�s33y��qWJ�Տ��k�4i<6���8��lc篟>xvz'��}ZFωM�mx�1�b������+�ȳNX��,�b�D�
!�3���B+
��R����,v&4nT��%5Tm��1&ZM$<@4lĞ.�ܑ�i4e(� C����R��ycg$�8�%wJ��95����:O���~�.����Bŀ�LC�4X�ҹ$�����؞K�!������F��F%�����I�z���J�SG;<Ed ă���vm�Zw��0�QP*�0�D�t�Yj�&!!��Gj=��n�=�|�z�������ӣn+�<q�|�������e�!�HύV�jkZ��vu�c��xd��C�?xB��`���E����J6Y��b��ف�'��nx���D�/�l�.�CZ@h�}�����:��rX�t�0[���������$j�r��*�l=xP��Ɠ�Cs.�r����~?+��aOH�6�9p�S�������\�0�.��� k	Prso�L���n�J6S�e0�L�W\�c80��Vm��ۑg�m8m�qǎ>q�1��Ǆ�,�!�C�jo��Cz�BXz��.�!R���dA�����Khѕ)Sc�xR�`I`�L
ٖ)aBQ�$�m��J|�k�А�F՞�c���,��MJD�;L�y�[u}K=KY_���� �w�<^ٵ�q	�c�p�4�Z�oq�%���r鼜%���4�i���Y��@,���������̩�N��V��~B��<�]���&��=JX���b]=�В�䆒�M��ݒ�ö���0����;wL�qq�M�JjzS�['eKZ�HI� l�L#�<Y�s��o��G19:�ɓ�9[���& ����<{��I���Y�j�>aL:=�!��m������}�����g/��=t����O�8�d��y$�h��%쒓gB����U*��0�̞.�wn��v��O��W��ݾ|��1�z�Ϟ<|�\߲'���٪����L���l��ҡP*�\��5-�a����f�
�Z��@���j�g
�ja�3��:�$�3v�&dߞ�$$��Z"l��������a,h�(�t��Xժ��4�O$Jpm����D�h3E�4񣽩*��ǚ��x�~R�X��UZ2��IbZ [T�PXF_��[4h�1�$%+!)a�"�!
��	l���J6Z���F��%�ce��Ū2��YmJ+h0�F֬u HQ	e�-�$B��Z-E�$aj7�h�;i(ڍ��"�K-(�9�m-H�����!e�ת���x�4U-��u+,ZF[�+d�TYbì).i�h''䬷"8R[�d,qQ�Y��0EYR��Q��Z�e���1�S��L�D�j\��PP����:m�IA�,62���EN�U���O;ob�$rQL:m���iѝ�zzuN�����[��YA�^/U*���k�/���J�k��׸����4�����st␕1��2Y,i�C����BC�UJ�e>^նw��Lz�Ӊٷ�M�m�	�?x���X�Ϲ��R���$���fC�q&y����}�e%���ɢ��4GG����K�5�&��ˆ�.Y4l��dM�7N�lє��O6�q2kەcW����M���~�Ԙé��-���g�y��=�(��D�$�㇄�Ա��R�S�ZKc������*."[a[6졄u�޽kԻ�kM%����F�p��9���L�i4;J9�N�R��UJ�C��.�o�tɑ�s]U�^=t��q\t��Ο��g�0��e�&�����,�l����>��}	������E2dM��.fG6�>��}��J�~��c�b���c�B�[5��݃�����'�����6F�J�i<�fd�*I%��<�.KJ�'=�64�x�rG	p�`)�a�8sɨMH��1���%%�C;�ZѲm082�H�.Í&K8`ܼh�ۣ���$���	$�[�8�}�*d�b���M�SP�m8�O�q��ӧGf�q�6����t�~,���,�!�'+�[O���۬]zKn�+St��V�'�����E!C
Iꩦ��pѬ��)Q�\6��U%����ɵ�Z�I�r���_]:�f��i4�6�1J~��@ �>��Q�M4�ǽ/W׫�%�F�ݝk�1�	K��A���Z�D�����Xs>/�z���VN�2<
JlF���I�Ɂ�zM���
�J<S�ɾ%��M���L�6�3��c�ĺK��fHzOT����KBC�^;zm��c���{���w�ϴ�"C�'J��.��]��s��#x���6��k*J$mEY�4���$&�%�zW�����]�̲��rp��a��E�.`��Н?<x�Ǐ	��S2�ZIj����$$��2.�;BG5I��Ci��&#*��]��LKA���K����o��v_��fU���~�j��J�)�����l�p�q�w.w$��*�I�rw��h��s;�7@]�yxm:��O`���:�~}zE�TVFIk��c&Xh�h�:�5������;�i2ĺ`ӄ��n$�V�̛���_uUsrBƶ��d��1a�R�ϱxAb�c��������0ۍ���	������Ǐ	��w��sZ���Nd8�^�$$��2	�\3��	�S���.��tу��)�:�R;�(�l�\�R��섳a����~{6;���,bN����k]h�!CGQ��qJ���{��`{�<�s8�v��q�zL���V�=*�*�tQ��R-׬-u�+���Dϭ�Ŀd��z��7�:Q�I�e����,qvBBҪUб�r��`NX��/X���iǮ>m������<'�K,,F�ڣD+�tUQUEU|��ٻ���ҭ%U����2� ���;Aܹ�̹�d>�i'�t���&�5,��[@H6�����$u��HI����N[J|s)��FUT�Y|�;��q��M�۱���J|�HI,���vto�-�p����k�E�%�c��Μ�����N�y!$�%�ы�v�HXã͈e;����k���x��3v�_���q�S<�]ۍv��k�af��Ū�Ʀ-|�-V��~UVյҟ��~S�����N��~i���V����-c\\o7u����ֱ����U�ƙ���mb����51����]ۍv�+k�aXV6��b�aX�qUX�V[b�Ir�$�x�x�I�>2Q�%��<P'�	�<W��~^���X�x��5����z�/����.�x�m���|�+ի�ƚ�qx��^��S��OO���4�L�'k����p/K���O���4��xƶƱXƽcX��:kLk5n�q|\��c��u����+�4ǭ=y��vƼW���tCM&��G�#�`�G�kWUŪ��U��V�ƥY����qqx��/n�Ř�S5ߺg��|�	��|&����>5l����@i(�T���ha�C#�}�J���u-�)�ҡydr�L�RC�,�LubP�\|)�d֨����b�)p'�*V�dR��� ��	4U�]�k�L��s)[]	�����E[�����c|�L��%�j��s���f
�)���B�X'�5t��V%t�2&
t�/Z�f8��4@���D���j&�7]t���0���1����s(���ӲRڌ���Z!>|e}�W���-��b�I��6L:W����E��	���<��AVq��l����	���!ۅ����MH`m2$ �YT�ݑa��0.ZiF>,b������r�9��'�z�,�FSZ�#;}�4=�]a�Kq�l��]bQ~�=���ǽ���u��6����6	�㬼�B�`�PF�8�ҡ�r�$�t ���j��%�8S��>|�����{�|��h����[�07`8:�sK�\�0���^a�lո �)��L�V��zy�d�me�7b�Ұ.�b�um(7�6{����W��9%�a%��X;؎e*P���Ma6\m��]4뮺�C�6J]������&VS��<b%�t���Æ���#&"U�G	$ǶJP�}PC�Z$��+���_~����g��UҪ�b��7��y��������U��}��~�ffg3=��Uz�]�����ffs3�ګ�W�ߎ4h,4l�F�6Y��lv�<c���<xy58�Z޷��O��Ka�e]�X��nlf������h�B�Y�,Z��;5�m#u,�,��#aB��(k����5�t��DvV%�$��8�WG���$��J��J�#c�vӱG:`ؼ�UC=���cVj]t�L�Q�ŭ���0�m!��0�W�ʃ+�Y���;b�_�O7O�~R]�.��;K��	�p�Z�2�%0�3�:ϰ�|&i}�g_Ý�x�2I$N�E	��֒L��w�0u���$�SF�yg��%��vh���>s;�j�J��y:y�v�|^6��d�����E����e�X��UJ%�Ͷ��w�,k�C�R[O���X�!�X%'�����{��3���6M��k/+-vsN�O��z��r+�I�Q��}1�����>q��n6ӏ�|��;~~x�1�����;�z���L�y����<UnnC��}�d��|p�zzu��l�%�bHe����I����	֎�N'g�%��s��!'��p�pB>#*�kV������)L,ٵ$��:4���O9t��K߼3�Y�����OZ$/3Z�V۶ST�������h���Rj������˓gzW�iU*IZ������]36l��$�"c<"Z�]r[���%rB�#wN!F�6�m8��m�c�o�x�1����vs��H�[�H����BI�����i.�\�Ò��=��L%.�OsF�)�X�t˄�CM��M77"��s){C�a6�Uɹm�[�[wM9�`���������<6�)0�HG�K�.\x�4HT53��hr������d0p�ø:�L�l[�6a�FM�Id�ޘ�P��*Q%Q�j`�E�9I��G^:�=c��6�����o��1�ǧ�ǧga���E�����L�\�rA��)L����]K���Ք�]����Y�(��جݛ3R�:Wl��6\$^̙�3��g\�ñ�an�`��<ƨ�2�"t����.�]�pwI��I�����d��H>4Jс����e��bY���t���u$��Y��}�̐�N�0��t�wbi4`���Nn{���g�!(���[�6�#��&By)�:HI�?;8m�q�����o���>c��@����%:�K����b�]%) �D�j>cG?j�]�l"�)�9#(���Yk$�vA�(����9x����x�M�h�xL-���;;X�0lHE^�{M�v���Mb@����в,6s��i��� q>n����0\��ͮ�Rk�n������a,�$�4���nv~γ�㳭4�]�ԢUS&�95�:7���֚������SiIb�c{�'-(�]����K�pm�Q��Ӆ���J=Ib㣦��Wh�p:]vd�ɖ<d�ؼ��RB��F��0$ˇ�xP�p��u��;!�q�+jB;�o�K-f!YA��̙�y�n&�b� �T0`)�0y9�s�f��0�	�(��ǩ<XT7׺�|:�G���txm�q�8�ǯ�ݾ~,���x�XY�rv�Gth��TUBI��d&���(�u��W�a��'N�NG[���ɷ.w���2i,68Sդ��lp�N�Ŝ����Υ���)g\�*�X��&�u2���0)��M�J�v������i�+<�tpPv�$���u�wk��N���`�{���gy�{�G�$���!��J��g�.��w�����ᶇg�Q�]�d*�IF��.�L>�m� i�Cfac��\|��;v�����c�%<�a��ں�) �@;�͛����ɴ�̦��P��j�2�^ap�e;�UŦ�~��M:�.SKJQ�.�lZ4a��%�?o�:���
/ذ�r4p�
!��6��1�DH���}��g�M���S�e�U)��t���L�t�N�i�̃�������l�R���;DۄJ���r��.nɂ�J�I�Z�Љ�;&m�fmc�-�.�C�9�f���R��|^e4��I��|�oQ�480��X�[�|�˝�uف�D%�V�8|�=�C����M��۳�n+�=q㏘��/�c1�^<<[5�I!$$�A��t�*ֲ��u�l�]0eβu��(SV���^�	z�SE��Ŕ78�.�I,�����#l���:������I'�=��2Å��9xu=so�|FN�!�< ��W6`�hٚ4bH�3�<7�\v\챓oq!$��L:N�pR\�l�tH���{	�<�e4i,�N��D4��<�$�0\�D봤0c���5��4�S�#c���Wt����1���c� �I�"s�a����cK c��M���̸�<Z�E��l�j� HDڊ0׎ܻ��E	<M<��AKh>V�b�<v�\O$�ģE��D���_�����,l�1�6v�Jn/s��͹D��H���J����$+�BqO|�-j�!`��54�n�	[�r/\��b�2HF1�
�JՒWt��?n�ȝ ��d�hǈƚJh9�Gn
n���Y1�y���d�yѾvI*�b8\��6��h21;�m�۳�,�B��!p�|yr}�?ļn�KQI�2I�Fa�$2g{���K!9le8��gTxoO��_��ա(�˦j3+�.�뺜�$6�Z�[%$�h���ϰs�J[�����#�id���drZHW}�jx��W���OHS�M!���z�����c�1�Ǐ�~�[��U�_��EUTUPѤ��ByçI��S2�>N�]h��R���Sb�JM8R�n��9Q����L���0���>L��J�r^�#�&R��GEչǅ��c�����<���lj��=,�j9y3�Г�q"��I5��Ob�<eݚ黭��;����.<���0�O1�F$���y�	hvl�!����� Պ'�=�H_o�i4t��00���"%�ӂp�B �tA4x4ұ�1�6��m������Ј�b%�D�"lDN�B`���� �P� ��UțBlD��âX�&`�&	�`�%�&�ق'=x��Ϙ�8�8�=c���D��Љ�,DM�AbhM��Bh�	D؉��L4t ��,D��&	�u���:|�|��4��6�[0����6x�ѡ(D����ΖYgK,Ђ~7�5�w�|�y\D����X0Tj���Ӗ3Xa�jm������Վ=��W�$���n�j=#���d���uΕ	�e���L��f�?�v�|Ӥ��s�]�/�Y\{Y��ֻ���3�����Uⴻ߷�k333����]��V�{���fffs3�ګ�W���~�������{�Uv��Z]�gM4Ce,�͖c<c�1����<W�߾�ֺ[��̕���$���1f����Mܘ$�#�,[��A�)��#%�ٜ������[:Ru���fϠã��	�aa��<�)�a]j�5!°�浖��[?P���+&�S|BQx8jn�\���&ۧ% ��QFz]��,:���I{=���g�cFfw���	a�*Q�K׷I��I!�񃍸�-����&!g!��UUΤ�wgR��������豜���y��Ҷ�Í��8�N?8�>x�������H��9	!$$�Ce˦�-��J�%Jn�7E$���6�ƓE���M4u�7�s�/��I��Îaīd�55��wMI����a���p�N��4p&)OD��5�::s�4{�K��H�0��6�)!�N,�]�:���T�c��4ܮ$aԢ�x�dƤf��O���'�D�x:!¸؉&��Mk����Q�_�"s�N'ɿ��I���Y7�N<tq�q����X����������������laݙ>�U�"��1��%�Lj�>WIeǒ�U�U����{��h����L�|vl�K��^v�%����/�RæĄձ^�sv+6�qmnf�]�Mie�]�NѺ�4ί_ɾq7�=
���qR[7UH2ԺS�F�9�R9��52오ah�ZcW2Tݵһ��?iң��=�6���m!��;<D��-�D�f%��X�}c&�ڕ*�Ȝa����WO&�5'%+��ێ��R�]�Gf�R���v�)z�2T
*HY�V%�&�x�`������u��R�&h�RR���^Q��%@�����a�����6C5M�fݲe����~�xy��0�?d&&q����Ȳ�5�Ҫ�����,��m�����Ɯvۧn<z�����1����<f�kZ�kE�]i�i�QUAEfHIc,a�ԇ��˵�yrPh��������0��y���
xXU&gG�C�	�]y$�f��S�>��ގQớ�U�p�BT�Ubd]�m��r�&.�.�.�Ū�eR�&2���Ѹ�}�^B����ۦ�m���)�ԩZ"a"B=z��JOh�ӂ�m�{�K�SFJ��ܽ���Mg걦ݽ|���q�l;k�m�6�l��G��!��^�JL���äv��x�r&:HR�������lW~~�X�~�b�G�$���\���EO%�6YÍ��8�O�|������|zvvvw�E�NrBHI�wNs)<ØL7��|"�z=�qz`�x���0U��h�0\x_�y�[axX���}��m��(a��!��&bts�s㖓���]��cu�kBi��O%���hK.B�ќ��I�!�)F����$K��'H�(��\�K�1�jc��������.��t���!I�������&�� p��lŝ�I�He<��:K&��6X��0`��GWq�n������lx�1������ٳgo[�3��	!$$�l�,g��"u�I��`!gf�Ӭ<��I��|B!K������u��q�{����;$�u�)m7U�����K/�$�d�d��i����d�LSCO`��@�B`��*G@����fǛ��t�q�4�z]l\�h2]nm(�
�ҍ��4�8vv��޳�s��s��DI�QU�['���%MS��s4��Ӷ����Ɯxۧ�>c?<x�1����ߺ���w�tֺ�Uy}l�Q��d�k5�#L��)��u�ApH��ra�DdoA���ĉ�PAM�{��
�hj+�c��uUl���Y5ѥp��$M$V�\5𽔲�� 		����C�5&v
.[n�l�[�"mrcGX͓��%����e%�!.C��7�fv'Ӧ��>W]�Nz��M����k׳���M���z9�h��3�a_f����qV�d�f7�Y,](.S��w4��8��.�iS��g(�(�ы6<e�Bz2.�ֳ�q:Ppӵ�g�4B&é�Ã�ϋI/G�SB[:����i)�B��.d;Ɉ\?�s��e
%��ɓ)5SK�����M4��<q�����1����>��_Ka$$�� �����iy3���^CZ�U��4�4l��C#v��c�/�BC�K����Bj�&Jh����ˑ7ɶA�rgxu���L�K�I8x�#��&S�:i���0����?��N'Q�<Ð:���J��mK%۔�"�f|%�Ϗg�tap��'����լQj�U���a�0ClO&Z,�)pi(-�	�\�7!��g���(�CO
��ϟ�?<x�1����:Ƿmi21�K�Ԅ��@�u���3�`�wG�x�1$<pX���<٦Ź�sEU��RM�D�Qt�C��-��-�ի�ӷޱ}%7�O\�5�UxR�a
K|d�F��T�(WiZ��Ѧ��a�z|�������<n!ؙ.��UJ��&�8@�&K'4i����xq�Q��䢞�P���d���UJ�(�0�t��i2],�2�8�(��}	�<��8L�]�Oe�p��-9���m>tq�q�6�=|Ǐ�,���x�Y}�{��IUI��UET$�3�t�R���ў�޻�9��{6��p�M=8]��}p����ժ�V��R� �4:�QB?���6{&w��î����C���ߜM�!l>����!V*��_%��ˤ�������K.W�3�e0��G���x\p���\4�ϢT�,�NPp�GL�aF',a�ΐ�I$�L��AI'���ɩD����=8�)�WtP�퓉p!����%�Q��͟���	�DL3���4P� � �ࠢ(��G�7�l�g�AB""`�P �D؈�0DD���g �!�DJ(�BlD���,�0L8abX��`�%����ĳ��DM���"&(,D�<l�㇏,��p�D��bl�f�#$D�6""`�X� "A6&	��&	�8&����BhJ���	�	dC��%	�BP���%x���Y�Ǉ�BG�,5�?bd���2�8��l�JO�(n��&PחؤHKc.�/�	��"u��Z7R�٢Ꚋƛ8��o2�u���P \�1��L�TD�1��2�2\�(���VB�H���;��&�(X�tz����0�v-���ra1��lv us^h&6Aa�OR���:ˀ�y7ٻ�[���7�<�v�*���,~�?O��3K2�GRPݔzٖk�U�BK�����U*%�}��?|���D���HFC[��E���i�|���GQgSF�	��i���PR��W$��L-�)�yf��:�'�Q�(��&M�BC8�$�D����)��w�5��5�&�,H�Z>+����)�"��w��D��xׂVVDȆB��HQ�iO�$�7T}#ڴbl�'q���A.�ȚFu'L4�v ��m���\����+=u�m%�i��v��Y4�1�t8)�����f�������s-�2�Mu�iB�6Zn�X<���T�Q�D�#�Ȇ�D��,[/xl@���=y_������>0��=��e���%f����K��6]�Y���~i���ŗ�CM�49v[mFd�Mc�C}lE/GZ���q��|��M��%��H`��_���}��q��W��V�{׷�����罥U��t�{��Y��������Uڮ������333��iUx��];��e<m\iǍ�v��1��c��|��>�dĽɪCv�L԰��hݱÂ��CZ��3l�4�Ff����QЭ�UMs6\�v�4�q�>��Zn�'T��+)�1�V�\���o������Z˝��`Ͳҭ����#��,fֶ�h<��6%�Fc�30��-xmh�=a��hFţe��=��@ z�>�'�Z����t�.I��;]3B\;`�XSge��i�L����9��}��=9��i(.z�1�t�d��FC:�0�t�l�撂�^$�E�����h�e�bX����r◍������[����+i�o��J��'H9�u�d�s�c%��:�lu�<X���M)2���n��6��}q���x"�C
Ec����Дm�4�vZ�Z���"}��?Ebɏf���V�Vv����V�+�����Ɯz��n>~~x�l�~>=>>=:;/Y�|���@�XA��_J���ƣJv�h���f�V,St�SV1��\���R��Iі[�ZَF�_���>t?m���ݔڪr�m�p��_� d�u2q0�3~Y*P����=ӁË�|f�!�}�N|l�xu��4��Q�ɻ&�ǌ�ҒѼe^��o^�&��2}S�^Ux�}��0\,D���c2t�A�c)Ƈ�:��]��
�gtc�T�z�Z��i�Í��8���n1���X��c�o���զ9�jBHI���#��7~�1=��� �FJN(�p�]�q)�.��%��2[�X#��Ѱ�6	�����~�Z��IE�Z����vr$e%rM�lGv��j���é
�N�4t�&�%��cy�톛�\&�#�vn�ŋL'�s�%%Ä<>�aߠ�8K�"L�s������Zخ�w��K��L�>�J]��[a��М����)Ee);n+�cӏ�1Í��8��n>zǏ����|�>v�y����eK��N�$�����p�&����q��!�W��K�"v%(9�L�	�ۦ䛦�����)/W(�ܽ�B�84��8�.����3���N8�R=8���LH0���,�x���gD��n��I%e��S�&�l���$a�v@��a�z@�e:ؓ�U��;#�q�Ē.���4B�!b�d�f����!Fpe.:��K�ѽO_�x���Ɯv۶ݽ~~x�Lz�>c;x߈�ϛ任ӭq~���A㋖	!�V҂P��j��rWqk^�Sޤ�/���E���ASօS^*I�%�(0�\��h�Y3�Ne���:1$�K���,c� �ԛ�·�	�X�WH���q�'��݁�X����� �@$#��k�HM�,%Ɨ��U��&׀�E�ш0���}=�����t��c��=.�J�!��!a�j).��a��	�$$$&$N�Md�s�-%��K�O<l������謴��7�}�$Dfn	�E)��'��9!�8�G��f&/E�W����{ܪ��$�
W&{2v���&z�[�H2ÙII<QL3M�fS��	��gY���:�쨖ֿG�}	��\��PU�2�b�%!��,b�!6�3�6x��n/�n�zӧ6�4��6���<c�c1���s�;�R��֬op���HI	 @s!��P��;ˁ�&���4u(ۆ�l/�S#��K%``�v��ޅ->�k6�-jm�ܘ��]K+W]�ƕ���W"���)ԅ6L=:���p˗��6��rBm.�IV<�.B�;���JS��C^j��3kK[؊��M����%��,�B��ݭ��l���>�:��\=�-4PB��s��@��<�xh���CN�a�M�X�#%�ɒ�v^���h��%.
i:҉�'
8��j�N<m�nߞ�<c�c0|<4tS�����Ъ	 �	 "%�6Y)vĝsJ���r�I�!��6�C��%�jT`v�m����$ɇoK�8�p�v���2f���7����%�ҏa4d�0�i
H�6D��F��h�L�~O������zY!q�L(��$��$0����8�,"o���s�n�\J���C$jz՜-�KZ*�
��(XƲH\�V����J��fj ����zY>Foy����v����!WGb7��aF�K3[(�lw6�$l	����?O�@�y�!-�)�ƥ�ӑ+J���kq{Ka�Yl���,n��|�bM4�Bʑ3iK���-l%�&ea�mt�ͺ5-�h5#1#e��Y{Z�B�ث���)�s�M��u��x�l�b�ce ZhRi�KRWix�esGZ��e� �Һ�����HUM&��A�,���i,��J���8K�QiE^�{�p�\0Dîn��7�K���¡3̘n�i�	o�InYq,X�I�L�]6���|�-b�nz�8ڸӎ�cn�??<~c׌c�1�ǯ5$��wPuct������N��5dG.�Cu�݂DJ���!h�"��#Pm�$I�*%�9�1AxELބbeC52 t�d�pNl�0S"ƹ�����J�T0505(�N����u�:���PR�EnrUQL��o�4�JaEși�m.����C	����U��y�g���i|+�[z�o��Y*#n�e�}��w������lj�c�D�YՊ�6�L@�n�Ѳ�`���j�=R���n�L��`S����K:xX<]������d�djp
u�Ƚ���8h��]|@0y;d�^������������L�;3s)�)����nM���GWq�o�x���c�l`��|<4t`�G�W
%W]��B����CY���2�y_j�����mK)t����w��̡[��^,g����x!b��	a��M>z�_xU#t1��4@���[k0�VcMձ�k��R:l[��HI	 C��x9Q����/��+�76B/oz����"�3kPm�;D�MM�����.�``����4�N��)�!�3̺
_|G��I$�T2�):���b餠�[��$�I��e�Pd��$�4I	%ݵI��l�$(�X�d�J��'����I]0�v�v��b���-˗V�/8i�E�_ٞ�uM05�
���*��<K��2�:�z\�`�Ĥ���Ԍ�rH�⋘�!Ɯv۶�<c��z�|�>x��_'OA���Xn�Y����HI	 CJ*�xn S��������!䤷}%UHJ��8G�fӵ4\���Y:](���d9u��1o�#�k��U�W�V-W�jx����e��>�~�O�c|V�Cïs�N��|\���>�v�KjVYl����^�$s5�&���qc�]�r�S��p�t���I!���(*���!���,�;D���3;%J<BI%��K�#�Y�4h��6~�4x�pN(A0�)�1���1�g��(�"A6""&	e"A6%��hL,���4AA��"QF�2&�Љ��u�&	�`�&	�`�tD�ĳ��DM���"X� &	
B'<c�1�|�g��>t���vھ|�"lN��p�� �8"!ba�c'D��0NԚd�(J ���%��(�A�F�GJ,�çN��%�4x4��� �~�@� x�v.חp\#�D��5��N�"��D�7Uē*f������h���(kZ �I*�f���q��J⇉��﹀��o}�0���s�Y�����PB٫^�*ch��VbH<�h��
��TB��9��Ωo j:��%��?1;zx��Ԏgwn8�e)�hb����&a�j�h&�v<��!��
����3���;3��Z����m��N�7�7u�g�+�����R��Wj�vo~߫3332��UW��WN��{�3332��UW��U�����3333�誯Uҫ�(���٢+rY�ͼx�<c�c1��=}�=ֶֶ�l}9�I	!$3��oj�@�<�Ȱ�Q�(l���2��H��@�ץ������#�DQ����.o�@��	������!� }7?|�+�Y�{�p{z�=�V��yh�{32�0җem�u4�.M�f���;���a�3�%:c`�=Is$$L8CFb�]���t�9���)2���a;V�����Gi��;T��Ī��y����޼J%��y���]�6�l�6Ƙ��j�\���6ǏX�zǇǧ�ǧg���� %`�da_l%QUEU�&��4IP�&Cq��&�����$�RH�R0R��	RG�݄ܖ�2)��T����Z�r��qt�K���*2VM�ѻ�׭�&���nC��$�M9w�ˮ�M&�����Q9j�*ҥ�b/tO%���H�1ꞫU�j�k[	F��])�_���L&^��c��t�ּ�����r�co1�<x�ŞǄ�	�*���sG7�\)���%KB��a��1�s��~�ZUM�`�lav�ƷM���4�j�t�Z����يV�,�:%�5ݥΈ;K������a�,�[��V�~O׈'��~o��bCc ǜ ��Zȥ��LB4e��J��B$c�ЈK���c��͗t�Q��x\�<�8{�a��ɚ~L�UT�N��c��`��)sf̓a<Q�&����d�b@�s����&a*�%����Itт�A��{�[Q��R�ut��Xz~�Y�~>��x3���]��䈗�4G�_OW�����Ж�4�֖[B��T�JM&S�Amz�a�ӸӨ��g��漷Í��r��z��`�~<a㧄��,ϩ�ꪲM�X�o��$�����s�ó��K���0�K�*�H;&Ӹ�e{���6�<�<m���0]3�(�@����3��h��yh��Ū�`�jF�E��)��ct�x�r!xl��
�5�&*��z{�V��֝'n҇�J'�%�@���Hp���̵�*쇱�;�'�O�=�k�c7c�̒'�e���Gr�t�K�ap���&3 K�N٥ͻRT+5'�)���k�.�&
L;4�=�R�2V��\���~m�l~z����X폘���ν�O�w���ֿ��H$�H����c��);�^��Q%J�%<k)!PN�_rC��NM%�L�N
��M���KK	�G����(�d��vkmfm�&��ΰ�������a>t�l]-\�5kY(�xq�t���l��ٳ���!����UYϮ�������Y �Xh�g3����w��=�������++)J"h8~2>����|�-���ƹo����Oş�x��<xK0�+�I�u��R�ɽ:ۦߒ6m�~6BHI	 h�x{�5!7$�V�&0I�X#&�4�,�����́���F-��7D����֟����]I�wK�7���'���S�JL�nѓ>�f��ibKj���x��f����g��O�!b�.^��r��ˀ���ξ�2��aЇ����&C�B9��B~��+�Y,�Y��>��;&@���N�㱑8l�W�r�.�-��z����=c�>c<{2�dHŦ�LB^)�B�)��H��!�tz�Y��ǆ���c��!��n~9
�8�
)M<�q��o�Ǝ��ר���R�o{����T�M�Wa\%z�"��%\���d��[{aء7-?p� �o�g�eE�1MjJv����25��k*�TX�&�����O�9�MӁ�J�X=���*T��`]��<�乤�忙0�u:@6�^��`�F��N.Ol�nC)p�a�>!���4K�ץ�<�	ڒGƓ�٠4�2��!g�f�g[�p��wA|�6d�ѐ�q��Q�*�e��d�;�)3�O���G�����Tx�i<�0a�efM���W����ba��ǌ<x�<xK0�*N���Rv[	!$$����a�{���$����&���f#$�
]���e(��gFrs�IV�X�g+��[A4垁h�3�N2Ӵ�X�q���C�R��4�ۮ�Hs�!�R0�	(�/Ll@�g5�m(�mXkKV��e��0K)`�����[˛-�}�t�{k�&4|�{Cc��4�+d��`.D���$��ݺ.��I��05�T{�OP�V#�y�xu���Q^gBp��.��M&�
vS����g�x�bx�a����4UQUEUbd�ٲJ��0auٜ�]H�8a:�P�ۣ����{f����i�&�P�i8ܷS1�2kWM�\�����U��!8T�su��&��IkT��bu4䃈u���L�'�4�N7KK���]8{����/*�`��G��f9R���*�1'X}��sJp�4t7�}�\��ѩ��i_���ƕƸ�6�Ǭz����G��������> D��5���1Z�q�I� ��'y��E"����8��N�W%��]L��rp*��Y����0`�����"hB- 3Y�t��v2C�?�y�H9��S�i�<K��HI���8^U����\<\�}Sf&
��$����Ӈ���\&ŧ�����zT*U�t>¾蟾����|�.�l�K�=��S�N��v�����e�m��!�K�6x��gD���,飂p�B �!��
�V4��.�qӧ�"A�"&	҄ ��,J0DD��pN(�� � �%hЉ�4"pD��L!�ab&	�`�&��nĳ��(D؈���P�aBQ�4"'DK<a���g�:x٢���"lDKE� �D؈���(�,N����0�(J# ��%�C!��	B&��&�萳�N�:"`�(C�>(�ɹ52Ɖc�D�d$����7F�PG�K�Z��f�H%��Yi:B�Y��~�f-2�B�j�LS9m���1IE4�⫰Ixݿ�ׯ��e��m����e�W#P�x�\3�*x�0�K,E,u��HD�큵(E�μj�Ț �IRu�@�rC�۶��k(�]B��z�g�Ԅ�-V�
mt�*N�X!���5[p۵��|�������㤫Q ��D$����zr�����]o�`���2�(e�!�	s5�bm���K�fEMi���e�J�B��	Y5N��9����@�k����� d��B*^Ʌ2B�-��-��R��A�4�0�a\��p�RФ�J�/J�Wv�v0��L�g5y|�6)�L4�Z,9d��	�����ؘ�4�9�:�����-�^ز�l��'�98Fʾ&�S��3d&(A��H0(���l�22\��/׵���ݬ�q���άH��ڄ�-n���;��*l�g��F�}T�[SM��}��M��/R��H��[[.f���x�#�6Y�� ��VA�~����u�am4k�s�-%S[����s�(i�)�}﯉:�H��K
�U餌4��s�{K��oK�WBش4���>̘Hm��&	���T���Y�!$6M��Wڢ��e���=�����UW��U�����3333�誯Uҫ��{|ffff{=UmiU߹�s�3333=��������t�E�6(�͚,����Ǭc��c�_��ә��ӄ�F���ֽ\��n�b�n�s5�1�ٲ�����
T֔j;���	oQ���-���X�(�m{K�	Z����m	���	x�����+�a�GR��=.�&��a\�\�:���-6�lՈgJ�`�X�֙�m��<�0Q��jiB�JZ�[cLP�IU�$��BHI	 ]U�a���L�b�8-��n��@a��T�4�([
R����e�%:a�2�,E����i8z��)��`���^�̺ɂ�c��,LQ�#����m��;���hդ
CXSr����۰�B���e=ԺX/Fa׾��0������K-����=��\�3dtl�l�[�8��2�[�w�$Ԝ�m8�zӦ�8Ҹ�n�~q�X�����8t��F�a��GF*����\�%&���);y�Qʒ���]4��}�)Ɨ7#�#��j=)�I9��FM<i,X# �Bp�͚M'Ėd*�dK�m��Ȗ(9��`���ˁ� �R@�����*���)E.��]%6*HQ`�х�Y$��]�}|�4�i&y	����Ӷ~z�N�xq�q�ݶ����1�X�O���������]i����բ�0��xi眕���ip������4������pm9�;��C9��w��!^)�����)~�n���ݗ���#!�Xu����h0�IF�SZ4�Ʉ�sno~��`�㉗�a�x{�$dC��.FϤ����G�|�i<��UF-��ss���xtn���<)��J㍽m�~|����t��|��=U��R֕ؗ�EP�y��ޜ�����n�N��I!!w�G�8y�>�ˇ�a�x��F1���F�%�6��P�$�6�:���u"�*M�]�wޝ���P������9P�*5S/�M'^�:6ܖ	�Ρ$�"j��7���M&얢Fii2L8Vp[���NOO$�I#�v��L�|�m�'Kvq�q��6�Ǐϝ�~c�1������}_<)��rH�6�FT��>�nL�v��A�R���������E��da��$J�4Z� &�HJ�M�ML��z�B�D�`�ֱq��K�
k/C9�2�dԮ���g㈢��U)ͅ]�U�ݿ���Xr������&��8K������cd�r5G�r��xnC�xuV�yV�e[�^��t������~à�Nu�I:��ٲ��p�Op�/����$K�&-*����$&�2��s�t<p��Æ���)=��s��M���Ʀ���M�R� �q,���v,n�ˮ��9�A%J�l�JlP�Ѡ�cX��*:	Ǿ�4��gWm�n�|����0�ǎ	��Y��;/{��3u��Iujզ6��~y�����tiP��lc��w���I�h�%l�vQ�K%���N�d�=�G�Z�d��$��O�4�i6i0X8j�vX��|=Fx��[4�P�T�FZ-Q�\�X��LlX�����Ӯ�be���_76K%�LZֵ֒�Ug��q��\UN����M)�O|��o�Ǭc��c�[�ֳ���٭�"�(w�g^w�²+ke�i8og�p�x}�)�sp�g�'ֲ�Y^�$��؞ap�>ì:��4��ov�~��e�G�.��]I�t���YFf�:�=�O��i���ɝU�Z׆M%݆W���Ѫ*(Ƀ��:(���
#�(�l4R�����Yd�]����t5*I
��"M&n#!���6B�,����	�H;Au(�֨M�p�!�q�!\�!��?UT�*20���zh�׆)���;�F����Se^2X.�92t�c!v��z��>|���z�8��|��d�v��CX�DQE9�HHp�:}
kAd�G$��̲����;��7g�T����b�d��f�
A]��C"�{�@���0�i�۝�'3|��L�x���Tv^�$��s)���&D�p�&�ۯI)�JCi��d�Mp=5�}}ڨ��RՇ�L'�t�t:p��.ܽ�޿Ll������o�4�8�|��v�1���1�ǯu�U�vs}����eB8̏1q�0&o'�K�C�+j���tŚ��'�����O�K=SV�E�\��?X�-�8֣d���R���B�34���}G��a[����F��P��N4yǟ��(uΈ{�v�5&m,��-#��6`��i�hV9a���
��уK�%ɧ�vg)M��g���=���QGO9�a�L`$�l�j���2�G3�q"��AΙ���`\�fo�?>�����2C��?>���h����[�� ��`n�6;G�����s��ÇyOC�Ӫ;���~�Z�L�2d�s���_���GWm�ox����=c|�>x�y-_�Z����.��Hd"Yu�$�$�p�ɔ���L>�����=��Q4��2<3���5��8k�<'5^��g;��������1'�.�6��Ks��řT%A�D�V�	$@'6�ڬ�K 숕M�>�1����r��~�UJ�UWd郧^�ޝ��^���[�M�USg��.S/C|,i���t����z��|�>xӦ:m�a������a�*�X�p��g�<h���"'DL�"%���L(D�,���0MAD���4CL��4"pD�d�,C�0L�0L0�	g4"h�f��%�A(�h؈�:`��'ؖpN�8ɳ�<C<p��0D��"5"#��4`�,N��6a�6CY%	BQ�O�A,����%�H�Н�,�ӂ&	� B�V�⬜nd���y�~>/��O�����g;���7�*#�ZkI�pwT!\�������
Kvu�����g�y�����'�-75�t��M"�[������O8e�ff?�UmiU����3333=�UU��W{���������UV֕]�{��3333�EUW���K4Y�a��l٢�l�ǎ�>><>>4������r}=��ȒYOBBB@�0Ѵ����
��~.�6h��>+�2�����l�����h�Чoz`0�(�v�z�%�X�!1����ԕ��ΚggCKե��{��������9�4�h{/m�e�$�g���g%�U/�4h+m΍���R��J.m<�.1�q�c��̧j2fn���J��i�{�t�mX��[x�m�q�q�ߛc������t|>}~�R6����{I&H�e0{2F^�UOU�6�O&�'93�Gs��ޒu�y4`�K�ԕ��,^��r����Y�}�@�:9��p�Ny���S�a�O���g�E�D�8?��;��f��b�^������-7<kױ���4G<��(�g�:�Tm����|�dw>y�w7��q�n6��J㍻m㏘��c�1������g���RU)A?����TJwq�Df� ��@̪%��kqɮЄv��JW_z3�����2��k2T@���d��R�BQ���|��K+
z�����>��y�)���h]!�E����m��/ɽ=6��]���e��^��%�mn�YvƄÖ�fsy-�͒�.�5���zi�O;%&����Y.�
�l�ƚ�Pe8�6C|0x�{Õ*щ�E�_^Ε�g�������6�����w�	���],�湊*�i#)��*.y��n�iN������?~����cDs]+<��+q���I-W}c�̕�4t�d��Kx���<z�Ӎ+�6�޸�������z|t|zvxIgv2��k9�UC��=v��ϝ�8�qI&`I�;������ivu-rF��2��HHIs��s���Һ�9Dڕj� �V̉b&<����rfI��`Bk��1v�t�Q	��[��ז:�Y2"ҏ��%�$�ԣ�\��4a4�n�=�D*�Аۧ)������&��̵wT�-kK74e%7X��㰂,g0���;]K��w�ɧY2��{EUJ�J�e������98�24f3�U�����}Ӷ�xq�q��6�Ǐ	��0��<p�aY>�f�5W�UO����ta�k∪'#:�2�F�ϰ�#,�5�n���B���w�>�/���+#�iCA�Svk�E���+�'߰�w���v�'�#�{���4BC.S~7$4j٢��zZ���d��%��>�l냧��;��j�U�y�N�=Mw�^��6�z$a�vxw���}?a��Xi�O�[tq�q�޶�����l|Ǭc�>=;<>�Z��x����{��Y���79�3O)�$c:_ۦ�H��5�BZ��*��n����cI��Hu-Ǆ6�OJ*�$�na��g�c��9��8{��#>(p�p����$���g޻$|>=;��fvQ}�ë!,�0o4>!� ^>g2gx ���q�o4�8���8����������G~'��t%�(��%yhhz�l��$�ɭ�� �EKvJ3
�F�!5&�E���H��=.�-�}�K�a�v�y����F0��[JPRbӘ[ZVi���*���&�cpXN!a��*4��US���zce�5�7�漚���{���Uc\셷О�v�ll+E�Nd?��\�Y�g?|�{���rK
4BHl�"a�ͦ\�3�0��UR�6�i2G)I��;��Diڊ�㊋��,Nɇ�{�ÇX@!�n(����=��ݫ���y��h�q����F�U$�:�K%K����e4>�YOs�t��-�gW���m���N�u*�NO�g��m�ƕ�co\~c�>x��|�cgM�KԒI8K퐤Ӧ'�x����'�:�-���O�pG�RB5v�p�X��L&�H28,M�L�9/R�B2��yZ�̒�)�{�+�}���"6Kh�<�9��>�F��s������#q"�E���Y�j�v�P��;8u�<�ɜ<�>���-%UV/{ު�B/�4u!��e�K�ŎCWR2&�pC!��4t6Q�4Y�͉��t�"xO�x|xx��B�M�v�UUNd��Ę�*G�]d��gG�ì�����y�������ও�7p�
S��>Tp��$�I�`��ܴ�3bԭ.�iV�2�^�9�gd�C�}(��*���s!�p���.�2t�r�P�^-�؝2�˳n�X�QNJ3���TGgn�����gWm�o�x��t��H��x·53U��z���H]�^OpѣI��Q�ܾq��P��]ʂ>�B���a����Kh��Gѧv�/�UyOO�vح�*���He��K&1��I�椆̛�t�K�M���nkd���$�+E���N�6��Z(�i�p�1�cO2�}�˔�4����~��@�/��rH0��'�$$	$$

�Q�������ɰ�1��,#����6ھ4h��D:TDI�c����sq�S�77�#�D*�UI*�(�[H�UUR�*��(UU,U�U��UT�KUUUb��B�U*�R��X��Qb�B�b�UK�V*��b�UB�UU,UR��IT�X�U��*J����UX�Xr��,UR��*���J���R�T*�R�eB�e*�)T,�T�K,R�YT�����K)UX�YRYP�,�T���BmR�R�i4�B�e*��)R�R��R����������R�YR�YJ�YJ��U)b�T��*X��B��b�Rņ�&�X���P�,T�YB�,R�R�*X�Rʅ*X�QeD��h��eIjRʲ�T,����T�U(�E�*�T���)R�)P�R�e,P�K���*�b�T,�U,�UK*U"�UT�4���R�YH�Rʔ�X��P�K*UBʔ�b�R,T�K*E��E�*�T,QeP��E���iE��E�Q-�,�TKDYI,TK�(�#H������%%%%%�������&��E%�J�J�J),JJ���%E%iH�)*R�I�Y)*RYIR��K
K(䇇
J8��8���P�i��),RT����)(��Ie%(�#P������J��RXRY))Ie�i),��))Ib��%�),)*Q�F�%��),�J��)*RYIJ5H�IR��%JJ���RT����47H�)))))*JJJJ�K"��)*)*,5R4JJ�J�%E%IIQId��"��%M�n����%JJJJ�
J���Id�T�!aB��(�T(�EIEB�iCHQb(�QH��Qb(�Qd�*R,Z�UR�4��(�EH��E�E�(�QP��Y"�R*T*X�,��
�"�IR��T�*E�R�R�LRX0X0X1B
A0X0X0X0H0`��EK%J�"ȩQRĩP�RT�*TT��EK"��IR��EJ��**Y,�)*E�-J�,T�%�(�QR�H��QR�K$�Q,$$���H$�i*X�QR��EJ��T���H0`�0`��jQR�"�UT��Rʕ*T��(�QR��"ȩEJ)*T�,�EJ��T��EJ*TT��EK"�(�EJ"ĩEK*TT���R��*QR��QRĩEJ��T��dT��EJJ�EK$�EJJ�T��dT��EJ��EJ��EJ��T�R��,��T�*QR��T�T�*T*TT�J�"�R��QR�R�JJ�**RT�R*T�*RT�T�*TT��EJ��IP�RA���(A�**,�R*)*T*T��*Y
�"�B�IR�T��J�K$T�T��*�R�Rȥ�H�)IJE*)d)IJ�))P�IH�)E))IK$�%,)R�)QH�)QJJY
T��)aJ�X)IH��%,JTR�,)bR����Y%))dR��E,�T���%))IJJXR��%,�*JT�JR�R�)QJ)IK(R����*KR*)IK$��R�����R�)QH�)P�
XR��K)R�)H�P����)d��)P���
T)P�P���IJ�,JX�T)d�T)a))R)P��)Q)P�"�
Y"�)
T�Y"�"��XJR)IK$���H�%,��)dR��
P���E"�����
XR�R�J�)d)��,)e))dS�D�QJ��%"�R�����E,��R��E),Bȥ�J�XR��������e*�R�*)b�%,R��d�E*)d��J)b��J�E�R�JJY��%,��J�TR,���IK���J�Y)aH���)b��J�T���E(���JTRȥ���)dR�X�E*)IJ)QJJE�K�R�*)E(�E,��)E*)QJ)QK)dR��Q�oij����R�X���R�JJT��%,���Rĥ�YK��Ѣ�T�,QT�YKJ��бJ����T�,QT�,Q*�Ib�EQ,�QTX�R���T�)TU"�r�QT�EQb�e*����bn�E�Ҋ��UE�U"��J�Qb�H�YER��ER�)T�K�*��J����UX�*�KT����(���UUX�T�K�UYUUB��U*�R��X�UU�UU �X���'���q��>�L<iZ)Jr�O���AI$ A�QI@1��_$�?����޾��������R��~��~#����}aO�����+���K�p?8�`Y�A�r���<�C/A��������C�>/k�O��x.��,|���r��g���,��(>g.��h(� ������W����@_������(����?�"������(���G��.�Q���0�?�J����'����B��~�?ٍ���!��O���Pa�S��A���0�"P}F�,?vh�Z����3���i �Ȗb�$�?���))?�4IxSB�ߜ��}�����F����e��^�! ��m�描�R]�CD�/
�QCQ�H�O���A kI�)bC�j�DE�B����4�I�,�'<6��%7&�v�Ԛ٩����ύ�W�\��O���H �@! P�ET"D�D�����h�H���I� ��T��ERHK���<?0��D���C?0~g�*@��u����!�� e���?���?p�o���7�~Ϲ?�
�* Y?�a��}ڏ�2k�����_�~`6A����������� ~2?��?���~��� n?�H������~�����|��/��9�F��O��EP�C��g�~����~����A����~���#��)D ��P ?/���R+���?���iA-e?`0����6�p�xװ���X ёށ�)8F���	f~�����$ @)JJ���)7t�vM��53ᦃ#A)(b�)
�E�����9Cxi��A�A�`u���7 �`I��pO�E@
S@���J?�����|�	�i�@T �Bߘ��  ~��ߗ���{}��������[���6�_��$���'�Z�~�S�h�~�������Ik�K'� ���������ջ��* |ϕ��PV���@C����G�(
��2~ݟ�<�����>A��>�~/�&��P�?V�4�"�>�ϟ�o� ��r��.3�#`��~t.����?�;�`�p~|���e3�.60����8P 2?�O���%���_�����J \<0��~��7��i�vH'�	�d���[���Թ�|/Ђ��+�?��F��s��ˡ�}���P~�����t.�����?�h(��r�?���	#֔#e��^�����.�p� �׎