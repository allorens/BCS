BZh91AY&SYК�d�8߀@qc����� ����bB��     ��mY�D�j�A�YD�4Q�[5�e�1�QUIQJ��$��m�F��[f̕����*BE(J��d4�P2��6�U���
�M�j�&j*V�f��[V�fKj�I���klb�SfҫUl`�a*Y��&��6K[&�EI��U������� ���m�S6١j�Cjʊ�$k�ج��ȥ����R��Z�-��օ���U��3&*�F��FƩm�X�eRcY�kb��Vա�ⵤ%I3    ��o�v��n99X[W;
�`�r�u�U�M�U��:;�[u��p���un�!��V��Gu�ֻ��H����Ф��R��m�V�m[p    �nT�w38
P�p�: n���Pn�ph( \uΆ� S�t K )@v�wC@����*Օ�6�ZMM[�  v'x wR�  z2��ݵ +4��� �{��<��4�5�ޏ@ �i��  ��
*�<y� =��{ހ��5-����i2Klٴ��� ws��@����OI���@�0]���^�� נ�\��OB��7��@� p�w� �E������ڕM����b��̭����[e� d� ^�p@�n�P
wG
 ����q�44���-u�@ P�vݶP 7 �P���m�T��Z4�ĕ5�!M�� ׃��Ӝ  �Vp�m��Û�i@3�����]F��
;aۑp� ���@ 	��Glm��  4mR��҆T�Z�k	7�  ݆���vU��45������Ν( �8�  t3v���r0�lt�u�"��X
 6���@ڕحMY5�-[I���[-�  �^�����'\  �X �0 ���\�G���QuӀ N�  �F �4�05��Ij45Z�&��  ���  �sp �P 賵��s�ێ��s]\P #�  -:� �g[� S���G�W���c!��(Щ��M� � �F  o8� w� �8 ��P��  ,vp ��� lLPP�    }   L�%J�@  � "��F)JR� !�фɀM2b E?!)TH      �~%)T� &��0&	��L5Oz��iT�G�z&�@��dh BT��E #&�M2j4�C@hơ���Fͺ�캼�l����m(��J�
�wŞ'���%׬�r��R��_}�UU}��H��" "��  *�O�>�"�
����� �����?�����a���PV��Uz�N�����?� E|}g���?	���L��ȝ2�vE��	�?F ����~��a0�� vd0��'L/G���� �x��(�dN2�S�#�� �8ʜeOO�D�x�<d0�G�)�� q�x�<d^0�vQ� �x����x�<`0����A���3 �x`N2'C���P�q������L	�C����"q�8�aN0��`	�8dN2'���D�q�8��8ș�8��aN2'���@�q�8�`2L���(q�8�e2�S���� �d0����q�8�a0�G����xȜeN2���q�x�<`}��d\�<a0G���x�x`2�� q�;����C�EG2<` xȪw`U8�(�T��US��'v�(��PW� 2�� ^2�<a@x�
q��"�DN2��`U8¢q��
��T�()�S�"'L#�G��2<dx�a {����N2'�A����� �dxȀ�� )�@S� �N2(<dT�Ƞq�Q�*� ��#�T�"q�8��� �8dN��P�"q��W�	�D�q�8��e0��T��`N2�S�	�D�q�8�a2d&@�(q�8�a0�e8��aN0��A�)��=y�z���[���T���3HΧtkt��1KS]�b�n�O]��ExAö2��x6a�����X�GY!�6���mE���l�B*#6P��sqDk4ʷ�b��$T�h�Ő�KRgh�z$;u؝2�Yڵ����9��7���V:X�n��XN���,2�yM�����1��D�Sz`��UA��7(�k�t�b��1䱇Z�`�������H�{�*�<� 0�px��B��;Tw6�z)\r�ݕ]�F�z������U����KB#M2�jN�[w)*�]�	�	]˽ƴe\ۇ]�ے�.4R�ƛ��,�֩�;Em�$�1v�ݬ�����̫{��@���Q{�d�vW ݡ*۬�X�Д,�+���������1�32�ɬ8�st�g6�+�ft1�F������I���Sc��%��H���ӘR�^��m�%A&,�*U)RT�����:n��.)�I\Lؤ)au�����rf:�lP����4�b\a�nk�$�ӺtU�۹q���LR��TkkQ�B��Vl�l�q���e��(�v7BaLf09�ff�rS������8�<�H56�nS��I��.g�-TZG�V�@�;)�I�[��ߒ����L��Kܦݒܩ��sA*V����[�Hu*���	��f����Z'n֠U�w��x�Њ��y)\z�#`��כ��޲�Ssn�YV�*�!���l�T��f:n��0DxT��u-e��Uy��&CD�����X[�ܝ��^�%�D��ݺ��3m�$�t�M��(�D^�������zVl�=�z�cb�7�
2�K�7��n'eɌ��rj�z��U��\�!Ȗ:���٫-nl���Pbcr��*Ƥ��e�D�W�*X���wNӗ7Vk�z�Uc*�f�	�{n��G$dui˂aŻQ�ܠ�j"]�w.�C9�Aސ���N���u�{zV+l�p�l���j���ȍ�Փ�P��������.�dq�ԑFiWE�̂��$��Z�1�-[P#p,R*�ON+l�E��ٶ��3qf���28 ��ƈ��-R|�o~��(��M�z��t�e;����R ��Vɉlȯ�6�Cz�,�)�3�`v+�_}eU
՗k��ؔ���ʲ-�7��w4��WN�Ҫ�2�팠�l�ma�6�y-�/F�3�E�K�R�T��4�qېBdJ@%��gK�w���6�nad��� �Z̶��r��׋D	�?d�e�^�RY���U�j��m�KW�5o��D��ab�5w��[
�t��}wN�tr�i.jح��a�V��k�4ùP`;�3n'&�	#oM��X����,ЙF*N�5�7F��y/���e� v�x�r��.ۦҥMf5v�g��� 2����6�m4�0M$UZ��zs�H�@R�ik�Owfh��Ji��mn�)���`��R�{&�w)���2Bޗy�"['�-�I&��f[���.I�/1�e��'�2�@g�V�����V,#KJ`�)�|�������U�S`ë]9j7e��e
ӠӴ䵒P;-���l!x����2��r�X��"��:8֌/0�N�0�n�������Y��c^V�����ޜ�j��jɮ��bb��*K{R����+3ḿ;�{x�պ��W�؎�:v�#+8�
P��y-X��K]ͅ��*ՠpز�s2li�2���Yv!t�]m4�m;����u��T�&�pa��2�A�����[� ��n�����w[²�[���c� �a�p�[n�U˫������ʖt�܏~�f����l1�ub�=�� �o�؎|*֝#s9�ؖ}C`����f��gEړx�����{t�ݐ˙��'���jdзPLո��.��f��Ƕ[�Dm�b!�j7h�^�Z�l6�=ZpG�es#�^�B�e�Iˀ�Lgk3R�V�MlmEwI�J�cu45D]�͌^c���q��#ܴTC��ZV�wY�]a��ѥ7�Q�R��JRL�naqb�Fl��[Z-�ؐ��-�7��ViM�GU�Ӭ?U����X4�;{��J��B�4��nl���-����L��m��r�I�V�I�����#�o5�r�����C�܇Q���r��ݺ�����xs���,��&�;���%�h7�)���>S�!��,�ύ������+'N\���B �GI��f:8W2��&Z*�-���a�x�x4f�,T��EfPu����a�:�1M�$NTd��cXA�E�lr�ǹW7�[T��A��U��'(����0�V�����J
d�W΂9{�6��O�˂J�k7me�NMCRd`��G*�/k+5̖����Ȟ$���.�ܹ0ݦH�v� ѬN�E��2S/r�c�VՍ��̱K`j�jY��-�0����m�^+k���w�uݬ��.�:��\�m#�fm�ڴ�g��D���"�=���۔2�Y�J8ƇmTZ��V����nI���P��Z�Al3)R*��^k�.4 'i��F^�B�&�ix��YY����4�͸��$�"�SyY��9�5o�"�� ��I�XE"]�kD�AF��z��Cݩ�eV��׹XI�Y)휛7M6u���$b�ڬwW�l��b�c��<�2�Ξ��x2f	t ��˭@$�[k%Zb!���)�؁h�˙i��^T��z7[�u��(���n��I��x�Rʷ�fCK*�I�}������vI�g7f�5�3TE�]��*��c7ĠEKďJimnĶ�ek�4��P��:MnӬ5%��)kD�)ZF<�bk���ϑW)�����U��,ۙso@?��*�-ࡶc�&��Z�퉌�ݣ�'ق�X���Ȫaׅ���E��`��`ЙN=j�ܟ2N����\�%��@,�,��v��9���A�(Q�]5�&�%���I���IB3��W��Q�(���廱�ź�˛R�P�u��u4HX�w\�cse��a�+(�Ƥǌ��`�L[��a�;�@C�b1�NϋNMih;�u��eUB��x2V�ðQ�\�T�X�������HB��U$6�JZl2�3fc+U��eӉ�Y��aa�����u��m_�b�#�w�0%��L��-�a����{e��j@q�� �K�2�]�Φ�!���A�V�h&�CaŎ�C�m���"�]�|֞cEv2z���!�F��"������v��OUk+tr��y)����hz-�I�LY�f�K��,���-dj�jLM.Yx��E<��r�x4m<�� 4��o5���I�3m�$�0�ŉf��A�7+D�#���c����1G����FF��މ1�)��\d��o,�g�}f�<x��r�K��:�*��k-`7��&T��
f^bWA��&Sobm�[�ꛃt|lİ�e���.��Vbľ�2��Z���];�ϕe"oWP|yޓ���/r�Q���uc�V��d�un5�\#3c�?��J��~���]Զ+ҕ;�M�*U[�(7l�0�b�e��"Y-⥫Ჴi����Њ<;��橵V�#�H�Z#vt��m��FS�R�\��.ѦY�F�����+*��oe�V3��nl-c8��-�v��6�!h�	���j��	�쬰��n#�C��:e'Csi���2j8��4hѷ���.�E�sD�+z�aV��ꑒ�Qj���KA�T��չm�&��&�-׸o�w�<coC�P�J�@%�S�NA��]�O�%f�gf�F�C����h8�i�gZ�b�f �<�y�V3��*��Ǘ����j���l&�0^��^��Q���V�TA�r��(�w6���h�1C�^��-˕���z�#~��t�*e�6�J���Ee|0l�:Ǚ�4�Jx�����f�͊��)�u9��It���2��l�U�^�F=
R�T�۽!�v����+5�>g�)��u���sh[#P ɚ]��C�'c.��AՇ\��@���Ń3�'V!��5���BMi*@wH��S�f��̉H*�@�0�Z���b�[)��D�-�S5aa�#u�Kծ츦��֍5ӧ.ĵ��A��{R���u�[,\d�X��ˣL:X��d�×�x�hP�[��E�0ĪĨ��t6�����YǴ�nYvODmfh�Yd=44K�5�.�V�al�����5�%A{�r�ɛ�C��	�ݛ �\� �ڳ(��)l�4eM�MMˤ^�PEV�[�˖��I ߐ"V�2��xݰ�s��kF�.��y���j¹b�h�3rm�� �ggi�w&//WQ!��Rk[�Ad̽˦�%�r��N�cG-��+&U�ʈ������
|�2�BJr�D��Z�ف�âB�b��t���Y�R�F��mֹ��6]�B��i�eMr��r9-Iw�wQaN�Ǳ�ʷ�-��w�D e
B���n��.�o~Z5��k$����90����Nb�Ӛ���ǿ ��0�b'�ۦ3����q��%����E��e^����f,y�6em��(�5�]��$n��ܢn<����� �7WpPY�����e�d����k���'&f:X�������U�4i�$�z5f%�7z�=�[���i�UɂVPT�XZ��1�g�Ӥ���1%��L����f�Uq��+j��c���nT6��JB�6|i����$+zV'y{tk7���b�|"����c7sLhކ-�Sl]���q�ZR׉om�����]c;˲��㗶�;#��Y�c�HP��%��H=�EX�з��dm��m̘��-�\�%���Z��Q��[)�$��!I*��u�I����D�j��X���bei�䨉�*�m�`SSj���z[�䵂��[%���٘o37E��M�1k������e��S��n��d92�3eyy�p@��0挗���+.�1)*JǏ"�i j���A4l��v��6�:ƞ<�ͦVX��z���:	�U�ta1�ٱާR��5n����ӧF]�J��Ӭ��K�w6K�Q��/r��j�y,��	BQ���S(�(�2�.�����a���m*�g
[
"#�[�E7fօ��R02(2I���Q�ut2O&nf��NI.HB6T�$8�'C�q<!7H\ͭ��2��y�k���:�6�+�����Qի
[x�U�j6՗�伶[��#/kF<&n�d�*I��b�/P���c�c&3�0$�Ӯ�BȬ�Cg�h��owX!�f��(�R�)\Il�3F��i�"��Xm��	�ߎ�[7^�N�#+%�`RѮJϬ$���v1�.�^6 �:SJ��k7 �&U!Y�f�F��v�v6��B0�)�6E�q\Aַ���D9��5�֕n��3w.�t���A�w^�Pe�ewՐ�m���&-�t^�WJD����ю�cY��ӶQ����*x�+>,%{������YRѵ�^�(R�)L���CJe�kX��n��Dj,
���ZJ�I����e�'1������Z���θ9�К��#V�'������fR�@�-�)L�̓6�
f\��y{r�j*��f!X�	��)ֈC��Ee"���s.Ķ!�V蒋����E�NìwK�`�$�2������ne��g�Ȫ;r^h[e+a�)���͖��l�� P���h�/�<xy��umڧm�5bLL���F-�����l�d�ޜI���3B��[�'c~x�.��&�ٟj#���q�x"Vu��#2m�*CP�:Aq�c �fJ�uJe�MJ�"b��H?�ծ�]\|؋p]���j={��u&
�6�f��I�$2"���ͬ���X��k�0�w=m����7p`t���O�$r��ҭm`�Q�2�cN�;�1�fE2��q�Km�[F��qk8��5Ǔe֠�^-�����`vT����ӓ2)��J�������ӈM5�v�%��H�HoI�*�<�۲��m٨��(D����W�-s{�d��Y�G:[������;>��o�,�k���dU7+J�	���KՆfR�M��2B�6�%�3�PC*]H�A�kI��ͧzm�"���T��7�̋�{��3FF�b�Ӌ"w��D�����(�n�MǸ1�]F`�m�MBԒ�Y�s�Vᒯ#m��W�MCg7�W�ZJ��-׽��y>v�<��1�g�xz����
�&*�L�3:�G2�5&ݸ+1�a8��Zƽ̼Gjz1P�cNՉ��O.�"��j���I���p��5��k����c�]�\�4�wL��[e&�X��*�,�r�8��"���J�%�÷ϝn �"�ֶ�)Xtj��YF��*�Y�|�GDGX���N��(E�ش��.�4iw'��R��(��u1���8V�3e��ō5y*�a���)�:O0��J:����ZPu��*�������P�f֢���A.�%�6�S�ý��z��{��NI&�Vf��.N;L摥Õ���@�ʽшB�����2�x�j!g]ۺ]�v��f��6G����W#��՞G��,���� �KڷE=��`��I��#�ڰkSgI�:��\�D�6e�VBj�|�i�:�ݰf�X�$0�ʝM�2h�e�|ڳȈ�1A3dY@B�Ռ�t�B�{\���x�A�<͓���>���v��	3¸�1Ʉ���f��8/�%J�d���h� Ird'8��7��_wsh������Τw3�a ���cɚ���A��9s%1k�6@Pa��:�U��h�V���p5v�p�QM��&�V�L+':��J'l�-�D�.����U;�^���~�����{?�?��K}7�����0�O�?���vۯ�N*]p:�;o���c�L�P�L�T�[��f���M��X���XV��O��C`�7�0����+��1�s�=+��꺅�.封����{�ԫ��̏GT�6�6~�n�\P��fc/fX��z8��a�-Us$5[�������Je3s(��b�{���N='"��4!�h������D��+8\OF�Zu�gc�^j�}!���y�\�w.mJ�1���'���Z����aZ7qj�ZBuv+�Xpv�_g�n8�R�g/~�&K�}Vv>-.�\�r��CMu�R�:�]�%u�̪�5��{n]����n�C[�Qc���ʻ�,F��8�wڳ[��y{i��<{�%�U�[ y�cQݜ<�M��̝�S5��*iY�DqL��o]��A[�h�:�ˠ��n�w/MJ�.���jS��U�-^�Rqw+��\3��`a��n�����q˙w���v;΂�nT�m��G3.�ݔq��R�g	,�+�n�%�Ͳ��F�v�a�L}*֔5)�nQ�"W@�v�pa�t��y�w�),2��}J�:3��8$�ε�����喊�qf|�(�w]�I��Hk�C{��t*VPF�G�9�/���*�	��;�̚���5��7.��*j�5%�#�W�.��}��o�[�X�1.��CětZ���+s&H�:ӓ15/sC�������/D0x	Χ�OV�5ׄ�r[em���sdX;���x�.�i���n*r��ϡ��Ư�vB;",��yO3R�ʗ������)7Ivm񇢧f�/%ʺ��������&�!�Y�yN�;��	U��c�~�3NVLWlc�6�D!��&]��͹��Ϻ,�"�$w�,��fWm F>�ܩ�6>y8k����wwZ��!Ԩ���a֛R�����+�8d'�A:F0��([���Գ����
��&oJ�����A�v�6�%H��O���֯��r�.d�����F��Q@a|ün��f'�*쮇�c�iQ�V4Y�Ǥ�:�6xl�X�ݚI�c�_w/�ż3�r|-\��dʻ���x�Y	F\�{t�m�uZJWVj�3��Se_�������r�4���b���3��Et�W�I�v�	���vGJ�:o%��DfV;i��1�%S�u0�E������,X跍��b��)��r�5"5�ZO��3�p�4��̈Wa<b����\�f��u�]�����Ϩf
ʺ�/.[�5C��ɨ�/���L���w���[���z_DB�{L��b��ـ��b!�p�sb�'P�yVa��-�N �v���u^���$v0���]�*�CD9�K�y.�4@��sc5=�_IhU7�j�y��rGc�Ƃj��w\�m�y�A�@Ԯ{�5.�S]�ī�v��K!����ý��˗�E�4�׬X����U������I}���<ֱ�����F�*�YW��{��w.��r����#m�� ��y&����I��;w>٪�_t��/!��@V�&=�t���f��nt�,ڧ�V�A�»�B�{1��`���L��먤,��E�F�4��Ι�^mM'��c	�7MZ��[.=i"��u���\�g���ޚ>�����(�[�x��=��U����xs5��x�I2�%`���Ř���^(���ҨGi�0o��k�e�C�yOss���v�*gn;o��S:�C����%g*�}G��+ K!����i4c�ʺ!�-����8ӕN��3��3�W��,4v�6�ۂ���	�o3Ō�gP�:�oـ�I�H[ۘ�� ��ȕ��(^o'���T�Erˣ�c�a��8�H.�ܰ1[�	��>v����[v�S!���8D�y@����b�nU`�
��Ȑkf�u�5tfjw�g.!�o��I֭�U�0��>�oG��W0%@P�$ɱ6��_ҧhG��w����)f���c��k��
�B��oM�`��prGbˤ��U���q��ine�9}���u7j�G4�K�X�V����7y��1����f�6X�o&�j�emތ��!����3 ��
X�:I��s��;mm�=+b�k�@����=��ɔ�)ۖ)sS8G�9��>ld�����5P��鄒���b�s"9�L
焞�ma�y̛�!�˝�f�MCz��5�iF�Ûo@���l`���g����K�kU���G��V��Q�X̀��݅�[�&⠭Sr���X�9�a�r�T��X���lYY�!#l1��;:܁ru�q��*�=U'ب�b�ͼl�����Q�	Zsu�����:�Ӱq��[h�}�B�ka�`�Y@F�f�s�l|��}��u��q\��o��s�#:�X��O+����P�{��Q��9L �jn�u�tx掁]�#��\[�w� ��]�jR:�s\�C�+\YOE���h�Ν[�8s����Z�ɭDܧ���|;vy��LK���7�b�������ղr�ʮ��h�e�$�!��17[ԗ!����ʧZLܦ�wp���^�&'�"o�/6g2���WWn��Z�Q���wy��g��8��7u�X���L�o��n�p؁�Uc�K9mn�o:qs��2��7ER��������va��
��E�2M����M2룸�B�]�
$�}�ӫ����F�n�oBU[�� ����8t1|aۣ�0<��_&-�,�M��.���Ǌ���	�R�F�<�U�A�Jf��veu�[����i�/�,�weg,�� ��w:�ј,mN�6�C;�e,��Z+4r�m������'�׻�����e$���Ǉf�+2�1�gXo��:�$h�d��YL����n-cNd�빜0wI�=�e=�nv)wܱ�:/q+p��9�i!+U4���z�䢪�GS_Y],��9�)	ٮm�e��.��7Y�r�H��t9��>�7���5�}�n�F󅝹K8�[]�A�r�Fc^��B#Z���fs����ë9��R8t�'Ϝ��4�t�}dK� SN��l|k�2�Q� ��-c�Q�:���*�s��y�tv�+�wwgM/Q���XT�_;�%te��Y;�'K[���0R�fwoE�{�pN<����,;xj���3�G�k��Xo�K�s2���o4%f���X7Mk�k�j��*�OQ���t�O0���-����C��ޢ��A	��*��!+G]��+#�z��/NS�5�N�V�	e�L��:w;���4k�B&2n	tc��Ǳ�xR-��{�z\9N��5,���hT���GXqw
�3��ٴ!��!"���AټSy_'����>[A���b�o�]���_�t�o���l��]S(-�IH�����V��Cxe���Y%��$M#R��u
�"�5��P[���T�ᒛb�*����й[��Bf�� i�? M���(�ժr��iC�K�l:r�%�Pݵ{�zm�����=�8�2�������1�Yy��ջ(gJQ�E�Kg1�U>�ޜs��8�i�����i|.������
�,s;Ƃ�j^G�L4��^�|He�RɆ���p�9qT�f�^`݉�.����XD-��T(��n��ܭ��u��s8VGy����5�,�\��(By7��o��;,�c�ފC:��!g�ڱk��V����lΛXo�lr$)��m�:�*��^Ic#��Õ��W4we�OT	��D��F�Z˳pS�Oc��B���0��-k�y�r?�G��Q��F��X�����=�SL�\��z��2�p_	��Z�-K;G�äOTsvfޢP��k{�v ���k�m��Q鰶��C)��joV֚�������D,̏�D��xղyv���{��i�*��o[N|�8�o8��6�u���x&,u��P�"�Q�������CG'|��XA����	=��|�!߮�v�k$�ݽ}��-���y��<���$�z�c������c�>6i�|�sS��ƒ�K��B��tWCi����Z ��f(m�1m9��&�_f0���X�2``�Z��3Ep���F���bKT��A	}�c�B���jfi)�Z��U�wX���wl�Gt���)S�2�@�E�Mwm湺��u��Z���3��Q�z�T�PU�%z�6��"�6MՍJ����;]a��\i�pAJ�cF ��T����,�l�8h�Aa1!��c쳅���J�
������&ǻS�o�ٺɸ(�]�U}��w�1N%b�PyWQ��t�n��k�Uu�.7������q�
��Y����|;�P��s�-�j�{�k�%�V�ty�:��-H'�ժ�ٮ�4��$aosI-pE�\��.�^�%��y���i��v�f���xZ�%n�R\���)8�vⷷآ�C�4�f�%���������ь)3� :1�L�L���p�6�#�s�V����v'>�Z���EM��r�s���oguS�'�K�JUW{/�����3���;�0�>�O��.�Y��&]��`�J�̈́sE�N�5PHLSdCG`<\��Ɛ
仗OsM,R4)Y�Rr�*�\k�83>��y�Y�"Ӎ	J�.<�>�0*��㡘Wݙܮv�L�ˤ���:�־�Ye\!m�j��U�8��Ǎ�3%N�u�^)m%|qB�*[��h�U��u3�m�vE^�c�JA�rWTf��)����A�jC_�Ug�@�a���?4�xǫ�O̬�/��-u���.�ݼc�T���{���V��ȫ���kڝZܲZ��/N��:5 �垗�3�]�ڴ�.�G���+Z�^[3���C޲����Hn�t���ot���b�i�� -�*���ë��.�wv"0��[lhG'7-V&�9��x��WO�9��<�{�z�V�l.���Jp�G�3����]���y7M��K��W]���$-u�s3/Z�Wv��m����F�Z���4���Q�����9����_'��kep��yq����x��/`�:П�I��)��������Uvٔ�c���Ak�wH�G����~�2��t�b���^�Z�W3�1\��,���}���{�pM��x��ș��9��È�Q5U�ú"���L�Ξ(�۰������4l�ڕ	6<��ؔ�$LI �#�p�c�wK7���w0��y���2��a�(�n=���� ��}�gS�r���BE�t����X����Ġ�Rȼ1c��,;��[��CX��ba��h�KiM$N��lY��W	��ddO�W��#NfB��x��N���B�2pvR��\�F������ʋ/��,��쾡)����b�po5�D:.�}������o��{lQ2ͣ�f^n	�t$
���0�w|N�+盷�	 � O�5��Eˮ�o,��d1�/��\���Uut���I-���O�����l��EG�k�-�9��7�"}/S]z�u4���;�b��]�])5r����� ��tW�\�:��̻�� Ӕ���k�R�7���[��AvޅtSrc�W������ou��m�U�����6}jD��2N��|�җ��WB	�9�׺5C�v\��]HX뺕��H����S�"v��b���y�ժ��뎍w`���y̱E��a�K��#^�B�a��o�Y��⹃�g[V�����"T��;�v�%v�>�]��)(ir�c�9k�8[z&0��YrR�ܣ��6{N-nDyR��u�����qӪL<��Ƨ�+%n]7t�r��ua���-b��t�J�j(jR`�]Xf�Z��غ�_qԗ[(�Zc���=>����h��eq�5��1x��0�2)��c�a�lchmY�E�&��,t;�
��8ލ0��0���Z@�r�C��ȝq����;}ڊE�|lj�2���S���6����gR�U�i��P˫P��6�nYCpؙȇ|F�F�;'p�����Ri(v���uݿ`�ѫ�bJ�l�ə=0J��m�+�鶕�m�� �ʔ@�e�Z�r�D�-����PG���%usκ��B'R?.���M���j����H��t��9�����G���O+9n�/�7Tuc6�\�h�)Y�z����J�$��.�b}-}}���=ph��:kɏ��a˜HU��R��h�T8�pB^�Z����ν5��r,�}�y%]�v��MLvţ�+j[Fj�k1�k�C�G�5�7�Z�CG��Y�r�)��!Y/uzcc�6�]\���Ѻ�����C8�����2�&Y�E�O��w�p��^�S���+�N�OawR��K�O8FI��]�.# ���I�x�P호��[�9����b�t�V�t����Գ�sՊ�:1�K�rg21l����j�J�;�vv��rϡ��Pɏ+%���;�'���o���0��>��w̍��>�q3�ŷX���'P��P	@ �h�s��5,`�-��}%g]�u(n^� ���>=��N�Zh�!B�qɄ���1uR%s�ө��q�z�tQ{���
:T�=\������Y��@��5�6�7z�u�v��j�$+C�/�?|�n��8tx����z�z��hN����l=I��b����J�Ԟ�����u���kw��{G[�N���>#�g�<E4	w�u�:��GRw���
Ч���Ǟ����{�q�Ժ;�~�u�w�h�N����X��ڢ"��_�w��E@=�?�||x������U��������}��Z7vhL-X�^!L=5C�����*ȞpU�aԼ{Jn�w$ҫ���C���N�coZ���Eiպ���\��>�k��J	,曉;�C�P��y�����)��5yg��{F[`���6a�1vzo�g7���/$f!���]m�y�r�-�xmq�Q�3a��%�M]�r���ۏLjY����yu�! iPYC&⽲L�e�7�J��bȫ������ӹT�C)��ͮX)b�o@��f�m�o����Yz�p!q���X1�~ǘ��5�i}·�wҳB�3��@{v/kF�1J� ��C2�XFٮ��@t�Ԇ$���>۫�nE���f��t��+�{�+[sl���.U>V���(4P�Iu��Y�u� %U�wճ7y`4��I��d�,��YTu�� ���_۱�{BVPA�;z
ĭ�0�T#12���[��+]Z�������nWP�� E]��6��)B�$2;t��m>ݹ2�,���`�U�	;b�j��+n���)��E�T�*k馺%�/��q��$�Y-^۵�M�oP�tl5�V����1�Y��ΪAv�pބ��&��H3D�;�ee<pH��!�u��*ޘ%�]IF�	k�:M������w�+��b�6�vՋ5�e]\�ؗZ�y���%)�ּ����]%��H�]Z�C�]��c]�sL��oQ-t2�AŔ�u��&\�N\�e�+yt8M�?�����T��[�t�}�Fl����5���QF�oq[�Y��5�I*�_Yc�l����Y��R�č��!�V]&��gU����P�t��]
�Ƣ�;H��D���ͷC�ue\=ñ7DgH��Fo]���p7v�#��M���j���;(�&h�bC�&�5s8O����U�Ȟ6�ܺ`%i	ULA���2�òw;l�j9	^E���%Ҋ��kdA��A%�s��#�f�U:��;V���3����d��+�HļZ;z^_#W��uPt�B��A^��u��`���`y$��,���FM�E(�]��%�`���._n֎w7샬���"��\.�\ͬ�ds6Y�8Y�U�f.)��v���w����'�l na��:�W3�P��"ܳ�2����3u"p[_*u�P�Y��ǔ8��/�Vf�,��>�;��Wnü�1�]p3���V�3�X�#�r�p�/�t��f0����k���d�g*��Pmr3���#GF`�5�e����7v�U��`�AY-���DN�«6����4N>���l���aVU[ćc|$ һ��(�����U{��n�\ޤ�_+��Z�G��9P��vC]�����Y��M,"��G.�]��W�y.j+8$,M��n;�J\��v(uL�¦�[N�c��}�+邐AoOH���*)���7/-yl��W[��+���pb��*K����ʱ�R��n�X9�-ҍ�@L��bgl��u]r�Qd{`�����Wۦ��J��5�f�c8�\S�:χ���~� ̤���bk4m��:���r���^����sT%swUn>����~}��J�O���"�"].�׳&�%Vb!A:�X��Zmڅ�RS��Vj���PJ�]ńo�Z���m����y%*�[E�U��fw'H����9nƬ�=�� '���-�v��A�AS��fp�+9㩏��	_h���9rٍ��^���e�Ɉl�ܚu�!+0�����ܗ[��cX�yԩ�+����%|�:��=����<L�sF&+BH��^i�y"�%wh�NY������U5f���̇�r3b�f<��1�/�s��w�u�"Y�-��C�8�s��rz��$�9o@�uj����zf0������P�:��2��S3�AP}F����Ia�{�ps�n)	w�n�ic3U�/�ݠ�۱o�G�\�u[���V;%�T{��ūl�L
�������S#4Vu����� ��]<�sN�*�0\Mk�2K`l��{}�9㵿Y�na!��b�V"/_+5F�uy�ב&��*if1�['!z�n����G���L�"���Z��P�y�`��Z#���[l��1=�f%�Y/�4g�x��-����#[���u�@o��rfY���#LjF������ࡨ��ӶF��Q�zx�$�V� �e�5U���u��t�u3�@B�����P)J�;�W��lt.jS��s�F�i���W�6��1 �\%���ǣ�m�p��Wl:坼����XbxqP��(�WX9o.��}uN۹��A�H�Pd���=L�5�����]kd!Ǚ��t��2!bó���C7��V��&��,�c�úU�o�2dg.�m-e��7_.��Z� ڛE�f�R}�{N΁Akn:yʝK��}S�_\ �=+u�^ؐ���`��E��ԭǝ���v�t��3/I#�rM��I��N�ͫ��UgD�%'T���f3��x���K��w\kq�M����[�T�;7(N��ÖI��ۦ�9*���LY�n�C��ڦ&��[hv�G
�-��8�5,]%fK�n���X�9�l�0�r�	��e��%���4���9�w�t���>�����\V���}��ԅ��<YI��P]�޾p����e(�ɛ]O`�6tT����3�#�V-���Z]7�h���0�MޭF:����A���;�|Szy��3s��t��n\ ���f��n�Ǳ�Tnd�N2��� �J�M.�a��rP�i���5�'�&��sb�Y��{2��]�f����'�X@�U
�D�9)&�l�Ϧ�8���R�^�v�[�Ǥ��ͣ�&^$ɩ�����c��v��ن-�Đ�4�l�8�o�-2؇�w,�����lbέ�YO(N��l��x��*A��FY�b���ok�Sx`��,�>�~�oFs��c:ci�;��lC�����Su�X���MD)���CV1���Ee�3�fGi�{�^�%J��c�O%!��jR���L�n��wX�#��I�F]��;�j���\��21]W�oߐ��U� ;1�H��&��2�u虲��i!K{eL�����P��U��[�&���.�k�E(Y$wuv�3j)�����ho(,nF�⭫�n�t����þ��$偔�^��[Sfp��%���S'$H��J*�$E6X����ʝi�*nd��ǖ�q�v4z�m���i��t�e�Ի�+�r�Y;i�����WE��}��V�V~a:����JT��;�z\{�%@���5Zwe7��s�FnBK.a��+~L�I��A�b,���5�4Q[�tR�X�����թ����v$賻�V<I�ۼ�}����TZG��`��V�coxP���+�;m��ozC��W��eC"Q��M6�>�V�op8�Z�Û[c�m�߉���b�V��[rh&(��s��
[&���]y���Wn��+(Bٿ�p��.d5|O���l=��Y������ƇX��2u�)	d�i����9Jl9w���c�{ H���.�V��n��zh������^�'����%s|���4�yx�֙�C�VN.1^\U�vfQR�M�n�+��!�m�q1�g��nO��iu����r�j�C��yO&��u��i���$V�;�(����.-��n's6�B�����KP�7�f�Y��5>Bj�֮G���P�l�Z���짺�/u@���Z�֘�u���l��77LQ�k��ȫ�w^���W�2jr�mK�b��p��r�B6!i��YK	n�ڝ6]g)�f��,Ώ� �g�{e:9�YW�-Pb�Y��H�D
"p8;vh�iR�%���1C�rLw�N*�vk�Nc�V�)ܬ4��f�7t��;�KaP��F�v%jy�UtTwΡ�Yn��<
�*CXX7d��
�R��
��nn����i��+X�$�p����D&�=t4�]�δ�@�0�l��� kh�9�]F[�\��_�����C�X�I�x�g�ہ��e�ՋX���e��o�4�X^>!�<BU�%1��oV�5R�h�Ht�`K�Us����K�\��n3v�W��D+��lCw&�f�*5���x�f�pO�
7��<�=Z,J�i��u����q3���V�s:l�݊��v���f���h�U��Ĳ�ǋ(�s*\|-����L���b�;I��a7�CY�1>Hua�Y�²�ۢNsI������3�� ���h&�p��)ؕ�jV��\��$S
lb�
O4R�0d��T�]������u�6PJhG��']����9�6��*�RQt�B��|v�H�B������:�&3h���p�E�c�d�o��
�!�}q������@�'*�ᬕ�DʼQ��|�t�	Ԭɖ�oLK;��98��G1ow1|��F���X8:��Kl��1��J��sa*B^�9�ٴ;��'6�&�a)���B�%C�ou��n`�����{S0
g\�N��P�͹�Mء����H
�/WU�ΡIU�=ݯd��ñ��8�|Y
M�QTW������_[��l2|/�ol�
�HrY�M���_��dR��Y���V��U٧�õd�3�68��':��%�:7���͈l=��	(T���^i�:eXrn���na5�[	6�է��	���xU,$rm��!U�fAA�(�g�;p���Ш����[(�.1��)(ms�HQ���p��o(}�fE4ٓ�U����ps���D�R�|賲��Y�v�
��S�� ]:��~M�¹�m�|�.�Z�R�a�7�W��OV�t�Q��Iu7����Z1n��U��U��{��t�^B��s3��]g[s����Yv��R7�9��:	�m��ڦ���b.�9���P�'ʻ�0頟nη�4�k9���i��]y��we�bזAYB�n2F�X��=��GwN	�����Y���Lw�VM�+6
��6;ϳ��Uݗ S6�5�bx�z����'[BQM<0]���"��>ꃾi0\�7��2ҍ䜲�m���9�8-�O,�Z�wn�̋����6��g�[���m��XΰRj����Ws#:J����M�7qS��QV�MV��5B��
�ִr�d�T�Jnib>G��:��6���ߓg3��,�\y��cd��0�vK{o ��gdͼ�&��V`�h�0���,|����D��FX�[A�o_J��kkQ0����]R֡���1��Nw:�CB��{+F�P����B(�$��k�*'&����3V!��\&����)M�̥�([O{���4w�"�Y�{'�k�%N��OmaƑK����31���@�zr�+4�^=�xtz��-�:�U�2��`�)�i4jҁ�[���1S���.�j���]�9O�x�Ә��A�V�B�.��b0�8�睒j���\(��#�\���ݣ��/b �莃;T���A�B��p��ڛI�쮰�!7�[��<v����u��cu>j�v<�Ɇ�]�Xzao�݊�.pKcO�»2I<_>��PARVm�
�X]�5��L�'�n�LJs�U\ �Y]|�܏C�ڰ��j8��.��$�ɒ��lc�o����bWr�.�fM�־\�P$t� �ʺU��۪9�r�	�+PJaر�H2xż�i��֍��썼�n]�Y�g-e�kQ��@Nj�۸e�
Y�T�iv��	�LM㢸P-���6yi�t��˽��HM��u�%��Y���;[:�u��ݳ7\��9�T�+7�&K[����ǒ�Sz�9P�Tb���]��M�:��U��e��l�=y-ҭ�D���O�>�E�����!^��e����S��/�u����9BȸUt��:�G_p��/�6MZvv�];�,gq1��xn�tfW4����W��������Kd�<��A�-W-wwc�0��y1֕��{_Nw��B�sn�._C0*}:�Gu�Tʛ�O(�ӓͳVв�Kaa���R5ё�Q=�vJ�&�]���"�7MA���fJ�m����ŵձ+���r�`ɕVw����	�i���\�4TQ>N��e�t��ȠwP�"Nʎ��h�q)F)��Z  ���gqR!͵I෷ot�┻>��5Ӎ��E�+=/�'M*�a��;5+��V]���iv�]w�x���� dۭ�;���0%в��
����9��f_F�b���ݠ5����D����V�5Vp�3hpJ��Ȓ�
�ǹF���Ě��eU�KI�\��oK���1(ا�m�feH��>0d�L��q<��Z;׫��y^V1'�Zy�ǜz=�l�XcG���)@�y��Ӕ��T��g�� ��!7��nf���xV���7TF�c͙*���a���(X����`��PR��g]k�P��ԄF�<��^�V`G]?���$�x���n�s[wk���.f��ڲ�� ��rr��PU�a�:�z��ʝC.���*(x��׆���\�t�M�� њ��W�߆3�we0[�.9Ւ�����5.�����E3y,b����d�/zD�QKVK��*���v�*�GT��}x��6pΔI�R����`���V�朳Rv��yZ�KK+�%����8)'
�✒H��s�!(벶�,�o�56u��̾r��@35��Q���v�{�!lWRi����1G�Z�e#n�-�i�����l�	هsm���r+P��Y�L����s��YOE)x�vi S�Aئ
[ȃ�T�������G˸U�4�����O� U��??���_��_���Ч��������?{�?��>�o�����}>�Ϸ���w��|�w�<5S�Pl�N	q��)5��J�2ʤɡ.�G�N�HU$�|$�����"l���-�~.R��A�  �ˈ�M�1�B?�M�'D�O���V��������W�S����oR�z��jKkzQ�ƴ�ŇV$ЬWue�4��1�O���'�փ"݄�EvwYڂ�oV�I)Y}���G##{
�]��Uf�6���r�Ig#���f�i�*�5�/vˊ�!�{�vɸ7G�x�&^]�H�8r[�F� �w`�i�Q�*����vj7�ҕ�� ��펷�]�S��x6�,@Oյ���7�
����\`��MNᨠ�\�k���űVS�t�U��SH�G�h8Յ��w2����T�3g)+�Z�U�ԭ��Һ�Z�f�*Uvݢ��FjuJӎ�����Ry��bn�e�Z_:kV�,-I���s��n�!5�����KMٷ�ԫ��EX5er]��q�W��@:�S���<69�U�!}����[�t�M>#~�"�ֈ;���E;�Ӧu;���̏N����E���.��ӝ��"{�VՂ����KIۢ+��\uz:w��y�.�r׵m�:9���X����";��-Dh�*wW_a�x���l���T)�/`]+��fJ<V�".Sˤ������G!�gv���J�7�63SK��{&�sk
6��	{�w���x��3Fj����.���`��^B�q�����y|2�E�
}}];r/�ْt�Q�![�[�����ު���ρ��"��,�,��%"aA��&|�P��!��I��%�Q#NH&�����
v]�5Fˊ\�)Ɯ���l�U*l� f�A��!:R$LU��L�,�R�*Fl� ���Wl�YA��P�����$�޸]0�$�H�`�X"�5M�	E���~�9Q!���?	j�b+�ꈊ4;gl��B**������$� ��j����AIMlV�*�� �X�*&��V�
B�tQ��m1TP�R�ئ"*b5��E.��l�3DS�h(&��b#b�	5EQZ4�A0��1TN��ĕ���U�E[fi�������(��F� ��(����"�����f�QARPTTEF�Rd�b�Ռ��ITUV�3PA3˦����U1u�Q4F؆��DM@T�)�(��b ��%�"��Jfi�J�(������*B&������
������JB�i5��i((��+cMCIJU#E	QP4�F�4S�5A�ĄUT4D��xS����ɋ�uwc���b�*���A��t��<1�4�9;�-��w��p�J������.u��v&�+VEmoE��5��	8�>�w)�d�)"Q�/�rB��|������L�H����u��cy�%|stԘ(�	.�l��2����:�
ިgi��v~Osp�~F�ǻޢo�d�fw���$��s�+���,f���mW��Ut���K��̹l��(/{����0�,Aq�>k�I�|"�Cgѯ�I�\�&4CLŽ���\]q5u����}�b S�EȎ�p��ѻ����d�m�����>�}Α^���%�gƥ`�{�J}�=@����'^�o�"يvry���L3!��1"��<0��c>Q���g*}�p������>�;d����;ϥ�V�f}t�]yP�&�����ħ�On���=����'�;����l׹�Ct)A�����&�����[���
�+�묹ͯl�N���Ǻ��lx�/�dnZ"�Jh�7u��ҏ���"Ǌ�0��s��ht���9^ތ�?�˷`�{M<+�tA�;��y��H�}��ܫ۔��<p�<����Xx�{���a{1/Ŭ�^���ou���܇E;�K;���x5^��Q��_w���ܣ��/4Z�3�1S� �ˋpM��z
R����'8�^��	*��E��|���C6��*��R�zh��ey������zѴ�j��ۈ,�oN�]�7�p��_`�����sྀ�k�+	� �􉷪�v=���J_����9r���"��g�����k�f�]���ɈE�䢍<����S;��ĺP�'�ez� ����1e�g*#�ﭞ��l�SÅ�����|���\\�$e���#�c^I��Cotؘi���z��k<=
��i��u{��y�ܧ��}���=�}n���Yb��J��.�o�V��N�ko������	7�+�U�����w\\�����s�1���ᛒG}T���v�VT�	\=�O�
��%�s�u��k��S��$�x$��<j��{-t�F���� �g�d$,��i���f��_�w�xI��<m�z@9�#��C[g�=�9Ux�^8��� ��V��[[OBY�փueuh��.kL�˘0�&�O��+��qɪfB�����-}o'ܲ�U���X�]��`c��~��.�G�kOI�M2��ڼQ�*����� �.lܚa�D���>�#���p�ƱK�j{t�2r�7��_��g%{+T2/��z?K���Ы��X�K�J{v��G�E��{�)�7ۼx����zz��x��[F$߱3W�c�~/*�Y���{�dg�H݁p����D�����w�;k����Lox�u���\"�������o5>9S/s������Y��<�Oh�p��#<��'�8�T?>����}t�ة^�Cȷ'/x>�-嘥��/�z�W��<!r�)1���Rm[��T�ڹ��L�3�ҟ����K�;�W�t�kN�ek���ITU���Q�t�b�&��"Y�؂����d�eT�~w�O�	�'O1�ȉ��û�p�q.8�b�g�Bƶ���u�Ss`�{�Wxzڴ�d�٫�s�~^Ѿ�ey�������:WX=(E��xH�����?��q��v0na����.��j�n]�܋{�v� �Awj���Y��A2�7���.����N�.�}'�v��*R=�rX+W{��F��TB�c�����&��VU̅e�I==�[]P��G���:#�|=�3W�
por4�@	�6�8fn�����z_*\�<�����R�#��wG?���ͿP�j�w�&u���z�k����/�Gkt�^��hA3 ��s�Nf��t�v��yܻ�8n*����[���Ms�4OE�ǽo^��#CLIEܜs������ 9"܎�j2��7h���m�>'����Y�>�g�j�/��z�l��n_2���6�l|���3Ǩ�r&Y�&>y���⃝��NC�2�N�)x{��u��?{������{�g��l�eY��<ߧ�?z!�*�	�ʧB��ھ����5�K��M�L�e�R.?V��n�}'��|߳~�����������Y��:_�K���������������̸�.{V��h���o'$ۻ��#e���tTÂrrDF���t�zmW�+\�R��?��������G7��Nfsڞ�p��*��L�ƚt\Ͳ��^V�VMTI�Vv��Y��]��6�Ļwd����pǮ�?�6{���Y�*ʾmk��`Z�2��Ӿ2���]r��\e9C�P/"̭,݅bp̲�A���[1h7ξ,�m�_wp�QQ[[�i#�U��P}�u�����S�����Uɟd���if����W��ב���z�V���eLϕt���z6�}]�핂����$Ω�2E��^�u�Aݔ�z����K��@�����b5�H��e�����C�$�xe]z�S3�m��Ɲ{��ei�����6�>������E�H�r�����w������n
7Z����c��]�1�_�C��nu�c#e������������#q���-�o���]���z�*�砋�A�{�g��:|��'�	���X)'�nC3��9����8��C��N	"�8m�o�۰I�q!�p��7�C�{���8�3p���%�}@?OKv�K���]��bS�מ�u�#�+��k^��>��-�p�4	���@�>9��;�}����Z���}�<�ni>�%;�]
ɚ�:,0ݹ�]>�@h����|�F��q�<nY�V�vde�s��3kA�w!I���&���+\̝�]8��zV��I�洞��w��l��8�F���[	�'-�0>�-x�ni�*J��w�S�{6GnI�n�����]gk��P<_� ���F��Tq��z��㾔�%xh�g���j������z����<���	M޲3���]�#�$1�����&�D������S��zC��k����+q�;�{mǣ�؞������J7����˜���Op�pm���p�[j� �OX.A1i�5���!��[.��U���ثۿfV8��hq
�&�5�O<�5�1T�99��\�ycß�/��u�mu�V�Uܖ�XdXܿ�=.��9�H��e��$o3{�ws�X�Ǘ|/~�L��oi<k�C�7�o���*?��M]v��,��Z|M4D��j�7��o|Y�&9/��\;ݞG�����a���Ll���/��&������ �sz\\��v[����B�*��h�e������n�q�}N���LcQz2&G��XMrP����_���3��K��N��-P֝��pH��sD%�5�U���dLocY1h靌}.o�f��lS �Q�t=��������x�:�D&��]b�3Y�����2-�DV�Gu�Vn�ޕ�&�{��	�7P&�8*=�V�z�p�zJ-�G��{:����9��o_}��nFǡ"z��O��^ݪ��VU�חT���Pxe�q�͋�tv�T�w8;M�M߹���w���
[z./X~C�WG#�0�_K�vl��G�A���o��g���'����9����}k����׌ע�(ҍ-�+�G$H7��p��f慨�\u��?w����Ƽ����Ns�繛S����"����߶��shn{j���W�����ϩrԔ��xr�}�1W!Yfp�5�F�ok{�'@u������1����ݧ/�7����k֪^1X���P���g��q�{|�6k�K]{�_+}��Ws��L��W���{�8���f����bW���j5J��y�=g�N��jx��f���ׄ&�����T��Z���^\�~��1d��% CЫo�%jw��bj�Vs�U'�L�g���R�Si3�is�����9a4�':�� ��������l��ߺ�@�I�����AV�C���Ia��U�0���o1���p�&n���=µ=ͳ����2���Q���d��R�^�y��t�F�O��8��!���$l��՜��#[=�r� ��w��P���¼�����vf�����}�o�*�� ����4��lw��V������CX/�"ݪ�DLm�@>Iݳ���G���v��r�n�����z+5��q�j��W���K�}���C{Gw��*����{H9G2����W74�n���S���l~���,W�����6��-gq��}�O=&�̝��6i��{v�_/5�E��7��	C�\~�ꌶ�ggͤ��~&�5t �}����E��9��ȸ��ngy �EӒ ?��,e���m������S����-w�D��H|}��խ��U*Wg�W��%5�<gA�k3�@U����Lu�����߮O(���V����+���3��0�G�����*���3�ܕ�{�_p�ʗOt�w�o=٘}�K��VuX"�#�,qk|'�~�[9�wh�6�[���Ȥ�Гi�`�j���f{'+85b�dȻV��}��W���E�m�qϤ\p��yۓ��nC�a��Y6�_$��'q��ݾ�]Jj�uY�n��ϙA�o����!�C<E�/�LB�������Ǭ���Nf�G�۫ة�r��Ǩ��k ����O��ғ������mp�8��v:q}��d��}�h7��sx�U; vP�T���1�Q�y�y�5o��n�As�W���k>�x�Q���^������2cJu�[����=���6�mm�q^}V��}��y VVи=�V���};�w��P�a��e��+y`o�5�OoX�gÔ��}��/ݻ�������R��e�E'�T�tj{Օ�}o��c��~�2���&���{��\�;�lU�ۋ���[÷�Mȝ< U�ח=L���@<	��{��k�}R^n?zf�(E�H��/�<Ԟ=����\S��X��r�mK�=��y�^�����tFF�m�n�,��{)���5���|�W){֤/����;���ޘ�[�v��PM[�.�4����Y�0e���M��`��>�U�8X��_�i�6�i�ΙzX,Y\�����R;e�5�r�pͮ��逼���q,h���8h�ث�fM��6�o+"�h́�Vs�ȶx�
�!)1�
���vi�i�uQ�0H�6�F��m �7g��33��^Ǉ�F-7��U,O��#�|���eh��q����)�^ɝ�������:�Kn8�f�~-�xߛdω&Cw������_���q{�3���[��5�[��m��=��u�'��s�j����W���l��Vk��o�p���ެ��t>��l�f�y�{�8��t�Ū͕���ו�U�S�WJg���==E�9���g�oݽ�sm{�?w������B�k�D������<�8���zM��E"�6�w��=��ǳ��[�>���t�%9�C>���e$��:����{L�ʥ=n��>��)��Nc1uHj��Z�Kb�R��v[XEEd��b���"b��yN[����>{W1��S��J����}����>�>�o�����|�_/�Ǐ������U�/pw��.��E�����ݚ�w�fGS� ���.�N*� ��yg�p��`�������I��FT��:�Ҥ8��.�]�jҠ[SY�R%��sD��������v:�ț�D��m�H!ن�&P�=�)�w~͊.����uC�k��;�Rn����DU����y�L�*X�S��.MoqX4�cP������J�ȧ=oJb���E_}o���uq�\������/��uӆg/׼��W�򠽔qVTE�hq�[)��+�ϟY� �WL��)�Ce�ef�s8�{j�8yl�P5�L�c]>����p3,��KvMgc.���KU�Eqb�<oFV%#/�O�[��yW/
DBYG�`���{+{%^a�u�B��K�8]�5ҵ�l��T.�b�s<�=�t��M٭&��8���5e�3��Z黹.)q��z�n����'HMF������r3�(,+�R�����Gd��sx>�Y��y�Χt��'t�H���v���a����L�q��0Ƅ�lZ��|��I`��)�I�L@���D�S�t6\$o�DCu�+��\�ea,�֌���v������G�v\�F�����}X�"�W+�H�j�y�ɚ�E]ø���v��@�U�O2��O9g��S@��ł�o�`�y����^��Ɇ�ET��p�Ԙ�ү�����h�B�@�GT&��iU�seU�S�bT���w���7m&����"[����<�Y;�su*
�Cȍ�fƙE�R��L �i2���.��ᄶp�W���xR����R>��U�.a�7Pm�����2�:_fe�*j꼆蚄�&Wd��޹0\E��|�6-K�Vcb�Js�y=[t6��Ɛ�X�5���w�c���5�Z����E���n(�:�$�y�^��tXΤ6Bsx^�i̷O5b/�	���YR���W��lY�wd}"|�V����NƜ�JQV�v�o-PZ��G"}XWT��El�Wڍn�x��	:�H9�m�T���+��tm�8���Q�;�:���N%�jLCihu2�u��uq+��3�i
�mg�@������)�FA���H�çjm�U����(�ά�EK�=Yd1r��ht\M"f��|�QS�P�|
'��<+V��U�.�=�D�]����J��;/LT�V���m��"j�W�6RP�58BD厷z���!ݾe�/�sAkk~s^�w�b���>YPC��� �͛gm�DP��AO3E6�L�])!|WS��f]c�s(BZu��V��3�Z����$C�O��$̨�]L���A�Z*F&Q*3%\4�bJP���vw�Ⱥ'��^c�c=��qU��Rk
>�U`�fN ��msK��U�S=M)6$��#(i~���ֹ�����'��1X��8lR�,N.ZYwu��ͼW��=����C+-]���|�f�w�(eFk:��F��1���~�A ��1M)�^�
hKmE�4QM�%�%,SPCD�B����	�*�h����
X�X�����jj�����R��������
J*�Ŷh
j )i&!��""i�E���!�"H��%�����RD6Ά�*��
(b):�كN'���h�Ә�N��64�6�����v6�j�b�Xֈ�h�-A�=a��"kF*qRb"bcZ���j�:",I����n��EE���E��Z�bb�bJ�64c%&�Κ����
5������Ul֩��C������`�E�:J+Z��b#f��I$��ͺ�����N�ˊ�8�ŰP3�i�VvF�ĽGU-u4h(*�6*6��OGK�$�Pb
�Qߣ����)1Z��MhӤ4Ř;u���:��ί��u�2��x�ާ�ƛ�u٣&pɡ�h�I�But���%)B�κQ^V�7��4�]%/�uL	�{������Q�y�vNN�{7��Q��&|�n�0v��%��C�@"I5>J8c��DT9�f�3����q�Qȉ�yY:��Ʀ^C ���.p+��ǵ�#w3E�-�cjn��dÇ�ɴ�5J�	qp�3����4���Zѹ�ڮ^�ν�5�����FPo�S��܈��jJ��� �\[y0L�M����͎� nmΌ|����;��y���4^�XE���ڡ�0��a�y�\zxP��%����M��ldG>r����,�ݚ�gP�q��^�g@`y�ޚi���/6���$Dx$}ݲoDF�՚mZ ��5\r#^� �A(�I���JT��&>�x�ϯ4�� ��Q%ٱ�����1�EV�@Ɗ"�M6�u{�a�y&q#��~���~��D�VH�T4���vO5>Eê�h�s�z��(U�[�S��0�Y�����dq��i'��)9X�QR�-��@���I��c*��Ֆ���}�>��E7�i�=���^���>��`+��a��&�t^��!��\P:�����D�U��pSnӡHnM0�>�>����遯Blp��}Y)��Us]�E�}�y�d���@�'LM�]�³�N�+��՝zgV�����"�u{�{[S0I8c�L�ְ��k���}��W�-�yw+��n��:���Nl������Y�~����yv�k&���S7X��q}Y�Ș��Y��ˀ�<`��Ά�L��kǾ�α�}�
�C:(���,a�>���:yċׅ��k>!w$O������_x ����W~e����n��2�X]O2c�b� z#��(pZC�D��#ߗ��~��6�Ȩ;�tp��&q�"%�!V�|7v��j'���/�^�=>��������ۯ��8���xo<j�&+lȼ�7�c��&�C�-zP|�]�P~���pS�8���+���-@��эn�lJWnɛ�f���gh��� D�� ߶�k%}��A�4"�2n0�[I���B���7��a�����m�L&~�� �.�{��+�w�a�j�G�Jݾ��<�]K=����
���`�)�[C/�v�o�e�s�z�{dS��|`��ȿ
��WX݊�͞ޖ�P�R�sͽ�zTpp�B�I\��QFu��f�qL���X02FI�1�:xm��t΂l���9x�m������d8�	�����z��ʊ��z:��ʋ�6��P-��e;���Wk�O��qq��]�l� �� ��� ��&):�F�+�0���-��ދ�S�)��5[O1��t�~ 3�I�j���P*$���e+}��޼��&?Q3
yoҁ�
%���_�:e�b�\|M���v()uMR�ym��u8�P�R�6tf��&ŕ�䷸;�ĩw=�=ۄ�y�W����|����9����jA�z���u�z^vL�8/�I|��Z��\͟��m6��+��~x�Bn��� ܗn���C�&I˯D��HеbU��˂X�"��1�F�kj�w��Y�iaӭ*oD�#ېqb�M�ۇn;�0���T�c	�[�+N=�1,��~ښ��PvP�~��A�3�v�xab�7$HA֘pNhL��|�`�5���1�*�&���c�k��5����8��|���J�Iq\�AY�~�r�%�?7����8��S��9�mл[ԘQ�\��,ܤ�iIc@#�?���X�8v�!~<~ܰz��~b�Z�rz�/�֪{��r����1'\]�TXZ��RUְMtl����0����qSIc-m������&U�#�k8е~
%c���+��PK�XU�N؝`,&��1������|^�`�3\�z�s[R̶�h��5�P6�����a�u�����{!�GJ|����C�p�B�~���_�ނ$�I���@ؙ�s�R2.lwK7�=��{E��:y`���xvZ���]�^��� ��g�9�+~����[|=�� C�|a]Օ����oT4�ik
buR˓�#2xoD��^g��(]G=��L�i*�&L�'��'�S��Qw0�B�n�����v�����Ux��̡�aՓ��v��.Pw��ɋ&��*v:���9�X�p��q�},
<����Ż])�s�\��[���h��+�W�L=�0�Ǜ�o�����pY�ǡ �IH$=%�L�H9f�T:&.%��g�`L�!_����h�1�iW��5���"NmZ��
���۹���h��C�W���J�!^�k�o���ּ���viz���V�6�#f���>'#2w��b�1��6�K[P�R��a�,���<����
�N��-v܁ܽ��ԥ����L���D.F���?�\ڍ�O�Jl�d&K�NI.\�
r��sk]om {c1���xeOl�{d�{�L��T0!�v)�nB��cU9�)��jP����j�s��9�R�T.�f�����;�amI��0O��o�wRzl�;Xβ�9��;��!�1�L�Y'C�YrJ�
�|ᮢ��։�DB`��b�o6�t��ԣGz�6 L��L��P�;"���E�y�)��0�_�����kÇ�#tB�1I=�1;�����b�E��`]�D�;JUeWC�zO��(-%��0�Ʉ8ps �;)|�F�t!Ҽ��=�:b�F�ى.��`Z�Ӵ.��Q��j;�M����޸�5˲�}gm�<sO�d��[�w1���\��ʫ\�
�k�#�%� y���l���Cr��k	y0�Iт�����\�!C����
��y�[�:�J�\�i���̴���w"�,��s)e*�km�/�M
̨������x���´�\ �Q�{����Nǃ�B9�͔ã�9�ڛ�������Uk
�XG��8Vv�)ک{�l�L��s���Ѹ�~���*!v|:
��'���4u~1�hUm5_��k���p�ۃ���ٚuͨ�*}���u����y��rY����}�����Lh���q2W-�շ�ۤ>lF-b06��/GMOy��9(�A�Z���I�h���j��Ǟ?�=uU�5����c
C�o�\$cr]2<�z'es�Tg:�M;����	C�@"I5%�[�v"���ݘ���B���e��ܡ�t���s�;S����g;�y��wj�h�	�*�z:;x�!��J���#��{/����?Yf}�
b�֖�&���sbj}<��3�Z��m;tޝ�­�9�T'#0J����8�X����~T1U���)g� ��,/�Q���*��W;<��~��h�շqO�k�K�Z��-K�{�daG�1��[� �d��%�.b!��Եm(-�1����5�X}3���	��=�(�je~T�5�����=����{�`cy�n_�=��G��8��I;�h���.C��&֠��Թ��m����t�+ޜ܉�'W�pN��{����7��Q�d7��л�{�5�ޗ']�;s��)x��Hr%]�q���Z�_˥��A�_M&vZ<��V�9�1�����^�0�x{��k.�����;6|&���vI�?D�'�)��˼������j�p�X��*C����[-�ܼ���!f���gݒ�]�a�oQ��<�)9X�"��,9�����l��>�K����j����C��@�t!)��n��-I�S6a7C�F-?'��v�����l��8��rn���]琫��a'���XE�2(֘r9���.~��n��\���xɸ�a|`v��n�'��7d�~/��c8� ĺ �xQ��X�]�|���� ���7��cw�FI�C-k@F�ƻ�2��^#&�lR��
�Y��Ż�l�0g!���\S��`]��%���1uo�LU�lz�^چ.�v���a������=]f����`O��;w;�.�>�L5�UV!'M�\����ٯr�C��Ƽ�m$�ߓ��Š���[E9`.r�9��Wu���;�ggV"��H��9���_u��L�v�-�f,Q΀��0*��X�1t8^8"��E<vl�wq�ߚ�	:��8�npwO�ٖi����{\p����l��m��ǳq��m��N%{O�p_�����C��/��,�Z�1���m��b3�_-���2a�b�6G�5+�P�_nL��)�����X	_�w/�8gt���9ʺg�I�T��qP�$��j,E_�����+�ᶳ1�^k;�<�>o{���!F'k���h`�;�˷�zm�j(ː,��)i�X�X��'ఃJ��-W>�D��6�<^d�x����< 1��H8��2n\����>lS-�Ξy�� �c�0:N�!&�l�E���m�sW�4��"�S�VժO�ga��/���������u�D|�*���d��\=������t-!\l<&����ܯ�6G@^����yN���U&���8�h}1�u�J�5;i��n0�n��P�������K5��N�7%ۄ��SsP~��9v��p�O�wz>.�CVgf̾h]�5�|�`����Uэ�L	֯C�3b^ܻpmΈn�R��3=W̎�f��j��g�t�yn��"��$Mxgם��n8�����r���A��Y7����tv�>�M�
 `ꔞl��E�.9�iy^=5������m  �^}Cw8z���\�a�[��Ç\kn����J�m&�e���E���������Cr;ѱA��s{a0��,fق��ճ��\p\��%��������f�I��U-t�)�u�Ң�>�sۇ|�˔9�a�r�]�t�V�<[��1.���W+ŭI�Wƶ����\X�`�ki�@�ޛ�Y�=s<�mzQX�����z�^+Y(S�Xŀek}�5Z�t=�'��Nu�\���}�J���2�{�gW"(ХW9�;Z��]l��;�ˮ����|?�t�" �Iۈ`�x���[X	��1��ۜdRO
�o6����=2
�����£6o�Y�Y=��GU�@[!�a�$l�g���9�mK2��Ú�v<��i�k\
��:�uj��Y��1;] ;j[��=�/a�ɑ.�8!7�;�^T�$�/���ګ)3��gj%�����G�t��.L�S���� �@�r���H��C�|oxo�5��7�Z2����?�N�*CT��C�A!���B&a��Y�}Y�^�π���as��Q9�vnWc�y�̄�JOb�/^���cNd)��/A+��{���q��t�æ�n6^2�[�R�d0��lnwfT�!������O�Q�]0��g��_���eХ`�<����uƍ��ӑϠ�r���y�<����Bli���U�.'���gY+�-�A��M���ɽV�8�|+^MVB�O���B{��߂��p+�ᦞ�� @Ųa>C�����#�O03���«�L���v;����x/��I`���B�b��_q�W���;�amA:A����!8���S4�B������K�~�.9HiAqR���$�i����T�Q{�w�m��`�S�B��z��M`f��ծR�h�U�v���ٵ6�!�����9�h6�L�ML#�p��u��o/�ڀ��i�h�3����+Vm��V�|۾���1s���=�����{�pd�sU1;L���e'XĲN���L�%޴���0�����'�}h3cyk!�m�J��>9�G��r�n��e��!`�;"���J.���L�i�n.eλ;���)�6ڌ8�r��<��'e�6�L!	��<t��hQ����YS��Qo='�IO���ҡ�ջ֝��<	��B:5���A���Z}#[��SIј��=0:f�qRaͨ�u/�-9�K�uL�6Ҏ��C9�:�`��PH���` �j�SM���E���J�`�j;���-[,�=У6�뭧Y�Sܺ��UP͝�l��+��~��3���������Y7Ц')�y�r�%����w�Us+	���3�עf�\�l�0�v��	C��Lh���a^�f
���6��lZB`�'ǽ}�ns���_���zHz���&+���w�X�c=�v�F��r4�tN���`ȰA��}�O~ڌ�'	��wk;w9!��@"A&����[��ȥ�����۽���?e��(\K<�->C!4��'���{9���֝�4���,������9����d�����!��Z���,���EO?H8k;ʣ��?C��G�ǅ@���z�C\�0�:f���Ws���A��K*��ܹ��e�^��z'	��j������2cv�X���9�d����x�1E·7��w�| ������F-k+����ܛ/��>W��(� �0~��x�>[u�m�jJ���H���/n�)����[�W��0�(�ћ6����{�S�`qmâ�L\zxT��	?��E�pt��ܽa�5s�G</-�$�ZR�&XbS�ҏy��-hp�V�8J�_�e�+�RK�������Z4��=��p|ۀCٝ`\��bY'H�S�JSS�S�h�Ξ}�v"�δ�k\��y�9�N�6Ö;A�'���Jt�������U�&���`5�ݒq��kYX��ۘ�=�����6��ϻ%�)�L8��4��yNRn�E�y5�d��)���U/:[Ѻ�<���P�?��0�a �#���Bm��ۗ��E�S�M��teֹ-�˗>��)�8���Ɍ�/K���21,3Ǡ?y��}m�s���,��ud�s{�hp{FP�l��0��s-x�^��61��c��3�/	ׄC��������w����&���7=#V�C]�౵�Θ�G*ƽ�I���d���*�s,�@l[�6��`��ħ�<=�O�����~�?/<x�����������P��[[����<%���}B+1
�Y]VPR69Ny	�f%�I"�]K�޿�Fq
X6g�ɦS����;��e��f�9z��:���4��x�aS���2��k�;�3�J����"��t��֩T{O�*�T��
9-�7�aN䮳]#�M��Շ~Z�=2n;n̈́��b�I��-L
���ޢ-�L9�+�N\��F�7�f�Ί�'krӱ�zB#��1H�:w"/3�j������o�������X�2ĭ0К���4�Aܨ���7������Zʖ�U��%�|�U� ��c̥��v����-�̬ͮ	���R�BR�ݐt�]n����#Kp>˩�����)�;:�n�[���	����b���{Llͩ��d;ft�A6��J��n��XRFk��<b��yk�eS�u�w.����!�S
��1�l�:�a�mN�Ă�n�L�ni�"��	_N�x�,��V�:��w���LTc������ܽZ�.ww��!-P�]�	Aѡ��ѭ3F�&�jA���;�kB˒����]�u�;һ���t*\\�nZ/S����y�:�tzq߬*���h�c��(*@�ݳ����M��5A��%�������p�1�Js�Y�����W��>�(|f�,w�L�[�2ʝ�Ԡ{�6�<�;iH3���cR�U�i*��0g_#�	K"�72��\�f���]'�NkX'S�yC�' +���H�Un��N���2������� ��X��B����ڱ[�:1,��:����WEk�7&B9��
�e�̙&�k#�5�v���w}�i�u�8��S�-J�z�� ���x��)c=��)�d5$�r������їn�[d,Q#z(����%Z(&f��e5������QݳC�U��ªG|�Z��W.:��]�ň�
�0Cl�̅��ӆY2�Wt�[F��z���
Q:}5X�z)|�A�T�J���Ȟ1�u�\�,7l��3NS�0����սUO#�؟K�4b(���j���4�l�;��F��(`:_pC1��11SOL3�7a�0J��P�@�[��0�]�2�XN�9���[�H��<��֭�თl.@�8�ۜ5��o�7�3Y�$��}՝�����=��C��a&PS��^i9	V臠Q��m\krb"Z���ˍC.�ng%��ֲ!�����2��/��q��1�T{�
���s�w\@r��3��5ّN��Rv&���455��vb��U�X��5N8���z	�qõ����D�K�j%���~xXyP��ut�2���T:�#��șu�ìk{vݭ�+���Vܬ��/l�"H��P��GV�G9M2��1��NȒ��4NB��7\eA�WO�J�V]�8�nF�d��Q8�5:oY.���u5�1pӭC�R�TG��Y�����v;��'V�U-:a(6�&�C��N�4�E8ڊ&��j�;Ɛ��V�L��سh�hf'mI�Z�=n�Zl4�MV#Cl���X�hM�h��TP�qD[!Q��ZMLLU�SHh�AM1#;h
)��z�GD5Hu�=IMUh�D�Ruh
u[��Xt�4�	Q%'SZ
^�H��QZCF�i�4)�:�M:]A��D�CCT��H�)))����i)щt#ԝ�f��-i(]�/P�Z�MS�1�Sud���R�l;�D�m��F�
�n���Z��(i)(i��!)B����%h���������qST���(�"ZB
����)�"�M!HQ���뢼z�21A1�dKiU��ʐ��w8Me�D�v�驦��VM�Ѣe�C��xeJ�/��Rºo,�ϣ%=��pl
\ѩ�nP WU����I�I�،�I$�iH2Da�1&��� ���hC���N�H�k��(��p�"#O�?��;����
%7�$��8��zt���_�?�uv���X��Uʖ�U-�nLy�xD�t؟e�b��d>����i�ũ�qhk�W0�\,��
��n:2[�Q�/̶��s�<!0��
LL,s{R5����w�	�.����r�v)���n������/��=�W..�vȗx�!�E�4zD�$�-�����z(ӵ��D��Y1Y=͝e�������	\s�zҋd��-�?4S�͑N�=�����!�-�E��]bw1V(ac��l/Q�y�C$PaM^*��
3��3f�Y����xo2�HQ�/��)��m�b�=�$e�Ct�br*ڴ&Cy6��A9��Ɗ��z1���2���{�d[D�퓨E�-�3/!�/�0�%�fzbu�F��MQ��۝Y�&->X�
P�0���6b�r����7��P�T�dTd:��| ���f�t��nK�	��sW��2Of"S��J���I0�+�z[{]lj�ӵ�ſE��zh<:q��A�" �a��:��v!���5y����Y�{Ȗqo�3�˾��v`[�p��q<p����68v����.�r��O#��� ��5_��B��Y���j���y-Wb�����ǈq��GB]�F�[���q�g-.��5�����>�4rW	S۝Y�[y�����3�x�R�a��B��_ ��P*�=|s�����^�=z�@��:���	�S�D�6 �^���N�!�!�!?C�9��\���K>���ez7��v!���ijRyoX&-�u�k�9�-/#�4^���: m]�l$7Fb1K��z�󎆬t*�E'W�hSyX��U��-f�'����d���̷!��I�3�r'wFj8�&�J��z�TW9��lu�߸�,*�O2�S�5=�}i�y�)sʮ������P��V1��4�
�T�m�2)pQ+u��+��T�[<��N�A�}���f�mЋe�a�H�p�3?���p؜�ږe��E�0R�k�(��o��&�ݜ;J��S���k�KsQ�^�/a��>i��*ǴBa�6߯*Y�uRv��݋;n˹�.S4��Z��\e���zF@�{C��B���Q&��$y_aP]��7w���=�^ޘ-�����a��C�t��Pi0�L��m�ll����ly�4빮�Q��Ĉ̕�b�/�u������^��W>W��O�2�6��<���tzoɠ	���	A#<����+^WlXy9Fw 6�B�����~V��W��A��h�p1���v�r&tQV�W嵜�3�;�}$�Ө[�v��>��IZ9���Rgo��ԋڝ��n��Q �����}�5+�\�㾽���UA�TZUP#㝻���]w��'s��E?�󢞆�/�B;W+ʢ�;�K[V�!7���aK*D��hx���P�Y�[7��<��=8P��e]v�s�)�?3���#@~ه��P����Scn�DsăP�'B�C��F�{������Eh��p���c��6���|et�n��fU9H][��^���1�.l)�j�]���׵�վ;����Θ�c�Y��h�_&�3���f
薀�qW�wL��ĲN����$��?E�w0����\��W�Q�P��r�ቚЈ��R�2�hpvQ��Ȣ酣R���E2������NX-A��iG;��ؾ��|7�����@�h*�:��� �H��z���ڇ@aU���1i��r��|��t􉢕YqųU��/k�p��>ߘG��Y�>�f��zLN6y�Y��.���cr)PP����3�i
��2�~�로�~�8ϼ���0?������8u��6��U�d�2o�=�N��#5�7{[��K7�{x��I�z�*�@7pv�����~��GW��S�N�_r���4�&��62^�DV�T�N��Y5�N�Nh
ê��i�����.Fm"{��"�U#C[��4A�*���EIab���^��E��4K��T�k������v�����7U�8rZ�׳���r�����{���^}�Ȃ�̂��� ���լ���Zڀf�|݊c�I�����ϧ^�L�5�f%�3�����z��3;5���B�En���t!弘��چO�7d3od���zHz��u���|�Ҕ�"=c;C���Ȫ������א|a���&%M�����2�N��i�C��D�jJ��H˃�**r!�GÂ_�b*(t,�.~k�i����������u����0_H��k����|n���bmQX��vy ����_r����2,wА!���d�����[�8պ�WQXs"���c�_S5��PcK' ���@͛OX�o
��)�08��^t_dzxgwJb��9FF���Nm��
�ǀɘaSQ^�8�)�����ɨ,3I�J3�+ǣ1�[ռ�|w����gH�Ϭ;��L�nt,��๏�T��svB1��k~�����$j�b�\�b#��s�:~��Gy�2��V'1��a�S������S	�����X@�+~sΓ�q,�.�,��\<����$��+�rx����w����kz��z<�[T%,�^���}�.�H�a��Q�����_�z�Z�\˾���/'��ʷ~���%̣䓅��f�"-�����҄TX�ʙY�a�� -���gy�"`M��R!68*LXI}X1J�v��a�]����\�J�Q�y��^@��I�b](Ȭ��EB�y�ā�w�Q7��W�Q=;{�w�Ͽ;ǿ���i
 �@�R�F��B� )���|\�4S�*?�?t��о�M"E�����~�#O�{�<�,-��G�Ȅ�Sd^�5:����ģm�����=�����p2�K�\�G"��at��d{���mxrS?�uK��pc`���+iE������k��R5�=���2�q���ѱ�� $�:A���~r�,�8��3e�UD^�תC*�V:�S'&m�7�'汈ɷ��>�S7i��W��y��e�q~��=ٌk!��a�:O]P��ڤR�S�^5�������5�^�v�}�x��hJ�[v�������'l�`��9X��C�azP����4��$���s4�t�3E��5V&U�-��Ռ�}���V�)��/����Q���ʃY.�����a�'�73S���"��;��j˲�.���ÉDY~h���`�1���:-q��?~U}S����?8Ug2ÑV[o[�� ��%L�A)��@%6�7#�o�i�sͼ��	��c�r��UR]F�vfl,l/3���r�Z�(D8�0�&��Pb�c>��g�cW�*K�����xw�P���T��Et�0Ǳe\*���f��,���b <���n�>�Ўwv���rv�d�x��x�v�{M����u3����������/���;๜x����<��<�TfO������~zn֞����������{��xx�R�B�
EZiB�C0f���7��bW�����~F'���½3r4ߧ'�VתO�}��zYYӌ��o�;d>b�!�+ݹ��Ԧ~��(h�,9�e�g���X�r��A�=�b��FD�B"3��p[W<Ҷ�9��.`X�Ŷ��9��u�[Р�5��Nӹ.�$�M�A�$맃i@1� C��>r%F9@�f��GN0�zh]��FG�e��e��ece�#�J��V��l7��i�%��o���dU�$MpgӾ[�	� .fN�p$'��VS�z:��:�
�ʆ�k鄞t��E�1�̴���\����f~vmW�uU[DXm�p�6��wU��A�ݤ6�y.�L�'%0��Z����O6�QgGfjxwf/	�dKbw��aF�m�:m�耛���oEs�5^��A�:���G2�ְ���ݥ�}u�ڢ�4W!閽�}`��mc�`�����R9�8Ȥ���_�s�b�}�F ;�<�ʍZ�-Q��4�G����a.�����ᯌ�����]��{o�}�_�Y��m�w�����ָ���6&1q����ٲ�s��� ���9b��Wu�f�3���A��f���h���d�P�8g޿�ye�T*�$%-����,�j��� t��ɛ
;j�;��k_ӵ<���N����	������#JR�"� ��@� �� �[BI&�SM�ߋ��{�P�;DԷ5�0��Ɂ���x��	��bgm�jpk�NNuZ�/A��ߗfS�(��bK�q�c��"�ƽ�-���;א0$l��L-��Ng\wk�yׄ<�2nq���f�����$:Ndz!�[.x��;w��[�-�݈�r��((Gc���)�����ƟfA!�_A�+��"k�m3q�f�c�8��l�lX��r˦.'�{��,:N&.��Q�]br���R����aWG�b���y�i��u���A$�e�yk���E����p���L���cH�0�^@nv�G��2X'*[�p�[&��R�&�)�7_�\ւ�	��"S���v@��z�=[�M=�ϞB%�'C�z`$^�+v��G��c^n��K��y�9BS^��RX&��B�6o���xOV��C�i}�9��9�͛Xs�,?;�]�؅HA<�ր��5���U$�'���y�)�y%I�s�9�o�2a9R+���z����Ls��vHl3d�����ݝ�"UvQ��Ȣ酄jQt9�-5���̃��o��eGϞ���æ9�u �(�1No�91��iT�����s�u�d����)�RD���"L��Q9�M���;L/��&f;�37F�+��5ْ���롁��>ǍS8�V$�*f�w����9𜫨����[�u�o=�����ȟ0(R�B%+�*�
4����ĂR< �.c����%����6<M(fƘBuL��dI9*IUt=1i��l9��̮&5���ޫ8ڎ�5��!������C������9��A�������˴&���WFJ��홐��)�삟�º�Adi/N��k�`�}!îsC�i���� �<�-l�/��366 eV�+�k�*��c��3�p��vB�:
��0��|]ej���c^�V�ɚ�M�M���]n�W�*�OO�	�N�fy��f4b�;�yXl�T��y���v5^!��j~Y�b>]��9��r�y?���o�1^��-�=aٽ�3�D�v8C�v������Lp\C�B�A��~[�K�Cqݬ`�#�	޿f�FkVm4<̌���%1��ٚa�����EC��,�8Bid�ŰDz-�~��z=�1�w3C�󔡹�	o��js5�t�����ߧ�
y/���3`j�1a�~
H���75>�zڶ�x!sZ�S5����}+Y.J���eU哌P(��fͧ��V�S���E��=�h��.��d��$����S�n����i~"���s@7Qb�\�Y��jh�E�&.�ǳ��1#|Ɯ��֔Փ9�߇ds�r�����о��������<!����a}t������ȳ*}��z-G�$ZeH��s��BR
D�D�4���)J	�^~9˷}�u��۞{��g\��|��i��S7�k�GҫXs�^��%6Y9�A�_���{���\�э׶�xO���99�o��.��s ܶ�/����ZB%�ϢA��61W5�A8�	�d��H�2�J�[�S�EI�y��*vuU�s.s7(g�IӼ ���N͕0X)�ivA����'.��)���p�.v
O7����û�k^���8ȸuC�� (f��	K6צ82�`��L8��4����!�_%��5�S�掑lk��<��0�]����"�@A�������E���7Hڊg���9�O=t�/96�O��]	�=b�O�H%�ry�K�{G@�`m���>��&��{
�U�#,U���+`*�u\�+�5�w�Qx�Z����(�T���i^C��������Ļ;��ǔoXɸ��<��k~��G}ȶ��k��'ֵ���&<���l��wfث͜v��o%	3Ļr`����y���n}��h]&Q)�W�Ʋ�'�Ӽj+���M���*	���Y!��k�&+��=�L��&- C�a}�Y�L'+�C���)�����4y����Ke����Ev4����Mv�.��R�T9�Ȉ���]���"�+O�b��/B|��!(o���G����W{=̕=�|��x	�9���DO��Q���k$�'����F]�[a�K�fA�-D)ߢ֩h�FgA�>��u�S6��D�\�xt)I_ҫ��W�4!J�% �PP��������<�ԝ�e�]~�\ŸR��+	ɔ�>(����8�b����],��q�W5mԚ�fL.#h�>�5��	�b��`É �/\�o�D�z%�� �íu�/6���Ս���O��c�\yfY�h��%ڂSl�W�v�|kO��pl�w��j�o"D�����Kz�V=pE�y�b^�Us��݊ƬPPq^�  ɫ����Ϲ�l�dgOEN0�OO3م�Y��v�v���nR�����=���L܄nr*ڀ�'ֳ��u���AWZϐ]^S]3�I��w����T\9��HvA8�"S��1%�uN�j�d.z~�c��jg�-�]-�ڶ�x�6���5�z��5�x5��,��|���01��ܲ:�����*��ZP��R�ۧ�֏ɸ��O�
 е~�E8���a��Ы�:�� H"1����r��oǂ?>�2���1��{�*L�1����%>�M�,���0�� @A�y��$�"K�<u�s_�3�
{^�'�n@�]�a����� ��E�y�i�Z^F��zw�~} G��������{��^�w�����{���O�������E4�����5�,�s+6=���;r[mIۼ;l�}�:��i3j�w泰X�,�X+C���N19'�٬���܂.��"1M�a�+EM�� �	��=7�u�u��vB/ZC�ok^^�<O��ԍ��/_C�V���T�p�
�V:�uݯu'��ǋ��n�WO7Q*V�7��:�������8��X�ՕP9W�7��/MU�d�+��\}(��)�J�HqI�}ݬ�Ά��Ñ
�
���n`U�s�-��N�My����=g;M>���ѭHJ2$���O,�.�w2��4�ң�pR 
�hvr$��B��(��r�̰�k9{�3N�f苅�kl������^�~wX�9Ԩ�"<��uT���r�R,q��\�.M&�/�G$�.b�<��/~�k:���)V�	��]'��6�V�h+tg9�����#7��T�=3~�ʭi�C�D��묌�P�Q�/w��i�ta�u�S�N�p��e�S���܂�t����W	7}]N�kby��Wl���zK����T��f��RT���h����X.n[���x��!ޮv�25��W1F6FΩ[!��pX��y{�j�;c�r�<K2��o+z���*�S粵��2���=4�@F� [�����Pe��l�dof�g5�t�B�֛U�����[��,�x��6��LRк�sL�:�5��zEШ9���D�G���8��I���mgp�;#����cE�Wk��c]��u���G<�!�W�!^�P�U��������Ү����`���a��PG�=.���k�k��z��u�h�Z���z�4�;`A����@Sz�u *^ψFN?1ݨ�V�� T�0XZ�V]�Yxr��Ŧ�{h�ff�]L.;@c�7)h�P�Z;�%�.8x[+�w�b*�-���^�+N��˚�F7]^��L�J�Ԯ9��:����9}��t]�-�U�n��܃}G�-=��7rq�'M���o�^ǝ����zU'���ПC��9õ�c7md!,���YtIR�;��]fC�m%����^�ʰ�|���4�5�B��|��;|�Me�R�&�p��|�VO6:�7Oe���3#�v곅����lĠ<��彭�
+��xk�ْ�����\p��=��6[*�haU�mC �p��Z�K��-���֞�e%��1�9��$K�p���n���f� I"�^��bcg�t\�K�C8ѓ�]�C���l��%���Π_j��}"AG��bod�����<�lNmE��`��nB���"����s't��Ǹp^��:�.V����T4���Mgs9v�Go@�s6�dR�ԹBi�����g
�d@�E��*{�e�Ht��Ɵ,��Ht0�a=;9�c��%9X��2bfT3N:L�<c�3%B��㵯~���v���)4T�Az�N��*"fR���z��B� ���(h�4L/Phi�(Y����N�M'L�)=N�����%#�i
��n�����OP=T���4�4�}����j$�`�)bR����))�@�T�bKm��
��[)�)AC�"4�HSl�Jt�"i�(�
!��t�4��*SJu���i�����DPh((��ZZm�04��҆���iZ����it.��1��4]&��%S��$��N��hCN�(-щ�.�] b�����>�Ϗ�,�۫�\�r�}�fەӴhL���46�PlT�m��v&;���~+,��M���GΛT�e�g��]��� �0 L*�@�"Ҕ�ăJ� o}���]CDsP�0��b���_zL�;㴘U��-B��O6��4چ\�
0�f�"Զ��Dr�ve�����6��s�-��uEs����1'\]�*�
��̦1�A�E�6�!�4�-�'�^���������:x�����Tv�q�j��V8��GoeZ��}ֳ]m=��zdG0�v��W��;����3��0��pپPr��j��ȍ;.�Zηq ��a�n0�@��
�~�ױ��I>�bѮ,��{���z�`<�Mm'i�J\��nto'i��X>�:���]����LIv�2�u�q���� ��P�M�#�p��oF'��r�S]��)
<�x�XP��Ճy��FdY�	�(4�L�L��2YI���,��.خ^����G@�E��̔����Ƕ��ә���_A�+��Q�=h�9n����:�sW�le9n��s��x!0����]��*��P���ߠ����"�6_8��d�)��sN�+MЮJN�~ޜa"�*�X�����|��x~��F�W�x!��5�
n�g�u���I�^ �jG,��OP-�M=��Ҕ%<�X�L���d��m��͢y�5��3�堉{Ψa"��$�,-��\��Fؙ����^12�l���-�p�m��Go]�nBg�Ą�j~��y��n&���� �� o0��fTh� R�=|{矞x��Hs�ko�P��~JBeK
Or�гј�=[�M=�� b�Bq$>�-Ƥ/��V�,d���w����^�S�O�JclbS���L|�*~��ǭ}Ǆ���X-��fܧ�/�λ�o!l�|��^�'췀Ga�_t�N�xd�&�TT�:<�:�r�����[���&y�HP͓�xb���J���.�#0���,UO0�K�(���شv�g�ws�ߕ�����A y?�T_��¸:nɀ��݆������]:]�f0���5_!�+5����cK���P	�A1����!���05���jW��Gdx̖_t�^��ML�~�Yt�3Hd�I�B�;�M�����4����n@|�HHä0��yí~�C���xdmDL�7Â�Սx�W5��eV��zW=�ߟ��+�񞯬�v����|8s
�m��|R��s��\p$�C��2نe�����\T��	���L�uɈ��{%��1a��i�Xn�D�nA����3 �@x ��yO��mC�vC6�d��`�zHzZ��	c���|c;oUp��Hx��{?
;�8c��(�]w5�R��2P&�,����'�8o88���	��ˤ�p���q)j�^Z-h�ΌG��w�q�6X�8��(����Z� �7�y�j�0��WOoX�c\�ާv������_*�,H3
��3 %*P��L���^z�߿��uۯG�Ӕ�
Re���|������[����ʌ�ͨ�t�A���0v����O�|���j콼Έz��Y
�jK�􍈨uY΃����Ai��=uE��U&Ӿ�-�	�g�V'�n'�`~������@t�ݼϷ�i�sͼ4�^Y�?45)f
SW�"��]\����M?g4������]x��j���l�/ά-��8Me.��~��|ǬxT6E;ǰ8��=Y=�����!�H�F��l���f��TzP�NV0]bv+�;���L Ɋ�4��(ΰ�@��z��x/�xܻf��N�A�]-ʝ�'ÄK�D��m[ �����N�j�2Oa#4���RkU���Y1�o�~�x,)�Ys�'�!_�:ǁ��� ���.͔]&Cݭ �'�ۣ���~"S���v����.��c�v�q��~��3��8���'����y���䦝����a��&.�%�"�/�v�Nc����{�NV�h-�Ú��/O���a�B=D&����%ߦu��:����+T5ۡܦ}ft:/I�R	z\�GR3L&H~��L��F��/�=��U�l9��Te�5:p�G�uCj�Z�o��׍�0{��
�V�3��v?J�����l��f��ug�[و\iK��@�r]+��se�uqP�YX��<��Mh�FE�vN�1���8�)5�[K�΀����Nt\ŻF��t�z�s���x7�0����Z����((=|Y�U�T>r�N>1,���M2��\׆�ڑ���(�z�,g Ļ��3��8�u��w)!����&��̝,�\���ƄX�{ғ�^#&�n��L�fE�uTy��	^w�p߸���&�k ��<�C��"=��I�������Q)�Qx�Z�ǧ�`}7�M=6�b�m�l֧���}����!�=����<x�-�/��X�w:��l�༗�P����vk�a��3;�u�/�ܵ��9��tG3��&9���%�aO}t)e4.��v� ��r�K�w-�8�i��#���=�ߕ�Z~����m�ߛST�m���8m���T�hY�MӉ�z}]���2ʹ;��jJm�j��M�	���p�:ۦI�rC�o轠��%�����"�G������f�M�P�qB� ɫ�\��Fu�6)��-Pј{�g���f�!�]y=;���2}�<���{a��9mC� �X렳�V��B2��`��J�W]���^y�_m�^��\g ��"K��L<�6��M����_�~�>���ǃ��{JN簓!��4z�oQ���X�/S��(�AT���6��'�ǳΙ��){[�a˩�Q���/��n"n��u��;ײ�)Ը:Y�vs��ռ뷆G��ip슇"ht�D��l\o�{�r�R�L�{��x���>@� �����$�B��I����{�s���ׯ��? J�F�*�
j]��C�.U�3�rޥY���N��p-�0��R���o��\�k ���|DM:Hȥ
x��ضvEמU��z�#a��a���v���W��b&]�m��u*L�1����%:]�9�@�^��[̸q�pui��W��;���z��`V�{�S ����ǰ�5�<�L�"��K����͍͗����*�"9[?:�C^�:���_�ul��UYi\���7)<�RX�`�yF�k�Ʀ�j`Y���ͩ����7\Dy�q|��W7"��ĝqw�Qa�
6By��1z�S�ÿ,#�est�n����c=�9���8`�~c!���@0���ʹ�~�[����n~ŵL턄�q�;���2��ؑ�4����a �:��a�@9�8/�c�_�����kع'�����Z���Y�:��:���q��;N�&��������Lw���x=E4�9��7�-�����w�,�9�n��,(]�ñ��q��9�lv�[9~�\Km\����u��w��k!9�u~����$��AD��/&F�%M7�V�z ����̂�Wv�ެ,a��X��u�u���4������s�!#l�ۯm[fy���v�Y��J=ǋ�V[g��E��"1$���.')��7�M<��5��"M����>HR$hZX%
3{�w+8�f�f��[���ב)��F2=�L�dY�� ���zB��!���Q�WhĪ8����優=
G:������s�W�0<���V*9�݌îC�U�]m���*�tܩQ���ۍC��ϙ\e9��uFC�1L�6��U(��jԖ�e6>XO���E��u�jlș:��b{_�]�G�4��RJN�~ӌ$\�C���3��F	��#��V�磮���;��v9i+Z�t�k �)����ʖ��v3}X\([0��^P7�Ӑ����쓅�����		�oW�n�����V�%:�%%�j�J��l�={_q�<��g��n&n�9r،%�U;�c@�H>T�@��ƀD��׻�u�1�d�`n�eA%I�s,����u�~�g�ԧ\/>\�z��HP͎���r���J��0��]0�jQt?�V�<3��ق��N�
[�نTr����M(f�~��`&��4(�;JV1j1��.�D���up�Ǣ��;��.�����C��!~:`|�������RF*>��t%�JW�z�z�eҜ�*̿�փ�,�!��y���S��eVz�W�{���1���ZH��q�)��X}/Yu�4R�G��8�K!^[����TΉ�!ԛR��/�Gٮ��L��>�W���-J��:�t������WmΞ���������`<3T�R��AQ���<��׸�][�N���a����9"���i��IWC��,��%��Ƿ!�� !ìW/��1��<1���4�4:�l-]M1]1�,�J��zV�����{V���N�g@A�ܮ�1Y��o0F�Wb�u�����NL3m{#`�1�T��OO�ǣA3=~{�Y�e�.j��P[�ֹ��!��z�38# 9Kߡ�_�]r����w�Q~,���8���Z6z�"Śk �����Aݵ�w!�
��\H�Se�j3], ��Tޫ�el�g�0z�u�6�~}�z���p�$jA}����2%�-�9gjd��E��ɠ׬-��Ov٨k�l�䩚+֤�4
�P�%�<�ٴ�9��u�,�	-MA
��\zY�Ȍ�^{����`ֹSS�/^ܙƢ9:�w�;(2Y�6�v�׳f�ױ���N�]�`�ssB�n,�\jC���3�t�X3�t##Ӣ��0*��W��	M�2�A�PXf�ܮ�`y��n]�����h��d�7*��u���8(8"X[�$>��G��e�y�PN(��I�1-��k�a�;n���bW�����)E
��S��Zo�譊ڼ�l82�^�rn��b}l�p	��v�����R�G6�xxW�����7Rn��v�m�F���3s-9����%�t�ЇSPdn^�	L�O�+�k����׳ǿ>|��nۿ^�����(|�R��Dxy�xe$V�s9�0޵�~��|j�t�R��d�A��<�����a��vOrnxN��N��(�֪��[w[�Tmz
�[] ����#�y��.s��f��JY��1������'��_YP��#Z��֬��6\*�%WH� �)9Y��im�Laz|�>ϘE�A�9�z�RCJ6�7T�ނ:���ntcIuڦl�n��#��P	r�<��f�I����ϧMڶ��Yw�`a��n5q�2�=q dıO`ud�wjL+�ϵM���#YCג��M��Ļ�û3*�FY��\Ejd9[ �g���vOǦD�z�r-� ƻޔ����ɷ���w��7��;*K\��5/l[�rd�.!�.����T:��;}BՅ�u�����4�~����d�e���j��GP�n�`ա���ŝ�����k��~ڣ�U��?�M/96�x��sT�\o1�`K8��y�^/��ƾ�|�Zh`��`q����h�=�����S_"h2u�dF�4]�q�b�0a���_�)��wA��y��j��E���z��[�ߥ���	a}��7���il,·Y���M�@��VV�=	=~OY���h���bR��se.#+L��Ivs��4��	u��N ����:ȇ��VU��4��Ω�)էr��-��{Ort�6��}����D�DH)@f�Y�Ր��H�ˣ���Վ���u���,�{��d����˵�5'�sͼ��3��]��z����K�((G0k{d�f��ۻ�Xa ⅘A��ʸA�1�������I�BƘ���5�R�\S9t����@��I�1�zf�s�Vڗ�|`;�a���kgB���q1�mZ�������*.��fpP.lD�A�'��ڧY5����~(��Φy1Vb_k���驘��3>P뤢���
P�0��d�PꋇU�:�����,�����{�Cș�g%"_sB�*��2����$�b%:�4-\�)ſE���Ы�_�hǮ�v뼳\ٺ9��vt����2��vA�Θn�2�p`&*�t�O@$M~�8]�)჉�7�ƭ�nf�s'��΂h�i� ��L9�v@�T;CH��)��L�"�i�.O#�odD�R������F~�_�K
�
�Z�!�n�K�~��B����Q��.xn�r�ɽ�M-PyflS��rn�\5�OuA)"kq�Q�aǣc��*N�~��tĝ�8�T噢�d�ȊD�8Y���A>��D��%F�P���G�Wu6�I�S�]����K��j��+����[}.�ʣR�!z��v���S�j֣��c~s]��Mʰ��h�r�V�gj�x�c�ٔ�tE^R���1���-ܛ���?O���f������m�L9WK��0�x�c6�"~Wai���|^}CX �����!ksL	���C&v+�4R���~�"�H�F%c�~Oҹ�%�*�a �4�+	t�C���\m��)ߖ����)57�e>��7;i0�:���bq��ћCިx��9��+X
��i5�/��F�$�z��:F0��V�c*Y�:�n��,(]���z�3�lyS}���s�_�,.�F���@ϕ,�|Dby���¶nq��a�̋!�� ����R���!x�jC]��GX�j�^�lk�mẆ�f��D���DfJOSu`��^�"�ן�i{��r{R���up.���p��y��]6?L�����x�	�X}N&.�̿��Z����̆���%��7:��G���x�T��R��p��l0\�C�yg�!64��,��W!S�P뛳P�v̋bc&Y��-i	�Z4)<#r+ON��ǨP�f1���5�~�9�u�_���]���ղ	��}�0
�7ex���%y��Ll1�N���1�]�ټu��>^^��{>���ǧ����}��>�o�������Ek`��n��S�uu��hvu��}۹�`T�M�n��;�|�-6�f����<��F������n�]��u��V�}D�T�ź	�P<7�b�P�y��[C�u�p��D܏���]�׻�5g�E܂wE�.]��@��
��V�������$��X��|5^�i5PJ2$ti)��ː'�a�r�
yT5��O8���,�Ex��않�aC"��J�2�އ:F�{`�=B�S\���h=ZZm�T�ZD�wU��iHmބ(�C��4vQX���q�{���1�ڲ��@s;H�sc��g>݄��ׯ�=[����邵h�Xk~��`v�soA�� �*�)=�7Y+����L��ߌ�:�Ve�q��-puo\��ȯR�O%���8����@��i[�ht��3��'Pǲ��Y6&ˉU��Q��)VF��C"�X�J�+�d�yQ��Zـn\<*Yw�-�iD��iE�w���&#��nZ�L�0[�7�p�7r�Z��:��k�Zk4��N����!&æ^�*-7U0o #����w����d�t(����|*����g��ȭ�
á�0lǜei37zP�Y�����Vw-�Ug,;"\���F�U����&y�`�U3Q5+�������L�	Y䓆jw�Tɒ�2^�{�wv�_q/(�Puw�����r���v�d��=Ӗ�a�w���)��K7Z�'$���%��y)��NVj�%X�Z�fb�j�'�e���~�����������+����o�[(�s�b�FV�sIos�6��u'+�U����O��Z�
�:���<��1����W�9�WKE:��4S�f���,Q����r�ϥ�t\q��*�^�R�3���w�">�*�t���X����C���INɣ��"fCq��M�K��dawn,�ze.����V�����k6E\����ې0^ok�0AyB�� �p�Ǚ���V��������5Du�LC��yyX���U���T��?�</*f�c�"���ƺ:�����9n�ۆ����MN�N
D��dg,a��n[�.,��cq���ղmǵ+al�|�se��ǒ�屮��MP��)���qBh./�ܿ��[�n;��1�;�<2�ޝl<���O��sKS��t�gZO�{�F���jr5�fs5��9�v5�r�s;�f䲬V����7�H>�jVf�9Э�bc�oiw"�,ݸ�v��M��+���}F���Yc�.�)ſm����h��O^XnR����,���ĉ��I��Jّ�"�5�K�`�i^��l:+8vXܗ�mt������yQ3p�2!}}ʱ]��f]0(nGe����b;��TY�^E������j��GHhj{�xnf��M��JZ&��l�b��\�7�~}x���u����t�i4�Bi@�T�&�
ѤҔ�JP����L!H��m.��b��4>z�u	ZM.��Ji4�F��]M]`���S�TkTPTF�:MJ�4��)Z�EU�h���Ѣ���%P�PII�+HTBP�j�%4EN���CCE!�Bh�K�^��i�R��[:uE4��QU5KM&�Z���x�:�i�z���&�%�ĵ�1:vΑ�����,c@L�KDT�N�#k4iŧIESli
MbR*B�Miѧ6#Il�44����Ӡհ������.ۢ��n�E��FA@�ݏ6�Ҽ�.�WN_�QP<�zyj��R���õy�͂a]� 8v��行�j�`Ŵ�wYO�X���fU�4�m�PF)E�K1��!!���cI��Ļ~	�b�#Qt\�b�f͎��3S~S/:����=!ŷ2A�<&	�v4;�;�Rt	�K(t�n�er^��M�Ց���4�Q��u�,��V�3�q��'f��B`���s�CuN4�Tey�E�y��o*iҖiZ^�tݭ��������{��x�@�h*����p��uL��dI��Mx���Aeqي�c3G\���*P����rPX�]&��q.����?�̛�Dh�n�_VOJ�No��B�gF���e� jm�nՒ+x�0��Q��lJ�ε�6��8x܀�<�kxu��+L.����q�W���|���*�����*�OJװ
�^��+�cu��L�X��Y؎����v�2L�0O�uݙ:m�f�}��VeRb��_4gӮLG6Z�B3��kƝ7�VE�v�p�^A@x!v�|/��s 3g{�Q~�^=%ܓX�9�K���lG[�aZ1áv��<1�
�-���ýX@��\<(��6�5��h1SV����2���r�ʋ�۝�Kd;��x<pF�jA}��y��xg�!���-�������e������hۆ�Z�o�s]Բ���y���_��򝷧"\7$�����kں��u)f1d9H��q���8��z3�Tc�jV�}�!�D8J*��y�S�r��m\#Gx��-[���J/s��qO�x������>�o�o}����>��L�@� �4U�B��K�y��O\�o��fz#�[eג�
۔#g/;rMqǞ�!NlM7�ӯ�M��f��!����	�9!�fͧ�z���5����Ol�������nB]�AŴp~/1q��X�+����%6X&Pd԰�'�c�]�@MsR���>�����z�����q}�,.b!�[ ��U�@?B	�/���k���{-���4�흟���p>0{��?�����񭘯�up�.ƀF�<�S֫&-ڢ��C����0�YO�ш��t	d�Ije��A�.P����(fܘ����yc�V�,�)���͔��#ҡēJ�|b����(Ǩ-�Ú�1���}�4[!�r����uM^�j�|����ٛE�=�na7C�1i�g�H%�J�F%���Uk^4�y�D��R�r��)��gd�1,��ud�u��\�`a�^(Z���ҏGs�ON��2]3}��	�md�=1��^���|g��@�P����vd�zdO?�%��E7j��zR~lF<לz���Dqz�"v�v�6��ޞsU�ƆT�E�T�����x��i���?Kz� o�~�����<�'�u�rO��ܖ��Zb��N'���6�����%��z}��ؼ�/6��ٹGl�vqM}DM�]K��=��o������x�/r��m�3_�]�O�9�Pง�����T:�彦E.Q)�S%VR��NX����}���/��O���\g��_N���5�Pл�(�����a}�d�Q��j^5@C��gp����s�a9�a^����j/�ܱj���4G3�
X�!�`��==vE�v��c���T��X�����y�D|}���!��b��?f����:zg
x��۔Z��ۡ�3���i�����q��`�Fe�f��t��1QL�o#.�o�i�Q��؋]�a�9��� �S�h�>B1� �ļ�G��&�ӤW9̂W(5�"��̩�n�V1��[���:����l�瞝��0BO0��L(L܂c����=�'��$�x�2iA��4�leh[�At8����{��95��+����O�fG9���ɬ�n[J~���K)��/����8;���c�`%]\b6-`�I�5�8�.	��u�#��H����f�Ş��fH�&�2f��95W;wC�nJnjЙ'b�%�(�%RN.�t�	�e��u��|+�;���x��#�������k�ӕ���NN�V�?8��{;��Q��ֳo��װ�7.hzb�>�z��S�Ħ9{���F�79��Xt]*��F�&�bG=�"�ə�;J�Fj+��%d�h��}ٱt��5r�m�Y��H������s{���3��z�8�!�e>ۗn#s�{�Re�1����E'���o�g�jY��E[���(�'����i�� �~��;��GjVW����E�z��/��&)�o��i�6�Im������)�3��p�Ѓ��0�7sԼ���Q�D���yg�M����Cr�3K��g���5<;�@܇ǟ8|m�&�p���TW:�YBʒ6<�8�KR�Z�T�\Z�q�­t�)�u�]>�5>�>�`�����#[��Lk���;�f�6�;[P����Z���:�~��`�%�*�a'lN�5~�t8G����Y\��Fn���`̋!��Գ-�;i0�u*�~�׾0�;^&����Hr�^�9/F̚zxW�oyd՞f�!�y����!����,�:�wK7�,	x�c�]���l���^Y(�]1YC�=�X��NQ/����|������1��u3�e⻤:���Bz����i�# ,��Ls�mᖸf����ˌ3%'�UE��^�W����6ܫ�!t�zأ��S,��j����wEmк
ޝ�]F�8$n]�M
|m����pu����W�=�n�\0T͒d�e�X>�44O=6%�<:�`�..����7�M��_fs�=�rrȺ�����eH�3t\Q�@Jkc��;�2��������g\��e����]׊�P��M�S����tS<XG�;�]����#g��v��sf��{Z�jZڇ!k��2YR%%=�6-��)��,��[\vF�WuC&�\;�9�dp�Yq�F��#s�-�O�!)�ѐ�U�B��7"����
�+?~��·�(&gb�=c̐�Ɛ\J|�LGd���Q���Jca�Ju`%%�e	H���m��<����h���ѸP���P���=F?�WW��p�m�zF��.p1�b��^,�\�5P�<M�U���l��~ݯyW!��?-ml3cס0\�.C\���ׅ+�mv�hn-�b�W�l�*�(�gu��K���ؖ4Ψd\˖f����B
��8Bn����m��`��x3�NE�ԡ�W���z����PXǨ.��^N%�=��C�G�:mj���Ps}6g5�UC�`TԽ�4�_T��t���Q��Q��l+���@��'��֫�׫�OL,�6���5XXÐa����ښm�����S�	�X����\��]zKWƾ�>�W���HH�KV�o	}@J��hL2cG%IkU��PA�{���FJ@[v�`#S�ܴ���Hv��t�e;�9�B�v*�����"�jq���e�ˋ�NU2f-��u9jQ���1Mfm�f�*���Yٺ�r�1��=������>�3�k�����:�؇mtӓۏ�:(]�*�OO�L�u��Y�w(�]	��ݑ�zq�.�xņvR�^����r�	�����Q��8�}p��n��i�'e]�Yt8��*+���-^��g�]��9a��\LJ�/{Q��$Wg�����E��;U`�����R���ۋ�G�G.�_E���a������a�~�wܧE鼜D*럻3�J�X�]uE��������h�_I`h���R]�ϯf��E<6�3�ɳ�N)�'ų}�-�_��|?z�~�����w&q�QM�f�;(2�,�`��(��ٴ�-;sm!�e�O�����S̯)� hqms�\zz�&��W;��"Sa0�&+�u��o&�+�{c1^�oj�v��ݪ��Yİxy��"�c�
�dFuYf/a8*k_�j�2_n{B}�SiuEM6�T�5�G[�W=���{w�H02B�.�6P�L����垣-r�6FU�Hk��^u�'��%:��)�$i5��;'���\:�������JY��W̷���?����
�VպJ<����|�e-������DuvhƳl|F����x�`����� %'c��9t!�ѣ�բ:u���M�C
r�����H���W3���8h���}I�p \0	���q�ѱ��}���9X��n��.�MG*u9��؀&]��nH
HޥI;����amĽ�����["o��C��N*a	�ӎM[�����suz`�R/dߞ˙Q޳	���O� e ��*GPFi�e=��M�wr=�8�H9A�[�0PZa��6[�,y�曯�W5��(�W�H�P�?s�QY��Siv�LVg;=�kR�-xlK�@�L��
��y쟍uP�u~5"�Ђk�zR~jV�v�qW#�j�
n�O2�����bauD���D���A~�P=偣���u3�j�M�Z�@*��f�9��X�(a���Yk�K���=s����˘g�g�<��O��ki����"7Z5q��4��";�MO�omTv�po���
�@���:�C˅����C�*h`qGCə�9���1Ï3��{[R5���A���^&h�P�.ŧ���tE���6�sC�K#"�DT���w3q��t��hlcH��]tŶӞ��̳L�^�]��M�\��U��m���*ɫxt����)i�C�bX��##ǆ��Us��ݬi�(H8�0��0�ݚ�z��/s���U�/�K5U��8�t2��T�O~c;/^�df
fX�r���DækU�G�;�Dξ�:͛�&��ȴ�/S>���dK�I�3h�d�)��z��Х]��*J�9�oWQ+YwXr*���..��sw馅9և_l)L�)�;�5~t���z͜cC [9~iw�H�����TE	2z����3 돏	fnKmx��I�^۵��Ad	e@�Z�_��eEÚ��P.E���(LO;wfI�[_�36�����l�͌�E�:���yN�,�j��3�q�uEê�O�Jo7Y=�|1]m��+��͋�	;H��vB�����L�ۘ���4-X�I8�:q���hWo�'M�si�w[t7+o ��i�H8�C��v�ۃH�醐;�Re�c1W��&�֞�9@�U�2�y����j���=Ju��-��#�!�!�'�pG>�ʻCH�%<߉�d]W�9��Wc�܈Og�z�2�漅gf�٩�_����Ð��R�{ƅA�L%���j���#�y��9�-�=r��ʒ��a�;H��O,;����{ʾ�u��{�\k��>�'�m ����e��Z��Ī,-ts)!]k	=��W=�x����`���JYM�}N�:�N�l��ኚ�ڐYVq�j��V8�/ҹ��<�Ҫ9�ןQw/h�U�|+�{"�{��A_�j�WA(��e�@��[w�Kv�MT�(
��ОS=MR��S{q4��~��:����Rݕ��
�	��I��fU�'�$R��ޙ�6����b�cTuӔS�)ݝS�ĺSҞ�	��5�Mb돫d�S���\ei�e�l�����^�Uu��Uj������ږc�;h��QԬ�'
�i���6�j�2��(�Ţ}���S��N��]�~��_�.�1���~!���^TfI���Ļt w(��LIv��]��J���z�z|�iGn����"�׺�奥����&�"�-"�\���wQ!�ȴ�7'%e����]n�YY�Шk!�:��F$k=/w"-�tM�1�63��	��@��I��Qx�׃��ьN�U�Nka#�c+=)?���ء�T5^i�)�P�L\:��L����8���꾼sP�m�pY�+K�MF5��lj��!k��2YR%o�����6�����3�F>R�yA�Ž��OϡC[/!0Y�:v�ܣ&[��D���2*�
O܊�zw^ʚ+M)NgEq��,ܦ^靴'���J|���$+�U��G6�!)���N���2�{M2�Nj�0���h[׈7�Ͷ�m�� ���!�����ƀD����I��RZ(����q�٪ob,�����䔦��+�w0�[[= �6O��^�k�+��J�@���avI�C<S�I�������z�x��޵X6�-��f�V�2J털�f�L�Q�E�'ƶ{�C[�S������~T�(���-�b9�#�*t�/�Iʖf�ۼ弸�|lZɲ�Lm�����)WU��C���'��;�������Im���QI�T��<��i�n�4�;�׏8zh�
��8Bn���|&B���^�M���ݴ|��ŕ��f-?5����2�֜K�w@~��ӹ$Ԯ���"6�7t�p:��!��mH]Y����h]�Ta�Z��Sa]砲4��w͝�0��<Mz���~�  �a��Z����U��-l��`OB�⠗�{
��Ʃh;66���LhW`Af��l6� `<!<÷;���j����_�X�"o����W��cs��W��v���f%�3� y�W0�/�H�W��{vw�J���3F��o��^=:�	h�L_��GǨ$}ÜK�>"�г�O����.77��K���A��d2̛`��t��'��i/��ӱՑ,�� �KÑ�Qp����d%�]�f��P��=��{9��ӻ�����t���{����o¿)�����^���<�����^I�v���u�|�8�4璶n�i�h,�`��(�{}�O�������}��ow����}<}�����|>>��E�ԗy!��Ǌjn�c��S3/r�(��x�Q.􉘁������U��1e���B��f��K��L+]����O�46�N���:��	hGt�_��7���l�K.�ꋣ-�{]a'r�S�,�!r��R�%t.���4G.��N,����/V�t�[t+�]��aR�Ց-�]�N���ٺ��I���a�e��'dv��{����q���TB��U��C4\���K���v�DPv���]�cnC>j�hMKF�+9Ռ5��Ĉ|;����X���楎�rN#mI�f�o*�M�D:�)�X���l�K�k�m%e��-*���{i��v)�7��Z.e�Rn��R����T73[�D��v;{{�g�x^�W�]�﹖��3���G�[{Y��0N�)]Ё<�� �ݻHj5���4t o͕#X�m��w�����ل�֒7A3rDA]�����bu�ܺͮʼ1* �in��OT7���)��eν@aYM+�]b�e�ɢ�������ǔ�; �H_m��X��'&���ۢl܆X8�Ln��|gv�E��C�������1h}�;�ݔ�<�ַW����������|�SY�	7Q5]��v&Nۧj-�M>��k�CI-�4���u���{�g��e����
�w�%.�;1�u�P�I�{+�&�<�F�"�uժ�7��a���@�r�'r�,�	&��GP�++i�}_4��DZ�f	�d=�+�N������ ͓�]՝ƶ�)�c_W����fט����v��g:̎(U5�w�(��H�B��y�V3mb�^ڧMZ7Z�[��T��Ѓ�f�_�ι����J��99<����u�e�PS�ܫ�W�Sn[�Tih��}L�J�\*#9���tE����>�v��hbm����(������,�fh�����H]�+2$-x�����V0�����L��K�p8���Yu�� a��ޫ�~�Ct��ԛpB���2�E�;��G'|�M�IH�K:�-j�[pB�)�yئ4E&i��n�3ά�؉
�᧹˸բ��CX%3*'��ͺZj�pu�od��k%L���\��T��K��v6j�Y��Ŷ�l���ݕZ����y�"Y��H��9(�d�J�:M9&���3�w;pT'p������zq,$�=z�ڥW[�Dy���;�ZX�V� ��\� �ey*L���5���}���V�>�ZA�E,��#�z�˼�X�ޭ�r��W���w�ɼ�����hn:�[1��%�CF�<���)�؄Tebڰ;x��K�36<�Tu"91Q/7�J�Ω�a+�r�X�׌��v�ٛ�����2m���af�k8�;4�(����X�����|��9Cc���1,��P{I�}�7���r�6��vz^�f[���(�b�l��uMo\��7k#5V���IW�>(����־ꂃZ�H�T��u�(�[VJ� 6�AC���Ө�֪ �i60Ub�A��mFڤvΗQkT��Ӣ���h��:M�N�(�E��KC�m�QDQ����+cZ+N��M)mE!��(��iI�%Ħ�Z�����,gA�q-h�IM,X�+qVƀ4i�[j��[*�la�t�4h����ضh����EIZ4klkK�ьX�����M�kZ�AlU���m�F�TPhuN�֭��gF����E�]�IE1b�&�6ӱ�V���&؊"�IQ��4��T��6 �К�����6v0��F65I��:w����u��y����3������h�w����+��Z��('!X�i�GmwI{��N%��H%c�*+2_��V�"����ŴXt�D\zz��ӱ^�"^��PdҦ��y�5��U��O	�S������M<s�[�(8"X\�C��A��\ѭӈ�U)����K���@.�D�粌�+T�5�}kVW�)ZN1�~sȜ������T��H�H��*�
es�s�'�)ծ�L�$i5�׹��_"��?��ki4�3y�T�uո��X�g%3Z�A��K�S�&<սf�>y�Rr��E��,9���e˶?�f������Wg�����#���%��n�}%�=�Sl�S�F-?,e ���<���ڃMZ�f������fX.��{`m��i�s���\�Փ޷{����EⅩҦ���P��Z�>�F�u�6kN"�-f�/��Ͼ��
!�c��.�G��W�UO���tǚ�����nϫg�k�.=u�os`��Xw�����߿T��k���5�}�<G��,������yl�_�E�|j�1f�dm�a�z�b1)���5���;�>���tym�����:>���<�Ǻ��U�na��`Vk<>^���"�q�/�'�ߘ��0�НѸ��[��s5�@I\��U�t[�Ǵe����)����x���dq43�Jv�c���DM��oE.���IA�8�;��lJ�R�J��x�ۑ��KI�[R����)��$��f�8�ӝ�z����h~ա��RNc�G���1\�_��b����̼�t�eD�MF��V�UX\��.9�c���kr�	����B(�����h&8��,�A'�}is0h�Uwk��g�YO�D�Ƈ�E�i���_T�m��wO��4��K���lf����|p��Q[�o5;/k�Yz�<��P��8�F0����U\����cbt�����3�[�D�-vU֦�����֬���g�f�2�Ο=;�.2��y��L*f��;a�2Y�*���g�7<-dzO�~�'X�h(ֳ��{k��s�����sb$���Z�ITlk�6�Y��ٳ����}�� ��1I���Jĭ��֎εQp��3Ϩƃ�Ut���l�f^B���a��d�d9Nٹ.�;!73s�E۞���j��:q�)u��5TN(��N��) ���.�2�i�:B`49�m˷�nt�H�I�1���n�I�zb��'���yz ��!M����L�7~
>�gяS��Wg���O~R|��,�tN��*W������1�ZDP}�0�f�CIbY�^�IX�oi���i՝-�X�����4���o�u�����
����to��
,씥i�M�R�ۛ��6Θ�}��t�v��a?B�X��E��4���rޥ/.�@"�u�c�h�1�]u*�G�{��{�?��f�_t�T�O�VX��� ׁ�U�Q?WQ�G�3�P��Z�,��*ZT���-\��%�a!<;�@܇�`���M��6�g݀۸��1`#��� eV:%k���Qak��IWZ�|���}�� �j�������dk$�	J�й�  \t��T��]���i<*qŶ�A/mj��O�؝j����z~2�1�M�ÿUk��o;_0A�B<��GG4�u��a���m��u*�����;N�&���t�>i":�:_T�6��{�#�K� �<h��#m���,�:������^�����)j�����pju���ݯ�6Fg�;=C���(5D���	h�/>����z���-Uөx�{�*���zTs��2�� ҉�i8"�WD���@vp\F�\H��I�f�)u�öZ)�[k��5��{e�;�O5�6��^��P��Hk��M}1p�)�0A`�;ci<��	�:�q�{聕�����wÎ�}�Zm^�Z��Z��0�*.�+�Ty��ޛk�4<k��>!R�'?~�?)x?bKD��!}%�qӔ��b{og���M��K�ή�3�������*�+�k���%A뚯{l�]�),��hS�3h��hѬ���DI0�Z{ծ%�m�g��n�ˠ��r.:77��'c�h����>S��)ˉ��P$�����Я��zp���.�X�եe�Է58�%626�
O~�r��b�=��C�JO�#������:-�?3���'_(L��vW�i�S�^~t%1��%:��y��׌2ى�.\.a����a�U�qI�ŬI���<�~(	�B~�pF�^�ҳ%�̗l���l�Fn�nY�r9�9M�~�W�&^��Wq�V�,A�N%��ܙ�<���})�4j��b.�dã�I�F�]ye�i�n�r��p���PP͌��p9�KTdݬ*e�lS2��hR��*�����'������a��T
w����`�X������f��0}b�BcCji9�S�QӴ.��0�-Gs�Uޠ��@�pL�R�g̼ǴG<q��6�8���ߘ(�8s��1-�z����J�� OJ�)�z��P�m��z�=��t�?Y���N�;!l� �Û-�P4u~8�;�o������˟�!#m4n+����v}:�b9��f%�3����ƈE�u��C'�{y�B�C)���J�w� ��jC𶮖��n��@�K�g����Ԯ@����M��ލ'���1���B�b{g%�j�%)�s�{�+p̒u7892)G����,��;ul\�w�%�q>�nRh�s���Y�[��aۜ��xp�ܖ�%���_���������	��gƺ�GӜI��^!�Y���4�N#]��٭j��]Q���}@�va�/p[��R3�E���Mg��@�{�~��Zv�n*޹�k�Z�y��!�?K�=.��n8i�/��<U�B�).����i��CS�B�^g4n'9뉟��`ZY���|��/\���CrgRR͜0��,�`����q������wG;�?H{�~Cy���ZV��\�zz��}�D&���yv�K,H��f����"T�{�u�ј�-��׭��
O�D��pH}Y ��j����p*]�4�o=\.�Yy� �RQ,�ߒ3L�R��~��|j�t�C�ύ{)~�v�yib�5�`�9Ct�_S!٪�j��$nJ���>�N�@�It��[��j��\:/�Ԝ�e���,����� ��8<�O���vDA�3z�$�^S���Q���j�g������S�$�1�����Ǽ�h�d���m�{<ԞΩ��tڞ��O�)�%�ޟ8�A�k�n�n�*�4j�f�2Νy#��r�6��低�N�t_j�i��/z�C��Ǳ;J�R�_Bgwin�mf�H�nj����;F�2���r�� �;�=�j"Ui�;�����3D�^aҲ���^K[���N䕁��(&�)[�#nۡKri���������˟��{Gk��qy����E�	Z���|h���=��|YæJX�ϏF�Ԩ�q��Ѱ-�D1�k]��w�A9~��
>����K�m�k��w�hY��i�O�،�y�S�
�Y��-ݛdl0b�H!���v�E�k��{��s5b����ݑG�@�k-{z}]`�sH/���!ۤmz\6��}���im�D��ݓ	b����2}�v��v�pl'3L+�@;^���/�����@�7x�ݺ��W�7�PnL�FxlcO�L~�*}�o��[���������]%"�����WR��A,)�Ɗx��!�E�4��N��q���G�2�3Gt�j����S��Z*��Z�����D�|n���2r�i~�������?ll�����o��AG���Tl���K�� �ԕ���g���U�-���y��,8!'v�ya؟���#��j��Y-!�����j�,�X�4�p*�F���c���Qp�p��,��߅��Lf�D�����2�NE�Mfǈ?��ɐ�ݚ�=�̫۔�_�5s��WӒ���8Aɕ���g4ʷ@��8aT��(.�BQ����kr�)��5B��jVL��꺙� v��ÕvrY�d�͕���C�1Cyx�̋�Z�Q��i�
�&�9��4�[(ɮ��8嘚����^��W�']���y�F��X��b��FD��L)�{�m��2SyS�Gp�v��.�W?Cr�t�oA�,���7%ۄ��M�^~��=��Jt��H�U$����,wO%��*W�]P�ʖj�h4�z���q>�rFܻpi�0��J�,�����ӯ=�P�:��ٝ �E�|��7  ��_��O�0��YP�5�l�kv�aY�U��;�{mN<�L�"���Z^���f�}~p�~S�A�G��&_���z�<������j��;�t.�ޤ¨�R����2����/1��L��$MƱp�������=��ݺ�P��kU:QE��eW�bN���E�]<�UN��'�}njp�=�1֜ܦ]�3�^7-sacw�Z��2����>��4-'��;�_�s��1U�N؝dS��p�{ff���g����y��L��f��m��@��}�ӻI֛zU��B�}ӑ�k�����ԙ����C�p������T�ru}����¾����>���;�,"�R���m���[nw �W\���]�a���Þ|��~���CV��wԆ���}/�a�?e˩�3�:���o���x���Vx&�pȫ�}GBCO+�� ���=A�O;�M_�w4�܏���}��М�s1�S��4����w9�����g��*x��PJfN��<��漻��|.�	톍��dn��x�����3���e�\&`�zxJ!�pC#A�c�N��m��i�V�J<ğ��!̵��/ڳy^�1s+]�6,.�U�mcv1�2	|��B5�q��t�îyg3�ӥ��c��fd5�#g����\! ]�c�Q�]s�-�@jR{[�Ȭ���<����W6�����~���1e��R�y�%6��76���6È.ܣX�NԷ5�%62"ѡI�;Xb74�⫯�,U�w��=���<��Z���[H�p�_$L����أ��MԻ*24&6
��}�9�\)�=PXs&E(ټz��	���C�hN�|�0O#��n�0�HݳBm�x�֫���|�L��D�N�<���������OC_Z$f���L:�0�m�c�� �t��U��.L:�N�_��E��\��7P0i�3׷MO����Q+1�U�L��(G7P���l�(qUeWC՘���9b|�L?5'�>a��zs��R�%4�c�Sx޴)�X��m^�b�c�"��|A(�Y��^�#���2bX'��+}��X�P^g��-��ѻ~��h����e{���E�|Bf��Ó�f�vu��bJ��Z�u�͛3� 2�'s��k�Up ΍)״�-u1	(��]��D��(0t���F������_y�gÒ(�Ta�֣�Ԫ��w=��]�,Z��m���"�zp��F�^��u����U�Qkeb�a@���fGc�Ou]đ�u���y_����x~���
=ʀ<9�x>򁣫������G��X���|�LTr���i�7s9��0=�'��������A%��'���M|/'Oc�1/K��L��A��ޑ>�D*%���/��@;@�����-]b�<;�Ł�y
�
�B)#9��`���(gg�Dr����WB̙�P��,x>��g�����kt�e�:3���>%Ͷ�7��C:BKHC�Za�zꋿda޺���4�}%�����R]û�0��d��[l2��R]{�m᤼�ň֖�&P�a��B��A~�Ưw%L�xeO{��m`5�:�����'^{H��J���Z~���x��$^}��U��د?Ke�l> �w6�)����@E��p1j��4��t��v��O�[� �Kw��0�-_�U�M���/4�-,���We��7X��F��,�����k.���u`iI���Z��š�toi�Ό�b����t�? �B�2Ӣ�T�F�rmtr�`M�/O1{M�Ou����>ʆ��~��R��4�������|�=;���n���,(�\�]�A1,��H�2���ٚ�]�#�����h�0ײ����&O�~�H�U5��=�u���vlS	�����ϯ�)�|1�Z�ʼ������~����p꫆�$;�bm�-��k��!͍0��t9pvK�S�&OuI��Rr�@��m�M�J��8���ܗF���<#����?G���2�8Lpm����TCu��>�E�9�lj��%�2qɻ#5׎��T�a ��a��>�Ñ�$lĲ�:�i�ǻUsX�g��&��=;����j�xC�Bn�)���|w&%ݵ�6y����?G�uؾuvaK ��ʱ���7������9n������O�x��yU�*�f�zwf��� ��ﲪ�0uw���Ե��z�M�T�j���Bը�è�k-{��WX5\Ŷ���P�n��F�W*;�T�Cuٓ�#F��\�:F5�æ�z��1}��A���N
c�G�v�8�sQ~��;�Y��j�2�`����5��D�؂�&9�mK������ �W���3E�;������{}�g�����{�~�w����>�W���m�cxż�ѝ��&�'حگW\��+4�a|5(���:����Ty�CP(�gF���oq���ݦGg[�5����n
�x�̬<���d��3�U����/�d�3̨�n7����WO�q����}��1�����j6��͙����Pr����N��7��B�?r�>�i��5��v��U놅X�陮��ŧi�]]���9w��Vd�wg�Ӣ�y�	�0��cP�F�2��sLi�ػ+3i�0�m��Ӛ���Ŋ����4��~N8=��I�%D�
��\9�d�m�&�������cPx�㘥�� ُ6��S�뼓��]%�T���;f��;�[�
&�}+�Ad��;ۂn�t�jG�cم��{+��z���$��8R�K�{%���{�a�62���+Ʃ���x��7����g��:��ȊѲ;��vT׏b*����L����]�K&��{)9uj�y��m��Wbs��w3�q3�t.m{zN&�F2U۳ypaa��pH8T�+&>��U9Y��^������]��N�^<MV�4SB���qV���էj���$Έ�4,X�Z�J7��qs6��:#���\y�8&v��2%�hܖuLF�H�K*�,�L�0r�z)�Z;l����'yPb4sI4�)�.�܁�
��W�cC{8����H+�7������J�[S�ZջI�Go�e��{�6NL�k�E��+h�f�4*�Wh�
U��.!�Z�弰Ϫ�
���]ΰ9Q]B�/��R���{'}��ҕ����3�a��^�)5�R�9�L�m!��]��D�]O5�5�	��%㡶Z����M�p����ڳh[{y����A*�x�Sa�ټ��(�[ӱ��,����YV�δ�s�#-N��R�u��K ��T<s���='r��KX�T��,��.�jg!է�E>#�r*}��J��w6`;5�����vAs t���\��Fm^��V��x]��YOGD������9tO5ވ�rl�z��͊�c0dl"a[��]m�鳲��z^���+���
Y7 rf�[��,i[�f۷s��T]���ǲ���<�RI�/��s!ljca<n���&v 
�����E���dW{��j�wS���]۩;��u�V MV-�A�e�=QǆQ�o���r��K��l���Ϋ�ia�8ĺy��M��5I��`���Y�2�*�S�q��莍�b��+q�7�q�.��w7�}��Ue�GT�R�鷒(-� ��(rn^c�\�{6Wc7�撾v���cB�.<��3�R���*��kp�L"C�%cM���4B�pcj�9}4�s�c��vDRn2�i�ԋn:�F�m��"⮦%$G���V��΃�}���N�M��|��;ܚ5:k�J���(_P�C�Q땝�����%h��
JJY�F�:�Rb�������Ck%$AA�V�u�F���6�уM�i�ڢ����ڱ:4����v�hō��&��N#A�DKIZ�TDQ�Z/{��M��`�mU6����cmc;cZ+A�F
-�mF6�mZ+gjvJ���1h�h�6�l��Z,��STԴj�lm��lX��m�����cj(������q�D�Ũ�fm��1�j��i��cEUF��*��&*5�%��QD荊J����L�Ej��*
b&b �Pd���U��SSQ%F3��Z���i�lF1&�*b���(Ѫ���f�J�i�QV�J5��""�j"�QQU4�V�,�u���Ѣ&���"�����նJ�b`���Lŧ0TUSQ3O���u��uc�]c�j9"!<�9��b���9�٪���Gs64JX��;��R���*�-��*�.U�z��4J]lǘ!��+��m�NoZ�����>f@�rd����e
I�c8Cn���L�T3]��=w��n��\�&�="�_/�i����!�������z=$?e%�ۼ��?{��f�)?LjS9��۫�]6�#��}kO��u����G�*�6���Ӊ�줃���=��^&�i#�cv�5怽
b��A�.�g���e�-��Kӽ�q����B�@i��-I�5��h��4��"��y�CT �Z�A=,�,���z���Z#pyWe]��!>�b��}��s��t-"K���NӦu�P�����2�%�9C�J����8���f��<*պ��Х�E�<C-���za'ir]�H�SsP~��;��.�E`��y�֤�����Y��[�Шt�z ��D:A���[p����!�wR��ه��P�O/�l`4Z����8��j�+��&�x�֗����{ BF4���B`�#���oz횎@�sv�������I�ʛd]`c�B��6��J�_%�r�e�̐��H���bS�4r����Ç^��Μ�%{��
�rW<�7)<���`�û4nC�l>_��n~�<�)����
c�;Op.ǀ�K�&=O/ �/���OoJ���xs�Ѭ�r6ki��.d�e�}�嗆���t�]�/�HϮ�����ʻ�bF�����nF��);3:���Kv���о[q��L)7���}���������5�O���6.h��`�����ú�����D
nǭ�Q�f�Q���.�E�Z��Sa]k�O��Όp����i�X�[���0dyl���kH��1�uH���i�j�Q+\u��\�⠗��Q��-1(7N��ﻎ+��&mu�J��� -�_���O{�0��y��ls8lNpmK2��,9��ULStV�X��M�Q.�"S=b�Q���vԀ��zyP�W���?�?��C�AKmu��$���n֜"_���ک���au:��y�F�����������+�j��.#C�}���¢�������ÖW&m�M}�,��^+úA!�� �3p=2�xc��������Tũ��GZH���������߂�w9����;����P���W!
Dךn2*G�b��^�����}9�γ/�wbv�,���L  ��L]�'��Ʈ��kl��!k��2YR%=�"ʝ޹�e��-���#�{�)}��	��#�cA�9��G���nj~"Se��	����j��3Fu[��?�W��FG������,��;@@Ŵ�8��S!�>!��O0��R��𡙔���� 5���ޛ��m�Sc��p�M�]����r{V{Β�:E</Y���Q;��!lv���xEԶ�\wx/��Vc��#����ĥi�w2���c\oj���D��wصص�yI}x%���s{�Lկ=ެz�?p�:nGba���=����|X�����,R��]�6o����z��;ćН �O�9l�lӓ<�ٺ7PaT�P@�H�2��/�:��T4�7=s�w0���� H0͇w-���#��]��Nt��uysǆ!��i��)CȾ�.�XF�X��ׂ�P�F9jw�:�ի7nVmCMj�t�DpN��d��BuL�=�����𲫡��^y\�:P�P�a��i:��.��FV {� s"���#�̛Z�p�n�6���58��;T�㊣i��L�z�I�S��/��Ő�Zw��ZΎ���U���M=�?R�ߘ_��uJ j�uRkeb�a�y�msɜ+	�辳��i�t�/a\sI��m�:-���AA���|���������[����n�z��U̬���Lz1���c��LXgc �f�\>�E�F��r_!��Fv�v�Lvr|o=��]V�m��0�t��IzZ��z}Ň	Ɔ���:%��~ˉ���T�u<v�VX ��8��6^��f�, �dn�0v�rC��G.�}������4S���r�����k���XֆJN��V+3�Z �gS�[���ڇ��#D��/:�G\���U�����G�{�]$>�{]۶{;ۗ0G�#�MM��ۄ<6��CvcBR�+rq�z��2��y� ��I���>�f���I���w�C�xg�DsK!��=�O���GGui�i�/��%T��H��:j�������S�t�q4r'��q�PЁu)~�P�}No�S��ɜjԕ3mP��-�,�B��n�Ө�؀˃T��7����}��?��J�����c�$�`�/QQ���%���#bM����ʝ��Þ�r[,(2j��4�F0�y�+2���-bL~���Ƚ�j���>���3wOɧ�P���!��1�8%�t�%�T�5�o��L��߹n��I?\SҒٙ�zy�:���fژ,�����'���:O�1�_�H�T����#�y��.��q��M\'��ָ\]��C�/@P�l��6��3�.�O�$É�I>DI���"�0Ū�^ʽ�Q��[��/Z���vFkל�g��ь"��D&k�f�y���S6a7Cݥ�k]�'����M�Z�~��G��<����	 ��a�Ϙ(֍xr�ܺ[�����w�����Jp��uK�k@.��-@�P��w=��:|�E�xQ��:r���w�����|�WK"��O{����~r�9�˙ݧ^�H%]���i� �̬�\2sB��	$w�3��c�Uo[�u'K9��=�Z���S������` �w��u������r� flr��P�.�G�Km�]�su��J-�8�
A���$t�5�c�J�9��9�|S����ۣ�e�g�w��r�T�b�͵`ޔ�P�����ϕL3f�;�`�`�6��O#����F�q�M��ס������C�P�j%0��Yk��U�i�a�#hFzyP�c�36�^�.�90e�`~mgd�>�.�9�\�[%86���W�v��ss���aۘf�~R�:VK�cPw��vr����<B��R%~����4	x.٬/ˡ�"����n�t�W�X�Ck-��px=�{gR�"]� ��_F9l�����؜�t���[6v�E\�l�>�hD��j*B>�\���؞��6�k�!������E�#�iM���X:�>���Ի��E�U�Œ�T�ڑ����*0-���zw�`��vV��E�*����������o,"*b����PS�X^O�Z�@TkY��qp�D� K�=r�3<���o��G��9��OEk�S���rW=��e�iD�:�(Х~�E��z���J����y�w�e�FhYP��T\<�{g�!���5ؘI�w$p��)��?Bd^Ö�Jt��7��^=B��Y�2.�6�盤S��XZ��Č���5u���� R��VF��i��KlM�|C.g�:Z��J�yl0��V�}�+�w�8�DZ���G�>�s���6�����ǝ�-M��t� ��$�OX�[��˛��W�����Q����k�7���(+B�`�"��oHkj�$rO��ۅ����=�k�]����&f9������1���n�I�$M�|���	��ς>�C�~��G:���ؙ��r.j�Y��Z6� �hU �JO|b�XtA�W�����\� @��$:3�C�.W�v։"�mO����^�T>q��� P۔����+�m&@�yj��Oa(,iq�`��٫r��S\4�#9�cj8�>�L@L�켧;������|U�]<�m]k	�F75��e6hZ���wq�9��8ÇC\0kX�L-�6�<��4ȥ�(��(���`���Ք�����{����`�;�u����z�y������d�2�ܮ`��Rł�=�bPF��t���]e:� 4�{���x����T<��0Mp�	��i���ʖd�p09�u~܄�qp�LҽܫXW�ힰ8ӱ磓��x=1�������@����n�zƭjk^?	Y���7%��aw~�h�#�=# �I���hE��x����@fC���|�A;Ɔ~���B��g�ڋDбVŭ��9
��o:�4�v��u~��;�����C��Ex{sJ��c��بu���/�,t���I\������e3I���v=��;B8�Ú�w���,L\Śs�&��T.�	s^�L���!KC��������҂�_�.=��{k��9�����%Ҩj&��q�黗\ˤ����;�śh�:O,�0w���8{����hʖơ��-{�2��Av��I�Y�5h>�i��u��n�"\tרtS���/�e���9�qN2V'j@a:D&��A��>sTMN0�be\�cP�(�Q{Q���<�_Z�L�J�,��������ޫ����"Y#ړǽ�g�>��-_N��W�S��߯'��M3�@7"2_es��4U'j��Y8���=�De�#�RE�.[&I�?_se:����_�L���C;\:����~�u~�:����di4�<o��L��^�؋�즜]�hf��mw�xjnA�8v@��nnt��������$Np�T^*'z��pˎ�i�X[/J�����U�_�-��:6 ��͞�ӵ\Qz�f��흣�_V�ߝL-�F��U~��^�C{���o lΪ�L���W�Ki���~���s�ս��[��ʴ]aR�0���s4J���&2n=�	�S�0��k��O>mh�]Y��;n^����C�!�-�l�yjC��r$���,�-^�����������K�v�Q���E˺����q�����ש���ƌ����R��+i"j)Tz9�^J}��pq���ʆ�bn�"���������ht�s���r��	�=B��w�����d�˙%����Fc�T��˫��P[Ʃ�-~�j/zz�/����㭐կ���6�܁�E�r۝���k:�~��I�kP�ѱ�/��Ŏ�a<&ن�'�͈{����%�O��AB���R謓��}̲�ɼ�!B�|\���5�fGniJ��ձ�?r7c�A	ک==^܌c�����]��a=����Gi$�TQ֜�]�]��"���Ez@<�bW���&`���w(�\PW�&N��w {2}sNg�TY�4�~j~��x�Ә���|5b��Bsi5���
�e$�.Rf|v�u[�\��\�]n/=�k�i�0�,@#y��Wn7�t�6�k��MU*	Y��OT�^�?`���0�}u�%m~.پ��
���w��K�r�x�Z�99�3�.�/�w%x5���*x�$vE��n�����]�K���G�ޣ��]�/�d�y�8z�S��᭥i�p)��p3���Q��9�[w����2zn.�ґ�z��V������3x��C���l��w���Y4���!p�����v�IJ�r�X޼�ș�X��G:b�p����}ىR8e��6�B����ǣ����#m>��ۛ��R4�z�_s�̜��Qp���l��|��*Gst0��`9��]F9�b�qN�F񫳆[��3\u�W$��]�c�v� �S��7/���[ɯ�~���]+�s=%�6U*rr�o% R��JP��a���-�D�8Ls�EX��m�p�����+L��_V��0�졍W��W2nT�F���7aƌ^��)�3�%�	͐�{�8�P/��,u�6!F�T;�]�����M��֑�G��s`!����V;���3]�?!��X��z��\���	:*��~fpka� �0Y���*��d�l��#Z�S���z��	Z�4PI!>ZA�{��t[���7���{���[1-BJ����X��uq^.�%䖼�0E�NVN�K���d�gu|[:�m���p�I�vl��t60́QgZ��"�L�5M�ʲ�9����}��C����0Z�h�|+:�2>�Χ��嘶�$Z��s��ti(�fd>Rqy\Ԗ��39�{6���Ҫ̸�|AJH'B��>�n��,9�m��#vM5Nl5����H�F��R�Uf����K/�<�TQ�u�u���������	�px�M�����a͢��Cq
�f�O���>��\lyN���T�8�{�W��o�⭭`(B�#�	��mlǟJG�X]?f�� f���l��;O��T"2��u#�"E�U�9:�QSpa�ȷ�GZ�3H؂�$����)"FV�k������V[m��й���zE�+ى�u�T4��m�-�ӱ���%�E����{�yZ���8-��t�
��=]�U]F��%�'yԁ)�z�LM�$5DaʖQ�VF�tp�n�����[2U�';+yr6��)���(Ξ���l5Ǝ��2X8����a��Փڨv�I՞Œ=>oG�����}��w��������o��x�=^�W��D�;�q��X����B4����%��"�#h�l�=5+�����[(�[�8�n���z��]:��L�#B����Ds	8��M &8�lv�dN[��c�r���ww0�d��v�纡mɦ�3o�3��;����i�7���$�[ʠ�D�}˱ҏ뒢��v�VkH0-h$:�0�Q�}s0�Y1q�x1QSu�8ajVdZ%�¯��Ό�+�h48�T��=dS3g&��0�)ql����ub�T��
C�n�t:�Ժ��.�g�+���w{�9�[&Le9�s�j5�@��TL��fLd��U)o��p����X�9���r�=x���5a�2��k��9"j��K
�诡��d�S-=X�K���\�XK�j�V޾���Jʶ����������U�y)>aњ���V�>�vDM�T�Gd�T�z�P�2�Y`p!��R��ʜ��eނr��ɺ�)v�Che������Q�V艨�l�9���]�o���)���\�.nuӳXs�N�-ٔ�N;9�왯�mP͚[D�V�>�V�%���u̩Gew������N�ݎ�=4q�00������/�V"v�Y����d��5qV�I�)͝e�6�{�]�Vto����р��QXh�mTt���z���8��1i�� ^���:�w��=z��&��� �zj���C�n�l�&Q�o�DѮ#,��M�)�9��m�'r^(�2�ۆ���7���gn�yV%H��Q��*H�։ڋݕ�+*Ot;j���|3��	�/��0p���Z���S4��ۮ�X)Z��=�&�y�Q���!�G��Xj�]��E�6���[�`�j�l�b�TG����VK��
`]+��v�*���Z�w�����)��﹎<�N�]%�pϙ��V8��Vh7AR��AC-!��/�::75�n�����~}�������D��N�oc��Fz����1=�6���P�꘨�N	�T��L�`�L���O�ܝ�oQټ��jИY�{�*�i<��p�m��nX�ٮ��<��c�!����r �"�aQbڱ��pw-�Z�Z�G��48Pd5��4b�t�fb�/��
����q�۾X�>jY/~�6lh�TGhG9��q.����LO������P���q�GQ=m0)/cw:�im���`������
m�;�A�5l�U`>�3Τ�m[�m���`n�zn�����z�7�NJ��:dZ�Vih�Ӑ sC�6"��wJ�v�t5l�í��l�2j�U�ms��@�ܥbq�.�7������'���73���*�ۇvesV�S#/!-R�d���-�%j���v�ou��
�t<FP��V4)1J� "#�zs�Xˬ���tE��%wJ�<o�Vl�A1�*N�	A��KY���3������-}IƔ���}̔d+�X$I?G��A%7�⦦(�"*����bт
ղT�[��I��ְ�,0�[h��b����i�uQEQDMhѬSEm�j���U.��E5ET�LU��QDT5Uk$�D�SQM1EMT�IE�Z4D튘cUlj�X��Q[b����(�X�tm
�m�a�"J������ m�EDUV�[:��
�� h�A�+I��jH���5�-��h��#&�:�Q��jӘ��b��
��j �'�IF�E1��$��� 
�lQAF��5���s���հmf����4蠩��hj����*�־��$�?O��SŞ�
��������g�;���b m�!H�p-L^4i��6��6��LDP��ݩ����_+�:������t�g���L����F��n���g#z<���rͼ�q�`'=|�T�Z��?n��U�߽�F���Vt�c7����_1��"��&!�y�N�1|�4sA��yh��'�@�>�ӎg���t�jv`y�����g�6�x��.�Ԉ$t{2�7{�$��%����^_�d�,/�)��f�n2AD!�EN�W��6�0��\y ��!gtu��[����e��~v��	5�����>Ċ�($)�	%��WX�����`�g��T&�?�Y����~��,J�(���ݕ���\��� HזU�ګ��2[ n�����)��Yޫ���x�ʷ
�%�,��F��)J���e��3��3M�5�ʱY6�nuE�ȵ��`�m�wJH���d��p~��5Ӭ�{���u4��;Ƕ������6�x?d��94�\��S�Å��ޕ���/f&���EnH=sؽ�����#B�
�����^t�@S�-c��Q��k��o:��B�>ي�3{��6>(YΉ�J}�L�3l����u�n��ܫi�={s�-��|F�(�zH0:�����rX�%������W%��q���i��e��	� ��/B�	�幸eO�V���Uzp�:�ۑ9��q�]�!��rTv�o�WC���p��D]1�޿��8�M
��B�'nެe��ƏS~`�6~�~���B����އ{b5Ǹ��3]I��e�g[I�#2��C�U�-�AD�XT�&E��O��`G8#�˰��;��Der��5|.R��*w"�{���i;���O�X���݃�[&Pj	�[��B�޻�*HsȣQ�[?E��k���jLg�마�SfNҡ����찇�����B�o���K����_�����j1[T��\����H�j�����ksCB�_}���*�鼣}�wD<5���;����(uG5��f';���Њ-����Ce���	ک����{m!�g�4NSN���ݙ�]q��馮nn�ٗ�L�����*&
����%�A��\�³VӀ��C�푉�S����ݖ|��l!�+������x�k���;,��Xgr���
��#��������.��!oM������o��֘��F��4�*���G�k̬��B�ע�E
$�J�:ٲ��L�e�����|��Ȗz��r�5��pY��FZ5�{���9h��d�ә�bzse����@���i牂g�C�B�(XӦ^�#ͨD�T��AI��ڸi�,�_�<��ˎ�����hBt)�[mûKjF�<@�k^���D:z��������_. ۧ:�!Y�HC�YM�=���RU��?mEp�bn�����|O.�NlǍ�!q�!l��+`��ݪΩU�{ٴ�/��b��R��9�}�*{���-��7�GC��''�m�E���z��b���oL�y�IEx�����k�!��# �	�̳���M�s�/[��<k�Q�'*�7��[�%��H͖�Pu�5�H�j�SBr��ۼ�P0n�p����;�}j��]@���3�Tgk���R*�w��lYQ�}���o^`d��	3�]/G���iE`1Z��IN�l�h���Y��2�bZ�*ܵ�r��������q��O���\�Y��t@�������މ0�hS�Msz"��k��u�����#v�>�#hk�طQ��qW��З�����R����a���z�_ef�..�m[=#�эS���[���q���Ϋ�\�J��Mk	��-�V�.�ɨ�#k�S�Ot`�nZ8�:$��c���然�N���x����CnV�6�V�w(�e���H(���x���ndh�\�fV�<NN�:�޳�\q�$�d�M��]��o��2T�$J\/%`�n��,e7ob�x�a����eۜ��ǁ�<�U	�]^���)f���jQG�l9�)�*���r��"_�5���z1���������ge�w�$���ԗ;���7UR���M<M3�zn���6ֻe�J����'����P�t.�QR䚯>Z�n[��ȑny!�U'69�CH����}��4��� ��"St�H�m�>k���p#/������+��y���h���Ƀ+r��ϟ0f�W/;)s�{hU�;	j��ޫ�W0�=�U�� c̜y��E�����8R��{��ڽ+s��\f�]�eʑqdTw��%�p���p �}�\�EĂ��3X��۵eÝ���
M��}"2jJd8�]3�w����E�����rUi���R���&=����!��&T�W^81�T��]fz�bUGD�4� �q�tq�Λ\�h�(q����M��09�z�̥FmyRӵC��Z�Pԣq��D%����}��1v��ֽ������\0K�d������B�J&.����ћ}��|�{ƕ�
a��ޖ�|�ǘ1h���+p�2rSYR�qo4�+K��z�˕y?NP�=ѳ�pѰ�n�#u	ݳܪU�{p�5���3���6�*�2D���1�#�M����s��lTĶ]��j��r�UIE��{j�j#��~��%���D�^<pSB��`��k]Z�%�a���/�ԛG<�S|[��6,����������� ��h0q�>Q�{��sS-�3�}v��	5�1ӗ8�G���+��*��{��C>�^��	�q��z^ׁ��|�z,Қ&�c
��w�ʹ��%�\�z�>%9�А�Z��;އ��Z�΄�@������G�����"�ԋ#$v�8��F'gˑ�\�(��7b_|c�τ�y�cTʗmt]����Nz�S�Y忻���T�E�a��ժ�&n���]'��7xs��":�RK.� ���әl�Y|,�;=(x���ͺ���g7�����܂���Ɖ�)J���}��=4�u�>E�h��Ɠntν8t�P:����	.�%�t�)������g��k�����$T�Gjx�[(�/��XD�ҋ��o^X�ӌ�=��d�ܞ%[�G�E!��nV���5��QZ�s;�v�6�Kt�ۉ<9��_��f�AY]��Q��m�º,nC"
��|UWoM�%:,�c4#�^(�w�Ũ�}�;��aی��7�Cz?o^�����0Qr-%���m�;n���2�mP�Kh���*�u��w��:9�<�P��)5un��75���3�셓��F���9��{�N������C{���O����'bQ��;Xءj'4
���ja��g{�FqB.�V�%ٙa���N=��A����ܷ.<��ݧ���1
?,8�s޺d^���)�{;�b��Q�&nq��j��5�e>��#d]qw^nT̷W�4jg� �1F�L����I�3�V�s6e�V��j�k�L���l��^F����zJ��ӗ��nkw=��2���(���݈Ӕ����uD��J�������D�sD9ȱR���,��$i�jʶ=�������t+��%]7������h�Ư;?7�'��I�Ъ��E�%Xا3���	�U#fhj�͓�U\�33�6�(����Y�wÍ%^(�f�˪�i����FCD���^�M�6��xw���苌�D,�(%np��PG�.O���eA�1�5mz��k��FTh�sD�}��ny��)PH�Pcz�����8�U�Na��ڋ�NW����M0�T�7�]-�����t�`���t��>��x+�_��m?_\����p��e0�ns��ι�|a�&/�p�̋���dyux�#1�� �ǜ��#����zo���2`��-�Y���+�SL�����7�Oz"�=�!`o\W���f��NV�r�Xr�۵.�ǂ�����=��R\�O[O��47MV'��d�&�[n�RB���6e��m�K��qb�<ërr�c�b��-چn�K3�oh��[TF�x�rJ()Zh1�9��ʞ��-�[�n�x�eP��;����!!r�lܪ�3\�l=rJ�����e�ƳV���.R:3Hi�ZC��;���Q�'*��R)n�Q�UC������d���C���y�@�%2svH��ըU������u<��Z�yӢ�r�$6�(�6�0bS�#���>����Y��䝮�{KKn�s㯶du0SKh�	��u�IUȽuv�Za�r�w����.��y���kr�Ĺ�&�S�|�zfu*h������Ǝ����Q�|{�q���NQ�l[��h��a�&�y01��>�6�
��ݭ�3WT3.�GU�x���! %�*�T��%�0;���E���%��>�}O���Z����w8�S�,���R���5��%SC��/�_@ǝ���j���OE?I���h��-%��si�i^�OL���9[[�p�&K��	$9��e�z�l"s�>{�cO�*ݩ3keL�f�k<�عJ$�J��p���Lͥ�gz��e�.�Y�
jC�wb�[�V7�8K�k��Gr7�w&�__'�s��#�-�È�+��r������ ƿ�����%U.̑�OL���|�^���٩�'[�\n�վ��%P�$T��l����u#�"E��B�q�w|qQuK��{#s,�����a%~n��;���j�2f��J��4��@9Wmڪ߆
i�}���a~�+L-�R���d�� ��d��%�����W�xp�A���:�A��3�;�U]�4���b8��f�=Ɩ��\$:rm�v@}[ճ%P3fA���\����Gp���uy����/ubW�7�lͦ�a��EOj�2��ݨ�gw�4ϲ��c�wx��IO,��-�7�9���)��5�g�kh��K��m-Y7R�H�~�����4����a�	#�n��MD�;l�i�:�q�쮂����Z;9���k�}&���Z;�����{T,%���5fſ����o[M��+����8���ꂬU��)�����V
��`4'-S���ą�j�3&]��M)�bR�ܧ��H.3�7��<�&���R��̨���U"9*~�3��^W�4�c�I���,s���Ӧ��lK�E���uʷ�6K7;E��ö@y6�f�M��f[n�D�Iv�Zm��[�}����ôn	#^_$L�YiK"j{�s0��q��|QzK5N�=b�N�����f]��^Q��Oa�P�!+{�5��ˋ��OM1Q/Cuk��]y�q�(�ƛ�S�sNg�.�Um�8ne�D穠��VU�[�/+�� �pn��T�ʨ^����}R��Y_O��G�}�����ҰO��Y̎�|�]����v���Љ<��e>�϶�׵�jy���m� �@%����|s�RE�.�[&I�w`�Ы+*�)LvS: �F�~�9� 9Kc����(e�c�FW����{�ϸ�K|c�������� �Y";�w:I��W����z��^�/w����{���o�����^�Q����e���岒���c�iȰ�y5Y�,���b�^n�B��e1`�j�i��Y�w`��gu�ہ(<���}V��;EvӃeN-TX��4��	��O;�9�j��x���R���Zss@���n˛���`���}\����=�kJ�v�h$d���8�u�,:�0=���6cC�S)R"��s"�vf�s�Ӑ������SV�WLd����3'��z��Q&a� ��NL�a���R������J�����:���cөٲ�u^��Z��>��¤ZC�h`�t��ٖ�R��%��וmu�u�A��ѷ�K�-K-d���s(��7tw��7Ɂ5��=��:
��姘�#�b�s�q=ͺ����eu6��2q��=̭G��A;�d����!�]2�f`�3��}0������6t��5vt���;���٦���|Q�ӗb77����6�PU�V�]wD&u��j������iGGC�}Rb��Dv�����qg$h��gm�D�]��`�,�ں���e���:�^�
Y��k6���O��)dĢ[���~�C36vxg)b`f�۫%1�D�s�ϱ_@gY��٦�����)a
q��\ R��+8�ҩ��.�y��@��B�Z��o�#�;y^đ>s��2t�nɋ���3n^=�������J�-d����0h/�b��e���E�`8�:'.���_+Kk��U�g �����e�7n�SRd��$(�4�Pa�򱎸����/8T}pJn��7�p��Ƞ��'kf�]W����|:%�vPu�w����%��A�(^��Q|��W��C��6��=;�1��`��Q��w�{M�ifwT]��lr�E:��%�K�W]r��s�&oQ�p��<`췌��5��:m��յ�a���6^R�w�9�pZ�H�w7���.+��qJY��I�w.�j7�{��7�"ZD݂-L�F(PѦ���*/��Eq������--����#_k��w/t-y8�*GmՋ��v��rjY��n�A�v�0�W k8L ��۩�f��`���`.��7�q��wWN�-��t�;$�y���Y(řx����,�e�l�ք�gE�0���[��rk�k{^�7D�
��*���� ��*�r�|M^�����[���b�R�#��p�+5�?��zs�]CV-Z��`9�Ό����q�YK�����v�t��ܯS�P0o^�lJB�Cs�&m��]X�M�z�us�C����6��{[�v32�SF�
%5�Vr�هQb�ړj���KEI0H��tc�os��G<�kV���/e�
��3��2��U�{�����u�tI������e�l��e��ޣ����Ed��wm��*ٌL�rgj��Kz�Ld!���<�%�;5b��TSTMQ:EU�LITlE�
i��)֐�F�6C,�	E�j��b������"�*"�h(5��*%��A��*����'`��A����4b�u�`�h�փQ�TԚh�+ML�UDTM�Pi�m�ADPD4D�F#QU	LM+c+A��(�F2�V��Xi���H��j����%��mE��T�-4P4ST�բ�i6�[%RUU6ƴ&"ӂ*1h4�*��b"I�
JJ
�),⩉cmS0�L��3����"��JJ"Z��ccE[��(h�*$Ӫ���*��������Z�Y��T�Q4ѬZMT�5Zq�h6����g�K��s��[D��7�O�׳G��ة\�n&_s��1�4�F�9%��0�4�}�u�,�N��G>��e�yȸ�LÅ��QK%I|D���P��/��B�Jͫ
�B��o�����>s�W�G/o��;E��eO�$֟�܉���HF>ӿO���0�k߿_�%�$uKkp���+^�]T�/4����&�a[���x0����.�6cuV��Uz2d��2e��P�KhME*q�"�S�{}���MS�`�K�����c���şhˀ��%l��4h���>��:K�����jf�!_,.o7�;&�@w Rg�g �a��䅓�[g���o7c���E�ɻ���(�;=W�0Y�ýb'��&��
����`w�㗯شaR�E�k��	탛�3�-�8�@��lS������`9ԫ��fll˺Xד�Y�K��F�m���[��O#^J��[])ا3��c�
�iG=Ë��]���ث�=2���r5$$W g�%E�ͥWL�e��=P�ّ!>\�s����ZZ���wU�hE�r!^�A+s�w���E䬸�-���Y�ηg�g�靡��U3|N��:�]O/DG7T�Cr��F-�i��ުrbĠ�U�/f[�T�����	�w\	��n�V�Ԛ���*	=u��Ƒ�Z]���>�1�{��g�Ipm��t ���Y���{VQ��Q_b��L.�٘I�bVm��z���S�}?e?x>�R��m@�&R�����Փ~qϡ�̛��ɜ �_r�}��M[<�ȩ�������#bx���-�_w�d�����*|)�箝H`t��~
2�P�w��9�Md�v�SlC�2I�+ȡд�=�	�8�o��B��=Q��fƎ
�F�FYx�IB2�M퀳�'�T���<��sn�;&�mP�Ÿ�j�9y� ����rא+�P�w.�,�y��!�ڌg,�����n�-�+`0Ft�`�P3���h�79���[�WH�n�3/��\��ӑ��{1���IL3��O���
3s^��K����&e�۬S��|����d�C���2}�wӾg๻�t���Y���w
h�h�s�\�>f�BA&;$���A��ϣ��'gU�����pK��L�m��Sj�a\4dx��*x�v�jۋ�Cm��%ɥ<�N�Li#�w���bj���۶Y���I�gQWY�K/~�h}��C#'���J�wH ��(Z����z�9���&tK�V��ʼ�����m�郧%ط��N��O�ҕ�[Ε)�z9^�T�����~1�ļxLu���=!1č������v8ƺ�o�C;ƻ7�,n�̴���� ��mP�:	n͘��{�����'w��A�5X{��f��+�#���*BR�;T�7�3K^[U����\qU��,��PJ��y�^���#"�%z/�9�Xs�S�3�h6�B�Tg���K�D��,�+�惺,C�zѱ�q�c�*�[}뎹�q�|t���*�̞�x�dR��l�HK�܅P$���l�ഉ�����0�y"�&�>P
w-Ԏ̉Lј��FS�����t���HB-y�^�@݂���$�7J�䉐�[!�����;�n����k��f�MC�'߾�������lm�Tex���J�2�XmJ|��@Ty�F\hr�aS��׽!�����C�y�X�1<�*�qtH�Iw�� WC�� f��R�݋:G�����'��=��z���Va��<���Қ���ĝk�Q:�X��Lm�Cq�[����WM�R��Ñ`��`�>Po,��\k&��),ܦ����!�{6�9�F�p�y����J�R�^�ɘGL�Ror|����ZϮ��9 >��ْ��s�o��Sk�;���h�>�����F+ʷe^��`�-��0+�;T+#GP��/}P���};�3@�=	ӛǺ�W�]hl�������b7��x-v�j��ǜ�57���o]ny#R4��+�c;�ѹ�p�6�#�.*mAוTDNV��뱬}�:���zF`͵�|L�<X��#݂z�ל%r��=�}��{����恬�4E�uF�o��;2�w�pD���X��&��7r�kvf�P���Q�t�B��a�'�6������fa!�HS9�4%�V����8_�n�a�<�E�)�E>�M��A(w&�Ls���Ò!�k���Ginx��G��Y�@�� \ә�gS��|�O���f��h��P��Y���Q��+��ya����sSNg���X=��W�WA�V�c<��@�X�j=l�1��]�,��tܵ�Y^#n�9�V�,�/5WV�CE�����J)d�s3�3 ���*�_+���/���Ȃ:�_	6�T9[����/���W��oJg����u�	��ni<y������[�X��Z ���ǽ9R�:،��DH��	�g��q��r
|z�y*R�P}����G�55��V��nv�K@V������@F�"GeRH��N����<By��|��F���U�O��z��Vק���� �/��@�O9��ǖ�� f�7FƓ���} 2m� ����r��ڤ+���n4t�Z�k8v˿gs�Ǝ�H�\�����+��=C��V>=�6/%{2�/0T���m���iP�k�/�N�k���go+KYqmv6���z�O�[ѿ� �vN̕C�L����rZQ3��L����S6ֳ��Ӌ���.����3���#s�Q��9��w)�_�]:bk����T6��7
�Չ� ���-�r��-���z�_�<b��ۧ�%;����HfB�t_O��8��<�0��b\+v���~��_���Y�(+-�5!���yR��⹸��:0�z6�)NЌ�n�����ov����"$P�ˑԱ��W�=�P���,�ҲU�4���3"�T�ج֬�B>ȱ*NU���স	��F7�2$WN˼�o��!�빩�YS�aݡ��	[��o�rN����{%�{O4vxQח��g��u ����x�{H�0z�j˃l�i���ϷyJБȴUґ�Ndd���gvc�.���c}��*z�d���5�i��rGJ�:�3iO��R��6�Μ���v�[��*Ѽ��˫E��u���*��Ÿc6���)�3b� r��%�A���D.�R��jW�����ed69xY-ȿ\oi�ٓ�s�V�E[<���EN�p�ػu���V�7�QX"�>a���q�ˢQ�j�T*���L+����!3dO6�]}x�XUd�z�sh�ev+K�2���ƛo�h�]@��M��6�B��ߝ���������b���^�RA�[z��j*(#K��[9�@��ҡ�׺2�(��
�3�|/;=�W���81�`9O�eut��b��r׮IG��v;������u�=6ﰮ�]�l3���&#(�fDˁu]�g��#�*�n�h��:k�|�SUݩܽ�sU5����{O��	ΠF�����/,.�;92���FwL&78T�207���,�?�Yw���?֋Ų�U�F����?cfh��Յݚ`}�������ٝo.s'L���SKt��dFͻ�Ɏ��z�'��	ā� sz�8�p͟�
=��iP0WG=gL�#$L��(͵��*��W�϶Ge��m���}�t��G`-��-:��D	My���eӦ�׶�;�c���1�:Ǝg�N�B���֣��=��8F�)wg���r�ǧ��y�����tQ��1솙���ⲛV�v����%��)D_C�S튾W�cٖC�q �k�嶹���3Iź^��H����}�vʇ���������љ��PGo��|�!Y-^��y�	>WM��W���A�]l�U����,'�=T�E��#"�RY7׹t�V>f3�N\ep����W�:�T
�s8Y�
�9��� Yh�V���^1��%wq�G<QbGY$���z��I�T{2zi�M2��������{�P�#5�K�� ���\	�o�����ld����x���L��r�8T�R�����{DU��������Tܺ@�J��	�8�]��m��yf�ը�v7:����}v2*�[�e���8ɂN�Z���Sk���`�M��y=u�i�vCo�b���T�	U>QܧY�̡r�[]�9�٣�O��ܧ_�k�!@m��n�GG��Jۥ$H���Uu�wtݵ�%�y��.�Ztz@�66̪�/�M�_��9a�!"��+jb5\�Q[��ͻ�'.rXc���G,��_Y��ģ�^8�4,l�љ�4U&n�æo7w4��)R�����XC� ս^ْ�Q����3��5cwkw�^(��*�r�)��!^�K-��3`0�`W\@��9y!�h#�]��׏u"���um=Ԭ*���#��=�mǷ����ϸ�c!�^�Ԫ8w�2��(�H���q�S�R�����������1� 3���}׸��n�g5@xVr-�����^b�aO����hm��k�e��B4�V�#�� �YgRpd�#}àf[F�+*���4}�~��?�'G�=Ogz�a.�`���S��bpb�� �1��>
�om��������j^��Ĳ���3nTL v�1�S���`��C��t�J�O�SCrJ�!%<�R����Ry�;��ܪ����Jr�G�(�`ޒ[Gj����+���s�hk˩�g�����R6j�uA#�R����Y��v�OL���>��{�m�)����J�ɱu��@����7���6'��E���u*�W[`��74�}��T=�M㽵�s�UB���O����\��3HW\���.z�Uo�i�V��̫��*�*3�L3�������9Mˤ i�'݋� �ǡ�<�)P�C#�3gXE�.�U�;�,�7D�<i�!(�[m��t���<%�����k�����ݎ�p/n�'��r�ưpE@���G[.�}�mvɝ�׷�5�*͝�츴��U��+;{ky�l0�A{�ʍ[�q��H;� �Dm���߰l�l�
M_��$�O����0�K��p{~��=�Ocx�=�	�~�2m*���ϴq<�s��mt�Ln5���O��ㆹ��g韋!�0m�|��,�_������wU�Jҭ���0�X��P�DSk�]FE���KR�|�m=�5�9֨��ؒ��^]~�é���c���a]��Wz�:��k�`�5vD��C���κ_�ln�������EW�U�el��q�2��sH'��r�+W�G�.F�g��NR��h䶁D�)�tȷ��~i�5m�;jzn��s>�z�,��HB����7$nu*��Ô;��e�Q��·�Rۺ�:kmvX�l�0�}�F }�#$,�-�؏��O���g�v:�Z�m�/��/����8#�c�
��%WO��O�պ/w����S�$o0sǇ`�#b��d3�����飝b����ؕ����M�7�wD=�w���	�UʿlS�*L�:8۲c��jYwsl���<-ڨ�	�}F�;c'��0��H��9����E8��M�3v�=|���A�{
���{��\�"������	S���0Mή>�_Y�����#�ߣ�k�?H����煁�T���P+��:��0�U����U�F����z��d�U�V�EX����.+7�^�/G�������}��o�����~3���{���T��>N�x��"�xA,��1�\�� i�''7{7�i�eY��X���v�Z\hA:��}�ӯ�o��Ti6#��x��=�Mm'O��^�ti�*'�*����Ճ���`3S0����u�3��vh�]�7���8��pW�bshS[j���G_tE]��fZ���!3f64Y:I�.1��fQڝ����S\oL޸.��)}b��'���$ ނ��@f٨N�{_+o�x,�������>ْ�0PF񣦺ڭx�5r��}Di����]�2^I3�����6���n{��a4}增]�7�Fl���q\g]�(tЍ����"�&�U��Y�8y��%[���݂���Nц�s�tFw-��Գpj &�\��Н�0b��8����3.v���b;��E���v3Dc��@�;U��Q�/{kv�/�TupJ��٫)�%���#��oa��r�%]%bލ9᪝�|U)x�	N�\\hV�*k3b�f־�)��di�@��){����)G�P�}�ne��5,��1<F�����xܾ���k�E��,�R�#x'w�1�����9�ޞ�F�S/�P��q%����8�#Y]5�fQ��Ɏ���Y�KvQ�y["Z)���$�8҅'�
������ll��-�r8�B[x��Z�5f���b?Io���M["�J�&�1�7�'ʘ�v��[���a��P�����/�
B�(��yYce	���%�}n��B���IJS��!�9ܨ!8Σw&wJ=J��q4�\���&�.ڗ��_��۠�8��gfǸ'���HU��Ox3��D���4ɴ/lX���vT�3��p�jzO.�;M:7RP�O����Μ�n�gp�0�w�4E��i2�W0�O���f�/�&'����q�I���Å�.�t�:�.��F�:ܠP˽mS�/
�3HN��נt�S���;��=C6mne%�_�p�8�v��ٮ�mt�'oUӴ��%e�	�(%�ǒ��Q��Z��D�R	v����q�8����!��wh'��SH'��R#a��L e�sxw���0'��ir�j���.��s��n^k�E���D˜�t�u�6�#�E��EQ��0�\{l�/��ZQN�;n���M+��w{�����╏�t��7ml�%�"":�;MU�d=���A�]E�����2���h��[��|)�\�=2�m�/-�q`�kU``���2���\��"�^��J��2b��]]�d�ݦE��h��[*���X�Z��DIƶVY��)�j�/�;T�ta<���ev� ��z� 8@��ќ������TԺm�Y��.��K,�R3��.�Ϲ��|2���A�b�
:��5ێ���}��e$!j,�2!KuXҗa�jP������:ZmF2e7Ƴ!�]v�ر��2��0`�ҹf���$�t���pw{�+ВڟsP��� mI�Z�
���!���i�.���BTf0�V�N�b+E�4QEkIE��ADAAJ�Q%킋Z�$����Mv�E�JU�E�b����*�4i��H������((hѢ ��J(�iu�CE5[:h��v��QAEEEU�T�Et)IZLCA�%kE!EDD�Q&��j�j�()h�(�Ѫ"�"f����F���"����V�Ztj�h(	�F��Th����DDZ�E�KAE4�@U	QP�0RV�Th53I�у��ֱ3%Ml:(�֢b��-�N�PTKE6�փ0�v�?��Q-���5�y5/jY�%��5U��u)�h3�Z�����T,ʹ���� �d�ʋ�/����m��>���>�&�{�IM�V_�����cП���U@?\{��ipEg�!�zp�&̽
�1����{�����Ғ�ܸ�����.�l����T�E3��q�i5�~Cz`��;m>
�TR4�[-��� g7�Z_�}9�⨭�7�xu7&���ё������-z�%�E\2���3w+���.�����m̌�EONz���&�x�^۱ƕ��-�B��1B���M�꣺�{�ߍ�F��?�y�ن�8*���E�1�z�a��6i����Q{����c4�P�+k�wU�졛!������๻j�.!F��z-��a&�n��'�l-��d'l�Pc t3��'Qx�3]��ۙ;�iن���(�����:ff�<�6���K�o�LJs��rD���ړ��3K7;B�#���V����Cϻ��1Dν���.'���56�3&XE�ŌY��!�,z��j٠�l*��6�$�X���o4��Ó��(	��lk�M-�A��U����(��h�p��b����4�:��.�X\��E�T�2���E����἞���ڽ�5�!���n��s
+�бc��*/���Eߣ�����L�'!�ѯL��{2�Z$uz��L��Z�TE�ݮ�s5��+0u�*}mӪ�ϺY���=T�zf�><�)bs��k��k}&v�u����3�vǈ�2���m=qQ.g �Üw�q�1|�g��j�������HG.H�4zM<���D��3�a���X�����U�ꓝ�]�,�#,����jH�I"���S�n����m��v��s���$1�B�B6ۄ��n�FےJ��*R&T���KGt<��~�|���˥��!��K����*��]z��`i.Y2�H\��(f��]r����x�.��c��@זP�T���3�;��"!S�vI��-�{&w/����;\{��R�	a�����2�ޡ�%5!}��.�t_R�O$^�Ǖ]�(*ݕ{,e�r3a�ߜn�'>ࠆ�AMm��y{G\�"G��@��cKC����k;�P;�Z�t�@nP8n�b��]j��z�8��IU�5�gj�e�����z�4B��Q5�u��I��A��ژ�@z.i���fvE��׻S�S!��j:�Y|����~�苍�v�gq��b��K�-4���:���R�] -��-����C�����޺h�A�Qp�k�H�~��i���#��*m�c�[�^b��7g���h5��p��/�d���0dm�4L�<X�����	��U[��/H��5[�_E�x�+|��xwxt�d���f�p��ls���k�d��ߓ	�k���Z�a�)٫��s�d��z����e�5�s�:���{���ה���]��;�H�k�.�\���elKvk�'8���ۋ����u!]Ǔ�E�)��9���&j^�).���ظW���(�]R�7ʄd@�!]w$�a�@B9'n�<�lm4]`Zj8�a\�fRI�pW�r���"Gb��y��y(Շ��4K;Ihڜ�@�^s\��c4� +���u1�ǺW��b2�|AY����f�wr�[T�v�9��r�v��e���2���A�����f3+\]�՚=ҷ��s���3ʍ��Ξ��5��添N!_��������X!
B�N��;U�E!�:(i�:�F�t|UX7;��&��Z��
S%[��#�_e��Fv`�~���z"��`���\����u�&���aq�����j�zKlC��J��a�L���},[}RA�pX&g���:s���+�9t���Ek�=G@V�2'�F`v��a]�n�/-Yz[��p�hN���v��(�
X^A;��8�w!�xЗ�U�^�n� ��r�zvgMtʐ�� ��r[@ME*�-�UQ�j�F�?g=q0A�� t�7ԇ8#�F�h>H��T-�|8�ϗ��wζ����%��^�)X�!�=Ŝh�t��frB���m<�1��C�y�_��q{�L�ݝϹ��}#�_�Y����:��LYLY�����o&e���#��������D�9�s��66)�r�	�<��H\nx��nvA�z��]bU�yF�\]����V|�r�*�O�)��z�z�D��Ȇ�6hl����X��3Z���՜pˉ@���$�gr�ɪ��$|+r�o�Jb���_Q�<2n�r-��޵2n�Oo���JWݍ^2P�;F/��t�6��Y�0+#*Fo7MI��4�'2"[\L�۳%�o.ݾ�� �5�j�hL���Ƚ)�rx�TQ֬qږM�6l^�ˑoˎ#i�,₻	Xw3�VM���B�₪��x������몋\b3���T^M�9�ASB:��j�f�>�i��n����Ή{��=.9%Һ�Q�B��Z��U��)��E	�nζ�\+��;H�iw��M{�	%J��UA���:^ɶ+��0q��V^�ggL_l�`��U#s��
Z�m�O.�Nl�X��ޤ�1�^�__hO/�H����F��Ͳ�}ZJ���a���|/����=�ʹb���e��n�O�����C�F��.��5�_|+�Q�;'PyV�0ź~��9X��Z��]����#6�q��Ԍ�\�eu�ak8�|e�-=�ё�K���{`�JP��`�<��O�d��
Rg��~���*o=��P���j1������E0���,ؘ�q/3{j��>�Xφ��\+9�����j*���B���7�1�u'[c��~}������7�]�����(�O�*s�}�rJ�#Q�v��]%�8�8�R�[t�d�A�a�己�[����n�A�&՜�g�e��`o�o�������{a3u��7^u�n���Hm�t��v-����UŎω��P=��k���s�L.���"��Ћw��(7M�.ҽ�:Y���y���^�E��N�B���]�s>��l"a��@Z��u�����C�q"J#�����;}�h���ٚ�b�;��ǝ�[�����g~��#Ę�ة�{����3tq��Z'����Y�V�GK?�j��Ozg�z�T:�t3�]n�������d�&Ԣ�6��Ohagqb�*�g;d�ڇ�ݛze�Q��!�W�*2=G���:fO�i�i�?ݑ\���q�~�Q�'�
��mny��o�b���{ʂ��+h����ͪ7z�Ż�_n;yۙ�W�(�\���!X�n��7`�~nI+���_��u��g���A���^H1��H/�r8E�ܚ�PG�1w8�QL�o-QT��vE�v����t��~�ek�v]2�{�:��9���@ wuT�T�Â7s� ە���S��ԋo}/:��.����vٵ�8M}�p�s��9���V%8I����」u-��b�n���p��Cn܆�u>�C.�AfUv��*θ�ׯ�_ðh�{� �^n�7# -��=<��L
�~�B��3�7U�6��=�s\�3�V���iRIw�K�8�l��]���x�t����l�h�m��M��ܿ��<��r���
��|h7=ևႀ�=y��]p[&�F��r�d���RN�NW�$ҽ��-�é������|�w"��Vo;w�!g���p���e�&�Ԋm�\c$��g��TI�l�<ڝC,6@���0#�/�d��`�\hd�BKͻ�zSVhF-����vu\	���}a�Q���{�C���a)s@�;;�۝����=ȂK����7́y�a�Ԗ�YdLe���{��l��!�*���nϋ�\zQ�rm��=�6�p�>5
�Ed���<lmN��G�#�pE�-&G/]�r�i����E����Yo���]v�#�Q4���ˮu�{ڣ�����p��m
&���G35K�9�
�:�#Ĥފ���f�P���o�B�u.��0�S�u��ƛ�6��P����f]r�{�l�R^n?a�~]�iz~��ڂWK]�"�Ĺ���ﱐ�7C�ut�C"� hހ�8O�bU�Ȏ�׻�U�U�l^�xX�<��TC��9���ݫ6-���@97.H�XD�.����%�ª����x[-�_�5.q����y]L`M3�7���J:؈|u�Z�򎇝#h#9q�\��gk?odq�U���k�R5�ȭ�
/��-ƙМ���l���^t���P��k������aH*�i��t�@S�n�s�����)�2�O�אz��H�\���m,/X@�iVޅ�T�����(0��Q��l�uv�������k�1�L5WB�����]hF:#���ٍ�
�z@ٝU�)���r[@�j��]��v��*(��ٯ�"�܋���w�X�8�g���>��Taj�x�;Q�W5��O�v�ƸV��8�����&::���ݻ�����Mt�tPL�x���W���+r��h^�����9���ԺݰS�w���(�(hK��T�K܈����Ż��sg"�/�9��r���;u��.�]�	
���xqa|�m���4nu���e/@N�Q��4�������m���fe@���G#nz��Y�}��~�K��1�[M�k�û;gce��\�����h5�D�Of����;�`vZy��#����(Φz����E������:^�z�OcΊ�7����wD<��JОE�U҉y���͍I�w8]����|O�&#��ޱ$�@��IQ�Rv����W�˳i�el���,�ła��D+&�\d����'��hSR�r�V����ލ�;����nM9�A�AO�\A���5j�2��lʹQ�{���^0�$rK})��tc۽T�i���A�0�X:!��SQ �@�k	[��.�F�y�� �J�H��뎺u i��0z��_"(6��bzq�h������] ns�t��7.4d�˸�({=����U���j-?.��|��ǎ�e"�Ajz]����������fg��b�h~����[FU��V�h���o�X���Mv�U-�ޗ�=7.W�x�\�̑���%0�=�";���a�޻�hk3*�[֎7n
v�w���۟�٨�\���<�����.�vDpء��m���TR4�[-�~��ow�Mf�[v�n�-M������L��f�UQ~;?0��o�3o;z�?U6�m'�H��W���4�^<���]�lt?�d��o�O�ZЖ�:�5O�f�c���F^���3d��
=Wr��L���[���G;h��+�ռ������쭰Ӿ�7��]�{�f����x;�c�q���y�u�p�g��*�Ŏ�1����1�'+b��W�:����+�N�H-p��h=_���IJ�p�p�#�5��s�X�+ƫl����Uff��������G�>����T�U�{�e���O��;��٬ǚ�M�6\X>�ǎ]f�b�H��G��gؔ�d�,�S�s�^b������i D&�ϰۙ�:A4�S��>O��>���M��E@]�`�/�?����)E���c�c���>�a2���  ̫0,��"�+!(�0,ȳ*̣2,ȳ(�!̋0,ʳ(�+0,�3"�2,�3 �0,ȳ(̋2���0,��"̃0,�3
̫2��2,��̋0,����2,³��`Y�fP&E�Ve�d$Y�f�a`Y�f�eXi�fE�V`Y�	�fQ�`e`eY�f�Fd`Y�fE�w�=�S�,³̋2���� L�2,32�ª��0�� bQ�"�C�C* C �C*�C"�C�C( C C( C" C�C( C  C�C  C�u���t8Ҫ�a ` d e eUa� !�U�UVUXz�( C
���0��ʪ�*���2��� ��B��( C*����2�ʋ0,ȳà��*̋2���(̋2,���a�zE�eY�f� �eY�f�N� �a`Y�	�f�Va_�x�샿�1���U�PF�U �?�����|y��JZ�n��W�����/
[�{��t.�솼 ӳ�{��_7� *�'������T���D@��C�����;��~���}ԇ�E ��c�}��>�]��y��@�О���? ��W�c�DX��QDhA�BI@BdT�P&@�� $eUa$UaH@@ ��U�$ 	Y@D�U�  	FUV� !	UX  � !! 	�P�H@G�?PE���_�Gڟ�QE�DZ�V����_���>��(9�>���?Q��� p~X>�ù��G��y�vH�@��v;������?(������i��1�ԞaW� U��}�>��>��J*��o�>���B�� 3�~���;/q�'�pnwN��=�<{@v�( �C�Z����E ~���Q�?�~ϰ�H���}a���	?���G
�
�>���j( ����;w�;�'ڽ������~����o�{z���I��� *�OP�|�rd����������O|_�ET�G�����
�+�����w�? �}����e5���wp�՘ ?�s2}p$Y��=�Dm����ٶi*� E(QE� EM��P���dԶ�!�ĥ �4Ʋ�-5AT�C$Z�2�(%-���-Z��6c{:W,�d�љ��%S[l�V,��Y�YP�-����ֶ�[RUZ��a�-[i����P�i+V�V`�R՚cmZ�j،ڣ��)����YU�-&�Z�D��m�fi�2M���&��ZmA��F�hƓ,�kJѴ�	�U�lX[&mc6�����F�U��<�U]kX�l��   �^k5�kmq܎�[N�n@�h6q�ڶ�5�+k�éU�i��)J(�.�Pt)��n�:h�J�ӫrIR��eÇWo��Ǜ-%e��5M�M��m|  �p�*�CCD��4/;���S�CB�
��|��GС��B���G�(z25{�,���:
�ZVQKB�{;^�4�����;[�ҩMj���;[6��]�%t��VQ���4Y�0٪ͭ�  u�"��B�r�E�m�ΚH�U:�m�Ӫ����*�ғh[}��Nǳ�(ж�\��4hۭ��;Y���gfN��A4��X�V�f-�����7�  λ�֕�U't��@���S�4�۵�T�і�wvm��R�p�涃n��*�W:��Z_wQ��G��v�(�;�J隵a�������l�¾  w{���	��z"I�n�
7v�uUM(#�i�Sj�ê�Z�� ���c�^��{r�����A`N���mZ��������  ��t��p���u�P&q�z�ܷ֞��H�� �Kt�CF�m��u��׎�
��6]�hs�a��lƪ�f��)���|   X�������E���#vp)]�ո�2@ M�����4�r���7x�.�kx��Gx+�mY�e�dY��eel�_    \�  z�F} �N�
N��= y� ��D��]wG�� Q��U� M��ր7N  �ޔ�e�5�V�٥faUt�  ��@ ܦJR���p= 
.���  3�y��(�{ײ�� m{�z  ��q� �{[�=U��{� �n��D���mi`��Y�m[_   u|=����]�w�� =���z�ޗ��C���pz �D�tP v�Wx {��otp = y˸�������&2�T& CA��$�����zxL��j���  O�����jm�%*  =JD��R�  1?���=�g��;�O��7��_֋�9�����
T�;��g l�ڞ�#?�{����������������%�߲�l��l�)m�K-���d���v[l�[RKl��l��?_��~��`���v���n�/�=."���Lk��7;���F�"}����͑�&^i�u7�)qh�Wvn�Ct��.�2��0r�ׁnh4.�w%���L�t��X$�Rƕ�+��S/�-��ۤ��Hc�q�y6�e�]ee]%f�N����Tt�V�j'X�Y�ޝZ���V�#r�P�D�:��1�
�2��{��D�LN��r�m�[W��0�J\c7%"�<��̘э�R�Ҩi�F�"Fea�O(6��̀�Сu(SJ�
�{
���Am�O-\��Y�u��!x�@mJ�^�R1B�ti�c ���^Y�kL܊�BW���tw`��F�[�h���%�	Aɻ���@��(�օSY�+�I:�>�[� �:��wy�>�-V1
T��a,��m��U�#�j��cF���{S��^Yݒ��7\K%flXvã5V�(��/u+j@٦���J&��yH 2�C(c*�K[|zx��s��Ђ�q�buy6�g��o���hI�S5��H9��zF�zt�h��cHB�X.�!�� �*�zL�%�I"zڼ��A	n��h���{-�E�����TQF��X7eB�.J�^%��q�n�v��k&Y�)i��4U��UM  [���x�/�`�Jϝzh�
�Am����G(�8�9u��n�l�/��XQ�&��v��pCnX�
[@�2n ֋�V̤��]�"�J�-t�ى"��.���<�yuԄ��0�,�q��7[Y)�kF����!V�-Z�@�Rٴ
�Wy �p
��n�n�Y�x��8Q���m�6���LmũS��ٹˌ��J6�-�%��UϢljY��+/ͩa<TI��wj�^f�)#x (jl:	:��)���G1�\�A��������p���S�-P�p;5��)-�FQ���Īj���z�T�ae
�AKP�#���[0�r��s�.�df�<H�n�^bz1���+k%A1�7�9��%�P!����=�1�"A�f���,f��!Z��j�r⧔#�d��IT�El *Tn�km�*Sa���t۽����vb):8��˭O�%)j�"+,��	k��q�ݖ5��t5r#�D��t+h�Ӎж�d��>���kP�%[�:A�A�l-d;�n-�-���n�S�*bW����TP\���ƚ�4#����U�jJ6�;�U5)6lBb�w�Ǎ`Lލ��nZ���t--��y�]$�ܷbmZ��}����*$��:w4�y�!�ڬ�����:�h�ފE�U4�nJ5{�խ�b�����f�[����"ܣ��t��g]�1�Բ4�f[)@��=1R��y`nX*
�VD*I���`�вIv� ͸%H��ө��R�ռ�H�K��`�'X�M�IǹV�T��ױ����t�m!��!�uk�Vi����4���1�#y���uf8 �������r4�yB�)k���p�?���-2��oN�Sa�x(Ck,]m��fܫ��0/LT T�0�I�s+1���c�^Mxۉ�5�l�a��h��h��^L�j�6R F��*�
$������ ���{p��P�e�N�i�n��W((-����4�������V��73XF�lEnb���
��db��|f�v�Ӵ�^P�hM�E�J�F���z̽���B�ܠ�Cj�:�3Cǯ]�8�b�����ղM �e�Y������f�q��a��F��(�����L�Q`�"�`�:m #$m�v��ܖ�u��h�u;��]]�WKv��bъX������h�'�`����ٻOb*�oE:Nx<��1>�<��=�FY��KV7M�
�7pl��ג%W����2� �u1;��:�<��-dpi,�4-�W{��ۦt��ZMι���(�
�Z��0�ލ�7R�b���()�:���F��i���n%GA٤������rh���S.��r�	��5�d��Q��M���
qJدj)y��]��A�.C�ӨP�/6`�kd����`Y�wi^ Lz�weT�q[�Nj(d� �{kvj�2�a��ܲZT�eS������y%�6�8��U�Ճ6I��$�ȣ��hQ�Đ:��uEx�B�Y�W#tJ��� 6޳��cr[F�7Y�A��[��!��(�-�pf�R�y�]O[=ht�:��E���4�m�w���a��:�A��m&�h��FdM�K0�J[�<�ɜS�MSg��ѝH���v�,���"�Fdˇ�����Dp�R��ע�73Z�ى�lB&�iyQ:3b�EZMSW���z�X��X�iS�M�a,�-+�^��n(���K(�L��Ǧek�X;f��K����݂���������q�u�u�i�v����Wha��V�z���0ڷWz�֤�N+#�f��Wso`Ʀ�������2�sU0�NG��9�0-y�f���~����e� ȓ1�7R�ʰ�K�I�	8nẁ�+t�v���c ����W␝��n^賭8�頡��C,E z�֝hn+x�[Ev��X�ɲ�j^d��o,���.=�kk5��ۧ2��T[-�ͼ--"�2�ܤ���5�JЋ�������T�V�%�ˬn=���以FS͘	.�YNԶT����tn�����Z���crHV'6�V��t:(��cC���a`�z�G�KCJ�8��ՁZS%�tAa9���{�����%d�w�0ߢ$E20�j�nӧ��%2�Y#F���Łk62�<)H��#�z��A�4EA�0Ka�ַ�%��}����t\:4�u����Ut�D!\�Q�
���vw%$��f�n�C/:u�1�V�+Ƞ��^�-���։��m���ځ<��#B頌�e^�bt=;���3���h��v�$Ч��+t����z#�g�i�a8��kq��&U�@��+�l<5�<�-�w{�r:�>Y���E<'^�ާ���c�Ae�3d���b��v���C5J�are[x6@�!����q�Z.�t&�ѣN1Q�J�6�[��i;r(z�o6K{F=ò�VT��59x#�]jA5�Q0����Q�D&o!��|PH�� н'@�����V�4GB-��Jґv
��E2��D����ŉ�����h��kKt�N
�-�n��]���-jNk�R)��� j�6!�u��7a�q���~�Z;q"v�Dԑ�Cj�����t���[LSߤ@��E'.P�~%�l�.�i�.��@
m刂��oSo0�K0U��i&sM����'G7(f�N��&kmH�&Cb���׃N�Q��,\���0�ׂ�9Aڼ�[�P�����v�&CF�0�xP�ݳF
6n�W��`��iI�Zr;3j�;�F��M���p]�*$6�4q8�c�*$�$�//2����x"�CĚeح��9x�:��m�hcG,G�166)�%�l%�^e�7��V[ck^�p5�;�N���D�2^Y���5fli� ��7n����<��jӦVV��Gt��g�5����a�=8``L'4�
Z���3� �oD|���b>�|�H�[��Gy8P�)tc����t���J�^��Z�����°��)W�X���+S� ��%�a��MK[&���I��M&�Y��f�?������[��ݰ�о՗B�C�$WKn�A��@	�92��i��xh+i�6A	�JS��Q�����2�a�7#R�F��W�N�[Ϟ��7A�p	�� ���SQfmò���P�ug1�ݽe4%+�m�AJX����W#�R�U��		xO��^�y�A��	5�n�2��:	!x*e��2YK�=6�?f)���j�a��/J�))�]f4��#���m:T�[SeH�o+q��܊�]2�B����莶P;	���j��hv��WX����Z:�)�fS�K��4Y�vF �S*��Wk�q�*إx+�#�Ќ�JVNE�r���KS>�A�oA�Vb>{)�;1�% �6�t��z�8�]��Yǹ(�M�ki�wZ���:0VF�Zu���	�1D�R�7�	r��v��\��*�nb�k�0��E�!!Y���E����+�fٶ)�(���N�)h�����m��ҽz�D�V�,ꙬJt�K�����%�W@E�G �p�K��ջÛF��ѓ\O�Ħ9�b������<g-jVr��^�j�x6�m9Ӎ:ږ��@��^��(���oU<g̬l Qzv"�f�v���ȣ���԰�8���0��M���ub�!���|ڴt���#{zv�e�h�9XO>�_��\��g��� 9�^E;5��\�E���33Z� %@jm][GRz����
b�܏l��>�Cv�1B�t���h�ȸ�zBKt`�Ⱦt18�+�CUb_6Ҹ�sA�a{)�l!�"N�wl;����rּ��l1�6���.F�n��,)[�4�p ���m�� ���;�NF-��S���$JJ��-\��i���wE�MF*��!���70)�4�G�Gs�N��.�#-�ʕ[���������<Q��,��iܨ�<����CVX�̥Oq���۩l�)S�qn���
�h#��
y�oQ�[�	H8�U�Xd��cK!�Z��"�5�A^�|A÷ܗ^\�IS���[�(e7.�(�G6n3(���i�M˴�,,yF;f�̀j��A��[aA�u�&,�N�ST���E�b�i�VU�9��[��8���ou�����M'��=�������#yn�$rz�����ЩP�W���=�h�Թ!��Uk2���%هJ�����7�j;��1�N�f"�)�亴D���C��e�5T�N���੹�!�KR�(I����課�)�٦�A�������%�Q�u��K(����򦘛���W�D��Ul�V^����R�6��F&�J�Bv��u�q�^]�Z����Z���fɥ���۠uD�&�L���g	{��j��6�DY��H�޸5�QI.�֚5f�Qe�����,㐁Y��z�]ZU�0Ԡ�cJ҂k�ZX�K�����8���^�C(* �,�7��7N����eŧV+�&v/�݀J�������d�5�48�?I�g���sve9S75�.#ha:���W�����J�݀apX
�ɢ���n�x����R��$�%���Vُ`sTj�A��`�����pP;�S5�2P]�]��K#Y!6۬#^�3Y�'��"W�>��ʍ�A뼥�6���h��ub�'��'�z@�$��N��l��,��m�����H�3/N��L�ůM�@6���Ԛp��Ś������(c<�^+���D��6���9��6���m�tjĲQ�]AW��f�m��g]Cw.Ӑ�����>�n2��3��c�@�2ZU�f �2��RL�6[l䕐Hmk�Sn�tʞ��:�6n��0�璆i͠5hf�Һ���Cv�CJ� ��q��[���=�:�.Z�uBj���D����	R�tp���g��*��"��ӸF�h�,A~��R{ Ӂ�6���۠���e�k �f�[�[�y��ԥ@!g��V�öث�m �VM/\�ed���uB�i��@ޭ+y�z��B�A�1j^kpS���a�6mZu��b�����FB�2�,�d��K���"�N-d��e]n�<���6x<���4�(}�>O`�%�QG��r����e�n�	!���Y'�T�Ȳ�؍;����V���)���.��5v@����j��`v�(��Z�0�cn�iY
ff�0��	M[l��GW�գ	����E�r�Y�(��k�ȍ� 9�a�,B�22��GJ{��U�nf;��������;���f)�w7,�1�v�\�l`���DR:jmE[3)��
�(��.�,��=���*t�4��
e��ѹu#��N6���f�eMX[���6Z)�7�����j�ؚ�V⼶k!U{NXv�2��q^5H ���20��*LKL�ol�5­�vX�2�y��vژ��P
ܽ�Ի.G��]�pыUio.9qF�R=ʷ����O%��Y,�v��\U�(dZ]Jck]�y[�tnЬ���-t�o(VS�ˎ�QV�hn�����7x.��P �Tg.ۻ[b�\����@aڑm�1�5r�ܚAɒ���)��In��nM��'����	q��
��W��܏����<%�c���������X���KaV��;�+K�����A`E��n,q q˄T�W�]��B��w����m��n���MX:�Ǝ��3,��X�3��G!$�&��u��'�t����*]*��
�+�O����D0�p��AZӳ�Z��0���`l��3$UXtk�������;�A��[��ɴ(h���],���8s����5�2�F�v�0�*�ReD���eIp�ac��;�(N�8�+ ` v�j�ɰL��89�'n�2nmb
��)�N:�t��T�CS`0�u+NT'6�`�H�i�n���Pr8�pj^J�ykj����a��x��������Px��Rʛ*LI�������3����J�N1�ȡxV���tt�y��*A ��1�ks]%��A�	t�ln%�0C:����h�^�sL9��M��sU;��jebǄ?�Z���j��U���������h��G�����q���J+S�:�E�z0	&��[.�3fN���B�=ѐ��!���;�k�;4XN�h�5�5���5����CYB��M�V��;BŤ�yBd"��
R�iWp�շx�=U4"�L߯d�6���s�L�/�qZ����p�O��*�^�����yJb���}s�c�7�}7Amw^��ۯ_��7�9�+UOxXoE^��{�B�n�Y�}�)���o0�D0��%���B�>�7Yw}�,[�wzn��*z�f����}X��s�6�xjűe�}sfP�c�-Lâ�/����ދ�=L�&?Ks}ާ�{�U�G�N�.^=pK�_���^D8�۶(�b���A��6��&Nٹ��S*!]6�1���԰�-�����gU�L�t>�t�Yj�o��o�,�r�`�3�2����RV`2zDi����J�%w| ۊO;oc�I�ݠ�^ˣ��p{%�c�ovM�o_�՞���qᏦGS��lc`]���T�t�g3r��(d	ݢ;�z'�he4ر�3��^3�	��k��1��Q�=��Zt/���1p}�̿l���^-n�`Md;�0���˘t*��E��}Ge�6��:��2�=�+��������u���K:;|��E�S�SOOT�{6�L�ͦil����� x�chaӴ�N=��\�i�����<9[��*���qɲ�Pک�p!쾮3���#S��cR����f*R�Q͡��6K���=����Y�m=�+9�qؼ�X�K�IV�,2�sq,�	]�����c���!U
��W���թX���f�r�=5������p�	��h�c]�t��v�%u�	�x�6�9���5y/C@����@�W\z�7��^�0��}�M��ݐS�`�~\ƕB�\�S��%E�y�L�=](�U7E���T%9.gQ�1�f�t��cSr��/��͏�ݓ��Y�>󬃒��Jd�M��4JW�_4F�u�����b�q̈́ZC3���n�:E�:t`��ws,�B��6k5d��'YB��Szyn���fU�o�;����uR7Z%야�
M*��<���O�V@����l~r�-�N��	:a�FX��FJ��b�q���ov�ް)�r���)z�5��[x�����ˇ�X��#WFky�e�o���P�k��Z<�
/�6����*�6��ه�V�\~�ܖOu騫�4oy�9y� ��w	�&��9��Y��p 0Txac�*�ő���9k��1���h2�%�U���ﭒ�����:!��,W��i����s�N��=;.��6�Igb�R̬���v�����Gr��>y�����0v�m�<<�?N����p*���3c(�f\�L/��u����;�c'��s�q4_t԰;���9Z� gX�P� ��K��k�Y���śƎ��؃+��bk�70/X��}���Js�י�e�푼���^���/v�M���:s5��kS��[t#��D��')�d޼����_�k�\��`�t���K�Y�V4���d'+��^w�Q�q�퀑u�����n�l�	�AE-��{���\;×R�����F"Z�:��j��u�g�k���V�����b�#�}�T��C�� r��|Eօ��V+���(�G^k6jv(7l̑,���tcؔ�<�SWP$쾯&�� 3�i�%��]l�,"²UH�ΓK�o�|�+����mL%.�Qgi����n��y󋼕�eQh��l8z���y,o5c�4�R�{*Uzg��6�h==�*�쉭�@m��@�-d�p�R/��^��.�-���>'�Rէw=�L��5n-��h�=�16���Q��1'�,;.��rI�5>o�y{[�E�W��3j�:� �Sg�o�X��^ �B������m��W ���j�Uͺ��sr��3�{�f2�ݸ�CLHxW\)��f��jEI|@6F)kpU:�7��l?m� ��1�LO�]:I����GS�/N������Z�襵]³L�S}Y.Q�`6{�뻂��A	���[V4�P���z�1{\�7����{|:��e]����5Ɉ���;�>%�V�U����I
�)��-IO�QS�Yzu��fd�Ú���'yR�ϻ5\.א�w�Iy�������t�i������W,��wó����is=J+a�[D]��"&z+9�0{���ѯ�����8V��Q<���t�&$������,&�5_e]��ȦF^LD�Ok��>og&���6F\�� �p�㛡>˽�樲�̫-=p
�g��l�H6�X��f�7i�y��o��J����4{.��S�����8dj��:�',rW�ŦY[�vX0�3�܀�����;W���=jJ�uѡ���h�y[FS����	�@ ����*rJ��\)�s��/�{���葪fue�ڻ�Ʀm�>�Ubu�����6��&��4�fɂ�9����hpΠ�*����S"�Z9�Df^vr��/�:��xg�ዝ�ǵu.�L�f�􂄮�b�jԇ�"��D ���� �������Y�����)�\���D��aQ=\@r���T{-3�����"��aPXݜV�f�)�@��������}8���WS�c{�.����SOU1�cxw��ڳ���3D@���Q*Y�6V��GD$���{�a�i�o��\y2�'w���XE��/�o�n�,�׶xה���y��C@�Z��$y ��楩'��N�zԦ�N�z)rWW[WZM_0ٳr�
��ċ�[��Jኤ���@i�G})�Y��H'`{
T8ٗ����F��p�s�^��5�uh���������U���V����^�8q���O������-�n�d�}*�c(�/*��]^I"�4�)�����7mS`�ʍs�:�mע=��r�9uHwa������>ʒ���/�\�B�R�Km	�����ٲ{�<=��б�<��체��*��@-��G=9:�~�����wnH�%��+�C�A��-C¦GvN�a��t� F���k�Iq uٮ�xE���m�]��]�݇�ZTV�"ӝ�X�s��1��,��8R�]o����i�:��]u|1c�/K��"�:٬t��N��+faf���EE9����)���n�F`z#>�'no��F�M����8�wP�~Q^
�����@�;&��=g�]���s�J��	t�=�a���$X\�vO�/q>���ؤ�ݲ�Ͷ����}<D�a����wy�X7����TB³��v��;��v��(��<�ynU������Ϻ�k�y{��u}�2�(y��vόzG���nF�Ց�� �&'sk�p��G2��t<�5�ok��S��b#8+W���}E�CfL���m���l:Cl;h�	��}N<�Ǎ�huj��Ĺ��G����N�E���{t�$��N�p����)P�Ҿ=8�G�ݒz��V��fE3�!ƣ�	�uy֚x�fʵ>\�Uպ��]gQgk���J���Xuk��+!Y�u�n�pZT֚��qJt�/h�(kd\����5�Lt��{���2�rn�eԁHh�]�����rK]^�h��Va�kX�)"�����=���Z��v��t��T�F�\�8���r��
�	V�N��絅f�i���6�[�RU���I��n,%nήaȗ@����N^!�J�`��/�*���P5�53p[���㱅�����S���c��x�q�Mi��N�u��K�Gh�*Z+57Kx���߱d��,xt��kI2�p�$���G���h�[w}����F�U$���2H��2�}ĭ��W'�d�Z��N٠7�@��m
������e_����t�cw������i�ֵ~���R�>[���ru%�59��M��\��#/�Entr�q��j�O�7��Ȳ��}��Ӵ��*�GF���o>U&��a���0�`�m�Y��6����efFuC��,�j>ۺx/\{���p����4�k�;0)�B*�X[]�T�Q]�Ƌ�Zf���"e�T=J�w%���X���>sF'�l��7�&�}}ض�>�&W��+݇�Ǔ��D�'j�(nP�C
����Vo�P�R��4��XFr����i�W�ےl��ĝ�M��t,.Q}^��ҶoRe�,<���k��fZ����F(�7���R3H�ǚ�󲶲�u앒2\���w�;s�679��>Ý�ß�MLv!�y�H�=���=�y�ņ�}��d�,�E�q��t�ҧt����5�A�U�d��C_^+��N�����5wp��Vs⠤�Zo��B�*S�G6'M;�!2���+�|�ث�,Fx噹�P��ugx�ݝ��+�c��
�	+3]*NW�����7R�6!�|�ͧ��U��[�x�a�\F[/� g'z��xgd+������V%��o��7X�8sQT�wa�y�?�S�˃�=�{���kpQ�]�3]��]P���e<�+�rܱx��I�ɯ���P�Ȃ�=��=X�Wp����/V9j����%����U�x�p�Y�ehS}o���Q	w�'-�g��/z�����oyq�F�����O�'� Tf�y\�f�;���j�س��d�r�Y	x������鯱�T�W9Wp]����w������,A��X�設u�a��b��I�1>9a�{3�Z��yԺ��*�q�{(�t�܁i�Lgh4�:�@3j�Ӝ���K�bKa��7⫤�q��ݩL��gR���[F;ᖊ��������1��jt�'�]��t"��+�#x�*P�d�u�����	zd�Z���]�KjL6�:t���V�5]C�5���I��r�����-��B��d�[���凐^�D�dp|}�:�3�_h��G2Ӟ���r��=J�m�0U�溛������η{J�r�����gok��#\�SH�S"_,�֣�.lXWi�Ն�!m��-���7��(n�P���K�y4b�U��{�:�T4�P����P�ƥ;�Rq2)Т��!фR ���D@�<���K��9��T[��H�p7q-�]��
���%[����v��ʹ�;./�0�l	6i���4�p=�KI�3�ÁE�%�3�ԁm���ki�O:���"=	+:ř�3n�L�d��+VX�C�OR���l�G��L�u٤|-(�����⫫e�1�'�\f�W�)�q@��@�f��(��(Iǂ0 3��l�H�<=��ȇ#IlF��^� [����	َ�w=�WL^��~:���0`L��P�v�}w(7V�,c.�֟l����s�X"$Rx������-LHcb]��'�P�劭���uGNى��Vo��:��M�h3g��	m�Tsݫ��lM૙*Gv��ӑ�G�#\����\GM�U<���y\�ܼo������Q��b������1�ְ��}��s{��Z�s+�tve�aS�P$���K������[)G܈�(G<�cɾ[�m��YGQ�3{�]��B����aR�/������lhs��K�4�C�_ �pXգ|-��(v	g��RbI��o���9z0��)S��noD{�:�ξ=���
a���,��b����%q]��?G��{�h==u�V{�:LP�tt�_�%��S�4P��{����R��0��ĬĴ2�fXېݾ��o����S�i�G90oLTpN�mL���h�#6!��{q��N}f:(��4;>�j�B�S�Qk2a��W����u�e�Nm9���7�����{D���ˁ沷��,7�D�2�F��j��*$u�*;�{$��w9�Y���M
�]P� r�e;��3x4��)�'�]lLDFALh��<@��r:�i���󥵵{)'[�5�}��3j�KO�w��~�朶'_�W�=��w(c�ߞ^30�J\g_6���n,[�<wO*��!����&�؎�4Y���'b�8��X���)��q�#l?�K�>��cز�g[�u>W0wA�râ0��%�0�:[;i.��q�Ι3s!���eu�,��q�lAw��wt*��b�Z�@�Ϧ���;5Wx}8�����Hv`�����/�[Z*CwnɏK^��T���I�����_(d���q�嗕l�eeI��
�I���P�@���D��P/�"��u��뺙Q��Tٗ�(��k {�Ǘ�z�ُA�ދP�r)�T�n��D��q�ȹ�B5Qy�>�-��ێ
X�Z�S�nb���߶P�E�yE�vL����s�qC�p+���(�Y3��`AY����2e���6��w���)��9ov��Q���.�����\nq�Ab�b�ڵ��
z�*��e]�.B>L��j9} �b��e.�+㳵?
�p��%����r�jz��r���SGo����!�;��r���(�� B�e�9GpR��&>���A
5�Wo|X��sG9�7W��ly���`�Swʐ�<���j�^�OW6�<�^�^?9���m��V�����O�݆�p4�A���Ab9���EOԇ��7��칫�7:��[`�#��MO�X��U��1�jG�����+�ٯ�����gXh����S�.���ݱŗG[o����y�fdᴜ����o$d>�;$��\-�j-�U�����_J����Έ�K>�gc�V��P����_�r����
v\UKo��-�[o�,��$���V[l�[����������:ݲ?�K���}�jf|�W&�MIe%Y̮4l��=����q/�{N:IC���GA��������u�L_����2U��S�\k�++Ź���ܲ���˖�T}�:g9O��	T�gK5y��1� Ӛ�SOcg8su�3z��)o�e��K�N�q�邺��Y�z�w��4W��4�t�T�K9�<�|t�E���k���0_c,Dpd,kZ,ʏ:�vl��}�
+�*�#u(pcY�G����.>�$F�iךd�~m�}���CcٗE��'|��.�u���hZ���!
��mC��2����9�����SYLp�D]Wj��}\�[媳�p���'�Î�&���:��bGо��	f͍����Zsu`콅��0Z��F���-u7/�GL�J&ַj�\��Cc6吒�oL�B��y�{�f���Q���:P���x/�%��嗡����dԥ�5����M���Oa�-]ݑ�Ǌ�X��۩�x�Yi�n�����d��D���9�j��g �	"t��ʹ����[����b>5����*�{U��{g������T���i"%^�9k�%&s�R�͵)2�;��W��@�#���e��T�R�`ų�V�=9�6���|$���޹���N�2���ѻ�qs?h�>˛�fݍ;i�k�9�\���b�����yM��{������;��U�����B�Qa7lp�nAm��(���{ܴ�u�s8�~ܵ�#�<���, c�"��z伮�}y\@�UMᶁPͺ�g{)|r��s�M����Q7�����d WO�H�evPHK�&(�'gn�I;��q�ō�c�lZK�x�[��$Q﫯ۯ|�2�&3%���a�N������q�}9�9�g"f��Q�:�lSo+i�}:�r�ƀj�朼�,Dww��jQ"�oٱ
֬OO{�Z6� �:
�&^���e�׈�p�T&���å�G���:n�3c����i3��c��w�k;ξ6�E�C lyo�q[R�E��ye��72J����F�D��V;q�!�CL����t�Vt�9��#]�7�Gl�e�5.�<���	`�_Q�ӳsU�q┋��d������َ����G�zLX�7ݣ6v��D-��Ҥˏ���[�������	yO3H���^�lْ]h��g��_��o�'�*n;��<��P�+E���eT�OdaS���9uJ�t:�mC�cT{l>b��9\�����o/+zocTB7�\�j��9}�zl` ��z��U��Ρ�v�4��1X=���:���h�K��:�?���u����v�d�;GR3�]�m-�xƱfa�{b��˰Ԁ�cF �8e�Srj�4�J�4�.������Jٸ/�	˛��`���Z8��]�4�Wq�fg;��i`��^7yؙ#�ӊ��CEMc�'4�H��G��6��9S���u���f�ŘH�-��{ٸ�u'�c�y�u��}fw^>�r" ��<�ԧ��U�.�zL�y)��ݺ���A�p�؜���ϯZ?\���� ��E��Z�B��]���i��dz��|Si4��}�rV�]���Ab;ϔf��V�$zK	#
G��[W�����}��`��v97컋j�0��j'4iG���]\e��E��:.��ysWQ�)����bz^m�usƯ�_{��o���Os�x�:q�=�X����j���)a������Ɩ�����;��j/(��W�z�e�v��
^-�D�ײ�yzv�œt�s��s��
��9�eu�����_:��*_��6F)���jP
ΆX�/*+���l;����q����&�
x�0�m:�
՚]��ɇ�����6r{٤Yhm�k�7P����]�->��r���@�˗����v�ئ�t�p5[`Z]*_���f���v����fz��v��H;���ߔB��r+��X�ܮ��T
7��'��Z)�o3e�H�N3ۋ*`(CШ�^ې�h��;�oq^1�0l�b�2n��Pv0OB�p{�h���;������YPy��@���J��AΤK�&��[Z�7'#�;�����]�z��i��Os�`��'{uw����W&�q���-0W�9��xJ����./OdY�r�4L��Q��X�:gŉ.�eJ���g����8<�=����=�8����:��N�X��8:C�
�|4��d�Ղ����I�I�+��eJv_V����	��(ի\�8X���1=�vޅ1�f���*�G����֒|�`ɩ��齲�wt�n�hC������({L'��I��:�m9D^�Hy�1c����y�(���0 ���j�A���1V�k�A��.&�E��Ǝ9���ı�F5�T�<���os��/��5t(�|�1�NkJ��=3�D�V�V�'��HV`��9�B_ri|w#���lX�й�g05���X�@d�X@�r�'@�7�i��G����z��	��$8��}�{�{3nBEr���J�����xQ�,��}��}#�yIx���ۢ�'QF�s8��yOxD7o����^����]/M�&�^֋W��ڮ�7�3,u��'�$��`�=��|*	j�J��{�ޛe�8Q�i6�`L���N�g`����E�:ąT�\LJs�&^Bv�	|����`��F��K,7F�αV�ږy�Ԏy/t��C��˗ݨWa���v�`|]�"�5�Gb�,%3��9оB��J�mM��u*��f�O�\Ժm5�Z�fn�'���)�R�p��``v,�R�
�*�p��;��;j�Q��B�l>�5��샺��'
���`G��ss�آ�#1-�Lm�P�mw&oV��mB�^d�[n�GS�o&ͻ�cH��zZ�2b�b��;��g(�>}Gӽ���z�o|�a6����F哾J��z^�T���<�+����uf�ne'�e'�=���5��ݶ��6�8y�z���T��%q�l���c�60'�=3���.�K���^l����#
��Uܶ���!*��)�0a�B1��f���ѩL4sJ�v16XǬS�8��@v5�yΐ�Kj�I��Pa�\<���k����ӧ�,=�8q��g^���f0v�*� @\^�q���-�d�{�/>'S�5Ot�Ş~��Ksv���X�+I�VY^�Cx�����V��n]V�J����s��3����b���"��u�FM���{<�oDp��Z�&�}�i�_e"�\ݕn=9��F#a���Y��6F:Tij+m��U]�|����T�E'�1�=�w�ښfuh	��U��U�6�4g)�k8l��S�Plow}��9�[�7�'k᫞���Y�c�jwX�|��Z/M�N� *VK��NIܘ�#�ޏ�0/l���*;g�è�F[%����t`���tH�Oq��8�箛^��
��-��48U���h�|�	�]͝�(>�Ls��pt�I��湊?ѰTx���wO.���X���0��hj��,�����#Yt-����ù�����T��Z�\O��%d�A��`���pn`{od�4c�ӟI�i�wP#�9Hk����Z6��B�'�%���)�˵�}�q:�"gm��Bvw���Q9��'�{��K|8:SD+P���ρ�݃�a��gC�L�KU�n],�����_<�^%´��s(�WY����E�Jm��I�(]Pr��0�_Z�d����6;cM�ޗB�;�/5J��$l�yOd�vZ�P�	��b{d���䆽l�̳�d�)9�y���z#}ʇ	VNܬ*�Y*nkƘ�Y�c#*�Z��ͤr��6qu�5�֛�2�u����]V��&��|���y��'o�H�zu P�N�����p���|�A���H���{��z1�d�w����W!Yݼ"=�xBL6ȨN���8��H��w���M�׽z����81�[f���CsI���C�pǞܹ�v� b;P�w���N��a�v�\��ʉ۸^SzvX��W�����,� ��RZ�s	(�h2��Զ����E������Ut8�+���2T{@m�]����D�ں0��q#�M��
H�����l�T�ǂ�7_N\�nxmq�r�x!�ɍ�On��;�ʜbC<Ca� �8ȼ5{�����s��*7<��in�YGi�k�Gu��)r�tb�W��{�O��U�Y=؁�j�魵[U�����r����_ D���݉9��[xe+�|=�ά�����7�F�˭S��(�ٓ���S'q�&u v����XΝ�c����*#N��k��B�&��{�}��E�)W�* ^țoۣ;b��a�w�BX�]>J%4-CI�-9�*3eZ��D�]���7����1����Y`͈*Ʌ
eZ��i�\((E��ا8*�gV�b�yot�ozoќL˞�2�/Gv���S�����M��O�;Z��yn=j�']�#�ɞ����g�� $()w�2JktfmUxXok�:I�E��뮣�a[53�rU֓w����	`�'vJ�Ht�,�^k������k�+H�"��2�*�gK��F��&^���Q�e
��i̸U�w�'o&zɬ��8
�rc��]�}�p^��M�Z;:Ebv9tn���k�B���A+n"�%���..�g`w��P��mЧ�Ν�Ͱ�ƭ15i���,O��Z|DS]r�ė6�,RTOx%�V���,�l��؉f����Y<�����G*��m�c��/�8[��Y�a��]]�hjQ��T�o	�'k�0���O=�{b]��=䇵�\�U<w[Â�'M�~ZҸF)�.���s�	nn��!��4�o�2��}�aI^#�>���BX���뚕y�upʣ�׽B�����~�v����^5���°���unŗ�\|�wt8Ağ�-�t���x�y�!�1;�F�fc����2��g-�5]�ca,�yC�VMr��'�iZX�PӜmkh-b6��1Bˢ��ќh���ٲY�Unz����}�u����A�����%��Ηs6���<f�+�:[�:��x�v!��Z�RR�[�h���S��<F��5_u$Dd>����6G�nzH�c�`N��s���&���ɐ0Of�;�y����}�c��ڦ2�nr������9�<�9X��Z6Z[�Μw�j,(�54a5�
f4k4tJ�"n]�꾖Q}W+D��L���ec*��yw�i]��Šј���==�og@72&DL[#����寃Z��7a].م_]X����s��GY�ɏ�X�Aj����ɜ)E��C�Ի��m�{�lYR�O������*��*���C�}��_��q,�žWQ���l�{�f�[����T���y�6��Yd�Ҙ����n�w�I�{������彠�1O��Nx�k-VF&�V��L^M5g�$8�wL
�6�֟�r�kzHz��e;��!�Qx����t�ܬ����f�k��<ݲ��y��)���i"��v��*��j��Ո|'B�:���eÔ{2��"��z9��i�h�5�]:}f��Ґb�ݚ5�G�Z��q�S�ihߧ
�^{�X��Id�u�esw2�iry����o���HSȕ��!���G���X�J�t�0��cTb��LV���+o#���S3n��΅�F�o��MjN]�ŝG?x8>��ϩ�G`��U3���}B��R��.�/�i�i��r�_wS�d�X��˔&���{�hR�t,e��᥃�c1�����ᑜ9%RKh��S^�ȣ�Co,i�-ZƩ��>Aܫ$�gW�o�f��0�Lo�p��[#���iV `+�Vu�k(����a�@y$6��	�������Թ���rׇ׽J��9j��O<�E�azQh��B�=J�e�x�N�,�%��,"L��k���.�����r��X[�P�v����p:.�3{[����uų��+ �ne����S0@��;���Hõw��x���L��G����U�HWg��`����g'�v�	�{�����3�.���a,�.��;{Z�;��D���)�
S�hM/Kү]ǉ퓦�p`I��������U�YM�:�r�º��z���luC��z.��l��6ý��+�jNݫ��ݝq�����_s�\�j�)���JѶ�;�+�Yx�T�Z!wQ+��-�w���7�p�8*gF���N�Xx1��L�ª �Һ�V�j�RݡŎ �k�kl��fu9��
hu]���1`}�q).�n�m;�=s��M垏�nv՞�oO�*���:o�hd��L�R,�ǽ|��_Bt�\�<��s���a�.�vva}�z̫��S��o�	�b��+a6F�2���iu-vs#�Zi\�н�ؖ�Bk�§Wu��;��&��g(1����4.܋si�D�9r`Ƶ�u�&-Ԭ��vGxlQ����DSS,Hd�9���ةtD��Vj(�ɜi�����C��b���$t���������!�X� �Hl���ܹVv��jTk�]�ć79�����ks�G�"-��N��z緷]��~��� �Xft�GZMd}Nb���+��}m�_!�hs�.k}�T:b�b�
#��!n(��W&m]<{��+�$�&�ޚ���zl��x�+@���Y�+ag�����v�t�ia)�t�A9��	yԦ��Ρ����!G2!���\��'��E�ſ(�؍ (��R�1������=�{�x{�@	뱺�R�l��A�3�f�
�Vt� �,m+�xf��+���~5��6y]J�nV���՚�{�-�v�񣨑�8�#�8k�;�0��=��#�!6[;�l� �6x�T�{`���
5P���;�25���&��q
�ٟ��m�<��m]��� ����A.�����$�]S���s�ǻ�_	%�fJ�O<��-�$��罳h�����r���x��_���X�����O���.֮rv�a"��,1`�
�^�����r�a���ʞ�u�lT�AJM�v�잷����R�- �����&��qS�̷dQ�sF9̍�Τ�������<�����/]��A�zu �lG ���½��B�KN�0�y�D�&�����9��QFhjs�=^����`C���\��>{���C
�w�Ȇs���P�z��7w2fs��,�8ܧ����p�8^���R��R�$��.�:���x�U��f���ޑ���v���pQ;=}�gg�����k�IB�!ԝu7RVo�ls�e�V����pP]c9��!.H���E6���E���7Q7i�|�f���z����R���Iv�ۼ�{a�,�c���4ST�p��n��Ė��f���`okn�{� �yl�E�Dq��]��}�b�1�{Ǿ��p����=ۈc[�������P�|]H��	�đUZQ"h!D	
* �� Sl��4J�B$�l�&�h ��"�"�Qb�6�T"BU�@�D��������jmI�@�$*�*D�H���ՙ�4�,*�B!
H�UDDB,B$�����UUD�!�X��u�t$����bA��"�!j) \��v��f�Mv��R	6����m�X$�DM@U��!
�)"6�ai"��U)�2̥D"(P���M����h�H�%BD
�ivԈ��M����!�H�$PB�B��]Qb%$�Q �"��@�@$�p�PHB��H�Q����O���w�>���?a��7��,���%�,"�a8/��x����y>~��+���Ǥ_
nP���&	���ݽ�w�}x4܆��Mp���{�B�E�]��O7�T�փ�x��V_7���9�;�� �8w�=�	C���']�atV��h=y�{����N�4���ޗ�J��Ťt�m߰���l�&�iX��3�4Z��(�.S��N�x��<�^U�$��<����w��d="�LWGjt!;����6kJ$e9����4��K7�ם^�6>{��Ǿ����ꕇ%Σ����{�D^嵇�$ '<r-�����)�X����ٍy���p7�x�};��|��{O�Ƀ�=�{�O���h��}�4�q�,��Q_@���\��-/�����YH��S�Oo�Ӂ���:�x�n0�u�����r4.E��$o�������CP!m�J����0�l:�:��0k|cq��$E�Z��d�u8M-<	8�K�UC��K�x-48Қ6�u�2�S��2u{��%��M�ð��`��ײ� ��������3,�`c={Y^}5"��F��o��u}�Pi
�J�=i�u�X�v�E�˫A�4�\�b�-�1�p�$g��Vf��+f�L�t�y(Cg3���Ox����l�Dw�bN޺��;�v���e���g�=�=��J��0��x��k�^�vܭx�|�UgN}0�ظ`s�iI��q����\+�h�{D�׾[�0h����?z�� +�#�uv�fX)�y��t�W��eF�;��t'H(��s\��Y�J���Hс_���D�[��<GC��b�VdW&�F.�"�#!�.���X�Y�d�?�S�k�3�]��Y�Q�:���h��[N���R=y���Z2/BT��L�8]����[l�����x� h��|�z���#�_�W��=�Ô�o�3�{���o��
u:	�Cn�λڞ����1B��&M��Ds�t��L��WL��LxA�퟼�t��8(D�='���'��+��S�r�wh��>dз(A�	�پ/�"#�.B�uU��U;��	RbNՍ����?
�ZH��.�f�!���59�#�ώ�d�붬��Kf�^<���o4S':���GX�M,���Q^���FY�g<�s"��j7O.$N���'eߨ����BMZN`5��s��V/�x��� U7���q7N�^`7��Z���/;Jẘ$9)��l��T6�ExtX���P��c�G6\�˥~�S��_,��Cʞ8%xA�b�	\9��/![�i�>0���,2;k9�)w�A�t{�-1 �gL����t���Z�z�2>]fh�u��|n��+��ռM��-J��˖U�/�mt^t�B�'�	Vp���s(����)��o���$�G0�%�s���[�8�󞁛n�D�ٹ9�$a=���^�^'�y��o.ߵ���y�/$wt�^�N��xm�l�n��+q�GK�� �+��5`����\d���RY&�(`L�=9}�Y��ED׵;q�aʋdGa�a��@��x�r�FCT����\=�&�	8̸�ɋ;!񶮁v�許.\d_<��|M��\t.�2��Cӻ-1�$�R������NL�"AJ��$s+2{����W-ؖ}�}����eq���.yz#=n=P�~nA���J$�舄|���`����w�(6�A��KzG7�=�r�]*���Ù��9��6w�� I�ak��&�4;�E=���"@�uپ՘��y�e���S����/�g/5��&("#L9؍��-�D:%�A���9�=Q�D�����^��L;�EI�vd�N@�p�`��fI�(�=u��Gw,g��4��Ģ��S%���n-L���r�J�C����&��6X�[#���;��uh+��M�4�|=��GyD!�0�Ց�zʫv�׋���i��ER�����o�޵��j����Ы�����c��Y����٧(�묳&������"�:�dX�T������7����x_f{î���k�6��1L�Y
@�s��n�0�����ǩ@}���b�W.,s�p,bu�:�kNWt�֗���� `�ﯕ0����U����#`��V+)�$��q�������h�0n���J�\H� z{~�Ύ�~��]j�6i��(�V9ZL`�F�����o���Y��.lױ��e�01�6��a��7�ddP� ��*�>���ȭ�t���mOoW;{�ě�͖6eD+�A��r�ppS��`���n�cM��P�T�r�q,%��>(�|7�@�<%4�Q� ��4��Y�ע*�t�Xn[=��t5��elok���rnvG�`�G��+����TV���1�>�Z�A[^��B��!�=�)�܌k�u��UuGc�\�k�$�3�a�
�l�ER���}E�xp�1<,��V>�Q7���{̍�>��hd���']V��T�>�!���H��W�#v��'�@Buc��B���2$�wbWT
B4������.�N� ���`&�7�s��""�t��`{D�(;���Xt�sؕk���a�y۸w�8�N��pu*�����=g���Ј�\Z��#t�v�-R��qZ�|��ya�����׻�L�t��,��o ���&�l!�i����x�c,9�f��x�1~���Q%B�&[�Z���s��5���q�}]S��`�ґ��F@��	����
d�^
��i��5������-�H!u�=T�]xe�^���9��Q�Z��A�D��5�#ʓ��5��1%Kyvp�6�t���d�z�U}Ga�G"�]���|=3���}A�L��ˈ缱D�n�HM�o���[p.!�mQ�v��1�a܌����:C���
�یmU��艴$m��������F�nz#K&�:>�,�� 97b�n���Ţ�)ѸD����GiR����ϟ]����<��>�����֕Ϩ�
Ќ\6_sQ�Z�����d_#~���Ҙ���f��n�jd=!�'Y���s��h5���j�Q�o5��R�Rp���:�v1Ժ>�.8���q�ʠ����qW��i���o�{Y�G��}�ѧ�p5����'f|טa
"}|�31�V��.]6w)W�K}��&��b��eW�\٪�i��3��{%��U	�De7}9�F��J�����������:)�+�ޫ���NW�/�1��]N�,����S���NO\d�9[D]�]��y���B�Ⴭe̘݊jwX)�ًb\� �N�h��t�.>�x��E}'s�ി�s�ƶ>uq!�9gr�{*^���b�o�2f��R磆ڷ��йU�:h	<�U�H|j6���T�=蜭��cj덽�G�%W��~5��i��0�Zxq��!�uȞ!��PS)N�7ֺ����_��TJ�OOs�9��
5�PQ��(EA�u�@�D���@�&���سG��zWb�}x����^� �z2,z�#�jN����(9
��(�ik��d_I��Ž�T@��(^5�Htqor���z28Kj�p�e��u�M����r��ȩ�u�I=L*�|I��g�����D�O:�7]#��B��ƫ2+ܚ�.���������;�պ�=���{�Lba�ӭ���X�����>H��12�����_*��h�ɳηy��v�3O54��
�D�`'��f�DtX���o�N�W�Gx���G��s�|q��0�'��G�^�C�C����+/޵<ɒۘ�huQC��L�vh��
�<�=�u��iИؒ�f7�F������7���HgD��(��v�ycd�I�|v��o���]b�|$[q�U<{�//R��o/Lصv�c;yJ׈v5��t6�u��û��8)���C�r��O~�|��@oT�ƪ8U��8\�\>�	o���l�����wh�\��B��Xf�ő/�a��Ըz�B�o��w	5�W6<9+�i"�eC����Ο`���"�����ȸ��j ���r��kh���E��'v�������rv҈��tX�:��u̎���ć<��K�)�<�m�����W�4��V��(��,��ΔUa�K�Nؓ
"'��Y��6��V��ʶ7W���,��65]��豝9$P�������@���T��H�-���C��/*��iz�^�؎~'�&��e�����g�Z*�yօ1DlJ��4���A,���)�+��w)��V9�,ÆҐ�Kj	��.��q�-�� )��]
,d�A�o`����j�(�Ş����8��Z	ž96����
�;����(���6�>��}4v�f�W���������R4�<V���C9#��J�~v���.2/�SD>&�Fzⷘ�'23��j"����e�:�
��Q�A��BS��eZ�*�B�����hG���%�rL�:�S����W�������6�&����{I�����9��48ĥ.��4��b+��[mUj����7V��ª=�I�Yd��'���I�7�>y��ٮ��u���O���
<��e����F�3e���iٽ��ßqJ�$������Ҏ&��2�R�D�88�B>q�*�#J��D�8��	�X�ż[��}&������g 6q��A�۾��9 �I\l��@� �����N�)�Bn���3o���!�fƞ$e}n���Ź�d��5��6���"4�3#��4(u�2sR�OU������w��Y�1F���7�N�=$5Ό���w
�
eْEa��U�^w$��Yw�N���Y�E�N:zo ;
7UW�hI��_�3
S��^ �e�W`�	:����|��ٺ=��\z�c@�^']U�f�/+�)��^ۯ�g�-��7��SƸ����} ��x�ff��ʄgEAl�
vx���9��;~�Ub�n�<Q]"����H���,�[p	+	c�yq�W@��|�:b����*���X�N�¨��_�=�V)p����˞'�
d	��VyT�e����z�W�?{��n��x
�3�zҒ^S��P����9�Gb�v���̨�`i��P�)� �M��k�Ͱ��"��<�7j+ҵ/.�a�1���,���f{�AѦp����+I�����"��@&P��E��c��)}Ac4�o�9Y�7�K������. c�;��v��4�"�{|��zc���^�ϝ��WK��z�M]۵o�4�VQ�����/�䮍�m�(e�g�p<�X��Z#�gip���c�]a��>�DP�(��e:�kwE�5���7����&���a,��P"��F@3Ԣ4�Le���Z�A[c���u��^��m�cF��~���t>�2E�Wt���W;(�88�J��B��i"�֮�dK��פ�)��2���ɪ�Ʃ�FO����>�kC%ss�N�� ��H�r�
cq�*�]���j�/9gTj�EY~W��\ˎ�e�q�p7&מ;���gܐ"�m�]R�#�7;۲����yé=]���{�@�Q�hb�����m���ґ�226�N۪fb��(�^�]���d;��ö��63���!#���΃��R��|}�ϭZ�˃�V�Lc�CP�=�5]�Z2仉���Oa�;L�\En�(z�L8P���ҦKɃ�ި����^��WV�`�w ��ȫWy���傇a�����x­y^���5�[��3릧R9:�5<7�i�䪢�q�A9q^[W�p�ڼN�~�.��6S��1��>�ϩ�/��A�a��nm�A�ϫӜ�Q׼�W� ���胱��˓�1m�wy@$�?�-��]{E���b�B2��}��Q=_��En��wr[�7�'x�h�Vf{ ���KfU�����D%�;��I����aPK��V�v2:?_,��wnS{#Z=\�%]"��\��4���:�roG���.��Ҳg,�tH7*8a�µ����������N��ヺS=����zCLN�˝�*��f���f��2��L�/]*8��w;}SM+~�d��`�`�����7��x:�a��%Σ��Fo��( 
���x��Ͻ�������z��l���v���)�`xJ�\����+N�%�gDl��1l^^;�Ω����j���^,�3ngNŖOu�� 0WO����s��!�T=Č�bu�#Y��{�4.�z�uۥ�K��n}���$�#<z���F���@�:���'{��tw�o�4�'h'�SӃO�<��l����`���D����L���>���"5%Xξ	vmeP�F��Z��89�2��lA�XQd�(EA��"<t���c����Os�_tC�x͈R����qۯM�FE��]�Z'�q�e9
.i�]nJ���V%f�8�a���3YI����v�
]tld����\n7]�Ǉ�S��W�C��{�S�s& ��2U�z�m�$�5�(������"�3����s�o[�{��`(_YMj�Xm��a����{R p��d���5�b7u�#�37xb����wZD��'����f��ּ��LjzǨV8�����E:޽��,�y���g�A`�v��>m��6tf�ק*�ձG��n�o��ќ���i2k�
ۺ6(�
^����HEpFw-V	X�z^VOv�7�'�D���F��娭Aݥ��y�&��6�?�PB�w�c�Z�L%���
m!���}��sэ̄kS/{�j;�P�y̤=ԑ��'f�����̭>�(�nltm;������U�v�a;��N�i�[�C{Ƿ�\9*��6���<�nj��d��(bs�Oϫ�����ᛏӪS]:��cs׸��%��#�;�Y��W�[M>p*����p�^�٭��4O���/`A^ |�{�#����(;������f�R���pa9E���_�F�r��Ţ5k��f٣�֍|��p��b�B��=���Ƞ��]$%^��m�f���vT��/��#dо�����d9l����I�}�'3s�q�1u�+fS0J.�A%s�=�O�>±#V�e��c:rCp֌tW-����H�|l��n.�`q��GL��-�<��ru*C��
 �_��r��78��~�#�|�t���]��8j��s�� ��.�ߩdrt���z�/���yZ��(<��ܾ7w�ihA&F�o��Y�C��&Å��v���<�E��!עZ�]$��e����b\6��z�����ʗ��&:x�P����=g@���(��r��d���`�=޷��8�-'��Gc��Xu�z��h>C&�9���|��q(�;���x�m����8�|z�8w�/{�nh�����ae���ȁ���U�h���0�)vd�Z�B��J�|���
Q��#�U�r��a��s�މ�D{��y�����M#��m���1����Ԭwh�ۂ�k'���XU{|�b
���c��r�(
�|w%~�Jso*�}�*�R�"��|3D�{u;0�Xie:����u�yl��+u�c��cy�YV�R�D��y�s��|dfl��s�8����ć��L�ݭ�A�7B(��#*���[j�%QυhG�sy/z��f��e�8vL(q��lEj��P��a�ҕص��w;x�J�I�N�]h�
/�2�4QaϺ=�u�E������0�$dz���o�3�s�4���hR^H�k�C6���N����t�ћϪ�[ɗ_6([��u��·(|7���Yf���@:������Nͽ7h}v����G(�1Ɯ��]@<yu������$X��B�rU�;�Q��if�x{��u�2LP���k�h�	F��/Q�7�e�2�i�
oܟK�kx����&\�����f�R"���!TFb�D�*  �������aC.A*D� \�(,ؚ) !�Ћ��)B�mH��k�Vi"�Qcji�QH!@�4"��+#eɤAH��B�B��[]v���$mt��)U�����m2@�2TTXXTZei�*��"P�X"�
!!
T�$H��I�4F��B�Ii�$6�)K"ESi��Cm"�		��R.�B��4�(A+.�HH�Y��%m2d�Q������m��XH�`"�*6�H�)""$ʐ�(�R"! ZH�B)"�P � ��L��ݛyЦ11�^ڊD]T5�<lBًڦB�I�Stu��D�ćC����� ve����z���E��9s�k��~��s�ݽ,�N��t�'��y��d�'�I���}x��i���'î���^�q'��r^���{����v�?��o��ϝ�rI��;����o����".�&=�[�0,����"��h�B��H���9I�g�Ny�K:_�k����z�����k������ӂ�K�N;�V��,��^r}Y�z���_��ܓ��<Y�����~�����\��;�<����䣊��""�}4�����=N��ow�y�v���k�_��9�_Re�w�<�$���2e�O4���K�N/I;���$��:�x�%�=N/|��΅��<O��O份�s�雭�2��л�c�>���"v����<哥����~~�ޯ����mTE���AD_�����"��H�7�}N�e�?=M�%�/i2�ˎ��N%��q,y���:L���'��gK�"+�ۓ*_���Г����d{�%���^���^#���R�_��}I�k���Z_�qgs�:���,/�?��ާş$�XO��դ$�8����yo^kK����N��{N,�g����[δ��$B�m@�/�;q�VU�����!�Ӵ�%��z��ӡ���w94�o���'_��$��o�O�~�Β��=[�}뾦��̾��?{�v����a���V���8�����;B^~Ӿu��n���:ߎ��"�����#��2<:N��N$��/�ŜO��Iİ/�=�q���'ǚ|���S����;������-���'���ęr��}����=� `c��{�#�@��5SW�����V����V�. ��t���~������V~Yز���i�. �8G�@��&=0@�L���_/�OWĝ��{�i�'I�d�޺�y��'��y�I<L�,��jR.�J�^7<�4�r��-����I�{?w�z<���K���yrX�ߖ�Jn|�ި t /��tz��=�4����/����_W�%��o��d�|K���'4�~�ia/�ޞ�k;x���!�T:�}�\F�������@I�~IǼ�N�֗/���{Լz��Ž������/���|Kz�~��rO�2X�����Iؿ��|�S�����n������8'S��%��=�����K����Ϟ�b��[[�G�e\���w}t��~�P	�I�<����;r�!S��(��Ms�VC2�M"�q��:e�=U��M��C6���b;���i�A�����o��`����^ �r��᳅�0S�b��z�F��`�9j��y]��76��B���@�#�ǜxT	��(i�Xu�O�z�^8��Ͼ�oia/�>�z���n�|�˓՜OR�'=��N���g����OR|K	?/�j|Y�ǀ�g��&�z`G��3�4Xoj\gY�Ev�s���T� �ވ����O�2e�>��o�~um��{��r ������׼� /\�D��=���{������:�������㻞��hq�|>������G�$�:�K�4�I��ԝ��zI<L�(�2(��� 0.z@
=�c��r$�,sz����O���$����|��W.�#�s��D[?|��#�p�~�Ǆ�5K���F��`zc�&����x����;�i;_���>M���,�ĜK��BHBOS����X�Z\�No%��o�>Ns�����y��o9{K(����X�2�YA֍_Zf��;~���<����m�_�r�9�i�x�����4�/��o����gIx�?��u��~if^�Ĝ淏�����\�m/�)��z�%��<�I��[�����N��G�D1h�joL�<���>V�RA�~�%��;Y��}��Rq'ia'�{�zx�Ĝ[�5��&Jx�-��ԓ�v��w4�}������L�=YϚY��?��N���s�/�|�ӵ�$�<q~sN>�>#�8ꮚ2�Y����DH�řd��9�_��8��]�}��,�/�=^$�>��Rq8��'s������'O��y�_�2_Rd�=�N�����q�_9�;I>�Y���v�o�&��r}��#�qzt��/����nsD�׷$��>�=�_S��[�N����[�r��;��,�'?k~���ܷ��/���|��;�K2���~�Y���K�����S��:IĞ{��HBO����9{O�a�� ��	��3Swӏ{��?�(K�Kx�O|�N/����gvm�����Rw��_�8�;�ާ彋��/���,�;OV�q~'�>�̗ę�o�;��,%�&}�y�V�O��fW���mo����^~����I��o�1���>��_ ����:_�,;�Y��'k���'t�/�ŜO�;��:K�~Y��>����a;�OR��Y���>N�rμ�d���g��ܟOS/ջ����Ž%�&^�ŭ�?�ת�a?����Xt���n��o���8������̳p�md��l3�Pe���u,	�#�6�$��xW-��6�&v��m���G�40M$=s�U�u�EN�F�as�$�����>͆y��+z����Q�E.���S��{�C����ｖB_�y�:L��i~����L�䓏�;�{�:X^�����|N�t�;��N%�8�I����>if_�=^&O�>�Ia|~�_��}_qo��\�"<6 0=��a����-;�?mZ�1J]�=���w�J=��xi��N'��x���t�5�S���:��N��7��|�'���%�~��u�r�Y��:K�M�o���s�N%�~8��i般1��M�?���c�gxvѥ�����qd���:_�>�q�N'���$�HI����$�,{��<ﮯk�Լz��Ͻ�K��o?i��}�$����/�r���$�I��4����-��䑈�>���nI��2�9���V��|��Οz��~%�&~XN'��������ӟ�Y�;�ս�o���O���K���m/���R��	'�w��I��n�y��/���'�����N%��O���` L?duP9W5�'V�kS���w���\�Βq}�Z���O��8�x�{XM�~��_Rg���o^����_v�o�y���y�Rv������z�aar��缰��k<Y��f>�1D��m���k�rɝų�}�w��֖e�'��$���8���~I���K�N,�~k8,�2_���,y��':����oi'����N�t����g����d�~��w���/ę,~8[��b<>���}<'z������j3����o������t��7�o�{��,����'Zω:���>M���g�qo�����Ŝx����X���?$�X�Y��8�/����>y��G����O���`M״_�{��ƻ=.>�'I`M��[ך_�8���Nm<[��{��N�N&O�q�{�������>��4��b�K�q�㵼N~�N�n�-�[��t����_�'�)}[�V���W�u��^p�Y�����8���~��2�O�8�w�%�;K�y:�ެ��'�I7�p_R���9６s�L��Og���oē����/�N��żK�w�/Kw6Y�k	8�o�@̰�����9LMO_�`�Jܗ�֟�XX\���s����qg�0y��/���I�ϼ���Y��O'^{���Ԟ���������|_q?��N���2���ԝ����S��Nӳ}""(A\E�A5��4�jg6&���=U�\���y�C�/Kf�l��(�=����u+���rH�7���D�����@U�-�t���OZ��뫤��w-Cm6=��ܤ��F�#�p�����9���=�.�\ӓ#�Kѡ>˧�#����Y*b��޴�t���:�%�x�#'�ccޘ��={I�X<���^$�'{�[�:^����r�������w�������~s��^!/����;K�M�d���=K���/�şۜ�/���8���g_��yk*��-n���~��@����z���־�����/R}�^�������6�~��$�Xwo\���{��'���y�������$�2z�߾����nK�L{����!'��w߳��q!)�_Vj#޷"0X��(�����C�����;�2X_�i��I�/�'S���|擋�'skδ�/��g>Y�OR�'ia{�y��gi�'ԜY���Yо�ϫ;O�~�|Ki2S��.�t���f����>�DDp�>|�[��{[Ŀ'�=�L�n�d��}�I}I�-���y�Y�'k�nI�m'��$��K�q8��O������N���z���'I����O��ߞs�5R�3�s��ߥ��}����ǲ=���
���{�� 
���pO����$�|����fO]-���r��d�k��'��/i2_�7��ޓ�����$�&�.N�7Ž%�&����I�N}�ev�<������ � ���B�}�7�,��\�%���/��}���_x�C��1�@ }��UT�lǡ�����M5X�1�(�#�/q^�~>w�|�+}�o�mN�#�@���b�(�M�J��ư8�:�a�,�;�7W������;�}'�j���"���z��<(	.���W��n'e@xA\�\��W*�OI�W"-Ҿp��F�V�t�������.-�	���ݱ\G� ��w�O2����o�
Wso#�2����e=�Yܷ*y�V���o�o�>��8]#�,�^��&i�<>�K^��v�<�s�*q�o��)wG	�:n�2[���L���3@ŋ`���B�����EGO.!Ы8�L�9���v<u.�����h{�,��F�'i����:�Yq������Gޝ�7���D|���i�vb���X?�������w��h�G��������8y~l6E�T���t$O��L�����pc��uw��;96�L��]"�"��u*z{��|F�Q�u�	�P���ޤ�����A쾥*c��1{��C��|����n�h�FE��i�è�>���"6�fF����!F��T�41	ј�I���Nw�N��-uѱ�[W�{.5Ej�y�y�+U�v�M��%����b%HDB3�0!*�N�&y�QZkG�hs���DA�K�!:�::MsWZ�AVL��z�"�#!A�[~x�K�GƵ��qg	v?3)��;�{�ԫ���]�3^By����"�HR[n���8��"2"B�Rf�J'� �g~>Ov��n�?YoTu=�f����R����<9>�X���-O2d�m���í4�+q��ɹ�]P���7�z�f���K��{n/HXqU���U�1�|ɫr�N��,fH�z��0Mgfp����V�}�@r�v�
�x��O)�FaP�٨�q�^���8T�d
����_,E`˫����,�ӣ���,k����%�}�C�}ɪ�Rѳ�|�M�6�#�u�M�1�r��њJ�C%�d�;�#I͏Ԧ^��a���R��r�
|;��"�A�IE����	�\M�!,҂2�賲Vr�ɑ�c]���9�{� -}1�������~��Y��@� n��VH�{��*�+Fz���mz�v6~���e���E�Ѿ2�uȋ�5� ����BJ���B���>���Ea�K�N�r)W����r�{ٔa�R&�*vͤ��Xmtg�4Qd�e�ea��l_7d��m���6�R.���ߎ��Ĳɯs�e��w��@���t)�#bND��c�1�iz{w'��%���OG:��"�A"��ו��Ӄ~.!��ۖ��Mߺ��%ug��{��w[}��-� �E�|�|C�xe%�|nnQF¹Z�����:Q��Gs���U�Z^��&z�fW_��??�
��'j� �*Ln��0R�x(%R��N3rť/:�0�M��i�8vʎ����A_�\�j<I��IJ��$s+0B�t,;���:���ڝ�[s�(����7O��t��zA��T�Q%+� ?x|��<��z6����/z���w#i��8��ƽ��Ey���y��A�w��*d���JG]�W��H;R�d����1/>���u�5�gV��*�W$>��#�Q뷾U�l�d��/xYwy�ix�� 
J�qǈ�R�r�h)q�h��ƹV�g 9T�/�����l����w�`��[�!~�lXyX�{d���33>����%1G�G�;���;�:[7��ϩ���t8��q��؊
m�.���H��o��8�>��W�k��(���{H��+M�u0�9�"��vd�@��p���GD�rs�4v�c�,���{�Y
%�'_�����4�v��).�0Pw��n����Nޅ���<��Y��{2�o�0ȈĻ� N��Vz��O<�Y]�c���U�:��U8}n�f�;0�6���H�ɩ�`k�p1�����g��Lki
�Y�m�0o����]e4c;��9�4S9Z�u37�(�\R,nڷ ��J���4,���U�8EU��Xʃ��[�v��a����3���D��2��<
��,��\�{��׻\�J�E(��yz��p:��k�W+��N��ʌ����g�]C��lʈW���\�2���g�x�P�,�X�v�p������$+���j�h��W�`�<#K,�8����DU��@P�\u�b�6�j��M����Sй��"�eJ7�"#d�3 �R����2���삵��DM����7r`�w�*0���.�ۜ�vF:��U����Խ���YN�OmɪfZ��:(��%���;��k�I�9�x0�r"��^�
�:��RP�Ї�X�F9R}1T������eQO��X�����Y]6�Ҷu;�Dto)w�{���^�ns�w.g�9_�h����	������Q%P3�a�
�l�C��������i<����njR�����y�Þ�0��{F�{�1�g�`�=Z��G�A���-���]]�g^pP8l�㫍⩪�ˎ�~.C�Ӏ7&�x�c�gT�mnx��6���z�6�3�K̅��C�xU�Q�qt�o	N�#	�)ddSn���u�i�8��=�mrF��P�L:���&&O>��ʃ��R�����s�p�����_
�rn]��JI��D�f�&���N��G%�}>���:�pyi�oR�z��8��.3so��n�a^Lϵd�R��5:02"S�`O��v� �-7�:bBk���
V�MO����C�$l���m��7�."Pˈ����X�Y�-^'X?v�����:7oo����X]9h�t%#b���:�'w��;�#a�����֕��Zv��o�TvQT`��h��c�e�k�Φ�FOK�t���m:�$<!��+�\��.�%tF�o���]}�p�{p\#� �K�)b�o���Ƶ�-�n㲺���ؼ���H��1�����p�\a��y�\˅w��v9;_=C|��c�Y)kB�z\���ݣ=L����b���_p���^�&�{kv5�����xwv�v��3�3Č�C� FNC�S�}^�����^�k�uJÀY�v._lo��eNJ��g�2�V����ma�@ItUpB��������5�*�ӼP�S�B�}^����������U[��0}�ˊ���,���ĝ���㕪��T���Y����椿�Ux0>�{��Y���n���nF�ȸ����/����R�<������,�v,B�t�]�Y��ӱ�מ�l���N;'+c�Pj�b����B�����O9�8lP�u��Ƽ'��P�Â
�z{�3�.6���aDE"�ތ�v��B�d�u��2AG�� x/��ռf�)X�U��7^4g�"�봎������&��{_xw:�#��yX����� eW�vž���og����w����F/�^o�$�gr�%��<lD���Fx���D�"D�u�:�*�o�3��-��M�-Q�}@��-T��t���D׃n�"�x�Mx����$h옑+i�����a���x�i�9�5z�3(
��7�[��^��Ҵ.�.-޽�j�MQ�Nڡ7=|��[�T�n���z�\�Őyy��C*R�-��:+���9�}Q�ܲ;k�o�*�{���}���;xf��1��q�S:�W�U�{��`�o1%���nүtb�"�	Pri�]癧
�)�&{�(�H�	�ۊ��wvGJX�)�Gk/��v)���v���|o�����b�O2d�n�9��EqI����zUf�i.�[v���ʁ^�
�Oa�	Ƕ��d-5�W�$���|ɯ[� �]�hD�+�ۑ����ej�-��p�"#�E�]b$d*�E\�I��P�f�!��������Hߎs�3���Х��o�my�f�ܖ����Ͻ��+�U�6��	˷&�S�<覎YB��q�u����a�k��e]L]��wl���o��fr�6lAyI5�	ӯ��O�I�/��$$O;f�J�T�v=�Z4���.��-�j�L#�{��%�����̑�S�F����
!�N�s̾�^q��@ͷC�E�ܜ��Wl��U�,�{+�bs$�"2�L�m���+�A"�Z����Ӄ`��^n[+=M߸:��o2��R��ibjSg�\xQ��z�8���p�k���EDLN{S�����wR���p�1�"�F�Y��,��(iY�ui��Ռ��2�)�>�|�cY:�wܪPC��p���S���i��]�bݪ<\��&6�XI>��gf�f�	����.�=�yi���_U��{4wM[��:hi'*�i��:��6.�`ë��$�+�^ʗ��{~���)#|H���
���Έ��Jܾ�����sR�T�Ç�@�:+�9�T��e����+�ur.��V���Q�8ksp��ĩ��p���{m଴��76��{4*����c���{E.��V:b�c9hZ�w	;eޛ5w4��-Р���N�ڍ�0�7z�k�y zK����>��W<\�;����[�9H�RP��^��_ނ���hMjϦf�<B����[���J���E,�i[���uMPv��i4������^���C�ץ,	L��,���'%Wh�I�g*�j�ڽw��N�b����{qkR���=��t���Uk)��T��;*�,��ֺ�_���V�z�\~���:$�*|l��溝J����p���*e��۰�����uyA�œ��4%n�Jܧ9C�TL���s:�z���k�Y3��j��U}}L��.��P�����v�c��7�+�P�!�v�;~�<�m�<�G\�:��|���CV��,��KR�c
�M���2?��h��5��W�d]�β|q��"�=�:����2U�)��.C��3����i`F�JUso�]tSj���lQ�G�~�k���e��ާP���Ͳҧ�����k���ᄿ2
���&�O�Yر%�mʯr��[�^�V����LK�岵"��^�ꃪ칾�l��7 ,����	}ɪY��F�ۊ��RiG����y�\|T}0�4��	:��'�cյ�(%4���j��a������O����A��=k����%M=ъn�N��k��]�>8�@<���y6x{��ܻ��/�bT��K��3S+!���� �+��e�v{	n5�a:���Y�U�M�0��d\{��V\K:���M۔��J#Hٽ�poV�<8�y�TGd�,�|^�vxR���H�\�e������7L$WC�7Z���V�O�2>�\-u�ҩ�=�m��[��=|8e`:�^B�uֻȬ^�-���jeD�j��5y��u�ҬKŬ��L�2�FQv;��Pޓ���=���4c�]���2�W�4��ڱ��p�1���i=��\
���o���.� G���$�/��$�S@��<a��J��ì����B�q*�y���!|��|�y�ಒ�Ь�n���č�v
f�U�}"���ݙ����U�]2@�O��}om֤�4G�&wdN��(�9\ZX�ڙ�k��B5n�U�5�1��n�W�+���䙳z�c޶�(���8��u������ƀǑvР
 PP�DXHR�!*BT"˥ $X��AKP��-�MSk�k��")5� �B6�"�ЄH�D!- I��*A)"6ȭ�R*���Fd"�P*�1Ir\�9���"�D@��Dq�H�B�ɥ�ܑ H(RH�!"��)	�!��R��H!LE@�!�"*�B�)W2�S�d�H\�(RD������T"����$$��j�4�,B���́`DZ�
��
!$,	4] HN.$TE��*8Ԅq�6� �#spd�E$!R,m&BI�$,/ECl������TI� �� �Bs���A8л\��J��}}���`�Y]�d+��so��k��uFj�l[���$�x��rgJ|6`��	���^t����"�O�>���<v�^�t]�Ќ7�-����P8h�'n���Hgn�sT}�����j{�{�P�tڇ�{��3�w�}'�r:
�qrQ�G��B �ZM�G2��>����a٭�/=�h]�O��V*ħc���>;�:Q��x��u��'\���H�/��͈����r�1<�{��=]ؠ�r�[�>�5��z�'Is9��9��6<۾��9 �H�ӫ���\�s�����1��
3��`OK㱻)�x��ϭѿ7#�8�3���F�"y��W��,��tﵱi��	���:�Akʼ��l��Xs��&碤�'fI�gM����	���i7H	�!����$����k�`�uK�ՉJ�����<�>�^c{�33-)��+ɞ�	ٖ�N����z��/��Z��Af��1��^�������=v�V�]�rkG���T��+mx@p��5��X�f�Ø��gζ�>�I���c6��y)$\����o�vո�A���>\x>;A��5/�P�S=a
�_��R��rs��y	�i��R������|i�bI�;D!��}
���o�]�W�A}V�gs��V��D5��߽S]�{�h�m�P��-б�i��|��1��v����5GK�J�3����!�GLR�'�,ٚ*+;��������;�{���ۤ��������r�n��L�̔xl��PjL�(�Dj<}�?C���f:�K��Q��~=-�M1��l��-�_kK���!�VO�M��S.�l�{-iS����ꋽA�5o՝3ML0.�p��W�ҢIp0N��V����iu����r˝V;�D��=�X���#�N��g8�vT�vD@�əz�_�gt�X�Fw-]���5�[rx��~�U���ưC�Oh����M��\\�48�J�>�S˽�q��N������kr�ϭ݂����}K���~z��>�H^�s�Y:� =���ֱ	�]��J�t@�2:`b���ڱD��=��8�8�k��e�4�
�ER�ŵ==&�o�u�P�
�Q����ʀ�(�5����S���M�H��U=�����Ju�q�~(?$|_5�1���;�LG���,r���>[��>������y�Jg}�,���DD^��ׂ�"lq�'o�29�N٧H��*�N�p���q�Ay��i�2���u�;�c�mE�ӯ��m���y�Q���ηZ�v�^��w�����kI�!�GC������3n����/r�3��ʉF�h���1���\�qg&�{���1�w#Uv�BzlI�f��U�`��{���������������f8�u*u���t~����j�/��(�ȉ	�0'�'j
�Q��k���f���7Я&U��$��
*�V:Om��]��!E7.#K�v�,C�螖OW��i� mvb���b�j�5g�$K�Y��v�T��fo6&�Q�}sa�Yؒ7�'��z�:�k��ڱp65;�>�n�e��\O�`vۿXS!�b�����B��y;݁4�x�1W%�" 0���j���Z���?��̵�\}aC�Xq�Lwlo;6_k�n����\o`j�`nel_�""�ϊ���)�`xK5�
�H��ǡ\K�V��N���Vf_+�X�M��R�f���3m�3�|Ot+�Q8+��Z@8[�Qǌ�A'�f"�ª�U����9ܷ*���l^z<6�[�q�.��N�<��D,���WȾ���/1$k4 h�f�Z���.���8v���bZ�}�]�`�]�]9ʖ����n���i��"9�W�D8�"P�bR�oM��X�׎�_���{��>lФ���݂e��=F��WR�u�_*���.fj��)�FKQ6C굙V8��ʼ�`�y��6�DtW��:����)=!mMv8p���C���R�@{�۷]����48$�fΫ�];�B����:Hϝ0����ũ5ۘMLj����磌�s_�~����8P���Q�3#JG�b��]9����:,O����A,8x]��zns���q���S��*���p1�b(2������; ��l��F��`��9#]3�p��F�u�M����} "!�J�t�3κ��WH�z��UlيT1G&��6��]勶5X1��T�9t��m��Xx�M Adu�;&/.���DF���Z��·Ü������;o���xkF�%!�mN�L3N":�������O�s]�.	����Y�%MD,��s�"�
���ޕ��'���jy�&�u�:��#jVޫ�.���jr�$�!�4bn���"?|~����8e�����v��s�Ib&.�Vo��+�U��3*P�M;�*������d.�2���l�`Q�o:�i�ڿ[�|5�u8�裳�C;�sv�u���x���qk2�� ٪���$+�ە�6�a�d����A�մ��-�Qk$(a�e�b�l���m��߶���&�p����-W�RS���6귺ts�S������h
��ũ	��b�j>=U����	#j�b�, ��~i׍1��]��ڷ����e��e��(#�t:J��E�y��~c���:�#�z��OIT�L��yG�������9��o)Xoj~������MƜ�B4�K�Y��`���;�\F�I*e��碥{��z�l��J��z��!���鵗��M� ��:�lWH��(�Y,s�e�ۿ8�s�3o·B-��u�f�
^<�n{S��=<�4�'G:��"}���0M-s�������xl7-�|^�Mt]�������`��>G`j��;^2�$A��׾76����
�<>�ǽ��{���TWr�q7���~r#���=�8ϟ��о��N��P�$a�[�W�:>��<c�_� ���7�aW��nz՟�Κ#<Iö�t*T�����G��!�R�&����j1�݀�r�r��
F��U�_X���t3R��y:Q�߱Q���O�H�i q��d�p��>�NS�3ב�:�6#g�����@b�^�N�8�rg���a�}a�
6����z_s�$�|Z�0���x�9�:S;H���nG@pɶKP�Q��8���[��[O1�n!���!׍(�^���a�U���ᩚ���CҼ�4~Sԗo��䧛�5v���XkXn:/��9�e�J���.��T��ַ��΢����[����^C� u�͙]lf�R/��a���Լ���B<����e&���t�!p�v����Q�N�m�ɨkM���EY���I��T��H���"�X� {��^^�n0��Y���y�Ӭ^���:ů��>��˵ՉJ�|�A�[�݉\�׫�,��g�[�hQ�n�_�#�i)@_j���A��OTd���}B\�y<�Vd,�=O�I�3��=]���n/	[��*��x�����ʘ{#B�Y�n��ax�xa�b'Iw7è=NV�d�չ�����<͍�V�=�A*��z������sB�Ӌ��,���٘��g�Nչ:��'��*r�ʭ7S)��� H�j��SI�L��w�ڿvv5Q]�*����\���H����.�!]�||K�	}���6�=�~ĸ��·�|x���:0�\����u��`��W�_
,�p��xV뢸G@�<>k9�=�ʡJ���mZ��;��ɟD?k
�N[=.z#9�R�F�dD�|���׀H��}�&��O��g{,������&�c5�2���=����7;qrx�IT�洆���������=�X��dK������s�d3^z/�>sr��߻jƁ="����)ƪL�=�[�+{�T#���$Pڹ׊���B��W�v�m&sj��"�����9���ڳax������=���g���[T\-s����j��J���ei�E�� /�k���q�N���	��4�9Z�0V�<��z�ub�g����.��|�E1�x���i���L����q�q�06����`��2DvLD��Ѷ�n��FQ0`0��YRbĥ^���ʁ��8�����%;l�&��r�0�9�"-�Rznl�j�V�*W���F����12y��]r��B. �>�F��8��ƲU�C
�n����e�h��ׄ�T&�ʓ���DOa6��Nt�^"�����)���},��W0���O�R�n
���FDO��`HQ;B���(�&/��;Ԇ�ܓ��L�62������5E."Pˈ������3���n�Tgq��.ļ%�{=|.l�1��7���ג��V��V����o;�#,����\��z�n*�$�L53��ڙՓ2�#�(��q��n\^
�\Oҙ��n����̩�7��s���j5��\ˮrN�X6�F3H��f��H��
Ð��(�������Cq�:ny�̭E����QE��^�������m�^�8VH��4�*�}�<*y�s�!��ۅ�V6�m�dΎ�RZ����������r˭��u����ůH�0���f���������dO4�풊T�Rn��ZIh�V�S�ࡷ{�Fg���"��c������w�C�]w�Չ���NhY"s�mI]���������s��-�fc<�;�\�l������޹�5��<g�N�YtⴍS��gx;�w	J��C[:����,�[�S�¶/=}�~���s�_���w���j�;���q`�׌�6��gU\]=84��Ǵ!KT�������^t�N{�r�=�w$���ID�C���Q4WH�T(��\���s�e����F'��V�c;��P}[6W ;����bH%DLt�3b6R>�UX�yۯM����ov���yW,�n������H�;���
J7��wQ���B�b����\�U����8�*bc�k�Ö����ˍnwI���}(�Fx���D�"g�u�F_���!ca��
+�:�5�1�\���D���؇n�� �:�����s<#�"���JB�Vi�)�Q�Z;|=��ⵣC���n��i�GB�q����wPS}��I�>�N2ޫ8h����{����~ޕ�ǹ>�XmP��y�%�;�rY�W�!&�a~���94p[RLF!zg�Nwy��B�@�� ���Ho&cow��ޤvm��*�:��H�s���^�|v����8�.?~����U
p��8k4�o���4��xY/TĴ%����X��Y���=���{� R�7�ClV�G�d�\�'F֊c�mm�����/$-:��$�W���B��m�VnZJ4�ϸ����7{f��3��Dp���H�P��U������	���mb��n�L(z����W�=���w*�<Nd���ʁ�5Ѫ�� e��g8����I��foIPi�j"+q�q`#,�2��!{��n����WS~�D���+�>��u������(zW����Kʰ4����DpW�{��Z��e�Q���G��YS
'<hX^���t�7(���Vv��N��F��b��&��2�}n���@��ˍ�}�#��=�����Q�ȓJ���"gaX���,W*�B�>\4�pl��^���;d�mzy�|8�&@��Њ�Ui�GK�~D���p'V���m�m\����m���ǥ�Nf�gk'j<��N3�G[T�3���T�Y'����"Q�[�߇�m���,xp��lro;1SY�a��
K���=����p�yR��.J4#����B/����f��t�a��n z��v�M��b���N}�!�S���K��)�W0Hp�-s��ح�:d\�s��K<�W�jޤ+��6j�er��ܺ�9]��+��D=LSy�}nwي��#}�˝��w�.���o�W���F�J���e�����kk5�z��;u����*ķc�Û��r�φ�=���^o�W$yJ�%��
�g�90�z�6���	�A����2'�Ʊq�W�:H�g 6s�v�n�"x\�$:象�+4V_s����0���t]���B�Zus;�����t[#�8�ܼU]��D���j�����N�kb�L`DF�$s�Y�R!S�٬�]�gy��<�4ow�Lh�|��sZ��W�$>z��L���*(l�(����-}�<�E����_?a��O��������\��],0�Y�>�>�zF ��?���	u�V>u���u�����;�Ǯ�t<X�6iaa�f6�V)ˁ݀oZ���r��:��1:�g���WyS�B��&���ާ��K���:jn3K-Ps�ђE���)��j�`�IJ|��?,���߷��3���s�3�A���A�(��s��VUi�S<�G́"��M&Y3��[��W*R��W�,�#l積U���Ջ��6n%��K�'�ض��j�K��X]xQ��|6�ly�Њá��@�s$�Ǚ�oe��w+U]	�	�`8�#������Y��#R�h @Bl7���<�a��&o�Go��}Ԏ��sX�#���aV	�S��S���\Ǜ�Yx�O}IՃ��)M�y��|{D����q��_��Z�:�K�O'.z���bgf 1��ٷ�����׫��<���G1ְb�o����z+0�\#��w(N���kۏ@�]��}�x8��Y�2lҹ�Iً�=��RC7A�7�d�����-���������l�"����U�I�np����ֱYQ1g���i+�Eȥmp{J��gR�U͜�bR��3V�,����6C[������<,e�m�/!�����vDB������
�թ%��ٷ|Imk"��U�T]�V����QM]X��0p]���hv�|��ut�0Qoo�L��"�x�G�yv�g��DM[�o�WF����ٮ��+�ݣ�����4j��쉣 ����̩�/y����ث�2��3�U�ŉs�3ym�B��=� )n��5 ��wW!�ik��?c�]�@k���ϟ�=��kI��Y񠅕ǈ��]s�o�$�kH7,J.g�dk�[ֱ��x�hOn���K���p���[���1Z��0rS��������[J�i�Pi�n�]*ά��B�YZ�s��w��O���
+tp�ƳEj	Չ�ܻ�lM��t��Ф��O�/z�
 G��o-��gR�� �|w#���?�I�{TՊ'Ҫ�������L垌u#��7�H�����Z �_����:1�<��q�����Gc�27*��z��Ώ�=/���{Xֆ�I���EY�[t�Tk�IY�s��5nݞ��ep��&�F�'�׼.s���1�mszY������p����д�Ț16�
H\�4�V�9I~�yø����;��wڏW�Ҵv��y���,���?�,4y
(q1���p���8]�4 p�����Mi���(�ù�Oru��b����wj�pkS��6�9Y^�_����i�V7ar�^tB{U�>3=�ոgY����v�|7A���>4��+�x��[���`7V�f�}75)�dr�8̽���8r�~�?s�h۞�Rᷱ�l>�~y���C����yqY��Ω�wdb�;�5ݎAua"t��b,��;t��l�{����_n�X!VV�b3��B�;;�'��,l��E<��&�O�Bp�۔Q�-+F��U�>�wr�}��D���b��M1�+��Fv�ܵ�!��HcAh���|��R��[�ʍ���i��w0�Q\���-�x���� ��G���V;%u��!��\4�tj��8���������3r���&�S8�t��z�GP�kt���uM��	����.`�BmU��Rl��M�aΚY&�͇�2�<���������>o��S}���tN2�T�ڠP�	�����MQJ�E�6�i��s`D@�*B4��\���T�"�$X��i� �8�$�8��Q"��	I�!͑�EA	8�Ci��	6�6А��UN5���Td��#���fڠ�Nm�q�9�^$�*��5%ɳZJ "d�!v���h�3�cI�e���D��Y�6ٮ�$bSB 9�26̡��J�i���.XN2Z
�"^0��\���.A�C�nm"&ړ!vM!#l��%""���2e2L�I�D�"!��Ʉ"r�M�b�m��T�S�t���}��ngU�1ۖn�l��DӳGV�5ϕ��!�V�N[m(�;-ZgkJ8�-@q�����or�.�ο�}�}�}^1�MJ��ԙ�vH���>��5>���xV�+�`�<'�/
,���sH�j+:��{K�0��DZTn[=.z g8���Fő6O���o�������ͯ\2Z���{h*wp8&�!ke��a��6~�;��8 �8رoylA=��UR��!a<e"���,�{>�Z��;�x�Oc#���kC%st2m���J��յ�+i\�Q&����{&:"ǡ�p*6+�gVՊ�&\wd8�<ܘ��wj�׈�m��z�(���V��=��F'ҕz*6S*
3�{l�;��
P�+mf���X�y���{2�W{ʕ��A�G���C
��jb
�AƄ\>��ID�1|�n���>�[J"��,A�D�f�%R�48ʓ�虭�l�<�-Q�O����K{��>b��"�n��W0��>���2[��5�2*�U�tE/�O��P�3*VcZ1�5k'e1'o.����l����
�ۆ��0��Q^n\F��&�;>��g�W�&Tg��X8U��ܔÜ�W���5ɨ):��{D�T]�:���{�:?2;�>�&=_5�MC\�6ڢ�mոt��C�l��X�#���Q�w�ۈ�t�7�O�ED��@>�2%5k}���,�)���\�m�nĺ�k�}����{ܹk�[WN� �xm�����מ��;�+𤋮WP��0'�ۿ`(m��zg{R}<��9�{�sa�VL��7.8a�ٺq���\O�́�n�aL��FE<fiE;����P�܌�:�wbU��i���6h(�n�p�j�F���#����|n�3��#=�h� �;�#����݆��g������5|��neN�����Dǃq;$ �9������3+|ɗ�P�!DH�v��T�z��gpR�f��{]7����d�`Ϯ=�(��66�M��0z� c.%�GUG�&)]:�n��K���r�=�S�+/�Ӫ��'	4\�f���	!�AGB�vqt��8ya��-K��/ft�Z����	Ƙ�P0�U�A'�lD�}AI(�]"��������0ϴ�k,5�/�����A���+��e��h����[���~�Jx�x�~΍=�|����~�S��Z�Tz�#�I���}��TT�k���L��� vy��2��m��}��7:%�]�mW{���Lx���l��%�<S�>�[*��]��0��nitB]v�|�����p�ʹ��9L�DV+�G�0Zǽ�X��S����zP�w���~wh�׀�3��"�xvet_-��� x	���}8��������(��Jj�~�{.5��'��bx�K?.48��(wQ�~��P�X5v�^r3�)���j��tv�"�{U�95jr�	����ۭ���ؚGZ����j+��k%���h�5�,�1"uWQ��h��+���he�*M�t�ӈ��DdAc�Cc��΋I4�\��q���~T�#O���vj���������ڑ1H�&L�����t@�!e�y;��h}T<�~4�+x�Z<�g�{�N-��d-5�W��Xў֮��^e^s��ڲ9q.ܡm�d<� `��DWJo�
�
�v0*��%�>̜f�/ޱ�zo1=X��Qa�}�S��9y�x�=����̩�~҉ݳ>r ���
��9�uqaΚ��b��;m�En*-gY��u�Q��Ͷ�~���;�L���-���ad�f�+=VFie��M�ȩ��O`aDE�Tc}�!"l;f�J������Z��d%�t�nѳk|cp�1�f`�}�	�r��,�u����=U^�/P�D�ɮs̾�n��{L��n�w'����T� IRr�5����BS��%S4���Nm�wW9�HO��v�h��;^�x���:gn���7*4K����)�0��b\�M�a.��[Ђ��Qe�
�aLL���Kۅl�Y聆�k��H͖���Z�]3�/ �6x�u[��0���ު���b�ؓQ&�����K"}�����g��c���k0���)%%����&� ���r�X)��@�88��Q0t*���׾7��g��9�vW5I��4�$lKո��AҌ��Gi�a��}B*D�qd��Q �<g�ws�+��C0'�AuC�^��^s�5*�Q���`0��뭂"�-+)=��kXod��4��h��Q!io=
��Ak�rݎ�st����I��TE��|M���ɠs�:�෎�����Ä���@iy`0b\^�}�iwW�9H�3�8�k �a�c�4�?%2~���LW�خ����S�6	Bg�+�Fo��3`i�FW>�Fj��0ĵsTsY��j��H���
7�����6��`�����W���jf�²Su�s���.촬^c^Y�!ޭZ5��2�x��t�l�1��#g�P]�BWP�ɞ3EX�9f��9��L� ��_��?]�E���.0�[. ��9�yS��'_��v��f/7��Ά|��w�dc{�>��{yT��Ênj���CDa��r���i�Bdm�Go@-�7�����k���A���y���/��hRtJc�O����Sm].�^�w����v
w��7i*3r)��0QxM.� k(�\C�t�˹?����j�c�L���	s�lWO@}����xM�~}�<Vr���}�L=�r�)觮����5�nzs�zA��~7�j��kE+�{�y�����/	Еyq�5]��Nm��r ���:Њ�s�;�b�*@�f��r���M��|J:H��<
��,��%����ͫ����wh&�����5�y�
�Շ[�lܪK��?lK�ؔ�8}:J�K�e�ҁTj�ʹ/C\s�s��2峱:E�ޢ,i�:|�wo�p��K�+��/�J���c�f7�7D�mŞh��Y�ע+�å�ܶ{=N��g8�]�(ز"Ϗ�5�����NANM�3iuLQ����(!��uu��M�ưC�y&0���&�c��k��+{��,ڇz���N��b9��ճ\��W`�qOg�Z����F<Dm�W�Z��5w�i��+qvew�Wmy?A�r��"���$B��Tl$U�\oVՊ%�q�\��y�Z�ڜ3U�e�V�M�0)��sni���`��p1ǨK�)�)�Q�kWG��U�\���>��C��ޛ,��/[k�f��lR��G�����=Ѭ�I�@�����y���9L��4�0�I��_^�g,w�K�S�z�����}�dȶF0����/3|S�{K�c{��>�7ٷ*�>�Ӝj�a�WW/-"������x=ʍ��َ��\DE#���226�N����IGO�P�BG}����xf�O&v��
e��T�E�b�e#즺�(��,��J�3^�J�׸ʓ����mp[y���hNIꍅ%ҝ�+zT45��pL�ZT�x2�9�`dD���(��P�=�Շṇ7n17MQ����zw��B��ݰ�jyN86���
(��ixڸ�eSYz�q�����NY?_���dm��H{^t��)޵���&��m߰5%�~�=[��^b~��l|�cc�zҹTk�j�;]��d�m��9=�jn��1���{Zr�˛a69,��=A�mvn�Fd'�������>k`}��4<��|�:�˻n��ba��q�^��7Y�oeQ�Qw�\�|�
�0��GXηϮ�ծ1c6ヾI����t�Ͷ����ӎ��Ww'�f�N㵣b�LJ�^�a�g��QB�%��K�ov��MX��$r+T7�CY��;:m,�2�s��;D\=�d�Σ���l�,5�6���7=�79o$�gX�\*)�&�N��Qr��d�i],Ԃ�pOǶɗ'�.�;�¸���'�s���F��h#��wVx��æ�����g9B�)��_UUUI���ݚ�&~�r�<�I}@N�
��J����a����x�@�i����^��Ƿ�A��V�7ʄT9�F�^|�JN�yR�\�taUU"T�f�DP�u�qMlr��u���Y�;�үEGH�>�*;��Ԗ)�UqPt>��w�[s��|�kS�͠��*����� 4�4��8�f3�W~霩���V��U�M����m+�^�݊x�ל�(��%gV��ķ]�v�B�����'��]X��M+����koC�cyR��*d� �w���*S&(��U���<�j��t5���9m�4��7��TJ�L��:�۱҉ocDrXV�Л�~�[����OS]��"��w/�,���)h��uɋ�f/�:Y�=�Bqk��M���_O{Y7&t+vy�l4���m��k�X����]Q��K�;֮�cvd^�9}������6�^�]�m�š�ew;��nu�%V0�9�_5J�r�S(�uԝ帝����<��y�JAe�;sB���b���J�d<�Yu�1�@M�J����_D�HR�3�;swC��*�ζ
v;*�[�����\�H�*�_}_}��NV�7U3zTWÓ{�oG9}`bc��7�k�[u�|$����;5َs�vX���~��R^FX�BF[N��^���V9���ʳzT��R��'k�]J�L������IN:�7�GJ;ҳ�껻6�T�uK��Y��j�
;�1��tvC�w�\�xN��ư�an+�����̺�Ry�,>T߽�	��5�H���N#dr �/�ӨB���郂�"criv������5���KO���ț�v���/ӷ���������y?��{��uuJֽ�mB�ؗ/i��#eo����d������q�p-j��wm�P�:{,�z9�]��6��R�ԇ ��vO����{���냫��o%��:���E���6�q>ا��F�\ہN�Q7ҋ�K�)�������B�����I�kq�"�tٌ��o#Ǚ[d�Y5*Q����B�_^犨I{N5�T�������zބ�]C���'��BCWr��s����W����6�&���;I�V�}�%�y:D�\�/h���),�9��n7�ދ��<�'i9���{��kZ�nd�J��z(;FQ��"R
}4'�n�rt>9{�<R�gq�7�.��
�fyb��8��G�J9F��VV����F�6�����qs�*�i�\U7�-'���аN�!}�1P����^���J���ͯr'X��1�����XI�զ�؍�s��c����p;���qMB5��jb^ezyk�����`s�׉�z��jw;�����qR^�sܑuNz1�';>�Ͻ�V�ma�������l���;=Ϥ��P0��x��=����#�����~������������=K����Y��=����l�(�/�g������8�BUSֲ�
���9BJ��՜-vk��R�z]�|y�4����ڮ�n�{:�Ч�W>����{��^��W��'++�t������/�_���3w��Qf�2s��Ɵ\�l�p�ÍtsQDo�vv医�|�jXX��Q�wYa�n��P��r6����?2i���^�.�g�'A^O,��3R�q<�Z�Ӎ���.�!�D������2�qvo�A�뤡v����
o���=�6d��5���޽w'�U}�9����Vv���(-�X���M�����7����q��2�����y}���ؤz������:G�e=c��}��O/�km�-��ڲ�Ҁɨ[���1Hu�o����]o�'�ԕ⬇��L��fe)�9H���O_�k�o��m��x9FQ�>��.)lTjk0B�2�V�c���}�.v���2���R�3����Y��))P��y���fWe�N�V���W�AS�WI�^�h��8}3��pO�#Ў�h8���:;g��BOV[)�Л]�cy�Z.��T�Ið��#�S�
3^-�"�\��缤��i;��bv������1b����U5i�h6ƺWY�Q��3Zrڇ�hm�5�bBq�"�Ќ��KKk?E'=��P��̊���ȓ�nN�[j8����UM�j�Y�:DZᘍ;:�1n����jut���
��U��P�0�� �ν�3Ge�m_��51��d����,
g�����>��V��z���kΧ��l�`X4s����ץ+���M-��Z^PY]zgI�þ�ҥ�O4#��V�c���tm�o��]|��F�n\6Pȭ�;�WYT`���óַ���d.��<̹�<eIOI4J�&W������Q�!�(��
�}��=�8�|�oS�����f-���u=vTJ�Y�e�d�1p�O�9� ��p�>���[4�	�R�z9�Ѧ��A���y�?��/	)�L�}W;5.�<�3ܾP$�:zkx5�}2@�{4MC�kK���0�4�bp�W\�-}�����N�BW�$l{ÃCD}��;��Ɗ��7����7�ۨ+�݂*M1jWr��9��f o�R;`���Sz���˝+���+��0WP_19�67��Z*wY*Z{A��ӷ��zW�ΖnΦgL�l=�QP���z$�'��o����3Xb ����T_u��w�K�m�鹠*aa`�̓w�db�^����xu� ���.q[z��n�'uӪ!J�7�����/B�!>�w�������s��<Yc��p�~PE燵M���V�<��_%~)��g���/eK?_,wsz���.�6Ԉ�ï7K֏A��{7NI붕7����NS�;�}re�C)�ӱ���.]��- �p�M�;�o\kE��I|c�����S� �z�2��Kb\+�N�ETH����_
��h%�=�g?e�D^p{B��/g^�]��zE�h���ѽ`�w � p4끉��xq�t�㚈ǰs(�G2Wl1!Y�5Xb��yJ�Y�&7��AcM���x��}h�]�X�/J�
����o�� �խf�Lw@�f�'j�A��u�0����b,�Ct�!V�нc�X9��/��8���W�a�S�8�V��hE��a����5���s��r&����>n"p�|��q�X�4�WO��u.Z���U��qs�8qSnr���`܏.�)tMu$E	*��;;a3fZ�!���h���s��\�v���Lڣ�9�쇠���M�����&����q�9����z�g�]p9)J�_2�]2����H�p|���{e	f��}��U��->��zr]>��p@9vm�7{�DVK�o�L�����#/Cb��}`��MmF��7�FPa-n�j�W�sK�$�a�RO_)�v�6d#�Z�0e"٫�`�ŏ��\�mw2Dܧ��W	#�p��L�c|�5˅���C�U۶CN�W(�OV�F�Ԫ\����9Z�0 ��]���4[��՞35i�\x�֋5kHK8yQ]�c��v*w|8�؀�p�]����	O	\����s�f�1����D8y�k���(᷹@8Nķ��b�I�'��n�ה�Tdy�yzݥ���oe����Ƴ�|-�n���k�C��U� m�f!�I2B��$�d�����8��Z"e$��3�DN5!.�Ņ�6Ԑ�Y��,�"m���R3JIXBHJ�af�HM�x�С�!fa&[��V�	�8�m�.Zi���#4�HH� 3JK���C-ː�#mi@� �T��̉�3��[h��l6m.c��m\HTHm������v]
V�fF��B&�b"m�M�&M
�D6�s���ER8ƛ
��4XeBM�\���l�i�4̑&�4�i�L��lTHF�cL�6.��m���4]�͚DD \D՚l`�m��!	ɴ
h�ȁ��.\�L�\���&l��L�i����WUЫ�\�l�W.H�U�߱P"]�M���I��z��x��4>�d+��Uē7��x�oyr��v3&s�u�ڝ�i�����ec�=�[��*����7Sܫ�D�-� ��K~�K�a�璗0�#�z�MU�Jff������D��}Y�����t)�M���3d���I�����Ve�q�:X�䙵]�Y�{��D��%(CuX�7t��k^��⍦\�*�=S�%~�-X[�^�y�z��(f;*��V�cy�.d�T��*�)Dl�Ԉ<�K�B�}�X���z���-}c|��#l�E����1��#d>U�%'b��)S*�9Ō7����'s�3�s:�0��{i�-�iTTt���(�ЍI��飬N��w�sVu!SY�mW)���sƹ�^;f�R�EB��t��'��ɽ
���S��U�yC��fzu-}�[J�;׭�C�q�eD)�����U�7�ۻ��UW�\8'���p���q��&�����8��oD�\�&}zD���#5lfeMz/:~%OFU��PX��1Z4��H��]��V�T����Ub�Jh4�.n�ļ�XI�Tg4�>s��kp=~�V"���kɼ.�����˚��f��qWS��j8�i>��=�����:�pGaP�A��\�����(�njC&�Ey�9т��5��W�ʵ��s����H� Њ�Ȇ�6���&>�����s�W��=�Cb��i��������A×���;w6�����W�2��\M�w
r��1<����v�OfP�Z�A��1��i4�����i�u�ӝ��.��ʯk�t5�]�3��u
33'CA�V<����~�_P�X�/�ؘ�]GP{�J���36:�d�'_C�����0�\�kB�ԣ�;�ٞ~����.L���f^j��#��y<�'4��.��|��nr���
/��-7K�û���U��:����m���Z�gY���,�N��ư�a~�cZ=RH�|6z�R���y����퉟^��v�{�>��_]f��:���1��u��R�+{c�1h7�o�KO��;l�
Qϑ�Fe9�B�T]�f���uxs��T��ջH����6{k� �e��!2С�l�$��ݠo4\�׽�F(Y{)�)��.���̊�K��^�V�бg���Z-=D��81�|����;o6�ɬ���*��<�WD�E�.,�@��%���� �����:�v���:��S^��ް�X{i��͵B*:G8����BZ�Y�M*�B��>�Of��<�j}��W��3�pۈ�/
6�K{��s�����D7�B7���N~�~����5ގԩ|oCٻ
�yEg1�"�ۓh)�#�t��R8>)l\�@b�94��''+�zo�ԢkngR��i��FTJCb�O�N�:���[������ O�I�u���5��o�����*�H�Gh<�G\�V���&��w8���sg6�S�K�S/��'61�G�k�9F�Z��^T�bR�D�jT�v��O��9ݵcumj�V���i�kͱC�V�,
��b���zs����~���Jnr[<��sŹX�s�׉�z�;��Rh��<R�ʼ�/ԄUd�Ui�O�ӯFb6�}%de���nRv��='�.�G#%aQXH��Et��0�P���d�G�����v�+�Ξ�E�7���b�P��wY]��%�Uy*��Ã�� ��ny�!2��bM*̴��z�����o'Y�7�l��6��ڼ���[z�b��+��)���oXa�BQsu\�������t�n����7Q����ﷁ���<k�������EY}��/-����rʧ�:��{ͭ�iͤH[=ih�V��b�4U�G˴��Lr�7�'��C���4�X��=y���47��6�q��A;�h�W�^<4�w+��1'��tk�cq^���g���^TdN���=�1f��X5g�Wr2"b�_T��e��
�!��c��yͧ�[�3<���m�|�!H��1}�u�G����G�c�<��*)<�ˈ�.ш:�w�����]F[	i�JBc�w�I@�	8���|�g?j�J�-��P��c��w����[����(�0�w��� ��Q��3']Aܴu��u�Τ"�&�.[	���,g2(6�ל�(�	Tle�UP$^��o�.�2z������7X��>i��M�P������v��W�5/$��LP����Q��^��֙�q�@�Z�۝O"%��3^_���t�[�x]�Mw����d��u
�=[텝��m�N��fz7���A}ׯj-.�V ̀:�Ӑ��wU��F{
�rs��OS��y���,E8[,�7�hu�w��S̓�N�Ɍ��Ʈ�O��y=h��}SA���e�v��ZoJ��g�9��R����a��!�V�0�<�ŋS�ڙ�i�{{��A�¤Ocד=�}K}�m�z�]ڨt�*�%������Xb
a�=�l�_r���4�F��;~Oj�;7@k��gҒ��-���}�燼IY��ف�y�b��O���'2�tl}ioä�M҉Ѧ�m��d����w�����-'aL�q��u�Y���˳��3U�m�Q������kk�s�$������7-��]�m���`�����m7���j��b���DU.z�PK`����V4���<�Sћ�Y���k}C"��/q���b��*y��k:���V�'��2:�)lU_����iqi�ޡ<�6|P C�BJN�uB.�C��b���nzN�a{�Eh{R��gK�;˴zx�^��TԽi�9Q��i�류����d�E�=�%�6�<�6J�VWb峷M!�������4�bX���+��dĻǔ�j+�M�O^��u�n�
+.����:��{��|�]���r�K<����'��A�{9�-�iW�Tt��I@�s7���wf{�MW;b�MC,�J�ʳ�S��e�x�c��xͲ�z*�oۻ�=� �A�z�{z��+=�^���<�:���`��u�87���,�$���pb%�i
�g�g�@�W}}J(�jus܅��q��&����qFH��S�EM֧s�߸.�m͆��g�P���>+\����ִq.s]PNe��[�������J4bl��H�����{n�sY�g��9��^L`����\�װ��\뽩篪j�84lk�X���ʝs,�ڿo��P^I�Ұ��.Ws9���'�5V+	:��f��#k��V�7^� E�9K���x���j`�f���S�cs[˚o����c��k��{�J��	���&�'��j=���V�\o3�f#O4Iyڇ���2��O��9��'�T�u	U��X`գEq�txKk�h�ʰݦ�Y&[ޞYֺ-YZl��8*C�i�|2��u7�MB�A|[�rҝB�P�����_�پά��o[��!`P��o�w`lє�=QނW�������gm����-Ri��:h����Gz�x����x��s�Nd��ݰz�*s�$�~P�|�qi��cY�]�yd�����F���Kz���u�|UϠ�P�=S�45���Q,��![�ˤ���fשnSo�]�a�O�l�R��<��K藗��[ӤVVt�����o4Ewt�BQH%i%�KO����Ң7A�Ts���Fu-Q�K�ٹLI׶+�J��57�5�������͵B*:>�Q5c,K�i\u�y���&1sR�y�٧)����*�����R�̮v=��m"��&,�R�	�Ne$�/��+�l\o5�_p_M�������Gg��ZZ������7*i��,�0����	Kb�W<�:�qȓi���H*�&C����jU�:�6��;�A����(��J�l�o�:7��{4T�k���q�]�����4��n-��#�U(��v��G^yM�))���q���U���v�"�)�E�Y��/5-(��>�mq���۪P���H���&�z^���J�s'��k����!qu������]�5ü�Q�d �=����>w�^����/S�&"�S��)c������Qx��<�y��d�އz����W��je�}S^i85���h����O(�X�S�10�fK������X�;�Y�8�Սյ��$�z��m��q<��f�rvش��:6�=��j�7j3:���^�Z�s�ܬv9���&��w!��u�Ҧ`����f�e�v�Þ������:��X}6�+F>����r#���չ�����Qٗ7&�.s��eB�7Zǽ_r��n}Qu��6/���MɁLi�qf�K��fw�k<����r����qϪÚ3:͞gkm˖%[��խrpoXPsM�[{bWf�oU�gj�w)22:s2y;MڞQ%Z�*��U���w���w���/�Y�XfV�8Spy���;�W�ӥ���I�;L��J�ky~����z�������_lJ��*���V��r9�t��>FjVΔ�v��P����"9|�q�K���k��4����:���C�d�r���g�2e�B+�8�k��f� �1Z�ZAi�p�ݶ�yi�V�޶ӺbW�A�u^��{��7k�=��P�}	���P�����s��W�X#����/Sw:���돔�NQ��м�����*�ܵa���^I�M�{s����B�۞n3i�9A�*#��L�;����{�w�i��J��SU�CΡ��l��$̆��Y�G-C�k��}����^>al������{�����P��Xe�;g+�R��g%*���H����ق�?X]SH��p�ڽ��kE��M4�;�e�u�)�/j0m�m�lm�am��ƈ��̹�{W�մ���کj�TVm��K���^��.�iKF&ʭxc�v��+�^eN-}�w-��ytf$�SK��R�u��=}]x�f��;a=��;7�8S���m��jj���Z���u3h��9�Cr��2��LsX��W��וٺ���S�����V�6�F:�p��K���C-��g����\��o����]�Q��5Q���n�tv�O�/��,
�/�.�6|�R�VI�7S;�H-Y�� ����ZE���ʀ�A���R� 6`�L3�F���Wv��wH��^���*0e�B�����`���nwfe�٫�D=�'*�]>�^�<2�b̾����o_o{l�Y3��-��w����	��K�aBE�Lߕ&��-��]�R�
�o٬��p&Iۃ7Q�UHGh���.��uP�=S�%~�l�cq���b��\�{I��v1�5ﳧ2ʌ���6@<�r�I}BuT�Y/ B�WB�U���+��dα�7�[��i��{�c�Df��ʀ���v:������ӛ��9��Ȧ:������b��z�q���Q��}>(2V����Y�Mv�l���_��ئ�O���sƹ�^w�3��QP�b�N��1��W=ۛ�e0C FoEz7�̅�K_m�ҿC�z����x+�=�:�r��/���n	/�\��� F�<�kӫ��,U�\s�I2�e���Y��qe-�S&�Tw,y�*�
T#`�����Z=���n�m����tGMt֮��̰��w���"dr���:��4�=��K-[�>�|R��g>�@Ggy��1\tx��hj�+��_��_�-핰"ēZ���} ����R�&����uő(uo�yZ�]��c)��S	��U��{|��Ij]�������R��>�f	�v��S���-;х�$f_R܇<�$p��=��,�2�ܤGa��(���R�<�#�Ok�;)gfTˡ��v7�)u-���q���� �h��xO��u�&*����S�����s����(�m��S���O��]8�G�x�E�S)�z�
q�XT7<z�<:�<��?7�XH�]��po�噠��Y�
e9zĖ�3+�S1h���r��_e*l�X.�0<�[�U���LVu��S0_+���O%*�|3�.cZ�$���+ �u�=(�%�6ƹ��jsx𖫕��C�������Se�!R�F�6֋�-�Oa����B�V�4�M�8�J��|qp}@ ㊚���Q�r�q{z��]�] ��2�괠��d��:�Ͱdl��Ƭ���j�iз[��A���	z�h���)���u/U<Nmx����w�
[ �pB\�u�U�Yn9�����ko-7a�ָ��.��vM����<d�w.G�h^�g��{�.�ޗ�O86̂��[�`Sʧ�Ґ��aro�Q�^��v�[[`��&�R�-�g�u�&���u|ӂ��ǳ�_�3�5�<n#΀����w���+���4N`w[*�F�.v���;{)�Ȟ� �
���5ۖ�I(���_s��%W���j�0󷻨�Yڴjp��HU�)|E�-���}�N���L�iA�+�Y��n���T���Ok�Jg�=t�����f� ����O4{נ���˛��X�����Đ:]s�]��߸v��̽��f�hn=����3y�*X�B�f#X7�4h@��/{�ȼ��K|M���;�X�ϕ�ƞs�J���ª�~'�x��� ���d�	9M���Y����r��x�(��r���7��,�O
���.�����Q�W��=�|��=7H	�XH��,�i��!�p:��:;PWC���8Z���	�=��/�z�:hC�K��1��̨�
ר��G�[�i
]�mmř�e2� �u��,4�<(����@����C�!���*H��}�Q�|��&���'��gO��5u��WPj-�|	�嚞���F��y�1'��/+�\��^�2pԫ�9�Qeʷ;�hES�]��#H����Ʒ�y��d�;�*L^~ޕy�ހ��ZC\��j�Da�	�Yp]`X(�,[:�:��r�@ǷL����+��n՚��SH���	~���~C�������!7}�9BK�G.�����7�x��b�iS\��3z�'�Σ����L�\�g��w�뽸"c�/j�˗p��*	��X`����`<��+f�j��A۵�N�����1�w ����m&(j�.�P+lbhm�#MEʹdl34�ܰ��5V�K�bm��s]!9�sk��F��^'3����#)ni����d9���h�#&�mr�3fNs�'d٢@���1�d��M�"��$&�I�ƚaL��h!t\�4���m�m�.+,f,�j�1I�Ɉ��&6�Um�3$˓M��I�]22Ud�&��"�Dˤ˘�l�H��]�d�2F��f�%hБS$�d�ɠ̈�D��ch��6M��6�$�V�]tړ(�\�h�mfA�	��l d�f����2		3$023R�h�M�M��
F��2�B�i�hk�&DPɓH�.ٵ�"�.i�іh�Hd�FB&M�L���m��	�3!rd�Xd�]��s����Oߧ����v��<:�紫�������h�6�铗l4]�#�i���:�qo��c|+��T��FOZS��;�_�U6�����B����O(�Z=�q�S��]���X���OumU�';���4-���xn��;Fmˉ��X�y��<�>�:kg_��//'����N�*���11�f����V&�������%0�3(�3��$���C��v�^������$��"�*�z���v睸c��uG����T���х	�J(8J��������W������5�`5��Gv�vP\�;�.z��o]n�(J�.,naw��T����s{����6�����yȃ�[SsW�S��"m8iB�9i���J���w�m��i����Ң5�ΖX+c�I��ky�R��+��;�z�)S(jou��=����m��T���mZ�����D��2@=��#K*�N��9�#<����N�A^���趼��/��P����u�&����G�����J5�.�,9���F<\��s��?�^-�ӷx��gou�����y�`]�p��?	8�����]Ւh�zu;�j|:%�3u�t���lR��喳�ğY88C�n���+��C���ۜT"�H��P0���j�u���}�0-��Z&�F!O�)������O�)c9@9FB0�w�+���Q��g�,�j�ȭV��q��u��d�-I�o[�w!���=ڢR���&n��m��K7"9rBT�o*��*��(|���Z���	T���A�Y6���i�h�u��Uz6Z;Yo�=�}�V7���ˠ�T�I����a�#�c�K����^��;=ݼ�g�=aU�����n��U��N����؍�t�a�n�.��[�dm�5�bS��E����*yk���{^����_8U©V���I�ѣ��9P}�6��[�	u�Vg�.x}7+F>��kU�RIx��Hw�z�̬�-�T5��U��"~����_��Xqġ���|�Z�=��s33xTsE	��N��n3��u������˳�9�e��T�uu#���B58YF1Aւi��ݘF���7�����ñn��\�|fSHk��6���J�K-:.D�S��:p���+���Xډ.�a���G؍�J�o
!��F\� �8�3o��\O��h�l��J�*�����@MH�Ձץ�C�
q\�qb[{~�٭��gitWVS[{a�^>W����'m0z�A͡%uN���+�0��wͷ�/�>;s3�"z���>��~��q�Q�Pވ�P��R�(cwh%i�SUxI�$�އ�����dQz�s~���O]�B�	)u��J��^�ĘB�l����p������am<㈥�*:Gy􂁅޽�}����{����c�:c��ʾ��[����q�O��daOzK��ko0u�w%_��:�e�ά]�	���'q��v���
�b�����(j�UU���Mzu���&����s�2������)�/gGSxJ��J6j�(�Yb5`���k��y:�m������U�ó7-W6`�!:��;1<�f
���rV��<���_y�}�&���b�f��`�}s8����Kn��®�Qҽ�]�t�sz�Y�!��<ՙb��X4��t�Õ5�P���*�M���sN���LA�9����e��[B��"j����w{�9������F�&���������W�4Yu�U�5�#
�fXM�5���a���1�"��m<�<��.#�wԨ`E�Qy��c]g4�{ؘf��Gm=��f�k��#1Q�����c+0%����:ܤ�L����Ϩ����7Z�0kU��7�K:p��W��T�M���79^��2�j[M����]a�ͷ�Վ�_b~�$<Z���v�7���߇\��l�zJ�(M�L�T���˭&�� 2�����s��9O:��ʏ��u�}Qg�Ө$4��[��Ry	� ��}�)��z�����Ǻ�� ��g(R����#��/��
q�#�F�"����/z�fV��)�A�zޠ%��o5�cW��b=���c)�W[��V{���Wf�U1]Q�:�M.Oo��[~a�)�����������l��F�n6�{�14��1"c�6��:}4}��x�`�6�3�� �8E��9���un����J��^L��ׅD͸<hNc��g��L�Nw���S�g��#�y��Љ�Kd@�4�gQ2��S�%դ�M�{g/�]v{������׽׶Zl`c���ʉ�f����؎�6��}x\gpN��>��Y��π~Y ��7�7���W�������^�OvC�]�U���ͩ�a��cnM�9fQ�>�5"6#����__i�94�f�lސ��کy��LV��&ΊM�l�E��*��
�'�eh�On9�9`��S�rB�\����1���o��,k��	T�G(�
up�$�\�];\��|�~r�HO{w���4��mTе�lc�S�5ى�"-h�ps��s��~���ž�r\^�{-����Y�o�I�_�0�hFכʡ���Ƈ}�N��ܩ淖�U�w�W:�ίJ̩屹��ʷ|���c��1�6��;�m��'��N�"��XWf�8̢��3M��IY}�N[N��^�T<F����\Q��4���/?9�����-
�C�Bnr�����P��,b��#�T1Ӛ�d�]`6����gj�r߇���{ ��Jns��������m���L2�i�*�V�v��9s�S�l@����
Ζb���Nv��ΈK�D 5���\��m��{�u�\��s��{+���0�.���#�)}ub.������Ne�����I�\��u�I懏��$t�a;u��D�a�����	�-�|�穷�z�C��^���(��u����� uJ�Յ)�/��1�<�p��k�cKq^�����->�{>�ٹ��7V�\�ޥ�ȉe�����C��k�7�5����Z�x�M<�;ז�U��F'.�~��������Y�U�=�r�_�����O4��tVR���Lٺ�l5�)JBb���p�Gs�7��b�Z�O٬�ؠ^�4�e�;=������yWJ�r��3�����PN�E�e�[�`EL���SqyT�vW�i[7�`gr+ͽ����*����m�����S��ROV�{31�'@c�����~g�~�Gk����7;�flcl�5����Bork7�{S.��T�i8���p�5��Vu��W٭l��z&�=�xt�l�B�/s.s�����<Vu4-0�9�Ѿ��]�)��t=�p]fC9�9�f��>���><��p���5�W�D���o�ޅ0���:��߮���ۀ�5jUu��r�݉���z�+����L�0Ҍ)x��"���-cj>e���w�[<�Tח��Ի��/s5u��#pJ���u̳�mL�'~���N\֩Wg=�'7��Z����ٚ~M�h[���<oj�by��t��ޱp��Z3|g���L�}�u���)u�?c�v��I�X5�u�ͯy�7ª��D}�b�1$}t���뵮��]F�s��|ā|��2���o�i�m�9CTfs�͎�H�w�L#y��}�&���[Y؅��:C�/���曂�Εٶ��ɛz&%Y|�L�ũOl��2�a:\�;%���{E�����&��nܞ�PX�_c)�ع���U�
Z��k�}�g�>�}X���"���b��6��q��h��Tfk�Ư��#��f�w})�[^��
�yY;��,�,|��k�Y�<�+J���ϰ��ESvn�H@��"w�x�8,�]*��:�>�-�s�۞n3i�9NT�T)��U,��#wM�ݿ�{kve�)�Ѹp����	6@�m+޴)���;Qڰ������9ecr�y'R~I[75�P�X�ܹ������d��LS����M#丫r���3P'�u:���#�	c���6A�A��dú��8�+��සZ#f#4jÓ�'��ݤ^f�ޤ���?Xcs����]��J��dPm��,�Dn��T�;���j��HɈ��Тٹ��pBSkM��V}Ũ����1V�U<��q��v�g���Z��\��������=��ϫ<���R]����c2�a0���!TAތ��ws�Z~S��57W�aW>�{<ě�΅�v-�v�4c]�f@�f$h�"��ȕ��ۘ2���/N\�m*{��U�c�����h[Q�ʡ��ָ�/T�=3����������b_e<�7u��N�9{m1�c�<��Ue�X;�o3�C��}���5o��U�E��"�e�����2�X���k%����Br����I�K[>�tH��T=��V���!�E{���U\�K�T���!�r��[vm�����ӎ
hAΡ.v��x45�0!j��/rp-؍�8����������.��<e�[P�g�Cnn��������g�}3�
M�]♵��5r5�����u�y�`?ypڀ�	ε�كe򸙏��q��2[����o���]9�DU�w�f����};�Y���f���3kԷ���}���9T�1��Q>�p�T=��gD}�w�7�"�IWX[�l7vo�KO���깓���kc��ڷڟ�Wbp�};P��]Sܞv���w��ؤ�EGF��3��^�.�Wq���8���|Ծ^�4�}���6�E�Ù'���p�(�RBbߟ��
>��*7����-}^�����unԧe��gR�P2g2󕺓7*L�1|c�o��B��㫞`��X����F�1n���Ђ���|�3�x4;fQ��2#��<�]�w�1�z��w����|��k��m�;e��
���'[��,����Q�7)S�&h�.Sݫ��o��k��lk�!d�d-�wꔧ�8VK7�N�9\�z]M������V+	:��<B6�ʎ�~�w����[ul��4F��y�%�F� �=m���>�;T*����E�=��]r��z��P���<�	���1����&3��9r�Ǫ��WN�\c�]֠�f�t�Mm/�����Cq��p_2��C��ǽ��!�Ef=n�i�M��;��󹗱�֔߳�܋��}���g��w���ͥs��?/_�?r#�}m�:���]��zc�/;\���5��
��_\r�$t߽�CO�m.Of�vu��8����Su'�kO�C�&u����/�����Zn3��u�����^ʌ�s��*��Ĕ�����Z/k��ը���m�(|����U���}>���(=�"e�eۨ��U��̫\�BN#�-��d7l5�o�[؜(���>�Y�F������Ri/��#�v�����k׭����yoalYY�Z#�:�W%��c�U�jDL9��½��I`�P���e;��%�L��ιqZ�s��;�F�8�)P���{'��‍�_Nt���aK����Q٧�9,�n�6�s��Px�S�eS���pA��@��.4��^תa��ٹB�x����`��xNp�ݶ�G{��F�XH�g���u�s���ЬX.�M�؆�VQ��Jj��dkq8�+"ʪ���ku�B��)�=�X�m�z��T0��������%=q3��Ԍ8j�po3w���vU`�4�H�R��h҂R�L9*Rye�7{�i����2.ڵYtv�b�)���o>�۾TyF8$���3:��J�*5%��=w��^���q�M�k�*s�n#�=f�hR��J�g	����k�HwOB8�6����'�R��փD��N��Z�:j�-�kl�Z+�"x-^�r���m��Ҭ�D�pQE";���[� ~�M�'���ʚ��Ty�Q�h��8�+L��B�*���xs���8F@�<a����U����XC(��m��t8)gǻ6S!�Y�֢�S8Ͱ+w3e���]�󧐮����W����$���8m�ji[r�rSV�sU1���׻A̽Q��5��m����0����;#����2ZX|�T�R���2h�M�N63��9��+�:�n��Ԝ^�l���0p�9!�a�.Ǯz�"P)/I�!���dy�5GrŇRa ;�ϩ�Ƈ��\cu[��Qd7����-�ZI�:��� ��_l�[Nt�x#�C�u�C��IM�|Bq��}ri�9�V���rm�$ ��j��*�gU�C�[x��fݴz��1m�\����s�+O1�:�X��W0��+��-Ҏ�q��ȁ��}MD����y�G	c�!��լ��B���;�cT0�&��C���M�)*i`�ca��nB;�ج�w��)vf�r���;����,U�i�zl��뛵���Gp�>�x��U �cz�b���:e^�S�� ��s<E�DU郶!�|���d���]Ç����\[�^���n�K�'l�v$g�s�P�4�X�9���K���M������ˣ����iڠZGzH�e��g�s���R�������0��t���x]Q�����11gb;c���eA���bE�m�w�����\���X�)ŭ��{[�ZZk+,��y�.����:�X��/� ]�o
��ܙ�mА$�R���vCX>�� ]j�7<�P�3� �9�o?=rb���}U�4/2��ٵ]�}҈��K�/nl��}����KKY�ބ�^��8�)��%�\8��}ӳ�_݇�����X��6{=��K��Zto��Y]E��ɘ�Y�2�ҍ�WJq�,���c�e�������fCބ���^՝�`��Q1H޺x�]�r�'����/�
}�f����G�__X�V	I>K)+�0�N����͝U�J_m���o��6;�-;Ͷ�͠��BQ=�۠��Zr1�������\�,W�ih�݈���.�샷fd�<����K���&a3L�BMe�D� 6���R($	�+l��arF�fh�m5�e�4L�&I�6�E�4��D�lDFI�6$�Т&i[B�LL�(�]��6,D�S&�]ٕ�i�MZ6Id&��k�˒6#j\�m���d*m-,�0�Bh!�$�Jm46��r�Yv2&m�`���#$l�̄Ѣ�FM�%̲fL��30���L�f�m�D�)�Dh��D�Av!d٤�[]�T
B6�i��	&	���J����a#kr��i.J@�1�c21���M����JZ!��Y��2�6�M��䍛i��6���I��lDEd�\̳&Je��.Rd�͑�6hB�2�����l�eBM V4%D�PCA,�I��V�Zb�¦И�\�!#&�6�e�D����!tXB>�7�IL-ؿ��l�;�ձ������[*��=�]0)�S��R���y������eʽ��a�,d>�7��x�c�?'�̫�����k�Ԝe���l���*DT��C����R�O^C/�������σo��8�Xg�Koc#M��SϛyΑ�u��:�����ɬ�u��A�����	��ͺQV\��6�,��8u��c��0�4v�:��y�9�j��Nsē�G(���#S�8�'��{r4��m7���`�*���R�t>^rNw�o��1y�4p�=3Δ���ׯ�ca��2�<�QY��Y�Is�����=FT���x���&oJ�~i��O��{i>k�����(������k���/�9�O7���<.jhq�$���B���S)��z���m>ͬ�8_M��4��}��[�Y�Q������(Ia�B|�W4�\��Įͭ���֫���nd�V�cw|���o�N����PR���Ղ���xv;\1� z�����cla/zԲ�A�&w�Z�b�����:����>�9wA�eno��~f =��жn��W��!ƍ��}Ws)����ԑ	���k!�,�=��}�-�/�  ���L���Z�� [�=�u�0?W�b���W\s���G݄"��ӡgݶK��������'\*U)�P��Z�Q�;F,J���75�=�3��o-���w�Q����F��Z;��nٚ���P��6�Φ*kr-�\esy|�[a�-�󲂴�EGw�`(I��DB�[7�\�+��*z�C�4�����T�a��Oq��ͧ��+�Cy�kr�=��P����:���m��A֮�o2g&��U����0�M�%�Cxlh<�h	��B]kM���p�=]O�(���tԓu*k�\g�:#�F�B�5���[ɭh�ͅ�Yǔ:�M&مy3/��v��� �z2}��_��W��p�y<����е�Z���˵XmT׭4h6ƻ�3#]�і"�*�R˒����O!p�ub��o�����*���xba�ڍ�'�^�f��� R>�<��ClT�yȹ�Qe�����Pg-�}8��<)pgx�zd���dm���"��r��rʕ��T%ʰ����`�����-T�;w�����b�E���hX�̤g>��C���o\�*oJ�9w&�y[ �D�3��7\-�34�*K'U�@|�a���NOv�p��Y�|���{�u:������4�N�ܨWӕ:�0/[A���)J����KKG��V��'�e��	�i�[���P\��>S��(���ޭu�<��V�79BK}xP�J�+�T��f�p�6���C�f�oz�u��q�
�g[�+܎cY�Qsؗg6779��O8�����}��gݶrTF�>VG	T��W�L=w�R{�f���`�����Kt-���m�-=�{=Q��#C�]��h��ɥ����Ux<��v����k����5^y+��[f�껧���c]����	��W��|%��ԒҧN^�9O,sֻ<�3rFzuZ�b�-BQ�\So��QӾ���Z�,�_P���TW=Ό�6u@�3�2j�gu���r��� o��y���U�g����׎j:�cǣ����+p���Hb'��Pk�K��W����=��n-軧C���[�|�����f��'���-V{b{��O����$��@�n;%>��J��<�B��8��N�.���gnU��Z������5�W�lǴy��^q�m���ki�Q^������O76��/�6��:����3ySM*��{�9m�4�֢�6}��B���X6$�e�-�7ݵ��L7�-s�ͱ�+���m�`�ttj�bIw*˺�q\�B�n�M��uf)��r������3_����%g�t���L�av	�O���fuz^eOc����[�r���LwS��������~j�[�[�_˭e\�U�ۇ�pEh�~Bk�8'8�Yޢ�9eS2�/�j�����k����=r-O9�t�v�+������ȡ|֎-7�z���ód]E�p�s$�ݹq�.1�0z�1�.ct>��PS��͖�r�Ͱ��^�ˡ�87�
2vKѻ��3�N��uϠ��WP�*�,�ㅰ�Xm��>�^zǈ�L��f V��hh�Lg�X7m_]հ�>���Kuk��sjU���f�CG�Y]�D]{�L>��\N�}y�[L,y�>��S�Q�=�;~��p� z��������+�c5�93̧[�ׄd���!�1�r,��{p`�9��/��Y{'y�9��u'�wC������U���kٓ#�{ȯW��{/= 1�1x��h񳱖�Z���TTt��B��zvRY�U���$��Yk���S�s3\3�s8��������9AJU����+�8�ԖJܺ'Z�����'����}�%W��k��:�3��(���kk"������p�OWr���=:�wl&�f�,�Ey�v���2�����5����u�PA��By������s�2��P�3�=�)fSJ�i`�w�;�d�tQaUPڰ^��6�j��u��L�'nb���3�� �o[���`�!:��)ى�"
��JԂ�[篼��^�-���b�Wz���̴��A65�,��f$q�赵|Z+?@�v��h-o�>8���_���~]��>�+��O�;O�Q�.�Е|!��;^y�j�o�VR�SC	<�˭����\1�cMqm5�*&��F/6��2����BC�q~���V��
�$����V^R�7(�<���y:�l�s��wg$�3"�w�0h��'�OI�u��	�:���D����u+��DN��WZ�{<���s�%>S/l$�5��:��6����3	�t��k�ZM�S��Շ�	�G�S�-��e7%��n�l>�=�{�뼪ŏz�F��4�Fe Uȅʀ���%ׅ��7��pGb5�l��L\��r��kΣ�N;���A�Y���	\l�YJ<d���z��O4rY���4�������J��<�*���P��[���1QT�]���̝LG'��v���->�oxLu��B��xX���S�����a��_J�hu:���cXkm�-���%�Q�y�����B3��6*���H���ߝ>��o��<k�>�׌޹KZ��y�����x�b�l�c~Y$Bo`o5};�����m���Q��=ۨ�jk��#Xۓh�х=�F�<�jus��,T1q��P �"� I�+�u-Y��0��u(5�����d8��ɍ&��v�盢���hRw����##s����z����Q��j�/WA˧Gn�|��6��9����7W%ffᷓ�f=�tfҘ]���V������ n�:f6�f��/�u_^��*�Ԧ/of��a7���E��!�}��'G�����:�죞�<��tq�|�}���X��#�l�
c�=��.)�����;��+����w]�	uM|��5�Fdk��6D�w5������Go�XG#�M�o۫kUbI��a]�ʭvl*�a��.������Nק�P�T��z��ฮU��iq�w��s�ޏF'C���Bu��[E�V�Ӎ���CG]��h�s����ש鸊�Xv� vy�aL�[� [�;��Pw�Y9z����;�&/���F��Ovt7G����a��e��s9�X������B\}g�';���Q�����5���:rOX���s/=A_��u�����u��G�a�~[����C�9d�9�^���g�O�7|��Ti�8.Ԓv�g�=�1��Ep�/�����2��b��.mk�C�y�e��7-����i��ۍM��Xԧ���v������]�<\Z',�;^�Ś�s�m��L���i��AGEc�7���!�I)��&��G~�֯cGFmR�L��[��V�H}\�����gN�irm�&c����.Ӿ����r��qq8V���}n���;^J�>�^�@N(;*�&��4��A�x\T��}}�(ڵV*�\���_=���j���c�\�yPk�/_"}jхO�e]|e��g'�����p��E�I�G=��OG��y���\l�"���V��j�(�T@��2�-�~=+��D:������o�P.��ou�+C/���Cu�I�x�F[�Bk�2T�q %!�
S���\^xc��G�y�{���|ߜ]���FZN�>s>��Ϝ�`6۽�fr�+���òE�yӦ��/t{/�F�s�v�4)ҭӣpt�o�����_����%���Sh�\Q���eE`}{�ټOM��
��Ƅ�Oa�ޥ��:����vd�r�k�Q�feC�?�Oʹ�k�W59�I�~�U@��m�^1_D����T�߷i�Wx�N��:
f��38����$A�4�߰X���D�x���c��f��Z_f����/���0^P�(.,�]��g�j���g��;�:o��_{*c,�NЃ��6wh9��%�8Y�o��¼�Q�z����ǫ���)��Ҧi���+5���ـ��dB�}�(��Y�t�m�S����Lu�E�h�ӭ����7ObP��B�-���K�
Jɥ� a�z>=_�X�e�t�'p{0�K�6�*�w׏�qB�R��g�������3�����js��;�/�Q�6�\;D��.p'Y����	���m�����'��e@�%P�T�e��Nu�j�{�Y��_�p\s��g���ʕ�����T6������G�!t�A�@u�V��<�}N�;�W��U�0��op���{$ߓ՜�rj�������fP�@3����|gT�Wiuaz0�`��Hg�n�=�oSx�����n{z*y��+�xG�.ʟ��,���!�`�q��R7[u���b;�w��X�1�wx'��p�&�t����;A�6ttQ<t"N�3
��
�f�+>�w����͖ "
O��o��z|⛮���Ԇ�^�CΩ�PZ��� }5�����n'���v+����5O�v�_��gfڅ��������|�i����x�F_�i���`�^@�+�_��ޗ�Z�iK���h�ߙ��1�t���]<3��N�0��$S��&�w����}�����.�qߵ�!�.:�1XTD�o���\���
Xw��F_>���_Yg�g/������ ��r��IOb��Y�p�Ne}}��bl����a�h9�2ѕ�e�ۇ5��J-{�h�m�No~��Ud
f��N����Y����6F�=�`�d]A��t����וp����V�x^�"�4����k/i����\57�X�1�'S?�P�Sٝ��&a���0Vˣ��]�{҃Z��a����r��G#I�nL���}Ox�z��<ٞ_�f� ��rGJ'k�~���hzcAּ��R��/��V��Yg6�����q�����n�R�00�*ƻ��'{�|�9>S��e��m�ݹ��Vvr���v���R��n^\w��������;�9q�=b�����pQ�.=[�
�}6��wW�Aʷ��:����;�l�n7-\5&^ԜW2��A���~��l�3�~w|h��d~��=��YR�rx�
<|��Q�qR����;iY�)�v�T�Q�7V3l�seq�Lz|����5Y��c��ީeO�+���^��%H� =ʓ2:�l�&病���*�{����kN8�\3O���yީ�qe��+>���+�U��P	z mP���9�o"sޮ�|��L�1�[�z)�8����ʘ��xВ�4�����]R��9�L��ٗ�{����wUF���c���Cۄ�}�1ޟV��D���@���;�
D�.bHҦ�����{�7\�3+3�b�4�̶��2��AW�=nN�@oe��x���Y������Xn>�UkT��9&�3��w���~ޣý5���;Nr�q�|r�^�5��4ǿn�p�G����S��=W���^��v8=���Cn�ڝp
u<�IAlG���oG8��������;������f�K04F�uMWNt8u��;-�W�;t�!�J&�+��N��.�k�
��%
!�
�o&���qK�r:R����{7F�.�[�!�|�Z'b#d�[{��cWR�^pb���ah Y ^�/�ؖRN[t_YwؕL��p�t[\e�PJS3D륍u�1�Yw�8<�U/�ܺ��i��ى�K_K$�{j����H���g���Ǧ	Y��i5B�Iy[�K�&V�������/p�y�B| ��磽������~E�#O{p�nŻ�]=M�2Wt�J�Vw��`���ڡ�(5_��纭��$A4f��=|rVEt�wT�DBۛw�����W+��1��IS{(�������Yǫ(��͂�����|A��eqY�����,pyA!'�m�u��*���pQ�w�Za���<��|�7�7�j��fÆOX�z�_/E�ٲ��<����qv��0�<˸�=�K�=�����d���J�N�z��p�Am�ㅁ�tF,�[�������2�+��$͑�v�f��h��GϹj���hb/�<��X�|�J�k@��&6�Ĝ�L�2M����H��t�v�U�-0�-�3{��; �Y���i��#����W��x�\����/�]m����X�̸�d��:�w��ޖ�����.�9k}I>�h8�˘"�o�\�72O��
a�ENZ'��(�8ML�¹�Yfr���3 �<9����q�l��3j��3U���_eQ���g	���<ts�x�cl�qj���� lt�{!�s+��dhO��*�̇�syj�
�*Ыҕ�1U��8�`F�ݧ����2�:�ڋ�]�CH���h��@�-]�[x{U`f��x䦷��,t��wX�q`ҕ��hX{�+9��%)������=�%[u�T����%.�0c��sj��ܶ�l%�V�"<���r��e�ɣ�ڡ;���~Ȼ(gV��dHп��l��E��V+1n��ؕ+t3�N����Ș��wZ7����7�r��%��weK^l+:� A���d�w��y/ Ѝ�2�wz{���c����{%+[��X�_�������fw�v;�oSw�\�*m�"�&04M�9ۧ�^]�Ɓ��-V�8�Ԩ9!S4�a�����n�7��934=K.�Hga�6�l\4�ˑ���5�;(��x�cD�*]��A��h9��Շ]q���djw�v�u���s+X���MPqa0�����A.�%no�eq �$t�h�d�dD���4؄�3T��4li�aQ�ͦF����Vڢi��[��mt.��јm�I4ؗ�ډ�@M�4&m�6�%�fH���� �˴� ��I�6V�4I��M#F�*�16Bj�6�h6�&k2��i�3at�"6�D.H�P�d3@ˈf���m�&�.�l�!i�ɶ�6D�&�K56�)�m�3I�26֦�f �m��16ȌеCf�0�4K�cMj$dm�&i��26�!f�����]��Ĉf���)&�`D�4�mv�DD������a I�ld��يm2sE��E�v���4ĹF�,�*"�4&d!I�e��$JuD!HL���kR.�h��f��K��ȅP,�2j�(�	�B��M�FL6ȑ@��@�!5��!"�M��HM� �a�i!�d� Ddͮ�\¦�A2�&и��m�
?|�7��o�ϛ���t��ǾV�.�-c���&i<��>�\������W|�o_%]4���%��J���Q��^V�L	�`�A;9?�~������p�U��Jޝd2��'�7�p��gȫ�l)�H�s�����W�|����F�Fn�2���3�W-�������O:���	���ފ7�h�b��� �Kd�;<��|��N�h�Kj����֠�z��c���;�t��'q:n*�@�}D��13ζ�������q��#qƙK�>�y�����闡�J@�q-�Z�;��2�z�	��Vˣ��\v�ʗ4�1K������/�6��ƣ.�tm�\��� kB|�Rg��D�3)�=>#�A�+:%T��Gt��>HS�ON��ڥ���������<��2nt�|�P�/�&�لv}q�̱��e�����[�	��#Xs��*^����Jµ^\/|����K���T��噍�l�%�ˋ���K~��^��~�<\3Ī�]8�KÂ�i;�i{�x�:}��bt9ʿwp����5�[\��bi�/���@�dew���@w=��]��j�+����ʢ�,{.�S� ۟���"�*q�Fm����n�R&�2�F��h���g
�����I�FDyM�ZTݓ�G0&�t2"�q�c*aӡ�h�ͥԮl:{pN�ƵҢ7J��n#{�o�Z��^�=��b�;����stS�:�'��.�E{�X�:�xz�d_t�s�g��B��Ua�����Oն��p:ț~k%%�{��Ȉ�_u�rSrP�CWN6�G5�ó��v���	V|gj8��ݥg�k;j&�uv¼7m"�N@�}e�W��&��<�܇��z�\n�_
�l䝊d��sH'����uc����Q2��:	����1qZ�7]XZ�z<�2���z)���ޛ_!��u��u6�׹-��M��3eڒ�(	�W.*z��E���p�U���s�4k�(y=�ή�n��H���䣦�F�8^f}����I���b�$Q����WP]�;~�B�t��������.��9���Zu�GO^:Pt߃�A�\�i�!���q7g�Y�Tg���ۍ��W�����g��)ľ~`+��9:Ѥ�C�R2�RJd�� Jp�"b%*�w��\]O	y�#ڜ)�~z���:��x��e�'i9�il���k�mހͳ(�V�5)�,K*���6KqGȯ�h����F����>5ϩ��n_ϡ��%��k ��6�G����"���G�l�A���v�����`+И�^�bz-6�o� �	����q�K��/�(g�v�-?]:(<��ռ��k���-�VӢ�]@<�gW^x�=�3� Đc��ݫ�٬��vW�ٽo��ʳ� \�Ns�$��:~dk
n0J�f��Y�.7��>7�T�7�tb�N̛�9p5��'�Zޠg�x����=Nْi'j�;o�/�*%v^Eb�����ޫ�y'wC���ʗ;�	�����ܱ�-���~25�H:Y=��`��s���Z_f���6�fs}�9k[�;ԏ_���S+K�n�3��~M��b��z�z�Q9P�3g2�_��|Kz'�D��NF_^�^�}S3x�e�Զn#rձ�UOI�r�ԧ;�v��s�Q�7��Ý闆Z���C%�͝΍���k�G����/��2�W��j���3̢e��ͫ��D5{����89[�+�˷R�U���ݞ��gJD����%���T��a@waV��ṵ}�:l�_\f�E�}�"d���:�5������(��W��:P��e�UW�K�х�_�:C"i6�E*�z�y�v>�7o��\zc#��(߬�I���4eS�%#���j�\p�tN�鼫�^��e�s�l��!�u�aO�GE��Q'�%�B����v{�0i~�yH�މ2�"To�'��b��?u�]h�y�҉��b�Us�3)X��#$\w��!�N(R�˄6����r�G_s�ׯ�L�8��9�	��[|�C8-����N>���r�6� {[�a��������*3y��;��p��(>.��v��!����zm�T�S((OwH��I@W����T��wE�j@����V3�����������Ӎ����܌�4�ҙ��5���w��/K�5Ua�.�����ll�P�
s���ᾔ�#��E9��o������4��6��{/��)��s&C������&O>��r�gp)a����e���A��Y�l��}�v���e>�n�2{�>44C�"qrz�"d/��# ����W�v��z�w��`H��N����5����L��{L��fX���I���D��ꂶs�>��gm��.������l^�ݼ������e�϶�mMQ���ݰ4�^��Rt�z��ZF� �����}����X]9|{�qXWۗ��N�' 9+��_<���+�>ҁ��S��|Fo��j���V�kPw�C'��8w��L�R�jL�0�q\��Uz?~��g߿~���"n߯};T��K,ϞɔP����e�C'��83ꞦN{���)�v�T�Q���c���B��^�!u��iu�:��#���b��R����g6~���2�\�k���Y��SomuLH�053cUu%s&���c������B�<��y�3���;�����#�%7��+��C�\]qq�����Ei����,=�2�+U�ђhR$���D�k��in0~����+�o?p��՚��T�F@W��i�6�P�P���ײ�*wN8�\3O�ok�u��ز���;P��u\gT���j���矎���S��;G*!��R�ϭ���ntv\��ܢN�9�A��Y�J�(����8[�n���N@:mk������9��ۄ�}�5Lw�գ��z�P$�]���z�ۯ;�WU���EL��+�J:�U�ԩ���!���d��:�h6��W���f��7יX�ܫ{��2��3�Oç��)=���NxWKw������Iø��O���'̌��;@�r�m���\�ƣ���F@0�[$<����q���HY��ӓk�W9Ev�U�/F��t����t����J��"T'I���[F�eq|�b^��wЎ.�5�P|�N���r<1j��\K���M��@v�'!L�������;$L��G�
39�F$��I��}�.�P�>F�q��Fcڗ[�m��[�П �])3Q(�fW�����3�;��X�sT���v��U�3�QeTl��Ǟ��1r����M������b�����+��ʑ�W��3Oy��,�̩)�/��r��G�"u�Os�aα�ͧ�H]�(2��G��A`��^8H��w0�s����F��S7t7���.��Sɓ�+����ק�ս��g����6��ߔ�&M�n�ք��/�'%t��Ny�{�^�c[�Yv��˃s��>
⧰ชǶ��v���U���N�bq.J�9P�\�J�=^��=���w���3�h�z<av|2�+�xpO)�swi{�x�s�ފ�v�WK�O����d_����ao��c�޻j̬>'2]���kҝ��c^xv� 2�_T_��[;�o`���y�}T�Q����W��i������V���#+�_���[XFGU�q��T�̎tM�O����f,*�ܜ�CWNy�]ϭE�z}'o�O����|�l3Ѡo��Qz1�Aڿ(�S<]t���;.���d�9�^���g��>��~����N�zK���a���?�;z�߉/�%���4�L\V�M�uahr������l쾨[������s7���QV��ExΛ�� �<����}}�(ڵV*�\��\:C"V�Pi� Pw��jϺ�����ϛ���q���y�*�� w,��t�����������䟩F��ʔU4r��G������w�r��m�Vl&{㺪G��y�{l|���"��������p7ٿ3_NY��e�u��u#>hd�o+��NtfK���̻JBL���y˦����܊6`�1�ǽ䙗�:���������s.e�s�l�>��oθ6��b�g�*2� �\M���{E[������k�}�*��*ˈ[��%>� �_�N�i7��R2��!4�J�� Jh�"�.`}"����ꓵ��,9�=�Fq��c��'iC����C���w�3l�|�I\U^^*+n����{��T�uO
�u>:7>)��ƣ.9��7�r��|�q�П�2�OW�k�sU��#�=,�ƨٰY�hM��6�ޥ��:���1m'fL�5��Iщ�/7�^���t�
��d"��<9�@����K�+�+=7��Co�Wx�1����<���T�����C���/��v���ו �d�L-��B�Wպn��?+y�G�r���-�B��5߭5T�����:�p�yV:�d_�%� �s72�鞒���y�?V8k�#$����E��cʪ����S݊���o�˕�jg�0�u:	���3~���;V�HGF8�Ua���d��dʁ^��L�(�R��z!�q�膯x��*\�����J��Mz�l�EͲ��1��8ms�˽4����a�_i=���V���A���gU��bP���
�3m���[��2���)VέQqa���X!>ciX�F#�]��s���,-��b��P�\�<M�N�҉��
z���|�|z1��̚!t�8O��gG]J��J��vJ�0�`�s�e�.[8Ř�'�.ӳ��/�VK���i����ŔJ�P�JS/��Z�"�]XX�G�C�����zAF�2�G!5������l��G���(.ʔnˈ���0T��R<+��W�^SZ=%������c�Ɵ�/D&w�آ[9�C����ӣ���_qD����yx9���։���j����o����:Z���S��r��C�!鸇�R2�U �'�#� �}]gҷ]�g��[��̥�5�o@b�h7�q~�X�>�{P�[���{Crp���r2��3Y^��s:gT�����6YPB9R���n����C!q�upҝ$aC�m�r΁�}��:����Y?�(��o���^o���ԫ�O�2��oV��₨�ۑ����7J8D�8|MJ�z�Q��e�s�~f� R�Q5�e�뉐���E/��6d��yʜ<�{��g��_���S���}wB��d�D#q�T'�k�����TT���e�99X���/kIއ7T��ρYv�ȆTWڶk��U4�j	ot.WP`�ܴ�VmA���c��>���p,~�6��y�<�Žgto_Dz���o���FZ0d��;y:SYך �u��Ac�7�;=���S��-�}�N'�����;N���Cj��Ǔ��7l/�U���k�OT��MDY��ӽ{��;�'=��N)����/�qXV���{����N�ro�;�9|��.4�L�듢g�jԻ���ά�^K�s���W���ZN�Fl�w)T5&^i8�ef��<ǵ_H�m?L��N.Xt��Q����f��3����|?`Ńѫg�����k�<ס�|�����S y��&���.��0�ٶ���+�4�?p��^[r��q^��u*�}��H�ط�r:r߽�����Yj̇z��t��E*�}�p���S��{���3�
��U��r��4�UH|�U~�����Q�:��E�a���;�>��23.Q'M}'���.22|o�x��e;ӻ��n�'Fu����Y�Z��z�xq���ʎ[.��;���� �=�g[����ݠ�:&�M�p5�u�L�=�E�j�U�jV��5�eizJ9�Cθ[b�q���
�yӾ���v�`���#�3>���Cخ��;u¯�n�`�<v��8VE�V�ʧ���Vn�,56
ݘp��V)vj�N��֕W�{�/:�by���>#����VGoSr�6\�G�Ly�)rq쬭h�ӶĜ�u^�X�P�y�ǎ����l�q��o����-��?N�"�̀�v�uG:���ۀ���SN�r��3
(�}�@� R�"��59�����q7�}wJ���=k|���/@V�F?���n;��n�D�#%� %Bt���u�n�W���IZv�˽�@]��ۍ��	5h{�.���g%�8�󸚅2�z�BF�;$B|=y0�v=�ԓ�1�.�o\&oZ5iu�6ۮ�,����ғ5҉ЭV��&*0/Mz��k�zh9����¾���W��vϣzV�O*|ڻ��y�'�t�&FC�xn�3���x�:���2\9�T����
|�Oa�8�����Zo�W�	'U�<�J�1#}�w}4=�Et��"���w�m�>:=���e`R^�U��i�U��ɀ�nޙ�e㱛���mC�7C���Bw���kީ񿰢s/�3�Na�u��.����Q<9wY��-�p�[�ǝS�fS�g�s��^O��Lb,��C�G�A��؜U�޸����h�*g���."8bn�XU)�9N����]紡S�z�.~%F�tgԟХ���3�G2��\��\�����I��tkAUÜD]���Z��]=�=��û�&�������.|��'�.r8 �r���V�94��ޒ����$�'\q���5�ׯ��g��f�!q��PbYRх�v�.&��LY[G��E���uآ�P��y��A�#n�7�qV�����;��1L�r)�(B�0m���KM\��[������Y㷜�r`n0o-&W'�x��y�V9�5�3p��\C��w�i�ޤ^���iv]�=��Ե��xk���*SZ�]GC�+^����y����:ʜED����H{�yk���˘�f��e�^,gF��\t[�˲�	E(t"���qM�n3Y��c{6�pr��� ��Ѳ�V�!V;��K03iT/,c ��]��,e��3��W�J}Ɗ�]v�]��S<����0��H�z�{��0�|}��4�3�'L��-/�u駈Ҷ �]M�����Vf"�=��-�l #0wVvf��D��1R]�:{��-�rS ��v,^>�ŭ<�L��F���G{Mv��S�6�[+�j����x��(�Ԅ;g�o����0���ˇtl���{�GOnݏ	w�>��>k����6�r������8�{^��� ���T��w���d�t�ܨ�=4���7�3ۛā��֤xxb�zY_l���cWS(Lڔ9*�ѕ�9��W����R���滝���\l�%�vܾ��P�Vt�r�}�Qm�U�n��M3,�%_�K7�w8��`d2{uP��g��x�:�()����j�1��B��=�Y��.MO���,���� �~^����+t7XB,=ܟ5�����p�N��T�;��Ep<���㠣���0yIC8=��k�|���D�vZ&�H��nr� <���}ހ�ƛ��T6����Z�\)b�è���4�@�o���<Y��r�A������x�q����:���O��n�ӄ2�)SL@+��$AJ̓�c���yU%�����ݏ��g=�H��)}R
�s���Qs[ҘZh��@�-�m�}M��`b�v����\��QD<{n��ś�4���ƛ�C��t�[�;S+���׷&�_x�%r�{/đP]�Ni�|�<}�.1�>=B���?[H�~Oe���i�V�6�\O��8�2E�'ܽvq�z4�U
�v�..��`N�g�r7ͱ���-jgv�N�Yh�G�Ƿ	_oN�CY�V�=W5������M��kANTai!Y��8kgԓ4nvWWp0kbΰW�J[f��`���YuU��_PLU)�ʹ^JY���:���@S/:M�Y��z�j�\L�A[d(�Lz�}�!+�`��7^]
�:�P,�(m�K���U�ܧ�ޣt\c,�v  T�$@�Hk��C!$`��L�ͤ�M�e�2 ���I�!l�f�4B�!��mq���M�H�h�Ȅ�i��Y��a�5�E$A	�� PE#4�D3TDf.Y��m�\�2���2L�&"f�D	��HTB�*� �BE��"���m6� k���	�X!v�&�2jA��"@�A�$DX)3
�r!PDQ����%�j�"&I�D�A]I� ���0��T��"#i�#&�Mm3&3 B�Ѳi`%���\l�L��2�mH���X��2�DH�"�D��@� ���M��H�0��(����Ѕ�	�J� E""PU�L,DR�)R�D��a�"R�"! �����u9��e�-6�'u�s$wOc
���Y��r�綔:j�8�d��vk��1�;5��!t���ӛ�� ��\A���ҪF�e�h��
��M��y���p��}Q��<��>�����T���s&�\ɠ�I%�L�UgC�����j�T�B�V��`�G�^�gN\r��5u]�\(���ϸ�;�,�[��@L@/��OW3��QER�����wl�(ߌ\������
�ѬM�я���ۄ����0��~$�."���1Ge%9�� kyl�5/Fɭ|7�K=/���5�����;~u��R���(��D�a@�)V��+��]^�e���V��o\Q�mk늿��� �_M�u#/�T��B�*j8�����i�C��z_M��!�6�A�=��DQ�qq���'iC����D9��m�z��3J8c����xݼ��ut�d���58��$LO*�W]K��Ϡt�n1������7/�e��K����5i���ѱ�і�D����~^*u��yWi��X{S������<�VFU�����f����fK��k�Q��ђ}�N�L-�/�
��T�߷i�W��<���y�.��+�<�}��ݭ:N{��H�J�&�~>���|Y�7�W�\j�];2��Zm_�:�ſ(۷Xk9�I܉�H>X׏���v��Y۾�:�uVv��	�K�Gܧc�Ku��2�9C��gCJ�d��Q��$Ɋ�'�v{o��pk���)���v�9��~�>�d�@������s�>9��b;��U��o�]T���7敱��r�ls�zz#�����)�hg��T�^J'(g�ϗM��U�i׌��6��9^���]�IxO�Dv�f�7-[UU��:��;^�B�rnsE������ޫ�h)���AS��W���)���2�{��}
��,��s���WՓ+]'�g�_)�ٚ����(��dˋjN��=BgG]K���U�0�;��`�G:�X6����^��yc�Y�xݵ�>Ս��"+;*t�2~\���qqS/��j���iua>Hzx�:S�]�ÎߥP!��!���ާ\xϴ� �*Q�d���FU8�T�F8|y�\�]r=�:���1���׬F�?��{Kg<��z� ���tu��ƣ�$�D���^$���������N)�$z�Tz����ҷ���CS�{D=6�FZ�AX6OA�۱j*gט��>�@������\��Ez1U���V��%��>.|�i�nN���g��v�:c&&��ᜍ+1>@4�[�	��yh�JS���eeM�YG�8F6�J���b�ݝ)͋���8�fE��b���cEt� x^��21>�h���)mc������>})��f�"��[������"?u�G�m��^-
�޺FB�C�u�J�&R��)�3 )�7��o��N�1��m"[�R��O�&��ݾ�7J�=ʢqêFB$�莩���s�W3���\�J���O�*�y�et�b�|���K��ÝvY�9�D�C5����2���&B��{/��;��k��"A��ss�߽�ï�|��!p�]иiS%��`k���`��A��D�@2���T�i��y^�����\��<���ݸzu<�:Utn<� ��`i~�,��d,��}��O��y�����M=��s���x�VOi\s�V��ܼ��rw|q9�^wPs�����WQ��n9eL����:
. �X�Áo��c/��ZN�Fl�or���*�zc�8�eV�p�􍮉B8a�~�]<F]86���~6��3�qŜ���?P���*}G��~';e��on)ɧ��k����c����ρt�x������|����:mN��+&���T��n5�jq�mT�*ٝ���ڶ��v��}N�;�U�4����^w�tݖOp0���B����FtWK�ׇU
c.Q)i4$8�j��7�4��� ����u� 7�l�������8�nit��͊�T��,
qj�J�U:%����v�>�U�|�v3�)p��W��Z���n:���B])ݥ���U"�_�)~.���u�TV�a^�͙Y1�U^���nv���E;��{��h��r�:v�������νo}�TOU�řʎ�3�o��p
7U�/t��!����>�jXމ�h�t�/1dԻ�z�nn�&��	.��@H]P�R�=}tQ�j�U�V��\�V�|�J;M���M�����������o\,��g��e?�fll�P�+�g���
���ႋ���f]�6�3Y2�KnN���r�uH¸%�� wQ�)l��js��s�@�Z�����+�%`��_;`;�C9��%㨜:��M|��j#���@�&&y��G�kJ���{�Q�F���Fu���#&�����M�n�~wP�\�@!#��\u��rk޷�'�Q�� �����o���֍F\%���j� ��F�
�t��m銬�ҍ��|��7����D#c�=����M����ZoSۇ����dɶ��p�d��0��tv���X#�H�*ө�\6�ǧ��a����	ۯ�eo�J�׽�N5�ı\�cA?Ó�n�1�u���N"0�`�O���+��~�"�RC݆�R�ӑè���H�xqU�}��q�7'��5�����}��2�;��ȈZ	��ei��ޭ�eC���'��N��1�%�.�R�ZsCrv��F\������M����n�IH����:���id�L.���]KÂ�V����A��dQ.��ӕ<�z�X���O���s����O=�

�f��D�_�c�	�0�+���ЩU?W5�����jff��� *3�[
e�3=�u̯}άn�F���e��z�Q9�ax������F��s����F׼��)�i�_�i *#ܕ��y)*�]8uг�֢Ʃ�=���%�}���ס_ۮ��Z�Q>h�	���9P�W��p>�;.�.�7�z��\n�8����'��V��YN���IB�$�L�� L�RK錭T
��k�C�G�^9�����*_�6��>.�����}a�s�{�bܐt�/�S�����QFժ�S:�&����o�����g9�CC���|��;6����V.O���4�Ex줦qؗ�9�u�d�+*b��>>�_y
�Sw��KGS�8v�θ7�A�%�#䁐�pZ�&e܈3�%1;���s�v�Z%�\�{3��3��}qW�{�����N�i7H�uHM)���.?}��Fpq��d��ފ��]�Ѻv�ղ�Nl���*d�C�xgKĎ�R��q,L+�ǪBm�������xBD��Z0zŤ���V�5�;��܎��$z���;Jd�����@+�w+�M<���Ֆ��gX���J�>�;z�N)�+���n�쿋�&' cK��
c�Tb�Q���G��}���9��[u�c�F?jڙ�}�^r*��3���,����Dħ\*���\tn�����Fs�t[+IE��.�z�|�x��e5|���H�p�`�1zh���GVE	s���+M�*|lN�<�n*Gܬ�]�(���ɭƈ������2S.8S����5Q;_L-�/�*We��Eb����y8U�ph9�[o�ѕ��b�Ѯ�4��\y:
f�`�~3�yRG�,��[�sv�3�wp\�>�Q�~�7�YZ^��z��{���=�:��؝g�Ճ�~O*�]̋�J'/��\J��B;=5��ë���o�4�-T;�R�u2�>��S7��aL��yLgl�WPr�{A;�-�r lQ�Y�{��}�d���.e��s��z��<��~�P*>�5p��i2ɖq0���}�,������:�e�o�W��a��p_98p�/�	�%���*���d��*`�n�V(�yKȺ>���b��h�."�${>�c{ u���ʝ5��q�K㵪�(�e#3Vz}s��òo�"�j��3��n�P����r�:}�e��.o�[L1QϨ�w�1�:��м�]������_�rZ�(��kp���ކ:,�P�B�	Ӫ澹���<�[�q���&@���%t�_R�&:6���U��#9K�4��pt�K+�nmO^S��:P!�C�3��6{�N�|��"��FŖI�C�ѕN/�=*f�zŮ��:1�������un![����������{m�O�ӣ�\�5Q'��p��ثɯ���z&����pVTm��I���p���[�o��jw���znuH�UH)��g��]�g��޹�D�n@&���O��`����b��S�-���;��'��^&i� ���*�%�mˑ�g�\t�<k��=R艔�A�)�3>
s�����S��+�x�Ƕ�&���Bk.ej-��p���s,�ϔ�F��a+DL�}4.+�s;�K�Ǻ�c��ϡ�w��s�i�ǯ��}E��q��3Q�)���eI�1���T��E(�?M�E�-`�f��4}��Ϳ��
�����}wB�T�~fX���P��A��N�!i���J����9=�'/���u�gq��ۇ��=�=��7�y:M�v���U��_�A���tw��ܲ�$g�;{�e[�:�����'î)Va��%�|r;�i�ܼ��Drw|}��Mǝ�g#��Et��`��m$S���W��*	�'T��إ���zG�&t��[�u�3@�J��c��zs�{�[g�%I���:ء��5�E��;�w{��q �����\�R��n�ξt��غ�������a�n�DFj��T�+�FX�������u^�������t�X�Áo��c.+�i:}�)���WI��:ﳡ'yL�5;��\8��?i�������K���,��,~���I����U���S�r�gX>����(����yŇU���Z�z���8�g�S���s/�0�Q_'�p��Պ߅�R�y8ޠo����<�s�̅I�E:l���:���ӶY=��^;�^3R}�=�v�в���vۿ8�N����@ڡ����:��[�{�w����>������v]��K�_�u��	4\�f����2�Η ���]���O��^z�7�-Kӝ_{}J�k���wD�ӱ� ')ON�L��B�����E��Fժ�W�[��rZn���ޖo��f�V.�����pgȫ��]�e0:y��)=�+�g��p���� �6�6�n{7��d����8�N�x�'�0��rQ��u|d�[$_�g����靟�h>���.�w�B�.�4� ���������A�,�0!���F ����:�����c�����N���J����W���9��i�[ih�Z�Ƕ���ݮ}V+}H�Rm>�RA�� F9ZZ8Cp�X�=a(K�|6����_!K�8n��}�37S���3�μ��B��f��� �v���~���^+T�A�}%�`�'��V����߶���)95H/���[��ۭۨ�S.g�7ݐM��c���F�pT�1:���t��q�p��Ѩ�K�Ѹ��p/�� k�5�N
����zl�k٨\�`w&\B�J �Dq����U׫��;�a�On�uS7�<ɓ%t�4`�q{�;X��u�
�PA���l�;5��l9�R{�}X�ؿF�-7���{Y��G��S�W��U��VBlJ��},A��yf���,����\�
��xp\Er�'{w������){�=ӽZ�[�w��5O��N�9Y�����ީ�(f�2��C�S�\,7��1U�S�N�H��r�� ���ʩ޳)γ��uct�#^����Q9��+\.^+�������Z���Q�^��$��]�4�"�7f-T���:�q�]>[|DV�n>Wc�[��nx�c�4�@��蓲:�Uq�(C���*���|�2��^�z�|cB�\l����'���V�8�p��{M����I�x/@�Ф��Z�7]X^�.�4�x��vr�c�U��r���E�=齠r^���b���jfX��tw{1�餵�T���Ͱ	n��cV�3%�h�pq���uY����{Z�r��q���t�P��
�.�۩�+j�9��u�`
C�J�|.%u?�F��zu�����Y�I�?y�-�����g8�=�Q�[��ˈ��\X*��=k(��`��|s�}u�9��{��S����T9C��v�p��g�¸'�I���A�$u/O�y��ǁGz�k�r��u�[��-;�������8v���U
�\�k�"��{��ؼ�����Q���F�Ҽ¨�7���[���9�>;��&�x�F\:�'��}�fU�1e��iWyW,�����I-փW3�.3�븢o
E�v�����-��ݙ����'�e������$��O�n��p���\tlqL������w7�y�x�u�V��x����Q9��_���M�EGvA1��6�*T�4%;��3y{���A1\���Θ��=}wF9�FOBr�k��TdV˳$�Nǌ-��`����cE��i�h��>>�3[��w3춬ێT��ڮ�!���tͷ,�װX�����e���f�F|YCP}�2f���r�i��9��{K��cܿ[�uO�'!�Վ����j��eLf������}c:���OE�`�w�׺�ۖ�@��d�}���8��7��`��{P�� �2��ǽ[-�)8�d����˪�2���)�IC���z#�_7����\���#h\�)=���X���зWv3�yM&K�vR�C��cm���Y�'ݛs���/������w%�j��*ie@keT�U�tgh�U9U�m�^Gh���E{���kmd�ˣU�����6�h:�O�� w<�2a��1��\��@�^;����V��.���qM� ���,��,Pֳ��!N�i����^P.^�ڸ+��1h�. �np��{�ۃ�Z��ت^�L�����į<��F{��ϼ�\�q� �U��ZIe;ДT/`@��v$��}t���.�ޱٗVC�շ
��D+�)��0�+v�1B��� �؎)�O���X��x+����I�d='�i����:٣}H�֌�M��˝sx��ð������1C 묆D��j>?_e�շP_�r��w:���6m�d�*�K^U������;k�zn��A�����]���F�ydh��k�8{]H��mn�6��`݂��̢�W
����Y��x���Ӈ)~�����D�����Y[h�%7'�r�v�h��Я���J�W�����%i "����[�j]f�4@ut�W}E1p��X�g����U�M(��,�7���5��|G����'����3P[��%��@iYD�/��Y�*F��(Ѧ55�=�C��l���yn��I�ة���Z�v��Y����g"�U�e>l
���%�L�cpÒ��ЮR+ؕ(hVf����?p\V��갆�N�l��Ħ��CwoټV��b�N�aG�@�{޺���ܻ�k�'b��@]kB���r���E���W�\�F����D��=XL�����������O��<�*��rJ��r_�/U���n:=PK��d����n�u��7Y�u���m��;/e��ĊnM
PȺ���gu6.�\H�bWX�����:�1N�j��vq<��-�e<{�k��0݁4���s:�X`��W2�c��_<�F]��m���(Aj�;z�M�u��VU�����S;�a���O]S@�S����㣽
і���n8�z<��+7۷g�9U���,����Ņ���K9t��w�^��#�ۗܶ@k�q�W+{��9�L� ��]ɇ���G9Gt�)D��;v#�j}���/��[Sf.��s*�^*�1>Q�#�{w����j�z��P��������k�m��p���!o������p�o��x.�/��ʍG�����W�)}�������@\X}�^����K���`�	�]Vȫ#B�[�sN���v�"&ffllo0������@h���8�����4���?s����w��w��"D@��:�F�F��D�!UR�P�,� �E�T	!�(�D��"" !6�2dD(@�HQa.]QT�������"J�X��!&�&$DI	 � B!
�\�TTH�m0TX��H�H�	a����dDA QQD	�����AnY�&DJ\�*D����&�,�!E��A	�3 ��HA"$6�!A�� ��&M2��hA2��@D�R�������˂Ђ��E�D!"��JD�6�0�"��&h��
��F� � D!UR���%@��I�6�Dؓ
"D�"I �DHA"-)2L�m�$BAJ����ˤFګ1\�!H@�������Z@b��Q�u��X�Iħ��=�)w,�`�l6���If���^����0pg������W�We�}�+��o8�.�g�����C{\uo����ҙ�WS3+	iTj����;���&n��{�{������p�}'����˃�!���2O2x��2�T{��jL�Y4��.�����|b�7O�|��3\57��v�	]�8O��	h�M~g����86e�!�w��G���}�s�\s��8�8�.�6uWT{7�^��T�(���= �C�T��*b��w]9�P]�U�H^�ʉ�c{�Mq��_�:C=�g���g�c��x��Q'k�0���4%3�]��;������|�I�g�AO��b;�7x=�%�����۴�O�GX�<}��b�ϝ��Z�Xw�&�q��`�W[5̬�WpY�v��%�x}�CS�d����T�J���|-�Od���}�H&��@	�	S�)����Q�+`O�ZGӟ� �3��j>�N�>̿k��7L�o���sL�)�Q��d�"e*�cJew�Nq��up�Tk"G^��MM�s��{����L7>w̲s��n�u̳#�F��a+DLI��B�W3�D�{ޭ��=�f31Wd�9ZU���y\6�-u˦�-�.�N��;B�R�[^.�kв�B67��޺5lPknn툥�eÇ�"޻R�B��]p��%"�X�����e��D�܎��&�V��vS��Δ�'��ac�ᦛ�/6��y������υ�J�e�]l!�/���3���Ǡd+UQ�T��3���1͛�tv���kcz9�;C�<s2m�R���ŷ�t.T�l>�n0�t�vŏ7<2���cۼ�2'��TTNufEd�;~�ۅ��5=�<ګ�~N�Spݰ4�@YV1�iኚ��{s���}e�/�:OP>�a��J��Z^�Ұ��ˎ���bt�޼E1���kr�3�5r����,���+�>��>�:�NW����ZN�}�)�ܵp�b_Y;���_�ƭ�n�a�����_�ךn�gǃ>�dL��0�N��gs��������f�S�]��V�[��<�����Q�Cuc7ϯx���Xg�
�[����V����!u뮅�*��'�k�4��r�̏B���t��R����p��T鸲���9�{�C�v��\�����\\|eP�s,�����
��ݘ��y���0��N�1ޟV�7]�/HF�n�1��̚�.E8�D�jO"L?E|gJ�Qժ������9�{P�ɘ�=�0��t�a����Zr�j"�7v]�V��%�9|��}�&�`����8��#K���[;�9��7�[�v$[�<�w�� 鏨�|$1�ÆmHpM����۝�8ztw���/�-������ҵц���x�cI��Y\�i�kQ�C����k�-���],v�e���R�=���ER���[�ϰ9�>�=g}�+sF�7�$��㶳��ϑW�6� >�(	<���H���̯	���x{-�c94���/�����㏤�ۇ��r�uH±rQ��uA�)l��^�lewV��-F(��~v�u���N�h����7!��&�x�'MçQ5�F�8�	B1k�:eǱ��J*��&Dۭ�u��^��]�/�MZr�~������u�\?;�ʡ����)�?v_b��,�ΰdb#���F�W�}�p��֍F%���n��i�5�ԧ����#.Bgo�66�e� �]93P�I�_�Dq��[X*����oJө�C�m]��Ǿ�������_ �.�Y2[���q��ɯ�a�����)=��"+��+�ts�)o�m�gծUOOm���8��|c��S�~r���,�i~3�zY=C��e`WR��y��<f�#��W�����L����A?�.�1��O���s�������-{�>7��pf9����%m���~@��W�8e�8v��cj��z����ώb������=&�&�@�4��	�S��[Δ��%|�{��a^Г$o#�]Z�󇉾�X�c`J��ʴ�E5��8`+����Gr�L=��t#1��(T����W%RV���ɿ������n�����歏|���3��2��ñ��\e��x��<�v�{��:�u]SD�fc�j ��w�7S)�ތ4�䨎����U�>IV�6 ���V�ɓF��"n�nÎ���\�<0�g�v���W��T���/,��y����U��ȼn_}{+���M��q�]C1���^���nI;Q3��	�
�*e���Z�7]XG���]�*�ޗ�z��K�\k����9l����ރ>�Q�|g��jH:
�����g���S��Y�xX��g�*R&���q��b�S�4z5ä3�h������ϙ�b����=��:�+>�?NM��{s������2C���g��WP[�z(lKN�z9�4{Q÷u��R����u�n��C��:z����b�nÁ'6����^�3��_\U�}��>��q:���H��~ؔ�<����{TuI�-	�O�� �!
S���\^d@U��1q����#�s>�ٝ����Q��[��]jd�K@����#4�I\lԤo�ANxW��qѹ��L�>5�"�*����(�]m�U�M�y��X��ϸ��n��;¬�����ו��=�2�e9�v��+��>�E{�kY��a	C��w���|�Ber�IzW@�;S�J�t�����P%�;�z|
����۰�:�@�Z6�k\���چ�)�冡j���*�ɬ�+����Ӭ�Y>d�'�(�6����3���忋�~}�1����//=y?N��x���;�29�}wFN��ʁ��N��ڿB�u���j��/�i�\�x�GƆ�ǣ2�6���qM�i��C1UxpI;���)�� ��.5����J�Fx��S��K~خp�Mo¸�?��a���Z_f����r�l{��T�����:�p���X3sǽz-�v;��nl%�g0���9P�f�eB��S�u2��>��L��c�*�zJS�O	�=�K�ږF]86�ny��\�O���`��������:s��OFL��j�]#���}w��/�)p�[�<K�;ǓU�U��x�7i`��9>��.����_������qS3(�e)����9��`�)�
�t��|��3T�����7e��2���(�350��姺�ݴ���8�iua{��8t�z��z�p|��(+�����R����6�KF�������z���X�F��Z�Ϻu�]�ۼ�Kg<��{pݠ��'ӣ�w���C<���������r��Y���ڗ,�|i�)E�'�Q�:�خ�K9�5���&�rt՞Q;f\������o5�#������,��ۥ2���G����v�|��Q�z��E�.�]������:�;�|�zS��o���&�4~����c�L�q�I�j�6���\�o2�_=��Y�뚫	�����B"�m����l�� �rJ`%L)��V3����-�q���y�~��w���TwJD��yT�#<g��EW��F&[��b:_���9�Wu���gF.=Ւ�%����0��$S��&�q;pꙑJd�]S	F��O>�623'�}�\i�݇Ro5�<Ô�>�qϭ�=��Y�9�D�3Q�)Z���e��H_ego+Yb������ؓ���)�.+һf��L;�Z�7�T5�L��`c�n0
�?\����Y��՘�w��ݓ�����z������[;~�v�i����]�'@)�n�Z^���D��'�������?�z��,���鳓��N��Z^���Zn7/.;�rw|iח�\��<��CMܰ:Kj�[y�W�}��~>�:�N>�=�]KIӚS-�c��}��E1޹�������u�Q��[�y��Fl��Y�˪K��t1`�j���G���Z��\��J��^���_�w>�-uk��'Vf��rƕӎ����EP[q+b$�j-�K 7�7��/\�yk�efT�jgx9ۘ
����ʋ��'_
$���2�|�"��MQ������w1�'����)Ó%u�ZY�r��S��w����� 3�\1�
���9�o����6���4�<<dey��%FX�k�_����'i�NkM�� ��i^�i�
��
��M��<=�a���w�t�ƈZ�7��x6�i���2z�B�d9s(�s�����P�)YGR�Qn�}�|�y�u��j��޺|�T���a��HW(������B��/��ʀQZ��v�O2~�Zhι�Ϋ��u_v�qt�[?S�p�NW�l���`��2����I)K�%�V+9�駑u\r����e���9Y.���!���(�D<녾�>E_��ƣ�����'��������"M_�[{����~=[<)�)��x�q�}'�u�uH¸%� wTm�eR�u�xvP;OyI��r��'Z08�ՠ�!��n�o��r�'!(Լ��W�Oq����ڪb�ɉ�U�n"�_�F,]r<7�V��ˮ%��fp"m�ZvbQ����궹���Z�s.��&%�:7]+���Be}������m��GC��QF�/��cs1�2uU�&�2`U,Dwr�B��{U��*g�-�]U��]׽�]���^�6�f��ћ�0�Z�;��]2ĕvl%�������s�^����Nop��0��nڒ�������{#�����<o�v�U��3f�E��o��W�������f�O�[8+"�\�����7����"���Ͳ�mm�k�x��K�-9�L�����U
����50��O���I�>���g?"=2�E���y�;��VqW�5r���ro�� �yf�K�����]8[ά{\�4�2�lO���i;����7.�1���G���V|��O[��b׽S��c����מіԨٷ�V�N�]��V���歏B�w��'\��s��ѯk���H��mT,�]��ܮx=7��O�r����
�U��������N�X
�7' �CWO�r�V�~7S�e�{7��_������S�?�j�b�	��:����3�t�Ε���\at�m�<u/E!.�5yƨ���=�-�${��Vo�|&���D�t��%�Қ_�R� ������u?�S��=�⩃�!���7-��5p��}�����D��e �(ln!"5tc]yBp���5e��6�Պ���Ѯ����;pڸz�E��_qd�~��MXtg=���V��s�"&��SD͗N�^We59�3r6R��}�����d�:!ɱq�����=;7����x� �s�V�io���=q$|�]�ە�,>�"vpާrNWh��W%xک
<<�@��t�N�����𔦶6b��
ɤݬ��9��oD�U����G�s�|��nߴP-:��yM��p�ǝp8mR�Ep2v��Dחf�~]f�3��"ʃ0��I���Vd@U�k��o������Ndj߷�-��v�������2����2zk�)��䉔�A�+��
�8�b�Q���G�@��8g�nO��s�Yn��(��J��34�I\lԤl�S���\tn�����]�)g�MTni�ӊ�z��N_Ϝ�2_���M�EqGf���;���Q*u�����<<���N	��q�g�MY���/�N�;����'FO'.�@U���5�N��=0�<��l�!p��z��_l�$���G��W��V�\o;��_���A'UC��37,�װX�~���Yڝ~���F�u�[Օo��1����S�9�t�/�7���~�=Ω��bt��c���OE��8���9�.dv{݌JU���{�#֥���f�9�
����L�'�e3{���3/	�{����s}�q�q��m�A�Ǟ�}s�>��
ϋ�
}3�>��d��dʁ�DK
����z������C1��o�Tn��Q��x?!�g�BI�
68׺麕%c�<{
#XRtI�����h76��srZ
��]mn�X�۪�C#Ӌ��Z��d<���8���mʮWa���[E�}���FWF��h��[ʰ�В9e|/�S]��9�{�ڸ��W�p]���O��eW�gG]K����;-�����#�B���WK�2��.�7�2��:l�W��b"���:lYd��.1}�v��8EoToƙ4�D����(:��o�����V��`��8t�7-�QN�>�����8#��=O��0�oO�� ��21����u2��m����X�����8��{�Cۆ��a��ǂz/\�^=<D�ӱ���H�%Q�P'���N�C�+��f��ۊ-S�ߣ���q��yú���b�F��1�~��Lk�p��l����D�%,@�H�b����\TV�L
��%y�|M�S�#h�D����qiD�����=Q.��J��l�P�����y]v���~weƮ�7�)�F���s;��ͻ����3!Q�*���0��	q����*���cxr�z�r�)�w�
Xw��F_>��9}e�9�D�|�F@T�'��P��"��ꊳH1�)�>�e�b�=f*':���zZ�R��8��T��2^e�u�u>�[m��o����,���Ym�Ym����%��e��e��l��,�����%����m�Ym�[-�K-����d����-�K-����d�����l�[|��d�۬��,���[l�[�[m��o��m�Ym�9m�K-��e��e��e��,����m��o���%�������)���o� jVl�0(���1#�{�aP��*ف"�T��AH���I-��*�"!*��UJ��ȣf�R�U@Kl���Q@�%41DP���6�v�C��F�E�[lml[mcY�k��IS%m�ҪM6�a��"��,�3KR��V��*��٭K6_q��[�˱��e�dg�ܑI�5���K5������bnS�VbV�i�t��m�8Ih�j�l�*��*�SFl�kef���mQkj�fa����QA��YZ�����   ���h*u��io]�J]vۨ4+�=뗳J�]�k���U[mۂ������Q�T
+t�:�J�x�ND�	����Z�6R��jR�J��  =R�
<b��;�8.�T]:;Z���������G�E;���G�4��袊�4v�g �  �z�� ��=&��4Q�x�����Kle�m�3c� �P�B���@����l����F�()ج���Β���wd���]utj��N�]E���(�ř�k[�It��2�  |(H���\V�$-*�u2�mͰj�7N��_Mq�[CN�
v^�v�ءz��-�������:�G@���)�ڛu�F��;�+Lۯ�  �p�m>�Ê��Ժ�>�.̊{s�e[B]�;��2���[���#WkF����넺� �����(��f�Pm�[6@ͭ`�����;a��\�lZekkj��  ;u����ݻ,�R�ݰC�i�]Ѫ�޸]��ۧI��ޠ:uh��O:b;[��0WK3mC5�T�۶u9vꁛ�;MJ�0u��YV6�$��Vڤ����  ���w;�v�6�����}��U랴J�Mu�i銐*]����TѶ�q[aTm�W+���׻]�X��C���V4����H�M�M3��iE+Pص�ȫVZ|   ;�[�k�f�9N�R���盶�֫kH���4�]^���Uk
ݬ�B��[v�k��֚{f7��Ս�[8��tֶ����T(F���gv���XSmd�[3k�  z��GB^�2Ъh\�Ժ�)Z��u��� ��3MZ��;oN�ݭ���:�{��M�`�����=4)חt�׷GJ�=/1�4�Zت���F6Զ���  Ǫ�T����{^=�"�"����c�%�R����K�6�֕훺��N��ޔ�[`�lN8٪u1�z� ���q==�:i��S�i3*�� �OhaJQP�L��O������S�A)T�1�Oڄ�*�h&F@	4�1�R) ��/�����Ϗ��3��<��/�O�=#Br=p���)������	/Z��U}���W�}��Z���@�`�HH`IO��$ I?�B������w������������ӛk-�$gH�FjSt�A�k3�V ��}jĲY�3Q�I]��%�L�e�u����&��N�����F��q�M�E�
oZ�,�͍-y�c�oQYY���`�7_\�I����� 8ɜ]$*�c���MH_b� �F�"}��M�u�Vj�/#��6>ׂx��Y̗(T�;�],�L�#9(%#q�{��~�aNTF]Ёɝ�W��hAY�n��#��4��v����1����r<�1�N+B���;���@n�D�P�A'���+ 3#̧.�N�V�OV��נ̫l�I�jGs!6lսUX���z��Fhy�Q{Z�@f�/��8���L0ݱ���v��H4'��y�'i�V��b'�|�D�=Xn�:�Oj(�XI�y����9��f�������  ��f��W3k@X��Q\ :4��Ͳ�2v�"��9�@�%	H�f�����|q;����e���RG1+q�0�'�,nA�d2F��,��pf,dY�lThӠ7N)���V�B��GE���6���SWH[�˧��	����5֯Ew��Z������F(��iT�����wchVԙ�c�,�[�RA�j�n��S�n�dL
� Q� ��X��A�#F&�D�'(q��pe�o�rU���:z�4t	���JZ1�T�^f�T1��jl�i�7�^�t�4A��T:��]rڸs��8:��"�e�����*s3,bn����S��4d��^P�ze���e"Չ���"�i'�fL�7�������:�ePs���:}��[�0A��L`k*����4X��
ks1�
�&f;�*޴��
���G�Kn�m�@캊�T<CPNR��I��j�h8y�&A��ۜ]�Y��1�^-�`{q�FWl:����;g�܉���2KCjGN���K
b�:+.�(e�����U�2)�-�$�V���i���ɺ��Iђ�]݀�p96Pв����8���qɢէhݬ4��ܙ!�=���팈�u���H�F����B����<�tȵ�u��5����Ծ8A��QS���{RuD*Y˛y�{�NoV~��ڻ&v"4��`�&]�1v!շ�lj]�6��tļ��$t�M�k4*�m:�)mm�����/f����gh��cՕ����۷�{YvH�㋴��
�/7�����bsr��Ľ$܁M�aC͙xkd�6��"+=�n���[��]�!WL�oe#�hص�e�hZ��7D{m�� �wv�ëMN�46���rȷ�j��@l�	��W��&a��H����}��%�Y�Lq5�-(��G�D9޸5���ݷx��8�$F6��FȬ=#6��5CP��^��@�"�(o�0�JE�pc�f�*5w�$��4�[�5�
 �P٩M\�:hf��㡊jb�w��Iz!fuš��b�f�Ӆ?:cf�	�z�u2�Bm�WLK�r��f�k5�j\\�ݤɧ��*ل]��f&*�k��5=�+��&����-�ڞ�=ǎ�ѥ���%^���њ�+\��ճX�p0�̰�X71���Ju�]�AV���������,�恁�e�t�૧�tH��
�]�ZL�2̓dU��ɶ^�٤գOm^��3)+�b�M�7�B�ܺ��!o
2��[�p�&�ff��Xj��n�IF&��\�����;�����ϖ�9�N��m|��Ǖ?su�^��z�@!�Ko��	�f��ʃ��z�5K���S�x�蝫����������I���;�r���g��B�J�G����R`�,[�WC(:�Jl^,l�����9oH	#G��l�kHP�32fX�X�f�ip��DŹ��J&�$;������nY�/.�Mj:շ�x�e!R�R�23��y�9A�g5�`oڹ3�v813 ǷG���D,%��4.�/�I���=N�ճ����
���z�*U��;mr�i�Ʋ�����q�n��;�mJ+�����uv�	�<�cH�ڞ;tb��|���č�-A��cv���D�ۘ�#:p3m����M#vW0�!ݯ�.'F��~� �V����4��Il�N3��nSk4�6�����H�襷zv
��ͱp����w(�+6bRa�̷V��Ǧ�!�ؚ��Iʩv����7E�%dʶ��R�j�y����bR:5AX-�q�t�P�ˎv����*�޻�y@��H���mgؙŅgҵ��ڑ�>��'�נ�&��w8�e��vK��3E��~K6ۦ�p��,�A��W��8���'�v6�-Ԣyj�H��4��5&�y�M�T͉F�H��J�o:�]�G�[�L�I��v�3��_W�E��J]����(�&\�.����t�p�UMû���e
i�H��r�7Ej��8M�Z(M��;��]EK%����@�ͫ���*�v��Gq�J^8f�	��+r�J�TU�6� T��iStlT�t�]zś�'wU#6���97��9a�i�&����sG��Dj��H����Y�wt����Vm��1m�5�*��O!=m�T^���ytE�F��y���;����C]N���OvJT��ddm��emc��ͤ�*ʭ'p��E��
��:��ZHw"ȋtV��7t��:3v�Y�w:�����\��p׽��z�SNv�W"jYk���k)dw�L�$�݂�4�j�[T�XM$��R���NR�v
����X����5��8�K�Z��	&7,މ!5a�;�	i
5N��x��x+J;�w���A��.�u4Ay�A�N�C9p�;�@7p�B�Z�y�s��M�u�N�w��������V�j&���X�OX�,1 uoMyy|�W�a��2Xч���bWҌpAd
�Y�n��e�>�$���,�q	����x�G^����խ�0~�mL�c+)ѷ�tg"�[���J�^ޓ��	��L��T�Z�l�X����`�l�Wب�Pr<�F�2�'r�ѥx����v$5��p�v�SY���Wv�ǔ�Y�e�~��}����qd瓛�
��Dҩ��3\�e]�kr��mٕ�nobwM�9d����m�=w�]3d�nJɊ���4�GnP�KV	���Z����݆]=�3LΗ�wq�셗*�1:�n���H%s+�)"lJT>J�AR��PG6Ыw6�kR6�*������mS�yO
O*ECR�P�x����!�'3�P��Ip�&�;[��823�,^�~!�"V�r�j��v�5��p��`T\��,�0`7n<�n%f�{�lG�k+e]4�VRj�ۺk�[p��S�֥��W�i�N��
�`իCo;�=e`cF�z���Es�ǻ�D�1��Rs-�q��ٱ��7h��4�8wKUߤ��S/C��2��(�w1�C
��C�)�1,J���"Hp��(ժ��I�Rr�;�<�YM���1G�t��7��q�3&�z>�ͨ�N�:�L�7O�Z��QV�.��壜�j�od/Gdץ�����;N�O4a�����@�X/�13oP潧�Ը����X��*s�p.�a��:�]̱A������lC�r!�ͻ��)��Vod$�ت�h�Wۖ�ح�T>y��Jò��QWy*��ۋ&������i=!�2�w{\�-2Fc�qfң��
������3���#W��m��ʺ�Yt���@t��Fq 3V�p��.������ا�y(��R�y�!2����r�\Л���#��vt{�\���"mi7u����0 �d<�UIE����`#���R^��A-����Ή��k$�©�L��1]m�*P0�R��p��Bs����~,��6�\��W��n�����n�+*b��퓂���Vlnf�n�1I�ԅ"u���\%�R��Ј����~!7n4e�׷��S�ΔHX(�u��L��V͡���fՎ5Ak׊�[�#��rvnk�H���D�rS!啮���ν����L�Ӕ�W�O`>��ʬ�Z�HY���k�f���� �$5;�snpo�U����ݣ���/Jf��G�Ń��w��U�����w(�]�M�N�֡ۡq�3����c6��k �Pn]�'*۳t�7�s��-�\z�ًJD�	q�>2ۭ�a�(�Psܫ 
�B��I�Y��If�<�0�q��[�A�������P0KZ���Өo4�ƑB_6��� Op\+�v�#�M�5ģ˛���
��e$��1�n�&�	�@��8�7��Z�3v̰��i�e2M��f��ӧ%�4$�q��{Ǩg�P�Ո���A�po9휰=�jG���uq�)9���.��m���m<Y�X�P�v�fV3��ek;`���*��.a<��)�OM&��5��^�xl���wp6������٪ˣ��T%�W�D��')7��!�m��G7�A���G�n�-�6SG2�a71���K��8�Jڽ���7z�$K)��^���{^ �^���y�pC#|�<ֳ۬A6�h�o�cj�%���dB�C­n.�WV��ŗJ�	�n6�_bR�iT��r�[�!���ks$K�OV�@*����ǒ�������j��H�d�+�t�w�ũ��Au/݄ܶe��X���Bc1Kv��m"�BV�w��\	�qܻ^'�F仛i�j��-�Ry2+0+�OԸ�][ƍ�iIE����`<ӰņA؆+�e]#��\4��:YR(Om�-s�<�ꂵdXê�!��q�M�̻�;�)�{�@�U�ٽ�Դ�*�ZF�yZ�hGI���V.�������Y�E\��j�`�9^�{�=�ubI	������m����Ũ�sh���P²ΒX�N���8�ps�պWv˄󁌋��XEMZ��*�۸�!�(:��<ނ�����I�Қl��քj,�	goY��J��:��m+�UbYK���c�I�l��=�bZ���h��f�L-M�se�7�en6Un-N�l��-����F���tր�5�&1TG!�4ְiZ0���C>;hh|X�eef�Ȟkv>��f��*b�P�T6I���Gdt	��=�A=m�,��Uͮ��:-��yu�Q�3b	������Bx
��A�a-k�[y��=���q:Z��X�{eӔ|N�7\�j�vmh��^L̰0���o[Kl`&������#9����V��� iƬD@��y�:o�kQ�U�]��!�{[G��*�0-�ɐ���͜vǀ@MrB����D%��3�,�ٓn��e�H �4S����n;1�3�r��r�T�+b���vh]�dc���ӆ�jb�-��N|t(Q�CZlc&�-��ugNf���p��w�y�F�T7L�^���8�P�7"�^qVX7*����q�������"єZ�}������g�@f�Rv�e*���J�t7b�U�XE�$���'���C��u��idY��i�u!�qѢ@���ф����~3f��d��T�+km>ŀcS躬�Yz����Z�m�2����VA�F����#1D` ;�7ܮN�����A��	[�F��(Jܶ��܎��w�k7�&�V�n�"7���ɫ[��.��ɮ62���L[�Z��X��h[GZ�~��x�p�a�[��X�i:sY\ȵˣ��5�"���۵X�˶֊��Ӷ2�:���K��"	Z��IEԘ�Y�Jݽu��M��$IuZ�Y�YX\JD��D����H%m[�@�����Y��c�уwR�!R-����֞Tp&�:8�]�K�5�,G���Ҹ�� `M�E�y�P��û�E�����JܓH�H�pfAzq5^,A<�zZ1�l��Vm���a=���g�.ѻOr��igVM���L��WMᵨ�ZN�ҫ�\��ݑ>[�PX��R
�w���/T ���)���p�Efd
�N��2�`��4�е.Z�7{�r)G��v@��ࢁ������J�Y|��ݢM2���LID�K��PX�f�S-f"��wOn���WAr##�f�ے�,,yҡ����3�����ߤ�	�{NT:�m䳄�Y��p��'m�E�"�(q�cC�*�H�D��I��pSr.�.�(Ѱ~�=ZbW�N� K���c������4ź��ڱ%i;&��X�ܘ���C3��db�����̵�5������D(�NU�4�R H&�v�_2+v^eMI�V,[,:9�w:6!�J�S�"�I�2�b[���*�ւ��UǴ�.>ɡ!���s�=�Z���{�t�qL���/S��dt��7�� �a��o,�GJ�ׅgrs�֐�5��-����%��#�t�b�����7"�hf1;x=����uN�_5��9ɶ�6-���n]QD�n�כ-�9]�P�-����]��Pr�0�ފ��>��9���he���IM��lh�J��dn,��2��{��z�e����$�4�Z�fn"uvt3f�8�Y 3g�є��`���Y����[��v�.�v $�!P̻�E�θ������@(%<ט�[�ie�Ǥ<Kk(�4V�%_ܓ;���xaG'e��Ku�<|1+烖��Ǉ�3��q��Ovb�ru�̼w�G\�cKv��]!;�1m��X%8�9mpڄ�9��$fǛ�9u#)��8w�(������{�ӊ������-iE��í���$�0䗼��Uz�>�r0��o�t)��\E�J��=�z[�f���u��
�f7�QL���yu�wHt�kh�3=Ӥ�ڿ��ذ�<��m���������i>z�F�A!���NY�����:�[	х�;ݙ�Պ̤ߧ����U֬IE�zgr~�-y狷��?��f1�I
N�Vz���ƜW�Y<�I?oO�}׬p	�U-��]4�z���I����I��js�S%9ϩn���-���*Ƈ�d�u�wd��s�wW�%Äl�3U<:����`�`��01Z�!�^Q�'MT���7}I��eáV�*��g�3|�b�؛�ctq���M����!3$ֺ���"�v]j;`�nf�8M쩣�7]dۗ��;6擹\�a�mS{*���q �*�+5�d<��@��F��O���~��IH7*�XJ+�R�ɛ��Ш�C� �}�g���BU��¼�� p��7*�Q�_i�=&B�A��[j�}/���ߺ7W�o"�������޾�gX:�i��.�z�V�O:wm`�Y�#:`��օ�:&���GB�{�|Y[�x�̈e�!9���Q�u�s/j�3:k��q2<�*�u53FS�=%��L�cPWKU��dU�4*1O��e`��'��3!r�8-z���luvӺ�/2D�]�q�y��[p�/f��Wv�A`��"���2����7�	���빺�^^"�2�w;�㏓W*>������Ӆ��-nk�]r�73(����Dչ)��?,z�e;�#��}��u�E ��[��t�w.�Q�}[�^P3+��H;�� qǝ��'��XUW�f�~����*)/�x�ޞ��Lܖ�A�N�8˷��z@�]p��Ə�f�E�^�탚��筍W�f�Zr`#��Ehgl<�4��3+���5��{��,�e�vo6
�����S�e�Gt��b��vS��t8l�I���j��ʪ�U�HzY��I���M״�p9�;}��+�{��k;�ϝ���/�.�7s&So�!G-T��T�x�!m��䳨�cV�6�%T
9Z귯34��0���YYC)�$�Б�)���9�둃����Wb()����h��YW�n�",�[m�Z�"��j����X��"O�͞O�i��[�\�]B�x��F|=xz�BDo���g*=�����2C�3���#��NX��a̛�چ���G'�t�¼{�U�#�!�m��렒��r�w�+�A��vu)��� F*A5+'��oJ�ϽOMC�^GC�h#�*�w��x��lfϞ
��p��7�g7�hdV�j[&FJ-�,��o<�º�����Oe�c#$=�f���;�wr;��$oit�
u�Zh'w!���e���Uy����rgO��Ԓǯٺ�4Ƽ3p�������|�}|�?1�Y�{7x�и�w"��r�m5�~4��d�Ɇ�>��=ˊ�	�y}�q"��o��.�ݍ%�)�r����i��Z�cĬ��A��b:������ѽ'�O�i�񩴘�ࡊV;%�P��釳voM�e�,)��oa7���̸����1Kj{�[w��:����ۭәu���յ�7�a�Z�&�G���"J�DƳؤu6��ڤ<)]�Hv���(d��1���*�|��o��r�V�Pw�zqx{�x�ǵoZ���3���6���Y���^K��9ێCwM�Y�d��,;��K���g�Z�E46����H9l+��B�=#w�b����`m �k��.�����Jjj!��*El���kŊ�a��er�QQ١���Wb[�˭Ү	��Ļ@AHwD8o>rD��y�W��#T�k�YTU2�a�d��7l
ݚ钅�Z�P��.�4���V�_-� �F�ݠ�)2�ü\�Z�X��eL��\w/c�5Q���������!(c>�8fz���ח�+;5E�RY0��;j��n��b���W-�e:���Y�f3��sٱKv����p��Q���ǜ�oT�̾�d�2�a�lT�:^�n;�F�� 2�9a�lY����겜����!�j�������xO]N�q{~�b��Ϭ�B�ܨwn���{���Y�*��{��̭��r]oke�6sZW��;T�J^ô�p���Β��N�ȃ'��>,��-xWN�$ژ����'���_^{���'[f���+��FO�X�p��$'��޷�*���=�|�j^��0�7�u%'4ե�	� ��e�'$�vD����#'l;����{n�E&�q��FF�{D}��u}���n�P�޼iϭ	\�ڧ��0�q1bq��)�Z�uc�{�䉨��i9%�a��TWR��e�˼�
�����)��bҩڳ�i��#해�Cff������0�-�e�f�Փ�2�'�\�NÇ6��&�ϖž7�7���|*��x��}����F���ӆ �칻��j�}>��R3�C����B�SY2Pz�P�ֳ��M⧜h�8훐dT��cU�����gV.�!����JH�R�i͡Mj�
����=P�������������ʹaSj��VI����}Ƨ<�q�Fb��ٻ�&c���E�4���1��v˚�Y6�V.&�3h��n��kK�tMM�F�F�q����3��� �7`����c=;���>�J6O�T�6���}C/J�ɕ1����Zhٗ�^Զ���$�,њ��է��$y�js�A�w2R��I�D��zK��9{�;�F<��:]`������~ߘs;la���厝��}[ȱ2u��Z�̔�I�s|8�D���&��$��3F�<3���t=cy�_��<����ëu�I��;_t��J�O��{�����[��=�z܂ו��F��>�o/(�]�$����%�䮴�a�����G1.5u(%�9
�x�!�y�gjܖxʀnS
���6�E>�)&�J�k`Ɋ��Yw�M㊓���pY��T����}��t�4�4җ��[J�V��g*X�z�\��GR���L�.���)�yL������m��(���v��#O�sm��4�WY�~�s5K�H���N��u7����|�V�;�cz�a���	=&��V�^%��!��U�s�@.���gnY�r�ge��N�Nj�	3����#/!E镒�=�x���MG�iȫ$��h���B�$�%.��um����3W�H �X��ĕ_c�qˢc�!g��{��+���nL���=�7�7�?;�>y��wy�I��bH��9
'��t��KDV�u�W�f`Xb�f�
��vq>�NN�	�M���ۢ,�uUo`�N�%g@����"�o�WWM�'Y-�83xp4>`Ωh�ob����2�0wS�&͔��(�Y�Z�v)e��yV�:���%���.;�H�V�qM���x3>�n̫�wG�d��Zfŵ��`<�'(h�������t�7�we(8��	L�Qzh��Ş�O�Qb�x�%Xw���X�S�րM������Ѵ�6�Z�!�y�d/�3n��⹞��rx��{C�&\�&�[�z2���=�nS�w5JN���2T3��C���o�����6��9`x\[<���E�n�����&�B#�8y�L�1�6t�sEՉ�M,r�
Y��ݎ,�IY�̍�̴oA���aj�}�*)�K�@2������W���9���Sr<�"��X��Ȍ�β?v���W��,ۅ���1�mk�!�.#����W�Qf9�=�w9-�C^>�B{��4ŭ����N�\K�;5�G�ũ3�Q�]d������S��n�k
�I���{�R�tfeZAR�bw��78ΣC4Q�b��h�Y�ʃܬZ�L�4��h};�<S�d�/!m���y���0QR�KM�o�W�cC)((�y<��˺�9���gJ�6M3��nO����	�N{\;��;6s'����!(��5�v��"�
��7X�=,��77���7ʻ8�u�E��w����=s)��n�6�L���h�����z{_�\Y��%C����{�	���1�u_u9.�hZ�Q�K4��*��jV��1n]���N˂����&e����҇c];�L�y��B �Oo��<u}�E*
�f,��X�q�$�X��j:��N�f�0�ꙮf�Y��H,س1T�)��{J�%+���֪�0O_3sJ�e����iOs�a�I�9���u�&r�,��m�)	BV����Џ��}��z/�~Kn���^�h�7$�E���=� ��إ�A��+�X��Z�$v��ݱIU��.�b���꒸�̔�^�o���'����]���5��ZB�`0��i�E�-ޚh�i�:{|ڇ�=���p�X�T�0���-�8���NCL�[ր�]���E
�@�s�6'�b�H��`a�X�n������tfSD�w�2JoN�ޫia);5��7���1:;��̄=���l��М��0j�gAv�V�w^����GA�n����Ó�Î�5<�覣�oom�ʊ�ō(*=�-\
�	r3�h0�U�J�ͭ��9�5,CP�h��~u�m<�S��h�=7t��^R�m}�%ƅ�֤EJ��|��w��k�*�tX�wr�J�qs�F��}Q�ꥳ��w��JkN^$�L���T���
i��$��t��]!�+ƈ��tش����]"�&$N��'AǕhnV}z�#�@]�L>`��3\�L�SY�f�5d�ޔ�IK^�w)h������n'c�_eA*$k0F��,˦�ݩf�l�-��t�,C<�8<�h���ձ�bxS��A�9mѮ��ȷ<�V��s���r���'�+���0>q��"Q �C����S�.7�0=����s���kF��UN�ϲ���Ŋ���\����<���êKI�V6��uN�5��l�'����Z�!W6�u#ھ�s*������@R�'%��B��^�S��鼌L[/r��	�+��n�EH!�3���>�)�����49Kr�֖C[s�&��R�EZ��VS�r$��W�w��Ŝ��ޅj�m t��+��g��39=CO��]���ZA^���:m��=z����j��Z�d�%�n�'�3'V�E
۶l")R�b�+:�*��ލּ�g���C�
��3��}����֊�%@�8��\��T<r���^��(�_8F��WK>]{�k*�syf5�$mK|�_�H����ѢSBW�v&�nh�{؟�'g��縅K��7��}C�]�jR��3l�Ov8�tT�$�|�ŝ��<��%�W]ӓ�R��7��4}%�\�Q�gF��7��nyzｬMz3q|�o����J�0m���ۮ��ZNY����$�mZ#�+J�d�g*͘��5&��[����w/��W6w����BB�t�n���
�/�[Z$��=^:n�k�4⃨]+۔]f� ��s�y��⦈-[Ձ;���b�%N�z^��0��a��ɨ�����:I|�Cz�����s��߇�3;}�y9냸	��4�T������|��L���5�t����^��xW�>�+͌I����2(R{Sm�\�sN�J;Q����R\/@ǻk�V�w���	��3B�qsgK�Lʱvf@�`���]�F�]Xk�B�@���Z�e�o#4����/�S`�����Ro9mXw��&7u�T�*_>Ot'wZ{n�}��M�k5�&[��V9�W#�[����!��o�G���4�
	�a�a4a�5U�[ĞP �=�ŹN�g�2P��zjڽ�Vv�3ik�9�mK�C�DŔ�3<_QO�-�����c{���p��A���|���j��kvУ,�{��C�g��ou���U��N�UQR+�i��W>9.��������d� s���D��h�Wڽtx��eZV� \��/�\[l>	��s��ƹ�u`6U+��Hq�ε(F�>hڜ��Ϝ����p�ٝ�e�$3��i��D�f�kN;������u����e�b�{]~�켑7���\Mj<֗��F�:k7�M_qi��:�~���^~t=�-��YS\{DQɒ�*'uj;d�u;V�)��.%�m<MtC�:j��
��l�f8��l��i�Sz?
uO��ʥ��6��c�7�4�;Wğ�dD��W���-	���K�=��݅��K)#yPS�hAy&;vi�m�@���Z�D�bWm��[�u�����3��M���oskY�b!��v  �'�k�E��T���M�{&oF�N��K7�#�8��#�;��u8Vw�����lR�F��ھ�.�c��hv��OV�����0? ��|!P�ksfv!vʹ�4��+�2�niu��],��Cg^F��鴱SM;���������|��	|�����=֥j�Et�p#o�[�]٢��a��;�NɆ�|#�t�[�j��h���Yx;fi�\�!��o1�Wr�Ε^�M����ݾ>�!���Oj��*ZS��/��83�J]W�G����[�9R��u;������F�/��q�o�N��S��t�����4�vc��y��ő&	�Y����|<��.��EF{�/>sì�o�[�B�(:�`�Yݲ�0d)ɩ�α�V�Τف�t`�}�r�[�!����! ����IN���_�;�35��L��J�q�ހdU�MjV4��7�m�r�4��'=D2OOB�q�m��D���{{f��K�%R�aD���W�q��a4�Lǝ� ������Ɯ>�=��O<���ɝ�od/ X��M����f��OS�� )d��o��X�
�S^����={+ u�%Y5����8ֺD౿DY��*�(��2��Ն�6Җ.@�����ҍ�5{"�YH�r�Wޭ��N���&_� Qܨ��,>��c��u�}>k�tV�����%�u�:2�2b�k+wlW��r��Ǔ�\�`B�:Μ�Q��;�y�J���c[%���e��KQR������eX�mlf���)ìG�nS�M�S�j�3���!з��J�.>���d�H�ǔ��@��$�(�eZ�%S[�#��i��I�4>�yKI'[eS�k.��4/c|��]m\��<mi�,4���#�f��9�]{���NJ�GeN��0���/f=��ʜ"哢������+��Z���
Tʺg��7��3��T٦��a��K܇-�鳜��\��ڛM�݇8�}4�}`t(mK�/c���f<�Knb<��<��^j8��zP6�Q��y��l2�		52>MbY3C����TJp�i:�ܣi������l��Vr������'n.+��&,�L-e���wIfޝ|��Ԝ�u��"N��Ө�Ƽ(�.<�HC���jS�%�3�c��Kc;HΑ}� Mh���ܣS��I��\��w Uݯ�\���������O+��5�Y��m��2[�b�,�����ӳz͗W�s-��77;kb֙a��f��+�ʺ�Zfa�c����1�7��â
��|�ڵ�B��]؟��k %w0E!�R��S���9m�*����w.�Hv����=���O�%K۶Y|�Qn!�[�8[�$ݑ"|���������+B,��i�i$�wZt��khP~Y=g=�}Q��U��-İf��C|�aO7�V'V���[�be��#|'��tiT湡]�z\��>��'�"�u��3�7C�,�*)n[3����4���{,�n��u@D� 6��#��t��D�P���˸f7fao%�c�:�7}�;���ԏn�oL�Z�7˔*�֞箵�Wr�Q�dd��Va5ئVT�}��/c���hB�3�����a["QcY��TR���Q�$��X�]���j��s��7�K��P�������������Eb�.����hW^
�t1b��J^��Z.� ���j��U�]x���{�׾�����y�=D�����OyA�@���V4���(���j�Ӳx�^�5j�k��������UOQ�Ev-�-�^�js>�x1NI4�Fi�"��~�����4AF�^C^]aCXޡ���A���µ����f��K�rj��n���I���G�hB�{���PgJf��{-g�<mp�_g-���n�4����+nwYv��+;w�+$�0�
�M}����<��%����f���h�YQ0Mxq�z�˃Q�w����9�{�	E�[}v����� �ƭ������d.�IÓ�6�0ɍ ��s��w������p��ۃ;�M���ɘL!�=��^	lcKw����kx� �ﻒNFD�����P@�8��*�o��
w9��2��NI����3�/�ڷ۽]R�!2�s����2�@�潦տ�f9(��+g'�r�4.s���n�9��8��a��Oʽ�;g�C+<�6]�ZVrEhV�\�����x��"�缺��ʍ�@�y-�`��Y��O��'#աг)��x�Z���ҭ�m7-u��v�),;�o�c[�)	浦ۍ�D��E�<�O?'&ueW!��ȝ��k]8n�!]AKqbYc�J��Wr,i>��24��(�K�3�\�R(��K'�cˮ!d��©�=���Y��V:�'+������@>�R� L��e���@V��������#������+��B�[ݾ����k�d�V,3�dMv�Ȁ@�q��u����Q���ky�4�YD�ٜ���jʽ��T���h"׳Y��q��J���x�]���18��3���26�ס�T`V�q�-$r�ZVXy\�dW?�|�T�ŵX�B��x����b>:k�/�g��{�	�W�-�ut����Q��|oS8�gt+��Bۡcrc����5�j.A^R���/c���b�h\F��}x�����
c�t�7�@g�L �kN��Vp�����vm�{��{د�����ô��e�|��ʧ���3��ٕ��� u�L�q�(�戲!�����8�Kx�o�j�򺤺�u��u�5����{�+�����}��ҜceKi:�Z ��=Z6��K9��",V,x�Os���M��қ�d��'N�ؽf۷�(�:�`�����/�V}��H0=��z"y�x\���t,V���/,�+�<�+o���;ۖ]]�tQO�����%�C�:˶����yW\�#�s-��5(�u1�f�:y���ܦ��L�Y�2�,�����F������Q����#�Zx�"��k���g�}�����,M]��"C;|z�]�2���@p�Ls��F\�<��6�ov��
�ia�:��H�5A��a�%���� �c)]D���	�6�aɇ2SU%[��mj����qtO5��s�}��Q�]sOӰV=@�S.��m���]nk	�'���C��ND���H]�݊wa�����W�R�ƹ�Tu��_�����l̼n��	��&ͥt5ev���F�x�!���R%Q���yu��&�Z��΢�:���w�'հѺ���D�׺:dj�e���GzIFn��e��lY���Β��Ecy�܆�j�T�?^�2(�Ku�����r-�U���WQ�t�Y�M�g9���N[�O�0W�7�k�1Re՗�Ak46���]XZetao��uo���O<>��������520�Q��l���)��1����ՖT6��ʹ�ȗ�h�e���t��+CDWKw�;Ώ�>i#Ȫj3r�^�$��ݏV� ���"~*���1^Q��!54��tK�G/^��LRf^69 ���b�3YJ�ֽ�b��|n�������su^�HZ�7Ɩ�c�^�'SBF��Z&n�Xt���S�ޙ�;��cUz�J�`�/�vI�m��"S����]Y�T8�P\�u7z(�{+�(6�t���2��{o�׉m���N;��O���Ӑ���y]��f�b#{�=�Z��'�V�XW(L.�|�+2Yk;�W;jV�F�r�\®f��c�p�q���Sv�d������K��wH�r�����m���2�p����\<x�+qe��	�ʋ;�=Bk�y�����K�s�Q���_E�M�N.��˾ج7�m�iz�����s�.�SӖ����.�*.��~�������-��p� B��۹S��T��{�"��u=�@�6� ���Op�ښ�*q��,')��Y�s�b8�21�O�o�c�"(�s(,q:I'�l���TQ� 9%���V�ŤU�^B��%�g</����Zm�2��z�Ȫ��$�h�4`;��=�6Z�2cB��t�!��`J�q�wHrn��V���x�Z'�&��':
j�
����R�4sK��DS�6���U�I���m|*�j	F�ea�j��\��>5�7Fwƍ,<BQfq����O���۰-����n�� r�����|�*Y5٨�8�77l�̼���حVj��Z@��4�ۿ�Cwo.f�L�*�A��dsCA��Um�#��-m����@�n�&P�n��Y�������4i3�^�,��闪�v�`�I�)�A�wȩV
}7}_�������F-lxb�Zߐ�WN��{V���ĲnxIMkO��.��6</�^�c˷]E��z�j�*���j�Y�9���Q���@��e&��ښ��K�L��7k��<yW���1��8ﾗ{��t���P�"6��k�"FՁ����7m0����J���TAǫtZQ3��Rap4g��N��ж�xe ?Lꐆ�i���p}�y�u�HSK�_=�R�B��f�`�q��F+%���I_V��/p���D<��ƊC�]ASݔ�WJ���<j����կC���ʸ�˘� �WfH+P����d��鐫�J����;�O�WS;�Բظ�^�ՌF�I\����c��oapZ�!��A��aN;&�:����w�L㻪�ɧ�NEnJu�3z�掙m\�D1(�8��tn�����3��$֬�'��O,�v����:2;xq_���|�'�����xp7���7���k �@��l�����1���v��^�E�����j�:'v�&�aVr�{h�6�N�K1���b5>fy9���	�����y2%���(�~x�3��P��ո�l��,��q�o� U�}��V-�u�ԡ�m�,��6�`����|�<g���s:{'K�x����n�$1����)�y�*Tr�ve�yN)%�!���\yvh�H�Җd���
������2d���܀���;Ut�3��S�I����n;��B�ie�Kݍr�g�t���M��4�\���Ww�ޓb��u�
rt�$�0��S6s��c�n� ���f>=�8j��U�oI@��m�[kƴ��Y�j]���>���	��%�/%t���n�����+��Y�˂^.�q<3��7&{��9�S�/�z��£='n�]Hm����F�DM���j��ݗ���ᔔ%���4ge8R�X)�
MWS���o6̺�75�I �C�uu#�{�>��lB�&z0jQk����˸�~J�S�w�W��dٻ��Sլ��N���*�L�Pδ�����ɀˤwB�ˊ�>�^�o ���I�Y\~eu���W�1ܪ�v't�9.�`��q��7���abΣ��LS��_dd�\��SL�|���lW�����f����2M0yNWV��!JOzn��X��c���g�ʼVFtIQ� h�t"�mu��VM锕"��u�z���u�3����%�Bx�D}��ۙ�u��	�3�v
�?/ 0,.��H�2߽ra�}�%����߶��:pH�Y��!� �ZN�hWXo�����Vm��J��חԪᳩkӥd�ωw)��Q�r��\!�\�kك��{�C��K\|+iE�
U-Ֆ�x�J���vx�b}P�$�1Q�������<yd�Rz��Z�`4v�QNI��W1�[��X�=6���:�t�U����{�	���H������K1�N�r�(;n�Z�c�S�R�T! ����ə[�9HWk 
����d��!���|�\�
ʂ�<v��֭�TGsS3:ܞwD����[�R��J��F,t�67���*��t�J��[Շ�
�J^M&�{�]�<n=o��z�	�r�;Hek7�T��*����ha_gZ�7�(
66}}h��;��̌�9L䕕�zǹ�V!����x�8�C� [�Rx�j�/�N�c�C-�_f��|���öݾ=<�{pk�_C�wf�7��X�	.:vL��	w �,�Vu�|�]�Y3z���݉��s,���kz?���K2��MՀ��ɭ�����C2o�����tX2�s|��A<\i�d6L��I}�ُ�k�z���g�H���[�V{��y#�Z`�{�l���ZQ	F���ܗ�i���[�C��Q��;�[]�\,���RѺT4Y�*�y����^_,r�9Z���+�S�u$��%�U&��1����,��w����aX�g �3==p���}�m,|L�g��"���ig�․�^� b�-u�G�,�h"z-�k��UCP�ɕ;#���KR(JxȽΧ����ٹ0#��3(��997j���V\yi�t4�:,�#s�M^�/�[Ҫ�j�~v(������˚��ū.fԓ)��ۻ6Ta�c_B���-��j�����k6�!L]���V��3���v隐�X���:U����JE|����>���wF� ��A6�{&ʻ�-_[���1�q��Vgp
N���9���r��[��A��^}�\�1�0e�v�5��~�,Ql������VѨ~��O/�c��Cf���sw�S�-�QmB9��B�8�C�Y�H���'�SS�WM﷮���ʑ��D>r-/�=!�����C�޾K�aj:��[]��vt���i�ܭ��0Lt
�F���n���-�P�P���K�*��YBepZ�0G�znv[P]�I�n���%�k�.�݇2ޜ6/�=�H�KT�,���L����F��A�T;I��ck��~�-|�Ż%m��h�j�tpQWqj��2�]v��{)Uޙ���M�!�NY����E�E�VV��:��uhA�s�WWI�D����׋�KVsڳ$��*�91���{W2�Su�	�Q�y}z]�i�U�PT��<t�Z��1��n��W�U�6��S��G&���I7�6b�ϯB�1���S�:��xfa��y�L��.	ل��J���K��x�^�}}*�v�DZ�v�V��F��yO;��X��5�/��ң{�m;��ݵY��rMGG+��^�&L-,�-G�{,k��
S�j �M��3��r�BM�Xn�(2Z*�TJ��j�������SV���Y#N�K���	�Ô4��ˣ����+s���9�F��ʪ��������\�ʻ�� �������Ơ��}�(�bf����ۼ.�)��<����B��C�n��y�J���z?2�.�NK�^�h*߶���M>�.L �j
��ˮ󛻦�Ѓc�tz��� �$�3GQD��z)�.U݊�S���z�]$vi�rV��^� \�v�F]�X�u���9�K��B�'�e�3k@��/>N�ǯ�鍷l?p�F{W��'�𨂉�������hn����v(�6�W��zSL�ErP��'&i�?=��v�"���.�:̠K:��#�V]Ԯ�[��/1�uܸ/��% |6m�3��z��g��[�qV��M��L��U0�wtu���n�:ي\aՈ1V�Q�8�w߻M0�ԶB�L�z��v��5�5)�56�p�\�8��o2��WK䮢�Uz_h�l1a���˾�,������gg�u�I:*:aX����+{UG�ܩ>�s��>���O"ct���y�砪������r�uԪ��X��!�4v��B��Y�8#K٠W�U:�!�������,8��˙9�Auhx�l^
s�L�I�1�t��Yz���kw�ݠ��fP/j-?��d%���T	��I��_�
�+.�����o8VS��<��y(nd��˸�Y�7����ĳ\A�y��*�u��=�m�O}|�Y57t{5\G(�S�sղE=������q�(�E
�R���X"UA��h�J(,��%T�E�6�$D�
"T��YU�FE�ZU-�lm����iR�m�*[�*�RAH�j�j���E�*
(�RT����ԔTU�����-��V��*�
	iiUVV(,Ym���ek"��Tam*ڌX��Tm-�V�%j(��+iR�DTDch�U�b����EHR�`TQdP�j�DH�TdZʬkej4�FJ-jUj�Բ�*�,�U�����F�
ږ��PDd�QkV�-�����)[�EA��VQ"��5���X���Q��VJ���j�U�X+h#R�R(T�UX�A-����R#E%�U���҈1��V*RЩY*F�ATPbT����+aX��T�YE��,+TXQ��F��laR����KE��ciiaPDPb���6�KjQT[eF�PF�
V���m�[QX,�Ab±�������7��鼸%`3^�B+f#Z,e>GS����)���[�<u�� p���mٹ����1W����<�5�9�|GB�f���Ն3yL7�����&t�[��A%��s-bA3}���3��uη�ʀ� o�g���\��]Dz�G³�JU��FI���*O��嗮�t�i�n�+��y��������h�
8��-�F5K�Peӡ�*���c�ny{5� ����eë)''���;M�
�訞����Pt�ޓWe9Y'�xS>ìr���=؀�TXBZD5αZ��\/�<I=/ų������'5�TF�6�<��Sw��O�uۡ�p��+������APs��	�>��:��<=�My�s���2����s����:�8�;�sU�y��	^Ş:M����c��q�����cҽ���vޯ#ho���=#ROOl�"&�l�.^*D�{�����w7L�" ����k=c��dM��"�K��W����=�Bqjbg��`���mD+��o���[�f��_*%ۏS�,wv��gQ�G��4�VjJ�-�r�1���2�T�^���y>���u&{zn�h�����t��x��<M7���/��j����ᳰR�+�������$�`����7K��2ovEA_S<��g�$<�.mJ��^]��3N�woLGh�{ǲ
,��0�$%Z���)���T{�^L��F����|�3�_"�E�[��b��a�DA�p.�ON�U�}j?�'o��z�[9�Q���^,�6�	d{�xHr���Wb�rM���z��V}�{��h~�qz��x����~�9���S�!u��Ҩ���}@�p�MƐ}�
���Ӧ��1Ǟ�v��[~]�pA���<��UO.g�}B��@�.�L��z�g*ox�*���9�yG�M�O)�hg-߹L�3��Ւfp^�y<82�6hP�O��n��Ϥ;��7���4'Ued��sك��Qk#����^f��70��#&(4��7gG�wn��/N�k�W܀�( k%��zYIS�x)�Xg#���/!��R|`mª��wNެ}�{��W��������c�u�B+ah��5>[l!����܄9��(���l�EF���N���fnc���՟8�Ъc~�ѳ�Z��+�|�6��%��{w�������g���k�N�\�UV�J��EN���'�,iU�����*�xi�yT���~n�gl� ��A�?����T8�||��B'��~��ˮ;���h���I�5|���|�s~�uj�vj��jg{Sr��`A�O�x�k�Z�/;/��� I�}��j%����[�]v��#��-�ı�G''G����b��`�.jx���Y�Ǉ�U�`}栻�{r	��/k�H�!�A�N�Q]^�M齮k���h��P,+�
�2�%:\� p���=���x�G|8l�{�yv����y�M�X�>��Ϯ�e�ZUb�+�]��[�Z��V�����m.�*V����%����
�?<%u�aބ����'g�R�u�w��5�%��=e��z�[��误���;�4�fk�LW�ւ���/n�&r���LQ}�� ,,�ll������K<W��51����]{K�sJ�,�x���DV�n/z���y6(��vtzy)Č�.���Dy2�_tƲ�j7�F!G�	����k_r�nG�ǜ}�'�oC�m3梚a��Yӑ=z��yࡧf"G��B_����\������Ш��tOC诬�馦�T�Pkږ��*����d��8��-�w����[�c}��������p����3�g�)���-f�v�ļ�g�����$���,��lr��>
ۋ�^��Z��1ܫ�Vt��*�-�L��
�s˟8� �OM+n ���0u�|=F�C��u{�3���$F�{��"��olaK��u��^*�6�8-�)�u�V��g���p�4���2��a��~�0L��E���%]�]e
cn��g� �{7�vl��Șaw*+���#�zu9y�mW��B����މ�Q� O��'��TH5�_�k��dz���7;�c96 ���(8`yP��eIdV�T��ĩ�w�^ӡ�1�۳������q��>�IV����z���aϻ� ��0�� < t�<�yj���n�SOX�
>����h��Y�V͢����*�{Uc>���3�;�AZԠG�h��@Q�[��"e�z\t��Rմ���0��K�#��[D��~Տ��T�W�bP�nd�t3���7�����<��m��n��
�{D�C��cC�����p?rR�-�+T���}���{xJq��p�%�D�p@7�o�����n���6Z蕏C)r�\��b;�ֿkyg�/����"W�a��'U����gWa��f<����P0W'y����9n�=ܦjזp��к���$c�r�T���S�ܛloы�9U�4�t��jns/]5o�ީ���Ʃe��Z�5�L�k|�a-�_6-踆�2B}l�	�3i���jӊ֏��O��L���ޗ���p�Bv�k�*�~s;=�z8ەyxCf�c�JZ�3C��f�7�7x�\�Cfr�&=U�i[��8�2�n���������
� ����n��t8Re���&�DG<�D����k��`{�Q�O����K��3�W>^�6��ؒ��='	3z)w/��ܪݷ����M,�[+�'(��+x:ڡ�
��]m}���6xftǘO�}����;|׫�}�U���ɜ���أ����<��{����<�[�u����ϣ��6�O!�^�;$��%��.T�vУZ�=:���{b��N�z���.>�^w]��>v��m�T�uK�F�
�V����㬃���G��ީ����/7�yHj����LE&Gu���ɨ/1��=�]�I7#���g*�N��GT�.�����wu�!R'N81�^�Z��j-��o����v=�ڵ�y��<�1��qu�$����F��_=�oY�&}��6�F�O:����Y�^��c]����*�����e�!��%E���YB�����wX��6)��F��ǹFq�P{	�Nˋ�,���v�+O� �i����Vm�|�I+gz��=k�@�J���=~�9�극�`t&-Ͱ�q�m�jJ.����[��Ů�u�¡��[����r�/85�%��wgB6f�6�I�Q�����^���b��䖯v�1�;�!�^�#N�/6�]�;����ϓ��_��V}��'���z^��$v%�9�M��7᫘����Fwsr=k^�,��'݀��{\\���q��S\��)����U}�_���*'�gԕ綁ɴ��f�%.�l'�/��1�<# uz�Q��/p��߯4��^>TP���}mQ;���u�� _O	;mf���^�X��Y��c8�q�#������m����ʵ��U���[`� ��ia�魞�q|��åL�$�U8>U�v6�WAO]9~��,��v=�S����}��?eC�=�F���-is�D'��?o	K�V�W�՜V9�L��ӝ����w.~3����kq��R.���S�k����M�5}�)=-,q˯�v���l-|��H盖��K��WZ��=޵X��u��\����2Me�Y�l����%x�J+X��i�2�C]b�Qۦxʹr�Qq+%�5_��)��rr�&��.V���S��mr���w0/��|&��&����=�^(�/���5(����j�#l��8���v\�5�<\�m���Iv�#�7�Reߔ�yC�y��e"�Ӣ��Q�����˸ٯvQf����3c,�O���M�S.*x�c�����-O[�i}��t_�u���թA�&��?V�J��յ]�����kHh:"*rC��Ozl6�k��g}M��(�P��Rcѝ+�^W9�[Y���Cc�	w�Bʓu�ۋ�Oq��=���ުRP�ړ�麫sf�����̇{J}�m��>`���_V)vj��-�++{~�=�����>K0�@��ڇl>.�=��ʭ�>U��r!<<����w�Jϯ\T\X�wA�wL�����7�Ҿ��s��۞Ȃ��m|}q��m��f篎Q���s�\��\�K�G_|ć�zy3Za��u5y,�h��Zf�7��w�fd
�~.۽������~�N��k�ׄ��P�T|3���#A �ʱ[��-k�V`|�]�HN�;t$R�
o^V0{7ub��6�\��:k��=��Z�7��W�ʴQ�H��ae	�]:�����	{HGv�l&�ځvE�nicNh�Six��Mv�=J^^wt*
f�콚�j���-t�;���ײKڈI�%�<��UI�2p�Q�cP�˞��Ѱ�}Ǒ^��-]�z��ߨ��x�䇠3�ם��T������K������O<g=���b�C���F���j�ߏ@afg����u�ۛ*c�Y�,Ǿ�-R��ES�
�}Ɯ���j����T��v���b�����E�ܩý���J�\R��S�hc�Q�֪���{2�n������3}]���j8�� ��'��-�k���ZD��q�nn���ۗ���GM*�v ܎�=늶����]�2������Wy5�w������s1y=��fg���9Bێ�T��UҼ񙂰vI���^}�{��N�c_\�*��=�S)�ѮPߺz_����ē=ftOۙ��+�]��}�3fQ�%E�X��yG��u��>�J�}A��3O�и3����������~w��/��i9���x��ps^T�_e�L({b�J���z^��fbS�Kk]�F[�p�a��ȷ/UXt�\<Uc8o2	ݯ+H�R�	�_�(�Q��Ә~��ĞMz(}|k�J0����:�B�;�!�=����!Ũ��4��&$g��|�M�:����j;����=�rN�ɽ�o���h6�'���K��ėUCg	��C�/����jZ�* vV3��y�7u>��OoA�z����W��9��ʊ����s2]���㝍���J/E�GP����~p9�3'��8{USO|��������о�N��b�X�0lGm�'Y�ܛ��SDy6s;�Rʨs�;��"�c�h>�dxMŹ}閲�ߪ�l`s�����_=���ex՘|�x���/C��{=<��yv��ܓ$e�*�]
��VZ��Nk��С�^��^�KΧwA����M�����ϔ�.Vˤەf�K^��7�Q~e�=Vc�^l���;�_!��_��<��͹��"�ɑ*�Mإ�p'�_Z�(>~:��[���3.}z�$-VW��oN�v��m�Oy�J���ו����v�b�\��ZĔo7�~��I�74VlwW�5�`7��X�T�n7�Z鸾Y�VU�W6��8�V+E<l3WWs�3���Q,��ށ�1�^�J��7��ֺ�Q���'V��V��_L�v*ħ&�ѹw�ۼ��ȳ�yz�ҭ�"�2<��)�W:�ny�}�d���~UO �]]�f����{CM�w7�3�ye��]�K��鱶r�[7꒎}7&���*���T�eWw{�mo��X;)h��O�{r�O�-�	��)1�ϺW���`���~3<��>�WN��J]�G���Oғ����OW(�/|LW�<��^ߏ�}C���<Z���o)�iԡC���]v���"����=�)�7}�{��y���f�[2\��J�����㚃���u�-�����qQqfk�rk�����P��B�w3#��bR�
���T}|'|��	)Uw�a=q:;��<��4����uv�s�s��^tE����Un�����rZ�L�A�A�v�j�[�8���~��Ϝ���Jc�Ս�Q:����@��=�~��׍*-�י���Ohɕz��q�[ќ@ej���ֲ�:;���Ɔ���=�|��Cp����
t���/��}��A9o��VSu�fЬ�&���d�f�S�p<t�}�J��qi+8��:Ky�KN;Q����][�(ͭm�@��Fst-9��ݲ�=��pw�2�zP&.������?=\R��et7n}b�����at0nY�ӑ�h�(yὒ:g�"V����0'�u���-�0
�'~��M�H�m�]r�������m�<�XsP.+�r����)�M"�����\Ō�d�X��F�Zfձ��m��/�Kx.��l��s�b�������ԣTC�.��8�����l��vYr��J�~U�������xy�4 ┚v�p��G�d��>��=��#�뭲7������*.�Փ���U+��:��Ӛ+�I�j�"�l�:�c�]B^��:n�8 �:��E��;�����u�V�o1Du�AC+4������u����e���y/��<u(��Mam�|���X�&Ћ��x�.Pt	T�b�U�G���M��&���/,l
�m�a��dLmҋ�r�R�7��I�֊Ǫi�nEg
�,Ii~����W�|��Z��]Q�Iwq~�9�'\��X����YW�r�m^^��Z��)u�]僜�{|�7���[�1:n�:{����9�ڛC��;jQ<�/�֮V�@%'��ڴ*]z�҈=1{r}��j�#����Q=r秆�S�"�}�+wS�s��wJ��^lW%��L� ����3_+���eL#4��ö�Ǧ�����m;!���|���t�8�9�f,�R��Q�F&9�]�j��J�C�BLo)�e�ڤ�7C���Fҕ例ʣ}L<�(=���Ľ��7\Q�Cp�٧)e�m3qܚ/s��Vu�RQ^Ѻ�z��I��0]��L��x��k~��&��ze�T � �m�u�Sb�3c�ct�0V�Y:����V��� ��ш��\އ%k�5��֜�
���h�VkY��G��b����M�ǐb��V�������H���h�x��n\�ˤ����m2�T��D�ͺ�ڄ�ü$�7W�&�(��gۘ�V��wu��2U���z��	��u:wٶ�(]51c9�S�=�=�;0DS�4Vᰵ�d^�ݍŬ	4N�s���f���k!b��S��:4=z��_I��k�v<4���؝��EK+w$�S�c創��:��ZYm�+H]u�YtfJ��m*vȳfM\㶩�k0�k�-��^���ni�;ټL{9���9J��ŭ�s}rZÃ��v�ε��rpڳ,��1���Ńh��ؼ���R��sk��(�ͻ��5��<^�9����ؔ��}�>��"2T�����T��T���m$Y*UH�*)(��
D`��A�+AJ6�)X(�T��R���`(X��*V�m�h�`�ڬ���F$�BF�)-�(-�*DAk
��cĪ��UH������@���c+%��T��*J�X,X�[*�eeK(#[ljF��J���QeE�VV��V��Qj[
�%BT�����XV
IQ�E*U��*Ĩ�TKK��U ��h-�P�Y��mV,+i-�E�bJʅ���Z4��J�TX�%�
����ҵ
�*+-�B�eB��Z�eFځQEU
�J����AB�����@�RU@��Łm�m%Kh�
�RV�m���Z�����Y+kT�[+-h�)��aYid
����j�eI��/ε������$=W�ET{�.���"��>Х�Rf(�l�Ν�:�^M�S��0�yĄ�>ɛV9N{6�5	��rI�O�����I�L틤�8>Q���������o��{��r4�;�S�=@g���7�ߞG�iL��+��*�NIyE~w��w�ﭩt��~��ˠ<��_I�������j-�:i�6m��s�f�hϱ
��.p�������L�k�z_A�[�Y╰n��':x�.e�$��U��v���8Ys�}oo}�<{\�r���}c6/j���4p���������q|�Z�b��Z�{����2�x���,r��;�^����9
�:U {K�z�j�5[S�}��>3*ݺ�vzN����ȷ&l�\w@.����&=ҽ�3>�ԃG���깾.�4��OLo��o�.�U�3���Q�Y�>�UZ�q�x>����z{��S��'�؂ޔs�Q��߻5I弥g׹q{)�c��@#�L�\�Sn�rj �H�!�<�x�Y߅�$��u
��
E�ͱ����V�H�e�*��j�=N���z��P1��u����H}[��
7G]��-Z[8�����`J�3;_S���ͦdz�[�w��ݨ��ձ�2������n�Ej?���|��y�ۢ���}y+~e{�ا��w�8�xzl\yL5���=��U��o]u-�+wA��ճ�2�,��\�ݶ;��_���s�ן�B]v�h��'a���n,���zߗ��K�4O��~�2��������m��f���Օ�g�5=ͭ.{2�[���]����wO&�{˞��!��/��\~z\]��O�W��毯�u����9�T�~k��W�͋��WS!^�Qq���o{�ˆ��n]��Yn{hS��/�@af�yߢ*ל#�a]�;a֎�)�5�S&�;��<�Q�/�Z~}�b �,l��h�m�{��ŹREו2(��u��Y~�=^|ӵ����o��6'��z��gW%�ޒ������\��T���:�e���ұWy�^��V0���2��}�ᶊ�7���D\�)�I�q�&�El��W��+������y �79C���D��j�;�����U]b
Y�e�L�י�+ěIDjhݭ��:�ˈ��5��=���)�Gvu�F�0�;Ҧ2s�~�g��W���ҚU� �nGu� {I���n��E���{�t��}��j�J��Y��}ދv��Jn:U z���جʱ��������^W��Um{9}o<�;����[�1�е��k25=�$D�=�-��ܿ#�\��V��`���m��G�K~嚺��j�� =Ç����q�}\�������m��m{C;�o+}/��n�/�9��.M�{�8�9=��{��U�@实w<g�;]�&�o��W�������ظ��G��'�q�t_��{n:,�z���\O�y�#����ʊ3Տ�G;�kK{�C�m�U���D���(|����EΌI��b�m|H�u�o:�;����TP�:#���ewv6S�'����l7ʽ*Iޣ�6]{u��=�ź�Umo���ܥUk��px7O$���?��2 T0�^pg��F�ܬ�B�>;w��<��s	T��:��dE����at�os'���˭A5�ڼ0��ة��떽g�H��w
��(��]���1&�-�����bL�^�r�a͜�r�=nԴ.Ћ��5�9��_}���;|=�=ֲ�ofS����v(��]qQ���w`�Z��M��շx�)���:����wzt�=�)&^T�I�wN�o_>�8��3�s1�O'Q�j��ꞓr��ח��&w���&E?|Ю����x?^�N�R�P���jf�Y�&b�V��ǟKQ�CorH���)�t3}��D�(�cu=�۱_?_�>LG6?}O����RdpL\�m�MLק�X]�W4�����u߱���~�r|�q�Y8�o�?$�6ox����^n����#�W�t~���sL~�5�c����O�&'}�2q��d*d�Vo�AI�'��0��8����W�I�YN�`|e2OS��x��C��j���_X��+��	iG?_����䖳[�����L�C[�a>aPPY%OyN�q�����'i�w� �����}�I�O7�I_Y'<��O_�;u�>��_|m_ݏ@�	���F��Q���8�~�8�̛a���Y��/��|�P�)��5�a�N%Bxw�$�M2��;�4ɦO&��$�B���������������߹��p�M��{׽���'��,>a:�g��<I�'�p�<d�O�d�C��A}?k	=C�y9̝O'����'�<��8��Mj��9�4ɦO���ϻs�~�������OT��yA�lA��k����)�ϫ���⺣ڒ/پ�b�^��u~hrJ�=Ƙ�M��v+�8�lI�Q��$�w�,�7!����qA��t2���yM� ol�;�l^������-�Ҍ�rq_������x�J��߷�������&���&���!�u����8�>J��P�N�?M��̜Ad�o�Hq��Y��`N$��u?2O���Y8���=��o�_��u�o7|ם?2x�����w$�$��<�+'�ۤ�R~I�xB|��:�e�a6§�q�k�C��Ad״�'m�������o���s�����N99��__~>��=a��̛}a;�a��L����&�N>g�%a�C���+'Xq�'�N'�)��Hu<�8��m?���'R�3�}�g���7�w�Z5��}%Iğ2����L9�q�I�fN���N2};�$�:d��'M���IRi!������R~-��:����`��UA[��ǿ~�����n��nFˏ/}���i�|�}���J���>@�'uC��$+'X~�m�N�x�ӽ�x��O{�!8Ͳw��d�O��$�4��TO�*���
�>��s�?���]�=�6o�r�|��w$�N'�,8��'_7���~d9hz��N�C}�@�I��杲z��'���x�Ԟ<�$�~d�}_~R�o�'\�jR˵���%{o_o����=fЬ�Aa�@�N��<m'S�ya�d�g����N�d=9�0��CygY>a9��l�0����u��1�!�A64�R�����V�����'O}�Y'P��J����IY:���m'm�XN2i?y��\I8�}��
퓬=�0�$��=;�'��?W�~~��~+2�T�����a/�+��@�5��<d�{�0'P������N!��d�+	��8²m+'��Y7��O���M}a���'��AW�>������y���#����`��#�Xw�a�2M�r����4���T1��js�!�4��}��$�O9�IR��j�d���Y8ɦN����!�>'��W�\+�Z4I��^ ��qJ� qgQow6���w��];dH;x@e66N�l�'EH�>ch<�j�F��8n^����k���fDj��P-��$��=^��������ssA�V�Zk�$ˮ�YN�vI.+�9Y�N,x����UUP�����F?��}d�'�F��Ğ0�ZβJ��9N��	����&�R;܅C��Ag�}�
O�~9�O�'o�%��8�4k�>��𪭐~���fs�Z�W��67~޷��'�''f�:ɦC��=~d��R}7���x��=�󬒥a��a�I_��N��
C��Ĝd�+M�"��_<��>���Lo��-��;/={�����[���m]�u<2�l�������N2��������5�>g��b���'�u���Ad�?{�:�Ĭ�{C�d�+���������?{���wy�>@�&��I6��J���M'L���$�C�&����q���p�x�ԝI���6���A���z�GՕ%��X>��O? 9��� ^�ގh?o_t���VC�_`|Ì�t���d�'��_�>`x}I�Y?2q+	��?3�e�d�%Ou�O���?$�
���4�Y:�|���7{������xoZ󰘓�:f���$������'5a='u�:ɷI><�@�	��}�+'���M���!�C�~d�Vq�|��>�*���{����Dߦ�Z��m��P�&�P=݅I�M%f��6��w9�Y�	���:����w8��v����''ϙ�IY:��7CIY?$���>�����޺�����ȑ�?~S\g�OP��?P�
I�|ʇ8��῰��Y8��>��~�2wvI��0�'�m��l���y�q���������}_�?���q'ӫA�ܛ��^k���x��t�CH~d�y�ē�u�~����6�,8�Ĭ}IXu���w��
��?�'ua?2y�`v��'4�']$��������w�󹭛��u�VI���쒰�!��l*N ��-!�:���2��m'��6��&��Y9��3�N2u��w�	�.�}�`������tW��~�5D��A�'vY<.i���Ҭ֭#��Twx6o�Қuc^{WK�K�jt��\�b��7ɴ4$�\�}ĳ���,�M�0v��#)����昞j�􁛝]�F�51>Ǜ�U� >t�,�[��2�t��l��M���}�����|��]7Y��V�_�;�����}_~�����{���I���J���Y�*N �Y6���O�,�i8���6��'��d��C��`|��;a�s�w8����7�^��&�N�y�v��'�9哩�Ox��	�~d��I�?s̒��3Vm
�Ԭ����d�y0��J����;?}�/�!�
��d���Žp?2m�M!����I��=�����0�}��:�� {��O6���(N���G}�RN!��d�*I��IY6��/��SW���!8fi�ʄi��w��߽$���:}�尜a�;�]2x����l��P�S�N�Nl���'i��{�X~I�x��d�w���+�S.�#�>��.��~����3�[ۘ��I������+'��*O>d��;?XN00׸?2u��}���'�5�䒲��s'Xu�s��?2q!���*I¨�~�����}���m�ՙ�U/��y��o�����OY&�w^�++	��'=�N i������q��=���OY8��`|�d��:�VT>�b�*|s�u��)Mz=��wo;�_w�{��밨x��T<ՐXz�Ӟa������/�I�5�,�>��y�Ì�����񓌇��p��d��}���'Xz;�>��UT=~��q7O��?G�|�����g���N%By�d�'4���H,=d�����u��~��	�y���O̰�$��x{CĜa=��"}�}PW۵�"�߿~�������}���� �������s�u���՝I�VC}�'�8ɭY>���M�y�sL���}I�Y4�ԨM�2~J�2OYn��al=�6���^��}[W���`8��6����`Ci:���Xi:��O̓�o�u&�Y�M�q��䝞s ��i�9�IY>`~���~~���00�@�G󿶥m\�A����ΐ��I�,~鼸��`���y��L�������6'�umb�dg5�8<�F��/��:�I�ط�3��h�W�5��S��0,��7�}Eb\�m0e�w�$��LA72J�J+�z�rw7Hw������_U}U���\߽�}����=O=O�(q$�*~�ìY&k�l�Ad�`C��J��	�a�9�S��=7�:�Ϭ'{N2u�O�8y�I�I���k���g5��w[7���k}%d���P������Y��'�m��?ya��^48�ԩ��B��'���d'u���:�u���:�߬'�u7��^_���;��g��N�d���u�m��0�&���|�������Xa�'�e�I�:�~��	����q'X�B��'~���d�d������;��{�y��o5�k���I��0�d�O{��']2y�2�i����J�IŰ�+'X~����N3ɗM��y�é��m�����P�����!�߷������8ɦM?3�\�
��?w�ӶN�x���p;d�'����q6���0�$�?s�IX���m
���i!�N����m���=��g>ߝ���~��y�{ߗ^��4�i���C����{;�2q�o�st�&�N��I�'���;��:����,&��&�{��'�s�IPP��Ь�Jɬ�;������������?}���@�=d�;��|Ì�:�I��d��C�s2O]�������{ïRz�h�d�~d�ɹ�rC�<I�}�Y'��M���k�o߹���o]��{�oz�d�(N�_T�eI�eI:�������&���Xq�q<���N���ē�s���Y'=�����4���:��4��4��<���u���<��Ͼo΄�I��ԝ9�IR�����&�Y?e'4�����a8����x铬�a�R�O�sZ���Xy�Ru$���|7��}�5�\�5��~޽�M2~b�׶�|���su2y;��'Xy9�IR���,������d�'����d�!����I�'Z��W����P���4��罯����d]��P��.�X�W��d�G@�xw3+�}ɏF�v<��W�p�����%13Xe��v��Bn�Dc]��B�X�,A/,>eR{%�D�-L#�v*
�5�����stk�ځ��Q{�}��f}�*y�i�ϝ��Y%J��y�4��&'����N �<;܅C��J�ɾ�'̟���'xoܒ��NjȲw���I��xn��N2꽽���s~��ߛ�׻�O�8�I;�d'��C��:�i�C�s��J��y�Y8�����'i�w� �����ϿI:��rJ�>������G�~v��9��?n�iv��a�����T<a���|�4é>�k |�2u����:��N�����k�q*�߲|��4ʇ�;�4ɦMyt�u��7�}�-���}�u�����w��8��&ӦXO]�x�e��O����:�ߔ���8�=�|�Y:����$���s�:�2O��S��J��߳�d֩<��}��o�׼ݿ{�`|ɦN�{�I��0<����ɤ����O��u�|����ԝB~߹P���O7�I�8�Ԭ���'u�߅A��X�c�ۮ�.O������~�|�0�7�8��M��l�d��3̒�x��7I������O�:�e�a6§��Ad���u��a*N$�*9�yͿ���������k�Ğ�왬>�q���:���Ӻ�l'Ι=?{�m$�Y+2
2�u�ٖC�����)��Hu<�C�,&��k��7�Vg�X�w.���:�*���(���k�T�I�T�d�d���a�i'Xzs2u��2q���ܒ|铿��a6�����!������R~-��:�Ƣ�_U�sd}��%x}��^�����̓�ÿ�8�Ĭ�������w���?w�6�'Y<I�{�6�'�����N3l��!Y&��?d�&�߾�yvy���������^��ʅd��ö���8�I��O���i��m���2q���9�2q��P����O�=�;d���Ny@�Ğ$����'�M�ŏ������b���Ds�Y3{�P��α	� �v�{���G�!�ub�Z�~����8��}o��h�i6Ņ�Ri�o����;&��'>v"��+re�N?H���.�upL{JjG�ҥ�e�:e�r�9�Co�7{U��s�&�ImA��=����;[��$	 ���s����=��
�c�߰�	���+&�X~����I�xaI6���ya�d�g�p6��L����O]!��:ɦ�s:��`k�=�}��ܟ�G�y{߫�`��R�_}�'g}�Y'P�s�%ABf�VN�d�ei8�l���q�I��d:�I�y9�C�+�N��;�:�4�y�>y�<O�ܗ�þ�Tv��������4��M {�a:�6Ş��u�<��d�C�s̒�a0�8²m+'�)8��M����'4��}��Ru��{����O��~����{�{�dI>a�[Ì%f�y;�=a�Iδ�N$�S��T?2i�s�!�4���p��:��{�T�&�0��|@�,�d�'S7|~�J�Lg�~��b���n���kϺ�OY8��w�Ğ0֯Y%J�\�a�ý��N �<�r2i�o�AI�N~�N$�߹%��8�}�}�e�-�<�����ϟ��"���d��~v�5a�N��������I�oyL�ow���a�)�I^�:��)���N2i+��Rz������M��?z8�d1����������s��φ�_�8�a�I��y=�񓌇�}���'�8��5�>g��b�9�$���\è,����a�N%d?x�_S}��_<��\�5��4��O��iL�k�~�m���rJ��L�Or�z���xC�&�����a7�>O̝Iԟ��i̝A��~$����o^g?~��'��6��=�n6��l��|�W��u+!�߰>a�M:I��d�m��~��'��|�Ld�h�	��<eg'�S���	�I�y�7��X�2=�X����&w[��
�}��~�'q9�Y�I����sV��2u�n�~��	��rJ���6�La�+!�1����q�|�:J������-�L��3ˏv.�\QǏ���&nv�G��j�{�b٫T��pUc��
b+�Ut�F�7��t�n6f
<�v'G6�mw6t-��u�ؤ�*]�};�!�ˣ]����n�2�2��B�1��^����6�
���r�������-�pn4�p��ӻ��F�c�_MT�f}�kw����kV�)�E=M�lR<�µ��n<RVu6�9��=�K�{�E�׈1�}�o��,v���ow��Bm���򆚕���{�+��ع�o>Ut:ᱮ;�$�&,Z�!1��r�|ŝ��*�����
�( ���&�K�,�kT�ß.���^�J0�xm4�U����J'��͖�ŗ<�!���Ÿ���e 3`��G�#;o	Z^�ˤp�[�����K�U9�x=�g�5��=L1�y{�V��!3�+ϱEV��F��nν�݁5Ӭ�ۚ�spBܕy�cT�c�L����.�;�9�qɵ���S�u35+��s3v��bh"ͤ�nZ�V���xczh馥�W5�V�}��&E���X'P�u��S�6�9v�;E1[9+f3g�7Y+SיCgh�
�gK
�����|�Z:�G+X��/cv��knm>�K�mǵ�ҭ��]�BT��˂�W�o+;�΢3#��k��!w�ȍ]$��l/<i��L�ұ���ʐgo���bNf��%�8���7�x�嵍@q��[ۍ���o�W.4R���d.��V4��F�z�v\=3�i��V{�$�X�X���{��+,�0�����kmr��^[�7M������a&���EV���g�*�g��8��9�ݳ�ُ7�@[�g�u�i������jnN�ŊZ�(�>��Q�?l�]����!9�|���b��cd@g��=�U4
	��j�2y>��!�b���ۦ��yY�odZ,�~��ѩ}��=�r��M�󯨞�׃@p��
�\޳������&G{o�w�ov�!��F�қְ��;QνZ �s�j(G�Hw��a(n�
�7�fT��v��鶍n�
`N�U�/v��}ۃ�jy���OFH�4���W;��B��x�
]ͧ�I��n�):uŬݴ��(X��^����U����9c)7cI���ʙ:�G����.��kj�G��Ey��K��=���x��n_=b�Ch�}�l:�_&L�a����EG΢|�5G���G������CF�a��2U4�9N�͠7��h�?�#�:�y5e��A1<赾���q�|�E&'K2�d2(;)ot��7��U���xӳa�u�v+��1�$w��J�/d�뙢���d�ƹ��R�S�֘	���Wo[9a���>m*EV{�o�+�W��4O�ͅ/�IcZH[�Ld�߫00��ǎo��趵˛z��3���A���,^VÒ�=	+5�1���h��i�rWf��z�kn�V�P.�+����4� ��PVAIZ�j�-b�a*�Ȥ��VX�d���
1AJ�����@�ёH���ŀ���j�)h%d�
�JȡZ��
���AJ�ȉX�X,*�AeH����
E�XAI
�!R�YB
EB�U��V��
� ��EDE���V�l[FҌT%d�%@P�P+"�*�ʋ����X-IQeE��ee`
RQX��X*�E�Ȱ�+m��
AE`(J��)�Q`,Y+
��)-�mem!\`���TdF*�E-�FV�eD����V,���=˲���|���HŰ��K���8!�x8�oz�0�N���u`\��1��������#��Ȭ��y8�=��H���s���y��[���$���ʇRm�XT�d�Vs�i:�s�u�0�a��a�N?0��;�@�;d�ϲN2O�3̒�u��t4���N3�ws�����Ǻy��<��������~�I�g���RLיP�'�<��JÌ�J�}HT������'Xz�:���d��$��'?Y6�m�s�f�<9�kϼq��;������}������VM$�<2���8�e1$�f!��I���2q+Ú�Vd���Y!Y:��{�����<;�N�=d}Ϫ���z���gG-�������˯��O��?d���֛aRu��i!�N�J�m'����I�ya�N{d5������~C��$*G�?s�������}���.�߸h��}��zL����J�u���t�YUn~�Nk���tk���w���j��_�wD����t��|��>�&,����wM
?o,��i��W>�ǧ�
:ڑ����$rW�=~�<�Z�e3�I^TȕL�4�8Ww�O+�=Z�L�);��}��S����$���ϥ�򡷹����b�J���ؔpf�=	��c^�>���v"�l���'Jw�@%7#Ϫt��j�AW��V\�2gV��ו�eN����3sٞ��ǡm{��]ឫ���������D����\���{oF���m���<ʃ���3�2�çح���J��KSq���Ѿ���7z�	@u�5�#W�Uߒ�����z����ʓM����6���t���qݼ��;4����#]�ŕ�MM�R�Y�w.�#2ez��o�UUU_}G���ݱ��_�f⽒�T����iQ�	��̯���G}����%6.�\��D�;h]g6��t����U]���E�X�l��'��s:&�Omw�ɴ�>�ț���0�����|�r��f�6��A�]���h"{9v����ܽ��D�;�ꙫ�*��Qޜ\Y��
zy#[]�^��?����^�th����/��Q�Pn�{\W�/���q���vóV"y^:���NŹ�B��p����8]'F�x69���@���Dh2�y��]�N{�y5�QCn��k�����W+�����=|���v�\�]�R�^��ݏD�ۧcn���'�����o��hN����\y��J�{�}8K�f�Qo'k���[��P�<%������q�{�3���+�o_*�'���>��F�{�,�$ˋ�i�l�u��g�}0�>���aI&��W�m�: ���#5�:VC�%onC�Q�e<����J�����ˉ/{ \��F���R���_�����ϔ��_�#p?7�]t���:��q����$˛�&;0�[j��y^3%�=������,�quz��MtP��
u������7�#�Y����F��np��{���g�ח��gyH��dG��j?e�����w]�ј���.�.u�{y��f���<���A�z�[Yzp��;�{��pU;NSژ��j�53r$u5T�=�%��qVw�ٗ/��7�q#��:�si��<_�]�E����f��ʱ�S;�Y%�w�I5w�����'J@�*�^�jڮ��j/|Z���ZX*X^���;"����/3���Z��UU�ҽ��?Qώ�m>����
���!���|M�Օ]�d5Z����T�y|�1=��i�������:��y=�*��y�Q�%Fz*��z��u׸����{ܥ���Z��K�+$�v�>���)��i����Gb��);u��/��Ӟ��D���q�1�7���<��)<,Z����E�N��BJ8������{���i��zJ�O�L��׺��緹����{�v%8��wұa�*��y.;M�4E���r�A�X���疔�u59�c^�nGʸ������}�N@N���up�7��ŏ]��Z�v�;�cW��Pr@�?[��u֡R{"��?}_UW�}�;��=���zF���������U�5�Cn�xF���'e��[=D�}n���/s�����M	�5���ߪp��|,{~��t�����d{=� �ɞב��'�p�;bꓞNz!�4�{k��zI�ھ���+�ԡ�ƹ�=�<tϜ���y��)�x���g`p�R��g��{�b��>�ޣ].�p}�<�iuO<�5~4�JOO�KY����Ϻl<�ׅb�T�jL�J_��ED��C-�v�Ȝ��^��I�����nT�udSʦS�hZ���Z�����L:�d��ڳ�L}}���y�JsET6�>�^�rj�qS�k�����n���9���߷�뗓/˶T�� ��*D�@�[�J��Vǫ�K�m�(��7�r�yS�{k��]�z�[��_��m�R'�4lO���,W�k������)���P���ʹ`ѕ��sO��9��D�����ӹ[�[�D���N��z϶��W�7��<5Q9�7y�%{9r�gx�W9p�C�.�{x�rh�/s�˸Ȟ�^Xf¹��L$�W�$�Bi.Q*?�}_}_}��+ӱ��~����qT��i{�N;�3����vWF}������gkbs�{�1��/��W!)r����/N{��-��j{���z4�1�9z�8��sZZ���	�z7��&�h^ۆ��cI�o�������V�����Ez�n��z�.,�q�Ms�� �8[G�8u��1���_�?ti�Z�ȕX��}K��=s��g��9�x�Jޟ�������J���ɿ�	\��Y��~�2����i�,��p����E�np����i�TN�Ur�}��z$��%<�|��`��<�mΝ&�k9-��ܚ��X��U__q��1w�{�$)�9���fj��e�w�k&]'r����sX�ɘ���D�y�~��4�������sJ(ғ9*��݊U� �ϙ��U׷�Q-@5�r���t���OG7�V%[��:DU���,U�+��L�����Wv�ٺj|��})��Պ�(�FjDar���Y2��M���Z����_�'�Ʒ�n���'�N���r�����fܢ�	��1:=������i=��l��\ʻ�Ϧv��*��<�kݕLŲK��*�M� ��^��g�g��;��7��L܋)si�[�y̖���l�����ݶ�D�ܜ����3�;��a���"�'|�O�_�j^�UR{Ӿ��N��&���9��M����s�0y�ߒ�vP���_wq�[^��w��!"�������!��A���cվ�U�{X}u�sǝ��*��8�X�+!��5?u��y6�g��B��(]c������v��U�N{-��Om��u�����5���ܝ����R���M��/|LH�S��>^�&ן���y�6��-q��#z���C��R��R���Qޝ�g8ª�sv߽��R����{�S�z�����${��J5�GK���3��ϫ�~��w�����9��l��e��E	����8y:5�8w�aS�^".��A�7u�$�F���z����Jy�8������Gf4�A��K���	�M�QZ�C	w��B|�~��{d�k�ٶPKs�خ2��.k��_����7��v���M�>=�$ˏy�f��Z"d��j�_L�qd
��Q��磌��~ng��3���S�T�g�.b����5G��v+�ݍ���y/i��B����2�{��-4�����k*e��r��^�nh��.����H����ҫ�8*��7�8K��T����Uۧb��tZ7Qm�Pmx4
�5�����U
S6dbNU���'���$�ʙɠ��O�����}ϳ���m��*��zEF�]npo�{����ywI���H��4�2h�Y����i]���R��k0��V����_z�=���f�{OgR�7���؋8�Q=u�OEQ�cG�����}��SR�{Ӣ6���7�D���C'ٸ�)�t�@�����@I��e�}q��"��N�9�}��lי]���B�N��k�zڷ�'���7F)�7A�{�%���=�j��c��뎻��r��8�D�7�z��gy�����L;k^�<���|l�B��8�s8������M[s���� ��4��wX���S�����^�{���Wx�����~d���Z��\��l��'��Z�>Cآ�3ð{,�
�x�Y��Uv��r|):�tW{�f����U���W�S�������zOo����Getgڧ��E�{�b�W���N}���z��Λ�|_�f�sem��8�l��)^{�>Y<���F��1�u�����F�n����MC�7�B����/�%2��� �]�`�����^�>��rr.��vܘ,_}�-�눾�d�7J�ǽ�NZ�g��g�����)�=�{ە��宫7�䣹�vm�J�O�،י�z�Ll'�@�xKnt�g7�=���@X,�	얤����t*���"�wʺ�羓}8K�glY���p��v�Ne?�q�j؟�T<U�v[�n���+��]|��?1�gN�y��	�-Z��r����igZ�+��%�~���{B����ϟ?)}��
-{���.z�I��w�ұ�gz���&rj��u�,��F��չ�.Fk���^yvi-k@XI;��@�gT+ mvo�}�;�|wd|�Qՙ�m�,��4�p��^��-$b÷����B��w	+ٔ�Db�O{��ˑdͭF��j����P� �NfR�fntS��\�o�yzf���سϙ�X �;1gXE>�v��[��m���jѨL�UU��]�\��qao�w�V��*Z�c1nIT���ʙSn�R���S�]�eW�[H��~�_��|��y6�'�ERdy���'&?E��@.���\�v�*�I^�>�vx'>9���[���U��[��2_S���UҼ+k1ș�7�^z6����7�,�O�Β�3=��]ڦ}� ���Pn:!ԗ~�~�1Nzx�g7���x�r���Y���;���{���J�6*�o��}8.F��r2��:+�~Kir���(������R/�Ó�5���G�Rh->��z�����>H����ěɴ�~����,�t���b)y�Z��r�1}J���p9jW8�*k�������h][	���_o��gfG<{�ԣ�t��������?l����ws���n<��XQK>�o=��P��5�8Uw�a?	u����m�6��ۺ�-���;M(�T��ݵ"�]�����$���ɻ�d�E�1R�75l��ـ�@\~�7�
�{��lՂy[��D��R��q�u���ZvuH<l���	�ٯH:��96��V��D��t�wٯ��:9���y�R�ǚ*6��cK2�m���}�}9u�^���U��6�xH��[Y���Kڊ���~�)[���K-��3��=��Lɢr���������ȉ毯��q�  ��O�N�K��}>�^֭�V�\�`ۧb��������t�Fsy�N�Я��yf5�㟙�}9��~�S$ŕ3��yN�w�x�+7����kq�B��HZ����T��K^�%�~�.�����߳���{mm��='���˿Q�w�Azf�H����[�Ӟ泌�{�ߏVu���ح���NwyVJhU�;{-[5��'��5��jOzk��N�&�>'�[Iq2i�F���7I]0GT��*�����U�ǡ}�6���1z�t�w�gA�8=�-��su ~ҽm\U�1�yM��yV'��-t����=(�ӭ�y��Y����Rr��8����_����z��_�4�g�Jℤ���(*U�muu�ކ�,ۺt�o;�ޒ�)� rZn�Q�1���eH��0�7����v4�[];���oWR���B�ڋ�*��p#ӵs��y��Rqjg	�v���;��\f�(]�hZ{]fh)��]�%�%����A��=N��2���tC�ZXv��� ����FЮ�X�Z�2��,}Kޅ�/�9�L�M!`ާ>}��bkf�,U�ךl�B��m"e��E-:��O'>���6F���e�I���ݭ#���&�,b��;�{JL�L�aǆ�E��j�q��TVQ&�{�1v-Kb�P�	[�����4RN�ھ�����-����Rm-G0�/b�;s6櫞�4f��T�r|�{=���u�k��<�rŵ��D���֡Du�WjCK��wb+�Ɋ�ҵ�\b]�W0Q�(�v�T�;w�>�E�Z �o�l��αJ�Ta�S�X0���}���a��h��Z�7fZ������ΚO�R�3L9��X���s��������%�~�x�;�96&�����+;k��C#����؇j�2��Ks��c��P?K�&��թ,�zڼa%�\tw*��]�q�D�����}����]t^�#��'j�S�2�䙋Tt�o%�v셹BZݮ�r�w&�
�&٦��Ω��+��mM8����"v�ܨ�����!v&���t��r7�{J˪I<,h�׍Y*�闘�	�z_M���5��+D�J��#�Y�ʹzt2|�XY[�*Ҥ��d=SJ�_��=��ޯ�����c��2��qioF2�Wm�|KQ�Z�p%�t�j�@�c#2�&���&�^�P6WL5�e����5��7`ȯ�y�K�z6��U�n�٦gsR�T�`�j�������T�1~���ޡ�ՠ�8x�i�b�wR��{����Y�$��CM!�gR(qʼ1�ut͎����8�4������`,�$�XQ��z�c�Ψĭ�MV�N���jِ&�5��5�����t�N�����)-�Ecj-w[��-j�-E�x3_yW��ʻb=e`꜂,S���8�!��H�������W�zs�0sV�.'��X��`.89P�T ^��<�X(R���K4;s\6��=Y�@��`
�9�E4�ا`�YԐp��R�\޾@FDB�u��:T�4�!��ua�W��F�v� �/;�Csp�>���u������7'.�d_GW��,�X)�5�%7L׋(�Q�!�ξ7�MXGh��ۓbkwz��\���Y��a�s��p�w=�l�d���J��"�o��Q�ϒE��K�-]C����4��1Zkڵu��gS�����r]���8�Px��u9��MB��Z�G �� F\����>2�U��ۖ@Ug��;�+$�2VS0k��mߗ{�w�?i�b �Z1db��,V��ȅeB�Zŕ*��DL��̢���QF
�mZ�IP�K��1���Uq�-�,EE�
� �����X�*�b̲�lb*�+"�R�KJ���!��b�QcREQE��(�9jVUkiJ����-@��ES-�E�ˁH�J�V�HV���U@U�X� ����l�b�UYV��1��W82�b[
 T�H��R���"�J�J�B���0�����	[e��#n51��%j�%LK��҂(�TE`,E"5+���lSTUQˋ�����1�EU%b��-�EJ��+�Ub�C2����JQQ�~���3��*��܉�ͫWBs/��-R�);��L��v�F�������a[���,^�6Sದ޶�0��*�����{�H�k�׿���<�yo)Y{�Sr��13;�nw.͍Z|�G��D���z�ǯl-�rFx'=٩�_�J�ފ��3�q�S�n��vVӮ���F��3�I\z��D�-ۿP��B�ߥ2��f����٦J3uP��Q>��w��nw9��X��(K��[T}q��N������*��fz��D��δ��J�ޏ)�=�Fyr�t<#_�خW`��}��sQ�)HeLP�Qv��+��/K)O��/e�,��r�ס�һ�I톷Ymo�v�y����K�=�=4I��貦of8(��;!WX�K�������w���t5���W\~�|�ާ��sK��/=�N-�4��ښ~���U���=9}F�^��~ss�^vS���&v�οd�<���`zI՞<�mC6�|����G��f��s��W��<��	!Ev����ᘉ�2�9[���Ȍ@mףE�]1��mܮ���oa���-���y��q�\��,�>T��.���z%˚HR�AOidb��j�j��V��(v�fus��i�Z�έ�,_E��ӖX�f���2%q>���!�g�����wŜs�Eo�{�^Թ��T�h�p���Z����61QmǇ�w9�0�վ���*�#�m��@������	u]]�T^�͈$��}�/������ȷ&?Nי� ���B�D�UH�]+�M[]�^���^�{"���ެ����<����-��~6�9B�u"~ҽ��xOOv�޷�ڞ�x���|f�q�ٕ�w��j;+�>�S�v���>* ��n�nz���������OO�Î��vCO���+ޮ��Dy��o��SP��>nv<F6�����N@�Q7�װ�!����X����ᷘs�V��\�������ڢ�����5�ۓ8���cE/t��l�ݏ�;�|'R���*z�s�S2{*o{N�yeY�E6�^�8 uB�2=Q�t��j���pk� U<#s�|���8{Uy�{q���S��~I�I����d�yՎ�)��7��ZFSӹ|�p{Y�
�Vy�2���R����ݍ�ц���2x��u�aG+6\ne ��gz�䫛��g3Mn'x�3�m*"��X��k�Z2�\�@5Y)�nKkmB�;����}U_\��\|��0m]H�֮_*���{�7ӄ��v�'42��Z���3�d}<z��_!g�n��x�)̭x�����>o��V�`m �5��V'���u��=�b��HEn�c�
����gM;�N��c�_��n���_lq��&r_<�m
5�Aty�oP��c��qr����d�t���y-{��b�����"�S)�4�c��'V���W���K':4ʕ��D��o�QS����>��ܐ^ӓ�2�5�^�d/������0%y�\���j���]D�`܅T�ҩڻC����nzq�l�쮟y^.��mL�1b���3=��ڧt��U���^&��%�>ݍ���=�N�Vמ�9�T�wuI~}���Sм� ��g,��Ε)�����_9-{���\�����wD^����k(Nίy�ؾ�p\�q�,T.�څFH:���q[�����g�%���}�\`d�,�|��p-�c�oo�)X1�q8C�qG���W������}�.
Z����j���p�м��W1�aĈ@��T�5����z;uq��\��Jy���n���?UW�_U�/%��Ó�]�ɴ�*�#r�i�aT����T��o%�e@�����/?wbP�vL���(��.,����5��R��0e����:��v�:���!����t����/����눸�W��#��_$�ƕ�f �{�B���ޭ���v��a{�"7_�V=/��欝�]u�vu�����uw�7+X����E�/�N�r�}]m��L��
Q��[9Q�6q��T��W�����e�w+�{���<g��ב^q{}�M��xf�=������q�S�;~��s��+tn�4D�w��$���W��z�}.OeS>~�;���&I�*�rUO)�B��O�����9�i���%�+���Ͻ!y�Z�1/�Kۓ"NNr?VR�f�{g�&�}�g؀5�1eε��G�3KZs��f�z�'�u�bi���mv��v.6���r��a�݈��g���R�4yOFr��o]�{��:M����g =�!Z�����R�=��׾]����ߓB-^�[~v^���EP�����K��:7RJ*P������v2��O�&s��ۿ�����1{=��@�p=_�;uSʎ��9i{-U�[��{�5� �/�������ao�8}Dd�r⭩�9U7&�l�W���K>��}�1N.��֐D�l%wF��>�{���U�(]7*�о�^vfvj���}V��Fj����ܚ��_�j�K����|�U>�k�.��$O�zW��ӐO�{�Vt%�k�_lv��(�5�-���o�-��>��ܬQz^�����Ν����]3K��}nW�s_�E�(�]��e�d����?9�g6�lس��ߐ�]ٰ��=��9>�7u���f��J���֡.��3���.-1�#=��q�3�L/��s���B]Wp����	��mj�f ���I8o7m�a�c|9���O���_=���T<#Tz���� ��0e���o=~o3JU-�=zh��lc{_���!���]N�4C���[=O�3n���Jck�P��j+o���Q;�a6����)�Ϫ���ţfo���'E�����
������.A��+\�J�v��[앝Wi3Qwd�ƊA�+c��w3Aɶqe��'��7;]�I��Շ��?�}���W^�z�ǩ�{0w��U��T��o��%�ދ&of|�},o��	]��7V�9�5���n����Ny6�z�d�槹��RL�R�w��y����4v{��K�أZ��z�t��87�=��ʙ���kü�>��K_�SםS���S��k2�N�oo6ޭ��z���]S�����O��m�T�udS�T�@�8]Q{-[�\����TZ�{�^�Oq�_v<�)��n��d�ۡ� �:�]A��$ �~DT~�9�w�i�~��^����^�j��P�m�~�����̢J��t7�,���4Ey�������L�yf��#B�˺�Z,f}10���L�zxj0gt\O9WG:cas+O#$6�_����{Ϙ;�3>�jc*zόf�MigZfz�,u}�����/��YyX��Ŋ�;���16�]�y�X2cc�e�{�Xz3Jڸ�Fg�q�E���PJU3��I�Yvm?F7˼�OC��޻��<�u{t��mvnY=S�n�N�+o��X�g��x����Pv �sT�ļ2�W��a"hWnkmBe
9�T���ctwkWVm;���f�4�X s84��r�-��v�1L�٬��v~�����������|����o�k�>�y�a�|�d���!�V`LtK|g}��C��uaEJko�V������l��q������0=9�Mj
�|���P(ۡ1Ғ�}hVn�٣r��ff�QjמC���ԩ���]�0��|�_[��3.x���kۉW
j�Z���|���۸p�Uބ�&	���~P �� 96�+�g��\�ߣ
� ��#~'�r�>6������U�(�%�_�}f�<Q �!#>����ĉ3w�����ᒟ���ޚ���U�ڧ���SD��!��W���WW���h��E4�^�+ݛ��y������!9ʜ;���	���ឩt�U2Ȋ$hU�(]��]]tX��)�5�ޣ��-����Z<-�W��gثE&���md�^�y1���_L�� ���{4��i[%���޹���I���>d��s+���k4��7KNT�0�{�U=W�`�9x�f�+��}�|v9M�S�ٝt�|�.!0�S����T��O�P�Z2K(�c��`;}e�,2�4��7 ��
�+m��Yٕ�5�|W�����}r���~��j�*e�զ�20;�)�7!�Ы�6�kٷ� ��΃|�$L�x",��PW�����eB�ÃN�H_.z��L���>��������<кf)� �.��%إ�Grj?����j�T�~�����}d���Y��¬�;J��؅�%��t'�g =@������zU�Y���x���~�l��G�Z�r�ׂ��K��4+������]׉�9;�s�%~�W��>8/����o�l���a��9��^����_{ګS��m �gr�h_��ǪUmׇ-jP!yǄeC��2��<�����jW��|�5C*=9�Ũ��b��A^���vj�c��ŕ����|2��L��n�;���q���(�k/��^���s��G	�ɕ��O�)C�
����9nfW�E���S}q��{Ja��/w��l���d�$�<t���߂d��w"�\�c�D =,N��YS��4�*�r���c[��g��h��Y�J����gȲ�����n1�	ʚ����i��A���2�kzzj���EXP��{CO���"9yF��I�s=&���7��qM���
K�9mZ%�����b=��υ�r�Y���U.PTO
��̟u�Q�b�p�P�z�լ��d����*�zc�
��c�1z���γ��"Ov>;��Z�F�0���d�v���d��Ѳ�'3T�;�"������O7A%5ֻ-��Ӝ���L�̌�ʺ���GqX�ǁi�vQ��oL[38��:�mokq�ˍ>��������ޜ��/�-�DU�%���>�L�LG��i���|'�#FW�@/���o&wpP�ͷ׳���ǝd`�h׃T&
{O_DL��U�V��q�k�=u���þ�k%�o~���~���5����UW|$9Ut`��[�Sf�z��%��š��aZrK�j�%��_o��o���|Wfw����"M�t�+�wWpv�]��}�Q�<9(�;��ms{���gvߪ�U�U{��)�u�Mk����U%�޼�R�S�\�-���^#�L�U���G�X���c6�@^�� �ӻ� ?m_��}�K�p_D�����}�l����W;�Y��(�璁�fB@_�ڮ�TP���0��=���J{kܔ�4��r��ϻ/B���\|�s�I�r�U�2�&4�LB�� �^�,�U
�㻻��I}�(��(6B�_���\���&�'�P�.�
Tܥ^ǳ9���{��Yz,mJ����]�2�<4N�|'�p����V����(L/��������~��ۮ��_�GE�}ǌ{��f�ث �C�ko/^�ڊ*^ ����HtRK��`��&��W���G��#�[h��SG�m�2�z�?nŮJ�������&-@G<E�ҽ�	�v�8���w��cf���v�9w�a��S��X�
�W�d�]�ͯ���}_V����;8҇lW�繰������_i�T9�Y�IU+��t.�p\���<�:�L�}��;&)�z�<��ۘ���׵�T�"<b�9gQ�Te�Ut�S%�3�(K�s��3�����>�-�r��ڜ`��yՉU�
���24?���3)��jr�Z��<��7�u�*�S�uq�a�$���b��<��i�3К�:J��ǒ]�/˨�㘳}��B�yc.&gS�Q�2�̏2i�L/��y0����S�6��_����8���X״]t���d:T	U]"Ɛ��J��3����3
�{����' f�?h��{�R,ǭ��h�CEBK�i��&�����߻ɓ2j��B�9w}�grT��:{Ԥ�S�gw	��pp�c���yL9C(S�wB�k�#��ԓ�ܥ�K�Ǭ�3k3��z����Sp�pڇ���qS�O  � R��g�UVZא�B��0��zt�v�G����_zX�;��:K�i��I�ʐ\P���rp��]�}פo\m�Y�Ԧ�&/n��y��~(&����n��ل$����}J!�y��l�SD�D�̇KŸ��7�a�u�,k���X�6�N�O*]����XNK�o��qJ�b\��`]�9�L���QE�ؤ5�7$y�8�|�( �Z����+E꺜-�z�t�5��S�>:Z4%e����z�m�R��\��L�ݛ{y8��D���V��	�lI�n�E��V����-��鷲�^wl�2;Ϯ�@�^��*���	f����O* �j���V�U�j�+]ʺ��j*=��m�Yy��(�0�c�R�p��\���\U���0��4\遭̰;�W%�'w��*�AE�b3@�,;oOgr���# ���k������쵨J���օ��,�X�ҝu��Fy�ܝ+��3W`5Y�v)��_Xv���U�g�96�RL����,Cɀ`�*y�ͅ#��ޅ/j�; B��"{��ǯ�bZE!\��h�\��;꺵�V�]�v���|��1a�fM9�U�F �*�V�]��L��r�]��<��5���U���2��ͥsf���Ӧ �^j��:E\ �<95�����Y�M+�,��1�2��kc���VNۻ0��h�w-�����.�Zh���앩̃3�C/-����P2o쫺��������1��:#)'��Ҡ��-��Q�|j
�4 ��M�m��m����ef\UwQ�{�A��z3��䧼6�K˶��c� gN��;^�'u���3Xp^���&��Z��ǫ��c�4�^�ihj3h:8#���s �'h=��ENt��)5R�k���]>����f�l;�͙=9� ���k�|��㊭�Un-ֻ�6�>���3gM2�Kl_.m����ww��y-����^W��j���0'��G�^�/�AWE�F�e�/�=�*�m�=�7pK�Z��w��]ꑗ���Z�%�j���aͮ��΁[�b訄����Y<���o�Vqt�ɖ�{��Z�N瘕ǉ<b�ӹ�:B�t��s|�>�����m�\EJ�I��m�(Z�����:W'k-��gc�e�t
��F0�)�I�Ͼ��(�������'����FQ�|�f���5U������AA��+�[2��w�u.�bB�%�aX�G(ra5^v����zz*JnR\�ј������Zr�'Ji^1z��C��{���?S"��QL��nu�{�z��X�&�R������hX짜��ެÌ'�̩��9���29aL##x�6�� *>�T���n�D��ێW���V*`�t�� ��G��z�Dl�4)�`��g/cڭv-w�\ˌ�/ѭ��	+���z{`IS��o{��@@�C�&�}���ʙ]��S
��2��ϩa����?Kj��|��V�la����[��hf������a�sss��޾���c!��K�1�+�2VE!YXe�EQ����l��Z,R"\�2V�P�)1�Z���AJ0���$+)Z�֤���p���F26��³Qa�b(�ơD�bfPX�صinY#�UPč���*B���Jc�¥e��
��\@̤Zʶ�2�\��E1%K�D2�J0I�Lem��X�
H��F��*V*�آ&2�3--���Xc%q*%�#�Tm�m+P�Qq�.P��Y����U`�[r��$33�++Q��1(Ȣ�T+b����0U�QX�[V�[+A`#�dR�+Q�jRյS.aVT����E�\��©U��Lpf8\�X�Z[q�-m)DB�lLaUD0�����D[e�k.5TA2�(ŹjG-[�G���5G��|yoUÓ]�:�����"�ƹ�����p�����.��{q����W$=���K�SC��Ӻw&��Y�����꯫��Ry�{��ﭒ,g+�,({6�?Uw.���D��l�(��3���<q�D�u�����t���7��w	޳��
�t CbaW��h��`�9J��EN��`Հ��|�-�W��39�C�/!����}֍�q����T���-��\��n��M|2��9��Ѕ�����wu�	ج�lu2����*�8{)Z��KD�V��L�c4���l�����ҋ�{�b�����ױ0&:R[�%R�#SG=�3���wD��]1W��hO����bq����wyҊ��xp����v���$�d�w�tb9*�%c����]:
��Yg�¾�; �;�i6����i�N��YXra���	RGsx��	G,��ބ�]����� 	� 9��0�8��f���5��=������M���T���&aa!����Y�H<��!#'j��q"];*�=��r{�����_�2V�Hpd�8�Q�%G�� �:�u:�t5p�SOr�9+���tFS�{�e��6o�v����YdW1�g�aL�ow8E�L�(/�[ՙC��(p<�׹KH��|89�v9Os��X�oA͹G���+i�c�f���.ҷ:���Ϻfa7J�#(fM[��0)J;]M9�]�c1vTޘgfr3�W�_|��Ko޴#���fW�q�Y���|~�eM���D�
CuTNi��J��5�`o�NHb䝿t�^���x�pe�'�5�"��}SɌϧ�)���� Ү3�˯L>�o���v<��WZʞ�S��xL��V�}-f�~���i�.a�LPh�F`la���x��^�>��ܲ�W2lW{�(>A����&S�B�hʒ�;�u�������|�>����6v�qW\����=:�B+ī������4��H>�{��ؽ-���>��Em���x�>�!��kʥ��\�)v��~���"z��;][��3���
�< )-��,�'^�lٮ���y���\���ͬ�ֈR-�����S������V<�ƥ�q��C��9]�^^Uw���!��S�^ŧE"Ni��}�oSۙP^�FSZ�б{'*n��j՛���G�������B�g��]����p?]���T���WB\J�h�XU<�����u]V�ܽ�T'�s��{���y����ƒt�6c^���m����Cb�*���D�O�I'Z���r��#�8��
� u��ߕ�坯�=�!�LN�uyk�'����v���a�&`V�'2
L��0�SvT�]8�[��}�}_n	;���{+?���V	�~�z
�ƀ���F|�T '��ϲ{z����g{0�#�����n熈�:�J3��`���6ϢX=P��8HǢ�'9�p���w�z�s�s�=��R�L������/x�L��Y�H�]KںX�������I����p�c&3�a� ���;hן�׎Һ�E��|�\g&Y��DpF��tN�`X��#����˜���^`��>M*�}�0o�ީ�E<�T��s�~r��Dp�y���v���]��~.Gz�6Ƌ�X�,ѯ_�Qj�4�|�t�U'<��
K�fWa�Z����]/t��5���]�$-�`s���*7H����Poj��G@�a�[��k8+͉���rC�C+��s���$q6�xs�7᮫q�
� /�F�񫼱��YE^PM�޶�����)�X�
��)}S*�'��W�_]��)(.�ךi��*��3'�7~�0�Ors0��=��C��@U ��e+���0����j犪���L����
���f=�X�ۋsX�9�A!�̫���M�Ш4r.��VE�W����qcz�ޅ��\�8팹�����\&��Sk&�����.i�f	9KE�ruژ�t{&�y�W��]�o��~�<ƣ���U}_Vd��9�]�!�+���gj;�Y��^y	��ޓ7�N��kT���O(�C��z��[���8�,Oy��ϯp�S�I��)Q��0��+��V���,�:�;͹:��j{k�+�C���7�{s ����2u�RnR�g�}8��}�#��z�U�N�{�k3vÃ�oD�8My���"?.�_�z$!�U�Rҧ6=�j{�����5�=��E�c��+�ì,q��\_�`�Ί����@�:�X��X��m��cvݟx��a�[�������jw^�MPw��ȏ@�FY�|]֚�����y�lg�=�f5���T�����Bt1:���=N������ypy��#�:.	��.��.�9'>�|���a������i�	~&&� A͸2����+���wR�6���:�{��5rkv���I��b� ��D̨̙�F��:Ͻ������0xf���v��ooL�3���e�t�z��Uo[!}���`������֥[MV�ظxh}I��ѱ�������	�H^8��ڷ�	{���Jќ���kǗ�y{�
�����u�Ü��eU�/����6`�O_̉`\��a�Z��82��YV���s�΢1�S3��R2�wR�m=hq5��R�J\����i`���ܤЮ�0;�[�Ic�g~������I�.�d�L|"0p�]q�W6h,:O�����WV�U�L��T��WL�2���,{3�s��۽�^[�2���3��O$T+�u
�	ګ=e]��{�=���k�����&.��EY�{�q�O���/2�)����	
�2b�s���A (���Yg��g\W��޻���-7�;��>J���n���T�B�/!���ϪApud��TĄ��������f.��:X?����	-A���u�҉/�|w=�껑л��&&�g	�/0#�w/Իt�T8l�Uj�T)��I<��:1�	�����Tjf@s-��n(��nI��w*�]�`y�Xe��;���/��_�P��X�,nv�doF�(]<�Ԯ}���;p��&^q9}�;ܪeo�UY�ˊ�`�2f7�ܽP�~�������u���Z��E�U=���*�3��,:�!�V`Lt����"�^��O+t)�o���[�o)U��K�`K�eq��b��ʶ�}L����5�
�~u�@�J���}|�g�{a�n��q�9](P�/7f��.Pԥĳ�np���x�CN�E�I-���k�/\���ug�*��5�A�iбbK��޼ܑ[2���B`��:�q]�F��Y�o�R��u�V����5�plh~���׾����i����䱞�p>�K�WPu����?���Y=��y��R�0{z$K��#����ʂ�AW�q>�`|e$�z?0We���Y��=�
fq��v37���1����=6.}s�){E��)�fU�d����U���D�Ɣ����]K;�brnO���˶��m�oo�	�*�pd�zD.�Q�^N�� �f���-����T5{ Yϟz1Ǟ���[z�W�9U���py�L��T�h�Hd��5j�Uݦ<2{�e�>�K��s�����S�M>�����ڭ��ޯ)eL��	0X�e��x$���iK_� >��j�_o�*�|�	�G2�����O��-9R\��\]�&�Wn�n�=���r�|��i}��Z-}w� ~|�881���.��OLu�ӗ��?-�m�dw��tvr��'�ޑ?�B2<J���K�[� (���vu9�b��ٱƹ�{�6'٩:���ZU�[l����kʥ��\�)v�-s��g*5���C/�B�9\P.l��w��dǣڧ�qR&��&��X�ž�4�l�@D/�2+L�wU��""1tu_<$s
4w(��Z���v�.����}�jcMM=�r�w2���1H��W�=EԹ�v�9݃�2`�������*��Ix밉�>��#}<��q����ϑk�_# *��t�1S�U;,᧽W�t��4׼�U���X�痯��LqVq����u�kR��<#*I΋�/*�;��C;�Z�:�6{�c�"+4w�����X����Rά|%[GêY��� �9�U�Á�X>�O}�J~o�v*Vz��g��%�	uS������h�TX�a.%Y�Qp�Wfu��G��enu��37��,����C@��KO�`�K��sUl�"v:��.Q]�QؠsU��)�__y��>��i����*�5^��aT+E_V|�'DE���n'���Wf���T*`�l���~&l_G9T�nM�6��b0iVt�>L}������W���ϣ�Q��f�	��x�4[}��"*��Z+��iz�&Y���Q�(63z�Λ�7ӞH��9xVO���M*�m1�7ŉ�N�*�y���|����X�SȎ�9��v�v��8�l�4	Z�5 �Z�\�L�}N�Yc��t�Ny�>�낱]q��{&|6[t`�Y�HL����w��W8Q��VV�c�IiX� ��n{��G_�Ѿ��F��yiv]�{e�o� \*^^gK��ݮ�e���ҡeў��>>I���<� Mc���[�%�Y�n�s���esn;s�n+z�+,�x~���U���ip�J����5���Q(5�j�1S|�!����7��i�;���'l�N��>�Dçt-`��몛��U���D���E�0-�����t���m��剎�)1���ႥL��Ւk+X�
���%u�oոȈP8��msr]~^˝�Ie߷�p@�Zd ��g�
���L*��U�!���`9�vfD߽j8�\�"����-��wL�W�@C: ������(w��2��9{��o\�F7//,�s�U��tKD�{�0tS�i9Z�**��A�&4�c�>W廮x�c}͆_�@bWg&0`�ZP��6ǡʯe�����&����2u�RnR�w�]�!(8��[�ݽ،{�t��1uq����>Ä��ҺF9�������HC���2խ�zA+�e�J�ԅfl��}��t�3����W&(��e����89ږ���yk��A��ZB��q7��幘3��񬪩�׹5Aޫ�#�:7
�>F�����Քk���1�ܪɘ��LB4!F�=�h�Tk���\|N��M쫊�|m k���cJ�Xɵ�k7���S����)$�)���[t �{���g����%�~�ޝٝ��o@kFc��~�^�~n��ԗt��ɜM�O�`*f�͹��j���p����ٵ��eJ��;c��.r�C}V��2�T��=L�7��D^^hmT�\&zzm�O�����ʬ�AJ��WZ��B^�騈snw{Ƴ��j(��;7vǷt-�������-�G��(p���wQ]حU�w�\k��>��f�q7=�i�����Iz���Ͻ�T�Z�D*�Du?���2�u9��*�jV�{�u��ˇ3���{�Y~���~���V4�Y�"��������[*�؋��d�m�+��U�s�I��-�!\<M�J�f��!��H���<�T
�4(S�Ĵw�B�l�)=�a�NKq�����AM�vxeM�ƕ>j�����f�<=�#&(7*yV,Y1=���k*N�ܓ;W4��8��Z���{yH}S�3���:K�i����՟K�5����+ַ�|���F��{Æ�$Uu�8g+���^[h=��wED��.
+�38���G9F������@X�F�'Z6}+P�_g�^��x=���`����b��x���j9bA{*���)Mn�.�W2c�`D��+�X�g�V��Ўș�g?=�c(o	}��W��i��be4�N&PH��a����Lw\#���������.嬒
�ޣ
/"K�F����@f�[���v9�k	x�A��SJˣ1;�&�=�ԧ���!~�%�?�:���s|�Y��>�j��L�r�i����m�mɂ��,To^\\����"QcÖ��/�� T�o���e�{���k=���A�t��~����lmlu0;�iZ���鹟
cD:�u�χ���ƌ��h4�7����3u�k�o��V�B�h��p%(eq��^�������NT֠��!^YW<���N��+Ӟ�b�&�&Uޢ�`R�u{���_o������Pq���i���8\�����0���uµ�,�|}��Ė�J~`*ؼ m�;��'�mk�Ch/���3��MS�pW{��g��h�X�5�CM�O���}f�<�)�!#��%O���׶(���a�lG���}��/ʷ���^aV2�XD�;A��=َ��ud��|�=8"Π�ԔOO�ꂽꜩ�Y���g�z]4T�"�١V4S���UO�&N��]�9��W[(T���ꗪ���ڭ��ޯR�FW���<��W��b��#���u��*sn"+���Y���')�ևE�U!�5�XɶA*��)��xr�s��WN�eho�֜9К��{��2�����`��DښEn�y:,�u�w�p#����;h��*fg :�3�KoFE�M�tE���֯zy�/�_���e��B-G��)������5+( +�R�L<=�D.�=�����e:���[?X.k�D��Fցy�%Z�2�/�iP�G���:�������	xq����(�}����B�̗I�gd<����3B譄�%�!�A�Y��������ѣ�Ez�����Ep����d�F�;͙�MΩ7+�3��*�iw�0� ]wuf �խ.V>�}$�Z5C�������S1V]af�Or鲖�H彶�{$�`�?\{�J�W���|ގHQ#,�]�f�QRj�;���T�K��,���`���t�)*!,���������\�c�ZrU���|����ҎmθeԨ��.uÛo0�@�n�����Vxټ���<�jŸ��}+��7D$"��f,�eF��̇Da<�chL��=��c�tͰ��H}�p>�(�x���i_<����R�N+1�9�Z��Z�H���O����J[�w&�l�v�EI@�(���:���tӃ�x����{�2�mY��x���/0�kv�UF�kx�a9�[y��F�lS���V 3�A���wB�կ�㇐��3d�!Y<�^����~�~=#�3e}��7��i�܏!�n1kl��'�5{H,�aѸis��Y�yi��g�Z�����A���*e�*�����ݸ_w1ۺXY�W�p�c�� j�_'��}��"���"O��R���`ڜ	�r�m�[u������RU��ck��<�e<�Av���tl�n�|%��I�V��3叶���&��q���z��)�ÈWcQ�.|@u���5w�fJba��()i��}�/�嫮�����]��y�t�620J�	���ѣSx6l�QV�� ��;��h�َԴ�K��A��,Ў�b�%��������5��復��o�#(��z�.���!ͮ+��������N
Ko�`wg�t�a�Kv1��i�����e��K]`<v����5�S�֎��u}��h[*ؐ��W��!sݦ;�ؙ��W.��@V�X�'tB����H�Ȱs*pS�8x�r}{G�Jr��r������S/A��{̎�k��ӝ�2)9r������9�&���T��_�+ҩ���.��f�4�]Z�n�9d�ݫ-N���[��M�D��S��+�Ki9J�� �9�s+�b��RѾP��uX�|�Μ'l43�1S˥�E�w�{��C֟lM5�mQ�^�>��w�^~������Y��l��MXQDETĦ5T+��A�ib�șh�Em���2�%f+AUKh�TR��TTX��Qm�d*"1e�����nfh�U���*�ұ�kf`TAU��9aV�A��*ĵ�J��7Ȉ�X��iF����R�)��֠�D�C-EH�R�r�J�m�r�F�Zʃh"-��Q"Z6�m�D��V�`�J�p��
Z�Kl.f6��&)Z���-�s18��-���m�ab(���L-EƘ�K-QT����*V�j88U��2ت&Z)K�ֱdmhҡYYF�T�n
 ���T�5jҖ��lŶ�2���dm�S-(e���X�-����jUF��Rҫ�QTh�9f8�Dm-F�[)"��� ^���tg��]
gQ�k<��]�T�Lp���4b�b��^��}�ސ)j�JBuoJ�n`�������u��+���M��@ �~5u̪�@��3�?��Z�U-f�p
���{��Э��X8�a�G>�����]jE1�F�گ�G���?D=������2����h�D�o6v�'��]p�l���6�q�`ߦY&�Y�*��Wu�FB�؅���Q�b��T��?G��hm�`�,&�t$$W�m9cū�~��"�}r�=�ʘ�&7�y�f�8�:f2��W��J`�\۱�.2��7�4n���#�O:�D���qܤ���ғ���q��?U=�+I[Y�[~�=N��-jP!}�����ӵ���yF�w�y4d���,o^�+�"Z<���ӭ���[Ű�]<u~=���^�W��m����>T66�F������/,]����L�s<����~��5��YW���3+�=��׏��q5�Ɨ�$�[AWG����KN���3�,�9��`^����O�`Z2�MǾ��m�;�_j�~f)����5^ϯ�
�W�}g��I`�},?w�>�O��8��F���aY��U�V\��	�XsW�ג��wǡ���B��0$ q��
�v
��ԫj�^psd=�D$q�4��$���`��v�_6`���	74:���¥�I�W>$'r<9�}�����L�K��@�[��K�ɛls����6�ڌ^���Y�K�o*^�,�,�_{=��]�4�}>Jc,�OE�7�;��Z+zj�>|.qʙdr����������rkr+L�]�~�Ի�L�{����}V��뿽��]3e1*�/m��������[${�������zP�}�#(�pQ����Z�M>�w���:�I�=��N����S~Y�S�t��jh��9믝�
~�' 5�Ƀ�}�F�l��O{�A�����I�%���:J�;6�JJӕ������]4�u��d���e%.�@uAҎ�ï�OL��xӣ�q�b���Rc�U.�m��Je]F��Z�����f�bL���>���oq	���i�V�ݰ"�p@�L� /H�0W�݊c��ɛ�Л�1/?�|�Wl���qށ���)���L��*�[�s�{_Jf�͸/R��ޏz/7�z0Vf��l?[�p�j�����
�����=[CL�z�W�hC׏Ö+�;�����ppn[�ҥ15t�j0�g����V��wj񌫺��$��̾O����.QC=�KEf�3�OG��wT��*����_�.�Ū���/k�&��5\�U��4{rx�Yx��H��YH��{�1�h��f�4��b��鷫��i)�`�꾀`ǋFP��U���Ep�qpuw�x{>���	^�b���^��L鍿[�u��d'&����T:4/�<�ʭ:M5����}gU�0�iL��t���Tr/���|���>~�Y��(��v)s��ө�gq߲_qʞ�⨂�vu��wDK����5v���	/dN���JL\�P����-LL�3}���Ԏ��ɪ9d`�p�ތ��o{7۝�ڳJ.�I�B��P��h,2��1[S�wxg�o��˃�佽��+|���l�b�Z#�>�e݆��֊UW*�W�|!*�نd�D
��pc��4�R��Eصz����vvz��Z�/�t{�$�ΒB�j]��x�N�*�<����8���b�yvf#^�*@��Q�M".���K�x8r���
��z{E:D�-�'w��OY�Y�b\��s��Ș�9���L�N�F��&�][}���m���L�,Ot�q� |��Z!67k��$(hR%�J�H/��Z��B�мJ�-��`�C���]
���e�Y,�D�ٚoH�����ܢ����l��f�������Q2�Vz��j�m\bC����.�6�̈́����Y�m��}9�J僱���Q�0}{[��5�+��o`O�w7��)O�H�]L̎��ܚ^r�7�(w�t֧\���g~���5�K0g�lq���7/2��!��B������dB^���������/{s VY:���Ƿ�B���̩�(������B������M�Ƹ��#^�`t���v���a������~j?.\�^��fQ&C{��oB:̏��}ݭP�η`xO�%�p� R*º�bcI>�qPv�z��.<��^���8�h;iQTڧAIxΓЏ#ygʧ�P��2��f�'���S���W�í���>ǫ<<&��~0N��x�w�長����;H�0�c��/�^�-���jz����=0j{��٨9T\(xg�c�&��;_Gz7>~챡QkkM���>��]9y��Y��k&�
�S{�.��Ƶ���12��������wx���U�����Oj�6�}�Lz�P:�	�O��z%����,�WP_o���ª�PcΜ/�F\��ﷶ>��f���X���]o������$�z?0l^ :�Dw��xj�qF���pm,�s|��6��q91��#Y�B�^��UQz�Y��h�E�dT�S,��n���=�wq��U���.	\�����X�g(����W.�Nc�n�m\`5�&V�Y^T�/q�P[�R�Zc�g�Ɯ= 5�R�G�
���������HЅ����<��$�w�uRi�
���o9�:w��L��5�d�"*���r�tƲ�j<�#�Le|J�)�A���|��ſM��N�\2V�GFE��ꂽ�ʮ�yk8=O�g�{�t�S,��vhW��6���zs���*�J�{KϮ����p�?54����-W
Rs��ԤQ�陸�;o�cy��M���,O���� p�(�B��*c���9���-f�~���i��x�6M���y�.V��*z��#>�e����&�p��������0w�yɿvd�٪0�n.��R���;YN*�r�z�u _��'��TNL��U��FBW�\]3|Ɲ�d��p���'BBEz����ĩ�w�.�0������{�GE�.�um�:���-��*�����>wDA_k�F@ک-�WK�-T��>4�k���^��ݿw������}�k�͂��J���<!�DEZԠB�8��~'k��W�8JG��4Ja�.�*s&�筃�$��gvS�e�j� �6��M\)5��k>���݀����&��Z�΢�0`�3"�2�.\p�	��VL�0���+�}�kYzdӐr.��V�T�х�����Y� J=��E��n�RS��XYN���Y�����p�aC�^q?{y%p��a귎��q��{`���.^�iqr�If�>�[�u�(��<u��qw-`_��z�Tu	��n����4mz�&�=����1S���}^3}m�G�٠n�����	U��V4���&�AE�߳ګݭ�� OK�帲��?	�(Ϗ�(鿑�}����*?Kf��廻�1���^�$�n6஢�eO3rm����9�˃�-q��W�/��5�w��·�7�Wh�b�
�ܪ�a��^K=U���/^HB!��Z���>��֔LC�XS��(���'E4H�eR�S�i���bo�v��yHb���75��^c7xL�A��n1�����Dhv\��W%
5?$:����������ڸ�<����>S�v2�p���u>��:�ƹ8�fLEf�!�>�i��,�ټ"��q��m��V�Z ��nyzB}��]*�]��y�Un�k)(:z盵�a6=A�P�g!�ʊ�{uԕ4�d �[zQ�~�`�;E�U�L�9�`Mm��>�:�>[��fe�ָ�#��Z=����"B�T\^��w��;c�����6yJF^*���v�����#�eˮ�.�j�d� �gR/���*�,&��i��_*%{��b3�b���Rc��ghw�2�2��x�5u�_M`w�Y�7���o����.T��5��yy��DHP��o���D0A��P%��A�|�M��痳_0l�U����[۳¶�/���1�w|ߺ�U��(:
����*j< �a^���w#|XB�C\��Cֲ|���X�Ȳ����I�*艵{}o+�̧���MI�r�X��x�X�2�:��Q^���y'������j�g}X�����8�;�sU�z�� �,^�Z՞�����w7�w�<����+�y�@��'�Ó�+���a�=K��ʑ!^Ǫ0k>��w�[�}�ְ�Ä���{�~[�7�R�^���;t�[�y�������\Hd����ʚ��=pk�����I��l�9�~�m#���}�h���UӡGP�P��l2t1:���S���*����[iY��d��s{�
�8O�be]�3,�p�Un��u�	_=�97�Ps�.�z�nV����T�#���O����c���Y��fB��\�LD4����IM�ER������F�>q�XkZ&�x�kCCA��&	�A�d�1v��O/�m���a��M
x�F�nM�٣[�Ԭp�,�鵙��-��-�r�tz���m�t�g��ع�+�Rw�W�e�g^;�!��9Ww�b���I�r���3KB�O�xYL�G�Lr�x�/w��嬻��P�t�1̞2�8�j|\LEX��n�62Uܿ-�͍<��׎^�C��y�_3��e�)ϢF������a髵�m_\y�ŏ�"��(�)�f�Og�T�%�`޶�w��pp�d���h��(Sf�
���t�-������	��=��	msق	��4�8�_�^f��3sP��#&(4�Co�c��#�׼��b �Z�UY�ybT���
C8�T樉%�4�P����J�B���s��z-��Z��cà$]���<ҳ�~1A�[�xɻ�D�ŵf��~�s�c�}b��]B}��=YN 4Ew����V�*C�|�2��X�B�0���/I����6�Sa��9�$�r�U"�AIxΓ�4��J��]`{M*+���U���~�Q���O'~�!�	�Z� U=PJ��z�_q��r��o���S��`�^�4U��^�7�MG���XÒ��U}�؅��c�o��u�P�C������U�ғ��Ѱ�%\wS\U��K���bZT�z��\$M1RZWu�O4�\���*A�⮟�!�N�f��n�CX�pQo#�m����WʠXWƵ
޴%?�#~���7�zp�#�H_W�;h�¢��=�o7e?7ɻ�%oA��V�\U�.��}�t8V�)�LL�ja�b�Y����g�e��q��Qr���+�&:%���'*z�/�]A�m��9�_8Vu��W��]�l]�__y����f�Ub�+ʪ�P*�Ϯ�&r��L��`� ���RfL}�vj��}�3�n[����J�;H�gS�s�j�4�L��K��l��w$�m_��g��aG��M�fg�Gw�ʜ.��}6ȏӱ�u.��U8_qϦZ�X����<N�n���{鳳��r}f�<�[Fj)��K�zu��+�u����\�ע#�{����P��;�o���}�hTWP�z�W].E�n�>�=��j�R�N~�d�x���*t�E��N��7�V�X��  _L�t� ���5t�[�
�U3�g�)���-f�rV�2̪w=�dO�ޫ�>{}���� ��OU���,���}�.�����}|�����f��3'�Q�b7<T����D�Ẽz!������M�2��`��v���G��W���Y|MZzO.�=s����S݈5���cnqW���`��v.x��� ���&Y۵������ˣΔd��BV��LZ=X.�+7)��T�x7�s���3ng^��op��TW'=�<��w�J�HM�V��qʞ��LD�[�GY��E&��r��~���������؃83��(8`yP��eIdV�T�O��d�7�<U�c-�_f-=�|�q����۴�;���8xD]wDA�K�$�6�X_Nͯ^_E:���½cq��!�E�
TJ��ڰ���V5M������k��*�;��]�ݞfۗ\���VԹ�ح�/��;�׽�S㨺kUzfP��+yK'ً���Vk����i{����¿^���[�D�a.�����d���Ez�ֹ��S�dj�����mgV%�D�p@7�o���=v�to#rwن��-ނ��}׊��{�990w����`��m��U����8{J�u��P�l���"�)R�)SOj~v�u��8��S�HϞ�����
T\��������2���/��B�Ώ����n�^�m�A�=T���e����l�DO*�S�\����eWޏ����~ʓ��h���#�:a�1����Kx�v3�ĸk��
J�J�@��+�ץR˷�n`���~�"�	������W���C��@���A����2��<��e��$��I���Â�}��=I�{P��+��{ް���~;3��_���Ě�_w��)���6xX�y�Ȫ,A=���@��w��T�/)��zf'z"�8��6����M��b���˘k� {��-��$�������:�S��{_ht.�-��W;�`�W-�6rv�R���zjWh��pu�,����ȥ W�s/q�m�N���%��mYal\�^R�u�w��ŗ��x ��7�D;N���� �H�$l��h��z9ۺ�ж�;�%��煒8B�x���E�)��oe�Q�y��>��z�q���x���K�8�W��D����!]�p���M��m�k���*3�]DKï�;BeǏ���:�aJ��[Sۼ�pe�cR��n
�=X�5������k(�^YW��p\{9�R���m�����/�w�ӽ�/f���<ͱۍ-�9I��kzg׭wH⺃���DG��w�G	�Fő�SEZ��xn��V���ب]^�i��q��6v��ZV8��-tx��+�[ʠ�/+56��h7�S�ՙODkl���y�������j��uOF�5�o�AV���X
�#U�%=��r|���k`����uz�jĢT���5��p g\��-Ь;G�D�Z�lv�E�s�,w�a�t��%�z��G���"����Gx�(7����g:Que�,�������E҃�-�Y���Lk�aW9��m�-.�+�F�;��R��ҍ���z4吐p'}�m��n5ZU���[�+5z�w�t��t���j���H��Q���x��7hflEj{����l�6+9��,�N�*�$��ѐ6˭b����YZ�b�k)�o��۠K�3X�f�ҁ��^�ۢ��a���9�q{��xk�_o�ΚA%�1���
���ٷ�Xڊ5.�ᑳT�q&�뷹R*��qO�杕x\�u��PiP���u��T
�)O,1�g+�tǽcW+�[�����*�6��n�8wZ�Ih
}K�Eؾ�x+��4��VW��m}�*�p�����7@9Hz�	7D�s�5�7Zu�2���n����=U&^V�N�j�������e��G��Э4������*����������6�0G�p\u�v�kT10�q!�=�j�D�I[1�;k"��l��R�!i;�����$��}��`iC�A�H��s7&�Y�w�t��#�8�nnv���Y�S�jv[u{7_\dQ���w���o�N�:�\�J�����Lz��N)v��ٝ}3\�S�p�{~އϵz�]{wr�H:h��X��N�\O���YS[8đ�*��f�:�25=���8�C3,M�立�Ū�(�Um��8Zc�(fJ�R�R��S38�Q-ae�lU.f9Z[j4mZZQ��*nea��Ehƭ*���X���K2�Q��X�m�-JTmcTmc�)��*����[m�F�VZU�"��	��F�mJ�-+kV��T���Z%�*��kmKlTj6�-����J���33�[����[jQ�Zʊ�kP����[EZ�Ymjі����imF�X[J��.9E��R�Qq�F��U�Z�6��+[De��V+emT��nZ`��cZ"Ѷ��J��-�(�Q-*��YJW3�*�kZ(�k*Q�KlU�-m(Զ*,m�eL��H�ɖ�F�$! �P�>���1�WK)�vjqm����ǨFGuk�J�^K���V�ʧ��MXu!h�X��˨�[PA<�NW	V��Gjk`�5Ŝ��{������@�TH�f��3Og@:���y�^��ն�?.;�юe{��SK��6����예�,2�\�*F�TA�Ї����1��'����DJS�gWhٸ��c��r𨧤��u�Ñ4%o#�Z\=�|��eB��>�7}���/@D���^������ܼ���sXʩ�0̣O~wD)�r&瓦=����Y=���{s̿r
f�g�����,P8.�ީu�S.
U2��VI��Y�zz�YAꏜ]Z�ð��C�RLwm�a����� }P�d��#>��_x�tA&��|wyoH��'l}t�V�^_u[�V_X���=�g���fwL�W�HlAa�]�y��g��K���%z6a>����<&�y��z�F�ZG�^�}��T��W7�Q��2�<�*�OI�x7���9�.�>r�`�1�JT�A~�aϮ.��d�5Н#nI��!z����5ފUZ�*�}Of2rm�<O�nj�>�^٧�����n�"	������=�ۮ�߆y,��4�'��Q4i\1o]�̺zT�E�x���}�h
�%�W�6��Q�=�8>��!$:�����*��!CS=�����X�.ʋ�^�vQ*\�:�3C��C`�Riyu`�9VD���G9:&`;ѷ7S�Ġ�L�^Z:�\�&T�
�=Q�Y5��;Y/����:J�\o�����ok�ֽ��Y�O��BP���9KS*���EOMd֧u��5A� ��:����t�����Z���^=u�}u(Q�"�;Aa�W��]�0uS������nFq�v�_�O�o8���o�e(���8��%���Z*�u*�U��J��aϦ�}��͝pyָ�{sۯ9m����k�׽�U���4E���U�����Q�T�<-��e����u���Ɲ���#Ԧ6�c�p73�S��*X5�i(���|	��ѣ>}�+=�_c~�982�;G2�
�K�soa��S���=�s>F�vz*]D��<L�'��S�����M��q�xd��O(L�pW�9hy�'�1��5��Ts���"�,���0;qZ/d�ό���(�FD�ù�kog���b,�TqV�UK���f��!\GR����D]n=��{{�nXJZ��r��y]����r:�9�̢�^AS��]M=��7�jɓY��q,ŐoD*��3L�Ui�:f�Ғ�-isX��)���Cה������.��W�R�2�R�`�lq�P-��̸CA���j�E�44V�H�vwT��6*v�3=��4����c@Ҧ��[�J�tmԺ�����_"Q���{����:��u��3��dXb�
�,lW���UCٷ��X�ff��Q�׫@z��p�6������n���m9`x5v�a8^�)CtPT&�7��]��Clƻ��	kD�����Z�*+�:ω��cN��<�g�q4�u�c�l:	YY�{�]ϻ�=�hx^g��~�Ր�Q���� ^� R���`�cc�����w7})��QS�Q�A��/��V=�}y�i�Z=�k����xL.<1�xF}7Un��{ܟ�{�����F[���ת�}���+ͽ�%~2R�1W
����4�x��<|=+&���1y�1'6-�p��G��iu���U���>��b�;),g�/%�w�)���e�x#���J|�a�2w�c�b=��ɱW�=i�ڗGsB���/~�Йʻ�@'��Y��X�9V��Ŀ76��^n�}_���gS�s���.!S!�L��`<�}�6��w���[�[���w3g�.�$wӅ��Ϧ�|�;�g��u����tϽ�tP�QFWu��q�=/f����A�'���r�����g���xh�W�̌�u��K���O�V�/��=:�Lu/�?{w������>ڷm�6����WzM���~@{������E2m�����5u�ݼh�"�T5Rb��Lt��x����r+,� W� ��a�_nM,cQM>�z��z�".�yk8=O��z�]4M�Þ��SO�w}���t�
�)в\3.���\��SO���֧�R�~���*Tò��̰�:=�����9>�(2e��2@u��VT�ߑw�8?{}ԥ@wEY+)-�FX��z��,S�!��u9����S�����ULE�K,�v�u���o���3���F�u�M����CO���TY2���D���mS�����}2�7��~9Ur�U��{W}�����]�=�,v����I�>�'C*K"��rǊ��S��$�m�,�px�7�2yY}�vgb��z����j��{��z�� ��d � U���I�yg)��s\���Cػi�R�b"uo��ꣽ�ZJ��j��Ʀz��J/���+L��G0zo�Ev���L�zݺ�>��zҼ2%��-���j[�X�J5�h�/JA]�%a�Fn�d�����j�����l�ǭZ,xw�h�����p�g��Lo��� 5gZ�8,��K��z���5ꐠ�����b�5�Ö�,:a\I���݁*�1)x�5h&w�D$���)��E��7��i�^S�_Mی3tlr��p��[c��v8Ϥ!J]ְ��^�ϞWJiU�yf�˵f�k*K�Gvq��s��<�z�[T�ʷ3+ު.J�y�;��cףDٲ�O���g˖�z���?//w��d�~n�\.22j��{lL�S�1M>������V�^#
­�(�|�����y>����$1X�Wg�]vp��	��*|\������-1���[����w��H�=�aT��u�Y����8*�%S�pM���yV�1ޮ�;�.�����:s=�^�r�WbvU�F:�����^���M+�UJ%]��'���7�;�@�z���q�yl:�OH�5v�Rr����"8(��|���B�?�MWo�!��3���Ƽ_���$	G��ܩ��ޗ�/
�W����<3�h��&�#9UtX�u�.{3�}=;&ݸ�{�;^�m�{o�(5�TX�`n^q�d���eL��emY��\�K��:�\~���%�~�S�5��@5�@l9L����
Lw��G�D`��WRu�i���n�z8��}�j{�,A2���^�Ly������%���6�����> b��ÂU��}k5�����b�ޤ�,�Q���xF�y��K	I:K7^���}C@4�[<q�	�>\!�x�'������WT���5���V���[��uɈk�Ի`7ŚoV�ĭj�d�`sه�o�G��v\ٓ^i.W4��
%NH��b�<�.��VgX���=�g��n�Vg��(��X�T�u�Γ�'��Bw��'>m��eqi��/�	|��=����>
��aqŎ/��^���c�&W�R����$<0��@0<��)�c�T��^�U�/0�Wi��&��^���6�Ś�d[���w���J��f2s�{�ѡnj�+}{f��z��粽�R[��>�-��v=�| �+���B<�xI.�f�Q�Y5��;Y/��Or�5%�Q�ss�3�t��V���,���{���K�]�h:�.�Z��nf{��������X��mtݭ]\��.���]�8d��#�v�P��uF]q4�Vؗ(wh����_[S�U�����n��~{������k�}�/./�pL��fU��]�}]lBU=�:��p��l��uΩüH��lc����N
�'��|�Z�x��xϒZ<����;�/f���)�O']�!E���u�UO>ɇ�9�ϧLR��]k�8n��:���]W��<2�u?d4�ӡ���kp
�t&
�͛���U̵����wFC5r��F�W{�n<��e��a�m�ޤF}�����8��׍V�Z�[x��Y���~GX�tX��9V����S3y�.�A���7J!MН�����!�������+�Cr%OƱߓ�{P���ZT[���1P�R�$h*;���x�dD�����y��΀6��6���泰�5AZ3㖇��vA��pp�I��L�d��wVo*JE���&��-�}
�I꺶9}���2��Y���f���٨3����zwV��f:�,�+H�ǃ: 8e ���������v�R�2��̢;ۜ����ڭ������oO0lmIu���3�"P�[G�y��pb�c�<\=�^�����;��N�j�L�ࢪL�C*K,�eS�]��� R�0�:��/z�������{��U���V��K&`)YY&S�ߤ�a j#d��\S(N��m����$�m�h�PY]91�UIol�ɸ�ttX��� �/ )}�v�`�cc�]\�zf����x�k���x�{�=��1�,�j����dД�r�E�=�lv{���u5fz8�+�`V���}T�m��=��.��}�t3�5��ũ���.�G֦m+���Y��ӫ�]��[�2�m���y�l�\���Vq��J��^�\,�L�wՎ��n#���8Eh���دN�a"V�B�])q6���K�h'r���h���*i�nB���D���)D+���1d,���gD����ǆn��=^S}t����zN#�K�	u=J�]B΁�w��X ��V{[��Y�+WѕnfA�[�b3��1^Uh(m�^]�L����B����N٭��;@O�p� _OY�{f'�K��U�j٧�wCM��d*J�؝�K��#�G��{��oCϓHLiHH�L=Sl���y����Ӆ��.�z��f1^���ɍ���o�+ NДO��f�;.��SO�ꂽ�"-疳��ky[p�`Aeez�{�˔l�H��lЫ)к'��WW\�.E�i��\n���F�&����#��O����{6��<���y@���.���WN����=�m�,%�R#}3�Fm�[�6�kd7KNIs/Od2z��-�a�L�%(k'���P�n��]vG}��9���s:�&S�)V��K(�g�*�s��L�M���~8�,���ԕb�G=gd(�u��1�xm�'� ��8`yP��d�Em�O�f�jy[[<fQ�����;���|N*���b��z�p��^��GM�5�
X6�v�㓶�}@X-s� �8p,4������{���r�4�ػ��0��o����A�z�fkW�t�҆1)��X���:���.
ή����t�f�£Jvw5  +�ʃ%�^�W�}"�k�i��eV��z U# )�::;�h��f�h?k�� �ץzٳ^����O����}�[�+k�:����aқ�v�1!�ɥ��������m=��C� $˺V�ׄ��u�xa<'�~5%�\:�-�SS/���ټ�3�ש�M4<B�7�v��Ϧ�c�j���W*���w�s>�cI_d�4�����π��]�'���JNاYUz���s2��.J�y�ӟT�z4AP]�-t��z��!C�}s��b�ז�@L�6���U�2�YO��SO����5ZU�@Q��.�'}䟲�(Һ�=���M�X�m!�-�9�����|���cc�n�ޯjS��Vi�nY{��O��J��|+��l�R�Cd�	騉*yV�2��|H������ݵ�O8��-�ɖG*��Q�r��j���d��nK���]����7'�M=��?QT"ً֬��-����-;����%k��W/F�F�y����S�����&%���3��:�lOc^�]a'���=�վ���V�X�a�x���@Ǫj�%s�"�!m���zVⳌ?G�1����[��o�P##�KL�s+����R�hM!�w�e��ә�2t�pm�{v��m j*q\yIh8�H<�o�+׼�;S�¢���]ap|Ѡ�y�،ڽrI��۲N�2����nB���]I���Y�X�Sr֕F�O�\�2�6�Ь���@t�.{=69�k_�HD����$�.�@E�@l9L�ȱ@�U
Lw�]Dz�L�+={��جO��o�^_ue9��$��Ap�	��(;��1Ϭ<��dG��<�L��Z�d���2�w�ڽY:0c��x:��_u_x�/��JCK���;M�
̮�J%�&���[�=��7�fd�P����>�00 G	�C\�Z���*��߉>������2���>�7�#d�&��L��)Q^s%s��V�)
c��<���Yv��&�oL��t��ړ�a��#(N>�uu�羜L�س�I��p`u���-b5ԡV)�j+8:��ٱ�M��6�U���^�³M�6������3��z��k��{h��\r��W�PȶL���
g*�
K��x�R]�h:�.~�U��=�u�Z���iVs�����AcI���ϖ̔�Ic6�%��9����״NE�[r�E��%�y ѳ��&����W�r:�o��/��X�z����şb�
wx�<�l�d�r��zT�Q�zU6�����C��w.���w���\�����m��G�ب���A��L�v�5���V����T��o>fm��$�<���7%Ԡ6��ޫ�Qfѩ�R��\�Ot~1�MXz]���7���l�R�js�t�@��S��<z(y�ù���cr�����Mt\}�������r|���,��3\³��CuQ[�\d���?x��z��=��(��5�b�Ý���N\��Oj>�1r�䄯 ��h�c��43�=��gIp�¼�ܾ�ktY'���&���n�Q$�)�<KU7��9�]�[7L��s�m�L��&J�����jof�4��z������.wNf�ئs\[0nW7��֭�_]W@�إZ�S�O��fK�S��1�x{�C�H�MX�%��9�-7��{{��[�n�.�v�Mu�Tͳ���)���J�z(�M��.V����ޠ�^���X�ƙM���ڒ}���j�l[�Y��\��'.�q4<�x9�,��$nM�_�X�+���w��$vZ�H�n>�z�S���xyg��{ubÍ(�a��d �g>P	�I|���@�M���|| �vh�ub��d�S
��]�W���I��ُ�"\k�h��Z�Vɗk���K]���Z3���p��G��u+$���o�Z����]�H���-�3/%�{��1].Eӝr7C�q���}Ϣ��࠿'7��u�2w����1v
Ǔ��s}V�+&ǝu��V=��#��}ŵ�ۑ���!�����,)J�jBotCp�}&uGIVik��Gb�d�z�L�S��y�ᐅ���8�5~���cK��"k�a�m����wb����/�2�ۘ�83V	%�T�����>Ų㛎J1����f&��O��f��Qb��s�7�Q�T򡴟7��-�6�t�y��Ŵ��W9�$"��Q-��6���--ɚ�Ѷ���F����ۑռV0�wR���o {>}��4$f��b���9£۴+6���o�m��S�[(EZ4�dL�±C���U�x�6� �ƫ�ot)�u�V����R`EϥF:�6���m*ϠQh��Wo]�e�Fcyp
�o2r�_f�0�1�Gs�q�zy}݀]l*^}��xE-�v������N�+(G�^G���*\Z��W`d���u��"d���ȃN]��1�H�[.�������3xS��Se�w}��$ܜ�s�1���IGZ��I�sg�5�#,fԜ�
e�F�6L�AOc:�YL��:�T�!�����N�1&�]�,�9*��yy��^�X'{�x,I���y��{�_�ÅtŔ��i2��̣Ⴖ�*ڥjV�m�ҫmm��D�#,�J�l�"�R�
"�cj�KKbԴYKJ���m�+mK[JV�m
�F�Z���5�lPYU[h,bE���X����iR�[m������Ul�m[KmT���J��V���QeQ�*��V�B�km�h��YibTmj�icimjX��*�mZ�E��B�X�֬*�(֢U`ڵ��Q�JՌTh�Rڬ�kT�V��UF��KTT�յ-%хJ�ciD�i[���%)J����j�J�Z6QImU�յ���F�h�)Z�J��-��U�X�*��Kj�U-J��6�h��V��m��AKE-*
إ-(*�iaF�j��TZԣ��F�Z�)m-����m��F��U���%#U�Z��,�Um��R��(��J6�h�0jR�%�U�R�b�V����P�IKmJ�hڕD��*��E[l-A-Zį���>&nJ2ù�g�u��l;3��I��\'p�Nѩ��y�(�m�ڛJ�պJ�C3͏7���n=���s �����[�g�7�^o�}gQ�E�q_]:u���'C����4���ۏD�SǴn'�e�z:R�����qb*�S]J����w�7H����g;ù�=z3�X�Aθ��ө���c�U�
��dB�����L����f��[��<�zy)��5�f�T�0����0���eN
����M#�Q�!�H�;�ɑȤ����>�:Ɛ�M*~5���ͽ��Os��E����������M���̏z6=����8��*�\*�؝�dΩ�
ѕ/���<��eSޓC�e�wlt��j���^Ĭ�J-�
kx\%U�g����ιf��Dޞ�P׳�[��r���D}�����\F<PnO A (�����ye%O���
C��˅gЎ�����o�����e3o��̤����jO�$ x	��ve���m���0)^�J~Oyt��>�3��+�eW�\UI��eIe��,������j����
��tG�.qU��x7{i�4�;���Q�}�up�	@�j���֒2�Ӡ�� �W�J���ژ���H�a������MWٰ
��ˤ>\��o�Ƀ0��x1)IKrdb��+wt�QFi��֏(��|MSb�0��8���k����{5`�G��t�Ok����T�*�/�z��w���6��鬜�R^�nA�y�ق�<�=Y�/��0�֙����s >w �T�����9jK�÷k�v�g�\�Ǭ�~j�o���m�%/:�������x��pz���?���6sa�h��]�="1�k]��Uv}ܴl���`��J�d^u��LU�`I��5���.5OD��������f���[���XzrkPV�E��*x+�Bc�%��R^K��B�bi����.�����O;<x��|�UnfA����LW�Z
]�Qyw�3�n�%o�伎�qwo��qgH��P�	�w���ǶaU�Q�o�z�0�x�AQfU�͐����>�s�ݬ��{N��g׶� �.]��iHH���x�M�"���c=R���8_q�]�9�%���{_<�p��b�|J���p�8yf�<�m1���}/T�ND<��8/�q.���Ǎ��[7y�|EL�v��4*�
t �a�\�"�|�SO����ڊ��F�,h^m>0�$���a�c	�H�GU�fO��n�q�媧;�P+�x\�M�F,rbO�����b�un6|�1=nl�A�&�ğN$���j�ٱ�3"�i����Y|�+�����72,�ȗ��GH;%j)�v˭+w������O&3'�*�,�
���4��^^�]��GJ�m�����$x	c�/���B���BC�1@���� HΖY*��,oYg��-ۗ�/y��`���ժ_;��m��<�r,�OХZ2K(�9u4�OU���d��L%Kkچ�m�N��^{H�e��U��.���g�������
N�T�Em�f�5��7Z�o�uӼ�:	��r�{}IS�{-��a��� �# {αm�*�Rx4��������]���M�:�G�}�W|w�(���?�a��=f��w%Zqb��$�����8_Tq��/�ۯ�,�^�~��k>��*Zv�}<]�l�3!�Rnkկh��̡��['�n�;�냇 �'�u�C�2Z bb�#)o/<����}峢k���\���m�Gn��s2����o��[aWG�٠n����Y}f�IOg�oܳ������[�FS�� 3��b-S�b�}B�|�*�Zҗ 9�_���8.�\�`�g�שc����f�c�.����<�	�F�|㏚��zT���Ż��ͼ�4L�j1����p̀��u6�q�Ց�En��:\mEz)�	�2�f:k�U��a@3�)�m̼�Z��ɩ��c��Q�z�®V|�ϭ����n2�������E�ʌ=|��*��Ϳm�l���ό�\*��J�躁P���Y�ىJ�Y+���ꝄK��[%ԝ�(Ȼ��>���R�o�>w�e�\�zdZ�)�Ij��Q������O�ʇs�z˃J���#�+D���=�)������a��B��L#���5��7��N�yȷz~�&��|kUy~����z�Ӵ:;�S���T0R�UC��-9W�N���Sn'Ě7�ۋq�q�*��!�{N�ͷ.��/�hʠܼ��\�V2e�9��]=w��t���Q9��n1W�]��X��%v� ��� 6e��TX�p]��R�#�#�u�ԩ����ڏ�Ǜ¢�.^�1��@f���Y��^�z'V��h���@��u�gj�;�ܼ���5'ݢ���.�@�x�U�}�aoV�+b/����W�W��Kų���c��{ب��nk62�� ��Ϸ�tXC��H���!�Y�xe��`<���S�3����3ˬZ�1��,�%Xr�$�Ŭ�_����Д�O�fjSNX��w�'܁no�si���H�诲����fo�U�y��Z��L�+]J��rv���
����m��ծ�Wju"�{Yȍn�r��6%:u��v�=��W7�'\���s%r���}��+�kγ�ՠ��ds�u��w�,�=�K�[~FP��r��~{1�4�'�ѡnj����B}��F�v�y���kMj������L/�V�{�,PI�
�}OT`�T�3��s���\:yEo�LLz���+@c�;���7$>�A���.�-LL�����WAx�D��^�k� �Ss|�*�-��Xt��Z�,�4����iЭ�.P��l1������k��)l_z��	f�yՉU��c/�oGE��,g��;����*걉�sk'��̩���Y��>��@���p3/��S�׶$���Q�,��<$>��V0燹V�w�ɽ�3|=>Wb��$�8�z��T�0���0��N
��`���GN����yԇM�m{�7�Z�/k�`ڇ*��k�i���w����00����ȹ�#�4`fΩ��=�N��{��Y�hey#B�O��
�\*�؋��3*j��C���'�1��1I�=��7/���㞧9�i�h>��J�&�]�&(�
�3qX��9x��IG(b�iӽ�X%rWX���ǕJ�'k����b?-�k���c7�+T�qB��N��wf�ş���C��Z�L��k���;!��+�_<�:	;w[3�gtG\�{��\��(W�r�B�1p���g��c�g)f�f�8�^�ū�g=:?\pq��p��
�2�(7'�*Z��rˇ��>;�o^�ö�2�*8�k�y����#�)�"UIy?B����Օ.��S<�|�¾���|��{���8�]�='����9s>��IR\T���Ie�����S�)�όr���Y��;�B����]Ժ��e�W��;��{\�FK�BB����Ɛ9KkV�Z�G�1����3���2�[C�R�Ԙ�%�C�jn9�_�E�<�@�� �K�i��4n����eV��9��O+|��BFi[��\aL�!^�BS����'�0���L}2��Ŏ��=��0��ɍ�`Lt�J�d��Zr��`IК����{rs�ݷW��&}V����f�>���Qh�ϥ�a�^��O��}��o��ty���AM�QKӦ2�{e�:����ǇTߜ*��̃����f�Ub�+��Pv���Sg_鸣"0<�F�8kpK�6��V���ߑ�q8Ϲ����Ow�f����?P'���/r7}a��9t���+S"Ƣ;Dmۚ�7B�M��3e3g��{B���"b>� C���ۃ�6�?�&ﲍY�;���D;X0����FM�?fa)4��-�;Ć�꧶aP�53�bz{j0�x�L�ƪ��t\�4H��㡆��'M��Y�H<��������Sl���y����p8�x����6nZ�w�6�{�2�ւ+F|K&Pa�Vo��m˞=��PW�9�8��8R�>)(���j��a�7�g�z�ã�9�b��k:�&&5��eSMM9W��OWKky��x��4wN�\*Ny�:�z)㞞Lf}S�L2nﮝǴ+*xg�A;�N&�{��3����x�ek���i���Zs�.a�����\�#�H�7�`���si)����ϩ����+,υhw=p��|�9�x1��E�)��J�eIe��N9��g�n/�_�U���$���n��`��
�X�(z�3��Y'��ۡ�%�[Bin�Ǘ#��d;ѓ������d���-yh��낑q9-0��;�o�,)���M�+8�&�1>�d	]�l ���媙�GƟQ�3�U����iU{ګ�-�a�����0�4�����Ѿ��x�É:��٪����t$���&Z��_�����(<ƦA;{�.ac���K�8V�n+� ��S@G�Ao��;�lc��L���z�,�&��+9l=��M^��~�܉/c^[ɯ>�t�{=}j����D��zX�yyT�Z9�o�lzg��+��g1�y=N{k�~��8Jŕ��(`��&NM��v�8*��Y��Ƈ0d��U֞]�=݉B�"}U|�?�{'P�x�W�R�[�>]�*Ȟ��l*��� ��}�J���{���z�ۗ���K�)y`.sV��#>z�@^�*�ڮ�-8}T p��4e:G��{m�"չ���Y���,Ϭ������#��K��
_W��1U�k-eG�ak;�2Zv
�����"�A��t�B���CŞ�&����ُ�����Gl೯*[��]��>8��#�H�
��@�@]83ٔ�}�ë(!e�>~z� ��Y�1�	�y���kF,p� p�CocB�ê��y6Oq畕�
��)�O�~.�Gt���簨`�}S2�S��@���:W����J�w��&U�d��^�[�Tf���Q(5�TX�Sr֞�sXʙs���LW�*��S�)���7�)�X���iqT�G
��y�@9%�n�ضpT���<}�k�H��Y�d[�wy�J��妻�-(��V�����\%]��Bt��
u����!�Vd�B�i��s�8�^�a}[�����||H��ԍ`{��j����*�L	V�����j���a�X��E�\��KM�բ���ɿz�����QQ�u�j���U��|��W��}a���DL�#���:��}�c��s�����v*�5=�}���q�x�d�<J�u�j	(,�:{�L���1[9�Q+�<��ʨPtH-�9]��a��a�����3MK�2L���ti�pƴ���y��IL���r��2P��;� з5A����IB��!��7��]�9�8��-��u�����E-r�{)��L��t���s�Q
`u���%�5�a��Ej5��i_��ǧ��	���o�E���$��OT`��ip�罖~�����\x�fy3���.$�P5Dn{��7�r���M[/ۋ��I\pg;��Nj����J|�i����;�O\�ȏOE�rΣJ����У�����)���3G�Kn�ǌ�������;��2o/���ʲ8z��&Uޣ5³ҵ�Y�y�k�{��z�r��{�FXT�ҹ*qz�*sYt�������:�s�ʴ9����ܴ��ʧj���G���k��G�V^�<��U����O�=��N �5;꼩���u��k��Y������~���B�H�yܜ{�:'oF̝�˭�~��8�Sl�T�"�s�e�5<�(��t�cl;!`�߫h�6�)<d��ۣ�2��<�]���&�b���S�ªy�L>s9�8*b�D.�xG���j���Wڟ�2��;�Bh14�ƕ?�w���puS���=�d\ϑ���t�����C�5=��=`�UwR�F�֖L������؊�ɓ3��J��w�{9�^��+�gR�L>蟳�J�-
S�xr�P�n�P�`�r��3�ulr�9K0eM��@�`���$_X������-���6�4w���xz��q�LPl��F���U�ޭڌVn��R+4��������V��Ts(�%�4�
O�����Pj�bB��d]+��,�v����Q���~ףڮ)zf�ﻐ�2��Q&C���jS��AO�Ӝ3�o%`���ks�GgX��!��P*�{۞p��wDI_k����S���gI�1k��(S�:λG���>�߄���gҵxi��R�Ɏ��<Xڬ�X������ g�^��2��@_L�P����]Ԛ5r����m�����Z�H���#����3X�F��)ZI��z���H�E�<jL܇U��o�[0��x�دBev�mz��w���]^�&C5�96�Cu&�.
[X�S�X���3���3o�i���'d��\.Ԃ��W�K���A��\�:3�ր�n 2RS]��L����޹���k8�B�M�U@�\,�b��:���W��VVwM������԰:�Ɯ��Wl�WH��fl�>wpwd�G�Ot'7z�����14�m������wB+���%b��/N��#��ypz��'�в��Ƅ�d�|�ܓyBsܜ�$x�#�e���S�NO+�F�Ut^�ҕ��+ܾWR�-c�� >�E�٫@V�-#�:A�2��\���5�t��4�WM����W���˥;7:|x�:[�}�Ĕ^�fﱠ�۾4�ۯ:o�[����/<ּ��"���M4��ӌc˻��*|C�#u�ę��o(B���;k�wZ=.�zZ��L�]�vh��Iu3`l�M��J���X�@�}#�R�G�;=�g����0r�����e�����	�w�'}n��ĭ�]n�����4���L�cl-��빨�Z��P���ٱhN��B�BN!1��l�u-D)o]��U����c�5g.�\j�M���6�Gj�&_�� ����]��`�eY+�� ����>�'���6�cT���f��M�,���bÁܡi�p�Uf�c�_<	K�ce�$�����OB���<�t��]"L��n�S�4��X6���o�1�B�9Z�p��o3�jI0	�|Ӝqt�{�X�@G���)X�����Fv,��C~	�dQ�ڭ�G}��P�w0]GD�d���{p��w��j4�<�⑮�n�#�T��v]�^Bn�D��@����L�RB.�uDE����7]eIԤϦ�w9C��Q!2��n�|l7K	�c�g��:��71>�D�yڱc���4\��Վ�w�^�k�;Y����Id������J<l��ڽ��y���c{L�/s�tf�e謁nyK�]2;�L���4C��a����қ�d�O6y≌��H��G�Իv�lx�=��u����z���I�s>=�s�$:���=��:�Yy9�d�G*�<�7;p��݇:ζ�ٮ,��:�b��h$]Y��Kf�!-���ț.#�j슘��E�׏+�oN��J�U�؉�c�X2�����"��x�xs"�ϥ`��J�(�,���{���}4�Z��RCw�҆T� Yͻ=\��֞��.�P�.���8�Mrc��RRt&�<v�z 'zk��;��%�~r����� �?V�{˽�N�#rO�k��J��ek�6�&��R�A�q"E�+q��L��Z=M��<�\e=�]f:B����
[�n��/&Y��aKLO��Dp��ߥ%g�^��	�r�vx^��l�¤���m]�Em��b
Z�*J2��J���V�P�(m�EiQ�Ѫ%TR�U+�R��U�YF�����imD�DF�h���B�ؕ
��h��(�ڍ[UJZ�TK`�бam����m*)jU��X�6�F�j�V�R��)IUmjJ�X����j���bVƍ�me�ŪR�ҫQ�-�[��"�)mm�*�h�**�kU�֪[j%���J�aR�-�U��)DYm*�X��U�[[eE(�R����-���Z��(�F�XVV%���QFլ��,��[e��2����b��m�YR�T�V��ʋiIJZ�E�Z���ֲ6Ԭ*��V��X��#b�ciZ���#h�U`�F�TX(�V��U���F�[E���T�Dm-��
�2�bڭ�%�(�[E�B�R���dXĕ�"6،��
4+�>$ ��u�M̻�8�8C�ڤ�O���׶�zb�\�Xv�:g�U�'o5{��'��763ԙ�w*�2M��̤0�[��M1�w_�ج���U2���#���p;�=��}�2�֣!�o,���w$��Ť���t�z�8�;>���7�MI�����a��{�>�	��_��R�.���%n�o��o?&���oP�i�˫�bw�����f�k�+�E��*x_��A��fz��N���7�5�^y&W�]]L]AWz�0�5󄸔����7�X�����P�����k���Jv�v5�wp���Й˻�e(��� 
��C`�=�
�q��L����o�#���Wc���c5�J�N�3�փϬ��$}M)	S���ʛdD�;�a��.R��~��ͺ-I'MV��U�#ڧt�jch��A¯�8�7��+h��ME4��z��>���oS�鮟�E�_���|�c5�eL�54�
�)к'��Uuu�b�Xǘ��ܲا���/zБ�ly��jxe+��9��=�OE<s�<�̩�
�띐������GGJ�=��s�ȵ��t���������=��塞�O��-9R\��b����LD:�%�;��)�GW3[Js#6�b�0WՠA���D	ժ�̼����Jw�g[1�R��A_k��R� 2'�����	��*!<��b��+vm
�"c�6w�͔
�]�y�����-w�R���M�7&�jЇ-�����i�K��-Ⱥ�^����Xg2��c�����
U�*K(�9u4���k{��A�V�f9�	~=����2��_]�zP�3�gt�O!I��Zݖ�����=9~�Ez���]tn�J�d�U�}e�/-��pU"�k��g�|�)�^y������Y�������� ed�[ *�`y<�^��EN��"=���xV�+k��@���ug}�k���޾=:�h*��@�8�P�zOK����-�Ҷ�Ay�.Y�n>���/_vc51�����e^�d=L�e�{麘�0h��W~�'�y�]E`�O6z9���9.؄��l'�̔<��T��]U��F�W��[atz���{#�=���MoSb�0x��82��A�`z��FS�� 2�ؙn,��f)����1��Ix��ˍ����묔�>.�h�e}g�̫����{��n3��'&�+�!����fvn�79,�5�k]���u�\o��Q��1;���K�:.�B��Uf�f|���e���0%f�mj���m�u�e������-�E�̂wa�!�r0��L�;��*X�a�l�}�M��@|Ok���CP�tn������0�j����F�a�&!�@zr�e�P�u$C�6E�j�闵��mb��;,�!�]X��*N9�qw�r�K�9i�>S�ͪ��W��w>8��#�TH�
����𦪈�pz���1��k��$��
��k�bo�v��yHDw����l8���B���vaR���`��)����ٻ��o�&
�OgD�PD[�T�{�ẩ��QO�%l=��mx�g��'k_0�w�W.��<��9���e�-A�y��.a�B��C]f��3<�w�m�һ3���]ES�u��d�`k~J]��k���q�#9�E�ֱ�~���i�e��]u����2��VI��/�_[�gԔ�yƘ�}a����LN��oGS��/�(p��6�>�[�2�j�b�T���{���껐Ԟ�q�6�/�����c|a���s~�L�x؂á� ���t@j��a��a��lO^��˼
-�Ύ��V����s|���دI3���1�o�HSմ6��(g�acOD�����}e�g5M�w	/�����|V��*��uw�xy��A�w��k����c'&����B��~�k�Ӳ���X�4eL�U�����G�&��=N�)�l�kL���]Z�M3]�7�yR�ŉ�R�\�H��a+̭8�z������v�˔�f��
>����⎖� ��d�����&$��7$�ِ�+��uL(Ӓ����������}�Yg�o�1Y����HG�/	�$+�O�lw.װ7��v��ؤ�ԇ�����mN`W������Oq��N�e	�"z�k��X=�������>�k�ɧ6���7����[5�E���x,�?�*��u
8�p;a���M���6���{�&�l3������=��&���/.*��|t\���yӏ�v�!K���;����+(���p�0��p�:��w3^�.��&8a_=O_vv�x��qZe����,ʻ�&+�]�m��ס�g�y�L>s9���)�5��Vބ����Ѿ�X��.�W�<Q�!���.�cH7wOk�'6�S���e��'���׼=������]�#�Ϩp��@�.�L��z�yulE]�ə��hʗ�V�P\/���Z�EK}����7J'��g�����(S��СGX�J��>��o�{����<I��K�ik�,-���Sy��ꗙ���70���B��������u��UU�.�8_�?̭kl�$l]�(�X�b�.]��k\�\RԤڡrW��܎y�<�ɁY���v$�V8Jr�B#v���g-g,��z����hp�t��5�	��[YS;SCa�V�Q�2�ێ�ՠ	�v$nٺS��o�������d�l����D]y�\�9�C��=Y�.gӬ3��DuIy8.ޞ��՟K�5TĄ�,�d4��d/��_Z�o:`[��I��+�Kn
��A�r�wL�J��ࢤ�t3�,����ܱ���kጤ����7~g�e�u���E��������`ʮ�*�\�EUH������G�7�w�ߏ+b]VF�J�Fϥj���N���U!�-W5���ߩ��R�lu��+�4�|��"�ǋ�wu��lV�69��M�8z3�uU�\aL��֣!�% �w����s�5��6�&�;���t#�j�ϸ�̘бف1�+�y����Hk���|�]�t�D�]C+�kxʽ�!w���ʚ��/���ߋ�ۇXE?_^q�1D��p��%]_`��z�0�_8U[��{�'����ݵ.���5�M�s����(���E�D�>1%���l�[h��:�,��+����U\�9-�p��Of���"�*deD�,'��w;h<���y��4�$gӅ��H�D�mt�^�M3�ے�����*�ZY�Ia�&k�ҧZ����_r��k��p���Z�f���}u��}1,f���a���װg�ޠR�ꧦ��[m�|C���X͈&��=�k��Ӵ�D��NRj�=�,�e����NFI�ga��,�xu��h?��y\����g�N�2���+h��E4�����́�cK����6"&z���ߕqM�c�!E�P�O��뉌�"��h$�����1����R�k��z��֊�9��==��O&3%�<�@-�@"�M_z���R��=���P�ֲ�zO��2\U��Z�4�P�-2�����0d�\c<-u>�͓�L��>�������� �'*co}p~|�9���>�*ѕ%�v�'�S�X3k���\�ǝM�Uމ�Q� N��q�'"e�R��doRgwDI_�19�	1S~�]�y=�L��Oj��X.�^ɖF�Nݨ� ����T��^[u�B�.,y�2�&Gvt/N�=��T�{٤�v�pl�� \ {��*�{lٮ�m,�����[�4�v���f���<����[��j�xx2�V�(��<#*IϺ *��ʠ������(^\s)u�+#��k9Ȼ�j���[�V�J�Y�V>������J
���ɺ��ڸ8p_q�K�b����A�py�]��+�i�#^d�,3�Q�ެ�<ڥ����x�)H�{����{j�o�y%*��q�Bi�����8�Obkdީ�G&!����h�P�6���6��o��1}����UU��M/��.s,���r�S�r�(���3ր�w�%(_�����WC�V�e{�\,�<����Q�+5q{ó�(@����4v��T��e��X�1y`.�0��FU=\ *�ؙ�����~����T�������x47�QY�<6��..��}>^z��-�w����IY�
|��c�of��i�e���2���nL��9��:�[�ti)���~��c;�}V��}1⨆)�hem�֔^2�l�e{�����")�Z �w�����b$t�#GQ�r����`�a����a�%�>ӯ0Wa��U�c'��7Ӱ�T�<�2e�z�Na��D,	E��ǥ��E��,�P60:�F�r��j*�1���^���S7�a�/�]�^��yWr>S3��<��b�����&���WlFr�W��S�t���Jg�-ܵ��}7��+5�}�c]�d4�f���t���BV�#�.^򒃗j�� 6e�ͮ��E�5@(̞���g�}�e�5��e�pR�e]EO&�X�%}n�E�A˵{�0�����z!���]� ����ש���Uo_w�1!:�~j^wh]mQ!൸(���4!:&�9F�����:_JV��h�N(�u��d������%�쵮.)',�r�@T��
�sbf�Ӆ�ҭN�����RJ���o�ӗ�]�B���8�&m��9s�-��z��dt���Ci�2�������b�O �������Q��롘&;iv�>�q�ۼ5+7�<��|+;��{�<��ϪRzNWD����qi��e?q�W�{ޒ3�x^L�
���^�g	�S�����r�U�2P��L,iΘ��צ���g�v�O����Omp�0V.�`��w�e���̂nr�2�g»\�^�{1�}� ��[d�&��p��0=T��{K�蕖����V�X�����0�"U;x=�f��Z�4��h�{"����t�T�t�����C�z��^�Ӥ�H�V�:����@;Qݿf?T�k��Ln۳�n�t����EOMMw7m��z�ȏ�Z���^.뎍p)_����<k9�У��ЕSE��/C��`�qՉ^�v2Ᵹdhtp/t�Uʛ��g�ꍒ�e�(W��~b�9Sp�:�ʧqs5����c�,ؗ����%�����F=�*��LWb�rM��d3�i0���0�����tH�~�Z=2'�(�=X&�g�'��\��>�e*�.��̂��7�WJ�Z����r�����Z���w����{u�v�2m���1s�,�X:��w��$�C4Ůat���hD����M���s��W͹�f��NK|z�eת��ח$t�$:���h1�����;�soj�Y\��{%秧fƭ�v�pd�R#�ET T�f��&P�=l<��b.�d̪���
k��^Ю��ig\�<[|�o��O���УKBꞧdR��s
�OI�ۉ�kTD��.����MG}�EY�=�j9u��^f��3sP��#&(7>�@0����
�0;����4&'��e)�S5����O��eT�	�����9�B�K�i�v����ʗPlWbe��':���;���1�JWaUe��RہUf���!����Q%IpQ_I��eIe�D�$���_�H� O�ܿR��s��7�+Ac2���{���c�����$�qQ�ey�*�;{����WB}޼��r_��֍�J��G�K(1��)����dw�X�[�Ɨ�X�ԩ[c?b� {��{v�\��VW{<�����|}�k�xԉm�ӻK؛M���U��.����ԹxL.<Ǣ��Ki k���rͤ�6��G�2���PT�ѻ��l�|K������"�jì�����J��fB��r�U�1���j�Ҵ�[JS��L��n���U��vF�̭�Bq��hq����-��W�J��bq�m�D&f��7�=i�������ۙ�������Y�t��Am��s��U`�u�u����e^������3ӓZ���/j�}^7�����m�V��T^��o%4�Բ׻霡�X���C��}#8�u�[��{�'��3��&6߳����򹞬��&T�I����,�RX9w|&(�� =޲�0�T3�ON_*^��~Sޏ��v=��g�V��	�k�l�!<l2�H<�� �w��L�">��=>��:�t_�Տg��T��pN���uʍ���e�̳|+h�me�#�sl�s�=�aØ�����j��^N:��==8����F"F��hU��N��O3&��)��;
>���7�y�
�jh�Ϣ�i���A���s��{�觎L�O  ��(=�V{�9�����=���2��L��{L�E2��Z�4�5~;��0��Od/Fy�L�bs����k�W�Nį`�/�a*�
�?1�������3�x1��Y2��J�n��H����l7h��$�ｵ���O.��O\�d���C=]gwDIUg��(����xFd��#ut�J�Փ%b��gNqݒ,\K�,ݷ�f�}ݵ	�c���b��S'oL9Ar{�,U�#�:�ӧ�gb¶��;�U��|̺}�6�}�*f���-!����m��ɚ����ԑ��be�3&ԧA��b§�0��k�eu�F�n�Ʋ4�ɷvF��/�Ul)a��u���;z
}%f2:u����b$^��Y����ҕ���,>��ׄ����yx�}0�1��$Ahη��n�r��$q����;��n��ū��L���N�]I����6&:#@����綗؂�6=�����I�ei��K���&ޞ����>��\w��Ʒ�6�I2����<�{�4ls����>l�����}-�F�6��#P2�s̎�{��d������BT�8�Z�lm��p��:I/�(LnK�除��B��ŗ��|��v
���8�5ff���U�Ɵ�]��Mh�f�9�:�x0H�6�V��i7�;��aܣ�- ���G�����:���6�|�e,z+&�I��i��*��ā���SV�C�w���3��0�����a�L���>WAJ�d�ɺ�B�;4pd����ӕ.Š�e�n����aς(�f9�U[-���Ӌ�YlK����u��ڿ�ʸhjd�z�L�M�B)3h	��e�,�I`xwi	;�bZz�e�����I+�[��!��r�\��P6vk`G�/��;�v���(ܬÓ�p�F��s��{�K��W�4Oμ�8�T\�{-����cF�Z�����*��Մ,=��^�zn��@��!�/l�f���œ\��!��#r��V���ܼ��hط�1Yvu�=�\7~��sPH�}=��ꏴ�܀mR�5�"�u�Ce��T�]��o�qVï�kB�v��ޥ�Yp��y��}�A������V(��޾�*��e	ȏaLn�N�OzcEl�.f�݅�DKs
oꓺ��d~���ܰH�r��Ҫlc�����P��Q�F�κ�i����7Z�pp���LgNͤ���s)�L���vޓ},�:�w ia�}MT�5��;H��t�9��d�,'���v�]�v�Q�V���`�t�Gwu����{�9 k]���Ǵq�G�i�в%n|�n:X-U^���FI��A��<�S"�v�7-��v����ܵIE�/�����=x���ȱ�J�>^�|g�V�L�v<��bJK}��i:Ts(����O��3���Q1}�ܳc��[Mu�k�}>�Ss6�q4x�Tڲ���b�8��0�dY��lvn8rr}����k����3��&��9Y���Z��)uKW˓�fG�3��f�:��p3t��eL�p��U��SrS:Oq�K.��r�=��Q��]<����IG��oC-a�u�Kͭ�b�l�t���7;$�{��N�N��2��,��lt{�J�M@�h{��o��JE�"�\�R,�"�V�J��b�A��mJ��jQ�0�ZȉR���TX�V�-ZQ��U�d���ek �Q�Z��B��
ְm���
�XT����5������҉mFª[E�T%Q%��%�+F،�XV-e��m�QUED*-�V6Q1Em��­iX�X�Q-Z�ŁkT+DD�AJ�b���kT*6�DVЊ���T��D��l--J�5*(V�j[m�KdU���l*V�`����VXԨ(Q
���T����%B��+��IX-B�A-B�X�DJ¤PR�b�"�ڱE!Z�ڲ�ITb�J��T���Eb��bJ¬��Y+*E�l`*�EX�J��%`�6ʖ�*[(`ȉX((������ڈF�Db�AKJ[J��"E���J"�E�)R#ώ 0�˧�9�=�i�&�Mlk`��,�d�H�2�N�|��#fK��O+qw&ŵ�^�1�*jX:�O��8@r�\��f�I�q"2��#vU��Pڧ,x�x�<�"KBa0��u%R����~��f�K|�Sd<
r�	�%k�F@���`y�u=]�|i������F�t��ژ�;���cS��X���[~�=N��uܠF�Ǆd8������3�<�?u��J�yoX������Y�����;�V���YՏ��WY�	Obd������P����cs��^2=�._�����hwVdJ�p'�̔<��T��U�幙^E��н7L��z�S���.�FŊԣ�^^>*�>���+�ڧ�� e^���31��^�Ey�2j�73k!�\�h3iugh�߮�ղ���\\C��-�Gs�ek�$�k���m��L�ؠ�E�ʞ�nM����Ө�7F�Q)���~�c;2}z�h������#�����(t<J�-����<�D�Wq��s�}2��Q"8#�� |�=�+��rz.��y�²Q"���U3��Mn'�v�甄g6-��\:}���y(HǬ=���_�y�Mi}�wZX����ə��Zcf��R���MnW#����&�#�:�:�-�ot����f�8���J0�4J����w�4�f\)�����hjk�ݤ���Z��u��d7�ܨ�݅�Pl���J9�-��K�.F.Jj~6H{=O�9�c�Gt���¡�����A__M���JZ�/���r��g�.d���f��b3�E���
�;�6߾��Ͼ��`�p���b~I�����71=.�3H{��9S�tڳC>�d2U[��J��e��Ay���s���~�?��^X��2��u�+fU�O&������G���7�;b��ڹ���קmk~5�V�/+u�&UK�ϡ�� ���9r��Ҙꍉ� �6�޲��r���k׻��TI驹�!��fWt�%W�Hld(:��'*� 6����;y������H�Ln^
^���{�C�Kd�q�_I��u7�R��8��0��{=�7���.��voF�y��91��qC�~7��{-�{R�?�9nC��r��n�J*�L?y�y^(�v��@��l�Ӟ���]��m5�ǥU��И_�`��t_���j�a[�'����8���tZ�,T����$��C�A����¬������Ԭ�t�7o<�6���{n��%���;��L<��eD��ʛ�����[Gr��J&"�k�f�Z����[DWwD*��G��tؙ:�WyL��څs�;�+6�Ɩ*�p�8��}����]l�77Y��:[��7�=
�綋�vv�W�t)��zaRu���m��a�=Z�_�'���=5�Mjw^�d�z���OE�H�4�Kj�X��_�w��<�BkhW!��'h�ϯC}mN0z��^z�{����Y�-��tR�-��y�=�Ie�I�$�(��k��q��X�C�pu;���N^܄����U���d�y�������Tz�!�C�w|&U+�\��lf���f���]	Q=ku@{"�sy궳�GsE�"Z��W�ȜR5>.&���nf���9�t>5w�ՇyZ��]N�4.�X2|���a��� T��#CG({���%�Dע��%I��Y7�N�������>f3���$��<��e
wN�P�`�r��<v���,��n����j
o���>�f�����^f�������	
�2�(7'�*SkoݨziF���s���y�pg4��%O������u�r8��
f�T)>2cj�η&k��5�DW̧#��[˱��a^�b>�<\����bϻ�Q&C�3�w����Г�c6���~�(�l�-,lė�s��d���ugUޓX��q1�>���L�,�Z{i�yz��O�K-�fk2^'����d6��q]��9}��^��y�f<;W��g��޳7�6`[#��c���Y��w�����f�3O@�glEv��i^��ׯXto�u�gҵP*������K4Z>�� ����e�Zgc��6%��(�PӔ��Ng@�/�h-�����e
g�K(p�-���Q}�*k� {n8���{�6Uk�_y� �&'��~���掂��P��m;妹йg��9��O��أk���+�#�����N�.<ƈu7Un�}���vZ�J�nF��A������S\k֎O���V*�]��P��eb��.�85��������T���c��J1Œ^&�\ �~̖��P���^���5�U�����8�~퓟��Omv{˭L%��G\*��p�}���]�	� .����d6S�0�<w�Ʌ��������AlA�yE	J�!aa��.'f��'S��OWpY�R��vg ���W��u��zw��T��pd�}�>�.�Q�Z,�%�TN�2��~��K�T�=j��{\���ӢV���}pVt�E�O<��	ư'U.�*�Y��
���|�YnF=��Du��
e4V�e��2T���8
�M�f֗��ئ�H��a{j��ʷW�=�F�t�,����7'�d�OR4��~�Y]va�2�-fQU��[7�O�x�F/�m�Wس v1t	32;�s!a$yΘ�3:�oM�7���J�Ϊ?3�SMM>�z��֊�9��=U=��T�c2y�m�����|�Nc}|���>�dt+���8w8]1�w�;j���k4��Ct��0��.ý�{O�����/��횵w��O*��"���65���8?>A��_�d�v6����Q4f�Y�v�{�6��W�g�� [�'��TH5��/q�ҙK�M�Y�8����܁�,����T�_��(�	�*�%O;Ȓ��3�\��|�0}� �yC���4��f2��~a\���u���dR`�KʞZ���"�|�O��KOP׬���q��5�Ez�[]�ua��S=j�h����p=': *���pmff�kù>��pr�x�+�'Ԗ���sƝ�ILz��au媽3(x'�2r�n�;�Y���܇��#r�Dlڿ �^�N{.�Ne�J�����%�¥:�U��[����T�իt;���N}�� %c���=v�to(�7 ��@l�����F��� 8O+R��4����y�Y�[�sGE��Ǔg��=��s����Ι�B�e^_���V4�����L�WRXܔ�y#g�=<ʬ�{���ְdOMyw�*��Jf��}:�����z�Q��,��\|x����x��v��u,�<�"�A����\�OL��Ʒ�K�x�~���2������K����}��P��d	R��zg;g�&H��[d��9T�f��cj1{�#gML:�[6Y����߭��!��7�h)�(��C�}Cd������aT�c�]���w�c����n�:^�����l�7�����)��J�+��Mn'��a*�甄G{/���hU�/%B��FmYw{��ӯ`-^�%۲1P� �\�Mr�����/N���Os��wJnr�y{ދ1�xn�x�W�t�Vh_���U����WU��Sϩ�9���Y���|�}�^3o���X+s���������U�ѡ7�J�wYIAݷ@7�:�=3�F3{��k�|ei��r���)1�Գ�:e�J�U�j�5�Z��%�^L��`+��<��Nw[x�� ��8�	U:��ʭֈ�U/>�� H�zT�x���l���J@OU��3���gvV&e���RNO}��v����2�����W�'
��R�7�/zd��u��ZfN;Sw��Qn��5ct�D�4�����̓IO&���7;1��*m�^�K��gz���]Z�Q�}ٖ�,D̃�L �A��H��5,��݇he%eo6��ne�Z�y�_F�b9;_��Y�	G��rځ݌�dw!�k26��'tW֯�H_
;O.X=|�h��$����L|+���'+\�G�)A�?���B���Jn�0���-�������/{-�^��A_��'
ʞ�]�W���&g���!Q�OѾ�^X����c𕖱�~���c��\|	���R��-�ѐ�ޛ��u�ct���y"B����Ms;�����Or�:4����𤨱^6g�;℮W�w4׻�2�6:���=	��'U[���.��9�N�ܚ��U����PͯU�Yъ~��sIw��op�	���W]��{*ڲ�.�C[S��qW�M���yp{�����y��끮:��0J>�e]�/>�uʺ���%S�0Óp�瞸=�
�8�/�m�8�q�u�]��<�Z�|C����TՊ��6���u�p_T�g>s{��w�e�a�4Hs*pT�/�Z�i(����ß]"Ɛy�J����eJ�]=�>�i|����Ä��y�/��,@�U.�F���ez�yulL�a�ڗ�٧@��'L�`"���8��+H�%y=KLjXI8>]ɴ����&��m��|�Rā��q,�di�ҽ�Q�|'gumi���W�ڳ�t�u6 �ɪ!`��	"W �B���Z�6�i��DI���`B�#��@n����Ǌ��n3��}��W�AZ2_��)�2����KB�O�N��
�M�l$��3�x��]�܎�]^��"�`Ϧ�Y��*�
^���<<$+�Ɋ��ܯ�n��\�}#^�>� ��g�UV\1e%O���>��̨�Q
K�i��}RC���k�X��9���ַ���c}��bu�B�����K�s��!�訓�\v�[	X���ּ���j�x�v��<$ĠxN�`V!��({���zxj0�c�Ȇ���-̹N'���hl�R�j���o���r�����%xBdU�}4�ش�>2'w9��}~�tLz��8`������V�C�_{�L��>=��C�*|C���kO����2���F���Z�C���W�r���c�����n�HLv���j­)�"����g�zz����C���]iڬU_`I��[�KS-��������=�(��;��a�;�w���,Ap=z�c=>J%VJ���N��Yfk�
��3 �����i�펽p���u�W]��pi�2"���2�˕^U�yU��w�f�p�ҹ�>��7���z��Ƹ����w�d�f�h֫Q��Q���*jǼ��(���eN
j�
���A_��4�i�o7mfE|�Е�uM�G���q%��bkff�t�f�
U�eN�gn��Q}��Wz�l�V�:��L�ͽ��^�ԃ(�§T؃U�{I����M x�U�����(�j��v5�<s[1�S=��'yL���u?v���Lk-_ݪwK��Ljb�����_vN��G�wFg�
ws�teE�ꗪ
��#�y��N5�e}쩣��7E_Ų�q!��<}=8-�x
������Z����4���7-W
��f��x秓}��{����<���� @�v� }�w��Ӆ}���3�d���Ե�i����i��^�r� �or�̻���Z���3����},�U]�]e
cw�.���t>�k�Q;s�jl3ۋ�f��FUs��ӗSOOU�$�K!����V��ؽ(z�6ߏl���~��E��1�F��&��:B���%�[AOe�72�g@����{��(
LW��8�i���.�W_�Vw�KU�p�� �s *��H-�:3���L��l�_�JM��|<�)�����W�(���2��I��<�XXU��we�[��Dr�8�,[I��b� �4���X��A�M�G�>7�y�ϺlB��K��C���s��Q��R�Иo�I��d�7�0[���"��mf��X�0��׫gBS���r��:yd4��U�ޜFw���UkR�
���2IΈ
Y��v��%G�wJ�}���J�.�~҉�&j�i|J�f�V>�j�>���E�S�yyg�Ք7�y�� ВͲ�U�ݻv�Y�{�a��P5����P��}
p����o
������ƣ���x�T��lx��o������ �6Fd5�G���`.�0l�"�	{b��{��s�7m� X���t�b�}����}~uqtq��+��'�Q���[6^
�3���9f�T.8�4	u.
����O�m��61{�>�Ui4��eK�c�x����I�Ltxp�Z��*�Cd�z.	��v�c�]���\�2�� ���Z�t��=��>y̯.��_(i(�OL��FӶ��S};�{��:�^��%:}a7�۫h��q��`v6}����2�ل/���B���<7�聩���/�ߦQ��-;��Y�7��Lձe̐�L_2��2�`Z�Ѡ��TN��*���U�Ukf���$��B��$	!I�`$�	%H@��B����$��H@��B���$�	'� �$���$ I?�B��IJ��$�$ I?�B��$ I?�B����$��	!I���$�@�$��1AY&SY0�� |E߀rY��=�ݐ?���a0��A�
���	J��T(I)"��JU �	�PQ@��� QQQ	��*�PQ%QN�Ҝc$TUQ�(�)��(*�
����	*���I) /R���*�Hd6 �:��c(H$SB�@�[`U�� ��k m�hQ6B�\P�m��M��CF��4�j
�R�p �� �    �    ۸   2�@1 M5�ʀ�3��7ph�;�
�֊�8 & :��5��݋�vR5�۠�
m@�5�U �UK� Π;5(d�ci
�b������T��3e
�*�
m�� �I,�UP�R�Ui�)i��@�6�)JP p�T�")�
��T%	����Ĉ�6�fPj�I
J����M0�� R6�����T��p ۊQ!DR(�0�
��(� �� ���0(A)U6� \�C�"%-�*ɂ2`�&�P6*Zª�� � P �lU)SQ �`�  4�S�)I*4��@ �9�&L�0�&&��!�0# �?�$���=	��`�L���(��hj0M#MF&�4�C�A�	4��J���b0i�Li�����OMk��4kN��$/N�Re'T��4nA�C�ҩS� ���APT� U�&�>D�*�*+aI���~L��Ƈ��3C��� �d�YQV%`��
����	"����0N�U�SKX�Wwe�~Y ��׈��T(���W��0;`k��N5	J�sK�
�GĿ�������Ui*���Y���̺��(��Oci>:V����x�����He�i��r�E���;CB�K��'�ꖦ�onB7J�Jå�+GF��n�U�7��\���ȡ���"Ըe����p��JH/���QI�J�w�l��.��n��^�e�V���pP���4j"f<І�KS
ᛴo�Kr�0y
�����;���].�8X�W�j�&�e+�D$q�+��{���.���=��߬V��Y�M[�5b�&�=f���4ݚ�N��k7FC՚pMkY�ôһ�n��8�8M�w��>L�z����/p!Ɲ>��a^n���6JEh����j���K����n�Q�2��&�qx���a�j��e�m��f��em��V�m���z��E��׊�Z�(�DEP��I�Eݳ���4G��cZQ�8�����}���Ic
��n�����E��ą����v�RLl�ks�n���4fiөQE�5�&n���^S�\Z�ګWn��-��F�#BZ-�e��ϛ���-e^��5���~H�3V�n�v��u{WLSZ�U�Ԡٴ�y�1K-�c���mg:��F����$ܥ��
&��+���I�5��.�G^]�j�Y���Q4^ ��/f�UV�a��P�*!�r��)$#e��Z{(ڛ1E.��J�W�c5�j|�7���bF&�b�kb�n�Db�&�:��w6��%2D*�ʏZ��Ƶ57qL��SY$�N���#B�pӣy���Ś�����\�vK��U�Ys1b(nVmf��4���M ��^�9���c5}W��::�ɻ�aK�	8iH�:M��$���Lk����q���զ���	�����u_5��/2Ν���u��j�T�M��T��XB��{Yw�v�U��;��$
a���워�X4��d��y"lX����8�wQ��ʹe	6���L��Z����<:�naa�Q�t$��D��l��YN�����)�F[ׯMƘ���E#�����wc!�5��m��jfnC�v��	�::�ʶfK�C��;J��<[Tm�*��UIT�w�/�iثy(S�4-����S>[��T��V�<[gVe˄��衏UN\9�D�[:�p�	�lᮅ��uά���,]g'e�Ӯ���ݲ�'���Z��%[K�wL۽m�h�c�a�ؒ+���;��8V�
kCg:�f��']�k-�c�9g�V��t5i\/)�i����@k)��L��H�V��6����:��|*�5eP�w��cOt��T�kDV/,�sn�wn�G��3g�PV��~�Nm�X2�U��M�l�u�-]T�R�ce���J��oohR�'w%9�
�KS�[��]epye8q��2�1jànw�|��▻��VuU3>��Y�d�A������ٿP,9z�Ef�j���ح�	j����^��*����ZV5ŭAy���Ux��#���M�p7��s/M��q�Z�µ(&f�i���/�d��Q�i��{�en�U��i��]7}��/F`!��(_r� u���c4V��yY���)�$��5��������'3"�b1]0���e��E����Z�O>��e��	�ͱH�Vw14�QB�4mi���;�\Vj�Ak/
�7̥�P;uH�i��g7A;6{�,�:���9%�9�U� To�D+�c9.9m�t�:�������5v<�B�D�d���1�Y�4j��n���h����*P7t�
���:�0d4�������kkr�l�F}�KMKSE���Zr��0��� �"�v��g�����UM'��Ť3���hM�r�P4�4�t����9�Ţ���y���͢r�V��"�PH�	�2a7�Ɔl�ܬ]�e��z��Q�A%PT�s)\l�P�!G*�V�re��5�Ui�űtn�^����3�����75���j��U�0�B�ցMv����K�m�����W�]�ūwF��Ӽ��^b%���mł>#�:��	�����CFUfXlb9��w�p۩.�#t1n"T�D�[V�74"p��&���f���Xi��0Q7�V	{(�1Ռ�*�m����ޒ���'Wh)Q[Kv���4�+pݗ�Z��-�-�6Zb�*s3C,n�܁�T��k!{QҘ��ĸ2�!���iѫf��P�n��^0ERD�v	e��Ten�m�2�fҒB��ԪA:����{����YW�#�n�N�Dt� ���a!�v:i<��=�x7\�f��o�ޚߣ�V��'�d�S�f-L,$Z��WV��"�,��h#��7��V슴־+JM�n��,ms�坴Z���>?$闠�ot�/(���7�ƅ#H�k�V�;F�T�5�]ú^X"mJ��㧶��/��s�����ёӦ�ua2�m���m�w����0o����;a���lP���̆�т �����x�N�\����Z�,�K�ii�蹭	��/kۏtgƩ�qYm&���8�[�����79|������YDj�ofu�+M4)j���쥼9>���Cl�F��$��1�x�#��RK3^-�m��V�z��8>�Z��n�y�ݱFc5��ae��HY
�Vb�ya���$��4��Wq�݃�
�.m��7F�E���5�Ϋ?k�Z�p�+��ѽ�g#V�Kp�\�P�K�|�M���9aS��c�[�'ww��1K�6�*Jam\/h=2���M�f�E�cmc���]�iM��7�t۽;pSN��]!�֍T~S�[��e;�G^��֎�,��8�;�>@r@�W���Xof˶&<�/6;�h��*}X�d'�9����,LQW�FhV2K��CV��QR�M�#F��=YI�&�Z:�_Q����#�p��.��lwfS��Im��mޡ)�t�V17&�sX�}���J��.�	/ky}�P�8�4t�%̔����'�Y$��G2C��u�G/E��6Ŵ~t*VK�m0�Ym��Z^�b��^L��R,��KjV�[���h�y��%���:V��Y��p��W)�t�U8kJD��t.QT0U\�[��n ���	4l�N���Y	'[xY���5%�4m�����k�W�M����^�mU��L���������Tq�x����p+�K��6�ҮlF鄪��T������³3A�l=��+�����-;ya(�i�Q��9SB��j��e���);���-eC�V��{xt�h�D&P�Z��7%+2K#4��.i:h�8�4ҥ.&�'��^�sSfl��-�IG��*"�V���ٓ���2C�ƺ��lˑC{i
�ƛT,mۖ⽕Pd������5۠V%�p+����g$(��^%����u�f���꠯B��o1�&�q�A=�4�Ѽ���*f��gH6�J��K�U����)�t��Y%ĕ�@�\�ţ.��������[Ǌ*�4~�������y�!�s��U��A�^��4�t�! �4_�*���?��E<?H����[���.���J��5<U'ל��z���j�����nc���uf�s���,�;=U�wim-��b���l�qb{�j�b�ú�F�X�+F�`���0CA�3U��OvB۵8�x-][�c��Ka*2�2����W�0#v5��_l�ޱbd� ����F�<�
�SIVY��RzhU��pX��Qn�Jj0�!��s�f�L28����}�A�2��C�t�V�T����	�� ��\�'�myܛ��������X2���#kZ�:�[قVV�|�ٮm�A
����Q�(,��A�Փ����t,Պ���N'�]ԭ�'g!\��G2�G �g6�# ��[�U��ν.�f���J �p�Z/\57�U�·L��ȧ%���2��oo4P�ƾǻnAH���tಖn��UJ�	�Aɦ-�:*�΅]��Y���K]�2-Ɉ�W�2����f���R��(�MԄ�^��r��N�,B���T��9�3I�{��PeHj/�j�r��+���Dy���>U��/y���a�I�6/��H�&,`����jD1gm3���<�Z��f\���c��r�/MwT��k+I��𓅍���L|s�[�n�0����n�:r�J���\4��P��.��>.�3�\�!(����Y�c,�{0V�j�g���9\�'�x� ػ�Q-����DU��D#/�N�(r�2���oc<�upt��/N��ӯ��9�����z;�lme�%��۷0��^�X��^����_!��[��p��cD�vp`0�%fv�4�B�!�o���e0z��%O6���1jk�l�yxN�|$��fl�Hp�;D�0��q��u7�+�*��=�g"t�a��G���-۷�����:�5�Q��=A�:���'�S�I��Cq��%��QGvm����`i��ǆ��/;�]�����e7�Z����F�
G%�M��kFh�W�RZpS��T@Nu���3uc�@�qC/�i�������<��G�m��).�M��@�L�X:>�Z�o8mT�1l�R�wRY�,�%p�*�AW2v�ʸ8��5;^Q�5��i]k�K�&�r��tYZ0�-4y^UE��+��%l$:������w#>����#:���5�7b��q�"�RU��,��q]>���DڽB-�KO�����75SZ0u�&P��V]��17x�]�(�� ��z�7F� H���lV���b��<�È5`��o>N^�S��pgQ�p]n�5���N2�;����YՔ��f��ߛǆq{D��Ӷ��F��F�5�����8��Z�6�Czoh']��M��t���8!���fmnG�5�a��m�U՟Yo4���KWPKɘ�f�X�Nƪ�M�o%vY���� }�W9�n\���)k��z���@�%�r ����d9�vK+s]�8��z͛�ǡ��Q?$ury���ͻ�E�u}%u=L�;��WLj�:���u�6w^ew5�͉�N��?7�p;\Ȍ��@�|���u�/%���4�V�b�e��}Xa�,��6e��^������vM$n��]�X5�4�e���)N/���]�h����:֏f#G�MK�+OU��\̼�g��{MX��X&�j��W&�z*Sz���*}V��"����N+����j�� ��eq'�}[w��]��r��*�SZ'-��ܧF��b��f�m�V��eG#�WIC�\Xf�e�&���i�\����OE�|uÝ�z4��cEri��U"����]%�����Ii}!<��i�����3�Ht��w�[��9�@#Lv�N�0b��Ml?9�b�Oxo�`�L��˔���n�W�Z�L{�6t�2���)�]%uk(K8���U��h'[�!�v�k��3k�|5ˁb��0�S��z�Lgt�ox>
-�yϯ{&c�:'���F����/��t�t��7��G��1���;����G�Vw�k��"��u���֜�^ꗙ[�v��5�=%s��SF�ֳvg�Q0"��t��'vs}�@#���z�NڹI+�ҥ��=խ��a1u����5j�s���%*�;�%�u��H��F�n'�,�\w�U�Z��b'j%Vч;�~��J�.��B%.�Dd]CS�xy,����ƌ-��NwS�̆��e���c�#QZ�̠��s%f����ƕ��Teu��G �olN<����a%U��J�NbՔ�ΜSw�@Ջ�K��3���nK�IO�������q��U��#*kג���m�U2�j�z=2N8=���]�pi8��n0����H-ٽ����T륭�,	ZÀ���_H�^ތ��6�7�`�dR�n��!@��(�S��,�p*��Z
O)�b�K���qv�]dX���N���N#0-pI���EJdga�u���o;L�0�:��t�$���1����z�%�2�Fi�2i;�&���I�f�˖A��[N�'�dW+3u�+C�兟����P����&B��f��,�G8fX��ܫ��L�L�^��,ǭm��]�<�v�],E�˱4���FM�ˤ�e4�F��Z���F�iY�h���h�(�P�X��>��]tc;NHvmdjɳaX4���k��`�|L���.�S�#{l�׻ �u��\ߺ�R6���N����j�b���:�־�j�:���[OTe��4���Y�ݡĤ�'��s$Ti�뿎ê��,��J�{���� b��q)D�\ݏ������/���2D@`@��l���0��`v�an��:o>��A�%��J�i��P���T�-uu�������̾H��mZX��6�z��#����9�9���O.�n
C!ZGI��X����v�x�+5�خBs)j#;�N����j!��@���!�� �;[�j�xckngUr8g\�6�<�\��shY8�VT��o-h��Y;�ZL���ێ�#g9C:�!f�|,�^#�B��Ϣ�$���
�yi���a��pB�3q�Edɔ':Gw��7��l
�4ot��rz��n5E�6�u�xl<(l�i^V'An�x�*���b꿱;쌞������m��%�}M��x.VsZ��p�t���Q�+|(���%ٳspI1YKz�. ��w�Gq�^^��Y��N����DT��-�(�r'%�#�R���t�"8�n�!8���*e��rH�*F�m4�m��m��m��m��m��I$�I$�I$�He'h���-:��q�Z�.E"�I$�F�m��m��m��m��m��m��m��m��m��m��m��m�ӒH�rI$��:�*Wjݴ�7��|r%u�l��ī��*g��	]�j�+�V82C�2�VZ����Sߥ9�μ�Y{���sܻ�H�V��ļ�o�p��V��x�m�Ԅ�|~�c&\��O|��>��WXj�9��C&�X�>��32͊a%p��������o�}���9fg5ul�r�1��@Ef����VATU�|�*="j�\�����*(�A�G3v;hM�+Ѫ��i���vZ�Wn4�:H�;�2^�+�+2�
�� ����+H��T+�@���L��U�6��L�0\��Mv�A*:���0f����릒u`iW6��Ȱ�e�zH��}���a���t��vDFJ��}uIo:��PCF�\��Zuf�s���1A�\E6Q�hf%�u��B;�>}W��[0l��&T�9���n�˅�q���P՗ٵ�f�w
�\��_]�v�0mGE`�)���QަRھE[;/���m�)��J�]�:5�	��+��sx5��g]S7/Dt!.�'(�[(3:nK|И�!M�kh�ŴB]���\R�M���E^g�C��H7fk�	���#y�B�e�ݰ��S2+u���=�������h��v�p��:�{��LW(%�N�+���v��ټ��nQ=*rYo��tp���6k��Ǌ	f�&���P�0��F_@M�}�s�d|�WٹH��8n����q��`P�v�C$�:�qFQ�7���cxJn�eŏ�v;s�~�Bn���k���'΋�.ےS�7N���%qB�+{�Гx���xq��i�u���ƑԖt=QV�uW��ԕqX�8,���t;Ρ	\��O-,�GL���kB�r�C���8z��.]s@�5�!��e���Qb8p�x��l(w۟*4xh�� �EZ���:�)��Ő�w'u����]�s�Ԭ'��6��K�*IPN�aI�VOU'��u&���}�f����ɖ��83bNX�ؕӃ��&s6�K�aU�xSҳ�6�\�B�Ej��M]��\n��s����*�W�&є����}��NB~Ѫ�#����j�rwl{{�;am�5eхR��(�K�	5�9XOs2��(��m���'LT_r��bf9d���O)u]������h.}�B.���xd³-��K��/����c�����9��K+d�޳�%I��Yp�nv-�����u�{t��G"�C�,V�a�³���Iwl՝�������a-WvnY�f�@oQ���Rz emu��/dT�e=X�À���=��;r3�R�Y�H�\��H�{,���t���Mہe��-7���I��w�LV3��h��>���,���#�ߥ��o�z�׏�!'eI$�؁��H�{��:V�3_gj�j�=�TC�������M=̾Fj�M�õwO��հB�� �7�KY&v`�{LNl�;'Too�8ն��v.|�)�X�J��K���33*t�J���Z7�������.��j'���u��9���}e�8�A�MT�tܢO`��v$�#D��u�W�#�sa S��e�l��!P���d�AY�C�����{\/΃�mra��wk�����k2ok��j�ed�lC'm�D>q}ۛ�[����ή°<�l�;����P����Cһ�
���:���"�tޭ��tA�O]�C6���2[����R�N�ӝu״��{�ڃჶ�=v���Ͷ���,����S�E�]��ɼ �.<)��ur(38��"��m�V�0��=��b��Z�aW�죖���cuՇ��ձ���[�������QQ=ď��㒺Wg�W%��y��������[���|-��'\\����d��S��Y��i���
������v\��^��8�bSЕ���1�\�n�5ՂKudar�m�n�pV�����Q�\-d�E°Z�'�)\T���s7���Gw�RŮe;x�����wmq�#O��Y�S7�9�l8�O�����_��98�{����w-r��{n�p�����H@����D���h�Ve�2�u��&n���'���Z�nz�\�ɕĔW8�t��Tl����t�}g"�C ݔuW;��6��M���wm쳦S�j�E�d�2�+9/78�%AHfM�g˻��//7!�f5/l�c�.�2X���mwpCE+L^]�e�]J\���#��K_wT�����c�L�Z�P��{�8�9��M][x�n���rVٸ�QJ��s�{ƣ�5�o��{4�c7.��K�L{ksNq|�D:���oV��@����N]���{���Rݘ���������1!Pt|.�e��NN[�+,<C�7���y���j�P�5���	 2�Z ��[�Ð���F+tk�L�x;OX�6�xL�1��Ř�Ƴ� ��ϫDw�YBv4,��kp⣧VP�ˡ���x��Ֆ�������t���9/p��͓3@d��$]�-���$��ڝ���6�O�;}+�x��&}2�Sk ��P�]�J�\����4�H��E���pnJ]Lq�T۔�����Z����v�*�tz�A�'6{o�����N5�Bv�2(��\VZ9�!�q�LU&r4�mGr�K��CX(<��a�a֘�"88��ު�ݷ���-QYi7�۹swD�;6>Q�.p���껦��[����Js�X�>;�p���&��\6�8�@�P�uWn�F��ü��92���ˡ�v7�*R��R��m��!�t�m�,��(qB���������,R���PU�;hvL�P���	��J�yT�s���гS��lD޴2��]����s{�@QGN�Ù���׺T��E��+Nr,��u]V�źX%-\\��y�v	{���nط�<o4	��X��;�7����8:+�L��;�6�e�H*l+�h��9��7ג��NN,��t��c3E+��oN9uo%ܫՖSꕐ�8H�X%c�����ڌ\��νy��r��͎8��-v�#�z�R;�rgf<rSR�5�q�@osT]�P R?�A��+DTU1��m=�eN�i�e�]WOV\��wgD!�M�tE^��S�aZ�E���t�T{�����C0�hǪ���\/�pf7��d[�޲��k�Kf͋k�!�&&R�>v6�M�����e���ɤ�B����'n������V4ڽe��1lr7�ԡ��h����[�Y5���^�S�B=��-+-�c�|`j}�0n�=��gx����V��z�IB��6|�5x�OS�+��1i<C|�q�x�u�K�o����/��"k��]+�m^�s����r���%�jn���)��MPI�b�N2�p�-��@��B�@�tl���SX�*����L�$��w&�8���ʰuv(���ZU%�A
y�#���Or&Qu��(E:��ɲ�k�9ku�A$*�d����,sSE|a,S֊�B��l�G���%��rԋaݰ���}y��a�wS^88&V���Q��j�wL���(wIm�V��=�hVa蜴75���0�,�nA�B�-X{tH�c0f�r���4�Ѩ�Ŏɚ��������&Ƌ�rMt�����LJ`�W֪���0pZ��;7�Q�x�iu)t#pS:j��[*[�3��;�L���:��Dּ��lޤ���bIwٝj�t�
ͤ�X�T+���O��R��������� ���p0;I(���5�va�U�UwX<=�����$o@Y��.�|�S;%�5��93��k LW|"69��2�SzL���+"�l���M�Nj�S����)ټ&1��_6"�W9����V�|��7RRL�·mK�_i�ۗ�l��k��z_LuB�b%_jN��N����ݦ��I]���b�j��z�[�S��/_@�L4���ΨIʴ	�	��Ԝ������h�i�v:�J��Swo�I#f}}j���jK��X�f��Bx1X���#�Sj�T�aA�Q���JEH�8��O��tU�T�(�G��5vZ���zG)�El�`��%ӎ�呌�r�Г���pP��\�˸B�9$�H�HbOe�],�7�E޺��w5��R�>=�`��n�S)+kec���˅���2Xŋ<Hp�
,��eLC�@�N+P��%E�b�s1
֫��F���r�(���AC2�[x� �%��"��mf��eX��b��(�����j�@PUS�Ղ�貸��h*�4�RT��bVt�m�E
�i�Q��Ŋ+��Z��$�m��3MsV��QQ�
�*ER,q�˼6�3C ���{�Nu���<t}a�r��:�זHD
	M�&�ڙ��tG��N�0U�������C�
�R�����W<�8������g�c��f9^N�����'^��\�P�g&��kg�з{��jd��R�Y��"�����Q7'�ãk��蝮8�8���)-{��-=b$�����YB�s.k'�?졽�Ӌq�cP��y�+��Sc��oWb�X���\ߗ�����Rv�;&E���X�g�,�q��ǘ�6����m��� ��һ^;�{�V��3�y/n��ŕ9��)�W,Dp����T�@f��p�}���5K9K/+!��Vr�4���h�.6�t=��+�.ʏ3�4k�^p�	^�蔧{>(b�����p9B�Q��rPۂ���q��~+v/(�'8�N,y��Z�_vu���+=��^)yfv��>�p�pߗ�UN����.H^�t#�h_`æc�'M�b�ާ�{F҆ϛ��	�SО�>لG�j�k*�R�k�^V�O:�ǯ]�rD0�M�\�Q���������U�2���ł�M�0k�踈I�'
��"�{ԏ�>�R��z�F�/S�@
rn�X�]N��6N��pk0D������9�'ӫ��.�|=���)Z����"������c�T��m7�Ӏ�U�W�6��[�<�]��N��{�s6ts�<n�q��C}�,�#�*p��5|j������Ng��i-=/�u{�o��܆�I[��ru�c�2���g�gb��dv�z�#���mN����h��]r�_X�������up�n��eu��j�6���\v`��A�>��&�XzJ�Ko_�O-�L�q�j�
U�>��w7t-]
Og\X5b���8z�I��WI��j̭*��s��[�z�=2t+��N��K�<�[�V���F����y
�hۈ���?5/�Gmۯ=+t�Qy���۟*�X�S��\'#�m{��m�y[iߛ*���{���Bς�΋u���������rм�
?,�O�#ik��\�U�6u���/2\�Ґ���l��.�Ï1�B2�o�N�,���hf���2�g�fy�Y`d��ʶ����}�ϺL�+�:���g&>������b�-�.��>��*��@�a�높�_���v.�%����XN�6^@�d�U,ؚ�W�ӸH�C�&�b�TY�v��x>εt|���E�{�8rвO˗�a���m8���wb��ŝ?3g�]�\�ǈ�!�-(a�S=RW`�j���}�`��_s���#M�^ܖ���^�O��tHu�`>B�R|�F�\���)���u�۵}|�=�AOQ�ܯ�P����Ry9I��ug��6@�0�E��B���ί3S=��tC#H���Hd|ȧL�/�A�M䛻�V}�Lq$x�^/�/���A�*���c��|�W{�>����'L��'˻�n/�����t#��^�aǷ�ٻ��k9��qp)ݛuSp�Q7���#+r�V� u��Q�K4�I�wZ�f4�v�<~#�H�^(�C<�D#�f�]�َ��s,����z~�O��A���y��k��r�G����E�_��	�X͔��:ݝ����Խ�t^��0Л�i:p�i�d@~^ZCJb��{��z[CN�dg�d����:n�"���7���Ҹ�	z�D,���K�=p�ç�:7MU�"�ߐ�y�������0�*x=���$z���)�(�<�l���XEO0������V���}��nnz�(�߱qdKL]���C��k�Â��\�g׵���u_�xD,�>��q�9�-!�ߦ})�b��9��'QÓ�w�[��n뺀��z*�s�⽹�7��e����}�w.MUa�Tw�e^A�pU�f������ρʧjȥgAM\F{7�EX��N���^����!��F$6���i`����}���dp?iIB�x���E����W(�����f�b�Ĕ�@���Y���	���M`\]!��}H��Ֆ���������C��ZC�
�qӔ�U�s�{�����-@-ZY㸾��R�	D1��R{#��+r���x�(Z'�qx��͑�:q���x=��Y��J��!�ٕN����s6��o�t�ff=f�K	"���5�I�`����!ebg��Iz��a�4XAZ���/u�Šk���D{�_o��cEƅ5`T"��I���^��NY}����!w�y���G|i�&����q��b8�A��2�ųpB�����}Y�(���?����^4~�>����W�<Y�!��l��"8��|���������xeW�|���������~�x�m�>�p��ԯg������c��Z���:h�DjK{��ه~"���=_g�/��a	��oq罝�����f�	}�/��,��-�#�N��!�4��ɈDF}.��r�e�n�/�w]��o����sf�{s�r��~���<��a�a.Cnh��]���ޯ����!<��n��\~ii<.�{ҷ}H�!��}��!�r�@���QѸ{xߺ��6O�&v�&cTm��.���
�Kn�l������j�1�+���ql��C�r�\���-��澇kL�-`�>œ�88��5���??���������a�W����w]������"F;M��ϗ�"���������-'-�������@�hCwRc���[�7N�\�s�Dd@M�� ��1��>$���<9T/G�w}�ѧ���1�A��j�PAf���oǇ���\=�>�������e#H���Ö6����/��:�<y������ۣ��Y�C�������{�_b"���Z�G�k�CG�uoIY����z�B�ƁʷS�}?ľ'k�{b��#_}ǉ#?d3�!�z�'�P���I$��UչІ�CH>y{�.]�j���Un�Gj�N��|{�{��ÁU�a9ecz��4:�m���]�l��_amY�k
/,Æ�j��3�j8�۩��p�-]xe���CU�c��*��0�N��wt4t�ϘcQ#L>>?qG���Y�=����&V�Dn!�l�cPt�� �����a���7~��tf{۰I�HG�"�#e<(�C���	G���z���}z4xEE��/����b_3�,X]��tx�{�s���.������/�����׉D�w�����!�X���c�x���k���HB��G��}���W ��C��3�d���4�,���o��_�$o��Hy�Th!E���ݿ���5�O�����#��	��-�_�u �_��'ԧ�%�r-��]$�ݤ��Y�t.t��A���^��Sl�}j�*9+VRG7H��`s�^c�8������V䋒����A]r��R�v1M
ʼʝ3�2�.�ƩW-)fCծ��aJ�j�GȨ2�c�Q���ױ�Q.����lgo$�b���T�%յ���[oZЬ����֌B�I�j{�l,��y�,YZ���=��'����b�P��w�*�2�mW\ஂ¹�û�/�od�oV46M_b���B�C�����̌e�v�k�}�P}�T�;0��s�.V�0��_DMA�8��<��8��T5�/��$n�]*�b�oYP����\��Y;@�;�E����6�K�BqmI��q*�u��9�W�~��_�%D�����~ҡ��(�Fa��kmT+C����c5�b8^Ǎ��r�&���:���됉����겴fG.%� ���Tr�����J�@��Z�C��γϖ�R73,V�[�bT��n@ �6���j�{�bwn�fg6A���RT�O��6t��ɔ�&��Z�IO�uyʤ���y��E��u� ��å,��N��5��V�5&����pyS��Ҽ��*�+�B���o8��UX�'e�6�G⚢�:�^R;3/�՛+xںW�4F)&m�&��Ħ��ݦT�\`�zڙY��R7P��Ae��If���CygV�4#x�x�$rI$�rI$�7��;��<������Z��"�,��Y�U��KmA-���2ڢ��F�"�d�B��+�E��c�W�*M�dU+
��m����]0������l�ȕ���kIPZ��X�m**�jQB��;�0-�<`T�)1�%�bE1�VAM$�SO9�4�q0�Y��QaRVT��TPUeM2�R"Ը�MG([k%`c�dQ�&+�b���sw�?�z$$���s�u��Ҕ��)�y7�O�^r/�es��ϳ�}�ayOM�u	�_����b|�z��ɹ��z-"���"��!��#��(�R5FG=�~P���ZX��Pf0��$<_�����ՁO���s_qz�4,����"��$���O��_���S奝7�/���8h���W�k�^o�´���">q��3퀽Ϗ�&�SV�:�����#���4t���O��\��@�ٯ�u{�y~ȸ�����/��`\h�:��"��=t򯫾Q�^�,��W��lad����~�^�Y�S&�d
���Ӹ�Z�R�	D_��Y�:W��U�h�Rߨ�e��탢�y����t=�����E�g,	LYתz|�I�鐧i���a�9���]����*wz�j{�~��8e!�<d��/��0�n�����}n���Yx�bl�!*/��f�1|��E�+��	ʾcG"Y�VIK�k�I瀰ڭ���,����?M�j�do��g�W��{�����9�6V���Wܛ��\YB�(�}[�����˒��_[B����0�͐�^�A����Y���h��;���by����,�|~#�Z]=��ݫ���8=a�*'�=�t���L�Y���Ve���yX���!X����1<�����F�z�<L���S�v_� �>/V����*b��/�Y�8��7����o�t����b�/o^���0K���#O����55��	�߱��S`������"b=��UT���������yZ_x�gH\�ꪥzϷے��Z��D���#�����UA�P�K�����_�����By��7T������t۽��Y����b�?x��R�t��֐�!�zg��Ʉ{�`&�Z�='ޞ�_b Y�+�]���y�׽�����!�i&r������,�?����x���z~�d-=!
.BFNzh����t����_U==�ő� FF%��<I�M
�
�kG��/a���?ma�$�5}D�B�������vB=�c�+�{<
�s�t.���c�j��/��q�Y��%%��V4}�Ou��?�L������2���Y�X_�R���BT�����A���vQwJ�Az7d���+2=�#���껼l��h�g���V_ �\����1�Qv�i[�_�#g��9 ,�G���^4~�_lʨHG��^������Q|$=|�O�?���Nr]��~͟�j���MW������H�W����]
�A#�)7�<���u<�ج��;�p�i���= ��?[�{�YäB!���<5�H�@?CB��+k�M]�x������#q���_��c�Ŝ�����������,":`[v/+Λـ�{����),_��J�	����H��<(�B����}�Ş���끇���/�TaR_3�'����r�t_��>�2��v�T��"]����M<K��$\�X:b��zkU�u��|�G&e���W����������������>�t�ea���n�a~XFE���&�k�e{$�b�چMP�<G5a�_H���*��U�{��A2��C���<]��>�G�#OԊsk�&�7�}�{ȑ贂E�FӜ��-���oA�d���>?y/�>7K�������_���9ql�{���L=^"��YG�Ai$X�xC�|��:w]ơ������KH�_z����'�F�*\�~�v��z�~�7=�u�mX�(�y�`�!b����v�m{#x��*՞x��V����g�MZ�ou����K-Xh'��>"��1!�l�|�s��m�o	#��߻��e����lo&x�ۙC[
����Xz��4A
�Ƴ�/���y+�x/�s*���n�(a}g�N�fs�������'�t`��{J3��O�>��o&j��ߗ�92�^n�ug�a�y�}uO&���x�;)�A�7w)=�hm|V�Ȳ�,O��l�}��6#/w	ٕ�Wc9a�D��(��Z=�8�T�����F?%�t�ߥ��ܾ�t����j��F�-������Z~&��#�7�Q4~�l+[ɘ5|�Efg���|���;儑��g�?,�?j����T����D�26� ����Q�������Q+�Oj�s��/'@H��u=c�x-B�44�/����ݸ���Uy}܆��e�9���+���(����^���:[�S�<�5|sOuc1�������8��T������'۾��/��h{���M�u_m,5����a��X�j�=����d*����a��Yh��1lq�diӀ�??��v�7����g}�4�8G�?�,!��v!�o��G�4������>���Dq��&��N8�����8~�#��sw2��8l���}�!SgM�5D;G������ƖEe�j�� �Ab>V�� U[���@|S _A����Y��n媿�/�ڨ��>N�}���fl3�,�;ʍ��>_h�fئ,�b]{�3��|�/�-�Hg��xi��ƞ@s�[�PbP���
��{�Uɑ���y��"��;B��W��~�^�>T�5�q�}9����/Y�y4`ư��yq��T
�*�{�ݽ����B����2�Y�xL��a��Ȉ���N�ӗ���.�1F�L��2M��wz��u�'��}s�v���^��	w��]�CP��1��M�y�x�[�޼�B��w9��:F����Qa������8�2!G�/���bbz���?f}���A9U�5��a`D3�ؾ�(�#F-5�ͬ�]���y��"����Y�ۣ��=�wi��ﲠ��Y�	H��Q~΂Z��U�yY+v�O�ы#�apH{�,C@���^���~[�k���Z�b�X� b�^$������A]=�+�#o��!��8h��y���+;:`����ܴ�"��S�S����<�%q�NU����l����̓�u�\:��},jr�-͇����������nu����-ǜ��4�y&,����vj�?��� �����G�&��!d�g��K���O.��6�z�p^@Y�<��_y0;�d������-�]�|~������$��
6&�<���%Px�JkoHs,{̊��o}_(��F~g����4[�S.��x�}k��<���daG�A��K=B���e�}GܾA��h7Q����8��}�s�SB'���~�����*L��d�8ա��@a`����{�=Xm�$(��F���Bx��uo�P��{o{)��ѳ��?(�����7�B+��|��-��ʡ��Ɲ"RQ���H��!�1/Ù|�*�3��WĄ3U�Y�2�U�.����kDU����yU\���}��\���*��b�ސY}�������}_}�M�/B���Y^�h.���?;UH�?������ۏ���?3�#��|���!B��s�~?����|~��a�O���w��lu��}�k�"'vzB��+H�U�m����*-##c]�2��=Y�<���t�#���,r�/�/�-90��C}���R�v���
��w���pw�|��l��L��Pp�C��������0�¹ZCۭ��n��cO���@㦎�������yY���E�q}��:|}Hhx�B֗��"��3H�nu��5Ãh�\^!��B��T��B}ky2>~�>>�	�8�^��C�S8�j+N����n�R<�b�/��!0Ω|ES�i�VNWyb��9#u�vH��}#�kF�}��w��IGn̄邧=�����V䛏;&�=����f��g�5-*q[�v���p����V7Rdm���+�9M��Z����/v��ڲ��+4	�V�)���ɵTDI�������E�*��m�s�v�E7�K-��|i���u��נ��n���0���1��u+�9�LΤ�d�􉝛P�ܛf<��K����;��^f\G7�����mУ�c�K���nZ2���E_2km5Y*aW�L[g79�Kw{v�.�=' j��wf�i@ިf5w](�3{��zΖ+��<��3o��Kn�Ȥ��x�sF'S��S�{ܭ�߳
�:���8�ɻZv��1�;��D��g(�ˠ�3�k%���� F����\)3wiU]i�9��y.̋��\qL3toK˃�G��j��ʃdY�5	N#{���̄.;�uy�F��f��3��6M�8��u}�V�+�YGz&��f��E��4�<�>̭�5Ɇ��w�l�F7���:m=ON�g�U/8���O{w:>�Tf��ηc��y0eY{�L�%t�!�J`K]o2��g1���֯w=Qp$n��ŧ2�cw��I,
�����5p�g����"���:̹i��=}��(ֻ�7���9lE����H�I#�I$MӀLW���E.������������Vv�-�2��,M�Ƞ��J���T���:@�

�((/-���ETgn&%E���UT9J��R�F*
<h���k+�EEY�d�Ӷb�,X��X��VJ񪓌(���SX[j���mC5I���b(�P�yh�Xă��[H����1E��W3��x�Cf�U�V#hQ"""��&��_}��f�vyۻ 
�Br��p��szTٙ�.!��>�����W��WN�g�wW����$D�w��$=�d`���?����u�����n�P�b~L� Pa��F�y�d!��w�0�V}���5qx/��.��������`�j)3d����<��e��<T@��a{��){�w�=ק>�����yI���3�<d��Ӊ �G(���3]Xi �|ʞ�^�aa�
����%H/hS�ް�_}�����)�E��T���0ڡY�%H)3������:aR��Շ�1���i ��7՚H(�P�J�S�^W�y���y�4�}�+T�V�Ry���X�,���B����H)�vO�H
,�%d��'>���%G�y�<�^k���~��L*AtÈbA@Qa�
��T������Xt¦��c���*��&�AH\�Aꐬ�4��R
M�[��{9�}�9��0;j��Ă��_ �<��m���bNT���*�AC�� ��Kl��t�j�$�֐PS/~�s��k�w� ��l*q��)�0�l�aH/��E ���1��T��!Xv�T��Rm
����+��:����T��v�`�z�7(����#:#.�\RE��9�|;w�z��1�	~W�)�5�� �̹G�������J۷-)�o]�{y�������O��8�I�	��Ȫ(m%He�~2^��0�
°�)��b��R�H=R�O���}����}��S�Ĩ�@Q}2��N2��J�m�f��a�
���>B��Qa�
��_Xi �a�3�(��6\������=���4����bA@�s)�B���j�YY+mI�TR>��R_Y=M0��C�� ��+�|�w���sސ�%H)��՝2cXT���T����aP*Afjɉ���z����l��$��LE �����*N����]oߵ�w�B��Y�
A}��PP��La�
ɨʐrÌ1�L*AM�LH,0��E����1 ��Os�!Xm�e�;���^&���{&���!PT�i���]NX�B���>M$�Z
�PR'l� �CybŇL+'̩=B�<�>�]���}�^�|�0���`H,5���a�o��A|`]}�1E�;dĂ��<�A���i��y���Xj�AI�g�:3���_k>�g�~H,�~�z��ά18n���I�
,�9f!�J�ݤ����t���1 �uh�� �HT���y�r���Z��{�a\`T��ĭd��û<eCE�}�+�o04�X�'�T�a�
ï�1 ����՛a�
��zo�s�u�v$����C�*AH,������WZ�=� ��TU'�T��}� <��>M�:IP>J�����O�~>ߝ1�^��K���!�n_c�R�us?8��e~�{]/߼�>�$ɋhػԔ��4������T���ﾯ�=ߛ�=�LH,���H)�~{a�,:aXi�I� �0�2�@���^�V�k!�����bAH.���4�Y�w�wo�y�}wגk���M!�4��;jA`q���1 ��\H,����x�þ�pt�R
����*���� �g̙g;ߟ}�y�y
�;I�v�>I;@��$�'��$1��������j�����]o��x{<I�!m ��
��@ă�_ra�
��i�z��sbIY�dR<g��
Ì���C�H.���}�^��^{߄�A`xԃՁی+;LH)P*�P�%H,�嘐R��V,;aS[�bO�4}a����QOP*A��E�k�}��stP+<��_XiH)��:�9�A��I���I� �3�
ANY=t�P��2�=La��޻믵�>�~N�
C�fT��["��+T��2c�T��`T����
��R
x��;�+a^���4�Pמ{�￹�7�}s�x����eH,�OO.��*a�>T4�Xk�I� �0ٔ��r�M��0�5l;IP*T���W���5�~��>��o�$}�2M}HVv}CI큮�$�}`bAC�8�rɾ���ccR
iR
Aa�(�#9�����7��߿o���JŇ�>�R
NЬ���5�CI�@��1 �E����A|M�d�AI�P��`xԇv�r�1��u�<'��/����Y/�%'U�d��k�N�?5Ewh����ks+]z�}�l�1h���#e�!��Y�>7�}n�:|ֹ޻����\��Bk3^��H,�"��癐8Ԃ��n��c�2�P4�ĕM�ACԕ�udăݞ�}��0����Rͻ�<�:�_s��N�M�T=T�� ^R�Ht�X �7@��J�%H,���H<�7��j�H)��bO��>eE ��}~��]y�7�{��AH9�Cl4�l+<�Ɉz��6��bAH.�d�Ryx�I�&�(bA@]Z���<�|� ���f��7���o�,6Γ>7f$�̠(��Շ��Aa�咱a� ��
�0*�8�
� T���z���;aR����}/;��o�H({�E�Y5�1!հ4�R��}���!�Y8���� ��c��ĂÙa�|��'y缺Ϸ�>�^ �ĕ��,ߖM0�I�*A`u��
)�~`T���H�HV�g�i��R
A}d���*Aa�������{ߚ�:��i ���1�j�H{���!Y��E ��]d4�P4{LՇ�1�l+����+5��P�t�$�Y�%}��\����;aĆ� �OZ��R[�H=Sz�i�L�1�0�z� (�=�OYR8nɞY+�5CI'��}y�:]��;�~$�M�T=IRtP+XV�����/�
����MٝR��=�R
s�sA�}�=��?��~����ҧ�Y�|ko��>Z�����rbZK�΂���	�-���W���Z�����Vou�1f��#�3�e��.xT]�6�d���T���'y��|��nü߿�hXu��h:d"b~WƳ��o}���� .Aڳ�L�,y x�v�+嫗�$�u�#����!հΟ�/Hh�M�7��;�K���,�a�j��%�|.ݷ@��=���.�[[G�U_��_�D��\m!�[����t���d�ݯ� <:�ҵ2,�l!�NSt{��_>�w���;$���j���<h�#HtM>���^{����ˊ�g?gs]�,�C�?=�Z(jn_Viع���!_]�*��~�CǍ�
wuզb�����|0�m�6B���#"|����[��q���6a[x}�.��Jl�v���-J�+pP�uI����̓�>{Ktq�o��A��kQ�c���~�����]��q���HY�28�Ô+�����29/ȿ#�'��F��?���Ӈ��r�i}�T��>�_��g|G�6E{Ϲq� �O��bfט鳺�=�dv�>����#�1���q�o�/��麶����y be��?�1��9Y��?/�4C�){�Y��]�i��<p���ǈ��~a
\���"���4�~䁈iw:�5|������b�݂��t �Gb�)�#�Hg��n�=@x�t�{.�����+?VDx�I��g.�=U2�a�;z��<e(X��H�0�0�g�A�TMkw<uL�+7.��[�I�̑�9�A���n�a����SwO�]J"���y2����@�e��>7���������כ�侣��8�c������1=_C�Y~���o�8��\���K�]t6�u�t]^4���{X���|����(x����U]/oC�gvV�z��4G��(�E�aZ������)�ue&g���w��7�l�7��/�tF�-�܀~Xo3U�����s�b���^�������ƾ^�x
ʪ�Z9�aVG����8����!����RY��{�!�y!GP����]!E����^ZB��aN�����A�����<D�0�����'�jd�m!dGm1iT9H;��O�ֽ3$m�Y��ok�����v{x(_��j�?���|�ǰ�eˆ�m�y�;��Ⱦ�r�ⶸ�0r�m�i�{��_}��A�<�������.��t8�6��O
5����R��C�h��0�i`�g��uЌ�t���dQ��+/�?��a;{�����Z��2����Dt_Y���ƭ�ce��8�XB��7�;�;�����}���Y%9C�����<l��p��q��"���W�D3��=�d�x�������eO/
}��k�W������<@x�/��e/���x�!^���Ƀ�g/!�c��ŤQh�h/E�����GRF�Eg�+�Zk�-adKL]�Y9�畲U{��> ���nt�)�x������DqX��l�8�7��ovܿ0dt�m�kA	ޘ���]]ɭ·0T��h�ԺP�)��T�͸���V��L
���֓뗜���Mw�o�=OS9z;x˺v��{?�/��oU_��:��0���	 ����"-��ǈ���R���7��ր��`#ZE���,������U�i�o^�p���������~�Vx�{�������t���Vz)����?J�4������]W*u���ز�F8�ȉӜ����t�,Lr�����	2+�Q�����4b&��>���W��ٿC�⏋b�h���gr��j�v��(�6�y�Rfr�d&����~$��3����eK쳀��� ����2.���ӑ�)�tX^��s*8$���	�V�ބ��Zs,�\g����|��H$3I�p4�5f��n>X�H�$v����y{��M���~�߇�� \�8�w��WOܻz��bO�����;L�GΏ=׻�|}��܌q����5ab��~c�Ֆ�0�������U�A����5��"������e[�R�m	��̊���x��{v�0�����-�`�A??��
��!�bK`����O���3�*�CW�=<|w^}y/�V%d��Ŷ}~�/�P#N4	�l���k�{��]���ޕ;�`�Qj6E{�r�HE��D��k��ovP� �+;)��f��O���}"8��4~�^�C�Ve���?B�ӕ��Xc��Kja�uӼ��ꝾuO3�}ruF�>>&���{��q��_��v�L�������T�Bx�p�R`�:�AU��ˮ�1`��g�sU�D�Dc�5k[�6yH�V_pWzp�E��ۭ�\ȢQ8
:���Q9xv��Q�[�Ո���&������n *}ݏ��縢�@��u;��d�iM�FP	;zjq߹�l�Gu�.��\�Q�W2�Èd����`���k>x�Kmm���0[,�wo)��_,�r�[��.܆w���v��v�"��F�iW\xNUZ����ϸ��q�D��sr�G68���-.�S5f<0[\r���2͌:��n�.Vs�q"�Ԯ�/p��r���e��v�����o6@oWE������V�n�Kj�ƪ}����C�'��j��L��~xv���/�?�.��#j��b7��${���16�/i�kWu¶����U\�߃G�����wj��b��Rq੪ ǊQ8D�������'g��uO/��L�Z� s[3	�w�+��rF3�u��}�tQ��\��`��b�3���дU��I����8g�ۏ�m�Q\��XFIG+�|#U�I٥ӳ�����l�+VfF�$�r �"/z��7�-.n�/]$("x,��{+����ra!�v���@�<�>�+�������{�j�-�3݈��{�f�6��	˦�LJ�7���T���{+s^�{�z�TUmWK#ݽA�+6�S4,u&�[3��s�qfA����rA%\�Ӿ&N���[�;w�Uj�/!H�I#�I"��K�.ιu�w���||>���(�����#�N�v�+��,����Օ(:J,A2�"�E4�Ci��QE"��St�8��f�QQ��T��*(�jʦ2��F"ɍa�QQwlQ5K`��Y��(�؊j�[h���*"��pZ՜��c"� �ݳr��P�P�&��u�*���fR�+��O)M�r��\�Q�ZÚ�6��[]sj���Z�U�T�V'4�n׎�y�B������^k��c� m���V�@����}�	��q���|b���D�����}��'<=��הD�Q��)*/������?r�z_f���@VF�r����I�7p����^��z���..(pA�?1��ƠvE�!+ή����ύ\�������� �(��V~C�e�s�ώ��\�E�Ԧ4�_v!=�H9�:ޫS}�{y�g��긄��,���_p�*5��v����:*4l�h���ő�L>^?8�Ů��o����b��0�ZFG�-��Ư�E�g��/Su�ޫ����R�;��ΐ,��x�J��]�$���+���P�V�xQ��jj�_V/��o�y
�f�7C9�&b�x�C�h�:�^����-8�,�w������ކ�Ռ�Ksy˭.nCl��X%��W�U}���g�x�2�����i�/�OA�C�B,�1�������8��l��3�/�!D����]������ Ahz����/��"F�zK��e]_s����y<�����]���k1���t�^^޾���+�����q��<!�Ť5m�
f<�UQG�j��y���� ]��}ok%wy��l<����|�]���c5������ނ^n��a�a�O���z�l��1������m+��9\�/��/���!�B��!�dgw/sC_*>�o���#�"Μ�Hg�${�MCO�n�O�Z����]�&k�[}&K����7۸��Vk���v�ۇS�}uGe"xd"ȴD˩�<������]�|>� 2N��e}�}6~�p���e���G�~��י(bGZ�!�@A|�"R@T����[��ǹ��<���"�����Z��KQ�����[��#�!GH����"�O�Y�.3��7/��2بF?y���ag��}Y�~��_E�Or���Ӈ� �ǈ��(�~_@��Q~��Z�TE5�C ����DY�⒇��Dq�{����p�8����t��?dVx�y<C]R�����q�zxn���~aކ�8'��S�ez�W�+x6,��q�ȉ��Q|�� �:[���h��&��4��
t�n��nz˷:�ߖd!{���L��VQSj<��:J���0���w�2)y�]���͇�����>��{+}�T���4G��!����ӗƈ��H�rw������oş��|F�A~������,��	��@G�P�ϥ�^��g�壕x���;�zu}�ۛ��uո���>���eD�p�/��물�Wǀ��������^~�xwʄ���l��	A�e��0Z�j�}7�J�����L�����F��?-B���([R�X�9q��׽^�t��4|��#�ZVO��j�vo�繎c����*���,_��f�?G5a����u߳����jl���q�M/W���{�]r���yj4�]d,�����"tN��F�T�|WGf�\�T�h)wYM\�u��t�/e�S`���]�����|>rHJϥ��V?]o����N�]K�7_��m])4�U]��T��~G;���x�^\Y��5�x�=���q�ؼZ@�w�N_i�� �u|��}]~����(��L+Z~7-]^e+�����}^(Dk�=�V���HB(��4|~����M�y~���^yu��g�<^��}	"�Zm&s���̓���Ͻ�h�(|<���?���$�}^��NI�~4k� �4�P�oA@��YI��o�x���$�ރe��̠����
+Cn^u��7�> *"-�Q<��Ƣ��_X�)m^Uc)��k/I
�a�MU^i	��WZ��q�T��T;��$2ar�[��v|�z��j�-v̎pQ�X�?U}U����~2�L���W��Õgo΄��M5�����wSo԰�A�,��+���0�CP��Tr�s|7�M��}{_N��1di��k�Di�s�eh�ͭ�+��x�O���~B˥��0��Y��+^~[]ߕ}ܴ���OH��98疞��5���3uC0�VA"������1HQ]�Kw�~���>�B�3����a$YH&{9�{~��辢,�:x�&�_m1iU�E�sr_^U��a�mg������Du�"��7u�+Q�����|����4���`�B�����������SR/n�gYyL�B�fr���s�7y-�[���w���!��Yu���1
���sM�Ij�i�1eI�n){a%���������/#��)/�RW���h�<F氭n�烜�Ow|���g�]/���������i���W��2�n���TB+W����X{Pqx�#Ůc�K�Gy��B�8}�#��Ai�D�t�Hw������Z�ow���ܾ�-�Ӝ5�H/�Y��}wso@�xĳ>s*��Eb�v /�äB(��e��,�"�x$(=zD�4�8"�Ȳ�Y�1k�R{�*{|�k���8֡�N�`���>#����zz�vW���b�H���v�兞;`��'�Oe����#G�e�	 ��-+䈰���RU���� ۛ�30�jCPygs�r2��Ul	�i�bt������w�P0b������r�n�s�蒱r?����y3a����|'밯�	)�G�ZE��?x�	�N��^����K�S��ޞ*��===���w��^��3����j�j��M����7J�X"Ϸ�7���\��<G�;WM�,�Ta�㔉�~B��ث������?!K�%�gO�<|a*�b�糲2y�p��YV}A����䰿!��Ci��7W}�0���8j�L�_#���6`��3䆉�䯲��uaU�g�V��!-<L�  ~�S�~��g���,f���^/ʎrܾ�ǈ�*��O\/��v\���I}��x���o��f��h��%R��3�.���.5
��vi������H��zn&��1�,�{\�qp�	;��1DlG|ytt���2��7L��~ ��:��C�����U��CL?/�P��,�`Q��h-<M�j�_��+����5~��_?w��r��ml<���������{w:�ּ��nծ��ʹ��m.���q!�g�5�F�hh/�^!v߮�ޛ��_-C�d�#TCCK�+��/�P���^�L���uT�� ���/�S��4;�ˏ�Ѵu�L��"P<E���D�qM�'!@�#NW;;ۖ�*[Yw���=�+��<~���!����λ���}����#�E���Ϫ�\����YKL��g�>M��b��@��}�ʽ�~��v|i��+(�&�B!�\+�K��W�Hz�m��u���En�:�d=|������[�U^�����#/X<7�J�W0����Ƈ|�s��Ō���=�Օ^��W�^��2����L��7����{���T�%����Ʊd�ejpg�vS�&��jK'r��E������r	+��צ�D�y�r���ո�׸e򩼲��M�|�x�J*w��n��o.\��=G�ww����;������N阙7Z�>�^QtԎ��y�GN��̿)5��p�>�^� #rAsx��4b��A�-ٲ��m`e��oQo6��:�E�797e�ӽ[yL�J5#����|����y������0��nK�G~�C]f���Wd	Pq�,�Q��sq�wg��I	�Ӽ����f8҈wǇd{OX]����=�ֶ8�u���eW(��Hc�����5����X͖��7��hɢ.�����8�I>��E� �Y]����
B�U�a�ǆ��:�	Ȅ̩�j�*�qɾ�B�^��F�ojA���~�*و�v
����-k��ˤ�7�����W<5�ڹ���'d��{ ��ʹpLѝ��
�\s��q�#��Ny3z!}NJ��p�������Θ�M
�h"�ޮ5[Vb<&^>�{���6����˛sh�u����L�:��9k9�u�I��R#ݻyG���ڀ�Kgv�w}Ԓ���l,7�Vl�aܳnú����Ӟu����v�::Yz�<!oo�4�Ou�q�m�t�۹�������1�:��u�7�"�-��)��
������F,��5�{�2*.��g��8Df�۫���8B�2�V���!>��n�T,Vo�n<�Oik�9���7EH�!�$�+�(��Im���m����:�(�M���^�� ���h��k�JD�Y�����,�̡�%Z�ڝ��RI�:&�.w[T�`}&�I)d..0��)|,�7V�q-��U�L��I�I$nI$�'�RMF����UW�x{���(��4�)��1�F�V]}c��dX�a��ƪ�I[�J����X����R��ޱ�x�#Z�X���)r���-*�m8浈����bꁤ�R��V�Q%ˈ�hX�x�$*[��elK�ӄq��X��r�qt�bU6�U�U�V+�M&�aR�����7V�(Qc&f9әyM--�k��pj8sV�8Q�KmŷiQ�+q�)V�h�fd�\]9�q¬mզ6�X�eB��˙���)�m���-榄�B�ڂ�1�hԭ�֪)�p���h�S0�5((b�ˬ���_�/�{�2x�L�Ur��j��k��;y�p��[%Ă�W��_U}^����W��i�4@٥���N5�V����r:g�l_��@jn������<�z����;��8�pgw���Z1��lK�g��Vq�SO#C�}�k���W��{�َ�vvjS&9+G<;�IT�#)*�y�y5���)��cTq����+��ӶN+�|���;�h�V��giq�D��;�:Z���w�{��n8ɻ�]m��4ˈ��v'�{_h~��1��u�<�@�Ѕ:�J���EY9X����gK�&�������t˸#��q���̊AL�:���Տi'���x�I��#b�i���B�_���v���Mxo&���!�\:0��P�ovs�Y3hN��u"+ҢXkС��n�ISMv��5�j�~V�|��f��S��l#�$������cN�T"�i�5]1�_,X�����Q�~�]�fUȆ�S/�K�w3I��EM2��Ӂ��kC�U����`���ǿoVۿ^\6���i�e�;��p�w�ʳs3b��)�����MU�Zw��g�38�e_��q�#�W`˵g��w]�TWo��)��O�2㛑��ڤ���W����4��zW��C	��}���fý�Q��R;���B��-�'x֠�d����G�$3݃�-�"�]0`�w1
���u��$U��Q��j�47��ev�0�$���,��қjf����ם%�MC�r͘�����IZO�]S�p{S����G�{^Tĸ`��_����SӬϠ��k�΃X�D��|��z��ǍA��MA-�O�cmL�{���K�1���A��u��^��
��Ǉ�~�R��6X��*�4%K�I�N��´��yb�U�U<�JD�V��k;H�*���m��f� �WS�!������~�����g�/�?p��ZFĻ��L�>�=$�/����aWM*�Tx����!�x}^�����\��(���xuϠ�&1��f�����VE�<�Ռ*n�͢&��E�fb?[�2]�@r�ʼ��gZ��(D�^����.�*P�\��c���٣���x}�IF�#�r�9��[��o�ua�h�Bx�븮�ej;�˖x���l��"�e�#�ײ]��%���{*�y'��-p�p��f�s�������J�9I^ �l%�Oݓ~3/G��vi.����i}�&m�uvI��ga-�l��UC�<��_���>����"/>�Z��_
�'wz~�+�'����j���7�Im=���&b��9������4~*
5}<�5َ��+sP��l�R��T!m�E����=7�ڂ�g&55����]Ԗ�9d4܂"}���վ��ϗ<���#y=�ߘ����["�������ծ,�Ƚ"���2���O.����U�6�l����͌��w�����3'�Um�Z��nc���$���ׅv�`�Q���xW]��0b�<�U��Ū��$�����g�$��D�H��f����%̕j�a����{�������zN{V�nl1hu�5�_�A�Iw��a����|���k��ʸ��ңΉ��5e���e��r��Lq��"�^��9��gc+�����̛'��B��=�M-��ו;b� ��5��Eb���\60瓮���ړ$�:����-����oW���2�Y�G�P��-���wL�pes���@FI':�P����>��t�'*
����I��yм�|,�y�z��>�y��j%
����ѡ]:['8\�/�e���u}ݬWov�v��)b3�hn:7����L�I,���O������~v][w��h����g��"�q��G)�u�5����{��g��@���n�yp��s�<'BI�2o,t�+�.��͙m�+�2#���j��ܝb4=���Ue�q�ru �a�A*��F�ҫ>����1F�A�u�����T���GF�
�s��9:�Uƶ��׸e��nm�uh��ol=�tg����ٮ̏ɱ�o�X �����a.��F����d0�]p<�ךEhUh�XGl��?�Z�k����y��-̔�(���՚��|b�<��Ύ�w����Dڎ��,�'����x���bЮ_�?���Z��와¸xXL��י_2S��͝f���U|mܺ�;m�9,?m��4ݱf�`<����B���X�;��o}�>���Da�;M�<��x��ug��Ď�*��3:�vA� S��+��}S�d(6��϶AoĹ�(1�`�ȹn�la�Y���}W��+��DM+�QF��"��9����K��	��-�2v;J�jU|W[�<Tt���3�ՙZVyyY�1���6^��>Z_�o��d�CD�3!��O5}��[|%��gW��� ��=�? ���Cv#A��fw���}���<+F�s�^�����3-�8:���O ��u�(j�\�p�称��:yt��F�>	�������B�-Y�)�E����c2�;��+������q۟�Eo�7b��|�Q��f��V�L�v���5��Efe_���K"{�Y��=���:�7�#1iC#/	����H"9�Rﲣ��.<BMM���w�(�X*��gE��$�܎�˚�-}���{g��CWwYسuÔ`�QXr>'��ջs�^����+?0�F������{�6.���۲�t�}{R,P��t3��q��Su�M��y�Mf�����gе�U���uCG����ɾW!�\���x��Ub^FU�}U�,t��{���S9&u��xqzr�>U��h`����2l�;��u�#&	����Y�l�><�-@W=���B��D���UZ��e�Gjb�����f�E���������\W�BG�=�ey[+��}c��;�QEL!��n�34e����Դ�ͪ[�U�;Hut�Y�����Js�R�?�yy��t�k��)�ޮ:u)f��,��n��/&l��$�MÍ����et�3��0�5gj���ӑ�A�jD����x2�:�Bd
���"���0��T��}��Qol��4��JPAǍ���F����Π�p�8�j�j�ib��dfPv��j�E�Y���,�6�g9^�!�	��	���ui�c���xP�E&p]�77n.�*��L��!^��+j���,
�ˉ͍�@�:�s�vp�;"@�
"cݚU�&X��J��FE�NbvuWk5Z.2��K[v�Ns��	U�s.��T"fA�s7���}/�36Q�X�Y�8��*�*L��LOL�iE�d��=���{�'w{v�Z�N�r���4ea�����A�8�]��A��V|K�̦k�N���'�[f����S]������źk�k��4,��	���'R8s�m`�Y|�X��(���@�h��MZ� D�Q�i�A�P�N��lPD���G�.� ���,5.j&^f���H��o.�lV�R(�<��f�M�/��5r�NRs+/�p쥨�T<u�(e6�팤iW}���.b�wZ`�L�!;vj��Y�+3,����5wJuM�6^��S{B�B:���a��9:�y��ɺ�.[=�5V�8�{�9����.KT��5t��[�{���y	�)$�HܒIR�ǒ����c�};ߙIJ�A�����UĢ_s���4y�j��eQ�leE�Y���4kK��\�na�1�PDS-U�9��y�1�[TձQ8��R��m-���eEYƮ��*m�Վ���WT�op�n�̚Pˣ+Yn9r��k�Z驜L2�H���ۋ��Q�k���Khc���e�.72�c��)�Sb���]-���QX�e�J
L��#ne�ڢ(�iV&%����(q�4U9��1�Ee-j*��E�QX+G������a;�u��x����S�]6�s7�*���UP�H�x��w�z�Χ�y�ȡ�M"��w'�Y�5�R��x�[�G&|=iѮT;b��J�1Y��iokm�u��v�gjn�Hu���ɋ�Z�Sw'/o�9��C��Z�Ɔ[Jk�<VOYGb�B�+�_��D{��=3V���<�;�ޡ����uk�ZT����&!U���&ŏ2�]w-<�$���v}�.s�%�f�X�#�M-R�7��گ-�A]Q�iVu�Քā��C��%���`�A��(gs~��s�-���N��-�\n=�[V����������}r�?�˵�J����ՃH����ť}���M�fκ���UZj�eu��0�W�WI��G��'�^�Y�]J�������3OI�|���6W���p�o�W7��XJ^��;UM�]�7��߫\��I�
��M�r������D�\Ϋe�Okh1�U{]�F������OQ�W'=��L�~�WJ�lt�k��|=������{x����Y��B�?:QQ̉�4e���o�F�{�
����\5ݽۡ#��A��Ͷo���.�2��Od5�k��RF�v���ζ�M�琺e���J����-���s{���+D���`�	��0����7(��U��}o�ǱA�[ds�u�ZJ�r/�g�5E��"a^��)-E�Y=&���Dyc'�XZEA<�~�K��Oe���λhk��Jؔ(�ۙf�#��2�{���&�Wym2�}ɝ�0R�&ߚq=e%f��U5�OJg��[�ͨ5���*�=��.榝m�)�]���3�;��{��Mg��D�����g��E��~����ػv	tʖ�*�b��P�I����5̌�~�ގW��cҖr��|nV����-��&�
3`q+��|L����?��'��1g�}qy_��[�Glz+�V���T��=�o:᳅���c�<��p�sE���<�͗AO�Œc4��"�w%{��=k���+��a�G~a�.��<�T.̸]�#ި非���e�s��;� ѽ�z�J�;�����%�ް��5��Ӕ��w��)�s�W�j���G�]V:��v�?k��J|��y7X�0�\iU��G��`�{ӳ���D���'���a�9g�t7
�\l�j�C.]�u.����yڃ���3�Vb��
?���S��^[�:��CqS�p��i��k��%z�$mbr�d�^�@֭�L��0o�2y��Q՛2��ꠀK.��F�w�:J�����k.��,AG$oq�4�j{P�C�m��Wc<�U~���g�f�}�0
�l�(��A��=^�a;�KwKM.΍�*�|K���r�k�����t�B�ؽ;�j
^�@�xJ���6�4��A�fI�^�c�mέ^�)Q���yi;��PԼˋ�ּ=C���R�nu���!��J�Ԅ�ۮ�M][A�V)��#Yd�1o����{�[d��73�����7�<�#{�K=x�H1���ڋp��:
C��z�*���[�Q�U�Z�����:�h{��ܦ�鋉� ����B(���9��wdj�)ί��E���f�{�=WX&�AN�f����j�"io/I �+i�]��]���=��	~nN��N�ǭ���S:��3�ߞIj�+�J��J23��)��gv͒�<��)�О�Jd�H�w�]cMb2�JS�[!3-z�q˛�\~l٥����eި�6��Y����n�ZE�ٽ\�v���q��\�E���u�3�_���7�7s����v(���V<i_j����ئ�!��x"[uٜ�R��nþ+��O[؅gp���չ��_�K���z�ʹ���B�Vy!���X�֍`������v;6$q�+Ҍ��o]�z3�FR�t�޿-�Gxz�-STfQI�^{:Fyz��Z�k{��W��'
��w�y���7JX���ض>����G�ك��8՚\3������T��K|a�;��{�¼.c�\�`w����l�;��f+��9b���Z'\�­
�vJ�/v���K���	َR���?�>k
Ӈ�ٔZ���>Ê�L��	�)����sn��\*l>�):h��L7�����}FM3�-V���J\?Ĳ��ph�����y)�sK>��F(yO� zW�H��2�Oz�͇��h��{�x��%s��͜�2̊��4B�끮�8�'�?]��x޽��"M���4���|��`�Co'����T;5B�jt#�5�Y0���upŞ����
x)�L%}~��-�M%z��̽�4�V�zr R�5w�;XgU>�~"@�i]بl�y����e�ݭ3�v��{�!�O���>�k�L�`���0�W��~Z�L��1��)��:�~�>5Z!Ӵ�;���fm8�̙ɴ+n.cV0���|L�^q>~�s��@�n#�K�`HgO f5� �=�:u��������^{I�gCw���u��}�D�'=o�����R��v_�5tE5n��N�p�Wwƥlk{(��#^geGr���g ���)NO����dhp>��Nlݳ^��E�Ʊ+���P}�=Y� �=���ov�uGZ��Gpq=��R�O�`�K�����۝ĥ�Fv�3 wx/�{���8"��Y`��ꪮ�A��C�Z7`���8�~��n��#���N���㊂��T��9�$ˮX�(��;�����V�m���k&��֛�4�'B�.ƾ��I�Ğ�:��K�m������0�&N��6^7=�S��e�HT8�Z�K���l��a��'H����f;9;��)��Z�&B*��y�U+gejֻ��(��c�^�٤^��	���n�Zy"�SVҰ��m<��[�_���i��6��c�&�������Fu��Vg,��7�5��+S�$�X�E�ܕ�����P�X;D��)k��q���MUW]G]ڷ�Z�5��=�6�fӬ&���.v��[�I5�7gjB8��[7eJWX����.@����v����YwDȑ���,�����ݢзtp�hRCOST�U۝ǐ�B�'{gm����t�)��S��k]"]�h��Y����˸�8��X5�:�{�op�)$�k�>�ڏ�Y�U��8K��q�ٲ��=n���K]�t�h��ƞ;������e�֬e��r�B�*�Z�k�G
�D4���w-���:����B�
�}ip̗خ�!\Y*b�Db�N�roR����=(S��:��ti�u�����R
u0`O��N�]�+u�Gj��,VJ��z_-he]����j�,��-Y}��@⬐2��e2]��b�$U��)�����vS�Y�J�2yٍ]�%�����(�`��2�<�<�5-��:�m���D�,c��B���9|��Fj]���aN�`'{����D�ܼ�l|.�;�D����7䳯oWr�ĕ(�|#�����K�Xib�)e���cN.�\�3]�]ǲ�e$�0��ӧ���p`��;-S�7�ʒ� �݂MPA�͒�n�(^�5J΂�:p��I̆BB�J׹/�ݔԴ���r��j�����$�G$�H�r���4C�&p��ʵԑ�����Z´�-Ly��C�+�A��L��+Z�E��TMQ����TUպEQE�8�D9��\k���1��p���Ҧ%D���UU�q*�Yk�cP�V�QUB�J��&D�\�m�q�
���&!Y1&��i���TƢS0R��ˍ��B��p�<�ӡƱ�**��UbѣmDb)V[E�*�*"�q�cS��#�J1j-fҫ2��
���D��hQ�*i��b[h��Ң�Q"�-�D��^���j��bUe��Bc�ق�}g4���g�u�����x.����Z)tc�ި�՟��3�nDQ���6x�d"B�:�f�e!�5��{f
ǐ�(��/�˪���z�&L+ �(+�R߱Փyn���C��9�)�̝��+�x��n�a��`0������<43���p�����CȮ��wJ�-�~9�[օgW�nUx�Y��)����yN�8��ǝ��3d�'��1��T0F�t7��2f�"}+7��g�zH�A��
v;�ġ��-#V������0�hQL�nYD��Y-@i���K7��$��;whRA��
Þ�@2Ki��{Ņ��Z?��c�|�����p�^<�Y�6ȿ�-7�6
�Q�~삱�Vǧo{�r�N�*�9kj7b���P��訞��Rcz��qY���4v����O��g�z�U���:���2�meN�ۃg�큅^U9�OJvz���#��{;���r��f�h��j�v�8�^��$�8Z�~����o��Y�W��-�{}�L���)Q�]���T�0[V�k7�

º����C�1j��HX��+��*zf�v���ø���� ��"�Hz��	��sl��̡]r��w#�9�-�a��W���|���e?�o��xY�Qn������Ցs1�A�A�0��_=v)��#�])wWC�zN����Z@�Xp����2�:��`�Ԩs�K����I����>&��5��j�U^n��r������Җ[*��D�N�A��[e����'X6�*j�����T!�*X��zF��n�=��qzr,4�sQ����<���-���*����"�M���Ƴϩt�f��~/�xUlu,�*�QZP�����1JSY�+�v�,�m�]�m̮仞]�Xh������jV茹hZu��2(�f���a��J������p>�V�͓�J��hj芳��y���&*S�7�rW����7Ҫz�^��z�̗��/���j�n�wUޣ���Y7�jE�q�K��^�~����2����\lK�Zz�:n��>�N��S��V�v�N{�=^��:~^�nP�Q�ޝ�j�Mˤ;WOA]6���p+������:�MމSXY�A#�~�^�rWr^���/$����Vb�D�z�1��mq>X�4f�~���{~���AML�����-��gv̓���v�qf����&*W;���mg"�|]�nVA�b��`�}o�S���N���,㛆8��M�*p}Ӈ�&nh�����Sv�J����/f졤dY��q�H�g3��k٬c�Y��e��	�0GY�6	��ni5�"��}�9'3TS(�{Mm.����|D�X�ܲRt�K����K�����f��q:\]�lR�Ҽ�N�p�����|����B���g�W�U�#}���ϑ�zH~wR�Z��>��w~�Ay|%XW��]3���J��{!�LC�XӼÇ�;��d�՗:I��YmƵ�7Wt�˓i��aYH�}������Άo�|k􎺸��؝���F�P��g��+�?�U�J���*���%0���������ۄt����[�]�)Y����ߛ��0�zE7Ot�'׻�@���N>!n����GÁ�m�I��}J��oG�Ô�<Jo�b���p*��K�8sU���Mf�I� ��7�,4�Q�^��^w��q�۹٬Vs���em��=��3S��}ff��M�N��:w�a�ޙ|��Ƚ&p��Iov��H��/?z�%j�M{1"lu<�P�ȳU j���kV��H�#^�+�	���X��3�5����9��^{A����S3j��6��>��;��2e�{m(sK>��^_�ދ*]3�L�3�����\7�
Fty.��l<���_�n�Zv.&�)֬�8�2*a��v0��5���l2^�UP#�נ��x��l*J�=�}d1��m:�.^���s&�{e�#d�z�W��j��!\��bd@z�'e��>I[��Θ��f��&e^wPZ�V)��Nŵ
�țS�kЖ�>n��#���{k���e�Ik:(�^�O�x�'��Y7�0���~���>��َ�	�b7��d�C���ʽp;VJ��S6�.��;�߲T�mIj���JG],�
�wB�����A���2��߇Ş��S'����W`���o2xx"��Y���X�G�z!9"=�F�Zy����7�9��X��С��FV��{h$�]C��E����Ub��8:\��¶l�6�Bi?4�:�6�^[O��Ʋ�3�۶�_����[�{3�V+�1���t�Xqj�z�Jl=f�;�w�Iۥ��y"��[����T�W�/�T��ծ���'�]J���֧[^���(�Κ�E�B��^��*+/ �qs�j�g	���ap�u�2�-�+�ʽ����U�9&�B��N�T�\��O{}M�~���6?wo��'G���DG��)뾥�ڶ�A9�̒�4����^TI9��݂Җ����;0bn�����SY��<*�J�'=�z:��M�o��Iĳ8�ȕ��<['�2��ѕE���Ҿڌ�Vfc�ڏ����0ݛ��dV��I���V����O�驛�{���Hd����y>��9cS;x�QD�4�y��q���69��(R>`�Ժ�J��^�К���[8��Ug��>�+�ɿ��K�O�'`�|��%w����<�߭p�1Vc�.�G}�Q5�m(�N���o����VA{�;�r��381�m"^�<��a�j�W�F3|��m?N���k��:#Ն۬��3��b���e9wkqu!yޣ�y�ò���91��34-NƜ~+u-�6Ͻ�+r�s��%<_@诡������}��`�F���]�����fC�egR�.��v����A�l�D��ۮ������M��Z+)�zf�oB�]��$v��&z.f�9����M����zƝxE��+I�A¯u���-���;�/Y�to<9Rҫ����w�^���.��JǇ����piR��b�]ʛ�&x��-Ѥ��w(���n(
�:�-�zyCt����f��f��P	W��7&Y����"���Y�y��'j��֮����$G^��%���M��/y���/�U{��[2�aWx7�֚�Gs�N��;D/��*�~�����u��� (=�]���v u$qB�f��92���ǅ��gH+R�NR�<�u+U�N�|pbt��M+�W�Vu�U+�x��Q�ځ��q��hb�����29F��uWn���<X�F�pL˽3�#M��p�w��)�h��M��H%�y����c�'ui(��)���f�y��V����r�R���օDg���q�ē0�����=���,�%�xw4wۈ����g<�;B��"L��k�ɾ�����F6�(lQ�1��H0^�f\��Uŝ�]��&�A.�|�M�u��Z0"u�ys�U�c�[®L�;��=�e�+�n����AVh�r���o=o9e8e��}�q��u�A�������������3����'��h�SMC��_�OyS�a�$rI$��$�"�.�e����D��m�������O4��P�UkF�Qb�J�X�(*�-��j)R[`T�ZVТ��st֬�E�Ջvc�(*Q��T���)U�r1Q�Ң:�,PR�%�iPb���Yq� .5b"T�-��T�t̖"�J��e��iZ2H�Ͳ\%�)uJ�*�+�U�T�j"��ƴ��V�KbЭ�]�t�ɷ�h�h(��IR���)]���"D����Z˼I�}�����{f).-#�|�Cqu踓���e���U��xy>��F�����ƭ�[�Qub>(Ψ����!���7�a�u��c�] �u˹٨W�]�6z���@~A�7iWx��4J8��&�T�d�L�*q'����7*��pվ���\^=�"�R�)��}_j�n�R�Ǩ^gG�?��CS����1��޵{����^,K<ϡ�{��u�N��wuaD�S���f[[=�#�>�@@y�#�����;=���ބa߱S֡K.�.�{��CC2��H�][Y��砍=�w[�&���n�p����T������ܤNK;���)m��K�����?p���enS��sU��i%����P�.dV�wՔ��c����wڅEI���Av���յ�s�M;�-�YW��:.\*e{��Ԯ��0�[o�����8��^Fe�C�#g7s0������Wi}�T��*˗���ɽ�P��s=�^�Ǳ9����kUǝW[�_i�I�=�Pj\u�8{ɐin|+�qU��W��>��ȈX�W��C�v�cٜ�Oj~���l���[���	/E\��6�k���q���c;��U2	r��#�{z�Y���t5�5ˬjf��������h�J�+B����]�*�s�{�v>�&�+�`�xk�s�u��T����x0��6��i�~~��R.�iؠA��:�j���uɹs����J
>����˺�{��3L�n��hz�![ݹ~:����Ƚ�0+%ƯC����A#��繍Ȣ����e^�$�a�\�AZz��L��8xfu��-6��cS���	���Sʰ�z���;)�U��Vp�s���)Gw��r	`�hy{'v��K_5ˬ���d��JR����EGR�k�yG�i\2��o�w8̃4��f贈w��|�ă�_�c�k�Z������!^3p��wO�^@�;��3
�=�G���>ם�h,���[I.a��%ȯ-z䦶�f����-������i���m�f����}~\���of4�g	u�j��ͮ��w�oص"���ю���b���;��bͷE��a8{F6���N�p�M����W����S��chI�1��i�8�8�>1�Ɲ�]ՙ�Y:ӳeڗ���~wK4���㕷E�x�ʩY���2|����������0��e���Yŝk6����Չ����>�68=�_���B�-���~^~��Y�([P~ޡ.�>��?z���^��P�.
=״u�6*���[b0u.�w���P�[QKߓ[���*-[��O0��g6�X�,c���{�v������Ӣ����\/1+C&�/NExm+�4BT�U�[����ty{���j�ݓ&������㿰��9ׄ�c�������k(��vdʳMv����L�s�Y��;�*W�Yks�+����i5��BK��rz��(ʝ�8&�:�����Ŏ%+��9}E0�n��5.� �B�L�s�KW������s$�_L����^��������������~]b���jY�y��}�L9���ش�嶺�I���\s 7'6�7~Da����Cza9������ޜv����Ͷ6u�΍V&�/}�1���|�rfOM�ģs�ɵ�N���j��OWP��O[�O[�=XM5D9Z���r�ޙ����yv��A]�8+m�xru�)��#ҧ@�&�����
m���{�:*Yč�5��������@x�T��+�i�kò.+(nl��$��K�K�<NC �:�rЮ�u�q�eC�e�ْl	L��'������������o��Ϋ�lV~��F�Um_O���s�����){A���j�V6fl@6ob�Ov=+���D[Wu��=�3O9����sN�Z}7����^�3��@�Z�lߓ��Үq�ӽ�W"�#2�<�D���8-Ųߦs�趫0h�l�u\]>�'�fV����-��h>�'`��nuY�^a�{�vb7Z�Sw$@�s��&^8+u�pkyo�!��M���ou�h�IV��zN߅-���WJ��b ~�.\�4(n]��[�=�y��ԗb�ra;��J��:h��e<�7��R�U�O�R^���V+�š��XV<�So���N�AƆ�_��o�ܘ9�AF�e��Z�r���~�ue�Z��H{9�]�y�s �ɤGp>�Yб\JPer���^c�Šҫ&�F�a�תb�eәc,b�b";�n��]��srɾԡ��S�w�]z�o�N-w�OT�"Ng�iǛ_(x��������5٥d��?e�N���;Z[�S�m���=���{˯u�s�u�J�O9P`ܧ�(�	��B�U�J᳦�7�뱵��g{5JH��*��u	��Id�ja�US����$���Y%j@������ٮ���4��~>Sȋ�<�r�������/��������~�+(uW��ݍ}b�-��49A9[䜋�A|,�%;G����ws9aEP���: �V�6����gsL{��E�9���k�H<o=�f�=�P1�5�}���c%�vmĢZ��O�����(߸�h��+�驯rwfqֶ�e/xՙ}�Y�$6;C�Tߗy�Ç��f���\�Y��o����yo�3�u̧:M�E�A����̷݋��2]q������7�)ʘ��>���ךÚzx�W����jf�8�69��n2w��͇hhX���od�w�kϵ(�v��,p7�U+�p���r��Z��ɥ5��S�ӺӔ*Q�6��2���5�ͱ���_�\��K�ȥ3:V���+��i���i5�]��d�Po
��몡�l7�M.��֩�QȚ���D���k|����M�\���9t�؈�s��3Wy=�=#�I�����цp;Mv��SsQ#3>4�d)�/+�V�caeށJ��ܲ�t܆�h�ڲR� ���MM>�0n��X#!ڼs��mc�2�5l��л�������vE��5�����l-ǝ��W��l9��+:p\��駔�"`�ꋭ�<[�ڗ[J-,��ٌl镢�U�z�]��q�N�,�ـfn�tf��E>�*
!w5x��WɣA��mK]�1Z�3�o�s��bF�7�T�+��"�ټ�]�CZ�\�[68�����qw}��)�v O3��h�b�v�ڸoa��T�LW�61���W�����,�W}����.�N\���5>�
���wEe�Ks�W�f���u&�J�Q|,_m��s7##I7����Z8���r��%�H�a�k�N��9�^ƓjsK;�dM����\0�YB�>�]e�!��O)�=�A��̾���%w2`éVclqyK|0��S.�E�]��e���K鲂�*�	���W�	��C�)���n:Ǝ���].d.��X+'u�EB��6�P�Z��P�N}u�lo]Y5�a{�hd�Dɽ�%'�쿄9{�#`�ˇZ����PM�9��JD�V.���*�X�p[��:��!�]u�7��5O:��M�z��Ғ]�vL�iKoo!;E��v7c�/��	�&(-�<Bo}K�Kt�u"��^�Y�̊��l�x>N�����wgn�:������G�Χ���9$�H�IT���1�R��T��]�_e]cUy��VUB����e`�J	c-)AeE�UU̸��(�d�q9��A�*��eb�cUe@�	n�c"+"V�j�+-�w���M .E݅���Z�X�RcX�(��b���"�%Gt�ݰP�m�j �Xc\f#E1+*&
�L�4�[����kn[1���c�����:�r6���(�&�4��3.+�`c-��J���`�"Q�!��@G�,�}�aUY�넓փ}�(�YsJ��Ĥ��Jw��:�����o�����!�5
�"���K��Ҽ��޵+d�B�+��,~��JUT8t���ܓ�����׏��{'���a��3&��uʯ��F�G�e�:�GZ7X�M8��J{��i�X9}y6�nݯS�:��_��Мa�Rd��8����'���++Vk-�$i�fn��	�Ty8��`n��\8w)\/J��q��v0�1Cͥ�a�CM�6��/k2�R�A�ӕ�1���۳	�7+�B��Js��r����5w���&f�Ю뤰ΐǭ�yv���2Vr�Ɔ�p�u�+��N��ˎ�%2��A�"v}Z�w�G��Ƕ�ɒ{'�rP���WA�i<�EOO�qیn�V&���`ܞ��Zv��j���b������/Vj�.�䱫i��F�z9;�b=�Y��r`ug^�K���t�%����{��ދH��k�G�v���vF�L·�U��wѫx���8���e����]�?��b{��ǣ�I��ʬ���᧪�f4�U�U�F�e�Vz��h�Ϛ��U���+�K��A�6_�����ȥإlZ��f�"�1tp�ՅkgY���Is�����f]�g�t�uiXʨ������r�̋5-U�fϏ����6xT�!<��璘Y�����(�k�qn�4�#�Nl���Uڵx�Y�4�$��˯:TY;�ũ+V+��h��v�˘���[�ύ\dk�\���^b��G�����naq.}^zn�����+)����ʮ����p�e)�)>�`�{�ak�3a#��Kp#/���KI:/sn��ӏ�WVb\FA�gk= �ԶŚ�]�j^����3ce�INz�A��6�e2����"�H�:n�:2��,�G�'s���޽k/\�Հ�dX��P(��hx��rw'b	��ڞc��W�j�"i{��<��iC-��5�w���(qf���%���{g���Qo�s��5n��G��G�q��O��2n�Z2���dqK��oJ��~�D��۞�7o*i�79M�Z����B��X��,�1k��i_�"����t2�+�~4�˲>�=���`�>�_lC�����.�E�R�Yyg^��]�	\ 8�E�ƜYķt���[�;���;\+�ӱ؁�l�p8[��u��K3S�x�|(n�]UB���L�(w�R�i�y�o�*Ρ��n��_7�7�o#�-��N���oP||�[oFj�Z�e��8��l����c���l~�w�hʑ�T�5$L����+3�d��4=WҚ������U�����LX�V�z}%S���m��?;�x�/`���������j�o&[®���s��i�
��Pp����rh?�����w����|�1�#ҋ���0.��c�S`�w�3��=�4���JLf.��������%�X&^CO>Z2O��Z�g>�v���鯡]��pkD/4x��L�/�9���
�HϰV�b���-}J�	�< ^iՔdcz9��v�G�C�}جB�nח�]��;Yx�����+5�����)�Mv�pϸ����=�u�/vcy�(�Z�\���C_:׉6�*�X���k�~Tqc��i��!��v��%��.D3��k�_�w���}i�#4\>u�Ў���kC�޷��w���([ǽ�lVCֽ�i��&��o����h��j����w�yZ��Tdu?z^^W���sMv�-B�4�x��<����y�8ۛc�P;>Q½��}D��x/��^�����{5����yF�D����]t)L;�H�c�J�<�Ι����n�B�'Ũ���d��]!=/'�VVhlj�=A����m1�{�W
��L�o{#�� �YW:$��}M-�Ϋ���!�5/��H������x��T���DK�͜��K�~[����PiuY�'A:)~��*�%����L����	�������VE��J�&�oxz���d��]��YF�gf������;���h�"^f��/���Z`K&�v4�d�䖬ގ/Uxy=������<�����0̳�d��)���8���:������&1�CϏ}AQ�׾���k8���M�bo.������і=��7<����ϺW�sv�h��5eG˖C*���y��1WzӴгq ���HŎS�L�>���<��鸙H��ۙ0_Ws��v6<C7Ჸ�lwl��F�y��9�]�<����@���0��߈.���[�>ͷ�������}Vh�E���E͎U���u_sV�k��,z�(�xQ�f��H'��e��H$Vn��C����w�eq3g@x{��R�@lr�������_�I�47��Q�u<�'w�w�UR�=>���[?Ļm��h����o�]�������[Q��J~5������=!�G�UP�-����3R;�^ҝm�
��L�f��UǛ������u�R�b����> ��'k�O�6#nta�}E|��<���#����L�Hjԡ�vԛ�7�U�8�I���x����Nw||@�P�v���S�a�k�Gb�W��.����N�y��W�Xڙ��y��*�s�jZ{��u����7x* ��r˩\+Q��7��"7��|��c�QT�-S�16(5]t�x��揄ÉQj�
^s�'K)��E����''^�PawwZ�W�+X�,�<�[�(Z�����W���f�l�O#��?��\5���-�AY;͌��|��u�5�2�]�6���ϑ���Lpm�0��b����Z��of'�a[�v����m�	��O���zɫ}``����[��i~�K:����gE�|�q[oh�[h�K��cl�vb��L�󚬘�<�n��.z�g]]u�y�K��@Gu��"��%�J&v��^wd�+�ʙ������i�5��w"(�@�0�:���9�p�3��ݕ�s�3�A�
KW-U��G��z�c���s##D���Ӡ��/�ν6�v��S�Vv��6I�8�f��o�8q�P�VĆ����m6��w�M���-���b���֯&��C��K\$O��n�<0��7�C�ߏ����5��wq��uZ[��Σ�e:Z�g��O&�}f"�3u՘]�-����h�yW%���nm�|H�h7.����b��,*2�����h������M�㣦4��@W.��j�ϕ.D�ma��ޟ�Pn�n�����So8��U���U�>��%'ͣK��<����	��wN�2��dr���r��nƒncs�4�vRrw$���Iu�V콩g� X��&��%n�ٸ������*ugB�P��Η˺R���5#�,��r���e����a�Ua�D;��C_4/xV��Mf��4�e�Tݾ��qn�7mn�d��m�k5���w�v)Lh���3oZ4�}wr�n�8q:�bX3@��(�TP�����&1{�A;%#p���`�弣��)�y�N�yda	��im��m��m�̕bء��WٜN����.CĐ	)TXiӈ�橥u��h��ՑnB�+�l�Lݸ[V1wq.]
�V��3,Prʣt㖄�+dKmf�1UTDE��,*i���Zŕ��6�4�Lq`��b6����%T�(��Cq��Kn2�WaP+�0�dҤ+�W�lQQ)��-�i����GMAJ�Qf�2�h�&1f�"�%�U�*媫�KBڰ[-��S�����j*Ԣ
i�5M�X��4���b�s1�mJ�H���?3���Eoy?Y��A�.K��8.�,�ink(��p�2=g�ކ}:�_�eF�˂OOy�=X0�	$�f��\������g����$�a�q��|�����w$1KG����.�T��e}�VSʩ�=�f�8_�{��D�?=����"b~��W;�3[p_r�����B��[�$��B��D��;�օ��k8��FFX�P��Tv���G��ckE[F�\�z0������f[�qM�kA�,��3����^,�~���8n�d�L&9wP��w32���m<�.�%�}-.�4�ʍ]�W�N|3�^�9b�<��*A��l����H�pm1��X�o�b�0�b��(xs�{Aer�~�i�u�G�4�wH�Oפ�x�g�Q8lBy'��%Z�;*��]3Kc�h���O_5��G��W�g1kO�Vut,�����&�V�����;���U�N��D�����rc#����������(�8��͑z�0�hX�"\8����u�(y��g��$�"��^�KU��V}_]����5�Zo��3�!	;��0�á��.�L�4+ݑ�,�E&e)��ެ�`e�R�v��rI���q:��Yb��eT��	j�گXw36)ܞo��X���j�d�U���{��>�O�����o��m���aK04���y�����	=����p����10�ib="�^��5�1I�q�G��(��+�9ʜ���%V����[P�*���_�8TW,�Y�"�2��Ε��̄����ס�(S��9�Wsp����kuC�q.`�]�`�r�1�j�:�*��l՞�uf��T�i��A&g2��R��{�bڍ��a���4�PL��Kl���O�^N��Le�.'��I��G��i�6*���^̸����z�a\FxkW�+]���gۮ���
C{(��7�ڼv�cՈ��	0�*��.�G�
�g?n����F��ZM�ƫ�FR#��NAw�m���'�d:�C�F�tw��Q�bO)ϥo,�H�0�c�ղw�u�OR����OlO^� ��x;z��zJ���*�{}����q�~~�J,�K/j�kH\S���Ѭ����_'w��Ka
Q�zE��1���HƷ�n-�u���]�
7ǳ'l��
[��� �������6�3�aو��6�$����CΑ*VP���9�%/�ƱV�2a���<���gh��i��<�j��d��n��PV�N��(�g\���WC�vQ�zFU��:5ܓ��}�aGC��x�9t���i&�+�)�{o�_dZ$�L@ۯ8Jt��$J�k+�?��B�hs!Lǃ���ky�8�v���8JU�g�
��y�&��"o�ވ��s��\���Om�*��&U�u7 ;�IRY���;&]70(3�$��f׽�@��Yx��C��O���]�>�3��y��#,d�Y�T7ƶҋd�WL���z*��Z-��3;n�{�:����&��RY7�S+Q'5���RJ��vN[��2�/���(�E�k�)��i��m���ڏ��۬��٤�Cq���ە��e^�(�����S1>Nv���K7�Kbx=:u��U^��u�_�ӝ7y�r^r�Vv�C͜��*L�C̾�w�,����H���(#\��{��<�e.�Ӳ�;����1��b�Ag�sl�WWWz�\���B��m�ViF�N�]��W��~����(�˹�x}:<o��y�G�!pd��6���_.7��}��=(�aƌ�a�U&p����m{K����G;>�%���RХ~ꈕ�s[�mO{�X��h����r�6GƦ��Q�|�
G������wf�ء�G{�Z���U��=�<��47��&'�L+�r�G�}X����q��o���9c�N�j�p<jK;�dЬ+E�F@�e�D��%���Ɇ#���n�;��w8iк���\p<�J���g<IH�A$�g&�=�ާ�:��q����)�ߧ�u�(�8����oXDW�P����{��߰�6�j:�|��l�[x�.ew#�pϱj���"�s=�l�$�<�U�L,W�J��Srh��e��6)O�}M�"V5sZ�3�d㎐^��{�
�H�NJ��s�<�\q�����wZ�HɺawO_gq�(7�|}�fw���޻������W�%nX6���uu���ۢ���;��4Hj���SBt�RXl���)��@92��F��iö0�h�:u��(�Kρ���:k!��|�0f�Vzl�N�98�Sɨɴ��k;)��\
Zm�T�|��C�<*��U֥�\;�%��
���+m�ݳ��|��jv���)����d�O~]P١/<w�0�{|�PHtܚ�߃�1��o����_�'�33�&�[��[|koV*�d*v��OU�{��M{�c<}$b��&�i�_ч2��	�v)��&��F���-d��	LдFR*�y�S<��V�y}�����~�
q��>:�K�Ef�����ut�;����d�g�"<���U�U�ǯ��Y�9V��:Hc؟[7���e((l����D{���{�G��G��<Ofm	ha�F�k���@/JC�o�"����������}Z|�VY9z�� �AJ�������V��л6&�ܜ��n�\������s�(FX��9�w�����z`���{ ��c��jENރ8����'~�hId��(x>��o����ߏB�=�凭U�o
7�C�/�����V�?��������@�?��X�Ub�!!$Ɵ���
�x�A�QWXaD�1!��P�0(fɝ_�P,4���~���Z&�k�=O�3t?�����A$�I	 FBB@I6��a`�E���҂zC@юi6QB�d��J'���DQ_�&0�ߝ8g}���5��*���>�B��Ń�
���C�D:���uJp2g��(��\��qޔT�kԖm��c�W�	���ЯOZ�O��X*(��qT��� $�E��8�ف�M
���n�O�������u�Ͱu���:�@QEr���|�ȃ@5�J�!�E**X�;a�Ũ4/�����L���,V
S���;
�X���pwA�3O���p������آ�(�26أ��l�J��g�!�ʉ!$m�2I<J�6K0���)�B�
���L�0yp6k���� ���[�r2H�8�7�n��w��K%+ϯ��c`�؜�[X�~V ��Yc��zg��Vc���l�1��(����QP8������˚~u.`>�m�Q��b	��S��̿Gc��a޶�A� <�`WEy��^G�17ʈ��@�"��q��<C��Ñ�X2
���
��Y	B4��lAU�
�h
(��P��!�KT�Q��p*���i��z2,�6@��ʪ
��.����*ԛ�,���d�ETV��ÈS��.�L�XM@D�i)�@<bB{���s��ڀ����t�h�I�� �K����j�A�w��8�Ш�+0	�v���������v������|P���J���C��aA��*M�X=:Ó��O4���nS�$����*"�����o��<D�
��`�$�*"��|��d�����xk���v�����=}�����!�������l ��@�ߙ��'55<��M<=�ULG3Po-��e�Ek��'.�rLx�IP�N�؉�^!BC0ټ��N�� hPǪ��a0 �y��;5��E�A��5} ������7��������^��w���]:��7Y�
��5��Ukb�lI@������������w$S�	�R