BZh91AY&SY�:����߀`p���"� ����bG���    @ ��)%U*P�*�I)@�J�UD�	J�*�J%��R�EUD���)B��*%T�)H(�ID*�j
JB�H@R�@�
�TUR��
$����"R�!@R
��T�*H�U(�B��H  �PD�IC��*T�� l�UR��D�*�D�*�*BH"� ��@��R�R)UJ�E$RJDR��P�wJ��J�U   �}
�" (k��j��J�� )F� R���TVB��BH��M�����V��QH��**R"�8   ��PP[0֔ j`@�` Pa�  ����  u̮p  A�� K��@m
 )�\tB$����T�H �  &�t ��.�  :�i�� l t�]�  �p  �>�@�р@��Os� rXS@�P�HUD8  Z����]�  �#�  �� ���Р�lk�: �Wp  � �4)�  V��  ;�� ��T��   ��� PZX�  f� ѡAa� 6�� �.Wp u�6�XA����Z  GN�  UXh�R�T�*�)
U"$�  �  �K4 ��  h�]�t  ր��GZf9ΨMia@�4� �]'p  �*��U$J)D�UP�  �@@�0R�h�e@�w  ;��p �X �&�UXf
 E3@ 1��hڔJ�H")A �   ,�S@6K���á@�� V���Pb` hX (,-�Fe`�4`�*�U�U ��DB 8   fp l�  6Fh�� �;��[EP
�`�6����%���L  ��T��U%Q��   Y��P � l� @T�Pd�h %�CA[�5��   ���   ���*� �i� �"�ф���&  L 4�
JRdyM�I�&OP�4�A�ȏD"x ���24�	��&b���M�0��    BR$~��0 	�  !��)�'R:DW�>@H���W�4�� �xo�=��>u*�]����%@��"���H^��YJ�W��'��k��G}O�%T�כm��zEU*��j�=	T��w����O���ba3	�L�f09�̦a3$ÙL�fS2���e3	��f	�29��a3�L�f2���L�e3	�L�f2��3�&�f2���e3�L�f2L9�̦e3�L�f2��̦i�̆a3)��f0��̦a33e3	�f\�f2���&e3a�L�fS09�̦e3)�L�L���`s)�L�fS2����`s)��fG0���&e3L�a3)�L�f2���&e3!�f�fS2��̦d3)�L�fS0���L�e3)�L�fC0���&d3!�fs)��fC0���&e3	�L��L�L&`s	�L�f2��̦bd3)�L�fS2���&a3	�3�f0��̆d3!�L�f\ɘ&S&`3	��f2�̆d3ɘL�fC0���&a3!�L˙�L�f0���&a3!�L�f0L���a3)�L��S2��͘I��&`s�L��09���L��W29��e3&e��fZ��9ir��S��-�NZY�̦e3	��fS2��`s��fS2���9�`s)�L��S2���e3˙�f\�0���&e3)�I�	�L��S2��̦e3)�s�f2��̦a3)�L�fY�0��̎ds#����09�̡�U�%�$�d.Z�吹i-!�G-�UNY%��a.YA�I����hWIr�.Z��\�+��\�%�D�b�,�rʗ,��S��\�W-儹jK���j���J��E�-e',�r��b�,�劜��-唜�S��夜�I�J֊唜�',I�R��S��9h�,R�9j+�Ir�.Y+Z���9b.XK�Er�.Z�儹b�-Qr�\�K�-"֐r�.Z�r�\���Ir�.ZR傹eK���k\�J�9b勖���29���as+���G09��e3.`���09��e3���S09�2�`s�L��2���d&3)�L��S09�̎e3#�L�LfS2��̎e3�L��S09��p3)�L��09��e3�&2���,��r�妹����n���U�Tߜ��r��P�R�a���"�+����&U��f��Kf���Q��EM��P�j�&�5���J�n��i^�:�r�P�0X�*f�M@�̫4� Y���eNn��;V݋�Iˑ�WE�ܩ���A	X�bue�kͨQ���j��m�hi�n�T��!bG��B�Q�a����ċ�Xkx�#��Nm�B�P��rR�sa��i��4n�7+y�[q��CTt��,��u��q���`��f�#l�B��)����Րe���f�`�iV�&��ٟ1$�&��4�I��jٸq1j�ZX���"٣��N�rX-ѹ2���Z
����I古3b�X�v�
KY��$�TsJ[��Q��*K���at/`�]#�U�`:Ķ��b�R֐�I3vV��¯!֊�̐��b� ����[Y�u֪	Mf�5[��3��Ѡ�d��z>�h�Ӎ��J;��]]c��cۦ�7pl~a�K����)m12iߦ+ĠZmhu#l��EffEWJ��rb:��t��X@W��,h�h�P�tcmhu@���%d�8�)P��Z��Y�q�.�q�Un[4[�Ykknԭ�ŅRH-'Ι��--�V��鹅��z��m��d��;��z V&�{h�u���Y�q�4l�Ԕ����U�F۳�3I$m�k�,+�������QA��=Y�V��۔��rK8i�3"k�&a��±V�g�;O���i���ͪ��)'����Vy�ē�1��PѸ��l����@#"���ug�KhD���N�a$�����@�� ��.��Z�eY8El�i�+Īi`@��-�͍�4��2P`M�M����j=�X��^�	Z�"���k3ݰr�a�ODQ�B����� 6�ҩb�q,��(��t�6�(+Tb�[i�o`S&�D��r�nU�me���P��e����75�%5�2Ȩ�u�Z�N��;7A'F�#�{(r��z�sI*�m�&���/��+E�{�5��* &�םV��۔��I���Z�Ff�ۊ�ۗ0�� �1A��]d���9W���70��*�h�f�s��}���j�c)!+r����P�*��!��ޚW����*�m�T���Ab�� ��Z��
P�Q��Ii�Ѽ�oE�9P�1R��2��,ХkT����ako�
���F�u�Z�f�����(R(I:~I�b�t:�.�l�uiy:�'��.��������P��$��Y�C:��q��,R�PZ7SD�o혩�����bU�(��0�&�!�v ˺b�VQ�JT�������cp��n��dI̹��Y8sM�[����ꭦi�~V�4R(�����L3E;��4��e�3u���� �A䭨�X��H�����SlD6��#Q��wr�k��A��P81�d�.��0'�+L��Aİ��Q�E<qɗ6��9j��{Lm����Ża�O*kj�m��Q�o+l]�J�����̒���t��$�%&�cN�b�x��$��;xl�A�1&c�H�Ӈ^S��#�yb��8u4�Vi��i�5p���K��`�V�by:n�L*��M+R�jZ�x�Q��K�[�`e�QT��4I�u�1�kV5I�9�x�)5&��D��ܪ�Wo(Ή���7I�GMm˻N��>q[2��/f��rR�Afdlk���n�ڎd���ܺ�:(U�l%j���ϻ@�v4&Ѭ,U�M[*=�w�$�R��j^e l5	�����u��9w�Аl��ܱce̔�mt*�1eD�vn��Ų���{+*��M��j/DIM������:"�
d�IX��+=�9���� �1���)�� fS�mK��+3D�ym����V)Ҁ����x;*'Hɣ|�l�&&JK+t���BĘ��#��ֽ�Zu&�]^�.�L q�mx�vՒ��`��i���N�2�֬<�q��f؏�7����b����s��&�h�5(��u�����\���˭����Z5��z�q,J.��d��\��'/U	a�`Ҵ��X��.�=0f�
X��n쨊��$�4�q�X�.�5��M2���J.ݸM^�.ٽ��Y�Y���Gi�x��N ��n�&7�1�a%�T�62����:�&`�R�4*2՘��L��:WY���/*�gl��ZeK��)�m��Z�ɚ��<�顮���7�P�����i +*詆*g��[׍�ʸ�����
�)2��ƷcǊ#�.j��GV��A`N����6^;�o*Л��e˦�̫��J`j�L��/n�8�,��ܘ�V�	m-B
{VY�ɳv�M[F] n�]­�+N��lGX̚��Ɋ�I�ֽ���CT�n�,p8Ղ�n�7���������>FR�#����컭粆�H��R;l<�݆�K7D�)E^�X�l^��\�:�Q1�a�S+
A�3��,��Y��������,G.�`��x�ڸ5$t���1=��1Jн7Ba���#,c"���´��⢯u6F��O('���^�j�%��B[Gwm�uI�"�jJ
P��Rr�=̚6�w�Эaj��6i�ɔ�ȴh�#i��&�����Y�m^�l^��$;L�@��
�f"�,�"ub���h�J���;�m�j��?4���˩JؙwXB���P3u%�[T���F̺t4`J�l�4�#�`�x��%Y���n7Y[X`1��`i�� 
XsMe�L�&�� �� �R���
�Ġ��!��ԕ�.��V���I<�j�n��b�i���6���1��7J魐���PA�-��*Z�%T ��u�]�ֶ�Z�X-�2��h!%�7^�	����)�@���X�&�2��
*��u:��w��	����FP',n�ׄ�A�m]�c,�@@v$�Z�A��%:wc(�w�4b8h=���ٍ������0��x���2�R�\��zj�qʛ.9Fz3����[�i�ʉ��T+,� ͞wҐV�Q���K��������Վ��E�VU�@������!�h�5��i��e4(��mAyt!(�3r����h,��x�
R�?��ښJ�t�L���§�3�5
���6�PR�QKN��pHt����!��,�R�%��V�mj���;h�#�W�5�E���T��>O�zG�e��l�@*��{JC���gP����6Rʸr��1�h��f΁Mj4����4me��b��6�O#*�X�5�J�5T8f�6^�xb5���j��mI�K7�J�e��ɳj�i
+0`/DmOl��[�QJh>D��mA��[�X�0� 9m�=̤@77`O��A�9�.�#�R�* ){��j��-�0�������0�U��K�e�K]�Z/Qd!{4��$�5�A<�p�w��б��ⵈM�ۃF�4S+h�V0dD���çF<2�bEAxn7�v��u=�&�M(�.�m�:��aZ�utqP����a�^��:%�у���Q��ޫ߅�-�T(9����p�;�����7)���#W.
��y����56�mj�Ƨ�T�aT2����`J�0ЫSw-fM�aU��P�"P�ŏ5���HЕ{��"t4�*56ӭd�Mų&:Z�JU+l� ��J�C)�+*���W�MH��f��,�2u*�;�a���ʛ���oV�55<��2:���$�-�n��Uj����${jRCNL͡Z5�����tl[��4e-��b������x��Q�	��Q��m�>ٵ����E�T0+˥Y���j�t0#V��f��\[��Zi�;k%�/p
r��ף:Z�LҶX+:~#]�y��2�R�f����N�krBuޖ�]M�H�gp�lcŻr�!7����ؤ�؉fV]#��H���%��w���x��� 3�P0�5\��5�[[�W��<5�Tc)�hm��i�N%CIu6!�v�
^�v��YyDQ��{��)�t�P��.�V�l�(��`�8eJ(�΁f��2�b�2IL�`dtЗ{�u �(U�V�H��(�^�T�Fj�����@�zw1�U�[��D)��$��ڳ����j:�Wz[V+��/%��Ӥ��IR<�%\+~�^ b{��.���(��B�*SR�ȋ
d�m�t��˴2����ӥNR�grh�5�ͷpIo`�����`U��0K��J�P����;!vX�F^�,'����:�jB�p,���B\��S)Zw��[onЌ����
/׳]=êˠ6H�t�8�@��/F�*SU�Ӡ1��Z�Q��O0P0Q7!��sN�bM��J�i5����cV�֌r��q#�n�A�V�&���/э������a��J��t�w#s٧����@'L�`M[u`�VՍY�yt�ОA�(��q�_[8�Vg��m;� X@Sw
K�t<p�&-�!��v�����,����$Q���<��-�i�9��`��ǚ�A�Lp���)Q������6�k��ʋh���� XVP��,���8�h�30TD��ʚ�-��& 5�h�r�ʀU��
:����U�eVX��)m��{.̢�{����kpma֪*u�银�/(md������l$Sz�ưb�V^���i`����J@�
I��FGX7U�x�Y�I�jؑ�FŊ�FRe,�re��ՙ��x:h�J�mJ��^Lg�#ٸ����ŷ�$�s�"k.C��z��>&�Q�v�y$̗���-e��j��f�ͫ�L�j�hi������@%,&�d��ER�<�i�e��3���DM��Ɔ��{.m!�n�!�C	(c��m&&���n�X�ɸĩ�-�M-EnhwZ�"�n^[�2S��,�^Ʊ�y�v�F����1�I�vU֬�I�U�p���&C#w�^;�� hށ��y{V��� �rEBMX6t�yFP�5	SX��v$߶�QT�Y;%(��x�E�ͣ(�B���R\`��ZCI��6��Q���4��Bj���3Xƛ��C%m�:U�kf&k]@�����۶((�\[gv�5vX&���
��V�(�(b��g,����z��A U��E݃{n��NV֝e�9W�.40�d�4�Mc��-\َ�b3��̂`�����R������ie�wX�j��v���f�04$�-b�,�_���Z�c�w@�^�雓����1m[W���v��9��V�T�E�6e���ȵj4d�j�R<��[X)�b�Į�-;�Sf��XFYg7q@ء�x�;t��zf��J�Ӗ)'�"F���r�ۗ{B+�d
 p���M4@�L)^m3OnZ6w�4!�[ۧL��l�ݓ-ZRK
�՚3U�)�l:�k2ð]����T�l�Ԓ^�U��-�wVV��ֈ0֚�#%n��6i�4v���t�Z`�n1MmE�b�=t�[*�
قXM��Ū����;�d���EZ3�١��EӦ�j
i�$�tvz�-��DIE�����=8��{�c�资��V�� Q9t����J'.aZ�����iPa	�3s:v��D��[�Ԭ�����Y�*$�M���U׬�'��9V�+V�hD���պL�#�͑�I-a���wzu[z��Y�R��(m�`��4��+wl֤p�7t������w��q�C�%�k����i'[lcV���0[�R���4vEt2�f�:�F�]IW�*�SѲ�t���T��i�)F���Mͼ��Uƾ;r�z�J�Z�!���5��f5 �����$�4L���
Fc�f�j���z���
�Pnn�rn�yiL���Fc��m]�k^��䘀��Jn����b��#f�6��uݡ���\`DcQ�-��l�d��]�嫹��njf��f�Bh3��@eKNk�<�J������롱f3z0k(fi�_���eb��{ud��^�-c��o&ěz�b�Ф�܊e�#�"�2���j���Б�2�U�h͎���XU�D�xі�(j�[��܎�A9#�N�/~ nixh��q�
��D�2���R��0):V�;u�d-i�u3�(e�B�������E��]*<�$KA��"K�B�����и����m,�DD�%n�](p&.$��U������P���:1/rD���wQ��ouf�<)��X��r&UչX�V��^��LrMf�)�5�6�V�=n�5q��8TR�ӇS	�a*��n���b̶H��oKt�Yo4�&�ثV-E�o�\�뜪���^��\����:ڲXCJpe$��j�s#g=9LR�ܝ�REU�J,�¸�w�^q[@i$P��V̔�%�i8��!4�xh�r�4��</��ѕ}㫻���Jc��,�.�ִ�ԋ����:	49Gv�N�0�yp��O-�VN
[Iɞ;�6+�WM��vu�ky�Ksn��p�>���G5M'�ƀ�c.�	@�vru<��`ͩQ�Ӛ�m�$���b;�
�{μ�T�J�wP�7!{\ؼ8������8 (�����֖��RZ�n�.����h8 �ee���;��s���.�r��p���[�"�jN��~��@@O1ژ�)���r㷳^�]��0�p�6w�a����u��pu�1}�;k�+��ǠY|�\:r#�<�r>U�J��]�w5�t7�)Yc�mh1�����pN����y'l}�h� 8�ST.(�(��q퇼�A�"�p�p�f;#4�L�G���r�Oj�V�n������[m=ZKc�֊�[2��=yŷ��]>��"m��x1uJX���wЅ�%<���?��������~�>~������*��5���z��V��EF��}��1>(���/��ik"��ˆ����C�o%���`�zf��t�Ϫ�y�)�0>�;n�e+�\��"nV��-� ƅ����w��=%�k�,𩤏��D�rns��'Wu�ox�kN�b'�;.��0]Dm�����`��2{�;]���7Kf.E����v0�T�Ƅ�ln�X�9�v���:	���36�k̜��!в��BR���}�=�k�S2�>	ZFڝ��l��ڛ(@�[�G\e�c��3������.�q&GK4ҳ4P}}�B��\�Z.p=gu"��gF6B0D���)�]֏P���'�g����ܦ&�W��v�-rxᔥ����6䃦l�<2EI�ލ>��{��b9u��؎	���+�S��k�D�ff�W&��c.�����o�mn]ڝ��O�@���,]�� cX$���F���%��O&�DouB���+�8elcJ���CF��3��_�n��Y5�C1��@���
԰y�>4.�p�kx#�ZqA���3v���[���b�(\)Y���f�M�u����sU��V�a�{�z��pYY��,11������ ���:��	%�*6�R���wtN���U�7u�7�����t#]�2�2�/	��^�s�ε�MX�.Vwm7�v>AP��n�P��9�2D�#v�Z��G�mn���8\�豃�>��^���z��	���yL�W��� [¸��2��M"�0�V�����)��i-|�ѵ�q�\j�b���IL"�t��;�f�1u�+��Y�WIdv��"�̣�VfޅV�0<`��p%�����Q��gsGz��'Y4nZ��f+���r|��b���LR;�y.��Ao)�����.�1V�!�9wh�}ݣ�;�NE�hq:S&�-s8�l$u�7"�����Fs� 0����{l��C��;�T���e.Ky�.�YE.�s2iT�������:|��bP�j��@�<�>�����^�7kM5�R���:��y/�.��;镩�2 bm�}��a3�����37C��U���j��$,=l]��%W-�{��zJ縭eN�p�ʵlR��Y��*�ӽ��Wn�B�F�C�ռ�˹˩a��):�%�	��\7q�e�I\�X�΀2�m�0���ݦ�
��yc�[�큩r�Z�W�7�1��]x�IͰ��Z��l��m��כQj�h�!�y�&�9y�B�m�B��;�y+*�+�K��dQ��e��yc����L�*�pYWf¬�e�ފ��84�l<����N��V%�.UɣN�
&B%?(ޝ�v����a{���yZ�z�kw�+����v�Wը���3�����A\�m���~D1���w�/sZ��S��R�o'V���bamG�i�.2<�����L����P�݋�};�����7n��[-�$]xY{z�.���v�=�+)��tˍ�Z���7nﳒ���t�1���֏��pN!��ף���O����^4�A�RK����zP�[�yEn���� yk+�>#��b��]a<�ƃ�о@'�(%+k�� �R�7��,��W0L��eq��/���nd����tݰ $�]��*�/�����7&Iϫo���G5bf���n��h>������ �#���V�vN$-��N 3]s�n��SaP���\����J8پ��2�P��#ձ��Iox{C�W��2���ˎv�'��N�'�~4�Ԍ��+����QE��R<O4����b;7E��W��Ns
����2W�z'kI�J��{�+rE��uV�I2XW����3*D.��>�����;p'z�o������]DSf��7�P���{=jP�3Z�/6�+��Օ���sD)m�"�+F�5�W�)��*�V�N,�B�ZY�{9	����=G��v����7T�1�/^n"!�{�v�n�]�8H�u�X3�ιc�2�ɭ��_";�!h���Y��M[88��PZ~�틻�H�k���.���s�SQ�ytk��t�����`ǵ�k��)S� �R��M�V������"�<n��垺�ndC,ev31`�o�����\±�Sl��C��X&�kWk)��.��!��e��4��ml�;	"��Jk�5Zÿ�v�&�52��	�Q���ֆ81�pdʏJ��B�C�����h�M+Jo���[���n��iRF��-˰zP���}ޚd����yF�<
�����w*��hפS`6��6t<%��sk��Ł�ai�s��gRn\�,���[:FWw*���]L�Zv�n�+��GPǉ����F��L���N�	�5��f�#�]n�HX!X��[�����WyA�͡v��fi֒��1�s7��w݇q�9p+r.N٧��'Os��i�[I����4�UŮ�Ր�n{��W}O(�`ou�eon��L��T�
}W4���y��b
/}�3!I<�3�	�\�Lk1Cv�)֮�A��A:ʓu�V�{��S-j=�s���{��ɱ�u�ՕXdGt�w7���,������;6���u��n����I��S3�e�tU�Z@�����}D��$���S$�z��u1�v�H���Eц������ݶ%��u��'R6|;���uyEܱ��J��)TtK x���[�����cl��+�T1]-7W{��Ϋ]3M�ϴ�o��𡶠O8�ؖo���$��T�ϯ�8�˚�(���.�
T{�һB��\��R�m^ȍj��v���ݽg��V&�6��k��n��*��z�ݚ�"�BUo�oC��t'���G-4�Y�36o��j`G/Y/���a�&���È�{�����\�
�n�iwC+��zEԷv��ī;=ʃ�ѽ֧�[�Z%�J����N���PY�D)�	˶��\�{|�')K)�kI��xu�}w;�ǐ)��3��vd@�����(Wz���S�2h��M�ʵmʉvm
�|$�y(eG$5�3u:��r���WO&�e�B�(7��ƫ��F���p�ת�Y���칽X�5
٘B����Ӗ�՛���_��^��쬵Hi\�A]�6�P4jԦ 
�K���X,��+���ŜDR�_7\;��Kv�K�|��aW.�Z�n�I8�%��iB�N�"�9����	@о���]�;�v�Lg�V�p���f�l�ׂU�Yk>1c\�5{�p,��L ���W3��88aO�����J&��oJ�s�.}w'��kW���>��۪A7>Zҕ���8��N�eg�ۈ5���KMg������K��P�ׇ�d.^�m!P�fG[�C.�C�A���G/��V��*��Z�,i��.�3'rujQ`��[t�����*u�Հ�}}[��
��:��6��}�y�g"�`N ��umWmK�oz�tډ�`��4hu�}��h1��y�Y�Q)]:���o���z(.�Vi��u{�(�$����F�SӡB��6�Tx
�K3kM�3z�p�K��'�>�1�4��9b�Ocf������ڻUW�_#`	*.t��;�5%�;�1ɕ����V�ʏ���Ϻ�bS4ZK&�9�H�7K�2o"��/`�{�J3H��%�lXr�2�����u���+LM�D��յ]'�;����W2];z���WV�m$���
=�1���][j嵱��=W(�6�T�Q�Y}�K%NH5�������7�"*�.��9�+�ٲl�C���$0�nQ���V���[�o�V�l���X�5�qL�t�&���!w��pl�\��8]p��Y��[]ݑR{G����m��C�u�;��VK�cx%�C���yo���r�q��('Ƞ�+aHԣ$d�[���-�X�C*P�sVuh��:M�`��5�r"�����t�ɀ�4���z{7����WG�Ƃj����EFV�?;�~��������*,�^�b�+���Ȳ1wb��+d^��-����Y�o����4]� ����8�ڧG�{���h��<��-�D�9�e3Z���W��&孩sm�`r�#�����;���E#�q�q�\1��E�4
���K��#Y�V]5�v�P�Ǵ�}�]vx"�#���hԈ<�|�E��sL�*��-7]hjZE_P�X�x�жV�1[)Z�.Ն���O�i�v�yiotP��&R����,2�fR���<��ݻ��v���'n�++tV4f���Q��Z鱀�A�92���hf�����#�G�f[�h������Ӥ���D�l_P4ԫ;���2�������݅�5�>e��JvY��,�x�i4���
��������+�,�C`󣙩�ϱ˙:�=mhA��Z��uA�i�c涶TeWHr�̜Gn����;c�<u�
qnx�rwL�\�v�J�:�&�;k"Tv�;�(��Ve�Y���ik�s�v�ZG�g�ˬ�^�X�}� ��jT�1�A��m<b%Y����D�
�e���㙦�h	�㙋�8SVnڳO��k8���\�����6>-[��!��������6��ǐ��/k� O!�vgP��j���=s�Z.7����9�U����ۦ1u%[�i���������ׁ=��@��K�+wz#vxU�:�b�W�|V:�Hǌ����N*)�YN֮��l��wM�9m<F�u�x��S�
7��q�Y�*� ��v,�+�>�ա0��N�ұ�X#-�yֲ����ܻXꜼ�P6���C{z4*��׳;]���G�[��,������a{�VU�V󬭰F��5����v���<\5��.^U��tIGX�]����Ӳ���>Q�Z7C�bƀ��o#�:�+����r�8�ތP��&N���r�z�D��Fa&���7�v�$;�|�*�q����e�KPX����`	�կ';�e4�V�@޴k��q5mX��-�s���*�>��N��]ĥW��wu7w����e����;Щ�u�]	ٹ7@өJ�XEL9X�m�̔��
�h�2])%�ތm���{k���:����41��+=d��*�nIt���++��GCd�9L�g�Z�X��7�l�fh��2j�Ao9��@�ծN���o~z��޴g�]/��7�l�ں�#٨��9EnE�{�J�3�厥̱�/z����72ZXfs5��u��́��$�u8�}�t�ƙ��d�PS�)���J�]�W��C�%���N�LcN�4��3!�"�s�&Z���x����F�c�nC����\��"޽/Z��a���Ԡ��.U�,�;��S�v���W4�v�-aXGl�i�`�I���K�B_J����	�{�v�GH>�1v.@���v���D���$�w͊+q ܬ����a��ݷ1nL��9�t����!kM"{�Y+o5'u/9��C����G,���t��w�7��q]v�e5)R����ά�ӓ��d�Z���:���hU�k��]D����p�,Zˮ%�y+����Bc�歛�bZ�8:�9Y]| �k����Ԯ��#8Py]oX�箷:h�Nq�;��QŒ�����Y\Lu¶�+��s���>���M��hVL�Y����zwF�Mu�}�*��}�S�s��A�(a4�S�1�R}�$����7���%>�8y	��v������:�^Ii�]Ù��0�M�-����R����S�Ci�[�E{7b��������W@݌��-3����6�]�%��.����6w��������x��ag�d�7q��M+.f^cZoPU�T�]�.Н\�;�ӎW [�b������:�O�tn���%v����&�Z��h-���ve1\��#�Sr‪)勚Q"�3_u[[R�-��������=�����R��y��i�,3���RV��]���^󻓒q?�xc�.�[Z�{r�%�Ǧ^Pu.\uv �S_B�B~c�R&�K_-�l���j#�zy"�ѓm��X��������8BL��x���g^p�^hӔ$��^ҳ�l�0ݸ+�Uͫ}���s��ڂW���)ݹ������T��z].��d^6gk]��Ϟ(8��_`�]t�j7fl���G�4��
F����s����0��EQ�}d��vE�]�(�좫JU$�o��4&]
ޛ���'ww��Kwo�ü�������N��=�@N������D��	n��no>aI}����VwQ'���s�����|_wwss�������������t�������������)7;8�:�ĳ�D%DyA�P��pF�Ic@@���,��`���	�J�����]�1��*M�U�B0�R
 �	S:M�������v#f��I��u�� ��:0
�Cj�I��HI��СO�*i��)L:���Rкi 
�V��T�R�B��i٩H�	"�T/ 4؂0E�4%R�8i[�n�
|q�J����Tr�uT""ch"]:֜��1�d1I6�袒 x�>LҍzJD"!��N��X�~�*��fRr�:(��P� A2��Q��R�Fo'RQ �h�J���i�)��T�V0@�*�E �	�,xU*̦��P�(
5������Q1��E�Qa���	�Y��v#�
 q�m��
f����Ed4�Õҧ��l2��� :@�O:�,IP6�m&C&���L	��i�lҤ���R֔���(Pi1�)R��~�wr���������JJ����?������q�����y��^��)��{_�ֆʰ3>��2�eB�)3b�>��^�_�T�u��9&��GD�ӆb�,s�z�_4�9WO�w3��Ws�OB|��T�b�+�A���	vp��H��׼�
�a�K�JPC%��+[����U/�]c�Uغ��]�69��:�M=��q�v�A��]�mUG�Vh
�=��k�ud)�I���Wݒ.��|+�Q'����[銜�|q��%�m����;&����.�U���AsډE{�_lѕu8q��B0�xF�Ֆ�ur��0Q�
�۬��m���[��.[��������Xͳq����"P1Q�vJL-<L�V)I\���d�L(��y/�?U^+�p_?;�;�h�2�vI�`3��T��f,dT����tO2��<�*�l\��E5fX�Up��Y}]v��PE���W_}��C�).Ž{W�R��uD�W���<����<���]�N�ܩ�x�������bM�$�>А�X9��p�:��Sa��W*����! ��ʳvrg������m��-���s��v��R5�{����ǁ��.fvI۷��
P�6N����!O��}�E�$j�AKttī�j�kz������ݪ7�)ޛ���.�F��h��dk5�׫�oh^`6�թ��
�3+m�xj���&��v�ٮ���B�/5����{}~���~?�^�x��ׯ^��z�^�z������=z��ׯY�z���z�������z��ׯ^�z����ׯ^�z��׬��ׯ^�z��z�^�z��ׯ���ׯ^�z��ףׯ^�z��ׯG�^�z��ׯ��z��ׯ^��sׯ^�z������ׯ^�|z��ׯ�^�z�����ǯ^�g�^�z�����׮z��ׯ^��^�z���ׯ^��z���ǯ^�z���ׯ�z����ׯ^�|z��ׯ�^�z���ׯ^��z������v1��+�=e�WI�t�K�\R��M���,�y�Uv�ʚ��	���<��@���[���Xx�1���陂^��F�է�'�dB���U�5�r׵��f�+ �}�=#�}蒋,��;	q:%v���v�n��=��ӕ�ukػ����X��+�Җ�|�N�Ԡ.����e[�ۺ y'U#I-]�J	�wJ�\M���k�-����e�	��:2�VT�q�V<�y�����
�Aj�9\����@�vQ�w\;��*��݇5<4�b�'!���G��5v���GziUĕ�7vL)�{�(ޙN��FMt��� z��̺)�wjY�5���k���Ԉtv���h���^�TX�B��A�����+tjX��4�`���֣�����v�wNp�J��]�n���-Q{+�Y�k�R��]�#1�a7����q7���9{���Q�M7[�CJ�J��*��:��Te);�i���#wv�*��7l=�5G'�C{֔SLHw��άW/{^I�E�x��X���ݶ��衡U1����
y��ݬ��D3&.Z1v��;eX!iY⺦IY+;\����T/fi��pXuj�L  �8�dUg$"z1��u3>ͺwɁݧM��U^���"������ʹ֠�L�j�k���5w��F*����˸�8~�������Y�ׯ^�z��z��^�z��ׯ�׮z��ׯ^��sׯ^�z����׏^�z���ׯ^�=z��ׯ�^�z���ׯ^�~=z��ׯ^�z���ׯ�_׬��ׯǯ^�z��ׯ^��z��ׯ^�=z���ׯ^��ׯ^�z�=z�^�z��ׯ���ׯ^�z��ףׯ^�||||_^��ׯ^�z��z��^�z��ׯ_׬��ׯ^�z����ׯ^�z��ףׯ^�z��ׯG�^�z��ׯ^�^�z��ׯ_׬��??o���<��c���?y�}�h*�u)����n��[�uD{�˛nPtt���uN�P�����,D�I�z���4�Dp}o.��V�f�C9��|qQ;r�ovp[��p>����`�3��Q��ym���H��"�yY���6��D��#�7P�U�5t�x����]V�=���]on��ػ��{%V11η�rJ�V^Sc�z%�ٕ�KT�i
�U��{��I�%�K+\�=/keb���YY�+F�í�mh�7XH,����.�TZ����EҼ��=�)�*wbu��m%�j	��ʰhRH��fS�quewq��f��b�F`.�a+:���Y+�g�R��`5]+���ƞla�Nt)v��靋C,�d�սѻ���wX�����r\�;��؆���X��ugv��E1��:���2l���V�e�3������ۆf�5�Sd������ݹ�I��ԧ5�T ̣�u8 'B��W��M��iE�=�@��@��}9�m_k��]Ri�O*�p��]jU+��D��,9QR�����Õ�z�隺��.ºյ3QK��0�ɼ �>��f��:��+�<4k���׀3�VZW���NWo���@B�͋.��#nU���z��,	�tY����t_c�n��2�Ϯ��wGt�z��[�Ċs���Í`c�����U�b���C\��"!�{Ƕ�yn����j�C;2�%6B��?_c�/�+x��	�B��#��MY�/���ZM���LˑJ�}9�E�����iPyl���+���7-���L�Il˗�^��ʟSO�E��ܰ��h��1s��I���ki��R���!�W�VX�5�!�n�J�1�e5��y�9����ep�s-�o���9KT���}�]`�n�XT�Bu2�����v�P/6�Z�]?8��s��;Ss�Z;k�W��V�.���t�	��pw�Z�3���x�����w���*�6�f"�a�qs%t<�Ú��\�����h���oe�����jLCq�K�U����wl���#m�Sk-rmb�$���g4-�*vAa���ĝS��RR7��}���eJo�[��@ڃmd}�f����<Gv���
F���yF���uoQ�tG�eis-��fQ��m<���pU�3:���ۏ��5����Pޱ'$�M�Z�E��>�2ɚPr>"�'���PY��q�U�������j��]��&P��H͓U:���*Vp�`To��p��m�D���wu�.G�z��PC�#WV4c�f�h�����5���s��	���[,Z�,0�G��v�p&#ɷj��̰��0b�r���fa�[�����ƻ�]a�V ��r}LV�uߪ��v�,F5e��A�3�WA������Rέ����ZFJ�f\YS*Q��;��9����.{b�fv�U9NUT���5�Y8�u�!+u�Aܖ7M�t��q���!���Y�B���3p:8�A[M��wX7���W�{w�f�|3����\G^჆�Y[�R�3�0�
�/$��4�a��ܻ��U�����f����]��n�C�U�Ef��X��S=xw�G�A�����M."��|��WН����p���T����e�C$��[�p�������뻎�#�Ic�i�U�`s*�g�rQZ.�r�=�9+�)"����k��cGX�g��N��i�Ju�uȾ���a��$�V]p��wX��!^�(L��C;�l��q!NJ�>7I��z�w2i��<���.wY�\�n]iu&4�z�T�Hbi�����K�EӲ��h��ɡsY�.��Ef��8!%S�^e>�4G=:5yI�C�E ���G�\����G���s�yж���d��qZt���J�;�u��l�I�d;q�f:����Ȇ��2%�!�/�;�W�{we���Bw#�����l�WQ�K丰��+�@_&վ������|�kj\�h1�t�^u�pכ���+��g+Q�a��G�Q�3ev�2.��ĉc���xa����]n�k�H̝��غ�t��R/,L�w�ĸ6�j����T��ܓ}��}��D�r�ܱw�T"P���>�w,pl��4 q��W��[H��;b���hA@��;�����X�S~�.Au(s���f�Vy6���3y��
˄%}n{��o{�������B��5���<����+���^<����5�0L�j}ce�9Z�p�3���d�n���U�:y��4�)M�Js8����痰� r�s[��0u�z8��78�cMa�*�̧�m��Sn]$�ٔm�ô4a�.)Q�۸ �ӝv�=�+l0�]�8��]B�ꯜ]MfvA@s��+�3Xm� ��j1��[���j1��5ԍ�/:�Z;976:�ˬw@�-��+M.�Ǜ�B��7���Z]��Û�����Pt���� V�F�p��&&R+��|&��hK���|��zR�up�X��Ǖz��!���:p��^Ix�(��[��ܤ��W�k [��%��MYA�E�XE��-���V��_mjS]�4�޼��놼ԏ ���w܄�]ܒ�Q����ҬSk�1�*dN������VVи�+=@n:5��ʄ^*׻����C��t��Hiu�x�bt�b���+/B��cV�c�vOpV#����*�*���rѡϬ�̕�>��V3Z����֌���d��}(�u�!q_H�2=4�$jZ��i�m#w�#�*��.T���m^kA��D� �vZ�N��Ǜ�{��^��i5�kv85<u΅�s��F���4u��o5v�[8�{F _T����N��.�8�����/F�&;����+����`��o�C4��սl4ң���f��2��ZV���{Y�P�ۼm.�wXޠ��X�J��/u�k@���T3��U�z�\�{�E�U���R���/h�,s��v�BoP��2,4�r��H.�������ze�����b{���ښ�4yb9֖`�͕R��S��8�W4�Ĕ�r̍d�5�m�%���H#�y�y�/X�1*5O���ĨM����jT�K�&6�[�	WI�ŝ ��&��3�,}�n�e�2�Zs��H'��*V���x)SNX �5eҰПe�Yd�;OD�V���k�q�)�h{܆�K�%�B�K�k�A�:47[�Sm�L���*�u=����J�÷�ΡdJ�����T@���lI�e��r�Q������l�����(�K�X����JV�V�)˴�2[�r��dW��Sc�5��㚸��x�M��V��lQ�WJ�(ݺvV�oB�a�U;:��hOgb�@d/X��b�zmˢ(��R�rv�Duc�m�]��T+d��Dp̹8��&��"�!4`sxp�lf�6�˲��[O��;p�d1�2)ٱ��d��Q���mmuk���-R�*G{:v��or�]:辯�Ha�邻�m;3���Um��
�Y<�6Cp�ݨ�,�nf�ԸG,l�,���	�U����B�Wu�ʙ�Y2�P������weffdu�bu���l���������׮���BoJ���)Z�]�=̳��j���>�e깙CT�=/ks�g���c�v�䬘%� H5�2��!���V(��l��ًo5�l] ���X�Z���K��O&�[4���H��q��ZH�X1�Z_v>�E���k������ɵ0ڙT�Uf:��s��IL���śDM� /�P��ew(�2�K��z�?SU�c��<����U�]("UN3upVRÙӝ�yWW|����Ux+�Ǖ�h��qVgN���Y��7YwQg�9B��U˺��Vz����>�R����Zue�Kl�<��,s�R!VYp�Yj�
4;�1,���u>c��,ͮÁ��g�1{��\ȝ�+�i�ʘ��۪�7��32̬Y��32���F���:��&�ZY{o1U���qڭwQU�l��g%&.��y%ue$wlM�Ksl���yι�U�+�	��s��<i����[����w��Ԯ���jw(`�Y�QuӰ��h��v�#HV�\r���UvOb�Ɏ_�	�V�X��A�+Ѷ���d��l�(q-tha��$�k�|����G�fΥXf>ƺ3n��t؞J�P����XA�j	�����p+�nً1�	�u�k�R@��}��@��J7�NҚ�����6�H[
����w��� 3(:u��8����;���;��ʔc)��*��ֲF��;�� �OV+U��N��--ʻ JT�v2h�W�k�z��s���3�K�V��wX�*�ݚ�8u-��sk�ƛ�`����{N�3rp�uy��<s�g:����T���Y�^�rc"S8H��B����1��U��`��7�7�o#����!`����XU�$�Ś/9璡O�/L��\kF��k��<�Wz�X�Vi�ӕ=�֍2���Ɗ��l3��K��.����0XMS�3W�����t��9r��� �̬
>͜�	\�
��mcSrD^쬨�K�}�����wb�"݇�����[�D����$��6mY�<0c���uQ��F,�ۀԨ4�hdSC��.2ݷ\��e�w;��']<���(���^�%o5��3m`��U:Өh]Z+rw7N���T�awf����Έ�h�b
�G�f�LG]��]��y����ԯ6�Җ���uWu�20�E5��J`%f	yLV)=\�W/��MX��5�Վ�;-<��{:8 �=�(fM\�sZ�y'U�ܤ���ME����U���.^f���h˨겒��l�(;/�z��	r��h��#��]�9�P�B@3[|~�sbΗD���S�=B���b&���r���i��:kt�2i\ z�2��]�\ -�گ���V�ˌbR@�V
Y��ua�Ym1���m����s^��m��"�+����m�#`\��-����u�(�tEq�:9���F���B�M�M�~G�G_Yw+��tSZ	搨_,Fn	An�����z�ah���#�/Ɍ'W;�.�޵�{\ ��.��;���O-m�9_P��y+E��m��wMj݇��2�p�#��1d���F�
����"���݅![:����M�ī�w�A���i<<��iξ�KjV��G-�����Q!\�.�d�kf��;##��*����ۧ����^�UJ��o��|������~�y@"3J3FF5�THTR#@441$�$*I�*����JP
4���y�lܥJ��2�_�ZY{��
���FsJ׺=QdcDj6���F�X��%J��XaDݼy�eø�X6�x��]bO�;��on�=�I>�1�4oQӓ;`C~ma�pd-�:����dՠp�O��ȉ��P�3:���M��^�L�6�'2�����+�-�S�·�'k�w���m��@';��*{��������|;�*��w7����K�ǦEc-8`��LM��������b"�:�ݭ�*Mz;�^ea���c;�xfC�>�c�1�"N�5���{0��Bts�W<;�(�}��SPy7���Y�sC�4�r�ӻ��W	�\76���[c����Z���:Jۦ���ح���Jb:r�me>U�.+"�ij�˩A�ب�k��y��O�t��*vs�� �c�͵��RҪ�ܣ��N�L��+��� �֟l��S��2ދ�&����"�N�7�rR��ʺ��
�v8�mp�d�
%FJ8S���ݩ']�c�z�*R�)h�]]s���p�7q}�0���L���WP����`��z_�j����K�4c��{{�����#�@(���X���{t,��v�\u1��ay]E�wg_wP˝E��A:�J���S/�C���)?�t���`Q�R`6�a�I�
TJ	(D(D��%�b�T� �*gɺ����f���Ü��W/8itV�HIQ�QM�\*#���Jo<�qы�1���"�s�����z�z��ׯ______^�z��1�_�w�4;�O6�"��
i���Z�MUQO����ׯ^�z�z��ׯ______^�z���4ŬGy�kDLPUS5T�\㦛�*�c��6"��� 5F��t�K`���/9PW-4�Q��QS$�o6��n��LU%4lb"�6�5��p9j�cڤ��7Ǒ��SE5�d�:���5�,�%-L4�P�O�<��h����*cll�I�����5A\�QEATlj����d�%4QE�T���3��㹵'��&	�Q9�{������Q�Ѩ�=��cĜIl�^�.�o3��4�͛k�#�k�E��d�Vb����,��nj�KQ���`�;Z"=y�F؊�i�4Z�d�T��h "ѶtDm������s#A��`�Hmb�cb�yp����(� ��ڱU����l��/}_8غ�|q�7G�_ftט�Qq�}P��fA�$����R�{א��.��Z.�*4�c������f4
�w@�V�0f_���Z�G�d-�t��!Y= d7c0�W8��H�C��n}�����i���W���^�m�~\�N��G�]�얱�[c����ϖO�`�֫��}�W{Ǵ�}�v�:�C��P�仸��yK}��T����������A�Ng����3�1;|�ga%>�+c�}<��k�-��,st-�Vu�~�]_TT=�3�؍N&�`��n,��ӆ����c��f�{o%���w�0i����; xWN��C������oY}�3�;>��C��}'�懠�;�ư`�<겻�Uv����^�w�{(�eE���;�Ư�ވo�>S9��)Z]h����]��5�wl�zlU�`�h���>���W�U뽸���ݙ�M�ϼ컧ؔYJ�c���o�5���.k@���<�n5Ƚ�����3>��n{F|�_�Q���m�N��'X��<���Γ�R�0�M#��Kj�)��;��ɹJ਼�v���J�z�g��^�W��c��E��I��z��i�A=]�����gP|Gn�����O6jg;�=�uz*�"H�+��uz�:�j�]���;7�/��r?W������Cu;'�S�~ʃ�z}A��׉�N�s]��r}�s������mo�����:��}�)��e�W�5K�[ڶm��s���}K�Ǽ�\^�銮�g�]�Aݮ_
B��yv��L*��y�j�������J���m�>N��������W��G�e����E{nk�|��y=��2nj�k�����#�}cj>�C\Nzy<G�s����g	�.K��M��C&S�^����.߫�-]^�ޡ_|��;ÎZ��=�p�p礞����]��}�������̡�Px�p�����>�\��J9��vx^5���
��]�v��^��*~��+o۪���2���w�!�A2>�n{a��f�9��^�v�>��#�H�y���]�>ӣ�o�z�_z����v�z�"�;ё�fQn뮎���Nuyͯw�:{T��~��� �-¯��4��Q|�@�Nm��f%*�^;;k)R��M�]re1������Q�tW*�9�����-ȳ%�7��of\8*K{�o܋��U�u���Z-՗��ߞ5:_w!2��'m�Ө���;�<����� ������Ɏ^�v/�k�OP�����ބ��מ)������7<C�Y��^�_UU��}��V^��<6dy�c�n��^���#7����}=�sL�aҔ�o���:A��ug��U�/k>U�#@�J?wΚ��f�پGt�I����w|���:"^߳����,G(���K���.��z�#Rߥ6�^��˲Vj^���>�<�2u�EN�>�DGwq������Gv�27�n�}[�_O���8N���q�چ�xH��޽��VSǶ/6	m���"��x`EH8=y�N��>e���յ;����R�ʂs��E�_ݛ��A���b�z���ӝ7W����8[���:\wm
�xF���j�}f���oL[��Y��>�nR��1=k�.+�j���g�GDؑ�0;x\;mɨ�'�dP������D��W����:+U1Ҿ��;���p�7�-/���u���&s����237�f�1uJ�}z��Zr��S)N��e���0*j;�ym>8zt `�
�Y��'��;}C�Av9����F����wb�"��9����֯��{���/�w�+/��״��D~����K�np	U�C�?J{]��d-�����F�����J��O�p^��MG^�������y���+X�_�ڡ�N޴���ƞ�ѡ�g�{��R��/�S�ǔq�������Wy�����U{)\�[�:��� �ןsɋ�[Bz����+|�i�6��y������[���߯+��ʽ�c�(=ͣ�b�����C��WQ�ߗ���7��u}��	U��ùq�~�����AK�g��)�=�v��H:�#ҏw�	�yJ�{ĿW�������h�>}�Fw�ä����Ao���`���NՓ=�_x�3��|���S���>�I����C�W���__���{��h����t�A/%S��ȧ��ѕ���B�������[�u��7�w3�k�\��]�}UrM̝��*���+������Փ�����(�g�_1�2�CF�e�����w�捕�HgE.�̨���&� ӝ��}]频�ίM�,�RY�U�AC�'�j�j���މJ��٬��Ö�n��u!��:&e$�d痖t$Op�c�wYES�>�B�]c'�X��7�1~���7�b�e�(�@AP$�˭����J�e�9�j�%�X$�T�*�R��³�F�l]��\q�U]uV�~��;kfb�q����9��o�/W�^�~����\��_������*�c��˼�<���0n�e/}�|�vA@��2y��x_4)}|1w�Ξ�y�|�Ufg?F|��B(z�{�_u-r�w���=�?�:\�X��]�1��lC��!<�vD�+_�]�2v��xvS:Y�լ%��x\�`�5�*�������dK��5m7��4�W����y�����+�/�T��^���m(���Z�M�	�����SÕ�����v����J[�ٝ|ڋ{�.2�T��l߳M��<MW��o�mA��{̹�mnX(�(߫n��GI�QEw^]XB�g=~�䶻�wOJw�j�>+G�R<�{k�yV�ҝ{����.����3���'=�7���@8�������]���5w�tl;˓1��b	릤Dg�>��j���%Nd��{���N��%:�^�C[-V�o�m��|c�:���	�re�䋭��ܝ�t�رbF�x{oy³*��6�V�Tx�R��y0�Z���P}�`�9=]]9��t%k�/R�w�+�ʝ	ytÂ�������IR��꿻^����3�Hk��f����\ٶ9����c/��y5����,�Q�g�w`ڝ�����D=&�)����x^���H�w���s�<\랼v��;^���x�힃��3�Ǹzu*�8�~�q�Os�ɖ��P}o�:�_�nd��Sv��z?u��I,J����|������(E�|�^� o�:U=��o�^���jv�g���q|ϫ����U;hUl���S�������=9eGξ��k����:5�`�����j�_o�r�v���]��������g������w�f�h�*�"�j����`h@�.�xG���L�M.>~��}��gw=�K�|�5q+&����z��N�"�Ʒ3ϱ���}=��gO`+ �-�<=~�<�Z}�߾2�u|�w՟v�j����W}�xa�~�t���eB�m�4�������|�e>vz�L��U_
n.�}��Hb��*gVj���"q���%M�6C��:�Q�l��'Bk�M�m�wl��t�Y���\K��;�' �V\�WxxxF��뙑�S���>�����-H���X���繥����I��w����[�ϣ���w]����Q�x�Q�<j��/4��j��L$���:�R+����v����V�7�[�U�6M?66�����]-�y��g���3<��[�.�y��ϝT��%^����_������,����Z��ءa��z�7����X�p�m	��Q��y�}:W�k����.��vR:��%!ro^��C�6�gTOK���;[���މ3zD�s6v�7�R//v�1����|�n�eǟU�[�G��ϥy�Q|�n�2%k�&�s��o����q�=�{���0 ��3Y���`���������<�nļ}�t���r3�̩�o����Q�/&׺g���T�<�.�}̢^{q�s4���W^�o`=��އ���o��N49���K�lXH��*WY�w��&�5;������?����_R����H҃戱h�C�g��U9�hh�A-�S>21� � �d���X�z�S//31Кz��
�v���W�ձzz��-*�J��jç����d�}Z�<G�q��&Rzn����){<<<R=w���d�w�w+��K��y�T�W��Wt[�{�hG�=��m�9\s���v��+�P�h��J��^uu|�0���6�?wT��Z���h� a���uM��;�X��z�a9�)W�Ȃg�GDئ�]�/T�m���=�\":<�F�x��NzS�]���nj�~��v�G�⣝Og{�}4�ת��ÝI��>�Z� d�]��_{�uqyN:'�����c��O��%��ڣ��}�>�~�;�j���V��qfp&���o���y����f���|q��/�S��]�G�WoxS����ޯ_�z��=����?Z{z޿X�=C|�X�j����{ӊ�e���w�#�����i��v�Va���3����=Z��X���m�#���oW;�=�/b~��ݩVD�k���,������1g�u�n���V�fЛ�vs��N���Ô�_�ϥ���ŝ�7�=P���]X<n�%K,�nezIc���|��U}�]��R�I�@�Z4���C�;4��?%�FfG}:gY���D��h��S�ԷS���/��F�6{��M����IT$P�J������SY'�9����F�﫣�>� �z\s��Gx[_m�
��@znzvz20�x�b�'�z?x�T��Oq�F�u����b����`���Z��^~~�9�Q�NX�/3j�Y��5�E���k��ų�������8�'B+��]��]��T��������Č�s���y@w���|�s�T]�M��0�S�vP�]�ڷ�L�;�߳�.Nfr>�ӈ��h s;���M�ꩺ����U)���<�=�Î\�ʪ��aS�,l8��j�!��,u�|���w�?oz����"<�+Z�ղk{3�0������~}��wꦧ3W8xX���N��^j���{je�Xf�Wc����0x��ҹ���ڔ*U4~�y�}.�S��q7q�=��4o��e1q�4�c��c��%�,
���zW�Pr��>���	�@}w����BY��Ϟ��wLT���^��M'>ٸ��}�����]:�ÀJ���u|��j�6v�d[��i1N��뮫��]�%;��Btu
��UR�"�MzFN.G����·�����ɸ�vuv��g��r��,)ܸ����B�d�FC�y�+�l�q���_
�C��«.�I��j]�~�cU�P��M;���_r�=�������Q����{K���Ǭ���$z�HUdLP�ʡv���}}�����(��Imإm�zu�˰���ӽ=��%���/n�hU|����]Dq:5�nrO|ؤ��,�'OQ�>��{����/�9,��VFw���:�?1� /�>�ʰ�q2Z�<�m^s�s|Ϥ�������j�WW��s�DW^��#��%sB*>틟ngz{j��tC�����s}px<{2�����9P���׎������M<>��+��}�H�4��w�:א�u	�����Y����g�|�}A�ڦ��w��\sP��;���U��]�[�Y���_p;��L���9��y�Fd}�i��<���3sǗE�:���{�j���[��]���,�};*e_�Η�P�xx~��cl�f�i�]UX���w{×6�Vy}ѳ�)��+�I��%i6�F)�nک(�B7�&m m�m�W�v��b�J�����ܭr�����:�#F�U�藽��5�;��w�॒���s��b��t�]��.wbN��6�o:�z\ܓ-VhVՖ(+�6���Z�;쎜��3 �k�$�+�Q}��釬tְ�I۳�0C�X�-�k�<;=��ZTX���Ǉc;{;l����Y�w78+5�*�K޷�aE�'L�C;;y�P|3nIs�*l�d�(�
4���C3��&�e�f]�������b�/Ȯ�r��a�=�Ӑ�U�Uŗ[�FW��k�ՋV�(m�N�p[����B����ks�dN�x��i}z�j��"��%gCY趀���&%���;2�RX�M6�wu��u�n�,yWt�Į�qyw	u���\�*��/��)F%;M��G��v�m�.�	6�5�o�&�4RJ�	m�B�[�{W�S�Z'yܤ%����7��Rb�$]��N�-)�\�s�m�8^�u�p�U���J�V`U���u�l��'�����d5���W)>����7��U;���>O=��Q��������l�e��M��u;'ub����T� ]�5��	Ws�X��[�!ҮLP��;��^�.�Κx�޽��7����u#�O���].��ɣy��4����3ٶ"�y+b[J�u$����2��P�{��B����G!���9$���ǑlVw1o"Q٢/]�VA2����s�̎e�Ww{�"I=mwG�"9Ӽ!�'��¨�Y�:�g�����u����f�ܺg�o���a��ml�Do���u)v�����r��i�����+U��h��Q�h�\N*Y�/)Y;�('���nRw�i'Wn-<��Z���yƥԿm�RWi9����6����z��C�jZ9�T\�	2Q��bZ��Uv����o:�:mQ�����İg�m�UF�ť����X��.��Гg>i�͜X���M�!k�=�����R+AC-�n�wZT���Q�X"�v�|�wEE2�v�fnhJ0 �-�i�43Tޣڢǝp�2<����Má����nv:)"���-PUt�191��v���9�w1W�]�
�"��Q��!���t[y�o�Z���fS#�f'�}�#^Z��IG��F0�i��ootfv�һ�v��ޏxg��.��4X��s:��/�l lOe�Y�2�
(oB�y�z�h�Os۾�bΎ�a�a��d̻ꓔ�ը��|\��a	k��6q�\65LӖ��',�:��&�<b�^-�] :�Z����Gq&Wo��2N��RP��꫺��-���m�ѢM��R4P{�s�P�c6"�V�9�`,mD?�5G2�vm�Fғ�6�ڳ�����������������ׯ�����^�z���~�m3��m���:1h�����9#TQ�'G��p<�8��k����ƴP�F.D�<~������~�~�Y��~�__���׿H�h�U�j"�ss��i5����J���14�Kэ�:*"&��61L4A�f(�>ܚ�tQ4�-5�D�y�PMA�֓^^G��5�>\�=��4��3���Ul��j����*��-D���
i
)���R&�*�!�JD�����ZM��IT��y #��r��Azd��p��Z�+IG���i��9���<�Q�$DW�O�(=�KATQ�ll!��/6��6#ce���78bѡii�h)�)�s�_>p�O�Q�0RU7͡� ���߿&�n{'d�
b�s���<	-܃!�a����*s�܏`f�Tr'ۻ��0�SK{	�_�~�������]x۽v׍y���c�t_G�@��p�k�4��c�pS�O'<DX.D���s�����#��#f��f=�Q�sOY3�և�HT\�&�ςؐ/�fex1�>끘u����'��!����l��W��bw��t�#���;�L�T�O���d�AU��i�`Ϸ+���)t v@��aD}yp�/sr�.�f��=�%�u�=7���w�������P=��8��-خ��G�]t��J]
M`��~�v����;8vIn���q�����D (�w>��]��@�|Ɛ.�
lx"j<y�2ȨY�k4N����3T�����CS�xȮؓ@���ȃ���4}]�lPK( 	t�r�����dJ������d͖���޲��e"�[�C���5�0}��6еNO�)�kI��x�Tϋ�Ep{:�yM_��z�ju��5�z��^u���p/\�DO��Y��$�|���[4���=��A��9��򷇯�}�Ű��/�t�'��Mk��
žU&��&�z\`i���O������8��/�t��\<��P��w�N�/d#��B�- �M~�Fkj��Z�G��ބ� $��i��>*��|�JIc4o���w�kOl3�o�4S��j� 4�-�ؕ6%�sڱsrC�;�����N�c�	�.q�p�
:0�H�J���K�C4���	82�5u������Čnǒ�7�,]˘��;s6_x;�b�W�����^^^@3]�j��C�G�e�z�G+{'ç�������@��Z@�oT��h�P$�v�Wa�
"�o� ���j�v�7� ��XG�����$]��Y��l�~y���=g�_���]���kc��\�C�9����L�uq�3�ܔA�P�������������s�zWQy�-���I�cm][hAe�g��C�Z�=n���:kf�&�Ĕ���)���,Uw�R��|E6�PS��kLWU����N [e��c�J�4���ԗ���k�]xm�|����E�\�洵4T���W��C�.��Z�̲F� @mhhp�ô�F��)��=q��v�y���kJ����|ӵ�����C`�K����_Zu��R�#�@��La�����=����ыu��tu��W������t�Z�8�jT��d�J��@��C��8���a���S��a��Q���j]��-e��p�e8���_ӗ�W��9����bݚ��g06]��]�N�Q������x�Vep��įK���>5���`,�z�=Z�)+�9^�8D���l�zvC+��.ɻ:�n�v4���]l����2e!CG�i���%K���Uu�p5�+㨺^ǳ���ٕ�PEz�E2b�)�xQI��?H/D��:��p�ᙵ��b�wk�'��q�)sz{�#���	O�f����yv�e��4�+|���H��!�>��^�9�������1bzO�����ۍ�gQ�=z�w��|;Z���k"��Ȥ�+���VRS�·;��2��N���^��z�ݏ��s���	��r�����QD��x�K2MZ�ݍf��*x~FWot����C�7Z��']����l�b����c������oX�O����l��K_>��j�ײ�y��m�&����u��'ڀ����齇�n7M!���2 n��nD��j�%�6hC����.��c����p�ϧ��;�`7L"���vyB�.U?+�h�Tps�������w�V!��^��G4V�	�ޞv+�N�E �@W}#V;Sa�lbċ Y����ɸھ�93ݵ�y�۳[bby����na��^��*ev�k/+}����Ն��g��ӡ�3��fG��'�i�;���O�v:s1�n�y*<�BD��Q�~�����Y�*�[Jv��a���ٛ��M��b	f({������}������ϥ���@a����	�Q�a�c��1���4���b����y8�>���3y�;�>�	^�����j��|�O��l"*|^��\�2�^T��|0�߄t]�c.X��Y�c��)u�E
�2�:��"a�K	���^�r�ۉ�М�68LMT�i���b���R.�S/^���n�m��V�p)R��ͤ���]�M݉ooWQ��{W[�{��$���B�Ea������{�w������q����ڮg#�8~�q\�m�8�{�Q/�g����)3���w�87���|�2���F�I�g�T�f�!���L��S����s�ܘ'�A���(�{z(��l;c)�\`�i�˭i�F����mM4�C���'j�	/]oB�ʻp��DvZ�[�T��0��#��M��c73���4����~C��鼼�~��-��e��7���`}�0%�ly��4k���҈y>���U�D�ePҳF]�{/Y�M;!�h.)�.��f�L�h�f�&�.�e�0���#��udf�)����k�1C*���,���=��>���Ӈ�]Th�kF�	�U� ڽ��k�W�ޓ���dU���*���LJ���U5����钧_�ؠ
;"�͑<��U�)|�0_:�\��"�������%�T��WV���x�f�x4{Tv��tD�IDR�sm)���&pi�<�S�n�,}�(��@�nmVd$�7ټgj���;+�a�� [�.
��ќ�f�F�Ss�m5寧g�B���bS���E�l�܎�]�����N/l;��_�
�s��@c�P-B>���>;�u5O�˝���p�Z���I34?C�7;c�a=�Fi��E>R��4�QVe��aܕb��V���,�3Ǝ�JZTi������)Z�<�{��eKn^lPq��<r9��mr�.o4�&`]��tNB�s��G�;z�Z33��\�Vִ��%�U��j��x_������?� ����h8�=��`�����,@-��HϤC��mzbU��'-ta�\�8�י������p�hz!��k����+M����7���;�O>�H�4i>M0�pǞ� �W|�Er����7���� Z�k����ݾ�)���`O`�z|�4�t�H>yasO�������ә�fU��W1���({L�-��g[$��'������6'�������t1��w �r��gRop6[���Vm����} ���4�8P;��>��C�aU���P,�6�s%��C�"����be�9~M�p�5ʶV�F�v�V�zN!M��/�����Kȶ&�U�$����Fa����'�`�"j4�顷����������fspV����0"^�]q�/�SQ�����7���@@�k,{f�m,K�s�n(g�=2Č+��`4,�]F�N=;:oH�X��aE��5z%��"���@I��k9��/�T��C��Y����c��;/b�'y\I�m����<5����ݱ��O�ˠ4:VF���:w�|��Ty훽���Bh`�L�L���dRx(ͥs(%���l[3�#�n�DQ��'�w��S���ԩ-%?tC#��Ö��"�_��`M�Bk֢Sd�R9�z#��崠���o-�!���|t��|��ө�5�oP{�Cͥ�frZ�#b�z�l��^������A����rIӕ������,,����w�Ar8w��~y�����ǏQ���y�<�{�L������vqeMa�Xw��>��p%0V�I�J.�=v�:�9���ze���
�0���t��m�m�p�,��F|�a�[�ؤ�Db~֯؞��i=q޿b�["��Ka5(�U �
�i^�К �Kf�a��e�F��g�s����$�-���q'�Ý�o9��t���c#�N'8���g��rB��#����YYִٖ� �g(ǧ��X��P�݅Zv�^�j�Cύ�ڼ[������yֲ�P����E�f��>0_u�M�35��n�꺻ӭz�3��r��f���T(i�>�>��R]V_��y՗�s�{fc��>w�末��'Ce�s�#�tΡ�9\�ZS@u�$�wz8��},�U��Wt�c��{Cl�{']3�F�M��;�f�������*u��[O3g8�����|�E�z��:g��_�ƗS̄n�r��⇠�h�bS�����p8�V�"���/֪�_O�ׁ��i��_s'�����C��]?v�=��l��4=�W��w�*���Q�|���g�~<��	·ّ��Qg76]M�c܂��83������R��"�Ń�͙u&^]ۤ_,�����rһ�ڣa$ZW]E���T+{���A��jP����;��l�8os+��u�����gz��h�sD��j/�u�c-�u�ء�П��6.됪z�眫���usW9����<�����S�<PT�ߗo�|��������t��y�8,Ѹ� b���g\Q���Y�O�����"��9�z����u5����0�|v׉��Ĳorw�P�V^E�aZ�NI$����uR�<�u�����Ə5t
����X3��S��������(=?��t1M��˙x7��Jطf�QN�ce�ۤ;�U�#�!�Nܫ��۾����m?x�";q��8jQ�z�@��WD�T5\�NV��$�.��-��0��j�����=��oQ�u��ͯg��ɀ��Ҥs:6��⵫֞S��oH��Q�"�@�����]�١�솊ak�� 1V�@[����,˷"M	Qg��}�:Ρ�a�qc��/Q7��-��_w��h���6j.�3EQ� �B���Qf]�ȸ���ql����!��V�C������v7h=m��=����/��w>��t���2+X	�3ͬӦ,]0�B|�a����Ǖ]�K`P��볒�l����J"v
�6��Tˎ����0�Nk��j�gp͙k{`�*��bm�Ї�4P�	5�Mb�t����aԧ]= qZ��l��Y�n�b۾⥺��z�a
�3��m�{1�4�_��u���q��v�M�+���4x���B�h��a�oq�E��f�ݙyC��$�V�`�)����s���Cl�q�>���Ϲ�r��sh�믞IJK����tP��GF��'e߹Y�Eʕy�?�^_����W�<D?|������?���8�����}`4Ȉ~�U�k�gP�O���/�m:jX��.�G������Q�={g�R�.�@^� �k�Er	)��
�Gz52�O&�Q}~�� �� kS��\��y�n�kaT�g�;f�g̒|.�Ea�],|KD����჌tC��a�|6Ț(��Q�����%�
�5;���^���<�����h��izl�L����=�s:������Қ�v14�m!k���obǸ��לC���ڣ�*ٽ�v�i=��ρ&|꧌�z��r$��N?��X����ܘ1aDv]=V�a�aѹ�c��4�g-�6����x@����oF��y�4;k&����\?`��yy��An��P���\��K�n8$�~:컼�w�Z���-�v�����9�qzP��yː�ñ�6�Z���Q�`4`�֙���	L3꽏�W8F���:����������E8�g��˩����"��p2j���G�v'��t6�r�q�ue?KP�U<L���3�<sm��bԵ�ri��+��dz�;@����<Naf ,U1�}埳ʿPv�.�Q��X�L
��g��oќ�a��j�B96Y��\��$����l".�NdeY��C���T�8h�b=-:�'�SUڣ����-�P�a�#�lg8b��fۃ���%�&���Y�#�_tŊ�y�z����߼�U����� <��o����Cƭ�qn>��z�	L�����6z��<�9=�8�fR�����D[��s@��ˣ�j�{���ہz܏��Z�5�9�mJ;ؠ	;)��{vzp�4�L�Sʇ��LYm����e����+ݛQ�>{Y�����w��7S��O;1�N��qi���t�
�/oI:\l%Ի���cxK��#��ǲ]�6���n�oEZ�(��bY>#�Φ�2~�Ňy�S���?�̨�����F����M5�V0W~#�m@sL���Ъ��%�_]Fƺ�d��� ��5�4܃4q���vA�����C�l4|�8�w��Ο����k�sK	m�o5�F�3/r�.w���bW[P��;�Y���Wf��\�1��j`��h� ��_ͽ8���1�Dr���vU��%���Z�� ��q�1ɳ�Ǯ�=��@{�����L�x�����ؾ�S�&1G�컇���<a���m�&=��m��@�\Y���i�Āzw�٨w�\�}g!�b�~�[�������rxsqs1�g����_y���܆9��3���$3�Y��OT&��4���F��T٭116�_�l�]���]1l�܎���Χ��S}��q�k�se�[�B� Ы�U��zr�;���k����<a�s��1�Hu;b�w'^bKq���0#�1���~��{������ǏPO���G{y@-�{��n���Ϲ��l$���A��q}��Fe�c�Wh��w�L`���3.�=If̬��y���$"�K�ޘt�n���w�X>���c-\�lK�f=5.Gt���z&�g�5�T�\�� ��<�iA���N7~�����E?g��ە	��_�#�_�ߝU��3�kV��&���|���Ȝ�C�|6�
�2���<`O8QT�̜��ea�
�����;��!���8����ƤzmuK�N�XT�����dSh�yL�^.�)7X�q'�i�J�V���������2�6����5�k�:(٠����p6*�a�n����+��w��N)}�/.���p����^�f����aC���q�t}�.aG����ɧ�j�4��RQ�Gg:�s����]�7d�c!��{e��6k%k$i�F��bV��Dد���Lg��8;(~�w65Z��;��u�6m��;��8춟a�}޾�O��$i $�m�p㙀;ia����2���t��{̌�v;ٝ_Y�gn��},[s�l�.�R�m��y�����w�ÿ��k�{ȷ�5�%�#����hStaG�ݷY1�Y�09".�vvs!d�b�كy��&�bL�aU��~�J;ky.���$�fS�/���� ���.�U�*�)њv��F
�M>�9�e�N�܍�jJ��a�N�	�\
��Κ�B���w�b�=W��H��m�ru�N��uf�XJ,��7{(���a�}5�_X!6֘���� t��̔�h�P=��Hb[;b�Y/w�����gq�2�8)��3+Vk�K5u
�ƣ&�rľʹ�v�YF�+��k��*�9\}e`SEK����AcĢ�c �]dt|�j���C۶�k@%��f���B���M���6���
VK�뚤�AB.���%�ޗ�^5L�X��)���lg+��x�T8䮅 ����|��+?j���w=3rh�5����\vS��˔�=3U���Xa�n��G����)h�o���iߒC)'�r����N�Op$Bvq�{[�$3u��j���=X�ʝ�����ER�.p�D���T�|��ڛϣ��W��%��,m
Uwl���	���qT�Wc�� R�\s^�wX*��:���K�qP\8�K��3,	
�_�k@[O�m;�A��4���bjcx�����`#;�j2�Od��%9���ڰ ��y՞T�aA6/��J�wP�Ѻ}h��p��j��v̺��t�f��V�7�Y��.0] �a�[NP�AJ9@�w�Vץ�j��E�|rDm�������,R*ل(����$�b����4~�P	��ج*y�}�Ҍ�i����l���b
ݲ�b<�M򺎸ӭ]}3!S���+���:�2��r�����Y�z���]9��qZ�x�D}��^ݓ&���Bduͫ�l���췍��
wi�[�.��ͷ����e���z�u5�H�V�ڣ���'%�U���+@aJ.�V�l˫ep��Q,ZU\s'	Md�Xվ�B��$wE��Qڬ+�#�D�ۓ%������ |M�8j�"���!�N�œ+��M�B�'WW9�c�.�.�ռ�Fs�?M�J�X�0-r`�I��%҆l�w+���]��&��4%dν, ���ڽ����p6���죸�ڨђ��`�5�����zvڒTuewN�/u��w<�y�@o�ɚ�[�ԧ|�"`0����/A��u��w|�����t�p�|�-�'FfP�q�]=%b�Ra�t'o.�}M�]��;Wwh�r�	�+�h��i�[Bp�n�<��c�	����d�����,�Z{M����8,
g^LU�rn��!!ݝ$��D��6��5�if�w[��A;����έdP�A�Ⱍغu�coR)�3�)�ÛL`Š�㺺#6�g���6��髿	YY�u��<Z,�N�a73vH˛#�&��޶�붔\��:/oA6\OWG�z�h��	{����{�f�𕄊�):	�Z�i�A:��E�-6�lW�J:%� ��E�MX�i4-XqE
����vn0C%�Ca��$FҔ" Jf�*De��ݑG���!�4G�5��E,ƌ^F�bb(���QDD�>���^�_ǯY������}}||~�_���Ҡ�;"�b	�h�m���*bgmQ��1,l�]H�Z�9��z�����׮z�����}}}~�_�~_�_����QP4U)AE!EV�-�����>m�j�)��i�R$�}��N� REJRPE@P�AE$KQA־Hx\���b���J���i4P5UNl6�4Pit�UC@P�Ѡ����i󚂏7��Ӯnm�V�h��gM&��mc�5E���ꭚT�>X�(��MitRV���i6sZ[c�	�j��{��Ѷu��h�*%3�[Pb5�Cm�M�ǒ[P{�s`�֔�R��{�G$��?~k�E'��^���ݧ��wVm��V��0�T3E\���
R��>�P�����>�e��ʶ�q'D�j����4�B�#�m�"�`�%�d��LP��ǯ��q�Ǌ��=�������~�&�g/l��zZSC�G�ϷT���c���}�W�z� ��.��z���G6V����jC�p��%�ųX3:���ҙ��e�lt��Q�"��c@{�<�:�(�I����?@�C�M �2���-ܖk��qc��em��q���a���:Ǟ�A�rĵ��P˱v�d<��G!�}�Hة�mP����r8:���r�V�@n<�ɳ�.�՚��y��"�n��̜��m�=O���Xͼ��(r�Fyދ�K�g�{cC�>����5M��֧�5�^�ּ^��ݼ�1C-�����x5�T�h� S��1<y�1���W�o*�QL�r��}V��h��}�Q�T㣅�c,���΄��P�3�*�����}��eq��wR�V�rue��=�؁݁,�}¡�4��'T�v���WlI�S���ȓ��Bgi����yś�AU��&%�S��oHf�p���o�f[�6S�cYѣ9�+Z�<�Cc�C���z̲�oV�T�!�zq��Na[�,DU���z>|� M�Ȱ�-���zT�Fi�4�mvZ�ߧ����*v�"��/��*蠼Bj�uv�{j�Eh��م=�3Hnk^:�#�䍗i�H�������Yv�`��S������մ��)x���򷯧;=5LY3����y7&�ګ��8�ִ�5-�<�8S�w����y����N���?��Ǐ�� ��ǈ����u6�����ˣݽB�"�cO�U�������[a�2m�Ê�g��l�{��@�L��D�f�x�Nב����Y�P�@���@��Z�`%���e軇�W�i�if��C ����yԔ�z��Z�s�P�5-n�_Y
݀�]�Fl��7L"���;�:������ζ�����%x6�հ۹�<��mC>0�H��F��x�"�����Eu)�����B�il1y��Q�՗��B�,X������P�~m2"�=(�7�s�F���;~���4�o��j�Oi.�Y��`<n���b�P��W����7 q�AŃ���i�ny�bt4a�8��o++/�i0{9��ݚ��c�$;9��粣��<�;00�OE����l3��ᷠ4tD{��>���m%c*�˙���OgZ���|�C�p���W'�R7�Hm=3y�;��� 19�؟I+�>Fߧ9��3k=U�گ-i,�Fƪ� �c6�=��9�$≅�<@��Pw�����|���"�4�/wʲg+���цQ���֗���mR�<�����_�]@���1��fM���mR2���i6�?��ک0b�o4>���h$���;o9Ú�ў�f3.�N�x��qD@ztz�·�r��� ;��$#[��1E��;o�e�̗a!�@B�*�{yN��6)P���;����
�����w#�O1��C��KkOV��w���w��{�?o�?�z_����x!�?����xV����j�[3cY���v���qb%��\��6n��U�q�e�do�|�P<��8�t8e�?39�s�7^Y!��w�3��R`$�۪i�f �z������������?I�B)l0ý�S�6Ձ������ ="�l��>�C�s��L��S��Ԩ��ɨ���w�X��y�Y�
����G�!]�_��
.Yڋ����>�@W�`�{�����w���HfȫѹxLb�=@L�-�"�WG�2V�^(�ȥsw��*65�׼��V;�0�m6-ǒ�6�;�70I�QV�-�5����kN��2"�'����Q��j��[�01�Ga�P������ާ6�n�C�DE���fĹ��o x�7�7[�3�k	מ�>�a��6"Ao��n��b�5Yw[yۻ��Z�0�Cѭ��_[����Q,�����)����q������@��4L��&�w�U=ݍ�u�;���^Ξ:�o�,@,��9�Oxؘtw�$D�Y@��M���0�4�{t��3[�X�&א9>�X��O���P2u�9��0m�`7��ǽ��y�orыv2��p���sN�GWQᾆ�l�{�-�:W�[ ���3+�w�{���$17������Mb�S<�W��������_�R=\U:�5Q�V�5D�W>7Km9�����]�'NzjEү:��/:�w���Y/'L�{�s�ٓ�����q�ǂ*������w��׈x�0~~ؓ=�J m�QŪCR>�;�w>�5 47q ��a��zcЪ�R�|D%v�2P�vy"\&���4�60�C#�zy��݌xt��7����'���/<��hb�f!���V� �Z�Y؂���ex�"�۵��P$���&��y�' c�l
8i�c9���#�<�����4�e��h��ڽR����r�v=�� ����B�� C��lH�.�1fu��;ހN ��s&��='�=���aOhzd0���U�i��+�#�C%��|j����������b�i�T�1lM�y�]��b3Z:���5�1t��ruA"�)/�ժ��H֖;�QT�����_L�W�G^�?KY��GE6�B��Ͷ��<L���<�\�y�t"y��\I���c� Zzwx��\��q�ynP,�[����!�9ڻ׺"�N���(�7������M�D	n��>�x(�{ږU�qfV8���0:����8V�+(��ϛ��]����Ѥ�푲�	�*S�_܁Ӭ�m>�yL��Л:�	8��0��Ct���ssʼ[0���λ �������Ϫ(ِ���[��k;㺞5���JƱ��6�y��L��YE"H��b��,@mȀ�fKhWJ��AC���(�D�e$�]���M�m�KY��ą�j�uCWßO���{{4{���E�+��%�"#
b&�Z���q4�(�s�gD;'w�{]�=�^��	�)��������#�.7ݤ1���ݽ����q/ȟ-��^y�k�y�Ἇ/9��/�����^ +���{����θZ�]<g%[��Ί#��]p���������9�s�~�K��4��Ħ.H�&�Ҹ���ɺ���y���A�����|�p����!T� GkύmMf�3Du�Z�!�4{���u��P�܋�;ٝ�Y������B<��2�
j�ml7��)x��fp��0א:a�u���M�<�T*Ocg�i�j���Uj��m�V�qt��8���ue�܌{fc��Py��ܪ��j�G�Yσ�FFk9}n��	i�>t	��<F_>�M�^G����W��[��{�S�̔�]��1�Y����-+�w�\���G�36��[Jh�'�ٲ�\�*�)L��Qă9Q�ș6��Y��{n$6��$6k1���x�+��߼F4]�{�͐70CK�3\G7H�3X�I�g�6��^6KT��xH��Ѹ���!����cV���.ܷNGs<��^��AfE�����z[����i��<̻��`̪�3��]4�C6t�q���(�>=wf���9C�tj��r��!;4��\��5.k��}��S"i�١�Ę]Ai��s��������wZ�v���R���f��Ɏ��2�g���4m�]?�;í��K�A��|3E���4�^��W�:����a�z�}OE+���<,;#h�s�P�y+HW3e��]�c���N��$��^o;�����������ׯ�������< �׉�T�o0���o��,�i��ԝ�zm��+����קg�g3|U^���yWs-������{f���(�y.*�%��h�4���SH�tCMs��>PK$M�A�i*�j�h0x{���(Z�gc}0�E�Yid��փ)�4��:4f���f�e��S*��\�h{��[�J�d��v©fKV�q��/F��	���x����jm�T�Yo��;��w��;.��ޡj�cR����=R�!��I���q{="|�Ƭ�#�x[!�'&�V�w��CĆ��+�4�!sW��J�c�O�>�7�#(GE���.��F�Fk�y��v�!�qv哇�k�i$k�gbB��Y�g:�!a�q]�9���s[�t�9^[vyB�>�-�)�h�%'9u��W����^2gqP\���sZ���K�@���a#z���G��Hn�ljP��	�}��·�̛:ŐfK�{)ٱ�;�M���G�=jf�j�T�0��Ld�T�B��f��j�8�\�=Tь-_F���w �=Ν��C8����'�9������@{�?~���U�aʊ�(j�A����FNY�elT"c�ټ����]�f_��"K-ӫ����u����7��׽�o���巁}j�+����b}&s��Φ+!��Hk����k�#kk+s͟�m�&Ω�s/:t֩v�8<<]��x����T�^wIK���!N�����	Hz�"�g�[ʷ1���i���ψ���Uh�)�Z��)Qѝ/�먦6��)��Z�hx�0S�E�������	��7=1zC�ۡ�	�iv1�}�Y#h�iU��*�E7=M�����i�rq���E@��1��qF��N���L�aSǚ��h�r������t��u�q���;��������L��Bq1�0 ����dY����	��k�}Lh��(�u��b��k[4�ˆ,��{b�=���f�%��>��%�rq1/Wm�m>; 1�[q�k\����m5q���Vw;��z�0��)�2ه"���c�L�p0uȷ��G�y=�L�`��bn�I�������a��*�6o��C��F�ÞX%��ߝ��1?0����q���L�E�󗾾�Ϊ׻C�[�PN���݃�"�ૠ���JWt*���>� ~�ɻ.����m}_��z[Y�Д�m7oV��9�*�w�@���"3���IL��׫OG��-�&.��M���Bb��#ʲn�d=��!�S��0�i������s"+�L#�b J��ҋ9�8*]n'.�T[<>E�l�[�t��S�����ӡs-��s��c��q�XXT�h�kVk���!��ER��ˮek3��돰�*#8:��/�(��.��"Q��r�����e�|I.ѝ�{g�lU���ǘ����v�� W���<=������k�k��J�^3���Q�hȅ��v`xC��K�\V��P��o>�Ks�l%]��a<��*o��C�PY���{XF���fMg#\�a�L��l��z���d�a�"qB&��{�ˣ5����%�!�:�b�n�G6�8��o<�/�Ci�C�g��0醯F����s���B@�ƍ��}����;�(wl9����s�Վɂ�+}�	���0e� :}�L:��48g���N�z
0{&��tkG>B��Z�\e��xm��'���0r"�u:-5U#��7��L �ڷ��:͍����\����?X~��ҹ��:޶��f��/������`�tP�i�1�v���� '�>k6{ڑr5�0�5������˴�d�>�%WۮY�t��.w�^h"|�!˫w-^���Si�C��[}s�͸��k�k���+n�p�Cό0��(B�a#���M����h3D�����3���E�1��&��y���n*�ȵ(y��NC��mxoA"�%M��Nɶ�����^�E�^��Pi�p��(�n7Q_��Ȁ�n�[ë�a�!�_�v��Տ]c�	����z-����]`�u	�5��L�tK��Ҩ}�`DQ^�18<��af�k%,�$R 4����~���or�2f<�T��[�R}���{��|9k�q���7�`����`��E�d:�PD���s�W���6��c\<�����^(��������ҭ��;�U][<����$Vs?�]j��i��D�JO�b�b#S�fo����ǔ?��B�tk��ȗ��8%y���T��<[�.uL�C2(��a�l/`%�'hr�>Y�3�=\ڣ�_6[�k�C|ϰM^3f���J�:έ�5�Z�i���|�IΦљ6O��xWkb���b�[Y��b�݊�/���E-)��6��S�i���5�Bƌ	R�1��F�x|��Vp�k��x��' N�gz���v?�j!�|�z��ɧ�^�;}��6�5���TV_&h�7����u�]͛�@�kB��>6�0��q[%��'Z�x%D�f˘�wV�������S�q+�@��Z�p�i�5�w�vH�`q�[��4�"����J���ۥ�b��S(l)M���)8�9��Ӳ袒���tW����܌{f��;>rn���" �ݵh�-7v�v���A:�C[n����e-��g@������m4��#���q����}��z��^�9o!��7@w�F�0.m2!�G�E[Rh{���<�]��$Y��������T�o_߷K������o�O��Y���kWo+x��iܝl�Z+)ܰ�'�Y�(���*�I�T4�W8*����eh����m��88�6��T�9�_Q �.��v���;����ݷ�/$n>�2m�G)����W��~�}� ?����� {j���!�"5����ע駘���n<[9��kP!�*m�.��D�ι�׉��uj&e���j�f�^��M>�}>#�+�O=}i���Ζpq�2p����T��]Ul�+k��kݦ��4��ە�����\H<MP����m.͝��@�}���dB~pZ�=�y�x�~����C�NϚ��X#��f�}%)�kR��3��ͩ�v��~�����]�G��������Rf��l��XM��w]�th�Hbݛz���J흙�Q�q��&�;�W��V1O��PzR7�����01P���5[p)�󢚧\�Z����s�*F��f��\��#rᝣe��x��[Sz^�~MW6�#GTBl݁vX�D�ifM=�9�Z�\�j�6�\�Q\������|^��_�F�6�a	������i놷������D�p��?�(���RO嚭P�jUQ:��@��a&�8�Qd��7g^f����)�U���tn�	�@g}M=�%crO>#6�e}軗�`e��5�����ܡ�[pw_B�[��,1�ԭ-�To%kÜ���A�5�N���_�[,��arknS��M�N��=�6�ٍq�W1�R���k���EXxN�r�p�e������U��y(i[�f�f�����v�C�Q������9�-\U1��`��Ք;��5�Q�i�m%Ӆ��+�[�5��V�9r����Av��l��N���T*MV���ۺ��'�
�+z�Z%:ޭ�K�Պ��<I�w���	�b�h|]ګ�4Z�S�eqo�7{��*ɩ
y�D1!�\�����;�K�U"�O:��W�Ք��xb�2,�3M5/��\^��Ȓ4�h�l8/e<�=���ᲯG���(}��5�yn@�ݽ�`�LPm���=OK��8�_}tpxqH�}Rwu���ޘ�,u9W���X�6�8<�<�˔M��V�;��I�޾r:�8i\�
�b�����<Қ�@	�iK������9 I�b�Ɇ7C�ᾔْ�,�b�O#���3Eh�*ٜH%�R��H�9
_"l�f4w�U]b�i^�^�B�Kq�K�촦^Z�`��Q�;˦�2��s�E��53�����!6�n�M����v���"���7WͩW�{uҦ�^�7{d�a�.dʍW
��s;�Ȝ>Ŏ�ۦ�pf�ɼN�l�*��ô��=�OI]Yj�e���1��b��4��(/��+g:���O�>�臋+z�I�_&��^ge����C����=Y��L۵�t�;;U�P'5��n��T���5le_Y�t�X�ʺ$�5YN�k��E���[�+`*Fn+f���Z9_fD��\f����V�x�D������ٔO����qR�:Y���e]t�֗�ˎ��g<mma��2)2�۳���V�]@>B*���tp2������Y�J�]N��`�ins^i躹J����Ϸ$�;�)���c�"��Rn�k:��|�Vl�z��y9�v;�ڟvM��ep����2��AT2��"v��������q��S���5a�[��2�X�!Cr��>[�>���iU�Q�|v�Vqʓ��<C�����&P�j^���m���;;��f�J�v�aAK���*����nL���Skr�lRcJʥ]�;6>ݥc:�Za�d�w�W��"�2M�����x�msU���\�t�c�{a��{AH���G�e9L�Q; �Aj�<�yfr��oE:,����*�ޞ�y]�p��ͪ��`���5��SA��*�1��
� ,r�!���K_G5�"���X���������S�e���2���ˍ�\��O�����ߝ?�i�o4|�V^��LJԟW_0w��*�n>�3vg����o�>~y�<�����D�Q���9�PP'#~���̮�<��<x���_���ׯ\�����������~��	�Z�}����~�Q͏1��"����.'����s9���ׯ^�~=z��ǯ__��������zv>˯�CUː\3���@�$<�l��r�	<����t�=�KI�Bm�g�4IM�P�Ǟ��{-�^ϑ�9�|�<�ZĴ��v�G �N����\�M�y:���#��Ϟc����Ɠ�ZM-.l�W6'�܊䦓O�G y��rJy���O*(6�RrGZ(�)��A���l�9���s'��O�y)�a�1���m�I��̧$)NLE4�E�6(9/ �O'��-��bh��6�Ӣ� (��$��VL��ڲ�m����$9����(jR��p����R����'�i���n��J� �*��8C��o���9��?C�?�׊<x(	5�Z&��{�O�e����M�E��Nt"0����F�}$섡c����g�N�ރ4]���j�����f,�i��ɇsZ@���K�@�ޮv:Ti�Ɲ�ڵM��X��e�mn�rr�A?���|�{�����|�m\zs��߸��q&�o\����ޞ����u�U������)56�^���8�F���>��0?�i�'�i�|M"
�u�a�n4G3�f2wUM�n@,_�R|���T3�CSpV� ����H� ��<.4s�p0:"�e���>r���D��Lfu��A�ن̅�(o=��P=~hf>��L*����g\���1�h�aeA鞕dd޽�Ol���ǚ݈4�{;U�U�����ܩ�ȝ�'��D�_SƼ;n������ɋ[s7�z��5��<+ud�1lVU%���	w����(4M�h0_bco��PAC�(�����D��Z�M���S����x��*�#1���׮E��WVf�3�;���G�E;����1����6�ux�C\#�P}�!���}xA��q��T&�vv��u�T4�qv��r˚�
n.�A^T�H�� �R���hX`�[��b��\L���0zj%�����U�_Xw�vs85��̈>}C3w��z���]X������'��*�x��?���w���=��~�#n�sB�m8�#֪ی3Q��F�6��[9@�mE��m�J�7��C`���_�"L�(<���V�ϲ|��K*��1+X����5|m�D978�3N�lX$6�e���Z��$�d*���;��Jd�kMҨ�8O({��E�f�m�՚۝5cJl�$fÉ^w|��ǳ�ݬ��:u��)L#��I�ƥpvF�I�'�nڝ����7�I�-E��P�@��ɧ�놡�}+�xڊ�M"�;�����U��}����kQW����.�1��S�g�G��6�8�L�ңO�-jǝ�.��d�Tf�j�t�J�O�a�mɨ�ӌ��� ��2$��K���x����x��e��l79�}RQ=Z�?z�>�7c��2p�Vf��'7YƂ�e�&7D��<?BsUj_���e�4["���x8;w_Ҏ��m+�1��07�C�����w�ʞ�)^���e�Sd�a�O��%�|�e6d8��c�jl�oG��Վxt��C���ؗ���MT�i{�����Ɔe����qC�E�nt��6��Z6��zgi�=¸��b�C���5��
ye�-{i�0(U�38P�����m��ʯ2s�ڳC�_��۵�w{	9�{8���]�=�Sɜ���`N����r��u(��Y?���y���xHQ�hs���:�p����(����x�q��<<��m�]w��*�0�5(�q�����o㯤@���`'��<���D⑲�p������8^3�C�~��GZ���B��(�'z��f7��@6�p�\�_M`�=�1�ˏmn b�1ǥ�n�6�s]�{um���7�q���Q�+k���ў'����s⃧k�Od���MENo81̣���0�iF
u��x�>ed��@�vA'ǌ{�瑪��H����8�cM����6�'�;�VvC?,e�����#��ǢS��+��!'�lT�Eޮ��Cմ�=����Z�u���4�\lz��n�
���5� x����s'),�.�$�����[�v��4����޼3Q�9P [��,*�Q[�V�u�{Y�"��l���u�J7���t�*�K]���D�<��ni4[����ܧ�-6�O�ę�3��(41�v�E��evl@�1�&�[ ����_(�qda�j��i�����c��Se��:��6˝��*8l2�=��goY��B�k�y�;�\��~�M��:��FP���g�A�;�^94@�k -��!��MM.lȈr1���|�J#���]Ձ\��P�����[K�.�)yVZ���C�Ɂ�)�Vxk>�a��a���@
��Ћ�g9��f���S��g"(Xz���ĕ��)է����)���]��Y�f���7��m�������<���y�{����`Ot1�K`fín�?�נ��s�\�"ُ��Ȣnd*Q�.Kַm5���d-g��}=�l��4�A�;���[P�4�G����/&�T��ެ�2ʠ��n�S5�؛��^lD�Ɔ�`�˚尽_@��S��*�4�i��>�D��'�ʧ��*i���i-��8wz&� �6kX����1���FC���2u�+���)����Nv�r�haC��R��^�zv�"��`p�NO�O3�*;*m��JKh�w�8��Vu���|t�ڳ��_�(�j�6�PDO0��B��|#��g�1jjƧ�u�2K�Y�$�|�9v���,X�H`C�T�^�%�+�Fb�;V���;�U�����6�E�N�3gguM]OSt�]�=9W�]U�;��<=��1�O�����S�,$m��":�:C�)L�j�v]h�1�5m-fzb��.w�y༃�P���?�)YK*mb��x�΁�� �gE��ͪ)�ot;��_��)�/m����h����D�ҧ�����rt�oCَ��e}7-2�|��+|��ƝB�@ٮ����U�� ��_�ak�D�]s�[��\˥:X��`�}��1Xk��������`���x����vmg;�-�'����`�S�Uξۡ�J
"�$8E�&5u屖��)@iε�2]�p?/��~~������y�s�9���^9��@�Ǐ=�x�X�seq���tab��ݲ�r��=���Z�O����Hw�.��i��S[��{��-;{����fڹ<��R̖"*݊��}C%�|�9�,9�27��Ԭ�9�z�(&'VŖM��3bl�LV����;T���V]ȞWfz��4�6�����|"s���D�����ɸ�p}~-N�~��mM��y+=��?�eu�ʎ��v��֜�Ǉ��wrs���N!�I�� ͭ����cj�1�y�C�zƝ~��.fzo�y���`���\��mL�y����#8���j�~�?xӃ�T���z뷀�#�L�s6�n(��K:G�Ӷ�t"!j��{�V�Q5`6<ZO��K��룟L�~��?S����뚑�o��N���d�2�;�<�1K��Q�u�6���	�O��y/���ӊ��5
Qj�o�kB�L���IP�5�)�+q/7���q �c8��m�����9C�95h����*!��>���鷮�9���{y�Ԏ����:foP�;7���Kߐ=���gt����3�m�o�3��W�8c^����F���J��-ׁu�2�X��ӡ��h�"Ot��*S��:�}�g_��SqI˒����G�u]7�I}|�W#N79��7F�i�i��ee�
�W���A3��^#Ǐ��=���ߟ=������0 =���!���q���?D�1��c� �
�Ӛ≁���M4M��"��C�/��j��r��!�����x������MC�U��1��mtm���^-��*�,�j9耄�}A~���>�;m�]a`�� �~��⿱Y�P��ï��L�`�Z�݇���ryb��G�Tz`�.��Y��(�jmM�i��6mK=�ȹ��ݔϚCz ��ֈF7�#x�H�jņZ�whON�9�-E��^r]mו�{�S�I��;e
.�8���<��h^(<����>�	]ЪYr��I���2�:)�))�Ql�f�F�5Jq��,��5���f�"��S%kP��y8��c6�]��vi��[z�%��8C9�i�ÈE�C+ןA�[��i���2"���9�zz�%�e3N|*��r[������E�Y�s
1 ע��(b!�:;4㋊݀�3�k	�{�2�o��k�s q��e�O�e(X��hL��k��,��O��c�ƚK�Vu՞�z���ά�B���LC�Tʸ�p��]����^v4�=�?X�E|�=<{��rwZ� +rwn��<���l���B��:��Px/@]���4wq�G^���1�Y�gS}J�_wg-3���Ƀd�C
���+��,C|�;���4z�:����A���At(�OÇ��Bx���x���Q�=�~~�������~�܌\}���rS��̜�YaJ�jgLlfw� Xû���^ا�4ӭ��Pz׵y	�*)Gxɑ�;0f��2y	>�X��S��>�21�7���}ۭ|�E��N���f�2M��5��s���$�b�~l�x,�+�1��	#���M��P�湙��;�V�t.���ds� ɕ�@��embH�>����@�-������z����3�&�e�eWL�v��؅�Tl<	ƶblki�k\�D��6�z�#[`Yïy�X�i�I��W��@�e�݁r�+�yށr#��KW���)�uqm�`�<�s��[̩�o2�A�UV俎/r7�9EsiwM`kC6fs`ֳ��ɼ��t9��|՝}]��UziQ�@t"4�ۯ; K��@�k�$��FF��L�X�E��[U5l�p�[=�M⚭�ω.���1�%������Mx��ybĎ��G�x5>ιb jzw}�F� ��.�s������A��L��i�bi���5�/�f�$��TA�ô[�v��D�zSd�[9���_����I3C�k&�\�O�^_����v.���Yv�B6hˣ7*�x�׏�� ���2�����<T�;\�����9mu�,��#��Fpb�<5�|��MHxQ�uos�V�1sw��?x�{�?����k+3��	�wB���fsX��h*q^f�a2�"�ϵ�[Mf��W4+���w�4�m�lu�ZJ��\���o�l1�k���o4�4d�Aq)쉍�z���0����^�mk2|`�׍���`��R+)E��������-D8�#^���5��mc}Y1��UM������ܠ�W%s��{�|�SfX	H�
��eGT��vS��Igl�xOCrfN��s?e�/���g9^i�N�c5�(7�����-{|�ˮ��8,�}n���&�	�I,��K����Fz����[�D����m��tQ���ڛ���AN�����4����W����$���׶$/=�QՂ���e2��8e��*�eE���]h���9g���|ŋO5�҅�a��j-��Y�=nI�I�qr2y�q�4��n���x�\�^��;r̲�b��"�̛_|b�c��_�y�8I&�Y󙌆�� @e-�z�39zg�}�M�����L�} �z����EϺ"�����>����c�~��_�T�C���k���^����K61v�徻t
�~G	~�]]QZО
�~���u���ڽ��l��Q%��;{�k�/7D�~y����r�1�1<s߷w��ͪ�
�n�:��w&:ùlr��},9�kW]|I�Z���Ν�PN�z���lN��In�V}��g��U^?���sW��<һ�굾���^cM~f���<��pkW3g��P<���a���iֆl�djJ����֭�B�k�`A��q�g���|�.M�f�[����|�L�P7~�ꋈYzDg:��[�M&f�o�����
��MB����@��c��~0���Ư��`
x���VC�-٣�˻��C��rq�Ĉm��i!�uM~��Lč2y��5N-�xw�@�wXC%o�$j�x�ȃ��p�Ѳ�rj4s7���f~L�K�d��fSx�D�-s?3��ҵ�/��e�����7���\�x�WH/Gϲ�z"���Sq�e��wGn�U�t�'b��ƀ�P oE�9~K�ʽ�D�@�Y#U=Cg����}4���1���Mc�w"���J����k�>���##Swk�e�����2+�ݥmp����j�-w��5i�c�ӓeΘ���Kp*�E���4gB#��L1�mn�Xۼkw����h]v�{fm��4�������eSL���G�N�~ƫ}X_�����?�wW�m���}X^Nh����8��y�S�/2��ŉ�%$��Cz��ǘ�W	�Lρ��L�NY�5�J�&��=elB�e%.�v�Q�k2�=�'\��&�����ٗ2!0���)���йB�Ty�q��<￿=�����)Ǐ
;��Ͽ����k-{�Nx��q]mѤG�=25��8�uٟ����@���[�[xң��j�xBfut��jM�'�at�q��a�bsa�`pi�d���[m{dz�쥷z0m���ΜeC�q�{3��������i����_����O1r�7�ƪߚ��V�ӥ����#��@�,�\��|P�֐���O���Hލ/m�+�� ;H�Jr[L�6����h��2��)8�?=�H�)����(��¯�l�+Kn��Ej��m#�e�9�31���x'�.�ɜ�4[��Ψ����rj&�eS�qwq��Vޙ���]N��3���8/.� �ފ.�}���C˴�o�1X�7����)�[�7��aG^)r��礠M�Y�e��okb��j�r1ٍv3��,��F@�}M`Բ=��oYT���2�ɦ�-�h7���$"��mX���Z�"b�3Q��F����G7���55͵wo�����SJ@<���)D���z0/i�bJ�E�bS�&��n���栾������o�v�5r���Yo3+q�C�������dWՁ�Ż�h)��J�OE-����d�̹y�7ݏ��o�1Kn��lGw���-_F��ųx%NC;�x���¢s��^�e�Ř"�u�x�s���������on��Z���ҸXK��܁t�r��f�_WA�qB5��K`Rc�XE�,N���<ܺqP����K�[�E�Af�nS��:�Ў���������ⓀN�r�j�V�p:R(������<渵�W�X�B�1��`�:=W�'�f6!�}m����a:��ʡ��e��_F�v��*Q���K����.'��Q^iƪ[��fug�[+�yR3W���I���t�ul��1f�X0�`U�n�bc���fi��b�BG��U����{�p�AiE8b�� 	$�*��Ks���&D Y�}Ǎ���N��,�����MT�{��j������3�V���9��=�8��S2�<��l$�����
��t��h��I���u=x$����Έ⻚�d'�ru6>��m)�{���֚l����J[��dYIS:���+ǋs�l���l���w�J7G�޽��OT��ܟ$d���*wV�e���o(k�(����l���2�r\,���XoV^�Ҁtxv�Ƭ\�]��Q�e��Pl�I֟sa�̝Ȩ�����~��b����v���U�k�M\B[Tb�:�x����S��Vf�X�4S4�m�Yo9�E�Y�ˀ�iБ�C]��r9��S�`��9�Ƿ�Ѵ_KGT�	�8Y.���n�ѽa(��N6�j�u9ۮ�=p�B8��D��Ή/I�U��QçJ��a��y}�M�%?![���j��L5�ٛ۬@�N��%�S�z�ٹY���$t4��).G�]V���gU�ma�['-wH�nҹ�Z��ZZJ����3,NfX�K]�U)��r��z�7|��w��Ï�Mu�b.�&c��P�лҶvh�|�ޛ�WN�LK��VMY��H�2,:�1w��h���5;���_0h�c[���[[�h�!������z�PT�Mo�Vs1s5�B�q��j0��:S����jΰ��S��㲚��9��]�w��j�+*�4�ι}��	��t�G$\m35���n9���Sf/��Z��hi֜�sw7���!�s�2�֘�>�Y7;c�M`12Vs�s��ڹ[�H��>���|�b]�O =�x1���*N ��t�PK`�퓜��izm�˫�k\��
�=�U����L��YVk.�LC��9?�{V�ut�f�7O��.e/`�.	��b1o4%�kr�"��wLڨ��QcS�O:�hS�Y�NI^R�|d�{�Z8x=�bF�n>p�T]]g-`�i��=�{���=�!M�?Q��o�A�BA m#�4/ `��T��!�RD �l�ӌJ!S�s\���	�<�xm�#{�C���/��X�����F���6�)��ѭ:=�n^3�_����ׯ^�x�����~>��_�קj>�4Q�N���Ɔ��!�MB�~���\Ĳra1�x�}|}z���ׯ^�z������~>�_����}Z�[?�~@h�GI�46���r4:��<��Bh��*�<�$9��"Z(��| (6���������'^ZWmI��ȶ�!�l��������h�֚E����C�8/2R��NO*���R�ml�t�/6���AI�-�4#��Ns�y%<���r��4�M[m�.�%�S���ql�h.�R4�k&���ժZ�#y��.h�i�4�'�r��4?6^F�퐭i����r�����D:
�  m�Ѫ�)f�Ym����p�ʶ_J�A��(���{ip:kE��g�Ӌٯz�6������K��83��O;�n���"	(׍"@�9�G8p������<x��~~}��>�!NJ{p>?�x���LR=���Wk����C��"�(���4��ib����:y��י�u�%�E㟪�����"���Az��)7kh�f~dEr��;KC;`P.����CQ͇�5�oM�賒3�p�0�`e��~N�K�tri�5��!smB�.�747�óws���-�)�׻�N�um�a8b��q;>,�����8�5�.��yT���O�m�����Μ>�V�����51Kϧ��ؚ���vfp+3�9�pa�]F�EA�]��m�:r��r����2��G���2}	?�{t������	���:یHLZc&����6txG�?sL4&�-<2��&FZ�r��ie!\���tb�+�oS
���4���~1x�1�8v�.4s���A�i�i0�ς1���������i��.��hU����OwOM3L��-�T!S�r���c16�L�Ȇ�}�&�l���`(���{ƎV��j��f�f���ol�tEsH�z��wc�v�Co8d 1*}>>.B��!���*�w�U�̪fg�9�*�2�9�Ȕ2��9�!ryO�zK�Us����+,S`��l�:�gٗ8�h��DE�����:	N�R�2�t���d҄zm��ylpI��1��O�M+oqwW2uq���^�x��o_��y��{#;�2�~w��ݵ�0k7����|k���H��m0���ū��f"�:SA��
'gg0�G�O�~����l&���Ǽ�!Uv��D���z"�).Tæѭ>f�#;k�8��~='s�?��+l�Zs��/$n����<ѫ�Q:���X��C�⤦�	aT�ش�Rww�އ|�c%6l	��jD8��R�����<��@�`�^o:�3_��<�{gή��ʛ����Ւ&w fs k/\��k��U �v��Yt���(t��l�L�YZ��Z�z��<�i��Z��f5�b���d���i4h?(cGA�Z�ʹX����X��i��Y٠��t��C7c�����\��R+$R�#�W=����|�y�j`�]��qQA:�Mm���Ŏ�b"�ϰy��]f�Ʈs�	����[eŮ�`f8�1��VN�j��ٸ������xd�G���j��[�G�ذ���]r;D�ye���;ġ,��H��LH��3�g(�S���Rq+_a���R����a�|���m��~#�'7���q/htl�5�u��p^���+�h�w$��䒛\��+��Zp��\>�{f���!$��5�;���#��������9���snm;��Z�1��i�S�;�s]
͵4e<۱�D����,���{}���^����T������7���z^
��m�=��d6����a�>v�-��Α[��Ǎ��g)��0��y�f��M� �#�#�i=��E���l�{%�8 �m42\2�x[Jc΄��n��U�.z�\+�� �p>C�o�S�G�YW��t��oE�sl���`�3kP�m�z������Ig��Xҵ��^*^<h7F=����t���W�b����pD���L���D<�nT]�"%��Z%���sl��?�T������8�_���;�t�~'y��K��v`���}���hGm����6;���Z��c�)7����vpW-6d�0��@�M5|5�ck�Rȗk}��������X��aF}QP2EtQ�n=l�p2<y������q�C�����I�W�#]Wє~�>�>���%s�Q��",H��C`�o��Z����[��iΎJU"n�N&@�p��6]�@-D
����^����-ݏ�U�j��fZ�8�x�cY�d{ZkSe둉=S	���O���{>!���W�b欇��~\��O��q��N�h~_c[�6�,Xy}�2Đ�d��4"K(�&�o�~��
ʿ��X�5�`ay��]]ғ��#P�1=�X�o|(5|z���zM<������sO�&���Ӹ:���s�u��!�/�����y��;�M�=���(� �찰�dL��y�������%[���u�z�2�U~�����ҧ5��k�"-[0�[��oF{��7N8�^��/i��Sgs�Xړ�9��6Y���m�V�N�SV/L8��d!�=�:�q���D	�X��{Z �E�z@̈́D�1Ŵ�y��z�.I]��kD�������M�
0d�\�5�30�$�A'���R�֛h�R��8uT��qq{�����/�c\��7Xn�"=:q�$���X�Ύ�,�wfZ1�����e��W�Wt��P����&�lƢ����N�&�$<[O�4h��Z���4�Q�L�Y�����yLl�������9���wH���,�5Kso�(p���vf����C	�p���v�["�JM0�Nc�acw�׹�����`E���Pˤ^o�?<�0Ny�	K��u�
qnF>sh�)��~�A_��w �j\�^�c�Ox��0/r3{S��Ml�ir�3�������@wO|���~M6��?���oz-�"���?U��o�_-�j�9uk��3�]i�ˑ�X�s�W�-C4�4��R��b�/�_a�ԟ�&��8�N����Y�l,�&�yuĔU�
��˅u�l���e��{�p�l-��e�;˳6�mݮg���R^�����~9�y��ܹ�y���y�g�x��s��?hV��}x������uLƣ�'ӓ�BO$�E�Nö439�M�Pv\��ji�������{%^O4V���m�-d7���� T�N���Ʌz�H�f*Y��-�K�cN���J�1�>n2A�v2��5!��M���D�!���v�+�X�V�=j�ݴ�5����y
q����l|!'
�z%��0,�θ�)��`'QF}y�y��ૠ���HJ��{���sO�8"n�&�!�[��S�L�
�P������5�
��o��������3=�J�2UflMF\-4���"{^��M[�K�'����"���AR��V(�h�13c�yEM�C��,;���K&0�oD��貧��8rX
�f<Z��(�8&8:;5�d˜�<��X˵Z�r�����y�5�É(X�hBp��\N�g�32l5{�Cs�B�0��A�Y��1eC�S[��O�v�|�S��2}+)�#�1����>����V~� ����U!���W��~h���V�wt{a��ҁRم�`�&Ýo��À��g�^oKI�z��&0�K@}K�{�LZ�������5����.��m46��hD
DF�=5��Y46UF	��u��S<%���l%�v��
%Y�����Ū�]��jho2s���MÅ����7��������oOK�����9��w�������+��5��w3��Ga�ᇽ�9����c鴮=�QV�ο���Z ]�M�Y5������.�b�fg���<^O:��m7�6���Վ�o����U�j�z-��6��k^��۰�ZZ�b}ͨ.�wk,m�O�1��,4T_5�)
K:����ͩe%V�q�>mz�7����~w�\��Ƹ��5�)��������R�՛���oB�����!7u�θ5�5{���'���O�]�ŴG�_@d�=t�w��է���Pxz=��G=T�_/T�f�@�oA9�f|9,i>U�5Z���F�:�ۭWƁ��h/~c����U�S>r)# w<z���]�iI��d�G�T욂$���F��<.���ʯǱ��ĤXU0�5� o4�8uj(ݷ���mĕ��=���ֻ/aI�Hۙ9AvH��L�t�i�j4:�W��XL�����+P���<���D��}�2�u5�q�d/�SeZ�''��ƸOe�5\1[��b9�с����+�����Bɨ��	W�d1Ziѻ'e)�Ǒ��]Ī׽���Z�n��P�Uu�3f8�ӿz(Si���4\� θ�ϊ��Y^�����-���	����5q��WX��er�h��mGm�nwn5������d�:������ۛ(�� �o7���cb=P��s�dh	�X0� �e*�Sq�@Z�YJ(�a�Wm"x���5@��c�"�p{��59nץ�n��y�)�E?��	�O����~�s�l�JF�
���+��L�̭Ks6��_<0�N��i<���4+����~���
R�eϧ8CD���@�w�����9��a�܉fa��Ɇ�B��{E��h��ell4��qF^��ggt�ۉ�X7N[���X�$��. d�o�߰3�F�9Ax�X(�m��ՙ�,j�\>Y�[��Ы����աX̰�Z��y�]�� =�Qo`&�.��E�1��y��0�x�'��L��l��V��w^�L2{�8�&�`IU�*;�3�������1I$�;��D���;���$�ْrr�6�7��(?�@U��f)�2�+z}�=Ϥ\��+�H�=}i��W
M-.6�T'�SuY�ol�c�.��3��ߩɤ�m��ft��>&a|�����r>g��Y��D�:�w��AC�<���U/qtw]&�;"����.�������^����{�\��������e
ŋ*�ԥe���cV�0�o��i����eCR�����@�׃<1-R��U��c�{�X
�ɔq�8�4m%������=��-FJ�0[]�]�y�h{�yK��Ԯ�pVF��<2ͮ���aw:��ӵG�ͼ��>�y////Uz���I�2 )'�ʐV<;m���x�v�A{h1���(R��IeM��,��ܞ�-�6_jGZnr�|�|�%� ԭ�vgߝ�O�8~�K����)+��O3г�v����;������XS33"|����i�|CM'G$%R&�E� �p�۾�s�ѫ-i��������cW�1M\�T8�)fthȼt{Z��SeW#9=S	�d��Wqn�S�D��o\�����}4�Ib�0C��q*,�}�͈I���yoZ�f�)]��R�~�-=����P�y�A�r����Q�]�޷L	�O��2SH�y+[rn����&��D�Nf҈l�^��W�y⡭��d43Q��c9�V6�df���5�Έ~%��T=[h�Uy����Ӽ���S���愡c	���iƀ��X�6}B#��_��{�;��S�;�g�7�5<!���� oR�!w?���7-�<�4m�c2��C5��C�0h�t7
|gy�Y����Sr��qT��P;���zݓ@\��-s�
̽���v~�;���y�c�D�]�`FoyAn+�nV{O�vb9M�Q�����+Fa�����q��6��z�=[R��1�Cݛ�2N������ǿ�;���Um��W��|��Ws��tp���쭿[GĀOWr��
M�m����sK}��wI�K>�[�/e	�|�7ƤT�e+�b`�D�(�r�����^������F<����~��4k�YQ��y�!�4�SL�K�q�x��C9?5?+p��0���~n��v~��&����q�y�i*�4�p6��D�b`�e�T���f@�7,ܵ58��R���5�Bq�@�97�	d��hf��$c_4b���Pj;�o@(��а�yy�j{![-��|}1�Z\�Yb�����F�Fs	�ɧ���K>
]��k��s�q��P�z��M��'x@��M�ds�dѰ����"�+��ĈM�C�y�[��T��t���CXc��\e�v�΁����K^]�V��"2�����7،�==����b��9����3��!����)�$eЄbw�7�d�+�6��X`@����C<�zS�5�,�ގ��S50��(�e�ƨ���L���9�oO_�J��>���۝ͻ�=6&k��M�&��-.��}s�x{$�b@�lf�E�����H�~"lB+7wO)M�\��oh��ٵ���h9�t���p�EYyM.�0��A�"������m^�5=޲�Ev�NRh�㹛{WJ�������q�O>A�ˍ����m��F��φf��Gʍ��z��6�7Zٖ�4�ɼL���٫�]F����[y�X��l�!(���v
J��T��7�`���;o���V-uz#:�H�%���/3Q�������8������E�JfO͌ϭdn��߼�N��nGlY�n"L&��|�&4:9z��"Q���h��<�������O\ǚQ�l8��,m5��Q�r����}�]c�hJ[����Fj�D5��<�X�k���j���S��J�n�����E�49��-d��&5a���ű�7�}���^-��p�Y�wtsjbG�@�V��׭����Տ~p�dtk���Jgo�s�Ad"��	mL��8�T>�9}dn{ؓ#1B9B�4����]`cG��N�=�����a��P����!�Yv̀�2� u����R��=�x/�R�ݔ��������t�WG='�{ G��QQ#
Q�1��0@Ox�T&i6ɇi�h^-���Ԃsw�+=e6��H��+�}�Ϥ�b�b1�1�ɷ)��6�����3S��"�
�s�!��e���fvP�,8�w#�W0��P�kC6�=��37<���ʞc�k9��C��������+|�_rzX�d�rD�R^��Wh���G����{�yM��g�J
��\�z.nG��k�A���g%���ͣ@i
���Fw�Rܛ��L��I	CdO�M�^Q9�u��s ۏ$	����}֤���V=��N�D�1�9
vaB���ZC�ͤ,> p�0�M���u��xJ�gnll����j�r�B���d13�^��MG�07�c�E-����S�4Wa�����$��ta��%�P�q��uxŰ�E��Y����8�XOfޠ+3y�-:�m��h��B�y�Z��h찫],�p�(e�CV������N�wq�f�Lb�`��������2E���Yv�v�L:�.I�ۻ��7�v�<�b�o���u�/w8u�����8b LC�
+�w��,��Œ�Da��9�8���}�t���Ϸ�%��ˆS��,���N>�o<�\�,ge2F�u&7Z�.Qr�ijn;7r�$��>\�u5{l�X>��۰q���w)T�c���Ƿ�:0�7@>m�}�<J���3�N>��vtS,ҚVQ��=u�g���駟Eؖ��f���!��<k�p�PVO�̦p_]7[Q޺�� �޵�C�úk9(��u��\8nv$�� �T%oj�Ո(w��i�m7�d��K�3���_�$�@�-)�������O
�)
`�a]�T@����4�y3�h�0���|!�ޥ�6���t��[���A�Bm�=	�F�V�|��ܺw��5)ʎ����^O��m�^Y�*�mIbIc�39v�jb�Xך-�U��`<3����U��5]q�5�]Cu���͹n���0��
�����1Yt��r��8�������Ռ<4.J�u[f��t^��_q��/-���P��U���>���z/�SoQ^�f��˫��t��C�.�Τ�*�j˫f�K�hKWJ$�כX�89��'^��bGщ����|mW;�A�e�Bb+^7������2O[�W"���VPLp����_(/o���;�sw��񫗒��*N�@L� �S�@��l8�;%����*�1j�=��
:�'AҳGk2����f����}����"�أQ����Y��nu�Tvb5��nG��fY˷f�����L
�ĩ�-���{��ߍ�v��=�&ȫL�+
mrZy�a�5m��Z�Q�ա�+-���/6�XΰWq�'Q<�v�q#�"�v$fWi�|f#�MwY�;}�#��Ҧ����cj����4y<�H��f��6��H�iyh��v�2�v�Q���57cy���L��˯�.�&ǯ���m����z�}�1Vq޺�J1kQ���u$_^��]�!Cq$�6z���ww\���n�C?~�.. �!�{�䔴C�jma�h�����٠��_����������ׯ_����_�������o�h��'*Jt�j�Hc4:ts9��}}z���ǯ^�z�������}~�_�W�}��%�J��H���ɣF�I��:>p[�_d(��IG���b)�X�lhy���r��Zm���'%�ˠ.YӉ��QP��^ۆ)��p�DC:�PE��[e�V�M����I�Ď��lm�F�ީ���.�l�i������9�'�T���[j �d5��p�CKCIQ�֨Z
��&��#PѶ���LLZ�X֪ь�(6�46,�s��gݹ���c�)�mLZ�j�T��)j�'��F�N���s�Z(6���p�tmj�y�y7�4��ZZm����lb�6uZ*+y�+/�����t+	&��ԡ����!�5$�X)�M���������|߾�]��>����xW<xLD�U��M���ߛ�bw�3�ƀ��L=_��j�LKɟSmJ��H�#`�D���L�"�;�s��s���2!?��^-�!kK��iLǽM̔
��I��SG�j&T֞9���{�a��k>�V��I㖮 ���ď;[�E.x�jUd;t����c!'7�K����C"��v�w?����+�a�'$o)�k�'��i����%����c�ϗSn�]�D38f�g����2��F5���Y�.j�N���|ok֧�>�Y9��ef7m*%)��ݼ���XFe��\�鷲^�y�'?�a���&���i����Ciֵ�m3�7�B2��6f��9^�qJ@/d8�u�>��t�3��݆15�D�g�3p��~
���	�Y[Y�6۠ʵ�Ba0���@h��l!��㠲�s�z�c@d(d������N6mL]�ٽ�8Pz�e�����B�t�$a9Ax�X)������\�6{��M�9��6^�fnV��!f)�2�}�f�,��Oti��j-��e�����9M�h��x�ٖ�����:�JPB"�:��U΄�k���m/�+zؔ��6� f�^�b�+F%{�HG��0;m��Y��}���)Y��N� ���Į�+��������e�.�����i��8zM�Arץܮ��%G�e�b캓���Y�S��`�oP̝'?����!K���P����Q�W��?�֞h�} ��&��)����Lױ����H8I&�����Z���u�2�f'1���eL�{-H�����]�h�������^�[�<f��mBm�׶�ս�7Ł�A�8b�Z��@n*��;b�y�+g�({�i�@�u�i��3��Cfê;��e�43nH*�#��'��ࢍ��s/�y]�f-�EC�g��FbZ�Z�Qy}�vZ5q6�u=w��+����[�������8�>:��i�g�N;�E.:��Y�\�+ ���鎒�Yo��3O��Ŷ���חf��*}'��ۙ�����z�q�󉷭���������+a�����)��n��i�tq)�x��6����$�9�-f�N�R��z�ݩ�����r�[ɳ�$вy��21� h���w6KBk�P/����]��c�$��M��3.z���LwP����я;b,
!��TY��Y�jA(�]@Z�X͗Wl_�gck�F;��x�T��$Ľ@��{�Ⱦ��ͧ�i����r�!,gfSKmF��Umb�҇{6�<U^�1ej�+�w3��.�p{���ǌ��{^JD��c��gnd���akB�Hb� 
]\��1=Cd�ϯ��|Nҟ^��Ryd����W���.V�bXd{:ų�,b]��vuv*ջ�Ƹ��Q�͹�^y�����\�"�������Ė���r�fҤ��}ܤ8 �oL�v�w�k3� ;YxdV��ke��pѭM1ɲn�e�^�o�%qSsZ�t�8���H�Q�̍@���j�%�#�8D�wp�Ԯ������^о���
W�?;ޥ:E%��U�Ѷ �	q)��(�=�����#xN�	��o1�n�:a���"=�/�D���],+׏i�$��.��#G��Q��9ԕp�J�μ?V�5e�����d]s;��r�3�q�ً����.�Ɛ��L�0�l��]ԻĿ9{dH7~��4�NA��!�a��Q%{Q��j�8���}9*�27A����r��9�^�"�,�T���mMO�v�������`C�DT������an�e+��2�,��qX˘Q/�3�y��-m��0�\��>&��Zޖd�i�ط��],�<���$����P�݋~<;ؗ�:��@���CTQu^}�ll�3��A�5��4ڎB"���8B%�m�-�G��Q�dz�|��9#x@�[�Tÿ�P��b�����a�qHC?a7{�*�W��v�IʓN�$L��.��ڎ�\��bBoJ�YӃ&
�o˹���"�����
�Cp}�`U�vz+���7�T��ƳE&�c|
Q���c8n!a��;M)�oDvl�]���#ދ	�Rʌ���q�ǌHC)0>w���O�?�U����k8a�c���j(�O�L�: \�@G9L���iO���W�;-t���s�䍆N��~����U" Ͱ�u��MLy�y�vU�Uǲ~��}�툆��/߹�I}6448�6z�ٜɢ�y���/�Y�Y��x����O#.���.���Y��;���;A\R`��a������]0*@w�i��`3��i{ZZg�U��5�"x�����>�x�DRS��u�%9m�k�OW��۴�X��H��^Xs���U,�AY������:��~������N�J6��1~�O4�$.���wz|�Z67c5�I�C;���5�"���S9�����]!��jnd�VStƞOgI���sW=˞3W��@PS�a�dC�wӛSr2";Kb
�	��O�m>�6�b�w��j�]gk�s�/�u�5Ņ�r�'��iѬ��8k�{d� #��w��Ur��4E��N�*�ZQ�a�E��F��� ��}0�t�dK.a����S\d6�jb�**����6���Y�^}}f��X�v��X�V���꧞�*`�Y���_3=Zb=ݙej���~�0!@�e=�G�!�ۮ��S�A.���4:o]��4i晾��pC���܇�Fʜ6e㷗�h�jݢ�{3��������|
��\���a�]G&�)�'Gc�����6�a�.q�'z��k\�O3�YN��yu���������Y����m�񳆃k�� wt�����l�k�Nm�� ��g�ی���:S��ó��X��U�G�u�\��8���ċ��9��2��jh�[
�_^1�(g9���5�ߞΪ����s��\���$Q~�I��Q�~˗�}�ٳD�x�	d�a�ǼO}(�|Y�P:V��c���PV��y����Q�l��f�5����>�&�$���_3�_x,�t�xV�g�K�*a��@�q
tދƞh~�\�$���!����9��S�d�r�ed�3� �{f�Pz���]�MEtٳ�+"o-�n[G;�㐝X�Ľ���|К�<x�}�.ڒ{�;�n�l��L���FGu� ����/s��Ζ�v+����*��0ͅ&G��H�ִ�l�;�#!�ٹ��<J��W}Y��@��ac�����<��5�	���w(�tq�ך��'�XP;!���@���0�X���Ը��k���g���ǟ���Pl��d#��<����5ud
�2��o��\�ץ(o��j��N�ѣ
�w�z�����Ef�NE�Îs��z�_w,�x�S�CC�g8������7�Ϟ�/|������ߟ��7y�_�>�$9���hk"�'Z�!��[J0'v��P#6aku�J�t���ĸ^>ԯnۯ?:9+�(K��`�e��نu�ޟC��55�`�M��b3y{趜ʚ�7� 㷻a���:kܺ.	�v���޵�1��`�'�6kg�K�2�˙Qއ�b_���N�'|�kA9U�g�"7M&��z��Nc9ǇևRy��*�=�J�i�/��i;S��a�S|��W����c����'�F��au�dYW��X�_�}����k��"k1�<b_;�����-��a�"�_!���ߛ5w��mND�����0�������b)�Vu�暆	��ĭtU<(����G����9��N&�N�|�h�ݏ
�9�����\��U�E��%��n<�?H���t�D����:����?�U;2��V�6�Z�QI�6�Y�/�	��$�L��������w�)�����R����fY�G��t��~UW�m2W��1y�ҝ���y�u�"��uE�xU��}1َ,��`]���Xƨ7&je߱�fZj���������ˡ��s[B.{ب�e�M�2�$iZ��j�s�/3A�B�F�*�6|��u[��e�֯��&_���;�5�R�]��Pι��6�E}���5���'-ΰ�ծ|��|��*��������q��s���8\5�����g9��%G����az������,e�`]��=�>�4�G���ϴ�.����\�䄪|&�b��6~��� ���t|Ӻ�&���|�'m�� ��R*��kv�����>�_�*��?��Ӟ���X���>�}���u�sԲb�v+ب�>�l����5��c��>��^��������1n"�T]�j����2�uT�p��Ml�x58{ދ2����`L�O��NZ��2�2_�u�le�ݍ-�r�lzW]�GE�>z���h�@BrV��{[29smz��7v��^��cڥ uLq�k�t�9It׹�ӭ`ɴ��X��z�U����ߡomW�|/�p�X%��b�΀֔�.�
��7��Ƒ�*��>��[ɟ[P��g�Y=����C;���������2
�̜�����zH��d�}�@%Dya�²e��*9��ج���:3�mh;�[%�]kLC�4�AP�s�Ӊ)\�Z�[}�l�yw�j�E���7���=��A������#�l�IF��sSx;����>l0jl���2��V^l��w�ʥy��>;X[����j����_�Cͻ�LT:�ʃ���f���;�8;���7_*�}�t�K��ϫ������f�n������ ���L��>j\3T����hU�_-�0�{��a�񋊯����x7���>&�M���U}?vƗ���`oHw;~��3�>e�#Ϗ|�1�'�,3�yo2����Իjm�+6�Ὥ���h�k�&5T�z��
�/e~�R_��~4���tR���1s����k�ꝋ����i����O$ފ.�Fö1,m�z�rP��7,"7&�;"�%"�����%�셕�!�[#�˙ټ T�N��U.C!ү*���jQWi�����d�Ӥ�!������ ���F$o@G%*�6�w;��}�92��D�W{�cH��	��M��b�xs׎�ip�D���5U3R�װ�v����ţo'"�ó��-E�f��ae�;E18��S@f�F�Z��8E�do�C����UQ��U�o��u�9b�Gr��Jִ�oW6D�Ow&��S�0`3�K�Ec��+5Ǯ��fUz9�̗V� {��Z"$r�Gv�Rd7U�ó�ݬ�L(��Xkƅcj�UF�L�i�7L��OAѹ�^�vCO:��M����v J�IÕْh4΂��D3�p�c���J43���;����+�U������N����kқ�͡��˒�z��Weh��v�JY���@U&5]@�&�6)c6�՛��w2{0���4唔7�.M�곽�������<���;�<�|��y��w�����>��s�J�$����X��,4���צּc��Qb��
t�W8|��Z�Z�>������	f~=�jy��e��:ss[3k�[q���C3#��3�
D�l[.t���q���|�|�Î6D';����������d�An�8�>��d\��^{ؒ��l:���k�_aĝ�U>c07cyq�����;�'5�O��\����Q�9��;7�w��t�A#�Y���������cë TlG�f�m3��휲�F�Vuj�YFu�O\��p�~֟[YQ} kl8N�5&�=�6CO�"���Ar(c���{O �B��h�v��ױ�@�.�&a�\�I���Ω5�8�o#�M�	�K/��5u��������E3��Ju�UC��ŇV~�睎����]�{o:X��@�LntBjW�.v�-k�dG$�_Q�в�����8�h�S�-M��D��Z�]|z�ţ�71���st�n��V��/b�'}��ԭ�r jzwx��\��E�$`LӉ4�3����X����c���J,!Z� �ƍ��*"�h�s)t�pu�P��uݎDr��В��l���t�[y��ʊԭ��o84| c���+~�w�{Qd;�@G4*.=�H������5u�ޖ{�p�5�=��d�k��f��i�)t�����ޗ?y�������?ۏ��"�n�.�iA�}��M m��Mn�Q����2��yl�+�fv�@�y���MG�� oS���Y*)��B�f8�a�	݁��gV��hEkV.oE&ۼ�4r���k��b��v�N�l���9vkq7p�;W�Wq�����į/.أ���3��xMd`���@ׅ+.tw��Z��Mg1������`�M.٩me��g?�Qk�����6Si6(	�$1�J4�0�Ͼ�׈�ik���v\��e(��B�L�\�^��r#u�l����Z�7��hN�1���C����7
�mu<�[�� ���^�F��-ˮFa���V8�u�0�w���w��{	�MKN�6]�j����|d�d��!r�Q�%��#����nqϬ��5��b�M�ɷ�[��{a�����*�(��e,��[dn��|�H/	��s�>�:8�cz��f;�+��R���,�P��y��kaB_'�n����#u�0����if@{���y�4�m���wո��5� �A��18�k1+_7Sl�O���zԌ�m�������^0�4���?�~�ʵ������z�f(~�7�W0\��}N�r(�f8�Ej�lN.Q��x�jT�����w�!G������{z�����:(oW�j>�O�j�Z�D Xf�&eLۇ�����v�aR� 3bC��3�l^���Ci���n�d��������5��j�H�n���Ζp�^:Tcz��N�^�z��P �Q�S|�\��6�ݲ���ehp���ZKڝuyuy;�V �*�+��J���][\��e���ե��ewV��8,#C�? ]��L��n�G�WbRܵo��R8��26�����A<���Gb�J�쏘ul�H�>n��u}��J]��Q�{5�E�]�p�7����jw��/�G�FY���u]�8�p�_P[Ov{p�6A��x��h6c��M���'Ne���`�%.CN^ff�Z6��
|%f��ڏ�Jt�;��˖�.���me=ÀVĕԛ��5�=�,�ZU��t�Yf��1��צe��$E)z�]����J�mɻ�M"-���ɉ}{u��Fr�)R�@�ym1�e�p�7�ֻ�,>V�޾i�B��ҷx	Lc�:틤�ڡ���}֩��2epE��W"�m��kv�r�J|@��TWE�^-�;wl��蹴ikfK�:U��i4Sl,�@�e� m`��\����W�%�wV�l (	鄢�I{̴X����t�Ȩ�<Ib��
�U�DF ����&ʺ3��DT����O!F�R�Xr���$8οh�`��EV�K!"ԸͪT��"��5[&+��4:�'��A�b^.M�"�8Fwۖ�kj�5�����! %+FW�F�����O-�{���lZٲ��̵@�s:��e���&sU�q�+���
ٰ�[/��)/Ck��+U�u���4��{/	ѡU�e}��]Z�R[φ�Ԍ��٦1��#�C:ֻ��x`.�7�˰jkn��0��vx�eϫh��ek�yR�۫H;��a,�ԎP���;p���"�"G�l��jv�w��܄Pr�b��^��d�*|{��c�՚	��m�o)���A��:Ԯ{[\p�Xhס�f�¯�<�-�*v���Ki��ev��R�:��D��x7@�qf��d��̦���>M�I�YvZ�S��;�d]%�֬���E0�޾9s
�)C{y��;绌u�/�M�*�-���
��V�
���,�J��˫Pk��Ρ {�L�7i%�wS�آ�ҳ+:f��3;4��B�`��9!�p�v�<r�O� �n�5d��6�3�;Gu2��2��b�Pp�N ֨��5j���7�$�����K�8͂�*L�]Z'V'�[m
U)�=\�E˔<���z/5;��c���6�V���/�����Q��h�Ӧ2t�;���ᡓVMQE+W0�Z�� P�<�i�A�I��h[4F�AФ&����
`1L���I/:!�4�4)�h���A���f
2��"g��9G�Ly8�Alj�
�hi�Mi���B��⠧l�͜�����~=z��ׯ^�z������_�������6�5@M���5�f�X���h6�!��hi�3���rj��IE39������ׯ�z������������~�?>���.G6ӧIQ!���uC�)
�k�9SN������E�Z�P��m�������!�$�^}�s�;h�X��\�bJ(
_1���j����٭���$�AZ5Z:kK�"�������j�+I1N��j
Ӣ�AmV�m�i�֠�C��y�:4�V���DTkmkm|�._6y(�N>c䘂"�v��h"`�.U�&�6+���l�����\�f�����kA%O���X�4RĔUV����n<�*
��[U'9��&����h�D�c�<�l[Pld�p�@DIQAr5��1U��Z(��=�\ؘ��ETQL�sbbj�=7r�@9t�x�ȼ����`b$Z�7�H�+�hs��Cj߻&�[��hOu�4����	����N���"�$Q�r�sks����3���P���w�w� �V �Q_��q���{he\�ዀ���"|U14vS�ft��sU�]�Sg��s���n�f[�8]Q��`_�qd�ЪШ�gҚ��P�&�w�VO���|��4��U0�����{�<J�[ְ�f��;���*�����_�ǝ�<��!��74����P�-�@|��.�f�p��	7,)��8��X�e�:N�"Z��ڞ]��y�%�]�k��ה�iݸ�;Jw���ҚH�s*k��L�����Y��!6D��Y.�bQ�*d���^�m��Ϊ��}�Nm��w7�׃<ܛ\��,���sU��l�W#$��w�/u��ͪb�E0���"���'��T�c���Kĩ��i�w�u�]�6�W����l���O�߿*P\ٮZ�`le֡Cת,�vEm��n��&Mܞc,FU�YU79xZ�Fû�p���ɝ�y�jp(�d���+��P���y��Q ���h.!�X���-{���lD���ѝMeg����8���y�C�l�};#�,`؝ݼ+]�8a�F������顙���ow2�4��er�VH�j��\�7��C{�N�[��\z���쿓��h|�m>N�A���w��4����>/�)���=yh�b���u��v:�ےg�R�B�+���}�{G!��A�������[@<��͡V���y���|<H�j�.��[s���x�T�&�N/ս�7�F��K���B2l���,�Ɔ��I��ݾ�ܧd0���P�"#�K��n�/������Wd2iI�X]%EFQI����QkU�dTW���^l��?����mƏ;bh�4z�>�C1�S�L7<�9��߫)�$�R��
sx��A�L'<I���]4��g���B=��/�~7����{0� ��ֽ�F3�+�ꌲ�`�=����XeW�>���eF:�7��U:|�a5}I�F3xͩ��֥���&֨��(��ͺ�I��29�������*�t����?��Q��~�qs�B��8+�'�\��ϣ�M��ٱ�hu@���1�]4�;cd�b��ۤK�)[P)��w/ �ۦ8�?�{^<g��]OB��Ǫ,=��y�o:>'7�-yvE���ƥ�q�\&h�B�7�x��q�:V�|c5�8��jN�\�F �p��1j�M�m��ٗ7�S��!�����wh֖j$ѣM�d;38ާ��	�Iexj��W4d+��J2��A;bV���h��yi�hF���3��c�VC>3�  j|���p�^>��
�������ǋ]Ӳ�6���u��[=*zdKL�n뻸f�����g��1ojSR�vg�^%�vE��;������y���G���n㻹��6�-x;t�>���fT5� ?qʈR�]���n{��M�7)��x��C^��.��H^�~*��%2a5&�}��!O�&��}��0Θ�
�k]�WY�cs�i�N��AB�S*n�[�#9ִ��a̏�ʘG6�*��{�7P�y�9�c5�YeQ��Qi�1U�-=���,D��ϩ��pՊ���Ѽ��SY��N�P����̂_S>���q7Va�T�~�>�E~���̘p�1��S9Q�*4��t�o)��6�T�L9�ξҩ�%Ǩx�g�9�d"[w���1�9ng1�Ά`wҙ�C�𫌫[a�9��u����/r�i2eF*Ѽ���+̷��+�̤!C1Q͹�e�u�O@,�U�\k�u^UM=��|jHm�^� ����=�mu��< �S�\N�Y�1{|�ի2�ܪ7��ukT{b�f�m��[�]�	x�٩�S�^�|ۀ�@���+�?�ݽ�u�] v���7L�ߙ{������U��%-��Ī!�<T�@r�[���@]D�χ�����'.I�5d�3N�Qt��lӤ4*�[oP�Mmv�v�t�l�!C��Y���E
�r5���D�W;޿Ն� ����7t�7�;zz~~�?ϯ^s�9	@~}�������5��s��'#��]���`�����}��V�S�/\.�kh�gt6l<�4�F������p��3�'���u�}>d���\�7�6��t�n�1��н}��I�lcݔC(z%?��_�Dͮ�猈�ͽj�y���}�NR�Qy�s��[L�w��G!�q����V�z��Y.
/����f�1k��{t��@Mp�<��wTr��Ye�֩<xM@�H��w����\�{�+�N�@�U�es�N�J�zJ��]mlrZ����Y�͗��M���m�����hhU��pk:V�������)�<ϯf�3�勜��uь��x��k��=u¼�<�N��Wgw�׻�WLk�4�v�h���|�ᛎ#v�_i<n훗K�u�t�wN��< 4A���ۆ�Iή����-�����7czD��]oESD�yv`e@��fP���U�}�⓺�1{vHU;Q�ǻPwn^-�!\�y9V��\��Z!w��iЈ��}AД�e��R9ސ'u9ƄK� �n�2�N����Ү��A;E��6��J�cj��v�ʴ�_���]Ǽ����f��vd�>\<ǜ1���/9ß������8y^�0���͜ߴ�]u$c�AStH��?�~���ǉ�JR���Y��0]x�3�^�^�g�ӱ�+p�m�t�	����ڲ���Vüv�GoY�����'�D����Qq{{{8���x�als .ށP����t5�U�Zi�-��R�B����gOf�\3m{��;w�9�_��0���ԯA�����PI,�Y�NDj��W4�Q�Ӱ�&w��	W����{��Uꖢ�e�ym����e��V�7�k�ʝH�9�$�ê�x�YYp`�c�TO\N�ǭ�!y��׻�z�7��(|$�V��t|pk�W[�zё����U��Y�r"6����.�Ѩ��7P��j�V���mc]7%�Ѝ����=�NM�MȟM��*�c`?;��uʠ�	��ʟ��>��1š�tڌ�g��b�Lz������\��æ�*3�Sߪ�v��,j��T��!+�pX�,-�
�=�[��k����9�إ�9#��!Cw��B̆E۽��,v�����@��u��.[彽���0c�r>�j.��|���c\��YAl.�۱�n7ܺG�RV�6��k�ӷW�{��b��nV���O����֦�Z�*bg�ʪn��
�� �>M;o�p�}B��󉈘��Ј�Uk<���fo�b��jrTΩ��`4z`��e,�	��Ä^�c��k����g� v¼�܀�]Y��@>��1�,�cQ���oD�2�Ǯ':sq��Q���@�+�����O�k��j3bN�=wpۻ�U��̷����$.�[�ٰ�hJX{�Xn�,����8�Ʌ,��T�Ƀ̻<c������4-�#q�t@��$
�QݙHح,̳���-I�'��Wc7(c̫QZ��H}r[�%��V��i�KEnϱr��/
�\��Duf��h��}��3U?Oar=F�i0ʻ��%����W���d���幾8go)Z������w�Е����h]����ޛ[���­���ˡ��nF{z�4��f�(z����i��Z��v�܌��֝7��Q���.bm.���;̱���]yp>T��:85�ȇf��P�8Ո����{�kU^�afrd؝���\�:ޣ���'7�w�H�>"n�f^y ѷ�-����5+Wym֐�}�|�?�o�n�<�M��z��l�j.����z�f��S9$w���X2��]��n_T�3�r��(�@xGUl��.���rxLK+��)�k��ׅ�u����K��쎙-�@�E8���ͨ:�;���vkl[=�ݛ���g'l�����t3w�d�CU9�&��{=W�-5��l�\D�����6d>������*�%w+$��X�$���gTJ˂����ڍ�����sĶvW>�,�J�:�)E��s;���u���=VT
�ؤN��[0񻅶����E����Wmǭ�'����������g7��S��-�H�����`��b����b[���p�I.�����7�n7���.�������I�2�ѕ7���zV����ܵ1+ǥ6o����JG��znw�;��G��`���5�(	O}rG:��n����2�E3d^�A��/GP�4���*��3��n��B�S���I��Wk{��\t����E����(����)X�q�\y��僕���>���U���w�u�˜�S�"���U�'I�z�/��p�a�c��J��w1�IZ��-}�^�o7������]\���ly�osl�����)����Gv<���7o3bM��V�S(>��V��L������>�m��ԥ���񓾬;VsOG������f��tO�� ESf�
�v�p1�����q��O��Ƈo|�W�Uk}M&��:�@�ķ� -ȻY�oc^u�޼��#d4L3��K��c�����2\�n[Y�z��/ܴ�.��76��;}�1�	�k/u�cC�@��wU���S�k�Q�{ps8t��uO���-�tG>�g�{<4��_76��=��{�Tr�uC+��Z�3உ
���S�}�=2���>R��h�;ٷ�z�r�+%��ms\b��~��oie=QX,�6�N�Ɍݭ�Zy��7���U}ʡT����Q�}l�>3K������R|��u��D{W?�f��k�S���
���9<��T��]�� 3su�UŅm��Dp{��i�`��j���0f����8��-��Z0Q�]�8�mUY�g�pX�$(
 vq�)2��Wz��r��������D���]���S(�֮�/y�I��$>�k�߽c��ƾV� ���b0�R�ES�:-�X	�e����^>o7�s��(0����LԓC���[���w�30�5ȸ�	��־�Uc��~�@�c�v�ywsY���>����23ak�1ȏpZ�.g����q����[�]���0ֳ9Sٶ3���v�O�@�L��~�)�ƽ�xw�W�hMi��������	,��� r�7c;\T{�k���We�YV��gV��:]���[TZ����˲�X�7��kܣ)�g#"Y�VE�͂�@=����D�|����=��r�����Y��w�1v�3[���WS�lz�ݯ�H)�pȧ�g>�B��������s4SHVDx>�T�ٽv�����*��`���
v=:�-c���D����y�o/n�XL �c��W!E(摾s/���I��h8Iĉ\�0W�oM�u=f�T\pWs���Z3��=��L�]�02�ӮX�Im�Q�0�/T��B�҈�����`�����W�_e���ٺ~��M�|�r�
ܽ�ё�������,.�����\�Ձ����k>M-��fK峭uj5��!������0����5�Q䮹���>�/��٥v2�y �o0��k7�GD�&{ѕ��-���z�-��o	9H|�e�!M'�J�r���m����G����&R%���)Gb��}!juE-�:��p�d+˷������^x�
R������Ff�����gs-�&��]Yt�ݴ����ls2��lL.N%������\�$��g\�d�����ouuU�xN(�m��gK��zU��rJʙ�x��vj�ۮ����2ej�y��~4ת�y�ʾ�YY�I����N_C�q��չ�u�;aW�;���^���~9�k��RTΉr	��zZ�m��mC�V����%9�ݐ0�O�n�oR�/�lw;Mq�}y��:Xk�D���-���%c���y[�/7n��g(켾=;{��i�;V{v|�lB��>��k��kf+�D���OY\=vDF�iSo˄tTWKqu|�1�����s�S��Zw��e(%��Q�t�f���A�·7��U��no���Z苿w޶s�*�>9��E,*Gr�e�w2�b�{���x/���|���/�`O�gM������T��*PnN�<��,�ϴ���Y��}0Y!r�oWSg1��A���L����`�	IufL�J*�9*=��t�?vA lw��[�^^��t�L,}�
���r] ��ٺ�n�o��w��/+{�M&����.��u��QoU"qZ�ܮ�Q�Bz]('�
�]�X�K��:�`�%\4��+S+Б���ɬ��-+5Hv\��&�\w(�]Q� X�Ck�����闚�q}s��v3���R���3�ͮVA��d�]v�{���G�#��a��7�K����wD{�J����`Yk[�@�t���W��m���*�̚�b#�ut0Y�1\ohT� m[4D��{
U�,=h�y̮x���d_4���"b�N�6v��ή��]9��W���l�N������֊sx�{s���'] T��ۭ�93:�m�use+�;K��b�^WR���`U�i^����b��r��~!C]Hp��_5ϱX��k)���[��hي��ܭ��l�hf�=O�7lV���g���%��)����g[�Bu�x'ǒf���@��ƫdSVu��^-�M�$(��Ό7b��^��x�,t��mc-�T���yP��e
J�X
)*>��_��g�����5ߕ[]��q����Z��%����H��� =��a��/!��`����k{�
.�GKȉU7���b躻���d��
벻B��ԉ�n��נ�S�<g����n�����Y�k�d\��U��K��*f�yf0-F�|4�lq�����x	N�!ת�n�.�·*ac�d�F�$-P.��ވr�Nu[cJ`���+��b�����t�J���.b"V�����&YD�M�VSR�Cm1/��uZ��a�[�|�0�u<���b�pJ�º��{�	�����-��:��'�ݖ����C�D%ۇ4(KSki@�N��M�<�Sξd�y�w,�I�|95�ki��{$��]՞�s�N��m�s�ͼξ�=y|�v4N(���&��+���ZD,�gz���`�Uw]{�ث����}���gdym��xJ:nA���9º�똺�Asn���U�Em-��N�����3�C4���p�E�}�ڀ+�cojPՃ���CX�}�j�
-�O�^��Y��ƽ�vek�
�N苶��^�9��y\Ѥd�r�h�\QMM�:��摔�<������#cL��OCX�� 8��G��]\g��U�!���{�L�j��=ɢ3�\�=A:�+����q7d����Yvw#�RÈ͜�c�����
?�yUh�
*��Am�@EURG�r�U1TU4�PE��j���s����z�?_�z��ׯ_______�������1�a��n�s�*�j�4]3�lS-�*���b�j�Z���m�`���}~=�sׯ^�z�������~�_�N�؉��SD}��QDTǑ�N6��E������b&�>��1QUA�K5EF���-:g�nA�a�m�|���J����<�O�:<���DQD��)ы�uQ�SDUZ�A;��DT^â�*����IL�`��_q�-�0m�͊
���
�D�͊'��s`�(��Tr�JKX���&J�.O�8D4y*-��(�b"����p�W-Q��h��G���+��[79�#��T{�4�[���3%�j�������TW=�J�<܈���'1嫘)�9h9���؝i�I�h��ITU�D�h�h ���bm��(�$��EOV�����aVަ�;����7L�Υ}�Vl��1��뜮W�m�y���ܝ�#�R�]W����MV��G����x~ *�9ä�CnW����r ��͆�$;o�S�ly�Ѝ_t��^�1�j�m��H_q��0���5S��k��;�ͥ�V�k��0L�ջ�M;Fc�i�5V�Lݭ�<�9�0q����;ܬF�Dwfg4��{���O�G�[�J�]��V�y{~�42^;􀜩���/:����`	@Qh�3����D_l
BE��O����E����q��m��tc|.�/�9hM�ä�릅w��e���<�t�L�ڈ��Yp�]���}y�rǮVA�k�C��mةU�1�OL]΢���cN��kC�ML,\p��W_�*;jY��= 5S��j�oC��=?>Ine՛w�cF+G����RuR��JWs!eq7���UG��D4�c����b�6��4�8=��f�ܣ��O���+��uR��.�h2?_��G�?=�fKZ�A�^v�'�����������Ѽ�S���@#���<,�@!YK7���i_n�B���ו��o��5�m��+��֝����%��:k:���v���(Ym���|%��w{�n��͵����>^���p<��9i%s����-�/C�;"mu�mJR��(�UY�S��#��m�~ۻ�l~�S�Ni::�V�@�l�ހz+����32k[9O���eؽϚ�{��'~��>����ᓾn�]�+����WR�Q��cVZ�ݧk����ۖ����1����l�$,Y�m���0��m�4I.���T��Mep/�{���O��WA�����Z7��r!��Cz@�B"�a�ﹼV�[J^���,K�ceV���R:�L���#}V���g�H\�����ݣ��K�W#s[��z��5f�N�cT�/6m^)��3o�SK.�����x��T��tUs�J��n`;}�kVP��&�Fv>nv�ƼE/ ��Cq֭����Ӑ��b��7]5p��Q#*K�ʽ���>�:s�LW���sh�ɭg���uH��"wX|	�:�~߬Y�2��\魤�3�-P��Zm����8H�)_ݕ�d��.�����N����iÌ�}�]-�� ��tWr�e\��LŨiՒ�oN�{
�kx��k�px�R�������xм��4G��e�mÝ�ӷ�^��2n��Ԍ���|ǵ��k�y���^���s��l�;���Y��&��.�3��z`n���<���6P��ώiL�����/T;u�>�m�(�M=�?��s��. �y��)�j�n�7�����5�v���s{N�9<��t}�ߋ������w+=���{{�rf��MV��Ͻ3Ux�9�n{ƭ�$c �<�ؽur1+���W)�bi��u5�" 2�w�����e��=�S{:j�/Ƚhh�����=��4ylI�q�m�+x��~P�,ޞ~����ʡ�,�Zt#�/����w�Z6I��e���W��8�����~������~Y��Ύ�Q�%�u�#��WM��ᝅ�5�/#��޵��{2}�r�9���Y�ǩ̼���E�Q�{�ͰnXk1����yC�*�cnՙ�ͩ³7�Nݚ�)��,^fso;tNX�����֛��Z�E��U�Sݼ�~a��OK��a�C�ۛQ01a��2j�h�YGd���M�=�ced�o�Ȉ�zv�GBq9�4�ߘ�����.������w���;��$�g1�K����^֩��;�[�zK�83`����e��]O@�����2�m�������y�.�m���j�-�z���kt1]͸�	�ם��w�RQ�D_4���2g�+�p�F���\6�/0�9�����N�?�t�U�(f���;��׋0c�,�7�<���z9�6p��0�&|�+�vC���j��K�m]6֊5\'S�]vP5����T��.�k���W4��n�O%�c�F^uLN�3�.�n����_o
��$?.�d�i�S&�����k򞜽�<oY���<R�[�6{��y����S�ȗ�;����O�
���!ހ�_���[0a�1�%w�<�Er�g���:����bg���2tf��Ƿ��94�Cn[)8��=�QRh�F���w�k/R�잵y>S1�%_���-�z��ԫ� ���ic��ۚ�xk�\5�����y���xZ��UQ��婻~��Y~�����{�����Ipq�p�5���& 7i�m����E���oˀ�_!+�Z/�}�X�O֞��.P2m�K�}��u.��sE�Z��mس��}�Q7�I�[�3����ۛQ���F���+� 6����2�,:M�w�x�����;�֕�ҩ�����O|^��c>�)��+�lJ���;�^�5�h^��ݚ~�睫��f��-^�h��o����Q�1�޿�J�ĺ�\K���*�+3TL����I�#��]��+�xWt8 �nҵ�wj��sC&9�b)ⶖqj�go:W�����8;{��-�#r�=n��}�$�v��*�7��vj z��,�:�Y����o����"��Cx�~���bpHy����'{z�#�d���̸ԏym�|�O����c��һ����r+�����:$u�]�dk���c� $���w�gHl�� 0�u2UȾ��2o3dl�t5hg3S��"���[�*���ܡUtsHe�SݭM&�� MK\�F]��&$�l�un�7/P�{�/}�4���h�������t6��M�ھr׎�Җ��q�Z��{���{��j{٧�L��`�mͼv�8v!�,9��~��\i��C�]���u}�oYPZ��Ӥ)U�Քxu�Ζ�*xws�Σ�]�٠�3���.��A��K�T�J/sk8����g+݂V���Vb�4��K��������y�s�ͅ�"�����g�:X׶���gc>8*4]&k��L���Mm�lCR��y����y�co�z_P�e��,��@�1����C�f̨U�m�m���V�q�Y�A+ؓ�l��C�x@Я�U�]w2Qg�A�<����/Mvw���m�O��T捾�m��J�a)�=wL��Wl�4�k2�0�5�6E��9� K%�"�4�{]��gԨ�fג�$���%�+w.�C�;U���!]H�Q<Fn��|Kc�w۹6����O��+sz�7e�R�[���Ѕ۳M\�e��n�{��4`�]4�ڨ�+My>~ݵ �uϛn�y^��,�nU�;f�wY��bN&�3J�h����;����Kv�ʌT&��6 �~�׌�#���zu���f/~;��_Nr�����֚��������;ɐ�/-����0�s��]e��K"y�^�#1߇�0+\�	�xެ�MZt`����[���c��P�"U��mo�"'�o�"�� sf2�]�ݖ�=ӺJu\[<Idj��m%Xz�g[�gW(\b�v�˾������Ü���Vy�dE@��;�"��!ϫ����{�L���Uim���J���.r����[y�f����V5@���˴�4��q��Ƚ���u�����s�a���0WYlU#�י�ڞ�Ȉj�;y��k𷝁�"��Fd3t{��<��Q����"��P��O��9F��g7��e��ynH�(r���,����=���<PZu��w��o2�N���x�_!��Ы��CT�̩۠�M�ͧ�g�1�h>�%v�\��&u�-���y
�ww��yu�@�LϽ�kqE�<��8�j�|�K(��
�4�
>���C�c�HoH��r�����O����E�w}:Kex�����&��(�ۥ<ޥ�tu�p����fg�żU�OflS�C�0,�����;n�Gm���~<�Κ<�	�
��n߶q�\x�i3��ޖ��ƪ��{�sd_Mǧ)d����2,c}��������=��Х�Kn���_�z�5�Y�2#���F3F�R}B���ox�#7l3��40����'���^��YԖG���j�O���gV;-�}H�Nb��ckU���f.�r^ul�V䑾ۛ��R%�mo!K��]��N��//~�nM\��ա�������J�՚#b}S�7�)��V~��������=�Mc�١)~z�;L
��3em�;5��f8����ީ����y��SϮ��y�C�������اו��en�N�S�w{i�X���z!s;4�ݖG� �;co��ܝ�˶��˟hU_N-U��TufT�A\�)T˿dPΌ��h�X妝��+�����g����qt�'lO���k5S�CT�4/Q�K��F?����;��a��\\N�NǧRT2�f�u$-��ٌٽʛ�7��;0����Wq��Z/���&�@��Cղ���E�D-|�摙�Sw�c'������=�1�S�'}*xgl�Ł�_9����||�A�4��6�d[]Qzξ�;7��!󥓶5�5���N����#��g���4��ښI7��h������2�E�z����O�G)�L���_��\�ؗYDZ"uܫ@�=<���<�����K���W�^9 qN^�x�k��uu��iI��p���1Զ�+��8q��Gyvt{}��NV�|-u%���Gk��̏p���o��b�FZ�*����09��v��lʗ�7�����x93:��5b���k�9���c��Ja���%5�w�:��^���f���d���َ��}l�탎˃����rz}=##[-E_N�>əc���g���aexyMX�L;��_�'s�i���ў��poyz�!�+�կ�{�y.�-ND����MSG��5�m��X'�5�v}�f�``��|��"�0:�+�j;v��������q4�
7uyks9���y��f[!����=�7�I�g���rf,:M���c���s���禛t������uǟ{6��=:�ۭ}
�j�F�uSQ�f�ɥ=���<yR�v��#�lp�t��.w���2�UF*���oø���YI'�3�//�a�sK���;�ic5]�;V����y�{�n�����J��.5
����o���>� �WW�.��E���k*{^ kw�ᱶ���f�N���� �r�L�)�%WZy|�.qeLpX�z��د�S��"u��%�nNL����Y�X��*Bmh��7�.�,��z%Γ�6��ے��V��۹��Qj�Eǣ��?���#�s�B2��8�}�O��O�k�W�����Z��q�!�=��P}l�'�vdҭ��B��j��8�P(Wt]�ɺ+`f���xe����čq������	&�`��c�3�����,��*]���硪���Ն�%;%㡁c���Moz�Q�����w`?rg���_�ꊬd��J���F^;O�ՙ��.�E,�/�,�d���E�c�(
�7a�c�U>��v��h�����u0�jY:��W���K3�d�UXګ%�A��x���lܓ9j���������X�Oc��:���T�<�D��H����c?b�G��\��~���|G�+W�_F6�f�X�D"3����3��PC��?}T��X4 R���V��[����3��d�Yu���cY�er��Ylu���އ��MDt��?/o�ߎ*�>�~.=��z�N�K;�F�����f^$Q�`���u<�8��m�Px��H�`]7�2[�U�y52C���6ګ۩$�fl��W��eѓ�ۇ�oZ�q�'�eEN}�`�!��f�[Vш����v��U�PZ��{<�y�7����s֔�����wA� c�x˚�x"CH���P��5�>rYu�	��Ͼg��|�r0h O]=�* �uB�ֱ}Y��뚙1u��{or�ON�r����o05N��@�X�Y����ގ�!��讀��.�I M�YǓ,�+t���n����{,f�N�ר���=�e���q79�vt�9��" ��3�[T����$y���t�w�l]Xy�ܙl���.��ZmU��@\�!s�2q�%�7#�*.RZ�v�M;�к�Z֡Μ��U�r^�^]��YZ�쨵^Ia����P@t �������Ʃ�Fe�F��@M�N�=��ޒ��U��qa/�2�D0�����w���z�..��RvS��r��f�C,I[BR/�h��]Q^�RO��c�����8�>�+ '�J��O.��2〱pH�`Ǣ�Pi�M٦p�\��Rp���Nb�Z�e�i$�w֝5���7[�ɋE�Ǐ�uw�\y�Y��]W����%2���K�����E��Ɍf�C�NE~���TI0b��ӄW.��C�I"�JE�L	�0�v�6ԥ]A-d��z��f��!j.nK'j�Ě��WA�B�Z����RwQ��	�ػ�:�!E�= j���hz�+�[�Q�=s��:�<6�]Oh�����QQͳb-��.�.��]AP�c�R�/��tmt��3��lNe���R�e���n=U֗po6�3�!�K��_L�DV��j^���gX��ku"�w��D��҉#:��u��5������a�^$�v
��ޕ�0�n;e��-;}u�<�}d�ΐ�Z8%��)S�Eg"�;�!Bv�V\�R�e2��Ϧ�ʍ�qt] ����P%�����.C��ơj{���4��n�Đ۩��Qw��@w��BmHsfC�U���j��7��f��"��r�}+"0kx��Jʻ���f��ȫ73�R��zڴt��i�q�q���<릗 g�Y�Bl�y��Ş�<>�/{GgnP̏��@9;��ܱX�f؛I��C/{/]�m��C0�D�x�*PH�k��q�Y�W��q�z�$�S��À�$��;.�<X�p��9����wJ�m3��ݧ�BB�AYʲeF�e�Z����)i1���`P���E�������5�U3DpK�q�������R��u��X㧱�o2�V��7Wn�L��e�\�����/'.��޼Q<����,P���N�a{�j&��s���u�z�ޜˮ7Rfx�1�`�[ԭ[�H�Z�*obf��7Wv��d���]��qw��,�X�$�gtV�qa�<���Ǚ =X���'gw[Ģ��ޣw�{����Q��rIp�/тi eL��&�&��4�` �Ӧ��N����x��i�l�(y �:E���B�(	@�d�2EI2���c���;jj�"��1之�s�k���*�
(�m55MS��������_��=z��ׯ������_���{�����EQF�?e�TQ����1.�-nZ����j3ss�5�:.��klQs&x���~�^��Y�ׯ^�}}}}}}z�~�^�ߵnQ�#63���Lp�����ba��cPD�\٫����y�@}��ɪ+��DPQUM��f��6ų�b"�\�Z
�R4\,QV����f*
���Y����AUD��&(���`�30k�11M1Q��"�`��DD�7�T��5V�/7�tQTEΚ+��T�E;j"gY�b���B$Ѡ���٢�����|�ZZ����y��">A���*Zf(����m��5Q4PPQ\�� ��lmD�X���%TT7��Z�ј��1:������˜��X������|�xI�"���#�Dj���:�V��=�m_��.{�4ѫf#g0�h_L溸�w�T1��sg�݊-t�E�����V�9���t�퓢�K�uM�
����Ð���<.N0U"EQ$$Ӡ#��~�w����G��l۽1/U����K�4$�Ysot��+)�c�u��׭�����[�|R��I4��<U�Km�o+թ����C>�5����)�!����Q���|������]d=��̒��lɼ��@�o 6
���mu4v�N<ov�c3\��A�TF;]�߫97�+���i���7��t��FV��㱺�|�y�AV��5sl�����]{��fVS��lM3u�wr�/9�^��ֽtE09�혵>���\╿��;6wp�KƘN.�]B�ٸ�����;�*��6t��7�-��}\��.;n��)��-=ӹ{]8�z�v����A�)����;|s\��mٴ�r��[��^OV�`���׫c�v^���C`f�Qʉj�Q��2��]��t�*Kݥ%�������L�W�l�:9�v���\vK(�]�r�hW��������O+!�{c��%`����jY-EZ�}�7k�=������H�쮤��*�,;9PzoUj�w�`z����NR���3�>��'%����V^k�n�9�3��3ب��������c�����Ke:�@�~�y���ˬ�Ύ�7(5�׀Ҧ�E�1Eu?��v�Cz��%/ʹ�c���9�g{9�6�C9z��,�/���3N
�XH;A7�Mf��u�]B{�M	��|~�ͭ�ٍ��r}�w2�h��P8���O���!�=3��ͫ���0���ׇ�T��Ż*F�gMs�n|�K$j�~́7|��/�B����U�p[�tt�4���,+=�܂�t��j�X���{n��g�9��t-���݇~�x��3���'��(���1�����]�2���a��Y}SS�.N2��{��\C�]�<B���l��>)�FyO�X����պ��,���jaV3�P!kveB��y�,��KS/0|�P�p.FH��ŝ�}�\��v{lC�m2�Ӎo����v�d��Æ���w6��G8��xR	~�h��ﻶ$��E]����ѯ�-���v�/ן:~�~��H��[��?�$k�Q,��5l�@֛M�Q��2oh/T������ް�t\��Lq�0i8F�ewo5@���E`�d����W)>X�·+p���f0;�t�ܯ�s�9�<����74�;�h�'FC�l��^����L]�kv�j��㪺G��#w�,Ź�t:��sHn���ۼqʆi�/�� OL)�����kx��^D��,μù|g��9GW5Ӥ�:T 3���ڊ�8�9#��}��p�s��j�.�ᦣ����WY�Ƣc*{�ڣcȐ|A&�������ۨ������<N�xW�c�������/vC��<�����u�+��~��߾�t/�iCu�<��[^@��	*ZP�y|���$�m��x�`�{��W֦m[3����U@�ly�& ^�{���i�*�V_GA�K�WG\��Y5��J�*�S3��eG���@VD��p����L�ut�ʺ�W��o0��t��,ݵ8�e�I�IȚ�n��k�R�wj���wU�>vǮ�N���پ�k�.�Uy��u�^�e��g�Q�9h����x�bg�ܲ3��uv�)�3z�{6{z�zӦ�!ꉧk̝�%oe�͎��R���[����;{9V9�����:�;F��O�?-ޮ�Y��<f�B��,zקh�z�����	�oa�-������WtX���X^K�P�cs&���n��xxx}n��0�����u�}:��f'�پ�,��<�<���\��M�+����m���v���>��9Y�vY�l�����LF�F��m5�;;{�{p`�u�h����'��v�uZ�^Xg53M�x����s�LoMX]�om<�wo*C��T^����O���f���ʡl��"�Ñ�����w^�>8(:�8Tѭ]۝�#���C��o�K�s��ߦ��:5ɂ����V��
��U٭ݺ	,�t�kT�7U��']���n�5�XՏBty��MJ���3��j����8�M�-S��}�2;,Hq�Ԍ��܆c��;��IC�z�φ\lL��t1��}�k7#"�L��S��#xK�,w9��,� �@g��P�T�XKy�{:Z��f��k����O�P���i*��b��j������Rz�q�cU��X6?c��m�OԳp>�t��QS���N���W%h��a��FV��/#.��-��$�s�Z5fG�R�0z�K�
K� N4#t�_@�]']��K^��	ڗTnU��f�m*s�eh�3N�b���M�9��֫�B��(%��8����~۞y�b"��r���������VoCm���D�^e�_�Z���tO:�;�mz����-h�J���[a�{wk6�/kD� r�5��x��q
���:y,I�](��Ǭ˪͗�ч�2��l̻��}v���w�gϦ_R��pZ�gԮ�m�lK�������f�G��\{v�w�.<��ȿ��\�[���Ci�g�.�*��jل$wl�_Skzz�]��W�AԳ���f��b
��շ�{��nKUTm-l��6�[M�K����++����|k�¿W�:oׯ� NF_�����;A����'eBy��c��R�WA�yQ��F�4�&̰D	��e9J߸lհ�Ls)�TDc��Fb>WTۅO�W�`of����9�,ˁ� |���h"ܹ�Mpea#%.�k�T.�c[z�������Ӻ����J0���s�N��$7G����`{��C�}�������:�wY�O�N�D�<�x"��`8@�ڱ�A����>��:��r�א��G4���wf�=k��LI��ڕ;18ዯ-�.��U�������]Ci���r�وwV񩩼�g�<{�\�:��ԩ��s��;z{7�5~����_)wG�����y���� ��0���-��̗���|��.ȧ�&а?*A���&?|�>˝�8�����G4���o|�<c��p�H�E1n�^.�n^�ۚx�{�ڵ���o����9�\ʋ��,�E��|�Y�1��o�^�{��/\�w;ݵ�V���uuz:%o����z��FcX�uR��x�zVΟ�� �۝f�ʂ�_�_��x���-Ɋ��ΩF���F�GNm.i��u���,�q�G���s��^�2�=-� _??�	Y�8\F�y����,��0,+8v�t�X�$r���V^h���8n��܋΃d5of�����צ�)��-ʭ%�5�p'�d�ja��+���O/��ʪ���/!mp�բp@��e��:�J����'�n�܇���U�����:���v?T��ί~C򦻯QN/!f{l�%�r�mc�T@h��م�$�Z5z�4M�+R�+ޟ���vu�zM���$���b�B,Ω"���F�MvnQ�j�&ªt�s���
fa}��`I^,h��D�S)��\;aƩ�;Oo�/*eL1�}�V�ɞW՝ִՅ `�.ܕ2%/¥��|}3.�7�:�PV�y�l[��R�G��v:ȋN�fof�=Ķ������݆�}��L�,1��rՍ���] ���F,T�ZJ��k�������Ѭ�R�k����8X��x�yt>��Y,�ZK�kW����E3�v�H��!d���>�ٗ�۾����d�b��Js��vsdMi����\�ǝ��ح@h��W�1[�� tWq�ϤUh<�a�v},�Y���utN>FM�@��+�;�Nק�= �^O�����!�m􂩔�0rۚ'F#�I���H/F�C�����}�U���i7[�`-���#H�>J��Zگs���נm�Wz|���2�O'y�G�^�E{����?L������Ws��+kI�a\:�T�.7��k��jCg��WF��L0؉�m�kzJ'H��[g�H�ڹ��Ș�C�b���i ެfك��ϼ_�>U�s�����yP|�����6N�vVvV]؂e�ٜ86��m�hh��y`WF����Bq�5l�X{{J�]�S��J����E,5�=�ٽ��Z�y��u���kY p����O���v�w+<���Ϥ�ξ���^v�|�|}��n��)8��s\E_˶�!c��\US=v_�՘��Y �S(�W��i�:�3l�Tg�Q�A�uקʱ��k�u��-�9UTj�u��YQO��q2���Q�]ļ�V+3�?<�+���e��;�@��dg�>�y]������7�4*�Ь�����/6�ܲ+?.�}`W��Oqqz�f�oc�=�"�י�U���mf��/�&9�N�fW�fͿ?�p&*E��$;���S�Bn 5=1�g�V��8�Z�Ӯ�n3I��rD;���FM���%K��5f2ov�+�=eGve*	s��a�����\ɇ��Gs��/2--2�f�#�뙶|Պ=�ܯ�|��	D����5S�����OM��&{g3�{w��W������EBP�}L'߼���w��n�oU�^��	�1D�0m�h�G�`������P�qJ������w��yM��3�R��\2md��;�'��v��d��ve��P� 'Q�6e)]=F�c:��0|z<~�N����,��P����^;4@�V	4#ћݤI�.��#/l�F�"=5(��Y��}y�2#�i��M[{c���5+՛{ �Pq&�U�C��IO.�Lf��@��}����T�3�5�觽�A�AlUǓHg�=},�繟ί�=r�P������������mۺ@���'����������-�M�5����~��Q��h3t�#3v���g�[�K���O�q��Y,_����X��A��'����E��T! O{Rh�z��(������Ӟw�&�{.�v҄a�[^t��V��E�̘�(��&��v�:^�J�$%w8Q��!���j����.�ޅS�2�͜�J=|���<�}�ey�2�"�j.����ݭh�B��ߪy�N���О*���������;��?y�I����%媻zq
j �۸�z2�ȸm
�x]כ��h�/X䄶*�������|:3e�5��@9��ٛ��[����g`���w�wz���j��l�.���6�>b�\��|��r�˸�^���(�Ɍ}kf=.s֯Dy��]��OYʞj���ҁ\��LvTO�{��{��0�@��8�7X��gk[Sm^<8�s�	������k$wP��ڴŕ���y�3n��Bwme�q1�ҹ��EI�n��.�Zf{ھ����cpN�T���w��R�t���W��M��\���I�[����a�=��o9���:�Z�#,>���rw:��Ύ�bn{w3b[�� �(V��p�������Y�_��2kіA�F@���|\���֮1�����6LĜ�9p�r�]˲��i�3d6��[AvϞ�C�}}�I�\�u�H|S�U[s���o�����䁪j+:\\w��k�9���8`�t�^�k�[יQ���\a� )z����sVOp��7�L2�sj=����n�2�|���ڱta�,)�����n��U�m�F�r��*�T2����b����=��o���"K_b�)sUD���w:9�r�^ٳ�����{����xV��`ޓ�b�vi�L0	)��7��l<c�؂��ME\���A[��edטΛZ��=.k�AS�Y�<ؘS��F����ZH�A__u��6Z�-=���A�����}.ENoۂ�"�S��=�x���6�ntZ~WH^@ťR��;sx�B�8WZ�Z���{/�I =ؖ�WJ�����e�]Y�M�YH��\�w�o&:"[�vL[)e��-�H���SXR���v��8d��Qb���� �C�	^;x!�y�+���-R���zQtpd��F�qu�Y��E ��(uvor��3n�2�9�'
��8딭3�(���6L��,to�c���EtwmvͰ�T�;��7L����*�����h���v!��{m���@7��e�ٗE\�Y��C�})��Q�{å6�dtL�������\Xb��qY�	�^�ɩ����3��z��	��v����),�3'[t��M�[��{���4&mM�� rgrsU�Ɨ[�j�����u��])���]>W�ʻJ��̉1���R�c�K/e����fl�I=tN�H��Y�Ot-㷡��l������s�Ԣ��v)}e^�V��{���!��O^0��'6��݂JsS����X�=YD�;[��*5A��;,�fa��!KMh��$�D$z�2��$nN�0n���(oJ�]7u�RLk«
��97:���{|u@E�.r�
�vf���lu�4 ��4@��E�˭�MFV+�y�0��w"]ښ
RGlԭ��'z�ir2�
��5���Zk��\釒��}7z��e�22��4�F��7g/���X�m����kh⽝9MX3g_<q�⧼��*�o+ݚp�6�G����n���~��O�?m��Ջ2�����*�n�ʒ�zںT��	�o{�4G6�(
(E�󎰱ƌ�Z���ɍ=����u�G� �_%��6���p��%�8���a:�&j8���8gP��ku��%n!�t�֓Kj
9$���.�^�Jp�xL�>�j�m��2SXu��9Oh9P��TC��*�`�VbUi��J�fӮ�R�aRTX+����y����I��������i����Zw~a����[����I�P	���U�F��\h&R! ���F�]�irg^��#���q��xō nͺ���p�*��eY�͚S&oLC�W�K{�(��os8U�.m�<�o��Vf.�	G�A,)��^�{9iX��α:6�VCɣ����CN��-s�+w��q���yH���f���@��$ν��2�
ӦD�sH�SuA��e�[5�}y�Az���H�����S�v^a{z��k,�m��X楞z1��E[��|wz^�"MYeZ	0��jl�}����K�\�h��ݱOFU��SƷE��K��ս��.V'�}��V��|t{0�X��0�\(x�	1{��*��U���Ѣ���QW�4x.�9�J��U_�e'�������~��z��������ׯ_�������hf+cA1�j�s��Z��b�y{y?̀�F��������F����9���~?���z=z��ׯ������^�����Q�d�)"*
{����3�D\�T-W"6/q��F����������`��W�t��F�����b�'1�R�9dѰ�A�����!q 9:clj��`����IEEO,lj�����<��`��j����F��kN�&*�ݤ���i���ڂ����Z�LQAM����������o���G�k<�S)Q�(���F*��"�(Ӡ���MG'AO���h��Q��O2�$@Qyjc�E4o���E����r��{�"��̚��{s�"���hѾcIX"��|�E�b��0TLS�M����b�.d��4�Y�˓As(?9y�r��~��������|�]),�I=cs��]��:qΆ�u�*G���Ǻ�����������Z��k0vڔR�iE_����=�h�ޏ�_n﫶�F�Y[2��E`��:W��A��ftc[:���=Q|�Iƭ����u���hGM��,�}F�ݙ/uwzS.��,��e�}{�����dۉ�&�>�ݫ��B���<-���I�f�`�<+c0����<�����1X�O;��<�l-�ؒ���7L�cry���n>SĎ��4�,Y�X;s-gn��}�C���u� �ǝQ[�������)砜ʛy�S��5Ä��P���_|�ط@����:ހ�>��o���'�^�5�Ӝ#8�>��9�]��a���׎��`Wt>���Z�j���U�۵-N���ۮ-�qۂ;�N�����6��_8-�i��S��dQ�ו�6����vG�r�X�s{(�\ǻ��z+�����������
���/��#Ă@39�9]�{v _���T���*��ά<oy�5��v���u'%�خ���y����s�����~N��t�hفBv^�� �m�E&oh�$�ھ�W]WZ&^�i��*��>�롕t�Rܮ���u�:>�8��`vN��%̜�o�͍>��WcKBi��f}�Th��F��<|}�*��w�����wb;�5�:��3W~.�iZ��߻��N�]gU���ݦ�d�7��Td@�¶C��dGY���p��v�
�����ݘ��m�4YV�m�p�|�l���`��am6y�j��5����^�i�{��𱅙󵁾�Y׬՚2ާ��`Q#�>�=Yv�@6�[�l�T5_�(^mFC4��CMZ�.�$�p3���Z]�����J�duŲ��L��J��2*�1\a�T���]�v	���J���֧#Ҫ�����{n]K5T�v�]c�aR!]q�ܲ=\N�x���Wk����o�r�*5�3Df�W�|v
o��{#m�|`�C�o�b���ӈh�lQ2| 9�Nn_F���cn}����h�:lvq�Y���|�#l��Z�-"�c���;|�ٝ�ѽω��[A��j���-�|`�_{ �@_矡9?@i^F[�̰8�o��}9�ٙk} ���ժ��h𭝒{˩h�^l��(A������k���K��T�n��I���;���T�M^�P�kDI�Hۘ�w	�Q�7��>K���I[����a�Ɖs5[�]� ý8����,�C�-�D�L����)$\�}�ն��-�	�kT+z[7{� ���wf+K���>5|XA�0OK�5_S\�nhhDe�����V���d�a�Z�����yS���ww�Y��]3c����	��8#��k�3�甆|����ֻ���1ݴ��l3�v��_iȎ����F��et8U�(V��n1���4�ǘ����'*���b��]=�O1�;tW3�����M�.9B��KɭM2+����g�G���!�%C�L��\���9���Y�`���lrl������]�U�b.c�-�Aa4����0��<��՝L������:ML��n�𗻜�Z���4�ǝdǦy�z����yd��/P�oW� �Z������i�f,����@�L ��b��:��8 G:�->'��论���o/V��A�����S�	����P�_X���t��ES���<�%<�LD����ܰ�;�=Ѣ�`f�x�;�Q���gx�}ĩ��e<�f��������Z�SqW ���Wc��ڷ�+�1س�F�u��Fu��޸�c8�n�i�[�I]�X���;HD�ŧG;/h�vJv],�@���|}�Sy��#vq�r��-{�c�BV�� f��c}�,�/CJȚ'`P�N�+'=�3m��@)�aI��S��Uq�T��H��~E�hV5D=n�x��ϻ\ӛX�2�β�Z�e�>օI-�I^�u����N�H5�p�R�˟�o3t�ܻ�X����U��r� ��۽�}����~�S�ÈD�n~� t��ٵ7��������]��s{��-�\�k
�8p"�bo��ru��C``�[�ؖ�c�^�����2�Z�N�l��x�qV��j�$Y�`SZ���K��[���2R据qP��k��]!���xT������ʧ�νO�d6@�[)�Wl �����D_k��2��[o�:�����j���um��y���}Y�/p\�d�]�㚺k蝥�;�w�A��V���MO���pgz�CzW�W=7t��n���a>7z�40�������Bq?�A2�~�#2�E�q��v�!r{���x���(L�w���zV<t�C'3z�wR����u�$ܷ�p_T��@̛o��ǠNLS}k3�޻�$wm�����]���)Vo�xxy�n�)�lV7�z�s$Q (ת-��9���lL7͋��K�j��g3g�	ݬl�5���7���Sz\�Q39�tuh\����.X�M$47ecާ�|0���Q���=y�	 �;4��0����t�|�q�KMun�E��[r+�t@���KR2��5C��x`�f���S������`�Pb�_�穄��oes�`�S���Ҿ�Vc'����,^��%Kkt�a�	�ތ�Z�]��^[�jފL&�Wo��o�u�ۡA��ݬ����ٖ�x��tE%`/N:���^%�}j�i��\<=>V辛�N�iF3��жFuNzz�K�q=���5��Ś�8A�}��;2nzڛ�ن��(]e�dp[���=��o8�͢��������"7sq�>6^��7��S�+3y��6�\i�R��h�wkQBe���y��^{�Y�3sۖ&�l��۞B-u�0
�����r;�7��3PDg����n��|�L4?[����� ��뿒�&g�^|D�����x;��f0�[��u��������kWX�Y��3���Q�u܀�	�y5R����}3w�/����KUe�}�B���#�>�9����a�ぼys���|����x3�V�Cg�����ݻ�ʳ�������=я�-�����9T�ϻVyK[�-7�ә��&N�9h�� ic��:n���8;�rsT��]����!���o.���́[�5��>ְ�5�X.ܾ}&�����|JC6.
C��N�>���\��i3.��yՀE�z��|�ۇ��ͽ��.���Y��|�pP���n���ώ�v��<N̊��d��'�3G�Ä<�q��$-�.5Kl�ں�v8������ۧA�M,���4u�����y�V;�*E���V����4�ZɾU}�U�{.:�;(��0{<�l!U_.����R��r��벺z�����L�ֺ����f���q^�m`Dӆ�P�0�+~#o *���%��S	�ޑ�����R?�.���$�o[���3w[�+W>�fQҨ*���:�5(0��1S�c�E��r6��$�m�E�y��gA�0{��U��;�e�ۗ}�\��`�9ߧm�1Q��9���̒�i�WÎC�ۏ�C�[���ʝe>W�m��l��W����ck�*4�,�^���ͳS����mU<4̥� ޼W���S�mvamP��Ŝ��+��m��5٫g���e�kˆ�PG�B����m����'���C���Z'Utm��\��]Աֳ���-��lY�R���樆��2yr�3?R+*����/��g��f�n��k���������78K<���PY�{7Ktͻ�57��JN.��y�D�5�b�K�2�	���p]6=��e�@[sK��v�6���m�wO��[�ܫ@妣ʌ8[cZ�s��M����̉�ێ�u��A�����.!����2�*+�Ԏgvp޺�ȻQz���l���<m����!�-3Z>�,0l���WE
�������B���o�q�8�H�,��h�pSj��\����sHl&�����\̯�;z�ܩ�j��w9�N��d�il�������A��GT��vl�,$n�Qͻ��M�em2��X�%VU���m��R���饻�ѐ��(^줕���4pӘq_�Rㆠב
�P�6���#�K��4�6�b�AIR�|�]����
�;�Ic��O\�&�*7� ���:=��fu��y�z���S�������r0Q�����M]���9�5r�lɋ���!y��.w�μ2��}�'N��śx�,�O�kˀ�=U]ү��i��;R��+��VY�/�$4�7�v��녁�[c߀*��-f���Z��>����TӷS�~�wj���H�����l��Xύt�M_@O�+�a
�1�{lSk���2R��-�r}����\�"rg���c<��S$5�L{R��<���R��f���^0Bh����Ó%+5r������oT��~C�>Y+��?�`��p��UiH� $Nv+��Y�p�nkd�V�zW���e�5jc�e����02��7�z7�/@���q����MG�O�,�7V7�d������
A�ksve�7s���9�a߶ݲ%=�ʉ�L�-�Bii��}}�w���$����0-ɤ���ߏQ��J�J#]O�1z��27i]f&��X���[ffn�vg3:�e	�N!�x�tk�V����=��fQ�n��"w���j+���X ��b����Avfv5[��i�zop�b�ų&�:M�,39J��8[���9,@�GΕ�HU���ƺ�1�����l����S�i�~z�9k���o����� f�<�m)u�>ۍ��Ԗ >:�쨥� 5�_�j��T�f�׳g<_f=lE�>k�GtG%Y|�?\�!�P�t��ϯ��ݴh�y�oZCt{\�C=ݒ�e�c�S����[Pw��l?���r��������z=�,��wg�E�V�(�__v�褘h�߼V/�w�vw�Χ�Câ��$(Fsf�W��ǥ�y���w%uKT&��=���z�/V]]��c�n�s��Q���xk�[u��4�6�����7����\fA���y��Ψ^��Vz-\��4����p���5H�>�s�\�{�m�؊��pzF��̅f邹�۪��g˞	����ۑ�\;��/+����Ee�J�E3;GFJ�&�gܧ|A������gK��oyr���
n�f�����n�Ʋ��Q����:�q]S$Ͷ3%._]�⚈ϲ��5��
��·!���X��0�G�F�j� {��V�=\�` =�żVv��ض��"f:%���b���{�J���!�`gj�'0���B�W�)��FT
��^>>������؍ǜ^m��z��Wo�R�=��:�X����P}��x�������>��n�P~��}b����|uz�Z/0�'Ô��כB�#^0��Ln&��Y�-Sr����!��S�J/o4uǽ���f]�r�c61b[^�ڜ+2}��X��6��z}1xΖf�|. ޅ�x���OFda��}�%7u>ݟl{���� �~87ǖP��t'l��rs����t�~�d�<w�v�wq�j��:1������yo'a~�����4h��>A�j6�>~}����w�s��x�܃��%J�cx�uO���vp̫��k�|��`��<��é�	��.썏@���<��՛'��H���M����1S'bt�|[>��,G�o��u[Z�X��:=���y���%��MycX��oLx�î��w�o.�Ξg�K�ۯ�N��xv�>���_����J�W>hR��o�}�)D�ZC������:뫷;�NZ�X:�-#-C-U���H�Ue���2ʱb2�Yd2��!��,�2ʲ�b�Yjj��eYb2�YeYej�Z�YVZ�Y�d2���Z�C,�Z�,�VZ�,FZ�VYV-#,�VY�2�2��!���Ub�2ʲ�2�Yh2�2�2�e�e�b��A���-#-U���!���C�-C,�ZFY��j`e�Ťe����!�����-U���(�۲�Gp2ʲ�Y`e��Ue����A�,�Z�-U�����Ue��A��-U�Aݸ�VX����j��jd2�X�jeY`e�e���e���,�,���VY�.�,028��� ���e�e��%�X��Yh��e�b��E�K,VZ,�Yh�Ҳ�e��%���Z,�������e��RŒ�IYh9.@2�Z� e�i- @@��<Hi, �HjA��5����0��i�@&& �Dj��kJ�Dk-d��5�FYDkk:t]Y�Uh֕�Z֪��Z���Z�֤�Rkk$�+�ijL����id0¼d3 ��7��<���Ue��!���Ue��C,�Z��.Ue��C-U���P�!�U�C-C�ݳ�c�~8��DUm)JMi*�f>~<����w��������_߿�t~��{?��:��:>S���׻Ϸ����U*��������HU+�����fj���'C�>:�)�פ}�UJ�����+����a����~G�O�Ϗ�|�n�o[(�A)m[
e14_�+���f�4��Ѫ������+H� 02�2��2��j������d5LV����U�!��U���U�CF���I���3q|_��?4)R�B��6 �B�k�s���OG��y}~Ӹ���>O��J�W������z}��u�ޟwi���s>����2UJ�X�3��t���*�W��R��=̿��P�W>�޺v�5Ī�]�^�|���/��w�yu:?��ô�WG]y��p�:�U*����}��UJ��|�v����O��������a������\�U*��?����UJ��c�ߣ��{�����xO�����"�����i���%T���k���>��{{���=��{'��y��W�{W[>��q
�|�s������?���O�1AY&SYZ��KY�`P��3'� bE��ZT�FƈkEkPUPI�@J����ePP5�6��-e*AR�Mj@U*�@���̪�m�QU�T�h�����֦ՋZ��L�m�MJV���ŖIKF6�����̶T���l��ʕhٗ���b��S��܄�6��"�ٶ�T�)��Z�e�ûZ���2b���[&3cTm4j�Z�j��U4�V٭��ݵ�J��bY���զ���kVЭ�V��[m�d��l��m*U�V�P�0�k�w�v�MkI����  �|���5�]p�j�U�˧>�Tv���Κ�Q{u��{�����7�tk9Å.��z�x�^�/fح��s* Z�v7Cm��[�2͛m���-����/�  ;}��    �>>���
 
>��Р (P
z{��� ���\��ݠ)g��JҦ�k�޵J
w{��S��޻�x��R�Յە�T����KfkZ�65UU���em��  ;yMiG�����E����G��4�h�y���QmMz�`�o+�5oF궦����\�: {u�Ү�Q��[�s�Ym�n�p�����[����M���H�V�� ���W�JU)��mP�Ύ�C�Dy�[{6�y�'�
{h��0� 7�� z�W�ƕ@=�gh	*s��p �I]���U�����-��l��  N�R��Ӿ�R*�G�5AU9:��ޏ.cU8�M��ypR���v;ʭ�A)W2�4�mJזF���2ڍ�f����Mm�2Vm�  ��}�K�<�t�c��9%�4�g�Uu[X����2�m�A��tq��oU(J�Oq���:!����=��\:� ��͵[6�V�5�43
��   1��h�ՎB��׮#�@�` )EMX  	�ˀ:P��T���� s��  v�� ��q�LړZ�m�m
��   <  	��h  ;��  ,�p@c�� k�p�)�  m:\h�Lw  ��  ��Y�M��������kL�_   π �p@�ε  �n  7[n�  NX  ֠�� �î� ���4թV  ij�Y�Ɍ�ֶV�bٵ���o   �<��i����  ^���  ��  ��  eOq�� g.�  ;�N  ��� t���  | �~@e)J�  "�ф���� ��x�<��Q��"��	J� d ��ѥU&�0@&�@ʢ��F ���������&�_��M�:t��bU�ص\��u~g�޺�&��=u��뼝�d BN�7~�r!	'pI$$?��BI�H@�$��H���	$�����'�_����W�-|ofa4ap(6k&;!�kZN�(�r᭥zQs(Â��OwX�)b�y�����葳�&QF�[ݬ93b����⸵�5��(��N�f��I��[��Ne��[�5m�̠b3�;�a8�LfLEQx/23QK2�Lh-��*�oN�BS+j���+e;�K��k�B�IboF��{��#0�{]ݧ���ya�44�!yVk9/��Ws�ǥe� F�AtS���峳
7
�Zp���	�,�I^'ES��Z�j*�E�e��Zn��s2Lv0%,
�1��;����E5�h���u�r���:T���@Ӑ81f�t΍�Մկ���Ã
�H݅Cf	3^�Qqd�w3�䵥��fhZ���=���$7+$'pn�wx���+X�%�Y:֭�cW�D�:[�wov��������h�XB�fܣ���S��AQL�2,�Da��� �2m��j���ɮS��-*VE�1��^�� �ť1���w(S��U�˕j�p%o5)�6�z��l�d��Z`+0=wQ�V7�XKZ�u�5`���_H�6�/�}ﷆ��V���P	]0Y�n�E�<Qk��E/30��cfG��4b��E���ӕ�0=q��C2(;��ж��ɔ�x-��5��.�;�o��C¶E�\'h�k�3V�$�m=tl�U��E�0�/v\	Ǜ�"�:��-B\�q�9�M6������J*�H����Ty�h�V�N���餶ͨO����0����1,Ù�f����cI��u�	րjQ��Ob�^�[u��h���i���c�� ���4���~L$^=4x��k�{���)�Ŵ��YS\ة�W5�X·{�����m��p�f�V� q�h6���n�ب�kY�0c����n����І�E�IM�+9��ű@Pc��r�̺!�����z�)%��!�Am*߭U�W)�BZ/g�*V��7�3p�@ $
8��j᏷���a���Q�����;y+�4\��L�6|A73���7u��A+u��9��PB6�7]� ����%@.����Gו�F9��S��b����{e�ѭВZ+2��el1	BR�e,qf�8�<�����e��{��:yt�
��״駤f�4yu��=��B�@j�	e�.
ڈ�r��,]c�q��{a�&ˎ Ȥůp�Ã���$�6d�yNP*�A�:Ԁ�OAx.��|ӎ=���q��B�nBJ��n���?��y��FI�lm��C����Z˃.�J�`P:�N�XYVؓ��5F��Ƥ��	�>��i�0�N�Y[fH��L��Z�܉�m���©<��v5�imC��ƴ�b�`�r*WH�̊-T�˕������U�U�\̃K���C� f�j^*�XՁ�U�
U�"u�.�;!E���ܥ��������ocћ���ĳ���v��%�<$G3�哽,\�ݷVQ)gٌ�գQx\)F�jT��')��ź5�oPxCy��Y/X/@ϖ[�b�^:8��X�U���Q�Y����ջ(&�;h�4Y�J�ܫ&�O,m֭-�+g�����i����Kt�̙i�n�_�Hc �Y�����'�]�{�f��d	��؄��-���V��U�'��[yZ�f��f�iF��=�XT�4Y�!mkJ �R�e�nb���YB
Б"�Z/X��4, ��c�����V�&�"��l���X2ԫz�i�KwH�oe5y@'>5v��&�1!0<�b���A��Z̦`��=X�m�`1"[+�E��,�P͑���yj(
����u�0�1}%d�xԺ
�&E؊�����"o2Y)[X��*ޯ��F8�V=�#��aE(�B2j��R4CShZ�p�N��x���IC��M]%�"CN]�4f�ɭ�fb��V���Ub�[�f}l`�A�ו����%Kͬ�,�"��5b2��V� ǚ�YT�W�F`dK��m�p��_�Z>x3�Uګ�{w,�=�Uf�G�kV�FM���u�E}���3綆؃v����T�H���ܣ�-�wW�q:��e��m#��-mǗ-�
d?�4ZjM��Qa��.�-9k%�5z�mbɖ�������s$��[I��u#*P��NJN�/%�KR�w��hl�b��Ay��[GF�ߍ����S��>c2�&��ĳ[�QT-903�茲m	��`Ǐ��ģRAh�n&&���7 ߡX/	�{�	�޳���0U�!���7BTj۬O/䮳,$��@k5�ٷZ����f�1G>(uaKl@��ۄ<Hj���t����[��5�	5�÷��ti^�=�w4c�U�U�*
���1=(P%��]J�6�vg���"��n�I���*�a,�V)2.L����4;��xl�R��%:v�\�����J��Y��@^)�\�0m��Ah��ZMX0+Z��@���e:�[��	����27�:�Jc�x��Ve2<����@EN`�v��m$=X�a�fnͣtw-�7v��� ���է�5L&R:�@�Y��e��<. n�Cq:��^C%�w�a��YM�Ø�ԭf&��:��5^�����-K`��י�odt��9�j�;9��^��e��:�5��k7���r�Y��]<׌XJ��Vje�b72/��T�%7h��V hf5ab����v�C�	�G��Ɇ 3`w`�")X��}��r,�Z�����6���)q����t����ūa8v��-'��j\�����s;�@s
��6hH�qiYB%qaú�^�5�q��<hQCgȩ�J.F�@q�%<�4�-K��k��"G��{a�B"9�N{��,<�q]���EKE,r��Wm��Nղ�Yy�1"A1��ff��h�:�KLh��j(B��6�y��v�A���'ԕ���35̰�Pݼq\`��XV��K�\%Y(+9��MԹbd/�v=���6�'�F�ks��Tᖢ��u��SZE�.;��e�2��3bMVD6|����C*�@2l��i��/h��J��=����k�f�6�ͱt�w����at�[�Q%��ǆ���A��]�)�
(�A,i���(���؈��J��4�XՑ�)]��2vi	#-���cmGH��8)UЗ�P�G4�U�yDDA�wM��X��� Z���a�tP�/1^ފӓ	�#� ]���-��;�m�A�����t��i��lc/.�j�^�ɓ'o�p�D���^���b ��dm+n�ǎY��ۤ�K@GuA/��n��V�3F��ò�b`�@�j��n<�ɤ/�{��f�cn%3v��J�ā���aR��Z"փ
��5�ǴH3,;��:j�]�S�r��k0hX�޻ȵ�)M�rZ7��2�E�d�����m�d����*��RA��L�N�Hg
Wp�=�������#�l0�/x��$
|�/��SH��Xp%��0���ܧ����t�^ŷQ]�	�ۭ����e��jm	�Ͷ����$��e��J��`��}���0p3��OsTڷ32�h�Z6�
��T�#k^`�`:�1��^7��ݲ�⦅6%^�2�V�ҭ5i�2)���6��FV
Tė���K��M��v��B�XD빴�T�Md�]�����D�	3A1�&�\�n�1��i9���K���nb$V�xK.��F�g+i�GKU6�*ژ�ڵ%3)�+${y�=h���.����.m-j��m��D�"Gwr̖�j�C7�T2��F�0l��Fbr̥��2�ZKV��&b��_Z��J-&�Ҩ�Ǌn�n-
Hh�/0抸�BR	�2�-��l[���.ef9u��VZ/��=�S*ނ��R�3Fz=����@�����2^b}������MPR�=��aP��wYnPf�)"Tܵvd�Jѹ-��D�rδ�)�V��zU��� ��e�hX����i۳�&���ut��ap#�Vq�̡KjŸ	;1�dCEG.�Me%ml��I��LN����)��%�#�B���z�&U����i�Xؠ����u��<0�XU�\F2��e[�Rb���y�蹮ͬ׫ �PL���'�����
�X�JM9��p���^�ni�r��p��A[ۥ�SIԂKz١w���XX�̥IDkVH)���ԛ���f��M4�ٰMp n���u��ST��J�-�n=r�sNʻ�4ʫ� ���3�� 4-4�՝�0��P�Q1XL��G��pLW5KՊ�̖�[Bi�@ʓ`�_�h'�p����F�[�R˽�����I��w�n��
�B%����Jh�1[X5-d�iP���yEX��ʭʖrCc.��P��J���������^�m�Q��I�sCdT����oc�,�[jܹHf0
�I�2�ɲHYDZ�`b0p�xv��z�RĶ�c��fe9�6yÒɅ%�V��A�)C��CՅbX2��]L�5��ܓ[em���KPsWآ�(2�v��j�6�x�^��N-i�W��&橙ʻ�;h�ah;��p�u�N�ң���	�X��*Vwl�M�t� ѱ������1�NXh�����s]LA<�*��hH��ڸs[*���ύn���ݎ��lMx����[w�p*XX&��X&y2��*q�Gu�l����q�����Y7DEP�t��Y�8S�Hj�>�����^�J��'��w�-˧�k)	�R���@�B�GM1��f��1AN���f���4�Z/$l���{Fт��cv92�XG �А�n��������x��{��R�^=Ge�������O�"6��pm�e�W���X�v�2�1����u�k啷:q-��7PG) ��藲􌿁�{SJݻDK��Z��E�5��n�e��vKRrbw���H�Z���4!*՝��m��)S��ɶ.�͇H��f��hF[�B'��ia�`�, a��� Ш�&ƙG5�S��`;[@��������2aRbut�ⱊ��zo�ؒ��-yvs`�j��r�^6�˦�(�t�<��/J��K'P��Y����k��R�c/*�	���w�`LЫ�)�CtCQ(vcZ�M��J;T��sf�P6؏1�8'hc*ي����PcV�;u7V�MeҊ�[Ak���o("��$43� ��Vݙ@溆(c���^���`�Ђ�l����p]���ܠ2���V�E���%P�z ��ݦF!�d,��-U%�ж 6 �*�ah���XԳ,��QG ���-i��:�K�z�kwu�-��,[���*�S$�s��Z�Yɴ��{z�vi��6<Yj[M�Y���D�6���-������A��A���7PI�\܎4�L̵�B����wM��^C�#�
2�o~4(��j��a����k5	�(L�T	�,C�YI����z�P
����+�t�S5yP��<�.R�ӌe�6�A�C�x4&���[�;�)���R*�+y���Y�  lx@"��V&�K(���+#�m7�XnV���/sV�Av��Vbv�����V��t�8��C�7N����e93~�bj�V��6:u��N��WoLp�i��ܹ>pAWI�y�V�#�8J*Pߕ�؝8��enZ�A-.�Xi-Y��Yբh.-�Sl�u�)�3(Թ005)	}�5�'�lcGqn�hV@�����@
���ɻ�+a��F�����Y,fS��O4�+:������mH�0EyK�T�[�n�-f�)��ÊZ¯\�7sxl~~^d���$�#!�7{��\�+h���l�n�D�r��% �)�;a����
�;��&��Yrń�����
�%%n�^���c��B�^�u���&�à���I��J�F���;�J�Q����!mπ↱v#�����*!b��n���|��5�-�ò�-���?Lb�U�7k���i�Z�Fc���4~��๏#;��������xޓ�2c�Xͅ4|��ٙl��
TX���������Q6���5���3h�5ـ������ Ձ'D�)<c+o͕�yiPV���et��4d0A�r>]�l��3kF��f�h )K�.c�*�7�/�3��
C7��t����Ú�jh�S�Z�	��T72R1"�0Hn�̄�y�a|��gY�����2 ^,tt����3Y���6e)*��W���t�d����4i8DR��"t:ņ�T�)SQڧ�S;Xv�2�H���>��Ru/k]m�ڍ$�3t���y��kU�mg�,,ܧ@L��I[�C��Aa�
��j��L,b̛Z��Ö�d��xFI�m\k	t君���_QE�܇���)0s�
Ƣ̬���
oi���VY{m��j!��[X�՘��m|��$α��V(�W6�d��mJ��͉X�9��Kh����V�֍��0V��-1]��	��h$B2��f뽬C~8v�Z2�Da�W�wuQ�rncsN��W�p(]�q��J�I���[�h�ř��a��	ݨ�"P.��Xe�6�SH�X7`XQt�4�.������̷Xݫ�XO��)�9�,�]iW�á9zs�N=Z�'�[�Ņ��QG�u���C�C������&,�"8�z�3�����0���$C�
f�R��G��e���gH�wd�����5D	z���e�m��%V�����ЩJ�m&Ekܚ�/�z�%i1�@��iҵ1eM9yb�o5`;�[�k��	�G�f�v�ʼ�۳�v�K�N�ص�<�M��:��^�=E��!�_�F�r�c��ezHu�T�-nq9I���� ��m<�6��B���K��q��=|OC��-���G��9{f}�k��v^�8�m���YN�����"�[�w��v۬�yR�O9깼�qp\:mv�T3����LJ�C�ξ�:^�+zx�K�A9�b�潤0������Tm1��8�m^CS��7Mc���Kb�u�k�ӌ"�)�����i_oYv[�q��e�>�`��]�ܕ��n��@0�����$�kt�&k�H���z7�z�g�
���c-���NcX�ٜ3n�uvE&�����v������շa���,B���ǣ��b��&Ų�s�\��Xp�6S޼�N}�ҩt��֙���i����]�Z���@oU]/�n�rH,2�G��"Јڈ&a����`kĮβ���7d�b�_m�;�d�|M!U}j����ö(�K-%��5֊�$&����Y����-&�K`�c|��c��R�}�
�3��Ђ�tf������1wp�+]o[Y!~�D����\�rd�Gw&M�gl��Z\*�-��!ģ����luYx-�c$�-�<'o�fsó/�,��2�'қ�(����^2�p�,�G/�XPV���YW�.�T������Z��� )��p���>�����b|���^Q�w�{2>��ty�+]�EL�	��:�4��dX�D�̅��r���b�<ˍ�x���^̇�.t��H��f����m��Z;$z$g���1Lz�� �0���b�����mqM�y���*�Ւ��U�=�:���y�<V�5�-rT�����Y�Y]��s
�Zw�Ћ�U�[�˛�b�Z�I�j2�o9ǰD��χ
��`4Ĳ�!����_!�<���=j�x�H��.�W��S���1�s����<h�w=�RT�"uw���{�w:������y����=7��`YW�v[k��{��h��>tt�-0F,W�/�X� ��g���a:�
uXϧGc�-�!��m���p-5�}�pY���p\�Ȯ�N���.a-m��z��c�*K⍧���w�J��KF	3�$���4;/o(�t׻�+|����z�ˣ��*H=�\���d+��Wï���y����hb��Xҩ�[G/^��=݉�X|�X�oa��ҫ���1��%�����G���;��{)����w+)��W1���S����[�i1��<���2�w��1�������p�fT�E�L���^0kX��ͽ7��[B���k���%P�V�'G2����a�oD�evb���O;��o��S2�Ϯ���},^ktgE��+�#,T}a�6	|�P�8�-Wd�������<�`���|�N�3�C�~A�0�k���pm�Cf�%�7�Zr�4�j�^��ޙ��,dγ�����Tt��0u��z�=�BE�y�}��e��4���깫��˳��
�8&ξV����/�R�X&�8�oIm����1hp�R;ժ���p6s�������v%u�B�&1�����ͧYG��,�zK{2.$�^d��Y(<��z=&�>��e2cpN}q�����{˳i��zx�GGpه�l"���gv�+1�㜎��nmf:6>�ڽ�l����gJ���s�	�j7�+m�`�n�,�᫾R���o2���]Ek�(n�wrCk`f��Z�a.J��m� ����ib�Ձy}�y��3&�o(@�-W��̣F�@�Cv�W��ާ��Z�V���&`�wC���m^
���E�p$M�����2�)`7�%Z��K.�ڶ���1o,�/5<1k�*�]�6�e��MJ��5dAz�b{Us�uP�i�X���T�I`����C��;��]3��:�ёy�8�E�CWS]�ix4L��u(��G�q�c9�FuL�o0�W���Ҭ����\|*	(c 8_Ji���[ʵ[b�
��0뱴B�2Is�� q�I}��{��������
\@y�y�]ȫ�z�E��w�We��[�#����z�I|�!W���q0U'��,�r���G��Io�J]�O��f��+ܭD����oӊm�ƨĻ."�6Qt=����{Q]<�����P��g��b�80��	�$ulMZ���R �|��x���%��10Z+r^fB�kh}�Z���7��EБq&�%���a@��XL�6��*����hq���
��̉[�"%�M�Ood�s��'*#��<M��%�.t�^��Ex=�D	�Jh�n����>Rʍ�u��I�1	���C4�Z�y���OqJ%�sIJ�[�-˗R��Ky���ݬU�vS�u�8K�D�}d�Ka�̼����V�}Ԫ��[��̹�_�gM�	�#�=e�@��]��圗�1(�w�4��es�Ķb\�'Vz=��`��T�'R�s0�#BK˼�t��Y)��=��������hu��[M	ղ˼�l]�PI3˱x!w�*�#nʛ�M�W�`#yKn��o�6��A����.8�ɯvK�H�*�W���p9����f��j��[��ζ��lC�Q��I��a���b��`V��,<�d�G.���n�n��tη�p���!F���RCWg��Ԭ3k�k�7�C)�mL"�E�ʀ]�͆�k�pve\l[��ƞC�k#�Sl����*i���֒3������qt��`�ꆹ�Ʒ��b-M�����T����%IZ����=����Q�}X&����K��̌[5
�͸U7���N;7A�̑�B����Ltu|nJ��d��ݎ�z.ʽ�@����<䘟\h����y��]ar<6���]�rS
�l�6����n{�1��v��J��\xy��`-�g2�C�/%�?`T�s3~9Zxq+���x��tk~���aJ���(��
rs�c��t������mjա���P�؟}�q�3{��v��n���د���R�2ɝ/��f��OU�0�h�U-x�����hk��֊�os�&�/�bv��iRK9Ӿ��Lc���b�%�*��a$ʟ7�j�ci�\Dݭ�j�i����X|sܴ��m˔m��+W{�����#�dcU�_9��l����+"p�Ⱦ8c�6��&"���Ki[ʊ�J���̌Z�8�!m�n�pdGu������|�h� hi���at�x���,b{�Oc��b�'H3YQN����(E�Ռ�����//���9�x�튦=F���L��}Gx̽��޸־q��󉌎˔����,�
�Jfd�2�<BŲ�r9=��~�󖐧a+}gU���c�Y܋�jSg��EGqҤ��xM���wA�lc/33lǎEWbi|��-6�[\���Z`t�f6���!i�-��ޝa�^Jk�e�M��]��D�DX�#3\��#����@����%��ר^hy�+8nR�P7e�tݴ�0a�Kc��uYvΪ���$'�Z�.}";H7�"���8Qz�_U��w��G)[g,e!Y��]��;�7:P��y�15X�`�^Ĕ�a̩�.x�/��G�K������{�N�S���Tej���� ���\ci�26�$��Q5��V��s�܇n�7{eB8]��k�
��M rd'�<t3��)���^v�T�X��a��{����Ѝ{�%�'}��T�TH<��Zk�i��8�Uֺxy�� c,�CTGtո8��h���"l�. ֆ��\�=tc�|d3���;�nfk�7��$}i�ţ��{��r>�[Ckrn��l]�2R-�4e�f����Rv������C�9�r�{K�����@�� #��s��W���7t��ua,�����^I�|�׆CT^���;�
��}tl��I� zd���ه�I�w	�����Y��Lh`�m�g���$kz.�O��z�d�H}�G�>si�<�T�w07��t-rH7�%�z�����n���p���4%��1�+y�ݲI��K��v��뫜���6�%���n:��f0v��� ���U�/B��%��_n�c�}��x�+S&\/�<�Lxߟc��S���dSg�)�p�뜜bN�^��R�c�ݒ��;A��|�N�Xj�f!���/�ie�э���V!�������d�|Hj�U�.��˝�e�]m|�9��8��뻒����Z�Q�u��vV���KUO�X3�u���V��k"O1�� ���YX��A�9�9��R	�T^��T�bZ����^qaYvuǞX��.̅�.v.T7d�z�gV�ˮ��K����&-ч򚚦�ł�3�KiWNe5���q�r�bg�`+h*���e�������ػs!�
]�m1m�QN�IPޛ�l�����R��$�[����S��x���}�.�P�&������/�(+���4�M��Tji�JeJ��vng.���Mn*EG=�Y���y��+a��K��s8)r6^E�(E�p�I��P�
+2�I�'	��=*c��%���
�9�YN7&�4�S�֤��n����jz���1�k4�²@�'��ɖ��Y�+Ɂ���:E`�����#�IN�p�)�Ș�y[s�\:}�U�-��s˦��D�ǟjvOF��˵Z�x_����haD!��-+Vb�<���^��}θ�&}�wU�kS���`�*��&G7�Ȋ�[�����X�s�m��+r��K�{A���n&�|����/�MU�i��]h��G��i��z�95���[���)te��Qӽ!l�F�wc��
����8�g�>3駛ů�ؕ[��9R�����J�={�ѕ}�3G;�(���_K�	O1p�}}D���.��`�����]��%����m��ξ����,��'W� �w1P�����1�V6���U&��ع�]�;�:NX�y.��4�t7[ѧ��W�l�
�xw3�`�-�ǭU�$]�i]�+�N�9���S��u����x��g����H�
a�-�4o�(?",���;z���<�>�x!˻��嬕{O8M=�v��m!��YVeuH{]�f�w�R�Gs z��i�f֝�D�9����n�ɛ�F���'բp��ͦd���n͜�E*yk�4_S��b�p1��v�S�u��4���G�Yګi@�0N([]k��{��c�de�eӤEt�����pV*��!��-[ޛz����6�;�+�M��)�(��&ͭ|����,&S]x�
�䗊��d:`WQj{���	�<��Sc�FD���z˺�$-�A���H �&��+:�0{k��^̫�Y�D�Ѿo�"���o�o>�ŢV/KD��iM#޻xp8��F`��r|���DE��\X�K�µ
8�����fh�ξ<�TPT�_=r���ڜ��cCxm�t{X�gY�8NۣS�|^_+/�gKŊ�î���9�tC��c4R�];��k���1�;) �`B>��늰-���w�g���:<��`ܲNSٞZ�
�X�� c�9�nq��r2����,��_M�6�nr�����י��Y���M*O�r��X'^c�����fF.�/v3�n�PTeT1��[/mgLn�f�$Te��IqYV�*C�R�_� �D�=ǈ��$2����%�-��f������w�F�<����<$�M�Fh*Wv豔,,}��'(��<�ri;����̥�k��3��9wկ����p�C(��w2�n��z�N����v;#��v����`tu�P�kjƚv�W�"��C"�r\�(>�v����5o�����$3�qW:N�Rq�qb��
�|y�ͽ��u��j�7�J�F�H�`�B�Jo4��̫)���߅,QiB�צnC�d3�I1d�$�A��5|��a��B.VQ�m�{X�W�Q��j���{g)��* ���zOv���݋����h*����-��w(�}��T��bU.w΅����˽��s.��%e?R��`%B�]˗����V���Jz�"���[��%�7F��) �W���'��j.����/�m�Y&]9n�^�.�6PM��F���P�<�[���%@�K0�R�I`*Z���ķ��V����ꮀ�(�7,�56�=|�KS �*K��������Z�
R����y�t֩��m�ƅl���2���Km�8c���A\�#n'Rkp�]g�4%�|�B�)��XUQ�b�Q�xұ�&3�b���c.�
�V�����!�f�NĦ������8	5K��H[5q>�&���w�Wz���g,�0���Ӟ�d���(��c��4�e��|�21��(�Y�ucR��dG�}�ʃ���myn(N�f��-�鷭���!ΣW�c;�'�jΫ7x�%b.
��lod�{���#x�{"�]�����`_b9݀�YM�g��t�5�vd�қ�&<*�	���F��짮|�V\h�U��.v�f]��@F���hk���}:(�F��ͬxpU3|���������{�(3#��,^�K��j,�3k�J��o�r�����E��7�� ����{	����P�a��^�J2:D�4�y�������µу��cymZ�����}��RH}ق??=��7����uF�^a�=׌8���nf��X����kn�J1�@� ��/k=�0A_:��p^��lUoS�>>�ێƣ|jى�J aF�K�����v��4���X�Y�����u�آ͘�=p�Νܮ�⏻����(�(���cD0i��Dz�*2�s�8�������ʪ�_Ur���>���}����I=��:����\�f���owO`?���m��:'����ZA�����m�*h�i��EeqUh��T�l��5gG���.
��;7��xU�׭�5(��P��i�&d���	5�Qֱ�0c���o�/ �B]Oc���5v��ԍЮ��;>k�NIS�u�����+���Y�f�ue�т(���4zy ��+��Һޜ��D,Nlԭs9�
-;�HM7m\����!��t��j��X������|��vkd��Xs�z�&r�4����Wh赜±�%���/kY�69�g-��
,u��cT�޻��6ꝺ�Ϲ��O*��;�w�O7@HʆI`+'S�NH­ Z��\_	�X-���ha�{z-n������ى68�|6g�۬�Z�q�c#�^-ۅGk�
N�>��}&�X�;�����"��P��7{��Z��7St[�ha�o���(h��ס�J��=$fcw�_8�D�-\t�qw��\���S�3�؃2,*F��F�p�ީ�Mu��pv�6�`�;��L��k�cf���et��ͶCX��H>ҽ�h��aEh���r1X�ln�-M��X ���=�I�ҙ�y�C�M+�v!qrT�g\����N�Y��Zʆ�+��\�w.@#̸�w��y���uqÝ&4Ⱦ���jV��rE��2f2��R-���C8�3.}�Ѭ��sx�ݽʋ�j��e&�V�Νn�����ၐEa:˽TU«���g�Qޡ�콝'M�����e�Ξnv���a���M1p�7��h4�����6��o��L~���mC���(��^�Rt܈{ԇ����� ]4��ve[��u�1en�o�o�h�&Xo��A���Ļ%��B���7��]��q*���g��JB���������L�9�Ȅ�ۤ@g0�t���{�8���KnF ʳO��Xy.��y{H�ʺH�%Y����fƍ'f��Q��<N�w��8/��hX",�����*��oI�^��u���w�5��i�3�Wg%
	�F����yhL�Ӿ�&_Ɠ�z ��n�ּ\_M3r5�	��,�Ǩ༮C��`Sͦ. ��|<Ts��3${q�Kݬr�٫�x�;��iYQG��H���o{:�v1�v��/0�b�K�9mB,�|j�5p����������iA���������f,ՇM��I.�J�g�W�6�����#����N��p�Ƿr�SW��3`�+���i�l5�Һ���NȮ����:��`�]V�E�#|�(i�/;�w��͒��իW�JvV��z�!���1�كnªG���N�9��ىQ��LԼ�^k�Q�#��0c��س���;3.P���t�Ӄ4��Bv���=o�".�krX�t7u9�aQE2�U�9zS�W����B=�@����7 �pɍ=�b�Xl��n�b�YB�l��ͨ��W�O����'+��g(�T�V��YWύwF{�[�
L�?V�	��X�K��k��V�o:��:	���Nl�����C�D��<�cy���΀�W.�kF������ΑV蜲�k�����T}Տ�w�q�m�_δ/1)ssU�₷p./�'�g��
4�S�����Rѥ��]MH^F@�٬v���j�$1W�#�ñ�6�E,͡�vx�N�[�E&s�:�[z�#X�Εu����C��+�� ���Z㝟$������J���]1�I���ޒ����cp�]h?^�=����%����XR�i�w2��t./�7��x��Gn_z����2p�h�m7�5՜��^av��2Z�њ�x�mU���e1t;�\h��b�+�;��V-:,]՚/)I�xwx����u�f"0g+
�z矻sgj'��S�]�p�T� �L�v��s7@��\ln)����*��g����1|\���6�����, �S��ԣ�����[ErVĵ-d<Y]��4� ��w]j�u�Ѽ5��>�HK�Z�X���h���Z	[��ugVv�-Ʉ���$m�u�`�]#9�Cܶ�2ё��fw�f�����U��g|5�7y��8W0h�6��[�������m��`/#�/x�Zv�kِ�[; �IS���v�����'[��k��*���Jir�a�!n!�����v�PQЫ1Y۝�gWqOy��m�ڼ]����&��:��ԭ|η_'tv�*Ly��q�E�	����5���g�T�u�p����z�Ӽ��`���pZ�mw/�O�:�i�#�[���J�\��HͶ*ͼ�2�N-k�@��Ԇ=���,&�����Osq�1!}����Y-ݵϖ�q�L���r�L8��0�:�Tf^d��S�l�[̦�nk|e)b��poa�4�J��+�V�:����M�SV��T��rq���B�[3����|��gN��!h�g1T���dR�=�\�Q��{�H\��R�>�|S���j�7�I��n��Z�j��EoCus|鋦���bK`w�PM=�m�:60���@7WĲa�G>�LS����<x� &��>�{������V*HDs`��pt�*��҄��֌j�m���eq<Ø�� ��:e:e+�YЩڌ�/�0���p`��S�Y��;��9�g��G�۳�h�]��'A��|��ʒ$��B[�Ӛ������Ф�g6�v*�#kVNS��=S9�C{�!��Kixm@��xv�wC��Y���@IJ�`�V�4Ӝ:`�ڰ.�P۔L+�܈�Z5��3RI[p��ۃ�L�=:%�,	F�mf�m��u�-lԛr�V=���H󡪬ν�d$�>�|"��̥�4Jȗ��ф��lRЕУ�V��b��)�T�7��S�G^S{�9�UV�rYǭݬ�Q�`ـۚ��{6<�;���Ҹ�M`x�zg�{��v��<�	x�l�F�m�i�W� ��Y�9.������/�a<�3	�2"{�����$Y�Yx���N^s	�mFh�(D˅��{�w����o��}��;���&S�#�����Y��a�2�Ԡ��+/i�=���hަ�j��Ea��}���7��X�^�TP�&�?8PT�����o��ᛌ�~"Ës��Oa5�~��#�w��Wg	��K�����݊�6��lu͗�N6��.m��`3Z�U���d/�t{�:.Ѐ���-=��Ke������x��A�����}��]M
��1��Sɢ���w\I�j���J��D�"�|Q�S�|��:�F.�S_V�5�d��'Vu����8�E���9�I���\�f�v3�)e�b��N����i�:e�ob%�a��ռ6�ڔ�w�7B�<*p�#�I����U����G�Y������C*��w��?qW�/�l0a�4r�y���WSK�n��V�f(H�=ס\&&i匔�iV�\ܐ���R�yZ�����n����R$��[�D�s5ՕG7e[+EԽ�uD�4� u�J�#is]�s��vTU)Y[��7v��:��#��N�eۙЉ����W}�k�E2X�>/F��"��Y���]���?U��w�>�<Y����x�.�fĿ�<*��gs���;��;p�+Xj�{��Ft4ۧKz�P��Qy�0oi�n8������ip����B�Һ��D�DmƵ����� %�k&��ʲ�!�g0lki����2P�v�ɂεL�"o�\�^KYN��`�K�j2�g:<���]Oɛ��=ɻ�	?:�ݽ�Ye���d/yy����ˌ�5f�S����t8<sd���1��h\�*��ҶNZmJQ:n�gcJP��]xYg�̡��pZ��ӗe�*mLv�-X'Ӛ��uݖR�W�q�ǻ�m�m��-9�Rd���ѵ$�FXsM��N�z��E�2��l��-��~��d�۩�VZչ�Ԉ�ݗv�,���&�#����a��K��|�[0Qx�2�g��x��� ]YWc{)��P�b���`��*9F@���̮��07�iF�l�� +���;l��i��m\y��ap�m�bvP3�J�S�f(��>�y�B��͍RgQ�@�r��ݘə�pN��3�(\-��۟
�`}�nn���C-r}0>*]��l
�-�"�Y�n���cr������[���m,�:��-��8����BITV���]v��^�d�FP��pl��ڐ�P������ޮ���EQ/+s�K꼖1G�:�����V�����E�i�E
pw|5�Wv���8.�ڡZ�z�~������-���C����K�3Ol�9���Õ��ǂ��Vsss�)�M�7��;J��}�
xc�kxV��S�`���Ric���������c��H`gnb$����0�}LS�	���j��v�nݥԹΗ��WFq����r^Vw\�jq�8ε�p��3�%����ÝT�aP�+b�z�a6]nF�NJG%ǜ�ek��Zٵ�e�H�Qf��5r��5�Xx�N�yXYOo0�7�H#�炥��XY,�\ݠ��qD3�|_�=�.a&�!��D �^�� �������;+�4x���v+71c��ޠ�t������,�Eo�����=�ox3���n������wipx�;��4��:2��`PT@���!�+�W���Zb�
�
�r�Tm���)aim���7c�l���x��M�-��Ί�R�=i���"����P�L��Ԟ��Â�f�;��4a���%��oս���p�
�J�$(Pߴ!�LVZ�v�|w���WnZ��z���:)�u�vO
Z�߃���+L���
b��һo��9��֐�)pd
ҕn�gB����yF�:�b��<b	+]ϔ�5���]��s��p���82.A�����W�EP�$YY��W'�k;��H�23pQ'�f�XZ��w��qx`�'�t�5�'ma�y�^*��X�y��`����jp�ݖm���Eƹ��e���mIԉ�~9D��y^*&�1��{Etp\�[�X�T;���}�B�[���^B4�F�C/��=J���]2������h��'c�Q ��ֹ=��
3�u�L�`��T�]{����iU��� ���*d��mN�VN��ny��ŉ7�|H����(�i��hs��c�8���b�v6�������ײ�ksɑ�J(:�{/�{i�W%���e��w��=CuZā����n�<��+�W[����-P;����Oᴯ^��wa�	+Z�� �N�2f�쩒#5Z�9�E\�F��	��ب^uW�x.�/jƠ�x����#)���	���ې*̩`�3V�_�]��y����xk�l�{DZ����N��%���n�QB�]h0��M�kfv����m��k��d/���%���y�A������Jp�TxE�k��eL(�O�1�^bB��u�#��["2�� ��N�ɂ�	�,���\[y�aAP�a�b�j�m��m���Z�Y�6�c�_q�f�����r�^�v]�9�1�[<��U��+66V�/,r��\-�q�z�a���B�h����9d9/n��YkY���Io������wxF��E"&q��[w������Ee9�u��Ҷ��4��j��7���oVfK�l趦��=�������8pk�D�w���.ŕ�8#��U�������VF*]�TufL]]�Lj����ped:k+��#)&���M�cr��Nr�W1}.x�W[۶��j�����d�eS��L��n�]L�ވ��:�l\�v��!>�����>�|9�D/��[���m1��kF�@�齡9�_$�ph���e�vD���eb�ư��o*��&���%F\l�\j�=����5^Y�SW�$��uּ�QS��g 8ZZ3�E}zE\��%�1j��ֶz����6�V��y��Sδ�9��v�d�Wt��ql�DG����/�'If3Ǥ�Qu97�tYrb�\�ia����hme���ˇ#5uzA�g��;	��%��ZH�Pф̲�f�)QX5�7异f짂�:�B���s-�ef �2�
�#���B+Uݷ5�h��QD�#V�f����x��C.�݂�9����-���&z���c���X.'H����!�|h���(�R����I�ƧC�#o0P�sc��'�E�|%Z�9[�H�"�ed��Jd���d�q����Y��ĝX)6��غ[�`�4[g�۶�'X����]^>0a=D�<�CC�Nt�6#yH�Ѽ�Z��|.Q�ٝ�T`U�t!�]/&Md]͏zR;����@��Hr�G"�Z�-�L��'�0`Z�z�^��c��c�h�H�����qK�ۣ[���,�͐� �Յ���\.��	�P�:��ᙱ"�Os��B:V��bqe�0xd�:/'�7O���\��k�ݓ�0b�K�KK>?3Q�//Gm�te�b��N϶���=�7a��7��^_D�u��xy�Z7Tt�ے�����B�j���'�F<�$��wp3\Ӄi٣(ùۚ*�E���>(u,M��<�]��\��;�/����;���5���|�S�VT,3���,�x�>�pŗ�n=C��ۇ�nC0]g�d#K��pA��n�n%c�״��W��n=0N�p�ow\����la��n��h�)m ���4����@t�wni��e�Oc�\IUV��:Ypu���0<L^`�� �����m����]�v�`j˱��"s9�n�����L&�"uoQ�nv���xkD�+��x�$ӻo��}sx(,eM�{�+]��_p�����:�}}\5����_<��[=�@���14K���. 7'�l��J�S���N���
6��9`+"Ϫ^��;f��.�60�ӗ� �+*]!��&�!nH�n.�A��7��+�����>]�T=u�Dtq��fK�L�QXQ=�R�P��Ev>Y� �g��K���K�����Ӑ�N����R�΄N��`Z]�fFv$�.���9��ZdK���.��OJ6<9��rY�ԭ�l�܋Wn�ZM�R�!��@S��@�M�6d��M�\��
�|jT���}�۾o��G�X)��l/L���7�s����t��챱�h������(d���?k��}���׸�D���nL�э��ͬ�{s����.� �B=u�)���O���4�0�óft��,*�ξ����yώ_u�*33k����{!����O!���Ѹ���#q���޹bx_,������E4�<x�յ܌�ț��[�|}W���ɳb-{�}�|��G��0M��<�����o'���p蝭�s�g1�8�ۚ@��cQ������e����:�;H.bp��Q�,DL*u���.!��YIas��9[̞--.'��@���@���H_>�VxJd���{�D�k(E&5kw�:`^\fˋhй�9�1�s
|TF��yx7��͉��PǚpR4�����6**���Z+JEf5��UUĠ��eW�+LnZDF"��U�V�+n��,(\֍":h��*��R���q��(���`���Z6�)S2�X+���I���9JT��U�***0TPUD����cR��Uj˙�*cDQE�US��J�,��"��2�E��h����A�˃-�,c���D�#��(�m������Am1�i!TTQVZ
U�ժ.�E`�5B��,b+1("�X��*i+1��1Pն�Tb��c1�Eb�F����YDR�-��E
�j$XKD�����2�K��U��UQUDuIGDJ5m�YUU�c[�f\`��P�UAAY���\Jň�"�
���`�J�%���lU�+�cj2�c,SV�Z�m�Ma�J�4QB��R��,(#�"1�,ib�Z�
�*��*��������pJ�U��TA_��������\8v�O:Q�&��lk�ꬴG���ߝ%:���Ӂ���Lsj^SU�ֵ�9Һ��{+�q��?��Ye�S8�0I�9n�y���܎�==��0=t�_\"o]��B��]��e�xfw�{�;����{<Р�7e�r�<��J�����S�bJ�<5�ihx�,ɽ���g�tG!�V��G ��쿌~�| �R����p�4�{مZN���#�Q�m|���Q����wɣ����rZ1Q%�E$;=p��9/0�s�:1%�ל�c5o]㇕z���T_�����ޚ�3�T�X�J���.�*`yչ��ůl��(\Hvu�,`�5�@�Q�����@ާ��N�W������*vi�T�.i���G�U�,�"�S@���s��n b�ڐ�n)8S6�w���=zZ�T�G#%E��:��]�{�k�X���Y�)�uW�|��=CF2�;zV͆��=ݩri��1"���.�4_��x�:$i4;qT���w
�3��DW��q^�茅-�����:E���Ģ��S=�[��
�b�!uAG���:@�ip�}�W���&�z;˦ �ٛ#8� j-�7���U�[O7W<퍘�D��+�����{v�<�hOJɗM9%����¦�*�}�#��"�L�!�'m���=�nm����ɉ�3�����5�-�Ϯ��cּ4Z�΁%��^�#Pq>�:>���G�K�<�pӝ����#�i������ӕF�(�F�H�ϲ�wu�Kc'\(�6)��`�nWF�4�h�m5_τ�Ϝ�0���2k����ﻻl��t�U�z+a�Q7C�C��^��l���-�k��)�E<���IL��P�l��_�C�c@z�8���b<iЪδ�M �]�%#��~bc�u��ʪ;O$	�J�&6��?;���8�A���8�eH�d)"��e��2����9��
��=~��s.{��%0zFU��;ި�c��\��r@����*$
����NE
u<�������7F4���3�6��Up̓�na3���*��Ј�[�<�f�Yj�d��˹.t������[����:6M@C	��è��(XR�Bj�1X�}�V*5���o:i�5��?��O\>3����g��H�\d��_k�j'B Oݲ�M24���n���qT�2�.w8��4���@B}�Ճ��ɷ+�/M�h��{T�3�m �.��Q��:�d�9�C�\@�������O��2Lb�i�uZvЗӟ`���v�V��)X������cO��и���3o��I��om�S�Z�9�Һ�	�w�ظswFu-׃��OQ�]S�َ�9t,���]��'zބ��{3�s�nX����(8s<�C<�\�b���j����P���0��܈���[XjU %��،���-T���Tip28�kl����y�o��
�3��y��Ug�JR���^�hf�{��'g�֖yP�R�40�2�}�z �����>�}����x��ߞ����p5��weW?�uօ�_t���sKp�i./��vi��5��a��ꌿ�ۖ~�ba}ǧ9���v�,|**�ˊp�^�����VzU��</R��p�'/M�Ҳ� �)u݉�x��f����w��ا��m��P]�	5o�;�![��|�
S��ݹ���F���6�{�����n��;%t��F*$�� �x����mBF��q�`Z^�Q�Mw�G�MGO�I��zLO��`V�tc��!ٿdt2�㑪AQR�ňC����wp̞QoJ�mw*JK�NbnW[��h�
]N���[��0���x�vr'��wk/������4��Wl"+�u�q�2�����K�lj�]w�Ru֟�R�]�k0t�&oNB����=R�Jz&�{�.��SA�%�םV�Z�Y�������X3N���I/��j�Q����gV1$�K��C죲�Ю����٧yެ�x��Q��[�/yN���/ʻ���bə�$l��"�����Vꨑ����	C	�}�;�uˡ=? �����]F��g�A���V��fVi�R��'��Χ�#c�yZ��~݅�2!�MP����Ö&�k��j�v�8`	j$���g�y�P�s�;�t"�����������T�kS|����3���uQ5h��ECt���>F�#��Ϊ+x��,���dD�V�2�}�g�v��
�1�7�5):\̟���<�&,0�_D� �,ۨ�П}{d˝�r6�{��o��Xp� �K�<�\���züa 6��.@�꼼p�k��"��(,[٦pa0��9�ԇ���V�y�^8���2��s�o��^��D�t����E��|��F��ŤᶗP�1*_�i���4eӤ�ӛ���y����]lf����Լ6Vs/��`�F~���u��(k*#�W�iA�[��x<#0)v�9Û�5�)���Y�^�{���}*��7�xʪS>�]tiҲ�+��) ��t�Jl.�nO�9x0�ɓ8X��y;X�a�l���}�v�/.�v�RT��¬�Ӽh;�UX7=��������u��]�Q:r5nv�ع\Cͽњ��us��#���*�����B�U�j����S�+h��q�qSzuE�� �F=*�9�<!�㑥�Ӷ2mJ+���\�bU!���v�yB�;���{�-
��,uA|tJN�0�
�9D`����ܺ(tA�)���Aj���O)�W���b����9�q�+��c��]����sZb�v�oX��#w�4�pz��b���Ĉ�\:7n����:���2�l��oY[��`��z��A��sH�Hn�� �;)�a�U��w�@{��|�^3��.�*�S��1p�U�qjzUΨ��x���=�ʰ!8ٌ u7�,�t _�C�����l�T��_Շ�����k��A�F�{���kk��3"��6�@l�:��,�˒���ņ2�~[s��e^*�ӵs�R|�FH�2���i<���Lb���GM�U��C9Sf���e�h�����������2�r�s��yI���lS�\
uo�U�����UN��}z�kyS�69��ӏb���[��*���T��X�Źu+�=���l�ؤu��kU> ?�7�<(o���d���5jn�$Q��@�˶���<���������K&��&g���U�]��́�@�<ww�����eD�a��W0��t��,nu��W�X��&���)۬'�9:y�t�6.�W�=��g��+O���۹D�W�j]tyvģh?��O�D�uL�C"�U�l�� 1VԆ"�_ӌ�ඌ��23����������hf�!���!�س��G���w���h8�!�v#��d�"T%�o.�[��wL1ۑ,Fi�����gڨ�ƃ��L���Z\~z���?b�QR�[����rUb��/K	��^����Չ^�>�@./�
�Ip�U���v�9�G7t�d�����q���Gҙzz"V;����a]3���|�����ѱ/]���rV�a1�����e��D�ɻ����w�3
�<�&��u,�f�<炻��Vk�0F�D��$pϧ�,8LpwyP��\p"�S��JwY�o7�c;��*ӱZH��Mq�P�)�Y��,�[֝S�ã��d�w�A}ྭ��K�Z�mLFފZ�u��M��"㶶�+a��SRD�4jC,@��>�S�����U�jMh�O_?oq��ᆵ�qi���-��.NB��9<�'a�AOݦ_�>�y��C��C��S�;�ش@:�OohP׶�i;�eIBi�f{����{�#k�r�gHQ���P]��K����5�u��)�o,�xw�'�5�1���
����-�3��
����BW^[u�h��a��]Ä��͇'L'�k�w\w1�|�ث�+x���u��ǎ��s<9r�6�O(�~w���B��T:J����9���[����=71Ö��T�YC��C�����*�����LaA�MIC`)b�T	���0;�n��O�2#=��ү���;;�Y7�3,0��Ѯt�� �mu0�B�,�Ɠø������O�#FX�vt�����/ɡ�m{ޭ��P3X���7�-U��k1�P����z�ĥ�\���+Ys��=ځ���fE'$`�界Q˲��u��jO�{�*��c<�)[;7��v)�������`T^��V���g�e!�ko[C0�/c�A�C��Lȷ2��5]�ָ���+�_�?<�O7�:L�xS���F���X��D��;��"�*�k�4�
��1�E��ɕ�g�1!Ti���ڧ�v;�n��埮�y��6n��!�NΤ��i�9W�����.:e��=�ŧ,h"����4�4%"��[g�5�g�O�`�5�|�J����eV}��	��ۆ��Cv,���ۈ�+�j��,�4l��v�S}κ���nm��p�Y�������t1H[�S�knU�Ag�fFl}����m����T��=.c�pY�f�mv/*���7}�ʹ��j�G5f+����g`֤�NK���i�eCE�'Qz������;^�⁧ `Ԯ���Eg��Jh��?9��e�:%��T[�uۿh���o�s<��3G�s����v����\7U�hԆ�;X�
��3��=�p:Y���8|�G	��wK��Ws:6�cDpL�+��ȥ�J�	�q�
�nY�:�����9�@�'��Y�<�(�u�_k�9�Nb�s��e��N�'�ˢ|�I���t��'�ե;p㉺�+�&&)uD�e���JPz��$��*�S�i]��*7���%��z��[��B�[0�So����:�Ky��S�ug�ybb�uAGF�c�l�bk�ン{=��
��S"���x�e��n��M�ry�%AN�e,�𛝕}����yۉ=��o�����=��VU�n���T�����z����L1~4E�V�]JzW�{=����3�N̷S�C@� --���}�7s�P�b� h�J����\���gr1�v`P�"Ը�(�[q�ۜ9�+�����p�=��
ߏ���])l�����s���:sX91�#<=�	x}��R�;���j$r�OP�d}�0D���i��]�Ii��ؑj��λ�8CZI�A�����x
�EshݣR���Rv�p�����)��� 7ԫDQ;:%ZU�� /�cC�+NN���)hW7��K�,��o��7�Uc�]
��d�H���l��(T\�#���dFg:L��n���Ņ�$�r�0n�cJ;��}b}���npK�#r+�<�7�����Q�|0']g꛵���E"��J1ٮ�B�'���1^گ �f�g�T��*�}���T��ba���umr����%�o��b.�84B��B: �v��OQE\�!
; v_�U!��e#�*�}͜�����F/��a/Rv�������4<,C���ppJ�cM�sw,R�ݵ/����&dL��p��.��c��_Ɗ�Ok����x��嘃���
��5��5}�&)��/����m�"b~���%q����U�XJ�L��z��\fu�UwT���	o��ȑA����yI�]OJ���fUa��AW]d��{�`u���o����"@m�b��}�V �޸���ъ������!l[��ZV�FF��n�r�Y�؜�:2�&��������j�����Qf-�[Z㎡6�6B��PšF����H˕Cd��Yy����n#�2�{'�{�T�O��[1uu���Q�����]+�C�V���:�������m%lݗ�.���q;�2�1���ʙ�][�����:d�.䄮?�d�ʆ���Ƥ��ꩊ���|��e��+1�.�[����gm�u�O�i�j{���8ta�i�,���LcD�-��nʛ7��:�e���ЧD�O1�9��U�z��zxFR~޷��G:눽uJzr��w�q
5#ΌQv�;���y9�t�(9���V냪���
����(	�D
�{l@��\;������,��9�]L���H�~�cd��]����6+��<���Ƈ�:���4���0<�9T\
�U�I-�(-���������_>�i��JŜQ�w�}c4E�}����w�e���!f*X_�a���xv�4\k�\;#UA�,h9>��	�u�{���������Ou1x�d埜i��FB�%�۔��<�C5Uʮ�G���0��]Z��c��э�ۑ�ϲmߦH/h��b/&P{M��#-��㌽%S��n��Л�뚺G�6Og�׉����d��3CY��F�1I։�W���w!��>��q�˒� ��.i�jV�o�ݗ�����ʷ�򵷳X!�7�ur$�v��áw�u�J:@���wBQ��mD�����T��Xv+}j�*&\x�Gd0�%�.&����������6`j��0��̻k_u� �������2�U��J����p�x��`M�^��2cC�vI3B��;煪�Υ�$H%+T~x����Y*�b��D����o4-,�6v��֮[�������r�3�Ce�v���嚅k[NPl��mݎ[�Q�b�ch"P�z��]d}�8��/F��ӠC@�|��?���.�F�r�/-��iu�c�] �����Qζ�;�ONJ�563n��L�J���Z������OeJ»RѦ��Tv�Gz7�~q�2%Gμ�q��2�8N��S-P<�Y���Cf��KwI,��@^T�5����㝄.��8� l��j��m��p�&Z�r��+O�x�p{}U��(���aY�zؤ� ��;,�:�H�f���'S����S�q�Y�X�^��`
��ie!|�R_{��z�4��)�Mdv�k�'���
us��c9Qzu�;;nV��W�ͣ�Ry=�
��su���n��L�m�u_vM�dƘ�DQj"[[����ٽ��J�nsq��w��D��(�);h��v�c�j��C'q�� �M�Z�ֽ�S7�F�ި�.�P�W�ӂ�Y��ݛ�gK�t��]:�6wPI%L�qҰ��_qk=P�tc9���y`jv�֭�I��s�~��K}C%}���X�e�D�P�YXy�<5��++q�e���~(U�n\�*mX+qK;ǽOWjx) ��0�9��9���K���Tw.�wae�+�ζ��8G���f[ޑ\��gd{�9�/��t�wL����v@��e젳{���obVM�,̫���L|�lX�mN�o��C@��<i�����L��!��XRw6h�*7���:+��DWi�+�+:ekI[7V��7��қ��t>�Q`�}y�D�ZqZlekf�u��e���Md�6��9+�Z�>ݙ�>p���+av�Î��MC��"��t�e����(nv�\ȝ;͜��Ξ�9��c�bwK�t��Z;�%*kӃCM������e���ݳ�R��:�ݨ���BY)���H
DL�;��طal�{Aky�w@e�a�q��R�4圼/6��D�38�$�t����N�����f*V�%^܌5+o���s��)�.�j�<�|�:�ҳݢ.���ɮ��4���_&���W�ܨ��5ض1�2 ��S2��$q�!�=_��}�����F{��+�A��[��^犘�n@��H2����A�ylev�w(S�&S��o+L�+qFҹ�8��J0v[CD�:��ǰG�D��Ҵh��|�f�����E��] �M���&M]���3; صI3��!��)�Fa=��ۦ�����.ą}��6R���|Αś�E�=�:�����xz1�F"�eQ��E�ea����"�QE��KJȋ$�d�F1UkAE�֌YmkAa����ҔA�mEV�J�J��V)4�����F(�Z��PDQ[m��ڰ�%.fDF"���bB��*Z�e�l��[TJ5QAV
#UmDTD�[\�Qr�(%���J�[Fڱm���h�0T�*2شJ�ҩs2��Q�V�V4imTV**��R�+m*��QQ2�`��1�Z�6�DX*� ���İDQm���QYmU�DV�Ԫ�Ke
V�b�Kj���
�j��cr �3+[*�2��*�)Xm(��T�EA�AFҨ���#-,TT�Z�k,Q*�EjWqX��
V���VT�#Ul��J�� ����+�{\���׫|���{�̮@p��N�͆�%���D�����+�{�d�(��Pd���n�Ɋ�̓)/Q�g�� 1�F��
詯�m ���~M}�q�t�U,�I�lĞ�CP���;� i+�MS�q�hx�!ᔘ�|§����>C�ޕ�$��=�u�!���/^��*Ɜ5�������f�����I�}�Rx�g���Ϙf�+<7ε:{H,�>�bbf*Ţ�������T>a��gYv���3�ĞP�m��=g�� �N2����d���w��zy��￳�v�bv��T9�Xt��?$�Ne�4��*c�M����++%W����M!Xu7��+�X�gG�����T{3"ɉ8��ΦS�X5v���x�|dN��.������\�ּ��������ĝ'i��@�>I��d�P� ��S��N!X޳]�8��N�c�7�|�2VVm�މ�J�d�b�T��M���>dϩ�L�@�TY�e���O5��:�}�׾s�|�a��1����X���8�G�OP������bI_��Y:�bAf�u���)1�H/f��@D�~f3z�c��8���4 T���i�gHbm���>�f��g���}���o�~� �P�NӚ�ht�]��w�+<IP=N��+�i����\�ya�6�x��}��遈m%��i�<zH,���J���IѾsAҰ�'��^77�\��vw�sgw.�����+�
��~�P���b���q����k��
��;q�1 �{CY�,�����i'�T�Hc�B��/~��<@�8�N�����r��+u��͗}����秧3���T:C�p�}hY�%I�/\�I��X=��=I�L3�4�a�<O�{�I�I�p�ßP� �;C�ĝ�Ry�vÈb�C���ҲVT˗�s����Mw|���z��I*}�z���f�T����AjzɝG�$��F�κ�Mg���{�!��O\VN��IP�l�&=�́�6��'~Xu�;H,��!����4����~{���]�y׹���g�3��(���U
�>B���@���tq�*VN�y����1=C�y�giP��N���� �C�9桊�RVN����I_S�L�\�=C�=Ir��VLI�+;JBk^5=�G9��)�.9�*TP���/�5b� vT�oV�H:�Fm�K/u���Vq���Q�&ֻr��K���˟������/,��D���� ����.�0$�Ѽ�.�5�%��e�]��_��?po�x��p�ObW�Fj�A]�U�`鴀};E>���ǿ�7�遈|����׎��q���b��l��^0�w���0� w<�t���b|������@Y�3��G� �v��Hb|�0:��� �n�b$'�y�~�Y��y|<�w�~g�:���W�ެ�
0�$���ĝ�뻉��>C����'ɠ�0�&�M���6��;g�o$6��N�u���������^���3]��{y��s�i�!���쒦�m
�E�^�>Lgɤ�:@�VJβ�_�bJ�N�q���V8�$����{���q& i/��c'�+9�DH�>�	��뙍D�u��U�K��8$�
���u�z<���v���d��4�Y��Ĝt�I�(bAz������T�m�*T:���L��C7I���$0����z"0G��l��z��hV,⏹�3磊j�RV�eLCi+�x��Ӥ�
��/&��D:I�+/�����!��\�YXmۤ��3�J���j�Ă�M��|¸ô1�B#���@��dJ��M˞�{���ﻹ��<CL����!�AC��v��hc'_XTx�&l���x�N��z�'i:B��a�d:L@�6�K�a�+���2�&!�L}Në"�2T�t��uǯM��[ηw�^u��7﹜��t�`r�'�_l�3�<�C�q��M�i�C2��'9CNk4��T�!S�� ӌ��!��{����u7�Z�3oI1%B�%f!����^���]��������f���ȡ�A|O��u�I��{��d�Y�%{������ݲ)6�{a���q;~`Vq'5t퓮SI��Z=d��q�4���1E'¢�}�>�(DBB|�]?]�5�En�xo��~��:C*T��L�6�'��5{C�������n�ă���0�Y���Xm4�W���hT;C�>��HT�B�oxq����>��K����<�K���M<�}��xy�7�x>d�P��:ҐR��w�q4����q�u��6�Ɍ>O^Ӥ�͡�;:��=C
vÌ�=M!�=�Xc��4�G���Rx���:q�I6�g{���Zw^�y'B��1	�Υ���0�U	��h�̐U�R÷F�;�x������t��%C�	��t:7��x�+(cG5[S�G�JQ �.;{�
y3=���V��#;/E��$�uU�aC�Z��U1���� 5Z��������_*O���h:aXWY<�]h�t���L|3̓H��T5>�
�'��ayCq����˧�C�=q;�P�=N�6���I9�d���A��<m̼�=��q��Ĝ}ߚ�xA|a��=�v���<�4�3ǉ1%N�u���Ug�/F��t�I�w��P���T��b,�5���s�:I�T���� )6�>�1cG�D1��*�%�54��߿u������_SLZϙ/���f��
�Cީ��t�]���xi���bK��5�L�|�'e���i �|�P�4��bs[C^4
��W�ѷ�v�����<�~�g������i=B��s��������2^��{<�5h�t�a�&3l�*��tv�P:��f�0�8�a�
��(C�6���w��� �H{=ך�OPă�o�S˹�\��;�_���|��&2��v�3��$դ�,��ެ�I�h�N�1'�s�a�x�Yזm0�+��;��Hi%C�z����%E���w����OY��'\�i'�_l����j�s���;�
���xNP�}���D1�y�X#��
vfx�I����Xb�v�'�F��A���:a�J�;��i�;I�;<�CL�eVm���i
�_;��d�vq��<�1�\��ԇ����ygWL��"0@G��ޏt�t��T���}�+I��;�*i��P��w�t�'[��;5f3�K�M�N�IX���gI��j&������k>g��V��|n���&��><�wz�u�\*��AT��0��M������i���g�k����J�����N�m
�ߘ�V��f����z�@�.��%ea���3l�*h�gJ�U>*M��cG3�k��4}#P�0}0i�P���w���;H,�yi�i�����4b��*��g��4CMaPY��wΤ�iRxg�L~dĜN������_�+�����O�t+*�/Y����x�WM*�|DF����T�:|d����Ğ�wa��ǔI�/�:�������i�M�=��m1 �y*M�I�(br_p
��%a����Av���:C�L1��
;�8�V�E:nk��=���Uf3����]�V�9����|�%EB)U��wq���TY�كC�+q���љ�m�$绂�]LN�a�u���Zꎚ48-YHft��)H�w���X�Ni%@��z@�.���b�p��Zu�����5�s�;˸_����Ԙ��
��*������B�k)��L���c�Y6�E��go�1'����{�x�&3�������l
��I��L�4þ{֡�4�x���t�^��Qc���o�d�7����<���Dۦv�^'�i�qa����fٴ�uN�hb�]Y��
�C�1���C����b$C>NR>Ԫ�tt�،���&Otw���p��f�ٗH1�Sԏj�H��x*}��^zp��FQ��Z�`��8z��; �j(ښ���4(2���?p�-���x��,�8��3��a�z�їȍ��)_z�<�S�f�5@4rUh��p?s�%h�b0E/t+|7�ʼ씨2�V}^�T��d��f�J+��#T�f+9�����6�5O�,&��G��\�y$fXM�f��GF3���8(F2�����o[�c9�\EƹG���X���r5aN����Jg�=��ܟ�eNT1V^�,`�5�@���t� W��m�Ժ&5kǞ3*Ͻ��/�X����w�.�v�O���i��R�t��k���I�)NT����}U��K|q� �r�����ݿ1�C�s�U���D�.���W�O��
���Z�1��YUbo`𾊊ķ�"��9vD�']M�gM�6����3�Y� �����B`�A:��g0UE��ȝ-������}���Z�Lu��Nװ�
[������]`��%�ϫ�
�i�M�a�`�p'�M(D����u����K���>��̳��2h���0��K�f�,E��J/^���RD�$h9�T���룔�A-����@��������\�Q���^�g����p����2���y������F�ܐ��Xf/AR@�L�R��=ň�eq��ρh��r�9�%'_j*�@b���q�՜�8!=B���f�UHU�L� LQ�yf�IΉ5\>�v-l���hu3�ٮ��Ǹ�[�]�L���X����q�4:[��o�kG��]7�ƥ��<#�Sz�{�}Z�`*wm0C}24p�pT'Nn|6K1�+�����^�	�9�FM�&���I�OӲ�N��+%Mo}!�!Q��g����ր#��T�_)�H�tYB,�c�ᵛdY�}��U������0�^L���0ɴ\�9 j�Ol
��Q Tt���`�؂����&����ňFi!3��X̀Pʎ���W�T��-��4�n�� �(�+���o��zRY�+�9E���*�u�-Վ�����
�n��Hs��LnE4ȉ�$�=��އ{Ԓ˜z.2�+1����o��f?>!wC�{Jzh�u.��bA^�c�Ь��s2ur{nH����n�M�$�7�7yTO�3s����-b�w^�t�)#����-���k8��δ5rf�7Y�ͷ]�����>&��-�h,��u�N\��z�˖�d���Evk�Z�ay倣\ �z�<3�y�7�z�6T�D��(�F�����?V�\	�=�@��߶��{Hw�˘�t�oa�������\qΪ�����T�0��u3lȨNH�_s[�Q�����-k57>�~�����6�xD^�\��U�Qg��z�-��z�c>�sXpZ�Db~�f�7�.�q4��:�1��i��Djx����g���c4�Bx���^����B�Y��L}��Ƿ{H)��PJo@Rc�N#d�)G*��i���-˖��I��_wZ�L�gJ̵��n�v��u��柽�Q�Va���5�@sʺ��e?�l��U3=j�Y�L�W5�lJ�2*��aC
�����Lm��sd�m��P4��j�wX���k�sts�}�z��q��ڌo��1�v��r��O.O��_�F���#���Qԃ�g�)�f�]gW�'��mCF��q���]�"�#Q��pS�WBWy�C�DwF���4�tv.�:f��Y���86�%�VJ��$ΰ
<���U�͜���"T����`q.ǆ�kZ��c�+�@^a��wg�݆�M��ɜ��3�66ayԛ��-�y2ڮ�,Τk{Q�IV�^�,#!���C�w��UG���K�#��Y����l�\�°�Wq�ڕ�����HNwn�ٗ�����C�Tn/d�j�.�xѩ�%���U��y`�K_*`��2��p5����w��v���ԽK������O�����zi�!��#u����W}o�V�eP�.Lhï�k3���ӽ7P����O,E՞���X�[L ��pF�;�Ns��NXqdC*�)��0s�<b��c�"�zo7j���"��h���n���Y�������4����ȳ#B�:�w�O��a��q����\2l�壹�S���u�5��&p�,.���~��w>�5́��7s'�O*p� ��o�1O���uvwCuG�(�,[�\2�ɡ�g>�R5��@mBۈ���z��s��j�y���]�79$����C�`�����e�.��B�氡����ԇ���֕=1[a�R>����0��Hi�	��m��P��&Cau�HN#Q��''�FH���wkr1�-�c�+:��h��0�pv�D��ʶ�ҏŋ+��*�z�t��-��ل.EU�iKo*mG�ڹ�I���]*�y�Ý":�����%U= �/{���ESJ}��7x�$��H���(Ej<H�[N�4�ٮ���ܣ��}}��׍>�pA����Q�s�N��s����õI�+�6����u�,$r.���)物�"�[��ph�P�.���K��ƨ�t��Yօ�J�#S�%l�;f�R{=;$:��w�=�]wy��2�1!�����#�ap�P����,vG�l�U��;/�pr����q�ְ=M�ms�A�U�i��uX��B�N�1�8�b���0�T=ӕk�g�1�;����`9���uI ����B0�td��m|r��x�ш�b-su����L\�¤�8}=&:�Ѹ0x-�����:�%q���A�-�&0�\qc:��ފWjjL���9@.y�+�rb'�䮝și�bbb�V��0�c�}�8W��
ʜ�/�]�B��j5���q̱p�0λ� ]~hP�(VG�_h���׾/�ys��
��y�7S%��i�qb��p�I'sgH"�>�[�=;�7LS��@���v6�LÈ�m�Y�<������U�fp�&N�J���0��$�����!��y�7j�Ĕ�
�;$x[�ҭ{[�@�"˭�\[׈:Tt��+����(��+4��l�{L��N�K�p��ܩ����l�>ooj�k��=`�\�����2x�A�k�3��2��t��}�cfY�#b��Pr��]S:<�J�9���"#�y[j{��Z��	D��1��g
���f�6����31Ι��xl�C���q�E!�건�׾�̂��W�����õ׿��'abl�'@�]�ɬ��c�)��d�w��q�|Gzﰽ�|D7�|�qV�,g�/�J t�继T���.�ޯl��޹�����^�k�8����V�����M⎫�G2��+/@H��c+S�/���f�NP�q�jx�E�<i�ƃ�ڙ��&��%l����dyp�2d}4xk7�4:��^�[�e�s*鋮N�Yy�E��H�� ���\�����t� ���!�<+�&a�U��2�����m9|Qj�+7<]Y{��{��<˥����!��y0���ˣzЊ�s�)����}�~ʭM޼mFr��8�um�wt
���6N�۔�o�	VkG��]���:�:[\�C�k6�LX!��4q�CG��c<_y�J��Eg«6&�0�3��oQ�����j��Wժ�C�iΨE"��k�sIz�8j�X�uj̷�U�����Ad4�^n���>��d !Z$�`Sv۽��/�x��{�|����q���M�����W���0��sw��{��߻W���:7�]>�e$�<��e̕�s�������W7�����5�쟴Lw4�'&a�Qz�ϓ���̩	���RB+�B����N��-r���z9�yLH%Vw���%a��:����/�3�\��[@u�{%z��댞�Y�X��:w�{�
u5�����]�:�,���[����*���l��b�mV)�2���(m��5�<5�]R��v�ʋ�
��}g��SG�P�<��jw����q��;�.�p*1�NRl��ٸ����gԼ��n��*jC]-W���:���]̞�]diؐ���s�a��,8��Rȸ-'��H��ƾ���0���]f}~_'6���<	�'�j����"��/� �t�+y�0/�u3l�L�c#��1P\��N-i�z���:����yzr�����ݽ�b-� f�P�q|�}�5��K��萻-�^��v�mw9zS]��6��tG���,�R����W�ϳ:p2�2��Y��I�}��sF��\���]�z�5�
�>Q@r|�r��88�񖗴���g��>:�"L>�]a����7ҷ9�F�^�҅�����9���q��燋{���D���g(@�?���u�\�>{GF��a���'�daP��2V���k�j'a�JtP���d���m����ވ\Ǥv��t� {K>�4L(b�]�ʗ�I�GE(�W`�r´�8E]���u��%�����sE~ٷH����?+�1�z�q�(������e=N���t�׎=}(t�}�c��o)t�����C:�DO��.�z�v��_ <�t�ve�����bK��ƣ-nWPr�G�w��^T���zY	�h��_'�ӊ5λ�<\q�՝F�ڵ��<���V�B�voq:˲�,,�G��vG{���pf�e�:��QK�����Ž,��q漨�U�"�m[xbn����^�:�v�ۛl�ܻY��O���Zw�Q��ʽU���˅���ΰ�@7_��j �<��VZ���B�3�gz�>^��H��]01�GS�=*�`�����u^}���=��H^,�a�'�C����t[|U7��)�H��[�Q��Z1�����a��Rͽ��Xb��pZ����=.�{7y���Α՞�-��iӝP})�'���N:���\�u���a�8Eq�#�}�L��e"v�,�Y���v����u��V�����)-6�a��ˋ�־ �>�c��z3Q�ީϢF�V�A���rj�'-Uz�=4(�����7<t��s)I�.h4+a%�*��(�zN�D�����wHՌ�W]�����Ղ
d���iη��|.��]p�1mm��km�T�VGm��t�[t6v�N�U��G��!�+U݅��]��m`�A�:rB�F�������5�'e�%��;��6���r�����t�7:T��*.�b���eS���]�K��Y��I�g3Y=A��KE�x�g3��o)��]�rY�7J�e����y�pٴ�Z^�S�v���`(s���H*�A�O;T��Ԡa���B�����@o�wh�0��D��F��[��k�3��";�0 ZmE���
,�,:eL���Y�&���Vt��ExX���6���ֹz-��vU���{��%�W�t=~�����e�ˮ�e��'*�;d�|"��َ�}�Wf�\�k,S�"���E�����Ö�k�Z9�U�Aw4��&����]��&v9V:ƾF7���1�*Zx��+�pU�V�I���8^[rf��<9�k&#:� ��o,����ᣎL�t�
�u����>{�N��c�#+"噙�����!�p��+�fۧ�J�z!��JڛcHv�&�7�&�D33�E�g.�t�qւ
��*b|0Ӣ�=��efi��"��s}h4�ٕ4��MA����*	�G�ʟJ'�t�m|��)�j�h	���źX�"�(dA�8O>���Nr����0�ժ�l����+iDJ��b1m��ڍ�+b|�9J(�D��U*1em��m-��*�*"�TT`����EDX��ҵ&!��+��R��b���E\K[�-**�QVETb��+Q�
��D֪�ҌV.6�*��*$X�X�PQF1�[Q���e�[ib��aV*(����e�D��[b#V"*�(�U��i�aR���&Z�X��b"��1Um�FD�TDP-��Jʋ#D�ҠX��dA
(�*�Qm����EET�J�(�DV#**1V#jTH���1�TQ"*
�,c��*
V ����j��b9k�H�b��(��b����J�8��b�r�+P��Y�b0�\j��9J�`��B�P��R���7�f����_g��nm�����n'�����BK[��'��yg�cT��_G���B_u�̓ϟW��}�W�Q�@Ꞣuq�*��j�"?�pU��xq6�Mg�TE��*.f5�Ms(P�;Өk}O����uS��ҴŲ�*�G��=1���,�j�5��4�Xyo�a�
����;��7�T��C���� �P�J��4RwP����`�I�LA?8����6t���=S9��=�p߈��}�;H�@�e��`s��THW��#�N��T�p���o��((g���b�ƣxS=������'1�8_��ҭ�\�X�k�ӊ�EZ}��	]}�puF�z:�'ʼ,J'!�,h��Y��9���%�����Cz�G<���"�OK�X�.��Sf\�Ah�~��d��-����9(`b���6F���`�}���v�(�Y�5w��h�T��}K}<��6��n�G]����|��P��3NhV[�Mu���VM��l�Ԁ�v6LX�3�J1pK�f��y�P�M̅{U���[��W]�*�$?�Պ**�.�6�x_sk���y��U�*Y�މ�2�U����1D�ݎ*��A}�;��k�.e���_*B��1&�]�C"���'po�����}�7��f�$U�8��b�ټ͜Y1	�	�[������pfB�9E��>
����{%��;4s4G]y��I��\�L��*E��������#7����#��F�	ɱ+�j�m�N���iL�_i�;��G,��@��ҳ�����Raj,��)���'�of�*T `��Ԛ�ܨ�;2��x�[���x�A�N�����@���I�ݎ���`�^�Eً�
���E�N�:�U��؈����@N��6�L�&��&�_���85�{hw)((�*	��3�l�M��X�p+wc���ڎ�rr��'��r5���S���������6�9��#W�i_�o��zǠ4�w��s���x����1\�T>.�|��1��KVF7��9�
���3Wh�];���qڽΪ��F�A�$ߜ�>1#��O�|��. `��Ӕ"��v�A�F���7{]�:��,v�EA��T�ן�QW�ӇF?�3�k�I�f6*B�"�Z�Z�^[�e�rN�>���d��=%D�l��3"I�u*a��ɍ���������HXm�i��t��#~��b��f3T����keP�^�(h��o�*g��Oi����k�c�3i/f������r�0�z�O�KV"o�|^X�L4�쮎]�1�EB�=��侠zÎn����`�S��.�TBe�e��-�+�,�j�V�w��C��w��e��dn�q�륯KA�MGkt�Ц��F��Zw�}}�G��rr��X*lǲv��g9�9�Y*Ɉ�rWN��M�c")u@��@�UeWY�'7S�����N��L���)̱�X�<�*c�,ȍʃ?p���c!j��
M�n,[[�|FY�*0�� �1Z�y��{X����0��v�����$��x�/��/ѿ*/�\9�e�Ryk�ewG��OƟ{���7���%�KA1N�r�y|���m�=g�9��v��\.Q������,�@f���9��N�w�'�Gv�z�{e�^�3}�dXjV���Z~�(��a�(XVlxW�������Ṹ\�bs�ȩ��H����+�����޲�O{�7K�Yȗ�&`�u<���eqP֗��JX�u<&�6^Tp��@���ǐ�����/���eJ}���r���U��F��Ro�o�?8���,���!��O�!��N��e�*t�b����͙o�']�ڕv�Vаy�`m�<$}�F�a��mW���N"� �Ֆ�k%����{�=X�%������Q��*�<�ԻUF�HAr��������<r�N���v�nv	�={�I�p�����^�^`~�9��Mo�t\W�s�%\���;���aōM��
3M�N]�]��G,����ʜew��Ag�YK�Lwj�j������Z���z���4W�
f���2�e�Gx��|P��}J�P46��q�f3*э�T�%ĶnR&*�E�v�}Q!Q��e@nJn���� &sں��\)��
56<3]���O�^��W�f>�w��r�)��ci��X��PN��!��PQ�8;̒(N�tj�ښi�&*_�,�
r�L�B��`�]R���t}7���R����ͿOi�|֍SP�^}ד�5��v��kص؉;�O2�WЌ�$s��k"���u(�u���%
�|:�Y2@������6�:���Wc��jM� u'9q"	���S ET���hr�Ҧ�掚��jH�l�w����2����P�;1p���h�s]�2�����ܹJ��[w��}����FEu�uc���pT�=n�%X��Q�6��IT�ܻ#&,�`Wx�Wl �[ޢ�����K�f3K2a�S���E����Ղ�ni�]:8s��GAc��n��W;5�k�<l�.�ǵ�^ʣ���g��>��0�ӡàD�Щ�"{���/��/*Ao^QW���7�n��AY.��.W<��f��LT%�j3���C>!=�o%�ۂ^�h����q#;]�n�\m����<��^9���F���?f��e�-�(�ܹ�Ú}�3��Q���VQ��є�R�����>O�4Ү��?i�;74�)��us�Ʃ�d_�΍1���j^7{�����|����w
�b"�ﰨQ��}X�w!:��k͸���ƈ�א��PO9��;�='Ao����n��F!��B�ET���v9Fų��=���C�<uMl[������}�_�7R��aZ�8�����+֓��]�1�*��Kg錔�,tt\�Vw=�ԟ$��o�Nz��q�#4���D>N
�|�⺦��x��yW���*`�}��GgsZ5#N+&vp�q�,`��Ը�2��.磅�6yVJ�2�X��B�n�9���i���/b�����L�^S�3^�]B�J���E'u��W@0��� F�I��;�Ui��;WIwM*ϩ��8E΢�6�#c�ܜ�	���7ƴ\e*�MTHN6{sv&{�jq5��KĈ���ۊ��i��GF�6�7�Th��f,F��rt���#g���� �{v���cُQ��
!U�q3��ш��y����T�=bϩ=�S��n�-����>D,=\�.��ㅜ��Ի��ja>���a���ҳ�Od��Po�1ʗٯ�!�zeev���ҹ*o�X�f�������fVN7Vqr������#���N�l��I�PJq-�JrѶ5�{
yW K:������UU�ޓ�ψv��b8O�6b:�ˉ��N���t��>&��c����2�*��w��h-�[[��y�z$ȄoUѸjCsrj ���U��SA��~ӥ���x>~6�'�C���ˬtC0to����۬Ýf�vj+K�Gɪ�3#�f ���Q����ƨb�0:�b�z޽اy�R��k��r2a�_Gwn��q��� ��¦Y�މ�1K����j�̕�\߳�v��F�c��zU�x�a��I�;��.��@��錹���p�U)M���WG���&0Tq�WӔ��^΢��ʾC<�i�:۪�V�o�Xn��-�^�g9�N�A�?ۑ��Ɣ�a���Ȍ�)yW��p�'g��em�.˵��_�����A[���>�@;uw��B�����e�S��
4��8j
ƕo����q+�]��\���P�v�I%�Uˌ�m�f�X�ϝl�ٕ�ǣ���~G�������Y.��Q�S�����J��[`��<%N��t�����f;"�1����z2!.����w1*(��wyB=?��N����؄�fao�_�<Y�
��;��4+��]r*BL�K��˽�G9jzv���b�j�~�G���9�{>%�򘥬�yJ�u�-��cPV �6>�G��WY������"�Q4Zs��:Y��W��Ֆ1�6f�ݮ�,5�S��c���U��W�ܦ��7� M̎�E:������1!3��CPT�zq���b&+x���6�mp��nkp���+rH���UHU�<1�肙�4Ӵ�d4.=���LV�u���Ú��0���)Q@h)���̉�u�G
�b�2P�]U�]���Y�w�����p�k���;�<8br��|"���7�Ӣpz�=����^F����H>xT��.1+BE��b/�ph=Bw�'�q 
F#����rd��Gz���N<�=ݱ����P�"��]m}�K�{V�)�b�ʣ@
��n��Z�D B����/*�=���[ە���k��!�[��Q��|@��t�
�'f����8�h�l {T`2�5�E�|R\�,�6��:#8e����3ђ����J�,��р�LB}Q�vwcFj=�Yޞh,��4\�.��Xo�/�T�:��aUs����:�3��y7Nj��;W,��Jw�VHȇ�,췓B�#��鋎p'���70��zP����g�E�;w�Uv!{xHʳ��^� 6�����\�i�X�	�jn5�F��FV����f���8�������g��fU�*`=�2�����Q�n�|���T1�����C�8�7����t[:{��X��=�{s��+2�#U�n\���)t�R���m�׎t�t//K���>� B��|%�q�1H�Q���6�����#��6@��h3�=���
�]/OS�}A��J��ef*1`Ǵ�;����g'|"���E��M}Q�hܗ�ؙX�-C�9��_t�v�Vv��1���\F b�#S�N3ff3Jc�^��܂��;��3�5q��:9��қ�&k�Bl��{9uVrc�Q,�6ܦWf4C3ن�YLv�x܉�c9W�t竱����.��5�E}r���L�wJ�W�S88���r�E�QI�y��^�ꑇ���e��O��0�jb]= v̠$� lQ�yf�X~۹�PYZ�M����*�Ak9���.��?'jገ=�_�0BD��d�
S������빫�̔KšD�ܘ�Q��)�q�ġ��쑁҅S��V#��<(���wZ75�뉸}���D]���z�tX��x�(�����K�H��F�:�g%z	�uID��|��Ĉ��3Q����n�x����W���d�'�m��*C���0�����z�!t-�����|����]�4,����4�Ë.5Wi�q{�>�`���[�5��Ǖw�YClh���f*���k�����3=VH.�x��̞x����$��[{��V<JI�>�:�\�r���W�TDDF-z��of�T��Ψ L)����t�U�"�?db��rC8�0�䕼J�����T��X���o�WA����>�0=����ёG]r�X�Qxb.�,e�'S|+.jz9�a��8��*>iPf/�32��{ ��*�o�N$+�,�1��KT۱*���O��q(h�P�l1}3l�̲wk<�	������G�>CM��]dhz��	����p��U1���Ua�g�ro��@	NX�UP���P0�3lȨn@�\�N�U(�h�Rx�Ʉ�heĹc/쭸w*�o�1�F�*j�,s8Μu��'��1�C��m`sM�ӹ�)U��c��,V0DxG�N�E���~}��m1���\����ƭ~���;��	OCiڍ��b��V��!q�(�9>o��Z�88�񖗴�֪C.��� �[�>���^�z� �@�a�Q=�z�d��}�a	��zk��N���L��JI��Vu] �z_Z��ɕ
�V��2���S�NX땗�YϤ�cS�*v$�v�%�a�z�6�;��l9Ă}`b�����f%�Ƨl�r��Ɨ|�,^�@.�ǽK�$����b�|u��J���f���ޥ�����y-I�λ��Ruh�Pi���K�:��i=:C����}܄h(F�2|��J��L����z������������N��=��g��]w�Ϫ�u.�zw!�dp�{P��vJ*���h�L)���.��Ri��UPa��� �(����ڄ�����'T��>�#Q����Q.\�7%t�I��/5&j�&
�
�5�\<���1"OK���9���|k�))�;/�Bs!a�F��
�]��,�-Ht��ht��4k��]���*�*��eOa��9������+����;�fp�q�ZN�勉�U� '���5�����H���EK&&��H�X� [s=:ٴqrZ��75�Gq�|��:T�r����Ҩ����2�~Ӆ���xOر��]�Ko��y�=HK����hwQ�68�R�fF2�0�u(�G�X�΋�n�ޭjH��'�̯2�{jl�=�0A�Ʉ�u�!�UK7�h���.2ˋCV���˖��Z����T�ӑ&<6����읭��(x��F���N��3����(�7�u��R���]֣v�v��3r��5 ��L����~��5�%�J�qVr��U!��!p����ݑ6ח-O����5h�֑GˀpQ�G	ُ� �1�c/�{Tܡ����΂�I
��&��\�˫QӠ���%��*�tث�"�b�*ɳ�t���R��죎f�����峠w'N����2o�+qSs�p!�i�u�b��	V-�����Q9���j�.�<yX�L�:9v�4N���ȼ����O���c�J]��)���S�.�<�\��ٞ<�������M������Eӗ���%2yue�OS��e*x����A��"��7�k��mV�U��Sd0][��d���68Tsb��E���N�޵C�;M��`>. }����$ٸ�;�nE!%����QmԘ��n�8��ޒ���zWæ&�7�,�I�nhۭ2wMp��{[t�а3y�:��%h�����G���u�-/4#��Н����� C[�F,o8D�^������G��aw[����`�X�Sw��x�8�F�}���:��S뙢+�r����Y��1�(W@c���z��WΞ�uy�ޖ�U���nHF!�V��%�jK�yC:�k@J��̕+�_M�u��r�&�3�$w�E�^0�}W�K�tQ��hW\Cw����[y�}��ㆹDN���cW@��0R��R��Ȃ$�a��6�0P��3໱n��\�ءؤ�Ne�T��Γ���%jks��آ�V#j�����J��Dǌ�Ϲ��q�+�5R�#�͎�^݇X������ @���4fa,QI�{��K�!��{fZ��B��Xd�VdL�c�c$�p�4���e�Z�Ey֪��Y�̝�B��t�8Ow(ۇ��dQǖf�a>����xzG�:���O4�n�Z���=���E�9Z���\篴PDܧ�4O��]O��:nN��q)���w���iv��Mt��D��Vǃ�:n��\�"��:X��p8(���X�[?s�"���#��	W?9�����$���G��_vJo�֎ُ+W/Q�4�b�hV�y�x�ZB��f"���!�E�T�,;�` ��B�Րq��h�
p-�9����E�8H��״\/5��)�V\�4D
eԡa�x���c2EUَ<���� �)�Lץ��Y=�N؊:@�h;�����-H�/���J�.�t݄6'I\/i���8����{��[n:��5v�o77,ɐ�F��g[r�L�2�H�侹��C`���t�I���ni�q�˼/�zE�MO�e>IX!�hܮ��ig!A̙뼔���$���S-et�|'�<�=[�;�5})�-ij9e�U��6��Czs�)�Qٺ����j��ӓHz:$�~꺺�b���Vj��h��km��b��"��""�AĢ�r�(-���R�W-�$Yb"���ZP���1%`��V
9J���J�AĪ�b�c�+�(��"��� ����1H�e�"ȪLeET�R�U�Ȣ�,Q�L�T���)�F�Um����\h��,b)\pjVQ����b��r��`�1ĔCbcR��� �eTX�"�i"
,U�*Q�q�&5YFUh[E�2Ŵ�"�h�-́F�����QUT�b��Qd*QRB��H�5$�[hȌ�f1@Z��*ED���IFҊLVe�!R���Ʋ)R�J�g]u��G�-�j����Q#�y�I��3$��˴�oݬ�=�^ޢ-^i�}KI�����Z�\��]ըZKw��q�>�>���l�v�mb�9u�<脫������.�#x��O�y�!*կ3*��L:�@_]���ĺh�_xb�����]�F(os���ϮQ�Ä�7���X�*�CY�j3y�Ƴ�x�[�^����-l�����V��n���:���?;~C%���x�Mh���aMVX�޴g�q�� h�\��r���ޔ��)��,1�*��ϒ��𚈵��U���J�{G���B!�QV�L��uDLE�V���o�|���#�8n��9bX�ٰӫz�#g4O-gNʮ�E0�8�۔�t����ыT|S:%�v���4$�oE˰�n/�]�{K]1���!�@�G�x�<��t�
���tyW��Zᣆ99���[oz�'�4��Ѩ�7�Ǖ׵.�|��w������h���0�F�����M,�b�<:�mq:#�����n�xr�1���_��:W�������?g��uC���9�1�2��1��1p�U���i�(ŀ;b��c���� $|ާ\�^��\rW,��i�wK��\� �br݀opA�B�F�,�Z��D��MK�8s�)��)�f�"���0��u��ڇ�UnM*��N�7�#�ig�4�ǟ)l��wp�Ͱ�D��3z�u[�I�խy���/L��ӹ�����fe�W�U_Um�R�|8�N7�����;*k�:���&,Lv�H�i;�/����-��Uwe:-9�;}j;��Go�W
��1�[���{
v�aKjVo��0���ή5>�	����,ۘ�ݪб��&��Y�r�ŝ�.WƮ�8�xS���S�|xF���Y��{e򱣥F�[�q���p��s�gX��+Ȁ���U�k�h�1�m^ ���om��n���B�8\@�s�b9-�|BO`�离�dY͝�����e�f����t!�2�}Ioj�F� D��(p���-;�	ܡ#���*{�;�|(�A�������;�OK�<6�+o���b5�@�nejvɸ�sn�K�i9CEIQ�cC�/Z�K�
;A��jC�6,�ĸ�k"�uE���yQ�������J�u�1r��!��E�dM��9�u}�o��+����+'��>�y�0zO)ӊ�6�$���m������+o�ê�*%(�=��Qw��^��������h���X�q�ɝ��zE���A_gx��!�Ec����6��*Dw�7�۵Ƶ*��DX�z�6��g�F�\j�aN�A�y���.�P �*�n���6�FXRI�nts��f�H<�����W�UT�2�{�=�4~O�\M����Z�麸<����ͬ�7��׊Wm���� g-DͭqK���>��j��&Қ��ʸ;�go�����o&-��'س*ӄ�}�q���5�n��;�g��UC�=sZ+U�.㙜�Z�\Ë��w���֍_�G��种W�o��
xk���Ї9�Iٜ���G��=��3џ��^tX��y�|r�M��3���=��#.w>-"F����]x١<���z<�s���8dKx��qG�%)��_��z�f�BnZ��h��u��4���}/_����t�����r�g�T�IqQ���yN�F�ָa�^-s@Tv\�'��i�⨼��XqF�Sn�qq��-�|�C]䉸Φｶv$�wd�NW�f���BB���Խ�>��V�+u]�'��9��D&iy�2�l�]0��z��Gu�r�^J���HS6�i�F�9*tO	|Qj5֑����:3��*<��H=�9tH���k�k@��\�Ү�����4����}�'���
�mؔe9���U}_SǶ���>��&�!6��6hz��8��l�����SO���X=�KV���#�y�Ȟ���G���<Ov�d�zj������C�bo��7[qU@�Zon1�۔�W�_e���]y�Cd�B����o]{y%�4��-.�mIJ������D%�<�7����S�k�w3h��W=��c*��X�»�S�|ZWBݸz����v���qg���Z�'Y.���Mn	��b��@���� ��E}��<�nt��OBv�3;J����K�ͩw���=	���&��}� ��:��Su��yjk���h�죑
�O\�U���@]�p��ԌpnM'%��	����J�C:���K����d��,�.%nH�o�����,�vi��cny2龧l�}edu'p���Իr�>�G� ٬K�\�[�%X�X�h0;p"��ř2���i��Dd�p��AEn�j�r�����h��婲�+��e6��[Z�wB�}�I���n�<7����w���tq�WH�d�\]�漪��9��� �f$1g��&K�8�es�e�-�c� �퉜�gV]�ﾪ��ގzys����H(��T���ʟz�~=�r��B�90U��ܸ\vm�v�o9M�:J�\1r����!<z`���*��r�����y�./����{���ﶾ��W����j��:���S�9���'������pw�Û}ͭ�W��5��츶��>�+�����y��lȼCK�Ŭҥx5�]̯>o�����^ ���n�Zc�$.�,��qP�;�x��yزce�셍�N���v�o��yg�M�<vព2j���'���,�4���T��r��x�w���˛�wm�P�f2�0��[K����N���"nSJ����ڥhN��\{�(t�:W��[$��Y��~�����4��.��vW����O��,)������Gf_G���UI�r��Q{|�^�ۅ�U@��.~��毣M'���jeΛ�H}aAF��J:;/FH��q��j�Qw��9�6�^���}P�̹cn�k�t���g�Fl&�(vcH��`nc`qb�i1S܆��e-X��n�"޵D,���I���ʻFηjbql�!�]H�iٔod�Ň�G���}ؙ�nT���h}��mC��w9WT:T��ת�.wj�������ݎ�=s/��\��I�Ry�\=�T�&ʡ���^OI�ʩ���i����Q��	X�q�nvT��c���c���<�?+�1Q�]�TzGiBɎl����j���';2�,�U��妦_s-M�T'�����zn�x�k@Y6kn�U���,{p�u��Ct�Ȫ�m���G��|����g��f��f�Et|��a.�}$9*��!=)��ʫwf�q@��t��1��-���u�^b�Ǻ�Z['_8���W`É���f�yS��끕����uoS��7Pe���O-��)�qx�֨����r�k��><�����	Q
4�-�y��	�¹��X��8��
+��ϓޮyƱ�ٙ9�����Jfm<�5l�W3�/�R��p���q�}eo.�%��w[
[�OH�ݹ����,4��z>�;�pܕnP����U��k�hN�Y:ŭ�Lb+\e�d�������`��̬疾�`4��Y3Dw��($��yu��΋g~������}^��F��~9	ȅ�]S����_Zo.�]Ƹj�n��D�;�5�;�]��#,%G�m}*kUqU���5J����x�*\�vrJi�q�%�_bx^�=�B{�}*ӽO���r`��g�=r�]�n��Oq�.��+ދ{�&Pq�R��Q�w�-ot2�p��=]I���V�.�z2S��v�\:0.�r�:�\��o5��*�f�}�e��]ƾ)�rakp7r�r�w�ۚ�>���S!8��6=&o�G��FfWӳ!.����]Ƣ
��.��[�Y8�+�V�����`ξ�b�[�ba����LW��ٖ5eG>u�{��͗�
ًɞ�x�/��Z�"�V�b�>E���]��Į����n���n��'f��q��Ȼ���~�P���3qΜ��/���ʈ��oHc� � o^�r�0�)vdƮ��>�7���1s�{zq�b=l0�'�.�1X�.S��D�+����۩R]V�}��-�8���;\ᗋ���͝��M��4�1CnZ�� :��}�4���U��t�do�����~�����9�����
I~=k�}jX��N��q'�4��e�}�����u�
��.�/+vsq����j�g��v�Iq��kyM
5��u���'���������]�/n�/
��1���}��q��U�B�_�銶��^vcJ���A4�<
:źعΨ�9_b�z���N�xO�6Q�'{����s�'.,!>!/QPv�<�u�1hvUq�*T�;h��P��_�P����x�:�os��oi�b7C���hԵ�p$��5ӵ��ƞ�o����1�X���[ƥA3��rL�J�wdCq��9k�Ƕ������+�C�}�M�j���������R���v�j���4jJ�䬭����ZV�vSŴ]�'^�Pj�9�ٵo�S�]��ᮇGe}%IK�E���LR�5ɥo�j�Jeݷ�G�N��N��$2�����2N;��2�g�ΎDJ;0�OnS;#�3s6
o���bJ4�c%�3�윅-u!�AGY��<N��Y0�#�t��o].��]�xR��.��*f��)jwL�w�k��_Z|#�"���8�y��[�?��;��X�\腕���*�`J�r���>��픽3W@'=+޵��us-�̊u���9���\8J]��=*|�B���V���0�sv^e!��q8HM�ˊI+��S���p�¯�a��l��]b���u7��wL�Z�#*]�ݰ�{�m5S�T5e�*�}
����k]��Q��!�����YZ��%�9]�ݹ�d�uQ��MC�M�,���KUa�˷j:5�U�Cg�k�����h��r����RƠ>�Sޫ��8t�[D<4�^��s.�|6�_��ˏO���m}y���b�8����;-*�:L�����]ŭ�[�5�x�U��p���|��R�^ӎ���5�����8��"���O���8�t��w�$Ag8��hC��,w�u��8Y�Z�}'�ym5�zyy��9�<�5�îu��FA��O�X}��#�EoL�)+�VCji%��Ĝ�Z�����+B3|�����[0U�C��צ���ֺS����֤*�54XY�[���p;j�f�s��O�i��of�˶�,sv9ldA4�\j�u��<|l�C��3�N�pi��mê������9�~��k7�h�T�L�=�1�z5������to.u�ޥ7�˞����P�~��綈�o�ҵJ�����}��+���3%8#�f-q2ԌJ�Aub��vTJ�ދ��v�k�|�4��e�n�wڒQ���Fv���ڋx�hW��*�
;w.�_Db�֫n��h��ƫ��l�����ۇ���v9WT:TI#^��9�]�r�䪛�C僦w;\W4��_u&�+��fҚ�R�����ԴE�=�BQ�]��\�R�Ulne�Þe�nyw�:ݳ�:��T�
��:N�dVSlu�,�i3-�W��Cy��W;̺�ո��B��n�WR��h���e��O0J��ђ#�>[G�쭈e.^f���9wz��ma��2z���Z��y��Y=����ȣ�����«�{�P���.׽�poQ�@X���(�ġ6�|6�J�J��Ἇ���+����c���%<,E�yVd;O��;eR�M5�J���dܦ��gVcw��
Y'nkʋ���kx8�$��0u�jR�x.;B��g]�R�pd�����-lp��s!�9S\W�X ��6i�5ho]�8-��W�Z��g���}�4�*���T�)K�aҮ.U����$(�C�m?d�[�ɹ�dCx���t��D��g�=~��eL��ʍ(�-���<�b]��b��īu���.���n��u�$�\��v٬@t�0�ؙ)����fvڙZ�+�#�6`Zm�Qxo�x;"|��23"�9)ۮn���{�z�wJJ�8��B�C%�A��������_N8�;�3/r�_�]�;+���J��λb��a�7�lŢ�r�@��o�ھ�2�%� �g�t)]�ȗ,���9����Z@��n��vNnұӾe�5 G��c�d�n�kJ]�l���Y޽�ilb<z��+2@Uv� �jb�[�������\Wٷp�5�,S/v��bl��X0nK�{Pu�I�;^���Xa���J�r�>��p�qT͚j�9j��Qh��z�&�Yo�b>�JQ!���WnǓ:�op���xZ�����Ӆ]Gj��d]c�11i\�$9*�n���9p龿Ofx��I�{OKֽ�c�I}Wܡ#6�3%hN�vJ8�i��w���t7�<��>`�����߫+�@��|3r8YzJ�KA�n��"��%W]��*�'�n���M+]��
ݍ��"	���f6��Ȭ��߱ohY�A�P�|���o4Qe�lS�ڼ���쨿�W�|�)ꗩ��2�¶���p촌ެ \���aoxv�TX�ؐ�㜱�Eݘx�]�c+[5��٤\y̷7l����ъ�b|_e2;Z�a���*�.�Oe��Y�y�/i�\I�����)t�t|sa]N\�6a�`Y�ռ�BQS5�V�'���� v���}�I+��l�@�Uq�{��𻧰�M9�f��J�fE����"L=�����)�����Y,\�郭����`�)4bT���0)^J���yܗ�%MW1��D������P�@-�[Y�{��J�r7�Z*.�����Wx~�B��ڌ]ȗN�ֶ��ޔqo�]���ؔ��v��^CJ^|)S޲��MF39���\#6�ӔKg���2+)��]���8�2$���b��}�M��d���(u�\1T|kc���h�q\��@N㶷��Y�[���7O*Q��Rd+5�O)5C����	�|32ѓ�b�2<}�=y��v��(�[5��K��3;��`���:ܳ^͓���w�{�g�0�7C������؀�]�����ű�%&�9R�e�G�����(���;}d��t����=�&��*�6V��]g[��E8+����3�r�v(���]mnM"A��.6;P�6̵���՘8�:�-ː�M�G����U�*,+V
�)-�,�E�ڊ�e_m��,X�1�b�¢����b�e��*�Q�c+b �R�F�-�Z��Tm����QPX"%E�@��Ȣ�)J����BT�TVEĔLAk
)b��*�.P�ZTXAAH��h�F,EV°F(�� X�eJ�ڌ�X(R�D�1�H, �ZŋY
�I��4��V)��R�"�jY+X���h#�*��ma��EX���2Ћ�Y-�UX�De��12ʢ
����*�Y�Qf���ypk��d�;^1�I�woINv(���$�/����I����zq��)t�m�t�u�W��/��]�QXNwj���}���O3A3����x��gF�]�o�����[x�U��3��,u5o3;AAq}�z�qoF6򧝛�+��ʃ���Gd�5��J\}鵦LK|�-�{��}P�Q�<�-T�<���>)o��6�c����zוvM�B6�}us���]U�(�[.2�TO�O]�k�9�9}Yr�G�ַ������V��Ug�8��:��;�M���y��{�p�X"��gQ�܊^է��XRCrT�j�⨲�^�QU��)<<�/	]���*�Ĕ�k;���p��c�םgm�mgP�++};�c��X��k޻m������r�ݼ��`�ާ��L:��D�F:N�QK��M��]�u��O]�-,�8kq�l9N�e+�`��V%�A����R��6�Ș�rrJ�*�<�]4�����|��}㽖k�G��.�K�t8�;��PɀC�sz]&�R��u��W�k��
l�1V:�q�������~���r�OZ�m�D�ʓk�Z�9>sT;�Guf����k�p��\D���Fw�OU�9���W^M�d���葲�WD���#q{��>�΄�Z|f�O���V����;�%ے�;ίxe-n��к�S;S#.���;��4�^�f��gLs.0��\�ypH�|q�O�S���ëR����=��"����̩k�������/�Mk1=ڹ�$���[|������bw;p���6���<�<��Kk��������0N��ݲ0�,��>�G����5�L�G�p:���lZұ+[<��jb�{W��]�W��;��q>���\&�t5.�9���v��MrV���i���u,T�-8���Pq�[�x
]�5�w�5S����$u|_g,]&H�~�W��ٙ╭�ҭ�����B���[�.��Բ��'����r��^7�5�bǖ�Ki����޸O��ɹ�*�qv����rcd�Z<���C֣9�*�AŤ�s�y��'����}kt��1���ʻ���-c�Z���:�I�k��]��g�a�fN������[(:+7���Z�ܸc��8ܾ���=�2r��B� �+����36��l�=�q��[�Q���V���:|��3�P��e�D+0:A�����o�X��M�jW>���!�MǛ8��qu���򾶛ܦ���ŹϹ,�*~=�dA-m��}N50�.S0��ܨ�Ս[�ք�^���o�⯕�;
��^�7]ۆ�׋�.GeOA�Z����a]��iK����gϝy����w��vݡ)%\�#gh`�p0%y%�K�Zk/M.c~����n���e'<�{���9�.#R1s�.�+��ʱ�*�*'�~������zh�m�}/��N%����V���7�[OP{x�噈W*z�0�ʯ���+^i7'b��2�-�ZT�8��0�s���;g8u�{	�W.`t.�
��Wʌ-i�H��.�f�9,S�u~9]̺�o��2���t��:��s�%P)�ڶ���Ӻ���ym�����Kj;���yI�{�
g�88	t�	�#��|zU�V�9����R��w�Bx��^X֩���މ�a�0��Rr�7oY�V���b`eP�עc&�vB��n���TN돑˃�{̫~��������+B~7�W�\�ڋ��pq�1��w��1�7�Ә%��k v���K�@��9��#22���uf*!�� ����|�������T�y	;��u������m}y���s���axo�f��is�^�]Cl�c���\F�*{���
�궼.Aq>}(�]���S��u*�Lt��wN;�=��^q�d��A��i�8��bj7g��8���V��c�(��Z��\ߣU����<;Qk
��T�T�E�9MK}�SR�R�SX9��T-���}��}�>܊y�Z�o��*��+m]���:���S��v�BxnJ�ZՎ[e��*�Jx����>���S"�������t�^�\[�GeD�3�O�k|��/iʬ��gh��m�T���+n�UZ5�@ɵ�{��Һ������l��ٽK��6\v%��q�Ӛ�9���X�6�j�ꛃ{wNZc^ӌ}K�����	=?;�4��Q�������T������g��{J��y�Y򙹓�\*<��]��;���ͯNE�8;ޖ��� �k�R�t���h��9�oK�0lR��պz���ኔ,���\���J��x[���4�)�]9vg�;B��i�o���W}זW�ꙑ8eZ��½�s����}��zOc�'a?�Ŕ�j�D����N4���gx+��R�nNn�J����C������ad�p2�2�'�p��.��v�&IU��"�ڧ�:wr�e>j�`�̻��s�̾���O�Ø��3��*��*�]\Ż�����/r�q��p�w~]�=y�ѥ�y���ŀ��ـUd ��9���eU�ʅ�'�c"�uM[��!co��|R�6��caւL���Έ1<㱟'Փ{��/Խ�O��3��I�l�T_h�:z�h�����&�Ot�	]ު+���>��W��_�8�M'�� )-Ȫ��ެ�9�Ӻ�|jj��)��v�Rz��n(��v��q�-�d��7��UԷ����7{��~����5�;X�M�rTݤ�E�i���iu�����ƞ-����XRCs�Pb���,⨲�w��஡m𘈼��w��2b��W�ċ8�ֶѕzn��XR<��Sp*�z�k'�J����y{��[
����N-���&�ag�:S�VGR]gJ�[u٭ɹ�,��|t.��s�\.t\�{qGѽ�A��@3sxf�-����+2����#聯4�sNk,f{�)e�>a�����we����u��6A�gV9Sیw��?PD��c�a��|�ϝ���;����{C��q��u��TNzJ��qw}�k��S�o"�k�u'��i=s���㸥
����Mkh��2.�I�-p�\��9+���Rcu_�Fk�+i3��.j�rWPɘ}��������	����19��w�������ƫ�*���μ�X;�wU첬��a��&"���j��үN9����w���W6ыնpͧz�|�2�Gbxe\�������x�m�GZU�~���᝾��mT*q	�u	:w�*_�rD3q?s�<,�r���<��ˊ��)���]�������jX�O�p/@�w��HG8ua�k��9���&��!F�n���Oh�z��ϗ{*��z������g��� ;�L��N>���l��5�vc&�vG)��)[{�~��l�,�j3�������ɔ��b~˲U�o�:{�K����Ȁ}^��t�rs\7�UD�j���n�B*4r�0�J� ����yl'�H�\6�	V�u��C.����j'��»��R����}��b�<�w3��
�G^Dw�|�JŴ��oϪ��v?R���+
�Up3�"e@�O���O��s��_*TqM>ſ.���]Y�Y9~t��+iB���W��-/;�NU?(6��{������Gm�ڷ�>=�\�Қm���c���e�lZn��]no��޸���~�߫;��ݡ����w��@�sч����ީ����cO�[Ыo��� �������n�`ܗ���h�J)�TY�_Yל�}�)�|�>�N`���.�0b�7bJ�f��18�%���pbR�|��e.�O��i\=v��Pҝ�#;�4�O}X��_������[l#�6�t�s}7	�)���=�7�n\��%���ӹQR�ۥ�#��ԫ��}P�ճ���+s�n�+�]�D=}�'��Ѫ�Y�h��a��wG���C=K���&�]X�Q�/��{ڐ�FАc]�|�<�{�T#�9�)���6Ǳ]�X���-�++�֞e���	,��OcUř^S}���G�D�R#�k
d9��T�@�>�Ǌm�\�K��z���B��\��=�*˜τo��w���?��'^��{սW�~��R�]Μ�;ez��^? V���E��A^���V�<Nw9DM��Qb����x{ޙ����:����J��E����h�kn�a�f8�ض��� �\��O��s�z�~��6lU	j뙉�����9��N�^�_mA����+�v1`8�w]�옮
M�[|��u�SFsVU��3�N]#G�z��O���m^c������r�y�1��z��v�i뫺ں�Й^Ss�AO�mx\(.:|��.���_P���'w{���O|�)��C�[U'����Z�cÜ��o���)E�SyE�i�n;��Z>��h���|��k�������8j�b^�^��p݊��R�R�sKHµ�n�<����un9W�nc9�xף��XUկnV�p�ބ8�}|�%�;�.o��80�N.qyTY|��{�y�F�^�)#䇼���h���Z�Ҝ�����́n�o�'_�O���l{��_,��{�c�SF��x�X��X��tU����k}���@�m҆�e_:L��e�)�$쎖�79a���-�K��ö�j��$�m`ۍ��Ư78P�Ĭ81�t�����e�߻�����կ�jg�5Q5��c� �v��D�O����%��5�g+��O8��Q��<��we&�hC�?\C��w۵r�����juցxͱ�E����]4���i\>��^�t���r��*�б�ި�&v��{.ח�Ԯ���X���Ұ�B��#�MG9R���׸j
��*��^�4�j��$�e\~5З}� ��~����֞p�U<K-����/�WZ�y��l5��\�̄����e����;�2�۷���]r����k��:�<K6��a�Wa�X��
�{�����L�s����
Fo
��>F��Љ����FhZR�>b(I��)[~h"/�kk��Uq�����a�
�����P~\��}S8n�MN���7��ڍZ���Ʃ1��o*j#���Pɞ�n:V�'깍̿`VpĈ;�I8[8^b��Y5ԱMJ��V�H�:gS T���7� ��7ص�}O��x�kl����*���pt�gW�]Q����e���͡ ���C�]eo:�qU���:����H�]�^�{#�Y�/�%���xu��}�_fho�K|�Eߋۨ��W����ޥQ��'���"�bl�iU�>&v57oڦ��8�]�o���Z{�}��p>�phc�m��e��5�i����j<�ޖ��s\5y�O �J��$.Ϭ㯱G*�K��<��fF[z�/z1@�+1�{����9��優Xڕ�����6�J�}�+-=N����UG�[ˆ��Ȧ�*��0��Ī5�jTc��J�T���Wr�׾e��_�S���z��$��E��p4,�é�y�on�!�q/(�ߗ.��C}��gJ��ܯRz�>��=�轄�هbE�6������tv�Æ�*K	p���.�I)�/���������dL�121ploz�mo��ܧ��$B�I�e��?_DWzoH8g�NŰR{jz�.�|�*�Utr�R��Q�W*c�kx�ɮV����1�����;`#ň5yS��bo�In)x�=��Nz(���N��q��4�	[��A@����.0J�;��v;�Ok�j����$yyBp�:2����>�9`x��,B��A@��򡛙s��:�%���3�j��a�I�݃���%,�����{��٩>���aXo2�/˝�����Z�s��^�`�n��嗺h⸶N�ѹ�d�O��1�so��ڀ�!,����2N�Z�KW�Zα���lTNl�g�X$�7����ݵN"��K��|����v����fPVs�PhWKT��l���,>���0{�.�~z���4��(�h�5X"ԲK:);�U]at���uf�v������MgU�F���FГ5��2 "j��٦j��\ë�vv��F�f}���P:�<�1B;�����Z,�d�sؙ�J�Vy��p{�m�띪�����m�y��`�����.T�<�9���!�.�^ҍ���q���p���k?{��[�/!Uݽ����Όn0uNz�rޗW�&,���4og5k�5�Ǣ��؀�F{˺��F�MnN�-���l��L��`��Ŕtӈ��#��tm8M�}A���Y��,��nѳ͛H��$+g���梔����[r���}�\��K���gLOe�Rnf���1I\�v0l}CV�= ���/�v��K��F��|]��y�pހ��n�>��[���j�z�w@LK�nˍ���z�:�匷�x&錁5�Q�6Fm�R�.;�R���61Ұ�Xh
nl�),w�h#SP#�s5�uJ�Բ"�����aC�e�Z�MA��L�;��y��yh�T�ބb�i�_bDP՜ر*��Ojn�Cծ����;{X���J�gy�����K�Ooq����	�\�8�V
��g��I��J�>��� �L��L�M��GV��2��h���6Fp���"���{�O��4�@��ר,B���.���ܙ|ER�v����l�9�h���J	����h�[�2����)6�A�@��l��J�ט�gg��玙5�1��W���`#��EYm�t^uu���d��sJf�܊¢j�ܙƚ�������b�*<��եF��gP�l�ٱ����om%�'챎�#5{C�܆�V����h1w��<��&ȐVXd�-�Ci�:7'K�$��tŸ|�Y�\A�Aາ�x�R)3�ӎ݊��IĹպ�J)��,���^�*c]���ǝ��#Q��Qv���2�.�ή]����>��-�7'>޺S4�����.b�q����C��[����v4�����ځҝʔ�]>��n�ņP��^�k\ft��f�|JU������;?r�Z2�<%��1��[^��l�`	CU��`���ө�
��Z��7I���I��	ƺ]L�a�U��w�Օ�Z�ւł��X�.ZE���(�Y̦ZVUAJ�X,Q�ڢ0����F�F\�r$Zŕ����EQE�h�2�Ҧ$��q���J�[d[��pkX
T��T�VT�b�
�B�)meE�#J)�U�*#j��*YiFAVTU�(,��j0�b�)Z(�X�i�T�T�̭�Fҕ*6�UT(��k
��YQ�q�ehVG��m��V��ekm-��r���ckh���hE�5���
+-���h�5+[i[K+�W*��Y,�mV�+X��b�0D��1,a��(-aQiKR*YAdE�\Ÿ��c�(QT���ij��kR��*�ժ���QDZ�V	iEjV*[
��6�\feh��m��cV�[emp�ܸ�	w��{��_H2�M.&;P+�"�`�y�)n�κ���\Й��+nr���ͨ��7�Z<�={ʯG���>j��
�O�I&�SC9�r�o��+��*�47�����V
O�	��kZX�)��{ۻc�{��IӸ�`����޾[V
�����v6�͞�[](Wr����/c~R`��C�MCYۤx�k���Ww9Mnr\D�Kn����Qx��h8�r�w������7�N^�;%o-�8����0A��Uô=Qm�h�v�X�y��;�UĶN/s5dJ.o��q�q��7K)��a�Kg��ڡ�B���K���A��C�nVc�z�oga�Y��Sޖ�����y<CO��*�B���-u�yn1 ���ⷙ����rOk�c??17��wM��LK�;RU�mO_�����Bf��}��{�zw�UI�[֞��|X<δ��9��/�|��x��r���P�:�sί}�zϜ�}����w8����e���4�Pb��{D�mX��e�������ٲ�/�M�}5س�[��݃�}ݳU���u�a��)�,K m���/����d��0I�e$��n���Rb�{=�H�;ݞX�j6ͽ��c���͑od\���<��g�Y�Y���}�ي��:�]_��Z�+N�aQr�M>K
�O���ZO8E��<����(��������YJ�U:;*${>���{�]��Z7B�g�^6�y�վ��R�@x�X��|#�T��}n�j�jY��I ����;����2�Z���^hY�uf���P�[����{�.�T,���%��Zު�����y���.�p����O!w�0����l>%{�3IL�ː�����*cU��}���j��}��˳��d��]ǒ[�Bq{��Eg�A]�i�}n��2����=�c��뿖s!W
�ג�����\�1'/�4�����ܿ��(�������)r��̳�r��A+痣����5Xy�\������}�v������	��9j�ƻ�".+��t���u��C�!�T�'�+\ʏ!���;����76����j��o,TF/�{�e��V�ב����6��Y�D��2����p\�ö��3٪�;]4�͵[�7w����$��ot��'a0��T��m��gHy�{���L����nX E��YT�,�G7�^H�AS6Ç�<7����F���X�}�}{R�kKs�_oY�3���G��Y���Q���[�7�bߔ���7:�I��3��q��<���Z2./w���m	�I+|�:��E���Q�C��J�$��6yG��.э�I�H��W�=�8�3@�{��g"��ꝴ�-����M�E�>��_=��9Lk��N.�,��p�jY�l7��J��TY�V_=Er�_i��._\��ħO67 G���^�� e�7�}Jx�_�P�B�lQ�{v�����R�'&n_>�h��s�97�U�W�ඖ�U��쯤���;1!WG.��z���}��q��=;4���ۇ�&!:n�c�cR���-L����c��Z�N-�����N&�<J隻�|S�������꧳�|��Œr�5��T�Lpj�G<���B�vJ�ӛ�v?x�'ql��Χա7��K��tӄ��E8��1�9���0�k�����d*Ϸ�s�vʗ$��%�Һd��Vۆǖ�cwAG��90�r�K�凹�vm�w7F�ZQ�y���w�	�y4�Ay[Xn�wvv��~��z�Θ�D�����	iO%0��=�bh�W�Ih��֮]ѓ{��^ŧ�N|R$�H/p5=[
���U�x\]��l9����J
��9y�Ӫ>��suÝ�����o*�7��hT��]���f�U�$u/qN���{'��u��ՌNeI�֩�M@�jq�6D��E��Y(���9������ݣ�F�w��<����F�[y	IqQ���yS\���@�ޖ�Bn=�;��O����[lߣ���r��<;�j��J7�=�x!��mC�,�/Î���D���r������4�n������Z�Ϋ�mx6������^@����ݵ:5���k8���D/b�Q%P�X�t�Z�WZ�[lW֓��y��-ׇ�-aHU�Pb��:g�Ko��l^<��N8���*����k�n�����D�ǲ�df��SՕT塋��Z�a�n�McN�'�l�W�<z;3�{PU򎲳��D��n�P�]JGu������I��b�����;�Rԉ��\�����9�`�U8��w��Y�m6����5ЧYȞ1lsPwÞ'�9҄�m�&Lx]�^�Tb�:9k<������5�)<FT�j�V�q�'�����.�����-��sSx�z��RҸ����:{j���]^�˝�Z�JS���ΝwB���y6�sy��=7O����KEk�N��áFr[��zKY^;ٵ]��N����P��b��s�f-��Ck���=�R��=���Ծ:ϕ�:B���y\Jו:�<�]b����53Le�'͞���s7r:��?B�s�v�Y�ٴ��:�߅���{k_wf�2k��݇Y�E$��9P��'��c��<S�&�]��#�ө�Y8}CymQI����?��I����~�uy������3e�p��Fb�.��PD8����:�E+ȼ�W�uh9��UN��Q�Z���2��;����~�'d���zF|���b�w��h.'ǟ�b]��n����QnĒװ��V���Ӯ/ZOs&�Õ��|\vTWQj��<��Vy��OpU��ٍ��8��0�+����'m��Ǡh*c���mJ�B7u����'�q����?R�6��3�7Z�ݺ�������:Ӫ�u�}��m[Z�����z��7Q�u}�ScD���ɱDwe��J]ْNgfs�0*g�)e_��g��������A��������8�'e��������=,��!�>ly5�r�w����c/�M�����㣙�5�/�p�g�Y���g/�^�#ӏڧkS{���M��]ّ�تl�pFd���kS(�?��w���e�Uew�><�|����їEW=,�vʝE�8����,/S���%A����%�+�#S�~�8M�z�����3&�F��}�������\�L�Ճ��#�3� PYu������:]o�م�7{��g�M*��w���wIU�[*0%�Օ��ڬj�H�_5C���`����.������<��U,ʹS����ˌ���!��׻#�Mr�T�خ����I0Ԟk�'p�����9�b�`�	����87h��CbV��b{�\�s-���|ʇ�ϳY=7��w�ِ�qxF��K!Ʀӗ'�����=��Dݷ����q�q��E� ��Ҟ��4ő�F�`��;���%ٝ����r����RYˮND3[Օ��2L�&� ���6'Vn��N��S d��->�o���]h^�h{�ɘ3j�u^�Ѭ���Y�#��K���yau�-�+�,ȫ�Ar�?�)&�.
Ę­T���c����⃮N�"y���>�L��]�ዕ���z�z`B��{��[���m)@�nq�Fr=�K<|�ﶨ��`�k�������1=���/�;�R�q�t���=�P�\Ƹ��,0�%���w3��Z�&�qy9_c�o�}�I��s��6���� �pU�۔�i��$��V�E�W78�-�Wأ}�/.7Rme�ڭ"d��K1��r�eVt�������mϧ���*��;q���Ȼ��	.�ۥ]����`z�����˙��$]c��Y�>���'i���T!�M׋����p{��6���5��-�W�`Y���QןJ�;+~���Xx�۽�ӧ��Kw�<鵩�5��wm�oB�㬬�*Gd�d.0mn�\(�y�"k�=Mu�r�g2��h�(���>?K�T	]�䵞O"no��#/f�y��BIn��ͧ6���V��5�{���{$��C�������Q��f�"���~���V�:@��yo��z!l{(�{��%�wd-
��R�8�WI*�v=m��Ҟ�M+��K�v��[�z�t;�o��f�syQ�Z��eI��VD��.���hw�5�R���aխk���j�3�r�s<�l�8�E��U5eW�3>���o�T���oc�����z2j�8m㞋�֜u�n	���B���C^�OA]�pw��P��SN��^�Ж��S�]O����{���&n!NGRy
O-�ܟQ�o�UOl��5�\�צb����uq��a���r�13�'�ݩ�hT\rxg�����"�,��L�[�ֻ��{=Y�����8���5Ht����S���5��g\t`��9�(�i��<�-��败4�=��cPs}�ۅ�ы��I=
b���կ3�y�}��@G������8�����Oƨ1�J7�=m�ܦ�/����k��y,ٱ]�6��-��4=EZ�TqM>���{_�&�g�y�a㸓���֬����:aӷ�ʗK1ngD�ʰ�@�kQ�m���w�
�f�Q��=�	��� v�5BV�`�x���F�-�U�}�u�]�G�O_����6Q��@o8V���q1�.֓�,)"���")/_0���z�6��}���Ӛ��/��Ud\⨳�&�پB���s�����5&&\F��ب����'��\ߐ��I��{�C{�;:q{�pDż���v�Y��E<0�;���7�+��}obQ�.n���خ����L�r��-�w%ѓξޥ�q)��;�{B��<�dԖ��]��Q��(�}���Ge}*�]�M���"��pJ��]�����2h�Zy6���ԝ�XZ���d=��
�\��|ﴖ�=YJRYo������#7�-g?�YuJj9ʗcU9eOL��� .�#��P�cz��rU�v������&5<�
���a��&�<��+Z�̩����iV���;s.���͖���d*�o���/�ЖԌO���u]SX���]��-{�ud�'�a_t��$��̨})�t��Jqe�k9����1������Ҋ�����{�r��:�|�#/�|zޖ��0�W��TZ/����'��P4v��wD�+oumN�Q��.�k��C��û]�� ��#�"k��g	1j��,���C�i_}r��Q��ڃ�^=����EX�Z�ry����5x��7�vP��w&/����G�1����'Rh�{���c� ��ݭ=���-c�wu�¢���.m�5��ߊ\W���.�WӉ�W��';;"Y嫹9�2��y�m|�S��l�}�]Aqٿ|����y�]��ȭ�����٢�ibs�/{|�n����'v���]�▮o�(){��)����R���UE՛<��Uw�~05��_�K'#hPN»�Չ@�܆[���gF8�Z^V�B�҇��7�_5�X��'=3�[�J�f�y�2��L݇_N���:��*��_ڧj57��>�oj��QѸ�����K�ʗ�1	U��QN�VyU��U,	�:�ߪO>�K)%�Z����O�S��cB�LOQQ�R��Q4�,+���:�V-̋�Y�/��a�n�a�!�[��mAv���)X���ʉ.J\7�~�H�淬õ�%]��-n%�C/��Q!�Ҏ�rS;6��S��i�HZ�Q�n��Z]��A���9iqUp�ݵn�P@f�o�U,�溔|��lm�֬3_x8c�Z+;fF�S�f+ ,LuΡI��"<�yG������(�]�����YX�Kx~��<�l{�o���җ��P����Ǵ�����~�S���>��+5��9s��f��'ɝ��`԰n�7m�{�	˲� 9���� w:�p�طAkd�?*�;wV2A-������ȯVv��۵}VbT�m���(�W��J�k�� h�t�k��l�
�ҝ�bx��T2ݣ�Z�G�t�5�;�^旑"�)0t�M��e���Uՠ%s�)]l����	Nt�����h=��8N�Χ��N:+��Ȣ+�[�n�~��������GB�p�<xø�;-���:eJ�,%K0���ap��%KG�^�Ck��G�0_Zwc&�ٰ�ߋ�gbhg	��]<'�{L3�}ٝ���yڕOf�
���y԰�Oܸ�nV�"]d�M�>�+l	K/-wP�y��Z-�=�}�b^f�ͼ�a}��a��m�M����9v��`��DhJ������d��{Y�BE���1[����}��E��ꖌ���w�� ڍ���g2�W7}HN������Nf��;�Rs��ҕN�����J{����5S�>�=�l[��G����זԼ�S���.d��/�\�ێVv���c��\Z�.�����9�d�a���^�[nw����dhʵ��1 %��������%ػR����@$��.��U�\03o��̓v]a����v��[����� �@�M<'�)�1��zd�����P��8��*��b�7���+J�}Ff��n3	����8��*��c���a���vc��^�VQ� ��2�Cf7C,�n-)��v�z�8FO�3H�k�P�:���!DZK0c�ȼ0hX.�;���P��ui�c�zp;6dF�w� �&�\��/�4x�����B������WD�¤ܠ%�9s/]�&���srfҧ¯� �@�������W*�k�<�]p���9E�_iecG��I7F�6R92�'xC��)�:�w��o�tT}=&[���gV�k,��;�/.��7���Zg$/%���{S�!���U�x������`v
Ӯ���<szA��M0���Ǖa�c����w���[ i�{��+��e��W}��U�B���N��v���萴%���ꩭ��1����z.�6��y=�]��>s���{�)u��.9�e��X��}�=k�n=���t^�z3޽�iK!�ˇW��0���]9��9�b+��SM�cmH]��W[�`0R�B*����;�<��2�ƅ�)�v�)<l�]�Pе��X^u+&�4�i����q��h�+8A�j.��G�����&N
νne��fv� /��z�s�,׿u��a7���ϵ���������*Q��+)V���e���A�iR��[h&Zܹ�\��)��Y*��������j�EEUdRإ
�ư����R�b��L�ʪ�jұceE�ZT�EKKZ)lKkj**�������32eT(��*�J�*�k2�b�%�#[��*.��E`�l˙Q���eE[n4XřJ(�E���A�Tʖ�%hƴJ�QDe�[m��X)�����X�iiG�Q��
#Z*���i\LqQ�Vj��ĦP�UE%�9LC+E�V�����A�+
��V�Z��h�)X�c��Z0���(*�[X�R��DR����QU�UKV,m��e�m��)m�� �Ɖej�T��mZ0,U�UB����Q+m�QV,m
�U�TbV�m����¶6�F*�A�Uk(ʅDJ���J��,���2��+D�V[cQ�US-1
���i`کl��,�(5(�E�-)X�u�yz���qJ��l۰�dQ�Q�ȬA�N�g�w���wm�!iX5���nQqm�)�'G��	u�L�8�V�Ju>V�s��k��J�Jތw)l���	LԜOP��G!�].[��KV��w�J�M.�PV�N�$�j��Y��Z�|%*=\<f�q��|(6���Okˀ�2�'1˹�T���8uBn�{�/X�b���v��4��0:7lB�A�ܚ�Ovg�̺o����r�9Ԋ剐�=�ʋO휎���WNx�: ���������q���~�̳$���|��S�;�T[J�m��dsee�}��^Z߯�u}�Wg�3���X�EA��	ݻ��!����s��5Q�Ж_��l﷏E����3PQ�8Ɋ�vNWؐ3�(1�M�8�_G>ۛw�Z�nE̕�aS5�.��V*��e��ד��K��-�_O/u��O�&HH�!K'��j��y�<�è�j��.�>{�.���W�wY�䏭V��&��'���Tj��t��f��.6�ʵg��-h�U˲I��q���AY�}�tT�!5?�8��C��]]f�:κe��o�m#��sN��]��R ��ɗH����(�*İ�J����m�˺�u�����op@..��Ik�%4�up�/�c���f�|���9��Y<zVE�v�F��T��En�F7�[��U5��y�܈�s_+�z{��BUA�R�������v��Uwٯ����hN�O�>������k�<26Ԩ��s�-�l�"ES����z�n���Ou��>�	m�{G���RZ��[c�����SJ�༺nVo���^�܍.���4ҷûn��N��=���]�}X��
��k�t<�='�]���3���_'�P��
�:�\el�y���<�ܶx�P����`-wٗ}쪝 '3R����慄nJ�'�^�}[9���*Z�{z�m����}}�9/�-A��VA�|����c�ەq�j���|��+�y �d�TA��Õ3��k6:�7/5�>V�p������&*�P���#qΜ��G�r��i��0Kޭ:7AC�纶�BT��7��\p|�
QLO0��~�qe���:�,V
��7.`"�*�K���O����u3�Sk9��L/h�t��*�4���-��+�\�9/z�Vp��K�ZS\�1�ɖ{bıƬuoL�<��*�U&�m"�"�E���������ήS�QS8��ו��n�~�7���RTR���o�{RS^�}�ި��y�Ao��w���j����X��y���
�z�v��5��=SǢ���r�Y%=�6�,����e�����������&@�#��s�C�����y��8��𽪜�dy+���Q��7,�4�٫5�S�֪�W���vB����vB����O��w�N�u�y����R.T�=0���9���r��{5�z����ф�=�-�d5�}��s�:��^F������|aGi����^�x����Ҝ��1��ޕ7�R~��@��)��U�]pc�_�F��;�������'F�O	��SR3�;>�G_�\��-�������
�ԯY��4m��=ґ��O��M�\��}�ʲ�{Q�|����W��,�e8%��% �n"����-nF�4r���(EC�{�񱋶���8#"���]S��>���ފ%�����|�0�X�ymA��4�tt�=gY�*�o.r�3D3r�w*�[�d��l�|���׶(]��w_��c��w7XfW6xZ��|q��F�KG!Qp7vR�\��'��쇓&�O��W�q{�Y^;Ӣ��e��p�U�/��3�J�W�ϑ����>�K�ػ��uJ0�h�E{��Q~J�K�����'��:W��rL� lB�2�&&�yd�-�v2�o����>�;�FA�Zw 2�z��G���c�%ze/]p�Q�&�D��I��I��vG�͚�Y�LLRU�u���M1���K�|z���qT�y��L%�@Yڇ��(�*��	>�3�0L�G6"r��FV�g����^�U�xh���L_�ꏈ͎�,�q���v��c��5CY���)z$��>��g��n�;ͯq�/��ڇ�Jh�t�$J��˗+�;�~���U>"�xj7���q�.f��z$�����Zoz��~�~4���O���u���~���.��>yN�ڜ�x���G���ݸ���nt��{G�Js��C�]����0V���a�����x�X/�����G�/:�ޞ�|��:�}�<b״�q��7�Ջ��g�d�v�3R�V<0��~�&����=�wR=��m�H����#��]������S�~���o�:������R�_vf�7\ўR��br8��y��d��7M?	.g6����z�j�I�u_<�t��f�8׷�t)�^n��nf;�ub�A+��s*y{n8���"�ս;X�F�]mv�}���Fy]��u�X6�|���µ.�+�F=�-5���O]T{Ƣ1]1dγy3��u:1��^ң|�����U��[�u�I�ǔf2�5e�C�9DcH�A�٨`LEw��L�d��9�C8_ow��=��$�^��fI���-�t�}/���[R�c�L��,	��\�9u��I~R3�ez��L�>�t}��Egʽm���7����sվ�+�e� &h��T�oF�f��x���}���������9���h�^��>:���tײ�����2�l��{��u>�[��9O\z�g��� 4]���^9�>
��Bo���cb��s�#��{'.(,��tj���%���/�8O���m�R&&)�{N���ǩ:H�zT׊�N�Y�7��W��7w��Or�`��۹=��*+��L��߁���VѸ��{�ó�B^5�^����3�����{�d�t�5׬=>� ;���R'f|Y�u�m�/ղkK��=) :��N_��5��F�)>��5~��ٿ���rUh�3��^>��ׂ㓓�o_XS
�����%��Ƃ�H���×�X��:*�*Ǯ�zI2�H�P^��;F]���c|��{�2�b�+��f�_Ǎ2�E|������ǏBS�Z�a�_Ѽ=���kc�{��IT��Ro�i>1׻�Tq��HTQ��Qq�{Ϲ�ӻ$c�~y-��/%��M~?On�L\o�x�o�w��띳�[+�S�Ǻ;�RV]*_�78�r!��}��]��7��5���^���u���g�D{��S�T�8����hS���^d5(���Ȉ�9$��D�Cˌ�ŋ�3f�޹}q����x��^�r;��փg���QY�/Gv�ܞ�	��kG��iqQ'pꙇgr���}���F�]�H�����'�	�ҟ�����i%�ǚ�;�J�+^�C�}ߴ���x��V,����J�����a���X7�g�]~�-<��[���?_���T��߽Q�kͻ�w��#]N�������W���9�$���'�3�l�[��ۘ��gZ����w�״�����ߧȗj�5��ed{�
f�� -��n��M�����^�������=�U��>�vK�z�?}O�ё�
��'J�z���]R�w�{�����U�y�Z�p�Y��;o�
�e���¼^�ڭ���CB��1q�=ǽ�FH�s��j�x��N�\OQv�v�g�N�Q끲|���j�!R�KA-fmCU�#"�%��'�N����r�)E���#����a�;,��2]�����s��Fv\��ji������b['T�bV�35�X�O�:���]�����mL3ʰ�F���O��j����Ln�:.mz���j�:��e����挞�������t���<�;�o��N+�W%q'`�Ds�8{)�~�MÍ'�T{7JhQ}^Ä�wr��~�{�nSQ]�6<�;¯M�W�};��7S��~� ;�n܊yT��>/��>Q���=�gzd�\vY���K���bo���'��'�Q��Lۙ�>����W�`S̯QG"T4{>��73�v��Wg�~\�F��k���^���+�o>X�˝yd�C��OM��������EѪ��Yo�����zK<��A~�יZؗ(t��s���ߒ�����~tMǜ��yj�0n+3N��b=<�r2�q�&{�_VM�2��^)�����n� Oܯ��sws��	]靪�]#Y묥�q3�~����i�g�#�q��� W��'��c���]ٮ@Wv�`�f�/�{�\��=*�v��g]��Mh�^ڞ=�O��t�{�V�+���=R�4����~�e�S�ڔ6����o�W7�3��\w�֢���o�tqLd�"G�r�����^|3��8׶etƲ�q��~�y�~=�oӼ_��oG{�Q�s�[;۞��ǔm��d�{�#�v�����F��>���]_=;_|�<+|$�;-/�߃�9���3�$���B�{-���.������%C�^��>h�<���Y�'1c��/�軬."�A�KO{}֧�����6�/1ާ[2V�='���v�T��^��&.|��;�q�>E�r���'>㾹��~�p���)�9���X^.�^6a����M����� T_�2�j�z��Ō�~��V��{5��P�`8S[�%��}��.�Zg��?
��% ��j	�n��R�]dF�4j-��<z�2=�q@}��Y��d̟b>m
�k{և�W���˦^���P�����@�KG��:�f$ٍ�]r㾖�ϣd�1�q7/֑��(�9���N�����p6Hl��m*�1�.,�nnS�;OK��Q�7��#�Ī6����#�9ģ���dF���\�)xO�g���ʒh{�n���[T��#ѹ���f�y�\�;�߹z��G���c#Ӵ�3�9s��L��	�J���o�}�'�@�ӱ>�웨[��cb���k��,^�J��5�~�Cޓv63��T{���|�X�~�ˀ*#�zf�92���n���V�y��:�Wuxh���W��~�&
ů݋�ͭ˳�پ�Ͻ5C|s�:h��%>��l{�{^O?1 �2�d�������=��������ł�ͬ�V#C�u��b� :�!J����rw�˻!��9S_���Y��&ﲻ3������Ϊ/�][����hp׻��/W}!�X�����q#��/-H��F��1k6o��5�;OC3��Y��I����^��FzP:i��ǳ�t���Q˟PM��g�C���S�����i��*���>E�雎>~Y~��D'5� w��+ݻqW�s�����q���b�����dl�JK�A����5���B���F�x03V��j}��������*����V��~"
�5��们���zFs(^��ZX���� k��ێ�l�cu�=����&��w�}�M�g�u�.�B�VY�`~��b�Ǧ�9'0�����X�����o��O#�ю�~�q���DH���y@��}xs�n�E<�4t{��Y�Ӓ(%;5	��ø�2���ax�pC�EoNӽ���ɷ�~Ӟ)��~�+�d�,�C�N��l��M��WJ�oc=�yx-�_Oi���}P������,���/���=~VԲ� l�����$����
w;���U�蜭�n2x6w>�aU�X��~�x�޾G�Y�v�{%��j-�b��ƺ�7h��D>>�0tn�R�PO�XC+���s�j՚1.����\�{��i�p�a�V�z��nb��\+ʽ�N1SUk�td�YPݗK<M��VVZ��]<v�)��S�*�wwZ4� r�	��t@��v�3����SvR�8�`��6����|�Q����%���ю�Vev��Wkb�v�r��R�1H˔/3Ev����st4����u�LGr5���D6*�14��� ���@�=I�G�"=^w�OM-#Ǭ��bu>9�*��u��){^X�#}u�=A�숙�������a�����`@���~�}���1��V�}�t�G�k@
��l
���I��[�gq�C���l��f��zH��MN��Ht��Ѫ>�>��Fa��նo��`R-L���{kI�|K�7^	g�9z�({����}��n�{��N���,i���>��,̇�ꏦ7�$�����y������z}���ޥ��f����KTO�<7ѓ�}q���������ǆ��/d���o�]x/��K�5���g��8���f<���q"�͝�yq��,\f�i�� o���?,�d�������p;�J���|�q�ǿo�$\o�֋_�l�Ve��}�^CV��_�j����}��$�~��O(��'n���}@П4��R���:CE�M��n�gng������<'}9"�KBg�J5g�������(���~ӛ�~+�����]���yk�)�����0��K9������6��ӫ)@�b�.H;&�z�K"�j��G�$�J#�Z��V��9,&#�S���M�9�}m�Y��g���E��b�ɜ;&\��|jY8;�k���T��q�P�Zl'����oi�Yr�g9�Ň�K{Qe��'d˥G�ڇ>3X�3�g:T֩��\�lvHY8^ޡ��lK�7k���a��0�������#��:�Y���c�qp��������9gjFB���s��:�p�׷������iQ���%�]O���� k�͉FX8��B�Y��L-�u�d���eǒѤ�;�oe�kwyi#}M꠺{��|�ɋ���b�Q�eңa���si5��Y�xy[�s�>4�v��)�$3z�Q}���&�ymJQ�<Z��0aO��^e�h\�*��lm����q@�����r��t}��BӬ홸>�'���\��� Y̆ �^p��l�9��;��$ܧq
а�������ks��5Q� j�py���`�CC�{�؄	̪]Ƿ(.�F���js�Ie���{�Ɋ�e:"�����G,#����M�j����\�I�*�Vc��k3<�F���r]Û�I=���"��p�؊���ݝ+U�ɹv!���ba��ِ���V��'oB���L�]��`�����>¹[�LO!v��%�B��M�V�w��i�<��;X����f�74^[��e��Tin�ʹ�5��Dq5��Cxd����L|w9�	¶�]�?��f��u'X����)
C>BKWΧB.��C7�+�s��U�Sv��i�%�4��7m)�{�fޜ�d��T�أ�xXq��[������l��u�������L���ԉ�{�>Ļ�ǫ ��J���p�;���fZ��P�rgk�M��F�M�%��3��&ƽ�q5GW�:�>�c1p��c�ݵu�p`�qB�z�閨vS�0u�Q����E��
�VV彨����a� [F$z��P�j�Э�Ԥ9�j��Ӏ�;9�)_-�o��\��L����	Zp\|J��ܵ�;�����z[og:Y�&�]��x��Vi�uٍw]I7�b��-�W()!(��P�/� ۞���a�i�&���DiB��X,�]�P`�Y���6EJ
��!����Wy����1���__v2pc�S��e���.{��w�r��z��k�i�hM��ـ��ng�ƾ5kkw~&�J+1�,����W:�
��P<���9v&<yX�`�:�ro	���ym!j����U�#\#7Y�	���ⳍ�Ã;J�DE�rKyd��k��e.��zY�/���xz�ٶP��={��!X�#x�CIcثx62t�� o�X�"+�f��ŵ��P��6)!y�#</"3
��XN���03���,��vS�P;�����u�w��`���eAdr�h��"�Z[[[T�(�EH���PP`��h��XV�b�E�Z5YkB�����ʬ��F6����b�(�T*�U��PjQAj"EU��PJэ�H����VҊ��J���+
�eF�����aQ�-�6�AUiiEm���TP�Teb���a���8�.dr��V¤U����i�*UX���X��V��eh�U��b���jʂ��U
�A(1�Uk�e�UDj�J��,F,E1���UEq3(�؊�ih1V�m��h�DDT�P+DT�eQ����VQV�Eq�E�hT[mJ¤��mj,Q��֖ڂ++DV։ie��Pb���*TEZ��T�+P�U�%Ɗ�(� �h�m�(�(�U�ˊ媨�@[iF�)bB��b��b)*TDE�0Q�)idXZYR���-�>��0GMvM��x����b��ص_*]�����I�f<_v#h3:��*�e0)��T���Y��m��m���/�j\�pr�%�V���g��/���8�������i�O�U�cTY������Ｎ�P�ެ=o=§�M�� ���"�G̨��c��RaO�ў�q�~�q���<��ΫI�n^{�^c���Z�U���˅+!mT�S-�N��F�
�?b2�1{���!�'�Bq�6���G�BY]pǌ�u��Al��O@n�!Q+԰���f�5n�2:]���F�S��^�*.��O�wmx��#���P؇���8�|�{7JhT��9�w]�lq�T�-��\yaS^�'ѭ���+Y�;<
�����ݹ�#az����j��*w(߬{�z���j�5^{�����8J�_rf������|N3�+�[@'�5�W�I30�ة�%jl�3��yF�sۍE\/1ކ�U��"��^��J�ö���/��9�9��NAr}�p�;�=ۏ��{ʍ��MΣ��oٷ��O�I��:�턪�s��� ��{<�@P�L����R� �z��9r�8��O���OT{o���k�o����F� Lr�_��b�ݾ�+>�#.��k�S�.OL�C�R'
�z��v����fBq	x,3�Z�n��J-z�`�����܍vd��W������│@g70<4Z�P!MA˻�>ǱM�Rp�i�mV�����3j9����*�1)F�əI�%wnΤ���#Ԟ�_������٩��@�~���c�xs�0�&p�/ǥ�[t<a�ķ;�\7����Pљ����e�����Q��q�i��SǏ�ñ;,e�V�)~؞O0J�3����Z�S���zn8��k�+�N�ǫa�㑵�W{��p����O�����]��}��r�~��u�g��/��o��+ʟ�q�:�C�+��ڔo�`X��33Jr����⻗�M����>��@Y�|7��p�"�G:��x�������^F}�w��y��h��)P�p�(�y�U2EqS�L
<�~��϶����2:i�4u��Z=UUj}Y��^��z�y�xuʤ<,�.��?Q�͒�[q5�7@Z+��L>=�lb� �Ofzuѵ����9��K��F����a[Rˍ%�D��ё��[��j-ג>7����\��X�yѮ��޸�9�Lg|�Is�<�Ǽ'E}~�^�s.O�I�0[;sg����qʽޣ�X���ǧt����Fϼm�Q%�{�{�Z�g�N���r*U: Nݣ�WW ��^����PG-d22&޲j?�u���r�ם:O����X��=NrO��3t��"���77	
�X'��l:���~��B<}�=�\�������ѝpN�P���}n��b�.=be�w��M6xj�(�z���s���6�������n�����u�=]}�^�J�n��2�x�=��������;����W�o�����S�&ll��ΐk�����F�$
py51�ܯSU�u���T%W%�o�~>uk��U���О[��X[���9�GT��� ȅ���"���dM�=���0���{K����Цcު�}7NM]���{3A.Ǣ+����	�$?�϶l��rQ˟W��8=���ڇ�>ӷ�C��0��3�*��A&vc8�����ƪ��\o����n����Ḏ�IG��bvX�W�Uؙ��I02}��|�V�߸^��-�Ѐ���G�9��:�{���D��Tp��{H��.$��t}g2}��j�\�<�Ry5��K��\���`f�-y��^�O�?W#w�\M���±�^�e��,��+�F;0���R0�ʦ2�kK�L��5�͎����^��˦�iO^��;}��3�?O�3÷��L�n�l�IXOL���WL\dγ��&��F���X���v��R^]�j�ۧ�ޯ#�~�q/-�eZ�Ӓ(%;5	��\;�)�/�]�uw�Fk��l��ڐv�E1 �ňy̆�®��ѥz3�7Ȯ���җ^j��DJ��j\7��M�m��r����c79Ιd��onۙ������ya�I�L�Y�{uh*dNQ��h^�&Wr����6�n�j����L�
Ϛʆ��{J�+ǻ>�[/�eIg_��N�f���8K�M��=�B;��S��vN��l��<��<��6r=�Y�9�|n}�������6Hl��W�����W)S��s�U#*]s&�'���F�
�ھi��0�î�Ѹ}�w���[��Ws�6|}]�iZ�]��Z7�ْ,���C+���>
��Bo�u�(?d��f&�c#oכ�R��y�,�[�^��iV^�[�k��>e|`����D������Z���Rt��6�f|�=�^m���5C$���6v�
�^� =��)�zn�*�S�2�__�����7���.^���D�_Q�kR(�pq�}��.=�^6���!Mh_����=r�����[�p1��m�+�_�鉊���*���\�S�41��ⴥFa�s��7΀�9��{>gh
^�K�ɺ�\Vf�O�m6�w�ew�{��U���;�5��&N�=�n���n�}1q�'Q����g*l�\ZT�HDmzo�u�Z���?���=���vl��d�7��3_m09W�<7�u��ަT���p��^M�������]R�(��J'��D�ؠ����,����kщ
���K�2S�s�d�f�8j��:j�b�s[ݫRS7��1��2�"�<��H(�p�85cյ��a���x'ݰ�%˗�j�o�������7Х���\���)�&��Tf�~���g���s�o�%���yy^���l֛�r����-��@k������ f'�^���*S3��O����s�8^�Mh�^�]�'�0�Ȋ�xk+j����7�n�v�U��3�C�w�װH~�=�Ѷs��_k�hp��B�ǵ,�}3�L�=�b��K���i�t�=���Y��w>�vG��͎~�i��*~-w��E�x.RQW�:"�4=Md�o$�P==���s䏨ͨ�}�>s��^9惿�����z_�Go��K�Q��]r���WUѨ�-f�p�|���v@[U &��-�mK���c����Ͻ
V����#�^�����#:��)em8�����q.�A�+��ꉖ�{�<���W	~v�%Ѽ~��o=����U�!�=�]Dm}�_�<0���<��nn	P̐�J�,9KGٟF�5�����g�w)��[
U�����#��]��~>�@���?{ٞ�嚏\��7� 7�qJhQ}^�3�_H =���hH%��5~�1�iy+�s�����@��ۑ_<�tE���D���/Gv{��0Ypb%�f�i�.�2t���p��bALڌ~�.Ot��εWf�8;vM%Ԁm�91Zx�uJ V��N��A��]G2ZM�����4���w���3��F�nb�^�e�侁�GY�-���y����(�4^\2e�:�g�2�sZ��;������t��^^3���ߎo���I����΀���˪"�3��Fm���4L�C��#��9蛦6��D*���EF�wǰ���P۟�)ϡ��E��׍��^����d+���'���Mϑ��r���n�y>&�΃;�ǹM�G:�^���긘����ɣS�\�#�����*Y���=1��0�ٵ�7ޞj6��ai�!m�`��iY����T|E���O{�T(l/i�~�#Y�o�8�����mx���W�������q����ݹ���E���3^��и~�Z-?u�+~�gFi��c6�W�3�>���y��ý9���nӳ�����>����
��|z���F׵\M�獧�#����ڠ��6��s{}*�H�p+�\2�ɭ*�&u�_��'<�lG?_�[�ң�x�C�wg-!iK�i�.�ŉzY���>g''눪`M�x�q3���3�_9���q�x�Ͻ�^G��j9���	y��N��ҧRCq~<?bL��>��n$�*n��5<�~���L�z�f��	��ϲ����7Y=�c� T�������p^��_���޽0s���m�ˎ�aN������0�}���Px�ܤ[I./30�l�Z]Ã����t!�����9;��4���s�J�{�qI�Z�8�+�m鎏� ���Q��LsU�Zac�\&vfiv��]�^CѼ%q�?Q�yH1pWq��}sd���"��-��h���[A��-n�*�z2��9+��JF��'û#�dh����}��,���[�8��FG�Y��+��~�h'�>�}>en�yҸ���H�?IG��p��t-���^|6Hl�j��<>�;~�t�,�u�=�@i�ob�Zs6_�Zm�NKW�>�E��+��ˑx�A{����ɮ~褖�^� z3����=�QN{�FJӹ�,er���U+��zv��vZə���ׯ��j�镯����ne���5� ��M�=��1��mg�w�c*��,NĮ�7y1fn��'��0�����NK�x�����`��U�x�����0�3��k�/O���
�3*{ݞ^�{��fٮ�Un��j���9�DW��%��x.ȃ8=��v���VE�N���Ԯþ�}W5�	�O2�2wu�9��}�UA��Q��IG.'��&B���s�}���٬H�DoV�q���iL��Y~��|��x���}���n�U����_D)�Fo���v��Vu�ޣ$�x���@�7�fU���c�zw���`҅z�{�y�n��<�꾥����x\WG�0��E�t}�5�6��,�
��Zz#`���ǔfa�	y�qo��B��[�gQ�QƬQ��:$R��N7�������.ZK�:ҔW�c�&N���`�}�-)c�s�OK^���Mi���@���zP8߯�Յغ$��e��Ig�*��~���c�a��0�2��Mib�ɝ���:�{{i�B|zĶ��ꕟ�-s��&�p?�������w���zi��I�:�j�b�b�&u�'�5�s0�/my��ԝ�`��}~G�ϑ�E���{17�%�&T�DI����P����Í���ϼ=5��v�X�{���>�	��T>}���J�Ko���ļV��,�?Q�@,��G���Ҭ����vO�W�Gf�
��9�l�h�?+�/Ke{�����>�r�^V]2���/{�UC���i�4���RO�ț��<��l����<���AN���$g�Nd̔��6�ŋ���L,�m~���Ԥ�ptJ�yU e�������}<2�Uk<+ vQ;�����w�{�z}��B�F���nY�V<'�ق�ۊ�LM>�i�Z;�%�]��G�f��Mv>�^���m���c'���=;H��|����"�W��\J��� <;~�����_�����V�y��m}�U�V2xy@�����S��7�s�D��i���P���(L�t�bMw��F3wPu>Nv����ѣ�\�>;� j�b����ó�:�+�^�[5�d����I1e8GQm��;��?C�w��e���E!ݧ�F�e�.~���3�Ҩ{!�h?e�ۦ��3���c���b��7��[�*�v�#}kd֕��n8�4���q��l�9�S���gh
�����Va�Q|2�(g(;^�JY���rxm�mh댝fke�35�i~5	f\<��v}1�Q'M{�Ly���kUV��Z�g�/J>��B>Ӑ�}����u�N���������λ�t����B�e��E,�ۃ>����V*�=����n=RQۉڇ�>���+\���`R<�E�-���V�w��d|����ߩ;Ag��BFy���k��O�aՕP��emC��u���z*��ϖ{�Ҫ�:��!{��Nx�޾
�{m�4��=�g��zn(��D�TVz�ϽعEt��Da�g��t�1���NF�_����q�}/��t�+5�ٿe�/x�Ft&���v�W�X+�U�L_�øɕ�ɟ/NBN�Ws�i�^+O��>�U���Ӿ�c}���>��zl��	gҤ�U�&*ygȶTmK��z��|���
�u�_���oC��rf�X'�i���>��Ź�Y��e,l���\��Ş�U�M�pu,t-ʏ���� ��uwe7;c�C+7TLB���P�ߝ��X�vz>�f��2��J��NGk�7W��=�fu�ӎӗ�
wZ�U���z.Ӹ$kP��V>�*�dX���_��"�����<c��fʐ�T�W�-�*�yK͖}z��H�~x�
�#"�^�%y@ɛ9�=�ܯq�/���d�7��[��T�U!
��Xp���al���}�c'V�})a�FM��=/ԑ�~�@��u�£�n�~�w��>s=�FG�p�ʊ��79yo�﫺��X|Oq���Ҩ�t�zJ���� ;��̺!zO���)��5s#:K��ez�wly̒=�l�����=�5�j=~����γ�9�:�_��`o����<�V�����G�윤6��tG��ZdW��|z4����;�϶�.9��)O8c�;������w���̦�g��}�Ito�h��ʇ�[��O�I��:��J�Kz=���g�������,�#=�A�����c9r��	XO��ӳ˜��}��ޞEhW������8Y����ǌl?UO����*��ݘ,c�8*9�*x�L�;q;P��g����t���My�[��W�Y�G��q龦 ��[�/���FDw���箅����/mO>�/��C=�;~���p/՗����:��
XB>��mg'�+.'ƶ�+��r�K&;j<�k)+�?b�$�����.  ���>��샫��c�-7��0��ʼrf4���v�Z%�U�E�Wpu8goj˒1��Y>�s��#@P����]�q�R�T��J]��T��q�N�L��E֌ɰ�X3���_`2��Ek��N��Uui�q%a�xu�Ö�sFx6�S��7������@�j{i�3U鏐C�XC�q�{4�׷��PPc���D1c���UAt��i���ee`nYę�mw�C�VP��vH�v��ڀ7�/�xx�aj�Ke[�t�Uf�b�Q�L���WL�o�h������Ccu�ң�:���}W����7��B��qa�eOAKB[��d��1��I��0h���Q�f�q�����3�vI�uo0.�	x���nU�:���]�k��E�%����b�	�k;N>�*��)7~56��n���i�3qRd�W���[K0"M���L�,�8k5Ba�����WA����,��/\X����01Gv�qŃ$�X����ҏ��O2���V�Z[�:�L��.�/v���|�H�g8u>�v��"$�����)R���H������)��x��d��{H�R�8]�6���<5�������B�+�����=��E����������˒!�e�G��K�PW>x��_j����_�{��%�P_!&��ۺ�5b.��:�eXif���KEg�79������㍛Ֆ��@2����f���"��*X�~^����ڂ�CB�<E��l]�H?e�V�S�T ���Y8IK�e�#���v�j)�%���/K�:�	�q�;�N��^dH�J�΢hUͻا,��u�S*�t�̰��]�p#��GW��zK�/U6�-̵����'<l@�����㒻!�<�۰�}����e���ñ����vǧ.��д�9z���H>L'n�WAǖ{0b4����u���n�Zj��*ִ�j�rv�A�Ӳa���-fgvBZ�7��
��%��b�(���.$�R�B�A����N���\�kw���N=*�L�:>� �i䋓#�_7��rn���k.3�or��ҙ�;�O9��}�u��)�����Z������7��:�L�s/k�L��Ā�}wۚr?���!��˪�<B3��|&u�݀J�g��6���nfW ��I��Gy@��{�u�lL�.�ِ0���qoe���Tְ��u*Ʊs6	�ɦ��w[�w��b�[А�-��$ف�KP�P�ԑ�m�����]����J��)͊�#�NE*Ǘ5�֤�O�]�C����t�5��{.-�m!��[C3�;�i:FL��c�*��*��D�b1A�[+,Q���XV*"֊*0-�
����Q+*���Ԋ��&Z�4b���cR������Ȉ�F(�B���EX�YF�6���m��U��h���X�l��"��k.YX�[ ��QE��ڌQ+�[�U,�̪�F"***�lFARбb��kU�U�"�FDV�K@��E����A"�"�b������Qq�9�Q
�̲QmE����DV�(���T(�e��R�)m�����F#��*1AEX)l�b"�TFVTk(���1b6�H��TLh�,1���b5,TTVҕ*8�r�b��0U�`�e��2��X���F)���Q�(�� �T���,�Q���AmYb�Uml+`�%X���Ub�,���*0m��QkZŪ�D���TR҃j\�r�-�(���R�*��h��RZ�J,U��5B��F�K�:7�)��� ��/Y\I]��֎�]S��ݽC��Ҧd� Rٓ,���W.&n7�z�B��yp3L:�(d�7�X�v�{k�����oO�o��@������x���f�5Q��H����d���;C�{�q�<�����N�Le}5���L�/\��㌏o?_�Y�~=�b�;�}ַ�ԋ��o0��T"]e��C���>9�[*''늦��crgY���/9�|g�:%<���U��o33��[���+�}�u����HܛeM�Sjy*�)��ɘ�=ɡ	�2�oe1��N+&}8pa�X=�{��=���7�`,.�y����u�u�
���Ԫ�G�F�~�+���u4��d^|�M��p�d{���?_��
��e����% ���qjt����y��e,U��ͽ2�}��i\MĿZE��u�h8=�t�}Eػ���f����!�G�h�ӷ]T(�h�@,-9�/Ƣ-�q=-_�\A7ģo�|[T�;:0�V�S��ګ�@���!�*D�=�x�8�c+�^�=�^�s�1��涗��V�뙞�c2�{vg��:���]��J�h�G�uo+��5;Gc\�wd	c,?[��t��W^�z�i7&�M�(�X����I����{B
R�}U\��y�
�[�;�t��v�L�} �+��\a��s�����\��9`�jv�g�s�j���
c�����'my� �h0���v�6My��{�����go���_�-�.��X��`���h��iVr�T�0{d�{�\|���9ߤ����\ �~�@�Uyɺ��[��g���Y�Q3c|5Y���JufG��W�)��e��T|_���_C���8�MP�Q˟W����in�g��Z>;���[6��K����mG�i<��Ϛ������~��`��{�J7ŕ���ެ�6����2Ϣ}<2�V�a��ߴ�{�nK�7���g<@�zN��v��R3ԹU5�=������{zY���'�g0�a��L����������M>v��Qj���g���n�_�˷�ֳgO�8�'���/a����udU1��ZX�wǣ\���:�{}���ǧM��o�1@���G����{nt'���u�1x��g"$��P�j1]1dβ���Y"��{qy����w�H���޷��^g��^
�塶r=�ƺ4���c���0��^�~�ǫG,_�_��=��L��w0�K��}ޓ�=���B�R� �e��$J̑�eSr���ы������W�	����Rr��47�?+�gЏ����,��t�7>�_��^pN��M�D�?]:���#����.��SJ����
YPe�S��eC�\����k�I��Dن�U�׉��G|�㑥=�w6JV�po��$��8w�A��"^����b��O���mvo�c�Z�$�{����]U��-���E�#�yΕ}� 5 ��p]̙!+��Kgr5S���ه����J�/����I��/?|ن��:T���z�T�;Ǚ��x�l�*��	�F4.�d������������t���ʟ}�9߷2$W���(�>e|`����>�i�%�����zl�Hy����J��7��w��>urn<���o@~ʂ��P������E�Lo��kb|�9/��U����GGi��	���I���U~9�@y38 ]�`S���'>���]:������:�s�wػ<��r�=~�����}F����Fa��ײp���	F�̱�g�`5}��#�E,��^R�q��o���>���ͭþ3Ѳƙ��ǒ��|�O��E5"]�w�s=��;�U+B�KC=r���G���O����;��FN��z��3[L	�~���N�x�8�5݉��g�{�w�S��U���+���q"�Ó�+�X�٭7��/=���m���ĩ���V��m>%B� �;�hH��i��g���FYUemC�fmm{o�Ӛ)6�j����Zx �N�<�q�Xr�����@~Xq%c�^9��X��&[���þN��M�������.�o��\yοa��n��X���/s�����}AR���E���"�;j���a7��T<79��x�w�|�e���Ҷ27D����>��!ӗ~�xM�6c�h�}�wy3�p8	�2���{
�������z�G{�QT���j��wz�S��������	��q댙Nb������9���������Ɨd��\OB� �HZ���^�~�+>*��L� ,ت`MO"+�"�ȍ�c��{և��3�y��ct{��������q�����z��Գ��S� -���z�[ TY��i�F��<2nҟU嬼Hz�+�=�޶=�e��>��/��+}7 l���P�T�*W�a�28�<�eZ:�E�5�0���Hȹ~��C������T5��7"�� O'$g�YU�D���^/c��7���<��	��U���>9<
P߱ =����U:"-vV>[���F.��]�G���`1��DS=� {�0�/�]�Q���U�q�����[@,�i�����xL�o�K6h�o�d�|�#�9^g��U��#Y����J��n|Z��kpje׏�D߂��4�Jv��$��xS��4�&I�G1ٸT,��t�Z2�}[F�#�� ٽ��c¼0"fxnxׇ̋}-�xa1��sdģ=[�\>9�\�(�7����잫\�/t������^�V^�3�v+D�p�@���B`/:,��1o
��ӍU�Y݄��9_5�Z�T���r�^��G���#��n2�K��\�����k�_�2��"��y���~wfm�U�]G�Dc����g*Aށ+�>�#�����0�3k�GB�������>����ō���>�@	��w�s�>"�}H��{n���5���PGnv��د�A����5w�w�J&�f��~�ڭ7|�M����݁��վ#>��Ƴ�h���օ��=U\�V�KJ�����x�Y�~��ۇq����`o�㏠m}����N�ǫ_�9�U��?�?J]͚9[���[P�%�!�ȕ����/c&���&w��Bs��f��x�+~)ʳn���F�5�n��Q��>׽p�IED[�%������0&�X�ɝf�ɟ"�Pw�~��'U��㓆w��z�X��Ӄu�㾋�y���r���G�*����*n*�<�~�ˑ^�wJ�f[ٯb�����p���BGO�X��v�{��Y��m��qw�x�L��%sP��3���'g]�{�y�岸�ُ#O�P�����������^VԲ� l���E��w��=}"��Ƴ����aJ�Z�M=ne_ݔ��5�ҵ�V��+��T�(�%+w��/+C��\V��T�[GkbҜ�;rwmf*�ŏ����?^b�Ž�Z6��Xb�	#K��6��{�x�8��ċ&-�����P��#*%�`��>Gۑ�iTN���\O#������=�:��|����Y�}5+yId'ro�:H�D�m*�_>G2ai��~5m+��}~����q(������{a��&�ׄߢTg1w^(��Ȩ�U* /�T0�"f)�x�+t@,eDr��������=9��Kk�S���|�u��;����pe�*���z�n�����bi��7�úk�.+���[�}���urt\y���#��yNC��=~9p$�/x�⪼��M�=��0�znw�U�3X��%K��N�չ\4t�ǣ�Q��PX�]���>�����B�=����N�nG{K�U�3�^��^ͯq��&ra��5U>#}(=�Q���r��P}/&ә�R�9w��H�/�TB�s�����v�t1������g�@��ʋ=�D*x��U{7y����W�7nt߼�#�n��*�?�i��k�xfy����w
��l��NϺo��;J
�w��:Ę��U?>5��g ���F%g�(�c+&��y3�7�@קQ�����p�y�,��B8Fn�]��[SNQZe'��,�To!�{�&��9�=�㛧$�|�8�Z�1���g^�s��b���HSj�l� I`���;vf>��x2�Ŵ����s��:���1���YӖ�c��ԫ�����6H��^��ztuC�;#��(���M��9���C��R������4�#0�/�*��y�1߼�����o�#|����~�r��џ{�)��S7��	O����B��-˼Hy/A�w��Z=2���yPi�t�����x��+�Y�y�я{���̷���W�.�g@[7P�p*����]V9K������m��>�q�D�Bd
���;��O�����=G���Cf���G�]4N<�(�a[U�{��m���ݥ���z=����(�U�#<��.�����mz�Al�0P{uR&	�g���ς�ȏBj�^Wd���f~έ}��;KŌ�\߶N�q�ˉ�7>�l�A��T��}>� ��Q���x\�n�	in�_����H�dz�_�zv�+��w�܉�7����@xW�=�$����t烻�����(z=�����{��0��%ޛ���W㞟P�� ~���ג�w��p7�L�OIR=Y=o#�3=�m�m�j�Mi��Q����%f��s��6��#��G�a����&<9�,��%ծ*�;�L���ja��yH��c#s��x��r�lu�AR�o/fܬٛL���Z]w���E�_N�r^�����y�V�U�]�ޝ�#�S�M�b����K�63���*��o �l�=jvK���0��,f�mhw��3Q�ƙ��Ǫ!,̇���Ϧ*�<��$ b�ٸ��g�$�<g��M�Q�_�He�ȏ�?�{'���;���Vv���<~�_=r`���U�#j��Ǝ�FS��z#�L��dЭ��nt����#�	���+A�4�kT�G�*;������ ��4���������NC^��������Ǣ{M��F����Ve_j�:�_��2�G�OB$�?Q�nҳ����q��F���z�%�4w{�!F=�g�:T%2��fg��ƪjy�~��O������w�;�>���X��s��N�K�]�Q�5~מ�z^I`1�ο_�wB����^�6=}U�/�P��Nb�g����k��i����<�O��B��Y�~�ӄ�_r��؏��n7>���%�*@[U0&���ϑl�Ա���z%[� CU�����2�D{�;h�w��n"_�=bV]3aĺ5�WR=Q-�,w�p/��C\�;�V�*��]Z$z�3�JG�=�F����Yȕ�P��no�'�=UA�����Q��ۣ�f$��b�&�w��w)�D��g(+u���9���'���y�o��[�܊ݚ�g��B�nD��+��:x��+q^	���<�ù�2�+���}�kްا����Q:{S��
�5����X1�C���w�r������_����%#����9�H�+��G��|<|fY>�q�1���c{�ս��'�<�_�M�]�<.����޸�u����p+����rǨq�8;��掕���F ��G�h��L3mQ���wN��/MG��W���}&_�ؤg��g�_r�X�ݰ*=�۪"��G�n���Q���ߵ����RVn��%��[��ٓU����q��yNz�`zᜠ)z��y�Q~㶭ײ}o0�}k��]g���dd�o��u���w���}�W'��A�/��Aٯ���|�\�;�
��O��nT{rw<�����]����g(p��}(�#T�ge�29[�s'�(�R'����@�����}��7)~c�e���X�ڗ���ʇ�(��J�^mV��g���'��^��
:�p4�G��"�����sf�8k�p|W��m�r]�؂�fQC~�YE�Tp]3�a@3_ip3T��\����7�lz�j�tS��d{Λ�Rz}�ݵ�W�cCt����&U��ҭ,��Vy�����?g���g�G�
����j^��+��V�P��U�4���ݓ��L�Oh��t�+Y�I�"�c�)i�ќf:kZS�Ә���p�30��}�aZd��F+ԧ�>�u��^��؛�6^�+���ݣl�57�uӋ!6��$��Wp�Q�ݡr�+1��wC�X������:��p4���+Vʦ���	�ZY�-/�|�<ɕ��7԰"���/D�3���"<���_��n%b��{j|c��em7T���D�n�1�Y&��+]�/wN{,��6i��}��z3�%q����8���+K���>��% �����D�{��ù|��P=�@^�x���4j/_�G�����wi���~����|{jQ��g�׭���Qۏ_p���G���<��
��;@��-n�4i�TK�~��?IG��p��|TM3�t��g}G'��u9>�$y����vT��.|�d�Ӛ_��i\M�k='y�F��_�E�����μ3�ģ�=;��~�#�2聘#�+�"e�Α3�t�82�k�Q>���_H�k�����WL{Ӵ�3�9s��M<��.TKG�n���x���h��n�j��d���VSGR�k�*��xm���?Mx�u���t(��)�0fgȮ���?� ���5�L��s�my�O�tق�Ҵ���	Q�69���9ə��+�:h�^�(����(	E�U�d�w��x{�rN�qG'I����u�:m�4�
�%�N�L�ۚ�[iA����w����tv
�=ܴ/PG���tq	ͮ�5lr�
;��m���?2S���sI�ً�r�����<��>GԵ_J��z{�Tf�����̰�2��+��^�9i���<~B�e�Z��Ԋ�w��s��a�峧uj��Y�ʺ�m�Q��@����jnj��Et V�F���ۤf�:4d%�.�uD�A�e;����D9�=�!]ea��.]�C��H�Kg�,i�52���՝�n��-�[�(U�W ʼ��oD��p�oFo��	a�?mS.�p�������VV0yL&�1���6������J�\_b�u㎮fv�����,ݓ���]��=2
:4�q�)@l��tS�;8�#iѧv-*,��x�\���ܻ�2��hȯ>�A��%ڽ�{��}Vi��6Owc�.�*���α�v 1�iGjˊ����y矹y��E#z0��[N9���hE2���i�'LEX���������+�@�ה��fnЉ\^P�j=Y6�w2DHMͮ�,�E}� �"���'j���)��X�yv��'c�hP���Q��b%�u������-�O��O]��!~m7S׬�5=:���؂�hy<o-��kj�q,����g�,O·U�ꂜȱ� ބ�L�<���'��m�����2�r!����6�@E!�AHw�C&����ҸU�sB���Dn�B�`ܫ=�/���r�x9����mpӗ,l���_A6�aE��#=$8W�c�&�n��X���3�ړIk��-������c���25�M�È��^A�F�����!9�us��'^��������b��*���e#���1yM"�WZB�ܶ��h�CE�T8��=q}|�\t���5�Ux��lq��ը��q��ODtfu5)9��Ͷ�Z2�v�0�-6����bVFiκ�$���P�^r만6Qm@�2!ʛ��g�������������!f�5USzR�ڸC���^{���{u�2t����*��I��P�t�h֛�s��z/wD86K�;
�NU��͵�>�B麉��Sr₆��v�֮<���x;�Q�&���ngSZ�@%��D;�5���5������,��<v���v��CN]�9�Ԓg]�[�RwPk���PN��ڽ�`��]�Ĩ�@�4����oɅ^u���5����g]z9)�v�G��6+y��h'�ۂ*!��3��,�1�c'�H����.ƹ�]��d��NVD��^<z&6�L[P�z'��E2P�Yz��٨7��Ħd��-rf*÷�����K�{ؼ�5���^[5ɛ&��r�|=u��[Z#+xd3ƏnZ�kzA�N��;�R%�b��Q�S�ᰵ]�c ��p�/cc��IZ�5�,u�P��B�K��x���5|��f
�
��)��C��ݰl��Tk.nL�����|���w��|��ߟ{߂��X��#=h ��Ee�H�2"+��c\Kp0PUE�aE(���r�b&$��W�*9DJ�1TQk?�*
(�G���P��"�i���2,ň�*+q
��`�EX��ڬ*UVJ�.�DG-V(���1bŊ"�*���iKhiTm���U�"���\��(���t�(�b�Y-J)mKj"����5qh��`��1bV���)�[m�cUR�[�P���X�[k*"��QjJ�)mT��0�J،bZ����+1�۬�ƶ�J�V1����U�*"�5�j
�T���%E�I��m�.amJ�
��(�,QKu�[lEPJVЭ�U���̬Q��q�U�1�l�U��KB��,Z�PE[JVT��%J�+2�l(�Ҷ�RڍB�L�cV��E+UmYU+%�
��-,-S�U"�k
1VZfQ[KiH��Vэ��T�U[h,�b ��YX9V�TA�t��1�����W=&݂7���_
oN������G�_d�w;Z~���"�z `;۶Sc��a��|�^sq��}p�/�v��T1\`����ͧǃ�g�j�{�~�ψ���~�����G��Va��t�3�C�z3�Q��J�a�R��r�+q[Ճ��%�|[�ǵ9���d���oĪ�()۹�y�kşGv��_���^ ���P�6�i���Ұ�N�r7�|X�ƻ���r��<���J�u]1�#}��F1��s�R�b�2kK�L�7�24�F��i�K�7u+K�ѵ!m�����{�o��s���ڞ0���d��T?�I���8&�����|s�����6eq��a{��͍^��s�:�߬�~��2<�:��{F�o�D���H��΢��aD������`�p��%�⣞T;���i��J�Ko�����le͑����o���^�wAG��u^�(�t|�Sw�|��2+��Ȭ^�ϸ�V����|�\uA�}�}��_;��z^�����G�S$x�h��Kgt����Ћ#�Y�V�㗅d���&�@]2����\=\�G�N��=��|=��,dٳ�U ��w�.W�w)t�������|e�?���Ǐn;[9��b��^H,f����H��דT�KA�[)�h�z1K\{��vzG����ȥ������9�Z���R�~9��s��U&��	]B�km9le-ɺ��y@�VK�l/{/��n.s���e�tT�iL�1��?�{��3/u;L���E��d�?m�Ll�r��>f�n*�1u=~٨أ���{�,��y���{��}	�G�=J��=;H���;��D���znʠ������������W��H���89�0��/���׊�u;� .��`�Y��N�-/k/5"��g�	��p]�gy�C��Vɨ�����^��J�C�~�e���Np�^y��y^p�]���Ae����yϤ�ȃuป>����ћ^_l��f��ꄳ2g^�R���k�oVU�N�{w�G����|=r����?��gD�~y;��:+M���n��*�z'�����H�Ő��:�Ѿ���;V*�����n'�ӳ�2�ŉy���~�G�����Y��{���}� j��ɦ@�^��'az�W�{m	��Z.!{Mw�Hê��-�V=�s*���ː�nGW��uu����#�4v�q������w��1���H(���H��G6Wr�7�g���>��(<UQ팙�M����ls��NDo���ؿ\l�G���$ �VH�e�Q��
��x�;�UQu"^M`�/�e���ү��U�>wb��em��O=�W�ӵ�*�֮p�{j�Ub�!<ŔbS(^�I�;4����W3b���TsJ��ќ+�l�Ko�� ��75ᗨn쳇o�l�YE��Ʌ�hՔ;�Ǽ���f�"�4=�T���CܙNb�ɟ/O3!�<��^z�k�.i�^ֱ^Z3᧸�����2��嗞����Hn*�<����-��jX���}���Wn��J|��}�=6W���K�?O��~���,�gυ;6T���z�[ y�0�!�`�~������Gݸ}�k}��w޴8g�鋏O�=��������A�j=D罕��O�t:�>*U���X�*����� s.��PպH��~���J��Y+�e��p�^������O�a����N��#�6}� n��t�ʂZ;�&�$�Ȝ�Z�I�)�U�M��ٷ9o*-��N�����s�5� z;z�q��7�W�j��s�w~;�	xj9x�z��w�я}��\H�ږ�9�;����Ȭ�Ӳ}[@+����y��!L�Gz')����G�"�i�_k���XΪkj��k+#o�;՛�O�����Lg���l��g�`[���F��Ȭ�ʇ��z��t�XQ �M�F{_�>iGo4�gg�y��K�z����=7�47�]H#{�%a��O��u�=�A��<辵�}0�պ!Ww��B�uq����L�\E��6�
�r���Y�� ;T�'Y�Nmuh�m��3�P�M]��h�7e�|���L_,�H.�q�rjva�6��&n�&_A�{�\���3�B�Z[�+3J��kVPg���k���u��X��t��L1����T���'���]�cy�*x�P�]&���n�>{ds�~8s���x��כU���Ǧ㩀&[�9zw�/��M{s�A�]fȩ�=n�_i��q�����S����t�^���
��򹸍,��uO�m�΀��:�S�T�{&��z_gO+�Ϻ���ϟ����x迧ʴ�Led֗d��b��No��oP9QF�~�Y���}ϱlldQ3���^��;~��o��;;�r�3�[*rp����7=����:��ȟ�{��Oo��^�6�dw�)�x���q���OĻUz�g��L��o�����}~���6���]`E'cׄvOq�ɘ�^�&X��X�J���^K�A������~���Z�WVâ\f�yk��j�z@���8M��e��j5o�q��M��x׃[Z4?W��a�3��w����t��~
Ozl��n��T�h-bچ�[J�K�$S��y��Hvk�GB�����j�xy=�t.<��@�!�)���T+�����ә��񨶕Ĵ�G�D�b*�tUwJ�D��F�"�ݑt��$Fm�P�L��j+���fP��WEs��� �A��9Óa���d]*uo�nz�H�	@_YsFX�"Moi�������n��^�;�组�lao7���ٕ��+��#T]��^���8�:l��iy?AIPܟm�l�x�r�J>ڜ�]�3p`�ʇH��=�x�9�/�C�]O�_m{�B��*>����z�1q����s�:~ˉ���� TJ�h�D�Cܟ�ǳ�G؄ǽC���%�ʯ=T}�)���J�K���>��R����z�4�誯#уz�G���Ӿ���wb�^����i�\g�����W}�ᢡ-ɶ1����z�sT3�2@�梠3q���N���S�Q�E�v�}�g��n�z�6�ǃ�g&���/�!�����=�RF�2��͝���>\;,���*Y�Q��QI���zp:���zX�L�`j��l{۩i�U2�L��;s��L�����z�7���ۏ{nt�Oa�BP��v��ɭ*�|+N�3��W��LXƖ:�絊B���=�W��s��C�r7�W{�9�� ���}��[K5�[(ݨ=��/�Ovj_�g�j��?Us˷ܿ��[$\cN��w:9C�Z��E�̶W�EDh�)~*�G�_���I������q�L�7�L��}�"6�W���o�y߯��%塣#��H)jE�m4�z�ˡ영%�=2���Qs���h��~M���-��a�� ^e���L��w0���,�}!Bv0�fg�@�C�{|9Ia��=�k!�M���UУ@QU�3��bJp����W�"�l�����z�+�+���mU�v�w�PK�q5S�65I�@er�x
f�c�\G'�}N��#�x���g��^��j�nFz{�&R����Uh��.��	M��Sw��Re�}�A�|��<�����߮B�	O!Mf^t)�Q=�Eύ���O��O���mK.4��@�_UH�}.�&��c������%K���m�S�=��>�>i���i\��؏����������n�D�Ox�:e�~1"��st(|�s�=��{��&�]w��(�q�9�{s"E|��,��n��O�G��'�s˳R�^�c�omn�%�gr��'I�*����`�	��A��7��=�&0�'� ���&B�Gús�2�ա1O�h�x�d@�xj��yU���ܜր���/X5��9��+��7����}��x����*�ᒯs��_�}��3r_T&s��&��������/���jif��gUh~��)�.���������d��l�&MF�=���y���/P`��}��˛���7G��uh���Z=��M���C/N~����=_�\f֏a�8y���ض�p����ӢЕ�J�m�*��%��G+��p ��2��T��b�U�ΐ*�_�3or̈́ay�]Y3I��'c�ΐI��=�6���nz��kj����'{2��q�o8�ۃ;3��Ɠ[4��������p�A�`�J]3��<��Nߨ��=^�=�s����\��hV�mΘ���4���q;0�/��^��ӷHc�z^L{��٭7��}��ߖU����~D�� �;�hH�����q�k��,{&����9�T2s7���7����'f⮳o�wR<7���b���w�GWy��n������Z����t=	mK=�80��Qa�خ��d��pze}�,m���No����PI�۹�{�Ve����Qt�3�v���}R���F������ި{�L�1y>��s�*t��}B�m��u�$�pq���E���m�r��uL�@Y�L	���>E����kW��V%ރ%W�_�v�� ����8�>�K�\z�,�>����UH�*����}���"���n9=\|���W�|�~�/����q��5��q��o����d�2�����f�{Ӕ�u��fz�F
����|��>چ��l�_K�6|���m����j�/X7���.�@U>���:O��Ā��qJhQ}^ÐKGw>�4�'��_�|rx�1�#mGUP�f&�c�&�~�|��7<:�s[/)�L�r��^�@՚����&w5/��H ��lB�Ҧ���Ai����i�.���N���R��0\�%�wj�B�e��Rz�2�]-�����qP��=z���f��4-�e入b������7[��- /зnEG��Q�GŢ`xfڢ&)�i��������zn=qT�uY������y�r^���g|jMǔ����ws�!���')��I�V����rTg�U�v%��p���'�k�Q��^71p��yN|�v��k�����>��#���C���.Us�[J������>�2}�:��_BUr|/�nϲ3��r��zht�5d=���O���A)��r�۸�=9�Ǣ�ѵ�af���灚�� ��_��>j�|F�Q;��mؠ��pu]Lt�E٩�[��,V�8_�'h#���y�w�U�C���i�*1c�.!zs�_˽p8�7˽�~�փJ����O�{c�Z��<3Y�n�X�֖=���o큞���Q�k���7�^�_��׿7��R�?�_�+�F�~�q7�۞6�Ԏ�O���U1��Z]���b��!9�<w*n�H�9a�S�/t��)���8�?{^G�um�%�l�:�*�=�����4�=��ś8ݟD)�edw���3��:�=^�q_K�q��s�7©��6��C'���~�>�,p����l�v�>����~7��lg[�w*׽'%�M�R<�L��*&cR���S^�jP=~��/ʴA���i���M�+yi6ţ:�5I�]��:��R��[-w�����;�޴�K��TS���}�-��@O~䋌Qjn�л�[K#;�<�O�}=�
��3q�1��f���t�^�^B�+�>��Y���G�����y��{��ݩr�8�,�A<ۉ�p&���ԯY�~�/��6}��ڷ���Z�K��z噥�\*�v���Iҽd�7�fA�n�8Z>��7�Tm���{g!+n1�O�Լ��K��^6Z8ٝ�~�'�Z$6n��*�Eϑ���26_��X���GSr��w-��rj}���9��Q���Oqܹ*�/��>f�yPՑL��s�2������N#����O�ǶeW�/�K��I��\K�� _�G�n��h���:!��s����ur�_��b����"���[]�d�m���"=.���ptx����zmS�}�LyĚ�RX���&���[�=b��_i��U�W��J�1o;��� {��P~"��l\�z=�<]�Q%�=,-��y���^�q��3_mC�̿j�|F�y7ޚF�g;r��m�z�g��P�.e���G��ZN�/��Q9]7���������&1}�z扭�:o���C�u=�q�қx�����kL�:��ܶ�S��g|-Q������}�ٸ洹[��M���ZD\�N�Ώ3�e��Yr5s-�:�T��d�	��'���E�C���L��+�#Df�PX�6�n�u����
���u��p����:}榸xdw����\��~�����g����\�oK_���,�BJc&�r}�ۯ�q>
����֫���w���o���o}�<b״�q��:�X�o^c�� �ɞ����>�h{fW�r���{o��l��ϴ�eh�~�C��\�_яM6x�{���}��MKI_�	^��Zk=t���;�q�>	�+�q޷㑮}�~�8��0>�Ϗ��Vcz��ez�qz��'F�7&�Rf<����[��G����]{N}�┲sJD���0z���os%Ҏqy�z{6�2 ����~�)�Pf�'�n�Y�r�l�h�W?,�C�w�6�e�J�#'$�G��;�<^�������R���Cd"͈���Mq,y�����*h�=[O�`>�>�Ư�����1�AW3��:j#�n��W��gD�o��۪��z��a�7U�՞���>XkO��G3e�QmZrݯ=�}>����=wLz�����>��ގ�{��ʯfi���"��XLVl�:KGw>c�w3���Sy޽o����]�֌!	'�	�`$BI��!	%	�~� BO�$BI��@�$��H����I?�H�����I?i��a BJ!$�	�~�$ $��	 ~�!	'�!�~� BO�$BI��I=	���e5��F�ee� ?�s2}p$�=��U��J�I	QD��T:h5�`�IAkUR�6ɠim��H�%T��[4$ چD��f��U$�������JSCl���զm[c}���λM�l�ov�5��m��ꭴ�kU3eM��Z�bkm�Il�lж!;�E�m[ݢ�V7��f�ضd�hi����b�cl�j��h-�-5�Q���[5��,��mj�V�f�jRZ[[`Ve�ڭYL�Zm4�M�E��̶­��j�5��Z�v� �m���[(l������  �y1�wwGw��.��l=���{��j�j�'����9���쮽�#[�;@v�7���#֪i�m�ײ�ZUY�*lK4l��B��� �u�G��n�=h��)�&��u���(������QE(����(�F�Q3޻�$
(��(��Wx��(��(��{���E
�}��yEQD�(��{kJ+-,�Xml�m*�x  �xV�_F[5TJ�wox� �t��֎��s{��������Az��@��[����	�s�T׽���=�ᥫ&[V�V�6�V�m�� �p7�v�u�O�uZ�^�8���k�y�v�{�w��s��H⪝�Z�h�����^��P�m�ݛz�65F�� �{.�۹�6k5Jeu���
�`լF�6J�kf�V� ���>�TӮe�k����ݪ���w�B�{i1�zU=tuǦꔚ���Stt�zK]k�w��q�4�%�z{�ru[��n
]�3��-]�n����s�5��ƩMY��Z�dM�mE|  ���֩���/#�z�݇E�{�5����wu����Z�V�]�=k�Hu[m+���x�����p�r�ۃ��������m�Y�jm�=w�w����]%��Z��d�j�&�5��{��|  <;�}gV�m�-�Y����^��U:�u�y��Ud�l����Ҏ�֥w���Ű��껊-ooN�6\�;�tu�[��޽�w[��ܣ���=h�[]-���kc�5����Skm�  ,���>ڨ�޴���� ӻ��k�Kk,�#���u���j�=�w��^��{ٛ\��z���)o]��u�m޲��4�[{���3�:��J�S������c"Ԓ�VZ�>  �>���͍�yw��֝ivwAJ����u]�ړ{�x��׭��n�kz]{������{W��z�7z�^�ukP��M׷�sT��Wt�� .헬�,�ښa�[TDK-=�  {ٯ|�v��V����Ы�U�wb��=h=�w�����N˪�<wWV�ݵ�A�y{���;�&�[�-�m{7��k����7Y�kM�zz�������eIJ� )�4Ĕ�!� �F��R��?R=@Ѡ���T�   j�Ę�UM d��
H&ʪ��f��T�����ҿ~g���������ݐ�j��S��ey.gup�g�^���^��~k��z�WB��aW���
�+�TAYD@QO�}�l�������λ�y���֊{�P�XZՊհ�-i�U�Dr�i�,i�ܔ�u�,F廂����%�ʼ�8���l��ĝL4��f���Gk*�4QIAR�WI� ���uxm4�B�{y��v����S%
����aP�edR���5�o.fû���Re�4���V������ևo(��۽Y/w2�٩e���J��Y��R[�DU�����W9/Uƌ�ރj�t�]�+蠚V1r7 �ɛ+��xDV]��k��9#ӷ�^�@�Y�j����	P��&*��A�����GwVP�S��*h�����U��bE:��R"T;xS]F ����2|�r�̶)e��m 4f����tfEb��f�۰8Y�vm�V�����X�%�ӏ O  7ki7blX�V(<�W��%*f(�D����`�Clhn�����R��qި�*V�Č*�suf�w���8�1nAmT%9�� ��i*%R�` ����L�n�݊f�+��a�[�V��6Ycc�u*!c,e�(i")Y[�k �p	��6�[��˱�/�:�w���-P/l�[�3���e���d����f�(Am:���Y��G��tp�R���vBb��Ո�W]1X�)���6��f��L��Y���
r�m�W`h �e)0PT�bz�VXU�-���ڙ
F��6��׆ZLwpC���.����q��v%
�D��t��S�5��V�6��:��YA�E:tJ��:s�u"�6�$��������(V�;#.�q@��7X�4�c�Q�BAN�elf�@l�Р��7G;,�hnj�[4���q
�.Qʰ%ԢU-�Bm3�p����X6��gu�3���Cn�hj��%;T�Ӽb[[��r��I�x���j9H���D+��.�]�� �4f�\2 7Z(���v�]�]#D䔭d!2�c�vv��ݒ���;N�5s*e%��OR?n�n���MJ*�/	K.Q3�����J2j�X�n[SUm���i.�4,�ce�%�u���^Y˺��0�)X�7���+Vm�F��Gjei�:���W�cd��$ۭT�݋x�Z4V�ʱ+U/s5�Ɓ�3rZB��Xj}w�m�$��K�R!Q�f�TslQ�\7DG�7@��m�h�&��R('n�v�26�)�/.�e9����76�����61�*QZ�yuj�=�n9���!� �p�V�]Ff$��Uڼ���lQvIuy+zE6��^��Ij;���9�Tu-�@P���ɮ-�lli	���&B��0ڻ�&�.mK��&��.",h�D��6ӣd\׵ �ӺY�*!W�\�\�^m�7���м�ݴӐb��%�5b��jS��Κ5���%I�,�V\���ꥨ:�M h���I����� �NJX�^���m��hB����t
�ޭ��t��$�Ϙ9�1��J�"��Jiݍl��1�mM V�V��mTr�-5�rZ��쫪�(;2�y�
e�ti�;��W����ЭdQ!J7���)ɸPĔ͠i�X7���U��p[F��U<��S�[D�{!���m��^Tu����<B�U�BQ�[9)mHe+���
ݠ��1����N��t����[3l�I	��v�bӧ+M酫$R����X����W�dH[��ы'�Ć�xa�\�;���(⫥@)��a;f���҅Ē�����d�%�me��=��]∷��Z���3FZ��J�on�5V4Vc`�׌��Nue^��lhʓ�9)1��J`8T	Հ泡���s�l�wB�� �VB�
�1�	Sǆ���4��lB�����IiĨe�WR��[���@�3aX�9������pX���*4wE2@DC�.�v"Y*�$�mF�I�a�a,�E��aвܫ#�ԃ+r\ձXf4vѻ��*��曖,�՗�m�V,�7#�P<�U�e���:�.��)�^a	��XP��A��wW�@�Z��\i�7%Ll�Z�@�YO4ٛFV<UGn2�p�*P!6��t��� #�w��3��X�*��jF����5&%z��S����)9f;�e=K�B�7JV�	]�8�l�Z�\����R�Z@�0Ņb�Ɋ�f,��u%�nh��ЭJ�O
�*��6Ցێ�clT6��!L�Y���D	W�Z[w��
t�k�z[N��Ӳj��+q� �]Ök��˰�����9zI��N�2�+3S	S~v]憵��LÎ�,�թ[g-5)Tqe��şi��J���e��\�b����&�bL)��5���q������ʴ��R�c����U���dڗE�T�:���8�I̹.��SYҩnL�j�S��Xr�SN"���.�+p�K�q��� (���V�wU�C,��H�lD-صV�����R��^��csQD��X,,��f�݈q(���˨�i��Lm��]%��c��kO��yM��ך^\���%={���tN�U�Fn+�X�f*�qQ�FZ3(=VnF���ܫ��l�w%�D;�2�ƪ�{�+��	 �y��i5Y��k^�Cr�R�R�V��#�W�r#xѡ�VPZ-��X�H��+[K!�Uw���pP�)�
��A�'��B�L�A���(##��Ju�	.�'��i����(�+F<ǹ/7v��n�%��������!1�g��l�V5ˣ�����K;�F����L��od 7 �����w3E�Z��F���E�/r��1MJnktr&lH�'�ofZ�ǒ�l���vZ��6G�kIb+s0�i,�afI+n!aDФ�٤j�%��x�S/� m̱O�K�@��x�j7�t��D�(@R�oŌ�JҬ��Kf�j2UQ�M�
�م�L�)�[im�<�Hګ����hc��,Zk(�v͝X�ХY/�R��2�ݑi�2��A�ֶQ� �)Y�vEFS�5 jõ���%r��¤X�Mz��y�S�2���#�J@�-�<������#�e����**�jAeO~.�
���U�%�K]�l%.���4L��,��-K(������^�O&(�$ 3Rݥ���Q.��#=�N���z�(P�1��F�V�k`{F��K��l�T����E�S
�9	7F/�������v�Q��\R�1@���+l8����j�fS����n���cO]��T(,Ra+*�m�[����r5&w2P��Ă'+fem��u�����h�IR�����a�@�̂*�QJ/f�UԞH�1���[��,�4B���fA4맢��TC���+wb�(J��
V[7Z�I�r武��u���%�;1b�-�#�4�:�Ղb���]������)^+��F��1�D+��8,�N�㣑��:�jr�g���MYaYѬ̓vmS����* � *��4,X�k �Ķ�ԫ_S��Q�4��/$�pj_2�J՚n��V���1B��&C�R��)�Zv�(��CT�h��n7�f��k���j솈N��*�X�8n���x��v ��Z��$��Ѐ@��D;śPH��[u�n&e2/�u�PWXN�,����ۙ�/@t�,�5�pۧY�
Fj'Z�@�w�zd�f�͹�Ӹ4�
��n�T�N�^n�o>:U2��*�X��㲄�nK��2�1�	ˬ��c
&9%4�Rմ�ҵxv�mA��6�bYWA���)�)`̣)���! L���ĢՐ�Nṁ3*��ncU!��-QvB�<�r�z@�Zq��m���)���4�����h	��
,	E��	�y@��:*�]E������ml���I������J�,1���GBR���-O]O�F��Y��V�DEY�ЕTE�f��U۬!J��ʉ+yy���j4�}Xس�]'��f���.��dÔ��-Q�)�mZ��XZ�G\_#@}:	�+^Ϝ�ub�tΊ4�3�7n�+k%�5�.I����Q�����VIb���si��jV)�X�6еl�0F鱉�#@{A��+V ��ѳwN�i[�tۆ�%�Ƹ�P6vn��X>J��`M�/F]	���]��P�k@���A٣���}i���n�򅒂b��c)mK*��@�&�0*�pc��e�nb��)]8hԣ�\�a�̏�R���Cmͩ�5���s��r�ݒ��3�I9e� �w��d
�	lST��n����iKa�[&��˻Ա
͛�n�%Z��,��VV���8B��B7H<�U�Ua�^Qا�cv�U��͏X7��\�28���f�1й�JY[���5��E�]Eެ"����Ұ��dQ�]ʼ[p��&��MF��әv��r�b��TPK�C�K�y@Jo+u(n��YX�����D֊���ZGe)�D�-��t��巅˛��=�7@�� nζ�����
�B�^Tx*kg61����G�Ybc�m�n���H�WN��h1�% �A���RU�.��ڷMꆡڭ�qӢ(�z�LP� �e��&e����T�o,X-���.�
���E[K!X�;��虲�����E��^*��}P��}%*��<�^!y��3R�cXW�aT�b鿱�R�.Q�ol��P���&��`Æ�6�aQĦ,αt�5�ҽ��]Y���C3
u�JP��˘���Sd�[�(c��V��%Ȱ��n$"i����̲��@*Vޜ����+�H���JVv�
�N��f���+�j�	m���w`��E�U,��Jh6�ء(I"!�E�u��{����f��<�.�t&`��d�Z)�b^��$�
�PV�X�b6%��:an���4��9L��n���-Z����к2\�7@��D&
c�(%�����Cr�Z[y��U,��Ć�h����1�V�]�d5�Ih¬���.�Ⱒ�&�R��v�8&Ʊi�v�hȚL�T�"AQ᷆�䧶��=�Ol[Q%�-C(�p?��$�6	�F]��*���H����ZiiYP�2rP�j�z�۴��V��܆�#�s5�@Ռ�\� yz�`��q
Y��	����&�(�9m�e(ة���&n��kh1 ��m�1L;�j���%,�ɪ$�m{��VKcR�ék��%
�v)hl�u�u����
n35[;3�6��)"c��m�U��[B�wi�+��雑k��mk��w7A9�WM�Jd�s��u����Ͷ��iE�2b�`�I�wB���u�шܰ(����8N��y����U�ˠ*L/��z�JM�m*�Wx��B&MһY��v�Ey5ar�0�B���CJ���ͫ���z��8�1�	�`�ͩ/k.��s�u�DT�QTi�3/�*�&;���#�Ӻu�����)^a�{�jEd��m��Wx���B�$��U�e��{0զ�l,�����:u`���E��f�+���e�$t@�0�q�Lնv����(`.X0RyB�e���1�
��*d�$߮&�C��5�oQ�y!R�ހ�k�0L�CR�چ�����d��y�9֨d���Y�ƪ�r�O��������XE�At���M�M�h�V�B�u��X!-�ɽb�
E&7���pD�$z�j��ۧ�*�� �����v`c�����:Y��6���.�^��L�j @Z��p�bn��m�
�J���2���n�h�7�2 �8��,hE��Zקk+5T���C�i����20D#w��ѣ7Rt)`�6�V�ed�5�����Q�����)1sM6K����9;�(	{�a@*�w��U��)Q��Ŵ쪶�F�h8෺�۳b��j�h���/���Ըi�Jūo[��^�q�w�л�7u[VK��#y!L��� �%��r�ͨ(���&��X��b���R��3���iG.�]���O#�ʳX�Bgא�4��	��&�ݑpG��f�=x��3�cS6���
�'�N��S�!t� �)�PL��ڈ�`[2�4�c���j��i��Xi�j���yfef�F�;�_��f�x�ө��;xo�1�`jC�%$n����e(�;�P@5�86�!�Z��el�n�a	P)�U�8YCF$.&(r�M�m�:�n%�!�;�|�C�lR�.�S�;([&5��8",�"��T��`m�`���j�ht���o-t�^����P6���cř�Ʀ����e�)�5e�U��M�&Gt�{b��ڧt�.��z�!e2A�C�{R������-e��!0U��Imjm-O&h�[�.�oe�I�c3.]CF��Mȅ�4H�wC���5�t�:�pF�	Y�hl��l���+q@c����$ܢL�-�7fPM���fi:5�Ol�y'=��k
�b�&�bWQ�G��MX����B��)P[��M83/~rP�a�)ȑT�����Z��]ˍ
: ���tl.bA�����n���5jn1*�KTu�:*$��,*9��J���i �"WfdK��V���ʧzfG����K�7X�7Nd��\�V�Z7i���C5[�wZT*�2���J{7S{���Ǵ�*htL��Uo9�j�+sY��*v�<�ȅ6�{�n����R�l<�uP#������H���nLQ�u�K�vb���5 Χ]��K�d�P��q�HB�hRa�6M%��i�������J�=�S+o,E �z�^����<����x��G̍�ՔZ��Ku�ۗ�N���l�u���*� |��z�\�\۱bwa�n��D���m��S�|�*W���3[rc����m[\�K��q)�1��(+��t4�X��wK��̶�5���ZX�m��('����R�7	���!�}{ը�ժ�7�6�
5-�';1�u����e������F��/��N4���^|tr�3T1������P^N�9pF���W�",a����:7����>#����sU�g8�a�y%:�qҎ�����͹i��61��ntzɴ�Y��4��O+X�]���!k��m�f���@ʇ3�"&�[�2�1�^0��/���	�b�N(t`���V�Cr��ctE�R�l�oC���,
��&#dh�A)��4�v�ԥ1>#Gij�5nr�4CJ]_f8����=̀����7��ƭ�Lt3����傹a?i����A&�6�j�����s�����/n䳳F�#CMٺ(�7&\VwU�/S�/6R�9��v.�յ������NV����e�k�x���� w��PФ���Z�7��ի�U��tu��
���i�e�[qYD���Ȁ���'/�t�s�Eg,v�f�&g15>"�NnsӃ8@���Ef-�;YM�F�R�C�f��{L��HﯱN����9�^��Ozv�1=ՙ�tE���R.��ׯj�cUq-�e�7,�u�.����M+�k���k���$���]~b神3�%{C���Y.�4�qq_e�WϨvN؝�օ+�!)U���k�U�,.nNn�7lRt��D`rs�u9���=���Ļ�˾,e���\ڴD@.�wfd$���ژ,G�6)x��ݽ�(��j�Q�V��jk-�M�,��WJ�혵5���xN�Pj��gvK(��YpR_-hS�%5��uH���sy.��u�`4mHh��G��T�Ul80&���' ��hU��C��Wە��'[@�EsWx�%�ΧSh����Ws㚦3Q�V��f���<�o|7�ò�mS/2� �϶��г]X��q�5�c^��+.������ᅩ���b�_\=(a����r�[{0�vz�7Y.�B�L5F���ffv��SeSS$̮V����r�Ng.Lt���R���b�G�GJ���7@�vd���)���(#��O�2=��M$S����b�#�hJN絍��)�yV��%��5(C�bf�)D�iX��1n�g;6(F���+����%�n�z�6��t�,�k��s�Qr�q(��:4Iv�k�Έ���U�*���Fkn���B��W�\)�:���.ŝ��(�,t)Ե���V��Z5�/�F��$�oL�W-�;*qJڭ�j�����2��<��D1��Y{��"N�U��юU�^?��؂����1���1{� ![�֞+۾V$�����7v��%j��=��]��5�h'9����K����K�c�`��¢:����<���7gv4RA&�PO\ K��V,k� ��f���-W�t�y�y%�Yt�P�͔�'&��h�C�Fwz����2�XNk�����瘦C�eKWD�xpK,HV^;�v�H.��,�󅏬��F�%�5:�5�]q�]�H�f��fɼ&�+#y�;�[	܋�Z6�so&
�AR�R�l�|�(l��`ݚ{���Y�A�I��@_U�J�g�iVԐ�w]��3����9\���J\�&�.���or^���+��7"�҂k�lڙ�n���-J9�с���L'E7�خ
Q��3�ɘF.L,�W%�G���<m�3����e1Ve<��r�ܜ��]������z�qGp�����]����gvT�}�+U���|�K�E����Rf��vR�4��r�v5�eh�nQ��.R,�;�p�H���8gy��eO��qܩ{#ɛo5�:�9�}59n�7Q�{��U���N"��J�:IL���kۭ+0���;�k�51A�Gs�ڞm��Z`�1�9��;+.�lԒ�nt�R�*֮�7;�A�s�F���V. ��8S��UK�H=}˩�qD���/��v��Zy�;̄��J����]��������z��$��@r8����lr����#Y�bJG��Mb�I�ՙl���U.�w.�o&p����:M�	�������Eڅd+����D	N�2v7W�Ҏ�2�$�̒E��掬�V��P��&34Ͱ�=Sr��؈H�8iN1ri�?<{:�k�AhR�Ղ�Dj�#w��.��W�I5����L�(֞�؝s� ���ܡt��*�Ω�Dh3����9p6.nξ��U�ukw7*R��'LJ�[C���n�}-&v�]�k��t<`�t��mF�/�b��à�e:�7M Z��*����[�0�a)Xjs�BZ7�`N�C3�'vR�[h%N�7L�=Ѳ�=�It�HBG������{O��D
�R��Ƶ��w�(�϶ܲWjDX�q��V)db$̝3�sz�<p�FU+�]>[b`Av^*�Y�ʈ�0d;���\i��$&B�d�S�w�aP��|�u޷EtN��|�\�J��6+=��v�������fme�KmV8��޺`�Jl� y��Q�!�McG���:L87�Ɔ�*�7�Z��*◛�m����=�1�x5b2��9Ņ�ā��E7b����X��Wq.�e�=�tb���FQk���(��]#ohϵ��ȵ�<*�#���R��Aio%N9��{N�5jܚ�7��nÙ�&&T�v�4p�p0�sP"�=�3E��V�I�*������i��\�vFS'7m�M�^P���<�S�^2�-�h9�,���̖�:�桉�Yh�v������T$�H%��X��*[�w��7���	բ�b;��z��:lg�"����E�Z�v��s;,�w��(�)h�ZXJ���Ա�\in�7p;�
:����w�,-������W*��v�B���v��K�fe�*�ѵ9WBhv��N�y��SƲ����=/Oi-�"��U�,O�ε�{B�^O*�Yeu�h�QG���bm��hC$L[y�k�5�$+!o�:7�p+�f�.��
��j	�v���N=��C4u_s�D��������޺���p�_8�1e�V.��U�47j�=�^U���-�DVS���Vx�u4����A��6�����7]-�,�q�nJUn>��q^��g��������MTc��y�pa���E���bNN5�y��O����8-%�++�K:��%�ύtQ�����=	�)12�� b� s3��Ҳ�Bd�����A��C�ʙc���V�+T�sݦ+�jG{�0��mJ��zRoe��ۮ�k��JyLjW��P�Z��y��"�ّ��n(īΣ�t��nVe:� .�N@��|����0K��F�,\�3��� ��J2����J��L{�r;�{���t��л�r���\�w	�O)2]]��Sf�'���#��Wq$�)�ҍ��j�]0(�Z�'r��iw�,]�V�D��,��wuѤxݢ�_G-�T���TcK�Z��z�l:���t�eK�mE���Ec�ݮI�5���Dվ8�����KZ��e嫭Į�J��$��
�K���W�;W�92��I�۵�kë!�]\�Gw�\uW�1m��'90���6��]s0��1Y�:ӭ%��*8u&Ŵ*�@�V���)��t}e[&�ڼ���o���b�BȖ��|�Zf�j�M��{%��Y`�ۙ��L-:l����1S�8¥]@D�^��cqݢn���F��:6N��B�"������J��>�����2u�v���������WX2@2e���[��x�k�6����tˌh�:�'S#��P#+Xٛ�W��u�J,�w�4�Mj�ךq���k
�ظ'h�QR�{�"K� h
)ot�6�Q.ᴜ��r���O2��i�7�P�z�%�� WYA��o�-���d�"^Jsf*�r�]21{�� ��u/\�S�6DD�}���h�鎍�g���E�
]�Є�[�z�>۵O�]�4�F��r�'��Y1���Q����{F�;Ff�es�h��t���2���	��m30��T��qc��
��X] �t��7�Pd@hҏ��N�-V��]`$V[�z��}�2���PLRL���p�[\�.1��4Ղ�X<U���0�u��]�wVQ��aԽǋ���T5�S�	7���@^V�8�M���}�=��P�k۞p�����.혰;��1js������[ma���qI�q'�I
��9�"��yF򮡋 v+�29��7��v��C����&�r�4�*nR�^�Fl��L\o{�ݧp̮��50��0���5{�Y��p�R����)4Rt�kp'N� �ھ�r���i�Y,gt�Iԋ:�w��a��2��ARXf9.�޾JE����̼��+I��R �W%�uҗfqt}fEib2ul{$b�id
�t�R|՗�J�-��9��t������k��C��Hu��{Bңl��\�˭��s
Z��Qr�r�l�-�dǄ��'�,�)H
5�U��[;0�"ɝI��*��]�mrK,�&/��ױԤeX9]x���@��W����Np#�V. E}@�w�#(�r�%j�/�s%e����v�[�9����P�٫�M�\4�2�j/��aj�l�&����e{2cF�uل��i.���1�%J��6.{	VVWnPV���JbR��N�<�lܣ8@L���ܙ)}/E��C2_�X���P<��dkF+�:"|d��O31X�fq�t� U��(iU���v:�ٓ"� �2���D�/��[�.����J��;��\0�s)䡊񶫋a^Gp�΁��$��+�v�n�j�u+�F���p����լ2Y�BX#��:��OW���v���Ir���ԅו�ގ���z7�4rB���,LW���VRq��[w#f&ɍ�@�Bۺ�u��o�%m��(5[���4�gAO�Z��s62�Mt���ͤ��t��rp���f�hyWm�2t�ӓ^����a��	��i93�z�U��wD7v.(�vL����!��)���);{�A�p�M�U����np�,iha�oGr���J�Yun�
���ڱ$��O:�7�\�iJ3A��L�9Z�u�\O�Gj�x���Qa!��fw<�jiA��W�M<1�{rh�1<��S�lJy�������-���<,�Wj�v�I�v�EV��c�(CW%}c7J�7{�X���!կ�l�֢n��EƞuJ�ፌV���󥛙��#���$)���8Ԯ��{�n�%����Ht|x�ϥً1\/���t��u�HB�-���S5Q�'4��i	��<Tms��w��a��h;v���-^y�Y����y������! m����o�]�[]r$˺,�5҄�i��s"�_U�-E����"�&��`<KZ4*���k��R��,�@�bG��:��Kd��[Du>�1�}������yw�wrt�M�L��8�-\��J�u����xmY�>56�D��I�r�m�7��S�����\�{_2�wI�Ж'�����&ҝ�X��Y+����h��5�0'(�\�m�(�5KIv��a��Iv�h��l����v�5��f É^��ye@u<�.YWXV���|���]�y]�xel��V���"�!�7r�{�R9÷,�z,�+HI 9`ND��ޗ ��0oa#�ޣEY�|ܒ�I�p���w/uDPy�p}{o�5{��u�׸Rj��d�)�خ�
�9� ����Ue��u*̤�0vPY�t���_�\���[�����"'i�:��sp��ف��TF�)S�k*��J�y��ޢ��^��{#஖T��A��1z����Q�wd��N�[إ��
�ى��֚
�-�4�]�4w*�=�Y2�e�]r
q��VpO��41u]#F��e��FNή�G;��>$��r�8Ag��&F,��9��yBjR��ށN�ՠ�Z/�	4LJoV����ܑl�DP˗fq�q�n�/p;�2gt�a|���'����G0���9eۆH����S�V����!W�iΆ��Xz�����'����iԺ&�R��I�T35�u�vv�f���I�h�s�]f��U�M0_P�<*�,oY=�i�j����w��d�H�pdR��Y���/h�N��AjWGCX`=��yʅ��c���ϻ1E{D�1w})�� ���e]�vL�K�y�U�I<wb��lP�|�Y�9PxF�>��]O�|�`nB��Hma��&1R��f�֯@91q��dA�%W.�[���7]@�[ u�z���=Ċ��,Luw��\�e0��Fһ;�N�
2�^�ڝ���`��7��L�Ϧf���+�	�Q�;#Ψ�><6+J��X� ABhI�u����j� UÅ�7����'�S�$��d�f�f��B���d�z�¥�)dB����^^�w�.����fS&���+��2b�owQ�q͗��ZC	nu��I���Y#�����{mjsV��h�
!8�3��YX��:����[��B6��[��ѭ�.n�i�塛\ƩsFL�%k;E�xr�lc�ҷt�u�9c˓L��k���k@�<�|�A�r�nC��d�|�FEѻ�tv�1s�A�GrK��]H�@0���)/�t"����֪m�d�[,Q܌A|lC9u��E�������MR���T�� (��AQ~���<���w���<�U�*���g#M����^Y$;.���=�,��0)yVx��a�����:�,Qǖ�wf�ć.�;6�d�|���d�<VTJ]��xu�/�,��+���F�j��rGn�����J[<���Of��Af�͝��ܶpiZ�{���b���\Qq�\# bdƫn*�ط�TS�U�mY�OxN���it��6&n�J�ӉW�1�Y'XJ���Un�r ��oL�����W�[wH�`��H*&����Xt�O6t��\t��5H�*t`�\il��A�G1�r�I��l��C��K*5Y@v�䆚�;�W.��V���ш����Q��˩Q�p3}�0h8�,ȱ�kVmk������FnK�긻0�&�t��뗹r�j�O'���3�vv[|�HM�n|�7Elǲ�ݡu+�}{yMaZ�k�����m-ye\�V�]a@h�T�_	ҵ���FU�]\龜��pfk���ҵ�̂�����z@�.� U�b�Rfl���X\9륽XZ&]�4ef"!p�u(���>�h�kӮCx:�ڗV�ӎ�(�i��z��$1cβ0�m�B�����V@n����:a��G#]x�#r��eQ$��sp�[ �T*��b`ܴ�[�vs�K�6���AZ�y��EE�).%)�uĻ�Uʿ�[s��x�⅁m<s��ʖB���v��h�۵�
�/mCZk���Q��.��b�+p쳇~É�� �I��9O|��c�Ɗ.���#C�#\fۇ����1�sV�z�gKT�괰�[�K�Ӳ�\hN+'TDU�{�8��be��)Ð��� ��26�M�iH�1R�3p%�{*WR��YlC��hoCH�J�}vy�Y�ضj��ip��-�U��oD��7�n���ڔL�U^8�ZڬV�9��
�!Z� cm���WX�W��7�1�����(9`+��C~�����0f�%�}��h̘v3��. v��OT <����o�-���zc��|.�Y�&s\�T�u��ΘqL�RV�u �{[b�ɪq�Ic��4l��˂��j�V����:݁�`��ͫ�t�T��9&{����t"��f��l#3�H����;Ź��ZvФ�WA?6�h���1�96_M��U�i[��W�5aYڈ�/��bIB���#/H�PR>�#F��������I��#�N��ܢ�OعڧK!V5�|�SGF��_Tpu������ɀ���&-!�ſa�J{]��Luc��W����H�l��YE�p+4�m2�ˡn��z��e^�ZI�O ��B��H.h]M�'0h��Z$�o|�m��-@�u�ѵЩ�ˏf�w	��T�Cz�,Rбs7,ة\�t)���~y��Z���So;x{�g5 �\�i@k�6�י�L�}�Wu�eG�; Zٻ�$\+i����h��]��s�0=5̀���1�䶢r7��a�S�Y���8f3��Cm���_^P���Eҹ��j�YV�<��굦���s�R:y1ۨ�S�DP5f���f��L�PSj#����c9k��8���;�Y���rWXuwI���Nzv"0��"UsS���{	}���Vi0��̠	uyZ:�M�V%&M-7[��{K��I�h̜_O���(�kU������,̵��
�RᇨL r�-hKvT_dd�	Wג*�f�՛�UĠ]м̐l��)�����y�t89E�s	�oV��v.w���Tl�<gJ�v'2�a��g(-:�q��͛D�n�7[(T�H�9�2)NיYd 'an���t�k<.��,A�Q��M�V�4L/i�l9�ݗG7�A�ɪܴ{|�j��^xWB�Y{f�Yw��ٲ>\�Й�
���g ��H�SoTʱ)�4Σ�w�Ňs#�:���),]E�Tr��)O��rj㘱f��� /"|�%��UM�!�|�i�٭���Č�k�u���q��`�BR��Jd�W���!͟k̾����73k6/C{ L��g9GwWfR������o�x�Vk�CԊ�2���R�cyX���8�v�m������P��h@�[8�" \�v����.�^,ln��o�-��aq��s]�s���.�1.����U4�����at8�M�-�*�v%8R�B��yg�Vu�	vJ}3�Z�%�왧@k@�ol0�/M�=Ʒ1��j�9�4���b�AN[{��;�v�C8�}��i�.4�Z[��%vj!j�Õ�AK������6�V��q]]K}ӽ �:ŗ��d �ݩ6�-��b�G�83ތ�Zr���솙�־8���T�<\�޽�dʹWd�����i{q��Une���5��O5�WB�H������ҵ�8n�>D�1Z2t��2mݪI���z�T=��[n�(�U��j���6�f�y���a�21]eֆM಩9p�=��Da�"5Q�*�ʄh�}b����V���(��3���˞�8Yr��� H�i,JI[+��S���*��)î��w�vN,R����[���K�Gb7�����7�
�\^,ڱ��Y;�N�N�^Rp���'Aq�Pε����}zM9Lӥ����d�m�D���A��-�뱎�v�V
ٵ9Mo[W�uj�"	��2��5y�ʫ�ա��u!�����>P�dj�g6�VcZeN�i��'�G�k�p�Ks/��MȉPyɖ��Y�X�n����r���T�}�ʓ��F�RfG;����'M���@x[f���A�7�::�f�xjTy��%�c��m�)6����գz����A��pV�į�U���g���B�LH��V�6W9.�1��:�)[�b�F��H�Z�֥ѭ�| �k�cfS�.,���/�2L�N�:ÝYP;�<P�1"1��ΗKj�Չ�Ss\��e��륙+/��&��3�u�ZoK.��ݣ4Mʲnfْ�|�4�l��u7�={��`"Z�)%�I�f�*p�ÓX�@ϒW ���+Wn�I���>H�f��q�C�)�m�m�LjUzFLB��o>x��W0mE�����cN�ؼ�4�aP($뮸�=\���`FYw�6ƺ3���3�p���)��r+��+R�Yf������!>QeAtRx��0ٮ\�l�w��`�g��存�l9ϲ�leh��������@��򶌺�*�x֛n�B��e�t�m������T4_\3FR��V�U�M�b�*������.�wY�	!�mY�ʙ��F��&V].�����\
�#�J��pxrg&��C7B��|+��혊t��A}�E��c"�z�{�U�Ք��u��-�c�;��Uyemq]�1Գ�ؒ¦0�C (u����̕�P����+�lm�E��3\���gL%L52�Ry}VD�J���	�K&�J}�h��tL���F�ε	z�m�L��_`�&���gk���2ʷ��q"��StR���nm�rS�ļ}�+�Z������RL6{ 9�;�2���'1-N�}�n;z� �5i�s��ѐ<!YFI�t^�b���Đ��U7�s-����������W��L=�d�*Y�왺���:��tn1��8�.$BO�b�b�ݦ�\hm��V�Sy�$�
w�lrݞ�.Lвt�[Bfe�-Ję��W�ݰ�bndY|�ܫ���x���ʺS���lԸ�	��h�3U2��&���,ƾ�]�k�휓�������*�o���ŉ+[�Ƴ�����H'(��m��;+o2"�-�e��k�[ղP�𵕸��4�"t�!K��j�Y��6b%6{�9xoQU>ؠ����X#mr+�d�RFD �B��V^5����]��Eܓ������⚢�W� �[�A� $؅Q�N�
�V9�b�Q�ݣE9�T���w��y�ٮ,WUݿqp��v6��t���dVw!��]�HRO%|��c�s��ƃ�e�y�)�C+p��=:���絡WjX���&��V��w�U �ɣ4��1��kOD��#��RY��Ь���Γ�q��%��=Xɥp���r���Q[��o�����"�:���f#h�fؕ�>�g
��G�o�R�IEZr�����5b�r�� ���ݖ��{��ƴgo��v\�m]��{G@����c��/��7�:m��o ����
�ж�YV��tw�t�.�+c뫬 �7R�[�B�>�k�|q�x�L��Y����mr�}�w�m#bzЫqfR�b8���y���c׮ƱJ�%z�m�HX�j��fl�b�#�K�@h��X���k��9�5�R)�
/c;�@NVyl�Y�`V�ި�Q��yu��ЬJ)��ڷ\�\#�(��ֶ��A����2ƺ��U����dd��^դ�� ���&�#l��N+�� jpp��N�}t�����U��s*>�]�/gm�I!r�,�#�3u'��rTU]��]�ud�i9�]WV����j.�P�:O��ی��Rp�9�6n��5enR��ξ��
��ɫ��%ee]\ #�i�l����/VS�Zx:��.%���]�F�=�
'5V��;SAJؓ�*�����̀nL[�i֭|\���6\ȱ�NbՕ{����G�3|��O�LyjȂ�:�1VQӊ����sbJ(vQ�p�J1��X0';��q��ܾ���K�wu�|�<����0]�֭�I�W{W�ƥg�1�p�J�0uv��YͼE͆�	�v��W�ܛYlf�k�Z�_u!�J��,����et'�9i$�Yb��&�"$����nT�F|b=y�//��^��2�e	y}�c��;�*"*��r����-�H@v=�\#t�����DG[��w��_ij�<4֖���-��E��$B�Y�Q*`��WR��=(���7gx59Ĥp�{�b�/�Г���b��ˈơ�镮������,fȯ�Ô�T��2�H(���YV����1�󅞻�%+�^����V�!��[WD�g�9l��|O������גuܘ�Y�E&
f�n�lh0�;����/K���u�3F��w�Ӂ/�.)��^�������%�tc�\�fm�����r$v�te�j�j�cx����,�2�g�kamm�#t��ݖC��R��g��V)5��@�fJ�q|��
�{�xXT0f���� u�C�ee	��&]a
S�/��W�h�⡧�/�X궻��c�ӧ0�ف��3���;L۬ɚ_Qʁ��㯯0�ֱȢ�a�F��s�P�2��q͍�"Z��歷;-B��lU�L���is��J4h��tMc�a�a/��X�e�\�XY�A._[��3�q�'�Ι�)KKɕڱ�L���(�7��-��gRM�+Lo�����Q���:�cX-L�Th_Ȍ��R���E����uI���2��P�w��ɒDo�ʋ-7�UhN
���i&/�9���P��X�/,9)B���6%S�m�)o���"^Dz���.���M�fm{p,�/�ܰa�5�6�S��i���Xk\���4�EVMͱ�����fI��K��;X��
�kn���]Ӽ�(a��F ��&N�'���Yh]}ρ�!v5}��["�-�*
�&�0i�n�J��V+T�[ŚkV�ucn^�6��3��֝�E/�2^�d��0b�-M��8��m6��2e�N�*+䦢��2�� U9wJQ���j+fD�M jnJ[*Fp�-��N5Y�2�ۑK�dd�X���ˡi*���R����8�1v]�Q��94�u�
ي��v"w]Vj��+5
�i�H�-b�Wu����#�uY�y���%-�4�]�e�����)A�o�\ݑC��ַX�ën�`R�]�;QI����39�:�͇+Wn�\GC�uyU$Qs;���F��b&ۭ��k��'K�䐼�9N�0�er4����sL09Ε�mP�CK�>��""IG/��$cVj�pWO�����L�*Yi]v�o��0�sh��ӝ��T���ER�(���2gj`�+���Sm�T��@Z�mqʷ�R���tO*�}�}&C��6I���ib��сj
ڎ�)��1!8
����&Y�����+�{N�=��b݉��ɬ�[8F�e;�4b�"���vv���"V&�ڪ�'���C��Du4чSV�eL�s���Zf��:����6&Ф�/T����˂*�,j��%!�(]`h$�`�}|�ބ}ɣ���}1�:H�.X�5��f��Crcj9�+����b����-���S�dd5k��	�7�*�k���D�����rԫ�L�W�����[X��h��fM�Cm���
ڴ� �� G��@-m��ss�H���d���O/�j�I-�WX���w�5+�`>��=G�4Lݣ.����g"�)�a�����p�)�+��ip�x��u����J�:���=�'f#C966��]Z�� �S[�3
YA�Y�#�	�݇�w\ˮ�Έ�͟"����.�]Z�[�6�,j���\�Hz�S�ӊ]�/*B� �E<�q�/����Ȇ��#�لG V3��#,ˊ�u���b+r�y�I�I�����wXN��0��d5�
�uJ��&��X3��s�!��#�*�3��,f�W9=���:�Fd�-fY3�!�k�eBS4]��Rwor�F�"W6�;�:8)�\(m���&��FN��}Op��c�TL:�����a��O1�֨k�	Dݾ���H-X�g%�M^������eW>��B]��/n!b������z�U�{���xθ�P�qK&�m��2��.��kwj�9@π��\���M�����ov=(�p�Tq������:�m^=�]+�:]��VZ]D�Z���]�����Pu`^�F��д��o��Gc8�t�;�5&���+ .Դ@[��]�щ��ǲ��(�M�,�/~�ٖ�VN����ܲ�;D�b���c:�s2��w�Q�v�Jy�n
O�&.���>C�it����@�}��<�5s�Vo��CZQ��r����ط���8en�Ry�L�G�Jd4e����Cc��p����Q�x2�^D���n���h��fD=BVZ#q�����Yj�3�G^6�	��]��NR�!�)�<H�ڛ[W�/�����ne8�M(�Ŵ�ʲ�V��\"�ыnc8���]:�ɝ��&�n��q3M:��.TpV�.���^��XA�i�=i͢N5k��*�Ayh�dwG�����&D��<��^|էw,�`��J뿵�V��.��!���m���
k���mZòR��f$�.Yq쮗�Mb�_t�--��K�sbj�FΞ�N�u��-����[�zp���J�G�{x�ݸ����mR -�
{��2o.̦5H��p%(�<;]4n_q�d�x�Z�1�r�4����J�a\�sL�cxҼ�˷r氡]�3�\�m`�s��Am [}�˙FV�!�U�	E��o�)j�*ǫ�/��bħaU��v�u.e&(��Oz��l2V浪��'���w��a1��u��fPULTM5U53ADSUDL5�I1TTŘ�A3AEQUTP�T��UMQ5P�4T�Q��IED��A�UfdVbd��eDDT�-T�3TT�f`DUD�YU1Ue�DD3T�LKEIT�U%TԕLIE�TPLQ��A4S�5DUA�KT4DEPD�TTUIRUTSK5E9�0AQTIME5PP�311VXTDE5UUITՖQEU4�%��USEFN54SM45SQMQQ�AAE0ED5$D�E�PLLUUQ�D�D��U$UD�4�Q�,S $�A ��.�SY�vf�u�+��m�+�����dɜ[ObC����H�)0	�g�L�5vT$K�y��a�޿x�\��CK���t˼�i�\��R�,�/�K}R�U���쉝f�Iw�%a�y�ng�'4��y�g����M�g�mh�:��5�R7B,�Ȑ�!ժ:`T���+�8J�mf8���O\�J�U�m������xlػ�W����Xp�ձZN������L*_{��Z"�^:�R�v�����H��|U�$�R�-�O˴��Ő����wno#1R��/:�:rD���b�Xr��9��Ra��1b��%��l���5F�<Љ�����;~5���	�&
�7�Q�}��^/new����U�:��~j�I�=Z.?U�u�h��e�:痦�s���Y١��/a`yi��S��PO��;̭`�n����F�R�{.wCس81�����gyc�w'q~ͼ䲩�6��L���6w��Ֆ2�cֵd�NM%�U�/;�M&��5��{��j��Sȼ"�:z��7�����d'q���̷���$����Kt��3�ƻY���?vN���=�A�h�p�6�W�+W(b]�x��N�^ �v����[�ZzegV���o���y���1P��1�ғT}Ĕ�M��c��^�e��L�gu��.���ټG���T?b�Y~���������@�؇��x���&�L��F��P:��٤�bGE�oF���r�Y. �8��{��VQ�Z�}�Vj\��!��)�X��y�j���;��9�gn��]om�[����S^a9�3�AJ�z'.L��h���y9�=Q0{�8ǵ�N�%�aq�y�I)���i	��p��{MϪ�r7	r䷤�sd�C���O^P�O;���U45P)5�¦o:��s�W�3��m��Kq/t�N�R+k:��<��:��n��^C:ENPf��>sWf��;�oS���.���E����X-�sӬf;�-hZ3m*�Զ��u���	
�J�=@6/Y�y+��P�쾵xꭈ��V�oZ�C&�x��ï�+�����ĩ2�±_�z��7 � �g��+O4|D�����ާ��ԫ���6BmL�7`5u�*�����䉤q=��D�R&���ĥ��2\�\��Hf�,�I7K�ݑ9��-�<t�[dK�^&G�|�_:I&D�-+����X\�:��o� �������v�}�ܬaebv0vt�׎��itt���0�����ݎZ7��K�Y��=N��t��I���ߚ����o7���e���	s��5���P�]^˔�rX�q:�	���\��]s�ۭ�ܝ�O�{�r�ũ�.r�ܗ�i�&��^yFe��{0����>���p,ۘ��T7�V40��J�3=�[x�u�mp��IK�m�՝a�ǹޜ�f�Dnӱ94��4$^&[�9�\M��0N5�W]>������J�����{s�3=�v�➋S��H0G�|��i�K�I����O>�ծ���V7���	���Wz�B���[�4�[[ڪ�_`V�]�SM�v�bT�t!�a��.Len��$ޮ�������WPQ�*v�==@F;ir��Kb����{(��-nf�m�~���p}W��!�@/l�<��˝띧C9=X����hx��s��87�a�+�.�@خ��Y�Z^ܬT�0������qڱuL�S���Z�"T�ܛ��,������j���g`��B�Ӆq��:>��W�)w)�g��ԫ�?%g/�u��q^�[,��uyZ�tLW�w�X[�{�Bzg��w"㔪 &�&C���BۯBڠZ|v�nҹ��ץ'֪��q�Xn�)y#U���ir���S�tD�-�-j��r��β^��ύ)�psw'<��!�`�d�S�C���Q�|��.��c�X!��>I�N;+��&֙q��8Er��׹����DmJ�W���A��MI����Dl��k��sV�WF�]Y9����9��_]Ȧ�e���ʡI�(:�V�!��LM1��v�w�V5�Zxs7���=��=�X�{$.��|���G����3~V���ͽ�$��p<7!�+�$4�Hc~��� ��3�Գ�>�8�֍*�Ms���}os!#w�3X-9�|1 ��������:�Md�c*�C9v6N�"!�-eM�w^�[ {���<�:�s��:���Fl鵃=g<{ϗ!��WKU�}�g�t�׺F��Ҡ���q3�[kZ�e.�*���d�A�:Z�+c��>E��n�sR��m$���w���k�3WH�����x[a���l��dg5^U��яh&��Y���9�T_�w��$z�T��T#U!r���;��n�M:�B�ohYTv�Aw�z)�"ծv��L�Q	��j��� ��=���.vʨ���W�Q����yݯN ȝe*�	+n�r����:�U�����Ml����������m��F|�]Մ�K��-{���ʾ{f�%D�4!��큹���~�]�*�m*��=���+n�[f�A�/��A{�y�:+����5��oe�}TS�Ÿ�n9sB]6�-S��@a��q���{�oVb�ԑ�~l�>�52�����g)^9��ph'n��lR1ј�hw����ɛ���Ϳ)�ˢ��!z�G�:fڛU{9��0ç�\v��tncB߶;c �7���=�>�0���RKb,
�<�v����km���{��j�j[��&�Ȏ��Ю��Y�S�����-̺V���:���;#������H��A�y��
g�a��56��i�Ѵ�F�9o�(S�'\+V֫�i.�u�}�n��X�I��#�u㜌�vlh.Ա���R7���b���6�"��T�ںk3����eV�)���]�u�ʾA��\�N�>���V�`r���m5�
;*�����pW��i�[�ũ�(<���F3�,OM��f4��s�����`��o��}}j��ypڛho3�W:i���dL�L���RW�ћr�s��k���	�w-_�&��hu�f�q����G۠�8v�R5:�y�R�T}����Qnz��M���z�����sS`�Tk݊E�K����j=s�V��!Q�v��Vȃ�D o	�w`�u�I[r�zV����&9�׎;�Y�Z�Q �
�)x���o��ˋxn#2����v��#��[
�{�B�SZ�����԰���``�7��r�5���v��x�q����۵6�+���Y�M���ʀ8���YJ�#ݡte��]_��e�ʑ���Ƌ]**��Z�cq?�� ���_D59�Y}L��m�/xT{.ݞTE�qEQ�`����\�C�4��%�0��EY�w���W/�����	"T��J�:�p��HT+���DQ9�[nƋ�R^�:�-M*��:�lp�e3˺uD01y�a�"�
���j��W���$�38�����D�z���_W�a�؄ŕs�qnwt/J��
A�&-�a����.���odPT�|��hk�nelH��-]qR"�G*w-��o��%�T�����41�&X�<�\�f9�%ʢ{Mu�KԂ�Sݪj���89	0��89��!�ah�پ��9�E�o��F��ᛇ*ߌۤy ���<=�S�Z7���=jp���W�$0ڮ����T���+�s�r�0]6+{��I7w�t���.��绍+ս����D��wr)���B�4-3���r�a�]Y��{X���9�9�ː~�^�l���>yT׍L�GP�l������sx�;9��&��9����a�z@]�+�)*^���c��΁e�8����vL�}P���ʛ�`T����dn}$�'�e:�(L|5uҭ���i�RVd��x�<\����3H��J�\c0# ���T����2D�R��[S���T�Q�z�I^ �D�+hG�k��<\M�f{_r�2����z��M�N�i�>L=�з`l��7���R]\*�	�#�ԍVء=*t��ю�B]�8�y��;B���6���Y�r����k\אq���*6"9WD;�')ױ'�pҽ���uw��n^6�j���N�Yn$c�d�h���[-+5�T���]ګz+�!��w [��"��Ei��B4�P��+�L�9�ٙ�Y���u�&�����b��s����Ρ��u��=���!sCK����t
�w�����Wr�e�j��q�W�́���R��Z{K��՛�j��単��Ɯ�O(��T2�+�DC6�d;��$�>w}�+=;^�ٜ0�����F���l)���̚0�dw��;���]�#\�	a��+	��t����(fX퐍���M��e���1���zNA��~�������ڴ�����0e��%j�RY1i�g����]���*����9H���ܖ.���it�Ɩ�wD=8��րR��';�`�Bt}Yl�2�A!��46vk��;���W=w"�yC�����K�������-]�x([�G=í�eX�
�k����J¢��Mg-�Y����r�CS�y���%�ށ죸9�y虅{R4������d5��X��ym�ϫ^�y�{�(^��\�a9aL^G�7�ӯs����씰ΦiOZ~�\g���s/��f�v�7��G8����|��x����v(_�T�HG�;�t
�n�6�/���W�.�b�[���C�rq����+���� ��{i\{ڨ��2�[J^s΍W�9�S�|���p;�=�hz�eU��'g�dy�I5�]c4�}��]f۪��;�����um�~�^��z����B����#�za�34�T�gk�\�	�ҧ7��9eZ�Rqo�X��5��q�w���M뿕%״��z��g�x�Z�*Ǉ�jo;�'�-���@`r�/��ڳ;����s�$�O��5%��-V.]�f�r��ov!�bsU�r��D���&�`��z�h��*�ɀEz��#�_0cE��{C2삶0'[� �{w9��mͥOd[��!Lz�:q��Nu��7���~B2v��5&���R�7��|���{���2�3���{��>+�%A�z�8��6Պr��!�tv=Oc�gv�.�-�j�^��>�.�n%�ؔ/��k%�G�gm)����l�}��� �$ħ�k��A�V^���3��7�[�;�^��	�ɛ��Uӱm��Ns���\meF�o��m��S������P��$7�_��
�ujF=�C����3�8'��{3-�^e�ۥ�i],�J�|����#8�U���^o3bi�M9�*V������t�F[�7�Ձm�z*Nu�𜙤6}MS���Y��x��,����}�f�:���7ܴ�=i�����~ǩ��z��Lx����v.fI�Jˢ;s
P[�v=<�["��ֶ�Z]��B���[��2�u�����v���	�'��ג�7��j�ӗ�#��|e �0|V�C��j�P�袸2�U�����-%��m�'�D���y]�.��n�8�Z X���7xa�]"��"�oix��ZiIc��Drd�>5��+�`�V~����vˉ]���&T��T�SN�S�޵�8�t���[r�X�:�:x7[no^�����9�nŋTw&��A�5:+�2�\�2��Ny���6#�wP�iV�n�;2�8۵����Ld5b��j���9�[]]ͣJ0��UsW�t,f��J­��3���)��Z���ff�k�Y�u�.��#v����5\\�3�7��XË� ��>���|i3N�>b(.ˬ����J�v�:�[\Õ���6P�gZ���2�	��2�\���t�����Q1u���o�q�b���������b�C�w�2����"�Q��;"�]���x��,Ըl��Vˠ2�	B�a��Cj�ʷu�AOVv�6e�\Am�Mh�"�71>�oh^���Mӄ��̆��^L�x�n۬�f9P`T�y��٬jTݝ��/�"q�L��I�J�8�ͺ�dZ��,��ZԒ�#!"�jҳ�01n��mL��+Jm>]�2&W�iH�mgnS��E4�gv$&�Y��\�����+&ƖΡ���[0?6**���]p42�c�{-��S%4�۷��:���n�1�a�fglu{SI6)|(��[�u�9@��T! s��Q���^FŃ�+ ]Po(Rv̤��O.���o-*k�B�^ܽ0�|Z��\p�Z����/f�Zy����тy��x�P�X؏򐥆+W�� �hի��,ͩt��j+A��}'L0O�ϑ���_�HzVf�B��eq/+�.��8���f��5�����&�;ls����w*�j��i�>TR\w��Ӝ�r�@���� |5:3�F�n��f#cWvСK�f�����Q����vaz�J��U����DDƤ��䥾Gv�v��P��+��4�hR���\.P\-��sY]�����k9RV]H�`��t�0�V�h��u{������ .�N���E�Ѱ��r����Z֌e"�QE�AmU�U����f*'wf�X�V�cp��ދ�V�q��l���;�M�/2\�GatbB���("�q�z��r�U�y4�yn���`ьm���]I"4���ZW�o��痌�:V�/t�Yq�,��T���5]z�Z7����0Q�6D���U\���6�7UuUz�B�JiS8�@
���y.����'p�f��\�� �.�vޕ����+A�Q#U/�f��ba�7Y}�4���g��CR�
�Z2F0VT�Z� ���],�"�i>9����Y5(��V]w�u^{�P�5QJ!DITD��BEDITPEP�QDĕQT�QETDE4!L�P�ICE�ACTSA0DPPR�%$UJR��BTBPеKME!MT�IQ̴4�S_�	��Z��Ȣ��"ZL̊�%�����C!))i����3���
�0���(f	�)�*
�r2)��L�
B���iih"�"������B%�c0�� �����j���((*��"��J"� ��!L�`}� {'�GfH��ԅҢ�u`yj��K��+٩IZ�c�6��ׯ4�.��4���u�(A����� ������yMt�R33td�8:��H�k�X�+/�gQ%�S��������j6���˩���q�v�Znm�b��1Ѡ���姻Q��'ꎩ0=>���|��|��q�
�tJeH(�|`r�Qƭ��ܹ�4��]����t5�a�t��ܦ��.rs]wl!� �ⶮ����̄�$���[�(�}���nx^5U�r�HL�\,o��=��a���gy,:sж�3V�}Ep�e��^�����N��rw[�u��	��I�6�%lU�ڢ�Ӧ�3iT��G;i��B��ܼ�ڬ\����O:���6�EN%I�^hk<j�le�7G&�J����I�/h��>|w�Xt^�w��C'N(������ީk
ټu@O�|�}~�/�{r�a뎳CX�3�ƍ���s2�ۖ�ouڒ�Bu\m�M��*�ܷcrP���L��`��[O�hs����D�G�y�Ssl�E��G��C/,���
�n�d?�m�+j3�^����Z�
���Mf;�s@���IqTs&>�D:Ꜯ�fާNW�����4���F���{٧���_�j\<�ڟ�����(!�����^z꛰P�V�����G���7�{/Vs]j2:5�F���"���؍wFv���Rɷs�z����y�[T��듬�}���7����z�`l���>d��~:o����.F�Y��acS2���[i7�=�2e����6��ި�(���-���%ʡ�2E'ؑ��j���X��wuZof��֩(<���'	�ו�, yLm&{}�O���2����.;���qqT�ƹ���M�e:��m��2#�}��%��=��(�h���ґcx��JRjC����lp���傣��ީ�e�˪���h�c=��ws��}���`���Hn�hu@�w��1OIo;s^b������s���)묫W0$sQ &CXt�m�F�Q�W��3+Uf��V�K5���|WD�	�9^h�e��gJ��2�]-����u�:�<�9��GZ���;��*�ٺ�R滊V�=���b�Ǒe� �5�SUf�\&�/@d�%Lea�+X%pր,��粣�{v���ܥ���7���;Lj��^�.1�Dm.�j��L�O`J�	��Av�D]�z�S��`M��;��ΚG)X��F��|�b�cd�WKǷ�w�ej��دu�S�&{���r})D�Yj�ʼ��A&u�;"�ut�����)�j�i��4��)�ttOP9W^��iү�oJ��9��y��W���[�=Uy��dH�;�����U�]��즃�����ʚ�|�P�j7�oX�>�~~�{�٩�H�I�tD�����Ŵ�2�{���;�{�$R�ݺV����(��s�CS��ͽ��v��zr�����^����mf�}����ێ��OFjF�[|��9WPy�����Ѣ��y�+o}J�؉
&���@��=Ƅ^{�ϴ��Y{��(��>o�R�K�q��&���=y6(F��!S;^��"����ij�އǅbB�.�*��D�&�7�<�-�B@��U����w���S�ʼ�� V�9{V��l�p����v9�W��"Uy��A+W��;N�h�n҂�E(�wum��L�^B��v�}��ԻW-�NK�%��)6א���w��U}Nnx/>Z�����/�Gﻺ��%H{�!�[b��|}���e�}Ζ��Oy,�˻rv�or`>�Aas�c��J�wbG��U����p���r�������ߛ������M]}�{�K�<G��ʏy�����>���>���2G����y/�����������5[Ʃ_���ђ����F�������u���K� }��L�H��aǃ�Mu�I�rGq�X���Hw�wӹ_g���p��������po�:�� �pH��Ib~=��e�כ-J��}�����!���H}�/F����b�f�9wnoB�C��i}�ܝ���<���}�r?I���4���ﾠ,��}��To�~��ם��P���}{�4u�߽�u/������:���\��x�$�x���GN�d��.��_`:�ֹ�?Jv���^�ܞ�Dr����| �������F}���~�'��GQ�xK�RoC�}��;wބ����Z3�Wrvszi<�B��ZC�r�^��ӓ��4��s�{ G̏`�����v����T��A��<���B����r�y�5��Hw�4��0:>�亓�}h�K�}����G~:����-�x#�z�}�_t�9�o[��bܸ�{�u��=���>�y��WG�hZGA��9RF�΃r�������09�C%�|9�{d/%��Z2}�����"V�o��m[�r�J_��]Hkx�H�'<އ�>��� �]�v{�伇�_}��;�ǻ�s�WS�����Jsx��w����!Ha�sy"��!Ϯ�Q���v�]i�j��H���IǠ�Y[�ѹ:e�!L�����l*���.�����+=�>���<�΄��ޔ��^��$��nԚA�ݬ����O]�p��6d�a�(�7p�w�U��N�DZK��&89��=/H;�/���b�\���kK�� zO��9	G���Sw�`����W�;O:��y߹��>�^��@{!���G�������?�|8�i���?}�tM�ʚ��}���q])�>��8@G� �Q�c���5!ַ��w/���u��R�w�%����J�w懒�)}��?HD�|=����r�����?�D�
�Jn}��쏒~��;�e8���d?A�z���iJ��>�����'��<�ǬS�:�����W�<�qB��Ͻ�G�n��ʶT�5���]u�|=�����οiO���m���N�?Jy�iO`�{����ѩ?H�l�:��N�b~��K�k�/!��C�����UD_�V��o�+�g�{�=�3���}�C�`����}�S��o.@�oI�O���� jN�u������}�%�>�w�~��|�L=��[�����8�{��c�������� ��|�y��ׄ���p�A�������D�ty�u��_�俌�>���Y�#���� || �[`���g��>;��>��fK��y��%�);u�~��/|֕�\�/�;���}�rC�7!�<�����2G[�^ߤ<��7#��#�I�.�:/�%J;�"~�G�{�p]A�8~�FE+���E)�b��b�f��z;��H�!ۭ�{���;�K���;��r'���>| �x�������h~�qҜY��y��8�C��p�|�~��z�p<�%��4QJ���K��r7�=���I�_��<;�C����X����/����}��h�s��g�y�R���:��}��N��{���M�ԽE<�zSr���+�z<٤?fֳp��亗r�깊�g��?~�}��$�v�����r�hLm�<2���쿷�Q':~D�*���ߙ+����!Gb�=��gݗ�L�۳�/*Z�L�ۀ��U����孹�V<Ppd8����=9�Z��21��:fR[�tW+cW(r��s�&=D,�8x�a�]�}�� =�.�i7�������O�������;:�}nWPd��A�/[擩|�O���}����sBP�{��+�:9���yv����0�/���v���;c�߶yqK'~����é���M�S�=Ht��S�����_���7փ�J��_"���iO%�bu�4' 5��k�}�&�߂I��;�� 7��27�n�����_s�_!�NJ}����/�rS�p�NC�����Pj^GG�hZ^G[�}"��v��=�|(/�@G��UƋrG�����c��~~���!I�^{ђ=K�P����X��<�eט��=;�/s�#�5/'���/�z�q~�J��?�A��z0�W@ʴr~���>w�j�	>�F)�{��=�˩?s��}��-@��4�?��NG�X����iܯ�v�֗�r��]K����^��t�}�b(�c�t�+�ľ����@y���x.����tK����O$�:��1
C �߸P9��K����|5�{'���O%}��δ���/$�_��ݿG����kԗ1�u�~��P'���~�#�q��7�#�=��}������~�Pw�i}��<���2_$ԆA�O���ް`(�ӹ���b"�
����π��}#ߢ���=�r�1�pI����@��}��䏲~�4���9�����}w�x�{ h�4d�Oқ��R�=��y�wԒ`Y���Y�|@�dz���4R����zJ�v���w��A����sԧ���oA��C�HDy#�Y������Q�f����7�m�\��o}�u��q��Wq�X��<�������Oa�^���w��y��ߺ^K��07	�;�G���7 |}~��2�#�3��O�R�퀥Nj��7�*�h�ȫ��Q���Qcn\[|��3J]��U�.Xk�)ˣ�n��+��d��!궨�{i���.���&Q7�u�xZ�j"��IŁ�i|8����m�(8j�6�ݣqgZ�]4J��ϣ}a��ͬ��<;�&�X�z`�{��Z�W4�a9�W˯��$���'�<�H�MI�9�FN�w���(���/�$w!��@}/�������>\��}�܇��~�����u�w]�\��$����}�޳��y�iy'�u+��5'�~ѐ���C�P=9���/��@}�=������|(�>G�ڵ����K6k��
���8��1G��� i�'9�'�jG����C����K�;����s@�I׼�E+��ߺrн���/���`@rN�����vg3��ֹך�����]��C�}������>K��_i䯳����ϒ��s��_`��x��ʝs@�K�o�2)dz��}�����y�{eOR��&���~���<�r�/5��'�w��$:���'��߸���=�o_���n;5��s�f�΃�}�����?��E��� �m>��GUU�}�n���~���W�;و}���u�>�/%�:�܇�z;�J})��4{!ܛ��=��������dto�' Gn�>G��G��Oꍇ!dď�V���߷��P�/Y���S���ѝb'_}����G~&���r�^��>��:�����&�;=��N���B�Br(r�����A3�!��}o���;*;3�{��M�+�����C�g�i�=�Y��0N@j�<��~�EW�ZC��{���&�u=��܏^a�{����ҭ�s��Ov�ھ��{p=��B�Og��G���4�!�b���/��O�怡5����K���dO�;�5����}�<�?M�K�tvj�a���5}����#�>�� �_�K���;��v��@���ރ�⺞�|�~��b��sG���ܞ~搥�to��S$>���|>#5?u�F���ܾ˺��ܒ�1��!�;/8m��nb�69��@���R��C+���d��m�l#ŀZàb�B��-S�M��v�R��|R�·���7��H�/I8��]�+�J�fg�ں��N��*����R۳l^�h��Ry_u�� xn�pJ���}�����9�䯰w�}���=��y��y��a���`9���^H��N��O��ѹ��w'���>����6��\���{\�W���u�X���>A�O$Ծw�?�C��Z^E���r�?@n]�����oO�!~���4���GG�J�ӵ���Ӌ�Τ��<ϑ�����_/��K��	�X���_ ��`��yJ��|��)�a׺_��b�����:�zS�&�����$UZ{Q���إ����4�{O��ߨ9'����䯚��h�?H�=�������X���_"��X'�y/{������W��w.���y��|T�9]ٝ�ѯX�#�t���EGz�cr���ޏ��~��<7�rGrua��PrW�ތC��S�a�z�Ȥ��	���5�~��?o��M�B�/��r�����=�~Ǽφσ�z�}!�|�<��99���/�r����S��5��ܚ���ӹA��%������Rk�/�mU������w��>��Ͻ�擻�^G�b������rs��>~ރ�d�\�G��_'��K�;��9y�i��>�MR�����w�+��*�������R��\���D������=��{��ﮑ�'z���9#��O��Hw���W��u���2G{������K�;�QO���_a����3w�S�Y��^�	�7���Y��f-�9W���B�C�؝G���P���{�N�i܏�r3�Aܬg\3�������=�S��x���_G��� ��|>+�=E=��5.��k���4?����n�5K�X;��wy��N���d�/pnO=�=�K�|蹘�S�n��s:��%@��@�ŗ�r���v���lR:�j����wK�+wj�v���c���;��@U� ŭ'f�B��S1.%m�t�Z�V�����̈́��.�a�d���74#���˵��+�.�E��&%Ԋ囕�5QW*R�� <=�,�u�k�Ͻ�>Do��G�W�s��_b��7��C���}�N@jN���:�~���4��^y�!�9{/]`�����p����}���[�T����wf#��s�j��/�Oҽ���8����L���+���h?K�R������r]I��ѝb<��>�I�{#�5�?A��/�w}������v������=��N���9/s�|?bjC�]{����u��9R���kA������M�^�r�d�޽���������m�U�
�-��A��8��H��4���.��܏�s��{�p=���K��>{�K�^��W�`�ø���9�+��0�C�%9�r�;����k���Y�3��/fq��|�d�d��(t~�g��I��u��>�מi䯲vy֗���s�=K�����y"��z�G���x����[��Y��D�}�7���|8��{T����pxs|�K�}�E/�y!�K��>=`>�Rw�t��L�u+�ߺK����7/3|�}��׿s}��h�/����N���O#�N����~���|������t��&�:��=���u�{R�w����z��>� ��,������f~[���<��~���!�b�����9����9=��?�B����4����S�y����ܝo�����4�=��&I�K��C�C�z��}~����ǽ��w�~�ߏ}�
WP�����W�仇y�i��<���y��Sr��z\��;3�>����7�Կ����^��.}�G�G�P�Ag�VUcܯ�~��C�^����Møz;�G����b�^K�;�	�H}W#��қ��vk��w/�r_y���.���#�D	>K(1m�wH�����j�c��肇ea����2������/��r)mӭ�V�og�9B�Q�+	���;k#n�[�S7#S�lƠ��L�J9��o����#ɭ�+.9E�{'��!u�nt*Fx��g.ģ;e=��_}U_���H��i~@D{�}����I�"<��K�Rd�9/\֕�_��/و�s�_��9!��r���;7�Bd����#�|��.����V�O�?j�r���k�����wP��$��2)]���4R�)N�1�?��1{3 ��u��t��;�4=�B�<:��N��T}��O����S�������g9����2G���I� ��y������3����y��Wpto�/��z����Cٚ�@rMGg���|�����"��N�g�7���?s�oq>���_#�[�N�O'�`w>J���tw	���o�'!�^���sΔ�AȢ��>��E/���	6}����G��p~Ϗ�n��\�[��[G�N��'����y��K�vu��+�=����B���;�ڄ��zNC�^�����9���Zs���υ���}���ŧw(�}�����;�=޸��du�{������@��샩������'%�:����d�}��E+���O���_s^�>�Dx:��� I^�u�S.���tvR���?FǇ��� e�u�g�~�#�zz�ܧ �����7)��G$;�rx~�(5/#��k�:�#�{�r)^Go5��_s޼������}���>���J�r���$�zL>]#��Iַ�FH�-�:�@�?��y>��^i7���^�r=�ޏ$�^O!���5!��O~�ZF��t~�X�2���-u��_WBK�,�|=߼�9/��<�w�]I���B��>�yjG��f��������z�|�e���;��5��9��$�]�@>��Wmeέ1w����oW���+�\=��>�r?o�`����t~����a�4{	��px~搤2.��E���_g�>I���S�����������X_lg	�W���|Om���&WmcPxi��ù�!F��g,tʱ�t����B�b�p5nU�v�w��g�W
��h�xȡ�R�`�"iX�^�Th�Z�Zj�BO��I���t�.���v%����z���5�b ����ݱ�梍"��Q͖hr��>XI.�>Wi]��&�����tia0��1�q�l:J�6�P�Coc�v��%'WJ�'�͵��ꛨE�u|2��V���Z\��Ea�m5��p\7����+w�G�(v���<K�+�4�RV�Z�+����oQ/�U�v�+Vj���ڽ��ݕ�k���ԥlӴ��h
��z�dV��H�ˢ��2<�O"��y��7�0�އ��
�"::JY��P��1��R��EbV�o��6��I�b��T�F�$�VkBE��ob��9�I�����G���nФ��mM˝Of*�:�K�Z���D�	m��n$�����WR����C���)��V��C�b��h��؝��)V�l����R�W�F�P�3�m;ٰ���\��
�8U�ȃ�R�]��K,���M�v�´|)�v�5ܕq�rF�Yz���VV@ۼ�C�nj`Lo���l��B�u��t��^a][��Իx�LY"7��S�ă��y�84gJ��1e$t�P����i�2�d�J;�:����� BX�6�_9X�����'��G�+��B������
䄷,9�Z��6k;-��+^�vb5̺�D���'VКb8�)mX�-���xf��H�;�q�Mɉ����
�tu#B�*0���F�˘�>Ȳ	���GU��ߋ���C�0�B��d22�A�9��3�X�i�d�����,��v��P:�wnӢ�i��F�J�kR^.���-�2V
�`���F��+�	��k1�}���k2���oε6w ��ZH�2Ba�]�\i�>�؈d�-R2R�6kJ���(�&ƽ��
��Ղ�ڜ�V���E 4����.�l���F((��ٹs)[B�+�k�(�#��KQv{wt77&u�t�yϺ��b��z%�϶�@1h�rYY�Ȫ��ڜ�w�K����3*+cu�Z�t�b�(��T�ly����X��;ʂ�v�{o�+��Cu�z��r	�ڰ��M�#]�q��zL���`H*�)�z'?�p4ګ�Yk�f`sS|�p��9��n��j�~x:dWX����j�f�F����"[���L/p��M���7x��me���9u�,���$�C.�6=�\{���%6��H��2�ໄ�R�F���-���`�����G���h�v.���J����Wb�mj���7Zd�.挶]Gw��(�Va��j��թ��qJ��ƶ�BέP+j,����u�ֵR�z�v�Tf&F��DMQT�-DD9H$@QA����QJ��DS��DAAT�	JQLUB䵓���99E5B�U�!A�aIA��Q&A�!Ee�4U4ST�M��!K��UA��EP��@VBPd5@P%-D�4a	��R�P�EBR���f% Pљ�!����HU�.FY�&MVHPa!If%9���e��d�d�dd��3&�ѐ�49E R�B��b.HRd��4� �`�b9�RU�C�a%-9CIE�~��ߠ���T��t�e<�+���z���I���B�G0�|����P�!קs.g_\���N���|侺���� F�^���l����{��#�}� �z�g��<χс������{����vk}���^��7����sm�,�K�bE�f�jF��o��y��ṇw��O��QD��Ik�%蘵�Ɛ���I��H�k�a^���K���޳&܏ϡ�9٨I�*,����g�W�=6���zN�lR�{s����7	�ӹ�[o93��>ʟs5��Ud#��^�����^¼D�L�wl��/w>��k��؞ҕ#����傺y>s��uߒ�1g����KN����{�>�O{=����Մ�K��1�bâJ�=U��E��s���E�Ҧ��_xJy���(=u�jۺ���9ޱ�V<�U��]ٝ.-��p�F]�=��6���P��TՄ�`�Odi��۽��+���v7���	dy�S(���^���m7�ْ���� �����3��\��xb>�,T�j�q�mo���M";F�.9�I�#���&�w�Q72�$]fٷ����� ���!/�ܝK�u\�J�rs
����)�� Tx�@mͭ�Q�]Y��c*Nm��*��xx ���u�R��>�{&���@��c��0�{6��iP��3o#�^�(�@��5��<9;a�4�!\�c�gX9y^��Rj:�k���N�v�ֵ]��C��I�)��1�u���������f�w'෯}ZN{�7���;�bE�b�qS��ž�<�e^�V�8��]a��}=��ͅ�u�����塽͔+-3\����)��߹n�M�$���C�����Ş�-z��"{�U�]��BE�6/R*y��E�q���؟)�)*��YԩZ��`;̚����YB6m�Fz����L��h��ޠj�ݻnE�cM��X��5��;����=gzK(�y�oʏSϏz��rWFߟ��jM{�f����rX�hC�C�����ށ��5��2U�/��d������G��4{=ĩ����o����<�L�mz���������29�*8QOtAM�*b�P�ϵ*�ٗ]�`w����-Y���_F�E��F��a�^�t��=�T�mv@�J�u�jj�t˭�{���.��T`��Y���Lc��.�w�VI �-uKkQ1�kwvr��G����~���_Oܒ��:A�AW*z�b���N)�T�MԻ=�$���]\�n�z{r�>XD���f����md�D�{�c���$pT<N���v���wI�>��ڰ��@������8�v ��qw�Ė�}hwm��s�ܕ��7Oܦ���Vƒ�*�mP��9K�iy%�QK�k[�r���v�8���T�A�ЬgM����K��Q��=o�ʜØ�Ც�K��C����&�f�u㢹Y5\E�Bm�Ko�mj���鞞��S�h�$g�\v�A��0m�ĺr�]�hp�ll�
�aA��ySo-J�����wt*���0mAEm���U,oh3�f���m�Ŭ�n}{(e67����n+L��Ρ�]��5��u�Wm��ums��L,ۛri�˔'�񠾜��a=�3N��H�U�T=�}�\�<"�xn�ptNt�D,�I��^B��h
ï�P�/P��!\η��\0�� �\��4�ԬPQ:ښ�vE�5�C5���-� K����:��t	�V����kT�ęP��|z�Z�q�]p������{��̶������+���N�q͜�,�-�J"��,Y�����������ܛ�����d^�hu'Q������1�ڱH��f����bsɋn����}���y�,/��cFE봫�z7~)��ȟ:a1�H�y����_f���ey@uX������F;IC���\��q�	p��uz5tv=��ӻB�>��}Nz�.+:��z����R�n �m�5��]Z4�#�괺.RjB�]�Ay@lo��t�|�3�zG=
�q5�3�}fj|�
�]_��K��c�ŇI[Ds���oֽ��%�1zg��yo�l]}v�zXN��YV�ԊT�9��!�!loMHݻ2p���v��+o������bw�ͪ���Н�nlPT�GK��re!gE;�q9����+��b{�K0��{*�PQ���^Rï�sy&J��SA[1�+��L����Ķ�{:�Ӌ�q����`�hoj;�dI�¸;�yo�V����X�9q3	Vz�g#zQ}6�V�3_dcS����N	����P�Ú�T��Vpq_	H�6�[����Dj���t�(�d,�E��Ǽ=��̥�����c�t���q�NL�Yj�U�T_c����Ȳ�rg���4f�Ss����ozǝ:�_�������RX���[7B]�7.��1���^>��<��絃�àP�ׂo.���{Y��Â���M[ݶ1Z=���9��N'QA��i�e���n6ۛY+�ؼr�o5\{eS,O�9��[f��:��������t�z�]=������I2�93Q��1���/�ϩ�^�o�Z��S����}3��J͑uX���6@��PĎk��Q�y[vZ�٧e��0{��+�f#���v�G��lء�ԇO��<��I[�
:��;r�;��7����l�f��NP]JG	m��j�Nz�qX0;��3Vru�j�o1���K��,x>�g�$-<�9$�h�*S�ղ8)�2.�E\P+|�ܭ��r��{��MhO��Y��yId�]9�Z9c�K��S�F�Qk����.0�X!�DU�=:n=�6/U��h/�f�<��s���)�c8�͖��b��.�{�SK�խy�]j�Tr9�ԙ��+�:�>�������夋[���2��o��!f�Ӧ�,��aC�nJqF4hݚ
/�e��|��/g✊�j�]�y�����U�U"�n�3���wm8�/Dܾr�ջqȑ+���/j�j^�rۥ3Orw���
1��tW1�{L����b����O�o���g)X��}�������w�ӣ��.e��ir�M+���>p�ʗ0'�`�/�i��a����'����X�]�Ro������|�f�C��г���Ri���w%:�#2{�\�;�'�,g�K��2�<���`���t�?	nxk�WZ���{�紉ZR�9�M�*�� �ޮ1rw�����\����Z�N싵�.[�����L�$�S�y����T�I�]7���b�~ק
���sbrdS}^�B񱹩
���A��u�LY��U�5�������"�E��sF�}}ghWN�s$fr�˥,W�3[2[ղ_K����q��0ӷ;4�q�጑�ëie� �6+�����X+h�e���,7@�I�]���e���C����*�'(��H�rr��? ���<��\(�i��l�����ÆZҞ�q\���|1|�ؙM��]xt�n�Տ�֖'���<�J�7�R��w�6lyHo`>l�`�#7�˟b��n�w���&�C���M�sŮ;&�șE^L����1��W����b��M��J�KOz��;��Ǻ)ִs��Ƭ*�9�;WIj�W۴Cy��B8���|iw-Ε�ٶ�t�I��RS:٥����DN{X�{�h�<�ºQ�-h{"9^^�'E�pi��{8C�6ѝ��	�7��-�3�[f�uG���+�{pe\�����CQ��[�)�uz��j�R+ʔ&a�4�.��+j�P0'4#c[:�޺p�FZ�+����Iq�	۰�lW�gd&p)2�4-3��Í8����;�-='1ዘ�1ٴ�A�G��B�8X�,^��Y�Y%�[�!�V�(�ŋ�S̝0W'���tȐv�cZ��@@1�Fy�T��f�Qv�g(�y{�-�6oWkT�Ўt�TH̋K�n�:��B�k�f�V�.�D�A'�����*j���GH��k�ڶ��z:����I���-��Г-�%��ȇ9���3E*�=]Vcf���� {�ԓ������ۆ���%ϖ:w������8�:������^��Ml0����0��
�X���W��W����C���A�[3�U\`ך��&(]�by�oE�-���k9\D�3m��˵y�n�����S���ǅ9t��Rzɾ�Й�S���D܎�TP�Y)��.P�Z�鍊ݶ�_W��6��V���[`c��4�oy�^�F|>Kn��Zv/I�ϳ�ݑ��֌�\���ھz�&��L�A`k/��4���d�v�VֹSLn
L�bFE�j�P���+���z�4�8�'��O^2��^�6���Ҳ�͊�T�J���J�MC���ug.�`ڵs�mR���s8�P]��	)X�����6�5|���^a����pخ�\Wf[��_�t-!`lp���R+�P�\�U��հ�PΞXN�(N��Qm�u���Ki�gT�`ӽG5p�})�|`��!��ˁ�S(�̘n�C���y����_S���Z8]���Mc[��u�F=��q��oP̣�� c���Ա�����|:^�j����e��$$0��x�Y#6�J��]�ǔ�N���gz��?��ȳ��N���R�27�R��d9�4���8'��4�������S�Wt2�ui�G+�ج���N��qMq�>[+q��y�#z��q�[+:���(z���L�|��ګ�/:��ojz�f�*��@j��V��r��[
��qv���`-U/*�ozς�Yu�ڕ諅��-����V]��o"�e:Lzԏ=��}y`�]����{��龦��O ���=�K����q"̳d�\��2�=Z�R����\�e�+����˹�Oe���l�F�e�y��M�0����yh�|�J�1��i�v�qz�l-ݹ����a�&'�jX�c��k=�/E�Ӟ�Y�H~��e�f�jF�[�>���_N(&��æ��6H����{b�m���U�"�ɒX�=�˦�EU��X}�%H�#���DX�uĉ��w+Xx�Ԕ�w׷����#��a;�[I3�tV1љ�}x�WYr�p�y�'4�˅]��ϡ]ې��d8o��]���z��D�/AU������m�n����S�q�L��lڹ�Cf����륃�.9ի�F������%�T�^c�[Y0���o�lب�"��L��H�c�*�rGNk���Yѫ{g�u��^��[�4���[@���;�N�bY�4Z;�����/�_r�入��8���0���1 ���c7��D6L�<������������}��Hs�!��զ�]��$=!u�o��J�˅�f$��[ݳV�x��*ɬ�9N��qG~�+�C�}L�j���w�w�T��ΐ��[gL��@���V�YY8'{U�[�]c-&9K��K�U8:VHj�Jf|�V5�/�cuD޿K}.��Mn�a�q���;�gQae*,=�9����
KBq��= J�VZNz�\��B���{�{����!H�I�N;��4��W/�Bο�_�,�v���Շc����(l��5����V�e.���ig 2��l���׵�6��V\n�ؠp��@r�7��պ��9ڮ�
m�9�k;E\���z�c��зO>����9�Z�n�&��Jl�9wi���6jՙw	x�U��:q�}�b�[����a9~otP�EV�'�2�Ծ���͎S��ii��8I���P���quck`G������ �g[��-H2cuاkq�M�L�X2���a�L�l��m�Z�4���e���.%�5+`j�;B��h�vE\���A�-�ᆗPY�ؕ�YR݋����Z�no@�$Haʋa�z7 s�C]:�('J�a�u$7|��vW�K3U*�˔z<�q�j2���lv""1'�[7ztIWX�+��c6S�gu�
�sR҈p�����K9��n�)�Z+�Hn��M����]��T�P;p#A��v�Ul�&�)JjB�d*�U�Ct3+H�OLO@���6���sEo�}۠�GIU*G��Բ�K��*Ln��<}��������g�sVd�BԱW��|7�<z�$`�jQ�j��&]u�!��v]�
�r�7Ь���ص�ܗ�ݸ����4o�ǡ��#E�w��Nl��
��1�2v'ۜ^d��M%ohgc��A[���9�\�����"���� �X�)NĶ+-�wE��̵'9�K�Z=��3t�PO����D��h��L���I=����D�}R;�A��+4����oj�R�bi���@��r��X.�<���TI�������vR7̦s�H)X�Aܜa[\ZB���,�H���H(Kq������0Kjef�o�Ԧ�Y��`&���:�
�'rܣox�d}b�W@��<�EJy���t�PO� �]�s�ѵ�bD���f��2(lF�^�Σ-:JW.��,9���YR�U��]�Ʈ
���L0m:?E��S���W,�������څjɔT�vmz8���[���;!�1|ʌ���w:��:��'r�= �.[�UX��u�˩��n�F��U�d1�=��]��gXM�����H^Up^{y�"kd�C�o���ٱ�@���қ�	��
�xΩGHK{n�)�B��,Wi�94�Y5�tM�Y�a�U�M'����V�a�Dq�U5�ն���!hIM�����h��y�n�k��)f�[�XP����܎�vy<�2�5���
o�� �GN�]���!�Jp�����{uum2�@eY�l�R�p>�\3�ǘ�9���5���3��@�s!�K�e�G���+G)�R�%f�Oz(~��S_�j�����M�$�EwƲݞ�Uf٩nqf�����ݱ#c����W�A�}+s�Wq�z����XA��Rd!@d�P94*P�C�e���@4!��9&IK��*�e���T��H���Y"R�T�4.FK���!%�&@d� d�ҤY��"d�	�V@�B�@�.J
S@���dJ�b��P�	KY���S��(&@�Md�d�R�J�efAKHd�!��SDIBd�H�%��C�S���I��CBS@R����������߿y�U�0���]��D�4A9�5����9�.���}Cu�2̎�G�,��R�	��{r;�
u����3]��ƧwQ��n�f��,wii0q6��U�u�c�C�8+��D� }s[y{.���{��\����o��
�lP�*F'QM���<̩|�
�	�T�tfa]N�IKA~���mwzwf���z3e
��&m[����ݥ����Mf���m�>ק��H���Z�{�Z�Aɶx;�o���l���ܞ.k�hM��Iqs��M��4i�8�➊�����Bm�v��VS9ݜ��,�㵨�*�V#^��xo&��{�J��[��T#���RM�v�UT'x�o��j�L�O�
��ږ����;�����d����[#�Y�=X�W�*v����Ol* ���\)�;t�NZ�w����3EK�#�|{lP;��ծ���>ʾ�ɝG��t�H����p�{�ӕ/��S:��gG�h�e�~��-���H�Om���3N���������e#B�s���>4&�RY�����b�/��-� Qc[[��v��i���^\�"�3�r�
�H��W{E9�Xt�푭�AK\�3J�oxf��h�J��whkǯ�b���<�h��+��۾U�8��U˺�{�cG!K �qŶ�*�D�P��xpj�U�-� =�"����ɌuT�l�����n��;�a�ߔ���j�Ƨ/�+����I7+��N�]"�y$�C���eXv�B���B��":9�臏q�yr���g}|��i��u^ˍBv��دs{"�1�)���3�)`��7f�W��[��Q��b�˫�5��L6v��c �M�'�4h<��#��������U���u;t��!���l��<���ՠ��շ)u��-C`��`5�@p�gk"�ԺH\7C6X��V�T�c��1v��+�b;��a�����>�.�8��O��⮩^ܷ�<c�Fɫ	v�Vэvt�;^Mx��~����0�o��sґ��[e��Y��ebˤ�"��6��J�]��_\p�����4�y]�fW���7=�x�6-�/n���-b�lN^���X��N�vF�5�����4-��e�k#JF-\��s���+�|jMŽl�+}zvcu�^s��{�9���ޤј37P��ðSu�]���RDޥZ#
��»�����T2R�)��b�Fѓ�8h��+h'���]1}��`����!_���z'�"�j_J�FL}1����[ƭK�[�����VT�T%e���J�ZA}M<ިSP� _n9��f�t��(��^!�X4&5�[ƽjTB:��p�,ٿc�^���T����M*yG'+w�=x'U�x6�lL@�R,#��̎Q��E��r�ka�U���֣:U��ںjHa�U��.��©�P�Y��p3�
t�QUGLZ>�>����)��53[���兜��6 S�B�,;�qK�dֿK4��������[��z�~��b�b��"�;6n�]H�Qy�|n�EW5\��Qзa��C��w��?wp�& �z��Ӵ�Q�iz��r�uN��O+�`�S�ߕ�"A���W����''svn�"��S�e�Co�v���)�6[�Ц.da|g��x7[��
e���34d^hn�j�[xl!��8�P�M�4��8�>K��^_�y���H��n�n9�z+Ӟ�>�K�[֨�+*Z�M�)#�=l�	Gi�im����Ny���C)�e=׾��+�`2���R~�$�Հ�s�[q��D�7�y����Z��{�����=}��^���j�B��H�y�!�ʼ���kY-�*�{�
m��r��*��,�ZAF�t�-]�����C�N1���su�j�j9Բ5y��h�n-9�{�k��R�u�V���ʆ5�P��'<n#��7]��2k��fa�/ ����[Ͳ,�E�yo7�������w�Ǘ�x�����[����9J_�i3�0X�fz���G,˗�l���<\߮ ��٤��X=V��X����k�N��X�龄�=�0gK�V�r�w�Hؠ�cV�)ٟ
�_��:8�Xxqu�|�6��t,�]���Nv��*�z�r0��V��L�nI��2�1�P#dS�P�8oK8�f7��ZT��r�T�\�\^�Xq�n�����yř�g�1:���tb:)>�ZP�[�&�HL`��;:zv!m۠�5+����*��Z5n�F��J��<p\�Y�`���8�ܱn^1�4G)p����ޟ�B0f��>�J]=����վ5��qr�������o���sr���h��p!�3�|,o4F}����̉U�#�����j��swVOo��"(K�K�7���
����B�X�����uP<��S�L��x߽�R�s�v����*�s��h��ش�3�r�`ҫ����n�R%�ȉ����(�jR���B�kn�~m^���wg�NEI\"��Զa�8�m�ogj��J)��*W4#�����ғ7�q&oT������K��������ӤO�vjN�����Z$���4<>��ż�y]~�����/�50�8%�Њ�c��z��u���L�!^u�`5�T�N��Pƈ�vi�Hf�ʹ=]�W+}Z�XHP^Kt�fT)xW2����/l�őGK�&z#(
�zcg����Ւ4�WZ���{W���P�L	�t&"�b�����L�*��dS6#��	T�:%_�Q���y��"�}F��yW<����{	���0z-�ث
%�Ԋ�*�(�Ѝq����-�ֲ�4�)3�&E�P6�z�ۋrh��8Ya)���]QM�i�ݝnfDF�4bs9,��Ι�ĳ�K��­<���>��Khe��1��m����4��xļ7�P��0�tH���J���-_{������&�]F�mE�2;D����ռ���AG��"�R�;�<%��Q�n�`m�<�I���[*t�[8��;U+u�nG���w��y�v(�*�(��;ㅨJ/��.��K��6�a�Y�{lq.d�(�}�+	��Ql�Q��k�u!*J���-�\��a��J_7.!��Z�r���^�U��N��wyvً�s��8K����."�R(�o���ŧ35���r;�J�n�HR���aܽ|csSԝYd�UΎ�֪t�1��dfD�$Ĩ���B����5�4�-�N�1gL��#V:�D����_�����_tvu'�0�����D��HŔ]��Yu8�k;���@��#�N����J�Śח���(�{^��wģ~�*!X�Ȳ�R�>�.��/��W�9��h�{
{��k�����3�C�3���{��F��;�sj�G�(Wx��rH����ڮ�ܷx�V��Y~��P����
���#� 3�w��k|%-S���+�O���TP��X�-�+z4w1��"��H��[ufC��[�
+�D�v�TB.����2�	�aK�z�w�9v%���m�\�V\o�:�B�se����3B���*"%���dޞ�}�e��Aè�I���q��Cv�X�o�А$�^�{K��G���K�ŕ�l�6nwz��	�Ew���X�geZq����V�
�98&���0n�٥m��9ל�����f�#���薋�*!�|n�2�Y�a����ɗx%F��j!�n��T�{�I$5�|��&�J�LN�V�Z���F3�.�4�x/�^_����+�if�@�+����2RZxӣ�8��5��OlXb>3�
��]��͖����I�����U�L\�*�W�^����5�.��˞y�5�]�(NCm-h��Ur&�_���Ы.7�.�������ر�?(o�i2�*�?���m.�Տ|f���z1�HJ
���E���k{ݽ4��`�
(�R�$��[х�i�~�0��B�{�v�~gz_t�l�/^�և.=�H�ci�3d0p�
�[�T���z0.}h��H�.|�U�H�n�
㷹�f���4q�}�;��Zh׭��Bܰhf�$�̝)�P��+^�Q��ƨw\���1Ac�,흾i]��^�+�pS��38��ÝKC�r�*��."��YV��������ٖ�vkU쪝k��6�90þ*��$H�����r�q��D#X�X�6Yx�)��ީ�u�������⍇;[0��4�9F��AЭ���<��E��ɴ&�B�oec��׽j�u�j��7�k�H��U#4�Y<!N�I���chc�;Nr��(uidmD���x����J���H�)̇�](y�!����������zj܇�r\��fx�5
Y��e�Odneu��=�7��%�uc�K,sC��D]�i{̴:7oJ�=o��ժ���$]�f �`��LѺ%N�s{,�X�ùWׂ���Mt^�St����#�_��g�Q��z����Ӌ�1Jz���icU9���=Vv�,�RNE�6��3Q�o��pqe?����<")��[��"#�����9·���+"�-�Y�;����M�g.Qu��7�t��$(��	ץwS�|%>F���hS�0�7C�tG8�sn$]UT"er��L%�mo���`������?}I��Y�Tf��GJ́ᣜk�Y�
LVp
�Û���}��m[���;a{�^X53�~��7԰"�����v���Im��;|&�nnif<�s5�(�Y�o��ePF�2��ޠ\W�1Pk�8�E{��9Z�:w��V��tT�Y����;���s9GM�۶pdKC#Hb�o/�OUíZ!����t6���ׯ��͚�q��ﮛ��V���T�k6Yb�p�M%8]�ucq�-Ss�n��dݺ�{6����*��T��=Y�Z'��h�
�U?y�[]AҼ|F{���"���[���y�δ�r}g���1�S�p����5�ׄ�e�P#i���������݅x�kT��t��Mk����H�m%h�Zj�G�GtM��"���#ٛm֋lu������ffB�aܾ���f���8�Wi�sw�H$`NJ��oL�ޚ<)޶�b��������ȼ�7�m٣���xN&�:d���SH1;��{�mXv��`��_L���w�@T��M��}�{0���0�
�5��.��_��Kt�|��9�WG�"�e_zB,ȗ�l���*�i�50\#�:�ס�8$Ĳ1ְ��CwIK��Z�d���M���-
�;�d2���!Ї�qÈdCG�t�-=H����ryu,V���a�/ђ�E��uHؘ��_�z�؄Y{9��|��,��/d�vk��ƚ/��%0�������%���
Y�
��$(�F�]�o�hV;i����۪�v}e��k�Yu�meq�e�D�"CY1�v+'O-��QJ�'���6PDC�uzؽy��,��2�,r��	C9Ι
�,����N�L�z��#�s�x�e��}:�U�v�D=J�E��g���o(O��`E��	�se�Ơw� St|g u�G�آ[�M>��O��2y�X����H�3c�;�bJ�Un�z����/8�}g�V3��8�I7ӥ't�T)hF�z��Ze�r��編�b/���"��^�_��ؘ���%*sx��J�z	��������J���l9�<ee�:�b����E���7BeEޭ��N8��=�r*�n7/��!�)�[�+9���n�T�Z����+�u���1�h%A����8��ʾ��p�
}DpϹ쬮�pEqX�#�0^u����q*�^,�z������5�;�u�"�vDv	��U��=�
�%�ū{�_��y�wyrW�x�3��C8�ϒ�����P�Yk��ݵNR:��{��)ރ0\��<d-�f��ڞe�.��A������l���>�.����S[h�.�[خ�3c�~�./���G�q��j���{���W�s���y0��G��w���.7��o+���(�	�F�QC��F�$��W�o��;T{B��
�VBJSvL�n�*�4�(ձ<h[�GVJF+!�pQu/2R��hCp�S�ccG^b�N'������zus�2�`���z�R6%ʈV'hYF��T;j�<VCܔ�]�v2TZ�#;����J;/���&�8W�p~���7BR���o��yN>��AN�u��|��������{چ�%�;�܋8���Vzx�^���VФ|�[�V���S���q�a�^^>���M�3�{L��d�����\7=�R��x�(p_N�!�`.�E�R�G.��Tb���Q���X�}l�CΜ�N�6!�\�n�n1c�4K��
FU�8J�{f�u|��>��*��{wŞ*�b�j�Q���j�8�ŋ��^kG�0��\���]-���N@���P�d���^Tc0��e��*%��(]A`gN���S����q��D8�-���r�C�ƌ�O������ �r�Z7 b�tf�wV���5��X&��E&�Q����4�+�f��i��-�`m�7�r�K�h\�CK'.�+<sQ����Bod���N8�4��P���LҤ�P��`ʾe�{p��;���kl��aWj�ʺ]�qM�-.\�y;����-4Kr��)�GOe�:�Τ���p���S�R\�L��sw�P�O�S��Ѣ�ђ+�MnW�A�fofIgm���׋.� cM�*�z�,湳TgKJ���LU�Yj�KsS�ޫ��ή\���`DOtެp�]�r�5�"Ŋ�:9���\�^�$�1d�w�Y}��<�<|�i�>:�%���cj��݅�B�*��y�RG���\;/��^�Z�1n��"���%t�3,��{&{��޺�Y�
�؁�CB�� sZ͹V��0�M�V�Y�-\(��`������J�-\p㠠!���干��d�B�q��[wR����-Ԃ�e����`�;��4�:o2�	t�̺�i`�aa�{��!���Ɛ��/u&&dn�X{�u�f̶m��'-t��)�E�p�w#wX�	�u88!�'��ph���)���|���ɀu��W��(Nu"�v�q�l>Zlp �ձp��JxU�Hތ'`����W�m�m�ն�6;xN���a��ZdS�Y4���ʇ��շ(�sy ����Mi䬴��tV��j	c������<jt5��阢1��e���\w�*��:t�GX.v� ��c&�K���Y�F�ц�4v�l0�/���sF�B��o������R9��Sf0:��XF�*��䬽e�ى���R��K?��:��0����0쩃�r_Y�BC2{5��F�;��'x�`�i�v���f�[U.��`��я8��; �ֹ��b�v�i�	=sz�[���	�UfF{P�ML�ǉq��svN���4�bQp�@�BEve ����R�oZ�ʝ��K�}ێ�4G��Y�t��^튖_���9�x撻��X\�"�;Y�x�8�ռ;�v�E>#�rf>Tho5��t�oXI���B�&}�\I�,�OJ���5h=�>[�<eLb�ow��[cFRU�J��vnS��ƧnD�Vp���Q��8yom%�]Y���@��q���� ���7UN�4gv����d��岯]g.�1f��s��crT�K� zf��.����Մ�:�;���d����I I�����vT���֥��5���}�MDmm�\�Y��DD��w%-�7!M/��vqw K�,Ep�)���pև"�6��N�ZK3{�]���3��L!��r22F�����rB*rD(�*��
��2Z2S r����h31L�)hhiL�R�r *�V���"��2L��e�hL����,̒���2R�V�ZL�0��p�r �Ƞ)(2r�
J��p�����'#'$)�02%r�ʌ��J
�hC'&3�� 
��#&��&�F��1�rk,� ��h�$2�R3��%rC&%��l�Z2� r�ʬ�!l�2L�Ƞ�20�� r)h) � ���>�#v7,�i]�N�]�K&�R�Z�gfQ�޳9�[-�]B]�Ǡ+������do�m)�kg�MoN���꩸��o��e��e��D�Y]V,���q3�~v)��r���/au:?##��rim<�����:�^��&�KC���p�>��G�$�QN�1a�q#Tl*��z;y�3thW�r'��IyA.z����-�S�E<s�q�PޒXn
���l��y��IB�$�
�$�Q0��vRk���6�~A��4d147ޥh��zz��cӷصF��ͨ.�S��FDo��f��&'Ö\�-��j�6(f:cVFe���u�O3T�[�xYʭ�P��N^��I{ӛS��1Ql�\��@�Ž��0x{c��$.>n�J��{�Λ�B�xf�`�ҙ���6�<C���\
�3.�W[��3�$�9�ݍ
ل'��Zh��4-�6'r4�b��"�O;a�W�+mq���������֠��lJ���8�B����q�!W�Yq�E�j��}K��]rz������=-B����y�N�R�����񞣣'.'����D6N��<0�[8���z�V�䶳�����^���t�3�>���;W?X��Ye;���cS9u1��9���\����w�"-I/9�jI^���z΄�F/2Xq�f��w�rr/p4��p�׉r�M����a:�G��:��CP�������}�k�-�ʩv�/\�Y/�Xӳ�;:f�IG�Q�P�"��8��ГD��y1/(���\��7�]��{�y�V�Þ2�T�����`�2!N�5矶ʗK9���{�պb>��k]{c�׫p�	���H`L�[6%�<mF?K&��p��%��{�bHՓ�+g�`�^�3��֣�+_VCb�L���e��s5aA��wweך�Q9�L�u�ʕ�Y�/,�>�'�X�LZ7O9�'y�j�Ϻ�eK�̤����ڝD��������2���*�_�OI�O���=
b���*�m�r>�E�[YǊ�������Jd�
p��8��I�:�eI(O|+B�#��叐���#o���zӹ�'{\X�z��+����W>ܰy*S�_����AE2�:�����̈:5 �\��L�K����A��#�HJ�b0fk΁ɫĺ�R�nVz B���2z#��a�Y��ɬ���J�-�3m�[�G�׭a�����wP¯ڝX�_DXQgTm��V%?V!����5;��C�b
&�OPv�U�Q����Af�3:�d+��ͼ���:B.G��W}M���Sцn"�%��,:�{���z�b.�����fuC���9O��*:��X�J}�vL�r�Q��2*�/���� �x\!j���wp0��u�R(<��o�<���u����LlD�vR��~FP5���#$����V62)L�y�Oi���\��][�Í;u!(�yY��K����V���=������f�P�S���0e��'=������Νk�d"���R�kNےk W�j�0zc
lӦ6��ݺ�(�b���U��Έ��㉏]"���]��{���h�й�=V���v����y5n�x&���V�j�("�l���N##o���5�|���=�W��ѫwE�.D Au؜���՝+�I�.$����5��_N.QA�9E��*P2�X�B�>~���M���毻�{`�*=@qѦ�.�������5���/!/sۃOy^\M�Fm�Zgd�k������a]�ӳ<��
�����d�>(r�G�����p?��[��Z�N�rEzP0K̠�C� ,*4��]YTq��5�}1�̅Ѽ���c}��C�ٽU�lV�E��W�a�4p��WH�z�[����,$u�0W�L_.�g��/-^rVi����%n�Zo�N:ƺ)�{\ES��e���{1�2�Z"7��մ�
���Z����k{�R��V����|$l�X4��۱�v^�V�L�{aUӋ5�3��ȹ�d������gL5$̅U�o����,S��K	ꢕ�n�	�q��H��:�4���h60t�PT�HUQP���YE���&#b�A\��j�q.5���Z��0rp�Q#ٱ�KeN�1:f+ʃ0[�=�����kc��!	��q�R��e��S/ �&X���PLH�N�L-�����\�έ�k;v�$z&!�B ��j
��ҩe�3��U��]^&:����%P\�X�u[*���9�J],���<�ۜ�$Ā�ɥ �͸�Q�JNur��^&:�h�ed�]Y��:��z��$yFi�j�K����� �����z{�%�6�k�m�e�C�;���Ǣ�+W�����5��eE�+�.��7�Va�V�RS�8ub�����!M��;v=�{'I�`�P0�.#�d�b��
)]�F��;��q�"M�:r��]~����$���w5=J��T?N�&Q�V��[�GW����(�s`���+3��%7����SkK��z����Cl*�����jy���ұT��}~�K��ꙅf���th��U���d9�t����9�M�O:�"��1rc7V38��ABV�34�=�AK�(�K��m��e������b��Di�I����TP䍙ӛd��C�9y2�+3&M��<jݡo��,�+� k)V�j�Ϫ��P���Q��Q�C�,փQ��B���p>/����L��-
���Ӎ"���݌aI1�y[�g<��#҆�	�wι�|+hR�� ,��5..N����R���򕝝X�\�C;w���9q�۫2cq��(�T@�C����@ڣ�>"v�լ���0�i��i��y����a�s���ʋc�4-�#4��o�M������L�w�A�U�U�
��O�v�q��i8�}ϊtg.��mx���'�W���}9���Cd�ڹW�v��A�yj,X�
���x�h/��b�˲�w��./��XQG$�s�%�0߄�ԦZZ/|���q��~�P�#Ma�s=�]N
+	�#��<I�bc"��1-i��5��zc�U�F3�./ο,�ɒ��d��s!�2X��UT�$�ё6ha���3��r�Ϻ��y��ǅ�� "�=�:��-�P�3fX;�p��8^�us�f��t=�|�0߁ �'9)o�\�Q��(Y��O�]�Kn������9xϪn�Ccs��+��k�(�Ms�I����-�#�mЁ���_2Ϊ��Ӱ�:q@w���KT����L�e�Υ��$SPu��i�ɽ�򓳓<zqͭʚ�wsJ/TWZ�P�P��� �*D�nv���\*GN	bD�^�@�♅P-��i�LLJ�̸]�߷lOR���V{(�����u#�5�4�ڭ4kք�nX5�,�@diHŀ�Qv%s�Շ62��:�z띗��ZM�\;��![�ƥC�+��eQ�e��������Z|��C."}}"ʑ�qGI�Q�zn�|��9�>?i��T[�vaPr;}(��^!#(4s���-r�x�k�a�g�{z9Ugj�r����S���xzx�yI(�zUG@�l�)b�t�����Z��C���'*�#��:�c�q>�!^m[��i�F9�@,׋�%e)����[�Mk�����.ŠQ8<��D���;�5����	���H�2:�ϽB���@��w= so77���`^$���
a�\�|=)����g�
vB�z]�K�|&s���j���ȟ�9S}�oň$��f��)\	j.��K�C�i�V:�Xo9�/'���ة��ت{R�,qX#��T�4�5]�s�l��L\ W��upv�����^bS���y��WtWZ�M�;q��H,�%+��&���L�Q&�A��abyh�# �p���a�ޡ�2��Xz�r�>\�Y0=�f�ZT�hjZw.�.���Fc��e�΀OZ�iV�k���0�ƱP.����L�׎r3t�O�k���[,���R�8��n0�AT�4ݚ�W�o��-8�������W~���a,��c�2Z��AR�E������a�dHS�%��ZR����<�%p��ޜS֣�i_'�z��a�</��*�R#>��'��;�@��t��XO-z�{���E+�K��=n��|}w��ld1��8���V&���AѺ$��)5T��,���Y�u��`�.AG6-窴��Zo�R�͆X�l�d�\�x.���C��>8�ǻb��շ�
�v��xL@���~D����"�ѕ(�E�T2rv�G����Z�ش�:�"ym2�ϩd#�����Zv�y ���cu��_èV*W���y]��-�ͬJ�t9��zYǏ-r�H�m%h�Zj_E"��J�4'��@�[%T�1}��Y}�Β6}(@E�ّ�1R��b�q��"��*f�wb�w+F�Ip�Dj����E^�zq��Ap��{Ȇƥq��C6��B*�W�j�3蔠a��m��5������BK�I�]�E�E�0�M���g,V/��%���\��$sy��]�u!�ѡZ�W;7]��X�"{���C�b�J�%F�]���o/����Ύ���5H*sh�ywL��`0�ף(�lr�O`Y�r]��v�;��҄������}��#��ΗPt|�Y�9�o�ROq��^�`�����"����|��І%�iW,�B�����k}ae�'���r�X�'Y�����\5J�顏�ꅛ�X�q���������d<"V�l@�J�ȋ���o���Qڤ�q������߯&]�:���\2����Ex)F&�[��b��$S3�6�K��uTm{�㝎ѹ𨶃�X�5A,�cL��g�꼛���_I���͖xG=��
в}���>W��ҥ�^�1�ʕ��2�xD�ʢG��Xd��6bt�|n�fS�gc)-1[�>RI��#(Є&�v u�W�Y�5�]Rʆn��`g*��t1!O=�b���O&�9�{3�����׊&l�C�_j
����K.�N6�yߍ׊�9R����攫��v�c����H}}�
2�nN���"�ז�(:�}���9A]��UHL�{��+��{V��8�/ݓ�ź^�u�E�<;�hj�a����u�sQ
��@���.�|��@{mdp�J�ZE{�:`2<7<'�˗ucZ5�[p�qYš�f����Ɛ�o���)�b�<���YPhQ��,(jgcH���Nx$�w��F�y�IX��Ry��j��b�����r�.��]k�}!��k���k,y��;�?mSQ��@��eEv���6���3ns"�*Gls���֔��W뽓�����Y�W��se�8�@�ђ��#\(�w���;ㅨJ/��y���^��/ٽ�����)jb�RZ8OQ�N	�)Qv烄]z^,dS�䰭�	�})J���]tڍ���GPUO4�ɋ���}�5���U�����0�/x߸$�O�w�^�;hr�V�\}�<�+�LR��d�
��u1j�qJm�
��mԾ3��ep���{�D?s��Y�� ���P�L+���dP}��#��tň�Q��an�Vm��؞m��F�F�8�
s�)�����E=t�\SsFG9��Q� �*j��WjDQ�I���,z�ۛ�ƽge���Ne'a�j4���`	��t����glgZ��z�^����Ǔ�0�N��G���ӗ�����1��˕���b�����=PS�g^�;�4�.�U�� ���%P��%��K���X�geZ�u�������{m�Z�E���Y)i�[���+/s��#jV]`9��;l���EϜk#���*t$�@�!\�r՜m!F2��9���e]���К;d��d�%�௢Zu�o�jZ7�S��ܞ��u��Y�1]l�ӎad%���
�8o���I�葀׵:'h�.!I�e�6���r�*+�q�㜧����V�+�/��(Fg
��[1đ����#FvSq��W#��oь��Q]!t�9/��������s�а�����]D��lEbE��tL�YPp�Ck����)���X�z9'�1����g�C�!x�
���`�r�cTg*���4�P�J� %?�EB
�Ƽ�ܓ�Fwu�~��G�_o�{T��3d k�S6���Q���oF�՛!��R��s��|����c�4��łu���S�h3��2�� ��o�{k�nz_��̈�M��ML��;uLB�ze7���f����@�do��u-r�=1xx�����z��\���[x$�.������\�
��vb��C�J40�
b���3���8��Q�MyMy�o[/I�ժ���S���h]֋8��ꇠ����v�=P�
��d�rچ�ZLv��b�Pw�t���qōrΦ���׊49t���T���Y�4�.^]T��̝׸��k��C��3�#C+�1���VgH��sw�fLeZ���E��*QW(����.L���gt|ލ��d�>{��+�Do�0���Y��b8Üj!�O��}�T�W5���P�a��٤$�IM��ua}I�\6ڼl.9�*�B�]���ȓ��0[$;=F�n�2���E\|��Ō��.&�Y(*;�ˠ�.���U��K	]��R2�)W�;j�#n��.�Z��wԻh�G
���4(�vy�`�*�[բ���R�G)�QH��w����1���]�<>�R#�橇�A���r�/�rv��]]K-����D:w
�(ʠ����k���i�g3rด��\��ۥ]���vb����)Aʲ�F��ާ�����w�@ƈ^koZ�pPc���d[��M��f�\�;<�P����v;,ҭ�=�K�κR�]>��Z�L���
7V�J�-��^�ƞ�bQ�u�������Uy\�C��du�ʹ��}R��Y��ݶ9��d�Pʐ�w>6��1:���t��XNӂ��6⇞7Y�ܘ�ݗ7j{��{vuMBL	��e�ヷp��XLu�0��:X�˵.N�D	^<Wtނ��ж�P���%��E�*).�:�q`x�P�݆�@N"��{��sY��:�$�L�Ăj�b�3&7�p�MMJ�[˻@]8�I�|��:s�@�\�N)�1�H�T�[���M#�P��H���l���z,pѯ���imH��Z��mk��,?\��K��ܔ�e#e[��gHt����XyŴ� _l�C���/���E��S�9�ܻ�0M7�hXt��)���	6�!�i���u�[�}����P�ں]��ҍp:F�]Xu%�6��q�,S��Y��Xt�VK �����P+ �h[燲���Q<V�^݌H�p}*��](�˽Q�a:�J�ME%v/)z¹i�eZ����#�|�o���)u�ت٨����n���<y�N�gcx�E�oÎ5�ᢒ�F�ݘGJ���X��-� v1MYzH=V�y��/�.�t��:�M��k��x*��iٽ���׈�u����IEodT$�)aA����;+��Q��_,�99�v֔�ը(s[��&��vX}����t[�u<�s��8ig@���5�Ҭ��.���8M؎��h��'����S A	;[`<�c��Ԝmb���z�v`A��V�Z�y��.�)����}�ԙvȢ^��M��$�\)(l��S�Er;sJ���忖$�Ϋh#"�N��M;��2���ZH�E��ԢB�h�]�C��P�Wi��e��Xy�!j��������"�Jv]s#���U�}YZ�'���a�5��c�P��#�vY	�"��ܲ���+k"���b� ��.e���� !�{x@�-̳z��� (�6�_ "Ʌgj�=`��㓳dnՙ����tq����-bfsg����{��ŕl�9+�>+�l�B�m֋
������~�ϰuI�L���D�Yfb1P4吕�@eB�PD���fa�dTNHd��IB�+E����IE+��@Rd-EH@(PP!D�FY9�PV�M�FI��19fE6`�Q�EJ9��9f8@��@Y�E�RFNAAF@P9��91d	K��d�%CSY)B�M!�f�CEIM.F�E�AIBP�C�P�C��46F4d�QEAB��f fafH�IBd�4��d�@�u��}uֽ��~�׹����53`y:
U�>��f|�}���o��������YT���C�M*R�����ltkv����FD&)G�B�$׌:�s��,���لC�p�H��6}-m�,8�#S�t5 �+-0���wO/���3��G"�.�:�?�3��v�_���*�T\�e�:Q���c96����.�hDs�)�����^6�ڻ��S�p���g*¬�[�uن'�f�T�`��(!O����v'�-&Sz���<f�ik�i�"��S�c/mv���G�	G���.�O7I��x'�'^�P���-8�����*�3�%{����Q���@ڹ�M�:���!��9j�#<Ι�t�Ifj*�o%){f�J���&��fD������r�3��ѽ@��50E��%�'�m���aoz3YN/H��v
�Rr���7����)�7�4��P�u�`{�����[�Rڅ�no�s} ���b�oB��U҈����5�V�5��ZleJ�e�,�,��f1��EXK�υ�-{i���b�E�m���3>�	h�\�TG�&�~��*��Ӌ���4���*jf�H�{�={���
��|Y.Q���˻#��.�CtZݖo1�	I�ҒG�����աܵ����(�A`�.�.+�`ћ�����dYGL��]>��8��/�g7�e'\�f����xs� 7�������K��龦�����=�%��4�נ���b�6=����NV@U�౱*�:ϬW�Wpjj�X�OX"�s���#F�g<�]˭#M���s��mE�fQ��i)��F���;�{�3��t|�
OԫC)�C(��)G �"�=�l�������6�xL�~��Emޱ����Ū�Ѕ<pX����H�q����NUt�0�N8"^]]TXq�c�+S�+q�;A�R��ͺ��h����7��4v5��p���I�)�f>�nȠ�_�����ٷ�>�P�9�$�HT;M kЧ�D_�K63��l����*/��)u����ZS�؅q��[�zo�F�E��Ȑ��j��%udE�S���٫9�)�)=읓R��0�ݩ�/۞:��F�~v�M	�Wr)Q��tj�x��ed���^�T�����눴vi��`�3{�E�O!���3�a�z�wqo�9E�{�#5>����ܼ�-'�5+Q��ՃN�H�؂'�&(;h0aP��;NY9S4�l�r쩽��E�gG�ajq"�H��x�]�(�NQ�EL���ˆ�o]ؑvR˭r:�Ε�D��8D�EZ��m��)"g��r�V��j
�A��$�X��`tC���p��-�6�[��=�N���V�1͙�+�^ݕ��o�8(7h��;j=�����ϩ;��k�-f�1��m+��mO�2����^U�2�Ϡ_�h�-�~^}������^(��#HT�Zh�hJ��T'���Yi��;S��p���P�ݭ[����]Q�VDw9����C�h^)�3�������j����4�VsJ���'�2�h�/���]T�%ꡇO-����F5�7a���I6�^�K��e%+�[0�26�� E�5�(��w���8�cZ���4[wn�;}�(Κ������a`�Pߪ���M�Z>�Zꯟ�:�Gz��5=���Z���阝���LvȮg�+��*�GLͨ�=4p\�m����씌P�N1�Qc/J*d���4��X�f�΁7/��қ��DW�C�P�؅ld�j�F��D*�QQ�����Z�*�㻨�&���Ҹ�\��z���TOa�j��7���q7�s�dًs�rp�T�%�҃�H���ܙ�m�jaX=<f��PU�H�l�D��~o�PB�\њ[拏_0_k�8�8�m�:D:>���o�'v��CB e���y{ی'45���n[V�7��6X�Z��;\j����xP����x���.1�s:%݁)5��7s��yW�q�2���OD/0��h7Ƒˌnhȯ9�9 ����ƚ(N;y�����w;GV�^$�O�]������9љI�F��\m���,uf�a�o)s�jӥe��fb�XK
 j�"V2�1u^��{}��wю%�Йb��ߞ�|����q�a����鍊�Y�!Ѫf��;���F�l����ӿ�E�5z�qBk�aV}0�9'$�8s�6O�GVkY��{(��}J��
����}�_�R�<._�.m��D+j�<�yQbH�.�Ber��֫'���A�(���f���+��!q��g�U�f�9FUeM8MbE��5�1�*L�a.�ݺիV�ޓ��!ywS�bx�`�^4��^�4��p�B8]�o"N�̀�a�o3��w"t�L�,��v�I�!EN��j��~��,_�}q�3u�1��x�}J��\=	�o��s��=��p�Z���y�
��k	����ÝKMr���,�C#JF6��#��fD���V�w�H��C+���Y��xԥ�fVl�*b�U����Wf�>��U�R@��6�qr��o�wX���g�v�{���A�>EQ�ة�Gf���CH-�� �Û���l�oe�nV*]ʭ�g旪g��|-:�Ē
�r��=|K�ל���B;_��H�!�\���n5>�9���N�G�6�0�R�|a=�͝��K|T�zgt�z���Eו֕s�l� �J���aP�ha�ŃBc\P�µ�ˬ���vd�A����Bv�"�7�J��躥�6��z-z���j/�����!�_j�1j�uSw\��K����(��*�!�6�3��#���(p���U##*�{��n��;����K ,�xѤ�����GLa�PS[8Q9�͈�?e0��T��ѩ]���d�G:)?�2kU�L�b:"q��(� �+T�z����_z߅Ծv�G�����ke==к�?c�i\����/�+�' Qm/-��Du'��]�(]0���d�i�]���Dx�1s����l�dH4K3R��V<�zL��>*��a�F^ѳٸb�9��Ll[��f�G8��T�iģ��,�%L9��2��7�,�x��wq�'�I��kJJ�����!q�i�%��!�� �"/��3C"@$���ƈ2b"=�v��j�"�#ԖGC��j�Z[F�=����fs�@;�:��%�����&��y�qIn�ū��-<���.�<�k^|Xi�}ݝΝv�Hڎ�#���\�E2N���从=�@��ɝ�0̗l>��A�XJ$�]�8��Rv�<%n�� �����E��lJ�3��>�&8�F�4��#�JFՉ�j'/��;6�,7�-��L\h)9Z^zf�P�t�S�lnK�Ő��V�kbxͥ v*/�7����=Q��g,[2�Ԉ��L���<�V�ޜ��E��mfWWo�v�$�r��)�i��}���8�ޙX��GP
8���FLH�뎭�N엻�y�ivuFh/vx�E��EŻ�"��y���(>u����i�����!� ]�S5&o��Wℎ3�����fC�n��%)�|i��gC�f�z����z}����A�����;"�����t��߫$�4�>�8�)��TF���Y�/����=�\��I0��kiU#Le�P���<p_�x���8��!DJP)EtZ�!��Q�T�n\��uOi���J�(jr������C |�Y�Ap����������Թ�\���xQ�`sۃA�+ˀ˘�GK���!PZk��
x�E�R��R�{��1�[�ˣf�\�ө6�mj6��;(�wYt�!el�e̵QL�L�b��IV�7A���i1�8黻���Y�2Ω�$F�}�Ӳ�9�/罹+�5��+�.Y���K�sz��@�N�،�zݎD��Y]������inZ���5����aWjfns��:�V�e�m
s
�b,k5��5n_9�k�W[�;D���8+��J��U�^,�n�X4�A��Tp��]Y�W�uj�Z缩%��xϭ�l3��+}ʸ���-�4pNp�Ю�����c��3�o{��~�|�{�@k=T՛N�� ���<o�o�i�U��8�t
�1ֻCs]�E�_Vv>g2Vg�ݞތ,X�6=B��Β�u��V�¼��\*�H��D�����&������*I~��O�:�y�;�~�\U�����p�f[\v֋����I�"�*ވ�oe��;��$eX����F�&#}�L��8:L��ɑy��^�6�v�R�����2ک�<�<X��֪�"�u�`X畻s�䘗�nHD��8�Ti&�0�ʖ�u��}��;b����}�T�<�C|�CU;���0鶟_l^��A���79w�}�=8,�\����ё��":��0E�7�(�UV]B:�֫��+v+�B�2������v�N�]�_�5g8����MP�(q����L�x�R��w:�����n�����/H^U�r��^k�t�VZ��T[�;�DRv�һ�_9�e׼����u��Oc��\Ieb��O-��
��#/y� 5lq�T�'8�±uJ�kii�*F$H���H�e�'k�K^;[���Z--�L�M��#��)��ڑy]Ib3t��n8��w�f�����A�t:�T+�ϗ&.�%���o������F�B�CZykT⪵�O1O\5��ދ)��{�T`�*b�e�K5�ׄB��nzQ\yX^�ڂ�͞�շ���88!^]��]��	�����ڹ��qdh#C���9{�cy��$�z�8����nU������l.�{|K�.dh��n�ȷ!�D5bJ0�K�i&�v�c�d,kO��0J.��k�׶��sә��#B������vŬV�s�S�CM�j���,��
FS��t�QWFϗSB�z�g��>��'�r���|�8�s�p��#�����h��ܡ+y{K��� ��~��&D�J�.:���J6��^��rj�V1����	��9�7���
�rL$���)L�W�x%��+�>�p�+��j�����݆l�7z�u�]x8�$��'$�Q֚�Rk��˽=�/6�H���!�d�+r��
3.Ϫ'�|̆���6����͕jN�#k�qG1f����2�AE�|(
��,d����V�ܼ�8�T0��p��%�a�}���
����#���GN�V]ܛ»H�;�j:-�r�������YyoN�Z�x��d�㩦�xϨ`C���ds���(X�d��Ԫ~@6�sךղjs�g�������+:�j�%���)�Q�1���UEf� o#1b��K����V�cO��)��n5��l��w�؀0�E��1�;&����iQ�H�]W�[��iX��l�y��*7xV�RR똲�]�X�euֺ���ϝ���	{�r���,��5V�F�+캢����K��.t���x;5эHݹ�rF��e�8��z�u:��Z�t�)��'��D�r�p����|nW�Fx���XR�+��,���R:�j�m[nO�󋇆!+�,��K��#F�qN_Z,�s�� =<f���l� m\����
��y��#D�(ӳ�sC�OD#�T��X��)�U�p�L�trf�>(�%���{�I�7h@(�B8�:I'�Ȏ0oP�m�=R�����2ml�����g,��\�� �<�K5�z"���2��L<,c>Ga��զ��'�}**�2�&�]:�/���[V����"�|k+V!��lj�����e����.�q�jv:�af�1��n�@�ꊳ2VpY���.^
�)-}Wp�́�vO�,�zlCuEzP�m�TYuή�n�$CY�'T�V��/��",�u<29��r�"�W�[s�e[��Au?@��[K��[[�b��~��gC�`���>2E|��:ۋ=QB��L\�7�[���"AS����B�eG�����г�܏��fW,��2ƺF��8��P�q�)U0]��:lFQfTf�����ø�2�G���-�o{n��É�����E��A��Ṯ��"
��-~&����k��'d�N���a�$�K�<%��m��rS��:�sƦ[u�0�(oH.8jb����4��mQ�����O1.Pn!��p�o;&O!�Rn��J�^�>����'ʺf�/'�"N%�:�x�t��sv$[����p�E�+˅A��=�N��8na�^Z�çy�>��N�(tY�N����WMz}��%�q_����Ձ��E���3X�y'���?	�q7�[����TE{:Yqj���+eoJ��oUv�NO��viO��s���w~�}Ғ���L2�4���T(�ޖq��Z�ZF�%h���MH�ݞ1;�Zv���تyĢ8��^n��xKe��.T]q�Yה-`�MI���n��	�XH��{\N-��ǁ�+���l�+����%[r�'���9A.5yCV(����*..	�KN�Q�����r���+�)Sz��<w"��-�gc9d�J�꼭��󫦑��C4��u�����!y]� S2[� �f��ښ�I�6S��4u�L����qT�3BN#����4�K[=�hs�ɇ���s�<ket�
�(�m�gJl�bкJ��:���.��T�M+&�R��M�yʉ�w/�v�H�ƫh��$�G#���Ǚk�ED�t������<*�'f�Zo X�v���5Z�*��o�#z��du�)�|
��'M�;�����y�X��3��#�޾�`�bg$�O�c�)F���f9G2�d���F��J�f�C@یi�K(bg\\ {w%�Χ��Y/3z�r�:ӫ�O�=
�v�|��E�Tʻ��9�.Z��7}J�<ޥ���a���42-����k��`����jĳ�pK&���k��c�,!��<�4��7���d�/i��Vt�1��pr-��om�Wr��R9��|�+q�(Hݷx�9�m��A˸�)dp\��F�ۃ�#��b����eP~V��w�B�ޡ�e��Y��7�V���:�A7.��ƱNX�V\�ua��N���;&����������F�Rh+7��t���L	ِ�k�ض���N�	�����9���R�2����)�vMЭ�X=G.����T�&(����S�-��(ffu��T��n�yT\��1lj�Y]!�j�V�P1N�!�]nF�vp��m0�M�ч�=ܹ#5�O�ӄ��N�f��8���Br�B@��*"�v�0u:Fl
ڍ�S�f;�f�uK�,��K3stH�t�u�����@�B/��U;��Q
Ѝ�.�/��K�%z�������ƀjQP�(z�LK�«�gle���\PY}�u��F��F�؄Da�
�j�'w��^l}.��W1���؍�;�����2)x��~�F�j��ǰ��*S�h�|+I7M)V ��wМԳL#.Fj���ɄҎ �E�bZ�[Y�*��-a�S~<�ə����CbIr�V�;��C�q��1@�#��5���,W8���mfZnE���FD�"v�Q���L��C6f�dX$KPl���&��w+������k�%E�%}�'$]�Ԫ��������#�_1�R;�sI˦��S$,}�����睷���hOs�����LZX�Y�&s�k@"��4�v��7-��[�r��*��BQ]��GJ%U��)�Hkq:.tM���7(��K��]�Ɲ�FaY&5�'�I�d���e�l��e��YXe��f�p� ��ݹ,�L}@}@V�2)(ij!�ɠ*�*��"��2������i��2R��ZZ*���((� �(hh������(��"���2ZZ�J���
����h�2��j���������
��
	Y���
H��(���L�3��*�r����3�#\�
"�������L�!�j�L�
(�)�����B���r$h��)��i"�0���"(*��L�!�� ��2J� ��j����̰(��*�����������Ȉ2p�J(hZ
���32��
����j������,��"2��1ŉ�'(�
2�#����;;���}�ِ�ҥ#�wu��B�b���t����3�mĔ�V����� 
2�3�7u�V�r</�\����[�ٱ��yL��X�L��p���܎tb�7�=C_a�	�f_~�ve��sX"��4��5♁�2���
��p�=��/t�t��˔�)˻���u��[J-��@�X[^��bҡ���C��kӓ�<:jn��:���*���SGY�|R(k�ݜp���ل��"�Ba���D���L�O���X���{����;;�w����޼��ʨ�WS�~!hXkA�R�D\,�规i�	^�|������-@n��.�[���Q�l>�s��|#�^ �A	|�(�5zV6d�������3g['�Fֈyxei�|%a�2=��I3y���l+u���]#7��P�h`X��iNk��	�:�ˣ�Vp	�&�v��gj�`��o;��g<�h:*��A���}��3���&�:<)��KI��\5��|&A�<n�
Ϝ�	)Ѣ�����:��DI��!���Ta�Ш3UdS'�H��Y����=�x�Ҕp�b[����ֱ"w1�$�LH�O�b,s��$��R!}C����ZU,�8��I��+��He���F��iL<�"�M�譺*̥�ٵ��{yhM��n��P�0k�g.�q��:���]9<->N�1�/����V̊���r�j|���Vs��<���Sll�������m�H�2�z�.��\�S�!9�04r{}�:tC�3'
'6m��t)�ܕTq
�N�u����2�JqC6h�oے��P��K���:yd���U�7*�E6܋�K9���z��Is�j!Q�Z%�?i>����U��ξ��eO Fõ���U����d'�
��>駠=�e�/�Ud�ǰ;��\1C�@��\�c��B�҉$��X�u7�+g���������b��8%WpSZ��'G�}=KC�@V��2"z[���j��m�:�x�d�Q���eB�����)Gj�]�
$؈�O7�y*�5��3�{/����=�!�ҽR̚�w���z�W\���D:��\z!l`95I5�NK�n�$;f�uLܹ�J6Eb���T�3F��i�İ�쮏�W�gU�<ŭaWk��r*�y[�F��ۆs�j��ӑ�~N�!�n㭺�!-�թa�/oP=}ϸq���(�'��؆]֪�6d�tϯU��G��O)B���j�xh�9X̨9�ѓoݍ�|�˳|%r�b#x��٩��ެ��?{���wme[;��Ԙv���%Q�+z*P�t�[qN��(7����kkf��MaC��>}]v#S�a�ת��N�vɮ�%��XԮ�ڷs4��]d����2W)O��´z�x��Px/O���XK\�������Y�>���k������ �/�D�l�����9},;�d��S6
�����Q��ue
��7�qn2e�p�A1���1J���Č��9$�6(�]]��8�,%��,"E<2�ˌ������R Ҋ�b�Q��c:Ij9Ch<I�MɆ�5���`�kO*+u���^��i�}�'��^���)E{"���;�
��T�$�/N��~D!�}5����^���������z��s�����5�^�h�ޫUi�^�T�$����rE�Y�V�땖|0`c|@,��~�v-��5�����S+6B��z]�]�cӼ##D��0I]�ɶ�k�!
�H\�Fx�`t4���U�P��6�Ui�V���\���:�V�K�Jf2�BV�!�}8�P��B���ȕ鍨��颢�U.Wv]-F75ok�CvB��9q`l��(gH��]qP��k�%(U���y�T:�u�pj��QUTvX.���-�hv��Y�8�om+���7���༤oqj�@95����g'*�^��{���Y���h\��rW���9����r�ƕ̣|�_H`�r.�BN���5�L�Φq��y��6/V7��=.�2x���� ��d} �d���ʱr}��6(�k��7���ԋ6�x�����g�*��o=�)���t�J �LH��r4���9�Ч��qƸgj��������a=����ܻ�C'L�.����τ)�M��P
땇�6�P�a�:��h��fF^�q��P�;��к�\Į�2hk��A鞈�n"$�t�GjcOLxH^��c��˄n�.�xj^��F¹w,t�y2%��1=R�^!�}���q��Kր;��Վyi$"ó<U܂r���:b�����E�["�&�]M�Ou>'��imu���6u�x'9�0�9���l�z���A�uT�5�������j�7)^j\n�`�7�; ��٪Rׯo	Yj����n?���-vH
ޡ�р҇�m��짨V����"|�b��BYS�˩`����ī|�T�t<zE=�6�>Ҷg_�t�F���N��2�ғ���6r�)62�3{�LG&���n�tv��uV��̣WLYM�A��C8��ֺu]������4���$��=�8ƼD�#����o�ۢ�!=.	��Z�*4sUv�F/4+�V)sd��]Z���.��l���'f�u�Kq*9w28->':�{�Ewo�x^�묊�:Q��r�fsm��4]�m/y:�+z�"�#�*/����\�ɠFlS�Ua�Y����	�=�a�SW�J{ݳp�,dq�C'�$�S�ߵ:���gJ��eN�+��d�zT�0�����}�C�Jc��u|��Ȇ��7�`׆l��/�zYpꬌ���	�{���Y���]=AdYz��yϣ~<���N�6&E�"�0xΩQY�����ҫH��U�d�=�z:�7O�Ѯ]1��Q�eͬ�8;�ɅPژ�'Ԅ�!3�(��xY�}���t�{r�$J�R�-H����k*K�hBx��3��AdJ��y�"]s����8-�y�4�D�e��!8{ӎ0)�D;=C���xBUG�E�_���o�<�P����Zr�r��qu������8��{��y_��Q+����d1����֒�;����=)ۭ��;�$�a֛qD*Ka�s��WEb}ܝ�+�������K�$9�nrGd��*:�]�QoVp��,�d�:�I��}5>&�zh���g�>]~V/?o�MfYǲ�Yy�5�����\hE�NZIMP��ˇg].i2;R�*0к2�;J��<"/.hO�O+E.��0�u���;N��Rk:+4�r��k<렵�p�Nە��^uܑ��޵�I+z���Qr�;�i����"d5�hG�-P�W*7;�������v+��뛵l�P�G��ƛ��r4q�ӷ�{#b�R<�R���=W�ʖ�m�\52��㵄#[�-C��>�<�}֟S��wR��9(�߸qu}�6��^*�e�C�����mp!S��[�������w���M�������q�0$�����n���-d����4:L��ɑyR���\%ۊ����)ͭ��6����cb�,pJ���]�J�[̊�� 
�m���$pt�\׈���B��v�&<C��Ѽ)mL��٢��nJ.-W.�]F_��ç�N\Z�
&,��E讼-�$��)�gXB��'��*$���2:�� }�;�(��w��#�8�cUvm�Ҟv�[�7]��v�2���P򣌃���uu(�&bH�
"+ծ�㩛��Ia�ūP��8\�KҊQV���Ŝ�pSZ��'G�T�-�
������FgcC&�v�D0��pQu�x���%7���"(:�Z�]�~�4pX�⍏B��%�&2��f�v�`�[Z�]r1ZO��sv�hœ�������Ő��e�o:�,�qv�2$�p���ū9��<�<�f#b�ΞX�CdۺSv5]�آ���X�Ȁ][�8k�!�wW]�������Np���z�;B�6*�a�Au�<l�
.�b�	q(�R�0f)Jx�"k�p�y+���W�e��T��\ڇ�(��VGg�P�Ű�ÂGxjмc��C�<X�}f�nF>^Bv=��
v��4�c��3�E�:��Z��'�q˂�}�����-�T����~�CLtQ�ZM*6�]⦪�̜-�^��}�\<sP�VXpp���ݞ�;��N|�j�nUu���W��Oʂ>u,%�TD��篌�H���姦�ۤ����3q��X��q����LlS�e0ׄ�3��h"�G��T��y�"/C��"�	�*{�E؃��c|�T�\jPY���<�|���;J�h��[�=�z������UO���i��(oI/D"�t:D�~U9&���)2�T��L�}]#i��^WTĿ}�'�W�=YG��8=�����}�#-�~��5�|!���>��/��-��!����&'�\�4V^)͊�c��UEf� o�ዄp�ݒ;5��D�>!�Zy�o�bZ��Q���e�ܬZ�%ۑ]�#,Ow�"������tlug=~��J�V��WVVn��B�v�#��nT�R�#h\�^:���YW���ܗ(:��WT�3@;A�gq���G�+G�j�!0�v��c�/�C�Y��C�2��w�1��B�{�w�X�~-z�e'��|^+��f��<��M���7mߨ����u��.��*�i�#U�Gp�:%ٳ[Ւ�oq���[#��wr�#��$��)���Qv%s��!�}7�|��}r���e#��'���<f�b7��r��ԱZmC�U�ˈ��E�~W��F�-yĮ��e���;
�fl�O*�S1ou�دN	,��LG�*!qn;\�f�9Eߥ���9��d���$�Uf!;�g��ɗ�N�k��4�>U(:���u�>�O���V9gy������({v�QS\pj/ry*ġ�s�]��3K�F�`�2!N�I�Da���*z�W�"�;���<�wv��]s�}�0(���ZG��
�]3&��Y��z"���`�"��F��jOL�ٙ��'g�Ԃ��=�k��-��
Uأn���!DJdK8�2L9Jɝ�0ff�w�.p���W>�2�S3��/"��1��-�`�\��5)0�&:�bݨ��:�}Q[[D7ɉx�31=E����������0L$@�b�md5sվߐL�􌢹G��\A���v��&���I�����k�4�7�]A�����Ʋ��+m5;W.w��5�BmhΖ�f)Y��[��}�	���|�g7FoKV��Ҝ�b���|V��/5�^V�ȥ0C5^�Nd�x)`�q<p�a$0�Xu����cS������_%������\��	��n!��E��A��b��ܘ��0Y�,®��\���s���`�e"��A^j�X:��v����
?9�YiW����k�h��x�3'hJ���VǪ�5& OV+Gi�I� �DC'K�	�9�(�ܧL���Az��'�v9H�e_�a]z�z���N��<'��bٙ�D_m"+�Y~K����GR
&I;,�=�xٺ�Z�d��'J0�L�]�S���o��%�9��~�X���!����i���d�bʞj
cغ�63T�n]����/C�u���z�J��;�����kv�p_�P�5��GYt:�b~~���TEf�3�@�Eׄ���1���c��c/V�X�L��w��B=�Ҩ��>Z�ш��kE��Zꯟ�f-NL��̵͘����~��r�E_�+F��ߝ	@Ї<pX���\�jW�ɥ������	���v7f�ZHU��Ɍr5W:�"� ʂ�FZ��yO��N#��71��R���3(|��v���&Q�����k/d�X��m��*��{��t9B�6�Ψ�lviU�I�\s�m@̹�Q�P��1��d[�Hzf��1�z���o%��p؉J]k�!�f@��9��`�,ے�Nou�<oS�Y=���ٌE�<v�R��E���sۃ@=�yps���s�
���p;�̦!P�3_v�:���n#Q#M|S��+�%���-�cn�Cc�BvfW.5",�3�&Ku2a+˽�O�.����d��d�ŵw�oZ�(<3����SW�8қ�Ӊ�kS�4����a�i����0���&�P�,l")��p�	;��A�*Y��YB7����u).l6�����������<|
���<%x�<N�.������O�{��A�ȟx�o������- ��#"51!�Z�1:f+ʃ0d*�~㴘�����Jux�
E��&r"Mf�k��\m�}�]:I�#T0.���G�Ga�Ni��.�)Lj��=Q9W�^�Y�v�<�ry$��L8�����͚(^�X���.�d��']�;�z�lUFz9i:�=7n߲wx�P�Y���8)T���=��Be�2�՗CU;���0�y�J�^v��k��L��i�o�&a�r�]a"��/������@��Y�_<��_N�^Sπ�+4�l�����\�J��&�! U�����W,��<�wD61���-��W%�,a �����U���dT��j��T�Ś�t7JPb�T��!�`�\F�u;b[�};���_m&!�J��ԅ�Vb�֮h0���H�E��P�=X��C�6�a�෕bܭH�>�Љ�y����h]E|.k�%�� ٮ�h�s_ɧ�Rռ�Ƶ��V�V�=M��/)70l�)$,Z�\����AۦȆ�[x�Qs�-TR�ʵm��Dݱ8�#��V�+�N5�M	���۝�]���o9:�j[�ظ�ǝ2�%*�YtNgtŝY{��O�4	Cl]�d���[�2�n�[Y]Y�H2��2"���W%'�Z
+�sSK��x�ǘ��ʝ�w �e�v��RU�|"������;it�j�L�B4�OpoL�f�ҀP����ح�aG����JR�A�ҹgb��Vst~C�V�����}wK1FBzt�*_kh�5��ʵ��P��;DS��[��+���gr� SRa���zs�16�����Oq��+�k�Ř4�F G������D���m�H�+m��'z,�)SXՁ6��`4wr���hV2-���K�]���`{
n�4�<�,�"�tl�Dp�ڠ��y!��t�9t}/���;�e%v��čJW�� %iȹ�(�����f�'��0�iQ��h,V`�<]�T���&�\���_fg8������kI����J�������A1Ini�d�"�� ��O�Zȧf����Dư[ ��[������4��3^*�4)m���m����xdY�/2mm8dP�@�����q>�/�Sn!rVb�u|�h�����w�=Rbl�Y����u�j񚒀�0�)D�N��k�w��뮧��j�[�I�lt˲�-M�q�:��Z�(���Z3o��UW(��kS��뜦o,�]L�wm���;a�m^�R4�B�����j�*�W��|�g�TV'���f�:R���~�x6H�����yp�u�ȓ�M륕�ή�����sn��a.���5{/����[�[}Ww]+S�ڐ�0o6T��Gg*�X��O`�RɪCR��6	
�٣�8�&1O���:�ۖ��k�3�I��V x��-ě�|�\�Zm�p�-&m�%\��}�̂b�eF�b ^��] �����&�F��t�|��ܬ�;{֣�����\I��c�u;x���2;)+Ep7��Ά�(�����0�cYP�� {��VR�����g;��n�n�yZ���[&���Ҡm�4���5�	��8������`<���i���,[�X\�=CwDۧt���)aJ���
�^;7����^@P!w�Pq]�����2J�1��2)J�$1�32��32�(Z(���h���22r0����#���J	���3)	���i�2p�(�)�j�*�*�0�������)(��*'0�*��
Z

(,��+3�)
i�f�� ����2((���i20�������,���0����1�)�Rf�"�""3r�&&*
J*��� ���F��2�)�h�������32&)rb��
����13,������032�
��*+,���(���i�(�
))J
��> | �
R���@��:��d���;�˨RG�Gٖ��3��􅥙E���	��V�m�%�V/�b����|�V]LEيC���s��S�X{U=��p��A��hiWT1�6Q��WT ^��sb{Eu51�j
���ۣ���]�[�e���ɅC�S��[8�@�ܔ�[1{�j�Tn��+��Z1!�.��δ��P�O��u�S�6pJ�
a�SS�x9�Zg��Ѧ�|ҶH��0�.��g��X������B"C��m��)�B�6qe,Oz���Yis��fM)�X�.!l
(څPߟTNx�����D��R�(Q�3=ҤGخ�MY��技�����{P��Q_������� K�b㡣�^ɩ5X���-ܷ�\��V�U�k���A
U���&�����o�锻ίo���r��������k��Ӻr���f$c�
5�H�c����Mx�!���È{��*����!
'���ޙ��:�B��3A��f���x�v`�Dϧw���p��W+Yǝ�$S��n�rX�mEt%�[�V6)���r�8�~�jZ�M^����s�[���1]�7r��rt����Up]X�Y[gd�D5670�/6�]�1��\+��e�[�j��=ϝ��|�b8��Ձ�E������Iy3U�@K�=��3΍�Z��ó9��4e�� ۋ�L
WeN}�{\Af��a���ќ��2ap�����1�|]yQcb��=ᘣ�1==�����Ϣ]^�a�
�uu)�cDICzI{�]8�$�b.LUX��hu+��uMooil~�̈́�GB;�K�Y���2a�u���(�=�8��í�R�ԵD\C����,d�yg�u3󣉄���&�tk����7��kH��ʿZWx��jH`����i�b�f��G����bQ�5V�6S-ԎW&!MR�x�<�)����<�ӿc��a�}[ы���c�x��Q�vt��U���؉g%�r/^���7j��a�}{(���(�QŹ\�qeV�cT;�i���dVE�V� K�Vĭ���+Iح�Jh��mK�[��ΑeZ��N��^�	B��#��샸l۬���� �(�"
�e�qu:���>'���U~^�)eߥ���aNom�̎7Q#�L�<Q�0���2��{eTp�T
ܣE:����տg/Cy���𡘒�>�4m���<� �Vo-9�u�% �wp�
���+���w�ް��Y�~�fR��!�;�ճ+��Y{�B���P��j�$3hA]H��Q7Y]jFD<���͗��h����X�Aݢ�mh+�t�=�O3������&�rB�%�vA{��[�4ٔb^��x�X3
t�B#��逍K�������ZD}�/}�LtN
�S{�Ɉ�B�B���.��@k����Dh��Y�
b���������p�,Q��;���g#W�wb��r�(X�#3ꕓԴ�0{��7׾�����x���qYHՈ��3��G&0�WF/�a��V��Y:�f��^�Yg&_�߶���/�$��z�g�š:��;#�*��7����xun��eX��ފ�սq��:����\��<U��Zq7��8�_�AG�U��y��Y���ܖm���K9�A0��f��@�H�%^j�V���B[㒝�	�9�Y�
��֝��7��sT��Ht�&V$�F��a�b����0s�*�5�0dp�'+K�L���e#��m�y&vM�5;U��:��p�$v��ڝX��:��
���g�����T�͊y�����w7.��J�F�,6�M�*X5�(�~���5�p���_g)�+-���jY\�<m�7#��n�d|��H�>S�Fo����twvfn�h��ԖwB��	]�����g�b3"��ZFh.���y����b�D��6k�-)c5��6Ӯp>�u�d+��"�VJ�����D��쓒lAs]Z� �����57�R9���y��tpz�`�2w�,�l��3zYpꬉ��O�\q��`��<��4+<�Y;�����a�E?X�9A�5�(N�nc�(�鋗���?9����~�F������׋Ioc#R�pn���G�L(�b:c��səX�Dk@ʚK��k΍[�Ƶ�%ac����n�_�r�jݫ�����<xX����2Gh�\e�y�k�
~���YU��$N3yzD�.��G��ulap��NEd�P��bfi��ߗ�J����gU|lMI(��uG���;9����'�やDJ`∿�(!�����4Ryj���2圈��F���5}6B��+U�o[����P�g�v�;CJQ�s�s�R��]�>��5�Hʹ�0(Os�G���<�&���~����G�y�4�E���xM���ҳU8�+K�\�
>W�Ә�kѭ6�3�d�c�*�ڷ�D��iV���EP2J���}]������<8�t3��_I��se�Yt�=���m� �ÇţLm�N{T�e��\tt]"k�t��
���;�(f���9�����P���O�.���r����{�+]�]E�&
�)����j)�0s�J�7i��SÚN\�O8�F��p���y�� ��S�"�r��&�z{���-7��!��t��+�A]�^��h��@|�V�F��&�2��B��a�RzaT�w{$^�<x:���٧��0xj�D����v��s�� ��\�z�x���/����������]ѬL������ڋ���B��X���G�t��lMxH��޵�W���#`5�L�z�ʙΨÞ�*b�+ҫ(d�ur�g�2������9Տ<��TV��R�댬sR+z�58��a���ȹ�(�#6Ur���Ub.�ip���`��_�Am!�(n�i�ڝh)j�f���{"�/�p��1�KS��pM1#O\ GT��
	&�
�Y��y[���ÊW|Q��w�<Z���eK��¼��ع飂��n좮�3����z�썓}�~�H���qe^���<��^��"c�y�V�,>�_16�D�ܪֲ�R�4��6�Y������>}�0EU�+|gQ�*<��S�)���L`�K����K�Wv�,'�����n\ڇ��F��
�.�����Co.{��ea5���o��e��fzl��CǙ��Vn���Z�{LlS�#eϋ�>V����{.p����7�va��!��[v���ڨi!��ՙttO9����c��\�U�P/�Z]g��Y5����J]���Fh�j����S���wr�+���&�3�A�h#�9�1q��K�>�<|�)w�׿���!n���o2����Gyj4�E%4d0�#䂎{�D�v�����}{h�VQ�Ҟu�^��!�(�ʯ#'a��j��Y��wL\�)1�e1|x�OEu�{��
�fs^Ү|��������%M��uV���H����N�R6X7���s���վgE�r��MdGhП&�,WVR��<��,C+h���bX���=����#Qfܾ�tA�z��ޮ��z��>φV��l�N/4M:,���8�$�����9[=$Ƿ:��ǥ�=L+]�%t��=^��(�βZ��ٌ��ń=N�u���)��ł��e��(3�@r,�k�c�T�9���쇢��X����x$%ĸT3�}\���s=�E�ӕ/Tg*��y�¦o��P�e��Ƕ]����~*i�&p����q�s�h����:�H;�^��^����иFe«Ɲ����q����o�YO#G�b���Y�{(u0]��a[��U����%���[mw)Ƀt�OP��6Jɂ ��=q�m�͝.�3JL1���RXy}�Ɩ�uڎE����<�J����%�ζPې�"M���歈��t�\�9V�3#���h�ڸ�¡u�@9F�yZ������c4N��(��$��r���·c�}7�P��h���|Uz�G(��ۿ{Lf�WX�5n\B�l��3�QZ��������"Kcɳ��0?.��ןKx������@�1`��؎4�Dq^�u�1�4h[�]��}��|OK�|�i��龾�ZtB$��=P��P>⶜����)�/����G�k��Ǜ��#��w��k\Hy�x�C�H��U#4T� X<�S��Uz:`#1W+|�E����rxML��e��.�O}�@�=�nZ�.z̹J�|e!=K	j.�6�^�������I�D{�g��[�^�z��o�9��:��,�c��QI�,�l����n�j�r=qN�f>Z$��c��Al�y��/w��#(>��{��3�����{ݲ��NVm'��t�S�ПԦN6��Qc3U�W�S�۽�!�"z���殓��qƒh*�1^Ti�4��;RӉqx^_��A�4�>�+ �z�*s�����D���wDݩ�����a���U�,,'{2_V���b���k��:'ڵ��sN�P�9\�3��V�+�n��A���v� �#;4�\�u��G��aWR�d��1s�����w��.VX!�jK�ŅR�A�eG�u�k(��c[��D%fAz٘,.�^�G�+&֘B��:ɀ��p�*{�?y]V�|��(�f�9^u�K��<!�o_�m�V�,���
�1����Z���؞��*W�&�t
��&����s�*��0g�,�\k�*jW^tq_��̼�D�gt㳻8��6�#~ܚb/cb�u+S�)zl~�b�oB��Z�X,��)�m�g"�?7��:��o�D�vi..���e����<h��hu������x�T�'�N�,ܕ�3��t���w�Z�F�"�}ב�W��	�\`�]ez3�o��p���;��8}6rs�+��[�-���aB�2k׿`��^r��C���,�,WbW��7Y�eOc��2bp�F��]|u��J��zĪ�lOM`���&���&`t{���+�̶s�̽�q��d�Kb�֨qF�+��F�h���J���G�4ؠ&t���.�5�#Ll�/Wqzw��B1�7�C��:�1�iT���J�L����'V�'���x�3:xеT�<T�T5�E�������p���5�4��&\1�]�2����wA�f*y-���!�M֛xe%Wg�9LwoT�:�eE�����n���]]j�xg�	���O�����4+9o����r-�疰�����O_�#Z��*u:������V�"�#Gq$E	a����*��R����
�9�l�G^���B��T��s���[����B�$;����3��D����G��5xd��4y�-���6���o��i�a]#4!�!����T�dЊ�z�Q-��q%HfJ��י�ꇭv�$K��
��p�x9��QgƷ�T�pΗs=����5gڋ)��������N�"͌"Xp��V��3�3ND�xD��N�bc+��Ds<���ٛƶ��5����h��q���@X�UC��`�[�^�^(�2/u�iۘ�+5����|���e�P\&��^E mF����ɢ���e�J������{�;m��qw��f'Ὢg�E�/V� �YhX�/�gIʥ�UH|�:�Y���T���!35ߕ)bIg���Df�4�߾�A�q�j{B(?��e�t�2�
��o�}~>���"7aX�N+ϗ�"�'o�C�xK~��[췘_r�{���C�l,��Z((�Z��:����8&���
����� ��v��5q�ޅfs��5�CD� ��*[�ͥ���&p{:��<����{�;CC9�}��a��mg$]��&��9�.�S��VV������e�+oh01s�'.a�0|ˈ��i�v�G�y�qNH�����{LQî]Wk�{]���J/�9��˦�8;�|N�%_�g+��*yg?zA����|��5��V���	܄^9�YEԼX�B���n!:�m�����<K�3QO���QɆ�mfu�?[�F(��dYG*���.��x^2A� �72��A�_HW8s��])R��a�j��3��>��ѮS�)��.�:�ܥU;��nr[J,�e4xi�pg|�C��,�6;�޶����)Ή�*L�kZuU�*�)�gf��vl�ěO��|$N�q	EtA�OL�$��b�B.�Ǩ"N�����+�t�8�W���Sw�N��9���o�z�tĖ�'�e1|��Y����$[S���gW1P����;p�Y��c��В�b���gK9J&C�Tʂ�� }j�%��r@��DY�#cf،��L��Y�
X��5({��uּ��=��^{t-����Gլ7��0����^��uO�(A�N,h�(V��`��nڲ����^�vJWռ��{I�6q��'���@�S��dz6��^O�K�iv.�laol&�d� lR�V%��	�M��,j��y-ʓ����Z� �����,[L��w��S�j;MZq���6�Of�L1�U��4I���W�l���l��!
Վ�jkI��xMZٗDл���Ǉ�Y��La���ì��-+�u�R�|^��ۘ�ɳ5�,��#T�8�n�]�D�r̂ֻ�N��[��*����� dw���Z�5C��]�
�Q�����\���
Ɲ�ฺWc��4�2�;5*�<,p��ebv������f\���d�£�������GGZ���K���V)*X@7wf��������u��رtڷ�Fn�uYEN��ʞ0�ݾ�*���y���u*�u_�5F�`��[4����r�,���d�p�E�<��U��y6�+�z]7�CpvL�h�5�(��o�S��ս�)��Y��R��3��et�[������Nc�I�S8�bȈ��I��P�{Ѝ��
b��Vk��n*%[qoD�b7�0��d��qYP�f�=��[!9�w�l�m�0��^hN쬣
��=D�yՕ�� [7BʰW@ �J�,>���t.�7A�z��ڂ�+vQ9	�i'ժ�7���[��˭�]��O�#��5%e�\A`f�[�l
�����t�SI�u5��;�����hIc�,Ԯ	����9CZw�lR;fX���5�����k�vcw$
";�8�V>�)"()�RY�x仳4�Yq�F�rQ^�<<����͵y<�<�c���D-�:�dU>��ژ VC�o'_g_up���d��Zԝ��Dw50Kl�6;��P"�������=u�� SUZ�J:`ݮV��*#���j����uv�}�p8���Z��ГyW봐�����2��o�;uc[�LZ� uxx���oL�B�]� �i�E���n����ќ@N�%[ݼ��&�t�d�Z�҈I�niZw+� ��k�E6w"�[̫�2b���R��?nQ�z�/J@����C.�Ζ�x����Q��u�|#���_�W�Y��<F!WZ�R	�����95�f����,�1S��vQ-]/�rX)����#��� ���L���hE �w�w��q�U�1�5�[�f�ċ�:��=W����N�����q	��'#YZ1ͻB���ښ���q���8�`/+�Vqcδ=�Rhi�.r9��Q \JR�u��F:*�����ر�/*�h!{e���*�jQ\��5hP��'Kl	}�XJ��vWU�;���k��{P�c��/� �y��q��P'W	4hF�LYM|���m���^�Wՠ�� (&�"j��2")(��"�r2B�(�h*&����)*�2&��
��)*�i���f���	��*����Zhh(������")Jf�)�*�!��*j�)��%��)���i��ʦ�j�	�B(�h����*�"�
����(�����*$*��bZ����"���")�ff��b�� ����j"��&�)��H���#!"�r�**�3*)h��i�"�hJ���***H�����"�H��&����(�j ���J"�( ��"ZV*))(���
"�!�"h*�����"i��b��b��b��( ��&�j��h�����}u�g����4�X��Rƭj��k"�9��Z2���*�r]�ťǃ��ҨVܕ�@|5�W��J�6�Lg8���Ru�*��7ڲI#�rLP|�f�|T��g&l؊�cp@�va��2X��Z!
}3�p{��Q�^��7R�N����y�ʜ�/,��bg/z��]y1���̙S�Jz�����V�vyG�~3a��#�׵S��~{ս��g�Yʿqh:�[]5���^���׮\��5*��X��6qC��1ņ��v���>2�U^4��}(�+���v�2�S��}$�/{����VK?oc�l�M{#JF/��bW<��_E��:݊i��MB�c�瘻xL�������ꞦN���^'����g�h��K�܏}~�0��x�$>��3J�"7�E��`���czvb��U�dY�SLk�b8�Q��8���,�F��#bg�=���s����s���П 8k���g�J������x5Q��:Ν���I�U�j�^�=�H��:'��j�o��H��mZ5nH,�`�%B$؈��3����mqC�b�qs�ee��T���:��	���Σ2�B�<]3'_��L�Gke@��!��ީˌ��i�TF��N\5�'v[#|g�����=i;�ʏΖ^)[����ӭu��ۘ�dП���D�5]��Ƚ�2o�+�L��ĝ���/��Y���寷��ʚ�$�X-R���N��QuD��u�(M��^ڇ��@z���Մ��������q}�j�{�h.�D�����R�;lӘ�r��[Ҧ�\�Q�3�Q�aC;0��[�����|#W�,	
���lj7}�Z��g�&gj"z��%.[KL��J�=�a�-��������$n����˽���Ġ��YdH*aki:�u-'þ|��O�BsmQ�8�C5B9�`�Q�&Ʈ;o~�԰w�;�x?$ʩfzLHx�{!`��ٔDO�=d.>ܡ���C��Tvzg���.;�r�1]!��9�ȋ��'L��
_r�������Kl��|�k��(Ou�R}�;f끷28�f��1�1�{S�qȎl���L�9喋�}ъ����f*����8KW�|Y��4�XC��U�N�M�}}h�bٟg�r�3ޑ����{ڥ����,#v-L�ã3�M��,�e����49uiy�sC��-�z���k�a�w��k��c��P�j��I�t�h���<�2=��x��6r��w��˕]]�_BL��P�u�{Բ���uM3sC�k W�j�6&:��@��N��z�8�D.S�5��C�kM��;�mw��z���aCF
�f#�v��~�gQ��_�+���B�]����3v5{f�rS�S<��3� w�q�D��)XFWZ�Z��h�>�o�wn��7�f_s���8T��U����z¡H麥��H���h��PsEԑ^�ȧ����\i������<
�,��L�v).V�_��p��ДC�8Ɵ.��g�WNmbl�QN�Hf��A؀�Mxd"��q��ޛP��(@؆��"�ʙ��M���wH[�ܮb���S�̠�h�K�h����������o;ˌ,���-Q���u1Ի���[�L5�Ht��\q�����
�j�`���À�(7OC`=��ҽH�=�{8O�5e�Ż�4�X4�A��J��Mv�&�B���j8|&�2�\���i�6��bģ�����v
a��W�B4p
�i�a�#5�a���z3	sv��(y�����O��zHyġ�$L�+
%�3�j�Y�0���<���3�:_zg�:�kv�h�V�Kc��:9��.'���f�,v�&��h4�b���U�Lكcq�i�#��\3���q�R��e�Y4��I2�V�$$Ĉ�'ױ��"_�ۯ\8��Op�ϲ�����;T�a�1���(.6��O	<��ـ$crp���*�GNP���]Z6bW�Ojr�]�@[��%Gǽ=�ڼ����%LSI��[��w
��J����j7�j*���{y��rz.W��VҜ�Zw1�L��N� �'�����~6�c�M�Wj%"�v,�ؓ�L����'Fv���{:k�j�׾� J�YhW��O�~g �v�e���P͚(���,�ŧDE{�^|)��͗�6��V�g�hj�a��6PkٲٺgC�Z�7�)D2���N,�#ݔ��1*�Y/��'o���8_�A]�ܛ�g-��C�-Nϑ���+�,���xn��2u7�+/�u]3�,�b��Ew��u��P�^7^ڱN��	��;�!yY4Y�5K�53���U��M�:X�b��pH넌Y��J9���_O{^��x�
-�d�Nv+��1���.��jcj%���\1yq=���������9��4�k����鞧��"T8�S��!Жk���*�[��z����:��R��5nBH���ٹn�Þ7^�4z�V��E:���],�ω�3R�T��I]��&�WtT65t�C�^Ǎ�DP]#�-��!�f4c�
+L�m����D�{Gg���Y��e {�1�1��DV:.Y��thfZi�c�.Ub�q�L���z�J[#��u:"�s�Gn)��n�Kc�$4#yf�f�ӜN�ҭ&9VήucCǓ�\�Rq(�m����"eB���Ո�9��y��Z����G)��^��f���y:Ї5p,6���1Vh8f5�3д%Di�>0ÇI�K�[��e���e�T)�|cj�Y��c�������lSK�2ESQ|MQ��rޑ:�e�c����K����������Qb���Ll��g\A�LPa��E.����6{e���uӻ5={3v�U�E�.�x+�<�xg�s�:����c����(u:�`y�����C�Z��cF���<I�NI3���eX��-R��wؗ�����*�b�m�U^�}�����ͨ1���<Uz��JI�GTP�3ʕ]u<�<���R�UӚ�g�m��{sܸ�<��l�8B8]j�q&��o@vl1���߂!oc�,9.��θ�^Z���vӾS��gNK76C��z��q~p�0��[м;'NӐ����ݍ�h�ߗ���>��z�b���f��d4-K3e�w�JF)\�w=�d2���.i��Fw#�KXJ��;AXs�ȯ#����KC��OL^%ު��tzRq^VL������4�gNvQ�I���<�-�q�'�v�K��� Y\\ڿ,�ewf�R����5%��2qsjT�0Z�,�
@d���cXA�hgg��b� ��k���K-��#�<��)-L�r����,��ی�] �t���4��>W�t��I�Y�Nef���G�՝���NZ���YT}���]�}��J�y��V����%hŃ^���q�R����Sutȭ75
��Yѫ'�M�qt%��g<����3AI(�J5���"��8��4;2��\kxν��z9Q�;et_C��X����޼Q�]#,)Fy��b8�:I�C���/-�+��fV�+��ٰ6Vs�فa�1Aܫ�X�dֿK1"�;�V�[�u3o��Iȇ;8r,�(�)f�c2����=����C~!̗aՎ�,��X�S���s����n%^���L��R��p-%�Z���5�S:M��e��x�oK9��Dx�H��p�L�U|������@3�T�zP����-&��:��:�C�t<V����E�-�~����q)Cz�Ҵe	C�8 �|�0�z�0�_�i���)�x���7!��񥅩Y&��RC�Re�����!��=Y~��q����)���u�/�dA�ZY����l1��鍰���zG�!�>��`�����@�Jڲv�u�]�Aw�j�e�sw����J��n�_�ca�]�y�iS�Ԇ`j��]���t�Nsri�pRknKu��yQ�b�[R��0�o9ؽ�+j������+OQ[7&[Qn��j��e)�^����.N�o�Pg��ޛ|t��,�͚b,laWwXҳ������\`�l�p��JG�2�ՄN��a#6-窴�3iɄ��,X���&�b�k�� �k�f����};�s�,�#U�H��DN���­O�{{�Zz�X��	�_�G�z����g"�������p��;�\-Ӯ	���v�3sQE6i��N��s��R�<UU�bkn�D0�QǏ-t�:�V��8iL�=`*��M�M`�FDb�-���,�]��Y�nȠ�H�ەJ!�Fݺ�BW+d����*Fi�mP�X��O��ή�u�W$�4�Yt.d�4%��42WӞ\dFf��>%(u�j9XV�vX�wG.��6�+���\)�~2�4-U#R,h��[����מ��+�'k��ݺ�Wtf�7R��lX��ڋ���P\,�yx<�ন+��pb�Xy��N�r.��-�w.�,^:���\�L@e���Tt��]YcЧ�ب�?�Q�(�W��T��_���ĸ��B�K�7/��;q��V��L�ͽ���5��z�q��3�X\�54K��Su�۞Gm��C�k:���Uǖ.l[h\�/x%Om�pb��l�d]5n������pvuf���V��wWo�VS��Y���P.�Me����o8���7����}���7�L]~Vg���@��^�C�?�é��6zX��,z��jo��ͱ׹3�	�"do;��C.&pPΙ��fkȐG_����>X:�Z���qz����}\��[P`��4�Y��OtM�Ι���o�/&�ܖ��>�y�h���&+c2���y��_�,ERH���	�a��c4^´�aՑ�<��J��_+�˜�q��J,ӊp�&�Yc��/��j��nHI�gq7C܌v*{ȶ�}�_g���/�Cd���C�/���U�:p��>Z\;�j��A�m�쭿eT�%�8u��ȶ�Lf�Vd�%�^PD2�]OmpW����9��%���ˌ��C�4�E�w���8�~֫�=�݊���{�Qf���ÆA݃$*-��~����=�(i���Q�E+��<덂�wE�u�q��v{%��k)�=�g����3�[F��8.e5lOpH��J"�x�e����ǆ��b]�����b5���T���͏�р5F��+��] �-2��3'�>m�=��s۶�U�*�MI3�f�z�ғ���rA�\�-����n�X{�R��m�G�yr�trͰ��k�����E��v�-���w2ͷ�ο_w;�4���s�+.�L�4���F1��6�Q�2��t�zmB�z����utOFMv{�}��"#@�q����m��Qu*P�)OE2{�Z��|�V��<�J6D͉ń֞W�z�dwl�^Z�'�t4vZ��:�^_m
T|�(	��'��f��F|�<4�yr��˳��U*/�ϳ�'y�J7q�ḳ!�1nH(�$ 
;f.]���;�Q�չ���鹊e��^�{l�yә�N�U���$o�tw��b�I��#)k�FŜ��^��7خ�o��\�� jآ:��R���xb�mgK��?���W�;�Pv�g��~6�����KA�r�X��J6�ϭ �(8g�)t=�Kc�"��h.�S�������|�A/=Ja�:%����H�ص�p�8�h�(o�q�Q8�5�|�Kv7��C��}G,��U�M�w�D��I�NKR��qS��8WL��V���E�U[��,P}PVr�(g��p���P'�y�V��~�Ǩy�L9��3��m�����.Zow{���S����z�>D��|@U� "�����;Ӟ�ͨ�<Ƣ��,5�k�b�4.��pm�{��>Q�{�@�i�kI���l�#�w�N��5&n�q�YV*m �^m���r�������,K$���Ӻ�ULn@B(���wl�_(�t�g��h+ׂ�'f�
�`*o���Y�s��Se��GNK7ٲ424�n��q`8uoV�g�mq�m�Ȥ%5`�ɩ|��j.�_���^X'_��bu;nX5�,�Y��#*t%k�����_U���5���5��K�PN��w�#w����8��z�N���^'�/�t�)l����#�56�{�.{N}9���~��\c�vb��U�dY�Ń\`�'�Z���	�'۫�{�Ugj��,b�E�J,�!�mC�zx�)�U̞
����ݪ��g��(:�M���vk�F�aODq�S�/\��W������2�F_LΖ"Ƽ�o�1IE�4�,�$��ODr]���=}66Vy���B�S��fIM�ͭt:k{3%<�|��Xhʈ�!��S��,�Ҏ��)��7\u
>~ݣs��W�z�g6��>sJ���16PR��KIj-���yDu'�X�jYa��U��u�9��Q��}�f�u��96�p������S���lq�ϋ��c��ܤ|��Ji��/���Ҥ�&�a�(9F���]q�D���Z[��e��+��J#���֫S6ub3�ұ���u�^B2���/I�K3��dW$u͕p%�ir<�U���3�ՒX�)P!
ߊ0�|ON^9e��#S3�N���7���6�tF.NX�e�0�p�*U�� �վ���x�]��A\hk�ZFv7\|4��e�b�)pZ���z�`�T��*���E�t�sy��X�Q+�#�O��6s�v.��G�h�i��9Y�+�5K:
�z��)s�[Z&���� P�ZB�9'�.��Y4�"@n�+��j����nEst����̋�X,nub#ӑ
�{�7-� �J���V��J��؆�Y�T-�.L�/�3���������X�Q�=Gk�Y����;��;-<��I)m���ӣ�f�mɜg:z��gN	�Y����Sn�s[*L��Kz��H�O��U�J>����R���"��w��ʻ@k��(_�W ���d(�o�ꝑ1{e��0ڴ�朲-vh�Ŝ^�,�.�*�p�MT��nǰE�sy�i���W�:S��eGT���,�W��-u�*��xV�Z����/C4��nM�Z� ;*'3L;y��)�.�K�9�u��'/���8-���LȧnS���**ȱ��Or7\h���,��G^��5�D�M�Y�^Ե�Gu6�W�$;vV��Ԥ-�('��^wëMf!p\ʶ̙�;�(�
y�]���]���s,�+MX���e=���8��5�0���a؁�9d����jK�P%�.��2�v]C�#y|s*U�G��D�(�Ӽ��>�[�읗g	���i�_5��d�=IQ�$���F��V�mEtB���$r,y2��]�D,���V�7�uK���z�u�,�h���M��0EG�+�zZS;l^�"��ſ֨��j���lu9�H�M3��W�k+)�v,��>��s�F�Y9G�y�
(�x{Q�5SA�Ma�r�,�Z�=�0P9㤺o���4`��9.�3SPAQ�WI���R��W�sS{5f�aoL{sS�]�q�v�����ʤ_�S���Lj5٣����7�+Y[��.�]��9��Nk�[[]�z�E�A�ql��N�5������,\���u��T�{/��;W&]H�Y,<��cv�]�-L�\���ut�q�vՄ�#0�%�9���$TV�ujnb�.��"�:Uv���tWryr�gF��.�'IWI�����B�<�+$Ut���kK�`�*���e�ha�4���n� ��R����XPK[qF9�{ZŘ�[J`U�X(⺷Ճ�,SI���X�����Q,�3(���P��H �@D�T�TMA5��EDD�L5ERMQMSD��ESPDUU�D�TAQUE�TTMUEDQARQ�U5TAST�DQAQE4DTEQ�L2ETD�Q1U4�USLVfL�A�TFe��Y5��T�ĔF`d���`DU��aX�Vf$Q��faP�AaQ5�I��RTQE�R�YTe�ŖLQY�D�DQES5MCMa1T�ETFVd�ĐUQC�DT$PfdUT���4�T���VXLQ4E3P�6Ye�U5DEDSUY�ELYeEQTSE$Vc�MPSS$ADILU5L�TQ1DY95LQPDQ1UM3Q$TQ��QL�EY�D��TT�QQ9E%�$��� OI�@��Z���"��ٴZ�޼�E����1�Ň+�c9ԷM�>-�:Q�#�+"�OnB�b�Eu��r[Qܔ���V�u�$H5�ĉBh+�B�C7�S�x�4���V�A��f��x�1�� p��H�L�^��:n0������u�CP���-8��^^C���>��Rh���uZ�$��H��j�J�ɛ�D�j��y����WA�^��݀�Z_=J�iW��z��aC{�1׉c`^�;.���ʲ�*��w`2%��{o��~�e��͜��GM�:f��SM�Ǝ�U�Q�W鷤����gM�y��]~���r�T����׹uI����n�%�����,P���5�p�K��Tán3�P��{"�j��(��)y�a��RE��-K����h��=�����B��׽�N W����6��-�ti�(�Բ�λ���Ú�Y�;T���n�L��9a�w��˸�Ur�6v#J4��_bUim��3���ap̪���jwG��C�EY��/غ�#d?bC4[0:��J"�J8��E�|���#�*�+F�;���`�ٴ+2���
0C�V�k��^X�w��5��p=`���k�������Y�MYݽ���lKЁ 3�x�7�+�lwKbD!zzF���X��9rU�)r�l�*M�A.�W^л*ILW2��N�q��P]���2�8IՇe)��wF�D�1��,Z���w+�p�e���8ϥq��5ѣ*YYӨ@s�{ӎ1L�!�v.0Ύ멕y�E<a�B�*Dp9Y����7�R,h�Ml>��:���M�aص%8SS9�<䧕�EL_���W��B���j�ȋ�)f��
��$-��>r&\ó̭��i��Y���*�R7B,Q��Pw�'b-ZM�Z$�^�k�t�Is׊Z���e�n,dQv'|^K�ȷ��g�<�:���!^u��^�i��|�88��d��,����h�� �����v:K�g��h�6s�b��ٕ3�5h�t��oV뷅��C��a/��R��R�`��a�B͌"X��ʜ1f(7�*�MR��5�K�
�bҶ��t%�FY��F�~��.%���&��6Fy&(F��Yw{�6�'���w��}�{X���H������S�ȣj0з6��&�Ya�n�]`#w�mRNz`���"n���1ح�E�^QY<mP�^���r�|ǬR}�f^�$W��Ř̳�ْ)�2U��l�ʇ%��T���8��Ǯٴ��W����uqLZ�뢨�L��	���,^�7Qƥ-�9��-�ge֢+��'��c���u��Rmg���L����k�	�j��0�K��8���M覾y�{y	r��d�d�~�s��æ�mnE�v��*7k���*$��=�����k���j�H�~�`�9Ё��eE��.�q�ƵXE��݊ī��j����[(M6ئj�U�l���o.�N��-�h\ GVJf(�p���nROҊQBگm@̎�ѻ��6�ff;�1M��&Ҽ6N�/䴳^�'��D��H��"��Yu/;F�5+v�9�CLk=�/<q�N&f�9A�t9H���*h�����R7.TB��e�)WԳ�-�`���s��=+�?9ӹ���"D�Q��LVŃ���k֪��sj�7Ӯx�����o!�놶`�f�����CV��S���hU�|��+lW5t�ލ�����P����L��9΋�{9:��z���n�ȿS��W��Q���#bz"�C��*v��;�B*_�o�i�yә���I�8��A�w�厬зt̚�:��ؓ�#^.�ŗ� j8���B\�7^�����c��Y��q:���n�o4Ek�JuȜ����͓�aZ�+���P=��,T̬�;fP��@}����'����α�m�F�dFZ�0�~�6�	��.�ڔ[�l����l���H���؛Rp�d�ѐ՚�'sHr���f��[�ej��ޒ�Ki�ŕ��whF��U�d;��\|�z�������]Fa�:���Qt��ge�0�y�<a�{�:�9\�ð�IZ�	p��q鵔�Z��-�@���Ⱥ�a�	G�L>��^O��|��0A��Q��9LT�\�v����q@���H{�8�3�LN�S�+��+ь�����qw��~w.nj���P�`�Q�����G�s�(O���I�i�c�bG,�2k���a�w�������`�G�ys�23j�7��(���9�'�^i��8 ���6��{����8�$��p��;uk�=��RȬ:j��GM�1B�l�fN��UqU^#�zbb��;$�=/��(�Q��=�o�`�/����kD��xs�h�>����g8�3���t{�{�u�(Y{���}�5^�f/vS{�z٩��hX7����-p{W��)P�N5�^z �-+n��������Yk�f���}~����C+SO1��AR����G<��Zy{,�^^q�m':r �:��S�/T�g"З֋8>��xzx�$��%Tp�B�����v0@y��v���\N��WG�
!���ޮ�:�Riޝy���k3#d��z���\�(���u`����w��\[��iշ���S9ty�2�NQ�f�޷/����g���7����CW'3��s5�y�}�`>&��a��!�i�c�w��>��Y�8C�2�Ou]��c�����m{���9�ۼ��Q$�8T@E˾������V��4��g�FeW��_;��,�u�؃^�
/��G,gzQ��g�(J�9e�:�1��zT�Q˿���U�,О��V��Kh�)<�!�z��>O����bB�()O锡,(�������Z2�_h��B��h�Ԋ���~��6y$�[j�����j+*�D����.�맺���)�6_��B��l7��|�@T"iɝ����GW�@��窂��1JX-��`�n4��L���HtI��� Y����I�K9���]�ޯrG�ӂ+�����1�KT_!Jb-~&��R,)R�%R�f�=�}���k��bg�6�YL�un�ʠ��e7X0�Y�#O�ı�/W��,�}1��v-���&7�DC'OX������]�g Ȗ#���Pµ9�6NދO��m�vc�kuwE�C�8r�Ʊ0r��PdFl[�Ui�@f:�~ʔl2�l�d��۩��r2r�;Sg]�S�eqbOI�h_(=G:����،�/���k�ӂ�]ƺ��u��K�E�r�ݜ:#�V���^L�l��}c[,��}��hͧ��j�=�q�Ug���8ﳍ�!�B�'=�Hl� �����y�O_i;:�\��B���p�N�>�n�ڕ8��4_�<v�G�P�(#��<R���8�(�Mh�1�VV��cc��ݢ)�S=��d"���R��ZvܓHPy��U��-9�F>��Q��d^RM�zTEoK8���]io�%h緛����W�Q�DF$���ݪ�Z���x�HH�E3�J���H��$"��޶r����h��BuH��utS��ˢ�r�����K�q������H�@J�A\jp�����>S�﫹����.�K�jV,�!1㎼����������2������@ľ���W�!7��Y�O35{~�]�3�9Q�%f�T0Qu�Ҧ(c�KMp4!O���Rͅ����9�q�|\����g����0K���P��#C�$:��:`T����
x٨�������D�����2�]k��z^zU^CpL�Bs�Et�ס�!"���$.�*�A���^��|b˻.���v�ƒDh�v:/�i�3�j�PΙ�
��B��sb��ܥ]�p�o��\��K#�9kJ�M��ı0wkU��1���j�����R� e-�\���<��w�|�����6N�&���z��tL���\��n�q瓮��r4M�g�� qS׷ �ޛ �zI	RD�;ɵ��eӽ��_M��X�x�:%�ۦ�5��|%ey?������bX��
.�^�/g�u�;O��d�/mq�*�)��D;�e���O��Z�>��@��t�)���2�V(J������LEb`�`�iY�~p���6'��^&:����.�B_��d�9r�;M]xL޵R�".�}{/�V��NI��k�͛q��H�R.y��B��Y]�m�ƻp��crh�7�(��*]T�&��t��Z5׸�g�!�<��٤{�촜ј�v+��0�24��f)`�͔TXWxYJ�+��un�`	W�8�z�mɽ�=��9X���嵁��N�P�`����E�R���s�8Z��*��j��,�Y���\{-���LR��♊��飂�3śb8�$����iN-ł�B�[(-��6v�����.9�nsa���:���~�4p_�x�s�𔼸��Lp���^�����s˾}��j5�����y����Se�Y���`秥S(���W=��Խ�m�9��R�)���_�C��!��KL�2�L{Q�6�5��a1���5�.�^+��zz ��N:�k9��_n0Nq����l��M36�XU�P�n�G�S�{6�߮��e<�:��5j+d�v�J��ེ���[�sVt}8i*��謇����y[�d.��H��K����&�0s4󺨵����=���#�W�%���2��{M�#����;2>�Y���31���{-�vgU�H�!�7f	GkT���G=Ns�0Rv�	�R�x�F���4�I�����]^O{��^��f��8J�j�5ѯd�.��ۅ�:��.\�CIV��Zȷ[�o'%�ؾ��Tv��_EwL�rexWPv}�Ih"�FJ6�ʴ����=U�je��,�4a��c�ǝԩ�>آ,s��X��3�-�a\~+�3C罸ړW��������yP�TJ��]đC�����`u��=^��%6��W�9�^H�$Lq�<X���G��
�x?�^_�5ٜ�
��8K��x:���oz��-ml,�|�C���ȻR1�*�"�mR�p��NZ��I�=�ތ ��	o+����e�et8�u�Cݦ`�kk�+*t�Z�t�S3` l�L-u<xr0a�خ��E�1E�}�Kue1��7�nk�n
��	Mwq�J���"��;W�ˬt���N�I��� vG_�2��f���K��ZHU� %<���
�<��$�^2aN�Lp`�U�m�%�R�u�5X�Rގ8���%v��;��4y�Z�������l��N�ػ�+G���
�����@aY�b������0f�Y&�G�u�����И�~�Od��%Z��ݵ4u�y�~�د��l���e��3<V�2u-���1����\��z4�e������'���(W3�)�C�p�,��m}哱ԻN�3}�7=Qz8Nס��r͛��s��OF�5㳳�J=J���*i���:�-�R�%�Ada����]��qz�Y���7�8��>�.���>���1/�xw��.�ө�d�P(�:I'�=�.��˺���C���`o��Pn�Iq�륏
���`�0g��,�0�7��E�Ap����g�Қ��v����8˒7])W��}��KZ{�\x��P�c����2���[KƔ[N�R�Tޭ-LEr��I�x�o	9P����u��n��rȐk��A��!W����J���o�B1���1�.�h��W�SH�.S��h�PT����q��T��Tj��zM�~����5K}���󔚳nQ�8�{��*!N�������x���t���3�6��Mf���ktsY�s�"T8�E)+//�=\��
%b$3�����d%��hCw�;��+�q�鏉�:�ھV�}�ṙu�gg��D���i�,x��[���%A���r"���1� �KnM��i���G���VY�Uu���FQ��E���a�<7P0�΂��q�"%mM��۹ļ�K;6�!Zc�`�p|�������`�V��/�yV�`8C�C�����'�<�<��c����紏DXW8r���L��T�dfżZt��u��ʔ�e��W&
�n�ej��cZ�6I~͜.�:��o^q�յ�k�T���~E�[B�� �>�!�����Ղ�y�G��Bt^�����E�UY�Y��{�'iEmΜ���'j�0�S�<�f�q[w��2�JX<tR�+zYǏ-r�H�a����MX�i�}�c"�s��b�jQԷ$�Qs�X"
"X�ǁL��R�7إx��,؞T͈r7b��k3��]l^N��s��>����ZʄÞ<"8�0H�ˌ�P�º+�i���kc����U���������JgØ�X��Š�;B�*����z%"Ƿ�ӭ~�>���+��W��W�"* � ����
�+�DTA_
�(* �� ����AQ�"�
��Wh* � ���(* ��Q�W�����ED�DTA_삢
���
���d�Mfc��4�5~�Ad����v@�����C|�TU%J�R$U*�BR���BIHEEP���J*�T�RIT����!@"J]j
�R$T�$*�[j�B�HR"(��JI(�AU�fַ��=JAHTQ(*�Q*�TD!IJEAI"!J��IIT�D��R*�*��"�E�  n�M(Fl���j�J�l�-T�b�QjZ�nZ�A�R��6*�iVѵZl�ت��u���Sm)TT�[� '"�v��*U��Q`�e*�[m��m�XUY6m�b�3eV�Y
�PkV��J�GwRT�R�J!J+ ; E
�g,�  (a     �w ��@,`   �.�Ve)��SKl�5��,5h�խmu�V��X�Ql�E*�Ip f.5(��kJ�j�KJ�ҕ���
J��c*��b�
*�mjT*���֕�hl�kXZ���"��Q8 �U*�
��U*����K	UQkZC	d�Z�)
�-l�M,���J��5HȨ�lhD*Dp c�Pvj�-�� ���(,�iYA��4��� �
m- �QV٣$� n�J�)E� �Y	D#F��P�k0��͵Hր�[j �)T����T�  ��r����C"FR��@Y�%H��l`[+�HQD��TD�  ��4f�T�a�j
�e�h�f��F�a�6�cIf�JR&��ؔ �0��"� -���jRUR2�E2`)4�60-����C,�(�C&�p     &h1RR�	�� M�LOh�JT�����&dB*h��Ԩ� h     �J��� � �c�bdɣ	�bi�L#0	4�Q24i6���56��mF�?Bf���}�<�?g����^8������]�k3�ky��!�iy����s�r�^a��  ����K 5	O� @� k�"/��L� !�A�N���(����?��u����0!�$�@�@���@��C �5��d p���oM�{Q?��������$�u��wɁfq�L�0�X���L�]9Oޠ�O��o%��H������o�����o\qUL5��.��V�Q��i4]d/Uk0c$���������eB!P]Lw�v['����(F<�&�� �UfIPָ��H嬥�'o%�zf�Z�.�nI���V\Nj!"��ف�.՘�(Z��k���dWu���6���^�y2]�t���Ú��
�ERī&^�Yw*�QD�4�[)һ2� �A���iGW!��l������mJY���֩t$,����b�ڻ{{Q����oP���w7^7+p���m!pJ�����1��T���
�I�leD�!N��$�JV��x�6è&:�R�rƊ0��H��Cvu��ܕ��.:Y
��n��!j��T+n�g
�fޤ��[��ͧ1�(`�f�m���Zu1pC� D����YZĖk�Q�P���� r�X�
��Lx�R�##��hX��}�U`�q�H�A��qk
��^�x6%�:u*GlL,�n�H��v��I� \�����$ŵ��4b��%k��Xj�,Ҏ�D,�g"`��P�V����DmnJ�����5��`����ú��UJ���I���Ze�Znޘ�P9�1�2�т���A5�i]���L�г1a�e�7偼 �ݭ�[�hJ�g*��-��ʺ-�.=Z��+("�*�[�}���B�3o5N�L�����1Q�N0���S�G�4V�[kk��2�cʬ����a%�+Ck%�h!���^���'J'�ݒt�eL�Z�Yz�G��eh�-�*E��ǲ#.�xl�*����u���8MKu��wJ��.��yui#w��=�6�y��u�`aF�]1��C/(ۣyx�8��ԫƱh�֯@ݒ&tl�Fa$���U�qT����J��f�֛�4{�	�	T,��,x��])��or�E����Z5���t4�Xk7-��ຘ�c7vļ����0,����lCR]�td!'�Qm�x�kUh�uS0YQ�
?�F�s۽*�׹q�S"P�t2�֠�kįT��r�����Ы�F��F`�]1P��P�V�Q$υ&��'p��wr�P�LȲ����$wt[V̬�-*ǍT�jl���=2�
.�\M��[ZfV�X��WY��!��V*Q#l�_".]���JR�IB�t�F^�k�@f�ӵ��1�XT�����X��I.���x-�T��v�ѫjDa�[u�w;�t:f�Ɉ�oÍ�`c��&w��6��n��2i�`+���ݧ�yKz�*X�˒����W�#&U�O&KV�4ؤNiI����n:s�6R�e�8Ō�#�'�
�3p�!Y��"�Ib��L�P-�c{���UԧB����^l��H9�(�{VȌ2�[�^8
jG#ښ�\i-���Q]1g[�e�y-݅Zo�ki��E�V}3)aa�� ���6�R�u ��qm̥Kr �F�2�N��.]+kFMjZl�r,�K�݌�f���n�rn"��ҏ$p��hV��.��(
����-�T���c��ێ`�n�X3B�x=�CF+Ubd��
�d-C#eA�U3r�a0� A�o781���m��4�2.jOb��Zfa)�Ab�V��d�x[�;(L��i��۫ߛ�Zqmg�(�q�����a����'&kə`�Im��צknZ�z	��㬸�JHTW�ucܻd�V�li�Y�kffS�n�&�C%,�uj���Ӧ�,`�2Ҭ2Xkeb�aL��mf�d�n:y�I�Sqa���RH���CvKG1lI�C����g5��	h�amm�LL���-[zP7�A{���-!�CH�hG�[u�ҵO3UmȱhV*Ƕ���J�T*�M���lq�-j`7E��zƫwm�K����K,5�5�dPZK@����o�w4̾ʐ�Z;�Q���m�:�6��������j'��ݢ_	�/$��;l'inJ�$sc��+D�Y,ڦ�Ԙ���:����+�N��l*W��$+�`J��^�_i����4L�1M�����}��!�3��a�|/^�Ŋ��,*x�z���yn`��M�G�Q��yr��m]d�n\`��WA'Z/��2lloACi
x�@��墯]6j3�&�BTvYcC�1�=7�����0�$�C ON
գ&��tI�7�@@X�]��hӻS"�K�x���l��e8�5P���yd��T��Ch�2<�oU8ow��n�,�*��]=��b�5yB%T�ɉ�짵2D,f��х�����ЧQ]�Y0��6Dԍ�Or䙑oJ7EDtʫ.ܫ21l�r�D!k2!�V�s2�@����g[�I�xt0$z(;�T���bb���c)����Ai7�^^�5�ջ��ˆ��
6,���r�:4LL$��w[EH}�dyl 6�Oqb�Z�z��@A`c�Ш�y��Y*��7vLf��0QQ���Y��5=�EY�.�f�2a�m4��t���H*�C��lnܶ��!A�Kne���5�L��R����h��@�k�W&uE��8[Ǧ�#C.�n�*��@N�f ���G����-,n���(�X��M�N��]�3$��jJR�U�m�gYQ�eemTE'Q"UE���%�ۼ�e��W��Q��
���
Yl��P�h4����N�a����5�1�A|f��,�-�]��V�}*v]l�H�\Ү4(�ӁV��n9Hʵl�[vg��TO2���,2M�+^"X��:4b�qe^�X«.K/�ù$pÌk7��(�v)��H�N,�Z�\Sߞ��%�v�h�1t����[X�#�ˣVw�
4,C1L�bka�6�p��{��M�mփ�p�NI�R�mG�m�,K�.�׈�I<���[��$(){b�y3c��+�>�R�YK	7)��f��#�2.l`�Cwr<�T��&0�ɹY2|��/�X��M.���Z�j�� �b͸�]l*MwI�wv�e�̀	y�,Q]6��BՏ��/eAt�t�U��K3PXѶ���E����LST<Ͷ&��V<k4s������g-�؆*X/Z����ڵ,�%
ݨB@b�n�G��sp)qF���X��i泉��lskQ�&������f�X��F�A�pHr��a�E2�F�0C�гw6��(�B�K/%�ɄT��]��xB`SP]f՘v6,Rʏ7c����Ѡ��j҂9/�mD�\���C�tc�h�;_`ux�[JȘ��]�gi��P�E-�7���va�����#)B*hf��Lzkahk���8h��F��V��Q{֛�����řsA��ޢ��@��Sm��#+#-�֦�YWFJw�偨<I�E�K��P�pǪݟ����#�]B�ѻ0��t܁�E5J)F�>�Ăq+�j����Z�P���ibN���CĲ��{[�K$Z��6i܏A{�(sQ�Ne�|���nd�c
W��{�cXlF���ߑm��i�W�v���Y2��d ��0���-ꖳuH��pZ s�nмfȨ��'��˰g���k3u�w���E�Z�-r�F����Y�5��b�sZ�we�k$-D�\��TqVU�G!�70���[���"c���TJT�/v���Ԕ�b�X�J����u�f-/q���ͱ�,!5��c�x���{krXt�-�Rת�¤�WN��Z�7�رz����MP"'"��!���� j#t���8��3��Z�\5dp�;`[x0��B8�2���ʚ����*ʱX���Y)�6E	H�l�@mE�h���!�ʖ���ye���J�����_Z�
�4�d�h�V�U�Fq��5/!ץ�先)@��#�*�4��%^�����[7*i�·�t
Ch�M����i4۴��#u��\̈kJ��u�^2���m���UWl�> ��ݷ`�J�s[�wsB���h0� 걨l.�[�	��S*�uF2��Cw5!MT�VQ�r��C�л�/ۗI� ���%��2�u�t̖�t|6Ƨ,�f�y5�mdF*ض����5�[��Z�e@2��u[�{�8��XEE]�^;�i����DMU��9#s,f�5����l��� ��憨���]��-+�T�ˡj�Y7R�SVU�޶�1�]�Ym�B
���
R��t�`ҭb3wrG�-ޫL\��7x��Y��2�aX���R�b��"�0̤�cehZl�f�rS�PY,�[Y�o(����i&��sp�N�U�������Q͖����Wt��fZp��,�yB�XV�!�Q�/v�)}��mj�R�AJW��b����٬k�cX�@�����٪߰�R�1f!m����Ҽ��� 5M�J�;��
ɴ>��ܚ>���//-�]�R�k@�#����n "9��$ŌZ��B���!!%�C6)nĈX�JzF�jh�BF1�5��&�EZ-Z�`+d)�dTXA�[olnVd�V� *Y:퉲��aR2!՘[V���ɣ1�Co��w�u�h����!��]�!V}�����N����l:���7�}!����ҳ�|��&� ��>�>G�����'6��.z�3�txt^7��z��yWu$�N�.�2LK&9]ݠ��_A�Acq�1�xD2��(��w]77���-�U:�΁����;�wg@�l����ǥ�v�^5]қ4s����u|/��������5�����Z6G]�_H�>�o<�X�>�Q��/!�RW��]st��R��rE���yǃ��չ;�Z�q0f.)�S���>O����ug���8"��_	�ͫd1(fs�q0z\�HNvEg����&�q�
ֶ�n���!��N��5Ō�%
�s6�\e��b]�W-zy����R�!���E��Y�W���^���"y�μ�-�<��]�}i)Ci	��W:���B�Wi�:�Њ&����L:�3j��9�V\<�Z<!�g�SU��{͎��F0����i1܌��Ú����[��e��N�)��&%'q6�=��D�|k��p�=G�� �Kf},򿃔k��sj��Tܣ7@u�˾��:�Q�ov.Z%*���!�	u���uj�'YQ�C5n����k#�-��%5m	��;B���.5 ��+{U�]GBLvD��<�X:�yrl�@:��H�R�=��r��X�q��A�Ct��쵚[;��9�0��:��,�j��J���T��3��M��v^
����f�ٖ�*�o_+�gnZ�J����/�@z��ȲXuz�]�*^�>����5�m�8p$����v4�UǮթ�;�	e"c�Fgo=Τ��� �*:� .G���f��k���|2ni���^QIm�ӂ���$tu7�]���v�5���&��l�RI���϶�����
3��Ԙ�jKg�j���(Z��Z6��7Hq�@Ӌj�gd9��X��5%	<�����I��V�:@���N��[[bb���6��E컭�JT�A/Cѻ3x�hV*�n
�bvO���V"\+�J�y%:B%��2�s��*�u8�ۂ����Ap�����Һ��N1X]��r��X�g�zt�9>bVgh}�;��"�g7�q�Ճ4�	�t�&�V�J�\(Qd�*[��QJ�r�t�K�Ƌ���w-�GCٔ�F��T�U��S�h7��f_� =�m�3ǫSnP�����G1>h��:����='��ܙ��4��{�B9py���L@hBݢ���ؑ3>U��𨯅��'#�䏄�E�*W��� �&���Z���B��,-׹I�ﻔ��Q#W ��Y-���`�� �%�aFR����b�s�=�F2�%��I���s,r�\x�;����Q ^Ȯ9�es��H���DF�ac�4թ.X�R�0�a/�v��Yӻ�m�e�V������� D�����Gtz���k��Sϸܧh��7c�}�ۚ�t]:�{"JmA/���$�.ׅ��3���׆�YE�v+y�6�bfwd�gN�����5$$aJ����$�'������:ʽG%]M�k�'m�\��̻Λ4���ӭ�:����au,�'�U��0�O{�\l�S�����*���#CQ�N�6�M:��Ic���ްŚ�2�N��k���ȼIr�\�T��nn��.���>xL]�L�e޶�Z��^�҂�Ƭ���yO�si�2��;�>�J7i`m�/tu%.��hC����D�F�I(}3���6D����1Rw�\�4���V�/d���7���Q�d%u���s_J�O����ۛ����;�^tPX��@�	c82��/gnWl��]���$N�Xy��퐢��me�s��K�E��m�鴰}�ukXh-�[v��ZVe�fM�\}Ky+�t�&U�,��]��ʲ5]K�8��ks�5&��8�2�,��g�k󱦗p��۾Wʉ���%r���y�:�¶m��f�޾=ۅ���P���NH`]Q˶�$1Q.�(Xǔ^e�Y��+C�t����[՚q���m]��h�[��|��ǃb���L�5�Wq�01��%m��7V��W5:������L,�v����Ԡ��]�����3� ���:�;r��k[՜��o.�4����ϊ�xq5��G_q��sF� ��ՙ9P\��:��膗+�v��:���2��� ;X�s
ǐ��(��Zmu!4��
-7&�*�&�o�[��Э����EJ�AY�u��|�cǸ��LUtS���S붖U��0��X��1Zc�v��B]ئ��9ۜ����!z���@y�˧�|	݋��>�ؕL`���~�t�Uc&M���8��ʝ1���n���,8g��w¯��;y�M߻�g�)���B�X:�;ܾjö��3C/xb��<��^���ΆK6w�y��|���1^e��1޷��%F�>������-�x%� �Ԫ�,��]�;Ru^u���F9��G��w1/hRٝa�W�4�ɦN��J"��f�6��Ʊ�����TyE���b�i����wQ�E�/1ڹ)]|b��ۨ���tBg7�/1�����ǩ�[+=�
��*R��m��"r��ow*�Ls��
����مmnG9]M0U�9�R�u�㶸��S�L�ΩW&�֞u֕W��\q� �4���n���F3.NDm���갇V*�L�:J�����I�d.�W��6�b���������d��ec�w賂��E���Mt��d޶��=\�
�uD��';L��j���,�P>&��$l�kk�|�ȳGGo,����>��6��+�7u}�{nJ����yW2m�xF��Ӎ���F���7}H�,������As�\T��)x/��k%��;s[�hr�o0��q��|�{ڦ,�w�s�oY�#��ǅsY3�Z�v�3��+α����j���Ի��<��J�k��O@<���m�=�����b;�0_	)��*f�Mh��-��*�&c�Yv��G���؇��=��в�r�����w5[x틭�C�S�OF��7+�wb��vn^�v�4%��p��3�x�J�h��n���҃j}܌I�I�(�JaIw<�gܫ��Cë�s�q��F�u�����D��lѫ���h|�N���8�H�vVŤVT��Lyvm��0�]��7���w�����릱��T�M�]�yth��l��2��:�uq��P!OnTU�f^�Pk�̾�.�ژ��%h��u����c]FƇ��eW^�!����*�T�Wk�Y�*����ͳJ?��/^�fY�Y���5b�U����K�#(|%#�+i��^%5w]!oyA�.5����kk�E�H�b���sZY�Etv��a}�b�<��=҄m�}2�7�g5)��7������q=op
�����K�]Ղ��&���^>HT�pU�|���u�t�����Kʼ5�S�~��+��S��x����.x�go�YU��2��4���3�swcd:��)b��m��i�dju�O��۽�]����x����}���U}LN��
��Xz��h��]1(�UغВ	H��*��ـ#D�ے�l7Ne���i�JT����c�+�̅|���;�Y��u����!�-u��2҅�l��t߳5AA> P�7�L�P\�n�	����hv�_iv�� ��O�P�����[A=4����VP�Y�qWm�|�?-�W�_bN�	P٫�F�ؘ�,�ԠõŞ�Ӊ �YՂ��cAk)Wgg�
��[�(��4�鹪h�H�z�t�������f���WR1;��Ӌ���ΜMa�ݔK=ڸ�q�c�hn�.f��X0T�I��6�3b*�@��s�ʸ�AS��Vك���j��Jp�96�[�[��ᴻk���8>91_X�AyiR��V�ۮL'�
�<��9b�f�)o-<�P:l�]�ˮ��u�R��ڥh�u�"W`!r�N΁Li8�(�5{u�J�M�}Dn"�)cm��s�R��1f"&N*]���5
г�:H.]\�um���껮ŷ��r��,��vc�6Q.���u�bR�pI`�B�TL�}X�u�a�6�*O.��gt��n�f���Ƹ6o���ۻu�v$Bb�:����,�A@ �XlY�b)���.���82eY�ڶ�U�dޜ6B񦲷.���|�_uMQ��fgS�+��/�[O��w&���lu��63��o
m4��z|{|:�i-���Eb�R�	>y.�v�o���"�Pev�h���m�5 �R���|��fK�j�V���b���}��w�M��.�2�yf�������+�ʸ��V]"�X�Oe�	܎��d�Ϥ݂KC�3�t�:�8�!�2v&6�\��6��T����}�巗�+b�53j����4�)��i�C��w�[�8�v�#����-�3�3�]z��Yo1�����"KчCe��v�gN��q��Y�Պu���ف��Gq���V#�چ��A���H�30���v��mn>��g>yyP��EB��vp�Ԭ�a�5&���������mE���'�e����n#��v2���9��K��AB�q��)"��(V����{�8�^�s�1:PՋŇ
.I�%��g.l�,�o]����fwP⻥ŝ�.`oL�>\��K�4���wI)B$�I)A$�ITm"Km�4`� ��  -Y4�$�#iǜ��c�G�� >�7��a><w�@�d;�	ZR���RI$�C��gf���?HO����fR
�э����*��ren6�1/� �DP���n�hi��c ��9��t�HTc8����PǗ�խ{97qL�$�<r``c���S���)[���Gbr�\;&>��E��9�
�N�,[]ԋ�;VX�[>�8fK~��>�o�L��͗����K�gY
k낤��q�M������S��Y;F�3U��;	�%Yd��X�f�s�`�.�e�A��53(Z�i,�p�Zc,�l��Y�5c#��E�G73�����른w��W8*��镨��6�e�0��U�"++����a��� φ)V)I�o�Ҩ�?5��S�����Zy����l̃F�i���!�ә��}����F�1W˹���ѻ���*OpI�x����7��A�(���k��,\��NM�S6JGrU�:�-�=p��8���N��׮aλ�h6���#���Y��x��Z��C���,I�7�z�:�g]P�R�vm�m���^3�P��O���`ϲ�'�MogZ.苜op	��Jd�H�uڢ��_��g��Wu�U�܊�7���r��۹'�PyyPU8�+��wbm=�;�r�$ͤXa4�N�C��'XxV^�$Ô趶>̣�Cv����ܠ1S�9iL䤀E)k]+� ����92q%t(f����$tn)�vN�j4.
�w__)9Ǚ��q)�:�,"���"Wc�n�%�L��(#��%	{/�_0��u���/�h�H!�;����H+ʏ���i��l�i��]�n��4�w`l�2�r�[+�a�0B�n���t4&>VS�(����)5-�`�pRMb��I�Glhd����cn��_#r����Tw�+�h�t�l�e�����ō\�u��`�K��#[������h�d�upeJӥs�f�;k�Di7y}�(*�1�i����F�k��X���cL5����3����;WZ����y�aZa�J[�7c;�TFލ=�
��ʀ>���p�x�t��N'i@�U��P��1� =��ehyu`�D�D��N<74��!�Y�Z���39�zD��Q���}y���>2�-̰S��O�`ꕗrö��nSN�������f�*��q�(mv�s��Y\LE�T��:�PѓhSH4Z걕6�mp2n'+���p��v�Y`-OTN��\sU�ܒ�F#��7Y9��X��5���%�2j��NWwg`|+e8wW��;kzf\�fet/���hp�ibg1Y�C;������v�fV�0�:�*����B�e馗A�Wvq�8�d�k6�:#]�]͞�H3z��9��)nb�ۗVk&8���:��&��Z�J�6�l��γ�NZ3uI�J�g]s�[Zm��i*t�"��f�s:�M����(�#��x��X<4d�4��l���p�%oe9A�3�b���n�.�w1P+���'Eb�jnt���� ގp���Ť��kT��뇵�*��/wefm-YEX����� �8U�N��֢��ňs���L�YD�RVu_R�'�L&�b�e�سo�!�̰��8T)�q��.���S{kx \��_�������#x�8c�6�M�+]��ġ2��{p�ь
�Y�s�yڢ�^Z�N�Iq��+��	d׭b+���,�)K�
��KRcS#F�[�Zya���&ML�=ͫ�Vx��y
E��=�(1�
��2���ː$���@��T�1�����Ri�ӒԷ�W��ʝ��ΒN���xQ}��6**�o�jI�|�i����P�z2��a���YM���q������2L����+���ѱݘ�r�[�t��E� q������Q��y4=���rF�t�O]�C��"#$uh$��O&"�
l�N⋡cp��ott��k^M�˼B>��i�@"x���x���J��|���5�7����<�a� ���Nm^̣٩�\�\/���s&	��v��us��͵�����/��A��#���˷�̽g��o��/���ה̵������J�lom����`�P�V��7�������`�P��'���)���������Ǹ-|�V�2��M�l֞���=��N���E�'�Z�۾Y�x���9p�Q^G�n"��v �mFڥ/��Y���t)�O��.X�Eݔ0�E'!�@$�`�Cy��H 3y2)r*�[mG�'a�]Z�� ֜�~���N5����}�GQ�}��X��w��=�bǻt
��|�p�+i�^��rd����E�m�%t,Ц0n�1cT9Y� X�r��,�{��]�H�PΜ�<B��j޹qm�t�L���Sj( v����q��ǩ3|ʈurn�{��iW+ܕ�Pݩ�i��Vu*:�����yV,@��4֎B�S�e�� j⚦2�Q�����=M-��FXT:�VsǗQu�B�`�N�7��p5/3�Ĺ��Jxz�]M�RB����VR4E�r����Tf��V.X�uJF���m��		����ԚFh�`G*5a�@�Qո����o�]Y�TPՎm`+�n�wbj�;�U��!�J��4S�y�$�\v���d�>�%U�*aI7i
�F
�\��DԛA�9�ȯ	�ōx� n,n����Xw��^V��Ց��ԯ�]�M�_,3�^��}���Rx&�]�m�^���T�b��%mGM���̢�w:�R%��s�($����-�P9Z��.I���h�f��aKEv���J>���M@����]����X+��u���$�u�x�]bƇ6I�2��`t��al��O'5QB���K�X�����v��q%Zne�6�u/7�0�c��[��{*�::pd(�l�cQ��6*�^q�A�3�5�e�2��ml-拺�:]�IMYN�%�� �c9uq���žL�X�ofJ{¯��#�{����©p��>����:�ъ���3�EB�9�]�A��� TNF�f�o��Im���b˘�ޅĵK(w+�*��G��΀,<����7��˗C%9wr�Zsw�R��n����ւ���2�@��^�"T���S7�Y賹�遊�zEJ��l�R�~��@�0]�ד�B(����5��F��JȢ��&�7Wi�k�5f�s��9�\�s�.��f�r)�������7I݌Ǹ�!wZ����m��t�Փ��]�n��;N�3�9\Xtp݀�%@�O ΩPSTV�Uc�w��]�@vb����n�I^�E"�L>,��ᑆ��즥*�O�Z��+WR��4�ø\�"�R��7�ه0];�39s�&���i��C�w2�R��%����$U.�u�q>2**���B�0;J[�����M֌\�3M�T�H!O�9F�{r`s���s+�vv4!\�=�)��|/�L�쭋M��w�'��h\J��Gj۱�7�Y��:� ��U��49���fƵ��&����顓�h�+�|��t�s�vv��;����+AՙWH.�-K�Ѣ��w��:�E�K��"�:��o)�,b
�i�XH}�˪+���3w^Z�MI2�������Q�I�VX��x�7)�t�^�PLz�g�_w/�gYu��s�%�6���wC֨h{7�e������5��AӔ	5���� {]��m�₝^*B�@@�K��p[&�Ux�@�Q���6�a�ֳ�$̪��n��4s�\"<ƜCT������rw�u&�-�eQ���Vw0��uV(馈:��ΫǗ���1�W;��dCi��H�qB��	�*�%"�\jn�zP�Hr�M�g�����Z������c�[���,iɊ�v�%d�ݔ�J�!*�a��S
2���ڤ��t�o<4��iv�w����֔ �ht���	]dބ]��;�/K�:%�����@�Je>��-�����t�i�m�N�a�+��)_S��.V�݀ԩj��2�i5j�u�#@Z�X70�w�(U#����s7n��|�ڮ�T*�ξH7gMv�=�/)ET�y7�,96:�G�!X�J���9&Uy���=��\c#L���R����eYԣm�����}�xSa�eΣX3���˭F����x�`ɗVa�.�;fK@�QҳW2�R�S�`�
��
�����U�*u��S�_ˉ�b���J��*l��཮Xo'v��$�L��*�*��:��T��hF6��fL�0�Gf,�T�	^�'z�)ëgV`�K�:{��X]�cTo�(o@�U׶n.���Xt���Y����^N^k;�4Wۙ����Sn�n��A�c�gQ�07%�1+�񼂵�,Zj�`�L�G�t6�T����MH�j�h���"ߤ���L��Ɯ���sV��kQ0G�ػ�VA�d��w]c,b��g3P5p������n������{J��[��m1Ho[@u���ܬW`L��B�i��'3za��Mu+y�%9Lg�P��>n��c�Tgr��]�U΀mս�Kz���n��L�1��$�,'�跒fif�k�G]mj�Z���v"]��]۫N��>,���[6�C��-N��oj|PXu�}�+�`�@ծH���qf�8V��{��(F��c�.����( ��IM�c��b�4U W�3TW�]�����DG��@ �(E�p<	�`���|:;2�4>�R5:����;?P�>j�t��!��c��ί�����ݜ�nR�a���c&�9Q�A|�"CR���5z�8U0{�ʁ������5�QК
+�J�T��1���#��&DI�V&M�e�6٤6I;.ص;t����,�Ye�j� kN������m�pGJyt"@�T5b�>�����+�fN�U��}�]ΡY��[��Z�8يm�z�����#�-n�xUqwغ�5Rm*n��v�p��h��6�Q�Ɖ��=LG�o��Z�ӋK�
�&�9�;�w��I��qH\X�������|;{�!��|�gk!I4	Fe�E�H.�e�
�²5y��%C�v�e=㒜��	Jo������^�AUұo��b�/�g(p��2���ꎍ+�yu]*
�A�x�Y��?�.���	���ڳB�*���3����ه���3j[(�[�sF���5��8N��f�do���鼺�������jWI�b����98�BS;'����D�������L*=�R,A��Q���*���1��V�j�E��E��+\Ah�c�*("��NR�H��p3(()ǅ��ĕYZ��h�b�Kjʕ�R�VAb�ưQ�&!P��V�V,Ī�5U�eC�0MU$uk1PX.!X�0�˦��\��f"*1Z��*2*���V�`�ZZ��P�l��`)-�V��0�FE[1���,�����1�s2V�UQ��j�5]["�6�8�,c�l�
AF[H��aY1&Z����EZ���X�bE*���6�q�mB��
�(\��w��>�����������[�C�v�b��k8�v�`<-[�]B�c;P[�3Z<{>�����w�~�mҋ����+�K/;�m�����R�Y]�#��>��ȫ�����Z�S�i�����g�ʢ�fo��[S��J�:㺚G�&_f�k:v2�����feP7���>2�*y�d!������G҂����U,�U5��������u��.����������0=1�U��zٞ�׶2��=3o�R����ǻ�.��>���}�����ԏ�=g�w�S�|��k*,E�*dН�R�ϵ�t�P A�i� ��͹|<�g�`t�����v��JtbD��g����0��U�[��gOmN9�%ꥅױ�����b����׃��[C������Q�ƈ_q���m.x��8 "�V|��zW루7�f���R��\�*�k�e���6�r��\x���N�$<��gP]9���|�Qc�z{���[�c��P I9���EX�����YW����-���̋�X)�U���U��8VZj-(�s;:<�"gٚV�j(7�.���0Ut���3�ZG�:1��<�;l�m�I�W[>~S��
P�A�?�h����s�[ʰp���yO��ɛ���֜�O�P4�z��
��x*�_b��p��=�����=�X��k���Xْ�I�t��nc�;>ގ3]Ul�cӝ�����A�ֳ�ƍ>�b�R]A}o�Q|��[��eA��[�q�44+���>���q���Sክh��q�9�ށ�Fz�����0�yΔ��~�W5�׍m/�`5��ƽ�qJ�U�����%ɺ�8{d6�F�Q=�^6���I���g/YM'Y�P+e�;�)�V%�3�N�c���]EӁ��c�O{j=����Hs�YY�������3�7�d0�T�[���xwN�Yj��y����� �wҴM��ei��v)��t5��]h�N�T��Əv��I�w^5C�k,��!����S��XB1�s�07ꗽ��e�-�qU][*xh��"tR�h
Y�K�^�[���r3�����.�;f�s�NM�{��D�TJxL5�ϟ~�������ݪ�c]A����F���_x�U�g}(1)/.]�4ne�ߒ�u]u�u[B���mxcإ}���l�i���7�:!��@�۷b;\,`��]����5`���[���ޑm�F�)V�f��)g�`�����}����h~~8���z-hz���`�����W����Z�6��~/ʠ�3�D��w��WU�����6-�/U�ϼV�ȕAYV�U���~#��d�'��$���v84)��K������l���>�˯p�n{�Ow���*Z(g-��O%	���Z�']��m�4pl�'VZ�I�C��iN�x#K.��7]O]iE�8K���i%�nU�wB�uF^��&ΥK�]/�Ԛ��v�]r�u�X�ueqp֯��8��SN�"nW:����,�-XQ9.7��F#�L����9��P���r�����,c�@��<_mʇ��Q2v��DZ|���]��j��}�E�i[�Ȍ�z&�gS[����Z��hC��.ˤii8k���5cbpF�[۹������K_QX��݇x��!���O^���<����n�C��f�c���P�5��/���9���V��=����V*�`��i60��3^��Hդ<*��;rC#^����
2�Έ��R�9���$���rC�0�WuW<��v�JTRq��}c�#Lze*����b��_t�!�0q|��c[��2
�C�8֬U���p����;ΰu��_Vg�#4^����n;B�&E�Nׯ��*w{`������U�ٰ�(�Q�Wh�Yk8sr�VGt����3\�Uֳ�����6�ɷv��V^8�>�y�!S�"�˕=3;0H0*�Rcb�.U�׹�b}�%��=1�L���T��ZU��E����pX��W��
�ɸ��Z�h�(.�b�(���f��/���֮]+��O+�5|�O,��'s;*���n�˗�u1�.ϢyF��I��=]I��5�~G�V0� m_�C:|
o���BY�s�|=���Z8_l��v�˯�0�Um�u�g�u^S�`���+5��X�5_��E�g��q���9y��Rf�R�tX�.���������h�y�&ur+E�|=��[n���s�2�ʫ�i0X�VĪ���I =O��َU�NU��x�ɅPȂ�LFJ�XV;��7�'_��7�n$V���������Ձ����
��;�-��������/+gѥ����h���eyk \�GA�
��I�Y�IB��m'�_1�ϥ"xKwK�,*��c���Ը���}Sct�X�_�CA'����ִ�xU�C��TQh��&.����ĺ�9�{=itu��]��L�oݗ�G�
�.��^��;Awڀ�z��Ysѩ�l��.���\��:���7$L3�쬯��]�����'ȷgC��Jo̮sO���k�u����*�L\FVJ7��M>ɫQl�gSb�!�B�W�K5��D��ưk��(�y���d��Y˓�w���w�WZ�2����ݞ��&v����ϋ�Q���K=�Z<k�,�Yc2��
�� �w�Y�4"!h��}}ǎ�I�d��#���E/Y��ӊ�_
��~U�V3vf�P�h�akLs�T�R�����@�B����k=���f�G�As'���["�
�
W�˖�K��wZOP�]���Z0�[�揃t͐E������څ3éb��V/�Cs\W���]Ǣۆ��ݗ51a"��;.��fh�Q	&0W<�r�ʾ��������U=�VBM�C�RˣXY<�iu��\�\�>��Pu�[���b�گE��rcTuF�#��.��E;��Ƹp�ʾu8����>Ն�Es ������h�reK�P�O�S�����X������	�󬶺��:��۷���(~�����t�L����������=ʹ���;���)Ô<�f^?eY��U�N_!ai�ß!}�ҷ.�����i�3]J_���B�d��ʠ��������+8���κ-�|�MQ(ӃP�n�J��IU���E�c����ݛ�pg��+z���Uu�z���
�������x��]r�n�:<95!�69ݾ��
(uYb���N�Xc�����X�i���]�(��S��h��yT���*!�/�Q�9��u��SsA����C�VP�;z��w������}�{.�%j�#���a\���a]�I��U{��x��?aw��L쾢��G�'�"����#�1y5.IOh�8����f�Ű�Ho��ڬ�C�o�[=�`��NN~�{ݛ�Т��c�ß��_���B�m�Qب�r֚����,2�=�?!]�È�3����W�g��W�T���%]dP��S����ӱm+���u�_�������rgs�B�8cH�6�w=�>�{c�������g�_�9
Bb�9~c�k�')������<��r_��Zۧ=7�)�c��.pF������׍V�5d��|���F
�yp�ol"71�z����k��Y��R�w�;fj mT���$���cd�XIr*����Z��k�4�`�0 �^�5u#eCBU9�'���q5��p��Ƙ�GP�5��|��	�Ƌ>��κ���2�IK`�
;+�,�/c޴-JՑA)X7]lMm��,�o.b�fJ�i,Hd]��<{6���ŚS�Xl��ˬI���"+^�Tb켸�l�}ܻ	=Qsf��u�M9"�܈(-o��ou�A��/��X�����La��f�
&4�5i1�S+^�3��=��kp�G�Fu�Q@B������:jetׯ��_N��vqv7�uHQ|
��5�u��`܋�<UG�O<;N�&����ἅ�,�,AD|I�5�kY����'yV�}4��8�̹��]ȅXx(h�xc������Z)��@ӱ'����=��	@՚�f��1����z�\�Hf|pX���8t<z�Wu-�O]T�e5^r�q�9^M�S�f6hi��W��(D��5a�*��0*��4/��v}�b-x�!{�߷��s��3X��D�����2~�/H�*f�82�ϗVP��F`����EȮ��n��Ӣ)ں����>����>S��#$���}���#+���$Y�;!vc��δ�=�zV^��Pưo2�7Ɂ��2�:ǃ�r�h����\�Lt���e:��!J�&aOS�F�3ƙJ�T��Ů2{3ܥ�c��ȫáᓓ�U*�Z���J�ʉbi'��];�>�����1κ"�J��甝GD�D�
`@~��ƸA�R6&�=t��*6<)U��e��Ӊ��h
q�r�
4�֞�
_a���:V*���g(<0P�%	��n�s(mA�M՚�7��Q��t�����k�v�C��ޏp�>���B��S��f�;|(1�>�Mm�.c��SR��D�W{9:��J�$њ���F��
��`��E�Z�!¯ZԐ�2�����n���ר*�Z��
�����*M(������kp�%jn\7�2���Q{J& �xg]yަYޱ�w���S��T?�~d�����8�d�?FR;q0G.L�E�U���E��RΝ�I�F����U;�O���듥��v�}��o*�ZEܬ��Z���9�Vum�9�D�B��R'6d��K����t�J�;3Fjr���`��m�ab����Rp;��H�ig9\1�;�.lZ��.3u(uc�n�
<����E}S]�l��m2�=�z(j}�n�t}�$��ƖnYE�ƪ�&c`n���v�	vd�6J'��ǳ�vT�.��;�GoS��X �6ٴ[���ƻ������ت9�L�5j�ͅ�X��d��]�(P���G�q`ft�b�������hRbr�:Z	[WF��c�7�/�����x4:V�~{��q
��m�H�T�+���ԭ�NZ6`l�=j��2!��-l��VU���\��:�vjk���)9����B�r�N7���K��b�tE}t�'N=SU�˭�VS�����n*7��j;�*���v�����!�x�p�
mR���z�R����d��U��3�g�s�[e��9c��̽�/�Gw�Ŀ�n*��! öVBQ�"�"ėi'\�gc���j���u��Ř�$; �O�;�᫺��Ъi3c��c	@Y�V�C�|��ه"��˙k��#uئʕ�VP�&��$z]\��iJ��ƥ�p-;W��v�Nϳu
-P'Ae黔)��u��ՕZw.�2v� e[�g�����0Az&��n�S�޾x̠fȮ��> ]J�1�,v�7\8𔴠�����iQ��]��v�j��7j[;�+��Ӆ����S�;�s���/tǮ�Ը��S�`��ggI�f��n����ۢ���7�s��M�C9Ҏ|��v7%�]I-�j�-��Y���<�C�仢��|m�E�YK����_v���[�<%���$�*��@��x�����׎>�bb"|�����cb��)dm�*[V�7)L
 �DE%�b��$U�
c��Kh)�j�U�+��X��X
E��Ơ�P�fJ�YQ`VV�"�6�fJZ���d�"1DV�yj*)�Tt�Y�����.Z�m�Q& 6���������,��bTb*"��$�2��b�E���+�b[V,U�nd*���j�qi*L�Ub�6�GX�fY�Ŋ*��P�r�`�Ƣ���`��Ҭb��m"��A&%�����*R���-�"��c�&�����/$��w�tɤ��ioE�GN�ĩCiV���Z`�^�?�t4q��������n�Mϭ"��8�:�ߐwN��o�>���eS���	}��T��W'peP��PhL�Xف���g�w�3u5���q���vaCME§.n� �����YyD���ﾾ���P}��{����|`�_��l;�B��T!�MF*3�9 (��	�q�x{y�ߴ̯|�x;w뒞|+����w�nR� �e�S��RoI/T��ǂ�신���� �]^�V
��P�7g�������T���/pT���+s�u��c�3��~�u=�J5�o%��kM^R��^�{�N���Ǩ��\/��X����߽�in�T�ދh1[��ה-R$q�j�)ʪƢ����fy��]�����
��Y�֍��2�ʉiY��?-Z;�˫Mtt1�D�t��V�G۾[�Y��%gS�e��Y�Ӆ;?p��C�kv�z*�2�򷷥��3�m�0�a_vХ�8��q�}��X�6����_�Z��˺u来kP���a��Z��t�#�h�5��#������kw9 1�@����i՝��Ui���������8<��������m����جy�s8C���D��2�"�Wg����ۓ�/~�j�G���kÛVZ𱂨J�[e�K����o�������>�MxR��4��[��c�k퀡��6������q�g�1Sŉ�p���O*R���]F�`\����a��x�]^g���Q�_,��~<01b���`���g`���[/�i���jPU�Q����P2�ѝ�V�t5�V7�@���Z�gF�*�/���Y�\�
��X�s٪uC^�Oz.V�u�@�40:��p���X4Z<<<,e�W
��س'���*����"`��mK g��|�w|������-wǚQ"*i�]��z�(U/��T������Sc�Nk˷�E��nyFkWy[�q��k�Ѹ��ؚ]:,|�%��Ŏ�5R��R%��k����ht*�˭=�[��VI�/ڇMƠ�F�R#ǇPxk_*i,QҾX�.��z�^���qT����p<�;}7]����Q؁���Ȫ��8�e� L*ebe�7LT`��j����0%K�R�x�v��������S7=��*<@A�^�x}>�)���~��W�����"w8��8=��ëq���8)U�4ad��U�^�+�@`��
�O �ԭ��:���t@�un}�����u����٭�R�yT�%�EI���-�1p�t����U�n�V�
����
w�pM���9ݛ�@�-�	Ӡ�Lh|xc$`�iX� ���cWc:��ܩ��h+5�q��i�XkA 3�Z-���c��+����n����9�K���R����h��ݢ��3��7�@�^�c�f�;��3�����"G��ߒ����)$sJ��	�
�Ѱ޻����Nr����!qu����+��M!R&?C��[*fc%��:F��r=iN���٫��T�PkJm��f�VK6l!=u�]GL2]]>����xUC^:���w����y���}��(�2���u������X��y1��[��s|+�̨7.���k�Yf*:�JN�OW@�Q#*���0M3�|y��B��3^�Ar�p��Ep��ò�J��u*U�%vҝ�:�����J�C�*���+k�\��Gu��o_J��z��wd�ǑP�~J�]&tVxϙR�k��FL(�dA:aZ��t�J�foq�b�)�	u��iV��
uh9������,'�3���{���T=C윴V�e
���*���0�0{��/+�����S�|%eK����H����î�Tb��/Yܺ4�j�*7qhQ�cg�|����-v�:��n�r7Q�gvq&l2��$���׈��ך�68?w���T�Mvev |��테 ����lC����q ���	2E���&�v/�舅�s�n2�~����>�яU,/�|2�2P��S��9HԴ��6���Ψq" �EVy��u�5�l�*�8�6e�c���r�r�D�����r."D��P�/�֬�F��~5�X5/�,]�1�~1�;V�V�W
R�u
T+x��g���s@./�T[3=�d~~���i��[��X)T?1+�F���T�k��l޴^Q8u�OLWq�2!��R]f3[Lةs��WG.�+X�����B��`a���cE���u�X5��l�h�}�
5�vw'��I�C�*�s�P��I�ٷ[&L�0'��L9Z���ZU�]Ny덚uӽNM���,ջ˜:��x�YXk�O{�UO�j�oF�c�|��^+2�](���yX*��E���o�ow�J�1�ʋh'~�#Ϋһ���uE��G�
���{�}tW������c~�k�,���]��^N"�bjD�5��tٽ7��NuC��i���<���}2e��D(�T)���pT9s��n�LZ��=J]������83��S�^u��	��S��F�R�6T����m�9��6�z\@":mӘwH���q��h��Tv�N�C
�)��IYRz�<=s^�/.�j�Mo��|8l��Co>����?�yk�{������ki1�U��5�hd��@��o*������6@�N�Yi#R�D�Q{S$`���oXQ7�#�GJTg��aU.v�t�w|���8�7[.n����]��]P�+4(��T�a޲U$7*�]�6�Ъ��b��d[���¸�0`���%��b��W;�9[SҲ��:���W�p�����a��1����YLvi��ݼ��6�Y���W$R���;��p��:5~��c��,�˭���Qʨ.�U�״n�����s�T��W�*L ��F�9��ŷ��n�U�����Ͳ �����f��s�\>]yw�r�����6��éwwyt�m�u������o'�5[�U����_�d+\:��ݏ	t����K�{�P����U��4���t�go)�Jh�J�DK�F\����;��'�u�C���6���Us���:�C��F���C�m�f�՗V�j��S�1�ȉ��:)N:s�%�ɭ��>�PGY���r�:����4�㒚��8>M&�IJ�%dd�����:tӘ9P�̹V���g� @�Ѓ��
�{\�x��n�\�����~#��)@�zòNj�+��/{�tw��a�t�b����=p%u9��N$��;���dp^�o/(��Tx#��������!�ZG���Fno^�v�u�|0S�<"�CA�B���w
���;9� !Is��AM�#�L�7�K��1�PH��5_b���jy)� c^���Y��[���
ሼ"_�OU��{����6�nfm&&��m�"��(�U�Nyz�}�U�m	��������%��~�w��ЅP:�Z����51r]�k��=t�y�LOR�=�F�H�mT W������L|l���k8+lܩY~���dm�׼�b���bkj���x�4�+ɍ��d��ثvr]�s�a��u�P��Q;1ʶ;9�:�K�2Z"��MRfz��~}��xg�+(�U��X�D�,���4��Lh��)��[��ν�e1k��4�VS0/�x`�<���)h{�&7V���LF*�JwX�؃B��*�$z�C���ў�%�Օ�v���O3Z/��p�go甠Q�����X*��
���~1?{Mu�Ҿb����[�X�.[��ꃯ�
 
��}���}��g�Ɠ�����\���mҡì�Ƴܪ�S�Vl��ŭ7�A�7 c� q
kF��1��� S���6�x0�͠{����R?����~Y[�|�Q��"��V�[�\�J}��}���Q��{���#�T`� �#���*gg:W��:���Q0��=�dfrd>�	ծ�X�#ʬLy�U�,xT�^��[-e������5W��Hn]��'�b7[z+h��ÅH��ut8p��#*#.�
�H\u�ޓ��
d�C�&�ז���DG�
�#���W�Nd��}����`k(h��K�%��U	B���zC=���B����kt�5�ѣ��U��s�k��)���}1K���v�f�7ڸ!�E�)���)�=B��U�������J��%�=8<����z��5���Ώ ����U�z��3~u�+"��.I�hBzTӄ=�`��?���PzU��?��Og˪�,���6��,���#9��7D<�~#3�˩Kq]g���)
m��1�oǶ^XYl(��z�Y��IcWtdAs��wB]k��yWWxQ��<+��;�y���.}ʊ�I�mX��^��F),��܌U�{|�rm;���j `�V��mF~�DDEҶ�Oj�ܫ0�B��Ƈ^>ưk�6T��dMόM���؋ˢ3'*-�nz}���{j1��96!��&r�LeӺV�e��֔u�b�~ʎ꼯��m]88n����,�4��0`c@��Q�WǍ�l��j�}�c��@���exӯ��nb���f��ZǨ����f��*��t~�t'��J�+p�;I�_����˅��h�����u��{��x�B��Sg�EH�������5�\��>�.�������]*B��
xEYG�<����z]���JԴ1���2j�Ml��1B}����ޚ�e��Ysu���29�U銔��=4̩[^�(G@O��T�C��N��M?1��BvL�N����i�ް�t!�����w�Bz3o�����|u�x���H�n�^q���Q��%v�	ZF�tЂh�/]��E�6H��Pҍ�ܣ:�5���E0���^�]���c��
�Y��,f�B���I��y.΀�75`|]g[MYyx����O%`gVf{���J�.o�-��ZER���	+R�ͼ���Sq��ͽ�=K�nG+��N�F��ٓkO+���Z�i"�{x��9��cG�Jm�ڙ=+������52��5lq�j+tu&Moegc�h��z��M�8K�r��&����<Q��	���q��ޖ��h
fk��)KȀ(�l]!�n��!ˊ�hU���=����� �ou�@��Nn��#�`߳=[�"�1*33���8̸�>ճy�=����,U��^��|�����s[`X�Q��ٹ�Y�Y=�JS�O>9����'P'�8{����βi��l����`d^;�ޔ�ɏBݵ}��k�un��G)�:ܤ��~��V�nnPbb�N.���z�]z�X���2f�z�~��3�\,*gi�������֥v��w��Y�YoKjUپ��A��[�o�F݉Q�ٜ#
�ہ��j��|��J�7���-޽E7�8��E�O^%h�"�����tێ	σF��o�ۭY\Zy�C�;y���;�oU]����p����ZzQ;9f�̣M+4�Q��lv�V����&�oR{e"�\r�vw��5�	K�|��N��3� 
ܸ/[��w:6!�8��싕����!����|s�W�RA����{�ا��ip�Eѭr4 k�Āu������,]�rTx�lajW�޾�y�9%L�Y�W��]T5�a�q@w�]�J;�1�5����V��NDm�P��[�3^����e:fl�[&��PA��9v�5��|�`4���69S���ƫ���;�1_sȩ�M���:�:iVJ_n���0l,vuD"�]묳@��rW;7Y6�.wX���F�x��YX��(���}{R�;�'7Ԕ�ğ�C��j�J�T*�,U`�T���B�\�,�b�gL�h�* �T�dDn\��DQT�U�F[U������1+�V�ٕs%�[˗��Eb">�3T̢ QDK���ks.*��Y��aT�9k���e�4�XY�TW-W)U�8ʪ���`��lV
�(��U��>����cQ+bV,��R+��X��+AU
%F�� �JƁH��%TX�YkAT���kUQX�b�ڢֱQX��Um��r��DQ �����i�B����f$_�!�-�����U1��ǡR��p�"�����"#u:4��c�ɯht>�������l
�Y�C���:��9d��&����Y��eOZ�\NY1��-I� ��x�n��Y�\o������^�L6�H(y�&:I�1�j�H,�'>fi��PSGT8CL�&!��'�o/�:�96Ö�8�z�Y�%N�TU����Z<���}���1 ��r��Xv��s�i �W2O2����+1'n py�)�����H(T8Lgi��IQ@�Vv��ä��^מ���3��߾o^��T=��%g(o�4���Y5޲m��׾`x`V�y'�E�2W�K�/^ag���7�d4�Aza���z>���Ϣ2���U�ϋ_+��=��`Y_*)�>Î0�H,�e��1�(oۤ��SoL�@Qa���g��gvb���凌*1����L��ީ���By;�<\-�4���Θz��'H+�Xv��i��z�i�mE�����i��\I�1N�L4�Y4u�M3�J���$�
�x�b_w�_s�+���x�"6c�1WLFϠO�Ϣ�E�9@��2�������i �!����힦yHT��9��:�E��VbOI��H/h�9�^��\���\�����_}�t�gI�C��"����;N=�i���<�IXt¦���z�Y�%@Qg�9�4��*CT�h�Y����\Ø��� >�1��9��x���硦t�^Y/�y�I�2W|��i��͞Rk��i'�T��� �]� (����P�+���:Nwf�
C�N�*�tr]g~��ær�Xyl<I_5�4öR^��Ι+:�̇���Y�8憑d�=�>0+Z����<��)��2�3l9L`up>�[��͏3߸Y���ؕ��&V*�V����E�ܷ���ow*��&���V�b���~޺ 6��}�I�a/���lޮ0_d\.��wU��L��Iw�O⪫練H�ӿ9�yH9d�1><a��Ι�x�Y79��NP��&	'�WǮ��6æ���!����sM *�d�I�7�Ol
ç\u��{�9�wϺ��9�zyHT
�����(�`VbNCT��J�9{C5���8a��J�����=�T���+���l8<�Y�%�v�:�7�/��4�}�d�D�L��}2g��}S�
����Aa��gl����0�}{��R1&�}d���6{a�z�!��&$7l���M (�:��F癜�9���Ř�
�Sh�hcz�!��ɣ9֢�*�-�+;d�֬���W�:a�+
�(rqMqHVc%}O{�)�t6LE�֤������ߜ��{���X����H)�9a�iEm"��v���*Aq'Iǹ�a�
�Se�啞2V՘�M�Y�8:�i'�js���i�fy��߾�/^o���^���
�3ިiEY3�c+%H.s�@�Ru|a��
�~P�i���.�T��Iˉ�u�i �Cfu��÷�1�q�b!�T��l�,|�|u���0��)_DD�J����S�H,7Ն=�IXc5�4�Y�%�96ɤk�2M3*NЩ�q��i�aS�
����x�^����*Aglw���5�q��sμ����]�v�Q`V�`]�q͆��@Rl�ᕘ��ɳ�1�1B�9�����19��i ���3l�]f�Vc%p���߻�מ����u�0�C�����T�gL8�4ΘT���kY6�'�H/,
÷�3�n�;a�b�o�3��0�v�]$�^d�TǢ����}r+u��V'�\���>�O�U�I���wՆ�
J���N�P1�L+����p�Y�Y1EXi
ͲV�}`W�whv��HT5�&3L��!9��8������|����fBۇ�V�)V�Ro����:+PI4	*= X��y���N�m�ô����WZ�y4��.d��7�b�h[S�{[r��d�+GS`���ꯪ��������9���Ag)>s�H)��ydҳ��0ߖ��Vr�'Y������M'L1 ���c�����Ă�Xrq�gl� ��J��+5��u�'<y�ε����x�N�h�OP�aS�Mst�Y�%{���i ��Ę��Qd��{���H)��-Af$����8��P�6w�s�u��;�<��O�� y�!��9d� �'�N�sI��qՓ�N����9����� o�U�8׽��]{ϳ�x�I����p���@Ă�����T�S<egl�e ��
��;�Rm ����<�c��c���z��2i �7����<�w�<���I�:d�<B�`W�y�m�0�R6���P֩1 �Hk�z� �7ohXt��'F���Vx��a�����i=}dă�w�=��o<�o�]u׾�=zAt�%g���H,�����%@բ�Y+;d�0*t�^��T�a�<CĂ��p[�,��$���ɧ�J����/�'����Z|�uƻ�|�$��̝ ��w�⤬5l��'I��m�l*AuՁ�풳VȰ�g�Ѯ�6�P��R�l+Y�L�!Y���py��^w��6�;�'�c:d��jgY��������I���1�0�1�~u�I�0�ީ ��!�4ö�0��2��e���+מ��k~o޺�߇�$zY�{x@����T�����VJ�\�f@Y�%B��l
��ea�Ձ���Af�:�o�`H,���r� �u��{�{��}�^�x@��N���xA@�+��,4�Xr�&'�����T���%y��0�̓L�J�]��x�Y�E�:@�o6��4§)���γb��wd5�6�3L?P�69��T)�#1bѕ��1_X׽'K����WZ����b���eԱ\�7۱^.�Yڲr�V�}�Gy�*�!ڮ�����W "n+�b�~��z=
���E~�d�r�����x�Hjk2r�_Y*)��<0/�{OY����[<Ae@S�H,��Nl��^�h����GtĂ��]y�]����}q���$�³O��bAC���`i�a���R^)
��Ɍ��O-Vp�Qa���Ax`s� � �6���&0�Vb)�0�[i��²�+�Ǣf=����'�s��ݓ:ef3^P��N^�fqdĂ�d*{x@�8Xc��)6qC�%@^��d�����"�g֯�|��W�A�l�q�>�>���X�VOx�zE �n$��Aa�Ն> Ua�I�i �v���a��
,�2�I�x��ĜM�Ă�ņ��0�H.���<��/p4Ι*�Qgl��!��H)�'n=0+0��� ��'�1��J����g�������^��:�0�;g	�a�Y�*^��=�޼����H,���R�a͝!���9B�t����XvºꜲi ��:�i�Xv�b�(m1��ی咳�;���풢˳��]��݉��%��Ǣgf=�׮}��!���:a�c7ņ"�Y�p��I�i��z�a�
�u`c'���}d�@QI��`i�sd��I���g<�F������|�0�6�̡��&3�Jɮ�"���k
A|`^��0��Ó��6�Y�N�����f$�Ă�Y/�V��s1虈���bG�V)�������}3��@Q|d�c9Ob�)1 �1MgX�l+Mg���TѪLE��Vx�)����٧�a�=��T��|dǖK�+o�����[���u�w~C�v�^�=:�
Az`]qޡ�z�9d�Y�*N�i��v�=LH)끰�0�Cz�ĂΙ�hiE�hUgl�=0<�\n��V�w@��v��U% QFl����Y�b�����av4�맚�;��Sj�㺶�n��(��-z�GC-�b�j\���)��;j�9}IQ��^�9���I�τ$�/=���/��p���m�!�K�&��ᒳ�3��9d��=̇����,4���m*Agl:L��H,�C�AM$��$�ô5|7x�z��y��o� �c+�t�H
(jZr�g{�c&��x�}yd�۶��8aS=�c<d�9�f"��!�����4o3�a�՚�LH,�޹�fuپ��q��7�=k��x��Eܦ2��Ă��U�OP�AI�z��S�����J����4w�M0�d�Y��ě-�t�Q��{��L��os��d� ���a�R�'�Vi9@��Z�d�,��Vr2Vr�_P��)��&ya�z�$���YY�[���f�<��S�o�{λ�{�|�������X�Yӫ�H
,*k�4�+\�C��!Sz�l4�	/sa�r�Y���m �4u���A͓L<AjN����޼뮽����{�aPR�S���
�$���B�N����3*�k�!�wœ��&$�
��Í���9aS�
ͲT߾�癛�qߝ��I�*�YS��]2{�4�Xx����Af��'y@QI�(c4��'�ϗ��T=f���u%���;����z�Sh���Z����ָ1\,`�ü�r�*���(@"n%�+�F`����o�z��<8���5���5U{����fWFJ�`��K�)i�L֯���g�Ӭ+��3)�W=���[�˃G��o��+�6H�+�C���豲N����x��lb���.�˹��PM�Y�b����u_P�g,������Y��5]�s�u��yq��7����ӑ��68�!�r����G���u�K��I�x���M�j�ř�
O+���^κō�ꬮ#�Xyt�<�b��[����i�\鋡�R>����:
Ѣ���Mev�e����l�ޱoX�*i���A��;&m�m��nʝ����NO����A�xX����_.��pU�è`��kץwL��m���S+G�NGTd���$��yNVW�@�/K#6����Y5� ���+.�����u�
C��WT���[㬮�/�߅���SQ.rL��`�ӟlKLt�~[ғ��8tk�ӓ������c�o��wR�.���3�MHh9��̰Ķ�Xp��)ٙ.:���W�F��s���*H��9�p�F��sΣC9��U Q��Fi�u�i�C�g��ϱV��W�Et9���(R���4�uǪ�_Lqt/�k-�e|S�b�B�4���iBltKk�K(Bp�ȑծ�2�S�3��vg��r���5qS���\#6�M�m��*G��\��B�=ʧ9�\�g#U���Ε0�0=U�Y0%��P�f��ȩUx��ւ�������վ� ����X�pAWJ�h�,nP4H�>���[�~O��|�H��2ա���UvJ������T���h3�����qb�Vϩ��j�)���ҞД�W�E����ѿf;��7�r�eMK��D>W���XS�ab�C�[x������4s���C�U���^Uch�����i����m���"��{���:�·H�\�1�7����!ì�� qxCˋ���=�]�E�][d`t>+�鍺|2������oO��_-kET�pS�&�6T��z��� ��f���U�q�q�EY
��E�u���i������D�{�*�]�h&ǕAvm:���v�;E֥�L���M=�!��R�G�	Ή �vgm��`N���ط�{��w|Zcw'��9���x�
��Z+0��Җ:���j��Nho>��M��R��LK�3**:ORU�k��9ԩJ'�)�^�(�1.5��O"U��ڙw�b���K{V%�(ukӕ^ιGu���qT&9f��:=C�w�5�Q��C�5èVX縊��g�9�-�/�J٨��s;77&b�%lcf��}WX�u^!Q��ҕqAB��O��@z�l���1�+5kGS񧖺�![�u��ۏ�}���U���AU\����3�<,V|��ڌ�6m��m���k��Ez���+��1Í��C/�@-�0c7&y-8�`�K�ɇ�B��;lAGM�ʘA�7�N\ۨ�7�Xr;������Ţ�D�G�A;U�V���2�v�j�^V%����ؖ��h0�2�k��$� ��OE�t�׊��ڼT���1��������s��Ǡ�.��u='�)�}��oC� �G�w.��u%}s�fٕ�Dz=��n�)��1�eB�*xm��3iX�v��������(�X��:7�n�I���rf�rD^s�v�/�?�2����Yw�����洔��a�ױXJ�Ԩ�3XEI��rg�vݰ�(�wr.��Tn_K,�R$�4=Ӎ;��
%ό:����@��Ѯ]Szt�r��t��{�����s�`��g�k5�x}�-W��nIY�N���pU�>UPV|6yhc� *�j�gF�y~n�󾓽˯n�E�M@V�ɇ�R��k�dɹ{62(�7{�;�|G��[�W�b��� �p���yI1�M�B�Y#l����T�wu(����H+�0�W5g�(Gs�8C	���Tɉq�\�_'u�t�Y���ȶL��z��b�`�ORL��WgwUUa;\��B�h�W�W{8!M\��v*}��qvNrBv�O 7x����p�7]�\�s��l�]]�
�s2��>}��C�נ@�:뮹�<�Xt���y����}p}�w
��Ŋ74K�SĐ�N��Q|����g���){���g��)K�láɘ�J�f�mx��δ�BC�/�T���7���/�KM�o�j�ܻ��X\~ѝ�x����L;A:���F���wToI�6�ݗ��gxW����xe���85�����V��}��^�y�	�z���?
^,�5:P��==���L�ݷ��|���#%H��Ӳ�H�7ǹSLUr�ɸ��Q3n�P��7�0bH�*�p��� �˅���/�
����xu^�Nj�-�і��5�g}�7�pV!}j��)Q�s��o��9G�=Rݨ��{��Y�	0�vWH�*9U�ҕ����sޏШ^˨�+W`�U���Yq���g�K�7�M&-v늨�7��g_6ҽ�r
Rsq=��\$�K.8�CO�[��K�͵Y�o�C%]vw(�cq��M�mP#v��=#�����S�����T^���mLa���#,67���5+�e��fbp�Eef�0ե��Y[WPU��:�2�e�<Jݠ���/��"�Ʈ��=x�t��&�5W;uvQ4�W��:�r�Y�m&�p}�ګ��0(�a�H�n���(+:�E�t����L���짃a��L�#:IN]������9f����Ab��̅ä�l�T%k]���@�i\	�v���"*7��=��9^i�4�av��.�Z�2�HQJ��]�[9�n����f��!F,��9Mѓ
����X��o[W���tP�M�x��.�X=	R�����%�����;�:Suo_݁�����Y*�c����(�hc�K�K���b̨*;8�P�Ow3|-1 �lg$4��OY��{6��z�7[���YN:�o㧷1>|���7�:��7/kN5��>�U�֪�;�٢�BҨ���KJ�5.]�v�o7f��e^�bE��j�bC�0��g&�TC��[�R
��B��B���:(s{�H���o㆞�+Gũ���8'.ё���\�tغ��ض�4`���YƢ��#�[r�� 7n:(��|��x��ӵ��Q�y���In�"*���XD�s~��`�8%�]*��Z-H4�6*�����9]����]��^f1bېa	!,�k��qh�����:ep����c��Q^���̩ȫ�`�ɦ����Q�T�]m�M�ի;�c/c��2�(�J�?��:b������ڊ[@a=׭0s�9��I��t�W��`y���'�\!��L
fGh����X�T��{Zв,X=��A�rZ�{+@�6�b�M���MՈ�V����5[A���n�� i<�Գ9>ׇ{z����O�;���h�R3���Kh��,UEV�b**D"�DF#ib
�Ԭc��2*)Tjkb	b��E��ŉR��b��TV�$P�Q�AX�V�X�TEU+APaiEAEdTPE��ʌ񥥕�mU�b\�®+M[ZeKV-aXԪZ�X�1%QAA0[EE-���\��j��ŷY����m�AR).��Ġ����EU��F������5w�J�`�YZݤxt����֮��H��\�)�(v���η�����}_h29���e�A��Z�
����ZV h�V�>]w�]aI�&N��&�{\W�W�Vi���kE,0h�lhbeDlY�da�`��}<�;�����v>}��a
�u��1q;*@��9a�;m�k�E*0�ޡ7�ȸ�31��s�3j��D�d0 ����Z��9�����j?����c]A;U�V5��D-:
�2���c��)k�ȘɎ~f&rJk�;a_*�z���8�xR�yzO>�����#�t���lfRX,Q�^@f�]y:F�V+�Ѧj[Z��ң\=�i�a�q��u�y8� ���S6q�����)�e�y����14>��_z�M/��s�-)�R���˹}�o+���j��+%C�'�P��C��L|��5ҵ;�=]�\Jy����Z�"��h������K3v{k�Dל�ӹ����̀1����ݩ����Y]n��X�VL�?�n�Zd�#2׎�+�f5X�[K��z=���
��2�\"~��v�2cgf���i���!J�&aO
��ݥ�-�"�U�G:5i�Y��I�`�|5�}c^ہ���� �5������\�@� �ڡ���쥢]>G_3^Ɍ�����˻�󅠺��bG�])��V4$pk�Ls��P6<+�>6oט��ي���k B��}p�D�@�l��>R��F<�1Rp��H횖j�n$���]*��R������i�~-u�B�ВiZ&#%�ˋ�<�'f��S;�l	n�[U2������힢zw|T�j�{��?*���V:��4s�+��Pnq��v��t��Wf  �8V3��Ja�J��uVkfWO�g7���E��b��P583_���S�P�j��Fʽ����]N˝�lSO��נ�T���S
[�-hzn���(��7kZ�*ķq6���s���y�d�l	�n�.V�{Ү�@�s$]�7��;��F���{���z�N��}�^:ǰ�bT�>��dMqi� �W��9M����Y~2��'.4s�hDi
����u�9,h�P*\�q>�֞eI��L�7�
u�["z%L ���t�ͺ���m��(AmFe%(���D�P�n�f�}-�^a\���0&�������Z�8׬�R�j���f���⬲�;w�#ϗ��xr�x(��rRg�GG^��01�</�V�����j���eq�u���;;���uq�-�����B�UO:�Ѣƈ�tkZ ˼$D!d�h�qx6T�їd{�co##@Q.|cX�FWN@�q���r�f.N���!G�k�����x:\���vE�����\P|�(��.N<���^Ŵ��WcYu�^z t�pU�kw�'����B�4� �n�ݳڶ��5Ӑ͸9.C)��V�uMv�Q%�&�:��MH��R��-fǴQ�Tg,-X�O���z]�_K�s�̳�MRԢ.�p���8���%
R�ѡjɪ��G���v8�ei�;#�m�UI�S0��yQ����"3Pڋݪץ�|��O�����Œ� 쪑�Wǽ�N�.���UF���<1�P�9�*��׶��gbvL��'3�ɽb�ކR�YnMF
��A[��9��`��A#�g��3�D=Aځ�d䩈���t��2=&�p��P��ꀭ�Y�5��--�*�)Ȩ�����	�1^�ƣ�(WN�N�6,[�擗�ҟP��o`%���%��C����|�|�۠D�/��~�or���Ã������*����ڟn�2�T\uN�b-��k�:	���@��5]��[��X�J��)�!��$�}�J���~ʂ�uQ��Qr{!\5��p)���R�Yj��{�ֹ+p��f]N�o-M$���]m3�m7GX����֦Q]ܩ�2	������ne_cY���"�b��Dz�4Rsq��I�#l9�Nzu�)�^�L��\�$DdLc=�E�DQ=٩���^wF|97<S�~�:�L��JTM�rB��7��n�J�7�26�
����)ި�9��P;}7��s2��-�>���d9ɮ����5����vxu�^4�+���qo6�HZ�}�ļ� ȴ<jh�ul���9�pXs%Ϸ��.yJ�oJr�;��]B�����_*&�R���F����]/]�򸾿o�"��~�- {{��Զ�Rv�Nʐ��b��#���A?y�Y�1�f�koQ�G����ۑ�2ڻüUq���n��WF��x��]A;U�V5��D-:	��g e�2%�鞩�S�U��0%�����{)�j5ѹH:0s��S���f��3�ԣ���㙤t�:i�i�V=S���F*�]X�;:��.�z������Rn���Z�G}w�e!S0�1u�*	�������2�f܃;1�S�VM!��:<s��ŕ��͠p}<>���%}�	4�Ɨ����V��^���N��°��T�	c޺��w��3Pz�h���~J���X�i��%���)�E)B�	~�$ݜ䋾�.���xt����%�"����>�>�3ұ;�<�����7�.�O�D��ȰQf�*��1�U��{N�
T�܇����jJ|:aK�Rz*�|h��9U%_>x<5�}c^ۦ�(OnߚG��qW���w��ܳP+�IX�A�)r��T���0M��6�{Ŗ�mt�p󅀺���C"�
`N̼��;��o���9���y]�Ovd����.l�Ƭ'�TLAޅfc�h��ͷ�<�BP/��Px:<��<2���CƴCԩi�/�ݮ���ce�5k�W��1g�0U�(��ur�k���*P˗��r�n^�Θ6�3L,���n�mI�rv�f�������l�z뭎��֗{|�j\F�/t3�2B�W�=���<�[5s��b�.j�:�C�@�� }��a:1�:2�Y�kp��=Ӻ"f��r'xh	������g;��@<�������	�kF?�B��łâ�*9S�O��,�Ж�����o����#�? ~�5��*J҈�6�kG��b��3��[Ŭ0r�|��!X�&iW�MU��;��sџT�M�칙��z>�=P�Z�k�?�T�s����t��o��u�y3r���wv�|�N��J���S�AGM�ʘA�.\�;��Y��������#.��i�(�D~�WQ�-<���uxΚ���z����܀����@0h�ႬYǨ�]�����pv���6�.��ߓi�������,B%ӱq�:�T��p��P:��i�6��Qq�f+�Q(�ɭ���%M�f��XTb���[MC�q����:�W+��-c����P,镛��U�˔�۩��/m� ]��X�dۍ����EӶ�OE]F�L,B,�����>�c�V��ƇA
��kHl�Mg!��U�#+���S�J]���<��zx�c�];�qWGm��k���kk���τ�a���xp��E���6�7'	�x�e�����
�4�����E�f�X<tUq�^����ӳ:v]T^2S��?�|h��J��Eg�?yu��B��z��kzL��|����C��W���+�'�L3(f_�RLAT�މ&'ѥP���@n���tO��0<67���ݙ˛ާ#f+i����S���J��Je�D}��)�x�>T���3��ȹ�;�0U�Z��j�����W�¸u�}}�f5�Y
&���Hj�U��}�P�qb���nm��'�l�}�uL|t��h�4�+[W���аS������f�o�]oM���T�-⏗f�jE��s��A@�S����1*�*ͅ��R��d�=�c�M ��Hڏ��yM{��^����#�lV��/
����%w�L��9&_��:-֭$�5c��%PR��h/�Wz���z��u�69�/p�@VVmR��zh��h��bs3>��W��;��U>�w�I�N��
��Us	��S��[�Bo*Z��G���H,�@�|�z���9aM�s�q�B�u��c<�J�"!�և(���m&r`C�ӭ��<>�:,T������¶�pT�n%��3I��Q/�Q�tzf��b�W
u�ν��W	Ϻ�"�t�5��Jp�z��V���U�:3��CΨ)��+����0�/>⶝�u����ʸ>?m��a����mxV���M'Iy�><�pj�Y��
&(�5i
&�R��H��[���L�*� �	��w� �������]G�gn��Ӟ�&�t�������r�l�"�.r5���H�:�8��G�Uy+�1i<n�ڳ:u	�j�G��}?}_WՐ$ZO+�o�����D3(��J�q�\"�ݩ���nj2ݥn�$��E@���U}kl��/�U U�#\�{^p��W^���O��,�vk�ح1'��(��0��k��Fb�H�-��1Çω�k6(�s�W5��1;1ʠp���4T�8u/�ւ�`*�h��e%��5���t|���}���r�#�p�mAY����������X��N�V0UA�o1z��ss9*zL�R��ί��o�a�t�w!_�A�}P�_$��8��YX"\�J|Ut��I����G�#鏕}1ƺV��LW\�eo7�V�)�����Q*�E��3XC^�V3(փ�;K�T�Ը�'�<�n�ҿI�z�P�'�4kl���|�:���/�l��+ؽ�+|�ۂΎ�i��
 �{9��]�����gEH����Ks+:�i�
{ǰ�Ɏ�KS��[+�s6��֥�M�>M��U��)��׌�l�pyb�$�jء�C�R�lu4.�r^eҙ�J�f�Υ�kӯONr"oF�Qa<��\�^��)n�+��ٝ��u�X�{�1T�俹"&�]��qm��[h�vh�;�]]a>��ї��z�l<��ۅ�9��cx+>�{�IZav����|�!�M��F h�Gz�P��W|�;&�Ki]��a�sD`���;c1����q��-b��<�+c�<,��{B�ޤMU��ŧ����ռ.*M8 զ��ɗ,+GGK6K=��kW�p�[S�|�5\
�����S��m�j�hb ��f*Bd�1cݦ.��q6_a=M�L%��9e֨�U��BZ�aW¹\QsC��!��ҨJ��R��{�+�zUJB�Ң�Zl*r�F\���Z7��n�]w�[t�k�A����q�8�]V8M�-QL�x����,�:����i�I�`H�d�t���t6gR�N}:uh�1U�E��L�ם��ǐ)��z�2'�XߵV�8�O�6��ڲ��a:��*�ȅH%N��$�� tm<Wu3�'gIc�˾��D⸸:�8-�W����u&G��1���=@�U��ʔ�Dg��rח�f���\��W��PMHku_#nĴQq<r���uԺ���n�d;-��>@Uţ3h>ˊ<�������p"��$��f4QJ��W���¾�n!��ut"����jԄ.[�gB����ѻ}x���kNڮ�p��.��.�b!�GhZ؍�#�:fd��CԖh�@�Ӵ�^�M��kU�]�I�;�qބ�<�%�J�h�WRJF��c�#ŃoS��W`*�
��J_7���wwnA_�W�"�������,�*+�xJ����*�Z�Tq+FTib�����*����k5Pը��b���������K#6�(�,UUc��ņ���B�`�T`���T�q,D�9n�LTMը��D!R��ڈ*��TT;�#r�V�"ț�t5��U��ETE������������V�U[ePkL���b
���*!��YEQ#iX�D��!�8烜�y9ߧ�����e� K[��8���r�1S�绽�[$[�:���;ﾯ�s|����P��zW)ƽƪ��Zlk��` �<~Wʑ�����s}���}L��}~u��G�ډ�1�r8\�<Q�f��-ɋqJL��b�V�A�j��|�D���c���2g�py֖�ޟ!|j�U�7W���pR��ZR� �5~U�i�*9x�[i�ϥX�4h���W���v�=��V��f֌�tN&�.9!���qH�Bc�uÑ+k�l']"TI��r2��=Չ��Q�M`�`�@�|m�,ȱ�J�N�zD��l��f[�*�K�>�2��5ưk�QZ�Ŋ�Ώ�s\ ��*�}(�\[��lLBu���^���HJ���p%��1l:x#z�y���s��b�s��2g��+�� �,׮�߻jX�b�Ϗ��ɾ�~�~�z�&5;3����γd�3����p�ۡ���)�]Q����Oz�_R=�LL���s�{���Vc�c��`��v�e���a���=�y^w�H�?�V�^\�q]�b�k¤
��Cdʹ��H^6�j�ɹ�:�a����h*f��X/ر}�,�(z����]/3�!Y�%�)��6T�rg�0l�u���fQC8;����)_OD��W^|�mdrv�znM��LA�W���'t@�<�F�@�[�(b�ڍ����1�U�TU9bc��3SL.D��;���8)�)a�G��u������l(��^0��3y�{c`Y�ǉ2��5>�Uk�F�WY�|l4`ᴹV���s��u͵�'b�tB��?u{�N���Eڮp�ƣ��Kˇ��ê}���B�wUrk���g�H�K�@��Cuj���JuO��qŝ���&m���'�h}�{�aA�� D����T��dm�咐(��9���8s�)��8^���HY,�6����\:Q��������e��ܚ�\�Ap��r�3�<uՔ�ھ+7Ndg4�bn��s���&L��0CN�goq���.VMJ�S�0Gވ��S������Z�P�����tB~�@�k�huv�2'$p(�}��Ö��)���� �=V�T>��^�;������W��浿9�̑�"�R�j�����F��(פל�V�������c��:��U�xŐƕ1޵Hlī>�yU�;���{	.�v��L�C�g�<�|�B��J��7�T�������*���a��eL��&�+~���Ҩ)P�����+vΕ٩�j��9�T�%���A�C=��~c����Θv*1p/'==u��K�,���g���yVq�[�l�&���I�;h�jL�����90���\���b�k��1��T$�^���m//wSU��T8�+�r+�����I)پ�өo��Uw4���d���EC���s�T�Gu`oB۔�Z�s*ڌL"��n��Crs�-�y�X�R��"xWR�C�t�8֗]Rrk�{�_r(�y�LA�P�W��TK�E����1�s yJ������;��ڻڹkC�����V>Z1��Q#�H�a���oQ���}vW#$Ɂ%���+$��\��KFX@�1�կ�Vck����lOO�'���3^�WQHxUA���3{K=���<a��3�dM�=�0�:�P��_�a
�rt�WJ�����ᢽP�H�'�땯aA���b����0^9��Z�{xM�l�#�ׇ�&�l8+ä_!*w�:ƺ����GX�����'��M��Z�4h�� 0VݶE!{�|(�U
�C�Sj,��\�]��ԸM�+o�b�
բ�M�(�^�o�s�{s7͊�#��c|sM,�bi�a��t�3Pv�7����&+�����1��̮�u̸P�e��] [����e,=)�����Gr�h��Ks9)���0�ll�Ք�:=igR�u?��.��uK������{eF��FULޏ,�ċx�D~����鸓="W^U��A��t�s����>�Q���p�Q�Pp>ׁϓ�;�d��\�P��>5��+��O*U��=s�[����>�%Y��{���ӱT�K^�:,H]��0�����J�tf�J{��gE�[f
1����|g��R~�y����TG��4>5V0<0a6*a��mv�����8�ɍU�t���<��:jTH�D��ډ�"zL�����MV�~�� lh����N����)Ut^���bd+3|���zSx�LA�ʋx�0�vxp^8)U*���*U����Y����_amK��NO��r��I��욲 Ca�v�\��>����5�U=��������q�%����BP��*���|�=��_U�{��q֒�\��iP4ޟ���w@- ��y����;D�u��0�*�F�7�k��S�Ys��`:�V��fi��eGƳ>�h�F-�ؼ��Q�Y�?��o\�Ԙi�
�+"!}�^��@��5����P�N��H�׽.�!P��w�Y̅Z~ ��X5�Sl�2͆�G�ua̹���榌�ڋ�10��^Ma
�|t�踣G5���~����l���0��YR/�c�\�k�?�uJ�s�XxQ�h�Ku�^��z�p�7� �}ARj�)�p�^U�V�]�����
�y̡�S�����Q�Tٸ�P#�)��y`���,_hm-�y\��v)+�j�CVʭ64hᢲ�
�z����"&:ю�:.qu���������ma�'j:A�*R��"��
M
��n�c�m̕���k���/�Lu��K���`�r%GT��3�	�%�m���=G�v�����L����	�w�K�VT����W��Nz������蹨�2��R�X<F;����TU���4�]Uk*T��PWID���-<A�f�v*5��vW.����S�)]�;�-�ғu�}?X�+�h�siOj9�6T�B:n9��N��#��g{ܞ�Y�Dz�|�
��#�^�҅�e���<�@���:I���{'~��c��r�X�f��b
S39�\6�v��l�W{����SƜ,c´2|9����r�h���� �V��zel̙����1Tƺ����2��	l�X�zĲ��~+�}i�8=�{���j�ߎK��u��)�K���������3+�c�&��\g���N�2�b��&�Mh!�&�����Cw��3T�E�V
1l܌{��@�YU6�!���`�Bo��y;^әզ"�IMn�gF}=ؒ����S���Ȏm/��˵h�$�P,�+��Vk�AW�o���
rW��K�K+u"�-u����eջ�S@�J7�y�,MR;���ɋ{�Y�lq��@h&�`�����{��/;vO�5���ܶw/ˬmO������|\4�q���hXrr(��P隗P*�Nd�K	�ը��q��5N������{�	��.E����)�
a틺��]Iq�!���L)㺎���XH&����z"��$�#V�)�I�JM�uz�s��jl����5���Օ���!{g��>�O![�i���4�%�<*�UQw[y��1Nn����n�`���Q	p�3Y
����m2�[�62�V��1Ы����Ws6��� ��ܜ>��mK/�Vx�'Uk���P�@f���.���]�ʑ�l�ڌ�i�����J���	�����]���\[�WG[.�:�[�����w���ZÁu%vx��pNӔ���t����"n��m������֏*=�7�,�̼Ox(��n(��6��y�qEJ~Y)��CZ<�x�m��I�*�ָE:;s��G'ѿqU�<s�2��	�V�Y�+��d�� ���n&o�������׆P5��w�?n���V�ӥ&x<��>]1�6�Ȼ��Zx�Zu�����&�DQb/y3Ǐ��s���nȭ޽���~�7��&je*{C���5�#׼p�������e��6ZE��޸��{#*��E�ą�6!No�m����U�ҁN�����:�
���@S�479��x�R�d��iA���?S6�� ��bܓ���^��X��<�u�����������6hu�۸��ϩj7ذ4�����n��^��+�՗2˔3�-���\��o����~�DqI���t�OS5*y
��A有��Dvw���C�z"���QLmfD���dJ�]2621
�kX\��;� TTv!��ta�m�C��y}Į[�L�*�W��Z�̦�][9�X��'k@��󻒚0�'�Gnx��rr7Nص����-Kv�ˬt�`g9ؽq��9�5q��:+��6U�b��+5�����Jδ<�T��u-�W�9�/v�^�c�A�1c���b1�'MSVi��=�o������,�N�RC�6�].�:��[��R�g�v�'J��
��M\N���������?\:�Z/����븻�',�l�r�!P�'u�z	0�*Pl�NI�/.*���n�����6����C�,M�Om���)����e<�r�Sw�!�z�F������5��<V|�&�o.�=�a��z3��f������5�t���0u�hEIY���f���T����Ҝf�!��m����ͧ��j����}��ݘ�V+a����їѬ��,�	�Q�ot��p�Ω��y�/g&u"W���C����,b`p�āap��k=��[��J�Ɲ�p ��7�l��`�lW-{��'ah������<,;�� ���y׌��𥛧��Gj����H*^dye+l��/�ɐ<5l[�Ū���F���sPH?M�R��Y��Y����I��y)�`��L�C�;�g�(7|m����f-qc,_bֵ5���B��hJ�0����ꄅC���$ؓj��i;H&�ZĜ;.�-��:�`�@]ej^$؎�彲��s��;���OQ~�t���=�Vu/m=�;�_wD>�:Py�!e�F����D�7[v�k�������]}��7qHP���51��_=g7�\��í��ŃVI�e:�n|����{]&;�N�ט��Cu�.�n���ű��.Khe�-ڈ]��t^=NF�Mu�-�xu�q�7Xs)L}�Xh���$v���M�����fN��6uۉc��#.m[����j�Ucp��I�:z�,Z�CB�U�s�gyɐ�y[w���h�uKEv��F�B�+5��L�OKܻ��
���+��^�c�}ai&�,���h1��ﶖ@ث�q�O��2R�EBͬ�S�L���S�[I`dI'#X�s#3u�h�˙���{(wmoVK�7�u�M=�`�ӓ�c�I�b�8��	�JJ��W�z��H�K�(�qj�o2*�:��Z��bTׂ�Ŏu-��3n���J�B�G�d7�Z��ur�ʬ˝B���gd�$�2La�n���ZΓ���y��w/]U� 0��J�e�R����y�V/T�ˬ1(��q�(����Ķ�Ȣȉm��F**�5�4�(��V*+fZ�EV�X(�K���*DEQ�\��0`��%j ��t�cwaV$P\eDb1ATX)�1Xbb���JU������Pq��E-�ҩ�X�kmB��+"�U�����fZ��EA`ZQVEuhLjԪ-k�Qr���i,�(��Re�F�����ߺǎX|3͈hc���-v�[���WWc0rҌ[Y%�*���\+�b�=2�U3X�}+B����etd^=��Y�����Go�9�;oN�lOJ6S��Wٮ�ˈTz��\˜�G��7PO&�G����rx^��őa����[��'*7�Wq�(�[��Ӳ�"�Yc+���e���q*�Nu��%I�(�����]z����k�xi�v��py�R�Ս�ϭ����G�+��h�D��o7:u9p�4	꘿np���xu�j/���߈@��"�̙=�W�f��,M)خ�R^%".�oI�P����D��'/��ޭ�f��.Μ}n�Fq�%'<������t��8V��j2�(�\���u�7�X͸[}�Ķ7�&d�GB-���'P���2����E�8����jD{��S����ێ�Y�Q��R�D'��V׬癝:���y�M�Sф`�/h�����.:�R��Mr��G=�Iv1]~׵J���ݥZ1���%��գ���l�Kn���ug��"��h���Þ��4��/��%�lH�z#�֙�N�N�#���-���]נ�4���p�Ð$��p�C�5����~��'w����mf�8�d���teG%��,��:���r6m������e�G��}���9hD4��"s��=Tg�]$.'v��-H�.��X�h�
��:+��d��TC�.ʾ�t�M%aؚ�ǡ��[�U�EX=g�^���i>��*|�L�;Nu��]�=���c�(���wc��.�邝rr���3�ݓ�9��������6�����w��Xj�����9���E:VJZw��
1��r�nRvC2aF�D%Һ�`V�0���.+F8�}���\���5�5c��8W]8���LgI���g ���)A��=�Gs�=�e��xÌU�r�].}���u1S7{�-j���/\�R襚�x߫ng}�ҁd�ۙ��P���o��A�6e�lV����Ž��[�6��4A��`�������"�i�].qC3�av�维�Dv�Ǯ���D�y��m��OP�"'V���g���3g���nz��o�������5|el�QR�x�+��܇/��Z�E('fnM��v4�q��ewi�i���5�9��R|����L�^����e̏���n�Rk�EӲ�|��V1t���}Wݴ{����̭��v>�W1�By��\U.��|{�u��)Ӹ�[�y��n>:l�b�؂(����n���/iCj^f��0#:�,�9��w�@d�jWK�ۇ<]<���9�.�<�k��n��e��K6ޓK�=uڄT$;*��!ϬS)c"�p�63�S��<hG2nGa�K�3����](�KgL�L��I�E8��%p��
�����8$ՏGȹ8��1V:�-�Ene����go�Y�КΆv-��=}�R���X��5dAn�2��3`��Z��0�T�d���n-�yu�U�"{�!|.�1�U�M�~ێg8s#���j0�ă�V�c�ٽ�� �`IbS�l����=&�u����96�DJ��ʑ����oTaZ
hAå��������]/�����^��EvH�l�K"�l]��\��I�n/���ߑ�C6if�.0=��[p��Z�]nKxG_,B�����2M\
��>~��n`�%',0"RS�nr���
+S��ko6*���䲲�Jǌ��}�Q�=f�!�^rYz�挗�2�찒��h�e[
&��t�7)��*���8{GU�;|
ٸ�,�0�%S�қ˫��.ɞ�ޭE�4��F���؞n޲���u��1@�=�1pޔ�/��ޞ�^gYT�f�Ѣ3�]4~��O9�3yF��<rc��H�c~��P��W��w�ʥ�x�,ռM�{�%n�D��7�ׯ9�:K�㬋�X �䣝�B����ާ(��ڝ4}I	Q��Ol@��� �oE�<s��)��ԷmE4i��D��@�Ƽ����u]�so�A��y#bp���s�C�W�����o7�֨�5�j
[�6�c}�"߱Bn������Q	�R���L�⸩�Y��p�$���>�^��s��-_���[��B>#��=e%��hJ��`ک
:�,d���]Ý��kA�r;e*�����mt���u{��N5�1�.RTZ���s��z����������s�mGK8�5Ϟ��V�<�J˃ �Dm�ν��Ir�3���!�
Sf-I�3��_RWC�GWt��]��¦%B�2�8��]o�j��|@=�4nH;�����:�[;ҋ�_qk��w�3�� -Sτjr�Ɉ&���r{�OV� n�[��ήo�� ��Aة��j-�G|/��f�kh^==
���ue7E�X�՛�s&j��>.�w�ٞ���x�{�v3�7��3W}�^���WS��w���<�n
T�j��+�Q�'e&�C��t��q(�L�1*(��0�aE��v^�Yѕw5'�����]�' <2�C��f]�/�\�S���Q���+)9�j^}�����uq�Mh�G��%g2�'Y�@��ަ�)��Єq�&U�Z<�H��"�'�l	rln�o��B��ݮy�/Ԯ�!�u���w/Fb�;`֒�^\�u'	��.��9%��»k$����=�f'Z�aĺ��e��s5�)���m�Z뺐2^�mLq�J$���+��E}b���H؎�I]��^�kv����{q��n#�h��VU�rڲw�o�ċFW'��2K�t^�5��#Qhj���/����|�oqL9yZ��?z8�����3{�~������n!f+&�NFv8E(�,__pZcf꨺JSk޴{R��(�FՕK��_a��	Ѧ �H�zl�{�ȅi�Ơ��:J4���M�A�\�i؀s�ZGy�j0(�9�/&[�wƻ���B������,���߂�v�`-t�n�IwT8���1p��{���Hj���x��x���<���/:��x�2ND �P[ENR!+��=u�x|燢r^xeݓ/�7��q�5�]D�C�\�������]��f�j�)��M�td��m��:'�A�w�Q���nh�_W�ل��r梨���ѩ��").��kn�~�rØY�ud��:�7T"�|�9r�1��j�	k�T������VJ���mU��W�Jw�G�85�]��J���g�|�b�

}bK�p��f�ݙx`�_5�`���[�EiB:�j�*���;Ho�j�����yu:*���Dr���E�׏A�I�
5C9nd��i�4�M��:�qT6�Yc��3�w&��t�"hD��d������y��X�ǻk˸��^QC�i�:� �4N�j^��o��b�5�d�kjvͨ�wwv�	m��2G�7�sw����B7���ڗ���W��&��6��t]�����U��u`̺��ܤ�#|I8�,܄ft�Wj
��Ѐ���k��ZH���, ����K{!Y@X�gqE^�n��P��v�M�b�f{�Ŭ��2�޲�q�Z�v�htcbTNp���9F�bգ/W=�����p�X���<��#�.���\�������/˃�,���h��s�8\�hh���7��n�l���=(�9�G����Rw�o����]��)�GO%�x�Bݶo����w�A%�3uo*'ݗ�+���[9�,ZO�;C��ѹ�I�a�J�Ż��Rn�煼�M�)�ʅN���U=�R�}>���EH�[�l��m�U�(�b-i{����,[�%]�M��k&M��Z�E�X���9oʾ�z����V�.h��yB��5t�.v%�E3�X�ʂ�Q7��������yz�Ӏ�k��>[wWF�C����E�"�$��v��F�����z�nv䃩�`[��|L��`|� �m-5|X5�*��d��ASЀ�X��4��Yn�$����[�����͑���9�w�+z�x��Q��v�����s<����4M쫓�����H�[�/X�x4h	����'ABP,��vjf�=q������n�������'��S��I�v�o�o[4�V�Su�,Y�G+�,w�o/���k�9+
Pv���{r\Nn��j���L���چ:h�-P&n\r�{C���Э���2�-�r���{x8s����w%�'V���z�93}x3�S`�u�W��L�N�b�{)^�/K�f$��$��H��QP�,<�R���x��)��	)r��T�`��Q2��U�n� �F��&�}��e��wi����tK)�D�H�Y�kZ�:�a�-��WMp���rRIQ8���n�P��=3�&:ccxd�jb��|f��`��;��{�8���:�辅L��$4�^�̇�<[m����cw+\����դ�Yjo��i���3u�$Ub�-�q�F*��ln���W$mn�o�� t!\�\w{-��;2B+��&��nIy�t��� ՙ��$���vU��NTv�R{��X8�Z��L���Ad�� �}nlU*�R�}��6��VMy�a��'Z��Z:���P���E�fR�V헯���z��Lk䀛�gn���Rb�D��QS�L_�tAze;]�'J��y�sn���	Q��&Ky����@2���Jsc���+u��Cr����\P]7��9�<��+�ʖ��(�E�F(�V��Y+%zJ�řeQ`Ԡ)Q�dU�PPKE(�T��U���*��J�[+��h�lb�ej��aZ���(Ņbʑed�)
�u����Pf%qQIR-U`�j�F�F0���aTb���X¨�N"��E�
"���eB�Im�R�Z�qRT*VV`�Z�`��4�b#�̰X��Ʀ"�Y*2�E��a�3(V�	X(1%n�L2��T+jU �,E%�%V�
�H�+� �U�D �%<�⫱���^�\;]�K+���l'�Wa���0��R���,�����2�3�FO�ˮM��~�;6gNA}�=e|_�S�k�w7w�c�ê�o.wW���ݝ���ѩ�d�7�����eV��t�;�ډ�EM���<`[
�}|�z��P�*�y��6���5���%'j�MN
J���)O~�2�v{ɺ�����D���ce�}
�4w���[7~F�n�{�:��;���0�smi@lݽ�@s��$@���������D�@�<j��<�	��9۔d�Ğim#̂"�N3q��>�a�+pm*	TɸX�l�@d����ʇ�� wC��e_�fND����
`l7Xɑ]�j�v)��s���m���O\�����rЛ��Ծ�3&�T���'m�%ǫs�Ū��5;8� �-5�/zVw>qJ�WV�iN���ɧ�c}����s��+������!��/.��t���y���t3��C�;P�vk�yf�[QM��mnE�e�✘q�>�5Z�;B�5�/�,�f�
Ֆ�h_	ȬN4.rL�BZ�N���ƇO�zs}��^�<'QO�y⧐d6*Bв�J�y}�[�]<��@�9��ƏA��V
�b�W5�Β�<�5{5�'ZO��=q���]�n��}s�q��,W�>j�fD^�͝�g���-����I|�iYv#��U��Ta�_7s�vS{w�����v9���P�6�*���8s�W�|���zf�tE��Lh-7m-����WV�m �Z�E�s:��b��ʹs)�qt⬻;�(��)���	��ЋFX��:��F��T�P7�7ǷI�^?�z�"["�&���-=kؖ�+BP8��m�D)=͞J�ungn)��喐;��yJ3S��{p��Z���\"u��"�V�aWX�`����Wj=�67[�;�ӧ"�.���te�+�����m�⌵ޫ�
�&{������6�k0�w⡝y�ćד>����u�g���κw�㶜�yB�~�������rst���fF��)�������88�Q����3LqGw�K�)�/�����c�Y��`���TTiC�4)]��2�`gJwE8�=nreN����yDnQ��y-��j�l���GUJ�e��
/T1�����z�Ed����%؞����+$��+�l�P{��y!�u���rg{ku�X��zK���G\�NX�٧hu6��c�M�������&�٥��x���"�[�m�Wp��_Cj�o#��J�=b��=���=���<�G�͋|���Ӌ�/w�\�9=�$;��
D�S<��\�>mmN�~�e<��G.SK��죞~�@Ʋ�=���.x�\V>�5`ۭ%{]�Y��+��Y�:�
β�
{'��s��a�N��	ڸg.���k=��X0�Y�c]�� �;��Ц*y��ޒ�.4��-u�9�� ��Q[�w$�%�ӽ�i���cO:]�I�3$�#ҊN�G${'��{{d�zl����]���Sɐ�9��긕?]g�ȍ ����"ʢ�h���5h};gb���b�9g�����>�3 /�|ͫ	E�Vi%0�#?F�ٽ�w6�w�A���s��A&�^�Q!���j��1�P�t5G 7�%��b,Ve��XsX��jx6q��^�V��&+��)A��A!-S=���yE��r�Y�ʧ��Wd]�������¶�.o:+V�uL��Z�J�ȋk-�M�j#��y�{|���u��m�j":���\Ne�\���m�x��N��1Q�[*��u�νܝ�Sa2�;(6{<�V�K�/�Ւ4'.no.b�Q��u��v<�(�]I�
����+^z�R弅߶�X$9GRv��{��NI�ux�~�L��'���AK`a�M��ܨ�[υ���Uor�1jj̫���cs����=4rR���ws��Lg�����z���Dvhđ�\Ҧ�o5^���7W����&��7�5�+�v��/^ͻ[�2x���Fc9浟p\�!�� hׄ��Ӏ���%�E[�Ę�QBYA���<hv�U���Dte]�M�X�y��R��Ѷ���z���Z?xLj�������9y��{s���j˵��9�ax�a���FO&Yi{޾�W�bP+}rZ�<�D�r�8G�o^�N��ҙ@n��S��)�#�鞹x���;���P�GQy;�����������W(e��[�t�o�r��ۮ�Th[�V�|Ha�Ӹ��u2�8�'0g�B��٣ulV�Mb|n�K��)Vfw(�vi����e��Q���7���^~�o���+R���A���0W@���o!�NN"���Z��~Z�-;p������w1����ɭ̜��7��p��o�x{T�Zy��~�Ҍ�;���>�Sͨ<�N}���ν�˴mOt��$0�����%�Эa�9�m���Dk��9J�:�s�Z��m��|)T�M�����>��Кh_�v���̑�vݢU�8������v�J:�1��R��N=��Ê�%A�O?��s�/t,���O{}�z�1��?;uD�!�/.j�y�5�Qu��F�e���t�R���;1�_*9��ŭ�H�m��2����J�0%--��.dn�6�(��]vXL����tTX�����F�T�{����{�i�.�iѬ޾� e���<ߧ��]��>�����Q�bc_$c���6Ӹ����hqp�&���b1��Z�	�5��2��{مxN�dh�y�'��(?��w�7=�Zjo��U�����y�z��\�o83�|���=e^�S��F��C�a��������k�G:�p�F��s�WΞ���m��3i�1<�W#�ȱz���do����voU�.ʐ!�c{��w�^��좷�c�lp������g{�F�{.�2�K:�n�(N�}�k��D5^��e�<��������Sn�0׶�y'�{�����+�dN�	:U�H��G.�k)��w�s �`ײ�Z��:�%��@>�Z9��]��	q���d�ޜ���o�ү����J�\^���<k�EYӞ�Ӳo�;�&y:��0�Nϡ��tTq8	�o)Uv�;J�E��5�u�S�4KO��=*�8�e����|�R�{5oa]��I�=0�:����{[C�c�5Z�dF�B��՗B6�R��k��;a(��s�lE�P>߭
�";ؤ�=����
�W��K7��8נ�Tm-U<"' �%��t�[+S`Z���1Sɐ܌��Y�T�����xw�8�\.��#��5��{y����uo��\禇��V�K��/S_`�u����ς0�F�e>�zU,T
H�)n:����'�R�tz��7mu�W�>�_Q�����f]E���{]!ۨ��::pv���x0�|����Ur�^���}���w�41#��7�g:n�y梞	���3�Χ�/���Ա����Ͳ�T��x=^UU��-2�_��[��h�At4�t�g{Ov�XZHȀ�߰�<�H�l�Bb��pw˚�	��Ic������v�M����m�-�ǹ��g_j�q�B��E[
��9׽�'����Ts��EUDm���{w^i>��f\R�x�U�ԋ���{j���ևDv�My���C�������,��vqU�H���*}� ����`*���"]*���q���1�"�^�=y7t�*�����w�g`���(����V��	i_	I.�6�ur�k�gD2>5r.PO+V y�;�"�!��D���m�芬KaI�hؕ�7}��;+k�_e�� o2"zH���ٳ���O�{�F����=N^DW\�u�_ta_Sޮ梥�/C�7jhe7��e�maά��+)���r鸩��S�$��{���ᦆ+�[�W�����p:i��V�
�e�]K#,b�۹H	�s�nB�E]���"Q�q�Hp����Hl:�W���Ev���w�"}��^�ٽ[���.�K����̧IY�[�b
ֈ�Cp����읃�y��S��R�Ԡ�<z�$�5nf��3R�*�����]nJ��M����gD��<�ǀ�4M0s�k(��:�bN[;�z�e�p΋���\q7��kEy�eF
�w5�	K���s.u�7����μY4_5���Bi��}]}ϧ<�ظ�7s�0��Y�@R3ueCV2!�fh#S�֩ѭ�i)�9N��;{�}��r�>�]b�fM���'эw׀���Y#��U�KY��IO`�eͷ�Ԫ��|�5�>[��0��]�-=I
���Z����zw������3�亐��af�f�pe��=�/pܡ�7���z݁�bf��vn��2�8�5���y�M�3,5��}��7�+��M��t���rZ�5Y��O���������M�$u�JscΔ���r�l����:�*Wϛ�Ւ.��CP��S+&%d�X�h�,�
���v֫�*=�s�K��K�O_Sh[�`S���ۓ���ܐFn!O:y�%�=Zr�us����2l���4��g�>OMh���wGj$�R�C������8�d�!�D�[dG{�v�L��&�C@�s5wY�4�-�-�
���v�_NR�$��v�e���iQ�5���J��폵ww<��}s�@60V"�3I7��ȲT�f%I1 m�T��E �KAT�d���9J�LLq1"�(���0@�+hTY[r�2[b�%AER
,1*E����i�eB�Tm�YX,���PQ�p@��- P����Pn�V*��ڭK���%J2ڵ��
�B�0���Cd]�1%M[1�V-���mid�L�
��ƭZ�
D��U*���%T*�¤�M!��c\T`��qb��r�lX�f�4��@�%��c+QV,��\����<�]�\oU��0�O��B��s�|W�9�C/��`��r#	F'}�c6˥��"w�S��Y���*����B�S�h�d�֫xV�QB5Ti��$ͱ��.��gVoqj��o.p��*ՌQ[�u�}F�H%��MA-������U�*^e�� ��7}C'R�W�o��}�z����X*�ۥ�;��|�e���'aHY�w�aoW�5~�|N/����5����u�j��?r�a��.9ڢW?�s��y����z�����)���If����{�'1
��4C�5)�f�i�;�#�.�x��uz�^<��C|w�+�T_�������e[��>nn{Aڅ1r,�О���r=%k����k�1֥�`��n����1+�{����E;;}��'�tУ���X��^0�,�˾�a`c8�������>���%zt�h'�&��#���{3���!����QPj;naH펁"ٷ�ǒ��e��i�**W��pP�r#-��\�z�y7��f��q�\yQ	a�~7Z)q`y���X�.��@��$c��R'�^&L�U.6c1���y�{N����z�B��ӭ�i��S=�$�Y�3�ӗ���^���J�)S��+��%,�-C�}�B�܍��i���),\�GN�n�mQ�'�7wv�E�S�lװ�����8�䍝�ue,��r�.}@y#��z3�"����n��3�ʓ��hI�9\�6�=C������2]b�xxc7��8����*OJ�:��;,ky���Uj�C.�<�U�a����e����d�ݽ^�#r��qlD3����u5�s�{�9[���F+���=���a����{��Iw�q�}r*w�R���nv{�"��a��J{ܶͣĖ�G;�<6�|�,���$�.����f�%�ɍ}ӷ'�,EC�G��:�g�&p�y�k��z�!���Y��P��W��oR�}rʎ�$͹n&���msOV���"�l]rLa�i�x�*O�(��=؟a]�8�s}xүn�wy:�,v�f����OT-�h�6Lқuz��[�(2�ۅ�����(W��g�E,7����J��.���i-��]Jʜ��3&l��x0�ݨ�sxP��	Z����U�ܴ�ot:h���P�8��j�����)���#^�kq4q莵��IBظ�yI>�,J�l]>�Y�8�m��c����*�-��P͎�'��m��7��}.�lK�@�z���a���S�o�b��>ո(����:��[E���f�=c��29�؛��ܷ�rb�X������Le��۩�kW2��iӐ�D�p�^��B��{�y�x�n�<T�m�U�����|xɼ��Y��UE��B[ٖ��V�Q�FiԱ3Ǔ��U�5:��Y�Y�&���l���e]����]GF����3=��PS�.�IU��=[4�ؐ՞�H0v^��-Σ��j�7q�ۗi��`��8]�\��\f_r��K��[lΤ�vLe�ιk.r��vgre�ؾ�������g.�a�V�����֭|X�y�w3��"�m�2"�E%�Ό�2������Ik��E�z�Wv�\X�̉�n/Uux0yq�<#F�?z��>[#����(bֺ�l�'�ag�A��&��/7������\c�O�^�c���*&�<�|��O�S�ۖ+8��V�����J�Z��'�5`�9b��p4eଷ��ul\>�90#����SZq���4^W\sY�W=.��^S��j�g��Hm'��]�ɯ��W�kۧ�Ue5���#��z�ٴ��pr|oB.���H��@^)6��
߭�<�
�9	9Q�\)uk]�nI���e�'b�:P����4bV!zv�����w�����Rdl�+
�������v2��K���j5�����R�;�:qO�N���f﫳�X����3�:�g�M�W>EV���w����x�w-�q�4�[�7�e*<�>��7��>��lF:���BC��E��+���v�>J�m�.��}S�;��T�"��I���*k��l*Vͥ �=�0�B�csf%��d�ܵ�9nxf�ˬE3
i�j�V�d^�]��J��NÇ@��k�i�r��xI�a�Gb���͵���"�Փ���ƟR�5rFf��6���Z�X[,P3V�3��.�+��]zS���W��Vв���LGr��H]��N���V���-Fv��ލ�z�_�
a��P�zf��@�.d�,���>���ѻPՑ��8D��s	��#��Ԓ�;��T\pCJ�E,�S�w0��k��l6�}�;=�����8��ԃ����뙽�غvܮ>��
ı�mw9a�wz�� H�Q�J+�q�I��ľ�s�Fmmƴ���cص;7_��Nd�|}�iܥ��@�=J��ʡ��-*��F��v�G7>;+�)O���pW�wR���ţ���Ӽ:��̥w�{�V���^���Osp��n�J�&7Ϫs��tMB�dew6Ү)Vj�n��ٳ�v�mu��Q<��ŋR+%$�����;:�IO�Q{��̝��)���0�����'=�����HD���Wd@@�6uQ-os�ZFw0�m�v�k�����R�V�������V����D�-Jރ�eGa�c��.���"��ń[���Rph�:�è�ׄ�{O��*{�'8���4�K;c-�v�a��������x/��᛺����ܟ:��}�)=��䝾��9��si��;�ɴ}�ѫ����:%ź���f�"-*
8�z��:\����:>'���7��~��=~*+&� N�2���Q�E�C�Ʊ��N��?{v5b8E�D[{~���[�4�rH��춟n8X�vlA;w�6dFk��C%#�.�n���ų��w�V��:�sy���rnŎ�5��v]u��dt�
j��_Y�]�om5�S����,7jV�[�T���hp�T��n��m�+��7��#D��"�c�#����w�v��
�c�2�P�#:���':���3y|��(�Kx��[P����V�,eή�\��eZ+�ZiE�1����u�[%�s�7�R�LE��i�񖬍{���H���/L�����=�0��U.vuE��JB��p��x#�f�n��c
9�B܎�)�D�n�q�t�O�(}�܎���8�5p�󞳨�\t>�=L�tGi��y�Y�S��o�[إ:�2��O8�!^��ͤ;q���+̊!�m�5i�RL�Z���[I��^�t�L��S���f�Ӽ"�SF6������C��<:��։z5 ��b˱+))��ՙ&X�������d]�a�{˗WI�&ˮ\�D�+�+�=͏i/����f�u�ڣ��Ԙ�4������;f�^Yo[���ǥ�/K��U�0�U��\��`�T1�4.�(\���p�;ZGt�X�}�k"�h,�5}"�vA���GI.��n��7�t�u������_>�%!��߽��E������_a\�RW[9(Z���i�=��v斘�Mglrn�ߪgH�K6�7m���geK͚�!*9l�8��k43�RU���]҂��3����V�)��uo�� ��7X�@T�Բ>������9��jy��pA����a�o%�N�br�t�t���$��t��!v�)��eI���j`J�
tޖ~���p89�5�Eԩ�6��:̸��:�;0"��:�]J4��g2C��G*V�Y��P0J��{Eh�X�͞G4j�a�pņ;����f�Q�t�x���`lf,cq��(d�X�lJ�v���y�qfGX�]h�$ݜOMꕉ�u
��d[Ư���s�p1b�ЇGN��]Z��McPm�Ǚ�֍Rq�')#]��>Z�[�Z@ba9��6�l&ՠB!Ѝ��y�U��i��Qx�t��30;��O�N�L���VC�\�2�*�9'`�ٚ�JRl�b��֕]
5��`V�Iƚ��d#{��uڣx��QO��*�p��8�aLE��z1�J'�s�{MN+�
YM`�����J�+n�/x��l�04 �%$ar�����gY{3'm�h��z�WLU�pZ�WjsFP�H*uQ���ջ��oWU�0N�+͹��Ƭ׌���Ss1�I*sg_n���>��z����u�p��5��LD3�:�xq Rٻ\j�_5yl�6���(>[���񌛼�EC��;�x*9SI���$]���ѱ���l��y���:��".�,E�l<��,UA��WD������|��L�9�)�q�;��EX	q���*�	����w��M��rJpvUA�V��7U3�uu�����1�BC����J��+L��7y��&E2�Ǖ���p�ޛ8&QYR����\���f�ɴ�+u���ӏ�9. K��.=�{Xݣ]�GRu�;e�*�d 1�mn��du�]gJٜ;+4��
&�|n��c��p��V��U�ӛQ�b�<Si��5Tv�\Y3n��1K����Mb�Rr̐��ڭ���ܕ��C�ḃ�X�b�Q���2�a��M�ʐ��u�)BY*�k;j�Vv\WM�5����N��U����0�t5,%eUjT++QE+*(�

DdXj�H:�b��%CV�TTX#Z�qSHCBb���,�FTXV����0�Af!�P�T
�kE�Hi�i$�%Imd5���	�Z��J���ƲVJ�B���1HVQ��4�1A0e`�U`�,*[aXL�
���Jʆ�\m�VE�V��R��
ũY1��U�e`c(�$��������k*EX��T�(�E����6�HV���Y���FV���Vjj�H�5�����>�=���ۢ.��s�$C�9;F�&���.�p�	�wQ%�^����3+�� �jJ֦���k�[.����W�*1P�6�^��ӈ{vs�`��J+j]�4�C����=�&w��d:�bt�E��s��*j��u��b8(�K]o�s�ɡ�2;bp�u��͖x:�y�%(�|Q�)�W;��5=�$�v<ԑ�F�u�<����r�5�Ol�踋�j���@ۦ�ESN��J�G-�']f�ȡrs���m *��*�%x����A������qw��s����{q5c�E�gyeQA	���^ff[jؑ�OL��x��J��W���/8��}���+]���}Z�He#;r�s̺�.b�+�:ť���~���1^[c��7��ڮ�٘�BJ6��%�,[{ff�2�Y��9gW�$1Z:��ѵ������d����>;/��^U�>fM�4-!a�
�r�Z{�/�oӢ�0��F�����D��㛬�YW�[sɔzv��u��,����eZ���wG����^j۸��x���ݳ9�]-E'�KW�?M׮��#��f��˹��&��.��k�/z�ܷ ��^��6�t��p�Jtv���:�[�c_>	�ɞ���E�CI�l�ǚ0_N��!�U��C�	#s�jm��"��q5u���2F�M��}�Ǻ�
��+�k��v,�|$8��߻,�w	�O�
�re{�^��ܓo�Sh~b�Y�d#�EM��,L�A+{�iE��<�?���=��Ƴ�M�+��6���d`9E�3v����%�|	¶����m^�Z@9��q
�w�R���:Y�v�S��8���^�_2�a�������$������׳܅�	�Z�Y�LT@/���	�ˡ���~��ݶ�MnME��/i��a�{�����]�}犠qP#5���j��E��)�ʲ���:P�8y���8F�	��OS:�n��ݺJ���$�lq�4a�Y7$�K���v�g����V�y9���4Wb�;�or�K8��-�H�ɢ�{<�䓗�C���W���i�Ɂ�㚆�3f]�|���V�n�@�9�EG���g����	^�m���eV���L�[	���{�m���	B�&�k�3�6V���^�dQ���m�"�` �.�7�6��Z�Yj�B���-u��nS���Jܨ�X����nI�t�Eh�[
wW@㚑YZIn���D��(��UE@���[���v{���HQR:�pa�Q��5�Ŝ��h���kP�zc���i/�'�ާc"njv�oK5���=��yE ��QCUF�S���j˙^�E�1���������SS���(,"QeJ4ݏn�	�b��x��������-�ߠN�Ɵ��f�5�I �mY:J�\\jl�h����Տ-�j�s�qS��C}ɕQ;n����R1����c�:s��������q6��s�у�kѩ竮�;��ol��z�8Y�/�n{�ͣB�+�6 �ON��uM�bU:��jN�M%:u�s�,Vf�Q�O&�!aV�-���`���9��m������I�g�:~y�>�AvZ�k;Uw��L�83�R{��ai�E-P�0*����5��oKOǻu��|srN����}�[�E��R$О���w���)F���v��A����x�o k��|�h�E�ɕ�Ğ�A�{�7u�Y!jP��Rغ䚽Q�*��'���L�4
i�}t���dX��&���S�摌�qo�ꅺr���i�Lϑ�y<�a{.��M&��槎D���"�w�g�>�o*F{R$���/#]�l�Q����\�޿6�o�M;K���O��Y�[�up�׻V� w!N�
Ps��tj�v���<Oj+o5b4�u3k�r�5�Hǹ�Β��BfN��U����2�c��l��W��g
�V|��/�d_ �Q�gW�XO���C�ʳ��Tw�'[(Ɓ}�{1���x��6��+7�+�Rb���S�<�+]�h;+��a�:DoI���f�6�vcq0k&������1��Z���f��O�R���i&x�^���y�֯8�l(�߭��$�M�T౛CwľʹR�!����4�b��<���-Z4"#�x�(J����ek2w��Ի�Wg��~f�8�'�t>x��+��]�K���
����V9cw���u���3.%	�J�g3��&��ѣ���gAQ��b�ӊ�h�L]�ʗ�@�Bz��-��*+9����̻T!Uc��$�|v�~ˊ�͇y>o��U�����ީ�qS}�������׿S+t&/̟
����++�kA���Oۇ���˺unq�=��� �-cPj[�pr��	g��N33�$U�X˺����rD�`�Tt�sM$̽�8��N�W�{�OMB}1U��q7=�=�<���
-����/�|�n�x�$w3����>��\�[n�������L�}�;[�4RY�ڮ��/���7��5��#�ж��U���F�?�o�c0�{k�����m#-�U��i+;�f�� ��G;-ub��$m7�]5tGj�K'w�l��_���/��E�w��@{�ov�);[8S}�]Nw9Ȼ%kG'e!o�dD�Wq�=��v�\�vp��$�����m]^��F�υ�k{2�\r����F্����Oʣֆ���0�u����n�{�~�{uo���ѯ7ћ�Ȗ��ΛƳ��m=��x[s��:�V�Gyӕo��ۻ��[�ܔ帞Wy
�aD�ܮ��iQki���Y��ctS���X�S���\y��DR9����֟{ί�>>@��)AՙaI�ߗ��~-��Hp�:���u�EU�����Ύ�)���]=[vf�uvX��)l�:1DЛo,����n��u����=5!�&��{K���+�n�ޓ{h`Y�Wk<r�DT,å�%Zјؙ������T�^"8�`��^��p�G!d��*�H��R���]� *r���s�u��kO���������
��z��W�_Ya�������osw7��9"1p��ۆ�[ݯ��k|���N&�S�n���?���Z�+z� j}������1+������c��;p�iWQu	��d:o5ߟY��!tW�������I�W�@�̔	OF7�~��J)�e���7/qЙ:��~�~�-��A�56�TH}�;��\�⋢$_<*�c4��6�T@<!9p/Й��WDV�僃c���K���/TU�ڍ.��E�3�-��C�:�gy������#��b������9�nh; ̔�=��;�T��NC�8��rf�l��4��Zº9g�
ੲ=M"��Y٬��٠�Ï�R���q�b�J軀7u$��ߥ��N��ʚ�y�2q7�J+�B)�zQXa�5��t3�6��Ԙ�{%=?S�Y8�W�y���딓n����D�+c��71<Ό�فմu��V�X�p��X�-O�H
C&�$:Y�h�-�i�pޓ3�.r�C��Y�`8do��>b��q%5Û�=;~��O>5f�V����{hҀ-NG[M��Y��l�9cB�J���3���b(��^F(�Q/l�c��*{T<���zꯩf�eK�,`c��ƪ�Y�QW�'b?El�L�U}���=�宀S�,�gϊJ�MX�������>�us5a@��I<��*���=vmv�U	5�|��ʒ�ɏp�Ә��a�Y;�[�I.6z�Qp�r���Iw�u�F&�ܹf����+E��s��޺Q*� �O5�r�PR�uxmq���u)�<���MQ|4M�Y�jћ��*$�td�±J�Y�D�s�8Z�j�R��@2�8ȫX5�4c�"E]�=�"ƺ�ݾ��=��q�:ٙx�]�Q��W'u�TCmgp�U��Xw�Ύ�H�%�U�e����޷آyh:�:�I̳Ri��-�fpB7�ҥAP���N�.���"T1�� ^�>=;�@�荞��<nm�� ��+�[|�B_r�����%�1B�]/Hp)�B[�Di�@�)m�հ��o�ˉY<f�p�0�5��]fV`c�ug(���*��U��B�(r�obS�a7Y�V���w��՚�)�ƪ��j�hmb�ԗ�6��Mν�j�y��b��X�5��Rӽ����A��>+��+�:f�B�����Չ戹��g�a��\��b�A�e��V%J4�Ө��n=c~ػ�xթ}Vn��5r0fk�˷�A�̩̹bweMt�U�m����5�wk ˳���F����E*������`�\ٚ�.O��Sf[j.tWG�n�.:��S�q�ٱ|�W�~U��%	j��U��t��"��90�
�w��ea�o�m��ee�`�nf�4�K{z!M��չl@v����hUݗ�H4�1sw�Բ�2����|	�-�Ήۡ}z9�W���ԙ;44bv�OZ}m����U;��n��Y�W9�9٭vt�*e*%S��G�J�9��0J�CL*'�F�p@���]Z���{]�ʙ(*%��d���ݥ{�� X�b���e]���/$oF����	�$�KNS"��WU����:��㎹�JB,QfZKi%H,
ʒ)Rt��b�H��$�ʄ�(��kjT��C-`�I*T��1�
�T�L\��(��V(�(,� ���R�YFH�T��r�oy1 )���U*Q�
�Q����i�C��� ��`�Q��ek+ڠTP�U*� ZR
ԊUaR-�a\J�B�"ɭXb�4�IRUE�i[iPĹe`TY
¡(T��Rbb9Adm"��*���ɦ�4�LMk+1�Y�P�(��b�����c�u��w[H��XTx�,����5�&a��.6�}��E�oV�qR��_��P,_2��7]�2cI�w�p�nwz���o�VQ[Y�n�#��M�>��x�ꇶ�r'*a���鈜�q�e��W�"*f��M�[�\�������Pk"�slm�x5f6��/���eK�U�M������ޥ����;��B*�U0�EnZ�oM��[���w��4�n�[}Ql��U�3��f��s�3jne�W��z�U�[��N���{LMa��e��i��F�������T�ʑl��r-���v�.oOYc^Iz��֝��Óy�9�WN�Ҏ��ӿhKC�%�ܚ���e�as)%��8���sy�";�I�v����L\#/�if.�����[�ؓ8��X���#�>xޕ��uK7@\E�����x�-U�z#�Pݗ�v#N��k��5s;���ط�U��?N:}������C��b��S�U����笫��c�j#{�hZsϹ;q@^�T��RP���es*�c�w��{>�����8u��낅��g���8�]���� m��\"�5�qTs��5��Kr� �&�GLvp�^��"��3_5є��-$�wϔy\}�+͞�-m�q��|WO7��{���aҷ-���"�k�ݽB�X5˸�ׁ5V�o���j�����N�P���[�}�j�E��E=�}f|�ˌ��3뽭�9]�i���)�P���p�b^+�����hJ��_@���
�������#�ŘË��>p�-!��D;��:¼}����|����+��p�+��3@Vqo.fgV���sU��X��**���!=}����F^���o�%��3�OcXZ����n��
���O��X�����D	44�-�{�������"�z,��צ����<�����N ��T������u� ��G;"���ӝ�������Ur���j�\�/l�ۛ�Ab�(8�=���Z5��v��;�ڳsV]U;Xl4j�$E�}P�ov�G}�)#k=��7\~�C|�'�P"y��+DWp���fL��m��>$��m��r�R�(���9�3W��E{i���;΢l�`V��f��^���Ϥ�V���$���G���KYG�c�V�g�2��v"jm�*|Zu��m�.5�K�{mI�k�睫��p��T����;46��P!��/�0�^���YxKK�1�#��Cb#K�~J(B����i�����b4Ւ'@�e\C�������3��}����\�ػ�T^��>��n�)��k,��׏���-�[P�Ȏʉ�g9e��LЃ�i�<���(y���s�'oγ:�['-������ �z�?^Ԃ��.S{�U/M�M+:[���>�ܢ�)A@�etA�^��� �-�3��p*��2�s�&��>Ze�i�1!��|�4�;�>@J�B����Sx��᜶��� 4���*�Լ��ϴӚ�&�V����`�uBV]��|��$ҬklN���^���L]q!�mD�u'%�.�H��sYד�\s��6\u�Q�wnD�ͽ����U�O^w�bf�@���p���'�j�pv�#�p؝���5���t��Eiv�L��t��k�oWA����|�w*�L�@@��F��F�Y�Ⓙ:P8���rVm:S.ːL��**��e��WF�[�Ǉ\�6M7آ��1[^�S�.շH�.�eS��IԥnU�P6���Yu�)A����9�-���g."�W���!(A����Ȩ5�t9:N+u���[: ��FNJ��]�TdGd_X��>����Ou�&�EH�J��}�m��{q�A��Q�W��_׌�Ѽ����N��)l���)'Z:S@�]��3G�Mno�4�NB�[�3Q��܂k���9'u���R�o�vc��h�M��[���Iԇ[�,S'�����&x9j���[�A���T�s��;��J�`8��ib�t����<��T�eL�_Q���Q���*0Hx�/��]���e3r3��
 <t�#<�FF�2x���}Z���	m��t;f�+zϣs�{vi.S���/s��;�Z ��m������fa�g7��I�Y�y��N�j(v��N��O�J��9�=}}�O�h�u5����ݬu�"�8��3�u��9Q�[�WT�\�ƣ9�5�I�Τ���&�j��]�tgs:�SX�8H�� �70���0*5��tywe�;�8�=z�;�V�����5�U��s8�5�u�d8\�O�yr
�5���ڳbh�$���*6�`�#8�^�w�,vc<��='{b��xF֗�"4�����Xt�����i�y���[Yc�xJq(�c��q�]
l��`��v��L-0���т.SOrC�9�Qǩ��8n���%�Bm���g�c��<�R�)Eԏ��p�5�~�����m͇���*����<Y]�9�Ay�u�-Q���C����鱄���;���
Xv�[(�{��f��hDGr^,´ⳣ��q�̋����1PՕ��x���`�=-(˥�(d�@0����̥�*�3�U��U��ׁj7RR��=���9tԪ��u�������1���*%0=�h��p�:�Ҝ5�h�«}�.�)�$}H(��۬�uK���Mj����z?�v�[ز3�fI��8��GdM\V��o�F��!4<�������%_Y\�Տ-Z]lD�R���U���Q�� o����s�����r㰢_:=��܇�Rי�=�=�=^pQ��{;=(&� �#��׹���U2�͠s�{�O)F�����I�^�픖������Xs���UٸJ�b6n�3�s��WF"�	f���8�]Æ�jHmC�Z��Tnu��u�a�K1s9͊�ѩv��1�tٮC�	x�^�����o|�;x��!�ULT�iG���x
%�ɫG��f
�E�įL�hvP��ƻl¶jl��Uŝne�mjn:�������X�v������l�(5P��fEQ�~T�8��1QhodT������&�B��zU����Ι�� ���h�<ngvru�)�<JI	�t�;��z
9F�76W�ff�^u�<&6���m7�OgL�ʜ�gS�����ǹ�x^��<��oX��y�T�N��p��r6���ȍ;�A�Z`_'��ى������g7|�賣<�Zy��^�$R:�	���/i��]a���7Ǭړ��_����ȳ%f8���`Iov�śe�B�����|�.�����Qb�C�e��=/uX�5'qѾ^U�����rK5m�W���&T�:m�r�#���s.C7\N�^R�gK�bj����κ�6��:�+�2���w�⮎-)�IaΨd��A32�1=�n澲%�|Hb��.��H�wn��^��C4~�*�51־]L���ub�M�Y�Vܞ���V�5[�ym�]��S�s\qrS��DJ��K�U������y�
�u'�х�9t�b�H�����^q2{����4�]��Ӿ	�=a7��3��Y)>>��{�'�,�n��:�����É��6���[X==[p^�:�����-`�o�"��q�֗3�#_n6�apo�p ��2�g� ���FU�;k�Ѧ����2#���{�ܱUG�X��KR��Խ�N���68�e��-՟߯�����u_O��EO����U>�6�@!�?/�I ��
N�I$�RX���aMK32g7�j<_������ׂx'iI��L�k,<�L$� �6XX&�P>xH_�!��A,�Fk�_� p%�X�|��I ��/�����[������>����<�Ԣ&pM��B>��tj!��'Bs�dρ�R��N�[̜����s�f��!$��������������$�I��I$�r ���L>�}_�:��|
P�C��~p?��O�_���Y�Mϰ>3�>���@!�������`����`r�$2B>قC�������p�iM�����[��đ��}'���X19�����q�f����,	$�A:>�e�F�.�lD����@!{�}Ρ'�ڬ�	f6��\����a�ܟG��SG��I �Ić*�O��?)>�������'���?�@�.��;�����>$7�>F����~G�d��?�������>iBI$�	dg���C�p}�?�I��0>��ÃAO�O�8��	�B�d����}�����϶.��r��t�:��g�I�N?p}ߡ��O���$�}�F=}_��"�P��p��nt"�
��}�@�-!��	 �&O��@!����);g�d?�H}&]�Ĕ>$���Ѱ�C�nI��p|p |�X ��d��RD?������d�I�r}'�I�k���<�2�%���	��@�'K?8	1��;����:���6BI �`}��~�y}2PI �����X�D>S��	>������'���y�>?Ğ����� �����'��#�!�!��>���������g��C_���!�k��P$�����#���_���O��2A��I$O���S��'������	�g�� |'�	�ć����<��d��!�?-"!��C�>"M���I�~��p����?y�O�~���d9'g��7����`I$}�a'�I�5�?W��~�C�?>B��s���[�ρN~�/�Ѳ�P��n��� �I$��~�'�L��}O�??��N����I$i>���8&����Rq7��)'Q��s���3g>0X�2�	�%�?O�	��s?�.�p�!.��