BZh91AY&SY]�lR��_�@q���#� ����bD�� �
        �}�*��A * ������0J��E%T)h�) �
UP%J%�$UQEH�dkZR��ĕT:�IGYHT��%T�f�Х%m��mDJTE)5�"kQ
B� *�%(UQB�N*�yȥH��N .�*u��N 1���ȅ��T
K�PR���U*�f�R�E
�T��UT$��%Ze��C`���@�QT�����:�W����3��cM��(���ˮ�� �����@�;w����뫀k;gm]�S����{��Ν�
K���)$�����e
Gϔ� ��|ת��Eܷz��(����
X�{�`�RTc�t:eJr�OTDRw�o{TPU/����ZR����������J��©��z�*�F����TD*\�|�(� �=�Щ%���R����E$(	Ǽ���ڥ�Wz�TK��=瞕@
=�{��(�{Ă�R���xk�*��{���}��R6�����T�m�u�H�'Ϥ� �>������{m�I
U]y���IT�zށ��m���C��*T�����B�e���TU{�΅(EBg=��"��{�c�ID�A��"@��k2�$�

�/�JH ;���
B��wA*�t��*AR�wM�=QT)׳{�ZUouJ$%Ct�v�Un+�R�,��yR�I���OT(w@��ٓ�6h�fy��/� �R|s�]j%c�۵ւ�ll����

T�u��R�*rX�TU*��;�J(*5��T��ۛ��GF�kO�� ����h[S�RSϔ� �{� ��	���$ g]��@ A�� �p�� ��W���P���(ۭ\ aV؈UK� 
�O}$ �����0 (�uW G:0v8� wJ�( 0��� <׸ t:` n�Pn��i�6�jTP�c�H ޽�^�� tt� ��A:���@z�(��/q��=��@ ���  g P�j����*���I�P�>�J@�|�u�  �\�x�,G� c��b` r[p �� \�]�@�  <|  )"��B�  ��2R�H�ML �0Fɀ��1)** �4� �5=1%T�Q�      j��&��(� с20M4�����% ��A���  "6��F)��� L(�z�m��������TFF��ї�S�����������B��jK�s�y�N3�g�u�s� U�ʨ�@S�
�*��芀��h�������������(��T���� �A�u$�O��iP U��?��S��
(��O��_þ��L_���-�m�Č[`�ض��-�m�[�61m�[ض��l[b���0m�lbŶ-�m�[ضŌ�l[b�ض6Ŧ-�K`F%�`Ŷ-�m�[ �-��`�؅�m�[ �-�m�1-�L��m�[ �	l[a��-�[؅�b�#-�lإ�bŶ!lal���-�[�-�`�1-�[�	lB؅�`Ŧ�)�[ �	lBض�-�l���^ʽ�{-��W��ͽ�ض�-�[��`�b��lB�%�`��-�lŶ)l��b�-�[���-�b��!lBضŶ-2؅0`Ŷl��`��b[ �l[`�Ŷ	l[al�-�lB��b6Ķ$`Ŷ-�b� �l�b�-�[���e^�^ʽ����oeVŶ-�`����[`��-�b�ض�-�l#m,b�ضŶ-�m�l[`��K`Ŷ�m�[؅��[��m�[ �-�alH�-�l[`���m�l�60`�ضŶ�`� �!l�[b�ؖ�-�l`�ضČ�-�-�lضŶ!l[b��Sش�-�l[`�-�l�6���JbŶ-�b��-�1-�lb��6�-�[���b�ضŶ-�m�l[`�ؖĶ1��lKb��6Ķ-�m�l[`��6Ŷ�-��lض���m�l�6��-���
b�ض�-�l؅�-�0m�SضŶl[`��!m4��)�[��b�؅�m�Lm�L�6Ŷl��m�le�
`� �l�6�-�[ �L�LBض�-�[�l[`�-�lX�b�-�[ �!l��K`��,bSإ1Kb�m�[�1-�S�!lB؅�m�[�1�lB��b�-�[�%1-���	l�%�Kb��%1K`��m��-�l[b�)�lZ`�ؖ��-�-�lQ#ت���(���%�T-�!l`�[؂�cآ����-��l`[R؈��#[b [[b�[B� ���-��l#؂�@�"�-�	lEKb [�
�ؔ�V؂�V� ��*��-��l`��[� �@�
�-�l` [[`�lm���1�"�� � �-��l b [ت� ،b0@�*0U� ��E� ���E��-�l �m���@-�lb([ Bآ��(��b[آ�@� ��-��lD`[ 0B؂��T�
��D-��lK`
[B����*[ �!l[b� �!lb�# �-�`��-�b���0b�ضŶl��m�lc�6Ŷl��m�l�lH�-�[ �-�b�ضŶ-��6���m�l`Ŷ-�0m�[ �-�`� �-�m���-�l��`��,b��%�m�X�-�lb�-�S �-�b��-�m�[ �-�b��6Ŷ�b�`[ �l[bŶ-�m�[Ķ!l[b[�6Ŷ-�m�lX���`�-�lb���cm-�m�l`����T�����H��h�����zL��N�}�
�|V�u�qњT
�ݛn����d�:��c�y���,�T��{vG�M7�M�ѡ���uy�dp��I���A`� �����E�@a�0Zz�j�<f�'1^�0ըe����T�\�PӁ��盶^�jYoo�v��Ӕ�_�h!X�Z����N�����I l
�֓��eBVm�N�[���3^n�A�D*��*Q�v'��OQf�����wz�)Q��o#�C��]I�LP���-n��Hp[�0��[e��r��k��5ff�E��-+��gD��4�^�2�/^C�`�LBEo�a�DV[[���4�Pp�$���T�;��V���z兦Z4��%�`'/owr��TD�J�x�u�V�I3(2��t@���t��j�YOFzS���Vl��Q�Z�<E��g��Xlcs
1�^'[��-PjA�e�z}�sn�Q��N-�Gr�[YR*,T����.S�Lo)����P��vf��~�M���&*��\����m�1N��׭Isc�NeJ��ե5��*m!u6�X���9���"�W� �� q�D��Wv.87r���.�]޻R�U��Q�5#j3OG��E�6]�Ӯb��ucLup*h<"���M'H%pfƴ,v5eU����!��˛�M��ä�i��1���7HݭMaT�/mˑ�ܤI�7~M-Ԟ�d�7 ؠ�����h;�mM�u���eS�+�"e�k�j��f�z�3%7�����X{Ugb��sn�#�&X�M�%�#5�
��(�
�'baV��/�l����zP1Rn�8#�)��J�i)2r�e_dyy1a0;��Ñ���d=N��m�pQ���ɣ)��3^)*��#�J<�l~�QZة�.�����t�f���2c�;�Yv�:Trk��fs�r�8������"MPv-�у�z(ᜊ�����ͪtD�VqЍ���(j�<�j�N��st\��ں��<�w��s��덌���*�;N^
�3)���NĶ��	�{t�P9�����"6T�+2�G
��&�re���B��n�\��P�b^CC[U���2�2Ƽ�,���*�^^�{1�VV��:!ů+�3U=�a9J�[ebn�-Q��dX�5N\ʚ4�c*��/ ]����oV@н��a�u8��N[(jÒ'MX$�9��B^#`MGQ�����Ӫ�S�az�e�60�siK+��U��8LKh�ӊ�Y��I*�
J:t�3��2�#�	�a�ҝ�����R��Z+l ���+��1t�4Όn�+�7$f�&]��j�������ӵ��V�塋V��T���A��rG�Y��36�k�F��,�Kv�nF��.����Kp��m�l���t�k0aa[���c��X��`�v�I����QQ�M�`J�ENar���i:%�u��F�ɗFm�O�1kU���*
�j�X8�l�g$É�:-V���v�:\���N�*5X�o
h+M��� �b��V�kB�$�/q
�E��SV��g2��v��O�:�{�.�FUՑ��5P[�q;�5my)�ZY��'ɒ�"D��K�<�7i(���Շ��嚬6Rǆ�X^���n�V."Dp�'7mm�;��E��H�)�J��+*�%\I�5c�SW�&�,a�yu7]�Y��w_�L���x���1U�dF��k`����Ś��#�����h��w&��]ed� "�F�4)�B	��t������rm3n��M�T�d᫧gv��4V����nI�r��k
u�x\�.������eޜM%��XС`�i7�[�S�!� q�[��]�2ec�~�VA�yY�EI��V���]�X��*K&m�6T�b���Ԫ0!t�X<y���A޾7{���C[O*�H�d<y���c�Z�ݍ�*��)��֪�װ5B�]]���̵QzH/k%�ڛN�mf��0�^ڵn�Ӕ[ЬlóD��F٘��.�E��U�cD�+u�p3�m����<35Y�|��v���IQ�)����򧈡�<���Ց�&�����FTe�ukz)���hB�R�w@�ǕL�n�f�]�ܒ���M?!���1��l/	ܻ(V
���̍3�\b�ħt��Z0�J̊��<��'*�.�SL��np���������v3GY�Az�� ˣ(��2ʷ�(2���Pf�T��0YS-�R6���
x�h6�q���=�j8���=�i$��ˆC��ͻ[��H�f�-+)��(���9"��2"�[�-��/W��r�kZ6V�v�l���N��5��e�с�(����Y�U%��b�A�n\�h:�P9��4궀V"b�$n`�5~�,ɯ"���iU�q״YD�.%��#S&0�cĥ,�W��HK�Yem <���8��B�&���M������mArH����N7�oK�<f�kf'�m�6�J���x�^]X�(�b���{�� ;su�E5����B�Yz�1
B��sojQ��i�FE�`'W�1J�X�O�:ޖUYJ�wt��K��ѹV�
�k$���.Y�hP�-e���sv��WWSa4�+�p(pQ���a��!t��lu�鰐�5�F�X�e���K��K��e.���uvI:زB��QkhnÔ㡘��[��a�ճkU,�	N]�N]��Ҳ��ic���Q2:Z|vŗ��;�m ��X���a�r��U̫М`�V]j��t&C�z�^��e��(�fH���V�P�n*GnTƚE�Hai �T�v��S&L�3(��Cˍޢ�<�m]�h�f��f���v^��J�y���l���]��z����f��pZ�t�y�y�3D�R�x2�˽�%�I�Ed��7k��L3i����&ǱÛX2�����N�Zz�6�n6�^nG*��&)�mi�w��n:C6�9!��c1P�J�4�D���^�d�Xe�	��f�H�4�J���vXY���ȧ(��4��6���3u�1�˸�� ܦ�m��(Fb�bׄmkc�s8��c���˙FI��L3I�nx�.MG)�6�;��oQ�B�)�7mZ̬�չM�3/ ��k]Kaz��Yp�w��ᔝaۘռr�
od��Xۆ� ��cI�g`��(S8ٳ�lU������ȣ#4V�� ѕ#�M�,Yře���3��ȭ��R���MU�]�&��MCE]�#��z-*d������y��K#"��46��Q6���yU���ují�����c�B�a)y�=y�m�{�+��=ƙ�'T�Z�-i"+�#lF��{�+K[7��]Zl\�shW%�rE,ޓFa�AZ��u���ͭ�j�5���av�i#YI�v�6�[Ba�5�f�tʵ�(�L[NW�ˬ�����ر7e�E^�Nf�˷m��Ct�Q��.��Ed	Rfb��R��)�W���gэ�9&	v�VU�mV:aCi����j�W�٬eMڨ�{*U���B���Õ�&�u�Y�v�!�pޘ&�4I�Ri��4�M<�Q�����-�L����#���,�X���0���B�	a-�`���z3ٰԥ�[��J�"��٫:o5X��6�L�W[�CEn�G$R��� ې�]%{qY��(�[��v/)a���Ѡ�`�Vm�E�b�!Y�)�b�.F�K:�Z��#����:"��
KS��V��D<8�&��
hXe���.��Ki�dʭ�JF��̺�n��bLLL���%�&���d��8��4S�0�Uz,�!��mm�V"Gur���,�icrj�U�h�"2���U�bzSÚR�B 2�w7wv�B������I0�1P��S�Xrc2�
�,<��� ��V��7�m?2��5�wVN���+$i�B�-h ��Y�A��Y�(j�˰f�"y��-+�������Z:-֘�h�����2��� �Y�&^�dVC$R,���(��[`-s%J����Xų���o�Z������)�p;U��(Ě �vRw(�b�f�(�Cͷ1�V�%fM�s)���N���YgV�h�GUdU p�/|���N������G]�(�v5�6I�md���O(��"�w��I�ܔ�s�V;Wx�l[Qj��%m+X�z+3v�E^<��i�X���Ϯb[�u/�%!TF:��<9r��Ǹ�`��,]�UI�Q��A�ɶ�*r�&UY�D��2����A�ɪ��i)jQ�VhS`��ݩ$Z�Ѥ*�;�܊\��9�r�:�w6�X#M%���Oe˛vJW��,�%�U�h�{W��lk��E��m��~́��N��\�R��F�)��e`5ZUʲ-d֖�GA�j'[�26/Br4���7��n��GD�5�0�:���uVL�a����6�+�.�m�%1kl��W�&�5�����*Dm^$"fJݛ�+��J�oM[�CV�L��3y�G��N� �0��%�u6��J�YF�wwtRdSʷx�(�iۉ)*��ʴ�շCL��ySu��*P&���kn�5`YB�XK�X�4�!y�v���kJ��5���N�s&Ԍ��u]Jz�V�`��T�嶖�N��9x�re�Sp�l:�L���w4V4�%�n�G6�bY�G��N��IҖ*�;���V�o����*�����'��1qQ�am�E[V��2��xqҢTW�6�چ3��.���wv��r���\+"���q��X]������[jXM^ܨ젃y�v�TrE-{Sv�EW�;��L�]1�K#iʥ�)#���2#WcIÇA.öD�q���qV-h/:���L=rCV`Ifb1�z�bc�U�-�2TUR��,\���`� �B�w��*�eV7��hZ�T.K8ܘ�aڻ��I=-�U��6�;tFZ�l4v��j5J��u�6��Xw�E�kki�n��5V��.�o.��l���nQ˭T1�.���4���yW,jŒ�J4�C���2T�ܵ�gL]�Y�;�fT��T��eꊎ%6���q�VU�ݒ�6h#K[*֬	G�v8�v�m��늉�O([LV[�RR�n�=�n�؂~��bJ�lZ�7wka��7G4��������%�LdRn@f彷&�b��t�,��4��t'W*eЗu���Ζ�A�(2(�OZл� �������(��ib�e�eS��K�;%���x�9vfhȖ����+<��O&m�E۰`�6ṳ}q�v*���V
&-��!k%�����D�hT̓���֬�+P����e"m�"Q�q�8�'i'uV	x0"��M\Nf�����U�(�t��i�Ũ�n�n팼-�$ҀC�F�#voq��Z9��9�fe4K�n����D��|�3 �Z�~��[�S3k@	�Y
A�4���=ӵO[1@�T���<�kZ��6��,z��e��4�����թ;"���B*�i+5�Q��L\T����f�ъ�ޭ����H߭h;%�Z��JKc���`���H��v:���ҕ�eY`^�nц�Ycb!�Yn�B�c�Unڈ�c�����㥈-�빷z.�����zi
�4̛Rդ;F�6�%w���LZaP�ݣ��a5���Ya�ZY�ġ��n�lG7@t���*�&T� �E�k4ܔ�M��o��	Y1ŹQ�gh����ˡe� ڈM&�fK)�T��ʗ+E˽f�-#�N\9@a���ҭz�����L�[�jM	�gJ�ޠ�+�/D�����A�U�Ҧ�YN҇m��j��sR������FguFoY�pw<��)RR�T$#�ג��#��?J�T�v��.`�+Z��B�w4����ǡb��\�)�-&�&���D�W2�!G)*F��Q����dT
J���4m[B�ڴ�q9�ڷG��N,��-+T�z�v��=����h���`î� 檤	9Ҥ�J)S�)�u�RTTv\"v4�K��#�=�|�N$y��+)��51H�	����T�-�e*�%��J�uw8�36��0F��5%s��� o6���ks#�x�WN�!:�]GAt�OKl;O���ׁ���԰�rں#�/h;�ڴ> k��$�S�a�������ڴ�%��[F�HQX�dArZ7�ϝP:��W��%���p�F�D�#��_&Di[7��b�PG��\�	�;�i L�	Ԛk�_-%��ЗKy5�+IY/�������V��bND�MrH*��I"B�"���"�b�hܜ�2�j5���i(�TBY:���1n$o��餖%����M�K�
5i$�✻E�P'J=x]%E�\B�iR�!�j�M$�\�V�&�Ė���b��
F��:���A�D[��N��"��Q��H͵�r����3���<H;I[	+��ڸ�%�,�
�_Y�_;j¸��5a' �{�������[��wU�xwv�ݥH�\V���Mp�����A�#��RK����V�I���x�&*Yw��%I'W���Ֆ�\͊�&b��⒵2��㥆��
�}V�I]�����KT����S�4��T�;KU�)����W�U���w8,V낙�r.tZ��a�@�s*�a�$�+p�����@���2�T-+���pJS�I�X%"6��'_g-�x�"�4q(�:��ZثP$�a���DLT���#'i6�e6A�wln!��u�B�(��1A2�"�'��x�Iq4��4�Z��ȳ�5ql[���y�����b��YUN2w*,It,UNII x�ԭ.a�_3)�4�N��Ydaw�-9���eӦ$�C��ir%1,X�Ʈ�p2mRؖ��{�e�H�܁b`�R��V��n�Unr-�pe�����_a��� ?_���z~�)��͢����C~&��7I"b��H;�t��w^RuE���[ft���sYF������㧪��U��DS��7(�5v3y����L���%*vE(���K]Cj���KI�.�N�0�I_Vp�+��T��ve;�`fR�[P�N�*2U�ṁVD�nW$J�oL�WN�{�Oz�\�Y�����{I���J���Ԍ�]��3��J���Ë�o�kh�T����"�W w2�o�-m���o��0��5�N���p.�5s�y�\�f��RR���p�׏@3J�"kH�.޺�'a�侻�����R�K=���J�o��In������n�wLz�>�#;���ˁer{����t�-�Te �}��d����kXQ��zۧ��V��V׺��̋w}�>��hFM�Z�)+�gj��L\Ùt�JOw��Mv�~�[��������yM���|:���H�<[����b��Nz�2t&����9�:C-ִ��Q�ۇ�e�wZ�1���2���>Wy�T(��S�
̋N����yM_T�k�ؾ�U�,�u�?$����l��*�6���a��k����;�B����ҽ���[2��hL��Q3����d�~�u �b_�}S�c/Y��}�󮫱����Υ[Ԯf�׭$g7�j�8ց�y�ݝ;u��Y�ܨn�E�ZJS��zf[-�;��]U`�Ҙ���qx�(�ܾ�bF�lT)5�C���]����V��f��K
|�kNF�^�x3E-w^�w��9��oA�1��صG�x���� Yq��;�i;Ԩ3�O:�z��t:�'��AG�5�(1ǌ�ҁ�/�h�F�&r�6��s�ܰ�$���XrG��ݥp�A};M�r=_i��՚|�%�I�l]rj��$�i�*;\��}X;��o׫g������ۻ�]��uq��.��d��l۩�d�s���f-�Y��������AՑΥM��qa�[��I�)��
Z����{/���m�s*Z�����A�H��<8�3����sD^����~���Ԓ��,ש�C�@���ݰz�*ص�SY�[Ըn��
Q<�[T]aT�4۹"w��:j:���eD^-�ǂ�a�S&�Lي�՘òS��n9�l�a���le��k��7�E���
<���ՁYG�����3�����*�xa��8Rc7a|�5Y����%���t�"�,�m��w�
(�=����Q��_Y]W\*f�KqI��s_�w���_^�o�2�Q@������8]�!i��|��)X�ڈ�3B��/M�e�=u�դ���o���I-�Suv�`�SX�k���ӫ6dR1��f���X����-�>a��M���F��2�ov�Y�y�}��J�W%�)��9I��W153��Y�����=��<j�8����Vsq����)����*ݻB�76�2����J�V��v��-�vV���8�]-ۣ��v4{k�=g��*)yY�NKS�����d���&3�Is5W)Z�!7��x{�N16�/���C̝��*���ڑ�z��{������f��N�R��ojċá�b�f�hhV{,t�'W
�����*���V]�u���};�v�3�x��[�8�\-�u�y��ef�fΧl]�:*;��B�ެ��)�Q�=#�+���/Y�[�qގU��',A��&�H�f�j�S��h��Ж��6�P85H���襍��t����M'�	�Lv�Z-S�/�N�Ꝼj�}
7F"������l�Z�K6fp�B��Eq�%�������.*���F�M���a��2=�q�m��<4�+��{VT\+[4`�ՊNoO><%�;�iI��t(�bc����R�(��yt����J�f��g>�Csf���:{f��:ml�$�cRwWQ����"���0,�jkn�x�/N�ZP5�8�;wj�㬫]P�o��z_[�1.˽�t�j5�Z:]f�ޯ25��F��\��oe_t�wnvr�ڎ�VF�k[�ݢ�2�������u)��:�+��:���c$��Sc�ۜ:H����z������ �%�����}��ǅ��!q�:�/�Mm���c���=wb��(���Z�}�_�Z�}��[�6Xj�}�.���ϊɱA-����`pVE�W�!ډ�ݳ����9^����9�����BT�WF;B9�*��3X�+q �bf�kR%"��HN�}"�\�6g�\�(���ü˾l��j�L�m�����*��zt�wĹi�������m��j�&(�^����e3oK��j�[�Y|B�Q��<ĝ�N@��t�qX�Es����,`���(*��j����}�'�co���nK���pǁ<N��-Z�v�5ńU���n>׭υZ)Z���g]2(2�]���!j)b��f��ο/(�FQ�3i_&�=C��¶�RZ�v�u�9R�:��Ww��):�R��mŭ��"��V��*�q���w�.�2�G[+�����K�O �-�5)�۫�z���9Dؼ�X����!w�<�,J���U,I{@M�/cO.�kn��#+�R�I��;#c�r��H��a���tyK��5.�����
o�>3Cξ�̽��X�zs�H7z�(c�ㅾ$a�Pv6U��jq�sF�G8���%$#��[��*��3�;ok+:f#j��E0 E]��.J�+��8f�i�n��.�ե�y�:�L�60ݡ��;����#cy�e-X�9�*��/�Nс�@�k'L���[��J5�N�]�yչ.$4*��	⥨�|�U���@���[~�s'|������񢩝!_?J���Sez.��j��bg^�9�ߦ�X71[/llti��G*����1;ck�c�F��]�Up��]�Hκ��Ն�6w�lAX��,5ͮ��_a2���8�v\��źF�h�dc�cp6��{�z�o�i,�#����׋\���챸��H,��נj�w�iAg�{�i�8�6�j@�\���e�.��J�9�\�nv+W����o�=q�z+����L�X�ص���Q8�Zo}}�����3C��7\��N<�����e�ܬo�C�V�C }���mhY�����dJn��X|�Ge�g�!nWvUͦ� ����)�e�zᴺyAm��Q�|�L�!�Vc��xC�u4��d�{��ӝuo^��=�FDו�yZ��9ێ���b����K'�F�T>��݋\\�[�YY�����IK�L��I��`�$h��u5�쩡�2�s7HZ'b�)�P.�׃i�[Z�N�7�e����"�6$sJ�u��VRp	�j�䵛��x���pt�uԍvM������QG�*�O8J�U��5p��k2�eb�j30���a�US�+�S�^7j@�j�c�u[86�R�̩�	p�x��ViT��9������[�V��N��_>Z�vΝ���\�b�V����Q�&ˎ�V�H�+D�kc;���/h�� =��t��aT�/7�T�.s}��"��p�2y��l��w{=Q_bb�g�u`î�(���e<`�v���Ҭ>\H�=n=G��	���U#��MTG-��jf�>�X�%jr�Y6����u��G8w��Vˤ;G-��_d�]
�eG���ᗑ�mj��,eN�UFZ��!�7�j�$8Q�tO���ik��+�P�]Ë]�-#�T�̛;�n5w�c��2���vhMt��G2�`x���6vڹd4Beoם�e1�Ih�efuL���]�Nyx� ����$6�|7p;�7�Q�Ni�1��Qw`������]��ma���6%$.8k_N	����:.�u��ո+{gl�U�G��w�MW�}��;:�|�@�%`b7�u����k�ꪝD�˺L]>"f���ɯ�c
�R[g����]y/F��,�mR̼c^�)WWiL�O]b�����Z�)�<���ʓgф��/�η̻�Շ=�U��f�����+��P����3���e�w��(��ɾknSћ]m-���to3Xjx�z��Ύ�p��O:�D�c���֝��vq��G$j&h����Ǩ�T�80����i���kz��u�
b!����l��Z��\#4ue�UuݱX��t\5����ԥ��:��!Z���R����fo\�\�b�'~icҁ�Sg2�w����R��|[�v�w]L���N��5�T��e��9w��gV E���+ 9l/E:��֝�BZKS��ם�h;��LB�Y9�6>���e6�{d��	��_ ��5{��{M��J����� �:��0�6��A���ǈ����rP͇mP�&�룔;8=Wعқ*�G.ʒ��b�;����r��d1՞��8�v��vY���W^�ƟS�]ֆ\�,m݂�[���(n��!�4="�Hv�W�lR�wEA�8u��� Xw(�z,�ݣ��dU�5������Ν�t�g`��;�C��,��Jd%�9�Y}Θ�Z�X]Oq\Z0fW�;�Zo�����$WI*�4󺺬��K��z�mbm��iq5E;��f�\bV�*&;^@z��nbF
�w��a�=�;o��yoJ�%�ӱP;�6�{�\��r���Po8u�m]D���6:J���X��ψm�Y�P��_���)�|^e��R�CA50j̱����oC˧���{rl�cgC++���r;;zoj[b�S���d��m�>����6���L��c�7�V5F�Ï��kH�v��K��5���. ����}%�e�cO'O��@��0�![8�����G6�9�OV�;�wi�,��d�wV����ȋ����{쫵S6i�����Эm�6�R��/4X;�ݣ]����*Jt��M9ٿ.��"��1�_��Y�!�N(q#�i���M�qպO��[�+�)>9��}|���Evf꽫���A�"�n�R~E�.��۬��<�k��ɞ��M�cf�w��RoI��U��o.��!Nɸ�r{6{�WfJ�⣗sQ����C�Q��;�8��a��H�*l��Ǎ���m���U�P�y�Wmܻ���������(u5�IQ�[ka�̺޼μ݆�s�Tcn]ku��{�)pC5e�ib��w�����tFc[���Gn�ͧΑ��C��[q���(*�r��&�D�c���=mZ4�ʏta
SS4]	5Z3he��3�gKɗ�Z*��E��ygA&P�J2�=���ıi�5Á�4)ґV�5�dn��Y��i7p*������*���N0*6eqٹ�<�[2��U���ȅ��0N�Bu�/�;$%d�<�2���)z�ZM�Ōgw	������J����������w�t�D�R�%E���&�8q
�k���,vq���1��]P��v�2b��S�C9�WiN
��<�xF칍�՗����bb�'�%��Q��\E�T�X�E�G)ͫB�d�Pfo��yl{Jb�U��*���Nu��; �aD�+U(�̌���]}>_8��ϰ�Pa;o+�rZ�������^��V�痛1Bۼ: u�E+M%YW{O5�=ѥy��m�({���.齨rK��`�%�eD�XR��A%p̺�_Ws�19�O�γdڛr�����Kz���kYGZ���/Ɠ��n�r���j�����1�2�nۗ�����s5s�k�ٌ`��z6�:��o��^Ζ��jć����ui���`Д|	!Sr����ϵ�__{:��՘e��Y}���*�U�,[(�V�W�k���\�E܊�
��)����:S�`���{���UI����pCvĪ�S4��h>��ʾ�K��9���o*��Ke.���DЦ�;O39w�P�Ժv��_T�������+�K�`�E�>��u�}��z�8��Me�KW@�l6��$��a$�I15ó�y��ȍHC.2Y�8Na̵x�`�e޽�3U c'L'*��	T(Q�!��q�ި�Rp;??�L�-�V(����E�X�a��i9)H�Y��Z�_*W0"��$.|ّ�S)"䃔37��S/o��p(n$�"��1CV9�&t��%�m��2!E�@��V�+Un��iی(�p3��P�&Q���Ad$ƣ(%VeU��,�� TB,6��ʞ���$���s��$�'��X����FA��7"�f�����4��f�f�5)P��L�B��,�B���R�9bFc8���l��X�D�55t*�`j�6�tPn��8��[ �UTA".=��2ɺ"��q��t�Mo,���H�S�ٛ��` [N,P�D=:ڈ�BX8�W0i�H�!E&������Ya�K��3IG���D\�	?��`�#1�
�aE��h<���,$,��-@j��	1���b�@��F�G)]Q�(:MșL�\�ɢ/���O`��C3=ct�M�2S�|@@�
�aƸ�5T-��_+![$�R?	1��
U�AI�QF�%���q%m�a���XD�\+8����6�fY8I�Qa�D?SO����9��)!�(�l�I$qIt��+"�J2JI�!JFU��vs/f��l%\�!.�J�eמj��������Ѐ��~�gۿ^�����TDH��_����~�~�����5��>��7�yϾJ!/~P�kI��d:m9���(Y�$�FY��r(�YU�V���@����&�m�Eہ�����wv�1�zY�ڼ���SH�ܕ&���}�F���(ѣ�f5@^�g��c1nٍ]e���uˉeR�����W��������n���s����\V>Yw,z��T����:ڶԻ�J������WRG6n��H���a��Xh��5mSz������x��$�ls�:��GBr���v���5%n��yy�ҡ�z�4ņ7�]�3 Rm��U�K�K���ihb�T]]�S��N��u݂p�9��<���$�]=�r�ʝ0h_RTzFS��+����4�g�{;��N�Br�P��9*�G�H�q֜�)�j��j�p��3%wfN,�L�Q��X����������ڙ�!m�n�l�qJ����S�[�Xr��CK�}y�.�<	���͝�JC����k�h���N�if��#���yŧO^k����sa��f��z�q�Flވ��ޭй�����t�2u�@�#��:���l�������c�[)���#thݘ�����ӵ��;&PU���osx>Η�K!v�T�1�GOx�������z{��8��8�8��8�8��q�n8�q�qǎ�q���<q�8�8��qӎ8�n8�8��q�q�x�q�q�x��8�8�8�q�qǎ8�q�qǎ8�8�q�q�8��6�c�8�4�8�>��q�q�x�4㏎8㎝:q۷���8��q�n8�:q�qێ1�q�qノ8�8��o6r��7��5�+k%���v�6UW��W�:�ݘKVZ�w�9�k�Ghy��f�`"��h�^���+.�>���-$�ɮ6��Ql�YU���u���WM^lL��r��z��i[���c]��	0�V^r�;3$�BWgS��r�`�|eЬ�ΜV�D���1"$�.�g�w���'=�i����!|��ge�.=�]���=�b�Tʼ�>ĥ��� i�O���(uBwc{���������=����8I��=�#��-ǘѾ�"���0����� �E%CKD.M�Kr޲��3�Hv(�r�$�A��b=f���m��o"�RYu���m+�8��_]k���SV��t��սg%J<�ڼ�"�u�֩DpX͹Yݳ��]��op����N�̇���'��$�}=2�Ewuu���u��u�ƨ\y�-�J��+�]��bSQ�+���i��+k'w!x|�hPh��]�W]s����G]�����K��{n���+.�vѺ��HfF�-��'wj	}+�Nyg#�h]c�dv����0�9)a��`�P)ˑ�ĝ*=ݫ6V�Ԁ�X��)w��p-ɕ];{�0PS#���.�4���V�,�UG(�O��Y��=��ǎ�v���z㏮8�N8�8�냎8�8��4�8��q�8�8�8㏮8�8�<q�8�q�}qƜx�8��qӎ8㎜q�v�8ێ8�>8�8�q�N8�:q�qێ8㎜q�v�4�8�>�8�Zq��q�t�8�q�8�8��q�N8�:t�ӧ�8�8��8�8㏎8�oc�8��q�n8㍸�{�%˚o��t���v�b�i���8�÷���҅v�c���M@~PY��m��Goѐ�(��,3y gZƇ�m�u0@�rXj�dԤc�ᰄ���Sqߜ���x��z^�N�j��֥<�ɏj�P�{j��&C�0�k�~���pl]X���]�&����.���{,����f��T�5�F��H_��}om��[ Y��ਔ�b�>X�����p��z�r��*Zcg_kJ�{�2�]�v�>�;(��bv��L�WT�����<�v����mھ��{���R*�3���m�jN�Vm���gqc���񪎆�V�˭�{��5��e�fB��V�U`b�Zwq��-m��-��6���U=��.3u}�j�p�Q�[�Q��R[���]�K(�B�⃨IVel���}R��X�C�M�1T�F:,{�[��](�ẕd�]5��=u�p�n&��WӲw]�^i}Oz�&ni/R�'(�0�t7�ep��I
��јc۷���V�e�����wz���՜��Xe�%�6�3-�	�DoL)�!s̀�r��գ�'U�'qA���+^a�%��oj��8�d\����DO��

ڶi*�Xy"o=��^��7��^;t���q�N4�8��x�q�q�q���q�q��q�q�n8㎜qƜq�q��q�q�pq�q�q�q�q�}qƜq�q��8��q�q�x�q�q�\q�q�q��i�q�N8�;q�i�8�q�q�8�q�q�8�q�q�8�۷n���q�q�88�8�8ノ8�8��4�9��{�~�w�������z��Y��Ud���_i�p�n�<3Z��yf�C�gl��%,�P-ԻUcK��It�H�W�һu��G�♥�=e[�/���Fvu�#*�>�J��m�c��.�OhT��ǥ�6���G��C��W]��͑8f��x��}םkD��}HBڼ��| 1��Yڷr��s�S���M�/2�I�he	��n�U�9�9}L��a���6�c��mj����dR��lAe��u�:��-�*vaK+Zj́V4Bp�p��[C1��2�U�Wܶ�&���pW9�k6����6��e��ܣ"ʳ�m���Ĺ��+.T�Ѿw�T;�CS��"6��h	����{U�~���;����dh�tk���uy�hUt�2�چ��f���(uQ���:���0�0#7��R��C�s�g�[���8��kA�]b�bǺ��HX��4�a���HZ�r9���R��D;�e��ū��RK�iͼ��Hu�*M)������f[��ᝨ\݅5V���[�d���U>MaS�ʶ���tɵ�J+�Uּ�������{���rۗ����P�U�Q�k`�-��a[|�S�0
�.�+�zR��#t�i��n�0�F��n��:bݮA�EV�*$�����܉Opְ�N3���f���;�].c��AwqKeJg'��9�+)�K�\ ��ٕ�������)U�����]��۩�m29�˵�+(�Æ\|ɬ��
�B4e��������^�̔���u���*���Ǫ�g�7���pR�:�������k�3��{aZ&�$�(���GY2���-м��vSonh��B��*'�R���'��zv�i��m�r��
���9;���}��(��RA���J#[�U��]qۍ����L���,*e��M�Y�F�)����+�'�}\eхJn�oy��&�Q�oM� �b��]AG�\�L�9�fd�.�J�R%�Yݼ��]t���� ��mʧ�S����n	5QĦ�ʗ]�鄦��a�o�#�7�	.Un5���~ն+���WYAWa����O�[Ò���=)��o���.T�4hiJF�v�Cڰ�hԸ7w�=��#ly!�B��|�̗X1�jqHj�ff�S�IhC�]%��(-�P�Q�빂�s�+t#W��
׶��B�i���˓P�R�u�X�S�Q5ǷO)���(AYZ�Ka��a�Z���f�+d~#$��_�WIk�����Cg���j���Ƽͳ����U:0l�Ǝs���x;6V��^TLg� �}v�	l7Z�u*�c�7|.���r�A�Zǔ	8n�����;����]�\:�/`k�ѵ}feX:+���a�K+��ܶ����Uj�[C/�Q3q�j�+��Ԇ���gF��]zo�E.H�w���1R����Σ�wN�a�4�7�w�b1s�����9n�mX͑Պ�>Z�ݻm9J\d+NA��n��\>�7w���_Uvk�v:$K�]��O�A���3V���٦�����-l'2��z��������:t��2��*��j~�#�'R�|{�7���>Z&�F�=cqn���;��H��V ��9n�E,I<S۬�o��1l�N�v.4Mn��ޏG^m��
jLɝ�캹&"�������G�:cQb��Owxo�yc���1@��yݻ~)`&^����{�V��t��'��$�uup�t��UUk#�Q�S眚����Yr���%m�5L�M��J�׽�7��c��TO��g2�EE_c6^>�=,�]Zu�u��/�l�a�ۛ��(�:��ƀ�o�.w,v�W����{��a��d�67��2\���A)��oRg��J�<�Ѭ������9��9]WZ
_H�ʳg*R��r;�'U�{�)��9e���B�[�k�ɗG�>
rO8N ��ھ,!r�к8�^ٞ�h4��U�����S��:�	@J��E��n���r��G���)K1ĸuѭ�{�D�] �`%���bX�=�����_.{��N���g>á�}R>��sY�wZv��{'U�
�����K��<���t��9�J��E�ʌ��7d�����#���8�5��h�J�=�(n�泟���+eC��������j� Ɯ��VRF���V�7s�xCѰ^Ӫ�r���y_�RT���"���42�ͽ�Ь�h����]�%T�"�-��ik7�0�m7O�SZz���\׋�{�Y
�P��z"���X�:�뙌K�p.�5
]Bg%�`k=n�_�58������؝[�׬ s����ם���Ͻ���W�n21��X���S��O.�.#��&�r�N�{�c!.e���4%u-��Y@�+T�%F���'zv��hw���W�X"7B��UL��w�NW]�$"ϫ+��J��0�vH!�;/^�Zc�Jl[�z��Y��egT�����pc�j����7E^{��߷܋�:,����X��b��zpxo<D���Ԙ�Tɂ����\]c�N�Z-�y�n����*)f�t��� �#�u������A�']��#���ѣ\�It˶xS{����6ܛ~�hТ��� �2�`�*���<{���^Q�ַuk'�x�����r���b�k�Ŗ�{Fm҈����(��6�Cj*5-]��|ok��<�a�4�y��G-�r+Y���c��([�#G�[N5�F7!d*����W���a�����7�{��9�&�ʨ�ɒ�[�8�a y
4�v��ވ��v:䨴֚����O��P��gz�-4�oU����ƃ����f;�}�KCg,�TУ�5�9Nk�����Y�)k�}ꮗ��vWvZx0��n�\��w����W'\���ï��y5^�[�iT#�%IZ�5�sG����T)��u��%:�:yv�y������'Dً�l��/�V�t�d�v��K��\t��%�%���7�d����N[��w�2*o{!���Zi,�]��B�j
<��t���kF�=@u���H*]5t�ѓ����. b�_s,ش�LU�o��9(v�ޛ��8s�N�e����r���Gc���Ї���ܜa���&{�>pov�ż�bD��������ok{R�t��j���Wovs�=���\P�X;(x�=3&��-v��7v��1M�u�*=�=�j��v-�>�T�)$M;V��/i6#c+`�u���o�m0x3��謾ӻv�F�h��y�5l�La�x)Q˔��1A��}�A�C`��˺���������C*�9w���ӭq���wn��M�[Q����vD��÷MA<�Iզ��ZUK[*��<M�k:��Y��@슸V�s-H�a欱�ʮ\��V��n�('�.�p|!}~����[F�ΑJ)���մ6�;�jud����}zv�Yf���5Z�pΠ}[ќ���z�{)�ے�Z#�Wb���`;���I�/��[�L�Ԥ5"�;H)�Up�4�ǒ�Ag����>6�f��/2�,�|�P��)�c���T}R=�tVt��V"
��r��c�ױ���q��Rަ��,v5��,�y���\��=�����|L��a���6E��lT�Дr�*�E!���/4%�[x���]=z�5�mއoH�ӕGy�.$���n�9��sNҮ��*9k|����!چ�n�w*g/m�M� �$-�_\�׵�Q�C��.��/k�8�hK
�n�{���:�]E�a�V�T�$�5K�u�S��c��m�s*�z�z R��}�R�L�eݡe��V^�3��Q�y��+.IX�c5��	�6ӈwb�rL�q���\�c;U�
Vö"�̠l5L���η�T�Y�*JR;�=X=�ۗ�v��\��nEc`Hm�c���^�!,�� *�S�7Y,�gcG�"qP�� ��z��T��j���P��n���N�_mT|/7��H�^J=s�V��,UH��+�Wz���tQ�I��"��M���N�;�D�o&��^.�v�P�p�J�:.�j��V2�M�y|�0v)�Ь/�n��n�+��s�2��Zv`L�Jز����E�Ipjn.f�m�#W�U	x辧bK=	�H�=��`��SwpW5[�Ԭ�0C���آ4�8fW&�dCg5�%=2�a��ExN��s���t�kh�)Q&	�9a�V�V����B� p�:���ƪ=���y�J������e���[��ٻ�3����8+��T�����JU�^�[�h=%q�c�޽��\gL�'	��u|���{��v��,���f��a3����YN�0��K6a�.|�J#(-+,q�3���i��if�t�] ��Bo�e_����e_k�K��M�1��q)uRU+[��+�"cx�U�k������#`u��?1@W�d?��'�~_���_��o����￿�t^��E��
1A��d��]�n�-�/��iх� z�D��ʑ³�* PDHpO�E�b|9F��~���X�)t����`m���ܘ$��t�����D��v��CK���yj�f��d�^ݾ+Ls2f1Z�d5O-��R��.����]ع�h�Q��rAs�0�9��o4�)f�]ԩn��L��C�E�����m�ETl�}]Om��eg-v)��Ż�+,�#ZL�`Ȝ���>	�9.�N��s��%A���Xμ �}��F0���;��Un��.퉧�E(+!��*�.q:������V��E9O8�oK������2+�����]�ސ�\Ò�gDй�k��Ui�:�R���V�71�ǷEZ��:��{oB��6������$ʝi�]9��F�QX���:VDtY�ƞe�&�_�5��\Y��ڔn�&v�_b�v!�Z��t�i��m���ǂ���9ݥ��qq����B�vvfe�r��te.�{*J�C��q�7����,�l+M��PKW�G{6̀��q����N�鈊2U�|+Z��SD<���e�
��#�Υ�,l�،�=,�X+n:��
1��;n�F�說ב�&ؙ [gJٝFvj�ʷ��γ�S.�^*�E3��wV��*=�=&Mq+��sΒ����Uz�&`.(L�.>�t#h�%PA$0�QB��tӌ�J$���'�[(�A��J��'��8`(�����F"�(�D� Ȓ#	����dHL?dg�C44�
�@�֞�DQ$�5��ۅ���hiD�5^��J�T�3v��㏣�q�qǏ<t㶝�d$ʪ$k��7����R$�8�xJ$�(���SRB$	*�q�8�8�<x����ePT�}�nu��Ԏ\�L� !$$�$��HBI��8�ǃ�q�qǏ<t㶝��$��B�R\�HNw;@�r.
�K4�ÒiHg3����J"㺻 2X���
Sv]K���b��?JA&�$�"��e��DH!�t�Zw�����wr��W�RwU;�]��q[r9���.m�O^��Qy�]�:h���p�.kk��w;.��-W����o>;r�;��ڵ�:�BTԻQ`�KФ�h�MQEU��=���z�˛�Ϊ�7t���_^�Q^�����r���]�o����V������m��[����V��s�W�z�S��7r]��s����|��*��˄�jR��0*aF���
���D�GgO��r��]tNٹ	�w߯^{�ݸ]]����.�]��-�d��+���tWgn)���u!�wL�wA0��uݠ�vL���?}}_�w���|6C���E��I�R�}u�K��ƇPDs��ͽ�\+���9�vl��o.�'����2׏qw�q�*��A�2*�&�$���O��J��b�:^���[o����S��u��z����<f���G���lW>�[���W�}�-�����7�%D�]D���\�1`?P��>�ھ�"�h��'���HG��I!d�륩!�	S��q����C��Z"tܼ�d�R����T��EגV�ŧH�(��!5��[���&Ay/�[8��>c$T��
[i�n�Ӻ�Od:�%�'��GfW����Z�o��>�?�������|�M>�Ȍ{d��:G��������.�R%��Ǫ1���]�!3��X[��a#��˝�F[30v�B+`�4J1*ˤ�efl���G��ݶT{9/6���HT���O�uDY���ou-������g�0�ۼ��y�T���"���N�3��HFѡ0�}��(�6Ց-���ir�t�s^ �4�G����/���t��&�`�pL�����"LuhUܽ��%��׳3�dBkѵ�4qG/!:/���;m]��ց�\zi#5����S4�p9\SȠ�y8v��ܽPx�z�:W7r����EX�����	6Y�_�(��«����`�kP��g��Ge��׃,��vF�l��r&�,�K�[F�Z��F-���vj�F����Wպ�pS� �U�R%IїNsY���5�A;lF[�K�5&��ڷg��h������� �u(������Y������[<o�ܡ��퐧�]yPH�Nm�h)�/D�l;�oz[V�J�g�T7��NT	��_��5GW��xy�Z�(�k7p�E���ջX�s~qKeSu��8�d��}x E1����92ͽ؆����TR$��)%&�)��{,�i��@Q"�uXI�sWKOJ���e����jRg�Tc�>۷S�KǑǁH�Ŗ�taNNǃ�^d[ۻ11�R>mEPו>H읳>kgʔv�ڋ�գDѡ�Ż���WK�QD��V��"�D�����T�$�ޥ��{�e�pM}4��t�q����4�|�f� H����q/1U~���M�KF��݊7���#��x�4�Εd�
$,����S���.�pa��Z���~��[����k't1�ml
u �ױ�FIx��[������k|��z#R�;�i�cL:��wd��H�R6�-����[��f�ۮ_n��7~�������巄��5��}DDd>i��ֻ`���D:�ْ�J>1����Uf�m�kA�1���nG��
ګ�*��V*�7���A�-��J���V_2�� g�g�`=��N�ډ�h��`�i�g��N�V��d�lf�n�"�*Óg�t�:�S=N�{
�t/��u�U��dǢd
�}1��ʦ2t�.�y��W!�KB�9�on�o�+�������`0�W����J����2}��\")�v��Y_1�pMgm�>���i6ު��O)�C�}�1�a�5��l�/T���bK��_�M�s:�t��n���d��r�F����>�S���-�-�UK�:.�c���S'�I��r���?����wD��]�64�g�x��v�}�6⭙��\�6�P��S��j��������T�{VT]����3{S�J�F�ۊ�������z���`��ߛ�xff����9�hR�!-��v�����\�Y������ZjV�V?�d����ա�$��/l�c�y��s��M�:�Nz��3�#f�i�w�-��~Ӕ��̗�\VM�}�^�DJ��[��	A$��AR���Yr�u�me�ﲋk���H����1�@�����f8�$w�E*m��+[`�
���|�P���_S*���Ʉ���e��.uT�L)���7�m.���cUHn�����S��-u�(��j��}�f��b����D�DBݣ�≙Z^|��n5��Y���ٰ�Z�N}m*�7ea�s@!���{�D���%V@5�햿A�1�3T�J�;�Z��A�y�1�li��p[h$MR����ٺm�_����S� �n*��~Hm�qY�����%~ܓ&�}�ɭ�w���-R��dŻKm>1Π��^��܃(��}u	�Φ�ۧ�]r=�˷�[ã����Z�9�1=�ɋ�C[F�UJ������g��v�P����E�ך��p�qWՄx�g�D���a�wJH�R�h�=H��A��ʺn�[
xNf�����e�Ԓ�z%I�B�˚hֵ+Ti�1�>>m6��{gkF�j(h�Q�NS�|�z������ڀT
>k���T=�r]J��M!�f���cI�)E��&r��u��^�"�}�W}�X2������s2b���SxQ�� ǰH(���k�oޘ��y�:�}�8�41=�yj�ʩ�^�e���������i	�Dz�
S�[葲�,V�P��Vя��AD�[[v��boH��dQ�:M���A�m���D�w������F�LJGD��ds~��c{w�:��Hʠ�܏�e�Ɵ\�TU�$�{�X
�^;	�@d�%d��a�7a%�0�׆w*vsrR'o���1�M;8�O䍺V+H�E�#|����*a�����R>rމ��������tT��c ��W���&���݆�9�W"�	�W�;��8�(�m�!a��6dc�f�A0��B�V�R���*��*��mB%�a�ʛ�;zIĝ��׫o�
e�s7���֥L��ͧ��)�\�f�˥��j$%�(���]��k����v�t3��YV�wZ��-�97� ��t9n^��<��ڹ��ö���g�{<|||||</��w�vaj���m����[IG�[0c�lOG�e:a@f8�ǵr�Df �)�܁��P%�X�B[��`m\fĥ�6����0m�"�ٞ���<'u�!i�4��Q��N#
./!F��b��;/h�+�#|�Dߣ�l�Ϡs�!T����rqgp�u߹���%|���|~�k�Fe�vޠv����p�]}�krϳqɉ����|���ݱ	�r�ft�=v-��s���fxJyR/#L{G�WO���y{�y���F�I��:���Ls=�ѹ���
x���2�ˊh�^�*{����Z4�t�O�{O3�ߨN:򘹍�;WٻZ���0/.t�4�F�X�TUC�L����"|��Ri�%�h�V�OM��xQO��~�h���N�?�2)g˵֏- �0ev�X�b�i�����8Ƀ����۵������^�&-��grk�Co#�в��&�}��Bew�Y�ѥ�3����ty�b�qЙ+�V��|6��Ξ����@o��v#��k����b��T�EF�<<<<<*� �d�뢵}>�=������ #�^��>���5=��NkS靳�)1Y� 	��� ��P����e���Ӛ�^{�
pM��ڱ��(�􅷑���ׂ��&d����G��ԍ��y���
��4�9jYn�OH�H<��Rwwe%~.Ȫ���`�%B�4=���hR�S�cx5U�"�e�\6��F7��J�z�|M-Vj��
�Չ���i<-91@�S��\�`eF�V(���&�.�{��\��[����G��ş[��Yi���K6�����K߆`m�H�����	~^�H�2��׬m��t4Ä��\\{X�/Fk+6�k���^nk֡��+��/�yxj�@@r��/m&���/
��*=[�(��G�%@��R����A=\�齾�x�!7��s:�*����9w7f�Kl��r�mf���wn��O��%�yw�qK���Z��1G#Y���g���8ƚ4�f�ft*��6�M�ʁ��p�[B_f3]`u��7km�y���u��ނL�6�K�:a�2�_�����]����H�,�g�5��l���Z4��Ӆ�U�CC3���&�dI�X_|h6����y�h\y�UZ��d��'f�t3����~�ݺ�}��f?�)�e�Y	�4�&$��)w��K�%�P����ZN�D���2�Q'Պ�n�v3-�u�Î���	�y�^Z���f�m� ���{=W���~B��KU�G���MVsi{�
E(�$�M����F���� �T8�e�#F"wN���]�
�ך�|)N�0�����6��e��H�GL��"��F��U��nּ%@$��AS�uss��DB�'��j�w��^�(aUA�0'4V�̊�DAI�N�N؇.�mN�nJ$��1�*��_$��W�����r�<�����6�i�DE8D^�أ����=�����׫�Z���� �}��~]�NZ��ߠƳ��<�!t+R��}R�ܮHꭵ�KJ�Ib�H���o����{�0Gלլ�	�t��l��z`�E�?3�����Pz?�%w�Wl#�0%Fa�x�-E�t�<���+��3d��V��p���Y �ۓ�V��Ͷ�����J�w)R]P�͝�� ���|��n��S½�>>>>>>q�1�̖�Q�}b�M��h�U�Ѥi"eix	��[_�H`��lc�ժ�ƕ����P��T���R�0��������k��Zj�Hy�h�퍯�á�F�K_N�թ'�v<v�@�m3-;�9Pw]%�6����,�����ꁖ�Ϩ������;�@��n�l=^$gQ�� �Й������k�
�Q���cB�XPu6$�;B����coa�sY�|Ƌ��V�)Ϻz��:�*4�iI%7����.��Ԯc�����ک��i���mn�N%�T�8
����н�%R���K�7\���s]�k �L�$C	U
������o�Q�H<}Us��E37r�8k�|Ƿ�˼�.��5�f���a�i�і,ߝ�}�Ͳ�p��FԊFU)6)>YU���^��Sc�؜�juo\��լa˘�Y� .Uu�YK�;�1J��s�0f�ԗ�����	$ I��hx��,�jC3��ʸAJ�&�ջ��	gZg9�*HK��.Y.���g�v(ق�Y��^��/P��kn��5�����k��S��`=!�O4��P���D���@l@�;m��Zo�O������|]��$"x�{w�mN����E�7p�V߈�fPg���4FaF�N&P�ʂ�%"23Z��7��6��׷g��R"a�FԎ�4[��t���d{�fXc��A-�/UY���-܂���$�q��SE��7\������[o���i����EZ�+�������lײ�J5e��e������5��Y2��e2�w(��1β
�n
7=��~=��¹˴�����KhK����֝��o�
71�#.|��܁���a�]0b�R�UL���}GI��;�|��wՓ#��N}I�>��К�BA������|�Ձ��ջ���Ep��T'a�Ϸ|7&��zk�9�y%ל�6p���`��;��x�$�����͵!���Ca�hc�p�������[׼)]`�2�u��Ԥ	s/{'1��y�E�N��%�)gKҖ��Rf�8�h]z��&UMnf��.�ѣO�����v�Jy|x*�t����8x4��W��o���&�d4�O��u@�����V�{��'[{�ͻ�ea"��j]ҥk(e�6�y��ux�ν���Bߵ��l��n3����S�m�]oY��ͨ�q�s��i�S��t�h�R��Y�0f�ځ�L���r:�k�єy]dR�*=KL�x�f�Jmʾ��落)�)r��Hky]=�e���˨�Sz�X����!=a+ܙ��w]2;��N����&2���Ś�:p�]��:���pd��mWQ���Bu�̺k��z��
�Y�k���ٵ/7�=�xH������Z��[r����,�ӽr��1��@�$i��Fuh�,V{uZN��NL����T�5��g��У�k�Ɏ�4�Vc���q3�Y�����y�s]�,����K�Pܒ�J�V�v��$��vw%���c���R$]Nc�����'r�4ly�T����E6���dW�Lvo��6�v>0��W�� k(]PU��ஒ3�B���0N���W1LH����Z�YO�V�6�e�Ij[Fg=�Rr�����!��U�*Uh�m�b��UKʌF�ʬI�$�߻�v,5+��>2P��B�������6���k

�^��m�|a5ٱw���������#r��Z:q}5��2���ʹ{zJ����MMǗ�2����zH-U�B�r�tS��ROn�6S�����âi�:%ҍQCJ/��Bj��/�Li7y���u�uډ�!���V`ѪX!��%�չ\ef��ПB��U������,��{��빋�՞�t�u�-K�D�aƄ�X/K͸����ɻt����y�����Q�z�wӤ�����km�Ⱥ����)��ĕ�N�BӖ�$�;"�o���x)JȄ��r�{�FT�^9�%����G�u� ����n�V>M�P��R�CGqwV(,���Gwc5�n� ��*�rܻ=Lgm�]�sH꺛@�4�y9�x�!8WDZ�i�f��9�p�;Vҝ��1i�pSd%f��/;�hW#���dz�Cw�=a��k�d��*��gm��iC<��vZ�7�g5s�:���Z�G�����65�]i��	����|�e�r��3o,�wr]��:�{:6r��IW|��"�_Z��m����֔L2���M�t�Y�-��n��pA�s�0�l���^Y-83b̖oW]w�]c�f�t]��=�tخ�]�gS�r��5����uZT?>�����������/��-DwﮚL��]�c2h�|O�a�=qǯ��8�<}}z�^�>66[�!�$K�� EO9J&i#�s$#I�GD�_^�z�1�8�<}}}z��O���\�A�dH�B-�����H@�`H��7��ߛ����w�~�ǯ^��<}}}z����m��$%<��I]�����4O�⌤�1����`�$����8��I�fyrIw\����ɘow(` �:�^����$�g�u��~{�o��("s���\J&��I!�H�&2$�nX�wN��$@�����ҙa��I���u=y0�L]�$�v���(����d	#$�B~;DQ�}��缉�t�2aM4����
��GȂH$��T��m�I��pH�8�t�Ì���է(1*ូ����Ⴘ�*�>\v���^�g��׏F��i��I����@ Ҁ.��z����_��-�4�����%.����DT>�D��q\��!�b���7����C�\�%�le����ޭ�L����^�'���I��3��9�U혚�	< 	��W>�ܮ���;i}�UI��5]�V�y�S@�=B�B�3�z��d8�x��nAp�d�|�x{޽ݐ�7'ū*�~c��a$����<����y��>0UW>~(H�t��p��OL;���x+3�-�> �����zЯ����O����&��1���n'�n����t?
�����c=5v�Q����xw�{ޖ�����F%�:����U�^{�+�(��kpy������cU�0g�������`��T����D��wt	dB�\���4��oM�n�#�֗*��H�h�ܗ�P���6o��.�4�C}s��.q~F=_?s�>�Z�%���L"���rø�..��f����op/�ZF�0�~ q�z �������Ȱx%}���&y#�S����^��N���\����x�&�/%��q��|h�:��D<7l�*��]��z�(��<1v���6w��!��PGw��
p9t���(��j��yB��{�#c��+��j7���%�ߴ�t�n�s���}kI�5�]SzEO/7��08��睋uꛜ�g�!��\M�Mh��}�v��[z�=�Z�|ɚ�>��� y���7������^8���1N/�>{(���W~ŭ����}r�4B�e�{�9W2$�C�`��f=�J�	Yy�<(�K!V�S��o&�
�W��@�X`��x>��������Z�(F���3q+��L��h&ـ�|��翽�>��?2b���u��K|hz�BmNn��:����W���~�|��|s�w��h~d��cZ���/�<كr~��2�����_�'!Sl�,�o��8��C8L�nr썴T����������у@���޶���2Cc��U�@��>�	C2i�P���*����P{���o���A����es����?3>�s�m����ᡱ�g<����n���9;������_FW?%����%�!�ϝ��ꖞ/�� k���\5��c'��W�}P��K*��t�MuNj�}��ӏ��d��d�j�O�H����:�Jj�b�_�3�	�#v��X�=;4�����x�������)�������=���2ojFu�9��u�_���:��l�qm�4i��r{�th"��՟k��>@ _-�cx�*�Ю��0��+�ib���U���Y�ɥ�ُ��V��e���b��uǁ3��6(1��
݆T���ZX^�m�|1�|\�"�<�-��YT��6Ї��x�m��Jb�'A��J��+w;�*AT�kA�ү�������y���%J�6�]�
yV^^�\�B��<u|6���s�Q&�F}`H�؂2I)A(�d�({���ż�o5UEmh����TKC�Ҙ8	��O��w������c~/��c[y��q���+�\��yꫫ*㧦��|��ﺾ����2�%��X��p�_Xl�ݎ�e�`�<�rw#)@��W��W���ӛ#�s^��@2<��2�]����8�Bߗ�Ԧ�ӑ�-��_gr/Ww����7����14�����Ũ�p�������7�~�9�:���XO�$����n���K\So��)��s�= &UǴ��Ih�X��߹��)���֙�;f�%��x�5������&A���]��}I��u���a�=����0f�6^,l��
��^k.�L3���0
qO�u(��RFx����kPXHnu{�fil�����,4���;5��
p�N+�6ZW��]I��
��07;�	�ֽ���ռ�#	����j&<��������Ղm�<|l���>���:��;(pk�'��C	���=?x�&�=:D�(�\�s��˞����=& �0�z����Tc����t5RM��pA����VB�ϻs���_��%��[�jj^�<6��gr<_��K>�7�o�˚q����cF6=���z�N��&��
K�ۢ�0���_"�����S;��;�"�cQ���V�A�ڈ�S��Vp,�9{C��l���~�x�����l���RK�K3��D���z*��e����k�</;-���	�?�	Ō���n^�������	|��z���s����<5k�j�-F���i�a��y�K?[��.���vʆ�(����������q�~�3��Ǡ��W!h���
�K�I�o�cr���;��Ζ�� ��{�g��څ��T8�鱻w'ۯ�������x�B=]U|�ƚK�g˳;9Ǽ;(0m��Ve&lR�=�#�|"�@Wǽ������>��=���K��l!0j�.�
^i��y�g�����ڜPⲼ�+H Y��<��ʌx֯�G�Z\Q�O~@��Mg9��
w�e��T����7s�-�U��\¼� V�J�?*B�pv|"^#������Ό�i�]�Ph�2=�6ny�'��Q�nO���Wc���!yB�MN�ǝ���Bl��#�'4V#�s��k ���'qI^��0�����JwM��N�*kfWk���u�j<�����I�0�΃�ƟW�? ��
�Z�R�/�n����{Dt�ً�����U.Tϲ�՗Fk��@�n���
SU-��ע�f�87N�э�嵔�D�#M�}�0��K�e���%�ݺAvT8,#��121�.���j�}π�5���y�)葅l����O
���xT�>;T�Ww�:�cQ |%@t����_�{\8ޖUU4��2%���q��-ᆺy;�V�w���g9����'�s/�\0��Dn�|P:���;�a�������F)�6g�u#W t]$���,���O��G�]'-�ٵ����|6<�Dx�y���m�xLm��i���.�40���;^��p͝�s��m���g�����m�P�aQC)Q� ��tXU���YZ�����;�u�0g�q�'&�ܾ7��sL�'$8))�N���8ݵ�����e,$P�����_���0ˡo
:{� *�v�����aF�׷e7�逆j��"|ݝ�=���jM���8���ΖUXw�+��H(��Ⱦ}�r�)��� ��wY�&���P�u�8���za������^���\+���S���a{��eEt[j��Y]�
p�[�<��^��`!�w��S��q�(#�V�o	홸s�Vհi��z,ݞs�<˅w�:�����f$'�q Sw>�� ���O.Z�ִW�� ���ow����N���󗭋R���חOzz��rrU��{�;Q�	ȸ�_d�O��J�n�F�+(49,��q��p|���ϮNU*�T��^vQ�(��m�qx��W!O��4�ߛ-����ٍ������{�G������KcIQ�_�̫�ߟ��h�����Pcʈ�I��J1��>ʗ*�s�_��;ކꪷ�\$�bn1�ح�����1g���P�t�O�z֟�������9��-�����½.*m�y7^���]�x�	+�&�Dז1��G?�?�g�6�D�<��렴��`:\���\�B���xƻ��w��qlu�$bXw� J'�y�a���C�����~��F��W\8��3s�`����<&�~��+�����-���A��;��Ua_:�Lb��~�|���=�T&D���s�h*[)Y��2y�$����w��s]����m�/ݦr|�L�:�zT����2|���|�/t��m�/���r:�lw�L���ޘl`�o�[yQ�,6�Ʋ���z��������_A\�M��8� ں,��:�犯22��#��p���!��۟$Z����pm9�`�y�,Е[Jp&+xsZ��ɵ�%ox�Ǣ��Y����3�l���ϣ>z�����ဵ�4ħ�� ̚�/�i=��<.�E�.���e;��%�k�l�;��\�:2��F�v��m>/��3|D
�������|��a�%o�\:���c̚�vȞ��h x˻\Ze�g�V���rUڶ飥u��6WF��0�L	�� ��s�ZSr��D��=P��[yt\Aor�\�*��4�X�fn����8*�t�[���m^����ڡ�A
&�8B**2�)�E"@�JJa�������T)�4i�T@$R�����rs��3�
�����?��y۞��Zy\��A���
ݟu\��ֵ�����S���=�����^|��A���8=��`�K>������g����x�ѐ X~�sl]�j���0�G�k/�;РW6�F�Mm@nB	׬xɽA#8�AA�똨u[ψs��ܦ�c#T�I=� �q|8D��vi���3��2lbͮ�O�c�L�_u
6'�0�F����L�	0
���;�ǼO0��O�tޱO��5�Gsȷ�/0o�uX��L�� =�=/<�뫥Wruڼj6t��ҼO��z3=X~7��d�b�P@Ys��y ���{$CM��*��z1fpMz�橢곸��R�2�Z��H��@�^��n0��G�pQ�0��D@A������M�f����J�~/��
/�tSvyGq�=���h,�/N��;���/�A���]��?3���Cđ������P#h�a&�K�jn�U�'�tɾﷱ��x��"Z���;�cx!�i��T;��98� �koDl�5����3�S�.�]I�v-�}t��'�֒� /��?w��]H����dNP��e���b�&����}&���I��'��3_U����)nQ����~x�Rƣ(�t��{�۫x�c+0���c.fS�d������4*���7�^��8J���i�"F��1�4�RA@�~w�ֽ�~_�;)�O����#���
	�Ln�S�]@Ĕ�3��:o&�]PX;�|a�=[V�W��\�7y8�{�Hq y��L������)yƵ�t��ϋ^�ŚC�a=��w��q����E�`OA����������<���{��'%J��
 ��r���}��<9澜`/�}	�T;�;���@k̓
ꚢL/���t�O+?
���'#����|)Y�{��EZ���=��sG�&��|����V^Ҕ�L^�P]e��C�;0[�D�Φ=�eO��q|�%��ud��Ԍ����c��=�t�b��z{���/zY-�������eĺE{�:@��?}��C���f�� �}R)����kl;7P��^���M�`���s�㹚*�����x?Z�K���k��ꢻ������O��MP{��q33S�U��?�� ŭ�/;cC�I3u��[$������n�9A�|�h`�e<:�ϼ� \{�^t�M����|w�^p���.� ���c�S��;�A�G���ƹ���@W��Fұ�Yc��YQ��V����\��s�����V�{zUj���閠VF([Hmc�s d�=�U�Mp*֩��ZDv-�z�|� ��ۡ��P�E��j�E��/A�{��V��G��^4b媃H�b�ZN(7r��s��4�E��k�أ��p�j��5��=�#cJƘ�A�Y������o�G�fy:��\�q�eK���%r�B
�k�@&��c�2��&iRrj�ڎ+�&Lt8�a�������naܪ{����01�`:�Ug�څ�l���W4Gw&��4وb�� �7 Fǣ��D�a̸LtfH����g�i�&^�Q|黝2og9wZ�7�zr�Э'b��n|C!s�wvWi�U��
�95{,9*??C��y�ait��B΂�t]9x�"m����n߯����F�� �3`�`�^�XÄ�1����F����/6t@���;E��a�����87ӌf+"I=�rbi���{�=�m���χua#�c�^�}@@����C�m���^���r�{o:�K���R�* ���<��q�(�y�����;)0�r���-����/��V�a^2j���S��rS���O�#�6�n�����i�	�s61[�E@t|���	KWx,4{�\�Tѭ����@lÕl�\����R��)�փ.��/L:�v:��w�5�u�
��D� ��>k�yTUj���=���ݔ�OT�-�zi����͹fS�6�gl`�<�u�`�6�guT�qgi�6�Iu:��!�#�����\��Yõp��>>%q���/��"5B�R��;]vN��&D�,Ƌ��ǣVg��.�f�%�lɶ�����S
`�ܴV���z�I�/|�>���Ɣ#Lh�G�w�Dծ�Z��v���ͼ4�,�ݤ�*1�q�+?X��"j�F��o���8�̑/��&jጦz����e�������}1e���|g�7��X~�l} �;��Z�����S3,^�{�Fᘻ3�����=�P�moX=��U��لwPk������S���gDK�`1���]��ߚ�#��N�� X\8\g�N6��fG8��,w�3�=4�b'�u�����x���ϩ�ܫ*�63�Jo��.�K��l��a��"�o5?l��ܟ����1���r�j<��t8w8�ku+ϩ13矰�}�"���z���s�F���/U�"�����= w;'C�uŠOf�ϸ���fk���.`7,�ק�}{aHty�p9������J{�L���]����yuL__^:�	����o�߼�W���<��}�DW����VC�X_�F��i�q�LKl��pn�j�3O��W����=��w���:�m�"|��=�SH6Q������Ԕ妡j��}�c��B]�1��a��1��Y0��:�4�B�~w��<�/ʢ�j:NB)��
�*�q��.1}_�dZ�v�㳰���� ���]��k�ފwI٥͛.��w��8w,�ݖm�F)��s�5t}R����s��Tț�I6�����L��7#pb���Lͭ��<�Q9!���`��2�F������(�8$��E�ٖ6�d�K���:��ܮ�wS�e�N�I;����M�*�,#N+bUZ��	���`�א9.>۶�DF�4]�r�*���f��]�^Y�`��y+P�C���SWGl��5�ƙnkM.�|ʇm�!=$�[\͡����y���mp�5Sp��٦�U���t�ڲ�(��\�B�s�veom�#�����uj>�|Ȥ��L��1��){�Y刂����nc�J��QSmtv;&����ǫl����ju��A���b�MK�q*u��`��UNU����m�hv*�7�4]��6(�5b�CKC(�YB����9S��B�PĞ7�=��Q�teګ���8��v᫋�^�x�^���5c.2�0��.��2�mC�p���4��$2W*��_3v$m�ZOe��9�� ej|�Ý&/��u��ӯ�0�q��^ݪxX{���YzF(�u,(�.�͝s-t˥e���\���49��y.<)�<���cH���]��bj�U-�����*�y�bTAiXM�Q��2)D�A�Ț�)5DRBV$s�	�u[~�w,G,��M�B��	�l��4Ed&�-�)"���&�cE"kGfך>&��iP¼�,�����j�W�W��
YVc��vX���V�r�gB��@��|���L�ٍ3�y���VrPMŗA�����#�m��b�n�lmZ�(��ǳjWDi��x��6��{c��	(@�݁;]���t̻���fwN�^3]c���ז�whx})�t(5!VzQ	���s�i-�6�Z�E(Ƹ���r���;�F^v�ۛ�c�gt$t���5C��3�]�`W�I�)�2kq^1��WR��T-�$;�vr�����y����}Kv�!�+��!���+D����f�[�LX�l�6����fvW�P��6ϕp�%�y[]i��6X�8]R�0T��W0V`E�S}I��I[[99W	m��&������Ѷ��h�
@�r��.٫��w7�Zٵr��Q����=�(=�%��z���g6�@��yCÛ��!�k[�9�ܱPѢ��";��Y,�g�s���D��^jT&�;�5u0�Y�-e4�*�>Zd65��Q`�G��7���5���m^�SW
V�ΨY�f,�Z5Տ�h�.%�M!-�@�N��nGZ�iA�njhd�$�רm�#�J�ܶaT� 7��ݖ�wNr�g���e�8��A n�>鏹˜�7��<a��h�&�0يJh2�����D�cD�D�)�(�(B�Tq@��I(i�F�(����E����8"`�n6-*DA��P
�It��Cb�2��%b!��	��Ӥ#$$�!�]"B,%�����+\K�E"�E���td�wu;��wn����c��K|\�&��M����ׯ_^8���^�z�Ǐ��^�||j�I$
�2�$;Ut�㱊�`��&��� C��^�v��[z��ׯ^<}}q���{�.�cF�&��.b���4 �帽ݗ���c��jrf}�?w������x���8��ׯ^���׏^�>2�S��@��5J~��8��;]l��<��/:�faݺ���]ܑ�]ې1���&;��)����ݓ�{�wu$F"L�D���)Ή�)���a1�Y	(� wn�9%�����),@���� ��!�C$��ܮ�>]t�6C%�r�h2Q!H�v��
e��]�!�(1D�2~u�e!+�qK빑aBɌ$��@ ���$�$��i_�^ah��җ�`˷���()��O���|g-�ę
�ƻ�.������3|�,�����*#1<u���p^x`:r����i�u�:�ӫܖU͟`R߃B�0�ЉM�]�W����O�A_U��e/(r_�O���i9�[���2=]���Jso�/�އB�;��u�b�v���� ��w�?�H{>������k(_`�]��p�~�7��	��
��ak��P[#�#*5,gz���5w�M!�rp(;�O^�����X��na�w\� ��`	N�wta-K"v*K=M��,vmn��p:�++���~>0�Ž(��|�KW:�ɦ���7+ڏS]�i=� �`�K��^��p7݈ӆ��ϵKO���%|0u�'�HxF,x}�זS`��$�{�x�	��{_�q�72�A��O�O�fۨ���-.�aE����/���L,��2d��!�8��½�\�C�q<�׵	����	eA#K��`L	���\e��7զj8�w��.�	�7&<2��p��k���m�q����02^�T+�z�L)��r�}�O�MB ���{Y��q�y�+�i'G2i�U}. ,¯������w��ցQ�6;��b'��=�dst�xH�����Լ�G�pS:\[�zm���4]{f�6@�y Z��A�����o�h��ɛ�f~CY�����-��[�\:/ht�Ɣ�.4,]�~%d޾^�u>1e���P,����K��մ��+BJ��-Gx>��5��B��si��W݉ձHtь<�WG����5��a黚������̾k<޸Bo�ЀSC@�M ��;w�;3���������(�K��|+��ܕ7��ŗ����������b�{����SZ�b5�f;�ذ���i�}�%�ە)=��p?����U���kN��;500��"�{�O��Y���)-�A�?K�kzm@�V�0���� m\�	�.*a�#� O�D4o�a����	��[��p���o0�n��L�З�~oT�����o��]I�+��n���	���ޤ�M�B��ݞ�0�d� ����`�1`6��F]�/G]2�L�"��WP1'���Q�~��I��F��ْ�[u���[��?�V@��E�W�`i���	}wR[�4�wP%��'��Zıi|�{���y���������o��i*��2jJ�Į��~3�s�a��
YkZ'��yujb�mo8�5��Mk^9�ڔ� u�(�)�z�\[:y�y���O�y�ّ*�ŵi�>��Ol^�ۆa�qM�p4���Ja�""�	�&{�^5+�Z�-�_1���<F߃�\�=�	}��@gҾx��f�{�`+_��8�v#�>`l,{m���`G;��ͮ9��2�U�1g�q[�� �a�s!ޢ��Z9:�9��j��4�ǣ��x൷��9:˓31쑜"j�ʂ�aP'����jݚW��M�%�GwW����-�-i��f��T��4"��҂SCB��	��Aw����'���>0�B;�W�2^W��PQy��5��A��e��ƛ񕼝ZW�����ol8\�C�lS �� [E�	���57v�'��K0�l�*Ȇw�{����s4���6���j��?nP�@]��
�7J�/�׭�/57��"���b�N6>��WF>���Q����6������a���>�ݮq��ߕ
V~F肂>>�.�-��SȻp�MC�=���v���}��0ɥ>��'�cYv�0�wO0!�+P�����** ,r�Z�C��/��o�Ct�#��'A1I��)�O���ڤ�ܷ9붚iv�L�w������~8)?�����*1Ӓ�gƺ�@���d˔��X��L���e�d�~����S���Sqq3����<���kLh��=
����Tkx���׾m�%�r}?u���p�n3fn�UV8V�d�T{���i�p8}}�8:�3q{�L��z Cp~ּ^���@Nu�a��4�-� �������O��fO�ֻ#`�(h�z�h�x����ǻ��$��(57_3m\9��X��\���� �f����ne#�"7B�8{+Eȵ*������ƭ�S���^��	��b��<y���	Xzb������P��u�q��x�^����{��y	�5\��W� X�Q
hi)��R���>s���ϒj_���aH�Ϝ��^zIᚇ�]{B`&m��?���	��k^'����MUf�X�_���k �=���!d�l����A��9�0��U�"-�PO���G@�s5ї�D��K�~�,�A>��>��Y7%����>�A!JR��Bsk�Z��v��ķ�C�Ë�i�W@p���a��oL��*�Y6�H��ｙ6x)���7l��~g��>�G5�Q��wk��GyD�q ^����g+,=0��ϟ�",y�v2��z`-i�*J��]Q�o����!�w�������3�<�b�����Yc�0Ovz2v=M����n5u��+Ok	�R#���D��0^{ˊNvŰZ�oD	I�{��/>��y�A�;+�"�]/swi�ż/�[�d��h�D&��}N��.������·����~x&���D�(E'��'ܝ��!P#��8�±Ƌ� ��Ds-�)������cln%��'6���׍3G�Hv8.���q��;��WO���PZ|ޏ1�pK�k��㬞e����UD�����^mK
^CVA=�퀏�5[�^z_}xi49X�`⩾��<9Ɂ.�,BpY��e1�f�z��$�H�4k�;�X �eJ�w���$��Z�E��/,pB����k`�[moB9U!c]hZ���qI�pRi� �8��ģ'����"�5>���Њ�CH�M(
��I������g�Q@��6�`�
�����5�[��yƽ���Q�nm�0Cl��Bz�-X������5��tZ�[�^p*���3�V7H-#�<�F �	al�d1�����(������om�W3�|����k�hU�����V�s(z������XW����~�ږܙ�ޕ���\��U��T+��6�n�k�=��^�2S��ϕL��w��c�l�N�Vň�kB�鰵�pu�0�P�o3e(���a�Ʒk�c�T��'�6у���u�Ɩ�z�Z\��;l�Á��Lkz� �O��d�� l'20H8Y�k:�`�YEf�A3K��g�j��`b�~x�,`��0�nl	����Ly���r��;���SE\>������Gg��0���C�6c��6Y[��D�c�^zc_C�$a�_ǝ�3�.��&�l�3��?
�n���=�(��T��w<y�6��]�{��ω����bOf|y��.���N7ew9�ö�f<S�:��z�#�f���d�5ϫ�l�@�k90�>��b����'ޫ��5���ۺ�f�=�w�S�Tz���u�<{��j��n�h�g@���CS���vP�:sz�)�ײ�>O:ْ���)��p��;��Ν�U�2����l�&�<�q�f�^V��L���ל��[���x��44����(�~fs��_~|����+���׾{abr깶��Zڷ!��ʂF���pse���ϳ�����"z5~`��
P8>���9����|f��>t�gc��e|�O]�
:b� �.{�U��D���`[���
ְ"���Ԭ�4>����B\���o�B��ļV�}<�fF5�;G�s�N{�P�I�!w��Ȝ�`��f�6|}���t�k�MԴ^C)eMK����Ӕ��7w1��W>w8M!����T����$H࢘И��i�^6��:)�;�[�����JSHܩ<�䢛��09�õ<����zw��M�Kw:pE��ĊZCfGCkp�!��K�S�R$г\B/,E��O~�ʸ����6.��I�W'a�	rs���a�0}b}�/7����"A���1.�aG�U}t|@q�;jt����W*x���OU����B��������}¤Z��WQ�)�$g��U5��cΧ��\���ŹTs	;��(�^|fv��3!�Y�o>C�u�I`�_ö���W��۩�<�c��eo'�l��ǎ�/��O�6��;5m��ySz���]��7�,�+7[4�Ql¡ؾ
��`)���$�}Vc���2W\�Y3�t]���i�{,��F1ڰl�3�w۴���9:R�i�y����x =��4���Ј�C@.��gN�ϋ��p_x���\��ԨoJ2Jz�rP��	����j;��le�V|�޳X��5�W����C�ȺU�	x�I��>��I@�LS,P-�Р�yw�$�l�<��ǟ:sA:9K߻����M�z�!!m�He�Ü��qV���>��-��Z�Ş^4�ͻ�g|L�	�%��b�7�L�Djq1q��Kս5Ϟ����}2�2T�H=R��ט��ޚ}�QRG�kf�7ErIl��T|2<juB�/�� �Ae�����T���-�nA�|7�s��0��uF���#5</uI��L�	���U�E4H�ŝ�#�~W��{�d�����a�O|�Pњ�n@�e٩���h��B���]����3^�oV�������z���^��v�K��eM��j���a���	����a�Q��.[��/L��|�E�a�ڛ�����N����7z�	���k�\��)�.���(������j5,������;I��7t�`v\$�	�u��T�~�y�Cwa��͸H�6o������GY`떾ug:.�lj	P�sQ���UG�Pb�����h&��[����/l�� {O�7�/w�s��ʭ�j�MͶ����(��]��v�vn��N.]u�u��xW�'�g�NL��5Z�&�O�-�P�@B�Q{��g�5��>{�mi�HM?�0y����Ƈ�}��%dv��Re�(�r�j�����o]�z��g���sc������W��j���l5�s���h��[^����"�<ʙ��E6��[O�
���O��_�^�4��I1�a?>������ĵc�|�jx�f{T�W��p3��+���{]	=����0�l�p���:`r��l!��2�V��'��C�Qz�v��0����J}:��ҍȒ��϶4���dֻ_����,W�_�t~�GudG�%�M��=����l$E���>�LZ_2���y/׽�Z�I��ACS:�G���8xQi�_��Hl96�ۉq���ݡ޷R<�ـ�d<�9۵�O�=��������9�&z}�Ϣ�����f?Rq�n��	׽���:��F:�p��ԇ/�����f}��=9�*���϶j}0�ڑ(�aG[l=��w����-�ְ��}��N0M�ݔ6,�}��_{`iU�,�,/u$�>�l7�j}/ߨ���
�i�m����I�X����aʛj�����P�OX��]���6o����b�h�mP4EB-3R�D,d�h#J�,���r��Г8��JQ�!�RJ�t>�/c8�7S+�����]�,���\N���D��dcy�q$�.4
'B6�d���U�\�}"-?C@)M
44�(j���^o;w�>h�l��*?|�0;B��J�v3����Ң���
�c��o	������?t��EE��̭Z+}�;�Sx?�D�<�v\cc�Ýqܝ�4�bOP����3=��!�%fw|ʋ�ba�O�]	�±Ɖuo�̓�xO��%��p�[�Wf5�őL�N�A�-ee�e����DwH�rU�5����Muw;�����[�Uu������<���u&�]�}\X���O�a?����z�h��2��Փw�M��uK&sR��vtst� <;b��g�����f���	���.��0����=����9���ˣw2��c��Ʃ~z%��/U
�^N�qC�4���GP'���Ȟ���3�y5����.=��oѬ�BdI~����Z�3�������
�׮-߁g�@)�V�=��5��L���	��B�1A_�h����qp��+����mx�kv��#>�L�����������|��V�
ЁC���X}�_D}ލ��^cB���s�0�a�wq:�k�~�$�E��l��$�2s��ի��߾�^�G넻�BN��j�<Z80^��aNP4�M���iL��_"JN���n�����ϗӑ<ϓ���D�DQ�Q'¼O�PJ�S�ߦ��#X�ہ��}�G�ֿ�����9�HBdWb&1�7����3���j7H��o��g����.U�@O_�Ҡ�CB>�   ,�Q������j��\���z`ꠐw�0!p@���Β=�P�N���n���ϰ�//B�ܭ��Βơ�"u���̹݇Za�m=��3�2%܆�-�zj<��.W+�r�Y�+:�����/_������NQ�n�-������¡�+��@����悛u[�[�y���p��t����xKIN���8��!�R�]�y�1�Tg�9eOv���':�Rz��2'��EK�=0�o��rq�:?�z,�!=��J5���yƷEl�Ϫ��cb3���Î��k���.yV����-dheo~;	�跼���do3bg�ٚ�g����TT�"�3����U��C���̥|�?�������ZEG6W��0v���t]��̞R	�j��������+�]�ٶ�Ȧ��Ʌkzh>4S�8�!׃ug=�������Z}x�osXo�@���L�p���Ȯz�P���[dR����~�>�\�����vT����@�ox�?�7`�m;�%=�%ܟ��n��7Q��-�W�c}�^��Ɩa�(,�'ɍT��#2�{iB�U�ၖ��b�+e�'���i��#��G��ͽ�eյ%��ܥ�#W֞��76��]zY��{Wr���34�'�u�^�)�Q�W�2���7àX�+{��Zz�u��cS51���Z.�U�GƎi41�5��3�8�3&���ql4�������A���F��.M�u˹{�@�;mRĔu�{P�U��ٻ����se�~���b�SiL���r��;��e����}e�n������AY�{e�]]9u��+D�:����S�x��k�<���b�f��M����Aq��qp��N�lK|bpuM@R����,[F��m#�yM�����,$&�Sy�T��ҫ��Wl�Qiۮ����*+1�ۅ��DCAt�an��Y�$�-Ya�S�E+��]�(&�eBAobլ���
[�p+��;3�&��u���A�5�Tk/r_w!�{Oew'�/n�5Z"�y�Ų_8ĽVs�As�5�:��;	x�%y�R,��W���@���Nے�5ѼS��r	X��7[�Z֏u#�7�72o4qh�3�M�d:=m��*�­4{{ptT�s{^GKj��CH���վU���WʥfՀ*q�ݧ*�X��v'i�ޗ*eP��� �%PT�n\�{��,��&�\��I[]� �[��U��+��zmX�cj؊6h�g��,J�2!<�Ydq�s��;�,��	͑���b&����7)�g嵥�MQ#X���Wod���]�7���#�:���".�1)E�Dt�YD��ݷ>�E�9��{��)�9
A��*2`��J���Ly�4Jci[6��	�gS@�����l�(k9��U���9�5�h��X1i�+3��ͧ|`������|�ؕ��<7Ӕ�hjJ"8����G�^����%��c��U��4�u�|��Ъ�Y���}�o��g��Pf��p������4!)�!v�s�7S��M�kE嚃���`J[�pK��d5�]�� B�Nn<w�{�}U��ö���ì���Z�#�pp��CL���q��r�&��}��Iz��;*��5�j�+|k4	�ͨ���	��iꮙ�J�tJG��!���ӗ��bpU��o!�	UG���v��Z�r�x���<4M��ujT���b��f�g%�R�%k=K9�{8=Mun���X�GD���UI�+W�6N:�y׏�A+eY���L�)�F���-a��؏:���u&e'F%X	xo���e�i�r�c�)�[���2\�ZwÆ�.�#kVS�������L�/;��A������^sւ���=�o�]�Xz@�n�3S?֨xU��LIoչBW��W���M���)2L'���o�v��6�8��8��׻�}�Q���W�4���w���BF2A�y�}�BHLq��x���m�qǮ8��O^�>4T��B0��5�I%W ۗLt�k��F����Io^�>�t��6�8��q㧯_�!	*�UH{
�HH@�?[�21�͵���tM9]HJ�롅�$�����W�� $OwB6$�I%m���^�j ���\��m&��>��-�b�a��`�<��6��{F���n`��A�1E�"LA�5>9 ��6�ƹ^�E7ur�4X�ܮh�9�d��+�ӛwu�DB�Ky�绹f$���i{��pל4�륈�Q��Uw-|^[��(���Ϻ��]ǜ��p�5�K���-�i��휗p���mR�mS��O�/76d�%�>�2�6���i�����{�^�z�hi���@|��{χ���|���o��2OR��mH�^k�U���U��O}Йq�a3���Pde�׫S�*N�:��k��0B��C���_����IN.�]I�v-Ք�7���������ݿ��id�kÆqR\ �����|C�7�=�㣙T����)W�IN[�J|��9�u"��s
i����r�V��d��\��l�9Y7e{���%��ߟ��>[�,� {�u��ۛ��.6@ ǟ]٧ɘCp]ʇX.f��ZN$S�TJ0Jz�`3V����9�"cC2P����I�V��a�5�]z�E���U���o�ޡ�g��Y]Pj�U��������m�\M����F=���^K0qWљ �<��CU��q٫�a�<͏�z��p�o�^y@b���Wh]���%�[�*��Q�-Ywp��U��S �0�V�L��@Z�]N�+�fg�6���;k�����?�! wr�� �/��v7]P�WC��Z�W�\��vP��V�� �a��*V�;�a`�����>����nm�~��ۛc����N��{)Ʊ�>�-�.���Q��֤���:��|�gk��kl�{�i	���ϻ%;*,�T��
�ʢI|�$��FCĖB�P�a$����5�.g�=�]�ټ}:��T�*>g4���Mڣd�1��+��N]�s��љR��wg�����u_a߰ңM 4������9��uy��t�-v���|�O-���X-U�gԬ��:���!��Y[ٗg�Ӽo#�a�����hhcZ_�b^9���S�;�t��9�C^�g�w�"�w�Ri�@v�M��G齎fV�o��)$�(��}�n�>y�8M��#3��/���ʂ�a^s_|���b�M6�gkq�~�}a�@��3����#��|�'�ʲ�?he��nIs��-�_k&�g��\�1p�@�ţ������C�*1������瓃��B�S�<]���e�7ЙW�Y}�^/�%�8r���`��<65z�i��OG\8-J�˔�BW�-�Y�a����wz��b}��}�`c�C�|�'��c��l�A�;��v�֨��{u�q�֪�2%���<^��ޫ��x�=u��}ϒ��tkmtl�t'ep;X7UE��"\gfl�`V�=���!$_�r���v�T�[PHgb�\�:tZ�1�U�J�{�g�xk	�(>yu���ypDq\�	�����b}Lh86L��"u�Ax�"��`�ӏ9==ܔ�=�6�t��}��n_�E���jT�v��E���̇ȋ�S̏���d� ���aٚ�UsvX~�͖-Li���v\�Ganc��7I<���\�냈^�kԻ����S&���%Ł�>A&�,�S
�����h)��V���1[�t��{D�J����*�E�&��ZCz�z_S8}���d#|��P����uQ-Ѵڷ���T�B|��ct�k)�0�yW��I3w��ql�[ѱ�H�3�:�C�_feE�V��yB;��XJꐅj��$^ŧ��o#z�0:hk����=�������/��_ƅ�ˢ�sw��6s�jg�2(x���W-��\.w��ttq�~}�L�[G'�xG5 ��nj��O@w)��#�V�o	��|Z�;�bWi������,:"�͎�A�c���� ��v%��`�tG)���B����/��"���w{~���ya\S�X�B��9�2Ǫ�����F[zG}��U9ȉO�98��Xt⯩IT��p�����7"Aȸ~/뀠[O�}�A؃��Aou��gKZ ?|O����Qt;�`�YWU�:�n��y��I�5�y�Ac�>;!�W�}2tOj����}�E�^��wP{~;�nBe/A(�s���ڞF���p��f@c���ևd,�������OU���i:���;a���l�s|�&�+3g%D���1g��X�ۢ�R6�9�F�flɹ�1����T�)�>�0F�q� Y����)�i��;B�W�<䌸��LT�%gC�n^4�DBP\q+;r���yfj&��R>���;CH44���s�7����>t����Ԙ�7�D��ך09�:O����güc�;���uMmU&���A�J�����.���޵�D�\&��i5�2��v��漫�B�����e(�(��ǡ�So�?��Cr{�n~O@K�dڑ@u��Ko����#>�x.�~l[>��{,����~C�Kix�j*6��X=O
#���ۭ��d�P�k�1ە��u}D������f����>��Av�&U�ҋ���kZn�ǡ�m�{*�.�*7%Q���;�{8�
�<��OO7���u�����r�Db��d����>ݒ�a~�}�
k��C�f���󋞑�7g���84��Q���V�i��0O�YK�v��*��_�������&y:C��R��u�'�Ń��X�=ճ����g�����֓�~�wg��y��u��xC<��x��;uF��A�lwj�yx��X7��^�@�Y/���L��힗W��;Yb�C�㦽_q�z:�����5W����(|���G�r��m��,t���:�<��Wk4�L��NkEo1,�x�ke%��k� ϳRI`�&y]���#�%t�����Y�i��4K���ʻG+f5�K} ,���@-�f�lWLk�)Y�ۯ �pK&���9�y�7��'�%�C@��ҡ^q������T���q��$��O�Ԉ�{�ǆtV��Vk��+��/��!��c��	{��U��;/g8�C[wDk��%?_wP^�2���l�_���[G��H{h�?s�~�9�H&��rސ��#[CZq{�k�g��T���"��*<WXl�M�����p��'���Ŕ>��D/} ݂�z_���J�E�����KOZy����5e�.9J�!�6	��մ�%FH&��|^K�48Ə'!��	t�}iz�+�\G'�"����%ACa�Ż��Ӭ�����|��̏ji7Z����<�AS�~�X�@��N+R\�����K��QySY��w���U5�9>W��;P�I?�,���O��_A�ha�}}����Q�a��2F��ke��|S$�;Շ���=�|=4wu���+ÏL,��z�������L���N.�S�}	@���ҌҞ�?}�?�gG�V��ȻQ�j������&�~�9�mכvk�[ԏ���ħP	K1פ�-,l��t��e�S:f'��ȯ.�]f��Z�I���˖�5.����+?l���*�@폫�ORi�/���8��^�0�k{��׃�화n�=������bd��i��*�������׻��a��)]��~���+�ǀ�\Vt
����P~�B���-44�������ߗ�h�<5�,,��:�����8_/섄*������1�`�{͚ƻ/���I�qI����~#�K;dM��q��t;����}Z�^ǆf?u3W��u���ޓ��q+�5�`�o7h��|_xX��񥔺}�����
b���	н�|�n�k��*�3��lB��-��n�� � �uB�($�ۇ��a�1P�XK3������q�mn���]�χ{kM��G��e�����,��z�U��#�5��Z��σ�[M����J�FLۇ9����������s��`&'��wJa�B;��؍�ǭx��s�T�2Z�lظ1m|;qX<��`���'�{��V�HaF=���׆<��\M2�.�aK��M֥~��xܚ�z�~^ʞ/�!X~#|�}�z�qNq]\ú��ܟ�f���b��k��*��j��o��P�Wmt�.6C����h~8��x�&�;W=�=�8����h��#�5���`���~��� ��Й[���@yw�.Yk/*���p4���� ��S{��a�u��[r�������Y���7r-I�FRN��t=�F7o�NE�� H�[vͼ��)�@C2���v�r���{�E�;UM��ԡ�fN���PtG�e]h��2e�����B~C'f�*"4��-7UE*�$DN8[ �� [�4�M �CB�h�;�\�g{0`:Xc|G�_r�/\��;���b^��H-I��=y׺�zG2���,����S�G*z�%�b6���aZz}���ޫ���2hP�dZ썚�.M�:��*;[lV�63�������Z�;4��yn�l�W�l�o9�-�N�	Ij	\�}Z��K�N���:Vz���8Te�H�h}��u`>h.P��A7<�K846Dx;r�u��є35�9RT�{��S&�m�v�cÿ����s���,>�8�'�uf�,�i7�>�u�S՝0�����[�����z�����(�/+�z-i��O����w��FhBN�K��qM��|U����������փ⮭.�<�
b����w����Z0�gk�>��y����]N�3=�-�ˢ�so%�6/�FG��:�2)�u�L�O5��Tv�x$��ڊ(��+[i&�~��y,_:�q���w�W6e>���/	�w)�1����/WmW�y����<B�Ä[�%ո���Y����%�?r�M7tO/��N,�P���>隸gw��|�8��o]jޣ��V�����]���]����;�P_fAY��yL���5�sk7��n����ZB�&%�U��Z��د3��&�F�5��>O���M�V�j���ч6�v�����y��8��8�4N=ꔲWn�^����Z�)ZLA�Ϗ���E���4E�S���Ls$�3BA�%����Ԝ��i��E6U�p��,�+"����8��|��=�&��� �,#L�;n5�l:�8"�y�������v��]���W�{��4�u�U ����X��A�Esnj��PN�m�ݛl��G���
P�}���A(�s��>��	�n�4D�alȖ��/���Ӭ?
5����F���'C?�����Ķ�8\u������e{��^�v3��9�@�zcrT\_oG�h�8��2�)ݭ��3^j��u0�Lj0�k���q]�Ky�?�ն"窯� #�W&z���R"6�ɗ��@S��<)����A�<"�w�>�^��$�u���ߺ�#�+
��l�CCA�5���9�ulWx��3�ur�Ӕ<�d�-���8��Зn|�}#7f;�x7�MAm���5���i��{����H�M�#�����3��.�у�������Zjzo/Kx{��x���i�
Ck�c
���&'��u��_�V���:�C����jx ��7ހ��3�+~\���;���6��������^��h�4�}��Sr\ꙷ�����7Ƶ7��"�%R4m)�6�j��F�����:N˹�k\�΃��f2-�E�4jI�dݮ�I'h��+5���o^{^�yg���M-44����{�v���T�C�_?^G�]ҡ7e'��84��d��>�-6��йD6�W<�ݠ�����˞�7����Jq�\B���Ƞ�ܤ6W(�y�U�O^����B���I�ð�}v�½������[X�� �F^F�V�w�1n�v��Y�{\�3����5�@���X�aΠ��^V|e�3��o�� 8�� �|�|���,�6u���T���iP�����N5����{�M��B���Ϋ�Ҧa���0]�Y#z��1�b�D����� u��FF�G9���}�����v�ja�M��NXq�^n���>�-���^��&X�h�u����S����O.ꯣ.��YCO^nlcMsz�����c�TA���	����|�]�b�1��=��h��k%op�mK.�N����A�&`B�˷��:�/��&��x��ބ^X�W<���{��l+���Sɳýi�Ғ�s��;D��lx�*���z���.,ț0��k:Նځ���c�!'k���*�24�..H_=��7*+Q�\���t�ۦ\Tk��6�����lk,���(�>G�qu���������3ݷ/8�t/�`��w�p�:��M�����F���ȇ	�.O]�^s�W��7d�Э�K#�t�j�%�GS�n]U��4�4444
�v��y�w�Ϟj�j���=���uY�@T��(t,<�E�\S����(��q쳂1��o8�O8�x�\�=7K�nu�U�����.�-/N��\+<Y ����Y���e�͢[a���r߄D�T���k�aT��k^=a)�)'5�)��S�gR6D;����\��dc��6w�?������O��։��s��(-��oK��������4-�l�n,׹7r�Op�N��_�O.��4=gE<0�O�..-�_i��C���>JG'��n��=���8�^L���ga�g؝&y��M��ף�T<>就{ˑU�4�7o��YvIF�֩��@�[p*�<�(wv�8��N�N|�8����d��'����l�Ϲ3�Z"<j�;��RhV���/j4̖��in�2-�r47Pܡ����W����Mv���ŗcϦ�g`=UsיW������rٜ6|�4�滄\W�7w�k��}]�+�^=[ռ4��;'5�e����U��H����)����l:u��	MA(�u`wJa�Q�Խ|�3��=��V��nE��u�^t�3��Y*�9�-���	x��Qn�9��`�W:�i����՛Iaˠ���������ǔLM�i>�[��`���rT*����k7��$��\���pNɅ�,S�kup0W^�{Ȭ�{�bέ�~o�J�܅0�Y-��c#�baAI��ϊ�{"Ǹb�٣�q2��'E1�kPխK��W:�ÈhV������w5�� �6�S�bF͌�xuPu;{3����|��pF��9M�ymi�(IZ_46��n��<�Tʹ�4�S�g2�����ZM��,�0m�JR����;��8��R�[�N��a,՝ݍۆ��hu�����rP �#zr��x��k��{eh��{�ش���s��7:�X֣iu�ܕ�K[J��ܬP��.�[�_a8�\Kz��ِ�R��,*��Vέ���<O���r��!ɇ9���Q�7�����;|}�*C�5���%�^Z��W&��[w���dLZ�u�ű�Jd��鋇;�lˬ�+B�/V�d���J�}����]��T��oM�]㘦�-�8�V�w����}X�,Z-���Fv	[�q��\'n�H�b�k:�J�9P�ѭ3�+u�$���g��Bk���/Js��%�sp7�n�pZo`����4�mK�vc��-o*��[������ա�i��X�lnm��e�Lu2+z&���څ��m%_M]��m!��	5\����Z� ��Tk�J���SIT|HƎ�QS5B�RhV�I<RQ��=!�U�`pd�S�H��C��Y��n���U�>������[�S�}$��|2�9������oWβ�T�N霙�zy{��ꌭͶ�x�6!I���]��
d�y����)N3��>����q���3�u���Ԃ>t����1��ڕ�;qL����0.��
�����+6'�v:��2ı],���k�5�a���t�Q�zU�Y+�Y�x*t� �ݲ-��hua�Cm����Z3_�(s�Fv^�9:�EZh*��[3��Zn�����s�Ưzf��"���P�<�.��d
��c����բ�yvĜ��=ו�`j�u�Ǚ����aBvzo��{0.�c
�u�J����2%y��t4˩#�F��of��C�`j��j�-��q��S�]��I�Qp�P�r"�'Κ�f��]�E�	"U��sOVp�9��=l�gqp�Q^i��g�����P諈cF�~�^=L��ͻ�Q�K�	Zv���� R�z�^Ց� ���Z[3����z���� ��_M��v�w#��S=<��
�j��յ�K��1oȝ}k)�c�S�5<�0�7���=[�jZ��p��}��X��}N�R�U.�t7\��K&{{)��:��ŉ��;�#7�1�AA~�RlEp�8�!�Ÿ6ZwiUb
:�F�"٨d-IURJ� �!��˹��B��ؔ�[B�����@�Kr$�HQ�f��	[�����H@��41��D�E�j4(B�~m[J�E��_mWLb�-wq! ��Q�"H0��㏮8���8��q���6����EA�4�-%�����o2b��r��J�҈�m~o��ׯ�}q�t�8��8�ׯ��]F��E���h��0]�����-%FI�����}z��o8㎜q�=q�z����B$`�)�3E�#X�~u�F4~M�L�f>v�+���wqgv�%��Ѣ��0��T�Ґ[��'��(h�6������a�X��+��A�	F��Es���,32+��*2Q{Zmq)4E��#H���~�e���	�|��;t^W
I~��Q�e�ۖ3���ن��Rh�%'ZW/�t^t��t�t�o������wߺ#�Lc?3d����~t�����4�m�)U:�限HN��kr3���譭�8OFj�%WJ�%=#)Ǚk)�m���m�z�P�8pt��@���R##P�
("!�%U޵�V��.Uޫ�?�����@�A	��mͿx�!2��-���{w�Hqm �|���+`>gݻ�O:Ĳ�����1��jk�{����PWq�P\3�!��$ds��EϹO�M�O$�o�s
�1�r�
�Un��^9/�>̓�QL@�R	P���܂����?���yQ�A{풁EV�;Ms��9}�w��z^��8����w:<�zy-4<�/���}�m��xUã0��fk��&����;�O>�<��֯����/B�5�(wW�/^�Z|���ې:5�Xv"
{��z���s��~����L�n����qcOO'o_l��/~� uT��6-��|����5�[3۩��a��%� Q���b@�{ţSu)46�x��pU�^�y(��@�⋺ҭ���VI�£�x��v���<�	�?uO��ΦO�R�e�ur�?����w�YF��rC�O_���Vp�BvKaZ����'��	gM�/I�-�������*�b���Ր�ա�6>�~���P�ۀ΅�@���,�_?�!�\�1¼F�zc]3�y��㻉�B����a���K��"b�S[�л����t�hqպf]�8�ȶ�EZjb�b^;}� ]IX-�K]6��U�׷-��)6���/��K���)9ʄ��>ʂ�:GX������s�v�(,��'��8��Z��̏�����z��ǜ Ei�/�p�u[�|��wZ����� ��9٩	|w�_j���)�bK>&Io�f�]���)N��T�0�K������A�t[n�rf�ky�c��㪹�¾��X*�A<-�Ckeޟ��-��ʅ���By�����3��Z��s�o�jg�ùU�O�׺���h���.q��^�=��>Q��P�&{�Y�IZ�s�]�˚��Z�ޔhU(8�ũ��|���>��@�O�]G�cS�)�U��wϼ���U�]e�#�6����w4	dB�\�Xc����W�;3��A�}�k���4��7*gx�,欬�ffw�L"��J�w>Q̺�y��I�jF1;w�=cX��9��c6�LwA�H,:�C�k���N�R���=������މa���W��"���"��Ȝ�o��.Bq"��LKmz�Q�]�O��so���BO^m�q�n0n;�3:d��[��C���v�@3��y���S/��l��.L��FW8��d���ђ���Z��h�w(�q�����g;�	�w�e<tk�����oc|�ll>Sr��?|�rύ�������rZ4�z�i�qޭ�-���k��/�S�ʬ^���ի/6���c�!���Ӄ��n�
�"�^f�i����y��q����=᫶ ��e�}��Ly�z63����="p-�>h�{����}�
��'�j��o�/��<R����2�{7�����Z�r�G�q�P���i�>7'�K�>n�[~��������J.�9oM0������J!�7�DI��!C(��E�b�7�W�MN��#N�S��M� 6>z�ϓo���)P�Y:w����++`�%\�d����ZF_���5�[��R&�p���|n�Laz���~����j�Q3��8�ǈ�[�K��~��-�I!�9'ν���/�C1	�!.��23<���zt[�/�'rbˮ ���շ������U9��Mfo�>\Xx(�'�C�!�>����5s�1Y��ʹ��{as�|�}wJ��mB�j������7�l�W¬y��[Q�qph�,>�Ez�V|Wd^[���VK�������ߒ��Wʅu�Ra����3��m�Vp�ʹJ����s��k�z�uO��ޜԔB�����qb*cg�4F��)��;��?B��8+��@�����_3���5%HtѦѷN᳏:�su����=3r1X9-ow��<�����"*�1�\p!�����c��3�WBJ��/D����žz�-��7\�c�W>�t��du�BH-hn��'��zޫܔ�t����-���׏��SCM44��r�y�f�w�~O���&g��S������f/P*vy�y�e����.{��b�_��F�
���S�/��������Xm��$4q\�Ku]x�hɃΓߩ���P>k-ᚱ����|䷉��\וɛ�̤
OT�_���4����;�G�9�n/R��^�yR$�a*�kϼݩ���L݄.r1�n�z�x��ЙqS^m��7\װ�1��y<�ۧQz�`���|��Ox�R��-�ZN�c*i��k�P�3/��:��Ҏ�봞'�|�=�|xF:�w��d�&sT�~W�Zv�N�l�RN,$���r���������Z��ey⁀��f8��h��^�X�`Zh-ހ�o0��sRX&��)�k��g�Y����S�g]�w�1�YWݵ�x��b�
`&�،��Y&�=:F��z�	K1/K Y��u�jkª�޳��o�;�YZ�ZT4y���J`o�R�|lKx}���р�RT���E�̀���G7��-㚱�f�0��hn+f{���'I��:��ǇX�:��L~�ݚg��S��ϲ��q��I�Mb���2ͼ�"O�~ܛ�����v+A�%�[rۑ���4��u��%�08�0nJ_��ДP��;�y��'�ު��b�-Cu6�ɋ�����^Y�u��}�k�������n"��ˁR�+X�ve�Om�fF8��^��I����4���SCHn�ߚ=���mV�;�3<���\G��9o�wT�ݙ��宝j��(S���G����S���$z�~y���q{ފ0%�pȶ����j�$�ۇ��vm�`��["��| c4*}�1�!Yי���oC;���G�}��U�#���Ty����Фb��=[�tooR����.��,����f�%� mVx��~~�T�~{^�KC�1<�c�y�5GwP�:����bh�T�w������w�V{�S�V�"�Oz��cK�8�v}+L��ĲfG�%�Z쓖��(k�����u�S��s�p�1�-.��=I��b�`w���zc�0�-�9�Tx��O�MBb5���W_qt�H"h�5�~B:��n���8�U'� �֥M�ķ_�_��N)3~�J3���t&U�<�Z�Ĵ�g�>nln��n�܇Q�]����Qp��0b:��:���	�t��g�3WP/^���+��/@v@ 2iw�n@y5����zA|Me���_�F����v�p�[�{��,$N�]���b{���:�F]�����X$~��_Bq9�unu�ݗӋ�rVe콬�m���ލ�:{:Y�����}�V��.��������:p�Yu%�M��J�g�U�L����ڎmX����Kлx�{���f6�J�	��E��>D��<$o|�Zx�����8�y�������8��߽p[�^�/I�K���'�r��������ě��t-FW<�<I��*��}˹�p��(��\a1���>k[�7>S�j̹��0��,��f8YB]J�r{�ׁ�_���X6!�1��<�����#���b,>�μ#p3�������M!�^S�a۽&0[��DT>�ĳ�p셸�fI�&��n
����~�z̏`���7g�0��h�o�:�����
�^��S�K���S99���Y�x��@�孿��|�*9��B��q�5��l�;E�;\�9��qj/��ǝ�<L�7�cN��?[E�I�E�����\���O5�����]��y!wV��l�q�{o3�#�ǘ�Z�Oʭ�GX�/����$�����������u]0�H۷EY<c��?wt�+�ޡU�q�~U���)ZPu
O�]�k�1�<;{�C]�9��z�L�����1�����`} R^�ۙ�wO51�r=C���P|���H�\����US�ν\]Fi{���$�8^%�c'r�g�|���Ҍ~
ݥ�M��_HZ�$����yٽ|�'e��;��y��Gk���NPH�Y�{��#n��uۈ��q���NT��HZ�'Ue��,���x��K�6KT����7	8�iWs�uˬ������#����B�x�0�MOl$H��P��-L��>h�h���.'6á6��&�z�`'<:<��m#4�W[g$�Z�^-s���|�v�'�4'�6����[r}��c�M
Y�#����'-��K'jz1w��ښK��{�v����gh����D�kvq��������Ϟ~e}-�f�Q"�vm��=�W>�U>Z���,a ���q}�Dz���00��Waa�YmF��T`���7�����Yk����F�l�����#a�h`�?1glnN�ҙ��ߦ��27�_3����d��pl'3L�j	i*֟'���_
���ӂiE_y{�8��_�9��pn��&h O�a#�8��jFbS��ŷ
q0�}"�^��9��~��!�ݞƪƩ]�7�� �}1𦷪ڣ}�%�S�VWi|]���@��(v�%�	`o.��
Q]�2m���./qKO���	>���6��<S�0TS@���W� �L����5�x���;.�S���
Y�9��k����n:��/�sm2�tn�w�q��L}��H&$��x�R����xnL�L��m��Ύ��\�rOT��*s��͈!��|�fe�������]5�N�n�����]?}^��^�.h�����7�>��n�ΞKӼ
X~�{\S
����6�l	���pb�����>�0�{��R4}��k�j5��	^b�'�/枬��m:�����p�7r�i13�-f�ޚ>�bP�U��L���]=I�5"1����K�?����zR�f�c�c�#�b3L���8Gx���K��~;�Ʒ<�s�C־&�~��ߎd��'�x���g��U:����b<���m �'!�2>���E�3g�e�`&��m�=�w,�Ô�W/��\^�J���ټh�#0�	X>>������e&5��n]{J)������nK;�4�]�cwUp��u�$bj���Ң��ǖ��T2�~;Y�'h�q|��<��]�|����闖�r���L�qU'���^`'�r^C������KԼ��)w��xs�6vNO_��L�8��]I�_-�ǭ�
,K��Z�'�=�!p�ꏎ��y�
�A�j�3��NS�	���{kPXO���@�c*@`r�us���d���4'��Ių��y����P)��{�^���Ql÷\�m
��,�Z�^1Z�ݫ+�:����(����̙��;�a!G8�S�)��0�=�}� ۓ������[�G�]R�.̪��Έᘈ�ʮZ��UL���1���U��.�M�4q�8BDw�}�秿Tb�C�#칆	�s�����k�S�7��V%�Θ	��:��Tc��HgΠ$���_�o-m�����n��z�EbS�J��R9s7,������߅���}�9�&��$����Q��dWΝ�v�BB�uϔ�pR�?���ˮ�,gwI��~J��Q�-�
���1�W�^��xNR�G��W��oM�N�f���SW�c%�ZM�ԟ�w��<�2�gͷn�ڨ�y/,� L#C�8�������u�㉻PƖ��c��q>�њ�[V�ʽk(*	J�Y��'�1P�)��a���}���u�	Я�m��1��=k�.�2|�t��M�܁�P�~�r���l{�*�s�Qj��܏)xn���4(��B��ޯ�~�6�𱏢i;�3��И&t��R��Zn+f�N�ƶ�C����1i����������,��b�F}�<�j��S:��T"vs�j���)�.���(��0�Ơ�ۢ�]��Ո�EQ���u�����~Jyz�V�[j��z��7|�諲X��}��(�E�V��n�}��V���m�Ʉ�6�M�܈6zf.�d�C.��������wi�t������E\���tB�''�r*�w�/.�(i]]sC`Q�t��i�Tlާ�r��&��m�V3߇������0JE'P^�8�wL8.�����Ss��ڬ
:jw����F����c����e߹o
i��'z� 3��9��]j��-~�Jeczy��Ĵ��-&�#;��Ix�BՉD����4=3����a�;�����R��5�;��s����CYy>���q��dJ;m�;1�(�[���]�j�{�]L��?�k��N*x��Γ�:�C���j�":�/5l��-�O�����/�4�J{�b�04Mڕ�Gx�4���`��-S�G����9���i�c�m@���3�ݏs���&:���_TӞUհ[�G3���Rk�v��kw��}L��c�˫g�7"�'=~�
D���R�ׯ�0��<tQv]��N�O4���.ϭ�(�sL/��l�����!PJ]���S�FDS[��� ��,��;\>ŝ{�����jjO��o]c'�.�P��ݔ���A���ݼ��-=x���ͼ59m
x{ѻ�o'�����廋v�AØ4�`L�Jz�ѫ�
!�]9�p�ܮC��7�����[�t�MSwX2�S�����SO�*z�+,}��p���\�05�fu�Ll����ySW�� ;S�9���c�1��UǕ�Z�\���{����cWK*���f[��U�V�tI�LY�\T�0Ցu��������.vT��\��Vj���=�,������p���d�5�\�q��U��Y)WZpgv��j��j�^�)Ӽ�J�%b|k�]!,	+`�M޽�w�6&y�o��s��D���	�V����Z�z��m�3q�K��$5�w�tѷ��x7ǊMXR���[���{3�.����B��%�ו�CtK�/%٩�m+��*rn`ڎ]ep.�~pK٣��o]l�>��{�20�Y���\p�9�21��[�4�1_{CxUK�A�nl��3{���RL���^v+�ŭ˰fg`�TV�rS)![k����n�J�t�	��v|��0X��\ٗq��I���P{G�g}|�MFl�����3���n૓K�z�ŏ�1u$������߯�3��{��g���
�]dt3k����CIV��Y�V�&��3X�H峯R�����IHQ�FΪ�rZ�=,� �[�Q�j���[�Z�3��^�� 3*�#���G2����s���n�s�7tM�u-����ޮ��:�q���l� ����G�w��l�ɩ��>J�.0�U*|)*����1�bZ���������~����^��/e%&��)7y5�l��1���	����]�Q��+V�9����nED��v�K꺸Qդ'Z� Y-�b���\��/�8�˭ս'�WX�L��v \��X0�]v'�N�������[Cn��.i۪����\��K�� F����wMWr龖��iͱ��5<m���x0ݞSi=O�y��g`ջj[xH9��������s�D�� ��j^7��6��-�\$��w�Rw��WQ��dгs��2J�����+4+�h����q�[�T.T�x'3�lZ�
R;ܜ��٣��ghw����,�Ż�$f6Y������l₊b���X禄�W-��}8��+�:��D��h�:Bz�s��X��������U���b�3}e}
fۺ_\��%l��6:��b�F���O.�x�[�^P��A!�&�Ⱥ����*RY.gpb�^�S������L�[4c�Il<��6�d=;ty}�F�n�U�šl������lGR���Zn��Pq2*�x���Ux�R�Z�e�&��N���ʰ=�	���z�l�b���8�u���z_(��CT�.s���v�gIqt9����>������߿����W"(�B�ܲF�c�?:��ע�d���x�Ǐ[x��qێ8���i돏�4BI!I$ME&"���QE���I�\}}z����o�q���=qƞ����B�2D�@�R5S�n\���３>]����z�	$��v��׏[x��qێ8���i돏�BBeT�§`s��7�t}�u��&(�aa(��v�t(Ɠd1���<ݙ�t���o) ��A��.F�#b(��rV�ܓ�\܍��2�i*"4h�Y#o�i �naΌʉQ]��_͒)"�ܽ�Z�yFг&Ѯ{ݲ\�ȝ۽��W-s�}�M�⹀��s~���墈$Ƥ����g����y�N�N��j������(�	�DUQ$�A�Px�uG���i�4��Ʋ�R��ą|�Zs�)V�\.;.J����9�r�s��\�2/rM��+[[�O���>>���]��c��j��>����]��(��'�v�*#������nfx�xۍ�]kt�Q:+k��8�z��[�=vg��,���	�>�	<�@�|n�����V��*��V�@�^'Ϻ�ܦ��w�U�(����eyr��T�-��\��b�F��<(w�f���̓���J~��ʼ�W5���m���<�f;I�=O���>n���f	���͎�g��Ce:a�z�K��A5�}ώ��u����'�0,��}���Y��E�ȁ�b���;�È����za��=�zPZ`[�>���n��5�ۏ�) `Y�g�YYI��a�W^��@�C�XX���#����Ruõ��(Q���mH�P��b�"���gVh&�w�(y�� u�ak�
"��6��1U�:�^����[�j���6X4���z��=����0��z��>�U#+��?�c�sTO�k���ŷ{��Yq�'�����^p;�%0TƲװ3�3^��Ǩ�\�v��8+��uX�{�e7�uz���x�+��6��7p(3
��xz�"�B��x��:@��y&���,t/��|6��݊r�.O�2j�)��Y���9pO�Y��@>�jތ�![��sy��8W^Y.�*@Ԩ��"$ *�j�|+��B�}�eӔrG�Dx?zx���{��V����i��K����֡�vW8V�ac�@��%�rɧɞ�������{���Yw�^<�&ov��(�f��c��sq#$6<Y�B�LJt�����A�;��xv���5\�r�E!"�$GO�t,�W�����Ox�!�����7��}��w[A��'z��84v�����
iDN�����^Z{_rW�:��VE�v}�b[�Jt_�Г���.�Y�Z��Z��.U��3|��]�ũ�g��x���P��M�k����Z'����u�M��7�������@���w]�?:��6{)�^�l�y�����u��n�ju�;vkK��'M�"���>��v9�z��Q��L)��j���S�=m���9�s��Z$t��Eυ�Ƨ��*:�����6�D������GJ���r�þd�,m\�a�b�.{��� �xt� Q�K�>�>�l�g�]�1��p0%9��s�/Ku����N���vj����a�y�ꏧ���j ϥl�{���F��F�~hݨ��/Ʋ]k��77'�d�K/�D�S�`�k�|o�\˔c��,P{6��w �YM�҅�ŝ���B��HFϽ��a�udUԺ
�m��i��)�:&3K�7O�Q��o7f�]���Ӕ�T{@��iV����}8�E��һ��y�=�m��(�P7�MCM��S�(E�/��<||\���˫S�~��țN��Xۮ���q���ėׯ@}y�{�o�A�U�{�	��w�4Rm�mq�9�a��<�Z��y?s�K�`��O<]ѕL�yv|'��.��n}>|�V�%��c�v��OH'#��h	u&�5�3�^�\�<h��I�@���|;(s۩�ZT�ܮ��&�kye�[�Ԋ��)�I0�.}�	=��,;��m	푙�R�h�kM���#���"��`:O"�\��������S�H�����3��DGE�U�n�՝�<w��Xg�P�y���E-�Nb��.D����M�@���M��J���0̔����^�ݫ��hvr��euG�(�Z�c�gTjyY;>����ϯ��د�Ӣ�s7�T4b�q���A%Pȇ���&{C'�"�<��Y�g&?yc����U߈�?��y>�L��c�
G���������Z5��t�f.u���ޛXQqMK�O'w���`��tm�sؗ��Sa��nC+�
"�,J.�f���D�����u�m%~>��l��]q����uYm[���R�@�v�w9ɣz^��@�ov��7q>yK�0?<va���L�3^m�͔^�K
/�D�9��^�'�[�oQ��<	I������;�Cq�a�5��8�
�����W�y��_s�J�Y�~��f��.�ۺ�׌DsR�29���
�԰
S��~(c��I�\���W�6��%��*af�5�Ϻ�6�����g����r�<�҉�^"��\s�����~4�ݬ4WT4�Q�W���5��xF}�K�!�6\1���\��������]�)��`��L������̈́Ls��t�QnV�3.:wO�c�(��~aݵ%?V��Θ ��+�_�~��A.|RM*,xy�F�R-Mu&��L��v]i�2ف���D��s�9�&���-}ЙV��j�Z ;�P$-r��U9��0m����w�=������!�\И,5�ۉP�K�,0`�s�twH�~�[!�ͮ9�<6Owy旮�O�צ�<�=>�@��[Q�:�U�f�X�[�6��ޞ׾�I�1z��3i�QS�����t2-�NƔ
��[�<^1�rԭt{\����b�aS!���4���T�&EWU=ﰿ�#ȗJ'�w Llv`�85��
{���}L�,p�t����q���m9_9�F:sUq������[�9������b��Olx�JTo��ŁȈl5pr2Δ�4���ܹ�VT��Մo'��10h;3�f����#�3�� �M���(���\gcD��ڍ�v蜶��~�x����)�Q������~��֟�H>ke�o�U�����Ul�&�|A?.�c�N��ev�f~j缩z�M�����+ 6`9V��wa'����)v���S�c�[W����"��b��^��o{c�0��a4��C6���yX��G�-P�cXiꐅj��&�->L;�M�5�}�ů3ϣ9������TQ��]0Ώ0��ɞR���zl��o1�A��[���vZb�A}
&b���>܇��gS�9���b�|i�0!F�����0<#;_+"}>��+�Ͻ5L���)2�=A�p]^��لP��V���L�$Dzs����c���1��ĕ;�x��"�����'��	p��?�i��=�)ǀ�]}���U��
V�t�~B�ݏ'Kn5F�ƨޡ�L;j��A��2�S>9w��{�����O*涸7"NE��]�5���땽O����*@��|*5�H�%ē]]ρ�u��ayˢ��û�0L��1��[P�ő�� �&��i��w���az�om2Cm�t�\}-.�ܷ'��_9��0W:֪��X��q�����UD@���Ɓ�O����]/.]'e�|ë�u�#t%���}�K�>�V�f��8�.4ӓ6��3�ci'�tkr��sÙMc}BUQymLoJm��Y2��L�q�UC�Hl���V�}�+������{�}&��-�t+�L$�C� �����O���0.����ڽ�@��y�\:�L�c!����*��z�S\>��^���O�VQ�c�/�ƽ_-��PN.�0\�foG8�!�D��\�bİG�04�z��WI��d���Ϡ*�[�؈(t.��\�>��v�����E�N,]:�x������	��>N�D隯��3�w�g�C�X>#l$w��(���B�zESE�C�eR�a&-�Z��6�e�>ܞ����4����Y1dɤ0p�	ST��5k�x2��B�)m����-�i���9�5iv�>����JOB���1�f�<f������}OB��[�}򯚣~]���}�,���2��׽D��v�k����۽ᡸ$O����z��y���ׁ1 �vC[��=���[��ث��}�|Cw�k2����.>���'�W���>�i߷8}�8U�U%cP�}�R��˹��Z����;v�N���
�M�a5�u�1�d��gO����.��5��/H�۩��oE]X�����x�m�j%颦U*j|2MΆs�5��S�V�ɼ��[�ۥ�j�q����(Cf�ڱҷ���3W�Ge��G�b15�o��۵b�S�JtJ��l�)��[�e��u��,=�a��(�T�6Ɣ�*A�RRP���޿��<|}p;ᳺ�ԩBg��!�^����Xp�XZ�����خ��*�'��Sq���Qo臁���m���.{����!ށ��]}�Z�Do�"?gH�jQ���B�+�qk�XR��~RL�Nf����F�Qw���"e�/y�>�S�!��͞��:�7v:v�j���O{�ڧ�~i�U��f�xa>́�8�<�>�zn]���W��#&�sz��S�QM����j�v��Hė�a����e��A�{��-������Pw��p��h�����j��t#���"|<�A�cX��8�!x��=�MViTt�Gx&�xh����A�)ťҷ�g)M�yu�%=��iw7��!�t��wꙦOot+9u��\��.(q��@�׍NH��Џ�cg\)w�?�f��W����*#{���Y�@_I�k8ı�Ǧ0����ȩ,H��l'3Z�<P;�g01vn}����R=��Wi��Ei����C_|�Zی��Y&�^�!�(������`���;7�*�j[�x��P���e�f�uX<���Y�{�����ED�A�*3���urN��6�?�Uh!�n���m��$�;n�ӑSd��j���\M��0ڃ�]d8������"��W��7�傕��N���ޟ0�y���	;N�;�l���	�<��:���G�5�+�}�O��a�}S槕��������"�#{)�9<���0X飄Θ��	|*��Ja���N�;X�+ìI�_K�
�/����j���3qn�[�zkm��ۮxb,�2逆j5�vn�x=�띗��E���6�~�rs}�ȏ���V��:EH���mCreG߄�
�>�6q����g�S�Lo[�B֥��OH��ϡŵ
H�^|�ۻ�k��P��;XFG7P�T+��J��WU�j�S�@�̿p�	�N��=[�S[;�M���Z������^xf>���ɓVuQ!&���w��k�o?�tc�{�K����a�f.}eY^PR��������VTc�Z��Bc�gq��:k!>�i�C��ٜN�̢Ys߸�2����W����v�T�g��tw,-��X��r���і/5���ᣳdl�{���9��X�S��<^)��H%A�MA�6�5Hu#��
3�Jݧ��V+"��s�m��wf^���fo�4ɲy8��&^�Q|��ЙW����PB�`HzԅwƳ���W^�m������-�wf��'O{bLvMY��S�!R���Y{�ym��EH�6�}�k2�Ìo�M�"ViZV�ݝ��Sn��#8�@�,��9�|�������|����ԯ�������r��{���g>�N����o��L;��L XkN�*itR��}��	{���T�.��Q��^O�On��p����a�����Þ�'~;��X}�[S2F{]�&�ia�1�s�[�i�[_4GjA��dr
� _���B�����C�`�F*]�.�Xq/��n�n���Vz5tz5�>��ސ`
�g`5y���}�\¥r�O����kU����	�"
�ݬ�~�?u��M^H@[A*���,��������2���ulk��Z9K������ˎK��ɶ׻	=y!%�_?� �jo��x��ğ���PJ���}Ϣ~���5Le~����e�z�<��~K{��ջP]�A�\�ԇkƒZ���=�'�w\^▙�4�DF��Vt�fy;�窌5~������^
�ʫ�n4�~Ż+�Fw�����,4Ws`��f���Ң��D$w����]��Z�1U���Վ��#+��P����8u�+2��N9�
/��v>߻�b�R��J���H�94v�U��A����1z�dnb�S:Y>XY1���p�����K�3)Q��P���VR��[��v�Q��n�yW�|���T���OVܗ�S�+����	,Ѣv�������Ҥ9.o��x(M����XF���{�F���>#�����3n�Y���\bY��N�7'K��u��U縰�P@�<�RĠ�{�{<�AN�K[#���۵�[»�(�U��.�B��Aǁ�7O�������/�%E��"ڴ�Kn��q2$��>������tv�ň�Ni�$���v����`�!�HXx�}/�U3k�k��)���M���z!��� �o\G;v��5��zv補��O:��'��[*�N��nƽ'UU�r�������8�4Ȉ���M��I�L��7������L2�!�F+˯��N<'g�>|�v�t�ҝ�4�=ԕ_�b���:�TҮ�U��4f�@���R�	�F�_� �Z��Q����_c�"f�����۠�hO�=�
3�`���2��緬H�X��0}>3��6Ƥ���H�S41����k0����-�F��7��T �1�B3ו��� �>�U��čH �j$[�6��7�.�:��L.cjWi�辔���kє�E�͔������-�����B�:[}}f�t���X��.ډ=�*2���j8nt��A7���Ŕ��R@���'Q����W������:έ��K��ݬ�R��Xg���iV�C�T˕ظ̵��@�
(�Q�J�F���S�P�rm<��8f�G��wUU}QY�x�� ��]��I �}Tu��`���R�vM������,�v������e��7a	Ib�ґ��]e�%�cx�&�r ���V����6��(��%��m)��������v�Wl�GQ���n"VMt��y`��mY������kFs��Sx+�����fe�dX��v	.�������\�U���G]�P��1.�rC�d8�m<��ܗ[�Ɋ`�j���iW�om�	r�[����M=:����W�J�Z���2�a�
5k%�L�yR�n��O�eS����
w+��H��]����ĨowRR�v ��C�0���YkP�u/p�֨�<���P�0�5�/q�яC�X��F�>n��6v�=	QaW[�}�l�I�Y{�Wi��L]::����d&�K�qQ��f3�?NW����M��9���`�|�Q81HsU�6᷷BՒUiT�`
��IRn`.[|�vȬS8�b�X4�*�ŷA�.�Dqi�ْ�0�"�g!�x�3�iEv�H�����4�� �
��L�i�]ۻ����끓�G��vA��!)�IU�w:g#�rn��V����w��%2`�R����J�f���(V���[vo-ɼmS����E�t��$m��s�GCXg�6C�
��pU�N�R�s��Dwb����V�MkU�+����m��]X�gl�#�;z�VIQާ_��7{C����V]:�w]E��gH���[3.%w�:��O���g�ث�۠�v��F�Suf��u���j�CŚGsO9k���c%�M�V��iNT�m)t.�T�z���|�X�9WoR[�8�.=�;^��6��>}j��=��F&>�7c��W�~�֓�y�E�}"���1Zn�X��n����Y�B
�L��}.��-.L�.�SWu̎�}�����J�>Y�Q���T��Ji�Zu��%��:��R�E�lˠ���H�f<i�m��l��l����Pr9�ǣ��"��wS�V
�Z�Ȍ����K����J����Y��m'v)>�KY[�׺������V�]WKsn���{�"��MgLH<�=��3%�IT}P]eè��t��׌�ʢiY�G��:I���m�.βE���ǉAL6ӻܼ�����f�ʾͩN��۾����̘��m�Ϊd�eD"�j���
��8JCD:tӈ��f})2aM�HLF��(�$mcv�����|É	D�S-I"\mBC
�a�cI�H"ݚ��PQmGNB)6��@�*!1(�,v�)D�d�j�{�;n_ (-�vߏ<ɠ�!��d�d�G�:|x�q�|qǏ?C��nڢ2�*���2 �.We�.�up��n]�Qt�&�EIUUM�R>=z���֟^8�8��<z=}v�j.�!#'!WI�A�޷��y\�w��.B�1�����֞<q�q��<x�z���KDdRE�N�jqnm�W5��y�r}nc���B��sr(�4r������͹�nj�3��,r�4���,mE��k�����^\��n\�G���[��gp�[�uyymʒ��ܯ#n�R|k��ܶ6��vŒ��k�2\�l����#|nj�Ӌ�5\��}��{�ʹnU���\��m��QҺ_J���h1�Z�����J��\��F��P�KS��O_-��n;V����C�YU�c�b�F�幷�n^�mA����VB'SXd�N��mG���Bk-��b�m���N���h���<|G���x3,5����l��m��T*��cߢC��vx��Uf��&Ɉ�p�'z���=;�LIA
1������
��F�7"���7C9���E\�y���/I~襥�M�qΠ��5yvG�B+/֫���>M/cdP���/����)�;�|IY�4�շ�d�p�*�@�PI�d��{���q�z'կ��Oc�W�q�;��Uw���pm,�y���Q�I댪�Us�4�eEAG�m*m�+1��L�5�h/�c�C�tWnx�,�wP~��!ӥ��sy��;x�����Rd*an�'��@�:(м�Ńe��+{KFUZ$�V.���r�moVϚ��Fc�Y��e\�OaKZbh�A��W){�ª0�٤�m��;K��2���e�G�^�$�쎾㾄m�^3����W_��1*x��[�
:��8��M�͙�JԹk��~�:w8�@��z�xm��/�MK�u](��Nɢ��=�o&#ZH���<�t��N+�|~S�=QP@���!xoE�W������NVb�	E�[Fp2qx�9W�[�Z����Qo�yK�*9���+��fm����yy���<�`*u�f�bT�3m�a���0oQ<k���#�<�lu��ʼ�	�c�d�"1�E�Lvi��9
��,��%-�cψ��>��/���{�'w��
&��QY��5\�"�j�*/�����0���4Ì�:�IS;�;�e�ۙ�SF���8q��l���*�C{Bg!�,��S櫅2ݓ�����N�ށ� ��$��.��)�ܗ�
�H�j x��f���U6U�[�㮴�s��x�� ;��BBI��Mys{�d'�\�/\e�xh>ܤ�����=���,�߁]
�ʞ�\�]�T�Ǥ�u4�׭W�&�3XM�TP�2uI�Z5{��fFX�12�|㕡�6|�\R��6��!�4�?\�	x=�L?���,�����_t�{p�����%����6Yk�����)۟Aa�r*i�����d��od��wI� Wk�kB��u�O���.�e\�nL���ydW8X�ۋ�Ա�S�'hc!uM[�Wt�
YO�t��9�|[�<��p�B��{��:6��{;w#�4�-y����f�fʰ�GC�}�c�z0s\�u�g7��];���:?����> ��߷����/ߞ�2�m������A��}����lW|Q'�^�]����)5��+	�!{o�6y+�u{�}F���4E���
�����7;<ךʷ*4�Ǣ��g�^��jH�ʹu����������5����nYA	{xm�I�CF8�u�nY����������vs�:����*��,ߠ�Y���{ۜa��kJHH ���8��`�Ƽ8�^�����.1�Wd���MFB��9�;6L\Ŭ���s�}e���p�@a��vh�U"��/xI�u:]�ƅ�.�U��m�މ8M�D�K=t���a��#Y�<�Q����x6=�ƭ
��h�Q��'�EP��B��a��ô���32z5#�B�L�ϡ3�9_[Su}��Πv&E��9&%yU�����-v�s3��t�M�h63B�v�J�Kn��M�P,Op�z��p'+�٭�輍Ԓ刳��%wq����lk���������Je�LL��Zc�cs\��7�k.��4�{�}ɞ���{IU�����h>�crQ�i�V�>�uɁ�!Œ�L��=�.��U x_+�љUd^
E?��\�;mӀ���;�։W��>��`��ޮ��T��=���ˎ#X0D������~��T-��_1�̞���y7��#TYT��e�[;���,(�+=|���3�t����6GÏ�?pţL�၁w�<�����Ar�ͮ�b��@����� z�O���Y��9�3�t�v��{�wۡYDq�t��|�eĺ��`��P(A���!C�;������m�^�P;<�˓zz9F�s�o���g�t���F������zH��lT϶|���{BvO�tr5�q'��ue.]T枒~4}����v�u1>�s�4�G��om��AD��G	��0����=�yZu�0fN1�gf�%w����m��q�#��?�rR>���c,��mӬ�P�x�e�qD�qux6��-�ɒ�k�Q`_%�� p�CU�h�r���n��^Fu9����0�'�S#����!�q��=�<�}�����j�z���fE�3yhܬ��.�9�чn�'bZغ�u	��U��1�:f�����R\z�5�gv.�*��:�n�ADp~���e���3��m�&}Ӓ��EN��;G�I'xC��w`��<�O_-7�ጩ� )�Iw2���KG�f�/`B7aƔ�3"���Er�F�>�c0vk͔W9��o;��,�_1�Jl�ﻫð���1�U^�l��f�d{z��:}|ԁ*��e'ۿQ�;�@}�I�j�����z:*f"v�\��'���%I�^�7�B+�˯�7`R��[@ؔ� �l����x�<c��h�{z8���^�_����?
��07Q�wV�j�A�Q��g���"��'�E�;c;����,�3��8��=�!�t�z���4[��T_g5Ĭ<��"#�R�1�&�,�K3XQ)1��������u�g0��WZap/I43���<;�@����~�e�+gOԺ\��dJm7�����@>T�k�O�=R2�⊕Idj^��iS�v�|mu�̙���\�5�~&�>W���u:N&�e{B�,f�>�Y��Us����P�-�������7/[�,5���\�;����sĖ{ǵ\������Y�SuX�"ml����Jo9_<�f��٪���r��خھ���IVP�̼͏]�]i	�BN❩w[���
�>�,,����+*,n��]bܣ�	7�lm��0�b�Ѩ�/�����Z�Eý������ks���p��l��`���̮�~軶�Ͻ�O�۔���D�p��@�:����T��t�D`k�3��l���.��o��]��"�9y�d����Umٚ'��#U�;���fܥCT�V��^�v��FL��.8+�]FP4Lf���"O	���뭭=T�/)�\�*�&|��O4;�q��tʚ���xvZ�MǏ�Ǽ��=��+�G)�ީ'��n�S��݇�g������U��g7�!��\��7��r.s�G`�G{h���`�1�
��CBx���=��͍�^ܬ���0���A�~�w�cj7;�t�Դ�'��'x��J��czF� �,Tƃ�Ұ{Zc/k�;�^�g���%�W�΁hb�^� ����7�5�V�v����
zSt�w���}YF��U����^[�Nh����	I<-�CO� r�ϻ_O 5V�����
��&j���nf���Y��%E����n�D�˲��2h�i;�׎��qy�j���|�Y ��u	�tfq��f�$q-��Ǵs'3g�\�fe�څ�a:�H��q��o��[,q˜�(�[�����y�o5=�Ō�K?!�^�עjz���y�[�E�:��m4(fqzzǀvo*��CWH<j H35D�'��{���3�.-r��܂ҸYύ���^��W�Ҭ�k��1ꎡ�ؘ5�J��O�W�G�:]���\9;k��n�gZ���fc�s.��U��>�SN��exv���P�����:�5"��v%��9~�E��hdE �*�H]ꃐ0U$�����^}�v��M4}��Q�6��gu��a;g�f�]ʯ%��.�	v�m���>�q�����<�9��{E� y�!��q�$�B*6Ҭ�L��#u�p��V���Я�9���}f:|+� ml?��}�Мj��J���SR�FQS�҆��%��0�#o��D��תwbr�t���Qm[;e�<"b�$�74�;��M{=�ia�]�#��'y���t���;�ה�<�Lj"f;'�#b-=�Ym��xW�Ŏ�oz.��[�qͫF��w+��蠦�ms(`���e.�q��܋�+�*�TppxM�{�W��3M�Ь_���ǳl�r�%6�c&���wU�7g[$���#������o"�ĬQ�_g���#�෦�y���5����94�z�\L{9�&�lD%R����,ow�%�������84��=ۖ$t�'v}Uz{�����`�S���ˁ\�}�@���#<sA�n�3��w�V�R�긺H�v#:��9���/�ػ�[��4���ĂF�����>��n&�+/F�fr�ݱO��^4;�0����M�Uz��R^s��ֹފ�U08�]�V>�����%˸���:^��PtU��z�}T�.K}}��f솆�*��
�xAf�*�����m���g���c�>d�u��Pl��z͠��m��[~�8iB����O��n3��y<w���W�X�G���*�ɜ��g"���#z}qQُ�Ml9���h�RVt�G#�#�'��Fc�y��M�u�38K����i��"���w�O�J�.�P�+�������-P��Ʌ�b��(@m�7��'��Н�v�o��9�nj/SrT�p��>f�t����J��^�#k�g;�E�9�m3V�Gq�,�z��Iæ:�O�L�A㩡|��3�Ev^��9�k��R,���d6���"�Q��aTW�O��Rey��k;��8����Pdo�����9�ެ��wXx�u�����ٶJ��v��v� ���G��DA�b��|�j�������Y�q΋�kzfsei����ޠ�I,q��c��i��SK:s�1w9;=�gY�n�ַ���E�;�G3]5h��aƹ�!�mM�f�����U�5J"���cUP'�^��}?/}&1p�6���iH#��<E�k�:"�#`�y�8<������ڞ.V����H�PqmW���Nt���՚w{L�W�!�a���Ε��^�܏���}�^H-�%th7��am�����l�~���0q��Н��T.=X1�(�"e��e�i�a7�&oDlF�]��z�
�4�ܚ��I�cy�����Ř�����S[Jm�Li�qp�V�Fި��J$i=#�ߙ�@=��������p�].�q��X�&��N��S��6>������g���c\`Z2��� �[���1�ws��V���i�	r;rӢ	��rA���M�%D!�B�>���'��n�B����R�!�#�3kc���I�+�wYB�/��C%�������p�U�VN���΀�etь�g�_������8O���yQ3±t��Aup��DVWoS���ق���u)l�K7�Cn	��=s���;�)����0�f����EC
ئ���զ�������;:~�����1�VcȱLj5k˧�U·s�]\���7 �{�g����V����9xBw��hi��&r�V�h�:u:+�v#r��q�wbEϠs���(�L"�FT��U�t�,�yw�ù!���N�����z��w\�x�jѶ܌�k!���)�Mq�nR�S�[ot��^5���p��'̅Mh���|�(�#��f
�)_�h^�6��\���Z_}���S�q	�[�վ��C���tu�5{5�i��aG��ު��z��=;�rÒ�YЩ�w���2Xs�!���w�������u)z�#�~�s�t��b\�I�.����!K@�����0wF.��8��2�{F�{4��U.�s<�e`�j�$xn�����W|�9��j_�&H�#�T�q��=w�{�!@��@���Kw^�slqȋ����5��j=Y��we�l�YЃ�sL��H�X]��2ӻ-�����a�jŅf9�Fny��z�������Б�$ʠ$��c陽\3dih-�SjM�M�3'}W[7_����6��t��f�,[O�].���e���-uWv��k��w2�L��wYe���hA���H�=�T�Z`�}���3��r��� ����p��nN	��g�6) �V�k7o$OE�`�����YQ�UeQ6:����+-��ƜEl(�,x�]ݫe�����AQ�3iTaRF�e槪JV���]՝���v�Xq��m��k,�뷆u[O9s�t�뜬�����Z�\+�9�Wc^5rs%������spAfv�f-p䩝�yV��CZ��zE��rq�ڌQ+�n_M���@�}�Z��F�"���.���X���%4��u�R�mJX:.����6�s�S^$�ζ�b��%Y�]���	�Ҭ�r ��;$=�2(yИmk���U2b0M�0��Sr���P1�|yl6z���VX�4��ջQ�3¬0�0�_,��u�Z�̢I��(��$��1a��]�W��������߯l��C&�o'J��Q����4b(���
�v=��߸���B�`Τ�]�}���e*8Q�&I�$!�V�fs�uc���Z+�m;yb�DV���%�X��n�l�8�-Ǹ����zj�wF�a9\�0���P)�.�q���tpz�D�3�����R�C}Dɗ���ZVgM���P�\��s�n�]+𩎊��x�P'Ϟ�1�ޝ/n�9c;|��]6)$X�u��\����:U�VU�	g^����kY%��΃ӎ}�Z���Ѳ��+@2&G�:����q�6V�Ǜbj�5�֔d����~�U���>��/q��Ƚ9j\�4.6O9'"M��XD��wW8J�3�wG^�B��Դ��Y�8�uk	z���)2G\,0��>%��5Go���/ ����d/x$�/0�#6����ܾ�˹Y�Af�&ɕ��Ƹ��*�(0��~�����9��f��8养����~�<V�Z��Jn���N�V���F��{���ð���w]a�.��0�t���5��f@˙%�O���lR͗�u�����p'��b�J��ݬZ��y�/7lft���{um����{Ϲ���y����̯��� T!$�
��-��n�/-��b� H�DBD=}}|v�Ɵ^=q�|qǏ=��v�r�"J��S�<���W9���W�|W�y](�5sr�j.���.�Y���x��8�8��<z=|v���%FD.�U#"��ȩpdV��Tj@}z���׌}x�8㏮<x����۷���;�����櫖櫅�X�ͷ-p�*��S߽�F�m�W�;ﶮU�w\��\�\���ͣh��j���k��ў��wm�yb��Ư���y�w���=v*"�[����+���zW��v�Fל�+�c�.��wj5�nQ\�>wUyY(خnmΖ5_�z�[�j����r�˦��[��Ѣ����xo"挢�j���U;���K�q���{�b����b޻�-���EmA�/+��\U��^�\���o9Hp���������gˬ'9��
�;k@�04����q�ê��z�,q7�Κ�Vr&�
.g($�x�)���Й�����㎢�o����%���|�t1��q9<쓃�[aTz<tI^���A�~	
�G6k/L�뤡`'��*+�*����t�3	������Q�.[Ua��6J>�r��R����֘h�`��7�a?�>��E\��ۋ��Z�o�D���Ï^��D�ђ��C�ȧ���(e��]�|��xa^�Bhܮ��f�y�����S6U%59�ջ�~���^ʵ�.�J���Z�_�k�֏�l��*�$���T�8K��蕓�ڸj��ճ�
�#����O�VDL�C0���������~�%��ݴ���e�������x��29���5��ڎ�{:m�xOm���$Y�s��L�WU��2_�cd]���׹m�ҡ�&��j	Vo�p����r������<��,�ə�niN���lU#wY�8u�V���6�5�I��<6�I��"�䷸�z�v���^�x��O�LA�W5���w����9��\/�������x�â��[��P���5y�)�Wa�;�ʹu���æ�|�f��v��q(�����w�4C��y�\��t�G���g��4�$���wMocj����q���j[M��N�ϯ��d0�b2섶@�J��R�-�����.��&"2��۴�L�n2nwf*����3�jczY�*���uA�������.�]�]�䮬u\�����)G9K�qV�I�3�';���s��}����;H&� d6�l�R1_�]q�D�JĲn_���@W\�ٛ�Z�drN
�H6����s�Ӧp��K���=��<lZq�b��tw�ږ�t;!���@������1p��?�j��b7��xC��wP��@]�Iy4���E���=�Eb2�Q& ��rW�U��VR��Ndd����9ڣ��xW(`�Gs+�[̌Jv^�!m��+Pe�n���]I��ݨ�v
/l�[�qwgNk��Q��[���3�ًB����o�JP&�q�IrFE�$M1��V����]E��N͹BG�Ɠ1Z��,D3�f�X�D�B]��9&M���Tv���v�Y�7�A�a4Pi��,'>d����ˤ�
�UUD�]}�� ����Fl��NLZ�KC<8���^� ���Xٷ�tݰ��xPW90���v�oI؃H�*;]}g��S^��\��æ��[|��D���L���g���U�D�*�u}�W�;�W���cM��(�#��۹ɪ�7U�n4Ť�OC��8��z�Ot^�]��5��%���z��BZ����魬��/��n\�h���G@�ޚ��3=���;3��Yh�z��$x��!��Yî�RA�n����w"j���l��}�>�k���<��� v1we�F<�Z���!F愍������u��vǲ�QSEL��M=�;��}�����o���ӱ5s�׸���wG��Tu	m�l���Y��'����5D���^�=�UY#i��S1v��'b2*:�N��c�+��8ԤF���Iݙ�6���MPS��M&"[��밼�o6�`�Ʒ�����k�[.�E�-"\!��5X�{�w��A�ڦ/8<3����<m3���5�Ǖ��_<8@�,G���3Y�e�/:&�n�f5vP%7��>t����{%�1e�W���U�T��v�%u�����8#s��)\����/��u[��3U4�������\����;6��tx������x���z�ps˺��e��h��r1���4_(��z��-%3�v�i�cC���:���U������rjq���De��{���@�Zm�zv�����pB�6ɸ�Y(��y��<�uS����B�+�}�\y��{z���u����gZ�&Oz�~ ��bj�ۋz����~�������}`wݧ:]���X����1�n���e�h�9ߵ�P_����,������4*��4A�dc�l%"�ظ��NJQy������Qy �<M5���<�z������S���3�����'J��焗wEU>=�˸�vFWw[�����,�h����wvj���9�!*����=a���JCl�S���ô���W�γ\��"��{i�����ybR	�n7�w]���bwһz���UVYbJ���v��h��j�͋nb��໶[�9��uuD�A{�1Ʒ&�H��^�KN��ۢ��T�pC���m*:�9X�uޯ7����y�m��+N����T�_\�oZ���=��_gИ>ζؓ�/t�6��M5Q�CGtx��4q�R���U^8�M*�]ĭ.��q��4�żƨ�<�l6Kjlv T0�q���Oyzߪ'c����<z���(�U���VK^Dln�����<��G�Yǲ�9��a�� �L����^G��U�2+37[Y�D2x���$��`�ᅰ��	F���{��A�{�M>�T;6�Y3�7�smg%(<Q��u��=���I�Z/d�^�aw0������i�^Ӿ�m9���HwL�x���5N*�xS�i�a$���U���t�Y_�}���c�:�V! ��v��V�pc�߳KA7�<�JIח�Ƚ�m���b\נE��AIؒO�Ơ��!���"/�}Rn���V��A7�mt�R�/.��}�����_>͠�]�'���������r��pW{�����\����,ߦ=l���\Q�&^]>�,/9���E���u��QĂW�.��\�o2���0���7���޾n1�uW�c�6��oa�͡O^ڏ�xl2��Z���Hk{.��h��:	[�
M���ԍ/��7�ߏ�fֲ4�D���5W��6�y|�׾� �(ͱ>t�^������o�Y�v�	��Ǯ�:��3^�B��.Igl�E�����H�aWB���d�w-�B����Ԯs��	�t���U�1�쮴������������O-3��.�r�,�r�����0	���_��l����C�����ȝ}�c�Ұ�R���߮���:�J=�7d�_*����>�3��"��n�[�MfUti�ݔ|wgj�x76�
p�;*7�ˬ���_�kmUF��uT�� �S��dr���^�s;a�-�g<�I[um��LF\��L<oZJ)b}Kv}*�KL-�j@���q�{�{��8�V�|[!+ٕ���x��}ܔz��S�������́��F�2��V3z���]"6\�@�J}�� �vQ*v�1�7&��;��S��Ѝ��D�T�K�q�e�v�u��wc�n����TT������ܘ��С�W���@�c���;�փV).u��H�ב�l��8ؕ�L�tW67�T��]��������:]�>��ّ��t��bu��<y�ň��v&�ڧ0�0�D�����h*�ѫ%V�*h�������lc0�da9�Y��i��������#{� hـ��� u���/��X�#l���]�s[\_e5G�8I���h3�i�`]#�?Rga]��-�ۢ�3��]CY�SD1_�����n����#�+�&A��`�Wx;�F��QW*�Y�q�l%�m'�U�w[έo.�3�KVJ��Nr���C���\�S�E8�~�7��D�U�M���AY�]�%�ٷ�.���@�qA]E�j�B���4�W��h�@>t��e� �z�q�R��G2nj! ��ҽ<�r��8a��C�{��ֿ������������o���z�r�!�wA�!L^��LEf�1H����
�AL��/H�Kc_��s�����v�A�}8X3V�o��^j�~��V�wK������%z���F����[{�S#j�b.(��A�J������#�f>k���o �;�j��qu�M|�m�ݷ�8un'��+�_pwAS�e]�v��>�'Y�j��Fp
+d�ҝv��r-�8�V��%���3����K�^��J�iGK���Bݞ�ZHc��K�@�C8�OY���u\(K��j��0����p��mҷZ���_(�e��Ś��ގ�m-������V���5e�o��T��'��e�0:���}���4/��Wq<q�t0x��곛?a��gFX��7���)��>����i������S8�!�����MN�����x��<�vU�7�G(qܤF�R���O�-��3�m���=<�j*#N�tn�{.�d7^�N�<�+�7){%8r��d�skl�k=��V}���UM�C{�n�=�ř��Cu��F���E�x�U;�ie[�6�ͱ�{q}^�`�HA��H$P7��1�q��Q��@S9�&v��;G��W�li���ꗻ�V݇*���5�"�z<��H�`�(� Ƹp��J���{�_���Y:/��Ɋ8N�BG@{��y3T��ڽA/{��\'�����[^r���Ǉ1u;���=O pyp����X�R��T���9hT�Cf(g|�R��*F��:�� � ��x`����C�*]�,7�\b*�Q�i��Q��������BJ�P�b߳'gu74��)�
��)���A���Ia!t����]L�O���P��[�핃^�y�QȔ�{YN��7��y���Q:v\�Y�ۭ�r׮%�<p�����Uw�̱K�6�5����m���&��fJ)4��#Vb_f��5Ю}2úl���1���o5��$کrsT=��̡wwq	�V�s��?K&�8���Z9���3.�6�ƭ��^`�E���F�{����T�>M-���N�f(u��$��[�e�4���q���Z���oGH�v��V�\V1�=��B2Y������N��7��`�=]�\ ǤKq{Q�1�)6�$�$�c:��s`hTZ�<�U��mc�a���{�<zu��2�D,�z��{�'�ɢ"�%w60jdޣ9�>���;��L�ו����(a�Ñs������e��ĜZ/'8�x���wg��F<��A���Y`Y�A�v���K�U�/:ޜ-��2��Ӌ�Ng���'cA*$*�C��X����C��n�9��Z�Yj9�����,���P]Yx���R���.]E�X��S���Ym��g5�����L਒��p���B!I0��(��=u�;���u��ԬƄ��56zF���Æ�Z@/f�16��`�ѐnt\��vK��f�0U�K�����y�����c��ˬ���Ё��v��-�D�k�����u�Љwnk�)۪2�:�3�t�3ʶ�o)Vz�z��f�!)'��=շ~�-��CW3��rfs�b�A$±"D�*���ks�}�������uov�ȭ�(�ۍ|}j軶�[�aO ׵���6}/	bt���em��8=[�p���Q��ún߷��(*�Im5]*�>oC�K���&��-��zι-8މE��8 ��w���OP�W^���.iԊ�~
�|F���Qjޚn����8=^_��n��u$��;����<r�g�KTQ�8XM�E��DcK���{'�4	�*w<g�u�/��IEW�_���W�6�#�,�(�i����X�"���_�nD�z)-�=��U˶K2��GY��9f"r��*�}��y[��v���1��"�(+��E�_�[��F��p^�l�I��v�NFv#�1yX�'/5 ��l9!~7��$�X�'FJ�Ci���Jvlʚ)66+�Oj�ko���|�;3w���wl��H��L3�k
ӂ���M�XŦC=���*i�3D�fO�^!x��2�cU�l4)��O�����/wRN�%:��G��5(_�B�����l���qWػ:��Ɠ��]ق�!�$i��S�W�ٻc�<�'kݐ�3� zXP�ttNٍn*�K��A����ɦ���G!7�Zѹ��M�p�����⸷V��uϷ��m�bTi��n����<��V����L-D봁����t��e�u]�c��صn	�*N�E�EF3��%��@�J��n
\Z�Ks�HP�r�U�]�3�̮��]���"��ʽT�](xmww5��� �:��\�KT��c�D;f���W<$�Q_cHmd��(\��씅Ҁ��ù��[�#�Q�USꓬ�,��#|����XƛB3��wp߫8�r�&@�ʛ�4
�1Y�Zle0I��%����s���K;��3�ݙ���.\�b�U��m����㯬�Qھ��˳�p��};���c�8�;sj�WY�f��\��]Oe!�mkB�U%�xؖ}ηz��W=��1URw%;�+I/�e�QȌ$�`*n�X8��"s L]�!����E6k�JC�e#�Y�$.��K܍�,�[��cv)D��<2B�S۸������C:!�\BR�}�+���5X&���ɵ�D�6��Q5U��tfw!�yԤ�c��ҾSy�؏vC�%d�������=$&#S�78Ky|+3;#�.��P:t��L��6�h;iM
^C��J��'�U��پ�f�E[�v�{��^,��v8Q�֥�M=Y�db��(��^e�JX��?���)C��|�&��::�G�6�7g[���_fr;c���&i�I�{��p��\�d-^P����!2����*�&dj���F�UJǇg,�)���٨�ot��m2rLv��z:t7�v�ZncTrٯV�5`���;���}�3��A.bMެ:`�,H�J �z�hi�-n��]�=	��N�t��������̩�T���pN>YSw�w/5�j�4��/�����3��5���n��1��i�����flX��U��ܣ`v)k�G���=O62J]z�I�����7wC۶���r�Z��k1Z�Y� ���H쏋�%s6��N�byQ��yaەp��)1�2�MZ�"��gCi�G2�ϐ�-⩴5;�[QR&�왬병���F��8������ ���&R��a�"�U\�B;��V�Ղ��6�^$X*�ι7��c5t��u��nf�71 e�\BP����i�J�����\tj�-F���EHT"�i�����i$7>�K�d> �0�Fl7R�$�a�TH�
���`��t	H��L��M/:TjV]�j���j����O�l\��st�GP��$C�Bu����׬}x��q��<x����ݷj\j-@�*�~�5[����Rk�u�������8�>���ǣ��n޷5���\�{�k��*4U#P^]�TjD�$�O�����}x�8�<x��׬v��A�@w6����W�k������c�nW5���y����yԛ�؏+������K�t��G��ƹU���μ���o_:�k�u˦M�;�V.Z5lk��E��w�o9�V���<����WO��u����4�_�ż��ዤW1s�\>/�H��u]�6����y���sE;�ܬb�\ӎ}v���.�D��m��)�c��SC�Y�t�S;f��ົZ`\!�VC�ˮ��j�r���M�jbqܗ�_]I��9pFʍ��fH�.(��1	��t:�1��~s�L��k��or��a��eO��1�S:�(�a�F�.nv��ʾ�I����u�<1��U%�3���W�!_Aa���֯qP?�����jVڌ{���A��DV?z6�t�{������f�+��;�;O0#�Ay���҅��H?�S�k���jb�����x*u%�\�_.sR�_.�j��_	��	�q��BQ���e&�cW,%̒���{�����7;*4�(�qJv�>;?�00G��4�,��`Xۢ��+���`�3�4bMClO^0���m
L�q��QS1�wR��E\e�l�e�wy��M�37ɷ.�A�s�i�|l`�|����B��o�0�U��:74K�;��ФU8�:J��{�����˖�`?��W��*n+=>����H�k��e���(uX|����@�Yu�{t�/I�j���=�,l6�]!N�s�!�V�����:�/lAE����IO(ОW.L�.��,
��2T���d˩�VK�V������S�
��LM��f��
ڭ���)�kCݷ*�)Ã��������=u���u�&�w�(G[�����x�Y;	�xc�͌�*�5N�JT7v2�����^p2Dtg�\�(��>8L�s���Qy	�B��L�ӥ�N���\���A�qڜ*�y��%.ᗜu����v��mi�sS���ĂEcF����qO�1�m�u���s/Fg*j�گ7�;��kӵ�l�)O���r�l6���vh��m?o
H�y�{�5H�>��m�Ċ+�&lw%6q�;4#���U!pl���c��ŵt
�}��0Fi����@���l�ߜ���=��SO�4�ōyQb+�q>����>��.�T�ͭ"���j�ڽێ;;!Hg��(ճܜ��x�[Y;A�7;b8Ü�B�$
W��C�R�=�����F�F�
\�.7�"����B�5�H-c�W��ʸ��E����s��^H��U��[��T�2q]ϙ��-Y��v�� ���;;�EM�o8���F8�1��Mc��l��Ĺ
䙬��/�t��cY�7�z�t��=���B�nv�x��Y�=��z+��~� 7���0���\��Q���$j)�8$��c�Ҽ<8)٧p��=��tg�^v�JE�] "�R��F��B�^�HI<��ƈ�}$�,�1�P���Q�.jkԒڽ#U ��w�6r�X4�Cܫ�P�M�&Z��C�I�Sh#*��
˟ ]�����^j� ����`j���;4�QL"aH��:��(w=\�����C�T�owd��'�փ��3OL�x���d��v6�a�#6l�	h�����l�yH��ǻ��S���r��މ,m�r��́ҕ��h�z�x@�{�\F�������G�_EK��Š?U���/+I����=�{�FA��Q1�=�8���=����/=��V�ύw��ڮgJ�}A���E��h���\��50��g�M��J�9��).��sm?\[�����*�J�{JWx3n9tV�,|��9ic�������HʕIJ��5W�.�=XHaݚ$�T��l˒=���x�d��n��UJ]�b��yR��#�S�Z�`�c���AVc�9��qW��o|�?�x{e���hwU��~�3�q�;��d޳Q���T%
����N3�\nlS똓R�����H�W��[xHC7�,O�K㵸6Z��3%��Ѻ�����F5HKV��-<��`-��ό��ֆ�Ј�T�4��G��n1�A���%q�n.4��F2I��ԛҨ2�v�&�|B)�h��C ��<]���(S�7$L- �,� tQ=�tc�V^���/�nAէ���P��X6ߤ��t�*�W�c��x�&|(�)8�V,���OTc�P�Ǘ���Fרw�(��ɯC�Ϥ��^�å/���*�X.?��A�&/���k���x��=`!�^{xV!Ͷ&����k��Y�-롹��R�I�4��W��@g�OC��R��&�����Jf�����[��m�9z���=Ш�ڹ4�E[p�"[��Ŧ��4�j2e�]��Ao��vh3��8���Ϫ��s6�{����q핊�Y��p3:�ӹǊ���Da$B:TQ'W!?&+љH�G�QdU�_h����͌�h�R�jV�_�w�$G3�׏r��m�k��wXF��"r�Z���.�.����#b�QA/QQb����lQ�^�۫5���1�cj�Q߼�{ɹ�* Sk[3	���N��V��f2��$�s�t�U5l1���&��"�^3���ϙ�	���펟%���8�`�:[]QΜ�Y%i�7��\����>�&���_�)�)gzI�]�����H�ŷ*��n:�΍S�_O�ɼ����*G1��x�(�,���|�Y��<��ڀ��+x�JF�1�;N��3�D�����M{���d�~rN�J�� �uW��]��-�|Щ��gZ&NTZ��Bk�N���WLF��^:2eݙ��'�h�U4:��졫9.iN}GDM���ս��C��J<�q�t\zy��d��e�k�K0Ŵ��]�:a��S�33�Vk��O5�ir��jD	�i�k�2�37��u��m�x��J��y�o�`g.�«�p%���t=�wh��&�\f�d@����Ԯ�xm<��ė*��r,[UǉWa�p��]|eթ��Ws����"�'_&�[J�ᵝ��93V�Vz������wTscB�;���C�P���]��2x�K�H�ܻ͝x'q�\k�����vV�kη���������M�msh��OӜ�m¢l�[�x���8:{�!vWw�t��S�uVlؗXNMM� s1�5�������-Y*Ʃ]�����} x~�'Z�Ǵuz��Q,{�<+�\H�C�����'�8e�C-�5wr	P�մv	�Z;=��T̕s��Y��R:��oq�dd�e��ow�Dt�m��Ǔ/�MWF�[ ��Ե0c=�r��n�E�L� �3�d��job�T@�SΌVf/A�;Uczߦ���uO��4@����A�.T�/J���#�ig`­z� �+�P\��U�37Oڮ�ݞ��g�xY|t74����}��	`է��&R<Q�Z�р<m����VwRcQr���Bˢt�*,]2�[|T�UǬ7lv�����,krSvN]Z޶&��:�o�ޒ]وnw�.6�F�آ�A�'�8pn
gQ�@� ���#�Q)��~�}V�2e�T~U�G����ݩ���BWdEL��n��]�qp��q�M<֥�'�;SZl�f]7J�܈خ���������;��p^\N����$��V����̽�^d߹��r|�R0#T�䠦N�0���޿���?���7žK"3��lli�%u��6Tƨ0��+Fb�#I�q��>�m��F�l�*��/���\�2M�ܥ:�&�fo�7;���Jv��>�8||�+�d;ʂ������z̷�әxw7[#����0�C(�g��O'<��1p;d�����i����W��=S㰉��gk^|hl�\�h��/��z�_�]&Y�up�Ty�L��Ue�����a�3�ar5�������^�.�-�#����_��>��_�K�b�߄�}�I���xDFdw�k��H[3g�lV!�u\��$�d����<���j�m^�3t����<D�Taܫ.պL�kˎ23/�����:}r,J�`����[�+W/�t�L����x�T����m�ؗSM��
#�Y�t/��:��	�}�5�m�
H�vQ��cD<|e۷��ʺ��Ai�Qg�Q��oT�9V�Ԩ��CE��:r]�Q�x���ȷt[[�v����-+�n�p�7��)ֻh����/68	�y��o7�  �Y��wm?�a��ǭ�xا/�+�wv2Jp�a����8������fRҪ;���E�<T\�Ǝ�V�p�N3b��l6��m��.J[gT���V�݄Rdd�iڇ둎��e��!ަ��-����Xj�#1(�3��͊=EO���SyA�ocwE\��ɬ�=��(���G\qdG�+��z���yfߌ���s�!��Ң�X�z���D�K��GK8�l��o�$>�{M��Δ�;<nD�?<������D�ƫEuo6��3
���W���q�����|����1q��*���X�J�g�nsƽ焥�(�L;�х��h����z|Bk�/��N6�h<hN2��#�U��ٝ��`'��F2I�:�ʂ�ʆ�=1�m9[wk�H>;!"����fW%ARAd��p]��;=m��AEn�<�i0W�����9�b������Ch���; ����)F^f�XOE9͜ϖN�M�L�\��p�?p6��fI0
E-�(�b���m8�
�(�)B��Z�U�a�O�י�Ы��(8�n�u�[�����A7F;�s��粳�n,'�~���,q�C��mY��Y���\�^�9��e�cA&"�P1M	!.��
���Z�������1�v��y~�,�(��=wLMI���!D�qә�Y�q����0�4��RSǶ�wC���G؛�y��A�a:Ҍ�oV��H�H��74����z��[C�s���<nnS��]�l/�u0s�P�4���}�V*i�x)�z
��F���#)@���Ю��@���S7�0'��5v���etԽ� ��=V�:���Α:o�y"ι��ޢ.��S�"�Fm�S��k���uI�/t�u©��"��χOE$"��F��D��(�4�5l�U��*����Oa��G������;*7�@�L;��k�.��[I�͠3�^�v	��P��S �y�C^��> 8"nx8=��מ���g��UQ����ԁ����V����@�8k4&��T����h}��[��Z�B���`����W\��+���-8I�Aj�oǨ���p�8���V���sp	V���� w���X=��mY���#y<	�=ݣװn��tU�� `�nr�L��5��{K�'_�m���V',��Hf1���xx��{�׻����Jb1O�:<���=�C�*��S�3l���7$�ks,k��%�|[�Br:=�3��|�sfT�vH���e�T��pX8ѷ1P�z�G+��eR��o1�p�r��z�1�e��]�G4����g�ˬ<�z;٣rWl�������9G�;���܍��9[�r(�R6$Z��t����m�X�bb�qۇ�0t(�w/�{�'u�`��kK=���W*��y�8��|�j-�a��b��-#+��#�|H�^"�Cy;gwR�T�����i!����#���O���l��=�;�4��C�:�%�4m�옓u��g:��`�fA��E��7�*}�=����ƜS��Z�^K��y�����ɹ��|���bf�t%�WA�LX*׵n�4��WڜĞ%��aSz�V��S��W�-�Su3��/A��]�w�*���?+\D�h(h�n���'����������rr�mr��\�y],8�g5�8�IWD�t��6���7Ҥ�c��X��%�:j \� rU�l�$6%
"��\\�1�x��Wd�+d����j�dovA�5b�)���Nz�!Pɑ��9$��	/iw�qۣ��o�hu΃s+%+XW_b裃��D>[t���V��cF�N�oZ��>�^��9J�U�0\�6��X����͜�۽����Jq�Sf�[�<I��e<�w��o`��tl����2^5.�鮻�����kN�ԯ��f��E&fo�P�/#Q��|-u�N��0�+�]%�`���h��ʼ�[��j�m,�F���i%+yWE�Й������(��v{���&���}�t��8C]� ���CN}�t��
�9r���b�x����Iᾬ��,��A}Ƕ:�u�rX���YR��������t��+�� �������C,�uQp0���Aop��{Q&��fW@��f���q���tWT��o��)���z-9��sC�t�������2	��i�`�u&V��N�hN��ln��i1����}�3��L_39��Zm�/Yv�D(k���Cl� ��k�b���+Bע�c^��r�N�+GVf�bfCض��E1b��X*��@���T�A�B�^Q�.���m�r���O2 Ep�YŖ�us82˩f��ŌKc2!�R�J���o�F��*�m�Wf����V��D�ܤ�ʏ�h��E�BT䕡����]�����;��g��A�OQ(���o]��&���<Wl�4s�0�8��C������Yws��cR;{K��∋���}�9i��M��ZwZ44er���;1�LV^Q	mS'Y�2R�A}(X���v�����O,�Y��C�|��>�V���M<$6�n�j�E�5t��y�2F��4�����f4Wi��:;ݰkM��Ф��R�Hu�&�ܚ�"���9�}c[�&�ڡ�i����+dlC1m��ݲw܂~�}�ބu�}�{mg#˖f�(�r��N:��7Vv�u�oX��wu�4�ً�a��l�J��`9QX{�m�ua��JnC����]�gu��:e���-^ut�Z}�Cv���WQ
�U��l�s>�,˻���銅>��Je�V��[ȚMf���y���v:�x�]v��Bm�&�,��3C����{\w����ö2�ފ���)dI��@ܔ	���)aűu+)��赺��t�M�x�6�J�.�j8Y*��hua��`�M�c��e`�&���SVk��G�ܧ����ӱn'u ��g�[�Vql�3, ��>���9r�)��V2�ZiދF��h2�	w�z��8�w�Qy�셗6����u�u;��V���(��D�këp.[{�m��NH�g���� �D�٧�,nUp�wq�'CP�h��(=�v���|�y�	7�r~ԳT�I�5��e��`��Vwl��d��$��e�/#�����q��sn.��]Po]�n[�������
%@��O�x�����8�8��ǏǬv��A�B檒�P����5��s��y���\B��$�=z������8�8��Ǐ^�۷mjY�rBB�Td�W��=�I�\��L��5BO^�z���}x�8�<x��׬v��Z�.��URI H\����r���ncss�.Nuw]׵�߫���Q�X�s��.`J<�]P���s����d5��֧;�?�{����b�¹�(�\�QY1��݌I&�(�\l!F���Ќi,\�����H�R'7Cs����R���_��O�_���ss=~z�*)�h�ſ=�t����F�Nw9��7���L��w���q�s%�W����k��Օ��:R����ۘ����E��H..];�š	�)��%��h6��?���������.˥.l�/E�7�^+�Z]޼����We>j��.��_�3�e��`�9\kW���L��b�ˁ��wW��!�nզ�5�j����k�ElƎ�U=�2�頕q�n������ո��۱ok,�n����a�`7�DvL������3�Ǽ��/y�62	I�d�.��{M�k�O�܏�=E��`:*b3�F���{�f��V�#:B���Uz�����pUY#i��p��i�.St���2^��n���z��-�㭧8x�5AN���c'h6��6��9[��9`��YXeFn����lDr��q�&]��(��e=�jG�C(ޗ��K�1�u��0C޾�#��饆�b�4eW㰉�dpI�c� 6S���5fog�JF�"}���-5ʬǣ�{���"4�g�ؙ�"Rx�� �I"���ړ
����E���1�rU&���;�賫����a��Js�.];[�Kx�M녛[���̛��i^^Dv!����[�9J�B�6��ڵn���yv���ܛt�Ǣ5�Gx7����{��sZeb�Sk������3��ٟv��i�V33^�Z�_����D2��eN��q�aj˫����e����4
��R]�K�hȪ��H��Yiʇ���8.ZQ���ꨗX[xUT�H��5��ñܘ�
����ƒ��4QL���3��Sob���_��N����D�K-����1���p���̒�|���S�ۦ�r)��kr�8�Og����V`������m�.�|�,��9���8�fkyT��T�<�:}n��У��V�ݓ��Q��k�Y�W�i��&���:�����	����6ØR+yB���z/�4�~��iȈ̝�
7�J���f����4����tnC����]0a�;9���U�U�^%����o����qM��"��9ּ@�HL�[1k�?PK5b�]�m.讐��K+�_}��{�貭u�Yw-+I���_sEͅ}{�*��P� ���FIDʴ��.�'Z'`�J�8���4&p�Y]�e�^8�d�/��H�Zu ��3�1��e�trN�Dl�X��[�D�B�i�e�h��FS���W��1�$bꍚ&MsS}��{�q���9��~�!@
Z�
ݞ�ŮٯmL1I�0��w,J69����r^ߤ@W�zNv�w�X��{���U��5���{L�$O������`wP�\�;�{��;p!�;;�U�3i��}R��(J��o��G`J��ԫ�|�X����xX�F��Y��i���&gW�=����V�:�����Q�����9m�
BN�C����aZM&�}ޞ$��+<̴轵&)�l3�;
�[��
>{G�7c�G.�B�{�0�z��QS{�3�u�J˟$m���ԋ�[��TR�^��0�f���tJfC�e9��C�x��:��_GO�+�՛c�۰�.��":�fc ;C<3��O�r:�������ΏW_�<�߁��)w@��M�`j͊Rs'��ԋ̣lzi�?��ɖ��oiTc���M�sQn��ѷ�f����%�ooU,h�I��4i
���Ѯ���ʽ��橸��F��[kX���rm�@����J
>�'�Y]0˩�;�cs*�I�r��_n��4�����(�)��x�*3w{2�\|�k@~��T�oxx^�$DԒU3Xn3�u3 �?m
���{����n�ndۘ���w����qu���vnn���wn����W@5s���{Xo�`9���ߑ�w���.u���F��&{x��������ws$�ϣv�j�3�W�Ή��O���Ѝ����ԹD��O!-U�)g�z9DV��F�-1�h�~)�1^�5�ͺt���~%M{��cD��N��j��ɼ+e��^�5�0�q|��'ʌ��}��vU:.
�˙L���,4@�C37+5�с|��q;�r�9=�欛��N�a�2�6N��ț|+_��r��Ma��h}wo0x�	8:���xnv��!��O��YPyq�_N�{�H,1�%�vCl��v�NB���>8	�ax?]���T�[�c
�O���M��ᨴ2���}Yl�n�:����»�p���+�������\��y,�WHd)�q՛sKKTL��m��z���A�U)Ġ<��W!u9d�vCw�
�����1�/��2�t�v��YW��ed���{�Y�D��M���u����������݃7�ܾ��xaB�QWI]��=�c��e�}np`��3a����<-�&�/@@����g�|�ŁǺ�W�v�g~��,��}���n�[}A��������:��]�u}��8���mT$��ϻ���v�z�z�}��&���M���`۴�J:[�'N���ðo@YY�ǵ�Җ�.[˧��|��^�n�)Jq�b\ ���������ַ_��ڹ/�+@�y8�ofEk"�A�3�:��N�>�>M1�=O�ۻnp%<@��=�����ꬵI6��*�����'û6Hq��aK��}���!Y]°w-�����W;h���]�e�ǖ�`����B�[~��GWh7x��U=�nb3� �Ү�*�d�6z�m0\^���08��.��u�3I�����em�Bm���rw0t�6T���S;{χ�F$�S3�i;�Ha�e�ܫxZt�H*�n�Ԥ�D��̮���NSΓ��S�UKw�7��^�Bf�$�V�g@�z���I���9g��uV��S�k���+�y�o7������U�߅A��jDɕN6|v�}tۧ�+��8���!U�\kbT#��)�8��=���Kl-J����-V�X'�W�Z��+X݉�z�ݝ����Pk�B;�����H^-�9�1{bbZMn�?C��u��Ӣ�xI��V�Kݝ ���P�5�i�5AJ������(�3�2^��D{}��]���]��xwv�VjX�+_y�wx���U�V'v^"�}������(g��8o@z�$�0�{y��qE���Z{ݼnw4u$��l�n�]H��C�v������!���!��Y��p�':|,0���w��)�R{=^F�}S�l%���k�޹&�����C)�`��%�V;���UA��!���@xۑFj��zݢ�T��=`:��oyY�]������t�-A{�iQ'�a�V�u��8~�33Hwrs6�4J2��@D}������#6��������2fbA��͔��n��d�\P�J��t�YXǤo������m�X�Q�Lяc��X�HX%��Ս��VY�ם��	�G�}(�ݹo"�����	�p�x42�h�B��JD�&�LJ4Ix����>?��Pa������ݞ��J�o���	�W�`C;�^г�G���;+�;e����m�2&jJ%��1�=�d#f[[a���(�t�����^�D��T��\��I��u�J���W�n4��c�Y�hU8j{*��-yw&W��N�_k���nʷ��F[:�6�L�k�d�
��I���ʘ�v�du��M��9�����L1�F֑0�]ӍN���'V�>^#�Es��2����n���^�^��w���p��$�=_3�d6@!�s:�3�\%�b�����("���GL��8�d�������Z}W�vp��i��ֲs�Ş�Z��:@{p��Os�=j&��v7����j�F�R�xh�hse���#���ݾ��0�뽾��M�r�:�7z5Iuo��ݛqX1��cO$�;[��.�-��f�s횶��p�o��H��4^�A�:�a����+K)U��0e�te�<�Kq�7>�t!������iY�-$+��޳(�إ�</�N�TKZ�8��_��m��5q�$'�ƕ�M��z�,�0��ѯ��@>>> �y��&����P�12��].p��R�4�yk�^�n��RŹ�[u튭��M2ю.����Uה��uQ����_����Y�gi�OESk1D���f��Pl�ŷ�B�{f	������SFڬ��sjN�������g[��'2|w��V��!<戔a�}�Bm���|<q����5x����⮟�g
���ϡ.��)Ʒ<�X����H��F�)]W�����y���Ӵq�8�~a���{]��x�ی˭207��*;vۮy@�=Mv����Q��{u�2-����]B6^`�';F.|
�L���I�K��Ԗܬ��6�.�ʚ�
g	�n,��`���s�;�@}ԩ�ĩsiZZ��?U�͙�ݿ��R��H�>��O��M@���nR��}�ͮ:`�i�z�H5�,�}�1��/��t�	m�Wt���
@w�[T.dM|WV}�
�{��*���QO�JD��i�[b�	�zs��F[ᄍ���	;��/����v.4�AKv��N�WGn��y�TJ�]9��w@� ����)��w�	��~���i��}m���=�h��")�H=W�=w�#����rܹ?�����_ْA�'Nɰh63G���b�]�9h��[Vɪz��YSݺ��3�z�P�։��c�����=>�LhF��4OX�A�ټ�H݊�/9����@7K���UY"�h <���sM�+A	!&�H��C�N�5?-W����e��Z_v��;d�i`�]�dl./eVgy�.ɖ�}/�X���(a�̷����w\��KV]���0�
�*���������D����TЃ��{���횚�9/�Rj�8#�iNWJ����;w���������v_f'(\�?F>���0I�(c�?���u%�r��� �=���]=T�1��G��*�3j0��l
3�l��W��Xm\�6�H����A���]qKm�T=Nf3�dXm,����������p;�*��S;i|���\sl
M�w��Ъ(ב�n��{�ԧԙ=�2ghf+[Z
Դ������ʥ#l�l� �u���JSZ��	S�x��O�� �ox�.��*]>���=�#������@㵧�Jx��с��.�u���N���^�] �(�fjB9W�(��oL�o������T̾]�xU��lԉ���ëq��N�%�C��dxqv~ك&DB^�*��"���s*��lD�ޝ�w���������L�<������^��h��}�q�L��@��9����ԍx�U�����읈f�$c��Sn�U���nY�6\�ܽZ��a�aj3���#!����s��lg�Y�Uٵ�1�Xc&��]^��{-��lU%n�x�E��Uq,�N�}^�m.����x<.���^-����(��l�ӝ����
��[���N4��P���NRP�����-Cﯝ⢪}Ke��*�\�Uf�?u��*����7
�+�D�Cx@����<�~�������ݵ�ʤ V������ď�� "/ *�)��(�(4��+MH�QL�L�m�Y��L�m��fښ�[5+i�f����śZmf֘�ږ2ژ��5*�R�56��V���ԵMi�Z���55��WkSSU5+SSZ�����MMjmf�55SRښ�lԫMKT�ڦ�ښ�TԵM�֦��jkSRښ�lԵMJ�ԭMKT��Sk-SSj���ԵMM�jU���56٩�MKT��jjV���55������Զ���jV��m6�j�����MKjjkSR�5*�R�5-��j�Y����55���MKjjU���j[SRښ�����Զ���jZ��Zjj����B���B"(W��O��ԭMMjj[SR�5-SSZ�����MKjm1�A��TJ�(�B �i��@���E
���U-KZ�jm���j��R�ժ��ڪZ��R���KR�T�5���"�A�" ݂��Z��R�ժ���T�+j��V�Z�Z��mU-J�RԫUwj�+5j��Z�Z�Z�X��T�5�RԫU-Mj�j[PB(�A��!j�iY,֥��������K�L�f֚�i�V���b��jmi�-i����՚��X�jfٌ֥���ɛk{޵y��e��SU�1��j[l���+Lf֚��c��6Գm]֮jmTԭ��jem2c*�ŕ��2��ɕi�5�1����2��7끿`Q���TAF1Q�QT�O��W_���{���~'>�����o�������o���������������{�����i�����?����
�
�����C�?��@��)�E��`�O��
 
���a����I��Ԟ��������>����~-��0����6[SZkR��֚�ҭ5�����j�֍jf�&�2��[QmS-k2� VEDE��A@ 
%j�KkU��jMTj�Z�KTʴ�jKT��M6����֦��Rښ�ԶkSfڙ�KSj�S(A EH�E����G-SVkSM�Zʴ�KT�kSV�Ԫ��Rږ�kR�Mjl֥[-��j�$ �B"Pݟ�!(~���Y�'���2
*$��2 �H	:~�/����� �>/� ����� �A�P'�f���yE�'�m!���a��;����� ��~(~���a��ZdQ ~� _���A���G�hTE��7�@\O���A�}.�������}xD�q�a�6� Y�~'��~(���P U������}�C�����?�}�Y���� �O������� ���B��� 
�`5���������bQ�(=O�������S��� v��}}?4���{���^�:�dPQ�0(>��lE����[��
C�O��PVI��X�	l����` �������_�����%-%JV��j-�T�I-aUA
��SmIHQ���أ6R���J��d	[d��J�D!Z �SmET���ى�kVՠ)
U6��&�j�KJ�Rض�ֱ�m�fƚ�ڭYm���eF��e5�L�����lh��-lH�N䙕�cM�Z��d՛��յ6kc5����e�ٶ�"���%j�P�e��Cm)��5��#� ٥�F�d�i��V�i�Z�im$���T��TZ���V��Z��M�  .���A[jwk���J�F6�ڸtҭ�7Qd�}���ݵ�Pk!�U��g:���ӗvht��qk���0w]θi�5i]ܩ֚Rn��V�mf��ͬ�B��U��  �p�>���FC݈�3���6�Ҿ"F�YkMST>��=�����ԡC�4*��V������v�m(n���mN��+g���ZuKu���ە�uN���U�g:�t5�+��m��j[[F�j��3YJ6��   .z��ek����{z�4��������[������]�[��k��*���h4ӛSm���k�W��l���hr�iV��ڛt����9��v�-�u��6e����Z�[T�����   [�Z���@�qՁ��[Z�i�����84(ѻ����p:���Cru�@:��-Tu�Q];,�GZ9�4ٴm�UJ����+ml�   �z�A�ա�TSUw5�4�ZM�����ܧMj�������5 �s�C@]�n��3@4�	��ZؘF���[[[l���|  �k�ր���>���n�F�L�:N�����]j�Z�L�:6��
�դ�p��96�۔i�A܎��
���`�U�4�֣UH�lR��  ��;b���nz���A�ѹ*�E)����(U
jn�uQT�{w�)m�S��{޻j���nػގ��J���u�U*M���T�iH[�b�K[fa-jk��M�� .����D��׏UR��7��!AQٷ�����J�=W:�D*��s�zdu�{����J�)޽ozQ��w����:�����WJ{���6��U�KD�-��[C
�� n��JU*FyY��T�ޫ�P�3ާ�RR �<��T���⹯l4�t��f��*�7=5V�4W���=ICm���+޽��`W=�F��Q��I�YeXH7�  gw��E%K��y䝴�UVw��T�+ց��{�U*D]��*Is{w�T�U�yz@�)�R���y�"�P�����)/�"��JU#@24Ѧ�S����   �{FR�   O�JJ�hF�4�j��A6�T��  OT�D�UQ� h3S������������Y2�0��T7V�-S�!M�Nj�4�Pv��_��W�W��}���~�?�յ�m�v�U[k��[Z����[Z��������kUU����m�������k5bB#(�)�4�Ԅ	�=�zXBáO^U� ee[G�F�i�X�`X��Q}���&-Y�Il�7��32���8 �h�P�=�A�ʕ,��m9�3r-�����	�(��ne(�"+ӻX��n�wFn�$�i�N�J��(��K4Qv\[�D���J��3M\p�A�g�6��z�V���7h�:�cE��`����憊�4�H
���р�vYGO
�d:3�\:�����N���l!P�.jL��Q�;�h���:pU�`\���e������FB�H��ojѽx�V�ʓJݫү�k���P65nK
��7.d�r�X
�)\�����K�yJ9�Y�!��Pu|�p��qM�|�;t����7��Z�[W�jXn�B�IB���f��1�4�!��}�V���44�w{��8��smA���!�����,+U��D��ђ}wu����d0�x١����M�:��m���+T;@�	�m]Y�(�k���2�V0FFa�s ׀V���c4�q'��D��@��d�%��Q�O�F��-�:���{��2�Bh�1�P�n ���ґ�ḺX���M�0\"����U��;Y���i�Q�)�Ã�V~1XnA��0�n�w�X��V�Bco�u�Y�K�Ă����r�+3X� X�z ���B"���y�O5��&�.[
����@�E��L�@-��-Swul�U�ޠ�
����sn�X��v�10l�0�wNq ��.Cp��Kf��t�ܼC�Y5ހ�:X��NV!��@�V�f�*]�܆�W�a �o�u�#��<�1#/N6����	q]f���]]x����O�� �ue
�x˽ذ����[XpZb"u:�j&�-��6��Yt2��������
��+-�l]��@�̏tQ-�fL0���X�2@\��@]*�Z� ���fYC7V�K'�{t
ikʁ�Ԏ�mqe�t�a
5䆻=��I�:��X��i��RT3s ݵoVPM	o�{th��iۊ��tr�N5�5����T�t ����3:j-��M�6R��79I�z�vL@�����pSZq8�j(�Q��)Q�S�Yth]�3^��O"��;��WSbYp�ˏ(M7�D�1\,bU��JZ�X�R	�vwZBKr��r��U�Kf̽����.��o`��
xӴ���HJ͹0���,��yyo!Kl޹v$�6T���͆�I��.����"��ʀ��3.!5�J&ha1�D)�7H�z�&Ɓv�gΣ!۴�&��	e������S(�A��OL� Yx�.�����v�P6
�F<�M��O�c����痢��}�b����{��˅TiS��1��>i��R��t�#awSejҨi�t�ޠX�J��G]ۀ��*+1de��v��Ѡ�i �&��j�/U!"Ef�5ب��MYF�8��P5�,R�Y�Cif�t۱�v��V��M���7�ѤХJ��^P�ީ�XU���Ӏ�EK��:�<c@�Em�&�˽	[�.��L�:t�v2�
6�Y��z�$�JS��KP�3&�Ck,(��"Di���ˣm��X"ͬ�nm˦�&Q���Z�"��m޴M��e^4 ��-�Hh�Si��5)�>Ƶ{MY�k2��u&Ҕ Hʓ�UidBX׻kJo2��,;5{*�:2\a��:(�7`�1��q��'�+��K�	7WZ�C��7YX��P'�欲`mD�a�U�ŭ�e�D�{j
�%���]���3K)a�0F�g%Y�ٙm��)`�˘&�4t��i�+aR��%{Z^�����scw�!LB����A�q��YmA��8w3�q��a��Z�l�yoY�ݏr��u`R"�b�9U��ahlߣ���*SM�c��o{��V^J3."������h��+st])�V݊Ϧ�KeЦ2�:��j�h� ���]�ӵ �·n���*��#����Ƞ��V^K����1R2]�ӍF�K~9r���Z;���ur5pem��J�[��ڇ�I�wu5���^VMDޘ,�T�!\(Z�$�0��+��
�U�t�E�r�Hhы%ѣDJ�����ӣf�R�v��DE��YI�ֈ�%�F"B�6�;&���h��R�i�`�A�e�j���в��vYE[�Yp��R �ꢲ�äYo�7)���V1�jw�s2�bR�]5���%ĩ�X��*��^S�Ĭ�	���sMOqS����B�:ͬ��l�
ܺX���A�4
i۬�dWWeJ-f�9�r����]7���
�M����*_':ۼ�T�a[�ʚ)�F�nՇ�XѨf�@�g
�jf��)�U���e�Z�m�E-���*W��=$X{VAb !��8M5n�Gل@�[�q[�jYˠĊ��^�5��gأ�r�iT�Lk']��['@�K�虇�j���fn�Q輫��:sBɧ�5��XN��W*x�V`��-f�e0�;�]�y{����ȳ�f���2�0��C�^V�MZ�m��
�A�#���U��3Y��[����f��E`�(f#AD�#Kq�z�b¨>�]f�
�H�e0�9�)M�:֡�C��旹Z�֓5��B�q�;�x��:�o�l9��_DŊ{�vR�	aU��(�Ŝ�7�܆�i��9�A�+3J$��>o�i���6�ֳ�X�#F�� �fg@Q��Z�0�ƭ�w+ShƲǉ� �f�l3q�u���Җ�7.}�#b�*f�
̘ 'ס@[���[߮b;s��¬��W+rĢ34����g1�����h"�ϳt
����K�)���6���MWJ�i�y�0�Y����P�hCJ�CXץn�6�f�a Hq,&�B��I-2Rj �r
F'���s1�K]���Z�KkM�qR��A�!��Xu�H�J��7��t��w��;�6ӎ9���b�k���h�-d5.�A���LbD� �+6�7kj٤	m�Ʃ�U��#3�20�[�-Fa�sUvV#�M*�� �;N���zo+�|�]��٭m�A��)n]
w�e�<�$�54��2,IL�p��fhX���Y��,�G�������*3Y*���!QS����rZ�ڗ̡��p
�E�1�,/\4HB�6�VfS�K�[�T�L^9z���;+
�m�+u��h,Ia��҇]mCw����1��VdS���%�B��3�ٍ�1l�BS�e���G$�{����"�+Hhýa�[|ƚ;�5���v���mZ���L`�67D]\s(��#5i�-#�)[�cVG�SŻm,h��	�wnE��d�&�6�Gv��,��3,#��Z���Ĵ�H���XM�wc2�
+ً*�%�H<E"�_)�X&��cR�d�VޖT��Z�̺���Ef�(�bX��o v��A!���=�F=fV�<5�T�tk6�R�U-��9R��yD_�ko[ո�$:���lbn����{X���bnե��Yx֔�7/�.^K���ުv�����Y̽�Y��j�T����"/0Z�	b��!c�F2`Ɋ��C"�6��5YJ����S`J�x ùVNM�[[mE�^.�	RI�Ԭ:�-�N��V[��Gt	3c�qm4�Փ��ى�(0��PJ�FǛGAOX��7v���9EC�E]I�7�TpWZu�4�[�X&�aFL�YWx.Kf�����LE�O�#Z0H5QsM��Յ���1��w����[9yh9[��Ma��LsZ)�"��F/a�we��R�U2���!�WSu<Uxh�R����Aû��{gJZ��հ��s&��
�1aCE-�'B5��n�-��^U���`vs7�l�]\sZ�@��[��)v�we���%����H�R��b��GS"�}��w� �XLܠ�u[��|�4�^�'	M�FV�j�����C��aKi'�M.�Z^ٸ1c/�1m�N�aT�4-[xi
�dU�*RX��Mne�Y�{�L��)�ŹhP�l�f<cL�x�h��Y���j�0�Dt�L��e�����iy\�F���4�d�{f�6���*�lֱ]�X��)�S�m+?'g>�gpn��R[(���V}`Rp_ХRJ'~Nm��eQ�+a�^@)�˭b��@���ͼ��˄C2V�P���=M*�Y-5��v�uVF���vd3V��e7hV��o%/���[
�M!�%k�c��&���Pn�0�PQ�!��=�2eY0��	����>zM!��(�*��R�)u(�I<6l�A��n�4Pei��%3��X�Yk  �Cf2m�/5��(~��҇)��54�N^ �e�-�yYtl-�1��.�)���k(	*E����hb�d��Z�f��T���W���Gu(��7XB��vf�a�v��ޗY�ô��ԟK�(��1J�2��t��dc��n0i��S�͉��Gq  ,U��[Go%k��C�#*M���T�1A�d�h�+����ލSob�Sn�l�1�i��)h�����j�hbV��fF\vܻ �bQH��*����u��<���x)=n��%�L����0�Ī+�.�i����^ފ�OVtؠ�̓d�V�I�F�అ)�f�q6��HM�UhR�;V�݉9{��v���2SƓ
���+EQ5���ʰ�m�Hs�=��4oHݪ;l,G�0����Q�t����WeǮ�%�(�Ɲm�o[ڡj�\W�b�u��d��K7f�m��-f�h�	@�\xZo7rS.��V�I1|D�����sWf	%�X����-�_m+��R)���{A�Uj[�ѻҾܭ�@�i�h�h�72��ػ�`^��y��[1�Uj���N\�%^6�Ssfݹ-�G\Fk�)�Xʽ��b�7Ko��)�&X�z�m�J:R/Iij٘"�ř����72�lUo,��[Q&�Y��O�f�f�Q������/ �'g(b&U�:���b"��*��E��D7�D�SŧD=�W�v8;.��0��V�l2��:5���t�3��ʈ�LEn�Un���цm]�F�� %Dִkst��@Q�eᦢ1ݚ��m�)V+2��fDU@��V&�Y�T2I����v�嚺�XPQ{osp,k�ҽ��&*��&T�a��̤L岖f��2�V1��Ц�����&�D�B�BGh�
��/
y�l����qmvFZrhU�X^�y�a��ٺ��4uQ�[�C[���4��q��Pٳ`������0P��4.�R���H���J�J�^�6Z2 ���VQ=�D�ܸ�#	Z@�۲��{���E���C-f�U.��aU"Jf������!�	��S[L۫C1f3x~�Zv�^�x-SsMdn�uB�jrj�*�5������wCdZ4l��t0TC=��Ц�Ӻ9����+YY�{�f����X�lY�"�+2�홢6�T1C�`VͧYB�iLd����ъT�݊�Rմv�壉��w�LGhP�Vձ6w�b��͊PZف݅��@��wSd��Ê��f��2�#�Y��>
(w+m��z�c��
3bl٬��C�L�Q������Ḷ��>z���*��k�3Cw��bV3��1��[�Y�Bw�f�hw{���G-nV]E���q$"e�Y ��{�ݍ����W�0���J]��xo3+h�t��xR�"	����5b�x������Xq���f<2i�+�8"ʷuj�-X3�y2�e�W���48�l�?��.|���YǱ^���6�n#H�;X�q��r�@[{Am[�����Q"�^��^^��K~���[�6�M��@|/�l��lbcif�ZD��	{n�t��y��F^ۚY-�謎�-�&�w.S�jT��bEN�G]^-3F���R��mn����-D\����ॄ��&3t.�e�j� � +XU�eR�XܣS�-iJO^j �\;�ߌ˵�)��h�(����;�=���>B�qV�K���5	0f|+��豄V�v�UEXX�Q�n���@ҹ��k%n++U��hv��d�i_ص�A�����P˨˷6��A��
w�]�a�۔Y������]Ͷ�Q2?���F�{[��5�X�� l�Ym�c�*4v�1�"2�7X�ZbT.��ʸ�Z�7j����h�j�[`�d��J��u.�N50�]d6�W+V�b�Q�P��Jb����(:�bJz��.���V��{��>2��v�[6��+u`B^�d��n�B�A��F4f#��˩e� |ɹD-�(|r�����E�>ۉ�P+
Ty�G�%IV�ۖk];K.�4��S"Mc:�(�Q��kE]$�i��7�.���:���h�X7V�ot�!�,&�'@�7���nV�J��8 ��3ݱf%���]�8̙���:��R$��
Y��^H ���xhYo]4En/!�����0�:���#�A��*ڋE
���]��
��{	�u�!7^i5k-�F�B���H��I�,��Gr�)ذ�VY,���5�(��5�5�����U��b#/v�F#@���[���Ѧ�Rķ	,�Zx�j�[q����u��ٓov�4���P7
��t	E���9Zb.�<���m`
���z�;1Mb�QW���2��"3 V��5�d��5M��wiQ|>�{^�W3I������5YWM��a|�a��\�7����M���QF0�T������a����	��[KfWI:�����>.z2ft跈�N�Hjl<�&!���&�i14��?p�on�]�,�hH�F{gl"�)�<�Ϝ�|��d�8�4w]p�B��>�L>pgj� �W���^̩8<&rSFs吷G�Yu��I[u�3�U�~��A�w�l$@��M9Ɠ�P�n�b����L��ՀM��6��sr��� �y�'n,BK��"=�վ<x� U�A%t��j�X/�!���FE%�����k���(�g,�g��5V��6��w4A��
T�=QB���0�zz*��Xoq��5T��x�$��V�}�77�7:PT��i`��1��W���u�˧	���p�F�W"�6��0M���1���ŮÕ���3�zŸ�C}�"=������%_m��G�N�!6��CQ���6�;��䵛ʟ���p���u|�O[Y��+�)�o��u��+2����V�h�[3��8�YWN� ��F8�^���&؂ۧk%�v�[�6q�\�Z���N�:ω�z�����DZ��0�){�I�U[��۝�R��kB������J��.�oj���>9�cC�T��)�7�d�bm�����碻�ۦ�{���+��\�Ckw��u1+�w<i�yA�x�r|�u�7���i͖Z��bs��c��]2�W%���QU(őP�6j�㏻[Եh:�7z� s�.c�����MNy�8&M���n���*�4w��%n��ިc�9���S��噻u�l���y���޼��Re�=ӆ�2j�e���tr��rtw|X�ـe��Ě��ޜ�I�SOc�VU
Lػ%P�am����-ڱ�:�XbZn���<�]��5�2z�lx��3���Ӯ��'E���H¦ݓ�� f�I /C���XC�`e�&��[U����r���Z؞$�-�v�<�� 6�*#t��Ǹ�h1Y���^̤���U�LI�5���*�b��,����ܥ�t_L�ƍ
2n�O9���U���'Pc`ִ�3�u��Z@g]��+ë́��4l���˓�f+��+�S����S+��KO\7�vgv�Ը��f�R�9;T0�M;�����f�ˮ���2�[tKŇ��+9,�R�2��3''���w�n�dPcf�u�,^�ِ�6�lo>p�ud��Զ0[��1az�d�w���ut��Vm,0�w|�Ұ���f�u.thWR�*�5�����ǵ��}��4��x�#��
�ķ��/7p\��Ғ�9���1�r]�|�ҡ)�+^D;Px@\�=�dͼѷ�#E\]�Ӌ�m�Yb������F^	�oo���e��W7x�
�ŝ)ma�͂LGq��lo篐*	�h�옺��Z26�f������K�_���R凘�2� w{wZ7�!
���M	Rd�g.��x��?�>]��(y���^������S��Z�N'y�P#a�M��P��t�+��4G����[,���m;�mIr��W�G���l+ѵ�X��v�P���
G8�����+�E�@�m�X7bk�Zx�j�Yv�A���C�>���8��z[v�An�wS:�f�b1G����V���P+77n�Xe�V7zX�wZvYM�Y�7�dD8h����L۠+�&�>�nu��`��&�ɫ3���i\f�Sz��+2��.HUm��VJ�n���n�ż�)�ME��ayYmJ�Vd�#��!��<�%�n.zM�RN�G-7u�wܾ4���f�Օo����
�٦�[D�#�
Q.X���dks
Y��i�N��h$m�օ�N�#hl��J���j#*��)��zR$��gaw0�-�����vN3Cq�����([��ʲ��/�8:�7D�T�=n�I��*3nXc�ܡ�g��eN���̘��B�s`��њeN<����o:�T緢��!�������t�h�6FIZ��:�[��xZhл3LZ�ۥ�S8��D�5,v�5�^��.�Ap�W��k3(���ofS�9]��"&�+l�����F�)�+9��]\Cy�7H�L����J�+�
�iӲu��ձ�5���w��s�m"Sv#{���ie�Z���b�'j�ү��aT3���f�Y��2=ֳ7������[ӆ#���W]��2�K�Azy�{�\�^�o�+����k�ya��P���n5ʲ^���8"n�ӥ(.�9�<���Li�6�Ә\��R�:���T��\!�\���wFt�{r�o}�J��:��U��j�롖�`N��[�`�+8�l�}9N�-;��-���w�)�F(0�0^n0��_>j�)��N����)}yjjI���T��0^GZ����q�� ���f�d�R�HU��l=��WZ��`���9 �Q�쮢J	nu�ʚCP���=�[�[�"��8ql�V�C�(�0rھ!���H�#}����͒��.=Bǁ����S���7r-[g�5�������gi�VS	�׀���V]q��f1L5$��TK]�uh��5TqZ8��Cd�<�8Q�'+��� Ui�S8	+�w0�-`�2vF�-"�hޛWO"�	�pM����[����:��œW:Z]�LˬzƱ��Re=m�e!{��3���FR�طCU+Mۦ���9�}*fh�X��3N,�t�Q�p X���=s0	uoKq�ݵ�`²XSM�f���c�R�2mkӍ��@5C9gX�onr��9ذ��-��:���J,zM9w�Jj�;Zj�#���M���S_^e��f`�Z�+;�Ʋ[�Ǟ+��I+=X؏�K+�Q�9Z�N:��^�e���}���F���h�wG�x������,J���:j&B�����S4D"��g��h�W��i�W�;��']���[Y�)�������۱�s���+(����Rȷ�:�Z*M�*ڟ�Ó_:/���Į."��-�)u�76n��bbvF���˛!YN�b#���N~�Gk�m���,޺[�^�W�]=`�p"u�wWf���=S8Ԩ�o*�ǛYɩ��2�,��v7��0�Y�J�92�M[��jѷl�Σ ���U�wO��D�	-�ԅ��I�%s}N�	�[U�[�r���f��v��׉I�D8Ԣl���Z��]O\�h��vyf?�R��]9s��;�e��.I�P'z���`�b�_�{�F|p�Z�Z�/�v�b�vir�J2��#���7V�Tl�TtN�K�37��.�����1�B��n���]��/]��k��eR�s��i�.Y\�t���}��Di�'l�᪲�)s�V�`��n7լ��hҡ@�ݱ�KH�iӳn�t��5{�C��	M�����߮]�m\�I�8�lM���A�z��e�{;���;�:n�u����#���4�i�.��َ�&�r�����,���S�R�$��UM���1m,'w�w0q��U�ԉL�����r�W�2jǓ���6���)r��! O���>�ݗS��b�E,�I�R�c�4�h�İt{��
C�Z�oqG�)0HNۣX���l]�E}�fS���g�T��t�����_AWn��e�ݳ�e��f�����=���;xq�\���Gv��Gv�t���8g ������n,��aW\ˌ5�S�q '�dh������m��֖���l�R�GT���6�������Ba�����"s6�8:q�;\생v05���׸���]
�n;�pe!|�rM�
�9 �1e.W��B�K��;G2���{��wMP�}�1���;
h b��-�ْ]�.��6���r�ǬL��!!�V�=�= 6evZ�8Ցm�Y���YEU��'�����;��8�kr��u9y4n]�pr�R0Э�l�K*����X>0�5A�n�J���sz&�e�ʈL;�F�kFp���B���bS�I�����-��C\�r�Z���r�-,%��l�aIt�`��w���{[�?��[����~���iC�sĥkܙ�\�=R
c>��=�'Ï-�goQ�(�c��kb��S+8�n�Y����y�f�"�]�2�U���U�W����5.��oH��Wwq�*c\�����.�`p��ˌX�E �3{����'�h��%)�	ϝ�]�!g��-��a��P��
�P�&12ɝ�&�o-#%���;�N|2�7�˷.�p|k�ume-��P��(�̢.��]�>��7��:MT��ާi�arr�V�H}�cL����6@H���3 ��R֊|"���ϰ�:�����GW^�:Z|�&�U�e �&�Y����3]$�vEmZ]4h&�|ɳ/sT<�Uy4hr��ZvCi:��mLɪ��%MKpJq���ΜZ7S�I�`���f��{�ط�I�B��8*���M�P�7y�k$o�-��TO�D�J�/4��#n�Q�9etbx���Ri��9b>��1�g�k}x�/y��0�(QTźB��v�&v�������p��O�q�d���w�2�JoVJ��%6�Ś�DNP�n
�Ϧ��K��+�2�fQ<�@���/CJ+��Y�Y2�!��䇹�O���,K2`(���{	bb�mC0ھ�$�y�s�Ό����g84#��)&�eu<���;�[�������07��=���9F�Ҥ
�ͥ����d���7"r}�>��9��3]8��Fk�0>�7t�g5���L���*ejO��x�n���P��E�I��eѭ��y�d'Sgf5��=,��Ff�sBn9��W�d�T���:����|�`Ұ�v�9�d�0
d�q炶��k\o2�����S�!���(�n�T�at��j�R��s�š���L*��wR�N���ݤ�\9N�3�9F���Ċ��ޮ�6�vr֢Z�F�I8�WwR��ҏ}�!�WCep�oo3���G"��� �B�p�ܫ�k'�X���5�.L�3�VV�4��$H7T�?q�&Q�,��y���U�����	�l���LŻ ��C��uɥ�Lh�.�71LK ���P��j��4����tX��؋��0�w���\�ԑY)�G��ćJB��Q�o�R:XN�/gk��a���P��yZ��I���R�V�s�6�R�K��������+�d�J�V��%&��4���A���Ԯ֫V�=��+���9�W&���X�][�+dݫDg�A;wiT��u�Ec��RU�G��\�T��%K�h�;qX�2'OGS1��l�t4Ḣ�1L�mr��[�;�L�A�+�:mF�М��2L��v���E���OgQ�f2�e��r�B�Vf�S�����?��^�����f��+�\�]}���I�r�l%��g�n����Z�Du����tD[5�f�H��mr�=W���*s���:7v6%���p��H��3�̾Ď�еk����_Qj�P8��i�ڲ�n��v�	�VCn�S�<�V�t�)�f�6;��"mɚ.u�Չtx�LoA�0���BI=n�p��ܜ�Q�*GKx0��!yRGz�]^m�Qd]���	e�t��8Uw]=����![��fP���.��t�է��a9/��emwX[�*w���筤�G&k���ĳ94'�j�]\c����w�'H�G�n��/�J*t0�����Ħ��&y�WZ�U��V�Ե[uj�f]]aI�SohX����c�w�H�&�=����A\�f7��^�����gf�"�h�)Bd�F�M7r��5����.]۝.���z[9�a��G\��k:��^,�
Ffu��j4l�uN�ٔOL��r���=cM��k7&}k6T����p���ĥ�[�^ͫE��|h�}����k�p ����u����^i%��}.܊m#�-�c����wgD��۶2�5H��[��v�>�D�]I]�0:�#��j��ڭbZ�sR����2mh�쭬i��ɪ83+B�*��Ӑ�7 v�
�WhN��� @R����wqPS�+�;��u��SK*V���/��;q;#pi����A�G�2�K��չ�kK�+�VCN���Z�6#Ȧ-�SGǶ������z��
Mo��]��n�/���N��LS,L7�]e=�A��$�LS�
�#d�m3��y���c���mLn��6L��T�6�!C��*���gk�Y���)L��R�G�h٣�I`��uYj	#lؘBYY���vLD��̻�#%^��h>I�ۏ��8���5�,�y��nХ0+X�_�p�Z�����Pٝ �-&a��A��k̦��N�%���i�K����+^� 3_�Q������7�Vq�xǶmy8
�oZ�b7*18nseu�e�(`�Y$oW���Yu�� ���-֏V���3"ߥ�R���h	Ry�g#k�!��*F��n��><�XJ=X�B<Ao� �k;�ĵj˓�-���.��Ӿ��jŸ��x���u��Y[%=ā�/��(�fa�����<Y���[�[n6o���)�9����Z���&������g�����g�I�H:��Ky�dЉ�y�����)<V�����a��Q��t�6kt�Z�#p�2S��غ�G��s�Zj�V��F��m��ox�SD}/��WP]�o�}:b�ð�O�����L��"aҧ:6��)��{I��CX �o-f�w-g9ք���A�"��U��0I�Vi✫��D�yr.�Ƅ��!m=޻�zw#3KΜU,��o4��i���N2k�q��ңk���YR]"W@Dj���wV�]OMo��Q��
�.�]��{�]�"%V���d��b՗���	�����Z��m�*R�w��u�c�e�]�jN�� 3{b�`'X)� �Z�vv�����='P�-I�����  >�������������������;�Cz�a��櫫F<]�o�+or�?Xہ���i��h5�^#	dAk{��F����h+T2���Xn��2!�U^e$\�6�b'�;��qv-��jA���E�
�/�D;xzj����j��V��i�%�I��5�v�zz�����]�qQn�xz+"�1"n�X�X5ҭ��\%��gC�w�9Ve45w5� r�C4n�;���#��.��sB��ӭ%�WR���j�B��P$�V�r�Q����M���sV֛	ERmu�EW0������)�A�ݴh�;:�A-���rޗ]6�J��{V.��pu�z#S�v�)Q77WUѾ��F��r"�ۆ��@+������ݰ�����ArZ�p�c:�S�=yP$.�r"Zӆ��C��������e^�4k��2ma���rshk�0�^���"1��ᇇe[)-q�I�
;�����M!��œY���>�ՀG��3M����-���1	tz���4@)�ë/b�&�v$���9/�\j���}�����˩v�rp��Gw�*Ѧ�Vh�wj��h�M[6:h�d�FmLu�sZ�ս�$]q)D����9����w�Q9r��灈�=j��;�ɠZ����{�`�+@�fV��y��� h���Y@�j*�R�d���f]�ы:T.JU2�c]�]]�K����?��ipY/rѕ���.�V��A��s����:�q�	ökEq��ٙ�D�qHg<ۺ2�kI�����D�(]�F�����p�R���_]�[wB�¯d�����u���,4�u#�9��}�-�fܘ��v6��e&/1�t�mŪ�D��k��P�MΩychۤ�%��}[�Q��X�.�r%FKӻ��ҥ���g;��=�D�J�S��ݒ����
�a	Bm�YH��|��%���"m^��<F����9t��G5;�ДS�Q�O�&g�cV��@�-`�L�	X�2MU�ּ�V�E������l�]��i�.��W˰B�>�5��q]�V[�V2]N�aV��\�ڲ�cl��6�
\�+!K����Sls5�e_Qي_vR�uzI$N�#��R�8tf،�w�a�a)���tN�=�)�ט��GT��λ'U�'X�W��p�^�$ =\P[]]W1�d؃�a�9O^Yp��Ԟu�MM�B��a�v�;���E8ܧ��),n���֫���inuNɱI�-�4��S��P�Gu�R�ZVG��坓k��ֵt�C��[����VTSR�1P�B����C+��0e�yM̑Z�=\�$뽢�\��s�-���gd%@��Y;�#gr:<�#ǜ�읗\�;��}ЛŴ�GB�k&'������a]��TUj�����rjv���l&me����9�GR�O	N]�Ш]v4$�#5����,��%L� ;0��vؔ򣠫5}Hv�A��3볘��h�9R�����t�
��Ao�C�m6[��lИ.g������C;Ua���d�nk�3�;�v� f�Y%��ub��3�iqչ\�M<�h�,'��X�I5ٻI){1j0\7N��l�g����I��'I2m;�%d�\,.=:���&�\덨��c�VØs$�Q ��ݕB��3t�8կY�wƈJ�=�/8Z�F�Q�Bu��Mt���S���# ��{�+��n�F>�Y����a��=G4�8{���#��2%W��v�í�ō�åkKgE`�(ҩ�2��_d�/L�yoR<3���
O�}1ٵ�=ٸ���:=U�!�dN�R�Z��&^I�mKK�=�of�08�P�k.JJulV�
�e�hY��Nh���э�K,u>+-l�)��4�p�e��	��P�P�� �y}J���b��t�F���;�l��:b����-7dd�&�cu�j1��)n�޷�A5]��PV:��«nw@F�3I7-mO�䄬=�h�:���6�I�ӷ܉�+X����R��[Γ,��Ԧ�LY�X�ĭ��`�6���,f\є˔7�؊z/M��7�<�1�^���O]i��fHs�v�+��Æ��p��1pl��'��qw\s�ޚ%T8b5�ib�N�Rȭ�'�f��S=3(�cV�#�%ci,�\��'Q�� ��N��v�p���BJ5}�We]50T�$���tL��i�ŗ��]rV���Q^G$R9ګ��ЧY�F�ͶQ�Gz�pbl�WO~�wQ3�Z~�s�v��ݪf��̀�|�k�Er�����j�/KE��3�ˡ��]U����ɉ��Ѹ�k� �ꔓPr&�Ȓ������2����t�JJGe"��2@&ۺ��r!`�0�n��l����[�:�T��Vێ��W�Y��D�#ͭ�v�s�V]�{S���aM)���r���,6/j�/^M���t���.lb�r����nU}�UԖ�'mK�O��,#Nk/.偽jf��J`ݺ�m���.���(�� ��P|��и���W am���f�\4�+Gh�s�.��	ه�ZU��F�z���Ρ�N�B��An�^�mG���Io{`�-{r崱ع��V�T�z!-Tᯩ��2Z�9Arr���,��n�B��53���W�,�������xEo�L�(�f�	][Sp<�טe��י$0�d��fpy	�?���c�nM�s����������:2��	}�p�F`����������TJ�+<��V�k��������a�}������lUt2�h�/�bH�t���*{����;�t&>ep�Τ_hoC�E������;��	�]�[{X���=��I��j41�8����GJ�i��7XL�R#�ӄY���p�w���Q�
��v���+8]�ެ����X��D`��v�0��qSL���zw�����5�'g};R�!֞e+L�ہ<��;��= �裶冰�'gF�Gwɕ��vC���2�ɦ+�]r�^������-˱�A������I�{��l���5Û'���}�ɍ����k����UF:�Ծ�eLWw�����U�ˑԛyʅYw2��u��2fܻ@w������4Nˇ�����6\m���iI�h�:��=A�+�sn���s}����Jڽ��u�F�#��{k-��*sx��;�	N�YoC��kxۜVآo��ͺԖX�;�$�n�Έ�`�M�a|C�tz`�u�hdB�P�2�W�#b����z7�";��$6���_Mm
�}r�� Hi4�����Gp\��S,(�4LM�ݜ^ja1��	�6��r�l{i�[�� ���v�;J8����(���¬���eV٣�2�!��YCOA��5�����L�ln�)nky;9@����j�7v�K��۬��8�V�yj3���C[̛N��/mH;x�n�$+��T����N�	Ղ���s�k�蒱�I��ݖ�q�
�*����q�Ut������Q�v�f /�VP��\±�*r�7���k��á�u5�SZ*@���'"7ɰ�r,�H�wNn��mHs7���1�쫝l�e�H�0LT�l%y��y7���i�n��S�ܶ�F.*62��M��4hP*��/�d�#���̠�n8�[�F]L��{��1��T�*Y�M��c�Q�*0�w��������s_ ���E�9����Ħy��t�µ�4�R�{ǅƂ��G+��@��e!��'ZkZOhG4N',��Ĭ܏�'~s�
6Q�!ʶ��K�  ��j8�����]�?�b��MȖ٨/[��k?^�i�h3g�c�V���tYD�ƈ�yZ�)rʘūL���`��/B2�v��Yuw:�Z|�'I���+s��ݐ��	� Zع����{3�LÍ�>�[5���_5�^���L�؉����w2�N��XƝ���䠐«U�::i>���6AtGo;`��Vڕ�!�'F��� ������;[ܫ�\� �`)c��}�_WJVM#eoZ�f��
`�%f�]�J�c�YU��v�g�g죃 Ɏe�Z�TZ��N�|EM�ΐ[%���D7|P�w�+��i�o$`��yN�l��k�l�.v��Hmئ�t+9l����r�x�^mo_(�G�Y׬�-ӑ�t�����ݚ'���#��M,#��f��;V)
6��XJ\���m����Xlm����,�r�ɠ��D�;��	(,ז�J����bu% 7����kH�3q�j�H�'k�.�Zf����>52�,��3�����9�&�\XX`Ɖ�G��FW[�Z5�O�o$
�J�[j� [3PP�{&W+�������%�n��N���St�4��Ɋ:e|jt6�G5�|;����n ˫qZ:b�
q�U��ss�.��G`ǯt��G�Y%�cC�u�kcf5x�t�����&�AvY�ݨ
�ѱ��+�Uv7fC��7W�xj?u$<�v��1pm]�����.�:��wY朧C�i.l��$�M���U�\n�K7��Q�0v���w��O���Rm��#ۺ
��1�q�h�.�!��H��!�96�7f�5��v�ũh��*��w��]�AV��(&�km�/5me lQ�+��_Der	R$�yF�֩��-�dXiޞ�o���)���eAB�);A�S"l]���++�5*B�H<5�� k�t��[tL���N��aa����A��_H�dg��{uV�k�!\���L��ܬ��M9�0�\�\S��/^��oZm�]�Q�!p�y-��� j�I�'�oJ��b�a��V���4���(��Z�l�#�v��+[#�k1��3F�^��e�����.]*�4m{O�pU��7,�z�)+g 2G��D=Jkbw�`�hu�:�ˣI���﫳�q5n�*J�d�o쫬��
W�_b����ڟZ�ޑ#�iݾ�f)�v�N�kx�DVˤ�R��l`v. �����'���U�7��h�'e 0�ʙ��e ���+L�u������@8�8�6V]�!y��X����w�ݘ7�Hhq�ݶ��Գ+q��,���}�e���0Zx�
��[��(�jP�S��H��4�3)���ǰf�R�,6�ꧢ��n�	���@�#T�����t廱�S��)���%���)����I,�|x�{�j�E
�;�$�>ݖU�r�,��z�sp+�yٍ��L�Em�N���o!.=��9'2_=��͒�h����}�N�1�ńyᛯ�IC1"+�/5�f4̨�i�U��E��I7�L{9^��
��;Q�U�r�W\���X)l:�KVi�0���d�1��&ġ�.bǛ��K�ҲӑX���4��f�|D�m���3���;ׇ�'4yK�GG�����Ip=pG2[��a������;
��Z�/�!GN>rvL�ڜ�\��W�=���x�bR�ّŏ����-nv���[} �-<.D9��d��h�Щ��^�$��kH}���۲e�aʚ�l��iWm,��]v-�Ы��Ѳ�cr��Cy��勊��	tR��l��0b����B=�fB�ƖK]%*G8ެʡ�KXͧ�(p��	�Oz�]��:%�cZ�]�}
���Q��Jn����b�{2@2s����^-�����F;ȖY��F�|�grȫ�*����Q�9��PY0�sS���&n
k+Ew�ot��K�r��ҴVKɢ�=�$������X:w*����C�K.��&'j�E\�b,vi[
���u%i�=�J�`�D$��Ý5�6l=�W5{��K^�n�'H�va�$��.�"ud�B1�n���MǤ+�e�Yt!|.�բ�5��ݴ��{��IJփe�i�X��h��3'>���%�J�1��ԉֺAt1��*[��z��3�u�P�4��i�"�m������C�F��7S�u^]��;i_6�i��8t�Xܨ��Q�i
�:�-S��N�l����G.��\pVem�h4U-����Z�f�-ࡽ�R��[+e���A+4����ӄcʊ��__h�(!�S�@��J��"f����`��
T��:�(
ݮ��yhY��6Bͳ�Ѣ�뷊Y�q+�VP,T�ݐmL�� �w.��{��a��k.������!��-ge�è���
�Y�5 mɡ_ő[O^�*ڮ�wBV^])�����Ø��.�\�pw���X�on�&X�j���X�7E��eZ���j���\�ykPu��T���Z�e%��]�k9=��R�b	PZ�t�<I���r�9J�{������T(���q��bQ�X�],���u�wɰgL��h���Gͨ�mqa��@��C���}G+���e!j�C)Gg+{���jێ��s�<i��W7j9�!�9�P�˭�֒�u��s��Zt�D�dv�틉�
��L#0�6�ݒv�o8��p�0�K�jdB�����f7�7#��q�v�[B��:j����F��K�l�r��`�%p�d'˻_PR:��3�3X/vm����K��y��;\c�"��\�%j�����sם���
�;�^<�lu�>�}I��6ɖF"��u] ,i5�,�r����5Ό��<)��M@)&�ժ8>�+�9��%h��S�v�;�
�^�A8�.��ŧ���Q�kuF�X�q�}�dCT�km��j���M`�h�3v�yv2��o��uڰ���*z�|0p�3X�Q�
V��jy�p���xI����叇�Z�����`=�Ӎ�f�>�Pb�u�.$�V���jH-��J*1��v�v�C/n$�X�ww��b�p���+=�L��q���6�%�XV����SJ¹� *.ݷ@m�!借,��w3%F&�3m�5��Q<'kA��������������>�K�X�-���qUv"�ѵk{�n��˫��s����LsBЫ%^�ː�'��ɭ���e����/l�&*'ٯz���U1�w>w�Z��l>�[�a�x+3�CmM$��E��Rwa}\t�Iճi�y���ۓ�5]7JT��ä�{f��tN�M���)��-Ӛ>�n���{	&t�V}�+j�6��W�V���魁I`�*����n�/6qS��.�ҟ6(p����:���S���\0Cնbd�d�5�D�1�d���3�
z��%�md+oUn�fh�X�(�	H�Y�/J#�%�Is�J�dpl�-j�^ΝNfGt��dl�˖2�]�.}{'�+���ؾ��At�U��IT��\rܷ1=7���e�)׎�+G%�e���_m֛�D���;�,Ӥ�R����̧eW�qfL�wdw�ii��w*n n�#���W$)�Di٫�â��e�UV�:��j@�����N�M$���)r5���\�*�k���(�z�j�d0�-l]�Y+z�)aZ�v��=6��UwL1Wk���'Jz�]º�6֠��g���"ͳ���N�i�{N��rM��t�����T�#2�U�UN洞�y�'!2���6m�m��]�t��7:P�8s=Yܤ�LD��C��ъ�<Z%�w̦6R�&�n�(A	��|$s+hͻ+�r������ݎK�����]�e(s�7s�K"K��eB�̒s�$wt��˚�ɺsK���r1�n1ntXK$�! "��$��	�"\�L�
Y�w\JfBCِ����@�.��H���u�f��M�lɤ�d�H��0I�E$a`�Ѥ��a���)�3	hM�C j�;�(�2dёw\4��Cb����4�L�L�$A5 f��C�]�N또�@#F1@�f�P���M2̃Ȍ�+�����D
>�h��m����P��o7�t���GE�
N�x3�ζr��d��F��Q�k/M�Λ;[�Z��Qٙz�"}{��VIݹ}b�����,�g>6l�Bj�r��1:�\)}�2����������YZZWI�؃Z�Fhe��C��#7�~�GU�[�m����3ZTkw}찭Ɂ����0oI�N �ߛ�k��7pa��,��2~E����'�y.T|N^W%���V_��_ɘXc�8����`�]�X��	��6���eNo���&�eM����*p����b�1UV�s��sL���kO�W3g>N`�ל��E>��Z�+9��'`�!2�E\�ҁXد�����c;��}�o��wܭZv9սf���g�������Á�� =1߀o2��ssT���|J�|��,�o191<����I��eZ�O�2Es��^���/	��X|��3ˈ��n9�0>���N�3�cymp\�Q�����	`eP��촄R>�gz`�Rk1�kr2IF_�ݽ9�9�9��kj���3���l��n��'@�<�C����ҷ�a\q�iJa��-�t�9�!J����9NI��/]�j ;b�;3c�Z�[f���c�.��l��g*�����T�e��P�&a����L������F7Y15;�z"�t�讕� aҳ@}�����jf��k%�������gWƪ��S1��)��Х0_���Ga�:z����:�!��r��P@�д�TwEבo�{�m��P ,��t ���[3��}����&ɞ~�P�\��r���ۚ����}-��Q�a��aQj����A��� !P�V����D30����Ϻ
[o��o�s� ;�}/^���8\4�@���(t;����df벻��M�#�h�y*=������*�U��� E�uL�U��,]�k��x^��.�S<���o`��uOj���)E���TĆܦL����!��(��c�ua�N�"�,O˔��[[¬bn�>�n[��b��)�K�P����$���3�'��p�;���u�@��&�5W:���kT��A��c� D�	�a��<q�؍,`�4���� E��n�󼪳�ŃhT�z�.|uX�������1�����?����m��C��H��Y�LQ��mD$tU�]S�y���ޭ���d���ϊ�����j�:�{��Ҩ 5S}3�z���CWȖ�٣�F�˚1.;9>�5�1�8��Cκ�`�:Ig��C	�z.�y��RXj��TC��ݥY�<sv�����	�S�4�`����V��rz��%���[9�t�t�0�RB�����xhp����b�\�8�>]�5y&�­^�Aخ�Pq���K�������ק��4���R-GF��fV����3U�/��IT坞�7��3�Rg&H��Rdg���6�)��n�}9GEY:`��3�I/�1YЈ�n	|:z�|)8@A�7��,�.!�l����1�i9B%����,�	{g+���6��	�M�m��L�1uR��E��
��c����smT=Fs���f�]gSx`)�#�3{���vI~* ���4���Β�;�,`��ы�{%������ʜcX]/�nTM{c�k^5�{h���#���K�}�Kj�W.
�|t=��C��w�ʹ0i�k=ƈ�ςu<��  �h*T�zt<交@���X~Az_5�λ�*�N�!�Q��[n�u����'�D�S�@��0U�<φ�ָ�n�=����ip�gQA�o���9��Ys����`�c4.]TQ�$.��c/�c�Wfӫȵ�y�#D�Fa���̆�
�Rb�I;,�s�	��n�*9�:1Ԫ�.K�S��y�Ս!к|�`�V��eĶr�ɽɔ:��	�D�z��u�A#�)<�B�������㓯z�h�Y��#�n]�}]c�w����{��4�,,텉w)On�5I�w��]�IF����ću�W���q8�.��J먛�q,��>�P2�:[�0\J����=��b�%wB�&C�����v�7&'S�S�b@2��}�Q�-Wu��~uJ,�t���eق���WY<Ǌ\9�0�pp�wy�$�:jZsB+��T��� �������վ`���ҵs��Qg�̣�;�T�[$��Y}<�˩�K���@�u�]��\o;Bb��D!L���5�u����:��-z��[���}F��>m�<���"c-���ӈ���ؖڤ�1���ˑ�ʆ��hܿTW��0��a�a׾g�*�p}qz��N�+b��f�����:'��#�_E���9���'���E�h��W��U[V"�T�{��U���b3�r��s��3�6 ʽ�a�H^�)1�0�C�4D~�Es��**J�:�����+�z����K��&��A=�o:;$W�E��ag��,�<I�~��>52�7�Ká`���{��@�=�qn@*H��9�0,Y�z臦�{ԇd���i�f�@���P���!@�7�
��Ev��b?�)���p��+q�X�Z��v�<�E��u�m� ��E��E� ǃ;�f���ϠH�U�xR�%�����U�YD?����.�����`��ݒe	ۂ�[��p�qGfVq�����m�}S�]�\ڰhG0�4����:��d�zdJM�3�%̰��s.8�H��x�F[�p����JL�$�:�=�����њ�T���4!��f{hy��f2	�/N|�ƈ�x�']U3AḶ� �� b����w]-&�Ԅ��o�h\R�C,:�:t|�v��E��Kn��sn�>��ݡ��y���р_u$�=�@Q�99�[Z�z�LC�g��q/�9�;�3����˹j��{5{ ���|���}�8��MNzͳ^�T��pO���/}�Ţdeh���Q6O8�<���l�05�9<��;6�][����ޘ�2�W��wi5YO�pn	����9��@983~n�e������X8I�C��}۞�j�ɍZ�7�|��y] @��L�׷���;��r5�1+6�D�s%�� ��0�@�;�]�MhQ��6�#�~0�7���S�vTx>���s9��s��.�L��r��m������.����
�x7i�~�����|���y ��gy��x��I���.�.f�D%�"?�������d2�^T�a�Y���[[=�ѫD��xc|hw,%*f�ѱ�-������Iv��]�L.-)v�d=��S���I�ԗ�B�V��k��R��{+��_1�a�n� �{kU�k�z�M�Im��M.ۣY9�>�ݻ/ղu��5���,�Ώ�������J�B�]�&��'3ĝ��:2d����1�q���1���<I�Q%#Pg��!��@�l�6n�s���+u���2�f�l�ƻn��czm�*�5�`$�I����e� ��Z��}Ze�U����DՌ����g+zs�rzs��m\1p�q�lJ+�/��$��i��xq~�p����(��T�kR��(1c�:�-�:z�9�쨄��a���ͭ�����^���|W �� #�ӓ�u�`b}����.�M�+��Jm�CI��l�Ny��4K_^�8}�Cф�d`2k��S_m�$� ���f�v���OZ�䁩"��}�tzW.��Aq4��{f���'y��(�6�	�<��eEO�^[�}���1Ĭ�@��C\#�'v��U��,�����*K�Z��!����N�
�i���>���L�=��3X`Ls��r�a�9eiWU�<���2�����8���P��;ŻםZJ��(j:��%>�ۛB��j�ͳA�Ӫ���ޕ �W���m:q[�p�<qsӴ�X�U���6��O��Y�P�iۗ���^�3��M��qPJ�Lja�h�_X�r6Y���g�/;�w��{�������9���po����Q�q�Q�z�"��Ԥ�D��s�1�T�8%�f7JG(�C�^�tjtna����i�ə��8Ԏou����f?@������']P��0szگq0x��u{n��*E�򥑊�-y�5�,��#R�Y�Ok�{���{f	��A��p�+��C0����M�B*01�T�RV6rIQ�2��r���k�;��	��Y�����~oJ^����c"�����gj�����U|��L�m����md��'r���ŉ�g9��N�����d����QU@�e��岲)����1�j�"Y�� �]6Vz]�bM~��A=��`��p]T�S�jhB�.���ä3!�v�W�Mj?o��Yw:�
6%ٺ���]*k�����X3�M*���w��4H�R�pZ0�84�Yy=��0s.c�s�Ȑ`��<ySD�^9C꜊�����uG�B��-���Ғ�y��*9��� ��\��0��73����ZZ���aÉݘ�1��ត1���&?�iN
�!ڜ��U�K��]��W���Tѭ���J�+H�\E��wx���^�n����r���&\��[��Owq=ƦwW[2�ӥ��9�1�IؒC���>f�ͣ�`S�/-�  _�2:j�<򂮇=���bJ�����N�i/�r��p���9Xn�oC��JbIB��谐(О0Q��>H>Ǥ�]�T�!t�� �5�&]M�c�1e�2S`ku�ȹuPEGL��F� S�J��лS�
�m�$TTal�guHAq�1��vY�c�nM�8̹r�w�cw.��;\��
���g�v�T���YvkL!��k��IUP��e��:���V����W,��c�!}a�P)��'��>�;���\�C�N�h��7��I��Hxf�|P��bzQ8�2�
:vm���ʑ�A=��3&ܼ+�1�0Vd�7���KZ�TII&J�m��2����9ԉ�������M�Ǩia�J����^�^��W��/LD�ڎ�3��C�n��U��/h���N�L��v�tZg��Qv��W"��s=G�Br��05�������5��u�c�����G�땟]��w�jS�{e�}��bXN��j{u�v5݆�̇b���&�Vn�m����r�>��Y�=��10W�Y���ͣ�ҫ�]l'w�K�t6A��9�C��ɐ�\�f�_k���8��Y�u��w{��I����yIM�b�Vo���\t[�b��C�X��X�tC̱�r��s��l4�v �Nq���{����z�G�㵆����Т��Ϫe� B�G��XZ�a�"ζn8�d��ssף0	l����@~�����P�'������R�����YC���m����o�Jyh�,�"Ɉ�������`kQ�� ���`
�>_	�gyv9퐡���g�r��q��M�G��ܦ\q��O��wV���D�P� j���x� ���n֪�@n� �aB.=3��<�Ӷ�d�^��ncDS�Q:꩚
fe��j4�z�rF��EX����S�C,:���*�I�c��� ['~m���y�*�s��.s]��t�A)E>i�>$�J V�F34�u�?��Ёg�m������OUҴ�*s�|�������o��O���tg-gY�N�����\(��x���:B���X��l��E�:"�����z�a�?s�rU���4�yպn��蟹v����e��l
PVg,�u�<+�g�Տ����i���v%�5���/������%��/t��F��C]Ϋ��U��H�uq+mn�<T��L_3$���g�2�Æ<Y��n��7չ8�p��J���֮3��by3z�X�S�+�y�=��#�| ��$3i��K3��@���2��个�Z�]�j	���%gչ�1����7���N+�ȍuLJق59�
� Ma~�.��zڊ�ǳ�A�������.XNa�m<�eA�x>Iβ�\�<�9���6��1u�z�L�U��1->�"�7l��
�0:v��,Q�?v+�E�����c:��EN����a�ƣԦ������k]u�ki<��%���0� y����k{7��O8JNdɾΚv���|0nzm���m�ʵĞ.������|j(�L�e����T-����FѬ��Ⱥ���0�����U��:u�5�`$�I�^��lG�;���_^�qҾ�!ɰ��%���;zr9�e��!mT1�B��^���RA��8�+��{��#��E��;�U�s1��ԕ|iJ`�z�#�I��8�z�C��Z�����w�� b�/�����Qjz+߁�S|����g�C���&�}���M竐)w{�3�XK%o�0���*K7z�Ъ	KvL�n�b������]�#�K�_"7~z�ʶ4���T���۩K`��3���a��6t�\ѡ�[|����}Z�o���{���žq�wШA�tݒw�� ��ܬ�%z�oI(��]v����v;�d�HÛ[�c)�+�z�ca��σG��Vs l���D�W�;0�tV;g>-e���WN�$m���)���Ov�2P���v"'��M-[��rq��[6�;I;��ə���9�L�H;��pb)�b<X�nM��`P�0��C��X4-�6+��ju< ��[�Ney]x/�������@mof�'Yq�6�#���5�N�&�Ď����������~b�E"]��vڗ(	��Iǎ�)l�K�{�iTXȵgq�/kC�\�*'u��S;�9�¦�&$5mɻ�6me�l��M��p�35�h���m�	6F*V;j�Gwr'�Zw��� y2B~���G�*k.�^�����G���q�]��bgHY�4h3�S�.�W^lQ�����/(:7��JX=p�K ��jn7��`���M4'Pqt��9E�f7�:A���k1��қA
�ƽ�C�y���~������]L��%�H>��*��E��kr���N>�J�d�U�\̭��f���e���S�6���o�}r
VYm:�c�E{�D. U��dt�+�X0����������g[r����"1��Y��ت\��u��z��A㘡��ͷ"���Ҵ<F#6c��y��[qb�Q\�ԮH�쿶��	��X٫���B@�_0OV���	2�a1�*G������z��
 �J�\8��j�7h w*���E���c�������A�CplY�H)l�[��c��4���F��\y��t���2	䝋�� ���B�~��NG	��P�yK�%��S�ܨ�wEcT��J�l��ї�ӓ[�� �eM����`M$i��k%J^=h��Cv(�5�7t*�%\�p��1)���ڻ��gnT�Ȁ�Vpr�9��-�Ѱ�2�XW�󻖱�����3���S'�F6k��](��z��Y�U�{��r�պ�g��kJ(y��Gh]�v�]J�L�>�O�}����|+�W�a$�v�g�7m�E��)DR �(����	:UZ}��%��8�T�dj�÷�Ŏ�9ԍ��>㵘���2wU���������g/Pμ�K\��yk��+���S����&�j��5�.��m��qEn�׷�<%��}y���ո[���)���K!���AXKmb�]�I^n$;or+맍�k���6���9z~���@�8����7�/V�KЭ��_�p���X���G��D֪��Z5�U��93�t7{�c�@U +�(PbF̄��) a&�qH�IM2�(fh�Hk�9Қ0C �L"�L$���H���$(�.](�i�2aΌTR���i��'.�!3�̈�&�1$���`�&�D
H��SHA1)D���l��#���H3&LF ٌ�h� B,���
d�BE��$���%$�&27u�L�� �)�	�62JiA�H�a`P̘be,r���B	ˁ�A2�����@&FD��J6fa QL��a@&H�a�JRdۢA�����
�;2��S��7�]��9оţ)Eq�)c�l���ĺ��Bc!��5�]�<wZ�{�u��F�9bsf�]��r5:��)�����_����׶�/KA{��פW��[�������^�u�W.m�nz�:�����+����}�z�:�->u�m������ە|\����������Dreģ#�i%����f�k��^������[��<ſU���/=���ݯm�m���}��~��գ{_����z��r�{��\�ux��j�W��z�|��׵����ߛ�W��5��-����ڡ�ʡ
�v�q���_����}���x����|����n�տn��_����y���y�E��|�����`꟪@��B����6���n_��s��/J������3�@��hWg��#�q��W��W�^׏����+��7����ּ^փ^����U�oJ�wϞz�����M�~}���W���_ϯ���-�W��s{���q�ڹnoU���j�[����������D|��z��6��,�S�|��O����ۛ}޻��v߭��������o�w�߭�o�~�k����=o���o�~�������{^-��}z؊��W����ͽ}�����?��_���m�_~N�� �yي�&�U�~՟='������W��ڽ-?:�4^�ە�K�����m������?[}^
��v�[���ߟ��^~u�o��!+���B4G���_}d�� ��<b$GӦ=xH��ku��)}w$z<Z|�_�w����5�����W���ޛ��x���w_���o��x�k�^->u�{�������{���y��^����|\�[w����mE�+��}���G�R�N��+Y�'羕�?K�(���nB��>��G�O��s��ס��>����{[�:�7��+�+�x��~�<�-�[ǽ�_����o~��W��U�{����[�^?��� t ��[�S��͋~����3D�q�� �`U!�D3��.\�`���z���c� �D�z~�X��#���Ei��Hﹹ��XB�������V>b�a������>���a�°}X>�������Q������DG�D�*@O�K?}�+�-� |��r���3�� �io��}m��~�>�_��i����/�|���6�߿{���[{x�ͻ������ A|D|�A"}�ӧ:���nO�l�+/u,��p��@-��j��ev_g-=t�ګ�Ύ ��t��^�̮�6�SI��+r��
�4�Ϟ�xPv`��w|�+בm���F��
K��V\��v�G{�3��au#��� d�Wo5eѝ�h�t���-��V��+\{!�3���S�_QF������}^���}}m�n.o��>���ۇ���	�)�����k{^?>��W�������}�����o�>y����j�|�篝\��}m�k�Qu����'�
�#�c�}�|�;k�_��_��?�ow�S�B�#�1C�W���1c��b>B>��3@}���na�����)(.j��=���ٸ����H���5����W��[��x��w��*�.k��w�__ͼU�r��[�ƮkǊ�_�w�}m��������ܫ��ʜ��x|G�>�����O��1���}xeܫ+����@���H��G�u0?�k�ſ^=�~�_��~-�����5�/��u_��z�-?ݱ�z�>-�W.W7��|�m���� �#�:dp>�4+�VBu��{�ڧW#������#�(�b(C�7�_w߾^�x��m������k��(�@�s��||�����T~�C��}׍ͻ�n|\�wj5��/:��؏�\�
1D�B>�/0dLx�5B�ܒ8�C�@`�D��~����E~o�����ƾ+�߾}�z�ur����i 2G�|d���q��  �ށaߚ��ֹoK�ν/M�y�s��^�z^#���}'�|G��x:sO|�3ӽ��~�G���׍�����^+�n�����|W�x���W�ţ|W��?��8�t	��ƥ@�����\�u������ݯJ�5���ޗ��o  �H
�&> ��V
��L���������9�zW��n�ߪ�]��{o�ܫ߯�������۞�������o��m��}�">�J�.�}|�}��H�,}B$G�>u��^7��o>�oJ�����3����mF>淺��A�=-�\����_����o��v��-⹿���������߯���oc~�������/��^7���h����oU�����Z-�\��|��o���s>}�o;����+�ߞ(�����_�=T��>����1�3B>�>��Cg�8b(G�	�������/Mx����ߋ�Ѿ/�u�[�x�_������_���}�>ur���k��*���w�ߝ���m⯋����w������7*^3�f�B�~����Kj?���û���̺r:3�7�2`�-���!E�M���2����_=r�wM�8�C��1/��7)���Nݙ{�����\9�]r��ʸ��l8�r�[7�	B�k�zl��T�]Y���ed����>v��,G\���>�>��4@1��%�r}Q������^��n�ߞW~��Mp׿��+�ܼ^+���:�7�7���������o���o���Z�/~{����o�toZS��:��ɷ55C��[1����k�� ��L��`t\}��~�hT `|b�cTP��G�1����߭�owϾ_����s~�����ڮ]�m��ڹo���_�u��_�k��w��0�t�>aNm�������ѣ�"G��#}k��k��/����lEz����W�������׭��W.��w�}no�����}�彯k}W�����ߊ�W�ʎ�c��>��]UAX*��@�ӳ�)��9 �����(�ypN(�}���ƾ����j-���z~6����A��c﨟�A���>����~��]%�AW��_}{[��W�N����;���׋�z��F�_��}���_志�>��^���麿gfbf����>������𥳐?��^v�*�����y������~{��o^�����o����ǟ�o�xޛr������kF���_�=z���^5�����-�o����ٱ羛��X�KyEd����}}��_|��_���Z/{��>+�ߍ���^��W-��->u�����/O���|\ߞ��ץ���ƿ-���\�;o{��KzW+�n�����ﭾ/��}�s[�T��ػ�ޛ2!�"��no��|��{U�w���~���?��_!!��0DR1�����$|�H��gx��x�k��{�-�E�+ŧ�ץ��||[�_�߯/M��7���K��7^�Q(ۿZ�o�ԓ�
�`}P���ﭽ��~�ſ�z��o־W����^._[�?>����{U�s�������E��?�W��oKϝ�����ݷ���������m�����?�-�_���غ��N�,�{z{�*����{�׭_���׋������ѽ/�+��`z>>�v�d������U�2���*Pd
�H�ad:+�]��Cd�)��P(�P���9���N�0�xy����Q;S�fD!tf4�bӒø��ȯfn�X�'N�Es�]c�?�:�uZӱv
+����7���.6�;����ʴ���RF��j�h[Z-�����u��q/���'
������(B���q�_K|�rk9�������EÐ�:���3����>�����o� ̚7 ���[4.��p
]:>T���-Yg>c&cӛ����3�ִ�E�g��r�:��9#݁�X�(s4��p��Ɉp�3���j�z6�wV�E=WdI	�^{~�"��w����3u��7Tz�59�6�xbc� Az{�]{�YR�s�Qw��q:�8`��
p��ˇ#sJߠ���Ȯ��D�C��Q������{D����q��P��V�S������z�n?Xif *Tqp��1�N9�4Б+���u�.��:o�)������釦.18�g5�1+>ډI�`�1P���1D�s�v(�,Gp2pu�Y�漰���P�ݕ}Q���<���\�<���ۣ�-A������K�큯�xu�Xd4Ff�P}�`L�*'�xU7�2_��Cct����ry]n��A�z7N4���q�k���H�1��ϊ���Rꏂ���x�][�䎼}���:�39$�ϕ&��-�����s�o�Y��g�k�<_��]��+�̯0+��lbfYŢ8m͑���Rn�jJ�r�+u��R3�ݚ*���Dͧo�Uk-ɽ��z(=j��J�4�y���������n}Iv�����g1���,ùbfJ�,�00���61If����ڷ֨��(�8)e���t:��_U^:��D�@�8O��@V!-�6`�������n�!&:��3B˝�Ƒ�x6)�޵[�𦏇x؁B�:xz9�e�Ϡh�6��p��)�e��g�Y�*g�R�m�{�[�̡rA�����>�U���n���.(<0_=v�h�:����j�WAv�ڞˋ�K~�uR��*� i�rt8T���,g_L�o�o��S�ѭ��y jH��_r��7��ɘ,�" zQ@���h򺠪k��n��)i0%�ʞ���W˕�'�/i��&��Z��E_�dHB�� .5�#L��|ͳ8��ۼ�~Cs���{n!0w�L�ks���p/ :��E�'v�S6�cA����G|hͶ+F�:�b�RV��4�5��|�L��2d���!��(��c�Xu�=1�Yg'�5lݽ�|�P��b��;;�눖�\d�=�uRwtb��?2j� ��;��
���=�X�+�~�װ!�<�
#�j�n��tja���x���lAwS쌍N�#8�5����ޕxr�'�k��<)���'�ֽ�RY7K�6l��8{;[_h9}\�&�}s��������7]0H�N����>�{�S�)�^l1C�v�K�R�g�(�y[���W�f�}d4i��[J/����}N�'r'3']��� ,�|2�W�G��jx9�IQ�ע��7	��a�A9V~�0Ժj�ň0x��U�(�gk��%]��ӡ�R��>�)�ۡ^{�{N�S�0H�ey�7�5kG�OZN�����䝮U٤ qͻc"UB�k��ok�_=��z�\�QѸ�aek����F�|�L���J���tb��.P(��*��; �1�p���m��1+G�r|�Y�Ó����N��/ϭ/EYj@��*�Q�K.�e�����P�64 �W�f�s9��f��K�� ��
K���.���������y��4!ŀ//0(��6���F�������g�a�Leh=�iT	sΏrw�~��Z�ޕ��X��w�Ն�(�Ø�p��۸y�������R�)��B4dcjDT���	�g�Jk�Q�3�yTpe�>:ܑ�T=�#���'U.o� &�	]�v欑*�^s�&i�υ����1ȿ��_֥�G���s���n�u׭ؤ�L�3�c\�"c�A�ru;�%�<0��m-��E.y[�3��8�$�k�e�t��Z�K�Pb�o��ۉ��!`�ܲ9��E��S4o7�jm��K;#"� ���^�me��F�ާZD�â�Ƿ۹h�z�L����8��~�3��Z���W�;�����
=+M���̡��/�F&B]ms1��ͲS`(n���P�F N?_��ɣ(=�=�$GujcUA�i�/��hA8�kjI�</©ybɴf�3�h��i�.�&�<� ʺ��p�����DW?��h�Uc%K�B���1i+��l�����46����:e�O �������A�w��=uB�N��Η�a�`�m�<�dfWjӲg)��5���MՈ�n�3q�vn!������`ߠ!��5�|Ē�?1'����v��T��aﮍ���;�h�̵W�9�'@Cꘞȇ���ʉq΀8`ǟ/q�[�Le@�]=��wZ�9�Ƙ�on}�5ȁ�%�e��#{]v^��C2��yEҚ�R��F�����ۯ�_Bq|��c�u�����fN��B/(4܂FZX�=ks���NL/�T��\�S<2���QD#�4F��61O2�:�ʇ55́��4�>�$̚�8��dA��0�ʮ6(�
��|>�� +��3ҧ���ۥb����UX�H]�=�0<;�y�\�3��+�-�2f�ث�66��!»�Mt4f��΂��3ݒ�>����G{�\\(r���+q��͍����igt�*����{V=ySq`�͓�ŖU�Ɛ�����@ᨲr������r�r/OV��Nh�^�P�_�i���秢epY �(�Џz���`>0���EP@����/�u�%��f�C�T��!����zn�!���j=��9_��)��3M��=q^�Z��7eC���n��a��\s��Dm|�܌�wV���D�L�,�~�	Խy<��E����$T<��xD,=��C�t� ^�����MGBĖBrH�� ��Tݴ�u**���Xϯ�xnP<%���'H �rՖwoG4�z��p�F'۾= -ﻥ�N+�N��?3u\�Q�Q:<��fi��A��h@������7k2��sݼ���ݦJ�X�̊�����Q[�7��6z�:S��ta����̀YY�ܝ��C���&���TBr����qFΡ�W ����fáj5hߩc���j ��.�����c�m�=�U��:����̋Z�l��`�t��&@�u�^�"B�ß�D�`˩ZN��<�^�_׽0�����s9���YQ#dd.�[h�k�x�V2�w�|�Մ�����̾��^_>���^���ވxt�"�1n��2_�Jޱ�p3�[�ض���V���h����7u�q���:J���T�Ys�'N$�8Kwj�����&p)i] �*�|TG��Cr�T���X�>�R	��0�LX=uMg����X�
��*��$�Y}u{�1�$�-� ��;����᷉a����eW��Y����R��(	��W���9��۽:�nK�ck$�� ���!��x�=��u�;���yE}�Qj�����g���n3��+�].2ʠ܈��)�R�k�۲յ�g��gn*9 �dߛHN�x�L^w:{&�>ʽ?:��L`TaBsq�6b�Z�;m�\�(�P� ��"J>�NiŒ��{ܯpEwS�.I ���%����rzr�Ci�p�&�})+1�{;�"�[ِu�M��O��*'@UB.�$UtҮ�r?�����g�莞Lpe1{[i[���L�G�x�Du�ʖT 9q\
�����0R�������BU{:ҧ&[�\�L����wo]��N/�T���=���*��aB�!���L�%��I ����2����c_6�@��cȫ2$!\`Ɖf
u�L7x��t�9ÑN`��c����e����3Dr��{�<>z��w�m��X�\/;��ڭ�˞�|:;dGZ��z��r��g�1�d����<��9��jV\�r��`�q{:���k�7�R1���(�q8�k.�ʓ�����������g�g&CB%i�🐘��P�*�MCn��ֆB(N�j�L\!q�u#��
-�;3�z�-}꣜�;kQ�7^��g턺�RR�2o�����`l"w#Gg����95�c^/LU��������u�����Ww�����~d��ܸU�ʩ�1M�kl�k��Y�([��t�L؂:�L=��+�+����F���k�Z��}�r�K$lO>�Җ��J�Oh8��8��+O;ʫ<�'����s+��`9YH1��k4�!3u7��V���J��G����s�Ѓ�O���Q�ɴU{Hm}���g?b���ik�XO@���ȅUP�1�g�ڗS�%ʥ�E�x��bC7�w��H��^���e�k������5S���� ��ǔ�LC�ٌ����*1��<0�.5�j2_\�Z�T��|t�&��<=���T���u�:�B||��ܶT�_i8�\&&�V��m�M��4 (��b�����\%�(Wb�#�Z����鏱Ô-��ڎب5�LNƭYQѩ�"��*]��4��R�l*���h\��V��)B�����!I�ѡ&q�e�U��ԏM�4p�Q&����u6�;)�M)�,"tpYT�T<%^ӉGtv!*k���|Xg5��4%�]e��M�$�\p}`�YA���C�z(�`������0��O��n�v1�Y�W-J��ݡ�Ga���c��H5QZĎ퉍��ԳL�[!ОeD��n�ɣ�D��Ѧ鏮�f�<��[�Jjf�4��毷y�+Q��+#ͽ3�xo�F��&��PZ��f�`唥n7kBu}r�=�/����(o5��R��Mv�)qΩ��KOy=6���əGWˠОAt�ޥ������A]���}�p�ԣ��f���YYy�Z#���[z&q{;u]2I�[R��IGd��F�bm�̡�D���*ì���J�hE���]t�v� ��WA�׹#�AS�ʸ6+m��#B�t�u�}g!!qj�H���x)n�{�q�۸r�t9Ҧ���V��N����m��4��[���M��(�ɚ-�4@��2��5pjC��r������)�u����fouW� S�Րv����3�)��~�P��N��֟ɮ=YuŞpL�k�!�`��O�:�؜5+���u�Ҕr	'�6���j.��	hVpO��^dP�<ޤ��|*�Ώ-�Y��o����䆦e)Vu3s/7䁐`Ǥt(a�hʖI�-��L��}�@�Y3�d �{�PXoK��ǁ���%yc�,`�hS�w�L5��RZ���ݓ൤�5�9�[�X������n/���\�����M�}�*}Y�q��!�V��qR滫|��zv
N�Ȧ�����7�`t��1q���s��P�z�c��$Wq�3x�-����=���w��������"ǀ�Z:����>R`J��b.���z�2�I U�����J
�d���|�&bTJ�d��Xr2Vm��@�H�n�E]C�n�F�����Ꮪ��0�� �<;�w�B���T{��1 �>�w,�ќMA�q��2+�t-·n8	��7��t�r�F��#� ��j�ż��R�a��J�/�7v�.x�:���bw��ś���F��}�@U�}��̧�n9E��yir�l��̨�cU�[j��s���w�at����ԁ��h<�\7�o�T=�]2���2�ص:*aw+(���U����u��G9CyQ)��>b}�\9|��O,U�] ��c�M�l..h��?*=nO��j���9���%��U��6��۷�Gz����J��s�`�Cٺ�=˒�d����"*�|&�ͱ@�0
җ �.='47r����,�)�O������mA1��6E�$����-�s-�m�m�I[���{�-27r�bse�u�]�����������L$��	1�)4 AL��$ DIK&�Y#��DfhLi"Ĉ2,Jd"�+��Ab2XMy�A)��EE����!E���l)�M�P��]r�I5�M$0��q�w5��������Ȋ2ȗ5ԍwt���A	�MH���H�b&Q^y��TD��Г��M˒c�Le�U�u��G�٠4EA�d��13F��B)�إ�p�pH�y���%�$˻�봐;�bK��]ܢM&�S+��D�:�,Q2$P�`FBY�2b�#h$0�Rd�����1��ȃ$���$э�!�����P�I�&(LiF��i4e�
SI7u��ٙI`D��'�����םHF:�&��!vNe���^�m�C-�,�MG��k�p؃�pm� ���R�Od��̆��ΐT�ﾨ��Ԋ��ɓRD3�����9�G끶j8�4�P>����K�{.L�"i���Qz��9�c����+�7�Q�sn����(��9I��)�.R=2��8�+�u�%U=c���'v�Pt�\M���pU���������0'Sͯ+�  T>��Er��(�{j9ms��Ц^�~����93�>]�|\膎9��nw#�Ո�`��]S����]S����7��$�KIzX���0��h�c�0��d�����5�:���]����a�C�sn�D��v�;<3��sA\Ƥ�D$��Z���b3�wn{�+z�Gj�pT��#8@t��o�]CQ��V�{M�����x%�
��NW�v��읭Y'�ЍJC Я�?K[W�<��+Et���� tuטԧt3�\��n>�S�r�՜	9���e��vn!���Q�A=@�|o���'��|�j��Y�첅X�0�5y{h`!�I���:�'���2(s�&.���6Dr*�T�vF�U�r��2�;ݜ��4�?��Y�0a�IM���K�&H�U�ۇ;�L����E���իp�y���Yl4\�R@��Y�ΘZ,�l�����cM��á]DS����N��W@\q������Iw �y��\6��9��}��_W܄���t���ɎZ�(N'N��Y��]S\�1��2�k�]v��(W:��r-���g�t�Uo��Y<2��Ғ�p_�!�Z S_�/>�z��x�_���w�
�1���l��������e>L(r�V
��+�]��_��(�{b2h>���@�;�'y���"�b��m@˙=g�:r��\�3�*����h
�~�Q\�i{��
����bRy�K�DP��"��ϵ��oi������U��d`��{L�;H��f� %Q��_�5��J��
f�Y�B��Sì�c�!鸇�HvD�����G�� '*ά*��f��E��",&s�2�g"�ۉ����yai_C�"6�;����Ol��'\j�V���۰	���*��fu��g�B���R�#	�/ND71�Dk�ג�5�vfI;WF ޥ�[I(}R�ʁhw�1�N*��v�-G'���#\�
w-E�[B�
�<X"�4ۿ��u�
����!+	�t9-���<���1��N�%A齵��:�WoJ�K�<}Խ�{�+��-�<�^h��e{tuq�"�+�֙��Z�H��)dlF��8V�yR�Cp�t�PY�.��X��X���b�l�d�Cx�jܭ�sb}iw��&�'@˙.�5���;�Vh�����#�-�i�qTA�8.?~m��9`w��V����ߙ�(�q����ޘ�ӊ{t9�����LZ�b�S~�C!%WGМ�4�Fhe��a�<���������n-2wu�|$U�:n����H*��s��v.��#PW�6�ļæ�	֙i,�9��b `Y���f-����|��Ǜ�8+�T�ޭ�	�wם	�;0��Vp;��	��5b����&}�5��XpLk<~0�7�� �y�ʂ$�}73�ao�5�Yݱ:�}Z�ǫ���9�b��o��DfYU�Vq��OӋ�����Cb��'�i�[:O ���T���5�����|��\k]t�Y�%h?P���PX�5�^Ĳѹ�����HF)?��$c LF�nj����m}^�~�^�v� �`�ݶy���[\�P�ߟ�&-��3Y2�^�@TaBsm�6b�c�m𿒜�N�v���&���c�^�l-��C�G�(r6�f�;zr9�g�u-ot5��1�=�����+W�z<�¯`�8F:>q{�Vލ9�f�:,���)�Y�9*+�-{xVe�Q�t�
������F=��'�{���ن��&hx�v�C��l�y�	�JQ;�ɸE�#�ǒ�+K�ZtPI'�j����ԇV+��U}��W���=wf�l���8%��l�H��h�ē̥?R,`玗P��p+�!9J�y��G4���1��^9�@�(� fz+�[6�]�ޅq�^]�mN�G=�jtcn���z�'�L��3����	B��Xb�<�z_e�=�1�)�:7�5�FSN��&�/k�������7�y_���Aq�'D�,+�����kx�ۣܟ����Ϭ�[���Ur��-��\9���S�`�*�u1�yn/�R��k�k6\��$Eag�Ẽ58�7Zf����ΐu"�%������֓͊�,�n��T�H@Ȭm�,�^`_/)���X/i�f]I<�53��ϣ�Q>����q ��{���b���j��U�?�{���0c��؃�m�u�����y�x�l���@Qna���V��u�"9�'c݀�WS�0m^G��=0���o}<���A�u����`���sB��ԝ��̎u�{���F�������ֵzp<+#�o_S
�*�0�JA�ҋ�T�z��t��>�T�\չ,R�Z���|Æ-�:SY�޸;�k��o{W����Qo1�#t�nJ@y�d_s<@�����q��J�=]��|���B^e��u��������$Vt,K/6�0����}�U}^�I�=�4��^�#�u�����c�|�������mH�yE*F�����Y���C�bXk���g�j}�oW2
�!��^%Q�9�]��O=͓����3��r�/$�%��:��cb��£1��P*"Yt[-�|-��m�^���rl�=H+����x��E/�ȃ̯`�P?����^�뉊�Z|�>FsN�ʬ�cG��;�qT"�j`3�ڸ}�����!���3�P�1�P4��^yV��lJMng��9��g�HK�0Zq-zJ9�c���:�ò���1�7�)Pq9���o�|�|�������rˉ�Jㅕt��rFiQf���(Js2�a Ajj�+���ˑ���c�m��b�=Yaq�������G ����Vp۹�hD�S6���}3�gq�e7� �&C���7����%ic >=t�T�[G�p�. ��J���6������`zk�(\m�I��a��1XS9�2DƤū�X��Jc���M���w�+8=�{�X2�Ǻ�m�8�o1�א��Z�:��%�\���9u9���v��q���lY7>}��fp���_�
Z��7p3rn�Q����1�NV�J����zI>4�xs/z�<�e[
�<;��n�Η��\���3��H�U�����#ﯧ�sK��Q�t���#U�5ɲw����\�f�)��}e�3�aEgD��L=�ɼk����w��U!���� ;�g��e@��d���]	�?TD��7F��e�@�{��o����q��
�5e�Ub/���C���f�nhECC*DW����6��&_�7���'u��:�Uo��kE+�j���v��C�I:���1=��١��$\�3�1��v_���q� pJDa��Xޛ�}	�u��_���i� g��o��7T�qC�[F��e���6�՗�2��b�ǅ��:w"e��?,�&n��RM�<�p}u�x��2�d$�Z�z���пZ�Z��{5�Ʌ
�R]��+L��b��C�P�
����'��e�]I�s�N��L�NS=���zaU�i�M��,�������Ծ)>w��@nQ�����j[�'4��!��ϵD�oi������VT����L�1T���hlx��4�f����6҃�ʲ�6/Y����M��C�%���l䕓d��u��O��}�7I��r�������W%gu��G&XѥY�EB-�Q�HYպ��(+7u�O׮�Y�P���]����q](��i���p�q./2 �u�jr�؉f�Z/-�o�mMc9_3e�I&��uЇ�������`��� > w����,�@ -���8|ǇB�\g�UɷJ�f�Ƽ9�2Eo���CTf��Nos^�d$���Z�@q���H�P���!i��hy�m��'4�.�S˪�%|=�����`��T�s|P�m�n�+�����.�U�떏�0I���_��.���|08/��pl��m��Nm�U©�G�!.	�ty�3M$Ǵ�9����zm�[��k�H��g���-,rP	�W݇}���z!�Mb�!�]{�գ��A��	�������:������#�o�`a}�dY��a���h�Ɂ"#���p��P��[�y��i��1�6!^�ӟjt�qX5��j쁀������R�i?Q�pG�k>��{U�[��a��է~��W��U��s4��0JH��{|��ivJHM��D���0M�� ��tY�������λ��諮�uOi�Ƕ��T"�76ۡ�R`�%:��4�-�kL_�o�L��f��P�3�)K=��A�X{���3��1���wu֏D��m��h�H�b,v7�K� ��i�%�׻R���(�ꮲ�,]#��!(`��Y�0��������r�SYK��.w�8���k�|re�LT�:�z�gW[Ti�����B�r���7R}�}�}|s�SMu8�&@ԩ<���2]F���u���ãZ�s�1���+��*?	wX�n���WQ�{޳���zf�2x b o)��[�#�W�m�Q���Ğ.�cH�;N�N�T�x\U���P9�ɖ;B�7
����1q-S���k�6=�n �s"����z����-U	Υ��
h�t7B
uY=~ӕ�A�� h�6ҡ����;ܩ�n��1c�䵙���;�/�`!��r����n�r?�����8�Yj���=sėT�}�Zrt��s��I�1��K*��`P� qjz+��1��ʦ�F���j�US"k��������t�z�'��*��Q	�j�� h	HX�^�'z^�ٹ�%N���h��
����+䚴2��c!����n�6���C@t8C�^��v7�wu��&8Y�Q�x��������U}�Ժ���۞��0E��X���)��\������b��4n�xR��E�!R_��V��f�����BE2d�7�ޣ=n�h�}��7��;���2���KpjuW���<6�I����q+��O70_�FQ輎e�L�O����Y��Z�>s�����/I�ChG;'28��33o&�>��lɂ�V�s�ɂ��o{ h+oE�����ޙ��1-��m���������'��ɯ@���?�/��㋅Xc�r�~3����4�;u6O]�U�e�0��3x'{v��N}ĸjzۈn�m�� >6(��jnPU�3^Á��ƯL3tG�]m�Noޝ��'��m�H�!�na����i��u�>� ��?s�sDk�bv��5��_�2�=����X6�b��8lq�p������=k�w��U<�f�����2X������E)q*v���V8?v>w
g�\AO_d7�����w����b����^��Q`Y�L��d�}X��b��|��)�M����~g��[`����u7�f��gv�t�w:2���H���;�~�)VN�n���),�Wحԓ����^O��ߡ5��+������I|�"��9�ݧ�9R�÷o�W8�ȓ�چ�����z���e.o���)L���� Wa�Hq4��'���ys����[O8�Ct�m��Cb��dn���	~N6����Y �sxe\����S�B�`V�t�V��|��dʖ�V��v��X���7F��˞#nfP��5�\��J�ܐ�0�.��.L�r�e���½�;J��6�aM]�U��*�!J]#��"��u؏P��b'��P;Ղ��E��������̒��8;�n߾���Es�P�wB��ؼV��t�Br_&�h��QMV���T�읈��dHm���l�ٺ�KJ�K�g0Wͳ��5:�Ӻ�R�0Nˍ�9�>�`r�Z���/�������꺵9t/j<��*h��7JK��D��%�j���]5oy쇂��kYFГ:��gw[�X	���
�7���l].��?��s��|f��T��Qw���g3�w+���Z��.�qi�5��h�S�<����Zp��:$�Z���ܧ/�^�e[�s��'��s��ֆ���o����Ţ�s��8ۀ�vU�߳��ej���'�1�=q�ۏ2�1�;��8�����9s�T�g*��X�w�?�Q�~�r](Og��`$����t��<AiI3�w��u�a�C�-N!��z���yUY�hL�WWK��
b�fD9AR����ɼ�WVDv}c
��m]� m����Y�{��Ȼ�� �tC�O���Z����\�Mf�y�:������Hovfto,��c]�����!�"����BsDs��o�t���8�
��&�kL���`�&�Zɺ�~v���YE��9�����w��U����R�H�]w�	��<��N�W�ht�=8*v35dE��Ϋ�c8;��J���-�"��2�fT�p�#�Z��T6��b�+{�]���^�˼�Z�U��&{0{�+x)���t��hӬ��A�z.��Z�E҇s�[�f���jM���GV'n�Pͦ屯\ݡ����ir<eTq;ߍM�wF	���Aa�wEv�?��G��b�V�q��HN���7%Z�WA}���Zf"h�3%�V6�iQ_I�tc0�$7��]z�F�[�]
�[��Fk�t1T�����XZ��ť=`,��p�QRx��Q��]�,S����8f��a��.�(�t�&V�&�]T�*-��.�]
�qWg���y���F�t7V�B������5��Ƿ굪��g�{@u�(<�������EE��.�A�������p8�#c�muu!�I:ځԓr�ra���ҷ��:�h����
t�QQ;��}@��=O:�=����p���P��nˡ�$��Q8n�+O�H2�u�ݍ�۹�����fkq٭�f(��^�,�|���w�l7YtY}:qa̽��h���eYA9ݍ��'��g�ֈ� ��\a��Nj��7�v�nT]��]f��%!�a#��#�LwPoV�Z
8CIu�+�y�ܸP���ɐh]h����DӺڳ��.��kiݘ�?	+�\�/���q���=U��fLޠhX�.g\�Zt�1�ۺ��,�YMX���{��x�Ƴ��d0����-������%����nň��2=�,8�	u�م�na�9��lFr89J�hظ��/�%���ظ���].��n��l��n�Z*�ڬ��;�siVK�]tu�V�T�2Ep�{+�{��"Ż��[��7
�J�;/�Et��%{��l�
T1�j�եC6��'i�bsw*���n�t(ІP#;��v�GYm�ķ���
�C�ٽ��[�A�r _e�D��fN0d@��0�[�=tjps���2a�N1�ޫ�OyB�T��� �� �d%�Yr�酽'r6���ս֔�KK�a����]����e�/h81��K��:N��e�Т�lb�xy�B�k�QwEF�5����t�g.��%VmJ��Ǭ']+����ȴA�!�u����rl��(�)	�ƛW���wXU��Sn`�r�L+J#%�ƚ9����xoc����f���;���J[�^��An��9s�+R碁�s�\�I�j�p�(�q=v���d�	O)��]�[����s`Z�v,��Hk�lȨ�Q��,bE��&����1���$*��h�����H-^u�)�#DhH�l	Awv#A%"�M)�E��$-$0�LIb��"6�vAI ��^uѳBfh��E1<��o:��C"2M*)$��$�%��Hr�f���6�$�1Q�Ÿ�)�q$ �&I!��	J4Rh�J%�&)e��B׍͉0lX4��.�yݙ�"�ŉ9�I�52b0����B�t4�q��AQ�5rB13��0
L�9[���M&�Ƃ�̍���wr�$��ܒ��9&�h���w%�y܈�l�L)�d,_߽������������B-�Ίӏ9���&r��`�;��p}2X@薧�t���+E�M��Z�٬�+�pBk5�������}�Л��Sv6�IY���d�Ͷ������u9Vn{&�WI�ɼ�3{���Z��Q�j�	ŷ�ʦ�\K��g&�{�*Q聝J�bx>�~�s_M�G�nk��N��	V����}q->���+�m�P��Z�ݪd���)�c:D��xs�(˙����N$�W�R�k��Ƹkm�{_<�������/H��sI�w�z^>���gڤ��O�%_I��+������"�K��띐{x�q�N@+R��4�뾜)��T�X�c��K	i�F�"��3������t�g�]��G=��Z���5��6np����IK�M+�7��6�o#b۔K��!u|#L�b�H�a�Kʧ��ܾ[��5Nw_r�[|ƻF�S�*ۚ�_pF��YNkqqHP��.ud���~�x�%SV��q�ќ�A��'Y]���a�{�V��8)�7X����3gh&�=^8�Ǒ�GRa-	�f�SÉ�͡�;U�I(��\��1��W	�"S���;~�c.ʔzE����8� ��� _l�(A����,��&���UwGd��t��P^����#�����������◎�
ٿ}��m�D�eK�5�&#��o9���jہ��c�;�S�`�|���u̅oTa���0-�f-��T�F��^���}^�Sj�����D�w6��s���f��_FbϦ��J����M��R�5r��$�p�Vo���<�~�{NU�a�T<r���ËҪ���@����������q��\��z�"���X��],+n�5m1u��8�5[
Ӟ�R2e�K�p���#Lo.ne���f�5�����եl5*�弹��q������%G*������A9m�Q->�sV͸ޙ�2��N�n�V7����莝uH�%��JQ��7��ǍMe�R!E�ہ�Em�h�����f��eR���;���I�w��im���ɻo9ּ*��v��6�q�N����}�N��%7�M�ŗ��&����yw���s��˚����1 -+ X�*L��3��N�o������B�e��j]%�h�a����֞K2]���E]�0��kx�i҇K偉Ə[lQu�5ǻ*��Ӱ0�f�ygS�wSt�k��bS���v��_��ﾯ���ƹ�<���>�/��ĳ���D:�5	�t�k�q�b��tf�׼�繀;a�;qM�{?vht�J�j���snk��Q�&,�㵴����"E[����^�\�"�J���i���xôn0�e�뉆�2�k�B$��^�P�Ά����^�N�b��2�I0G'�+�f��;�)�v'�T4���+s��Pے�2�<�œ�V�C��t]P��ܚn^���&l���qƾm�ڮ���K}`�k��f53ڻql7��wu���z�+���T�m���18f��;7;ήk\�o�f(�'���s�F/4�ؽ�H�VyZ�S٫_�L�Va'���=q�r������ݩusNn��
%��{�!D�agTM�TN��P~�|�	���U�'�<�x��>��5Lح�s�OV{N�n�����^璹P����SO�茵�8���t++;�6�5"%<�5��V��J�i�q�Lso���n�e�u*Жml
/�j��Ċ�U�Yx"�x��ǎ��Zf�X�X�h.w}.;}3U�	w5��S[V�b]�@�:7��+�p�EU���7�k�e��;+Y������}�d�8"�N�S��{��_��w3-P;>�N��*�{k,�gi�[�@mL�[-6����+:�潕p����g]#%�^�mY�++.��u�qQ�MRp�Wx�z7�8��UB�ب���7u��s��.C�'{���<㭕;n�U/M�)(�+a}Ȋ���p���;�[�rj
�̄�b��+��,}��·��K�[����m��;�z�yfc��e�ئi��H��l-��U��pjX��	��i����[��kQ�1�%r�L�]#�P#c�M�ח��}�TB\֯�;���8�8`�C�<����a_l�/z�\K��9�j��'���׷knA�ޭְ�� ��RR�ƻ�n���G��ԕ����..iBT�s�ùJ��c�Yf7f\n��W	*������ʇ�"c���)nk�[MfA���N�'Gyu����TN�j�ʇ��i���'4jݹ���s4�bؑ�m�3GD�k�U������6��Uޫ�Ռ�l2{JH��$zvn�wΖ��ͧ�>M�0goB���;̶����x��ގ���|Mq����菣� +f�[-	=�Y�;�n5d�U���u��2�\�;P��C�����pE�����Ӯ���TΨ�쨕�*3�d�؎�yi8猳���j��Mq�IO]��}�wӖ��� f*���3���t�ϲ%:�����<��u�=VL�i���}���SØ1��nr�C�Qs�vB@)u�wkw5&rI�ܤ��i�K�ۆ�������W �s��ޑי��{W��p�D��K��c����̴�/OL��.���P9���͌^]�ϳ
쵔6��I�\'����Wq�ˇ���O��]l�_u;A��i!}4,eA�i��[�/�ҔkyF�km�Oj��:.��{NǓ9�y�Q"ƟU�.���`��$4�O'qIa��+���t���O!K$�א�{]��� d��g+�TՇ��/�I�!(�Ϧ��Ǭ�j���U���5�,fS*aRxp7���㎜zj��z���˯_pn֛1�M�N0{W������>ǻ�y+�1[�|b��=#}r���1�4��.)Sz�oi�喳�s���qKM�*���0v,�i�8�ؓy���j��
�3����1�ޗ�����c��otW�ڗLҙ*��\��	殗?m�),Ol�ͿS}EΤ1�i\�;f�m�o�m�B�su�b����Fߝ��S�_�@Mh�ܸ���r�[o���k�n&�+�6��s�˨�t*�x�T�$HZ�
���ԥ�X�w^+IT�L��k���[�{Z����r������[��υɶ���싖G���{Z�W����}��k$5����Bq!��,t�oeCWP�U/2�`��sYV��>��4��'������6̝Ĕjx垸�;_'y7��{�3}6��`��U���{g����իFa�6�ÙX-'����׷n�mBzwl���J���p�uׯ�쯮�����#�p��_8��z�>o7�9�cY=�_i��Y�Y��s��>�E��Z�-(]X�b��ys7+��*y��+T�r�]x"�-��;׽(Ln1�DIZ�:������>��j��Lf;Ѧ�1��P�Bv[@Y�0(1����'�9��4$8�˽�S��:o�*��5t}��on�D�$˝:��`��`���G�i\��ABQ�U]`�
���ﾏ��y�b!f'F�^��%�W%�D����Q7�'7�Վ(��U0�Z��ֵ�"��9�����r��=:ђ�/N\x�����
!q��N���������q�=�m=�S���*� � �� 4����.��O
�ݗܦnI�,���<k��y�*��n���ߒ�����PJ��zƾ+�,'1֔��Wu�c�o0;g:�)���_/)�5C;�s��rDS�[���f;4*I���C9����_9�#;1m�RZ��֫�oNf]�ݡ`%�_J��	���UB\�Co����VӸ�1��B�wں������u�^��q�5��7��I�N+��W.�P���3k�TrZ��]���F�f�_���nz_FP[w�)��س��-[jbEPY��S��\U�;��SV�3M�Q�r��ȝvT
[�b}�'1�ӡ.i�?J��N�b��U�>�͇<���s�D/h�O>��F�T�j������گ<�mo
�ɥ�u�-v ~=�o+�0亝5JF����k�+�讇1�[�:��s-uN5x��Ҭtۘ�km�(p��A�6��c��'G���}�}X�sq��Ѕ�x��YW��+o�N�,�;\�&��p2`[���W,��qͥ4)'/6�����++U�L��笳��r��V,d�-�k{�xJ��ݐ�ÎZObnr�Z_b��v>h�q�S�m�l��/Z)�X�>�Օ@O=W��;���˜�P��GO�Lo>p��Y]u�{��U���wc�y�ެk'���_p5\���uFK�}Y�!J�w��2�fp[.o�_>���[.x��A�R{���W3�B�S�m��?W�,��:���B��΅9��m���amJ�g�{rd��>�L�hz�R3���<���y��St��6�qNMJ����i��⃪;�(U�����y�R��,}��·����_�7�5�{$���VDu�}����g�X�}��W��E�k嵧o��^s��0���������:��wx�������B��C�}r#�s��6QǪ��q��"̧�T�cI���:�������.9Q��jW��뭫�(�Z�<�#�{Y[��8k��pk�KKƧO�̶���ybm�D�u�E�ę=�����!M�������z#q8�����mw�Z����3t���ʤ���z�r���gXW�
ᜉ~���'mvo��N�h�Չ��Y*[���N!�y���&��hTd6.'�v�}!���������3� �l��q�c�cIL�p���k���T����2v�NR6�{���gZ�ʗ�u^�YV���bp�D<�;mΪ·}�ڇ)z��܃w�)� �{e�:�����j��Z����S�L��u�u^��3�i��\��z]������������>�>��^����rV�3Ufu'cf䕰�z�/7��TF;���=;���3�M�TD�|1ӡ)�vneg5Ԣ��8M�P��)���6�oz����ܚ8�ָ��}�~q�{�5J��˛���}q/�\�P�52��~��/c�%R�n��+�I'׷j�5у{l�Q ķ&H2Lb��6�e_A�����y^lUH�\��}8�c9*�4�V�,фZ�O�|,��u���ۑ�D�ar��m�Y�����F ZAis���L�M}�K+)�jt�.vr�*�o�t�{9�.7�Q��#ﾌn����T��
�%�DJ�U���꾾�n��}r��o�*��"2�\��|ϕ;�`r/�Z/�Ҕk�I�Ƹkn����Ĩ�Vھ��l�WA^k��B��ب�~F�O),��N̠^<�ҕz���מ�f�����x��J���}�F��(����Qx���:�:{�SS �8RҸ5�C{���:\���J����!���W���՚�oծ�/%��Wu�Z�s١�M+�w���snj˚�'H�q
r��j\X�zG�3nj'�MF7?gqU����a��#p�1SwS�M^�vv���рV��3j��{�_Ky8�"3^$��DZ�
n1�|L���:�v��,�\@V�\?��]K����7mv�]oj����r�%X.�`wkL����]j!�ʍq�Z�t�]P3yy���������t*��ڙ.��Q`�R#��$UŢ��Y��ojU��^J����ӏ��̇p�aPr��k��x�r�9�cr�Ui��C�WS�=��(��+�e$�s:FR�1��{2ػR�s\kx��'+i�@X��[��¶��7��۷v0]�����S9�RE�E�t���k]�
}	k,��J#��E�7/x!�	�Hؚ�g�Y�����bm�&T�G��ٳTt� �EnC+o7��f��d�V6�J������4�$n�S�y�n����H\vV������4`]�lX�K������n%�tQ����p0!�sg�Ħ���t�$*_u\x��֌�y*ݶ����PZTK ��m�:؀2YU�y[�-5�2⢭bcu��B�)=�{�3i����L�u1n\ Q�l�,�n�U�m���,Co*�F���xT�tՎh
Z�T�[{�1rvr�X��7&���*�E�������_�1EW�#\-ޓ�؋�jv�g*�ʂ�#M��IF�:���qc�Z?f]k2�x��8.�wi��1����"u�Ǘ���ޫд��(-ً#�mbv�VǼ�j��tU�����3�He��}wO����b|�k�wl6���n�]��+ܺ;ځ��{��N��4�!����Q�)I�t�u�aZr�� �f���͆��}�Z�fs�ݞu���l+N�^���Д�Z�{&�C[B�M]ԞGS�ve[m9�Om�T�,n�z�.�2��\u��!�R�T:[@á�se��s(��rӎ�J7��P8}ږ�йcBg:� +�˼D>:)�9��Ŧ�gw:�8���F%��Y�\1�@�Mg}[�ĳG1�f��䳢�,�c�Z�νz�O{9��eɱ�` XX��<p�=����`ga��x�C9�O/���d*��v�]�05��T�_a�T��4:��2Y�Qg9G맘�ģ�ـ�|�e4!$]E��,��C��>̱e�A<2u!O�X�\'�5�X��V>R�	�m'�u�K�Ցm��A�����)*ؔ��7p��ϫ���p}��Ww �IMTԆ�p7pf�������Wx�	�/3!M#q=wڒ�	��;��<h�v��sMmv2
NjT����3������$��� �\i�4%^R�]�k4B^�73g7e�kE��K����oE{&G�+53P��;{4�F�T�"-ݧ�o^�2�<��1�:�*ދ1ܖ��R�#����[�>⊼���]#���>�m��5���M>Q��m+����6�:�ַ�)'��T+�,��}Kmop�6	 S�O��\��W����uNs`D.�����D�lh���yi��nsۥ3(����Q�0pSpcU��IJ�Q%�|�8{7�q�(+c���՗��&����LS����_?U�Q��_*Ŋ��\�e��|%�@��f����q�X̾o_9Ӕ���l!�2A���%SK wv ���n�b�(d��5es� ������RFP�B�w]B]�FH.q�9�[-	Z5�h�m2E�"5E��$��f�l3Hh�����i�PA�H��I3Q�b"��,��kF�܍��p0T�d���j4`Ů[�Q��h�5�˗(����Y�*6I#�r�	6*$R�����cb�eJh1�TRD�FX�A��,VM�p-3%�$��m�t\�wvM��чw6��"�tź] �I�g.ۤ�,8�;�����u77';�,h(�m��)Ia5K$�"	�7.̙���{�?�����5%Y�h� ���%謱���2��*��n��O{[��aۅ��8�"9E̪'+�Q�n@��)e�������gsz&�������7����c���0�U�~tOv>;2V����C{�͗�n1����t��p��q��dF���x�]�c��ӭ�N)��RI����gNTO!أ>�\+�󋂞�n�z9�V5��V��4��74�*Qt�����������������Nt�ϗNy]~��-9��e=���.hO;�U�pX:�|TrQ��DaQ?_ ��\�&P�m�F6��2{��Z��uB��S�v����Q2�_ԥ�h�K��=rX���yz�P�=;��ۅ8ݍ�� �:%���3�vi[-h��� ���˃�����|3k�r�N����}��'N��uog�xݷ^�߯�>e9EwpX�r��uJi9.���' ��l��؟=�}y���m!�>YT9��Ы�Vkx�`m�Yy����0꾃�P:�yʒ��[R���9ۏ�Bw�ղ�2W��v��.�\�yF�����u�PM���;+��ɹ�v����5VJ}�-b	I�OAX��<��S��"�j 9ݧ�qh�L�.3Y��Ix�m� �����7��I��t`��$ߺC��F���J�ˀ��}�W�s-��ƍ��͞-uN�O�Z��0N��P㕡P����'J�%��bɌ�Vp�&�sՖ�Zk�p�n y(���n&��nj:�W�nJ�x����0��1�ӳ����mﾎuyq���Zp�ns6����@�@���#3��T�K�l�KbO�����_d�U����6��nv������Q�F����Y��%w.	O����}R�eF'Y:�:e`��|�#\�׏rD�^��[�@�Io/��	c1���y���*'��Pc��3�.
z�k�t+�D42�
�8�g)ƽU��v㹖��U���]^��R��w��h��yßS�˙=��m�}.�[�o�vhn��P/����ҙj��9	���VٻMm���o�_>���5������ו�~�'h�Z�<�sXm���'勄ˮ2�ut
��3���>4��(�̚���������O�fS�3�Mw���q�r����=N��'C���Z.3�� ���ٽe�f�0����|�!�ȴAKOR���{����`49Z�g����=�7�l�_���wK1v3��w������j�Kwxᬷ�mCi���9X�*� �/*&K��<tq^�(˙�p9]D��K�t�Lt�|�OC���n[�}UyT�D�r�U+e@Ï��T�w��ilI�\��)]Я�{�T��H��&�����ߗܦi��H��nَ��p��Nƙ�f�@K��Ih��X���p�;N��$���
g�=�~���Y,X����T�9e.����&\ri[/��gV�D�lҙs_q�I�Z�h��Ț+r�.	!r\f��⫗Q�I0�7�!�l\Ls�5C����M)�}�I)w��B�K���s�&����v���N��k�g)���g���7�2X��G6S����.��Y���|]j��{�s�i�9��k/9�<zl��O�W\�V�p�M@���f*�xV��sYZ��G��Ϩ�Xh��D�5
�h�Sx��-�Y�ة�aS:WnJ�E���!�N������%=��՛��x���7'��Ի��*h!MX��'�`֣���ݱZؒ�"��d���\�x�C��ةw`��J��O��H�Uf�*�}w-s���ѻ���?�S���OW�b.�������:����*��u���ǫ�T�&�Ùn,��k��8�̥ⱞ����U�ۇ��WdEhoF��ǾT{�/S^���qe4�>�y���5��V;����Pz�B3f9,�K˗�/W��Y+*�ss-=R����Q	���P�H-�ժ+P�8N�:�+�Tr�ݱ��_G7=o�%��x���b�'ewj�7 ���N�`�*�JU%�R�bO/\5�@��"�F�K�Dn��$���k�m��)/�I�?�1�Ry;��ө�%�)ר]�ϧ^#`�nֻ�x�S�J�<.�ܦl%7�N%�r�M>��[�{�Ob@ap��I@y�[��t�~7U���tB�q�����j�.� vrҰ�c�C��i\�;�fد�{Ӝ�2�����A2zP�ċ�wW�Tߎ��An�����+z���Î@�f�\���1<O�U�Va��>�&�)ރzy�i���E懣k����6�טy�7j�J�"u�([�ڜ�ȇl;�v��l,[��+��������3p3AV�5�ʍo��D��@�#u�KܜOc;����6�;ƻF�e�t>(�r�s�~b�����8Gs��ۉ��Y/>��D��Z�H	l7Y����S���=X��)�7P�ȕM��O���e�J�5�2=<�׌�үЦ���G�� ���#_[P5�z�����jꁘ�%�����o4���֛w]{�(�t�Uj��9__J�}�C�_dZ�;-�J�]�o�� /)E��[�r�܈��+V816��vg+=ޞ4��q?E���X���p@�N-ݒ
]��B��j�np���D]/fzz���缜�R
W��Q��9�N��̧O��n��w�=�*V8��b��O�Ӝ�<r��W�-U���GBM��W[�9�6Z>�JWGCܬ�ͭ@Ӝ��XK��oP�QT�7���E���\��F��]#%�%��o���i�G�T��=��ˠ�&���d��h��X�ãמ�^a~U�y�x�i�k(2)P7M�M����y�tx ���`p��YЃ1}H�����ul\G0l�y+�+b�to�ƴn��e=��������;W`nu�K�Lw\fg.R�ĸ��&����\k��ޅ��i�n�m�P�'`�� 1��7T�o����{����ܜ�u�I��ƻלoa:n��u�/�,k�����q�5�K��pvN�r��oq�{��9����.f���W˳1v�2���g�E|5k�f#�B��Wky�`�Ktġ�ֽ���t`u����H��{� F���MD�̸	�E��P�2hV�R��fnmYo{��*�\5��+�n%;b�۞v��\�ɬY=G�Q6�y}��x���y**�&ާF�m0i���Y^�j{}��o�=?�j�9m �/�W;�n̸ד�V���E��n�6�\w���KC$�##����{���9$��K̨�Ƿ�&+*�qy؜3Qn�ۆ�y��N�KH�ޚ�.0�գ�r�b���t39��j`Ǔ���ī��q�Y�]r���N�G�(�cEX�\�88�-g�:�K��Y�#���u.���o~k{%dQ��%�[�O�4���e��u|m�A�œ�G��j뿦[�J��N��TO|�B�L��׬�T7z$z�_1���f[ef���n�[�ޒ��v�c�Mq�U���}�	۽�|V#��f��K��-�닩v>v�y�!Og�8t��kGc"����x�_�����k���rÃ�/���X��+ĳjL#�������ɇRq��y��z�1�����us�:�$���dr�S��̸Rr
}/k����������Q	��<�3�s7czl}��yGoH�J���)_�[�pը��mCi��W��)
�ɶ%Uj�{������UY�"���D��t�OO7|᭷��<�w3SUPꧯ8^f��d��_?����`4�O-�vv�뀱���[�6`�ݕ̓r@�}��R�'%���S4��F��al�f����T�W�V5�p����9���v��9��2W���Ϧ���8��tNet�w8�p�t�i����e�w�8�b��k�2��W�kgt�^V��f+�+���kr��5��\�d�8�RYZ��ՌJ�:�u
�i;�R�0���fn��$`e��HQ�A�+�=s^۵�H��n�\mcڴ9�arbCm���w�_n�x�j
��N�Q�	�_�2�"';*�P����%(�� ,�s��Y�;�߹u�$Æ�B7ظ�Nj���K�]J��+�B�O�w2���kOk�q	*���mƻ�g4��WwNB>����UΜ�a k�����q�Jf53�u�';��}������ܦ'��p)ɸNu�fr#\�}�3D�ʕ�3���#���[Z��۩q��2���o���/@̣�şM�TOxf��3:�J�5����>m��3�. ��ۗ���j�X���?�:�=�Լ�M�!����=�qظgK�4�"]淝o�vhn�E-�Jr�6��Y����qRw_�gdJ��/�(����E4��_>�+:Q��fرh&]뽐�9рnS�� 򯤾�Qʣv9��sw������vU������8��t��wl��v��"!�QJQ�Ğ'<O�p�hkݽm=�y��S�,�� �:�?e�򂾵��e:��IyPۚ�����=�S�x����".�=¦`t�b����hV��n6�e�L5m�Q���W�ˑ�z�`Em7^6���/'u�g>|���[IQ=���+��0mK��qT*��kjr�s����ܶ��~*�<�	ؓC�M��JW%3tL�p�O��f���2��x]/�I�0����qtаqqԃ��EUԸ�k�-+5�y��3�.��S%W���B�v�F�Bs�8��u"*'<�\@]١$��-	�6�Cob�͹i?�%W������<�ny���%�f�>V�����*��2����][����n.�k��j� u엢�+��Z��7Sز^f�V��1u�'��qݺ��M�����7�#�9Z)��Sٕ��+��;�ӆ�69u���A�'-r�q��5�l�F�ʭp:`j������n���~}M��_��uf��S��i���3����׎v�����2��]�K�\��⳽Ld$����Y���X�ͽ\J����z��k���y9�u��j6�V.}܂�$��=o�+�8���F���Y�Z`m��m��`�zV���h�K��͞C��EV����t{j���8�kN��ݺf���/%ь��1�
-/��	t�-����˖��+7F��x:�gu���1�޷)�����$2��rz��_���k|����\+��=�o7�[��6�3�캠8Զ]�¶�܃�Q��P���F(��\�2j9�H��V��D�;��^6�Tc[=u�t�]?@:�$��Qʣ�@��͝�Ii��3*&a��M�~�ϗ��9l�sW(Lzu�#%n�*J��Y������5yR�/9<��e�ж�Oo�8ݍ�� ����������|�Yw�+h1ە����,5�I�;k^��8�r���	5���b\��ұ���pv�!�4Lm�5
Wu�X�r��6��q{�ڵ���Ua�j^);Q�5��J$j�0�b;4*�iXy�՞3�a�ɥ��`Ԑp>�_%qBLϹ	�V�=ɩ��=����qU����mN��r�f��x	���
���q)�Ӝ�F��Z��K��;y}{�f��Z�����9��&o-h�KI��9H�l��"k���LP��lJ�����|9ǳ{Q�yOn�X�F�wt�WU�*��M�����#��a;���u>m;�hM�2B���)��M�Y�;�����w0U��Ѱ��]�9ƙU��x��pHt<%���67�-<��y�f��	W������_:��}���#������I��k9���-f��t�,E��&����^�y]��j���,��,���-�0��4����z-A����K����F�7�;>��V���KnI���Ǻ-�@���hG[�F�[b����S����j����D�(��|�gçiz8�V�eO��yYE/��J���y;J9O����5u�B��q��2�lc��w(4<���7�Y�����\�h���U�P�.�t�U�"K�I�/i�[����f�
�DKS�J�L�z,͗v"�݃�������sVm�Mk/$��!��u�V�}d�Pu&�eX���"EX�I6J�)-�����E���xq<� �j�f��{{+%58^d����2R��K-�ݭ	�U�n��C�n��yw��㵬�W��fjFZL�;���5��]�7{���(;�Wl�㉨��T��zj*ݻ2ƨ�W/�lm�}�:��:L�"����E���~�kSP����ѡL��2���&$@sr֛b�,�u�T3R�K �afیh�x�'�N>7s�
�N��u��}]K����:��c�_�k���`�_.�(�oXf�Yy�s���w)t�u�lMb���e]��bL��"@k��v�q��=�[v��e��[i��y%�l
I6���zl|�Z�]m\ccP�W���oe�1t�֋�3����!�V�ǻB���B5����Sn���5���1� �͓��i_e֮�Q��J[���l�(2�+��V$����FѸ��Yg"0���U�Ozd���"�5V0�W`흡�t=Q�9#�,\õ&]$n��2���z����,ݝz���`ì�L�b[�)H�x�qO��훵�q�L󼑮tM�@|z��Z�S$�Jtn��U�z�6����r�9�0= �KC��w;7�mv��j�oR]1K��y��&]^&�	-K`k847'���Ss�m�7��W���u#'`�~�+�H]w�vE���prG㳅�0�F�q饯���Ϡq��C*뒬��nZ7{{%]�u��u,%���c�͑��q���p�O�	�PL�G�+��D�* �}Có��6�Vhάե ]/q��Ы�Kǽz\�*��GV�k���I��}p����-U��y*�(NSÒ�]2�
ݑVb�NFQ��Ǯ.��(��uY�ڳҲ}l�9�o �Hj��b��{�ڈ��֩ԩG�R|�4��3xZl��C���Sg	[+9�f��E��Zh��4#w��6�q�R�&Zٻ �|*ɪ( )!.\Ɉ��6D�[���VB
4F4F�"�r�����L�Y5%I��lW+�l�!�PY9E����ܮR&7wF������q�2���\���I+;�uݹc�ͻK7uĉ'v���.q5˘�!�dL��Y���.ni#  L��#b�H��cc,��Q�rN뉓��41D7�s�RD�9r�2F]ےFli��4كF��Ak��"e&+���2#M��,��I3Wu��1�$�!��d��d�e!�v ��P1�w(R2�Db)4�Kb$�`���￿9�B�|�N�7mm�ޔ9�gVR�f�ڜX���pb�K�<��8"��z�Ώ�3hY2��,=���rɻ��T�*\�6��|�`�n5�#q1���>ͩ��l�c�I{s�{<�����r�핗/;'���9��N��p6����em?`0.ڵ1x+��g@�|��G�$%� >G��%��W��k���N���:��88h�!9���ޣҰEeO=P2`Zꁘ;�X2���\J��I�˭1�+��(�Vu�F���ʮm�<�f��U���'�������Կw���(�n9\�l䒲Y�U�կ\������*˥嶺�6�}�x�V���t��3	��c��4�%�m�7�������Q\�:�n:Dde�V\��֧J�/\�=��]QL_ ��ͧ�����P��w�u����T.�b�o-'u�.��/�\�)JW���Z��[M���-�t����V@y�*`��z��~�D��Os��V8�|����j-�w*�CO�x�����FK:Y�9�i��*>�-���!���⻫���N_]!��)\������K΋���gv	��9/��R��VXh��ަ�o>�����,^�d!LYrk��ۉ�,\r���+�	!NCx��l4�f>��]ї�z�nQ�SvK�I��s�|�@�
@�廇%�Đ�}S�]��r�]#I�t��&4���M�[����[ru&S��SS �8Rҿ��i������s_)���.���Ϧ�"e��@�I�ղ�CB7k�١�%�\2�6-���L7l�B�s\B�L�R�W�rA���*%��d��ɬnc;����k��q������"��&���j�i-l��3j�{���Mb��m.�V�3_6�X+z�Pȼ����w�WY![��Ș�����j�%�W�+�l���r껼�m.��PC��H'#���t�;Q5_k��o�b��xVϳ��ߩ�\.w:M7ª�+��WC�������Oy����b�ƍ錹�6�U��z��'z����Ÿ�$���̝F�y�������V3�a�C�l�,���1�c3��ƞ;w�]�v��l�B��u[y1��̺g�a:A"���FŘimf=�rTa�O;y��N�8���<��Z�7�w8�GV�5"�}��$��MrzHr��u��a�N��[�St�����e��t���3���U�%;�鱠��.YQ*b���Ë�SO��w�p��5����hh�S}铖OV�l�~��V;j\�J��_E�ﯗ79M>��ϔ�<�Nf����ֲor�2���u�t���g髪v��]���lG��=��F<�������A��F]��w��|S�������qN���mC[p�-y�9�7p6ʥ�)�;wik�qe���3sP��v���t���We�ֻ�x�WΩ+��_r�쉦��R瑦����o��������-+5�7�*3�.�D���*7�Xx����"���\���=]N�{�W�o��fبm�nu�2�Mرnw3���L^����ЦG���z���*�
����o��Ḙ;.�.ki޸��֍���9��6n
ܒ��b��5�94�i�=��F�)�;����Xf�/,��L�.�:�~�ɯl����> l_mk��,Ov�;���ܰ92��tW)�S�eب�ƲN���DƖ�Nܥ��l�ˮ�����z]��g.�v�	nN�i��y�;�c�zed��כx�vM�z\CZ��Mƻ�V_��6�Og�R�tz��=�E��Iġ�m%|���s}+ֵ	~��͝�S�jځ��V�ʨ�p:`j��k�@�z����Ҟ�̗̈˧����+(��R�T�^�W��Wx�%��/=�I|��hV����F?�ͩ���]�؉���e`���=e���Ŷf�ؠ��Q*t0���}ic��48�ۇ�w�Tb��b�]/�YO_Bɬ{-��,�J=Jjz��{]F5�Ҭ�؃wz���C��#ή���O�ҭ3�a�s��2z˖�ڧ�p�*����:J�uT��G,1Fə����\�F�pQIR�o�Z}p�9o\���8lT��N�+��ر��km���]뙴�Y���k��Cж�OmN7p6ʨ\�8�`f��q<���ɵ���E����s�t�qa�)<�mj|3i�����z�Zpf�6�%�E��6]�ֲ[�����x�M,�Aat�����v����ί0S=��H!Ʈ�5�Y�6;��>,��e�%,8���9��جq^.�3���.{��&
B/;b�;�B�i�'wh�P����t�_]c��g��)��~��L�h,��niJ�o����9=�pA'�))
ż�t`7�oS�#��P�"JT6o��q;����t%�~��I��=����3�k�so!�r�S%WH]P#HO��M̱=��Ӣ�rg]5v�=��L���m�h<a�Q��
m�}�.��9�9�+�PKn���Sz���U�Ǯ.�I&|ۍw�K�q1����1ǹ�@��r{�������;-nL�NeWs���8e�9�O�F�wo8���kp�G�b��y�f�]��^�m��x���{x�3nY̒�ZZ��U�j_]�}O��k�V�����������կ�rS ��oK�Z�k�t�bS'�}^�p����iªy��K�aŵ��5udmP���GE���kk�L�&��7���L�~^ӏ�����!�<����kTBkug�[�T��SޒM�>L�;��=�,�G��N՝R�^+�E�/o%Ƕ��r�4����z�s�N�ŋ1v�A��l��\¦���W��soY섞��hnT�&� �.�8&�Uz��׻Xr�]J�(�סP��ٻ|���~��V�X�s����dK���tc[=qV;����:[[�D��e�����I�_K��Wo�M���i�|��Τ��ͧs���-s�kk_E(��p�p2;�����Taj�1Byp�-m<�"��h]pz���pۈe�����|�K"Os�C":y���l؇T�@�L�o&I%�Ӕ�7ªܤ�	D�i�g�����+�Y�v��x�l��.�u�8�n��8�֟��������^c��f�j֡E���jZWkY�9��gi�9��L�Q�T|#b���9[��� vl��Yawf��	sW������3��\У��n�F��]�\g"w��v���ygq��s.Dÿ�q��F��b$f���eڡ z�e�;�eħ�X�c�㴕M}i�<h1�r�0&6�W@�JL�A��!Yug�w�	�j�旾�Մ�K!IN:}�������V�j5x��%��;g����iN/&VmgrSU��P�f�u�ؕ�����;'Gyr�	U;��G�� 0�d�1ѾO��8�sv�b"V�D��58�+i��sfį|��B�>�`�@����E�o1Z��B�r�>Jx��{��`��ۆ^K���jk\�{�1TM�+�V3��l�ڼ�MPT��l�{�N9������\���A�O�1U�����jܵ�WQ�e������g�\�����ϵ�V;��ON���,�i�+{�r�$tr�79Q�����p��|��i�}>)��Q���X�T5~֛�]X��EX�E܃���T�]���Q7˛���|u�ͺ��4>����Ae���5?\�7�}�J���<>d���d|�8�ghfӝ3+-����)�V6ʥ�r;D{���J�b�ǯ1��B�5E�6���m�ж��-f��eR��ub@Ϋj��]&Uد2O���~���I���冡J�Z�c�P�uI_��u���l���@�}�-?^�ݴ�8�!����O;�e	����9�#�{�I�27��s�A��Y-���mp%ϸ|�)�j����u����J��mF��/r��TU�32U�(`X�e�}�V��(fx��ʴ�K��r*��{.��B�FVs'/1v�d�{�J&�Sp�c�nZVk܆�E|�t�Qz;�U1]Oq�<]8��>�3cWt�f�P�J�7��Lf͸h�]��$߲L]����?�\�ЏK��~V���������+-�������<⨎ѮQ��f�:c"ۚ�F���5)��,3p�Ya�T1+�v��QtA�m:�����k@�|�dO;r�Sꁶ�{1	�b�{�bn:*/+Ϫ�<�{3��&�w�=��6��nr�5�UF�05r;P�ШG�8��M	���R�ecsYV�����^2��юv�N�nܨ˾ۮar��L�#3��1�yZ�ՇϝL�V{�<i�<�Pƨ�^����IN���O|��G���P㖹9������£�󊖅�b��2�uI �D��?���{Սl��·(� \�^R�W����ǛX11*朗g��K4��g)���� zs��:��;�t�74�8�|�[;(���ѩ�M��:ݬ�Y����y�f��F�+H�B�3�C��9���8ޗ�9�����M�y�*�Ҏ��I���;*�sN�ҙ�Go�]&���8����s�ĭH�98�sZ��mb�kg�����UI|%����S=G{���p��\�Ҷ�
��A9��nb�zq���\�mKu�}��xu�[a,��;zE"V����+q�ǡg|�{jq��*L)�u՝�$�������0Dw=���w���|3jpVs���op#\�W~y�HO����RvJ&�4Lm�(��iڧKH9`��Os����#����r]D/�T+jO�o�L�vh�;�R�wy���U��l<|����iKS%WH]P#LP�Et���Z�Y�T<�������X:[L�7������<a���Jv�4�#�]P6�Ln��=pUS��u�͗+2kLf��9u���q�Ѹ|*/�v�X�U!�d��s+�.a���̸�[ɬY1�V���SQi�5�_s��t���|j��;�i^����u�?$s22����;�8cvՊ���H�����śN	7��+&�<i���q9|�dS>����n��R��_l��ևH�>��:��c�9+%�Wwԑڵ��jݬbG	�F�Ǝ̹�aڷ@����V���`@*�`�oj�/mg%����>Y�O�<�.�{�s�ޝ�k�}Z7x��/��R�9Q����]�j	�����;@V��|�a8ha~5{}l�G�����E��K��R�%�ӏ3z�q>��o"���r������eٌ9�+K|��^���ڍ��#�
�;���TZǛt�+�b.y�e��y�z���7�v,wj�:ME\L�y������������W0�k���B,o�y���w�wC6�n�������8JQ;�����0���QR}�`lI/�]1��2T?P��_�8V\Ϭ�C� ��`?)9��~|x��H�Ĩ�6�O��%W�a�
�2*e#uS��EԄ=_a}W�p�g-�1�J�J��nUe����_��0�.�b�덵,�y#DI~C�#=Ɣϣ�خ�
�yz�6X��@'U��;rB��������#�n#ڪF���~�Ӳ[ ������EE�A�Oz���c֥6���1/���˜g�q�8v��SI��7�B|n���:~���JL	����T���XgEe����Dm[冏!j����,4��qg�;q's����?.�Ͷ��_K���.tc446y�&q�A(�"e��{����oK�7�к�+p�J뀅����-gr��w8��5d����a�4�v�m�t�H���%9�W��\�\�$+���jl<850T:�v�5܅�4Mt~�����}Y�TX뻋�B��3s>U��d�E��Eg��z�(�-�O&	9J��ۉ�%F��ma�{��E�g�L %f�ôm���a�r�)ut���	�P�"����ut�@
lv��V��dum�3�Ƒ�����뱢��S�(�ԫ+$[�*��m{.���Z�ܧ���\��7C\�d1����)r�5WsV݆�J^�ob՗-�78S�}��:�Zgr<v��)l�q��M�^S���lgC�oem�a���#l�6��U�QoR�M�S'k�ս����VYA�ص�\��dчl;�&;��e�v^.����\��M�:���*#G��MrPd����-�խ&�1'ܻ�1����u���6�$1m5�V❶��C[��*f�	rwZu��Qi��R�]�ए_c�!����C^���|͚�n�:�,VvU��vکf�X.gm��.�Eڗ}�/��[�7Fu��q��Ȯ�5�4��Y���p��[�]�#�Z���[�L�f�����;W���NF��Mj���`� IB�iIO��K���Mqin�Fz�>�Ȓ#X����UoJ������a��%�
��F.������2��ۉ;�`�V�<����R՝@�ʩ��!6'8^1�쾚��S[��y�P�>�1u�+J�S� �Z���ueeol�N�� �+��GSi��b���l'Q��nr0�H>��b��zR�=?��&��w+Vu�GI�)�z�2�jP��H���"e���r�>Rw��5c���}bU��k�V՚�Й�Z'�V���[d���h����w�eY
2И"Uw׶s,��T�3t:�U���g����l���m%i��)�P���9]�Y��0��:��ٱZ�d��&VZQV��L)J��N.˧�B0�Y�tIoz�ྐྵ�����������Ku��t��zCΤ2�	]+�������G"C ���G�N�^��R�fvQ	�x����:)�1���+�>cx2l\���B��Ǯ��b1�W$�x�w	Z�A�dI6�r]y�kf#q�6:A�CRe4�ur��J�JƫF&N���.�{]�g�1��O,�� �(��G7�S[�h*�PR�}9Y�]L��b�T�����O��Օ�Ǧ��!O� è*�+�	!��:�l�U�����
�X�&�W�ec|�����X�*��<�T�+5'ע��n���������6�cg�]"K.u3h��EL�k��\wY4$h�]�(ؐf����k�I�͓$k��r��(�;�S��H���H�w:�J���黮���b"��bƙ���IRr�D!$S��%�dmsvnr���B(��(,X��Bwd���d�
R�F����ٚ�76�L�]�b�#b1��������wtآ����.m�sc��1��s���k��F˜�NF�
6F��nk$[��n���.j�Wwt���t7\�;�M�rH4nnFc�������9�p��J��zh��)�	X55.�.;8]�8Wiۧ��C�]w�� �/r��F��}��������ຝ�����F���f�~�W�ޞ��븋/6�s9��n��:�eErJYRHj�R�W�*�uNu�{��uC�_������T-�!�ͫ�c#��gœl��e�4%����;���i��y�7� �ul�	_�hD�>�F赳W�Ǫ#R�\&��[n�O���w������S�k�w��� ~�%[�:�2��{Ǝ��r��3k؇aC��_s��J��6�Ǆz�2���Ԡ�8�Sθ+�3C/�!���ʰl>6vp;�V���OqzNOzQ��e���ػ�yY���&�����6��yI����o����Q|:0�ss��HtL�Mc����fɢ��(VV���J�"��ay�N'߿*���L��`��}3�=���v�ܙ����L'ИS�r'�&�%�J��:/�%���|ܦw����yKM{/��8.�e�^6�P!ܜ�d<���(]d֛����{L	�Z�.yz�X�O��W�nz�6�uca�������TA~�7�i3b���A���:\ό��C�X�@V'Kޚ��2�r=�+�MU�9ڃ �G6���g1�6���8��3/C��8�C�*���&�݈�s��d�0f*�Zr�n!��N5��ҏ�c*gwkc�[��ǘ��.��v��<"��-�uv���?-�*�̑��o!���� T����JI�|�g��_��ȟm�p���,��Q%��ѣ*��Q�#qE�L�F̠��|�؎��5���w�݉�P��3�oh6�>�:�Y�:�A�ç$�r�%TD�#�C�L�H���%c��.����])���S�c\�=��{'����V2�6pK. 	�A� �XJp)g�R�Qw�+]A�rS<�خ�49uz2=��i��8v��Br�Uqb)gս>㏭jO8�����z�N��6��� �
��]�W�W��[-���e�Ӎ�[��hNƽ�zo�];��`��J�5� yA���AO�	�����7�la���_]��tw���`ԑ�Or�Mz�|�j}��߉�2{SF��8�G3�=�/]�c�hӿn޻ʸ%�K{��놜Dk�*�ÝӃC���W�K�όX-z[�kߋ����y�~Ʀ�-�Q�P��oZ��R4/�̙<��c��[��1�y���lԸ��PО��K�%�uy�s|";0�0��C'�}��x=�U�^s	ɯ��;_7J1�M��`�ZƬM(��%Cɉ���D�s0Q�F��U�x�c�I�� �T���_�J�VW����^��Y~��K�t��kh͋�.#,U�<6����q��K;��8�k��]�m�Z�)����y��Ĵ����B��־��<�����79��s(��.�*��H�����V�Γ����ʫ��z^P�sQ�o�g���Aie��V3�rrʹO��WMx�v���@N�_�Y^�S�vXk=��|���-ϻ��Sb�������Z�f|����"��R��kd�ِ죞C�ZXhQ~%\m0�j��[/}��G�W�-z��/��Ӎ�N7�c���ע���QT�$��9��Y�W���.����R}�+�7nn�wt��>��=ޤ��E:��dC�\og�{�o���$��aP���|�4z�rS���:_���|�c��}p�Eo#��a�l����f��Ҵ�4�<ꩢcoFq�>ѹ˼������-z))�t�3;���F���I���}A��:V2"
�Y��X={�H�����������&(��
e����/�oף>^��+cʎ�^��<yyf�K�v�7ճ1Q(�����F�k�� ��C��f��ö�GSX��3��R�b��߽6�����}��Ꙙ����[K�3�:��U�)sC�D>�Li��r�����#�˱nB��)lQg��#DTCR �����#�=��#-�x��թ�u��`v���f���~�*�9nfb�/����"�Jz<۾0�wV�Cx��|H���� ���mP���>*\4�nd��Ӗ+u��t�]���L��B�l��{7fog2����:4�~��λ�3z[<��5�m��9�eg$��j��7� t��B�������ipV����j0Fx���wz����,�.q���[&:jZ9��Lw�~⧱�|s��"��gl�-�«%�Y�Lu}��T�@ws�&�r�k�8�a�M�2b�KY����[�=Im�h��"v�B_��,'/
��ўԪ:=撎���s4�v/Dy��^��彿V��p�/���!�#'�"�=��GPMf���F���+*����ziL{�xX���ۋ�cb\(�sÌ�4:v[3��-E������bJ��a:t?�������"]W�=QUD���%�M��y�֓����o"�;X�_�؝;L�(��ԭ,;sqLLp=2�w��,��Փ��b'��C���3by�f۴3o�X��^)ؾ�S�I���EXE� |��ۨ���n�z�Q�,����G�gP��u�Dk��;����#��ix�`ӇbC�B{,�ʍ��P��+?�P�Ґ��2��L~�7�@:�t:p���3��5�~�]��SH>U����w~����'i��()ւ�gӶa�QO�m���Uv2t�-&Kܫ�,��9�+Υ��3B��$ʝi�=���'�e{�bC��LQ�'Iݛ��Ӱ)�$�$T�n�؆GrU�ȵ�&�"�8���y�\��Nh�yu�
��N&L������'[�ʳ	1�^����JCm��{>�����׃#\K���k�v_N�n��3#�e�!��zm�^��jx�y|dh�~�����L��s�yPL*��#�m��c�{�9¶��_t���Q���yLe}ΩǲN�w9 '5x	�7P+��lχ�Ÿ�����;&��`���K�;E{�	c�.�x�=8ϴ�rp�<u1�*��iD�\x�ҝ�������QW�x�J�@n�;�P�Of΅�^��doS����Bs~N�����6�{f"��e���Y�/ ��;\Жu��>
�fю���N:~E�g<�E����"#J�WFj����MA��%�R���4"{�^�tZ٭,{�+�������K%����d�M�����P�
^f� ��.D'��6���GT�D���ag�v�yN0dp�cɎ5|����{�4I~E�j#�_s���Qt�B�Vf|!GiÓq��,�=�����)��4���M�}GyR��V��D95�yI���Q�#�5Z�A�.=����&~��mZ��ͷYV�2�lᵸ��rC���w}w�"-r�R�b"40����"�p���~	gKۗJ&�}�cV�Ф�h橜ybvu�N�K�NÝխ�yw���Aa��i�R�0×Ջ�)J�Tb�M^�u}��5m�Y����w]��� 퍵�r��g�^d��3?ǒ�X����ay�s.'|?~����S;ߤ���5��##�%׈�{��Q>#��w9GD�D�}Y��cRy%����r��`�^�*uU��[�f������+���,c���fGZ9��J�a����V�@��W��s���]vm|9�܍�Ą���u�G{���������pf�=P�T��]��c] �Q���s\f2���;�.�K��S�Y�z��Y/m���Ad\�J5%�FUC�3�d8	�֖�]s��'w>
1�;�ҡۘ����{��'�Y^����.�����y���J�y�k�R�u��/��y1�*r��H�3�kw�9ޑ���d��y���e�5�G�O��ɯH�5=�7������K��$�{���h��;CFB}�h��W��\NWΪ���݈������}u}�b-�/ ����� ��
���)��[���<�WE��N7[��+�������9��{<�މ�讽��I�g~�D* �2.$�>pa��oa\7�l�n2�kC���\=/A�����<^�+�aycc�i!i�.;�&�A�*���.Е͚��2�_\���:ʍ���'ϭ���ɫ]����Z����5y�kd��}�/	��h�b6鶦�z�r�=�fr����Ptu�l�+�U�8��Z�ߡ3�x�'>m�����aWÒMM}�$��|Li��jto�/����??hp7AQ�h��[�J%%����=�;�4�#]�WΓ���~j�'�\yXk��5vzV�3����5 ��{�����v���q���6�Q�Qu��8a5p�M�R��竡o�����4��hH�P^�ztOl�\2{
�����uZE�0��g��jb���7���ӝ���ɮ2!��c캿�N~�j���v��\�U~L��p����>����sQ�o�g��#y�U�!�Y��j�����)Y��`��Gy��:�+�o�s�������c�U;�O�5h��d�L�^�X�Z�D3!oNk��^(��c�݊�9�ƫV�G�j� �]�=~�m����p_yw�M�7���bZq����F�y�z(c���r�<&��o��/�q�}�����~��Q�m�������u�\�/�u	�ϝ:��/��}9�迫�I�g��ka�:N{L��ߪc�jf܊Nc��g�B�u-n[>����ҳƻei�e�{�:/�A	@�5^��ܥF	�KdP�د�q<���o��D�H�l±V�l��{���p��
J<ŀ�]��5
����Xuh`�yM�Y��wx�Nf��3[��Aΰ�<�G>j󘹐[�T���M�x�z�d�=�C�����3� I�M\��IS8�� �|e��ʗH_�RӚfC����dkz-�m��^��t2z��*7��wf�zl�{����D��X)(�[72��}m��V�#���#/�+ʵ�ra�)�ձ8hyӠ���:8��r ��r�@����vZ�	����T^߇ֲ��W#���A{^Gp6�4��f1��iK���cL�n�P�|}X��S���V��ˮ�ç�b��p���w.sKg��-���J�U�)=����1�[���Z�л*�w�y@��Rw���\j��94ܿ͂�/�j#9�d�=i��~��78D��s�t�,��DV*zu�O��=�f�1�=ު�+��-�#�,L_D���ܭI�Lq�}S�}�a+�b��oF}N}������,{ΩE�s;��"�xy�w���kl�{S����C�1Cz���Dv�vGjk0�G�����!
ʺ�h�M̓Z����1PK�-����j��͆�Fם娻֠�B�񣘇PV��#�N�:��'�w-l٦7��.nI�zv���P7��?#�_�)MH�XhU��Qp�k$��$�]È͎��+o]T	V^�6�D[-�5���+��f�ჶ������ɂ��+�+w���*s�]N��X��ي]���R��5�cs�HV��믭\x�����'$���/��]N-��	�ܜy�֓��<�߶ݗ���Pͤ�i���W�\�~��)�f4j{�w��^����{;�>�:�G}<ֳm��6�qv�#��N�\�L�<�C�q�/c�&\:S��P�!)�>P�p+��x�ϥ�ߊ��\o`n��}���N�\�ǝ75޸S\]']����S>F✆U���u Za�	��3��S+�}�x��Eu�{�\�������3C�=�1�k�2����R7U>	��RW���l�1tq�6@�1w{�2 :�o�{@7]M�ă��,�2�,��a�Q�����}�n�Q���c�3RN0[N���};o��q������~χN�v� ���x	��s��4�m��������Q�-��vP����g���nN����5)���>. E���Wr}��5s6KLEj��#��V�X�븋 ��|p9��i�BvZL�MQ��&�)���ne%� �4}�$wA��SB��x�������Cޟ+>9���'u�{��
'XKr��ha�F��`+\KU����z��mk�QG&��l8Ƚ����A��3��u\;�t*�T�:k�@�K3�T�ޙ����Byu���s�<��YҌ�1�*4��p�5Ƿ��/�{���m�tI�#Sn*��2�Q"(Ń�9�I����Y3����^m�92��#��M�}^�!���ǔjW!�M]�����4�}4��yupHƽ'X�>�޶h\B�.�!�tѯ'Ȏ���պr���ه��cFoY��GP���sv�¨������Qhw��q�C3C/�!�zḽ���aϧ0��¹���j��w	_y�>��(
ʺc�{���sQM<��m�J6�Yid��<e_���B�g���%������蘗��&�2����<�b�;G���w1:�i8�_�����i�f��=���kz��;��,��,:::NI�ϓ�'+'���ѣ�{�E�:�l7)���v�'|��U������~\G�ח?�~����1���8gNӐ<�i� {:�+��؉�u���f���::���8�j�4���c�K���pf3�}2�Ӑ��
�c����u���I��|�)��E�������^���렲.Q%�Ѩ2���5Z�*���u�;���J/`u)�:��/�-�A��	�q���4Ԟ�\	<L��=֍Y�@���fR�7&��5�Z��/
�W���\oP�wg�B4a�oH��L������o��}\5�8�ܹ�U�N(u���g��0A�n��5��f�t(t�z������P鴬����<��һ���:��i�H����U^	�/Yozf����ܙd�M'7c��� �;dh�oj<�i����H���^`}ˢ�w-5c&)��1a�rF_T�+GC������r��<5$\��"osCCl��ֱ@lY�\����S�4�U�M��)v;Y;�ʳ%�CV~���Z8�pѧcT�4b[nJ�f#:��[�ejfu�.QÄR�z�[t�d�����f�,+%+�2dB�v���\�XUҢ� 3Lu�NV��K}X�S��C|�V��9���C���f�2s�U�#B���;B�Jìö$�T�śS���Y��⫳~�x;X)������5�wa4�u'ql��1�z�F����=�"0sX��u�ufI�V̚Z9t�t*�%�}B�.�Qޚ�$�v�%��S�ʷ��F�T�Թ&S�6�ݹbb���
$���N��Nj<�rID�m����=��8���n���@Y.��4p�J��{H��˱�L`В��gDܕ1r�_���wJw&	��D�[+I���e�t��r��D���N�y;Ր��̛���J�!���i�&��N�gwn*R^V:|��ћ{�P�YzpN��r�a�����뼅^3�¨����%�:f̭��G�+���zeA���.?eah�\��5�e�VHd뛲�P�Ij�䋞��f�Ž�O1�z��of�2�u}Е�K4�7L��}O#�:ɧ�M`�q�(�[�귮6�A���H�w�qDH��'���X��:n���XIe�کa9)Cv�$�ƥj㑉�;��	��ע�V�LT�Bn��*�A��o���oh��j�W.'8�i2�uG�������b��쬏m�����)����QR���ت�vb<�:�l��-9�R�S��6Au$s�.�<҃�I��{o
LTYԮ��9�iW9�S7w5�xL˩+m`g5�8EF%,Ɓ}@���N`�ܔZ�M����Lݩ�c3:�s��ު�[���"�m(�<J�C���������B��^�'\�zau�b�NnoX��U�I��UєW¥*��z����䬢g�Y��$�Zm��\UWx�Um^#qD����(M���:�����(�s����㢖�;Pe��4��d�s�&n��kE��)乊t��X�Gomڊ��>7��ԐӨ�o��:�*�۲�m*�,�I[���9Y���,̥/����`
8z.��L<����X��g>W�7vE(_7Έi��j���hsΣ�A�'i�w����'��r�j
=iO�]��X��Z�R�p���5���ҭ���];	\};8}T���(�]ݺ�v��cs��t��m�ZGw5!�gq]:9�n�p�Hŉh���r1�-F�9��V湸mʤ��݊��ccr9]*-�뮨�u��F�"�rṨ�.hۘ-����Eͫ��1�sV5rł����k�k#ws�W8m�F���t�,QIͮnN�Xɰj���s��Ƨu��-9ۑ�r�Ȭ��Ns;��h�wAr�j����(����������Ь �����{̵�̌���#�\��j��*���v��{Z�G���H�4X�/-�}�xVDM��ن]UՌ��J�.w2f������S��n�W���0�izO��P��e�ѳq<v��U}�z���w�e�"�}1s�*�H��S��Z&�;CF'޶��8w���9���ᑓ��7o�'�Q.h�qاM�� t���J��X��o����Θp}�~�^���6�HڬG�RC�'�;��S�q7���D@j�� p�"�K��&[�C �_z�:�I��݈���v���']�/S'��N���Pj݅\�jk�I�ƙ�4iӉ932�Օ��'.8u2��~�%�>��CN"5��!����Jڑ_)��7�Ʃ�o
��;�MT_�j@��{ꗧh��^�����ex�)���w�(��?#��Wt����=I��s��2�������Ӣ��LU��=�t:��U�_��'&��S�.�t�'~oR�w<�V$x���� �C��Z=qS�:.)Γ����ۼbU�����V\��}3I`�D��3ls����yJ͍s�A��GW���_Ӑs'�"i��"��iH��F�y��T�`�+ 5a�D�e3p�F��H('�\w}���Ƶ�U�odd��+a�VH����-7���.:^�8޷�$� tjnZ4���c$��-�+�IO�;+����y'C�
����E+��K�����aa��Df�oK���{�2����Xm?9�fl�ٸ��e�['vtp�AZXf9��V a��]��xUQ�ۣɯq��N5��{k���/|먪s�X��g0ў�P�.qؚ�]o-�����a���5����P��^���=�.7κ�^�O�]�&��U�g���ׂ��1�φ\T�SS����g�\iu��ϑ�ܶ}i��+<Q�}�٫���Q���Z}�ATg���c*U!2|�����_����z���Qg��l��׽ֹ#��v�yN#	���G���:8����?�"��[2J��h�q-��5��j^���*튟^�}zq��y>����:���,�Ì�/��'���1w�W�S!����y����T�b_&��x���kcI�񩍯�Ut*�R�"N�d�!���e��bf����<�I���W�a��q��4�q�,�M�؊��l���=<���V�:�A93j���/%"���|���e�l���P����_�f�'��!}�[&/..�ɧK��^��A��wITdTy.�H�/,��ݣf;{��'u����P��g����յ����Ù�o�Bvp��jb�#-���څ�+n�T5}Ù��� �0Ֆ��5҆���]{8Ga<�@WX�o��:��g���2�tŝ�m��M"��b���к��5{/M}�����ܑ_ws�&��#^u�s�Y��+�Տד� 8�[&����F�\�W���ތ�s�5q���.���%�mE�+��f�:��E}�o��i���!������"s�	��A��g��a�0��C3=��k��@�{����[Uvo�ܨ��z����P�++��_�xթ
��:D��7ۻ5l���B�����]��ù8�:�\N�ʸ�m��'Nؙvw{o=Vc��V��UƇ����}	�%�c�>;���c�I�f"���f�n�ͽ��k�sx�c{�r�g`�J31��X��s���~�L��>����#�o�,_w�z�",	�\ϰ't3u\���W�n�^󼹠=4c��]3�p���P�b�g��!�ѳC��� ��ǯ½��Rۤ`��\o/	3'��,>s�z�]~9Va&2��,��/攆�_��DA/�%<�ڇ�y���]�:���-�1�A��zlr���6��>$�F��� �VWzP>��	4�A�{��H�j��h<��@��*/9w#"��-RZ�ݲ�{�;R�%�*Q�W��Aڽ�Q�N���4nA��w@B�s��{�֝e�\n�Q�}5��[�w{�E0��t�9gJae�=r�`SV���ڎ���nXQ�luh��r~��5�E��@�^�f��};=F��j�o�~�9%� �.O _���2ݴ0^�ﲶ�x�4��Fx�7^yBj{��6M��8ܜ:��*�sJ%�j��L��"�����N|�
L�l��B��� ����V�X�븋/6�M�:t'Fz<�-pQ^�o���TH�↤��#��T�L[���pQ�޲j�q���wd�3�Gj9�Ï�T�s�������R�5��Hj�Љ�}^�tZ٭,{�+��e���#�}i�V��:��L��\F��*#9���;��x�/Ɓ�AOj�7�<�+����8��j��o��(c��7��c�*F��C�s���eE��ѕ��ʸ��pvp5��ң��Û7�4�"/����ƟaU�t�y�i����\,��(��ɚ��D�t�6�����9�C�$/H�Oq��{	��|ʬ��ޓ.�����2�w�~�x6��?��%P��Nz�W�${p�D�%����ꜣ�Q�9�����=�b��<�Y���R��bE�H1#
�{e�Szr�uJ�\p�z�\����� �}&��(���۷��2&�DzPv^��&롲�(KguR=�Y��W�(��3F�M^B���|FG�у�LF��������zb�[j�&!�g�I@+�K����,����i�|�kL_�6�?OI��1�:��d֛�����ծ� L��4m?m�L�U��Tb�'��0%���W���衞}t�Y�R����Fz��z�����_j�S'<b�.��X�.����D!m�w���Lyg޻C�dK�B����Y�\�J5���A�P��t]/��7�n=���g���hdˏVU�cŻh7鰟W�s��_����(T%��ζb�E�'�����%�C�4.��9��6+�q���xls�����|��;m��Y�a�{�Fϼ��a=��$!�N0��<��ncb�S��[u�mӴ4dB}�h��Rt���T��i�W��}2�Mz:��������p@N��0d�yMp,r�WO�!rϺ��2$�{'\L���1���k玄��Bk��f�� p�"������a��gTrq�Fq։٣y��iI��(s���ľ���d�m�����aW$���{�"4�ǵ4rv�幮S�,�fb�v�ϴ�x��C=⃯w�ɯ�k�Xr�#�q�8=3MH��K��öA�f1�w�T�-n���l3��M�°�gx��,�7�狅�Dk6�3O�<_	��9��[�`b�ʎ0�_V-�x�,D,b,����yL�����M�v�ާ-�6�v!x��-U����5��ԕ���*����k-�����e3�\�g�tcܴ+���Ά@���꥾Y
��F����X��j�|ɓ��F>�����1�7��Y��m�_!�:�|nt+8�+N��{^���]yp����~����=.�Ηo98� �ܝS�2<�z!�:l\y�%T�򸁵��O�踧:N��(z���	O��tz�'W���=1~��>"uǽ,7+����Ai����\�9�d?�GN/���`������~�{��5��I��?�K� ���:��͜{7�ҋ|��ݳ!�@��
�ü�c��Ңp�X�r�פ�ex=�VE����φ��G���d/u�{�]Eg��d��ݚ�('�z��Ӹ��Oגf�b�ab<�9D!���f�\���Άm��诱��}^�^5TW��+�l�[��)��&~�+�J�ґU�!<��+�<�m���h��g��}A�T���~�b*'usŖn���J�^9jH(E�*x*��s�nh9����ѝ��1�`�����n�
���Ra�+��+�nT��$��� �H�>���L���m�DǛ��l|�w�"�B#�V�j�>���Lf�,�� ��W0!W6���I����;D0��r>�u�������)&�Q-t������(�r�. VY6���h=�b+,Rv��qX|N����	�W�b 6,�&�!���+w7)�\UȯC���y,L��?{��q�|����/D�9Ӡ���R�0#܁��$��ϙ�J+EV�R<�ĭ��Dz6O'��U�d��{b=��ļs1�ꫡW4��q��Ҁ&4���qɝ�0���@�@�R���1�4�a��]��s�[8��-��ҶU�)=�E���8�S�y�^#�\���ٍ��P
^���<�������rh���l8�}Q�-�w��ҧj�B'���Y]&�̐��ê������zk���Hw	��0��#@��g�槯��tB��⅄r6by^�j�<��-m`�s�5{,m.���L+èx<���U{7=���:�w�cf[r�����b�����*GmD��Y��=��n��Z�_�g^hu50�*7�.��ay�C3Bڨs�mʍ�ސN/���l��>�@�U�3�����`[�3d�x|ʬ��<��&��N<ι��Ƿ�ΦѼ�[�r�nz֣p0,������\�WYU���Ȕo�,D��~��L�1>�ٶ���z���}/$ۜ��dɚ����(J�{L������.�^��*�Zʃ�ah���盻�v�yE$�7�	��̓vS�U��V}V��kw��9$Q��H���A��[}Ju�i�w��c�f���q��$�X�8�BNU)r��"����~yk��?��3~KF�	�
�]NG��i`(�P3��x����s>ɻ挋;�Ɔ^��$�ci�z��/�o��Ϭ�)��<X���#,�V�5���gN:���ݎ��ʙ0���Oq�^���x�}�3蘒A�� �c>�����M�{�/���z���.ņ�UcѾ�~;�{�����l{����,�(���@��P��J�^��]�S^ճ����N��3q�lW�����`y�>���z^zf/y�8v#g$�t�G�f�ViY.ܠN�>���\.K�<-T
+�⌲����w-߼l��>ӟ7'�jbڕ�[��JΥQ*&����w���%,��f#dChE�҅`/�-�����0=�Mzg@ߢ�-�!�?�o��Q��j��g��I�����g�K����MvB�����!��?κ�X;�-JyEQ�:X����(`�9۠�����1�ؕ@��ѯ��d�=�E�Ӭ�Żow*��uS�Y����.7ܔ�o�%؇.#]�4.!b�BwM��I~1�E�=�0��dC������WY�a\cUn4	�q֪�V�{��m[=Rtν��������Q��~�:4i�p��l�+N�Y�N�/*�gZ���p妧�����D��i�T}WN�i�B9;&����=Y9U�s��!6�WR�aoC��	�4�ܶ�K)����׾�,!�OP�+u�twt�|/��sq���>�f�\y��fela�����:�4��#rkw8��0�G��r�3�����P����=�U��ri�'?~���XicG �����d�v?��B�8|rPQ�B�)�����Ҽj�_�R�c���li8�^��M���.E�����ڥ�?l~�������I~�Z=mc:/��;j�	�����N��+2�w*��F�0��n�9��ֶ���ʝ7�vN����W+.��있�D�j���X���I��]��9w;r��>���i��z1�%��6O�FGY_�:�ix��c���q�Թ�L��[�]�1ьF5��������~�U�q�Ԑ]�r�(�Ѿ��ˇ}}�����}j2�֌�4���ɟG�-TW���=�ߦ����6��f���[�zc�!�wW(Wƃ�I^�e�?u�2܊
Z����k;��s����=q�p�{�34�y�~���9�����鳞pO�� /W�xEp������4����N�О�������j�o�F�J�^�������S���D7�Z�鸷��I��w�h(�z����)W����c��̠E��pg�p��rv��� ֍a��L�v>�u�#j�0��O��.���쮶\ս�)q7�V-J��MS�u1�;��P4�
t��z����u�����М���G\<R�#܌�l�=���5�K}|<=��ׅ˓��+�o��>�c�F�mn�A�:e���Φ���� p��R*$�>k��VoN�o�g7��uF(q���<���=�D��fn4kb+��]3-N'�b#M�]��L�)��/<g[�;=�dn�F!�9������CN"5�q�����7���姓��}����R"=�*AOq�ka�v�owU#||ɓ﹵������>/�^j&���&���Q���8��j	t9`��SNE ��C'����=�U�^s	��w�sf��ת���V��r,���	�{���gֿ2�_�%�5���xښ������ƽz�yƛv�`6�k��)������έ*:�w=��:n^�� �_�8�h&al�y��$Z����8��]Y��O�o\�{����"��yJ2����!�_�%zz�Ne`��;�nW��Q����׀��1^My�=.1�s��ض/�8����I�� Y�sBL�.`�̴�Qł�:���"�WX��WE���(����z���ت'@�v2�+�)м�P���>��.i�oB�dZh]kV�����m���C
���z(���-І�x.ӀƈIk��j,6�����MgAڐ��_wnd�/U�\�s���9�{01��L�[�e�+�5�Q:^Ɛ�4A46^N����oTR_-�V-,fl,�'Y����y�*nPqK.�6����(�q�i��N�%��k��3���\�`ʼl��ƹ��ef�p����oo<�(����9ei����+b��xe�c�+ld��M��غ�U�Lc�ӀP���ܠ�X�P̮�뮴r���u����H���،z�����c���o�:
pm�Z�mq巵�0hY ����uN	��+��k�]\�-���dV:\�{X`r��ML
ȼ��Fȕ4}�ױaB�!�dt�q��^�X*�w���l��Ou�ךC�4J��eu���C��ye"�,.A��$nt
�3�O,D.�{��~Ȩ4������:�K�J��m8gU���D���G�b�t/�\ʷ�9�ِF_t@ՙ����!�Ӳ6�.�%���殈hin�YjgH��Ѓ�[�lxG(���e��7���@��"̨���������Vh�u�ԭ�t��"0����ȭ2 �woN�!w05ہ� vh rX%q]N�:Ռ����]*Ԧ��Q�.L�}���$�o�ƛ��J5u}7su���Z�ѵ����NB�mBѷI66�A�{�)y�������xlr��-��h�*��:m {Y�Xd�G<)K��)�J�2�e�E��vy���;HX$��Nym��bQ���ٝ����C�Ѿ�]X� �VEoF�ó�)+�$��%:z��{[�Ef`���@�s�Fb�ӫ9���4�P��c��K]�p=��AEx���":iV�s��Ĵ^���F���\V�k�݌�8�L�D$O��V_pǵ����BW[�	V�ǫ�l�+2�lE�e��]}�J�Ɠ�	��r�C:m-� �{E�\o��[�3:��R�3N���,� �J����}7�*�6�Ё2!§F����ZtK�K)��m���p��J8����>Y���&NK�*paf�����:�Z�4�*��D���ͮ�0�;o�G��׹�W)'F�s�ȉ���[j�|[{�{8����|*Ϡי9Lp�Xz�9��'�fV`c�����9�R���[Bq��m�:�m��^�֖^�t��

�ӷ�s��⭙؉ݨ��Y�5S�Iz����f�����<���{U0���]���R=�@Z������/8^fV��7\���"�<3��\�piD��Ř�d�<[M��Ic�$�Y�A�o�r��V�OP��k��f|�ns�!�1����R��δ����:�e��8
��DPG0)��%]�,�nl辪A�D�M EP4~"�"�D]�\���֋r��w1˛��Qp��7Kr�N��]s�sni"��!\�ۜ�E����1�\�"����������.�G+����e�\��;��s�mt��b���d���6�&��͹��.��n�+��uݸ����2��k��r�7:h�+���\ú(�wnF6�wh�!1w\����"�L�k��d`*�p�r����7"��;EsE+�.mݺ����\�Vg:k��-t�@G3��5�;��T�D�$�.ns]��s�˨��)�5�.��C�@U|
�K�p̙��b�7t�1<[B��M����trsb�Bs�p�TX����/�ê�N�d���p`u�z=|z��������.F����
��x�E:��e?\ody�1�oC�.ifv^#�w�DAv�C�I�2��D��PS/�(.��M}�Y�|0���G�F�r���w�v5�ؓ�s��L�b�X�=�aL�H+��0�b�U!qS��"��s�Ӌ�+��5	7yQw��L�	�[�y���o�=����q���q�'�3��}-�����qeЉK�;�~�|�jI��=ܮ<O���;@<^��C�:m̳���A"��Q/x(
&pb^�x��ﾯ^������Mb��mli4񩍧U]
�改與�~�n������/>f���}P* d��$v���C���q�������4u�V�t�;�����ɻ޻[�7�&��*Ot�ā��*�*_���;����r�K6�d�94]q�;V}�9[�Y�N ���oI�^R�jd�+��b��xП��e��T�&����w&�U�]ۺ��cq�,yτoXe	�1y�hתC�D퐄���,.��a�q�W���D+�%���n#F��ߨ�;��\4*Sk���m`<�pǕ�����<����ءv	�t�������c�L]7 ��	d�h��>_�]];�e+�uZ��Ե��t�1�y���SUމ{8���Ы���Fm�T�3m�y�IX��l��@�����1m�s4ܸ��t&���!k�2}_EH��:\�!<��\h{���̾��Czk=�������*��y�C3_[Uvl�F��Ҋ�0M�A��me%Z����,c���w$(J�?Bk4�/	�@a�UemtX�K���N<��I���Ƿ�C��G���v��t����nL\G\Ns=e|rr6�V�����<"G��r��b9�|�3sk�[��ֽ[W�=V�C^/zo���OϦpd�eO��r<���@�p*9z׌��f�^vίVO���ph��}N�f�n���}��lQ�}�z-A�=��c���نf�}!R붝q�w��L"އ^�a����Mz�Y�Ϯ�r�$�c��L\T�G]]���8��������1���x3\K�vޣ��u���,^�S<tq�'���7�f�g��kEm8�E�7S,&i�����l��s�o�����1{Ωø��.�����G��5���Yga�2��P�{P+��L�E��^ۉ�n�8\�べ8u�S��c�3�Z��C5yY?�5���p�z\~���v����q���t�����vOv�O4�:ض��w��=�c�:7��6��j��/TJ���;���)m� ��ZwR@�靋l�5YrQ��Ry��|�&Zm�7rcHm��x�ӽ�eEY�5��T'��(!Q t���҅`/�-�����0��z�ϸ`��#�L[ˌn
�p�;�Bv�UW-�T����|$������8��Uz�r��"�c��W%������	~���]m��'��P�s�AWܥ4hzd�z�T햎{�+b�kӴ���~��9p�)�Φ=�)�ܙ.��.#]�ƅ�.b�B�h��_���׺�L�]`�A����y�{�#��e�^�Y#�緲�wt�|/��sC�8�.�ʋ����ՙ�Nvi-D��ܭ�1���;��\�u-Y��/i�=�}YWC������u�]�T��V���@�x��s+K3��@k�:=7>�^����ըv�)O��s��1ojv�9f1&�;�Dl�y	�~�x+ޛ�g�� ��?�/�·T�J������d1]��yg�������)��b��x���g}�]{���:ls������W+�~�z��A��E�4���p�-D?��pb�?u����ϳ����7�z����D ;��!�2mz?�컋ܨ��&�.����� v]a��Ln��ͅl�[GC��c��ڼ\Wb��Yժ!-�u-w�'�����wG�=�}�qצY��i���d��κ���gU�Ҳ��V�Bl*eJ�.`�c��nκ�J��]ぶ�d��Fٻ�ؐ���jò�����Ւ��j�
�k�+�N��5�_��/U!��^Z���,�D�c�ݥ�4����w
K�/�-�e��p�qܙ�z��*�1�݇���O��t� �+�&~��U��6^"�rv΂J'"�;�u)����+����xls���:���čM]�mfR��$W�/���t�����<�R����s2��-��7��/#x�W�5�x���2"���'��Br�Uq���S�p���A�:d=+�k 9���N=7��yw�jd!c�:�w��79�����T���*x� Gx��>hzo��ï6&%]��߉p�b$y�6�8����/��Yv��M�؊[��fd��$�I�W���Ҫ��!쩽�kҡ���V�Ǚ���~҇P��94�^��CAƻ�!wNs�!��K���d\C�RL�+㒡}/�Il�9����Z��߻�̙49��Г~baJ�//n�O�"8S�F�/��qeQ��/���Â��??�ޯiB�ˆ���\�&=rڱ��Vmwm��\����*�3,�	Oq1��u�E,J��m�Ċ��Vmc�:�V���j���J�^9w+��[Њ��>&��7al봫�����T�S�+Z�T������󭖕鋍���8��ۮ3���XڂS�wH��S)d�5'��*�z�fǕ1� �a���}�E����er��룈��3mvg������Ol_�چh[���Ai�w��޹�p@~���:�����ܟR7�V�<�K�pm�%[�AL��[�s�fC���V��ۡ���t�����,"z��6�=���vf�G�N�����!��י��ƿN7��d/u�{��=2�Ɏ~�ͮ�{�ʋ�*!ܜ�TY�!��iB�Ozn8F�T/J�R�=�O��{Kw���Y�Kj�ٹN'ys@X�jU�X�]2ǔL�u)���c�e��,�_^��-����(����g�I�/�6�A� 泍�r��9����@�,g�R����s�nh=I��yH����\��"Oz.;ç�l=G�����J�1L��G�*���>F*}-��Gk��'�p^�s>&��S��&(O��E�����x�|�z't�1�3�7���&"��w\�:��5��3C>�a�Co:\���؟��hf��S_:��T9�/M�k����c����2^�����"���m��s�:�b�m�n�2�5'T��5�w��bW�u2�u6�]7�4^��B�h�o7�5y�!x\���J����I8�H=�A���ܲ9�
������Mh\�pp�!���v�[ *��oc���y_��&4�=hB�-�@�ӿf��s��`��/�8�m��=��maܝ���H����I#��F�讉����54��A�P�iC�wz�W��~%�����K��0\�;�F�
����}'j$G���a���ŋg���~.��4=q��s�������ɸ%�H?k���,F�⅄F�G�KG�~_D����dX��T����v�Jܬ��u3jY�*���uJ+����r�6���~�B*�̕�}qtC����&��:��4�cQ`"𽿵z2+!�����j�����r�hy�LV��|�9W��1������H����P*K�p��������g{�Ǚ����}`c���U�3�x��pIO��x����3�(�ⲫM�����ʡ��/�̵�F��@���u�q&X���YƆt۵�zZ�W�5A��E��?E��z���{�1�]+�����-T���-�g؝�Ϳ�u�-��Ӵl��3� ΐ����d2���u2��#9FE@ځ܊gZ����J���`��l˽�Ү�!�w>��4��Wn�XJ(嗶�H�.𳂱�[\2���b�w@tQ�mH��ox���A��+yt¸N�+�9.X�i�wlY�p��XU��J믚mNkz巊���>��p�s�9ЈB��q6\ϭ5�~��<E}����N�dv���Q���k\���I���KF�S=X{���p�g-�����rm �e���I�/�\	���<�v�]L�b�!t3��S.=��t��g���a��=F���{���ދ�f����V[�>���BI��L@�$p�	R2�ֽ�[�:!9��cޓ��S]�f�}�E�K�� �_����yN�f�����u��i���j}Is�3�����K2ufxwu��*�C�y�a4t'i�S*+�UR͢U@�{����9����o�r@�M��Fn@>"��~��O��l9�d�"�g���T9Jh��Ɏ��>�Q��t�P�>˯8p�}��5����z�(wrd���}TG:B=���G�I~2+;w�atM�����ߏ�
���EI�6�Z
�y];�R4/�Ú��iv8ʋ����*�O��f�o�ߧs�:�N
��@����i�����e]��:�63��rh<���H�$B�Ƥ�4V�X"w�+�Õ\^/+�9p��x�f�L6g�۞r���Y����4�񏎮8b*���7�@\.#�x齺�ml�s��j��NO��/��k��4������f��kic�:���h���G]��-��;�V��/R��i�"26µ��W\���~��Cfn���A��sq��qx�����P��:�Ҟ��u���Ro7��:����_������r um�_�1�CF�����;y=W���;Xk�3u�(�\6.�ۭf۔��>�^�(=����9'2�2�	�(]d֖f=�3{��Qٟo�,�:�ݑ|�8�ƽ==��K㍵q�o��!o�]#�p�{u�X��ŧ1�zsZ1r�ay&i9�~��8���ܼ��ߩ�,�]�~yh[�력ؔ��[p������:�z��Ę#p�)W抜P�7�reǫ�-�Lx�m�o�i�q�wt��D��5���;�BP��r]|:}��.�{>iCN�����®�~��{�x���z}�ӊ3��w/�G�]�}����Ͳux	�
P0<�F3�i{��sOHq/�����e���vd�1�-t���N��mA�~�f@���ۂtf:Al�PzW�֎�S�������d�v�sؐD�<�hE��0�:q�[���Bt�Ω	C�T��9A�G����][&������o����YFj��^:W'�1X�v�J�ׁ|Y�R�B�_(&���=�9�v��֑�]q�#�]�����S��wY��e��d�a��b�����_��H�x�hy��g?-�l'V9u]M�P�z�4�c��v�.p�����$=�mq�ϫ��s��fn-�ȇ4�.����a;&������kǶL4MY`���h�Ešr9�;�P������_}�&�W���0_���ĺ�P�-��U�S�9��i�q>�Ы�<�#Ca�r;�3Ǿ�2d�ߊ�]�ד�z�@W?��n����)�ς��N
��p]/W�\l�5��ˇ�n��~ɧ�5�ϖ^^�M_�0���-�s~n�c��#>�0O�ۑ�#�)��G<v�0���{�7�������q[�Tt0]�,g5�2��hN�yJ�똌�&��2�k�qG0u<Z�'f�`[�,'92C������ud��γ0��ɨ���e�['v5��k��ٟX+P�kbp�}FƧ�zr��cL�|�-O�x��u��S�{�\B�Z�*m�s�N
3V��L���/I���3P4�_�6��������<s��]�?-��;c����l���E~�����]E
�,*<�S>SS��Agrϐ�K0a˛��9F�n��������ý�}�VW=]9��,��V�or�-�o���jet���e{��^nx�<8m�0���7K��+�m_4pk�1��k*Qդd��{��cC�/��y�W���8�Z6�ޙ�3�.O(v�D�n�ڹ{&s�5rjd�6z���~+"�Q�5�W��Lˈ����>�p[k����,����T�n�-�)�7]Þ��h?;�v9��mԣp�UA�A�1��ױ���U��ݰs�N��7�}WOs����_���^O�l�MF�^0#}��!�O9���qo��MIb�0k�B7>f`{
�ПO��8�'������N��w�D��1��y���]�ܰ=�S`���#�`X�L����_-�m��#�8����kA�͉R��݁?�͐�0�U����K��ʹ|"'�.�@��%i����b�P�Wᇹ�J�RmJ�77��Dy�x��u��&��j��.NL������*(v̯�|�q�C�Eo��,$`��`{�T�_7ΌSr�k�ChوC��F���D����d:�� �N��Y��xW(��ȹ�1��E��uR��C����hM�~�B�wFO�*Gl��6sf�����I�^�Y�����Lh���7Zzo9�fmʇ9:r�h<��߾��3�������/��3��'K�Ъg<��� �t��p�r滾\Mo6(�[])��*�s%%Y1vtj��E����.��}R����J�ݡ�e��wIR/%Z�0B�9q�.c\�'Ε-X&���7)W �R(U�h+�kc��:��"NY�*�v}�D(���]u^���( 5j���F����#''j���5�u1�C��ͽ����H��e`�y&2���F�#��z�LT���ot�}ˁ^f�km#݈�.w=��L�d�]�����`�t��(�7�#K��:\JXѼ3x�m�|�7�c�!T�]ZM:lVv�2�]Z���.��SH�Px��F޻9i�V��b��/������
;�֛"�upA�%cx
�C�y��{�����H(�s*m�K&hDS�*_Mn��]=�L�
F[2ځiB�S�v�u�fk�ym����ӂ�Q
�vѤ����+�2���F��K�I�cf�m��*�c3%��$b�E$���Y�u��'�/yu�s�J�L���a/�'������e�7$�u��w�ޭXYiP�nl�iS�w8��:u��Kv�9��Y�lRn��Ԭ���P�����0��\n�L�}��Ī5[��Ņz�K�.�k,�̾��;��AoY�Ӿ&��dv+%̶ 
��)���w�Q�C,�֨�Ίiв��AKw�0��P�K���e�qӳ���A�e.�Y�,l�WrP�"' dl- wK��	�V�h\$/sz֘aQ�a,�H|^���
�u�WEf�c�>�cL���\�6�rc�Փ;�v7y"�֞wF�t�)�Vs��f^RDL�H��wԠu�e4��샗Ӏ���Nی��U�c�`��:yP6KsxWS�s��yJjfث�R
ѷ�iͪN к��T�y�����0K� �����F�۽�����[A�)uӷ�J+��V�f����� 
��K��L�.������k0VիR�C�.8
�Oṽte	�	�1��%-T�3{��Oծ�0Q8���PdWJ��u�Sl��'O,%P����v�g��A�E����n3W���B�]tWC�t.dkO{�N�V���Қ9�q�n�G�R�v��K[�K�Sķ��C���+�e�e��c3������Ҋ�����[�wn�Běrv����+e�r��k@U�uӡ%j���o;"0Ԭl�J�)@�0v���7OCysTtU*d/�v��Ck9��)s3�6������B��9�D��s�jf��7t%5����]�r�Ǉ�[)J�N+�N���q�5be��up�:����g6S
.e�B�֓ۤ����bu�+�r�:��������W�p�FT�)7�ps)����WzR�e��\�)L�O����_(��bV��X�]P�m�Wn�m�
��R�	�w74�G�2�V���K����+y:ӬY��9��_p�B��C� ���]���wn\wh���Ź���'w�������Ɗ�ۺ�79wt�n�rFH�"�He�ˡݹ\�L"�Gu��e�:#F�iRh���@��W���]�������s��9�4Dș]�˥���\��,�sQ����69r�5˕
H�Bh��+��qF��(�7.P���wnQ��"2X��9�sp���\�卲@�.0�l��� t���w \�G+����r�d�;�]�ؤ�f��`�ns@3I(͘�LN�qۮ�a�WB)&H��Hh�����L�띍ݜ~*�A��5.�'���m+ʹ4ۤ������O0Ծ��[�t6�g9c���kYE\����\�g�{��h.�Y�>���-�tO�P�v�	�t����/	�a^5{}hd*������x�|'��,�mc��]W@SC�s��;��;pZ#N��VUq��H�.���jL�@]Y��m����^���O{����x���o�X��:v��?E�ǩKG"���0�E`p8$�@�?_�I˸���372X����b[�g�����B߲�����@Ϣ���/�Ճ�<3�v����v��C<(�|�����t"�s�6��K�C��<G>ģ~GI:�Gi�j���gi�}v�)�0�m��{�)�G�a}W��7����=�:�A��gم*����{�=��#}*�D�5�g��S=eq�g���a�����O<�o�Ϣ�ʇq��m(� ���d��� ^���HS<R9g��ȵ����Ns�qo=/G�s�"s׷Z�I�p��S��3\����E��0� ��	�V��O�,��.]_1���x��}7���u��0���꩕33��";|LF�+�4.����S��� ��)}�g3��#����C�c���ՙߎhn��zV}v�v�t��	�x% ܼ������=�ɛe�r�J˺�,v�/R�8m)[Y+���n�:ׯ��tf����np����o]�D���TLެP|&�}W�3<=p�[��k����QfÙ�Km�[������!�� F�`���U��ǳ�!�:� ��FF�M{e�T�:^��z�>����и�t��t����>[ۮ��;��>~&'��Ԃ�Ո���$u���cuto�6�~���f�d�2O�W��+���uW�H�=�:�`67�:�����?h4ǘߺkʧ~&�sQI�<.���Ê�=�nf1�Ӻi�ٛ�tF�K
4�}�z�m�R�5�̪ʺ�<mG��{N�Bu+s={<2��{�0���4�O��ߩB��g��gn&P6t;���ǅӝ'OB����4���n��T$Z�y�a��]�����޹L�}���W�o*p�9�=�f=�u%s�xӷUa�R[�9=�;�7'>ίA�O��X���N◺��=�EDY�V�����0uʙͷ��Ic4�-@,K�x�w��|5��/zj�,{�����{lq��?U"��3�������"5���K5'�ў�r�ߨ�	����Z���cŻ���jg���°���q8B�S���b�\�qJ˔2 I��8d���ӻ7x�kdFR�;,�]��h�,���$��7Py����
-��q<���+��л:�dN�e:�}]�Yh]����P�v(�%�r6�4�8ȉbլ�s��u[H'qL5��{刻���I�؉��:�S)L]W�3�晛������+zB��|�L�qF챮K;_�����c.�l�K-@�
P5 �������#�S�}S^͓���o�jI��ӧ9����8v�z��uL�6�Y�8�r3���]&�z��Z"�k����z���z�ul(�˽^�=�����M<t'M:���r��`C�蹋<c�9Y��W+�<�[ z ���	��{b��tYx����F_6��SV�-�̊CU�og'����ʵ��q�K���4	d�J��|wr����a�ͫ�����(.�5��-&N�tg�adOu-y��^�?X-�1+���#�+��å�����F���Vk(u�U#���U+���q���d�q2}ʀ�x��&��M\5�j\z�l�)���\�B���H��7�2*���׽,����	�l�<����8b��|����Q�#��/G���=��s��ǧ��#ll���eUǢǼ�l^sP�k�sL���Z|�ң��	�d?[���Ns&n�=��m帉Z�6�����F�U�:n�X��_vpY��V��b񩆠�
���\8'���t�@:��qbR���լKn�m�ڍn*J^J6��a��H�2��z��ċ�ݖȺw٧����A��cI�Dƻ�Ю+&���7�U�����\�EzvP�*���亲����Y�s��VEw��&־�-F����ε����X�쓯��xF��M��أ�J���V?S���^fK�{-��j�㏞�Ϧ�����n��/����E�9'#6f�gPW^��!��=��P�@W/R����������<�����o��������|먡��QW,e	��|�%���S>�`�Fm��5~-��&X��ޢϑl�w���3~:9�aL�zLAq�
,uJ�.{�R�ܦ��R'�.�����K�C�����Ōa���������dC��a�ʖm�Iux�+.y���v��Z�O����3�n"�XO-��1S��"���퇨��x���:t��SſDog��)�7��v�Y��E�F���b�Eϸ��L��:���z��>GT{�F���daw�P�ywsY5i�-��� ���]T�� NzH�1��Q�����-�y�m�>���A�H�7��:��2�GyRA�����SLә�,(U%� ��HUԾ>��ҫ��ҵ�U޽#� ���R,P�k��K��N��c�u���t:B�x᡻3R��SR��	�-�{%���7O@������ߋ�y�(<��6c�],���[ISJ�Y�3�P�w��.>�54��µ3����%¹����N	Ǟ`x�B㝗A�;0�ql(�sw��%�����'�3l��*��ղ���I؅2CW��g�hm9Zj��|��̌p��;޸+�,>jc��T�_ws�͗,F���f!�i��C���0#+�;]	|d�E@Wu����w���p�=�ެ�ܒ�_5f����D��!��^�2V{��Z����HI���0�p�i}�u1��o-����7��35��P�fە�4�ϲ3.�uݩ�p$OLy�('�n;Ǝbn]����:�}{}l)��� s6�S����ϐ�3�Bm=�	���� t��_�a�驝3d����'�ohv�s�����U�����ɹ%���%��m��nr�}�o�X�t��2��Gg�m���i���5r�LZ�R�{�K����n���׸��<���B�Gc�G>���fX�x�Ho'�A��瘽����g��F����+^�
��?��C� ��b�~}t�IS���cn��ўĞ���� ��$�>� '{RW|�}�%��|=��[G>u��!�_����o���bm���^陴b�zH��溃G�n�r�e�V+z(���ow���:�W9;̧[m J�{��e��
;ؤ�K�#�1��UK�n�/ΰ�j�ԝN[�s+�4e���s�Xn�QP�*Wq�o �[�����dhJ�,g=R0&ƹQ�Ӆ��O/��?�H�q�2��lW$
���l��0�v�z�=:t��ېf��9�:���L�^�~�m�X:vO����O0�1�ِQ~.�ۉ�n֓1Nz�H,�G{�t�_\����~rp�Ƥg}�e����pB,�:�9zxWA�/�U�.:N[E�v�3�)�u�E��OKg0�<t'i�S*(rJx��1W�@�{�������O�ww�[��=���8>���m}�tts��,ۙ�Mǽ뎁�TS�>��L��l=̀��nv{<�G�E�����kO��5+����Φ+���.�ˈ�|h\B���؆T�^��~�Z�.!=E���9���KՈ�-�U�!�P�y]�ʑ�}������}/�v[^��ù���f��c�M���Gإ[��>�z^�]yp���L�]���_�{��&�G���� �|�(��d�P֢�9,+:��z�l�����y��+�#���׺���}��lk�)����oLJ�߮��ƼgǾ_�����@���*s��վ�1��p����m5F,t�݌��K�Ĳ�`��t�*�Z^c۬�����������e(e�ڝ�����32�y�U��mb�hښ4Շ:9�dDG7���Y�a��ǟ]�	@��|-n@֓dqI�W���7j�\�ܕ���գ����ά�&��C
���zg����^f��g}�]{���󝓻:�:���Y���uԇthz�֛�,{L	�k���y{ X�O\�>mdo����P��K�]����J��a/�Ny�d]��!��|s���π�k�99^�Ӌ�1�z�^��2`���w}>Q�J��>��Ժ�{.Q%�KF��=P�������ٟit}�#�o����qsF=�o�xQ�>��}^��Y��m�ʶ���%w�<�@�rJSU�L��晚j~:�\���bƙ����x*�%��}0�a���<z��q��5�>�ӂY�����0�hA}��`KiR������i�T�\�D��˩�E�������y��Ω���v��ۂu�-Hu#�O��,ε\��@�+\���}|(9j�P^:�n|��&��Bt����K5�4po����O��wV�#�焁�K� �{�L>���0ߝ0��k�}��:4�m��󍘬�qz]M���� ���ڒ���x�{ƀ&4���iәq#�@_���;�NM6נ��I���dDq̬��L��e���jp�(�`״A\0塢��1�D����쑬u�tߞ߆�e%�Wx�W�.r�"/>ѹV�6�bΫ�������B��ɕFg����n;I
�ۥ4�����uβ������S`��ڰ��|�_u*�ބh�����'���U�����ޚ���!=� ���5���3YC��>$<����,����|�d�%�/��d��~�f�
�ʎP�X=Jrς�62\�:2��ET����xD���{�7��r��~����g����bzOq��7�N6;�	T6a�l�u�X�p�&�[~{}�0a�i�3�}��W=����3��3V晝��-5�yJ́�`�����h���ՌoF�M��G�V������1�W���*�z|�yzs�4=*lcՐ�ۋ�'�9ۘ��bk��E�Q��u�{��<5v��eV���J�`�o�8�Iy��<�k��{� ��U���~����/����q���=��I����a�W�7\#��\5����^�3���]�7g�M��~��hw�h^h�1{�]E��J*�e��x<��򘸧1ޔ֊�M��=w���V�v��E�`qhE���g��	�������{
g*� �W�*��q�<�(:�5��8}�S�iM���*X]8���5і�;A����Vx��jx�x��s^ዹ�����ҊJ_gF%:	�T�A���jǞ�@�P'+d�g2������gZ�
wOu}.mhQ�v���y�:��4!+�j)7��m��؊���in;���%2k.�.��`���V�zD�[V��N+;�%k�9Iv��R��9�{��[�~�(r6$�̒�*J�H):�|�g��;A��N�N�#�ky�+�s:�|֫���8X�7���'�ڈE�q�GaŭК�{�~�=i��ь�6���������9������zFz+��M�UK� 	�}$q�-�
/�V}a�[�P�νm�剑�s*wdx<\�r�3����VA�۩��J�]32z3�)=�LF�9𬊗��`y��Ē�~���g3��MH�XO���e��l8����qsVʃ�.Nzd�z�UA㬨�����yx/�U�HM^�5���kR��WrGw4Y���c�ͣf!y�h����Z9:~���f�;5��HP�яD��џ-�¨d��=��X�T���P�k���v
��\��my���$��o%�(��N*E�}�F���0�</7WFEb���9X{�桙�j������DxC,�]�?c�u�2<�zr/�A+��Ѡs�
��_#�N|ʬ���L˲�e@Ǹ�J�=7�P�'\F�a��'�=���k�j ��~8rr:����G̜5��o�H�芞w�U���I
��q4nИ�f�r�e���u�υ��p�2&�m�M����x��L��"Qs"j�'�aCָV��PU���'��n�D;�9��*f�Bf�Z�yn8b�*O��A����2�����ˀR�ˤw�y�wJi�o�Γ>��-�e��y�:���7�v/��Ӷ&\Z��GI�9����14%r��Y�t׾���cK����`����".y�3�;��m����m/O���[kj��*�/����Q����3ń��d����pbk��[�~+"�Hyau�����[`��⦝gU�]Z��Eĕ�3�u�u2Ѹ� 'qRZ<��0y�=N�']�s�7�3���2�����p�g�ʟ��ITf:�j��p��Ǹ�r@���6lk�};���G�ǲ8�b^`��6�ݖ4���;%�9 '$p�5�ٺ2��ȋon&��O�w95V�1��b6�Bs�-"pꏽ��z��x=:'���@��7P r��T��+ϟ���
=�}��A�:u�E��i�l��:�U2��fx�U@��5���I4&t<��7������:���]z���߭�3��g���M�_5n��R�/���	���3ОxL8�\L@���mܕY#�3��!rtE6�y��TX��������z�����6��km����kmڶ����j�ֶ�����m��յ�m��Vֵ���Vֵ���Vֵ��kkZ��Vֵ���kZ�v��km��mk[o�j�ֶ��kZ��Vֵ�����km��U�~�m���Vֵ��j�ֶ������)���e�� ���0(���1$���P T�EB	P�"	P��
*�U
�H��������U�E$�RQIQD}�T���JEU �)*�R�JEM�((R��cJ_Z
P$�UI�h�	SY	 �3���hҒ�����!*�H�RV�AlƙQI�ܡ;Y��HkbkR*�kUHZʂ���I�*�SM*��-d�J�SlJ��KF���Km	�e"�((�QZb�m��IJڮ��
Z���   �x(��L=��S�ݙƝu��i��M(�ַi������+lu���@ �cWWLu��!�����ƫ�:YB�Ʀ�T�i�Z��R��  u��p\ƺիUf�qGN��E���(��(��(�U�P��(����(��EQE��QEQEr��Q@QE[���(��(��-���F��9kM[+#V����Nu�   7^h�ڍp�rSFg\�Xc
]�]UӮU5GN����UGZ��4j��q��B�]��k�[7j����5�:���IT���e��Kd��Kx   �<��tt��v������:�4�XG.Smn�K��r��V��;n��s�쫶�ݹwmݩ�ԭ7t���n�չ��]��ݺ��m�Av6�t�Zdj��%�bR�x  ����-��K8�-V�m�v��5��n���.3m.�s�-ٳ�u�7��W�5���룻nu��:�S]��]�)�u)�l�ҹ�7d-΁βٝ�%U�j*����H�x  g���v���'wVґ���k�����YB�f]������u�[+elݻL���-;k�����Ɯ��mʗ]�-�9��n�v;��ヷf��g]��i3h biI^   1��.�esW[�k�i�&]��mv�������ͮۺ+vUMEM7r��KT�[��[�:���5s�\����Mv����ݶ�t�4v����]�������kQZ�ͥ4�[�  ��.���:�Qj��eh�Ɣ��kj���[��QS5�X;��ڧmծ%t�kcMv��k)Wk�j�v�l����n���kin���ң@�i��R�T��HF�   =��wu�7]Z�-�ۺ�gY+��E�l�aˍ����1[*ۖ�9ڧuv�m��wN*�[uE�'sS��vuӻkr��[u�WmR��ӭ����!ٶ1V�Tٕ�j&�E�   !���8UӷKLm�ܻ]��u�mv��a[�a���;�(���6�]�KiT�V�̻B鶕��ew'q[����:5mC�3��B[�|56�ʔT& hS�0��h h�<L��  E?�� �S�&d�����M%4OQ f$j�p9E�tU�HBK&� ����A^��������s?o��0$�	'3�`IL��BC�@�$��H@�XB���BC���ʢ�O�+�Î��m
(�{ ��+�n�L64�ʎJ���MˤCz���<�ԍ�nK�`G��ya˗���\�X���ռ�X��(�)��ڙx�WJ��4��lƓ�g	���flͶ�-�@C:�N�!��Ѐ�weY�+r�b�b�6\�d7�Ҹ4\w���T°���Mi�F���\S%��,}�KݧW�(Rm&.+gM�L5�S���n����]Z�������fhyV��)J�c�{
r�K���ٵ�j��{�G�]ű7+1�C#�a�,e�C&0Y��[�h���d����d��ي�5��A�Z��*��=4�*:�-���[{��@ )�Vjإǁ�x,nc�1� n+�ʉc��AF֦m�ɂ��N�-V��֖�9��a���VH��v!���Xr�+@̸)68��'��\C(7�"W��k"mdʶ�8d�)}3h�.�
gL�EA�q�`MKV^��DJӒ�+��a���]mJZ��9�&�x�
�����ISWE��j�ܼ��n3�-R8�x!W��im�Ca�t�V�Ztەe֣7Nm�Gw��q�NƫR�2E%Q��/NLT��b�ܣ� ���Z�V�2�7��Y���ZOh_�K;��R�eӡ��z�|kPqi��n1@l��%e�E�WE���{�AnP��Ϩ|a�4�2���
E��ݜ���AtM�F�hX���3�	�ܫ`3uP�Tj8YI.ؚvNәD���,�x4����dT�~KT�NL�ǳn�2%h���eh[����N�b��m(ZQ�ni(�J@��kR
�M��P�8�w�>I���v�♭;f�c�/\w37�FI�Z�±٢��v `h@�Hq�B[���hKs�EHJ@t����E�Q��ݑ�Lbv$Ł�(+���e�6X)]��f�#��jV�R6lem�2�(�iGw���j:��<͠4�^��UYf��M1��It�6Iy�`lc����)�	�����@e�!�p؃2�r����b�P*+nЫq��S��w��lG+l�-9���]���/p����_/*F�lMM^�I��M]�&m=��ґjhJ�/U��e����
�ҀܘpݕZڣG&�gee���.η��Ah%��)�孶��i,84RƩ���He
��e��Jf&�Gn��;2��6�ʹ-���ǎ�)陯6����)3(j�v`�/0���0�l���3pEB�m���%�#jMd�JD�ꉛ&�k���|�f^�t�	�E} Y�M�K
lMe ��!�h��oYv�[�n�@p$T�ti*��Dkq�4�z�W��5��֧4���~����WZ�n�K�gb�Ϥ�d3X�����{���A��[-����e�o�eT�]�t��4\y���h�H	J�ŧ{�(F���H�O6����"Zf����݊��Z'@#T�Xe��/4m�.<���r���\�M�uR��V����Z0Y3@���*�iat�w/!���Hʰ��V&uB��@Փ�5�t2�V�!x����մc�&f*�nn�:���[[��@@,��.T�tn�m�J//gЩt�Y�c �t�;u��x�T"T[�0�/u� *튇0e�l�f0�d��c6��phVu"��ci
"��77%��(�:1M����� -֛��V���.ժ�-��+-Iʕy��ƛ��u{�� ��'+aM�֌Uv$ь4UK���ٮ��Ǹ��Ыa��@84��$n����z�<7ko���%�����ԥ���[Ɨe[r�7����2��{��rD����ڋ&�.;�g�훅���F1�#6�^�{�2N͖��qM'V��7��n6]c���13��@Xԯ5�
jAIkz�lP��l�	�BXEVkЪL��f����镏�Z�욵��mc�ݗ&[��įjU����#��YY�Y���%Z��oԆ��MRϘ�2�YopZА#j�R��ꕚ��j���/^�lI�iִ������V���5����#
�d*�[{�N1�(Yba�iA�
g.�������S�]�+R����V�m�O2�{���Ƭ3^]+�uksh�H��M�h��Be41w_T�En#���J��Y�/2�S���t]�i&�� 񸕵j}�n%��Td��ka^�>5n��f�ޓ�*%�Z�Z�FL��)`���3��lL�7]���mc`k�oUj�-휌5�� �-��a��&m`ł�d]]��r9�r��A�</�{� ����q'mb�u���R�۩$&�ҵ� ���;V@KB��QIY���	�<U U7��Ch�u�%����୔�Jl
d���d Ȗ��[��8(�����Jot�;)����v���wHK��7C\�4�{�&���/v9PYV�`�*�6jS�CDt\����0�6-MJ�U�c���p ��a�s$�\Oo4lͼ�J�i��ݫ�K�G&�oג��00љND��I0Q�Skr�Jq5��+F@�cl�*�v�F`�h%�ceޤl|�l[���	��/S(����0�*�ܤ��Y��h���
���[��EI��F��j�x�U��,�sC�N6cʹ��\Sf���h�n���x5,t�a+4!��OwFԩ��[I��/���o�I��m΅�)��To*c�Pz�-�D��5�ݿ�3��-���a`{;B��%���e�]���i�V)EwJ$�]K8	4+X��D�;�!lkUwL��k<�������I�Lem�N������Ь5j�豑,����&�ӡӷ���Y�R$ XR�9��k���I��������l*���%��0JF�:EŲu�*ݍ�r��H0��r�3p�$�$ A������i���Ҭb�#����0��Kv{���~h,�-��i�c2�h��i,�Q��d�6*���#����Ո�� �)�	��r���͍�[Wr�!Kp�,*X]m�v�:�����eڭ9nSZ�)R�u7e�)}1N6m�"kh�Vh�1��Y�魥P^���h:Oi�%�׳Cvv��g)�%ҫĔ ��gl�n��Son%Y�7�n�5�m�LqS���+��a*"��ˎ�Y�:�X�A�if��l���9.�vZ{����'(�B��ˤTB�Xi��b�V^#�;h6]E����$}�j�+����Ň4�x����1���k6�K���Y�M�W�8������Ԭ���l���8�K�J:�FA-[��Cz�n�`������*�
�*Җ֌֥A��us ��]�V�i^�xK����^��[��+U㷮��J9"%�0]�Xo
�^�[����:�eQZ�iiROW��nڳWO&(#Ze���(S�V��K�9*:Yg-l�2�Sz� �&�QhX�1��Ք$�a�N�t0ψ�H��l����-��j��le��jq؉(9�	����ż�(�l*�K� [�H).�a	�գ�����v�ࡈm]�Zh7&ԙK�1�0[�N-�ʻr��K~����Q[�5��wjn�g�]@N3��@�Waͼ�5k�X�VG[eҀ���ղ�a��x�V0�,-��$�ȮJt�\�lS�l���MY@��Kl]�J�W�.���:rP��T�I�VEXeJ��:ʸ�H͓̽h�����NdF�#h4Lv�!�"�꫋*\;mU�l ��^�`CFjk/+��b6z�'+\0��I��u�z�Jw+)��|�Y$�orK�5m�Oa�[����Y���ȝ��h��rl�R\�m�z��V��V�1�.�4�u$�J�h�3u�����r�T�����6�̧�����6�n��Nd*]A���ٕ��l�`Bbor���tf�������RJR`�r��Y �2
8�Û��mJ��VRѶMGH�/X����C���W�υ(�[�����N�ǀ$0+$�P'+׃b�����m�6icrh��Av�l���4�: �-e+�x[yCv�1[V�e�*�V1�T�om��EG{K7v`	�����r�ǂ��"��a��5���z��RT���̫I��cri�=����b�%��QD�b,�jVTj�Z`k�x�&�-k��t�#I��.�?�/1��oNϡZ�*j���/E.�5{[;g-?(�n�ǔ7{���E!N�^�aB�Jw�4�[��$.#�Z�B�!oAljc���)"�-`��c&]��{K[�`�X�e�f�'�h'`��jk`[yV��={��FᙐXL�Q��(T7n��%;E�a��:]c%���UmEj�ٸ7)��+1�e�TwV!S%���«���\L��n����WkhP��b!���߃I���Kfd��a#r%V�Y�4���x���Q�a��9B����,��Y���B�ӑ0,L�6�{��ң�F\��o1j!��n����=;WY����0jὼH����Or���A�V�A��8w2&̭Y�n�G �GR͛-��ѷ�,��Z��,$%V��m�#$W*�JJ��a3L��䡔��h,�3 �(�!GM,]A�Dq����ƶ��u���J�i0D�*f��iA.�Y�i�P�YA�� �q��[-�rT�
<�Բu�Jї,b���bm�B�؅:ښ!yO.��h[+10�h��E�YQ��R�B�WzFBh���EOc
��w��~7kM�f�n�۫-��JV�Ԕ�v�Յ0�m��67���*�s��k��~�&�ķV��x̊�mjSm�WP �VX�4�A^�r̫�[��,k�Wi�U<-dŔm)^U�,":[z��]ೡIq�R��KAVcX[Hm���N[1�uoN|�n�Z��eWL �u��Ja[�ٗQ5u��h5Zז���$�+��(,�᭳�͙"߬$b�z� H��|u��FN$6e�̬6d�U�97]�A���t#u�f�ڰ�6��]�	 �A����G�i;�7��Wu�;��"6��nd85�´�T�h�r�hL�f��EU�%[d�Ɉ<����m� �:��,��L�/eEyxVU�"����U���DM� �67^J�B�3N�ݚ�v@�y���-iԃn+��"���f�W�kɥ^�$d��m��Tu�fn�(Y��ӷq��A1��j1�&�ƌÂ�2�J* ��4of��xt$��wd5�$����C+6$3e��Fj"�R�γ�J�`�!X[���1m[��݅d:�aC0��q�M��4LG� �1����C\gwN%[]г�<	;�(Z���q#)��7�ʸ�h�
b�ŔՔէ��ii:��P	au�qme�
jd*L�9j�eɵ��3q�%�ypL�4�Ɲ����Hԕ�u�ZV1�Aq]�{���w���������\�oSWE��lmlySv�|�e�T�ˑ�c�5����M9�K�
p��0^��[0��L�-L��ȑV+rF�8襂�[Yhoa�f?���-�2X�N^��1X�aU����-c;B���I��5��KVY��F��P��D08�a�Z��g��+29r���y����.�-�JYQb��2�'��s�)�ѡ*r}�����NЫJ�s^#�h�W���2�W�����ʠuK۷�G.R�4h$���Tu5ȵ5{b&Χ�B���4nAhe#V���2�mҼɻn�͘�*�%�5y�*cMÈ�y�CN
�)�sm�4��������́!�I��+]�;Vb�֔�ҭ�LR�V6͇yZ�U�5e3�d�N��q/)\�R�vԊi�����v۔(J*;�CUF4�Ս�7
5s4ܒj�5�Y	ƕj3 �> e<�
bۺүdw �4Z
�5{
�����Hf,�Xv��Y�Ԓ�J�t[Lb����k^�kr9��ҡ��T�%{0c�T��=�oUn�hT���(�~T�Z�F�;W(}{��E�0h��[�AB�3d�1X��꠮3C����\u�u,�e)̷��R�]ՓMT,�*�&^�P򤆱D��͸���J'l��A
)Z�w�*�4��KN�g�u;:TtAZ��&
Y��0V��#(�@ʺ�P�vۂ�7qǃI�)�2��U��-��7l��Ӣ��`kB��JUu,nҀ�ZT���HV�rVT��/��F`ܩ�������te[T�2`�*h�� ����U���`8��U��Y�ݻ�&Oǐ|�`��Y��.aQ�5�n%SRqE��	w�j�E�9�3!ʌے�k*��4�U�2-c�vRC��:�ڰm�KAݫb�Q�M諝e1S�	��D�k*5�����b�Gm6%ޏ�e�EiYV��[��5ڸ�bP6�70X�m�=�VP��D�Z�>�Rqe��l[y¾�̵
�3�.�]��$�-{w��o&�5�"��Q�jYr�&����-A��Qbf�`�.2#"�+V4ȋEݛ�F�Sx�����(�F����N8�f7�	��n�v�Sh�n�^��ɤ�Y�NaB}`3��Ը����M=ro.y�n9ElZ�rZ�5K'6��|�����[�Q��
���VDY�
�:�3B���j9W�^v"��E�&P`LF�B�Ei��q^\ș�!9�P%i�*AE��I7E��rhthZ72������xK��m9<uӍN6���M���RRW���lՍnE��ڂ�<ʵx����ُ���@f"�j��Q�R�p�d�v!9������<�C�
.Xr"6��r�K��T�}R^Іʷ�w9�`����}a,W;�7	�[W����U�@km�v�ޜoxf�f��C�Ӭ�����[s����Q��j��x�G^s�j�R�vxn���tw8��I����:gV��=>k5ܩ/h�M����4]%%b�E��L�3eq�r[3#S3aZ�Q!Cp����N¡�m�������I�ۗ�x��H#t��X^s��:���bx��WQ��təA��plM��pd��#�E|6O��̑�gbJEVWe��lz����m�u࠻�k�F�G��6>�wW����q�FO{w�u�C�G��_n 9��ֽ�ˮh#�dre'\1�3�����,B�����;4��6�V�&�G�+����1����(U�Nm����^�U����ы�ؤx�TG.c)���J
M���_��YFm�t�v�sEt�:*����C7�l˳-^��_<��.I�t�%c�唗��YX�&G���ZM�V�E�d��W,�V�A��a�/�����i��â�	�R=�O�J�:iaa4��I�"ez~�FOn{o�x�iXi.9F����j���;Gj��W���D�R�!�.���F�R�P��E"�˒�D^�u�Ϋ6m����Z�i�NR���\�^�.WJ�,�;{�wR)uǓnB���'��SH��嶈݊`q=59q������(d�e�������Wj�,�o@��*�Ed���E���o���[��1�������>���V��"�l�e�x�����>�	�t�@�+�3]F1U�F��D�o�nP�9�l�|��������:���V�rr�b����uJb��1D����V�&͓�Օ�Ru�{���W���[A�"��Y�	��j��UΚ�Aw��|��L��J�Y�N�:\y�[����:V�5�0��I�45�nj�e>';�<��W<T��/���S#6�I���� /�u�Mrm����ux
<�
Y�C��j9 ��.ܺ�`��&��r�H�cu��
	�f[;�\��aO�X��:R���8���,P�6L`XΝ3]� ���]CQE;+z�b��c8)�	'�I�d���u	4�꼖E醟3Xt.q:mK��Yy(�y��^/�ǽOw.�Lг��2у�T|��&6Mo��9VL��VM�naDWoZ���o#o����U�O�M��	��j�)����.*��B��o
ϡz����n��d�A[����{*��dF�N*��W��u=�_�F2n��ǯ��k����N�rt���<0;V���3�*�0��Zh��I=�鮗�Rh�QT��ts-f�J�:�y���#�RL�QJW��7�w���^�^�Cݔ���0+�ch�j@FlO���V���w#寴%������U�u�{�jαJ��^"��������5���y-퀂�}2��C�z�D�+�`e�f�bd�����w:��mX��XƊr��L�5Y�]=;e�՘�9�{˷���*��e��(�y��k6ɾ�%q�N�<s��S����7i�_ǣ��}�NiG����x�LH)��vI�Ԯ�s�*o��Rح�i�yQ&�i�I�X��$gk��������A:��mI�xNb������>8�g���
g&����[#�;��d����e]�
',��n��vZנq�N�-S�t��T[[��ȑ��-�����v��,2��vgk×��]����ӫ1��hx��F����F�����,^�O����i�Fk7Z�6s�f똵�@�aje�by������x����t�Y۪��%`;���o�n^ҭt8V�ݬ�W7�T�/9L�wD@�2�r���f�1ԇ7��� �m�m���Y���8�2o�L�+��C�,����yV�Hp=h��x��)3����ٔ1�Skr��WW�uw�1z�٣��Xh��GҬ�-�Ep,�U�+b�ͥ'A"�ed퍒�ʼ�.���PB����y����MM9e
YI1c��u�� QL�mĶ�+�'-�}�Qn�9��jT��(�Y$�+/f�+lֹ���P��kjvBwo�#1�w۷�nѣ�5<= ���� ڒ�˓�rGPy|�7�W�S�-��^��G/�%��;i�9��SR�9ڻ7jŬ'2W�RFZ݁i]/	毢R��f��c�:��/�Jv����]���Vx���k$����Z�L7tȳ�����R�^�r[)CWCF�0r�m^(��R��qRO�{�*G&�᭞�,!<\�5��S�-;;r+��(��p�%h��C�����1;��8�8W[�P+}��^nW>B-��9�%�-�k��k4��t��GL���z��p��7�)�_a��1]�����X��m�7�7n3)Ww���ʩrG�*W�6�!�Lj�ge��j`4�5�vsɉ�;��U�/�-iZl�\�%�6�v�u��M��G2CQ�޼���Պ�!�0|���ػ,�Uv��x�j�\��7����X�P����b�A�����o-(]���b1Õ���1��4�X�4�v_Е�Z���V��p�7)oV3�`ZMf�!��HT*�8�2<�:��Aɓ6��qӽ�)�J��O�yǨymE����z��-ם��vV%t���<Z��ob�Kb;(2^wR�����]Ca��M�}8	�eG|f�SU]n��V>�iؔ4��a���ه�'I�_Ʒ���hL�B|4��]������u�|�e�V˺��q��A�_#�\�c�˭8ҳ38Iӌ�Qo��R����a��|�͉Sޏ>���[�c�ׇBb�wJ:��(^/��:y����N��S0\�j4`�Ib�g5�m�R���o.��o��WR\����k��a�yC�_e��ƞ�(�+}P*��;���B�[�t�Ʊ�Y�7�_,҆�{��aqY������\d�"��j����#第E6!�q�#������HC�R�� 1�gvS��ם���&F��<J��.�|��n��({Jh��DR�����'�%J�*m�9��sz*�ɠ�[ �I[i�=a�:�+���OVf��U�o���W�9������p�ta�eBKMf��v��WN fT�/��s۩��y�U1KV�P�<&����ӝMV��G�᧪t������Rw��u1a�r����w\��M쨣��u9jB�f�p��0�i��uv�X�X"w�����9Gkx�$�y�=�Sm��Y�֘�!J	��ߢ��b�2�ӯ`���O�lAmW-�d��[l���nsj�Or�m�[�Z�sX���Hȥ`t"��W�M�O]�㯓�t��q��>|Ɓ�Fs�D��᮷4+��R�\�y���(���HLy�Yq!���\h��01���.�5�o)�%˓y[����/;]�qfB]8pԀ��8^p�wBQy���	��m�υר��:R�f��e�ޕ�
�
�Q��:����*	����Ҹԩ���5H�t��8���iά%1��B&v�`�%`a�I��'��-;� U�Y�0����̝�������/rn�(��6�g�nu3����R�1q ��^� ���En��뱇@��9������%F����}��*/�����Z#�|kD�����|�`�k�(��V���$��T��o�6pð*+`�;��t�x��b\����[|�R�Z�
��GZG]n�~�l��.�6-�%�(���+1H�	mѼ�wR�)�������.=6�2�N�a�I̓6'�˘2�Ɛs������UP���!�KU�w>p3�y2����x��K�����n�%;.|��ЕVs���1b�u��j�r���%������C�LKB��ƒ���&g,�M����`���%�Yo5wPה��Ń&E{��跺���^h(����'vfcfMq=��s���m��jn�A�s_]:�Y�`�o�m�������%J:Ρ%M׮I�aH�X�)ԫ�r��L�E*�:��T$U1�s�~
كv�0�	�Ѭ�'b4��B�n�E!��zo���+�*Pd㜹��^����k0�x"�m>�}dz{<�)e�7D��(TA�#�P/-���ܣ�e�X/���X�S{:m`�c��ЧXs-��ۻ��)3z:�V���/^�Φ]˄�����e5�oQɍ���]��ƻ-�q�F�iF5mC9�ݮjZ*"௧qH�fZ(���m�9���m�>�����f�G����s_�%�4P�ݠ�CƎƖ-�OgY(f�i���m������V�k��kB44��*����P�����6�|l�9���Ůѡ4�Yk�f�j���޷��m�b��av�U��հ�G%Ƶp�*$L���YFԫ��`��Jq��a���q�Q���rgA0k]���q\�C����V_?�fŹ|�ԕ����`ȓ2�t��er�clX}Y��7���SL\��Dp�p�8�$�!��=N���vO���Oz�MٛI �	v�;��|�:�<��D�į�qڽ�0C�:%;��żp�wY}�+�b���6vݥc��2鼲���h�6U�[`���§WD����91�3u6V�np��5j���f0�t���5�"q��w{p���YZ��/�z��&,.��&�i���۫j���� ��S�:�5�Y�*;��������!:ͱŋ��3v�Wt��[��u�0���療��֍݊)`�2�az��ӷ��t�i���xzF��X8)��񜀜Dґ^�*�So����+B�N��]]���]k��ۢ��z�k�V����ʱ�����IT6����[�]B[���Bފ�u�zq��b�M�V>�cS
:e^^���%�`�̷��K�:��nt�S+c���1���'$͕v6�`=�Z�.[����X�>욫o���N�o�:���Y�N�쑺�%�)(�[���n��)��^������$�
�]]en���˘���!C����bȼͱ��:����D�"��Y��쬺WSt�s56A@���|	,R/��e�R�wJ3�� ��v�&��L�;����p�;�t霮����@��C�%Ԛ�iD�;FuO&���
\!��:e�;��&�Q��]Xn����K7�*ˮ������4c���E(%y�:ޙI7k5E�������/�%C%'y�bb��t�7�Y2�םl'�t�,c�˨zTnʅU�$�E��=����2�{ه):�fm4P���i�×��\F�4vހ�a�y��V7mGÊL[V�sSދs����j搡��[t{Y,�:H-�&,ս���G�\��j�b$�Wڡ�׹��
�%2�-�4����t^�e򃷃x��+y�T����lw/�օpML�l��1o]���Y�;vI,t��q��Ȣm��׻�i9]���g��3v���.�})������d��8��Wc`?���M��p�E��q4�<�Υc�;�yX��*x��yt�ZÚ���k�A�Zg%Zj��3���$e�$]�m��KXx�:v��;�V���Z�8�aԅ5�XF�\��]>ה�5\P�|��fs�m�b�2�ً�x#��N��q�ޙI²ѩG��jE���0g-oM][a-I;���T��f��d���I���=Ó�!����3>�p���Ԓ*A��s����VB��93���f�޻ٝ[ʹ)(Ě1�_i�8����:*u(�U�Y��@�\tV�l������fu.��e��c�x�鱮W����-��E;Z?$��$|��ű��P?h�V]�� Y�Ό�ʥl�`K*�W��	��� �����D�^:+���Нk�r1c\�C�>˼�;�������Bi���YIH�-t=�Bv���Ǉ4�{�I��5M����LAU�2+&�fֵZ�W�9Z��ᎊ�_T�(]�i���S)5dVĞV�.̻��,=�� m�חx��f�p�+R��\x�W,�3\	��kޤ�{�)�v�jHh�9oX������JqPf���8���f%/���U׷������{����QC,Ҧ1�.�^�娾�NJ|r��%0r+����յ��Q��Xw:�G8��^>7C|�.o�.[׽̪4t�)$/]��%����Ә�E�zyVM�9d�C��aZ��1U����z˺Ď�V��+l�Vud����a7�2�Vfe0���7���{�9���\)Ԭ����(w��0�λ��\�0`P�؃���V����[H �m�>;�4,WRϓ8�7q��.�]�.���5���c]�7���`�eI}j�$k��m�ہ�����*oU���]j�u���lrsD?��������qb/s��a�-�N��-���3���b�cK���O��W�M�'%T�M�̯��K:Y��l/�f�̚\<{Z\��2!�����Ei�X���A]̮E�_;˺�S����Gn��{h��яz�"kY�u�mN��`'�٨�5��ߕKӚ�C�&=�|�r�K��H���GW�W�ūi����wR�Py�v�IE�
�ϵ�ɞ�n�Vc��s9Χ'v�:�r1A�j^�IӲu����#�Rt��֮��fV��Ä�*TF	���;p�At�n(`]�!nrTX�\�����}�qiV��
��N��nTܝof�Y�6��2�`։�����ԫ]CR�9�pY�K_�g/�Z��NS&Yٹ�V8u��T	�͆"F�(2�n$��K1I�Qj]�ą�loe�j�=0ʥ��0VV���,ʔ3�syoxx�x~�{��_}�e�"����'�+��F�%#�^�[1�z7��Xb'�����\����ĭ	*�Z�ʠ�������֣gBêMsS&��E��%dݍ�:��}�.�+7�J���oSq�4��v�g3���E�5oq��i#ӳv�T���n$'7t�n���GY���%tQ��6�HA���g*ܹ#U��õ*��s7�r�c��y]Қʆ����E��]�������:���g �� ��/�d�Q�-x5�J��AN��8����Ѱ��^%bj�t�)�+�ms|�X�� �5!E3m��JY���W�{�$Vy�ڜ7�9I	�ƴԇHDب=(gRq�%{��*Sy�W'�k;XK;8���m�SB�����\�ۧm��#)[�i��R�R����T���X�5͹7��f�%uY7�Oc]-��i���aW�1�o���$lЙ ̫nTQŝ;�����'{��2eӽ��fGy�J.ImX�HY]��-���H�����v�7~86�eڋ7���=ղ^��zx�.��+p;��9}�rg*M��U1a��r��1&.]��żmk�v��j�'6ɮ;Y�u5��n��!Nܮ4!)Vn�����A9n�[�C��(���kw;7II�k��2�I�+_CDcF�rc`��7��x�Z�Ƿ4�����ws8VRcL���[qS��`<Ф��v��C58EuB�k0��"5�47��2*��B�O�sΜ��1���1�i�o׽h3ۥ�p�a���PY�� �tq"��"�k�z�m��B�h�)8�v���%�{�wQ��NR�f�=L�dn�.��:v�[k�Z�+��/���V໐3�+�^�8�ퟏVo�5�>���@u^�[x��	%��c�+y~ѷa�ݳF�<�r`��Xm����X��6Ⱦ̨hn9�"��T�«Ŝ�t�~B� �����Y]JfTltO��2B�G;N��h_j-�u�*�u� ��@^��h�}�W0y
wL��q8*܎^m )����(<�H���"�͸�] P}�y���p�7q�z�kp����Ҡ��ˬ�¹h���%^�:8�X,44�[��ѻ�3�-�� PyH��ZO2>��#z��:��H�ѱe�Ek�O'.�FwI�Mfg�#�{5s)��sEw�Z��R�����ǰ���*����C�6d�S��i#�7vF�n�d�9nh9[l�.����<�÷e�
�����`-wto�_!7Uɨ;���D��L\nZ�T��������I�|�]�^���6_P��sj[�����j�\��QZ���i�3&,8�1��w��;�ŭ����vhlwp���i��k�=6���|�	��`�rD������r��o+wx�VԠSv&�^S'6�6�|�W�� ��+��Vl���qΈٚi�K9X����5ӵi�����ܽ�V��i*�v�|�u;��Fg!aɶ2�kڻUj	�)�/��SX"�(*��tܸ��es�#L�h�v(�{{Z�I��p1��à���F.�6�k�U���ܣ4HH�����^tY�����w
�kv�jI}��ۮS9�t$�K��j5Z��5��C�ʷ*��V3&��Ua�D�i��yP2U��]�����ٵ�fu��g\4�c:QY��VIX��Q)a�#�y�S�I{m��+�;e�$V�wOt����n�����1����cF�U�W4��U�*���f�f��8�Ʈ[���^�.�7��o�6sK��5j	xX��H.Ġ1u���1�	����n�
�wa >�Q0ZU���P�@J��q��lӘk3���.��л��R�G�Z�E	�j���a9�A�зq=�Wm�]W�vA��E���������D�Z���$)��σ��\��ڧ]q���u�%����+�JnnL��xۨ`'�N����.F���@�F���]�^�A�}��D���dI���%\s�����l]2��(D4�y�����v�#A�eZ�{�\��_2�F
�B�K*��᷁��G櫨ؐR���E#��ZV��i�{�f|��o]EtK�jk�z�A����s3��zL�$�L��@��)g'f�e!�{�z�����Q�(_RD�9��-*[!BQ��-��ͫ6��<�P�9���T�G��y@����˭K���A[Zr,��Y���Js���'M:r��\;�BE�m��R�d�/4��.�����b��`��f����[k���N�3o/�4�/@��\,a,%ap}�E�6���� ̘�&G��j�m:9���Ҟ���ҝy�a��=I���]�ө�L^\��⩃��47��&�@�_v��gsY�=|��l��S��&P�Vw�]�]����aƠ��T��d�Y�z�\}�M����u�2���=w2Z<�]�vu9��hl�࢓@Y��z�z^��B��*����VYx@��VN���mv���6ʆ�H8�ڷ$��Ǣ噇Mw�<�`.�s�=��R�RA��f�K:T�C[7i6<xD��n���(���'|�}B�8Z'uAiވF�7]��y�r���t�6,�v���mA��jsΠ�ѻn`y�C�f%Ѭn�U�9Y~�➖f��EJBK�F��l��W�A�j�.�@72�v�eV��`U�jjs����y�ֹ�wׂ�p�G��1�v�������Q{�f��d�����j�,��CJ�P��F.g:�+��Um�4{��.�B�J�wI���MP��-z�'/����WN�t~RdV��fܺ�����ә�JɋtzX��3jw �j��X��]�Gn>�m�EW�lIkei�l���E�+{���&��\HQ\7��eZ��	���T��h��-��Q⢋I.VlZ�s[yz5����*[;�zW`Hh��Vp����ѵ׵�J�M��}
�*���Eb��7�a�hK��r��c7�:�.ZH���SK��2ﾼ�lFV��s�p�*�SIt���J�������8���y��=��)��o�/�n=.�EF�՗JPE>WZI��aֱɫ��y�Q��vUhf�%5I�g\.<$���|i�[�[�[�����c�����^~a��[��Wܼg[���4ѫ�j�\��WU�7��wkn��p�!�B��kI�:�B������²r�{ɴ��V�{m�h��$9m&r�p�����9Q�f�2�apX�9�j���6_��2�9�uϦ����u�X��R�	 ]���0&�W�V�#^ZZ�b�R��>����p�T^M�g�z2��V�J�Ě�h<5���g�ר�hZ�]]൉���9����W�U��B�V��+n���I�Z���a�B��d��i���Cw$A�i�+�2�q���3qJ�]b�0��Bԡe�
g���ʂ��8����[t�T�Ӹ�Ȣ���ch���奈sy;��|�J�ͫ/�7��[�E��ک��r[�S�o,��b�ʥ*�/kG`|��.�q*`IB�;�92%}�4'\Z��:���=��f:9O�Ԕ�J�/^�lm�9.�Z���퍎�5��?"��IԲ���Ǖ6���`��n�f��5s�"���ԅ�b)�(3�t[X���ҕҷf�z�~;�wR�EV�(�EJ[�,K�Gu)�q̏B�>4�xv�J������C������nƩN&h�h�K��xi�&��.q.�]�ka��X��j�b.��[9(�ae��Ɠ;A�)���7���3`���t4��w׊���P{uy�P��v��
ڜ���Խ^+hϲ�C�BxX��`Y�L+�$�6'�8����t��*b���
�ɖ�m��/QV�Շ6��D�`41d�y���)i�9�z����;�y���Q� ���K�Bm]��Y4_G��o��=u�v-��b3���]�.��eWwD�{C���W�6fұx�䮲ԧo�0F�>�i�,�e���
�|ʾ�89ݳ|x�����^����cW�V�7I��N�;;��X���M��Rΰ�1^s����hc�ܷs�Zw���U���[h��/�\	N�����O�,o*����h}3��7����\i��軲�;ɥ%t�{�Q���jY�W��30KnSUqM�8L�l��^��YҸ�N�U�Iy7Ll�D��#O���{ f�;E5��Pח��95sNXp��Q9�Iv�p`X֝�˙=����ɍ��خ��n�yƴs��ϒ,
�)�s;-;�m»3x�*���Y|F��)n�������\��Ӿ�qʊ|:Rq�5��A�� k.ᕤ{Z�dy��`�Rm�־�{Ǻ>4��31��hi&�XU�q�L�6�r��g^N+v����'{�����]������ύc�6�C�� ��fVe̓��I�sV3@��Sw����� ��m$�Vu��������=��C�Cr�Ʈ��\"��L�3@pP�U���a��:f�J�b|)R�)b���ɗ�Y;�.I7k��K`*�v�)�*UQC5}��K�U���Mk��:�����
S�p��j{�m��{���c�">D�vk��r�O�ݙ�E�0B����M�Ed	c�s��t�̷a��)�]RԼ�C_^7��;ͩi��i����&�3w��	���k~�2����Ȼ`8��⭇1����u�W4t�x��z3��=ϫY_v]�IC:�ܛN��9 ;�gصat]*�N�t�B]�te��(�
cMP��#P�.ՒM����5|��P��3���a��.{D���?8Q�E�M]��w�M��d��S�K_[�Ut��x5^���Nᗕ�ri���k�&�0��2c�fT�.w�B���qZ����T��i��ػt펣���Nu"���0�=��yR!r"���`=�|7��;��
"s	^-��ٓwiKhKMғu!*�`��vm���Z\�.�Z=���{՜L��J�/�j�4�XK��'ov�f�<��a�[��֖#γ^��S1c+Vp�(�,9yZW>�H�*���i��9�=Y�)�=�L���b[7�#	y���{���mf����꽐��Kuņ�h�y�Y{|Ԋ3����c�U3�h�̥���0V%W�����"�6��JUe��@�5�t �K��J�����kx�h+ok��9[f�T�h$6��%n�1]SE���"�8�b1~}2�v(�V�em�����T�1�ُg9&�Ky�Œ��7�h�t3��+����t������m֦�V�|���)�~��+�;�[o,�\m�tjú�r���uk�n��o�{�FQdk��nd}B4�˭���H�7��ҍ�˫�)���^����t�a#�ڰ�tĢw�cɜc�k�B�9֞�7�]��9u�-��ś��t��)������s�W*�Q���ςc�i�o;.�w��):�q��fD���˅FB� �1`
\�Ѵ���o\�'�n�}�e�jL�ڔH����I��r�<�{�Zj(zςC_SX&�U�����_ˋ�UN%Y������E��uԸ���av��)��KmZV����$]]�o���J�wT]�wS�PSn¨���+tj�����9�K�����Ѿ�A%v����ukѹw�/���Q�Z��S���}O&To�ZY�8TQ�f���7�Y̧RO�ܠ%�wt�̬�i��)n` ��㔥LV�{�U��;�n�X�=�'���YA*�cÆ�ɺu�܅�J��C�?e�kkMl΂�%��k�=�ٽ9�[�,Z����Av�فL�c-`x�2�iv;�9�<a�����d��X��L�9va͍���-Q��சS����9��M�v�m:��fۢ\�����h��W_+�1F�8��)`I��قӹl?��򡰔�Ky,V-=]T��B��Lw�a,���2�����v!��x��1öӤnoos</yU�+B�r����	���!��1%�
EjB�-�<��P����p�8�<y�b ����?c��SU��ǋ66N0Y��i��t��}}N�+\l�"�YKm;�*C���k�V���m^JEe[Fyl�1��Ù��8��.�DN��ʻc�/��_.CV�͹�۩i���	�t&ʰ�sv����KP�yy�M��l��"s2����Z\�hFt�[�����0X	�`�:ꇭ�7�0�՛A���·�·o	�Ee�4+d��m�1�d=��G�kB�ꕌ�&�Y��C�c��v��j18vME1���tn���&����`�n�4���
��5b��fP���uZ��k[��߮+����}�_�ߴ�}HR�[,��d�u���R�^�h�Y�l�,�t�m�V�࢐�K�+�jJ�炘�yjH����F�]K�#%C<�Sse��F�R�ք�z{��m�9�Lh�vA��rv�f:!j�$<4 cF��ӌ�v��u�lp�W��A��eהc>d�_�x�D�k̳���h]�c���h30�0G+,ۯm���H��J�/�$��X���:�ڥ����jS�;8��
MnF�=;\�N(�7Kl�6�h0���aJYY}�&��(Z�ˣ��6�BSj����7E ��Ϡ�(��tU��܊uѹ�c�W��.enL�:��qҬvu�R��T���؂�Nߐ <�mIqR�o]�;`�U��c���X��w78�Ho�Wil�^�uw��WU�FN�B<��+.��,K{�7VR�;zxwc�Mk�尭�*xj6�[�" ���Y>8�nR���U�P�dmM��Cz'b]h �+n��<���{'��F@�z�X�Q�����N�ʞ��+��Łs\tL�)n,��T�������X7{7�~����<�������e8Gj�&ad���&S;�t}.αB�ҕ��;9�[�rp����k,��0�O�.��M�o`Wz�*�� �+ҙ��=�d30,�m�!QOY� ܬ5}7���)u�����F�.�V8��bۺ�Nm�ɵ��0`i�ӛJ\�w��ٯ!J��i�o���s�8���v ��-�U=��꺆��Mm)���D���:# ����k�f�E�
v$�&�T/#�s��l<�T��(�t#W>�W��,�d����ɼ��x�u�dޠڦ�J�)��2��*H�P�w�Lt ������w_5�����E�9'fT7*YŰK��u���/�J�\^Ww�yh�=9LS9cR��|�H��_PM�Ou����b�����ܩ�콶��/�9��]e(�xT�FET5*��Tj�eaa;�1��H
� %PG�\l�->z�9�k�ہ�rJ�ޚ�wv����J�T��o/�n�^W�pܨ�Q�l�^�evW^��r{RW.��4T&Ɛ\��7�feֹq�n���Bi�'5ی#��%Ƹ��oCCE�/;bQ�rm���es��; .�ua��-�-8)�E��9w/�J�U�58@p��PU�V5��W]����Z$j�OkP}Ȳ˨�,R[��T��ռ�ܲ6,�<�U�r$04��p΢p��i�gfj*R�(6�R��Ҷ����F��(ZU[B��"�UiZ�PTF"�U����j(�2��Zª""[Z�im�Z��[X[KKHʬ���-m[DT���Tc-����AQe�Z�0QR�@`�[X���h(�ň��cQ-A-��Q��FE�T�V�ъ��Fն�ҫm�R����iZJʖ6+-
�F���J6��T�jKelDj�b�����J�ŋ�DZ� �%-E#i*ʖ�ʨ��6����*�X�ԥ�(�Ȉ""�Q�D�5�6�Q��J�+E�ڪ(�����Km��B��*�-
�m�V*�(�5-�b��1T�Q��-J+5m��j ���h*(#��b1UP�+J��X�ZX������*�m(���T�[*�jU�PJZ���-�e�҃mQJV�T`�X�\&��[?x�e��F��ǎ�;1�y̌�q
��Lj�u8�VQ��O_I�����;�뮖p�6ٕ;��]ow-z���:�|�Q0ˇ�>�p��٦����]�r"���L�B��?�������ܺ�ǟ[���{
Τ]]��p���9��D^�ؽ��'-�A�:�W���^�3/�qϯ!M8��E���b�btPM�5.lF�#/ԫ%j��p��T��غ`��Е�.�^C��c��4��;��b󺯱*V��+��Y�Ya�pt(�z}U��2]{5����O<��9�e���̉ի������C7Ѯxq��{"^X�D�}����CJ�<P�����ٛM��;���]����w��8�s���Z�m,��g��+����z֍���U�\�oؚ��owfΧ�u��I�*k��<����IU��ց�R魔(^6+�\�Ǖe����4�্��7bga��v.tC`��Է�g�A���u��$SN�(_'�I�N��>�{�{eo�g�$���}��W>�|���D襎�T�:nZ�V+�Xa�x�_|�{�ح���]�gF�3[Pgu�.�B�S(�9hED�f��q7{�����I�:��3����1u.��w�RS�{��ʖV�Ĝ�Y�;�s�E5;M�>���V�S�[ު�̯Q7@ܺ�:�ҁ�N/��!�O��{Cy�o��mS�KyA[�'�i�E�cco�D�,��"����e���9�b��wf�]�ɍcy9��+�;:�bs�v�x�@��\�t�%t�x��ެ�׆p����5��8���p����D#���-ᴨv{�Ɋ_�k"y5����K�9U���9,�m�o�ם7ua��X�"Sh�[�&5m�u�-� ����V�N��Π����u_�������i��}o)��B�˗|�,�n
���[�Vճ+ ��X�sywԎC�f��*e{�{0�o/>}l�?c�n�U�ګ�c�ax"�[g/�]݌#:($�Ld�;�h�\:��m��B�&n�*���Iݡ��4��>lCI�A�[�d��{�|6�ב�s�ԡ(%M�ͻ�*��]7 4K�+[2�b�kr&�k�/�j]�_��~ r�����3U\�*=���9��SĶ^u<t��36�~(���S��*Gi�:.OE�t�$�w�b�����r-�s�4��'�������Ƅ�X�<X���&-t�Y0K:�~�T�ے��F�y�����C���O+7%�3X�*��U�R�G���n��*��(d���n&���M��jK=���+=��deN� 0�K�yT^D�j�����[�β�MF�]؈�n"�:�ȧz���'K7l[�Z^�6�L4.[�{'2�7��}l>�J�uE�{=Uy]����m5��o����Xg�}��E���Q�NWo�����K8r�v��)�	�����y�Y�/,'R�[�������_�>�H�=,_5���o]��oa�[�=I�uM^ �́�����u���sn����k��d�k�]��1����wj�ށ�ܫ�����g����WJ���G%ػ9K��Q�3�F���Gݙٹ:���w{Hc��SY�[2��Oqw	LS�m,�:�j������Iс�����P+uŇU�-��j
�Z�_����*�o��٣���<��z��/Jזlq���3J�ҙ�c���<���܏F��e	$�]j�cm.�ɴ�z&ʃWXw���i��:��m�� �ʓ��.�������+u^saW��'�tI[�^��-�f�J��j�yŧ�iQ���}���|1e��pr�#f'ڣb|V��%k]L�侅6�օRR���:E�*�[��2�&�M�y��Qf���a�C�f�3�^J���)��˵T/�͚n�L,��1��Ӿك����&�_L�H�=�!� ���w"�ڱ�.�oi��_zs�a����^�r'7��{Sjg)�,v�47��/d}ybiV�2Pη�y�Q4!X�LZ�Ye��#��qn��ߌ�'���ʾ^�{ڇU[AKaB�}q��뻊\�Ͷ�]k�U���P���K5;�Ǜ3׽T
ȚnL�����c�kP׫E�ܔ����gG)�\��ƚܦ�J��+�Yg%��%t�^��\mۣ��)�l:bw���p��	��|�`��oҰ��L��˼��;B�C3ȱG�0�7j��su�ߞ5ƞw.̝�O�f��s)�Q:�|��%aA�3qʬcY�\��U����酺Im� ����:�����YY����ba�'1K���kK�����Ft�Iǽ9��(~����mn�U����KUů�]�l4j�/WXJK�T�'/��Y
R|�>H=��d�VZ�y����<�хn����!��u�o�j�%�W��Me�����f�UN]�J+A�tum��7��U�� ���;^[G�,P/z�r�Ӱ��9;�{/��ܴ���]^��u�j�;��>��
��D�!o@為�v�Q���ښ�Ŏ
��8v��Y���U�}I�z�"y��n	9��L!�K�v��}��O/��f�����E��J�)y�ͅIኌ�ޥ�U�Xٞ]���C;nk���S��������2����	�L�\p�<�S3LM�s��!o�j~��Q��y�^#͖�ٛ���;�t�D�2�b��Z�62���|����Q���W�.���4"aPF3��cU�-�Y(C�j�A+[�cdc�5�xq��zV`��^��ka`*�ʊa�+��lGΒr�d�X��$!������jk͢��T�';;'j��X�.�5k���"�m����)�;O�p\R���t��{�G�tMږ��>�ar�1[��6a�
��\���.:c{_9"T���m��ٕ�v`��e�q��w�1�ԄM��@'kb�<�לkذ���y"�.�c�k_k*l���������^i�\�K����+v�Z��y�c^�ȧT2�X%����]�����[�n��cb��W�*�	5�1��<�e7�6�Ɏ��g���o���k���|��,y�7�q�]��;q��=�a��h��[�۶%f.�QEi:�JN��G ��3]\������iܩ��v-�x�Le���ʢuW��Q]
M.���
��Y/Е����5������-c�y�NK7ۍ�fp͗�7�X̂v� �Ƕ:r�����m�MU�y쑜��w�2�>S*�iꦁ�N�7����]�J���t�47un��r��Nf,�]��ty�w2�$Q!��D��Q�B�������"�����~�����l!��ܨ&��]IŽ-���Y\��z�x�ӝ4���C��#�7�i����1T?.n8ޝ�s���֪��tz��r���ȳ:c;0E���fP��K�5vwU�sȕ�%��p�-�k�ݗ�kW�S����	��b}�R�7z�L�RY���Xڝ�s�<5�T���/>�h��n�FNj�x
��9p6c��d�Y]v��]OøN��k��6bF�ۅ���t8�Q�����]�6�=��wJ,CϺ�FP�&�	�N��G:��+o,O<�J��`2�(��܊5��u�W�昜hD�Ф�خc$'tyٷ�*��0V�n]�t�MS�g:��%g<��b$Z}��|���N�����J[����XztU�۴e`�d��P���1����n�{�}:�]����c��{3�/*�Y�z�P�xЯer�:�-]����o�yѴ�d���+���wnK7o����ޗB�j�ȑHօ^'M��vR������vټ�yR�K�4���J�Ģn,� ���"r�eVwVŃ]b��l��=I�z�p�0�[{:�{�+
��J��N�0��JS�$cC���sʊ�M����]"ժM6;"Խ���4�֏xY�<��j���툜���
x�:�kE��M`��J[���b���m"�Jwg��=�9]}�3E��X�j�Brr�Q���Nnby�l�n��7{�z�33�j��>y9�V�K�������;aJ���!>V�y�a�	�g^��^Nǣn�<�K�A�����˖��N痈%{ӾT����m\����3!���[����
Ŋ/z�r��R�\�]}���<�7�
��R�W�v�^>Rq����I��v��f�
k���fe�-��G^���&ţ��C{�ɓ������������v!O�&k���=�}��}��{��^�qU�{�2o`
[V̬mΎ�ӛ���6$�s(�qsU[W�vb�zuO([��e���#(W�E&����a0�ΊS�	\<�~��<��'���kuTwΤ�u-��٦�����b����T�Ȍ�����G5��Y�U*�У�r�|U�2]ױ[�D�O��1Rx̲�9�c�Nv�M�}%55�S�^5]E���W�\�y]<3*~�>�X M�(lYP��0�	�č��p����T]��+o�r�矲J��+ �t%�p�oJ����&��R|l�S;ˮ����Ӳ�"%)����s�hK��W\�6H������+W�L��wǸ���$�3�[ޒ�#.���A4[ڝ�x��I�/f�~�&�`uX�fk��X�iH��2sr���vg;�mC����v�.�V�[cؚ���nRͤ�^t�f�+�������[S���n#��(^7:��Yk��ƚ�os�fR�5k��)��:�����=�w��y���b��Q^ĝ�؄�c圩�ӻvnE�_5�a�+��nԛp㲼r] N�J"���J)d)I�_%�lsB�ýђ�yL�u09s����D=U�s���{B��]���7�Ry�F_5w�ΥL�;�W�.����h�C��k��k��ֆ���n����O��/�C-n��[�SηVZjW�aT�ȱ@�v��W�ޅ!���I\>��5;��X��y��u_��Rx=�$e���^�L�����౽����7�WB�[>�O{<Vu"��4���S�n�t������ͦ�0Ԗ��5�R�$�(J���<k��k۵0�c���[��ǻ#���}rʱ������n����W��Й���ey�]�]7��*}�m��uc��f�b�wa�έ6h���h58���!ʞ�&���u1��O^K���s�	���RZ����/d^GM8��Z�z�������u�ޤ,.���V�A4��{��,Y��=�Mv�}u,y�|B����:x%�T�,nv�*�Z��o�I�'t�Y���\.��N@��V3%�z�4k�Qn�N��5�h�0������~�6j�����J/*�s�q�
-n�θ���l��(?�t7��O�Bv�/�m?(7��,���
��Ÿ{4��t�])���3e��Y�ζ�5n��Y���ҋ^�D�<�Ӆ��@�Uw�{*D���B���9M��4֍ǛC��]荥�Q�$}=�g{���X�B�#)�B������8�g�tގ�*��,�٨�����g������]o�:�s�u,�����P�Rj��!x�w�&5��݆Z�af�M�.˨�܆V���<�6Z����F���Rhd���s'�w�݁EQ˺��n�e�)���$F�ҩ�淒�
�v�1W�5-w�fC�V�b�:��a.�,�"�%OBޜ��gG� ���+Gj�[1h0k�ed`�G>n��RΪ��U�z�32�jR�RV�[���.�ϴ2%#��s���]���fιW����>�zb<.��YD�Dpݧ�;j��A��[畇�19�E�6F�s�`M��ⴺH��Z^��ݣJ5.R	�Y�L�{�N�V�D�qP�:�u����5��Wt�ٺ�ӣ�<��.��'��N�1\�^�GY���۱�t'�5j�U�J%�̉!�������(ƶ��muuuG`�G����q��|.Z��gk�j�z�N��ji7.�\�S&i���&�X�7�ܳ�]9Co��:�ZoM���xa�.j%�~5�O��	�S4`���
�RՂb�܊3�2Y�3]B���b�ș\<����.����*yS0U��(-�k��ܨ���eF�=FԽ���eu��{Om��c��Z����,�9����ں����B���w��3�:ˋS�4v�q�^�؊�W9)�Z�����0nk�%	���~�@�U:�#���!Q%Kq��ѐJy��еN��:��
�����2�c'q�F�ۙ���}]	��[����M��O���`mN��1 |rr�R�\�Y��3ux�lү�F�]�dhm���1L�/�������q�����^ˡ�{y_Q�M>9]3�%7y<�����.����5�3>k�`�����y�)e�ݕ�S�4����#P�{�f�D�l���Xq���`������u�ڝ.���֏>�ke��ۃ��7]�����C7ǩO�z�0j
Be�Й��9�Z�j��#�پݘЂ��隗 ���5}�G�A�����9�Z,�6;J���2��=�E��&=��NA)�^DՕ�V3H[�m�y��^WL��kYu���B��bS]��RfJ�^�̓mkʻ5/.��pD�6�Gy�uhܙ��)@�{��U�ci��u{bY�Z�1oN9N��:�ŷ[�uu��d�/	�ꍞw;N��67@)�4�4�vX�Ơ�+�iv���f[m���lU�=6z�v��Z0Z�,o�C�\&�
VFE��a���J���[N�y��y-�k��̡�ᬕ���V����ϋ�Yԛ�pٌ��l����%H���*����gr�aTS]0�'�S3�2.s���1q*!2ᅼ���x�V�l�l����Y;���9qpyk0�awoM��3]����N�st �o�x�ȑk��Mrܙ�f�����I�q��NY���͌�\)��<Q9f�����Խ�ҏ�T�CW��Y�И;zLu�騩�t8X\o\mf���N���m.�T9oQ�a�i�Ӗ��}�>�d�
��w�}�'��vy�����s����*1V"*��mmAm��ĶX��1`�����B�P�YT�Q"��Z"��iTI%)R"�ҥm+m�A����%��UmQ)F	Z-lQ�����X���h�(��jQTU�-(�**����hъ[`�����TTKh�eJ���PX"�+Eb��(��+QDKT,E�*�ڈ���jTBڪ1F�T�DU���X¥UXT� ��-(�[[dX�eTc�����1�
�(�JQ�mE�*�F1DR�(V���,U* �l��DUQ�����Fڂ��EiV���"ZQUle-���E���l(�E-�(��h�������[X�U[k��DE��R�0�Q1��
1Y��h��[(ʹ����j�AXe�"��W,�XTQEUE-Z+l��UAkZ�/߾�}�����c!	1a�}j�wdҭ���k�q�)�����[v��Z���0�2�0%7\��}��Oe�ג)֖�Uʊ�k�X[
B�����;:�as�v�,Q{�g1J�wy�i���σYN�`���r�ǝסs�a+ޝT���&���=A�sȌS���KC�ܻͥ���Pq��鮕@��_#m��My�wV�d��J��X��H��x�����	���/s������1�^q�U���]җ��g#5�Ul۷^bv#@>,�S]]M���Wٳw�T2Hg����DVb]�/Wo��M�4lƨ�µ�	]>��Ʒ�K��Z����!V��s��ܚ�3(&Ld�;�~G::�me��RsFDfT�sYc
x���3���^#��JM
�alW1��Ѡ9��7x�q�|���L�ڱ:g:��K��@o1�F��l_1��*y�jZ*���T��q���bÓ^�y1�j��KVl��O1��MF�)k!]Nr��ю�
���NQ��ϝ w��+#�]b�r��L�FUm���ݼ([��lRU�@���r�sZ�{�ۮ੓]\PWe�Ic\�e�:��%#2YY̜���k�n����X�jDfc�.y��S����цs�xL���j)ju3���[��Y��Ύ�#5"�P�ƅ�Yછ��S�\_M����w݋�	��w<6&��I_ei[��6P���Zj�sc<����w�ܫ���*)R���i����L��C^��]k����f��g���v��wc�_.��j*�tS�p��{����9�v�\�����#��I������2u����D�5�ar���	�������da��:Wk��g�J�,��͆lq}Ĺ�����5��2����/�Z�۵�	���'�f^�#��:���s>�R�?Yr<�#��ddj��U�{*^<RmK�V�Վ���F4����lʽ���j18«��7m�B�Ze�W�盞v�ӝ�
��(>,�S]X��X�8��%{s�;z꽇*��Q^���yЩ���u�ç����z,��t�;�����.�Y*�z�F��	쎹��w�ה"�5u+�!�q���=��^�uc��3�Ь�hv�Ϛ���{�J�L�wҢ�@���᱁��P�Th��o^5���lK�ס�ȹ�7:�2=����k��K��ķ�v��N9���zD�w�f�g�8�]b�q�����}h��Z)7��38a-�����X�:D�h��˗)M�*�uW���9�A�B�`��C7�]��_��Ut+�̬�C�������.U�S�c2]ױ@o!�RN@��	T�����\W������!{>�ח�"�Z�(_#��/��3�R�oM����r�x`��{���ͪb�,{)23�gFkf^8�{�F�v&2i�s�QV��y��m�kޙ���W=�"\ǝ5M�y�ˀ��|�z���]r�yVZ��4��{�%f#j��;���JKSV9�^��5L��0D�b������؄�X��S�\�3�fL&�[�Ng{"��T�V�}��82���S^Xq���8���=��N2q*js쐬�a��0�I��z��w��MvW�yAa@�GG��� ��d��&�M���|�u �����!�>I�l2�$��S����n���M��<��:���y�^���𲶄��&#;C
yP$ܠ3h#<�Q]��{	��v����(��I,�u/�u���ެ="�n��r���
*!j�r��\�bg4s\�V+��h�D�a�glR̥U�/�@�����A,'�V���]�z4��\R�Z��`�_+�ۙ������u9��������������N��I��'?w��MN���bI����I�6�~-:�d�Hm̝Mad�a�y�O�(#��F�k�?,��[wzU�ͤ_�ĜՐ�h~d�'_P���XCG~�oO5�a�'猟0�>w!8�d�w����k��䘂��t��h, ��K��ѓ�*Wӻ��U9k��&0�wT:�I���w�!��8��l>�́��h�p�ğ$���}�:�d�'��!6�$��~�I��m{� D�;�@�6�!�ݪ��O}���㸒��*J���d�w	�O��T6�I���+�!���@�O��}3��z���M0���$�i�pG�;�=��=��x�O�f����q�tI�����1*I�봕&�Y<�N�~d���	������m���ԕ�����8�bu���=Iԓo�&EG��à��\�l�L�^l��%�P�'�,�����4o�|4�8��g�I�RO?^$�����Rq��'_P�`m<����	����%zɤ5�.=�Lc~��U�Owl��n}���$�	��sxi��\�AC���Y���'̜��u�/�&:d��7�,����)8ɴ��'�P�`u<�����p=(^w"���������}�
m��>��$�T:}�8��*y9�:����Rq'�T=�p���'��0������c�$�����Ð P=���/���to���YԨ}��L�'�8�����N ��o	>C�h?o��J�{�:ɴ�Ms�=Iğ�P��r̟�4~��m$�}Ϩzcc����)��7A�}��-��Ds�Ka���8��x��O�S�x��I����2q�����8��7���I����:�ĨO{f�u��?w�_�u���X���c��.�aiv�r�2�z��[��0G���74��A��m���Z�<O��#G�A�ϒչ9�ڱD�'��~��N<�-ޔ��g+���s+;RT�6�|�.�9{�f�P���Y�.�����VA�x�+�����v¸�7�{�D�n�u_��}���`�?xN�0�&�l�O]�i4e�d�%g��ԜBxj�8�ɯl�!�N��yBm'�3y8�g�����=��y���o>��y1�u��z�|���'�Mr���@���Oϡ�~��S��O�$�O��'��'SFY�I�*xj�Y&��d�&���IĝeMsq'X}�޽>s�Ӟk�j�Ϊ󭫟�����<>.G��(����d�O�>��I��?9�p��Ӕ6���PіC�񓉣)���MO(q�a��2u+����7��y�ə��|��e^Ws�(p=����}
��o�u�I��̝I����r|�d��rN��Mg}�LIԆ�C�+'�!XC8�Ld���w������w��j���ǰ��I��(q�iX{I��d��9��VN0��p����&�̝I��'��d���'�����6�9�y&$�CE��VM�����w������^������=N�1��N�0�c$�P�&�2%��M�w���HVN0���i'��9�:��$�5�#�p.=�-�	�{�=��g��W��"3���?f���}��w��'}��+'�,<-�?$�(�m'�Xm<a8�L�������d�O]���0��a��ͼI<d��a:βz�N��k����ʹ��>=��sss�3���G��v������	�(O7g��J��P8��M�F��O5a���g������CW�`u'���g0��&�;�����}��C7w�}��=�� ������x[�=��CL���$��&%a>����iY<�@�Ơ�<��d���u�'���̆�kg���?}�T����j�u#��C���
=�?N�<d�O���? �\�Hu̝�`,'Rr�$ĩ'���
���Yd�'�N�La8ɶf�5��ߝ��3?vAc�E����=�cUuެƌ/�����X��	n�6x�F��k8�Q��)ׄ�s�.��͡�m�Ȏ��W$��%�:�5n���$:�Α;������v��-��P�\��`ПMr��֦ �oQ�P] �8��Q��Q��[����:�ڢ���LLN!��é+��a�~ͲLJ���0�$�[1'R킆�>Ag	��'�9�d�$�N_rLJ�uٺE�q� ܫ����[�Β���{�*>��=�I�I�M�q�՚~I8���=g4��^�LJ���È,���I��;`��O������$��}�i���S��)������*~��{��Ϣ����,8��O_�������u�Ĝa����'P��y�����è,�����m+!�w�d��}\��)?я-[Y�m_��~��
��;��5$�O��$����vE'��C�Rz�=�Xi�OS��8���'�<d��ׄ���9�:��{�sJ�W}?NP�ڲ�_j�Ïy@1!�|����O����'�M���ԓ5�~�Ol�M?$�e�d�%O5a�a4�3q��'�u���5���T�m���a_d���3x{`������i$�r�d�VC��Ì�d��'��=d�'��w����5��'�N��l���ɤ�2�2O����!=���Y�w>���W,Q�@� ��>C�'��km'�f��4�q���d��	�� u&ߒrk�'XI��yϼ$����8��Ğ�Yd=�T{�@��"�\U7�|��|��}�� ��u$�/�6�Ԭ�m�8����q'P�s'wd�a�ì�~a=�r|�'�;�u��'���}��8��v}7g?��k#k�T|@1�TTJ�����SN��k�Aa6�jÌ�J���M��'��s�HVN!��rw��u�����ē��rR|��-���A�S���k��=L��zc�i;��y&0��h�6ʓh,<-!�?2q5��i8���:�M��6����8ɶN�!��2Ad�{��
��+���ߏ����B ����/�{D������@��k�_?R�{`�[�^�Ngl�֌�Fk�"�\�a4�*�~U���=��l�o!����/%F+2R�u��4t�q���=y@���>ŋ�Q��"�ʻUb��f�;OD��-g;�� x3=�����d��I��'�9	�m�G{�1�~N~�$�'۳�T�AI������0�M��i�N3��M��5w�� 8Q��P�Dn}�sWv��_x	�����x�x��Y:�d�M?��B~f�4o�ya:���^I�(M��VM�d�(a��i�,�i:�MXn�'j�Mtsy������>c�q�<!d@�O^!�9�>`|�\�m�'�? };�I��&�i�N��'���C��$�'��ԕ�iY<�@�̛�����j��o�͝�fwc���(��Ƕ�I�y5C�+�!���N�8��>��=I�I�N�<d����	�i&�Y�u�:��N��9u��VMb�õ����>�r��q���{ ��e'�OY:���XN�~O'�4��u{C�+�	���	�������M�ˇ��AHs�
I�?�����f�SuU�ٻM��{����hzYXM��H�m�̤��>&�,��O=��䓈h=�=N�i��~�$�ʇ��������p�'Rk˒6'��ҟ����<���� �@0�{��̞o~�i�q'�ϼ�=�N���d���Xq����'�Y0=O5COY=ağ0=Ld�~�a>B���?o���}�UM�Ld��}y���O�p@�����8��!��d�'?%a�7� �������̓4��I�Y'_yH�����-�XI��{�$�	��1���<!���S��y�)�.���^��	>C�4~�Aa?3�YԜed5�4�l�%a��=d������d�ɯ������x�7H�����a>gQ����������w�k�;
�l'f��x���^�>C�8���a'�q��o��'�z}̝I�VC�ӌ�d���f��|��&�;��a?0=���o�'�S���6�O���Ng��W�VV_:��=gzA��ꆯ�����CZ��q ����5U��!�&�[)h�J���]�Y�=$%oO�<�'��(����f'"��h�l���
X��1�}b������m�3[x��.Pj��X��ͺΙV�W���]�u�X���2x��P�I�*xj�����d�'��>C��J�>�Bm�]Ӊ�$�����N~���w2u���v���tl︌���b��7�sg�|�О�;�N8ɦ!�Y��N2�l&Щ�jÈ)&y���A@���i8�ĩ����a���I�/0�=������wW�qY�ekȟ�����O�6���s$��Oϧ���q!��m+&�|��Y��N2��~C�La�n�aĝe`x{a��d�T�g�=�+c[�~5?
��f�m���$�æ�$�����I�����$�	�^�$�H}l?%d�����C�N3Yq�~C��,:�2M�� yG�x�þ����ݮ���9N��rH�i���?3����xs�6�a<d��aԛx�z~�,'l���|&$������La�AN�Y6���i�����$�2�ӹm߹��Mk�uׁSL�׹a�M�d5hq���}C�~�`u��a<d��a�'猟0�>�;��M2jwxLa8��k�1	�8 Ǽ���w���7�S1��<ީ��I���fI�f��Y'S�V�;��wC��I��d�C���$�'���$�i�l4�����f��m�{��uWCux�b�2~��w�y˻�1	�~�$�>eIP:��'�,'Y?3Hu�����+�!�}�':��́�	��:ɦ�3�8�@�Ϗ(��K��Je��vo�|�q���bT��w�*M��T�d�ɷ����q�y=��XM�����̇�~���4sr2���(7�VRYz1��g][�g���Q t7������Y�s��~d��=��$�g3�$ĩ'��ĕ�~��N2~d��(N06�Ohi���P��}�@�
��yV0}�=[S=r��m\O>#;~��#����س����Y���]*��6���hJ�cK|��s��b�ͻ2
����'0��ڑ��$Inj��y�dۼ�Z�㬭��o�����n.���e'z���� w�q����|�{Z88�4<=�Q8�ɫi�ޏ{� Ǉq�<&&�O6���Nw ��O�,����2xs��i�u��ϼ�Y'wdY7���'�}M�P�`u:{��������k��~�n]���c�8�䝛�>O:����d�ʇ�o �J��:���wԜI��w� ����}�|4�c&����c�$�y"����ۼ��lw݇��/rU�ﮜ}��P=qq��u��)�6ɦI���.����!�4~�Ad�<=�d�T';f�q'̨~��@���&�w�6�bW�{pb�?J��}�%K.��Mχ�	�tݑI���l?0������8��=f2u�Rl���8��>�z����u4�?3߹�Y8�	�l�{���H���D�|n��r-���z[��u?@�O;���'�����m��5=�)=vɤіq�|��C�8�����M�d��u����I�4��ǽ�'c'\��uwq��d��RX�&�0��6ɶM�I�,Y>I���~��G�p��I��2�>Ld�~�8�>eOP�$�?`u��,�=��y����:�rj�W}Ծ��&����jO�;�É��=�Ì�~a=�p�'R~x��5ܓ��~s��'��Cl��0�L����J��~C��q�{��Y����ɘu��%ZG�bOԜIĝeMw쐬�a�y�]��a��d�N?0���8���'���:�u5���1'R���VO�>B�:�Ǽ�J����3N[����a��{� Rw�������:����&�q��P���B�q�����Oh�2u&�0���2�|�����1�m59�y&$�<:i��mOONƾ�t���x��l c޸�`m2q;2��q&�^Xm<d�u�8ɷ�CR��&�;�y�$+'y9�~v�xɣ�é?;I�O_�w	9�ލB.>�>b�3�m�Vi��L��#���-��f��f��2�e�NV�&��^��7^;�M�_Z�&���@t��d��e,��
Y�lx�!D���i�3�})k䮍��Z�v�<�GPWl���L�⣹Ú��Ehk����`����4v�*g����u�on�;4~���q����" �u�B�m���ğ�u��RM��i��N3�������d�O]���a�:�G{�x�x�g�~����s]f�-L���?dyG�q�q��H���z��d�C]����'�vq
ɴ���?$�(�q���Xm�'����Ǽ,���P��ekϋ��߽��Hc	��?2x�H7�'Y�M�����i�G|��Y'�}�1+	�u�d�VO�q'�M�M���@���xy��~�ߍ}.����>��+�C��a��ğ���9���$�Zc'|���r
2~Af�;�C�&���Iˬ�������� `I��{���FR��}H�P���y�N�q��Vi�I��é+�&�{��$Ĭ?M���$糷'�8���;�P�'�js�AI�Ow�&�N��9�y&%a:��y���l�t��<���w�_�k��oH�i��,��=I���yBml�Vi�$������C^��d����o �J�s�:��)�AC����Ѿ�'�=�5{�;�����#oK��������xzc��{{kޘԓ��vE'��&Xq����'��	�C<���M$��=f2uwz�|�a����$���0����zc���z�-�����ͭcջX�f���O�ږ��v�M)�Ռ�B��l���oբ���^��C�EZ����W<��gx^U�M`��b��53�)f6����.�P)VZME[O�)f������{���I5=��޲&��,��jT����"�a�S�wG:�2��<��N��n!~>��]Y�ߣ�[�Q��PF���M����xz2l_B�A�讪�X繘�P��oX9\X�j-ަ��u+�.�9��CvK�m\���p۠7'Wk�	;��H��`�w���
���*V{�M4�݈�Z��9%�Y�͡��D޽+��]�ǉ̋1��́�y���j��]GA�����	bs'*}w�HSG�J��
�9�`r���h.�9ҽ�u!R��[����0���;��Ԣ8 餅� �un\�5ԚT¦:�U�����ұ�ӨK�����*��� j������Ƞ-BR5s�gF�B�:����t�V%(lCX���`�x�FV(F���+�N�tl��p��!�0���[�k"ݻ��,=�{��+z�l���dQ�묜��@R=Z�b&�+�5̓Wd������7�����0,�C��ZZ%>�nG5���u�n]�2<��c��*o�ήm<�ޖ�_��d.t�fM��B��Wu'N��[V��3��:2�-$P/�k~�,@��7Yd,�ӯ�fP��L*�]�$$:'����v5c�o��<2�l�m��A�<F�(��`5�|�vEh��;"�X���e��N5+3��e	��w%�b^�ȷ�6�Mu;�zޚY��K��t�3�*y�)��Ј���ݯGilb9�o�;��Q}نI���d�p]mouj4]gQ쳘�{���i��6�����f�Z��ʒfPڏȡ�5i��ْ+�B�E�
�]"��E�#{T9����^���RJS40,�����!�p���AVrlvY����`�R�b%�Ck5�[�pS��hX=�M�8��Z����C���U���xM�.Y������hfIZ�_�j
�+�p�%'S�>OQ�S?ϰ���åg�
��8��*��r؁�a*����'Vj�X�#ZmjQt�k}4!�n;C�l\��6����턢�ݧ��v��u�X7[��}S��+�� ]v��^!\�pXw�m�]�8'>ȔܔOW[�kX�T[�T�ٹ���yyf={��)�I�tab��%�-�|+r.[��95f�h=�t*+o���u�Q���ls�j�����f%��X��7)�ָ'�ݝa
l�핅����%���L�!Xpl��\%����ڵs.�{��(ý�U��[�u�N�f7M;[�(Lޠ6����[�;@��+'w������I��D��@��lB����'j�%p{OI�]٘��"ٯTv:TL�w=�/�ɼnJ�}���Z��>v�ة�ů#��3��Ǝ�O�-i5B�(�؟������5g�ݥ���ꆃ!E�)h��!�Oј�^Nu���ݶpse>*q���:��wԻ�u��Ki����jj���]
�MU����X����siJZ�Ѳ��"�不elEkQ+A�(���eT��@�X����1iD��TEQQ
����KJ�-���BQQF�k\���%lR*�[b��Q�Ae�P����б�U��TPb$QE�����TD�@R�1��+H,�PdcYm(�(VT�Ƥ�[h��j��"���eX(ւKZҬPQ�����dUPV#mTQ-�%�X6��ң�QQQml�"��)mb�AEjUTU����S�TE�X"Ȍ[J-J�dX��VڌTQ����R,[j�`���bƊ�lQV6�AJր�0QʠS"����Ub1�b�X�����R�J�b���#l(�����4��FE��
�V�a�9l�Q��� ��F�DX��¬Q`�hUA A�C�}�p���gv����U6�9�VV�If�^n4�d��՝�O1�F0�a�5�v�]c;з�[�V��o�����U�d����@��HW���W:�+�}��kr��*�!V`wz:���zV���j�S��_%-'	��Bk,=�����[��rs2�aqX��N1;(.��BX��7�e����'���ꨭz��8ʞ��G��:�X,�_��I����>��,b	r�*b+��Ie�m�=�U^�����f��-���>,Q{�9MF�	�yO,߶"�ڝ�G���o����r����{\��{DO(�V�x�de�!�����Z����}9� �s�t�i�u^l$��^X��d��yj�}i��5,	�"�����O{<U�a�X۝=�6�us9|��/o_(����A=uu�@z�����E���4&�<�3Q�1����(Î�9�~�Q��ds��;-Z�(r����8�ܤI�"Z̰Y����Cd^�W�F���:���}�g�=�lP�`�e]vV3d�
R��9I�7sB�^��-治���k_ӻh֜��	��bJ�D��GƲ�w��x�4Z��{@�g����Ӫ�<�k�p1��\G%�S���� zd'm�Y����xn�B�;�a6�uBھ���T�X̗�isn� Z��2��w1|�Rv�/���zhsÍ
݇׆S"3-U��"%�Z6W5���t7����U�[��ߌ���oҊ�u�� ��\�CN��t�Ւ��b��R�[~��[Or��	��}Txs*L�m����}Q�fʮͻ�й�n��d�c-��{}7}�OV�dd;�k{�'-�9������Y^��HX�l_%���6�ʽ��u�{�؟c������T�/��	C�8�|�l����y5r�,���n�|�ü�>J���FƉ��n{'?$m�Y>�鞂n���t?_s�aO���$�^�����h�q��cr[�Bۭ����K�g��r��g�s�[y�y�������V����I��n��e���U2��>rf�nS�X�q�N����v���O�st���rF����&��	������ܓ���e�y���epZI)��E�圴��anjy���+vQsV��7nmsS��"b�Ҿ�zqE�Ÿbֳ̩���{�QܱM5�2,}n�Gt�B�ה#��±������K�_hs���^>�8��x�|�f���!6����i��uB'�{O��o!��}����tv�7� ��U�9���ɚ�L�av	���9�}����>�/<A2��{���HN�	�����8buG]�kҺn�m^��w;���V�����jf'�3M�	��G1���Qf��r
�ŝ"�"���Q��/u;X�V�fJ���Ns)4('kb���wG��o�iı�����Xݍ�v�`����P������M��I�ؿs��"���䦫�q�ŌXrkE��;U{iMd�y��f�ֻ�|�3�����Z������]ٯ�r�<ٛ�
ȑMH҅^6+�\�6WT�x��8-u�<�ͽ瘖����4�˼�kv���X9.�
Ȥ�.��[�5N���=�����syV�`��^�����ѮJ2�m� ���s��ݡ�sAe�0�r��d�X��m�6;�_c��_p�i�N�S��k��B�)];�	�4�EV��^ue�k1 �V��Zo�xm!)zv�������  ���U^�'Z9lR���t�G>��i��S{�%fP]tʢu���u����\�����|�PY|��~E����m6�.�m�l-b��� fy���9����zz�}|�_��J�δ�>����{3,�p�tu���h�hdX`Gj�O*����w���y�eqs6�|�/=nȼi�7�}O=o6uU�}����_�!��UwQ�g`S��9썅b�C�R�X�җ�۫{T9�ol�Q���@���R+su�r��C)�m��U�\��b~/:�.��Uԩ�4;0������vS1��)��G6so��6�9����[m��I��6�1z�lg���f0n�{ܺ��p���uq���f'�ͫ�2�&���	�5�S�Y��-��Z�ϪR9A��cSU��v����"BM
	���vY�z�3� �a������+���6��e�K��x��e�۪�/�4�_Zbxm�����<��(R�V�E_B���N�a=J��t��]�$Q��o�u'��mX\�P��z*��P���e�˾�\[|5��F�kB�]]�&�'G��f�~� �Ь���R~�n�Z_^\���J�%�sء��)�z�{K=�^8����[���y��bq0�
�ߦ��VKW�(3�؁w��˴�����G[r��N��><������<ٚ�yTVE57�\��"Dfw8�ƞ�<bb�W*<�,����l����k&:���G:���R��)W�����6�'y���er�ʕ�>�	��)���d�T�\ŋ�ڽ�3�	{�{�hN�/��I�O��Me��uһȻw12v5���x�̔���
;+ǥ׉�R�O�tH�k��oX��ϡ#�.]差%�����'s�u����ϒrĹ��]k�C��w�ù�i9��j��g���iR޴�u�v�������v�x�u���>�����|k������l���h�Qр����[dE�,jආ6��fœ�Y��]2�v�&�'�n�[��k]��<Y|���F�^�擛9��YŚY��AR�KE����N�*[��N:�ned~�5����P)��W�FО�� �Իp�L�뺒E�H��E��b�jNr�W��~��=�7���T����?��9�w�Q�gg�Y��<��u_���:�$�!w�Skp���Ν��B>=�v��څ>���3S��U�l���n�X����^��r���]���#X�f�w��>�gUG���{zC�:����p�fݨ/�x���ǖ�׺n��7���o���O\��n�\/3�7$ޏ;o���y=ŏ.�	���HN��E�S]P�P����Skw��:*��J\�Gc��HD�|+��ر�l�49��h^ȇב0��잤�lF&�U�Y<����T7����P�kb��my��^$)������*qx�żk�e�J}Y(U�B��P\�lbj*�}�)co��������g���\��!����.m�&��](U�q^��@U�����ӑ�=��x��a{�^��K��()t
�H��_%1'��	X�P�m��\������w#��#�\��_\ȇ�~�/o������Ѯ�68��2M��V8'�)�\
�	�쒻_N�t c�$0�̻Q��mCۘok[L�uu��{��W#���Ʈg(e�=�t�^���q�7�< ������U��Uw�˲�.Z�S{��*�,�8�%�u��w�+g�s��S��r���>w�_+��y�%E�t#c|�a:�S��zd3!�]�f�b��etZj��aHW�4��z��{gim�q�xk#/�|쾞���	ܼ��7N{�ٝE�Ѕ��ko9O:�Yy������8:ŏ֥��C��"4����V~�<*J�e�{�3����o_V�Y5<웽��;����{0�U#"�O\���畾��h��w�����})*��2޺+��up�Ok�l*	�qў/zjVȼ��q�-�,b�Vq�c5x�p�y��yAY�LN�M�5-E��Q�@�sB���#}W���wNd)N��ƍ|�f��(��C��N��8m������{Zۛ�7sּo˼���*�s��
���I�^N��1���̉n��d�� ��޽&Ἵ*[*��� %B�ٖ���t\5�#I�����FVIvhؙ�����{�l-3���r����^QW_#���J�(�^'CU_T���}B't��a�<9|�wv���v#���@��	�� ���j�����B�.��dN:W�(g[�t��ӰK}���3ӹ�+֥�W�re��F����ɇ����Kw��C&�-��K���ĊM��w���#�3]��f�y�z��hX��dSX+�
��\�{�(u���xɛ��o5�򬴒��[��v�ݯm鬰r]�$
C�\�
jZS�Ԗ�n�8��J�����::v#�e��Ղ�ݰ%f.�QE	%�֌���}G)<�d��y�_%����-e���i���Uwwms�8w;�e޸��~*]_T���]|�XN�+��o�ӏޗS/��̽�˷�g��i_v��(�i9S�as����;���oWr����&Ld��G<o{��s��<N�m
(����[ް.w)�{�|��J���|�=�-71�SwW�{U�{dg(腽���Bgwc7�F�����-w��4�x���rz�jYJ�gXp��A�=ڽ-�{����"fi�G�c��H�:Z=B<����3X>��}�����2n�0Gr���f^Ȇ@�03�	k�i���3���**`�ZZ�;Of����6�fe_^31�]�؞~����nMrfn��_�,x
ί"��]V�L�Y����+zu�^`��k���KB4�ا#5��jٕ����O����/#T�9����lG}2b>��Rľ�u����z��ms2�&�	�5
��nU��Gr��X�Z���c_�[��.|�ɻ|%P�̹~h���=9~��yC��r�Op�nZ	�x��m�S{"�^��[e�.�M�Rx�x���vذm��E��:jLE�s+�x7����)�x>�Fu�8Ӷ*�Lf�x��=5l���
����gs �s#�hˡ�5�aw��+�z�y�w.xK�y3���ZxneF�8��bn����:�J�*�E�;
ʡ�؞wcqK�M�.7O[L�ذ��PԺJ��M&�V_{���Y�C�^X��T�{�KX< uV֎�-Uad'KNBei��cd�W�M+�h��2(��ޖ\�W�(_��z-z��
�L���[&�:p(��B��C�w��]h�=S>A��n�k��,�x ޕ���7�L��[��Y�Aj�0�.Ʃ�(�)Qƕ�h1��1Ѵ«�.nsF[ՕM�L����=2\YDf-`�u���Z�;�=���������� ���GEw��`���J�"B�9�����B{hd�}���*=*�3#w�z�gޥ�(��"���I��e��Q+�{���n*���D���QNQ�U��	��'j3�ĽS�sn��U�x�f�6�"ZD8�}}v�*�P�C����UY��,�i
������F<�f���g�ۈh���'%�GEGB
��M��R�YX/��|��"'�t��;/��v���:.V�v6͎Zi���Ԉ��tp�E��w*p]�z��kP\E��`C{*ӧzvT�m��sN<�dT[�vlX(.ʒg�Ai||Q8;yO*����A�|߆�T&��gf��u���o����9D㏨y�޳}�ܑ�^��)�`�Y�p�\�y��5թ���C�H{��.|��>�;�҅l�����)dh�
m|��UDq����[e��q���.c�f�1d�VV{��ٙ5zދ�_���1h�!�����Pv�]�g�IZ��yWJ�YjB�X��[iQ�K��y����W�O��లu�X����'M�c� {+��!��X�L�D}��WJ��;6Zd��p��/�X�aV���a�ޕՕ��4�H*��!P��uLw��`��^�������N�(���V��
��q'��YՈpX�v�cN(�ɭ%f����=�y�vA��k�J��.o0�Stj�+�]/e!���������}V��H���1Uu�9}�Vf�-*��sFf����w0��i<���V�|�o@���:�ݷk�*f%j�Eh �<n��3����8�7s.!�1���:�Ծ-�Gq-�5���Yƅ����Ӄ��%:8o�#:��9�\�I�F��v�3&r���=�Y��Ұ�j�	 S�o.�_��`��o�:�}/QY�g\K�:l�@�=ɱ��V�M��SZ���c�6�l*�K�:Z�\��S7�ˢ���J�����Wڷk�(q����r���P/��Wqz��p|�B� �m4�4�^g`��6�j8��ʹ���i��Suo|o {���V�#-Wu�o9d��p߉H��Yw�s#U���խ|�"4��5����-��¹�� �z�9Sdy���mFd�gIN����{��m<�!\��۳�Uu�X&�"���T��U<4��㤫���v���K��A�T��3su���ug�J�p�H�]�WqE��][جeYֻc]�u�V�mFl�KQIý.��483b��0/]2䣂EH��PD�,o�D'C�BB��Tc�u��8�C�g�K5�6"7���؟Z�I��z���/��iC.rXn��9�C�ܟ>���2>m˫���ϓ��6�*r�8��M]/Wh)����sE���3���'v��l�:���w�&�v��v����������ĺ[hm��#e�O�:��+e���bI	͹~ vV�̖2ЋV���B�Z�R��{�0I�Xvޞ;�VD�wm�άN��]Suou��
떕��+XVc�I��]���N���6�Lt�����1<5��9���J�u)�2��OT��ބ@�����v:���[��b�=�LAOL,9wv"�:y��<���ذ����N��Pu�\9����O�Sг�]������7� �j�4Z�Pdc~(�&җ�Z+f\U�)}w�l>�wN����H�z�2� w�Wm9�o���a�l��8�+��	F�j:x�|�}݀άv�g��.�\�;w�i��B�J="���i�&�y�ʉo��v�x�R-̈�Z�B���4�ǳ ���gL�IX�#Y�=�]Q���(O�&�&N�gR�+��d��^7ak�=D�^ܞ�I",�Vu�Z�!ۡ�R�QW�~�d���fU�d}�>C��w(Ρ��4�=�T)m��e5�N�-.�=��bJq��M�CbQ3h��c�T�Ft�ջ�yV�fps#o�V��V��P(_9ƺ���;��w��J�TŸ�`mb
ٙ[�Itܱ�9����'�[J��mQ����PH��T��ªUb*��dPF6�"�S,���q+Q�TEUk�PV"�Z�b"1��D�(����eb�+TE�����Uc�-���BҢ".Z��`�5���*#q�ň�b��[fZ�8,V�U�.5b�ڪEUj(���UQQ#��(��(("�m�(�Um�`**�ʶ��Qb+TX�D�%�´F*�U���1��L���W)ar�cUQ� �E�Ŋ"��EVZPQL�A�*�*+b
.Z��J*��%h&%UVDjTTVV�(V%��(* ����E�#�P�T[E��Rڈ���",Q,DUX�QDT�J��b*e��k��ZZV�b�Ō��qDTUP�V"�0DU��e((9j���[A\�V߼�~o�~����G
N��ɺꙧ��-s���U�-fS�v���ݞU�^��\�O,�`�f��]��3��}_UW�R��g�����D����߇a�}Cs�
u���N�61�3���ء�:�1=5iٝ(�𭔒��� ^���w�A����k�D��z{����Oo=û����;�U��=�<�މ�}�ӂgc�X�Y�M��VW����Lu	x���gz�k;��t�y��َ�.E>~���j���n\.�S��^�$hR�H@G�o_�uZz,�Õ���ƔU㈛V����ORe��d^>���y�n��Z�\2RXϥ"�E5ԫr�����-�%_2c�c
���m�QP�K�R���'ٶZ��xiŃ�x�.9�۞�Ve��+Xwԩ��)����e84 6Vd��uT��zą�١���x��Z��E�vw��[��Y�
�fĂ�Z����dP*y��D8u眰U���;�D8Tr\�8U'��p��a;WU�����܈�d��]L�P�zǪ%�L��O-N��u8�����a�w'x�g~�b6}Qoj�}�!�M,�5?
�W%���j�5���:=��.+��Tٮ�Y�76M�Ȕ�d\6D������2	u��Se'�aٽ�F���{���#vqg�ҩ���w����ab2����)���.E��3���P3�O791�Y���sphU��	�u���7w+�����u_m���ҁI�����2�s��� ��`�-�6nf+�z�F{�6ї\s��L0|{"��L�{S�c�ߓ��囏��9+�,�:�*wJ�"��f�����]Ʋp�,{�qޫ�<pJ�h�C���޺o6��T�?t���*�lKj������]	%qpn����a:�ئn��
r��̷���:����s����h���,=9%�o:�hjb���"�sh�9�a�r��!���L�nd��6�XV)�@^G���p���C���'تǝf� ]_? *�ի�5�Xvp���Ky��W��x���޽��Qa�k���4�zIl�l�!cn��q��7l⛽�甊���vb�<��q����F|��X1�nĺj�(�(Cֶ��"�t͊ך�_�]�B�+x�j�Ø+ݾ�y�6�~��E�j�v��2�Ij,5"��Mg*�Yj p`R��U�e��	����g�:Zq�5S����/ˤ�ʡ�1�&��лR�b�S�Ԓ��O�	��
��(f�:.��9��Z�܇sw8�{�� ;T� �&� z��9%�+���*����-q�O7��r�R��r�jTxܨ��7r35ؾ7͍(}��ߗJ���J[V�9|xռ�-oF�v��ȶ%b�o#�e,u3�?����S84��\ف֌�(���	�a���c3]]د/,!�:�!߇�< )��"�K'�ؕ5��B�3D�D�"���0�>�\�>R%B��<��!��2]�S19�,Zhq�C�<���OWz�3)JP�S��dS��0��2exof�qi+�[m��#g���sGP�����ۺ�F����9m�QQs���-PYϧ�.��YM$2�E��s[��+��n���.��Dq��VK�p!�a
�*'OK�^e�뢞8��/ܫ���8ե��V�Vo��Y��,�`��bG9<O`~���өi�e�>�X=4*tx���R�v3T61'�A�sb\M��Gnt��yֶQ�%�I��`S�E]WaY�<�mY��t�|��5L�����T�[� hoՕ/%���E��c�ÎԒ�Vw��7*�	�XP�B2���^o@6-\ۼ�����sn�7�1�{X�$ܔNX���O���<V+��|E}{B�gԹҧ����Jn퓇��3��l�=�
��G��=�5'�H�^X��X���Մ���Nx�����i�~sqϱ��F�h�h=���Ŷ3�-��[�ky؆=�~�z-�~j��?6�S���Z�W��@j%@�ȵN�n��D�n�]�l��=����cg*&S-p��E�CWKS�.��<�p7�2>{rӛ^����1N+���xZT��J��l���;E��]f�b619D�<��������0�x������oa���9j�(&8�-ʊ�LE��d��w�yݍ��DյN;�,��������ݦ���-��T/����w���l�K������"UZ����q�N�h'KK���1�JF�)|V��ʽ�u5��&+E(Z1�'���w�j�&R��>����3fʾ�#9�YYܧ��}C�p�k����fTCɚl�J"��
�#��J&�.P�붛~�[Kg8㚝ɫ�md�c�,��k�JmQ����S4���"_��}v_����C�p��+Q/�{��;ު=��Pּ�P�~�,���s�Dl�Y��f��tY����
5�u �S��g�"��yʪ����ya��P�OwE�\ m���/�ф��_/
	�V�	hoeZu�5g��:����dT[�vV*��q��NO(Sw}�a� x�����.L�߮��@�B饆�ػ]g�2����蛹��{W������*���{��Af��Y�L�b�ױr���	9/�(OL�:�
�^>���m8�Q�4�x�� �^�^-��u.����t�m=2��VJ\�+4Q�����qv�W���҃R�A.cY��2�Vb�0�n���%���ؽ�� {�α��z���u���5JuҸ�D��I<ty�S~����Y��K懃��p�e�L(�����g;���F��;}TG��-��ӎS|<�1�����Wo�}�pF��ؓC�fL!	��Ny~��<'$a�J�6�G��/i�*���v!���ؚ��E��"�UK�_'\��S�'��~��aD�<��W���"�(�'q�1��d]��W*/fT<9%��95��;D�ά���Xt��w�d��U��u�2E��ms/��e}G��O�>
�3�X=�6�!�U@��MA6�����q���[kG=��<<{�(�,�6�zQP0�Sf��!3e2on�4�Y�l�ZO�\�f�qs��Q�H�"�J{W/x_n=��m-�,)A���~�U�H��g{���S	�wl����Ѱ�U>.0�C"��-+mӎ�ys8�\2%��|��S�5/������,agR����Fs�>��X�/�%{g��/�i:C�*g��T��8r�C��F��{��X�͓�$X�n:�H?��V0�¥�=^�Le��R��w �Y�Rr�e�;�	�@�"w�"���H��t�M�R�P���"]+���W:�k7C�CkH�Lo-=��EM�#G}cpfs휳�����~� V���nٶj��3;�L��/����~[%X��,Biż�>�+mmL�0+�w-<��NQSf4���́ �v�ah�dQS�'<�p���,�{�����-*����ȉ7=�{� .��2r�`�6�����R����Z*ã����灌��u����V�u�����M#�p�g]�^ye+7��"�s��k�JӱRᮢ�>I����&z]Ž�eŻ��/b~�G[2��c*+�_�Ӎ���8J�/���.��q��"��B	�˭�ۜ����ݐ�P��5�S6x%8�N&^�LMGC�sUP�2Ep�d�K��ײ����s�M��k��T<���'J��f�My)p�Ћ�F&'Q8x�.7��Zf�ϲ]���ˊZs܀�Ѱ�k��L�:�3��&����F�6��U�\`�Dչ��k�j-�K��������海a~��ϗ��ʸ��C���O���ǟپ�(f����
��p�Lؖ�Hn�0�V��%��ˬVX>���ϩ\VF#�x��<z)�ҳL���C<����"�)�V}".܈���CGq�y��ך�0a�-�,�6u��l����a]�y{Tl��:;���O�����ʹYf��Kt�}�s,�U�|-�� _S]n�y�]�7v5�m�V�;ү�Ƚ�61g�� �3Z�6��h��'�g�S��4���
����y���yJr��'�ΰ���P�s��^��)~��l����ָ_��fz��;�L�7�j��u��s�utX��Wic>�����v�k��a>�R��W�.9zT�	N��Ζ�
g+v��>]r�6���t�~9���K/�%a��Ip�~`/�� ���v#�����]sVf�ֺUԄW�����a�_[y~�(O<tp���'J�"�t~l�
���O-�Hɜ�-5nS!�
m?e��$6��>4�Ԙ�CԄ$Ĵw�T�𺖡�uLG�"�k�[":�������Y(�gm(�a��Ȕ�����ޠE�`�SWxP�勮��e�tϹF˷����d�E���k��=^o��_��xo��n"h{�ɰ�"M!����񙌬���}�P�,c����.3�u���3"��r��~�����H����c�L�C���ט����&n�Plڊ�x���yV;5Cb�nb���N��1���DmSekdFr�ճ*Hr#��*߮�K.�������e�)T<ءXV�Ь�4KJ�9�[�����c�ӂK�����s�+qX�]t]���$,J�㒄[{�j��l�k�J�u�����oN�~��7n�^���6��d��߽�  ���}��<1T���[D��Qd�襉p�E�B坛����̸V�R�ޝO�����˛�߽�p�m��ے��4O�>�=e�-��
L�<'� �/�~h�!�6�;O-�{��qJ3ܲ;���j&Ă�&�Q9s��+�����<Kì�[��{�yG��ݠ�n�y7���ǽ�v�Mg)�J��G'KE��SR}D�u�,5o���ͫJ��5�Oi�7�5]����HAZ�+��=Ez�E�7��%��u�,�L��;20��^�G<�s�bd�^������`!C*�#byݍ���&��w g�ˉ���h���4/t�@�T5�y�����r�s=^�� -��yU����oOta�^
W�L�����kѷO�`�B��F����rJ>��ɋ�M�t��9���DiQ|�o6ҹT�p����ĽR�8��R̨�e!Җ)P���͏J������S&��-������yu�u�63�Ü�]�n��U�x�f�6�"Z"��:���Ŀq�C�f�wZ��4�SP�vO5�k������A=rl�A�v^7p�F�Q�Xs��ՋF�{C�Q�ɕVDC��3w�)�ȓ��1^�����\��;:l�Rz9�k�rͳ�F^��慤�����������\�E򢷣Vʼ� x{��9W�EPϥW^�.滈p�Ts�ק����e�����Dnec�T���y�n��~4y��%�[���R+N�qqO9]E�}N^;��m=4�B{�mnw�$#v�9W��073�ā�`�hB7�X�3]mJӾQ�f�%��0����x�q)��,u`�<�P6'R1+��e�q~@���ia��v�S��zQ"�r=�4����v���'D?+�����$W���%�Z<�7ᮭL<%�VA�w�^����7m��ZɎ~Sq�֌�1bW"x���8�h���Fj˪g���դr�{�-r�rE���
�}�p��m�fL!��s���8AL�!�Cm���{�}�����_E��9���*���#s]&��B��NЋ���@0g��<�˾�)j���v�t5�}�C�x�<���Ō���X+9����o���Z�r��ʍ����_y����C6ֲ���K#�ǯ#��'�KX=�'��Osb�;9,妐��۾�-K ��L-4���^���v�=*��F�wX
WbZ�_�Q��39v-��P�k�T�g��DP{2��`{�������s@	M�;]�8d$��le-�Mb���<�1��`��E/��KA4�%z�	���T�gU�'0��xxL��\�Z��PG�M+P:>���@���٣l��K���Hen�����P���O[������k�t�*e�l�iު�a*H��S];n\.�Opi�ݍ_�#�����P�����D%M༲z�95��J�oh(u*�
t2,c�ZV�t�=ɇ
�Q�&v�ȼ�b\��;*���N$��ı!W��L��"���
(B}.sȠD�6��P����{�AYtm^t�=pp�C��U\e$CJ2���鴢��.�l����i��_]b"����C�i��s�����j�K.L!^���"=��_�GY<T���C�^y�ap�	�ݐm<I]����6�Nab:4�L	�w@��D�6�3=B����X�20��v�������F@w	��G.{�����,w}�U�<:��@�q<MR=�gʗu���1�7���م9��'
9�>�7�2��g�Q\b�Ӎu�&=��_>�ʺ]��q4��5v(�M%1)Z,)/��v*ܝ5�뢢Ҝd,f��L���]�8��=����|�!����l�1����v7sR�%�Gf̤Mν��m�^E�p�[�΂d��~��f$.�l%p�� s��JN��uz�j`VX���g.v�ӸQp^��ڽ}XC�-Q���8�̻�t�[�λy\�:N�PՊ����v�hF�u%�2���C��^ٰC?,��i��^UFr&��&dz�h���X�	涱v"ڇ�q �!֣��w�GY20����k��V4U����_`�{T�ƀ�т-�5h�Š3�[|Ԡ���*�i?�?;�XEAuZk���VJò��F���1��>k#�~�vX[�r������a��f�'/n��H,ڛESNW^Tю}ڕ�n��r{�X��x�rRoR]����{h��o���A|e�+����0��e��k[1ry�Bs�;tR=��t��ͪ}��+��k3��D��4y�4��,�8�
�`��6�:� Խ`�(��B8��z)��\砱S����U�&��O�@��R����m�4{�5�T\Whۮ�r&�Z��WZ��5�1*;Ա4�;1pMp���ou:�B�g,͝��]brZ���	�+�ZҨ^j��V9���Ьܦ,�Q�|KP���]�k���w[tR�|@3b
_B���sz���k��ǧW��8;��1�����tK��	�u�Ae*poh7��,�)�ʦ�������ӋO�f��L}�9 }�dDnԍsn+�z�\�F��>��W���-��w$�,��y��7;���^�)%�b�����
���g"��(����!bWVv�q҃��7�w���~]��K��[�>������-�r���Gis��(ХvD�n���rY��6�/��kQx��^p;g' h�M�����ˏ;k���� Q��"�`[M5�[]ib}ݣF�� ��̀f�Zٴ�n�	F8���A<cU��'s|Բ�vid@�&�jU��`{�.+���/���2zp��7�����e� �Yܻ�f�\�+��jK�]>3�"�՝zU�T�w���Nrr7�7�٫F�FK�C~�xBG�D�t2�hD�l�7V=D�z%�8iAX���͡�\�GY�כ/"F���+�y��&j�/�/�g;�\�C�4u����K/y��u��4	�=�Ev��`�r^��$�H��,��Ҕ�60������/43d����W͋uW�:�ɹF�6ZR���i��} t����%*�t�sLt��{�x�� G]��b��,�-*���ռ�Rŉ����S��}ٹ|�l�a�M4�v�b�*_vY�ev��M�Ү��w/XQm��!�r�M�cp���ڃ��	��ﴣ�GM�6c0�0\{�V��`Ŝ�_X��'t ��GU�@eIܻ���g�t%r��<�}�C���-��|�h�ع^�$e�@�7���^��h�١��~{R�դAQ$H?A(�b��QDPĕQ��1TQKJ"
��cUDƑ�Us2b1c&-,��Z�	����R�ecKA`�4E2�*�A,Z��1R"��[ab()iJ�QH((ZPX���ER��b���F+֑iJZQG�S)U���9h#��q����eQʵPĢ�RbQB�Kj1�-TT�Q���X"!��TUX�6�F(�-n%F*�R�R����r�lƊ�b�Z�+Z+���2k�(�YEUYZE*"�mQm ��*�#%ZX���AX����Aeb1Vc���
("�b"奵�V1J���k���b�URѵP��X�r�b�!Z6�ũF�����m��im)[��h��(�Eh���QHU
�sr)Z"Ԣe�+h��_
>I���SpA%�v��sM�}u���j��fe�V��CoB�]��cw[�(�լ�Z:`b}8��˓�w�5�� �Y~�;�����-8�n�GW��±����O%.�7v�O��qڝ����N�S�]��m���k�ح�;z����n|�92X��gh���RN�$�p�vcE��<r�;�kUds��@���pm>D�������/���s�\
��x_ۉ�d9�}�]-k�Wa9�{�䩈;��WK`��;��=V&ƽ��Qa�h+%R/��U��w���҈��..��K%��:��w�f�{������N�X�F|��XɌSw.���y�b��\ru����W�2�e�C��VveaC�e��a��WG_��ơ����|NF���np�{��*0���"Et�"�g�@Lԧv�:Zp2�Ƭ�n=��	WTc)��ta��Z���g�f�%a�Ė�������twkd�^e��t����n�Q�t��o�J��_����+&���N��S2����WD�D'��6����Uɶs�l�ONf�U*pS�	�D���kM`�!�x�O�Oiv��V*U|+�b���C��tB�ޑ�^�j�&�m�|�Ji0���Fb�ˋa��ii���]ݷb�M�Pa�s/�Nm��;� �F���1�;�#�k]��^�ǋ��񽹉A�ύĔ�-\�oX��]q7�L�ip=\�$��Y$j���eO_���y�e�M!V�g�[F,�訵o�lf�"Z�����@�����ޡA��m΋�7��_���mb��T�����GU�z��u<���n碑��p�ᨊ�&.�C���N��E=+������B�$*���`�����N�:r�M^G�l��U���YQ�{ғYݬ�Gz�D��NBe@�5�6m�@\���!��r�&WcOr4�Y(ɞL��g����c��EM����*I��Lv�襟%�],s��qA*�9�k||8m�7��S�	L����f�zl�)��]DILa��]���I.-���6W
ϙvxA�ĕk��}�쀻��M�+���3"&��P�a���V)�T���(	r�7S��*6��!��yW�����F���r��y���,A��Љ��=��<���m��%�r�Ku��j�zT�p91�^�޹פ�4��C��ôP�e��T1��6�z7z��f�S(ҋ<�V+�ꔫ�-Ԓ��?W!x�K�	s��b^��Y�]NۭF���R�mK��us��i�jgVF��� �f�v/&q�����!�zx���a�F���s�Vt�/ޮ��%=��$D&��h��݋�C!���^j�xSx�Oc&0z�7����i��oY�ݰq˕��@Cx�������Ƃ�os4ݝ��s�)��h�B����z_�M�g7tv�|{N�#I�61�\��N`=>�V�xh���Vz�-�jD"t�]O#m뒻�l��ӂۮ��Kob�
a1�^ˮ�e�[���ܕ/+��}4�z�����i�݀���<�9kdf�/T�!���̨�e!җJ��WȞx��y��Իݚ��M��K�*�}f<������:�tg�����4������,۬����!IS�u�k�/�n|7�O�s�z�֘�j��=E��Q"��k#.���Ι��3�E�x���.�t�]u�^��H����Ǟr��].۪EB
V���]+Ց���,���C��x�Ixo��١��`N��u�+N������ܽ�}��^0�>}�+o�� �5V׍w��lN�bK�2�]�x�3.�Xl���m�t^Z�	�>��w������r�S��r��Z�x��C����^�i�f�qM�$7쏴P1vLhzUj��Ϲ> >�.�'����b�b��������V�	3|�D	H�GҀU�K��歪d�t[�70�ȫw��FK�]%o@pu�i]���c��*���򲛩�Q�m[�Z/9��*��Fe�2���\�}���4��H�+%J��Hz�Gf3P�������K��K;�3�峻�y���o��unp�WΝ��1�u�c6v߆j�'6�3�BA1+I�u����8D�!��v�tDq���ו��VKU�شKZO��z+i?m09մ{z�x�`��v&���+7�W�C�>��͈z�Y�5q��og���<�v�����6�'h�9F��̭�ĭ���p�}�{N(r�,�6|@�2S��n�P��F0�6am�CK���fx�4�(�]+����J����ӵ�@�;����ѯk��_��T
��}Tپ3Ei�>�yn�-bn�o.%��ùn�5�C��tr�vz��;>Pia}��� ��v�%�6����@��!3e�66��T�.;�:1�-+@�N;���ËD�ԍ^��"�C�.�Ɉ�<�}�4}�+��%Pw���x���7��`�u��W[�>�gٷ�֡Atct�O���;�Q7���MB�z���]Q�*�NS�iE2;����na[[U��wo
x��޴d�����۹F�T�^�΁ �u�UP�DaS�'<�p�zcV����Δ�h���h��r_V�K@��������yT�|ύVL�k:��vܣ�2��b�tv����e�~o��ԗ���|���+B�YG��!�6ڱ5�h����]`�O�]��n�������e���Wb��C�^�����P0N^Ş|��򭛒:�_�<e��H�c�ޠo�L3h.u�Qh�Љ��f���'���Vu�U���n29��r������8��4�����z�P���6�3=k}Ť��Ԛ�+�mK��w���'Gᒼ��|=d
�Dw�9�4U�m��zr��?Uf�͉Q^�'M�]	d$�|p��p�!�ӫ��_ �g±Oc�M��� ������j�3�����R��,RQ����6�Ό<����B����\��1^73�q���b���)�6G��L�:�m�&��(ʣ^�	��D���+ڵ,Qj��{�}�������a�<:����y�^���l�\��>�FߪN7aL뻧�:�O��Y�?3�m�Ya�b�b�k�'�՝��y���v���]���_�M�����1�ӍN�_=X:3�)�Xb�״�jn��ɮ�]�*Q"�PP$WU1E���Z'�Y��Beiƥ��~v3�	�3�ʍ�'�g���kz�뱋���Y^��`�����Νwd72��Â��.=v�m!�5����o�%�C���:(l��X�'/i��]-��v���ibR�U��y57�5����'srG��E�,���"�}}嫵�x"�a��{�Jޕ�zo��O�k>������Iꮡ�g�*f�;��Ζ��5Y��b珑o�Z~��j�Զ��r,ܤ�?
�g����>,�S�G���A�D���C|=����*v�*^��L�"�:���$�x�TfҦg��ىtHN5�Λƴ,%��Mo��g�$F{��O_���E��'���AC�i,���>�"�r<���/�ƶ�hr9n��l�d���P-l�]�}
�+��:��sˢ���#A�0I��x��f�f����UwS�`��Rz�K�	ˌL�G�ު��xo��NDC���5�k�2M3��z�� ���J���}��<�ƭ�u�����ӗg�yY�qb���2J��PV���o�R��{V$�}��J�P�Jȇ}Ƅ�S[V5wz�{�I��i-���򼎚�e3ԵIP���~
�S��&�ȍ�*���N�.�9�^8��^sDp�ۀ�j���KT���Z��Qa)�"�si<�;RK�!Y�s֚�޺��_<���D0��MM��C�:8g�P�os{T�xH��kw���"w}qo;kֈ�˷p�;�I�X<��s9��|@�e9��U�>F���g���y52�`���3�x��ޣc�}�I��&;��]Oc纥;�]k�{����>{t�螬���>R�n�W��r�kS���)�9�Q�T4I�'
��}D��U�}�X�A<K�>j�R�7ޕ���ZqM�//�eH**�y��,A��՘�vV�|� H�2R{JxV��>w��`Z:�~�={͌��N����i�n�%�g�}W_���t�N����˅��:YoZK��ifK�X�6sa�P�RR^K�^/j���B�UF���\"a@V��NJז��/۶L�J<��v=t{��|���C,�9�������x ��;������oc���I��8N���!2��s���[{�P+�m�J����-��;���Zz�զ��^[�;�jv)����-l�`�u�C��\̨�e�Qҡ�+|��S���:���q�F��(��.�}f�6_�}j3X��p���9�0�:��E8�aco�GC�xu��xgL��u��)P�Y�r��w#x�q<6}��:�09R�e��{ˉ�=�b=�P�h �-!0W[���SV����׽�zk�Q�V��Նa�Lz�d�y亷�@��������%d+��;"���$Uh��Q�׍�U809![�T :���m*������}�Z�b�t��u�gSMv�%^�O���k;����#��d���,»y� ��p�C@��5Y��=ݙ�G�=��������y(��fu-�c}~���J$��P��hK��	篜ǝ����^[�uϸb�ww�x��S�_�'����v\ؐ���ȊNH�]/-�~�PΓbccv��؞��H��J���*1��txE�8�)�Ju���&���i-r����p��XO�Ԝ]���]R���d�3D�.*���p���<sG]�|%b69���xD������ε�F[�S|<U�Ӌ��.��v$�m�f-��"�bV�+|����,xjEX�>Am�ܹ�s�`��_��'�x&�����#\N�,⠼��r��#�>�fp˾�{r�!>f�t���P><�n����<z=V_c�sՔ�.�l�o�y-��0N��ڷO�D%gc�\5R�<�zVG�a\FZ���kd��dv������:0���۷L���(�w�@ϱ�|���f��W.���W}��Y��o�&�\���o9�ڎ�t�NԨ}�N�7T�x�5Ӿ>�_EU�j��������������Q��C�ہ�Э2����Ƃ��ǀQIv�yg22�9���^M r'�{�m�5'֏�ƑIe��v�
��!�RMٗ�#n�&e��ðcq�l��0���uwu�n9���N` }�c�y[�1��X�#�T�.֎ނy��>���Ƽ����&��Ą~gJ�oh(t%S��<S��cRҩ��}�G������̄���ո��^hB0�䭞���Mz�k<<J�w��m�QB�qj]r8D�7GZi��.�铽�{�,�p�<Vς��7�P�^T�x]Q�Te_�NS��iEbd~���w���5��K+z9�p�=�Y/�^���n�I�+�Ts6$��"GQ
�y5�U�R���kw5uk�P1�ol�~���n-<e�i7�ޠo��I�Q�D\�_&��H��דV��B��=e?K��ny��n�b�<�f��#�h FƚWJjd�T}�v��*�-�D�\�\['N�:��)��F]���<�:?�w �^�
�z[�+{J�m����rϜ���]�^y9�ZbJ�Bg+�k�VX�8�WV�q��v���~�h��XY�
�Z>�
*:�����.o5Вx%.n��^X��Τ�U������qc�c<'+jϯ�@T
���\=8;1c>:��)��v�����#w�3W�cq��P$.r����t��n�y���] ��RA!MY�X:�N��t�V�:���h<���<�Hڲ��R��?�y���m�ҊݖrwS����yF#�8�Q��&p2�S�ݚ8.�n�|.������l��$���͉�왽|R�g,�(~�����@9���Z�#� L8y},��Z�<7�Ou�`JS�~���/����Q�0���ī�%8����9�w���bo^��B/N�\�tPy�v��P#����}���t	���,�1���3��П�۳��qiym61����=X:0s�6+r���&�g+2^%b�ni�t4�A@��B22�e�B=*�F�eiƥ��)�F�ld�Jd��該��x{!�1��ܙ�,�M0D�BynT�N���󥦶!�G��[�%޷3gc�ھ�m�Yy��Y��V�����=^ ?����C�xo�q�CVғ�Ծ��s5������u��i�����O�ՙ�Eh�����^�E���I��2_Ik����~[&��+���H�D���Zh+�tC��xE�]�3Х�f8����7ڽ;�c˖ه��I�ȓ6ٳ/��D.�E���@�0�u�:f�Z�;I�$HN��������S���lz��u���x�.�J���~��l�ai�U�j���c��q��Wl��j��ʰ�D�A����+v��m]���K���;�.ވl!��R��׌�l/�r�y��r�x^C�`��k�mv��V��{A*�Xg�7yS��M5Vg,��p�q�Q�+gv9A�Lq0�<0՘4SC��,�w�-t�t��X�����p����
��v4��hn*�5�݌Zr[��s�Ο�^:yi�8���έ�;|�����}7z�<AN�ى���{w��������"_��l�I6��3e�7{-I6��w��t�c�բ�C=N��e�;��޸n���c��yx�8N�ۣ��*�)!'Ws�b���PV�iu�i�S&5�f藝.Y�=�ʧ�JR���,`��)%Ñ#���#[��
�����Z5Re"��y��F��a�ޙ(��Y��'=�iA�m
�-��V�Y����@+R# ȡZ��]��or�

V�l8����Q�:'|�^	F��z�����Y1%�K6�L��9���,���u78�1�}M�n��8����л��G�q��IHV"�!�{
N�;�2f��H�8S�+KxV>YY������T�f�.8�N�dsj)�R��2�ݼ�)��j���R����&�Yhr�7t83�h�%ɢ�*8��F�"�7�Pk�LPo�#���G1PZFZ׹ܝ	�C�b�W]�-Őҙ�df�u-��YMY�{�C�˾\d�dOEL�9I}�0_*-[�,�v�����I 1�@il�E��:jE���gM��3�hw;}�6i�ǘ��ՙ���[]�E'q���W�Fz^�2g�Ed��xT5f��S�n�ik�R��SB�fq��;�}���c}_7�\RW� l���W��jFr]�J:�CK^��JF��ё��`�n�8<r��\?
:r��f����UO%yڟm^w:]�f��k{������r���m��Hq4�����;�aUq"����j�/2�];+�T5���F�ݏ��vG,�������1J`�+���b���Pqٗf��������]�2�j���*e�W����i���SN8u����p3շ�6���j ���u�r�R,I�р�ѩ�L��]F��UET�*9���=�h�ۿ��=���_X�*�{�V�t�k`X�垥�e�X��9�U�`�hk��>][�M2��S�-<�s�yF 9d�9pћL͐v����ݎ;ʸɆ��9rV	�V@K+��0�"U�G���)��"*W�� v,�Gz��M�pK�aǌk�H�eՕ�G:�os��~�[��m���!3%pR��ψ�+l qՉ�Ӊ�����UMʜ�;���pnfS>�W-�,���P���(�t���WU�vDv��SRj�"��8r���Ī�kp;c(B$�*��;FZ�u�V�����狩�p+�k��Of�t|��E 4���R�m�-�r�b�آ%F���W"�s)��e���j�Ve�b�\���PQc�s嫍mkh��mW,�Qˊ�8¥�b��Ѷ��h�,�`�1l�mj"�*"����*�4-���
�U��R�UTiF�Tj�j��[U1���
�\�j*��-�m�(�YUmKUJ9�A(����Q�řJ1�`��ˊ�e[��iTUW+l�Z�c�`*���ܴE*PD�EJ[iUb��Z�啋iQU-�
�eQUZ�-+eJ�ܴ�n8eEPQb�ڍj-Di����Lk�-�DT�ƭiD�Qh1�W%��Z4�Z���+��V�ֱ��((���m����+D�Z�E���,QE�,���(�([KQT�RĬYe����E��ejı�F��am�����TU�#Qj�X�-����m���߼�}�tb�۝���}��A}Z�C���U�X�,��Ky
4��;3q���Ԭv�\�|C4���
��{=C������)D�E�1���Ux���!U�n��8ե����̋�a�vz�}��T�����|���H�c�|&�$��4��:L�v��ı�kj�wz�^x�u��7�J̓/����%<�GJ�lĜ*���N/�r���91�K=wªhᖹeY��Rx����'�9�^7��%����WpN�F�N���yv#�$���Xj\�f�R��2OQ~-�hͼ�~�𴎏5�/:Y(��'
��}D��~����;+�m�8��{|�vߢ��Ğ��,?��0+89ОÙ�n�w��7�9�w�
W钐�f����o]Ȝ�-g3��Aa�)��٢z3�dm�PQc�C*E�����&�ǔ����30"�W3�f��f��B�\w����LO).K�^�����*�8��Vf�X ��^�fL�o�z�-.;e����������-�\�U9��z�1y;"�Õ7(V���3{m[ħVBt��!2��룰
[{�E(mgҗ��P�VE�X��{0Y�TF�ˤ:[�{!7����{Ugofn�Q�wKzz���P������^�w�#=Ɣ��gg�ɳE�-oQs�����T�V�qz��ݓk�}H��VH���d�]��m�k�����O����S��Ƴ;��UѢ;����2Ҟqb��ƜK�����?k$!�K�87e]�":��'����ޏ4������:��P�����)p� }f�6YO�F>�z�<ִ:Uy0G��tј*deֻ<��L�	,��ڱr�?
��ȡ�c��qA�+��;��l'����!6��l��׫H�:>=��+&��QB͠�2�t�]Oɥ"x���=���Y��i��������%.�v»ͷ��X}u �J$��

l���?��3]��on(��m����̢��Vj�]DTw��vm�

��܈���DЗ=
���P�
�o_*wX�cz��5��EQ*,+\�e8X�q��G�[�p)�N�8�D�����Ou)�.������h�9i�/L;�Sp���p���\x�UQrV#c�����˶���E�v�np��>���w���g`]�hf�fb٨B(&%i=�Ny�+f�L��;�w�k��X�f\Y�:�x�u����^�
t��j^బd�@M�R��Nw��Yě�+@K����V�&�n{�v7�4/����J�,��G&���:���W��
rأ!�
�m��w���f��4�3��E�/Kԝ?Rg�;V�;�U:pQII�
�c�g�RK[tw3�K�S��*������V`C07a�7�V�;w.^���_�P��F�됇(xlşS���߇�3��傌�U�s�c�W��] ����lc�g���3�ZY���*�T��+���{4�q��h%���B��`���]d;��m⦠�i�iC��x�g8�X׵�j/�^@�UA�k�U��q'�����l�ۥ�U�j��,cT�Nۗ�S��5zs%(iE�9�պ,]�R�Se�v�e�D�,N�b/�ҡ�
R����\?c�ZV�t�d!q9.ذ�������� �����]�TPPfJˊ)7��fs�>�W[��*}�f}A��y�[�}Ts�|����W��:M+��g�]Q���52���(����NP���6�Nb�U*v��9��X����4:�{w(�Razs$B��UB�&GY]�\ѵs6�2�I!EfO@�O�9`���S���t����P,Ę:�3<(T=�ۃ��΢�I��ܙ�U�mB0�Z���[ÞG#c;�������P�4��qu]�瘆;E�Q�un�B:�7DoA�/�qPo7j�w,؇l�j���Q����uo<��t�f��!��.�d��� ������M�8��S�1��r��J�������י�'~�>�
fQ��b�Q�ӄ�K�؁{CF��sf�-�r�*�%�v5Iτ��ur�qW�t�ν��;+��6/ǃ�%WG��;�p�Q�ۥO:��qO*��ǉ���6�z���sY�C�{�j��͗%g!8�v��VX�h���j�Vy�8��{���s��,,�<+a#�y�g��e�`d�sy����J\����WdWdēh��<u6��I|�8��#G�G��[V}j�C��r���������q��W4)�Xf�=�$� ��"��GI�s�Ӯ�1�����4T���(:f;���ܹ(�+Q%�Z4�;�f������ �S�[7�4ﯝ-�dXX���a�s����w��^Ԯ�~�b��R��Ĺ�ͫ<,��Vy���MQ�w#0�5;���M��_%��vЮ��b��Lf���5X��U�Fr�`g���KXw��=�}~��X��<:(�_[L߷I�=�N �����٥1y�XϢ^K��T�#�E��3R�ۍ�S�L���1�u�	�Vj,CEF�t��Ҳ�,.�F��X|e$�z?0���Gp$�~�9�iR���zK�k�rx���@�n��BQ|��F��_kr�a���+Z��V$y
�љ=�]\�.�Fbt��T;�ꛐ+�oi���a 7�̅�.U�Ab�,F�������LC���8f�"���f�Q�2>U	��Y{v%bGj4mZG.4�)��KN�*7�l�9r
/��=�禡\��W�uP�u�;��6HPݛ�T;hӤ���+-l�T��*��>R-�OoWLT!�B.I�a'����CQ�ӭ�ܧI�����EE�R��r�]����3|͙|�� �w<�/ß�@�ؖ�A�h�<#s����ا@�{�J�d����0��Ĝ�Ǩ7��/��<6�Kݑ���M�`M�eN��|�����x��ԉ?qן!Br�3BX���*q�K����fEᜥ��X;�*m��5>�e�5ګ}g� /*{�µB�b���E�����+Tp�u׽��G7p��iY�N;&���7ka#phN���ĸ�9RMrc�ؗ<)?���Ŏ�w�Q�}{(b1��wO�^$�D�;S�&��p���"�s4E'1���]���%ŠV�7(t�mFS,i�t؍���H�
�' �T�y��x{��K����D�^�"b��K,����Go�ߊ�{+]�UtdU�f��(��r��bV&��tV��D
 bq#%7vW)+�΂D�-���(ǲ:O��BH��P�~�SҢ�e��4��*��R;q���Sm��&00T�!U�ź׌��/���ג+%i����)��OS��w���5enR��-/�<ݭ�n>9s�W�6��#{a;V����W^�᜙N��̃�.��՗���?T�O4��f�{T_��2�[;�X��NQ;�]o�dx�>/�9���4��R�C�yh!߯#V�x�K��yx9��7��T̩��EQq֤T�o���,��K��_��m��.էyJ�Ec!�.X�����q� ���}ku��D1u9
�����N��d&f��;S/ ��/9K�W[*��uQ)�ŗ7O�őgJD��Kd����S�)kdg��z� d8ݰ���B�����ҫ4椽��1z�"��Us���9i7����ds�pg{&ڮ��gE�sq
�����x-�S(�}Q|x.��P���qX��¥�hR��>�(<�u��<���rn�U��3ܐ��n!�;a`w��3�af�Aai	���/|�H�������Dv+wF�޶���͏l碮XWc�߂ziE��ԈL�N����etHT�Ud��\��t��ܐ��X��\�m���iv]Q�ܻ.lHZ�܀�Ȏ%����7��c��s5��t�:��g�}랬GO(B-�Ŗ(R�{���	�9e�撕j�8��w���̡���r�@�uH��=��E�S����\�'*�[sΧ�`Q�"�H�^���G�T���F�{)�u��Z�����M�Wu{�H��Po[�Y����//֜�H%pډi�c���5N7p����p�!�9T���i{�����2ta=Ƴ��6��;S�ׇ%�C��Pxl�'��]�C��ͱ^�+Ό���b����q#�
�H�����9��5X�Y�٘�3P�PLJ�h��"u���;��Vӕ�/�-�eIf��V�ś�\O2�ˢ|W�a����nuhR�O,��-pwy�k{6%1�͜8�N�`y�؅z���!P�ً\�p�gh���u����Q�Դ^�$��jv���� ��V�~~P��f��@{ �a��çj�2���e��2o��t���L�}��=�do�K�HƝv��s�l3�v/^�Q���RSyeR�k,s8��S���hׯ����)���C�N�7T�x�5Ӷ���T�
i>yC�;���z�I1�C.G��:鈼�P���|\Br.>��i�u��\ɻ��o*�4q؝�hhı�DUh���U���*��}���{W�����<w	��]F��q�<+uǐ��Me̼�0_Y���y�(��a���"����睫�k�
�P��cn��#-mzq�^�u�w�bU6���H�������zhu\��n�WK��x�]�z�N���S�)���x*;O���F�YV��ds�v==y�g���?g�_�4A��mU3���v*�*Ȝ�n�$s#�95]5r�:^�wQ~��#`kРX}��=��x�0��|�0���vc���Wm����[�l���vy��!àr�W�uܧp�e)Α��Ϛ�0o�)�sx��d�}'��e��ٮ�r]c��\���Vð���ǎ��<�f�<:]��t:7�܈{��o�D\'�ݗbD����%�z�N��u���U���p�ï`�\w�ߩY����1����Փ��x���L��ڝ�֌�P��a��^ٝ�¹W��WjNn�u�Y�q����i�u��X1��H8_,,�8V���j3�]̕��X|��"R�`�;��O�˜�����]WB]_p1hbu���z�	Yu��D�0�,�����B�)Պ*,u�lU�kE�;ru$ֶ(�t�nm'<9�i���9}f���*�g�9Y�~��#[�b�^�~��e�{vi��2󨃣8�����sOz�M�{s����]�YW����-l٣A���������"�&�nft.crN��f��:���!�ko;�]bQ�c�.�Ʊ�g,N�W\x�������-�)�����f&�U;�|d�@%6��n�:<@ZXrR�k�px�Y�śc��P�D���YF`�϶�vs8)�R꣪�	�/��V�x���T��t�;��E�MY�P�8���z܉��S/�����9:~�/��ΰ���R��}C�e��]t+��gc&V�p^� ����Xg{��Y~�a�uޭ�V؜�܉��ܪ�]�*��V=� 6\\�!��0��z��.�g��Io�ǺW㓱C)�ӂ.5S�®�]&�\�C�)%������������k�9ozk�һ�y\\��|뚳�f�ذ�v�S�Y������+g�,U�`�j��*�ob�W�Z&+���ɅK`�C�!>����5���D8�dʳ�^t|�XpZ�N,N䳭-�2F�����a��R}|���^MJ����?���7�n\-��睙\w��n5��+�G|p���S/��C�)�a��8վs[��]E����}R�2�"k�^5=2f�W�}���o���a�D��ן!Br��hK�����٫�N���}z�B�<�LG;彖�v��հ����;��<l�o��]%µ�e�O\�-8���-���i	��;�$�Ki�_�O�s�w�qx5��������:^���d��+[�q�KJٽ��(��F�=��~�Y<hl�A��J.)�P��t]P��{��P��EwRS�{��͛M�j�WǬ�[!�7;��q���q�cG���p��j�����ddhnb���N��n�?	^V�.�ȍ���M.��e-�O9���[��g 듯�\\U�T�XNb���0ד˰�d�.9�����u�莫�I�ʫ2����.�p�<< �_���/�ހ��@��RQC��e�Ne�q��KS��T����J*/v��Ez�E�cQw��8�~�C���B �=��o+�Կ��H������9)�{��4�cu�U�g�}q���>���;���3˼��Kips-�������>�e���i�%�	�>S�	guuk��>}�Y&m'���.y]���B&��N7NT�z6ϰ�g�j)�V2K�9���+[�+������C�q��0�yt�NU���sV}�NSU�V��������D|N�p�:�	�)�k�'4����S�9rS:��9����Fb^��C���(��+�+E*p���g!���EW�>o�4:�������ï<����}j1�K�5��n�f��r�y��r\D���aeXKV��P�N����_\���ڬ2 �I��T��9]���+i��Ƿ넝�0�E�*B������M
Ԧ�.Lt�B	 �k������OgI�<�����qz��,�����s�R��d�tp)�w�z�A,�C�[bJ����NYj��4gt4��gkd@{K䎝�MV0t#)�����!��z�
W�Y��4�<ͦ��8{n��r�=j�
���T�F��7]L7bp�|��%X�ޠ7ib2C���1U;��;�e�{b�{(����v�GF�\Hw	�X�~R�G*�8-���
�՝E%���h�s����뢀�g�.���h���s��B�E1W`���H� Y:�}N��e���ib���§bk��,ȒӇ�=�B�b`�p��{�KFV�,�kGN�=f��oM:�b@�m��J�F+v�Tc+��!��!�\2�����e��F�m�9�����������9Eo;�jh��	ʑ��j}�FLOl�kf�O���ٌd����\6Ԃ�7׃������l�cu_K|��y�_��iP�K��N�ݺ>��Ĭ8Cb�
��ˬ~��flГ�w�U�fMk�8��i�]P�HE-��)Y��y#39e��L�54Nk��d,,�����c#�mռu:.$PKwS۰����)皭��i�K.�!�6�]e3���z=��W+��5�wŢ�ݹ|�j[w����qed\��=F-�_m5�><��r҆fm(j����o0�i�tlG]�4X�h�p�W�WΰM�$c�\E�{�[u7jv	υ1]t��D��]�X+�u����xX8o9jz��xN�������B�.��*;� �Eb;�< ���IxG�k��(j�3bR��Y��5�7aqF����C��@CIڬ�kK�����j�]�V��.�Uq�h�൸1%��ZZq饳�@�y�;�oč�˱���|Q{�ܔ�r�ޗS�n@���h�������]\v��9�.�=�H�{�p��w�x�1�̽ K勪�3��M˅�ϩm�@R�#Kv�k{1�x��05<��I+�W)\�^�-�5F���7�+1Eelu�;,��8��{�$��XAd��\����k�����h0t�2mH��F7�s[R�tn�������:tj����M=ցho#-������]Ȭh�rެ�w9+�0��¹��u�Y���%ݼF+5��Y�]n���[�alv�[������mBL��j�m.޽��QƋ}��]ˏ�LhZ�-���7�6��k�{Za��T{��dѫ�b��%�Э�o�@�>4��s]f�rr�����e�!�]��,+�S�{f�J�^��7x��0��膷޴�KY}�j2�P]�����=��l�~m�R6�m��X��P(т*�����\+Z�6ԢPRҪ�T�"1jTPDVڔ�J�U�"�[m��jʣQkF�-�����UR�k(��c�эj԰TPQ��J��!V�Z�6ح�����PQ)mF�KiZ5�,��J4b�Jԣ+mmV��[P�����J��Z�QDH���-(���Q�ԶU�-�)m��PmJԴmaZ�֥��`�j�mYZ�1kն�q�)XĪ�Q�YJ��Ŷ�h��F���#R-�U�̥���EQm*"5+h%�X�eh��ZPYEB�LJ��Z4B�4��ʪ����-�P�*R�mb�PQ��Z��m���V���QDF�JŬ�kJ�[(ZU�%E��ؖ����������j�&KaKe�ƔJ%�B��6�[edJ2�KD����kKj�j����Z�.�ɯBM��5k��Y
y�Y�ev݅�/#���F�[%�}4\�>.l����2�;X�rt��x���W��L�|:\��;����}��0::�tN����uC�ҫ��R��y��q^y�����2y�ֻ�W����%
��D���tY�j���Dl6��	�� hL��ѹy�ե���y�ONZ�S����7�H��55�cz�z�lN��U���AB([4%�te��c���v�(�CL|�K�����.���;�f�`��'�")90��sЪjte
�[hL�n���z�~�EK'"�k+zJ�p�5N69:#��\hHxʒB�2�+�a�8LZZz�]��>�c�*���V�	Vha_K懧ܠ��q;ԻH��31�:�����1�.��b�n��r���r����c�K�t�����ň���=ʻ�*��Bݥ��'K�F��0קچ�t��Hp�Rz_�����i<�[Y��t��W]���;m��(;U��F�F��q�y�1~��d;HC��|6�]8�:�߇��.�ʵp�lVf���pE��vHP����߃x+w���O��hU2�b�'*ݻ��t���{f�=c��{5L*��<�Ҏ�}�k���ۥ���g`�u�`�̀�Z6�X�!��U�}F�m�׷��u�t3�o�b.7Sn1�Nߍ1,��&��O_�x����,	�ݣ�]F�p6�7�7��8Z�.N�.��P�r��Y�YX��Yڪ��1SPE�N�����>�nՑ��_x�0�ޫ�N�w��,�f�Y�3F��L�t���7�PZE�T�N�n\.����]�
Ï�NܜPt��3P�`z*�WU���"��*��:�O��)���Ѳ���;m�_�{�S������������,g�Z)��U���*��Wd#���&����r��R�Ӻ.K�W?q�����l��/Y~�:C�|7�$�y$Cʨ�g����p`����L��7���{	E�]u	�F���P,�hu���ČT/��M���2��k��<���B_��6�-G����;�~w]�wp��I���܈�(�l��0�ˆ�c�ڮ���;&1��йD�="�*XyL�5�<�GC�U�n稇`��n��+n���n�Z�� �l+%�>��R��Qx�5/7���<��X��~��b�s�`�I��E��ĳ���(���d
[�t���7]�4�o�śզ�Vr�I���J�œ��K��s;D�{���ŵ4[�E��t����eL]�c�9��-�]�AV����;-Q� �Ѱ�[9�f�\��Gy�]��2��'D�0kl[�y�*�p�V��z�3��(���to�ecq�#�VV�ݒ��]�MwW,�Wڰ��/�MGC��:��q�tѽ��@���̾�f��c�aA�;�&t�ʿ7��It��V$��>�ŵ+�����τ�mY��)��p�m��q�cu��Q%���aN�q{Τ����M�B)��t��1����eV�/z�4���9�/�N���%}wYOɗ��/��k��WS�[9��s�bo���[l<��Zt���VX>��:�ϩ\VFR��;��o��n�.�f���aO��Mur��ڪS���у�)�V-�%/:�p���}C���mǣ����u�^f�y�V+O�w2���Q8�N�ܧY�<�WE��5q��K�%[&�WPp�����&{ S�q���<��BR��CEƬ��q�J�ȵ�h�V�$�WQ.'��["T����a��ܱ�'.�:�.<��:�.�C�gǹi�����Oj�Aen[[����,����q3�LS��Jd�␰�d ��
��>R/Ϣ{zp5����ׁ�>�WT�M�*�����8m�ȳ
m<��kK�j�sS=�N���J�wcG�h#\��/�)�u�ﭭ�B�X�8��{A=/{n7XO�w�ǡ�k\Ի��2Xٙ���C5�Sf:�Jݥv,�ӏ1t���o�p� /i�r��m:�J��'�:3�]m��I~S�WJR�EuL^]P�d�c�̽�U�ӓ���WhG/:�C�6�:��s8�3Ff)��ȁP�p��%iw"Gs�Y�t�����w�����э�/Sn?=Gm{�Բ�y��h~�`���R$��B��~f��;�^r��ktkY7bĘ�n)\[��l�F�V{�����qqn�S��&'��&�T����PIh�}S��F�zf�cgh�zFB�*m�N&FC�st_����u��Xs�$�91�lK��(O'X)�S���R���q�r���檒G2�p�!����8yvv���p�.zc[Su�d>����-�L�<%<�����^o@<=�ޥ	/�>�
�1�=ο�Ywl��܂��۝!琞�B\���*�dU�F��-q|��u��2t�(U���,r_��V�{۸&��sEҚ���Na��,�~%Fc�5l��AE��(^]g��9R�W����p;��]�L�[\p�a�h"�1��i�������c~����M�b�>�p0-�P����7R�efn�˷$��$X�9���������rc����:´���y�{m��9c�T��K��w���-���_vsE��m0,���6�"�C�Ә[ُ��c�{@e����y���G�j^��L@K��,^7ӻ��Y���V;`hwT1��������q���h���U������Q�ER\w�V���=]�Y��յ�ҧ�XY�N����Ӗ�tvxR�ظ�QN��
�~{vN�����������\\"k��cl���
>��-d��K�^�w�}{&o�P�ە��6{}9Z�q#"�).������Q:1K����:yCał�Z�/Dnԫiü��zU��וFp겏	�`�L�$G#^�T8��w�{��Ç\n/˻����^ݺ̞�u��B5!L�y�,�G�d��Qag Ae���������5��&�9��.� �ț\^�6;��].۪E�҇�2!2x�\o#wBsN=�/��;�ngpW|�yV�Cޝ�cas���"���f�`��'�"('&7[�&c9U�N�u��[僚��o����i6���z/��S��N���\
sb�Uq���U'�'g]je�C�J'I�#в�u�j�:�{%���p�h��=En��K'/�T���v�sY
m_�����sE]��5��r����/�"��wMb)y�>k��ǽ�p�7_Rɔ��oGk ��ۊh��r�gw����ƅ�7}j�u��K��"�)�ݬ����c]�R՗7{8��.���}��ͱX%b�t�im�;N4�xw�1�Kł���#x�� ɗxu0�&�y�(X<5��JJ'5t,xJ�5�����#�o�<-��~7�h��d�Y7'�<3��E�%��C�"ٸQ���q�`;"��8!��Kr�*et�\ͽ�Z���Q�N�b,j��Cy���%c�g��3��_g�b��zˆ�Y�0Sf`�(�~�<����Ӄ�h���D���D���jfo�SPE�cN��;������J`VQcӊ���=S�	�-Y�]��2*�4/���)��ۥ�;�֤LBgK���e��Y��h�𸫣+3�9�ش�=��c��^�v���q�!N�b,gJ�vB�T�*.��'ѵ��͵2�x�SD2:x�{��y}�G��5��mw�*�a��'^q�t��ٖ���Fݷ��6rr����#��}�a��Qr�Ӌ��<b�ͤ�z|���o���Y�=�K��0�,-������3���@O���{w)x),�_+��ݢ6u���i5[wE#Sk2���h*Tw۱��/�J6u��G�Q�&L[R;Y���GyI٘p���Wݏnd��tL����(:N[�91�V��O��2dk�����Q�R]�[,��`	|�a��o_"�����B��Q!'��������4�c��vE��J�᧝bi�n����O��T��D�v����%O3z��8�b	�i�;�S#	���;�xײpW-W���Uyo/2���΅g�l8��v"��iX�5?P�]���}'M�^�«#�#.�CL�ڛ����S#��g��Y��Mw �B)����s+�'y�|
{�f��T����ؤ���m�f�q�f������a�q�����)�F*�RTk���]���~'�Н1�������jN�NĒ�p��ЋNa��#b�f3�9[V}z��+��}�������D��7�+,�en�\V-ә�GՕ�%�+�jX"8��h�^(�ǯ�^U�X�cݨ�%�+����ϭ\��¨��=���ha�_x����4	޹�g���*��F)ה4�^fMW'��;D�j�,m	�(򱠅��Z>�x�����+:|2t�'q2%���1W?K.����H���u�Ճ�>V&�ɋSv��K��SԺ��*�}N������E�!�,�е��f�7X8((`�ͷ3���&�2�HZ|�k��q�
ܺ2N�gwVb�l�W%&�$�l�5۰k^�Y6��*_�yl��[!i��4g �m(S�G�Y95�l;�hāw�!}�be�_^�Â/vR�6��f$z�2��5N˘.ϻ���ˤ��D�0�=J��]@F�eb%gf������r:X�Y)�8�y�ӀCEƬ�Ƕ�e�.%�X|e$�x�{ݑz�}u�]�H�L���jd��ɞ�xd�ˏ49��5s*j姽}ar��Oh*�iޛ�3K��ǧ)�OR+G�$;)/q!��i0�c�nC�"��ޜi��_�w��w��,�v�x�4�L����L���Z�º�/.�G�K&X��{g��'j^�#�<xnS�i�[�%�w*a߇u܈��0��$w8���j��G��3����%�Ax ;t+�/��^ߑ��{���/���V ��VM��"M!�hP��y���u[C:�Y�ݣ���wa�w7���ea���ȼ6ܻ=n��G:�N,3���rx���_�C���ۯgho������q!?t��CHQ��M�	���a��:-:���
q`9ʒk���7��C�OQ��=;��yzoŔ)y+tX��&vn,f��j9�
�f��'1DP	͡��Mz��xK���Y�]z�Y��|��|M���Q]n�1��Fc���0B�JS�Ǽ.�oyj�s9Ű⬿O�[6�%-϶��μKq�^&{$=5�#���/����@!7`�V�bl�����Zg�����@�Rշܦ�M� R=[�Wy������`=[G,�Z�^]7�L+<,A�e� s6x�DL�%�~9y���34\3$��m�U���P� ���ܺq�B�E��r^�g`�Kc��J�6y��y?����6v��Y��9�i�B��粓�4�7\%�g�������~)��ӝE�A�n��;x�o6�����E�ca��Ըa3���(�r�[�y	���5k�ZG˰��wcs�\"k��8�:�����b���E:��C~��ah��{���|�һ��&���}�V�$��t�NU��뚜�a��c]-���(smS)�W�8Xb�>�gҗ=�]A=]�E���X������B��Fk�Mk�����yT�"S�̝"�Q#"���Y�7��fǥD�d�=����ƞ&�Y��(�o9��k[���:�S=����(��0l$Ȗ�+�a����%C�v7�GP.�r���_��&RGO^�F%WEY�w���m�4J텀뼌F�*o�fXN��vׇ+6S��y=�q�زC��� �	|g"�6����;�I�u�"�ޑ�J�Z�]�� �衉���#�c��<Y�wSK2b��[����, t�E�16v;���:�Y�,L�q�鳀�t��
^���2�\-�K��ٌ8"{�iY`��^��\ ��[��/�fw�������/�7���:�
L:n���}�0>�Hu�;����9=9�+��%��j)<���GV��wAn��X�1d�7	̸��ʺ԰�;k�2��]|w \z�n��3¶h�͙���X�dp~�ʒi����tz�S~��P�s9���(<6W�׫���`c�*e�ߦy>�F�Yŋ���p���O(�-��>{���^����ۿư=5��m����^u�Ǻ�*�TxEgA� ���'5w���S&�v:c�h	#o&Ǩ�:�w��M�Wf���ע�Z,�S�Cy/N�>���`u��C����!��\I��!���s���9�G�'h��v�7֝q6s��8�FƳ7-�{�����s�KS+�&K+!��U������b|e��#�����Yx��"�7]�s�w��1X�8�d̮�Jt�cӣQ~�}3�T3ꦍ٨����z���p7Ai4���k�sY{hߌ�o�O9�z
Ku�8fo(چ��}{�b0�:�Re����Wɕ49'^�39���pYe�wB��X~<��;5�v�{Ȁt>/�.���9�`�,^*lI���M���g�$���~�?f�%�w�=�h��%9[��K7R�g3�!���h:��}�Hp�<HU�s�k�U^n�M�z9�Ȫs��b^'W��k�+�pBvW=C6^Zm��E�r�԰�`���QK��8��.bs��	+��*�§(%r�g9�)������N�(5ƙ�H��+���q�5��<��_�������ʈp�y�2h�C���2cZ廳���7*$ZS��8��Ѵ��8ҳ��p�*1���o�-�^��/]Y��u5��C�kS���&2L��l���8#���*�\i�L6�� �ztf��A��=�w?�fb���r4݇5�3+9̋>��2�N�e"�꾵׫{i�0�|�:�VC�&�0f�O��QM-���o�z*�Z��I��X�D����l�����깻�յ��?�GCS�"Ub4v��]F/�(3��<�P�hKw1�#�; 56���ڍk��1S�z�/=u��ukH��A���*JF�T/�@�<���<��j���C���y��m��p�����f� 'w-%O��t"�c����s3[|6�nԣ�@{�Exm�E����*���oH�eĞ!(�Õ�,t������73��۔ī���㻰�����ۤzJ�4�ޫ�l�睽�-`���;77���W�ed>�u��M$�eU��b��j�*9�{�Ωc��z-n�l�3�������[��	pT���6�F�,c�3H��]�cXh��<
�����{z�<��D+������^�H��k��E���L�b��R�����Kb�٣[��L�cnAEA����b����kGǳn��Ȕ���3��
��{��ZV����
�H���on��۳Ė��h4�fmadz�e����y&�Kv�|���K��R쫦�R���C��GǸ����,ݩ��N�0�gJ�PҡY�f�9$
�;��%;l�t�\	�;�2�[�0�Ou�r;��eR�d�4�q��vZJNXK�U0K�Q�1���sC�Ģ���a<+�5}6i����n��*ȭ(��og�K䳺�uz��V8�jJ�{^u4�����H�:���{NĲw;�ě�tkZ�;�з�pI�V3^�|�I|]_Ś���#d�'��T��z=vY%9�Yn$�7,�=�BE�{�����m�S�b�Ũ�S�����rˡ��Sh�4�|���\X�wn�*���\�4h��x��s�G�GTڹeP�Jo�R��g1/�C*B>�:���]��e�M�*������M�jY�]-V�NO���$�j�V�:�=6L�����k#�����>������$�A�Ѵ��K�Z�-kTPj�ZYcZ��
5iYPQ-�X��j�A�Ue[-زQXT(�Ս�hV�]��U�QDE[k���V%��)QbԱQjTZR�J%KR�1
���Um-k�ܵ\Q��ڪ��V��ڌ�*R����V[m���P�KX� �[IJ6�-J[Z�DKJ�m��d�Z,��+ckl��*5Z-��EXcr��J%�aQJ5����KhZ[,ke����Z��[�E��b��
�4���դ��5�X�B��kJ�
U��Uq̫���Q�Q-j��as*�յlZb`8����V5H��F�Zص��V�jZQZ���ңj5A�Ak(���2�R���E�h6V��̴m
Ֆ���ʨ�Z�[�.f�b�E�+kim-r�c*��J�Z"[m2�	Z�mKe�D--��.(̶Z��U��9kF�)-mj�եF-jPu���o����A-��a؇4`��<{/L�7�Ge�'���9�|�m�W���{��9w�V:��m΀L�"�-�*�;0�{?Q�Tf��S�3P`z+G`��@"q�y��͍���ux��R+���s*��rTt3ʅŎ]KJ�[�-�ܢ/��w�[k�A��CA��c��輺܎�d�e���qj�7�����.�=��N�(�xi����4K�f|����g�f���5������%�z��^�x�c머L�:���=�Cm;�F�T�B]��K6%�����,�����ڙ�H�"�s��j��U�t�V��j�:DbO&�>)חL�.���'@�ؚZ	�� ��L��"���]�Ul6y��v��]pLE5�]@I�,���{1-���T���]d���U-���eMXf��{g������h�&"����1rF?hހߠ���+��%Y���61:n���-��a뫙s�f�#�v�^o$-r��No�X�Zs͉��a�q�j��l�:#|��z�~�4,{[�_��їk�8&�},���V$��R�SuHBfм�����q�i�����Ԛ�qG�������/�v"��`˻�h7�7/��U�ǡ�З������3Ѕ�8nq�n��@ԱO<�U�̩�wz��!����[Աu�ۣ%mPh4��9�� ���lP�qU�52�[ӻL;�v�[9��\�K�8�h������e֔f���v�`�8a-�͵����|�92X�U���Uf��^�(�t�nTi<�Y���a_Qu$Wn���� t��Q��W�W.�F{�i�FC��q�S��A;��A�k�K�BX۶��W�5l{r�R޶���u�<lU�+��Qq���������g!�^o�k)��i?f�^��G���e���ì>ٟoc�ģ���������
�=S�a֙���)�p�q��m���sԬ����N`�Y�=���g��Niv&\i4�!ʓ�8o;���!�L�P���';��l{��//�Rۖ7IFbV��o�<��N~�f�m�н<�T�p&Ǔ2�q|���uLO��v,=�J�G���8��s������[>\�v�p�S��\�LP�!a��aPX��o*�����ojC��t��)�̅_gx�eOQ�k�@�
�',���e|י�)yp_�
���κ�hc%;�H����D�/�p���{��-ˆ�����!�_%��
5���;]]��^m�x�X:�����m�ݯ5՞%s?0yxa��ja���:M?�D��e�����6M��f.TT�����S*�TÀwk�y/��>V[�Pl������^�]��Gz���7�β�E)tJ�Ꙉ�rga�-N�Z�l�����QHg[g�DN26���I3�l���w����X}��x?��X��@pͳJ���v;TſU�x��u�&�X_��Q�Au��mȼ6�g�[�����8H�rx��ʁ�],y�{8��O'�`�p����qBh��XC��8�v �PȰ��h���ì���RSЏ{{f�ԇ޸���
����X������]T^8�������ҫŸ�H�vua��VG���z������N��[t�>�LK�;��f���}�♃����
��E�acn,[��Qj���}h&I�蜶��ʯ!�AR��yp���,8i�ugҎx�;u1���ͅ���ɴ ��m++I�5DR���HJ�a�R����<6�S��Q{s^��j����f���\N߭��>0?���+P�R21�y����;U̷ؒ�X�X���Up��B�U�ݍ�)p��mS�㶶��q���,T�U�qm;>�z����oDg�/,j�z��%�"+�*z�*�a'KK���([u�Ӥr\+37CG��,�˷�0�s�Vo�4J����U 5=RA�nj�H�s*,�J�/�����+�������̬��m�ٚ�u=,�9���>�̀		RΗE��8�)��Jd�۬Kʸ"ŕ�y$�V-2.�e�J���5=On��8:��v���ϸ���>P�F3�c�a�������&k��S�"�O�Uq���c���o�T�ȫu���;�3*!��6F"F;HF��dױK�`=�#��$�ߦ?	~~躐�3y���W���r�G�eh$�����o��z��a���AF��㧖y$�b����a����!�9ơ~��Y��	�4aP�a:U�ό��a`����*�i�n���u��V��m=4���I�Ez��-��j�wk��Q8H0����ʰ��X)��5gd�"�ù���

�
�Z���˓;1��{H�K�3EW�	�.�,7�ػ]eL����q�L7w��K�{X�j�����6+�ҥ�K։�YഗK��8߆������9����W��+$\�Ьֱ�_j���a!=�,��I
�VC��r����x�"`m@χX�cXj��L�t^VIm��5Eĭ7�b6��M������3���B��Ԗ�ꕺ=oY!h�;ׁ%ns�V	�6X4ޱ$�M�4����>��<p�wA�1ַ��J��\Ҭci�-yb�Iw('' ��v�]�X����!L�G:Hu��Gz�sܝq]�o��L�兒�������u�������ũ�Ra��d)9���m��7�
��Өx1��V��筐�����B󤖆�M�l[��d��D��|a�,GS�+y�-:�m9�x��lk�0�A�{�=�/oY�� y�k��TmX��dz&�p{�cP{=͊����R��{�z����v1��ٝ�4ϫ��3��,J���TxT+���aChe^/x�<=���y��U��!o$q��d���(r!��%Ӷ�v�oplXx��V
[h�"��/6���>�(�/�b&��625�R�
T./��MS}�ż�ܢ:h��]�TPP|L�q�����4Q.�&8��qf�[f�\pR�E��>����Qb^q~~��3h�6Q�����{Ƴ���"X��U�!~V�O9ݗ�Z���=�Co���#&R�B"j·e�x�%�D�h�}H���īa��}$�{Z�|�p��QQ�6�u;�:��u�����$W��A�g���G�UC����S#��r�'�]��N/�-<��:����@�4�s��7����S��~��Bs4R4]O��s(λ��z��[��45y��>��o�"{-fN�z'b\�N�%n�w�y������t��1��x��xE��d�+����XË��0';����]���c\����E�Eq�^~{B�/����9-qx�SVY�^�D:o&��������ű�z�F>L���'��8W��|��E�V�nW�.�Mb��j�ӊ���O5�89M�����Q����)�F+Рm����u]��oq݈�y��`.�X�(���BIIK�A��"�sv�y��׌g�r���}��.�p�ay�~4{��������#�K��YV~Ax8��RMjb���!�N�ss[��[������ߵ�7�-Y�D�L�a_9*�p?+^�E��~2�Տ:�� �*q)p���H�9��±�U)\�����a=��Qa�h9�2�%�~͚�6�!��V0�z��X��;�	�~�)_��"����c�g�g�{�b��SZ%��@]je��Mݲ����Z�5W�GC���r�Y��L���Qr���`�ޗ&��%�מ�Us7�gӛ喢JBV\"zrN]�w���z.2�����{�t�g��*t����}n�U�,w(��{Y�hZ�)��s`��KX�)�)-�mSJ.��:�Ǔ����B��ۓ]!���]�S���93�k����s�>�Xڔv��~��U�G�p�A�W} �C��2��Op���%ĉm�lt���賸�� k{�e�xY��ǰ�U�����LFWK������.�!��1>f�ذ�-;�GBe;[yK�XwErT�8b;e�T�3�K���D��B�al�T���!�z���j�1��u�2�#'o[2':�{�ˢW�'A��∭/E�Z�����P�d�a�u<������ý{~���ۯ
�X�E�s���	a�(k���].^B�LLB{���O;��Y��|��}[��]C�.ͻ��^S�S�5�D�"v�<��)�#n�e�w�[�%��v� �����l����vz��-�Û�|�'��'s�9n�:�O�o$�&t��=^f�kVU�C�뜕����Pȿ�Br�6%���^�v��S�g(���H���WU�bƺ����c||:x��'��h�+���n�ٕ�;6��ĦUCo.V贉�ߺ�Yk�FO��I�	B3�v�=���ס�z|k�'�����V�dD�'e�x�u�v*b�^\/��!�������#nx�����I󫳇�IR��I.\Ko���%�u$�^�^��L���5�Ҵz�i8����cz{T[�4u�݃��m]���EPV�Է �ɣP�uQLa��3;#3���e�_qʆ� s6L�4�������]y����6�b�2��V���!(cJňvV�mQ~x����4���<6�t��5/��[␥�ϭ�i5�&������3cȱ=��&��(�.265���_^F�/sҳm���\|.,����_�ʊ��b/�v2g�;���D�R�t������i�G����E2��O�-
L���%��j�qlŬ<Ic.���ņ��,��5v�{jX���.����>ɂ| �Bь���<#�]-�c�M��S��q�W��%������4�H~nV��C��3*!��?=J�uTN��%c%q��Eݾ�ވ��58�oZ�7�o:�����2�N�bx�(��0IdL	
뱨��^b��Ggj�8q�>t���?#�Б��ZvG��τ~V,�Dt�z߱�Sb��zk������� ✎���z�ߞr��w���u	�]H��s%�uI��/����� A8���zux�y4H��<n-sxXy.Ȩ�sQ�^[^;�C~��?b�=��}�&[�رn����9�>7+�󈃕� uA ����߆սU�+�zU^Jũ��8���<Mj���p�ȭ�l�n�>�,c��}@_ ]m[W
���rݪ,�ɋ�!�i��za��uk�L]�ul�0�X���au�M���G��B���M�bJF%`WS3�\_�&e֥���>�V��l��ႍZY��]�t}�E�]gmk�Ƅ?u���BD�J��Z�i/��G�o�]�4,����5��k�ټS$���gOS,�^��F�>䐯�d:��g�~o������K'��k��*�yh��z��5�i�>��l	¦� ���֨��T��4\Y�5��?Eg�w�9wC�/�:�z�4�^�T"(g1@����7�w�Z�P�d\6pj[6�Pb	���b^'f4��b�r$V*P�gh��v{y��N��	�3ĸ�Ȋ���Oz�{~ۆRw���{3�Mhz��	���c�#������8=�&Gc��ج�/�Cؚf	��������\]%k^����3���%��*<*߸����*�[;EC�I��
^Wd����k-r�J��=G�q���{�U�G)
P5�B'��v"�2V9�������n�w(���6J�,�qa���h�\[�/�(�C�[k�A�����6�s�<9`�`�{nA39��y@Of���l>��ί˒�u'�G�Z��s2IamH�0m���(��Wt^E2�\1��(SY���ݻOp�L�Y��)W��l�l]W��>8o�물�U-8�V"<��3�ꂱ�핢M76���v��޻ِ�3�p����0�'�゗J-�O�,'jfXè�ԥMP�]�$��cg'���u�VG�a�&�s�"rֻX��=�#x�v���qT$q�U�r�(���I��2aC�j��L��(��N#�*��U���w)��*a��\L��{y�H4}Y��Ym���Z:*\<���Qh��}gr��ɔs[~�4h�9��y-�Q{�S[�gԲ�����A� O�&D�÷"z\�\U��	N_���^�����ؘ]x_�Wya�9CmK\s��L0؉��	cp+y�n�a�Vc�pzK�h�w�Rd$�<��W�[!�|���������8�uvX
pр�m�w8��܎n��ޛ�m�3^Qܮ��yK�v$�	K�M�!��<����7E��m���$�"jj�b�4����)�0d7��Rd�bx�mf��]gz�-�B5�Q���=�u�5U7��f��ݹ�a�l��P��ȫ��k���+�pՏ:�� ��Y�G�
l<�������P@>��3F�u����=l�rT#��B�x�І"%���/ɼl	׈G^˥��7˶���f���ۧ5<�x�9A���W�v�|\]�v��j�s���F���������(r�m�JĻJ�R�8�v�xXk�Σ�Ɂ�b���!��Xt�)]��z��ع�o��֬R�ڃ���ul��o��i��
����W�f\�Ԃ�.6��%w������w>F�J�N�؊��x1Q�s��fMB���8�Y��3s�Rzz�.����f�F;�U�ה��m<*f�}��Xlr��:�u�up�*�B���i��S�,#ב�qZ6��t�t�]�݄槂l����
�-X�˴� �]/o��U���Ǌ S�]�=Ώq��.^d�mLYy�6	���n��J��k{�
#�e1�CQ\�|;�g��L�B�����T,�m2�-TJ��w>��v^�V�<Ά6�:R�s˥e��'�o�>��(���'wc�Eb�Rb|�sG�@��Qܴ�>�9�u��ؒ�ǹ��$���_tr�WM�pq	����;׍��f�sh�㉽�i+�Y��u:��j&�YڕM��
���G�m��y���i�r�X�X�(�Wql�J)���3���r���nsGz$o0��!����oov*a�t������Ƿ���yBWN�j'�Δ���"�����.��(��,U�8��gW7e'�;�3/� ���vR�ʎݚ�i�DV`/Fm ���5�4Y+F/��vd�3���TX�wD��Q�3R��{ёH�dN��l͡1dv��|p�[Q���އu��K�SE*O��s��7�,Qj%�J����ou�IxHC��Y04�ኋ˥��W��q�������3�v�����|p�h哝G�wc)LX�k�Ծ���գ�qY�W�X�]*N7����R<8���8v{۱Cq�y�	��_�d�Y�Y�'�b"�m�E��������x�^7yz��<�+��k\�7��WA��r�0�ۑb�셺YiRFz�BS���I/���]$��-��*�^��nRW��nc��n��4����r���9����j`��ع��>���ycE�N*5z���%����V�_Ŏ��{�V�r��
�¸�3�E=ώ��2�z�$Վ_Al�z�s�\]���	ڶ��%.�Y����U�#N�D�va:�0s��B27B���d�_>��mfR�^`s�j��fȠ��Vءl�v���Uj���a�G�:����蕗ڄv��V%X*f�2u��J�I�y�!.����3u36��_��T�f2�{m��£�8���F	�.I0�s6vf-C�YV)��!!��w�� �;e��K�hTI*Yv�kP����n�E��nA3N-\� �ܰN�X�,f�#�����m�����Y�4��*����wE���(
�I� �Z�KB��m�-�*�����KZQ-E�V�T�Dh�ѥ�Z�F���D��R�LQ�DYiR�b5�ID����j�h���j�"TE(�T��2��b6Զ�F��������mZ�*%�ԴV2�[m�F2ҫ�1���(��k���iU�ڊ6ֈ��)k-b��m��4��F��s+�ƣ��E,B�R�ڭkm��ZТ*�-U���B�űikJ-YBƍJ�-˘��ѭih,�JXT����իcr�pKE-+R�m����b,m�e,F�X��Z��J%h�E�me�*�ڵ,cZ��T�ԬE�-�����m�QJ�V�TTm���ֶ%DJ�T�J6Ѣ�K[Fڔ(���KJ�A�B���m��KJQ�-A�-��+-�ڊ�iJ �j�kU���ZҶ�ī,�����)kbZZ�J�KD���J�-j��2�>��D�������nv�\�+eq;�i���<�ם��5/�zY�����ޥK�jS��:��U�g�	�+���m�ؖ�H����ҳ��V��`'�:j, sM9�2�%�y�Qü�ec��ʗk$Ͷ�^]�	��Y���]�wO>_�0ӕ\�򒗝aq�
���S=�C���o5����_���өk�9C��Qr���`�m�px|�aP~7r�]�u*T�E��_���1,�f��r4'�ڌ<�i�
�ӏe�켇�g��fx���{3�ie�+�|�9���7��fB�2W���sW2�ƨ�?pY������o.�tY��V�X������+L�+�e�cqHXl-�}�����-	s�^Y�y��y]��l���V]�1"|N�V$��_��<"����.6�U���Ί��8�9�]n*-���BF��*c��܈�P8D�rzD������!�c>Hg�ns�ʽ��ITX+�C��ly����y�̿[�'+���X�� *ѽ��y�����qK}@��B��zlt�T9���7"�]�yn.,:�N,3��y�!��>�PRcrs�F��e.�Z�f����L7{S�X�ܮ�|;�U�/X:j  �!��15��$,*+���n���ʃ� ��ɋhm�yj��q�g��������mej����t�OD�i��
s��J5��'|���r\�:"B�*��0e�fOjŠ���&n�^��f�P�GNM#�뒭�H3T2/��F��=6�N�ݬN��Fx��/[�.�O�r�d�%�bƸ�qA*��c||:Ux��UkP�샰g�:R�%D	�n>�%wH��z�Yk�F®�p�<��ۖ)<흧ܩ����<I�9dt9i���(IߟQ9bv_������&��^_��X���y׳j}4�S���墏e3�kU!(bjňvV�Ԙ�Y����т�͠:���37:��:�ZȄ��T0�^��a
�1E����ω�E��;<�����>���FT�<r�:B!�s�:����E{T�Xð�ePQAs���J������ ��U�y8�Y��L%�}5W�N����8Nt���gְx ���<)��bOj���/n�t���R���{�y�L�(_��}<�\"k��,R�65ӏF><����^T�u�T�p������d8ݺY��C�U��9|�������i�; 0��7�{L�#M:�^�`�M�Yꗵ�yʶ��k<�L]̜�9�NI�}{�8n��Z�H���������5��lJi�};os�u���86���}.��ge�W�lN����iL .�᣸+͓%�zj�է8�a�%w_��V�i�O^��{w�����[F�l8���`�^�k$%�9P=���"ZDCh^��^L��)��ƣ�T1�W��x��8W�0ۑ�l'��>˘谺�
�rQ���9�::�3��ؿ$��Hr��#��ؠ��@<�u�z�:G�ziG#��,�SwVv�'H܈y�t�8�vAP&�$*#^M�;6s�Ӑ���iǒ슈Ꙋ,�����3rJ���pX�s}@��G�k�GJK�\T&���gf�]n��E�����{���g�X�r��/
yJt���4��Z��W��k�������y8�NW�\��mN�7ܠ��U�8Th�.<w���9��F��[�t����x�a��Y����+����U�X�^��ņj�	�Zls���\,xJ�5�#b�Nz���o@��3smx]&׾g��I���k>��_!@�I�~�(�|�#b���49��RY[�-w��|��*�Yw"}X��͝��^��7��i���2��i��X��̿L<�m,�d�}���尻Wz(�=�'"���h{��wG��-�ގ`��1�z���yQ=e�� S�@k���wX/��=Kw2hu�ܕ������%KF�f3m����O��&L�7���ȗ�kD�דJ��3�Ӯ��v��+�h�=[w�	��*�2���L�C�4���l���Cjf@��(�
����\�z��PC>�ҙ�<�qؽ{]F��0L��Y���x^�G�f�e�WӤ,B�����Ł�x���q6�����K�nGm��þ3XtI�"��B�����l��;�v�ɮ�J�oh(u*�8�r*7��-+mӎ��������r��ʮ��(��g�v����|<�Z֚�{�x�θ�%ҋ{��N�(�K�N;�WBH8�H��3ܓ��l����/���.Я�)��m(�s�,�ż8DEY�5U6R�,���l�8-�]�d�T/����˳<*��'ޭe��[�!`~l���}�<�ؐ��֯�"m�����z�C�R��d�7�v�J�$;���&{�N\�L�r*-cw�n�Q�xod�'����*ܢ\Cw�--�5��q��x�qa~+k��Yh˳����5ae8��½u�GAh�o?7;��z��ߢr�����vޅA���u^I:���1NP��B#l`($խ��k:]�B#�b��ҥ�J��7���qr����U8��S��o����O�c��v�e���W;�. �d{F�c�ħwh��BE���g:5�<}s�^�'Mo:��i��5KNy�5-���^r�9YdP�eb�+�a�V�͹�����p_���k��+�׎�>���M%.��Ra9�xXN�6�x��*Y���7�z�|�q��V�;>�@�8�9u=���{gY����I�ă��꼆�<`FW���f�u������ﻐ���D%q�l�j,�?;5�++��ǵ|��¦t�OLP��Y�r��&T�V�2Hn��\��[�v+~��abu�ϕ��_B�q����C�+�H�Ҽ�s�R�n�H�����MY��<��s���s�bc���M�F/f�����)�k<I��,�&⚡�WR��uZ"�e
�]t+���d&Q4�N��V�]��6�+ �qc�׾uv���{��eƓ^�$WHB*�"��@�k���FΖ������ǰq:;]xyj��Ȣ��zZ��<�7>J���
�� :;��˼b>�^���
��H�b��N�}3�!v6}F5�jPQhI��z�Y��L�u4z�$r!<�M�g�J�*�
�{����K�k$��L����
Ūv��pQŋ�Tbd�乇�WXU�Vvd����f�jP��+�RHL�����pp�b#C3a�����b�m��T�M[Fc�^�#�}}x�R�oc{�1��lܜ���/��:�#�]gt��5l�1�I\���.�h�,��V��`��F*fR�P�uD�[|*��ڸ�{m�i!V�e��.�����3OcS�]��ޠE�C�OWxPU�t�����c��]�˰\6��Õ=��*p�����+��;t����qx�ǲ�ܤI�(uW.g��]��\%oj����HLо������N�j�[ڡ�qܻ=x��\Xu��\"R͋�)��7;KS(��$�5����帠�\�٭!Cޜ��X�PȰ�g���\��;7;$���&���R��U�N�$i'��KRᎨ�ca�ʳ��됖�ͦ��6��J�3n���T��7� h�J^��]���I.-������vxA����v_�
�د�Mۢ�7ކ�����¡&�Q9A<�FL��T�Q��N2,Jt�m���N�y�tr��|�sz�]bj�.���j�u�&9��)���&��ܿz+Yy��o'�9Ɵ���Z����t��03��k+�7�Z��_/U�oeˆ��#o�00��L�3���Wgw�pKIR^�(�u���4� ����ЇLڴy^�:轮0�Kt�Q�f��E8vMqG����s����(A`J�����˔�sҵ�kn�^�[}πZ���u�%�`,u:�Æ�d�ꋵ���/���\^�7��
�v�Z6;��6\"k��8�"W�-ũ�R��w�zz'�=�c��V	U��QP��s��O?S���X< �tv-�+ukU.mާ7����Z��Xd${����0O�)و�>���PZ=�w˳����cA��%]�p-�~<���孑�K�5Fc��(�=0��L�oU@Y��ƈ&���W��D�l��X�*{F ��S�Q��v���o�`��3LI�0�w�D'��pu�u����/�ꂱ*�5�\=�>�(<]ur9}��ϲ�:Q�h^��%Y+�l��g�Aq�D!- �
��y:�v�/W�zπ�.�]�\C�P���z�%��ע����t�Ԣ �q a�	>C{(��J,=�.r�TF���n3[�}s�ڤ��*��YK�϶�Bd�'D��W"\u���7y���mj�{7<�Z�9���
j2�C��:.���ĝ�I|j%u�̿�.�V�$�޳�0N�*�<|��!��,Y���F;�s��{�yr�:l܎_'f��L�/ӝj�6p��Q��%��z%����t#Bu	��u�N��	ncN:�6�.J�R�{�6��y�v�;��|d�Q%:\j��Y��[�k�_����Uμap���­��ǎ��#����ر��Čk�e�9�����hF;�N��b����ɁU��bMw[fb٨Ba��:�� �5-L�!�1qy��L����K��Y���Z:�h�W�a��?m`Xࠤ��e�\����{0׮�v��=�ϡ~�����R�52�{����-�QB������X��;y�E�|Na��J�~�έ���v�j�N(r�՝�ab�ٿ�,Ƹ;+���-�J��!��r����+Mgc)��-o-(�J��1ۭ���#a�~׵�j/�aB1U�Ey՘ ��)a{<�]T�wbj�o.1u9	�wq���X�5�ϱ܋ފ��j�[C���Ӗ���R����7ݘ�@��<���.�
R�`�m�zV�t�)�LlX|�o�U~�����l����"���LP���+�qE6���3�q����D�6ӷ"b�!���&!���/��,x�9).�RKG�4�i=��̬6�F�>����lz�M�Ď;�n�9�G�M�������}��b�ù'<&�%ف�ybC<'��^�[Yd��]�"�RX���J=���B2SRV|}n^-^��W�f1���r5u,�wn�v���ُ�i{�C��AM�νX����&N�{ֳ̨�a���d���a��;�f0��
�f��˳<*���>ʄH3_dAc4ۛ���3k?+����
� �I��f%���3�({}R�{�G��U�x��^��|l�Ou�C�_pp\T7�^E��D;!��D9D�5%i�K��i$�u���63�IC8�*�v�#��˳����5ae8�7Pa�Ho�2���c<����.�}ZrR�~��b�q@Z���󮎌M�����ؚ��!ƹ��q!U�Hʠ��J�A}��\N᢮��֥3��@�d��w��bI���V�R��tmw_cK���J�=�x�Ǹ�pLV�2��W��X%��,����.{p��j̇E7`�'�:�Q(p��N�&�/��ȇ>��x��|���kШ��4�M]�#6�ཞ���;�`��f��uKy��n����e.��\"��>�3�[Yf�`sJ�"'ug�����C�Y9������(n�	��ﯥ!���)�B�F��0tK���@* �l,��D�6���.yZ�;���Ӓٟ4D�����B:���|��°ǋ�=[���y�3�5*�q�k�M�5v���d��V �^e��:�[�,�Q��\.h����b�qp�����.:,�x�q��K ڛ� �����z2�L|��>�u��B�����V'����	�MzڧeM�A�����\�g�4|Gct��gZ��D��s.4�ؑ5����E�P9�'֨Oo0�����-:AV��w��7�Z���Զ剜�7)+�/.��|�x��v�w��}�����Ŵ�9}.�O=�J��ӉQ������ΏD�;d�C��ҟ����Hwʺ����8��Yf�v��Eӽ#=�݃��3�v�銄=HBN������Z:S^g�=���~��5�`Ka�Jm"y��T���yf�EE���͍��_���wt�`�OW{�j�ԞkP�T��uMS�`�~�tTX�/��8[�5}���:r�۹ؤ�aײ��G�z�d�~²-�;�_D�W���r�.�6R/���#�7V�3m�x�egj��{|��F1ӧ��t�V*�����EW<vhi
����N&E�֢rݗ/��ˬ�*�\���U#t�*�N-�T��ȍ%�-�\1�bƿ�����.���ׯ�S/)��h���o�9|�u�M�Wb���u��	6��Z�B/�h�%�5�Q�wR��J�) Us],�t�����K��Q�����������t��}BdI�ĩ�1|�%$���������2[W��1����]Y�E6qw� �6Vv�v%+�}֐��}| A�X�y��n��#l�|����qZ+oP��D��Re�B��H�Jm�
{�J^�W����!i���U��H�ɍ�ͣ���<�sZӤ��<͗"�)�X̻;�{| ;�&n:�Bho1�K���s�['eK.K+���D��:q�:h��I�ӬR�Y)�մaLCZ�P�[�Lnɖw���gf�)T�^���o�y�Y>X��ŕԳ 	i憍��m��[Q�Ѻ$�d7+PX�͈��md�Y��]�ŏ���ܰ�7���PH��H_f����-�N���(��]�c�T8dvef
8��x�����Fܰ�Y��qQa�����q@��Y�e4XU//ܖ˴�Ȏ m���y���'`
��#Km�ѧ`�]p�t��1�st�n����Bn�X�z�v�L�"j�QMd@p��YW���zo ׆��[�W\�&>-�A���V��`����^bA������oro
�[�M�u:½YH��4�vM��hW���h}IX7���\0G�݆)��g���:�coX�s�X�@�Y$�뇛�,�K���|��֞�5虇ڦ�W�#c�h#ZV9x,Č׺���U���2s6r��Ԯi�NNq<Z�mWwZ�[���{�Ny��B��Ŵ�=P̢��:��&xӡ�}G�kt�V��+�)�d� 1���Y�8P8��8$�ʺ��(�Ƴ�S�7��SP���d��X��#�c%91���Ӂ�^8��}�.5	���&�Y�7�묋�k ͡=�ƥ� )Ԑ�h���7����/�_������NƋq�j7���X��`�0+;P����P��I�C�#�]�q_G�J��Y������rX����j�#d��Q�m!L�FwM�F��k�i���n�`���-�pf@xcw1�!��$_]�0�j�1��贫j2���h[�R�������M���S&;�/{��\#p���)��Fs9��;��B�[l�\]M��<��@4$�3��+aȃ�h�m]3�"��'�X�)dD>���#�+��j�8��X[ZG��,7��wo �Oe2�4�i|��|��2烦\3V���{f�&<�p\�4���+�i��)�[�fԮ 7ר�ٛ[ک�g��Z�u�-�sN���!�P����ǀEP�4U9`��CϦP����&�!n�.���϶�HMjux��/{;i%�ٔs��u�mw{&g��1TTi�YU95�����,m��c�X�{|R=���E�YG����^��m] .�""�PV�mD�
�U
�iZ(�����KklR�ԪYj4E�"4��--�YU��[l��m�J�`�hդ�`��؋j�B�b�Z��iA�)V[V�V�+j[-�E���mj�F��(�*F��U���
�F�������lij�Q+ik+mb���V�m�%����F%�-T��-��օm�h�V�ڕ%mm,Fҭ)TDTV0m�ō�������P�����%B��h�J¥b���T�����D��حe-�+*�*U�,e�U���"��e���J�-Z�֖�+Q���DeV��YKj�(�R��m��R�E�-+A-V�bZ"�U�1��%R�,�VT�eTJ�DiD[V1b�,m*Q��j�*6�Db��ִm��m���X,TEZ�imkhѶ�[U[e�-h��iX�҉mcl�PmV�RZ�U��4h��Q�V��V��UV��[F�iKcU�QEi*(�*��"#liEQ�X���[AEDYutָ�o6f�ӟe"=zfK�}N�X����S��G������N��o{��j�(2��-�v']��ζ���C��Z��w�Z����Wv]ӫ�^��<�I.�g}.z6�T��¢C���¨���|pU���!ix�IV6Oq�.76'
������~�-��Y�.Tf�Z�Sq&o������~��l����;��LA��&� :+	��������������-]�ζ6�u�$�'8Ә�xJ�l����b6+�M��Q����Y8��A�3�KAru�s�9[L��3�f��B�H��qxLK�2�஧��S���x��z�,2܈�:^���_vb�s��c�^��<�QP��qr�_���q^#>���mh����z���;N+i��ʖ��!2��]���F��9'(��]�P��و�V]p<�Z9W4����ܸ�:�
}a��-l�֩��q�t�%`�Hȡ$�k"ڧ$�ǵ�wR�i��J'p��a�t:XR��c藽8�p�g Í�/%\.���7��_�1���|�Q1ّ�K�&��.����CnG#a�J��>˘���6g����OR�T��ÜBB�Xp�:"�`���F�����smWl@J��j;�B��EaU�	�`�ǣ��)���P� �~�����{rm��2�۬�B}�ÓP�j��h��+��ggWxw���u�N]\$>@�@�se���.�ַOH3��.' M��xhf�fX	����	ԋ�h/W�s�|�t�4T=ȓv嚭+2�w��E��_�t�'R���Ŵ"����ʰ�C5�ԭ=ӽŚ��#��m��l��&�����EGQ�/���>ۑ;Ȏ%�-)R����61��|�a�)��ټxj�u#|V)~�c�2��0�Q��r�S���$�pQ:�f]W]�_ft�ղ�&B�P�@�@fˣ=+ǋ�TXgZ��q��vG��<\=<ʞ:�fM5�͵�#-����?	�^")���H����0�a�ĭ1�b3Avjl�z/ɏ*��F�ꔚ�J;��/�Z�=b�o�;DVk�$׳��i'lC��z�z� �j�llz��}�{�ۑ
�j��!�@�m�C�<��\��P�դ^�;짤�䈪�݆�͉C �v( 
���{O���1
��|;�����y�_S�{�e�o+~��"7�{��{�����IvF�
ggy����o���׵�j/�@�4-�"{�j��C�j�˧jM���kt_�m���j�mZ���Dh����+iR*�eh*.�Y�|̺о<�)���_<��Yz�6�7�G�>��޲��bjw];'��h�Ҕ���A=\��#WyF��aK�.]4�C���w\�U�c�Bα;�ޮ��v��>�L��҆S��nGa��t[�r/z*�b�K�\�*e��ūP�Ŋ�n���hbBm@{C��m�z�S��9ȸo�a�n�w`��63e;|;��Ϧx!l2b=�Up���T�œ^�ȣklÀ�K�
]-/���bQa��՜ÿQ�KЭا��j�#����
�o�I�۪!��Q�`��b��QmW/C���X� %��s���pk�	��a�֝ܳ~.L!B
�f�3*�.����z�A:�[ɍ'K�mg�W5t�H����º\�p�8L�j"���Pzx���-��8��rn�Z�E���t�����q�E�Q����U��9�D�y�w�xWY�Xt��Y�����#� m�s,�Is��/�d��s�oǝ{;U���g#<ʊ�VS��e�(�@w@�FA��'-��*�2��9�NauuA�Q.+֤��]��	����3��Ύ�}���t�ȹ���n��D��VC�h���#��g�����ώ��y�T����WpZ�=�����Y�J�Ԯ�z���rc�ޞ�yP=�D�^%dWx��h�"�L���iَ抲���;�
�b��7���i�gH{T���M�]�Hⓕ�d���jY�N��+]������U�n��}��؝�a[�O��4��k�Lg��m�Z��+���L��lMY��7��e���q�.���kN^b��Ák�h�����1�*��" 0�H�_K�����xE�;]}��^�5��-]�:�w֬.�/ة�@N�df4��:�߂{s�����4\�dhb��h�^��Wm:���2N�c6j>Sp�Ǿ1���FaI��_=X&,kޛ��<��ش��>n�lޕD�����R�m�	��ꡗ]
����!2��j��U��SSv�۱[���xA��N(E~��6�~Y�d��a/��T�z��A||u1[��ޖ��KN-�zfL8t��w��l�R~�4}�u��n|���|x�`'����e���~�݁��S���Խ��T�|\��>��;�|.XQZM-��:R+G�?0:q"�.�i�{ѳZ�J�wy:�!�n�L:`y>R/��9��W��O�(�Ҏ��O+<O�D��LRd6{�X�Ji^J�3�d�e��3g���$�Le�2vȨS�7���^̊�)ϱv�kt1i�Y��s��'c5XBӗƦ��y���QZ��4vic��8��F�r�$d� Z��=rF~׽ ��1�w�x�T��޶R�uk8��ʹY�MqnRV���-�DM������S�ܱ2ʡ;�c�rl�7�]EE�\�6N�-���z����������I�����OZ��I��Ġ=x�U
��f�o4*�W���N�j�9T3K����I$��r�~�?t�y~�R-JZ0B@���P�K "��6%��ڽB�X*g������v��h�����t��I��K��i�3�+h��Di-yh��.���c]T^8�C}�A-��ĥ�{jv-4�a�j�<'Q#A���מ��r�..�ץ�FՊ� ����8d�-nE�r�3��ڿf��/�5��&��*o���˝����W��LYOӺ�3�L��\:1'�o�ÑT�,�=+�;��1CWp�&�T`H�;�YL=0�"·�O֝wH&'��qՒ�f���Ez��(�9E�5���lV'H��q8�Y��9S�%��s����k����0�j���:φ^�1�;
T-Ψk��faO5U�Y<̭K��x��\�N�.@�=�j�z�g�j)�ήX��ʩ���k�ݾ�w��2�Y����[��p�R۵C{���f�Ӻ�!�8�1i�]�cA��*���a��ܯ3��{��˖J�蘴���l�S.����Ս@9|Gh˴A���]&8�ݮ�f���8��.r9�6�B������ނ`��"��r��Jx��9�)Ս�۷���Zpn�;)m�_���m�J\�Qu�Ic�V��p�z�8g�C�)�~����Xa�B֩�C���%\`��V����f�◾����ςuo���92q�{fy�}J藽8�=>J<wWYaM��y�����gD��Ĩ�LƽN�uʮ&�)p��0�.���r9�Ti5sZ��1��^�y9Zt|xl�}��Qag3,'H;���/|�H�V��q��=gM�9��)'��k�`�7D���э����u(��W��P���0u��y��\�3�NNZo{l�Nœ�j�Ӌ%��Q��Pv�nDRrG|tv|�xk�*��4��V�='��u�]�5���Q*�
�8%N�Z.�2):!Qp���$��Q%��K�.��
��N��
�n����D���@⡛�G��ű\Zrp�h�q㮼��+���d�7yR��z��~��y�<۳�w���pus��"���&߻�V`3�����N�7KO}z�Y~{[Z/iJ��F#�s��C3̎�bX~��%��F�./�%�Q�}���ŷ��ƺ����|��3��]�Oj-gG
�E<��|BSp�J�>��U����v�o��s��s�͖�'F��+j>6%-|�f��T�����U�%����{�Y�cؑ��}Z��!�^�U�l�;DP�t$��B����>9i��5���Z6S����͡����VmȄ�u���C�x��<��v=�/��ץy��IC�za<ZyH Z�|M�8��G#b��\Ł�iar�T��<�z}��W�����$I�c1��։��0�]d;�*�c5c�[���Z9�bƽ��Q~�rQP0���g�;���G ���/JB�a��P�S���7Ai1�k�E�ؑ{�T�Xٝ�����̈t�L#̝�r0ԍ�t�_��C7�2��q����zVۧ���������ngzZUc����I[>����u*U�&��E[fT'��KN)����p4��2]�S1��~�},K�N,�:rR^�RKG�HV��A�|z�Ģ�Y5m]�sw-�YY�n]J�<\]�bz6��a;�f˓T��ʇt��_�GY؝h��x�e��!jfS&t������'K����Я�,Q��N���1m�O���R�Z��6�ݓ�|F��,�Ws�Ԓu�PB���`U�G6Н㘋�
�-%�ϱ}��]�!�O]�R�" a�h���+עj�m�<��s�t��q^R��h�%l��Y�v�fQ��(2ُ%�ܪ��M���M��}�!9\~��r6��S@:n���+��G(�u�)�ᘴ=3��:�h���v��]
v�cS�³�W`4�����9��O]�DS�'��(���ᯔ�W]��2�2�f5⭫���:*�yOOd;f �S�za����oU~ͬ�\�7/�_n��y�g��⊭{��sk\����7BBөi0�u`+o/��@��Wn�2�SvuWq�ŭ��5ܴ^��B�7b�1��5�xq߸m�]yr��s��8�/�om�I�KF��d��b�����+����3qޚ���x�Yו.^�K����)�bk�Ւ��͔+*�ys^��P�kwޮy�E�/��2v�VN��b�|/*�ȑ\�VJxС�ʏ:Ě�m>�fv��h����5Iۣ;��X���G+�ޡB�����q��ܰ���&�Sp�#պ�|�ã�
��Ӽ���
>6ҋ;9��̺�M�m�U|An]I�_C�Ҡ����<(2e��f��i��:���+L���[����E�$�b�R���\�UrkotU�z�/l��F)�x�#�u�,����Æԩdu��+SM%�)��]v�����}�>�T����;�$[S�U7�ލs҈�V���y6V�:� �ݿJ«���G�P']	c�\̆^�"fX�RӢ��疶�[�p�.�����K��^�`��wY���yco��v&d����/R�MyS�N����h��I�Y��Y���nb9+t]\^�B9.����.Z�~sө5��X⫺z+�{���f�g�D����ºk��^�Ve����7���y͇g���߾ٍ֩^u��(>,�S]]M�q�-���;X����^4�Yc2/�9�����I�/5͎����頦�X��=x܃ת�
/�Ό�W�=
�
~�����ӛ�h�\:��%Yg�y��L���R�����۪��1���7HPL-��1:��6�{P�De���-�ٔ;�_un��ڙ�q�F�ݝ��U�`�u��ձ��$ZJ�^G9�J����~I����[���u���3�]Ǳ���Hb�_Y,Sv���%lo�e[�g(�5蒦��	���Z�i���M���U@��e�l6�Wm�wh�L�>��5�V�6�
�v�/�C������|�fx����E��ז&���Z�(h��y���
z�z�ޡ����շ��nc���'��W-��Y����U��hPV�T*��-�_�u�s�76��ĵ��[Os�f�O;o�^���L+�܏WJMZ���X=}P��7X5l;�P���m�i���:Vd�U�Y]aF]���nd��ߦ3u�]���U�%��|�e7�~�����iϦ�oN���õ;5����=|�PY	'ϼ|��<���s��rlm����mÌ]uW��Q]i̚cy�I�e��V[��;�b���k�F����{i�0�E�_�9@[�a>��I��v<ri��w���r�c9d��<�鳢+�g2'<��Uq=�O�|��Ϸ�`IO�@�$��!$ I?�$ I?���$�B����$����$�	!I��IO��$ I?�H@��	!I��IN@�$����$�@�$����$��$�	'��$ I?�	!I��IO�BH@�|BH@�~b��L��F%�T�o� � ����{ϻ ���÷w��*� PT� �AB� $ *�R%Q@$D(R"�PP� �[�R���R���RUHT%%J��	
m�(� EQU��QARP	EEf�
(�
P"JBJ�R�"���*UIB�%T�JT*�)��U%A$E"UT��=��J��X  <�Ha�[emlf5a��P�eT���F�E�5-E���!��4��b�Qf*aamT����6ձ����H�PD\  �h�cV���Q�i�������PkUIZ	M�"���)�ի4�-��b�Z�#j��� ��BGL("       �b�  ��ѡ�����  .��:    7#    �� ��j�+ ��k*�H��Ҕ���EmcZٶQT�"BUW  q�ej�PT�m6ԅ��V��*��[V��me[X��AlT�Zٵ�l��%J�M����2Z��[Y
������Ip p�V�d�Z�f���[4�b�i��-A64�����M0ԅkV�i�j�Q�����[jm4�I!R���%S� �馨5-klm�6����JPK2��՛Y l0�2�P�XA�XԊ�T�P�**� �]0UPT�J�l���(L�CZ�1�(#`6
�T(j�
�(*�)(�� �@, *�a��Y�U ��ͪ��i�����R�F�@M HAT� U�\  �
г@�l�@��A��iX �i &�(c0M���5UT�U
R��  p(+��A�ª�ؙ��Fb���5)�j��4i`̪Y���@    �7�2�J��щ�a�� `���%(bM �hdɦ�  S�=S���P4 ��  E?��4 4F    �I��	�CL�F�&���#OA�	4�&eR���i�#$��N:"�XlQ ���-iR$��(A dFk%����������2�=����Z��K�a�$D	��i,I�C��%�|
�^IV�?�~
�c���$���0!%-G꒤�&���E⤕DҢ$@�Q��.k~X�0+����n9�"���Z��[��b�geZ��ս|L�X��Ui�w�����|���RY�y�]<Z�n&u�	�m����ؔ�2��д�Z'ٛ�L+l(�٬�Bni	edF����0c�N�[�����8x�����ŧ@e�����ڹ�V�%��7�n1,������>(���	�E�}����U�Z����޹P'�����fnCLf��T/e�UԻy�h]�.�j��_���1�TZ���z����k!�ٔ��40ɦM,vZ6WoPCE��� ,HӲ�3 v��\'���77+sY�mMEX�RdѦ���ñ1ld`P@٣�7U��<�q���r��f7V�A"��Cp�O7��8��e��^`GL�5�+mj��������ܥblm�I4�yM�J��%!�Y{�*�MWk/N�+r>��Ʋ�:Od��v�[B�%�٨�=���c��̽��U����Ip	mҗ]�ׂ$��XG���h��4�:�	�Ⱥ�G��`ʱ�& V|�i�1�faV��Ik̸խ�еoܬ�m�U�Jێ����\��7��dڗrf����C�5'��0d�3siĶ�D�줋��ے�� �f�^�4)3�.FkEJZ�*܂��<�V��c��A�Q�����WM���N�$X6�s[�����E����w�X�^<r�L�Btк�A`XU�ĪWl�u�'k�����"6�ڶ�)����d���n!Hͬ9+$h��Z0�Ȥ�R�,T:�zV3��Y��RF��g�9EQݦ .n^�3Z�<ܵ[�L����9<OP�Q�^�'Ma7��b�W���l����P:Zja����Z�Xٔ��T��$:��͏b/1f��à�^��@�mU�*{i6)�+�r�8��Je��bҊ��:�c�A�q]ɢ`*�on�o7iHF�u�m�tĵ�_�u=i�rm)�*L)�C\Hh`L�K0h��SiѼp��YN�s&�T�w����y&�[X,M�1���ڳ@����5[�����
��,�j��.�%۰��c1MoTZ�U��"w"��A����5���e��iiu�bM�����-^H(��j<����d
�%-�&�5�4��ɒ�-5{aYYC4SV�ي<�5JI1D�[�d"�O]X81<S[5�W,d ���shɴl�z�M�t����[��i�-6H'Wb���(�acpR�<�`�4f�@���h���
ی�5��ɛ��S�A�t�+̛x���Z�㧻5=C �p�C3i�7�K+6uu��4�.*	��;RɄ�̨mK+D�n�
�4�l����Pi��)��4**�7��E�\��xX��ҙfl���������Md@��]f�e7z�qؽ�"Nf8�0-�0P�F�p�S8�ße�yAwHf`�"�r�;HK�Vҩ�c�������^A!�{pUӑа����̐� G+4�S�Y����2�ȥ����G�%���1]�yLA�)n���������S�u��p+�2�e�A�ީ�����B�
�%:�fI���U��}�i���-��-)1[H(\�J�����WW�T�?q�����9����'	.���A��m�F�i)��E,�L�e6-�N\�lk���w�b����m�����Ǎero�b��K$��U��7������h��ӎ��v�ST�a�Z��*��wvk�(�C)��]�Z��)���A�Sy ��m��2�,h���4��B�='"(fqn�P8C̥�e�)Z;�:,}�([]b0��NM*�.�Q���"����w��u��h���ZD�l�Y`C�\N�iMy`@K���AdF�^DnF)�ⰶ��(ƴ^m#��4Q�᳸�Q�e�Y��n�dL��L�J[N��P�j���Xn�m!yC��ZXu�}��f�9z�(1X��XT�"m�Ր�̠�T��j,��Te:�Tzj�3oL�u���@�+K�Z&�,�{F�i�\��GpVa�k^��ՔMc�JU��;�ku�J�O�U�
)e�o�n�嶰+��� ���D+E� �G*�%�Q��z��$�V��LX�s^� ݰ������`�I�����Zu�jĬ�-m�i\�X�^c�cL�bKEZ�.��W�	*��%���2򆪶!sr:���]]��T��b`V��h�'bm���n��I������I�xg�C��8A[+6��J�N��d�0�t+��e��w�����u���J��v��&��aW3�傎��V��@:�r�u-�����[Bɲ���m�503��2�&��P��a���X�N�C�ڛ�6��,�Y�wE��hBF<v(@@���Ϭ�:Y#kKM��Y�
��|Y��Kq���bݼuzF�,L�KKˎ��O3���Kn��ƍ�<p��¦&��[��bR�$xY���[x�j��]�%�4�*��(�i� b�R���n�"0U��y��$� ��H&Bl�8.h��Ѣ��Ǫ�)�����[���E�T�t��ec�k^<v���m�eZ[M	V��G��xm*̑K��h��TH�����v���2���z�p�YD��r��ъ��f�E��.	i��:��Z)����0'��Zː�e�1�jWm��N��*�e����-��w{�]Ӗ.�dN�j�x��&������kr�[v//�6��ֆ|J,= *���8�����,#�Z�(��`���ΰ�.[ܛz��߰�(,n��,��Z����*;�
��)�Ш^�4��\�R���x[WCZ���Y�da=D�`'ZMW�[9H��h���zK%�C4�W6��9dI.]��/���C6��s��'�%5����o �N�1��kj�Q�+'Sok��N�E=���k3	��Rǅcyk++����\��ld�(e�v��T���QYv��c;vF��n"���Z�63GbZ���2l�E�2���YP��l�Ҷ�Wv��VmK-Ұ��F�m�����-<a��u�{)��@��W�t�}��^�!wF�)jMg\��%y����)�F�]kh��M-�U����v�ɻ%Ӆe(U�v��U�	�M��7�w��sctuXY�^�r�����r�ӿhoI�L5z�қA+ܽ=��E��o/�e(a����hb7|	����i/�V���kj��[��W u��IY��6o��,�t4���A8t��ԍ4N��E�lJM����ϕѧ�*�-��.�Z��m��^ �h����Wl�.�^^��j�,3p`*�E�J�AhB�n�`���Q{�ȋ�,��|u�IZ�=a7y�+]�^�-�����n͌��(iCv7Ja���zЬ���]������c�� ����	r�FE��n��y��)�ի�����y'zp�3l"����L���f�����^H!Xo�W�[��N��ָ�噇/a!�f��S�[�u��u���QrMՀ]�F�nc%Qe=kf2r��/�q��.M����	�e�Ϛ�>kb��^����Pݲ��LQ�g^��tz�W ��	F���y�޺�j��[%�fV��V�*��Rb�5�Wƞ��k��L�q<�w��.�5�Z.ͫu�����`�7�HSu�m���f]fReD[�7Jj+�N�9(4_�{�I�*ěR���Ӻ����K/tZm�,U��yD���������{����ҋ'-S)����4��6����+�gP�����y}��zM�{�	�v��,"��k��oHڦ���5���GhS�*d��N��K�m��.κ�õS{� 3�FX͋bBܴ����ڷm��S,]ˣuv��,�x�*ӶSƳ1�����b�_�G
ibR�EP�ҵs+)�cI�#	�kj�-+Lֵ�V�n����s*�U�5���U�ڛ������tnne^g�չ����B���yM�UY] �A:	�������jn1��ժ����5�6�Za��k<ǙD7��Wg��'f���ǔ�b�t��[I��.��N��T��i�`��S�m�щ��t�	Xj�WA�br�I�x�<v��&�B�'l�l�����&�:���BDo��,��զ٦�Ts����щB3%�^�S���A�)b)��]��v���+�n��@�Mr5��,�����S^$���`SgN%�N,�u���ݑ���v����0ӣ`�:�t2�CƷ/-�P\�P�A�]�O��I������d���r��-�7kLQ�Y�����.`֛S�r6^�Ր^V��D�S�z�ahhF���kd�$G�h1�"9��)oh��^��(k7T��i�(�]ղ+r�8I�iV� h^��F|���K�ޓKjֻZ���b��hNқ.�`'i�oQ�ܬ�J왘2�9Y��V�*�;hѮt,���&��hq6�,Ix
�pi�b�Z$ύ �����+&[5![� �j�m�nD�Y��X^ѬcI���%*&^Ǳ�/K�FM�w��4���5����˳���1���[J�4�/hV�ܥW�S��x̘�K"��*6�F�Ǘ���`���X.�n���Z�#q^(`���<&��\��ߜ,�*�i�6q�]� ���u�Ŕ۫o����"jL����2��yl:���n�b�ܨ�p\�D[��Q��[�se�h�W�Ἣ���髦�7&^�xKL�&HN��i��2f:�{�[�v��hO*��%�+ZΓ�P1�/#���MY�Ř����n�����GRǚv�d,�sWm�7&������*��#�7�49�� �3\t�ݘL��Y
,{f�d�ܵW�V��E�`�
��(����-��4���nmSyu��J��Yԅm6�Y�-ܼ�V55t�qe��%JwyK+)�J��.&VԸrJr�����`����:sr�n�&��Y�n�밬ڳV"ùa�(��ԕ� �`xM�Ы�@�aՂ�&!JX���ee�l�p�v��p�`�5��,:XW�wa��B��67KH�]e��a��G�g
h@��k	[4�y�+W.T��8�)+)��6E
�*k�S%��h���nXl�������Rۨe���ref`fV ��Ж��ؒ%��; 㿬�sE������ބFF�PU�Y϶-�-]�i2�ʑ[ˬ�� ����V�i�w��*�W�]��2�h��Ǵ�X(���Z��4�7wf��x�����Y�עƋ�v��OZ�E>$�YhqE�^��{�q4�ή{�sJ��H*�[�������B�?mfѵ��W���`4&�Mm$F%w��<4n_�ޙe���3S���SVb
�N��ז����E��6S��efH:vn��SXs)���D�[b;G.�GcŐ��
�4s��\�m&����/PvA�A�F��Ɩ��`�T,"ILG��h��òM,��ފ˗�NX��������_Ѫ����JJt8VZ���o���&,-�������Pd�i��>,F�o��y�N�E)�Y{���sD�V2V��7�J��@"�;�e�L9�k������;-Q2�}*d�ʔ�y�]��{��a�-�<i��ӳ�����v����*����j=�z�t�9P˼��}�q�8ƧH{k4����xU��c>�B$��5\��шq%_O�[g4wA �WQ,�֜�p��d8�7����Kث�;wkّJ%`U�+�Y�	��Փ�z��S�[��d0r���j�+������v�'o�9��I���r�a��J��:�!��+g,ʕ�+��|�ڙ�"Wo*敒�l록��IS-�+.Ժcnu;��*�a�Ts���
�)*���[�9K�7L�ZhGi��]*�ҮH�o�&�:������'��V:RӚ���([�Wd���tL.�4�P�p�t�BX��Nw�W�*�u�#)N�j�1vյih�G{t��Y(;�q&������b�:�I�[�f�fۑ��U�Z�����2y7z���j�ZT l�[Ά��m�+�Yt�4!��P���F<�\e=ýD�����C���E��;�%�#��v��Bd_n:�ֻ��Λ3M��&2k��t2��%��b���X˒Ų�ǯ)��}�6�Wѡ����G9���6����[3fnӟ�h�;s���U��'�+�n���q	הhJ��yc+,�/e1���-�2��Tm��+(]�����Q�c�U�;�V{25�T��IN��\X[��.ghC%ۭ�ٱ啚Sy��Їi��h� �v��J���֨[����/� ɝ�<�Nu��(���D&�F.�Ig螎kr�#�'K�-*՛�ev�?>���k�|e-,��^���YK�R�gbJɫ�}�a���  ���>���:��C%�+��U.��{�c�i�ߗ�����pm�$���L8�=���/�����hV9T�N��]%Gv�U�9�a]l�ثvt��Z���[I��h�@�����Ƴ��Y�eqњ&"/�h,8�%0Ë�C�L_ֽn���~1^x>��[�ԛMl�p�&]�5�g�gI]ɪC6:���t>krvS���4������>Cr���79G]��\�������S��J�ە����6����Hn<�Jx��{*�mK�)��koy��v�cCPù2ә7�{&P� =C��&��6��K��3#U6py�6
�>e<:���v�QG����+/*�����nm�
'u�CrSx���CY�J�g`[f�i𫝢Q:�-�۹��f�\�HJ�w{��5w�6���Fbj،E}K�q�ZV�[�h��'���SE��u9l�c�bo�%�m��䷤�Ļ�K6�΍�F¹�!��8�Û+�_7����*�MΎ��¬��ѓۗ3dK,tQG�;�]՚8��Di����N���[ٮ��K�>�s4&0�8�׸n�[�Aڅ�tk^� ���� ��nY���b�k	Dg�P������^.@MSo��NV�X|���CF����)�����#����TT1H'T�UaЅ[U��q�y`���ى5�J��><�}�#xU&n�䗽ʎ�[p��@������Ic��<�Ԛj��[�f�Yj��Y�:o�W&meb�_e��4soL��H����د'	;�2�u��J�D2J�(�Jq��	Yj*�k���ut�4��1�Zj|�-}�%�����"˒����\S��8e��.����R�Y�be�X�4�@֧u}�ie�xR��v5.c}�eJ�۷2�������-��R֍���s���B�20#T�:`�7�4�����YޛNA��x�ʈ��NE���/�9R�D�=G�`}�	=r�� *���ZR��:/cwYY��DW(PČ�tZ��Xк!g�塺`ޣ�ħzp5	���^h�C.gT6�"�r�<�`�6Z��N�J�<{_W��i��0��DzX�cyaK�>���а�N��US�Ʒ��zwp��lm�[]m �7O-kPȃ8�4�T���t�'�|����V�rJ�,��	�p����%:M��w4���ikU���+�@ -��V��7�ޙOۣS �!cV�P�g�^�s0�5�]HNn���� �{��Y��1�@�3�z[�����ʲݮ[��)w����Iu��o��ǻ��b�H�(�<�M��K�:��;N)2����^(�+�r���d����_ZZ�x�ՁNaP��˗�$O:���Im3�w<��L�̳�ϖ2���q�%������B��/���3SVw]+�6soK��j<�Ce�&��"�+p�ej�v�u1�����X�6����+�k(���lW�M�Ԝ�:�� �gjܬP��(bD�V�]��'hV�����$�8c����XDq��G��^i\���Hxn�(���5�. ��=X2���bRL�B�s�z�� m�젫 �nL}�V#�r�y1�n���t�
�)�RI��D�*>W��=�:^�}��7ڪ��æU�R,�הw/�]����)*z9��N���,U��4l�\�]�gt��Acڴ���g+���ZYKoY�[�F�񳎧l|Ȇ��ԁ@5J��Ŋ����I�Nwuc�m�Z�>���*�D�,[{b���D�}i��{@��;�7p,�d5��w��utU5���;�*;)n�����\���:g6�9ة�;�顭��M��W!F�4�����1�s;!�u�����A��wFf]�G�k:��RV˔_�����v#I_sa���F���C�W��oqO5H�Y,v�1)�V���	�&�{��.z��z_������b{�/�A�t�pƘ���.��)eƳF¥���]2=;��j�r��t�[Oz�͈ �S�VX[��ݸDMZz+�'�e,9��7@,U�#]Lp��c��ם�Ֆ�m�ܒԻ����yQWa�Y�wW��a�2���Vf�
C�#�)"v�b�Gun[l˧%�[�P�HVy�
������V�B���7�����dł�Lap�b��Ŭl'DJ󹮳u��ڸ�gm���Ƴv_>@.��AM��+��v��bBʺd��vo��l�7��]��2nrz�����-�:m�wL}J�l�S�e3a�2�Q�̱:��̫JV�`)?�&�l3�Ƞ�sF��;),B��FI�͸�qGn��G8'�E�k{/��˵�Z᫱�.˜v؋;M�A�1�.e�P�W\�3�;`����6U�ss}��2]:X�;`1ux��ݹ�ܮź>����x�f��(��e��I��t���Wg2Hyv����x��QZ��C���B��o�������N�R�N'��r۷�/��;����'�٫��և�}�j+6Z��J� x@���1v��[��	�& c)���f��ӧ6oS�s*3[z`3�r��mJ΢Ө�`�������:h�V`���f���N��!zJ�Ct\��	\�Н��+*p�[��P�3fLբ�&
\���뗋p��L�A}t�f\5���x�%{{9(�L��o�녊O>���f�l
j@�-��43�9���ǀW���%�ţ���I �����b�PΛ�{%�����^:ۦ3S��;Πa8����n�)��*"{�,�tA���W9]>֫����7x0S�	d���;��ษM)>%�aK���s�e�(͹zx:P�N�Gh��Uv�-t��{�E2�����ܨ�Z� n����p�+=M
�A�z��Yw[7�l:���n�^��]���$�k��id���y�qr. �#�t�^���j�k�Vng$я�Q[��u�ۓdjxj�㷘�=6*
��:����%�,�˽%FAXd�F�h��.nMQe�)�a��v�����!��46/���#r۝66�+��@������Ƣ`�x�k��S"�ϣ��hm���x(�H��-T���[y}����^J�{�Ս�6���yB�K��t�MU�!�owA����rn���h��[��8�x�@+�zbPV�.}̀�m����x"�Ғ��G@im4Sk�Tao^m��ڑ;�rU��n8��|�6]SaЎf�j����mm�4�k�/�t�We�ݴV;J�Z�nX7���oV7/H�P�����}��.,uY����഍C%C�����8��Vi=��tVL��M����	�Q� ����r�޼���Esr�d���Ώ�v�ht��n_�lG���s"���w3	�)�%GNb��ZR�=�n����'���-�J��Rڂ���]	H�[�1d��3`�6��"衷���R|�8i7[��f�Z�=�Y��,�u�v�
��ވ�%ܲ@�*Z�����xQ;y��m��S��9̉ܫf�y���c��|V��Y*��+$Ɋs��#H\�y�_|���'��+ݠ�L wYTp�H�W"�H�&n�p�X���7��w]j��3�m�[�6��0��
F�o���eݕ
��&�h�Rλ�*9��n�X78��Y+`[[�jNK I�ٛ����e'��I8r�_v�3���acu�m*9Dӫ�t2�@E+�8�w]�V�ނ�Y8�p�`�� �:�%;�mws1vDkIk��U�]liaX�\��L��	̚�w���]mE\_5�tZ�o,u�R�2ȕ�ݓ�Xʶ������}��=��iڡ8�œ`E��;/5��+s��jtxb��`�����8�wuGY٧���-��!�*�VŨ�˔�(_3v@����h��%�(!|�M��v��j�霪��2+�F��,R��l*�G���p���Lx��4�6\/hwF�^B��=jm�4�b����Ⱦ����,�=�ܪ�f[����F����E:��|����!�VR���X�Zɫ���XhS�#�bv=HGK2��G��lCN�l[],7r����� Ol滓dOEL��1s�XA���b��s ��Y��8�VƖ���YOqE5�B��d�#]�V�Et �6>��5�Ev�3�+�V�tx����X��<2"
�1ũ���}fe?���uȪuo+�v]��Ʊx�uL���TJ#1�{�.Xl �<��gdO���N�@z�竔O糵��Î'�V�J���^M��/���r�C�6vC4�l]��}3����ܒn���k��ޓͣ/�]�x�9�3��I$�I$�I$�I$�I$�r7�:��$6�rX�*��t��j�}�֪�0�v�R�[]��|�����9+�)-��An�o8�{�zzʝEi�R�=Z%�i6��L@�����@)zh�x��S)�e3�d�X(Rq�g(�<���;�6�N���'�Yx=J�6]A��zC}g��YG��{��μ��M���6��`y��X=�e�<P�z�-_�;�!��X���`{z{^L��݊30njC7ZV6�ܿ�����ͫ�M>�i���o�X@4k���1m�DD@�7E7c}ؤl��!�&�F���?np���WF������>�J۟k���W 6��]˘����u����Fi�X)�r� �Oy���V�Ӌ��v����Yk�zuwky��6��[�[�7r�ȍٌ U��i��X��]�[��M�l��smT�H^}�8��Z\�	YW`��&���:���8Z׿%X��ٓd�=M��#T�m2��r3�E=�L�U�;k=ۦ@\T�p�K~ESmN���Y���٧�����c:fJ�b7{��vX�h��@���̔�z��཭#�؎X7�K=x'r�P��߲�_fj���
m�ٻ�;=�yͤ�GI2Y��nH��y��Ek�Z��  f*&�l�k+y%%��$�o�ѷ9��5ؤUc��Yy(+2�OE�ą<�b6{�l�����#��C!ݽ;��ܧD�Euu>]���@���]3�)�F'x�Ҽ�y�����[5�l�|���F�E�qfH{4|,җ�7Z��d�%��:o6S�N���+~�m��a[/��lU�3G+��Tg�γ�m�s�g�x!��&��_
���]���J���	g]��v����2��⺮��l^.Y�����\������2��kZZ܁mefJ�v��;�͝HY�Wo�XͱK:wn�ώ�{I���4�ƮZ��i����;.ҭ�)��E��^7�p�n�7 �Iy��\J����fzUݕ�4jV�f��J��Q��!�0q��d�\C˾��+_�Q&�C58�ޒ�;�ǡ�=2�2^�/��x��/w,*Y����ḽ[��c��kT)�����:[����4ǆ[�|�N��$�s��	�d/�mZ�,
�ǆ������gj���u*�?fm�C}D�g93���8����Ua3[���"_)����brl��gv��g� �����`]/�+�>�/"�c��c*��z3I�����e��)����T�m�ǭ��\$Ƒ��S�y���ַ�H�:��:Ū�&��ncX�$x��:с��C�F�R���1�L��Eu�4kN���Q���+4�,g*��
�ܣ�VeޗL@4��787}��1�����v��`�D��e殲��T��ѵo��~ڀ��@���Ui����%ͤ��5/�����87� �C������(oV�/��'p��/��n�]�/����(Ao	��ü�(�"�c8r�K�����!K�\��@gy�)�)!��%�;A���V$�J�j�u��p��3��ﯪ�e�K��D�j�����!�f�lmv�@�|XkID�u+��b��|3qnF٭�4�ʖ�U��fTZ�XdG��X��X��J� r8�rWܷ�b����G	1i�U�q��_fe��p�T4��e��0Q
�󰩗��l�)5K��q�q`��5��T���5գ;� ��w;{����f������lL[8V�Y�2�����e��t.�k�nJ�����<ps5|��N�-ͬ���9Ӏ'�)��`wb�[Y��(����n*�����u��B��H�w�]�:ڰ����/$�h`i�Q�m�o}�d�B�e��Jjn S�a֣�y&S��@��{�%�ju�v�AMh�YP����-ȯ�k�wF��.;L�֡ۂ�ma!c���z�+��$71uĜ*�t1�X�B� �]��U��Yo;;�#�܃fK�0��_Ej�
.���0tV�t��3���EY[(��!��Y�G��8�@h7�2���L�Mг�ͮ}��p��C�L멠N����eҒ`�\�'�+y Z��)���`}���%mݎ�TT) �X��ؠ�6�罼����Һ��j�"f	��hc��@u��Ki�EG�<Utxcgw:ӽ(\��[�1m^˸<;!��[Đ�>�eY�ntƠ��0���F@���tή�9v�j\=�V7.�n���b�Z�j��O'a�aS2�O�f�s%<:˵��XV����Ԡ]d#����b��n� Fs��Չ�s&[=�ZX75spK%��{:�C���qm���3r������O)�y�U����%k���K�2u����� ���vt�l�.��Tlwa�1�屨4��mܫW��(e*y�Ek��kV����rN�G犔�5��º�x�geo7���Ĉ���Л���N�>�!�7� =����B'J�v5��oM�b���\���m��*�n�k�U�n-iRW��Wq��^�{��*�Y�U�����v�޳'Z����f?����znǢ��#���{��m-X��w.Y��rޚ�5�F}"[�c���ӾWB�Ρ�U��j��-T��ykBP����s����l��n�0�!�8(�a�����.�j�7�����V�3���m^U�8�k��9��f,bԲ�Ŵ½֬�����\�c�X�$�ŷ�sz��5�,ҜXM@�d�s�]m�\(Q{m���u�:ro�X�վH�V%w׈AE��V��[��l3EB�'S�rr�lg���_L�g̨q"5��[��х�v�4 .������}��8�2��u�P+�^�͌X5fx^a��c��IR��ݾ�s�h&!ӊ�"�T��ld���M���m��t��ݲN�r�����vށb/]t;r�]��3�]����xf�a��im7�®;y6�-5&^K٠���� ��n�7�F��d�6��-ʖG	�������!�,�X{F����,z(ś�����!R$��\un漫�2\��tM�(�=�9/2�ї��2�b�l:����Z�uݻ��m#y�3�����ڼ׷.��Ra8��Ԥ� ��t
-�Rmع
�Y�����T���e�Ob�
�!�s���sw�@X�hs"�FӷV�l���V�Dwh-܊�䬺��)]W�m�J[��{��f��8���r9�c�G.�!7����Y�Ff8H��@S������U1��j��\�a�;�^4�YA�ϺQN�w�8��+��T�-�)����3����U�u^r�&�*3m�\UN��[I�KN�U�����t���>��y�2�e�c�LX����A��XY]��{��9�=��i�"\+Wu�K��������杚wvdL�)��[�w���`�2١@48�uF^���-eٴklC��F^u*PD�ڊa��P8&�|�������;H�PP��"9�ʽ�l�q�$�$�U���"�ª_f],��:� �����W��+E��ڐYVr�:�S���l>u��0PW����Z��7W�z��f�D���Y؜[�V3y����FK�r:�:��7���,O��.�rbk��R�H^_[�
q���*]�u5ѣ�b��vl�>��7�T�xF�� ��辘��9A_#q%\D�|>�/R��X:�}�f[#rcDbb>��Qڍn ,gg�����|�<�mN����wv�}���&�ug.d)�%q�xn��3��zQ���K�(5̧�:�u��:�`��g�;����^2b���OrV�0EҲ��:��Xe�i�OU�Lȹ�ʴe���[}]�k9���7Z��:H�:`��K���T"[Uݺ�xU����V�^Pi�)b?*�|s��`�5\�}"{@Sw�)4Dk ��|� �}O��YUb͡�Y��	��p*M����Rrq������*�8"j%vk~��͆�Rڶ�'�w�ҭ�q,�2ՙ�tՂ�o��k�������H�Z��F�򳝹���}Yt�u��	37!�Ԧ�%��G!-�Fl��>�����M4k(���Z�Lp�T���Y�ˮ.�r�gf����Eff���S��w�nvP.��o���n],H��B�ge-�'{�K��X��ӻj,j�5�6���vɏNMY�X������$�s�I�vE
��c4����Ym��wݻ�v
Vo(�a�}�,�.��Ld�/.��F=!��8�]��h+}\%��J킟+���'Z�����w���Yu��Q�y��B�3�`��R���o��[;](d �e��Nnwŭ�\�n�8��k/<xܗ����l�MO�9���W��q�)h��|�f��z2j�����!���h�	�[jR(��׊*7����<�`���ⷕ3[���Is�F���nK���IY[t��`���Ȉa-U�ey#�%V`���Ni�#+wwn!b��c�7hо�C5J�����f��8�ZV��(Ļ�G�c����%^;��5 E��U��ʗ�uh��Г���5ǝdȭټk�x�[���XP��^h{*#.��c�,��KTR��T���s�n=����G��� Q'-��%ۜg`��sr�f��z�(``��J���Αj���p;I)��ۙ�}(wk(3v�V�mwC�N>�����&����}7l����"���s1�Wj<�Uyq�i����BT2}-]�(v����<�E�Ku��sgw�j���!�V�4�ԏ)�����vrs��:����:�����
A�W�
���f�أ�Y�}O�ʀP��M�V����I 7P���e��X%�����+�HJj�<F�Wo\4{�åe:'3}���[�U��b7l$$,��/FU��j$
%Y��q�TUն��p�$��U�5_��{1��`p���zIAαXU�0!B^��W���Qc�5{�q[]
��7F�� ���"�._,(�ku�U�6�e��/����o6�_	��1�\�:� hD����N�� 7-i��H�[m�{���nu�v��˜�9+����z�W)���B���j�c�Wշ�ϝ!�a��mneff�e$\�b^4�$�|i�ZE%6�t\,Q���s{A
��8�\���rD�pR1��0��]���[���ꊊ���[-��o1�0_:h^^q	���Ky�s�p�Rޗw�7���`�ޚmY/O��]i.���g[��)F�Y�pP���m], ��kop��Ew�c)qчF�͡��Z�C8�599y�p��f�{��yN��z�u6�	6��5:]�:�2��ep�����5��3d��Nf�K;�W��ĺ�,�s��z�AO.-���/�n�u,�46։m��.=�L��޻�g��bi�V�D�h���n¶;�s	&ѷi&�ʶ�vmb��kZ��W�5֧f���W��ZJ�날�5z���"I]�Ɋ��e������r�궩�e��$�uNPv�%\���i�vһ}m;�{$��ow�~�t!}��m�΋k4�2q���c�ل�H�`��jq��\	b���|�[t3 aG�7Ok��a+�VGS�''��r��饳��{���oqz!W�+oK��C'e˕�P�*WK�)�͊��u���2�vnu�xhnIg-��/�b�xi2K1��qӻ�d���W�t��G�{�U�D��c�J�=�ebc~�z�8�
K��7��c�=����5�t���VE����R�������������_�&t�~��Rq�ɇ3f��V�#������S�����T�W(���ofcn��� fr��ȴhɷ*�=������,f�Q���B�1y�Eg����&;ql=g`B��/+�1���볐�y�KMd�l�j[Ǳ0g-a��o�h�(��f�n��:�.�V�P��n��$֩ї�9�HvJIڄ�j��W��泔^��koi>��_w�SQ�@
��äu�lCJ����5\�v�n���m����&K�܌�{ R��ZU�挆V�1A� ��Im�p����>K\Ud��2MC5k@�Dm��k��)�WR��-��y�"��=G0���۰`\���a�WX7�<����(�wj{��6M7I�b'�1c��9�����X�U%�����|p�6�������/�Dw�$��+�����\m��Κf����;���y���p�Fѵu�I5֦�[˲���XB�����= +������:�rRv�8�3im�9�����M�:3c㮻*�Mc�������ueӡDg�ֱfR�.Xҕ,��F�[J��12#[V��s(��e��r�Bb6�V+�Q�1T�fR�+ZUb3-�hZQr�J#YD���,U�+KDf[ݗ��Q��
�T*�ڢ�b,Vs�X���2�(�E1*�P�V[e��m�UV.Z"�1*	�V��k,��P�j��e�e����"�-�֠�[QT`�Lj��+�V�e�1"*�8�i
(�%�v���k+T�q�����-hS,�VLh��إJfc�q�ETQ-��%TUAU�UX�R%��r�Ī�T%KZ�1X�ܱȍLE��[��
(��U���TQ4�UL��Ǝ5��9lJ�2�m�U�r�U�Ք���%���QL0�2��C����]�ޑ�M*�k��V���ֻ;�v�>�H���/du�;T��M������r��)�
��f�N�g�W�/�� Sا��"����9}���!�/��M߆�:�	�;�\�X��?!�?���A��A!ҁ]ྡྷ;���z�~�e�ŜE��Ǹ�V��fU�XC�%���	&��>�#���*���T9��!�:a����{z/�p!��Uw�����C~�Bi��49{H_�*�
�vPҽ��󮫳��Ӟ�Oz�H������IA:J�)i�+U�n4�a�y���z��>�@�[]�`�?V#%�����{����;�QJ*����];$��_�+��a�X��B���;]�N��]J�B���d5;q�W��<���<x�>��E7�^�Po:o�I����q?���l����ž���{l���ڌ�!H������9�]��S_Q2Ѩp���H�ٕ,���c��6E~C�.�����l��?��!��9F��#���O´zQ9y��pw"��xU�껤��JMf�X��(ktC}�/]	h.C�B�]�����T`��e	ѢP��cu�Y��g��aut��f9ȱ��m��@º��E*L�Y�;(V�C�{�s���­�������v6}�3H��`{6���~p��^C*mr�����zM7��;��}yS��+����p�kx�<	~�j�7�3����*J�ٿ؀�vl`���Ze�A<o�$~<��]��_
��Lm4�R|�:�ei�Z�A�^(tb��w�۔���{x�b��(����r�!O}���v}6Φ}K/T��75�̳�-[��d{��Q#�������~�[]���%X/����ȍ�hW��ߓBB���q��/>����֗i�Am9℣����ё���q\c8,�
v*��g���ߑ����|�> p��}����?u�!?e�,�@�v�+��G%���DF��)(SuPy�/�.��j��V޹����6�C�D�S��y*z��z�>􆸍��p�aO=�p��)YE]�
��#x���*:ӛj��veG!�un�H� &q{�离�^�h��^q��[}s7=���^�����d�E\٘���Wk�T��퉸X{�1�[������a.�s�m�U��zhb5�E��
{���	���G6���
�v��0����ݙ�9�{،d&ۥa���B�uC�q��=d>����룹�ɰ���i�W�������I�������>)��К"|]�<��:
�syƧ��PP�S������|s��}h���Ж<�[K<k_*�;XK���_�u�W�Ѓ�+%1���r#U��)�C�=VqE7ϩ�����<����
�AE�y�۔;�����f����4��G�1��fO9Ԫ�OW��;��*H��o`�c�m��}�赙�#w��$���S]l�Q��^'��?��[d���	���mp~R�S8�ݿ{Q��I�U�Ͻ�V��5����F�5�4��P?`���C�^��"�T��Su���;�j�mb���w���V�3�}�)�>�'���\�w�e�E����'�o���u�n�e��y^w�d�i��e����f�ovisA|Z�R���ʖ��}�;|M�ÛsB�.,�yp$�f�u0���q��Rq��L���-�v'���|��+��1�'�M�-�H�!yt�~*�)t����ɲc�C�O��^	U��?<�{�f��<:���s�D�WzN����%�c�}���;���8|Ǭ�}F�}>վ�+����.��{17ʷ�8za���P[K��P�ʕ;^���S#���{2q�c�����k�1�x
�V#t���qX~���+풂7KƋ��GO�N5���*���ۼX�C_���Vu/����J�U�}�^�w�{Å���Mw��k_N��X��t�1�&�<}��Cp��9
Eۖvm��{/�;}�pz����c�n�9�?�b{<��/��?6d4�"�_o2����gm�ڻ�VP[x�鹤�%�:�X�>��x�wA8\Q�>=;�hǆ�A���+��R-�C���H��W�/���Z;B�p�d�r�~^�{��7y�o4���$�\�yy&ARX�@y^����Lܰ3{ۯ�0̙ȏq�hE���+�][�T/ 9]C�Gp�V^S��ֺ̨��gw�%�Eu�1�:�z����
�:�[�qB�q9[Ծ�ԪT*���ep����h��G�t~�^�甘�O>v���0線tyΧ�@���������v�dȴR�iy�QCX�6+�o1��o��a\�J���bWV;w���6ʗ�����՛Z�����;�L�B�~��O�o�(\>���k:WV����o��և����[���OV����F���N5��ښ>�Vv~�nV���9;53�{Ǿ?�m$:P+��;�B%���g��5�t�<&$:Լ{�z��$�%b�l�=�E	�����	��!A��9G��/=�:�TU#}�����~�a�4��up��C����p0�\��"}��5�Ƒ��)��۞��}�Y��7��5|Y�4�������3�w��]�PP�-ګ���κcZ.��6�U�=�`�?P��d�j���Pu��V���>
�@�}� �;k��j���=+83�6+8;2Zʮ���Sn����1∷-�P����Ȭ}������Әۃ[Nl�-xe���z�6l��闰��u:�r���1�lԜ��u��*�ۦ��|� ��Jϼk+դz�`Ck�T��r�@�e�3�V�"��\ ��7�
Nv'���<+�>�~���λ�s���ѲU�{�
c�˄$t{��C��k�sº���U:��)��ΓX�qo�W�_��+��Z
��i�3�"��]�tU�,����1��7
<Z^�t�^y������^*ޜ�/���ث�Om�/��cf���oġc���cݳ�L���ڲ�ї����x�S���w��.���P��-l�}��s�=�Շ�/'�F�������u DV5�]Gf�(�';<5tS4�Ɵx'��!�:���Qܥ^�A,���
�i�t+B�C������ܕ��W���=�{Y��'���8<&y�#�\��?q=��9V�m:{~����Oud��`H��a����0�y|Hp�?t-�W���Y���iʍ��|*-W1�Cm��r`
xu������L�A�Ke��J��J0�#��ֈI��׮���՝�n�˝s3��u6o$�����ɂ�\+a��,���������y�n�/����m���O:�_�e��Q�T��E�a��ޘg6{�㲙>|=��4�z���uB!������ʮ>*o�~�ǘ��&so�~�*�?$4���n�,�ڵ�N��ב�G�(7U��t�{��W��Mx���(�����#U�� ���M���>􆸍��XqC{�w�������M�`��y��g�p/��g��=!�V*gH�����"��q��������Aw쥀4=��}���ѡU��a���_]��ͮ	�rS��r��DN+��Ck>��O�_w?�gQH�j!�����l�1:#��vq�<��
��d���P�k�����B���g?�����U�=˃���륶���ߧ�)f��J����<2��Lz���W�q�,E=�פ�2��*����?A�	ӔgR��Nu���k�]����WC�\��.�m��*�:�]�;�|i7(�O{>�nYߒ.�/�N�1���R���R_e��Z�[� ,븎�	�v41$��$ ��r�X��aʶ }���`��M
t����K�mZ���5%4Iy7�´���
�MV�,�Cލ�clk���s櫕��o�9��NU�$z��=87O��[�����\+Z���GP�X+�:´߯p�������<��[���"�e���#������<0�����K[si���K�o٠�/��f�r@bl�.��X����<�YH���֫��f9���<(#�����B��Ԋe�����-ʴo����D��}�`q��p�����~�l�/�А�Zs���a��f����´�x`�WQ1�+���b�9}��4�����/��PK�!~�za~�C,r�u�$���MgJm�U?d
WҶPc��L4=t���|4��<͈Ь2�5o�UG��z�oo�.��`k9+�Ck�s�r��r����������w��>'�N�������T�lpZr��w� eb�`��gR���|&Ѯ||�5�$0l��ЭI�ӊ�KQ�"7We����*�:����[����w��6��}»��:�A���8�'sM�wM�j�}�E��#V������ԝ`�����]�sMY��Kf�!������}\e���A�+JC�W�������{���M�m�4S��7�睖τO��RŌ̥��2�z�J�V ǳ�8���P����K��-�gUnq~��Q:�]F�ߋF�z��e��Q�m.�����۞��XWB|�O;m�����J=~ZE}�
E�hv��es�;�߲����_�V��<iyVNq�<`�^�����r�v�e{��d����g�G�;F\�z{n��e'��y�Un� ᡼�C��iz��:.r~>��潧�'�(3W�:�V=�:Q!�}�rW��C��k�`�Y�n�� l��b�Lnr��m�����A�5~K��o��ü�A�+MY�:�|C�
��,WZ�/c�k�MpS�a�����iW�O�/��z�S��R�v�!8�+U�����-��x����g�}(�q�e�B�o�㠱��@��TGyD�ջ�;skJ������=�b������+X�L�~NS��{��x;yL�7j��[ؒ,>
�/���Zw�&�Y�F�g��]�GX�eL�����Ϗl� U�م�J�|�����币rj�oho���ޕ�C�p�e��BhO��{�Gi��
y]��Gvq�Qu�A{���F���7�Ҟ�n����OƘA�^�+�޴-���޸����]��|`�^����x�g��	��$'��3*i�sq<�+cv����T�-/B��VS��0D�a�2XA-P_�o��e<�;\�p/y�ٴ�g��u�����|�������;^�
��C�ر�>�ܵ��ܳ:��^�TvE=���=�cjNv/�pvW��ݶv[{��^U��F}�2:
5!p���}����X�޼ɕV����o7İ�՗�Chz�*�����y�u�J��m-�\'��9&]��s���I��)���׊�ӝ���6�U���W��x}��O�G2�ȈuN"�9��6�~c�e�X~}˼:��w5�[���/�?p}W��^�b~����p$�i�%X�$��}�ph�m�6v��V����l���u�T	��7n���v3���K7δ�d�	�yI[��\��p�)��ɽ�D_Q�ж�ECk�H���D���YE�����
N���
�3y�vqJN믣vl���*$m�&	�خ?ݣ�	���k?-K���u���)��d��o�4X�#���i�%���]��᥉!6V&h�}�M0��/!�7�+�-VUҺK �4%%���έoR��O7�
����yVV��.�˿��n-�t��d���B�na�A��$5��*�h�H�0�7�&���(�-V��ۼ�z�Y%�7�v�y�Z:#� I��2�T�U��\�Êɽ��!��9�t�
�c
r��o��W�*���ӗ�j80)O2�b��	�u��\o�y^�#�|��S}*��|���&���7��`	$F�\b�� t����n����eiue:�,�2�k�[5��L�.,2֢�c�;	Ye�#xlu>`���Ʀ�>�+����؉�3S}{��㩦�2� �YVӱ�V�S�� �2-��I�׸��S*��Kֹ\�u�AN�N�ה�?u�K� :�;�
7��4�+5N�����w�=8~��Q��]�Lȶ}o�m�p^��T�2��`0�:n��c/���w;�"2	e��mfS7�0L�!�n!]`��3E������rmX�=ʊsz^m3�Ӫ^���hqb�+�aS�e�4��sM��p��P{@���}����)m�ٰEF+��=��[��(�x;E�ϸ9��s�t�Keۆ�5�H�7xf@Fr��V�b9$������L�<Z�ML˙O��y�1�f�L+��:+���*��p_T&9,Q�#V�7��_[*�^A���i�S8t��<&I����Zh'p����'�cU�k�����5�	�uN�{�Z���1�ްT��5v7�T������&�N"Ƶ��i)���£��������z�'�7/+,F�����	�ë��Ui���7\!j`V���3��[�cF:Ώ�y��
���G��к���[���v��s;�q�\b���G�[�QM���ή�Z(QV�5��s�dLT�[.#�jvZ�$v��I�z�dWEk�q��s�<�6f��f���?=N��eވ6���1!9������������DDD�E����+��Ģ,Q1(���cEZ�n7E��f8�(ң2�EV9h���3*����D�QTFbUU���+�D�n[1�30��e"Ʋ��
�����TQE�ȥj�R�,����b�+
�\lkA�4Q��
�*�G2����Dr�*bUD�X�e�q�Ģ$2�`�(��X�Ƣ���J�Dc���1�R�Eb��ԔjQAEF%�B�*)��X�d���TF,A�cU�����,E-1��F �J�1cE��"VV�DPKj�E�DDKkU�D+�,QDQEQG,*��MR���
*�5kRЫ�Q�ƵP�\�Q��b����UUKB�����"�kX�6ʈ�u@��. ����3����Q�B�>��ݹܥ��%t뛧n""��{=�?C=�Bj�W�6�?�Uf�ͫ_�b+M����~����l�M��.����k�ٙ���˽�xai�-�ޔ�j�P��4��8*?�>�ׇ3���U��I�~㵖H��T�oe���a�g������|O�A�P��������5���Js��>�=�g����Ⱥ̆{��	�CA����p=�׵��=87��>~��^��`����q}�9[=��E{@x���g�����=��Z2�Jy����;�C�)Ƒ	{W�ř�3�	�����=����y���3Lo��"f_����Y�e���P�[�C�)��D�Ch��J��S��̵����~����Lz�3�Q��}Ըh����|r��'մu� {��"�b�2�Ny�a�C_y���Z;"�Ʌ=�X^�yzC�aL���KT�6�b��˪7^����/��C}��r�����x�w��*�˯C^guvӰq5��2X�j�[#^�eJƥ2o��ε�q��sJܜN�,R�W�~���_��s��8�Q���W@�S��p�@�GL��b���<)\��f�Y���;&t�rgM�>�p�v��LuM@<
�p΢���{�:�{�j�|���9@� �
�C��%¬V�b�uJ�Ɩ��T^��������n���=Z/|r�w�f��a�U��*�c�(�ǀs���ߍ+�f��A�N��k �R[V����#��m���h�C�p�x'a�6w2��:k�+�u�_O����ZVj��:�U�6�!�%�ʲ�8xka;�=�k�	.jϮ����}L�w'Ƽ.E���Z�R�]R(u�5��N�;J���J�o�����!��eP�M��y؋�����r49����Q����ʌ��3�A�ۯl�"5|+k�E�޿��9�n�M�@H�3q:�^���^c��<�,8�e���!ð��\!���t/��:�>,���m�n*G�GOso7p𛛻:(k�����(xp����kB_{P�E�E�yxd3nK���� �j����y�I��Wny�V@���{뷕u-���X}sd�ͤ%�h��|��~򆺽��k��;{BГ�����wZ/)oX�v]_lP��p�^w}4�sm�|�19�o�e����cN��}_9�0�����K-�G���4���?��}���0�|�0�W��e#[Y�8Ѯ͖���ႎzR��k��A�Yڼ����>��{Y�pz
(d"ݜ3Z!<yu n���|����E��-
Pa��#��b��4���׮�����>��I�T�>����`%U�p������O�1��`l�&����!��N���5z�4�~
Ґ���(�����R9w�p�onS�ɷ^���v��T�^�j�:��ՇS��N�c��9 �޵vJ���*��fk�:�?\=����'�@Q��7�E@�۱�N�Vs�D�]S�߳�iV�y+����9�6:��dk!#���:�?&O�˒��O�x>��x�Q���{�۞[�<��Of��+�[��m[+���%s�`���b2�G�O��g��߿gw�|~��i�V����1�a^R7Ԝ٢y���Y �^�]zo��.�v�a�Ӹ.��������
۹q��:bT�D;1�*�^3�s�)�4�yq���V����Mr��U�qko����R;�q_R�XUA[y����h�8�Q����(oNf�
�ﭧy˽���,�W�]H������m��y[;_0�A�&R�\�����x�x���5[��U�p}(�υh}ʠ8r��s����Y�3�R�zd���va�~^�i�a�h]�����=Z�|���-���f,_���^��^�=L|z=�.��B��P���FPƕo�Z)3Z$'m!�_)g���W��T��:����C��e��(MO�<}�"Giں��;`ծC ՞�9�́�o���iOn|�\"ǲ�ŗ�0�=���"o���z�F�H���ůq�q�9��7�䈐�y�����������=F��E۹�*̶0俑�eK7�dޠ��=�9�]":�L�C��cý�mf=>�b��=�#,�kٟd��&�J����u/�:����n՝�����"dM�d(Gg¸���<��7��G��d�Qކ�X����9tCYQ��).U����z����XyP�uz�nn㘵��T�%���W���,��148����hN�S�C.��wQr��^� �_{�;��n۴�7`Kf��
?�ﾣ�Ɓ�x�g�x��� &o�']��3���Ə�ѸO��v����u��[�+zy�}KY��Ǩc5�,X�kc�iʬ��Q�ͥ�x��{wW�$]���Eѡ�f�>�S�|:��U����͊������7Ϻ�f��,��^�=�0#��U��u
Ux���5譜�m�V�1�3�ݥ�ޮ��U��pm#¼u��?o��;A����'��wO��ƈMgy?�P��X��� 坺T6�%���¸nXN��;�9���M�<3��C��<+��vC�c�"����\�S�>l�Y�e��U��|���3��Y+�ؑOj!�w������瞻����7+����Աg��P�������V�_��K+��;"�3_'�䞡�Ư�M�_����I�A���ř3�T"�p��Q�L�7ҿ��ty�����xG���I�����%�b�禌�g���2��>4�L�����ϖ�|�Z�@��,䧓nv�T�h�$�ޱ;*<��0�AA"�ԧٓ���s�������l7{��E �Z��Pg�B���׎xp�<;B"#Q[c!��a�ܫ�؞U��S���_��L'�����0����6����6�շ��-����f23��v����F��� C�av�!�o�6R:�{;}3��n��Y�9{ɚ��z!�Cܤ6:/{������J�!Uf�:G�b�<�k�l��4T�U��8P�Yi��Z����/�_QH�j!�f���[o�g��(�}ア3���V����@GP��=XX�.��}{0A���~M��\��>7����a��,�#cΧ���*�n�����{�r�w�����F�|�k���Y��'NQh��;�q�\��W��0���R�/���s�7�eֿ�R��?����H{ҩ�l�� ޽gx@[�0�4u�<W�s
�|7�;��^$\L�~� ��"�ǣF�Қ��`߇��ZY��E��#�r�\�
�nQ�}Q݄4r�U8a�L�'h�>�:��(Kvz»邗��Ly���w�!SM��W���\���{��_ Cֵ\km��Rs]����P+M��Y�Z�UUW�7�ܧ��R��!���a�Ty��R�s���=WN������g}Iv�'E}ɗ��c��V���Fq�X�P�r��6E޶a���I�-����+�ܧ��Տ}F��|׼_A�_`���S-�<��l���O6�S[-����hϵ�^RW�_���}�4��kB_U����^zg����S+�l�����t2]�e�`׹||8miu���ǅW���ca�\i�kq��׺�"{鞿p�+��߱�s�P}k�]�P[K�XD:ҡ�p��/}z}�ֽ�Y�%�|�/���M���Ǽ�A�槀��b6)����>Qm���Ѻ�ӣ���3�҂�80�>0|G��+�m�gQ���>Uv�ej��|�r�y�������4./����)�+�P@����Wo�û:纻Ts� >�$V ΃�j�:�ua��?���]B���n��Kr,�<!X3��	z�67K:���;�o�@.�*�w��2�ҡ�Ne�kvR	�ښ��ާ���O=��)��܁�>+2��h�GXs��&����6 Y���ٹ�9l�4�)�mL�� }��m���䫧��{a�k��D)l��~.����y���U�:ͬ��$L����=�LpC8��ټ����M�u[��~\R6Jo�:�f^zW]�����n�z���cP~Y���Bt�W7℡c�U�K�}J��=�����M��P$�0Q^���q�ٸ�3�����!P�}�sf���y��,=�7Un��{�[��/3� Ǿ�3E�+���q��)�Wyq�6z[�_�ѩ�\�Z��7oƞ
~~#�{�[�;�
Щ�:ueau˰�V�pzL���ˮ�n��iao����0�j��ƕw��ա�!�?^����u��̚a��~�r��sN�L�����@�l{k�Jw�ff�/�4udy�k����{��Y�s����D�m���}"����������3�뗂��(�{��8w�|�!��*�����/��&K񧹃���pɧ ���T`L٘j�ʉQ�Bm�|��`���w-�t*��b9B��b���K��<��Ǌ�U����+:|xw���pb1�+��/*gi��c�]}��j�:�V2��]IJs_ϫﾪ��qrw��:(�5�HҫO�]�8�K������H_�U��wU��W��e��
%PR��1Z������o��u�\�#%��f���0f�y�*)��=��NZ��{�=|FYw�!��O/^�)ӻ���|�u��^U{��hz3�>N�(�_.����zJ__�ۡ�b��e��^W:�M��L?jz^<>z@?g���sySE����6!0W�v]s}=�{}��	�}���(mqW�(�k�شR��8��Z&��[���zm
^!�޶s�l!RLxU��=XGJ�-?W��C�X|^O�{�5���z=3E_�>D{Nq�)��g��_p�D}ϟz��w�{a��>z$9;����l����5�KJ����{#B�+l.���~��	�Iz:�z�_۫�zPҵ��ѸZ(m5��6b�Kf�ה�nK�a=�0�Q�(������єp;ytk;6��w!Qm��Ka�R���-i�5+ϳ}�#�W"��/�5�{�ݘ����ә֬L����/J�g*�s��8���s��4�ޫƧꪯ���Gw:?k�y������t��N����h1�/����r���
[]��q�����|��/��BJ�7"��C��`�ׅ:7�l~������^cp}3^�؁Y�3����W+d?DW����费v��UL��v����i.�H�����*�
�F�ʵO���Q�2�w�X��#��H_g��}cRVx�u�`�xg��YVg��k�mK��ۮ��CZL{\C<�������ψ�2���Sٻ�C��r��h�F}송��G�p�#_H��a�י�
I_���z����.�u��|���M2b���&��@�O̬�&����L+
�2s)�ed��~��*�����M08Ԇ���<f�Ϭ��Y���b�޿?����k�?_~��������|�����V,�߸u��
M�`Vk�L@_�T�h�`V��|}I��d�lǌ
�I��͠(�`T߼0^O���b�u��������|8���N!R��OIĨ���bx��6fAH>P5���$�dĬ⤬��"��T�)�hi �3ۜ����L*�GX��m��B	��������}�d�`I-��L�}���^����e�X$푔��N��\�È)n)�N��R
�7�r�q�+�7�9>2�W�EG�UɆ���2��7��+�WS�1��qѦM��v��y��eZYN�oTj����B2TΒW`����d�V��q�;%˷e�� ΅	goH
���.�e]����G�ɝu��+��gTyvT6iQ�H�ڥ;sF�;�s�����w�W�!��K�e���q�YXMv=��5��a+�`��u�!uw0K<��p�Z�Fr�w&�txo*��7��vI}��mD�Y�91�ܔ]2if�A��n�K:&&��)��j�
[Y�Ŭ�Hg#� K��4�%j��7�l<5�!J?��l�z�oz��f�U��T���g�#�VE�z��0�e�g]d�B#�wմy�IϹ2���Spmr��3���g1f��#V1�;,G����*�9��Y�m�B򲭪"�4;��VՉ�w�cX#��Z�\���8hYh�ڹzWO�U���`��y�N���Б�9S���=n�Q�}��m��t��K�K^�>cb�2?��Ha�:��O]�׮��UP�MI�Ҹ�پ��;��K"˝���& +m����1cC{�����ěG�Vg��1���
h�	}�*vp[%�"}y6��
s���e�"�����lm_vԮ��<3L5 �v'��U�Q0�v�5W6��]Yϓc��k���i�W�ɜޜł\�O۶;�8m:��/�p��oV�r�U�[��v�D��b��KT�93���m>�l��� ��Zy7�mD���V&�������sn���K������nlx��iu�NN�?m�;)1Xw�G��s��ͪԨ�=����ÖR�V����`'��5�5x8	9�v:�K1t�[��6�71PŶ��\��&4^9{Ň;{Ӧ�djGn��yR��η@�S��Hh�s�,�y��L�u�.���f�d-� ����7��K��vƖ�k��»�l����r�Z������O���IH�Ѭy�{f;X��T�p]��G�;')�s9��k�ЀZ�y�9*���n�YN�����րJP��V&꼾�ڕ�L�c"2v.=kh��O��O�<`��h��]�����]��e�uC"�w͚���[��02���{�|��r���V�o���CE������D�������h��#eU���2
������2�UjU�ZyK�s-D��̽��ƌd�EU�TQU��V1Q���X+4�q+���MR��LlU�AE1c*Ȫ��F,E����������2�1QTm�7-U�,b�����,iX�Z�Q-DDG)E��˂�U�Vky��lD�Y6�X�Ȣ��5�����J��Ŋ��A�
!h���X�Q��F0ETU1�q)mT�(UU����S)V(��Ī"
�UL��0cV�SV�
��3V�̔`�6PE�Y�V1E�F1Q�UF"#�1\(�F5[h��ܸ���j�"�VcQU
ѕ�R�Kc-�r�E���MffcL���QJ����
e�a[
�3*"&%R+7aUTDQ��Eam�����Ub�QQ�
�T�J�����QF1F+A�^�o��5�!��J���u��B+�r�D��˅��Ў՘�	֧	�E	k�+~�>�����$��<��{��u��@�Af?�?{���c~���
���0����!Sz��?�<La�+?2W�����)? o�'YR�7����qP�6Z
Ag�{�߻����߯;��k������u��
��GV0�w߰6�P�9˦��1E<?QI�� b���~d�s$�n�0�³l��wz ��J�v�R
xǹw�_��i�o���y���+m@�i��+�������é��>�I�f!�<�X)�J��}���
���3^Y1&�LE��T�l�t�Xc�>�}�{������o�}��}�8�6¡�J�`V|�O�iE�Gu��!��Ϩ�!Xj�!̤��@���i�I�6�'{�O�1�l;�,��&�E4��,1���ӏuv�������w�J�*J�VLE��T�6fI�F�Ϭ�&0�?]$��<��iE>f���OP+'S�N9�C����}d�c7;̓L����y��ۮk�us��y���������Iܢ2q� ����>T+<5dĂϙ��h
,�'���$g�jÌ1�_Xi ��n~�O����;��x|}�� /3\:��y}��������L��l+�+1�X�Y�O��%UH)��YZ�;a�R��>�i �7M0�6��͚�bi��q:�$Y*s|��w��������3���g��H/��CLެ��{�"�l*k�w2m ��h�բ�X|¦���`V|�Ն�^�k(��!�s?R������+�uB�䠺롟��*=��k�����Rx�O�zoH)�'\~B�R�7�&�wV������f+��E����RbAC=��g����ެ�AHgs'̕E<�N���9������ߵ�$���a��b|��P<�SL>a_�<L�7�1��W��XwtR
z�����e@��gi2�j�}�2�+�(b���UD}ԇ�Y����}�\�;O7��YF��v�����v����,�֍��j��F�.��5l�]z1B���]�ŻU���k�:��jÉ�a��o:ZƇ} y�UNWl�	6Dx���-����z� ���f�n5;~m��~� A������k�H6������a�����O�Ld�-QC�J���R:ɬ��P4���M�����a�/0�u%UH;�4ulk7�d��!Xc��m���;��7��oϵ�>�}� �wt�i�Z��Xq�����4�rɼ�g����~���Vo�LO-"�aS��g�H,4��ٮ�@�>a��^0+/�oΛ�����;��o4vN (��}�!���P7�9H=�+�a�?!Y���I�?s"�S4�m��H9tyd�m�{a�x{I�J�++N������j�љ�{�Ͼ�����~OIR
{�����La߱�T�ɝ�M3*��0��8�@��J�2u�Xi�0�
����Ag���y̓���SN��M�~_E�U�<�~^?��|w�Pb����V��
A{i�|� (���	��:�<>�M$�i��,+
�S�RW�u�y�1<I]�0�vm ���y�h�a�
�����~�^y�{�=���>�ܓ��Ag��(i8���k�16�X5��wHT?<gɤ���|����s��
m����s&��6e�z�a��5f$��f�>��=v<��F~+�~�������B������Aa�Xg�P+��4�_����b���}d�x�Rue ������Ri
�/�YĘ�
�xW��>�� �5�~���?G��y�������&0��'w@�%g�癄��&�f'IR����d������Aa�l1��TOs>d��~@���1>dӞ��O�w��|=-��~�͝�{�}P}D!�~,TT��Xh9M5�ܢ�]e�����T���2Î�H,Cw�u@QM�@���0���1 �Þ�����|=��J��V;���]����Le��Cԕ�����+�G_a
����OuH,�f�M'�*�J�OP+��B����8�H(o�&3L=LdI'��5�\�JV%���}\Y�;'f�L��w+�Ց�R�t���1�Z���Hu��i��ګ߶=&z���[�AS�IXjcGy�`��oT��s�#$渁�.��S2��>�f)��qQ2�^��L�k�\�{%�߾��ﾨ�ߜ׿s~k�4�S�����������m�:�a�<3�$�
�r��ٓi�a��a}�bAf���<��X~޲H/:�ϙ*A|�r����9o~�[ߑ�<�8�3�|H���Wߏ�i��~�N��$q'�?{a�4�S���d:��`�o�ɮ�?&0�h~�f�
J��U&$�bx�Jɩ�bA�βa$��㜹�|��~����$Oi�>����qbI�'����~g�x�=g�,8��CY�$�?�ąCS�VϷߞ~������<��+6�$:fa8�XboTH:��d4ì*�S�J�:ɞ{�1RWodR:ϐֻ�+��s�m�2w)��&'�}�������1l�i�n�N�w3���W�T���\H<�:�
�S
y�ea�1v�
i���M!ԕ!���+u8����Vo��}a���L�QN�����o9����{�s�x�ߝ��r�g}�0�At�f�����G)�`T������A���I��r�G��i �k�i:�H)�œ��,4yI�����=����}�N��g'���Y�IR;y��b|�J�g��i ��L6w�xì*Awl�d���&'�ON!��$�ɯ;��!Xi�w�'����9��8�^��^��t�vɴ�N��J�FN��t�m!�S^��CI����i�gP�N2��1�y� �Y��Xi�V�+���鴂��+���<��q��~k�v�� m ������B����f�;��n3�J�d����T3�:H9d��d�3���q �L4������5�i�+#����������wﳒ�d�Y�x�����׹&��k!��(��~�0��
�Cl1 �O��&��%I���S>��!��S���6��
D�`����{�#��F��k��h�Ss�*�52�F����V�]��������in@�Ue��weMD�OVƯԐf�jKhk�g�Rm�jWEG���6��:˹ne�ֈ�S��{2e��>������inN�=����u�]����8������O�0X)P/�S~���1 �hް�8�*��fI�T�)+7?Y1 �gY��a�
��i��d���V�����������9&�N2c����M��h��~R��x{t�M�$�����̢��Rb~@�&�ܚH>���
�S��g�1���b)�{��e���u�K��I5���>��=��C�6����Ɉ|��OY��6���C��Mv�����&���oW�3l��O5C�%N����R
z�SF�t�}��tw|�����y��~�}�"��<Ld�� �q<�E �o!�6�RV}��,��4�3��
J�tw���@Qf̢���I�P�a~�Ɏ0�¤w�^xs���{�޽�^r�m��Ӕ1��o��Hv�����4ÙM�C�4�Y���;IԨ�n�%OY:���� �@��{�?Xi ��X�3�9�����s��ߔ��4�>���̘ʜE%zj�ă�7�I�aRl�$z��S���� i ����o)
���{�o̟�w��u���k(����)�aޛ�����繽~��{��tYă�����R��:Ρ����3����A@�隰�a�
�n��8��Nvɤ=O~��ǈ��y��d�kW��>�������|���y��0��d�P���&��J��yUT��@�k ~jA���L8ϓoV�Y������a�bIY�&r�X���ɺH):���w��M��kZ�u�}���k�g��b���p6�i����s���P�y��aX�ư+8�QH��`T�<Ri!��:��B��/u�z�H)���N�E�����{澾w�k�o���x��~q��ꘐ|�u3z�{���9�&��IR{��Y?2��Cy�*AH6��Y4��{I��3YA@QN2d���q ]}Wu��e.]���[4Z����ߐ8�&Mx�,�tW;[Nǹ�[,庤���L��As�k���\�ͫ��T��9>n����Y׺�+��5b�PVآ�������.�_S�B%M*�Y�WV�����>������l�=��������'*��6�ɿ�c+%z�̧֐S�
%a�bA�������:�T'��I���3��1����,4�Ra�Շ�1��^g�����9����9���$>I^��>d�57�N�P1��+:ɬ�@���aY�N�>@���:ϙ��>`�f08ԇy�D+��o�d�H,�yy�/w�5���s�7�����=@Q@�鉦f!�J���X�_��$��`Vk�L@]�\a�;�>{`c0����Ri�aY0��x��Ě>�6���S�k}��������{�y�?{�?f΁��[<�̤+'yc�O�T��2~I�Ğ�E��Sl�q����)�����l1 �ɉY�IY�
�'YS����H,o�ߟ}��<�߽�������VxɌ4¿�X�Y�y�h
)�5�p]� T��J��9�?MY���̞&0�Ն3�%xɳ��B�S��2N���o�����Rs��������=���{���
Af��z�@QH/|�g�6�P���:��a�s�`m �Xk�͵<d����Lt�ީ1��7��<7f�~aY�O;� ��J�������}������y�:Oʩ8Ϙc�vyL�HVgɞ4��Y�Xq4���}���3�}���%b���)��6r��ydě�1aS��y����]f����}���H,>a~�O� ���x��`Vz��������=@��7�=�+ye'�*�Sğ8�iQ���'̘�;h�R���'�kO���;�o�?w;�|�E=a�Xc�W4���J�jɈ�q�=O-&$O7fv�2cP���AH)�_Y4���3~���z�Y6��N9�A���}Dh��)�1o0Q޹��?7��y�>g̕�:{c�)=IQ?2��X݇
��VLH,�5��mE���O��H.��3Va�x��
g�ǉ�L@]w�~׽�z�j�~��~z�%�c� �H���B4a��;�,�����ټ6�Zڽ�P3�3D�fG�Ù�a����	��|�L�(��7��:Cy(�r�&t���t��P�31�z����[�������������b$�1?��`g�L��-��=aY�~>�� ��M}�*J��S�FY�;a�R��>�i ��4����7�&&�q��w��|��u���^k�ߵ��׺�x�r�S���'��]�w!�6�5d�<>��a�5��M�9h�V0���0+>La�
/Y*)���w��7]q�c<W�ߵv���ǯ.�
��s��A�"r��a�A}gi ���T9�]7ڻ���f�8�/�{��g���7By�hy2=�ۑf��@�m�t�W������j������(J2��ުR��5<�?�9�ayuwMsw.��h@���@�iZ�*�l秓;����]��z{#��_p{Y�����S����:����5q|UJ �R�����g�u��=�U�Px/���=����"�g�"��۫w�˭��*��gP=�B���q|G��2�*�P��CH��rBU㺃7=�~�����>��Ö��V/��<01/�ӡ�[H�a���ckX���exx�{*m�ڦx�u8O\jd��4kIy��ѷ����vV6�,����n�/)��n�..7}�
�ۚ���;%��뒎7��!��K �p�>���^5�.�5��W�}�U��sr->y����+]
���X�'�j��\h]�V���<��ZG�y�Js��}���a|n���+ꅏe��摚w�E2�M��)\1�~��4L�����s�����'��aue(�~�g��ꄉ6�1�7$��f��_(���U`Y=҂���D�X�ZX>D�_�F��x�*uvb�z����T��J[�̈Ζ���5����#��=��h����ͺ�}�YoT�[��0�_Z�q������98e���� �?p��w���&�-��|��p~Q�-"a�?d.��e�$#~����	'��$�ٽ�q�k������	Ƒ	y��/�F�����S�ڨEbq����f����R{�G�Wih}��yxWxFha��}_$�m��~�3�H^P�D����I	����ۄq>�{P(;~]x�<ߩ�V��tged����y�4�4A��+��Dǵ�<s&1�����������uCYg�%��^�LC�c�����σ��$�+�]���?]襨��4�p��#Nՠ��s?+��着;��h�[�����t���{����U�=�E�.��Wɞ��i����FVz�&+P���+̭��!����C�~^��>}�$�ע{���gM�D�U�7��֟�<>i8�{����MCGˎ��������N��Й�k��*�}B�~2�A�qWaba�lz)Og�ԧ��n�S�Vq���M���7��OP��è:�[��<p�����u�,��Yn��LA�Gq�H�TCh�1����x�z�/nt�G�_z��4�Y���1?����^6�zz����aL��W�v:��/��� j�>up����@/�+_�Ѹ_ȡ��z���:�,ɞ���!�`�pxV�Ɔ�����s#���;�s���ӗ��7�
=�Ԉ�վ�dm�����~~�Y���+���o���%�F�`��z�����;�&�VS��R�b*����: �ma���T!܂�xFN�{��̎��&Q�|A�n�<��N'Z�v�S��qԲ��NZu�e��9ا,i[�d�'C�諭���ww���d��R�fє ����ک��x+˗#�o�t
ǝ�%EN�t�}'.�0e�������4}Rt���D|��C<��#�Yy;{n�:����?g��xQ��Gq�X�lxpU�b�5o	Y��/k�K���("3�'(Pn�Xq�~��8.��;�;���W��D������~��2��x�#|�p��B-��0FhM���or���x��.n���!�^�~�*�G��֐<�Umi�3����{�y_InYh_�X_��B��C�ɑB����1�ޱ����Y�}�S|=�ϸ^Q#՞D7[J�����D?��N�"Ǐ��'������y��&m���Lh��bh��0��|�e���Y�Ш���eK�8m�����΅q	�O�y��~���6��O0v�t��e���yG$�kc��f��f�n���袬V���c1J�����82�u���H�e�;�+��e�bm�<��@H���OnbAj!��g3$!�n�mC��brۤ|m�~���fN}R�
���a��_��ӯ�w*eq��s����ެb��~���:%DOB�8|1��W,�p/��a�j�,T����9{��yy��e�Svh"����VPTy���/�����T:�CV�����Ueef����4`�]�P/���PN��k���|�����]�R������#��0�j��Y6K�O�ǁc��)e
�<�y��[��n��ix�2o�A���4�w�FUo�0�x�EA�޺v���d�[�`r���cU/�+�|�4�u�����}.#������~��;{s��,�5zmǎ؂���{>g�˽�o�G}+�}��=_<Rˡ)��@-�%�?{�P�Ԉ�;�e4����P�e��U(:jx���O+J{�vo,�}X�ؔ+��>�̭h)�a��l{��9>��W��H��^��k����ݡr;|���n������T�S����Xw)\��{�ra���*T�QET�(1�_�v��v�:�r��Ɖ�N�*�bs�±��Ye�E�;�5*r��J��7��t�`���f�י�7Ew�dp�U���ˤ{�K5�0m�H;�Ack�=:�ک�b0�Y�l8��w+:ګ�;W"8���6a��Ye�5��^�0�.n�U��o*��]���mWD+\��K�*���kJ6	�#$��ev�Y� n:G�}õZ�"�C:[�E�X��hKۭ��P�^p;b
j�U;�`f�Q*d|Z9�GYE�����|{jk4ZSf��Q�)�͎��r����pM��7���wc����z4�$z,j+L���Z��e��dD�v��]r��_d��M���a٭.���vһ�Xh��ۼ:.J�n&��`�ʈ��Z��ǋtV�Y�݄�ΰ}d�a�h�&�n[\1��Y�K4ʫ�(n��@�|�U�-Pp�h���}����e(,��e�L�&!��/'p��,7Ge�|���9M�}�Ӹe�L_7յ&�5��ZO�e(^��Bm"3"�����I\o��oɟe���������|�F�S�֋ɓ$,�04�&�#g.�}Y���d�� �
t	F��%�Lٓ�
c���y�s�G�B%�9�ū�4���Ǫt��Prܝ�;]��M7���y�-�	d���B�y��Kx����]K�W�0l��Ĺ�\�[I�D�qF	��.n.eu+��N �{:G���՞�Gdpm�6��Wyw�T�:��aZّ���{��l4���N
�h������+B���@ł��:��hG����+j9$���<�7^�X�;�M]sC$��/��Y5��ͼ�"0�s�Y�(%���%�P��b^�eJ3F�|>Q�d�u
�0���4ժ
]ඝ�H�ɺ89�>���t���
/�E�����l���NW�������2l�/9]���Y���_q�Vh�-U��[�Zӗ�!q�f�vPQ��X�Q���>�^�R䳑��DT��&�������]
`6�*��>���"�;�ܹ��2-�8�iǶ�b{�����洓icٲѨͮ/sH~D�}V ]Z9�����UX�1TV,Qi��AbV;�������E�j�E��b��* ���TAQDkUD9K"+Ơ�V,T�(������J��V"��"���4�5���[*(��b�D�
�1b""��(�"�Ab���H���*��5+1,Ab�X�E*���`�֠*�+j3MTդTe�"��cb��US)EE[J(����6�A��X���+�2���r�*��EP\�
#R[Xʖ("�"!m�.�Q�AV(+��l"j�"����ŋX��d*1#�Bڢ�+_o�ߘ];`�m���&o@�G����*AD^����Sfd��v�ʼ,���nG�|> ���QM�c��?o�о)�?p�~έ���xh\_*P�!�3s',>����/+��  L<<)��^ |k܈�ZD<�=����X�a�]}<�C3��,�}L�G��)_��/�_�ɵ!�B[����o�E�����rH���xF���g�eu�=��,x`b_k���ƒ;�J��48��j)�o=���gԏ���wʙ;BC^����+���V��VN�O�;$���%�?w�K�*��s�~]B
�g䂻�R�{Lg���a�~Ъ�%�9�v=�B�}�a�Y�+<y©3�o�uXw�ߞǩ�vRO%��� ��`Y+�(/Jz4JU�������C��1�}�J{C�{���]�#+MY�m]w���f�-O'|k�!��B�!��VM>�J7��/�7����W�3�_�M//���\SLf����݋��l��U�k=/_�ێR��t��Юe��i��,�����66�<&x8]	[S��ۛ������ط�)�5�#S���;���uHZ�I]�sx�C;i���%5�؆���7Z_���| 9Wo�s0y~��;�tC�d2�`�حk;Oh�{º	t/n�x��	�2n�{�x�2� �}�{ô�!/r�?OHxi�g��Oa��1]]���z�0W��o��,�1�WvG���~S��xFo��nծ�e�E���3���H�d���%I	����ۄq>�Gj}YS�zg{Y]+�x)}�����A-L{�=���Zϣ���x]���U2������Q�+�Ӷ�*�Њ}���=
�`Aw)���T8'����5Vz�M��ۻʀ������9���e���.C>odNen8T���"�u���]&
�E�����/x�(mqWaba��N�/�Z�艺��ǵ��7�ѡ�!��w����g=!RN�����U����:�[���خ_�5d�}�t�82V �9�W�6)?*Z=r��.읊]7�2�=P��FX℗뾃��1����K���.�8���cP�7�p&#��5*nt�ʷ�KY-�N���}�r7l�np۟쑷�������U����d쫽�{V���+��z���]��ٍ~�����=�L,H�9���z�<����|tb{I@�V��G���WA��[�f�Iy�z�:#�P�ڀ�����\�=��������wOMx$]�����a���}Z���=�1w��wH}:��~�F�C�#}l޲��������z��W�)l�g��;>dF)!.Z�{Y
����#AV]�n�=yUK���x;,_'�u��TS;�_��_`�F�[�hr�����><���WFC<x�9��|i���T3�ӷ�Yyε�ڭ�˟U��|~��uQƐ4�σ� pC�M����7�t9=�}�q�s�9>ɑn�O
��B_�c�C�����f�U�.��eG*���M`��[��{����y���_o6Jm��ǏJJ�*����e�3ҫ����UO-��O�l�1�|׶ʁ3m�"��2)'3��"�`���.$�T4gk��/Vu��%Lb�'��B'K�K2�A�$��/r�ұ�َ��ˉ"��7F1P�0������t���C� �O�_}�}���q?/�w0~n�oԾ8U�1R�s���\i�({�!��'y�n�3�;�Ӈ�gXG>W��:D/j!� H|+*��.��'��5Wk�l�/wk��h��k��LW��n�ܾ+���]��VE�Z�g���S��R��t��y�2�Q���:���YT��T��Z
�t7Pg�WEi"ў4����^��Mx�Z�{R��*�+�^Wo����eo/�����֛Î�)[W�z�EĊ"��7Hc�¨tf�u�CӁ���]��[9G-OK5}u���K���Dϰ����h"�������Tk�|��y���=�n={�����A}K�T~�X��P"�S��3�jX���g��g;��~x߸��t
��18��Om0��Uj��ᣤ��#�O�ד33gc���Ea�~_al���q�T��^.���4��'��}��� %�NA��s�Щ���4�(��:L�U�kIŶ��o�!���I�*5��ޙ���;��`��mp�\D�cm�K|�ȞVVV�����s�9ac2�p������>Z���HC��;P�S�[�{K��_���矑�P5ھ~���RVp_�w�t̿Qp%�g|�~�c���6(�)_m7Bz�)���e�w�jv��/��c��~�Y@��.�����'C(J��s�S]�]�CL�E�p~���+�{�z|��,cJ����oZR��=L��I�u���$�RG�m`�>�]�J�R���|6�p�x���O/��MNh�>��"��xK*���[��> }�$V��"x�SPZGM���Y����y��wj�Y�a�`�@8~l�v��=���_����^lj��\�)������8<0_j���[H���E�����\yb����9瑿�}ʮ�[B���_v�=ƞL6���om�q��u#�;_�\����υ�!�(�:���X�Yf�+��.��b��(.7v���|]s�6W;%K)�ہ4!��b�v�.<6"���W4�|xe�`@�]�1N�{OJ�H��$\�t;\+��v�L�
r" ���4D��F��*����#'�����򪬛Q�i/~��=a��zj�P�^�j~k�����I���w��J��'[h�
j�f��g̍���9A}�OF��k��|���^���9�5Q�c��ڒR�Y� }�+
�����x:����/�����A��zFd��w� ��kټk�C�|�����U�i���N5���X�_�SG�=���+S���N�^N�����Hn�S¼7��,��2�E�����!!!���]����麸����>����i���OOHxi�v�_,�m̽���1WdS��Sx?Wk�j��\�>�\�4��W��^�b���o�#��r^d��myz�/�#x�����PT�3�w��Iz;P=�d�'����8����1�����Ai��_�=C��;����wG�x���r�72���ay58Sҷ����,1��O�'�o`A�!~G���f{u����1��f^�+�7'pN5��O��/�"��מ�ۛ)��䰝"o:��h����.mmo?�	ΐ�S��g\7�=���х��jgi ��Nz���p����K���:��1s_��꯾��)��}G�i}x��7��O����Z@#Z�6j�Í݋Ϊ��<���"3�WR���+4���?�^�YCh;���;Eq���x�8HEm�R:��c�F�|��0x~�M�$#$ǅY�c�.9��6����f$*�����:*�S�t�82Ubң�<j#b��۽���w�_�x��f���<G���~X�������>���,JV��m�I3���^e{} ���27>"qA�����o�	��R�^��=+W�-���oN?f��X�f"����V��C�a�}�,���T����u�"��L�X�uƅ	B��<6��kU?<�T_m�h�r��̌CI1%�Y��z�
�dw�`����x8t#�V��Y�m��U�%�U/eͭ������^�tW�4�����Wq��).�Ѥ�/�� �(�AfDZ�߶���c�o����y�R�m���O���C+VxM̱�]��b�*bS��4�ɘ���f3KgPm��"�]��j��z%���7����̩���`j~�����In>�b�����T��҈�B�
:~���ƓaY�޲��_yPyx-�x��Oj�
�p�<+�8�>)(SuPz�C<������^���m�7��  a�ǂ�K��(b9dx�5���l���F�`���arc�{�y��*�ZC|��g��2���w�� ;%o.T������'隽�F��*�/�Ұ�W����dW�W�6��0:�1۫V��{yƀ��>r�z�]�����.υ�r��|��F���s<�-��k�zGz
�B�������vS!Yx5j�"�&`o��f{��t���_c�=C�8��9
��L��y��?p�S<Nz7���c׍�Ŝ�R����9�Uo�^X�8>\�u��+W��A����y*N��
�H��UHy�*�ݵ^X4=8��^�_�2���A^�r�ۭ�����E��^���4����<S���Y{�m�`0���̋�}l��Ut�[��ŉ��>W�SoՕ��|vwn�/z}-����N�s��v������2�hR��r:"{),�1�]?}_UW�3�$��c_3^œ��5��o�W��D����Z�3�g1)'!y�~B�a�7ڍ�x��@����ǫ�CU+�G��62�����a�S�͘�0�#d]�fd�'��!�r���C��`N���Q�m�>kk�EĊ���z��yO���y9�-�Z8�{rwC�
C�KXx��Jg��Fj�t}�|��U�`ӯs�qÏz]�{�����g�/��/�Y���}��l1�k��m	��4�[���d���Z�hzV�������̾#j)�������˽A�Ｒ'j6^U���S�T�Kř��k+
��$x��TY�q��q1ʰ�����ξje}^���������X_S����k=h��]=5��ۈ�{�;+a�p���<;��a���H��C��<y�/�
s�X���#֥D+ٹzΥDbX���t�/zf��V�m�B]��uj.ɜR��-EjZcv�yYZv��id��M�S�{t!8_a�p]{�����A��(����c�ս�6h��T�L韕_U|�{����W5��1������y��fC��R��3N�}��\�.I��5��Su���Ī�βb��Yc��0_j���B���Ӵ&d~Ǿ�6�VpBP?o�TK�����d��� ��W�^u�0�I{>d��C����c/��%��+���0�W��+��DǪ��kʎ �Bas��糧�ï�c����.��Y�a�U��g�@j���i7�}�{:?%����&�k�%�;���-���X��x�#��3p���(�yS�L����~8e�������{���+L��a��p?y3_f��2����k��q�g���<*�D���_mc�PqL55t�-͍�m�z����5�
��ƽga���,�m��̢:-��IO���.�0W�k%н~�M	��a�#��!w�����.�����5m+D�K�|	�L�;�J��WS D�r��=��0o]�g�dqC|�t�SA�w�����ٓ�W�=�DH޵�Yu
�?=U��(�n�]k;�kP��n�#Vax``,Z�r�P�3���j��!�(�r�Ept6=��}k�6fɒ%@��P�����ɀ�rr2�KC��E^�B���5+	�6��v,(ooM�mM3��_+E�8���7V��;�6�5����c-�����'Wvu�.�A/�GO �۵�v��&%ީdgSŰd�[`��Y4vڗ��zH��y�zf;X����֡�U�X�#���vc�!E_v�2����Ў�mڭ��>vgk��9)p�&�Ѡ�$wC�����E��*kk��ub7�������Ft_)(�Y���[È��
L�MkW���;�T���G(vvwcה��2��lqT�Mv����匥w6��a�:�qw`��D���--:+L�yk�v��]5F��xٚ���^��7�ڣlį��of`o
"�V���sU/4���-䫺�hP�j�H����b��~��jd6%Cy��q��9(�e5�A;+�KWU:�wH�9Ai�n4����e�&�d����^v4����_|�Z�m�J�;��;L]S��>��*� )A��t��[e*�ʚt�d�u�\���]�+V�z�(
<wY\�n�к�[��H���!0��g��>��Wy�3,;�/�ԲB������iHd9�S"�6��
;�	�$��)�MV�X�	Rt�t�4J��]�Yrm����*q�ÌK����|.=]Af�S�[f��J{�xGP3�aLL��*�����>�7��o�ӊ��t-9�Gr�v ����#s�E�Ȯ�&2��Ә��ɲ��_��Z�Yc��*�s�a�/����h
M�v�lzLd�tOj��P��8��|\��%�Q��EwçJ�.DKӁ�٩��f�\����!�o��BPl�:��1�87�r���ȅ4eŨ�o�%�J�f�)n�89>ZĲ��I���wט:9Ο��2�)S̮j�ڰڂ�)��tz#k9uHd|��o��iJ[1������m�$�e��	��tii5i����ݦ�VLY�+�5�:���-��m���݋	6�R��B�֏*���s�I����߶?O���Q]%���ڭPQQD/�U����b�(�U�bV~h�,T����EQQX�
娈
�DTE(��CIU�UR"1S-�b�DR("**�R"((��%�VT
DX�4��j��0SIQH�R�AE��A�ª"�
�YEH���G����TDcX�X�f�*#VQTAA��")�RQAF�-aU(��� ���#U�P��EX*�R��,E��UGM�"�#��UX*������ߜ��I�y�sd\3���� j�n)�a�]�Vh&P�A�F8'lײ��Ђ�O������׿t���>^ނ��{�	��<^�'�W���������tOt����{�2��Y|�!�uPz�J�<-�{����/Cw_,;/�}��V���_+>������^�`��b��|'�3}ouo{6���t���C��O/^� �����z� ����d;�����&n_}��V¬w�@��Ny�UZ~/�0z�wwԦP�����Z��#�B�����V��^�����_J�{�U�4z��A�r�r^��/f�O>��y��+�'�q�J��-��g�L�ǼiU$ǂ����n���m¯�=>�l��i�����{n��&3F��,�DX�q�^G�3<�rU��
�]u�TG��߂��������1:�J�|���{&̘75�)3=��Y�|����w�ت��|&��K}�@_���O*�zr�!=\���0���*#ct$`��o�}g��ء��yi���)��7nFo&����Y�Z��Fw:������-�/���t�\e]n�*��\���O���s"�ge���睊[����ܕ'ߴh�-6�ԕ�T�`zk��8�.��	
�Y�x�M����oo�9ƽ���4�!��K��G *V�����_v���w�RN=��a�yɷ\���v��}��-��	�,��xw�>y������.�2
1�\�l\o�s�p���F��e���Ѭ��{M�I��6�0CK�!����fǩ��萙�+��n�#a��B���3�?/|m�ж)��ܝ���\�]o��7��Dd4�)��=n!�B�~��jf�!���+\v8�
?4�S��S����ha��5�o�1���}�p�����yݲ�ћ��!J��$'��?V��"����ށl�4<�W:����J��Xb"�S{K��g�R�*χ��O�P��Q���Z�y�s.{����.�D+M��Ԡ,�G��ѱtM���p��q�ݵV�8e�@L���pK���)���+�z��*&��Lk�R��.���
�@��i����kV���ʋ��nk�g��{����ks��m~���}��-+h%m�(�����?�U}�^���ڒ"��-��W
��Ք�xe���U��*�)���<+W� ��X]G1�T��$�/l��Y�y��Lx0u h�mk�b�@ɷ��MiS|���~Sw^w��$ϑ�v5a���N5R��q����ܩ�״���sڿ��uu�F�Δ�!��V>��ܫ�[�j�����P	
�/�c�n���<�l�Ey�R"y߈^�sq���)����*���e,� �S��Yc�}��k�X?n�xi��XD4*W�OC���,�z��M��V���V&ȡ"�[0�%�>��9}��P!�רK���?>us��_O�)_WȦd!�p�E}n8��*at�t!CEbֵ3�s�w�w��hkx:����>���z~�\����fئ~>���r$H�����!�T��<>t:·^7��Z�l2�����j�������V�sj�� ���0��"�5�;���3�O��#^x�Մ��p�g,�n�/�p������O��w��R�A�sy��PZ���Ǭt�O7�X��a24�hӃW)�g�}���{�1]��Ֆ]	N!�8/��}eG�S�U��z2���M˕T�XngQ~ȥ�����MOa����5�P�#4��[�(<X�a�%�z�P~󥇨m��^)Y���^�-��f�q	�c'2>uH�|`�
���Ҽ�!����Hg��'À��/ǲ5:��>��:i���꾕���C���8~_6�7�
S(=~9�z71�xA��45�M�*��k�^b��}e�������{�G��!U�}U�ȼ!#��P?l(s����RP�K��~߳s��-v��i�ٓR�T�W��Z���l/���<3���VW��s����f�2?GsW�$_-;��xoټ���z�(V*�0�,ׄ�=%l�6ۓ��v�;����\40�5o������lt=�X��z�CP�B'���>�k���JU��+<5�I��Ϋ#���.L��)nY��i�jj,�'
/����V��Zc9���j���C�ۋZ�ʈ��\讆����P�um�R
C3�V`œ�e�2n��w`��}��w�<��r�aZj�ˢ�]�U�#���_��t����D�}�����ߨ���0{(|��_��˽C��T;�'���1����ςUG����jf�|8����|~<�"GJ+|�P����2�E���8�9R��5"�WAMBq���E	���a	��IP���{�US�-e fN��wP>��o��s�Ap�-:m� V�}b��C�=��Ay۹�z�P]�F��w�W��BJwIAPHOϽ��#��b��#˻�������
�V�{��__�̛�PZ`��E�#�*97��!w뷽�`�3]��5W1hCQ��W�}�8�C{��!��
u��J�x���f٠8����0����t7�
r���+S��Ǉ�Z@��`xu^7�fvV�;j3q�H�����ț�����|��D��,������+�[�v>N��3s��&����>��}H�����qj�>ד�k՝�k��ŮB��#;f%7��8wi>�ĺ� s0Ԋ�y\Mopl2�L�yc����/wf���������>.-r����fZ��eZ4�!��w����m����ѢA��!�ν��=XDu�c�<������Lf�g�x��1cR3�����gs���?���������k��>LM���c�sA��tS�i�p�=S�X%����3������ho�q�B�@�O�ܟ��2[T�>�y-P����F�uH��M���`q�[!٫�yB�O.�:JE�ܗ^�њi��U����B�Р<:����:����EG�6��>]�75n�>�ս�]�Ċ{Qü�l0�{��+h`��g4��e�������J;��%}�m��^���ѹ��d5�A'��=wǢT�����$d�/�W���P����7U��!x��� ϼ��][�7�.��	�.{��r�� ��ΎK0� �d8���P{\C<���@�]��
�ddv�{���>�w��]�����Sܨ1㼗Q��}���"�]��Ƴ��蹗a\�6�`Lh�&T8��w�ݜ������s��T�ak����ɛ鵰�}��r�#�t�=���+��&�_��������H*xU���ta��5�o��6���_�1zԳk3X����?{C|l�"{�?/�3c��j��:���E߹սO�����o@�5OÖ�y~�N���J��a���O&Dtt�ug�;C��^��{��p�#��@��wW�/:�
�Q�Ұ��>�8lC�ǵ'κ�W9��@�����=�C�5�z�_��/B>���_�wV�_�Aj��r+��|��u�Y��&<����o���@��97�/v[yu�?Mq�r��5a����U!����|�����`��v���*�T���_tA�7�!_��B����G>��V����8�.���kZ�����ׇH���A��_ȡ�5�ΡT�g|s5W�d�ce����6�����x���B5�4���+%/>�����ۭ]��L���h
�7��5�MeoT,�:��4[	o|A\_ȏ-��q%L�z���yq�������+��%�1� ]��� ����m��`g�m�c�����T����=�U��:�FD�����aw���)�wT����>�<�ޛX��(׮��|�J���~CdP�*ѱ�
�wnZ���i�WM���P����%�*5�j�*�럞;��_��TG��Bͧhg��ْ��Y��=��4~�!�I|kN������=����ա_��۫��o��j�{�؊�1L4=t���:}eG�S�B���G>���_N��Z�H��cځ��3���MO���?{އY&����κ�6o�9ƻ��y��n<��=V���ԡ��%���)��|��ˡh���y�f��6.S���1_!��]�Cb{�><=s��j�e��v��G��,]�v�é��N�x+/��5||���!��Ǌ����c�t1M��]F�P-�n�E��ߝd�����2��^��T2����cĲ�iC�]Y	v����(�}|�9�_]�e;�Y�NQ��>�m��#��U��*��<I�5��ӎL�1*��O���ח�_Y�xRX��}����A:m������V�{�~��F��=�ZE|�
F�l!�~�R9�i||�Cm.�!�^I�S��w�Y�9��k�f�3P��exg�:�_e|����d6(�Ρ_y�Z2��E����f�{Mf�W���z͉����z����?#�O^,�+��}6^ok���҂��~�N:�������#|�Dv<��\4h��S7�˽�):~K��O0V�+M}g��?�X-O'h����m�I��~ً̏X����]�D��*o�7�u~����?�X~j��T��<�}�ð��qt�ƶ��o�X+4R��
�;��:ȧf��>"����u���%B2(i�T�B|G{�kh
h��1[���`�����l��Y��w�@�}J{p7W�����|��ed,��N�y9-tr���Xn]�z���/�|D�6�Β����L����j���Ѷ�'���#Paۮ{��~��¥n�Jг�Y���Z��&-�y�	S�xX�0±��wz���
�w �CK ������3M+O�ի]����:���h�BZ4]�_t�3\�yŉ{B���� �ղ�9�~	{J�YO�P����>�K��$5A�:=���3�y���n�v��v�^@k�\;>j�Wӟ��Y��f�xD9C���}6��7՗��3�����ip�ǽm���9��9i����T���/S�'�q�;�N{�V�SE�-�b{b���|�u�����v@��Tt0�W>�x�f��P`�}�襞M�Z�ih�%��|J����Q�8�/w�4R �׸;�[�[ε���dU���B�i��g��n�\�8=�&DE�!Z��/�x+3�h���{��l޶İ�E�]S�{�۪�n�e︉���w�����Q��3��}�)��np��X#��M����E.�wJV���4n�M+�qo��D�a�g���X\�x�n\�s��������^�k#�KGzzU��)�Y���g��
h��~:m��r�\���3Á��n�`h))32/�.d)tf7���'ox�ټ��[�N5��5�nF�ֈ�<�I�"�­�������-���������Q�g];�&�g9���0�s;z����9+!��s:ɵt�:չ��1S��6��Q�!����!Qzs4��-����u��2��Z�mgƟ�>w�*�HwC�9&X��^�vfb���r��G؇n|�2����IW��h#����]pR>=��-����1�	���f��k�:��=HS��trlf���!q6Efٷ�H�t��{RV�͠FҦ�bYWي'@�a�5gj�#W�7{4U�1�2��Ä ��}�F(��JL�h]��a�4�h�2���G��GG5[0�ŖoL�Yx�4�w�5KI=���5t�&t�e�U�����C,4�.�\��V�Ρ��2w6X�S�w�Q�:S��� ���X��w�X��6�<[�g�Uv�*'��i�p�� W|���71��\\Y�d32�܆y�"ѻ��rG��3N�9�c��{���a�6�}ݸ��MZ�r�Dq.oN���#�׈ɘ�j͋&GO�E��dqf;�����MurT�y�|�`����ý����ة�vt��ɮ�s�F��	�0v�r��J�f��yf�Q�Z(�4Rb�����/�����*�`�W�nV��/���n>MBT�P7����1��;����5��8����<�֯#GK/.��V��Ǻ�m�����+P;�T��n	����G�
�>�	���r��Y��t`�OD�\�16�����i������ ���hs�F�uMH�]�·�JͳjЩz�x|A�%J���+�8��Q�*}K�ͻ����|@݂�&�!g,�F�t������uv����m�6�J�)��x��	1k[�<;J,�ʍH�1���xxJ�VR���ou��d��,�(%�����h�7��s�9Wa����b3�h�s���xhm�;h���t͔t�+�LGx;)�踃Q�Tn��kHr�ȃ� ��mj�$��,^[�t�^�W��
Ý��
���2���2�q�{�]�N���˹�Y]w(���X����Ã��N�����GU�W��� |*�PG�B��*5+ګ1�dQ�1,-��m<�DU������%UE��ʳ��
(��TKj�UU�����TF����1DkF*��""��*0QV*%��+j
��b�Z�UX���Y��P�UV(��+ZQ(������(��1*+�U���j*�)F(�@�-1r��k`�U��UTb�ŕ�A-�j �AV"�fZbUQ�S��*�"1�� ��E1�H"����+��B��%Aa���KC0�TX������(*"ŕ�V-�QV�o뫼���
����^�j�g?�U���k/A�ޔ�i���o�q���8����ʏ��&]6����eV�$Ǔ|���?�;P�z{d]fC=�����`����$8h#�yhN�&�^c]*��񳞂��K���V�y�Q^���ѐ�?Z��I_
��u�w��i3	�_o�=�_�w�P�n�7U��^!��T���z����D��q�4p�<+B+�FCJJ�����]v��z�]��=���@��i� @�e?
}���Ah�"���+��-��D��v]��=�C���tC	��@0����D��Պ���Qy}����d���qʱUr�j�u�����M���֕���7�Q��hEX�^N����DN(g�6���|
����H��B�J��a��]9zav�vV9�/�羥����z�'��@�.���־6�G٬�T�VlS��N��7袖m��}_eZ�+%1�����#�����_;p��.e�n���0�s�6(+��|����](�2��֮0�n��|�Y���Y����U[�T;�4�ҸS��3�
�Z�)55s���a��k�wS�23��$���Fؖ;�knI�?|M�et�6���6�g����2�+��X�V�Act�o�^l[�OS׮�y��GʙW�/���.�
�|�ƾݬ����-iϧ�?��������V��kS�xX�q5�ad$��`�=�������y��~yT*�g�~KU�PK�6py�bJϖ|>�JS�3ު�<��ų�a7k�(�VW��M�!�S<b�]�}�+���rJ��dMU���/x�^���P�/���Eq����N���h8��2yėW�9uj��os>wN���:���E鞺#!�}�-� �[�M�Lr�#����� ��4~�!Ɨ��}�x{�C/�{��<�[�/i�]T��)_M�7r�a0G#E�D⤐Q���~-��.Z�8$�ճO�w�� ��B��L{�~'t�1��c"V��[�\�)��G��w�s*RjԾ�yO�� ��,���}�p��O�7ݪ4&\O�:Wj���jv��z�o.��
բd�[���=��&�X9��I�7��I%���Z�z~�1�<�z��1J�.��˲���_��L����rP��!�~�_�s�U��]$o7/�h��p��wj�j�(�T��k����^}��Mܜvo�X��E~#�Dn�(@�wB�̜7�Kq�?K�m<��F�j�\�Z��[�5�q3eI����T�זmKý��;eK2R��`fZ�J�(Q�x\�r`�[����OgH׹�+�Ă�O&��U�N���<���ѽA�jߗ��OPIo�?.o�fG�����KN��h{����Ol]���p����o�U��s'!3!��:�䧲�*f��O�1|c޺�������[�wވ�����n�KK�^�؉�5��̬5�Mo^�~y��ۢ0}��a�ȹ`vM�ˮ��o�ǹ%c����ʒ�������9�gNC�E��N���1P��A5�S�&�z�R[��0�?��w��g�w/��]?�c�����莕����zf��zmڷɺ�Uut]{|�э�O��,]�Y7�K��>���M�9�$��ڗS�kj7�-�a������y��vߞ�����显��J�H�ٔ_�0O]�ԓHl�8|�#�I�a�|)�����X�w�`����;wW��3�&�T����\6�<e.GZ\ ��~UCW�mE=�{�\_]�����ʍpw�!WT�j�q��93$Β��p��|�}��<,UN�*�^	�y������Q�0�>�G6��0��**�)����N���MB�,�۸�t��s���w
�,خ��(c���u�*�e��j �7zGٻ��d�����	*nk��orD�i|��	��ٶ�󝢬�W���y�C��U�
|�T�غ��w\.9��R�0����6�u�[��-�C`���ʯ����ث57&P?���ZīuSaq]���b��x`~	|�rnnt�8�����^����,��T�/�C�n���ԝwl�.�������;|.����r�����[����<��q�'�ѩ7�b���8�X�F,�
o6U�W`�y� �r�Ս�}']I0�����ux>�����q�)��E�	�Rj�jܣѥ�O)�ֆJ�����w�\�N�O����y�:����4���}��w0��/=qĽ3�ǿfJ��&]n�K��e�>��=�՘�;q

�#o�!��VI@`ĬI�us�%s<�y���������G<�c�o�,l�
�k�+=�%VU����H�ٴ��_��dZ�@�՘��zY��غ���B���R��o���S��>�&�{��V.H�7�U�2��;�= �;skH~��a}��*��^nbU��v�Þ0�>Hh�|j����nM�}K��ɞ���3r���2�R)Vc��]��4K��C׻�B��D����/�����O�SE�ӭ0:)�ܛ������o��˼�3��u~�ؼ�4vlo�&�1��h�t�!S*p���ſ}S\0{vbP����zF���z$5�m���bAv�/Ϣ���}T�f��$�K�1��c���*�lc�=��v�J��p�z�n�����y;|3^hȖ�A6�h3_J��cT�b�h}o�	:ؔ_{<,y��A�0viZ]\�o!���j��wi&�=Y�(�{���Mwy�^$��Vs.�rq�7B;
�W���<�u?���
�;�����[�F�%�Ot�K��Z��o�eEӕ�����xJ�jt�ۏ&�b�JH�BV���$q�O�O�U}V;�-�������?O�^���x����e'��d#��:1<�oE����2���8и�o������Ρ2G��Q��^+�+:_[��Ȯ#���A��È�dx39h��^��Qӫojp�}wմ2'�p�^�t�<�x7�E_���vSs�gMx:��-��'z�^浊(>~�xSe�	rO���^�r+��J�GOy!)p���I���Y�w�\�]��n�$�S���IRG�喼��չ�����s�vc�G-�޿�dF��5N��̜:<���w]y}����ѹ��k�}���ѯ�^��*�*�ǅ��lػ�����c���v?&��0�d����Ey�t3S6��W薈��g�J/[�sy8b�b��
��e����5���vQ�9�����Z)�������,��HL����t�@��}�͔ml�0����3eCy�v�w~�mu����?��n��X��g�R�O|�k�\�F~o.��>���@}B��I�}�ܱ��}�z� �VZ��<��:72��M��� �˫F�,�Iֱ	��W���
y�і��N���3����O��󩼅NC�j��~�����ݹ���]^�nGZ$�e����`�����*ީT�K�qη[yPVΡ7P��}!�mђz}���m�kKp��*v@�t9=����{N��z��n��hjmZ��X��Uu�|�`_\id_p��dR��Hȃj��߳v����r�>+�#��i�.��o:Bk�bI��7�1�3��8�{Y�fћ"bYn����(��փ7��p��;Ʈw�+;�]|;�3����A7X�	8�q�ͮ=��d5��Vj}��z&�i���Jp_d5$Yfg@�fK���n*��e����n�,k�ܴ��:�l1(�hbd�*���I/s�t/��v��f�=�1U�vШ��g�{K���I̥%t ���kE>�\0]�1�s�zs�w��y�O��X`�,�����z5hפ��kΰ�ڳ�ʹ�0]\agD:�u-����9H����s�ǖ:�=1� ��o���1�wK&���K�y��������hp4��@�곪��t��i]`�,������La�q��(v�#-x p��N�ͽ(.�{~�{{��)Y��{y�Uϼ�X��=�L��6�9�W:�>w�Z�@>�2=���&3�a��`,N"�_�㣩�\5hV/M��ɻ���s}�:��*^3�^g���m�Dь5����5�#쿺��rc���b�_N6��[��M"��]ƹ7�xc��	���E��*�;�K�v��E�u�,��S;q$�\�N9܎�t� �ˀm�q\�}UUUc��"�W�}�k�O�ټ\��F�)��'|��yL�nd�l���@��3���C���d�Y<U歽wF���q<�s�p�:bp�ȇ1��`�;}=qi'���o(+q�_c�קOp�M�vCt��U���^�6��]�c�426S�9Jё��~͒��I4� _���L橨�Zr���~�o5����͌�c�����X!��N���,!u ����v�go����v���,f�wTm����je�c��U�&}�)��g:-᩸�Wϼ�]ch�f͊����+J��w[��&b5rb�C�����9�cʍ�-�d-���#u%���^:)��i�)8S7��j�D�`bvF���K���b�ot�p� �������u��+�OI@ڂ�1�ͧ��g&�=In����4���p��͢d�-�tk�Cu�vGd�6Bx�������7�/A� ���vQMŃsr��8�n�ѩ��J0;����x�ζ��W���H�B]@��t���5V�e�&]
l��ٍV�p`+�ңY��R�-��7�t<&袅��G˘��1m2G�)z�-���wU|�U�SM3���F�DX�N|Q�f�����k��;�"[�L+w3#�]oL����,�Ծ������/����Il��l��^���������*�S���Jy@K⻝F�uә"�+x7L��W{�MԢ/��D:W:�����K�og21�W�A����e(�3Zy����Ll 
��wћ�ƆL�a��m�[E�����z΅�R
;���Հ�%ֵ�b��h�ۭ}����t��wF�-�'g~�{��ç8:�oq��Whyf�[�:�	�6:=N�F����,���{�w�f�V�M Q(śL<s�>�y9Zu�Y�X���§əq4��=R��*r�&�K�w��T�@s݃f��v�U}{$_�,g0�s�e����[U3�ʹ� *ݩ�7�U�r�P?&��J��ue��t:`⑘:[�6�!�&�D���^�+�"6b����xl'u���qP�����R��os���*V�v]u�Z��L47�/f���tV蒞`Տ��kw+�f4���C:��k��3��}O4�������L}�X���:
��;F���ݐV_d2�VEO
�b[�F�<g]<ŵݶٕ�I�$�Z���x �u�DӜY2)�{�vB��ت	k>8�	���u�{uh"�!�8<��G5p��lR>�VV��RW�p���o#�|�E�՝�+i%��֧��D�X�ފd�7R��9|������\w���q�ͪ��8{����Żjr�pN����G��u;la9Z� �γ%��R���G1�$[�˗�uFj&�+r�rt���i�s�@���Wm����ED��[MC��~�x%f�(�K
fa���Mdܿ�*�ݱU�E
EM��n�@��e[�ϊ�]���xҬ3�2u^�;Wu+�}0�=���n�P�>���h"Olm��T\eY��O-,�T`�T�U�1DkU�ff
��[E�)CYYXU�R%��"�R��4�kZR�&4C��c���
��[��Z�1Ac�0nQV�\�-iUX[Lʸ&e1�EbV�Ȳ,��4�aU�Q��][j�P̲b*�)�P�	�b��2�L��TEKm�3 �Dr�.Q`("+F�Y1+���pjbE�.#i����Im�A�]%AMZ�]U+CR2�L���mUEcs�/������)��f<�Mǌ΢���AQ���*�Kz��"��n60>����4�d���0���}�}����S�����<io�qb�W�u)Kx	]�_s^ʞP���㈛�akyY^1���#���h�ڋ]�w�XJ��v�r�lϺ9����~�b���#s�V�~4��`�����{t��=Y��AkY�M�q�Q�'�=O��V�l�y��e�<8�b�Gk��M��]^��}r3Vׂ�7�����r^y�"��G_me�s�][�����ښ�b���4Y�my�d�OvOKq����5]cR�R��C� ����1:�S����j��x�@���rVD����w{��()cվSM�߻�~H��0��쭌SF��+K%�NJG�x�����2.�qT�x�|�$v@�n�W�B�o�QGl_{e�m��ă��a*WU��LV�7b�셖Q��7��ҕ�pp0�dĹ"iY"�S��ܱ�9�f'Տ�z�h�%��ݹ��y+��c������n:Uj��ƴb���Z꫾F��G*�M�[�;�p��� U;�ja����4������%E+7��-(��!�Z��u��t�rGF�=��&�Κ�V������ ,��l^Pa/�Vݡ�J��fI(�g�(�~��g�-g�A:�Wh�+��\;޹�aA��'@�@YNmwv���.���dh8Ʃ��P{Mm
+���Ҧ��hY��Ǯ��z��֜�������_{=�4�X�sz�N�7�����������j�~���gM�)�&2�\,�[�y�A�U=|ԗ\���+:P��{��m�y}>�z�_*�,����Խ��[P�s&�P�]��]�_��F]�3kH^�˸	��!�30t�g����$`.�3j����{�I����5G��e^¯�r��]+�/���7Ӣ��.OE=B"P�W�ݜW4]��V��/�����9�'�2�l�@d�j`�A��L@���-���UYήs$��2<8�䇛\.:ȥ}ڑ��l36V_c�n��ݯY�/�1���g���	$z��Y�#�\Y��Y2SSn�Od�Bu�#�K��̩
�nF8��>������l��*�8S�+�ʍp{rpU}��� �f��O;�9�SǔwεկX���0Ga�����a$��Ë�U��}3�m��pa���_������)��x\�{�y�>�:mP�Tm�[h���H�c�E�.�3gO�'e�|�ֺ�nļ(@�f�g=U_[���|��i]�۾�����
�ӳ�}y:����Y�\�y��]*k9O-�GFw{��+g:d`�'v���D�(f��gd��%�&ۥ��6����7<(�Y6�k�Ĝ��oخtW�qa�s�ᶴ��p��ǜ>=[Is��̫���݋�b�s�}ƫQu��^^Knf"8(�m��~�{i�������{���������I��|�@��������r��,g�-��.�s��������O+�چ7�$�Y��y����TMn>Nf�d;ʵ{��m��j�h[�5�n@��{A���K��w�W���ğf�ԅ�j>���fp�#����z��9�4�#�w��Hzb�q�̔:�p�.����U�s���|g,k�t�����o�	�
�1q�Y���n߻������4��{�װG<�i��6b�k�6�#��׼�#mLg�y��l9��|������}�ҏk��ș�k����Td᥎��u���MA�eݏ(=��4�+ji0�3�c.V��n�7�'�b��԰���-��։�+��P"QC]ћ�)cN���Xԏj��&�P�3J�.O���;:/$�1�N�{ɷη}t�w��e��4C�,+�RN�º�V�k��E�^�L�}�fm1��" ��u�3#�2����+�$�l���\kU�-��k㉛*^T᜻6p���קfB���*�{��b�`�Ԗ�xl/_����&ʗ�o�\��Ӵ�.�;�K�Ԭw��<���!�ڲ�m%��K*)%�z;�]j�g}���Ux�������.���N��n�{dYF��o�s�ʙ������BsU�۶n=��fb��OU�ݔg4�B�չ�����5�=hy���Qyū�b���>�<!�zKʟ*堊��f_�g����������Yr
�v�{.ט�E��bvV2c��d�7YۻW�;��2|�e-Ɏ�K�$h��nӱ)Nݼ<��H<U���a˻��;6
�yX�]�V�b����%^�Q����m�n�~�;��SɈ,p��	�)U�4A��G����O�x}�-�G?2��r
����~\=7:�b��nmtn�E�!�;|��dO�߸�����v����#;v�k햨3�rG,��Se}R��%iap��k��5�\�vg]	�:��p/jp��n�}�N�{�J�&�s/�L��?�TrWDT��������Ski5��Q~�9Xu���ց���Z5�e���rn"��6�B�s��k���LO�f^I\}�71s
$�1g��hzϓ���V�>+Y)��o7(t�P^��_u�GP:�%9�/�a{�}�=P��)�������]1s��#��}��̷V��{�y*X*{�Q��b��N�{��c�Vf�d�;t�vS
�(n�d5���ڳ�s%@�n�f��{�{#��
���۴&s�Y�y���K��ŐH��@����)ꍠ,��k�V���Iղ^R̃�]���;�8i1f�;�_��[���F�5���9��T���	���X�t)X�_�nIe�̹�n&�E��ͬb�CV��yO�������f�/Q##rpɴ�Si���Ɉs�5�S޹&���hlg֜BK.:��R2p���2����W���@�������9�A�$���kfй��V����Aa���q'��eHn��j�ǉr��=��zG�T�� ���t��.�I@*�>�n�ڮ�����jb�8n�;��N�K�7�zy�f��fG�qW���L��i싺ַQ�C�n�]�\���r?D�_[��{O,v�uz��L1����q��S���$�˩��C���ۡ�E��a�3�h�B]N9(����ts��g��]Wj:����Q�9�_����j�&<����׊��7�X��gNT3��]zV%�sGN��Y�W>���8r��Q�n^>�� �m�����U��K~;�F��N�:���K���U�g�'�9��1̮���u�%�����=ً`μ��������}����n����y�T:;����]��)�;�M�Wެ3|�ܞWӵ}��	:�I0�g�r��s��E���{�66�3�o�^�mԚ��ܢ�h�yx�۽6[�e�7{�}�@�D��d��;�����_�9�ކe[Pv��������1�=1p����Λ�Y�@�Л6�%��Ccܷ4Q�9[�=��JU�%WDj��cE��Vmʞ�]3�w�P�yf�/澷���񷝀�x���\���Q�������q$�nCu���N��gv�q��uy�}ooo"��;ɵIh4nV�71�U)�`�炙V.�YÝ��cR����p� ����`c�o��|���'�Ƴ��}W�j�2'��D탇;�+�^V���%�I��u�G�ʥf�-eWg��S����I�;��.��|�o���&.Ǯ�M<v�93�`��ACsF�w�+�C&7�ЍE�uEVƍ�zڎ��̌+�LN�{&u̹��ʫ�G�sS�k�lWV���iT�7{$�sQ��A��_�f�{c��b��6�����~����L��R�!2���虦�-�8�?yߺ�'�z�gy�W)fǍk�`�	���,��!����Ii���P�/����6�_=��ՓzM
P����C�ld�f��fQ*0]9-��,eg�f��ת'O{������Ղ��Q��W)�z�[��q!3L=�T�G��i�7��-�m��J�w9������ǝ)���2�TΎB�)�����G�w�ݙC����|�sU�G�x=Ր�T�[uz��6�;4���q��A�(1��Լ�ֺ/>��;�G�'ۂ�B�$��}���n��=]'�}ݷ�'!�wdt�ӿ�g�n7R�y1
M���N�WR�s��O=idt�'����##�5Hk������ܬ�������㿈��PV�`�����}lc{���]Kӑ���A�(��}���e�YR����7Ac�mo�=7��̛��t.H���,��� nB�����Y�����%t ��(7%���8d�b� ��=>��A��1X��d�yQ�͋^ʽM.uyI��:������m�u���.2"B�7id?�N=�����q{�ԗ�y���F����� E�v��imaޙ.�0-����	��}4���(�P"l���� gq��9�юb!�V��D՗���K�4Z/q��;O�j�9��x:��Vޝ�DȮ��M�����t��*q�2��;)T���W��c��X��*� P+C^�ۛYï*>��'p9���NMof.�b Xc���E_`���M'L�vu:&TJ̼���vd�}��3~��lb�٤��4s�E`br^��[��W-�ʆr��@J�f���ûQ�ٛuY��r��
�X郥����*�P�F&\�52��Z��F��y��Sh�y�B��Ӷ��-�m���.�ǰ�)��ə�S�|�<s��wk�5��U��Z����.m�r�(݌�r)n���{Zx�5B����yj�x^�r��*셩�H�v�}2��-�|g%��M������,�Y��q�i���h���;��R��iG7F���VkG:M�-Y�*r�B��z_�him��U��px�jP�^�)T�N��]�Rn\�Yzy�Y��=O?�ɹ������Yh����5��/����xν���0��-�O��Ha���nс���6^[S7R�{k%�UlAѠ.Q��&TI�Y0�j����	�^|�V[�J�BPc�ʕ�.����ԏm��N��
�_hy�����V�H����J�ȗ�hj S�چm�ؗ�)�9t�c�mL��w]�]Qb�J��k���tt���MM�V�0��F���C����ܖ���u�	��KF�{@�Ң�L�ŧpoM�ɳY�I�Jŏ\eA�z�{h��}��TU^�o2�9i�J�����t#�Hf��p��1:����I�x��ԠB�m��8<'kLW@RϞTa�̚rl��
�)2z�-.��laq�J�
���O����/&�(b�NJӋ�53hh5o��_h�[}C��7+;J)ř�- �n�K۲P�r'd\��V�zb|pσIN�|��;�7R�Eft��sn\٢��+Ta�$�qV�ż�/� j5�����d]r��vp�4�m\�xi�2V�Bv7����:&id�F�<)  I|Q � 4��)K\Ehc\���c�љ��d�-2وb���3���EZ5U-��-j�%Tb���PC�j�DR��\�[���Q���e���3�˅���)iE������LKkeX������h�i�f6�e��I\�mW32՘̙V��icZ�����Jʘ�J��S0�1�¸��rP40�,�,�TDī�(��.Qh�mT����.+m��e5R�ڰ���-Ƃ��Z���b[bխiE�eJE��2���*�V�R��-kTD�[Q�qƎm��a��ۍDb�iq�,��K����R��kP�jde��j�Z�e�QqmZ���pnZ��Ķ�Qq�0�����s.9e���h�nV��[DӉ�H|�#�h�T~B����pO�E�@��U�<�of�����n�S6�k ���v1 ��<�bn�Ec�Y������K��L�z���0�`o�-�{�b��:n*��|՗���j��������}�f�-r�&J�c:n�NvX�B>����(Y�*1n`�}C����j�2���N4˝�ˬ^��#��Z5��L�؄�����M�a�y���u�%�#/h%�)��1���λ�l���)W�������q�������J���2��\���j���k�P|�����']I0���2�3]e���}��-.u�e�\��3;Edu7P�}X�x�P�x���g�M���l��`���Č���j}P�M���r�5{G�$ي���g"1�C��q�d�b�z���U��UL>�2�¯*�K����@�q��[���]<*#����e���f��{]�`eu]ߜ°[-/�[���{��,.]������C�ps�s�7\|C�X���Ln4oDӅA1�á�"�c�ۜ����pѩ�ʻ�ͷ�m�~�(+q���~��TsɈyf;�!\��V�'���w��{F;̵;jV������3�$V�Y�M>����^͗�>�h
j*���c8{_�st���0��b^��ܷϬ�7-\B�e�7��|�|:��U��j�m�J�j���=�o/�eW��2���VF9��~�����T�e�|�ǆ���v���~�O*����7�6Ɨ�ꓽw:f#W ���wS;c�� �Z`�ԗ�����K+e�[���W����cւض��	;��a���bnJ�����|C=N�<�7����M���?{~�7�㼩M?Q#gA���u��kq���9*�x��i
Vv���/�"��Qݍ�Os۰�1/G�k<���vo��}%&�VQŭkO;�fӊn��V�[��t��x�r�n���E�J�A�fu�U�{�XA@f��u;��Sk;V7�'[��-��D���;�M闷��0s'��4+��m&��'m��;��b��(����/�9җ�3��2�G��'���!�̏gr�U��孺����2S4"m��rѡ1�y�R�X�U��{�ŧ�Q�����@�Z:��|�gj�rڡu���OvN�0����8��喜�s�OK����M_�G��)���8{�C��k/%l���+�(�DU{�WQ�Vd�p�p��<���q���]�>Un�x��\-�2=
���0���v?xʗq�T���(���2Y��~��>����װ�דL���Gz��*�b�#�U��M��F�}M!I5��s�\��m�YX��9ts��n+���q�FQ����cx_���&�mt�7)��f�F;��U���m��͉�O�������g����+����k5�M��G��y�t�g�4�s�N����+!���N벙�����a^-S�{W_����:%߫�}D�'�D����U�-�ϼ��}ݏ��LQޕ����>BF�RF+ښS�^���ƶL��($m�
���a|u��՝_V���������t�����.X��q�.��0j.s��T��'��u��)Oo�s�!�6��.D��a��cl�@�W�ʔ�|���pE��)�+uu꾐շDI=��}��bީ��{�C�������Ỵ�z���\�"o���-�X�\��mα�;��y�Lby�<du�C�b:Q�in�;���!T���5��g��̰lY�r��Z�Ќ������
���P�`=�T+{��U�@�X�{�.�%�r��kN�]T�{͞��}�KM��m�O�����^����0:wVd��\6���vo�Җ�~o�W^�2P�0�G�xl�y��۱��vc���,�+���Um.Hurx��K��/���V'�C�9�Q���c�rWʭ�����xo|�Go��{�����Å�7%����	���ϒ ���х¼_w�C���b�c��y��2:y��$e���H���d�ab_V�E��/5�Y��Sꫫ�ei[I�9NmZ�� 6=���'~ܨ���B��t�O��/v�=m�:C������
��X;�s�s����(Q*��H�/[�:O��u�O�3ޮU�*;'(_�`(�������̝}+����e�Sc�=��w��#��#�k�@��`�+o��܆mҟB�t�+�~1݀��������*�otC��#'�U8��&u�e`��#����؟dɁ���ep��nY����k9}C:I�r�e��-�vL������W�۾6*ѻP�ӣH�{G��/�����$��=����W���w_>\���>�S7!xd�+Z���f�>����.ws{�x}_[��"O�PI,T�wP��4�Z��~M��I�W���l>ᜈ�iLC��Y��Ywٸ!Ok�ɊtΧ�{2.!s�5���謑�p�\�*�V�x)p��j@�ä(�s�1����M�Y6ۮۑr0v�X�o�Ak���r�:S7��mp��]�fXw�m����N�)�L���jM��}���~�n��t� �����3�����ܵ|���V��1�Lfip)|�#�: ���O�=�8��iR��q�O�t�_s�S�2K��qw�.�u��MW�
�Ae��^܉x.M��yn��x��wsNA����Kއf��wU���a�|��S&ѭ�.����,E�fvо�)�e������KS��9���n�>�C2���`!�Y�� �ӵ����nQ�tR��f<����ο�J��L�����SY�%�]}6��W:qUwc�r�u��	���i��ˤ�t���}Au-y���9+�@w+��9�3��u�Jmy����S����s[�~p��B� C�|��+���߆v�{&�����l���-=W��E� �f�^�0o��=�(��M�s��h!N�^\R��;1F�U�cE�%����|�佽��䗲Sܮw6��ֹ���m��m?�3��ː{��������8��pA��7v�,hɴ�AO&!A0G:/����u<����c��B��3~"�ڽ:ǺAB9����=��O�{�.�[K7��CWQ3~+hp�e�x!�vV��F�`���G�V_Q��#o�ۥ0�=FG�o�S���΋h�a�J�R���Y�AQ�ɭ���)ѽY���X���]I-���=m���oYR�'X�8�p��m����H�j/ڀ��W����®�*&���3���z��O5��?~�fvP��:���D�%�߳#�x��S�V&;އ�5�f=�6T����qQȫ�>�S�d{�I�~aʹ�.L��������G�v��tP�Z��� ^O|�����vE���3k�Q3y���;~g`fZ�+����\|v瘯S�ʫ[��=�3b:����@M���i�'&5�  V��[�_���o��'��8u#Ec�ٹ�,_w�]b���˺u��9:?/�v�Fj0��S�Iօ���9��������8��~sdw����p�@�P.s��MU{=����[��
�q/,H�M|��b�|r�K��>��? ���n�E�X��}&4μ�c���X���)��5�T�����I��v����Ϳ��#������,�e�&���^Uw�ݎ�K%}�{��A�Jt'�S�Y�~��Z�!J���@���v�/"y$�޽��n��{gڈ��o3�:f�|���1���Ӻ��ڍ���m��>]{5��s�la��I��"�������^�1ޢ���K\L����)���{��gzo�D�`2{u�]�h;�ktI+��מ��|��-�W!�G��T�W��D�v�HA��wIC�����pƍ�J�ΖV{+�;��Z�k��j���pWk�7%tFw���t솶tк7�������{cW2��#���5�n�'\yb��'z�n,T�Qb�
���zlJcw�չ����]�����MXW^�z���NQ����lG���U�3f��\��-�Qf��Ҿ��K���+��j��y+;-����,��\gm�,7of�Q��yr�I�r�V4�H�2�Է��U`��.��Q���]VW���c�ɮul�с�ܰq��v/hpV�)_����:bo7�uSC�ˁ��a���=ϗX�C��+p%�ۯ����n=�T�b���(��uz���؟3�c�xX�����Ns�LJ�������;��߻'V�0����S�G�ogd��f��彴�u���M�:�P�,��mJ��ף��^;VZ���>�1����͆F�.�8x��A�t�P�V�o�mN��Bd�(&��u��F���q��)���/WM��r�#�ك:B.y|�nu�c>�����/���k^��Ƥ,Nt;R0r��TsɈyf2>�]��%k��l#�
=3���gU���V�udzڶ�얊�`3�b䀰��eʏr�����n��*wbR�i7*
�ʺ��4�t�8������ـp�U��l���2�[��7WQ��o;���ҷp�]�؍i�=���7����9��Y�	��;�U��T.�-x�Ж�%j�{Վ��Y)J��3t�Xڽ�ۦ3�k�m��������-���+S�q���co'k�k H������(� hO�����]�ظ;�w�`o�s�r�����&7�Z+MH��tƄ��0N���I�{yή�T�u��*T�!�&_+h�#��Vջ�!�0�w�k�k��썥2Cֻ�Dܑ�Mb2�o�jud�}���k��%���4l24Ј��w3�e �wbq�	�{u�w8�S͗�E��P�
Ӽ�u��ʺF>�;y�lc��宫Œ���.�ɶvM�4[�
J8+��K�CL��h/Yw{����ܶ�q����E˘�:l��/�s��d"+����"��d������/f�x��7�W&++���r;T]��ݭ�h̥ھZgj7���}��W���SD����b�r�V��v�o��;9�MzWG��k��N.�RQ̦�DsU]�ub2)o7���X]%�U&�*+�u��?$�y<��-�s7u��d�&�.Q�C��\��0�f��v�>bm��ʁ�*�-��}�w@�i4e�n�k+��#�ͣbº/z'�q�:���&=›�xR8ca="��b�T����Nt�l��jc���ɻ�x&��6�5��6����"�:��ΘzK�5�B;4j���ܓ�RuIo��/��d����ՓW��swJp��Z�i�
�\���W)3M'}�̵Wo��x�jp��7�r�4�\BͿ���ˠ ޢ�X�1��C"�7�kru�af�o/��mܩ�jxX؞d��X�A[��t��u���c'.��#��
+/��U��Dq�@\j>�7_`�_/�T�~�a/�/{�ǒ�:�vc�y����cJS9A3{%�jA=K>� �Z
����@�ÇH�Vp6��YO��'�͏4HuVi��U'"k�0V��<l����\�����3s7W%J�y��}Bz_�P�Cw.�*��kVA�S-u�P��6P�z�G���kO��U�4�q�)�%D�_ P$��-��f\�r��j�,���-*Vm�Y���,s2b���UJ��`�Q�m���k������QS̭rы�LR�.5[h)\ZW)�q��R���Y[��cU�m�)�q�+ZХ�]\I�4�bJ���D��*e�����r�V-j,h�eL�k-J�R�W�̥l��l3r�.�Fi��
Z�G13���UKTjP­A�B�Fe)r���s1�j�ƣacUi����-��m��m���1�X�n8�F��EA��ҵU�2�.��tܔ*.5̪��Z�DDEL���T\���2���)U2Yb+2�-jV�Jܵ�kU2�aq�Ll1��F�V�AC-MY��TqmD\��eb(8ۘa�X��DQZ��i���j������ �8��'9�~���Z�3�c/K�j9}/�3֧T�k�e3�a�Ϋ|x���{V�)���������S��1a���5P�!�`�=�tr59��2���s�l��-^+�B�j̛������~�l�y����*:q��c�I�>��4�ё�b��T�^����vc�Fni|������eQ��I�i����λ���3z�*���ռ�S��W�h�v�!Sn���:Y���7��Y���fɲ�d�o`\ԹսR���{�3t�\^8��	�y��������;�Te��f��=BxX!�z4X���IG��o��񩞻-x�^�V~�Q]�c�ʚ�wv�3�c{�^fm���0{֏t�S�Kv�IF�|'��ז�%����#[m�@��G��S�h�]Qf�����|4l��9IҮ�t3���p��Q15m��<M���ܩ��C��6r�R�d��h�}/$���q9ђh�E�77/
�K�b���1w�{0t���s��|�q������W�G��]'b�����r�<��ޑ�;&�/���o"}�5�;L�����2}g	���N�z�m���z-��گ�D�A���LB�:fOM>�}YJ逯���ct0bt0E(���=�
�9�߁�{j��32����}Dn�V'p���\	�9v��'.��bmc����+�㗦�Tf�k)+K��W���[y�nU�n��f?h��>��ߺ|���{ʟ|����o�3H5�@&�4r.������2=7�6>�Qp)�e����[n��������kZ8ؾ�	���ӚtK�.w�&j�Wg����[z�����Y��J�+��-o��<W�!�]B���1�X /+x��!k��W�m�H7���!G��1W��75�ٹ��J���k��<h�J�0ֺ�QU�s�f��+�Ky+;R"�lZX�e���䞸�S>U�~����s]�S>�x��x�Ʒ,�~JU�~�K�n��+Zs��v51�����߭9�}�g&s<MhSq���vթ��q�;q�*��3}��7���e���]-����z�˂�:�ܿK.��ἁ7Χ27�7�k&�\�F�i)�ޡ��c�\�Nd?��oQ���O���K�e�@��u��,V�^ྐж�OX�^ٓ�o�w�������lA���Y6�����L��UnW����B-�@��|1��%1:ȧi��+���gB����:9�c�ڳ��Go�W`��U��NN\�m����yA[~��ՊV��c���7��aի�7��W3(V0�o���s�����.���G3ЩĮ��W��N�6F���f��S{�%e�s5BRD��%�P
U&��W{Mu��S��V���4�Q̉m��V�^9�T�4��J�,����#�O/&;�b�C�gUj��&���-��� ��
nJ�*w��yժo������2VZ��]}iͿ�p��m|z�(�ý�D�:�ڼ7��7��J�_Qb���~��C���U.���y]mq[��#�����v���"�/Q�Yj��)�L�j�����\��v?;�h��г���I�5]蓚�"�CG����x�����DQ�.��ȱ-�-�d�fv�Y�N��h	���>g��E��d�F��.��<����/y
�C�j���ӷ��ᓮ��c�+FtıS�^�o�ϸ���>����S��Y'�ݡ��~���:�D_,�R�ƣ�t�G)�n\��:]��{�J�TK6}�N�+W������4�m{�WpZ,t&�]�|����yt�w+T���D��T��r���qc�L���)ک�Ȯ�Y3����J9���Εt�S��u��}��LOA'z�Ю�mfַ]W$�3�<�� �a���^��a%Ő�Nq�98$�����8�����Lv�YV9�kڇ�\�=l�6���S�h_��~�9G>�y19XC�U]�{=��Jf���Ъʊ�S���v^�(tQꣻ�����oO��/�yv�j�I[i�=�ǔn�!Vi����9U��E��Ց'��\�n���Y�Q���Qa�I�6��7X`(��ۣ^�T���r?M�u�^��W������q	:)Dg;�Mk�[�0&��;�b���I�D�^R�nN�z���3���~�S��̹:�*PԭmA��#�lu���kN��W)�ڒ�*��ǋ���T.�M�ڇ��Ч�t��!�TZL��!���y�w��J��MF;t�u�cl�"�Z�}2�4�b�΀;m2��4�R�����tK�����{��0pY[�sg�,{T�[�s�~��^K�.퓦�X��;��{Q�;�gg���$���>���*EύkPww��v�F_�,���wY}}���ꥰY75tu��gl��,�g����P.#�W/n�S��׻��N�ߪ�|;�q[�k��7�e����n^S�<�9�\��nR��h띍CL�p���<3�t{}��)e�{2_K�s�-����&����b��b�k���]���7��
ܠ�'CR�j@äǢWg�U��z��9~c=] "l��e:�J���F����Q=�=��#o�p|r��V�2�SU�M�l>����]�^��f\X�tC�s�.m`'��,3�����ℏbG]���ׇOٞ��x@��K�=�|d��q�+���BL	�cr�Lw6`���K��f��0�դ��s�Ι�-�^�(���<_y.�̌�g�v�1����ot��-A˂S���\)�DpN�2z�Y.��Ʋ�w�|y5ڡG������f�F19�{�MkG�:�m�s��[�eP�ԭ!X�����wWY���D�u0�Ɠ�t��[�{ճ�z��~�>�u�<�y<hM�=�+e�|Z�Ǜm��M�K�W���Œ�}�mW��>��r�J�3)fO�����ӑ���Fo��օN3����;�d铯���Z���H�_��_q�.��|�Lm.Soݸ��;t�w%'	�w��9f����Aw�;G���N1���{b���{%������tF��z`ķ���lÀKx�t�Y��inuY��O�ܡ��ָ;�ޖ��k{63���RX�3_\�"L���w�K���;V.`����/p�f9��T�X���U:Qۋ�Л��@�`T�-�2iM�"j������z�{}}*F2m5�A��U��*��3q9���Vc�;q��xa���$��'��R����/ز�I3����[0���@՝_o���w�o�<��ϱis*��� �<�+��P<=��wf~;+9]#;h���<�p�}�%tc�8>�Szdy�<�ƽ��Ws-�Z15� �c\)�+����//ǷfǏ/�h�ʇ��]jM��FS[X��A�����ek�������P�9h����,J�B�|*��ΝB�qכ�&GY���`�����fHp��h����65oT���e�ܮ�:��@��*ur�u���z]}8�����ֽ��*�g�K�� �i��#P���ϥq�}��S��Ӥjg�A�
�)WE� +hW%��
������P�sC��W�Ӧ�T��!������*'Rim` >v�ވ������ֹ�}Q�g�ۤA�8�?z��ѡG�����B�[��J��{�y�t�k����N�9Mn�����C�ܛ�	w[�4��8Z��*}�o-L�ӻ~��'_�#�>�[&�]%��6]Qf�Ӿ_O�����;ʷ������M�����뚲���e]��S)'�υ�/�#6�RNAS�1RPe=����*mv�u<��m��3��dg0���n̙ї��u���̔֜2 ڃ�#�y��ι�
���o�J��9��U���}�R������ ��y���~ֽ�u=�cn<��P�ɇ�5���Q���H��������w+��ӓf*�Ӝ�^!v�¢j�ICm1\0](��d�ך�T9�������������l�7��J��I���o���7Գ����g�O�\��5�w��m�A��#�P1>�V�9p�p
�l͓V�γ\A��]���w2l��40^s��h�܉'e�W���8"����/�s�L�yfK�����Y:��7c�����K��DUhҥ0�:o��W��Ӫ_��F�|�� dw_vSU��Cb��'����,Т�����S��_���W��H�ɛM���y���h�Y�!�y�!��bc��b<�W�6�-�i���y;f����j��/M���#mx s�qӳ��:�����vA+����,��}V��~w)�B�+����ko~9/cN��a�'Tr��f����-��a�F�	�s���i&�<@��>�s�Idۏ��8������'̇���ne+���e���/F_���n���uΡ��:�^�'���� �U���7�G-��泰d�n�+�U����v@��$�evIk�ki�M4i�c gT�T;���� k��ל�-{(ZՇ37#��zЧ���l��c�d�J�Y-q�N���Z�\���2�$��&����*pS�o˪U�Q�VA�f������u�Sw��ڡ}��.���kR���,��5�"iXZ$l��k ���wD��7�r�횝��n�����cqIQ��d��e%�3�]Z�֯���Q/0��Э�|��|p�9�ݢ���om�ܱ
�Mm��67��X�d�M�9����[��ӸQ�4�r����)�X���ஆ��"��1T�"e`n�hZ�]M'�S�yWՒ"�ӭ��w4s�[yΔ&��z�FRYo2k
���tCe�}�%R�4����Pv�.�K:��[\��ul�c��B���M�!�]�unus�|Ԓ��&&rD�z枷0`�P�NM2��2c�3	qt�70������O��'��$	�6��]~�u&K`��j]��om�����DH��GI�}@�6�y\��5m[�3up�gVvp���w4�nӻEu�Kd�5�%p6�1h����\)��� F�e���I3�N5�'Kc�tl���'_'A�@�V�+{���;Aˉ���<�YSl,��u��ȕ�&��e�9�8:�Hv��g��{ƍ�6-X�����`&s��tEE�M�`x�oaPX6�ܝj�S���-D��l<�]��E��n9{����n����Ԯ�[�^I�@�Յ�&�W|�LNRU�$�H1� KJ�.k����QI)m.ѹ"��w��Ffǜ͊
��8���PE�L�,�g!ni�2�W�GY�Ç9���F�.2�����&���j��pȁ��_:�bF���q�k�ɭ��N:9�r���J�ۭ.E��C�,�p]�C�1�Z�Sb���*9zI�[��wn�I��d� �Y��/��kJ�2X�M5���nόUy�;���Ԅǫ��*��
t��jw,�����uM�,�u����i�܍C�{��IF��u��k�y)-��Qk�Z�\B��d|�-çn�ݛ�:p����L�f��E|$�>��9�>!N����j䳂�.�e[u,��9�}��Lܑ݊Y�ޭ$P� ��f	QR�[Q�pY[Keq�k1�(���K�\nK���A�S�U�V���UTS�Eb�e̃W+ba�*�c�j�R����ժ-k�\l̦*V(�R��m�ʱX�W.*�l�&0RƶᘥB��T9���J �eLfd��IBծ%������DF����q\��� �.\.+����q\lE�Q[n2�-��b�(���Lkn4�ZUJ6�����[Z��Ơ�U�5J��a��neR"��)n\SQQUV[KlUQe�sZђ*ꥪ�s*�D\�� ����&D[h�3.,��Y�U]!nU��ň��J���m�F(,-Z����S-DEF%��(�Qp��eq���Q1�F"�Q�[KZ(�j#�(0Cj&cH�䢪�h\�\�Z���P���e-F�~���L�-�>t� �f�)��B��d�Ժ�*t�ܼ�+o��.�E�ی��i�2��[9�cw]��5��B,�G�Pd�7v�d���7PSɈ]�+�&��Λ����/�C�+����`�Wj_�K��N��H&�c�p�Ry|���"���dO�zw�l/c�]Ҝ���e�H-y��(��:�8>;�]FpT�����X�^ZyG����R�xc4��wg��2�t��#��3��p���<��9LP,�w�r*�Fw�NG��h�����XQ�՞��x-L�����U�n�X5�E8f�����n��x��EiS{B��f��:����畇�s5r�I3;_�Ax��8�h9Z���Ñ�Ń�(��qL^\|�s{�,jm���lz,�7��0N
��+��b��6���u��g���.qR+̎���R����X)D�S;���s�G1c�ܤ��|x�m���P2�^�[J5���=*�Z0�ټ�C�����-�@�n7y�}&�Y��w.�%�m5�
)ǵ�ت���䣬Q�/��Z��s��(��C��`���{��.wWZEfZܷ*���:�yB=_d{C�A�JX�pN�ժV����G����[�;��αOd[�ר}}!���dJ�5Ԇ�t�wE�7{�}���ڏ%��)rVM��j���s��;�ʶ�����L@�����rLcO˂�=�7�NX����z�'7��~�_<��:��v���:��+�T�^ԂK˾\�y����{��%��-��=�ܞ9��ʧE�V��&��'tT~O-v{�[��I�6SܥV��-��b�����Mɻzǯ��WZ�V�J�J-1��\���c}�V��^��nLʻ�W�6���we�Y�3�[��8[����4�-H�u��e��fXcr;n�v ��)�d0�8�ԡ�8�R^Lf�9���S�2f����M�R��j���t��Y����P|9�7��"X����T����ۙu��:L�j��Fm.�eP�~M��Іd�˯g��G5�v�sy�sI�V�Iy��3{��{C��)=ff�g�m�e͛1#�Bgڣ��m�'dj�x��_{i��&�8��V9%�Ƶ̰�D�y�[���^�4���Q{ �^Юc�6�kQ��½|,E�|�B�/�hZ���g�ۤeP�&������=�P�Kw>�Q�����E�+oس�x��n=�)�]^�<���t�I��63��@��ڇz�ת��ι{x�GN鞩��CO% __WڽF�#Z8.Yq��V�oב���:�[c��ǥD-�7�]�V��V�f���N��f���Ke�B�ӃR��9ݩ0L����J���ި�Q��jl�2#� ���M.1ɹ��gZ��t�a&t�m�2v�ᖪ�\y�N�HȾmA�Z�sɆ,�������WL*}�ۦ��n�jBĒ����>�߽O�2� ��i^L�Iy�y#��-gQ�5��e5�<�#�9>�ߥ��}N�������W�b��܆��ۨZ�jJ�LgY]Y��=I�q��WA�.��	���>��jU;�%Z|�:�5�+�٤$����F�(;gZ/G�F�hʠm���INR�}�L���\2����9�&�<������d{<���nlh�q5[�)���8�kt�5��	�s�8CR��f�<=�ub�u��\�ycߚ�+�+����M<8N��֟s���}@��K�t,ꮝY�����O|�4�+��C,հ,��[�k���.)���n����c qjiD��gU�k(���m��iG~��Jʒ��Ei��9�v�v�t���`�r�߶$։v̾�ˮ�b�e=��QRq����H�������s�v??OTo��4EW�Wg�Uknъ����kcN�_���{�O�3~�k��E�s�b�=.�y9U����)�N�з(��'==>m�.�:[c<Y���[�\���0��\�s�CVׂ�7�y��[�x�(��>��YS��7�,d���dFMmA��V;��c2v͘��-�s�G��1:���U���ǆcV=NE�W�{
�Ny|���"��e:��3r����s��n@sC�=�XE�\829nQ��͙��+/w�Q��)i���=�P�ޝ�\-���6{ԥK�N�^�\�L/��;\5�r.���g�����w���~ԝm�XV�)�]���Y����wa�Y(�6�_h(&��1��%��+��ռe]B���*CE� ��Ï��i��g'Q��'��-F.��d�������Y�t7�,���y�|�X5��K�t]�������-��ַO_T��xg٢��fj��I�x]����M�~���}E���S4;'��/+���KE�8�1�3��v��M��m�}3�#�ܼ�\i����X���8��Ǣ���x����ѓ�?k<���ZǬD��[Mg��u�w��v�ώ"N�}��������_{}�p��	H�.����f��B��.�I�G���,Ӓ�XB/�9�#}&�����8j=��y53��ȷw�Tw"����/n����<�����yҤ���1��zevS���C9��tLB�~L3�����=��5��y@tSy�r�&`W�Xo��z�6�G�V;1k,=�Ѥ�b��U�7[�t���t���--�YN���Է����>3iS=�y\y��X�}t�+nH�;���g����&����Q���u�=^X�=%\�S���=r�,.���u��]ɾ�r?o�-�u`.w�탇H:
3�b�v����r��=�+���*��ܕ���F�{���Y�i�V^���<ܿ9���C�O�e�w2��EC�_����T��l����V��ȭ~K�Of.��Sޮ�yu,u�bF��z�H�[���V��Pu��QA��4kF��*�y��x�>��Wۆc��wI[Rem���c�hGْZ��ZV�U}6S�[�%���Sb���/�ʝ\��gM�厭�Gv����Y�]:�7���)��l�}Y(�� �Ϋo69��.� �;t��),���¸nU��Э�������Z�C�V���c���Kڵ�͖$�F��6�%�QO���sT��G,��6<��9���f�ケ�:�	[��xCwj�`|�FU.�j����S(�.ܘ���M[�i�j�f�t9NӴ�.k�����t�W����M9@5u�.U�)���߿������ǭ�ݯ߼L����\��W����lt_���dw���$8i�
��_�=��b��	X�ŧ��Ϣ��{�����5�#�$��D)2��⧻WZq�k��B��,U�\?W��Dxx �r���}c}���M�h+�㛯��3�C�O
���d"u!�h)(6����+��<{j�^D�;�c�{�i}�5\km�A�/������ Hhq����PxQ����<{y3��e�!��~�O.5�ZC<��?!X����K.���(i�zj�Vurݰ��\�m�3���e�r���X��|p�r�xIʮ�x.4��xȬ_ �C��������r ��Ws���:�E�j!���v|*R3�y�`~7�1�f�_�fY���p��(0w�־9��+��	BZ�X�ny�o��f�~�Rqwr\VH�u��wS����j2)
�W6��.U�·���3�tl��I��j�(�kM�RN�]��.�3��4�\7n�@�i���k�sv����L7�y}��U���U�*���C��uW�LM4���C�~���;���x����I�����j��W:9<4�r���dߵ��1V~�j5�v�:{�
��GO��H�3��l�+}B��P��C�\s�;�ot\o�܃���~�k\�x8x��?�٠^c���w�g���e��~�z��M��Y�O�T���c�w��Ƙ_o����Ǐ����u�x��.�|�zk��Y��"Cަx�j3>��]�%B����Η��,�f��\�|�_/��'��dW��Z7�
�wOxy��5��o\-�ί8�Q�4���o����2���uQ1�p����ٝ=�ٗg������{����A������6(� �}���6�7y�����ǧ��p���C���|p�t�g��Nϼr��;`y������z��ْ�����2^��(=��}hخ�/r�$��X�2����٣0�`D�	dd2�Mg)��nv��Hݨ���� �u�:�DH���%{�P���M)�,�J~r����#����P�(*�ЦygY�����=[1�8�ת�P~� ����_Q����M�\k׀�f�ۣif������Z�9j�R�[����1D	�wC�|D�|Yc�S\��{(vor�a��~�ubl_+!�p�P�r���͙oJ�(s��-6�%��g�}r��Cp�L-J��o�	V��O�����=Η�gS���r�doӪ���$q�Ca�xf{;w켭��_Q�!R�Y���(�u<֦dԭ���sP����9C�jR�>�}����P�J��Ɯ�O<����H��A^!P�i̚�;V5|״�������h���^�RU��n��q
r�pw͖H�����]n�!O��X�g�TU8����(�P7Z򫲃l��l����(��_�W���?�u�N�-V���R����/Vy|"y�Ii��7��R� �Ŀ�(fW��S6�����5�=���&��nBIbI ��HBPO�|��tP{��7T�}��������" O*�U�gI�sW�Lv���|s��~��k��q��WuB�(��g���:���e����x����1����D	�ɻ���}��E�����T��"����%TZK����xGM���C=2]O�u��/_���ռ��Ą@��G��7?oET6�/��������yf?��1���ܶW��8\��eǥ=��⪩�m���Ljܔ���bV�V�i{p��y�$�#�H���x�Jª�&�%�[-��B׿�x�<X�ۏ���B M�I�"��ӌ�s/����x�ҪoK;j8�ᄓ��c�w�0�����^�m�T�B N�SKJޜg�m��'���p���Wj�D���O>�]���;#�&��Ӵ�o㴜�z�}��7y�9�����ZU>����CK����%)ChI%��9���OzJtV>�NUb�t\a��m�=��ő81����"�d�z��J�/.�8�'
�$�T�1���Pt:fF#�Jc��Դ�����)R^L���T��֏nlᥣ�s�b��r�S��pt�Q�0���?b�\g.a�I�}{G׿�a�5tG��:$�'�w<߅�u}ʗ��V�D徼�̏��ѳH��"u90��*��9(�!'\�l{J�w��O�^m�h�I����xg&8Q������JQt�t[��\;{��F�z��xN_���M58��ɉ�:���:�?<U��^X�4�,��S�>}�E(�lz�?;	%�db�*EB"�%$���]������f}=|!u���NeFF�:��⬋I���i�l1M��I�}���k����ܑN$$&)>�