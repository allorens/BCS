BZh91AY&SY�OJS�_�py����������`���>��
�*� �   @  9�            P� h h   c�>�� Kzռ   {����q��c7u�R��v�l��ݲ��E{�qp�}Ʈ ajV�v3n�	Ѳ��wn]�����S�   |�;��-n�u��C�tnS�'a�mm�t0A��Yn#�K�{���@KR�lwn�7 �2���c��x�  ������Kmt���w6[]�u5pfkqO����{���`�Z�\� s+�we;��_5��   �}��3;�nf�9t�n�5a���O{���szɬ6;�鱥�Z�Ú�nv�i�   r��<Ͷ������ۺ���v��z����{O6�p1����Հ��r����� @ � 0 @A�            5O�b?R��	��  	��1%0��T��D`M �4��i��%6�M=%U	�M0 L   ��R���Q�      � �Bb !�OT̚�DM&�D�A�R��di��#FF!�2 '��|��QL*����|_ y�_���H$t��IH��"� ���-{���?������a����?����i=��?��H u��U-�`-�d����$�� ��+n�۽���j֭{�Vތ*��v?������o���9��,[R��)r�տc��TzL�o�zIk#�_$2ܤK�fH_\��+��5��Tpm��%c���o��˾�t��H��.y�����0�Y��㑭VK��r�"���}b�����$�Z�4���ؽ֙�ݧ�^H]�H���CB�ݩӖ�rp�FH�$�8/'w�,����d��Ym3t���U�1eԅ۔���q��(��K��89��.�$��ݟ1t�t��IT��b+���l��Uf_��F�d&�#N(�Q̓�\ w��.�'z9k�Ӯ�6��co��L�n�y!}r�=&q9�N��$WNZ����%e��8**N>��,���)�Ipv�m3q�x��u�D$ ��׾�H�Ӗ�rp�FIf8.�&��%�o��I���K�r�u!v�"\ML5�(��M���I0����b��7��^�p�B��h\�L�f�0��FkK�F�d4d.�QȤ2NpT_�<��N5ގb�6��~蟏�m
uH�E��|T4�t�xq��ٔ�/��ZE�t��B�7�7�7�Cqy<\X�!1_¿�L��O�1�gSxn�&/���v�E'��S|8��$D�lm3���R��	�;m����>�:�<7^�8u<L��5X���D�����5Hh��"�r�]�����p]*L-��Y�&pXzL<��K�r�u!v�"\��&R|G��	SMy��q�<���ȏ�Y�H����墮C��E�����s�CT���$Pr(d�:���<9�ޒw���M���#���3ꍡN��N.�>.�o1x���'�ZE�t��B�7�7�N�!���W7HLV��>������:&*���O���|�Ͻm����|8��hi�46��g����/s������ؚp�ᜄ���a��p�<��%`��$Ą<N#�3�	ߓU�^]�?'�R��$*bb�	��&*�q,�D"א.�+�pL^>�5H�h�X!y	�g�4||,E�<����e�K��%7K���]Y��dW�3֧8��g�T�V
g,���;�<Β{��穞�;i߼�.G2�S�3*N�_μ��ֈ�<�����I$1>ە$<�$�S��ޥ�.��me���[�N:M�tm�^�]��8��嬱>�Y]U�;��|�˾|��|�7-��'Ȳ4�]�?y{��e�G��&�X�֜���&8�����6chT4�k�7�i��y��_�����b���|�\:݉�ə^N�byx'O�wV�{����'�-0�&��.�Q�j,�;�	�po�q	����c�7]wn��]�Vq���ﳸ�����������G�'���`�$��9�L��U#�6�[�e��!��r���sԙ��J�%Ԓ�-6[%�<Βy����N�?Scc�����&:1���N�m�i�~l��#����3��v��V`�c�;���-ю�99�矧\���'���օ�أ#u�|��GDp�:�#f:�ݍ�$���r����hX�67o�ru���I����&��p���wq�؛G[��v9��G;ט��s1�G��coc�ϓ�Kq�O�n���r��}n�8��6��Z<����;������z�뗏���;��m��oט4������zC��=!ι<�xy�����M��֚����g_8�t~����?w�a�:zOs�I�qԹ=�I��8��1���hCBmW�k��6�6G����I;I��
���y��o�I���$��a$�$��q�ݕ rJ����6u�vꌧ28�w�r�����ד�N�o9�r����A{�h�ۣ��GMk�օ�>ӎ��,k�8>g���c�uWrU�p��8�������c;$G�t�>��O?[a&�u�d��U#�6��[1��fS�?zԮ�s��
�L�%Ԓ����lv��:H_� ~����u��|���F9�})��26����!��c.9^g�O��ܻw�v�n���}���g\���&9�]k���\��|��G^�e1���cn�ݒJ��+�q[�n�t��'��ɜ�q�[8���7��~o��&��:�ސ�uc�>�s�y�1��(���clo�1����%�SL��������㉱6�֏8�9�w���y�f:1í�s
p����[�v�yM`��<���s�$9�u�uט[�{�X���ߛ]i�sj4��:�y�w���9޳�E�{�w;'OI��o*Os�w���d�'\�օ�4!�6��]mco��|l�w����$�?���<�p�Ҥ�����'*H�FN�N���9"��9��ۻu|Vr���w됍O9�}~]j�s�U�\3�8��˜��Nw'4Mڽ-<<�Kh	�<i�fT�?'��zA����,�H�=
Y��vb�����\�/�a���R�PV���_�z���۳��7�w���=}���}q���r��B�x�UN\�7Q��>]:��JX�i�	�QS�-��Ҷ��B�}b�G�֊�h�
>�83M#m_�	��c!H&Ď�!ͺq��r�B���y�s��gcPю$E���(=��#�	2����G��n��C�:(��1^iE`9rcX�7(q�4KDCb+���KV$6Ʊv��i���=�J�,�R���h�LrL}4�͙�Jp�!F�6YE?h�!�|3�����|���:N�Zmf���;����:�N����	Ⱦ�k��It�2��n�!޳y
���P�AX�{ٲ����{I�Ւ�Rǎ�?�Q&-Bّ2D m�hC(�B<�Y`�iu�h�#�e��[2��f�o�-�)�E��	U$�,�f�w�5�-d>)���;�����HM	h� (�5w�i�#�ȱm��6���� F��7L�M|�j��
pJo���""�D?t۞��f�o����L������_�.y�q�^L�i�Ɗ؊UE�>�>E86���R�'�Z�r#}M��ĥe ���a~�T\f���=�vS���Kg`U��$*$F��=87�%��J����^o�Ͻ>���C!9��7Ny��,�����4�q&|<hgu�h�H\���J�L��>��Z�s�B �)O�=�1b��>8�%�ӥZnk�
F����Û-N����.�����ǟt�j���>~�s��m�>Y���9������PP���Q�����"6� �E�&���x����o�p��Xź�?���dA$�N��f�DDG���K�T��;r�e5��s���4A���K4dM�D�A"�#1�R"�n~�\i7�:A'������:m��u��8�L܆�frb�ý��f���R��ڊS�}.C��>vS�Q0eyE�F�"���ɪ�A2�~~�>ݣ���	'4�]�	waJ��4Y�C�����7�|ґo��[����MsG������8XQo,8F�K,��qҕ�����:w��A��eVA(2�3{wV�jL4xػ���I�R�uw�x���Ƹ����M۫q6�ȥB�īɒFB[(.֍>��B���4�~��Ço�x�w�ǯW�c�(�(22tD�|í$1|���b$��X�N7k�5q��?/B��0��B(֐�8A��)6�i�x�����`���VR��B������4KHT� �P��e!1���)'ד��s4V�)�5�!��~���Q��p!e��6Nґ�-X�ȓ���hkg�7p�"��!=R�a��5�ȟNYR�t��Y`�"DA(�(��d+ե�! "�(�Ȳ֜�iUpf�D(�R)F"�-����&�ш��b2c�]��iA`P���?sE�Z��$c�QD0%Dj��ꔆ���� �@A���r��_>��I#��5�� B �b���1�^�#��@�FpD/#u
Ě�U�d 2fS�4�3��1�QP��Jb)�Q��b4وH@!A�!F@q��US��Dh2p�4��A6iH�V�"��!��(���כ.8�SN�p��Aa|A�y�ƒU!�R�c(1(;K�
�c��h0��#�
����U����؞1��i���U Ka'�y�:pCΈd!��ˆ�a6�y�	� �A��JRca)�Ԣ�<B�r���\FR�ix���9�B`��Tn$P��M �4B"X��>�}��HAF#��!��R�m4��:�4����(����A;��ns�RW�j-��(�:���|�kL�ch���!LB8B=�����	[�~���|�:�S�WQf�)�J�Wb������T��'8"{��
�z����U���"�'1�Y�u��4\��
�Q�>�Q��n��+!Sʤ�p����I�m&鱯���l��*]������ۈ�Ҝ��4c9�����x>�Um�p��U�8��*E�g$��tj�2U�CZ+��ռ���Z#�ik,�d���Q�����I������J-z-�{}�ٳJC�a=���}�'����l)\GW��������ӃԞ/rQ���}P��k��"K��4ٍ&���k!kc���)ڻ5H�,�2F��v��e��Z�Znk��?�/����{W'9��z���7�����ع������T[�~���|������<��Ѿ���K���s�Ȣ���,Sy��n��/�}|_��6�qc_��.��t㛫���Nç}��ۺG!����ƝOS��5�m��cO�ϋ��˴ަy��g�y7gYr߷��ܾ��<�jHI	�]�Hݐ5�Ԑ �'��:V����T>ȁɌm�BLmĜ�wv��q�ۼ6���i]e��{�X���Y1�����sW��Z~��f�}h�J�Ts��^��NOx^��I�oulW^�3cP$p�M%9��c7ԫ��{�Q9w���
v�W�WlC�$����){_�ל���{���o��c+�hDGL����bIϔ��!4���B��$�D�	�&�(}���E4��}�۫&'��W	���i��YK"Q�>W�Rzs-C�Y���V%6�%#�=�۹lR�mZ���fO��{�/�23�.l�'��?����B$��wTpr8ě	��������q\�.�z�ƍO��2��+&����"��y�ۢ�6�[\"�BJQӴbN���_3�\��USlQ���|w�^A,n�B�)c_��]鸻��4>��t�F�I�-WMm=n5x-��9��^U#g�8��(�j!N/^4o��B
p��v�oN���L�4Q62�.���Q�d���H�aH;�o<��Ҹݭ��r�1�)DTB�=��r��]��|�7T5�k!j���{u�k5��a�\DM�Y%VF,x�SdPD�I�0�}�ۛgN��7���ӃvZ�"y)Z��^�h���b\v>h�Lm��m��C��N{��	s��ޥu�"M�$ې��BL����6�C���Ȣj�BU,T�*TJ^�o�q{]}"z�/��u!:�CCi�q|���/&�qMu뒩�AT�YitRj^�*�ުG�̲7���V���D�$Ity���M�I'7v������,�)vj(���r&�VqJ���?ؘ�#���=�Μ��n:�x�)
�T����JBJ�'�ʖ�KFG���V(Gk�7S�ʤ�';�s�,�$^
:�q�5d�t �"!F�I�ϭ��m��%�bY?k�z���Ib�|�q����~�Ԯ|���,�Q��A���Gx�gҩ�R��؇��Sڗ�|Y�	�&�6A����SlR�!�Ȕ�y�n�#���ʱ�ڙ-��%-���*h��H��\#湓�R��M'Q�8�b�r4�N��<Ռ��A�Lm�6!:H����Uƪ�b���YR�R��je�R�{!�jh�Ɖj#��of�y�y��5���ו��Rs�EJ����b�H�s[����@�>?+虜m�P��zBz��(���[�C������{�/W���	T���|��=���>?/0p�9�s�s��
 ,�������  ���8 @  0<*   Ѐ `�: ,�
 ,��@ {��%�/�|�_}8�PH  0 0������P`� �]�Q� �`� �  @ 0 �� � �( ��8 _|�K���$;�D<�������>�   B ������t( 뻺�    �(��� <  � @ � Ѐ ` s��4E�Q�ｖ�{����9�   � g�=�{��p((�wu`� <  �  �@�p 0 ��   ��  �  ���QBEA��[��_�>  �   {�����Ѐ ]��,`�   � : � � �l��8  �   �����À>� �8� �`��/{��� t]�P@�    � �( ,���
 ( �   �  3�6��}�)$$ �>�g���U�5�>��/��� ��a�>'���0{�y��h��\^B�ŋ���,^]B�����/!뷍�m��>b������]��f6a��,�!������M>|���ӷj���zzzc��HHBh]HT�+T�.�X��D*�>>>>|���ӳ�n���aZ�Z����h\M				
%�o���_���[Z�q�K�ꚺb�����1f��F����2 E��"����fR�\���k��t��i
��zW����G3�$Y�O�9�)ז\�P����3b7�F��C&̭�%��Uj)%�AȕY2l�'r2A�D5d��eY2ʋD�5���y1���d�# ŐB!"�-��d�!�(X2c �Rb�b)�4Q��2���FB@��#D3M#�C!��1���I�@eD�!d2�(�(�(QB(1��-�(��@��hBSr>�%CM%�&<�x��}��T���mBK^H6���o�g8���qn�V�;���4�ts���J�jQdb�M���)���X�ji^l�1!F��i�+n�N�[U���HB����ё��W�+�Ʃz�lNj��M�v<�N���\I��i�*�T��F�{ki%Q�$Mڐģ ��Hַ"�:�ܱ���m��LN�[fVG"��}��Ii�U�ʤ�V�*;��d�N��2z��nk��/{ߪ�M��Q������{�U������{��UU�%�Z���[�wvꪵ$��-^�nS�{��UUԾ�[��r�����뮼��۵Wl��f[���z��\�K�d�B;�bX�Kq
�I5��(��A�����SHd#�
!cP�����ݐ�i�F�I9"�2"U�5j�Kin$�#jD��lǂv�OP�Vb��$l�j7�rj�	���
���:0}x�=]�4>��-�x��3� �D�]!��gL�l3�L�x�
�#��`��k�t��f�j�,�zh�;<L}���Y;M'�6��.+�a�:�o�k�Β����t��郐�yY�aѾ���N�`("S쮕�»VyU�}�)_��١1x��c���1����韌�tn04ٺq�a\�Xt�l�U[�m,��WN�c�ٶa��խ���\VRH�8P��!!
n�U$�bLA��5eý�؊�W�UE�*萦2�h�j������Ix�(s��Æp:���$.����d,52�+m���1ٳl0�o-��u<�'3a���p���p+ʖ�b$���"!�RB&��R)*�-m�K�+
�sg�[(p�BU�a2�B��Ճe���Mi��874<��p#$��f�k!� �3���>����p�憸#�$�r��~�!��b��4N�p��3G���1<��ԆF�<w���m��v�*ŭÜ��Փ��#�[�M`��c@�U��7Z�mVԐ^�*i�H��Uƙmh#X!����R��i�F"�i�+L��ԝω��znV>F����3C�� ��ԌB��C��ܞ��h��;��b�-��y�zl{*ڪw!�֍���L�!g(�FN�	7�l��d����ٮ�_��Ƙ�:;6`��@@�w�L��b�Ss[��U���lNR�@�n�����8=<쵀��nBH�Sk?�#���,i�\�L��A+��$L�1 �i�����U
�UJ���B� �3��уp�FD��F��ދ�I��B2M�t7���x6%�]Ɍ4:zI&f��N�~2�G�,�̄ R�%
\�<btx����m�~b�4Y�ܶ����1nb�s;�;$��v&۸�>jŉ��HgV��<B�446�5-�fi��cJ��%a�}�J֡p����x�%#��i��B�}7���Q$#�G�Ѷ�#�i���l:&6HN�7�ؾ'����X��˖\nx|�:�e�Ş�m�M4�M�MۆFMl�s��;I��ɦ�G\*�d7��!p�AiG�pB�g`�Ǣ�c(�i���!&��O-�w���*�@�ށ(�4Xa>�B*LN�+HD�8 �\O���G:7&#��v2,�$Ɛ�DUch�bDiBI��cr0�1��::5<��]�Y$nkA�tv:���-a�F=���I*���T�P���HYj� A!P��HXhq��Î�C�c���!��!CC��0x�����P�L�h�Ӫ���������5+�ӻ���kY�&��SaT�f�Y�%ܧI��ƈB���Aєj䌬n�`ĒH4'/�3���D$��n:��֎A���Xsq�xV��gUzlxO9"a�`���	ӧߪ����s�=8�{"t�C����:za}�_M��;䎎�Bt�IЛ:0�Bt'H�G������=��v�Ne�4�^����^2���W.��.�NOr)�'$�tUq�1N��\b�1��g嫷�J��_�������'�\f׊��qgn3���\^�՝��r')r%Ȝ�'R�M�'keU�U�{W��.8�]�gǬt�/��ӌ|�_Vx�t�/�
�Ux�x��3�����'<�{��ꉟ�����.����M���R�� ��y����u������{c|�LX��o�l��Z�z�8�Սv��D�O$�O{���]�W~�����=ݛ�wU]KW�]NG��wnꫫV�q�ݛ�wU]�V���vn��Uj�ls^��n��Ugʒ�j�!P�w8� "dI�,Bi�ВիV�g���ƴ�j�'Dw,�7�鵒rRk�NKs��6j#��g��!��c3�V\e�����YTqp1�j7=�w$!$�β�3e���E��p8;�3��&¡@�"��`�Sr�88�^+���h0]\�0ln����`���l6����,�$~OLM؋��S4�%��ߚB���B&D�h�_d$�!%�V����'���m9�I��tT�)K7*a�c�uH��e8K��H#6Q����H쯋,�KZ�` �a���� ��[�����Pb��D�ma���+}ְ�&�zl6# �:�4Q����|�5�zM��zI��L�� ��J�`���ۣ��1��Z�;�Xv���M�d�T�&eF&�A��B���q&A�|K��i�%�����pp�A�4�iM8KH[�7 ƃaÌy4�H��-(�����dY�CS֛�H#Ao/U�i,K�n�)r7���CS�%�u�H��	ȧΈ��#�s�P_!��Ɗ�YmI51O]4*ݸ�T�cdw�BBBBBX�+F��=,��E�YD�p�ɒ:LL!cZ�3��d`�!�1���-��0�p����(p�*U8�s��aq������CQ�K��96H��I0����p�a��6�PFQ0Yp#2�ټ�7 �P�g��uNGu;XS8i�؀[��6H!�F(���2�G2ϖ�g���Tǜ�����X;e��g����T��E�׏�4�M(h~�	�����jfإJ�BKV�[���S��`�X��ʖ�#�������x4!�C���و_FJ���m:r99��24�"��8�A����A�
C0[﩯,�E��)����0�rZ��v�����f�}*��J��&��V$�+���;IC�b6�m�|`HBdppp>Y�Ϛi��tzqڰ��;�mWrիV�[$�z�h�K:M���r��!����Hb͔���"وXb�1CԁF���t���VC^�+����̖������l�1myʟ��oN�!x�L��خ�[�su6J;<sN&<�������¤ï������T��a�������^��J����,X����DdD�H\*hUj؟LLN�8�ۇiSݙ`�{P+U�i�aPצ�%�؈"I�#���"��uM�)�\ deƞ���w��T��s�F:e��|$f�Z�ݴ0��A���f�]�ܰ��y^g�:�X`0N��Ѻ��BF��9��C��Au��<�E�3��������!CC�0�U��$\�mթ��X*$�&5����R��߶s/'JTVu���>�vr1�	��&H�D$(HF$l,E�b�(>|��0듳�Mՙ����_S����F࣒�յ[�Q�d�R�x&��`��9"�d��"�whtYӚ01c��%���
��Y���{Ͷ��Y��.�N���ة�鉯���9wUA*�A�|FAz0kMA�`��:$��@��w��w�vĿ7ݠP1
(p1O���w�?��-�MB�i�pωV<�İ���'�X��ǩ�M'�L��;<z��M4ӣ��j�LT�ܬ�jM���������0����ǖm>LN�]��&�7��gJ�;��Ȧv�P�p�,50sq�a�@��c��,�C9�9�nA�cDA�J�A~?A�(HBXXmaP���FHFQC#�CL��;84-���v9l�#�2��rZ�ik4�:',��%�5�u��m��OR��91�2��imbt�Ӽ��'�ɳ����i���j�L!b���Z��YS�d�
C�{T�SE4f��$���qƂ��������`.6s#a�'*y9>�������c��Stf�[�����W�%�?���
Rc:U�3e����z�2��uErv�MK�����~��9*��42�HH9h��Q�әll6���끁���D�]�cӣ��j�LV���{dV���SM3X3��`��K0����F���AǍ�?%O�t�� �7w-os2$n��.K��ti��\�6<0ؤ�!�����ܶ�M�+Ī��D��L�VyS(�*b��o���J6�,-��j�l���ni%Gm�!C�����t��W�$!:����P<4�zv0fڪ.QP��:p{�/�	���Od��y���||:�/�����\Gޑ�0�!�#�����/�A���ƙ8�1x^-^��~k�׋���X����Ț'K��N��"�^��8���3����~b�З$�tI�r��w���ut�-YŪ��x�\^,�2q������t�x�+��x��+���[W1�ƙ�¸�x����y���x��'y.�[���i��1�.׋���4����q_/��v�6�/�
�j��x����sC~~�eտͣ���?G�f�v8Ȓ���D��dc�Sh��(�=P�J������L�*����.AW���ckH*?Cv���/��3|+P�З�)�� �l?�{b�t�)ĳF���=�ɽ7H
��Ē<����|Fh�>���ͅ#.c����-u�cE./�k�|Xq�N"�$X)I�z�vd��Q����,:m��"- �-~�F]�I����^/�[��mYi��2aD~E7�\��iz��8���
����[X4$�[��4C��!d`����f�Fz1��d4F�H,��-�����P�A����2�Ht٦�f�����>l ��8Ct��.";��p���	J<����4pԛ܇9���H�XS���׃ⲧ�)�a�q^8>��
�n�DM?�?��7��w�j��rL׌B�͟M�ZG���oW��gӻm�����k?�uV����^:�o����s�+rBIY9|���U���z3��G��g-������Rv5' ��-�^���osO�}��=�5���Y�[�"j�$Tډ�[/���TQ���qo9cl�2UV!���nE�bm:V[]�GD�r�Qm����m��G�kZ�EY4d�R�c�Sn�M&�o��V<�J'!�5pxƓ��I��YT*��I����yZL�����"�F�暂bKb��852n	���]����q>�����J��ݽ-秦q{ߧyڕ׻����ʫզ�)���ss2��i��{����f]ޭݒS����s2�V����?~�9��(i��c!C�ӂA�C&����(�1�B	+�N���HX)YJ$D8���D
Q�B��ZC �!	��*��C�ʖ*�Ԭ���Ԝ#$x�2娂�N�1�Wt0T����F"�!J"!�E�HƐ�!Ij�ŉ73*��춭]'GP�UL�g�%��6i6�,�{qFE�E<�NG�p0m|� 1o���T7l���ȹ񵃃E8C�K��~�9J��֠_� 84�0�
����`�d�C*��3��`����ɭ�U��E8W�_��)cRIR��mZVK�BW�l؈�h:< �,�XrTiI!$#%��0�M&2�/i��綊�ż9��u`��O��]���la��oO�u6t4S�~���٪,�)h�
C�7 wp��|h���Su �q�$�zg lh��:� �Df���v�%������SC<���,f���<vI�yP�fƆ�4x�1��O]�
�Lc�t�I&��d�Ş���Ch`Tt�j2�r2�]t�$�`S6�
D��*듓~��5Y��>4jTnfF9u�r<�x�R�#%����P����UԪ*��y# �m����o��W��B�OM�Gp5C��p���v�$�`�m�p�oe�p��D�1��npǗ(t��P�p����G�C��%6Q]��PC]Bx�cCl�G��	�û�&#wVTcLc�smV�w D�Qen��Bı�t����ͬ�,��l/���_�Ke��D�����Y$%�S�����@�R��c!CQ�<.�I^Y�\l-�%��r@t5�蘖�ɉ����H��x�N�S&�S1یctxv�L3�8��Cwg��E��kjQ3�.�tyS!Yi)'g{Hv>¶8>��a�QK��%:M�9�g0zEe D�ժnnl���*~�-���'�<��D��jA6?����l�	�܏"�j���,L�G&I�nL�j��6��AK"��*�Yb�18�Ŧx�f�sfj
�Æi(s�#�� �g��V�,q��T)�G��F���a��kc]�F��j��op�%S9-LOқ��X[��HJx�t�^�QTT��~C6��I���z2���P0�a�8J�,h��j� �-q!r�*�V�QI�Fd{5BU.e'Sҧ'��tj�1�ת��:=;v�+M1��f}�'��gI�Nt~����.2M�K������&�����u��ĩ��*m�4=X��j��!q�O%w�)p�;h��;�k��H�!DH�(��qiz������I;�3,??���c3+A��b�={��*ˉ�>J?�����b�ܛa�u���*�i���aZi��?'�s:�K�3���`�7C0r8!	
��*bT�u��q:��L'�hV
�P+
�\�F*D,R!T�;l� �&ڦ
�b*dt@�zh0<l-�lڶ�_ɣ�F�;Oq/��x7p���no��U��z��0����,"�*�ElC
P�WH%a16�.!�É���Wg��[iCC�0D �O�i$L2�x�XS�;M����'��t�a�Dfy �Ӓnd/����lǌJ�F�Y�j�ie�'�a�Q������P��v��Q����ô�;J<�iU+�u�jTƺ�%[�l�*sN�*���bu(�xz��R������My-�����i���V�t8!�}��։;1�A�3�6��ގ;d����dg;�JIRe,�9�w?w�F��
ɞӢ6M���K6�����b_�n	M>8��B|(��#?]�6a�S��Φ2�5*�h�ܫkiJv�=q8��fs�zG�ɩ��N�����S��1'�Q��t���0ܣ���ZLGi�'�ssG��%T�L):J���U[r�x�0A���.yѰ�h/7�?q��"hR�fZ0d�c��p�1#�|��)�=8�U�
�D?_ȶD>ȥ�%�Ĵ4S�Kj��I�Q������ż�Z�)0-��˪�&Mi�d땄�=ߪ�:��ˍ�6gX���HHXM���a�5(g�3�����#��{3J�sr��1��|f�ό�~�p�<
𰇐n�hhp=h����MP��h���D�y���'�Ƿ:�������'L�	��l�t����||t���>'O��>=��t|&���%��"����q{i��f�1�|��;^�gJ��y�s��\+������qX�~gˋūŕzU^I9;ĺ��'"{'$����U��Lq��g���������x�+��8�^./���̵W�9K���rI�\����^ ���W�z�z��ҿ/���\x�-^,��q_/׌v�9���NR��ȗ&�����o^��oI۝�!Q�:O�#��ߏ<�>�;}��t�?.w��������y�^|����� �LyOH�xO)p�B��j�%��㯼���e��3Ӟ��������]ڻ�w��9��s2�V�������eޭݒwwko��z�vI绻���̽[�$������f^�ױ����m�3/��V�4ծ*K��aX�9%#i���٣^a���r>Y� <�|���fHz�k5��btv������I��L��#NTL�F�QC�d��T�%5`�-Q���������T�����^�'��aR���O�=��pˁ�^�2�$�72D��[\6Y�Av��Z՟+���ڽ��S�Vݪ�i��۵aX�>y��]٫5���GS����Fң�r~:�4��~����L��h�eC������r�VYQV�����Sf|7#��z�6��T����0:�<
_��4<B��~�Ÿ�#�p��le�@ptpl��.xB!CC�0C�i���+�th�B�,�D%�M	�Kr�0��H!�"�l�v٢c�)E�	���je|���٦�)cYЈ����L��*�k�WJ�&S�	$GC�5�H�Ƹr�h6�G.KGkȓ�&E � ��"	��USR�Jn�d �2���
2��[U�A��[��-QS��[-v��OGؘr0�r�����h-�ޅ���w���i*h~J���hl�SSI�t>�nnY�lw?�1r�U���!C��!]<� y�GE���p�`�#��6�S%��6^� �gn���ꂄ��!���R�b�f���<� ������$�M�1ƨ�B��e|���9_R�kAf��F�Y��-����a/�U|�i=O]��&�Ə�C�X�"5R�AՉ4#��5䎇V�J"#��|W��F�>�N&���zsE���&�|z��:+�j�4xvڰ�WәYz3dd;O�'���M'㳴�=�i3GGs^v)SzG�~4��k�� 6�t���?�*�Y.ۗb2z�eC�����پ�ʲ��1:�����z�l��!UMRiz8��6v<�N�����g��|�8V�Uv���j±g6��3,��6EJu��kiN�c�ɤ��{����|UP,b�iJ�		*�BN�ep����=1:{��zx?y��&tv:?;�.<1:����~r�k�������z9r:���l�o��7� ���4C1��>�:$�-�8��B��8A���)�2W��!��{�	�_M�r��8Q��xMe��
��Q�HH�B�G|����մ� _<�GWf�}�qr߬����\�9�����iJ&ٔ��_�2^<l��! J�DĊ!(7W��GC���;#!��^���r��b��Ǻ����4�9�Jh����8��&�c���y�h��?[U�p�p4F|g�LO=v������g��
�v��U�Lghtd���8�Z��I�dk yhķ�pt:�xN2H[sR�88��<�Y�x<M'��{����gVcO�vө��㣕3uƵ�-+����,�x?<L�r���h�:�6;����Γ��+�:b�h����=y��+~��N�hD�^�ρ89|����H�I#�Á���1q�N�=�����@��/+���}�^c!�#��^"�I	�2�Z�kZ����|;�0;���q?|M�}����J�~߷��1)]�2�*hp�'��#�=|��1�G[V�1n��&�rڬ�(�@���*��r�A.���p��H�����@t)��>��0���6��Z�9o���%�l|m#!,ӱ��$!(���8��K��P�6���:k�����<g�������z`�����6Ώ����=���γ�ã�:`�xΏ����:K>�Ȥ�'��|�p��8>��\�4�ק�t�]+��1x^��j�x��8�^/2W�*���X��U_-Wk��W�U�j�-WK�m��j�^1�[8�q^�K��[��t�<:Y�4΍a:OE�dN�%ȜÑ9��%r]��ux�Ld��T1���c���|C�nO���`�!�ٌ�C�Y6z6u��<a�Ȝ��y�z�e�og��6	�I$Qd��u��;�lc�^V��<�D�̚�笠si�6�$�JZ�P��@h��%#d,�*���Q����`ɨ��i�[�Љd��'f����"��!�asD�aIi��Q	Ѩ�Pղ×sM��!T���:v}�&4&x����>��H��bV.��"ǎ"�����6�	����gth��Ѥ�����M�)�"�MXK��H� ��4eLtD��)
�1��r����N�2�"���!��A� �=4�F6��� �p���ʍ(�	�tctCH�BՐ�b��<��5�,�H��Z�w��8.r%�$�wlZI�c�� ���ʦH��]�]��۳Z�g>]�v��T�	c����/?l�=EH��tޮ���������5l�H+S_�!w׺4��yb޾�"��[#�e�Y�[&NZ�H����ƺè�G�9�{_�4�Ї���g+h�VV$���6*r�
�:-#�&=�N$48K�Wd�*�c*N;R1"8�MHn�K1����r���)���i�̉>
;	����J�,�A�7�ɶ8�9byc��ce�G��Ս��Q�<�WU�_�Om�3/V����wv�����u�~{��[}��պ�?=��۾�fj�{������35n���wwv�����+V��+\K�t��{{1��Z��Q
X�.B��"����W	&42����h"FR��H"FQы�"`�2�H�2�2�h�	]J�A��r��D% ܣ�rɑ���,v!	�H'rV�"Ya2�M��<�x0��HJREX�.�K�ce���hv;=67Aq�C�� ��+hW۫--�_$��ob��h�:N��m���ۉ��X�>����#����Y��v��o����`�pC^�!q�Je�;�c3񋒜OF�w���gM�c�G���
�yZ[z#ä�hzm)��WEF�!�y6l�M�6��,������A�_��YI\�g���2��J���<"�(��ċ�}oQՎ��^'��;OE���ˁ�O	/��r<��Κr8�
�j_%ti��1�����8��"��7�"�l�������8P�qk<�B��R��$3�m���,6��4�n�.�/-̮��!/�£�y��~�|p9�~����/F490v��<��z�	TSUQTl|�ɦo���� t8h���<�Z�O���c+��>�itz���<p:��zjob�@�C��4!ݥ5�nfGUF��Ȇ�%�׸�u��tΤ�7;�J�=�ܖU�
A�N���HHƜ��C��c�EP�YN�.;�Yp�r����v8�N��&���J�s$�{lWGIܛ�LS�m���1��IF_ܮ��8��h�zw��,��Id5�6�pC˻ɫh�Uf��D,!��FXP�%�1��Z*�j��B5cNƍ�kX���s�@�zD��Ll�d�'H!���B�|�V�b�o�{Q�FACf�`�yX�ݘ]hYEy�3Fv�^<.D�I�LN�!!�����ls�ӱ��߃u�����NC|�ԩ���vC��!�9��̙�xp�s����̦���oN'n���O����-i��+&2Y�=7?|�m)�~ܹQi��eA��
�!�8"&<4`�{�?m���sw)�] �;@�z`l�m�$%.���ʇ�6���a���a��[o?vv{�nyi]'�hͦ�ѩ�y�/���\��K��m���4SK1�fb1d�� Z�#g�T�U9`�t;
����><�p2>K0l0��J1�����Fx��2A�hy�[�^��0�,綠��e��B�:��7��g���Ce�C��<]V,��SZ�վ������ºV���_V�xI8�SRU�lﾻ���|\��b���S���*~�xF��}���z5�I�|�tق"|@�<6 ��D���$�J�T��.����m��I��-n%�(B`�������t4d���2�'M��l5z����c#�ӛ���u�F9'd����������o읟'l�<.�4{��z��ԯ\t�c�<;m�1�O=���X�h �OȈ�ljc��Ei,������i&"�3��%��1�6������J�Q�x��5Qo�Y[�x�O�*u:"5r�b�TQ"- ��Mc��I��_���1�O �@��*�c!�K"y3������G[X�BG*]�vь:�g�G!◷!�q�`���B�9�/����#����.BKQ-H}2�����^����hщSG���)c�W��+�=;m�1gsw匀lx���p��8�!�& �3�@�1CCaڻ���@�ߖ{?ˊr��K
E��=�W/{�b2-��p>���x0|x71�@�j�xu���>N�nYb�N�� ���\��Y:z>�q�=!�h��g�ӌ�8==gD��h�tp��:`�=g���M��vˊ�6�p�Z�/��L�\x���4ttN���DN�'Bt��>!�N�����h�"L%Cѓ��x�z��L�]I�%�~]�-�����'g���^+n2q|q�=c��1����Ý	ȗ"r'"r]���;����}UW������˵���m�'D���a<'	�xD�&�$��zD�K����׷����K��V������S�W�+���Qr���K՟���s�7����z5������
{'��MK�K���3:w}��[�����ݻ��f���u�����s3V�z��wwn﹙�u����ݻ��f��������s1Zi�X�k�O�a�E��}�v����C�Ѡ��A�Ȗ��A���M�������c,�V/�A�����m��+�ݣ�~U�g��d��0�é5?&'g:<v���ǗV�;N's�V��^;���_�y�R���ς�)�Æt&���Ѯ��J$j�ݻ��b�d$!����ݛ9Aq��x0�p��h���c�|���S�[VU��?g���ͥ��Jh�4�䩲��[|*tgf���r�U�j����a�w���>��	#q�i���:�Jw����#��q�%d��f�ޫ��8q��)U :@�BC ����jᰛ����������?��,^��;�B6xi�\�d��]׸ĚVF�fT�k�!�ՋDFi1��G��$5\c�!��Fx�x?���צS�P�ho�\�
gة��C��_���I�����k����G��?��$�AH�����~BĆz���k�O
zv�N���|d������&�N�*ve3��YѴ�[mU����l1�r����7;lΔ��`dp9�pɲ^ͧ�6a��tv�ϧ�M"A~?����P���D�N��#IJB�K���+��BI��wR�	�PK��&�r��m�&,����W��_>����Ͼ_�Tn9�Һq�LF{�g��>�� fY��Ϡ�p7���WUf��;��?Z�<Q(�!�؊;�.!"d�<^h46v6ǣۅ��0� �6�g�����9�"8�������y�y��l�ٴ�h�}ٍ��ҫ�cӵ+q�����A������
d�}�ږ�!2"7-����W��)������%\6s���<M~nk4պ�i[M��Ē�� 0���1�I�Ј<d̝�%�����s燃���iM'}��K;>Mvzly��1�o�O�i���Z�%2�$UD1J�Q* ��e	z2��cI(R&�Z��=2p]�T�܍�i��(�JD�1�B����L)G+�]e7^�a�,Y�][��g_J*���'%��B&���8��(����F�*^ �4�G��Q�(�!:ꎴ��K&!Z�Ŷ�jL��U���O��l����SÝ�����=,9?*ޏ�r7��!׹�w�C����C�����$��j�SQP�p��e�wIt�������ʄ$ԏ������x<;R�����4�&�ҭ��z�;M���i9IY|��U�$I���a��F��V��:N&�<LF�Si��}x��!~�-ȝ�R�˔h��S�<c�r�_��Y3�t���:N��ԧd�jT�V�Q�i���5QB�N<����v�Or�+FIN&&͡����&�P\�s�N0�RIN嶅�+����Aa<�DU�����|������K����e͛M��{*o��g��N��ӛO���=B��H(�aҲV�JѲ��W�gjV��<�5�U���7
>��w/g|��y�<�Z�Y�`�Oi���3%��s?e�93��NA9��b�w�d%�C�j����h�9�m�޸�6xx4��w\,���1q��n8��&�6�O�8u�����'�酗�d�g��l���'NOY��t�&Η�G	���O	��M��'F�:N�'	�Ǆ��:��yoN3���y��^-^�W��}"t�'I�W��a,��HLo7����'S��x���� �����^n�9y��g�zNKn1�x�W2���<^.��S��Iȗ"r]oY�Sv���I'�BzJ�Y��d����k���W��g����Ӛ���d��$��$��8d9�.����┨�l���l:�8N�-!��[��iJ20��%FS�jF��1��_ԗ[F���̲0��A#4R����D���2�s���ܱ�߫�)X�Y2�.q���ӆ�	��"5:�
�h��j��^�A"�r�c���+�؛��i���di��Ƕ�u�P6�+���b-���ǭxE���k����Sc�ʄ��S-dx��9,��V)�$P�=�lm�v��@w{S�D����g�A<h�mX�j�R�����D�D�D!��ˈD�(�@�� "HPb����F� ��p�A,�?F��"	,�x#��=��I#�%�e�2B2H0�S8[j���(�WPЩ�F6K�J6D\�,��97%��fԖ�4�ǭ��T�ys�o�-u�z��ґ�D��5�Z��ƚ#����e�wUH퐩��8�v1�:�Vu�9����i��KI�Z�άe�Ҫ�����|�cic�F�X�i.cv2�&�U����M%�kK��j����I�o����b5��q�IIu6�#�WG��5S��%�j�R��cȅD��&V����Zn3Dj!+tƈQ��o+�!Z�Ε��J٤~�kv"b5�U]�Y��_�����n���3V�{�wwv�﹚�[�{���w}�պ����ڪ��Z�[�{��UU���[�{��UUY��4�,M5��ڕ�oƾ��j�u-[X�(��'��
4�d �! �2���c)I�$tHX1"B�L�i6��Q*�Q*�J���\r�u:AD6��| �CDh�b�4)���i*�U�i0'ƶxu�z���&c,ٓ>J�4��Ѣn5�xT�m�t�9��08Xv�
�Ѹ\h`dp�,-1����`�s��V�A!f�o+���ڙk��A	�D�!"j���*bjvu:4�:8��V:Ux���J���i=O�����Ppt6��s��Xr��h8�%�	��܁Ҫ�Tp�*�ޭކ@��A�Y�Mg�yT֢l�G��kVd���%ĞR�1m�'S}~:jL9��4T�o���O�~�<Uc����jT��	��y�7a{���J�����C�n����d.�|[txg��}��Bs�x�HE����%�5m�e��^��F��J�}�J�@�7�av�Ҥ$Km�x8�ڽN�;O�u�14��V:Uz���J���kW���<�i��;K��|"5�&Ȋ!5l%J��lЌg+���	� r�H�xC �p�y��U��Xt�\&�q2M&�<�h�ܵo�:x��<1�1�~v<;R�s�̯ZF�!��	X��TX8������Yf��, �A2�R�|���b4X\]�A��Tm��j�w�n,�!�cI��7b�Q�S{�Syv���˔i�E"QQ���؆6F1���<F��J�;uY�]M3/����*v�t�7�|�~ӵ�Ə�SN���'m|�91�Un&�u<ݖ���8�v檳&2�؛O�:oϳG���ۍ18i:jI���Q��]��%��jۑ&��wP��#��pJk�HHg��[4~c�1�ޏԳ��Mh�,ZF�E����l���pkS�N*lѶT�:K�i׮��|S���{yY.Lf/ɤ�xT��4i^i_�6,D?
�mP�EI~e�J���X��CLbw�YXWJ�\�*Bu�$%͆Br4�m��#���٦=c����J���I�ѡ��Dd����Y���躚�K��jcs��s���m��ִޝ����j�ՓFE�8��0阕��zp�?$�=�{�˻��#O��<y�x��lI��zc�DY�4Ye;����N�5�������ރa����J�V����S�y;OO�6cc������ʁ ���
�"����m'G�|�YYs,�=G���䯃����ք5�D̵�E�wv�1j�%�4I1�GCա��A#���0ls�գ	!]�������ev�M��ʭæ�^�o������{BBd�#��c�1���NԮ�=�1d��"%ܣ���۸_>E:1�L���nI�jA���B�A�#&Z�!��&���%�?���y*��j�GmBM
�2*Q�%oP�U"B��*	�.2F)ҥ;ǉ��N���I��vZ�w�e�m�\Jt�x��u�e���󙕙r7:aڦ4�M�h�O�Ő����)���$�҈��7o.o(��x4BD��0x�����DN����j �!̍�݄��z4q*���Ak1���hCC:�gL��d�ɡ�w%(���qΈl:�o2Ht�͆�aǙ:D�D�J=7s�E�4h�ӆ��:qy���V�!bP��/!y��z��o�i�O���������n�p��,��```ed�x�ϟ>p������ҽ8p���ێ4㍺c��q���ϗ��4����>>>i���ۊ���N<q�y���ߗ��4�����>��|���=�DC���I���֝{�gE}�PG_��9q^O�^/<Rv��7}�w�(��峛��SX�'�WƠ��Q	Ѽ5�'h/jND7����kTW��"��QsNoZ�|t���W���E�u�߱o�ۯ�{�iUUY�V�{owwj��7V�{owwj��7V�u�wwj����n�n��UUf��n�n��UUgԭ6���6�v��J�e�'��zN�,��*y߮Z��ta�kU�D�>��K��WDj��fͳE�$���cI4�^e�?�!1�L��d3�S?
b���"BG&V�71����V�l���������A�ޫ����	:px:,�ki��1�x�<Uv�_f{SN8Pɏ)�IbYAL�����߮Ҕ�[��ۑ��Ԯ��Q�����&f>%N%���Kg�M���y�-��d�2��m6w���-I07ۮGCa��
[���s�Y�:�qj���U\c�1�=N�N�g��j8��K6�H��D8B�3g	ܦ��Y^�4u�&m
��n8�&Ѕ�Ӊ��Ga�qk)h�Q���%���7�6�]A�J��j��65R��u3�@���_6	,K�ENx2�gI�^�	��Һ�:��:N&'������v�;p,� h4�D��c��`��v{��+��UbQ}ؐ��\
�.jY$ɉ&��d��������[�9-�-�M'i�g�Y6{S����8�;Uv�u��\ɋul��*j�j׉�G���{��.�'B�+�xV�s�g���7�a��s�	ÂS������
%#%D��#�S/L��sh���B��|n0l]�*J��S�ܶ�xҫ�4�1���U��|:���=������:�n6n5ݎ��O��.���In�Y��UXI��q���<}�%<g�É�*|�v�뇼�5*�S㩤��Y�]�y<[_J����c��WjV��.e�s&�'{N���F��.�<:y{��X�24�3��~N�O�����T��S��S�Ogǅ*x~�Oq8il����tl�,:l��v70B(�C�L��p@�ߓ���BF�l���͹�[ed.|1��iI# ��K��-��2�$�c7����pf<�4�}8t�iSGD�ds͈ћ��P���#y�-[~y:��/\�\<���%�	E�Bu?����;:9+j9bRTYjKW�,4
�A�,oǈ�Q�Ȗ��y��!2����ǾR��C��������x]&���!rH]��!���y0~��/��:p&cw`�(�v��՚4[H(��E`{aY\+�xR$!�pDM���x@�ΥgoU��Hё��(`t���ޣ�GM�\%�������5A��F�� p`ݸX{i'"ڊJ!Ohj��T�a�dt��01�g�����7<�KmN&b��8�rcJ�1��o���a^{<�6OS���2	��j7��-+К򄨟w��4���c�8�:�S���!Q�k����awK ش��J�5��r����	!豏��5�d.����a󃑰h|x���s'~���X�lc�<UWl!��X}��~K!���\�HK��-��u��P7�8g~��/�CȋlN�Im��I�C? �|����.=��hh:=��������]`U�+��kcL��I'F&��6�5�V������&v�mT��6���ϛ|���<~|��+\T�B��!y�^B�V!-�m��>b�>>>>V�i��޼a�f�0����&,�|��j���Ҟ���\8||���*B��-Z�!b���8p���1����͸�8�-�8�|����4��_�>|C�{`��3Ծ��56Bh/<7-�ǰ5+Ki ���k99F|��vٓ��-QU^1̖�2�]6̠�Ɵ�,�i*{!�.>M��x4-��^be��KB̬6�&Z��z���Rƈ&|p[�6�GHi	-U�fUxǨ�cv��!�Ʉ5MC7��~�.��7q�3KU}r�;.T3�Ȅ��]��"�ۈ�r���l�ע4ҕ�h��X��D�B�B�!1R�(t���)���Z�4��G�I��c��B��b.YB} ��>źq	�$D4d���D�l��$�K*��K����#��GPӐGׄ�6N�o�Y����s�آq~g�G^���E�{���'�8Y�2~����式t[���5kx��֝r ��nb������z����u��'I�6bn5�e;"1oy8-�*��i(K1�8k&ǔ�S<�I|ؠ�����ڴ屡��qX�O�*�,-����n�a-#TT�+DYU�m��"�62$-�i(�����Zlc�D�q�j(i�D�2�ڣM��U�YJ�F�ZH�I\���u/��߾���ۋun�Z�wv�����[��ݪ������wwj��{�u�j��ڪ����o��w[m��2�c)���#��ǑBy��5��)!�Ebc�by
5�	ph!`4��A�B����" �R�an'F��hN �H��*��
�6(����W)TL!J$!.�[y'-��� �2�7.�����
�R�<���z41�	��
%�w�[a���B0��ߌ���գC���p>�wQ��a`݌��� ��$�bH9&2Q	5l�7�"�7d3�'s��'�n?Kb֣s�*���>zv���V�x̜5��sa��6�,CRTUT��������];���hr˗d�����j0��4��Uj�Ｔ�,K,�U[/���J�v��Ȥ.��e�ѬN�^'�i�l��Y�Q⪴�Lc;;Uv�?V]i��i6��d.�ǫ�BO�ͷ��-+P6W�9�d��b$$�������hɩvh�nO;OS��O�9�����M����Ż	0O�Ru����X��oO]��J�L�pI'�,����=�@��yX���YbA.Y$�d���3 x��3���;�}��"�Z�c��X�p=+�y\Bp���|˳c����N��2HH4:��c��E�C�<1�����pcw�M^�
ƿ'��<g�ɼ�?!��d�梊�1��b4��(�bҜ�s5:엶h悫�ă�Ad?��K��Ki���{H�2���	�d�e�D6*("!��+��]J"KD����G�H���t��(�HHI��Mbg,c7�/v0��������| �t<�G��kM��t�r��5)r�aT�gg]��x�'�ٌUz�lc�;+�a��v�K���Z����J�y~����A�	Dޱ<�֊)��Tr90Ė���AϚ�E)r�´��.7)E�[.�to�٭���=NI��?��$NBK?|`��A��g1�D0K����	�y>�^�N��ݬ����e�-�p���;�-J����Wc�����-�t4j0�z�EG����4�t;Ou������<FF�BW
��{��o�rt�2�o�67���%�w1=1>x����z���,���8=L�B,vtt;�2������.;YBԭ�����T��^�֪I	e^����^�����2�N	��GO�:&n�8��|[���f�Á��db�cM=$���7��PhT�Ӧ�r�U�ڠ��sc%X�s*!�Ҕ�J"��d�)�.5��U�a��7�hI4�B�+����b&Z��i�˖��"1H �&��oJi���U<N������m6l4W�`y$X"|�U�ʅzC�޻��av:�6�	;f2e�p4r�!/���yb�h�1D%�lD��L$�S:��2GD���<�$�OI��K��рtH-�Ga��z<g�U�e���'�io�'��yN�g��;�'����9�rѾ��,��i�u��1�L	a�X4��;ϛv��͸�ۇ�>z���i���X��!5�/!y�]X��
���4�������m6�۷��mZ|&	�a4Y�a��6����zzzc����;c�5�b���.�^]MZM				�vq������qǮ��o������0�V�0�ڕ⏭���~)���V�kw�I9�Ye4�>צ�|�|q#�p��wB	������ڕ�J��Q(��mW�ϓ���f�'=�.9{8/�=ۯ��~��5�գCj��{���ջ��UU���mj��ڪ���z��n��UUov=[Z�wv���|�����~����l(�Q�cN��+#4�x{V+�6SRB'�び�3�FBF�k�ŬU�$���u+P�*?���� dy��z �2<���cBV��׎�C��!U(��âB;BG�]��1�_��h���K���I��l�x�Ϧ2�WE �%P�
$˒��)�䭱��f.����pl-��#a��6�iod�m.�ʙ.��G;�I��<�h�Btvq��rz;vRyGвЖ"'���x �y��.|�{��1�t����iZV�� �h�!� l�͓vgx���DsO�1��e��B����+�g?��� K3��s;�n�5�2%E$���.$��qIB)d���r&�B� X�"�*���A��e���C���d�ac�ζ�	!�C���BgcN�]�7X�����3Q,��@c*S��,����Ӫn�J��x�U����8���Aﰂ�q�j��W���o����gG�<N'�S��,��xx^y'<�������`�d�20\�|���E���\*@��G��㒡�ca0>c��`����6��1�xzm��ͳ�V�l�m�d�T�j��<�px6t0�6�!��oܒHI$1��


, �M���w3B�{\:I�F�:�+��!6m1�s��o��G!�p�hp�mC��^��Ǉf�a�o.f^���s1eĄ� }��!�H�,B$���lZ�B�kC�t�z��&�O����q8�N'y-[���$B�-'�~ެT��<xHC^��S�&�i��V��c�ƌ0�&���e,4��L��p�˜Z˺mfn%�J�J�N>o5��E�y�^n#aF�!=�!��(��.�״�57�����Y� W�kp��Lyj��אT�e�U�a
�d�u�!��� �����BnF6��%ޙ�L�{B��$c \^,�w�n�v6���P�l;�����K�����}sZ����K����?fV+ϰ՚$��[wv0��Z+��i�w�����V��v�U�4�1�80`��w�����f���>ē!/4ݐ��f�;Z]�j�,x�ǖ�Klʨژ�HO�a+4���eϑ��4b�I(HX�Y42��H�Hm�P
�����{�/��.�QEF1��F�-M���2j�dx�G����o�FI���z>LV��g���,PbLaCXÆ?H]3L�Qp��Ň��a`��n�-�=�1U�1�p��1�y�Ug��٠hn����hn9&�Kc�űj�q�Mf�J����$xӼ��a�X-�:�`�z846��a�e���PAېla�ڹ�^��ogӪ����E�4|0�m��ө|���w|����|�����mbF;"*���	[M��s�FJ�Ʀ�v��UVR�o��"�R,���"�H�)�"Ȕ�B��,5I0J���)
���%I),"��F
B�"�%�#P��QRJ*IE��ȔXY$�X&$���QRJ,
*IE�QRJ*E(�TQ�FH�T��$�T��B��Qd���QHQRJ1HĒ�$�RTYY�$��Qd�D���
)
(�Y$����E�QbJ)e#"(�B��Q`QRJ*IE�EAEI(��f��@���TT��eM���T֕-���cU#J*%$��E�EI(�(�QRJ)4�����ML]�Z_0t�h�E$���ȔPQI(�EJ(QP��IE�J,QB�XJ,%"��I,%��#�)6Ҧ�T�T�T֕5��)%������X�Y$��QI(�Q`���
,IR�T�J((�QP��E��YT(�RJ)Y"�$QP��QQ)%�$Qd(�TJ(�TJ,IEH��RJ%$��QI(��T�*%T�,E$�QRJ(�T��%�%$����I*E��%TJ,%RJ,�Qu�#���Q(�TY$��QH��EB�Y0�+)�R�(T�i
�KEJ*P��L`e�JU�V�YeR�K	�R�h�*B�*))AJ�J%�R��*Q)E(�!e
�,�R�(w���hT�d�T�)B�,�R��R��VYX�Z�+�T�JV̩eL�eJV�ʊ�TVYU,�eL�el�)eJT����(ZJPR��)EJ)a�$bQJ*QJIR��(���(��J�T�l��)JX)AR�QJ)IR�R��������E(�E)%(�J��E(�I)EJ)EJ)AR�R�R�QR��),�eJV�*R�Rʔ�J�J�%)e,�,�JYe*�)JR��Z�R�RY)JU�R���R�Ҕ��R�(%*��JR�D�``���0JE��TJED�R)H�Y%IARTJE�(��)$�TJE�R*IH��Y%"Ĕ��H��0��d��d)�P�Y%"�)J��B"v7���>b��zҔ�Z������$$QU1T�$G>B�S��
�ɟ�7�g>~D���C���ǹ���y�o����쫊 '���}?<w�������9�}�k#JK�����2cЇ��M�iTzm��7���G�s���xY�~��}Qꊪ������^~P?/� �t/�!�� �t���0AG��� J�_�'�~�s�?�?7�!���A��%.���\ ��e=�O_��������������UQ'�J�̏��x��@L����S��N�<�u�,���Z_���RR�o��i�k��]GާG����s�K���~�S��ݧ�j���E(X�A}�@E�ؔ  �D@�"���CM?r�p��O�(�����M����Wv�����ѿ�Q����(��KEP�Z*��P�I�,���h�� Z��h�DK���&���Q>o��Jq����`���� &ߙr^���O����^��/��HC�Q'���ci����EUD�|��!`=_�ݭ��� ��C�~1��^���>^������� ���Oئ�'�}#�����}��ߢ~cG��~�UTK{W���2����~o��'8��������D@�>/�
���|�V+�q���������9C�ҽ�t���������6.����P�Z�Iy���$���G�K>�QAF� 1,��'�l��p%��ͤ��e%�4�����D��P�z�w�>�6$Վ�����M��o�}J��<@
P����I������>z/�U����X�i��	����'�?��'�~���������`��}%|V �����>����i~�}_gF~p~���IG�G���h���tn����)_�z��	>��[@���W�~��H�ȑb�TQ�Ɗ1�E�F4Q�b��h�(Ɗ1�E��h�1��1ch�4Q�(Ɗ1��cE�F4Q�cEѢ�lQ�Q�F4QE(Ɗ1��h�(Ɗ1��h�(ƌQ�b�1��lc(Ɗ(��h�cE�F4Q��1�DcE�F,QF6(ƍ�lQ�1�cE�F,Q�cE�F,QF4Q�cE��4QEh��Eh�hŌQE��4Q�cE�F4Q��1(��EQ�4hѣh�Eh�Q�4b��chъ4b��F(�E1F�Q�h�(ъ4cE�Q���"��c�F4QEcE�E�cE�F4Q�1�1���F4Q(�"��F4Q�cE�F4h�h�(ŌE�Q�b���F�Q�F�Q��F(ъ4b��(ъ4b�(ъ4b��Ɗ4b�F�Qc,b�Q��1b�h���1�,QF1b�Q�1��F1�F#F1#��Q��b1�4QF�1�c,XŊ*4bŊ�lTQFƋcb��Z*(�Ɗ��+,QcEF���bţF�����hѣ(�4h�F�ъ��F4X�bō1�,j,hŋ1�E�Q�h�F64TQE�Xب��61�QE4XѢ���4X��(�QEQF�1F�(��(آ�b�(��QEb�Q�(��(�QEh�EQ�1�(�F�(�EcQE1EQ�Q��(�(��(�Q�(���4QEQEh�(��b�1�cE�(�4h�EQE(�4h��4QE�F�(�4h�hѣE�(��1�F�(��(�EcF�(�QE4h��,Q�(Ѣ�,TcF,h�bƌX�hƋьcE�1���(�F�ب���cb��X�cF��EXьcEQEQF(�h��(�QE�Q�EQE�F�(��(���b�(Ѣ�(�E�Q�E��(�(��(�QE�(���4F(��(���4QEQEQE(�1�c�b�Q�F�1EQE��F�(��(��(ѣE�F��1F�4h��QF1h�EQEQ��F�Q�Eh���4QF(��,lX���F.V�o��}.�~D�
 '��c���T���������[�8�}� �H��B�C���7/$o.��"�x?cj� �Œ/�}\S��?U|��C���)�E�lu�;�L��e?��C8�J$`�����R�[�����������'����HD��o�͙ �:��*��6;�O�C�{}��PP�OX�a!�� ~�~�S��lPPr|�]*nW�K���f�O���q��I��7�H}�T!���O=S��rE8P��OJ