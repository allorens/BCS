BZh91AY&SYm�U�uߔpyc����߰����  a��                p  P����P�   
  QA@	�T��T�$@��� t1 |���!%
��� <�W{W[������������t�r��w)v[F&���gb��}�t�002KL�T�A!��4� d��2U٢C���E����<�8�����A�N��Zj���(Im^����]�g��.�:i5��t��m��Z�%A+F�Ѻ2eV��7feL�F �J��I�D�Җ�u�ޫ��^�{��B���sM�������.��ޕ��cu���8�w�m퓬�j��:�  �iPy�^�]�l��F=;�/f���A'f,z�Ald-AGn�Kc��Z���
���wG<�t흦��j� �  �Y���oN���i��`-/f�Trd��9�i� r�L�K-L��C�RA�ӱ�1ׯz��;֐�K��嘢 �(�   �ʤT��klDR���  � i� *���*P=C�4 0A�@2d� ��DIULD 0�# F m5J��R  h      	4�4jT����CLCF��&@b�)I  	�&�I�<��ѧ�i���M@	J�Fh��&#@�����y�O�B�bJ�Jɭ\r[$�2n��Y�y|ܜz�K�)L��n?��$�p�DN�J�z_���3Zi��;o��/]�S[~���^�7k_�q�ه�ˑ�e��_���%)bl���������f��r�)o	���$2
�����d.T!q����י�o���{s�];������S5>�ܣ���n�	��,���gDN8U4Q�J(J�SDgM��
�v�DN�p���J���0եA8P�#Ҩ�<�ob���_a�\�GR"pg
؉�u�x��<x�5~���~zU&�F��#r	�0�ϞԮH�gG�Bhn�"l~D�0�ғ���m��j��l7���oU��G����f��ڨ�ʉ�jtM���}jYΥ'9SF,�eQ����p�]j|�|�UL�HrD��Kv��=ʛ�Y�%'M�BB��J�N��:!���e�>�e��Vp�5;�)�FΛ6l�9�ģ�I�9ML��uh�4&�ԳGMt�@�M��GbQ-��>��GITsf�c�F�(A�QBd�L4&p���Q�F50L%5/�S�p�Z� �T�7Q(A��L!�v�tÇK�TD��l���}Z$AUD��N���jv�h�r�%��	'M�MO��TDs���:6H�tGXW4Ib&�╆��DD���飆�O� �97QG2�p�;�+�f5Κ�j}f�B�D؍�D�Z��RΔ;�tFH��)4C�$D؏�Ҹ#�����$�jh�����m��"5ʚ�bX�Re�����7q3�P����󫨘7,���D�8l~�({����啲�~~��M�m)6��keBQp�<��K��O����<��DL1J�a�[J�ĳD9iV�'�ӏ�!o���2�A!�n�}B3�ڈ��%�
'))4'ND�G�,�!�,�jpD�'��/���J�250��%"gZ���bP�n�&��L:�;pNT١!4��(J'R�5YR�'fH���@���$�J!�t�~�O�GuS�Ŝ(�ژ#��q�,�ڟpdÃ��M�D�l��Hoqcs���%��'��";�FUDٱ�8#����˩�	7ȉ�Ȗhwu(r|�hMH�ݔ��n�&��Ա��Q �Ѷ}F�&� ��TD����N	u:pG��Y�ԣ��J83�0Dy8"v�S��|�!æ�bib.����lO���"�Å��UBw2UYڝ����"hYg	��a�,y$��>I�ܤG�L0�e&Κ����WJ4;���JL�.h�	gGZ��.W��0�'M�D�;��D�ܬǙ+d�WJ4&�+��I��)bd��pMD�JL8p�$�,�:�%�}>��[�0�r��¶&�'�.U���l���cr�$(dHt�R��LJ颷'ȑ�H�gJ-�DM��W�hI>��L�BpD�r��F�+�t��%|�}�U	�4�Rsb%��2��E�]8&��W�?,��4&�JD�/�B#0��F�UT�O,�ɂt��}�Z��J��v�ȉ�ܪ�e=��%,��6t��N���RX�rR&��`�7�\���w����N��KL6h�wSF�u(�r'�'����D�͵I���e������"X�UF}E������Ue�ІnYF}e�ꪵ;Ȉ�lM2a ���ڣ�-V���S�i�Uni4'\�����"�V��=�Q�:h��%	DwU�9(�2��}p�"B:����~�U��}�0�#;+� �F���SB<��8V۪�&ܪᲲ�pGSbpMj��X��Vt�$��h���n�&Qu+��]���r�:n�Vh{:&,��E���/Q��S$��Ju*�JȔ[��D�{)8?"9�Vs�B;��t�4c�_"G��hN5)bggDa>~�v@К4�i"hM��-Ԥyo*��8nJ:$w)6�R"9&�$wuI�9�Wm���}F��&��u\��U��*�F�"&�T�0��ӆ�٢�wK*�MT��R=�vW����7�JN���.�m���Ԫ+����VY��N��	����&ı�U&6py�4&��W�sIPPA|��m�`�K'J�Dæܕ�6Yߓ��J�� �B�n�'0F��L} �67��蘝4h����9��M�؃s�/Q1��(ѳR&�{ډ�8.T�	�"Y�jY�a������&�		�8Ԥ��J���~�gk�'L(��l�m�N�WI۪�ʣ\�'n%��W~��t���V���������Q�f��l�W�؛6�WS�۔�4��UU$�ڪ(؛6�V�'9U�(Y�!Se5�J�UhJwU�:,�F�M��&���;�W���#�b<ʬ��y)4s�6Cr�|��RP�J���S8B�䢹4g'����j��"7	��UX���P�����TP�URY�/��$N���U&�UA.M��w:P����{���[4?�u+��%&����Z�".�|��,N�Dy%|�IR�#���H�l�_;���D�e5,����	�",�Fߢ!n�hN�_P���ԤN�)Ϧ�(����JD�I�c�_X�9��'J��YF��n �W)(J�WM�6��f\�nV�8b��6/������ �IBP���8A5�J��Y���މB50E�P������b%}b%�Џ"#q�L8%r"9KU�u!�}e�X����vN�ѭ�,��'�;�Уdu)(Jw)6Y����I�d�u�Ћ$ϻ�M�M	�����'DM�r�'2�N`�I�	�r�D�9˓�8�2lL'M�k�N$4we���͌�tj��pѤ�\
xNB[R&�8Q��>�2l��Eh����jh����6���ٳ�l�M��NJ�F�N"h�E����y0�gd�$A��]�g�ʝ5�ErD숓���B��I5�� ����
e�/�C�TG�Rd���?���aδ�\�����E\�G���߿��ֽ��V�2�_�穃�4l5�/�`n&|Qӽ��`��8����ܵ���5c��&#�=)�^����ߖt������1%�)4e9����<��_fb;[�~o����1W�OD5��'�������}�8�Ȍɴ���f�ە��wm�龔C!��X�/.�A��{��H��3�/I���ƾ?�:���%a�O�}{�݆����KWr�Y�=�N��wf}9�/:P��&>4p�{TE��b"/���s���u
��ǳ(�ҽ�+��������n����H=:f3`*�Ǧ.�t��(E�N�5��B.�=-~w:����T.����~'5�	m���?5ǵwz��v�5��w�ǐ?;^�Ʋ��{��k�{��Y�z����i�a�י 9}B2��)�g�v�ݯ�V�p�l7ھ�%��f����YT�1�I��ڟ}�U��e����!��w=oNޮ�5/��ܟmϚ}#���^|2�"O�b^!L�_��g�/h��:_�����\/�uϵ��A����z�1,F����4mzFG��W�OY��n��?�OY{zC�O1~�����t<>�����Je3)��^�B��/�;�_Y�ꮎ��2s9z͝���XVU�ɫ��ݙ��ϳ�ڲV1v�������t��/��c�.4I	66�6��}@�&����O�2�@�zo�|g|=w��g���اw��:{�y
�u����oY�����]�s�����n���+R���5Ye���9˹���ۛΞ����ɧ<��s:���_.�u��H^O;��<����P��1n���>x�������wY��;��c�>$�{����5so�S�F����w<f��$������~����8�տ��. �M�'��w���	�x����;�C����͐��л:�81S�T���xYY5�P-(��G�{��Nź>Cw3n�fÝ�o
������
p֋�k�Z~�|�y��%H��^ώ�y�^����l����<�/>(��P6���4���{���hݾ���x�gG竺&g�=ˊ|X�	���ǵ�ރ7ɇ�u��k'�u�����t����k?5ɛu[H{�W5��^��ɭ���?}��}����y��ه�v��wYp]�L���gz��:�V����fe�����L>��Რ����~}�����%>a�?gi":\�4�Holc�x2t$�A���v�@qa��'ݲт���Og�z�o,렐�ݚ��b����'��Tv�s�FN�;��^�m���2��������B�<i�wL��B]�,��tovɮ�J�����:�=\�޽$4<^�߷�WUǳ8)���E_Si��a���W��<F:�KuB�x	�צB�{��!WOQ�֣2F����q���[mVw%Zʕ����{u��UY��sb����������ɍ�l��lj9��	(��k�֨E���=�=�Nyc0����Vp�����\Ɗ��꯺n�N|�d�w%=-�Y;w2V���d��N��3����t�A�Fn�	�8��Ӂ�������NֻWj7����Q�����X��"��מ��m���l���#��=�vF)!vWkmsP�����W7�8N���C��ك�����G�m��_�6o���)�ž̝��^��~��i׽2C/���ޫ�_h��⁙WIa1����C�����k�3���n��C➸d�\Ѹ�~�wUא��834[[J�zȏ�vXzj���k���Œ�J+\+NW^�\�[(���yI�Λ��_w�X���|t"C��<Xe)�s�ې"1�b�J;��IC��֎�Y�F�.����I&�0�ͺQ9�ҌǎNQ��*D����xIF��}u�gJB'�7.W}g��o'�'t�iY����ˎ5[6oP�	��Z�u�$~:�v�q�=�Hz]��:acDz��ܺ�,;��ͮ<z�d?_g�^�Eu������$Fy�od������P�S�P���iP�3gD����L>��}���x��`�E��־���E�8�p�(�k���a��.��L�3gQ-�`S=�D��'v6z�Ο_��s�sن�;۰t����O�LZ��.L�����z3z01�C뱜�R��ێ2c�/�&�����3��������7׮:qF�9~��N��y���97�s�~�Kf�zG����ׯ�u�x�zv�2jx��;ܘEc���՛Q�U�K?l,L��7�YӐ�ܺfOv���^wO�{o�Q�y�=���s�Y�)|,�7�g�#x��ӧ���aoN�<}}�]��e��f)�=�i����Y�֏W_��C����]m��p��XQ�Bu��$�~��w����؈13��7�ݻT�_����M���:t��]���Z~8}�&y��Ň&�Ƴ �T}��▗���,����
%I��1�����4²\���3Iˇ(��9�9ㄔJ��)���	.Z*�1�ɥ�c}o1�'�ڙb�x�(��X_L����y�6Igt�����0�O�>u�\&�����Ѯo�$�o��}~2S��r��/ɑ�~~�a��N_������m�4z����t��ڬ߯\xK��+���u���}3r�I篺�0װ[P�`�L�gӫ̡�c��t)����<$���I�Ub�&DS����}h����~:d���z`w�}�Ldo��;݇xv��o#O9.v_J�o���;�{ �$jo�3�C�y�0�c��_X���;N�{cQ��xp�'Н�N5 �%x��O�:;��I]���E@o�;s����i�A�Ӷ��ni|����{��o	�(�:W�/H]���=܏׺���w;*���}u�Zu��5�C��wiï�ܐjԀ��uç({0��L��VƲo��>+NK�	����m�e�c}=7��+�9�\G���A��I�]�2un��}��vy�+���z隩����.T����Ó�Oz�������$�'^��D�s��I�WzVt�KO�/�iP��hV��w|��p��u���u����ms�mҏf�����5z��{�s�xq鮧I�,����>g��:s��Sy�\f�R.��fV��vTd�Ș�57��/�9��s��Gg=&�.v=���~��=��^�~X׹�m�;:���8�^���ǿt�[�����fl�1��]�&�&�]�~��ٟ{�(�4���I�as	�U��iIkՔ[�M�����6�l,6j��/�����F$%����nƙsv�3.�5Е�q�:\Jm\[��	%"�f�a6�L�ID���l3K��U��}���l
�ʋ$��>F݈�Ũ"R��e���\��m�'��q��=+.�ֱp:tBt-�2z�1�'�y� �w��K��nB�l��m1�r���5�0�d�[�F�%�0XFC,�$-%�6!H�� M ��4	�\�b�Sj�J�63��S˞:n ^֤���	f��إNi�i3
�m���Q�`�J�u3L\����H&���$r�P�l6í�����+�|B��7���"$t�P~.!6�8�o6�\b��*h(ԀM��7��f��Ll�2�ʺز�e7d|c��+S�28�T�*\{V��m����Y�E�><5_�
��C ��r� ȉ��O0����Q���j��pH=��$h��цP�!teC�CA�M�ᢀ���F�D��z���3 �o#
HB7d��6���}%�ڰxe�V����3L4��">40BQDI�9
mr50�H�`���F �l���n����W��;�7�^�c��vBc_��C�a�Y`�f)���$I�(�0$��!���%��F�%��nR�אR4�lBQ@�>rD���$6!��H7����CG����xBju��! �p�̂d@���-�9�`r@�l�$��;�L�� i ��a�I��0�4�	d���	�8)kc�S�$�����g������H˲K�X�Vf����0�����"M��yJD�)*����o�����*�@�.11���TF�\E!�}h3�Sg��6�$Bi�lp��;ʊ0�q�Z��FSvC�Ȃ��,�7"B�P����a�լ�:n�J����W�g�@�'�4��^(А��LJ�Ě'���K��.f�Of��A�Ť��#d7���Ҹ~��O
��4�8x8�agO3T9�KeOY�b.ٌ��OR�-�H=Q:n��#�<� �����m��&�����|g�n�2��	��|�W��!�FCH�ɛ6f�7��S��g����3ënA���uf6�o�:��<;��i����s4�?o�u���w/c(fP^F*�|�{�?S��LUW��WJ��iU[X�*�*���UW��{�����]*�U�Umb��V+�z��]��Uv��ZUV����������>6�m�"���*��t��Uڮ�W�Ҫ��UW�*��{��z��W��Uv��WJ��UU��Uz��U�U��v��u�����|�I��� �^�k�Ҫ����1UV֕W��Uv��WJ��]*ݗ�����U[ZUU��U�եUmUUUmiUx���|}�}��*�,��E!ѯ{�������}��^,V֗UUQUV֕W��U^*�U^�w.視�UWUU�*��t��U��U\X�����kK���O�$>	��2�$f%fP�-`5�d��_gr�JXf1��,fo�������Hrx;�Ž�������sr�0K�pN	g�ᣆ�� ��J:&�"'��ba�l� ��Ć	bY� ���
4"	��"%�(�4A�D�b'6"a����%	DA6�!�D�Q���B"hDLI�(�"%	����8"u&�L0D�%���	�X�'KF�:hND�"lD��N�����"Ce	F�#�N��νUXJs���ej��g�H���Rƚm3
=�h�6/=�XiQ+��l5�\;g�6��Jq2�e.�S��A�(�ʅ�Q��&��,�l#�q�h0�(�"P�5�R��(ą��6[��tE+#fU���")l�$����!AY�a��#� -�����5ի�n
����Y`��]c-㕋�
aЌ����a͵^!a@����4c����#�,���zx����#�Ɍ�5)v�/��k�脴�M3h��0LӴV%�BͶ.�Ԯf*Dn�G	(�.ŦI��>�=���ۓ�!�ĝ(�(MFDd d�#MRB�#Ym*�M�c6�1���&j�����K]krSV�a	�b�1u�Q�5�l��k�U�L�88�*+���v-��뛑�8��"D(���A%I�Y (�0�h�!0C�Al�\�� ���d����I�K	��b�.�\T40�� &�QFa&F["C	��S%ٸ�M��]J.kL�e��YZݝ��nV3���h��Bi����,6���Ά�,8H���Ȝ'�&��
 ��Ɔ|4f�a�j��D�`��Ѕ�-�eVh�F��&q1oa�1��}}�,6���!4����F��JL��"&`�!��
aؐ��H0�����H��:<l�J�:���`Z�+Wk��y�b�lE�ʀk�hM���Iu"R�emuq��K�A
0���g��I�$#0�H�=3`��.[ck��N��Z�*	%�\I��i�e�����AP��2'�$�`A�TƄ((E'ƒ�(B�d�P��
�īen���]M��5��XY�����d�Ktٵ������Ml66�UHʮ�%��B&���]s�q�Z"f��61�|��Qmm���,]�l�Ia+LT6�r����^�"!�oTk����-��)�I�Лk��T6�{��Q~�z������z���T
���{����s���`Iw��{���9�}פ$��{�������}��*�f^y��y��tL,�4&�0�tM��[�~���47���!Z�X�H!e
���].CY�e�n� ���\��o[�؅�%z6�Y(,Δ-%;`�5���J7�ó�C�����tu�5Ki�l�!a.h��q�;Ƅ�m=v���R��E�4�\�kt��L��J�e�`ᚚmH�[���{RP cJhSf�jʕ!6%B�L�51�d�@� @�נ�-Z℀��ci�(�"�F�(��כÙ��"�?�7�U�l=�xQ�MC���C�j)�����*"ڌ��0�4`w�eQ��=����q�'�=�2�!����S�yC~���[���7��P7���C�.s^�/����Mc�r���37=�P��>����=6~Y�b'D�xD��	�Bh�q֝M�۲�Y{ԋ�dv��nn)�y�����I�Е-�0����W��[�R�M�㼴����B�2{(����9o=խ�N�[m�]`��F@Z�����8�<)8��07%�'��M���D2�-$Z��F�i�]u�u�dM��Fp�:%c�R����tm��a>�������&�GxlѨh݁�Ո���sv�l�2�	�����
��|�� ��ȸ!�E4�����6[Z�&|S7�'�ack�$��i�+LVie�&W����_1�Ә|r`��E��zp�����\/��/Ǽ>�F��0�0��lDК0�GG���/�5"
$�$�&�����obC��`��sf�Fot0�3m�.v3��]�Қ��ԉZ������˾��!��Qd�'�=(���!�<߂�Ȧ��2�#>�rj�p�s^Qo�@X{����p悓h3|�70��4�[h�f�֗�ƙZ�C+�Yba����b&�ц0L���d����C%	�A(P�XܪN's�&�|���\i�
#�{xkY`�wC�휇-�+b� ��!�2( �n�O��G֗l�Fw�و��OZ]��q�ٳ��ݾ�.ͯ=���%��,f>^A�ZB�u�\�KL3J��÷��8{&���c5�ϜF��6My�EW���pE��VC@���p���G���Hj��V1$���"��M���̈�37�Rm��L�[�SY�J��e"z��$�Ǆ���-r�Vi�b��j�]��4��8&�M	�8`�(X;�I��*�1 �J�N�%�8oC�̂'��sK�=�|<-�&r�}�2�1Q5�e�7y��bCk�c肩x�"(������G�rJN?��6�Oa�a��2I��`�S�����b����Vw��ӟ xЛ�0�0��lD1��GE�:�j���!����م9�ZvB	=��X=��j��+�ۛ0���0�����|���O�6{����:�3Y���Y`ͅ
P-��
$FJ�z�����j*9z��hok�c �;���s�7�A����	dC�I�F�̗.���ϓ7��r���`���<뮺�l:î�鎎�:<0:� ��YH.3
�ݫa+(���&Q^QYf]��6j��8&.}�ێ+Ư˯9M�ԫ#K�����e�Zc6Q�ߍK2�!�醽ޫt���r�$�7,(ok�3�ۆ���C$6�u����I90��!�9��g��<X��&hM��FQ��.��M4�M]�D�W����8B(�6k▱mi��kЩ\t����(�D�Ҫ5Ĥ�؈.�ImF!�#���0#�l��;`��j��vd��.�5���c.�2����M���Փ6ҎB.L���;گ�A��Z�-k�{�8IƩ�ӽ�m/|yA�=��3�氭����A�&��+��9��7���vE�(l4y4&��u�V�{�0�)zYuuv�vs�H�!g�Ð8}G�'���(�3*\)���l�zh7����A���ezq��Zh��*�˰ˎ8�K4&�M	�8`�j��>�T\!�Q�}�P���h�,$�<}�W�!�C��3�5��M:��$� b[dI����0NÎ��Ӭ�&��ީ(v�7��zx<��yY[D�3I��-3N"�]GZ0�y���<=���[P�A�p�a��C��j�Ȗ�E�=>����$��zx_O����>8g���'�O�&�*Q]'��:zy��җ}Zh��za��zOZyk<��yl<��u}<��[��xJ�'J�l�8V)&����<�ym���O4��Z��y弳byo6��O8��O%����ż��]����y�ͽy^[μ����ż�	z=)h��>�Gc��Q�ؽ8gL/L-�ݘ^�^����z=;]3�ӥ�����kK����u�L>[/���o<��'�[�-�o'^[�����_-Ի���"l��$<aL�W�+��U���Q��w�gKӅ���/G����S��Wr�;1z=)ML)Cg�D�D�<��y���Jg7}7=����Z�kŧ�J۝��Y��z�����a|AĠ5�{��V�����|���.}��'}�H'�Gi�Hdk�od�s���f��X��^yY�醞/!�!��E����ّK_[���s>��d�Y�k\��O��:��Tr^���}!x�qc�OVZ�ẍt����+�|���s�/>�z��Yp�����~}�k�~�����3=�s����z����=�����z�����=�{��{��e��߼�P��6��μ��.��:�Ӧ�����^K[�U��H��ϣ	�	��,�`h@�}yB�qM@DD���&��8*���DD`̲��Q�=�Ḭ
��NJ�d$���6xY!�I2K%9��_f�����:ʸ��l�e��CpH�N�'���V�����@���O��#al�ϼ\��U�DD+�wjU�*�ӽ
���0��!�%%|03B��	�v���DD�'}[e,��0>8���J�=4!�0�%4`�i!F�;��Q�Z��Q�2�O*����|���4뭼��<�0�8�Nv�^��}$�T"�K�9M̫&jn�91p�Z�%XNl?"M�,����� �\$?_��B#l��*y8��
z`� p���c
�D>�	r�X�<���f�ʇVݗ�}���C���hX�d�0!}�����(�Q�3���i�R����u�O1}��-f�Y0d���-ޤ�" T(�����ђ<�Ϛ6"&�O�&�Ht�Bn5�H0d��-�L<����Bi%���c�<㎼��u��y�yva�Zu���j��_�L�8�,Ĥ�ejR�	!(�El��4�P��X��i��#Q4L�2g1��B��i�	hD�J�B"�<2qI#	��2I�M�I'�AVW�����Ӎ+�_�GyCCdm��mޢrt.�밆�#u�ySO-�1Zjp�ͻ�D����,�K�r���d�:��s�b 0a��	"��t����h<��q����f�?:-0hD���D�2}���y.䟣'�d��Oj�|�Ma�2B��<��F	��d� �J3E�gH�%�zF%�!)���UW��+I���I��	1��43ғq�'*J��Y�O?M'D�l�J:��,��H��P�etF�ս�jE������1���F'�L���5�w1�Y�d��n&�p�G/�̢��+���z�hd?Q�i ��<p������F�Xh50�ՂUTE��s�(��u��:�Ɲ�Y�y��e�]iכjyN�/ff�3Z;UV"!?�N����XR�=�,���n m9����F"bO���I�DN#!�EGA$�)�+ ���1����'��^xd3e
����*��Hd��S0э�D�"0����`~�|��F�؅�Y��~���!������60�P� �P����'�	���"w���˧>�3{�*]n�[�(��9�[C'"��i�E;��2ȥd���±��g �C,OߑTl0"gn,�(����"�̡0�/K�q��Vb��X�#	K�(�*ȫ�9��dS�5�%��N:���4˧^yg�]�Xuׇ�N�i�f\�ʪ���`$A��0���7��`�
R���(�e���2A�M��`���(pDO"K2�!C�z2Y'�5ވ��B}ϭ�B(�)-U��R�˞Y�TJe*O�lL�
�PCad�<��( �:;?"?I1˅B���&i?��N���e�E,<T�	c%����)�>&��Ѣ�s$Q���N,
q,t�*�"Ju�9�f�r`����0(�l�`""}&=7YL@5:��%�l�H~8	��t�DՔD@�
E
��f$PX
�3Z���D�DH_�%M&�&�l��b��W��X^RG�h�N>q�ϟ�4˧_<��.�,:�N�یm�b+��P��k.��bgz�����a�A`�ߧͷ����w�[�+H��B	A������@X(��j�<���Gm$K$��"Jm$E	Ip2�9,D�U��<��a!C���ZC�0ȏ���Qu�����RGY�0��z2Y>�dS=�Le3
pCZ��������D��
l�����{# k&~ZL	��E$Ђ	>��Q�Pѹ�I(�����x��>�#�����!�x�~�JDPXF�r�E��$J�dc �C�I��1�P��LdQ�FC�?2E��OF$���� �'�,<�FB��& �	���q�^u�Ϝi�N�yg�]�Xtx`��h1��f��N��N&�)|�f����)��3���D�%��t�Ly��D�����i8�($�\��isS�+��]
�Kq�<I$�@���P�e ;ˮ�$�beX�2Gk1
W��tr�MS�J�f�M��bM	�$FOt���,���'�!Az!�?1`���1�<	�!`¦=J��y��h�4���8RA��5ߋ��a 	��ȇ��ZO�hC�d���3
�\���sg��6�;դ�&�'�1 ��H~a�%��P�=-H�@F���$�!�X�d-!�V�1�(<�06$�6�ȤY�=�C��FI�����h�@���0`"§ ����ԇ��N?/>������7Mr����%�8Ȍ��>��PdЕ���O�I��bI�'��y
M�$��I�5W��U�J��Zu��y�2���,�˼��ӯ6�7�.��״a{�Y��v��$�����O�`��
Q,	K�`$(P�����gdq��,�%Yc�����Qhl��)��襐C\��||�Oa�xz	D�T؅AL�X��!�R��)����+�Za:�5�(��DC�I�<��/>Y,����&!"�}ϸP�uB+�L֛vM��o�j��?	��EY5Js���t�r	)?JJ'����M�(���7Ģ#ƞ�)�d�` ���?]kF�ӷ.�t�-��&X8�8��i�N�yg�]�Xu֝y�mw�_Z��k��Z�m�a�*�!�D��XS�~T�v'�O!�a�'�lb'Ԃ��Y���=Kݵ��4�jpM���B�֚�Ɂ�(2	��R1����gQ�1r4��R��:���_�E��&�/>��gf�Z�6d��?D�
^��	NM`���H`�%�I��-:6�f��<�ƭ���p�
�C��bg�hb)��kd�����>7O!�)�t��J�&�D��SZ<�S�d�&���Q&�)"�K.��f�Z�����s�ˑ�-���|�ƙt��y��e�]h����F��3����P�R��󪪢�(w�g��Z�h�N�(=�����&"�<5��-O �L���r�Ս��uʴl�:2'��,�
��i�O�GQ)��SXt�za��ˡ�V��ӫ����9�#�6�U�����R�GQo�<�dB�y�\!�i�e0�yIM��
�7�!e�so�ɣ|�̺qP��U]�L��*?-Uh�.�0`��;56C��u�����V���\N>�Uv���uo�y}>[��/��a��{3�/���:��OI��yŴ���e尚]o.��Ɩ�弲�<�Ly<��a����eo'^�����x�8k���<��qo6��)�Z^�w��y<�h�:^�2�������K�z=].�e����yo'�y'b�ˣ:	��K��G�ڨ�6]�n��*=z��/O��Kҗf��K���zw���ӵ�:ah���ϟZao�/����X�.�Ϝ_��(��'��D�XO$��<l�OjeM��0�BL<V)	e��W��N�����zp�8w�;����zzd�[/O��(�.����*��6��$}i>K0��t�}u9�1�$h��
W)ێ�S�kB6X;�w�AΜsv���-��:�`��Sݙ23G^L9S�2���\�Py2!�N�*�Y�SSBgrdU��m��L�,xś�mJ�5&
�W�I��&�()�z8�Kz�)�]$��_K�ȝ�ƺ*#H��C>a3\L֮��x_'+���Æ�
T$�57�Ae�	`�7�V����&36�3	�NaZ�����"����F�u��kS�\��Lc"��CU<��.��q"cF)g�5�m9Jc�e�Lp5�<Î��a��U�V3t�=�X�X�s���;=Z
<ƴ��m��W����1�	��L�1�����] �G.��X)ϸ(�exI0[.�J4�Fc���e!sŒ�q�Wb��\W�ח�z��Y��-�#�W*��iDq'%�[$3�)3L�\�YiV�i$A2�J�����oJH	$��L�\$��d"���E:ٕƐ|x�l,��j5`�)�ʉI[(��u@�C��R��N��H�K�e'cc�Zb��qJA��*��������v����̻����U_{333/�Uoٙ���UV��������	�,DL:pAy�yw�a�Zu�ܾ��^ZJ�_��1�e�k�SV��i���ڦ	�58�ДR��T�^n@�F�z��+�Nm҆�,��� ���m��,�D(&`�� �-��1JD�G��ɰ���ό�
ʁF[l�!�FȎ����1�c.k�ftx�� ���"I�	M���T��Y*&	%�
��5��,���KD�LB��I$�v��1��&�lay��)uAc	��8��P�+U{A�E ����`|��=�+'��<���9.����_uL<N���֩jxy3÷F&�����B8`{3�ԡZ#�I��I���77���;���)���ն-�kb�#g*��>��E0h�6�#��� ,��e-��G�!�0C�ɒh�y��np3k�~o�R�R�T�ڍ�b]e�3�}�s��گq�[�u�[C-t���1����ƥKXgt�X��iƜ|��2�מY�y�u�^m��+�{��WYnsgj��8~�8"y���{�{�BÛ���e˝�������jh��	0�/3�i�-�Y-�d��W�~0f(���C�F��3���i�᲌��h�K<����A����^r��#_���{O�b�嚭U�[t��]e�ȋVz�nT�^i��6�=O4٥n��BɂK���!FW[��/k˭N�:��㬫Q&��P�ζӭ��ƙt��y��e����ᣣI�<�|.Q�	�cXg�3e�y�ǕxSfiUQ���蘦�if
Y���q=��8G���g ��Y�vBD�'$$�<������D�"`%�3��?!�����_��]�PB�o��4D�������B��e��	��2_Ñr�{>��
'��^�O��[2���LR�bS��F�/���N8v�D�p�f��0?�Xh�}m��������=h���>(|ڙuB6��Մa�θ�i�N��g�a��u֝y���csK�lb����I"����	��O
P�tò��:2����@�#�	R2ն�-��af�Ӿ�Z����I�~��h�0�8`]����><�o���m-T�]�G�Vj��z�Fk��\��w�m�|4�p�}�8�M�������7�X�/�-M=��o��c�#���D��S_�d5�g�4���#�4�OUY�f��V8�MU��4��>u�δ˧]yg�a�͟8sf}��H]�c�&kk�����C`J��D���1,aM�,p�h(�+�a�3Ǖ"�H���I_l���%�e�h��ICڋ"�L����N��$�H p�pտ4���9Z;Ǳj�̈́[�.d��FD�L,Y��Ԣ%�`��3<�CxHb��4��kz˲q��T��9�v�a?�����[]�OD�&����'����Y����D�Y�����1��.��s�Stőz��Im$�k����߫F��s�j�n\�3'�NC��=/��<W4n���an֯>��|�l^��Gi��ޒ�gM2�>u��8�֙t���0��:�N��a�bObֵ�W̒I���Y^��_���m�z�3�Q��p���ׇ^_��nd����M�CP��&���3���ILS�ۥ��>�����W�D�w꓎�1��ORaū�m!���,��2���X�ű��.�܌%�x�����\�N0-f-��ϟ^ז���8m)f[{˪�'���!'��
�]�H�A`�mZZ���#/6���>u�]:�<x�ƍ���񒹪ٚ�r�z(��U�=:.M���:a��i�x��u�v���iůԾ���3K!zl�Z����ֻ���[��	�AA�c@bp?0��?D�=���*70�q�aS�hMG��(b�ܻ8֩��Z�\장�gkd'�ٴ-�V�Ń�/���w-�6�m��=RIo��q�Z�w�|5]��rpC��z`;ܓH� �BWִF�jѺ��em��<��Zd�$<x�ƍ����n�>�jju��3�nmUQ������T�њ�%X�!�v*�1K��c���l%�{E��@��-�!d��+I{\�/�����iu���q��f�9;�|��=V� ��m��Ї��O�2��{���R%X��8쩖�=��
�٩�t�00�s������������87��rh�$PI�J-��>�<6�,'��e���l�ܬ��\�0�n�i�ݦѦ]u�0��!�Ǎ�4lD�7�W��DHUI1Tr��@�Q3��R4��nQl�C���ٶ�0���L���Cm�!��P��r��J��D�)Qd��`"�H(ऒI �?L��@�-L��}�\�,Zz��pٛ�����I]�D���q��S
�qǽR�U�Rz3YDb���{��_�N�L?|�xi2�0�~�f)e���e�2�M�����eh ��0��?8`�w.%3���s�?�a��>�O7����q�6p-	�<כ�/����r��y�70�o�������?C�k��z;()�����+�tB���TDL�&�@�ߎ
97J���iu���;5M8�0�)�ZM�z�x�Lo�4kԳ/,�.�8�ǝi�N���y��`D�1�Ǫz�:jsuZ��}P��z;��m޳����Ҫ��7烨K<�?�����^�V�'��Y�C���C��uiioSZ�Ö�DW�^�r��r!ֱ$|�]mgu����5������h6!ߗ�-�,���B8C���"� ��tQ��၃��h���?O��wa�=�8ᖞ�q�.�y�&�[,+r1��T�[�v���+�Xg�w�]�V�帛|�-�y����yo'Y��4�igM����.ǣ�م�J�C��N�җ���5���t�6pΏM�����T� ���I��i<V�����Ҝ:_c�OLK^��k����/Kӥ�p�M�2�A�ѯ�L�e��W�[�-��qw�*x���L��J'k:Y�v�*l�;�KҔ镵�~)z`��/G�Ӷi���<�^[˭�ֲx�<����>f��1�V�>_��kyծ�=�U�L&(��$�<WK���Wq嶜yn'���Y�����*y�=./ó����xtέ:g���+ze)Q:�Jt����J!��������wu�������;�}����l�������XfE�2�H�>Ί�b>�ڳ49*��C���$@]���cJ�'8C<����Dt.!�.�aW:�9xx �Ξ��|�����Գ5c�T�S=�����&Y�b���(i���4�[��=���=���	ӄ#�G���Xyىa�H�qY�:H7�����o��������_�fff~{�U\�fff{ފ��333��UW/ٙ���t��<x��xǝi�N��<�.î��̽$�H�����]�|�1Z4�|azy[q��ku:�]]�k4ac�Գԏ�����)<�|�UqcT���)��k�χx0`��*�e���8�HZ�]���}M�]���e�����W�0t�T�ēU�.�a斚m��0��f|��ִrD=�,fO���Ob��mcF�u����#��y��y�]:�<��<�:ӯ1ɽ�wR�f�u��*� ����~?|~&��@@@:�@���6��5G��.Mb��-2��F�)������M���>��q�Ś��-�i�KRԵ&5���-��Z�����y�>���.�i��������1�����(k�ޗg��d��m�+j�YcLU˻|bM��ea�8㏚eӮ��a��e֝y����|`�g�' �I��h���ik4o�QK�5+�,ۈ��ݰ�(�4�H�*��B?��(�l��IЅ4�B1�Df����#@7l����0��fH)� &5���,�-��k�,�����=2�w�I$����	���O��N�<Ծ�U��ؒ�R�F���C[�BR����}��"��A ���o��N�������x��6S��L^��k{��8p���4S$�v��rK}M�Ӝk�Uc�������Q�Jd��^���Z�6Ѫ�W��k�����0Z�MӬ����=��B���aэ�I<P0P�>D�-���S���=��Ȉ�3s���P�im5GӅ�쉇�4h���q֙t���0��2�N���F,�UTHɼ_�6l�牚���/��ѐ����ESSQ���r�._�������D6q|0��4��v��kYZ�iwqm۲0��J�yh�""��32�G�¥ˇ��p�7>'TDM�|~9y�ҷҠ���t�@�n|hՓ�8�&�Y�'�N��K<ۯ�q��2��Q�a��e֝z������FU�ӆ����}>������7O��I#�Y<�,����RW�3�-�W^������)����LL-m̮I����������2hU'OU�l���%;>ן��a�up;u����)�P�>��D<����6��7�?|����8_T#m%�i�4��<�l>qf^q��|�.uy�a�]i�Ѽ|po.�FN������@�R]c��Z�.�fE֯R,{;g8����i����#gܬ�EE"1�1X7^v�B8�{���{�oQ���늹�7kU�o]��{".O��Ȗ�5�R��{��V)ߝ���8i؜���P��L�J���3�����mʆ���St�2�_ywYY�^q�|�.u|�0�.����Ҥ��q��i�E��q-��G'��)�:AD��ǋ���dփ���ʑؔ@0�L�%�t�I ��F�oY߷[\X�y����ԳsL��8�XIo$�t�;l5PG>$j	���$�qt���'�޹�ia!����4Oϕ��K�@��e�aXul��������2��g4��)�aXd��}��m�;���,uj��U�w�SI;���+�j7�k��`
gAo�!�4S�nx��r4
��:��T��	#�^��Ye�St�{Jev�D�3��S�[af�<ۮ8��\:�:��a�Zx|t݃��ō��Z03�U�U�UM�9
N�A���_H��^����q���V�=Lz�7ǟ�[=��f���s3t�A������4B�엌��Fi��3K�K
?��<���{�>i�����A��$��eq�t
<;߿P4v�%���ib�s�g���l2ӌU�;�I��י��wr��g���|r�å�uf�u�q�L�u�u�y����<x}Pj��tV�Ԇɩ6VID9ꈨa7}�[M�OC4���*�>���(���ӂ=�����n�=ԟ6�;��U�8��Z3���Ż>I-|^Lb�Y�, �0�.�R�w��@g8������t��6d����Q4`Q��$���2���ͮfanfZ�e�]���ֵ�3NR�zinq��?R��l��o��8��\:�:�y��|<0`��Bt�`����p��G����S���$�$���|�f�v��kIg�����\�lE�-2Jm�_p�C(V����t�r��ْ�kQ)����
��-K�Z�e��L�9$�j�+�55=�y�>��9�i�x'L�	�||~�}nP缲۳R'�(P��6��n��+t��gt��um>[O�u�_'_>_Ϛ_���O.��[I��֓�,�u<�l��Z��D�<�Y����兼�ךy|6Wd��Z'��H���ŚI��kέ�m+�q6�����F-��y<��O<��yn<�Ɩ�y����<yo,��y|���i#�-���æ'J�/Jt�#Jt��S��X��w�e�tS��K��*�aN�^��ӵ�|:^�N����iiҧk:T�z=ƿe�3�������o�?��K���N�ӥ������K���<L<U��5'�	���tʞ/Sée�|�C���zh��ΝǇ�zt�G����=�J��z=���N�C����z�9m/��t���h������[��o{s���z����N���N�l�f8kUŪ�[m��6��5��\jV�WI�TIh�#~>�ѐJ.�H�gc,��B@�ņ�C����L5!�%L�U	$%PS���L�n�Ak���ҫ8[=�4��6��j����)'��WK����뉇�J%��1F�����R0�KT���+��c
&�"���[�|n��yL��*	�	���҄ׯ5�Br C�]�Sa�׭.�E.�����N4��@`�m�\�/gd*D��8S�<=]UVza���2=�F�Zﺞ���J��;�]8B>-����$nN���^�P}��>�Ip��y����k���W2v�K�5�"���x���fPI��2�P6 �C j��,9gj���D�.#��Y�4G8A��{x��d
6|�Ǽ#UdL�]Ds�@"^����|<I�����*%�SU�Ȍ�Bk��*��%���1��F�h2鱴R1,ͨ(9
|�v��p����p����}��}����f~{�ʫ�����{�ʫ�����{ޥU��ffg�x��&	�	ӆ(��0�:�N��wU�Lc�Lg7��R՗Mǵ�oS9��Mfءx��B�0�Y���e�f��ٶ��ƴ	]5�m�nq��nB���6�Mt�.�D����P˥�)���-Q+L�a@��D"�1��@M�b��!ㅑ����O7-�v�b�v�b6U�v��]��\�%2�*k���6��	$���w�'�ye���*��m�Dͪ�s
�10�]�꺵�kܑf��Y�&���k�֤�U�8������MC���Ϣ%3pB�H���Ui�~q����,^��,ba�����f�%��]A6�?Bx7a����p����9꛵>�
�h&8�ܸwbW-�^m�����!��1�qw������{�kKߜ�L��2ӏ<�4ဉ��g���D�کʩ(�Yn�L⪢�e�f�XxSގ/[X�<�R���Uy5H�[/!�?!�R{?>"�jǂ�V����I���|�m��;��dCs�=+�>��.�}�UX5��I/j��p��e��Zh�o'�����������|�k��Sa���+S!�*�1�%�z�4�;����Ye��<�D�çH"x��g���<V>�z��4�⪢B���3���k�iKL���9
P����E?AX�Ύ�����XI6|XS����z��e�?`�5���s34f�V�U�_�M�Ӊ��Ca��C���Ǯ�Y.��xo(�:v����~:�k8h��ٜ}���Oj[WG�/�nH�X+����'�kNf%)V�G$A'��g=]���{���4�0�N���y�\:�:��h飧�����V�`TηM-�UQ��M�S�zw�z����`{�դ�`L"B0���Y��WƜ����>?}:7��?	b���Gs�ke�8��f�Lmzf�e;[�����5YEϩ��mmC}�t�MhM�N�XnewN�S���*���D�k��yzb���r-�Xiv^igm��8�L�u�uא| �xQ��{c��"���V�$�q����)ah�DR鴼ˁ�����0�Iq�-�\L��,�Ŗ�Zm���� "I�����I�|�(a�kȞ��Q�UX���\�s/�Vd������7��+(a��]���"RC��c������R+;�Ě����0��>��������4��fęZ���]b*�n��LTFH�Բ��:�s��ֽ��i�'l��9_Y��aD�f�=�l5�֍z�+e���S*��~I�L0�3�;2��O�X��m<�y=OՉC~.��,�,,�ϝy�i���������������q��Q5 &�I%�D�R��VVjj�YbW���؍���M���R�Q��މ>�}m����n�"V>����4�u��itp�}��nYG�xCpaC��t�˩��a����f�v��Ĩ8����XS��K4�d���|�LJb�r���G~��r��$˹d���,�g*�Ԍ0�ytFW���|�1�i��q՝y��\q֙p� �����tN�;�7>�I�K�T�Ȉ<p���$�A��.͜�v�CS�'�����4N��f�oP؅���Ut{{��vpDC��h�,C���jh?z������b��T`��H$��=�H8hىg��Oba���a�F ʸ|P��6!��K����jx*�y���)����JP�)ِ��ޣH���9J�>�֗�v��^Sn��]��L8���ͼ�:�.H"h��g��9��T�_ӒI$B�3Y�֒��_e���4�w8K�.p� |_�$�<D�L�h�7�f����[��9܉�L6��S��5L���"�"賄�D>��Kh�<��`zC؟��Z�V���~0����a�ҝ�g::�a��MxQI�����m����FL,,����O�z~8��:�.uuw�a�Zu����h9K.���4�G�
!���&@��s�L	��#,�Cm�)02E1�J�`�DD�i�['F$[2���I$�@�h!�{[G$R�R�GA.��q޳�&�Wh,���uU�_���k�R՗���v���t��VY��C��G��S������쿪˅_C�G$�F0؅s�x��̹�fa^�����&L�w���.�ɰL�;�'P�~2���o�D��wE<��������x}7�æ]ZbMmq,`�r��t�}���=�e���f���������yfK���F�R�|��o��vG���Nm�Ym��u��8�L�u�u��<�δ<0fi� �Z��dp�C,���Ƒg�*�!�Jp���5�ɲ�0�������|8p�҈{+�cZ2��V�}&Q��S+�j���{��nrJ"&�}����!�zPA���a��s��YKX]]f�I(�%Rd�'9�F���NR��!�>�}�-������h�3��p�M~�ܹ��V�p��>F��M*�E�m��y�ʹ�n�㮺ێ���8�̼ͣ��<���eAġ4hD؉��	�ab"t�(�0KtK:"a�F��"""tDL�$(� �b&����(AH%�&���6Q��J�(J�:""'!B"%<l��:x�g���"aBY�,L���'�aӧ�"Y���$N�ZDMt��|��EA�K߄߿=뭿������ɉE����D���:�FH�����u/+��դ����٬��H�i��UFN�)ڡ���,�
$rWrg��F�5��{���=�(�s�:����:����CR{u�Q��l����f�ʫ�'MH��w~�̷33=�z���_�33���ʮe�33=�{�Us3ٙ��x��Ƌ<`�`�8X"AG^a�Zu����DI#ؒI"��,~u�u�3�%��/���Ŝ>V�B=�%4��n�������>�����PC @ކ<���ě�FK`�O/]{�:D��|Yq��r�SkR�V�j�wM�!��}bZպ��L�W�O�3�>���:ee#�0�0�!�/m-�lD�6pJ<tMa��'N�DО6|<0xQ�q�D��Xd-�hH{I$�!������.%m�Ð�J~4PQ3�8� @3:�'�5F0\���H�T���.�4���Ӎ��"����L<�����2���גjq�Y�ǁ����cZVa���"!��Mh�(�5
!�(qMhl�Xa5�q+*�?	Ț:S`�ɰWSPѾv�m�ܥ�|�]��>q�Ze�D�&���tN�9+9��k�Z����Qa���-�u2-ƒ(�b��6���y	��q�S�+��%�	eR1�bb5 �2�0*���bB��PB�-�$�AnL�P��e��:BUp�Kp1RJZ�����\��An\q
����B	�Iv�מZ��)f\����i��4�|�ʳ�}T��a!�a �0SG�*'���p:�&��\���ݗ*���J�ZZ�r�����Ѹx~�jO�E<4*h�8JQ���.�
Q3��<���<BC�ON�����~��?p�}aCs����]��KYkS�K8�N4���u�	Ӆ��DО6xN��5�Ϯ�wF�������=�t��h�D4�6&��"�LS�I��z�Y�
���[��h>�˩2L=����>��z�m�v���cy櫕����?~>l��"Z2��(���:��)��;N,�j��v�}KS~.N��ᰰ���),a��-0���u��>uȭi�ߍ>]g�4�fx�������	�8{�����Cu��W-�̥�{i5��ߊ��{i�M��M��Z�[�4 �O:�*�a���uj�e��ewi��gB<�^�����݁T�1a� ���9��1����f�0i���l�`'�?~Q_�F��y�8�����L&	D��X�d,7��c^_	e���5IZl��ũr��y�qe|��8��^u�i��uM	�g�K8o�r��R���$�!��u�n�k摕���Y�Yg̖m(<7�{�j�EsT��PTֻ-������	�d).բ�D��}v$������.1��yQ�<븥�N��l���s����2�+.d�9j^��S	��t�������=�Zp~�鳦���,<��
:'N	Æ<~	�	g�(DО6xD��}}�|��Uotk�(�d��G�	y�Ȳ��(���6 �:�L���02;�0�8����I4��I�Yl�#k��L�m�3m@�"Q&՚1�&68K45ʲC��I ��wF���I���_$��ǳ�3�#�#$lĢg�g��3��ys%P��x#&��/n��<���!��}b���O>n��\�+��ԵZ�����l�4lJ'��r�8}���2�}�a�r�Y-XC��%<�[�@|�	,l~)A2Dd�-�r���n���^�8y�CP�;����#5��]�8Î�q�[d�%����{�UQ���}�M�ie��*�!�Yߏ��SD<�v�X���2�Ȇ����v���[K���l�!���r��n[����s�i�zC%2Y0ٲ��Բ��
���GS�4�L++e�J��mZdE�̉0���3`�@�R���M��2q}j	������t-Vd�8`��f���斒F���vO��*:�ii�i�v��i�-�����6x�<a�Y�0J4'���8Q��CN_�UTC�Sä?5"�o�ONIkW������r���Ze���Gԛc���[����b�::G(��(�A�#eP�T��ov���{���im�K��7��'Y��'j�2��B"!�57>�٦�J��S�_F�]��p��:>�����"{x�L���u�k��Ӭ<��<�.�J4'��,��7鯸Ca5$T+n\�3�Z�=UTC�'~�ʚ�k.����\=�<���:l��Jn���f|�S�}�o�����,B�	���!`W)uV�Z�;Uvk���b�6��#%�QϷơ�,<�dLk������><>!v�������ͦ�mYr9��+j��L���W�$��ү&)�FUUf#L�w1[f��ޔesRK:a��O���gO"`��c�����:��0�/0��0�< ��(Љ��&��0���0��&	btN�p�%�f�:$!b""%���!BB�A��DL�A	D��a���C`�$�&J��"'DD�8Ad����<x�ǋ<x�DИ&�8%��a�X�a�0�bp�,��B��"p�:%�&�l���	f�(�	"I��V�R^��I�\K�;��R���ɸ����
�k��VG�u�<��Ԓ
���³��Ad�	�<e���5�ʎ�n��Uw4m�f	���&:�j5���O�=����6I�SN�<T���;Ym���mny��fMNK�74��3οiנ�3���`��:RJ5K&�I$�B�or�]3�p�K�r���K �*҄(��)�q)�%���ĹHt��z�$`O� � �v�۸��M�,�����`Q5��|n�œ[k��R�K�,9�r!��Ԏ�U��'��x���4<"7�2���'	j.�{�����n���D���8��p%*�L����,U��kj�q�H�Kq��n<r��c�ev;(yw��78PkKh�J��rI�-,�۝�:���,ƺje�@��cZMv�/��;������9M��!*ϼ�,h.7���5�h(g����>�E�"ɾ��[.d�G\P]�b�� \���R����W�՚:�lN�8Fu#��`n&��I,8��j�X�a����	2�h�ؠ6�I�z̭C�>�����eg�|���s3=�{��f_�3=�{��f_�3=�{��f_�3=�:x��	�<Y�0J�4��}��|ϙ�/�v�>E��TrK]��X
[�B�Dn �:����T��퉛,&�&�Ԅi��X��$6�p��"*��(]�Z.�l�68a�b� �6���a��,۵�f��\r����hZ,I@�XC<�k��E���d�6y�t�.�iolQl��E@(A+���	i��OI$��j#�F�I)�<��F �:U��'��pM�.�;K٫J�鸚a#-jD���F���+�Aة�1f����P.愽��>)����َC Sh�)���̳A�g��0���QS�m��M.���˫�"�F6�O<�>��wwE�	��P�B���r��l>0�[���a�*C���Z��p�8vݎ>�Ụ���U����Ls��|-�'�aT}�%��U)�)�I֫��2�~	f��Ǆ�ŉ�P�h�G�������q�sH�wt6�mXa��u��UQؘ'F��#5v�eWF�R!��Z"�i��)��0�����_�g�p<�����5�fj��V��~�寯�ͫn����9C��=���6�(!
!)5�f�U9��dzӐO���84��kZȦ:�4}�a�oi5K�b���3��|��n=�����Ѳ�2��|��m�Y�qw�q�ю ���B�!�g=��I�{K�f���W7�����_�'���>�^O9,9�3�M�p!�S���������$.�����>�>j��nI̛���/��@�L*��mJ�y���X�|���FW�QG;kV���Ϟ���;�Df��S�1P�js�Lĺ���.�2��u�o]eZ�,�UѺ}�n+��-��6ï>uǛu�]]��aǜy�<Q��a�4������O��Gi��f�1
��]z��<��û�kJ�edq��C��VQ�/&�6�A���&�O|�/Ӷ�b$��)~�9�0��MO�a�ܧ�W�i�.��K8��ɄP��h���(ʹ��ٳ�>!O�[��4��ō��$|��M�h��U��$��9lg8�n��[H0�̰�O2�:�ͺ㮮��0��<���t���l�0�/,�DRf8�H��Q��a���j4���AB��%�P�!�KM[P�%��2�SU����ۏ�$�xA�=u�<I���6�h�2��&s#�em��o$I°h�M����iD;&�����+�Z�˯V+�ZF�S���S�-�]r���ra�d�0�y���?�3.]�+�r����r��#�Uv�e�^��K,:rny��F�Ǵ_NB"0OxY?h�y�߶:օfi��n��6|&Ϧ���}O��tS"��b$�������e��:�ͺ�F0ه�<Xd�P���ItkM��DO�ɮx8���C����4"z~b(�dS�Ap2v����Z�tj�O��7*|f��L�|�FD�y�Ƹ��a�"{��}��'��Q�O�M�|�j��ĹMRD\�J)���<�g�B�!������`�l4��R��*M9Z�-0N��a��u�S�҈	�Ĕ܌��lS�R����a$����<�gO	��Mh�f0�d����-��0ent�O��U���-NI勢%v�Y��5Yn�e�6M����0�>,;'�����h78&	�nŸ�0L���z[�_�,�>y�����9~[a���ѥ�:'�"�,��2"w���T�'�lD��C0�l�������<D[p�=�^�m��W�iv>q��>uǛu�]]��aǜy��ڴ�n���&n�E����UV"S�p�:��Ǎ����â&J~�g���Ȉ���a��!��BmD�𼉒�H!��gu����YeN_]���*��Y_�i���!ܘ�����y��8K�Z|l��N	�'>)���<]C�
">���0�ߝm�4�9�������Իk��/�2���\y�\u��]����>5���?T�L�ce�K�0���&�I��	Q�	�Q%4	b���m����EV.]�i�Y�a`؄����ܮ#D&�G��i�$�xA��sw��{U^3��36h�|'5�ݶ_0�t�TԼÔK������WN5�r�M����e�jT����.������荒����a�:mrL>��Q���ꋣ*�wE��VFi�atF��EV�jf�y����.�V)F7J'���Z0L�(�z9߼F�"� D�Xn�٠ِ��Ȕ�Q9�4�洃]j���o�*�\�g!ӓ�h��}MQ>���FR���k���M<�˶�ͶN��0�bX��l��,�j�洗�0cuS1����>�aa���n�P�<5w��k'"0�e)����݈�ú�8�a�R���-��0�"��a�1O.<���K.�f*�Sn��6� `��v��T�;29��4�|`*��M��!���$L2��M"�V3æ�M�O$XS� �g��}J"_��E�8������YZ��K,��4��<�O:�:��]I�:t�8&�٣�h�F��Ǐ<�,���y��i�[u2�&��0K�t��tN�l��!�4""'Dw"h�'� �$4��DK�A	DA6�4QF�H%L �%�""X�bl�:u�e�Xuw^e��m�y�""l�6Y�,Lĳ�����gN�"&Έ'D��`�gN	�"QBt�EA#��=��`��F��u�*��2uUĻ���CfW���ut��G������3�9��1=�����qC��0�Q38�)�T����0P�)���<g��$���̐ע�G�ϵ?w��ݷ������Ra=�n��T�a�^s��^컹�GD�l���ߝuw��+Z��k�Ks��y��s3=�{�ڮfe�3=�{�ߕ�̿fg��{�򹙗����<t���:'��ŉb&�4a�x���UX����2�>��̷���4�&����u��>7�L<�i���pL3ť�F��ί'�͉�`�ɳMq��d�z<-��[�S,�������ϲ�#�����?��.�م��z���2}_���dZ����6a�]����p�xk��(`��E�~^7=f�摷m�i�θ�n�뫸���:t����E� hf�"�t�Տ�*�D3��#�ٺ�^��G�*U�;�q��{v��-�+YԮ,	"��8A1PykM��X2���N���i����1���U����C�2�w��*S_�)�7�C���Sލ�Nl��ȋ%2�W8�)��f�dF)����z����;Fܽ{�q����avq�y�\y�[u��]�m�kS�@R��Z�ՋE��$��8����&CmIe�(�Z1�
N����<�*U�B��E(وĭ�kw
.�m;��0�X��I�o���E�W=�0:A��5G��ɋ�Kj�r�V�}��t=Z�b�j��Âp5�˽�����fB�	�M�OO�ȡ�����a�������#H���cFkJ��Yfk���I�OaO8"�C'��D蟡�p��`!�D�i��	a��dB��F�F�"�|p��Њ���(��R��9�U��ag=�y��6㏟4x�%��0ц�,�����Q*���J`�5M����N�f��M�两��G��4a��{�م7��n�9�r��rxpK��mD��>Γ�>єr�|�x�}Vծ�:x���p��-�RL��]>ц�����{Q����S��?jnmv��ET���l��&��r�D7
�2��<6Q)�K��Um��c��|��>e��4��\y�[u��zh��ӧ&Ǐ�q�{��ta��w��6X/ː�aDJ���<<���Z"f��~)��[�=�UL�SF��'a���^���:W0����7����4T{,?��{�n��ȗ����%�m.��ܙ8��OZnى��z�'�R��O��:4yF��^�Ëct�|�nD�Iq�џIg7R1K՟4�N��:�<X�"hMl��,��
�BM�"�NC� ����w�Y��0��I�;����n����p�L�kF�G$���,�o�` ���r^����Ua�q�eË6�)���Y#�s�!�j����oze�4��k����;W�1R;\����Xi]g]������X�#z��7��]�:Yb'D�x�,D��c����i��mTڢPm,�eI�ԍ
��$+/rQ��!DH@$
1��)lAS���,��,,2��1^0V2�bH%FT�,Yt�H�6�mf��Z`����(��(i$���=��3��lm��*�ᣫ�gb#�zcI��pf��U�O&��u`YN�	�N3&3�n�g%�穚iv�j�#.>�韪O��#�[�Vm�q���S�	�y�៩�tOP؜��M���o9�,���福qxxldR"d>����ƹ��Y�'�
DD�c��N:�֌�ˋ�d�'DADJp�>�i��a��#'g��Z��T�ߏ8l؞�D�x�,DК0��çNw��q�LM��D�f㇦�N4'�?eTB
�<6n>�.��q50N�Ô~����iGc���zuߵR�p���z4��!�Q��#���Q=Pa���	)2u������r7��XS��{V���C�Q�,5�S(lO��Y�������E:Yb'O�a�ıx1�F���A�A�C�ˌ�SDa����ER���S������z'��٨j	�)��/oE9Za����e�f�=L1N�,�o�ֹ"(J�����"H� ���e)]�Md�6��ũ�������F�6���^�:��U��>�ܶ��p��/4QtEJ�Z�J�.�VQj2�s��if�a��㍾i�θ�n�뫺��8��N�ҍ�6�">*�Dpl�>O���,�%ie��2��i��/�k���Ȳ�6��m���#���vϊ'>����OQ��L�L���ᆍ�7=�\�|��O.C[?{���^%�&@��Ӛ�Xw���'�.���R��ϩ�����������]^Mjw����i����q�]m��i�\u�\�,���4pJf�	�4P��J,CB#�<x�ǌ<'M<h����,L����4pM"lDDN"htMP�l�$bX'DD�8A �Aa�ٲ(� � �A(DАDDL��D�tM��7�x���0��L<"&��0�,Kl�B��gD�H"&ı:hK8"ag�O�D�4!DB�K���G��ʫ�'o��{��Ѫ�~�{Xic��P�F��v�Mȣ��7M��h���n�Yx5R\+a��5�Sl��SEq'�A�][�膡�����^��`�{��2�g���p$p��a�]�|&��f��mR�@���cޗ��fS�l�1�h�H1ldF�h�MA&�FS�71��`�{_p��_nK�}6-�Rqa"3�����]x7]��[ f��X�2Yx�7�iw���^�Me٨�P�Y-��#�"0�"MG;��H�۔�F$"���nc�$�5#�����	l݆lOH[#W;;����Z�!%��!O�ru�����V��<E�aQ<��xCa�6*#���2�g�zW�o����E��i�"\`��n`���d8�!�P)C�7�rH"F��"S�(L�Sd���6�i���i�HBF(%�\Z����n���V&���s}Up�G,-��.��w�7DH�n)��3I���;Ĝx�f���Am �ʁ�A��\�K�
�!l��DT�k6��7�n���7\��-�������=�{����߮�{���Ż��]�����qn�﾿{�:i�y��uכu�]]��a��y�>���o���	���Y��-�2��o «s�wY���2�eS���Ўq��J�"�`�"�Bc&�LJ��e��l�S40c�N8O�0�i�b��Hͩa5�ىs�Øk��4nŪS� ���6:M�$ʭ�&ٚ�1�!i]�h���[l�Sp�HܡKL���� �Ֆ0���iU&, ���XA����z҄Y�g�NE�|I$��;�请�U����̸�"!��\�v�����0{=��RC�$M:r��Ga��+�L<�ܼ!�O�
hN���ѣݭ6%�
_"�M�h`�=����������5I���ݴ����QD���|�eE	e�UEw���	�NO�����9�oM�n�F;+6�Y����1�Gp$G����x{4t{�:'�)罾���2��{��t�GN���<"x�ň�>0���çN��㤕��ӃRr���ٖ¤�X�U��Y��s(�erZZ}�]����5g���������adY�va���Ϣֺ�#�k�rg��K��J++Qkh�ܥ=ׂM��J\�\��pop�%�ob�O ��a��m��yM�z�
h�n��,�=��-y{�n"Dm�b��M4���u֟>uכy�]]��a�Ν8v���������p���[]�T�|[q��1�濾�C�<����ja�a�Á�w�̳>9���3�	����������؇��k
�Nj��Ѻ3�w!��g�ȳH�<����ɤs;b�K��4��m(ú�I��_*��O@����lx��}�����kb}���{b���߽��[���4l�0��<"x�ň�x1�F���F\z���� ��+O0�x�I�fJ�c��p�l��U��1L��H�z������d	���B�T-��M�`3�`�y��kz��N���&)�қ��P��xl��/�6��3PN�;*S�B}��|mf�#9�$�,�ӭ���0�a</M=cH޶�i$}N6�]�Yq�>y�^m��uwWq�[y�ݧ�gq�+��6J��;�J�ǖ"q2ۍ(���M6��i3D%�I��9�_#cd͉��'8S��k����P釞$�xA����|Zyf��mϗZ��.�cG-o��u.���DѤ��t�HEWz�9-]hY�c�ɽsX�V�PH5�K�]�t�;�NJ��}'�K�����-�#�s�B&j)_'O~�O1��hũfZ��=obȼ��F)�w	�erSu�g�i���kme�QrvvJ{JhN��=�����X\,��]ak+(RҀKm�bbZ�i�Ҟw��E�c2}L��\i�̴��y�^m��uwWq�[t���{�K�\�#�4w��<<�k_,�)�YeѪd��i���f��Ȍ�[���n�Y�IXc)l�,�S�7�r׵����,�ӕXC�T;�6Q&7
������"��O��hN�0�u?!� ���ak�z�#��YZ��,�"R�����۫��M�>:h�������o:�ͼ�ή��8�o<۽zV!���d���p�3Zՙ�U��<�+��)γ���e�:"&��n�������'�����^È�E3WX�O���eP�	��$�	R# �Bi1�3����ډGF�6'�A�"���D}==����O��D�ϗ'�g'�~!�g�)D��Z����7KZ���Gڥ�S�K�ˍ�y��:�ͼ�ή��8�n�9<CɺLJ���W�V"y,��u��2��#�ӄ�K%�O�ϒ%��C���D�"l��h���Kӭ��m��k�q�L�f�D�ʻTX~��}WÂ"z3R%��ŷ��4aDxzRʥ��M���[qɲ��JQ��;:ͶithMUz�ꐽ8�M�q��t��S����v|�M�㭾uכy��hMa��,}��[�3��z�7�����C%|ㅘ��\�Ũ'1�,���2 yL$�[�����qD��\��U"����fω$�EΩv�-s�3A���\�(g,"D"��N��wq�K��JA�'q�Pu�l�`lfi8!���]��� �R�ӯ��,;4'FP�mn�m���\|�;�g�J�xh�&�D�=�=ܶ1�٧��tu�syuuټ[[0��e���D��8��"Ի5Yg=�ۭf��l�{މ��N�&C�≳�s��.e���J6ː����I��v!�kb�.4�+�ӭ6㭼�6�O:���zl��ӆ�i��ʩ\���U��GFJx&��3�ϋ����&���߈,����:3��HM�>m�f������3O��0�1H�m�|�p�l�"���g�y�#���1A|H��(jc�RNb�*NmզSg�=)�5�~��\��>B��4%� �f��<(x&������L5\f3K,��u��y�m�0L�,K!�8tN	�GQ��D�Q���:"X�"o$�Ǐ8`x��x�:'N$ât�F�R"pDD��%&�P��N	�6a�D���D�QM��f�h�`�?$���B%��'D�D�%�bl��<Y�ǄO	�,L,��0L,K��b&�:'N"A6"p�,��&tC�H �lM�P �P�&�fɬ+�T�9_[[�v-U>�����cY;��}Ƙ��-�R��{1�z�wFla&����&.��|^��>��{J;z��w���W3Cu�k�\ޚ{�Շ<~��Q��yw��
g��L���z��-T8M-����Z�F��iE�RR<H}={�<��w=���g�<�u�Q\�m��ɜ��K\5���;�:i��Y�C����ёΦ@�li�;�"�ҽ�����
>_h�{��fjj���3��{�����������u���������{���߯����{�n����{�<��8��6���<��㌸�ͻi$��6�^斴��|���'D�2N�}~��4y���ga���z&��Y�t؏�-�K0���P�R!�fj�\���$B��,�~�?-���C�DOޔ���D�j��Q�{�2������a��a���'_:_z�0uNG������]�ZMS���o<��6���<��㌸�ͭ���cd֐~/	�pA�gI$�C��L��|"�rt���x%2�__�����B+I �esDH��I
	�3���'����ؘe55�̹��*�.lD�_�Hn��Ȗ4'�����ihq�A�V���ͻt�-��5�M"9��^�QFj�y��k���k/�ɐ�S�<����L�?�%�&	g��g�<&�ц0O��Ғ��F��h�xx�!R�A�!,G-(�o"}R���cl�EHyT�:��6�)1����zQ�M*��s�T:�qZ�u��j��ΒI< ���1-$�8چ'�h+�B�ET^�=��Ņ��-wN{5�v��Oo+���ֻawh���ȵO�$�����|s�W��M��חj���2�0ˮ��[���+#��Y�v�^���"4��uL(��.ѳ�0�FÐ�p�h�V�i�&��V�u��ASa�S�^�����1ījʹj���E�/'�L4zƠ6i�]c�#˱M>m��<��[y�[y�uwWq�\u��=5�m�43���%b��Xkf���!�)���kw������!�AI5{��ZE�����N���}�&���0N���m����FhU>>2�AD�{�e
l.�:ߪ��$&F�޴�4�������&-R7L2���uw1y���e�Z���lɗ�,��<�n:��]m�y��]�q֎�HyJ����F�"��7r�2�y��D�},]��KS4�ZD{Z�⤽.�=M5ՖgT���=�IL@�DB�)[I�O���9�m�h|9�f̜;��;~���s�M4%���rha��L�ږ~��~9N�<�hN��'M��'��$��G���e�|�>q�[y�^ywWq�\u���ON-m�gɖp��M���n�I< �:y�oA�0pM磂o�8';�s0k5�ѻ��]�Ӭ�,���?v)���y8���`���S�y5��p��]�f���lO!��5����'��~Ӌ#��,�n���*=_g�:�/M���aY�0�%�b�L1��Y���{}�JY�]�|���:�o<��.��8ˎ����o�75��O.��a��'Ru��vAU �&�b"�h�5PեH� �m��K�9�ĹM��zÒ�"V!]����u�a�<oBuɍ���I�sĒO"�t�>�VLG�j2���3/�����<g&n̕�/[o�+U{f'K�u��a#ܽ��%�^�8aӰCg����xy.9r���C�e���iu��;)h���1�+�$N�[=����AÛ�3.2��k������Sӕ�f�_�7NSf)�|��%�<���0��3��:a�ȝ���fT��8p����0��<x��Ƅц0N�+&T��5��UQ��5�*�a�������բZ~�ԟ�����ѝ�+�A��K��f��^��-dS����;�{�:<p��e"�)8��jh�^��٥���Rq��G[Ε)��絾�Ă���"\Ħ�&�g�ל'd&�����4ۏ:��\m�y��]�q֞[X���^���P�H� ���`���-C-�����h�u��j��j��k�Q.�e��2j�a�nO���К�i�O4a��Z$�hv!�wR�#���h�K%2���RI���^����+�L�:�'��qd2�j�G�+\��"Zd�+ӋUycfR�O��$��%.�i�e�u�]q��a�uwe�Zy1�.��i0ZD�����H|E�����4�]g �|�(ܲq��e�Nv�Z����{>��f1Vk���lv&Kc4��	��2��C����CP�M�f9�=�u�c��5�=�ʻ��w��۩�r{U�v�r'_R�$�������5�kQ��CfA��(���ʼ�~����	?�?�?�"(��X����!"�������'�97O���_;��M�1��M8ꪩ7��hɽf�~'Md,I�3@x�X���� �BQ	HD%B�� ��A	P�BR�JB*�ы��0���`�&��,2��0Ɇ2��a��&0ņF!!*�J�!	T�0����ba��,2�b�&a��ba��&0��&�d���R)�BR	HTB!*���JAJB��R��BR	H*UA*�)��"�!	HD% ��"��	HB���B�J�ABB��!*��*!��!�T!�*�B%!*�JD!)�b"1 ��"1 ��dD�DDb$F"$�`��$F����A��0FAdD�ĂD`����� �	� ��D`#A �D���H�AD��H�%"��A��"DdDH"2"�FDdD��F	�Ȉ##"$A�$`���ED�A���A� �� ��A"#DH"FD"#D`�� �`���"2 ă"0DF"#AF	"#A"#""0DF��I"#"���� �b �`�� $"0D�#""2$�D��#	`"Ȉ�`�#��@D��D� #H#DdDH0D$D������ȐD`�"#""0� ����`�D`�#" ���1F	F�$`�#""0H""2"1#"0D���0F"0DD�@�
1�$F �A �A��"1DH1 Ȉ#A##DA"ȃ"A� ��Ȉ#" � Ȍ"�#H�D�"$FD@F�� ��@F0D��D��@FA�AdD�2"D�##" ���#"$HA��ȉ��A"2"A"Db$FD`#��DFDdD�"0"A�$F��� ��DD`����`"2$ �UQ(�DA�A�"2# �ȉ�0� ���0D� �Ȉ#"2"#	�# �"2"�FD4�T`�R1��i�aYaX��ɅkM*Ʌcd�4�h����ac
Ʌc
ɉcX,�cVX�b�cVLG兦0�`1�e��FWXzaJ01Z�0A���"�����!)��Z�J����B�JA��^�0@b�"�
������T%/b�]P��DDD�HYU!J!��BR��ؼ!(�!)�BTAdAT��A�`�0A`�D%�PD� Ȃ �s��,BT ����� �A�D2$�!	HD+vX�P�%T"�JB*�P��!�B��JB!*�P�BR	U��!	HB*��%!JB�!)
�%T!	UB���")��aj,J�EBQBUB J�T%H�A��"D�D%!�D"��%%1*�Au!)�JB!)BRP�B�	D"	UBT"���A�T"��J� JB!*���B!*	HBD��D%BT�"��B,2���&�����P�BQ�JB*��L1a�0�a�0�+�JB���"�A��$A�!AdA!*�BUB�-B�!��ea��L1a��" ȂDDA�JAJB!*�*���B��J!JA	UB� �JA
�!)�JB!�A)BUB!)AJB���	!)A*�J@�B��% � � A�� ��*BTH����!
�	HB��% �%!T���"	HD% D%BUA)��!	HT!�P�J�!��!)
�HB��%A
�!*�"�DHD%T"D ȄD	`��JBJ�B�T!B����B��n!*P��!)BUB! �A �	DDDA��" ȃDB1A�b	!JB�HB�� �A�DA�A�A�A!��������Xb�Ɇ2a��0�+�20��ņL1a�ea�Xe0�+`��"HD%!t!)BR����!	HB)��B��A	HB�D��J�A*P%!��R	P�P��HD%A�P�D%!�dA"ADA`��0�a�&�1�LB2 �1`� �R�b�B	U��"�*�P��B��%B2 ȃ��A���!	P�%T*�JB ���J���J�A)BT"�%!��A*	P�HD%A���D	D"��BT"HTA*	P�%A��EBR	HB	HD%B�HD �T% �JB��B�JB�A)�ԁ"��_���i���fu\6NE�i8Z����<�B���%3��2�o�N���v~�\>�.=�7��;�7�����i�w�g{���nc�·Է,6��71��վ4�����^�Nu4�/ï~���}wb��n�x�7;Zis7׮g��_v��:��w�=��á�)J_zu��K_)|��b~{+����L9U�%)~3X��2Yh����3s���yQ��p/�2iMW������1]s��{/�e��1�Ǳ'���ĥ,==����y�a�a�4w���z�i'��o/�vV�ɵ��9'��d���N/��բכ�.Q��*x��߮���ڷ���e�c,���z�>Ʀ�F(���6��H��m�T�r#vU.���v*#l�)��[�����C'�9��U�~���on-뫢?��uu��tĂ�aūD,�T�1�L�B3i�*�V��f���r=K��X����w���]�L2�q��.�躇8��a���G�9������?�����������Z,ql;,����?rq�uo��ޑŃ���.Hꜭ�ӽ�`��py/C���g�8bn^���������y���_���{��t��TJR�FT�Ί����>��������澣���MS�j�᪡R�8=�)K�<W�&U�g���X�l�6ڞV���|�Gj�W>N�fp�&���פP[���{���l�m$���$%�aa��p�j[���l�⹛��54�~٨Ҽ�Q�7���WJ�0��?b�J�.�r�MC�}k�T��8?#�S��<�J�xD�.�o��_;a��i]v�G����9��s7t���t��N���g�z���^����e�V��i�KK�%�/'d�&┥��:�~��|^�E^���ļ\3Ǔ�?5�g��Gl�;�ju)�\�w��I��9L奧%2a����[��ݙ�74i�u�U�������1=��{z�FS�m���zl�6�8t����nY�>�)��%)b�,�Wb�x[�Y��O$�vb�V����V�.忑{;Χ;���,9�G�Ɯx7�4[�ٗK�~�Ȯ���w�1$�,��פl;�����?oÊ�;N�4�]�j�:ףӪ��p�Z/#��������k�3,|sF��aa].�r��o���"�(H6�	*�