BZh91AY&SYA(�(�߀`q���"� ����bK�               �	BIR"������
TU�P*���J$UQR�� �$P�HH��*��5���T)�})��
N�E5��iE�
�T
�F�RJ�!%V�TT��%U*A�4�H��يl�EJ/��Z�"Dh�R���^�f��. ιP����p uCF����9�V�RZ�k�Yʔl����hJ�7 ��e-5��T������(��JE�ꔄ��`(P��@�=�n�[9��mZ���KU��g_Yz��<^o{�n[��ƪ�����9u�3���ڶ�mgz۷��zi���sWB�K�!m��kcR$Q��)Jm� ^v>��UG>�� z�R�<��T"(QNu�T�)H9��mB��;����UB*n{;}�U*�I�V��OcJU^��ｰ�J�N�=QR�9�T*����D���\J����� 73�}T�T}�W�� ��T�w��l�T��ꔪ�J=�>}��T
��7���묻i%R�y纅P�=�����%U�Sݭ}���T�B����UP�O�T�
)�E���S���)A��s�R����N9�{5R����3>}��U)U^�٪�ډ��}�J�U:N΃�5T����>�UP����B��N��*�QR�׷���U*�^%D*"AP���*R�(�gy�U(}2��v��R�Hǯ=�UB�e<��;���������QR��t���U�U*���R��ޛף�[R���f�}�*���׽�T���URU	P#ehJ%��RT���� U_o{޷�*�RT�{3�*���p�� w���7�qJ���g���������v�:项;���8`�UTTUUP�� }+픥 w����k[kt}�w��i
49�� �S�t�t����N����^��Rʠ�=�)S��Y�T J���hҔϕO@���h�[�� w��x�<��+�q�s׶ 9{��4Dj�CM��h��u t�T���(JD�{�R� w��>�#��@V��݀8�wM{�U �k�Z�n�p(.�ᯠ��<���� �s���QT-��U��������rH g'��P;ce`�:s�J� �˒:d7)y��+� :�w
�bC�w6�*]�   �     S �J�� �  O�F$�E@� 	��& S�A)UM�M  b  1$�PF  A�	� <�@�UO�&A�@ 4 �Hz��*$��=��C���z�$y'�s����?���v���,A�� �	�&�s��yL��[��ΫhCs�.}[��|��
"
�λ�����
�  ���PAW�@������qS������ʪ���U���%O��_?��/�y���v�������1�c�c�c�1��1��x�8�lc��c�3�1�c8�3��8�7�q�d�|c1���1�ǌ��3�cx��1�c�cƛ�q�c�q�cǷ�3���1��8�1��3���1���1��c1�����1��3�1��8��<1�g�ǆ3�8�1�c1���3�c�1���c�q�c�1�g�;q���3�c�1�c�c�1�g�q�c��c�1�c�q�c��c�1�x�1��1ۏc��c�q�c���1�<&|g�1�ፌ�=����1��cc1�g�q�cǧ�3�c=����1����1��8�1�c8���1�c�1�c�1�li�g�1�c�1�63��ǌ��1��8���3�c�3���8��1��1�c�1�glc�1�c�q�lg�q�1�c��og�q�g1�c�1��1�c���1�c8���8�3���1��M�c�3�c8�63�c��������3�c<qፌǌ��1�cx���1�c�q�g���8�1�8�3�c8Ǎ�q�c�q�i�gq�c�1�c1�c�g�1�a2�SSS�*c � ��8�8ȸʘʘ�8�8�����T�T�Q�A�q�q�q�q�;`�Q��q�1�1�q�q�q�1�1��)�)����#��
c�"c�!����A��A���D�T�A���20�2&2�	�)���#�����0GSSG��(�
� �"2.2�2222x���<`aLaL```\dd\`x�02'S�A��A���C���D��A��ƙSGSG��Ș�8���>0)�)�	�������)����8�8�8ʸʘ���8���0�0SSW �D��Y����T��A�P�P�A�Q�G�GSC�T���E�A���P�1�q�q�1�1�1�1�dLdL`L`�D� �(�
c
c*cc
c*c(c'L�02�0l��#���	��������¸¸ȸ�0.00���ad\e&S�S�D��E�A�T�q�:eLa`eLdLaLdLbeLd`dL``LdLdaLaLa;dq�1�:eLa`LdeL`aLacGGGGS�q�q�zaSG_Ld^22�2�20�0.2�22�`e\`\dLaC��T��T��Q���U�A��鱅q�q��GGG��1�q��W0�0�0�1� � ��L(c�§1�Ld�@<ed\`8�8�2.22/�(c̆0�������������CG�<eG��20�2�2�+�#����l���c(��8�8���8�8¸Ì�2�22.0.0.00�2.0q�g�|`�q�1��0c���8������8�3�t�3�x�ό1�c8�1�1��3��8�4��0c�3��8�3�oc�`�1�c��q��1�`�1�g�g8�0c8�2c3�d�g1ǌ�3���1��8��c�g�q���=1��3�c8�8�1�c8�1��1��1�c�g�;`Ƿ�3�t�1������g�q��q�L`�`�q�c�8�1��3�`���8�3�c8��8�3��2c�1�v���g�q�`�0g�`�c1�d�`�c��8���8�0c�`Ƙ�q�c1�c�c�|q��c�c�1��:q��lc8�3�c��c�M��8�l�3��8��c�7L����&0c0c&7����1�`�1�i���1�g1�d�:q�cl���c8�61�c�1�q��1�Og1���g�q���g1��cg1�g�`�q�1����������`�1�1�n3�������32�	��=�1�g�q�c�q�c��3�c8�1�1�c8�1�c8�1�����8�1��1�c�g�¸���#�R��6iZ\)m6K����)T�9g2�J�T0	k-c�2V���ʻuNG{Wt���+R�#[l��CH��uiͰe,`�bݴZz��e�����ɉɣ�6����Ӂ�O5�Pn5n�3%�LC��Y���N���M�YAn��Q�n��շ���5(^��e�\6��R�M����]��-^��@z��̫���f#� &輂�J��qQoc�VU
��m���n)'�i�JK�R
X�$x�ͧ&T-��h,�`4-�
�
�n:�a��%YVk��������j���ݻ��o��Dh���=۰�����Le�v��U�Қ���س�"�	r-h�G�t0^P#Y[Yh����PCw�����+���l*�QX�ۗ/
�t.kYyJ��&�4Eq��Ы��9/����yi6���Ӽ;i����;j����$�A<�ƈ�
^�iZ:ý� ��G#�f�4��m���*�9 p���dA4�K�F�)�$��J�ϴcƂrl�B��Qɚ�����-�EC���D��-%	u����SD	�J!N�l)m��0�2X$� �NY,U��`1�����.F,Q�ȩH���̕pҥ+a�A�k2V��RA�ʼ'���yuƕ�Р[e���2��:�S�9�t):��j�K+d7`*{I�6�DPi�sY�$˥DV64հ!�W�d�1�v})]9�n�n6m�á����������#tY��7�^mg�݇q��ٔHsU)��-=.�ҚRk�����Zؑ�A�B��t�P�`�Ub���@-���+�����`�O�.�jQ���j[�q�l�de�ڃ�I�]�J���("�0�v�ڳg_�dZ�˵�� �YDSx+]c9F`m�P��RaǴ\Y�g.|3mլ�V��Dڛr����{��ط�#Jt{C[����A<��ү%<��X�D7�+~:�[���X��2���u���̵F1�F�m9x	�kP��+��	�)�G]ڱb�"�Ix��=���:� ������L^�Z�z�{���,-t�a�W�JL׮d�ک(k�1a7a�����+2�/h5�CǗD��Um���WI�7�Լ�e�JcG/RjYL�k�̲.i"Ri#��^�ݐe��1pÑϔ�!�ybU��n�C&Y��A�0]�/O���#��C#"�E{QLt�U{s-)Ia�;�L)��u�JY3�X�t��iP�b�R�RbGc��^�����53nJ����}s0�ɊӺid�
��b��U����-�L��d*
ےc]����b6�419Y��K�1�>6,�ߦEn���NUەy�N��5�-��f��qYp ǧ�d�9cj��X�fzL�f�[��� X�x���T��X�<�2���D��eeX�`ID[�����#0^*�Y����X�� �����f*l�U�k4�_d��S�Y��Ʊ5����,!E̸ �CEYi\c^��4�A[Y����M�6�ӕ�Y4�6Jcd%<k���cnT�L�cW"�mՋT4L��f���&:9{�n���q7q��J��i��S�ĻBc��2�YU� SX��hoeV�F�"S��K�IİX�t�U�qV6eQ�;4!ˬ�znӖ#��ۅ���I����ۼ��F�كM��`�J&kH�+�����C6V� ;L�W�SQ�]нl�.\@�8�(��#˧�/jt����l%m�"��wKN�Te�V�)L���Oα��j0�W�3$�b��+pU���4�4����Cv�Ţ�­��ai+--�����2�&LOL�����A�2��pRp*�mѧtl��b iՕ�s2B�j���IYN���9O+aUGF�aJ�Zs���-�OT�L�]�G�V���SU�l���^���jZh-!���M��+q9@�[Yg�8#r�̖��U�MV@�U��X�݄��fZYt񪆚	35�>�t�1��L:��J��,��36�0�i<@�%�I�4��%,[IfmiZ�Jwt�0̚����D2ݥ&��CږY���W6F��5��`ںD� YQ��������5veFZN��2qԅ���C"�%PS/S�,jԩ�������6��4�l�F�|�rG:7w@}��	�R歷|�]��}FI/��T�%b9� ��"�>�����XF���N��&(�if���c�mnS��5�j[�lJ�F�C7L�;K��Yw2��p�/Ȗac Vs��X3I&�\Ў��oyF ��ѧr^�Q���=���Y�5l�p�׉�R�d�%c���Ŷ٫-P�N-6(\�* `!,�I���KS���ɔ��ܖ���Z��nS{�S�q(l8i[�Ԗ�4��k�D�!�+Z �έ�f>؜yK��X-a�Nխ�5�5�֚pB���NTy �@(� �5)�ɹzs[���;CM	�![Z�[�U&K�4a^��D�Sv�r�y2���n�k-����k��-:j��F!�+r� �(�[+sKK;��5�JYu�����Pj�VeGVۤ6����2&l ��-�Ʈ�l^�lU9rf*n�lUp//2,:�Zxc��Z)�lk�91J��n��*�/wY�cd��A���a|�A���q��Z�ں�6D�*�&%��Jn7��{{Sl�f}
��i��VN��Bc (z�2�lQ[�%�LQ�Dֆ�.��U�`�d�J���՛��V,� ��f�n�@�R�Q�e`b�Lr����\&�#p?��&�iPt�3z-�Qɭ�Г���e��&�Ù�e���-/��{	(+f�ID[;b�
�D�G4ѫ{����s#
��ou)��M4�9X��P5L�4�E]���*�e��4G[��9����i坛r�J�YN�(9�%6�V7Rj7�wm��"h��A]EG)�-��0%8�Vӡ��3)fՌ�v�:1:�j�]չ�D���dƯu5e��� �p�)e,N�6*eM��%
�ѿ�H5N�U�r�\Q�Ռ�B��j����7�dݸ�Xfn�iԼ�2;�-�����ԥ�G�̩t�T��1x����e�?=�.�B��"��q�H͘�*+QgN�<t�N;�2���&����졷�1J+*bu�2.��p<$f\���V�A��>˴e�^hƋJ=ݦ�w�Bom%o��PJ���E���X�PV-�H��a�k(\2+]�<u�rٻ%Y�����6�8Ѽʊ�U�ښ�yz���r/���&˶2�kd/��@س�f܇U2ˆ��wp��V��T��4��OA�.Q���H�1eX���פ�ZZ9��j�TĎ��o��ٲ�T�7j��uL���J�ͺ�6�{s4�+3�%TZ¥�^MڛyM�p-j��y16���P��.��pDQ��	��4JY"�4�T���N��0/؛#��c�ͽ4�$��#(f�9�L�" �,�����jb�Ȅ��>x�ٌ�sth�y�%V�����N��.`{�t��G�CA(����Ԭ�%Y�Z�+�PP�Kw4���<d	�;@<j��\��5��!��՛lapi�iU��Ҵ�f�Kn� T0��)Xg0�tSA�f��@��/c6]��&�]�n��@5o73@Eh 
⭍/��"	S�F���Yu���f�D��`Z��^�r���U)Fґ�[e�` 0>�h)�%�I=(���w�/]C �%��
H7�F�F�5���n���{�C�`��3�N��acT��I��
T ��*X�霵knؚ����E5=��D8C�+%X�2L��U��ck3��\�f�86I���pn4o-Se���-���[46�j�j����ݥ&)�Y��`�Vf
@Rp�,��8��,�������46Y�Up#շ��Z	��svV!$d��h�
+	
nT;xˬ$S��G5;5���S�.,�Gif$�:����vrЬ�&�:u/�R�9��EF��
�X�c����G��LjՇe�ˋ+J�71�U*lL֯-%�UK��l=�mEo5aϯp�R��WR���3j;Y�Kݗrk�\q�eD�w6�
���Nء�a4c�]�7pq%Ӻ�[y����͸�M�jPBш0���ʉ]f��FR͊nM͂�5(]nS T�F����7uI6�ж`Y4���:��vխ��KU$�4��n�%q�V�uG2�&�GK�%*,{�^�8�Iu��uJȷ+i��r`v�,Y�EDI��Y�.���rX����?Lo �UѮ�hRI�-�k	��l[�7���䭋(	�hN��0��
ܑ��b�9u�(�m�[ge+��c����.ɬy�٧򔴊�V��
d��Λ�q��a\+([���/���ғ�umѥ�:�(��ιS�r��ٸ�����G��gu�ҕZ���dM ����,X�i�LHEDVB�&�{Dݽ��E��cZ��n|�lXn^@�2�T��K+Lj��.��nXu���3����V֙�a��`��h�.�йIC0�0X�a��u��耿����4#djX�U�"�[�n���kb��\ҍ͚Txf}��W��(��%��OR�����U����f�@��f/��؊�niz�E��S]�ǰ�N:�b��*��MaMɀ�I�oPEjZ􊐂��fP��D�[�n^�ŕVi�����6b�n�E1�Z�
���͢M�Q3n��U'��mIAڒ���a�^�DƚoI�\��|��L[	�
��sV溂���n�yxַ�Ò��<�$+U$K��;x)�t֠j�P`�s`�3F�L 2��[���}o0^V�Z׫*��)R���.�b�Wn��[y)��]���Kx��t*��-��wu�jI�0H٘(@#��*�S尒����)��>����U��v��l�d��rDi
�(��j��7����m��ک��	�0�ə{{�9/����ۻC��Y� �Ttj��BmAL�qݒ�+T�fc�[f�eW�cjV�����2\�-5j1M�N��k/X�a�ŭ�b�ы��*c
-;C�b���I�в�;�
Ф�ڲ���[O2Qm|D2�f���3��"�hl��#r4�1!��[�nٺ�+ �Z�kS8`{����Ѣ�H�jb�b���e?�n�R4i�8P׸T�!�m�r�t[928�m퉵2'��g����/i��*����F����DT�Q�V�s��9�o�.1/A�/�=��N2�����\���
�!�9�Eh>�N�ĒH�fM��5�q��;�������>^r���<����FJF"�ò��wg��QR�>}���{<�������LW�&�/�Kҽ^ݿ������/;���{�%A.������B��u�����ԭ�a����r�����r�[�*SZ{3�Eq���������밮��wO֨�k]��U�1�=����Kj�n�"����Z$*���wy<L�]p��~�|��ͩ���K�%��n�\�9+���B��c��'[�C�:�Y����]���Y��jV�7s2�nY�@�Y��u
��d��Et�J��|ﯪ:v��^��5�`*y#�5|j���ќ�yQ]�6�3������,�����/k��Z�&��/�-[;���d�����V(���E�t��S��n��������"n��ݽ@=��S2�1�!#��N�.�f�t̓����jS�6ЮŪ�� ���y�y�����#�W.Ǚ���z�Y�w<:��|o��u����!#]a��^c㲭�d�o�B�\{V;��6�o�]o+;_�,��U�]�}*��:^,�6nև.�FI���^\��v��L���#�w�A��E7�j/%���z�d(��Ü�nB`��,H��DC�3��섽�цtm\��n�kNF�tE�w�l��N�v	�%0�u�O����bi�y�)]����P\�,�7&.B�iE�/������i�L�H���Ĳ��B`Yf>#}p��ۖ���x_Xju�Q[M�	��2���<8��p�ZV���i�Eaowa ��t�������աݞ���4&�ٷ�Z�{{�m�����j򕭴u9��9ɂ�4���	4(���bx�✤0�XF���߽~SԨ�$�����8�!~�@�oK.��٬�o3T4r�ް��7�i�p'{i�*H��;vlj��>}�x�n�i��"�s7\-\Ρ,l4l��l�$��Sm1�Mou��c���L�o��Fn�_d�|�"�8��a��~y~�y?!�P7Y��҅�V��aj�mP�r���Rzg��t=�R�\%�^�g��⩶+=�l�N��t�&L ����y�\hvK�a[C�ڧ�y��G��Bsau��:��x*;��B+��L���N���UБW�$w�+Z4d�����\���w�܍� ��yTOv��z�y`k���;�L:�6��{;���%іrגM��N+��{e��"�$��V6M����z�������V(�8I/��W���?�|�Z�܆��@�i�m�f�����u��^��",ˈ��3��oZh�d����2�r�'^ߓ�ni���G�ul�sv*w��](�J�g���]�p\vy_�dWڟXmP��q��<=��kdw�V�R��2슂�h˴�;5�_�U+�6v���P�Ne����k��r�ߵ�g��_P��������g�t�
տ��[�����뒲�;
�_("���뭚�>�{��ē%�$v��
�e���W�*pOi߽���uf��m��m�S��W�z���L��L�(F�}z9P��5�j��J�ȝn��S�'j�n��M�������r��׬rnϰR�RX'�epk*��x�X���B�ʖ�h�>��O����V�{���ٞ�~N��t(W��,���y�8i�Xx�Yٲ��3��5}яzj혦.� 0�Gl-��d�]�9�l"6Y{��^��G����Xfe�o~���!�OxP��{���/���g7?���J3��dv�<Y[m�}P6N��Ә�eL�b�,ã7����͆^YZ9%��;�˛��ʾ�V���+���#WӺ,w��Z�`Ty<Z��ה��ju����j���NVq��<����wEf��s�.��O6�p��7b%VR��ݼ|i�}�l��xn]�&���Ղ%g�;�cSrSU�ǐ�@J���5��7B�6��zC��]Z�S�������1��9�.y�},[�N$�NFZ�V�i+t�ut8ٻZS��f�,�u�_p&7ͥ��a������Q�Iѓ��YЍCy/�j+�|�.���䤰>��d����p�J�,.�y����Q��`�}�k��ȩ�6q��w�W��c�%5+��ޕ����Z�Tm��Z�����7��Ֆmg�1�OA�ةt�,u�5��	t� �κ�3���1�6ӻ�U���P��S�> ���X-q�2PN�:�ͧ{��'5�[��j}��&�9Ʈ�[ȸ�Z�8"n#u�O�t�s�v�y�.����v��T���[�,G�Sg�1�[�u������e��9�������*���Gs%��rZB�(��l:�F�nJȁUyb�f�0��|WV�F	�٠�~.�����a7bu'�_S��f�ΰΟeK�C+~��fжjD�^D�MJ��^������왅JF�<��w6T�M��.��ʙ[I��n�w�gP0�@;F�ݽ��x:��nZ�tٺ�h�В�i�+�^�|(���z�`�"� 	�y[/V����n�Fu����M�'N�[������h�';����7��w`{���d7����Nw=(��JRh��B��ok�KUt��(�1َ��Y�Wg����9pT��
�	ӄ�5�Xs�r߉9�'�k�ڹk��v�"Rs�g�n�Y]u���¶>�娚��f�ܬu��X���c'�αp���v�\PԳV2�2v2,��a�a�#r�A7N��i8F[��_��kK/Aw��ꌩ�suE0�XV� 9 ����R���v<}�fH�TX��;���C��p�:�ѯ7��lM/]��r1�n�R?^GB���;���Y5�v0���-��z�����Zb���()��rwF��]@�a�7u�nXAo#������&�'^ж3V����� ^���;B�4�׵�uDk/�4��(�)5[˱���o-Ř�J]R+�xAx�W�:��i�؛�0S�4��X))O��L�
��f�r8�ѕ��u%Np4ڬ�w�@�6eu=��1{��x;��d��nRF��#0\��Zf��?!B�d}n����=0ড়e:z��w�8� ����Ъ�:�c����u���gB��0PQ@�K�f:�BoA�Q��{�:�RJ���1��H����ѣb݀���io��WT-���rb�)WT�:�ʾ�����M��"?�����O��i\��������ܦS�z��w.1_���A�Ҙ�=��oJY��#Ye�n|�+q���K�����. >�n�פ"�]Y5�G8Փ����[d������@І���Ύ�B�u	'ʄs����NK���j�*r/�n�(Y��E'uvl�bͮ=Ώү7� :��@��M.�8�Ku�sQޟ
G��u1�����!����;�e�F�������ɢ�V,���Rړ�� �����V��V*�co#�f���,Պs	,V�73B���;|9�r䌜a��ٓ.=�ofӸ�! uf�j��4oX�n��쭵!F��R38(fh��㣀,X�}s#���]2��oK┐�����gI<��g9O�������jT��6��bg3�h'�4Y�쮈�i�]oG�&��ևQ`-�T��h|��������%L�L`C�1�PWQ�7R�dV�lo�F�i��TFTIc�Cx8(���+!H�d(�s����ki#y�g��V-j'9Ҥ�ʌ�}4�f�5�tm����^�z��Ȧ��eZ���s�#����Jq����(I/Ec�u^yo������2�`��mlӕzө���r���[\���:�&ʥ՛iL���Nf�T���X�i|5q �6_w����K�=W�4յ���Q��vm�c�w�����D�2�u̜��e�8r&=����HvT����%v�!���`�o��᧧p�)�7̊�S�"��d��O��Gt��,����ǅ�ꋥ�۸�f�g;Y95v���po�u�BF�t���,|�h��wJgY<���7��l]�DVCh��zJ[��' ��z��]D�[���D��o-N�ޞ��ijuz2�]z�&ms�^;��Y�sʶ�H�������b�.z�Qdic~fi�EALqk�Rm*U:��Y/Ӹ*�*GuNdiޛH���V�'E�([̕,��O_�`����ko"�$&7�m
�\�7���F��7����W��hu�A�"KM����f`�V)ݫ9e%/D���	N�Yy":�]ua`Ð9v໊�w'2�n�Ļ�-!9��/8�;
��Wu\U��V�u�����b��'�2��X�+�ݴ��b�Xv�<�5�d �OCy�N!�\�|�勋-��,�Fk(�[�ٸ�k�#Hv�<��7�
�a�<n�x�q����=�V��g"���� &��/i��oܖ�W�'(a�������뮓��`��ժqڂ�;�������� �u�.�>wx�R�"�k5�Bz6�	{g�vo���X��SBMcgS���-Y{]�P�Ǒ��
� �7+�䣭��%9GR�F�a���_]�t4�.�����7�7j���M�J��T��Q3���nM�//;q�q��Y�D������j�ԴG
�$Z8Ud��6Q����1B,�H�ǃ���ר�5ȥԺo�0���c�L��s�ZEs��Zw������ҹ[�%I�}���$�LJ.�#x��^��q�k���])MGp��i%�q� ΰ�5���ٻ7m������-t-]#�͌M��9���gw*�el�ܢ-�.s�=O��`с*��-`諗)5�Cϙt��G.�e\A�m>�b�Yc����L��I]:ηi�+4{�D�O�y�଼���o)�X�E#ō��qde/(Z&r�\��B�[�f�I��w��4����`ɤ���t��;����wA�k�P�T�늷�Z�Iv��-pԧ+Z�ҵѝ|�Gć�6��k�Â�s,Vm#����ۣ�p�ΊmR�_0�g*F�M�aڔGe@/���%��\�m�75��	�8��Η�oZpŗ�T��q�ǚ�����J�Vn�X�n���
.!�okИ��@3���w��R�������1���Mͦ�;BjA��a�·�p �)һ�iqɕ�p�In��;�[׎�.SO8�/�MV�W��G�R[�.���cRX����E�@�g4��b��ئ7E��wo~�vr��2��y�׎Mk����V4)�-Iܶ�]�
]��_alo����d��e-��k�2�q�2H��ЁoV�H*�Z[�<юĈӆ�����"�u@��f�g�N���tE�^E��t>��n�]�5�����L�s�
SF�pѭ(Z��ݳ6�p&Д��z=���cNsOn�t�/f-,�����]0�H��XU��][%���d�t�����!e�H[�V�O��1I����1f�Tr^-�iZ���Q�z-}b�{7�A�Eh�s�F-�.��\���t�9+��0e�F��Z�n����9,Ou�U�Iή.����ŗ�a��D�d���Es�b,��r��7,��Ớኁ}�w`���IK^�c"���*B�)��ޮ��9��Fɗ�<x,ؤ�$�8Mi홃�,m�~'�t�:��մ>e<�ŘΗ}ϡ��lA#�6�2�k�e�v�s�Ǡ�f�p`'�b��^Th��j+�/u�����}��A9|by��8R��S��Q��*/|Z`���+E��٬�Ib��e�o��Iq{�*!��H3�c{�k��j�n)��"K\�����cC�9�@;(U�iiTsn>鬄�����ʋ`�����i��wRS����V<ɺf�ވ|/��S�y��@����a:Y���\�1�cn^�/����:����'3:pN/��[��ʳ�P��3��5|���r��X�
����,+<Vz tF�"�<ܫ�
�������p��
�Q1�G�gu+��׷kHjH��ȑ+����2�f�9��J3��x�K�}��ޅ6��g3:�ˎv�ڑe_k��t��n8@�ݖ��mY���d3\�6�cӚ{��S:�̓�,yP�5o-2�,:N�JH^�fr�Dֽ�L��㢇k�������]g����:o�,�Рh��6�V޾wk�5ە���3�a�\�\��#{��Mq]��Toq,������1�ɵ���n��ɼ�kN�x�=/M1�,��9��Z^l�O�Z�����W]B�g%I�v�㎜�<����_R���q�*��]+N�H��Y�]�t.�6�J�)v�*2��]E��E�.�_.�Th����1tі�B^V�Zq���!��%���{�D��_n]��o�Wұ�f�}��q����jŵ�8���,:�J6⻭�a�b��qi�]�p��,�X��I�e�׭$$���яv�@���u�(���՝��h`c����n1����(�)��a�j"&�(����R�fo���[�*%zI\�����!�}��b����<w�۫W&ڄ�{�B;yԈ�����ChT���[;&s;'o<lCsl^!ӹ��SQ��a(;h��с�쬱Z.���D�U�Z�|o��q��T�9]׳���i��M��f���Od� (M�1��l��v�m�cyv��pO�ɽ䡙[ĢX�}Նq�֮f�-��ue]��n.=�t������է���J��w��m!���(L-W=��b��u�p�A۠y\��VgE}Q]����ܥ��Vtt�ǣW&�-��텍��@��J7��_oNnk���H�ʀY��z��9IQ�N����c��\����.9��imƷ�����e��`���,�Q���q�L�=�S��Â�9�5�GE�{J��.Z�
Vh��,�A_:�������}�&�q��p���*ES�t9�:�Nc�C.��r�����gL��ڧ;�mB;m@�A3���.�&p���e��Ծq��u�*>ק�m�uu,�p���54��(���3�{������eXF��Q�(�m)5���K��z�y�������\�m���]v�Lb���k�Bh0]�Ee3Ә$�MSEFͼU
V�(��.�B\��Ԥ)*���6�][yF��M�"�!U����4��!�+v����:��At�]�k�_{��!;�ot�.�t�.n��ɚ��7�H��E�,c�S��D*�[�Zp�/)R��E�J�L*	��AX͹�JLU�@��� I1:��I�t� m:fP�A���*��]*4d�-��	�B�B�&�)��h����i���t�
r�,{���w^�v��ַ7n�n�}�l�
kGh:>qQI�)�!�I ��dh��(VB�e�#+Hm�ˎ}3t��UCہV�	�n��IEd��+V�*u�1��ݿg7`�p��<�yͰjF�x�f�c-).��sc5_
4�WчG�&�]�38'*Qh�O�tˎPu
xq���paITn�]�+t�E*%���$�L�WX>yQRJ: ��A�|�
l�ҒO�j�A�tI>0q*Ӫ��K��k�N<5��L-ԳO�����Ή��K�ѻ2��S:M�l���Ӽ6�&��7L���I�	M�K�`�r!�2�s[P4����*�z�.�5thو�';Q'v]����Kt#��M����P�0��[������|��Ä(A޹z�qS�h�ZM�ʕ���N�s����et�(�\�ˢ�9�q�tJ%B�������M�*�`,
����n�J8�S�e|����L6�L^���mk�i��Q_6�Ȕ"ݪJ:H4RT��?��a�B�E�\�>���̡a���%�i����g3�5����n�ݴ/�6h�Q3��k�B�eX��r�Ud"ɥN��v���[!(%2��!@��T����1�9��)�2��wS�e��H!�KD�l�$[�r��Y@��E0�*�
�e�E���e ә �-un^o, %!-)2�:y\䑂HlQ������m�D@i�����eCQSb[�avBRˬ�wwmݔ&�5�]��}���K�M�w[e�l��cs���W��	E��|�nz��
*/���{PTO����������
*��_����o���_�_��u��p�7W�o�����Q��so{��[�\�c��`RZ~��)9 3뒻���PNe�Fs[v�Vw�s8^}tL{��۬�����Y��Ef�i�G��v��;�V�TV�<Y.����+N��gyR\���`ut8��&[�*��&ޕ�r]���bbjU���@�Zpl��&V�W:,6��ԣX����󮵜X��Ik
�����m���,G$�A=̚���ǋ f]d�)9�%��U�L��X�9�R1�ΌO�.$WrՏ���}H�T+-�Щ9��c��f�E��L���jّQ�]f���}�Wv];�9�Z�	b$��!�z�WN�� �i����npϏ��\C��Zŭ��,��� #=�xC̛L �O�R�lP#;n��msqk��؃�{"�\^Wݰ�wi�,	��=7{.�zt�}�+�^P��6Pv�q\f�j��(^��9�O���^ŉ�]�чV��.a�/F<����PZ��#2��f�)�USy�l�El�#̠"�ʹ� �r_�LR�]/��>�t��~�?]u��:뮺κ���^:���]u�]u��]u׷]u�_u�]{u�]u��]x뮺뮿u�xκ�뮺�뮺�ۮ�믎��N�뮺㮺�Ӯ�뮸�뮺뮺�ǎ���n�뮾��뮺뮿]g]u�]|u�]{u�^:����������뮺��G]u�]u�_��>>>=�:=w��;�Ӧ��Zf���u�8hdE�w�O¯#|k:ب�v��2%>h�P2q�����H��lz+�i� G�Y��m*F��_�K��Ȱ	j�el��/�(D�\9s	)3Ž������U3W�c����4x$�t�l�����ƹ�u���Q��;��o��Υ3�dN����E���d�����os�]ս E��X#����ea�f�Y��[;ϳ��m�aq�2�thK_��R�Dl���*�4\%�h�3;���tfP���	x8u}Y��,B�.*ᷴqûwr���&�ɀ��Z��yȄ�Ux0b�=1>j9b���Son�=��N�,�\�U��©�V;�)�s�!�[���v��������Q�/[�7{*������]�<h�GOU�ѓ�m�>�t����V���+�Ҵ~�Q��{n��}�UM����6@@Y���UH%P��JȦ+�֖C�1g���:8�v�vS4i"���d@�gS�F�M���5���'�!d�ln�ֲS9�S��
I�{��t�Q�;��Ju_ɋe^۷L_Y���o�t��2�EZ[I�n��{�·���� ��.��Gk�G-�l� ��u��+����� LL8��������뮺뮿]g]u�]u�㮿^�x뮺뎺�Ӯ�뮾:뮽�뮺�뮺�㮺���]u�㮼u�]u�\u�^�u�]u��]u��]u׷]u�_u׎�뮺����]u�_u�^�]�]u�]u�Y�]u�]q�]zu�]zu������~�_�O�]u�\u�^:뮺뮿_��������Ub�S�Z��	����D�"V\a\�z�w�|	���F �"�M֬�#:fO!UON�+4�ɞV���4qҔ�;Q���8G���Ԁ�U�u	2"��� L�2�v)ś ��Pu.f��c.��A" q�Oe������iF��:uc�*k�A�w�D4�(��z��8�<Gi<K���T�&)�b 
���YDi�,�1ӍS�98�u���ʤ���������'PQCe�"
�}�u!��v�P��r4���DQ�R�hڜ���9�!;T� `[��muS��q�e<�u��͹z�rP�#�!I����ȩP$nb�.�Q����h��_-�;7ޫ��8��M��`�zd���"���U�3 ݙY���Ʌ�V_N�c���@��=:��$ʂb	��ߛ�:�f���pr+�6x���"6&�fJ�d���4��ɢ`9ӵfn	%��:*���z�;,��j5�g��bu(�!�{A]����y�d&5�V�r��xv4ͮ��IwSD ��V܉��u����u( 1�-����k��Hru��������q����K)1�stN�_V9F��Gz�fG�GC}�W>_W3��k^��W��ْ���gf�k�,{ª^V�Mbd}ɵK5ʣ]vw�D=ش�![b������g�[��
{���W+������h�8�}����P��+�ɧ ��9p��UH��VN]�O"���?|q��:�:뮺뮿]u�]u�]u��]u�]u��u�]u�]u��]u�_u�^�u׏:뮺�u�u�]u�_����]u�]q�]zu�]u��]u׷]uק]u�]q��]u�]q�]zu�^�u�]u�G]u�_u�믏u�]{u��~��_������]u׷]uק]u�]q�������^�9��Ϲټ��GK������M�Qv)�v�t���_a����M�n�!q}K7t�u4�û;{*ɮ|*v��� �9e�7��Sxn��Sﾮ������Zln;�9u�Kբs�{6��$��\�H�FC�7�k�Q�-GF�3��%��2��xt��^���ޫ ��m��	�Q��Kif=��"�u!�k��H����9�w�7��{w9	$Z����}�ձq�YQ�/N������Xy3*�{��l��̺�g��M�b�
�5��	���޽5OY���!sְ�J�mْ�J�M����_3`�0j�_f��޾ɇz�e�\��eF����CI�8yr��z�:nG&֬��+j���S�-�k��mQQʂ���ŕŌ��n�;�7�#���z��P*��u�h&G�&'z������X<��e>��T҃�xbuV�r�v��㼐�L��R�ٌE\5�z�O	bձ;7]�Ps]�&iĮ�<���d��L�����̈P�������y�e�kw����Y΁ъM�|�֙:�s�T�:����=���k#p�N�\hg�3��Lhڨ�渲mH$eNi�K�5�8�QQ��.?��_u׎�뮺���Y�]u�]u��뮺뮺뮎�뮺뮿]g]u�]u�㮏u��]u�]tu�]u�]u�G]u�]u�_����뮺㮺�뮺믎��n�κ뮺뮺î��n�뮾:�:뮺뮺�:뮺����?^�������:�N�뮽�����Q1�QQQQ"'1��22�5e!=4�=M
�n�ܫ�E+�xt�'N�%ѽ��Z��+�F�rn�-�l�.&��Z���|���+���w*���$ϔ��(�}�OV��\M9�8����`�� �@����%Y���5���u�r�:��k�6��"�u���1S�։����n��5�D��{]Ig�ึN@'Q)w�be���>ʹ� �&���[���2f��i&��9�5��7v�'�Z'E��m���I�ӭ�yu��V�֥���,�K�7�>]�֪�Ǐ:`}r��V�٬�3W�f��"(�i���U%[��y��rVΕ;�%�Mn#ON�t:�0�ؠ��	mHk�L��4i�i�
Z:�Z8+�,R�3!����R�1ud<oA�0�a��pb����s��J�Y�s%��Iz�|��zH�s�����	���F�ǜ��W9��n� `��o`�]]<[�q�o!�>}g=����yލ�Z4�����\���aސ�1L��ǔOa�/_�c3�:�G�$)#ȍ^S���M�u�g�.qٓM%'& ������F�_l2�܀X�sT�ך�js�w8���������뮺�ۮ�믎��N�뮺㮳��뮺����]u�]u�]u�]u�]~�κ�Ou�]u��뮺룮�]u�]u�]u��]u�]u��뮺뮸뮽:�u�]u��k��믎��n���]u�]u��뮺�����������u�]~�κ�뮺�㮺�������؉��;���޾�}]}�lڝ.�����[ޛ�S��� �6(*ͩ�y�a�Ǝ����H{H���.Z��wi��:��1&W>=R�r�[=Iq�b��1�;{"��iΛ�<Ix��&�;Ñ�p:����)��4��1�Jċk������]��$��7R�f�'ј��!��n�\j�4�Y�6{+�e��{�{�e5;t�6r}���+b�!YBD�7,�
���8ᷡXy3^(�S+Mp}qgR6��;��Ԡ�eݜL�=ݽB1!�}q�����n�z�S塛�ל�f-���lU}
VrT`���*�B�8r�jm�/I/����u��;���#w}���ۤ�zw������ٽ�:�kG}� y5�W[��w"J;��e��w��LF�SsP��;4�d4+{�'���}K��6� �2��	�+����4�`�'tOH���S���6��`��vb�e]���r�:Cc⻄	�T�Ԯ�h)|�,�g�S�U�z�5�-	|x�z!� ��.�ҫWw�t�&�ˡ�7�s8k7|�U��ࢰcAj�\��(��X�}�У�(��ں�.62:226:ttttk����n�뮽�뮺�뮺�뮺�:�u�]u�㮳��뮺����Y�{u�]u��]u��]u�\u�^:뮺��]g]u��]u��뮺뮺�u׎��N�뮺�k��뮺�u׎�뮽�뮺��뮺����~������u�]u��]u�]u�믏��on�����GD���Z缑�#���)-&@z�ڜ��ۙƮ�����c=�<CM�&KB��J�[.�lfJ|zN[8 ����Щ��� A�Y�'r錶�j��}Z���'GjP�sV�7�8�8�+�^��]%]O�0[p�3��R�VA���NY��R�M��1��ŷU��C���Juuzf07�Z��X�P�f���%�����������d�5�����Ʒ>�굮>:��ݥ�b�Y'����ϫMA�%h���{]��y��q u��;����3X���rT��e�sI��ӓ:�T�����fe:�Y��e�w%�5K���9N�[e]�ٮ!�u��0��C����Wd��wV8���Z�;��:�̘�;�"�*�u>����������V���{8��2��@�ƕ�Lד�=24�%1yۻ�+)l�6��
Y��VoN�P�j�+h��q8w�S'��a��Ĩ��o1�)��q��nT���#��Rq.��;{ǎ�W)>�L�n̍mt���6^;�Z}* #� �Ɂs�]p2ĺ���]Ξ�^h�rNL(��;�t�4���븱�P�x���L�����1��Ls�D�P%s-8Œ��Vj�"���<݈���*Х�<F��@��wƬ��s(�ߒu�i��U+��h ��x[y��Wi]�4�r�P�f��	�$9�H�O,�g]�;{1�mle�-%�>���dAn�jз*�oY9q��y';�յy"E�=�Ы��ua�*sd��H��f��8E�c������z^ʀj�'tU�����̵��؛�����/�.���v���婼rm�u���T�Ut��^U�ND�������NT2�̸�X�u
`��ZHM���%�N#�r�t:�6�ѩ���_EY9��*X��|.2:�PNY�n��C'.���f�s��)ћ��ͮ�3W)ҁv����컓t�T�HN� u�͗�I p�ܲe��m۰�e0�j�1J[�����残�q0��ʸ!�Dz��Yк��ҮC$�\���a'*�)VV�+C�\���*d�nr��2��*��R�V����s����=��1��afꇺJf�ɟ%�Bl՗��4,�-FkiU�F�F�v��uk��7��|�-��Gf�7H
eM:��N'�:�u��6�jN�w�7U<y�	j�\��y��X�T���z���G܈�����}[wB�*n��HpC��u��${Y��ܮR[����r7IXt0��(,��űX(t�K�k.Pв�1�T#̌�T���Bbaʴ�Q\ڴ�ڬM�jh�ڣD�ʪ�}}2�j'���0wu.�N��B~/��<;6�[��糍������֝�]#����,�&�Y��G�����Д�"t��U��X��9c��":���ug�j�<�W��lu��[��/ST ��|��UQ�d]�ȘـN{�HҤ��/^�������"-:�.�þ���Օa�%>��u�}�{
������ֺ���x"�D-���Raov�Ȃr��A6�g_ a5�W��/��jݘ��U�Fz�)��s;6�97+R�T�}T��%�g�G!+&S�%��lL�N��� +�ժ�c���Պ#���F{
S��:W��Bkx�33�x�k��5c6��*�8���8s�Jsݐ��(N�8o.*�E���Sp<2�n���mmb��|���|�%��SCM1{��ː�J��[`��֪ӊ����>��+@�NT�#x<�����.�7�C+���yfho;V�x��vˎj�Q��gQɆ�WMcgN��V����r���˷��D�7�}�9���k#-l��D�Fr{���|���0ݺs�3��2+��ǯ����S�+~0���Qy�1�a5��g��9K�(J���I��f
���խ(^ec��!�bΡ���E�e�3�z.�N� Ij�ӵf��YSA�r�e���A9�6^��G�/����GG}����fI1���b���� f6��6K"�TfjK�t���u���蓲
*��N�ѶiS��_>���D��[�\�8�^��ʦ0�-�r�n���w��`Z�젢E�YR�����bVh�{j�����K*�EM�V���W|��Pս�P ����m��:�v���c�5�4�E[�,iՖmw3u$�lջ�K��6�X����+�G��Yp�='	���kt��˭����7O�>�����7���_�S�����������s?Y?s�ߙ��l�/�0l�Y���jM�]��ݮ�ZM�sG@�޻�C��tf��y�� �ܴ�Kf�l�]n��q��]ڠm����a��8�Z�-�ޚ]a� ����@�H�_�����W^s�[9���d����0�i�]�6�SR6�EnME�T�umw	�9|e93Ό�m�-E9e����(�݆o^he��9�b�b��6a�������= �3/���̥*居�G�S/Μ`2܆;4D:wM� ۮFͦ�c (�έ����Tjk�ԑ���.�_<�p�k,vZ.�����Tm^��;g:;N��w��cҾ�R��*=/*k�]�3�E�J��IV{�]��.fT�m.�n����[�M[���p]�����b�U�v�:Q�݆.�Z�9�]8N����g%3�F��1!Su�7i� �ݛf�IWv�.�����a,��U=F[�˦��<ֶ��L<;)p�����#��o_-l(Z�]*p�C1П �
i���R�H^�)�\v��C4�Q�-+5�r�eou��Q9'�m�I�����6�5����̾U�Fk��;3�b�N"+b�5�Jgvj�[�k��/���uHƹ�#}�q��uy�k������*�BAn���rS�Y�	z��!�^F�w]�$���ݔb���uv�+��,�8]强2�44.�*�ewnlX�)�'/.<��i���ťe��	�G�ٶ�K�4��4��.��E�v�)���h�7Pޘ��QU�eފnlm�s���uP4�P���!�U��"�Q�4�JT�M/-ҷ[��f�D�L��&�l&�����6�q�[p2�Q$'�$��<md���XE�����p˛��������gy�{��^���Ґ	�ܬ��YT(!�M��,�5噤��s)$������&��HdW2D2&L��@&LL����o���������~>��<}6P�</a_Iy����� �w �;��T��9�:�h�\^��� �"��!\�T+HSGr%�:���bP��ur���S��B�IL��EfES2$U3$~�&il�RIJL���M�����^������|{{{{}���a�y���'�?nF�u�,2�Ĺ���醰2&��6VET��\�񦣲�lHe� ��6���͗�vtia�!���^s��������������~:��������1�zt0�e��*���v�r�VP �a��.�B��
R=��XU��u�r㛝g���.***4Fǣ�`��>J�#Ș@���e�!�����
�ȑ�����
F/�B�.�===�|q�����������<|}�!���?4����r0Í���ª����J��"tI`A5�2�EXC!B�2��l%S � E��T0A@�&0�B
�\�nj�$�ό�"d6���4Ά��8�B&F�\�6�v�5!�CH���2�g
M0�W�\�2�c�d@#�Q*%�YK�)K|fTJ���6�}�X����3���2^��1��:����}$vt�I;�۫�|n�f������R涠9�w`��nU�m�l�'��NDa��D@F@�eYh��*��H�jh��x�:V�+Z�Q���D)�Eb��SN�S�����^+0|�+��O���]��x*���bsgٵ�❫:�Q�x�+���[��>�	l�����츭����}�C,^T~~i�@�5^�(o���5z��מ������]�<-I�4���Y���；�Z���+dӸk��5y����&�9h5l��A�-��S�w�f���м��iF�
W�<�9��kgNO�	%!d{I�<%>�)-5�^�L��+��ʥ$��6J���_��~�5 ��c�b�ɦ�z3���b]JU{�מ�$JRx��dH����ד��SbVi�گ*1���y���oƇ��_m[�Il�Z�z1���5�o��������\a��W�Z}X^y�PF��:���3GV���n�� z�ܜqd��8ڮy�\[��/Ԇ,��6o��mh�[�%�E��f(�!W�z��J�-�WwT��g2���3%f�x,� *սP����})0 ��.�����fnT>7�^�6��J����y�F�
M]6��V���8)s
����x�y��^�x�f<b}'b�>�|�x���d3��l�Kl LG��"��s��T��7�yx���ڥ�XܪS�`��}�������73��Y[���,�V�;�W�x
c��K�s��&��`"M��r��!i�z6�+���*+ތ���p��~�(c>�:g/��*q���Eg����6Lr|'ԓ��S���!T���:��}�~s�ϺU�9q���A�vի�Mϧ1n���]D��`e+x-�f��9F���X�U�4�V=T
��5�����5.T6M��Ţ_"g*p�� �ǹ��iS��F���2F#m� g�;R�����	οڃ
j�Nm��g���Bp}ҥw;��d7�P��
Cp�3H5��!�<�^�>w�ҙ�.��rBh�L�Ƹ>!;�c�̒�dA��Put�	�cd]ς�v�ް��;m򘎸!�!*}����kw�=.��'�潰-�'#&VeHυ��N�����ޢ��3g�n�����2�Ҡ	�j�=�Y�ᨩ��M�oKL��Y�^��)�ϕ^D)�K�D���k�k7ٟkS7<>��:��a�S�=�����ޭr2�
�5�����(7YҭN���:�!./�=�n� ��E�����Oj߷:a�h��{I��|�)o@lE��OB������,�u�����S&�붻��P�N
��;Vv�D�.|�\�-�ܸ�a���iaB1tvV}�V��jm?Q��*4���oޘcu����&:�����WZ�A�t����{磐z���}���L�< �ӈ��W��45��Pt���c7�iX�*�.��w�u#����B�3�K'�����q<�DX#{��a���Хˌ��f�w�w�5�2��Uv�E�6%��2=ji��5
��n%w���-7��O���oW�(�Z�̷��^b��$��wp��Ճ(�Ψ͞�`�ќfv{�@�)w}{�ۙ&����{hgi4}�K�U��wǨِ���I�!kY���oea�.I����Gln��FvL�Y]4��q�5�c�z�ò\ 
�CT��� ��D�`��ڜ����ICH�F���e
@��u�LҼ)e%����
���.v��btwbbn氲N����11����3�	w]{@��V��+ɱL9��ܪEgG˰Z>o>@j���u�!8��{���]a��ӆ��$5�Z��4����\~϶���4����y�G����Ok*v|;5z�p6�J���n�H�Z푔��� B�p�jg�h���Dݑd�ݥ)\�K�ϔfnf�������+
�@#X�'M"ƶ&�X�qi����9�+s��k����QL����7O��2U��;�o�ֽ�Z#��������C��yB�)��o^aq�Wv��͎ĵ���V��Q�>2�hqa��C�Po&uk��]m�`1w��-=�3�A:��.�v��TY�Φv���dq JO��Z�߅��F�a3�gT��|�/�3��,-�R]3Qњ}}�G�:��H��y	v�D�M�e��k�-���
�Ժ���*B�d����4� �h孾���oI)4	)��e�?u�wŝ�C+i��`6��x����b)b-:�]4]�/M����)��5mOB}m�!nV�_�'�b{�)�'#s]տ��!�>�h8ˏLA�`Fb}*L����2oe:���l��k!�=D�q�����y�zu�,#e�Ow� �m[�[�{�*��=�ek���5�n�/v©zj�fAG���x�7�����.0(A5M���R��Y���b�|�wBߐ�o��vG����v>���e��U�Rr���q���s���-lDS�|cxs0��_��Q��%]QR+=Uz���^�J��s��5ʽ@	�D2�����\�
�C=^�2�O���gP-վ��[>�`�S�E�A��0�u��m�j� ��[0�J���M�ɩf����=��h�D��'w�:Ƞ�yp��u;��ޤ	�oqQ�<wk��_��oP�Y��D7��H���?f�C�Ck�w�[�lu�Tu�8M|���:�Rv.��W|k�U%�}:f�y[4���~����@]'|[R��MeZEm|Ex�������Qhtp��`��@9&VRN5�%��0����g+nZ���7�E"u���Y�3o��Q��>�o��޲�W����"A�{��r�vN�j��)Й�o�@�>KT9�1s6�����]�&0�|���{�OF���ӂ#Sף-�f�
�¯V+�˹wQ�N�q����f�?�� 
�M{�l��a�E�$�,	J�m��(H��RT��>�́��{e�Sbv�3;Y�W���J�J�����z� �)7垿s���b�05�R�r�1��`6��o�?!�O�,}U�sʷ�]�b��`� أ�v@�o'�K�6_�P���W��>����l՜���и�@s���Q�0{r��tN���o�9�Z��߱�qH	�&����ka�)]�+��ew{��b�k���G<����j��ɤ��e�+={�����uc�V��09�3Ef�T�*)Xk5X�4�f�[/���p��o�y��p�X��stԥu�K�fP�f����;��wF�s��5����Zd�a A���������~<^ml7!��Xtew��������K��u�3m��j�#0 ��ۗ�yW�Y2���h[TSlL�����զb`̍PM�w�X��x�l�����O�zM~W�9�f���s.��҃�j��yir��7|�r1#���3dN�e�WXLӓ�����k��J1j�{3��焪%�D�A�=cz<�y�j|p�f�&Ve%��b2�a�8�O'y{!��'��>?<�=��V̪pd�����5�}Ig�����
g�u��P$b��Vi�ٳ�\*���݄^������Y�&w��oZ"�کX�����OH��f-�OLҋ˯v��'�w{�����1��'����H��ڍ�T@w��F'c\�>@Ҁ.6�)ͺ�Æ[� �>���"�Ė�����>�i�s��Z��ߧu[=e��ۧե���MGu)락K	�
����r�>j��>5�h
���>��S흳'�	�g�[,��tX�8mj�M,�/���OMSo>�15�iJ׫��D���J��B$�m�xw7�;�շ��#�d�oS��[����P�5���;�����P��Fx)u��(Vү]z��m59>"vB!3j5,��fs�fWn���T2��]�7��k9��*��^AQTP�ۋ˹�q2�7��5cJ�P࠼D{2`��F�,�"�"�	g�!�M(�eY�������KL��e��jڴY�M�fC�x��J���]BSd_z�'���s�:�	��wK�m��2�'5N�;U��S;�~�cf�qb�7<D���dQ��N3/<�k ^ݢ��&�����h.������G���ϊ�^��ߕz{���m��͡3yM���F1���� �50ݑ��cW�+D�u��#�}q��V 2v��t�E��4��W[5k!#��6g!՝`g�q�3�s�X������4:���Z��Lk]ϖ�
�׎�w<��3�,3iFQ�q���2�&�!xTÈ5V"�2�9j�D�f��K���4�q����΢N��~���6�lpT��l�;��Y�j�`�n�3Ow���w��6D�XM���2�����A��R�&f��,7���spr��A���ћ�f����$ᒎ����r� |�2Ck��9��!�����l�9^u��)L��l����޻�k�I���*%�P^���~ly�Z���ĭ)����1�����<W�ZG۞��cR�Q!Fg����y}�]x4*�H�ö�K�����{�2�v��`P%��͉�:���P�W�����J9��P�n�Yd�u��1��x.s
PR�&Pɽ��A��e1�h}̘
�Vٶ �}���M�p��7����j41�c_�F|ܐ���k���B,�0�b�!����m �=H��W�-`�@ԡe;��q�e��4�	m_���mw���J  i}����z��J��Ҿ��S+d ɣwi���Ӌ�y�����/�{����k>�rS�L0,
�z���U� q!�^o��j�Iɴˆ�q�ɛ��9�����d�]������&]�eڑ�[;�$�a�`��KS�, ܐsR�i��ܥb�!����O.A:J�l����le���s�ES�jf��>я	N�ں�D�,��7:�'zSK¤�T��t=�USw�GS��w����Ƥ����缹-��4�QVeuo�U��E{�C�Rw�����b��3�|��>���[�w�\gS�G�Qx/F���]�GdTS�ݗ'˫��C�*�c������Ys�L�\�Jo�� ����K�:Un�Y��妁��[�^���o�1�bR��g�nVS��F ��gg��Y�-���Č�b{*��Ld{ A�^��/z��5y�.��}\��ݳgF"H(:޴�(5	Ϗc��6�1�(�Ixp�ܔn�ۗ�_.[O�/���;5�\��rb{y�IJ<�}���k�.qB���]X���jp�n�g'��d�Bǘ����3FR�|�Lk~|��;ڼ�ڭ����uNf�͊=e� z��`�؈b @?�]���j�}8��?X[}�&��v�쬮ޜ��u;�8&�2����Z����X�̍�'��T���1Ր��ElKV��FwQ�v@ZP����CMͰ�gwt�_�cT��̋0�� ��Z*؄�#���0�Ŋ-8ޙ�su�V��]u�&�N��w�AC��K6P�������E�Iܫ�}n��,�X|+��R�TE��OvWkb6�Z�={�e����Vt�6@y��[�:��m����.��y�;�dnEЮ7/d̶�)�[�g1��i�A�������o���ϧ]H���� A�rKj��e��ۄ
���ڕ�ˍ�ΐ"��*mp������Ҵ���t{���\�T1���m�zߝ���3( �4N��	O��t;S
Q��\��bKWF��}��ǋ�qֲ����1��\m� ]d���N=��(f�X߻h(���OtP-�JJ���e�v���t�9��W[�7�*9t�m��f���q����s�`wy$���;i�M/�����XZ��nfξ�ˡ-D�,�wN$��jq\�ي�V��ڸU�d�ά�k��r���|�6:[yg!lbEqR��V6r�?D�Zf��.l-E���To�l�� �J�Ef�vib-���"es�6�bX)��3$e����� 2J��;�1Xi�Z|ɯOmq��F���1ZZ���{�5fP��v��*�H�bl�k�P˂�g=�#{9{,�z��CPWd�N�b[�lf��1Sf�7�[X��)b��pqh<Ɉ�$�(��Χ.�tP&m��s�wS=:��z �g�,����w��!s9�9mf�n.J�^������9�r�c@ �t�����Ϡ�#
�R���n����d�586��r�fe�vjH���9qjg1u5�.��������fv^j�m�ua�h���pǳN�,C�.N�]� h9w4�*qf�5ow���t�x"����ZkWH��rs���vcug�"�#�:��as��PR���/i��;�6�+���t
�Iy\�H<4/���-��l>�k�� J)c6���.`s�w>֫9��q�9;j�u�2����9gܦ0������]3�57��dՑ2�R��d���R�Seh�Ԩ3�t�>���祿(�IvМ3b|�Z�t�nG�y�#��=�g`�y㍛ޖ��e���.��.��u�wh�9Y�)+�!_j )|t�L���z>Y�ȣ;Bd�*��9��L�E�����q�w�[��o��}�)���r-rҔ��c��*�+�@��A-A�D\(p�EEGEED���ǃ�����۾{ɋ�9�E�.��eܖ���`���քc+���ٕ��.9��}�>=�����}}fx���xz�s�.GϽ�n��$�� ;r��2�98��
�\\'	�^<zx�~��>=���G_���L����|�+ X1E>���X� d �FR�b�r$EL2�2�Ƿ��������ooo����ק�r��� !��#h�b�1'��Xo}l٫ X!$&@�?�`��*�q�D���C��=����]xϯL���[<'���V�+�H�@�[hz�}$� 4갅�B�+�Fu	�U( �B�*\dTTTLL`�FǡA���� �	>���\�L�͆2�"3�$� `@1�*#>�1B�Va���B)Ԭ88D�0�R�Cc�Z����0!�:m�ц�p[\�+�Ձ�a `rZ@��� ��X�vP$	�n8Dp�IX��	9� 8DL'De�s��a`�$�䑠uƇ ����,$�Y����E �'���G�;-߳c���	ی�s���ǰ��W�_m�cgpMO]�3�)��j�Y���o��\�;��~g~w\���a�f�����d
���� ƀ�_@|}���$j@���S��0}1� q�n�1>�.i�JJ�:c�'�M�EF��~�]�-aą� �w%��.;=�@��� Ǧ���he�8�
�:��� 9�@ek�}�t�54���f��5+ |�56�S Lyq���>��D8�]��P��>C��D3�C[�d�rOW��4xb�T�z�_j ��N�6�I��Ǡ�*�`i�1�f�>�`��1���+�/۪?{~}c0������ ,�s!.��O���>�`O�a3Q*�#~H�f׾��������<����z#A4)EùD���̭�<[���F�q M����+«�q�l)4���UW�����  J^�,+Z,��Z�����������FE�8����6r����,��}[���t�0/��\K�M}�{R���s=��θP���p�3����`2,9	����o����c=c����xkr�>��L�٦A�2_&z_��5�� ^G1�<~�� �s$�C���O�` v\��^��<��@ϵ}����%���>�W}��K�1�}W!$D���_(&��=13D���@Fkޓo~�2�{(F�" y��ߕ�<�j��pT�����V����t8G~���ߡ�Q]�B�ZѺ�,�������n+�=�t����X�osI�	Jd��R���%�&	$��~���-?o��_Tޱ��-�ʞ{��/#�vʕ5`T��F�fls{e�Fn��p>�可���A� �b��P�����x�@EV:~v@���}��IH�i6� 8�ـ���҈w��x���
= m�����R���m���@@��j I����ңN��LEp@3u���2�BD"D�L�����^!���#h�?��{�NrRAL� � O¾ف^���	4Xl=�aI��q*B:1A$�0�`k��)�W���W�.��&���7�� vw���Ԁ1ɐ�a���f���#�Q^��yQ�ăQT�$q����p���@kN�o35( }-�T_�D|����%z��@z�67��fKxVnu�l���uQ�8��p����� ��AM��+b��ҏ� h�>?lfH��ߦ q�vr�'7����_\l��c�מ�A����~D��Kn�8[dgP���0$9`aϖ��s)&(G@aW�'
n<�&�k����z]���Ȧ�oL��KY1�A�4Y�<���T����q�0�P�yt$��P�r�z�h��"����@l
@���� �S�J����n����\{�0�}�J�?nv����q�fHW��	�vb$5q��P+�����@Nk��!�fǧ>!ړC7��_6�l_DF2���]��t�u���r��b7������<^��O�8i�C�����oUL3�K� ��d�a�]p{Ŝ�)-�Y"���]�O��0&��l��X�-�`壨�����$d��9��;��;ţ��m��V�Օ�f��D4����y�Y�l��I���L3�,�	���VHug�<���;��*V��(�OG�����b+&�����P��X����I��`���{5�;���sW}���jzt��\���v+�n{=�[W������'�> |M�u�i5��>�M��og3���T݂`�L�k�q��,;��/���P(/z�� M��]���?2��@� ���b�7�E����]��ֻUH��ziFH�>�����uhTَj�@�D�{
���Z`� 0mn`5����K��c��WA��٫��}@&�0n5����uq���� �c6@�z-��BJ`u�?�O�Cp��t���������+������P:~z`h�~�G���vt�\��(��WתKF��"h��p��!�!� Z�w"4Ç��O�\�d{�����E�0u��.���6U�η���K�0 � D>�v�s�dV *����~�Q�&��񸕑H�>0 ��}�����[ߘ
R��M*�jw�gL���ͯt_H&�a���!�@�}.ψ���r���z@
N�>"C7�r��
���#�:[�v�|K�{}Θ<�G�4&�y�$�DƗ�%�����0Ԣc�X Y�^�[W*���hT��m�n��_N9�5:s��)|a�#Ӓ�ϔ]K�������f�(*e%��|l$��'fi����j�Τ�F�*P���խ�7�:��u�f�[�����vwt7a���S˭����=��EA`�1�B� �Bu�cݝ��`�L O���8�7���d�Q˩3e(��6��^u�^�gey������Y0�p�[�p1�;��$G�jG��f�ӁFa��fv����O9�`ۻ�LH��ޅ� �Y��&��V1@���D��n`�u����zX>$�^����G�|��|����3�� ��(�5�y
���"� .�pc�TK��gaC��8g�0��ɀ=8��J5G��}�6���m�>�^P�p��m��z��^�W�q���� 1��O����o%Os���ʹ�v�դG�캁U�e ��H�Ƭř* Y�׹u�p@��x��'���I�BO+�̂r�5۳y�������<(��Е��Q��&��/�l��6>�6X��Q���o��a�j�8T��z�0e�\r��¸	ݑ����ֆ�o���5���g�7�E���7���90��E�&�t>�J�����Y�~�u�vF5xM���������8X( ��pv�k/��n���;gdst�7��ǻ5����z�b�l3������z�{����3�b�p(c� ��O���RX�[�\s��ݐƭ��lP�d����q��Ě��|/���^ۂhP��ﱋ�ڰ!w���B�& dY�A�4��w<;o*���nL� ��%Y\��y�K���SgU��u�VsekƔ��ͳG���T�A� �!
��ζ�}��D?bRo����:G�Å��u2v�sZ��-V���i�0z�!-��dj~?�`v��5�u�f�k�)��ߡ�gߍ�9U1�{��P��s��O^�s��Þ9�\y4�Jq��ħ ���r4�qsPz����`O�q5a�˼������V���ǟ�tf��U��&���RO��"m���]��EٴZcn���<�XO�o�nd&���D�{��S�����kj-R]�ȫLzzz�G\;/)��5�h6��,ٛ���u���Ihh�|���;'л賙B�F[�2P��N�0xoϋ��;�!j�2��ݶ��k��?ywFBL�hY�g"i��M\V�Fj\B�W0ӊ2K[vE��&�'��ײ�9�<g�W,����eI�"�v����2��9G��c)�����2ݙ�Afh������XG�Q��n4|�Y���-|f<�[��3�������@�$�'��̷\&\o<�f�����3s-Y��󻲵�B��q�}�O�f��&��bWo��^�[,^[3^'P�L�Ẋr%iV���H����J�I�
4�?e��rl�P�C�o+70��9��� �$�$(&9 ��Y,Nx���>��9ʎ��x�趦Yu՟���I��B�'8<���3����h�`�C� �`�1�6w��ऄ�9����zb�\� �D��žS�~�L�Ә�k�Z#�x�Ыs�Z�l����{��Q�㼅��ϤM��d�b�1��ߕ(~d�M���kK<�
�����l�����ޓ��)S�E����G_b��ZqS��=�F"s�!��Ӎl�:�5���>��%��'��[��&�w>�f���P����@��Ey��B�"�^&5MwJ2/v.>�>2.�˶�r���[���{˦���7|v�p0u$YM!��a�>�z�Q�T�-�W/4б�6�qWn)����&K��>���>���u��
A�kă��(�E{ύ)��OZ�g���~���x|u���/���n��6����d�X���֘J�^Q+��'�&r���|g9�4�y�y;�%�����{Ί�R'v{�e��-��Y �3��(�W�v����(�m��.چtf�����YY�FW�D�H/�^�.	1�Ϥn��^4[�y׶	p�������ݛ~����WC�v&�w���S�Ym�d<`^���?8�rM���dz.(sxvsa] ���jK;e���J�Q�O� �WG_���>9�u	�wm��VՅo���2$W-F��`R�
�!!�m�� �O�w)S������D的w����gv=O:��{��<}���ө)�oS���'k�w�b���-��y��JmJ,�i��\���l�b�9�u�F���/.�9�?#�8u'C1�82��@0 �,������JKp��/�h`;���:?�I�(i��!��z��
Sly�C�y���l�ʻƽ��㚇ܾ$��Ic~��t��4y� j"�@@���'ѐ��9�E�X�yn|0��RX�'���R4��R��(�a,P��=����{���}h��J�H$�c:��P8�
��Uj�q�Ύa���=�܆X���5�ջ/�)3�P�:q�⻐ۻ���T��p��z������)�9�bZ}N�}�r��ֲ���c�+M�g^A���ja�1����7n˰��v$�0��D�+>B�!x��4��b�j�l�<5Q�b�v�c�m���8oX�.˹;�9*�ь*��W�Hȭ�S�L��pd)�lvfAbh1	���;�f�M����^��v��Iz�|�2�����K�(9I�!��|~�y��<v�f�5���t��g��U瓹<x&�M�L;K��`�֦��0�l�m/f���8�c]���\H}���_��4:����3�����ɥ?���|��pg�$f��D�q�?d'�?c����I]*����"�L�q~�EgFxmM�/�J#�!�n�w����:J�\��97Z�����0vK�|@��� �����;O�-��S�x�,&��QsFҡWjr�W�\M�����7#2�U޼�zC)���D0$2�2$0�2(rP>�{G=��f~���݄��~�P/Ͳ/��o�G5N&�=�u��Ҙ]�>5-�#&;�-,�=m��e)0o_�L�os�=s�侉yn����X��2�n�?�����(Єֱf��a����i�v~5��P�B���g_�L0��Ձ4y��L�6M�V�Qwu�����mi�c�^U	H�l�fM�o�!�j<�)���>�Ŋ@��^�̝J�	��D�g�� �I��v���fY;$Ŋɢ���|2=B�}S0" �joD�>2��y�CQ��Fbց� j��C�>R	�gO^aɎ���o���+�����l"��E ��z����P�T�Ϙr��Գ-�� ���Ṵ5�a�X�>@��k�V��][�oۄ��G�[R���Ē�g"h��&G΃dU������=������w6�GO��|�7Ϝ�خ@�y��̥f�T.�p�ث�#}1�_/�ѱ�l�ӕ�wK���vnN;�B)�5�>�>��c��MM�~�)]���6\O|���3�#�N�P�z˸�q�L3��z�.��C.�=C�譻9&ǋ��sk��tEƹ��E�;��c�K����Ӻ��������o{�����^�@E<P��+����f�r��on�bgk���)�W��9@-��޷�?�'�dde�T80�� @@� @^�w�/������ъvXR���B�;�M�:��Y�E�5�����=��nC��W�5���?����Z��\�F�>��WE߽Yk�0Y^�vG�n����+T���ޓ�����֚�}����&���ץȁsP9�VEy��u8����^/���\wOc�w�z3�Εgz�+<\_����9�bd���x�`S%�q�b�<I�5yQ�M���L}O���{j���f|m3�b������%� ��7��	���X���	yj�ΠU���p���Eè�s$KMv�g9<��..gK�-��������>�o��d,52qDF���Ȗ42�KM���^����S���2��rm�h��E��`DD矇D&ʶ���3�ޝ2yt+�n�1���� 2����V4T�T6���΅޶�$��!O/���b^��k�.q�����T�Ƈ@�h���!� 5����͒�6�n�nI7>���z��R:1=�FV},�8Ŝ$�����G�WZǒ�f��F�=��?t�ޕ�\��:ΰQ	�]sƥ{�X��LfTa��h#�m�~63[��q���׊~�t
��7^�\5�ܬ��lXx��X�6;�c6w�i�����b3�0�&�DM)����w��7��k�
sI��g���ȟ<�*d}7�AW�o���˾�H�u�{�
y�" � �" A%C�2��w�~����^��!�:�j����a8d�ߙ@��P��`t���:��Ϭd�^��v�P!��1U1
Y�`��a���D����y�{�R��c�K|Ӂ:��4����&�X3�}R���\qL�����O;��]z�I ��3֛8���d�-�Ic�Ǫ}�R��;m��R���q�:��`Ѻ���Yn��{� $�G�y�u@���qn���L�,�jM����ٝ3��ɗ�ʍz�d�,���+���npX<��d0��{�f�*�e��逶,u�v�W����+����ف�kZ�5��izۺ��tF����{+�<S�y���fCj�j�����,2��O�_�y�2�W�P׍Y\����k��xl�c�����U�����-@���Ț�(>foW8-}l9�Z��,�u�!�r�Q՛��`Cz�����j�YC[ڪ�;n�
��Qh���j��%��]���?)����M-�>@	Y�^n�E��|��Ô<>#�$45t6t�6ѳ�f�/~����=\�9��w	�3-����H�z|L$�z ��}�9�:�#�4eG(^�m�	bظa���"�5��Q�?'Y��?o04N�<J�)��Y+i�6v�{Y�s�-���<cs.���a}a�]Y�5��w�'u�_7y7\��IZ�_8JJ�k��#�u�Ӆt�u6C�6����w)j���Ԟ��:�Ʋl8�C��_V_N5��M���sq�o'�����)�n�>+�W	ΐ4���ʚo{����'�J��YƸ_sTX��P�������V4�m�vM<m��X8�\�q� �:f�K�j\=2�?�bmfT������a]��K�v�,�s�v*��ƚ�U�!���/��q�l��:���
4���� U�����˃�E^f���wx�S������X��MY��N�b���ö�(���4g+��[�V��W�z���E�7r����WF����5���	���B�9���7I�t�+�e�ɋr�n݋|hږn�cl���QXXM��J���N�s����4s��gX̬�^vD�	�7FLUq#*�WTse��5,�kkI��fn��lq����h-l�}����>\��m"�D]�ɱ�l�Mqb����7\�H�R��n�`R�(.y(hn�R������{Lr9���e^U�(�� �D!Hn8�1��
�y{(�N������.[���k0������H
�Q�yНV.�Տ��BRɪ��_� �4#n>"�=&�^�;t���[��	L�Hj��p��4�	b�9[4���� �|>��[�x$ AǢ��	>��A����=h;��E
�Ydۢfu��<�ì��@m�u�������,u﹦��N��K��C��X��g_<}�˔�ctSlNg*|�5wv�i4���d�����Fé�gI�N�������n�X!U6��c_Z�6�˽���kBs���3Vv����� c0�D塺�YF�Ҝ�ʡF�yz�u1u��=��w �"��	;�Y��}��Z��ĺu�X'��˫�R,+8��nv��'��&s*cov���l��9c�#�:��V��7ǯN��G'i��H檷s>8+B�Xh���QRW+��y�(�1Ǵ+��h�r�V_]�{/�+@U�������1+�G%Byݠ����u�P����p`>y�6�SIbx��ڝn���2-Mc��m+1J��E��w�M'�Mo怷E�ZJS\�-�|���ӯ#K:�	���c��Eݲۨ.��Ab��l�����]E
�����c�;��r�)S���p�����]�]6{
��gq�Z�o�+�M�F¦�ݢr��_��΅C&�{�:=�Tnau.]�lu+i��5��1�� d&��e�8V�9���BoM��SP&ސ(�KO���u�ەy�jqd�RNtGA7F�,�Wy���h��QS,�	 $�BI��0��o!�Q����%�m����zͻm�n���WK6��݀͗X�ei���ܤ6�Mb�3W���e�&��)V<����m�%����H4����)���WŨ�@�@$�}m�m���m��4t�hB��H�B�(\u���P��O�VVt��Wן�*��/�R�1;c(�9m�"b�B����K��0 `��R����.nx��}|||{{~����>�����)�,L ��+��k+l�
���,1VA�ā���� ���.�D�Şa�<�γs����u��<}w�x� ۑ@Ec >-`�@�	�m�d2Kcs��*�F�����{~?qǷ����׌���=�"ǵ�@�j�m�@�b���'�p�! `��0@)r>�Ƿ���q�]}x�}��
�d$	>q� ��C�0>6�AN,%�0�(��������~?\q��������x���'��WeO*j9q�A�0�[I;3r�Q�'K5gP���+ `"(��9яOOOn=��\q�G__^<x��>f|��`y]&�( mh� �@�����j����q�4Kդ		G H�@+� �	�;�q@	�"g,�9���!��=�:^)��(E�\l$�,H|& 0 %G �d�xR��]�C�r��2���$	��2�=������ J�BB
�$@2��*��m`J���+��^!80wqL`"�=�/�.6z���C%"�!�N�q���@:��<NWڼR��WZ�xjb2cser]sRuu�z�:u��$C�B].�S�>黶���K,6X�d4���%ۮĆl�6�\�V�i��I��C*0�$0�r@�eBQ:HE�y"��e|���w�N�F� �> '(�W���1��]%�^�������P���6��:\M�ihfm���NĄ���|����#\s>6!�y�*�L=�0f�>�zJ��gʫZ�-ƅ���)������T�2l�FZp��<ϗ��%�0��no#�NuCk ڲEk:����|h�]�0<�z�'&m�}��g�w|qȝ��6B�"C-��r�z��8�4=�ϙ�ʔ'����Ű�S'2�X��eE//�����!s��Q���P(�4��c'|�P��2^���%r�m����=�8p��� km����CH�z}�iz�5 A|���X����7�����MTg�Ŏ:��qmB���oҌ�}V�A�>,�����]��cĖ���C�+���%o�D#W}��|�dF�K�o+�`Е���D��)�E�e6����:�+b������ڭS�o�1��ݛ����,ʲZk�VS�US_��x� q�����d*�gʣq��5uƚ����?k�]�YyW7ݽ�t��	ڏ�n+��ӳy���P.�1����p�݅4���9_F�B5*=~(��?~�zS���)v�d���&(�u�^Q��<��r���^�1:�Y�[����p,��p2�Z)a� q��Wf����^=��6�x7�>Q�K���-o����75p� .��t��˙Q�K�Z����4q}X��.�W�Ԡ~Fa�aQ� �P<���@ �߽��}�y���d8��|�y8�v/��3*���N��ũ\4�7�N�!��,����z�m��Y�TkyJ�8K_�[�<c�q��ߟj>׻�K#����][n0s@ݦ�$�pӭ�r~�>.fX&�yӤ(�y�s�:g�U�H���V�����e���I�<��=��/J�"C=��|��r��%�D�efht�s0��g��fG7x��g��?C�ۙkNS�P5Ӭ(��zܼ�;-{��5�9�][.ۊ���v��u$G܊+�0dTw��w�����5oD���sc�~b^}N����ӻa�Oñk"
���@�l�[�v�����"�G��!���N���'�ϫ���f�Ո�{��v�EL;��q�ba��E�$���<����hÊzW��:|@�)czf������]Cɨ�\��5�6Mca��]���;���#�ϋߛ��=��!<D�G�n��Lk�~�hOޚ�1�F>P~ge{7�q��~��d}�z�
	I\�M�w����!uI �rU�J1��GL�4�ɢ�[�X��=��l�\�� Q|�V3�a��y�1!��%)����/l�*#��sNL�tٸk��ɑ�>����VW$*���Ĝ�aL��E�5�t�&���uʴY�ӜhdA\��e�sz3QQ�]��up���)����߬Vf��-Õ	����5�����muq�P�u���=��g����ə���{Y�e��#�� �!�dVE�a2�A	�{&ޭ��}�)D����p��������c��:�t���èl|� ����PHǻ��K�/&Z^�=Y�z/����t�A��J9�3�W3=K��]ʺ=�� T�����zR�ov�} 2��ǹP�(�7�b�fgD�S�����@3��v"4�|��G���]�r������m���3G�c#�;g�:��̱r"۴��E/�v�T��7�>1���:�;頩V8����L�'M`�@>}��$�J�8/��kU~/.y�\St.����#����ژ�y���� s����??78�8f��18~�Ϋ�<�ˠ��HD�����z�~�V~Hh�����}�g��Ջűi�A�X8�`<k�w��*�"M@~x�NK����q@�)�=s�P�H_	�g�M�a:�9�+i���v���0K
�S'�c-��M�Ĕ9�X�t���{��e�qܛ}�;��:q�=�����B礣K��zL4,d�XX/�'��{�:�	f�8j��n�[�,�����Ad�j�8s�����{l7�Q���$p�_6��yH/ˏ�o�z6eV�k`�+�='��2o:Z[�J���U3R.�\W������&��쌎U�������w�<p0w�2�n��2Kp=����Y�u�07�v(tޙ��׽��#h��wt�SAeM[]5K��S?���=�82 C2��0�(� ��;��{�����_�<� ��n�v�F����Pd�@k�bG�=(��>G��Z�c+���^�T�����/6�]���yǢ�+}�3"?R�,�dRV`w�f+:����$�`n���,�N96�h�����K��&[-�N)X�������=��XTL}��0¶(頱��b�a/8S<j=��1�l����1�j�%.��zy�]C���d�͖P�{"���uc� ��0"�#bB�l`4|dn�+G�=��������IO{F8��v�Ɛ���0^cT��RȔ�z�%P���h��Ly�]�xDC���U�ڎ����k��?f��S$q�?z���쥊�"w����Z� �i���w�uֱVv�n��2̓�tL}��/z��+�����"=�.f_�G���T>�D D�?6*��\����[Ŗ������7�z�\�o��tF�dʼ���7�>k�8η���;��L�OB�qC�7��� 
6s|	ږNT[��	O����U�m�g�RoCח�L\�^�-L5;��0]Y���9�!�^©Ýf�MH��dl����7� ~�W?H�k�rU�I����3���ܾ<-.�Yå�]됾�R��K�Ƨ/��\��N�z�k��*TO��Z�:	F��߮4�@?�\�1�.�eA�*�I��L�q�X�������N^f�5vZ��!�-��o��u�k��u�J���M��o)V�t�:v�>�vL��ˬN�n��J�H�m-J��t�(c������,wwe�K�4e³kw�2~f�2�!�dRL�X$@�H� � �--{�^L���h��i��E�_��8��Wޙx�=��ג�2�H����(-r�YBޒ��ٟ��Z��20"��n�t=�L/r
~����<�5� fuVP�5!��2/H��Ie������p�@�z����y6�W-��N�yK�r����6��/>`�������hkBa����(n����1J��4�A��Dj����"]4&��h��UO���Z{�|$(*/��5X ca���ך����~�G����zd5����V���T7�$tm�鯕^6E_rj����I�#��|ŧ�y�~�>� ��(ۗ�$
�>~6jP�"r>��ϖ岉�2�dQz�nz�ve�K�՛�W$8
��~ǳ����݄��g��H�,����oU��C���m��H��f(������FWz۩��ó*�
k)��x��.��yJ����s�9lH_����������	���"}�ջ���p6��a	ạ>������Td�d�X�p~{���.ύ��o6c����_G��> Nα����k���v��9ܱ��-G��55�2~|e ������lC���$o|���	��g������kP���5W[`�Z^��_g]>,�4�_������-�,3\m�u�t;���ZgН���q���V8.'�a�&�����W��δ��onU�����Mnz�Rk	G���ڛ˷���U��2�DG�D ,��	��(2�����Tx$��C1���/� ���~v�J�lYb�Y�?��"I�ǚ��N�� ������m�(�O,���-��{��)Jߛ���5r���  ��U$>�h�}B��~�����~7����j	=�b�8�-�����fiY\��(���й��>�r�H��K��j�z�zg�V�j!�z���+��%9�L���v/!���o�u+���	�Q�+r\ ����=η�<�٠����I��U����  �`��1��BՋ篳2�w�93�b2)�x�2~ d�=�F���y�[��$_���@͋�lV�.z/0���D5�?	`��Ͷ�q�(�A�@�/Pkݶ$%c�I>���BF��d�[2ʟ�@���k�~=��s�yO0�l�x �K�~n�3~/E�t�qQ��݀��0�Q�xB���;J�����
`�LwCw�/|�~x~�>~n�k7���m���,6Ĥ,�O��4�f���Ϸـ����W$�1jQ+G�ټ�q���t����9O{�I���LT�JO�9�c��C��3߻�{h�L7�< ��|ƈ1�B��lT��BK�������nTL���h���wm8� D��ax��W���Q��o=
�xqe��J1��J��O�}�^�I�Zݜ�_p�a.n��-F�p̊��jU:�k�k����`P������^N˃{�|�O���0�C���ȁ��S� '!Q(���Ϊ���4�H7�L����P����Tx� �8Oy�����-3�������=K!67Ql�a_���ᮌ�=3�v=o!B�P�}b`v O�
CJZ���&���bfk%��^}����w����R:�"p,?H�� 2�+(�V���O(Oy�=,�0RTž�wD�J}3�ܓF�g��}��Љ���8�8����o��k���@/-�&�~ޟ)����1�'�m�xq��}l�%���EQ�L�'L�߄	mG9�����@k���*�o2a��>�p`�f0�f'��k2%"�m�<ϫ��A��8�U$箑��L��	����f���p��*)�ty&k�P�NI��Yy��밾-G1�b�r���9�rbe1�ȶ٘J� XIw�6�fM|�x��j�Y�K��7y��z"Lq�>i�Q��Az���սՍ�ݙ}�́�Ol�����٩��ϛ��	f��k��w�=M��m���X��׏_?2��C��V���s�o\�A銳AvNCv�����~t�U|`_����Jf!��1U���#��Vj���}PSKitfM5qm�Ճl��!�n�뼛s�(�F�˵X/u�(u�M�T�C�г������k6���?w�5��݆���2 �� AT�twY�W
v������T�V�\� �N�<�K���l\T��V�S��׎�Z���~�0 G�<aXHW� 0����� �1 @FDE/r�}��u�ݐ��|h�S�a}���y���>�#�1�E�r��I�[)��e�w��W�qYȯ���30�=l�Y
�\y�miP������OL ��ސ�	_o�`d|�+k���klĭȒ�d�	ZQ!ί�]\|��,]�>�Qӣ�i&5����a�sj�S-��tw2�,�ӱ��w��ߔ�B���&Ӑ�B��p��'rvF�!c{�c<�i��M<2ia�"��������̫=&)|/��WB^�.�Q���G��M�2�\8|�ݼ:�z"������x(J�i�
tQ3�͗���/X��va�ⶱ}v�zt�@�i��k�gj��o�n����I�b9�뚩"C�w�a��ڳg��G�:��iq@�@P>� m@�v����� �Iܴ���^8	�kt}~B�⯵����)����ь�ϯ����s�4�1��%2i��[���~�+�ap����x�YF$�P�-�.�D�%^�f{�$Hr���1<��s/T̺�紌��=��ݦ|$�Ǒ�	�>(oݐ�{����O����-)Xş.��_`����;3��`䦱?ܰ55�+h�zp�8c��Y�_YN�����6�y��:/[�r�>h���cYKS�n�`��$8(-�e�P�Df�V�ټ�.��]�_Wi�^;�躜�.�Z�Q��p)ؘ�v�i�Y!Rh�����-R�۵WMU���Nt�î�*��e8$�pdF���dP�TS�Ԯy�2����������Q$7��K�)�B��j%r�O�\}9�R�B����B�*����Ӛ2k{*�M����<l�"��Lכ����7���9��,�K2��hWn '!����6�����ܑ\=,f���޸������!���gCw� gUG���~_W�Lvq�E�+��CMO�Z�D7`ڨ4xa�Q�/���mYLUâ�(^�+b_�O��tf��{ֳ�m��Fz�¬�Þ���W�l(S�Bs���K��VP���d3u�N'�?}����x�qp���j�瞕t0�j��`0,S��	@Mh5��jg�ο_i;�fo����@�ؑ��0~���_<!��/�n�G�}�(4�	ae(�2���;��{���7���%�Z�Q}/���\��)�t�h9�� �q6�V�����t�x����٣��x�
X	���	�(�1�����W�l�-�R/ޜ��3��*�X^|��qR;�H���ˍW7���0�(�\.�K�r
��g<����:��8��jD�ȟ.��F�{_�<����۾k mS���l���/��ҽ��,��-Z�b��'8��[�"��#%b�rI@˟m�ݐd�0P�d��m=���۷[�38���.�@���F���S[/���9=\�P6�
�t�z�t����& G�a��@���N		��BW��OĂH�?������`�JK}��ik��.6
�$eg��̅����џV�OO�	�+Aɺ��ý�쮩��Ω�_�hN���,™1�_1.�TH^�_;7�/���|>��'�1��{�)��WG�Z��]��.t`ai_d �~��3N]u��yy����%�E���]�h�|������q./Ӑ}��^�ϼ���3SV���<����NCT�Q���^�Yxmil�T�{�:Hq�����Z�P,�ww;N����L�o�gB+���4Cc��YMC��M7]�*'��j��3
��t�t���h���=s�]ۗ�V��|w�[�^�S5.��H����_�\����G$�8yE���W�)���h�3aX��jE��q��9��+�@�oA����VGn���SSq��P3F+'f�S�G�!�����=�̽���	�d��O�O�B��'�Os.������hP]s��[c��f�=6�|�49�y���j����ֆ�q��_�*;�o�c�QK�]��H�񎻧3�9m�H�X"�@� P���@��
���g���]7��4���aڽu�tsi���`���)=��J_Z��>����K��]��o�[z��Gp#9����U����U{\����Lh&�+{��0�尊���T�� �T�a���Z�®��� �:�DyWQ��3;��ƚ�r���]MI���-pp�޻k]�T=.*M[~��\ْ��<��kw�h���>9d�鋔�u����H���*�v������ljyp��i�|8�JrQIӢ�9�r2'�VQ�^R�I�6�[�z��8(�DK��i��uJ��T�g�s�w������k5�b��J=k�T7;6V�
��4r�-@՚fpz*4rƁ3'�CF�q�]�,t�V.ΤOQ���Yb\d�:�NϭA��z180}�j]5CA�2�/o��@˖����,&�S݊�q�4��6��7��{{֢����i��{�m�ZM�=}��t�57��?T9�#��5�C���^m��sQcUk]]t ����	w�{���h��kp����X�Iw95����!�F�WS+L���}m����]u��� 㧃�˪޻�-=6���G%�9Fڬr�T��J#��,-�j��0^�wo��eY�[��	l�J�J��N��fҤ�2�һ�J�)l�5w�i�%:B6�Iedn9N��r�}|N����Ѱ�ݟ�EQ
�QQ����[Yi��*{�>��i
��&��e5AYr+�I��٧D�/5�v�B�Y����6)H���cozݤ�R�'���	���A��c�3� +���r:uYAl=�\z#;tT���Nwv��P�|��i����%�jaӄ������;S��!S(�춅ʽ��c���s�7j|�d]���x��� ��x��w����
���9�����v�J�oo��]�k�A6sx�]��[���MJ�+�=�6��m���pO��
K���T�Fa�N��&�ؘn�O�|mq{�KX�d�\��ļB�=0����u�z�];!��n���tmL4_e�+2jx6.hJV���r�z��e�7t��q*��ܭ����d8�3IMJ}�t���:n���]1�y�^�V�=;u�Vr"�':��ޒK�)�+Z!�uj�Rvy��&�'�"�6Q���i�q���G[�xlX����7r��58sC,G��8���+��vl�I�K\�;4sW�Af۹�u	�o>��xLwE`K7�dR�l��{;��ͺG�����i�˱-Ƿi�N#6�?ުN�t�m.g�mt܅$ Y%-� JZ�bC��Кr�3;;���x���ۏ�q��G__^<x��DQ�W�QA-煚�G�
Ap��J\Li��5��@�D��
\\Ldl\\[�������ǎ�o�/`��Ǯs��T&!��� a���3JMP20� &3�%��JE�:zzqǷ�8㏏����Ǐ}��r	�#�FD�r8B�@�<�g�'=d����D�BC�+���:zx�������q��>���x����H_��ژ@��! Mc�$�(L,H Q  .!� Bj��9�����9�gY�u�Ϧ{�g��y�gެ!�)(��D�����$�a@I0Z�&���L\TdTTlc�8�:��������(��s�	�>901S#��"��z��Rh�cLr+�����"�R!1R/N�l�&8���(��TG  ���"D�kl`'�61�cXHDH �$�e1�+	�05CL�9��0d�@��7�%� `H&�F�1{뗖^�g��a�������̽����:�e�+�v�����[�k&]-�ݙ����γ�3w����U���"�0)/�82��>���m���ya���^;�(���_G�y�������pԯΐ��*2��և�j{z{z��H�G|��0=1�S����	���`p��b����qs�� �¼�R�{ix���l8�;��v�/ʎ��yD4՘3�䁤|I��b��ǳ:W��H��2ե_m����:Ǣ�f�@�}0�����j z�	����!����eM�ڐfe^[8&BLH�Ϸ2�{�avd�D�E�ĕ�wp��ʔ/5�l�p.\*Ĩ\�ya�$�v�$0Z9���L|����Q�݊%G	k=�4���W�b�C�{��[
�\��_zM��U�ޠ���B�6���h���ʱ�B x��7_jd���4sE�8e!F���=?=c�5,�X�f�f����{��P�kg���b70����(/��,h�.����`�wo'�`�;AS�+�g����xH�Q�SОF0>�5�Rg�����k� ���8u���QH�T`s�w��ܨ��I��pt�7{�);%�<�t�,Y�= &�e���O||Y�V իW�N3��0窬0	�;C.#h8�e*��}�������կ�ӄ�N�F������o�r�Xg2����/�
��-*z��w�x%׬`x�v+ɳ7GGO����mz�,F�{�s���/�2/���N(y+��dF^(B�@ ����ǽ=������� <i��Ļg8�(�[0׌�F̈́1I��h�BI���o���}���e�;2�������d��a�i��?7u�/��av�y��r�	.��P��������~IР8�ܬ�ݺ� d?ԁ|r���Yb��� ��j�&$bg�͝��뉳돾��*=��̚��t��xF�>��,���;�*�]ŉ����ap�X��� ~��##�y��P/�lm�J��t��U*db�m��k����J�|>ɳ�W�$7��b��������?��1M�~�P�J@z��ٮ=,��_��H�z��-tٵ��zʄ~�Yж�K�ùW�Q������Wp���[�|���Z��_!:EG�$�������E���`9pY� "�[��9T:�9t�i�2Z�|�rϡLF�N��2fz�L��ey�gqF�6��.FO9y�^��t�F��Κ S�>��X�g��U�l��8dik���l0a���L�S�7��W�l� ���rgM�熾]�0�]��TI�7��j�C��^-OOjj���A`���Orŵ�z����e���Ê�yz�S�]���T�~wV�$������fRM�2�;2��dL+�m$�	���'G[oVN;i�����Ts����/xS�w���f�sx<�"҇Wm+u8��ӝrW>ŕ��wi6x�E͓]w-ͪ!%�$P���ꊤ��(*Hv۩ �>.��e��qr����Q�T�S�C��@'Ta�H`@������ @ťj$=�Y��U3��Ә�)eg����n��%<"B�x~�� (y����yT�9�B�1�����k�x[b����MI��W	���8�3fy���I'^�d�>zY�:���ا�!ݳ0t��0h�`�Z��'f�������E!����H9-r��7��A,��C�B��2�����}������ךG�#���B�'>�Q��X�H�߶�޹T��D�d�L���k�0�O0~�����&��F)�`���Q��$��=��DR��� VL[�zǄ��;ִ"zc0VC���;�T����%��<�����l��B�8�mL���xؽ�k
a���W�Y	�w���? �����������S9�ѻ#L���5�dc��W�����r>�ϳ
<�\��t����x�#u��ꑞ�j�n̼�ˁp%Y���T�4��;$�Z���w�H�	F�iB%���N�ӯc�q8����,�����Ei-��>��%��J�P�6�]}���z��G:W<�q�9)M��p����%#����P�>�.�3]�lkF�4"(�w�e����L��sN&JtUv�YY��4ȇE�ze��@PޫD��hb���m����j�qW����8��MqByߛ�^���l4#��+z��2��Z���p��O�:�s���o��6&��#��S�@= �*	��H`C�A;�� ~=���/|�������`��(�ʊg;�m��!F�h8?|��3��[b�5�!񡳼���ȟN��;��`ҍM�Em�m%^;��&��뮍硵	���.���Z��>tѺ��lv�Z�{8M��84z�1��;�^�>4|g��3�Lk�,ݖ��<���E�����m�l���ۣ����ډ�r��P#�,��ƃ��e�C��C�����d�WPr��<FD^��U�<p3�N0��?���m%2!�h/�P�X1��Ŗ��7A��.��Vs�d��	��]KV���lp�{e�oP�'�9�_<�	z�S��M��܆��}�yn٘wl{�t7]�E���n=�xw�a��?B�y(�א"���:2��pdcӽ�<i��[A!t�5�A@
��3n���%��iU�`�KГ��B]��)��9��oL2t���t��W0��P_9.�o�8;�%���^���[[�].�ɝ�s��1��
�������(�K�)I}�M�$F��K����>b��g��	]^�V��[%p(�;}�����ڍ��'4;�/��֦oV^vP4�|�̐>Y[ �t�CR�4K�&.].Ω�q_:�n��
���2���v��rMs�]w])�=] ^ptf������wWZ�w.�{63�W�������ڰ�A� C
�=���aT��f  �Vta]N��5uЕjT9��[����1��Pu�Q_b�M�\G� g>Ӄ��q9�&M
�G��Q�Y
t�[��ɽ�m�At�?�ߘn�;��n!�C*-�S�|!���z�^�#�C�>xo6���Y����2JW\W�f����̡��Q��	D��_�s��z��]۬\��[;so`kow:��2c=��	鸹�s{��Z*o"6S�Y�$9�ۯ=� �J.ϕj
dǇ4Ol�L/��F~Z\Vl�G}_!Q�b^�j9��Ic2K�FI���Y�hy���+��7��Kc�)��3[0`+y�Ͱ����t�sܛ��dM�ʝ�����)���ŀ׸y*0;^l�!uD��ԅ��~a����B,nR���W�z��A(\���iq���;�.,�D�礆
�[��)��������k�Å^�cS�-�Ĥ^�`p�'��>�4�tB��!M*Բ��}�;y��[�,8C�wWf�;y�7����Fuh� �&�dM��b��Lz{�o��OA���u��o��j�f���l�Yc�eN�#��
bZoF̀lg	Z]��4�I�m>�OM�&0j���|���;��O)f��m�%6��h.��qE"_F[��eC�.����@'v�k�����
�*���2�02�(C "2�Z�k��c��U(�XG�!a^��Ljm��c��ǰvO-
��b�t7F"��54�7yg�U�����f�~�(e���+����Ȑw�,'!��B�}�oŢOշ�{��Z��E]
b�y�ѿ:�OU�Ԁ�%�b��[��������wrt򟇒��Oﳾ�:��?X�wۂ�m�L���c?�}f<S�����f��{ks����^��m���р����I��UDCأ�L��B�����3Ɣv�rR��v~��6�?��i����X��kyX��v\�>{]�y܎���]�GuV���������8C�&�q�������L��>��rR�/���5��t��5ۦfz���;�8������"Ib��phR�j���s��*TE|���;�C�Y�&u)�����c�=6�5G�'�Y�9sI˛a+�Ɏ^] ���8����ͭݎ�h���9����j8餺n*��fR��M�E���:a261����?|Hs�����%ßМvs7���xҶ�盚�k�Ζ��ۂ�%^#�7`A�8mή4�`��hE+D�n���Wɒ�>�e�F�P���A�;1��7P.Z�o�#���{W���f����\��ܿ���1�Z�eJ  ��-�p�,M6���]�����!��̐���C�0<NC��!��!�yM}���{�>o�� ��#6c�1������9��s����ܸ?��^a�l=c��t��E��9��,��U���@���޽�-^����)�;�{2G�- �{L�ts��Ds�r[�	S�.��n�uX�F{A��y�C�X����6[��^oJT#!\5��9�T�4����{Y7����6�z$����xK;ic�-�1�}//��ʟ�n��Z��8c��t�����㢅2K"������� ���!��7�*|���P(�%Űn̵���1 VL���cs>��`z�|:g�|����L�`��h���֖����^nJ95���y+s]��#(������"�������qi,Z�A.%�0�6��ѻ(�ɟ}��=;I|�ڏ��*��fE�H�\�H�/A7�t����М	���\d�Y]��Ŵ�m�3���>_M3�J��7�?��&��uD��<;�Z����� ����FR�^kK>��FUP�!P�;�0���A?S5��T����sOex}��*Z�cu0D�F���Ν��R�!��.�#�Z��M�mU�Z&0��[�ޔ+R̬���z՗��@D*�`���;��}�'׷�+Bca�.�g:��.{��K�ܕ���t�n��N�uL��*�|�.�����eR� !������R��~�4߿���ރ����L�U��;6�%�K�|\Vò�!�FE�9eu��~�������kp�Wq�TyJ.&�=�lD���k����4f�j|C�f-aV,��g��:āP�~A:��_��_7�y���a�dj �"/ա�F�O�ߛ)�5��Sж�̾6%K1q�ه=Z�8�>bR9�Z����4'C�	4BfJy&}%�op�a������A�I�W�zS��6�>�T|��}ܲ�3e���Y�ڭ�v�o�C��!n7�c��(��ϤO�jm�*=u䢇T�p��{!{�LK�*���Mk���?oR�NZ�b��&@`-+�Bw�D�?/�I�շ�z�����L���'*$t��C�b�`��g_I`/Q�8V�'ih!�H^�f���8X����'�雸����~�G�B�E�u���E��ϙ*J����cg��0a-3�wc���H��޶1䰽�=�㛸����)�F[�F�R�dϞ�$���ƛ�4��j��ϸ��f�!���	5��+Q�k��lhwf%Fd}��WZI�ݵNd����5�ദ�Y
˪�i*�-����.I��'ϱ*�w����8l����
�;9�}�v�o�o3�.��^� G�D(^��+���x2p ��j�[gP=R�S�S/���D��ô>D:��!���}ЮtFw�k�(����Cz۵��*�yaP���Cӑ�|A�oyX�JA�@�b>A�� h\K���C��kӬcl9��4�uO���>Ļ��������+���}(Y�=�_J,Z���rL�I�k������1hO�xb���ǫ�Q�kVP�0}�"�%�|� t�2���<�'���q��	�'a��@f��Y�$[��c eO��ήob��s.�f�cO��@"�~"{�wV�w��S=���O��!�a�3n���m��.Ǿ��]�"N�!�c7$������G�ߞ7Vj��y�ٱ/��U,+]ggT�UT��q����vϏUȞy]{B�z�%���������W���W�������=]�YM�C�?jƻ��S�s�(���ꡨ����k>��w���W�[�rJa[&O����N��F�㩓C~��
���|?�|�M�o[�	\�G�B��i��'o�,�3��Q#�S-��q��|����c������������m՛UC_K�R<tﷶ^��G�2�p��&/�[+{.�]�a��)SC_VrEPQ�A���X�o'%�g.�b�,\�м��mĄ��t���T�կ�9J�M͓WW����
�ۜ6�"#��@ az�80 ����&B�x=Z[{����ǹ�.���=6��H���Ћ`�;#͐��D��T]̑�U�{$�_]������.N<�i^�za�i�"�Ӥ�ڨ��J�u�B�E�L}C��y��}��KD�I$�H���T��?O�+kP�onĔ�-x��R��^���zfz6��1j���j��D����m��q���9����wo��k^������O�)O�%Q�`G
���F�޵W?`�������P�~XDڳ�)_�&��YL�<��^�(����ΓJwJ����RL��2U�%�#G ��� �^�n#�@���>6��D�c�i�Y�kU����2LfL8n���Z�G4��Z� Ȋ(��"����ϊ�����&��ۖ��^u�v��d��1�O$�]"'}Q�@����i�T�B�å�Ec�u�u��O(��P�ay��ȑ�
2<\4;�}��Gz�̨�@�l�P[]�9׸�~��߾�[(TºC��d���E�|ͣk��=�� ����.���ݵ��� ���韄�?[�n���&x����22g`�G����w�k]%t��L�WA ��t��Nu�42u2Mo3���z��1�s��oT6^��v&y0�����q�^��J57C�m�c��K{�%l��SYg�ٛ�Qڐ�\��t��m���C�v�I���!ݨ��vS�3NF����v��K��Gl�	�񧋁��Kg�T�Wd�)�
��i�����������!n���]�٩��n#�]]5[R��W�Y�u�e�Rg.�W��l���D�i��*"��ed������X6L�r��Ŭ�$�4��0�8��^�]��g>�E<<�s�bK5oBK��^���s-��!e�|%j�n�^wkZ'a�F��}��s�+]#�*�z�����\���7F��sJ�6C�KY�r�$�utZ7�q�x��Z�A�ˎ,�����u�H��u��^����7�^>�����tUx+�� tֳ�0�ȭ���<���:�)rz]�vwvpcm���sݚ�/y���w��Ai��<���2Iܑ�IL|.vm�&cB���qwo�� \n�
���q7�=����}fX�t�`�c�P|�!��a�jRv���g�$U��D�M>('f`|ңI��қ��V�|��7�H"M���V��kME����e�#-Z���ͻ:B�����E���J5/.� %�qdT�X�Ӣ%B�aK�Wb�	�2��T3I�3y��I�=ul�z�a�tr�P7�D�F� �^M��ԏ�dW��^�>�-t�-0���Y�㼣(GH���5�dAj�ӽN����qg��҇�71��s)�+R�gZS9��B�xuÌ�{u���'u*��Ү���5�R`��o�;�ʄ�vUg7@[�S)L/m8�x�ǡ��حםHW�;���p����VGX��}
צ#�$Ϣ��Ϊ�̓�Y��C�g_D�D�{J�2�T^�ݸ����:�;�Pd霗F_f�� �WVP�;�R���jJ�uk�<�
g��j�����*>�ʡ�+=��5"��?���c���|м-�Ȏ��%[�����A;`��r�uv[��a��%�z���Q�s���h�̫,�Q�e�7N�٧K��n6��KKL� db��V��.�u�#�0��wG/n���Z)
c���rc��sH�0�i�W3���J��l0[�'���Y�Mѫ������]\s�2�OY��ᓫXM���g[��vU����e��y�k߀��8�%�;Dɏ[0�`}��qw*���Ω@�;N��$�\s��qlo(�g)��廕�6�t�h!U1݉h�n�$�Ns����!u+EћH���x.��c��n�ݕSU�����MɱÝ4��f�|e��o�(Æ\��i_��NZ^V��vꎓ[]�f��bG-�;yȚ�[��a5f�]���[<.�Fs�7�BҮ�����E�V�b7]i�GsQҬ�f���Ҏ����}Cw�,7	��t�vq�I/ ζN��2��
3+p!#�^��q#����o���s���9���c�8���>�g���8Kr8��\���HCL�b JJd��b"��Ǘ#�8|x��������q����>�g��E�^܈._9��	 ��R$�Z_� aFA��x��������8㣯�����ߔ��%#ۤ0��	 ,!:
2?3M��yϏ���_�8㏣��������U����C�$�0�$�ۏ��l3�k<���������q�:�ϯ��EG���!"��$>l��E"��}n�#��<�rǏ�}q�����?G��}x����~t��{���7��L0�b���"�@� �Cٙ��Ϋ(�E�H*@�4���IxbA��F��"ǚ��%�P=�j�D��𒫢T՗�ފꐂL�YX�2+&�XD!
ڇ+L� C�|>�1�z�ptv�u�ŗ-#�ݯ;�澊>�yוx;+KG�l����9�4[��P�n�����aG���V�i�۝��E[	��!�M�"����XV�n��m�ś�:mH��6;�e�n�j����0���Ü����.�'F�9���xp Q�ImV��*P�;�j>cƯ2��͝�R}�u�/؟2�*ȍۋ�D���}3r�7�K��,$���2-!�I�v'�^Z5N�j:vy�u�ۜ�y�)���ղ�d�[[�]�j�À�
L�s�Įd�a50��*�=[�ڶ�c��^d���`\z_O�����`�����CG>3�q�̆T�Sd>Z4yi��j��)�6-��υ�ѥ�sw[)1���<"o����$Ж��ϼ���n{�͜����Մ��?�pw��2�"�|%��d�[ϛ��6��ƩSƃ5b���u���:���\2��ގ/B^K�T��Za�jΎm���y,a@S����ҷ3��f��Q��U���wB�dn}�!�kr|���"2=2/F`1�e�2�Ms��;��J��&� �i���(%�oê����;4k�%��	l�:0%��	c�|�Z�~9�Vu�-�]�U�rCk���Γ�܀d̖�n���!��ɷ�,"ǭ�C�.��'����ܩ��1�R����[0[�*܃���x1GLd�70o�,������z|�d� ��F̰��DX�2�yx��wQ����k�vc7�p:cUha�m؟����k;6xL��Z��V���� � ~`B0d���	�Xa@oq��{��,�m߀��	 F��(qy�c�{��+�W�R�H`7�}.�š��މ$�sOSp8'X�ڐ4���1���	�Yw�=�R���خ������j�{Y��� ��o�*N&����L!��#�$I �	 ��v�OЮ��4�N�5>�S��!y͎Txz�xE<�2��L=4;�5���	�w"��7ʥ
��F�/P�˞C�8�G�3xNR���B��g�S�)9����(5ԅ��������	槮xӳ^+�����>ך~��V����v��|�h��v�M�
�f@}������ӓ����)��^u�f��鶕X-��F]�>�>��@�g��|]+ˡ}C���p�g=Sr�Xdzp6�1���l��隮���k������G3G��cI]8��py���ϙd��כ��\��+�m^��z�i�����䎦2"Ú7W�D�V��=@_���_9���.��"�s�s�B��â8�d1��a��� ��
���UƗ����_y�v=�Hy�
�Ӿ���h췇>����A�#��h��fi�n��έ6�)\�5�|iR������iڃ/������Q\��`V��t��1N[c�Y<k�K̾_q�w�5�,�Sfe�@�r����W�O�ʐ����Hdd�()}�>}�??�����������q�XJ�}��[?�r�}h:���ނ¸d��.W\bd��{��{�r��b�w�N��f�i'o^�CX+�|}Ьu��R��3b�ۯ�L�5��:�p��w8�O�-���;�d�|o���+"^CX+�[Rٟ~�|��lq0���f�ʡ�o��=�l6F���/r�Ԏ[p�ޗ��3	Y/��y�qe������fo��u� �^%�Am�l�eت(.�ݝ�t��T30�OyT��˶JH�����9
}x���/�.��l��xE�g����M����pů�a1�N��
��˽�y�|�*��/��7tE^�1NH^^�dJ�Rl�퍘�v��n��N4�iLX��3ߓ/��ே�=>�'ZY�8����3�aFlJ�EȈ��.e�S� Ն�9�W5%gOd�w�42� 1Ɏ�Jސ9��޹��00�b>1v���4?4����"b�6���, y�t�YF߄�؜���vM����Q9@���qo۔��c���2m��S;���Ui���� �b�z��2->�X�B=�V`�.k�%�NaY�7-nڱc��%�[�V����4��oY��夺5�m�>7ֻ*���m�Y;2:St�K����:�k7
>��tK��g}�����������CԧR��y"җ�����nx��ge�>�"b�4�g�&C��	����ly)�V/���r+ǮL�Ć�����)��W���c���;�zm�����]&`?�}�������}��G��vs�r�
�����xU�d]v��݄��6�[��c�#gb��H@�8~ [Nl�`��M��k��]�!�*�O5?S_-�����:`3A�m�C����z*(�kb����w��|n�)�W�|6�/V�*��]<�AN�8��������	�L���B�:\�����Y��d�z�

a���K��ڽ��r��a��Z�^�����3s�)?���܍�ON?	�����F	ږ�c�5�\a�>eW�7bY��C��.��f�F��7U���ސ��#���f����$�:5��^�8��)��`���P2o&���{��w�����3��><�N�b����?�͎u�MAn���/��j�n>�j��~i��c0��G�keb�n1��Ho�A���؎ ��3("w_�r~zZ��Y���b{3I�qL�:���#�^X��]���Y�Τ�"v�Fp�DZ!�{�+r�%�]T��3I�Ӯk���.q��w��9ͫXp��Mp��ۇ6�.��t�efq�|��ZЍ&�����Tӽ�啀-�Ӝ�yBpi��6���$����L'����� ��N��W>����|3I蔌A%'EGӫ�	|l��n'$&c���m��vDÔ�DLQ��4��m�v�TS7{�ܤ#gH�^�� ��⁻�4�ր����ѥ�']�ߥFݧ<�s�+���o��ʼ��3����I���5d��W1�oR{wƌ����\-�nm!�Å�G�іk�=���K��T�o*��)��b��l�3/�g!���<p�R��(������P�18y��2J�������>'�۩�Q���,VW���b�����(;��u���B"b��T�1}=��3:6r�� �(�,;��@�4�d[v�oM�C�L �L��>>pD�H��ڍ��9�OpVU̙��R��Q��=q�A{�dgJ����ĸ�~h�76^�ǉ�:���߯&n,��$KB�wt̥��kd��џ����^y�[�����xDǖ��1c7�?|���o��@�!��wt?�}�W��4��������f~͞�R���4��|�?1	c5��]� ]J��?sN�v�c6ݨs�֩C/�X*�}���&�5����Ohة�b�m����Wkn��7[��.��v���g��4�tǧ�˥�Y��0�We%W�Y����&����~V��0���!!0�FDF /���z*q��	��A�},����1C�~��c=�e}�f�(y�D>��n!�}~��g6H�k�2v.)�����ŖRn@:��Vn>��9|Լ��ϧy�&��v6Qㅚ�/gn���1}���_Hq����|����zg�?tX|03��x�ņ+Pn�8���]h{zg��tਜD�Jd�?0B��z�Dgl�z�������6t��(GR�PAxȴ8w�#P��S�u{�"�5�3wd��u=�'AqGѭ6�~r����
�.�o�A��9ȑG7�!hW/��3*�h���v�/B�5�
	#�)�Jb~%O���d}1+~�+�/!��ed�l��IO�F�3�G34t�2���w�h��7�=�;��\<ֺI�ʣ+�X��b����X(���q~i�ɶ�}�3��54c���U*�ȓ�Vc��&���j{$ΐut%F��G��%�W@涿6�T���
�U�%�.:[��͘�:Pvvw�Së�>R7��]���3`cG�vc�)�BX�~bj���~�՛��jӰdV�m��.�Ϗ�g[�?��_�<�v�uW<|.��C�o@u�^���%�]h�V�}PH�7�$"�r/x�G�P3��k:7˕k�E��e�9���c���9ԫdz*�U�ͮ�w7W���s47��/���0�C	 -�0�=q�K����s����a�u��M�mP��_V7�TE9��`g��˚d�c%�(�2U��f���v���1�k��!��|Ĥsu+���St��h��0큦r���W�3�5�N�Pk�!��c����6�E�	�\���ιGy:�Z\4�E!9r{�GO���x�L<��0���xl *_�w���þ}���ssT�tt%B�����DU��������8T}^ro���Ƶ�HR֟]����X�a�+T-��"5����6����ΛS���#�>&u��a��#Q:��'I��p|��Д7�^�$�j���}������'��as���)��X�ko�)�����1�gpń�{�7�r�)k�=���1Ä�^���cs!71�c��Y;�K���3t�T0RϠi�:ծ6lb#3��#��T�
F��������N|��:�*2���hz8��X�0�����,(��~Lap��C�>�"Z�|����-�'����=n���}�e��ţ�Tr8.�O��$�#0�s%�ɼ�*;=%v�8���6Ӗ�O�P����G�D���t-����]y�pl0���s����<)��z%�b|i�D��&y7SM>㼋[������x�� #2C=t<d9��~=�߿��X>}	~�#��I{89� �Q�a|��{�q����v��@�ihŻ�w����r�Z�"�y%��!c~�����gg��K/�4J�@8�T<�m�Ni�t��*���_V"QxH���a��P����Kc�鞜>y�i������|���;]��m��`'���q���%�
t��:p��^�	\⋸���v�ONFm"�S���k��ʀ��<7k��Ql4��{
���t7��T�\��5Y��xwz��[�k��닙�5�H�(o}:Q��E����br^�P��}�͎���Q�X`kE�MQh}�}���}��&qk�<�J���*y�1�l�Ow��惡�M�wZ�4��g%P���]Ae���Oc��5�v�z�)r��lx�-���c���꺽K2����p���a^��]O���TPOIP4n7},��Ë�~�{+�c[�ަΨ�5{B�|/-��K�gƫ�n1�&C�����O��zM6��}��C6�\�-�+�DEM��Ym�ax��������2�LV;u���P?_n�c��Ґ�@
�,��e��܇3���?w�;�)��j��ݦ�u����#1\����cId��Ӻ�1;lj�k�8	�t-��N��Lf��$
�P(��a�Q����ֻ2�r~f!a�a����%Լ%<�7�H��g�w�Y�,S$�
~S�ʦcSЗ�2#$��غ|/_F[�F�c��䋻���7��s�;pǌ
�yx�
O��HkM�@������|EF��[ K��r:��km�	8ORЅ��{��d����Rb�0�/r�G�dM�=}��)�L���C����<��t�7���R��_?8�L�)+�Sq�Ӆ̙��9�>�9��=�NL��gZ�=q�Y�O���$=Ϫ4�r֕,ܴJ���f�nys���SrB����Kh�����pb�C�<�Ba4�4hpc6y(
@�DN�s�98,d�7������~�'j�Q.%��ש$����L��O"�i�4��b��ϳ�O-�;���'䆗�O�ՑF����C?�������|z�Jm�1���d�)	R��lo�ǈ�II�/��VW���_2}�Nb����oҫ�<@�X��?��
�,o�ڗf��;�uUv��ɷ�}�}u�W�vБV^|�4#"�^������&�����x��hy��s�p�ߎT�05Ë���H{��ŧ2�k`�F�׈��g��NP�"=|�w�mT��T@1x�R��A$��`L�[!R?{�6���TJ~���
�/��w7�t�*"�qR�c�ga��!�t:t�Dc#*�q�����d�d����g��������\�c��-�m`u������S6W)��t�&��H��XI���y1�7={���p��q�C0c.\o:.�z���q��+Z¨�LxQ����C���=��Δ�����Ц53�^�&�}��[��z/̺��F��l3�>��£s_�Uӻ���+��\G����Zs~l�R%���%����6��Aܷ�4���t����B~0v�'᪠�2�Q�/� ��W(	�/�#�-u�>�oN�+.��سT�ͣx���F7y݃��1���~N}.[��=sȍ��*1V�mts�s�x4f� }�k~��.ȸu,oTuT1����I�G_?/a�|ŉ��kY:��:/&��oxO[_%;��nu�Ny���Ps<t��3@��'tXh~5cj�QO�מ�f9�yp��ȿ�k~�P�+�``#��~� �×�yw�Į��'���ix��q-�Da�7$T��w�6bK� 1s���_|ƨb @=�������_��,v[]�d.��cY(a�����ΧE�x�s�LnK
���knRN�5%rR-���3;9P���-{�93W2������^r'�ﳻo���J}-us�h��7���{T�Z5ˮ�y:�����^f_7{ʮ�۩]v>'J��<���s�}�Wf	19���+/��-�{����ѕ�	���֟1��87���4�ΘZ`+¥/�[&��Vݔ��\�Ҳ%���K���u�9MG�\��h]=XVv���)�Đu*ܸ~Ƶ��"�W�)l��®I2-��� |���p���V��	����-�Or���_
CTg7�r��U���#��O�D��ʛ�������rν޽şm�[B$o!�h�F�]tu�dp��ށ5uv�gD���,At����U��9����i����`�k>Q�86��Z��m�;@�:���g%.�`�q����;N>��S����M����iR�w����ww/�mD�d���@W9J�Tf��nd5�1�m�Ng�.�Prwn�z��w�{*ت�����&��G���ù��=]Е�b�.��vcExQf)�2(�a�J�7Ej�Ӷڧ
��ޛ�[��t���}�ޯD���JYKa�@n�aY;�ڕ�]�Q����q�|���$�#��M���[��3DZ���C�dl�8�</�y��G(w�����O_�����=a߅���\��r������Bjq���i���$�o.�5�Tev��᡼=�z�R�w]a�|gf �O�����,�/�`��阙���h,
�@Ȗr{����n�e����˷`�jYf��׼�A�q{׌�۶DSF��vN�M�o}K���=ۂ;��龸/���oimo:[�d<�8d�`h����p��R�f0�Q��Ս(�N��f����,��S�GAD{40=@�C�P2Q�V���qKk��G�"
��ȷeּ��a�f�,}�)�M=}����Iw���S]:�z]����:�Kz�i�a��ũZ{����.�w���q
�� 43�&/-�;	���w�Y��]Z!X�H��2��#ي�i�����7+.�YQ�Hm����2���@�3&���v�����eW��n�;�յr|�!�8��t�&���RԄ�D>��Af�E\N�n�Q��k�ꛑv� Gu*
����]u�\� h;EM1��9oVX�*�٨��qug
LgiYE�v{5rA��)���n�����p�n�\y:�ޝ�K ��6��[����	 AHt�+#��a))
*�C!�H���3�On�_Î8�:���?����!1R�@W��L�3�# �! OH���r�O��q����3��~Ｔ���g��<����+	8��C���������OOo�����\q�G��g����ϼ"qR=���΋��1@��2� ���� 
$���JB*��c�7:γ���\q����3��}Ow�Ȥ�y��j!ܕ3��ȇ�d�ac�>������g]Gl���������8�_Y�_���9�
�{r��p�"�
8d�`Hd+��RaFQLX��=�ns>γ�����>���>��>�o����<8Z���t������ P��Ba2p�8 i�� 
O�Q ��"@�a�#H�$�CG�k,'�	��((v���a 	�00�B��!8RÞ4�d��H�T !�_��<���˽z��z�x[�K�2���t���WJ��G[׽��3��0�L!1p2��(� �0 3?i���U���w&'��pտ�N(ӊ14���� �}�(�����;��I�>�x�;�Fu4����$#ԎR���5���%[�&�^!п�D�zn-V-'��=�s���m�;�g�w�c��M��w��Q��9�Ug&�0��-�ˊ�71;'�;�v�̶��=e�����霾��ńqSɯ�U�ݮ�񇥐>�Ǝu \(�&��*�gЭ{/w�=[�2�m��^|�DIp=��[�Rq"�18�op3�Y.�����3f���?k���g��t�"���Ƶ*�n���uy*����^c��z�SJ��εO�۰��f�1�J�gl��e۬���[����ջ����.�^w�5��ݧlU��D�g�i\�!*P+
?ߟ�g��e1����P����� ��Q�]jn,��lx���=�H��ՂҲ���e�~��r�6TD���b��:2�
���)g�*���tN���mT���BB��!�Z�|�6�磚���ۛu�o\�|�SŨ��۲n�NPw�h8t�Mq}Ӟ+=�
Vq	�F4�����I�����
��&�<` �|�F�2v,t��^T����]���)���`���n������Ҹ�����zŧ�m�vm������G����f928�?�`��$���w���pz44��g=A��I�`��!�}O�d���-��m�\�k�'X���/u�%߶]٦�8e>�6�6�[w�7�V���,3>����3��#|'�V����LH3W����,�	"	�(������0ur�N(
�<�BB�� �&�_�0b�>��
�)��oeU��s����Ԑ��͏,8���gͽ#���(%9��A2��W�R3�'ջ���ًu$������/��ɯ7 �SI�?9D�.��N��?O��2�AU.}A���+&^�;i��9gO"OA����>�IH��HLt�z�Cq�t	w���N?���ѫ�v�m:i�8�C��j��sjD�����-�|�52d$�~��>�f�9�8���j8;�M���Q��Z�0�)�K(W���N˰��蜥֭�:'��3t�@ciY��ڀ�4+�I@�P�gcʝ�	o����G�M*Ί���΃+=�\䪿Cօ�J�����?�ܑ �J�}��77�]~�F��nFߵ��p}�e�-��=3�#lӹ���W�=�QhEn"����md2��+ן_}>�6�c�z4����l�X;J�Uv���@��.������v���QKW�vK��K��Xt�;�ڕ��9ӝg{���r����n��ˍ�(�-��'��&��b�K��w�2�l^*Gh�]��=m�)~�SLa��B"Rb��C"$���2��Y��ϴ~h��ʙ�)m��>ú����P��_?��L�y	�-ar��\�2>$34���ħ���Ӿ�~��!Fgi���cW����IԿ6�t�4;��=�T331\GM��CR�E�b߇{�}�Z��'$����D��d��t/Ant� G|�����a(�
��i���K0[��X'1���U��4�#�&|�gˠX���'�qt���y��ִx��^���3��f�\�ު���⣠����1T�be����Ͼ�u�=��!�T7������]?W0��Y�"4��"z�ak�)���֛�r|q���|��+��\��D5���������q�]��>R��|�0�R��/�2~VF�����=3�1z"���e���0�|c�ύ-�$	�!�x�ۍ ��.3ҡs�-Z��n��\�+l��B=]-����Aj������=����V�2��;=sW��c�]�B�2�3\����!g�T�be�ކV�+�3\0�'�r5����$�ܹ��>�:.Ź2m>!�y�ʘ���\�q���E/��,1K2�r�W�L�C�&�rkN�8]k\���<�n:)r&�-�7���J�����d��>��G��3�WC�Q���r!�Tਫ਼��<�*"dU��Th@Ę��GO�9}��Pa�T�v;��_��&�ת���ը0�I�n��/gul�ӓ���3��Ɖ�OL}j�����Ce���.�'�1���N�>W��u�����U�u��¤��3�'���ўz���
���0��0��_f���	�o��ݏT룔h,��Ѭ!0����W�;J2�uwl�{JKA&�>WFT3cj2cgx�.K;ƻ�;%���*�@R��8O�9̒��kVh��ت��$�cptb���?�|��m3"��\�2
��qw�5�����!D���4���/���7���k��5#{����F8���u�V-J�%wzp��m�<'�3���fCO���e^���܊��aޛ��Z�@�9�ĻbR*`�8�[LObG�����p�5�$,�=�'(I�7}z"0�1���� ��Y<$�,�(N�&��v��Nr^Q�Dfry�bW*)|˒��v_���yQ��5�>���G�c�3C��C��]C �]{ԝu�Ïv��[��ǎ������հ�̐b+�
l��N��2�^}fl5wc׸6}xX7�l�^���3���e��v�	�y�oLr��W��P\�ٔ�36X�!Zve�b��;`��&[+N���� ��'����IP�T�����ۆ�D�8�PIc<�W~��Ŕ�a�L���V٩s������g�*j�9e����c��X�V�=`έ�n���Śսz�;8n�3�|�>�+}W����Q>��k9��S���5��TNN�酖�N5�����P����4�e�Ք/�_=����}	H���u���v�^<*ی�=*Z4�Iʦ{[Mݲ�+%:ȼ"�-wC;�y�ug���l���{{wb�z޶�8����j��g���X�n�D����0[���Ip��}�\�S��V����.�E�ۓ�Ń�F͙�
���j�J�Vw /�c1�u�5��8zn��遈'��t���9�����)V��q�j|�cnS��h���9X��n����لM��3����d�R�? �0$� �!q��B"��wd� g��_/N�5�e��;�^�@Ǻ�R<z}#'�EDF37&36������VZ+�y��z�>�>M�o6Hu��>W}���K K�7���u5y���;i��/R�tx
��9����,��O��e�v%?��&V`��q��{h��T�����G��wq{3��X�F�܍	�����ݯ�e�����~���3Pk�y�m��Q�InzRqj�G�_}��U�Q_f�~��"����k���0���[+c��d����Lۍ㵝O���yLj2К�8�͗�;��h��+��Sp�]���`��96�Y�޳��0ixԀ�zFg����uݯ��ʋ=���'/�F�} �����cg�j}Q�f&�Ǵ��� E�&�e&��=c>����f�M5l3���!�Q.&z��e��>Y3��a0�e��#�WhW��t��+���m'�����_r��n��MOl�F�z/�ݮh�����n60T��c��:vⳭ	�˼�rq��k���_p��kKY���uw�1t�N����ή��krh'i���j���1�;68m���h������Y8ʮ�6/F����'8Ga����+%�a{U���$$)tRLge2�	��{� �`dפ�rX����������G`�����9�/>���Nw�:�M��HҮ|��]w��Iު��8J���JL7u�8�6�5Ǹu����]iY�0l~=ss�$)f����5f z�[)���3��
��3�O�� t��:�ę�U�B������Qz^�����H�o^ϵ]����{��u�c��,��dn	͉��2vR��x��镞�=��wd����h�7FC\5��*�weh;��_Nm�Jv{8
�Xm�WY$�>[�:�Q\�c���NԲFB��ڴ�bxǯ�=��}B�t���	b�����Y�y���B�B�n�Z�f���<*�Qs��3�>��iR"7��9����;�Y�¤T&2D��k>^1*.�C�0g��u���{�i�R^odK����~��|�O�y�8p~~�ݏ�Nnv�YN~��<Qg����:�jB�{f�NK~Z>���2�K�)8̦
v�h��ϰ�����Rn_(DĜ���D0A8��ͩ��i����Ӟ��J�p�}#Ȅ�l��;��%�ŵ.�;(���v�^ݳY������{�[��/߄4��)Ǜ�<���`��������-N�������[�:���2�]kU/�3�wT�z|St܆=�{�����>cQ�b�g\%�箤�U��2����M�3��.��E�!7���垟n��v����
�9B�VZԷ}j����p��l԰��{�T���A�y?���<��~+��Y���;���a�����40�&DNǹ?��q�@��}��u<�U�.�w�l��2Z��de��V(���C9���z�w�7������d�i��h��(�r|/���=�e��>Qn��F=5�����,q���(��p�˓�Q�#y8��귃�]�;�r��n�=u��ƧM}�u�nJ�)	ޑݵ9�9�ʇ-�*���MkԞ!������+Puʒ�r��w���֩��+�8���^+�l����mz}�WT�ҽ������ԭ[�X�-��g�h �o����~,��S����`�i�W��^ן[�<ne*���TU�	g��%����T��5��Ӵ�J�N�ׄ>ķ;P�*Z5�u����m���{��a��s��=p�/~D��(� �! �B@��χ��������?�6<�v�}+ں|�j̀�w��|>m
�<��nM�9+E��?o�!]`�5���~ͯWN�{�����CҎ�k����f�5e��|fӷ3�W���S��^LE����V���[_!v�0ḁ��/�w}��Q��ܠ��<��7�y^&��p��a/���:��mf$����q����P]����G�ʵ)T��ܿo�'�.��[P1�4WR
�Y�_.j���>�Ļ�^L�	�v��IF��̋#T�ʃ��pD��\q������S`��H>�M�e���VD�l�~��Z��\��[�&�@� 5�W;��uڦ��G)��٭��aa1����b�6Fty�!� ;��e���W��N���6�$J׺m�;~ņ[���ia/~�aƯGAw�^S�p�]�=彠R9]�dN���]6�=[�5��ӻY��Ξ:x���p묻M9��U3�^[�|���+�6ݶ����_q�qR�q��X2�Z�Y0�ׯs�V�%�+K"q��9k:�O���D ��hB"`"w������«�>�i�������Z+g��+�u�턇=�/4lݛ�ժ.�P<��/FTm��� ��V݌�M��嫷�^8_T�R5n���S/i/�$(I~�@s��[���+�;7�Yޖ���ϔD�l�m��?#�������~�"�����~��g����m&uE�ۅL���u��#2=P�F�J=K��1Â�T��9)�����bd3��=�������[_�yՉ��2�_9:#n�+���#����ͫ��ۃZ���iUL{�7�+L�u�m�
�o�\�M��X�F-�g��T���f�>{*I�
T��Or���v`�{�uH0mMEL/v*�A^�0)\�4��Ŧ�
9�;�-Z�Nu)��Ud�J��T��pYa���Q�=�1�b}�+ �׽��<�h�,�!,��"$�9YOSw��T�pR�2����&.#Y9��@
��&m���@���%r�Yt�o@��^��Q���+*N�U��Y�9��]��ǎ�����!z�=���mf�K/����k:�C�N�n�W�!���o6���صEW�U�ь|�V��8:Z;"����]��N�B]Ԫ,f]�;}��]�ZxSW�6���h�KT�@��&_��7���ʡ���� 6gr�Z�tQ�rCS�SNX@�Ų1pUh£ݎ�l�B��*{��e|I�%(a��9%���CW|G��i�|[f��~j���sp��Ծ���U��e(��'��?���cE� ���[.[#[�D9-Q��@4�q�s�<�������Gq7Wt��k6�n�S�u�!K��4D��r�a��v�<C��ىn��*2:�7I�H=�s$m!;��Y;��\!���۝��q�^;0�e#�X9Q�ӛ$r��gG5Ӵ���)-���HWCxM��+�9�Y�)���l��e��E���re<�1�^�e�3l�砑[�'�pX
dw:�b6��{���:�t���J7��51�J^E�VW>�+pT,��r���])'׉n�T�T��/#yvd�꒟�U`�!�X�)̘��
�D����C8��
�i�
��]��2Z�-��@���ˑ�zr��Y1OBp�3���*N��ѴmU؃�����5��1��I��[?q��m�e��4�T��+̫��9S����4	���Ƭ5]x�`�V�.��M�+`�Y������%`�v�l��oTS:�2k��글�����̘i�jm�SeYtT"r���	ǃj�X�ũ��+��R��q�0�kVw�$��d���ԥ�D�i�P��wI���X<kZ�J�,�ɺ�Wfay�����3N[��I�����,U�Ԧ�0@��ZV�c ̭�jf�W%F�,6/wϠyt���&�r� �u�qeD�ۦ��0�)�Sٗ|-�N���PO�ڳ{�U�iH�&m�[\�l;��Y�Gst{�n��f%i;R��zn����_o#V\��w{�%X:+bT*�d���m�oIg����(P��a2�&���K8���Մ6|Ơ��ub��+7u��z�Ҍʸ�3ts!��e+F%qq؅�y݀�U��p�ʇ2E%���{�8*��GLo%SZE��'�Y���b�J93���r�m��Z��̻�V���%ۄ��!t���n�\	٧n�̹�gVJ�: m�P�4S�{��#K.�}E��.��T�d��V�Cr���xz�}�jr�⬝�r7T()2T&� ��E�asV[��6K��[�����;w� �\�S����9��ݍ�ٰ�m�f�n�])��Mo8,f�?v�f��b	m���2ҒAvӫ8�F#E�4C!	�	��sg��8r�l��ie�\�w�-wv�e�͕�`�����JKf�w�9�yۨ+-���m�]{��V�2�w'�N�7n@�Ob�:d��i�X���J��+V	�� �d��H����������������g�_h� >X��йeB!+�	H����W03p�77>ϳ������G��g�{����rs�{ �\a���.I�#"bpL�P>�bi H>4�Sp�ED���EEG�����������<�Tw��i� b�Ik=cg�!>��yXd��L�1˛�����߯�����g�{F��uG\�>dd�$�88��$0�%���  )�J$���Ϟ���ߏ��������隣{���9�Z	�"$HĖČcR$BKl�8�gۗ779��{{{q���}}f}q���� �p�|K��&F]d� IvٰیDɢa\k�5h�Fe%���k@��sY�%L�R���SC�	����@L��rf[�"$W"=fM&K�5�*0��Ph��H��bd|�ͱ�0Ȓ5{6��	�U`RR�B&;�3L�Q�6ۑ��� n���7KaT�t��F*b�b�i�T�S!>\mv�`�N+h��C����-#����vB����e��AFj��}u�.tT^�Ns���F��`�y[I�\f�뺦��"A�D:2��,�bt���G�D$�!#AD�:�4줼����lc2v���37.EZs8�ō��h�0�~ �����Q���{�OQ:�\���]TՠzF�ײZ̽�\3�g�Y��{}�2���f���ޡ�f��pB�~RSw����ԫ���/GU��W7�1�m%�n�����v�����X���� 5@,�Mg�v[^ގ}�kݬg)E2*���W�>1`x�˕�/뎏�ކ���F=�r�Ik���d� �����1z��/EG���|�p�׽=�7�MGP��.&�-���zƘ�TS��^���wj̊w����-�`�i��ն���� ԩ��Ur�N�_���hy�$���-
j�ژ��3�`���P0��<H�*i��зR4UW��������O0�-X{��t��u[���f�hޑ6^OZ��c�-MVr�����Y�ɖy1�D��l;��J+̋qcl=\IS2oHu5�]km7��T���AՎ|�3��n=��r��=������m����k��dC�fs����u���ym�����'�{	?���A� � ��TJ)��n|�T��Mj�j��{v����ջAXY�ʚ�ى9i���=��@n<���n5�n\�$�6L�pX3��Ӻ�S;N+�q�\�[�޸���2���ÿ�[g����S�u �?Z���͛�u=w�!�c<`���F6������ܐMd�����u�;,�N��������(��eql�2�Q��0����o��$lu]����o�8�BE�u %��w���)D�@`�y&��v��{y]c�)In�u"N_�qq,_�1��/�����Lk���\�����Z�����,�S�Kf+��
��?����HW6_�ir}_S��\`�x���13�%x�k ��;�d7��1W)���oLE�ت�����_�X~�=�f�b�N���o~a�}x�q���O1��MuC���;�2��m3��{~�Ws�PQ��O�uG�o\ڴ�p��6�)lc���F�m�6v*�z��U����2�[v�GV��ut��[�)���1�ʬ�K���5G$���\� 58^��;!����:���/����r��7���1cs���˱�X�ٷ�R]�C-�X7l��1�mWu�u��rj�X��T�W���X�	�2�Uvyp�M^7`��jO�h75W���N5�:��r{$+�p�ί����_^�4^
�b]�%�I���4hܹff����p�h�)?��q��s����� ����9�M�ݰi�Vkm�z��v!@�ZC$��-�0�)�	+��]���0��GHl/��M�h޿a �uV
XS3�enx�����Wȍ��}c˝\���0k���6k&Gk�*�bS�ݵ�ǝ=�7����nl~�S��;{�Î�O-�}��ޔM�������՝��.j�e>;,_�<�5�·]DW����N�����&8	��W��9���&��`8#%����6�[�K�G<�G�Ny.nff;�9R�t��a~�6(ɜ�j�i
!~��//yjڷ��lT�كs���f<��x�G5��z1sx]�vO��o��sKpU;x�2'#2j��Z�F��I1@ဃm�(>��~�b�}.�r�N�X=�����g8J������ؤ{3y�4���7n���d�k���"	H�!DA&���3�zL��c�v�跆�X5�)���͑�#�ɝ�g��N�<[�F�_s�[�>KT�5�� ��~���ޠ��H���"��z�J���u�ޟV�%A�
M���4��:|h��{>u2��W'���Sx�e�M��2���Զ�k�ȞI�U�
��t�F�Rwa�Ur��SS|�ڽ��T�\����@u)F��X�UݥN姀Y-Of�� X�(d��^�U��k)���&�(7�B��eK�-t�x�Mry�x ���nIV������Y�/�ש]W0<�(���$� �����������>n��b�`�]�Zӏ��8ON?��n�f�Ul^��4o �5���ow���[��U�c����{�y{��%ZM7k� �������C�����`0��1�R���=�RWg� �n�{C;VU�I�.M�*��4W^��qQ����]��_���G���3���6@��4�(b߮e�7Ρ&�8��2%�}q�����;��y_P��;���}K��;�#�|�1B�
nM B��v�	t>8�]�n��j���/�ɡ�� L���:�0���gh�d�"�F���-S�� �r0��4dz׫�ͅ5Ԗ��%5�59�
Lb�4��������r�$�tVH Km�e21h��*P�њ�����l��>R'��lg.���u*T̕�\���\_J/U�W���|i�<����ݷ�=k�]vdT�ʱ��L��zn2��[�I�ޏFn7��e��lR��k٩�v�o�k�<L��GF��KYk�Xn W�D��0���xZ��UYuٶPa�
o7z�Ϯ�t
�f��y#-kĻhl��|Bu��̭����h�z:���I�l��8��	Ě��S7��b���v���͒�2C����r���L~�^O�.z�Ԭ����2��V�+�Ρ�[P�qXW5lÿ�,�sRO���(�����2�aK]�6;m�f�r��'j��t����Q�q��{W��=�fb#S��0i�k�F-�{*�K�V1C�K�Q�X���ylV��K��&ɺ��(���uk(Z���ԕ�WLʹBkG>���3����y��DQ`@0&���B��~麨��B3�1.�w����d����" ��$������S{�3��k���)q�����|z�'�}��5��w>~�E��z��Fֻ�9G��rH���J�̠J�±��Ur�Ag��_��~Ku��z$��G\Z��5�NyqEO�U�{��ܳ��Cn���"�Ns�ˬeU�v�:�g_�;�2a&��Nٟ��#�=����0aU�n�	m�z��X��J��n�g��1\hN��g�:7��Er�ݮ����D�GjT�e����m��M1s�r5��c=�R�R"7�#�LY4:y��϶,G��R�z����ܟJI�kz��2L�r2#/g�+��L\\�U��;��a wYa[����	�g��K%�n�9�U�a�6�wx,���<VB��A�>���-�z\�I���*aȀ�oo��Ae��qֺɪ�k�rۘ,�B�soo��w!�X�\��&M�YU(�VK��� �-���wzʞ�70���v��+e��nX���ǃ&q����[�΂�:���fka������0vs�rF��z��P��F�n����蠔��'�v����r��+�Ȋ�{+�ZZlޘQ��G��S=j�0�i�.��"֕,�]��GK�w��<���}��\��xI�o�������n���Z�j���J��U;��jR��zd=e]uz���r9�(3ZqO=gYv�wq�ꗃ��$� ��\�y�F����}{��%.�'��ov��z���V~��a���EF�Z��.�B�z������Ȏ�gnʘ���n��^~���<ג��X�#@ʇ'=J��T҅���3uP�D�{�|�����a���8�bd3��e����[�7�R�9ݫ��`Ǧȷ~T��Q�`��W��G*Z�G�G/�� O�s���y�Ia�>S�|�x����{�Y�	�%�˯˪��g}�8۞u�#�`WF_�:�ku�^aJ�/e�6����ͤi�a�[	�c��u�zc��].��e��ٽ�3"V�t����<@�)�K1h!�O{
��ڣkô�(w.���P띜f�s*kKC|�aÛʵv���� VwQ.����I��=<s���#�����q(V^�.���^��M��:!��mDH����c���g$�W8ZiVWn�ȪI)��{�y��q~'#�KQ����ȏf��f~Yޢ>�)y����{�*k6�	(�[{�Y�.��ޥ�f+Xn�{s����S������5�y�Q����,^���p��q�_wVa�Tܻ�mN�:��@�`!dMijp��	1�5�iodFwX���౽W-�-��2����_N�s��L��3��%s7��_+E�yLz�}K2j����7.��۔N�=qf�"}��5(�U�]Q�|��= ް��)��m������/O<�FI�+�D�ݥ� ����N$�U=�kR��w�)����~�$����������_�s��f�ZU@J�RY+)��6��s� �YxG(��ʠ3��_�Ng���v�Ғs���ϐ�Z�n٩��NSsl�4������v�%B�@�ȫ>�W��ʐ��`�ڶh��ى�� ���=Gce6`���K�`���ɝ�c3�ʔ��,!$6�	�c6��k�T[�t=�x���n�KS:��Iw'�!��L�-r ��ݣ��+R�.Jr��(�Ji�J����#�S�����6�Ț�Z]rL�����+��d�F��4ܝ� A`@"	T9���'����\��<�=[����L��~�.�U��v\�ښ�̩�ۅ���Z��M��9�-x@Wca�l��y�>���.;��W}���u���&wٞ1W�T�0�A�⭴mr��'�qU�x�l�N�pY��1,m���8��+��]�0o5�4sO!�
��ͤG[� aw�E��Ӣ;�g�k��,����W�<�M�VE�˳f�a�e}�5��>���5���5`�������+t�p�}����[/=��`$����\ly������W������Q&ϥ>Vȼ���PoH<s|���k��1�s�pT����&�5����{B�R��3z��f3�g�B�:C=�2��H�T�� ��B#lL�$N�2���+���3�3�P S}���<��[�B�E�h_��.i2�juҜu���?M�L�����`}*��|L�y5,[��f�:Pӵ��T�f�q$��c�s>�g 3n+c=]]�qŲ�D�{���GU�E.�w-sݠ��Zf��g�2{�A"(�A]�{�Y鲯�T�\���ƃx3��-�54�d4d��$���v�����:g�)͘�����9�؝0<�ϰlg*��,L�3L���]A�H��=e��&a�ޖn~��G���X����8���K�5���ypR��Z3u����.���U�G�k�5������|"9�S�L��fm� I��e��F��H��U ղ7c�����h{�X�]PA�w[���^5�][������ax��S�{�OF'�!�g�e�^�L����*Z�.�4���.�yydw0��%q뼒��D!�kPwb:�s�n�
�1����硱���D�w_j�S���<��v�%}�!��I�A,��x�6�Uޯ6CO��oï�r^�c������9�k!�
�˭�%�d�6N�;	�X}�wk�4$�����"�ܻ|��T:a�E]\]q��o9�Z�!�k:���;�M��<�*�Y�}����3Rar���߰�'vӊKj�%�=�f��Ȥ����KwqCXKX(uG�<:�n���h�
�����8�ͻ졥������f��wY�!+�f��8����A����j���q��%�-ͮxo�Xw]�T�t�ѯ�J���nH�[�@_7����P8��+5<�k����2�<��uo�]ǳݬ�q�:cvV|����l Xi�!��i��Z�պl7z�ϱڒ.2�]��w��ۏ���4p�v�d8pv����4�{(�QI&s�Sk��Z�9c�"Sm28\W[x5B� �:��]�Ր�^Ƴk�#u�D�W��ިO]�Î���vTG���H^#<muź�LvҶ�mp�������l*\�le��7~}�����@���Я�R���tÊ���VA�Ԭ�8]\�ʖԩZ��p�uv��P>{L˼��Q���41�ւ�#�*�M�9Wh���ma廗���jIG:	�������s��˧��?�!��;�*�]���+��9b\�!ض�Wg�6�b���h2��������{�0��x��g`�7�]����feu=���K�o(��h7�P|@7�a!y�����4F� �~o���*�n!,RT~2�2	Ov`��,'�r3��8`O�7�k�W8J��3��[{쳐��H�|/�rϜ��2����n*#Ug X��wv˕��u���{Fl/*j�u�l*fĝG�Dx�("�C�%ۇ�����Z�)u�vv����)>y��F�˙�/5�A΂���p��B�� �嚉Gw�5���ۘt���n��zq�L���
2F������=��C��ܹGu���¤�W�a|v`1:9o6��ǵ������]K;T�Z�鸕u���Q��t�R�S{��k�[�����h�KY���:�4/h�!��)��v��Y�#�⮕d�o_CO%��n̥P��g�kVJy�.�����T_%2Fy���|V���S`|U��Ǒ�6��REJT�Β�M��=^v�ӝN��Md�7��'��'0ee���W[��ڎB��\�]h�cf��e��8�f��2]���j�/�|�a|*����uػ�����"m�ubS�t�5��C�Ψ�Z�k�0~�.���K��ب�7%v7�sG�)J6p�4�����rۚoF[g��9 ��C˹oU��K���\�"���o��ϗ"���\��n������P{���*�!Ȁ�d28qb��rr�L���ӊ��e�u/�29Yg�^Z)�ZV]��؅����B�JDĖ#0 ``D�b8���8���!	�-`<z|~=����������o��܊�F�9� ���o�5.lv�L�H0۔ɗ�D��	U���IK�Hc�7>��������g��f��|128�,��0��ԕ�rʓ��|�,L c��Bc4P@�ZP3�D��D�����GF��>����f�|�>�n�B��1$2֤'�ȣ�H@1�K.�e�f9���Ƿ����_G��g]-�
cے ���c
p��Isn�@ᜬH�]���F!�� "�^Ƿ��������ۏ�������{�׼�,�e���JP�d��� �'��%*�kHl�,����q���������}}f~��Pĉ��I�XD`y!��ے�e�w��	66Wz�nD:�B0�ئV1�+�(�"�� ^�����خ,�0��珞�k � v���#�l��Q"��Ƹ�
�3JR ���V##i�$�B�X�"D�d��H1H�Y�Y4f��d�tJK���+�v�\G`6\�9v����g�ZI�U��T�qT�;����=��+1���m���8HS =���ctP��ϗ:Ɯ��6Fo��	#&w�t�D3�~~�7??��i���HϖqS��d��zϴ{��X#�k��'s��wN՜�}�Iߥ�b�w����+��Ϩ6Br#7f�xb3�E���{3=�a��[N\��"`��Y�J��s����^�x>�uR:�QE����J��
o�ǰd-�g-[��3S�9~X�7�3��˱GG��z4U{��Er/-Dc�;��"��g!Qq93P�%Nf:�dy(@:K4f��g`x�d�U{="2`4���&�Zṩ��{���u��ю7�;�v|�o����f�)��葉j�1--�b�]�s ���w���)4��g������3v�����5��C�Ɉ����/3��e<�m[�[y�agu���������8�kT���^���z���BHrhT�V���\ן��Nrm
S�=u�+	���W;=���Ox�, i�aƖ�V���f�줳�E!e��8����C�.gt���l���ߥ-���μΥS5jFl��ٝ&���Q@�� ��j�ul��3+'�Ư�_��T��o�
��եo��nf�+�st_��hK��_�W�^d��
oOv� q^S�-R��#O=_1�UsT���q�!��1����MsN�xzW�<�#C�*'��)�
\��s.��z�'�J�'�g�������r0?<�lг@�����d�]J��=���u~�'��>6S~[��N.�m�zx�6~�������ֈwpӧ�vۗ�� '4��}�9�^-�e79)���<�#DV!Tܨ�0�קr��U�Xˋ�l�73�Rml���wNoM�\lz7`��cN�E:+��D£q)��v���|�UQ�����9�q���a��)חm�Kb���N9����Y����`�ii�����HX/~�Q>�d�Т;�ΐKU�g�S�d����9~y:5����)�Xo��JyI'���]`ԞT�2�m�'3^~���֎�O��l�^��RE�$�o�V�77u�?d��irܮu�V�'}R��K&��s�s�^>X����p`O:�
Z�	a���׾!�gv2��wƄ�n�1whKFXƏ5�Ö��L?`L	@��8��o��yqkKM=7kѣ�w���e$b������n�Zi�Q7wͧp�����<�N��g	�������;Q�
��%�K��L����ŵ�RL��n��Nv�W�t�z�������'��U���7�e�G�ʧ[�wz�Ǽp`޳�d���z�x�I۞q���R �s��\Nc��5�h�Ec�[n�v�1��f�
:Y� ;¿U�ޤ�	�+ّ}��7�j1'2�-���/��o�v�P�4(���}]��%�-.��xo89Υ_��W��-���Z����b�7���h�i���a����Gt���M��9-����w�����t�����Y�;33��;�3�O�O�o$/A�����}Gҷ���,�\�����d�O[�{�tv׸୴��b�������̞��/�lr���b�ArY�Ũ�duKꙘ�N0��c,�w�B��A� �33�Mf�NrׁZr��@�(�j����@`"��$���sn��Y��3;��R�9ۣ;����d��w_ugu�.�6s�(�.��[�QƢW}�M\��43@�{��{��yÿ�D4?��F�M�6�\޽�5�.�ӣ��۪̞e���Nk�����7U�M��]آ�Ʀ���s����v��(�7
�����zN����3<ܳ�Uz�Z(]���5�D�\^�K�z\_�a�n�<D�N*C��^�1��Vz6)���'3sP��{�f��oX59�ي��X�e��,���H�1��R���M]�Y7MC��8�[���Cȯ#�꿶���w�O���+�ĦԥJ���0��~q2��K�s=� �;��ˠ����ȍ7w1X5{�XƫB��:ņC�k
���.,��J����2;��[���Rw
{��\O0�����e]zߏ��>l�Us��q�<��t;���j��d(����`M�?�l(��D�\Kղ��Mw�Bm��3#�b0--1�Tik�[�!Q:4A��U�Flc|�/���[�$��v�
�K���OeG,x{���:m��t�o/�7��j����ovF�8��ssn�fh{��S��}i>ܹR_ #�A"@���ٴ�sW��=�+�߲�F�$(��%t��y!��DHgͨ{�
�)���B��ήb��G��P\g��-���:��y+��0�I�|�|("�d;Ƿʃ��#�+�����0��s�z�,��鈖��Hv	�p���7�O�k�X��p��o��6��gih���,ˎTB�Ƈ�+{�w�8夂D�\��xYWܣ����H��g�p�l<"3ݛ�//�ջ=;�ں�����_R�n�W+���L�폽����l=_u��I0I$G�2͙��ow��uH9=���4�G�a����u)k�K����K��9�e���W�)�3��j�,6U�mQ�cQ������=�+�Z���h�3���co����Ř�{K%��#1QsA������s��Sz�(l�{�5u�މ�)ф��=����
^�>n��nP��|3�B�f&�zM���^���γ�] �3��Q+n�Lf҅T�����2����7�C/��^���:����^�{(֤J�7*�J��&��+&�/�&���ں�<XC330�Jte�A9o�n;E����+�R����U�ðʨ�"�?^����F��0`sh֞�����@D��MQ+X�fߛ1�2{��,��j���&����������4HNTHR'�LEb9�)�� �3˺�Y��O�����È�ޮ�38X,�j�����S�7Տ��s��J�h�����.�w�5Ѝ�v�$�֊L�d
nۭW����	*�ݐ�p`��.�%d�����ӫ���cff�*Z�U�>��W��� aE�F���9��c�����z�K���[�`}"��6�ż�
�՜��2����䉝EHs�ݣ�{\Z=��i%����CjE�I�D��H��RD��W.�L�;3kw3s�®v�<l�u�r�q����Mot�5�v�[�'f���TMoH��jw����9�(6YK��>��g���Z;��{����A���(=�3r�� 6��4��6��lӭ؞I���$��M�.w��;������.�EJ�i�W>g�iF�M��([��:�lP�f,)���=�=&�ys׫�ढ़��Zr�;9���N� q�;���v��K�iڌ
hς�*B�[h�-�[�ئ�)��.���5!g�D��DA~�[:6ߵA�w�o5y_@�|�P���e{[-��d�CB�I�1?ڦ��~7����`�y�0�%�)����O?�-\a�G�Z����і��jr�6b߽]��&}Y�g{�C�N�y����,Y���v_:��x�F��稝�Cr7,"=Z����v3#R���>��u�9J��ǂH���=I3w�������Wd2�|������f��Sc�g�cD���z���g�!^� �ě$�r�i�`\�8�W;���O����L'M�l��$��I�{g'MDb��Qb��vu\�4�7<XG����޴�_S���^�u�{�zt��Y#�vc{�7+�
#���Sc� ��ʣ���H�h�^����\Ϭ�Na��5�F���ד�eyq�j�z�X�Pj��g�ǟgٯD =���_�yw6o!�mL�Л)��n��������mő�q�uu�G9q�����f�����&P&�t.��I���ip#g�})���e9�wx��huۜ��Zy3��ۍ�)e ��F	L������bR���3��Lvf���Q��W�]<��\u����h�@?�ju�:����q�z	\lv�Kz���@�3Ү\���2��sd>�������^]a�Q�]GLf�q�on�p��>[w�@�q�^6(	<g�vzz�O-��c~pҮ4'^�Nv����9S���Θ�Y���E�	�� }�+����wp����0r�:���9̩�>�}�-3|J]�`%FA�>���;}�Y�w���$�|��H��LD�{��傹*� �H<��U�S�I���q�;r���@zU�LB*k�/hVo�v����o!����3Pe����]r��Q��C�-[�Q'NhQ��黩��-�SV��� o(;S�F��" ���u�c�����4ˮ+�&�f,�Y��0�Jg�ݝXp|����ia��]#Δ�I�۝��L0:]�2��6��ܻ���q+�܁���#5z?
�>CEYn�N[����Q�T��fZ�-2o��	0�P)�b}���q�}h����ˏ��S�Ô�HP���W�R�FN�[��o���p��wf��uA��̷��}/�NxL+^|������&;�x��+w0�MTk<_���y�g�f"m�9R���	0=���z�Ǔ�ڍ��`��U@��d�5e=S\O��MP��9�4t��Bgz���0���?0Z�Z��\�2�[�\y��u�p�¾��})V���\��A"�Ue��o����E��sƩ���fp%ʱ/w�������v�I2�o�k�U�=���t;z��|u7�f�w!ݻO{�Z�V�=ä?������<9��U��3���s��0׏aծ��5��tzb�xfǨ,Ս#���Ϟ�9�U(�����~�������(��x���Ezrtc�m{��2��q�!U�٘�x�z4�үvra؂;�,�T����%�2�vH<Eh�^Y�%5���ۭ~	V!��Ki��q%���f��E��p�u����2
��b����˺�ɷ*S��,{%�FCa'o��Y�o�n�y��s��_�֟e�:U��sE�6u�z�����]wu�c�7���U.Po <�<�<��R҆e��-+��;�#aݛ{��Y>T��d?�K�u��6fe��~���=�q��,�Eci�7���z;���\���
�ѭ3E�MB2i�4�"����ז��ŋۻ�z��T�S�SH���%����!�܎Gh9�&��)w�	�8�1�;��ʪa���ӛ�H�A0g4�+Y�U�p���0mޓ�|&��03���V���q��n�7zӽ/%ޭ�p��&)���j�W��a�3�A������L�_��c��Z{�	��/�2�J�j]�뱠`�B=�*��[��kLf��57�n��ц
���o�iW\7
&�Ж�TY�T�R�r�fj:�zۜ�5^�m��/�����0�"�EwnX�䗯�����=M���yI+3�=]��K�"�XW�����ڼC�����Dzu��������Ro��p4�4qe"��C5[.��&i���w,���/hWZm�:�״`c��N���f��@�V�L��0�L��d)K}���L��xbR�\3ᅣ��3���hn��6�[�-�Aǜ+VBv�o4�-����r)�� ���սx��[�.��dZ�T�]14,EQ�պ��UyT�h�k6Q����lT�\[���ͥRR�PVByp.�^ۗG�6#�[]Gqˈխؑ�y�W҄:�Y{�sy)�4�A���2�H)Ν� ���,<e�����-�5t2|x�������;^���n.�5��#%��.�r�����}�;c�s�0u)9,��W+"���RoC�b�.�o0��g�zw�Eσ��;H9j�Wr��ո���ɇf�i�G��Soj9��LK���R2��4��K�& � ���wMǛ}}"�{�]�:�&��)�P�p�c��e����Zo�����c�\:5r�N�8�N�ϔ��W�:�n��Գk�-��Kr����TX3XTt��\P���s):�� ��u�Z��#�vX�s��׌�&3�0��|�r�N�eX�lTb3J�ax��Q�ض����L�a�/��_c�jT �Yv�؄�L��L��#4�eW�al�f�s\`ڠ�Sԕ�yI���]L�P��_�~S�#�:�
����xJ4��d�����e�(d�~
���
Xka�=r=��	��w4e�W��L��������Z �B�?�	^�kA���
���N@84�t�|����0�� X��+OP�F}j�]=�4/���n����F��y�v������Z�����C3�!YH
cSQ�KV�m
ôf:�,�Lj� t.�qk/qbw��� 6�N����6��l����;f�V��˞��Rp܃-�,��������C��y}��^w^ƣ둣լ�ݷ0rN�U��s+y|A���6����]s�@�p�,�y��;�ws�jtu֝p)p9�y�9^��3�|(��V�Mgf�1VOw3�4�Wzr�ǌVM�kH6����=��IZd���oJ�� �{X)�|�n.�����P>k�Xz�`����v���רd �,G0l��˸�v.8�\�oTo8!R��o���)�시���y�t�@٬Ⱥ�]C4�_>c�=��hi�@l��v�bNt��SJ�r��M�Z�ښ{��/�@�-�fìq,k�C�C�.�Ԋ-^��Ӷ���WDgE����Y��Yk-��Ȑk�#��z�_p�qb{O�5��53xc92�w;�.���	��k��;x!��y�Xz�FB\��dѡ��)����}s�Uӹ����G(����1+el=���a�KYI�wyu��.��g��!�v=�6v�%�R$AL��5و�-a(�T�YId�����k1�ۓ��Ai�݌شP��G[Y�t��"[%�k��MLf�7�.h�a5�n�t����N��,SID�&�Zt���Q8���oW`N�r�m��i"�bУ��������ɰF$S���T��Ы �Iް�we�@H)@<�S�4G�
&.*.&&&&&.<��Y�7Ӆ�{�}|�����c��\�B<�%E6�#
r�f`�3F�0f���������77777:��ɟg�a�}�'�$�q�� HM@� 嶄���Ո(J��K_�ب��f���3���ܘ��dxGG�������q�Idy0Y4�/���X�pǡ�Ep�v�S%%�����nLTdLLLLLddh�G�����8�ܣ�b1�q���'�_���W���#8]@ȝ�2�)Q��A1�
LddLLLLLldxGG���g�茄��Lp
Ğ��0�� A\n?B2�X�Z�AT���]f#���i��������Ƿ���������3�ڟH8?A�H�#I$h|���0���XB�-�хɑ��2$�YQ��^)��'�)���̌�Y�eX�tZ[K �#5���ʤ���mA1K`@x�h`��&;=wz���a ��<�[��l�v�V]&�!\2�-bIL�m L��E��ZkIE޳fNq��\�0 Ij˜��� �
a�q�r��H�/�k3��
�*���QC'fÝ�"kv�䗜�kP�e��Fp_�H2�ԛ����n�"�#t]to離����t�5|9�-��]���s��'9������ L	���]y�"��w
D�F���U2���[j�c����~��/s���O����G.5+�c�f �d�W�1j��k�'�\ir"f�uN���VD	���wt���ꐅ콆q�/����5��
W;��xɋ�k���X�lگw��Gg7�kx�S�{KR�m�5^2Y=�l{2��0d���>(��{��ɲag>	��ank�l��|�k�>a�ƒ��� v�a�#'#��~@a�������'/Tn�j�0���Tk������V���.�/Wm*�zm#���3�?f��|v���Ƴ�!p�R��֟+?�Qw��g}����$)T�� G�;Wr"}���$0e^umRF(�������kl�1>���dM͎�����l<7�5z�S�����*�'�Z�jy��/j���AL��~}\&�ǆP�ClV�L4�.*ܦ0Y�7�f�N:���@�97���J�P� Q�OxV^�P|��c��ѵ	Ǚαǽ+kz���&"!���:}SC3wݫx���"�� AP}�=�~�e�з�9�E\<�Q ���~���p�;~&�Iߠ*i��*r�,i������"V�i���>bg���E�R����ٗ����.���{ؼx�ҕ�S�ǜ�~:��o����3�^�ݻ"�w9�̜��ؾ�e��Uڑ�+� �\H8P�=Z���+4�k��ͼ\&�M�W.�9opi+�/P�Zh��ݟ7��vο�D\�|�6N�~Z���y�@?��o�;ux�q\��W��:�8��f�~�ܴ�(={��^͑��]�(�W����m]&_"N�5��z�g�oƋy�S��]C~��-�
{y*o�O�sWf���O{��oPN�in��v@8Փ�\nl~I��������P�l�PK�
{�����	.���-��}[�nɬu �E�6+i<��e���s�joMd�2qԔ넡ZK�
�4��9a��E;{��ùR:��'v�z� �U�еKR"6�u���[������\�n�}�U]do�rb���}Ht+��2�rC�{�/~�fɇ��󿮱QGqJѮm*}�#,�L���í���A��d���j��m�LGz�(�׌,�k��k�k�>�úo:��aߋT(��q�N�e���L��ʛr��Z��>Q�����"��B�D��c�� 5s.뉣uq�L��sG��=��^Ò��*/=�~[}�캹$RH!(�h X ~�|�z	���_��C�Q�C��Lߛ����#g\Lt7�*�j�Ʊz� VOp�m�gc����gw��o�=`M\ITy��}z�XQ�1���޺��G�Z�jꩿvcuϛ���uqk곦XL�Nf5�.8�ig��.���]��Q�}�f��ؚ����^0�՗�[��_ԣn-	⍰��������:�+�4]Q���Q�����1�!eE߷{��V�R����.�T�K�8�j�e`�z"�h��Z�����K�qs�UБ�:�J{�:��<ɴ���C3��"kY�`a�w�yw��8V��-�B,0����=�����-6����'�jo�n��Z[Gv�pK��� گg5��j8,��2���ʩ��
ü��A�1@�1G�� ԓT�9SE�c�ܣ��U���:�Xh%�����z����P�Mn�w��1�����to2w��PBD��I$�$���4�<�%@�u��Xӓ��g���gt� �es&��{|��lJ!C���y{����A0�{I�}���4y�������I��SP�ĝ��P��p[��*��]{N|3!���coЕۭF��vxh�e� u��͙�p�=��+=��1w{�R3u��
�Β"�U��T5�K�7��u�U.��p֞3��v{b�6z�-SQh ��/	�j���,���h���ⷯ=9�*d�9�Y;�B����,�v��ag����L���!U�g�Niۑ}]�Q뭂+Ҋ�*jh+n"��d
�,������&��ݱ��D���7��<�*i�5�1u��.�g.��t�on�4��Y��m��'�J`9�ɑ��H"v�	�TNa�Zt?���K������"�V�L:�{[�|��i�}P�Ԇ-���� �\� }3+�=Ӱ;�rưqV����4��%�v���ܺ�
i�%��BZ�wWr�t�q24~H�ApD *�bҹ�:���+�ePA�ɗ L	��fl�T���ں�/?���Ogu�D�g���v���U݊[���h�����b ?k�|�oQ�)��y�o�avY�OH���-	,�dY)j��~���sO=qB|}+썉�N/z�c�T5�k�9��n�<?�-{w�M[���3�PC}r�i���|�!Nc�ƹ���v��&Vwv�v�b��S%6�IO3�p6H�4�M�e��f�.яIQ>ov>����2�2|�fz�~gm�dA��sSYW����yF�ĸ�ww�9"���.��M&a��dU�U#�t�m��;���Ǫg@qVfs�=��y:	\G&7�g�)�)Mq�^�}��T�$(�m�z���*n�E�}l����_G�`��������G�-�ᰭEىw���1E�_^SѦ��`���Khq>�5�^+�i�������d�ۗ]����)=]0�w�':�A�ǟ�γl�e����u�s�\�^�0���|@�a#$o��µ��M����澗Kz�0�x�d�Wv3yܷ���a�XšǨ�7y���鲮�6��G��D3�7��$�ױ�9mրpQ���_�����lڶ�.�j�a�U��{a*黀��9�Ͳ�8�e��+]YjR*�>��+[����<͕�T�y��Ȋ��1|�yt	��8���xRM"I��{��"�H���T�V?�7/g���M�ynk�h�Y�rn/�}��C-�s�Cz:Ղ������]�Di��O(�\��Ϊ7`I�}T�ޯx[�����^����*���Q�y�<��WTu�hhv�^^)M�%��&�F燫=5�>�wfU��*ٽ�f���#��|ç��^�&q- �����9�x`������hҕw���h����>Q��n��bv���Z���+/������Qxby���Sk"7z��n�����7:�8d��q�Ƭ+�;3������w��_����u�(k���HSAc�z񭻾���0��M��|�I�u16�6�&U��[A�pgwS��#����A�v�o�-�l�ѹ���ht�/�u�;Fr���@��\GWuIX ^�&3ji�sgI����qT�K,3'�ޤ#ݬ'�����+�9s�᛺38��|�7�m�n��u}���R8c���j�#ǜ6�Ƥk��U��(�S��r�w19#�wR�^��{K��n9ż���>>C�p�ˣ���5�59���LO�[�J�g]K
Td'���^q�8�VQo��)L����ϭ������o�l]����YR�j�-x�X��������UG��<UH�۞�b���UǛLf����Ug�M�`kԦ4�j�w�;9H�=T�}D�)Y�-�T��&�yƂ�p��.�֦$>R����������.���i5&�"�;i�U�6�wڦ�2z�Зr��|i��͇8O������+����"�;����\D7-ʟE\U'��)~�^r7�<���c=i1�q���#�t	S�B�Y�W'?EG�Bǲ� ���7n�bI���ol�*��NQ�[��t&���b�� �f�\C��;�P�'���򳯯�5�։�ru�7���5����0�w[���]H��B�y�[��9���0�3�X�mr�g�=؝ó�0r���c�߶�Qa!���gF���:�d-���ʤ��+y_q�JzW]ϏR�M�R�TH���[��s��U2�!��~����V'\��6%w�����Ը�.�ʻ���y���L�ELUS\����i�@J���M�#ES��H�1\��#V��U1Q�w�^.�]O'�j��W�J��0;�jC��ث�O��k��ɋݢ(S/^I]�>�N����;����IWZ�6V��\m\Yͣ��l�Id��fn��GLm�"�q��a�ʹZѯ�������^Jt}�7Y�0����D{b=�l�R3��hV� �4���Ή�[+98�^�����L�t�a�p������
�o6,W��z_�^sfSܘ��V	�&�'J�o4]�Y�},�` K�t���%w�~�9lod|p�.�UM�]���]��}��pz!��gs͗q
���f;�5Y�xf��wTJ�w(�X��v:4�n� 
��e���{�����F@-7�]��b���'`�ٚ��ѯz�#/*���4��8���#��/�\�s���T�c
x���	˻7�wX���r�o0����a&HI�2@��q�Tc�!F�ɓ���'V�;��4#a���!�y߬׮R��^̑8�#������o�F���.�1����9T!��(�wadסd<Q���5��Unm$�t�����.`D�7�&Yh��:Ȫ3��;��YDڎ��o���	@<����F�w�LԞ&^WV��۶�`���2�C-t����
�d���Z��ʔ.��x*�Sd�B]�F��^n���7ػ}z}������F��fųo5�쳦u4Y�2���Ǌ��n�ǱU��'�O�D�_���؈��m�Y{�����B�{=��q�4��uU�}�/y�	L[��̑r�^&O�0��1?L��k�����V�{]l�O�čn%��і�-�h�cxZ��yO1�8{�����pZ�d�U�in�cwܺ���L�r�o�m�5�6xZ5�����ӛ�<� 0����և]^��M��t�#]��ǲ��r�K�,SC�wFsy��ڑx`�0(�]1ukz%|vC�u�����m,b����N�ٛ�p�Hq��1sVf�z�޺�3���=�3%U��H�8k�+/c`
1��@�?���9�hVn&�fx�ka�wab*9�t8h�ŕ��^7��uף���	7�o���g!G\��U���]sf�����P��S8z�D�^p��/^�u�Fwc������g0%J}���=�������ߩw0��ݤ��DiQ���vƇ��~Ε@E�0�3�ވ�*2`�gڬõ�º/� ��a ^,�Wx�;����Y>��ݐ���ɷ��n��?c���roh�+%���- �a���4ϧ�`3v~l=��4���0jNi��S��R�\�}˹��t\o�G�Qpjh�9�V~)�R��Mt&>a��<e{&g>{�*��I.�.�����Z���"/�;��7ckM9�u�%��y�q4��yPl*{^�[T�����b�<zo� j����")='e��nh����@�u���OO�-X �+{q����=u��l:z�;�d<gEf����䭨;*V�ң�L�p�T�"�,�ΚTTe�o6L|R�r�H|*I��l��V��3��I�5�9Y]��rQ;�I�8���QPy��Q���K�N��b�Ao=��WL��iWT�f�\��u�L:�$6���C=3%%S{�����!������W�v�Ꮐ������%]�Y�����s��\Jʐ�җVB��3C��u�u����v���E�Y��#[��(�;rRw!�V�1���P��+t��wT�H�af���1S�!��Z�n��ރ1��M[��&���U�R�V�8gA�1ǟn̠FmsxI��<��qs���K��z�9ٳT�|WZ��J��%�������q�����4�y����x4Q�}��u�r��ъ�3��Z�˙�qV%^MPX��\*�&b]N_u���h*7�oT��Q��@F���=����յ�7w�[R^�����ւ. ��6��N<��G���hs��^���v&t���G%M]C:�<����jl] If�<��z0+�;�Իn�F��gkR��PV&�Q&]��HwQ�PQ��[R�����Jo9�9���u�.^9��DMP�"k]<��vS��������էz3J�L���s�l�u�<�	�YT��zܜ�}�����;F7"��NP��D��>��R1b��==�4��F���x�r�m�U���$����2�\�@`��B�wG1�;�;�η��S��O��dT�J�)�s.v�sz�t)��ޮy�2`JI�Vl�y���6ӆ���Sp��g�@s��h�9��*]�[-Ȑs�q֭Qּ�A�}Ӟ��Tw9�kEB(�[�����#��n*�GfLGT�g�h{�Z���[ Q��u����Lc���^���	+�㭋s]s/w���>�r�݁�Z�O���-#5��O*-�1e�t}P`k��l�颐M��YՂ���'X�`�1�b-��ɔ2�f	��u��}Yf�͸Tڗ7Y�&�]oWe&i�(']��WZ�ܬ���&D��<����*1h|���wYWQ��l�ꕢV���P�@	�]z��˦�n�r��S�_��Jܝ\z�$:���Fo3�}r���t�I{ǲqA�7�uJ�Ooq�L�[l�e�<o9�2�\��;�n�-qW��t����ѹ;4;7:���$"�)e��]	��Ha!�;7����E$�����x�a�e��?��#��1D�5`Y䕄�z�W꒱���f9s��={{{{{}~?^3���6*���Κ���K��@�@�aJ퍭X��["d@�M,%��I-}x<{{|q���������G�里TFD�����8��"gՒ��+V\�WAq�!	@���ڎ{�8e��g�������;ϱ�>��y��FOD%X� ~nJI�G
 H��I��gV�2��#k)`,s�1�.ns=|{{{{}~>�gG�C�k�z�D@�ۄ�O8�0H��q����l��iH	��3kI�x�O���Ƿ�������>�����|(0HYm��u}z�7V0�ZJ@�KhH1A�zm���
8��Ȩ�������P��=��AfzL���ౝ�Jᬈ	S�g���	�	YbH�ph`�)�9msK
�QF���nKL�^�rXbA�"�0q@@A$����U 5k7Z�F�HHHM7b�E�n&6�%�BRS�Bh��Lدb� �4%" #�yo�x�9�<8s�ŗ!���Amb�z�d�]}��T�ĝ�7��٧�������H]f�6s�����> C� ��˲���1���0�WQ���۷��S��I�u�����H�	\{�#OQ���r�+�OS�̌ky�t�"!�\r�\��ڨ��_����<�we��`c�6�u�3\��'b��v��:v��A��+ٲ�:��qX�������	n�c�C�Tf�x�k4Jdj�U<2�<cO�߼m��_I�@oa�}4*{��3�����׎ؒB�b�t@���oAڲ=����&3j&s���1�ZM�%���ȩ2��nkۏ6��o;�=���h���֋�+9cY�_z;��]�.|�3�RP��Td`�l�a��oSۚ��WR��8�j��[�34Sn�r��O��'ψ7`ev�Q�����ǐE�
�Gڨ:�_@z*|�7��vO��/G�Y�gޡ�fb3���L�ʄ�H.�[��w��pg{mM�x�O�涶�kҌ)̒��V���yl|F�.n׹�2�54�q�g&e.�K�9Vps�k9T�b颭��p\��/����KDU�H��&Z��X{7�'�$�!�=�{��>������k昛Q��=���غ�"�����5<f[�8�Y��ӗ��Q��&̱�l��C
4)�W�h������J��oU���W�=��E�	��mh�(_q�R;��9�#sO�����2/�C�A�R��y^��z�-��\�q`��1�y�9��/'MZc}1~7<��ئth�������
��l��e��|A�����ѥQX�b��ky�;;3�;�>�ޚz�W��������Z�V#.mi�l�C1��櫐g�}{�⫥���`�z�8#-�.���E�.U�oM���6�M,�2U4�Fr�7��ەp����7Y�|�^3�Or��o
p�fi�ff/��n*��.���dA2.5-$���f�ń��0	*�N���O��:�!��<3�t�k��Tk�IE�4郅�ݗ6J��<�g���%F��j�{[�1u���n�L�N��#��% �Ub��8Dja�mtʀa�r�A��o�KΛ����"Sꓨ����ԕ���O3H�X���ʻ�rw�O9�*%�]\ ;�@0���k,і�Z�-��۱����@�DQ'�FS�Uu��O�H�I���&vh��_�;{+�}=��B��y)=~P�g}�UY
l`p6���޷���XD#ގ��������g����9S���wrBp�n_{.�S���c�t��:*Ty��5�:�,�'��f�զ��b�TP坛=�M���K�D���c��E_G�e��������5��vX��U�g���M@m�]�ð��L�p1�`��I�%M������moY�k+�C�q�Mϝm�G&~�U���Nl�;��V����g�3�)�{��Z�`%M��0�{&������]�D����[�[�^��U>2;�g5c�O���wy�$�b7�|*�߸�T�*�Ԛd"�FM}�_G�Ϩۚ�ߢo#�iO�I6�QM�9����y�B��:n���X��k�:�a�9�Qe��{ϼ���d�� ��9-.�;3�Pt*��jb^�K��r���z����^�{�;�1��Mֈ�	�bQ�ڈD!<=�);�{�y�k|��۞|fq��,j�;1f_
;�ʕ��������㮬R	�	DC;3,l�ԡ�k=���{ي�.��d�����V���k�@���6��"7�y0��x��bd�W�,���y<���mOk���u�;�auFZ���=<;�U��ɞή���͵4���`�s �C�_��VVc>����Iޣ�w��gǏHs��^-l�B}0������d2bY�e	�2y��35*�~�Ʀ�yu��Z-7"�*^�M9��\Nw�v}^�lq�2����dgGW���߳)�4��;��b���gJ�fK��-���Ӻ�����g2ŵE��}�Q��α*�Y-���>.ٲH��q('�LQ�å�-��@F��8-�i`3k��N!/ꣻ�j��z�����^W:\��V?�� ���_�q�+c�!��ˇf��˻�EO�5@����;<�Rk%���ۆc�62��5���sf�j�?z�5um�c��[}y���N��7[�e�\@�'���$I�	7��[�soړ�M&����&�3��<�O�--�.�4�����\�;,�����߄x�0D<��'!,4�Upj��C	N�h�@*���@Q�A�L����iȁd(� [�9�o��	����=f�¾􈚩YԳ���!���z��wp�iW/���Ӿ�d�����A��1�Y�MA���J���%��g*�O~����R��W��{�x��UC�1��Ƕ��iB�w�{�di`�W��x;�f��f�)u�Wv6�sw�ӶdR09�T�E��e*��+���Pz���u����h�w�U�̗�Ԏ�'�m"�zl�wF��jQ�>��<ߴ�nn ?e�K��y>0��;Us$�'9��}FD�8�.���>��oi���vn{Wr|��{�
�m�-���
G$?g�F�*𰍗t���:�;�wn�\�Сb���%'��'|�Q�%1�쬟gz]�����0�Y�Kш�E�ġi��Xհa�<n�B�>D��_v�ԅ���^�i�$J�,�,:��x�1�@���5����3f�	����9�G����iw��D�C�rw�-��{>9�<Xj��ov���� ��$A��~�y-<���L����RNǎ5f����~�~�a�e�ZјD�8-m0�=�yݾ���Ko�W}��vϷ�4Vd�F8�O�:o�u:�%h��df6���H���1���Xom]&eϗ�nF�S�;��W8����w>�Ϡ:a�B�ʯ\��w��1�1@����VLvEa�/>��i��O�������'��ն'�z��5��^����<:_�c�F�w�43�����bh�Z$n�{<knx�a�<9�pqG�w�F{��f���sbR���
L/���S�VT徛���b��J�/\Z��NEN+w�-���]������e�,nCU?Ϟ��F�Rp�sfi�^.8}��%Z��u^Y��#�FA8F���CBn�4�e���dǱ�թ]�wp?��~8
)K������S�.X��/Z��*�ae��ޏ:s�RlS�՝e��%ZYmF��)GG���0Y�X��t��g\����$���<2`
��񁹯�ɂ��:�s�/��%�y��A��ת	�މ���ɛ����`ٶ�@v����&�vl��(��]	[u�Մ+V�.2�Y��3�c	�2^��3�l����b.!��B\������������߾�&����SK�����!M�� �lLn�v����)Mk؛ܕ��U����dduy��>�=��O#q�m�[U�^.�i
���JL�H�ݞK8
!��Ϛ�e�	���登	[a�٧a�&:�-SM($�����/Z�����9XU�����Li3^�]x�6�H�:��V[�=�=<��^[�|��r}Z3�N;i�����v�c��GG�,����#�a%�]�S$䖧���I��^=����ܲ6�ܨ����^�]r<g���oxӿU<��L�ߎ�Fy��5�m��fZ�}�S���&�#S��s� ��,Ę�">罹�����u�UY�-3~����]�"��vԇ�k��ۇ�e�����:,S͙�=�C���8��덍h�!�\s�&�BvJv�7@�xݪ�ֵyeM���Q�%���7���9]}��� �����X�,c3x^^vz�0��S�;21&*��g�,)Ϯ�q]w����8���oA��:V�[9J�Jmd�Փk�,[�(۾��9�˧n���@6�ϿW�Q��x)�U����`�g�����?�0j��PPM2��a���NTJ�<n��p��Q�0�S�'CG��T	�8���\�����r�X�&)���͝~yi�*o�/�*��nV�wu���Pc����kX���:0FJĻ&|r��h톪����l$pS8�N�vk�E��Q6�YY�ݮ�*�vz�8�cu���Χ5���4��V��3B�C*������ݷ\�u*�>�e��V�͎T�ӑV�L]�C�ܬϯGX��R�E�D��(��{�����?�^��fz���V��5�yQљ�s������"!Q�9ޟ4�����M�Z�k��P��vN�c;5���ulV7N��q���Fm�����*��@�d�M���Swq��
��P�\Ȝ�HV&��4\33nv�_�58(��=��bp��;���l��{�)�m/�Җ;�)v���u �9�r�sW0ma
�����7��WV�́�3�]Jmf8Hk�X������w����N<�����}]+�b����0���j�N�W���;�D���<�E׷��+wvt���`"A��欽��U��iQԲ�y��ly��^��f�
p�0.�0{ß�Mt��Ul`þ=�{�d�߈3�A4d����ߧ;v�p�E7�Μ���l5v{[k��6��;s�;���
��N����}���=�wP�WJ��S>2x��w����0a�\���6��Q�dm�']��s�T�ߣ�m.X�A����￾�w�`U|�6��b�&Y�� <��%���}}�2ʋ�c� `Ӆ��^C�<Q�<��%t�9�j��vfG�ʙ��T�U��y��:�H���}<r�J��gP��o:T�6&���/�=t�<�.��"�����[��/{~�X�#�w'�}�>���ݏT2 ��1��ʮ)�S:Sl�Yg	�a}-��<Q��)O�]�.�L�8���Ь͉�٣v�������N�q5g�J����a�qت�OU� 2�DOv������8>[�:��1A��30���B�x�)h� PS #�Y��9�9�7b��R�sUNǯ���Vc����>������N��7/�t�.+�әt�#�(��#;{m���	��d���{{5���0SM��oǝ�/.�[xe�ֶ���{R���E�>�����.���˒�+�͡���>RA!���Ra'q�mG�T{���������ls�-��Uʖ��7m�ڶ���BuF��y����岻C���l�al!�;����	WFl1U[+{ȣ�r���]�noa��Ѭ�eOd�����J{<wf����g�����Cٌ���YB�W�-K=Iy�b��a�u�0.��ǋ)dC���'<���_}Ә3�ؽ����I2 �U:؞��{Q~!�>�Cu���z���>��FBY!n}�b�n�;���;��h#gg׮~��8o��k��+�K@�wo`%�:��ǳ��5L@�q���M���n{�|=[2vM]WA���}���<|��������?�����s���DAW����������W��C���ttH"	��:�<�g|2�XB�%F%! F%F$V!%�^pQ�+B,!��*��
�@���� !�BDD BD�X��!�@��!�@*!"�u׃�v	$J�� �% �@`BQQ�E$T�`BP�!�TH�Q B@�B$A�D BA�B �P � BE@�U$�P BQ@�	A$D�P BErG�!(�@�
��!(0!*�! �!�!*0!*0! ���t(����������������"��"�����*s�!�F F !$!�BaQ�E뮀C�F%F F% F F %F  G�A0!0!
�!0! �! �!"�!
0!�!���ϐp��_��ET�U*����?����ߐ��������W�~P���/��{�����������Ͽc��DAW��������U_��Ȉ��@������ d�O�/�'���"��*���C�~���ޒz����?����}���?��\�^��0+@(!B"�"�H�B�*ңH�J-"�@�@�(�-"�@��@��̂ҌH,�1"��(ċ@-�$,��-*0H�ī2 (� R,�����($�,��H��̂� �� �"�*�!�,0,@�0�#��1�B�
��*�ȴ+ ����(H� �,�J3̋
H�@��,+$+@�ʒ�2�,2, H��!"��
Ȱ�1�0(�,���2�+H�"�(�J�,�$�2�*�B2J2@	�̫*Ȱ@���	�#@��+$�0�����@��$0,�"��,�,@J2�-"ģ@�0�(�-���*20��@���ģ"� �@),� !, ��R�@
C�2*% *P1"��%NJ�J(J�	H����p����O�E((@hTT�P�@�����~�����C�t�|�<��"
���~�����X'�v��?����������U��P�t���~�� �
��U��?V��DA��?p���
���������΃����s�|O��y>��@vh����!����?�U�C�P��h?�~����~���?'�~����<Ds���J" ����?n!�R~�������|O��I��A���ߡ'���" ��e5'χ�N ���A�_���M�@��l��j�//���w����8��O��PVI��Fyl$�mV` ����������oEQR�R�R�D )��TH�JJ���QDEE%�T�
��T(���@T��RI�U"TH!UB��R(T�A ���IPBJ(�T�!D�RTTT���%Q%E$JAU"�D�Q
Z�H%IIIT�)R�"T��� *���)
��
"P�J)%U
R�*JR��������B�P�� ��Q   ���m�l�����Mmj��ڬi������ե��U*4T�m+f��f��Ջ1�Q��4�	j�UKZ�[m4[F�m[L�4AD�B���RUR�-�  CB��fB�
t���T�T�$D�S�t*wYj�[!e�֐4��+mmcUcj��,�V�3R�ڴ�"R٦�R�h�kY�ب�j���4U ���IT�JUU*�   ݍ���M-�Yk-a��a����F�hʭj�S)Sjb�T�$el��*��B��a�6��6e�Q�T)	T*�
JER7   ;��m�����B�X�X��֕
�[Y��K(��Z�5+ZYkA��6Vֶ,2��UV�@�������T��DQ@�U�  .�44,�j���lֈ6���	M��Lڣj5JVm���kd�[V�	�T�ȃ�j�Pi �V��*�U*DD%$��  r������j�����"E��4�� j��(�-�P$�
4� ��`i 
��H��DI8  p@��U�  MC@�P�k  �)@ f�� (*�V � �� � P LI%J�!!
 ���   ��  3�l a` ѪM (R���( 5�MP �0 42� ����E@L�  ��I()QUD%n   w    	��҅
1� U6�Қ �b`ZT�  ���L�  �m��@�(�UEQ*�PU�R!p   ˀ�  )�р  ��eh ZV j�*� R�L  �`
P�cU�h
Q�0  E? �%JR �Oh�JJR �ɉ�LL��JR�  S�L%4~��  L���UQ���jgU�h�˵��>�3����7Y�0\"�,ֈ4{���X�?�諭����}�>_��co�60�����1���`���`�� l`������T 솇a) �� ;X�3*�H�KM���2»�ŀ)�iюⲒגѪ����^�*������.��`X��sI�.s��,6���fA�2��+�¾���ń���]�̌'����f�O6�r޼hLwzff���Ӱ�4f*�R
=IJ�r2CЩ���n��Q���%�FL!W�osZd�1̬�ؤm��ws-7W X@��x��f�3�E����)l e�c�M;Xuh��D�v31਎
�y	�C!ɸb6����V�JAڡ�dm�Z��ج���v"%��mE�U�V�h�]��Z�+���!Z�R�m�Q"�iz�I5��S��下ۣ��7kOۖ���6��j�s�� g(�f5�K�@����t�{���Nd�>D��%�A�Bq��T���Ђ@�{�Q�j��۵��A�MX7O ����L��6C5wZ����"k�	͓�&)yW�i�h�YN�5{Pe��l͹Le�(2���(6��/QZ��'I؛���6��m�b��Y��:���m�"�U�j�Vz\�r���T/w%�`��٠���,�-k[������vV�����WӬ���ǐa������V���Q�mS��)iԡMn N��j`j�- �MYO&c�p��$ {w��PA�5�X�F�n*�[8$7qiC,b��$���x!���$��۷�^�ͻn�K)"!*Νٲ�
X��H�$n�3ק8j|���fى"�kE����N]3� �����MrL&`(��we���i��55���ͳ�V���ƚ�x�ws�Uhe�ש�̈to5m��$lm)�.y�"ΰ�$�i�ux+
���b��	�yL\�Gl؈��5ub��n���cA�f�:mVn)�c����SW���mEr���b�R�LE�*��:��/FF�5Ռ5�b��K4�p\�����d�����2�̀;)M�u �-��f�O-��S�O]��"m�t[̩� �`1oJ��ͭ�3)XKT�l![�wx��
�R��y��35+CE�Ii�Al��J�ܼ.ACr�Ukr�mI�[��$4���ʻ"�4��M6s1tr%C)C����l�B�mVȕ=YcI8e�3i�k���6*�Xp���	m-�͒1�YV%+�E�[3r�cw695Y��B1������`��[(��8j	WaŔ�9Tׂ]��-�%�X-���Yb�̀�w���hn���� y���T5N;�M�x)Ї-�QP�3* .#���E�gF�א�l�Of���tA#V�m��$���X	��`j�(��ʑ�G��X�-nb��Zw�Ɠi�6u�DYB�l�T��T�ʏ.�J�b�媻d3��T�%�[MR�YmLH �[$٘�7e�	`f��OU���T��70n��TI�{���Y-ڶHu�F$��Ƒɴ�XؕK��m�n����wATͼ�4�襉ޙ$d���I��[c�������ZwB��ʼ��:�X���y�p�L"G�Dz��DI��O?�n���[Q�Y�8����fP���a��0�R���{��fU�kt�n�r9r����	�-�x�09Y+�ӽ�>TC��0����r�J	[��f-'Z�azjd씝��3-ޫ��J��R�&5�a4�[�ú����	eE�$�l����̏&�E<@���M(]%WhLdm�2w.������Ոp����Ĵ��u���Z�Z���[vƫ�w{O)�E@��؈ln21�{��j[���~�j��4E�t+NA���Ĳ䦷5�]�hMkJڍ��ܸ�L��sr�9T!�b�}�Tm�ۈ8n'�6֡�̌�ux�Y�\n�V�K`�x\�R��LVU�t;� Y�H�^Btjb�&,�*�+k�/q`�o�h1���ٻ/b�
6��΂�4M�n#�l��֪� �	MMcs-�*�q���--8 �CJG%�6bfH�;�q<x�KnkjQ�z%� �1\���+�-�5ux���L�4��Vn��F�lhO/E���W��e��C
�ͽy��d�u+IN�A늶��K^����^�t�CN�"1C"ve�(�����>.�r�D,�x�����tX�su�s.��ܬ���K���|�t��h�U�V5�E�;E�ͨpY�fJ�݁W�Y8)��{j�ێ�Jb;P�B7�kwJ�V�^��C�{� �����՘kH;A�-6Kt` �9�v#2���ZmS:0���臮P��O�P��e�G0)����F�T�Z!� ��L�{6���:3H�Ul4�Y�k�-`�Ŕ��H��:��[�Px�jn��0J9�΀Z�1���S:��n6�m*2�S�j^QǌU����N�úU�cin�Y�d���V�J�hІ*�t�h2�z�ktP5��,��i�V������19f�iQ�-ل�R��Z����{[| �Y�V�[�j�a�#���[q�1�i�RŷO6K�lLG,���6���F�M3aNޔ⩧[���k��X/`�	$ʼ��W[x���j�sX9��I�����`,FeL�0[R:2��B�E�����[��M���ƶ�4wv0�r���o6�pK����J�3��4�
U�f䎭Vn��W�:o�&��j�,*j�+B��9"���N�i!/E�GY&���z�:��F3��S�]�Ɲ�:v���ۥkEGj�F�S8�8��x1*�����Y�������|P�s%��Q�yl-�+Z��%����.6�w"���K��R�ۭP^+74[��AVȱ�F����tS�V�R&Zu{$�F�nA,۵�HRy!jCn�;͂}�O��ͨ�!I62A�Ԑ �XX�td��2eŴ���(�t*콡�F�������e#�N�X34��6���n�u4�Q����y8)����4���z���3�]Dp��a��R �YN��R�I�<b�r1]7[�ȸ�*�Z7a��B��3X��bwB�L���St��F=mH���/6VDثC��ژ
��T�C7r���%!.�kv�$��Ӣ�;"���[���ŪC��A�
ٙ6�P(Ջ�:�O�]X9!�kl�t�fd]��I�� 7x�)͠j3a���e��bǋQU�b��:p�\�wz(V�ŷ���/^l��چfKPT��`V����=�O[[d�J�kJ)X��֦'�Y"��*�
�Ӂ�J�[��ϝ%�m�m����Q���{���$����$�Ԛڼ�l��RZ��'2��2�@
rc���"�n�<Y�d�u��&Z&�
�@�U5x��C�OVS֓㬃��` ��ذ];u6d�-�6�T�[��,W�T]	/1Qr��[�5ۂ�t�p��#u�#�y{'��r�ҫw��t�j(�i�nM�R�EC�0��b�2g)������A�	3"˛Q���Q�ۚ)�����ݦ!1k.�*�uw>1V�=ͩ�M.��V
���mJ6K��v�k\����Af,�6���J)0�H�Y��K����#fhF�8�T�3{�CH1�ڂU�lY҈(����j�94�s*�ܹz��R�c�̸��.��(% -K��]���J����,�(�ޅ��Nj[P�w�u�eS�y�U��v��j��L�P­Z�WH0�` \�P�m��@�Zb���tp�� f�� ����bC.�
rJ�u*�wYe��m���-'�Q��u��T�O��\&�/7�A�-�)������:i�����{�5��*��j〵����6����Zda5���&�R,ɩj�(n�5K�ɫ�{BP�p��[�*wbV*�YL,�SˤQ�'�Kp�l�������v������dd��tӴ 1��r�H�G2��˭a$! ѵ�k�@J�dGB][�(�ʍ�;�B_�W��Me�k˷�՚sT0�gn[�p�P��ކ�YS�n��0Zr���(4�B��f�TpF��X�W����h*�٠�݄�f�H�3>8%��G-���Mb�oL���P�C�J��wn���g��)hC/�F�4�7\.���ԕFxZ����[�6�*��-�4F��em:��>Y�(�v��J9��L���)9��M���A�Q��4�2T��)\�Y.��L����xiQ-��0-T����qR�������R�d�1`�d���pF���Fn�%ӡXM���`6A6;#�t�
wJ����t�Te鳻j8����ݷ#5�(���և	�4�n:�U��9��EB��j������(��Cm@R�T�8��8ɰ��R�t��WW��o�&��K�Fwݐ��c ٌh�l��wYQ�M-�v�r!�z�]�5c�������9M����e�r�Q�k��ڦ��#:�J�Zа�p��lv �Lej�븍uj�m���j��lj�5{�$��,�f�Ǯ�Q#�[���˓���҆KO5�V���4mC�ضR%b���%t8�E��k�WK#�X��ƤUXY2�$��Ӊ�Ub���rU��*�7H���P��G�Oh����Q�0f� q��u��D'&�9�bXze�L�`wJ��/�����#l\L!��P�� <��׸�CL,��Br�S%�D��n�p��*LG�GP����	�Rm��[x�$Z&A��]�:�kM%O�V1�%��I	���%5F�ʒ��@��x�{Zhg��c�zo(�mI�PR9L4f���i�a#!_f����ĥ����F�?
RT�"����/s�u6�ʊ�t�nMQ,KĲ���LbE0k.�Շ��J��`mO`zѼ�4-�v
��+�Iҩj�Յ��	@ ��%��Yo6��F��&��uvID��fL|K�iǀ9�oo�-�����B�����Tn�0�n�$@ko.a&�d�*M�I�#�R��,�~��� ���N5��D���Y-d���E �5+s�mo	��S�L�<Р��"H�ߵ��V'�R�95F��e=��JF���%nlpU���yc(E���B��ώV���;���ň���l��@�M��gwH��!���XƩ��`��*lT	��r艈M�_]1Qع�S�cU;g4%�e3�d��*G6��L��
�V��k#^���q��6���ú�S)n�iy-�jmoȑX*G�K"Ԫ�me������%\V�T�╧5d��ZCv�_�[��цR�SZo~��9e��:�Q�y�")FPX��U�Vd`"¯Y&�r��T�Z�e�ܩ�3�� �̠YP��jl0�U�ł��:���^e&[l�٫V���ܒ�Flӷ�mJl�T�p"o1P�����kCh���dV:�IN (��{�m�v.��ڹ��^<xR�z��/-Rˣ"�["Z�30Ne����]�)��QF-��!D&־�@��Ru�
V6(��*�&���N�ԼFЈ�C/>�nc�rM�NTA�7Q� \qf�;.����k4&1�m�_K˗j�D^�T��&:NV��-��E&Y�.^���z.ؤ̔�Z��1M�Рv����[�;�q���2�E�ǁք���x����2�m�R�Ѻ3%�& aڸv�De��Ū�&"�1��[-�v]�ѕي#�2�b��ˈ����4 ���fQ����!�v��Z�������%�^���4٠�*�r�e��-+��\���{6Fw"��6Z�K�N8#�Ը�h;��d�ZFZ�tۉ]�C3�«�r6�fUn�G$�WV�5�e�@�� ;JSƎ^l(i [�4jx�Z��:�'z#���ܘr�Ŷ�b�̻��+i�d%p�^ѽ�4��u5��D��+�Khl5���Z˕*�
��xx���	M��JM����Y�VX��XbnE2���Ɂ��0Ř/6(cʲ�MkV����,�F�]f���w�F��z���`�$�j��*�:U���n�Sߘ�/A���3n��4�e�XL;Y,�ܫ�z����52�ɴ5D�Z�Gj
�u{Z)lW�]1Km��]���n� mX�6퀁i���m�7��Yn�Oڀ��-�hT��q@�e������H4�QYQ��̬���Z�����'[��ffi�'�8��s6V 7H�!4��"��ܸnd��*�WwH޵J�N&��,U�@G�*q�O.�W�Rf�Cf�[�o*�醂�֌��n��ʻ��˖w[�ɩ���٘��Q�b$�0VU���
�i���W��.�̠�3l��bpΓ�k]Ek��Vʎ�i�<�"V�断Vި�f��X�����R�v�ɏB�n�q��W������[��iRy)�29R��Gͭ&���5^��:��C ���Mt7@�7�F争��ta[VX�2���$E����
�0\ݩ7r3+r��J�]*R���q'c��aRV�hEޝH<ݖ���P�I܎��Pk���#�QP������M�љz�L�YV���tU����١�SLۘ��q�O�Y[E%���3I%#�ۊ\��Ug��pc�hr�,���[Nay-
��X�A6�墴��Ln̩���l���/K��nۋ
u XNՐ���VfK����TNG&(C��q^,�޽0�ұ9��kzRr#z���#q<r�ò�R%婵D��&�/lm�l�"�`�Y,�(���#��`�p*G`{�(��Y8�(�(IqI�1B��X*j�tR2 �F�)�љM�\B���/U��[S7�
'W1e�p�Q]�59F�ޒ����kKuSK31�%	�L���2�U*�!�����>���]:�(�P�I��+g5b�^Y��c�+e�s���D]ܧ1R�6�3z����s�.o[`h���	�%��yյ�x��&��[�o�5ζ�;WN�ͮ�m;�k�!�@i���К5�-��l&R��7��k(������Ved�t3
���'r�� Cǹ�]JLN&��tH S'���j{�1�V3:�������k��zֆP�#C��|:���:m�{Y�Jg�5uՊ�H��T� ��G֋=��˾��fjP��&-X2e.V���v�|��M��.C����jqA^���h��XHɗZ���b��t����"&{/�w	�۫�R��3���b��� �2a��T)�A�7���������wyۜDZ��d�\��×�[(E�m�[�q�s0I�u��n�
H\�i��)���&�/i],+�+�p�j���[��4Ƚ� 갎�g����n-��|�p�d��S��,ں,n����Փ+�KH��2����YR��1a�ֺ��{�<�T��$��-)�'}��Sv�٣E7Ue���3P���t %j����d�45�|�����o[��49�F���4��op�G���N;�|��,f�G�y�v�8�7H;���xE7Xv�4���7Y ���u����[�RN�I*��L�rD��ܵ/�s[TAE���w|h阳(���
��5K��VΉ  �f1��łV����"��Z�(��v�,.[�����0�L���t�-.���Nf�6`���>v�U����-2���)���꼺	�^�ee5�8��m��e�]��'���8p�BJ��myI��]NSwdy������*㪵b9N�{�%�+\�DU:S�w-�su���hܳ���>�ҳ�1���V�9qҳ2Q�ľç�R��/���W4]���9:���ݱ��,��
L�4r��3y������e�����%t�W}��8�ii�ډY5ۃdg'=�����MC2��X@�*c����J=:������|
��u �R�(�B<���gc?(vU�Ixr*`�?�R��&�7Y*R��o/_!Q�ZM#�F�c�R�>;���t
���f�v*:��K:�+��]�T���lV��b��]}�g(3`�N���G�ݼP��h�2��>��q�J�n������0]#R��y�'�v�v�錡=�l��ȁ�|���`Y�A��rXZ`P��ٷ�}��Z..��f��"V��1W.R�G�������9 �8���Z��f��������^�,� �\X�q��P���Ȏ�m�,36���V�=9V��m<�#�n�Y���mD�U�`�ojBBSD�:�ӛ�޻�p8[{� Z���p�]lR��{̼6��V��|���﯏�[�����w]E�p=���eg003d�G�7%��=v��uf�r�z�1g7-����w3#�t���+:K�#�����&�����yt��ژ�;,v}�t ���^��i��#�ٗ�E�y�m��.�ӕk�[�3]��8�msS6�`�t���c�:�����Vw�/']���u�0�yИ������j>s:U�},_zv� �i��l3�;�s����{��X�.�U��_���a�oR���5�IV4䶺<{ƭ�r��"*Ԃ�[G��'%�|p����E�l���[�oEtMҠ���7۴��*�I�r�v�6������ ���o�$�B��_,;)ޅ[3����)^��c8�Ѽ�#z�Z�*��7kFR���Եb#vFq�:}��X���n�u�u��_(K�/j�[f�)nU��i�ќ�)9���Di�ݸ�A�,mʝ��ۧ��0!�5��'�;I�����'L�⺳�mS���_ �
���{�\�O���`�{�C�`w�vS�QU���"a�8��������L�9�c��fPҟv�X�3�U��7,ǳ�P��>���c�O�߫$�~��h�3�%_mrاe<�+�렯�7��}��׹��Gs�dx3t�r-:�3kˣ�� U�As�9*Gp�cU�oox��є]\:b�+)�-p��4�'An+�%n���s�u����U�\���w�}G��7���N��]Y�����^��}M�6��]<c���]�ޝ��C/��9I>�4�2Yڬt���<�Ar
n[<���y^�Lg������u�X�[���J���2trr��N��˔ݤ�/>�D�̊�=�6k
�(Ism�v��=��΍���s��Õ[��ޥ2��^���u�5V�ժ�R��~ƃѪ����ض�pÕυ�Irm�[��W3MY8�u1���A|\�u�餹�����s�ٗ��k��*R�3y��rk�}u�eZ��HA1���+��-�ksh=%5�nU�B.��n)`U�Xu�Q��R7��+��`�\2��뛄�S��������;��v���F����Jwy]��u��C{e�+�	�:]79�g*�ct*��'NG��X��fl�4�>T�1�M0D�q�Naū����#�5�)�'\S��ĭX�=q���2g!7��JF��0+<c�.��Q��mc��r��p(����.yV�☰5���	�p҃P�|�^��Ճ�\�#ì��c*�i������V^%����ٻ=��X��N�������>����k��E��L:��.��hv���\�v�o��]��j�FWJy���v�p#�q�Se�\µ⥊u�q�3ns��5��-��$n�Y�Yv�A�pRu8u�vɡ�s,r���E�N���g��l�p"��ǘ�%qi`�{P��	F�Ϝ)u�W��p�
���M�ch���n*yc^a�vR+�7�4W� �%��-�{Ư;wQ{����ruKr_}pua�)�� �	�Vwřw�D�<�/�(S��Q�Zp�\�d��>�7y6����N�����A�������@�qw'xi�̔6K3�B�&�yC˕�������؄�77-�쾙�4�
Z>jgsz�%�qW]�7{�tXNq�2k�3<^VK���=����g>��'`1+��z�7����M��ۇe���͕-�����K�r��&'�}R�p0�'-Z�]������VmDfL��5p+୕v,-���eV�o��,���@���-Z�S�ץ�~��wSF���{�sV���"��ͬ��7��S������V;�98I&�&%�K�.�h}y�2��ъ�YpӣМ7�;Qm`��}R˕�>cZm�5�0���Rֳ���ດf�����u�����{|ne@��r��&.��PY�G:�-:�w:�v]��r$0w�8m�Wu�V�,��͎T4��f}��6�����r_,��F�wwoib����C�"�D���-���r�΄�ɩWf��GBGfdz�DX�*�Q�
N��d�]_ru�� ���-��e�@Ί�'�u��6�<֩�%��:4�f:�mL�	�ܶ�E�<c	���Z�ޜj�%�4���;R��81V�����Y�rīЫ�>]�WyI�oV2�%���X�WMZ��}��D��>�4��M�nq[��^J��{rWd[]*L�ͫc)Fͨf�<��`j٪���J�Y��6{�7�Ǝ����%�o�E"d�f��ˬ�+
�͠��]�B�D���c!ޢ�A�ݸ�+P���%
UƯT�s�O*�
��CO�%��\&-�1y� �f��{���M����)�i[�3l�9ۓ
��k��p������V��袾��ŗ������*v(�\�ٲ�W7)a<��t�U�H�>=O`}m�od'C�Nl*�а ̸�݇�<~�~��w+[F���9�ЋU�(�"�i��-�Qcju:}q[�ٖ��>��8�`IKNH����#��^=�o�k�p�u�p�=A� *�R�U}��έ�Ad�F���wf=�J^]���S�3N�����ݛ}{Rl����Bsv���hӱ��&߲�jDZ���߫�ʖq�X��I�IoJw( ��/j>�"�(��4�΋�o���խ���/�A��gg���e�U�٨��q���ݺ9Me��S,xG�-o���i%m���9A�|k�wpW����=�_ƒ�7�E�	e_9ڶ��ތz�#�c]�ƀ6��Νu$�i�=m=��
u-Ox棓FG�\�E��T-.s��F�h�}�j;�M���͘��n��ր����Eh�փ�hZ��k�/:�W�i��w�1f 1	�O!A�z!V���7�-˓�%C3*�$�)P�1C���OGA�'|�:@ֹn�WUe�b\���f�6Gi����6�z��6��t\�m�oG
g^
�rn:���u���cN'Ӹ��u7��Z��MN��T}�+x���n�3���_W�g�e�"�[��[!�7��i��޶���+S�mIR��
��kj	}��)�9Z�{6gKJE��{x�����m7v��2�s��D��\ڍ��I4��MU�q=�]�*S华�����Zn�37����3�^v5��ң�!�Bq����p��;`b1K��m�5�Ft�o3��$͐][�9��N������B�#��(S1Q�u�B�D�#q�Sf��g��B�|�t��4��Ug��#��.7]���'
_a�0ˬξ<�V�D�B�x�e�И��2V�;G}�M�}5��c�W�]��n)�˫��'w$�/�ʅ<�j�ѷ}ƅa�tqq{�l��݈e��*Lh�
�|�F�����N���+�i��B����Mi�%�	ko�=�wp_g*�**��!�Y�dC.^��#w��:����F�FX�pm��xe���x�3������d�אTvl
:V%j��w#�}|8�@��� ���6��:Ό*��4G�І�iH� �����M�ˮ�N��D%��od�(gp8�*E8�*����Z�^���m-2m���u��j.Č�E�w��	!=Qeɘ~&�	��u�'b�e�K�B(>�iDe��kk����W�bx�3O:,�=Va��uo�e����|N��Ts����#ɚMh��/v����Q��,}�hW��S�Ya$h1��_>pü���\#�)�[�2Q��ע�Cbk˚�Zc�K/�W�~[Y;�aG)ϣ1J�Z����$+�AJa����w0�X����#�����*�)�-)��T]h��n��$m��&�Dֻ�V���Md�q>��}xk�P�yLorg!�~C0ꈑ�k!�����td��F�<l_f��K�Spd�l��Qp�fƩ;1�i�M��R�ڳ�D�eK����ˡ%�Ţ��;���v�ݮ�0���48��w��:�����KS;6+\��z�M�����jśBؤ�]g�Z��b3��9�m�FI2���E1�Ӕ5�e��q�;Y��,�k��'N�SsS��1j��!��G4�}/wA�d	QNʘQ=.kA��}υ>�:��ޜ�vT('��7�w��ԇ��'k;;dV����i��0��g�)#��m�%�%��Q�6g#8s�m�,��Q��3�1�pr�4��U�b�O��v�+:eaIRemt{nZ�:��Ǌ�)*Į��,�c]������U�U�vVC0r]���Sr����V�qDsgps3uw_U�z��)�X����pF��yOz=������`�υ�a��jA��N�׏V��V�023@�.��ۘ{�����R��\m���,5�i�ʗ�;�N���d�uٷp����w݋�d4�Q����Y�|:ÙN�,�4�C7iM8i=���Ƴ�g#�q�(s)G��l�}wv�f�K�ջ[u���
�R�άA
j��aJ3��9m`�C����|��N��꠳��O�����U�]���O�@�c�T�\8�Վ��Cw�<Z��[���:��b�"[W�nt�]�j�r�j�
U�-���z���`B= ��\�G)M�sA.��pw�O_\�%�D�»f�&�G��o7���׼)R�M=m��M�y���z�
��sQU*��
��t���/���.����tL������uv�p.�()�^7�z��`�����%2{
WG/��'�c�]5lS�������5�r��0�n��*�M�R�.�ۣ(CmE��wjwb�C�欦�����Sqpm�Lk��"�Ӈs���v����I�j��F��}�&�N�"�Kl�u�痩��z����VLʗ��jY�Pݕ�@�1P
l�z�>�*�����iJǴ����ʝ�Ve�$�k"���Hk��������ػ˷�"ⲳ��&�MƆfitٸ���\S{�@�Wf��wk{R��3x�N�JX�]s���v:��eg"7��M�F�*�}���UlA�����s�]r��W6��Ή�f!�m��ϑ[�g���v���4�
1�_X0e#�8WD��i6X# �a+���}��,s1}��v�U��R�� I�rJ�R���Yl�����e�;����2�8���s�8���)<���rm�W
;�uwX��.��{g�����>!�|�n�]Z4̫�t�=&��xc9���b��w�g_ �<��r���V�Kz���pe�h�-i��3A���,���Φ���j�2�]�vmwa�R��;MԧC�`�!'[�R��LjkE5|�97y�%��|γ],A����>��*�	�؆��Ĵ^f�[����J\�j؊�:������@v4Q��dqq�'$�Y�N����r�#�ԃ�s5���l���ġ��%�{!������ܞ��ז��9�t���82s�˹�'����o�<Z�͜5Źs7�>�N�=�N�)�8,u*�p��V��m���5}��7�<�Ʋ:�3���;����c�;�6�����1��uz�s���=���&Ɔ�l�61g�xP����ڸ;��WtSK�Jݮ��!v(�#{��*�T����s�]��KWb�(aR�3c$HK�;���W�2�Ɵus@�l�e�r���ަ�sS����m���hX��w��*m_t�΄��ʶͩ�%ag�xF�W����m���n:�ҽs싮�!��4���V����(MM�Rv���ucض�*=2YV��zu˦M��/as&F�cʏ��m�	�wT:��.o��LEtη+Mc�G���;Eڼ�r4i9��+4��
�d}�E�A�ޜ�u�Md}Auv�t�\����*PS9%؛�����u����Nͺ1e����<�����;m��g*�e�u�g ��]�9�s&��n��r�(���S�]N�ui��qVe����S���M(+[��|wy��틘��e���+*=�h]ƭ�����ѽ2����Yb�$���geَ���j�+�63R�Ni}ǃ���.	����B0z����w�[��[�m4���y���Q9������l�d�b��t�5�|q�ws{H]�6��5��(l"��W�#��4�V7M��ֹo	N�,�qa͈l��WM��k�6�:�]�Q�+���a�Y4<ie��D�jW�v��M�ջ�u/�L@��Wk����9C�7,']�pe.�t'̻T1кʵ����u6m^ZWX�t,Wv8�Kbښ,��Kqe��;aƃ��q�51�x�7DV�U�h=��,.ܜ}�ա%f���[�:�Iu^�����Ȯ��z�J�s�q�B�1�m�}dn %�vI�V@��\�y������m�u_�]	�U]�ڛ�Sc�}Z�vi�b ��ܔ��w�Q���"0�]����m��u�m�ʼ���.U�4�
k��feY%��*�X��\W��2�CIʺ�]��)�ۮ>w�k�9feܭt�
�h�Xp�'b�S��-�;�� v�=�2w��u���*G�:�'g����(>�6��(�)
�[{ג�wCfД�#C��P�I]h=9�ⶸ`�_�tr��Ǌ�|j*D�o4�{��ՑZ{�6��SDL8D&�_s���G��7R��q����i����`oE%b	�vƝ�n_*	M�笴$pA �CŃ13�����͢�J�]V���8ؙ��ȵܸ����6�qR���N�#���Ӻn�.Z�>�3�Q눥Ǹ�
�]رF嗔�z�1���������%��α[\́�0��IW@e5|�KA/:
�����ߛ}F�J=A:�T�&��@ŽD����4����9��i"vPr�m�YI���U�Q�2ͥ�Z�nc�u���a��^��E��]��o�r��BBR�⣸n�ߖ� ��*�2�5�u�Gb�'��*��$�����|���cW�X�?v�A_I���Χ ��
��ff�������6A�%:��k
YG�mgE�@�Zk`�%d�Uf����U�WU(|�-(xT��P5�)��t�>��I�VSYZ:�u��2������&�kd����a�J(a�6�����,��]V;������KLv��q�#�8ᛄLw���4�v��_e��K3�윖�`=HL!l�ɂ�]6�Y�n��+:؎�N�\�
��i�wn]����_h����\7��Ʈ˼�ա�B.�B���);!��4R�0�Z�M���nb��ŕ&���Q	���T(mp�&�JL�˭oAi��]�LbhW]�ӟS�u�.v���ή��}m˵t��b��7���_RH]O"Z*��Z�.m6��uy�����R��WAZ[j��_q��l:��&خ�$%�d[毫�(��|n�J�)�׬�-��s���C�a���A�6Ň/&��C��&�t��U&*
Z!+�lJ��^��B�ޢ��)P�{hf�f�p�R������!_l�Rd�ӻ���v7���.v4����9��BC&=o����y)�f�O)]G��a�;��;7��o���p���ʼ;��B���+ؠ���i��&�!�R�!�B�.�i�X����(��j��yқ]�[[S�[]�a��xe�Q�]����9:�j�X��ކv#}V� �g)%qӽPY"�en7n��Z�`c��	0�*Ba5�(��٭s��*<�o��x� �T������y�=���͉P'/~��[u.����,��7�uԊ�a�n���ܼ���1B��$���ǹ���V%��s�.��+�Nv҃].�L��L�kN���Y$�����r-�l�=�Kꗑ�ԏj=�5��4`���+�����$�J����p�x'`qF���\ۘ��3&=n����^�G��5�����y󃴷n����w�LkrK(���\����k�^ѿ�V��YS�+^[�QO�����ì!���(�'n#7�peUփ���x�Ґ��q�-���1k��w4��.�@vJ�� a�E��X��O,}��T,=����'e���;�o%A��'6j^�v��v�tH4�d�Q�X�e���N��:f;�v�Z�ܟ7c����b����X��V����Da�ˋ,L1�ڟ1�Rf�_�����Zp�v�^e-B�!%G�#����W�@��ujR�F(�0�GGL�8R���Z���L8-S!����ꒋ�IP�a	�e��u-��|�7.�M�,��3$�������k�f���OQ���x^8��+Ų�нT�)���%�d"�w����õ{S��Qu� #�X5��iL��·�Cn��mڟ-��s;sq*��ՋX}̮�V;k��e�h.������I3P�s��f�Ą�F���{�݆�rM�R����(@�����v��±w�0��R��9Hk��eʰU�*4�u�d:��q 2��F9��أ��sɠ�]�ݡ��z�j�kwB�R��5o*��u�1�cμk
���5f������ݱ��g4D;�A���3�A1Uyn�8��]vw��L��pf��갑�%�F���зr7.����5�NЋx���g] ͭ�Ӯ�r�vq֬��y@�ue��*z���LT�]��)�y��ln�$�#�(A�Q��ɭoZ��J��7�ҡ�V:I���f�z$��u�(ccA�9(*U��7pPR�I����Q��[���U��pvj�C�C/��&��%v���[��Y���\��܊�ue��:���+�5��-�S%�k���#�o��u'@���Ɛt�ɒ�voA�[����I�P��+\���ʳ�#�� ��<�$B�{[�-LM�el���0�$���}0U�e�6C�N�ѹ�i9+���뭼u�0��m�v�+r�.R͚x�F�5,�x�:�:ދ��I����x-���*f�!e�JW��7�W8jثM��3�^vW(&j���m�ʄ��(���7fv��N
�.K]��^-O9���q��e�I%W|qV��E�����{¥j4��qV������.�2S����쾀��#ױI+���7[�����5Ν��O���f�!*�#�09\�8:�;�8Q�&i�R��"�B�ݳt��{VCs#i�a������2qG�����6�ŀ���ǁ|)���]'gS�*=X�a(�`uD�-�`��%�K,���>���h��g��UЋ�X�����5�{��}w,�ݸfE��]<NI*Ë���e���̚��[��D���Q]NPjԎHw���{�_;/����t.
X�
k+j���̚��X��3��;s�h�z��gj���u��|�4��a#u ��r�t����Ҹ��;+��2�mպ2����/`@[4w��eZ��Պ�,��V��i����M��{�]^(/'`��'e@󶶳 �6�!�0WC������d�S>�K�[�r�g@Eu���c�y]��!^�����:�)��hN�����u �+*ն��=9X䶭�����h�Êa���DѰ@�uݺ���S5��S�֮��h������^�=\+�hl�+ ��ժV��v�Ok��Ns	�ޏVŦf�ʶ4Gjn���oc �����&$�裕2k�X��Y�w�����TZ�/.ָS{�Kx3lʺ��;�LJ��������!r����;G�=�Fr���Ԍ��ܱU�⒲�B��z�Ftt�:?�tB�rӐR	��{.,��Wn�G)'��:�<�tu��Ȃ��#)�����]3���b��Q�I�3V¦$�m�g�=ǟk}@��#��+ʘ��.��vQV����1ə:
4v�j��R�l�^));
�M{�c3^\�i���������p�U"���y��R�;y��y������X�أ�f���9�<�Z~RNE��Ju�����}%��}A��u����\����wcx�oS�"��]�s��W��inZ��gK��L
_m;��yj|�q�9X�+{qN��sm�V���-1W�*�M��ZY�:_�W�x��w˴���[��V�k�$�@������ Hl2��S��⤷q��׆�
�m>\D�t�Id��rX�{zz��e<�\��pi�<G�ۧ^�^;DrhRt��'z�(X}���RU����FwM��K���4q0o��}1���ⱘ�=	��o�y;��Na�������+�����JP�Z	�R�Tν:�k��ݬ�ͳ��ۜ�#&��t�ԥW�g׽ݵ�#�w�3�x��b�>��]N*kJ���֫�ݮ"��0a*��{�kf��ub7k8�P�C���Z���F��c�]}��s_[��«bI��d!e� ��20���J�t�t7��CH��Z�����[-՜.,��T�uىnd��^[�`Ws7G��:��e�"��<U�ѫ��$�Z�nd�aC�e:�\�5٬�hgo@�ȋʐ'z�=�O"���.�5n�B�U��Q��;qtn�)I<fVtUiΑ��H ���mXuCQ.�(1L7l�C���"�Q���!v��̽���<�2�>W�\�Y����7y��������vV҇�lP|�ju�%�����T�eL�����3��0��:8@�i8㧿;)T|Z��6[|���Ż���v��(�����&/��c[�����$��̅�z��[J�9�(Q���e�{�,��i��r��{�m=]��z �B����u::��7{z����X1\����/�m_%]�eZ�}:�]��ޏ����C#C���jnwN��`��q.\.��w��N%e��*S�0���8]�.^�Ғ֡�Wr|�w����9���n��9,�U������qb�5�miE��d�������u%8:��7y�X\���`��5Є���N�7gN�n�@�A˵FC\�>��2�ʛa��R�g��1d��g����V��4s��s�\]��t�F�*Y��h�r�y�� $,w6+����z����Nv[����ۋ�BDo1�C-��&�`�FsŐ���@ 7\7:W�9n[/~<�H;]���s�Uޣ� =T"����yG�pQ;Y�#yV9u�c���Wu�p�|���ƥ�ʍ)ud6Z
�
�9a[k/��G+��\ʥ��>��/�� ��x;�ھ䌻��E��^ɉ�f��>v��T��-�U�|:{vk_>(�5Q���u�(���
`i��Z����_D�r��헙�H,������w�#�����r9�x=��t��3 %cC�f��<�˵i���0����p��K
]��
1�So:���*n���D������R��V-�27�� R�{��T)�a�֛Q�<̩�xX�W���k�����]�}������]�z�7�`8bu)�j&+�%�J�N�+�X��ۼ�,�Z*e�k�n�E�����9+slv�+����h���t�u�Z^�8�QBq[�&�f:�q��Qg)(2O1?�gA���K5jp�m�At�Q�W��Tpu��=���V$�!q*��-�*S^uo.:��;��+L-�#;35�)j���ؕ�9�&r�Y�&WT����c��xħdU�(�p�1�uc�a��!P�_1�l�	�e�9D�Tx4eI�el�����Z.n�:шb1e�=L�����i[��)��R�錖�1��2�%�����ǲ�KDSE�^R�pEt����@[�*�8�]K��op}I]Ld�0z�t�a�f]��I#w)����:7�Z�x԰"��:21n��F��M�9?���wN����n�С��vf�%�	��i��������Ϫ)�7/y>Y��vɝ��͙G�����9% 8�Ķ�Ux4X���5��o��!�P�{:�
�isK!TU��{qK{�$놊�5�a�]oo����'��maAT��]���R���띹%×�FP$��a����A�+a������ۈ�{�Nm��l�krh��WV�hScn("�-�.�՝F޼�üU�5t�4Xv�Ct�D�s����hR��	R��4+ܖ�K���J���q.���k	�%���]�I ̒�g:��\K6���b<z ��'�/tek*˥y�bH�����켽�υ�WbPh�򲻵�x��]E)x�[��z�bW8ؽ�<���,����&ZiR��Ō�$]��'+�� 7��5�!u5�2X�X{�R:.�ۜc�ΰ�H3^�������t�[�Xz��+Gc�MǄg�=�ؖ��'@�&<9l��v��ڟ<V`�[�+:3]��Sx��1Y;���:=Ƕ��f�0Q�����L	*�%�\s���}�Uہ-k���T;m]w!�@���b��s�A5�=d3z�ٓ�(G+�]u������Ga�J �?���_}�}_}���꺒��[L]�#���2}D��zu����v;~|�p�4�ȥgD�Z@���(K�^���n��.Ε&��B�;.��ݾ�2Ȗy�&�>����B�)�����q�E��8�ɛ;_^��<=�w8��`RˠF>�����N��S�O�oj��j�--��У��7�����|�&���THZ�S�޾�+VN�u�v�+�d�������-�J�3j��.�q��m�烨�����Q��Bʽ궝`��8B.�G���c�6�#�atIr'Gt��TOl���J��H�d-�x[mlg]��4��7���L����2���is��m��Ӄ���_n�NS����}����o����.��특�JA�u�GK�6sŊ��
a�>��WjU�f��y�5%�F�m���4���E�[���}����7�OGVa�qk�p�wʞ�7t�;�T�ƫ��0�=�v�\n򄓛uՆ��c+�v;PwW7�ثI�;�wF���aONӬ�-���ngvSՎ*E��[�	�V|-dݭ�B�;���D6��Iܬ�>�g%dg5���v��J]Wwr9)����G��L�i%zћ��5S�ֹ�N��4�E`�h��Yw%m�W`Ҩ�5ܸ>l75��1VB�u*V�rk�<�y�-�?�_	Y�G]��N�N�G�tW�(V��Y��)4C��/SȓB¢N��Y�R>u��"V"i'�N��VF����9ir���gL��ӵΙ�覨eUI%OP��1L�鄙�-���Uȏ\�Zr#�\$�V�Q�>��GdE�qR��e*�T*�I}n\��+��:;���3��<
����s5C��FT(�l�M2*����+E�|�C��(�4, �Q�W;�0�V�W̴B�H�iʑ.��QMM
2s�x�ye	�GM�լ��bZ���ggsz$OJJ�妩�UQ�NR����r�K�E
w �7K.\�Jy���X�By�w'�D�HTNB�W$���#�7�xfba!��y��=�N�F˗
���'t�<��á��G4��C�J��^N9� L�+��(��R�$��t�B
5Ͼ�n��	u�gAqL,�ٝ]W�ɣ�P�|������i�W��m��e�J廗��S�ⵍ��P�xї�m�5���!��5N�U/��sĀ�2�չ�(@�ePU��e�u'G
/<o�X����^2��@�����lQ��݋����>��.ק͵��bF��.렦�_8v�X�Ϫ���|wN�Wb4���1Ѐ��������������N�){8Uﵞ]�Y�;�v�G��l/�^*:iר��7��_���D!:���J߆��U��ޕ.Ŷu��\�� �tP���綽k�AU)���{Ɍ~�VU{����~�z8I,!/i�ɾc5ʴz����Pm� �zP�H�_O�[>�P���a���`(�i���7A�gZ�y�v���������Z�^��������y5fv"5S�0T/jf*˟V�����7^�=gD�3�NZk���gW�"�}�_��=CEp��y�=`�@��8��U�e#�',h�"	^se��Y�x�w���ҳ�H�N�����ˢ�g��'�0��/ش1�D���h婆*�1��}��#.����o���/q��kÕs<g[�.� W hJo2�w��6�����#VuSMJz�
�]6�d��o�R_�6wMh~
j�[F�Iߌ�r45���;�����Q�m�Ž[��=�����V��J�H]��r��6���H�28;p�+������t�2p���<�w�O>�k�!�;�2�[��~�k*��q.�\��5j���?\j
7պ�f��mF kx�V��:�X��_mg/i��/+�>U�S��@l����q���]9��Z}䶇��c޶f���;e]G������[����1,g���EN���)���+f��:�}��T��+_ ���Ͻs�ok�ٕ�+���x:t'[R�}�t��k��Y"��芊�"�gǄ�J�d��U��Kt����\^��ٱ<y��^܇>��rZ.NDK�5�Dz�T+f Zj]\��@��\5�F��=�K���y�nl�v)豽\���o�ok���oe�����z���R�U����-�<F�{s׷��L_�U�"�p�4�Ō�٢P��C���#���y� kIHv�6_G����;��M��=M��4�)���?cu���0߬��zd����A�#r7�rW��'��]띅�ū����E�ӛbc5�y�T���XuV{�����ԫ�Au�����fy�G�uw�mV����o�-�00����@���]�����hɽ*�+� �X����p���Pqw��8w�GV����A�'.Xk�bi�����s6s���r6du��յ ��o 6>d� .��k5�.f�6���y%��͡6��r�x���g����X0��0Z.��@��B� l<�!=o%{ر�j����Őō�Q�ٕ8�j�����.=(C�u���5��޶Fa��V0J�DN�𼴳�G�Ϛ�ĶJ��g{ˣx}����^�~Y[�vV��"��~��=�:P���g��W��W�-o>��zE�mh��gY�ɕ�i"3��c� P��;�I׼�A�󬮳�q���K���އ��U�x���u��Mpȗ�ヸ�4��j�.��oG������ޓ)��Ob�O}�a�R�U�*�� L;y`^d�8J�~��0�ƌ*X�c�l�7hW���t�7��=�n�C���D�ܟ��jk_[��Z���w��������m�۳^~o����А{&=/K��b�*��H�d� j9��lS�\�U>:=;E��^�0N���r���sk�&��}t��݇s�*�D	�[�J1F���h�����~"��LY�ٜEz����� �ei��w�W9�]NOȁ+X]�b�ge{�9��#	&������ϓ���BeR�s��)��{Q�7�-���-rS�8��������ͻ��uh!�O)C�e�$g 8m�w�4�lꮌf�{i�p�ݒW�j�7�����ε�.�b�w-H{Ъ�3�er����\��%&��m���뼋B)ª@��-�3 �b�ۉ�����������:��8��x}',������o�,R�U������Z.�
����<)�@o��H���Rb�{Mf��d��� ,���sG�e"��b*��]�#Ն�QV��7�N�֓�!���A��������1IU1V��TC}鿍Ñ�Ḋ��
����s���(q�H���E됥y)'�nE�s��'��� {�'E���*��m��X��4[�<�x�
�\�ߤ�س��Ћg�g��)ZxJ��n`_ٴ��C��nle��"��s��j}�����^^u�)^I�F�Hz�}*��앯�
���N������'����WZ�ɳ�L{a���ʱ[5�6]q�Pu�W�sć��b�R��}*�yXG������.�io�/�up������p�\��#������_\�	��K�|n�.��㽸�lUnaUũ^���-0�V�[����ȭ��`>�|j��ҩ�3yADwyd��Zͭv�o:��.#�,�^�δ�N�s�Kz�8���c~ց0����V�S�'ٕe�Zy�,�G���x��_���g�^@�z���n����E�<�NF��e��:Wp;On�]}!p��h7�����em���I��c���D-:8і��¡1��op߶a���#T�2�U��n���>�f�6�'��=E�UG�&<.�ո�^x��1��?˳�[�65m=9���	�!� nS���Ǳs�
�q�h��JSv�����R�qٙ�~�/o�h�p���y�{��13���TB���ѫtW�M9[g���L�|}�K�����+�X��M]�{=d!q��O��}_j��f�]5O]���X�P@E��R�$?-���K�d
�p��>�����ǨR۶*�/93bs����M�2��\7���7�陖�v{��T<
�kD�=��9�i��Y�l�3��l�1	�93�%����9�9��Y�R�A4�n��VO-���G�z<f\i�T�W�`3�If���y�CY�U��j%��6yuM�u=�7���CtY��cj�S�|̞��j:���|���ݗb���zʵjX��rW�??S_u競�B��Z�yeߗ�X�����	Y΀�c���awt��"yx\�;2���\I]L\c�E("��%�Ɛ\����O%wM����.���~�9���*v�-SX�n��Z�v%\���e����5�{t<t�gd��P�]����iM�2����ewTط�ԱVK�����8^fx;�v[|��u9���Ƴ�{��i;��z���x�p?1��;���7 1�X2<�	�U��~'9)�3�L��ظW�<6�'c�]�o+umz"-�x�p�����7���hr#E҄��0��ș�^	��@�f��]|th��.&z��=���+��`��L�v];'��/b�|}/wv�j��_�ꝣf*�.>�U��Y�� '�h��0:�w�����ȿ$f�/�1p���R�������Y�;�����}�؄#��;7^F����P��%���R�Q�P�U`?�UXƷ��k��{�ok��ӗ^B��y�!�2���0-Vm�X��(f��lW��'�{%V�ƈ��*��^���X8Û�G�/`��>���׽W��M��"�a�2+ʙ�Y�!�����m���4�|�ǫ�z����{�;ڣQO���߽�<���h+ *��[�"~Թ"�d2�}�,�1e��J����U�x�W+N�LTX+��|�4���}PrcEA)�&�S�6�o,�Q~t _j�;O�Y�Y���8;����\0����}ua��f�����#t�tە�zֿfh����~��7��e�>h���X�+�c=u�S�Gع���ʇ^$h�:�a:�͙19��s#��\{%s�ǼE��vԩ˓z����3��:{�%�-��Ny+�|��WY'��#�)'b�y'�°�Xʈ�
�eҘ�'�f�ݺt=t=�ڼ�ຍh�2⭾����S����gl
Z>�i�?,V�W�_��,eDl�(Tl�P�Ɠ8ۘ�uOd�)���\�;�[ ��e��}�O�ppfXa��yO���A���A�$�/����$�gsbN����_�3H���p�����;�D�B�d��e{�̟[5��S ��m�]�T��S!�[��;Q�T�F�F�I��,5Fg���w?v��G��^T���T�R�J����|�i�;'�'.[*��m�!,��xW^��9G�k��l��s�<.��u���KG��9�e���C���ҷVb�o��O�o=(-]�H!^���z���GM�#!#D��V�&����}�n�������@���W�}iv�^�+/���
}O�x�_���w��?j�y�ٍV*���*�x0Ţ��� u��MpϢ\7�U��4�
����ȥ(3,zD@��}[X�eb�2V��Ʊ����r�앯�Azz�뵼eZ\+D�Ƽ;9V�$�]��*
�iزyB%�b�\>I��=^/*�^��۷]�r�]]���z�UNo�=�]�p`��B�w1��m�v�,�ԫ;cp��-�B���GC5�ʭ����5v1��N�R�y��hq3���N}2X�']����`	k�\�dڷYlV�#��K8z7�Z���,�|�w���\�g�зUo�@�O�%�q��}c:*��P�n��D�c}R�}�^��U#����K����m�/*$+�� $l�5:��T�]/]'%g�f���"�۔ �/%�9�0����#�4+%�x�Ȩ�T���Crbt/`nO�	��oV���P �^�A(�?Y��We�#�qj�w��+����������;�s�yM���8�ʖ
�m�aО�H9��2�����3�25��C4�سcW������Z��]��X��7Y��xO�R+E��^OX\4xR2���V�ߏ�f8Ven�LOU�Ǚ�0 {��ȟ�S�Y�y������pF9�	��r��+V��p���s��~�>5��1?'T�C&��x�ƾ�C��m��2(����~!V����Ov{�o���TB-��U��w�!��צ��D�n�F�A�-����J驃���cdԸ��Ncˮ᷄{�2����suX<��]�����\��`�N���Q�S��^ޤ^�T��5����t�z��>;�yu�������ќ��,ݾ�kTV�]J[
�n��+�ͩ����wj�X�7Ϸt�iX0�_gr��+��M�q��y�r�r_F�ڷ���i޺��L:�<cY�E˺��y�e����1|@�h�^��������OOsۓ޺lVt����gn>:k�f��o�j
�^n��UǡB~9W�sć�&3{���w�,	~-��\�(�������6\^���G|���X�⬑���2Ƴ��`�#���Q��'���Uzv�)����d��W�� ��\t�l��J����8}�NVS�H�g����RۗR��^��ۍV�ߌ1�7�r�T)�lVmPGfs��^l�Z>���cp���"���@?�0�Qe#�b�u�tƭ��GDx<,C߆˒��M�H��1kۉz���X���/TG�z�X�ͱ���0���#�$�=��W�w�=�L<�xm�)��h�-�Ci��Sx�Qʒc���2�R��y#'�j���j�y���X��[W�V���sQ�/e�m�҇%��r��NOƪuq(��X�է;mY�&�.�Ug�����w����bҶ|��aA��A���`�� ��= �����|r�03ҳ2�6;��][�$E)�&�3;��*7���x��%}�iwΎr�Yz��{�/z^�>c�m��ۛP��e� %{Y�䫴�˶��u��q�_��Ȭz�V�	����Q�s��i��[���^u%I���w����ͬ��v���z"����x*���KN"����S�>���Z�%l�zx���qy^�˄!N*4k�r�q
�O�Ѐ}�Ļ�g�'�A�r�2}�;~�J�aٜi�;��\zt33Q,:�T+�����K>S,=��@Fɂ�b^��L��7��Cӷ
��}Y��h�O<���
��xNAU)�����a^�V#޵�܀�6�;���ݿ:P|²q3�G��h�j��7|�(�\�T�yL�����E0$%W�����l�Z�n{�U�@�=�����{��{j��k�ּ ���L�IV4�8���O�Fz���(�vv�d*�{��-5Y�v��U�����H�ᴇP�f(مj�y���P�v��-�����`�ƣpܡ����Z-��B�p`;~� }��L3D����3��J���[�g��Tߌ��X�1�ꝣ��B���'PY�~�)�YHA�����9Z��[�ٚ�l�!��0���#��.!�����a~sg��yY<il�ނЊ���M��E����=��>����[�Z�5㽋��^ӗ�0D}�ZS��ǐ11@,�T���:On&F�c���Z�K�+�����m���=��4�貶n]�Xkv��!U��]<�����k��)�B��^�r��:�V���k����Z|�FQ��u�M���y��c�(.�bn>kU��FZ򔄚}���gR���j�]K�Xzkxk�5�3Fd��q��c9jT(s�B%=9�� մk�r�]�s˚��w��ٞ����k_���l䲺���ek�A�:�Y�3~���}q� �ǯ�3�6ܥ�&WQ�y�[��%>V��t���K+zh��%�v;������l�5�H�aA�j��,.��*baa��`���W@wx��cu�����6���B��I0vV>���
�׶�=�φT�ӡN����h���E��K1�7�f+�)u"s��M%|/qkHQ��c^�%8de϶!H�<{�rZ2���$��ɕ�ۺW���_��L)a�d�9����!�/��ǺD�����r��Pl�8��9��.����w�=ݼzu�jd�F�W8��S���ۧګ_&E1s��{ʅ��v;�g�Bʔ�܅���a��Y��+D�h���2Vյ��Wq�e,��7k��)��ւ1՝o�$���=JL����6=��ՓV$_cwUy�v�εv�}}4���_gn�ڜo���#�)�u>U(fh��c��;�񣖊7�2x�n��.���u�*�#1�㯅���u��b��vj�@�anc�t�^2n_ m���0J���"w:�k�Bm�
\
�� �x	][{�2�'��P�R'�*L��	˺�Ř2#Vټ�N��ܫ�+�G��K�M�[�voq��&�#p��S$��,TC�q@�W��\�Sih3�-1c��S�"5}�kzM��ʂ��_���K�[g����Ԧ��}'���Mz�g���49��|F���XrH��zo% v��D�U��������e��]W����V���첮k�+��/��F_VA�i���r��rqn�ڥ)�Kh=�;%�C��x��)<�j� |-ۚ��c�Y��+_�V�� ^q�ɷ�[u
�65]<�� v*��rvHxۇ�G�%ݩP���Rk�]%W��Hs��,XP��Np�Fr��r�����â;�9,.-_IT�]:�A]���v��:����|�I�v�j�\��#+�fTl
$)1��KG�#�dż.��p�Q��͜RS59`+8��8����3�/w^�O����1��Y[�6Ջ�?*W%�������f���tƩK}��A����m�v%a`{}�x�w�-�Z����(�4�\���cH�ū4F
�X�G�oZ�]�P���<��H����뻌��@w|��qV�?5l���QW:�L�pRh!�J�T+6�Vrܘ�
��$~�G՚�^���qf�A !l��J��S��J�C�HŻ�0< "���D��Dz��\w��7��%#[L[�w3hU�'e4��^[��Wr[V�u_S*P�o���\/�S)]'�_t��wk�-�W��1�(;*��P�� AF�"$� �"I�h{�z��QGTe�+���*l�?���<�˫B�aJ�UTU��#��ݢTfQ�wu��#����K��=�k.ms9���ioWR�0�-ֺ&uU+�/v8�&iYҫ�UK�7�NTUQ2�EDUV��gH�"��!����!U�:��s�f9x�̪�˒��(����#�����m�J�".�&$��QR�{���D�Υ�K�)&�I&��$�3�]Z&�Bd�A���N�]%#H��"��#���#�ӡ\��㫙AUN�8N�*�tQ2"��S5�I���,�sÙ�U̉�/}Y�9w73�)�Ģ�ǫ�3ts�(�G3����D�J���O9PAb�ˤY%Q���IhDJl�o����{�v\}�b�P���WsԬ��u�`�����v��(e��B[�{Tޣ��r�i��/�PW��>�)?|����
���wl��_�ro������������돤�8>�������h} I!����<�~8�w����~��C��_�i�ԓ�������}"#���'���5�]���E������9S?�I�����oϞ�p|w��{����0��?>���~��5��W�8�O���}v?�O����O��$���C��C�����&� ��|CtFG	����#�;b/������������.�~�s�ο�ɿ�I��o����@���+�}}x��	�����?��r�o�����N\���e��(~��o����W��T_O�񏠏���	|��*��mߕ��!�>�
��$�A1`�������$��U���'&�Bpx����r|㟣���O�ӧ~�G��o�䝿�ܮ��i����P�O�~?}".:��X���" �煮�+brʚ��/˷�T�}|G��`����G��y�p?>�߈y�q��?i�շ!���|���>&~������������&������������}pyG��c�P��A���
�D_b}�po�D�G�B D1����""0QX++m}`�W�UW�^5U��#E7nE7�H�_ԇ�ě�	�v�?#�.pr�����q?�����i$ߢ@��,�@>��
��ʵ1q��ݼ����� DDH���_H����H}}��ߨ~��}����I��U7�}n�t��?�ra_��Aw�ݷ!�>��O&�BN|�9@�I������@�!'��=�`�'�_�-(����s(��΋�b�n?{��"4DJs���}�q���>���﯆>+�w���܇��8�~�|t��ɾ��ߜ|L.�M�y�>�v>��>�
����y7�	7��A���9��}�@�I��U������T'%9y�]!��DD�C���������i�����7�����Y��iߎ?������ ���q��~v�'���������HO��s���`�i���_�}����&;�p{���(}������8��Z��ZC�Bw�ܮM�۹�pO��}~q���	'oj?Y��� O����������O�����i?�������ӷ�����|C�O�}�w���O!�M}�##�~��}" ��A�������Z�jZ|��&(��5'U�;���/�{r�wU�+����Ob�>�A���%�S1�����_�fs�ĳ�=��]~��آΕ�:�i��}�K�����P�9�\��B���	��֖־=!T���96G���v]���r��xΞ��p�]6dV{C-䶪��O��� j�^Ԭ�}E�$DX��F*�Dk��0�_q���}�����nL/������}&@�y�w���$��>������w��~x>��0�}���0�D���!����>��>�#�=۞\������"��j~�����+�������M���M���d��n�C�����������w���w�~L}!�1���>����wS��כ�}����ߎ������ݲ�M������F�b$|�P�쟰DG���}?]|ƈ܁�$�?�<�!��q���M���'��}��>�I�S�;���|v�������}�#몽3?IЂ��`P�{>�e*���A>������c� <�߽���?�Ʌߏ�
s�?�ɿ>�~�>&7������������~!�$�����|��~���_���ߨ�!�1���cp_��Y��Es�{���~8�W|M8�>���C�4��ۏ|���b�B>9~��,G�"�e}���������t���|�����v�M���;��wþ��O�y0��^�!���P���F'˄it�7VT{�A����
?!��#���"�}�~���O�9���n\H.�Sw�}�	<����>���������'���c�r��>���'��`�r�H��H��쟾����" =�M����/��=�<}�s)/(�ފ�1��G��;�1>��s�_����?�����0���G��7�~'8>�n@�I7�?��#�D�����`��G�^;��|��DD1�~��D1���S�� r/�o�쮔k;�"4G�D�#��~�M&�'���P};O�A�������眻)�P����}����;�7<��{�<�[�������<��F�" �#�+��_`��	iBu��`�(�++_��Q*��"�D��"�럾/����9�����e> ~���?ǭ���^~w�n<��i����?�O�}��?RC�����I��"���겇�>�<#��!|�P��s�5�`,ڙ�H%���"��w}yL)�������NO����ǿ;�Dp�B$}�UM��@G�"4}�yQDH90�ϫN�������?�$��C��|@�I7������;���ߢ!U�{�;CJU8�]]�lj�q:��$T���T'�щ1��jjE}Yז�H�Q����:I¤��]u�!:���N��n�~�>�y��{i�3u��z����	�ʌ�]�3R;�:w;��>�*3���l�������%~�$��o���N'��m��q!���'?���t�!�����]��������C�,\��;��q�|�g�p}��}&~�n?ϓ'����H� ��DC��tz�����L��e��q��'��������'�9������>_�Nӥw�k����<��	�O������M;㾿�O"���=����������������B��=����D�n:Y�w9'�Y��֨ލ�<���<��?�;����������s�h�2���x���_7�b��TɌ��d*�Uc͠�55x�E��V
�V�vo��-���/���S�ʅ�.~�C���OU�+ܺ���*㒇3�������\���T��s�����W�+�T�덤 BC%/�D�c�9�hj#1�T��v�:*�eΘc0�r�X����ÙB�%~2��
�$p�<�~�K��FpڊE�wuχ��Av���W�/{P\��q�'�__\�	��~��x[�xa9�p���r=�J/q��>|<'�w�׻�g���h��(X�\@Jj�L�h��z����͹̖ ����a-�+5�a���7���#�e��L:>��+8�o����˝�y�����`?��)�)��[�65m=1�s	Ɯ�%]ua�^����d���+�Pd���C	�����������!SY�.�z#�����E�?{�6+�����v�V���Ço^�ήT�N��em�磖����ɴۧg��!�-s��� ���:���\�ك����ݼ�ڥ:�X�?�Q�7޵�����\���ͱs�o����*/q�x��X���ǎ�72�Uמ̢(�Z�^����n�q$�����;�����`����i���ۋ0�xP���nizs�����z%~B݌�F]�K��{_�*���a���S5��⹬AU^p*�H�h�ǵ��g��A��O%� �� m|���:�(�0°~L���۷��Y��ד]�%p������rIV���"��A�>th�k�5��T��B��"�c>??�C8�I��V��G�if�,�S8k����d���
�t�f'�n*Y�ULSR�k��]�}�u�y���.�� ���3�jƓR�֬p��X
uV��?J𜂪S����������fЗ���\�V+��%�2��E�y+�|m^B²��U���z߀n��Y�����چg�3�J�����u����6���c�	�U����k�ُ�
����x@�\o�O��Y�;2��o߶������W�߻���k�&{@��^|n���'���V?X��j��T���tA��b���n�͠�RG�J�:�.�OX[�f<�q�K���Ro���,�m�NƠ�;k
����X�#��'���ղ]��6���\�G���gY]�t�ϜU�]+���Φt��e.�|�}_W�>��;�~���@!���	�0������r������f�C��6 ;+�h�R��1�m�Kr�j�S�ٔ~�0�O�	$-/T��0�|�錿��,���@R O;q43;�ߎ��:�����m�y9�ɘ��#��U�B�m���5��6ĝq�M_�v\ZC[J��k�ݍ�=u����{�w�յ��zrjL��|-�+ Y������U֪b�?���x��p��g'3bU\U����Xᗤ�:*S�[����s��_�΄.ڑ��3p�>t,}��W�b�Տ�v.���X����7���2S^�˖�/�����W������!�߭�(��HeG�&:�YT��٧�}� G{�ձ#��bg�a�߳��fև�=��ϗy��޸C�n��P��9u��d�k]|7���iu����������b�p�Zî�N�c��fv��vP
6*�Q.�5JҜs���=Kԫw�VKV1W�[4J�EBr�"��u�n�������$Zՙ�ڸ�*
�Cvui�#�����)����6]5cŊ�n�F;�e���M0N�<�����jr�4��cB��`�f��	-��8H�-�NK7���娹�nٝ�4h54����P����ݮ��U��Q:�\SL��}K�<�����IHjw)�>�l]�����U���U��}[�*���yS�S��Ki�RBQ!mj;9!^�:�B�O�`��-u�;�2}>��:��8�x��èm�XO���m� 8�G��}��,�62MCs�3�L{.���Z5�b������h���wu�H�ˈ��F�vTk�&<X�E����/��(xG�{'�pxxSB~�B�yYϲ�b���ݐ���-,�F�e�[�y>ڵS:{2�h�.�^�g�^�D!?��gһyߒ�+z���n��@s�!��u%|g֗���Z��y�c��l�4i�b�/|�=��V<���P�on2ߝ�?_ނ��Ct�uVD+}��V�p���n8;��M1}�q��}���b]l��*���A8u����l)�\7B��bl�P6��/2u%Ѳl��:m��btj��B�Lo��
u�p��t��	d�6K�ڟ���M���w��m��p{���~��ƓJŲ��ܯ��s�n0�~���j�Ȋ>�Ht�(� ����Nbm3���yE����l�r��U���]̞�֯��ݓvIc�QÏ���L�VBc�Uk�ӗ���j�G)jdk|�2�a�3V����vڑmv���\�2U��}��$��V76=Z���[�ݾ��Y�z�3nӬ;:��$���	�_D�}�}_p�jI����Wgn���e����ڄ}/N��Ƅ.M�����9()�U��������Nϼ6g��Y��J�xj�cz���=>�|g=�!3?{���gճK;7	�B�׭F��W����ѯ}�xHX^�+ʖ��H,N�H9��2�	��+�m��NRI�3
uz��p��л�:P�}^��t�@�J-V�_�sI�3hݔ!�}�Can�ɴɩ���鸭"< ��W��H�`԰D)%���f����eB���ə�kD��*ח�l`8b��ۺB�fK5�!�N���#�C~5�!���a����d4�\e-:��t� F��{�b_ͦ*��mx�A���GǨb6)������^�Yֽ���?T:������}����O�@�ϯ��)��W7T�8�<�^��/lP�޴�(ݡ�V�K%�<�Tf�����}Ϙ�j�E^�0�_ي�w��d�| \X���}���������0�a���泅�+��q�v�<9�.%~2��
�X��y��&
T���Vqm�p!6�lo ��|�C*����醡�m�:�0��-�;����掺��m�p۸�i�Xh�T��g���.w�w��.��,�eN{[�.>�|���]¯�Y%dBƺa�wgs�ʤ��Eȫ33�u%:�է|�qBm �_n�%�Z��W���W�[K۵��/N՛���l�>��`�qZ3؂��8�9�u���@\�̔������T8(Of7���x7���K�<���-�X�p�����������@�T�@�廵7l�O�E=}�E�-����x��{3	^�Xo�c|n�"��yC#riϣ9�LqǬ���|�g)�g`=�H�ļ,�U��A�wM1�-�kk�y�Uj�^}��|�����#,Bx�����T��b�d�6��o�غ7�����W��tk�p=�èY=;�δ=�"x�����>��RɅxbZ>0t/eT��@�50yo	�xo��%ߖn��������U¦�wg�V���Gܥ��U�Y/�(p��Z�}n�#2']7B�7�y��f�B��Zo⥈5���X�Ӳ��3?g�c@_����e��pO{ެW�R61�dŉ�`��:4s�r�bY'} JwNL�Ig��o��;啡B��U�fz�d�eZ�)ծ�Qa��\��i��O�Ėj<��x��D�J��Z"���ܯ�D3��)q$.�<A���V����W�hF<~����1�����uK���jD�mZHn*�v����i��d�鹎�Vp��x����q���6뮱L���O���{C�R�o�gם�>�d��x�U���U}���:1��}Az��/�Wz�AG1춳�w�����9(����1�nb/�Yyؚ�;�e��L��l�]���M׫݅�1�[��%x3
�õ|�(��4� 7^B�����x���s\2��*�@~u %����yX.!����r0�+�:��^��(p�2����Ûdz��ޙw�M\1Wg�����d&�>[�z-:M�uoވ�f�/�W���3A��=:Ē��c�\x�f B�<�	�S��gG���*t�?z�1qيՉ���yY!��OSNW;v�\��K��xo�;�x1z|�k;�����(���#����7p�תg�;����(kp�UZ�<,�����}����=�-�u�^ҮPYy��{��DY�/�W﷩�{X�]%��k� ?�[⥮�N�c�w�|5�2���H��U�z��>k����CB���,Cf�%�~�������s\��la3iH�=Ƽz����7/�gc�gd�Y�4E�<�!�/]�P�����g�b�?e؝.>��W��]ܥ�[�<���],�V�|�?D�
I*�0�O���~��r���^d��4T����u^_]{���S���Y�9J�n��z��by�n1�,��I7z��}�+��̵P��u����Ĝ���{-+�JK�tׅH;����3�GQc%w6lcw��3��}����Jo���jUv��LW�P�"f!���d1���*u.HD2��9U����%���jm�Ϻ����O2�*�gca��m?M�Ж���;�w�!�ꠀ�Q��Nś�k�� ���;�W�48�-�Y���[BaT}��L���ڗ��93��q�[���;� w���X=E+�7�'~`b�Ō�٢P����|�Ԏ�*(9wsv'P�sR(�s??\� ?��-^�=�n���$5�j��8�3�A���v=/G�V�bu�7:<ޙ8@���l�8+k�{f�KR�zC^a|����m�OR[im_?wo�<~���a�~� ��&��e�3c$��ʠ~�Z�R���eW<hZ�!n��������}7���������P;���@Hb�����8+��¡��3a�}��3���ީ����"<�0�'9V�!��a�uyҀ��A
�vu{�~n��;>���7
��'�����b�v�}����J�ʴ���R��ʷ��YUu�C�g���uPl5zkt*��(we枕� ���C�g ��F[5�%Ջ� (h��Ǫ�1W6�;/D4f��14"�q��}J�ܷ�M�dR=+[z�Ezrb�6��T
:G΃[O�9;0=]��+�X�W��b�(:�!�Ս侸{��x�T;
Ve���)�M�FV�lHs�p+c�m5��32oZis�=���3���3�V�kz+��@Mu{C)�=�����nDF_o����;Kx"���& |9Eg�7���^�28���J*�Cڡ�a�vn��6�eZ�������6��2�յ}�Q׆���#W��a�z7sU_�G���ZO-tr��7�G��q^����G۪&pղ���XwXx��>�ADc�x�ZEu
��*�Y6�����`�p���]�ԖQ�/1�_j���#e��%�Ú8�]�6�}Sd��m����_;ÎgS��(B�)�r�G�r��u�Zk����-�QC��O���a��M�
Dc��:�Ϸ�<-Ev�g��.Q�L-����M�xP����x�(f��[�V��<�{�g-�H{#���+��^j�+��ӽ��ak�S����ȶ��y���J�p��Db���:��×@Wɝ�g%��vV���5o:2��.�b�X�p�7jm�+.����+Uu�wq��i�U�2Q7���k�OX�<�$Bk�-V���h��1� �d+����(6q�wK�]�;ɗ���V�]���"�#	J��ݓL��E�o����uEY� ][��� �%�,��T�=�[���)g�Wp�ѓH(.R�VZV�X��j��3�u(�h'1��f��sY�\�u�u��o'M�k˚7u����I����,�V+�tʐr\*O�vJT�Y����o/F��Lʲr�؃ڽj��B�����P�v7�[ۘ��"�sd�b��W�
9n�=�Ӹ8�;:U�P@��ϲ�z��1sZ�f�U��|��t�H�/�&y;`Ь���7\u��]	��C]� a#���1mJf�h�jгE�%eIg-�Q�<�[�+S%�أ%˺���9�j�o2�����/O7asv%aT��=�퓏v������t�yXQ*����oۂ�.�JEoRšB�G�"�����ُ���@9j������d'��e����61|��2S�T�K��I���P�m,���`	�\d:�ߌ�!	�.��B�t�^�K�*�Q��j�L��'�b(�Y���czA
'*f]0��E�����|kOm���At&;�c�=Ŏ�廙
�w�� �]�S¤��k�����R7۩�F�[��ś�PQ����.<En��Cq`��
�x�O���-������`L�x1���j�y:�4-K�$��[A��8��i�2�1bް�lF��ǥ;�Xk������+�8s��֭��t��NN!p�Ի֗wTټy��|�+֑Y�u%C��۹u$T���Xat�C;���:�j��w�{�r�I�EEWIk�ʞ��Iwwq����$����$R�QrGJH���r��a�\�uܖ�VI���,۝��H���3z��t���u�QeY�b7Du]q�L>��U�<� �"(_#��������&�\���G�9�'IM�B��Ť�"ֵ1H��#��.�"!�9�R)�ui�sSD��UJ���"?=�oWR����.N�;�I��G539�o���$00�R"̋7�z�r"�+�TY�=��D�t��(���FF'��BާV�M�>8!�9U~$�6]ZY���Kڜ�����Wq)[��2��ؘ�T{���)r�!P���	�UWQG]�C�EV�'�<��QԾeɾD�Zj�<�s֔DsER��r�;��>��&���[�A퉽/��#6�S��
��;[L���g�iOo�to�Yd�sv�3�2i���M��i��U%�o��}�Wգ�;��r�����N9�%�:~�~��* !h��rX���%�\!<7ێ������&,1���Gt���9�����f�xy�Ƀ��5VJ����r����x���N�iێ�3;m=��Z�˺�������X�׶��u�N̄V�r~K@�Z��,�va��d��∲�\��=�T=�V������g�a�x���̬
vX�/*$m�dE�������e�x뛈�xw�t/�ѱZ=��U��/��JRmqǾ���Թ��^D_q�/J��2�|����nL��7秏8����J�;T�v_ɀ-zz}�ڭ����!��ي:��>�����2���A�
ĺ��K�.ٗ$
��ۚ^���,?��T����r��b�+�|�|�������ohj�껜�)=�c�ޯ8~���/B�ZǵD����8���E��^XM�ž��;k�,{~�F� �x�)�5�5A�����)���{VRy����g�6l�^�Xve�S�>�5���U�.�G�>ԋ0��s,7��?�g��G���4{��`F�|�L��ɠ�av�k�3��iި�[c�2����,U1����b��h�Au��q�*�QdǢ� ��[[פj�V�]v�|[�ް��;��3l ^TNGG�
gl�Fsi�3(Tӝ�z=rf77jpv�	�!�������UjB�}��s��;��X�`��G|b<\ÿ�f�0&K52�Tk~���ӯ�Q�onw1�Vi�Z�1��FE���y>���/��)Zx��,>>ʳ���׫zD�㞳:���\�5�O�7� ����He_ -zHy﶐ �5-���f�����g0`��/�N�%�j��W��2�䘱_6���̡u���]���.�gF���ޝ���~��o{�~��zy��סX3��a�A�g���_\���yt�j�
Ԟ��7K�ٖ5��fP���u�E*A��O�47�����2���nׇ���Ő�S����k�=���G>���ͮ�����s	^��Q��E]N���U1h�=v�wU�TnrB�y�!瀵~�!�{@?d+�s(`s�	�1A��W�cV��ajHo�x{0�W��^�|N�X�}�Π+�{�=�a]�σ9�<��¼ó�	WZ�����W=�����{�~UO�yx����^ㆎ����<Ո=�����)�%��#W�+��saF|������#���x֡(T�I'T֏:�M��͓��fS��3{�W����3�)>��<���Ҽ�OO�Vux��xȶ��j'[�]�zK�͂����o^k���Ĕ�0^֞r��7�C}9b�֙�]��"ҽ;��_T}�}
ec텒�m��>y��������
�T�|��O���Tj'��W��g^���Б;y�:�+�����nMi����(� o�ˊ�n�~C}����^�~z�K��X="1E70Г@���J���:���vG��������t8��<��q��}�%O[�Xj���3h*��9Nǔ�W�ۉ�O3Vb�R�'aʿWz�1:���-�I�Iy��g��{�H�����9O�0�ྴ�{�Ŵ����@=Qo���j�]��=���O_w��K�<��sޥ��	eW��^�2��;��FP�G��>��H���+��e����hO}:��;='y��/6��{�V�*m����j���-njk�����Σ)�.�3{C:����m��Y�m���@�2�{�@{:���{y�8���#ӝ�����Y'l������~"�Uƕ{����ள��/Zȉ4�������F �K�s�)oMkT�or����Զ8fi��-�J�*����ܥsZ��u����f�u�����+�`��Pz�?e��MX,(�����ZNU�w;ɋVݩ�6�K��>�ﾃ���Tϝ�sF�Wugh�@j�Mx�D��#��2{�݂�{�7���T��<��L����4���_�U���z�-�D�io�V��=�g��Y
ŵvDhI���m�G�}\ߟ2���������0�m�w�q¼�x�ơ���v��gT)�c|#T�,bۇS�J� �����*A�&T�`���G ^����)�cx=Z�Un�Ҕi�j4
�kΪj58�~�^���K6r&���SΗ��,���',� �_�����l۟Fx�3Wf�!��o�*��%�;ِ3�����Aƻ*�t���&F�zq"۳0�Qy:a�BW�����k���Q���|�e�Xx^�1ujK���Z<΍q���ڙsP��b���(�O:K���`m�Êf)�>��Xə���ۙ�]�'8�,���w����'�����b�qu##|�ݲ���#�U�j^�30���ە.��_f�w���c���"I�:��%�+`��c�Ń����Wm�S��ғr���@�ܡ�'_l-9]��:<�s�
w:����;�k�Dj��>�)+Z���f*ex�������{�Ihq���ٱ���6��O_�Ϟmw���h�g��S�L�Bs�׽>�{A�HV"�z����Qo�PuA��^woӎ��w���� �"��pWWge��Z_��g�=�溗;�T�����5��+cș�hͻp��n¨������-����:����-~�3f�D��hפ�z�A��sg(�y	�goǧ^N�l�N�U���/oa�U�:��1�8v���Y�sZl��G���^�.E�]����	��Yם��$��9oŧq��*��q?_�^���w��
�BU�^�'�gqf��FEzYk"�;ײ7Tv>mҏ�;/�ݷ���'�{��P^����gYޫ�s=�u�"~��o��+J�����sy_��%G��G�Ӄ<U�F�b�CI����X#�=���rU	�wc��1	폚�}�,�I�Rغ~�Nu�:�SR�t��N]b{{lRx6Y3pw���p�*�8	�S�t�/y��� %��Y�4-�����i�k�#t��(n,��'�CL����ܻ;z�F�Yr-�#e�ܳGx��Sl��V��aK3'O���}_Wױ=���������s�*|�*��^5��V�ԝjw��hQ�=�N.-�Θf�\
�����z��5��>�}Ꮢ��^ϷH�j���{�������>/[]��~/י��OmLn���j�5���ϭT����]ʜ�X��Q�X�3������ҡN~^pZ���!��s�FĮ��tq�FdyS�&w}̫���6�(�n�Ңb��nr\ʺel�^ֹ��-ŕ7X�'k��/"�>4�-�y{i�
�Ք_���SkEP�qf�?�����U5�#���C����㫏�=R����{�}}�����N8y�u��F����/W�{�X�����Z�2)�f<	��i��c�2��5=G'SM�YI�CSn��W^zC�O���JS�lsT�Nmø�z�Dp�&�nT��;�>�-���Y�@���T
�Ez�;X1o2 �E.md��Ȇ�ỉ`q;��jP�n�>���=k��=�Ez���Wu���ί�JF�O6�j����ˉ=
�up�N�h��Uh:,a���
��k�>�'�h�3N)[������Lg��A�JO���������߻�C{�U�5������ΖH�"�F��g=2���vu���	�|_)��pI�c��uvj���r�;<6�t9��z����W���V����c���y�t���Q����{qk�Gz�>-�����S#}g����v�dx�s�Z>�����]w�����/n�Zܛ�Xd(�wP�65��O��uq��SU�E$#Xz�ǲ��.pU�U�@+5��ך���NF*��W?y��ܝ���)�
᜕�ĹP�T0�5�AxV�S�n�*�1wd�O!W�J#�g�q�������ק]^����Y�o�/�<8�ｖ��>J�[�ϑ�ϗ{*e�Bp��岑�~8�w�\V{Ih�k+q��W������)y�v���=2^�UY*����r������S��W[�@=Qx?'��Oy�ˋkC]��v�@P�O��9F�n���܀�vM|hK|�w�.����==&g���W�vg�$����ָ������JRPU��]�6�c����8gm\��X�9Rv�w)sVl2�`��코����z3Z[+x�T{��y'6Μ�G��諭��lY�zf�\��Qi�?C�SQ���X�ip�2�b�y��o��1��'#r�z'Mڊ֝'�3���ޚ���}��4<T�Ј'��hJOܡ-*ɫ9���0���u
rxo��ϗ�ʣ�fga��6�e�Kg��oT�}=C�\54�.Y�.�=8������I��{1��j��=4x�W�j9��qP�5A=���yi3��+]ǩ*�*���yslmC��P��^���_9x���+��Ln��z�&�ȫ�v��g3Cs��f��:�*	8�o��{�2a�N��K$�Ũ�L�͸>�gj�'X�e����ݎq����ߋ�o~���M:M�+p�T0j�:���B�y�j�j����%��i�^�����B�r~�S�u�u��C��u^l�L�qu����+��#X�U�/?0�o�޼�ꝶ^�;x������`n�v��V�{��+ĳ���i�Sl�m�tR��1J>�P ���y��j��?x�+[�w�.L������pL6�)r���0(勆�qF�-*{�K�ʹ�o�h�ua=Ą�!Y}��%e]�U��4��G�D}�����lae��u��ɼ�[K(�Y�{��?_O�y����Y�ݶ&G�nwm7ꨶ���T�Q�4�u�u�-c����S�=�[��;kgwu�q�.qƪٖ�Ȗ��wgs�3�6�5�'�`:�:ܔ�y�۠_�vw�j%�p]���x�l���W����AIAqHF�� 
K�kTW�7o�s��ؠ�[��j+�ܷt�D�ʨ�g�Hm���k�U���b!'Ȃz���S:��/Q|���Ot��~�.�X���]�b��,����0ߨ���>X��'��.��Lym>���o�39i�^~嚏��mFm�W%q����9���(/���o:��qb{��Y�]:��5�q~��Q����^~:��TÖ�ᔸ��"w�ĕ��p����3���'9\jc��ow��b�O��|�;ht�s6��bvb+W�>�#DK�����d*ֻ����t��P�Y��|��Gu,�כ�޹���H��V9��ŎXD�%�y�d83r�]-�9;��y�k^�\�����R�^��8�A>y�v݊�+���,�7n�m��+R��S:b�^(?�ﾈ����j���ܨ���E���,^���c�����L;ȸ��ު7^�����^�/W��:;�Q��wk��dmG�W;Y^��Ӝ�?���N1�o�>�盘��^�V�y����y�����mo��կ�\���SCMe��u"_ثMA�V@���ǒȓl���ks2s�o�g�S�ަ���L�΂5�j�k�¨�x&)J1Z�Uc_�*2~�Y7�Q�n�R��܁��f'��'jh�q�����r��>ws1O��k�7<*7E��f����i+\k��^�1җ������h4<��t�^Wut�Wix��v�$�R�c)w���~u[ހ����h\�υ���9y��pq�Y�G��&|�2���������_i
&�v�j�A�@>{����BT1�R�õN_T*��?#T�>(��]�5�
���C4mz+މ��Q9@J�B�8���rma�<���n�U���KDb}�_Keܼ�ხa���t�G0e��U�9���*�tcm-�Y0]ݤ�j�DrȁE�I;�`����<R��K�q�K2w\D���F�W�"I�MG�b0&"�{1i����Ҵ������u�r�jy��b1,[�������s���ե}X�*&:�$l�4R��>�[�%Ҿ4ɾ�;���M�x�{	�e[c��O9�>S/�`���ĚZ�=������V^jL#�Ղ�<�;�k㷊YW$1��!��mcab����u��˵� m��`ο������ג�m�_gq�:��z��5����tm�<Q��*�s�����8�������0�d�D'U�r��N�7��1T�m��h^�jr<> nf%����az�.�;e�.�7�z9=�^�e��)��쩰�(k��HXr@S����dͭ)�X����6u�� ��z��w_�@}-���꧜�.yu�~�)�@���w�P���J��n#g�Шr�]�Z�����;�
�P*�@{t-��߂Hlio3�`ǲ�@�TC9c��E�&WG�ۯn�ވ�Ԟ�Ό�:�jH��S�f�>"�/�I���r��V�G1RN(�wnqrYy��mn���(6���[E�����r�]�H)�S�Lm���Zkh��v���W\�n���`ܼTa�|� ��Ǌ������R	d�F�\�F�[j�t$�|B���t�0��w5�E���D�c���ˠc��b�}�X����\�6J�r�q�&�M�В����S�tz��u��@e���n^Sa���7w���D. �$~x����:���s��4�`V��lJE��G�V��h��k]�e�Ɗ�a��"�����/*�R��gwxw:?`ciwV�m���f۝0�.AH(��L�n�&�W9Ҝ��X�;�.��a�w�u)f�|�4i��o�P�U�f\nV�|�y7��@'rA.�����6�o��MS��|�R�mގ6����R뛹nnh@s��������e.�.��:��Ǭ�0��/(7I�C�vs�}{N9�As(�<��q˟`LRYg��w�Y�6�}���(�\���.��kL�d��u�a���]�d�]��ʴ�M�-�P�ok0`�����m·g.2��U���ق��7,����y��w�ܫ3�Ŏj��c�v]Ӡ�b�Q���pl��*�dّw�u��٣��w�t������+�Ш���|[�Ë[BS�;6\���;�Jvn7uZ��f4�U��蕋�0]��@J�
�uELh��Kc#����<#�23H+�}�**�R[� !��Q]�AE�TE2�*��=y�r	�(���GY�d������2��0*��
NS��'���.]ε�Ҫ�UU�:㑗��DW.z��(���>Yr2,"�DE�eYЮP\ޮҢOw�wu��=��f�I]p�
�Ep�E�݅�N��4�����J���"��³xdr;{�����y��/<�������+��,�t��it)DTs(us���������VY���2��*9j�E0��0���vQyޤZ9�^빯��="=ރ��y���Qȹy��$dM.+�#�0��Qz {���K���w]��ZТ���9�Uz]�Tq����Έ�}\�T���*H��yz�$*�Į}w�<qnK����r�}��Џ�=瓨���oy�r��+��]��R�\i�PU$����Q>�C)�'e��<Fg#j�n�3gƺ+�x}El�}��
M���4 Qi[�R�ob u���y;�Έ��:#��x�r���ﾪ�*��S�j���߻�{��v�2����寍%7~�Խۚ�o=�d���>Re��\T�I׾y�'zq��K�=�V�J�m��Z��v��z������fK=ӣ~��?y��Z�D������������6��In1�"\�Q���Z�h^�=<~c�~~ܨ�;�V���5��CҚ�ػ�u4wn�(��'�\�<{���\x�&v����v�O��2�sw�5;����|��W����u�z����N��,��g֖�]5S�wj�vT�װ؏T�}����(����l�B�mxuy����J���>_v��,���<2$�������ի�\?w*s��a��0��yu�����)>�z�9�P%�M���U�H׃R��W_#�&!0�|�w?��=9EKڛ��`�؟����}�����������5
\m|�
E�Hz�u�
�=~	��s�\��h0���WJ]6�:�ڲ�X�c�y���ۥǭmD���5�po�T�i
�^�:�7�4{ω
S�ȽA-���yP�P���J�o�x�!�4P<^
T��ou�1*�WbO�	t;�]t�� �+3e|xR=y`a	���N�����u�9k=�}S�)6��%tC4�_=���fmQ�7]�e�U'�ͯT�vz�����"B�f�X�K֢��~�5u���1sU�o�&3�\���T��/κ���PU��Wy82���|�;��C�_�4�e��f?yxF'�a N����<��ݦnw��kPt�u��M�����h?���X��N�c�5�n^��/NE�Ϫ	��ߔ��יY�{��{�_��ciC��Ν��;�#�s1w���ԣ�:�������ʫ�3��l��}w[1�=X�O�ҋ͔�{e�x��ں�k[O�}:xo��\}��fk�I��z5�������������.�D.ڢ=9�&��:p�ϥ�W%@�B/k����~ƽ��TÖ�95
��Y�Qek���n ��5�m������=T�|��{}�x���z���wW34���\{�ϭ_�\���2�K��iU�|��V�l�g{N�VUg�i������ǃ!q��8�����LuO����p=�3;rs����l�9s(���Yq+�u����g>ZU�L�ǘp�7��F:��&��Sׇ'$ǈoF$�:�W�qޫF�V 4�v7@������/�3��ꯪ��^����;e���>�_z3��~�a��̮������Q�:a�bƎG�˒����P�լ�Z[~����b�W�2���m�q��U���-A�Wu��>A����>��MY�4��Jh\��=/�#�>�[O�ml������鷾G�9�5��*s����7�W�ϛ~вm�����w�-��yt�Mf5L�K��S,�F�����kig���=��ʞ�;�B{�v�]��($��7�I�����
��b��ڂg�1׃�Ñ��WJ�°E��5q����Ns:�]F̷q]��g�۔J��v�˫R˷�m���/<��Jv��F��Ӏ���q�^��^��=��9=7,m;X��5�7�iÜ͸˜�ā��G�{��c�ߧ&����3j�ct�hyU-�dy� t���L|�I��X��Խ�����~��j�؈�۩*�~J%��$�ߊ�y�ܐl��5_#S�����K�e%6�i+86U�3��lA�
!��#���{:�a��sY�8����+Tk�����9:�.�b�7)E-<T
�=cd�i�J��}��D}��嫵f��y�S��4=EC�m����I=�]K��^Wў_Y��	͸�{�}y-�E�I���#k~���hrW;/W.8my�T�Sۇ�k{|c��J��\I眜x�yG��Hj��:�z���k(�!uT�*�g��-%���W˷�:o���ӹ���P�7�U��W'+T�7�Rl�����q½��^��U��i�4��_m�{��)��4�^�`��)q~�k՛�)�vW_����uӏ|_ӻ_��1-��o�۫���;;��)l�θ�r�Iz�/q߻�K��棪��'�v���k����dx�6�����=���u�u:�M�*��U�5{$�C��b��d�u W����1�-�Y���su�w%W8QN����E���	�]G���7B��j��Uy8i,����kk����I~ʋ6�h�l���2"�3ak��Ƭ���K��&P����c!8�Q�-c��.�iW�X:,��3��K��ܡr��Y@�c0�n-�W�'zz�b����9���鹽F,ͦ�'�ɬ ]�l�"�:�U/78_iB��n����hCk{,+귛u.��u]KZ"�����:�'��I:�W�cҝ���_u-R�$;%v19IN�����>�U&�b~S3��Y3�b���s��Sbv�k�.��vI��E�9�8��}�T��@f�*���ʥ�'�-�!�p�yKw�~��^��2�wo8�Su�ë�	a9؎f<��y��=-�i
.��j��.U-�k�y��U)�zk܎Ԉ<�ޮv���'ƑŴ��k�^�'��ך���ҪO!�W���V�r���Voyv�,z��ƪ����E~�����H�ߟ�kJ��өeIGU3��{Y6�ㄟ�����h��¢��G�=R�Uo|����]b�U/+·�:p�����>��	�o�{O%v$�G���QД�8�,�������q◞E��]�ϻ$Y�p/Y����,m���i�=�K���u:>}��M�o�>�}�G����T�~{]N�PR�žX|��6��uP���j⼮2.��Kw��,*�i��4�EE����`�Ȓ��
�n��5s��>-*�u��N=�Ct�[�Ԡ��}�18�s5�ToX1}r����^�L5��:�u5k�N�5��ɮ�Ḣ�$L3�V�q��P����ϭb���g������̔�띷u���~^��Z=P庍:�	l1��jn-��V��6�)��{�.�K�/z���A�{ѫ�~.�L6�߰�X#�=��u[���8V��Ld���Z��-<��jb��1�}��F�պ�1��4Ŝ����m���+��2b�e�@{w
��Σg�4�2S�n�Uޜh=^���t�P��k�A��|���2�����+���5�ף�@��cԅ%uu8��a?����i��j	�,�zߑa�^����t\޻]F緒k6��r]��:�f@�in�����1C�\���������	�ن������5��u�
�j<B�L?Cs�º��I�����	.�.�z�5�\�s�I���(V�u��.=+�ۿM=�j�̲�a�3��:e ��C�Rh;^B��֫�����R����:���~��ƫм���c`6�xhy|���K9J�i=4�}Κ	;���*�W�.��]��ƽ�ݷ�g.I�_lP>��x�F�\�0�3%�U�h�{�tV�˛VyWd��L,�kO��z��tT��f��Uӗ״�Õ ���:u�f`����Z\��sxO���5�o���[��<�&�}���G�*�^�vF��{B��Z���]K���-�o�:xfN��l^�қ�V�
V�F���3U������U����N�P�za�u�z�Vp!�Tw+η|\KKMz�^�^�ARG���b��VuU������72�{f��PI�b����[�9�7~qCsП�m��[�@�C%ۛ�t��u/lΜ��۸�RU�Q����6�wl%��eG=�}�K�l��_4��j��wd\�}imD_�TF��խ��ʈr�Asl�z���5��Bu��[��z
��{\#b�N��v*wz�7����oX�� �L<Վ��=�ka�B�C����W�S�V��x�������m��)ב����;�{��㓂[ơ\a˯�f'�5p!<���ڹ�����+�9��ޜ�����P/���	�q�����T�Q�{Dϖ9���	.k��`���e�}�]���������¥�ۊϳ}�ϸ<)cU��-�eoPC�^_���e.��r6�k���%[w�N���%۲l=}A��J�u�{*��q��p�{\ӛrћ>�U}�W������w���O}�����k�̷adLCn�/�ھ%{8`��+�q�K^��������f1���Zȴ�:�9�ae9�	����p)���{s��5O�َ39��˜�lQ���Nͨ���xT��`ՓܷtfuO4���z�;����oȂz��>��Χ��{��s�[�Ş�M�>]�~�,����P�^�m����Z���K�v��yy�׃˓��(8�c�����p�������^k0o�����\�W5q����VeK׊�N!���E����ר�%<w��f���|���Ѯj-�xX�9�23��*{ռ����iN�,�W)W�N�[���{���	�>��U�9H���:w/{w�d����P��҈��{�C�g��ζm4�n��j�+.j̍�b����2�[��W������~�i��{����q��Q�?z��u�ř1%���Dl3~(���E�$�C�Q&�ڼ�Tb�Җ\;�U��sqԖ��We#�+�~��Y�h)z�z��sʲ��-��cc��q��v+r�wu��]ԩ���830;2e�:�+Qӎ��ݷ@Μ����-��F��cgK����r��UW�E��k��KDMz}���r�BZ3ay����D��7��S��GW�[��{Ҵ�����[���(f%�5�.�`kjN�����Vz%n�=�3��,����C����Q�����S�V�E$#5��C�kiC6���^�ŏ3�{TY������c���-4j�T��f+��H埏Q�z�_���kMT��)�nz�֩!+�x�a\�l�>bf#\k���
��q^�&����R���2����}�ߍ%�ϱ9͠�9��̧��ʺ��X���U<Ӳ�ݧ�ȟަ[�Y�>�Y��q�ި�??b��m�s���)��j{WaLu����S�f�{��B��z�߽����>5H�]�ٚ��o�^͗�tjW�:n���z'��U���%pc|qrr���;�~β������/?R�r�?P�v�mN��^��W�{]�ۿp��<���uS|�-�����
4l��s}�OH�:���f;w�Ⱥ�1i ���!� �ox	{W$�}Ϻ��͟4��תL�*�+���
֚Is,Rbj쾟EZ}�]�%M�t6'I�����iE=�Je(���X8n�2�e]Ᵹ����
n�0t{�S��ۛ���}_}U�3�伞�-��~�!M�J������T�?{�N~b�9S<��-���B�r׆��V�lb����^�T�醷�Ū�x����d��1Kw��ԋ8v{��:=7��r��]G��?u=��}�����Q;��8���Ŏ��Q~��{�N?[�~�l��\�����ʴ�f����Y=�A�����v2�A'���{������	_ц�T?\mNQ��l]��k6��Q�z�]&K�mT_���z�W��~.�M|[�VJa�Ʒv�	1����~N�����eض�n#�yj�z�U�M)F�D��+zg7O���cW��)Fim-�W�I�9O���Y6���7�ިѡLl��fie��e׾�+��o���-��O,����?_�|�#\�t�������75H��\JT�i|L�c�ǿfx�й{6�����u�W^�෷A��R
�Y:�ʆ��*�j�Db7�ח�XOm�u�^fj�4��FDR%�Kw0h	��55��C�-ɕy�}F�n>Π-�{�SBu�ꕠ��3)7�.j ��ž��������dU�K�[�WV�c�ʀd�i�%Ց��f��BԎ��^�V
Mw#��L�����v�@��K�Z�3�OXn��K��!"7��O�5��T�u���Ӆ��=09�C��-b�lǈ�6� N2o�X�J����,�!B4r��)�:ޞ�Q0����u�ǯ_.�H��[��5���(b�hWSn��fc3�t���rkC��vQb�sr]؆��d~`�8m.�8�ë�}�g�[�T�5�ʞlڕ�#tJ�z��	v(͕�]q��uoE��7W6@tx�����h�Na;YY����pwZ���[�@��g(@8��3����+���x��fɓ�F��u"�tu7wT������.K�^ԩ��.��2�냉�TW�nP����Y���c�w���F6f��엌^3	��0��K�5a<��1H{�%t:v�L6)Tw(�B�"a��}i�Fs��:](��G�M��k2�X� t����ɠ#�[M�����M河�)]�@S�2Aq+@M�v+D	��]���јf�S�U����,$�#6j|t
��ؖ�黩+�\ƺw����W�R�;�a'u��!�5K$5���M|k����/N�}�a�*�͟��Hf���+]���r��;q<R�ʹ3-��V'���2.�1%\���)}P�㜰r �Y5bY��يJ}[��w����R̡��{]K-�5ђ
�37'@�sT&\�h�6�n.��'��X�7ĵ�w��\���yu`��}�X�����ԅFV��]�V�e#tp�]+z퉙�T����)��\���>�~�n.�+a�,G/�P��闹{�6��n�)�n�T]��wםa�spތ�7[y\{Q���RQ�y˳���4�t)V,��`q�5���Wt�]@d�YY�����셃I���ub��v��.�!�U��˯V��)��K�Dv��^#�m:�`e���X��j�5λ�	SH:���`��͈�w)Ǻ�If�{}z�I��,�M�2q���X�����lf�eu�]��s�R�n_I�Hg3N�3�86hjyI��w:��\�Qd`��lou/����2��[ս����0_$�:v�Ю���v��!IХ�KOɉ�&&
8o��`���:���̜�&QV.��ae�8�Px���H�;�w߬�}���ö��:�՟556�R��n��U��f־Y��ܷy���nc�U�^Π1�]za��"�٭�ʳ�˅��8ɼv:��X�;��,�%dWU�\�>Ur�a���痵j(�'u\����pSg�+wvw]՗��/o��vDٳ���T*��VVFi�S�����zۚE��Z6�J�K�X+�	���2����99�0��]'	���'�����s�"Aw'�E�2�y$'
C6\39DE�:H���L�J(�hjI��
p��2+��O��i�S�z;�.�ez��!�QfDr=Y^���͐T�"�B�;*��,�Iˇ��i�K.Rz�DBH��^c��5������޹�b�\�R�r�,P�e�}�뻂J钅Q(���(��9�!�*$��D�Wz�W(��'PԮ5��k�/�2	���K�+��s�L"�Sn��T\9*��y�xBB&��J�rq6NN�LU%�%���8�:�NQQS�dE�jg�Ȫ��wXS��*�Ps�����G���o\�{����]�j-�%\�J�
)!�teU�r�J(�W
���ǯ;�s�*/^�T���\�Q:(����@|?
�P�i��-��L�u	w��
���MO�﹋�6�uZ9�o��K�k{B6�����%󝽨��K������.�`��UW��ǐ��%�b�{��������/CRI�j�Y��h$���X�xF�<�f&�K�N�����cj�i&-0��v�=�NT�E��~X��'�A��;4f91�W;����ſ'}K����*�:��螟�t���gM�dp��x��M�g���k�Ib�]KϨ������}��^w��j��n׍2�evs��&s�{�3!ڗ��m��Z���ԻX���:xo	2n���K8��=+�=(���f�Br7�~&�}�ˎm�~�=8�بj�u�������x�27#��f�8��:�EZF�uq4���k���%Ac͵����)&s�Sޚ�s��ѭ��װ�a�es�z���rsMeyy�ɛcP���G�ǣk����Gt/}ۏ�?T�s5��~��P�i
��r{i�L�~93�<͕�2�\Vlz���)�U�f�ݿZ׻k��Oϻ)/rU�y%x�:��{����:��3���7%N��Η�5�&�VQYj�Ѿ���l�å�s|��G�X^�rvy�F�0p��W	�L*mdy�s��Af�����9�jb������R@�Վ�]X�:]J*J9� �	NZ,��D}@c����ﾈ����m����ϐ�{�`���Jc����oJ���W����ޮy���3p]�nY˫��SBe髨e��a��+������D��D��~�kzi�Ǹw�'f������*I¨��b���ׅO5�UQ<�y'����7T�_��f'��n���ƹ�*p��-��� ��د���	�^e��~��s�2Z/1���l��N5��2�+�j�5���1Sk˱m�[;�0���$�P.@�؞̫��k����	��]:0��^�{}Awճ�#!ǧ�-]��ǥ��6�&�zۏd��W��uz����4]We���l��T�-�u_�u]W��k��mz㞓S���������f��
�i���A�͵B��{ƒz��k���):׾�˝�.(M�S�$��]+�Vי���\f���~���N���W���d���&lt1-�_�z���W�G8f+Ա-�v	�!��rg]�</9�d��i<D�����PT�->���ƹ�%hF�q���ee�E����2d�*;������[�]�r��Q�'IW��e7fN��=Rj���ޫ`��r�}_}�_�R��{��K����-��s�ӆ�w�����*�?%�G���-��+=1H%{���ZdC��ߝ���;���ON�Uow�6��hi#��=`������k��}��k��yV�3����{ݯ��]��W{�AK�3O��8C&}-�?W٬;����jw~�i��{����S��]���W�Wpn�[%����Ϫv��7�Ґ��+��n8��i�Hdξ�C���U���l�qyTn�
��Ӥj�U�05G&5{$ܹ{gj���t����޽��2��J~��� �P�{ѩ·c)J1Z�Uc_�\�c�yhS�7I��ڼ��M�d���Ve�Ϙs�;PF�6u¸y%_�>*d��{��஗{��f*������TZ;|rz��L�z�wғd���e[�(:�&��Cv���̇^��}`���ZG���*��?qt���DP��w�|��Ѯ�Cwk�7�D(�L��EWv{��K�v��S��Reoq��$*^Q�q��~��{	�73��VuH��kV#�#�`f&�֖�N�A��t�f�n�rӰ��83s.vի�W�ײ�T���\����#�x�l_�~sP'�K��D��Q��W�f��BK��O��cU�K�P�]����V���<�J:��f����:��~�?$��8����|x��j��+�c����>���X������������׹[W�һ<�x��Q+���Rq?{��]K���I�*��᳽�3y�/ ���[h}>���k��5G�]Jܫd�Ԑ�ޯm�k^\�]S����~���S�m�lx^�*�EQ�2�[Ù��X�����ŋ&�����W)S��E�݃��f��)�xZ�&#!�TMU,p�=��;Gm#q�p�\eު��ߩ#�p���(���ٵ뻟9^M��Ic��ޕZ`�{���uvMr�Sκu�/oWL���]���`�&�oW��P�O�Kv�ܨO�ԥ9��j��,��6T&4��U�Sr�L��0�=Z�DZ[Q~���^j��d��-�V�J��/2��9֤��F�hܧr����o!�b����eA���U��4�8̻��xַ����uDZur��Dr�K�����.��)7�����$F�W�
n07����B��}׼v��ܟ]�[5>6�k��m�JOﾪ��[*`�����ų9އ
j+�C�@�ᶡ��ۑ^1�'�������U�ET�q�ho�F����M7r���;���mmw���<�i���/9CٙY�y^��P_9U�e�"x�*��̮w�vc� �0�y1݇�g��t��P�:�{lQ�^��������Lg����|)S�X)w�@����}�VA���u�wJt;�3k��$��{�Y�I����=~�3�mwz�<
��*���4��uμ����a3�l/B+�+�g<��v�n����(~K�sT��n�M���|�y5��[�f��ki.1��:xuE�k� �]K�O�gӨOo�w�t�i͝��͡��+֦羮���Ĉ����,tB�����WW��b�O�)@;j����9�}K���晧�&�rW�~J�m�ݣl�ߟP�,�a�\��=�7uά�uN���P�����WyZ���Р�AX��.9\r����!#�'x�F�i
�o����G��
�e0�Sk2����c��c���#��p���GS��U���g��+h�Z�Ӽ�77�(^'}�5��\G%�qα"�p�������d�:��/�jpp��1��n9γ����5"R�gހ01�l�V<}Z����8�K�z����ߖ�"�uo]ƛ��.t{���0E(�i�w�V7��;�x���Q��}Ͼ{���oϽ���}�U�W��n'N�my��"��Rpʇ�&���V�w�tҏwޓ/C����,Д;ѹ��7'Z�̈́*g$->q��<����D՞��jR�;C���k8�r��ٰ������&)J;q���5���uoގ��ޒ�a�'�WÏF*��qr�i��n��	�,�Dl���S̭�����'C<�������>�ݞ����W1����]l��o"iS1Gc�蕝q�m��y�%�Ӊ�s3�J��Ǌk�<��N�W�_in���j� 5Ҵ��!E�-��B,.o��zɜ�9����<��ڥ_iӀ�	��É�b�J�n�����X���-�y��C�w�F2��gmx�`{'�ig�V�0ѽ��6IDWu������aZ ��2�[���}�݂�`���}ZڳW���
�x�r��&����ɫ�*�E����5����|�5���K��zlg�NmѬ=�`LǶ�����<�[��XϗP���Ԙ��NV��Oݨ���7]���Y�7:>����_�'�T�-�]KϪ%�=ù�ͭ�m5˞�W{�������^j�j���#�T�_yk����W���a���g���O1�T������]�w�䙤o��Ep���oN�4��|�g˽�{�'��N�9k��ӧ������B���t8Vz�y�,	��҃w�:���~xlk����R��q�[��!�/�7�϶�9���ܫ��/-�}U<�����k�^�t��uw�>�Y����f�(e��l$�!��y7墂�}�9׺���s���ݮ>��׍٪�LM�*񩭷[�{�V��y���s�"vW�J���yЛ=��#�,�#�����-�k�N���5�m|�:r�bl�=��gd����l~�S[�R���|�@Yۜ�aϻnN:]]�WT��EX7��xP8n:��M����A�>��ʝ��,�r���ݼ�H`�R�َ��W�;�w����W͌:���⥃��}�^_-.o~�mZ�A�s���‍��Uʌ��G�G�v�,���rs��������5Q���p�@���,�:��C��a��ӛE�C!\��Q�j桻�
�����	�[.6���%�3�S�z�E��z��%^p\o�4���^�!*���EZ�*��J�վ/�׮�m�<���ޱ��=�WxzR����>��ߍ$�R�c)w��_��3���=ܵ��L�s�լ�=�U|����s�^��w�f;��W��R�t�����)�`'�)^��/�Wz���U�G~� <���h?�����[^W���Y�j��4]<��Q�.+�;q_f��|����G~�+j�ZEY.����-���"��D��i�u�y�U�G�d�A�T�F�~X��bߏ���nd5��mn��)�;o����6�r׆ן˪v�ǖלZ�})⥨x�l�g}�c�p��\���?,���Y�\�g�MY�Qe��y���2��0�^ޗ]�Sˋ F�ìݷϵui�M8.T�S�ιd�'0Nj�R�]]�نk�6��=�4U�"H�z+�+ ��pQ`L9�B�x��.J����9�E���NWI�skV��� w0o��[�.+��Vujv��w��}U_`�2��=�~�ݽ����%��C�|8���Y^<�h��Dt����Y���
�y_�l�7�]�;Պ��vz=�g��5�W�o�����_*�6;���zs���uf0�z��Qt���������7zl%xa*eC��`2��͋�^Q�9+��E}M�kv/<C��,k~qe�)���[�z�f�1��?���<0�ȧ�=�k{�*s?v������kro�yj�q�4��^�;>7���Mǜ�dC��������eFS��~���9����S�����&�^�`|�wc�)�qG���j���
חݾ/}���I֓���C�2�qx����_�g(l'Q�����L5L�l��L�f:o�&+�7�ӽ��w�g���Ə���s������a�L/Q-C��L��-��{Wq0��-�Qi������^����LZa�m�+�{d�q����jq��B�6�԰#&R@@����]����p��L#��#�U$��9��dѹ�,;���5ӊ�]�N���L`��Ӵ���Ǖ�]�(]꽩�r������g L���ɯ�8��uҮ�-��r]��S!�t��h�����fO^���I�g���y��%� �T�S�����މ�m�r��n�����>�y���Qm}���-~?RX�1F:򌘍Pc]88�G��9�z�����8a������~�+n�Zc����K�v�����Ps:7~�+/uy�CW�����PI�k�'.m+5qU�͑��̽~���i��^��nb���7:v�L-a��k�u��P�8��N�{��i��s��r�6c\�gG���Ӎ=��۔|�5_l���䧍���;�wR$r�ʹݷ=�9���R�L5���[Tvq��>{��}#�E<��k~Oa�� �����2�y�T"�z����V����7��OHyzw,�K%�3`��{y�D�"{6�Y;}+%?3�[�F,]�	�\�_;�pf�uE';gy˭�;����U���}n�Ҕvن�0Ƭ�n�?z���}�0#2��NM'w~�Q-��%hJ��Ճ55�M��1},��XUܥ1[ �n�7�$	h�uN�Hn���u�R:��.V�ư[u�=�ÚA�����}pe��cdV�7IIZ���d3oZi�p���ѷ]g�/OӢ��ܭ��W����!�K2gf��7���Sͥ��Y�N���A-O��ȕ��D�t��Nf�7{�5*�C��*�����L5o�}���*���Ya[�R����h&��F��LV;��g�@Ib3�w`c0
���|m�G�)���pp/-'����v!��v�K�ʐ�]LU�����d�a�{L�\�=74qf!�sz^�N��B�s��d�|��\���ٝ�gWP]�`���̆����U����;뼮�� ]�j�1�0=���'�F�A�+�BB�m��RՎ�\�2�����b���f���5`O�gn`��P�~�0wߍA�sJ�LĲ��
�^�ͬ�r���r2�1x���sx��Y��߬��3+�����p�m۹64�W�Qkn[���v�Μ,Ҙ�Gk�L�Fc�n�L�̳8�V�)�L��Cm�3iҥ�f��Z;��ǐHΗ-3ncc;�"]��;��Q��ru�{.둺�#�v }W�S�\�bk�[��n���gו��"�1i[�Fpw�`��i_NΔ3��N�Fw�P�X�ئ���A�S+��WE���75�K9�u��彦7����v�6��ˣ��$�]��$��/F�G��@؜�*�(��awewq*Ӹ�I�0�f�fV�����|�.(�v���=�C��6�̜V�Qqpe����P�n�,�ӎ�鋵�0�e��FK�'.?�(23lɰ�,��!������`5 e1o����e�h)O��ƞ�hs������9���׷�9v4d�*�K��v���U���c��X�6��7�>��Q���eA�KGWN�]HHG�l�>e<`���Lh<����J�2���+tT�ʚn�Ė٨+�U���0{-����3:�P��z�8��w+�}3h�s3 
��ەΘ��ˡ�1���WS�iB�e�t[�Yj�h��a�]v��u5۹�P��m��+WI��G��_�Sb�pf�����J8�u���ܝ��J�L�l���#]$=�=:Շ��_!,��&d7��Wqv9ui"�g+�+�х�5hi�.�3�1�k5`x�[��@��.��5��3�uqTI�Ԑ��7��ޣv���ˏ-��-kK����涬�;b��1eV��Ѩ��r�WbG;|����f���/Z)�6�e��{߽g7l�/	^06��ևo�P#��x��X@��Z��ju���E�Bɽ��Q��S��9���	�Y2�����n�n���7M�ƃ��X��w��l;ºf�s��v���=��[x�B���r�Ʊ�6}��w{���D�G]C�=��r'�H��Y�P���k�p����A�b��S�/�v�Xf�s���%YW
�af7�<�����UDr���AsC��=�z$G)�Ar�QTU=J��ˊ�B��u(�l���QQ8��G$�rtJ����r*�0���N�9r�E=��*
�<�+��I��a�nW�®�y8jFar*��D��H �EQ$��w����y%�2��P�瓞BN(�:l�(�';�T�6���	��U��쫔|�(��{�|���rz%:p�f�8Q��aQe�Du�ܻ�s9ΒU�M��J��/B����W	ްt�kT)$�9E{����
�J� �sϞ�����P�]΄�+D.sB�̪�t�P��ZUPUp�
CJ�ZR������LN�޸_^�J�D}w��}��&oji|��Т�Z�fW`�rJ�(ԹҦMSw������q������������udSk����N�{q_��G��<��2������W�'h&=Z�*��&)1��G�TE�x���kHs��˯e�]�T�fy�6j��O_��ɡƺ�e��y��ώ�ܹ+�6pVx��U������h�����P�������[�w�Az<�k�5����7��0�ĕ��gn�;��1�ŀ�bs��*�ŧ����K#�3Y8U�ZB�T�\���Wu{����.Z
�ޱ���y����x�k���d�]%�Us�{�� ��\^��O�V%�|�Ƙ�����/6o;/��'^+]mCՕFzxסx�F��+l�=EN��^Z���ZףM���:����wq����1�P��]�|k�Vי��rW�7[I)�f��wC���h^��Q���ey����n%ۭjq��$�	�g.��{V�����'Cu��e�M5��4��G��1��ON�}[�ಀ�-���W(g�s�=&�6�\�7��[$\'�l�Gp$�aX^E�cA��݈�=���J��]��V}��C��xڱ�&R�F�z�D�o�]� s~�:�8Ex�V��Ǘ}���,���b����'1�	�Ez5@��*�5T��%�}�7��d�ܥ��El/\m\LC��_]��#���v����^���Ք�����js�2bjv�ש>{���o�������\���Ү��S�@�txc񔎧;z�ڕ����v������/g���%s5�ů9�ÝW���..7���mU炯��1��ԃߩ�ˆQt,4��vX&yl���X��g��]<�r��-�̀���-�Tjp��	�(�F�.�����u��ڲޯ��V����݄�,+�ۓ:�2�8P<��bj� ��W��x`8T��B܄k�}0�HJ޿d��Uj��pe�����:�̵�j*�9q�
�)d�m�L�b�k~4���K�����w%��K7bT�/G�x���J����*?Ui]�9O����K�/��S;f�9K=���j|���yA��ZC�L?794�]}a8��eזz�'�D:5���l��wj���ʣQ�/V۱��kk>�{-;��\ѮC�����e;���ɯ5ZH�]r�;pp�p���6p[���}�0�i+��k���N��q7R��0��cۺn����E�w�$v	;���S�g! ����ֈ9=���s���2+�N�\?����3}��_�Q�~��q'S�
�ՕO�մ���n�5��i��a�R�z�%DԼT=^��>�}]���/%.��~���};|'yt�LD݀���Իo_+����&s�{��5B%s�{�m�O�T�c���> �ޗ��	hau�^�-(��k�U^�}q����~&��[5�Y�Q^��� <xs�����w��d�9a����6��~�TU�vj2!�ȫ�[����{Y�b>��&OW���z���۟�N��ga�es���i�.���zU�����-</FѨq��E��MV���{��~��n�M��BNק}v��>�S�+6.�ʧ(�Ȩ�Zm��ċ���խ�]x�e�����_�P�÷�p�M��Wz��kf��PݏS���d�w>�f�=>o�$N�vx8��;��C}�#�x���ȫꮒ-u,_�%3��=�~��9�	xj7���S�wa���5�����;����m�j�Z	�d��HR���f��GΘ��⡨�,����ų�y܉θ���l��8 =�$C-�%�����N�Z+ubd��9]�"���՚������#�����{������Wًe?@�^���?����7�u����`�u]$Z�!�q�t��ԁ��~�B���F�����)�����3��1G�.����:��s�$
T'�����~��w�x��j)l��/ۗ��W=��W�"���t*����2O�H����*��� ���5"���:�3<�w����\m�,�5r��AU�^�^;���f��1�p����~������yV%���GI�9�;��=;}�^�Pm",��]E\mm�����p��8}����� J��
g8�)`�.L�^��+�L�'W����k0�꜆�~˾BW�nZ5�������,t�ip=K]��Ǻ_�	E�Shj�99{w�g{<GgS�m�~�\�~dn�_�Xο�HE����*��ʦy� �AC�o.���>�P%J]2%��=�ʏ{��OC�����uQnU� ��䋫�FS�Z+K�����vxPX�����O6�g��a\?ER7*q�4���3/'-����Zf�@���2.2gx�d��h6Tk��-S�9�ֆ?Wb��_-��jk�gf�qz�#~�q1��m֞	7�\��u��5֎��q5a��⶗'���B8�T`7sن�*��^�XXڊ۝j� ��,Wrt��N�%-�۬6���9��Xo�Њzv^�5٩힣�.Tk��zz�Wj�HS':K��Ҁ+��y��IN,��>��{�
����zX��2vw�̔��EF��s��,p��ی hQ�:�=*mо��3�ܞ�]�u����t΀���懮u� ^]>3�R�3r���H�I~�8��^̆e`�S�(vx���V����=E��#��}��T=q���0e	���+�MM�EuS�����ܕ[n7�]k7
g��q����{,�J���M��D�2����v�Ǥm��>;�|�ʖ�ʫ������ݝ�L��ŗ<vo��w��V�H�KF�bP�G;@wl
�fc�����T�a�eU�1KӰ�B�'�/M#�����W LEwa7�dю�F��ݽ���g�'*�1���a�E����ջLx)���h�>�#2;����Ku���\���}�"O��ǈ(~��fJ��Y��/���{��'}f�0~�R���Df�tW����`=�]�^��V.ʑ5�ė�"&g�嬻�x��c߀��z�.w�������u�;ѽ�s���<n;j�*��Vj�r��U_����j��������?s�����L7��Wt"8ג���N=OU@�U-�a߮_%yO)(!�V��2Qݤ��r,��%\�� ����F����ԄY�uR��B��풯fD3U�/4�^N�Uk��h�sUsGmf�4�j��ʕ��t�ZH���uC�ݒb\���_W�༽ና��%��`J�p*6^t���9��k;.Q����m"E��ꈽ��fhM���W6nW���z�c��U��<�#jGz�i���9�i|��lv�0��9����kz�#F�U)��L=fB����ΔK���o�]ɟq� &��1��９�&��=�ֹ�'u�Z��x���Zޣj����cr%�uuxq~��b�Y��w���,5��.���p�c�[��a�^x����:����X�Y��ޣ�v��L���pǗ�8��,�+na?���\��+?.�Y~ڵS�����_�}::nܱ_l��7�@�� :�db�Θ�<�Ȍ}��/Y�~9-�U���w�`�s�b����{'ơ���^]%��LKf�;@=Ϻ�C��rY5��Jo/��(��>ԡ=�d�Vl�jg��]:T���GT_[ȑp��n|<'�(E��{�W_�h��C���xZ����%��Ac��;���[]F����w��7�S �G��D�s������5E���Jo� .��\LM�˭ >9�a����^�D3�ˎ�1�����f��b�t�ř���8�>B)J
̆�.�����*�厗W鮛]N�QVwd\�`������Q���u����|35^;Ì.M��<մy��73���򻶮���Y��,W��h�y�(E�.�<b�ν�	k�Ox���K�@�2,f�̓�+8d{�7\����nŤ�� +�����\�J��\q���#n���3.d�/Ǵ�/|�f��geld���-�F�߭�6}����U�Q�������t�u'����_u���O��zX���Ԭ�s]���q�&}��+��'�}���d� �4x?W������a���ǭ�Х'�������W�5��G���5��1��/Up/�]�9�t�ڶ��Wܰ����Ͻ���V�fm��5x�+�kȱ���t���`{�4��<�ʙ=v�Q�ɱ���t�6��x��`s�z���ʑ��r0��kn'����{%Q��=�\ �G�������k�`^H1ތsґY����,�!�{ݻlc�:����b���k�a�uHc�1��?L������QHL������(�>oL�S�<�|��C7�R�{$��9�����.+�3�1��rbl�͵1�3�ۑӜ�g[/�Պ�J].���5�d?Gz���"�Q9,9�Wh
��~"^]H�s�*��r�-9�:|:#fy϶l7��cu�9��.mT4.K1���Cr�W���U��2��i�N|�Xś4�e����.���^Ŕ�A��\�ݓ3�d��mC�>���E�Ȯߗ�F�ɻǹ�ڎ�ۤ�Q�F����,�;徦7n��c,���͵Jō2�#�*�ʣ]�p��z"@j�A�N�5�^>ޕ�
�C�Ž�������<����y���+w����dW�@�;�������l�����j����^�Z6㫮8\����x��D���U�3�{����?}U#N�`e�����^>��Ntsϻl��>�������{fs3Ѻ:�ˠ;��~2��� k�ι��˱�'�W�{����s#����R�>���r{��sܐ�ϼn�.H���D-�\e�__u�dF��/�K7�������$qT��]W������}@+��,��U�E���h�\�v�m%��m���ިj��U����ܟy���|2�hTul�)�=!t�*���� dG>�2@��A�j&j�=p�A������,�8�ϴ�r}s�����<���)QP�B�Rdwh~���5#u]�x�y���^�.�ԏ����I���F7}�zn#zt���UO�R�,�x�������}�-�2��J��=�(��i�gr'j;	�ʇ��Ux�x�;;,�U����q��)��dUR�̻�"｣�s���ez������➠����G���_�ǯ1����[��*�o�e��u;�rtk�ײ .�u�u��@.
�����켽�����9�b���m8P0*���~��l}p�5k�r�Qs���*�;��:������1�-ެ����떴i�����˛����fw���)�#�TǸ���D�gmΛ�9���9=��#���~��XO�a`��4�3�t��G��+�7�6_�~�({$%pk�G�����wo�7{*Qxp����x�u����Y��Y��E�W�V�k�����#�fZ72�y�!�����jX��I��R���D?W���b��-�L�4&dZ�ձe�;/��
���#	L�,ozh$\V��q�-S���Ύ��}O��xi��"Y���c0_Ft5B��K��5ݝ��%3���[s��k����x-�ُT�_�}C���^�xX莬�ᐧ(�y�x�no�`=�W4=s�ʭ��Ȳ����q����)T�D��_�=��g��{�k����ϼy�GA�?W[�\�<�d��|%3��]P��;���i#Ԧ���N�*�e��Tuϫ��=��o�x����d��t��>0t?lG���VO;�B��I������3�xq�]��@<����Um��ǜ�R��3Nk��q�%�%�kݮ{԰f�R���ǭU��eUΞ�Xʅ<O
�zi=!t�ʧ�W��'�M�y从�9%h�8�5�U�-�9�x�����.�b�r�v����bQ޻�=��:��ٻ�L����^e��J�n���65��[��oD:�f��(>�����]k��<�z'�[[�Nw+��ӹ�}>�G��A��k"C-�reh�،�>�2�,9��>�z:�XmRCQى��n�����U-�3���?�~�'�n���Tk����1���>ǫci��e�q�5z�<ޠ��\]{㻳�>ZG-��A��
��QN�A��s�~��������/��z��wLf\Bg:��07��۵�����G���m�xv�q�H��C�ӕ[\7#���~79>�c�����
w����-�a�Z��(^�W�ḱ�oO��r��y�c�f��Ǟ�~�����8?z�`�����hQ�^z��#,��G���P�������O+��o��8c�	���|�����jk��Cf��n_]�u~(g�;f��@�� ��O/��']��M���{'LW�8v��<o�ٱj5)���t��ϛ�����KK?�����5LMӮ����GϦNa��3g�w��+�2�B�,+{B�ܹ��Ϋ���D�)�'��{2ÿ�Ղ��L�s�L���Y���gy�Kﯝ����z29Ie\w�ȵ�`=��\�*#�� \d�s���g�xzg�G���[�A�}����+NC��7���)�,�y���K����w�7荾z(�F�/�l���RW4��*9v
P��5V�g<1\D5��n�Et6!U�Qak^oʊ�!�r�N+�:��~	gYi<~̱y�\�@�7��,Y{��qN�(�����������v���x����a�g�	��%��(=�%������-$�D[ݲ�˟<ݖ�K��v���Ğ�X2���;�̘�wv��5mف\a>��z��9���-k�;��۶�j\� �l���ٺ�K()�bgv��'N�	�sb��賕�փN�Nz7���_,FW
=SNY��=����T�ק�F�k���Q࡜�2�fT�eS�okB�T��;��(��$��v�'@>���5p)`�F�� 4�o۟]�A]s��ʔ����Of1�S͕ȹ�9���ju�	z��m���G��j�[@�٤�:C����5$����f�Y��:���E�4��ɺ�VX��w(�mӾ Vv�zi���7{�X�$MK��/���v�л-<7B�V����v=�C�2��"ܺ�����G؁yh�\k�z^��ͳ�`y�oel�yՇ�KD���ҵ��f��gvV2�Δ����8MF�9�������s��x�U9��6��7k����Ƅd�o<�}���oYֻ^�t`�UcB�va�0w�s5fZ_�1�4REp��x�wD+39�3�l����d��u���m�r����+PL	�گ�NUDۤ�����jx��@���7�ήV�oi\��gg����Sᣡ�rf�{L �܈�'e������B%��ށ�\�+��EԠ�i*hӏv�ܔ����J}x҃wh�h��v��uf�T�L��"���nJT��S������b��(a�S2���L���t���2�V���潻��a���gX��5�}4\.Tkm �b��\�y�-����lM���a�Ve�L��+3����us���T�w�� ���!��8��d�|����p��W.�ø��N=�%�u�X�ќ�D�*j]�wl���� �o��D�����U�v��.��̤3J���G*��L�2V��c��\1Wv�ڄ3ƕ�n��ѩ��c5s���,@���E�ZBUmo�G�n�ul�Z�����CF�WՎ�j��(��I0�۩�
h��Dr���]�j����eH�ǵ)j���oI���d>�r���3����Tۢ9�k��/F=͞v�%�uj���sy�Ǜ��os5�9�,��X��#y|�q&���G\ �IK�ѶsZr}p����������kId�%��o:��3�X�l;y ���1d
b�N�_�{hX�c��{�N�{�a��'���R�(!�����>��`ʉk�M�#�#9c.�S�H�s1��B���Hĥ	�ک1��k6��x��=-7�5��-=�6�`��R�w�[��f�gD�̔)���R��Z�V��� T��N��W]ݵ��rAM_�Ɲ��ܤBd ��eq9A����α�P[��t�2�Ft</�i����C�t/��,�$�WG�+H����U�as�t.�Yr/U=���*&P�y��������p��<���=Ź:�V�,"���B(�9�#�AE�͑�`$QjC���8���s�\�O���(SԂ�(.ˑ�J���z�M�B.;�ʊ�Dwwl�s*,��P���j��T�ZK��:��U�'Qѩ�	¨Ԣ(��(��<�{9E=�]�\��.��NϘDUE��!� �dU�z�"M:Hz9��WC�/=�N�^�r�LH*�.Q&q2��Ѕy�$�r�T�i2��$�r��Iwv��Hwfg���p�Μ���*��Q:��\�&�3���8s ��.��	S�!����s'6nE7�ȝj��<��Y<�֐�J2}������jN�sa��`��{dV��6s�j&���_N�y];&վk��� ��Tn��""�p�7��o�|lO�g������5V鋏-���8v_\vI^��Ǿ0[=�Tv�z
��^{���Z�TNWh�2���up��l�����i�.�*o��#�/��H�}]7�ݎ�W��k+ӇT�R�L�LN���{*Ǡ�}�	c�v�1q>�f�O��N�����W�7w��G��W��T�;��.DJV[��@���\Lmf?ea�%���Ç>��~��*���D�tR�w�����t��s�t� +]�����*�+����v��̹�H�ӐKºM@�<���s^�3[�:OG�5_� ����ԁ��L�+�����g������i�3,�F�7 ��3�b�cOi޻����>�P�u�=0�	��u\;�Q���Y��'�;3��z28�X����
+���6�T0�8}�|�GA����8t)�TF:��q��co��G��H��;k�g���Z�%�J*�#]>��w������5�y���i�0�V��<b�Ov�-��o:� zg���g��ן��5����s��,��l5�~{6���[�=�< �k�'���ϼ� �Q�U}T�ާ�z�0��Wn�3h���AF�np�ײ�J�����3m���	�ʅ�U7����;ڔe�٧�9��6y���j�K�SA��
���J2�O���+��{�0�Q�i�<�!��8�ʾ},͕ut�w,��k�C5Ĕ+�q\�#��/���q������Yr�vg�X_���\�_1�J��=/�W�"-�&�9V�~S���&n6g���s\�n�owؗ���腮�L������lod�*;ޢ�s^*�K���5��c�T�ܾ��^灔�J�S�d5k�rr���/��U^}g���)�����Wx��(=��3~7|����nU�z��S���^���c���x�y��R�h\�a?��+���`������yv�ޥ6��=j���U� \e�fo%���ɱ��j��s��l�;��'sM���uc�{;q�e��jQ*�B���q����-��_���X�;������Ǖ�=v���u��W�Ŀ{��ۖ��!��F��d�z���mw��O�"=P����7q�\�������.�zw��D���8;��*-�9!t�,a���*@��X/��s�y��F��cׯ��<k|����/T;�[wF'U>�}�D	��	@l�⽷@o��j}}>�:�;��9�����;�R&F�R���J��;`vP�H�O#�Q 7���Je��������ߪ�7��a�Oqҡ<����f��{�'���w���.$���m
�d��gJ1�Ol޽�S7�yGW����Sp��L\r���Rˎ��Y헭W]�b�~�hW7��v��lq������ԭ�=��+?������t���l��O�U�p�D)�X�R:����h���� �)��1J�3���W%���%N�M�/\�x�g�]��΃5�8T+��)�Ȩ�\OyTg�L��j);�ښ��!�l���ԉ������n;�әP�=�^7���m0��L��=Ƅ�����smX�;��:#���|�+h�4=Ͻ7Zw�>��mH��^�w�NO�X鸞><�P0ҹ��{r�]�����	�3�s�O�w����"@��b�ʿ-my�N�Ξ�zʣ��B�����;��LtoH�N�oT
Z�t�纽�ߗm�>Ke|��}���]�u��>V����ru�d\dϙ�ɖ�i!����%�N�6�6���y�����eJW��{Z�=�{If�s�VD[��"�e3y2��ڰٽsb�;i����1�1!��:ok+��_���1��6��s�՛s�PmU]��,�l��s�޺H�W��{\Nı=�U	�K�����r�49��
r�/���t���Юhz��~��o�n�W�����^�,���ÍS��sL�����
��G�T�S�3cQ$y
n�>������3|W],�����2�opѡa/'Z.dVݱ3s{ۯaT7 ���T�+�p�=�e>�%�/�uu��ݜ%wT5��pΓ9��y��A��/{Y�����=�����x��e����>n�{Yt��_�V�q�-����W����=E��!��D�:����p��$-sEo�w?_~\�x�oA�2hOG�Q��ިW�zo�i(���.�3�ȫuNJ`�*=1(=�%R��&H���J�9kެ:�w��1�v�u�L��ŗ<vSs�s��2��t�od#!��P�{�(;G�b|�z�
�~��c��X�/WI�x�4zB齩�����w��c/԰W�Vlj���O~���k�$�g���i5�]�E���F��K�M�kK�R7�}�7�u�MPZp��
�}r&����3C��J�������ߘ�׿�� k|R�p��T{v������-��7�=�����C��ȗ�:^���k��e`xrrf-rM���c�|,̸‘�W|@�y�7�^q���q�����Ρ(z�:��y	Oz���eMU]W�I�x�O�莟
��#�p	z�@'���U7ӑso��1|�+t�� jc0��ݕ��mE��4�����}W����dojG{e�='u�m��/9�p��,��͂<|�"���-�֊Ys�)-���*ޤg-/ ]B3Qs�nm�ǹ4����L��|����꽾��2Co6y�R�k����ۀ H�ţ�9m�ea�n��_V �z��+��&��;]۾n�gN*&�4���5���*�k�ﻼ+t�9������O�.��L����w�!�oM}��bV`s�޿3��q���:����;�ݾf�(.�L��*p2��� ���}e3y3�q͙aϼ/ֆ���슮�禕N��V���lp�X=ޢ���)�t�{9
� ��~����������oJ�c<;F��+�j����aQ��9՝t*�[-������Wt=7�;�G2F�9��m��:6m�d�VT��3}/Ž��O��;�u<`�{��BKG�M��K)
�`e��U]�:Bp�)}�Z��iЏN�*!��~�����vzj\�z{3�Uⶉ�ހ��Ӑ`���˺/��x0�}�}X�;���O3��ԇ�Չ���Cs���]��U�q��s>$ޝ��Ǫ3������&�x7��OA깺���e������g�� )�݆�!��OMX\T�9]��5�/Ǵ�y������[|��7 ��:4it��ڮ�:�� �s�&�����k>�^ގ�*�nz'�a�������̠�n�D�Su~k9j��-���`skG��K"y���;nj�:N��@ǫ;�L' �v�71�u{X�W��Wr�W2TD33r���Y|�ޝ�{/������v�<ĝ��:� �w�$����WZ��;��tb"��"��a[��>��<��<��d��<�1��=1O�O�;�������~��vo���U�]~��m�Q�خ����������3Q�`N�\p���P+q鿻��j㟯T��:X����c��v��A�� ~����T�k�\�M����s�f�i�����W�,�O�mx�;�N�m�#*8.B��w�Ʈ�kO�JA���X���5�M�_���3]۞�O��1~��r�UO,Ô<�x���+�t7X6�������Ȟ�9�$e|�{�W�>��p*�kM�%��렒�U��gj�&<�K3nxy������B��!����U`�Ʋ+ʨ�ޛ���Q�w9=������>��2�޻�'*�}n_u�����<Vv����a�s����Dꮭj�^�ȟ-��%ϗ��>��#��7&Z?�6l7q��*1�����T;��v�1��Fo�p�I���Ú�q�u�֋<�����^���.W��J3Ճ�h���{N�Gm����Q�ܼ��_j�s%�Ȝ�/��=Q����ze@��wC��_��.Z3y<��+t�sӺO�Р�G���I�V�[ә�r�Ѫr���"]$p���C�?���itNv�*�S�t�c�bw�eL�"�^�y������.u�Ѡr��H_2�]��m�JV�2��%�;�ո����;���t�k�݋�s���sg:�B�n!����Ed�u��-����w����_]��P��2�~�U���34� ���|���1��>w�\�*}y��Y~�%���>i;#���-̹#���b����T�����x<z&j�������-��{kڎ��R6K���K�_vY�H��Q�\v�V�z�X�k|������+��/hмR��@<2���;=*b���zx:t:��y.�=S)��f~��ɞ������۽��pl�gS���SD�P�uE|�B�SC���|6�:޿u߳��ꛞ�O|�	��!)��Tv(����<�����k�j=LpUS���A�#V����2�:`5^I#�7����m�5y^���� G��y�X�5ɽ�����J [9�Ew�k����_�/Fjvl�h荙�q���+�n#�Ղ�����ð�jFw�n9z}^���F�����U��$=� �<�Z�+�����;S����^��<�7���8�//G�8������?�8���؟�����'��#�tٮ�i{�"Qx���}q�޹F��<`{��]_�?�t^�ή��Z�K^�ҵ7��+ʈ���9NSv>x*�$��YS�?lP�W�=Z���T�A/Q���M����V
Uԯ�F4[܌�q��oۓ���¦`X
}��Y��ʏ[�X�E+��V��bu�q������gz鴌��g�L�V��<�}�def��"�2g�o&y�l�{{\,/5LJ���*y����*��6'��K^���ݢ�˝��@U�~20�����6�6n5͌햏�{�z�i�3$��{'��O��n�c���TK�܅W�;��d�o&Xh�m�����7�jϘ������W;�g�z�k���h�]\.%VYex����H�Au���O�k����$��%����C����ء���߷�_����h�
��lV}=]%�I�>��G]P��Mt]��Y�)*{��*�z��g��Oi�����<;��7�<{>���2�Ƅ�.���ѵ���7�{'�\���]*�7�X��t�}���ݭs>�1<vo�Nz�ʂswag{*�i��������)��U�H�%i�S��U�ُ�To�s�v�<O�(����W�G8��k����Ӓ��+���E���Q<�}=Wp��1��zMx���c�H,:��cIU~�:��gx�н {mMP�9������ț�t8��4;DJ���zNǋ�3�a2"b��{1�{ۅ;����U-������k��v� �zl�3�Hc��k�&��JCx`�iz#�c����A�"�n�+֊LU�q��h�4=�l�:��.��]:]�9��IX�Y�ك�(���7i`Ւ��/��2���j�݁ ��'/Q�����z��p�@<i�S&���B���BK������vi{��w^�K�~Zo��8��x�'i�u�8���Q�q�U�W޼�=;>u	C��I�TOM{׃DG^55z��匿ȼ��W��ӿi`J�p+g���S�J��������R �>��<Rw�2� �~�A�n�-��O��l��1�Ԏ�����'u�m��O��=�'i�~����e���T��xQ��������^&�����*g�s�	��z����~qU}K����2�v�{D������{��R;hS�͆V�\`�7��S6O�kVl����{��ޏ+��C���Fk��⽑�mVoz�+�@�����W8}���&���g:o�����x��ӛs�]�7���9���:ξ
r�;�t�}.�{U��e��1��J��Uy��]��'����E���[*�Ձڝ���oO�f_\v@�S��_��i`�ݸ��c��u3�.�{�e�㎐���e_ٵ���=�E��t��~�8�Rz_^ʏ_�������B[͠w֔���(�'1/a����2�Y�#�d³u4����u�5`��U��T�X�"/-����d�}�����P���4��WC��l���an�0�L�{D^�˥OAz8�|����ƭ���z�hB�z&�f60�}���=wC���׃KG��:�wK�k��_��Qw�w�з��ZG��H5pE9f�g��{��2���ǫ1�+�f��xZl�ٛY�rr�/T�A��3�����M��� ���[���Qe_���۠:��˙6���R"z%/{azW��^��z@�=��Q�ӔioP��ޠ:�e �zL��(ZM��/X�^��'�3�n�~�l��U�W	�C�g��Ô���d���'���u\:H���R̋ʿ�H�=k�ݜ������ER�7"}^�Y��zo�ޝ},����A����o�U��S�*�}��n9Qr�{�;��&��DI�}p�n;�ӚXQ�Mx��y������@޹�=5۽�&������߇���x��Q��Ճ�	�;?�a���n'z�����Y� glF� =�|a"o�3��綊Ve0+6o���}
l=+{ƐP�N�\:�cK�/��{�W�>�v�6+�M�_{�j��=�	��fxz�at�f�p�9�v�B�z�5��!��5��Vu߀q4�[���$ñ�yl�m�������F�h�h���܇7{
`���}�.�
�;����zU��Ҥ.Ѣ��~�]Fˑj�X8EXP�`{��\+��#w&v��P�a<%�Ίvu)���j��VE��X�"v�݈�� �t����/\�T�쨜LY���炚o&>��Ip5yMޮ�sV�qި��ٿ+�`���S�q��3�+}Z�\�k:=Wϭ���R��k�n����=z��Z �SWa;;N9�#Z����2SW]ɩ�$��ر��y�u=٣r@��Zd[���Lv�+4��:���m���;�{�����6��9ڈ<̘lG���Vv;��NG�;�r�YxB���-��`�GX��ꣽ����Ȇ̷p���q�X~b�I��gR������M`���vZa6	�Yi~{��2:s���t��H��e�wnoBz�'�+�K���1�����V�b�l�/f�������6�����������T��ktw�N%��}�f� ��_y�o�˝\l:���+��%�H����CG��Gr�Q�o�iJ�On.�Y�x�yOH���b�<
���3ί0��4�y��hȏB�	�L[z�h�.������s���+Ɋ�΅�yKw�mt/qr�c�c(���EAP3�Ε,�Ԑ��ռ����-@�ξ�|7�WZQ����*���1T��wJ��O�#{�5������J�aҘ�� �2�ч:�h���B�v�ɂ�
�% gX��V��Գ���r���5,�;�/��M|^���ф�bI�F�v��3H�K�"������"8�pi�yc�u�^e�)�t�I W,&�.�T�KǶW@��h�tm�c�����<NP��Z�EH����p��x��]����·�j�n :�4��t.��+;E��J�o[ �_�:�?bLE�|^c�|���ʚz�&H�BI+z�<�e+�J@G�t4��7��P���{ր2�+��K�vl�B�Ҽ!֙Y*K�^�܇�j�#��u������6����x�7E����x+������9��R�FKI���0rθ��с�h˝yDc=�q�]� ��NB*�j��� �O�aj�t]� Uv.�2�.{�JJﯷ�[D�8l��Xu12����wu�ȅ�a,��ٷ�]P��|!��}�����I���Duf�ц�C�����y��:���L바��!W��;�r#l�5C�\}pW�V��ܢ�)\G��.�� �������f�}�|웫(6�ȥCGk� z��4��J�p��q���F$�
k�u�!�{M�4i`ہC������Ʌ��n#D�I��w�=��\��m��;�8OVnYK�i*����v�̂�p�j���Y��R�����8��]یj�;�VaW����e�3�J��D�h��c��.��6������ s���wp��J�Z�7Y{�����YIϮ��(���UPE�䎂T���{���rv�nH��E����L���2�{���A��547��ʨ�%�Ή�OWCW%�#$�OD'
����Քw]�D�3-j=s�O����.]�¨��������{w,�(S���w�גuwGT$�.N��NUs�AK;�w7�p�G�q긢�De�V��{�ϼ�V�9������>>y��<��i��9I�R��Qy�qFR�Fw�N{�z����H��W9�*��՝D*�41k�<q9���!Y�p�8�"�\uū��E)�9�S�nw�g޸N&c�^�f���L�W2r��>��G�,��;�.�Qh��!���Ԕ�����Na�Yi�>N�p�.��<��ክT2��j."�ەV_G;���xu't,��*Ǹ;�+y��1��'sK����Huo3����+3i�E�#Ot=�z�#�Hy�<�䫓��E�8�]4K�w$�p�H���R���P$�D"��ԧ�>�+o3[������Л����2��$���o��[����V�])���وe(����N�i��f���Z�G6�tH�����W�i�i���]��y9Ts�n�}�q��?	�=�L��l��h%���_��*��e?y8�2��4_m1b�1��N^�6�;��9�N���]�5��3��WY��� ��Q{O�����U��c���T�ƹ�wˏ/Uў�/�9�Wo�BTȮ͵��D�����E�R��誑��T��7�����,y�v5�f&�$��\u���;�GY���D`��wB�����!�Q��ϣ�h{g��mNW{ǨO���V��/�j23��,��{�Tu�������v�N���3����d�U�<X�0u�\F]��9�ֲ�^�2p�No��{��9�>%᯷���}T��K���K�w]�u]$Z�!��&�3hj�ɩ���og��9���c�Q�y�Z7 1H�y�Ԧ,�P]9�������~�>�wI��$��nf�G{��4v}���5�>W\=P��a��B�����W��*��*�;fP��n=u v�&�Sr9N�U]�{"��0��z�N������J�j�C��S�~�f��38��5nZ�I�����C��˕u�r��Qy�/�^J{�1!�]A`��� ���l��ӭ������*T��u*j�m��)8��ܤi��Me\ه��h���}i��|,noV6/�����,��:��	;PC!��I0{��ϫI��k�����̉�:(��~�k�����{�=�LB�b�:U7�~�O®Fv=�� ̯V�'�ث���s�}�X.9����x�ّ~���Gz��@�N�6�D�S�Ѭ�K�<��P3˨	�t�'\5���V��eL��z ���b��9���U�Sh���o�?�W��*��U+9�P���҂��k�FE����F��Q�ٳ����W���)�-�pڢ.ԫ2;��7�L�/>ِ����b�T�˔Ɍ��1bs�W�)��p�Ό���a�Obe��s����n���ɔ���a�u��^R�]�gO
��8�$�����\:��HpFè{�)�˖܅W���X�d�o&Xh���OJ�U�>�X{p:���Z��r;m�Y���^G����e��s�sC���J�{�^�t�7;嚨oL��zc����#�#_}�/Ǒ�p����<\��6|%�����55����-pn+�_C�~�@9Ǆ�Oi��z�\O����J+��<]�vY�\�+�3*��WE֙�ֽ�c ��Y,d�	��]» �6v�2r�c���Z��'�А�fN�G..E负�%[���e��qC�+ymnP桳����{�}�!nP�����o����<Ѵt�9���x]bqw ��>Z!�:}C{��kW�.�_[;�չ������~��~��v��/��ܬ9���nΎ�U�S�٨)� �/u�}{On�X���}d�*6
F��N�Y�<+1����xn��X�x�^�F��䋛����)�s�S�+�����|nĪ��������1�s�W����c���t-�/P�#�1I���ڪGq���X��M}]�	P$u��*ǽ]%W�uNygU�mj����3ѵf�]�
d���㯪�:MG,5"j9����V�c����q/����6ƞ���U�x�Ff�Ł����2������h{���N��nߨA�Jn��֢���G��WD:V���X�O��X�y��x^t;W���LT��#�Tm{�.:0nd�i����^VeT�9���[��,�ߝ�ޚ��cޝ��@��#�m0�w\%�y��ܙ�ބ�������mw-PW�9�]���_�*��5��ˡ����t���e{=Jڝ�6:X�/*�ó1IS�F���T�R��ػm�27�i�"\��s����q�Tc~ț�2��Ԟم&��c�49�SN�B��]���cm����۶,��]t��7�ȡ����ߓ:�1K�U�O�ˡ�6$[��:.�Dң�O2�ۨ��j���[:�$ʕǒǚg7؎۾�8z�LޮJh㝺��a$>�1�����k����d����]�3��ƺ�K�2��n��ub�
�����d[ �*��8ϣϣ���+Ci��Xiet����#��m�7q����i|{�:ξ�(��r�K�s�7�0'/*�=^Fv&�θ>�o����ľ����;�d�U��z�t��R���O�_WTtUw�@��}oxm�:���by�tl�闦È8�	��e\fևs=�E��t��S
�����q��]�s<Ev��D��������7��%��]���%�O� ��;������ȹ�����~z�|v|��y�v{�n������ .����SK���=�7�/ײ�Ĭ�QW<�����؍1q�(�s����p\>��m�<��*���;�����lw��W��˷�9��O}��+N�T�>ޣF�t���ʺ��(
�w]&m](tJ��A��������]�������O3Q�~&O��
�Q	UOL_A�5���d@~�:W�RK�Y�b�{sհs���<r������a��X�w��;����,c�]��
!Hu�q��\8Q���{�ͫ����/_4��C�FJ�+�nG�G�J�P�eQ�dw�,z�~�냮�)b�x�cj�|�)�`��,U��~�"}��I�Z��]�3.���W[IU�jp��x��������y����m�H $F̒��!����u�\1��%B�.�>�����&��Ĺ��j;4��>eY��/�T�~}��7~Q��s�'�yzUҍi_h���������;�¬���5톱_����� �H�{)@z��7^�e'����ʀ�Jm������͏Q߽�5��������W��י��%ɟ�'�`.��w|%.�KL�O�>��2Ǯ7�	�N�3�[\<�wk��J5ب��ׇ�Y[[{o�fi��4��d{+���ȫ�&|�0�\V��F��C��E[���u�����<Tm_7�'�	�0�{uL�ƕZ�zz{)��WxC�~"�q/&Z=��s�bÈnw'+L�k,�K��ONO��N8y�Ή�uLƨ.H^��WxE�?/.W��K�ɱ��j��xתv�vTM��{����a��Dz���ᐧ�y2���UH������8x5å���jqv�^�X]sK�fԺ���������j:��n@�N�\�W��{0U�r���>�3qImb�>隗^�H׽0�'�����;p����vY�\��]G�0S>���F�@��J�*�������=Ѭ�-�2�n�i` ��ke��/ɻ��Hg/؈���z���-$�f�&-�=��Mtx�ga��P9��Uk�^շ��9��ۑ4=�0�u�K}Q���W���6oK3Plh�	Wlv[x�]�/�]�	�+�₲3���v߆d�� ;>�ڎ��U#K���:��*"���H����Oя�!��aD��s��{���Vԁ��Th\c�Ӹ�P�L:��S�.�U=�yM�ȫ�o&���+�5<�~xH�m.�o���n�׋��<�u^�T)�X�������1��DƬ����p��J�{���
��5!�H�.V�̅�����{%��{��k����M����������>"�i��T=�|<���#2�����~�k�
��k�f#�\-\�WB����x���{��OF� Oʕ1p�s���*`���>��`�}�G}3�nmH�K6��J����̰�w\Yӝ��^>S�z���	�t�'\5��YZ*���7��F��YC��S�#VE��Qy�>�����U�ɟ9�21�ƙ��s�鐇b��;��6��1�mW�
����ٚR����������١�ɟ3��-l�{{\,Rj��߼|�([��0��O=�9���,�z��=���(�ǱT�˜e�u�V����S;�L��f�g�z���P!ڭ^e㮱Qvl��F�机̠j��"��Wgd�VU��d 9Y���0%e����L��b��fm2�v���]0h7�s�Џ�p�\��,��k�[Q7Y�q<�˻�hN�{��Gy�C���p�hδR��+e�2r�e/N�מ����G}i�q���N�q��B��Xڪ� Wgz���%3;�[Q#	S�����{��<������X��;o������Y������ȅsC�;ۯ�ީ���^	z�5nY��ѷO��Ԭܨk�"�^�g#�O�E��ceu�@���y��5
��Rr�ܒ�he�xo��P���P�����酽[|�v��y'��yd\�����G�=�'�f�����U�'B0wOzbP{�z�Tvu�`�àX����>�1e�����Y�D�ʔ����z�����_M9 \*���Ǯ���~��c�ӹP�]'��J%���vg�34�-{����#�*�̀*��K�~�)&�}���&�O��#��<8SO�\�UTN�p+m,�vP�+�M���fGq��@�}d]�S��\���rW�p��q�*M�����otvI��f�Q��+��%U<o�����Z*ګ�ԉ��C��%�V������:7�����_��O��q<ɓ�����m�{���mW�weX؈=f~ܭ��j7�M�����ٍ�����O*ʱ����a�c��SD�`�/��L#��.���,bLg<���{��U�j��c���Cn<��[��K���+���\�:l����jmb�F�%�����_,�V7��0�o 壝8�JX��&��gf7�ŕ*p<Y�3�9e�x����h�Fr��=�>�i�O�x�y��M����N�dΘ�V�IR��_���p8bF+����S��b�W+��_����ș���^b�eVy��kC�l���M'�훊퉫	v�Q�����+�su����0N��� �!���O�.��ϸ���z���̸��FM\�K]gPC���F$��ʞ�����c��xJ
���������Q��"_v��~7ф{�kMi�G���>ٖ�k��eyE�c�M����QegmN�`=�{��=+��UQ�z�{ӌ_H�>�@�k�p�/�}�0�ƻXo�/�G���n"WW�Ye�W5�"�ӕe</0)����*�e}>V��ɴxM�U��~ڝ�
}3�y�j���L��P��9W�f~�tR�Y=T|��	X�puk׉�g3�6Gd��=�x�����r\!c'�����?�j{�mH�y��#G3a�\�|`���˺.:�׃KG��	c�7��4hfՋ��d���GD��7��������z�3pI�+� .��񬧩y�C�G���ថ_�Ic��f��F��� ��ET�w%'���;��Uo�S	�7��;D
�s>cJ��CH�L�鳞� �+_tKsD�(�[ZĮ�ܖso��5¹�G٠��}�5����8�}����V��;��\����՞)V��+�|_�³А��H�x9ߔ� �w�
���rʨ������J��3ӣ_Z�s��sW2k���=��	��&NB�q�]@~7�{��`�ٍ��1D�������_���^�C�'�c����c߆�	�Jd���'���p����˻÷sS�G�7<���xظ��T��g���W�{=>����3^���\p���P#,�*ب6��Sg��1~Y���vm�5?4��gh����N�v��a}�Mx���K�zW	*�쭥��l���y^��ݩ=�6=&���X/��o�D�>�[u���^k;C��]XH���z���	�����=P�0���N�K�u�h�C���5�=EY�]�ؾ�pZY��'Ż���Ϗ�S����p7�<=� &u�t뇙��x�a�{2HH:y�R��Yyn����q9�-�`�~Ȭ'�1d��ze�{z�\NUeq�U����ݦx�4���B8�,��Ü�L�K�a�+��)���'b�e��6��b�F7[�}�I��kQU8�UMmݔ{��wi#�ʇAb��Ot��v�u �j�'D,\" T.�ӝ��5A������{M�n}|�Q�e�ܵ��z<�|��"jV���s91�`�f�|��.��&၊���n��z��%-�'�t�p)Oz�z��;�<cr;��͖�������r���Vzls!f����b�N,�F�ݝ���P��y�2~���¨��!���p;q]����(�g+�rf�`�oӋ.1�t,�t�]�lp���7�s��Gm��Q�n����d77��@׳��4<�~��r��(m�:qo�U����'O�#��^�C��V�Q�ޝC��u��\��'��<,ԝ��/N��k!�7��Zu���<�aωxk{j:�'�H���7/�q�de ��n���g+��}�#�������������h\F9�;����n�=z��
w�g����}u7:�{����^�$
���D�Rވ������5s��mp�|��b��ګx�C��F�}��V�3�z9�G�n%M�. ���5"���;�Uw�>�x��z�N���bؘ1ؽ�̭���3;���ʩ����#��u��9�lMw3d]��}qշ�O���'�����S
�>��yhQ����;7��
��\)��/ʘ<n;r�F���`�熧O�"z�^3^��k�E=F����ͧ��z{�A�Yڶq��c�����b�ԫU����o35�!qݩ�Z�L�:����3��U8WV�1lU�7��T�������m��څ�U��k��re� pGc���g"$^��������
f�W�+���M�a�!H�	^@�=���M��Ѐ
���1��9�e�;8�ȸ"�Vf�4r�3c6S��:���mO�m�Em�:*��El����Sv�]7�ZIJ{���`�aʘ�7�.8�[���T"��Zq��Y>�6���Yfv|��HL�r��i�]M`[N�;b͎Һ����wd�k��(��@�B��"�v|�x�޽I�9�5ݫw��(/3�)H�(�٪�����F^�b����X\�r{������4�;����MRm�yǚ�Z�[�wVw'���҇EIs��m#'�7@�Z]���x�}��^�����)p�����J˷�aB�n]�[9Q���I�S��#��}�{�F��G|wazri��2g�Xa�G��7(����]s�Y]�� h�U�(�!h�u�\*�݈��8���-�;��f�FIX"r��v�s��ۚ�
��8_Th����DhAK�uycKl�[t��k�ٰ��[�N��$�Z梠�t�3���w�����	Ư�\�}Gr����x��V��4hc�(�gѵ\�m>��r��8��K�E� ��,Xs5'�K�Q�nm��U����!0�r`�t�v�.��ts���LӍR��mP
f�\n�|ԭ��V��� �cl�{[�,H�h�,Yٹ��kd�J�5cv��E�[Ui�u.7%�6s���8s�6pޭ�Zf}r�6�a��k
��=.^{Z�����D�I�{)�:��@ù������EB,Ս�n�oJ�p��/���`�t�V�[�eǨn��Jrܼλ��z�6�ۡR��r���M8�VƵ��Q��Y�r���ݽs0:��4�L":��#r����T/�4��o*��3[��B����p��qȻ2�sE� L��v��2V=�y��L�z��X_V�k��|�
Z"��a�7j�x�Y�H�1rv�T��ܶt4DӘU_v���d�֭v�q�#ID�<�ηή�V�[����E.�56��:n#ڛ��%v��k``����6�/�,y;�]��m�,Z�
�v5B�U���J�6��.Ž��*|�����b����A���z���rL��u�n]�`������+Y�������Kw�{�9Ѧ�k5ٲ��T�u��t��,��ܦ���+k.7sp:�Z�fƲ���v�c�I�G��̦��51��|���;nl�s��h��j�;X��N�V��`��V�BUjI/��*�L� ^�׷wi��)�(�Lu$21Wq�nN���wEϽR9��.Q���Iw3K�Ô��U<ɏ{��iȰ���8F{�;]��$*u;�i������uuq��T�'R��� .DnN��B��p�eH�΅Q���+��"�Eh�ҝ�Y���QT�z�/s
r�w\*2N��5 �J��TՔYV)H�䓝n������C:q$��%�:/>�
��={����
%Rr��u���L�w�Q�wn.��rK:�dx�҉:W��G�.HS��;���p�s3�QCS�C������ù3�{�s)0�*9�AWϽ��y:��O*zzw�c������E#	κ���n|�Qz�G�<r1:�NVs���r�p�Q�*"����s�^�n9�C��YE�p�t/+
z�z��y�h���;�Dn�TD��UK�n�/]�f�[�Wy��J�N�da|�O>8��r�w9:�UMO����S#�(�s�}�������B���;��U��;)����A��]�vU���r�8x$��cH��\�V"#rD��6W1̳��t�l��Ʊ_�l�B���;�d<�=>�Mǋ��7���Bt���#!:�snXۇ��(����B��7���/6<CG�)�x%���9��K?*�g��)ZP���҂�^���_���w�� ��Y�����޹f��|Kg"'�^g�vF?K�Cѓ>f�&y�l�{{\,ug��)�K���eN�<�Jc��'�+<Wb���:cW����-�;�h����FL�o&X\�u,�R��T;�=�6*#7k��}}O��e!����)�e����� Wgz��b�����35�qֱ�9�^ٝ=�=�<;�Dm���F�\�[��lh���ᒫ,�� ���� ���W��,$<��ʂ�uf�]��[�@�ɾ雌�mM�f�C��RG���\v��Li쮢�h8��uT�NV��nUϼ�Nq�@�}�ꇶ]`���^����~<;���~�����=*��X�&.x��S%�M��p����˰6�:�0g�/zc�gGlϩLSQ@���O����o�g}�{MO/Jge��[�� \*Ѹ�C�"=v�Fc���s�w��>�����D��;[��طmAq3��AV{aZ��Z\y�pE)umY���Y+��/�<3U�{Z�E�1:�d�>}Q�+���9uɦ*���ju��1X�	Hou����06���زNT%o�%Ki֗r����\+Ut�T/	��������ud���&Gr��8�>��<��Y U��p
��vz��v�Mi1������~��߄�VV�tk����Xv�p`�BxT.�E�v���w��@W��D�DS��\���v��@u�m�w���,ݣf�3r\���x���C�J2x�>���w���ZfD��<�+U�M�u����g.�EV��O�~#����p�3��>��ρ�@��x�v�xW����Ͻ<�W�N�41lYsU��vT�^9
���[|=������8}r=�q��0��
��Θ
(��2�?J;�o����~������B�~�/��Z����=0~��B�]�L�v4$�]���lwY�`��Y~�l�=|��v\�~�>�x��;�>5�.��ϸ޲��QN;���}yjs�O�*G_�U�\�����x�B��P��B��K����ێ͞��+����fmWE~F_�y2�g6e�q�w��zKS�9C�ݛ쒊��)ǅ�{�녶;rFw���R�q���Tl�����!�����kǋ��>��:ξ�2�U(�����_�����v�`x. �,�ʄs��΅���ҋ�kۛ���~��Πi���AӄG�E��Y\`��j�^E��|�nK �)��	�S�cH�{hmcsm��G�띺qwʤGt�t�A8ˮ}g'r�ܵ�QUԻ��nS��heq���@u��ˠ�B��눝w�/�G��l������z{����NE��u���+�x�Y˭�]g��q�ٸ���UH�F�?q�d�*�ͭ6-o��f��9�*����C�>*z����q#�>�����_zbPz�;n���ʵ_����0f�{cD�N��.ŝ���T�;=Gc��ڈE� �;�	���-H�$�;���`R���+@�����O�5E��?|�W��+xO�(�������Ż�/�TY[����j�Ӹ�)u)���Hwu2y��9�/
�a�I������] u�`r�;�12�.��Y�ϋW�'?}���;#rx5����5筌�~���B��)����=��s�Θ�*+͓���`]�@o��dz#�D�gsꭿ�O�0�ǧ����zt��3k�8,��H�<�W<�>��ڞ���Cj��������/j�l5��\�M�[�>}�|`s�v1���V߳�ɭ Tye0/θ������7�w��<��x�>�[q8n;׷����R!װ��âƊ�թ*�[����Y�b�`.a8�]�9���i�{�}Y�D��Q.�ܥ��5V����C������=�\��]��X��q�@��5��S5�����:"��)��k�/ ����� y�{z�����7	�iy��m��v��N�9�c�ˎ�����θU��W��%��v{�������P7�����P��f��3��Z��Qqn�A�ʺ��ǯb�h�
d5�5��R��=���E\dϜ��L�s���o]��NU�/��"
�&�ޝl\��V�w��-���A�»@vK�=�N"�����~񩾳a�s�.}���Ĭ���8�R��i�n{M�b�����nwEu�-�r�{/˕�n2[*��m����Ӿ騿v�_��%L^�\�Әv;��8b��猆��Ϊp9z�F
�֬lU�?uo{�oؽ�=4g��N�w��X����':9�Gm���N�wO�����zd�}�B��}s#	^�Cb�EwV�0g��9�dG���j����=>m'�8v}�
�-�9"�-w�{bo�н![S��e���;�3�o��2�S�|K�Q�p����5�/��r��]Hܣ��w]sٷ���O�$w�TC@�{��:�v�m%��m��9V=kj��^u���V������B�bS
��4�*���$R�z���0s�j�峲�d}�zm�R�5
��G�tᾌM�����Vڽ�u�Kt@��;Sg�w0uS�k�Y��M�!��ԡ/9�j�J�N�FZ[iiU�Wع`�Y����C��T4�y�D� ��\Wmp'����-u6Ε3���Th�+�f�^Wg)�/#����`?���"]K�T�z=�_��?��`�_�s��q���[�]�uyJ���~���\��~��sҦ��+���ɩ��V�5����^T������y�fn�V��{{�ϧ��S'���\O_uP��h{��<�9���3]ߛ�%�Q������`�8L?M���w���}S9�\j����}����Μ�Y�Ǘz�Ct�b�}z����J�\ܛu�X�J��3�i�}���)��N�k9�+EE�?y������톶�.�h�����J�c��_?U�'�1��r���k�%�L�|"+��n������ܟ{�Q���_<�Kd�N�:쌨~����ϙ�y�6d=�����0���v�7f�;V։��M��+�ϻ�eY�lU3r�s�w�W��ɔ�Ӈ�w�����Fv��j�F�]`�-Q�hq�&��� ��s�6�M*���+wַ�YS�~C��3=/`�l�{�a��m�q��7�y��4t�W�9E��Cr�|�ި�Ɍ'Do��鳖YZ�d@��թ�v5�g����W��9���.��ou����׉Oj�8]��:��[��ڝ�k�����]�N��qN��fv�u�&�@�c��ηŎ3)Koeu^V��v_V7�Pc���Q�-u%�ԯ��~�sC�v\FM����mM��C�]I�L�<Ϻ	����o/���Ы����J���+��'z]H�8`�;u�q���2�P���Sf�C>�҇x�.h��ko՛�N�c3�~�yT�xѮ]�EE�R��t��>0P~�]������-�Ú[���S�3;�.cr|Nv֌<�Ƿ�0<��O|\��A�EwU̐/`�jz���vm��wA�{?\�ޞ5,��M�*Q���;����}��F�H]*O �����H�>���?{����,�Qv0�ލ��pc;]\<)P�)t�5��u����q��)��_;�Tf���s~��H>�E��m	�P�s�O���)5/��G��]��<j1� x�Ϫ�9��c��{��%�V���^��DY����1���z�i�v=���a��R�3z��d>������i���y��o}��S����u�_�������}��23�cKK�
�<�awS��}�{S�ɽ���x�oWk��cվ�d�_��d?e��}�E��6�)������(�SlMOIe�����d���K2G\��ܥ��unJu��47F�gVo�
�
9�/n  ��V��#��J ��$�۾�����tAw��{Yېl*E��=]���4:'U�r�p��#�gD1�`Ș蝲8�Ҙ�e]D.�=t.����j8�. ��N]mgv-���!S[�����ݺBy�x�Sa�~��d�������k誏x�;�Ǽq9Ȧ
7Y`6���[�K'�@�ѵ!�_��b�T��S���]���eQ�Lܹ����5�ޝ��.z$՗�gY��&X\sfXw��.���N���W����C��ǘ��@d�5qu��.��{�z�����\�����NF�T7��Y����Ǽz`��;��9g:ɞ�]T8�Ǖ ���*�{���z�u߀��G��Ke^M���#�64�dNB�L�y٧���������X��ĶoҨ��t=q�O�}!7�O2�"_u��+��A��g�ػ�%V�ѕOK4�vO�嫊�]7#�'���1(=�T�������]�Mf�܋�W�'��|zh��,:����ϧ���O���;��{ ��L�\+��L��d���NWgQz�oR�6�GE�wo���)�z;>��q��(��\&n6� ���`U��7�Ӏ��]�fg��/[�r��}fǙ�F����dɨ�/Ǵ���P�{�d� .-WP��DĞwR/�m�Q}�v�N§�Ú=O���\���;��U&N���[њ Ջ&��XŽ+jC��\V�Ή���g�68�(��q=���]�+PwP��v��'�'	��d�r��Y��ߵ�MC��3U���u�����L���3��J�C����7���Z�yꡑ}���e���Up���	��u,ȿ���Ϫ����{ǲ=>��oN�>�=�#O*�q�-%fθ��2`_�K���yV#ܰ��7��}qշ����3�zk�oo�#�|{�R�������
��`/M"��{2{�Vi}�c~ko�D�*���N�]�L�}�R��O|���}��+7r��� =Z�	�9�3i�iy�:�4���}�	�s�=�ճ9��~�d��!.��\W}�>s��&W�3����:L�EOf��^p��'ً�o�>��#��\��ͩ��`+�����"��9�����#L��z�R<��%UG�J��#Y�b�L���#��5�gY�@S7�s����xG�'c	h���0�}�<3��Oh�۩��ut���Z���>��;���/h�7 O_��*�.�Vl���	z��簯�ߊ�M���T���y�3{��:�|�C���ʁۊ�Eƿy����*�7g.:��k4`�<�b�
��0�-	�z���{�]�*�;�������z�%�v'�1Ս���j	6�7�Ǜ�u��1-uf6��\�z8�f�_w��Wv��,ۗ��jrv�>�L�ǫ:��oh���#�g���+��d�����X���t�tsqܲF����ޞ5In{b�/�;�K�|��yS��h+T�� �n}������Y��;'dpw��A~/Н^�g��s�7!�qњ���GG�%3�����}}��+���%�v�q��>���/�k��3x���]�,�*ۻ�"�H��\V�T��v���{�� ��D���������R�ބK�ߤn�[���u.G\���H�yft<�]����w���;�R�5���u߷o�k��%
�QO�.��SC��}�	�O���*����x�痊�@�qQ�<�J�w�2�|:h�F�@ϧ��w\-L�F9�{c��{��b��5s�T�w`��v�_��c�j���������U�q��voi�&up�S9�_���>��}&��`q���cF'Y�bg���eD&<�\���o�u߆��U��k�d_��y���T�ޥ��{�N�C�b���Y��Dn���S</��z\���Y�3�}��7ҁ�~��S��O@m�g����n=��
KV6_�xcV}Z����I�N��.�룙W�% �B��٤��7�,��U���\��i��t��^Ѕ���������W�����Cc����0X�:��r�܀-�Y݁\���,�5�FvEs���̿��g>���i����>����DOz�
�-�4,�e�L�-�#ޙ0�OK�����a{�m�R��S�]9�*���E��T�Ĺ�\�u�O)�М�](w��Տ�r�Z{t��g��ڰ��h{���"�1�7Hp�8��D�*\��%�x�2���vפ_D���`e���L���̮�������5���9Eށ��|c;f�\�:��[�J�z�\N�dɷ�7�L6��r��.��ǋ���h�������"o�,^��L��*N�I��u�lG]P��m;��Bo'�M��C����OW��o{����[����r��D��}8���tDӪrtg��7�A�dݿ���6�/o0������K�+S̞�.w�_}2���;:�z�ʃL�I|�KF�bP��P=��uD;	h���ܰN%^w�c��<�{��KKԤ��(���������
����T'�$nV���W�ٽ�fs���|��M}��U^�
T%��]&�>�#2;��^0~��Y��+�������E?Z[y��Y���iv
	���6{{�o0ڜ/f,b6�����hG���nj�+�u�K�q�Z�ޥک�_b��l�b����`��m�mr�i\�����h*��;�㦶�iR;g�J��)E�7��Z��n�6��j:�y�8�-м}(����U��X��I}/n=���F����,�)j�ʹ<W`��6�e��/H�m�����%�ލ�8͙�<3��EC�\�h�T4)���̬6�D��:2s��=Х0��惝e��K��r�.�Ը;)��u��JWW�/�W�`zt��e���Fث��J��ʻz�"�`��@�u;Z�}/72��H޼����G>^nv��-�눎tn�^9v��竇uKp�8ч��Zɥ��5��]Cp̹Wd�E��5�
p�@:y�+v�-/�;{��[����l�(e8��
Z�c:��Y�P|{)r\zY�)R�%^�St�LfB�'��̰b��v���2QƁw5n��i5�f��̖�<�]�}��d�Y� �������a�ڐ��Ċ��l�k�:5%>G����ٕ9�/0��������;ڿH��v������11�Wks�_Pz� �[�H�u=H�<���Žq���` �}�8uwq�m�Ạ�xN&d�vr�3�Dn��f�g���5e��oO�V�׎j��س�\nuG�Z��^�%�){"�t&��u�nr��]ԶtoYf��]y����ҝ�b��\��K��,T$�;γ8gZ��Cx�	@h놼'ub¨��9��,�[7b1g+���z����������-���d�`�� S�q�%2��7��K1Z�EN�ZBd;N����|(fֹ}}P[��ţ���A'\"��ZGR#Q�InhC�c��(�*��d��.UÎ�N�=�I%c@�5 թ�s��Ł�0o݄��38�q��ɠ(����ځ[Hu�5���X	�HD�꽼Pe[�VѶx�j7+�]�n5.���h�u��n��膆.���k�fܣ�\��ol>������H(�!���Z���tPW��Ox⮡N�0��E��,<��.����f��dfc�!<��MwU���ó{����_s�{��aY��n*�	��*�ueZ:�\_J��,�}�V��{�ښ�zQ=r�$����w*��:��s0X)���:�9v5���ɘ�q�g
����:�ʔ�F���.8�&;�]Z>�Ɣ���Zi#O���v���ʽ7[�Xm��'Z�h�2�N��Gfz���c��]��
LF��!�U�G���ذKc�:CkN}w�fp����|���>�	]$ �ut-U�EP���8T/`�aӣ:��,�gK@��`��,��*>F����rf-��4��	B-��5wP��iX�]�))�وD�e9�p�L.esu�\��}`���KL���廵yf���u�ce��%��I��.�3K�(�p������me*�N5ͩ�����
9]!`��x�j��֔����S[���cZ�p5z�s��\44(XJ��G�4*�;�GI>�u����rv⻷\�2�0��nd������=qr�̂�4�rJ�P��%��F�$���ҥC����>�OS9�Y�Iz�9]"sg�z���w�
{����'p�=���"��VZ�sQ�������gL*rs��K����J�>�l�y8w'�.t��y;���6N)�x\x���>��fA�t�땟uz�y�{��q*�hZ�P�GR�$*/$̷Wur*�I�"�[�����s�n|�Vt�s�(��z������s�T���;��tI2����H.V���<<��gԯ^��
)!Y]��9R:8�!.��2<�,�ws�U����+�L.�F�n��x窎�<��-�>�y�����{�%���S����O{ϟ@���GR�S�^��w��;�V�����Q]�m)
���}Ǚ���&g��iHK=���Qu��ޞ�r�_n�%^eB��y�qv�"��Ԥ���$+'[�yTPc��J�Lz����H�p�̔�"��Q$�2��Tsۚ|��ԝ}6�ZJ��	��9V� ��Ğ����,=Jø)����u;�N��5�b<���%E������gqf�.;��eM��z��{��f�okf�7�����&j=P�һ�/䪧�Ǻ@����Emk2�uC��]�u8�Y=�=��Ȼ������gӕ��NV����g�����Fq�2W�3W�c�ß��U�^c�����3��5��r������Q[|<}9���¼o������^���ĉ��5�坚�����@�Գ�)�t����{},R����l{�u�������ytT���[|�{3���*��q� ��Ks�/������Q���
zr#�|��_���&�{�����3D�����ф�=���{zhy5LL�]��+�ưP��bԩ�B5��n�;���e�GU��|��W�\o&x.9�l��]X�ҙ[�v����~�9�˼����m]d���9��r�~�W8v?d�����o�#na�t���/�ӑu�y�e>��������W4϶���E�+?UHʉ�h��G��Ke\d��ˮ��D�/����W�^���\����|W��ϯ�;"�u3��ĶoҨ�u�^�?ܡ0�������u�o�?<z̱]�$����}�0	��f�p8���ᥞ����#23�������3#<�qdt{�3WNՓD���1�ש�J��J��|>呢T�}-iC�kjA�nMMi�WX*)�-λT��6��|�"�[�\�H��{����Lq=�B����H����E@���j��b��0t=�˺%{�ǟL^t�ru~�u犵E�����g��	��gt�|y����vӾ�Fw���L���y���)�C������X�t�n��e�u�ǳ]Y���{��[�xR��7ps�g�
���`j��U05�>'}9��q���gu��:@ﺨ��*j��R��L��0�ӟ��*zL�] .+t�^��̂�j�(g0;�xW���E~���<"M�~x�~��z<f}��T*b���#�UW��N{V�r*c�D�5����'���Y�o����_n��qV=l~T�����1�J����ѽ+��L�ks����P*1��������	��x�s��������:��.L���q�]����g��xl��H	S\@޹�=T��ٱ�}���s��>��w/||b�$*�UgD��Y��l��׷#ޥf��v� 3Ѯ��'Y�q�x��U��o��Z3�ܩ	J��U�cҏ�E�*x��N;=
�~���dϺn<\Γ�=��)��<1��w){��غ�tRA�],~�h8�z\�F�#ǮW^�D^�x�蔃���������wB��`��t�L�����MP5�� nJ�?/y����.�`�����6������b�1W>���\;7U�}�ң*o>:@˱[� ��(56��guVס,�CZ�.s�w˽RͿz�o>s^uV��슼��ɞNs�2���ܲ�T����e��T�\ʟQ�)��2�z�ϻh
f��0�!]���E��,_�2������w�����{c��o�ԅ��ԼWϧ��V+�ϑ�,��tWY�-�UU�轧���,���S���o�3��f|[/�Ձ��J.{O�H�/�8aЪ:��ٿ�g�v޿(�3��Y���^���r2+�P�o��e�q��a���,\}=;�3��z����n�\wW���Sןfc��N{Nz�I�~�nzI	�㹡���f'�VG��ݨjv����:���E�KԻ���z��J�#�R8�Q1:�������o������{���}T���{��n�9w
����=����"��WI�!�ƥq������F��>����s8�*�}w�w�W��Q(tOG�k�:���Pe�n���]](�(<���r���MC�LVG����e��9z�}�w��U�Ԧ�a��.����. �Ď���ܵ&��ߏ��֪�<E�[�6�2�P��|qi�m*��ǈ}!C����@���j����k8Ɂn��+�u��ؖfR��.1��l�w�^=�TRcՀY���yWeR���G�q^���<7�r�޲3Oun������r�/KJ��D܋$Q�ң%v���-�(��lǺ���F��g�Ç��w\.�dc��<�U�CSb��~��:�-	{�~^Tnw}
1�s]�:ۅ��̨{���{L*��Z��"�����������a�Kw�[]����%��U.`v���m��ŏ�t�.��
]��N9���X�RV�e��=O/E�7��rI��n�+���o��>���Y�3�iC�o����~��G_f����_���2;�S�s��3QO���x*�����_���|�'̛�2���#�����G_L��,P]�ĺuϧy\mwPF5v�v�I�\�]�6Ǽ2fI�Y]5�ޮ�`���f�١�g��XMmXl޹�����t�_VZ2�w��)��������U3 Ϫ�ڢ��5�w���ܙa��s��k���u���0t�SQ�z)?v��tVۋc+������0�Eu���ɷ�70ڛ�ʇk�#���3��g`��uY?���������c
��Eǉ�����u�^ӿ�l�;�ܦ�v��]R��Ȫ��=S#�7���Z��ީ��R�e$�ͭ��XgC�h.	W�)ɼ>�t�X}jq%�Q�wʟq�Z���>���â_�����ޥ��>;�M|��Z;�X׬i�r�r�|�ܽ��MY
�k����Ԕ�/tInt̚b׽M� R��ػ'��N�,�{SǽS��n��C#�'���Ġ�=v�;:�0a�K�ӂ��(����
9igc=�TC*c�\�ٸNxq�����@��BZ7�LN�܏]��n1je	�/�Q����F��݂��O����M�*�\Gw� ��|nĪ�Ϟ�B�����clk~���;jT�OF�9��0�������꿶��BX���l�T)�� �P�i�p,��[�Y��y~r'����F����~ڬ����Jx�ߋ�������}@,� ���r`��*�n��Ӱ��87��U{�~>�t޿�m[����zf8��x�&7������f�7ז�����]���I�ޙC��V=��N��u	C�շ��Ӛ{	£�G�Y�����5���2�Ƒڷ��[p*#ec���v��rʍ��w�p�<�;=#��"�ޫ�èa>�&����åk�:{�=���ڐ�{\ ����q�v��Ճ{5YF!/Ǥ��WЪ@{Yu��>�#;�	ܧ�7�t/&|�2��!�\F�XMK�N�ǲm���C}�����p�͊kӞO)��ڇ(�V���)�٧3mA�I�t�=J��� Їf$��fF�����=RvV���_�K3�i�Vfԉ���f��;�3.�Nֵ�0փ|r���˯����8��YN�S���j���d*6%m+��k=�X��J�F��g�zp"��X~~ȫ�2��ɞ���_{]��^�c�8{�<žQ3y�8S�ukVt,�gx^9�+�6@�����p
���y���C}+���v��t���e��,��*v5�����^���u�ȅ9E�����t�Wt<u��G��KeR��v�������q{k��l����#����K���2lSg��]�WT�p;���(��7>�Y�Nk�t4��8[+�kC��Ӣ�t�SC�����(\>����x��>0P~;�w�@���̸�mn�PE=�*�|ry�}�c�����O�����Z
�<�!�]�� �����a8�K�.�J^ϸS�������rp���l	��x��.x9Fx ��}˼��l��o���^������w�d
ڢ�`��>����ٗ9V}����}e�
���̲t7���kF�r2��=[�|�
���S����]��l���iO��^>΃��x:0���y��n��h�|�NLT{�O�Uá���u,ȸ��gr�o�6�d���Ń��vx�g�j$סE���^����`����F{o,�Ǣ��R|�݊/�����$>�A�k.��H��5�3�>x.�����J2�p���$K�#�s�u���qN�,���*����.�\�ݥ��fe�f��3��iM�OT�^�2��ɻz:�	��pũP*1���#+�s�`���~�j�}'��V�w��������״w^F�����Pt.�ptw��o�(l�ѵ�J�d
���<�������7���|���L��:뺌Z}3KV��iϪ&�}���~�Tq�3��\ �k�&1:�3�{��*���y�$�m̊���Ҝg�zUL����:w>�w�K�Q��~�ȫɟt��.gIឍ�S���h���:�gw���va�׽hkɔW{�Yx�<
��O��dϜ����L�⒙3�w�x\{5��gw�ڬ���J�֝.��z+�+�@�TK�a�+��)����X�+S�{���by��\�C��;Q}�X,H��u�>���j��aMcn;��͖����$�\ϼ��Gv�Z6�l��r���Ke^M�f�T�����$g:wwЧ�y2�q�7��\����ٝ���/����+���\�g�V�b���8Ύw�#��*�5Rj����{�����(���oC29M�I�s�hz��ـjr�=P����3�x������%Q�4ߡ�i��f�'��fA({�ڌ���{k^ߋ���\-we{T��������"��6����R�v� �22��G@n����Y�%�S�t�֪>Γ;:���թ8�WMbᓳ�5��t�Oj�;���3ϥ��Z�
��Ve�suʸ���GڶJ��(W'�EE�WI��.=1)����������s�/{�*:,s�cXc}�)B�;��{|E�a�<�@UݖE���=����M�㾍�j3���s�u�����8ǆv�ڍ�
�<�g��&��08���T���@sā�Q<���W�������c� �⏚AN�='�ޞ
�����SD�T:��:B�u4:�m��ɩ�9�g�c5���p<�3;�
�W�=�����/��:�G�����\)�Ȭu���Uq��MSQ�îv���o(8³�'�~��d��'�[5�Mn�~c߄���]�U��
�7��+`��{��~��V��Tv{{0�����N�g���u�#/���Gd{�^7,t�ip=Q	�@t�_;��y�>�U��y;��<�D5�����i�����6�R����'�</j���.<�yϻ�
��ꜥw���J7��I9��{�n;�w#��Ey���D�pq�d*��xhT�8�<H̙�����Ԟ�����3ȼ�ِ���X�MSt�N:�����aglU3q.q�>��rd~&��
u�z���l�A��-���y��oN�ܢ�;�jS���3�P�s���F��u�.��v�nZ�ivv��u���L6(?S{��L)/&N�[���|e�P�wԨjᘏ]��o.nۗ�c�i:��_p�˫�f���$��v5ܴ���q�Ĺ����5�s��y3�o�av}�a�q��g�SG}���Hp�u����/N&�Ԡ��Aռ������j.��.3%3y2�G6烸�Ig���4m�S���*�xG��z�U;��C����~�W4=q:��/�|f�a�9�0�u$S@㴽=��-o�x﯀G��n�l��ީ��]`�2��k��Xǟ�n<��T�����u�������Դ�#�J6�'����"��S��}1<��bP{����~2��䫚�%��INe{v�OR=���ݭO�Lx��p�����A��깒�-�z������׸��J���y��+)p;{�uF��/N��#�����7���T�lw{ uƠe�d��˟x�j�ls_�n��S�k�����5�`u�/��4_j���]��������/8:�'�)�]��IP$od�k޸y�t���Jx�ߏ6�/�H�7�lV�3QGlȷü���}ު���_/�5�qzr�k��NVq���x�&M}����p�+������l����X�{��Z*vz�U͏Ֆ�z|�Ǘ���;ge%���aʾȝ��X��{��������)mƧ{z�������3ǥ/QN�|�q��k��tǛi��.�W:��Z��'ܲ��s���N��ǈg���rfftt�q7?T�+�q�s�:g�k��W��T�����:��{>�z�w�	�]1��Om�yvxd����細'�T�l���/�=�1�{���.9�V���|�ݑ�]�׬Od�_?ma+R�+]ic��U��<�jG{e�<��	n{���8�_����
zw.0�Ɠ�jp����/4Ϯ�FgJ%�u��v]�ɟq� '�!�~޼KT���l!���fvad��r㗶�C�.y��edu\x
�~~Ȭ[����Q��T.����l�at���t���[��^�h���ο��+;h
w��6��~�m9��,�9��T7*Vs�{�����V�^�ч�{N"�iU��9EϽ��q.�{�+�;�Wo凇��������a��7?+�ez�:�WG����H����9�|j_\u�U�X��1-��� �:h�S^�
��S��3�yD޺���p���ʿ�kC����CJ.l���*�G�W���þ��|ϧ� v���g,��4к�w���7�V�;�t+��c����{�������?~x�������6����A�lcm����1������6�6���6�6���co�0m�m��`����m�m��m�m��m�m�v����m�m���lcm�]�lcm���������������6�����co�lcm���
�2���a�r�������>����������B��T��%!�J�,�ziB�TQ"�D **�lҒ<�H��U*T%Q*�*HUm���٦�M��R6�3KT+�SVTD ��l�38z�G�I�����a�f�40�
ppvҋ�R���9`�Ű�hK-v��-�T��)X���s�[h�C�i$�݋��j�LB��l�4�P`2)U݇E���b�X��f-�`��������DNZ�A�,ų5��٫@����)�� �[$ړZѵ��U 89��[i����l�&XV�"@��F��5��KM�F"��Zi6p��&+khk4bf�emaCKw�   Ob�U(       ��R�� P44dd  �L��i4�M�F�Q��Ƨ���~%*�       4�ɓF�� �0F`��J�I��4b1=ha�&p�n�˗L�W,�2�7)�tܨ���s�TU����� ���H� �T�Ȋ*�Qe7~�����?�� �>Q��dATR@��U@�#T�`��**�^_��)��`�㳷�؊
�cA�uJV���R=��s�cu*E����ߢ��d;�������[��7\��r�
Qسhޛ��)J�
��aU�V�qS�mkѭ, τ�2�`9{t�ӣN4��5��OT���4�`��.&��S�_n�(�U��u.�����ł���f#c]Ի�H���e�CK(�!�465Q�b1�Q���^���+{��Ai&�����ɒ l�,Є������G1)P�n���C,�i����s���5��+N�ոi�(�h�552��JtYJ�
�Lך�ܕ�V^ĉJ��T��j�w���b\,��#Z�7�o2T�P6�k #,i�B�(��fe{�1Ĳ�M[t�I��C�k�SS��Q�SEk��fr�E�ySh����-hĮ��D4�<ۆOiRwh�����q�&�[ s*���Wr��#4�^n��z5��4�s�eH��Y�YiO��(+(�)�cN�f�VK.�܀���uJ�����b��ź)�VL-l]h���ӭU�l��bV�B7�dU��.��U�њBxZ��W{n��n�c&���jK@�ۭ�a��8���ܑ�CD0P�X:ln�ߙ)�2Z*���Q^n3������@KLi/.(L)��ز��@ ���iKͅ�8�� {U�K�V�_���5ږ�n��]$Mn6��#G#GAפ��ּ:��0�oF�n �n�Ab��]]'�y1�^�	��"��AL�`�X���g#�EJҤX�����h��Y�\j���&�_=L^krͭm3[X��0�XE�Ca�1U��k[Ge�6mIFR 7��G6p=U���Px%ZY��,���Z�Yɶ)F*�Zg]���7`����S!�w.�rʁP��1R��	�r��j�R ��&����˷���:视��̫�TD:��h��Ў��*O^��0���Iz�Jw-^書�i�Tw�鉬l0]������\!��4\2����ۤ�ϦQD�W�[�o.4UOVj� �4��!��Tu��ӢVՋu�h��f�A����<�w]b��L1��-��@R�W���'�*�/�LwN�kA-�R�G[{m�\eTq��Ac���/�	��eʕ�B�>��5/F��`���BƇ{(�qX�@ Ž�J!mE��Z��V�m�"�R��z�5řaEkhv���i�q�)̇��=�E�/El;nSc�&�u�t�����3JT�,<�X)TWz���e���"d[9���06�Aq]15g+vR*�*XB�8��4�^QPiY��30AkE'����mh(J�M֌A������Mh�
�U'���p����ͭ�y�Af:���Q�L�X��1�F���86���X�'��
7���J,`b��y�/��Lr�F;�E���ެ�kgҊ��FLZ��$�~zsUCO��.VS���s��'l:�䙏Z�SS��l}�$em��XK܆�Z�fE�(����B�?�p�%h7%6J˛���^mfO�)��%TeӲ\��53u�gt��ZA�ielwM��@���"/
�gi\�����ۤ�j���9B��pX�*�۷�*ӑ���v���x�d�`CV�/s&YA��m�*�
m+W1Qw)�ZJ:X�([���*�l�55R�OjЏwv�Ҷ�Ԧ�ʔ]
%E�Cy	�onyy�m��fӣJ�T+i["b�h@�2�ƅ'X��Y�0�u�[���J+X�f�T	��N���pa������ n�v�,x�+�՗)��Z
F#e�*(�}�H]#�`'d`i�9d;�nT�#[J�KU1-�͍�2��۲c�k7v������B 1V�dK`��v��<袎V�P�+eKQ��k�ok$p2M5YxPZ��MR�����f��>��z^���*�nv.S(zmVXZ�G.ɸ�(�#!���5b�eh�H�ɳrT��-��Aئbx���3����'(+8�Y	B�Э�Z,�pM��B�k�6�J����$�ywi5z��=�θû5��������9�lJHy}�JrC��d?�lE��������xV/�>X̤�D��7[�V�P�ABt��سo�K�� �tw�ݼv�+�޾�e�1ͬ���ã
��k�{O8[�˜�q"P��q�r��­X)�8n��1�}��"FZU5�Z�k3{;Jm��pn�������"����X�Vо3"�HU�����1|��z� ��FD&rs�^h��@Y�v+�][Cj���7�E��1�шy3r���YZ���#:*�.c���(U��X I�����d#kT�X���5�(jY'_^���8�s<�����a�^��άH:��f�5ݪ�a(L�'�:\�SC�:[W��]2�z�WH����<��c�j߻ƳT��aR�8m�4
�J��8on;�4�N��pۦ�63��2�ۋ��k�h�(���*���wՎ�.�7�2 6.�0�}���̬ś�qz���Q�N\���nf��0��2�T����X����t�l�s_Uǆ�+I�W-	DNX��3���\�Y2%����pdE|�f��ﵶ�'5�aG@�m@腚�\�a�apɝ���fq�Ä�:���%r�|����-��O�Mc��<z�pے���&}��]��B�Y̡��O&�w��C.ԭJ�,7�Cb�˸'N%<;�܀�p';�5��p��R:��n�N"�PE�ut�y���\5��w_��(̫{��� m��m]��_�2�i�-���9�a�%I��݌#2������pw
B�f-kE �F����wĻ�L��Zo{5�GM=�5��^���ԭhѨw:aW��>g��`�V��vQ;���J�Zp�:N�n�=�����*qv��A1[��K��]������egBz�j�=�ŖK�ݮoM�Hr
�ݶ
�"j>����;�1�ևYU	ʵ�y�i�J![�6$M���f;}Fm�� )١Ewj�]�]���4j.a�@��T2<��GE|�(��м�=\�}3bn�7Fn�X;��Q�Ee�ݓ\�0�e\�Y-*�5{��%��S��B��~:��³b���c���-�w)��|!�cV]:̈
�5gn����j��&���o�FcSoz�Q+�]�>f���EK�/��u�ʙ{��5Y�r�D��7�%L�+4�]�.�$KmV�G��@��#4�	��_�Wv�ب'�+�XZJ�,����dx�I;�PI�p:&^y����IN�XW�a^ے�3��D��v��A%������N�<8�v��j��K��j��Bi�0fB�x��6A�Cz�t�͎Gb����cJ����ge��m͕�j���6�VzS_m����ދ�S�Q�T-me�nd�F�f�
l��V�۬xɷ``n��b���wN���V�.H�Uцܽ��3� �������yU�J��Cr�`Qp��R+��:ޠ������ӑ�WE�ֱ��I�C�����3��@���;�2�����Ӻ�.�Ym�u� r�.�\�}ƕ����U�H[9�ܡ5�5����D�������:<z���v����o�͏hI�����	wi#flX�G}`�VUsW�a�{3>�e�B���գ���]|�SR���H�'�^٤�⎻���"U�R�Q���	VQm�]��AHkW��{�_:P�{���$�.Ь�3�+C+��������m�2T�ٛ������@�
\j$�[N�m����V��)��\�N�Ri1φ����}&���9��67���ŧD�;8ݦ��v;y��Ku�Y��f	��Q��w���s�k�L�����619ܡ���e�j��i*�zz˹�r��p����>�������8[B���>�P�����V_�:��2�Q�mQ��V�8'v�b��r��e(�\��1][�9sw,=[)�����v��[6E�t��s�_p�*'s��h�'�)�:s�K�4���c]9d]J����J���&.F�u8vqf���gS�ƙ��[��y5C*�M�{xT0�����YԘ�������KN�W%�ٻ�%�.ty⓶��]ϻ�����k�N��6�]~����EP&i���(!��T@�LN�*���t��9۝i��Mi�J��ږ�nHs+�Ҵ-�R)���݃��z�+4q�Gq\'�ᓴ�x�'B�G�]��ua�kdst�J��n���e�]����2v����k�|-�з��i���0֗��"�*EB�<���=v��v��/�^j����a�2��`��)��)W�Ae�;ج掷��0���D�_F�q�t0�=*S�}�2	/{u�=�)_��|d��!��c�˷T��j]�Tne��6e���)��wU���gT�be���2��Ӗ� �ljq��[�ك$E��5>2l��� ��^��:�G4|4���������ݹ��tu1�-�UG.��ROk�Qq�z��XM��D;Q�:Wi�ܹ��y�yX�mn>��o��*�\n��hdBVښn:�C@���6w�vn��=�e�;A�X��C��%_%yYM���7	8h-�wN�W�&4�m��C;Px�y��������X�E��A������E���u��H�hv�Q�o���5������+�,��!�K7@Ŷ~��NA��i�+��a&��l�Jn�X��j[B�vx7�T�,��2��64�G����dmj��;���6�pN�p#�p5cz#��33.K!�r׼Ѥ�:�u��`�3M� ��j���Yゅ)�����w1�u���!AȪ;���8_Mf�<7Bqi�wf��a]չl�%\���yWs�
^��#%�Sb��\�ܴ*e�0\�[�v
�4[�3�;�0���e�s��ꏧ=�М]Re����KY����e���˕���z�l;������2m�Nq��Oi�頷�e>O���<�������ME�U9mw_5c�mӢUԖ�F/�:�%�3w{�V\�ZQ�錷��]�qٸ��Y�Rv�&:^�܀ (�".	����V�q�{e��g�qWi��� �=�wx�.*�<�����	����Ol�F�!Vy��U����»�*�_* �6��$��v�U�(U�g^�R���ؤ�9-Vm��Ѯ�A��R�Γ��t;��k����qv'��kp�B����#Z3��#�ה�������1�a�s��WAu2���;c�b��*�d�����jc�Zh�e�MM�մ���\��Y 
�u� �@��2���hh:J�Ȓ���n�r�6V���H(�e.��f�<�t��	�j����Be��1ܼ����PW��XÊ�K
r킘��=
�T�%��oR�>Ƙ���X���EiKl�kpV�Ye��(�\֫�Wf�F��1Z���$�m^oK	�t��*9̠���"�u1GH��-�a��flˁi�bA��'�9�Vd,'�Co�3˕�Q�#�i�s'R�� ����'�}�h������By��mi���gL����QVU�u�}R�F�j�OP��KM��K:SK(*@�.��.�t`�ʲ��ar�]s�&wm��#��rȥ�l��{X\�k*t�3�-�4��g>	Nf�^�Z��ڵ�+��iKn�����w�N��j�[,�W@
�*qr�VZ���m
rp��h�����p����"ܷ�p��X������؅�A�
ɵiK9]�r���	B�T���Jb�Д�c�ܽj��XmE�/v�>�~�5y��Yu�fi��J�V��`�E��9�q����!��tv���W���6�;m��\ِ]7��]�J�S{J�*��ے�ې]nwۏSY�-���2� ��K�oH�p�a�g�A���wZ*��/��W2��=��a����E�b��Yj�)��PY��gQ�b����2�q��] ���u�\]ZN���Z@�m�j)��Ѧ�|���Hg]�]�o�譠�̥kK��U�m�5ֻnV��i86sknrj��X�J�b݆��:�ʻe��;��_=d���]v%�6�,�k����f����b����S�`B�].sGT:k"�����
�t���Cp��Z�/�U�v�G���O
��v�Q�Ӹ�#�[�{�l�vB �H�}(Xj��cT�:]_�_�Z{�/���#���~������������Ra��`���i��=�9�@]L"<���+<(am�`E���,�Ubt��QIU�{LT�L�X�]�����>����O�MJFI�P�XM�ն7�F���U%��Q�:��d�U��zU��n;l^IQ�->��s8�4�yJ��4�Xt�Ƀk��FC1oV:�i�{��{�`���rK��J:�^4(�}��:m��r�n��j/q����}�N_�[��}����մ��v[r�E��R��0E�Dq��%L�.[vت7d-���\�.ܗ�X��[[��I$�lq�c�Q3V]�31F����1�n\&3,�f%�"62F���[�f`fIrB�%���j�[u"
���Z�����B�Օ�o��ܿWkÓ6�����:�L����������cfn��bl�[1���j���G�ܔm�a#�x(�ϴ#쮕�D`��)��!N�XK�����&�6�X���u)�k(�y��ڨ�*V_�'�y�yw����
~��,�u��0������r�Q5���Oa��~si(|<�����6���}]�Gr\�MP
�x���Ow�%�E�N�p�����a:���V�-�30?mh�S�����⌽�|u;5��F�������!�S��_��oϵ��Po�T��R���`�F;Z��ed�dSk;�__�B2�T����bv��3����~w��	����!7hL�T���gd�kpL�J� !�ր����+-�W���`�FP���k�tަԢ��� E�=�k���p!Z��Ӎ[N"yZ_^�f�A�{�Lk,��BE��*~0:�ʻ���+P����o�Z�� 	�<}0��z,B��\��w�f�^��0ߪrߥ�E:c{�H'x�Ey�N2w��V߳3d���[�msn u[�:�A�G����Q�:��sY��Z�k"�&U{#x ��I�u�S���h
��3$MvC�u����
 ���އq�5}�U���.1&��
�縂��.K�y��v����}������Y�_?c ���j�/��uΝ5J��Z��]0����jG7O^]��U�|rAXt3���{��Z��(�:���B��cT3eVC(���ކ;SM˄:~��>�9ۭ=`]�r߆`hR�r�k+�7^'��[�q��i������Z���0<	}|��}���xؽ�+Z��m���K<�<U�$�]��S��C3��f�y����q���Pt�7x��H�e.�C��$��;O(��*��9��Z�F �YC��1ו	g���:k��|1�
�Wy�"��ѯr����L�c����cF��O�u��~[�sY�/��rz7C��ύx�79��e=;T��a����z�a@'�\�V���Z���x��fp
��&αIR��`�ïB���ڮS�ޗ���-�-Q�Jz��]h�\�~��N�i�X�p�7:�R�m�1��"��;��{�V����^��[+ժ_���M8�>4,>��<p��wܳ���.�Z�{%Ԏ�cY���j[4��U/;θ�(����`�vz�a���e��K�VQ�{�#���l(��'1����/�{@��zjÌ�ƗUF���0m��Ol��������f���r�R�����/u���h���=�#J���[/���ù�����צ��y��E,�>f!u޵���Eg����4�VU�D�m{p`��uNz������e��m@�;�gS�?yr�WlXɿ9�U4,��Sw�a� W����o0��}�3I^l��у�!�0�wŐ{s���l�o0?f�C����קF�Tň<��j�U�b�ÕWr�1�A2�D�T�J��"�U��]J�OSohl�4�l�fQ�K�������;����Z2F�9^���ү���[�iiK�Q�Zb2�lGم)�i�~29��!g=:�e����zo|OxP���Z�b���kφ
�+��?2w���zQb���͢��^��e���8��G��0���R95�l}����ɹ�W�{�����C3C_�����	�-|kID�f� �X�	�\��&��n`�c5���\V&V���*b�w��R�V%��\�)&UьwLa.ڱ>��h�+�5o_<81��c��"��	��o���v�=����6� �\��}�v`?+O_=́<w!�6���+�K�9�3���]���j�/�>]���@Ɉ;��;M�֋��:��NP����d�x�����}rU���'b�᠒�Ó)'Y�?Y(bI��#�F�Q*˩@XIJ��� Q�Y[F�.������4F;VHtռ�D*
x�'�ڴ��6�m]�'�aP9j<*�%������P`�����R�!�8�*Ѷ��R�`��q��c��y��h�q�Ԕ�eY�a2¶��ӡ�Q6XpQ���W7Q2�`���ڻ��p^]��ѹp�F
]�����[�6]�˶X�$�]]���Ж�V).����*5��0�3,���\��v���icmZc�2��J�H˸]�j�e�d�Z\��˫n��f^\m,��,j�[%�`�f�K�Ka�����AW�im�6�Ҳ����EE���e�n\\q"�-[v�H�!�[�$�1�F�7pH���K���_����^~�7[�yw=�������%����T��e��0�d���=Y�G����'�廢3�q�^��r+�����cE� /���~���Uˡ�=��gr���.�uaj��V=�gl2��9J�܄Xr+ܲՅ��F��A�5tk�m�zB��P�e:��NJZ�u��s�ٗ =`�~����cK�����T�ǈ�;Wۗ�m��ďQ��l_��tx�U��~������ܩI���}�*�7�,����׈�y�c��18+xx`&dU����z��Q�rel��z���Q�ML������w��v"b�i�����{� ��ݾC,w���R2�~�l����w=�J㻰��wlD�����g��ww�Ɠ�pI�_i�}�׳��~�����i+h� i���D���i�G���w=�{����@4|�~�UG��(�۠�Ebh[V5T|�Ui*��t�w��UJ�Rg!x@Ž5��qJ+G�j�5X�Qy�ӟ�35�悪5K��JE/�:TC8��KP�(y��}�}Ϸ��W����(�Tk�G*������>J���s�r靈��!m���U���?%Pi5@ZZ���F��j���{��J!�}���X	�SH�U�X�a
DO��7oy�N�](-
ƨߥV4����ץi<�j���IV5T)U��4W��S��ߟڿ����W��r��Uo��Of?'�7D��m�+�g�o��{�Ϩ�m���6���Th�(1��U�Fo� 6�XzQ���kܶ}�?5UQ+H���!�ƨ�S(7���D
D�**\��l�Pܢ��u���(�D�� ������ kr��+���������T_���QR�a(H.pB�L�"^ Y�&�뮚k�j��*g 1���UX�Y�UD��@��kmQ�ETh }�|��>9UDB�����,j�{>@Ī�J+Hv�P�Uu���L�P1����⦑�4��(�J%U��u(�EW��Pfv������@8�D(<�F����?&��9���Qփ�U��j�ky��Tm�?%UD�h��
�Ahu �U�%UO�j�;��۠�UcG�Q�-"��H���SL�!�Mo��� ��߇�~c�ӵЯ߫��`_�����y���.��j>�}_qH����B���A�1(�j����V6�QhJL}��n��Tq���H~j��C�4�|�m���Pu
�j�mW���l4�Q�(�A�+�A�_��{=����/�K�:[o|)"�#��{�7h,��c\(κ�A��.
S"��+�z�ֵ{�:�2v�
zk�\�^铵��n�S~f��.v��ۘ��/i=����~�$a��J\���n�� �b̬l:�7����[��7Ӗ%��}��M���V7W?E���f�?���gm�n�)����Y`��p��E�>u�i[�ʛX��j1�$��Tٞ*�b��-���@Ob�&�6S�]d�2^�m����6�-�I�_%a�nhj������{`�;�<{Ul���qJT�J�6���]����9�dg�󼓺?�U}��a���]��kj����e����k�=czթ�n�O�2���w.,����$]X�.�{���d�U��X�)�"�s�3�)�� MO_^������`� yVtI-�r�\�I����<���T9�i�^�N����c�R�������>�����;�*j�x紴��c�8G[�µ������J�.�OY�?�}��U@ڈ��P�����덨9l���7{yڬ�pNgKof�̾�ءn�l�#㯽/���͖ό�׸�g����%G��GL���v4/|�-����~���2�b��w5��O�.QJ��.�j�T�j�	��wA�k7/�~�^f�;�@w����R_82����2>��}_}�Z�T���/ߴ6���+=]�_����S�X��s/�N��f�̋�HW���Ȧp�z?7,C�}�������S�ּ��啑�~�Y�PͤNT	��� �:+�ӛ�B�jn��1��
�{�7��D8!O�S���]s'�q���-�*T��2OK��~��K�?��}_Q�W�fײ 1i��ޏ��0�p�Dy�A_s�+���1�?ؘ�BKk�)����V�*$[�\���1�E��7����ۗ!�Y`�|���NNS�2ǭv��2�c��c���vw��n�Po�����u߼sIɓ�#��/��֕a�h��.$�^	!7�@������z��kx�3n�K����{X��pX�*�
�=��n��$uky���LY{��ᗯeC͋]����F��7<jWº�C��d�R��8�	�j�V���h�@�Ȝ��%d�3_Q��h@T-���B�K7\w;8���S�N���ޥ��=Rm�(��y�ݘP��Ԥ�mR�8������ߪi�ͩ�/�eJW1ӠQ�J�k`��L��_6��)#����V�9f�<"7�a�6�WW�#�wN�%Ѥ��4�l���+,!�+*����A�
R]�r�|l�c%6�գ���$,�(���Vn�&�h2
I�I$�t��iQ�w�憑�]�$In$Z�udܥ�!��Kf�6aF�P8�p�H,�D:92	r���w���t|q	 Չ ���m�/�\L�k.cR�fJ.H8�s1�`8H+��1�,eK�˹m���č�������	`[��]��ٔ�-c�L2�vʗ/%�܌ˍı2cWV�mn�Ӊ��2�*U��E��yvd��̸72�	# ]]�D�*dd�"�Dj�1�8�vˬLr۴�G�[$�ˡWB����;�]o��d����B��' �>�W��Q�s'�n������V��sW��Y�^,r	��Tو��W\����P[s��P��H�c���5'��D�W�]��:�&Z�~�f_vS!嘈�=��8���;^��&���Wt���w!а�ۃ�'7���<�:����Qhy��2��̽�)�y��*uپ��*����v�ҥ(]�����Vz�-�� &B�<���f��$�Z}���Ƽ��4F��}�� %�"c�=[�c�Ҙ��#��mx�H���|;a�eW���T���`hT�����	a�_ԫ�_B����-\���Z7����N�ugU�|rk����'P��߾�������߷*눃=�c��eor��U̙�W����w�=��[�ێ6���oP�z9>�&�6���ڂ����
l�6�ǲܻ��~��R� � !
��=���^f��&��P����������6Ò��R����`��y܊%������X�K�Zc\LCϧ~�\5�q�|��Ɏ�hi7z����t��tϢ�Bs���lp�Ab��w�{�)��7J(�o�9gt�;�қ��Dr�+��.o��UT�Z�P�Z|�����\oЇ�c˼<�g����j��{ҍJ�������Z&���Dv{;�ucG
��EQ���`�����a����@�*�.�ߥ�}z��Y�m��vҞM����K�ν8dw�w�[�x�j��16�m���v��Χ��ї\t�b�3c�t7w��A�'`�V,|ժ�����;�X5�}�kF���Ʀ=�z8�{���[]�V�D+(ATY�+�Vz��Ѓw����}Vʠj����rc�����o(��T^��4w'%~���靖���������Zy�X>�j�Տ�{����Ⴜ8R'�ڪ�/m��^k���j��G���K�=��^�n�n�|�ʈG���Ϲ����<k;����Pm*ݸ��g�e��u�L�ga�+�ָ���p��z�|�{��z��'qa&<����тn3MR�W���� �
"4=�f��C�ε��4����14�Ml�u�h�B�`�ĨtWa�f�QZ���ξt�ʏí��r/�+���s�m����ݏR�$��싿W�}��pb���pO�v/Z��ۦ�\�^n��}vD�ֿ&�'�4��^�_f}|����sM�c�[LkOZ��w�Y�&4�Þ����}3+�g�ف�|�TYPp���}5/�:�>ѣ��ԫA����[Ǿ�4]�_����ZD���k�N?k%�ޖ�ềlE�杧���~���riI�Љ�-v��w<ڹ�^﵆&��q4C��X
7�	(a�����Ʉ�noeY�y7�KS��A>�6�>e�^.�w����FY��1?��N:O����gaQ5wdO5�M:k�<Md&�u�S-%���)���W��k®�n��}���яÎ5􆝻������t��S�BH��OZ�d6�'{��g�Ϧ��e֓��B5�M���w9�W�C�|��6��J��֜�{��g�>O��P �*��B�4��4����I�V>�Ih�0� �q�3�k��٫�ܶ�E>�G����G���u�����u�}Çq�Ev�j�r��pL�ᯟg;9�M��U�'Cs�KN�_c�z~�&kz�Xq�����J��H~*~�˖��d!���k��Q&��Ah��o�o�[\�9�:����CW)�����k7�m&E8����l��v٧�}�霐_sgi�p�[�]��sƳL������W�C���,W,���z��6G�?J�2Q�!�%�v�f�gX��\4Ɗ�\OԀ���&}�J�M?u{P���^u�R��;���Z��<~M��B��؞}�:���������Ux�{P�'�B�~������g��#_�H����*�X�O4jD&�X���7rӰ��MYz�I�'�ը��������q�Ě�a�擺��۶��5݈d�x�|lS�ק�njm��z���N�sF���ǽ��Z�����W%s���͡��կ!���Ϭ����yӪ����*!>M�q�oһ&�s�szLm���D.O15���L��x��N�	���Bз��Fܲ���u �W�(�kB��I�X�\��
Mg���8�ޙ��I�ﾪ���7θ���_'�_&Sčb���߳5Z|����߾�}�;&������75��t���X�Ҹo���Kk�LM&?\>Mw�i3г�3=�s҈���5�uԎ�#;�u�{X�]�H�X�����J�x�ZW�*���t���������{f5��6v����Dy}��Ue���[���<qО7&:�7�ڶ���l;vs���m��%���~��o;]�f�u;�.�F���2��4�5/���\��������C���̋Ö��K�wr7���m����*����.��]�["�T:n
��v�i��lZ���+��\eX��X�&�L�����m٩���u�<�yڣ�d�h*˼d�<��>���}G���M�2�8���t��Yq[ـ.f�6U6(�j�[���Xh�[w�kRf��sQ�z�۽i�?{9a�e���7y&%&X-\��h�ad5r�Ym����À4$-�AYe�-ֶ��+h�a{��1���1(*e�IY��T2��i̬���|!�M[�B)����i�w2��<�CAb�-��/�0/sj,�;Rք�;��-����R��0"@�v٘kM��E&�R5m�I�	��%�-[�w	VʉKV%Ԋ�.0�d���Q�21���j72%c�[qȐ̙Y���̒햲�NZ�lVr�!i��vF�-̘�նՂ6��0-Rd#�Tq�qE��q�V1#�����ԁ�fE�j��(G.���Fግ�D�Ɇ+6��.Z����Q�L��sߵǳ�4ߞd�� �.���U_7�N�u�7�$-v�C���s\~���	��ƢkP-*\�׾��5�oiz�ϓ��Y>q6�R
_ܰ�Ď���Vhz�d14����W{"C!ǯ���Y�\lWӽ�ֶ�V�P}��~�(h�ѣx�ma�~ܧH���V���5ni�L{{ѿ�c_Hh�[| ��^��u��(��*}5� �H�Pp�����w1��Sյ������5���������ps��p߇�~J�\�x�ƫ�{iC��c��I���fK���7Ӱ����L��
aF��Գ����*�{�[��B'�A�1�}pӷ9)�/\��Vi8՚���f�uķ����܏x��tV��5N��� ]�'v{{�91�}�����F�O�ϽϽ�t�@ǯ�m�_\4��^߹��G������/�M���&�"��s!�ʝ�܆�p�˝L쭣5�:���nM�:�E��7��n<�٣:��s��[cM�zWa�	��ݺ�Mo=�i7��DP�Hl(T+�O�@���K�c���-$���?}U��}x����:�4|��i�5_6���k�陸i��Q��Y����i��bP�b���Nͷ�J|����}���G]&�N�M�u'�o�{nOsu�������^]y,��6�����z�'d=s��\kN52T������ۛ:��K~~c\M�jswD��a�枱��쇏Lw�Z�;*��up����%�kr��H|��{��<���k�f��.�[!�����;-<M��K�����J���|\R�%V����ۭż�H�
�/�_W��j�Cڵ��a�m}��o����s_��Z���KB�t�x��Z�=�:3���z�m")sv�Bg|s��]��?jnJ�vg>潛S����=�Xxu>��ʫB�^��A�zT���J������0O&6&�s5���m�E毎�;m��s�����q�Y����u8��;����?4y4�����GK�s����G�Z�HDϧ�|�8V���N3=����Yj�]*�=(<-sdk�����}�a�����?�V����9ڄ�Y���m�BI�����~�,֊"P�(h���1��ݿ���̼׮�i��3!������n��|��?16�5cV�ݞ���>u�tL1Hu��)
�4x$ON������ʫB4j
�>C���|����Z�,4�r�Ǧ�n4i��|�����}��[�,�i�s%4���N{��F��$�^��T��?Q�]NR���5�L
��0`�qQ�)����}Y��r��S���p#�$sK,��S/��u�u�;';�=@�#$)���Kߌ�O�Ps�׻_�~J��\��^�~����m�rH�я�5�_{B1HZ4���'�ef�T��Ɛ\M"��M?5��r�:����q�f�=p�|�=e��|��j%��[���M�:�����Hi1�:H�4�ܨO�19��wZ8hc�'�Hj�?xR>ճ ���kzo�k=j��.�.��7P���i��6���4�%�Nsy��k_}�U{q"�o�h�G�%CƠ��l�"Q^F:�B�5mxU��	hq���}��ӫ����]Nr{7u�s��Z�{ o%�6�:=	��tt��{��;��Z�%�rv�n/��z���v�����
X`�	u��J(��MVx�+Z������׻��S��r��>�u�^>J��2x8Aj�G��e�|�y5ٶ��S�.���Y[q;z�m��]LNr���^h��ۆ��d���1�\�5\����Rq���u ���&K�7���NbJY:��-�ǣ�Z��K�g]Z���W:vs�:���V��o����Ҷ6�M��ɷ�MJֻ��~w^?�?'�m�F��ֽܲC����_��&�I�����B�Kď�f��6��-̝w�x����D 4��I~�o\jrB؋lt�~u��5~ܖy����HD���.v��}����C��8�B�}u�۷���,��]|�_�����c�CO��}���� ��\tl���pKU�6v�V���k��g�jK��>���W��G��bc7(�5�j;t�Fs��� �����:>�~���`�^�Km�.��L�V>��n%D`���zn�޵��0�"�:>��u��L����ˆ_�����1�-�z�q�='l5���)���K�����Ë�%AF�Sf��@����}���I]k"�U�Hw�?{Y��a�S�����1T�Hj�5��-�����«����QtY�#�K>W(���7k����c��jn��ak8\|s9��kW(+���}�����4��ؿr|�;�I�̟8�vѯ��y�@��l@k�Ǻ:�4V�
�:Y�G���V)�Myf�#�>/���N�V
j��\t魱��v9�o��d��i+O΄�5f�I��+����q��Cᦽ�X&�<��r_������xv�=�y#�Bj
��i�ɭ�w��ɷI����q��s�čp�����?!�֢f}tc��[��]��w�|��y�q�1�ZCI��=ߺW�b�mnQ<��RZP[�XƱ�� ٣�JM�8rc�Y�L��>֮�[��,��q
<��{���s�K�m��\\�u�{�qq�M�"��qP�o.�Q�����Prf1]ENhi��}�$���mr�>]��*c��ӝIt85�6�����u�ǸX�������"�6}e9&�H������ڊ7��N�8��Y��D>�/)�fC�q�]�t�Y�˃�tr��8����%+Mߔ]S�RN���u�P�b)��Ք�'���wy��:���v'O�&��n)�J�Fh��G�G�� z^�j��[ƙ�A���2pg�"�%;˨��V.6�:��q멛ك���r�~#�^�Vmb��q�k%JKV�D�0��w����Y���t#�Q�dO&Pzp��-��e���ȱ�,����	�����6�C��w�.]ܱH�J����E-�2�[��6�q�����B7	�E��r�rQ��E��2�ja,�Y%e�(dV7d-����S.]d��mb+p�sr��� D�L�.����da.]��(�Bf�֑	m7R�>�h�A���>s�tUP4�X����u$"W�+������;�g�*�;��}�V%����yr�kH]ʓ�����\�Y����5��'��U��5/fZjC�C�Ci�m���沑�*��E�9Z>���O�]��>�kɧm�7�stZj��S���m�ݜus^�����ۯ��m"˞H���}���]zF�[k���� �R����9�/�I{!�4��-����K��Gʻƈ^4x�*������;�u"j��_�NΧ�oj��rc�x�h�9�F5��:d�g;�����{�Pl9�������o�꯾���q�i知i&�!9�{Tu۴��\č~q��S��{ �������1��+���k%|���Ms�ݡ�s�)��汻��{;�U�O&=K,Lh�g���'q��'��ߖ����Pߦ;�-m���j�^bc���f{�U���5+ύ��vZm*��h�W��6����|�rWw�b/p�����~����>1Ab�B��B���c���N�o�!�X`,�֑},�&�Lmw�7y����<��UU}\�~��~���\�|�m�DK�ϻ��qz�������u	�SLG����y�O8�9p7�������kڣi�c�t8(�a�Xkզ�Gs���}N\+^W��}�N��ihY��r��2q�:�,�K2|k��f��-�1�S���R�-��~N�(m�#��Ѭ���9���m���hs�P�`���wc(�͑�[6E߾����;��0�Z��7�����Q}C�ƕ�#W���X��Gq&ܛ~mU��r�^��9�C�o�O7Ho�5�"��8^���?�u�t�$Fxni�W�0���U8G��s&�MY���%_R.�+�r=v���B�Nd)�u�C�l���o+���n�tr�� .��S�{���>�~����ǡ�N˼b������?�֮Zܾ�j?����r��Ȏ�v�Fq~qp�����uϔ�!���Ԩ�f�$�9���X�d�K��5���:�%}�����3��lvT���u�z�:����րG�ˆc]������p3݋x^����o�z��ma�����rN�}U�x�`��7��e�����og��~����X�Y��o�YC���.62H�+��u��9_(t�u�)�<���vx�����Q�Ĝ���
�f�P�Ѫ�8�g>)����zp�d�ˬ��\�z8<"��z�w���凁e���۫��(�����r���Տ�[�^)�V�93"�5���UU3�k_�u�����h~�ҵn���Jv��Z^1T�� ���d��{mQ�A���q���٫c�͕E���w���]�-��}�M}����z�"����N1�O����Rj��¯�3#= ���[^�]�����<�b�v���8k�ѓU���IWc�G��`�f>�;�����q���&'� ���<nc`�������ސ���e�ڏ"1�2�����w��VY1vg�G�i��EuyD��9Ӧ��GF��K�:N�q��P�¯eǧjY-_1�F�w&R���wϖ��*�%X�e��'�e�g�p��gIݘN�wSbE߾���3�}��h>_*�a�U�����^�� 94�[˸[`����<(�@�\�Y����#C۴��ioM��*Ѣ���F��Y���_VH'����mR
V��9�//��t��i6p�W�:�
�K�~V+w����3�R:�D	˞�O�>{,�WmF�����}U؏�վ�3��w+�`>��?z��Zϳ*uzO�CV��3C���j�>�/�@[������"��K��O1��G$���Nn�>�b���q����'	�G���l�2��wȟ�*���<H�y��T��x�+#vwks�؉��I��y�;8@�&�Ѯf�{||����ޖy���6�Q�<�N�k.=�bf:�>�Kf���c��_>�%-�����5�PwC-��f㭫Վ�2���RhFȧ���;{Gls<�=aa6�14����*x��/4V�]�Ďq]�i����n��uee����7b��a�q[f��GT��sj�*W!Wt@Õ-f1ڳ���r��N�><uj�;��QK3�������Y$�:�_`�95���|�Z��6�|�v��I�c�2 �ݭ`�� �v�a��\�L{u2�T�GEMぜ�9��+L�`�8�
�OHLu�R�����i�'Zt��p�2P�A��Y3;[��P��:���BB��o72�3C�;��3'j0�2��ͩB��'�)�Md}y�,�ƨ&r�]�δ*�nm+i�a��"zzX�*��S+;��2bQAs>�MV���e��sEN��W1-}���;w=&9l�Ƒ��A�(�H��m����o&8�������L���(�̺�c��V�,�.�%�!.���%���Q,�WcifBP��AYR6�w�Zr�yq�����Վ\�@a$%J��K�_�����׏�smt�v�_E��#������Q�g��L��1H>1h����tF�̩\�M5�ݪݦYc<��y0h$y���r��f�c�P�Ӑ^�f������#�{�/ړ"b�Xi7�8*D�U��`W�K��$�+VgIu1�P���׷*��v��}�f\��LI;�uX;D����e���ݻ��o�4��G��}UZH�ſ϶Ǽ���{�f�_��z�2�����D��ӈ&:�m+ͷe��L-lQ�S{��5�����֫���ڏ��wj�`�q���Ѻ�>��� ��ZPr,�/ۙ�$͓���vL�����$�V&���a&�د{�]�yb+��J�hP,N�Ei�v�Y�6b�5�Bwq�/�˹�q@g���UjԆ5�gb&����|if�w�.�5`��[i�~�r|y���T3>��3î�9WM�����c�;S+P}���<�y��j��GwW�~
���26%�7�4->�^g��"9(��	�Ͳ�y��>�`��l�4>�t�VvI��l.����}�m�?	���|��q��k�$O�R]N��n���մ�	R̡���BVX��#�D̶zE{C�<e=n�G?��ۿ�Z�>�����K�i>:	��{Ź1E*�Mfi��������"�������||)ž��U�<���Ėޞh�{9g(��I7	}�u�Dv,M�.fN�}UU�O?˰7��/���y}�����s����x��Q��7@8��[�q�
e���^3�6o�D�-_��FVM��i`�vT�vV$��<�:w+h�j�k0U�#��]ww��=������&3L�齏�E��dq��"�6��)�0��}]@�x^�Ǔg*���W��py�+*�˺	|��?�_W�4��a��cs���c�J���b��eba��9��Gj��N!3��LGY�Q��k
�}�E��o|i��G��<bmbױ�I֏+�X�ՐCxm�\o�i{��uN�~݄�hX�S<�����^9��@7E�G��Z��{l�ҵF�%.�r�����l���ҷ���ǪPE6����?W�| q�?X��)��.ՙ�?v�U�\�y/C�ߖԉ����&��N�����8���w8{*�o	Nݣ�z�����/�&���)������+N`�L�����\�to����ݥ��8V�N�z���%ܬ�:Ռ�y��F����=���ө�����5����z�J��Y�\>�cތ�B)��,�3.���W���4|�~X�����7����/P��CAS��n����ty�;:�!�X��P���-��{.��O-!��.���E)��"�A���8��{̓8u��b�s��<l]2ו�wy�ۯݵ�-��m�t�"�v��ߪ������@�^�z��X։����ŵ'�ϧuh��k7U�(|�?k�Y��	r����m+.ߺ���k8ww�;�S�^J9�уi^u���#5�.R����#����X֍@��t?�'3��=/�ч���[��mc�DZ��钶�Է�k�
Br�A���ˮ�ڟ�����N~�+ `Z�'5����dbKU��ٓ�m��r[oo�55��zԫƫz�4����|�x����v��=Ge�WbwJ��+8�<�)���OK��U��1����C�n������0n�/��=��s���F�NqJoq���C�OY77�L�p(��h���9�����!�
A�%�bD�;A���:���QXy�t-�ʏe@�>��n�q{�ss8T�1��,���	��K��U��gAJ-|����(�Psume��+n%\8��Xٴ0�v7s��;r]uh�Ȕ��zs���:8�[F.wa]�.��K��O*G)u:�&�|la]�z�VVQ��RP��X���
YU�1�*���P ���X�[�.�ZA�`�0(,6qS,]�XI5Y 
��1�lR#�Ϛ�Zu@�:xV')Ϧ���"�X��4A��du�!-�f��h]cvi�h�镔Z�2�`�2[�̓*}�Z4�U ��L��+f�g-e��*��1!�&}�P�,1J�<$�9���܎�7���"����@*ܐ���cv&8䨃#�v�2�r�"Չ���ڌ2.1&F���j4��J�-�/��idČ��%�"��A�I1��V2���.����.�i\�n-�Զ�L��Dr1�̲�[��PtJ($k/|���;U��>Z�6:4F_U��ٻ�5=��3�b\��B��i7����72�R�O��Lg�Us{2ؙ&�xs���Ժ���da����Mw��'|��I����V&�
�W��v�":#�}EW���c�ʳX�����I����Ӡ�=[��<k륁���J��xW�>�۝q���'.�^���}�F_��O� pb��}�}���o���V=������蘙�Ys��z��sA�QϮ�ޓ|�X~r.xOS�Qz�֖$x�W!�g>�;�%�4|n����첫^Ж�z>���y�w�O��(~�۪��
�6����ِ\��|L��MS���cj|m-.�9���a�����C�4��c+�t_����M+~���^�]���	�ñq�n�z\+��X�Un#���a�fo��u0�n�z�[-�QwBe١kےċ`w�j�Fb���۝�t�ڭ��p�;O��ya����͚V��<~�Z6u]�O�6�gd���yzt�/v�Ԙ��:I�I[�g_�V-΃�㓿W���a�:�^���Iv�z�7���+�]ک��|���_����e���zϴRA� �C۽k]f�<°�n��u����p��.������K��C�$�vRl�1-���^a���@[\��x6�yxI��;$,4W:�=Q�a׽��d=���^������[X��J#x��>S�Yk�}��<'?e�=�ϳ�R���ھӜ/64}0d&1��.⟲��%���o��������k�s��Mnoe�7&f�=.}u�e�:��*ݲ+�\O�^G���Xb��T&����<G����<��R��
S�)ڬ�;qA':�zͱo�d�49v;.�⺠Z��&��䁅��D V�>�c�����a��7S��J� ��ˬ�h���6�ҷؽ)�1��Q�GŚ���Z���>|��S&�T���h�\{˔%�ۿ�O)<6_w�q�K���w�H���nj�5��+�ݡ�N�����YҐ��K��7�j��]�&`L�K�{��kw��cݾ,���)� �z�ٻff�.��$4�KvB������ϙ��ź��0*�^����8��������9X"+�A��zg����`�M���|�S�D���n�ٷ�e���5���'��p٧J���l�Y��Ռ]a��{�GZ�c�1�u���puf�{�G�3�4��s�P����|��P���Ъ[�O*�j�w$5��׋=����;X���d�󐌨ɇ���={�P\�;�q.�X��Z��um�eE�}G*hp�qvd�w�����HY�iʛ��d�y���x�=U���zǻ8���"T��J�״����*yʸ��>�&���:y���l�Z��1��6D���G][�����+����dVI��f�Z2��w"�	��g��f����Ŋf�ة��]��v�b��Cp�¸=�ArlzX]�"T�~�[��d��v��\pR�k3f���Ͻ�y�����ԑ�u7��Wz�5��er������}Ҋh�z$Յ��fr�.o��U��}Am���Y�&禳F�����w6�`ӂ���w�u��W~ڹ���F>*���
�9�z�tP�����=rV^�����ױb�V���6p��
!�bC/�����������ݴ�ȫ�H��nKh$v�*v;
�^o`=�<�κ#V��+u�0D:���]�H��q.l�5�pp�0����J.	oR���Ё��.��#NUѶ4$s=Z0�"z���9S�I��27Qm����U�vsX�W���imv꫌��@��N��W&y�Ͱa礌q�ari1�Sf	�$��y&Z�)�U��ѫ��IyZ�Mn�d�C91h�_�Э�wH�����i۵����F/F�T�ѻ[7]z(D�p�E`Ăv�e��2^X�ƪLVIq������\9*���15$f�@��L��;��H+<�ƪ`�6�7X"��L��3t��Z�� x�:�ʻ	@�bBlPF�Veʴ.�LN��H���,jSfK��1�(Z���%ee
����!e�'j����ws�(7��c��\q�d��%*�r�lRa�)�%��2H5o2�o2\��B1X��^d��F,Y���J��U�bK������%��RL`�5$�0dX�ZY",X)*��2�Jd��4�-�"�ՍHː��d"�"4�I����%HJZE#MʉlY���˙�����#������aby�]��$OJ{[��{�q��X�5Ϡ���{]ق���V^	�����L��(�Z��Ƅ�W��-�z���¾ek;� ��V�;�i�R���@W,d���*w�$�����Xm틦��sq�����8	Xz��Mǜ��C-��`��V?9��Z5����M�[���x{�[c�m��4�+�Ǉ���&l��� ��؋��ݗ0�l����D�+�x7}~�پ<2{�E��=s�g�['�u��� �U|po,�s�*Y=ԟ*T�����ɓ�`g�+ܭMV!�}�~V}�\���j��9�L�b�V��U)�ܹ��f{ϙ���}�X�a���<���nOi����'��[���|���/Ҍ����9�������ESݥ�n�&>�l��gf��d�F���r�h���7`�X}��1�]m�יx����X�:瓖#�IK(?B˗�Y�Kʪ�8oz�<f�ܶg�f�Q��fx���s�>��|��B��1W�iP7a _�n�q����������<��/�x8��Ɍuѕ�k<v^��`�$<�ZC���l[�Dx�OMN!axu��p�4ņ8!zϯ+��7��<�n��.�_�A��p�pѯ�����{�
g���SA���n�J�s��S���Ӟc ��ص�M¡�|�;��B���n�k�0XUŒ-an���b��C&�P��)��]H���Bv���lR��û�6�O<��N����[���Q)=|#Y�����$=m��g
��OH�L��K^>�e����a�6Ԛ8��Yoi�{��_[�����m�7�����������M����'V���m�oI2�}j��A��Yd�����˗;u�����޶M�76��{�z[�x8�l}w��|���EH����2�n�]�
����N��b�x�J��=���lJ(�y� �g����`�IC�5���x�yԑu*z��{z���U�T����6=e�0��o<:{����Wx�1�
7oM�k:��F8��!�0���^j
��ir��o+�p��	�q%^3�Ʊ%e�y쑾4��b����oc��\�ʓ��{����Ħ&ߠ��8P��Θ�)��K���Wyڔqȟc�wgĴIβ������қ�}�lfA�h�ے�<~�R=��~~�/.�u..�a�n�7��_���N*.v�f���*'���Y"�Nq�Ƅ�y��j��!w�'iϽQ_vXJYZi&rw�pw�ŗl�zy1��� @4.�
8��P̻�U�B������|�����9��H�|�?L`o���7>�)�r�w�&F�8a�i��X�0�kq�l�������j'�RN��Ex�۞��؄����:&\�ɧ{�{�ǽ��B�D�}�y���i����z����R�����-�ĽK���թV�r�3�"��Ԝ����u�����`Y��uׅ%a)�Wk���X:��0̐��¸�c�+�{�͞��ᨫ�g��k2�+]c����6>h�M��$�W�0f��'�������A_(����f�]ee�O�K�=ǰH�E�2����}F�����8(q��m�ioVJ2�x�����[�8o�a��t�˅
�x��ەѝw��J��z4\�Ulf�ڔw@�.|�WH.ܽ�s���MsI�S8�#F`��勊X����wq�aj�����R�ZNŘ�0��so7Fl���u���E�9u�n��O��4�6�R��70�M��ff�T��Z�n+�.�L3O>=.�g�Ȱ��x�b������]5`[(����L*Q��QW-FF*�]�m��ypѼ�YJÏR�L����h j]��f]�/-��k���P5g(�S"�`j�̫��@��@��R¼81"�#IV��m'�(�tX��uC]"u�tj�8��F�R�TeH�D��˨yuh)s%܂��5��1"4��d�V*�ˊF�0m�R�Z�]�"Ĕ8%����e٘KH�bB䪒
�Fɍ䅷l�r��d���L`cX%��%8��.��.��Y�E�c	�VYwR�ne��KE*h����	?�����}	�^��G���VmwtZ�.W߾��׳W�(2z)u9�%jvq�������S*(�iyyj'켺`��Fu4���������β�i��Ff��礉{3|}3iɌ��	��?{K��hV��Ƭ�W����@���c/�����v�;�o8�ms�k�4!pP�@C����l/��؋�f�����ĘiS�=$J�=L�α+gT��'z����h���ߏ1�z"N�T�y޿1i�Y.�[d������t��bw]���s2{,+���G����v��C�|+®�S�{G\ɴP�Uު�W�4~��v�u�7N0���I�������6�d�Q��爺�ٱz��N��7�`	�ʜZ�K��j9�r7am�����D�����m-/7uW${-��(��?8x]����=�W��^ib�g0P�C����Kr`B�{]1KN$�	qb�.0�{�J���^�^u�#�,�|��Xɫ��[���.�m;�3�=ޝ&�߻�=�a�|"=rd�U��7����#]���9�k��0v{w,�.@�r��-��Ѯ�cY�r�48�����M�qv��
mq4��j��v�j��tщ�5��+��[��Pb嶓1��0�'7=��K~S)M��H��,ݚ�	�P��1V#y�qa#w���B�#��싅�^�ݎIRX����K=�*W���b~|�}�
y�5u��I���el��댹����n�F�[�z/q�G%M O[��S3;5�����vA����r��2{J�=@KVt��K���혧a��
\�/{<��d�X��g�� *=ѵ�Q��m� el]�.�OpųS]���1�4$��;��'��܀�;��8s�:�\�:u��X#�/Z�>$�gr�[��	x�<��fA�)��������/�鷁=/��v:��[�����z�7�׻z���O�9wD�gNÅ��f\����l��x��
��]!�/�Ez��;�%݋�����ɯ%�1;� �:yӽ� .a�1��Nw��X��=7�yI����ˮU2����6:>}S��;^Pc%ղ{��jl/�J�B����uS��,gXz��怮�8�w�l�P*#�p�>v�1�^���=�Tf���c�+�7]h��ϻł� �s�6���\ݯ
�w|��o� �<k�h���v��Y�=zݸ�Oe���P�e��&l�[e�?[s�Ŝ������Qk˭���}��d+VV��۞a̫S�������f@i�il�*W�D�[�
��ŜO�w�qڍ]�!u���z;���XX��&��$��"��e�b%�$����k��ز�/S������%��유����r;�a�S�_�p{�A]b^U/��#|��YfhJR���W�Y�^?>���"���u䢏ӵ�h�)��k�X�Z1gm��*2�,e�noc��{|�S�0�v������k�N���2���za|�ik�F}�6�u5�1�V��:�����O�ȟ���So:(B��P�|P��#��Eu&��O�_ek9p=��ɯ�N��_!�m�/z��\�����v�1;�E�Z��]������p̮����U��XC��ɶ��]�w�~6j2u��{ϥ��_������W3�q5x�����!�'8_9�p�(*V�ev��z��Kl�z�Y�|v��vp�G�vM�(s�TۘfrYf��]^1S�6�і�C��⡥x�7}�h���јg86�t���!=N�hpcj�7�GP9l�>�O��)�5R��Ut울G�Y�=��\��/�%*0V �]#�u�ק�=l��.�Y�4�';��R]}��I�Y���pk�+�!��w[��s�&�$��iMdX=���b+e���i�2��m-���:��3��J�d�;2��b�wef]I�!��02i�\��NGR�s!�x�/q�X�@��v+�M��:L%K���NCD�Ӊ�wwJ/��?��GM�k�9�7*I(T�l`��A!QE���u�eE�^0�y�]�c�f>)5#ir[j#kr���w�cja�e�Yd��ALUX���&-�Լ.�9q-�����I���Dl���qYa����K.��2B%��i,���K�U��n��vܰne�KY#�J�ʘe�W-�r\#-��m��#Xҳ,��C%�f0����fY.ĸE �%.\����ń�%��oz�'V_4��3K ���A������3s�z�i?p��~��|N�e��ע�=!6I�"E�#��<���ʱxW�r�^�|�\�?&
C��z�p�/��[�N��ٴ�Y��tkŦ_3t�s]���-�_^��k��ok3i�Q���x��z�P��/��
*���P�v�v��{{_Z��ź��C{Z*��+=��Q�11�z�Z�0����iϏ<�VI�;[m%��|��=H2����Z":��E���<�wm}�ҝ1�W]:`�(��Y �}3����U]opܙ5���٭Rқ�~����;�i�G��]�;�.����������9����P�>���h�.֗s}��b�
*��H8�{;n[��!ݥ�.G�_{�=-�7P&�a�=�F�虲��Un��IezƘ��Zє&�^\\W1�����V��M��-o�8��L��W�Dn�s'�<�M���S�e�5;Y��޵��;C}�m�9_U���Ɲ�.΁������OEn��5l�^�RH*��]a�;����;΍�#s.h���{ee��4g�y��@Wxe��(��NpU��*�eMEK�����*�A��b��<�]|��<�����O[�BkY�=��f���w$]h�3u��������8vE���=�֖=�~!
3,̝�n[�:����"Ji��v��mz�*��'�1�Y='[�k�*{�8�yCƒ�^;.U{>��H�W�B|��o��N �=-�\�~|�R�V ����6L���X�z�㵣յ*��v׬Y����^p=��Ҏ"��%�ر7}͙8L�@��w�uf�ۭ������o7<`^�¶�ux����T<�`��Rl���w�%;E��H/�?6l���t���<��
�]=��������DO�k��+�~�R�t)#f�VI���>�'��*���n6]�ĴEswHK����W���J�����/��E��ӎ��7{N�&;:S����L*l���g������sL*)DT�{�~��I�Y��J�����������ʄ��q�XW���E[���(1��L�H��W^QI$d.�P|�������޺Q�[�(�P��4^ۺ�J��M�SPم�^�Qu�RTOn�:Pl:�T��d��]9#�7@�w�p��7Y����^�����ؘ�'�ʆz�z�w�[�l��mG�v#�s�Qg��j�u5�\���u�;�^F��@o���"~ng�k�sfW���P~�>��;�+}Խ�!e����	+`����b��:��E���<�oZ�����x�ta�U��d��1�\V|Iu�~Åp��Q��]��ֆ���.��1��m@P��i(��q�c���2��v{n��piō�8�2ƚ"�����ݞ�9T=iE^�di�c]pOB��;S��6����3�L	�e޼��޿��\�{nժ�;�̦���V�@�f�N��:�e�x���귮Nz�`��F���z�dȟ��o{��ޑ�܏�[��4�S�E���Ub�\�S���GH .��\���[Z��vQ����/�CVĪ��	�NIJ��z�i��UϞΕ���;:�Z�o �����k�U�:��B�?��UU��AUT����ʠ�P<�R�b���P�|�Q�0(��t�m����������tUQH�U@"P�fY�t�!�a�h"���-���,�i�ޛ�b ���&ٌ��+m��_�j���J�-n8��p��	���Ƞczlɩ|�� �xQe���q�.�(*��&���=�uu�� ������~�ꢨ�qFD���5�s��@�����OK?m����r���[^h�_���_0<���� �a���j	n�����07@�L��RՂ��� �;kt#m��;���mÝ^밽+̃��W*(*�3��֛�=��	� �e�`�CFa$�ia�R��1iZ�zX�8�N�Cど�@����IRpm��a��>�pJ��� ��@�L36�W�ha�}G�4=����&����4@�kGJ2��=ɶ�i�����Թ���J�- ��?Oe;�s/����Y7���ǣ �6�b����'���sD@�y#2���2?#e�,�9T�����O<�;@UP,ʽ���L=�;�RQw�pȚT<܌K5,>����"���Ed��hթ7P'�d;f ���b�c��������w�����A��������Zĥ<KX�*��*
�f�;x�ǆb�N(��3���w@bz~���4�l�hpǠw�A9�p�Q��*M�Z�k��k"y'���ܕ�p�b}�yDAT���m���O�
+����I=H��_K�Y�S�螆{�>���D�M��jm^�{&$n-R��~B*��t��G����������	<���ʦ.z��{]�D@��q,�<x���u�]2!�P�Fn��h��q�1�zpȰ`-ؖ�P��"���nA�<�W���ǖ�TC��M��ˇWU�˴\����}^u������Jݮ�u����w$S�	�MgP