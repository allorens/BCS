BZh91AY&SY��.��|߀`q���"� ����bX `                                      `      :  �  �    ��4  P �4�      (�  ���        �            (                   �    U(>�Ӟ�D��d {��&�p 8�;tUC�2ɠ�X�h� ʁ�$��9�vh 	U�   Jf�rÓB�r� s@
e��P��5�f��4WW��yU �� �I��q�*8�T�ʽ��y5��. @P�  �        ��^6��:�0k�IU������ qꤱ�)d��h\�I\�8��7 �R��q9T��S���  t����e�&�R�� �
,���һo=�S�h�ڤ9�r�%C�� <��й�s5B�ҮZ�sd��W&*R� @�  �    P  �=ʄ��y3Z\�K�C�.Mw�
��;� �U;��-�6���.,Eq�DAr���R�b=�b�p  �x�	t�`l� `  {�94H�5C �� p��=�@5Gs    <t� ��        �� T0 .�����@�2d�u{� �C�u��� (�t  ,��@z{� �#��`r r9 �C�� �@��2@p (  �       �    $ ����@;�(p���t@1�w �	�2 � �x    Fv p  =��C�`=�C �� �l @�F^�>    �~CI���2b`& F�2a20�~L�JJ��      
J��O���#B�)��S4�S���B'�U(�hhbd��� �4��CQ��R� h   � �D�
�$�'��&��	�����=�O��_QIۯWN;���ӷ}|w�g����E%]����IWY(=�{�1)*������|�����3̏�QIV�>6�GJJJ�-w��"������|���F����T�2��U'���d��2b��5A<�!�K��夹iW-A�U\�Z-I��-Ur�9j�����\�Z#�$��G-!�.�Tr�\�W,+��r��YC��NY#���$�r��W-Ur�-!�%rʯ+(r�3(�9i-�"�VEGV�.�*'V���i2T9j��bH�S���h�}/��������W*ؘ7ú�ˇEk�|1=���gS��f���*���	9�T搁�3��{m�w_u�e����gN���%U:Mƀ�|��u���eU�㣂�=,��Y���)��'(�^���St���v��Z��D���gX14�Ct��j� �,]�;�\P��q��BU7�Z'n��w\�e�g �����er��Twk�[�7�Ǯ���;�r��rq�+iI��9ȭ?]܇�g!4+��	�s{�<���n��5_uW����<Y��vko�ir �.�PE�D����DJ���S��a���rwr���bLJLsI��8y��X�,�PG�l���Dwcv+�ob�6����N+AW'.ږ��ts��[�l���dn��t(SXX�u�i��98��y�Sp�['@�f�g��v�~�׻׆0w*lv��1=M7�a8@\w+΃�gc����h��T��m�K��s���a4`��[qkc_F���Ƀm���n���p��������H&����]�nn�+�k������s3��Ҋ;����8sE���ฑ��y�BM��8�E��QGu�eJ��^��#��OR����d�Ӵż�AP;Q��-圲j	��`��Q�vL=d%�N]�phG�M�w����S�wF�幃i�����@�sd� g;�Y-t�6d��#}��2��}�z�uSpm� � �n�A�wH�-��h��č�����D�i�V��k�3�{<{c35���>�n^��`���0�J�[�)]�-������ i+�.VΟ��5gv��1.��D�/#Y��"�7��F�i�sw&N��ܝ\)�@�'�ۂ�l�3��.<_Gw�wj���k#��Z�-�/"�Ɱ��[�S��������=�ೞ��Y1�+��9�s�'�^�c��.�x`عц�թf7��|V[���d���܍��pw63aV��[�B�Mlɫ��d?	�f˺7p��౧����]�����L	[�Py���xᗚ8]�uF"�A�{���z)�;c�ȴ����#$���Ra�̆���:�{��Ԓqui-�7WD/spω�Jvb�������v.�\VU�;jp�#�ܱVR8n���
�\"�.��-��ݚuguY�a�MX�}�ݽ���]�Y�u�[d����-��sxqΙ����~�S$p'����\����qbX�ݜ��]�d��)�f8��}1�u#뚳��$2�ѡ�*�lО>�'�z�T��%8�8�bl��A���۠U�Ψ0�>	9:�0S�;x�r�p�ֺ Բ����Ý�r��U���4o�ge��{;Z��2C��Qr�u���A�[�p����'��\��Jz�|Žy��p���ղ��/�f��\���'��0s[�T���|�\���h�a�UØy��	���
Kfh6��<�z7L�Ǭ���㉞�-X+p@ז|��vq�SU9��G;ɒ�e�&����Ӧ�3���
�Ι��Uw��b0���3ss\{�:�a}�DqM���%�l�ź�3tN�����r����*_.w#�e����5d�����w��#�O�2�o�jQ7�zƝk��Y�pv.g;��5+��Z�6��A�^�MB��r�{��=O���O<�q0c��hm�y���z�@���j�p�q����Y��ti��Y���M}{�_j���z{�$�zL�lAՓK���+e�M�+��n<�Ӛ��$M�7Y`�j<�V9pa@�� �#OY,Syo�E�1�q��qŋE���.�\�8`��vKx�r�-f���H��'u����}�IOg<�0��Y:on�#�B�8�>��v�C���!vYh,��euO�^�8N�C]1�ǜy��rۆ�y��0�O�c�_t윸#H��ssJ�fs]�X�sx�ܻ��4o�2�a!�U:4��X=��n9�]y"�>?N�9��jeqnz��cmD:H�˷B΄`黺5"���ޞPt�W^[)�@��JF�1@�1a7���u��Wndd�����T�=� 9�;��r���nw>��b=~�c��ģ	ʬ�h�(��N��$ҥ˫yڮ����Q�&T/Ю���y�B��-=^l�!ۧQ����E���1�Np9��f��7C U��ɧ�Xm)����9u3y�΀4���~\�1���ث������8n3��O8�v�sPi�uDw�찮�s*�ԭ��~��*����կ-�nj�gh��B=��@=ݳU\��;�!���|�ɥ�T�V7%`��f���wM�t�B.��yvk�v!�H;z��ˍ�2v�K���6k�d[��1�+��ϾC�\�O$D�r�:�Ȃ֜���.���]���% 9-�k�v�ԸŁ*V�ݬA�s3 ����7"�l���ԘF�ol)t� ������U�s"�g7�@Ya�Fr����{�X��lc�;	d�,݋��l֒ ہ�h��E�\q�)bl2�'���vU��:p+�isbG�Uˢ`O�ig��i�N�^F�}�n�8���#�f��z�,���<P**^u�ڄW����#�n�tZ:���ViW_L<��@˥@���D�2:�/��,u���K��q>���B7\}ր/�����J���dv���w���c���LB*���:�W~�c��v��yö�Gr���uC�w��Tg�
�ʗ����`5u��H��enq����j���p���^�=o[���m=��ҖYgq�w9N�W��	���ĵ��k�f�p�)��u4M/�ls�*�rG��ڐ:�(�t:`Տ��q ]�92e)�]��|��|��L�^\4��i�kM��,����xC� ;q����[�&�:���d��u<�Q�{p͎�Y��M�^O;E�%Pkvs�>�]�v���y�A��n%�q�˪������f���3��s��D*a7;&&a��jX�g9�Q��k<�w��� �s�I�1��Q��)�Un�����ƺ�V r�ʝ��oxh[�L�:�U-�.�	Ю.՚�V�\�'�`
M��%�ă٦j��	�L2^�z�����ά�d�B�Z�:&�I�4�����X+��"{��7S%s��[&k�F����F�N)
O83dͅ�C�4����+1EI�Y��4��U���vLK m|��m�����q���<5\�;�v��K*�<�knu��:-�'<��vu�����w�]Ok�_vp������!��$ ��$��Y��6��ױrɸ�*�H�L��}�lf�l�	�v�98ok/d���W�&�v�p}{N�	��ڀ��O�`�t-Ԉأ�d$���k�'1$�����6�p�A����Ŭ�Ǜ�
�~;�ҋ������k�'& ��زܳ7Ʀv��`Ɂ��x�xw��~}x�����C�׸ޱ�h7&�@��U/�4.�k���v;�$�i/a�%���lr{ٻ@���� ཚ�W�x�ּ� ��j�w�gT]��V���ۘ�7�L�Do.$�]��wA֋�(��<;�ɂ�/�-��Kpޖ��J������䊵ſ.Q#ъ匥Bv�,H5�2�4��'E��w��z��f��vŪo&�3�Aŝ�
,�ه��.ź�&�ҩ�>�ם͸��{x�VH��dZw�$a�g=1��H'��;�Wyfs&)m��L
�Eq��gB���ˉ$���a�!��!��c�bK�p�-�-l�Ⱦ���]b�N��� ��6�;!b�:��[!efv^�ؒۜ^�	���ּ!,jg��jB���Zu��% b��IA��틶ak	c��9t�;o#&�X:\��A�ټ����7�v�1��jov��V� �Kז�P's�.5��'��$c���:�s�m�ֽՃqǿX�6�ڶ1�h\b]�5L�h�B�0�۴��t�wHC���V�Uus�g5�M�[9I���d�ǻe�Y�[Z��e��W%�rX�	�f='n	���{�Q���C[�-�k�j�of��7�n�yggN�yMَf���WeM��(��ln��zf�
��s�b�GgSа�gt����ۧ���bɺWkP�-��{�ri2W�Ǉ�d���z�:��
M&Zq���`-[�gqi�gw�=��n�맾����8�*���<���� ����l��oj�cAmVwd�n�޴`ŪcÏE�װ�Z�X�Ysob\��@.h{��V�+8�+�@Z����ȡӐq�>�WIy�T8W�TWnoa'$!������;q�o���%�T9�l����Nܠ��aw��v񛃵��J�˸�m烺���ŝ���k���q��m5BuGh\�ō��f�e,G9ݱd�a�c�d1��-sx�&��	�WKK2�Ǩ�5�dZ���R��N2�y:�+��ۼ���ǝ� �=GHu�:��F�D��b�ҳaIh�ul�������yӵ+)Ȯ��G� ∘�(�}�p��������[��8�j�
:����T7%�q�oa��DOp�d����S�����3�,A��y�`��c ��ȝo9�Z��'[�wlaC�C�8��j:3�,���:ð�S���nnd?u�¨q�wN����4��wf���e��ޜr��IbX�w;���~�Ya.�׆��N#Z��Y3�ܣ�w&�qL�/ �d�Ǵ���1�s;,;��Ɏ�62w��}� /���P�w=g����x0�Pu��gy����;���3"�v�K���y���}ݧK�P��婗�9F��b}�'F�;T�cc9�:�	퓀�ɽ�v�N�*@�X��� �mNn���c�7�A�q|F�ϴ�o_8v^�Cd�B.�3�t�}%�T�d�Z�0bC����˹y��6�ݚ�+�K-��FӼ�$=���-8�;������c[�*��t�8v�t�[T�9�sE�)���^l�����3C:��;@X����<���UA|s�hˢAsCssyo@�7��F��u��;����b���cs��8>%��#��z�\����b��J	2� 	���]�g0�g�L�'D�*�ػ[�G^�׎�7�#���s4b��s���#�_@U3D��sAM.va��0Y[�xF�V3����-��9���κ֮;�� ye*�KB�ɡ�&=��H�NU�,+�,���P������W��<�'Ŋ�����臎�r�n�%�"�Nyb�m�&��61�������{����c���w;�Wl���t��b8xi|���]:���.n��	<�":�����<��"���M��%���U����9��� ��L��l�Ҭ�oV�s��x��2�v�Tw'N� �{�e��̦S�m	�k2%��B����c�ݸ:�F�On�wL�{C�5Gr�+g�(i�(ga�5�:����'��ǵr&�2�<�gv=B�B����x�uÂ19���NW@�ͧ�FS�[nTu�ΐ���'�Ͳ�(�%7_r�q\'�ta���{'f�)��`ӡb(\��Y�6-������ʓ�l���Zn�܁�{����v!3O,�����1!9�cLи)�ϊ�{M��\h�]8�� N��W#�dJ����ע!Jp�N��V	�`�FL�Mm�a����܂ť��;��X���ᆦ� �xRGocc@�Gj�����	S��9>��`��c�y���r��l׷��pU���.�nM��>���<�f�m����U*�����"].�h�.ˤ�&+8V�O�׫A��0H�̨w�a��:�@ݡ&p,m�;Յ]����10Kߟn�@�ٺ�g�L�K�xn�o�"&i��05���,�t!�旅*���;o>'8��v�_\|濶gQx�:4FwM�{I��bYnNON��J:�P2�7�;:��w#bd�sX.�Z��O�������5��d���8��̈́a����~�A��މ>��/�5�Ny8���vӖf����k��R1	��v��[��O"\�c�F��.hh7g&j�6.��:9�˂�r38:95Į�TI��걕e²{R�ѓR�lz�l���ʗ���K���]�t�a]H��;.��*��N�Ѽޚʌ���X��PZD�It�~s[Ůp&�K��f�y�<��:�D���3~휭�Z4Rsgx��7$���s'K'��9�Nǝ�Ќ'r����� \�NZ)����{�q`�?G��Wh�^����B�)4���٠7��SҚx�Nq+�7ˤn��]����n��$B���u�� Q��Ârf�,�\on\�n��oS���gu�i�MIr��t�^�"{�$1;]�'�gU+
SU��ɯ{�|\ �Rh��mZr'l��кn�H��{s��A�y{a�=����N�~;�ZQ��X6���bD�$��!%�2�{*��,㧶�(�U��Ku��w`���m��
��w�;�m��K�٪\�.Lf�ʬ��\�[!�4V�ݪo�-pq��C$��n�iX��bK:.mW�3O:�+��TCª�3b�hs�&���"V�,&��������դe�:����G
O>1\�z��'�ӣo>t���pZu�/xv8�>�������%��^���yn������q��Ӥ%��U�Ul��-�6*}z��ʸ�*lT�UF�-��6��8�+jV�Ƅm!8�V�M�[*��I��`8�ؓ�(ڨ8�b[)M���5+h�V���m*m��B�2��V�q���m�h���+h&¦�SaIM��6���lI6Q�ڮ4�A���UW ړd[*ڕ�+�U8�)��q�.56l��-�#��I��J�0��C����ک8�e8ʥl6!6T[J[V��&ɱ�QƇImE�*ڕ�$�$* H� RE	���2����:��IHR����\�.\��"��sQEɧYs������1��iͨ���nsu�R�?�!$$	'���WU��y�|�n�?})E_������<����O��1�����2T9>��<@��������Q������g���;���8���}�����i�y�z.��������zc��7�.`�����=�sݾה��\0�V��|���Ts���&V#�^��)#����$��6�[��/q[;�E�Y���9�����|,=�{������&���P����=G�5��B�ؗ|��{������tlq'=�L^�3�yOh�4�{Ɔ}a���'�I{ǻ�VF v�GZ=��j�U'��{8�����Vw�rp
��w����qYſ���W	8�7p{��{: �n��Ǯ�*�����1�gM���vr�T:�������s<5��꼎=x}V��8��s�9w���&z��2|k���d���o{{ݳ�3�07��������o��G��m;1�/#�,��3f��?_q��!����<h�f{�]��~P�\d ���,}���Ɓ��/-�Ľ\�sd,K�5精j̂U�;�
Ⱥ���<�n�_����������e�s{���-[��Et���3ܴX�p^�S�b]���s�r�"���P�Ojk��/�h�9��ˢ�㳳��g�����Y��Qˎor�|�7rz=�����4eX�� ҉[�4�����`�~�xT7���yt��������Kb�&绞N��A�`p���H�)c�b���w۠�`#|�W��}��|s~ۮ��7=k.?M��|VNz��=�;6�=yK�X�p�ݧy��jw�Ŕ�L}.�=E8��雗b�.zU�Sh{��R$��R�痽�Xw=�"����>�y��ӹ-����k'	�;ƍ�@�Sg%I�Z�V�:�}�>����|����3����8.sY��~�dU�FW���+��gw۴��m��rqNW��q��7�,,u�.���
Y4i��80C�r9=<2/uÓj.�����YGl��a�v�	=��RË�y�Y�r���w��<��~\l���ܳ��rʌ���6w�6S�5~z�G��e��ܮ\���d�L�|{M�����z��o�G�{��p��\�٥ִ�ݣ�@x����Aǆ}�8�#�P�|c�xV���B�8���ũ�Z�Wפ0��/S�yQ�|!�}6��{���sʐ|zN���� �p�d$0�OT/�M�W�-�!0t�O.>��>Ì�On�����ie�y�m�lP���i^l��^=ڟ@�ʷ�g?	c/�2�z����}��isxn��"�z�v@T�9i��nR��6]>��=�~���3��ή[��w�5h��O=�@��6��3{����p�A��ݳ�槤ó�>9�þ�ޘ�G�����VKH͒�7���7<�N�5z��qN���=�;�H\���#�Ђ3��$�w��_���&������Ɣ�%��k�9�;�p��cs��>ѓ<)Ѽ��b��9_�Ӱg2�NS�%�Cy~G��J~΄B�{�+����a�_)�Ԋ�j7����=�� �}	�M��X����X����u�f?���鑄��s��3����t��;�]��;{����!�c�<nY�=��^��`��G�����m^�^zi�^�i��:��p ���]�\<�^���B��b0��&����&��D�������9u�s��oBj�yNE4y�|~Wmh��ʌ�ٔ@F�����}��{�ݔ�^�Q:|w�p��l+Q�lݙ�E�-K�Tz�Mz��ܴ1#֐��1�N�q���J󞛾{]cH�n@{۷��7�ycf�mg���ʮ�w�f������Iޟ�d`�T��A����z��{�a���"��}�i��剿�I?
N��6po��{Erf�DE�{�*�ND@�ru���c�����y��y��N-�S^���3p깽�z�����%���fz������X�N�|��gt�#��l��E]O7��ɐۓ|��$�o]�	N��vϹroy�yr�<#�#y�$�
C�kU��pbvi���P�:���fZ	�zl��t.ŕnX��R��<���V%��xx3��˪�B�0׫;�~�/tTo�ӛz٣�
;}�����^^���S�L���hW��hzp.��28r��ꚾ}���V>皟��v.�=k�9�v�9{Y7�/�����J�����ޏJ��Qua���7�-���=��8�֊.C���v��,�6[�8��=|t��Ȩ�xEV.~�ђ�f�3��;��Y�V������{�g'��k��-;:<0]5��9�✓�_�菧��{1����U����,�����xn���x����4�Gb�k!ް����{��y�K'g��kO:4�>��=�h�G'���7���}龙����.i�sţ��N������6w��݉��i�Tw�����O�.\ߛ�M�#�/{o���iM��`����n��4;���{"�?��kމ���W��Qݗ���a�|k��[�p��wOYPW�?M��t.%/h���2�L9�z�R��o"#����gy+��]�f�нۋ��~�t���J�K=���'o��u�}����ݨ+��{�tM=��ֽ����o��j�<k���3ۺs�����aR].Q٤B<��ݏm���u\3���T�:��p�O���� L��y6Ϣ��i{g{�o�|����d	�>�l�.�q�����h�X�u��C�e���/{����H���C~޷{��ȕ]��=2�C~�D�	���Юg?`�v���������ղ5��K�� �|pn���mB��7s��ِй�w��i�߳V.yg�d��C O���Vpy�y�[��d��xg��}��6�T����{�4'��wٽ��լ��3�ov�tʄٖ�dk>=���_B�h����ٷ}�Y2E�9��?t8V=Y�r'�uX}{;t{޾�����azw�6�.��^A��W��3����9���3֝`su(e�� �@P��g�B�˘!�L�3^�m�sۊ�i���a�-���<Q'�F���O]|��w�D��޼/���'��{�c1�]gw�=��<*(!\:���^�Sun�(�8�[��1&�3�q�-����]� u�y�Qg{�ewx�"�(C�$��o<�ݗJ��T��1��������-��=$y ��9:d��w{LO�^��k}_�>���WWޏ�n��wqx�!��uo&7�{x��w��_>|�������3�1>ɐቩ����n�~W��,�����K�6��U�<���J���v���|<�}.n]�6�w]:�l����Z����+�������hnt�/s=�����D��q��1�4��N��7�9T��建������ʎz���s��%�,� ��ǃ�]�qwh�V���K䷹��y۝��E_�8!m���ۻ��.�}�ş:w���c�&��ۏƐx��Sܨ�2g�6�4B��J���p�I�kG�A�H7N��A��z�����n�JǇ�l}�U��=;���y��Pt�2w=<�|���ub,��HMyۻ�O93�O�������>>oL��%|2�)�A�(��]�8�F����:m����k���?FfJ��s���T���f���4�&���=���\ �z�;��4�9��ѶSsۏS��y�}����>W�u�.��QNE�K��2ø./�3�=s�KrFV��|}�F.�Ʀ�v3�3���+7g�Ӝ���E�J<�t�=���.�K���[�|%���$rq(��Tf��M�)���4zn���y��|����#��=V
CH��ּmN@0���,���2,/�D���/����j����GK��b��{� Cu�⫁z��n�����o�K��	���e~;x�M�#[\OJBd��?s�o�����ֳ]�}w�����Mc^6.����"p�H[�~���<��t�����;}���p�~{Ko����ۇދ�n'�W��F��A Uڧ���@|�{�M����c�.]��)ϰe����QJ���e���ݻ%��K�Y�e���Q�zzC7gvp%)K��n���������ދҿb2<ؒþ�u<�d�Oڔm�O�{{ލ�>�^�����{��{Պ��\~t�>������A�M��^�T.q�y{�ny6�����1yZ�w��T��������׾�����!�ǰ�f�=�*Ǝ!=��̦�ﹾB4�� �������wD�{5�.��]��������&WO-��K{�yģ�I�!��ˎ��o����}.7���2?h��ʗ�����C�7�ڼ��3 +½�<���;l0������{�t�M/X�e�#'e�����Fz�ɋ�������Mܕ�
rVt��e�=��x�݌9�p>/z�K�2���Io�ꧯ���sO����A�ٍ�
������]&��g��,s��\Қ\�emsY��پ��+�o�I��|�4�MS�S��vj���h�>I�DKu⺥��y�;����h�p���ۣ��R�1o'��(!�i����#����[0NV�y����!�;��x��f������׃pD8l`�������n�{����W�_��8-ħ�0o!]�9n�Kx�b�0���_v�7{O"��a(����-U�{�޾6s�χ	���yHU?zT��qg_+��Cv{�=��roS ސ�<_m�o8�3ޞ#=�_u�zi}ݤ���`��$����!�K�<}�����ח�=̏�Z���veӈ̞\p�o�UE5ٺ'�_	��3E�e����g������C�t�[���=�O�xJ���j3�b��뛻��^�W;�c�;�F�����T7=78eQ�w@��^����ܬ�n�5:�_��xo7�g����bBp(N���ob������e�n�=Ȇ��0��x�����۾�!��g���W{�==��rz�^��o+��{�<��W�j姣缷�؆��j�zɓ{g^��+�'zv�\<E~ӑ��m;���o��÷��<�����'�o���V������9�������Wc�E{��Q�_93�� ��٫ͽ<��-Ml����6w9�称��ۅ�P��'o�rm�Rٻ���V{:$�qU���=��R<�zZ�p�No�ܾ+�5/<0s�u�`�ӽ�Қ��Ώ<{O���_(�=#X����.'�<��z|�p>~\~�K����x�<�k��}��c+W��[�LLb��+�j^ƚCxH��~�I��f{d��cc�x�ۗ�ޢ΅^+S��j�#;u��4q&�LԮ���5@f�5�������6	V��{��.�-��=2�����X��V�����gN�ۉ��>�7�u2�~���~Y��d�,x�$j�혷47��]�8��M՛	�/�}�OvG���s��{�H�=���y��f���0�k�6a�hΞ�b��;��=4N���eVK��r����m��r������-ż���qc�en��J���W�%���WZ>9%���do��B�w�)e�'�p�a�LĲ���ܠ��K�@��nVw'@��$�t�,��m�F׺>��w���ʳ�ڏ���&A�� �׹{ޏW<"2嫭��5R���,	[������4o�>���l^@w�ݗ7����=ܞ[�b���r��w��eз��wl{p�vu��u=�� ��Y��?��;������^��_m�7D}ڨ��p��.{3^zK}���7=��d�^�/��`�c��^'�`βJZ���T���$�7��G�������������ϸ}}����������.���
F_
�M��^�[����P�ܡ�B�kT�,P�<�X3A>����Ì=�� ����]�`l#[��􆶼W����� ����}U����0�s*�̠�Pm�d �'2�N7y~��,��wҧ�����_�4�;�q��b�͚��S<���{��aT�^���sp�h�h�_��و���p�V�_����܃��YW�Yؗq��]��x>�M�s�|�=/�k����胵�����I�ix����.JΕ�W+�p%��Q�7VJ�`  ���uU�81q͡�w9���:��s��q�ݬ*�?P��8��Q��br��8`]���)�ɷo�)��ԕy��R��{j�~Jm�E�����귯����3�X�h��}S�ջ��^]q��h�h�Onx�t�6gg�ByN*�k��X	8��k�y����n��6�]0̽��HP�|���x,��/U�����y��7���ח�����r��{r�H��f݅D7������䚎�NW�/�}�V�클�5���_JǄ��`_t0�ALǶ�U��܃�i��҃u7��i�t��
@]ǽ���oݛ}��/���=f�D%T ��Դ�ú�?i�=Op��q���0Fpq	rW���6D��λg���Wa�|<8�l�jE�B(ٳu{}�7�v��v�)�����)�پ=�1J�@<p:��J[ӷ������#�\�/E���bĩj.��K���}�<�cV<���U�/��H2����5��b��֮��4K���v���W�i��w��={�,ø�����0r������Q����]2{����F�e�=��� �5����ކ߲h�g�������E3��}i�MeU��}e�Y��X5{��U�;����p�-�#6������y#{�Wn�j�짝�M���<[Y:4���c-�9-L�	����Ǻ�=�R���xH����o���a�f��������̲X��"ZSʌ��m�|�rX{��~�=�sU=�=>?y��Bu@��/yF?<��8�I�����`�z�%�7�=T�s���c�w��h��݌Ľu"y�`k�1�Ҏ�ër�}/�E%_�}_���}L�U^[��S�O�?��g����P���876�ni��iwc�e�ȣup�������y�:�=nzf�%�9�؎�>c�����^��-ǵ�]�N�v��ܐ�-�:Y�F����F���n��V;j�I�;7R+��e�ݢ6Iۓ6.�h@�����u۠�b�M̋��;�.�շ#�;��k��5�Y�^�����s�^#u�Xn��R�R�;s�rN�\�y��2����ܼ����1�Ey2�wc���ێ6��8������7VcWM`z�g�'���b��m��:��n��W��q2V%���3k�Wu�:�klBv!��uO=�i�T�u����5��n9!�t������s����p�1��;q<�um��8��N8Ͷ�{i��\�uV�k�u��7[�Sldz:�sj�e�j�t5i���v�X�n�l��;sۆ��8��kCcۖlyz=��q��j��׸MX�z�]�;�2gZv���*M[�mv�u��U���,�<�n���x�� �=z{q/�N��y���㍏c�=P�/l���=��Gs��[�m��siu�m۬��G<񝹱 qͬl�^Nذڶ<�q�f�h�٭ڴ�%M�C�wK�z�n3k%�n�Ò�����9y��ݥ��Tq�Fފ��u�tá����y�A/&J�CE��D�s�����n|u�d��qG<��h��9۶�a�u������#[=���Z{cGMN���F6�ۏ&\�ӵ���a՗���j<�s��g@A�7u�p��mf8Asg{�3,�<U�k���dq��7V��9����w^g�;�<�m�A�׷s��n� 5����d�GF8�i����,`�9���x:���X�1��Y�v�<X��k�&*���x�7<�z��@����v���qֻvv�x-q�MդyV��Q�wOM�[&�^72یթ��]�;	�[c�
9y]瞼7�n�՜q�K���ڭ�l��r�U�\J��X���F6�h;��]������1U�Yz�G!�r������9��]��	D�ۧnl���XE���rc&Q���r���;1��ɬ�{��γػ[��d��<�cn'ϑî�q&^H{'d*x�����0/iz���>-��奸�8��`�G,�ms	�yϳ�s�y����v@��vn�׶xMa�؎��n�ֹ�B�Nݴv�W����m�v�����`�[ǃ�m`v{g0�����Y&8�ױ�3s�W�u�����8�U������d����۴�u�\��rC�=����^�\L훯mnS�t	ج&r��<��CtR.s�؀=��<�ۗ�ݑ6�)��p�7�;Gk�ɧYG�+�����.|=8�q��Y�٣�#\v]v=3��g؂�gZodJ�u�O��pd����'�\��ɺ��98x����u�g.��Ϯ5vyz����OBRg�u�4;��X�"t�myN���!oo����׎`�vCn\M��kWi�ٖ�A������\;6ݺ�{��պ9�l�2cW";��v��{f���m���\�Rr��8������vv��t&����6�I�I��y�����qN��\�G\=4��ƫ�WN��&�p[Z{��P�-{`ۍ��gqp��ٹ{C��y��r<��l<7G�Ìvt��I�{-��b{Aqg���p=iL���O8���;]v1tpp=����	mϐv��up���6P��!��Ti����ln<�����/���e�a[r{C�����s�r�ON۶�w<��d幻u�ϭ��7n���
T�pv�w^��:9�:��8�Cb�p�v�6vඵ�.q��܀J��Ę-$���{t�8�5ط'�)�j�av1�=���$X[÷�D�ۺ�	n�v��n%8.��4�]������z�-C�������N��>�N�3�m����)՝�;�j�s��Vœ����/
m�f�o6��g�v��y4<����F�뮳�O�ظ8z����v��=�c��۷-�oD����'vp�уڵu���,�b����[���9��D13�X�v�z��H��2��d;�ꓴ��G����v8lq���u�����ک���=u�m£�ng�a�<B�nӷ7cջN�0����^w �;z�۫�q���v]���b�x���N�v�ۆ�S���/n���������՛����1݌��ۍv��8ڎ^P;5����,��Gm<�N���C�ɞu�MA�;�31�u@���0Utqۮ�jݢ8�i�[�6{ulfy�`��T�F=:�8�˛�xr7�5����ܭ��z;y��X�>�&x���e�[��w
��[t��˕3�	���M	�coF	��q;9�\�ێѷ]n�Qې�g�Y8�K�y��k�WG8n���+�cP�yt�d� kvy��= ���N=[���x��/g�N{#rO�
�]]]���8u��;&tq���/;�.9�:7k�7�{�g�D�0\�u�Yl���s���V:z�Ʋk��n{�s��'m��vq[�sh�a��7;�Ż;x®���z�.�;���6�"�ۊ5�n:3�LN�n��狷��A��-��#����ml���;�8��Jx 솮սmm�6܃�اK���A3��v��ۚ�m��7<n���n�g����!�ӫ>���AʶV���n�ݷaLny�Pn�G���L��3�=խ�Y���ͱ��g�ӭ2��P��:�\���T7��v�!7`�����ۮՕ�kvݢ����f�q]�ɛ�:%�
�V�bqњi�{.1�e�T��O+�uCN��lt=nH�:pL^�mƭj�5[p��*�)Fb��n��!u��pq��рz^7g��뷵��=�g��w����s��=5���^3�sb뷻f}�{���v�;C��E�B����t�<�pNv�P�q�j\]�r�U����6�+y�m,]n�rp��]��z��vK5�΅�5=�(�����vN�����u<v݌g-�m��[A�7=���{s��^���p��O�6����:��N���kyƺᨺ��a�5��9Ab!n7[�g�/4v��j�5y�A�=���˸�k��:w��`s\UT���k6=E�P>���؝�#�s�v�䞲�y�=�I����Fv�E�qBP㭻r\�v�V�)�g���z��u�C��a�c����GH�q�p���)f�y�F�
p[�C���˙v��^m���{c�c���>L�k�`�wB�us̍�c��%L���j��z����6��wbŇ<4�V�9sk�W�'K�.����9�Zw;�kVۍ��G�����7�Ǉ�Q�p�6���r��2���뱞ծ�F;k#i"�{���w<n����sխ��
��`��O'dG�����r�٦��tc���G�G���ÌZ�����]��p;g�����M��ln����z��&�}��q�fv��ܸ|V�q�^��t��g��X��= &:��z�w'])����Fx:����x�vq]�p����v'���Ͷh�����wm��v��@yհmɸ�(Lс1���2��l��í�M�;9�ɞ��n4;w[�=k��̦�#��a�Y��^�y����ڛ�v���u�a8�K����η�t�F�i��s)������@L��^��&m��n�۸��պ-s:�X�=s;M����W�M�no=n6��n���om���I'sl��)���܌�
����U˂s]����.z泻<����rqrY��9v�8�۵�n}��	���ѝ�[�gq��%�)�i�m��ZxM��o\t�����F���1۱؞�;��۸�sq���I�Kh���h:��lq6�q	�V{�U���r�[uX�e��k�lկQ���:�%�6��K�rv�ME��k�A���K;����-b<gխӓ3�qƉ�iNM�4���Ju�˯;����$8����S���ɴ;�k�����<��{s���HXp�i��Y��n�r���,ףs6�un��ۢ��ۓ/�
��ك�����Z���n��;p`�	��[�������n�b���of1��l�����m�\���ثh�M�t�(�[ɣ�fw��j��E��H�{n1�]Pޤk���;t���X4���O�o�5�&#D+���3�n�qӸ2I\�[sی�+�V4�y��M�h��L�O+��ݽkl���fGc����v��u�ݞ��i�۬g������uJ����B��6�;.:�lW%<ܱἴ��l�ݮ�gEsm�x�GnX��ĕ��:ָC�ܑaֺ�O��=����Xn��J�ƱFOi胉6ۮ��F'��Kd�	�zv v� �8=��񸵭';,�y�ү] �����:�r���ns��e+�{uq����y�-m��p��ų������s���յ���^��ܜ�:{=���؂�RL`��6�ɲ�8�A�|���..���!�#˓m��H��p�@��"�\v����Ӗ�&����9�P����ꇋ&.$�abl��c7.p)͙�nG�V8�l���Jփ���y�U��M;�Ks�����l7n�2�q�0��!�v�n��:�]�k<s]�J9�[�7�@��6vu�N��l�<����8�@�;�\�a:ݺ�'���t+;:)4����m� GG<��c���2�����u��%m��j�v�:���G��ka� �d�c�x^��϶���wD�3x�Jִ�F���1�l���!ݎ���[�ƭ�Z�$y�{�n��V��5�����p��LoLg�E�u�]f�i)ӭss"�p��Pl��)9Ph��^8�d���k-$̂h��H��4��:e⭷r���l�v+���z������M�r����zʃl�UA��jh�Q��U%J°�`�ʹ_sS-�K*1Q���(�f#Z
����Yl,-mm,cZƕ��ٸT���Q�X�ڃ��X���"��-]w+�R�b*5��T��e��Qb1�e*UQv㈈�m�Tʵ˘YhTQ6�ZZ��:�UDq
�*ݳ1����[j�����Ķ�Ѣ-�JdU�ؗ��[Kv�1��q[Uk-imRҒ�f0ȋm۷0�ܸ,ZذU�8��F �Ub�ŔDb��aid�[n�u���J�cm� ����"N4�X�̘օ���yq�fR�iEDD[�r�)R�lZ��LbQR��eh�J�����X�%J�")5�1��[UDQEUFe)�B��*�m�����jZ�Z�����(�J��+iJ��W[E#X�J�0��AQ��-�u�L�UNYF"��FŪ��+U`�QA�Ҫ�UR��9�$UJ5i�Eb�QQ*յ��QU5�h)T�(�E��FjvI$�Ch���sne�ۺ��7#�]��um-Ʒ';%�jtp෷����<�e�P���Q��n����72.�eu�
v�Y�`�2s��=�r[U9ƃ�7g�э]�7L�s�Fk�&y�s���-�����wͣ�E��铭;�x{u�`9	���b�����v�i��=���ɷcn-����MgqSŸu�m�b;q�x4G>�/�IyT۱v������
y/\dNM��m�!�b�أa06T/n��Ȝ�>Gn�? �c��E�r�Ë��;k,�sV�4�\u>i�r(\sTqt6��aG���vx�C��.���stp�<S��.��I�ջa�q�v�1<�qm��*ɧv��,�D4Z{o1��}lϟ6�o��4ig�=I�m<y}DC�qpKȂ��\�^݊nwojm�a�]A�[�y��ums�.�{l�i���y�T�;���6���v���^	�m�n���/ o=�ks4�>{#�z����+�y�(6�uv��1��M�*-��:^�� �]�h�]�όT�v�h����o'[q�'�}��-��Ӷ(^������8���WJ�����g���Qg�����cH�מy�qS���c`�9��R�[;d����Ƿ����q�˶�P�jK��0���ܮ�0��2��j��̈F�8t5���3Ɏ�z�q�j���u�F��P���8�ݝ�v� ����h5�M���x-nݍ����筽�U�n����ƶ�s�s��.Ȯ�v��q�,��4S[��i�\	ź(�����֗/7c��� �稗�c�v9�|NU8�wcV[q�\+�^�������t���;M��^��������i��Ν����m�Ѯ���t<����^5�.�u�6�s�m��0Ʃ��tu���!�Y�-���m�����;'��0�{]��g�g��v��qɻ���4��v�ar5�y�ڵ�uLS�N=T��E�g�j�n��p��[�#�x��;���{��ニn6s��e�p[pQV��J��"q���|�s�W�� ym�L��V�s0�j��U���.sȀ�vM�le�1���\;��evǐy]��G0��̫lV�0Q��i�8��E�U7d���.�|n8v2�8v�ȇ�˅��p��<>8v6�/g�/n\�;/�/T�>|&��v�/g��L��������(����U
�U(_��w8�!ud<�$�~Wd�~ݻ,f���b����I&��|+><�0�&QS*�6ֺ��W��b�r.~�׵@�HW��7K�57kf*�ܺjע ��	)@�����B�$�=B$��ݯH�t��~;�_q���1�+�rHP�Q�b�v�Ϫ��˂A٭�D�׵Q$�������l���j�To��*A?���I�^�{��_�N�p����,&HٗU�$��|��;ohP.!�+U�TD/�v�&d��&Q�s���:�yάf:�۳��������'�O�����jf��b�s����o��|�
{�ۡF}:&7*��B9�)��Q1�ǔ[�8�������?upVK��&���.(���+��H���&�6�,�2���ɹ7A�h��y8_Xw�v�8�� �9��D��d�gl�hZN��T\|F͖s��`��y� {tJ~K=�f=u��F���D�
eV�m�t �N�\�?/lQ��9YQzv�	j�TF^܊2�eBDFIHBĊf�<��Fܲ��KշP��]
'�N��\������� �7�f0%�O��
%�ȿ��״�d\��]��X���G�}��#�~;�h�Kg����R j�b%��^;�3�v��4����pɷ*���SkW4p��������һ���6��z��y��9B�ݝ�>�Z�6}���Ջҳ�I�z�P&vYa���%������3�޵m}�V͈~�Я�����ڠA�R
��c��c�����宓
�b�
j���V{(Q �ǔ(�M�~�����Jس6���^��N�K"'y������.��
�]B^.�7X�4�������z�8+ly��r��+&�X	${Р	f����1�&�{�b"L2��׿MV�死D�}6�W��I"��4H*�u\�ػ�j=�װ��E|H����	HBĊ98�
?V/mE*��Fq�$���P$�q����n\�&%���\�<p���qƎE'�\F��v��L��ݢfR�"L#7�),d�
%��o��E�ɠA
�u}��G��/Ӳ0~#|��H>X$�̙�B%����_A۱�2郤4)^ק��O�o�_J��U�?݃�	��b�>���ba"g�flV��Q$�-��T��ܩջ�ު�X`PQ������Gݽ�M�f�w��[���~?���� ��?L�0KZ����	$��/1�)Hg��>��k���\=��ӵ��D-f�c��}�aա�lK#�?	d��^���VcY�]a����M�*^Q�e�{A ��У��8��
J
e6m�t �N��DJ&��xqDρ��4	���@�[��c4ś���nM����@0z㧸�7km�Pd�zS��`wKۭ���v��U����@���(F(PT� LHߏ�P%b�*�H�{_FNG�D� �;�*D��P�Ȓ& F�Dnk��G��z��=V�'��Փ�Q �̟#m������c״^�ml?f
 D��E�3(D�1ƚ$ߞȠH$/jB�V	�����|(��B�����(�;TȂbI&~&e��Z1�ks�D H/j�Q$�~�(��˩�U�i�3��y�
 ��Ɉ ���;�D��U��s6�� ���(�H�=�_F��
�8BB�D��H9�ʃ��?]3W��|�Y��R�-H���v�a"����n��(Kһ]{O�g�<�;��߄G�ۼ��˗sh�f����D��Qy�<���Ãa���8we��=�Ξ���ۜ#ړ�;���l�ݣ�[qg���7�w|��Vl3rtp�v��4���]j�x���n8�o]2��&�Uř⵬�n˝����127D3�a�M�!X6ɪ�9#&���ݙ{v���q�;��Od���Wj�U��\j�B�`����X�yp�;N��8z�5�X���6��Ɋ�&{]�.^E_F�c]p�w��~�ZP���U�r��|H$��~���١l���J�ݡ@�N��	�@[�G���@��F6�����M���P�5/�s � ����|=��y� �N׍����/st\��x=TR8	Qe(�ɛ�@�w�uD�����m����9(,��N[�}_wv�Q��h�(̙�B$�Efܚ{ �@1EX�_Ĝ��D��u@�O�{�1<�f��{�9n��;TH�fA&~&%�v��L{�,Bd��U��|��o� ;ޏ�͟��;�o��??��}󾫚��R��+��d��\n-/J���u�(y9�>찆�������Ә����>���ࢃߞ~�qQL����f�N-����w�;  Ic�`g��>��P���U�s����d���~ï�}Fh����3\�\Ν��y�=;���C�v[~P�3�M�5��_�%��ۮ�[i�㽀~��#��o�ត9�A$��?��	!z�*m�?��<���v�#V�Z����
�^�I�5����F���A�x ����<�$L�Aѯ��,WF�
�'p{n�[�I������hy�P�;���ĝ�:�Q������12�J�"�=�@�pˑ^�\�#`�������fN���[���;�4	w;��{WP�L��y��x9�&=����ݹ�8�w�7 UE!"(��h]"�$�����uH1�5�$��(�=���P �����c&��	��&�'�� �P\n����.�����(����A-bbF9�ww7UE��P|$��IAD�.���~;�$Q pD�D���no��Q{퐰�g�ہ=m��b�6o���;�s=c�� O'����̘�p��7��!�`%�T�Tb�7x�.񊝩z�=윪�"/gM|I�{"�� ����	�mf��ows$k��_g��Q ���
#"0z�ω��c�"���ti���G� ����dTG�ќ������|A~~�����W�3��:�"�H�T��%	��ⱬq����9׸ç�v랛��s��x	`s�����~�	�(D� �8�"H��EA$����g&bv����
�O�oh`"+i�B��P /��߅��+>y��x�6vX$�O�������t�3��4���1�J�)fA�����_!�ʪ �<n2��|���ѠM�m}@�sv�Ŋ��$(2PQ*��������I{�o
E��n@���5�?���߈�18��bK8�w�;nn{Wgz��mc�ʃx�Ab�v�?vr��������j�2.�^#����z��{bL�>��6���n{���a�I^0�3��L	��d��'�b�f��H9TҼ��Y<�cǃ���?��W>oϠ���_�����qn(�m�Ajv2�n���e�N��!�㶌���a�|����6��Y�DG�!��	 ���.�"7Ӧ�	��FVCw�ff9	�����_Q�>Zi}��(D�1YH�h�Q�=�dP �N��Q$�zt�&��ӋNʛ�T���Z0����"R�3�1,W����1�H�R�����a��c	]����i�gX���( �d�=�'��ޢ��6r�?G��ب����<�cs��ρ'gn����H�2PQ)�����Y??��,�	����	���{чĒ6�УrW�;@�C�!�F��]��;9)��C���V�!X�>��I�`O�#rsn��{'�x	���7o�����V:�<��7{�%�<���Ӧs��'s~3�9�Է@$�;� Ps��L���������+�����w2�cQS��Cr� ��5���`S�����rp��Wms��.�v���M�o\��9꧛\�ۏl�j/vc����N��=ۛ�ѣz��t�q{&<x�F��d�ī�)�=a��n{D�϶2�j��^{��w��z/V�]��n@��/aLP[�$�W�E�Vm��ΎwY��V�1�.9;��۪\M\�wې\z�")�I�k��پ���Q�@��#Aɬ���~�{B�����=�{r3i���xɿ�?4	b;�V�����x� 8н�f\)��&/Ӧ�m�
��8}���+��N|�j�Oۣ��E��o��	{�	$�ޯ]Pn��v��w6�$���(���;4n$@JB&B"%���y>ʽ�U
����t� �Р	#wn�z�F��"B��46 #�J10DL�_�m@̺���B�8j�p��H��f������t*U��S���1�~}g����ո�ɻ>.}��Y�έ;��K�|��\&� 
Y�wwT�?��Xw8u��@@���E� ������7��g���M���GB1����*G�٬�D�.~�|XZ�p�C?��9ӑq��}6 �V�a����:HZ�z��W�\���,ʭ�VRq3��6��r&��3�e���T�<WJ���dx�c�	�ݺ���j
���� �@?b;�-#w��JOė�u�H"�OrA�H�A����,Y������p�k��m�����"U ckZaR7u�Ӿ�Iu�"� �=��|�?/��㷺�����\�ְu�D����R�����b�k$���g��5�훁��c ��cx �g����{�G����A�ˇ�-),Y����<��j
�q�vv]�*�sgs�y Ӟ�9V�����F5 Ĉ12��e
�~9�r(��`Ĭ<��{0�< �t�g=`m�Xw$j�����K ����0�$ ^��H1���!J���ȓ�:ߘ`�i��D̠�J��7��Ts���N�������?�/��?��!��7ɳ���}��̆���ꮭ�#�wdhu�]ڰ^�Qdg�ĚSs�W�o������'>�h����t1���#�b�zg��u��/��{���]��ޙ;��!���a��{P]��Ns����(���bo�[�O���r���4�5�m�I��;�+�pל���r�v�������"gN��s�X=��>-Nrk�tg�b�;nzV��p"s_�Y���i�W���]#��'��n�HP<����J��;� �����,���;`~�w�H'��'t���9��vi�.i�ͺ�ډ�A��&x�3��&5��&[8�9���ј�y9��^�������7}r�}�q��oM�zh/[��}������wOx� On�����h_L8K��[1�V���Qc��#vt*Ɖ���v��d��"�Lx̰�r	Wci��YQd�H��.�!���w�s�~O��>���U�QN}��Yu�O��N"T�Ùw��V�x�����!�k��K�����Ś� {��l�{RY��a��u<�=j�/���
�ǫ����/����vw^�o_��.~E�r�a�?`GP.�����Fw&{}�]U�h�>�%���	�ˁ��Tvw�_w�\���a���r^�{��w���J����'X�=r���=��*���"��z��~�$����O�T�l:���;��{����J9u�����t�u���,���s���w�ރ���y���[aķ�I��� �w{�lɈX�����8"{�pL$�bL��#"��R����j�Q[jX8��Ur��Т֨uh�7
��EĪ���&�w0w)�*�UYT�61r��X��yy5���ġ*pn7c+���۷�7�^dv8��M��@��z�{˄�k������.9J��b.R�r��������"��KҌr�3
Զ�QKs4tV�C��Uj˖P��N^9�PE�Q]�q�my�)�mF�mm�8"�u�U�nJ�-^[QЮ�����DGl�Z)���e��j�,���P*��+DL����X���T���n"(��0k2�#13��DU�1Fڊ��k�C-kq�1G)YXQb��b�D+Q��YhS,�e�̪[EA5(�2� �����eAUQ����mDTU��fR�+A�
5���m˘M�Z�Thԥ�TJ��ET�h���
�X���̱���Mn���eDI�D(�mV�R�na�Lrֵ\�E5��XX��
"�֋�c��T�F#Z"�Dj��"�*���Whjǜ�Tc�ѕ��AR�F�Y�)��9�vp��R����w�zC����o�y�	S��R�u�U���lB��b,|<G� uy�'�kc�{��j��| T,d��}�g@��d�*J�g�o�%dAd��w�M��Tgl�Ps � Y��D"u���7������3z�'Q�7���!��!m����ϻ�At���_�o7���
�s����D
�}�|�*FJ�*'���\Xt�����gE^��=`����aLĠ`/�D�Q	 \+eF�O�N	�^�v���4;�;��b\A�����主)�L߉�O�;�����*��+�������,
%HY�w�K������j#��f50� ��a!>��2 �!�{�8J�A�S~�i\���t���N���qgBe*_>�/��O��y߻;d�
2V$�.��>�'L*KVJ~,���'� " @���eufg@�����G��Ӥ���K��m˹��Aa�>��C����[H}���HV�+��~����}�o��}�����YA�����p� ��d�~�qaВ���/�i��u��z"�)�s͆v�����:d�!Y)�;��s����J��R�ﮔ�CR5��h����z7���ZT1�NizǑ�N��������aļ����:H7�x�^����Z�i�h�_e�y�ן��{7�	��O�x�߭Ћ �\�m���nf��9����{���P�%O���Ι:A�����i�O�!�7�	��D"Ͽ}�@����z�8������=E6�5�X�r@8�`v���U�6:�W�0n��v냊セ�����Ɏc��ݹ�c ���y�C��B�!e�;����BB�HT��{�G`�?hYq����~�%���
2T(���za�IXo�t�{�n�a�L����
�w��L:dL��gy�3���:��s����A+!bT���t��
�B�}�ߴ�GV|	@��7}/����S�'k�C�C? �fw��\{13q���'�����YH�Y<���::B���IX>v����o�ϳ�_��N�%aY+=����AN�,���}����!�o?�	J�R���������ώ�G������d-��������HV�*VJ~�����:� VT�������s��}����$�>*']{��ä���{{�q<+�����*o�g�2t�d�������e`[��<}r���ö�T�_y��!��Ad-�����ud�
�}�8E: ��R����5�+�݊ٵsO���Ruj�q�^1��n�B����ɝ��s]��u�����`{S�,�?nh��{�ʿk�L��@�F���?�"�
 8D��2��umun��b�\DDѣn�-��[��0p�`7L����i��Ӏ�3�mc�06�ݻd�p��z�<ݙ��g�V��[\�O������B;>;���iw�7 z&��X;u��[ �ԝa�Σ��+uӷ���d����n��N����ݠ�W������2nՄ��J�W�R�hm�{���]���^�/<v�x�ヴ
h�%��؝��k���č������]��-���nf��9�����9�,���Y*{߹�:d�
�Y��oy��#�~�����U�~�'��e`T����'Q:BSN�9��1�nk�oX��7ϻ�!�Y-��N��u�����;���/�!Z����}�~`q�Y�D�����׶LC*�{�Ӭ�|'�:��XuVߺ�Ϸ2���J���O�
���~�����������e`PJ��*C��y\�׼\������ąk!m>��Ձ�VAlHV�7��u�)�)�~��Mܸ�:���~�޸���褴�����?2 D~��{��d�(�����κ"��%aY,g�y�\Y7�����zn�u��(���{|���C��yٗ�Q�5��o_��Xw���,�V�)���8�$+�}x�߻���g<!SсS����'C�*o�����*$��|G�׎��2>G�뎟{���	�)ދQ\�Qv�u�v�J*��5�,\E�_Ǭ����\�_��g�/�<GK��۽���1�/^�d�!Y����A`t"#��yTH�?�#�ڼ�f�k�~�jB��}`q�^��o����C�W���
%L�1|,�}M�??����{ssZ��6�*��s�:�s�Ղ(�����=颌��=��_����\�sk;ʯ'�Q�:+|7 �Z�7?F"ELQ�sd̥���#uV���>���IXS|�޺"���Y(��x蟾`  ~G�#�{;Ì����M�ߖO�!t��;��:��v�����߽Md-��y��qzHV�
�`T����<��ﾰ=dAgɽ��\"�Q��Y*޾�Xt$�,Ͽ~s͹]��m��� �__��߽��|����y�<dN!X}�s��V�*T�;�ߺ�Ht5!Z�Yi�����9�,�_��g�|G�����`T�����q��e�u�|����+,@�X�S�o�S���.�}�½���~����P���?%aY,g�}�\Y:B�Q��bR7�5�̆Gð��x�GtQ;ƍ��/���E�<�'=l�s;u��[���<Ce���7ww4��f���_W0�n~����9��y�u�[d)i�{�8�$+ �
{��������|�/�`Vt�wκ�:d�(m�~��qa�$�.f�~�̞��[�s?d�o?P��3�Ȁ��tk̳S�ԽT|��˗_xc�XJ����{�JC��+Y�>�5�$����*ȍ�w �i�K~���&'c�޾��Ksn�gD?'��}�,�@���P�%O�_��?|��~�?}��ܟ�^:�����;�nh˜���Þբ��N/{��aa���'�;^������0�}ɉ��x��E5�/��m��<��g�3��
��+%g_{�\Y:����S���ud�:HSN�ٍ��pݹ�c ���u�¬bޛ���~�pK�#���z�lHT��>�>���:`VX�Ygt�{�	�oO//U������5FJ��z�XuV��tg�r���[3z'䟆>����C�(�d��a�3Ϲ�t2��9��������*����JC�� ��_z�8���I
�7}����S/������u��o���������`kN��ӈ^�"����fmӞ�g;��=��(W�����g;��h[p�'������
�S�o�S�N��IXXy��:aH����j�6��|,����7�����++ ���:�t�$)��?|5\�]�m�� �w��rL���u�o�����畭��w��qz�
��R�{�u`t�,�����~߸N!�2T+%Cλ���Ǿ�'�}�8��$�,�{_s,�n�ۺ�D�:T�o]��L�
�D+�y�	�IXJ���m��gw=ϳ}Y!�Yi��3��^�/|���"�L�ڝ�x76��1�,�:|����O�g�v[: ���
�*{���:d�
2Vahz�4�Im�1C��\'7YTwG�s�����z?/{Pg|�6�o
׶�76��o��n]��{I�v/�[Z�U���D�Zc�J@����Y���e�
MV������UD��_<��>��7֮/��ʙZ���?�K��p� Yy�l ��i�-�y{�{��;G�4���7q.+���pS�^�6�i'U�nu��<�p#=������Ӻx>����7��?�$/޶�����/�/���Ӟ�[D���w:a%���~�*!(�`ϻXm ����zV��s윪� v��l��n4���p4w;B���o�MX��I1UI7�_w����Zl��_Z���,��G+�薒����J�x���>�*9<A[�ñ�N������b��Ղ s|�` >G�m�ܱ�y�Gh�^$����-$%��萢TɃ`]������PK���pj�-�ٵL{�@�����0a]�0�E �{��_{�q+f矎#5F=���)F˺;Kv�ǧL�L��d��j���UL}'��#��8����i%Yc`�B�%+0���eL((Lv���h�z��x�V��[��y=j���k����t�������c[u�٫�tn'���n��*��g�q�f��ml&G8�A��s:�ʍ0���ݮ���r�A"{$O7Q��\�`��F-��X^��'��k��us�D��枮whݜ 8��vS`ҫ�sr�᣶T�\2m��kUs�U�;!]�ގ1[��K�����gu���ۮ�{q�]��$m�z��6K�د-��yw�����"��?~H����  ��v�h�w�Y�G��#���z��	%ל���#[�`�&_D��[ݮ	ˈ��ei�R��9���P  e��a#����M����ǧb/˕��=j\ḌB�d%;ewu�� f��[@|Ŏ�KV�;��� �;�����wo�q�Ԙ�"&~��(o}9�� ��̉説+������7j�$��To8����ͷ�lT�u��M�Xr=�ߦRH�sς��ֆ �}n��@r_}�'݂�߃+�j� �o��q��rAy�뗳�o�
�Xtf�>D�Ć1$nQ�I��Qݗ��*y�1�L��		/0�����o޸�UDά߉��M0@w��3�,��0��(;��ٸr�hQ6�[�L��CU�����*����Y�n����L_��٠�������b�?vT��y�Ev2���2,�����p��{��ϥ,���V�����:��JU-�uFjBG�f�ED@PϬ���읺�	 3޷��e�k���x����5lG�f%}ݥ{�o���^N�R�R�=��U۬�䵑�nz�\R�?V��6�ē*z����?����c
������I]s\3�>�י��Z����E;��RI=�e��x��\$�1��#*��z�-$���5u�znqg,��]D�L�ג_$��d�M"N�e��b�p|�;�ӿ1�:���9{� ���k�-�N;r#�S`L�c\%h/�������G����������O��|���ƛG�����]�r��������A$קZa)z��:$LI�2�w�A�6H��g3�*��}����\_� ��k�?I��a�MF=ɺ�|��1�|���V� �������N����s�A���$�y�.
��.�}k�-Өq4������I3����j�4e`~�o:f{�o���r��a���ݻe2v�5��baSu�!��������j�9~����nZl'[S�TEM
TD���_t߽�/��_G�u^�˞p�K�F��($��m"W˻��Q��wk\���3kX�]�q32�&>��	N�~�a�I=�-��~���4�G���r�ƀ��M&@����p���]�;{�ӝ���n�M�7���b�>��D/F�qں�ɗu��x�m7*������߮��H���V9푨���Zi0��p��{�a緥�^A�>~��9��K䏹ݴ�`śL,J�EL�9a��ۆ|~Օ���Fc��dx y��i �Lw]�Cy~���W]�ȥ9:�%����:$LI�2�,]��|�a�RW��J	s���[��UQ<K/1�1���L'Q�� IU%T���׳ױ�|�τ;�䉞��m$�J�΅�HO����BM�m�9���H�U��7��^��nRbb^}��|tTL[���u)h���HG����v��+Z6���n�9w�~���
����:W�vX���N����0�[9v#J�fe&>���]y6�d�9�4N�<�ޥG��:���K�!��6�@̷���ۆ���DEg��ب$L��*AS*LDk�m:������t��w[�n��s!�^U��߾�QS�a3$�^�^{�?� g�M�0ʻ�n���]ͬ�mr�����l6�(+ަ[K6ˈY�1��L#wgo�M�?oc��gܭ�|�kX$;v�m"T�u2�I����j��/�w��]���rBay����{��1 ��� p�x�u�s��F�_!�� ����\yvb�R��QQb��{�t�vM�&h]��I%N����U�e�i@_��e�=s��]��`�k�
MW��$���T���f��@$�}͵p��T�`��U�>l"[�[�� ��u��_||F40ש)��9)��&�D����S#_'�T�=�O4��G���||�yǬ��y�%٫�ym��T~V����j$5Q���"9�O����B�#����������
:C�*s�c������N���v�����X��ړ��&�ĳ��dg��GF�݌KJ����7��k��A�?@�0�����|=�|����z�;����%3��^<%)���,���a�7_h�tf�4Pkb��Y9yL�N�{�_d��i��z��pvs��dzG��ـ?x����i
��۫+S �L�8tǵOS�7"=��7�[^��v�ޚ��qΐT�����ߴ������x�>�9�����7W���L��ݎ��D���29x�1�|���{k���;�N 8ˌYS�tȺt��0.�7�q��'D�v�N�/XOd��K�x�`YV2ٱ�/����Zw��7�I����e!��y�n����O������U>C�#�b\�Z��p��7��s��۷G�î���|^��X���ͷ-���3�M��&X^���+������᳁e*G1�M,4� �Pa[�j�'��^'�<T���x�]�۞�@{�\>X�wd���m��9O_a�>�Hh>��
{�N}�w�ꋱq�e]n�ߞ���b�q�V�z�O�M�e�{����G�j����QS�К������NQ�8����'�=����*��7�����E��S���p*01�*��uHy���jD�͙?E뫞Zc`*��""�l�Srɀ�+-EK��5��.Һԋ-�E�®Z��` ��i�[\��L�R�q
c��u.YYS9K���Sr�su��Umݠ��[���R.R6EQ����v�uܑQ[��f�2`�Tm��MK��[j���kW]¥R�֬b[*��V(ңU��rűT��U�f6Qb[b�]���p�,�T6ՎV�f����-�
��-�[L���V�-����(�+m
�
���AԻ�#9e1��e��E���X���5F�ֱpf��ԼLq�����hT�-�R2+�.R�tl���h��q2EYS�Z�mP�X�ˊ�j6��2���PF-�F��D}h�2�^2�vؗ1��C+m�n&�<h��V�w���2�ED\�x�p-�)VR���QMJ%B�D5�Tb��[E�̺��b�
�TPkVj��*J*��,L����TEQ�[mc�V"������lĬ5�Eօ��+hZY����/Ί��:-��V�n�b[[Ks��"y�N@�)�u�8���'[LD�&p���ݷn==�F���1w�^}Y��Η;/�W//cY���#�;&���r����y�X0/nd(%��<��:Ō\]��Aa��,v��p���v6wS9�Һ:�7b�����r������̛=
.�:�7m.�H�S����7Id���%Q�u�G��8i�2[;�(�g���湪��v�bY^�_2�wg��ׂY�؎��vC����k;]=&�g�3p> Ş�Y<�OQ�T���C'�X��km�����O9�:�z�^��v�`��SjI3ϸrƫ� ���ݮَ�"���ɇq��e����am��}��6�lM�kkt�n/&���9�8�N��\q�`܏5��N�v�Wz�`<0{[�)t�=�܇n�чI�t�{K���\��N�m:��s�iCgo�箓�r-�r%��ͼ��WN���ۍ��=��m`Xk��5^�(:h��e�q��Z9�m/P��q���`��;M���k��+�G�m�Xwl����m�t�{v��⴦���=�7n�;pHg�o;X7mU��B�\�r�ݸ��2ݞ�۷Y�q\�Y�bwH0������ujNu�;`糮K��	j�2g��I�I�^mOc�ZL�ٌ0���n�z&-�cU���!��m�Z��魻W]P��h��_c��H�39w�%DI㛎ۘ�s��`_Y��br��7."׫��C�ܯ5���7h�O�[]��˭��@[]�;��-tݷv:��R�j�d����S��8��G"��F�jnug�=�l�F�:�N	���2'U�8�v���λ۫�=�4lt�������v���6���;�'U��8���g��qݽ����z��筹����Ʒ��@���4'dv˛N�Υa��5Pku΢�w7���W��&��Lh���fg�[���Q�v]q�l��*�[v�ݞ;��7,Y��<by���p�Nv���ݷF�u�d���\\en��k��ԅ�<�\�.��(��#l�;����L�S�\t�)�8 ����ě.z�u�r��8��m�wmm���{K��]��'��4�v�sٱ��+��=��g�MţL/���q��y�q���q�Yn��밻�=Q7w��t��|�rO�n"�)��m�ݵ�s3f��,��<�F��v:������rn��l;J�s�g������vژ���S�ֿ��O���Y�� @}{�i������/��;�F�oK���+wi�HF��4AFb!D��"�/9��	{���vG��w�CA"gwf�$����6�'T5j]�=A��GF喣 � I��&��ю�[I��ݠ�I>�f`�}��_�" 
�e2�H�^��i�NVl����&�O�y���
��o%�Fcum �@+�y�I/�=j����"+��!��L�����Q��J�UEKO�����|���Nt�y,��f�ݠyy4ZD�^�l�����mS�~J���:����� �J\/"��v���d*m�n�olϵ�0� �|��~���Zfx�������	 �	W�h6�%oOZd�P�s�L���o�� H��l+x��eLT���&��K�:؆�Ds���rBKƮ�:�/	�v�yz	Ąѽ�\����ը��i�ni�{��5����F�^R�	v�.]��['�+uｋ��Q*V��W�|����֜D4B7kxQ-)�����F�E��z��,F�7�a�1D�5gy�i�"3g�iK �[�o���J�.���|q%��l?�Ȥ�zz���h�*I�"ff	���}-��]o\�%�~w�'s}B�-���p�Y�x�voYsʾ� 	׍6	X��
7�MZ
��5,@ �o��
�U��e{��<��l9��� Vn��AU�^�'>������|�9�-��sF�j���u�v.��wnq�2�[���zœ__[���N�]�5sQ>�Z0��5��qL�~{nZ�uv����3/��5��y���	310�cz�<">�1V��+�y\�����|�"�#;��I$��� u�懃S�f	�ģ��%�	u��%%�4�A"o��K��ۜM�^M�UX��xPo��%�xm�Ɵ ��of�o|��4K�d y
��Q��a�Rl]�m�;�/���a�y��}��������L��?~� �؎L�+�LQ33C;�֟r)ז���w6|�'����ͷ �/{�}51�}�w9��v����GT�L��C5����H �$P��Z�n��S�\J݄���a��S��r��wm4�R��Wrf6�\��n��۵�X&��㠽5�ӭet��#c��A��f�����g�U:�r���	�\S2 �{j�nE>x��������%
��eń�Ό:���eUW`��Y���~���Ȉ$��{[|PπA1����"��i�Ȉ����>WUׇ�P(G$DDL���R�����m$��gP4�G�=Vz�q�޵<����b������� ~��a�m� �&
�B}wa'Ϫ�W�4J�[d.���>@���� 
�u��=�XN��jfw*�]G�����2���}G{�p����p��F"��JK�7:�=�oj��m��{B��^S5�7Ӣaa7e/�|�|_��ΉlTq7��	�1�+���h�s��(�}~�g����$�s4I_#����6�]��Uzj	�
�)
���+m�B�̳��l�n��Dmu<�a;]-M�U�}��h��b���_pNm�I$���i� �����׻�l���b�^��� �G�7l�=0J���
�r��忔1N���V�D�/� @'��M�7^�� 
�g� �gzvo.!�.8�T�5AT\���:�`�A�{j����&��h���~��@��6A�F��M��j�dD��UU5(���=��{y���y` ��֛T�P�����Hd�U-��0N˦}��֘H�vP4���0J٘Q0 G�7d��V% V�U�v�1�>矼~�0�i ���I,��D�K^Ŷ�".���D�\w��}&�0��z��Y�A��dy���e�38�䆙��R��}#j��O�䗐+�'��ï��$�;�{v�f�fenk���F��̜{<��Üg{&��vġ̚7V��gs��6���yw0Q>םn}Y;EKn����OFzv:��V���lm��@�����$)�r������y۝�r�=�Ѳ��W��(���q=q�.��[Z d��K����q���G��,�e�t�ۥ�z�ظ[r��k��ʴӳ���j��]�ۋY��g�]4h���\�b�;#�ǎE���)z�'�`ȕ�~~���^�7�r����.��(�'u�?�I��;�XIb��[1f��h��WϘm-��1�3(�ړ��$���b
�#ͳ���m���� �֛ �n� �y^�=�i���t(ؤ3 �g�e$�e΅N;�0"=�m+ _���m�\1�I ����E���I.��rL��TA��"w�j�fV�8��ɔ[�j*R�.s\� C絡���z�a�:.���/�	V��!A���Hɻ]K|���Os�Q�&�H�}���Dz��W��;�_�>n�lU����񏧯�����s�x�m�^c�ȼ������C�6s�kno�C�|��p#~����@����?��K��
%���j	$��P�	;[������JEU�� eN��T9�J�)*X���� ��K3�*zd]x�7��z�����tӽ�HY>�ڂl�}(:P�����q.s
�@�4�5V���񥗖�k��ک�����/�_k]��|Q��,I;���$�[�\�vty��|xL�1���7f<��	9�OݴH A�y�K��ۓ<�����r�D|�i��B͙$}1AU.b'q�v�<G=h7�v� @'������|�]�ޚ�˓��I�;\4��pz!eD�UA4G8K�Zi�	7�n��;���� sι�`��6D@��kM�<���}S+�Z�I3_T�Ċxإz��A۵����)x�î�ݫ�s�+�K���ﯯyL�SS������<�Zl ����ﯼC~�v���1�{��[VL#�2�d@_D���u���k�w�K��\��ס/�D����7�Ou�
&�Rw�z��pw�W�\V�IH��\@�>D"�%1wz�Xm�Ig=�Z�%�DG2�o5S�垞��տ�u�.�i�f寲3�����,Ã�	��{�ǡ��UwOe�=����2����<�X����d��&<~����}���~�sO�����dDG��m1�]�<#�f(���j|��O�d\8�_� {�i��� [׭6�A���U^��F,�Փ\ַ����ab�I&E�LEMK"'q�T0�ճ�rw��d�z��sް+�Zm > �=i�@C'��%�F0o]չ��1hDD���mS�	i"'�=ۗ��V �<�zۤ�8�0�j���"<�b��&�՚��u�� ��{B�I�N�4�TA��1=����n�z����JY�Xm@c~�0���0e�z��o�n_s������>`�!��6A,��K	I���M����i���;2ffD��O�N����H%���i@��-x�ȩoEP��|����?��/�n�S�Lǀ����L/^s��Ai,{�D�>�K? �̷��u�[~�;]�ٵ�]���I� ���tȑ[��)��Ǜ������U�ww۲��|}u�]y؎s�yyB��
���.^I����tT��������| ��$P[O��k=��UL��Q5$w�Ec�M� ��5��ꍋ[7��_{:�d��@]fS-%�D"���i��N�Y<�+||�~�?�mՔ1��9{nl:8�H�����p���k��u�1�����)ߝ�F�6~���_NV��	 �(��	-#o<&f�Q1g��	@��L�B_�'D�32�$�j6���rql�w4�+2�:ږ ��\0�m4�A(�NE�#�[8��2lx�	�SR��]]�l$I/��_K�;#+�6v�!�޵�'g�h���$�s53��"fdH_D�O8����F��p�چg}^�򭀑� ����OO��aU}�8��X��ᯀ�)NE3�}����3Z0�·���y)LL�����L��%�v���#�U�L���L�f�'��"����i��۝�f��T�����g��y���Հې���X�U{`������0�$�=#K��h�{Z��o�n�#�;U�X�> >�&��B�3���e�����u������N�a���t��:ͮ����פ��:]Z�l���Y�*&���	����� ���n96�X���ϕ�_����\v��Nu�g�N�l�W\7`K2��t����ø�K����;Zz���٤�[�Q�wj��:������֝����a�N.�����^�t���V���7��	8��1ӞX7[�z]q��l��˳���&���v2�DDAQ?<ѡh��Q
$��>��N��������$wo�s�˅��G���pn��4y�i�T�Vx�bQQ1j�S��p�V�[\
��̙���� y�ӈh�OF�}��M����B]�'D�33M��:��L�se�R��9ViɎ�߷+=�	� ���� G���0����\"L���[]�z��������HA9�i�	 6��!�����Dd�$���jf�('bD�̒��l�Ȯ�����l�Kb���}M|Mg�2���"3i�� �ڸh.������ՙ늅`�Y�m��/8�9�q1q��(���sd	^U�����H�����'��_ϯ�_$N�=b#D�S-+,=fU�`��{f��B��W�\�����B�Q&f�1�sXE/������x��A;�H��7��Z3�i�(.�����g!�xu*�<R�[�F��홯&��B�xOb�OO7p9�Ɉt��-T�>�����}��4�%n�~M�����E��5o��I�z<h��cZT��B�@�DR��m�x[@ �fմ D:�\��z>�� �7�z\C�ڸi ��i���FfT�I6.�u�6�+WVr��A�{��F@��.{�b���m�����I��>i���D��SD��&=g5��!�}i���s�]}�����X��[���eN��� v0�kl�����p��B�����&{[	�s�=�sM���+^6:1l�ˌ;����k��zx���LG��UUDMk�}��� 2�z���ƛ@�yT�I�~�����{[�@�(ܹ�za2aL�"�J*a��}�?�I/���-�&"��&��, >��h ���#3����N��5E�`^1bL�#waOM�j� ��i�@|��
W�X��߆����b�^v�]��s�]�=�����g vT�v]����g��g?����ve�iM�Y�팜��	MU�@�;|�K�ty�C�-�?t=_�d�w�Ư�DA��~�zv��.���Z�i۹�݌��>>��j� ��������{��E���v���o����T��}�}�~Y0x�9��t�N�Ɠ�vt�%G����^Z��ȣ�9Ly��i����F��|�͏=�f���Lu��<=��z��� �4�4h��0zwG��h�F{�޳ǭz��\�}�g��tB$�@�"1#��e��A%b��Ze�H�6�Y���}��!���1���Lu���Wؔ� ;� �{���C�|�ѣrn�>���u����Ö���r���A�ٴoc���ƕ-�I�{�rh��kua���H��Oqw<ݨc����w�� {y���1w����9l�[XŌm�=���jL̡`���j���w=�x`+��ٳt�����L�ɹq��r$�z��w�w�9�2�߼`�1r�@�^9�����	}w��ˬh�;^�� �x�b��8�u\�˥��ta�5f�L;�00�n����^#�8�-�	� ���o�ۇ�b�&���*����5m�v���||�%�\{��O�q��i;�NR�S=[�/m�-�f�o7�훅���NK����gr��I7'�{6��ּ�&ܺ�R�{���E?nk��c���1��;��ЃշQ~��qd}���o�s:���s���I��J=!U��"�R��B�Y^��D��11u�)U��F�k[e-�T��U��F
�`�"��EDQ5�m���ER��X�X*��*��eEQ[S�(�"�K��Lcj*���b"��i[�0�������31R(�EaPF1�U-*\�"W�kXc*���PQ��v�X�E!Ī�0ܳ�����c�EV��MA��Sia�^Z��DT(m��x�k��`�TZņ�Z��X��cj*9J�q0C[iD��l�(T�X"���)N4�T�+��h���jEf��*�u*[QL�\�֣�0�Wl��n*V�[IU�����bbb3n�1�e��*��R�m̅5)��N[l/�E��+Ə�R��D����LH�a�A2�f*":;��1QL�)YL�J���̋S���H��D�����N��Hﯳl���ϵ�� ��4�.j��Q����\��.����t6�ի�� �'���� �/��\ �7k;�G[�r� ��m���0�(�ʘ�&�ڎ�bŁp�D@	u��z�f3Տ�٘ >�O1� ��֛ ��6S�r��W{U���$�=;��٘Ir��<Oc�w1���qF덼��n½ ���{}w����.�߻���A� }�ݨ�h�ֱ��T��%x[B�GS��9h���W'�('�"ffI_D��]q��4�٬�^��N�	$�w��-�[��6�HH�]7��4����O���s?"�D6?��5��Fo���`�p�f}D�ԓ1wO�����W� ���a�{Q�
:tj	iL*����y�"�_�=	ۼ�� ��4�eO��*���>�B��Wt-�()�@4**L7^$w��	���&BܼJ���G4�T*ϼ9�59<���<;Y����y��_��| ��G�A��P��i��Q5,��-�@|��g�����W5�ׯ�G�1s�Zm �7��4�d���^]�Ѧy�L���|L	���&�`�nM��ֲ��\j���˙zup��ïY�j��CA�fJ�xYX�i��V� �A%��	{;#�oS����b�%��z�`���Y �)����g���M�������O{��Q`$�����a"V�v8a$Kw����k9�s�+]ࠜ�32J�'�'�uh-$NJݧ�_%�y.��7޶0��з������r�ur~�E*��M��7�l��*�>�eg�� �9;�X^�5��TS��"ʛT�ߐG[a��7Ĩ�R�A�30���z�uؐH ���6V���}��u٥�g�:�l '������q��^w�������a!�,�4z2}4���m���_d�r�M�d�����ݻs؞Z���"�R���JO	�Fʨ���f3:���'��O�����n˅�r�\�Ǘ��ϑ;|3v,��9֊^{3����M�u[�Z��C����O'��㶬�޷k7����4Rm��V!��n;��7>W
n7k��۹�^�k��^��[8ܛ�i��p<X���9�1�L[Wz�7f�sѺ�m��j|�J�<T�Ń`.B:g�3��	���v�Thی��DAX훜C	�nCU��n`'Hj͢�Mwf!X۷m�M�m�Ru[�n��5ʅ����!{�`�����Jx����~�w?��DT��Es�C 	��V� H�{m-��ٔA֡��j��0�h��}�E����D	�*B�w�a��Kk�^�w���]�-|�	Fv���'Ռ?�)'��z͐�u\��[PΣ�*D�2&aNw���H��m
���I-�fҍ���es����İ���ZD�[��!��8�B��%}3wiu����q{*C3�6�0 �{*� /wXl$�AoW1�|2���$�D�����(��N�BJb�z�K	{�i�^AN+�Ñ�~D���S/�J������z�L�]���s�j�\-h�'�l^;<.	��m��kl�q�����Lk���Cp�R
����7�'D�QU$=�-춒I%[�B�$����l%^֠�g��϶�$�gc�8t# �(��T���������^��{w�v��������i ���"�z����*L{�|�O�/���Ѳ8��U�����%��7�*]K�w��g��;�k�ݧ�D��'���{��l�� $�����G���6@�/j�^m똚��iВ���8�fd�
Ř��{� �vմ�Y2ע��o*���D���� �֟�>^U��#�p����0�ݩ���<����ʱN�b}�"7;�M?��k)U� ���SN~~A\���m��vq�����HI ���'e�ih$��͚ig����lD��
��i�?����4�d9����o�_w}����X.+]4X�/iTno&�`ݎ-�7��6m��E�5���;����}�~�nFJ�#�ݵ�0� ����8�9�n!2�j��cٴ����u��U�I �^0�,��z�&eU*�#���{M����On습��o���|���թ��%���2K	{�]�+p�w���N�m5�,Y���EC��崡�������[H }7܉���wg5v��#��_�2v���.ԟ�͖�j7O㞒[�A}�^e��(��A�Ü�j��>[%���d��[�y�����}��2� >��>q�����	�����J3��e����d��f��U��<�3n�*8k�K��[���j�*~>ݦZK�o��I���M
Q�G�$���?��(�	�J�fD��L;���@$�U��F�o����VY��f]Тo�ӛ����wZi��z�v69Ǫ�o��߾p�a�bŞۍ��vxo^|�J��nk]�k���`	UP���D�n���Q3 ��{	�������z�!� 
���aۥ��-�o�mW�;v�a%�a+�p��"�c;�֚dGT���w��n���"��e��&�:�����s��.o��DD	�3ݟMt� �  ��Zi���ї�m��S|gy O���!�E�5��2=,���URUXnv�nq��}}��<�2��>�����{{w2�s������{����n�|䟽X��xn�<y;��᝞.�Yu�u��tW��}�Vd�Ga��.)�4�����U	�n�Te�B� ��g��/��4ZK῭Y�5AQU$�9�Z���@ ���hs=����(���N]�h��_$�wkK	%��ņ��;�����W��Q��#)L�C��:"ۗ���`���ה��4V������6��t���&ao)����H$���4��okb�^z{�4=�,���2�H�]�B��e�ȒdJ��>�����-��6���5sˬͫ� >��a���#��ŴPJ�3�>d>F�I���H}�L+@ᘑ$#0��z�Xi���W�� {���5O݌���#�|^�4�d ��������qL��	�*R���O���fo�f!���H�����$ m��.!���O�~�ǻ5w���j�Ēʿ1FN�j��fH�aTb[��4K	F��0������[GZK�[�H��˫+K��_FoS,$D�=�%a�j&6�
i��ҟ���ALy��`'���HQ؄�>�(.��M�(��X��9���C��={���ݣͰ[�f�~���ns3����~�������|�T�G��\�IE�6fx�ͱzە��џlV�!�WU��m۪Y;V�q�\��e�9h�\<k��(j�\�2Z����@땱Yݳ�]��{g�7�۬y+wl8���9�s�$㞌v��K��v��p�ȩ���3����N��.\�2��*N鷭�dnC��=/����� �uVݫy�tTn��mΌ]!�4�g����s�|zg*�حY�=m�a���4��m� �JO�&	��|dIPTEQD��g��ƚ`�^W�Ā�	�m�`dd����u�d���E$n�x���:qD�$̉1
���K`$�K��iòw�{˫�� z����S���""����?�ײ�)w�`XKpo�I0�y�j�DNfհ �-���e�C���y ��u���ݷ�$r:	�2B3<�nq������vIK�ۆ|�;�W<�~f�H~]����F��i���'��ʩTPs�H��)��@ ��Zi��^z{i������E��i��)���?� E�kW^!߁n:c� �B�@�QQ�`����tph�s�cV\�QO8i�p�hD��?��"�UP�ULT�:���-�g���� �����	9��l_��z���z�f�CQ�"�QD���|V�b�H�3�&f)6#��B=#+H�}�׋�N���e�s~�ٴ�hŧ������<�����v(��PNHe�Gb�}���Z�ۗ��b�ͫ���~��d\�-DF�^�W~`�A�IRL�����'�$���6� ���ϧ��7�W�kޫ���{��m!3��2�
fG�8=�]wUn�-��)�YW�o�	 ���M� G�u�ܻ����� o;]c�����UT"*lgy�4� �*gk=nے��Q���v��l�.X!�r�;]�(Ǥ�׺,��_0��R��ݓ����=�v�=Lc����]�E���q]�U��k����RL̪�En��g�C@��A��H����%^uۻgm��s�z�@���4ˎ��@��ʩ�����-�3���܏o( �|�h	@.��E%u5��ڳ�g��&�QQh��TQ24�V�4�d@��j($Fz7��H�W��8q媟[To����3����S&\�J/Wٸ�W����z?��zώ���R��-lyσq~W�M@�^�����������[����3Zi� ���Zi��N Y%I�?J�mm.�����Ci��BȊ��o�k��"^y����7nUI��|��$��[�3��2�beLݓS�X%%����W��sk�'k5Ҙ����~R	S�q�>;}֮!�2cy����zy�_O���$L̤"m��`�{О��9v<��	�ǵ��7t���}}Db�QTP�*t�9�i�� ���?�]����ǁb/��9/����a�J�uv1E��&D@��+�S��`8�w��*GW��<�;v�`� ���7�	�T�\�u�=[��u�=�M��4n�д������I/�#iv�I%깇�X�Sq�27�@r��6DFQ�r�{C�z )U)Q
��u[Iܠ�Q`ㄉ�wn@��9�Z=͵j�y�v�쨄Ysj��n���݇>P�7�[�9���g������k�3�v�*8.O���.��~�og��GRyE�@vq�W��}���H���A�����E}Dͳ���ڣ� ��?Zl3�3s��L�'�k����+��εp]��{�Q.l����QQJ	SB&x؇�&���X�G��5��I�fP�����~��tD��U^z��}r���޷@�@|��Zl ��ʪ�Nߴ�fb��dDvWmC	u�pc�TIf88����|ZB�y��[�#ޘݬ�u��RH��p�%�9�$�~ߊG�*4Us����{�S9P3*�QA�D�����{��E��J=�ڪ�S���^}q�OFR$�=�r����z!PM)��S#���������}���vԂ 7-[A���b{C�׬�Jk��4��KHR�(�8�µ��r�m�u�9Q���o��wμƂ E�q�� ]�0��0x1/)z��蟟��坉T�4����޷���ar�Է���4no������9�:O�Q}B>w�Ǘ�9�ӍHp�r0~mV	���=,Ǉ:O��� ��}�E��ۍ�[r�eo��ٷC}�'��_E�1~;{����%�;�6*ƴ��׽�;2���I����[g��E꙾�=������=N�J���{�yN:�Ia�N)�4�<���=4k9T����	�C_����g��E��h�;�/w��ś:��}�r��m�D"�:�%��Q�pw��:�T��o_�w���k�.&m��s�����x��pӋ=�V���_����z�{�do|�Y�Z�{t�����&�瞁���<<���|}^�s��'����/�^�;|N���yz{*�ǰ�c�g����*�;�x�}�LRc�HJ�Chs%��;��x]�c����ǸL�QU��K�������;5��Hq��+��><�/W)�w����n�Ff,]$6g��&��X\'�F�oq}�q8.����o�����~�|i}r��xH�ޣ}����j*3��od�R���{���_uG��G�� /�{��_����c�;~wj������\r�f���E֯w�$w��D =�|�������9��^���l�5}޹f�	�������A�7p�5�7��	C]�ݼ���w�9Z��у^��}�D���O�yf�(l�wK'E�W��o�R�#����˚�{<�㛌}y��Ƌ����E��w<��f�Q�^��K�(B��0Ƽ�'QE���{T1�E��m�
�ۙR�aR���0�m�z���sp*K�J�n\��Q+SR��q�e�(�U\ef5D+R�m�6����ɖԳ*��(��V,�px�Xk5ąJȌF��qr�(��2�-J�X֩Fփ��eh��,�L��eq�,�E-N�]�R��"��(�(�q�XV��U��9\��ƅp��[J2t���u&*&X�.��+2��e��"(���!�f�6Ȏ��L���XR�.�+lu�Z���TUA��h�1[i�ƱEb&�k
e������^�Ŵ֥-PPb���ڣ[1�Ϯ6��E*WKCwUP[iR�p��+T�j1U��ũc+PRZ�aG2ܴ��Z�p1m�����\�]n�1�`���K�Ī�!��]-�e����?�yy�\�]��=�Qq��F�����n��Y��[rX�t�\ss�4��;r�M�m�ul�v�pu���W�bWd^�S����Ѵ����+���ͺ�2
h��ny9S��������9�9��.����3�wf����\fKw=k�zg��&�G��<�x6����17�7Vw`'�#t��nMk;��vk�gllN�23KnOd��T�Y9ҷ[�>ۇt��&�í0�g�Ц-;v� \c=6��ka������2��!ջb��B���=v����F;LȐ�z�ڧl�����v�5��b=�762Q��/"lq�v 776帳�j��=�ްwn¦ �G�����=�kx�N.����km;��N,'$��Fא����<fw��l�kv���v��k�������n�u�σc\�l�s�<\�=�vktn[��Ksi�fs�8��x�v��v�^ۍE�U�b�Փ]���0nxr<���r=7a��:�������N�\���Y:���]8v"�۞ۣp:Ν���8�d�0l��<��{y��ڻ��u�Gi^E46��{V�]���:�D�����u�W��\t�/�+�v��6�IAu�h�豻���#nuu�m�//g��ѮN�`�;�M�nM���ig7l:�p�ǎj�71ڔ^r�U�w��;��<W6`�=s�[���r&��狄��S��@������6�q�ݶ���.P���'7��:M�n�pu�9���<��/'������m��az�nΉ�.۟g=xدq�]On�Z��^7�7+1�R�vK<[:��]m:S��(�yT �7`5p����M�G�����=|S��bƄ-��uץ�!�]r{plv�&�u��swZ1��9�n����hvٷY8���T�,R�dn�7U�\��m�y�X2E�qj�-;7'oM���:6�fN�ѩ�Gm�R�9��<����>;s��c\1�Rm�6a��X������Gf��\��4��]N+�r�g=�]u��G�j�o�ww���-���n�.��u.7k�:ln���,�t��=����p۲���5䝜l�\mv�磛v����!��r�p��q\��<��)u+s-�j�S[E�u�՛2z��8:3��-qv��h'�9y'	���d�]��齼㈒�.����q�]�(�h祢�ap^��m��9�[�t�����;O[E�Yz�tb��Y�n�oe8�]b{\n��z�.���9�ܛ����\�sn\f-��Q��������������L�������  _}�M� |��Zl$<��t	T�:Yٳ���M"PU��i��B��((2f��o��.!V�{ӥ�z�vԂ@}�4�$v��6��,�y�u��˗���!t�~�'��P�*urxgoZi��zհWB2��g��9�a+� ������֮ndɊ�*fjH���8����\�j������m4��o��i�ԄuZ�쟐1cwq$����HW�(!1!`�'-�]2�&7'm�#�t��ry����`{�֛@ z��6A���cr���)��J��?��=;�ɷ��ۢz.��N��W����OD&`��bL#>��%)*b �
u�0 ����3�>Nmkgs����+�#t���(�	 �k_�L��QL�0%H��7��+��`�C��CT����5�>����0�/w*=*���fǟ��;�sa�i^��{wu{ǲ�Orw�\:�,x��oխ�{?�ٟf}��ݛ��I"P�[�;J�����"G�Nztn��}��pj=W�`���
E7�o}j�+6}nO� �qo�z%�U�8 ��Z�����լi��~�R�@�3B�<l��d�N�o�}�}��j� 
�W��A��Dg�GU,���%���_�a�{2!`�3T�7ό��7� /s֮�w��ߣ��E�f4�
��p��S'��֬�����=��je%D�@(L%�2�ݫqV��E9���a7�;�q��k��)���_|t�AP&L��&򮸵�K�sf�i$�ns��̡�1���ƍ��x�vP֊�$"}���K^KJR&T�A�w��k��� ���A�wv���a�w��> O�i��I�U��D�=��Vz�]C�Ǻ�&Q� qJ�������M� y�i������躧H� �׸ߘ��>�zJȎh��-����/S������߼h�=����L{�;ﶇb�Xb�{c�����o����� �7�����HF~�d��.{�Q���
�L�҄J��j���!�>�~s��� 1�*��2�{x�c�Il=���)�$5={���%��`$�ɏ��e*d�3e����X�W��j7��M�m�6��%��UیQ-%��{Ѓ���+Q^�������l�&5�.�{N�݄�n����ڌ�;Z��q�h�G"�������t������+n[	 �5���I/��6�[~�N�dܙ.}��"��i��zЊ��AJ�*G-���1j����������ʶ �2հrv��$�ю�f���J�:}�H~0�R&Tb�N��P	{�
i"D��h�"��͏Z�K��	 AW��Q- _��*�nD�q���'��^��b��ݱ�_��M0 kܦ�H�';��<�^Ų=
�j�D�y�~�4Gڞ��b��{�N�B�3֍�_����pK�����śl�zk���.ǽ/$x�Y�>���������.�v��A�
T}0"T7i4�~�`|��\G�ͬ�M�9�.�q�������iNwM����{�y�8w������0�U��՟E�34�����h�Q����Ĩ�J�&���oI�I��$�R����� �t����ۆs9Uʑ��:�u��mA�{��3�a���������|���6O����ZL�Tv�s�~����> ��ˈ�Vn�$���܉��H��T���&�h �b�*���1�m�
�m[@ ,dk��k�sRA$�y��h����2��/�׈ƒbD�P�Xv��gG���Z�vzE��&����@$��i��I$���ٚ'��h��z���i�C���Fg�&�
USH��Vs���|Aw��1���Y�>URO�����@W�Ɏ��ܽ�ƅ{����y1���S�=�4�����-�)�ǎ�t�sr��z��j��Kg=�p�?w�{���4�<񺺳Dר�a ��zv$�!�C[|��r��l��cw�:�_e�u�b�:Kr���q]F�%��Gi;8�7=�v��X���{�KO�q���џK�F�m�x�F����v	���������{z5X�=�nv���ŏ��ֺtn�jok[u%s^=b���S-�4b;nN��ßs��q6K]������p�pYݑ��� ���me�ܢ���m�'F�M�Mv[n��n���88�&���<p.��O$�&���Ѷ/�v������vn"~�SD��E��� V{�l �/r��gaW9��*or_̃�+3-�)�yzL�Lɓ&!���qm ������yv�1 Ow-�C������g��F�S�rW8���݇�4T�J��8�޺o� ܯE�@|����.������=� O6�"- gk�B��2�
f��L��ᥪ���h��<�Vϯ@κ�A|�l[@ ls�������	3�U�2�\8�CI1�*��qr']8�a��w��g0�|��r�
�yn"��M��ɸ���:o�ߜ��{}��`��������Ҟܾ�8�97 �7��`��p7WX���������ﾱU4�7N��f��/��M����%��{:���K�r�8��5��ky�T���?T��y� f�_ʙ�B�ξ���'�������]Ŧ�*�De��4i���ɻ��!�h�;�{�鯦'�X���,?xNug��#�8�v1�y��\��_������y�D�I�o��6 �?����/�|�oo�1�"}���f��"A30��M0�{�Qa"yfۖ�I.�������6>H�Q�ޠ�����p�K<w�0eLJFeEs��ٻ�܌�w���@ �w��`"UǺ���O�HNl�W�d���Eq���i��4��ܤJ��$�&b4��:`^��jG���[3ܵU|�8� ��M��=�K�� ���Zw����t�hG�f%D��d���E����[n�l�[����m���iB�#�������ވ��J�P�f���W�p�rm��O4�[<�W�$*��ϻ��ޱD���%�Uk��r����&���^��b	f�ݷ[>�E���I��{�[ �+=Z� b�ҹ�ݞ�b����j'o H��&>�*��I��1- �����!�>{�Dl1GoZ��u}��Sq�v��ob����ւ���6g�H}p�B�rn�s���<�.qo�S��ê�ȁ7� >��7v?~	$G���[ 
͟�DN�ɡR���TIg~;�֟���T���� AGz���:�H����{�v�t/ �H'�^x�
`����@3t.��>�lI$�ܠډ��&���哿\e8lLD|��ֱ�>�wm?�u���U:��.ț��?�is���u���1D�dGi�65��j��̽/
���������+�quԿ��c�����>��D
��i��{�����*���)%=��4�?"�LH��;
z�H%�L���3�d�����KU��(��[ۨ���2��Xg�6�|�]�;�ED��4����N��> /����"�ú��o:����\�P�V������L>��vi�d��%Eݤ��
�oOT�wMO�Z�w9d4+��M� F�{?Oj�͜}������k�����מ�N0.n"��J��yG��N�/���v��Y��<�a]���^s�$�s���_|������X���H3�DB��U �u���a�?~t���{EID�;S�߃ܹv?�"��j� ���m.}Y�B�*����	A�*T�b$c������&���-�6:�c�\Ȗ�k�okخ�ZH�����T�MQJ&TVn���ڐ /��W�_lk�l%io�c��~�[O� T��8���d4�)�UL�h4��Tσfn�6���q�o�  ��Z�� 6|�_́�Gx��62Z����V���LH��;S�l6�I|��|ĲPK��=~�r��|�gzyx$I��Pa�
! �:�6��#��bf��T8�9���Qܪ�l���W2�L g�e����]��y�*n�#;�^�\5��;�J&����UQ=�~��\� ����2]�����'�э�δ��|�OK�hͭdD-���%�qYq˘���*��̻��1cR���;�y�b�{����f���Z�x�w4g��&�;�:n�Yq�vR�;|�p����G��}�h�#n
2"I�=�m��ϛ���A�Wl!w9��7f�q�D��`�v�\Zt�6��방�7Hc��}�����w]0�*���Wp���R�,���6��t�k�a�Y��۟i��Wl����[C��������[=OX��[�MW�zvۺ�8�n���Y���q֞6v1m�[cu5�ǭ��r-�Cdn��*]=[U|籃�9����#��m�k�n�&ےѽWI�s�t���5��F�邂UEB�y�`��/ſ��y��?���x��T{s<U�i�ƉRFd��L;��
Q5H�&n�WEV��6/�}Uvsn;h4� �n���A+ͭc�"=[�VJM����nm#12I��I��pOLe�'�%[�ԋV">��S���,��� �����>@|�kX����$��E�1�Ћ�#�bW81��G�[;攱 �����4 �f��;�Ѥgg��'���i�̓P�̈����h���iH ��O�c��${��V��q���` �/٭?��=���������O��qfO5vn��������������׳on͙B�������1���U�C�y�Kz}nC�T�.�Zm}�/W%OVVW�yO�>읱��zH��IQ?ETT cG^kM0A
���~���_���]�8shT����b�cS�#ƤVxU�g�:�9��1T����т,�4S���݌en�E����ٹ��ALW���W���h$Jzy��"���3��F�uG�����x% ę�`@��V�R8A������^�Hw���>���` ��֮��zȩ���ER���,6�3��ת���w�vҐ�"�kV�A%��u�=VlM������,4�u��K�C��	��R�M��;v���I+�|���^�z�tY�C��I���$� ׷[�j|���O�q�����#Id���\r�=�pk�3�c��؅ꔎ�,ȔT���+��2�D�p�[�?��A$�Z�(�>��G�w9����� �u�~���I1(ɏ�J��"��
&${�w!��j�g:�t0���޶������9�.6NV#�;�����nI1*>�*HJ����0I;�D|(P�E�V\H��5��)�*=4*����("�Eef5s���`�F9Ɖ,�B�� �3�O�ʇ���N,L����8:���$d��xB�_g������3�ږ���4zI2�'��bm�o�&�I��jF�������ϼ��{B��JǗ?�ז� ���?yQr򄗯�vkq��/o�����~Ẁ�~��W0���=-�h���M�j������?s��ES�ɝз|>���ڳآ�����=!�Rg�nN>����X��g��kΰ��O�C�H��zw&�����9�sA�gz^�L��`Aj§��x�o�̒�r$�����Ǝ�mL.����ѯ����v�^�sw_�,���S'{��W#3QD)O��]�GoMKz�z�\��������w>Ԗ�"ƙ�E�"C�5�}�2��m��d-%��]�Pk%@��,H��i�@y��z,��Λ������Ϋ��)e%�c=Ȏ݃�,��8�Q��gc��k7�y��S����{��������d�o�����������o����vxz��T���h�����a#��ob�7N�۞���� ߚ�{u���ow�(w��/��D�"A��#�a��'�����0p��	�;��/���g���ɪ��fA�́���'=4����<��' @�{����~��4�=Љ�;����Ըy��N�@�l��δĚY2�ʾ�V{}�מ�pq���f�^�{;����J;�Y�����p ߩOg@��V3�8X�ㇻ��;����2�O�8| T��}�Ꚛ�2��Ui���%x�D,Ӡ���H�>&9��<��)����)�.Z��B��*
��V)iKj�E�-%e�m�ʭQ���5
�e�9�!��.R�w5�JܵU5�Yn��U,�0�2jbe�s*�Fk��+na�0��ظ�]So.渢�Ӟ��ɎS�X�e����0jje�ѣSR�����bW9���-EZ��G,�e&Zax\��PA3n �g)V"��ڜ.&Z��+�-�Q���`�-�DYX#����(��[Kh��7X)R�j���Q�8�-m˘T(�Z0�̲�h�*J8�S�\�%k8��/6�31�Pmҙ�����˂�kY�0jE�nٯTĨ�\�76\ov��n�һxw`�8���'�cw���{8� �L�8�+��^nf$�D��Z��Qy��6�b9s�ں3-��TUyJ3��n&[F
2Ѭ�KT��2\���� >�)�������m�'�M|s��x% ę�`@����z���z#��A��m��4	���]	�#��p�I��<��D�V-Z{�d�u��'���=���������n���$���Ă~����1|=��b]k� \�pu��\�3&��7/v��qs�A��=oog�{1qԻ60�ӎܮ���wo�.n��W�|�;�:b��l�&3�)����e@��w��$�ٯ�" yj>1!DH�-���o�OP��DMP�c�{�k̐	��$���˰I���V����]��2�{�%)&L}0"T6����f�$���[��z�FG�����A�t�Ē#7��&9/zI�Q��RBM�=뼌���̐Gn��~0��L�+w�
�w�?U�UU���W�1c�/��˹�����6�}��o���*6>��g|=�v�Q�������]���O�|�}������~�{�Y�3?�����'�u��>|��;-��1@��~���k�����ķ7�Iz,��D���I��o��MB�2;/����	�m��]�.��B6��l�g�<�m��,�s�v3�k�p��-{�����\[M�'��^�$��ݠ����L�{P�t��gՃv� ��XgCK`S&T��1���AJ�҄�(M!c���1��lEn��ˍ���[�q�D�J$D����A��� ���r|נz;�,�c��L5�����{�%)&L}0"T6D��-�G<�W�"��={ZH$+ۍ�A���|}ڶmFU�l|L�%�H11L��Л���[d�'�j����
"+2o�Ñ!�{[ �����`�	���G��|v�N!3�َ���>~�喯���x7���gu�b���{t��1j�>r�{z$#�	~�����?~B���dz��u�7RE&ex~�}��J?}�_c6��x�:u�@7��CoO(�C�۞��S�ꮳgxԇd{��7Y]�칁zgv�(k��f3*�Vq�ٝ�Z�֏y^���R��e��A��#sK�j�̇n:���9�p�
"�Y�$�Lm:{i,5]n��u���A��t���۞������d؅׎e;�Lx�_>87��L�4dId�۬�bq�l�P��tV
�y���+�6�� u٘�ۮ}v�v��V��c��8�l�uȶ�����߼j�yP'���e�cwv����@��Q��gzjwTo�o5������ïv�bfDI3&&0}ʽ��9���1�np����h$����m�"v7�A��m�ʣ>�S�՚|υ�Pb�%*	���o��mo*$�դl�}C�1}�`�j�[D�o*$D��DIJ$D���oz�E�L���3A �s� ���KNoS{7��xx�<�ș��IJA�)0f1Kv��m3w�=�u[=�=����������$+��_	�3}��pz���~|�/\�����f_O\{O����]������%7�weP���*}��ݥ2Q��Q����s�5wci���}�g�,��uV�;]]A�g�8hx�	H3"f(�~�����}~�18Qbx�k��#;j��4b�l-�>Y�X���O��o7-=��=���{��1}�t��'��S؝��/|m����/�g̑9Ѧ��O�u��`��������3[�ԢfDI�&f`�j=H�M�v����x��G��]�߉�zx� ���6��[bfĥ�όu=�	N8�B6�߈��t ��]��A ���QՐ���{:h�1���J*$).:^׉$�vQ����*n|��!�{h0OƷ;�.�7�>����\(߾JDDf L�ѳ��dǞvF۶�g����I{{���ma�<�M���~��ʃ1����"k�I;��N���;kP�HD��E�I!�g0�	gU��u�H��A;���tB;;������c��O�[͒I����>�����S9��[���o��R�1*"�ך� �"�w.�?du�풉g�2ߔ3��ji��C~�����T0��S̥�{΂v�9��[�X�,��8d=���x!�c<���%.b0_�|>�w�|O����lGƿg�a׷Z1"T�"f3�Q�z�o6'_���}��﫾 �+ݸ�?ճƯ��S�0��`� �����r��)D������S�� �ս�;�>�ȍ*�蟜_s����;[<h�����y�MX���4���	�Jb����<Y��I�z�Sq5qv�Ɔß��������Q!H���~��I�f�d���4NOn�V��wV3M{�$����dL% ��L�3�jv:���t�Y&s��-��:� �+����<hYxw�b藝3��	�VN�/�$��e}
�V��v�i^���슡4c|�3ϻ��H5���T�7��2�1*"�O/�ݏT�����C�}=~���F�$��o�ڌ
} ��Fz����s̺=J����S��T;�`}R��BT�*"����Yw�cV�M�7C���k�i��k�=>B��T���z��N#�ؠ�����߀'�y�������*B�13	��O��P7�����'��D+���W�luF$^m�`ǌ��}�Q]���,/!332�
%㹭��-������4���$^x۶�hw���Z���ɑ1&!�7�0~;ꍯ�$�̓�ц�j��b{t�Wy�~'�z�M|O���3)(��D�%���&������ܳb��3�$�Ta�H$7�̀Gʣ���h!�[�DD�+�T�f2��6|�6�$�y�L�I��F�Fz��d�s'�Oz� I!��l����D�_J���s�:Ю�\:I�äI'��0H3���>���&�w��@���A�&�!-��kl�~3ٹS������ǖ�&��	��{�� ���?��yΔ�O�C5R�~���^��Y����k��'�g��}0-�+��G�颡۾滺��:��t,��u���;�=�=&��w�eٛ�n�ݓѬ��q�ֵkq�rݐ�Mfnݵ���#�u� ��}O0�����e���:���23��r]��^�D�;uv���tڤc��X:�$�"Z���W���0�.ַH=���l�Iݘ�K��$��3����v����5�B8n ��]���(m8S�=�m����5�/���ui���Ô
ե.��X���@��c.ۯM�6[\�šH�z�t��5���Z��f4"Do����ɕ!L������-�m|�����fa��Uޝfoá���}�l��0�J&$�#C�o[ �Ԭ��O�l<�O��[�͒I���`���D�}#j��【*0,���*"A�2��r���O�|�"�wЖZ�Z�K�n�@�nuI�������?)�LL	LmLtmtOJ��D�{�2A���0H�T�z:o��'9k#4��7�l���y�)S̯�6��(0s�m �k����}j�������g{|�':��qw�_>��}�?����L[�`�R�����9���j�HlOS��m��QA_�������v�&�!=�;��$�;��?	�6���w~����������[d�O�{;����T̙�J`��T���z�m��?/_`���d�K��}�p��*"1�%G4�No$�K�6��0z����<�}�C�pOn���zW�96}�yo/���|?:��?|H'���6	 �ڟƀ$�M�MW�!�ɑ�fk�������2�ɉ*a�sx�d�{Q� �xz*v���	���W�v��D�J，�P�>`Eo��N(��Y'��	.}�n�A�!��f���Uek�Y��� Ú�N�����0)�*�/*:��g3���o����L�����Q�P^wS+I��竐(�F��@ĩ�	D"���]Gks����uv�fN�v��%��l��?��>�q� ���$��w͒7Uj�H$K����8s"C�]���$^�r�z��`�2"
�K~�se����q��9��r�uB���(�H��͒}��3
��]��X�Z*fL�%"̧�G��@$��u?� �!���W�V{k���v��rXqҹ&!U�ҹR�A�yK��6U�X��^�I�R��{�"��a�u�[�Bo*���F@�z��z>S��� 2�����Hs�	�o}��H�;ZA�&LIP��uVeF{/o��@?z��&wٔ�g�|���*>���W�dt�+��J�&�o�7�'�O�}����b�P�{��� ��g6O�V����)�^�������~���;Y�m�hy�L�4>�gn��뺝��l��z�b�[vh�,�g��y��0%w�N'#v��k�|��ԃv=��#鞑@�w��?D���SbP��Ϸ�2
@�3,>κ �gs6� �G{|�?m����ݒ�I��P����o����0I���n輁\/r:��?'o9�������\�	L��IH�%�������U]�H3�L	�fy�I����>��]��E���Bx����R��FLs�o\���-����yw�1�Bt����Xs��ڟ���{=j<�����M�O*��s,VB����  ~�H���9��
 �&d(E��og�~"��I^��څ|��&ns͂	����A��@0z�ʥ�3 ���"���AU�
��p�x��ώ8��La��4sT�c�mk�������Pb&S=�{]�A��m��#�zE,"�@r��GF`]�� ��[���Ob��&��vC���0��6���=����A��� ��k���BGxE�v��%��f�*w�	RT	�BJl���������H�>ҷ�����^޿���ks���յ�D��"R�	lz�9���X�� ��|H3׾�I��b�O�����O-�K�yQ��$��kg_cL�0��
&Kg�{��ٴ�wWp�[��DޝD��6�?�U�[�,xpa�4;jtL��S���_H���E�v��i���� ;}���7z[�}7{���q�u�������O�_oX�}��z��ʼ�q{M���Z�H���ޣ�o���g_o������r���7C��!> n�$�;�v������G�M�o��6�����>'�xɍֲI�O�EUF'�{&DFt�3c���x���	��%tW�i7K#w}\9�,^��9����°6������A�C�;:o�/��cgy�����_�{K���y&/�����I���!��]z^��ַ���7-{��٦��<B������U�6o��}W�uh%H�i�O��h���_�7�X�m^��ҋ���Әj+��zn(��~���#W��۷BhUV�� �\%���{O����{R�׾�>��а��nJR�w\Zi,&���0G�9�,l�U��^���wu�6���e�#��{�&�X.dЃ��hGq�/8���%/=�'�|��ޔo����om�s������L��7�ޯV�~���Zv�5{�"´|F���ȉ%�|���r/`�k��ļ*�ۗ{V��`�|�;�/Zv��IΔҾ��*l�"���G?\�n��z�_,��j���֧}��-���g0���o�s�S7�����D�W 1r�w]�
g���<9D��.[�:��U��s:�ZVm��m�H�or�s�n�s����9���׻yC���/�6���>S�.�{u���~}��Oz�>y˲���㕐7���h�����G�u���.�ҷ6�m�]�n5x�w�f��F��8�m�1v�GiZ�[�L��x��X۝�\q�[�<x۵�} ���b�0���
�u���E�imv�]����&��0*�X-eZ�@�7�;� n�"����RE���\L�0ģmq�)mmV�x��X�R���1.\ULj�qrr�
]�����
�$R�77C�u���."��Q-A�w2G���
*�2���̢񨦴�c8����-]²�aJ۷��,b8Qe2Q�x��[mF��sR)b�+�b���[C-�XnW1���PM��y��KJ#�c�np̠�����*+�S]R�Jӌ̼���a�1��ժ�+R�kR��
"������ԦQm��	���cnm�{c�G��䖖���)piU)Eܘ�j�U��kF����W�W[��yn6�ʫF�h��n��������������0��mj�h��Up�9�Ӹ�!&�Ǵ���{����lۃ71�y��0�۰=cj�c��5�������܉�n� ��s]<��^<���^c��0gX���x��Z{-�qř�kjM�8�wZ�I��-����n�uұɕ6�.����Zݙ]V�F�T�����|{��\�����ûǘ���R��nNۑ-��Ֆ�����2�Tq��d�mǣ�[g8r#Ë�n9��rrg���e������Wdݍ��s����]&�ny[q]]�놟I�V{�4]���bv��v�kv��#Q��5&ŉ�vDѵVEٝ���cb�����h���kv{���q=����#���Fq�z�l��qi��̊��2Q�o"n�.'�kG ����v6��&Dd0W䈻^նP#���-�F��1f�t7���c��W[X���<c����uύ��[ɹB�[ݒ����Y�;���.�-���Ҿ����3g�Lvܘ�-b6��-��ɸb�۱J�����n���"���j�k���n�i��qb]x�۱$��g���Ջu�ٺ�1�shN�χ��|p�;��v�}�rXt6���C��9�n�B]���%n	����6v.m{�Mn嗖ݯd�:��x|��UVӮ5�iMV���u�<Oh��T�m�	��yJ/PB���V9C���g��ֵ���ӭn�^��w����E�c�'-:=�[j��n[uy�ͣY��C�m<hܶc�v��un&x�X��ݺq��'I��{
���3Nԝq\Kb976ҽi��W\;��w\�n�]\��X�Ʈ6��0���Y�r?�;�=�ջeq	u�ձ�E��s�����Nݝ��q��ձ�着� qƬ�fآ�c��88m�y;aw[p��w8�nJ�Fs��P�s�:{�Dn�K˩���˱�n2�'������q�n�u�q�\�»�:�b�vwV���n/����:b.[���卸6[����~���������պ�)�.ub��cy���sonN;3�V��K��
L�{Hl�F���y���tI�����v��ţJX�s��i��9x^q�k:{.K��p�%\]�[IE�]gm[��<��B=|Un�Ms�z�{/�-�1.���rv^R�1ݳ�v�7]�����>f���9�=��mn�����xL����TQ&��U���f�n�^�4m�u�m�c�{�����x����호��sn�]h3�����"P���a���o̂/j�A��sr%��=#v.���^���_1�~Q2LD�Je����H.Ay��СD�>��g�A�U�W��w��~>ɓ�=;/7��]�M�zBS�L`Jb�N�ď������7^��*�Ow���7�Z������ ����*ġ%SϷ�ݞ��?m{��3�f0����O�!�#�Ή3K֨�.�F�Qk�gk	$�f����w*�*M�."ڠA�ws�$+{|Û�N��~���xO��v6�O��.�n#��-�<�+A��mG�`v�s��E�������q \�2{���� ���i�OĀMoo���g�^�o�[{X��$�9�cpz��"dDL�)��7��?;�!�U:T	AU���q���Vzڻ�&n���x���gZ�QԁI2��|.��֛�����1�\�˜�1����������A�;���OĚ������ͩ�<��ȵ��1џ�0�RSMt�a�I�v���?Xq����/s�hWv��"{���0a	�)��W�<�0맰	�=t� H%��6O������	]���ٮaĂ��	R�	FL�ٯoy�Aʶ�o��x�ǲ+�	���$��>�W٪yg�fY�L�<L?��g�;ٞ��9���-�mq�i
�iI�s��&f�����&�f@���[�Iכ��������xOoO�Xd����׺ɘ�T"�B��L�/z�XAw��(��:T
^����A ���|��FtW*$����b��#�������%"dDL�	�o ��� >^��٨U���D���V�]��
��z�j�A�����^��x�	5WuP�O��z(2{<�(|Xns)��s ��>�^�dY�W�� |��?����~� C?L�5�"�,�|TH����v+��������u�V�ĀWKm��'���k��S7��φ�H1=��NyE�0DH�"`J��c�>@�k��O�n�o�mX�vg�k_�2uN�@+׼�S�bz=,���Q䎭а�����`I,�%��j�\9��p�-�m�)zwvz8�d�ϯ����t@�*��{��d�Q�>'�Lto��:}?D�	9�8h�0�X2`(&aD	oל�d��xa0}�[���	��S����VQ<U�g���=ߙ�o�ə�T"�B��َ�x�?�gS�3"i��*5�8�;�h����{̓�6�!H�
"J	���W������b��M_v7�$�y����Δ%y��	ؠ m�T�<MU4q��1�E{м�T��-�RȊ�!Y����/`^��L��N��j'��ee���}�~ �����%�Q����2��q���� ���0�N���NP�������v��`�}�o쬓{���⌯	!E�
B�:X��l��yݎn;tv�]4��[���jX�G+�v��J3~��6Q�"$(�`J����4����� ��'�o�,��:{�����/��t���q�H�^�2���)�^�����1�i�l�Ă�H`���a����pzk�t�k�{��=�D�^�	�Q[�{[A����_+�_�T��y�A�'�|�g�_u�(�EH�&�~�]ϐ���"��i�~3���9�<k�&׾��#]���������2D�/��Y��}Q����*:z���4�͂H���FmO�����l�(��f)�l���$�{o�?�����8T'��g�lwUP�nҋ��L17�/2U�mcɉ�(8N�7;�y��nЏ���}��`�<@԰��Om�)�\=�8��k�%<����;;���6�4��y��]��)@����]�qm��އ�N�z%��z$�rb�7j���	�軜�nK��8�$G�����x�ۮ�n�m;);����n�q�u�����ې����M�����W��z�;��r'`'s�6z�����]�n2����ϰmT���d�D�U�ns�!1�1��c�]�:8v���9�Xޞ���/R�5�ډ17����D����"����$c۾3�$��4>1�yO�F
�|�:�c���ȉ�G�aD���)��GP�a矣E�O]i��m�~Ω�DZb���{�`���t!I�!2��=�3�?ꍯ�WFǦ�f�]ǺjwH �n[NuO'<��$�$�3	A���U;0��ٞj���A�|�d�H��\���;-v�O�D����_{"���3!(��B����;��@�{z��wu�GQ��$g��� ��N$�u�6��B7W�#��ft�&Ja�+X�5�;�;vcU<g\�k�{mhB��YE���ՁH�
`Jy�l���Mk�y�H��;�Y��~>�co���O5�w�DL�34���`�����A��]۟Ǉ%����'�U�G��\���:<�^'�I������o�$��Z`�4���{{BZ��"3��-/�ޚ�����ߦ�`�=�\��E~���$ҟE�y�+{n37>d)�L��
B�����U�+�v�$������������	�:��ަUA��A�J0e7���/I�<ʵ�yo�	 y�A��r�=��s�s4X$Z��	Zv-�� L%[�ݸ���1����;�;�k4�gۓ@	����$�Xw���pT}�R�
ą	Lm��=o%��+����Tk<u�V�YT��A����3(�F`����P�D8�m0H'�~���zژV#��ܐb�� ` �����c�֬e�(lY����^"�+c�#�,`��� ��]�6H'�=�m��)Z�px��ǔkS��5�w�DL�3-������gݶ�d���9��t�ۥ]~��>�⼯'.}�7r,������-���~Ѻ�ǺH�(��
�s�靂j�,���g��A����#r~$W��͂I�~�l�ޏL��
B����u�;�B�_�bkt�e[�	�Oս���WN���%)�J����_sd5y �2bAQS�ן	յK�j��A���d�OƯ�ېQ'5���}�}�2�w�/Y+�mVz��M�m u������=F��uq#ڝ�^:&S1�)���2	D��&�;�y���vm��$sk�]]u���4��z���n` |������D!fO�o���0-�����S����>� ʾ�l����)Z�~�**��#3�%)2�%1��LF��E|}�(��9޼�I&��m�H:�hP��Q"bD��l-��g�y1���*�3�����}ճD�Y����}W}H\���"@J��� �b{����s2�m��<�;���`�jCu�12SX2��8��}Jfo�De�X1����ۊ�X���ي��}��&y�6DOdzd�@R}0%?��z���^��O�ٞ��V<v?���m�I#������o���{��ߢV�|H�翝�WZ����nv��2�nܠ&��u�!��n�زJ ĕDD�ҳ$LH&!Lo}����;[_	$�f�� ���Vd��{���0~:}Y�9^��g�	A��}��<���K�G�M�d�|��+�~'���7�A(�(S�棷�ޥ��������P���S%�w��$k}�A�K�7�ɚ�;��metPaͮlez��� ��M@qqq��2ņ�`'�Ǧ�� �~����� �v��*}�һ�!W���H���%��Ukd�A����=v�*�0H�Wq@�k��l�Eom�O�����hD�V�5p�!x���8�[�����;�o��([��1�p�)�ȋ���������-�;��be�;�s?��sU��ns&bR�]�mK��ۭN�ծ��5;/v�秌�ny���&^�ƚ�vs���6�,p�uh]Qa�t\g����u��j�۰��ʑܙ�s�����s��uC=�X�rnw$��:ི�Z{b��ch
1�Ax�FZ����[��Cfa1��CӘ�]8'�v�g��m��%M��hw�K��OL�6ե*���m=�0�F5n ���2�g����n�5����1m٩P������6W������v�u�@�^��d���`�>���ְ�]~��U�E	����]} Ȕ&I1
b����d�ϼf3��{�������lH5��A�����v��s�F�7�0�&~�&�v�m�I�6�̂J��:W!���E�	�g6$V��O�DP�(�2"!L��܄j�{��c��?�ܠ�$[��`�qutS�Odw2"ݟA;���=��EA���E&���0N�WT��qp=���#޾�H5��?�?�y��
H���A�����:�vZ���.���7[��ZSm.�+U2H1e9�phF&L�H�=��Z���	�����I���4Wz�v{���o*�$~���3^�D��G�S`�t��i=݇�asv:�q��T�����[�Oߐ�5�=@�r��>�ms���OLgz;D�&�gh��`����=��h��໥k�`E����S�ē�߷��8~q@Κ��\�Ck��~�¼��J$��1!�>��A$_k�?$=�LV�L��H3��A�>9���s��b
&~�&o2��{��v����@�k�L�G�ە5�$�z�0Px����%�Sn���)
	�
d�G_�� ��u��ӽ���Ĉǘ�Ē��hKy��m��#V6ft��9O��^ˢne�4�%��]jj:�]��������d�f���빖��||�.��ԷӁ���	�uD7{=@��ʝ����9�|��r����312T)�\� ����C%��yh��Z��Ov��~'�y��$���ί��|�����I��0T}0%0�_:�����`�`}Bŋ4Xy^��Y-}�A.�SN̹�Yڭ͹���l���7/����}�;�9�����g����~�{��{��͈a^C}t�}lC:�.��@t_T�>��x�M�E���k:���u�v{cq���W�twR�`����|��c%��(�����_O�u}ܷ��} �4���=��a�x��B㧅5I��#��n�������!���oo�K��.w�ʘ}J����� {�E��e����4鞞z�(�V�{٫z�;ˎ�_�Iz�
^��؍
�����eլL���e�/6�I��4ך�to)+Q꫍�2U�`�*g�\.<���'t�˶�a��nO�j��ӡ�W�l>�q��"�ΰOb%?=�r\.��|����&c
��+�ں����}�3�ۀ�"�d]��7 ����9����ZQ����_^�(�.=�yg�1�$��R���Ĳ���Ȳ^,�Vii����6�qc��1����
�9�)X�e��&���Wv̅xw������z����>~҂k��q�7{���-<�,����O����<������C}l~#����]� ��)7;p��}�J�t���,�-y;}䞫x�B:��k�޷��h��z���л�\9QYܲ�,t�O�#T����q_y��mmc|��6}C2C��{·(��6�-���%~��ppǢq�x]�p���Ss���5Y�����7e�ؔW�+��L�z�Tҩ����΃S��톟#��^q�!h�{�u��Z)3N�W{aγ�����c&G��C�rk�@��4�XQ"d;�r��6�Ԣ1�Tk˜M1�ml���V�R�D�DFۉ�
�e�s&�)���pyqm����s0Qˌ�U�\��Sn�WhUX�m��v3�#�w��ی&<v.A�;r�X�B�9n�b�q���cks�.Y*���(���%�tG.!T���-Z��,D�E�R��1&���T�U̸���1����A�]\��pjW�6�5���ai�D�������LL��Mjճ�E�ZV�3"e,̹�U��s��#��*���MfD֢�s39����Y�*�J���7w�y�5�f�1]�)����rR�`�l���ZZ6��<]�ZZ�4AR��6�T��ҹJ֪*�Z̥�Ѥ�q1��-��K
#*�V�u��UD�.0^5�B�E��e���\�yl"	��X��s�nk��0^R�"�\��X��79¨:�[j���iY�wx�/��-��]�nS]�E�DԬV#k��v������H)�~o���!D�&H2�b����G\K��AG=�(��{ �g�="��y"/�~ϼ��
׎T�DȂD��M�/������|��ojc�sq�h��EM^��H"w���z{�����:M�s��Qٻtn���VwPa����#]��v��ۅݴ�ً�Z���?{��&D(Q#B7Y�&������g�46�[~z݌���ȁF������hQ
DȔAT]o&��7/"�V;�}Y�~$��w7� =�� ں�1=
�*��]�.4���ə���Kj6��~���0�$���ڙ�����.zp��͍��{3[�c{|َ�G�LD	��BP��:n�/f�����8H;9���'���d�p�t}�ila��=�n�a�|�wx��xz�ı�{:��1���Z%Q�=g;On;��l���4W��=���.�5x"}Yu뱉P����> w������6DL�&H2�b�����	õ�4�P>�6h:��>'z���c;m�I��(�M�zgՂ	�s�"T��Bp�jƳ�S��r��]mJ�H��ˆ��ꓢ"%�vʘH�H�1+�7}m�I ����A?b�裃�uo���^���lI��[dWb��Ĉ�dB� �/]A0���	S�^�;W�4Oѻ��?r�T	3��,�� ��u��%ȅ
`Ș ���x2�*��	;�ތ~���W$�f�|Ǻ+�|U3�%���)U��۱k׻'�ߚ����߮k�� �H݊ԅ ���U����xk��Y�1&!B����U�4�=y�L��w#/���+�ܾ$G��l���SƁ 9ﹰj��)'u>gn�)q-��p��Ӏ9�t�l�:�7_�ﴪ��Q0rs�ܞ����t�"ܚ?��|#;��������Κ�;E3��BY���\+],S�het�钝�ٲE�������u��=��V�c^�ՠv9�Xkyˢ�e��X�J;�����2Z.�\���.� Z�k��s5�$`6:�����sB����[��W"rs�iC�v�����;>+��g��]�]�ыZ�&��>8�����(H5�`�7lU�z�0�t���$x�7\�:-$ut�����T�m�Қm��T�;sh8�F��<�k�E�;��;b�?������t�ӻDLW��u�O��Q��?N��6f�E�Һ.���?�z�|H��2�	JB&`Ħ�/m�g���s2<����I�6�MO=�S�H�F0�M+��}1ӕ�Vr��Ĉ�dBQ��?"I������X3[�<N�N$9ﹲD�(n�D)�"`��_�u�X��=H&�o�.'�$���I��w$~5ݶ^V�8���~wR�|Oʬ��Fff&�
[�b���;���ǃ�����
{,��ٳD�C}�o�A?�����O�j{\w�v��FG��0�/�LLHD��0p|�-cv{gj�d����X�������s�mߟ߯��U��������{��^��ϟr�^�yS���UK"��{)�f�\l�P��R��ϫ��/q��y�M�AK��Q��z�k��sێ|3���<Ԙ�c���h6���֓�����v���a@�wJ���Qdߔ;
������Q�|���H续�I��߶�`��ڍ��c��4O��l��&&
`�N}�� x%񾝶�-���1���ǩ�}�L}�t������ Ȃ�$6z�=l��MWC�	>�nS������]?�'��]1}^|-DO3��Vn:r�Zui+
���������3���$�U�})fDE;lK��a�	���M�o�ȭ��ط�B��~�$BL��e�{u��n�7dM����t�ZՍtG@���vk�?߯������R���b�����0A ��L�c7���N�`?A~�O/zdʉJ" L	T�u�Dm��.�nVt�X$�C��l�Ot��tV�
�\l�\���`H0�(�c����'���^�����t�����+
����������ga�}��&��Q���4�޳n�����/����h?~>O�߷��鉍ʏ��>����I/�m�@�~9]�k�H�Ͳf`��M��w�O����h�1���r{&��=�7թ��N��ݰ	��Vc�Cہ�� �СHU��}���&N��NxF�z�C���/ݘ�������MO���òb�����}��������K�vq�۴���Υ�K�����j�k��yE�ϯ����F�s{���^���#g�B�{�/��{�4���������==�_U3�)I��R�!	o�U͒9�3'a�K�d�~>�t�$�#{�����z�fu�Ӯ��3��0�J��3S`��}B��y��0�������d���g���N=�6|�ǣ��0$R�L� �w_u7�oRɤ��ĀDV��Io3�`���D_M׹?S��u
//�+��p��	�{A������P���,ۻ)���*x������Tt�3���t�2�ߴz08k����=��׏ԃ����������ə�JB���o��w��A}�l<��>�S�z�#��~ʾ��A/{�����	�B��U�(�F�")2�l���G׆��Y�������ۧ.�l5�Q/����߽& J")�<ۡ_c�m?�'�^�[`¥�:V�Aw�4H�o������
$	L?��S�����5�:��-�WƯs��	5���`�w#�yE#K��}S��O�%&dLə�%��\�$���a�H��,�{�:|	�Wy��I��� D�ǦL)�DJ�0�m�n$|����n�$��LA�n���ut�G,	D]%b����d�.���bI)JQ2��v�d�Ful��!nym��;]��?Mo�����]4��t߳���C��DO^p�V�!��b�ya����k����w�\у�]�����n"�O����z��zaKcвH�~�|�߶���]���O���h�յ�8'��q�k�c#"{=��xT�]=��5�Ѻ�s�\G\�!�N�����X6�N���U��Y�u�<�h��-��ѵaɊ�^4�U`}���`��.�{`Vās=r���R��5m�!�\s��N�lg����V���FS˅�2n�$p���j��+Ss���5�C�ź��&e�m���Z��{NN�ޞ���6I�<�6�Eh��ٞ*r!___x����~p��l�����Nmt�;�i���i��l,���$�{-�CwK
%DIHB�"��uD�WU)̗�޿e{�I��+=��$��]4H=��#ڣ�d�Q����DH��+]y��$o��� ��H�ɘ������ˠ�$�t�;=�b$ȉ�*P���]s�x$f���|C��2A;յ@�Ev����z��tn�$���	��͘�Z���"T(�P&��[_Q"�7i����B���[��~��6�$�ޭ���]��`������ԗ��@�5��Z%��לy����r��Uoi�v��bɥŇ�o����1jq����ӕ�o�I��$�w���}>��M�O�X8�����["��r&&�L���o���%��ޓ����０��b(�Vsý�w\����(����g��r�y�q����x,�My��5Y��<<�$�(�{�e���+9�	�V�uﹿ�=w){3ET?/w���L(�%!
��}t(�A���� H9X�t��c}������ ��u&4�;)@�2bA)�W:�l�Ue�1SxϺ|I?7~��?��:U�\�������Ss\A�B(���k�`�7�o�o3G{� I�ΑD����'�=�u{��y�\�Y�\N�s�mƍU�Kgn4����|���N���\�V�p��D����� ��P&;�9�Q��y�L	3ݷC��h�W��Q��~�$�e�P&�1
 �H.7+��~>�}&w��VG���� ���s`�g�m����ݨ6c��W2<'���beH�*bT�/|߂_t��e�Q�yڪC�l!ܿ~Q,4R>h����n ��#�sk���mF��d^g�->Jr�/�I���̙� Fz�v�"�¸��������s~3���474��TL��(R!��ۊ[z�?|S�t�$�g{m����M>���+9�`�1���D����ן̒Fz��>��0՞A�>�kݞl�D�m���h�;�q������@�6bJ�~� ���&�C�����´�$N�5*]��5�����""LD��(Ow��lO�o6� @>��=2#o�ђ���=^�� 7�1#n=*R�2�L�e�`��-]�v��2A0����'����(�b� ������{�k�6�J�0R�b��� ��յ'�Ez;��DOP��pI���O��T�@��
��� ��P[���j�q�NV�6A$�^����N��8�G�>ʯ9����dk�y�ag|�����/M���<4�}pD���97�;N*�<�q)�F�e�;�w���*�T���;�����39��b&B@��<<,�<�H>}�L�}0���+��� ��mdP$|yﺙ��3����E�۾A���*D([a��6�u�\爸u5���c�۪��m�۞�֔/���6R�"DĂc����� ��m}$�#�����J���W���˶	���U�$LȈ�2�	n�k�fz}~˄���g��`{� �<��
'��a���ٞ��'K��Ԕ�j�UM�7]�=��L��1>W��ib��:�?r�آ7/�A�m��T����gݶ'P~��&���"�{_I'�{/1�@#_m��|LǬ>'O����%FD�P!)�Pi�����6v��˲�-]8��ν�`�~:�m�?G�8X��&�qѩ����������~�s�ݢyM�;9���\����hp�3ٻm���|/b����ʈx���{_��'�������hw�m�"��@��J�d���C��\}�����>���t�ǝ���{ݢ��h�$Վd� �NJ�1�霽��읣����=uw<;y_1Dn��5�|7}�;���Y��o��x1��yu��I�ˁ}�/���u�?e5v�3c�^A�7����N���{β�0I*c�Vf{7��4y�<{t������`��<�19���[tN�i���c�G{�����-���9>���rIs�+�Hs�q�h��o��^+$�q�8ي%�S��y8 ���K=N�9p�n��W�a/;���M�ȣ�r����;��[�{ee�}o��c��p���w`��܏�M��,�_m�6��w��?@:7^�F߼�xt�����Ǉ��o6���L�����$�zy���6"b�I.��ħX�F��50�
�^�m��{���y�R���o�{��ݷ��=�ϝ����iA<�x��G궋˳�;�+ήĚ��r�V%�/yoQ�g�����=�{������_d�&��m��g�F����to��yx���不C9%�o+D�S� \���#%����|
�^���&�Xǰ�<�xo��{�KB ��6<+�Jvq�[3��%�	Ҡo~���=�u�9^�X��;�vn�컔d�����d[通�<�h���k���3�^���7{�l���c@o����s[���µ�Ǒ�o)�	+���<��+�I��s,�}8���R��e�tn"&�E5*墱XԬF�`�6ʣ\ʣ"�bQ��2�4.3�e"�*�R���b0����`��E�C����j([rً��5Vm�F(ۖ��q�X�Z(�J(���&5\�1E�33K�0AƢ�k�AU���԰��UTm�Q��J�V�2�j�*�&9P���($V+�2ڣ*fS(��������m�m\�B�PD��H�0W%�UA��M��.���UQ�FV�i�P�T�*YR̴Pc���)��LU-l�֠��7
c]ª8رU�Tb֊�l�Q����h*��A�[U�eq5���Q�V��)�(�����LD�B��7���*�[q1CK����[R�Ye�E(�Z���ҍ0e���(\�Kq��ҢV�ɆZ�ĬUG��[
Z�����1�2�S2�5��r��UTR�kE�QF���L��G-[(�Q�Q���e���
����"�����T�|[�nV�M+pu����u�y���{^3[j���e*z��z��}6�u�{v��jɶ�c.x�:Su����b�b�u�9��Lv��h̙�h��l���:���]���Y����Zz�c���o��k�q�}̀��[��̎ޝۂ!^7����7k5�ֹIn�N�뇰Z���k��S�͞S�0W.�Y�䲇!X��`��Ψ-=����q���;��Z`;f��x���6C��M�۶}��ڝ��i�\���ޝn0v�;>y=�ݮt�Gk֎���oZ�/�;�d�[zL�y����$�(<n�J�X��9�y͑�9v�r�]�� �q۵%���m�K���t�Jgu�N0v�<���&3��F5�]\=Z=c��;)cs�u�ۋ�bY�r\%�{p<�9������vӟxz&�H^����9 ŵ���d�_>���9�ۭ�@��^�g���y��c6�ݝ�a��
��]���@�%Zv�b��gjwcp����ss�U�Os<m�'.@Lt�M�h��n���7&-��@��Wf��:S��v��-�n��z���#a+�[�2�vs����8@]�coݩ6#0�鷧\m��ՃdJ3���=��8 ø���MW��g���c�n��[c�.��L���j����2v�q�C�<��+�qu�hӀDp�sd�[qrUu���÷���;�7I��s�/8IN���L��V-��ɥ���,���n{p�m����OG2�z+`����\']�K�c�nӡ���d���$�Ŷ��K��|] sRwj�puv�P�y���;�؇��E��V���ć��g�I:�r:�ܷI�4E���ų]�s8݀�;um��f��j��6�;pd�⒃m������!(u��<ϣ��@���v�ay��\�9�=�����l��vҼ�X�@ݸ\ة��BӽP8��x}���#N-8�tv9�[Ivn��X"���tF�]�yÂ��Vߙs��7ϟ6��v�[�z���psClVzt�p��N7'-��8��k��9�����6S�.��nNm��5][a����%\n�И�ֻh��=����=Pq�Mӊ.���r��nc���{8�A#�q�[Qa�X�s6:���;��������Ji��ɳ��c�v�"+�+���k�N0x��Y�����T�8�����i�
�y���K�YW�\ah7��:���f�ٲZ�q��I ��*Dχ�3�J&"dL���Y���H;�ͦH$���l9�5/���/]-ڊ�}{��.x����!L�b����l�\����}����� ���`�Z���o��;LB���D̈��*P����I��?��V���fk7�H$^_��� �_m�9?B��L��P"i��]��F���A'z�Sv�n� �lW%��%on�y�Yd���6Msp|�J�0��9���Иi�F��A����7�$��m��$v9�Gñ_q�ݍ��
'�
Q���&��!j5�,�{
l�]d����>.o-Iʵ߻��"e(�Ĩ=»�͂={�A�7񯏮�T{y��F�{�m�Oă׹tޜ�R���!$6g����_.�S^�h��=��gܻ���/dL��~s� [q�%[��<Cn��nE�39�b��/ S��V�Kh�Ea>S�OɗLZ�Uڑ��{��	$��l�;Y<hf;=�7�g����>B9$(��Pgb_�`�u��o�j�z��-�������Oǯ��`�HQ���D��&dD)�	v.%��y�<A3o`�~�~�	'�Ȟ_P����uL�$޾a��i�)JTə�%�5�Q���i�ZFeۈ�2��	�=:�$��v* ���.��xO�P�Ga�����v��fLf���v9��=�/Ot���c���w�{IJL)��f�$bT�0�����]�l2H2w6��G����;��Ϗ��nn62{�(��X*d�@��%An�;͂~.������Nɭ����A��	�]w6	��v�1������������A"���Ԓ71��}���c�E�+�P�H�6lx�WNT"W&�ݙ,U�匹�q���b��[�2gew����.{͍���
+�u�ē�,�@�O��7�.4����!A�!���:�B�b� ���$��>a�H��=yJz�� �)�ETܔ&$D)�	n1�6~�ݍ�����]M!�w>$����	$}����^p���MJ��/�T��IS�F� y�v��\y8�C��σ��]�e���j����}�����DO��C��~$�k�d�y�e�}�F�_^������ǬEˍHĩa7Rw����ֽ��xo$�g��]�}DFo�6	#�v?����qs�#�4�7�
��!)�P_Om�|H$y�� �o��b�{y��	����H#�v0ޜ�ѕ32$!$S�y�p<�����Mt�I ~�A��Ч��"�-&��R�Vk���XFe��x�EV�n�s��3�ɒ���8 $���l)���d�̺'�{��)6x��-dW��G�����Uq�S��&�@��S;Y�o:���/�m`��-��w�m�	^v?� ��ntQ�"��44E=�{�*LT%""L�*�I�.ݮm��ޞ�:��2����s]�������]��=�+k ��ݯ�A�@����^(/w[�E��6DH��)B���P"[0^u	?]"|�jy&�����$�nc`�tQ ������!OtV�H�V�""d"��Q2�/�����`�lP$��р�Ũ���$v���$]�	�m��D,�!)�P[�9�X��<��깖}��&7�$�}�@�C�|�k^�{D7[�o6�e��S3"B�bC~�rܒA���|s��qGVnwv�c}�o�	;=	$>����o'���(5�"|[x�v���U�����	q�_%�,��:����c����#ݸ�����!��.nLK��Fw��>��y=ۥ��s�����Y��8�׃;�%���e綶.�lid�ݐ�h�е�m�����˃������Ų��ظM�x��`����5�xa���xl^�:x;P�u�.\>���sS]��ElcA�8.��Zr0�g<�w]^�ϓk�ĝ�<nwgCKp���.��T�Y���K;of{rgquԭ���[��n�j ��E+n5�h�f)s�M۵Ȼk����Z�����j�3gp___{�{��2$!L~��k[$��hI�_y�`�\>�1�Ѷ�p�{��!v�Q*��2����%�!�sd�m	e[������0~a!*�����|� ��~^���u0�P��bTB����,#]�~����|��|��13ؼ��{�@�]��f��DD�E#0�f�vs`��Go��{���Y��O����d�>�w����5��Z���"ol
!z��eA{;�X	�y��jn��<g�
K��@�H|��	���a�5~W~��g�6n�M�@vq���q��5��eof�VNu��;n��;qVI�__���V�هqþu$Nf=��$�����k�,)�P5_�K���}��}v	,���#"B$���U��a`�4:F�aH�u��#o2MLa��jĹ�jˣ8��c�τ�׭��(� ���sQ��P�J�Ʃv5��یN�E�ć����8~�}Oď{0�$��>�뜵�i=�y7z����en�
AJI�"[7Z�����v?�ѵzb�\к��A~���$��c��������L@�l/8n\wVC�c���B��LZ@�O��V0��:	:#����a���lsA�DDIE"�D�`�v�2@0{6|�eU�!�2&��	v�$n����0�:+�_f�����1�-�nn�,�;9�'ΣY�hm���D�[����;>يj��B�y�($$�ąU�V��mDAo7(`�����_ xi������˦	����� u��ѕ33$��W^��ܬw���W�$���2lg*�}���׶u+�� K�)i�!a��V�1k:�u�};ʃ�"����������rc�����HU�*��]W�۽N�}����4����H��,�g���3��(7���V�6t�m*��e�e|������r�3�$̑/a�U�sw;u�$�m��Lr�*$G�_<����:�w�Ao��9z"� �̙�4�5�����7������^����*����#9ʉ'��{��k���������@��Nwe�x��A���O6:z-�;��@'Yp���{������������k����`L�z|���M?	��#�G�=���'���TL��	ό%&Ks��l��w��s0�7�ו��N�j�h��U�GP�U�v�T�16꟬{
L�ȑHl��_?����B�Y����w�enc2t��=�2�JY�$dHB�r����d��ls}H�Iu���~_vo��Q��`�����OH�ӯ=��(�z	\s�}R΀V��_���׽ߨ�p_j>�[����hSu��ڮ�3�*j�`��^��d_$����b�2�*`̑-���I�݌<��=5~�n�h����	>��>�����;�7�Î%�`%�)�f,� �p�׻c�Q����dz�^Z�??��O�c�1'��c��[��#��ݭ�P�K���^�Sgw9�H$_W��H�T/�""J%1W���d*&w�=�Q�9���'�O>�0A�#�����������X*Q��&L�������y�� ��w���)�*�.f�ĝ��	����a����aI��&��}�|x�������Fy�$�u��n�x,�!�;`﮹�*,���FD� I�;Z����;�o�N�����6	�{�A�Dn� �O5�c���jJsq'z�k���[��[��m��:��c�dWF/p�Z����+fw����w�����~�3��埧m�-�gmr,��UES}E�g���ZB2t�����n�������Nûs�K���C4/��:�m#��9uڋ��7G;�Cy���n�;��eM�u�`*�z���V�arb�\뇹���!��"��=%��5y �g��G8�FՓ�֗p��P[n����Ƚ�MDq�@��O]���>�ݺ���ݥ켛r�rW$Y� k\�u���O=�C������"Ө`1���݈��˝ĹCts&�&������:d���G���A&�n0� ���x��f��=�^m�I'�ݍč^VRFLɘ�L���D�f�8�zZ�.yt8�v���'�Ln�$3��}g۹^^��ݟ�o
!A��BaLS�v�d��4I�yW1E�nj���ݍ��?F��L�l(ϊQ&Kf>�~Y���ʮ� �t�	�Ϸ����L:::cr����I�����̉ ċ���$�s�L��]̬���VI!k�lH���D>�l��\p��p�o��|���eH��A8�����Ցۚq�R�Ʒc('jI6�]�֗)��7����}��D�~��I'�7�ٚ�^$����#���H�d�J��ƈ��S'�lDm�`�,�ot��r=�vn^/��ͻ����|Sȶ���"���W��/g��TX^�\u�d�>�3r�O��9��P{����	���Hs���?�X�td�e�S ��-`̙�-��_"I���<����w��}�8h�K�o6�f���)H$����s��r6|5Un
��F$���s��ܾ�3�)�u�G�:�k�k����Jɒ�s�Y�$�z�q���z�_� �gMK��l	=}��ϳ�w���fai0P�
c�j�}��0����+��������8}�n�r,D�`�Fb&d@�$w|G�]
$mfm���2��(�����U�4H�w��C�)a�!a��g<5W��k����w	�vD����w]���g�`�a_�zl+��M��b��Q*b�-��7�2�}L�v�,t���0�i{+�v�vE�ED��T*b�	63�3���_��0���|8�,7��S�I��I��>�9���c�#�v�NC{����=U��N�`����J�:��ey��a�o����o��k��V缾�wZ�q�0��2s[�e�Vh������~������mRr��J6yzٱ^���}�{����B�^P����f��p�=��K�ӽ(�����+)�6d�U;{w�����Vrvl�ٖ����̤��~����[�x��}o{I�JL�S/�x�Tv	�p�&p����7�d���{�&!����S��)�ҩ<^$t{�tQ��#�"�O\c=��z.��]Y���x���w��J`�sݎ��z�&^]�0����/��g�}f)���#��gGb�}��r�����}*e>�
�t��7ڮlY���~�O��
��Kf�vI�)�������"Y}�k��{�=^h�/�7K��'��9E�-�;�������*�:��|�����[�d�f�M�#I)�g�M�v�f����H��t��y�w�^��>KM���ތ�8w�����w�ib�7*ٗ��}�:�����蔎Α�ɕ�}���{� ��O{|X��f��u�V�v�a�=��_{���R|Y��������3�;�?R���˙o#�&�?:p-�9<�.��I��9���,97=}7��vbJN���nGK+<�l����=�'�˄�U���V<`R*���^O���AC?xA�QZ�|¼�J���t뗟�~�A��j�ϴ�s3f�X�Z5E��&��ܳ1�LJ"��D\pp��k�.2�(ъ3)����p�l�V�-h�Vۉq+lkJ�B�5r"ָآ"�<h�.E\n�(��S.6b�+�L�X��3-b6�Z2��
�m���PT�Ԛ�h��`��b�f�"U�T��D1�r�(�3b�Tl6�Y�*��+F8�1�֣ZV��-+iMu�i��c�kr�����j�Z6Z+h--Cw2�,�X��eqԣ�1�L+5�m��)w�2�R��ʅ����%���U�+
��X���TE�#m+c�S5���4r�
�"+�q��h�,�Uh�1�iQX�QZ���1W���q1��eDƋ[�ш��q�(��6ʨ��\ITTE*UQm��[�PYR������EEb�፶��X���Z+�Mʡ��QjD���$Ѩ�%EF.&3\�h����\���Z��X-�6˭���6�
,�,b��t����b̼�ݜ��Xw�o6H�_{|ى��>���0�ۮ>�t���+����	�K�m��$��]>D{���u�'��W6OPo�
0� P��>��0A����}jfC�X'��������2Nmt�>�>���&�	�3�R�H�P��fP]٠5�A{X���>E�n)���qR��~�~��	���,b`x�[;��Asm�'�3k��>�	eF��c=�C�խ�w�l3���ҘP�L	�bF��<A�-M�����ve�A~�[`�~$��M|	���Y�B�������&`���0	 ��u
$O�h��3�	��Ź�h�Mg����]4	
��&J%)�?Kkn��r'ԢXg�]��I �WM A��q���j��.�wӅzQ��-�U\.�F���E�N.����#��ku��h��+{�]ė�r�}���(T�-�ۨW�G���v5�0�����|3*`)�u��O��f�0}��[�\��2�}]4H�]���;��|�o����s=;eǫsl�qɫNʇ:�����>us�|�fh��0��w��S���>�\���J�|^u��=��D�+w���/����E���7A�H;ճ_9�(�""J��[����Fz=���8�{k�� ���o�IT��TW���噾��1�Ԩ
"b$�Q!��y�I�׽�L��3>�OtKk�]��'�F,�� �}��$DjHaЌ	@�2��3#�,F0.�6��?��	��k`�Lww��<Gu�����|L�+	�J`��v�������H��Q�"�d���I"�;�`���H�Z
�j���/�D<���bC#�mɆ݈ʜ�~�I�~�Ԇ��H�ǣ۲""'w��y��O�N���6�
3(����.N�Ůr��6��ާH���z��|�{f���(�=��kr�q���\�%c[����p�vш�\M؝�y�����h���x�6,9:]mzu�5��ϙ,�I��O 瞕C\�.N�]`�8y��sA�6�Wk+`���@zp�lB<�ٱGmn��q��v;#�m�h�&[m�/c���O3�Gf��g��b��fY�}h"1)����'m�ƹ҆K7a@:�mv�>u���jg�����DLĩAO�p�~��&�wi�H$���6�_�u���F��c�P$��S��r.��B2�TÀ�^��P׮��xgF�7���H��c`I������.�5�'����們�B
<DIS��{��	���d�}��,�N�k�hx%﹆I�����7Z�DJ��*$7�\럔d5�;gl�a�����o��##y���ZZ_ta���6O��x#B�D��Mcd���*n(����&�hhF���`������|y�b�z�*����7d�ߜ'�M�����c�H�v��vv���϶�d��)��nM���MD�O:Z�P((��wQ/�ӈGӻ�d��B�����2����`����͑	��l""bT������^�J�}��#�dҿW���qU�I0.�A�=|k
͇A�����}��l�Q��-���D��M��
`g��b~��L�G��R�����	��~��y�	&27�Ue�$��f�R����c!���0�/���d�]�� ��v쒳��0���H���`�H���qO}���Jf�)���[8YU�*�nWz�	.굄�$�^�D�L��o��Ǥ<��W� �>�� z��J$�ȅ6�:$��SE�����=��Oā��$	��6}=�U����n������w��tp�m�w4IwnK[;l8�07)��d0m�Wa��c�Z;��}���f4qȚ��?��T	J��͟A�} �uǯ³����23U&5+��@�F~��ۮl�z��>��H1���q�G��g*$��s`U��8��Vc��t� �&�"&%J
[9_P���ݯ�/{��Ѫ����M��ռ��Ƒ΍���z.Ɉ����nj�F`�G9��Ѿ���)䇯�|/��y�_��h��.E��2�E�^�^	]��I�܅V���E�lp�"������w\�dz�J�ì;�4I9o1�O�����9)Wͻ��_��ƀ$��Q��@��
`6�n?�=y�É�(k�9���LߧƁ$�[�a�O_u���I���ֽ�Ne�7��R�c�Sx�j���[j��<�^.��k��*>����oϮ���J�ȕ;�=�Ay���~'o�� ���w3���G�K��!�"��R!0�=^2>5�q��HR�{��	�{��H����`��`X�w�ݽ��v�3��P(ȟ��sZ�$�#}��1�J�eg��Zg|��� ������A%_u���$���?DĩAKf2�.�yp �[����^e�$���qk��wh<�m7c����x�{'.J�s�L�[����
g�{݇�j~����^�x{Z��rMʶt�ȃ�whV@wu�j0�'=�m�1O��">���/���$G�6��~�Nc��=}�����I �����D{g��D�p}�l����1 ȈR!0az�t;���ٗ�����T=���ݒ�2!_��߾���+艔fu_n6 v�|���D{g� jd�j��U�����ě��Sc�
*$�ȅ2a���@@pO�o��v�nU{�I$_��Q?E��A#��E��񨛎Z��C�^PF�0�D�0�Me
$�c��	f.�=�=ْ��Ќ���{2��"�yS	T�J��%������cV��]���:��P'���>�O��[��I���Fg�c��?L��!K\i� �vޱ�oޟy��u�8��v�}�K��~=�����](�.��4zŰ�4D�|�U]�V�#Ok)�����A�c������j/y˾��ḣ�Ӂ=����5���6u��s����._7�pqsn��n��PŎ�xۘx^Q&�tؽ�ӻ^T�����"�m5�pt8.S�Udg��������xnY�0O��{\�.{x�X1���1GMx��l�;x��x]�t�����c����7��x�c�[B�5�}�]��n�
�4l쬙:��F�۷5�|��l�@rq�lnv�iw�^x����r��V�Vz�]1��:��v��Gc�睇v��c��B�AL�=v�, Lsȍ�������(!LW�ξ�	3yh~'w�͂��{�N�b��.��S��H�s���3�Dd"bb`�lOn�g:`S����՞� ���I����0\V���R3�w�Q�
���f$�2[���@��{/�0I{v �r�h�s�I��D��_S��A �R!0�=U�����S@�O�}|�$�ވ�޷���	��=~�4L�$��PHȟ����H>��
{�*t����F���Xdow����Yח]"<��rޮ	��:���vC�d����t���خݵ:N�w36�s��������u.���~�|�S�״�?ww����
�^eO���s�4	�������A�
PA�d�0�/���1���w+��B�;��Ү�:����W�mʛ������W�a����m�r���ύ٥�c�)ْ5�^��W�ڧ�v/=D���1>ɻ�i�V���p ~�^S�{���hz���8�ė�x�,FL!&aJ��s���ĂA��U��a�=��7�;?���|�$��wz��9��K�D̘�-�r���T@�QW���~�i�A��@�H����"w��}�ì�C���$�A �2"	�a��Ml� ����z��6�l�e���3���@!w�+��}������k_k����]s��yӉ�V9���t��q	�kj7Ku�K��>������@�DwMֶA>��Q��H���9<��̟���������zk蟎�'B"$��-�����ֻ,r"�ǫ���O�=��I����Ko|p�u��?ka�D��$�Fa��}D���$}�{�=w�D�},3^+U�3��GE�ܖn��*z�t����{�΢o<V�.ӂP�YO�0^v�/:� ��@�/4��z���ߧ����Я���(��`�Bb��*B.�l�8v�&�� �ĐUS�$�H��ȯ�'�|�{]Ǌ�|_K�/a��1[�ٗ�$�A���ʳ��'�Ztlnh'�ڢ@&^EA#/_6kw;rkG�����'k�[��\�������Qlڧ')x�ܨ��i��ۆ#6�!�������;��~U�(�`��	$��}L�9����=�{ْ(
�"��\��&J*�"��͑uw�j}Q��w�=��D���ّ_A;u��ě�
��)� ��{��(�����Q&fP��+��$O��i���v3i�1U9�o4�D+܁@���� ���0B��)���u�������;��������r��~�HD�t�:����Fa��~���o7���yA׊YP/.����
�O�ȍ�A,SX+��HW�%~�~M�.� ��;'�K�������E|HY���Id��w��C�rq��Duu��џr�dP$=�u�OĞ���y*���!��HQn�a�4�k���:tm�nus��.��>��b�"'0�H1(�I���u�I��<�����۷k���v�/�ӄ�̀���l�؂2�@�0������[I.���V$H�}��I��P��X�YJ�a~}1d�1�/�d��HBٛ��$�wz�O��|�#�.<nu�Ǿ$���;����Oǅ�H#fe�����n��$�{Ι?{��@���h_u�3��}o+̓\�^�"$�2Q3�y���L�*����Y����yCo��$|}��+���#������O�W�''�E%\}��U�_k�t��E(�|>����\]��ΉDf�Gf���d�pԄfJC4U��f�Y���WN����¬¬�+2��U�J�J�T��+:k�+5J̥f�Y�Y�Ve+0�4���u�Ӣ᤬�Vi�B�ih�C�%fR��QYӂWJΛ��IY��Ĭ�VbVj+1+2������çE\1+1+1+5J�Ef���QY�Y�Y��Y���"3.�	���k;o�"��jJ�l�U5������|����zn����o��8��~?/���g�����WOӧG������|�[����+�}��_����RU�񔤫���iz%��>m?S���}��_��s�}c��5���q�|/��=��zw��J*��!jP�-(FKD#*��������hJ���f��}��Q�ԥlSb��K�9^�=�����c�|&{��0��{owWcó�j�}.������yN�=��szk�z�ו��yu%%^j�J�����y;9p%%^�w�))*�Yqz�'��;.�qy8���}=��4��\�n���QIW������O�����c�����'����'N�-꿊���_e�qQIW�����|����]-�������|ޟ��|���]����v<�mw�&���8�2���<痕訤��u�8�^{��E%\o��o7��������
�2�����x�� ���9�>�#� !JP �(U ��(B�   (O���PP � �@�(   @)@4h�R�Q� hH��)E$%@�AT�(�R�����  jT��EP	 �J $D�(P� ��                                      (        ��[����e�T�b��YhK �-�R��EU���mͪQ *�wdErp�
�@
 P;��5S�9hUD` Y��"L����.��ĭ几 xx �J�0�YB��iT�4�ЕS�7�("RA^�zT��       P  �.�#�f( �jT�3E.`2)ޙ�y�TPC ��@b�P��yb�4�s4(U�)͇�h : ���Α Y�����@Q�Ȓ��9��АdT�� p��t{��,�Bu��ol\ �6Sك�!^��]a�AD (����  �      ��U�U@�۪�W�!��*��� �	�eL��+&"��F��7 �Ъ媥)��p��U�   8��s��k� �R�s�fX�;sVY%���Q��ī���r�նܵr5�{�����[��ڦ������@��  �        z��M��Lkkr:.5{tVf�n��� 8�l���J�=���2�g!��Ͷ��m��k� �ڔ�!��677v�(֍
<  �I��vU�\��Ip 79��r�3k��\6�nwv6֦��v��8 ݫm��#�՛��71�#s��R��@��
� )H   (     w�a�\�s-�g�4sj�l���ƨF� svY��V�nZ�kM�4,�`G ��\\�U��J�D*�<�@���0�]�9��Z�� �4%rӓ(\�T ��6�vU(9� a��m��\Xۖ�i� < �?�� �O�bJJ�S S��  =��F�U=P  T�����T�@h2d0�IMJR%bg	�LD�Q� 8	=f�z�L��M�=}� �$��N��H@�l@$$?�	!I��$��	'��$ I@�HHs������s7���f.��3^s�+��:��َ�YP'Gkl��Y)X�˽F�wy��6H���!����ᖨ���r�e�1�q�Xp��z��W�f�-wwqж�h!�C��2nѻ�f:��[��^+�������mG� e�r�w.5��n`-:��65�vs%�� 6^��9�m]�ԗl�v�ũ;&�/bV��ڎ��-^�n���]�	�(��f�N�t7DIr�˗/l���`roҀ�yW�A�mk����N�& .��2����	�gC��+붫
ɍm���Xw+1'#B&`��ԕO�4���x0��i�79��:�JWq�YF�8�n�{Kw3M��bǮ��wlͻڑ�n����F��24�୘�[4���u��y�e�0��w�j��w���uf��˘%�4S�i���ւ$yP����P�u'!wyT�S���y(iͨ^�Y��T�S�ͬq؏l�]l3�ڐK�"���m���	��BLPz��V�f�Tn��ٯe��*��P�sd����a�j��1غ�Qǻ��3O���;Z�Vf^9�X�4�Y�T��u�	��H�so]�b �ސ���n�^�ñ�bŦY7Jֻ�Cч4�)�M%^�[u�v�
�@���kV���Z�qL��"b������-a2�PZ1mK�͛ݘ$��,�4ejb'R��Ze(�ʻYW���VX
�i�j����+*�ޥDL����d��*��B�ĥ:ѻv��l ��,L�Qp�8�b�˦4��6|��mMX�'p;\.��KH(�Ӧ��ÖpGg+`�n�`g1R-�ڶ�3k���B)�y��cY'�29/ ����DA%�d���FV�uB�C-ӄ]Mz�t�X�F�"�V�Gf�A�m3ZO)�ܛ�pj��ɛB��X��wW�CWS^n�ˈ4�*�Lcb̹�sRd�ҙi��Y��(=ݖ���.�{h�-��V�0f,���Wf��Z�9Dc�]Rش����,�i�ZR�VhC��q�]p�=�Z��(bF�nXX�K"�{0d�Q���ucx)aT ��G���"
�+�4�(ܫ�cQ0a�T�l�`�fR����M!�ۃ���X��Cɲ���[�m�TX��Y�Q�i���Z׸���m���F�J����v��l�5�wAk�6��+�)�1Y�b�����K3E<A�ڊ9rj��J�y��+�M0�x�^Iʸ�EJ0��.��)oDW&nT�	-=��a�a36��4p��[;5RwhbC*���5�@d�$�ṷ�z��=�f�N�)&�W`�J��{�-��2�u]�+,M
�m<��%z�/@Gi�z���i�&R�V�����k	��,=.Ͳ4d�n�����7��.a�@Z�ɬ�d]���-��uȳ"j��P�4��[͗�������Fdd!2��t�H":ܖ���zUʛ{�����n&��R�-;;�)��#k��7m����퓰�e-_�-ɸB�Y�[�d��a��"7rܒk�CyN]���U�,IM�!�û�CWWQS�Q+w��'J�WZC��bScv&���r�]�K�p<�wA%����4b%ȃ�M�
�n��F��J��ɷlR��J� �Z���yb¦�[)�Z�hE7Y&�t:R��lf�X�ELʻ�T8^�n�~��ʁ�E���Îe%�lb�*lwK[�ӽ4չ������'yxƷ��aР�M�Zh��ue��i7ĵ�^�v�uXù(3�\��1��RE�A�֬h��W�8r�5e�H2���ݫ�7 �bb�Lt59�e̊�C��n�/uȰ2j[7.����ͣĭ6P���bݭ�Ø�Ef�$�WdR��+E�jk8m�d*䕅%V#RT���3te�EjE�^�N�4n�c��X�]�2���Y͘�J0�ުu2�������":��
��i�#�)�3%�wQA)����J^�i�d�`��TEO�U��pD4c�	Yt �������Y��&�P�J���8�k�m�ˣ,��p]K�C�^V�����ؕ�7)�r;�u��P]��9S�gn��̸D�~I7������ûj�U�u�BjN�
͏z,�4B��������Wm橣�͇kRR�b߀���n�&ʆ��^�*�&:/+2aʶò�e�TJ{-e"j�)pK�Ȏ�²���P��u�o)SJ�"e�/H٩KYL�2+����˃)
ɷ�%��6����n�,e^�h3W�FhP���Rt�9�+���;k2�5o4
�&Q�Kr���q��ܔlb���Z�Vnm��m�QǊ\�(�`u�Q+^\�|��<��H��g%�w�M�V�xQ����%R��8P�#:�M[b�6�\r�陕����Fc���7b�l
R�BpYgt��(��̧����EG�n�;�Pc#&[Tڕ`�h��������t-Yt�ȴ���%Sb9��ՠ]̸��FCiVnb*)j�xi͖����Ĝܽx	j�B�/#�7Ot,{5Nj@��������<:�M��+�D�u�YOn�`\sSֵ��,��B�Y*�8"w'�p�J�K�4��feJ�S�63r��M#�VA��Ǯ��7H�P�+�Z4[+NY6��^�=7mJקe�n�*�ˬ����lL�Y{1h�F;�mR��0�v�T�m�O]*n�H��̕+4dscE�D��\u&�w�n9D v�����D�i�lk���ٴ�;��Q��&�&u�����$]sە���� Md ��1m�iڔ�ɻ���T4��5����d���:6�����f�6�RF��6[e˦�4oka+C��NR8̕ll�nU��h[e=�uz���+m�Cn����J3�廻ƭD&,Rμ��,C
���DG1�p�:&�T��\˹�Y�j蜹R�mF#�`F�1�QF��Ֆi�
�9���f��
rY��.�,����Cͽt/ )�Ғ�Y�.�d�W1(�jċ�
˘��F�f�CDU�\�Oi�n�����ʗ	\�Stj��u���!x��x�l��\���<.��QI]��*��1Gb�i�6�SV�����H�� ���)�ݼʽY�-�*)u.!�RZ�R͗	��w0��+XI�k���2�p�Z��6ج����8 Ҳn�V�gj�D7-K�<�Lek+�,�t�6�y��H�jW��n
�Y�ɈU�qar�[��6��Ȑ(�����n'y+@i�oح(�ɣ\Ң5��3�v;�͌6�!���Y�Ť��xXA��9N�'�hM�gbBG�yۏ���X���{��n�5wZ1T��R�+������3A��-Z�ϼM&b�<
c�\Fz��ݨ7�+TU6�Z�4o.��ЗA�z4��r�eU*�~ب*����Y�rnT��Ph����4,չxS�BR�%m�#�(��)�t�HQ�V���<�F&~u��w���Ő�|*%H�[��*M{xIt2��"�Ǯ7{����McTtf�L,dۥ��KF��s'@V��xb],��!��n16Q��
��-.A#Z(�*�+�Srٲ�KY�VnȬnS.}�]'��0fe���H�z�ui�2�ɤhc�w$�ݡz�Ĭ)�@.ʖ]�{gb�e�*/�]= �v0V�+o*�2=���hH@���]کu.�V�p�-��Br#f,�n�ֺ���<t1�a�tA�G�4-:F� /3�+*ȅ��M����T���*j�B�&۬d޹$4�m���on�7n���k��YL��5�K�hChn�<
�oo�3q}��x�۳Z�sn����G�` E�XӚ`x��1���2����!7h�N��[�14`�ST���^ZdlK6�y��o0V�h͒�� Me\�vu���\�o]�]�ߙYZ�_����R
P���Aͫi�a���bEU���ɷ�ɓB�[φ8���*����Z��>�a&��Fc�Vַ���J��+MS�4�� AZ�؁���Tue\�c~;���*�n�P���]X2ͪ���,� Ԟ.RI˳.����լں�ѲFi���ׂ�^��-Ei����L�E=���ͼ���?�jm��vm&멸�ӑ�4�ȤXv�\�/%UɀJ.� �8�ͭ�V�e���{2ܽ('pd�;!ߵѢ�V/U����V�e	��+�7oY���e*���Z�Z��WWX7v�+u�t����\ɦenb.�tSzU3[��"m!^o���Y����aD��1��4�v0�X�3�:�kuh��e���R(��t��J�P`�b�t����e�F��]`��f�V�����Sne�{m�Uk���n��h\�&P+hl���Q@Gh�
52�����b�4��Y���Hnml%@�[�3td��hRne�0S�t��%A�j%P��������}�Z-��4��-�������4M!�VGŰ.�M�D��u�)��\��r�l�եd�֖��U�h�Y���!\�P���j[�+`��/e��j�ٕ��H����f5o,�7V)��P�6�ћy/!��c&��]U/�Y��8S ���-땖��u;O
nm�mdF�R���JjVcuuU)�a�f�'y�f�m-���iI>�0jZ�Vl���z� �n�a��;1�elZ�;ɚk)��wB�ld�N;�-��f*�����r��`+۴\�v�l;v.��P)�%�B�rfn�*mn\{Eݹ���<�"t��]w@Ul@)�Db�@��M���n�Y�^_�5�8S;��$�1�5��iq�h[Ǎ��W��S@���.3F �쭬�4�jc�j�	��T�B��uUIovĽpeV
�I���ʣ��o¬]������n�zj[�av
�&U��@�o����XR����F+ٕ�݄��LP�Z+(
��v�T�#i�u-�<ݪ��U]�J^I�N�73H��9	I�f�n�r�}�}�>��J@�
y���x�T2f��u��� 2�kn�u^ԘA
�ef�[��6IX�G,PyF�w&�ק-c˔�RYtw�ô��z�J=�*�:$��@���uovbe�	u6��i�սi\$,G@���ܬ�S�M��e�Z���iqH��Q�j�DR���ջv�@�Y�R��&�v��.8����DnS�d-�� ӄ�YorV�R�)O.��{V�)o*kSp;����[�(�Bm���ѳ6�N���zn�.�6��kF����H]�N�̭���@˭Y{�V�
10l`ꩮf�`�@3��œ^��H'�m�p�ݙib�dx���w$��ךs,���pP�-ـd���y�WCov�Ũ�	/1ɓj֖h�����H�E��Z5Mӑ���x��{�s~��+�Ϟ�RD�n�V�)<:�r�Kjm�V�W�f�@����2ݐ��4ǚ�֑1<u(�3�5����(6��ր���؆:�&<@X�spމ@�V���C����$L����Q�%�v�D� zv��*�7 �M��İ�Q^��1��䷙7$�X�j�V�E2!S����i5`lڒ�4'Aɩ�sm��؅����j-�D��b�Ls5#������N�T"�L߈p�Tɽ�b5�(��q�ӵ�[ۈ���Թ�emVڎ<U��%]�Xna�,QVZ�T�UJgqǡ�QȨ�9��Pӹ�=�s�T�R�[�+&H����F��S�Ǭ	���yj�׷QC+
�w񤃸�^�pҹ���Z�^6�Hf�+Nz�K9�e�-L��f���]�W���^h�%՘���]j���x�s�g>��6����|�i᭖3#��&�7w����ۛXBH,w6�٪�*�M�:7�5��������M�lۍ�Wd`ۺc�4��b�
�Q�uLe"�0\{t���Ui�Y�+�0�b�[��MkMF�hI��xډ#�B\.n�ۉѶhPt굩b�]���X�-l+���7kN$m�[�#0��c�&�(l�Vb�&&c�P��`�2�`��N�7{.�	M�n�U�yP1y7�7d5e��X���B�����*J	uv�z7$T�gׅŷR�����w�D�N��<gM���z[.ѷX�
�ŌX���M�[{zhC�-w���u�!n�eɵ�K՗M�Qh݄f޺Y��$��|�w�cڋG����ۃ0M��ͺ��- ��"ǣLb�,���K���JN�Im�u��ʫɻ�@�#v�A�q�=�`wu*��h�j
7e�F��m��u��q�4���3v�Z/�k%K�-d�`��r�8J�M�7LfX�/(@�)	r���z7L�����AnGN�S�­��XRh���j%��
aٖ֞,������L�fhw�v|���6�l�R}���[�Ռ:3�"U�R���̂S:#6�0���B#X.��VJ�w�q�T�n�#c��I�O �5��U�f��J�К�a8��nk[b���\�Mi��nҼ#n�c��馝`I[3A������V��Ŗ�&"mS�C]Gtr����Ә	 �y2���I�S[:�ؕN��p%t2嫬T��L��"z��;����*�Vr�r��R�D��w����[+k��j�6ܽ�qf��9@lQŚ�8wS[�0�5Ԣb%Uϲ��ܭ"qR-dr�[��ݩ��(�Y@�"����6qXa��1�ʌe��f�Sڛ�#ТgM�u(���ߏ��)�J��*�*C*S%޽�R����l�H-Ú5�0�'QJw*n]т-�d[f�sMMҤ�e����۷Z(�[5�I��h�0ݔ�.sj2l�[Թ�w^v�7�3ζ���� O�2H���E$�����B�BI!R!$�I	�@
�R�,�����H,	B
HH(J�R@
� X� �HBT	
�Y BV�I , ,�	
�BB�%a@@XBA@��IP$"�� 
��$��B$� B	�� ��VBI"� E�$� �$$�H�"�!��`@Y,$"�$�%`IX!!�B�V ��!  �HH�	��"�Y$"�@H@��P!H(H$��T$�AI+$	RPT�
�H� �E�H[d��*�P�$� ��� �$�s�?����w����{�|K��[��
�ܐ�r!T�˰�@����*
�j���a��i�Bg4z�����V���m�R�;*^s��T���kwkm�I�x�Q	M��.�]�^}�f>�����W:������y�M��1�m�<�Y5jt�"��b=W@��N��c�&�WJ�90�G�$��T'Uq��'�uW�'V��n�N�u���I}Ԉ�.���ٯ��X�{X6Q�r�7,�v���]�_�V��i�OVLy��w�.�1�� m�����n��E"2Q;��®}j�k, �ƻ)d��^�ogi��2�􏵺�MR�n��7�6�IO��BU�-�{Igה��F^����%���-<I¥�:&tm��b�wu���:�[�)=V,om�;�4��q<��]ϩ��$si;�#�Vs*\�/v9G;���pлZ��4��α��y�w\��N'�:#usnF�u�9ͺ�ػF�Χ�x�>�t�N��0u��t��i,�Fn;Nr=��1���aN�*G�w����;Y�m��d>&Y�r^��N�b��s3C졼�E�Uf�fc��K&GD�>��������R�d������m�U�u<�/\,��f<�W%�oX��$��DWVU�ƭ�]_;3G:��� �/�%�m�у����#�;G��g��Ô]Dv��ʝ:'v�U�w���i�)2��,�7�S�LZ�+'V����u�Y�/.�H�ĲѦۼV���'�_r��wg�o(�=y��N�U�/6e��Z�)ͩs�>ޫA!]�-��"�	�i�k�8���	�r�'cۙ�+3P��(�;dul.6^�# Y���;�;B�P�;�ӎ�/{(��x#�b �4�n\����a]5��<�e�A��ξ��ҒU�=8����>�boC�/Up���=�:�+v�]����sF.'�U:J�t��!��%��q�9�0�RŃj\Ѥbv�]l.�Qם�e���Ф�R���+�bU��3]uu�U�LҺ�U�,��վ�8�,u �}٤�H�"����&6���5���B̀Y����9gOlØwtGl�6#>/�������:s�y�/�X�w�k���`�,o�JSi��qW�i]�3��$5ǎM�p��g��"�������x��3*�٨�Eu�����Xc����Vr	u>	L櫃짱h,ν���q�
%�=Du5|��{Q�K��q4�c��I��gh�Wc/%��Ky�3Sn�̊ф�����351�{�+8�����:�ދ�;��ܝ��F�n�X�u�f�,en�}��f@�VǫR��ea� ��j�� v:����V�;)��)=�W]��)�]�����SU��e"wt�2��k)�FU���n�q-�Q�J����s����5�0l�z$��T�V��<m����#�4���Z݅Bފ�:�C2�x��%��.a���F��w[�ݏ�٫N�:��$���ʪ���ۮ摻�M�O�#q�����-G)�>���-����tS���:��jU�n#DQк�0�}R�U�u�Y���9�L5jT���9�C��CQ⾖�"`	��j%v^��WP��;-_
}���66����. �Q�u3Qgu#�1̗B�����q�B�^_@����>�V���ej	����/mOmϺMӽ�֒]J����4];��������W$gt�d���n�'@:o
dn]�2�4�4l�r=������>�F�j#®a�plޔ���\�u��9�����*�5�����E�hvU��!2�;3�U��K�D��w���r��L�N'X�����:┥��&;��2����.Ħ�`Mε�Vg^α5��-M�a��XzV.4֦C�8#�+I4,����/����ӷ�:�KspR����I���Hs�כ:(����ΰ��d�;�{m.�����G��Wq.ͫ��8���©^��Ru���C̜'_*�ov�Ɣ�!t�-)bЪ�W��V��"$!�q:���gfޛ������xi�.ރ���l�:��9c��:nH��P�f�ޱ8��z��['���l��3��IH�쐻ƍ� �l�m�4��Ek�I`�}6��ZT-]���m�v1P]p����]��<�ѐ�I�7�VDY�H�"��mR{-�rw.��VN��5��#���Mi��m��u��k�\�Q;f���9WC��Ev49�O�%Lڮ��Ӣ�q�r|����^	%�DӮ�+W,�a�@z�=��-�̋//�+�j�8�uԵ�pQ�"a<C �:=�:[v���N�q�T�1N��]��9;��� �X^����o��dz�3u Ĵ�X1EA�(�@
���;Y���gG+3�)���3rG��;��y��ͤ��kG;�O)����I6��u!��;�2T&�Th
�Zp]�|i�zُc�w��w�I�e4t�P!U�1�zB��9:� �����9��t�ϳ��7 �層�z�^���W/3n�q�Ƽ
���9�>H�t�v��N�S�,���GV��9��\��n���4B���ӵ�2�3�g}�e$t��l]��|U�jo�2P�����,�g�N����5��8n����vdwj���i�yB�fՑC�K���:C�}3�d7������T�S�qȑ��m�������m�i���&��V�>:Ut�`��:�����=�˨r�%l���]��z$|�t�yDٜ+���s�ڻ"�1Ӭ�_C��TŐ,��q�w�^iզ�P�`=s�Ú�ꐪ��#	��kLwo�}�LB,"+u�f��u:���Жd�&�'K��I�����n�t
���iw�8�R�Q�6x��*��aQ�W*�y��X`�=�k!p��|�'b��\�SܷE۷�k�7i��Z�m�\/x�m�y]h0���%b�%�8n3�c2�Y5�#�N���4�tg'�����kqZ�Av������8���J�LxI9��x�-�y���r��X<��{Ysu-c,���#G,Ϻ��Ieҫ���K"�Y�j7P�Zi nv����u:�״�AQ���U�����|���f�Q;����U]��Y*A�#����	7^�UrM��ξ�h�w�ȗ�.��� ̶���;����va�Y�ن���qWN�2u33)s��J��n�SM�E1�듫����ю�t�O��Z�墛X7���N��A3�[5U��Y���B��'f����;GZ�Vya%Jԥ�E�3+n�����k3��Mya<�Sy��;�9�PWR���#�.�q�5�<����el���� hM���zU�v�8(�ɺM]��X�w'b�9ۙQ���Y�s'=�	��PO5u�7n�'&3v��:�rAu��Og.���:�1Q���yW�B�],�RaYjn�u� �&f��j��\� �����������N|��c+	#ne U��r���z����\��tn< ���%`��dν������)Mޣ5$��ٚ)�!X���^�Yx[�;6d�wrgm�#VH�k��ݡx���9�����%�ӮZ��Vи{�͋�#'�XtM��(��:!m%���sn��⻴w	�月l��w�T=ҧX׊r�|F�PDE_1���F�����h�gf��]ZAP���-�PǙ���e!�񪾟U8P��j�<�nUZ˼+�1U��b�lU��b���%ݙ���Z/Ix��M�++WZ�e1K�Zu��h������HT9S���fv�A����F�۴re�ps��a�{*������e������8@G��2���]�N�(����H\�++EG��Ƶ���*p<�g!��u���.
���f��{.���y&vi9�҃��r��:��Q�]]<	f��	���0NCN`}V[�f쥢�w�*��U�u\��D��5�+��׷�淽��%�f=��k�.����8*�*�w�g�u+�]m˽G���^��N�uB�&���;-=B.:�zj�gW׺��60K��bDp|�B�iu*i���٩�Ƴ������WFcT�ǼֱR\�ҩ.��[��m��8
�%��km]tߕ����*p�����㱛}s����fm[������ͬ���]��M���1b�.zv�S9�6�B�+ŭgv*�(5]YqՃ� �eo+ŕ�Q]����bKWp�{2��Vv�yx��=��]t��8��f�ӱ���.]밻/'<��&�@��;���-�t�v��KՋr��(�Wi���I\�wG{ce�}*4��ڒ��(�A�"���Qi���vv���\Z�v�2���$޳U0к�71��( h]Z�����T�u��՛Y���:`h��v��olu(o�7e��,�y;��_J���d���7ٴ���&��Ǖ� �-ff\���<7�mp@���^BvV��#y�#1�w9������M����X��+8�0j6I=}br��%��t�]����S@܏(CvJ,��ձL��C�Yë��Co1gN7�K͇�ԋ+�Q��W\*d��ܷ����TL͋��L�ª��/{WbΜ��[�u��ӷ�i�vX���}ل^���ޫǚz���tX%�؜���N����^��lc�!���Ť)���ڭ��ٹJr�5f�q�ӳ�̮x��G��ZP�eԥ���ܝ�x���M�%�w��g�`�j��a�(���0���\/��C�u�9λ%ô5%}��r�΀��S�N̠�<�OD���4R�����sVݷKZ)���.���7�h�� �%���_V8+E�4,��l�y�Zs���x�������W��R��RK�j�.f(D�5�^UL�4��v@c'-^ty%,�[\
�#�&*���|%�ep;o�)��Y���H�I�Ṭ��X�v���)�v��꜇rӘ�*�h�Ȣkv���E��o��f�NUv�;|%Jqԁ��{&��W�й6gr��f�[w�����Qg$U���ݔ+��J�:'m
�f�F�G��h�r���)�&j/�,O�$4Ӭ���@.��t�Z����[��GB��/P���m����u�P!u��E��V��+'��Z�����r������S2���>��-�؉�\�L��-���Ŋz�Ky�I$Xj�˵����<��y�nl�:�� �/�H����u��ј:rYx��V#�U�V9�-�l�07\v�躠��((;�aU.�g���IZ�[ȟJ0.g6��[%d-Y��T"��|YHb"7Vؓ�4�"�q�X+��N�Übw)��\�T�l}әXf����������3mdDpΎ����²���_e�=ݠi�U��K�I�Y�9l��uץ�wղR=[n�vA�q�b:�ݺդr/e�Cz�"�P��S���9^��c�b�:d�h�X�6�P[��@@ �����X1ǽn]���h�tlL��+o1Ͱڵ�i5ٺ���}�3d��w�p��bT������-<}�����:���t�e\����e.�g)K���7�&�v��:sz��W�'^���u)��ng7fmX�ElǱt��H��a��\�u��s�v�3+�z�����x�&��]��:n�w�΅�4� r�����
b�'3��1�G>E�B�v�r,��(��bU]L�2�,���T2*74V�wM)���r�o�O�Xii�]Uq.���f\�;VIY�FػGt�� �:�.�d��8�����=vIIn84L���a����Z�Q=�ƫ�KXڕt,;a�ή/#�!3:�ȶ��#�>�
��M9�r��ڕJ�ׅ��:��ʥ�F�$�m��˫L��Ov��(j�yV�z�C
�M�t&���-��)��[��.�S��S���,gU�T���˄�!���4ؖ��K��c%j�F�T��T�T��!�N&Ƌ�|%#�(�5mw=
�����VR�k5�d3�JW��XY������9rs�秩L���3y���r�l�Z��@�0n�ˠ�Y�7�������n�>EU���s�f�`[W�Vxd�7��U̸��;�a�ar/ms�LLM�nMzw*b`0dc^b�;���mB)n�g�ܷ�և������EÎM{��L���E*���ݵ��oc�ݗL%1+�����f�6ng;����b��k��]f,�9��a��P�]�i�[��.D�j"�$4�m�H�����ӗ餁�o"ﶅu�o��wǝs^�	V7��<�:ڃsyЪ���Q2i������tGrvE����6���׵�h���6�"9�����\��n��hķ,X�|G��vTt;�.�H_+#L�aoY�o�.0MX���̣RȹW���]�3�`�H]�<��%�*�f�|yι�=�|&�o��\Ww�G(�YJ�t�0[ޗk���Z������}e�M�Z���U��K����4K�� ��&oe���Z{Iӕ�� ��;�y�Zz_̰֘r۾.�N�+�u�qL�J����BMx�
eqp��ٺh
�4z��_mf\�;����;���4!	�(�}X�
���ٕ��F�&��q�w����	��������v)��L(n!��fgeN�m�}'1w�g�)��wy��n��a��oa�d��nt���G0���O&����� ����ͦ�3�hW,��D-���+�+Y�ϩf ��h�c7$�)��Z�msOu��ben+�V��5���z�wsJ�6���V9�6�t滺���,�ؤ�)q� ĳ{h9�uh�5�C�c����s\�0{�0V<Yyq�E��v��ـ���f�x��-�h�.��@��yh��2+�[W[\e
���,�s�/pJ�BfާG7s�S�+1(�F2���8��P�z���]�t٥�3~��{�N���	!I�$��[���\\�y"�{��bYy�́-ή�u�Y�}�A�$����qT���bܣ�l��ue�Ose q�۝زf����[Kֲ�v���V-=�9s����x{(�5<���yr����m������=<�`j֤5j�g=�M��:f9ʍ���tH[:���,g�q�`���c+�\���#,�È�u�Fl\��{u�vZR��P6nݮ�v�1��z�7���uͮ7.��؛��۵�\�mc��m���{�4a�)�si�u�s�vx��s�g��;v�-cO\�N;(lQ�m�)�mb=��U��2�=����\�g��x�d�a���JgvJ�[��"N�g;���j[��R�X��vɊ�H�sj���h�m.�[��ma���W*�$��wm#� ��s�)�.���ix��dqr�V��lk��V��x�>#���kOdR	q;�`�q����c�rc`��0���{��+��ڳ.�[M�c��<�v��=l�Ɍz���%v�p�r�)�p�#�p8h� \în)�7ZǤ*6���y�Z��6n�j��um:J�uC۷���]���L\k5�6�L�<��ޫ�U�Ӊ ܏@��=���cE�������	��&n��f^{l �3�v�����Z�`��y�Og�����9�wV�#]r���n@�#�'�7JM����>��݇�<Gl��<so]�[���&�H����ۜ����7G�6݋�����(֘���'�n��]<]B6�4v^���&��UGWm�c���{p�m�!����uq��j,����4wl=u.v�t��t]]�1]t�$&㡹�0m���]=D>:�)�I�p=M��E�8�����[#�v�@�tvڕ]��<�h�����6 �<Q��Á��:��\�N�݂s�'<T�-��sú�7G[�յt�۲�9�ewV\Y=bS��f=�����\�:������#x⍣����ݶv�����4ݻP�sa�W���{=%��1ȑ�l�yNqηN�Kv��'4u�k�3��Tƴs�7	��e��*ݽ��]O���/�ݲ�X;V��ċ��62�͞;�ta���{E�3{tzY�kt���)K���Z��gn��M�m�#P���1uֶ����n=<i�ۛ��ӦK�ȣ�(N�s֨���`59:��ъ��uͼ��5G��ݷk���0�^xrlݳΉy.��	�<0ƽ�p��<��H8��v�$�[��b�`zy[e���D�y�=�mv�́����m�6ڴs밊>h�\Go:��]:��+�l{�[uV7O#��62e��q�\lW���YHz��<��9���/طR�l��t)��D��u&z�ۙ�K\�vG��;��n/m��b�m�G7F�xd��x�/l�LV72�����T��q�&v�M��-g��6�)���3��z�ϝ�g�x-��Cn';=�vM��nۓ�P��9�^N����A���5���I��<֖�a�qg���\ε�G;x�hB�:A�Ou�u������u��#����1r���;�8۞;kW��W:M�D�{ ��̹:Ku�H ;��1-u�[�q.�p��Ƽk�\��f�k�vu�'OPpx6c�ќu��sv8ͳ�%�3�����cy닫z�nx'n�h�y#w���m������u��ˆ��M��Nx1 V����Ys���ۛ�=:8�+�{��|)!Hn�ʚ�0�y;.��=�ɲ]��)v��\�Xcn5v�˫��W�&�cn�ŀ��7��Gx���<��9ݽ������lv�Yf�[�/a�K�9�0�K����z�����H�We{p�ׇ����cn֎S��`@\ �=qB�y̔��
����+��k��̜��:���vr�N����s��Zy���y.�b $��e�ջb����m��|
�����cv�t�q�ݭ�ՠ�[g��v�`�{=��=q���{Z���L��Y��������޼*�Xv�����8z�^g#�X�h��m�Ts�Vq�H�� �����[xL�wE�k9ex�ݒ�gc��Ȗ��Tl��6pțF�8����筹���v��YM�C����s�l�bRG�ϵة��+N8{�.<�q'm�p�V�����d��a�w;v����r�X���o���mm��벷"����v����k��e�Zy7�'ZM�Ӷ���;\��;q㞺lg�5�W\���k��.ٻ8.3��<y�ڃ��^�=Ǻ�m��Nv�y�1�:c͹�u��:��M��iI
���w]��n�;v��{�mC����iI�Ecz�]�Y�u���ͻL����95�u�.�n�S�mτ�7�Nw)��ܜ=$�/�K�I���9�fØ��Yn8��3���n��<���͓]���f���ށ�۷K�-���w�xu>l�� �9���ĲNy�{V�+s��c���s�Gf1�^��Y�-ѯ&�2��Ƹ��v�lkV�A\�M�ޥ��G:�	]rv��˸i��qh���5z�v��r��4GvA㣚9�g�Y2g@��u۱n�ɺ��9�o;N���Wm�;�����v7����=�l�܊hy9�Gg>�`)��a{�{nڣ\s]�s��9*����7>9y���j2�rl��rs�vD%�v�rWg��;�u���c1��LW�(z�[�=Y���n�'oցv WX�<sֹ��Clr�u��:qt畕,�b�X�3�����;���R���g�����]��W��n�;��8��pj:#���λD�u�Fܴ��]vN���W���W=\�On�nf	۞ݍs��{vV���`;��O��9������s���ubJ8v��;m�s�z��۶	�m�;'jgKv۰���]�#[�E;�a1�S�m�GAWd8#���cq�܏[G�-����:V�{,GN��ʔǮUy=u�=�n͖�u������d�6�c� �ٴtk�ګ&^�u�-����ݶ�s�۱��Kxć{\�ݢM=:�;g-x�z��8������p��!$�a�b͎W]��n\91৩�hv�^��5����k�K���f��n�\�d6u=V6u�4���۫�+f���n1�B��U�*�cH�W.ݨ�1cC>_��8�qҷ.��<n;���{uĻA�cq��)�7,S��*�\`N���A��۞�g�z{Ek��L��ƕ�a��z.9�dK�6^xzW�z�9�=;q����\r��m�`��V�x��ļu��=�����^����\q����[qtm#����88N1�{r��81�E�;e��ȯ\���'���m5��<�K[:'�]<W�4�(v�bN�z���p�ܗa�k��\�����;>��5m�r���'k�E7>9E�J�\�\��e�`H-�Sc����u�-���7n�lv���cF�\:����.��͌Vx�<ѫ�v!BKt�xkq�Kv����v:�]v,����a��&ዳ�NܖW����u㛂�ي8�n�u3c��{.�N.�an�����6��,�n�E]sѼ&���g�r=��H���;�v�W�l���{^�Bⓗ1�n��T7<uu���K۷T���Ơ�٩zKl��`��rh��6:���Gk��RW��&��R&�5�m�!�nbG������m�����[�V�� ݙF4�9G��+nq݃��F8�@�*rv��q�nj����m0e�=F�ع�n"���ܳ�����fNy�wn���=���e��g�ǲ�.�c��c�{b:w�kc�f�:<t��{pM�\d;s��뫗�Ň�2�2ݢ7�wqc�+؎ ���Woc�[�N��vk�)���h�m���^��jy�ys��c�m����λ����q�]p��3�[�Y.�:J1��6��D�:�����\ F��[���`º72L�IxH��m�,��N��6�pY����:�ڱdS�k�g\���q<����@݀��7^��e����71�]`�O/�9���W�9X#m��u�X��<v�K�|7����LݘM\�j3n]�I��Y:y&+��{Nm����|�����M���&�$7Rݶƙʂnvz1�琱������+:��_7=��
kk]��O\x��Ƌ{�x9�㑻z�p�[v{��+f�6��r��<�v{s�\� �1��u���>�!�0qi��5��m���.�WF�x۳�n���T=<��K�=�d�'>M�;K-;�/h�<�7vIx���������o�h��<���h�us=h'�,��3�;��]l�U�y�����wA��'a<�0�<�^صՠ��k���; j�SzI����p�6��J��v�p7�C�ٓ=On�P7&y�vGpO=��Wf��g=�tn�t��m�91u��8�����5˅�c�1ƥ���:zݨ���Ѻz:����� 6��y�v�^����49����9�[��L(�М�'�P��N��̹(,�u�4ݪ]�+�c��cf�L��Y�y���nAr�s�<�&��.��%
�7l�n��<�e�b�Ƭ];�� ݇�pƌ5�O{un��q��V�G�k�\v�^ڑzt<�Lw5���d^/n'�f��'�`\F�Ȉ�ԫ���ݹL�۴y܎VN����qً�����Y뮀�N`���qs/m�4�׎�����m�Z5n�����f1���q��,��4��Z5f^���em�3�G[�/b��BV�s������0v�$��=uJ2�.n�p�]�izNܩR;v㓚�������ԓ�ϋnn�a򽮲5��붆y,�۝�8�]a�gN�%��u�pB\�EY�f�K�]GO5�ڛaa�),��Z�ګ�om�����ys&7(���.5PDr�-�pf9Zi�T\V�Ѫ�Zp�)m���YiQ���U�QVѵer�m��.LLIKkR��\�)F�c\�Z�L��ƈ���`�8
�T��eaZ-�*	V[B�aLsiR��e)r�r�R��5[k�\����\ˍdS ��\��U��m���F�����2UTfapQZ8�-̮&eb5�����6Ur�&��eG2��T�h�sUQU[eb%n%l��.5C���q����pm�vGx)��\q�s-2�l̖��ղ���r�L�\���-nf��jԨ��(�ˋ�K+[j�UUVڕhTU�`�9�b��ѴlQ+EUbc�jb����&\qQ��c��VYR�%h��\"�q�-Drۗ�Ym���eC-�&YF����\V�PEE2�f\n[Lj�ebcLLr)�����jUs-£���G�\@�DJ%jZR�)pTŴb)Z���0.P�$�g��A��'{7Edx�l���<U��i��ۍ�&@����W<����>|Z�p۝��W=�u�ݵ�uj��`��n�=<k��v%ؼ�l��Ӽ�K�ָw>���p=C�+�\��g�\q��Y^�$s�=ru�xϞ�y����ak�`�)^��R�R����۬uqӛ��ڶ�n�kŗl����;Z�9�i�=e�[^�uclm�v�[vϞ�Wq������v�a�(Nu/k�s�V;Z�7%��vtOc�۲kg��痗L�]d���D������q���]���m���[j2W�::��Gn�Vs�;���B����b]�W|m��|{YC�n��r�N$�v��a�v�)��`�X���{{�-����i{M�z_<�'��xמ�t�xnve�x;�&�;�3�&��x��<�Uu�ۋɓM�휀6ݽΞD�ֹϮ+�v�v;Ry��r��
��b�#��S��xʇ-mɮ�Ļ����m���J{c�ۍ/E�qv�^ܖ�..��+����;=�3fG\DF�p;�����Wm��1#�85u�X�L�:Ӯu�g��O��҉B���6i������h�4�8Y�!����S�5�5��U��l�u��ݣ=�ױkG<�b�l���bx@���[Z�b�Z����m'k>����b����m3�]�0su�s���{i��<ۤ}F�76�ӎ�m��;WA�W�͌on>,���ڷn�u����xc�rq��N��үh�;MѸ9z��N;�P���v�Ӹ�ݮ����7mڋO����Eb]��x�zzC�X�{-��f������-��9���X;y��/�:�>��H;&�h��{@��C����X춫�=.�<ݼt�lnP��rX�Ah�<҆9x3��I��u�8�:����n���ܷ3�c���$l�m�X�^ݼ�j��H�un�ծ|ώ���y�]Yd�k����{ӹ�:�W��s�y;q簇'gÇv��P����`��L�J�Y�ڔ)�!�.�<�����d��N9��UrP�6��(��2�WyD���ݼ��{�<�mQ��0mi��L̪�s��y\����d8�������[�ͳSUqTG���<p����g�qɶ}�����y�=�vcg���n[����D���^����幠̬�.��-z�hP��j�P9����#:O��Vl���?f�zŋG=�&�-8m*���U~0{��w��m���w��$����I�ٌW��	)�x~W5��o�wKuȣ���7|�wZ	$�tH!n:���W���A����	'������MH�A�	^�����~3I��~�OČ^�b�$e�=~�;�v��X磌n�����R��<or���z��z�P�ǟ����ٽV	�����	9}��>��z�w�L٧����N���v)S�S����Y6Oc�i�ƻW$ �D�3=��26c%�/���1�� (
~o�}A��P
�<V=� �x����p���>��j��b��j�v�����$�9���G@��jW9��n�w��,���˖���*U�웬�N���w/]�s�m�FH���3k�g{�Խ��g��� <���>o�
g�]�C��?zN��D{�a���p�n��������fm� ��c��2���p'���ʀ�����"��s�o0���i{��{7��ʛ�9g���� 
^oʕ�w���5>>��ڲH	r$�NBh��eY �N��,V�j@a�.�
�����}@WI޻3ß�§�r�5�$^E
%�q@�w�:ڶ{t�v����O1�K;-1m굸�Ͽ����B�R����e'㷗���$����H5�Ycݾ7�r{܆/���
�א���f
1����=v	 �]�m�>g����
6�_P�U�w��~!��wd�}B�v�q��bBV%muݾ�_��O��Rp�+P^������z��{y2�g��A�����=]L��Ud���+,��X$��k3~/v�d�E��6���]�����@P^kڪ������D�M	�&���<*��}���X6m =o���+ޞ�P��"��{^�M\��M�f݀Ht������wt�e� ��Bz���=�*W��n�  ���� <3�˷�=���~���������R2H���oni�UhN-̆M�,5��1�WR�F������Wlу�XT��� :N��� (xgK��P�J��U�vH7���X�9���(������P�޲�/{�zm�Y$��U�A'�v?�5�Qt�������6C�0�b���ZIge@~!�"�*�>���I��z���>3���C�L�?�� »�/�A���ޢ~.{=V	$��;b��;޿nn�#b=(���Yב��U��������h���@�$�ⶃԛ��믏O�"��3 �	�����
��bF�E���^���o���{�bl&�p8�b����*\=�x�g�t�j�EK�>g��$���w��g��v�W���<��(�ߨC��I��צ}Trv��P�n�60\���p�H'�˼�M��Eȣ�I��d��k(Qoy ޞ�`�rq�q*(�B��drd����������nĿ{�?{����A��n: �׽vIk�F�V�jﳼ��fV��/@`�����|w2���v�=VB������v�'ܡ����ɥ�:B��b�{3���(TZ�z��=YP����^wz��)Kv1�ί��އl��GA�vkk:��O�s���]'��o�p����>��J�
o�볏��� �)��$�٣�׹]Y�uhW���������mި#KVg��Գ�+�y��9ʡ���=c�C��rs4$�����n$g����3i[�sא����S�Whc�y[�o"�Y��<�Y�h�0����+�;�o5$��ÐXƣ�E�ܧ��\����7k:(�x�OS��ۦv��3��>�y%��x��yz{�'�&�g��ty[�m���]���h�N�]H�-�����5��m�]��G�5J��QB��ݽ�ۢ��&n��)z��ͳN��9�<9;Zk�n�F�s�x�[�y��wkOmc��ݸ�s��I�[_����鉰�B�1�ћ��]�,�����r�+ē
t9�7wBHu���y��čGv罗`�Qҭ�����
��w�C�?2�}vA�ޱ��{��e�T1#y���r(�RDJ3 ڡ搯��s��@U���ԗmg�[��נ-��(
�����KC�`�������oW�����ԳI?o7�Y�}��]�A ��mvO��U��D���K�Kӌ��>"%w]������=��t̮QU��ޫ$�������=�*�=ư)7{w��ey�'U��&K����.���lsZ�7.8u�\ݘPP��0��x�B���$H0�ƽY6��>��P 㞗�0e[RYm/y H'پ��1�4HTF:4g��=P:����{�]�*Y��{�!�h��?�ԒC;�`�xj�+xICvW��Rk&�10{��o�*�J��ʠ��c�]wr�>|�ޑ  �{�P$��մ'֫���&���%ݭ�G%���9�e� �㵴!��6u���.����K��o�v$q�mB�g�H�D�	�{s�İ{{��$�߲�� ���������ׅ�W����Woz���ac�`��L���|or�$���_��wwo���/3���P�O�M�	M^�_�^�{�"EQ��̠j�ȱǍ��&��]p8�V#v��NzgX9�^	�v��/��}��S�����ۿ���>���IW�����b���U�H}�d߰��!bI�"w`���� ���V0Ǘ��*ڭ'�@$yzk�6��_u�M���~���=��M&�E�
��_=]P��~�~#iMщה��<�83�0����Y0��y쁈�nѝ<�論�<����E���	e�	[��o�f�^������.O0�6�@*$[��]ɯ ���P�*j�%���-�BF��s��5��I�sU��U ~����7�ݠ���+ü��5W���"Q2Bh��$�������3��ؠ�z�@ڻ��o��utscg6{|+&l~2$e4�l��qQ��lC:�h�ėa�6�]N��]��t�vn�����01 j�7�$��]�3=ޫ>��mS��m�����`�ſrp��4��.�V�I.�.,�������=��H��H {:U���K>�+9�̚�(d!!vj^���N��H$��;�w4�+��S�a=מ�$���H�f�I�Rb#2zp�V#~��������P��j�h���}2�-
�i[����x��H�`��zߣ��&ۛ���1�����
���(��3q�\�Rݓ�'9�@9/����WD%�~��<ٙ4�f�J�7w���]�I>3v���Vi??:���[�|���@��:me�E~��ཬ`��o~y�x�Gm���n��E��Z3�u��7��B�p?�!	+sB�?8�$'���ąP��j� �!ΗKy57_{ۻ s{�,z�K=��5v|w2�1��yX�M��l�Tw��@A��  �S���{���ɣ�-�'� �J"�����$p�ڄ�����\fz�.^� jw���A�7y�+F)%ȈB]���R�y����D���k���)��� {�=y�y�;쮱�SI�b"2i�=�  �՚��8;�ׂOѴ���I��(M~J�������x�u5ۚ�;�����4�-��R����7�v6���X�Ս�s:���3����w�Hf��9�3
�:J�d����F~���Ŷ�iݞ(lw��꽷g���+cYK���5�9�A������q�]�t70ݺ6c�=���a豻0�UW�>Ӯ�\s��-�K���Gcll���
LX�7n��*t��H��l)�44��m�q-m���\�h5À����nF1�%��YF��M�v۳-B��S��&��ny/l�3ha�@k�
l�G��B#���d��)��x9\��/6��_\�H��o�zF��0��7�+r쟁'�ݨ=�����n��5��z�I�=��֢���\����rœ�z��v��w��^��#�~$b���>��P��/(�f�T`�ު�p����*�.��<#{�`��
k��
�ڒ��/.�
�vЀ�Oݵ��e�rp"D���*�����J��{h_��� �edHP|����`�c��Z�,f-��E��d�#(�b�oh�	}��_�(������bj����J�����p�^�e]xK��94��0@d����뫯g8�c�s��K���z7/Nb�lx�����߿Px�z"2{�FfЀ��ͱd����s�"�u�lW[���O��g�_�v��i�JP��������D]C��lz�otپ|��SB��u3%�&�5Ý�;j��A NGL�L�n�$��(]����	E+����0��ùއ�B�{\H )�w���Tו�]���d6}T2�P"�e�BwF� t��@P�sǖe�?[��_��_ �{UQ z�+=���5v��^��ۘ����gU�	��]�A'L��R���KƯEC�_��ou8"�B�Nu�z�P��}z��5�V���� =��]�A'L�#�;{�4:}����e��<��^۷\]=�t�W:�(5�:;=\wT&f�fI(��&o�5u�_og�^�I�k��mo�t�/|���Oč�{�`�m��A&!2(�E�WПGא���{F�z�dA=��]�H$3rW�-U�������͛�Q$�HLR5m����O��nЇ�/�L��W~▹\u�z����H*/n}��2�V�4���Jwe�r�J��;�K2��B7اM�tΗ�Edj����F��ϊ�w�\Z#-�WwG��u8h�*�nV������q��X1p2>y]9\�bv����M���gf��Ë;	{�n�T�N�)+��CU�C��R����|GJ���'X��Q���	Bzb,[����;9	���h�X��aw7./�J��qu:W�GZؕ*�b�Y0�^��i���&t���[؋=αN�R��R(����p���t���Ŵf�v+ ��e+r�gUq�Xn
��A3,۠x@���)-�ժ2`��0���8��y%���i��h�3"iA����3�W�qӷ���bR�}�o_E�������A���C�b��Հ��!N|3�Q�_�Z>7ad�R�vŐ�� L=�R�&�p�ʲ�ob�t�#Yah���%��Xڝ�s"�����iQ�G�U��_:D�l�5�ں��ɕ� }���+R܍�c_k�|g	0)l^F�:�1˒�q钮��[wQ_޾�|�U>�%�����r��k�%��F����x�,7yw���wYβ޻)���u������M��0a޽{��r�o�3�N��G]��5%m�h�P�4���w:���cbo��M��C��#;����nK׵\��������]ֺ���Jf�κ"!fuN"�eּU����ձҲv%�U��Zmj�h��[;���(�nn�מ���[n4�[iZ�mYA��1��S���n7;�'�Z�[Z�U�R�����0p�\�ek��Q����aRZբT��QEQJִffb"�&%dơJR���i������Kj�ʢ���1ƊVV�8cq3"6�����3.6��T������Ō@��̮.2�eJ�cf)Z�\�d�W-3#���ZV�\dm�#�f%J�D��2��@��S�g�ropy�q�ض�UZ�*.+Dj�iEQs1,��V�%��q-���KmimmIm[JZ9h�U�Lp���U�խ���7q�e�1̱%ܳLr�fU�B��4*���RUG-��r[��66ҥ�\��Z�+F���VX��DTqh�ֶъ!V�h�Qh"�,j�B�`�e\p�8����2��ص,�R�TE11�)�QfKS�Kq�*[B�X�-*\�-Je�LX���.
�*�e��R�6[)m�-�V��b�QZ6��TS�䢸�)c�n�V��{�~X�����A 靵�1V&���\���va�垉4y�)����+�=/E�k��e���
���Tu��*, ��X���W`��ʀ���V�[��>�x���P�=7(U;_��Ð��\Ј��J�q:�1v���b�^�C���{.I;9�۞sǮ�}���7Eń�~�fm� �p�ڄ�H�Vz��U�]e���R�Y�ͻ�3v�d�-I aEdʳW[�*g-xg��a�
&�ޫ$P8gK�C������x��W�����z�L ��r��u� ��6Ő>��p�9���� 8gK�v�$	���M8K��w����D�E]{X ��� ��_�v-\g�ɦ`�9Rl��qj��^��E�[v)�5��z�����ހ6�Z��Z��T�9��Im7�p3\��|l��Hk[Z��[Hh�f]�;;�VP�d��Ih�U�1D�=՛vH'ᙽT�\�s/W��"�v8hAۏ&��8��hq���{[��`7 �<Sc�Dm6�<�ޅ��F��ٕ����C�C�缐�2��]rR=����뿉-�GP!�b���X��S�;�MӁ����H�Vm�'�Ff��`�+�(%����ͲԎQ�L�������F�{�`�H#*#4���]�]�J��>��s��V��&!.(���mq=�:�� 3۫iU�~�����G�� �YA>���ۻ��sQ4�,�4߼�@��v�nC�����@}W��� �缩PSk.�OtoxOp�j6����/,ջ���uM2M�d֬��7:��KY�K�;�u��y�?m;��tfd�)��s�����|�ǂ�0<��M$�Ę�&I1��h�< ��
���b�j��z�ҥ��
�s�v�.��:y�'&�n��GvMl�u�M���Ɗ�/%��7<�	��i3Ӱ�lSuq5�[�^��wnM��eSnNz'���O�*�ٌ�����2�vyqk�uq��`n�;&� w=cDv�V|���� �[n-g��-�7e�A�;�/m��C�<��|>=�)7@/n��jV�F[�ėU�u���[p����qb���s=(�;7���~��2Ka����˳�'���g�5u�#�C���~K�+������*�`U�U�]Y�<=��7Q�!��c��?7=޻$�^���;=^kr�;Nz�qo�$Q�Lm��ٞ��F^�$�����W_����~>�{�g�>��}��5��#m�.�K�w�ݧK��٬r{}B�?j�����]��E~���$-���[Z�L$�����h�v���3��멜��);�� ��W���g����f���Dl�o#����j{tk[���<y
�s\�u�Y�Wm8^�� �K�'�������a�7�3rŒ㷻X*��&��A=��6p?u홵�=� 	^�-RX<���f8h��r���ݮ�?Y*-�i�yD�M�}lu.�U�"�Z�߈�®#kj�D���Dt�R\+���ᡳj�ӈ�G�w�(2o*N�P�Q �r�7������[��8��,TEc�Hb#P�]{�$mfz�Ab��1z�]ꗃ	���ڀ�v�����I#q�E������%��4���d��W���*O{o[�r�P~y�U ,kv������#��Y��������newx��y�'�n�:�H����<�Ӻi���>���_����b�v�1�x�W���9'^�/<���.
P� �1 �����LBY��L�>�vm�d��n���ʍ��mv�Dp��� չ�D�Y�i��EHM؝^�k�#��˓�5�#��
�' ���H
��J�������C�T�� �Dm54�ۗf��t�j���[t}�g��B�YC��^U9*��q�4���i֔��&�m\�p�-���J�v},$lf,���GҫÖo� =�ߟ�I w��� ��� =�Aw��ʺ˫)P���u�2�5P��w_��ݽ�@ ��S~�~�9K�W+sOmU�����y�P.�������k��˧X)p�w�_�sZT+�=��9ͪ��Ϻև��,�9��o�a	��,D�F�W�z�9漴�;e�-��n������o=���߼�C
F�p�;=�������$�~�ٮ�Ei��Ψ�����������(����I�L28��!��[��v��u�~�$���,���h@L�:�{��!<��EU��e��E8�O]㗝�*�o��@�ݳu�/��������hB��pB#i����.�[����Au��A#�>�_���!H,�{�|�p�5���������ww{/�A{	�c?\{�L���Y�\��fe�m�R��S��̱w����eh�n�y
Ċ�r�l��<��U}��A��P�����H,:~�-�g�..�5�^C�;W���n�pB��Q�ts�~�>�.�oяw���1UHQTn��è�������r��KῳW��G՝��{0d�K�%`�+����<l���c[��zqۦ��Y��v��ْQ*~���Q�e������vq>+(�R���vq�hT�
���}�>�:ì+�ǻ��g`��s��ݝH,�Y(��}����M�_��}0�ֵ�ֳ3\:�Xs\�퇱�����=G~:�rK_k�x/�$/�с[>ϻ� i8 T��	�>��ì�%eJ��=�~�����?~���l��+
p�{�e�������pa]߷�a���X�H,?s�=��βVT
	P5��{�<���7��>�����F���}�n�m!m���Ϸ�`V~��c�1��/ u:$��s͝O޽�s
���-���4φJ�2WW��l�ɴ,IP�J����{�u�F ���߿}��3�׾�����3�~��VK]�y��������9��ff��e@�������XjB����߾�ă�=;:��}��|��ہ���Ry�ngFJ�2T(���~�b�������8�1��܊�.�ゝ��.wT���]�wt]<5�f���	�4Ѣ��`�E�vn�����<Y����k;��7���������>]�x7� �.�E�u{]X�Bq;bM�;GU��sv��vݑ�1�`�k��^��ݜn�j��.��1]K����rs�KkIΰ�88�.y"݋I�˻]��ɼTu����w�݆ٗg��`]�������2\����x�خ��Ѱd��%`�ݳ�c���ƻ�38�N6�z���7^��=v��"垃�|R�s�g��I��0���m��2�{8n���.�u��&
�U����m�r n���[�����=�]�p��!��
���͇H)*���Ϸ2u�Ĩ}���:�ؕ�	^��������~�4�W�X���B�ü���ïc�Y�~�[��s1���dYz�ߨa@��?+ﳮv����+���l�2m
��D���s�=�:ì+
¤�y���l�N�Y++>랯G��}gg���Q /���XRMeu������?~�8��5!e����P�C���>���������'������R(�s��:Ό����y���q ��}�..8huu��6��»�o��s�����Ci?!RX�a��y�gFu���Q*���}èJ�R������o��~|߿�)�a�^�+�=��[�ta�����M���l�t@���������gM��g�sk���ޓ�J�;����+T����8��VJ2�V#��u}��(�.T��a�߽�!"-0����x�9��"^Wt��֩��{S�qv���&4ֽ�����k35���P>��ϼ�a���!m���}���-)
�o��}�'
���~��߭�9�<��s��H,�%B����Ρԕ�zb+_�F����~��|EQ�����������aw-���wC�#��x�;X�s ��#����TJ���WӒ���.f�gjnPXgo#HX�ͪ��2�<S�E�ᕕ]�H�<��~��3���Ĩ~�￸u�R
A|�w���� ����k}?���/?W��O�"�nw8Tj2��3\��ğ~�϶u:�YY+,d�������B�*IXf���������ϻ����a�
°�(�y��u'P��� �_����M�Y����ֵ����L����~y����?�Ƹ����-�y�y��t�-)
с[�{�yI�
�+y���gw�wX�a�6�*5��l�VFy�S)�eu5u��4À»�o�Ì6�R���vu�d�����Z�sۣ���S_���:��+��Z�����p7H4�-�������^�
�:]�v�7�O���3<r���G6мd���j�7<�K=�Z홤�c���M�w�ϡ���ni~���&��l�u����d���}��M�D�
$�,=���:�0�G���}B��������G������:�d�������wH�����ff�������{��� �5�Gt������P�>	!�E�O��}�$��	�>��ì�%H('�<I&_CZ�s�#�O��و���Uњp��:ñ�^��a�IP����϶t�J2�Q*�>�;ע��bQ�T��O�}R���Se5evVd56�!�&m�23�%��Y�tT�B�����Yťuy�}=�Np�ޗ.ѯgҹ]�i���;OPմwy�����o���Xk�}�w���A�!ia�?���:��Y�~p���ڌ��@���F�K���8Y����%w~��82mT(������܇Xv0��=���$��3�Ad���A����w'"m�����kV��fb�P:��y�n`u�
��g	�l����u���[��~r���T��y��ԂβT(��{��:�Xw��0�'����~�h��6���@�2�7m��a9�l��A�N�Я\S[Pn=m��ߟ�nNxCSWZϡ�0���p4��
��V�����:�FT��d��}èJ�7��;����V_�ď�:�z��!�(�-,;����ױ�[5Ǿ}m�F�m�/ u:�z���:�Yђ���>�μ�7g�m�ַ��&ТJ�IXP=�}�u�F�T<���8��
ϑ��oU��3�3�H���K������ Q�~Bۑ�`��'���m�
Ԃ���߾���BҐ�`V�����bW�i^�J�}�� G����~���:βVQ��by��l�IXg���`���u���~�Y�{��_h��!�&!R~��6tgR
�Xy��}é�ְ(��������-��O\�=1[�b�(���s/�^бj��7����s�_f��i�U��H�9F�;���X��b�V�l��u$��Q�n����着�����ƾ+{��ۇ�n�_߳Kt:\s.�� T�O�w��N� ������vr2m���������!�$�;��}�q�XVaRPO|��u'D+%ed��>_���D��W?��ǽ��߁�C�8��W�t��v�v�f,DeM���s:���ppml���k������jJ�_�����%a�y��`V�-�{��}���HV�
���}�'*s�wy��W8Y����}�u�+(�P<����:$�,��^�FS��j�Y�i�Ww���pa��B��c��_������k��nd�eH(�����P;�,k �>_���!h|XY�ʬ��3��5~�����`V�~��n�2ۚ^@�tI�~�͝N�
�2VVJ�}�8ɴ(��bJ�s��\�~�w����F��IS�?~�gRtB�VVJ�y~ί��EDޏ P�6�qP$`�~�����˻��.��g��(�� y���l�iJB�`V���� i8 T��Yb{ϼ�p�3����]���f��L�%B�wsݝC�J�?t���Eth�8fna�����0�AIP�=�}��:ɇ?_��:�s��6��*�����u�V�_����H<�+y�Ϸ=`U o��}þ~�����P�e�Tg7H3�ml�atz[�dݨ���]`�5�A�D�c��<����$�|iC��5v��!�}4���p��˫}�p'N&�˘�Y{ۍ��'ܒ��[j��>v��{f����l�uXeF�}��/÷�d� MÓ�o��/&u���� ׉۸	�LZ�$ʓ��-��gU;Ը&�;.�P�"O��XomtR���mޤW��B��{��kt4,��*�cu��]/>Y	ɲ*����=[�M��e�\*�3�t�*<�觽�~��T�H3m��k��,��t���������s*��o������ٶ�^]����*����Z&\Ӆ���O��W/G-���Ʒ���Y��ݻ�ӆ&M�](��DY6�(V%�I�lѾ���ib�	˵���e�ê�
�j��G���d=d�s��!XΦ�مA`։y���p����.u�
A�U	%5��yփ���=\]���=V��(}�o�d�t�4u�x92��{3��5W��^�콜kZ�]���}W�W*�!�K5�JѳTgu�!�yV[˅��s�m=�eN�q��[�5�����1F5޼�]��1KF�E��*��؀�tf��@���\��9+U�*��!V���YfdtӘs�����/�	U�5n��))�Ԩ���ef���Y�_q�W��N�/#�&N�k!	��'9Qޤ ��GR��/;��H]�;n'�ٲ+q�,lw�����L�4����KVnu0�q�E�dW�1�mk�&�Ac[�Z2g%�kL�.�V�f��cl��,݇��>�^"�DKb���Y���*�e��%�W-�R�����"6����ҔR�ԥ�˙hԭnfd�S13&J��ƥ�`�m��,Q-�)�KQ�B�����i�qQ2�J�Pq�Ŷ[-�n�q�`���q܏' a�isL��1�2��R�q�n\�U�q�1Ĳ��ڵ
�Sc�m���L�<�`7*5���f[lR�*Vъ��s��lx�sò��vCe�<�Sl�q��𫳱����r��.	J���j"��E**����+TL�k���be�˙�).\)h��֍���[[�KmjZ�a�	�v�px�6��U-��S)��ZZ�kmPkc����Եh��J.(#ikTj�ҥZ�Z&``�f)�iV���
�2�)U+F�F�m�e̘�L�2�cPJ�a�J�h�K�W(ܦdl���;vl��{�v�r�0�JTj*Z�Q��*R�Z��h�q�F��2-�TD�[[h嘥�Geom��|?,�t8϶�ո��tm�S����kr�Y����e��qۄ�8�Y0y�]�T�bDn;&�ڐ�P�ͱ��;��y�Ɵkm�s�/g�v�i�V�Ɍ�ۨZ�bM�j��'��ͻu���/`��I�x_V7i���;�睺P:��d�nA&TVAM�]�2-��q�v�A���-�l���z���ͳF7Ftaxݞz���bxc��A�����s�H�ep����Ӷlqv�xg�ލ���	<k��ݧ]qy6Lu��
���v|�k{�s�Vv�z4X79�y���N�1�F�]C�c�u��x���N�5KJ`�]�=1�^��1p����ƺU�OZ��u��f6ۛ����Yte�iZ���v��YNn��"��e���ۑ�6k����c-���ͮ�<㷂���.��h�pd:'�Mݣ�O��ݵ���8�=q��xol��}V)��8L��	kM��[v���1��{dN�%w7.�y���{dn��$M�z����$�yܽ���ͽ���8hNʀ.���H�MwŻ�bӻ,��u^�$;�ڳ;v�^x�Js��#�v�{n���0��Wn�Ldw��vv�.�V�{n�l\�:��V�q�C�	^6v�:��l�둻]��E�9:3�۲��vX����i|�<�΁!v�`wn�=�1��V��gX�v;Q�9�/h47��䷲u�K�7D'�Om�ۥ,9�f���\�a�'l����9�s�W�7diz��=��`�l��u��w0j��Zw7g����ܙ�s�[�zwg�������*;R�2�F�1maZN}�_B�d:���)x����ݽ�/	&��6�����[s�Ϸp�ˠ�w۔�A^Y8�<�'Fqk��=�ܽvw%ۃ�g�r]ծt�ٴ�0�oZ��`͞��I��������cN��=�iԻ�����Y��<=���xGim<&;<\q�^�U�q\�qۭ˶������=��ɛXl�qT��7H깭hѫ�j��&mu�v���1��9:Jqvݲ�Q�˲\�j��t�������d�u�����v�yƝv��X��x(�J�.۝��(88���\�=GH�=��V0/7&��XC�7��DhK��C�u<��v�8�e��li����ۇ��\��E�q�<Bh�˺�F{R��qn: ^����ͫv��۞Oj�z�nW��?����͟Xiw ,U��[��Y5�X�:9�Y5��Wn�.�b�u̯��])�3G�>��hn�K�e�:� T��~���u�����%|����2m
$����y�!Ԃ�s[�_��7�ޭ�<I�7�����N�+%eH/��}� p������un]f��t��;���`PjC�e�=���y������+Fh}��� i �����q��� ��Ͽs߻Żc�ۿCg;��;V͚��2�榮�������l<m%B������:�P)�2i���=/?o��C�y�i i��,k����7H6R�{��}�u��՝���I�k�,�#���:�k��h�k/�z�Yc%r��l�&Щ*Aas�>�:ì*A@��~�gr��y���>����Ă��2��{���"��a�.E�G����۴���!A� Ivw~�v/�磎']�R�����H)�Oy��gFJ�2T<��q��3���g����<��h��dLn�E���q5Wms��ik���@+�g��3۞f�v����G�\k�d���|¿^��a�Ib%�V�߽��βQ��@��=��@蕁�|~=|��>z�\�����A���|;���s������D`P�[Q�ND��y��:�++%gt�?��������k+/�m��-6Vc�����YnC�G#�����
�Y�Z�[Cs!�[��Cz�g
����P�ܭ�;��޾�=p�!>��ۿ��C�IR��}�!��+
*J�y���H,�ed���{s;���{��W������� ;��a'�EK@��{�߶�!e�{��}����h���۳�|���y����~���$�Ή���ì�%ed�T<���u�+8k��c����ra�����q���w���nk��bO�%B��{���N�T��g�?}��t�(Ԃ�w�����a��~������|�p�с[9��=mn�5m�/ u:�z��6u:�YY*A]����C�p�o?p�CV�����VaRT��}��:!Y(��FS�����E����������.89^����뛷W�ۮ��A��1qbbDj���W�����ǀ(8�r(�	 ~!�������!m����g:R��h�Eu�X C�¬�������x���p�=J�P�y翾�Ԃá�t����isY\�C��}�v�GȀ��J�{u]}]��L�����ޯ�>T�_|���:��+�~uW����#�g�� ������|6�e|0��SsA�CmFe�
���{��'��d�������96��J�IX0���O�ۮ9��:�{ܱ�0�T��G����\�0V��~�e:�N�L����18kD�qW���������b]��oA�`Z�������=��R�%��Ͼ��ԝ��������q��?v��Uպ�R���|	�]_�P�g�d����?��y����vR ����m �
�����ì`短�����#5�_srq�Ovyx�+�3.�m&��P?|	~����}kOݯW�K�W�~��/;������xu�+�X5��������}��Ԃ�'����!����Q�����3#�Q������NX(��8n���zVvLӈ6����ߟ�1YѪ�4}��I�w�:�+(�YFJ�߾����(��RV����C�:°�syޟ��ׇ�~�I�>�{��:�d�+%e}���Nq���_��5qִ��P8%a�߼�a�� �=���y�Mq�t߷͜�������q8�R��'���w���R@�s7���OgOuw��ߪ�i�#�Ol{�3�!*4[����>�����* ��~}�γ��P(�~}�y_��ϣ{�3_��x	R�}߾j9H6������p��l�׿h҈�b�⿀$YW���a��~����%e+�}�FN!A%B��?o�}�8ñ�aXT����8��_����g���I:�N�՚Zb͗����$اs�+Q.70s[���޾B{np�(��o��q�R����yٔHژ-K{F����R�����dI���}��W�����e_{�8�@��~��s4�[�e)�H,9�~�{�(ԅ@�w��/���Y��>h�*��� i8�R�����w3���g�$B]�߼��#��g�Gv���Y*��9�nm+��v�n��7{���x�Ӎz���]�����	���O�~��U�@\a��
��Vo���d�ʁDD ��w�X� ��7�~�Z�����t�￷���K7��w��Vw|R1�҉& ���0���C	؁YY+?k�u���o=ǽ8y��"����g��H(T��?o�}�:�Xv*J�}��u'P��ed����w������̺��)d����� L���L�\D�=��=�u��R�?{��s���R ���7�ܦ��5��I�H,�����é���
!��}��u%a����4�k��f���+���<�>�]]�����8�Ib������:2�Q*����@�T�����{���{�m�H;�-�{�:�p�E���EQDq�_ I�'�~��N�VVJ��_.��gM��߼?~�?s7�	�$�7���Ì:°��ID�����ԝB�Q����������|,W��e˯4#���ABÒ���y+���o;AC ������+^������@��z���e֪u�����a�6�vQ�[Vם�����ww�o�[��ʵ�ύr�V�t%��9]����F�y���n�8R�T�7g��u8�d�Ӯ-i�]�j�n��p����[�]s]F1�=�<lk�`k�d�1��q�9����h7<�à��s���s����+si��V�kqH�y:�l%�偹ɶ}:���6�ȅ��g��;�y{�=Q�8���s�7W*��Sˋ�ƏrF:�C��/��sEc^�WN��j۱�.y8��e�5��(�(�B$�7��E�%)?�����y�>�tz��R
�����H[HV�+g����'
�W�צ�w�|L��<���R
A@���}��|$�/�=��ar�kNk��Am�߷I<�T����o������}�;��gY+*J�|���p�D� �]����!�)���s�]��p��쯇�
����k��u�1��N�M����ԂβT����ݜd�$�Q%a级�9������a�
�RX��{��:�Y:2�˿�ܜh�=��
&c�+�,����z�ם�;�֧<��:�������9�B�B��[�o�����H,�<��{�u��{�>�S����6�PЇ��߶uĕ��=�i�:�7Y\�C�:¿_|�p4��%B��~}���N�������<�@�T?}�;è�
�k���w�t�JB������ïX����߸��g�Q7Dvd뱬���M8�uJu՚}���r�n88������`��5����'���vu:�YY*A}��ݜd�%B��<��{�q�XVם���}�P<����$OY++�������
~מ�2��%�e)�:�Ԭ;���p���>�K_~���Xr�?��
�k��nV�{�)L"�y�b��r>kye/.� �/:�U#1��8���o�q�5�B�����g?�!m!Z������ i �+*y����:�Y��Dv���V~X0���V�q�J�Ϻk�ja\�֝k��0�]��p4�R���72z2���{���~����=H)��_���n�m!m����w�`V����k��u�1п�� ���dK���������;�
?#����_o�y���hT�
$�=����a��aRX�~���:���Ϻ�;�Y1���Wۭ��8�@�g�L��Y�7��X~�����z��H[@��߼��/�B�s�M��B�DS����Rp@�P+,N�߽�:Ό��d�w��CG��?+����*�H�^{�nmq�'m��^p�D\v{qJ8��m;��)�ʁ��/��P�̌��o�#�O/fl>a�������w2u��P,<���p�D�>?�_��<���H.��p<7H)�}�=�p����Yނ(J�!�*�E�������'�|G�Do��F���b���!Rmu��TD�Vw~}�!�aXV%O<���H,�VL��}����{?:�����m�z��[�%�e)�8��Jü���^�+R�=����� �>�w��W�1�6~�^��0PQ
�Ջ[���V���Q����CPe^ǝ��[�)s��\�n?+�j��y���$ ���@�D
�@�?������J�P�<�����tIXS�ŌD0��8$��?��U���o���~�{|�ID+}���βXʁR�}翾���X��k�W�?{k��������R�_~���p�����K��2�.��:����y���
��YFJ���ݜ��C�o�}���f�&!D��>�;�!Ԃñ�IS�?}�Τ�B�VVJ��~结����|9��:mY"�D�QR6_�$��]�׎h⎷U�M۷���#[�o��������.����J����͇^�+R�����9Ф-)
������}�"� "<��{i�uw�����}߫��?J��P�{���l�Aa��~���q3Yn����R���wI=*G���{��3��������%��J�O<��u �Z�~ﻁ��)�z�z��߇�L��a�����A17 ��Z���~��l�v VVJ��_o��g#&Щ*IX'�7�M�����߽��x�Xz¤���}��:!Y,ed����=� s��{�+tĹ��3�HG��}@k���d^���
#�H������*Ah������ i ��c�:�~��a�¿���]bJ���:D�0���V�+�|�jǝrKe{U��������gc��(�օ�WY�������p����'�*�@b�}�|>�}�3�d���}��;Vl��*a\���!��+��~�q��T*J�?^�:����ܮ�שgwĀ!������֤���w������}��ף����׏�gU�j���2 ]��c��'7E���[�AV�m�k�V#��H�g����Q��1!��a��uv��u��������{���H(T������:ì+�׹���k����y���Τ�H,�e|�y��i�G�yllְ�֋�@�V���n`t�~�չ���GgW$�:��O>�� ���=ϼ��4�@�P+,Oy���gY*AC������m�C3�����J��}n4�4�ծg!��+��l80�J�H,=������%e@�T?{���|1�������X`V��>�p8�R�w���z0+s7��II�!�E H�G��o�D�3�>�}��߿�x� ����82m
$�Q%ag��＇R�*����8����9�v��d���FW�|����@��?=�D��aL�ԂÛ�߶�`PjB������)�Mo��g3W�ސĂ�s�I��@�;�?{�q ����b���l�Aa��^}my �o�U���^����u]�����[���[�k�{�A�a�[Y��[��<iJ�Pڽ��͘��)s��m
sp���<���}_W��Y�]���{�W0��Z�,�]�� b����>;rr��z�Q�[v��Nl����Ӟ�uj�R�� ��8�<+G6غ�s����S�;7Z.��v�';Y�Nh+`{�������W�X�qĚ8��r#2�B���펷]���7��=�(ɨ|�v�R����s�q�k�7�Q����;�r�z�^-�<\	�	��@oh�6��=�ˎ-�V���ѫ��� �s(�u�=�]<ь��5�5Z�?~p���Lѭ��Am��l?���T*J�a���p�'FT !���c�_Csӯ�����4�/��p9�A�!l������ױ�[�w��0�sE�fa�<���_���:�@�������{��I�Z��i�J�IX^����a�¤}���8����VNf���7��漝y{�wH��j&�k35�8)��~�v�X5!e�~���l�AH)�n��\�{����>��O*X�YD�~��p�:�YFJ���~�gRϵ�}���(��&_���iGȎ���¿�g���|�$�B����{���:�YP*T
~���p�R�k���w �p���r��o����>	/�V{��Ç�j~�A
���W�,����u��� ��>�g�h{�߿e���I�x$�/�����°�¤�?}��l�N�+%Y(��|���țD���뵞���j<�1 ��	�
� Q������1Բ����Xͦ�dqr�q�v������٫�Lu�)~=@�+������Z��h���q ��+X������/� Duz��EUw��x��|Fo{����YFJ���~�g蒰��z��qk���Z�4Ì+�߻��0�JU{8�'s"�UOι���\`��\�ʭ�RJ4I���_>�,�vЧ]��J���L�G�F�>T�`)~Kݛ�|���H �7�<�g�βVT
�������u+��Z�|����A���ϋ��u߿S^����n��Uy�ͅ�8�K�#?՟�a��d��|�ݜ��B�%Bĕ�����?o���[��s��Aaх@��߾�ĝ�VJʐ_/�{�@�w��D�Mff�g�V���l;���oO���08Ԃ��}���$� ��y！���R��O7���g|��}�W��w�<���Lf�*!��϶u�+�?w�\�[���ra���I8�ID+w���d����������|y��
����:�ؕ�Z��~�{��st��Xw��p�с]���?{���Y��J���%�E���sIv�g�/t�8��&���v6m�g���w�������*�.k/���g�
��Yc%}�~�gM�RT*J��}�!Ԃ�8��kϳ���&�g�w͝H,�ed���|����6�g�z��*�k
^H	�]_�P�E���~��y�p���g?JB�B���~��4��,@G�FW�u�ٞG=���6���"�EϜ:�Ig�ڿ�?��R]�w3^,��d��`��x�l]�<r0��\;��z���ioqސ^κ���U��Z��U8x��c��R���x@_Ak��`��ܻ� ���%Y�� �S(�������үiAf鹵��_i}F��8�̮&�����q��y�we�_c8�dV���,�(�����b��� I����8�Y��5�&w����ƌ��ͭ�.����h�O��|EqD�����g��#Ϧ�ݼ�����}�J�*��.m�+|�q����D!��͞g�Ri^�T`nt�ݟl�ǡ-њ�����˞qR�/�y���q�5�sk;6�����V2���^���s�(�ՠ�B款�̹-s��_s����˔%0UJhp�|P2�=�h|:l�/��
�Ӄ�pTL=˺�P�Ws�:��>�S0`/�9��;I�o2�^�b7N�|a�ٻa,Gpv)�.�I4yf�n�����,s�y�-�"a�IR6��X�4ޚn�^Wh8�5�+�L��;��c <�_���S�>WB���p�U�R�ɩJP�,&��B|F�g"w�Nk�sFڎ��"��;��X�+]A�/;"Vi�uo�=޾ٷD��ŐK�w�`��3k7�9Lһƴ:BT�4&5��y��;�םVb�2�����־�R`9�x�M�D=ʔ	���|غeQ�U.�V�R��s%�WFh�����I�t_XǪ���=�V4�|_M����.���8ȳZst'���Iꋕ[/N�w�Z
�dqY���p�]V"���E�����V��h�mj�YJ���J�&-ưs[j�J�d�.d0�j��m��c-K�ƳC(��5���jRTQ��a.����q���-��5������ ��ʽ���9\/8���rU��09��=�����
ffF����R�[���1�ƹRᘦ��3+�ĩ��1W--KiR�r�6�9�Z����g���n��)�퓅���`�8�ۜ'.9ȹ��.aLs+���m�)R���2�\h�#1*����8�M��M����;q�an	��0L�kp�m-��Lp'v�;���p8�@7�"4�ceZ,TkE��j��㱶��&��ɰr��9�i��Z���ZW*�j��k2�j�c�h%�UQVՖ�+*ڣZ�ҍ����E-[-T��V�lm�pLZ	e��Z	Zŭ*��Z�ek(�iE�Z�ƭ�J��D�KJ�F#A�YkV�d�-)H�X
R�����S��I��|���|粄����d�W��F'q6 �/{n���v�!2AGz�A=����{�8��]�gg;�e��}A���>���"6�P;��� �{��V|��!��;ʬ�"�y�$�/ջb��wz�����\ڼ��tTh���M�QŃ+�ݱ�v�]d�[%ָ�d�7Z+1��J͸�~��ȴP'-��+|$���ݟ�������8�YBy�����|wg��}��)�*4+�޻ ��>���GnW5�!u�onPS��@};�� I��b��$��z�kŢa�!+U�ZI�{�VH$��uح�T�)n�'������P����p2�s���(�r$���q�>�\a?R������$k�K�ң�:l�Rv�{�ï�`6���i��9 �s7b�����|,�����%�cuG��6�*�n��Ϻ�t���� 7�~�w~� �Uz��18���_�Vݓ�?9{BP��ޗ���JwD���b�{����×�':�B��<n�h�$�A �rH[e7����l��4X�C�\�����י���}����ܑ-�#nA�=���dww��$�9|�#ǵUxD����{��vOÜ���(���ܡ[�����=�n竾��wz���_T�k��ת
$�~���Ύ("MHQ��;ՠ�v� ��m���u��>�����F��}XkAaB�D7`��]�T���W��ω ���B���tg��<3>��G��Ϊ�rHo���2�s���Gk΀$�ݻ�|=�`\JS˒�
]�C�����k�omj�
w��Ne�RW��u�]:��Lh�ӘT�ps�/o�2�`���F�q~�;���/r4�i <��8y��$ Ǿ�b��tf%t�Z�L+n|��f����ۑ{=�<:�qk�E�k�B������Xz�R�77fzvv�cp�>�����ѫ�9^Nt%�"�D��u���;�wZ:ײ���85��c��a�r=�xMFMyy���&�xz�B��-og��k�tl���R�ev�rnn}s�n^^��SHn3�1g{[Gf7�q`�{;��r��6�0�-q�Ff�]��ut\u�ۂ����n��[s�����Z�G���~mD�E�Ђ_�ݭ�$��ͨA ����������d�t���� ��YΌ�1��dH��
����œ<Ě������֐A:�9����ݒ_Y=�.�s��·\�hذp�u�n�=�B<�_!@P�{�\�gg'��vI'�f��==�d���G���Сһ�Y��-l�}č9ޡ�7j�9��\ΙF�{%$=:�V���"�4n���u�,�{��G{#��ǽ��=Ӷ�I����5��w���fH�����(Ȓ1�1���ڞ� �G8�.�z�On�q�f�|��?9����`��e�BI�M۲	'���]�9o�ZA�/���$v�۰	W��Q'��c+��lHT��/�)n95��_�w<$0g]Z��6����nb1Ts����d�O^Vҗ�2u_;�޸s�����.;�|��I!mߛυSO�w�'=�����f�4:eA�ɿB�c	�ȑ9�on�$�wz��@#%J��\ft{��7lX';��d�}�	���$�&[Q����3}&�}W��� '��P@Pc_[�J͸TĲ����ud���lȌ-�Q�]+�vI'M>�W�m�V������PI�䀠>k��2���.���������YC��շB=Y�f�<t��ˎu�q���v��u��� �@��7w��dA��z��I�Y΁=L/W�o�W���vI#���Xv�} ��(���o���k�*�u����	gT�܏�i�m�Wwj�_�Q'q�`�az{n�q��	?�Ȝ�;4M�ҍ+���.2��/qz�S�lӻW�u�
�KWZ]���|3�'S)V�-k��.���nk�终#���ߕ�֝_�&{�������7���`�p����p�-�"r(��{/�5v{�����
5�T��^� zg�~AU��ة�^I5E�.��	6�=��A��_#!���e*����ͨ=��W�]��W+E��'QU����lKI���J�[m�)֤�؋�����	{}�9��*4=�����:c�� }鞉|=�"XX��%M��PL�}:�",P�^�߈�W��m��*�ծoP�T8��P���b�)��7leU��K�$M>��l���H$u�FoT ��M�~$����7޵Y�'�I�3��	#�{n�'��ͨ����0K���U��q �>$j��
��ľ�>��y8&׳�ߖ5��o'~��ؠ~�_�v��wa)�՝q��wc�M�F��LS�\�r�|P��l��~��.��ޢ�`��ni�湽s�H���ݚG_��p�a����ߤ���.��N���NzۯS.+߅��T 5��V�w�Ұz���|��s�������`9�=q�4���<���u�[���
L{�x�*Ti�"2��ٔ! ��3�,�O����vЖ2x;����N�ƥz�=�6����0��ЮڿX�Q�YV���y�+��� ^�۲��zŚ�%�7e�(o9tq��#"	,]��޻$��{�d�G��p7*g�,�ެڿ�/}����l���H$tB���<��=�xϵK���>��y* 
7���|�t���|uu��>~w<��f�)HR��:����jb{��V	;�ޡ`���_ms^3^�C�k��"�@/U���Ѻ���W�ő]����r���{�+!:˓b7rC��wQu_�-�Ѷ��f���}���Ң���������>Xq��n���� �Clvۊv��ƃ�����839)���H�Ӵnɝ�A:�]��)��m���@�.�Δ8uD
pjܯ�j+�љ�ouÇ�<�mڻ7+��H�.�v�����ntu������<�rv��b����5�<�h�-=q�ns��ֹW���um�l�Ar\�����B>ێ��.=u�Xn,��s�� qK�7!m�n�r^K�n����ƫ"<u��	�n܎����k���SY_�zH�����j(T]3D�藀WS��`�v{�d���t�YQ��iK�=ג�Q��[8�9�����Gv{�I}�@�{��y~��I]�Ħ��rH��/,����PM�ETC�f緜��[��۝�$m���\J D2X�5u����g�5@��<O�V�U�OĂO�v}_{�=m�����Hy���+����1���pC��!N���Y��}�=`�A�z���>#/�B�#�Y�M��߉(�TK�(i (��.78�����3˘�{3vNl�=#����}�����r���^�2kK�>�\�� P5�*��~�p�����f<���$G�v�����[M�O�ݙZh�eo��ԢϽ��M�����L�εA�8��7���(�)���/.ͬ��X5o%h��]fLQ.c��dN�\n��\�.�K������τc�����w}�|Q˞<����ɢ���t.�	�_
�7�Z(����T�}��}���� TO����g��)�sI�B�
�u����&��	"Vz�O��3fz�	���������V��{.��\(BD2X�*oW��v����G>��q��$Ft�]�O�������/ז/5��������F�K�u�j��S�l!�½y������q��]M����p�94�.`�|rd� �L�I$o{�v
�C�}�Z�� c� �;��g.�P'+���*}��A�:� I��| ;��
�W��Z�}��LL���耶�����sl$w{�VAO!�76��1�Q9���ʷ��N~y0^��өq÷�:X�Qd�о���M��c�2�0z<��^��V{^-2����}�������?|O����ݒH�~�]�;��T���"j�
o���ld�1rQ���,�	����A�ʇKə_{)�D̻˲[~��!1':z��A���z��|��<���ys���)��䨒@#2����%{x{H]- ���eu�`ۭ��2[�m�{y�q]������m�Ꝼ���7�H��K%L� �s��VI)��߂%rY�s�����%@���M$��$�[]TO�9����˛/E�I��]�H'�3+���;N&7�W^z�����S��.�f���޻����(�Ee-���wC��{����]_Q W��i�$B}����{ۓ�b�힞����]'�Aܭ�@�y��tG<8��6��!3jn�{�9����^'p8t�e:*z��OM�B���=K����렩�U�j�+վ0�:W���R�sf������*�����n423$�˲?^�l��,��N�'���,��k=]vH�3+��	��v���ד7���P�TD�:�H�t��w\�m%�w$�4pL��F��U�v|/o]���a�"

q��w�A ���@���=__��IJ.�5��� 
�]�T`���"	,]�W^���gǐ��t��=~���/ҁ �d���H5�+�������^��{�|��Zi$\�$��[^���}�v��N�"������u\I�2���I���q�J8�G+5���3$����J�nM |N�m� �}U\�l|}'�Cs��{�TG(-h���dI��=�Ϳ��H=��U�=��xҡ�x�{�WĂw'��N{��K|��n�O_F��WIU�r=��+�6d��]*����ݛ֜��ۊ�_:b̦l���]nL�����ʾ�G��u{6Ӵ�h �@����]��:V��2���O#��X���ⷶ�fY���CM�[(�<��;o^�	ن�+��g	Y��U�(�`]������,e�K�}��V�<�]�l5[]S�C�� ��7��sR��y
�:����c�+��R ��a�g�|��ǂ��V�+rI6�i�p�G/���!n�L���5�c(�T��D���-][2�t�L�ʵ�C��û����&e����W/��p��ʰj��]�F�Y�ʬmʳ.T��tԌ��5����|�T��j�mJ��`sgi��#ZI��>̺�Z�*�St��et�rZ�2������)�q.�%����k�����M�����xm%3*����o����0�\��,�����qi̻�FoD^z�Q�jd�=5Ϫ.��7�{�,\B�f5�����wo:�ɚ���Qh��mf�݋�|73���G�����j5�h�a��q����$��떸�őf��WK��f�����xY�BCY�_K��juQ�sk�V2a#��ρ������偺�V ͨ�X���u,M�卥�f±mL�B�=��8��TF��P�2�`�8�s��2�o���#��)Y��'>�K�ogduT���2��-�[Z��=QBv�
P��9gy+�^��q�:��.�J��V7���ze���boU����w����r`Æ�m���Q���4+imJR�j"6�[j�)Z�2�V��Tj4�l�ciERձU�Z�4��jU�m��TF�+V�k(�X�(�h�klm��FJ�]&e�6��J-k*
,P��UT*�U��QE(�KJ���Ae�Ve���&��MZ������)m�֔[�.e�,V����U�*VVҵ
U)V6Դ��(6�[[���1�m*�[F4�6�,�(������)[�JVUEkm�*�J�("�l���X�u�LHV�����JYal��e���+m�-u��3�Q�Uq��1�J��mTU���)m
�QVVW3"�+mE\s)�f-U��E[j�%���mhZUiE�L���-�Kj��(ҕT�mb�(�E�+YF���j)B��-�������j�V��,J�*�KE�(ł(�bQ�m���T�(���Z66���Z�V���ZYDl[M2��(��jЭ��AF�V�ն�P����k�un��/l���6o5Խs��U������gu�n6%M����f�V�۠Nt����`�f���q��{]��=�4�[S�mڤ�qx�*�`N��w �	vcn�m�,����n�Mǳ��6ݟN�W[s�	����Uԡϣ�V.#%�8�Ѹ6�j�Ո����N%|�nC��q];:��7g� �=vwV�t�l��fk�V7)֛�7-�{v�~s�v�Up���aZQ���xM�uq�N]>L㛎��^���.���ݜ;ڸɝ�nzv���p�[Wm�كj�=-�\��݌������Ӯܝ�,]!�M�0��<���`�9��糫��J��ļ�Oa�3��meL��^���s9�C��˭��c��I�wl8��>[|���:�N=Yng�y�|�o��lm���v]7m�R�k�ݛPɇ��;��Żu\#�TΞb�$�u�ز��� �Y���h�:1�)gX��X;h�XD�I�&z�V�7vl��;u�Tq���m�3��^����ݵ�5�'.��3u��t�m>���[�D��Y<�=��z�Z�r��knv�guu;=���)�6G�y����#�ۜ�ŶE��GbW���cX��r�+v8��;�C�I�#��l�3`w���.{�[,U�Z)�ў�%��=�Żv�Hl|�w˃��v�1�`zpY�����;{n��-	���8�Sӥ)�on簑�ov�㱒�nF���=Z:�����m]�5����Y�㶳ǅy6�����v7n+vgY��k��ۦ��k�v�۞�b�[�d�\s�����ݝ��%���F�e�x�͞Wtrk�C-"�둎p���'�n�5�ɍɖv��G*n4�>oZ.�U�y�Sr�q]�Ln���6�ĶЛs��ó�P��}�}м�krks۱�v�s�]���΋q;�9�v��[l%��}*��U|����۝/͞y�ne����KMذ���(n�B�zΣs�0�N�ӘkH�IC.]&e��1�hp�C�Ye0�r�[��2�yC���O���ۉb���v�]=�s�t�M��͝L'<����E׹�ݝ�p�e�V�u�ڸ{8cv�=�/<���v9ŋ�A�,��b�n���|���Y軩���%=s1X���7W�xR�u�sQ=,l��0ro]v�m=^�y�;1���xE[�������7�5=pmn��@��.A4=�6��'���C�7	��C�����7Vύt]�C���K����ѠɆ	W��̡Dsg�ŐH'��<�x��n�w%�����^y"D���2FP�B�hW������͞�����Ղ�$臨��N{��dD��GF��̘/k����d�"	,]�j��vA ��U�@",�t����6m{'�H��U:{UP,K�`ݒE���!M�V�.�	�D�9�vIWN�K� ��vw��un������\�!%&%���	 ��ڧw;;3=�����4� S�J��O�v;��ގ�u�$�H4�-%N3"0>�M{,9�\�3��+8.�ּ�ʼN�������v!o�"�޼��;:����(���^�Ĥ2g�œ۝���� �@�!Û��I��w�dʹ�ڽ^��V�!~�u�j�KA
�}���Uz��,0xRb�A�|�(y����Z��CV�i��wo����sݟ�w��Ծ� 0�mg�g!��=b�W�J?����[2BВD�hP��e�ĂA�y��x{�y{��=�����z�	8o:�!��.����Ibĩ�yZ����U꿉�9^y�Ē;����Λ+O]�p��'�;�v!a��H��I@�7�$��v�efzWN�L'|�� T	˭���;k^7��y�ގ��b����C�F٧�m�0U���b�n�s�1��('�QB#�;�ڂ�U*�O�C���� 	��vg:�.���y >#M睙Ix@\M��0����6ŐWݼN��Q��9��KU (W�r���'g����v�ؽ���C�Ց&A	y�x���7�BM�H| �_U�(�Ed�T��J^��r�ueoٯz�qG�k���b�;��M(�{n���Q]	����35X�{]w".�r��^s<�s[��Y|�����>Q���_@I�o���/����9BHbr!]]�WPg��t{*�~>5y@@A?f�ľ����rX�G)� B)���{L�$�0�Ib���u�';{�7.rfp�Ӝ��Xq�뭪�z$ r{ھG�����X^�XLz@ӄ%)!v���K��k�p)Ʋ���q:;!���8ٻ_����?�P0Ϡ�]ߠ?unز��z����y�j ���@~$fWm�5X��(JBJ7X��^K�B�`wgxN�X ���S���ѣ���ܞq�(^���v��ݻ�P��iΒ�`�`�S�A̼�_�f�z���/d. D�9���ͯh�WY�A��]���ozőǳm.Tb�W{	���"�P��d��uZyn�oU�X�fiw�.�<�r�AQ�������p�>-+�f���à��wi���@t�[���}��p�M绮�$Fvx�"h9ND+�W~˿�$���k�q�ĩ��!?w�4���� 
9�α��)/nx�[��߿����O�LY���ju�\-ՖŲ<sWWa�/�SX�]GJ�<���m�t������@ �;ڨ��*���s3��A�|���A?{��vWl�M��s��g��C�KqcG����� ���X'�A�ٵ>��Q�W��(;ͽ�jg�ƠE'%1.��^����mBI^�qP�F�z�9� ���%@| ��7�FZ\ .&��Ƞ��_�O�s������P����E��+�|���(C@��uY#��"A�˳�]6� "��(���TѾ�q�����?f���z������J+���2����mY�)ڥ�.�W�.�̻�Z����=�n��ue�4��	���zg<�vF�mzt��#S� ���LW;GXe.V�f��oNL���n�ܼc�e�kvv��Ӗ��s�N��m�֗h�8���Ӳc����;M���ޖ��9�\�к�m��^וX��F۰=�n|�l�p���p�:��r6��m=����+fz;�Y��r��`'�9u�H�[�k$v��)4m�q�pskoc{a'��qr��.m��z��O99�h\�ƈ���3K�Q�j�'��Q�ں�m��\��
�v.~�w��ܶ��د�^�H� *9{@�^~U�vحA}6��>=�P�c�������{�������S^��$��f�$�g��'�o�^-����sA?-=ěI$��'(���=~ͻ ��V�n>W�~��I�[�P'/����9�j[q�S�uUjw.�G�n�O~!�ΨA?�_��$f�z�d>j��#��U�ZX .7!�8�{��b�'����Y���&���@R;�u�}�ג�)�w�
�)�y��,T^ʽ�z�?�`P�H'v�tc�kR�������=�}O[��z��7n�7���ޅ��F�r��׮� ���ő� ���볓"�M�g�Q�z� �n_�_ѝ�-�EhP��m��y穝~���7���C3ٴ��3��K�a�˫ۨ�{�"�upV郪s����7;�kH�˼���v�où�Q�e=ڝ+
�+���| g�߄$�����
��ߒ�(?uq�8p�]���v� ��t�J?$>����mD�W�QPߝم�J�@};\H �w�Q+N�q$�IHD	���9,�Y��X��8���
�wyR�ϱ�a��+��weY"�y�jZq�[�)���`xl��^�l�X��7r���|�����| ���Ek�\�h��t� rɎ7!�;��2�ԝn�e\:�YC���ғ�m���f���9����H���V$�����g.P��˰	�޻���^�\@�
�.�>={Bko3�g��~��$o��H:k�Po���j�!��W�32��-�O⌉!���w��/��g��
 9֏��^��:�>ܛ�j�݀��sÙ����"7�bcپ�S�C�sy]�5mZ�8�������q�X[��.�*O�W�W�{} =�߼�	L�����z��`�X��vn�|8&�il���M���dH�7] H$\�z��+3AVpX'�Y�]���>��I�����3���N�f��<�1��ր+5��P�l߲��-���]����9B	X��*�E@
�]���Xϝ�"�z&�����H��������-�e�Ux�O������g.�a���^���	����WH�@d�G>9y[BOH�C��N�=�`�=�  >g�/E�~_{�F}�>��[�R������Ы�r�_{#�h�T���B�OU	���Vǫ*�I�����	��z�����8�"HcN1@w�z�~��x������8�[U�A���	�����=+����UYw7n�eMWZ�l�{mg;�Ҟ�u_�.�Y�ޅ]������e��^�N���ĉ+$3���U�H�Pf���ߴy�ƋLN\9ς�=��>w�jz���������\7=�b�;��W�镗����n��fy>�x�t�e�7k�:�\�9��끍��{΢,%�� �hǮ�?7���0�&6��}�Wm�A ��ڰOč�{�g�U�4!��r�nf�7���K��ؕ�w��T�i������~�(񹻵t S��%@P��'�㗔�G̬'DIs����۳� ��ޫ$P%/ϼs=QoN���7�Ń��z�����3P�V����������|w�R
?{�T��Sk�E�h3�����]wP��٥8�"HcN1^�� Q�c����:�Arq*� ��{��!G�o������5�q��?y
iv1��4m�/�
6��&���%<���v�����P*�,�m��Â�Q=�gG;U�U�W����^�7���w9W�`ԭ�a�����;=��ri���Y��۷f�y5������^[����j�[m���d�ϑ�ϴ�]��������ƞ��Hl&w9�v�v�[����nՇ�N�ɯn�t�E�%��t)�nyp���v�l�h�\V2��:(}Kq���`����9ѻm��ݱ�c��/�ݶ���ط<,ci�k/7�=W\r�8���.�00z�ƶg�j����ۊ�)�Lц�r�U�~���Ʊ��F�������98�H9���������&}��������d�H�{޻ ��c��,%$H��[^��B{�CtʲV_)T� t�y/� Ve��璩�Vߞ�~�x��zu d�-�v�]� �;/hQ$��^
��t~ʺ�|<	����Af_���t��(��8(�{4bt��i�A�[B��׳@���Kw�5�/�[�tW�K�H����f#"N���B�$s�|�Xx���h�y�)E�� ����hQ��mY�s��uo-�c!,Ƒ�8��i�9Ӻ�U�s���3��N5�5���cʛu���{�p�D�Ɯc�&z�Y ��� ;��T+f��r���R�sstM�����n�7W�d����.�7���糒O�zs�����0�U$�`��[c�U���ʪ�x.��G���J�w�0}�t�a��������r���	#s:Q ���g���WK���7��$/)�XJH��� ���@|%�M_Cϼ��/��/{ޡ@Wfm
���7�cQL�ؕ��^��x���:���$-�A@5��v�����藩��9=�*6�e���GgfزH=��P�wvK>����2x�_d���H���z��8N0���󇶼��V��/;��5ӧ�3N�exh�����,�!)��n�W�!��D���}v���n- ��9an�N9�{�l��6�̃�6�����+����R�����9�@��g���� -�ݻ������^ A~�{��2^�z��~�𴁡=�A�L�DM�
����$���z��%�J�ϻÉ$zs^�n��>�R�㭠\�����MB�-���u|U�m&-fV9J=H�X��;���0[�¥ŕʝܔ+��n�'왽��_R��La̢��/�{V��xv�r�F�p�C��O���i�.�1+�;-sM]��{&��:�*S��/�\y�5����NnU�P�WF�쫊㮈]gS��GnWWNYW�Rэ��|a��mvEeSԝb����e���ְ�Y�w��Rɓ�c5rƵ�փ�v���2�rT��6�0n��u?�5�H!�i�p�.�R⼻�kp�E|�o�Ӱ-����x�Y����n��z��t�.�9�Vt�i��]8�*��(b����Q}Vn�f(�0�Y���Fv����e�됡5�jƴv^T�K��n�t납��V<��������Bc<E�v�ηv��N:�jK�oEZ\v���!���F>(+�T��h��P��䴩Z[Uw�eA�G���̏R"\�*�;.�n�.���:��.��#5%:�\���J�b;K7��w�l��%�Ѫ�>\+�eN����G�Qk�����0p��H�s�{[����'7�#�쾾���nI&��D��qu��L媼�O#B`�� ƨ�)|w�}�{��Y���S�6��˭X�5���&��S2`�Ù��Cx���lwl��SÎm�X��5��@�A؆�"�(�2*�.��h�[ֲ�d�GdZ�r��S�	c��:읚����1.��x+J�34M�k.p1�5G,�/w�[̺+M����3��r��[�~y�����TeT��r�6Յ4b��(��G)J�-�5�V�Ҵ��mKiZ[Km�U��QD��l�)*Z��KKR�-��[kiE��%[J��XQ��-*T�pmDJ6�Z�lU��Z���kh�b"�V�iU�J�[[(�ekX*[bV��AV�U�-���cs1�J�Tb�#m��Y�\YAZR�F�,m�6�%������ѵUUZ�Z�K1TkDYRѭ)Yh�j��MՖ:h6��jb��)A�Q��D2�J����
�U-l*�Z2��U����R�T-Q��\1��F�\r��-���QP��D�F"�JU*��mV��ʊ:�Qq.U���1��-b�R)���U�ED�j�F�kUm�����-����R��+[m�(T�%F�mkh��(���q.R�(�FҢ[E�l�Z�Z���j�1�6"�(�"�h%����0X��Y��G)im��
R�U%V����use[h�*ţPӬ3@�j�\M&[�Z~_/���y���չ���@##w�~	�®"PUE)~h�t�<��	�vη�� ?fk�`��h"!c��V��wW�8>W=ۻ��n�S$�UP�eP�1���D	��Ǔ����/����ۻ� ��o�/�Wk�~��˛6�@�$���Q�3i��;RvYy�0/CG�k��R�q���;7���xx@T��1���w�{3)/��%�H�m�(q�* ���[Sxz��f���mx6l�jhP�&�
%6�.�cM�*�C�moL��]e��@�w:�`!c�m&@��e�X8��y�̞N�d�2�5#�k�W���_$��6πͯ�ku�γu��߈ >�����?E�LC#����P>ؤ� Tw?5� ������n�j�?*���]�:gi�gf��+��]C$�T7�
�}�l�!�J�������Kn�ӭp˖D1d�;I��7���}I~$x{�դҜ����%R��C����>��~��2����B���}�b�I"�I��=��v�õ=u*�쇂�j4�v�=l�j�[��y9�륯fև�ckE<�� ����R6�2Db+�ɜ����H��RG�I&oO6ɚ��J,{���<��e�U ��Ԩ��M�n�m��6����W���� F>���g7`�~�0Q�7��]6dښ1DM���i�����ńE�:@��J����7�Q��y��k�ل��t��r(Ԏͅ�=v��b��w�v<8�5����5D��ӛ$�H���z�;��o�T��y<(��\�m��*��HS�MH�T8c�ͻ�� ����oۻ��=;~��79��g�9� dn�~=�ĩ8�鹪�G�=�XgE�᧥��ͥ���ֳ�`�	�q�����7�6re�ڴ�J.|��C����з���V)+u�+!�r9��u�����~�}�ô�G���vԫO�Ѥ^:�w�ˮ�٬��\G;��nN)�X�,�,���q��oF�p�\�zz��ny;r<�eOX-Խ��X��(��nQ.u�i��s�d�܆�nʙ�ey6�dK<s;�͢Ν�n����:I{u�k��R�%�t3��Ş��G�.��t:���b-���1�v�63�C��ܯa ����X�!���-=�����1v�Y/; -�1���+�c��^��$��>��Ep�`[_�B�v��@|��w���f���cױSgfQ����l�H:��`�9�he��:{�T6�sŸ��=��Ā�7ٜ�E��i�� �Uߺbu������G�Y�0FYkU ��SJM&��۷j�����As�8�ȏU�u���'_uova$�徦|9����� ���٬����}T�� �w�ݥdDA�;�X	 �o��\����*���ė�M�2A��\4u�T�c�i�S��u�»�Y�@N�v�� F��|���<�_�I�I�U�I��E �"�H{:m�ɮ�Kl�P���5f�ṟ�U�F�Ҧ��￫�S�MH�TlG��_X 8������y���Q�{}�wf]� �r�]��ñ�Ep�`WV���Uo�W^�<��n!a</7Q���)����'ˢ���{�����_�߱wg-c�͕�%���l@��^�!� !�?[o
EM���}�����7���w���o���lP�ךw��$��`�#!�#@�"�Oʽl�H�ܪߒI�w���p��̞�t$��w�� �[�~��5��Tҩ�
���s��9��7(�&��VI��A�E� ����vl[iz�P�~�<RK	���D�x ��]�/� 	�ܝ�97��^�[ =��� �Z��D���6�4�����>�09�/.�3��v\C�K�[�ի)��9#��mu瓛]�
��w��DCr4dtO5:�"_$EE�HK�{�d�]�S�;�������q*��
~��Q��n�S����=2��{� ��{�"�{�	����҆f���y|U��� J	T�(�����ĀA���j�	�i�w������aC�4q�#V�)(��1t�ϡ���s���t��|VKӎp<���x.��G�X.�NfĲ�gJ���,v�������"PC��o�@�W�߶����2j���UH��P��{"���C��y�D)���� �]��' I�����&7�9�q��ВB���Z��RCGh]���	 ����Dd�弦�d�(�g�}�s� ���wh���r:鉨��R��lO/�L"Ltm���=�v�ֳS�@l���:I�;�z�o�ϧ��y}Z"*�߁o^6��v�� ����<�֭�Lق��o�@�W�v�� �}��"ی�����!��¦��؀�n���dCA��q!��*�fL��� �s����p����.HJ$�=���� |���� [�{wa$gt�Hz�jl@JI�!0]ZB�t�x��*�4^R�r���3�|���� +�c��<���~����&��U�W^��佛~]�Wo�wU;���p_N��>���R�v��
{TKY��뭖f��ѹ�v�m�_[
��t~�����}��oR��-�1_�'���$��ۻ�����UT7�K�]��$;�~�!���1�E�x�c�Y� ���#�F����'pE�'N�Y��&:1�&��c7=��s���&8(�gm���/����j@��/׏�":��_��[��� 7��R1����S?UB�U-�[���6���y�#afď}�� �_{�=j�D���ͺ$�>VfRk~������%��ɸ`E���6NtM$
�����A���'c\ӻ� ������I�ۣ`��1������.WY�۳����舆��j-D�_ysw��`�r�Iz�ċ��j�=�;7(	A*�R~y����$�\�5��з�����PD�~��� ����]z�r������3�)�7�)*2�i
K���һ(�K��h#����=�vhJ-oXb��F�Q�d�4��:�S��L0�9R''�N\��8�����{��������4Q��vc�������k�'I-�`��n;	vg\۱mv�$�p^2��¦�1�mG9�'��R�&�����ɞ�k�����C�bM����u�������Z�d�nյaZ�Z:����;���V�E�����p3����q;�����v���:����y�c\�A�[۫v��Q��]�����ӷ7a�l]�g]��s����� .yyq�^���Li�3wߗ� e3#@�"��O6��	 m����{w�7yz�s�U��a ]~��e�j�U�LpY�v����%���J��\k�}���H"���`$��n����tb��ə/R@y�D�l�� ���$~$�2o� �:wU� �N��ձ�ڽo�@�n� �T�x2��w�����y��� Ԥ 3M���� Fv�z��/���D���.� d>��.�XA�sl�k�g�٪���L�OzB@(��~` >��m�� �ަ�ފO24����2�m�B�$*&�\N��II�����'M�<]�����-�F<�������EjBL^�!s�Ua$����  v��0��;��2��{�{ϛd���	!w��HL��1���OJЀA�$�<x���R��S�U%�2�v�(�-�Ί�AЉ�d��X�iыG��p�h[\�����=���j��/�G����� ]�w�	�z�vS�1��MP?b�{��,���J��"f�h���qG�ޕ$�$�5��7i��S���ϒH�v��#3���f�]SSS�҈��5������{�cj?�4O=�H0��p�]v;��NDDj@{=�wa*��J�DHLҀ�4w[��$���K�/�o��Lt{�D�����w� nwSi+����=ʖ�ow��FUf�K-�+��r�z��n'���3�ۮ\�-m�8�7�߻��6�nƝ�ߨ~y��� 37���> ��~ �ݹ��y��˟s��$�$�f���.Z�Qa��$�tH��԰^wx�OU]�� �;��	
��!�>�N���]p99:$�4�̫�e�u�}�� �MvH�H &vp��u�+���Y��W��`5o�ҵ�o]g����b��kW�|�Hd�T����v�+@�>��0lt�c"&p����C��"?|��~��@�W]����&�H�N���ݖ.�s���twE �y��AE�c�H�=ݭ��:��-z��;�k�0����S��
�U^�/� �3_�6l���6S�s�ʫ�� +��� g����$����+8P��<�>d�d�m7h��Ռ�V�[O���^K�ƭ>�Z��lz�����$��B������%�  ,�ƛ����{���xO�y���=�v����Hd�	EAF���s$h�z�+���}�� ]f?0=~�L��N�p�㰧e�p�@���!��p�Q"�o��+亳�y�%�H%з���f[vb��չ�D0z��0%sNԈ2���cU�矬<f߇�5FDD���m���n�3��8+��?�H�ol�AH2�NP�*��)XoR�v��w����������W`�5��[r*��GAB���Z�r�b	��DL]f�3�9 �����^DR��A5$I���ŀ�=検U3ΰ�-�r��D���@_~z�6�FgOy�ܹBɜ�}�m�$J#�D��[���f�*覺y{J�#%�����мu�f)ي��LRM�.���@��v�> ��r�,)FO�-��etzH]UTN�Y�vNP��&�D"[���#��{>�,�]��#)f�{ր��$�I2yX�|���|�[r|���}�"C&*6������[�ޫ��m�r�%^̫�$�He{}�h"0�m*�$�J�S0L�(�O��݋��FK���PC�	w��� ��-| ��gDd�N��F�����?n�U�T�*U�M�a��mf?���kn�m����݀���d�I�ۣ_a���
��x�z��wvU�4�F��b9Fd����w�m�]Ja�u;�ɇ�\TE1��t/�%N�}Y#v�'S�5���[ەt8/�d<��$�;p�<9wb<��p�CEޱ��*���!��ҷ��N�G|Gn}��q0Tg9ڄ��F�qG������$u�I,h拧V�7�'wa
����ff��;I���MH�L�ݸ�E���)�c��!�׎���.+}.�p`?1ۯ�d��Lשnp��٤q
w�p�(��F�s�J�Fʫ�g)7v5`���.�R�,��1!�7윸��XI(�	ׄ�` �u�ǇNX��pػ��u� �u��&�V�s��;hvB�j$�<5PG�Ǉ�k�]��M|_��ѷ[km�;�@ƶ�ҫ(+`��8F�u�{�!{Oq�|Y�;"8u4v��ܷ㹁m>��Y�O��GUE�T4L[��.�m�QZ��J3^�xo�)��ȔL����v{6AA֖¹�.���#pd��f��ev�rp�J�d:UЁ��}[ żmu��e�a�βq�=t��b�7��	��mC:��1*�q+�].�	MT�̮�#�z]�k�[�3)��9��
�=|��|����ݩ/��gA�H淺���eoP���v#�{������.��6+���h�����x��98$�vrH,U.�����{;��p`�¦�o�!���S��-LgN��=|��[�P\�[�u���-����#V�j�T��Y��R �Z�҈/�2��LD�E0V
�*��Tk��1�iemJ��Q-�ŶԢ+m�ci�ain�L[Kh)mm�J�DYm�.� �������kQ4YEr�iT��EKJ�Z��Z�TĴlTK[kj[M4�FTkr�&%�j�.Tj%J-�J ڨ���#�M�cF�[A�����E��JQjTR�F#i\B���+Vʔ�j��Z��-���[)XZ2�Z��\�(���XԫQ�b��b�
���Q���CBU�B�Y+P[�U�V�ZEFV��#�Dn�-�+R�R��eH�Z!R�FѴ�X"��-t�V�kj���fZ��
V�c�DX�b�m
�j�cD
��jѴ��QʩKm�T�QR1U��j֢�+jԨ�+q��Z�YsT��f�*
մ�+JV5�m*
�`ĶԠ�*�)XV[ekm���TPƢ�QR�֊���q���l����G)Y��5�J[Yic�`�b( �SW�<�i*�3.4̹^�9�|v�۳��-���\kP���Q�W\O�\��݇g� /^819糎w/��&|v�j۶�Z}��P�v6ݶ�3�kv��<�FJ)�)�09��=�ƌ\�=d�)Z���1�8�}�j�����Mgq��i��V�\���*���u�cqW�)���a�#���JJ�[m������\,��a�OF�r>9�z��ۗ����c�m�hu�;-��m�q��3���v�3��>9�f�s6�����ڞ�v�q���3<��vO#nz��cur�Ɲ�[���m͎x�')��7.����es��x�8�n��:����X 1Ξ�BnӴk�v��طn��
�S������8������Α��"���i:8��x��۴c�C��Tg�qڌ����c�~c�;v{��s�p�k��a8|p���\���0t�2m�r�p����쉻p��:��;8�Lv}�Df]i�t�!��ф�*�h��o�/o�����pi��ۮ����I�nOn:�R�sn��[���dA$����;��/��۱�4qq�r<����>gt|��69����9}s��-	�c��u�7a��κ�{������=�^�<���۬���� �c��0q�����xpO���^,	�']�9û��F`p�y�s��[��u��^�:�K�\lt�ӏ;��yS�۠'��\�Ax� ۷X-�.�[��F#ƫv��bޝm�Dze^����F1�ݝ��n&C�	�N�\��-���v���J,�zݱiR�7pɰ�ָ8�{ct�[�vx���X��c<v��r�u����/=]'g��pG��m<�ۍ��.����ķh��͚7�P�n�S�.�v�rы/���ǭ�[�����㱶�1���$k�{Q������l�Y�\�0���5��R�)���vݹ�Nx̩�n��֎0;Uo6N����E��8���\��6;9��ꗑzy�͘=�۰4�V�UpNn�Զ����K��PS��7[<X�s#��F"	��Α�c�N�����vn2�/�Knq`�6�O2%��g��.�mӵ�PF�ۍ��\ �K+y��΃N��d��r[o.���8�c�ݪƚ�F�G���i���y��-�n��.�{I�e��s�v��x��]��NR���v�2��vɛ+��l4p�6�A��X�դ��N`:LS��p ֗b�� ����=H�N�Y��r���;46e�����`1��Q$���ov\DDu���@.��{C/�7�2����߳	ďj���_kŁ��A��Ciܼ7�W�kNc����s�}`�@,��r��
��""���j%wF�\O��jH1O�M3$�)\Gq~�%@���q Qkך��+f�S�׀ >7�����<�%G��	f"a!Af�׳����]�w;�v�L4.���,�v��;��jc� ��=XO� ����n�(���'[�&ς#}������.�feos�V���荮�nZ���d��u�4������.�P$ӉB�"}����U��[�8��w<�:�M��@v�@h�x����ڡTL���_Fcj��Vcl�{�n�"�}O�{�#Y|ڢ >53�$Ce�C/(�8n�+U����x�v6��\�#��k�74ټ��'T
�Vʳ�>�*�`0_�˃6��8�@�}�c�g�-�p��Q��4�
ݱ�?]�7W�I��7�Ϳ�	�D-�^q�N���sw2t�L��)
�S`�/l@ �gk���@ �\�.յ�e��	.��6A�]��%���qU./{�ڪ�wz0*��` /��w�	z��Sx&On�gI�Su%�&�玳	2�$8,���z1 �-�?U�N7�\���}^4I�rZ� �.�v 	�<ړf�z���҇��QT�J}�ٶƵ�<u�]�j�wn:.�8뎞v��+jV׬L�"&�V�Gl��	��D��u��`��]�` 3�����XD"[�rd���ݠ���A1E
6#�Ny����]y�w.*��
���7|s� ���ԑ�'ѝ�}�3p�2�������4�$�JM�ove݂�ܞ�@ �ê�����.��̮�YK�G����wP*{����]�@|�ղ�`AP���	ش�y�r�]EX*v�D�C����S^Q&9}3DKݻ�Suk�@?{�F� �3�y� �m̝1R�SD
jSaO���7^Kb�������&����$��=��M�<^��5���)�_����Ud�L�TB��" ��9�C ��o}5��ʛ�O`���ww��ܞmI�!M�6�n�*2&~��~�����{t�=��a���/]%�e�LA[x���h�])�1]����:WTҙ��Ǜ��V {=� D���=���k�\;�ٛ�I �����=��I2����){��/�˻���|�/Orޛ�w��D}\Ȉ��7��d����v�:o׺��uB�&(�Tʩm[<��D ��l���ͭ����ٝ� ��C� +���fb�&	�F����øg�Q�d�G�+ԒI$���I��f;؈��)����j�a�M��eI>��T�ω�����.U�/�j\4�*�m�
��K���V��zYP�.�w���7���A�|I�|�����̱�Vj��MJl�g��A���읞����t�
��u
���2�K�;n��:�u�o��dڰ��e��ш�IDx����M���;fz]�;Z8�
z��C�;?{������f��<r:6ׁ /��b�=����B����w��H����І�c �0��*�GR�4 ���/�<�G��z��K��mU��	/���-r�Nʪ�7מא:T�*i)��/�� A���j���&o·�]�vIs���%t�nf|���ꊄ)��Tʩl��sէ���^��em ���� Y�w`|����n�5H�.�]��HV�[L��E*&�J�)7�ٗX$�����=��'/��w�u�4 	]f�݀�F�_:�4UMĩ���}k�N�ו#kr��w7�:n^(�����A��b�����ب`�Z��|]m"���Φ�KC2����f��Et\A{�\����0����&�R%�z�v�ޢ��U=�S*�ڜ O�<�h�]C���mGk��Y'��w�=G0iWl���ۚ�ֽ]�@ݻc�k��g�k[�Xu�p/#�[���;�\���Z�wZ3�pV̲�O����4��l��[��pW;��T��z��3��
�3��nX�a*�� �s���<�n���O�u�ö	�<�������� ��āq�=�W���'Y�C>nM=f��fɶ�����_�g���4�~���g�$Y���ӯ�0�½�i*�!{}��� Y[�w`}0�qP�%��*ݯۻ�2��ŏ�P}^��H$�M��$��q�z��D��}ٯU���{�]55y�KQ$!!�q^�x� �2:��x>@ D�˖ta��@�=����D�骫I����"M�,]_���<DN�W�y� �������t� Ww�=�߸��_7Ϳ�4��fj�a�������%Z@?\�_%zr���@���7=�w`|dm�k�]޶���/��;�$J�����T("�unq���2�F�\�`LY��]*u�����?>���]DJ`�yw�w3(%���X��H�o��}�a+�fr��e�9�y��@|��U�<��D��$MJl��I� �ҧ=�S�?Xo�VLc�u�=�|F��'U�����/L�p��
d��*>n�5��ķ3CU��Iu�M����S��zk*�<:ڋ�� �|�> Ww�� �q��M�N�n�MFOAQ*�5@A��u��|�$�H^�6^M*��X���fl[�� ��o��]�i��W1P,�'H#�����m���$�K��/�m�?DD?��:�wy�L��k9%���C���)�e��W��slWg;�˿.�um��vZpTuߩ�� Ww�� :�:�æ=�����y�:7�sk��U��n�� ��ǖ�5׬n�N��]��n�]���k�������9��S*��W� ��M��ks�d��=��c�fѱJ��D�m�H���"�S���&��חvO������~�F]�� ��:�"�N籺O;��f�>=�u+i/�Tƞ�&"I�H������`2�9ݑ W׾p��I�D*7{�S0�T��*b����<j�����J�-��Z=ǫ:�J$��mdX�Tި����g]�ovK�{�T��ǀ�s~Ih�ݻ���$���FL���ƻ/Ѭ��O���B�z� @%}�ۻ�><:y8.W�{�憒+s��7��KP�(�f�Uu��Ē'Oo��e.�Q����rO���[� /��ݠ> ���ׅ?7��O�d�P�*"���mbu�rH�P�g�]�
�y\�<I�\y�������H�Q$�ĭ� O��� ��k�` lnw���^��:/���ߵ�� W�λ��V�%�B&��S5�Q����9Q���!⛫^�����@�ګH4H��+�sH�1�(ac"TR��ݷ�X�tvw���5 �{�pm��f�$�}�sl�H����/TƟ����M��G��6)/&q5wy�D<��iX��,79��Y}��:�Ϫ�CYe_��^I�6d�>s3�Uz>����]��7r�v�9,"�ګ�*������	&G��n/f;��}m�AJ�z	�TB��PJ�^5�wI|I�ڤ!���}uuD�Z��`2I���H ���UH�b]Zw�.�#
"(�j�|�DW�99d�
{f#�Ogƹ��W];����~���K[)�UZ�l�I��ہQ$�'8���]k0���˻ 679��Qt�X�mϛ7VB����IWT�2LuD�����<�A-;9��s�"Q=�Yt��Sۛ��{��T�+p(Bp�#p����b�$�nm�� ��i©�3���Ā@��� ͼm�C�mD�S���&���0���mmux"�Ho=ZI$���z!�9�u�q���]�[-��&1�t��Ɵ�������G��~�A$>F<�we��lSw���|���j�@˧����D���t���1T)�6�0_s��l�Zt�5��(��jo�����~����@y�n�v:��5ۗԺ�Q��b3��m�������6H	ۀ7Z9�Ģ��R�;���q��Yֹ9ln5���)�xy��WKks��8^Ά����;]��{sє�l�nI��9��rM�U�.͝i˼qWlF�t筢㎱l�{=��c�qc�5��w��clg]6C;�:�o�5q��vyM��T����|:u�P���.$^�{A��DW.-d�y֢�ô[��<T��4!mб�ط�u��e�U;��ٺ����]��~����v�m�?�um�lH ;o:���F����I���KH$��tqh_�yKP�D�f«��f%�C�a~8��~�  �3�� n�u݄GT\Yy�<�_I[��yb��x`�nk�~}�m� ך�DZ�=U�vfV���c�:�:�Ȉ>ͼ�f$��i��'B7��OW�#Ĳ�*�>��֛>�7/:�����{���N�S���@!ue���ǰ�f.��{7,�I�}ޫ�]G�_I���7� ����@ ��]� #w���u�l6��;�1(ߛs��Ot�q�|�hѤ�F^��՘�yНZ&P����'T�ąDԅJ|�cM���;� @a�Κt�;R�ȩ���6:�����ݠ>�]]�)D���o��\O�.TT]�U�^B���+�z���U�*��BK�j�M��5ީ�V7�8�:��|"�s@=�#�بmT7���������o�WΕ�i�&��� {y�v�@���PK�YڋMI�����I�G�%�����N<��v������ ���f���zy"{s��	%���R@�:0HYI6�͛�J�WO����\.[I��ɲ�`��q,s�o�o�t-��M�m�������*5*���2�����^7����Ѳ��Ҧ}i~�˻@ o����o�t��U5"��ѥQ�ː�i��b����S�yW[#�d�c�s7	�]��r_?�~��H��"TR�����qh�����@ ��n/���5Y�#l�Ǹ��Ua�x��q�cM�ca.7�b��s��a��s�" t�9�`x߈��{:�T~���<���0TjM�^Ҽ� �tKMQ$���S��+q���G��Q�˳��l�ҍ5�z��Z��nw�/t��>�o"AФ�b�����9��C5D	�^ �%Yċ��Rr�7�LgKXm�ڼr��5BD�c�̇�6`�a}�WN��0�a\]&B��A�a��+M���ԜAP.ƛ��a�;z`�I۷]7ը�t�t�f��l��,oڂu�W	|l�j�Ҷu�Ӕ��ۛ���C/v֖�
šS"��<4�Iѳ��Kz��ff���P۷�&j�}�ʵ��A���.��ʵ�Z9���&�+EuN�t�*��E�1L�C�wc$J٢�%��錸%���ݘ��
�;X��U��2iy�m,���4�o������!F�*�T�fN�P͚�fF���}�j����(>�uu��8Ɏ���fξ���j��``�7�E����F��%��:���^�ka�ݝ���QM��7P���B�2�W0F��4��E;bu�YC�������J��(�O2kx������F��a��t�. h�і���%Q��w���W���ͥ
��H�ͪ4
�Y���Uk:�{[�'C��'�fv;SUp+:-�BҾ���.|�r�ٙۗ�c�]|�x�嘪gEY�K�k,
����^m����Z��6�I�-l���}��>��=��@��	��yC���cʮg*d���L@�Q ���1˺Ε�L�Ǘ]��+q%8��Ge,�QGrU��h�k� e�����4��ʡx<>�|�\]뉏��+���3-�*,q̅��c�FԊ�t�j����F[TQ`�mhS-�Ʊj�[ej*���*V�T������V���kXc��b[Z��-U�V�kH����J��Ek,Q)j��Zت[,V���
�T�ҥ���kB���Qb��K,PE�UA�R��Z%m���Q�KT��ES.�VKJ���R��jT̸�b��ն���Ҳ��jTQb.�QUC[��1
��-J��V�F��цR�$q��f̶�Z�JQ�f5�3e-Z�[q���LB���.��t�X��R��X��32��������b�����\h���V��UU6�cb�2���kZѡʲ���JŢ�S-b����FE�Uc�����0��V..Yq�-
��)�Y���&:L���Jぎ��-R��e-�0j����s�z� ��q��q��
'�F*�� 0`�j�ٓ�z���㭧�'�g���@X�0 W϶��z�u����XNT��a��`e�ہ���%fw_�D����x$=f�U���iy�m�t�9h ��D0�}�v�&n��E[w>&����L�@�en������cG^�u�̜[��� ��<\�X�n������)�D�P�j��H�1����_- �I���ۢpK��h]u�;���y��� ����!���IJ�42����k��D�S�˸[�D���I ½*$��ͲM��y��[h�ss@���Ɵ���n#�|z�~ /���� �o�v�q�gd���` >:c~ H~�ۻ@)U��	�*'&����u�����]4 A�N��� ��ۻ��#/�Ly�ʬ��WX�3��b�Zz2q��j�E�}:�TeKu��&%�0Cn|/*��]�5�WwϦ��Z�_R�#q���0�$�뻤��Ap��gЖJ���I%���b����QV"�o�0>)�ݻ����?����Ws��J���m26@c!D�+�t�]�ڳ�d����.9�u�;�6�߿���4nAj�I��q~��| Ov��@i������A�<�i ���$�rݶ�p��G waC޻�H��&D϶}���~> ������ͯ5�[W��W��-x>����)R%E*N;:��� |���� �ڥ�Չߋ���X�#+7[���7��j�&y�JPMRm��mI��d���pYw���A%�w:h��a�%�օ��V;T��4�5~�h@���ɣ�x��ᴉә�E]�k}�E�I�F�`2MQ���� TXo��-ͳ͙b����i��9x(�"Kͧ��R���%4q�1�w�kox�AWzWQ�9[P�JU�Q�\7=٦P���ժƈ�#�nX,��/8�^	����u��u�QsA'��q�	��R9s��=�;%�,;3��n[p(E��{Cp
r�ʕ�����'X�>��ܼdV7�9�� ;e��s;���ju��㌾.�í�î�0v�}6�e6�"�Nob䋉���G'	��Fy�vX^Ϯ^<[=�ۣm�]��i�Aۛz��G�KvE�	ٳحr\ٶ}aޡz��;ecOqfbl���Vnu�z���iY���w[�N�[u�=�
�иBJ3�K&�__�"RZ}�UC@e�:ao0�+��{1+q���� >6;���ˈ���*e�Q(M��$	Z��	���n�k��ğ�{�X� �Xo�}��7yn?\5���x�ו��!	�a�@�£�]������Y�ֽ��H"���m/ p�^<��&���H��8��o�{��n� �Ww�� �Z;�Qu��u��M�:�� x���y&�(���*���m��I/\�uL�~��=7�v���\E�T���� ��u݂�������q �1�3$U$*�)�B&>'��d[�D��+q��m=x'�;b���?{+�Is���GC|߁ �!�z����n�_;5�r�&�P�p/ݻ���D$�b�XB
���� ?I*�<�r��w��;��"X�ːl��Yvp����r�E�������}���3i�i3���pz����|X�0>��]��f�Y������W�>�LDD�0�U���u�/�I.��H:$��<7�{˱��c�@&�X�RJ��ل���7�	�I�Tw������ޖEM���_4�| >}�v�@��>�~�zۢ u�~>��&�fiL�JEv�]� two�^3����D�6����t� '��`?��{��$ۃ��nС�~|?���.E��8'n��̌����R�3�J���9��H���ſ�@�e'PW���ږ�o9݂Aa����\�Ϊ+8���u3*�i_��vN`��� D�dٵ�w�I#-LCWd���� |��FF���i��\��G�=RA���BE�J6�+=�]~&�n ľy��J�W�弞�W�-���ј�� У*��2�#(m\>w}b��wO3�C=a�mu�u�#���ÝonGݍ�m����+� +��wh�27���TZ;	3蔂F����=�Ѷ��
����9�k�� @a�Θ#��zս"�;�1p�	!�~��	z�kpHQpSUH�o6ׁ�t<Ɵ��n�{ݯ� ��#o�I$��y- x/D�ҙ�'h�־H�V�N��`�~��@�V�8��Ϛ��:��}q�w��gq��Ͽ���p��ҟrGcܷ�two����c��#y�=��[�����$�L�X�&���q���ך�+L�~̺����~ ���M  6ck� �3AHW��ݛw�ʳ�L�AM(p��޶��$�� ^옷���W���x{ܖ�I4x/E��CdB�q�b6J��_mE�.��~�z6���@�\=�S@ >��{0���\����Enme�t��r�܁�ow����$)��K������.U�:��
�H��6�.�v��RP>�N�/���`� g�Nef]Zm�D�$�?rC�����\t��3-�CH.y��@�������-���o9�Uh�S$��|��ӻj����ǙZ�������NbGkmuۑ�/:v����JU0D��EL�Ǣ����1�I/����	vS�}S��}��0�U{�-y���n�&���13R�њ�-ņ��ۍ��>��Ǉ��� $�����D���� ���eH�nm���xt�[Рn�Q,���v� c�ɲ���vd�^����$�!k�o�@����ox�f���S*3��u[G�������|��������sn� ��v�K��({Rm+�^���]ՊH�CdB�q��2[η����������Vq��Q���� ��o�T�.z<-�f�gRѦ*�<U!�[ᕴ���Y?wi:^_wȍ%�����m��u=��*��:�N��.�u�{��7������etZ�-{k�.ն:��a���XCQ=�H{D:��;	��� #a�i-�Y�[v&�Q7m�&�T�.�+&�z5���^4��I�m��:Ɍ<�1��<n4��s��
ݷp���:�ɑ홹�8�6�^�\�c������i#D{,&6����맞��o9B��x�U��{O����	�)]�[��ֻ�ޜ%��yWlh�iu��F�:溍�N� �@a�Olι�Y��`_0{x��L� ��������|
��v� ,7��Aǩ���{7��I�&��A$�������j�2�p�eQ�ު�I$}�G/��L00�*Z~$�s�y�D�D�Q&X^���~^�_�ܤ��>e����
T�7z��Y�ݞk��ӽ��h�.[H��w�I{ӛ�h�ޗt���[�P7D�L�{4��E���������]�| lwg��I���.�k�֭+��� �puz�N��C�k�/no��m��^r랼�'='$�?8w�� /����񳓅���3��<��)E�!��Gov0n�9��a;buWQl��oCǉ�{s~~~��*" ���E�z�帿�27��x %��t�0�٧����B��j3f���@���VA�
)*���uV���R�����mt2��bo���.��`�y���&��&g]oH���MfJ�.M�ݽ��C�[���g��d�Tr�1�d��l�藩��{4q� {}}�{l,����s�`p�J��U��?D W�JP˚�Gvv� ������$�m_ԐWz��LfZh�.��ݹy}U�{�E��Cu�I�\WE� �:{�K�S�J��6���W:��)���M���Ɵ�����N|�J�/G�逐1���ۻ쎪șQ�΀�����
��XR�M�:��6��+/���Vsƍ�7f�߱��T����(�q�o�� ����I���vf%C�Z�~�I4�ױ��Lo�̨�@�EV筀tm�ǳ�g^��~=���� �)ŀ }=�%��X�(d��ϡ�w}I	̮��R�TK���� Ov�"�'^����f�Twϕݘ	L���e���%�ֽwO|Y��F��Z��6�X��ջ%�]'�T�+7 \k1DJ�Ki]\'�$�ͻ�P	>�rN�5Q��fd��0�R���%���ڝÐ�p�~'�lKOĚ$�s�Ͳ@&z'2�ϰ�q+�8�i�p�TQ0E*q}}oR�H��㭪�(η@/�退S}ݙ�t��V)t��-�HD�am�GY����q�v.kZ�۩<�dֲB����!�`QU�v&u2RJ)_ ���� 	��wa�Gu��<���".�6)�k���v���}�*i���*X�ϫI��R�B=���D������s���#c��D?��}�5�n��ղ˩��%Jg)$%$i�	��"I��e_ԒD��O/������Bb��� �F�u��{f�QIMUD�~��m\(��{!���w`�a�n��"��9=��{�3�y�v�h��n�.L���f:��fb�RWu9������.��������ovҽ��C9J�sLof�+A���W���wv����R")R�*A���X pj*[ؽ}��r�5$��D�O�Gu��A�����㦬����lyp
c���t�n,d�],��j����p�$��R�u���q��{�g�!!i��0K�^�컰Aѽ~~" ���A�'("����m�^{�v�@�߃*�&y2R%"�a�y���㽷�M��\�q��'�O��{�q|I�C{Ui M�y�!��;�v|����0٤|n���@E�z��\fΑ��w� ��->�݊E ��y�P��#������<?�뽾oj�TN:���y�� �|�!�;��~dI[5P.5�]�_Np�X8
`��	Y��� o{[���;1���Z���u� \������RU�=4����-\}��t��&Zr�k�&�u�)M��ͮ0[��^1eܗ2�뽵ɹ�Q�nV\M�*q3��;9�yTyYUU��k��eп����p;t̄�5z�!�0`�/D*����\�icl`f]+˸��I�r��1[�0�iք�i���;I��gi���谫5�qhU7���R����h�GYz�+yy�ͱ�i��Ɠ��fS��d]k�����U}��:)���I{��մ��!,e��Ŷ*ڑs2�5��^����igR�(a��cO<�gcVr�e1�1t�pc�Cڜ]��!O ݅m�/ [�ݛR�λ��ɠ�������.���hb��g�.���KL��ʗ�5\�\�y���%�`��T.[���<�p(;�ل�Q�C:K�/H���h���	lwX\}r��S:�� �avq!>z嶥++ �ʎV
���uýi#�.����Ɲ����9��Y�m :����k���P�D��[�8�[u{C�;-+�3-�Yz(�[�y}��;�e�vs9 F���[�L=q��h䮷���*D��+D�y���4g72�n2��{�a����6��6�������0��9M֋"���5[^��r����	�Ύ�9b�����yǪoT.���A:�-������F�VnX��8�e}R�J�v5��2s'��XheY�6�a�G�0s}|��q���Z������m�Vy��|��Z��v�^a�u��GWB��˧�=+1�*���k�29���e����6v��U�œ+UF4[m�m��8���m�AUS2ܬ����lS.baLV�խ\����.�����A�K�����c��0EcA�;{%O����mm��)՘���b�����5��[V)"(c)l��]̮:�nC��wm���ېr���Er�]�ۤ��i��i�-�5+�V��L����Ҫ[.4S)�
���8�)��E\l*VRت�(�ʶ����h�՘���T���օ���F�TtYV��AB�ܴ�il*#�V���Q��PF�AV,�\Aj+\�ܦ7E�QB�����,r�r����T�-J*,E��魺�u5s*�*%*�����Ԭ�""(Ո��1�w`w�u���p�4Qf�J��q(�i]6)�Q��`�V�Tm���*�Uq�M�q����'�<ex�w;��{�lU�Ve������F��(b�lV-�b���d�ը��&�S��Z��\�cl�ع[��q��T�;x�ps�#�c�#�|���`�5�^z옫=�7l��g��qX��0�6[���RA/mě�#��S�[:��ɥh����sv.��ѱ<�� �y���S�"睻nkֺ�9�Nd�ɎI��Av��j���b�q�;=�d��Y0[	���^�ڵ��˸Q5�iw5���ݭ�V�s��5�s�x�{��z<��D��O;��fC��-�41�YH'�a��qv�9�ۂ��m����][O�����`�=������&؋��{=qÌ&�*j��5�"<[�e��6sk7�Fܼ�֍N�A�l���SϷl��8�*ۃ�.:�6��8]��Z6xϱ�ۃ#�GnN�-��v�"������7���۸��X$W��յ�v�O(��@g��Y�9��8;7NN��N�\��1����znw;G�-��`��t��)��Ƀm�a�/y�+��"R���)l��u��Tit҉�Y���Ӹ�p��a�<׎ty�=�l0u�z��ku׭�nLt�;�(Gh����/n�8Mqf�؛�v�z�J��k
����l۶����4iS���طVݺ+���%���j^nM�wX��!��[v%���^h���D���wj�;g\h��㍹����](%���k�k^ݍ�=�g����ki��������Аc����Am�^es����ݹlv���]��pR�6v���)��v�/#�[��l����ヶn��V��{c=nެ�gg���ј�a��S�q�4�S����9�)4 ��=�x��V8�۳م�<<,��;;��j�sւ��:�i�:�K�;u���.�Rϵ�C��ׅ��p��ϙ+n�^I+�Iv�=�=%��:�b�5�SO+�/!�s!�2�T�ת�$<�;<[u�Mv�kZg��<.ݳl���[�0�����7n��v�M�����;C<��'�s]6c���H�V��n{<�Ȱ[\ۅ��N�������]F�s��-qs��{vsb8����:\Ŏ$�d���5�8��B����UENm���F�yΐr.+`�8nW���S����Y�vSY�# n��v�D��v-Q�ܽ�=Pojx��7�.��������=�uqsz�\��c�=[a��YweMg`v�ms�n��U�;����u���ҩ��z�/^nnWWXw�6.�䧃s�l��&�І�A���x��AE���Yͻ�I ���؀M�u݇�{#��~�=P�|�y�J��#�L�т]�_G��D��!��517�{7ei$��w��7��v�s<�p�59S.2f��=Q�Uq3��JR)(�M���m� ���� ���S^��ٕ� ��X�d	 ��z���}�*���;6�r��C���V=lt�R� ��m���븋@��q~��̓�IҊv�$܍Q%�e���#{|ׇ�;ޕ��c���~`$ӗ�wi��]�F�m�^.��-�D���hM����7uأj�N�j�H�I|���ssA�>{b������JSSJ&b� N�[b��;�@���a��w��81��Yi39�"!��λ��YJ�(�3�J�"fF��/�Hb>�-�]���	��uо;
O���k���S�Q��<�Z9�����5�G�ou7�e��ު4kVd��p�d�B��Ե�� @N�u݀���~ �M8�8ڴS�l>����B�)4`�ag^�3+�}�mD��]�R͎�ۉn��ހ�"^�D����^uW<�$�"�����^��=�TӞ�KgWĀ߽��d�������U덎�̈��fm���79'F	#;'��'��^���������6���HI��{ܰ ��R,7d'҇>���~��"뗺y��kl1�Δ��Ӹ��Mv�y�8;ms�:;l���~����vV�g�%�e݂ 2;��x ���-���Ì�DN�^�)�ww`|�ݾk�b�ԥU4����u��lA>��vl�ޯm>�Ϭ -7��@/�HZ�L��򮞮j��O٘�KiVdT�>)M(&dq������1��$�ck��e�{o^�v�d߱��WUL���o�u��A��V	xf�*��S�@l�e6���&��\���.+K�f����.��Dw��v�� ��6�芒�2�J�њ��=&��|�y�8����D@�c��)��f0��F!��l���b����3ȢjbE5!I�[���؀�+/����*�(}��߃c��4�@!s�o�@���������ƞ��6�lZ�S���C�nҾ{j�MLY����͵��U��sk ���$�(�$l�G�x���H�����w�wa��1D?_v�S8�3}wH������fg)�܎4�K%�eڰ
}����{/ܼ"2��D�N7�6�$�Hg�7~��i�A�Z����{���i�H ���j� \�Lz�:6���+@q�C������ʙD�*b�L��ѽ�&l�̝Gm�� �U��w`	-=�7s�u��YR;"���2;��]�laN��ҕa�!��Z!&��R]t���=�F�w�l�ǻֆ���i��w(��B3����������dQ4A2!J�f�����ݾ~�VR��4�^k��W}��@dw���x̼�C��	;�6~0�U���ݍ��6��;m��l!���Md����<�&�&eT�K߃c�~e��L���� �˾��+�$�"����J��{3 IW~*DP�H�.͡�m�]���w�[k-G�t�y�O�Wy�w�	,��6@
3ǯ���Fd�[��	����kkf�U}*f�(�\��2 ;ݩH��OO֮���A �����	 ������T�T�`��(g���ʞ	� Oy��dD#���!�l>���{��l2c)�yw�Y쩔L"�)̍��7�h �y�?J�G��D.�*�q �S˻�����̃���ߊ�6'ץtŏ��lɧ�w����Aw��A ;4��fV l�r�Q3f��f���5��Z��m9���L>"}�����eR������Ԉ�d�ۍ�n4�+u�λ>��l>�(��5]�4��I��۫�����qn+]b1rq�l벷�\h�%� 1���z4�Ɖ�v�㎯�u���f��k]�}qKw��K!>�4m�8�[�s�v���+�>�Vv�ǘ��{�q�۲�;Vg۳KUv�c�iw(���5�\�	������b�yí�vE��g�0���.uu�s��t���F�Y����aR����3��cv�3�?~��l�2�ߗ�f�ۋ����� c����a2g&+ֽ޻����~���M�(�e6"j��{6�9��H.?G�{c^d�j�#��Q <������9Ǜ�������U�>�*�*�������0���4�Ax�����x����Q��$��� ����y����[�ĭ�u{�"���ͪWD����D�$<�6�6�{w�s%��겞֟ �}y��+�مj���S%UZVz���@$�J����Y^�x�i[� �U]�4� ���Qng]�q�w�P����>v�W�g�Bݮv�^�"��j�nc�3RN��u��^y'�[_����2DL1H&d|��cm� ��Ɵ��ۙ��/:�ߡp�o=m�#��^(xp������
U���~d��a����5�5y�43Uj�|�[�O����|�|=��LS�Q�C֔��ߵ�B�g��Yׅ�f+Um�n_�~+S�0�w}���ѷ����kzO6�Z�o����c���6��
'M����ʄ�U����b@$�,mM�ĲV:B��F�6I?9˄�J����_<T��q�U�!�S�S'ּ�Ҟ�Q$�yR� ?k��d�I���~�B�Y�-�}��$d�"�nC
�\�볩'?n�{r�װމ+|IғX�vt�qm�i��6/Wnn궳�Dʕ���M�2Ɗ.�9���͛kq[���i'5�O�'{�	2WW�Vr�]/� ��k�� �6����+U���fAǳ� �I��ͺ$�&̻ X+*�ݔ�.�$��[J]��l�3��h�۹�q �o�d f@����k�Y�K�)s��1�ci6��-�fۋ@ ]ݞk�Do5unC���:�E�*��p�ϒ�3*�eFG"�p���o:f�uWSC������ծGF���I�\6|��v��S�;)tu���� ���� �B��m3J�yR���B(��|k���������i ��;V��7{��#��#�y��h��D������� T�jf p����� #�~k!{z���T�u���D��m� dvm�CUk�P���K����8J��:;wl�����	g��^ЍO��^s�<�f���\WngML�!L̕T"�E7yw`����� ��@)͘�;�������� �{|�*-dµIQT�b��s�4^Lyu���elG�|��`��w��VH����&�]��4�MWE����{�1ԄD��`�F���i�	E�?����=��'��ڃ��� !wvy�""��x��Њ����$
T���n_���w黜�c<�}�����h ����ڛwk��ڹa�3w���)�렷�x�M�1r��v���w��OҞ8]I�]{z�fe�L���	�c�V�̐�M��+�@#�N�s�ω5��',�'�2��M���j~ 
��w��]���<g���Aq��H��������J-��&�C�9���k�n6+��@�ۧ���؟M�p����\\n�ߟ����@���TN���
H$�Zs=b�|��$��ݙ�-��W��ۏ��U�	$��C�s�m�$A[������"w5b���={����{W��K�t��ۭ�XLI2����b��ժb�%ER	�=��{Z~ ��w��ҹk���L���$ žo��۾�@=��R"��L27����^�fv���UZA�[�?D -���	 ���m����|��M@��ȷ���]U(��$��7���� ��	�UiA���<�ޔ�b'��$�%vv��D�u��RK�oW���9OE�R6��Î@)lyg��=�2٨e6���2�5܎�,0���W
e��H��
�'St�TO��ki���"���j^��zp�:}�Ճ��I��;�]7\��rqA��{r�"�;c�;nշc���v�6Ųk���%���u�;of׸3�6���u�'L%���ǟlmq��#��>��O��95�1��l:���O�×�8�y���<�C;[d:��՝m�ojum�*Sl�������^y8�Cs7.�(�vy5j�sí�vr�h��&w^���{M��x�Ny��ɺ��Ųv��nv�l�Pċ(:�S�P��
C���Q��7�&  ��n���&��~�ͅþmx� ;3�h��>��!R�˰
��%U�	�s܏�=F7O�D	e�� #c����������H�e]%Q��)6�RD��^�n���I%�޺�I"G�4C�k��9�	��!��w$I��]_ԕ,� �@C�;<�Vgy��H�WG�$�J�z��D .7��2-�2L�=�:&�=����^�1!"��Jff[oZZI$��Z��t�:���i�M���~���o���$���v�?�x?N��ǅ�8�[M�����WOb3��8�|S\�^n���9/����/g�g�����m�� ��^TDc�O���j9ޕ�¤�Ǻ��H��ʣ|�'�P��
C�K�7o�t���_�Aҩ�������GXp7$���hu��f�N�'Y�
�z�p��PC�N���S<t}Sj�or'[\��e�7��Z`��o�"�7� �l��w�U�$��W��$(uiP@�1��TH���$����8$�W�W�u[N���@!_u�� �ȷΡ���f���E��a[����]'��a̓�HW�^�@��t� ��nf��a;�"���4x#b� ª&�Ou�	 ���͞�ْ9�>���h�?%XA'�����"�A��z�L��hF9v���]��躡A��y�Z���uy�o��t��`�'���)�T
�u�gw-� A�<i� o9���q��:�uNW�fV݊E$��W��7���*�$��y��c0AyR�	w��J�8Ǿ� De��, >��9���!���i^3�,�=���Ik�߄-J(������:���@/��;ކ�D_�q�/�G��N��X�6U���s�G9�e]l*�]8�^*䔻��]ٗ2���/5�WYM�DS��E���o�̤����vY�<��MPc�}�h� ���x��IS�m=K�����J����dk㵴��g)|�a*@�;F��rO�ݙےډZI����*]�VZ<��|r���夎[����n62-�49�Y��9*ʼ��K�A�s�L<Ie���|�[r��iA��f`B�t�oz_����`*m��a%`�SV����Vn�P5��@�u���4�W�ػt����\��m)o� �G]�&��vc��icݼ�c:-�"���XN�P���1L$ub��fQ=�*�Θ/#�a�x%�fI��v�EN֋�x)�P���W[�ژ�Z�W:�_f����of���uX��%�u����:cOVuud�@�U�8�!�L�cU#q�����8^A�f�'z%�6���c��총_�CL�ୢO&&]���N������n�#��G���'.�fbu��Ȣ���zq�i��Z�!"�L<����}ø�}�k�*��G��!�G�C{|g�´�W85��x�$^�"����yw���&�휰R�.Z��H�{s�/�Q�,`�ƖS��\���p��������*����׸�ʱ]���u""�HXA�K���l�����%:�ɫ��ɗg��B���%��s�����ٚ��r��f�ٖ�Tge4s1���z�ϸ�0;�q[
Tq\��Ļ�@����h�BZR�(V��K�QƷ.a��G�ۅ�*��G-���v��{)ݓ�����[1�ED��lm)[�f\b�q�n�ª!Pnd.&d�2���f`Tm�J�S.cJ�bR��\�--h�6��F\e+b��E�7��Ej��q�n{v�<aG����v2�C�
��,��5̶��+�qr�W,s+��aG)A�Qn5PA-*��*��V"7.
0U��1s&
[� ���`�iq��QE�Q�j�#G\̭��j�A��\�r�mb�*�K�l�r����[(*շ2���n�l㓻���qܜ����¹Î��ds�m�)#�L���Ю[�**�W0��1Lm��ej`��1������ګ���ĸ�r��!��r�.*�R�V��+F*(�,�1�f[�-�f7lFڸԹj\�2���w:���z��DA���G�g&8�*��	��fȫK�~i�A�{���������O����>2���>�M��MI1*J��C��>�2 �����j��Y�]X�SS���sm ���׋��U?I�5(��b���9d���et �;�
{5�N�Cs���CA�=V����k�������������� �o��0H 4�M���]�zz�������m�kr�I�aADR�f|����|�X��������i _sm@lw[~""�t�nJ���K�pw%"��Rh�%�W��� ��6����A}uѕ-�LF|�{�� [ϛ`�}s<�$��d'O�n0�`�����i$ܗ[dDA�_� |e��ec�XR���>u����Ҕ���p�S�{e�qR�	���g��WeC�q=�>�S����*pޮS>��jN���޼�69 ���`(���H�4R��B�*D�&����ƢV#���&���@�v�A$Fwګ-ǯ�u���&UӟX���[a���'�ٍ�N�`1��v�x��DE�D��7M��F?~�m��|
���` .}�Xn�n��=w�&�ȒD�Mzo���u(�Y�*@��]Z���	[^��υo�z�j���������@|e������%�CV��ׯ k7�I����)I3-�����u��� �;�+<���"@&��$� �c;�aV,��TE)�AJ�G;���q<�I 	��4Ȁ��9`���o�#���69���@f���"j��w*���&�n.�K�7l]�Y��G�n�d��4	8$���j�y*����UZV�Yy84��Fh�3+�w_�u��w����?K�J:g�.�qd��=;'*l���'�R>�pAFׯ��!E��x-+��}�/��ˠ�4�# ��v����ʒq�֜�G]�3s���E�$jv�f��:��UvU۲����!�
���)�ťī�v� ����"�oO7��y�P��G��G�Ք�P'v[���`�\X�Ok]ø�m�)2����݌u�vG��V�r�P9��,���1�ܶ�t=v5.y���Ōg�nׅ�`v+�c�Y�f����Kv3Sf��6L;�������;
\1�[01��8�k�۪� *��sR�1�T|�ۻI$�|��@��n�/zT<��M�Q�}L�d_���K�7�51S(ASU(r�v7��7ޝ��ܤ�=���"�+�-"W��u���H�k0z���������jR�8�w��u�y� 
r�ö/� ���� :/���o���-���$�E)&g�'ϙ�>��7���8~�SA}׼�� ��u�'9�����I�%V
HK�<��@�*��k�=tI${gWS�o>A�3	xyn�u����7�/�)%�y���vl|���1*PB�m�aⶋ�}b����j+Tۮi���������a����%�=�tI9��i�H�s�A]殚�q��L����D0=��	/�Q�5!*Pd�M��I*�^!C�X��OQ�֚W�:*�\��)&���F|��Ŷ��#2��%���-�5<z�4�[w�i�������zr�K;.�>�-��I ���]��J����r{��K�5�A�MT��C���`}��& �eK����޺� ���� �6�;gB8$?&""uiY��>��
�{H {oވ��Q}����Ežu7h�Lp�U[��j��&I�
��$̸^�~Ϙ l[���6��P�R+3�'� ���[�C���{_��ȁD-f�A��.A����Ƿ\��l��]�� ��<��8cvs�~�{��W�����z/��ɂ �6	 �[�M�GV��{�������r��e�"a����%�7jX	VETߜ5�'7��_s~h �|�!������mvR���$��jBT94�pз׏���|�������,Cx��ռ�^렯�S=m�&̧��ezȯ<U��6��4U%|�mԗ�Ӽ��W24���v�t��AH�Bc�'�";�uD��%�/�t���@�
��C�>�q蘬��Z wo�����u��&r�v�j�o"o� ��m��5�"Ȫ��TB�?0q��TCA���r����Q��z��0>�������u���ꊥ��Y��ۃn�:9�ʼ�n'uwR.m����k�v�~�����x&I�*TR�f_	�[�4�x��� �on��+5���v|�o�z��2�o�NViSH)TETIJ��}���b�uu�]��*��| x�"!�n��)�+���ږ�y�2��USTJ���I��b�~ @�ݪ�D�=k\��i�]��q'�^��=���$js0@���VmU�w�$K�:4� ��y� {�}�C��H��s��t�x7�o2�س\��4Ѯ]]��k��ꪕuB����-�J�I�����;
���';Y�v>�O�c��yL{�B��V^��&�$��"��P�����}�p��{�X2Uj���@5]���{������u�o0s�Ny_ kt!�$h��,�1�@�͞���d��v.�b��`?1���)͈�uy+�i�����C��	F�c�F�Ns��Sћ4j�)�ۢ"}��@$��&� �6�����K�eU�|}�筞����	 ����"�H]}��/d��ֽ���o�_K�<�1!.D���uu�����.��6�/7���0��� v��w�u�6�.���I�O�n>�b� ݖ��"u�?42��0�Dfo=�iY뻻�Of)R)T�M(B��{a�2��:�7*H%��P���r��^��DCFX��������Tp�
e�rz]|�dʗ��n��'�ʥ%�+�z�NM�ᛃ8ҏ�������c��(��f��P��Z��ǳ����N�묉"P���ի�����b�2�>�����F�Y���۶x���Z�ݡ}s�V�X��C��n����+e�������r��5��f멷<�;'��z������m����n�v��ǎz3�i��ghȞ�mٵ���\�]t���ּ=��g��������^i����B6G��{��.�;k�nÂ���áܻ�=��.���lr�玍ݲ��έ����n&zP���ƻG���y�����~��m��x�����ۋ�Y}�l ��/��m=�,���m�so~@ ������b��i)�H�C�����|�LC��Lz߷�|� ��=�� ���VIv��{�6�7=�������PR�S33����� cƝ�v(�od�nܜ���@���Ih��>�T	��l�E*�������ٗ�mN{}��w��oކ�^�h"�n�]�:����j�@!f�7�deY3�MTҕ13J��u��:��w��X��y� �u�#;�~h ��m.��]��_����	^;䙨Q1$��yt�k��m=�z� �Fn���e�cn�q�0����F�n8
���U���I%�����ۻ�q���'���y�m2 �Ş� *>Z�-ʍD·j�;��?&-n�w��[<�����X+9�(b�lgq{t�P�m�72�]-|�9[W�^5!�.R��w���v�!�N�ۛ�n�h�vӧ��ԉ�Oğ�u�H�=�����	B�ч�%�}���u�ߎ�ጧ lO��ҽU�q$Ooo;� �P��������U�� F�z�!��n�]�Z��ffR����lO���=��}�n�N �m��@ 7�z���]ٞz�A�zz�aБ����H]A��Q�#J7ďg�m��׺MT��\%�ʗ7 'f���ٽ�w tvcx�!�Lɶ<�Iy��_{�n�
(n�;FV�D��*c�Ӊ2��r�A��u??>���7.媈�H:��� /wyڰ���t�^,Ț�Ϳa��mQ 
��Ҿq#1��*����H��7����X�/��V��Ѐ;���- ��َO��n�h>�{]�����ZQ�J���]� #�<�	 [g����CywQVݲ����'I�wf�"( �Ά��a�<��}(��9@eJ�����c�i�������ɽ�y�(bW3*K[~$'�ͲI$�zm�$r��i8b|�7D֩�M�����QH=O-�� �f:h2�y�g��qj:):�y�ݠ���&eL*S2L�8�� w8��^A���&)~$у�,~1��Udͣ}zǫ���j(�("�"k%��%��M�)ˬ�^��y�Wi]8/���~}r(�
#���+�s1Oݫ��$��"����a/o���s&�����` >6;1��W��JHS5Q�����"�Ǝ^�p�}��, .71�@|�2�{�HNۮ�VТϦx���A�z�0@�Q�U�U��RIǞ� ��z6��`��W�����*����� 
O�d��l�`J��s7zo� ����	w�'�F��ןY{Y����9�V�|vMCEr�tw�'=�b�*�v�1�Cq���	�(G��b��3��s���_����6'�vkfz '�����78%)���z\��Rww������;oE1���`2=uڮ���I���S��7\j�q�aNk���"xv{�m�R��^�mT��uY �7��v]p��)�}��b����uG|�Q�Q�9�~�e�&�W���6�������޻ �}�޿�*,<�����<��&�i ܄�׾۲I���X$O��[�����}v	�ww��'\�#5X���tl�z�� ��]�d�;�ޱ��<�>U;}U�z5��	�]رI��2K��	W��޻��H8}�S�~�M����vUOٛ��`����f�H@��HH@��H@����$�BB����$����$�����$�p$�	'� �$���$���$ I?�	!I�HH@�Y!!I�	!I��IO�H@��B����$����$�@$�	'@�$��1AY&SY�CV!��߀rY��=�ݐ����a�  ƁB�@�  (@ �  �(�)@P$ ((��  �  
     h�)B�
 *� (   @@ %$( (  �(�{�J))P�B�H�EU��T��*EI�TI@����B�$R
�J���U@�����)  Y���DJJ �U�T��t���r��Wv�U	�*�G��TW�)+!�UX�h���J��URQ����ʥ
�Δ�����   �y���J����*�m
�L��ʃ�j�Vc(�u
�ʔ3U%S�:�JYiJU$�( �=�

�U�	QRT)W�(U��H��
P�5UQe�H�q��B����,�Iݹ*�WwHS�<U��&Y�3j{�� �� ����Y��Y�>7v�!�E_y!FO�֊M\��؊��4W=g[���q�}w/�d}Ͼ��Q�u{�pWZ����yw
��ݍ�Z�w&�i�)�@ �  Q)U!*)UH���B �qTEW��w˸��ɪ�<�Ĵ�:�-z�N��Ի�H�B�Ts۪�Z��uU*�ʪW�(ʪ��袮��(�J� ��Ψ�b*\9@�*�6�UL���\ڪ�=۔���%=U34�V-*��RC=���Q@*�O҂�ҕ)TJRJ���*x�T��L���R�j���@Ȟ��z��j�X�^�'���tĜT7T��
�wgQ@B�W� �=�}�	UwnRUX�9֓�A��R[���Y����R��D}k�����^��P	U
W�  T$�$�A H�����U\̚4�qȊ�d��/Y)q��Y��$��]��B���7"���Ri�g�)%  �@@���p��W�tp�ꪡ�P���E�R+=�P��ET�qT;�ɢE2ʪ1�O|}�      ��4RR�1�0!� ��ba4фS�b���10�a�C 4i���P5*� 	�     �ȥJ��Ԧ�IL       ��Ҥ�= ��S `M44�M0�M�L��&���iOУzH�4��ړ���|��|~�����u�"���,�ɝW�j��&kP���*8���L	A��"*?���S���|�
���k��XRT$�TEG���h�`�������_�?�?�N?렯x?����$d��DQ�LC�)���(
����:B(lb,�"���S���C���Ƌ�(#�ߏ������k���:�s��9Ü�9�s��9\�9�@��qT�(*DD�
�w A* *w ⢉�UU�*����(w@�����w$U�(��@��(�PS�;;���u� ^\%V9��D��'�G�
�D��~��?���e~���4a,(��'���|d߻�~m�E���Xر9��
5��M]�s��3.mTt�uQef�Fm�=�b�@C,k��˫+o�7E)��3>��b{Zn��J�T�k�dH�ݦ�%�SX�NJ�(�Cm�xp*�*�!�u�K2l���������;�5��ע[�:��ga�;-mD1����R��f4nF۲[�{[�t�^+����֡4k2� �4ݖ��b����G����◲�^h�uĖ����i�
�Pq�d2*-C���B�RJU5F&��3�f�Ww�����BK�kD �%y�e��0�e�lj.�9 %nA�[�fi��QV�� �ф�b���!�Q���ˡ�2�p"�����)��̃j]t���~�a�82aO,,�O�i�Hcn�]ۇ
r|5Ltd�+��_#���;BJ�r�s�(�b�p��������6���i�l�CU�}qˮ�H�N٤L ��c��<���"�f=��3[Pj$L.��<t7ov-p��y%�)�nCJ�%NLN0�B�l�t��sAOv�\�ǂ�k��*,F7ke�Ŷ�f��ɹaaC	SoV����TT�R��[x����L�[l��*�f�@��Ve��`��c�i�v�i�����.�Y�5�(����C2���� �l
,16i��ɉ���h�k1��͔Y�O-�ie�n��!cw����v��R�r��-�;�]������j�C����Ys*�{KV�X�{���f�ɅUgf�qhySm���M���7)�䦂����g �݋Oؙ��.���X�0ݣ�lͨ�^nmB3q?��j�#��T$�m��N��eX90�ۼ��P�G7r�|���S�2���Hl�e๱Y�v)0n��p6�X��*V3DZ����K�ܱ�2�!&I�yoE曺��)՚g��hG�=��@5I�yA�N�a���a���4��e��w�2enk°fhAԢ$���q��ۼY6��T(�m��;i念"kd(l3Z�b��V����HԼ�f���xʼzs0a��E�H�6싥�i5��aʘ�<�v�q���2�<�U��B�H&[������.d%�Ɉ�n���S4^4.��Z��ہ9l�ei,f]:(h�6�l��Z5-�dӔ-;�YN�d��Z��il+1^�v�XB��
ֹe)�e��L�@ڰ�H	�]f5VVT����&��n��
̥�yDX��x���]2jC���۳L�GfIP�n�;���t�e^�1*��q����nZ�a�/%Kk3f��-P��Kw0�kb9`�ʗ�f�e��s,�H�On`��7�mL���u����M�x�Պ�S,X)<[QmER��,-�5	��I�憦E��4^�����ɕ,��V�f|��ê�9x
C@W�7M�+i;�Sڦ����`j�^�Z4IZNC�B[�1Tm/K��L,d�m�B���Q&-E�L�J
��mz&d���Z��PT�3.$����W�%� iH^��z��4�Q�@���mᙑ]G*ڬoF���[Ӕ%��n�ij:�9w�T�\ݓt\b�.!A�tU���u��DD'XM��5�ۤ�H��,vZ ե�m��������}u�4e
�ysw0�C9�7t�A+�ԯ%���͙I"�hsN=�niǔfV��v+9.+7�'��n^�f��`�p<�`�mM[��X��,F�hO#�̭�-� �$�@Z�N:v��+9��N��gS[m^Tɯ�%io""���5+5u�V�t>�u^�x��1��Т�ZSH�[k2��!(B�DK�	��2n��.`�l���)ܴJ�fh�-�ѷ��`He86�ŨK
Ce�j�ne���V)1YR�T@�fU�5�q9�T6��⧫t�a�����4��]m�`5��<C���*i�L��X�b�z,֥�2�eJ�fѩ���-�ګ�����Mc��ec�Y�L�?��乥���Sݺjo7��g��bь�b���MTv�Իd:q��ƴEwF	n����w�V�D&f\7�B�;�Z�S]��5�eL��X���m�o^�Wd�YY>�9�#űS�ʲQv�)(��_3��: �.�����e`����$�[XsAqLѳMC��6��˶�dUy��5�9O�D�p��V�ݰ��j%��n�n��r���[G!Uo(�ut�\z#L�[�j�7�
)��sk	�U`�Ffbј�Ć���֍k@��PZ	�Z��:���j k3r���KM<x�&���o
�Jd�(TKՎ���nn��Nޗ(v��j�%�)�yb ]��q�W��򚫤k2��&5r�6��w���sm�6��f�sn�ǚ,j)��^k�(�L���(����3��+2=��+���G��r;��4�%��O�v��&i�t�hʺ��2�(v�ޤf��dἐ�)��6����Yb�d�u�۳�λ���m�E�ل��;��L�)H� �j�I,�-�6N"uu{��{8�a�Go�S7}TpT�ӢA�2�T��m�#����7���V���ؒR���<j��T�3Z��R��� B�@I�A����y*b6�o����۶��@m;4�e:��� b���N��Qtlm��X 7%[I;�Q��1n˼�#y��Z�����7�Kʄ�E�4-9%���,XG`�wS˽�w\�>�M��Nmar0N��-��߅M�whL��b�ɖ"cn�2(��1��Y,���i���H^<o_�Td;{�x�K��[��ӥ�U�*ֳ6TX+c��e�%t\��l�r;��y�X�2�8Q1P2���S`ҳ1���֧��K0f�(�9�|�[ M)m�,����JR�q*�ʀ�j�&��b��PɔNHhq���"�oً����z���N)Z�7-���+�L��K^F&�	B���ܕe+�)��+7Vշ��f��1���Ǌ����ݬ��� 7a��b�2�sk�sM� 8(0�L6��T	[N����"�D(�i�- ���"ŧ5�6�3�Fe�x]`�-^9�ı��O"!�C*�X����J�6Sd%L���a���B�9�1�^m@�\qA�������a^�IcS.;D�t^lG �a���w/HX��+h��R�-�b��ݸM��Uܚ��^�wi�L�P�[x;��oXgw]�l���2�͕{.� �&RW@�t��wy�V��7�Xɼư��`S!�uL����jc�Q��%��GjK���X�϶F�R
��U�"�ZDj׊'c�b�I�7��T櫽׶��Y*�������'���r\)�9���h�b�X�R�*�6�x�&�
���� �� bR�Ad�%�%��lۘ2l�a���2�$e����Aʜ�
�@�`�v+��3�2�]+̔��a�Y6�Hϳ$��G�e��^\�v�-:��;yN2���Pѥ��^��Q��dn�䩚ݼ�4d;.-�;v�)^�Kf^T�]����V�[a}>	n�\` �6]k�d�X6��0!���&IY�Gi���֘lڳ.�%`c^d�[LI��4�R�0�q] (U�5��"� <V�,�s1X9��V��to崱�S��L�r ���"�5f�h��-V<�{p�G	*���*(�`�q���W`�nF�6��zY���2f�/YE.�0�Jm�K����9!b�q-�b#�2e�����o0(r*/cp<b��*�Y�-81]�V4�G�e�s[�5�IZ�[�fV����5���f��ˠT͐�g^���f�{j�d��pP2�˩�n%V�kW�L˰��wYoQ.!�LY�Nc!3�SC*U��m��o,�H��R�c�I!Җ��a� 9�c:�]4�HE-�ً@�y{6�86�a�AcX�{`Z~܄pd�U*�p1\���˷N�b�]<Iٙ0V�36��]���DG)�X��HZ��d{�Ԣ��W����˖d���LӺe�ɺַ�����F��,�L�]�m��9��Z�C9��к�}�};a1{V��P��ʖc
Ȅ�3P��2S�q��qM��Si۫-�d���Mv��˻��W���#���0{�Qv�Nd.�ҳ�ЭSɚ��&Q��
�e`Ė�u�[�b�����L�1E>ZE���1=�<D�J[Yb���#f=�UcK�2�`���j�f�Ď��S�jd��i���CL�U��y�[Ֆy�����1{�f���'��L���^Q�hX�����6�B�v���%��vl�����e8��^�r��q�V���m��q����x����%�WD�`چ����!���6�K[w�i�+ ��7,Tp�g�^k� C�S-�ѳ.RǪ��skjI{�Qf ���F=�E;��ma���hdwj�u���R��iTv�ݜ��r��1��Ǻ���z{��B+�-�o.V]��Ջ���k�I�u����ӗ�4[�����f����'C��x����X&n�x��wM���b�y``��f�wki5cC�i=8$i�A�W����0��bar�]�*#[�zMLc.�d�]n�v�O���k*�lyw
�V��}kq�FsHTM[�5n��OҦA9�T4ʔ2��N5r��ͼ�7�b]��"�Si�,ī�-+�̩NLeM�*��aYa�<�,U'��.R��mٹ�W���6e��5C"�V"(i�l*�z t����N�g�y@9@�9u�5�Չ�X��G	�rlwx�9j��b0�*k��KX�3�n�3g�ЭYA�(�:	L�IWp�^5NAGda�cN��%�+5���x��0�F�+��nΣ6�ܤ��ī�pٱ	Z����dlzF��ޕ,��b:S�kو��̌K-�E]ؼsM`��8�F&�yYo,' �}ۚa�����&s�[���6v��A��s.��X7���Ҫ)�QK4�C���h<HX��w1CV�`u���fʻ�ID�+/�X��_[Qi�6�倵�ɢ��&]Y�Қ�`)2�GET�i^��i��2è�f�&n��B�vaJ|�h�%d����a,l�@��-�Y4���)��$Ne�����d"\�����ʱ.�`���q̆<t+2�Z�D��Z��	�z��ұb��؋\��r$A�V	m:�C�GSZ�f�R Dƈt��/�yF8)�e� c"U�qjX ð�ܺ���j�T�]�CQK<^E�/VR [ǘ)��jp��D�Z�����mٙq��@{(ٵ4��Xw��f�70k^���TrL��8��-TwG�u�b�t�B�P{O�ޓMҰ�Cw5/�"E�ۘ�-Ӭ�-�$�-[6��+Y�o4�R���4�f��B[�f��N]��1�x�Y�K�"�x��K;x�W�
���n,	�6��m�
+|S��	U5��b6ܬfe�5�`�F3��ե�36V�W���nZ�#���[n[`��wvU��Ҷ�2�Ԩ݋��튕��Rj�kU�M�7w-���e/�:�Z���;��L�H*f	i�iB �F��[[X���XM]�Z��.oE֝�vM�d�n��1X-b��x��4�eO �-�.lx��/)�#A�>�坿�72���Ѵ�3�+2��;#	F�!��,O��5c%I�o��2��
�3C�G�:n��6Fǚ��X�"\���4�	ZΆ���iq�%'B=����c߭�]�;tw��hh8�׀)�d��j���ù�b��a2��n<�i�nQ��6��Ɖ_��(��l�Q.!dV����r�P����Ub�Z������p�ӷ�a\�6��͘�j*�Ej�,U�;�)#Afǲ��V���
VD��)�{��V��W���T��jײ\۴J��YPk��t��gBm�P�9)Qъ]]�7��j�J�����`�4-R�3З�by��n�%���l,ӛ+a�l=I*�ňL�aB�V�j��,yHT��n�����k�6Xܘ��GBݹ��R�0a�z��;�AB������f�yw�H�M�ϊR�@��m�Uy��ϲf����/3wc2;[Q�����6��=ٶē*|�#�3pn��'���(�#9&F3K�f����Xu�f�<y�%-o/Z�إ�E0+�Yg.�OD�@љ��[�θ��1m* �LfK�:��w+l�1���3**�� inf��k���=yP�y��5�ܶ���W�	B���.;l�1�)Yɏ�E�v;XM�L7Xn��o���M^rf��E?������c�>R������$�P7�{|�/�3�#Kt�[I�<�pލj�lQ�&���*(�< BD��
Ȁ TU�$A$�AI * @�T�E	���FE�DD*QA$D	@@�AdP@ jQA���DEdIFA�J��"�*$�	Q@d���d 
�� dDI A	�T$DDdD@Y�$T�$ARD $ �TdD�UdP��PD* �Ud@��5dUB�*d$TYD�AdQYFD �dEDZ�	"�Q@*(�Q	d�T$$@R������B*�^�������	������c_7��b��� ���&:+{�k�� ����pց ���ת�*����T@�����|���gݏ����b8�e^c���_�{�Q2��$"ֽ���ɥ�|l���ӊ��<��q�9ʃ���cŭ�ϭj6�H�IT�%�_}m�t��]R����\Q��]��r��v�*�e��Ph[����r��QޭY��	�׫0��T�u�M!+ΥjW]ʹ��pS^���-L9�[�W\WV�Δ{�^]ft�����8��9�#=���Y����旣8���-,T6�"媚��|�4�ֳ.ڬn��C�e���NB���c��o��Q��&�Ϣ�{�zˠ�u�|��%ϸ+̂��s2�gN���^�.|`�Yjg7�̒aS��o���S"����f���*껖��ݣt���e�Yf���o]��r�z�b�M�}w��y#�`��zvhY&n�t�VM�2�/�c���j�Õ������oFB
BĤ�WJ��a*�ݥt���8@\�GFa��PY�J�!��ٸn�9���G�Э�(c�3���gH���ݧ�j
����RV��Y�W��7�2q�b!�QV�������WKާJ�ly]�-���d��6&V�Rف�8���[�&
R"�X2��X�:63IUҙ�= �q�	��3�6��J���uc+�7>�Sjlɽ�6�oF0b��B�#1�k��*��L!gj��R�`�x��
��V��s-���\��o
e�-���u�wW�]*nY�̖a|ҽ���.^ee`����Fr�΀!W��&��g{��z��:���k6�iLna�{�e��j;�2�#'���G��6vj�5Z�ٚr���,\	I��骨��.�Ց,�o$��aQT�7�%�X�{��]gZh�T�����`�i��Y�3��!.1n���3�eF>�^N�N���膜��dCg��&�,�:��u�ޫ8�Ո�ۮ{P�[�DZB��Zҩ/ڹ�;Z����8���k���j�4G��.��<�p�))� h�KG�2���Y]]Q����N�9����YAbt)�ǰ��P�ʥ������r����-�:-u�^"+r���ّ�V�ͨv�;�����`J*���p2(�	���d�J�mM�R�^�E720�5j��@i�;$��Kq6L�/�ӛ!�T/T��D�@���t��e��
V{{�����r�b��it�.nڎ����hY(�zis�$���퐡���ҫ9;vKa�f<OJ:5���CL'j��Gή&��tlƨ�h3�k�f�y���Y�i�y�h�W��/�`|��u՛��1NV3gP�1U�"�1�"��1�R�����o�vk)�����fa��
8���攏eu�If�LWA��{#��͌���X���7O]����V�� *�������7���v�}�]�lS�����P*JZV�fVJ�ff��ٕ
x��)�P�Q���F��cm�R\J9�B�$LF�ԛ#6�(��hmA.�>���4e��uyM��<����U9YW�O�*آ����LɏT�BhX/��]�nfu�����)1�N\�`��1�7w��5��EE�t�AN��ou�����.��X2�C�{���*�#�@`g5p�w̅��ST�K'y��'[�ܻ���Jj��]
�Ù�&� ���nd^a�z�|A.��z;,��J���Qz��ߑ�B�Y��#,('ᨍ�ŸƧ��;�o����.R�w�=sK�f��\H���9:�n#����|��JYw�eL�1A���4��v>�k�ѥv�>W�Vjc�;s�Ĥ��捼bm*ھyӰ=��+TB�nWs\N՗C�,��Z��ݷv��IM�sXa}v&ԗ�uKOp�.j݇wz3�e�fRWS+�d=7r�gH:��w{*R�{9��*�ejۼu�g����]��v�طmv{�m��ۗ���l�ɮ�%��b���V,�2^h�*f+�� t:�օ���
� ��͵L���"��,��J��/#�̷y��P	i)tv�)Iqg& F֫��O�䲆 �V�\�nŁ�&��|쌂цp�}Q)+��R�7zB(q�Dk���?�Shi���+��8s�"��&�!�z�X�&��.��a�K:+�68��uv��V,�+v�uNdLa�,n	2�FQA)��s��u�W�hab}����X��y
rŜ+�*���ыj��М�57OU�[;]��3MH2T�:��|2�X0X�����&�]v�k36��Sl.�G�����Vk��F�ݛv^<��N��]��bĨX/ZՈ/	��ej�g)�[����.��5o��V������3B�CGq�y���r�?��ќu�pô"NT��/��P���3�,.�qm똯�KU��z�=a+$1�g�`�th�]-3��FQױ�u�u;+Pb��.�t��l�{2�dY��[5�k��ݭ�Ձtv�\�U���U3�eX����,S����d�h=�`�Q��"�3��:&2��W���!�i�쫥Pp�vP�N��&�׬�#3�R{��,q��:�g�%�}�oXY�C�i�"��]�X������ݔ�60(h�&u�v@k������hL,JcV�f	��^}:Bk���G&Lc��=��{t��o�&Q�O{���7�5ա�.�s6��r�zkCf	�.Rԫ.�)M}�ͮ��QI�Ю��0nj��i�c=:��E��}K�9��):�T�:r
�%L��ҳ2���G���˾�8vӗ�/��k��:�z�YεMi��k@bR=�V�h�֩L��9L�{ׯ�t�s��Blŷ;��5��f*�h{��k�{]���!��{��X�����6��WcW`ኮP�R6���c�
�}}j�݊�b0�����+
�zR\Mj�{����=wc���hm���[�]����3(	�w�%*�[�8�Y�\d��}�;��;X����,X�:�7�@�l��Huֵ|����uZKڅ����CUXK!�oqK�a
��͝�a*M�e��J�N[y|{3�����x��
��|���|/��㿭���J+Y|�{�4�)2HچJ)CUGV�"�PCD���Y���Fi�'�{j��e��!k�2��o[\Vq�k�w������%�ڻ����l��y=ѮRv览�S��`�����3(�@̇w:e	Wz�y\�!hۮ��#��̻����	�"W�p�6��w�u.m��H�A���A}�Q�����K"�e���ޮu-4'*��ެW+�M����C��#'*t��c�F���m�)����q�D����� 4�C��rfQ�ae#X/Jw��J@cΣx��A�kE���U�oj��PIZ�_st����
�G�`����((6�Tk�P�՚ލl*���#/eG#QWS/:��6����b�m�T��ٟ!�������Ìf�z��KOi���j��x]ۄ�0��\*�N�6�3�i�G+�ů�WD�|������� ��	R[����!�ټ�c�[yWs+�Xl���uV��y0l<����_G�d�݌��Z2!�{��R�Ex��t8#M{��=)��Ub�hV(8U���-�K�WX%NWj�+Y/��*��`��̰dkM��D��0�^��zW}k����
�����tNE��x�ܺZ��9������
����{9�Y�p>l�X���,��'%*�#�I�������N��WJ4�ˣ�\E�w}#�k
!ږ��3�`��ᨪ�՛��6Cl�r܂V4z�U���R�ƬY-��}��[�G�:�u\\%��|�<��L�՝��E��wF�J�V)q�'���L�4xRǵcz�p#4�H5�/������J��I����Ѧ�΢�>kwjݷ@n��jww;yh�YMb(�D hZ}}��'V1ל��X��܂���g��^޶�[a���;�r���m;����Ǻ���um`�\��V�;j�fR�����lڷ{���Pή�eqJ�]a�:�+U4V-�]묡z�[����&��U����APx�����(_5�f�}{[Zx)��_s��->a�7;42�Pq��mۻȴ[�r��2uL�/���fn��qۙ�zq��.�6��!�Y�;!#����ט�c6�3q�]^��pvV�V԰�+/;dvp�%� �ۮ�k�7����,�uBd�{y�c`w�u���`At.-���zf,f#S)}eHG=[��C6�_[Ѽ�jЉ�����z�94Ժw�p�+���aD��j��Y0���䍕�D-v!����FP�헶����3�6\S�8e������b���g2�o#�j��$\2�gmd�xV�o#��е�*,����7��6�j� 4}�2�7f��,;��Z�,��yG/6�"���7v&���=9��V��y��*����I�ˑ ~@Ы˙0�d���\��3^�}r�b��!-f���})�����Ϋ��r������"��KL��k&EAu,��;i�V��n����"������Z�m�\@��gm��o$:�5�[���3Q����E������F``�b/e�%�h�,ޢhaC���	�1�ko�(�2;*����ofp�ak�ӕ�yool�.�}%�ٗ��3�K��"�Y�a���2�����/M��9IPhQ�&<D&���A �N�p�"U�[Kl���6j�Y���淖��V�sOU:ޕ�����H�:jv�j���*��]�Zk�sW@��h��k; ��� aw`۽�c(=�<'V]��b�N��s�
�9=�]'`�`����nu<����բ�)n�����,�AGd̶�;ު�Gp�/"%�|S,�-͑:o2���ɋ3�Fk's6�˞�V�:ҩ��39�_e�ü��Wt��eܡ��Nw`�5��n�tى��&k]s���c��o"L�Gf�/vQ�y�Q�;R��|Į�ٴ �a��֒C�i�I�q>���N	/~x�ֹG|)�������t8ѫ@28峃qΰ�[�v��׸oio�4�ڍ�Qq�2�2�'oAV�E(u`B�3Ԟs�׻�fvp�lнϰ��Q��4LL��j��x�Bp��ݖ*����J\#-VԚ�Lg=��!J�es��$���,yݖ��Riu÷�1FاW�[�l����Z y��� db%y��E�n�:��|��Wƭ�*cms�^�(N3�J5�u��[��`[�.��!�������U���p���N F��a�I�n��W>��vuv1��{v:A��h�/�ѭ�/��)��̸�=D�e�ϴ�ɽsx�Ȟa�8g7Pv��\i��ܐ�EvX�C
y���a
Sf����2�{zf�d*��F}t����ݬ�����i��3���0v�[�y�z���]X	�`$&���[�̵���̳{��:�U:�/���X�����f]����?*�rG��9��>�;��:J��ՌX8���
�RU�U�R��_q`���ΠEvgã����$3vjHp��h�mV��:�N��bގ��ů['v)D^���ΠA������bϝMw]�^�m9x�f��vKޗ��g]ʱF1c�R�C����+��ՈE�J�[-.��8*����A"�x��.}4�1��l�,��m����I��{8�r�[2�����o[�����M�Rί��E^c媛�F�c��Cq]Kltrn��Pc���H���{)�������m������N}f����F�	���� $U�O/r��@Tv�����[��o^�wk�r�n2"UX�Eup/����:�$.U�ð�cl/�l7/.V�Zn�~�����fŜ

�U���fQ���n��}�^��*D�n���'Kı�X�@@��o3�0*�g"���/���;�� ��/Nq�5�inn�XQp�.�[��Y5R+�%�pV�ؒт�ڑ���,͋�M��Q�!�k�%�7��t*���t�3�v�z�C;�t3`��t7�uk�܃8!�yx\1P�b��B��M`���k��@�ؘ܃�jx�2�����\�z#q=Y���ë��Զ�-�����Ѩ ���q^:{A�޺ń>̳��I�{�_=MU��CǶ�8p�KT��ȹv��4�:�;ٙ:�U����v)wks;���)6̍&\�1cFFސ�Ll<��*u��:i=.A;�6�뿜o�8j.%�IӷPtͺւ�}/m� ;�d",3�n��л��ﳶ���JK�`�|�3��M5��;�;��+ˁ�fi̻cK��ө;K���Ii|/��YgY.�"
:�ݓ�5��̃��#")g^��޿EF,a $�x*���׻�����S�$����<������W��'�s�O�7��"��"�ݣ���fɜ�1����4&�QY������f,���z��0�6�녽�e\ԎqX]�afEm]��Y��!68��i1��"Q��6�b�����Uճ9�Y�Sk��f��TBmj�űt�6ܶ�Y]�v
.hSch�Զ���Pv��D�j��M�1�5�ce,.�HvUѱ]N&�YoPZK4jh��ԗ`�.%6��6���qn�iE��I��rEr��3�B�H�R'R���6�6pSK�Z��Ms�m45��t��7 cDCm0b9H`6�4a�!Zͦ�p���`,D3rUځU�����--�&��k�J�GGZ��,�\kŘV�34M���v��A�R:��E-���M�*4%�U�Y���
�KA\��\���ڥ5��j�l+Pt3s��IHh�nn��B,ؙ��4/�.Ąf�k�.P�2�uK\vH�w8&!���l7=�j�A
�dњѺ����T�ab�]s4b�f,i�1�S�Ù�be�b=�����meF�k��%�r]v�p+s�l���Zp�5��]��ބ
�Mr���V�n.êa��[��J$ȸI[{:i��K��ۡbˊ��שEP�.�%i�]T����p�0�k���/1MFͨ����gm��4��Ҵ![�"�1S]R�ֽbK[��m��Bf�M�L�ApM\�+"k���<k�+W8�1J0�*kX���#l�8�V;t�.�Reͩ\R�XP��6!��z������S-!R��E&���T�E��[�j�Ro5Jm�*�� v���a���a֦I�*��01�Mp]���HM5u���Xd���nMsev��s��.6�Q�Y�M	�Ž�Y�Cm����K����JGB�]�4�cV:��X�P��u�,κ�H�l,�K���]LRQ�4�Rݕ�����V��f�a�MD�GV�]D��Q2�mĦ��%YMl!�#�Mt� ��v���v�� �`�AiG[0�CB2�S ]���2A�f%�Ųד��:��gEZ���6����*��2�1�C��u��[4t�l/
��i��n:�+.��Y�iZJ�����(J�l�ΰ��j�`�gm��ͺU"JݔsD�мrK�$�I���.�I���cRk[�k�/2���L���t�nuα�j���͆S��uI��Iv���ؒ�5(Ff���(q`�v�T�v��/,ае{!,v�&Xņ�ĥ�Z�t�Δ���cZ;`��e�-��&K�Z*ZjQb��fÛ�21"еVT��RY�Y�8J�jm�����tv#en1x\���A6e"�Ҫ�-�L��]�D Ue�X1$�6"�֚-�Z�٢�rK�$�IE��5�����r�6���(X�]4�u;LJX�CJe&��S�eZ̮�U�C)N�h3h�"ᔃN�s1&!�C�F���v��\����r-t��m���h�l[r��DK(h�9!u�2��H�l�e��ⱀ�Jh�6�fl�aR�jM	��5ݖ8�&!��(]r���Vn,.�n�!,U\L��,4]&�������B�˛�-��d�$�.�b�YM���,T��R�K#��%���Xk��f@1�l%)х�p�,9ٰ&�06Ӯ�ú�/1U]�\n�%ZG���V�G[R��,mJ�,!��U����s[2��M�0�����)4R���$	�
E��#`ds5Ke �M��b�åWZ=m�9�J(�+���\�ܹ�76�{k@��K�#6ЯjMi��J�K�̆lS�q(�\ٮ�L	�M�R�[T�A�X�e���J:��W���[�f�v-YGmI���{[�heM͆�e�b�L9�ZF��4x��ڍ�%�6rL�)i3,J��F�b��ij+1�¸�44,���D�Y25Рٽoh��I����ŉ�2pFhhK�j+*�&jZ�eʲT���b0�K���{i����í���p0�Zm�-���m�a�J\�s+���-�ͱ\��1�ՇXŔI��.ԍ�֝�2��K�\�5Dl�8̳b�LQ�eK�=L���]�(��3L����9Y�,�E���h�
�Lʹ�lX��
D�ңib����6�W@�H��W&�V��7<���X])/�T֌����\�ݺ�	H�/lf�X�qK2�t-4ȎcԣW	] �l�Yl��kh��k3ˣG7kd��YP�Z���e���Q�i�Ǝ��vڐ`]57d�J<]��Fv�jfEw4m늎5gRX��̷B�U�S���m��L�5"F�e3q�R�ړ6Rm�e�Wh���7Ar�mK�&&�1X�0M��jqcf�I��LD���11a��6�lE�@��v�u�-��Z�2���iZR:Yn�x��sBKm*�
K.5(͍�d�QMks)D-�v�B1�+šAꖕ�v� V��h3M h�c���j��WJ�#њVb�K*�Yi���h(˓d#gtY,��v��n��y��U7j٪�,,�4Kf6x ;]b�D�]�k+����%��Y
b�imBVV�j1�y�sjZm��70�t+E�0���F�X��;�u������q���U�\ٲ9�k�F�*�PC 2�.�)+�
�b+5�sD�n�a#[�j����κ��6���I�iLV��@Fkebh*
��4��b�p�ki�Jn�ƀZT)+�����sX�F��0&�[����^Zn�WgU�ٰ�6;vY��ELmZ;st����k%��0��X�x�j�lŹq6�-����������8�" �����%� �B��ia+R˥�.a���"�(��٥�������\i�]C
8�mJ�8Rݣ�K�]�cSZJ�.q��7!�ݬ]�������ife)q��;8�3yp5��A���f5�B[�P%
����iC�`�`��Jsp�]l*�-�馃l],Rj�%�I���*mك����6cT�Z���h�Y1��r�n��m�MF�EJ�/h�s��h�ZJ�	�n6h��g5SV�R�')���gW�p�\;�0��B�ۭ��
*��L	���5.p[^4EȘ4e�[���L7�T�s�%���]`��*$&7��x��q��ml�d�E��bS�����n��I�ZԦB������.!�f���`���5�Y����ر�XR�3M�VE!�Wh��jA!�)�\�
�mѩ�-�9\jF"����`N����6�u�:�BS��R�@�!	��!��k)3ce��Z���r�8�eb=�Sk�ڳBޖP $�7[J<��mԱG-�V�:��nf����l���f0�l�D�Պf�Ƒ�XBf��If�����6��c��\,�rd�������űz�c���(�X��Ճk
�ZĄK-�k{.� ��7�b� [�KaM\���5�1*�����n��M��I�I,�ĖV�mi^R�B)ڀM����%Gb�v�,t��)�y�0LM�)�]�Bh�6�bQ1]�6ѬM��ó���WM�� ƺ<�t�cP�c��0�(K��+�P4X�2][�ԙq5��Yfb+a��;:WX���6q�����{T ֩�I���ى�޷:e�Ԁ�o�Xh[f�[W������I]�
���mkq0A��:�a�Lf�[n��h�Z͋��!3A6h݆��,�0��% h�\k4qR�6�au�)[���]�m�&f����؈�e�����%tcg����k���4��]6��z��b��Ĭ����"a�L8h	E����.Դh��3������q,F�7k�HFl��ri[� -�F��eqp�Dmֵj$.��I�s-�)FA]��h�KTΣ���^�g4���@�bJ�)�T���.��L�ašP.�w\J��c@���"]���f4���C\�h\*fd��5։R6n����`�s��.B\�ͳl�Qm�^��cZ��܆�qj�Z�&h[HA�VM�&��uڂ�KP��B��k �f�x��Ѷ; ���6�@H�hp�4f�.�4&љs,3*�+
��`���t��DPy.��-���e����vx�N4�+X#�F7fZ�6�%@��M����U�.��x�#%c�,b��V]�Wh�(�r�Hi�[,Z�-��%�0V2�L&��i��a�pR#ٗ\���ͮ�KY�p����{�5��*�4�l]�%�1ږ�;L�����,�6�̰vb���u��J]*�2���+^p���e��������frp�
�W*���S�aa���
�V��h��"͢m��\`��J�Ғ�e�]e�v��Huss��tp�k5�����[���V��KZ�jԢ[�4L�9H8���5���s4�] �4�\��[IJ)5ٶ;�+rXMqB5%2�ț�EL�D��@FZ�#�W``��j���fM\�VPf�,�0��b�Ϲ}�5���b�A5r��եF�b8$��rDdN	�1 D"-4ҾIbJQY"*ZBƠ���bm�H(�"@�BU�"H�18!@����0T��4�JR4� AU�UR!ħ?% �?�L���!<s�$�B5�x��)�a�1�����2��HY>	ϛB����&��!J�l��(�$�@�̾R�"�щN��E�%��@�e�d�T�Icb�H.%�mz�L�e�����"�[`T�J��uV��
�u���!�*���M2`�����bK)l��ev���|֖R���W�z�F������%|_ �X�YF�e P:��:���kI*���[�8�$�`V!�N���g8;�Nb�
�1��އs�U"�UU��5�z��r]�Lc{')�����&� �-��V14hEs�fy��K2:j�본�L�]�-`�4L�h�ڏ"�e�3��W��V.�k#(,��L+,�Mf����K'�^F�n22��n��4Ձ�Jr�Pc��k���c&Z8̱�N�&�l�-�u�f��fX�B�˙�Y]U�+XRcT����o�$ts(uΖ�d1�5Vb.%>�L�Q��n0�ElB�YPڌ]M�L�4.R�	t`F��b#�qz��)UM�ػEG��JB�j�#�,�4-�a�I�0%�x\Qr���n�3�λ6��݉�����Vi�F��X��a���hb���z���E�v��������b�݉m��9���B��U^ƚ�������K.���R��밚L�E�o��j�i�5�[�j1ũ�q�C��0iPJ�k�e��Zc&e��HT���Kdю����u��v�FX�jh�Y�ac�K�	JKB�.q@��70�k��CV
9�U[cwZ#6w��.�h]m���+n�0�BgA֍��MVW���il�jIB:ǭbf��K\v��kvCc�,kaղ�6]2�Ś�N�9�cJ�Ltmę��P��,i[�[�o	)E)����%ģ�F�p�Ym35�=��m*ˍ�z��=O]%�k� �XSt1-��0͜m[B��\�D,v[t c�3f*�ћp��Ui5�t+E����-#�T�֭sD�XYEŅub&�Gk���M,�]�p���<ܤ�Tp\m�����Լ��n�Q��7�b[Kk�2�MK3��5[.5�%��툌h��ɨ(U+	R�s�aÝ��Rr�(���YT�fW7��l�1E�)�)
$�]v�V��-@Dӻ��CrK m��5 ��T�ex
X��ZFZR�=o) `ҰP�J��6�X�j��R���-![ Q����BKIT(�C���X����bRV��xH2�e�� J�IF���ȥHPcachֱ �%�e��h��hYm��)�4�k@	��CX[���,������*�K(m@ƥ�����[�.c1��O�G�{3n� ��(	��I�"%'���ն�	���r��r��֮���� Մ:��R^K��g%�b׵��+� �ŒM��Bh$��٭l>1J���B~��4=�ZWv�
̢p�t� A!x�P��D��VEnˉ�yt�I^��O�{]'D� �!@Քq\��TTDp�+�� ����)$m�� �g���f�'���2��Η!4
���-�Y�|k�:l�h�v�]�!����7�$�=����H�Bk�Mj�g�O���{)�������VP�����%&��#.��m�,#
[֖.�q��έ� �Ȼ
�,>&�L�&�9Sd�=���/���-n�4�OL��M�t�>�8����E�t�a?Q?��F��[��U@�U�j8����WŮ���)M�غ�ݣ#��*vڊ���^�5����ז����x�"�H��КH��άE�t�G��3�r�)A^��YAQ�(IF�<��$�D���%h����ޑ���G��'D�$�g�J��6��	+H�B�e���wTd����)$�Hf{d��M��2{��	��&7�Mۤ�4 0RB�P1�s�0�wѻb.�y��cw�H�Bh$�A=�wh�/��Y�J�ԭ�P�L�!!�fK��C*7��ڍ�h�a(ݺ踅�uk�A���;aJ1$DH�U<�vP�A"{[���R�w����opݶ=p��B�t�Q ���%j�,��*P�l�e�(&�Ļ/��"�$�	!��ݤ�I��\�Grͽ3�Rݴ}ۗs��b��*��i\�{ْ} q���D�EO!qD�k��"2s귑���C�]C�	隹���(�cϧ���ټ����'Q��<le�sM���E�l������D��uD�H'�(ˏ�����!��u�*�.~k�2�_ ��Z�ŤA%���ɰ� �s���>a�b��I-=��4���V�V�
��x���I&�5R�5�|�A!4�@	.�ۻ�D�,��(�l�u	%G7��^L5EP���R4*�XH�YF�ڳA��c�[�%�&��V4�IH��0������"�v
/5�˺$=�)@ #3Γ�{[�3TЌW���R��ذ-#<C�R�I&Ǘ#r�RA!a�Q�{�d�7�U��$��i ����I$�|�k��p籱>2V����B�I�M��?I��*l�MQ=�.��{1&N���1�X�IΡ4^ٺ$����RW%~���\�����w'�I�en�͠�#��M$J�{��J�0������`��2���g��WX��`�q��Z���V��Y�jb�Ջ��Fq��ڱ���;%���S1��Te�.T'뒴JI]���(IF�<��L�Iy,���1�C����$�ļ���(��"i$����wk���Z/*����u�8֤%�m�D�i2��1f�M����+�P[T��Ct��ʘ��	5}�6�I�B  �B}��^j|��Z��Ϩ�̖řf�5RuD�
 0���@�*��:1	{��|go(h�MfyRe$�Y���[��e^�WX�c��	�:��e(�ڤ�R�_c�ɪ$�N�:�h��>�"z许�XHn9A#D��k���WPB�!R���>̜}�NKk=�6��4��?�$�sݭωA"�>��}W�:4m��褆[�47��v����J��쒪I'������56���&��'s�X�W�I�{�B�������v�fTk$�ﶍ�Ǫ�7�trnVTL�5f�u3E���	�����b��~Y���g7~�r��X�W�F����q,l`�R�;\h�]]h�Kh#��܋R8U�#ˉn1���m�SMZf��ܦ��A�mgT���i�3�j�9]���)��Y�,�R˝
�0�ȗ�r��J�U���.[bͥq�B���.����-0��5(���4t1�����F�؍� ʷ�h�%!j�.nZb��%K.��p�UvƘ��3Xmt�B͈��ڼ�3��~�󼂙�Q>9���RA$�suF�D�\olU��>I�~t�ĒI�v�	h
Uթ$�Q$v���6��Y���^H~�Hy+|ꉴ�qݱ~�W�J7�2"�����A@��HJ(����%Bh�KO���A-��XpfJ���$���;�Z)$�olQ�dqk��)B"Dʋ7�#q�d��'��$�zؔH���rfyR��fs���?T&:��B"�"m����$A�H�Cֻ�f��I��H$��ܘ�3<�2g�=>'�����Ƌhm
��ͽG�Z�hF�T���*��bK�U�.�ݩ����YI_x�̒=��N@#3Γ'١+�.��Y���%B	&���R�?d�ϲ��	m|0T~T���Ay�_��r����r�b@��)��װ+ �ɢ޲.����� -���`I�l�N왋lꈜ����+��8��$��r��I��&H	�R��iV���К��]I!jT� �$�^�ZH��ȡI$�ї�`D�*v�77y�$�,z���9�t�t i�]��J(��<*�Y�X�{���k�$��4I �9�W��M\�O/E>��xq�We�H#ShF�
�%�K���Z��'��dٷeNOb��I��2@'�풡���_~���|�o�`ޱ+i6h���t6el�喰�1Jװ�Y�����ZkX���mO_28I����h�g�ITK�����>Qd �&��t�o�MڢW�RW�ǰ��r�{��w�Ǵ�@4'k��$��r� @��/j^�NF��>uv�+ ��8i�:d� L�6 �N��kwROyy�V<�o��2a<�SMWx���0ak���J�t>z��h�uwOF�gs��,���S��;�=+:��.���d�H^9I's���Ȋ�N�:�ZF͊ ���v/��?h���O�OĀs}�J$�h��j���#J�����I�I���j�X�Q@�^ۢM��>w�S�FΜ݊�w�&�A$����PIy-�s~�\-�pf���\0A��X�ΗY��]/g;�bm���x��eB�+�Y�{ÉUhU�A^5y��&�%n�Tl$�H.�sv��;��Y��!�s["XH��u�����(B"�"mZF�2�ɞ�ށo\a�s�Iԉ^����"W���7h����C�+�D��t`i��+�)+���I��H��G$�#q��M�O|t��'R%yk�w�D���sv��+�0�L"�|l��#�v��η�I���I$��뛴�D{q��ԝ��ļI�)<�X�3�ٜ�V�����6t�	����4+�-{zz����D�6�1�5Kw�M�S{wF �H��QA�=ٶ*�Iy!���K�V���y�ܠv����zI� $�u��+�#�(I-�JF�\ƨ�F���+Io*��8�ᔖ:��e�p$�Q��ט<Ꙁ�:g礝_��J�%9�+��H$�Gj`({q�d�o�I�����N��ۢl$��w9�i�pԤ@�2dچ��O�I1W����xV�;<�P�HIywk���(��A"\�^kż�ю���&��]Hп��J�2�vJpIܑ^��D����fqՙ׸�H��j���^�T�~}���i\��s-BJ�;�+���;�F����"Qz�I4�nv_VZnې`�ˢI2�e�Y
���VA���5��M�D�3��3R�[� �ǂED�����I��W�$�s��|�bL�鰡�̊��;��~>��A����W���e�$��LǕ�k���o.�cm�W}�2���<������q��B��y�^VSG��v�g�)3�c��l3�\V�n�2A�5au���EG6��ZJ�J��cf��K���.�*6XƘ)���.@HT�Jė�����p�f�5e)�!]cD3���WC�fQ�%c�mp�@ln��h˔@v�R9�K�Q)�.�R8̨%b*���#n�u�]��]�(KLuJ��ʹ�h�u�e�ج[��&����,n�.36���&H&گ&�a��`�жD�J��|��ͺ�PH6�I��K���()�����n�%4�lZ+� q�MIk�D�%I��MGm0- ��c�h��[uk� �|�M�In{d����i����Bh/��Ī�B� �S�W9���	>����կuXj-Ps��q$�-�M���;�428J=ȑ4�3x��٢�$�A�Ƞ) ��K����	/$�K�9��tuжo3:��$/y����`H"�v���vdbQ'�G���3���֓����I��;�O� {}�����o�.��W�su��i0�.��Yk�s�hg��bhе(ۊ�+�����?D�Mp���C;(W����W�D��Z���AО��q��t�d���%BR�C��J�+�(T���t�	1��W�zc�xT��.k��DsQ�ڻ�";F<w��>�bp��WYg�@{����1b��n\,���$��Ew�qRC��O$I��	'��O�4I'=�S�A���'fq�2�&I�p��V ( b�b4I$n�o�d����!a���7LKH��8��I�{Sg��Ut��A��\�ZA�iNb�� ǏЀI'��RQ �g�*�.�am&�ďOk��+�5dU��R�-�'�@��*B��7xK�=�I<�wa%䗒��n�A%��I��t��o޴��)X��A*ɻ���j;�u(i��,V�uK�tɵcTu\�~����k����0f���~${ݱ�I�O�3ΐb�u������$�>��>��d��H��!�Hb�Kr3�t���㫴�$�s{T�ѢH���7)7</Ņ��^N�	K��Wʕի�R;���RA�$�b@����/� G���< �-?�w<��7?ʆ��{�)�Dx`�|]+����Qy�YhSOj���b(#��I�I��ܬ�`m��t4�C�`"�s&�bS}F:c6�)��ͭ��t���.c��#@�Y���I�Y��� j=� r�P�;�:��M��ɽlѲ������,wk]J�ޖyu⡒�#;�M�Ja�׌Q܆��E����0��3
�#pe�z���k1����u��P��>7�sެ[w|6h*���゠{��[��.��(a[u�nN�gnN�+gwe�D���fa���Z��E���|ҕܴ���\����`�kj�*�+�������ql�����V̌������JY�@;�<�:�fԭ�w���ƫ#�@�WME����"DT.�OZynq����j�Ǚl��)�K8�AJ53{4W�V�ۂ�^�
�v���G�]e3�K;7q��{cLK�<7�5i<��gM�����W�� �`�d�ٟ?;	_��5�Cd(m#��S�2,���{:�r'{s;�S��u��Knv]���Me��L^q�.�	[)�k�s�#�i	�k�.���4��� �V"�^�y;6�N��闓�ǣ~뮲�ݮ���+|�.��r�]���,�%N \ h �ʂ������9WΔ����嫙���_by��uy����^�^;�Q����r>݋d���y#��y��l��us�݄��9!��I�B-����HԔS�@�R�)IW�INI��X���B�N��nz��ف�	��NħC��a�3�!�X1FcĤJ�b�N��D @�:$ ���#<j�學�	)�I�[a  �� Y��Ýł���N�%aq���	N#g���N ��au��C��K���Աh�R��sOV$����kBOW���k�8$�)a�<�l�G�!����d��K	�HU-��rH!�^|M�/q
D��Y�'Á��U"+�"NHg�̱Hppt�R*�X�A֐ @�9&) AS�P�;�t�"JZ�RP;�1�JS	�
0�rro� �g�2	��B�咒RXIHe�HC��C(��u��1�k,@�����a H	 LJ���eN��Wi�JI�ԗ&�'N�D�Z�$��W� IH��)&&:��
w'v: ���"ڝVbA{�V'1e~>HNsd��%����Hft��$�Jl
�X�@���ޭ�Fk�<P �٭	$�y�&������t������I9R�q�w��@�2d��@�t+ԒH%�k��7�El��G�y$>ٻI$�^Вh$��;�h�&*0z�t�f�5�@в�MAl�h1l��#(�tK`����.2�����F���T��ȟ�$�NT�$�k��$�ѷ{���}����D��Γ&�p	B���,{�li)^J�HzD��k'�&I$�}��*��i��w��P�c�R$_���i"o9ՋK�!�E�|�MÓ�c�f\�y$@��Bk�/$��;�HL�F�C3&
�I�ޜ��;i W"� ��K�]ݤ�'w��K��jh}�Z��}��a�ˌ�X���H]N�]uu���2p0`+�<���6��������evR#M�����"�7�v~I�m	������!�%\ߕ�mش��H��ߪ�
x0<'H��V�?=��2Ēw{�{��>|����L���CfݘeUfSd�-hn�xu�W�l�Ld�`0�>��g��f����4<��z�A'�ՋK��o9�	c��˚ȓ��&�Iy$swv��.tJ��R&�&c�=V�Pxve�p�����"Lp��Z_@7���I$����a)ؼ���vj��KI7�(aH"�w��~Η�H�H��;�Z	$�*����V�u���K	$���wh���[���-^ץR$_l��\8�Q|$���V-�C#���	$�9}BHq��ؗc��F�21�!��uj��T���:��$;r(Rv�P��Ui$�[\X�He�'~6jzl�W�X��u�	�^�Q�)v��;�g��	��3�\U�s�2��������V�Ѩ����Xb��A嗴�ٻm����'h���#
�&&�
hPn��8@�5c.�`4m��"��Q����:j�BPsq����!!jYE�u#jkm��ֲ��A�����.�u�ƅ����J������D䭩��WJř&�YTUn�M��mD�e�e��Zk�R\�p�դH�3-˵؉L�VV�2Jv	��	�s��eYJ�J2��Z����6��g��kY59줺:lፔV(1,D�����R ę)��^݁h��'�|��Ođ�Γ&���E��=��{�A$a�m����E~�ֈ$�C���_1դD���S�V- �	/���� �Γ���uw�{���
��	�j�]��T��¿H�$�5��ɢ@�=r��9��oo��BA$��]��5�ʓ��/�ҐD/��"��fJ'nZȔ37�D�`�:I�g;}b�.|�^�>��??��)R$�_	(ן:uL�I3=���������XH��ȟ��	T@���v-u)�S_)�&���'�pB`���d��Q�v2�KH�Z�'f��Ji��U�m Keq>�ȣV��g����$��ȒM�g;�H�sVѼ��ݱb� ��t�&��<O]�Š����BI�^���g߉���[J�������s�n��]Y��=/��Eීs���8�ܖ4�c���W�`�i-}���M��I��&�I/.�wD�[T��Y�9r���b�
���(5Ư���J�K���Z%%
F�ՙs��^�x��IԆ�5䗒�|�ۣ���(D��P�O����Jn�����H�*t)$��Vۻ$�#y���,��I��:O�S�'JAQ_Y���}��!4I	j|⧺P����k�9�Bh$�^]���+�%���\�ڍ��p/W� `��&ֲ嘍�,Η�v)u�n���(��>}����"RJ'��yR$��^nU�I ��.ǒ�!'�*����E���ݮ1wC�U~E�`�)�>3�O�$�4 ���T<�{!�A$���%'��2���~>����h��7Ò>X�,��
���y݋H$�Mv���	 �Υ�$ �%ѿL��0(�,UM����M��n9�ՁsY쫾��_
�6U�΅9�-[�w�%2�|��/~瓡ǘ��иȊ�1�r�g�| ��;�eJ�F߶؁�WV	$P�1����Q:k��Q��F��Hd=qvI/MЀ�vdbܻ�E�$�Om߭!vrc���&�)m�6��	q�(Ԯ���]�XW��/��o2�A#��q`Z$��n��b7g�v��1Ys-1t\[�v����D�#f 6���A�5����.��!O�D��n��Iy.O�ͯ$�C�t �ל1�]��-h���F��#M"0H�����jC���h��,\���,$N��M���&�A4��O�`�]]��L��D9R�L�NQ<g�R��4N�MI&��Bq�nk%,��h�\���s� ��i8��tN7��f1Yf�$��2��)/�r"�I#��_���9�Ak�B���^9�vj���ĂZ��.��"�n�|���oq��ʬ�3D��[�'b��ű{Q��0���G���-#\F��H���MD�'�n9�B�8ꬍuA%�Ob��$�-t"�%��x�U�d���UuJ�V.�J�+���Ca�Gd�HݎɊU��g�w��ɠ���(O.��A-:�P��# $��e݄�v�+xnaL=qb�%b�B	�UI=�zL�� ����h���_Su+>�P�I5�uպ${=��*��ly�-lN�Y��9	���"��"I������DL�c�B~$�����e�|�8uȂh$����3 �&P���EXKU��f�۰bP{)/%g*E	K�$��n���$K#y���5Ty��(�ul�.oƏ �XI
?���H@5D���Vi�������9*�T%;���A$�7�X���{���ޏ���4+ dL���3Hm�] �� W�8J(�AA��fv����A�,��a�ԃYda̝��]ok�<���X�L��`ʭq��MX���_k� �e[�f3:$W]Li��IG�u���35�Msl$fb\W:\�1�a���T�;!�Ԧ���]cK!p�&�3�`����ZYb`����+�Jde�U�$� v��R��Bf8��m`e3e�WL7[�ƹ��4[eH����kn٣L��XJ�qU]ef�-t6\&H�kD�KY�,�k�ѶL�Z�.)�����:�(1+�[��~��Հ�I1>0,t�I'u�Q��+��.�"+�goLD=������$���Đb�Q��(j�2��>ˁD��	��<�a�����J���6�Y�/֊�E�:�f���sw�HU	����ТeY�뺢�A-_k�6�%�������^H�ܫ�IK#y��B����H�m|$>M���c65���IU[���C�#c�ŒM�MЃ�u��7.U����݋K�T+2e�+�f%˳nl���P�WK��s{�$��Hc˻��	/-����0D�K�B)!�����@q.!D�,� �x<GT�-�5� �l�5��&`%�_~~��o-J:d�rj/k�i$�i�6�I.MЊ	9X�5��Ӵ��F$�r���CK��e �����:t�'�����=�G獾�5z����,W�f�s���q�^b�J�>�2I�5\�����`��t`M��Üb���1�m������i �	!��8�	$�-ȊH���:u�d�~�L���v��Ta��}%R��A.:�A���J
w��wR%����Ԩ��à��ƈ��Тe}n>��&o��i��8�K��m$�K��&�AvvZ�T���_�H(���3	�nI����ܪF�K� ��:�Z���R��.�I$�I/$��9܆�_�Uܶ�:H�i*"����S��RlWm���6Ι6�y6��GK���|�g�]�}���h$��iȡ	�I���Ӈi�Y�9)\wt]��H�t$�,�Q�����XW�lm�������s��V�Is�ARV��G_�wh��2(�2�}��jAp�8Y@+I%b�[#$^K���H$���Q����T_�T�k
�(��\��2oS����`�\ŵ�k�6���.�F�뤊G���3X��n�{f��	ݼ��~�����"i$��݋H]����D��Q�W��7����r�$�/�*ud�$����$�Ido8v����ګd�W7�����aQ��B���2|{�#�Ej�qU�!kv_]BfK�6���	%���z�I/����	S����^�Fܕ���;&�tK�V#��6�k��r������TG�H,j����|w���B�I%�:��I�G|��s�2nG�fP�	/$~9��ī@s#�$*�Y����[�Σu������K�$��:�H��y�h�y�b�f�U�Z��G��	}mB��Ѵ�M>qW�Br�d܈ԏĉ����D�=�	��xq�(v�HE(��u�꣛���4O�u�I �.��	"�П��2�_|Rv��y�W�
(�㳦��&�1[/�dڞ���H;�/y�a�����j��/$����l9hLN&�����5��I��%Bk������D�Ta�ٟ�?h���l�(���D�)$��R��qv�#9ȚJٌ���Wf	�]jLU�	F���[����k+hb]��M�b9*������J�DDL��=̺$�\�]ͤ�K�=�����ӡm��xm�g���@�^�6*'�p�%%�v}t*�&���]�3�+b��xZI�8�I$��uI�Iٺ��(�B'�>�J@s#�$DH��.��.͹�W�����K�Uk��o�Q�^�IѺ≴�9΄�$yg�� �K�+�>��fL��<���+۹�A$_:A$�]��ōEv�<��:��N+v(ߌ���B�f-$��Q|�)�D�}ۮC��wMo�/5��%�-��!$�?vКH�?���U.���*Sa���v�?P�g32�ʱwݸ�;P�䧃5����:X�h������m���0NB���3Ou�W��m�ͽ�@��	ͽ���a�c�|�+d��a�0�x_dw��2����+h��Q�#"�$F�h�զ +�18[A\k��{�H��{Z�0-o)��pB��Ҽ�쫺�K�q��[����/'p�:�Nƕf�8nJ�f��<��$ek�(J����BEtoi����f���>��=��i��IPh5ك.���ѴF��a�2������k\��#U$�,�cLܡ�W�7DH&a���T*�wJw�4Pc[���30�4��S���aT�8����25Cw3\�op�9b���3:�a�U��bȷ�=���%���}[w�ύ�{��-Pe�1���t1Kt.僛�gSpn=L��oSf��W�jծs�����	�N�f�݃�kHp�R���7C�r��˽�7�\�ݝMl�Ұ n�uαgs+)X��o4�͜K���6�o1g\cf��dv���4뀨���:��.���B��oh{m�L"L}ӣ��w^7��U�e3ƕ`�%ww�.��V��iE5�c�$kh7�,SG71��D\���[�>�݄�wu�R.�`LV	#,��
2���/��@fMf\��b�J.�[G��hVy��B�i-5`[@kN�n�vМ�q��і��5��um��*ܥ.�JN]�מ)K��ߗ��=�>
G����#V�R1�i[�]C�@&d]kl�y��U�@���@퇱������#�:9A �/ ��������N`	+,	A"*�"5��F�a)�@�� !����	# ��	2�NNAH���
)JǕ�$�qE��{![h�әv\#E�ՉJu"i�*: 4�'"q�סW��������M�N����X��:�)�80��ڶ&#
rCZ�Er�S�v9m����Ō8F@�N�!3����m��k��R�Z�`�(�V��-R�
*",�0�$UH��pc�Fh�B@��že��;����H�@��vXB��]XBLrB1&��a�P��X��V@�	�@:Q)�.5����D"*���D����TI�{,!2�P
tI���Hq!D%"D�\v�c�iI	��@8ĵ�CPb�ְ�$
Z���0��~�	�r�rhR��%�Y
R�4��f:efb��.���ג�tզc�E�؄bU�,L�
Gl��6�j�����J76jă�í��5��-��
��t����B�*i���ؠ,fkm&�у�].��2Z$В�D�IGBjJ
�e�hZA�j3@%�
�дvf&�,V�r#�a.��%��8��ИF�(K[5���`1�ԣ��LĄ���3�[-�d��B�4&����r�k��.il5St�U�9)H�F�5�GK�������7c78�ؕ)�\$��`�fv;��XE�B����)�*4-��mɑ��5ҡs�v�PZ�� U� �����c��(�e�-��Sb�R&ap�72閩5�u��
��#����i��j]��#I����76�P��hXd&n�`9���K���g���X�v�u�a�j�,���la5�p���\-tYW8��5�I�����-�@��=dV�:��ZSRb�n3E�k3NG^��B%0ˍ�u�"�-��B�bnl�*]-���`��ĸ�Y�z��06u�K֚�.D��ˢ���X�kw\��#��*MCA�ͬ�݅sp�t�+���8+�E�)�%�p�t֐٢��m,Q�j�1��tV��C&��a�j\��vÔ	�@b�I��s����5�l"Z9��HԤI��T�Z�2��օ�Kw!���jf�J�-ɓ$�0jᶽL�4��es�7b�)C;p��n�A�%�MZKCs�%.��7W�iSh���
�F�6�h��ZpJ��e�eMK��aP���MM�MK+H����F�Y���E�m�jKrp�a�+1���CWK[3%ŹP����gV�\���er*�e��uĢ�e���.�T�n�i�4��n�
����b_R"©n����uSlP5D�ݶ��KXʈQ׮�Lb	�4s�n�m�kZ�H�lLѹ�h4ћ=pP�X�Be*�y�х���"�ihmn�u�*�3hLX�̒�+t�B�: Ue[�)5����"��"��+�opVa�2�h63J�Ŭ3U����êX�0jE�WD\�0���ެ�k���+@ ��h�J�[*9Yv�n�aZˇ"6��~��?ʺ�JɻT0�U�_�$�]�"�/�	!�n��K�`�⾯G1\T��Q�H��Bi$Q��8)�(�DʿZ��.�$�a�L\3A����Gw�%���	$��swD�
mo��<{��,���%D��1ӦM$M�uv�D��}lu��d�[��К	$��]ش��&y-�2DH��*�[ћ�bv7
�����iy"�$^Iv󻰒$9�Mҝts��鄐� ſ���%��*���*G��Z{;|�}�h�'S�4�I'�wv��I��a�����Õ�P��2�WaPʺ���q����W��Y�nɒ���ƺ�0D��_��J��I ׾5sΐd�����	$^��2wЯe�]�Ŭt��~$��{d�L��u]]�dݪ�Z�Ip�?��ry���A�7-��7�šɍp`��X���� �2jk�X�m��P3r5�v�(�1B;c��lH��=�=���I'�~�*�$K�د֊FS��e���.��%1u�yE+]�J���?Z%y.�ܸ��,.̮u<xk�'D��$�;.���L�?5v���E��IQ%/���z:N��渢M��*	'5{�I�kۊ�y�W�ܺ0�c�[���- �O�$)!g�Pz��"F<�T�[���6N�λ7b(,sجZ)!�ȒFee�Zwf�Gh��̣vɵ��\ˊ��)�-��TcmE��
����;�@��I}z�^��BI;��~iL@��<�	����#VŚ��t�}��d'�z���$�I�;�Y'�0�m:�����s���	���m$y�M%uK;���K���-�ą)(��*ck"�I$;\��H%`�G�&Q�J�~*1���K�l"�̯Jp��h��~�_H¾Ж�g�W�,Ky�N9*
kgJ*ц�I��UV�pe}�{��Z��	 ������9�ЖI���w�R�Eݤd>���F��v�V$�ŕw6�D�\�A4���@y���B�W��Hb�UE!0+T# ���b�BR	��T�8yY�έ�D�C�i/$�7B)$�]��lȈ����Og�(M�U�&h�S3h��ZDR�9ٺ2���ToTh) K�q�<�Ф���g��ù衢MQ:7U5.쟉>�� �ZË���/���r��u`2yg���"�%����!4I~�^!-�ǔϔ4I$����I��ݢL��"���wt_� �6Z�j�B C�YT���D�;]�A$�;�8�p������%�]��$�۲T7��Z�J�B	^bU�D����F�$���H�y󪴗�K#���H�������#79.��f����a14��hj^��u��^�#�f�jVڋ=�g��.�Y��0,ÅLU�R��D\�j������#�䗏ﲄ�HU)���I��Ua~����I�~ܱ7/AM�`A���':���E$J=�����>�\�/{9v�Ey�W�RF]��
�A�������X+m(Gn���b�fv_��[8�Y)|��W��I&v�	$�J��ȻJ�ku8��*�PI��ǻ�	�a}���/�~5 ��:��d��ʱk=�$$��˕$��>�J6�Y7j�I4"���"�%��umش�I4�"������t-���$�K��l$qod_�#9�j��H��I��]l����U�� ,��"�oݷ! >�WCۏ)?��d�ێ}
�sB���D�h��j+A/>r(Rk��氩PB�:�̄��_G�lQ7�:IF��yfMo?���y��Wгٓf��`���ž8~ zYމ�3�F�e�w�x�\���4��ge1<'"��ɮ�5f�X�9��k�>���$7�ؽ����,Cuci.H�n�MW��X�)�v�5aIemɊ6mM �j�F�i䲄�3L� 1��5���t\R:��2`Q�Y��,�;[v{q�͕�h!#tA�%R
�jh)Ib2�2Mc��ZA�##jGs��+iF+lFͭc
F�Vf�Y��)+�h��p�չsZ����n�kKKT�ɐ��ŬX�Hf�Z"�t[���p ?~��5?��)��[�f�]�<�sD�	 �9КKsٍLEa�P�q݋D��k��B~v��o�*��_+|�!�D��u����ty%�v��m!��M$����z�l�0�y�H���Q-u��I$r(RA%���m�H�Ux��I-����C9Ț�KǧH��T�3��(�.k2���$�6V�?�RI$߶��I$������f}tPHx��*T���`ժV�$1gƮs��I$�n����N�XN��ۋ��H��M$�Ks�߭:�"EW�C��>#��2�s�Q��6v�Sl��{c��3X�_��z�"�$�T!����'�I>��?�$��=� �����.!.�z� �A30��*JF"&Ug�neѰ��8p�{�f�)F���9;�?������s��C�Y���Co�C���i{ih�y�b���`��=���ՄK�+��{����V}�_�H%�����K��~w`B�6�'c.ȍy�BU�(KЮ��K�!��ՇTH=�B~$��Om�糙{��$�.t"�H${9��芓^��D�D�^B�.W�}r�s�@I��H�@$��� Q��m�Q�$�}έ�$j�'�v�F��Ⅿt��j�����%��^ ����ŷV�$���;�Z)#����.NJ��q8��I��0�5H���[K�l����]L�v�)�����ϟw�ȵJդ�@�{�I$���>�~��m�7)tp�$�7V�I�ݒn�DZD�j�2���"�c����!fr:Q$��wv&"Idw8�If*���pfclG��Y�eIH�Dʼ�O�.ů�D/%�~ۛI���zH�����g�_L{>pD����eH)������K��Y���7ܵ�82b�jfr���q��ʙ�x�,z#�I��u��$���8�-J�A��1!L�զz�7S��T�����qIyY����m���utH���ķ"� 5�B~V���Tօ��HO�6�I&[�BRU����H�Q]�v%���(��Њ	g`�u"g�>~�ͨ߁a��Y
��c���y�)���m�Ѷ�טl��0L��o�/�f��9�*��i�n۟I8}���.P����Q$��؁�vl�EZHE(�R9�Q,�P�l�N}mu��	j�qV�+:C�Әce�ųю78Y���2LL�U���M�I$�'�j��$�Ay��)Ov��I8�qb�%\�EQ%���%tH������x�,���&�H$���M${9���P,���GX˟�Y�=���S��91C�t�ջ�ȡ����8�m\���qxCKlq�V���{T�?���G�K��b�U[��*���С0�z:h�h���ʨxȅ��q%��7`$�\[��_�>�݌~�^R��o���xt�wM	4�HU�[�{iV�l�`�D3��v�M�:��/��f�~�z���.�f�Ȃt�ȩI%��]Q<>1�C�g����Ġjݡ����h��&}&vv������J�9���i"P�Њ	�������9��Ƹ��*��mO�!��6U"�$"��4I {;\�M��"����9a���ɲZK�7B+�$��n�ҽ��H�))��'����J����Tw�5D�z���.��ލ�$ ;}�los�f{=����d�mp��IY��FJ>��! �3���u"N�s>�=E������@'��0'ĕw�4��6�xd������3H`��9C�N'Ǆ���K��ɹ�7�ǔ�샣kU{,�;����b�Nk��4lD �s^�L�;��QU�[^j�e�Q�h��+�m��J����:�t�]�����.�u:�3�8�X1׉G	v���lͩ`[j�iNX8�0i�i��ͩ�Z즰ָ�
�cwiKFV�qf⛌��K�Zـn��`a0�R��T��b�.[u��H\�iB�1��D��Yp�b-HS
�-GD��t����kqS2��6SQnn�di64��v
)�vKrئ[��h��	j9�?[.����@���9]
�I^�V-$�G�dՄ������=yAPI$�z����54��&`������
��Uu�U�j�W�$�Ixf�]�H�Z�&�d%���ɽ�$���]V~��������{$&�$�wd��V�yn�˱�Y�G�H�~�!�D��b�	��7vl�D����:ܜ���M�J�{V�PIysܛ�'��
��S��Ly%�v�ѻ��D�ILH6������ݚ�yT�X�#{�np;8�~�h�=��!���E�2���6e�����5��k*h��J%%�����mƎ�16B��2´U�����u�I�n�#�����H�캲BK99
��O_%Y'g�b���u�� ��K{�ѱ�%k������Dm��=����H��wq���v�A�l'+�J�A��(�8�]S9k*�q���J@�	M����V^�'�I��:��7�� ҫk���)$��ɻ	$���*�I��l���-��[�#u�� ��>�GOt�p�I&Ӑ��J�ez�t�ʪ��I �K�rh�s�HM$9N@�`���˜�̼J��^>ͲI#��� ?|}���I�G�߻�Q����lwĒ_��R���x�ٲ��"ܣbs��$���V-p�BQUاK�s͛�%MЊ	�g;�Z� J.N$!.T����a.8��u�\A-�U&�&е#�k)�2�>����)U�IV�a�/$�I<;U?� ��uV�8т2Y;�O��M���E|;U[$��]r�J��H���B~'����ų׵ui%䗵7B($�Ivs�1z��z���vgq�μi�j�,�h���%�ۼ�q��r���y�d���[����l�[����]�	Vե�[V��swy��/%���a
���܈=���d5���U�Me�5Ԑ��z���ȺQͫ:�E�1j��ټ9�|<���������ޱ1r�u��nL�(Kg�&�yl,[�o(^�����Hg&�ǐS�ݹ�y��٪S�������w�Uu,�+S$��6�t�U�50�P�+Պ��uy˲<�����s��]��@K+���Wן=M�g	$E�%��#*-Χ1��+.�"M���Ь-]��DFj���"�!Nix2��w6r��ƙ
5�\�����D֒�5�r�|���viu�c��j=�� |��f>�E���sI��8[�-^�2�q6�֍���U����Y��<̚M�ui��ɹ&�wӬ���뾮�-9�w;z�:�\7y��C�[��@Y���/�ow��X��b��y�aƷWuB�9�v��s�T�t��ķk9"�� ��W[f1��؝�Z�s�3��b���>�WD�P��I�}m-�k�S<����v(qf��f�[$k�ump� ��Vt��h���޲c�1��:hV�C��wFT�E{Yma���]ۥ�vr�77��&F���mJ���;��7�+���+u����`�{0;h�z�P��+%���;�}b�A��箹ճ��о��!�k8ۮ�:�鼈w%���N��p�y��!��}w�T�.��73���I�ON�V8̼��(��ΪXG^���N���,�'��D$*�Bs 	G"ȒMc:c��IN�������)$�k�f@�3���C�r ���ń� *�d�$DU� 7#!��h�45a
�jI�N��@�C��@��:�)�Uz# ��JA�JJ*� 
rR8��x�$I�f`���G���Q!u�bH�@�K	1"u��$�� 8H���X�R+IU�+��
�	m#T���҄R�^IKF�R����,P�[TR׭z�lx����� �Y,�����"��m[XR���!j��
�Z���Z<��{ՠrb��꼒��6@���+ؒ��)(KZ[��$��-l[D89"D��))) ���"������!m䤶��JJI@�8�,���\,��׹���u��c�xD��Z�D�W��I@��Ũ�,j�����q��Q���G����#�ҰO��������Gf��m�7�Q�Q���7���Gjh�Ÿ�Z�^��gqw�P�.-�ˢ���e3��՟��V*�{�|�x�A�Uu@��ĸ�-���C�1p�a�&�ph�޾�q<|�j�%���I��M��w��s��!���K!q��u}kZ$qA.7����ts�9���鸵e7吸_^y̦c��
�[�o'��W������kR2�QV�Lmnh;����-���������������d]�ݨ�Iz�9$<��q����t�y�`��q�l��ȗ�uߜ�f:����|⥿�ٚ(s�$�ρ�ڠO����Z�@�7u�1��a��K7}�9i�f2e���V��ڴ��9�4�ڮU�A���_rG��T�o���TyzϽ!qnXB��:�Ƣ�5�Qj5
}�
>�^�#z��ר�NXePZ�r�-�K���>�̱�w��-�'�N��3�q5mX��h[Vդ�{��uq��Kaq���	��y����\$s�\nˍŻ����]���Ք�[���}y�2�����,�䪕[	�����a��w���۽s����t��P޵�jm��ܶ��dK����sI��"\n-F�l+�9�U��v9�IOn���cq�Pn_:8�op'@��d�ڲ$�罹kM�$G��u�,>��UwP�}w�[5�R�1�s/
�� =�{�3�D���!�[V�w�s�N5mo5�/���LJ�kD���\n��w���w�QlB���@���z	��\���W�G>{�B��-�[�;���Z��\[������vn��R�7�����H��ş_�����?{�1/��W�؊�c��J]Fj�P�̴ҥL��vL0���U%���!������x��b�3�����|�q���p�w�YL�Qj5d.7���#���yﾻ*���yˣε�n.��qj�n-�\/�w�S3p�[�ד�˻�0�&f^��m8�FNwzۦ�ڶ�n8םy��\��/!�<����Z�E�r\:�9�ZL�qj5�.7��ȵ�ljڴ-�j�����������U��G�y��z��ɗ��ƭ��D�����u�t�Z�D��rH�-M0��.��7�:��3�W�����â\[����n�y�YL�Qj57�r����е��h��7����fX˻��Cq.o����εuw�;��<��.7�P�w��l���F�q.�}�9�8��\nˍŲ���s��7߷�s�o*5S�V�[t���s��'�K�h�gd����W�m���Hjf-���e��7�9�M�w��f�본f����!㋴�j�;����ḗ����n_9��8��7�q��cp��s���;�r�:��ޱY�t�@�1���ժ�UK�׮�u�7oAu:�a���G2�+㮵aα�N�5&q�t\��
��no���RJ�*�Y\a�V4\i��]��J�e9�+�-�B���Кj��R0F��a+-s`�[��[]B�X7#� ̺�e���'����s%H8R���K-&�9)Ǝ�k�[�y���Z��#��c�M��I]"ܮ�����3�͘$[1��M���t�[�:��%D԰hљ����0��AjhbȇX������qb�4T��6����ԮꍹU~y���\���U�~����q�u{���w�Qn鸜�s9&�s�QjY�p�<�3���E�os�&�O7Qn5^ș#���jY�r�r��H�"[V�v��qOm�Ļtq�'�M����jڱjй�u�s�����j5�r����9��\n7�\n%����8�Q�ys�[�1�9���j-n�>���sf;k�B|��$�ϼ��|~�m�0�2�|j��m�';�X�F��-�˥�y�|Ơ�M�n7b\����k߻&n����3��	>����2�×�k$�"�j�q��}}�q��ƭ��o��L31�/g���p����5}��o��u�:棨�]7�י�#��5�r�\[��s;��n\[����m�:Ǟs)��\17���|��l}i���X�F�kY�>��Y*���Qj�{ƣ�q���qj5�s)��~ѫ�y���s�Q;<��։E��Z�E���9�n.��qj�q�u~y̦&�n-�Y�O^�}�,�?�[��uD��A@�U*����qq�e��	��rb�`ܿ}�6�����,�׻�<�����CS1n7t��P�]�� �7.��lK��α��b;�Q�{�3���>Yq������Zƪ5P4��p.7��1��!��Ks�4U���rK���\J��V��}�Mq�D/A��� ���o,ЩI|-�bg���h1r%bȀF��ۙ�mHj2�e`3fol�J��;>�����������J���{X�B[���{����>��䞊s �a�q���\���%Ÿ\���:��M�f�n5.�Ɇ��ȣ�~�ܞ�O��>}FEt����fS�8֚����6�m��E���^s���w��n-F�sZ�[/�9^k�GvK���\n-�w�cqvVSqn5��&�ḷ7{���]�0�L��x�m<�����zh�3�t��D�J=��}�3N�h#T)B���0&��-D��̢��;���M>F��ut�!�kx�M�7�~�����[������V��6զ}�e���.��e�q;����8�S'Z�o�u����yٸ�F��5���.�\[����l�9ߝa7E����r�_��B�5Q��c�����������s��-uv-��UV#R�����{h�Z���@}}����f,�wx�iq�-Cz���@�n-F�\n79�X7�p.7�Q���~sZ$qR�pqɏ7�6Hf��^��~y�7{��մ�[���u�}a76�r���Z$y��wy��U��mϹ�q��������{ϕ��u�����n7b\ny�XMGP�K�Ũ�N�γ�G8F�p-���k͒�ֺ����;^�/}δ|'��ߺ��[\��.����\no�������ql� �ݪ��P>OR���7��p���^W�LXg �ڇsb/DW�n�]����wcj�e��{�"��yн�Dkf�6)�E������  ����� �z�TD�y�yLGLZ�Pj@ߞ���	"y�t]Hp�\1xfSQ9�����᩼>�w�;��\�Tj4ng}�1Q�$�#^u�5�D4�DG�Hw۲ ��⁝��ޏ�
#E�{�Q��Ԛ�ߤ�e�7&e���lJ����SbJ�5Q>��+hO~����;�e�)h��!���b&��� �~s9$]F��i��Q;���[M�C�N�N�ke�y�:͖�!Eڎڊ��f���kV�v4]�� ���}�ncs/��.y�h6�(����;�)B�h"P�;�����"s��Ľ��r�{��ڨ�J���u�h�Dh��=��̱�w�i.&�T<�{���E��S.�n{��=�U��}�u�h6ƂJ%Hw�}�4�)B���w�;��z�B��ġO��<�pcwy���pJ���SbjTJ����i#�� |��������wy����� �A����5�E�j-1��Ɠ�{������p�ykwW�h6��U��,���LR����� t���DJSA}߽�M�D�V~��!U�t�?��؉�H�G|�ۭW���̌6��X�I��@�B��ح��+��"7����j�M���B ��p=A�@箻�IDJ�G�g��C�x�b��&�n%C>g���L
�Dj'+�7�Ds%�fߟ$�x�(����-��B�QTy�9�5�SBTMמo)�$�o}}�D���~�����f�Pm(C;�]JA�	� Ku���D��C�v���U������0��G�I�k~kB�)B�)�=������TJM�~oI���P{9��{�:��+���f�淽d�ILj-1�s�u�i^y7�m�s3F�F4\���,�	/xVv�t������T�x"P�h"O��t�bH�����	#��,�@7�,� �L8s�(��B��Dh�ٞ{xY�2��7E�
{�w�6��Tj4{<�z��bD�����rϷ|�E���B�)�y�f�B�,C�߷�1�AWu�L�"Q���` ���:>׺HU7����Gȵ��0`jA$M�]�)��"T T�}y�d�vu~u�޻7�=�J��5_sx�6{����2\���ش����tJ$�U���rMP�<�<���������P_:� j	!�P(�\�5���P*@����"j%A������ή���̋󜳒!ԙ:����]�0X��,h�"��Ld8�M�T`2'1wfs�RUx�ƶ0��f]w��� �����tU��
]��(W�q[.V���``eL�j�����⸳B�՗+�u�q4IH[P�&��&(]@�(Ҥ2����%��Tu�F���GU��٥�Q%j4�����X�S�m�p�è��p��f��u�ôģ,҃,G���`FWUSY�a�&�1�*�c]�FZ��&+34��B�T��K-,v��m	Lj[�;h��n�m؛�l���ʙ�߄"x��Rb|xi��R�@�5��'<�k)qtF��G��ХA�y�3�ѭk��(S]�0w
B��;�}�QnƂ$���ؗm��ɛH���
x D�jϾ}�<�o�9�R�w~a�VЂTh��(�w�%��J�L
�L<��IQ��Ƣ�=��<�O!�:��jZ��_
2���f.�4cE���QiF�(��}���C�Q��F}�{�Wֳۚy�@�6 ��ϳ���ڨ����C�~�z���of{ۘ9�ww��-(S��p2�5���s=��CIZB����޺ɢ8�LjP���ȴ�ֈ�Y!�5����w|�|L�
P�C�g>��h"C�h�y�xe�w�l'+�o�Ц�#R��5Qjל�����W��Z�ߚ֎q9�V��z�\M*@�4î��H��E��Z�C�y��j��;��穾�>�f��v#��l��lmf-F��5��*7�m��K�ߟ>��!�q���t����]e.	�T�U���rCE	PIR}���M�D�]�WƓ��ϳ�����
`�
��<�H��Q(�Z�l}G3!.��Ǝ4Dߟohm) @D �,���lr�f��=�B�2L�99q�kf�_}������A���K���!�ff滬�C-�s�:�Ǚ�s3sZ���A�yy�'�V5R��H���b�m�bP���{�l�(eB�˷}����{��z��A��	�;!v�[�/��J�}��SbJ��D�~w�m� �&�;z�5����9}��)�9��C���Y$]F���Hy�����m{����-�.fb����fP�����ղG�$<@�ʠlQ4(RW7��i��-D���YK���U��g+[\A$[�y�"�Q��.`���^���"}�������TNu~g&����굝2	!����-ؔ)D��w �P�F�v�ި�mKֹ�|����e�K�6�[��qY]��h��6I1(-��.V�	\"��}�����r�0���_w|ޅ(R���Q9���Ҷ��Dh�����E�l>�]af����U�Y�E���O�gȔ-T���o�¶�@�k6=�L��2�� �'3~s)pI�:�+Ɍc{���C�(����<ߝ�J�kt';�oTZP��*!+_�����y��4-4F�}�x6?#���N��F��5�z�h��5��j'<�k&�����#�����i}_M�돢�7X�s���E ���P��2*m�yX�۬��Ŗ�c;o���vj�/�0M�#����6�uwNwU
�u�?{ޠ����h?h ġO7�p%��o���R��k�yYu/1��Lh@3~w��]s{��@n4Ũ���s���Q)�Q(�x�ZK��%A�A�w�9��/5�>y���N��i���L���m6�7�}}��o���7ܨ���yLA(�@<��I&'2��B^f��V�>x�B�m �m$�O|�w�-��Q%D%!��{�Fƴ�Ѿ��zvM}40�]���4rG�ԫBk�X���lXD�1�B�ݘTrT��tﾷ������iB��y��J��Qh�D��Y4�j5� ^��n�>�>#�F:���9Ǒ��|� �P�FR{��TZP����`�n]��į��7�J��F�־m���V��3���*4F��=�=ޒ���T�y��u�Dj.;��m�g�ml�(�;�S`�d�D���b�m�n��c�D���>�Z�h#�&w~�O=Ϲ9�N��9��YK����5�w�9�F��4s�����s2��h�>�\��oy�y�e���'ޓ�|7���m�J$@���A�4�x$�}�> ˸y�.���$�ϳl�N0����k�aL޽Oeeȁ��9��0���q��l���+l](�V.!.c8���o��r�w�DG����@���ڢ��A�}O����w�lM�o>��)B�ƪ%
~<�pؕ��
��5]�pq�%D���Iq5����C�s��"�5D��ZcP��� � ����Zc���z!�BeB��Kq7^2mupT�����B�+#X�.��W�����.cx\����A�Ƌ���-mĢT�@=��C�F4��D�����H]L�z1F��J���R��-@� }���BѺh�s���0�������ƈ�������D#Uz�:�{��q������k�$@�Ͻօ(R��}�@hx��;�<�
US因����ݍI�O<��rܻ�vdy��$�H$����ΰh��$h������_��}��:����i��Q(R�;��V�6���C�"b"$>��(�m��@{Q6*�vp��E$ʠ3��`�i�T��N{��bH�9���Qm}��=���N�|��D"ߞa���Dh�kݭ���d%Ӻ8�ƈ����J�E��Ny|�MGz���7&:���	'7��6�lcA�BC����p���2����5E���._��~��Ϻa��2� ��zN�������u.����x��v�L�ȇgDo���\�Kj���� ��\�-�:�(��9�u��T]AvEVNH/u��NW1ܼ-V��L+�H�R���l��eK{C;n�T�
��,F��s盼��ZVP�k�M�RdV������[H�l�f,�Cu�� Y�Q����o�uf�G6�d�D��;i���w�q�N�s�wG��jk��KKC�w&}q��$e���,Y�"��3,��'{���:�5y3�t��R2����r���U���-�cH5�e:���2��p+�J�ĺ�̘��{k���-=q���`s�lF�A�R�7;s�ej��n_?�ü4=܇9�[\섪v{�b6�#cF�}f�;`��m^n���3��s�D���ׯ%��ކ�+inu���ܜ�MhD��sM�Wa�ӓvڙ�<��N��+q�%�z�(l��7K���n7bʚ��'U��o\��ؗ��
MW
ǽ�+�/0Vm)�-���"^�:r�.������a�����(����̛���X��/nl\`���Ѳ�H ̝�3m��|��{R��B��E�9Q�|�L�W>0]dP�Ӛ]�[��*�Zoi�t*]p�6��:�p2�o���aήMv͙�F�Z�ܛE;�Ϭ!�vC��H7:S��5�{0v�W;{j7n4�j3&n�q��{��hiKQ������:�S�5mn�H+TԔ�U�D������X��NjE�$	H��aN�}�k��H�[�S�DTQam ���K���@��@�:5,�C�JP,UF�D#����u%PD�^� t��ֱY@�8�VR�p�.`�21�@�Q�^��H#,#^X�����#^�X����^��BPY-F B��=D�<sYN�AtI�$FVV=H���Ԉ�;�H�m�D�H�a%�Xw�cVP'���8�EbwB4�TH�y+�	Ia)*�2 $I�H�W���I��y�ו+)H<2[���Ū�e,�`�cD��" f[`�Qq%�2���?h�jO33q�	�c]��b�yЉaf�Kb�K1�R��r܅�t��\����A��m��K)� 3.l6bh�v%���a��Q&�ITK��X�ŵ�������ޛ�Y`ʳô��ehųE���̼�Vh�K��a���G	�+e`[uB39.:ł[�YBj���h���u�f���e&X�A��!�\:z��{�k��}_^��H@�C`SA�V�6!�׆W����lj�fm\9��1j�[���Kr�L�	 5-��:��]��ؙGhV	���g����6�4/=v�r:m�l�v����΍���Fgls��j[��ثؕ74Y,M4�]���
��KxNJJ��k
K��6kƦ!�̓��wr�Qٹ5�o=rK���f�خ���+�����IK(��Q�)tģl�v��� \jV�cH�:�2䘱�	B���ź:�H�$ЃRj:�C�b��hʑ��L�)�ԉ�)h��`�:��+#�i<��$XJ��6�[��a1�s�3��me)����ك`�J��t�&�\�@)��٤h�(\�a:��m��j�@���eSB�׋ɰ�֎L֡�b�6�Vݩ
�v�Q������PU��)-���Z��-rU�z�؛���P��k���f�M�& ��b��v��*J�R.mQ3U��X6$�lK�X�r:�d�R�&j�b�!��Lb&�r5+�ٸ֛��ٷ<ݑг,c-a�O�\g�-�J�%�X�tX,y�l��a0��	���hͦ��é�j�M.�7A2Rm�WW�a���J[p�X�:�f�
lv,�5`k.F�lM��a�����v���,�`Ɣc6��Y�ᴨ�c�fb3^Lc�-�R��UUEUG�l�&.v�D4�e�-��Z=T�1r�*�;k_����һ�}�dQ�4������"���%jf�X���y33�i�E+�e�]FbT��%�+�X�F	v{�Mtm�%�Iw��V۶�iB�E %u�Y�2dc�-��!@��,̸��i����X�	��Q�҅�U�ö1H�<K�Hmv��X��B2[��V���֘�u�A
A[40UPv��f&�P�Q����õ�l"Sk�qitV�\�a�Q������eK���o�&$��v�'@��wTj-C�y� �0j	"Ro�y�%��J��1|�nl3D7�:����E�Q��5�=� ���'���\���#��B�>��A�D$(���{�z_9�����F49��`M�D�!����1jA�3��r�w�p�T-��k��/�7.�r�h�D�z�x05�TZ#Q9�����"�5 �޷�o�35��Y�o�ڭ5�(�Cϻ��(X!���5E��kGo�2\�r���N	_w|�i׿:k�y���Z�E�s:�$A$JbTJ��w�%�$@�4C���E���^Vz����N�E��Djּ¶	�	\�h}����eM�A�4sW�2f �T%P��`ΨJ���W:浆�8�MI�7��؁'~_7���-@�@��y���!?��ʜ_A��	R	������JR����<�A��!��[A[�����϶��-Wl�9�%C]g���A��';�o&���F���<��5*!�<��{3��CȔ)�g0%
P�R_�sTc��$�s}Ol���/&h@*��Q�|DA���7���2��'�R�zZL�(Z�z�^� ���5�XL7���+{�u[�+x�+j�2n��A����b=9F�{� ���<��部$�H�z�y�&"se% �@���p�U��P�Z��w�4N�Ӵ�w��@�����˘\��vq��.w��m�Q$(������B��	G�"��Zz�m����?�`�'U�7��@��Q~y��H�o=�fb������64D���|�9��W��j�Q�s{�1(P6����4�n��F%C�{� �N����a�ڋ��H�&� 8���`�C֏��0��̗�@m����z���F���ΰh���M�Ѭ��j%D�W����MD�5�u�0f.��BеPj'�{��6�rM���ɞ���jhn,C�W�m.��f��b�����֐�ԕңmD���o���n]���T�F��ģ�B� �ᤡv�F4 }��dA$5�﫾N��TӞ"n��LA>���C�~��F���'���U�I���Pי�APjE�rp��zs��G�{��5 $@���5Ԩ$�STy�:��	*��°��f�e}��Ծ�{�xI�U�}%���y3@bu+y�p�l@�Jj�Q������m�#DJך��ޅ�N{G�v���f��h�7*��%o*Oj�[�/��u�Zn�o��(���qQBݙ�����h=5�jB�Q�k���s�\ODJ��4ÿ^��iB���յPj'ߍy�iy�/��s�3�h81���sA���,�}���3���T�@7��IB�h#)��Q�;� j	!�Q7����ƺֹ��yy���5 �������:��wX��#wy7E�m�'y�06!���k��O�g�}�{(aW���#�^	h�y�iB�lbQ*C�w�{�*Fr��5FƂ'5�������3�f��
î[9��F��� ֍�����+�����`6��ݟ�����0�l#Q��F�';�lJ�*%D9}�эh�]���v3��2͆`톼����5��Z#P�]���I�	����ے��s*lZ�h�o�	#��C�G�q���,D���#_�2��h"C����P���N_�sTbP����oz�4;��aȜ"TJ<φ�!�1x�[4����y�`5Ph TZcQ9^sy5�	 " +�6s{>���_�''s�G�XƂS�!�y�n�
�b����mNM���v��/&h�16%\��,���{�%�jq����rh��A�$�����1LJ�H(���"�b�ϬOR�Z�ad2�K�'O�8�h9i�P��WRbG`���F��+(�11s4�!�a�=/gX�Rﺒ�\��騾��Z�'?�W�p�3�{e���vqCl��^��� �	��9�9�0I3��.o��P[��'~��IB��������ڨ�(@C�}�J�#�?�����}�$�D�@���(��(M]s�]��P���1е�#������U�f�;������߸�TB5Q����w�cZJ�wϽѶ�lh>��{g�<�x��{���4�;���o߷�1�A����.�q���N��w�6E�>Dy}�f.g�Y�}9���������]G�ns��v��Nd���TDI3>A��\�A��"�.���v:�ex�	����I#��W�Ղ�3���5����`��r��� �F=uD�H;�%i�t�Ƞ�=�o�0�]�UiE[w�n������%V��CT-��dک�OsuD���gߕu%���B����Q���~�c��;ƛ���3o9]���ޭ	n��u"�������V(��$�5�3�6�n������{��SSv����MX��B�]Ii(?���m��VP��ӌGM	�5%f�$����X�ܬ��Lոv�j`�0�aH1��v�^���ѳ2�V����+�%C� �"节@�gJ�*��Uɡ���are���-�-�S��l�nй�uɍ��X��FX����e���:�`	J0��6%M��V�	�c�.����^�Zj˫��V�3`3,��av�+�ِ�E.B(��~����fPV������#-��sD���T��s���(�dg��箭��H���D�N��&�a�;ղH#��}��s�`�X�����W(J��R���v�M���*��9���v��r��,	�TCݑ�L}� 4�#wh�4Ǝ��^�+��PRj` W������K��nʉ�f%@}�z��:� ��>Z� 4g��v
LO+>���~T���H��(������އ��6Xᘤ�ِ�MX��K)��J��S��6[��Uv-XJ�x�Z�B�;�>��A�!�_���q������x2�����Z|~�_������p�,l*�5�ېz�����̋THp��[�O��5�������86��vl�"�.�e��{����n~�7{&�$��}q@����=�[@5#��6�v�����lh ���uH�ܹɳ� �߹�N/��T���""HAZ�+�8���/����]'�Ǯ� -�H��κd՜���KpAۧT}�	p%DD�S��v��^s�3�^��W��7"gn��;�I#s�P7;���������?(z�}���#��7���x,[�qs��e���s��ə�x��~�������A%��� ��uF�Z�+&��Fn� 
ӛ-�
��Uv-XJ�m߹�V���}��5�>$�n�Q��4	"�3c�N<�%�ޏ_�Z���V��~�� {��@�-�gشG'�At/�3��=���w���+��b�����`�p���\��X�f0�N��� �G���su�p��_�EK����s����oγV�X��v����g)2y�<+�+ē��
� �<�ۊ�B���p�j���J�	+�=�7@|*{q������c#�F�T�+ē��uD�sʭ{�{��A�	-��%�\a2�fE�kmCH���lk�ņ(ʠ��}������eۯI� �r+Ă{�PT,�0:�nOn$��t+�8(A'D��|n�����\1�C6�����]���$�<�@�ͣ���Df_F�p9��4�صajտ��7@
�v'�J~�eՍ��\a$�k�$sʢV�&��Z�^p�2�~������@x�޺"�u��?w����IB{�U�� l�\����}l��Xx.cUۉ�v$��h��m�����E����;�M��?�����z,�������R�"��5��k> h��ҷ&�F����(�κ	"�u��mWϏ�}ߑr&��RS�vm��U�K�I�Ao7j5
�f8U|��x��*���}>u��;c�� ��-�V�gn�J�����gEC�$�&"fD���,���O!��\i��� �m��E��G�^��Zgyt=<<�N�ԍ���P|����RH�=�oo,n�	�{s��)lVxҫ��`%i+t�����}�Y>ыz�����g�Rd����o�94���h��".ա3�C�hU 7;S�qu���t�M�w	'��Q�<#�<���d@q�\��{7 ���D�q�q�'�@�(9s1� F��St�ڇ��ne8��WA]������z�^!-�]��>����,��JZ� ��֡e��ƃkf�6���qa��+�M��B	�l����T�\�&�:��Saj�z�5Y�ie�B�iaf��Ô�ݵ�(g���K�����+W]�i�I�$+�@h�萂Vˍ���e��a���11aww!(���,���V���[��̳5�#2�M]��#��&k�m��� TG�?�o��d�TB���W�Q$:H��L}��:Cٍ�j5C��~�;캊��TmI$�}���Xۭ�-z���b� �θ�I���l���.�2�]+I*I|>���� �j`}��j��}Q�7��A8�n(��hzpW��R6���H���X�o�`o�� p�t
'���H$�<�/Z��X
��6ݿ��V�D��E%m߹���ٹ^;զ�nB���=����uA��o��R�
� ʉ��l@*䎋��X�K��å��##Vl1��r�����ٕ�&$��eАK��P�Cʯ�%��+�x�7�'�P�j�"��*={t(��͏���59�_Ԇ��g!��kE�{S�P����XKՕ��k.�!��u�G��]�BU�EH�Y�D�z��7]�<<<<�����@Q�H�f.��%4���a :���*)I$����lSۍ� z��I����R�o!�{��	y�z���숙��$E��.�b���^'��ׁ 	����M��UݓךO��S/S��yiP_	��4g��e�T�"4�=T(�^vH�E��0�����h�Jo�������"A*��M�&)4���b��y�4G�s��G�?_θ�G5X��I�eQ"�u���^�B0GUr�@o�����V
��)Z�~wW�G��].w&(P��?�����Y��$��-oo
�\�"=*��w�B� ���H&�~��e�x���}�韔H�R�귶C&h�ɼyw���ҩ�J�=�P˽̔S���cv%L�z.oq:���+^S��j�4�D6��X6e�W����m"m^f���V��B�33S�nP�� h�}��؎�r�
癴'Y���7}+�t������R�^7�*&vG�4�h!pk+紵�����m]Vy���vHn�1Q5�W��CQ��	:��YpM/$��eG*��\�e�YA�:��E��Z�].�F�P[����U��/h�ugv�!��w�*�M�b���SL�+z�:�T��/���V��� ��-��{�ٓ4��Uʛ����j�nK���Rk�n�l��x"xs',\@���mV���:˜ك
�X��ܯ(*H�Rd�wq#vPyCwtk5ےmW��Rs�� ��&�bS���u�-�*	�ʬM�As��È��5�ddР�ԋb3e�lL�3j��۶y�շ�5)VA
��)؏K_f�o��W+]��:��&:�j��h�4��RH��B���t��NΓ�,3�eL�s]dکՓ-�lf�!���L�qgq��a�Q�\�b� �G�H�j�NW3���u|����oM㕗G3Q8��v�t�ޥZx�l8彺��#�\��
�+4}5����޾$�{�0]h�9���K:�ث�ҳwd�C6���խ��0�������9~��� �A�Pⴒ�̢@!+��X��X̽(�D���NQ!%:�Y�E@�(�+ւ�RZrb�=N�z�Z�P�F8��y�)1�P�AB# F�aI2��'#D�bHE�HR<R�c@��JY` W� � R���W��X�J ��Pzb�F1��dC��z��H��"V ^	8'"��N@�#8�ȠA[e' rа��J�''R%���H!�R5�Ae�K���8����e9��R��#9z Q:y�%�KZ'D����q��!d8!$T�# \�QL@�U! �U ����� IV�F!V�����F�$!*��k- �=#�w1y�@^N��B�y$d�Ԁ�Q$ᬥ%)Iͷ�ğ���w�7�}��|I���T����qD�jB[�ȕb�IOsk7�3���i�K`U������n�`t�.s��V ����� �O[�$o9�x͕�}�,k���O�7qD�w9�\�ꉌ!���F��s`��5+�6�
�h.���.�H�0bg�����
|X�� ���Q��"#B���X^5T�
��≴�ylZ�J�%h��e��׾�G�c̑�Ľ˻"� ��΅w	�S)�=�n`����UAJ�|��(��O��,�ݫ8^Ru�9L�մ�G�9��Lj�"=*���Ѯ��<V�;ez �ۡD��o|�fگ��A����;-����u��on�vX��W@ÒYx��=�~>�qrC*f(�ˌ��'������":+~�J��V�$���� ��5��>�i�ГD��j�'���Ou��8e��)�������߯��hi���6�&f\Tq���mbp�Y�vJ�Q��T_߾�����,�_~��=��\�$�uGݻ�s�ƕ<�Z�	-�����S2�݃\ꀠ^�owk���	�� ��t(�0#�\_`u�+:��(Rf`L�Jݜ ���	��=�ԩ�	%���
��5��x;U�Ti!(x�0�e٢v3)��kĀI-��A>�����p�3���1y�D�B��D���IZ�c�Cp��k�Iyn�����oc�@�/c�Q���;��_C�b�ȗ��f�E��3��z�)�Z��ݼ�F���w�;�Y�[�Z�;6<o"���mF'M;�jd}c����#�ADv��m~�\'���f�q+L0��Y���E�JX-"[�cb�V�\��U�a���mu���ҰB0�]2Fg\V�ЎR��8Jf���^�L���&��h0�`kiuղ�f�G��l`-j�S�:VU�aI�6;i��j�֍��Yk�,�]4 �}�v��sq��*1-R̬�#i*�@i��5�q�؃��Z�)�.[�� ���E�D����y?��媻B�IO�l��	٭�<|�3�Wö��k�׭�� ����P�)�B"H"�t���9|
��>e�H�sq�M�u*�����OlGX ��Xt<�IQ_	�5Lo��b��<ݗ{f�g �y�(}}HU��FQ���WI+ܫ��f�pfvP��F� 7J� �=΄&�Ls�@�b�ɛ=
$	D̚`�Y�� �nh�eF�\�R6�5�:�?���k��O�>y�g�ǿ�>).��3b�%�,�I����Hn�[h�P�#��������Kc������t(�㸶�<oy��t��x�<�@�V��.�������JO��7@Q�R՘���#E��s��aDl�h}8:�BxL�W�z�e*٬���g, @�˱��M�Z�z��>A��T8�(�����In��_���{��ϗօ|� �/�W�Mݙ�b�m� �ҍ������ЀA�nhM�9�e#��o�M�B��=�N��dQ����p?N��l��	.�b�N�	��(z�x����c�Q�ؤ���������k�S��C��5�<T	�n����N&��.�#
�鉒J�"A�d�1v[@����m	ٶe�[��W����)6M��řPI���4��ni-ȗ�-�ԛ<�Ꝩ��/_k�SU.)
A�(�==0 ��3[6�0ٚX�Y�u@�su�񳹜���w4����,��I)+ϣu@|
��t� n��|v���U�"��

�����p��ky�Œ���0*jv7Kȣt�lD�٧��sq�^��Q���{�Mt���^��4hZ{��hӝ�D�ɒ�w���t��ơ�n�zh�vH{Ψ	��u���7S�H��OUmW���D zJIQ_	*��Θ���ue� �管��
�$�7T��֨��rڵެ}\O�%��3D��90��Nβ�),�%����#hD�	-�����a$i%~��_  ��tA$��Z��n�����K�t(��)tM����c�p:~��lI!溢I���^$����I��`I�m+
���Q0t�l_�п��;8�-
��7|O�9�רoWZtr��"�H$��7�7[sB�׼����_� �]PI�7�ֽ@_s���^��G�emŸ
!��6�Ɂ/�>�2��GU�U��eKҮ[S;��q�Z�C�oy���
���8���F?�~$��^�H"5J�"$�+��\�G�3�ڮȷ.$�H}�dQ7��(�����(���ьe8�mMA���*z�݌�˷:W�u^�fZ��������
|_Ʋz�Az��H�Ϊ\wd"g|<��t;��`PS�.�7V�($���n��߳��Rۗ5�B�fzl�'׹�^��AW}0�p�=�jPD��{�3�û50	��o_J�έj�(�()���6w��V!*��m�\@�،�-��"F�9�A=����w���>s3Ɖ����B	$��q�>=���Y���9��RHx�$ێ�|w;*���F{���5�XRZ���;WD���Z�o���Kji2�.!�Ь����R�(]��告�Dui� Nf�z�럕e��u,Ŷᐹ&D�-�:�an*��,�%�%�.��.&êQ4H�j5,]�m��3]����(��]����ʜj� �J`4m,p[��X��#k�ڍp�8��e��æ;���Zօ�]XA��]e�"m.��S2�k6\J�#�R�h�ԍ
�N6F���SPڑ�BZ�����t�c]�6�T�]�5�Ԧ੮+����4��TϾ~��y�h��.3��&�6h���� �Kw[1"o�O�f�$+�H \�3!O�٨�^�y��<�n�*� �f�H��_y9ó�k=�%P��� ]XT��1Uj�$�וG�i�F$gF�xE���f�P���S����6�����Tv���C����S�	1��@��yN���,G�b��eP��u@Rw���2$��*=�u4�y��r+�Gq��M���r��ޜ4(�so���~�O1��z��dK��,"q��U[t,ݫ{�w6赻ՕH�*��ڱt/�R	$��� 
�3��@|��C�g��8Tn�C�dסl�DR�� ��u���I?;3e�?��4�t��a˨U>SfL��9/�u��K����Ðq���&]"��ͦ�fS���CuϿxx{�Ϭsw(W���a�tį\F���1�.J���Ƅ�s���"	0.��)o���;��§y``��n���B���"�2G*�c�� y-t�P��Og9Y3�M�Sjv~H���f��w���6���� W��L5��Y�4���D�C�4 �Ψ����A�Sվ翷(3�#0h���i[.5U���� �&�Q�>����ʷ;y/Ͽ=���Y�leI ��Ψ�m9I�#je��^�Xs��|����^����Bڵ�:I"�N$��u^$�$%�n����F�\�B"H>s��"��>����ԶՄ+��<�r�v�>��|�m��-���r�]g�T%��K4�y*��Z�G˲}�i���s�U����{����xxf�4oK4	�|�P��( \�3!O�ߍG3��Gb��V�$�/�Ψ	�����0s�m�^E�����`P[�"��D+)+n���H�y39�2�ފ�^'��n�gd��nC���s���m#I#h�)Y��6D��E�f��K�!���#ŋ2�-������l+}����^�t ;'�wc��}:������`P���i�_XUj��D׹L��8.E�v�R�K�`�<_s�@��}^�H�ܱ�]�OW����37~}#`P	���(qW�[�跏���sD�|{/��]06L!$E���]�33>Y�#�>$���|��(�/���֟�!�{��WR�oI��\ݪF�� y���m?�*c��(-`,sM�a	����!��H�fB'�z�� ��&��TO�GiA�f&DO��Y�H/��!��2��0�eh$�ڢI �[���;�
�G�(k֋3�ns��җeb[i��<Ꙁ�(�����l�&]�e����
�����J��o���
x�Z	�tK�� �w/�Q43� �
����2�wٸ<�a��I 7n�<l�`�:�YLZ��%bz��j��D�����t�P^�ڵ�Q�J�  	���P�������vE�|��J{�NO ůP&nn��I-gd
�:w�%Ry�O㓷TLl�$��0�D�Ex�t'י�DBވ��N"B�U�s�$���s��N��ߠN���]��8{i��X&m<4r��r��j,R1L���j>]�Y�+ӗ�0�/� P�;8�n�˽S!@�f%fAJ��xy�^��H0X�jkl�ֽٸ�¡O0�{�e+��v�r��h���nf�Õ�`6:�db�t֛t35���S*�:	�<�x��M�qd�
�n_U�f*N��.g@H�_HM����ޖ�����Jm�9��W�6V�з��T�W�ԭqW��JB��%=l�4��/c
�z���G)D�����quq����z�Q4���o��H�u�O�{n���u���S��#�W����8��X
,ز�ޱ}�o8_6�E|���8��0ة���ֶLT6Y������2��պ��N��n��.���F�B[�{2��:�;��Yڂ��w�e�Ct����s�ٶ+q�`���tf$��5���QY���E�=B��YƁ�w��fs��o݊G#�1�m���(���Y�sC�W��wu�}.�;��"��-r�"ؗa*^��	vd��W�Ά�\�@WD��\�:[�5B�70�"s sX{>fX�WHcX�T~�E �-DХn�n�r��S[m�;Eh�|��}Յ��wr��J����9�˞���uGʎ��,�IX�BvEm����J���ֺ�tU 	n�O�O��۫+j����&�˭ [Yf��V���~UP%dK�N��#z�c�*ѕEJ��2���H� XסC��H����ZF�9� l��-:�`%� B$xNB�	 9�
U�K*�$`�z��;V���e*�2�--���,��������JqX���6��' �@��K�R�r��h� EE�[Iu��:S�� ��u$��	 cU�a)�+��Ҍ ���@�NN��V،Y��sd��gP��D�"@b�ra�cR1�شZI ���APPQ�IN�XBX</D葋9�P%$s�X��V3�8 A����R$d0�<�)@�aG�BU࠰ $AE��J)el"$,�<����������1A�a��m<��@}.&�+[�ЄԎ���t��.̖��$�f�*��uE�!�,b�Q��B��$)�f4��G.�th2��F6�-`M�(.{Y�&�Cm{k7#����p]�uƂA�A��MG$P���\�ʛ��6�i�x4
T"�����Ŏ63�ʖ�,Ԅ�^t��f͝�%3�`HF99u���M���lH�[�գ�e���^0����P!5�Lhg���$5��ݴ������Q��ģX[��Զ$� Elԥڕ�0mlح�P!�X�6���2��*]�uis��Kr�.�%�Mc�-�y��7�a(��Sۣ*ъ���qv�6$9�hE�c�%�¶�;5#az�"�BD�ZK�A���u��ҷ9�&�@R�M�:��Źf�CL�	���u��3f*WC"]�����66�IF]�a(2�˥P�u*k��p�hl�l��VfÞjdzY����l116�b�G[��.�5�+a�-�,X��e�ؙa���S:V�I�B�]G�Ye����2���خi	��9�q�`�K4ˇ2�km�!,v�E�R�պf1�m�d��t
��:�L;mn%k6�@�ՀB�]�n�<����)X�[1=��j:ͳ+�2M��!Ը�[fJ�:ݲ���LQTh����\�2����C��0��-F�[BP��
nL]1J�kE�q�������+j���KXl[�h3u2v��B��,Z�jZW]�G%�9)2���S�,I�6�ژ��	v���Ĩ2���&p�
mJ�"ε��2Ẹ�-��k�*�1)r�d+j[W\����a��]sP�Ae�@uG��r�a2�
�"f9p�*�����e�e0��8���bט���N���Z;l}t�����@1�i��V�J/e�,��ue��!��f#̰y�f���GL�Ycvяm����Va��,�i=3ؤ��ٖTl fm�!�%`Mf.c��F���xF��e�u���\�`cv#%](�1�"lqp�6)��fZ ��.T�mh9Èb;-JD��ᔎ5ښ R�,��\�4ʐ���1`�M*���pؐYs[�,����e��h��.�n��n����}#2���|�����F�E�y^�	�:h�rK
"�GU
���W�3̱ �� �D�ħӞ'ƵFwa����*s��@�����F�uy�}��F����N���HD�H9T�cD|{q�x��y���]�o�W<�$�fy��]��)A*(�=������'*H'ā��B�'��v�CqT!�]�t���<�ן�.��������񿀠@7��V�flL�J��%�.(H}�TI'����K�*GH�|`��/IL[\�ΤΨ.֌aƅ܍�n ڥ�����W��OɄ"$�8٧����d�A��#���j��\�����ɘ�>7f����z1ϗ�=[�+)�����y���!7S�]�S'��jS%X�-�Y�Y*حڗr��21hAus)�ijM_���fG���t�>��Р@2Q4� �>���gt�aB�f"fb���P��{[�D�F;�N;ʊ�� �����*�g��I��H$�m$%�g��YfM�M�l�$���x���4fm0LC��5:�EwʂAR(J�n]z�:s����Ϩ�sD��P'vE��{b��e��AHē��l;l2�P�յu.,�E�����n�`�]����qq/�$DL��M��	 �k�(����"��j!�7^]}TH!b6"CD�A����8x^��ݗa���/��GvE����{�|
��\����L�nר�Ig�T�O�=s��`m��X������\��R��m�Vv�g!$�r�RH5�G�hJRosC`�>v;G���)��JY`�aG}ײ����z(F���5�`���Y����Xܹ��y�l��!��q�b���sb��p�K ���3m���>�Mz鏓��H%AP6�P#ٗ��j߄w�^L�Y�@��)�o[�!���Κ:r�Vu�o���b�6-�Us��X�Xe; �n��kl4bCrܑ�#e]���7ʑER*�&�G�p�ƀ�>�i��V��[�7��Xs��k����>�I9�x�|� �K���VS��� Q=��D8(e�3Yt �ɣ� ��""H"�t�8�I�Α^$��3N��y}y��sn7Ăw3��!E�@�Jҫ_	>��|�/�_M<��*���w1�H�����q�C(wU��#w.���d��Pǅ@�%�&u�]^�NBuV���d(N+���4l8I÷	�gљ�9V2�G���@��� ��Uл��%i+����
�q�s���z_�.܊��:���Oge�rm}���y�<���IU�r�nQ��T(H��[22�bG7Y�%���E-������m$��hN�9�I �nvU˶���9�b�v�������7ʑER*�%�vF٢�A����v�O�9��D��"�����c�����p5���]���<n�3��I�7���A\�_d�=��D�|{;(Qى��$�I�fؒ�G\�zѢ	a��H=�*�ý��`�d��O��/ѷ@|nW/�ZUk�%z��A%�yv���a���/��.@���t ��e����ty+����a���á��ǵ�Zsz��I&��G)e���=\{<��셓�6�˾��xw$^Z!�������&f�@�M
 @�ښ�$�m�1׊Em%�[3-��b8)�J]��k�2v[.�f�X0���rfTҽ�-��3jl��/�K��S�A*���gL�$.�
�@�]��¬f�e54�6f��&Ó�%��2[a�Һ�@n��oY�Xd���B0�iK��n!�*b�R�=���nu5�%YEvZL틜m%� �	�5ZM4�M�+��:���������Z�31)��I ��(�|HŽp�f+#�R� I6�>ݏ�n�jB�
�6���cB��+�ZzB������ٽ�@�O�w\Q�k8.DN�e=9w:$)��J�����:�I ��B�E�_�{��1w\Q5;^��Q���JJ�<ohe�뽶+Ҙ/y��<3e�$��U�0��y淀c��/wm����D���j��9��=ie��ڪ����>%��$��O��ײ��ϴ����MŖV�5��؏����;'d���m�D������_��D=~�K�����Y�t�I"�:�b�zѥLW:n��bt=�iP��`%i+t^���?ɯ�����f���]cpĠ�T�k1m!�qgkF��M�Sӛ,:���+5$�U�a����/��E�X�&C������D��,[yB9�����^W��s_P$?���g�@�ڗd��s�/�G��c�8,����'��4���y����!�I���T��؟§�����U��Z��cӣ�>\ڂ�}뎨�I�:��#��۲6��t��d��?r�x��|+��I����,���~��˛�8iNho:EA�n�vy�}������o����;Rd%ث�4�Iv�ͤ%-.hj�p��\����Ͼ5�F4,�����͚$Gst7oz��J�r�M�#w6�����LLD���];!f2���jN�y@�5��{��@�&����r����P��`Z���{͏���Dw������ld�_}>Ǒ�4�C���+� 뮑qnt�Ƹ�X��;?nLݳ�0L]x5�C��;�'������/�j�$����E�2g)������{�/^'����QE=��L=�v���޽[��m�����YJ����:3���U�;w�3֠����jA�����2���k���<�j5ԩ�&l3�1�*82f�T�.G6� �f��U���
��m%���n��;u������!�]�#�_T��9��;�����0��"LD�E�5�^�[�k�]�6I$�k�� �]JI�DV��˸�^�h��Q ՚�٢Ag�����5z'�d:��${������+�bA���bbf"���CmH�gpe�O��]
��n(�}�?��/UL�~�6���e�?�[�,˰��S��on��|�9��H��ͻ��h���Ȩ�4FmfL�zi`Ģ�5�ר7E5�'p?ʣ>N�_d��~�s2HIyy�)����٩�����0����:>�����Ʌ��Õ7���ڲ�*���@���b�Q����f��
����ݞGf��y������ᷗTA'���>�{�U�1B�:���n�"�����P�I��Ej��i�1𴔛�ЩB����W�F�����.���&,�wI�Z3��0b��7�b���D�����+O9�ᥧ��/���x�Sk>3��А{<� �J�u$�����^�@���LX����73���s�++gE���فx�}�F�bA��"bf"�=�P=�С�MEC{���آA׎kĒ{9�����ߢU��������`�σH�Y633?>4������CH�����-��e��(��,t�W�u�cd�U�.z�n��@�p��c�7��8�ĈS�$I�.F�Ȍ&�nm��H[��clx8�Gg۵�LZ�5ъ]��F�f��� ͺZmJ��.ΚƎ��m��`�1.h:嚒���En̶��j�f�.KQ-��i\a.F����V8eMG[�-"p�K�uVǬ�	�
4һ9
����h�qLcJTڌRW�v�u%�u�����ʁ� Ѕ�ud`�ı,q���v#!s0��h?>O��-Wm6&&�5w����wq�I�s�QˁK#���5i�K��5��-) ��V�"Gm�D��u�.㮡���4}�Ψ0Y�c���������]"��i)S���đy�h����ç�Z���P$=ͪ��s�������� �:z�@�ݴ����Eؘ ��o�(`�����'b�c^&]�P*(�O����8��������)J{��'�q2@$��+��_M�o����"�(ʔ��ZJ�ї�]��]kM,G�S0E���b"D����Q�T	$�$P5��O�zT�i�j��� +��t�'S9 �Q$�V�d�u�����, +��73%�9d�+pf��V��"U0\lV۲Q��2�Inmɨ��*�kX����a�{���9��'7r�x�_�^#��輸!�+�yz
�/JH+�U��{r� ��u�k�DУ���l�A��7@
��<�M���A hZJ{�Zz[e�a9h�'!��I��h�}��Z���R3�mm
""4��a2�$��lQ�&�:hs"�NM�����|w��	��ίh��ꩾ���F���]6���3;,�3c�.��l`S��M�=��R$L��!��31���ڢ ���I�fuQ�(dI�D`�ݓtn�L}�iP7j�Z��۽�`P�IG^D�*7\(����vgP�&��T�۬U'Y�T�"I%+RP�'/��V� }����J癨�~�o�w���wXM��i9�ŗ<�Y���qе�9tl���3�&-B���X�'a�f27x冲��td-|�e�t��Np|���7���,&#�Duq׫�M�->Stا)0�wom�Y���cP�뀱ʋ�he�"�N�A�K�̛�fІ�u��^ۺ��q�`�Զ^��j9�
��8m���R�3��H��6eRz����#!��V�Cڥ�Ē�����;җg`���J�z73v�^ñ*۹;�{:_fl@��KklVuI�m�q�7_=�F�5���r�6fYFY�Q��P��+�$���e�6���n��O+*'Ã��W=�Σ�7_p?����V��Vݕ6T+�ݭN�*F���H�~�!������U�����3��q��akV���:d�k�����n�!O9���Z��� ��S5�HK�ϲ�"����
�Z�r �y���rˊR�c5ȷ���ǣ(添�Z��v^<H�qWXgcC��,>q�jX��ܖ�P��[L��$c����X�{�w�ڗ�e���?K
����걋o��mlh�5 �������7�{��a�Ѝ�8Cu�9j�g���oF���u��S���7$P�

��A��on1-���!ĖQ�v�v����u���g+�/����).�XG1�cAU�'�B>*���+��ؠ*�(��)��� �G����#�IlPŗ� ��%�	��K��+ W�ŋa�&"B�z� �*B,Vք�8F��L�����D�%��qzԳ4��@��术 0I���3�TE�I[DHA��ā	b<� ��1p<r<D8VD�l�Ǖ"0G���ʜ�$ ��!$`���C�9 E�rA:b��;�^9Y�yH�8�a#�$���RFAX$DEUQiEH�HABE��EF#))B
B H	rJ�����k
��(A�e�� J�����QW� HH@�$��D��y! ��c�8J3� 
��8��� �*BpFSEG>�C��z$����1�BO[���E��Z�j�%��d�P��G� +ֱ: {sS� �{}�k�+ǡ6�<�eg�P�&�M�]t-Q�i)>ެ�y�^�|kY�	;۳D�:�U{�y�n��r�x��L����V�5��ɵ��MMa�[+���K[tk��ߟ|�.�$+6��$�f�H'�e��� ��u��$����
7�O��U����@���tssS~)96��s�������:�ߊ-��P��W@ݪ6��t�y� ��N���߳ܮ�6���N�}��0�L�iI)Z�Q��,ӫǜD˺y��ݳ@��ɢ9ݓ�>���6GZ���-�]ڳˈ8�:�WIe�M9]�:�/o\�Tw��6�1f��piT�ٽs+����/����\���Z�A�dL}��n:��b2�"b.5��{B�O����x���ޞWw����/�f��d*�@Ҡ��y�9q�L,Ɇ�"2�F�i(s��أ�r����M�њQ_^}������� |3���>��S�wW'U�ר�G���TD�E7���A�!GP�q3D�{9�I�b�ܤ�������~ﶭ%v�Pw�t�y�@Q�w#eسW'��I��T'��d� �2���HF�SA��-��"�%�B\ʰ({W&>�� w��/��m]�]0�f�QH�	)Z�Q��D>r!�:��2L�A ��& �ظK�S9@6�Nem�y���L�LDf��73��#<��#I��{<�@{3�`ds��6��tA�R�`4!
Uy�5���&��=��39A��F��UԎ#l#X��F�eh��D�UIqU)�k��kBۉb�k(��hds��;fWiJ��ѡZ)r�B�u�ت��b�+�&�5��t��������]�-Ȁ�ˣ3�nDn�&�!���D�� ,ԩ�`�lu��,iց�F����ζ���M���Z7[��ա�V'���,��j0%�vu����eژCWX`��i3��p&n�F[��J�ܻ$`������1���˯Q�$��B�$�Y�UO��0\ݱ^>8�&�&��{�ѵF�����7B�Es��Y��t &�/����?��]�KA��ݑ�@Q��� �nۡDr��9��{&�:��$���h}w�U�}QV��y��������1�(!����Hٜ����^$��u��"�h�;g��$�z(ĂbbJ��	�ꢢN�rTN, zdL
�7��(��n�w�٦5��vz���B��
�v)$��q�Hb�֑tn��hԅ��PHZ��R���E"�$�jxQ�c�A��4M$�����ʎ��Ǜ�yh V�y�)��v��Z�j�%�=���;7�$�h� B�:6]Z�Xh]!w������{&0N�쇁&�̑Fe�^b!ҍ���L�!ʇ&�{��<ŗ�T��s��Iz�̌>ϝ
�[�jsr�{8�6o��E:Dt mQ�i)��Tƃ��������}�.3�.G�6�đ�νQ�PAbTD�@��J2��^�o�7w�@�^�sD�O�{� �����d�D�P�-��31�bz5����P��+:q�n몁��P$����x��.�w~y��'�)��V�L�u��t���B��e�6�r�n,n��T��NwX�B@V�^���LV湠H!�\��{�O/dT��U���풫;�DR���ىК�mZ���L�Wq:�7���{�0(s�{l�F<��wj�դ�R$W�5� ��J�	"�j�a�������Y�8�u!�w�ڸ mM��ԶS��}]�|���<*`�bܜVr���w���Vd7c</71P��ڪ�F�΅H?��߱:�|Ȯ��4-%'/c�~�7G�t�>@���D����{Mf��	6�ר�A<�DA�*"H"�u��r����*�cx�}�D�G=�L
��u2�8*��1��$��b��R1��RR�{�ư���v4:����D`h��k���s13���� ���P>'�}�@���ی<�O){:?�P��N�����&&$�.�p����Q�oZ���@�O��0 ��tĂߧ����m���E�$�j|=&0�g�0>9Y]���΃�Ή�N�:�RwK�wj�V�$h�u�:�X��&��̪$�t(�����tJ�v��a��8�yA'2a�� ;ƩAԝlf�Uj<.�=��Q�<!ST�r��ws3���!�>�	;�mBk,�j�I?yE[B��[�^��9)���r{&�>'{6�@;�Х���[���O����_օ�*Ҳ���A���8�nqnt"iq��6��������ؿ����,�Z�$����n���r���7Azy?��Ƀp�\m����s����w�����_pU{B��!�m
���x�d��E���"m��Q�$�Ă��,�����}�F�;W��K��F�u
�#��Q*�l�d���M�!vd���1�#K=ʲC'Ďo*�$�Eo�������;�
�5�<�mY�i+H���vz:w�G�<���ʸV�c��Lm�/S��C��pL����ݍ��R�q�06JAھU|�Q��w��:3��]e-N���e{����>�}�[~���l^��f�����M(&�������	e2:�j80�io4��B�gٙ�)kM��`���i���l�6�4��
]���4]�1nA��.�Z�n�L����s�k+�f2ܱ�.Ms�հ˭�����ʙ��i����K�3�`��X�̴�,p]�A��s�n���Z��T�-sjek�a�R�SU\��-A�ر��#�L`�U�4`p]̈́�-F���~��~5�t����}�J*��;q?�
���N��;��+<�7D��4&P
�b"H l�*6�9wA(��vM��I����Nw\׉�&��
���F���u���$�>Z�!�wO���7s<TT��^�9�U����-����-
�ﱙ�!:r�%��!���	&�<�$��kz�=��N�w�	 IJӠ=%�ݚ�~��"ѽ����
Û��'ۙ�F*TWg5�Pd��
$�#Lh8˕.c.V�Lٳ����֍(f��	������앋V�I�M�: xgcB��
��:�P�+�Ѡ�^ȠO�\�(�su��T�@���dܰE{źNqhW"�,����;������I6��p�l-]6J��_'�[w���Uid����=���z�
3r����!@Ȳ�e��� �P�A5ν$����w.茫S��0�̀H6sr=[��@��G�NL�D�n�u}��хw��F�S�s��(��vOv]w�ye�*s&�!)��@��h�T���� �Ű����0ăە4H'7:���e
�g�;i3_{\��]+5u�Kģ�Kuה�2]�r�b�׺�w*6 ����/P�5?�����~��s�1��˹�A��	��#
""&A�wB�$>pT��v(�M�u
$�ʠ|['nF�f�'�~'�k���4JJ�x����N��\�N��争{�c�w]{y�qP�+P|`�A�8>gbΣ��v�u�p���x[���j�e�r��v��<	 �c��$��ʣ���h����F�=����l	��C�ɠA�9�����tlJ��S�4J�]AC��DI��s��>|�KP���+�0V�� �������V,�b{�C�Q��R���A ����s��f&ܦ�����uL�a��w�M-
�;�6 ���c��ɣ�*M<r1$M����TH"��A��� ����j���ts������	�n�
� ��6	���ut���#��7�>O1�V
���@������+�4���,��I��T$�{�*��G��������j����Ux%���M�LVvyL�d'��wP�3���=��F��3�*���R^"S�2�%�7�����߲f��8u�g9�+�Q�~_�ٺ#��5�+�B����-`��LS��ǉ�	{�k�	8�&� ���^Ί�1Set��z,��6.(L͢���3`�\cs5JeZFa6�Pl�D���m��Ɉ���P�����+�|A�_uQ�,��A{��
k��)�d�!!B�@�vy�L���	�n֒	9��A󪈈�wž���}4ΐ������ ���Ho���XZ��\dMn�>�$��ȯ�ޗ�w5j�) � ��Ǌ�߶op���a�I ��z�vg+��Y����n�W����S%33n+��^8�NCX{w���WG�ov��F�uz�zj2����{+�r�"Y�de��ۛp�!YG��YZ������R�O2Q����Q%̽��Őfr�6�1��X�{WȺA �#���v�٘���λ��4����pbR�|k���u|M�>���pw}��N�nwB���Tj�L���k��J�Łt(���lf�pVj�wsue��{ֲYj���\'�n:(,ۺy���nN�.oe�����J�Y!9��!WD9�*�s���ۍ�����n���F�콍�g{(�ۭ�ӭ�y7�S�=ln��st�-�l7���kR�e�nEe��;���pH*�/�M�܏	}T����og�*��
㋎�ֻ�Q�r��ˡCz��ubHk���XT�X�2&�+1�^g3Ԉ���ԇ��̺9���X LT*�Q�4�D3S�5v����%,����ݺ�~�i�0�ͱ��A��i����:V̷5��<p�U�*#m��c��]k��2�d
�����S
�9�J`����>�r��G]�ƻ�kfnc�qqD����hĠ֔�+mٳ�.��<�X�%]����-�k�>�a`T�[���kJ�)���ӧ$'WDet�v/�w����};���D��lVЖv��fۙݹb6ƭ���^�9�u�BlD��3�����8��,*5T�*�ن�9�jy?F����ϵ	Y⦺��s�N�[����pD�YO��b�Tjuçs2jܼw��)�PQCx󓁔l���K��ޒ*�X�Kn�M"�	���Im� �a�-���^G�q`H׆T�	 �"'#m��"�KXpX���<�%�Պ9`�rF@(��p��/<��5�L %`D�bFU(*"�&�b"<�9`bXP���1�(W��`�t"�m��P�!6�<�N��d�p��<RD�P��C��L�^"D�S��b� T&;�ԯKB*,��pդR/�%Q �V
�H<p�Yj��yRb�ïJ@�yr�9S��!�d�HH
Ϊ�	J
�a !c0 1#�QB@T"r�P�y�F$ �F'EH��X��C�  @B�JD��< �!я0̽�	!
0�cb@$at�����=���%���Yn���ì��saĤ������caee�-�X�UcV�)1���(I���hMrPC#�b���y�Y�l�F����Bh֦n�\m�7(H�j6j�Y`9̵-x1�-c���ฆ�b7M����Z5�W;�`��@�v�M\�XD�ڴu�й�b�V˩1̭t���0U:ѱ��n�I����s��ƶ��ЈZ���(�m�
α������P��n10H��D1�ݴ�e�n"M�������6��-�	v2&���j��d����3f����@lS,A[��;a��;k�3�mM�E����mt#����`W6S]͋�$��(Tf����M��,GW�K��&��:�:#�1v&fs��K5�X�p��-��f�\]S�� h�:�R�i�md���:3 T¶�.��Pו�a�nG2܈١aXɡ�t ��楋n�c7;,Ѕb�)����8��8�mv�5^-�����YE�]�Qs�2Q��
��e��s/j��f�ਅX�8F�v��dƹ��j��z�i])��B�ꤵ�S1��Tvr޶�m&Ձs2�c��*K,�F���]f��܁�`�582�������gK�3J�@��3F]�Un@R�L�
mPv��Ḗ.�6i!L�<��(�BZ�6B:��R��Q��F
�WX��;,&�1����L�nf�/X8�@Knufv��nVg�])J�Z5�	��WpK�CX���K���f�n�+/Z��r�0&��t�R�Ƞ��4�:Q�j���ىA�]�cL�K�%a�m�
育�0g[-8k4�t�mk6��]��\��ih��1�n������.�+A�Q�EQDH�Y�@�f��iܘ^)y�]�cV,5�65��\�\�;Q2&���u�2�Y�s\�b��H\��ִ6#֗��.��h�\�q[Wm�̈́M1e8.��U�i.��m�ձ�sV�mF�0�U�/���z��	�n�\Xġ��nZh�bX�b�b���t�B�Z��I�!������j�=��#Pmh4��Lܲ�.�:�ŭ�4��gM��Y�F�D�%�x��#\�q�ҕIu���cj�X��,U��S���.�>v����No�0У�s��Hy�Q�*�����L
��x\`l��� �F:�y��L�9���-Q��$|]�"�=��(�f.⻜�]J=�M-
��}���:n#�(!O�a�\܊ �{/�����Q6��+R=���ݴF
�C��O��n�Z���T7���C�u@�Lg5j�)RV���GLC�{�'D4ρ*��A'��P$�����iy��ٱC��,DlлFՁht)%ge�3W�fք�Q��(���6�b�������GiU}kw<&���G����vEx�$[��N���s�B��#T��$i�o�(u�{^�H�2�ڙ�����WƳ�w;��%�r.�w�5�{�03��E�3o:\�k�ʆ��\���#Hܵ�mk��|H�yT!��#4Ä����=|}���+�}R|he��@�Ig�T�E�H�u[�Ms��Nn�@�w��}��H̐`̥2��=LoD��"�����z���1��.��
���N�w*�IJ��ٔ'�z捳� I��Ψ����W^uW��l)��2�P��#ff""&$@�6GL1Xb�:Z���c�"�B��7.�u���<L�mR P��Ӡ8gc�(
�y�CD��9z�c���P��*umP�M�������2T�)�n��7/�I$o&���U���K3����ڟ�F�)t$�#��Gę3�`P%����i�^��C'��nf��u��+1 ���W�8gd���/w�Δ���J<6��ew����Ig����a'Bb{���"hT�߁$���EםT	�Sc�LDD�n�G<[v�� �2AݕDN[��α���ۃ�X�@܊��OD�HY��M��P${]שj��=R��I������@|;=^*��P�EWZ(f��W]*�0�m�y�[6�R�լGG�����\�,������l��@C��0T����>� k90(
ټ��}�DB͢I�{k*��	`Glآ	��P=�t+���^'�y=9<HR	l�1(�I)��o�B�z:� �����0޽�J 
��l]��ݑ\l}vM���R3c��$�>��$޺�A;�vEz��g���FڣR�$$d�1��1���k.�S�^G�?Q1�"C�2q57nq=��l
�s�&4q9m�T��h���_�G:A$<�uy��\�t�fP�|{�Ϩ�vM e������*T��JQ)D�BUt���6��iI��ݳR(1?����j�Үϕ�덀H{r��I��4���������*^��� ͍���������B\Жu�����o/�
wmЯ��E6�n�O{O�zB�ɓ9//-�ȯ����O^��4����"�^Pɫ�	=�t(}��E*��(�D�I)<��Χt�dx㎝�ۗLy痌1� x�^� (oMPb �PTl�F�E{V�͏d���vE�\c!}3�TA'ڱ�
�gU\��R�s���U���|k6X]�!;���CP�ʇ�d�:�9��8�s����꼽7���'^rÃ��nVγם�M8i����b�)+��v�l��í��Q�G�Q���ԍeR�-�aҩ��G��g��J��L��Y���\i[Y`��f�����h0���.�e����y���FzǪB���<�Ɋ��8�a�Z�R�L,�K�������M�M�
JC[vs*�U��q��0E�\��\�qw)�`�Lݴb�l�ej�-��c]�r���V%@�8[e8f}���P��7R3\BZ�� [D|����<���w��Q$e�T�H'�:����V'q�]ͷ@xw��м|��D�T�y�$}�����2#��Q0l��X�>=O��H����/��]�4&���
d�IJԟ/�����N� ^��k��
{��u�l}��ҴAV c��H{	8����24 ���:�����dY� �ՃD�t�h
�
*�4I����� &z7<-��
�0Vp�g"�$u>�κ��T�#BX��b��4���@�ɝ(�J��%i.HD�b&�(���(���P�GF�|��p�E�l� �ι�hj�}9K�"�]k��66 A�""$�vG:mQ[Süy
5�ޓ�Iot.v$��F�,���3�U����W�w^�]��Z��|��p:vVy��ZqY �ܗx��zǛۯa���H'v��I����@���ygn>{;I�/H(�fR�Yӄ��הIỐ�9ב����
�$�v:b��g�QJ� �T�=p@�{aїN]�������{7�C�ݗr �,[ 
�~l
O����V�*�{���;?�o^gѰ��B��O���^�I�ۑ@�ml!���˽�mъr�C�L�����#���Ü.��@�9ɥ�-rV8P~��Gq
fQfgm��@$��GWs�f.:&#$M��<uDgeQ
!P��R�) ���\�O��a�ͣWf����|I#9�P${�$Q����E��l�B�P�A�5�Q� }�B���Ά��ڲ�k#��,X[{�Sn��v�ޫq�d��o%I(..&�v����Z�<� X;��X]W���lMf���q>=�s�;ۓD�8pq(�fR�����'��,iw�T	>7݉�r�9pБ*�������C����'��BT��S��>�z�����8\�+*I����wy�x�x��Z�-��r ��IZ�W@� �1�b�e��\�����qpKF�+rX�b"��|��S+EX�k���s��(���OhY���������;w +�QH/�I?t܆_N�#�ee��`P ��y��"�:����;��;4�jQ�Q�$@��u�Do3��$�V�5�}8r��M�v�$m����uQ*,%�
��(� ؕ�]�7vZH"��
���t�\˼�]���ݷ��&�Q��߇7� �k;/��gJ�-�L;�˫4Ca�G������o1����Nz�~0�&� �|4�}!���C�������w�|j-Ϩ^gUOgex<ݘl[��뤐^�NJ��B쪻
΍�QIuM���rJ�D��̚�eL���y~�:��L��!fe
 �wqȠ	��ʯX8w�;�ȏ�L >��l���6.�Z�� ǹ�u�<EZ��'����� y�@'���s��;�"�h Wp�j��$���x� �g�S�7a�����n��R��ʟ�v�\�7f���j�aIQ\ı�� ��A�n��A�wٴ5a�F�L���S��*8$:��D�n�l�زH#m�
 ��Nj�{v�Q'��вK�ɢǮ��п ?Gbr���-E�v��m��w�*�v�z��8%�ouwBM�
���,v��f8M�s��P>���9�m�%��(�cYq��k��@]06]���v%�g3!GW[[�nu"�g�%`�[��]oZ5(�TS8ԍf���d���ta�5�T�/$�c5��,6w�\u�5��]��薑e2� �p�n�Ͷ����[B���*�n��iBTJ�d��#3\hh\d��a�v�Ŵ�	�����9tN!�V;=�46\]�B��A������,`�f����7��dI(̥?
��%��V ��N���n�{��rF���������ް��J����f'�lq����kޮ��T�$������ɠI}R*e�x	�ި�	 ��Ok*���ez�$�=j�j� �n�'����Q®�/����s�iX�Z)&r�{�d�	�/;$W��έDV󻉉(�۲T�!��0\�
H#<F�9o3f�]B{sz�W������ǒ(��C����:�|��߹���i�.fvu�a4M�c69��U��m� ���&
��EpIA8��>w��
�́��鶱��[���y�{�+�y��&my'�pŎd�����j���%FN�R��܊b:C`�!40vmӼ�c�z��:P����/%��Sk:��/6�X��f�t��2�#Q�����$�vH�OfuP!�y7Q��'X;�*��m ����vj�C��E���2�9��f�t ٞt	Oj%ABDI*A4
��k{7�1��.v�P$���Iz��@��1Fy���dO8�xe9y���u���ίc$�X��V�ϯ���@�>v/X��O�/avQ/	�� L��	xƖ��p�cK��ԃ��,1lf+(���Y�b��d�8���@7��@�I�;�\X"gg�h�WMI{��ī���*A����ᒐ�zd�w�� {ś@��|�X+-�*�Q�>�N�ȉJ3)N�=��3�]�$߇�r��Y�ε����K� B��\����&�����l]�Cv%�P�]�ge^jau��z��0m�m�g�6�H��9V(����w�K1���[w;�)k�7�틬�q��e8���n8�@bb�j� �������j���������bwf�w�eBY������5��]�.��I�ԪLÌ���6�ڌ8!Ðr�+4�ne$dbMy��P͔�4Ȕ�TU�������=���G�F��e;O�;��:r��o�-'�ڶ枺��x��z.��ܧ�|�C�l����Z4w+'��:�����䁠{R��H��w��Hf�QpZx�-�S�+�m7�̌.1ݍ�᳚�\���k)e\�Ӑ�X��=�b���
�U�J�W�qm�����|e}�;2�a�87X��8��Q���Ԕ�c�O/9)����ҙ��9*�ErЖ1��p ;5r��W*լ�v�������u�ha��\0��D!BF3��_.�I���m�Ε���k���9s�g���j>=�_m>�J���ͨ���:e�DQ��*
d� ��Q�\��y	��=��_ �yu�c���[�fG������ӝM�ܙ8�݂op�+8�4�ڹQ齫s2f�Z¦d��1M���5oh󽵷�z����Z �p�U�����H����b��XUb۔�X
��%�$�'cW������Π@�H�ҶEA@c~KF! ƴ �
��X�g��BV0�*q��`��S�sT	�+N
rN�G�m	H�a̕�E�bE�#�:̰V'����B
@P�a��<�g�֬uH�-"@�H��P-�U�U����*�Q�BID���"��� �1�Ba�Q��
��Ҕ��U@�9c刜��j��d�5芄�U�"HE��P@8XE��	x��d�D�H�6�9���BQc�NEB	��$"E �F-z�XH�"A�j(���H�дT�)��,i.EU �F��zJS�"�H�P�*��q�BL9���d܁�X	קR�㭌!�+V'�+b@䊧0:'B�8��4y���ƴ��V���*Ɩ�1�"���{��z�f��(�����/`ȉ3"TI���󯳰d�/*�!����;w�߉�>/;&5fV�ST=&'�Z*�D*"��$nvP��nm�ml�{63��$C{}�P n{,��
4�{����bˋ�-Z:ъX�4{M�"0��n]8��i��FJ���Do1"|b&j���UA��Y ���@Pn��C���Fs�I"((&����m��3�;�8��I�|���A���$c�:�ٗ�W��/ь�:]��;�>�;��ڴ��*�.*�%�rRWt����Owk���^vH�6N%ȉ�
�%M
��pe����U"����I@��O��<�ڮD���aiw�56��w��ޏ^|�OF^$��H�V	ҡe�Ή�R�>cN��+�=<K=%M!�*�:��!ky!��W�«H�Wh)���n��ݎCN�N	��zn����������������</�>~sLf m�m�:]6��MA���Decu4R��l�������歱��$A�^_�F�t+�s�
���_V��ksv��I5��H��F�!'�"f�n��3�y�������Y'���74>��ձ�b����79��$6K[zas4���֚W|E�7X��t�n�|Iz܁��/��Y).DD�n�;ۙ��-�	Yr���H��"�Ff�;��71K���'I�)!@��S�w�l w�eIY�f�>�� =ݍ� Cs��<9�����ڕؾW�ԌkX��7�`c4�%fN�x띐[�&���U��*�@�.$@6�tf��Q���s��jvC��C:�i[)+Y���Q)x�M�pZġu[5�hp�B�Y����T.�c���ج��n�Z2�ƭ�ڎ��kaK@��N�4�����)є4{v�ݥ�cUMmz�7P�5�V�l�@k�L���Xv�:��.-H9�+�jRZB\]rbYAcq1l+ګ�l-�;5��n��*�+W \A��޽[J����+m	�����(m�7��7n�!cZ�q~>#z��S&"LW�t^UK�^$�C��vi�Jw����@�gMx�����4��
�T��0w�%@1J���K�b9�|O���������[�'/��F�}@RH�]ժ_���E�P����TT!�e�l�'Ď�ڢI��~�
	�BRA��Օ���on��;s@�Ay��X$�윝�Z�R�7 �5�@�(��C��"H4�T�ʀ
;q.+1G�K�����  �����o�h�LlU�.iw\ň�8�i79��iL����X�4л4b`�JE!��I<�� �RT��T	��uՂA ��'���VуΝ[���u��p��
�#j�з*�u�t�G�����քd���)D�Xp�s��V^ܨ��x�t���͛�w�7�U�L�k���<:3��=�u��EoO��j�^�nv����>:6ޙ��	���4ڔd�@�"��.�>��D���Е��Ż�Unz^�M�k�`�o�E	H�wV�|.ғ��
��]�|��8��ɢI�Ψ��@��	��ܻ����bBRA��4E�t׎݃�3���R�ʾ��|^vM|OfuP1������U(ġ(ǑH&�VUΰ����oL����JgXcYc��m��ۮ�C����R���}��O��fu����(��t�+sؘ@X��QV�H�NV�^rw*\��'�rh{3�1��������>�6�����v�DNp>���QY|�h� �8]ZY��q[W�x�i)lP�媓0���-�n��t���)�fmh����I>=��+Ď��4��3)"`H�ڴ�7�秊�\�>"]]
 ��u
����;Ղ�����W4Jn��v��(��(پ�7�ۗ][�����>9��>|�]H{B��>����ߣ�.MJ�Gb�X	�6�cWe��K6"fˑ�̼&7y��Ծ�I��M�ey�>�C����^���l1o�{����t�5�z���B��C��H�F����j�0	� �^w;�A��0�{vdo�3��]L�Ă��������� � y��Y�����A�զ�H:�����f�D��*�;W��N±��+� ��h�I3�w`��q{������U�Ue:�b��To�"3E�C���G�"5L�d��-펬e˻���-*Żˉ	���*��s���|�`*Dt�U��3�(
��n&��_I��$��ذs�;�Jqp4��w(!#ȵ�Թ�l��[�\�@H�q2k�:�1!�������qP%���(P#��vA��~Xo����6��vʂ��,
��
b���1A=��B�Q��<L�A��Ő��$�=j:Vu�B7�w��(�&�Q$��]�����>7���w��/��'�y߬H���	�O�"h��{�#��� �������sD��Όd��;�O�

y�'��UZF��D�(��Tω����'=9����%d�݂Isڟ�|����q�v�x�{���]�k��-!]]�iW��F��^r�j�a�n'jM8yV��߳u��q,�H�Lm�Qj��B3*��H��#A&"���Z�/M�M�F��K�5�����Fd�l3e�P�[.��1+R\�0�3s6J<[����5��f)K+�h@��n�3,ZY��`)� չn.4t$��VͶ��.�fh��a���\�$E%����Pn҆�,{]{@�%�
m5�Ɂ�&��i���5���cQ�n��@�U%3�ֵ�������5���e�ʌ�j�$a]k�aF��������
�~k�� }���|A��������Nz���r&:DiP%񈙬�˪$�;��}�v�=��$��u@����4֎�)�VDz,<��$��;��>7��$����=�v����nk�D��t���\�DDD�i��=���H�$\v�>]7B� ��uD^�a��cA ��0��p�1%K��@�s�]ގ�-mۖ} 彚�$���>$��wC��}!u	�$�A�*3cX��ŰKlsm�;'X�� E�׵fʙ��Ϸ��V�J��9��~`
������eX,R�9=Tt�׉$c�U�b��&D"	$�>��g��0<̑/s(�l�[����Rqj��w63\12;3[�J1S-��b!���Le�UO"v����;U�2-�p�uIo\���vX�A�٦;�ʮ�`���J3�v���VЮ��8Dߞt��S�Ψ�K��Y�&�&A� �!�kQ���1�;ٳ@��{�vO�9��A�e�{��I�`+�$�qI+��(IC�]��C��+F�1�#��Q �y�˰I �s���y;�d_� �*�����%�B$�&� �1uEfڍ.�,`�f�翶�+D�%�*xU�UNv�U�I'3���)8į��v�H7������S��VQ2
=1�;�v����\
o�.�H���kĕ�]��U�	C:��D�4S�ʲ|C�u�$��e�fD6���DW
T	�8ธ��*M����u�j�sJ��2cňVh�m�����<��-z��j^-��t�O����u�3��=u���(όD�`�˩��/�OzG��bω$�� �ns�C�{+p��7��و��g 4�B��Z���3ڝW�axV�̙��B� �74	�'��W�U��e�ɱ�+JB(H�LJ>"eT�`˦����
���ڳgm�`]p�p��>m��Ȫe���ݻ �7TI ��Ψ�Y��H��I���P���2�����]�Tw�n��q���X�.7�C3ڝ|I>��U�:`�ٷ�'fa���yo=�
j��a2��N����lJ$ ���S�W�QO� ���I4�eݥ걾`*�(�*T� ��]����$�O�)J��˲l$�q��G��t0�آ�s)�Vz��P�ͤ�P��y$sN�77��z��Vp��J������J��kք�ţ��3��$�\�:�O�Gc��D/��FJ>��!?I��آ�4K���"i$���TM��[�-�y���NgXBvJ�%ECM���i�X�#���Kv6j9eK�1XEr>�|��o-�h�;ƞy�d� fv9]��z\�^x�t0-���I� 	��*�H{B�i]�*Bx�z( ���H+{Pt�D��I�]�-�$)��F�݂ID�X&(B���F�h���w�$�jq��um�}�����0 {�}	oYUv��a��S�7��:�RIO=��I+�\]��H�:8�A�D�$���V1�2!�R�Q6_d�BI&��������9x�
t���zHH f忙 ��|I�����~���@+����D�Q1Uh�!@������ ���K� ��b��0a�p�f�K7G�`8&�������s�8��;$�'kZ�XŞ��+W�	�ڸ ���F�	!$$$��ҋT B�( �"� H��( ��"� H��( ��	2R� TP@	.  @TH���"�H�fnʶ�j��תC+��i�J�P�J��)j���}��*dTaR�C�M�ge{}5�潵{�;/��?O�d2�¿�d!F�.C�c�} �VZ8��w}'TS'K���,�#G��z,^h=��Xxv�M���]B�� DT�?��=����>�?����+J�C� T�E�C� ��?�$$P�
F���?�1����@{���?�W������ac����S�� l>����@%_�����O�����>������h��8���#�(;>�q2A:l~n��T�"�'�g����T^8�4dɅ��f� g�~�>o� ��c��m?$4��O���~� �Ǉ��O��YD�1����D�@D'	�P$AqEP�>�� u@��ddb%lh,��zi�R�*�'��n�G|��=���'��� ��!JT#  �$R��*�H�H��?���������>�x=?��b�B�.���)��y�{)��)���}�	k���r���J����̬WG���q��A�z��b|�_�>Ο���} ��f��ï���<�,?^ ��h�~G�m�����h~#��"��>���<S�xY�@�Cg�o���}B ���Þ�>vY��~�!�����<�Ada� ���I�4�FO�0AQQ���"������D��'���L�'��0?_�q�y�����4�����j�
��H{˄�� ��j}+�΃�TTTh�J\�����8t.�������,�T�O��>��H5�#���}�Ÿ4J�hg:`I�� p�("��~3�>���?��:��A�����?�@���q��������d�����{}�S�����O���� �����(	��,�q�
�=��'���C�|U��%���Z?�}���?ȡEG�~O�&��|AD��h2�?���G��*4�א4}��?�`?��}���������l��?��f��0 lB�??�Ő�-['�{~�>�x�����x��ǧ�S�rX~O���k�y���#���I����B ���(|����jbC�Y�>'��?#a��p��l(��>`�=�}#��H>�� [I���G��0!����dI����>
 ������a� �?��������{;���
 ��W�>�����]��������3�h)��
C]_�b~E�M��$�?Z
T�$	���s���v��.�p�!ۈ;x