BZh91AY&SY� �B�6_�@qc���"� ����bF��           ��E @ �@ $ (  �QAT�P  � h@   4P�T   h  {j(IED*�l���Q 4�
5��*%�Z
)�@�Keh
2�`��E-����
�4��J+��6���p��kF�4tPm�� 3��P��6@
�V�h��*�iB�5���Ti� S@P(j�� tMQJ�  璔�  a�=����l3ESTCL�U2���4��j��m�ARSZ���mUIa��Q�qY�i@k��� ����Q���+_=)I  ����횠�\����(���x({V3���{T�@���][UM����K�>�Wn���ݽ���z�ǥz�@=�� =��T��ot��vP� =
({`�4R�(���� `v�
�i�W^<h�곝�{�oa�Mk]�o��3v[����mm���{�慠��wh�޽J��@��������黻Lny=�ON����@��E�P%�[`��mL	|��( 7\�w��)���y��A��s�������{Ν��F��Z���4)O]-���D l�y<w�A�hG^���̞��ڞ�J�I����֍2�gjQmM�(R�m�5Z6�ϩJ�=���=h.�-v�ݯ=uٺ������͢Pwv8���]��ݱS�m��B�ŷm5�4�������s�G=�=Q�fv����M�ң���N����6j��j���6¶f��ҥ@�|��բ���ukJւ;���2w�u��P�����=kӠ�8���[f��S��\4:sv٦曶�iq��v�ZɝO\�e��C��aZj���})I  �ﯡEV�t�l
��Φ�S�ZuqҪ�a���=b��^���s�ӂ��9[���(�ѹ�QT1��tSw@��l�[Q���@��T� ��\��qs�H��n�N�)j]��)=�,��]�s��-����Z6v�@�.����x���;��6�AS[!ElcCA_>�J w�R��V�^��@*yѝհ5]����֋k��^]���ۇ������$��L�����Э�;v��&�u�\4(i@ ��f�GϥJ@w|�S�Q�=��
4��8k�P]ս�j*vIwi�5[^���Q�;��E��u�nn�հ#M��m5x���  � � �*T�      T�1%J�` !�`�~�A*��      5< RR��@!���`&#�J~�))�U       �j3JI�!�x��L�yM���=O�����G��$|�W������K�0�o&���_/F�ߜ�{�3ٕ��Ҩ ���ES� *��������@_���y���G?�� *��J�I'֐^�0"���@���~_���LO�Ŷ%��$`[ؖ��%�-�lb[#�6���m�lKb[����%�m�lK`��6Ķ��b��%�-�lb[٦�i�lb[�6��%�m���b��6��-�m�m���l`�ؖŶ�4��-0�`�ؖĶ�-�����-�lKb[ؖ���0m�l`�ؖ��%�m�clKb[ؖ��%�m�l#���%�m�lb[�6��:b[�6Ķ�-�L-�l1-�lKb[�6��`[�6Ķ�-�lK`���1-�lK`�ض��-�-�clK`��6Ķ�-�lKaLb[LK`��6��-��%�-�����lb[��b[LK`� ��m�l`i���%�-�lb[�6Ķ[0m�lb[ؖ��%�m��lb[�Ŷ�m�l#���%�m�lKb[�6Ķ�6���m�l1�%�-�l`[���%�-��[�Ķ�-�lK`[ؖ��4�AlM0-�lK`[������cؖ��%�-�lK`[�Lb[Lb[ؖ��%�-�laĶ%�-�lb[ؖ���-�l�m�lb[ؖ���-�lK`[db[ؖ��Ķ�-�l`�`�lm�����6�V�(�b�lTm��� �-��0�(6�Fب�[b�[[blm�1��E���ب�[`�lPm�-�� �m�-�Q�`+lDm���E�"���%�Q�:b�lTm��Q� ��Fب�b)lV0�(�� � ��V؈�b��ؤb�lDm����(6� ���Fب�0� ��F�"�`lTm����� �F؈�`�lQm��lTm����(�Ķ �Q�[`�lm�-�Q�*6�Fب�b�����
6���[`lAm���V1R�(�[`#lm���Q�������lm���
�U� ��-�!lT�-���U� �� �"6�F�*�[`�lA�*�[b+� �� ��@-��lE#-���@-��lb [[b�lm�1��� ��F؂���[`lm�SKb+lQt�R؄blm����
��i��li�-��"�U��U���شĶ-�m�l[b[ �i�l`��6Ķ-�m�L-�lM0m�l[b[�6��cl`���m�[0-�lb[ؖ���-�l`�m`�ؖĶ�m�lK`�ؖ餶%1-�lKb[ؖĶ%�-��lb[����m�lKb[0�0-�lb[��Il0m�hm�l`�ؖĶ%�-�lK`XĶ%�-�lKb[�6Ķe�-�lb��6Ķ-�-�L��t���-�lKb[�6��F-�-�l`�ؖĶ�1-�lKb[�Ŷ�m�al[b[�6���m�le1-�l1-�lK`��6Ķi�lJaĶ�-�lK`[L�0m�lM?��">���/ݝ��8���S�&��O+R��1	k0�ͽ�Zo+^�Ar�0�bn�w�Q���%:k&]R�J4/0-�H�o(hT����2��(R2�KJ�����u�zsd�t��n)�ՐP�̖�D�i��GJ����c�$�S����kn�[ڔņ�ovf��R��aVRN��P4���/��,w�N�!�*�����ѭiۢ���,���j��K���Li�1��UbfM�"�g�U�Y����i�̪V(L��kK	�L^-��F@�U��+.�ƭ[�D�-�O��L�&�6V�y�۷�=�׾ܺZ'��@%r�Q���jGiЪ8���u嬦�U�3��VlUVKX�X;���KA���-��<���S:%�з(���3.���n��:��Z�7v�J���5�7b��\�MM�rdr�6��7�E))@��лWe3[��j8�K˗(fm����Y1F�V�pf�)��1`���4¬O!���EW�q
թ��ѻ�BN�/	�j`*[M����Ef���^[��B��W�tX%�d���׶AM�n-�h�Yt�XW�DFFd�I�*��D�5-Ju����Of�] �c�e�n�Ok4ռ4H��o*�Ғ�y��Yi��f��6����ƞ	��x-��TN5jȤJ
�G5l�Y/uTŘ���<�f�W��!з3/4TX��[�kF�f��;��صP�u�m+e�U-�'C��V�-L��	����V嫅j͹��l��ͪ�^�1�K�nUSl��x����E�^�a)y�+m8�����W���@��2R��J�C�f�ff7�mL�͋qÆ��^ѩL�ӥm��f�ZG�詶���(��cں�V�����ip\����6����vػ�c&�i�Ǧ"*��1,�ku��JRA��*e�)ݍ�6E�b�ԓ,1r��-^v�ںlݍDAF��r�mZ�J�ڸ�7�n���j���ȝl��^%�d���ӊ��%�rγ.�timhM�Y��uyaj:NE���Õ6��VkVwn;�7�H�Z6�^�F$�$c�b�إN���KGU+���Yj�Pht/U�;4b�Q�P�:�ZT%ާ���F~���3.k����t�.�a��
�P�JFX�&m�]]���r���t�f��&��p�'��f�z妎5j�v�i�4Z���5k��7���Od����F������Ƅ�U�0����V�ۼˋsU�Y��ͪ3-`T}�ӭr6�%ȝ�*L7y�j�9�Y�N�4EXJ�oh;�D`#�j��X�N"^�����ʣb��,�+0�OAM$����6a�`�(Z[��5�����d�P�1l�sud�iM��d�YUXn�[J�p9��w�%m�*^��{p�*��,&�fv�fH0�Nm��gT��!��$L�b�"*�ʭTeV�7vؕ��Йk/h@jU��T��[7f��uMBb��yFҵDml����PZ�a��+M[�B;)�Z�DV�r���J�����,Y���;j:�7PL*�إY���7b�˔��]e4YX��CS��\�ߘ�t���ʻ�����C]�e;�������P��X��˴N7	�s3)�RU��-<� ��ݳd��{���'2�e<BZWFԱ����Gh�9�5��{`���L�uv��i:ckeʙs�Q����獪�fcCi��P�[{��	���
�0dG1�Q�Y�^�B
���
����tڡq��K6]��e��U�Ę���Y�M��K˺�Ñ`6�:��S-[V�����Y��dVlF�"+Jm�^�.��W��"jŜA2C�q*+�uX�[��\D��Y��6�+2荿n�ZzN�l7��R�{-N��L�g/5"�A�hR�NZٹ��ǥ�kR5=(ڂ1��Y镻��x�+��ɔ�]<��@���M#�"f�n�@ڱ�b�+�7��@un"V���¢�-���r��[�W�0��C�[X�P���e^8�!Q��+-��/x�a�9y���n�e��
Wj�a��36�=N�J��!�Kqj�u#�Ӯ��Zf��[�X�AW��3p��Ѷ17K+
L��7(�5#&��*�lL-
��ҋ�D}oTw�oF�f�.�kFݍo�Z������6�2�fQ�鴱�shV4�c ���t]9��)̻��k18�ڵ�	�6��ĩ�5���L;���\�L;n���SNI��9Xݩp�J�����*:Lۭ��&f:n�1[�{h��ȋ��I\Ai>4Vj�Kx#��Q
\�a6�8�l�Y�F;nЇ�&�!xM���D
wvR�3�u�fj�XB �W���݃�^UM�eh[�Z��d�V�K8��W4����yڹ�Yt�Ą�fd�O*�p�&��+0g	�VNʫ����M����c�%��uIS'!�.�i�1d"�����j!���Tj�"�e����R�\�6^�m�ղ��ҙ��!���Ib0aV��첲�xF
���YSZ�xJ�*)��V]�$!��Tӛ0={`���7��D&�"b��~h��"A�NV�U7kD�V�J-�f{u�n&Vd8��8LͬԶK��f�AU]�e\��,��:��Mt۵%��Bk�1]�yY&���f�fՠ����步,l��=3`K.��t��R��j�����"�wc�3Τ�qej�f�㷸/EG*'i�Nb�2B��v�V��B� ��$�/n�)��T6����½���^)�̵ͭ��kt�r�n9T7v�ud@�!�6<�3�_<o�<��lYhI���Ŧ��X�E��˛{RU�6]�h�VrLJ�U��{4ex�rȒ
�K�V�d�xX�1:�n�U�REvm��<gp�~�K.�!"*jw�e�ӆ�d��t�h�Lӧ�`�!DT��x0��&�Wi\;��(-�����M]7���`�̅EY7�b���*��BG�Ƀ^��Uz�F�P��A��iV[���M�*�$�^4�!�!)�c�����!x!�W��]�����[M�A�G0L��n���y�\'F�
˽��yh�R�0�*��7�Ĳ�Ң�֫N�ڔ�2�I!*��/e�֤Dƅ�e4fl��(Z�D���̂�Y�n���M��IުzH�n���T�X�V�n�2;W����A��fV4��ԝ,���T^%�ٱ����Yq��^5V,U	sid�x�tV�7f�vY�=�x��3��s*&1'q�����a۟�L��Q(d�N$Ö1�,�0�.�bD*1n�L�nγ=TT�ThV�p.��n�-\7�5eXq-�NZWa]!Q
Csrī�ZNIM�@P>�Q�&!�.�n�UUh×M�L(����e�l�qQ�ym7��:�)�U��c6^*F��7k��Rd��i��hE��5�����*@��"A�1Pِf+حL�2����j�!r�\�e����E�����fƄ��M�%�����Q�aWU{�u{qnk�u�������J)z�n�X�%��-V1������!	�����`��7y*��Sܣ�#{E�f˂E���ҞS��*�ך����ʖ+<�w�7d��O>uL��7(����V
�U���(�r;W9��j\��m!B�2��Ng3MD�%ti�l�9Fm��+�!.ȕ���oj5[)����u��77q\��Fj��2I���
1Cj�8�Vd8ʇN�$������D����M]#S�9����4��i�r�u��֤���l��d�fZ�ٗ�H95��4��/dF+�r���{F[u�LJ��4�	�U�c5�e�先j�ꝑTaɨ��U)%Dv^Lv��ʕ�.�h�3�&g��'"��]kV3Hbr¸�����T..0��Xr����ܪ�X�t�u�Y��e�@���YkfA걵��X%��̥JG�c9�CV��-��q�����H���t��eS�e�R���%`E��N�y�&I�D!��vh�9�%,���suՈ���w&i�vE0��#�~Z��Ӻ�EC[�i�q�wtj�ޣr�w�n;{F�M��k`[�r�Vum�pj�D#8U�@�k:B����,v#�d;YZ�^��ڇ
a"�{�]�7Q3L�+V����zkp��V�5,oY̨}t�ݎ�̱�uW6-2�aЪZ/QI�)%�cV���2ۊ�*���L�2�Y�ȳ��<���Po2�$�:B6B�U���Z͝0�Yz��P�V�tt�����V3[^ch]��F��n���^�#�B�Ct4e����{ݺK�VNlk����n�u��U�EǸ�ul�-�́�M�;�,���̙�oAg%b��DЗ�M�M`����h�I)�q�����hïPu�^�Z]4�h����{Ԩs�^�E�
ecCfY�E�0�=������=x�֣U��3��P�կڎ�]�5��N\���Ԟ笻's.��Yp`���E3�Oj��Tv��N���Ʃ��:���S9���N]T�l�F�
ܪ4�t���VT܃�G7���'.���+J������	���f��<��J5*nf
��m�^�Ǘ��Q�:���5]Z�ZUv]`�uD;z�ᚊM��$�crM�3�,��kVfd$��3)c��80�b^kV�4����'wIC�nEq�r����v�
ZDPm� �;$JDe+ �{Ib�H(Yq�flݻ�vqC� �Q�C12v1%-j�U�E?���f���[!]e��T��t�<���ѽZ�j���aM��5M#:͂�ɣC:p^՞UW*/C��Uy~������Y3,�U{.j�v�5ҶD����ȥVJ�x� ���ZV<�&�ݵs<jXͪ��:0�CV(oH��70��Gm�K*�YM���*c��X+h�n��:4u1�r���S(��ՌĶ�a�M願�v��,��U����J�l$E�����Qh��p�vn��	D��6�U��m��Q��Off�u�5f<čfI��)Շ����Ī�I�pY�Xb�Vn�2U�mfh���q����ݴV0���[[�SY�����
RkL\�5h��w*n���5��[�bn�h�)�ʉ9T*���F2�"��F)UF�Ѩ��aYѸj�)�2�6�Ō!�yf�Ub;xn���$��m��Lf��r2gI�2���KIƌl�TiTU�zꖊ�R񨴭gnj�M:��c1��77/sh�Ѻ�!�i�軇*�f�MZ��r�H6�})ʧ*lڗ4f�dT�n�Y����K`�W�6�Z�d�t�D�m�9Vae^T�D(��1�4peY��y%��-왷5T�GE<yR��Xr���,r�Pwr�,�,�����-�G�Eb�GvD�t��k52Ҽ�F�ڧ$X��鵳^&e'*�XQ����Z�JљT2Kݑ�u��,��ʔ�EQ�{�J9��u{㭷vK^{���R�S�t�	khU73 �ۼʑ��̈Fe�TnD�e��*������y�fƮ��^Xc�BVbu�RmU�H(�����9(l˷k
S��,;5Z�!�5UNz�w&��@�p"�(\F�U�8�G$&U$�݆l�9�AdA�[��/UXy�/����oJ9YTn��(JєƱ�`����QLi�Ei��I�e�v�7�ܗ��mh�#��t�G*ɭ/&Ӵ�А�Qx9�n�,�b10p���x�Ӵ�Q�j���~Q�r��d��wpX�T2n,���#+�������
�YqܩPcp��5��m�Ҥ��I[�Q�p۹	)���o*�0K1%UI�y	+
:ڧ&Ai��: y�K\�&-�B̥n�j��4��w�+S�0�'������`Y������R���jM�{Y��W�(�,�NS�akO$1V����&��K˜0X�)D�*�����52�@�eMŠ�E��\&�����Ȟ������31d��%mI��n��nSv^`�X���j+ae�-M0��˸m�tCj&��(��f���0�̹�8_��63#�n�RN�`݈M5�6��Ŧ�I�����%T�a��^Xs)f�Q��{Z��2h�K����T����]Jj�]�[GT���N��W˒�J�MZ�N�j�%ں*�)l�r�+V�ԻRwef��✶ҥ���$������-^(�$nh�)�jf��t�$����Չm���V�糉��qt��WGF�b��.���k�5-J]�qlE%���W���l��\��+��])��`�H��r�R�J�Z�lQ)x�F�]4��eu��I'i5t�'jEqU�����b�R����oP'j��ޡ�DSj�@s�[���*��A��<�W^�4��;I�������p����+T��Υb�PJҪUK%��4��R�E1\Ui5@֣jZ�o��=Wb劃^��9�u,5<Q�I%к��ZݶD�,I���S��w-�A�G3)k���.R��ikY�j�]��+\���<R)žAS]�����X��7}T���4Zi4q^%�ibM)�:g^	ԱP�f�K��NJ	/M�,� ��%��WD��Z�R���O������WGhһY��q JF�f�Z����u��n�R���֭���GWuz�omk���rb	�K�QU���B&ҥ"6��쫧i%���!�&ꑥ��mL��Ω�;r��I���.���dq���W+�;V�+�I�r�V�qKRI%t�*�QH�-�t�meU'���3Uj�z���Q���uΥ��/+�\'Y�=3�I;E���\�)���U�5�v����ud�W�)V�qu.�R�FPC�^�Ij�Я}_.�ܚ�I5�-W��[I'j$�If-J�@�[��N^b�flӵm*�4m=[j��N%��8��
Եi�ѕy�ىj�Yk�`�W�=1�k���\���_#�J\�M$�-H꘺.�z�Q#ڣ�Ź�Tl�o1�+��0{�$�$�%�֥Q��qRY�"`�g#k�M$���t]Kq�Nꕘe�QP3��ͥ�mD�I���\���q�]{X�ǽ]�B�2�[	�]��P�%d+�1b�3�)1���RWI�[Z{-j���\��,]�e(���KJ�ZMZLﶮ*���S�;RD��Uk�X�}L�kqlJ��~�����ߒog��~g�B��K0o�.�W����~9��sC�	�!5.�4��I��n�1��W�Wz�mb���_�J�q������3���
m��Rb5T77V�U'j��m�ӌnR��R9o��z��l�2���οpW��l*��c=6�ʥ��2���]sk��J]r����++�7���4�f��x���i����;�����Lj�c-D3}�e�:�;����'u�kmS��l]Խ��.Ыg���P�3��cɩ۪�6zK��R�;{�8��#���j��V[9�^�qh��a�⵽���-\�SF�Ӈ�a�R!	��Z�r����%t���/�u�ק��l=B���r�`��{vk�h�QGk
����up�M	ٺú�FY'N0/5[���-1y,b�Cu�V�n���"�b�-�};�T�z�#�Mk&G���[�Mm�wץ;��*����Xɼ�VZ�0����P��\�ьZP�d�P�A�����Q�yMJ��$�Th�͛]t���ӥf�WV!���J�b�qԚ�mb�Nŋ���+�,��Z��ө`�	�Ȩ�bZ)�]�{Y�i�ВD�9#w��cQ���qzL`�=�(�u�9�m����u�o�'w(5}��b�C{��j=�v�R�8k��:뵩0�O(�̣������݊r�
��ך���4^���w��T�K���&�or�������ceM*,fv^S���� ����]��p�����Æ�RQY(%x�X��먯����B���$#��-ʪ6�d�2���U�P����P$�66��.Ꙇ��+[�Ag��ӘZ96���P�&v����\V��xM��;37�iNb2���c���Q������'�yIC��T�ee�
���5��7Sm,�ڙX�N��
[�z��������'(G�Cƍ������s�2��ĺ�9�t��V�Ѹ��tɍ�V��`����v�v�R��{Q��ߨ7G7
��N�@�UNKi�1��.Z���\T�nU�q�*�iq���!e�pq]�\R�]Q�'�U���oK���a�`2�ת�Kub,h��V[F#2\�wP�fS7�U�m�ތcx�gs�ބr� j��hA��2�sY$1�+�P�����6��u��c宒H��wU|A�V���w�%���qt&�ڨ��EJ��қ������{�n�Rڻa�GV1o4F�qn���d��,l��)����18��M���}��N�����|e�;z�6�ư����'�a.h��h�������p�a��͹h��&�ɸnh�k��v,�a�YxS����)��r/N��|E�Rt�U��"ʂ-���(�
'�۴�M���W`ׇ�tgeӘy�9t�aE%���f��<�E7mUe�gxVgdˬ�.uY�3z��¬(���0ɚ^_h7jr�G�K^CzލJJ.N��v�¼��YmE���X�6�T�RA2�ȕh<���ȣމX�;%�`�I!��,գ/YL�-�r��-fP0Cs3�8��t%���k��Z��YHs�3�&�;�M��2��"k`�)Nj&���'t��r��s\|�p�^���5M0X�&2��yêO6Sd2�Zɘ�p�����率i���)V����Ru�qu�{���w*V�y\̝[�e��w���i��ռ�&�aX��t��5��H��zj��ǵ1�U��]۩���h2Uz��&�:L�S+_G�[%�����n��9�w�y�ŹՃ	�p�oέ�̵ΆԺ"�:m�+�9�3���GU�9�ɐPA�
˻�����#pa��l��P"�{��r�MR���!�HmU�V��o��^�v���N�p�+c�
�A�#:�Nk_[�zf���Q�12^e�$��J��-=݉#)i�CR�N5=�r�j�#d'��ܛ��{����7�!���c�%]���wzf�M���[�Ό�;et��Kqr3��s���y>��)��b|)�%'p�5GقՕ���"s"r�ma��X��B:󃦕ٗ�ku��CM�ư�P���7����v�-�����Z��"i�,�ۻ�ڱ�� r�����]�t3D34]n������,�.޺T� �Xݎ�Ǯ��%g<5�r�e����+N��&E3��Z������2`�����Đv�����$�޴]�f�&"�ĵ��ʕx�q��Uv��)��n����O�eٮ��e��	e]n��E[�;����i�k7�Qa�]9��dD��X�t�=k�Թz���h��U�uVWa�ڹL����[nË�T��e�S{�d�J�kG+rq��ٙ��ŇUoEnv�b�����f�[-�N�Pi�%i��Zq���R�R�r�2~�'!i�3���	��u+ҩ�f�tqR*2��fh"+#C���i��|)k���n�^y���d�F�Ъ�1{��x&�Й�{�kfް�+ ����;8�W�J��}�8�0ܺ��q�#Y��a�ܕڥ׭ᒟ7�w�E���苩�rֻu'Fխ՛x��H�����:-+�%�7NDFB��W�o"�=�����;.��:��Ӻc��45�T�Bh�7���l,��\��5��yWt}v�:�֌�R�/$��z�%���}����pfOE2Y|���ɀ�o9�� �S
�n��;]+*tR3�k�:��W�cٔ�vB�S��r��EVᮑ�L,5Au��껠�NL��uL�BcUcg�;�a+w`�uL�VmU4/��^�d�Y�3���Y3�:-�nɗ��m�fvh}(q�:�Ի�ܫK*Y�,�ژ�㱝%v�i�u^X{F�h�B����Or0⬇:���Hᒘ���/3&���^mvT�&���=��א�o�V�Y�5A�3�<�s�52c�c��e\2��۬�qU�����̪[Ķ2oQ���u�O6��w
-�

�k2�Zxc��wZ7e���9$*��A�5*�Z�n���&��n����]3�3v�L��!B�sJmN�%̍n�yL�J�|�Y���NH8��{]�u����6��c��K�R˶*�5�w�6��:v��]���Pm&lvFMVf�ܲ�S
��0�J�f�к��y����ظ�	�/Q�,��"�m���w��T��ʵ���{Ntx���Z���a"��R`�^����$����Vm��'��fXŚqL����Y�flQʛ��WuU���+��Q!f1�ّ���.�xa���6��f���[��y�R5X�C2�]�2�j�TV�p7���cJ�TP7�j�uë���/���6��]Ʒ��9U��T��.&�_��%U��w=u��KO2��[Kb�g{)��*2�92�ve%d���ɪS8�T��aTb����b5�2@N��@��ɒv��������ĩC��&d���u��[V2�U�"�bscH$�gj����R�	�\k�&��Sa�8��w%�d-5����<p��S��p�b"C�d����8�Y�l6��](��Hy�s�R	�����Y&�tI�+be�W0��,�9[�A$EAʵn[���h⺻�J��Vu��i���L�f�b�ɡ�%�
�uL��]*G�n�c��<�l��	qo�[�&7y/{e'gޏz��q]�]�mE��j���M�D�'cm�dݎͫ~칧aX�(tsM�l�(��r�Q����������v�:ͺY��qt��ќ��2�*�}���
��)��}��be9Yr�ZX���P:o"��3z⛱���6kb�aq��F��5y��A���ID��"�빩�ĺ'���V�/�CW�dߩ���J�'%k"�{���$���dV���;meE�Oi�N"�L��՛�)�Ŧ��`���6�]Z��*�K�2�tr�U��U��f5w�nVޮ��{��w"�͏�maM���iI(�X�f�J���*T[�0�}�$�w]�Zl��B�r�|5R�-�W/[	 ���FJ'ecT+�l4P��j�7:��ۆ�9�/d�%�S�����rۜz����т�ó��/-�gsN���1Mȥ�3N��Y6)���q�ڛ�͈$���"�YdY��v��8jW�teS��V�c�w��Ԏ��5��Ȣ�ͻ��9���J�"5e����j��yʗ���i���m�U͍b%�ք�W.ޗ|����V�C��ٍ֭U��wͻ����7]K�x��nCv.�eEł�ۇ`�ˮYRb�c�:���k�m�-�4��N���T �l;6��ˋ(���L�QW}��O�ﷺwn�lán>=�z�vqQ��ɮ,��AC�Ej�7\��+��sF���Dڏu6I5�-ĳ2�Y/��!�o���&0Һ3.qӉ-�����<qf��]��{sc�:ס���n4��%�^:R�6�G��yk+mV�������/mV���Ù��nCv��3ۀ,�Kuܳ+v��Z�ڻ2�ԑ)E(P��hLZ��coQ���cl��.�3:�*���q��Ж
���dH蹙gj��,[���b����FQ�(R�%�WY�۴���`d��v�ӷ	�I�q��	�bN��+*7���a{�U�4��wJ��,��|�nsf�����,˙h�!d'�
�y��1>#2�1<�0�i���X�����
�̘�p�R)���UV:�QlVy�_�a������j=����ố�h��n��E�$�k.�K����Uݶ�)��S�����[5�cU��pWY˕[���lc�nnQF�ʘ�<w�9��Ƴo�MX�&	{xęW�՚�n#qf�e�,��"�M%�;�%t/3:اv�>��&�fk��vMjJ�+H���RZe'�E�v�%����N�.��9��cþ��I�iha�-7�f�}�ǒ�(�[v��:TF�5wvrnf]o������k/u�W[&_8��f�x��+h>��;e����;��jז{jW2J�]oe�Y�\-�s���x*n^Jٱ�᭼(d	�UN޼���%k�r��������\�z��ض�51GO��
-4肴ꮔ�e�"oZx5����b�#.�i�Z�-�Μܕ������CN�U-�H����!�w)9��n���4���\v��YxӍ�,kL�)e�*�)���M�yLa5�6窮a�����^��;�Ǽ��q�vWq�A΃�{U�^Mڵa}q���T�.&���K*�g%\n"������[4�*�1a�/A��%z�T�V�;�I1�ŨEט���ie�w�v�`1Љ��W�7��7��n�PRջ�{(ms�d����n�����˼HTmty��Pl�͘&��ٚ�[��H���o2oq�;��c�u�ʒ���D�p��udT�+�Rӣ�jE������[�A����q���[h��R���n���6Q�!TȬS�灲�xF%q�_P"��+5-T����
���������vm9��^��iڻrb��+%���}T��N�V�!�z#��v�x'�)���42+���v7.V],G/8�W��	+z�͡����z�nǻ�oo%:7��AoMraŴ-�V�����2��X�Udf�f��f%���A9d�ƯKXE�Y�Un�ΗX5:N�YAמd��2�n��Ǎ��(6��e��n�g]J��(�Zj^�+S�]�>S��]�|sg0/�7�u�M��fYVnUB�cr�Cs��UX���ru3SlmgC�{t��XN��|�S�(Z�K��\ԩ����Ⱥ�7NX�c5r��[3����[{n;�H�q��I}zs2�7p�A֚U���v[{�W{.�۳U�3���`���2�ݹ�Y�9����v���Nᚫ��/uË��R1Ncg3wn6�xw/>���1N�q�ڕ��Uu����*UlRn���W��Po�3��F	�i�e���:�6DUdۦ-�f�f]h�Nb�}ERq_N��j5f�H[%�	Z�k���B�R��
�כ��,QL���y��c&0�u��k$UnN��	�T��:�Č�Z{�5blX�gk�lm8����A]Aˬ��z1㜯��]l��%ٖ�������x��t^��J"oSNdR���|	e�ƃ#���G�#I8@�jŰ��Y(�	��܂:'�<��<�n� �!�B�[ם�r�4�n:���-(�Xw�����z�F;���W��b����<,�}t2���c�7��ߕ�|�2����4jxyW. {5M��] k�9���GuW�UJT����o4)3�������@ 1>|=�f�=���F����{������d� g�i�4�S$`��x|@�I#�#�3�� �r�F��&*`(d�G.�}��K� �_��2�ʮDjH��rjP��7�;����`כ�H'�P���&����PG����6�"�������S�?a��(#������>߫�$�������}ߖs�y,��y�w{�]J�5¶�bͳc��F"ت�s�1�]hԒB�
����J�vt��f��cy�/�k*���X7lyEܧ\�ThD�n�ZQiZ��I#z�Fmi�u)�nن5b�p�G̮ͩ�x޵N�h�]�B����K]Vi�]i7��2�iu5R�-Θ��`��,F�Q'R�t�U}v�FRd%�iQ�������N͌1�[6KBe�ޒ�HK�\R8�5Q�a]�s-�˨ݫd��L�Z���b���33�n|V��׹A�&ּ���e[��&䩛��8���L����vS=���+�9cYW��BMH����M�^R�]�X�9Q_lմ�U�h��l�PT:L����ےv����%ɮQ�i掾=-V��.�F��2�\�|춟#hJ�Cc�$�6�:�;A.�e��Y}ݘ�.�&'�7yC��J;Mʘ��0t�[�&�uG�*n�ۡ�r����eL1̝�{��)��n�m`�dα����T1�����F�x��4I���
/q���/,������C30�,�
���T�׸�x�O��/N�ᣢZ���wʏV�\uޥ�uRi�{��u����vu��%)��7��snof!KyiN��s������@��ؚ�ޮ�j�����8��q�q�n4�8�>�㎜q�m�q��q�N8�8��4�8�;q�8�8�<q�q�q۷������q�m�q��x�q�q���N8�8��8ێ8�q�}q�q�q���8�8��qƜq�q�n>9�sw�+��Y�lВ�+&�L-D�Ep�,�#P�7�i$[W��Lk���;�.c$f����Xl����i�}�����6��O�L���� ^ ����Cf��rY��%l�õ���{6�4���j;M��Y2��ᚎI/�w����]��/z��|��'�79��׾��8L�� �Vu�t������e֞J<��=�83e,��,���+k��.��.�Be����-��[��,�Il��B7DJ�Βi���_l��PL�0�5���t�T�"��w�)�HFm�ΤmWRܗ��F
֚<E�f+�c��3wr��4ߒL���)�mòq�ê���=Eu�غ����"��ֵ�Lڡ�2�um��O��kݴ������sv�UAyj�v�ۥ'J��OC���)�-�S(*ͤ��M;�믰�.�VT�)<�M�nNACv��L$u�f:ʎ=��S	�&������:�7hQi<H�p�g!f:-횢kwAO���GˤB��CR.��UNe����M�Va��q-ps���Zׇm\�wfZ�l!BXʵ����.W(�k�p����CJ3�\Ž4�$�kW�k�s�78۷�ǎ8�ێ1�q�qノ8�8�c�8�8�i�\q�O�8㍸�8ێ8㏎8㎜q�q��q��q�nݻ}}t��8��1�q�qノ8�8�88�8�qێ4�<q��q��q�q��q�q�|q�m�q��qǽޯw���i6M��}�f�|��+1�<�P��gv�_ejl�S�����K��*����S<BO��8����	�8uSz�i�:ʲ��:��M�i�p��ݤ
���==�J��+�\]N���
��D���\���#��Ooq���{l��]&�!u�͔mv];��E]���R�]�ynl�-<T�2m_ƋH�y\�ݬq���N�,TP+)�̡��N��*�ۂ��\[9��Ys/�j�1�m�1>�MXw�伽���Dc;|�e����(��6�4��Uz�ob�n��F0���H���#3��gF�p#�9	4�����ν���H��r�ã�}�q�W�U�]�	1�
k�j�⢣F���M�jX/�k�Nl�n��z�����ܷ�:���,�Q�!IL�/m���37u�=վ̷���e�a8�bSR�E�Y��+{	E�͇��
Zs3P�C�&�����6�F�������{*�1�:�d�\k�ܖ�f��;Ί�t��ȧ}�*�1����Kb%��5ڭ6SZ��Q�m��/Z\���a��`��Ԙ��ŷyBȹu��$V�z��4QQ)��Zc��2��Ɖ�0n��O'&m�e�9Z��z���{u�ؗ]�����=��o����:q�q��c�8�8��q�q�pq�q�v�8�8㏮8�q��}q�8�8�;v�۷nݸ��8ێ8㍸�8��8��q�\q�8�8�q�q���N8�8��q�q�q�n8ӎ8���w����y���qU�����Dyζ��|Nv�@�g7"�g�Q��J����/��5Ct��� ������{�A[�U`vE*���Ao7f���ݪ��Ơ��6Y�;t��#��	�i<��w���9`S�۱��Gk�i�8�na����I4�ط9�f�A$F�:ε\�6M�ĶV<�I�d&�T��9'�xe����\�yA>oO2���I�Te���Qw&�z�P�6�Vj�5{xE�N�i�!����O�qH�qa������Ib���V��f,�;����:��F���䊷b���̈́�δa���S{�x��h�����c*�4�o�aǎrr������j�x��ͱ/hT�4�u�?hF6��9��x�:M:���7���Y]�n��-,�{�Ŵ7gL��
�*ɮ���D�c�PW(��Y*�=b�H34�h�W	ŧbي����F�ph$�s��%)K{/�lz7�t�D���h�P��}W#�: �J��+�\��6�p�/�Z�ڹ��,<��f�gE��/�5{d��R�H<������	k׉-�*�i�2��L��݉ ��u�[�#z?x!
�ʷKe�\S�볘�i�몂@�˵�74�C��*�
�Z����D�R����<���z��8�8��8�n8�6�8��8ӎ8�8���8�8���q�qǎ1�q�qǎ1�q�q��;v�۷qێ4�8�>�㎜q�q��q�q�N8�8��q�q�x��8�8�8�8�8��8�8��84�7�������f�6�8��2�ǧ^�nU�#6�el8�y�;޼}�BL�Chc2m@o�����q�f��ggnvٴ����>�)���U-�������(�3JU�7/�P=��Q�GzꃿX��P^�Wi��ү�m�[u�t�T�Lc-tw�t"K(�]Y��3Ui��9v	q�Kyލ�N�eK�T�U��c�R��ً�����Yq����y�6��n$2f�n�W^Vn�ڳ�&��"�B��U}Ok�Q�32�Y�y�������\i�.�2�`B#o%���r�miC��d-�r��I5��7dᭁ9�� �cA[�=]��X�n;<��W�k�/U8�&��p�c:�0�dld��� A�kg�wo%�m��t�		�^�\)�J*��Т�*և\׺_,��b�3D���ٖ��ʨ�Ui�� /P=[��Rj�B���+
@���{kB��&�f!�v�����%�!^��mkmGib���)���c�=�Ai����-�A�*�ߖlV7���N&ܼ�c(S��Z^�L�BM+�OQ�[���O� �Xl���]=$��NUj/^�WB���O��f�#熩k��p��]�����`��NB�Ɍ%ܶ �;�r.v�Uf@ 8��G/M�`� �eԫNh�����r�Z��u���%�M�|h�p�,ր q�+���<.�������B��qH��)�X��R�]0��=�l>6���8FX��x0G���*;!]iEK��������v��Ob�]��U������vQ���]�*���(:�X����Jã��w/�j��r4mMA�[b^IѤ)r�V-���^\����24��	h��n� ����>��N\ݥ ����n6��R0n�'���e'�S�b����N��5��oj�6f��/��7@���5X�P��^mc�^ܦ$��#c����FH��z��\���=�-���n,�޻;�l[7^rqOKY%VP��VHD��KYA���^�x@�������t�����O"Wj�㗹��S0ΒEUZ"Yt�k��lb�=t8��&��.�a]5v@xr�Xec-pΔ��s�(����k���ݮ�n�m��"5�L��s��c�V�o� ��|��VF ��3vֈڷy�}{�@syv�Qy,�o������<��k
��{R�&'5*�i�|�0c�{Ǯ���&�Z75��ov1Yw����U����r�v�0��=[W���%#�/��HU*�<�y��7���w���_�5 �!w2d���BտL�o�$�)���ј^`�9y��{�1��}!�{Uf�ͦ�m�1�)/i��K�֐�E����O�4�M���j':�e]|6o]��Gb7��r�o��u�p�:�.���^�=(K�yFʴҭ�d+eJ֬+Qߨ�]
+���	`��9ZC�����_J���
�DnQzK��B�UuB���I$N����t%�E�I�݌����Nf'LÔ���¬s�[�+DuT�x�,��y�Q�*�mM�`£)��WBk`���Њ�M��!�k4�QuU[[.&$f�v�L�y|r:����7N���zbx]�U�rә�gn�Se�� �������77EZ5vN˪�&�K��L��Dr������D'۷T�ޣT�Br�]ծU��TtD�pmUa"�V��}#�w��Ti�ไ�{�
��㇀ȂpeU�8��U�ma�]�����0�;G�҄C��9V���ۭ˾�;Q)j�li�j������<+-U㹚Gmc(1ά�\�R�WuV���Mo�2���Λ��8Oop�V3�J6��{��-�bo5�-l&�:{%Q�ov����*S}�+W\�C��r�MU=R��iYN^^R�6薲�<"���`�H���d��QmU�I;&�}�O�vT[]Sy]{��&
C�cc�KT�\��n��QwV{�/95si�n�؝VL#��!�PىE�z`�KSU]�'j��)bڋG\�)�]bN�7lYvo�t�B��Y�y�k�5�t]{�oK��y����A��Զ�z�����{6�3��Ώ�ǅ��R�z*�#�af�p�V]�/sm�j�V�J��`ޅ+TV���A����G�v��@��b�;��>�R�\ݪv�!V���9rIJһm�U�"ڕ+:__��W<=�+YH�&#Y;^5_F�8lde���}���k3VQ��,�E��|�LFD�m�Ŗݽ'� k��2x��ҥ��:(�89x�I�ڌ�����&�1��KƇ]=�j;;q�c�o.[��j����^ݹiһ�����s)��Kz�7 o����G���Au�m�������;8./��uKz$��U�w��I�s��!B���×B�D�e�z�"��)�����{bh`�f�*����`]u{�jX�V_NJ+X��z��&oSG*�\PQ�'�8�ݤ�^F����yE�6��+�gj�]�僵�����m�]tfz��}n�U$��U�K���[ٽ�ץ\A������0 �Y.�淚a�F�N�OcWڕV�ӬG�R���+�Ȇ�Q9ܺ��=A�NR��
�΅*���(V<�֬,�u��ɂ�)�OH��ve8��wT�'�ԣ���l�ۗ �&.�
�9��)<��]R���B�ͭ��9S��촩I�F��8IalF��)�ݵ
�'ej�v��c��wNf��pB�u44d��J�v��:���5����ٱY����&ˬ^���֩P.�!uu�2K	�F3� �X�L��ܼR��׈�a�3���r˥s�ڣ׶�������盪��q*e귪�@��J�R�Ow	������N�8��$9V����i
�b�#�s	��d;��Ϲ�fyG���;5m��3{��4��E�)]Ō����˘����sӗ��7X҃�&PqG��^��kT=��%#�Xw���*wS�(��[ke�(M��H5���I�r-4�N�v8_(m=Z�΢��Qik�����E��!��,h+7������**޽=%���t�Ñ�e�=*��tsw��gKы��^YeѲj�b����a#q�M-�(v҇�%Y~�vɒ�\��=K����d�o-G[��GP�7��L���)~޿d<%GިV	ȴ5;gNVM�W	��F�q�V��4q���Ṹ�eAgoLU ���Ĺ�h���u�yv&�ٙlQY�6v�9TR&�a���{y�p�e�Rb�YsEeuJx��u4�ǻ��{�A�b
i�gn�o
zӭ���e.�Kɓk[Jl�t*٬X���U5����c��U��F�]jV���]/n�����@i��f�j^V�y���Q��avX�4S�!��D��^���l�Nn="�HܩJ����Q��N���,�Uӏ^�+o2�ޜ�tI�m�������6i�7vmi�rܬשQ�Y5�����k�F�R��k59�+t�56gN�2�-˰�(�0Td���)���5ë�uJ�; �!�Y���e:�����J��Q1��l�ʚ�i�D.�]�u���hT��۹�_=�2V
O:S�)̭�g���Tv< ��xfd{X�
��Ěuw�jn�cNX�r�ܼ�;�ݝ+���騞�1���ֱז'J�I��X,��)9պ���l"�bə�j�Y��d�E�t�
�US}�_�sm��l�����X�١�ǎ�<���yYɦz��i);k���U�I[���b����\�*��vV�S�V�!�v�bL��ț�u�֦�N����,���.�<�A	o���v��͛O�PC
�kf-n9��
��4���U&5�ܾ�ѷ;,ܡ��y7pȲl��;��4He0�U��kQb��B�#V��A�Y�6�2�-VKv��i�;�+o�J�M�w�{Hn駚�wS�r�����( ��2��w�_��?��_����~�������H��8�nZ��һ�f�A"cF5`�D����S&~J12 ��f0؉�d^@�HH��!H�p��	# 8�"j�N2"q��0c*6A��"0�^mF�	��.A8�I�lQ��(����"MXHD���ꈨ�.D�(��" be`i����I�P�$� H�:�MTJ0s��J4��aB����i����EH�$��XL4��T��S�R7A�(���,��d��АQD��L�1��_��\6�EH�lE)8Ψ�Ŭ�ZsJ��vsܼw$�R��Y�sU������!�3wݔ��v����va�D���,�]X9yGjLؔޫr�JIk�y��2�z��
�C�yj�{]U��`-��h���cm��7a�I�P���j�o�gU���ӷ&��JЭ5E�X�A�«�C��Pa��Eףi����Ƅd���9����-�d�S�2��k��2�Т�=��\�Վ�ۋ:9[g,�ٔVӬ��<I�u+*�GB�������f�#���=p�.N��U]h�ܙE�ݖ9��rq�`����8��W�F�!*�S{%V F���02隹��q�B��V�fֺ�6�۵���l��g�ЎR��$s�]�ư�ҦRx���4�ƾ��CJ+˜T�'vr��v�Cu�Z�5����A�7iz�3���Y-��2�YEjk��K�ݪ����x��IP2A��x�T�2ٺ&v��u��m�g��s0�QP��v��f�ر&ۊ�����Q�f�d�+;
Y�mN�yn�4��EwM��Y֚]��]��(�n:��ٰ�[Sgz�.��61��>OOoG���U�N�:�;�������GJ.⍄����(�(�M$�R0S�[m��G!)�K(�T`�5P"K���p�בm�ɉ	P� ���.!����
6�iM��) VUT�Q�8YE�T	$��(�2�KŃm�a��-�O��DQ-
J'�<��iBa�-"�ȆZ�H� FQ4|d�m&��F�((�
7b5P2�@�̑!�4�&�M�q��DЂ�e�>b��A��&]RT��.I�[g̒���Ba�!�yy��TX��:���ч�"��M8a1C��-��1�

'��!���M<[J���j	�CiYd@ꑩ�i6"Q?9䗛QA~0�d��!h��i&mԎ�eP$�"�M�ġl�b!�Q�F�f�*"��I�QA$M���[2
iF����AXG�4��e�b$��%@`�p8�4�l#����, �0�P�	8P�$e��.'
r$mD��D>��oo�ϾBN*r9��(p��K�E&Z�%FB2��cO��\v�۷nݻq�<�B������4H�գ����H�q���me G;w�}��}�۷nݻv����fJ!!	!�oG	m�( ��H��s��[b�(q9��q�nݻv�۷�1��F@�a8�S����~5�g8�{j϶��m�v͹��V�!UQ��RRF޾=z�۷nݻv�ǫ�.����m��7�Z/k��۽��[mlZ�gu��{��֮���f���8�m���3�"�Z�]bۻ"ò�dw>�]��b��L��.�ٸ���wv�vq�n�N�㬛T]�Yֆ���=�9�Z���kq�u�q[kv�u��̺5�m�m����,F�Vű���w�pq�V����8G5�Zٶ;GZ��ik3��+XH�V��6�ݜm`���b���<�]=��M�ҟ�8̢�"�ִ����pW�h#����IGw�ok;���.��?M��$\�t8C2mX\��|����(r�:��#�.8����'�v8�9�W~>��޾|�N$�0�Q�(�N"��6�����$�[M�MB	�@�R�q�e�#	5����Y�Zї��{�r�"����������K`�Q3��[ې����^5Da�1���
��Q��'ŔyH�.cNR2A�H!όE��,@C�)fz@�""0�0�!�q��q��E$Y�����(��0�
�,)�m��`���i��)��%���x=W���|adՊX�<2���\*19J� ͦ)���4Ԑߚ���a��M���+*��/�����*�-�Vص]��s�,<���|8��u��恗�n~t��n��w�o]spF���M��pp$ݷoX�MI�$䤑����.N��ޡO�e��>̏����d����G��.E�j%���jj/��݃���� �]�ܺ9W@�V{�F؛ڜ�����q8r�(�xqD��������|<�[x�"�ジ���Y�~���|�>I����o9gsw��uHG��bΠaz�*f�F��N�)���hH&x��g��F�1>s}���Hv��;�[&��_�H����[s�W�JL$�ZD�����J�W�jx������;'��]-��V��y�K"m&����|��:p�}���N>�$u+��۠jg�×��J>Dmej�N8�ͻ�e=qv��x����rƬ	T��S��(K��0�̜E:�ۼ�B')l{�b;��-�̦�xԪ��P��J�O[V�LKun�5U�%��k/:�%��֓��/��ӊ�5@�N@��A�Ru��у79�5J�
�v.E�V�����Ӌ.����T1۟P�!����)�G"����[é����D������k�|ʖE�3r�j'��\�3�p=zü�/��WU�y���S�Yn�a)9���89$�lm�Pj�*����bc���10���_ck�����~|~?8�+g�j�םy�����\�8;��Ņ!�
������&;�λm�B�U|� �R�f��법t���#aF��76n��xs�OP�����+��î.KIanwa4_K^�x����?j�NW���>]P򗁬wd��J����XK.7	�O��`[�ٟI�nO(���rqr�y�@��r���f!ca�q�7eW�x������6��V�6(e1{��oS�U���&�q\�a������;�³zV��R�-U1^�����g_/�I��}��Ζ[�Vj�X�EY4�9;vl�BC�O'W[�A�:���s�2�L"s;��
�໖�m�u�]'Vpz�-����<�_c���Vv���b�ğ{Էv�mwZP"'���k�Q
�M}f�k�WM��������*Qq�o�vfs7�<�shn�Bg�ң`�]��7��o�$�ݚ��[K/�C�J�b8�M@EX����vG]V��J�w:(@�2W�>V��]����T�X���2E�@��[�gZ�w��m�g;���g4"�H^B�.�˱��?dXA��J�I�ɼ�2i�c\�����k9��j�8[6�5�،3Q��8Au�Nή���B���{�0�.a*w�q_+M�5�A��o!�������h|FѰxKC8�S�]m�]��C0�ܻ���J�+��J���1�V�t�Ђ]��S5\�ݵ_`ۊ£�-[�F/w]O�YC�F�u*��ڀ�=L�%���&8��Q���r|��N�_]�m��6n�̭���Ӻ�v�R��e�u\��Fu��&�_P�����W>:��++ucĨ�|	�8w�阕�V1�+R��L���:�}5g����G.'�E�o�Eq��K�A���,���I޼z���;i�[qJ��6�ߒ$�nj��T��W{	�)]���i���޾εv͵y5�#7EsP��B�yɍ��tW`�3��1;��n=o>��g'�d<@̛�퓳�|R��f�V�3�e��'�x��!XU�Uws3ϔS!�a��㶷�%��kW�
n��Y's�ڗ��0�;�8iruɇ���i��c�x�/��a�V�8"�1��r�\�~t#s����l��٬����Єo���svy����"���{�"�2�{�-6�0��x̪mWˉ=���0�o�@v[�U�1���w�����ױ�_H"�p�������	�/�x��u���aT*_v�\_E�6A��/�E�������.�79���s�&��Ǖ-���=h�9b�`�=�΍�f�[��.���P�����3.wU�c�r���%o�JG�wסI2'@�Bg,bv��Ʌ�J�*����CŹos*T��$�']���L��E��q��0h�5oehꥺV%w�����	fI���/ҝ�3"7]�u�7	^˛�!eٳY��S�����7S�:Ԧj�rBS�Y|��aH��R?�Lʺi�g�������&��FrԾ�Ż���3E�Q#EE��ʢ�j`Ҩ�m'��!��̃|����_nq<(o9��(�������م�����_76�J���X2�J%V"��p#�m��	�ύD�0.�+.`�qݽV��ܘ��:`IA}U�S�/GӮ�{{��K�t���c�λ46�����H�"���F�{�{S����>�F�Yma�M��a3<˩�T seO:�/�6XIOr��;]F��o3�o�;�5���}I�c��[�;��LP�#Mq����oA=�m�ٗ��t�T��� �V��Ϯ��3'��Gl�.亓9&�.��Ҕ�v��v핟.�|5����bD���r��p��3��A��������Q�,��a��[QܐI�fQо�x�G�Skqb���r�)�7�r�Je#�>���֚ǳ�nn�~��:�3�B�qfn�Z��kT��t�5�ީ�[�7v�X}U�d{�k>��v��J�&�Tܫ+���qX�M���w7c�+��P�[b��e��:��vtQ��@FYӼ�|��'�X�T�,�j�Udj����=�@$������B�:�RV+>��KJ|q�yY�!������K)<ú6o��j~��k	ԅ���S�={=��[Y���k9�V��b��c�H9Е�b��Ӓ���L觤��I#'�=Z) �D80��;Lr؞�D8	-�ʮ˿tp�5�"����}^,�^�'r��e�]�j1ܘ�o���;I���P0uU���Gp8�Hi�S���*��]��������,�Us�]܂sP��g������-}�f|G(I�S�𻯨3�a/�}��dt��Uv�����9vk�g���]l���xE�O����{�4��t�/�r���b�MÀY�]p�
��u�+�;V�+��QB�9b�UZ�����	���u�:��:����^O��U7Qެ�&�^;��v̭��P��.�UBsx�ӢK�U��c�-��&�k��y��6�Do��礯���h���=�5#���q�8Ts�z� ��`�jP�w0:@]o�h�7k6�W��ڸ��7rJ�>�wC�1�j�jϭf���$h����{i&���������KI�s��/�)��[���-��甯�����W*�̄v��Na����X��n�tRv��s�
m�䚶2
��.b���&z������P���3�g��ҝ��s��s�F���sx]����{��$\�}o>�78%Rá3���F���b�9�>���qȥճK]��m�]���G��O'b��ɂU��-���sn2%��#ݘ�o3�w��u��>����BC��ؓ�������q|��Pt�۟&�ĳ�_�b�}�5rj�
�֮ԛ�sܦ��������[X5w�p��j��a��b�;ǋ���%lfug)Mf�
�
*;~�]JȖ�L��dr�:ݳI�D'�i�;ҵ\'`��߭�7�1�}�ɪ�}u�c���'M�<Ul��q[2����{��
ms�g*�ob�M����z�<:��o��ל!�6:� k2V��vH��
>1���o����?;�������PN7�db��7z��f���ޮ6��(��LgPK���VM[��
���Eg#uW��Vx��J��������+�d:g��R�R�E/�k|�c��x�!�wh���as6��C�E|�t�UP�b��܍�]��e�No�{w3��϶��F-�ɩdh�ق^�T��uQW�B���U7Oqwɳ��<��W_����K�:J$R7�5�U
�㭗}��3�LA��v��-*����S]����}fN�aK)��z����<t5�\ޮ�6��vYB���ʳ�;�Ww6�`�Qrvh��݌�{�mO���KvI��'�(}L�'�S_a���ʵp��F���n�AZ�թ����j+�#��9]ʆ:IՑ���ycr��UD�ʩ/�����=uGmD���*�;�t����9[5ײ���T"pxy[��
ݱ܄�:�}��\����ԩt�w�E9嗉5B��გ���Ad&6�m#��J�2��ճ"��˱�RF�^*��7�x;s#)=t�ޅTQ��nٓ�f�|�RX6����Hմ���̑.D�@��a�U{�6z�sc��D�:�:�*y�]4����*���n���9Ճ����m}����>cK��Cz�0�{�����Mb���Mqϟ7�\�q�ad+,olOӗ�l�Q�ψRH w�.�Y�mf��HG+��M���2&+U�yTS�� �p�Մq8:�{z�
�D�v�5`M����N��_��4��q������3�1p��S�O#+��δ���ȼ��f���ٮMk�'�EI{6)⋠�Gl|��?��4�!J���f����S�k�� H�&I�$����dѨ��Yb9��+0]�ľ��cO}<l�u�ܣ�gPv�V�1zs&��h�tU��[��o#� �Е3��Lݻd�A����2Li�\y���S�iJڶ�G�&f�jBı�9�Q*�sα�����Z$�7�scZ�p�A�u��*�*,�o��tK������W��]�h%Jmd�3���ye���������m�>E_Դ/N�ÓF��m����#��ǷYb�=Ƨ��'*9��#�}�O�������u1`J��z�`�{�u�B��LG$R1!@�lU���/�LV��i�:B�����.f�"q��Z�K�|�[��bCʞڒ5圧z�����UGva�y6d^����'}�a[��7���c8t��.j2��G0��W�/�SW��տ<��<��9t��Fp��usV[���oj����r��o1>sc����X�[p�8k�^��!�R�]X�\Oܰb�}�S;�m�_�e_�q寀�ʝU�*�_����D=��>�οg��H����B��l�}��+���W���Pe4������*��r�mP��y�g��|�pn����<A��h�"{��{x�u1"Ӆ��rȵa`�ٔa�O��}D>�/=퐛�<����y�{�M��>uGY�E�7���Y8�_w���!�R�-�0��S9�\��dL�]�s�;J��w� �Л��*W��Sv�-���L������֫�J���/�V��׸m]��x:�Mĕ�Z[��D�¤�-�pt�7Y����υ�W��^7��c<�n-��=V��e�F�g\��a&SmPŅf��m��#k�S�]SE�]���9ZeuV��m-�CoAWr�5eڋv�9;��n�vۣk\6�)d��$zOu����)l����b�2��[������)
��N٧���	�7]Yo�3]�A�&�U���.�4;�蛱���)S2�8�p���;+��x��K̆�8uIx'R��B-<���,aJ���wT%�;�D��ŵ�D��)ט�MQ�1�h=x�o�>��6.Qo��75�Dt�<��v�4��{ug���,ʰm̈-������,B�����Ն'R�V�u.��f&�1�M$����z��5�4c;Jfc�ݩ�C,���/m̽-U��R�+:�hͤ��56�{
j[��e��C�]ר��sBra�	�Ob;[�&�ؓ3�T�g&p�U���{���9)�/Q�']��u�]�Q�U�0�Kn*�o�_u.}I �M�7k��SI+R��胦[c�綊&ﶳ��^���Xt8�3R�����$�/1�Ì�Sw�c�M���U,��y}�;u�Ր��Q'�S�ݝV+�L�YЩ$O�Y�Ͼ�Q�<z�$�zG+Ŋ�y��Z�^�����73g����Y�슢��R�V�(m�D�:�ut�U�mLB-�y;V_0�k��J�#��jeիŝ��Ӽ(L��Ù\�;lr�5s82�L�Ν�wU��b;�H�)M���Z}��bV�n*�˘9F�jBO��]6v�w�k�;r�
��NZ
����eD�΂2i��
��-��c��h����.�bZ)٠ҍe�-�[qI��K��Ƨ�piE%A)�2��1��9��n�JB��֝����o:\�f��y�g��r���[��p×���]�9�eS2��S�[��N��k�&��;�%�S��D�WRtV��t���2Y׺�<��ɤr��Xk[���4ZhA���c�J����)�j��]�	�W��;Ztcc:��&�M�J2���ޫe3xi���l��a�:5��}�o��HkQ�жNL���_;�X��E��F�f��uy��Z�͗�I�a�j��d��[��s,j05�ۦ�P��}�؟L)�t�ה��
�������n�i����v)QG#0�:QZء
n-Mi�E�qŦ�[����۩YwV�H�K�y�7�b��J{B�'1OI`�y5��=oh����M)U��7���I�$~;�gBr#�%!�wI%rDT���÷8�ۏ<x��ףސ��$)�k�Jpy��ZB�u��L�H���8����T��|q�v�۷o^<x����q�k�y�[�I-�u�;��o�i�O�ã��~�n����nݻv��׎=�$�j�$B�Tt�3tM\�Cn�g����)#$$�A����i��^�q۷nݻv����$���$$� 5!-���#�m��Z#����i���Nf�I ��I:HNA���2��Z݈$HQ�΄IV���.J�I''^��?5���wBG'_���P�q'W��XH8'%�EC�m���!�r�W�@qЄ���/$�JD�/08r�
��rq#�)�N�͝�g9�$w%�%�݉�G8Hq���H�7m�[[���^���:�A$0�[��:U[�2�8��j��3��}��;�Q�8̺�t��K�,�Ţ�^8�x��P�\k�8Dw���cĻ�y�y*��P绬� e���	t�k�!����w��z��>��-�<7=%��5��cً�.�t᰽�0aL���	���/~�x�������^͐	F�z4�$c�}�ފ��&�q\�'�:�>���i�@3�Z�1��?�a�떜�����y��F.p��a���ҍ`[��py'O�5������7�f��E����G�2�X wD(�} ";�\�� &���}������p���=�f�$���d
�C���=���ۄ�Kջ0��,-������Y���T���o(�%wRt 5�͌��h��|�V�(|V��_�O�xR~���9�t�)����ך׺댹�~eN&9i�Y��yo�����p%Dc"��]7�q,d����ё�a����z%�1j�/��*����
q̄R�	�a>���0X/g�č�T������"�)���a�u럩XL"6�ܜ⻠�;�S��:�e���O	���'7�xBy��P�;�(zb���S��4�H�P�>�#;�� {z�+SM����]���^�t��Ð��`r=*za߫�ʼ*�"����q��	�<=�e���L�o5��Z�`8�9*����P���4�y��c�!G��q%bЩ8���s����}�^��" �Ft*��#j��M9xr���`S³ݬK�ut��ɲ�^�Ųj��-ÿ�^bY���|�{�MU����ߌ��D��B��ܩ� <8��p>܄]6;�.:�e���/ܑ�~@w͇��A�7�����Sp�� \^f-��=�;v5���+ �s�~��nþ��\�|-DY!��G�p'����-�K�Jb�R+�24�^�'�8`ދb��9��:�a�=?�^w�O���>YHz���D0nH��m������
4|&'�.��7��7Jq��K�D0h��F���r�P/a�"m�:�L��^B��=��δF7�탞<�"cm�įO�gU�/�ׅ{�$�+�Z����!�01���Z�qN�ft� <3@�.�ao$|d_���oq����T@��<�tj	��I�8bI�.�Ŭ��%g�V��a��`�(2��[Z���p�	`���w��]y�/Czg� SF�uG�c���Ֆ��8�e����Hj �>>����l���9���a�y��z`�9��T�YQ���9|64�����Y6ѽ�-�c� C-b��-u�=�	�*׆ǃ2ϛD��z��W��ʈ�����LB*���ˈ�q@#�����T�G9K5���0U^�E/.UZNU��J�5cz���[��q�4inX�ц�,�3X�-�v�9w�qI��E��u;(�[�[|�����-�Da������,��X�u^�A�RQw�K�*&��1^j�N�sը�k��&����%��ܩ�p�}�+��Q��)��Lh�!���;�:����]�g]t<:^�YWu��FY9S��Xw�������z����O�%�\�o��*c#"w=����a%!:��U���,ѕqqnS���28���:�
`���F@��	�9�	�2��O0�[�5��)�Xμ�ĪfQ��{����ɽ��n������g��k�8a�f;�\T"Mσ�9n���?����h�����R��5'�m����<rco�ѱLY���b� 'k�ʼ�:�~J�������&�w	�2����b�s�OHC������_0����45Y�E�p�ӷ���^�b'�p�l~���_o͡^��Z��^S�N�y�i��N.��-�B�O2�S�4'�Zy��[��b���rСV�Y%{�CZ�� p��L`ّJ����W�Ϻ��
��d^�"�������Jgծ׳���}�� bS����ǉ_��1��ߌh�֧O���{�k=�� {�*�듒w������s���{͓>�!�j�_�Ot��x3�S�� �O6�׶���z��F�p��x�ܯ{�-�܇`;��-�aS��Ǣa�/�|��@�*Y��9X�Equ'���T�f���ԑC1R�u�L'G9qڝS��Wmޭ�]s��TG��fZ���{�J!d�(ʙ�����fp�ٸ�Vf��I��k@�1K�$��Ƕ����me�_�]ꪡ��w�'��o9��뢟Lj�hd��$�MQ������fgf�_�NI�{׳VsvazF<i���p@��/��� \G!_����uZ�i(��r�Ӯ�52����+�5�:
z�rF<[�Or黟��:��C�,=P�'�,��_��2�$����~��P����_��\�%�@��q�ю?h����]�$�f�7��&��Z�U���>9�����H�$P�`����Q���H/��� &˾4�ܑ-����S�.�����{��[Cג��I����IZ&Gt}����٫���GT�6�=^�� 8����қ�5B3���6sjgO���v�-�:/��	=������ͅ�R���C���� �}>-�ޙ8��xY'�QLhi7�k�.�������$\�~�1�,���l���v�t�%{��څǱ�M���E7�&�]t��7@ƽ��uܰ��>���X�I�<����c��/��O"uzc�V8/�;�M񞇢bӁ�a(,WB��3����p`�=��:�+���=փ�`������p!:�$a�������8����UD.��Lu7�/�n��Z�]�Xvd�WMj�����>e��*�+0�졵z3G\��j�ÜUًF�P�{f��N��;T���RW�G�tT��a�r�>�|^A�q{�l*�r�r�2�Se`I������k��uodyK��[w,��~4SM%4�4T`��t��>k��i=�.���4�ҹ�9TQ��1-�#�>���R׾WZ�
��ܮ֪���%�|c{�ѝ��.��탕�L���!�.��逹�[�e��+�lK�M�<��H�CMq��|�zq�q�ij|'��#�X'F{���/�^������N�a�Q����R쭜3�}�s ��l
���k��~<���m׻�ϴ:<@��6`�
��#o�X5��1���.���N�({��k�NR����^X��r�2$���x��=�5G�XȊoCtصg����J��/�����]��Ht�И��:a
�~es_BkP���,$#r��C�.�%Ls;�)�7kQ~�W����E<6�3��	i�`5���y̿����0����b� �����TSy<�m��]���ڳr|پzǶu>F�-�k��ay��L�E��4.|���"1�uE�;5���/V]F�qT<H`�N�`b�dIp;�6F�.�%��b��#�Ht�K��K�WTGr��n#���/\zش�6\O񁃦%�I�'�K"�ׅ%��緞�^��A��y�?C���mg�vbJ9�uq���$�SM�+bIͭcu���7+��P��8&�g5P������ofU�P'��ӻ��ߕm�qd*��X´T�Ӧ,�"V.��;�^�P�="�kkl��g�S�o��o�<ּ�I�_�!M4M4es�k����������YI��E��@ {���.X}�s7���Pq�.�}%�Q�,x�I����í�\*M*Ӿf���W����E��u��p���a:�g@�^�>�T��(�9���"�x�����l��
7�5�Y�]���?��\85&P$���i/���G����p��!���������9�P�8ŧ�wm2���������yx�xQ���0}��;������c�W"bc�@"��kϽ���`���+����|E�,���J�����ns����s��W�흂���`�}�52']]�mf��14D65,��gtP-��2�0zo�S�U qyUAUO�kӸ�����,:N9O3�;�%�9�}�ۤg�*�<o�(#�!;Z@?@z@�����|�Ӄ唇�׃Gf���+:�kV3�̿J�p����6��t�<3)@����Á�ţò��i��lY�Z8Gg5�.�����l$?{���߆��}h�07�� 6>�N��o1.k緌���u�ï" q7*���ֈ�L�0<�P����U�x2����ߕ8E�ޞ���;\��v�\%�z�1d�o-.��r�W[�|���C!?)sp����o��ū	�O��}�o~�E}O�k��o�H]�i��W�x_��x@�3���f]���Nga�"��}_�f�o
�ʻ�:뎯�ק3���6JT!�X����٬�'n^�r}A$B?M)QcM�M
�MEA�0�]�}�K+}��޳2��T8Mir�.0�x.�b>0����T�����:�Јog�g�0�O�S[����m�����v�_�(!�P���k�z�z.H�nq��{w����le���@nGMId�CW�3��y4˜S;y9�=����'��N����r���j��(03n ���
|n��aX�*}͌�aN2o��n/�k��m/}r��<C�����=���F�5|��V��|P'�	�[�FDh`��AcAb�X浊��#�"˵��|��θ�x��؊���{��] &x���:�ؗ��d�n8"*s#"9����} R�@�U-w_2[9�n�����/�W�N0��I8��]Ӈ�pE����(��_@��T�7��>k�LC^�q��M�1���2U�a�!��7!��z'�sȷ��n��|�xm�U�������fT�89@�<akLx�u8/C��Ӹno<C���ψ��#ށJZ�n��:bI0i�'�P�O����RؓV@�����j4��)��k{����V�A��fb�^�ݾ��G�����c�e/:�
<;;'��<3��-���̩�u�P= (.rg�77�f�����[�+��?BRtu𚫥tN<��
��L�"��ŉޗ�!fN=�Zk��%a�)�NE���	��;�z`�U�J���M���s���]|1qz���zXw{���FjgT�Q��%�αn���y���H1�i* ��
i�Zi�* �����H����۟6-���ނ�L��9`����G������s-{*	{`.Ts����1�a֪PtA���-�V��g�0p�xc��'Lg���7�Mn}�]{P�{f��!�ZI��ي�+�0����f�ƞ^2���3�#!��p����~���z�7�n�.�� �2��m�~٢��k�_��9��L ���R`�/���k�|ϋг���?N��br:݌��r���_��f*�3${��A���wT��1*���� �C�M�d�^����	}���l�E�ǡ9�{k�ƁW�=/B�zJ�p�J�sj<vaL/v!�Y�������w��q�����B!���n���j�R)���o���C����j|v]U����|���y���E3��@�[����C�����ܟ>o	-l/OzBd�p&��7w7�-�b@x����;����z��xi��z��1�mܙϔ�@����is5f܅�z�� <t��C�$�*�Њ�o�v�5��Oo>�ËdȾC��Vul9���ן�l=����Wtu�*��1q�9[�q��Į����f�l;v�!젴j2b4�t�~��O�X��c-On��ͫ�S���UQB�9�#T��6��˸��E��q2��� ��8Y��ۙD־�����h ��()�R�iR��� ���Ȋ�$�����,���=���R�89�	b�Mz���F�מp�Q	�\@.,t�B܉�~�vj�қA2�����s/K�l� ྔ�;�E��Qu�n�c��wx�ܵp��qn�o2x��Z����CFG��B1�	�ͷ��
��*u񞇠E���ƗJ��맳��*f�M�DI��0ƞp��@�2������"Dk;:ub`�5{^�@��`���0�F�����1�N������='\@˯B������G֟�i�C�ط�9���T�- �\:F�&������<�S�>���j�N�ﶅ{2��*r?*"A�a�$�^a�]3���oL��v>���yk��1�6��S����q���j	ʁ@��+�9�/�����i�n�������(���D�Ő����G/3�P���^~��a��4�u�O��o&�e^�Py�|��L04�f�ؗ�J����2*�Cf�7�b���T4��-��l�����"V�������p��%� ��$KO�\&v,����\���|/,Кޝa!�D��ӷ�|���=����]%ԗ�Fف�h��	��u�!1ֆ'U��뎮�h޻�vm�a�z��}�oX)�1k�����د+���r�1:�9wT2�*)���R��Td�_j��ܚٺ�w^/o�����Y���9	���i�ȀF�D��iT��D���(ȃ ȊH�)"$���o{��;�����;]�R�8YU��|?0ջ���=����йu
�7���bt�f�5фx�ey�0c����:��8f���w�Xqma�{��L�E�'e�?o<O�M.���a�vi����Ku��x>����d�#�-�	��'��U�P"X_�5	U�1��b�
�����I�iq�d{��z!�ĲOa%(���+ъ݆cЋ��y�7�q�"T�#ӺM���ba�P�+ p�P���&%�$�J��Q�~vk�!R�z�4��g�h�����^�����ڣzD���Xba��3z�$��1���Y~I�Lq���b����q�J`�,�?��{ʖ?'��|>~?����p��;��P��e͊�=A9�=�Y΅�ļ׶2l�i��#h��	�ଊ��$~�����g�������ū#m���<�xP��x�JBn�'���6;���L�>o[�L�>/B[�I��?v�^����*ܩ���w]<՞ޔ�P�������U#5��^;pC�iT�{7_'r�=����r�9�W��L�]x�����7�����Yt�Ms�Y2]���u�na�v�vߕ
S��iS�Tw[�Ǝ��������r�C"i�Ɲ��7:i��Z�T�]�:yM��2Cm:�K*��"]�W�c�B*{4��,����C{�WS�WJ�%Yo��qf84̫��o�^U��8��	�1e�J�T�'��K.��:fք$F�'�F4�,UǻC�m�Nk����kOU��Xt�q�5m���k�!�\ʽ�N���6�wVIL+}��	1�훗�c2XדY�"A�{�^��a&e#���`��7%�jq�/;�Z���a��ӄ�^����{��Kkqh[3������;(�V���41Ҕ�_a��_5����(��t5�"��ۯ3-��7��6։�K�y7���T��ٻu����*���K�2�q�}���òn���m��,ܨ�6������*LH�̧���u5V;�T���{4��8M�9iEn�Ҧ#\2�������a@�s��z�u�\r�����J����H]q��n.T+��a��]m�
z��;y�Y��KUi������$�泩S�	������+}8$F�v��w-ʹ����f��۬�UlL���g,��V@�	@FK����y��V��k�2�l?+��u���!����5�Щ�P+g��mPȽsz�p<��d��{{�a���Fߑ+U�U��"�u�/]+>�6�,�}�x�h�v]�+`�bĈ�iO8�+h��N�%�mn��#��%XR�~)�WTW\�A�^�3�+ѣ��8y�ηX��/���6�U�+�]��7���qM'�#��!9	Xq�b޴fYHc��N�U`ȼF�����b7�L�E(@�Ɗ.��8�`��IT�3{�N7b�Um�ɮ6̼u�9]v��|[h7��"U�]����925�5����J��|U�����Bj�`��w�t�����a�Ly+�����+���i�ݘWh���յm�:�V,~�c�	j�X�Ca�7���y���S���d�k�� �n]e9��{��v����<MQ�qb�,z^\@���5�l$j��z�\׋�UV��/V���:f1k�5WlZAX*�E�T؛�/%�f#Ldc���z�����wV��+��t��/��q����Tg�M�]�G�j��!�乒�^e��_k�`�ݝ��$�{Jl�2���n&�5�1P�B:E^���e�V�۝��ѻH�oo��G	u�Cf�Pe/i��yY��c�4����kٗ�,��w,�yn��df5ps�F�aܫ�],��/���B��3��-�U5UԈ�o��M���������:��NosQ��-�bM�D3���Q��fWdFt�qwv���ͪ��j|���US�oGڣ�%�U��yؐ���f�L�j�޳��[)�p�ɖ�ESyx%�>o}}#��IqNE�'D��;l���פ|��8�~�u��|݋+ �z�Ǯ=z��nݻv����@��J�������8䢀�Ύ(����ΡCLiӏ^�z��Ǐ�v���=}����dgvq�ZH�6�I�{Z̒;pjБ��P�`I��t��=z��Ǐ<v���B@�%@��֩��M�w�r'[o�d沊�T�I$��SP�d*M4Ӧ�q��x��Ǐ=z�����Qd$��a��e��
9�ڲ���ř�E�ܑ�Rt��Sn�&k��I>��e���m��G�H�o��:�:,0��D^vwyigvQŶ�8��+���絧gd���NJ$�Ì���aq�_Wt�l���L��̸�m��Y�zt]w ge�q���]�㿂����\���$��#�d���Z�GLF'�h$�@N@S���ls]�bY��yG�9�'���x��2�)��]�|��l� ���BV�i�2]�g�Uܚ�|�s�P>�d�|�.`n��nQ �@�@�	���FH$��DSh��.4@.D�����DF a����mHa,��ȍ��`�?�,i�������j2H�F� *	"U�� "�"�" ȡ "�#��s��t�^Wy[Ǩ���5�4FnF��U���ji��\�(��D�ϗ�K�d��P�nO��u1̱�tz{�gZ|W�m�^��	��ĭ���j�͚f&�>��=�&�}nס.����<���I����.��5>���XPxg����D+&��V��k�:Yڰ�
߯�2U���}^�c���.�n.�P��'9��������a�S�׶u;"$�3��[��򶨁�׏��aq�a�S��8�����������3U�{  Ș���֞����Z�C3�;�T�a�1�{E�q�;*��L�÷��n���m�d�&�IE{!�؟wՃ������T����Լ|}U�IY�D)�Ɋgv=�`6v�	�,�,J��r�N8\�C���;,�3kM?u��KK/PP�\H��y�H��27�����Ab�H��Us ~������}[����
���<�����!��0.��O;�8H	���1�ވ���:ڶ�����k�!J.w\]��D�v_s��+,~~��|�)��i��<%2�{��C��-,q���ńn�:IK��n�
98$�1��*��3����#�J�/��B�2\݆d���qL����}�uUO�3��̋��	A�{�I�J�͵1��B'�_=̐W�5R�����j���k��/Vr�7y�7�Y>���J�2#hV��"��R�hj)"*
2
�"���
�{��=�r{#�5���r��I}(��tQ}w�xa���AF4�r��� �r�Mo-:�ɭ�9]��ݨK32�����߸�2.�!�៸���+����T_����f�r�c�o8b��ӯ[���2�OY�熲��E�%��.�Bxw����3��KD�wm��P���EL��}��S�:���q��*�
Y�̪�V����Y����uh5Rs�+��.`ρ������7W�2�2)W����=��zg֪�Q�����t{�C�� 4�`Ӳ�F>�i��i���}̮EO0M>�J�mh}�4<G����/�)}YZ�Ѕ��n���*��4E��͠�@�-��/o�0�Sڗl��T/��j�u3�tXi�D���ݎO@��)�5��HƂ���a��@�d��w���C���`����T�b�'(�]������W�Tz�#�"i�3 �e��&����B�&�}3��IJ(��No��E����\�Ș�Sܺl Ji�ةTZD���C�s$�O"^���Ż��N�n˽��/	~Τ��s�����u�6�ĳ��w�G:�����0���ģ�!��G�Q��c�^<B7r;K]�he=4>ĺ�n�k��]��k"����B�=)�ͬ��	Q�\\�X��ywp#gy�@����J��iA)��R�iQ( �H��� ,���� �H �繿�=�|�p�y������<x�,81.z�i<���3y�����=֨l=Y�e��y-�
���W�6��^��"i�4-"G<��J�����"S_�ؔT��<�/#Ք~�e�]j�Al'"�4Q���f|�7^oþ^�_�M���>�̹�Y�/�Fb�A�F���u��`����]���}jf���������O	G*.jX\�����y��<�v<2ogٱ��<K��	U�VQ�k�ܪ�?)��c���3w޺��/�w��u�yˠ,��.�8�c�ʥVvQ�~����8��oY�j~���ڝN0��^w'�#DG���^��M�}"M�(�C8�C��N[1Ab��v��g�D8r���ǶE��a��+�P'�4ƈ�vr��:��Z�Q�X�*T7�M�g9���p�e:��W��؉&=�׾x�������;}�!�9���8h��q�U���ZP��΋�%n�k�f�c�>��1r�N0-{b�l���P��(����}�Y͟���T�l8�3Or!�ma���hN%n�������F����Jm�\�P�/3!��4E���;Vd9*eV�]�v�F��O+#��[n8T�,2�Ѹ�D�1-�_!����aۣ.�f�T�]��߇2��*�yﹿp��� �*H�i��F�F�A����ȑ����Ȉ�
2
"Ȁ��Q3j53Q|�ϡ9�=���j��>?lb�*��	CG0�kL�
."�f�%�N7=!U:��I���.�m��]�cc�6>�21�����:Xz*cK9����S�G���0!�f|Ĩ�R&�oI���z�8� T 
��- �'��pu�g%�:������P-��"��%�!���4�3��N���5yyu��!J���s�;���'/����b�և��|�ܥ�g�B���
=ŧ71��zcjPu�B��Lw+���B|��<�Q��	��OT�u�3�j��A�RLXG���v�Q�u�yN�Iv[x}��QJ~���%��������g�o�������6�$����q&C�9�Uid[����:���+�֑��1,�ɬ�([��4*��m�|�9�;E�,Y��[�&i�}�>,zŇ4�N}��2�͏D&%�tD�V��cEMm�
~�j��5u���Hٔ�uF<�g*�[�o>��wҥ'������,�흒o?uĨ�z��m�7z�{�4w)�R�o?0�I_e���K\S41x�W�z�Vn�]>ݝqN��Ue�'Yh�x?�q8�!�������`r�`���|/:�����%y-59r��Yw������iJ�Yy6v�����K�|D�	 R?M"�4�-E�2�4�AE@�RDA	D 8g7�<�{=ѯ�^B����G^8A滁��7[HD��^*��$������c)�d�o�e�˞���y�sӌO�!�wL�n=֙u�܄��a�䗛[�����6ˡ�]v2��>��;�c�,3���[AF�����]��f{ԫ��k{�^��f<Q��&�t�w�|�� <;���Ɔ
\w���0�u�i���tR���"S�	�-ϻ)�7�'k����\������,c�k�)��Q{��C���vj�
�`h�vNSԾϟ,���?N��<���~�z�?�զ�� C��ؼ���j,[C��u۞��sc�k�@ ��3���0�ȼ3'�0/oe'c�z��#m(SF��=c���ǔ�h��<z��4�~8Y_�?�/�?>�^�X��Mʽ�,١'0���u:�ϭǆ\����~�E�	[�c2D;�A�4`���&�EDz��-i�gR�P�ة�>�S��>��kNJ�K�(4�fAp1�=s͹��{d3?�(E��N�e�5w�g>oj}�-t�n=3QLm�q��1K$�(�j���n�@��M�93�����K�[���j�U���aK�q��D�_j�<ldH�5[:�F�<����s.O�g�9��3�A(Pu�Ds�L�rA�g۶ƪ<���ܨD.���V�Y���e���+�(�؈�J�J�%uuw�����Q��* �$i��wuYU�WE]WH�$�2 2�2����Ϝ����!\An(�%�y�Bgv=賃�P/K#�X笨�g/��r�⺓[�[�����{�c�6A0��鉯@�t6Mw��w}i�w�Yϖ*�_���"���}Ʒc8�n����K>R��Y��	�
��0�|`�#M�4��w=��0[a��Կ��wu���;�B���ѳ�7��oD��L��bb�:	�N�Ɔv^W:g4yv�xy:���<�_<�/Eq��TlO;5����u5��O�;�[Q��!ן��dT\���i��I�1L���p��m�\���٥��#:��CNhCY{�ׄH�7W�Ȟ���v�O<5z��/iAc�˰L��]vC�n33���e�:�C;7�y��Dm熄� �#�vw����*�
Y�̪T���Y96D����:Y����$��W�^C����dRn�.8�,zU��)��n��Z�(�zv�d�:�ƀ��È݀F���<2tԈ�E�&�:�<]�Я��G-����j��K�-�[�3l6Ⱥ�t6�{B��Ć��u�I=��gU���n��m1A�їKM�U��t��p7���3�=��N⯤�x/���"���F��qȨ�I�X�n$�oh�y�F\���5�e��)�=�x{}�h� 1���!i�# H���
����ʹ�r��Z\v�K3�C~]5�z�NP}��)�O[��H���}#]$�{�m��Q���m\��ڙ����L\B�6k�}�0_�c�>̐pS3�l�g/<��  �2����I�9O��e��Sb�q
T�|��!=�Y��C�����M�,኉;�*D/_�%Rz�9Fo'"�<�7q����z^�"�3 '=�@Ot!�:��J,���j,3�6�+�-���<�����?Oz��tI�;2(��O���rx6(ڃT9-�h�S�x���-��
���"G��T�<�c�S�0Dlz���yu�;tx���t��q����i�9]|ݸ����1�L�]*�^= ;�'k����|D���w���ndD�[��X����]�m~[����R�&�EP�����:1�<���0��n8Ҫ����w�ܧ��S �Ϭ�����>��2�����o&�QLJ2�p}���s	�ѻ))����!��k�a������}�7���ʥY�~�cy�C�x���%8��)1TZ(��T�hͫ�S�>���֦���
��h��x�n������X{��|p�cFp5+	!F�^ww���zZ�4mi�M�B��Nbߥ����#�n�RO(��t����d��ފ�����<����<�\����H G饨"Ȭi�R��h)��� ��]q\wuq��wT]B� �{�ff���ʛ��ͺ�&���B�>M�0l���B����|g���o��H�R��{^�3����[�������̅���{�L��樅W���ފ�;�ب��.sQMa�o^*��8�:��O�Aα�6��\<��&��(�_T��R�j���Q�=�Z����#.���A��S��.���e����BH��W	}11er�&�iL��bhye�veo"�)��U�g�/�k��f_e8��,Xs�&��X�:>��'�V5#�zX:"��:lO^�n|�\�r׺1����i������%=w7�`v��W9�Y��l�w��AS-x��,!<�}�5e�^�*l�Pw��UwN�C�l�j�l�p%Y�i�:x������g��������/ƍz�|�
�z$��u�}5�Wi��Jȹ��U��]OԱ�w!
T�8�zO�����`�!�xo����������E�ۢk6D�fk���g���[���Qlh(���6�����0�p��4`t]G�_�����$�:A�J�7�&{uU�)�x��U�q��!��o%�9�S�%�y����:T�ktg�]�(���Qpr���»��=���%w��U!4�O2�.�˕�ّ��d��;DSK5���\</c�טl�D���wߍ��@M4�T@#M !PdQ� �QaI  �oEO�lGK�Ʃ�xef�0�̬܇�I�N!�Ĳ`��j�P�[�Q����k�s�a�	Mw�2�&��%�Ӭ+ö]����+��_��ً{E�Fg���2�6�,2}�#a�d7M�;Aq@i�d��Ji��4)>��;ˌB�Xu%]cݶ{���2��DxP��D�8�%���'�^|�;|�w�u�RqB��%:o]hت<���RŐ�s^j8�s�c�,�?�<#\�ZG����z�$�Vvv=o>�d;b{���5{�E_��^���ϏL/��M�,#�4hWLO\��hF{ݞ��x�}0vL*�(�����i��n��K����u� z0��'J0�$Ly�>��]��O �Ix���}�*�jW<U�������� �;�Ƕv@�N�E�1�gTsX��
tB�*�Ȟ~�&����V{z=%8�+��Ŧ�ȟ2y���wW�ݮ���o?K(�@k��
ä�!�ܧ�%��E������c׏|g�^zmG5�4㳲�+j�M�t�f���~��� ��p_U�4��>�U~���[���7�"~��Vl�A�9'�)���Ƕ{�n�=Hʏ/;�_�V
k�:�˨�5c-�aTw�/8���^m�y}�3��=�a�J��_nE*�xݥ����ZVy,wL�ڦŃ��Ó���V��I�b�T�I������v�=FTk���;��Q4��
i��iE��P���! ���o�w߯f��r~��nV�˭~?	��cC��Rm[���P���˰���;-�W�+��� �bK�wnn.�6�ξ53�"]��H?\ء��j{���Zk=���<;�����_ʮ���k���x6�F��kR}^m�yX���C��j}�C��ؼY���s�c/lq�Ъ)�m�.+ۑ��PK$�������:�tgO�:����3U�g�+��	,9ןC�v�pUʹГ�v�	ϖ@���%�zR��,A����D�xǯ��p��z���^l�T�a�B{d�-�dF�6��X����Τ�."	l.۱$���n���>����\����|'��Ô�����7~��E�	���3�Kf⫰]�˦f�%��{b'���#�RP-�-�nE�<�����8�rt����e���%���2T��j�I�x���_ z{y����KQ$1w"|:l��d��j��,B3�_��@A��>���C3��^��{�Ⱥ�� ��4���\��_ �{�x	�$�*lC�FS'jW�����p;��oj�W�����0s"�4�Е`�YGZ���r���Ì#me�K�f'�%�[x&q�3b��A�Oe�N���dU�Wu_IZ%�:i����'�]�g�,�C̾�k1Q��6.R�>2���[�o�k�V%J�8Ӱ�i=u�(�ÇoN�A�ę�Mq�y���nf���Z��[���;�A����7�IW<*r��ra�F�w�G�e��;���Ę6�쥳r�zY�T�U:�U��U��yt.um�U0��֮�����gtv�6E�}÷mRͱ�]y���Z*X7aV�e���V��kJ5X��lk�5�#p�j- �
0�f��i��v(�{��rZ��#���X���ǯ4�Y�-f���Y&�2��O��Ou�uPŦpa�{�Q���Y0�K,�V�ou�Y���`�7+��$e��*��B�����@RO�1{`����珒�6��gx���:M��z�LE����*�Ƞ[�i��K�����̬]�_;Ux�����ΣM��!+�G)wY$svX�lTy]t�=/1#vz�Ҷ�s�z0u�_q}22�^Zo�n�Vnc�+T&�����͕S����q�I�q�z9�K.��͸�.I�I�)9��cq]f��7U�'7�#7�^�F�&�vkZ�|V=<n��P���^���]�O#�~�-O5�e.Ax�$m+YՔUs��z�$H`��r�ܸ0����p�{l�OD�M��<1�'�3d��3�g9N�8�"�u1�9�����Ηv\Y���0�͚��d�C6�2��]�[kcҩ���v���U�&z�K�-�c0wV|u�D1�DT�����<��:\�T6ޕ��h��n���wbV���=H�gk�9���s�>�t�c-�}^�n�򎮫0ť�3{�������9{o���]Tf�PT
�ǻK�,��x�#�M3˶_Z�|�Ӷ��������Z�fw����+]G�Q�4�,���o}�P�m5�/���]k���j��>�N�j��-\yC��V��ztR����]#w�#{��ŝp~�n�j�e]�2�t
��� ��<pV�E�8t"�&�r�l@����ӆZ�bH�զm�w�	NA�����4�mhq�e�a-�r鄲(U� �ȵC�ɓ�L��9�*/
{[�cA��u��Z��;���iV�9Z�8J����]x�+
���\�ӵz�z��O��OV��l�p���a�d��J��ɺ6U]S�KA�Xևl��J��Pԯ��_	���y�dz��We!ڤ5�x�9�Q��JڍQ���a�FKi�0އ4�H�5���r�����L��-N�(����km�Ek8�[5ontlF�TJ�R�G��~�)�wŝ~�n���l��8���YtuLi�Ǐ^<v�Ǐ<x��צA�����D��^h.�T��D�$tӦ�q�=x��Ǐ�~w�~�/�n�;(��0�s�μ�Ӣ���qj�H�"SN�q�x��Ǐ<yߝ�߷�Y\twIw�h�N��.y�L�#NÎ9$�FF�Ɯq��x��Ǐ<x�w����}���QNI�AW�$GR��%@rV������o���ﭔEI�ݞ]�q�q����
��*҄� U��p* �(��H���$wIqӝy�b���s��~�trw�"Q�Z9��;�8������^դHfA�n�.f���^س����s�m)Nw'�ܞXt_ ���	�S�N1@�fp���&2i�eF�7�a���7]��2s�k��c��쉅�Ks���t��ɵoq{���
������J�"ƚDi����H� ����:��h�oƺ��uղ�Mlv�1l	E�%�Tn)��b�����]خ8Y���p�C���@�[g����\	N�*T�S��R�Ξe����7k�Fk�K��ş
6:<:r"@��g�t�==�"������Ů�V���8�v�uG^��t/�of��ބ��ji����@��ǉ_|c�ݙ��'�B2�d�Y����ꎦhxw�.��ܨm��{���0'kLz�5x��^�90�h�D&l�y��T�21�Q��{����^m���������8ñǠI�}M������^]�Z��2"^�C;���Ӹ�+X��Č{�_�S�dW�;?�"R��d�6�f�zn�5�O�OR�ڧ���6�����4l	���ۤ��[�'�M��lP�wF�y��?L�0ƅ�D�oQ]�ˣ ����w>7�p�d�dp=�<%�]���B,nPg�bݞ�W��Xx�l?��"J��do������*Ƈ�e���1��O���yL]M�=�%�����M� �]����<�a�9��̝v0¶�"�]6���m�sl�����k��@�	Բ�[�7h��]u�P.�L=Jn��܇X��[X&�G�L��v,9�D�9RG#K`V����g[�1V(�[h�D&r�q�����i���(Fj�������
"�k�{�>yU����(y��[W�ٲ9�,T)=�]�(�ǯ[ռ6[�; ^�0��ܞ%�&�9�
��BJ�Ϭ5c�^G	M^�%Հ����%n��+ͱQ��9�<�{w�nV�U՘|Iז��
������>��	���lB.tsıOz���F�
��qP(-,�Ч'F.m�Ε�\8�o@�}a>ǆ��A�	aq*x�'�>l\�O�0+#�D����>ka���/m�r��p���7���	���M�}"M��P�
�����j���Q�S���݄�]&��%���->llj�5���Y��[;�h<˷��X��7r�6/)4���>�~�hN(w:���ߕ%ؗ���������ݦ<j�j�|���̯�j���D�:��7��r���r�*�Cb�n�`���T?�Fr�|}�!�1�/�T�)�ȖX#cʆ�tj}�X�^�z� �=v�l�7
J���i�z\��`�ߔkN|�D,��6�/����~�{x�ƷWν�ݖ�y��� ����[V}�*���zT��/h�w�#'� �(r��7�ZF'U�ZwUm�f����F�̫��ز���j�Ҡ��w)f�Rb�UZ�EHÈ�I��MlC#3v��ɉ�cAUk,�\[w8�1���n�}(?M*�H�DH�B4�AVA@�BD6t�w/�Q�ʨg�����x��ص
�6��n^LH�?ig�>���OڢW���C�"}�
WU�I��s�/^�D����do���<(��؂ێ�+*-�����s��8vB���:d���[ѱ��mw��N���F�F��X~Z����ޑ[�C��v"���}+"�QF#�#ZZ|E�H����CT6��y{���z��p:���[�@��B�;!PJq�{�W��
��Ȩ���f�R(���*���;2kn�y�j�L��..���z`y\��g����lbD���u��9�c��Zl���W�L:�̓\b���Ɨ��
mN����,3LK$�
R��� �֘�u�o��V����Qg�\3�P�(l�=� !�1�~!�;#�}���9�x��EX$��έ[�x��Ͼ��s��Ѹը���ŋf���מ�m0���pe5�M��:ϝ+���W�o��D��˻�.�@\L�~�F��a�@�Yz��y�l[AG�Ȅ��js����l�bۉ�k�nKN�BK�y��7���2��1i�g�H�b摴@u���آ���@�]�3U��3�ŉ�EI�ɸ�Y3�kR�Ǉ-�TE�FwC{�E]�6��;D���K+�,����8燇�28D r_CMn22
��o~������5���;`���^>d��ժ�f�.�+^�GMXD��Srn �>�.��{������
i�B�iR�� b*��΂�1�D8�C���p^�B�=G�la��C������g�ü{gj�5��dżʧ��I�S�w��9	�؝uB`Kk��5oB@8B�O�Q�UR2'�㩠�vs5�
깷xx� D8B"
���� ��G���Qi�/�+���1p������k�{�����ÖR����������A��E|x���߮afcK�힕�^լ|Ȗ������ܵ��k�>��v�
<B�����3%n��s�D�?Z�z��G�����
w�I��&]���a�qjW};�;3@xH�Cg�����Z�G�\�ri~:9��הű�V2<��R2�e�Pi����֞�<���6Dy�c[�D�_['lj@���7�t����g�S�}�:y��r2o&�k`!�Tm�kV���]zw�"X��0�"!�|{q�2=��E�,�!o^ KF3�sj�_Rc���𷶄��Muk���|�i��<��ɲ�g�^�;�_�������DL�roV4onЂT͞ ��Eh�CW��׭��Dj_���]��1L��r&���k�>����B7|9S���{u��F�e擊�Ѱ�V�qf�m'-F圲�έ;�IS��oot��8~ ���璉i��i���1��j���{�f���q~
�u<X�xe��~Դ�Wc�;P�(�g�����9�=�#d1�q��jwWx�6w�.�^Jv=q�o}%Մ�^�%8���a>܋hU����	�p���ه�WWYg��j�ݏm~�`@͞�� �Y.h_A��y�#%�!�I�"�Y^���R����f�@s!I�	���m�2�ާkَO�b�X��b��m����:�g��g����މ� 0t'];���Ŵ��ЗM�fD�_Ra��&�#����.�y�5%?c�M����"�`e��н"�و�����U�2;�8��*y��i���C�_��#�.G9ֵ��q�p��Q�1�,�s��ǡ��uxT0��F
�U4�z�V,�������:�
�^��*9��� kW=��s.Ġ>�ܨ@���V��[�J�3fX'j+d�Ƒh�lzk����ÅʇE���W`v��C�J�t��07�K.i40gy���C�k�O���&;�	/C�;r\g���<�zi{�Ǻ���F�SXU�#��X
��\�[09߆�����J���ν��H����I�r�ѹ�yG\�8�`�/������r������&�(ha�4m;�Y͓��J_���=fc��/�SH6��Ӭ�;s;�v����xz����Х4Ҵ�B��B5$$ d׹��e�>s!��}����4/�@��d.�<?����޼v@{�	s�} ��I�l�q�;��o��g���FH����C�3G��>k�>��=
�8E|�N{b�y<~�?fgh��1ϩ�#�r�n���n�Ј^<3y��9�WR�0Ʉ+����軚��N�h�٩�sځ���֍^�����}��N��yr�
��T�,���K�p��х�	�f�U����[���zN��և�5�-��C��,T):��^����oMV�Ё�eD����zA�Mm����|�5�Nw����k���]%	�^t�P.�f��^���E(7U{�e�h�g���Cd1�\�
z�Q�^D.~\�,S�yc�Q��xJPۃ�k��U��e��U.� �0q�^f��2XKL>�+�*�.��]0�r�E��T*4�I��2��6�v����H(��-A�������'�y�Bm�0l���Q��N���1�֩K���v�u��t7b��XJ]&�~B;X[�2�pZm�������"�?nKU�����V?�[� ��6�\�-���z�a���n���X{�!N�ڠ|4j��<�۹��{��+S�{T�̭��k$����bT�;��&匥�լ��6��z�潜�=�o���I_`c��Bd4�%4�T4�T	�=��h�;�{��-��w���ڏm��'��+qL�ǥz�����&y{���]�.��F�F��*�s���^������F��s�\���U��܇'�~��6������o(X�%�^¸e�� "9؁��صs=�n����|ޱ/���m�[(�Ny�{�}8�o��v�<�K=�y�'�v�0g�1�W�|�~�|�Zs�Y	~Y_y�=�BO�1�KH��6����'� �xb9�y�ş[�t�<�</w��^��ǉ�AX^E��%M�ؗ�K 6WMw�Kk�l�w�OB�o���9n��f��٨k�xƌMDT?VD��B�ZB�bja�z�N;���=�*&�3I�nn�����yBk6y�5 �<`�e�f���tR�5`Eb8�@xzF-]��Ԯ�4��*��zk����U��o�9����XA�d�C��7A�6m>53���%1��6{~?�^��w��x�(�hz��q�b�#BϫЊMv4��c�}+�o�,�}�/�mEM����=h��:�fq�`]��b .s��w�Z]�.7K$�R��T5�p19�G��/�fT3��Y-��ZT�qn��+l��o<3�y-�t��/�w1;B��Q�A�+wYVv1=�tC�8��1�ʻ�Z�Y�%���U�����Ӽx�=/:Vw!L;���rj�gҕ?������hx;{��v۸�2~�@��=��ퟞ���y�)�5ra�u��a\��uo���� �(��m���{K��u�v;�L�I��:�O�p�� ���JD��>�8G��(=i��]����c�S�V���D&�c�EW0>/q�eӰ��gF0�
=r!6����ڕUx��n(��D�⣺]��(z���R9�tU}�dO��t%N@w�*󕝊~���ӓ�������N�{"TI�{�Ą���Ń	�?%�I�߼�^]���E)�g1u���-�	<���`d�r^D;��.ţ�{r ���Ic?IN��L�}9쯳�i0�gSٛ���̷ڙo���w
]�>����~�za����ۀZ�]@ds��m1���j�*�L.2�v���_�_��9�mX����
���75C�"�̏�w�2##-��ĺ1k�iv�Vג���@~�W����W����9�А���C���Wy��g}BL(�����lq{d6<Vk·�K��<`�%
`s�VWA����8��n �����l˱�ry�*b���𤕨�Xstv(�օ��H����'�yf��R[B����=����U\\��7�TW0��P�t�f�a�gU��\u�%u��sc6�9՛ŕ ���Վ�/�[���|��l��2�4е#L��4�B@���n�%q���{��y��К�&����Q3>/�i���omκ}f���7��tL	��H�,�Ĩ�K�*r_�-�1dn82(�c5ؙ����oU!{')SqL��r�\<��>��nK���c�^�2�'��c��_�L囝��=�s]gN3� I�2b���cG�.aϔ�!��	�Y�e�5�q>�5���N����rݧ��̻�?�6=�6|�|���ZB=_a����)��C/-�Pd]	�����;iw�-��W�\�!qLZF�s{�N��APR�S����,!nK2~��g���3���;��%�7�[�N�g�`zcAu�S�A~��eRc��Z<��z\�ds�W;5��;Mk)�پ.��e���G4����&�-�2��N�{S��q�e��[":����Y�!w?zk��V�y^��0{�r �%< 3#�W�-G���5�i�ª��xj��.����;}�����~1�ֲ`[��?E�����2�0t�>�	���0;n4��� ����F�Z�
���3����UU��i�=�����q�Z�r��	�.7U�u�L�Ke5o��СU�����Q�{_���Gy�*��JPJ��7S�2�vrt��7��u0gՔb�WQ}b�����"n.�Z���ڣ�Y��OO$A��Ji������2o�W>wy�c���?�k��|ά?
�3��F�����@&�8��H<e(�����D�
9�7�����k��1��Bڝ49Z]9�8 �
+ᯏ�gc��X��u٬M:��$T��n7���Y oEx;��1�!���1�A8��;��L��r����L���f��n�p6����/�ݍ��K�o�5T:ݒ�{�[`�=hK<=�;���y�F���QY�}��$U�/1���4*<�.r!���D���;rT6�ze��ƽ��pP&P�.$k��D�\"��S�أ5qu�R֠K�v{��7Գ����K�Aͨ�م0�oҌ��"�G�t����K与��P��0�ܜ~D��Ļ��۰1����_�2�����}�6�@���:�΃�j	�nZժ.TF9ԸtGr]r�f�z�k�Rl�4<|���������y��(�`���W���)��#�y�*�~��#~��lr#�y�:^JS��B�F���{���b�@�j��aO��a�rDe��)7*��H�v�e�f\w�f�0^1!i�Am��MkN���f�R{!ʚ�UH60��f�q�&�G�����>��4T���`��<�0��-�泇5*�%N)�x���ʘ��\�*Ql��&r�~5��;�u唧K�:tAna�0�uJ��Jt�2bO�ۉaT,@���QS{X���T�d׉Ҹĝ�0t�A�ÕVe��[��ׇC�Z�}d;h�w]k�w2��ð%��*��T�S:�����Qƍ^�6��[�ll:�Z���=�,#���AGjf.M����Q���\d˾7K��tp6XՐ:3�l�o4���ꋉ�0���dp�Dc喻��T�2�,nY8�np��I���#�`^Ĳ^�;��9X�J뫖����)����Zf�PԂLͺ�ʴ���!e�,�40:�XRTj��?f<Pb�����=��B��S��Ø��0���8S[U҅�����|�o3a�5y��"*���'gM�s�%��Y���:*vK���m�l�Jٯ�.٨-�����e��n툽�}��!U���ɠ��8��͏$6�/5**��{�D&Q�էx���+�b��.����r�H^��4:5!�Wםۓ[�-���!U�wҜݣ��#"���^�D���M��YA8�j��5�����&�6t�_���3�$;U^`���lT���L��,�B�*�:��.����Gdj��iÂ��i�{�ut�0�ޓ�(F[�1x���r��2�V!uA��ӌF2��r4�%��ņ\�D?+�׵���y��ިRU�J����Uu�u����x`��CL\[ս.%e� g/!c�0�X���OX[O�T{�k���T�f0��[V��5}\���q
Q�4�^_3��t�<��_L٪Cd�C��W�:T�K(�Rc}ʟT���Ԫ[��e8���rw\kO�B���.��/F�2:�Y���SC���S���f�FU�3y�/����G���5�B�TI�:�8�W�;uU9묜s+cZ����,�bf�o]�+-sg	/0�hl\��ѵ$�>@��I0d#B�m�?u��B���.�G+f�ҝU�kƨ\$���Ԇ
�Vܕ��C����nk�1�ei#E֍ۉN��!	��b�к�ps=�
�˫�K0kCt��9z�-�X'�����Q\hn5sCiΒ�5]7sD9��f+l�ȓ}��{a�UV�����j2���pot�՝��eɁhw�E�Za���Eu��T��+��}�,;U�e,�KK����S�J��ӌwtR�9*�حZ�n�WF,�M:�+��+c~П7i�0{��v������׶�.;��I���iGq�W(w�9���n�=q����Ǐ<z�v.ID˥�GtE�9t=���D�$��I�Ɲ8�8��׏<x���ʊ�!$�%��*;�E��pR'�H�(��ƚq�q�Ǐ^<x��Ǯ9BI5
�"I$� BPttupQwC$$�M4�8�Ǐ�x��Ǐ\o��㭱�Xa�.J�e��;��+,���:�#�9"�.�*8�Σ��8��Y�]u�E�E\�]ͻ�/;��(��ó��N�N�Ȋ������gG]��㳎�;*8��.ˊ��,��N�PVr�gegGte�Qu�Œۣ�8�. �:�٪2�mv��":������%��R6[n'�R-��-Ȋp�d��,��B$8�1�<C��6Ȉ��IRaX��Mu���<�J�a���fe�Үi�
/��sl���͹��d��ּvm��5&�q�����.5E�#EJS�!
�QReDR~��	"N�fD� ڌ�\�P(��f�h$�DZL�Zd���d!��~@(�ED"�O`p$�p�_`�񠦚h���i����r�>]|<�S����b]U�˧�����l�ݶRen*����k�{��?@��׻�(Lc$�� ��>�f�0�\�>�gO��������l�2#���np'P���U{P�9����+��;�����K��EW�&�0��S���ዺc�m�n���[���jw�ޚP�cD��#�(=�\z�x}!.�+ǳA���]��=C��m8ؔ�t��5�_ka~�_��=9����3MQK��B��vg�|3�Ya=BV�X��w:��ӽ�G<A��XM��3���]�bW�_���1-�^��)�E�oZ�V�M�y\U#(l[�)f��v*��dc��n�$�8���y������to����:�q��q��fP}]�[5}lDnnI֪+�TCy��g�3 �<� "�!���	�C�ʨ���_l7G��Z�x�آ����@�~��(X�yopx�����;ק�#�ĆE�/���VHl]v�Kq�D��U�Yֹ�2�8�rhI5~�|�b�%��o�2�?`~�ʕ�����'�v|�u,�z٫���YQ�r��5��k�ۗT<9ZɊ����d�"�U�++V��� Բ���<ڪ�	ŹiN��e�6�l^Y���!T�u�+�U��k:f4*�%ξ��]�bp1T�n)V-^sE�ܰ�5���T��CQ�4T�4P1�4�L>��K4����[�"<�[�ۘ��^��g�3��فN��!�N$�<H2��X����Rg�5n;�n����{�Q����f�Q|kl˨P���W�X���z͛O�3�o��ܬ��ز]��}X���4׿��@���;���g�ŰF�s����b���k�>���"���ʈ�4���X:�+�ŚQ.%:�(`�a�"���y���~��db���_��ڄ(�X�W��{������K�\^���TPZ���|�H��A���!�r0(ۅ9Κ>�-�Q�q��\��d����N�"y�P%��&����fzd_����|���5���������3��Ծ�׬��5y���wJ�_�D��IS��3��)�OO��<�������H��e[b�.��a�za�r'���R�7��a��b���U��36j�ǢXzW��?N]��u�#ލ���x i���)SP�Ӛ����*��s�Y����K==]	��X{e��u�W��/�X�� o0�[%�_�~�A5sA�[����~B�׼���(JK��-x��5:ee��F6	K0��UN-ll*�� M�l�-�qq9{�4�ŝ�Z����M�:5=M�7m�gvV��m]��բ�9��E��J2z�Ne��)�&��cĩ1�Yj�]�;&Ik[��q�Md����G馚hZi�)���2
*�㥚��|�x�ν����V��9�2`p���S��v�TmoX�`�n�R-�sLζ�D�u�k�C����/]�|��6�Gt� h{B�����B"�.^��W@�ө9��;�y^�ژ�"��Zptk�<P�"L�0�:��4_���9���Ŀub��{���C�{��Lν�'W��f'�1Q�NXu!NĻV.g5dlnU_`����*�6A�fË>��u��Q�G��������!W��,��&a.�E�e�K�Zt�]O<F��q����~����J��*����{�T}6�>s���x��x��fj�-�;ٱ�Q���%xV�8�C1�CaDK
Xt������=qMk�'�I�&�wy�g�z�c��dA�EH׌�Ƈ.�N��S�	~���?�T72O���B{d�#�q��xi�-�w�9��������b�)L�	bۜj��o{ܼ�����a�y:�B�}a�	�ن��<w/�(!Q�64���\��]YJ��RS�� c	�m
�N7��u�/n�/�F/�����>X�l֭�"׊|p��O]GOgօnk[cx�d�a*,�v
��S�i��Q:n�HO�l�%.YB�Ƀ0mʨTU&}�:̧y׉����%���]��{_�T����h�9 ��Yz��hKR�j.C�!>�y//'��o8v��Zb�x�����E'��?6�]�����;J��x�X�E��_�ط��~���^ˉ�"��ub5Ft`�0&7�UH�ȃ���A��Ω��^Y7�$���V��[����oh�~9��}�p���@_8���D��e�
���2B{=�%�DUПR�/t�Ŷ둟jW�����e@Q3!�֨���h6?5���|�����*�9r�Vv�� �@�QaAgO2��Z�G�e�C��ڞ�(|��-!���yԮ��/���������}�!�v`N?�hO�\W>��T����Q�%mN�{K��^��K�;�vX����qo�خ H0e���=0N5<W�M�W��8f����s�Ϙm�>��^�>�y�UD�5���������x��,
�c}2��#��]3�0z��Pk�߶�����1���aZ��L�zD�d���^� ���g���$Rn���s�b\�;�5,�6�46wr�i���!dJ�<�A0�U�/�E9����a�4 ��A�7���܊ېK�7���T���lv[ow�$����&գ"$4Q܋qC+0)8�W�=Դ�i][B��8�`�r�EA�h��f.�\�Q2��L�GRU�i��B	���VR�����\4>�7��(COunh����������~6�Y6I��Pk@y���3q�|�Qd+/��|!��r�c�[i��тk���eb&~�۞� ��?>�C�{��4��x��s�F'�'H�4>(sE��P��Yn��NW��U_Eǂn��&�#��σ}\dJ`?���]�Uq/�\��_�-~��l����+�C����ٷ���*K�這X���c�q"{e� �8�g4Lg�Լ�),�R��B (��.6d?u}�z��?�s��Jt�sx&!IT- �m�$�߳3�Sp?�4��V/�K
,EIz�ż��>�P�8:�����}=����z�8Z���|��1�[]�A��N|��=C��[��`�L1�C]!_Aw���/Y���<�Z�o��3i��7a��`ۖ�p���Mt�~�Ϸꀛ�ud�h9X�M��h=q(nV���g��q��(}�D�]��q-�Ez3_�:im��g��Nm����A��0c��T�0�y� �����똠U�@�s�5�p$v�x�f����v�OK���R�RnN�-��4-~�1-��D�݂���ek�`1=�����9�tOv4��Ӵ�f<*�EM�M�L5dS.ʡ��� G7vqM(��o��.x��P���Nd�CWvy���2��֯��/oV
�ݽ�ɋ촐�4��-�ԕV����� �E��YN�d,�γ�U�D�9[T$��{�����aFw�U�+8�~��@�����GW� h��+���#���ֽ.�����9�ON��',��ƸUڥ��1�3��k@vp,C���2^|�^��;@���|��~ٟv��,JVGc�2����@8�z��D[sU��*��^��>0���p��/���J�J6�i���jי����kމ��`NF3��O��za�Q���闑0u�C�(x9���WM�W.��T{��j����s_&��;��(w:;���فAܾ�6)ě2c7�\�#]ھ�o,c�Y@h����?�>z���C��d�[n�C�3f��-����o�se�AOl��#dS�hqma���Ǧ}�p�����q��iyA�Bȉ1`$��#T�݋S��	l'����m��Ƨg6k�vf'��r���=��ڝmw ��o�%52u�^��y�ͺ�o(�eQB��Yca��PP�$P�融��
|D�-h�u�P]2�t��i���u���~w��R)�iE�3W��z�gl\G���#�3S�P>)�w;H�Q���k(�G1�9��j�ԗ���B%�l�̶͍X3{H�z�ֻ�8Nv�G]̚ݺ͐DZ⿺��,U�j�(����+*�fM� �vn�ڗj$�L�U2`Z�ƪ�&(���<�fof�wY�|���-��0#�y�w��s���uq�2E��ޚ4��t����R��Aq�vd��]*h��wV�����%7W�,6ȸb�C���s(~-���e#�s��=�$C���J���|^�a-��F����.& xe;��}��
���_�t�/��t+5�Rc;yL�S�.�	xw�|ga3���f �|�ũ�H�R����N��
{]�)��kit{]u���>503^�1 A�t��.�?/�,�NAA_�|�qw�A��Vյ��Ѵ�����쟬x4�|�������D
-�A������a��s��É�Kwj�p���L�lڒ�u�~�a�@�MsH/������p���E��ϟ�jU���a�-�����ԋ����Qg։ޚ�3���Һ ���0���:j^n�eg��x)�h�&P��*U�L&���2���	��$�K�2=ϧ�`�9��l{�*�8[���5�Sq;C�I,�x>�~Q����%ק����r\`܎%�Ԟv3�T�q6��\M���"�k��M*�5vQ/�r���(�]�*�R�7}�+�j�h�5��'���d���pً�6���j0�xMKό�Ȉ��a�0�I��d����8f�66�iFیG&{����ߥ浢W��c�s���
�Wz�@w�t����E}�ı� ��{�_L7�%��n��Y�9ԑ��h�v�3�h�����t@�4WV�����O�:k�C�~�fß }|�"�`���9q�l������=�h؎m�S�X�T))�a-����z���{Bzm+����;����h��t.����5����j�.*���tSyHO��{�*ȡXMԙ�^��d����f��Q�lIw<�����Z��?SQ�7��fofʤ�<.�y^�]�u�1��2��e�CɨF�<�;�� �{`�z]�6��ɸ��~�jU�����)ջ�Su��p�Ƣ�y#i���p��ޡ��d�s�n�2'���	��	�U��'�������r狤��i�HN��܇ǐ���`�5@L��B�
���u��2�AI��[{�aw{P+�Ӹ��r�B��i�ʵ��, ����
6�!��D��������&��u>�٩VX�ӁԷ)h	���j0����ҵ��A/mr��Jڵ>s�.å�H�5��8����c-7*�Z�&����P�\J�-�ؼw=�c�m�����P�wn�\Ǎڕw��&>���	��ad:�Am���}��B����Eݑ�s�cDÈ�T0��l	T��b�3\]ӫ���kb�ϕvhgjl9���>>�//��$�z���Y�ә?��LT>*�Bv>x,@	m�qs">�#\�.���
��K�<�߮�s�^�T��:�1��}�Q���C��C�	1��9�R)�L�O9������L�#�9�o-u����4,� 6���W�'5ӯ�c��b�lTdO�)g���8����;���cW�iF���|��}��BT�� ��w,�Ɋ��Qz%b�F*+�m��u�`܌Cp8"�@׊xnW ��>�,�9���������ۛV�U��%��w����M|�BW!
Dך@��yN�1p���-b9��I�'Y<?o�{�L���݃���㞞(R�B",b������p��'���H�yL��Lr(�6�r��=�U�����	{g`�"{d�d�f����Lz����^Az�[�.�k�t�x��<�5d��r�7n>"<24�F������dh�'�4VyN�l6��	�yz�G�y��l�NE?X���٣F"-�(����?<��D<����S'�`t$3^a>ͩE�I�S0e�Vq�w5��a�]1޿M�(�b��_�*������(�  ���\���r���S�Qq�DH��H���;�Y	v���3&�[��l[V�"�g!C�F�2���:�v� �:����� ��'���[����\]�:fak��x�ӫuȬDsS���#}:���muP�Wp)4��Wb�or���;Xrvя�c�W��{^��}��{U�x�Y�T�t9�]C��r��ký4 ���&ڧ6r�(SN#Z�Vv�����	n���N\�(���OC�zO�ܓ�L�OI���g���?��u]��E��`���#���f&=f��V�㐘P����`��f mQ��Q�`���o�G1jw��gZD�(K���A�?�C~~a�W�3�߰)~4Sڮ"���k�PKܽ��Acl��*5En=e2�i�����d�7�P�g¤p;��G�m�[(�c�?��M�F~�@�k.&��ݫՎ��Ƴ�^몿;����y�U���?��:o�#�d�e0�F��T�-��Z�������i��:�����<l��K�N4���/�M)�q���("����'�9&��_�l$K��c��q�$�6{=~3#�*"���D���@{އ��{�Ss�U�lvN�~��0��̊��s��k��ɿD��!�zz^=7�c�M�S�]2M��2i���1��xH���;*~���D(p��
�_�%Z������6k<42?xx�.l�!%`����j��c#>��L�f=N�)��-�D�%�y�N`�19�Z�R�6��*��l�3']��U��N%��X�k�r5l�[��ّ��j�t2��ʦp�d;'5���v�!a�{ɃT��6�?��C E������]�RS��p���L�؀���an����ڌ�j|��n�,8�6hΗ��Y ��ډ9;�&d�:j��T�ziSH�
co^����8�D��e9�Vxh�&���d�^�p�I�ff���g
ʷlK(�Ω5�3��^IS:���
�+3)C��R�Fl�Ǿ�;�:@���"hS��u��7�Uz���hge���-���̳��CCO��ᔡ��-�𓩰����N�
~��U_%�X��Z��Zͳ*�j֣RԌ��n�!��I�hi�F�6M�@ԍ5����̗c	|кґ���S����g_c�j)��֝A�����)�MR�x��p��2�9��t1��V챗�!�G���k/R�[b�C��L�.�Z��U�(MkM��3���W�y�B��~�o�r]����GK8V�/I74ud�ܪ"�rޜM��Jn�靇�.�ӵ3.�
[�6�<bi6�gn���Q�9lט����	3-����=ǖ���a��(-�\���Us9N+�bB����YI��;ݗuYp1�P���92R�	11y\�6��&;�S�����Xq]�� Ƌe��ݻR�`�!�Q� �!kL�W��2^ ���U��\�/�����ղ]�^����JK���a'.0���&�]�v��a�O4V,͵Թ�E�ty.�^pF�뺬g8u���a�J���6���-�Di�w����;�v5���.K��t�D3���jv�b���@㴲4+U�̡wch̐��2�І���I�b�N��(FS2id衂���o`���5�Q��������3D�*7z���
6�tLCq�F\���UX_^�n��ε#���f�V�ͽ�zv��i�>�l�KS=���-Ÿ��4� !���`��u9J�Ӗ�R�&���i�ˌ$��
ۘջ�OY���au��1U��FN's��ײ��H���46�
<"�{͝ʪꕼ|:c���솆��;�M���j��U�f�X�N��Ү�o��2��#j�,T�u-.�-��$ ���Omd�{Ȫ���q{XgT�JLŻR��a{�d��Q�u/%B�kt�؋���AFV"�g5�����$5��<�&\���D� �H�jQ�0P��7c�����T���u�T��;^�x������LKݵ�5��+mc�l�D���=;�U'��r�i�E[��z ��W>��ٹ'j�����|�e�?X�BV�.?��e�k���{d�k:����wy[���{\ػ
�J�Li��ǎ8��ǯ<x��ט���[;8��m�GG=���Wgetu�nݻ��q��o^<x�������H�u��Ge��C�l�d�	��F1�N�q�x��׏<x�9��TB�Td$*)%.�:xj��l؎�l�EI*1���q�x��׏<x����W�m�m�vI&֤���iݒ���7gbg�gE���(�]�a�[n�N��G[k�+�������Gefgemn㳠�:�C��f���Zl��ܜ��gXX�t\O��Q�۫,�������Ȼ��ѧ\wgg~����vQն6�wmn�ʲ̩ʢ���V^�쎊�l�f�d�g�q�Sl.�Π����Wfq~�x�Y �G����Dv�]2�T��s}�a[�﷈'����wr�j�37��|
�O}V����fڮ�u��ߖm�FX�1�~����y=���.땭J���������)6l!e�����0��O��&�|��>Y��,:c�Z*:��cl�6�]ǩ޳��~�c=x[ռ'�v`�����@#���~��i͵[�V-j@J��6�e���ؖ8�(�t���$��aތ1�AC��#�:u>#{���^>T�{e�Z��%����O;�t^z"K�JE1�&���=�r&_P���0�އQ�߱x�'yq�H��?�����`��w��$�Bb��Ww��ݲ�\�3���E��h9�2�9�����2���v�By�R�"ߙ��	��()�>/���Jw���H����e)m�m�X�	1 {�瞐�DO��G�&bO�%Ĝ���%�{^犳>	�;�v9��[���T�~�u˒jzc��c���������P�M^ˡ\�
�7���D�ގݯnPթ�"�Zoȯ�P���s3�;��'��ރ��H<I�����������d/�;�)�l��҄�d,q����G���4�r/l>+׬���
��?~�.ބnv�	���3.![
	z��Kj��uGGM�{��`�R�le�'\ѧ�F���r�}�eF���Yڋ%���fQ��6�d��/�e&����ǖ���ʭ9��oR�kUN���b�C��.Y�U�(Jɢ���,��rf����;��Ւ��_J��^��� ����ݭރ��iǅA�]	@�J+���H��dm�ϹѡѮ8���@��D���(�RF�f��񎰥��K���Íoy�.7篐C6k�oL5�0~:ĭ����3wO�N�n��ٌ�J$K���-W�|�5F�/�zT�&�B]'��˂�,й9�/�)�#r�6S�dS����00L���!�Y�<S�,TS@W�GSn����9�ዚ�u-���t5FD�����i��l�+f@St�{���!@����*�(��ְC2/_���$;�qtե|���˧n���	��~c,'�(������n�M��7���������C+�{3���"W����R��)�
Ī��/�	ǈ�Zf�z�Bv��S-�'= k��{!�<T�0�f�b']�"!IOMq��+t��W�յt5sb1�5SM��މm.K��;��[�W8��T��<�_<�/�:��fY�dv�o6��
:^����_{����jc��N�#���p"c�6���V�/��j��g�����ɹ�\�*�f���5�K�-�T�\bJ�e��6T��g��V�FM�P���j�(]u.�q�z{�l�#���9_��+I���nf�+�Y�n\+:I4�X�y�-f�%�B/5���z�eΩ]�T��x�.�8o�x���~ ���
��е�V2̓I*x����3�]Ė�]�5ͬM
�\ �^�h�Ē�Fȯ��L��8�8�j+��H4'!�g���p>�Uv�P��[Ԣ�_ O%��m/t���sQ��E�~n^�i�HO^�>�]�m0t�16���c"��f��]�r_�m���Y�W<��7���\ݧ;=@�ND�g��W��"=Hg/<���� �{؈�NP{AyF�ǥk�PH����}�n������W3����y�Gt�|�΄��<ͣg�ć�y�fOr*��i�jT:��z�_=&�q�̪�*r�!T����X����/����9��gA@x�	�;�:�}�f��le�qn�tuMY�sT�e<�K�d7�uASfG�
�x�lO���O��+�%�4g�d[4�������V��|4ά~�ε�V�����I�i8"-�^)���G���z.0�G�&	�PZ-����6�_;�;������c�@����E �{�b{��HA��|�x��.c�A��lzP���x�+���2x,�
�k؝�@i1�m���˝��Y�{�l͖F|�@S�NE��{����(��,��Q1�UZo ��L4�����L,籍ΟnH(l�Q*R�W������'[5�92��I��"�e建6�S�z������V�[*�"�n�	Zhj!�/Fm*����|@����~���qY-+����5��!ך]�[%�"<�=��nh�q)�F�	��"S���Ծ�9X-�Sx���j�5[�l'P��a:h��}@�z��>�[c�ݽ�ubl��kL�z��j���˘3�u��s�� [�E%���@G���'�+���^�T\�&*�q���G�hy�����ģ)�?Es�v�} H�#�;�8d�|IU~F����庁@^<�<1E��R���7_����9�r��]�����:�몜�.�a�u#Ld�	��$^Ȟ���4_�zb��iAc^]&&9�8�~����AG"����:EB�#Lʕ"�*����h�˘��B�H�A��;ҩ7���u��T;���ڈO��r���լw^`>��tz@�^hLKg�]��)[�B~�)��wM}�4�C���$���o��.ː���)��8���wf�L�͘<Ê�����S	}1�he�Z��]h��	�N���v�ڑ#��G��J���67�?5ӟ*��Y�uk1�6N���Ȅ��k�EڡKn� �)�^ұ��O���M�Ē��!r�0�����FR��̇%=��)�YD��ki�m�V�s����t���ʸ+W[K�syB��|��o2�ɜ���z<�����~1�c�Y|����M��2���ߟ�C`�n����4:�m,Ny�>�)"�� ����uS��k��X���Ъ�	rڨd����[i��^�g�MCo���:"��%�'C�$��&R6&�[6p�A[��6jc�zBp��u�Z�^O�{��(���Yz����N=q[��\���O|�Z����g�E�)}bo��*���T.�]�C*	N0,�[����N'�X�P����)�1�<GXʪ|�a�}a�w��?�)�̺2|��MQ�I.���2�n���WI���6$�.�a��]�p�OBpL}���D8l?dh��g�Z�u�%�J�V��cu�w��R�ej�KS��|�?5���[�DH�	�߀�wח���Y���kx�<w(`�"�>c�~d_��]XJE1�Q���r;�!s�+�\P�����1��#�G"	���	? �4A8GPy[�*R~1	��sȣEF�3_0v<�]�n1��gm�9��>u�	�`@G�>�-�1���:y���˜�O�(�=6_��7i�&�T�ObX_l���S�x�w����tz̘j�5MI��򔆩Ql(Oa��jN� M3�%[����1���S9�TkڇH�o�q٭��.� ]MՓnL��Ԭ�����U͝ǉ��n�g=����b�VZ�5����1�c�]�ߓ�o�>�q��������>�փ�x4��U��wڽ�5לԞ�%N܈����R��mq 8�Z����|�O����������q��:�|��p̱8~U�b84�UW�:4VtC6{T4�F�k����\���hd��7�D��D�=��,mw���}�v�1ZdVө-^m����U���x�~���}崽�=��<6Չ;�a���u�{�!�h�	�|���k��H��X�tx1�Y�^�\ź�ǟ<�`��y�&&L�������P���X5������Lq��6�k��8�L(q���@�9�<1" ��~���>O����~H��l�ynŀ�J���8�	�z�9�#o�z���0���]���[������	��2&��J|�9gz�)uД]E(�����#�2�Cs"�$�(�k�d�-�cц�"X�zʥ�""	yʕu9�~�á��~�6�N4{�ݮ�w��Lh��g��q>1P�_���A@����7��&	߲Թ�Ʋ�;�g#bƲ�<��RVs�JJ���%��S9@��o"���u�;<��B�,}���
�e��d�W�4�l���b-�W9k���u���ӷ�!��z��e��n=Sj�]J�����2�͡o*�h������&�])�3�\��+5YyUv�~��4�~�a�-^<�GV�3����P���yŵ�nN�����w�K�N+�F`�,����/Ljy�"�64��7s�DJu`�AP�%?�ܺf��g{r�����h�9��l�F4*	�8�p��]'�2�Q����^�5fҤۚ�$��c�Fg7�������{�/�%� I�n$������'�`�>��EoS���8���D�̵}U��vE}ז��G<x���@|���I��ݘ=�!��Z��yd�a�`�3'���S���I�BJ�mk
�����/�F1��Ӱ���#r�o�6�pңO�e��"Z9�ə�>L��O�er⤰W��jL��(��&k�{��~]7�WxA{|�����G�(����	X�<\���Z�T��%G0��:N��>SN��y�����P������� ߡ��|�H���CY�I�oH�J�UT_H�^eE��5�Q�(��O�;��4?�4�1�����-lm��o����Q�Uz(u�8�(��\�J�j*�s�eC��f��nalbՕ�N,4������4ZjQ+jYID{�l\,UN�+7�&/�Bf�TnһK��R�"���OJ5�6������U:�r�p�F�>q%5UÖ���-{�Gc�r"���aڝuk�&|�L�,�}�\Eds��5��N�0#�3�����aB*-�/+6�
��[�f����ȶ��8�/���� 1��������3t1��t���f8b��_'�Q�1�Q�a	��^Y[�E\��/O���J�!A^kss�#\�s�n%Ǆ�D\[�O���&=�{��7<�8�JR(�z~�ߤ�.:�
x��������\Gv�^9F�ڽu=��ձ@�>�P$S�Id�3��~"K^��ȬT)==$��)�]���mg�w�	Ě
��a����L�g�|CG�F6?���A2�{��z��]��5Ut�fxnf��z^;9�p�ªT.�7�^׶t�On�!�ۦE���	=�)�u+"q�gKl����/^Lֿs<1Kк)�x�I�j��,�~��5v�|ť��6��mosH�^�
N��ג2@����_�t�� *�G�����j��TG��H��+���QS%!�z�������پ����)�W�r<8�ʎh�PX�]&��Wė{ZI�n�����4��"�	V��/������g֖�p���O!��.�E(c��Ji���;[�-�yt��MU|�{�h�0v�0���h4���ymWmf���P�m�Ìŉ��Z�RN�GZ��b��K$�S0����{�|��ԧ4�C���23��zcO��@1�\C3�Uz���0T��i.�^��;���n�l!^���p)m{(D�ý�����6���"7k�o(X�0BvI��/n7�����s�'$;����P�l�&G�!�$��Q���Eߪ�e�P�'���y��)��׸�1�s��zk���~�g�ӟ/��{�'[
���`�ܡP�)O� ��3x��]���=^	�I�~�5Z���v�hj���Ơ�U�nO;s���=L�9��ށ7��:%�[�[�T�.��D��'��Tθ@��ǋ�"tǡW��p�`eO��e:�)|3�0�nA���������-c���4=��i���+��~��i���?ǽJ���y��Ә�W�������,F��!�C6�}o\@~}�7���{�$�H��רE쮌�u�O��"C���p�"��Ռ	���Fی�s2L!���V�M�p8ܻd�MAdIz�]:��ս4��zfmA@�,8E�6>��a�l������vқN�����Xc���6�:&�&a7�T�M,ݷ���}�o��ɔt�,)�^G�yZ��|�����V�ܲ�MP�əOH�U��r�v7Th���p�I���mYy�Q&GMo*�y���o����|c�1�{e��\r�_Cݫ��E12<UǼ�yyU�R�O{#m����[��A�]�OU�v7YW��0XEt�<b�:"K��R)�$i5������Q�.�DSԉ	�0�2��w���}����~�R.%���wҥF!1�̽Bҙ���9}�����Xo�9�\Ժ�獋a�9�hLpm��-u�]���~/I��l��*����g9|�[����_�X��<A�I�1�`A��[4q<��w��st��~����$s�I���㸂����B�!��y����4몪zѓԁ�� ;v�+��>O4@gBۗ�v�Kٞ�F�L�T)�,���g�#6ބ�����Y���F��1+����q۱)yd5���z>]��`�@/�K�X���{O��������JF� V�jG��nԖ�ۡݲ;*Z������N�of�]Hd3�,�	��g���E$��ԧ:���~>øeL��Z"���f�ӝL�w+����ݛܳ�5�:3ә`�8l@�����-v�%�x�b��/MJqs�v5HB�����YE9�'}StdY�9n��5wT�}K!�Ր�N�[�->��a�ʬ�:՗�[��!�<lc���Us;��K�pn��s�����0�*��શPJ�����G�5�C�-[-�Eb(n:4)8��!7
�⊦��r��H�/e=���2��:�ԙ���=y�օH��Xwt��ȸ����0p%����m�s)�q�[��ˇ.
▄7����z��,���j<�9���AVd�ha�I)e�9�Fj!#$Q�7�D���gU�ɋŎ*�[�Oo6���{s$�T�d��YY�o��A���Wں����%#�>s�c�!�c�7{\)˭Qj&�ec�؝��U�=iXW�*U��-:��e��3q�#p�v�u)we[P�C�\ާ�,�<��EK���0�!�b�*����M-�v�&΋�c%:!d��T���}�*��u��e������i�J��d���]w8�G��>�����s)�ߟL�ei��e�;7�ʱS&�n�GZT5۫��������a)D`"7Y�nQn�ote�3.^�i�U)c��	��!R�l�����C�No�U�WM@��j�i�w"lH���j��Y,+�����Gf�Iln�9��f�Cl4Xŧ^^���GN����-��Î�s;F��DD-p��gٝ6ܲ]5�{jr�6R�F�E�9cx�]���ȡ�z�/c$ڪ�%���M�ȑ@�dW "���OaYy	u^{��Z��|��aۘ���j<��.J�6i��/CGn��`��SH�5��f�!�e���R��h�+z2��5V��y�ە�q��]���%�ɌzZ�I��Lmb6���SY��m�ζ6"V�
�*'.�2��(ت�Nfb��,�����/f�%=�*��zkvG+��3�}�:v���.z��h|:�1�lqX�]:k��)���p��8���b��|u��Iwl�u������A�,����6*eFu���{1[����dbfb[��L�8��u�_n�k^��Sڣfr�L���g����W7�^�uM:���2����'Nd�K*�Wq��%e�����X!����ҽ��:��pJ�k4��8�QX0`L4�0�!�Ӧ�,z�*t�q�c���l�N|i��Nk��7��0	���'f�,fj��E�Z�光V�Mn��۵�ݷ�3�����Tr�:Mg�y�v�nTt�V��;U]�ukru�����ڕpА�9*��t�XFCͫnfP[��㼛M,�H�4��{��k�{��Ͷ��iθWJ�ڷ5�b6�,R�Pᑎ�r�n�c���o(mq�އ;��$9����K;ܒ�)���䅖��yS�B��3_?����E5�N�"��;mݗ6��ˎ���.˪%E%4ۦ�\q�Ǐ��<x��?/�fK�ۻ.m��d��+f:��Μ�8��F��q�q�Ǐ^<x��י!��YՆڈ�8�������3Q���GYw���EU$�1�N�q�x�㷯<x����VXY�QFւ��+� �kmfn�m��cIZ��4�$��O[m�q�Ǐ�x����{THQEH�$��vegvu�㴩�qY�Ft�p���Y�*]�y�݆a�S�nγ������kw6"�#B����,�c�m�i��e�uifڋ�����:���#(�:˦l�h�l�g��eْu���;���#����e�w�a��n̲��㣳m�b����mg��l5���e�P �����r#lDRh�Le3�$� �mBD!�d~iD��B��"$����%�U������[�5���oQ-P8�X�r�LނҊM{��b�#*�pK��nfgm�BK��0�����nz��,�e D��15���A�����D�B#d�
2�j@���*p��!��zA8��)�<�(�+�(YfF�m6c7.EJ�H��c�ed���{�.���be[r�q���ۗ�AT����gu�lf[:5�����B.�K�ƺ�%��=�����0CG1�y�l��qɁ�v�~sbFt+K.�̮~��+}�̲4�NZ�t[���G��v�������rힸ���KY��q=g{�}Cs�J�¸U½V�zY��h%%�._�V�q9����{�%!6^,T������I�&�WkI��ȹ����j֡���u���pFC�G����mk8�}\�׳9i���4D/-[�d�qu=�Q#nݜ6Z�d�Z��~��˺�<%@�������ո��^�[�.|��9��G�[y�)[�������5�m^��~�������95�O�۾����W�g2�R��t�D�FN�6Φ*%��})<lKNETD�x�\�ǟ�*�^{����7
��\ซ��-��I����q��4�ʈ|���7|�)r��2���n6@mn��y�K�N�3�.E@�r�!ַ�ZQK�#�����(���xۓ
�X��so��Zy�$㹯�9�&�[$�h$E}�}>Uv��;S���73n��Cw��)"���j��p?�.��3�[��kz�q�Ws�LJ�m�/I��>������������ݴg$X��֥^�ޘ]צsyr���MzV�Ζ�;�׍������u,�0CA5��	��1y�,�n�ue{�GR�~qT2����ً���U��\�z��6�W��<��{�S�@����I�k�P$�"�=˭�NFʭ�m��Ț��G6�e��Y��q)4'�r8h-�d��wb�y���4�����ny�l���ćd���6`��O�<f�ZE���'p��b�>�ɩ���t���#Bp*��f"I#A%���|�w�LC�$�j������@�E���P�	�Da��R�ٌ2/7�M��d������P�q�u�7��j��ǧs��$W�D���y�.��x��c��[籪ݧ+P�������2���i�L�?�c|~gs]iM��{��f��Tk���Ci�/*���԰}�W�h�k6�������73Օ�%f�,k���Jɭ�{��-��阅a�r&�+0૕u|8�fYSTp�QaJ9��Sz� =�o�V������7������*Ѯ�S�LF�5*M��z���M��DdG`���Ln���eb&ݥ��ӓYqIxu_`��b���h��x���||}�右��[���z.7� �T�T����Q�S(=��	�gܻ����PHi�����s�X�J5IFю�*�Rd����k�\-��ԝN�j����XsX�3��N���o�ʼ�3k��U�7I�kw��l���C���.m)��5Ϛ�_B�M���񇹽\�2��b��V൘8Nmh��w�Z�Y-bw�ۺF�wJ}�{H���O5��mr{��}W��%�Fb�mp[�X�b���p/ɑU~��D�ޟ5���4e�5q�}����߻��EmG�f�)_����"��j�f�F���꼕��Rw2���JAX"�n�e��؅A8��q<=��,��'�[��1݊��U�C�o��.���;M�+�ş���~\-�z�g��"�ym�n�l��9վ��X�h��3ŀ'��A���<9��P!I��Bib�F��wc�قEAE��x�&�^u�Z҄$��	��md蘁�WC��u��B�n����.�"�T�<qA~v;[X��T�k
��Zlm�Y�w�e6�ni51gr�f5�1J�p8�yX6�oQ�v�7�15NH$�������ʾ�_WO��)��P�<�����J�Uɯ\��P�=! ���඼��glR�%���ܥ졳oYa>���k���O�˨�nlS��i3�.q������~{��W;~(xXF^neY*����#�،W;�֪�]/f�@J��;h�$Y�\Eȗ�q��u�ɝEz*�����l��.�R0R���ʹ|�#��۲��ȴݪ	I�;�2��9�;��Յ
�7�EO��OޖK�<�	T�c;� j�щC^���O�Д��c�d��S�M����뎴g�����Wt�Ѿ�#A�zV�-U�!��m��o<�.��>���U�F�?P���匔�ڡ���>֠�W��#����~�#N�y�w2jMn�ǲ�Aך@:�c�;��~�r5cG����c���w���&f'�U���W�	b�r:�r\�s��3xZ��*�l�V�9ۊ���s��R�rG�FG��{%	��MɊe�_,�7��d�8wA��K���/I��=���p�o[��p�ML+��Wh]<
��NYS����Bc�c��/����y�;��7t�}��g�~hs�O�!�Xn�+�C33vӘ����R>�x�H
�6[<Eǵ9i��A���f�j�K��w=�']�J���$7�k���˕!�ێ�au���|�ƾR��y�q�H��NI������-^�&a��+lv���ѷ����%�΄��`�gU�],����}}_0]� �����`�F���r��"�4�f"g=��"@�0�}����2,=1�B){���;��h)>�>�E��ﰦ��ܿ�u�փz��
 Cݣ-�n��<�*��H[�W�����޲
�VD��W&}�吨,�
�2`�3qW�w<��X\䧽:/%�e���=�x����÷�ӄw��.]�:����4�ݧ:^D�8�O�p_�ٖhȝҋ��Yt2��{UA2k�uUKZ0��*���p�{f(� �y�������+"Ĭ�s���	B`�IꝣGM�*�F}�V[$L1��W"�#�<���]r�ݗ\R�EX�*5�����r��Z���F�?J����<��Ǖ�V5|�\| �ڃV�a:�YTo�1�c^�X�6`����ͷ�nu��"�^n���.�ͻ�*�w�mL(���5�~1�c���3�{���y���W����~��4
�bK�b�EqNܬ�E����j��	�L�4�8��8�_?zG{ ���fO�ЇI��`����C�v�ve�f�|x����L��[��ƴ��~mM�8��A��1�}޹B3��)��Z}��7F���ŭ砪���f�s�~)n�<�Vz^=��ȽfV!���K\v�+ :YϾ���&NuU�ʼ��MzV����>�*��Xj&�8��c^�_�hE{l0�O�_U�)LJ@r����J�bb!�%/�QK;�������;��%�'��\8��P��K��ذ0�U����_�W^ޑ�:{�>|FKPs�6�a�QC�z�/�ΙC�ͶKCj��%S_��#��]~���c�Y�d�
�.�)K���]]3�w��oJBh����|��	$O� ��\��R�?��^ �c9�Q�zPף�s�ջ-���Pdw30�Ё�����+RA�&�S�5��>�; ;��?'x �uRz
�UuÜ��2�
��Ѧ�a{nL�IT��P8�%{\Ժ�w2��]��K��3,ի��T�TK�b���s�KgS��������γ+����j"E.��0�	���X7>ݟ:ы���j�]E@9�y�<|s�^=E���|au����ѷ�\n�P��^�3���kw86�Jܚv��kĺ���uf�0��K&��M������>GJ������G=�[y�ev#���b��+g���M9��p��Y6���,��<�&tgc&�}n� ̈ ����a:=����;U���},�Y�=`(ܯK3�R�v�Q�g'\�����Y��p�=<x���Z��瀪p\�7]�&q="��o��˩8K�u������B�m�*��������y�wK������mh��*ߡ��)ߗ���Q�{1J1�-�����xS��n�6Y��z��*�OH��UQ{��"��T'�n6��Ov��B��#AgY��_8[��6`{6����|y{iΡ3�:�$��6�-U;�ʐ�TU=�n4�鎺�bw�;'Z��4�4u�\���:"V:���k͕�����|b�
>��u|�g7�u2��뚮ae��s��5Y�����W$u�1OL�t�&�;ׄJ��]�P~�x����||v+9xL������^]jI��=Qg�̛�J��s�����|��S��>�c�H����~�|���o�.���m@ߣ��}?,�A�׵��9��BR2q��U޹�T&xM�X���l����v�o��41����ж0�?;���<)��o����Y�IT��f�2�}�O82���(�1J{���S2K��QP�1�Q��G�|ITUɫoMOD���7��Ƶ�U��P�q��}�)ǜ��cf|�Nz~�s�r��~5�w�����L��_�H�(�f��.�l4�7l��A���BT'MW�;^��>@@�B��)
㧎�=y7^�s4T攉�����UF�R�q���}\h�7c�=ߍ$�B�&&�j�X��3S����g�Wo���;���g2Dj�\�����{=��R_�'�!�;U��j9��ؽ]PX�U�Զ�i[x�-�MQ�0���'z�A�OdŴuY�:����v�p�y�[hKu]\����s���oRZ�i����6{�OkP'eV�K3��p�ZΖjV�F��Iq�fk�J��������c�';����K9Œ�,6�N.�
 Q��#�`��pT'5H��ބ�θ�U%��mY����=��6��[��<�-�L,���Q{Qy^�C����|�-��ݵ���*{������a��V�__��<(�d�7ֵ鶍>��yݯ��#	wpՍ�����b�H`�ͯ�\H��eI�6f"j�j��uW.� �Z_��>T�t� iB���S������s&>6s�wa��X,�z�-/7tf|�Ѻn��f��&��9#i����їt<Y�Vm_0c�&��"~��AQ�x'=dxQ��Ki�=�k�va[�msO7�;*�)�&�{��q$t�ϡ_?�z4��g��:�7,��XFcj�L��ǥ��}��z�SD��2�݊��δt⻫�7xϒ�&9�e,��s#_��@B�[���z'֌3ҘF���w�]�M�y̋ȶO��Z��Ø��шO&��Y��6��qέ,��Ҕ�(���$Y |}�Z���.Z���.�ռ��˒�(z�	՝Qs�o��KK���TAv�U�Y�Yz������x�	�{��o7����n�����/&���ݾ	���p������l�5}-�x���5l���b6]ұ��/G�W;�<��lv���ay�D��Ucպ�I��`l���`۰雋J5}o��g"�^������j���Kw��զ���ɱ��R�r!(���VdW��(�m=7��N'qs wk;�&|�z�.T�[�́I(����%��x�!��p��]ٱ�樼��o"��ɐ�#'o�T�ُ��"=h�F|��d��I�^L�v�v�bq��j�+L ��j3��d�����N�QG:?GF�4٬c��+�Ɠ��#WǜԮIp>K)
j����Ľ���Gl�}�Q��\��!=�o������$J�gV�TB�g9�`&�@����=B;�2��G�^4>dL'�	aTκ����;X�0s2ʫn��qL�f�_S;\�t_U�je.9$��-M�f�ܩa�.)#JJ8n���}�4�IsY5j�=\[���a���e��H��E]�Z�bN��6C{7dmB��b���V%"�y+��I��T���H����V@ܷt�X7[3�<�� ��Hqx.��֦/���F@��o3���KRZ3SV
!���,����\)���Vp&n��������#}�T!c��o�h�Pګ[{��nPJ<�P��yw�w�9���Yo҆�<�s�����i"chd^ʚ8M]��c��м�cd�.31yF��{V���1�»*�yep�uXw�r�NV�uV�MÝ�]�,w.�[%89G�w$�T����ѻzo0�Q���ٶ�ZŌνٴ�Y�On)K����m.�wLf��='��o9Y����b<�I�8w4��d����}�z�ĉVvf�J8�en���L(�qZ��5*Ũm3(�ݢ�qY#����Ɉ釕r���Χxm�۷b��TB�;6d��'J��g+F�z�IC,�Z�,�z6 Z��K��T$#D�Wwx)�u���]�z��7r�Oo^U���;�i�v�hA�G*Y׆�*��2�[�-�-VTe阆���9�t�7�U0���������.���2��'���Aks�]e5&�[6��F���v�
�v��U&����	-��|9T�Ӌ~I��Y4kB-�k`f�K��B�U!A(43TK���s��}�3-|���K�%˻�v����E�����(�&bco�0��w�UΈ��yL3)Y�}lf��u-s��R������ܦ���kMV�(FV�ٸh���B�����.�إӆ?w�`Δt�����0j��X�fn*�vom)2���0j���(7�jX]��qL�7Ԉ73aYp� �f�LI�h\dx��<i����EuX�F�3���uU],��8�熽u�%Su��w���w��:e�VPt��4NY��{z�i�����!δl�^����#8ӈ&٬fޙ�H</v�.��Z۹��>K�(�(ORZh�P�y���M�<��N=B��b�roW3�qfr[w۵{�l^�I�G�:��	�n���A����r�U��tL[�Dd�
n6���Ο��^�e!wQ�7X���&��Ԯ�6tV.�'M�$z�wJ���P���A�
��'ЍN��w4�P�K1���5�\�=:^��a�/��av�P���p��^ T{�{%I.lj"����w%݊ai�kAY{I�#{f��j�+��[�RRv:wM̬"�:�4VM����n:��T�dy�(����YwX�lg�h�%�cd�"̛YΚ�L�c�M�[O4��ff8��������W4r��Ǹ��G�"Q�>D�!�\U�f���m�tڳ:�D*IRFB@��Liۍ���<x�Ǐ<z�t$�d�B@�!�[X��n�3��ˎG-�HIF@�i���q�<x��ǝ���~w��N�6�H$����̛dD��[��r]�B�Li���q�<x��Ǐ={��Y���cQwfwb\rP�Y���s�ߝ��;����Ǐ�x���;(*FD�E5+�����meͫ;�yn8���s�nӲ��m]gvu�yy����G�6���YVYGi&i�Y�5��J2(K���):NJ6�A���Q-���.ʓ2R��/��^q�$T�ʌ��@�k;¬����;����̏�w��Im�w�ОV�ߞ�����j�68���f�p$Z�[Đ	l�:+�T����y[[�T2���f��E�8R��u�
�^x���g��]���2��f��SO�|�o7���Ù]�Tq��f&�7a�I�k=Q���#�Pr/���U�~NJ�#�f�'�U=��|׳u�.w���`����:$�:�:�{�>3��8�ͺ]���؟�N��}�;��E�F߼k��y0�B9^�l���FĻ:�s����Ut������rlT{�\�՗
�m~���S.w� G���)���"�,:�P����eZ؝D#Z5�I�.�|��%��Q}�����^��o�₿d�*�NP��3T�y���FT_b7^��oU5
\����^J��Y�w��0����ۯ%��=*q�Φ����������)G^�r*i̊� md]�%�9��aSD�ݾsp��&5�΄�g�)(	m��:�D�<��tb�8�rݞl�ޭ��BuEﳄ�9{�g){�s�A�����r|i�����7aQ:\�nlF�J.u��G��81Ղ��R�vz���a���M�n��zvB�r���\%Z�Rb���Ȱj���OHv
E��T�&�:Y4b�`�yº�mo@Ӯ���e>7LWq�}"ʷ�n^������t��������`ר='��C��ZZ=�<�r�J ��J��gX���QW�צ�<��w�>H�n&5l�}Erh�:�KT�I���Vs�zg�zK��ȩv��Q���`����R#�gۈ߮����|o^w�+�+�={;�>*�>G��vC1��3��y�����-�U�P�7�^׍D�w���U᤭� ��D�XT�f�)l�0r%�3t3�J}痧���{��hrp<%\WOK���� e�o��}��؅@��ɉN=���N���ͨ�a��}[��W���Zk�+����ƄAy���Xt��،������>ƨ��X{�[= n��X�4ᤓ{n�C�;=�+�r��� ���}Ra(�	����*��Snc�]�͛YͽO�ie���])ا��K?��`f}H��v
t��Z�C�>���;MSߙ6��4��2��d�RgV���O5�v��R9H��Z��N����_�R<GdPw�oQ��XS�jwf��7�S�v�f�g�b���^-4����N��lF���#{���D&q��;`�����������-.��c�]�.�Ժ$M�f�ڝ>r4*T"��D��j�oh&ѠWj֧�~��>��qak*��>d\��`}N:T!`�υ?�����q��qW�^O�i�к������u\�<y�+]�7zxȄdA1�ΏU���Z\RP�w��3�l2�5i�&)��,8���/hig5�\��F+3�$Y����8�IS{֠����F�e�����gv�!� �\D�x�&�f(�=`���ީC��KF8rkwx���j�u�7^�� ���6��e�^&4�Ff�l���s� �O�}׽����=k['ݲ�����^��":��u��2i>v���5�:��(��Y����<�U>�xϮ�=)�r�&�Yܙ�h��~�>�<�6�7����Kt�x҅U>�m�����Z*���X�����#ހ��R����K�kڃ��yS�UKK�UeXE~-�@�.�#.�dY��Nn7�^R[�Z�c^��q26�ݻF���U�������	N4�Cjħ��7�/K8�opp�5����\����sPr��6�X�ot�U��,�㺛�9���R�b&��2V���1�kY﻾��ww�~>�N����?b.`�qZ���$���B;��g2� s�E����S��PC�& z�J꣧�+���ں(8�,d��(��a���-�}şhA�u�ݾ�g@�`��O�[�W����hٛ�����Utcu$�a�<�w��g����O4��H��q��e���b�W55Zޏ#�6��VFx
��7�����꣹�������y7��bbA���nߤ�/���C��x+��[��C����N��[�U�ܪ�&ܯK��]>�{��c!��\´o/A����r��g�`D6���ط�}�nuUג:i�=OD���]�]p����=��T����_{�9�8��9�T=v��V�2E�J��!v����-����s��U<a�=����L������NgوON˝����U[Z�@g�'�]I�5��ET��F�nVi�������2���% W;5��Su�ܼ�e�NUf���5!�:��'QX�;��\�]Pb����綧Z��L��k���mk�O|;������{���0���y�&8z�8��������y�Oٽͣ��br.-GH�M[t�oo6�>�Ͳ{}]A��%��ϙ�u���dǮ���z�9�4,���)wv�6.}w������n�d'�A���{�<.z ��[ˑ:}ʘ�Ʈw=Q�3_촇b�,��`Fm0_{����ͣ�����'����i8�����T�� Y|9��=��yZ��oV����_��#��۩+����c=����j>x#���p�{��C�H�"$�<�6\�ɍ���+t�2��y�=����<�oI�ưx��Zm��W��9�&���F��(MtN�/�;���)Mi<�w��L�K]�)�Ԫ߮3K��2���(�g69X�K=SMj�'�4���o|�&!ݪ��k����'�a2�,:��埝��3�J��MC�ĬF�t���W�\kIo������$2���+r�>!��{�VE���
�y?�9y/�A5	ܮI՗t^C2���p�O(����;�O���t
�v��3�m�Ϸ��U�//��>�z)OS���ʫ��74�\3߼|||||@4)����m ��{C;lӵ�s�)�,�S�F�>
�z��u�mv�7M;ƫ1R.�^.K%d�\�ә�[8@ߍi�Fb�D��J�O�(�x�[��(b��Ф�*�)W�����^z�c�[k�/ۻ�e�?Y��2���xا"�
���eb�IZ���I��$��T*�hԥ���]��*O��؁{)�����3g���z}nP�0�f�L�vc���3�e6ͽ8���f�ɹ��ޢAs�Hk���?Eg�?8mꀎ���y��N�:%��������!����W@`��W��ʑ{���61�1:[���sI����.�{��lO ���S�H�j���v�?!p#��_qѩ�S�b^�Kk�K�oNfn}���#{�_Z7�q�4.�u��P�!�j����Q0�� �f;�Ͻ�Ѕ@����<+�mY!+��E��9���SU�}���S0](%�֙(���^�~�[j�s�1ռ����k2��	$ 	�|h�	6QS;3�i��2͗�o[&��w��v��&��v��6�R�V�T�����ˀ��a�˓;w�^F�^��������]�Ծ#���R)_)��˒Dfn���oZu�0�L<M��Wz�F1bbL����N�>2�9��s��ϒ/h�ۢc������HН�J��>ήQm�D�b2�G+�v³��=�p���b�xȕ�/�IE�rHl��6���%NElv��o�����^w��K��w���3���V�嬬�W�r�'ǹ���&��>x�*�R���~���L�ëXg���[�� ��	z�%�l���*���w��W����+;�zd�>r�}��5n;�WZPR�:C�}���o'��o�n.R��j��>�A`]����1Vk�~��$�IJQ�I��.��y�$�vU>�=A3#hk�tf��(��g�OL��Y�v���Of�a��F����uә��7�a~J��S�e����������
��-q�i�p2�`Sn��烞�&V�=�<�V���ދ�ƥ��W1�C�Ym���\�.ؽ�;���g)
ʃW���+KD��:Wҩ��X8�17���p(T�q��T�֋��)��/5U�d�N��jm��Z�И��;h,����j%U\"��ؗ����U�szگ��y��o7��ٗ�e��ߧ��4z�q�O ǽ��<������kp�N�T��t�E��Lp��	�$&WH��\c �Z��仧V1f����|v
�h��8S\�����a���z#T�^��~3�yR�0e���NO$j��l����Ͷ5���^ik����mǦ�M�w[�gv��6�3I�})s�Y�jgC������7�᱘3��0�v"�nQ��Gz�)�Z�Lct\ٮ�׸���#�tǺC�Kz��`�Ц��+��);VZ�񇀓f��mwf>����Tuz�B4Z�	�>7�a�/>�e��6@�SV���v8O�_��@=]�= ��ؕ۝��]�6��f4�����4d���E\Ϫ�����R�'�p��~"�3Ԗ����'�^��Ġ����a*�������[��_Z��č�U�Uک C���ˈ�N<�! ���3�g �ߖ8S�-��xb��S0����r]t���n�*V���t�!1��pH��!�̴l�=ܦV2�MZ��5r�^i|�3
=�֡�U��4g"�f�;��`��*�{��������w^�Kx�Mf�a�Q5�^/����uDϯc�5f��mNh��Ǟ��7�}\��y!���QI���O�9P�=\:� Q�f�+za{��v\�d���ՏT��3�v�n[�́Y��e,In�8f//-jg��4�X����i���)_<�K�����]=���em:�W�}>��Mq��2EULUA��%UPV;��f�^��b����>X C���jj�,�Tڒ@�}�u͝4�������]b�zz��|y��k�wS��!ڭ�ɚ�������TBPrq\�]��c	�����x;��&�&L��j.3�.L�S�{-^�������0*�Gb�Y���Ȣ�J%�d�-���|���5L������ו�x��8�	����=y{����.��ލ�n���ߺ���q��;�a&$9A��䂻зG�cj�x�ôpe0����%T.�ט�"u��H��՗q�+]�K��b�Uq��ĭ,���ݡb�Y�ܟ���#�;o����7Zw��ngc$��׵�\HV3���G��jޔ�;����C3LV'^	�Y��3Y~�z���1�c�������o$<��ͥ^��+) NxoI^��d��gU���riG�f��yz�^3Z����fW�=x��ڶ��%$^�UG\��ц����I[E�>�<�п0Fz[��5u�2��gbkK�sN����iDn���f���Y4F��M��c��1'���KH�=2�;�����������������b3�[(�p�T3�l<Guq��Z��M[3vD��k�I�v����S� ���U͹�U�����~^j*��D�� :���u��2$\�����]�w���$��t��JD�EIU~z����)�~9�	�ǎ�v[��<�����o�v���k��9����q�6�nF50��:�ִ���Ԗ�s#hǤ���ٍg����%u��)�T*l��{.��곝���g�4�۫̚�����|+Vྂޚ�|>�<4�u�c�̕J&��f�y�S���v���μ�T�I�V*'I_b����������B�-���kE��*6��U3���^�#YNآK�(�'�hc��t���Y��jZ'I��j0qU�ym��n��f��=���ҽ�vKWM���ٹs`�nH���T;�4�]Ϟ�=	��u���o6��6�\Ν�8�Wy_$2�er�drL�ٕ�-�E���,)�4��y�	��c͕�"D����8XgcD^{/k#�B->�*t��Y̝�����q���|�m��e�Ķ��ebw(�ѝ#эK���2Յ����l]R�}�\څkA7�r�̛��\�o]�
�:��SYP�.��n|��	R+�잼�v�Oq��h���IUJo�R1!�j�%s��s�O��K�c�&�>�Qj�T�B���u�{o�.�PUD�)�'�)Y�)oj�ƕK���^%t����a
f�gpbf���j��+i5Nn����<6qt�A*�Pѫ����3W���Ջ�sm�2ݱ2L6�&Fp�N)S+0�ԭծvi�7|`h�J#*[�`���R'Ơ��wb 1�z�9��%^��f3wNek4V�2�=.�R�V�#T7F�g*h�n�AM�^�vNŽ��j�Jb�]�hH2!r������k�eˬ
+��L¾�S�� M�%K,T��p9�:�-5�$���(��s�,��S#*E�@�%�(�5�urθ��3v��*_���a@����W6EC�e��"�k׷�7�
�egA:po�շ5�ğXd�푇h�;sGؖ�p�*�������{�(�2	S�l���w���)�gm=B·���P�^�#�
Vk��(<�\F��'{$ٹ�Yyyr��4&�neZ姙��j�&�m,Y��E�2�[��b�SS�ܗY�j�����vѮ��"���F>�U�&V��d�ݱD�w&*�U<G3�
���jn�b:�ɪѳ�bR�6��6��n6dh�u�*�Z�[��)l�N�c�I_�݃W(*n5"��T�T�w�hq+y{!UV:�*�v��}���x.Y,P�*S���u�\But���Wm��\�ȫ�򑦓՘���e�x*�q��gH��Y����ԝ��CϜ���F��Y�v�q�l��]�Ja��2�o7�_F��4N8����r�y$=�q*+�wr�wm<B�!����nT�Q�-�<v{�8���U��.\������o(a18��u)NT��yzF�p�X� X m��.i��3Nm�';�QCHct4��{��K���\W[�8wvwdVtf����dKV�]|k. �F�s�NI�&�{�㪯.#S�qpWAj�a]�Ak��ӊ-�㣺��ּ�jJ�j1�YS,�����P�H'�(���G%9�ݒ۶�Z@�Z�������}T�n���viێ>=z�۷n߳�o^��d�2w�����gV�[5��EBHI	��^�8�nݻz�ۏ\��J�*��F�f���u;5��ݩ�v��(��&��PF4����v�۷o]�z����DGH�~~{��^6�.��8	vjD�:z����v���n޽y��H�Sn�"����B�����2�.ś��u��"Gq��K���݉�^ZwgiF؄q�k�vDV[�KY�.$�:�ӣ�@����եm�hm6��i��P ��tF�V��J@G��-�8�m��%I�8E	�D$ �V��I;����ku�; ~~~��>�f�|��p����Y�A��a��- �-B��r(g�Q4CQ�1�մ���:�N���i����o4�9cA�����uA��RK}�T�Pi��D����)���7�k4FE �F�& )h&X" �%&�8�$6�2��ۊX�Qp�4b�BYJ�q���1���A!P� �I�Y.�)��R�p�jT�Ǭc�3[�����{��V�m��L��/^�FS1{����������+�겉���HF{[l5�����<̑r��x9��Y��0F�<zl�v���Ł�;n5�Y��5UwW��B���s�lþZ:#�n{
3Q^T�Uf�������J��K� ���#�	� D���lY��P�L,����gkOA�P!��w�bjw����r��g�=I��*o|jB˶��s���'|,t��|g���,��}���a
��GOH�Ly�a��l[����9CX��ԩk^����01��\��r���W@y����y%������8ޅ;��ۭp�����R�>=�t����(�2<5�랾�����t�_����c����O����=��U}Ǳ��?z�GӔoN����9}�s�!�Z��ƻ� �Uv$�,YAJ��㸨v3=,q�u;橔�@�s�M9�3YXd�-ܧ*.t�[�P�/��	�̷�1�Rx�3�)��N���%��|�aoFˆ��[7Fe��*�/�)V����u�F��#��E��#��\�7|��-b�\�x��4�ÂM��ض-��1�c����W7�﹪͟��~��f'˫��'�m��ެ�&�R��^T��#��n3�F�o0�뼣S/�?@�N��}���6�m�A���6�����Z�A"���������K����+�D�S��1���8���qyZZg�i-�=Ǘp]df=�A[��d�Į�	����GGs�����j�֮ģG\�2ص���+���w\�A��'�W|A�n�R"7f:6+\)�Z�X]�)�uZ�����"%��`�Ö���e�<y����0JB "����b��0v�ISKt���P�a7_C3L�H+����"�Ϙ81G�	�����)p!��Y��gT�-��8��ꗣ2;'$m��6�������7NP�Q�淝�D����Ws�˫��GWƢHq��ƍc�Ӟ�{��E
·�ZϦ.>Zy|H����C���fn���_�}Wf��;���k-�>�KE��4I�UC ���U��/W�ú����2EAWG�gK�ꤢo�4i��v�v�y�V�Ы%�y(i��(���x/߼|||||}Rm�Q߇9��⦹b�
V�X=]a����)��u��:���z�Ɣ%s�>����W��OW]��G��XD���E��(�p�[rv�����8&9�����U�J�sE�!*"|W����ދ�Aݾ�aen�ji�nk�F,yb���a��ܟ?e��$(	}X��oЧ�n@�b�r損ED��^OޟHY"��J9yI�a+�uI���q����E&�����4�&��`(7"yJ�١���)����z}>�c:\RR�W��HܷSْ,G�����W&���C��K�p�Y���җ4	q���U�y�k��I8�v;�=�ip<4�2:��W�y��uP�+�6�G�skLϞ����]��]���$Y��/}A�$gH�(�ȭF�_y6#�X�~_1���ՊIY�ஆR{u�s4�޶wZݦ��`Z��NQ��h��s~yPʰ�K-whx�a�uD�5]CV���#��6ٸj�k�ˉ+���J5mc�x����yf쵤��n×�O/�^uP&p�Ju��7���Iv�':�[�J�K��w7�0�-'�Uw�W:z�%z+>�;����ǎ�s{�Y�҄���zt����ݒ6>#׵;~c���~.|��L�i�~N����>o=뿚�ܰ���8'�q���5#큸��ġ	�BW��P�ߟ�>y�s�ն�g���A��SD32���	���Ĩ
�@�p3���3��ot;�lg�C&�-~�����m�mS����{t1?��u�Z9^l?;44����+'���;�ЧK&��h�h~�M�<�,Ǟ�����u��/k��Y�fCȘ��������8u4�R��Oa�wD%vޓ�QY��t'hn���s.��h��y�.��F�:Q�6��r��Y�����Y�;�K{p�ܠ��6m�HU^�)PX�(��w��iä������d☛�n�U�Ӵߡ�Rt�%5uTh8�<�쪑�k�!򴪩�[��t�_P����3I��-�����^�=��� ^�� �n.�'D�V�Ɇ^�4�6�K%��4����-���n���҅U��YÏ�1�c����{��Dٵ�;�u�w����t�T�@�ɩ�QKV��t_4C���j�c�����GH΄�Ĕ�Kx���vI��ˇu2`������n�xj�=��6+�Zb�G������+����8ͨ6�e�7��`�e$�����lr�>��p�,#6_�s�:$9��Up'9ƯCM���.<�僞��iί�<��Z��� Š ��-kG)��q��x�i���&W/(����ÒV��G������TXv�Z��bx�Ւ\Qp;԰�����g�g[�6��;j��tq۱)8��#u�S�wP�+k�QJ���_��Lޡ���/J󛥎��p0_�Hq�P;X�J��O����'��wJ���_f��hm��Z�QY�v��ͅK�LAdFl�qD��Gi����{2h�}D���Qgs����d`���7f�#�Cd��/�N>,F;�&h�˺H���CID��;�cp�׽��s�P6�"�J�0������OVP�j1�!b�vP�lB�8�������\����xw��sE�ų�)0��J�I[��w��Fq';�,�ȕ-��7>��E�u�WWn`�~��y��o0x�w�Ɍ��
��&9���lI�dU�ЈgAܹwvk5�2�˘&)���t6pp�^ĩK�V�P庲{�ݜ9���AVK�n'C�j��1�;��6�\�I���EP�襋z�`fH��@�!I6�Gp����c������M�� �1��������wc0bo�XR�:G�+�E�\���ɭ+&i�{�mMV�,P*��7��H
��(�����Z�<�Y�iO�y�xs>�g��+���m�]k<�m�kPO��'��M��\���Q�~�v[���z�n�`�޵j�l����eK��ugsK�(
�E�5���x���g:�ق�ܥս�n�g =�"�bp�V.1\ir��@�J����p�A��u�>�����DuL���5�屾�)B=ح�УOv늌�ۉ���43�3��驔ج�Q���vir`]gҷS�<�uZ3T�d�������Ss-�3��|��6 ����sr�C�ț3��^طFe���R��Q7s�ܶbV�za���̖v�裳GH��}KS�y{X#����y��od�7Iۄ,����7,�~���\f#��cz�oB`�z�8�3T1��"0�a��k�/��e#-^�G���~�{�	�k��)r�.	��F(�q[��q������̯>5GV}�U���?�"��:�@\���˧蓎ո���3����VY��+�u�=:z�D}4C�#�}��Q!O"K/��U5q3Vʹ?x��>8K�?'�F�"ݬ�lv�M`��s��ju1��~
��y��i����]p#t�K<D��YjJ��/���]/œ��P�����_x7"�R�PJ<��<h��6/m����Y��uF�T8��>�vƏX��yꧪ,�t�S8�[��wK	[�fCE���r���M_ԧ�qp������g'5�;U��x�re�]^i�&I�S��6s��]���W����꼰����y��nf�j��U1f2m�6�3Z���-8�[7
�x$�LԞjNLW�-A�)�%Z���8�"�YZ;�s�O4ͷ6�J�)�A��"vy�+x-��]�7V��A��&�!��m�k2Kf��>����ɧ��1���7���Z�GYv����[��U��HrM0K6=�
�Y�%���t�ͽ��ƛ(.7ޱH:��\���X��B\w�ni��o6^DKG.�*��9uW7Ul߼;�8��k��N��y�c���+��c3;i5�e����6�4.l�l����ӡY���/�P[�'����(R�hTn�D�ݼt$�F]�#	e*ܯ>Kk�[{[���*�C�Nt�A�k�\�gv�y���Z`t�����;ظ�'���*p�.����N�bj��˺^��`#�8�PB����9�o`9�-GSV����׼���	r�z]N%��K��H��C�i��ܲH4�_�_��!����˞�hr����"��O�[�#�7�χtv�E���Z��Lױc����2�=�ga�S���E�Պ,]������N�7�IW�-U��&X"��!�S.݇���n�;�Ы�Xeb��nk�eUs[�k�w��O��N(��ڬ�����|�g�7�7������sku����Mr9����w>����z�fdWf٣�c�wh�p�hKρ�~���������l�d����E즄9�p��IV�	A����Z�z{CY��W�m���<z�-I\Zff�f��܇E�����d*�:����^W}�B��@ߚI�^Q��O�H��BMU�GA�����p�qʽ���42�:����o�k�Ҏ��'�2��8�7w+b�g�.�k���/7Eޟ�ˎL�3�!m\���0�e���Hé%�n��(����ߥ���R�b:�t%D�3*.d��댻�����e�0��ٺc~�����Ʉ�w��{��M���.���O&�qnrv�����A���N��v� ���UmF@Q\[*��kl�7��f�ev$;��:}%�g��b�)8+��!�n���Z(�Z���(���)�����'.����_F;���.����j	��P�� :w4��-)���4q<�3�Ӌ��`��O]�!��=~z-�M����so�U��<����I���2��z`i2dfq�6�:��}i��1�Lf�;s�)�R�]��+��{�+��1����֍C�d��ĩ7�u{�on��cv6E�H��qq��d��Toi���>>>>>>�3{�W>���aJ<�^ϣ<�\�@P3�����+�J��U�ws�'������V��B��|��s�vj遗~�4�Cn+��l�k�=�$ߥeZ��<��Wn���M����FC홀��Ub��������h�߯7�k������[�He}~��g�; v�Q�<.��Vшj���'gpghrg|:n�.ҧ���L�S��4B�"xN]U��������(Et�og��Ln��M'��^Z�9�����0��E�b��v�i%Q54bj�#}c>Z]:ک�԰U���F�:ٲ�&u���Ϲv�q�ߝ��g�e��zԇ̓�<���Oq
��

Uǀ���	�	oxFu�U8��yW����F5W���s��}_f�0���9U�'����'K���V���`�S8�c�캏�Ҽo��խx��W��i{�?����W7�Ox�d*���mw�s;�&Ԟ�j�&��\���Y�E���4n�i���7��a��d7KNȵ8qCKn�;�2V���K^����͖&B+,�&�ى����^v���n�D*�uAK���$&Ajt�riʩ颷�C��0q�����YF0i�������qI����sr���rQ���ힽH.</50�:J���C���RTpm�X�ļ���m�Cܖ�qf����/�s�I����v���-�,��10j���Ι�sY\�T���TB^}�os<eY�z;�ko74��]k�^6�-�č)5G�G�B�׳%�q���X�Y����B�r�j���U��B-��K��<%�ͭt�ɻ����8����U�U��U�J�3�(n�(;���Lʹjsyo{:�#�����q�H�\�M�[o��W$|��;<���'vA��5��/6�����:�����HcջuT�:��N��z�{s�t����AX�G/C��m�s���{�PfKeS�5�u�'6Y�WGKY��<ọt�3}���Ѳ]��ܱx,�o���]���2��*�RK���,gm�"��:��'�&��MC݉M
{��/+2�WE���/�gN\ �~	����~��2�����^�Ȇ@e�$��f^�֚?^���ʨ�)@�4�=���YP���
e:��ȳ�Kyr���O��+����ʗd�詶fk1��Z�-k�v֭�NHA�����r�oLZ���U32��l�w!{��T[�C:�R��*T�ִ�^�dp4+����x�-s݊śY9¯&�ݝyoʜ/�6M��+v��Y�-�E
Q]�Ǧ�'s�^Tӵt;�,\X̩�l�Wr���){�C����eCڭI9��nSk6���6��[9�}6��ls]�e,ȝ�,fN��H�LD�L��ҹR����b޴�s6�r-TF��Y݅X�ڹ"Eu�WuH�n�&m���S�z0��3fR�A]�pShZ�l٣�I$v�V�&p"�a�k.�!!&��۽�L^&�f*����j��z���1���+,iF�9��ݲ����
���Yx�ւ{��7�l��]�hAG��Z�՚�7I|��¸��t�Y�JA�YX���]��^[ޢ��.��@��ܫ2�p%���%d�d�".��r����/���Vu��iםW|��ϝMg�j,��TM�&]�i��SS����3��UX��bOS�ٽں��VPT�ؠ�g!9�mB��WԐ�H�jy ժ�ٶM��f�zX{_v�"�Z7qjL�yS+�{3�����}��o��a�BOI'��}+�c���R�N�.��9"$㴎Ͷ�Ӎ��}q۷nݻ~;z�Β@���ݻ񢒈��-�NE��佴������=}q۷nݻz���:H�C�Q
��AJN���,#$$$��J�ׯ^���۷nݽv�띒2B1�!Q��jUU298f���Ս�D�U!D%J�TI��z�����v�۷׮=s�$��HG���B0�G?5灶�j$'�Z6�ɭc0����@��է!!��A��,�w� �k�_N�T|������:�w�#��m�"�-'���m NBN���n8$���'!H�[��q(��� �5����˱�'N�'(�%9�	x�H=���׳�c���В�����)��ƳӚ���l�����9��VT&�F�i�s�'/m4E?E�c#	��1�c����r���T���ϧ��:��� J�IM�}t�F�,޺�4�-7�4������k��UV�w6����6���9���怅twȷ:�S��=$爄�B��b�ǧVw(�Ɨ �ֶۡv«�2����ף���G�~"�Vӥc�ك[��Y�Q�	w4 �s�V���f��0��!�|���<�d����<f#�ۭ���J]LԱg�r1OZ��WC��^?�X�ᛧ�
2#}�"̪j�N�G,����v�5_/!En}��?q�`,��>_G�yЖ}��2�ދ��5�Z�t���g>Y_���s��<������s2r�'���e�{]gO-&���Ğ�^+��!�zˮ��>}8�v��}�n�dmK>VP����]���u�ٸ���{�nrzp�I��Ŕ��vLW����}����;q�e1��K�Oy���V�d$t)�8ܙ؊��j�V������=��(۳��JJ�a�{4tA:���;J
�*�doY<)T괯��Y��gE�pX�V��w!�`F1���=�����w��~r������� >����BWɤ�>�O�β����|����X��!��xo����w�T9z���yf1��Tf��d���U�S�=��s�3�8� d�^TrZ{�ciڊ�s��U��w�|�#!��l�wp�X��^��j��FE#&��U^=y=4�4�դ.�^S=L���LVC���j�p�K�⒗$�;����a-����ocfm�9�H�K�>��8*��缄���%.h;�W���4|1J�w��%p�R��#��F}���|����j�X+y���i�Ū�ﰻԱ���u�g:��g����ͰԂegβK������82���,�|����<qN�a;�j���@i�<��䝀܀��� ��Hee�/9F��"��i<�;�ԭ�W�4�r+ؽ�áF➐���9�b�-��#a���6y(�����-*��a�S&�a�wB�Z�*b�e���<g:˩.9m�E���|O� ��#�A M$of�Cw��:�+/)�rbD9 �Vv����ǎg,p�wJ�n��[:��|�=Z0����UZ�V�r;�W+H~^>>>>>>>���du!�S���+�áo@�u�d�����BPW6�]bgզ���V�?�}-In�N���(�WB�m��gw���h[<º���vt&�<���mDK�Y����7;����c]��V�6�q�4g�����R&�>��Q�	�i�6n�a��8t�^�o\x%������x��2	Wo6��^���$���N����)Tm�P�`�>���o>^_���J`�HzJbjz�mB�3-�Nz+��	;#M�TU_ܭ��i��#�=q#a�X��K�*�3]˝%���:��뭡�?2����;u�Ϟ5䚉s�ʵ��4*�i��͸��Q��׻�
l_w�zX�(�F�B�4��U3XFn?�w�)U��(��#jȀ)f1`gBU�JY��y����a�n�!��WF�lzi���KPx�P�����}{����n�5�<�:�-:������A.s���BKf��UT�ϳO��h���S�y-�Y�u�_L��4j���:��G��VV٢?��w��3�ͪS�H�'5V�F�/T�W�YӗWp��1�y�~V^F��1�c�ys~�;S������OO*�k�]�g�Wc�P��~Ф�˼���~7���������sc��+EXc=>��#��X��jAKpXT���w+;��bsD�D{�~\`�Y��QZ�/�j�������D��m�M�D��܁Xsu�v��n��;�Lr���y���/�y����%�e2:�7��/�G v�0���LF'uA�;��䷽e%qsv�vQN�ˣ7;M�p+�E�Ѿ����|$x9��BA�k�/� �Y��
s6��篺6a�*�oX$!��A� ����4��[��-�{��5k�~Z��v�D�1?pl�xVL�v��u�ɤ0��1U}�r��W�;������3��'_ov[�ЬK�Y���>��ӳ�G�7=�b���<Nm����������j�Z���J��#|DO��x��f%Rt�Nv�ǎ�6:�.)TA��:�¡�(8�C�\�G�r�� �iWT�鯣e�71j�Ց�Ľ�|����8m=�/f)���4���ڈ��^���d]��}��qz�F`+P�f�r�Z�hUݔz�1����޷�{�p�P�z���`.��B����H�!H��֬�d:�233�����U�>p��X�c��-��\��3��+��4�
�=�Dm�5NG]�F��3{ix���ө~g+��=�=?���9T@�e4T�t��d�~�ܞ4
R�wzt��V� V{ �St���wL$$�f_O?d3E�<H�wx{���c�U�P%Q�����N�i@6�&��/Z��)�C��S���4�I_�������Ǩ�1��!�f�Or�3�F�L�G����eBu5gr��^�3��6��'B���in��<5<ڃ[�0��qf:6Ej�7˟��7�I��g<���w|=�d>�Yz������O�Uz'�[�^��M|��������)�5�^�ҝg`�{0�"~?��i���Pc���עT�-��`�2As_���f���n6�P�o;g[Ô,��,��56;,��u��ϳ*��V[5���*J��5��ۇOB�Ŀ+{]�]p/���k[��T�k"��2�8WYWb��U��]��_����V����1�c�gs2j������������r���u��W�o���fl�W�5�5�"�s5�ѡ���@]]s˳��O��z�!�dP��2��pQ��L۸g������o�m%���lvY���y��e�Ef��ٺʤ�/g��z>0i�-`x�>y�o��uѫ�}�p��PX��ވ�-��?2�t[��k
#�Q��Gb�dU8W�I�OdH����Z.���Ȉ��=��}��,	W��@��&^{,�R�w|~��u=v �Q;gX�{�x����(dK�Y�W M�;5�h�Ր�s�F�w?}jE�r_�9J�N�=W��&����J���GM	+5�~�(G�k�R�A��[����O^I)�j�-�!��3� Q0F-l'6H�Y�> �����
+H�V{�6
69��`s��iF��v��̴�>�Q�����
����TQE�ƚRʤP���Ծ6J̺�m�� ���C7/��qEoɦ��h�YDx3��[uE}�������L'��:�	4cJ�Y&���%��4��,&	��L�\�ܵ�A��fQ�_ L~1�c�xL�^xn�k�ATN]�t��FHu�J̅W"�7&aҮ$^س*$-�#.�(��˙T�F��8�i�b.������)�h�1�:���݌j8n�w�3��H����5��h�n�"���>��!��C��э
�6�g�ye��4� �t�%��C�����p�W_�Cf
�{}lZz�r[��R�[�	��x�U�ސ�{9�a�5y�׺k�=W�#�-�;
!�g�ץ"�?i�*�q�j����}�fh2��C�=��Ňx�	����.�W��{o>]f�+��������h�n�0�n��28��8���X�O�z����0?eK'��	���g-������x<*��U7kR�5ߜ��8�eȾȆm����(��I�1�v��"���t+�,�����6�/
��9n�x,�~�`uZ^�L4y��:�dҡ���ͧE�۟�J�(������1���h�{�a�j�wۮ�A��3iRڶ^ez���+q_P�,+b��/1j1�oM���7!�x�cEB��j�̜�I�Q�v\p���A�����Z��oiH;�k5pr��]�Sެ7N�)iŞ�������z��;�d�ն���U>�ng��v�.��;v˺�q�̲�P���O�+<$�����/cΣ�%��N�U^�)g�u���2#�Q���G63��P����ҭ�:�nC�V�Y�C�3�	޾�͔�Z��u�LE�i�g�ٻG"k�Ku�4��뼚�抓Ǻ�cuT�j�d���ǍC����|��ܽ���]B��S��3���Σ�/ݻ��ci�k}�O��sђ�d��ޙ�o=�Cbg��T!�I�pޛ� B����V�$���/;Ե_��[ϲ�on����E�ۜԛ���`���!���O���;:gys�^G�6�%�e�Dڮ3���j1��5�����_T���Q��z���?z���iqtT9܁虍|Uf������#��r3��� @��^e:�2V���D���q>q&_7������s]�t:��˂��uO�9e���5U��h�H��*���]#�����WS{�'��{U���oz�Ñ�b:���EH��)*غ�C�4x�#X�o%�QaݐoLm�cS��8��"t�w�p������(=�g���.I+�Y��\���T��s�d6f�o��C�3�ծ{�8+�K�l���%����ж3y��tu�z��|���vr;�Ԥ�9�����6w0;���Dю�b�մ�[��d�s�|n���s�ۚRu�0ݟ`ф`�2g�R9�5=��Ȑ{��]������V�^�[K,�%ϐ��F��<��H��B�xe�ҍ���4�t�m�̬�^yC�:wG2g谇��;����rY�~�2�L$rms�%z;�c�o t�N��W�M<9���ub#Yj�I���O#".�2]��h��^-!%)F�\�鷁4΅��7����E�1�b�g3�s0`�c��*�O�k^
�J�	J�}��u�\��4��YҺt�9&�#����%������h��@{s��w~���Ѣ ��H�E��&#�kX]e�)�v��w�W7u<p���1�A6vu]�fP���*��#[t���Ɍ�hS����O]������0�R�.Qz�P&��Q9GU���Dl2]�חe�&��Z�v���t���\_O�S�};1>�����gr�q���!��n�q�[*��{E�˫�8d|T~��K�3MuѲ+T֭s�_g.r��|�h%*�r��٘�!#�<��]��vq���+��/YoX�*`�7���J��;W�+����)��7ף3�ÿ+���w#�@w�}��YJ�����i������	��w�|+��˵>o0W.4t,���~Ws;�r�ȩ��u��)�q��+R;`��'��x��[8�;��]�X����I��H'�#��{�N�J��IIu��w�F��a�r�ƍ�؈V⠊������·��M�v}:�f��Ķ@�����^��q���ޑ7�ym����?�1_C�2"r�fG��E��븢�(�7�:���p����پ�Z*6s�{M]�?�����������t* *����/�?�J(��?���F��D�<���H��Q 1��FH�0�"0��F�HPb���H����R#�V�cHAb1�u.��u+�\\�������#��#1�Ԯ�\r��\q���q���r���rqs��Qκ�\��rq�s��q��1P�1�� �H�H�20��E2'����u%��p�cH �1�!H �1T��!#H�J�W.W*��.�uHĈABHQ"�U 1��R�#HT �1T�H�H 1��RH�)
  1	@�E��A��X�4E��`0F`1`1`0F`1F �E����Q���A}ף`6� �
�@b((�@b(�@`* ] �(�@`��@b��@b��@b�
�kZ҈(�@`( ��@�PD ��P ��P � �( @b��@b
�@b�(�@`)�h@�
@b!�$
�D$b!�� �H4�@`	�$�@b��$*��@`��hH$(��@b	�$�@b	���@4"A�`,�]t�U��8�]+�]!��(1��D!
����������U $@T�T�O������|������/�?������~�����{��Q���5������|�o��:( �������?�TE�E a �O��@���b��?�>�އ�E �����?ս$���6��P�a9`W��C��Q'��UF*�$b	�$��F(�D�$R ��@ �`	"V
 �D�`�"@`	 E"	H�Db!H"D`�HEb�H
F"
@`)`	" 	"	"D`�F(� ���`)�$`	�@"�"��A�$b	D��`"F*� �(�b� �H�H�$�) /�A���($��]]WE]�IWIWNutU�Uӥ]]WA 	
^��!(?�����T�@E$ �@P�����>��>���,���7�T U��j������>��p<���}O��G�������x~��E ~��O����� � ����
���A���QUk���Ђ��@)�_�(?������t��� ���}�G���h�@Y�!����"�
��m$�����w�?w�~!�~���"����
�
�7�����PW��C���
C��)zs�M����h?�����o�|Np"}�~��
��䑉��R󅁛���>�^�]_�
����(>�,TE������^?��!�'�PVI��Cbp�L�` ����������T�	WL(Q�D
)J���V4�eST*��	)SM�مJf�E-1P�AI$�5�5H���R�!-��b��R��+o]�(��i��αƋ+T[PkZ�ݻ�J�F��ն,�����d�e4�3V[V��Zɵ��6�I�Z���-�-��ٵ��m[d*�\u��l�fSj�Ƶ
�T�Z�m����5�k	l�l��fY���SiB��j���ݛm�fk-6Vڵfd���Z�`�l[j�e�����w:dGe�k�m�  �{��Z5K�h���m����kR\��n�������]���n��g[m�Whw=�v���wn��wN��wg:�����gks��^����j�����o.���e[5���Ȗ�d�&�Z��   ��P�5�f��S��w����S�mb��֔(�}��or���B���͚�x����j�7JZ�n�n��m�=�V���u[YL����p�Ǯ�{�m�w]���N�em=v�v�8���ήGl����m�5�Yj�4ٖ�|   ����Q�;��oO<����5�M���ǌ��P�m�����-�v^��Gv���;]$p��m��]���[۫���i\�uݵm������ۺ.�ݕ��=��+Ս��aJ�4��Y����  x��u�*�鞞�Uۂ��������Yolz
���;٣@�G���]�5�AР���ްW��V�5�RmfUV�t슪m��  w=��Y��K�U�<�O84 ���P@�*jj��ږ��A��u;�m�`j��wzg�t�j��ӊHO{�h��tp(Y�TƭfkZ��n���_Z���UWi�`ݭ�E'��2X��X�N�]Ul{9G@�k�^p�d��m�U�N�v�8D(y��M0�Lm�h��h�� ���`��zp ��p
������y�ם  ��  M�p�ڔ��p�0븡@����Ph�ڵj��l3Dֶ[��2�� .�}��������e�t0u�9 t�^�= zs��z=h�zp � ��^:(�g��h�+�:+@w�F��Sa�IF�3G��2�>  X� � Y,� V��P��@ n^ۅP=w��P�� � Mƀ ��h W\� P��Y�Vll�[�	��6�   ���h �8�t)x�� ��k�  ]ˮ��
=��8���=���Ӟ��  ޽�tz 
c�p ��O�LeR��@h�0�{FRR��  5O�<�UD��0���R�   Lh2��C� h Iꔊc*�  f�߿o��W�����9�9��9w���Y�K&*l�#���3��%=�߾�|>��l����=��km��UU��綵�m���Zֶ���kZ�-����������۹��ş�c��p�'cVe�y!R��E9l��'F�7��5eZ@ ����d��6��VXn�I�O\*�C[�n��R &�����8E�b��,)��f�1��"ҹ�U��9�t�Ւ�hc��KN	��G(�a�*��l�{�(¢�}z����־�2����K3 �y�.ݔ�!-��tN`Y,;n�##J���L ٩��"�8���7�M7A�C)��:.��T8"�7$/�^���y5�.���Ve,���gU6���('!�۪�/^*N��P�=��c>ŵ��j��YhE����Y��+���@T��	��S�ca�M�������-��A�Wa�ͪ�>���yyG@�m'�;̴��33p��,Uoi6�]FrP���;ld�ƒ&*N��A���sĲʬ{��)� �����{�2ћ>�q��Sn��뼄�ȕ�{�IA8eߛ<��X[�/q	��5���.��	��
V��ÛyKh-�[b!�m�̿��w�n)W�b��qI0fG����Z�A�XLm�@`�N"�� :�,�h�
�S^��Ǎ�wm�M,�(Q��]
ӳ�J��j��&�
�������Tx�6^=X�0wW�D1bw÷4��B�%�S����+�P襙Y��%��l�U��k�eXU/TWp���+e�yw7��9��t�V� �ͥ%Ão�@'���&�)S_Gu	TwE��\�d�bUՁOL%����1��K9W?�$�zj��N�\�;KK-R��R5���Z�Q9)O���\��D�An��3�ӑ�}���g����od�{X�XT�wl�l��\��q�cjلJ��R�XT�hz�T��oC�C�H!am^RB�v�G���×�K�ġ�2:�fV�I�8�J2�1���hi��x�M�z�` �R�����ͧQ]�#+�1M�eѫ�(5����X�[;�M^��LJ��C%��z�R�����pm�R���]��� ̳V�n3u�BE���
5"���M��*��˗�BM^�����*����-J����x�{7H�c � �T�
T�N��W{7LF�U�kġJV'��cm	��P킍<u*!P2��L��SYh�Y(�=0^��īk.�q8l��	h�6Dt��`*������U��P'UDXfH.�j3@���]=�-�8ȓF1BVR̢�3���Wm�8��[��sm����8��Wsђ"���e���[�u��t-^�Slzvac"�֘�h�+6�v%:w&�M̃[9�)�&�w�X�!�-[H�N��ul��G���84�҇Hf�U:�����0��"�j� ��n��xB�R�
�&�Luao�Q��@��R�sB[M�i��6�֗���	�:�����5�aF,�� �!��/�(R7VOs��]�N�1Y[�l;a�̄�m2�ĿG���8�{��F`�#9�`c�l���5�7�B��`�B��E,+%ȝ"c�����)�i�ˁC���u62K�Z
�3��Յ�I��V5Sl����	S"��iY�Ad#�yF�A�x�*��R��7+~��n<���X���l�H��ٸPx|I���y�9G����B�<0h���L���Җ���h�x:A��gvfr�}>��&g��:)��֛n�Q�dV^^�k�U);�J.]X�u��i����%�@cE �����:k�JZ��Ih�[-�
˅*��ĉ�m:�kT�&l�+���0M�M�k��B�n�ZyM,�{Z��ݢ����xC��:"Rfɦ�H��I��4\Of����i��z�"�с�<��o��8�����86���~�hM������C����i�1q�f<�!	&Y`Քu7����fJ#�]Kٛ��2�7VpR��(��laQ,�<&����'Qb��VY���/C4�Z&\:,i��	�{`�y�*dڀ
)��t���۳Y�3NbWiƚ�M[W�4��6�.�����0EB���{���m@ҫ��8KE]e�^�-�NƄ�ϭ@�bPI�A1Ǟ8����"q�Is�I���E��*3�:{�BqgOoF��)�ę������R"��%��Sp�#�%��pQF���wC׹ �(BrG�T!���ku[���&�^^�*<�@�90��"4���s3Bn��V������%���Yv�eB�f˳:��d�u�H�-�z������3��P�CYKMd���i�k�i�[�%�;�S�kU��R�M��+IW���w!�;u�/� ��}V)R��$-��w��+���VLV�2���r�\�F�p�'
m^Y��!z� �{���piݣxɊۻJ<.�([��WE|��`!pƩ'���-ݧ-ԫ�/i=Д��L[i�b�[��泪��g1�_3�f:qe�y��(��Z�F5y�qn�W��K-�䧙qޓn�Dmm��,7hMK{fee۔kn|@fa�X@Y0-��� ��:��dh,m&�����I$;���I �OA��S@�Ȧl����2�x
��*@
S>;����I���g3v�V��!�Um�m����k{F��cd71ؕ��\8�b�4�*�T�S,�@�m,ۭ9��A��/V��j���f"�}��.�&�H;�y��>��[L�� ��N�5&eF�Kl$Y�UmR��V��jֱ��^$.�B:6-	�q D�22�0Z��"O���F��	GXKA�Po(f�q�( �s7��͈ͦ�ԧ��>�4�Fm��IP�lxi�����b�1d�WRM�n�ׁS�7�T�R�.f#�������ґ���b��`-7ll��n���n�V;�]��f�(`xU��1eY.<�-�� `�v԰����JՌ��Z@r��&�-<�Ր���jʧ��gU�UEt����ܕzF R�6x����\�ɋqcf�g���L��V��ɯ.�rC4]F#Z��n�QY3fA�@��Y�a��:�=mLPMv��aҐ��AP�3ٛ�.������r�Zh��7E�e���tK��*�EdT��XI:GmӔ.��8Y�ڣZ��"D4�`��&��8d�J8���b�#[��k(ջh��VB��3�Z�t(��p!Yo)���A]��D��y3C*�8��3^�1��3wSv����A��b����x��
tl��L*�y�%֥��)-ڕ�>�q�7��֛�r�JJ�L&�,U�K6�� ���}���Wa5V�TCb����xPb����L]e�ɼ�7�!�-W��黅�2��fT�s^�Zm��pSrZ�� ���V�����#ـ�@M�P`��RA��1-L�"�
ЧY�xNU���+
��&�f��p�e"�"����3[ʔ�kqV�S��\�v[��gƱ�"��Pkxv�������`�����PN墡�Ѫkk_'Y��d(S�w�8��5��i��e� -��4\ �՚&U���7I,*Q�1*ٳ�ˣ��J�f(�Z@�O+n�,޳�v(�XP�1i2�d.�n�������nH�7ǟMΑ)���n�R±-!�vס�$v����RS_�%�E��t��+2�`��z�va�{�I��Tʼ-Gx^ћ�{���p\ �ۢ6��Y��$�<\,��y�PB'?&�8��Kb�V&�V��j��aAKʺ�h�LL��,�@��paD �tU�gF�e�wl@���7���
�u�fK�jJ��e[� ���4uj^P���+6%�^�W�$�i���'3�be-(TE\�{o&�`�:T�BeO��Of�Rj�e�Rb6�Ri�z�a�>�����u�a����� v<�f��iA��T7j�Z��]F(	)]H	W6���Z�O&T��A��Y�[��G*-��K��m�̹a����`�CT�Ö	
�$��e���F��yn��E��z���f�gv�Ad?��&�`-V�e���z�!�Ǭl�*�wNR˲�Dbܫ[7���nJ�4��
5�E!ïA�D�����P�j�"�U�i�m,Uvݪ2 �3h!�-�`��$q�"�ɥM��������$�۲�Z�/��E�B�Fv�>��^]��(�d�@ό��.X�FYܵ	�;mL��V���ފ�ON�7yV&��P��pM3	ӣ)+̻���FުPN�K��W@(2m��3B��!���P��b�]F�#����n�M�Rjb��S�J��	��Oa���"��۵vʟ!wAh2�yJ�S�&��t˭���O.�!kIO��RR��+����h4�&eP�6(�X(�
�kX��5�b�SZ�Cv��qk�����Kp������Қ����k�� YX��je]�KGEĜu�
�J���`���Ʒ�b�;�pݼ���&��,œtCm*G�u�,cuw�
¤�m�
�g��Q=w�L۱��1�f�����H�b�p�!�x�f�<��x�DdF=ZUI��H1Z��j���
���*�2-V����zt�E-�,��ot=*�J���A��Բ�miq�;���gmb1QI�{�.��n��B��J3��ñeXV�[k22�RV͕�m�RŒ�Z�@c�)ВF��:Ǎ�lG���@8m��lU��efA�_�1)��V*���̨�^�p��m��rf��\���,-I�1f�wNk��QԺ���j�Ú��-L�����Z~@*�u�RM�`I50ƛ4�5hdƆ�H2�')����j�B�F��350@����J���c�P��(���(m6`�pbӐ�s5��JV�Ä�J6u��'��:�V�v8F9���&̙�U�C]+k6�vs��J:�c�	����g7.k��O�IƶK�)��y�A@Q�:��v�I'r�t�TM�Z�IMY��]52���k[X�ၡ`��xp[vlh�tT!'Z�V�T�L�u� �lYV"ۚ>ej�+6��Ď6j1m�P���9�m���-�Vc�R�^p$f�<�}��@���_C�@���el�!ystC��*M����N�j��e�a�Sn9��D���Ҽ
�u�.�c��S�'�#'r�رQ���X�@;(8-��6j�v­֞�U-�i�fm���Y�^�d�k�v���+/Sܥ�A�w���.�䒚��:�c�%*/��5��*LJ�\�!e��n�r�&���Yx(��%j��˺6�<��j�ی�`Qa��W��ǆ�6L���1�d��a���u��l��HnV�0][�Nլ�W�Xc�#���F�%�ƪ4�N���l{Ȇ��j��H�E��F������*�i��ѓsj�$p�񹹦���M9J,L)�05��"t�.��x�z�����4K���N��\Bi^7�aV�s�(ۨ+w^�I5��"���bn��e�y���JT����챱���][�(IR�SSe��Nb����X���m�V:#؎�]��b������������zl���ҫ9�1�T.Xߥ'Qã�!�tbb��nVSlV먃td�fn�x�t9nQ��n̽ŧ2n���L7�<[���k����s#���W�(�)�b�Ksh�K�=���q�h+ŷ&�wa�2�Pt^e�WX�S��JX���;�TG��KmYFVՅ�N�Be�.��Pd��fC�� ]ZlS%2DM� ;���ʟ-�jo��Z�F:�Jn�@f�v���*�T�N؋-�#r�3�9�� ���Y�`;Q�z�^)�c�~Z�Â�yq��8JJ�ԥֵd]�n�;�� �p�?0��ei�e�f���ӱ[NeIW�fʶ�:���)�b,M�Cq5��/2��`���ѺB��H�r���,<$^�W�USo�j�F��U�}j�Qk)=�!��hCBܻ�j|L�i�"�����&eG��kY�ku�k�u�HuweM�#�R�[a;��w����@i�ʰ�gu��y@�ܬ�I�P@TF��7�֗��P*�]�x�,��jbp�ò&��p�@`�{Sy	�_�Eh���X�w�c��?M��`ǭۿ��J,H%m��i{ e����f�E���Aխ�q�^�h�q
���wtƭ��K�T �< ��e�⩅�d݄*{ ��u$� �Xv�8/u�1�v�i�Gme9����V�5旪���C'�k�0��wLR���J	OfOdC�@}�)��b��C����B�2k̲-h�(iN��+n�������%�f��/ꍬ�6�.���j�;B�ϖ$���e��R�It�M��;���e$���ȷME�fkL�^���eZ:�L��4�ĝ�cq�{%hZ�!ʼ��$�Q4���x3#66�ɕ҃cW����N�Wn��Ъ�������v�K ���0���_;���l*� �6�2R91ԥ�J�-�lc#U=:&��Ѭݍ���u.^��	��s4并]+	B�M��o�/K����t6�H�@���n^��(2U�zZ��W�|�6Z�i����2E(:��YV(K/��A�ee�6�
�l��h��譕��Ī5�wv��eS�nֵ֭1�.�jA[7!���."#E`z���v'�cN:I)��'�1�hĞEF�,��(Cr��)�м��P(�j��w��fP��.�(�چ�����Ea�%ک�V���jf�r�OZ^�)j-L��ua�nO�e*x��t�J,iV@���8�Cj W%��4���LU���wDE�%yHמ|F�L�1�ad2'��4s�����3׹V؎B�r��:%ؼ}9�j%�;�pr��D��Q��t⍉y��\��J�M[�Lv�����?��J�kv�wN�`�e@��ᖸ	��t�f�U�*��~s_ABˮ�qN�\��C�ZSح͘�xw����:㫕�Iҳ�u-�ˁ�*��E@�4��b���*��[��{xv�p辱7��,.�ȃ]��*�g3E��v�"��u���q�د(ʯ�}��.��
�Bi�uܹ��<Feu�����żM6'm�8���7���Z:��!���;��Єղ5��\��5���2���=َ��,��K�9B�IQ΋v�s�$�a�/��R����Գ�-�0hӦE�rgS�v�9"��3ӛ��[���b�]+���Z֠�MA���u0�r�Ė�E$��lU�C��V��b�o����n'�R]C��S3�j�.��%���S��ͭotEc���M��$8uv��c%V�ݢ�j���r�ӎD'a�ֽ�m�/M��)�=���gd��:�u2��v��vb�bS����U��g#����[Ae����8�ֽ�0�P�p�#��B��"Z�N9�@��9ᦇ<qF����p�:ҧ�FE$�VR��R�S�Y2�ཱ���9�<,Ѐ�k�m�oQá�W��׷�{r�o��=ss�=b�x�t9��r�%]2�=�i�ue��VP����jikN�[�|%��:�>ǖ�,��iN�.�*�7��u4�U��n�uK��:��7qM ��+�v���R�Mڸ�Kx���ź�nQ���`=��P;�m�����Ń|o�$���#����#��ck�/!;S�Gt!���m�����i�wZ�=��;8u��tnhUȜn�wn	��,l�j>ڕ�s�췚j�IQ�4�:t��+&��\�2wh��0rAhJ操e�s��a�k�F��H�n�TǽxOC���e�&�{-�����_B�i���wv����<����9��੉.�_�OKn�<9��n�=�+)c�q!��́HGk�6i�)ը�S�P8�a�9�=\C+��C[���{�۶���Y�F+��h�������Q&��5/g�v4e�?t���5�i���35u8̗զe�u������;�Z(�5��=x�p^��X=Zo�sS�w�#�9��OI�61\-q[O���,�"��Q�a{����Ӻx�F�!@�K�:�.���<���jw7Әɾ����]�-���(�\:�l}���:��T�N̝s5U�:�R!}���Ԃ�Ȼ8�b�N��%ueN�wZ�î	�r��:�)�Xn��6K�Y̓��h:��ZU��k�*�>X�fv-���{kZ��ۦm�-V�km�����Szl_X	�|ƭ'��ھ^��z{M��.I���A�K�]���5$��fE�:U�����ΛB)�]e�X���\*�Lq:�)^����[�k���Z�j�B0<�^�'��>��gw@Ō�QR�q���[�M���9�q���)�CCc�>��Kw�uGs^���w�oN*B���n�Q��3L�d�R�m���K��:!��-�s`v!ʦ�w��:��k�׆��h��m���ͻ�:�s�#;I7mP{�E����X|Y��}e�Չ��jV �lM�����Z[�st1s�����[��9���\Z���\��sb��UsE.���z�ݳ�em�V�t^ӹQ�RM�k���v^� m����v�TO7�Nw�=����?��W=���m`��tF��	Q���?K��)�篃�;[�Pۇ�tzQ(7c��{���?PC�Ni�3�=R��xq����#p��óe�7���_sxO{\�u=�ꦗ��Ӽ{l �v]��h�;Yl��P����}��Y��3��|��¹�!�z��J�0m &X^p:��[�drZ�0o����Q�:�,��յ8�+�5�VN3q�.�h��S��nסD��W9IrKM�\��\C�YN>	�ŊyI˚�eV�lBR�-�B�}�:��nuhm��y<9� ��n��	6n�޻���]8�����3�Q+4-<}ܪ����Ro�<�O|U�ӮYy���$8k9^T��u=����Ky��>ލ�Bޖq�8��+�SH4c�[H���Y����u\n���eF��˓�po�Ş� ��2���&9u�Ը�N�s�S�/m�g��y_!��@vg�'z��Y�Y�On!�Z���|����/Vy�-KF4�Q�5�CVg��n��L��c�6�$Go+�V �}ٓ{���l��txo���y謴:v�f�l'��uA�#;E^)[N�8�cM���:��W�����0���gzҝn��)�d���e��v5@��bW�NՂfLp�C5��Y
����W����5��+��Ǌ��"�}�x�g:{N�Ok�(��g\���%�M�A�n����6�[�3�P���s���� ��j;�Q�&H]@4Wu/�*<$'���'ͩ�xp{�W|6o�����j圸�]�zmt۫��H����`�q]���U���	m�dl�(���wҎ��TډlE�V���#��Yؗ��OTʂnL�i��ګ���V��l�����J�4c��G]�#��vm>���p�w(�d�T�Ȋ�vya��d��<�m^E{�;��:�̩@��f��|�20^[Y&m��3��E�w�W�f}<���HD��f���#7S7:0m=�1 m�HŜD���߭��a�EZ��A��J�.�O�k��P�e$z���b�u��6t�ǔ�]��S�Gd���j��*Č�]�\�kS�DO�ތ�Y�ݺ��J�8D�s�$6�L�]�;3{,���~cX@�u�L*���^B��n��0y�;ĩ����Yև�z7ԯ��CMW;�� �(��:�:j|4�[���1X�&=1��im���͹�>$���<��9^Fs��qX�uЦ����^�uݸ)E/�V~\�hY�m:8��]ޗl��m��m'b�kR�ll���e��&@O5d�(�_Mя#X"�ic�J�5��-9&�烜��π��j�ux_n�XFMF����7�k�!�����ml��Dzo����+5�	Z�n��V�	F�EIMS��xp�J�+Om��9����nSlh�xM�n�wSC����+5r��1Q���$����"`�dvƛOf����/w[^����=�s��a۽(���9G/SM=���y�HZ٢�n�2���
6f^��{��zLY}�c�����>Ї��L��mVnl38A���&�{��Җ���=]ؐ<[���]]�ea�9�jkhG���CH�ˁ8~��}�7�FV�VzN+k&�AV�b&�;�3�4�Q�fE:��C��l�x�m�f��.��b�bK<����x����GB����G;�_t�<��
���EDw9c^��ĴV�x���[��\��M*��1��&Uݴ�rv;�
V�Z��N<J�t������?�t�X@��������ID��n"�^u���(����2�@������qɛu�:,��9�o?7�a�@Ǣ��Gn�Be컹�����������bDq��[(������wa���w_M��3���S���a��6��(��3O7]oxRY�漙��h����ss�x��b�b����ی�S�[Wv|�Ÿ����1��j��Ab�S���Hݿ�t��uY�2��y ݙ�t(r�xf| �:�5��%c��ojl.�Ӿ��|�Y&p!ޢ�M������W���,�Ў�-乚�zJ�s:S��/��Rjȥ#�÷��r�*�@�{b�<�C��$�v��Od=�$�;V^�Vܺ9��g`��AMޏ4}�m�k�����oPo���N0�
�T���V�R���լן7���I�ݜ�'�fΤ����,���{B[+�G{�����:�艹Y/�W���Ņΰ��`�76|u�4+7�
�9���D������E�E���gQ	Tx��b��=�h�c��[@��^��ے�nG��*|0��� �P����;q�rl��wS��L���(.F�g�ؓ�ydT��B�-����y+LS���b���z�f�ȿd��3�z%B���ut�U�u���᪳b��sXT�+;�L�/W�0��br]��N��W��T茢����.�֤d{N�^��u7Zܳ��K�k�kj��ET����b^�k}��m�%q9Ǘێ.��B���y�*�k�����S�#J�ۜ���b��O����{�7��Q�y{��f�esO�#[��n	�q�z�s4��Z�Y���n�4�Zf�:�]/��]k�"��_en�����mnqq��3��4��k�n��!{��pZ�;U2ư6郊B��v�g %G&���8U�7��zs�H��
7y�:|mm�s��ܾ�:Z��P��"�!��R�J.�Vm��`Th��q��U!rVuEc3��W!m�������)S�x7��f���7q�թ�����L5�)�GD�����v�;�s��C�x�ڮMѪ��g���^�Il\6��zY�pI��;Vw��9x���厢X4]垈�b/��'`=8�`�YA��i��\ݭm��{�����]���p{���ֻ�#��	_-�7_gn�wn����g�j�_h�rG2%�s4��ć{�a��r�v�E�Q��*&jӎD�<��'<6�h��4�}��v�[�n�'�t��a�xÇ����c�N�����vi�/֧��#���9N6�R9��*���ǩ����hI�#�d������9w\�2����0�b�����}�#ȯ����,Oo#����,Eu��p�s���;a,o�3&u��� ��(���p��0@��=P�3D�|Z!G��<\��;j���"AgוΞ�r\mVdD���ͳ�����ӹ��'y{S��C5޳�R|yۍm��w���=����������rkD���
G�����2����h��ȟK��6↗��!ٸ(y�L�[�
U��7.C}G	�֩�-24�i�dt@�8�Xʴ��[�K��wkkyvH6�$,*�[��>�����K�+�i��^����<��<��9�`sn4[�_>���b�a��|P�M#�F���$<�_D��M���;�T���q�ſ����`�*�	{�pݛ�z�tnn��7�U mSOk���vvģ�O�{�A��%�����+�Qq�syW^Wvd�t����c�f�k� ò�ҥ�E���i:Yף�!�m��C����C+v��]5�����h#�u��� XFR�M*T�)�0;�u���p�Á�n�Zag3]�a����	����Z�x�3�yhWi�쮴'�m�,�9�h�;NkG�����6�ݧF�Xy�*�)�s�.9�g�鞬�$��f�v�[���˒zùfzz��۶o���������S���Uj���������ݩcٚRs�]R�H�귓Ҹ^��%[h����)�ZD{�*uHu1d���z���=�G�F�(�h�-���r�'��Ř�5��ൡ+�h����5����7�^�1u��[�<��S����7o����HXy׸���u����1�nA��XY����a|�MKC|�w6"B�F�]����>'��	��9ՇgU�����v:�;Kd�Rv��_c�Zյ���ޓ �O��i-�MN�u5c>0R��2�A�I��%C�F��ΑN�84�]�$�`�TW(��Sv<��K��Wښ�se��İ��38Z:��tZ (���X��=vv��-NФ��c���.a�-��M��%'w*��˒F�4?��F�\C��wW��r,F�s�x9X��ͬg��E�B$��R�����RnR&��مZw�N�KJ�c1F�(�Sh�f��B�aN���2�#�o��}�$D�}�� 7X�9��oM�����̼�&�D|������ת��Bu����ú��,:��b�|�S�dh�Ygv`��-w.L�ч�_*�x:�6@�@G�ېXs���Ã=�G��k����lu�bS��M�-n�)4���([������Z�揁Ԇm���]��U.<�n�j�.���cBb h
��П,�W9��*�f�/B�t�[*ݜ�י2æ�I��f�;o�����)�L�ҟӃ���"Շ���0wm�|�uw+=,�D�^�)K7��4��9[�8�e��γ-���1^G�+w=ݲ;QEs������r�µ�.˝/�����p�q�d�J9K-�����:*��n_So�gslE^��їt:�+콅,pҫý�WA嵙p�B6y�I�[w;u�{m\ةw.+C�
p�v����,c�q�;�V�r�ɑW_K����-��/7�x������e��[wA���g>R9�������&�N	V�jw�;�-�o�[*�|�m�)/�0�=��qd��
W��ۉ�WmYm��v�t��g1Rd���wNw����K�����&��6��2�oe�%�3��dv�O��څ5��-&J"��)�[�C
��}�]kb�;3U .��sVK��6��73�,-�%YoM�3�������CM;Σ��ݽ��[�S��q�f�l�K9��{�7�	WՋX���6%�NR��W��jV;1�Z�u�{���z�\w�Rq�xW�ҙ�Zy�ie	��wl�,��ȓ�0$�xk5L촫Q���c�8��:��J��`�w`���gIԧ�`[}F��_O�|��R)�|h��jW:PQ��۹����	J����5��w�y�f�\�'�Q���H�'+���N�:w�{�   ��?��{�C��˧����K��]c���RW<ָo�l1���8����y&���ֆ������`nЗ|+і4���B�����*)�ٶ�Rt֕�M���'A��:��M�[�c֧8֤6�0�i�ܒ�luͷ�s�a��}L�{)�2��W]��b����۾�qm7�@�n�(���nG��5�(�����'�C�RY���RW%��#�	/wi1݆6��Ӛtn��[ �������A.��5��&>�@����RȆ�ٙ�)�qBK�a=3w_��<�6m��F�\�93����BX�;�l�V&�0a��n���=[�B�b|�n��[F�nЂ����(�i�?s/x6A�#��n��$�1� �#�j��O��:�����(m�
�cV��]�Ԭ,���i��>�=�uݚoa�h9���Yކ�boo�q�<�,��`���!xz�"L"C�Y��~oN�ف^Pט�m�<�Wu�I���C�;3-r�j���dru��ŨjiGձԬ뛻�"��Ĥ��Ů,��n����smk#�ր3E��^k��<�^)h'�u7�w����47��.P�1������l�HJL�F����twP}­3i�G�7��M���1�Xr�	� KW��c��<n�f�wXNm;;��
wlD������HII����bی�4n�(Q�uӓ��,4�y#L�k��O�^����2�57��o���3��+�ɬ�+�����ݻ���U�H���F�ᤌ���v�U'F-���^|mo`�	����)g��	MӋ��MEo>b�������p1����-�ʔ�<4;��4Gg����Տ����Z=L|xs��a�nrݗ��L��hS�	�n�=��tS��ׇ�;�r���59xj��'��&5]0CjmJ:dV̴NV\����0'��r|���Α��e06]t��+�5��N୧��ZB�A�b�CN��x��$=L���p�����Bz+�ǐ����n�(��:�����Yl-��0�ph;�+�>^U�����%&/w��M��`��ʊ��a 1���:����i�5
_ܪ˸Y)	�"�%q�5�I`���f������I�zLȸ����sG��>�z9?��ǡ���6�z^�՗w�6�"M�ɂ�vp�ʝ�s�4c�#�Uȁ�1�a��%�tm��b�N�ɥlg�]��d���ˆ�h
,(-ZGY�24]�{OyD^pS�>s�#��J�ɞ�c/�II�PwI��l
�����n��*Q��v�2n������ܫ��J��Eh�W�a(y�|Ou��p	���(t��ɓX���cKm1e�K7Yݓt�mP��l�u��"6$\쫶)�V��4�1�;u�S5��N�;�����9Z9��XV���+N����V��뛭�YϠ�Ɖ�L[�+D177�޻ՙ��;�877��F�P�N͈���3���&��ʴ���ƻ��B�M���D*�rz
w�:<��F�>_2�`W����`��yE�`Ǯ��|�+��n�Q�Y$�βš�6.�ִ�Z���/9��<�*s���(6{}��@Fges�{�ed��kUlϵ�����˟y�CJ�����A�\.��ٞ4��4��v!�X��{M�\Yy{�l���EW"z���F�FJM;'�dW�kT��uǄq�v�{�)�}�o{�`�=����\Sl,��ށRKy$����͓Wt��J�ǧ�f����7i�dMü!y@I�s(���Z����	���[�)�gX�1_��^LgT���`��s�@U쫢�v�`�p�)�+V�\��&�mv���h���3���p��9��7���S���=ٙ>u�U�� �Y�^��&ʺ�u��D���=i?��v��$U�g�_P��9��q4Z��O��;MZz�!�S�[A�g,d�i<���.W]6�͢-7Հhc/ 4�n&�k�u=�z���#}8��;7ЉJљN�t��N���	�.u^r4�<Ř�8Z�tm���C��c���v�m����a�Rܺ�w)�o_l�W�"�z0qC�v�}9f���.=�<�o���I�Z��X嗫����U־��76U�И��t�E��0w�y�����(�3��r��9K�O��(��=�b����E}�]���j#ufQ��Vx<�oU�8^'��n�q3)�nrV��q��d��WŃ�a����K[nxMvb���
���z�Vm�e��RC2���g_�h�q��(	������_.9|�����
��v�2�y�g_G�趛�*�3�7Lͳ�K62��D����~ް0�h��g��q&n�'��J�Xx7�����P����p�׎�w:��=r l�����p��R�٩�Ҵ��*W-�CS���([�V[@�)`�{O.�B r�N�thf:��<oĜ���j��<����V�����
Kl������ZŻ�k6���z���OL�\i��'U�V���hXD)��$��{��##}{�F���u|�}��������ޡq�O#nnP�ۦ���Gb�D��3~��ɡ1�S��h�{�+NIz��W���K ý�c�ìi�o.Wm^�ZS��3*����u��.9{,�yR����.��hL.�XA<�7�X��R���=�5����7�Y�I]���x���[���L�Y��ܯ}z��g�p���h���q9�ڵ�l�iv���U��gg�R�q�$,�ٮ�7X��g��q�`�Gk8E�[�rCs��lt��a����`���v�DɅ�[�����T��:�i�0\��̴^aTHDW�w�ܢ������Jl5c����N��ћ��/"��s!e�z���
0�9��Yٗo��=�o4�;s�(Q��{D���W��g(6�g����Q�"�j�y��TWZ�	U��v;s+D��Y|Un�j�c��m����:H�WWU�?�5�EIF��	���s�<�=�t8;�
DC��3�c��mݠ�ш6���n��YN�,ɳسro�||ȧx��\x�.������L�څܞ��p&��wN�=���y+�ik@ɗB�y/����V�G���ѕ8ս�[�rה�JL>}[B�۫�(��elo���&e+ot�7M�Z5� �@����M�Z�k�ph��'�nT��v#�f��2�[ut�w��V/-4]-庎�&�������v��l��]�=�]K|�۾�+s�������Sdʫ8e�]-��{L�	�h��N��S���VK�����u�ɩ��y.�)*�{u�J�Y�l^+o6�t5����qAY�k�*�/�]�Tv��������*�Ts9c��pa-�a�� �1i5!�>�nO�X:�%�6üV�n�i	b7Xw�D-l�|�*k�{�*{B#�}��y�qႷ_7�.�����9s$������v����ឭ0�p���>�6_kV���3�0�*N�bZ�
C�O�CES�Y��u�n��=K�����V���Z5y���3q�!�s-@Wd���i�;RԌT�;���1�����s���[��P�0�-��0G+g\p�Y����k(ަ{l��F��t�)LժTrQ���kq6p�[���� !z����f���:�F==e ��b����w5Z��8b[��+��q�Ɨ,qf:<����tff��M`�aG+-ަK+�)K�������y�z�S`�5���m\�N�̋%s�3�]��|�_��Q��n�%'�}x��
jﵭx1V���R� F��ʎ�\I�ʅm>ݤ�}Ϧ=}H�j�e����9���`2]2"8�ӛ<s!�|���ʵݭSa:J�˭
j��ZX��6^mre�w���|h�W ����`�)aU��}�{��Y��q��N�}�gT�ײ�8o ��"��J�
q��|��>�hp�Y�%s���/�l�S�|�뚥�n*����y�ܕ�2� -gQ�z^�hɚ(�8рt$��|̊#�\"��y����f��0�t҅�	�-<ї����>���{��X�vvN���\��;J�w����
����l����@X�M�����@�R��./.Զ'&w�j`��J���o�=�g�I�"c"�F�Q�[\"�c벧��n�y_1����˚"��ة�"��9�ޏ�b�ݍ�e^Zb�fW�3_�o�����V=� ��̕��֭S�k3������-w�9>�m��띆pG�a���9wV�M��	j����N,]�Ġ��]*G�7��:�d�{kt�S��SW���ԂOiiT���<HsY9�m�ڔ/�Z�
��s)���i�J�ܴ�šY�$F�"��CU�b2sOݺP�Ss��Y,;]�i	F�]Ң6�o��f�#���m�_k�M�}�.�ō��6��6�p��i�^t��b�i z�u�d��qe��8e��i\2�\���5��)�{*���Q��r�`��ނ�w����5��.<b	�A��h)���`�=:���h^��$l�Z"�:L��+����C٢�鋕��xe*�bK,������6S� �1��`��Ĭ�{j��K�;r�M\m1��nm.�}\A3D�*�7����sן�'�-O��iA�z��bͦ����Ϋ2R7E:r�k��Ge73iį�P1e�Y�ۀf]���I�w-�>-0nm����oe����ڝ`e*��3����bS-�l嗻`V�0%R��	��8 ;�U<o��"�=	�7L�Q�`dj���v X��v��⦫!���ڹu����"㐴�dtj<�L�d�I�
��$���va�&Bq��&w��pi�K-4�hpWyRv�S�<1�'�WJ�t��{n��.��[�����Siu�[�1�g2pY(F�[+9�M�;0�!m�|��>yh�9��XL�X���g����)�[�u���w;���ns����5uB[Qۭh�p�Їfkz�q�k;����n���8{�2-��ʪ�v��
����i�lR���u���flj����c�Y�!��Q^�.�.�c�=/��:��T7�t�`�o���kL�75��FMv�{�
+^vu���0;��#�i���[#9Ԓ;{-�->�K*ζl^S��C*��u�\񳔢��r�Ж��󓶝e�$Ǖ�b=��o��:�2L�yM�nw1��Nmй���]H.��,��[
Ֆ�<mA�y��r�}��y3)�X�Wk6Woק.�ϯJ��B(�f�̝Qu�kM "�zv�*����X܉d˹��t�٬'\��Hi�J�->ܽ
�-�ߠ�Ԙj�y�"7Z�7V+����(B��"7x���>LU��$Ȟ��R
���ʯH3e&�
p���v�s5�뮯T�.*4�ӟ%�j򙧉��V��I�T=��Ƈ.�Jv�$rn�1��}"��n:�ie�3
Uh�]�`<؉m�{`$떵u�r�řΦL�m�ӊs]����֝��i Z�޼��H֟D�&�n����u��C:�k*�/*[KuvQ��W���b�mW�L�;�%�/u�BB��H��a����8Z���2��+�oXW�$Z6M�V�v��]鼮|-\@h��%لM]�0b<�!8L'{�9�-���N�
��̑څ�j`@���(_�ݽ�^Y-~�����v�XGd��.@�֪�!��v�+#"���h��h�5D���tU�Y�n�-wɡ���D�:Yx;Ospѽ�"Uݺ�X޼�m�%��M7�gM�"��'�0�˺�"�{�o�C�~�p�[�X�y�8�h҄L�i���2�(��.�9E&Gs�˕����+{��F[��)X����K����� IG�4	�(����Q�!�qn<�֠+��K�5��l�8������-{��6ocv�ǞUMf{9�>�K�F�O���`*�&M�H��ܢ��i�Ή�hg��V�W���M��*�����Kx�r��V/���ai�+��o>2�|f�:��v�r�h��\��c�cj�.*�H��;s����y�rj�h���e[�s��[o�+��8q���>�# �d�$��\;{��ԙ���n�0V�8�vY��	��I�ܖEZ���sc)r�/S.��r燶�'�N�c��C���;�F�Q6m� DE'�C�pOiӁ���X�\fV7ô.3���=���k$V=&�d���Nk<
�̂��vvRw&��2�Q|��P�FqMx�]��bY��^�f�q�Ұ{�-�����ة�K�[�^ {� VxUq]�*���$wzJ��N�H{v�z>�sMi����ԥ]N���Y�E!Y�[6��γ'��4����f�SI�As��V�]]�y�W�C߻���NoQ=zoka(���E0 �\�O�,����J��flH��qQ��Z�EwΚ;��C�x2�R�]*]E�U�s��X�0/���`�f&qC;P#K��0�9�YS
�RV�����S���}��ErSf.����ɺU:�`:���+�5.f����ыn��� ����"'(S�$L�e;��+�S45��b���5�X౓yV#��hN���o���.T��9�Xni���|�����ٛP��K�'{[Ԡx��*�6�Y�U�"��Wt�]1,�K5�c_]b��{�0՟��`Y��dR_�=b� dŢ�x���f�~��X��c-��b�횜��O�V����Y�,�r<ӹQ��-iS�y\"�5�7)�UE��3-�W�E���+��Q����wS mT�n}��qm4��X�"��>�$4x�n�=�T�7m���D���� 	Ot�/OΣ�Kpi�B����<�
{��-�V=5�h�=p(O��xxxx{ޟz\��}Ҫ'����޽q��g�mV�n�C����Ģ���-ڱ�z�,�Z�� K/$�|�����mfhO���Nj�6ӣi�f�4RVV�Ѳ;��ӗ>+�=�}�"ʧ���_Fc�����:e�zP��Tڌ������4pY���gH����#Xi|��]�{�j�Sr�����#���{I�Ƒj:l\}�0q�T|�̖p���-�%R�`�;[xe�{�F�5�,�V���涣�#�A�e��8^�B�ԹQ�x�����֕׎�<Ӂ�>�4q���t�V=�E�L�d��9fƨ�/Gm�5�oM�/>�쓔\�����e��T�j�1h���2m�x\������������bѱ�)�;4� ��B-���1���]k#>&��&rR�d�j�z�=���B�0FǪ_{��#��t>̫�Ζ�56��)����@Y�N;�����o>�N��u��:�:Q>�V�_�aE�U*�X�ڞ�Z�y�@��z�wHF���a�\^��uȑ�ܦ��h�Tt�!���WEj��D�>.���{�R��ъ�j���T�ʾB��N|��#���&�|�K7o�} ��Th��T���D��7GpY��]h�,}�5�`�yE�h�.�i�-4]���njẞ�yLڈ��i�l*Y9^�:��OFc��3b'��3�Zy����`��$�)$ˎ�bBI���h���ds�\�;������w)���1���J(1�bi�d��"$�RERI&`dDІ��.
C��d��3$A�F3&�Iwv]�А��wW
B"���(MwvJa�p�ԖLQ%��,0��&������6�C&6!&h��BbB��H��d�E3��!��Q�3L�$���$F�r�Q"X��I2c��h��)c	!��a��	F*�l�F�,�2����1��d���t��"��,�Ii2�ɒ4Th��l�S��������+�u<�I��'Xx�3�*ż�*�OZ�VIW�zyM��_x�¸���� a ���r�̠sV���^�܎uo����o��/㊑�v�B���F	�0���aU(��_��!ث���>��h����B�[μ�P��s�G�0�{����-�q�-�_yM�a�0�ޖ(ȓ��z��c��l\�<�%!�
Ш��e_s��FT��ɋ���3&���W[�JX켿Ztȿb`�XZ˂�V�E'B��&����r
P�>��,84��N�5����fr���2�XQ*�#����W�o��^��_0��
�I-�^��$����$��r.��.7G&ʧd���b������L�s�>ޖ��,�F����m�u�i�3��+�8+G����(c���o.n����DĐ�a���
���܆'�v|���k:IӨ�Ek��^��!��\.�Qot�����-5�e`+�L������qi�+�FE������U�M!��>�ט�`����Fd�Ѹe}~V����CpʈK����+�'�x�t�@�,vT�?<�D�.Y+]==�+�855|I���=���T���_Y�a��3LJe�D�Y�އ�b�^u).�>��3�l�1���[���fr��,:�֬tj^6�^�a���Y7��re�9��Y�s��C������"�����{�u,i`��յ���l�̓t�PNo�3�2��ȱ���R0�����B���o����x|z�@�=�޲�;<�ׁ������_�V�q��3o]��d��s5�w�mFX&Cy���m#g(B�2D��H)���]p&;+r�˫�AYZ�z��5��u��9�ګ�L|���J(!�֚��D�*�y�2���܊���!XH�2,bi#W݆�t��w�e{gA�鱀�@(J�q��5R��Y����?��fVÖua������P�C;:%�\����4TrT�B5�T`N���g��u�[�yY���*�7�ͅ>�����ڊ�/é�6Cԝّ~��d����kݡ��]�k+�^���:?X]������}t�7��^X�Z�}g�����T<���2+'}�v�K[w����f�z�T��%	~�}o�n�b5�88X6���yq�	�q�f���^�1G���=���͏i�`�3G�}�\��I��2�C����)X�� 
";ݏ��I#8@swQ���gt[��L��q��6�Ȳ�vMۡ����/ex{�s(�l��V$���R飈n�3$���Sr��]C�}�Q�)FV��vR��-`})����]�����ւ��^�v儱o ����kHX�Z�]��P�y��,�1ֲI����r��3ni���<���e���첼�3S��b�%�YX�W�Ô�W��=Cn�t��&�Y�Z��m_���U_p�(G��r����ttU�� �\&pt���Uާh��WI܃�{�KΏ@����Ȃ'�˖fӦ�g�W�Q�%yp����+�f��-����f`}�ɀa�"�ɦ�b�0���aӋR����ʎ�L�SF���|������I@��sO�&�-%�^,Y�b�4�"�1MH�����t:'&�eִ��dc�A�����->V�3OuEOq�~�8�D���q���D܁�\|��,x�����P�����%TT� �0>�~=�0�;[y]��?X���G���t�����*��}exI\���V �O�{'IGDT���:��ڴ��fj�wa_ cj;���h�;����5����	�� �R#�}������鱧�s���{�0��h�4��x���!q�2c7�YEk~�Q褨��[�~f���4��]�3�*=�8�X���Y{�2Et�ɐY5�)�㊲r����dJ�m�r�M	&��#ue{�1�mv�o�Ni1^����L�Ҳ,��ժN�*���I�ep��v]8=�?�Ӝg�=�����n ��`돑��e�'qP7Z3;S�ʡd�S=r�8���W&��v�����@)��� W�~�������D�t��+�G;�W�^D`f��IA���L�T��FA&�E��n�k0�P���]Ep�kKl`�׻Ɋ{궅??����q��o�:)]+ߐ�7o� �A�6���w� �2g*8Zʤ+}	�\7�z㥃��z-|�V�D�a�m�W=�OC�}�N,!6h򘌊s�l6O�֝s`C����',U(����{eq�����6p/�d.��
{+G��ʭF�;Ǽ9�"�?w����د ?]� �ԜS���m�/E��R��U�س!f���u#��G}�*д�z);Ir�o���!/T���C�U�{˦��j�M������ٸCX�C��H-&�Q�����V�Dm�tz��s��o�`>/�:I�W�~�\�]�ICx�����Gj7��Q���ރ�¦xAK�]�=�9�qg��Ʃ�@q컹�Rt	G��5gO"�./���=;	)|�T�͗vR�����4o�E��*y{z��;)_�O�+VDB�ebٽ�w��|��k wZV��/�+�,4[�N�k��PwM�(���֪;+	u�i��w[��У4]N��e�n��{m��<�qd�Y���{u�Ltu�:��w�ު�'��IL!�}�@��^W#�����F|��#O�*A^���b��[�&ݠ��["�v1�b����m��3�/g��xȭ����XD�ShL@�FOR�.^��_�m(��_ hM�Ǟ*�p�V���_���y���
�q5����.?+y�kS��s��bDn���Zpy�+dQJ�s
-O9�6ze�Ӂ�-�:"�-�7c�Ǻj�D����&����e���x̦k�ӫuf���6eEm�2*�Y{
w�t�d�o(�S�a�q���ڪ���~Zj�(<�e��{����g�<4�cc�v�������,/Omߴ��c�y�s�����
�!�-}���v��ݞ;7�ת�#���Qg/׽Al�LV�A�.
�V�E�\R��	�tk�y�k|f쾖��A�\�j��̭�S�>t�&r�S��e���'c�:�(>�����cg2k&I/*aM�B���ˆ^��"+X�
<�\`���t�`���+�_DŁŧ�2���9W٧�W��.�]�#&��"�A��)���x�%�ɳv=�X���󡯳-\kR����9�ԯ|� d��:����`�Ώ<={�[�+h�Ɛw϶:r�m��)��q�a2�n-[�d�v��n���V�>w��ݙ6�t��,R��v��ub-M��]�M�zU�,.�K�;�!��3�yD������m��@��f�jS^�2���2p��R��;�*ή/�ݳ������:Iӱ'�ѝ�����#�oɔ;��#[M\F����7f��s�k�׾^���&��V�o��$�K C��V�\�}L#L�m��Qq�#}���%�r��Q�0G����#��.3�B�p�۾XB͏=�v���:�bX��t/ƨr�)I���献�s;��J����lӛ����i[1m����� +�X���寨��P+����K��
�tny��3oY�����@k��s6����4�>��yCMi;�Ht�x.߄�eF��*j�d�<�ǌ���s�v��N�1�/��x�Ґ �����0�=�ϙ�W�z�w��p6�8&���5���3��}���U��"��%v����U�]_#��k�q��8�K���]|�+e�NO�\EG)Nd�و�x+��*�8<�]�>����}�%ad��K42�j�O���QB�H��څ.6�B1��TL��P�7��b}�լ�e_n��h�{�7G_�m�0���mby�9�ӏm�ZiX����6�����H�lv�Y�+w\u8Wj�K��o2
�̊��ݖ�ܻ�o)T��_-��.ks�Z�ެ����ז�ّ~�^s$鈝���e���+O�l�1y�Y��Ύ��E�2��r�U�E��RaF{x���s1�((�L��M��|��i��:����zʷ���	�B����^��}$B��ÅC���!E����M�E�qV���u���x��5��nR���z�1w�	���_e(��G|N�\ �|\Y}h�1O�es�|�{�
�plC���nL]�����+�^�?p@+F�9��:�Y;7� >�fd=C')�j8����7�=��Q{�j#��_p���̾R�_�FtmKGM2xGA,���xj��OOE�D>0#��w/h,��~C��hN%F�JG����<=�����F�d���7Ox��bё��q)D"4��	�ʳ�(�W�ˏX{������*:�ׇ��(�8'�E�栶����d�e`
��>��uI-����b�4�#���<�S��\�����)P5t�r�@}�iV����0�W�}9����H�t�٪�D�dV�J�D��3S̽�����xy��1݈|k�>�)y`�T�0v��U���\t��؛�ҋkͭ�1��e�8߁�i�wcuS�q�M�nu0EN�-�����H�b�N6x{���4>���<����.�`,����ޭ���˃ڳr9Rsʴ���0�ׅ�^�{n��^ATxM|�QSq� 8D`��P(d���y]�O�+69!�9�x�z�\�{�==ǉ��Ҡ��p��qJ�A����(�(���W�F�ɠ��go�������F=������1���M��o��
��E}2Gi8* �Y�	\yL�-tى�6H#%�1��Gq�2c7�YG�f#˄�ǒ����#����g�3:�^Gvv���@��2,S��nB�����,$��XR�Qӈ���..�U_8��Uy�1�"��ۅ�*�ς�?5�vg��
�4��^��u�=��Vv,q.�^�m�^_���z�8!j��B�[궅<�xE����!_��`##��ղ�����o�}÷��U��(%a�ԨB�U![�O}�Ἠ#��K�(=#�ý����DКC����}gz�>�N�@�V���G��dS�Sm��\�z���֧t��QT��3��l�~J3ax�j�<�ǣ��|hZ���CH��x�)��/�,���.g�5ͯfl�6��N�Եn����|���Ooz��x��ޱ�ڙ��h\�7��J�����w�ubhgx�[Օ#�,�t�f���Ҝ��xBȁ�����R�����F�X'{qu�|k�r�o=�kx�w�ͲL�2$gL�Z�-p�2��;�� ��t3�r䶻]�����`�~��D~LS��q��Ƕ��Ҁ���:���rT��:J�[��h�=�z�[
�z�fG�p���ݥ���_N�Q��P�l�y�A�۟tYzƷ�.����������\t��⾢=���+�Ɨ���R5�f��g���^���.}��3���o�\7Ҳ�W�|Oq oN�� h�C�����=�ע����7;�F��X�c��vM��t��QHx�,�8���WP{>H�+��6�R�l/y�p�N���"E���f��x˶�g�se��n��x�ViwnjUR�љ�v��#'s������"`k�ܦ�ҘC��<6�����_R��>�G�)'�e
&����8����\]ԭ���"=�@���t�a���=̈́p�uϊl�˞�sJ�¶#r��:�`��� U]��ι7�eiD�L;5��Lׅ����K3�8;���k��^���\�o�c0�!}�PW���ˈ�h*�:�=��Y��=y�S=����e 6��G=�:H���GP�!G8�'n��+v�ՃT&
k͋�o���u���0�o�>>Η!��4��p��ݮ��n1�i-�4VV����t���m;Y�hY̢�kv�k��ł��+��⧨��)���kʱ�rd��"7ɼ������a�6��V�á��W;�9<���f�J����E��c���Z���k����顴���>�}[����'��Q����*�&9}T���*):�ƺ�����]�om��B�h�.d+5�|iVL��)DV[�
0"NǬ$�9����Z���==D�u�|Z��骚R�MvʭW��n'eq�"~����\�}*��x,�73>�`�]�!�Չq�?M��S�we�Y�=�~�$����������@���B5pJ��"t�s+Qa�P:�L�lo=>��\cn��N�;����H״�]Cx��רS�w3]r�@���Y�����e�Q�>P��;Ⱥh��Xz9r:d_��  �2�m�����h̊K�n�"��+�J3�T�v5HEa����]u�+��X�aq�Ȃ-�]�D�j�v��~�W@���Y���H�H���E��iN�������sl��T^\q��\g���� gQ�A� <����P�g`��]~�V�p6{�c��./H�ϼ�c3	v@;�W�8JK�9�g
���w.�̧���>Of.[���tE\]���n8�J�}Ʋ�sU&p����V�L�2����St����&�H��]�OeAr�q�	q�G=��Q��y����'��"�;�"N�ֵ�+��{����}珕�e�Z�َ�
����"�syF�����x�V�t,�v1���L��S��/���%ӻ#���u����r
c-��5|:߆����!m}�E�w��}aӅcV��ͦo��D���ۓ��
�.�3�̒���r��2n�����{N��Q'�6�c�X�Zb�*ty{%#�2��:�7a,ѽ��8�a�����!S��3g�IxpL�aJP�����+1Q�A9�JʇM�ww0V`�N43:���L�Fnf�`v���� ����p�璷Uk][�-���{rW���� ��n,8Ot����k�m��<��t�m��Lp]���&�j�2��/������P����g8�53��|���.�g]HZǵ����+<)T�,3sy�!�>Z�SX���~發�č��sX�63q"!V9��#˕^�'n'���b�ᗇ/��,�֚�A�,�^�C���݋�_��/5ҡ;�<t4Dq|o,��0)E��G31�/�0E{r���B<}�:�:�]�����ur�Q�8�'c�^:�-�wj��@0>��m�B��yqP�f������'���	L\���T�F�ZV���fnt��ؓtv�;��>S/"m�1�3��ȊT�B�>���ts�0�{�lHx]m�s��:��D�
	��g��ċ��G�(t�+ͻzy���qI�b!&�m}�c�9JMӫ�8)VOYI��v�:C����Z�m���nL$�i��\Bږ�I��lܚ\�MAU�:X���Ft��M�Z6M�y�Q{��	�O7�8m��:�mF��;P�Wd��;����'��B�&N�n�nI��fi��\b'r
�ke��M�:�}�l9Z�Z�f���g;:_}���l�`D_C$�]f:yud-:�Ͱv�gt����״���a��v��(s\K�c.�I�h��Vͭ7|�@r�-��}�-Ը㙓D�������q@i%��l�6�h�/Nf�Jѣ��t	���ۢ{V*�5wP��7��Qrܻ�,d�i�>wH�ӛ\U��@�"̝����\�a2�|R��+�x��+Vrk3p��uc��lN�kQe�Է��^]4r��?!�7M��(�XI�⩊��{B�꧍����l�o�䧝����(��$��*~�X^\({ޗq����j�ݻ#RĐZ��̚��WI`�w���CiwP������S���㌌���w�RS8E ��H���[Vl>ė/���X���c1���B��z�yW�l��*�&ݬh����
�R��m�G��T��O��j�A��QF���L���M)D�#Hͦ0�&1&fF�-!�����Q�eh�0��t �lP(��w+	S
-���lAlXB�F��LlF0Z"��Q�����j#��#Hh��RQ���P�I&$�Qb�b��APh�A���a���-�cC�����I�(����
"��b�#`Lh6K�hC��$��I#! �6���@ll��d���hƢٕ�$QF`�[,cl@RFB0�0h�$X��2i"Ńh�!����DQY*0S5
j	
��Ĭ�oxֶ����ݐ��!36KS]M=y�*^����3}st��,���8�R��Bs�ܞ�Y�m�r'����7�ݺOZ�1����|	�����5潷��h/��k�+��x���^wlno�����J�so���_>v��r�r�/������ίKO�~��.��z` �L�y�G�{� nV���
RG���r#x�8���B$�wb��s�����|��ݯm�ۻ����+��~-��^z�]���ʽ�u૜����;W�ڿ^7�Ϟ_Z�����[�������~���������s�����ȶl;���DG������Տ���6����M�ۼ��g������6�;�m��*-�W.o[��+��}�\�+�ޗ����-?s���m���ߝ~��j5�y�����w�����~�d����\��]���qc�",}"#DE���O���:=Q����"#��U�oJ���瞾u�����o>��W���_���|���~�W7�?���W-������[��������*��k��S|7<sG:뇴�B�-qc�>���}�w�����O��忛��ߊ�}�ߝ��8���`d�8���##�#�ţ���׭����x����o_{csx���2 c���WO�P ��ޔ��rs��ng�/<����q G۽�}���_��u�o�ܫ�{���m��r�{�|^������ y�����<&<�ޜ�w�}
�ѿ7�ﾶ�ݷ=.[�����*��~�z�eb�m�rQoP7�0G��"����t��p=�* �������u��-�h��_��i��}zX���x�}��s~6�;~+��oj�@����Om� y���}��<&=P�����}�h�S\¼���8�oJ�߿|�7��6���?���~��j=o���� \N��� �@���^yzZ7�~7�~u����h7��_�z[�\��]^u�����o��*�����Ӌ��w%�ny,��DY�]Yɟ���ʾ.W��߿V�}�\�;�nWջ��^����[���_˥��k�7�nk����{���o���7��+���z�^��ߏ����-��7���mX�DH�#1�����5q8�ּYUy�������w��y��77ǻ�>����soW���[�}�U�Ϟ��������:�����~7�����nm���/K�����m������o�࿼�[�1����qB'����g0U��ܟ�>�5�����ے���.�/wDH�����k��)�e+��ic�oqMi;�88��bJ���x^�����Y�!���Nb�D���R���K{������I���m3�{\Ea��w͞'�&z�<i��O��oy[�@FG�Ǯ<>�ϼ��0<"3�#���ݷ?�7�?<��W�-���;�����������}k��ok�Ͻ�������_/|����W���<��k�^5{�}�`z ��=���[�+}��l埿?�>[�\ۛ���v��_�z�����&Ǽ���S�t(Ae {�V6Y�� ���08��9 (��f8}��D`�L`܃m������b��|oM��E����W�|W+���y���^/U����sN������._׾�-���z�J�������=dl{�ޘ \	�t}�����=�}^ E3��}">�sQ;�)o�X[ٚ���@�G�Tt�Ї#�c��u_����F�����~/mzo�ſ�u_��z��KO��ܽy����+ߝ��������ޗ��~6�w�߬{� xA��Of >_�G:щ}����7�nk�<���}m��~��}���W.~��^����z[�s�{�}�^ן:�7�������}^�|\�ۻ������F��+��:��;�o׍�1�H���k�M(�w���:�>��2#�쁱�P>z��<" �3��q��
m���~ur���/>���{o���_�|�������_������\����K�o|�\��׶ޗ�|=76���4s�Y���Fn�L��{��Q�E�sW�]����x��w�~]ڼo�7�,N�`T�8�h�#�G��Q�4W�=-��[����^��o��x���kү��~�����[x��ﾼ�Kzz�1��v��z~Ӛ�X�P@w�{W�������*�������szm�}�}]��~7��ۖ��^-����W�:�7žy��5�/�������׍�x�Ͼ���DW���|���i�����4΃�b��Z�oZ���#�� 	\��;_��߾�o�o�F�Wۻy���+ŧ�|�[z�ۛ�z�|^��ߏ�抾.�~~����}W?�>|>�@ˑ�1��>����A�`x�s�QUx�#{L?���Q�LϽ0��Q���6&,5^�����-:����@1�Q5���/KF����]���o���{�u�oOƿ�_�}�>ur�������� �L{cޛ6}��T 	�9�U	�qM��5n��Rv?li����*e�&nS��dɡh\7\"Ē���A��F;K뮺��~lw>IWR�dO)�x����8���2�\D��ڜx��4u��9k�V�A��§a���4Qyg+dz����u��EF+9r�杊�K�D�g��ɘ��� {\���}W���7�ܾ-����_~���{m�{��|��^���~���n^/���wy��\�U��/��~��{Z7�����ֿW���ﷃ_���)8����/���aoOJِ�����W�P>ǅǽ� �ǆ�' 8��� ��E��#�?D=���E��#�g�c�~��~6��~�~/so����ץ_Wy�~7���5x���x�w�~+��Z#�>�2�����3W��Yۗ�~��?����|^5}��������x�߽W�b+��������;o���׭��W.�z�o��~��_�|���h/�����G��* '��6=ꈏt{Ӂ����>�c���T��J~L��~z�ߗߞ�����s�_u�/CQo��������Z�����޻���^���7��3�s�*���� *��/�
��!x�6��7������{���F�_��|������@u�<�w��m�74��[���=5���v��W,~/���W�����y��o|\�^���׾�{�v��K�|y��~uxޛr��������ѹ�?>y���z�p�>������"DG���rԚ��u����Ǽ�[#�c� l�ML��P<"�N ���������k��W-���b��[�^z����m�W���x׋����~�}�/J���{�?|���\��w���o��x}�q~��܍51q&=�78��p}�~}�~;77�}�߾W�_|����ᨷ��x�k�5���k����<���x������5�������y����^->v����7�ż�4{�G�<���>�R�Q�3Rr}�t��"D} /ξ�ُ���=�P�}�DG�<3~�p �ǽ�Q���/���|\�o�����_ᨷ���y^���^|�_��76����^��p��LE�D} O�8����{��+��c��
��f��lT{ 8����������τ�P=�* �^���>5��??~��뺹c�{������ ������8�� ~�=��ML���#����̐#0�;��{&��P��g��ʕ�c��
�^�:Y>~��3�z�X��#z��J�\�8�d�n���n������"��ŝ�����c��!��'�CU���=f�fgaJ���g=�M�p�37�����^I*)�w

e��1�`�|�XK��|�U�2�4ߟ��&�UPγ����a諾�S� {ެ�㋝�;�7J~�1DDh���ϫ���p��ʸpG�� �"N�w���ŞO��-��ox�1;{b��i�3R#���py�=�����G�<>�ʷ�c}�\H(����z�����;�DE�����G%a�P�]��ׅ����R风��;2������9UѸ���0�G����|����ig����(�=+���5��q��4~���Fv��'�j���ʄ���1Pɛ�� F��y�(�']�N�h���~�|����e�` �ᥔ~pW��K�[<��yUc���e�M)'�L��Q�>n�^�����BՍ�_��yY7g�˞�
Ud{Rg���s����7�4�w'�f��^��Vf��U�U
�<�ٟ>^:��-������h� R�����UBp�^m�f\��
�a���ߒǢg�#�u��>+�U��മ {r�? )Ca��c�o0:�Tчz�Y�֨�x\�]�O�5�c��]3='p�3ソ �v��l��yA�x�����f56�͇��e
��œ =p&�[�>��j��8��n�O2/�T�qK���X�Gc1�YGv(�Z���É=u�̘ҁ��ބ���ҎwA��U�sn��k�5�Ό�|=�he����}w�B[݀����t�xw�,�2|�;N�r,SE��;}�c5�΂N��|�'�(H|ȥ��}7����Ū�"������o�/���9F�6�8�V9xmdR���R�r�d�~�ፐ@
�����^iV�ʮ���⅌Պ��j��o��?x�p��̏?�����9|	�t}~;��.���5�qo�;����1vϠ��:��i?O��^��G�#4�U�H�7�G��)��Gu@�0�ɏ����b!G���Pw/�8S|Na��Bk/3��RF<�xx�IV U���b����@�0w�h5��mT;�[]�G���S��{��{!�pB�$C�M�D����&�@��*���ðrb+{�=��%���/�E�?S^��;�7�}��R+zyF㒠5z���T�G�r�^�v�UyZꅝ*�‭����A���{���'vd_�ל��t�N�;1���L��#��q�FW)3�|L�0n�pCH�3�O�᪘f8f�d�� K�k;.�+"w]�*��d�\�I.�̈́m<���+(���w(yjiz<+�瓗qn�"{�!�:��؍If�{}���OCM�ǈ�|���3w�Ȭ::�O�f�u�{_���;t��r��T�,�{e��E��SO=��Cq�{i͖y�5ot�����y2�*�B�?7`�߹�Gf�|�8�Z�h]������8X6���u�p��Vv�nҗC*�Z=x��&�6=]7Ӳxe�BUy���N�1��]e�c������;�z���DΚ�s�/������$�r�ƾ��;�^��R�ע��k3�����.ļ"L�n�b�}#׆DGa^*��E��y�*�(�T�n�	�PG���z2�mi�	0�3k��p�z�D��g��گ�Y�A�w���3��r�ū�ܨΞ�<���27-����,R�����p��(W�������b�0��\z��.3%�)�{������龅!_ =꘻�>��<$��/�����i-�,1��xX�Id���6�ѵ���(9�ar��8ƃg[�a���Jn<9T���DC�����A{��;��DbSCB�&Z�����vYWKNgܨ�,�#�I�)L�=@ExG�&R";��t���o�g1.�۞,Er�������V�jr^���ݡ�Ɋ7�*D�kG�wmݛW�Rx�����]b��g�+���]bz���A��rge]l���wM9���A�b3o(�>.��iۤfn�ˤr�ݬ1N��hy���Q�����w[�s�k�|ˤ��#�2��ї�h��$�=9r�d^iy#�|Ö5�����rҟM$+�>�8!��<=�i��:�{mq�S�����#^�J�����[��[X��QYd�P�c��i����!Gd�2S���a)誑�rN��y��"�"��I기m��Q��C�\g& �{
2�}�0��ZFE�T�M�B��g�5%vb�V����+}N3'M�9]�9/}�\ �\W�=�*��9�"��\�ӬɿPޕ�A����tO��
z���u(*r��^�V!b��qB�VշF�1��u<DM���!X8[��<V .�Ykfh=�~At�����y�a���U+f�L�j��=���1���NH"e���W!-���)nﰬ���x��2��͍�,�!o���1�:���f�i�73$l'��#;�nLw^]�6�g}�\-�_y�Q��!�S ����o��{�Bf��m�:�9.wCs6�&��_+�
��]���<#�b�.C�Ք=�3� ��[��\�����s�y�J&Yˮ�~(�]�R��{�=7���W�k�������ڨP���<Eފ5)��<8T*�E��S�:�����үF���˳�$9���
���Q���xEm�t�ה���=[�r�P�TS7��|��}�u8V��3��4��k2�Є�ꙗԁ������wMyq�x�^���e�vlu2�@ ���_�����'�ҩm�s�u(����1Ӈ�~{7�p�, �<xi'r� -1�g��+S�6��z"!�Ǫ�����^�<)�e�!*����Y�~�1�.�vO�K��Q�L@����o7�C�&����N�O��vM�T.�� ix�,�jV9��>��<9]�Zv����x���GW� uz7��"G9�l��ga�.ۑ{/'���猊̇zy	�=1��5C��/�({kL� V�@�ؘ�|���7ݑܯ�)]e��[�*�m��P�q*n�׶ M��!�Xk�7��Ԉ�P@Q�Ӄȡ�i]�u���{���^j�7]ˀ��O�;)��R�5�A���*%��t���� �S^�Z+ְU=ن_{������G�����`I3`F)q0Ct�6^4c%y47ʼ�`?{K��0,���M��2�_14y�W���<K=�~�o@��k�T2f�
 F��Y5z3Μ�t4�(.yˬ��i����9������dX���8��lT���u�{S42���N��;�ʛR���(��v4A���Uo85p��w��w�MZ ��z�2gj�ܼY�e;JGq�����žD�t���ui�3n1+��P
�o����xpM^}���G�rboN��(��(HFl!JP����I�'�� �%Gn�����@��~@��k�՛����.Y3�2�E{-�'c���5���.'%���pk.�U���Hbt�EW+�x:q;2�/�m��@q��%��*�iC����~�	�͠yRa�gɎ�����dLg��<��ִ��nc9= ���=�g������"�L�tt����F�������Tr  ����\��3�4���0���L�D7$��Y��A>P�d7!SEƪ��ˑ�"����㵑�I�c���ص�]@!�Q�28EI�xA�[����Ρ���F��q�Uc�{���$�z/(+:��7�KAC��D��4�7wL\T�j3�?��P�OǸ9�&�p����$r��{�i��X+=C#\z��Eh����jt8S����l�������1������0r��_*ݙk]��%O�n�9*`CL 0#��uDՏt���?=�w�o��+F�Sҷ,Dd1�ݸ�i�#�����`��pdH�Z`�PH�'�mb��{������b�-����2�Lno\Щ�G�~v��33n+�F17�[�r�*eeOF�^�wS�;K)լ[�V��ڽ�3����"�� ��D�:e� ��p��I�d�7��:�����o^�cf�Os����k�{v�����sMG|<=�{�V�9�{�w�;�Ey�f���)5�%Z
�U���,	J�}Uj��+��e�m],w�#ol�z��A�z�[�WS��°�?dwmH�<����P����:)�<�W���u�F>��������
�r�?J��;�Y�ݗĝّcy̷,D�L�N��:Zܼ���rR�	���=U��5P�^�X�􇓐AU�E�eFFT�Q��/�OB}�w��䡛�;T뼾"���N5��Ρ<,*�}6�$+�W�w֬-�o_��طY���"2o���hJ�x1�Nv&�/�`�F���>>O2�f��ݱ4I��>5u��k;`l���2��b�9�t� 6�+F��p�Cϡ,�p���E?��Z5����Ԭ�c��wn�,yR�����2�9(G&T�P�g�ª��N�aAƎ裣a��Y��x������x���zUT�l��H(�a��x�UG��-_�+&���q؁�z�Y���*�Ӗ
\V���h\"Z�$}���8aӏ<�J-{�R�V�Mv���t֚��
�Z�k��>=������mh�U�#yU�;�_�IZ�u�ZNw'��k�ܳ��8zXV�4u����-�a��nqods6��3�"����2A�<�{gzߋO�����J��<�v!Xʥ��=���g6keѴn�T�%�H���[|$�T:fZ� 3�%`\"QvގX�֐�m�AV���o��)�:YV�Ïk��1�9�9��aD��	y�����&���%�_��R,�	�lNr�}yL8.�9����Ş�o	���Q�庥.��K�� Eaw
:����V����w� ��o�MT֎���
k)*'�c �ȷ�����8h2��]JΉ;p�N�+,`r�W�VԂ���V�9(@�vg`�.r\�5�z�];���^� ,�x'Уy)��%��hJ�癡.U9cկ��b}��0%�I��������߻��.��%�z[��s�:������]�~�˨w"�D��e��
��r�x���۔�ٳW`�N+j��b���sP��7s��	��@����;bZ��"N��}��t)�sm֨���w��j�68�=�r���� et;�x���诂[��J�4ɫ��Kv���˥0QG��G�B��G��~��%]ǎЂ[�9nt�۲_>��`�ي8
�fР�h��S�^����+�'7lv��M��ҁp.h�4���ʼz��Nǝ��CZ!����Ql[1n�=�[c�0�v!�,�C�2_���T�:��n�B[̬��r>Xz�J���L�z����Ng���W�n
��T:�C�N2��=�])��C���#7yw0��=�2��ǡ���\)��c�����t'8]meƝ�V`����7N%ۈ=�+�fڰ�*R[�s.�S��Ս�Bt̋vբ�Щ�b��]�Uw�)�O�m%u�{Z"nM��#�ӥDu�pv-���
�h��4�8Oi�r�d,X*湜r��G򩕅��}��dK6�z���]�4�R����{v�k�D!���v����܁fN�%en�叟�X������:<ޜ޼�V���/���]M��T�u�Ǡ��̵� Җ��Kks�4tV��XZ�w�	O>��)�{M����B<�w[�w���K8��vy�ڒ���1Y�C3]�dxM��".��q�>M��"��'��7���$�'�?ziS�5�rB�[�/k:m��iu��Sm��ݲ�m��/~�G������@h�,�Q�=����D �#�^^��]trg�]\�
�vV�F�Y�e�pښ�=����__X��� Q�����E��g���NX��Os��
wsL�F��X#4=�:;I3L�c�oo�+��Q���Y��鋼坷p�{&	�3�ujjZ!��0a�wv��ڈ�Ɍ
uB}v<�{�������N��ò�7��^�\0T�<-r���/T���{%��$ O�~$�2�cQ&���$��Lb
2S&�m�LL�-Rc��KIi)��F���̘,
H�2Y�$ƌF�ƋE�J-4��(H,I�Ѣ�Z��h��#cFDH�cDH`�dA�""ъM�)�%1�5�h�4I�*��&L�ъ��$�ʌh�F#�,a�l�(Ѩ�KF�XRJ!0TX�X�Ѣ�aM���ƌ((M��l&(�*(�H���Ƅ��lQ��+2���F�@Y4d�Q��B�4bKI�X���B"�"#bɱQ3AB��(�;��w���O�O�Q&�{2���=�nv���?Nt���S��8��Ŵa�����C��N˝=lM,و��z�#���Ｍ�V���9ӟ�%c�S��!C㤞� }��&�_�-�,0QI^ ��Q���Q�s6�v�h���!��K��C�rKv�<��Jo��ʦ����ʞ�/ .�����{����X>�`W%b�2:8	V_N�f#zm�	�%Q�5	U< �@��{��ޫ�H,v�ByVՈq��,�P}'�{�֩���T���+�W#/�UbGLI<&M =\���k0դ��;R ���V=�V��c�����4B�{k�U�V����!�=7�=NxKxe��!d�����Æ٧V{�sQ�F�w���~r�֮^�|�˯M��M�{������d��W%����A��d]*y&�!FWk�8Բ��Y��P.7V����
4�:g�@�G��"9ٚ��E�\'n}��2o�T�\�W�*�;�~'�G叺����4�fOm�Z���paVՆ��#��P�Q3����̨��a���';�����.�j@�y<��^ڌ0�O�f 8��![�����_: ����q/'Q�~uؽ�t��i�#S�ݢ�N.�Ooe��ĭ�B���<��V�G�����j6 �i#�����-=]g��������f���%�<z��j��9��"y�p��|���qV�� B�i.� %0K��7_��{����kA�غ���C����g����"��=Ə)�ȧ:��l�j��6�F%Og�vp�u�'�$k��6N�_q1�j���U��}��}";ԝ�+��`������%��"��fx��V�_
��Y\#�����1G��-1��@S�vˏ�KYe�����s3e@n�)��g��UFt���a�+W��Ҩ�|%4��q�ng�ŅJ��;�M�m�t��Ʊ���kZp�����p�,�Mĩ*zfx�k�a�>zsޓc�ذv����/�Й��u>�}�}9��.F߱���`=⣲�ߖd�t���S�8��x�/i�᣼]2�����Jq.fUo*���QO�;��,ڔ����.��X�N_�����@��%P F��2v�U+H��x�ܦ0Ej#O��(��C|���ޥ=Od҄���u+d2`Y4/��=`�ڈ;���|8s�ŋ��,5z����""�e���S���K�^g5";�@QӃȿ��4��u��U�<��=�%��˩���H�
G:����pVin;W�OVF0"�E]I�iK3mӰ)��r}�2�e��^��w#\4��ޯ���{�ҳ]���8R�����X�^s�w�{�-���^�ng��{�+��u���KO{�9�qr�I7\/ۆ�A������|4'D;˩����߃l����F�3�(6\x�%���S/�8��\j7��̕3�Y�r+6�1���(n����������P"����42ԏ̇R�D��� Z��/1��*���7k-v��R�l�f��Z�V+^gH%ns��@}��"C�U�{���w���d����� R-x\������b��'��Q����(�˽[<��{�1d�%��7��o�w���}�+��D縼>Rλ�G������Q�ҭ[m�;�v�N�U1m�����M�g2r-H��"h(��x:q;3����Vx
�nc�q�zԚ3�w�0�����dk��>ޛ�V�O�ݑ���W�"pV�>K��\�ht�65nw�oz���CԀP<�"��<��\�g�#q��kl�`�I:]#�eѬ���M䵗�:�_y�>b���\,,��(N����]4�2���;���#*�ߗ�9q��5�L�%�*ν>iG����K�_z{��V+D��Z(���7�l����7�|�1e���x^�1!����:�\&�ŷ|�>��ƌ|�9���{��ϴ2:��|t�����Z�C���r켌w��������Jü[,�q�M��(�'�T$j]�j�Q�����Eyk�vny��+F�:�rU�� < �6����Q�of�u�x��A�' _Z�w*�*�ܾ9���z�_q�0/�I�#Wq#sWh��4�|{���B���o��|g@@� [�N��m�``���?M���V�p�N'��y�V�F�L�L�z�'M���F9�t0Y�(��]�v���2������m��v���7�_|�+Q�'U�\�/D�8:�@v��#	��Bi��ެw��yZM���Q~�1��Q׽P��S��
�"q�q6��hF����N$'27�3�c'ћJ�N����F��"�zyG��1pU�MFt(د[�fy��3�|�h����Y�G�>;ؓ9���H��;�"�ל���}k;�'��:�@�%���m�����B�vJ
�s5�6ϕ������n.
��'k�3���ɶZ-tN9^��0~�\J�Jxf�2;7�@H}*��r����
C��^}�4�{v��m(�~��8�9���X9с;6��O2�ful�퉠�H���)��?v5x\E�7�(W�~뮶�b~��4�9�G����N���%>�e�ܗ�s3\�
�
57hq���KF胗�p[z�]�L	�hC��t���
_f��ٝ��r�{[���W`κ�� ��B'��zZ����g�F�	��!]�Į#G�� {O�,�x�*89=��� ��m�@X�5uczz��=��Ч&r2ӟ(�v^��Wf4k�k�bU�d��2�9(GD)���y�`D�Fߕ8�5����i�Z�_����C�|V+A��%�ѥ�U)�C6��lr��w���6�7*f�íl'Wc��7�Ni�K��z�:���@�\%�Dm{�b�0�e�uN6�����\��ў�9��]p���Y��f8W$�@�O	M*��Z7�~��nX2��^{�P6tXP�J�	��c���a磰қ�Q#D%#�Q�B��:jy�Cꦗ�gt�t��~Ӝ�a腓z���j�*n8�D�S��4m���D19�AծQȠ�H[�~�L�9.�S���"[f�)��
��~j<�ke�3:G��mh�ꓙ7� r:"�OaC�i�`1ٽ�_�K�]�l+�SB.����&$��̶ژP���Z��1�xׂ��Hw��4_��{�������'��B�r�{x#�V��6��ΰ/Tr�m�8'˾C9�M�������L��ٛ1w�F�j^�%+�o٥ﴮ�	�]��yq��=�T"F��ɞt|�<�+�y���7����s>g��VŮ����4�"���}ta�z��v��{�}h�M�ӝ�*Tu���6g& �xY�
��DN܃�KHȰ)S�7!Ff�šXƆۺ]}4�C9g���ˈuD7N"�5�F}p��E]��,��^Wg-k�OJ��r�xs�N�¶Z�	���N�A��:rm)��=R"��v�����m�B�'�:_f�js���	��ٳ# d�rFe�'|�1�ڦ+7��}��L{(tZe{�W�Z���h���]Q�c��xe3��a����kT�(�:��d�]�v�t)��}x��5����b�}'���@S�4�6%>Cڥa�c���-�����C�WtهW/1qS�FE�	^��ai�
��]�:a�>~LS\���Aj��I���DzyѻY /mk��N{g��z�3���=9r F����&v�\T���VU���V�������^̣�j kZL8X6[����A�_������ߑ�а��R@S�3�MxK��	�ܞ�]<jn�M�z6�#5 �Fo�����r~��v�+IF=��@v���o���`�xDۍ
�bJ�W�uu��Zh�H�<ĵ�R˷r����<:�bEOO��ͮ\B$.ҷ,\I�!솧Z�J�N�v�N��{�7��4������8;���p=�Uؗaz\]�:�w7�&˾�]^#��ڊ���R�ɤ!uJ����d�K�Fm���x���xi'qn�;0��������e�_�<7����*�����^9kz�ԧ']G�C6�wu����`�(�2�u@�cQ۪��{]�W����1�0,L�MLs���w:G@c"���5�I�g�D
� c}��O�x\����u�Ŵ��*.�*�r��|o��e�v��x��D��+�(�WuM*72Gt(���7��a���Q������$㳃;�DhC�O��V��J���*q�
�fo��_M��!q�Pq]野sq:�Ve�Da�^[�I3~�q@���lq�p�x���P���mإٽ�]��eZu
�ʥ�Up�wd֏1��W�����%�]=�~�i�+�ضסXK�1��4������0��Q��tm�_y�;�a6s������;���.�y<U�$s�H���jP�+�,8�&/>0��P�c�W���ɹ��U\��p��|.�tc��hT�w`jg��Qsɣ�jąC�h�UpB������������ӅG�x�A�H����e���I�6r�V�D�ͽ���̰r��mNj�:��0Ύ���1��Y��CjV>��=��k���*b�w�w���� 0兛I�']�D�W#)���p�g$K��m5`�J��͠9R�ԫOT�ݡ��x{�No��,�}Y�۾��E��2��ɟoKW]�kox"�ύ��;��=�Fn<Mu�����6����*�@Y(=�	�ޭ^�g��s�-[^�~�^�v��� Ad�Ϸ�{�FΩ-�������{��W�s���`�f ��(M2�/�F0�2��;g��S��.��Ӻ+�Z�y��!��Ѥ4SG�x�4���?Y��e�y������E�W��>����]Y�p�=�rW�o���w"TNZv&�KJ���s`�}'Ҕ���QĥB�������G�Xg�����!A����xW��x� 7���\ G�S��xG�	�j��1ۃ�z;�]�Vؠo��n�5�ݙ�=v+�̕>!�䩀A�����.�QW�@)���ҳW`��`Eg��C�j�`��1�d�J��\N8h�;M����'�)�ݨ�s6rN S:�3~u��z+�+�`�c����D��C�� �g��q.j��j댕5y�7��h�����,��n/m{N30����}��E}�<��|���YԲɽ��Dq�t*)��{-R�e8dzr�({���&�m���c��"Z���)�μ�s#�'�hx���z��%���,�E�#`�p�t�+���U�A����T��	�������#�rBZ����-�6a.�����%�?{� x{yZ58�'����Ux�ת�\>�Ī\��ý����6B�r���譠��1B�ή��v�N��ݬ��Z�`�롖��4|ص]�j�
�0o��_�`�~9�0�ہa���Um�q}�<�����]x�w�k�l�
���{k>�a!\h�}1"cc��eec��Ȝ~����Y:iN���_:�Ό	ٷ�|S̳�[3�~�&!�ަK�v��V����e�y��T�3�(8��/�[�C��J������֞��=:dW!y�Y�F�>�7���d���,���^��;6��H�J�eLE��9�D�Fߕ8�'GD����r�RV9�o#.�Ucӱ�>-4���t��^�Q􁢏�ۈ��Pw�EQ1���ϖO-e��B�2�Ut���w�	Q�%:P+�S�A�|6�+�K^������+��Ӽbq'*4'�����>�e�d�8�%�}�Mg�e��Qt��r[����u�=�S��XQ^mC����}o*w��[a�-y�z-���KܴN�`K�L�d�3�NX׭"7����i�"������ʙ�4'���,#��
+o ��Լ��ų���w3�'G%/
/J�Ͼի���m�Z�(�1&���4wP��zL��=z����h�'=��n�!�e���n�K(�	��8���<
������� b�m_
�N���.��R��[�a.����/�9�L�!���.�#"����Ƙ^�~����>��Gf갩�p�Z�y�Cnr���NX��t���t֎}`���0=��&�ө�s�5W�;����w���_����������lإ֤��]�}kҵѥ�G�ޅS�cf��HvoA���F^�=Z�ߜ��qb�ۣ��M����'�G)UU�ڼ�aV�Y���������H�Xâc]�Ma}(w��
���]��{�v�b}���M{��+p��u����)��1�H�#�.u��w�l���b�*�Kȼ�tp�Я�G�,�;k�{�ى�"�FW���o&`��z�+�.%�ֶ�P���:,��bz|R4�����9S�=ۡWI���a-dc̭�Fa�t!�>u��}�g�B#���[í�������͜��M�y4Y9.��U*N���\�l��=��N�k�n�H����{\�ԥ_���C+[K��ƪ��n͸�j��<r�b�Q3Z&Hy��ບ)�q���H$7tn��q�zG)�5��r]��$Y�9{���A�p�M�|P����yu-+6����xZn��|-;��Q}��Zk91u%�<*�8m�/�	�/�wyumB!�V���l,�ky��bQn;�����Y�9b��Dr��x���$���7� A�0U޻��cb�o�k���sX���N�������3�̮�g�w1־iX����J=6���Y����d�w5�BSh�$^A�_iy��r�f�
Z�Nޣ)���wW�E-�o*9����5�-kYTxbZ{w�Z�E�큼}�sG��\� XN4V�|VM�jS����P��ƞ�f���G
��-د,ru�۸���^LX[���)��Â��/��љƖح��	u�FT�se��!�qV�8K��0QK<���C`{`\̽�J#N����*���fj^Z���ֵҲ��D�X��{��YW��+��H�D����\��˓�OP�&�m����EM��o.��ۺ�i�ygt�)�ѓ⸬E�Z�!Œ&soj��$�	OWA�@��
k75������w��M3�-Ù��6t
�u6E\���^2򬋤5����#+!�;
j]m��*��TL����R��u^��r�i�{�{l�ǯ�1��VOq��eQ��o����}��:��]�ˉ�mR�1A�v��lůgIʄ�jhrh���%#�����]��ó#"кf��z��18̏��aKq�M�,bU�oY/��$�U���s��[��5.����&J|��C�˖��7fd������oy�~�Ju�R�su��8{"P�c��oܵõ�b�&���J_;us���m@�GP���]U;2�jL�)R(#��Gt=�7�D�Tr�b�.��wDn9�\�L�jض���n�xA�����}Ƒ���1����kN�1�}噛�?B�5ï2�)�����`�w5����g=��aA|��`�c�6i~��ZY;�B��z�|��j�C����wu�BQ�J �Z力;"v����N�`��;{��c�㬔с]دێNw�	9�q��0G�W�l��9���9���՗��}��z��k�W5�9�},N��������� ��F�oh{C���*+�s�S�2���ɭu=h��N鱬��k�L���V`�X|��J�Zz�R;6�Z��G:�3�.�p��:�`Z�D��Ǖ�V9��$-qti6�V8��E۹�2u��w]������C�S)��ЈP��S����[�o!/��N�,�����F,u��Wj0�K��I�@�
Vd��KF�E:�w���|c�Bw�^�%��'�C�H �B�Q�"	 �ld"Ѵh��t+!$X�Aaݸb����1���F36(�j)5
DS1h����`��lQ@ZH��rۛQi�&���-;�QT�Gu����F�7UsE�,A��cv\�DIF��r�b!7wDbƒ��Dh,N�]"�k&9\�0-�ݮm&���仹b.](4Nn\��e˅ݴ�Q�]�F��3�n4�l�+�đ��4�&,	DX��˻�\�	sr�L�!;��m\,s[���5�]"ь���X˻t��Q�sC"�L�%ݢ��\���!7:�9�,h���������$�&��7읢�d��Iu��:���r��(s��D��>`-��՚���9��f�x�j��$��w�� )n�sE8��8~����jw��eu�q�D����uƐ\�{mA.*kU��&�-�������
|��S{ܲ�w3��,N��ηrl�J;'Vo<���`��˲W=���0�coPe=�W�i��]�Y�̪p1q��p���tԧ0�#2w[a�5�����O�����a:�r�㪴��wXz����mN�������Zʄ��ܱ��c7��u��O����z�;޻J�VMlɸD/r�#f��}Wk���)7�Z��^r�x_j����l7�ފe�UJ>�.�9�J�}�!_
��\rA1,3���{s�n6�9}��z�ےS����@ծ�DƲ�V	���ښ�+s�gi�:��e.tBo��žSa��G�L�ǵ�mF��+_V���b�+�V;�7^$�R�qIu.�p��f� N�~�@�<���y�Z�"����2|6��/�����n�z�#�a7�JE�e�Z6�k� \X/�ݒ�a��n���V)���v�3]N��3��1��s�Yxs��s�@,��*�\ނU��K�?L#mY��4�ݹJ�1�9��of����_}U@��I�k�[W�^�|Eva����ev�W��v���F����n7�+8�+������X�I o��[��^Z�V�Of�<��}�9)��8���UsK-M�uu��^n�U���Fb>�{+"�D��v��RCgC��T�/���^o �s�^,��*�C�k,�b�6�
����~1\�Q�^�z�1	��	�����]wq���&�'/���E�y�{�����zm�W�7�7H��_^hkQƶ��=��۝=�zk��TE���LT�"��B�j�X�h$�oP���v�̌��f��_Xjݭ�U���ar T����ҬM�kf�t('Td"��m>މ�^�v�m��%c,�v��>���N��;U����kf�i{NT�_s���k�<��-؍�e{�	�$���3Uو�6H���k�ܚw��o"��M[�WI9,�j3[�2�*�"�ܮ�6FR���R@:0�3�|�i���	�a{�7�=��v�Q�E �ޱ��A1V�����Қ�^n��7t�\��X��
��]��Q67+��H�Tn��x��Ѫ�{M*ݺF��������7��1x����IL'����ov�9�)�$7Pϗ���S4��b��.�F��h8�}p����e&����=�>m��\��^�3su�hQ�������?Gs�Os,Bt;6���M�;�n�M�y��EK�uw�R�9J�=GfF������Gز�\"�G�q[�����ȋ���ױlx�6�q�(.�+���_S��H�0�G��{��~��9�3��Oy�%6#H�X_F
�#�F-1��<�����^���1^��|/��O�$���n��լ:O
�NsG<ʻ�,��Iwi�^�9
�2�K�����c�q:gU��[������>O2�����kq���'6:���]Ӆ���O8����ª�.S����z�i͙Q���Jzǌ�'�^�G3��-�wQ;�R�>�C��z��G�b����[S�Ϧ�E^E-�0z�,�Oewy�ZzW+<1$M,�+\�ӧ�}�ONu���o���
P���F>ͭ����T+{�@Rg%�u	V_ZfW6�d�9��&0olL��;���GᏮ�^��-+{݅{�ޔ�p��p�t�캴���F�uN}�k�x��z���!xh��b bY]f㸉WQ:��|E �d�ܔ3N]S�t����g2�vr�9���m.�|��}��=��}B'�=�U>N7�Xх�x����t��[�ǲS���o,aki�r���.�>��p����1
���*ȟ��S�������E�b����W휄W�\4W^��diR��d��(G'1ق�92�u·ژ��p�S*Z�/:tJ:�N�_bH��T&7��$l�lP�O�-��ES�
�%�y�f'Ղ3��se�u�y�]i� mT�:��>�����E-y~�ݛG.k;gp��E����jkۣ��/��LBV��@����#��xTjb뫿tG�c�8>�.�F�'���p7_;tx�XȨ�]��k7���yށ�����>��v��Չ%U�c�lkQ6�,w;]�|!}���z�h�|�e��.a����{$b����`T2����5�F<8qS��S��7vk�9���Y���U��Z���D�qk�k��6��1�$o��Oc۔�A�Ŋ�s:�V��O-�a���-�7��M�Y2?x ��Ε��қ������[γ����*vۭ�.j(X��yq�xmr�����E[�y�9�8u_��儘�a�:��u�G,y=��p�:#���z�-�V�o�qnOֶ�P��|~����\Jp3�_vu�n��1ok6��;��Y�	WP�WXE ��CD��{z�bbE��t�v��z��i�3y�y���q��G����=�����{�s����cVGs���1������|���뭗s(t]��+�<�'[��7}X'S	���l�w�7�����{`*�W�du�q����k{��Vr�|�x�O3R�_����o��ko������ v�C��ݒE������{��e:.�ܾ�;��<�GtG���,fj! �5C=�X�n4v_t�ūspϗ�UP�/��=1�8��su�<�΄Q�xyhY�R��^nf��!|���AOAS7 e�)����>�M�:k��ok�yL�T�y��4�V�z{�J�H�/�U�QӛH�%W+*#��=��;��ȃ��YS�Ҕ��7�˺�X�cp_k6�!9*�¹'�C��d���)l_7]y�BƷ{����\�U+��D�#���-y�����{_,Oz�n�,�`�<�I/��<���­��SZGm@�Co���_�0m
Uu�m5WF���s_oBЗ:M�5�lcPF��T]ɂ���J�ʝZz���;�T6�6����Y[�J��'[c]�5��LTN1�wg2(���Iy^>3��6���Ȑ��k�)���j����G�b"�.�f�;�"��Vj5��#������a�,�9ΎW	��&EMIh�j �{�r����W���`k�D��*ޚY��>�dZ��3�Uv�{�qbn�l_�|��=�5�/%��+Khqϯӳn�l���%_��v�q�`�MB c;A�|��z�*����S~^�֛�77R�R厙zJ8�ڽ	ô\KF�q��v�!���^->�}�~kUe)���@���fWs�a��)����_��c�;z+�w,��V��آwCR�;or^���b;�Ms�[3!�����+_8@nh��X��6�����yZЖӱotf�|�B�oʣ��N��t;��μ���*n9���pR?Zi� �?#�u[\���5ed�a<��U�����dT�4�"�ka��i��W;�I�p�� �fe�*�{{)�莩� C�1�N�9٫��&ͣ~ӣ�[N�O.q������nW.Y���g����}�+���a˳w�.����BS��/�mcv֡�f��8Ce��,��U��$���>�%�Jy�+=V���h��[�o2���eIn�����Y1]Z:nX�k1¢� ��!$�V�5���a�.��ۦ��(òW%5J��2Fe|#['��Ö�g�ڦ��Ь+P��k����{�XmN�oh5��}�z��a�4��ѧ�X�=������A�\���]N�N�Ej�:�}W;u��/���2�I�b�b�bk���vn��Q
��1��[a�؍ s�}0b8b܌�i�`'�[8�Nm��j8u�CUczgp�������O��&�8�#7�v�Ct�ݐ[�Q<��M�i-��8g*`�,�+��7�QȄ��S�i�����������9g�5od{�����Z����C}ꔹ��z�\a�UX��B�xz�'��3�����jÔ{7�j�'�V�u���*�X��>�,�v|����\�7�N�d�~�da�����U-��'�ƺs���e`]g3#HVD>ө�q��I1Zī�����M��M��aUs)��o7��c�]��aX���;=�:bǲ.��c2����C��z�n�5n���h��ᮞ�o��2�OgR�a,DcYP�i�7��,>�����mg� �nj��fW[��c)�%�;Ά��o��=�W���b��z��@�4wO)�Ѥ����u�5Z����0�w^��(�K�����,�v��r.�*v�\��YX����,T�5/���eBN��kl=��<����n�rFe,Uոp��ŕO�o�؝�o�=�Jå�>���/��c5���AU��,�ꒇs�7Y/��G7�S�0;�Frٿ�d��3���ػ�.�'|u��Srgj��Na��/`���(7�-Kv�m�ta�=��
��AVw���qzp�X�n�gf�k�p�	kwwh��`�}c2��w|sGI���Ot�t,�wt?#e����n�	��R[�I����7�X�Z��;�I��	�=_����|> aq��y��kOGؔ�*HUR���a��d�+��}��aV���A����&����{{��B�s͊nܐ��t��#M+]R�N&�ݮ�(��q;s�����Ba.4@�;r�;N
n,P���|4�ql��D�����;���9G��G;;]�I+t[c]�ſzZ��xؓ���S2�-4x���8V��<{cVQ�j����Zâ-�:���2����w\$eh��B1�E�1��[��YFs�p꾪yi1�c����8�u�������-��!��q~�%�Ғ᠉��]@�*5䵫���6���I7�9f�7���<��qw��a�ʺ�H>Z�cdnŨ=+�wՅ,i}
_!Қ}���N���eu����V#T��)�vx*���O��w��FR��b����i����Y�5���nXS�Q�(F��h�8�Q5�óE���.�<U�6 	���WN�gqT�zb9/l��5^�����6��<:y�4ZZ�6�t�����i%w]u�s-�/d�s�	��ـ��Տ;C�^k�)��i����\�u ����w}���h~����ޗ��C�?z$�-Hr>[IX�n��co����a�5F�m{(=-������� n�}ڮOq{#�L�.�,���pa��v4k<|�uc3��Ӿ�R�k���ﻠ�i�Nլ�)v��	
j���pC�֫H^5�p�S)[��|�@�!!^���~���Ɋ�[��ܲ�T���Y��m؇z�݂��K�8T�������{0�6���װ㭇�k*��g���W�,�i8};�IX~�nHUN���1��S�j�o�@��o6��Q��z�Γ}lc�6(7n�:���i��V��T�a����ܣ�o(��u�IUr��m�|r��U]���p�pC;�]�{"����W���[U�����4��ǝ(�	�o�+���.�WЩ�|#H	V�d��GP}6���G&{�T���/j�N8�����4)�pb�"�Y�f�Z�Bӷ�D���l9z�ދ��G���B��\A�4}b5+�A�&˜�_���5��vIU�̽ǉ�cU��n���;��jlAw��V���U��q�бR¤���	�Qo��%�Q�֬�-���S:�:��t�)L�����p�����8-�F���'�0�9R��Xf�M��N��י׿0��]w��#!{D�ѩK(ƺ���؋c7xT=**N{ہ�Ɩ�tt���	�᥷��ա������^�����*ď�@T��g��;���Ն}��v,��-&M
��0�݃��a��(D�v�7"��w/�i�]��ś�ac�:�,�eL	M����RP�Rtw�����a�*���g��{7j{�Y#��s`�{y�!�|;��*�냲�R�kc�'����+h&�1��ϑ���X>=����;OZ����ʴ��͉����>D띹��X�!�qF��Ae�X��+K �1�ε��L{�{����j�s�b|i�n�uq8�9�x,��SVo������ۃW5x�މ�V ��(��F�؛�kӏ�m�M����Wfp���/z:��4�&�,�(�Q�۷b�a���Ɩo�e�Ѹ��1}9����Wt�%� F�k.����ˊ�.�^�Z�m��[%]4g��l������.��U����ιV���>=�.qn�ON���)D��9o��k�S�G�yd�(M��<���7^�.�p�qޡ�#&?Uxd��m�:�o���h�<j�;3z�'�p��u�"���ݮ&>K�y<ݥgt�'���i���Ve��+\nB�x �R}\`KF��&���h����d��x�bn�W�'����K��e��溸8���K3���n�D�Xs���M��[>���
�@������;:=�F+�3}���8xǵ�Y�Ч�p.[f�.mr|�YZ0ʾ��1�-�9��[�u͓q��֨���`>��IM|DE�ʇ�>�h�/{��؆z�;2��:vL�4F�p�{Y3��[�$�>���q���F];�s^֬�Q��g��ӧm�ȴb��4A	{�8.$��D�j��
�O8��<�G�3�S�F���3�,jc��q�7�
��J�͛���|{�'�Zx�%��]�R�����R�Ce��[kn2.Dh��v��9o;�m���a�}���@��^���X����=]GwXʖ��*ޗ�	�u�6XFg�<�u����O4DO��/kF����[��x�lL�*�P`�wk�������������(|Y�7rcZ�Z>I�凃Do�(���LM��v��/ͻ����Jp�D{�=���+���_f��R'q�n^b��
,'xę��7�.�ٚD�S��o/�N�wSɵ8�V�A\�ӯI�+Ķ�m��Bޱ9u��Z�/���W�,lb�scd�t���r�:�
˗d��QI�M#�e�ssd3��d����#˅T�����F.����9����r�����ѵ��d�A&$5s]6�r�+sA6���$�����m�nU��;��r�Q�!J61d��,lE3d���ӎ�\�j-3���س�Q����#FŨ�gw1�lc��cb�cRQ�\���s`�4`�nRX��c6�6�Ŝ�,mstŹsr�6�L�06�Hk��b�w��y���??߿߮����;�Q��)h!��v��6/6����[��]x��jׄAA���Œ�ڽ���f�:K���������
�����Y~J5Z�S�BWg���%��F��.:�>Fia�/�ec�܌xŕ��T�z�}O{<�p�ee����V:�ډRp�)J�}h�xf�]a�'q	�]��)���7��#ʙ����f��i%2���+o{����@�](>��8�%
�\�am�����
����^=h��}���o<ke��3��K�!ȭ��e����=bŋq��vb�������D�{�Np�M�r�oַ�N�+{#�zMZ�T��uȸݽ�g6s}��i`쯒���Y�����#�+��G9��Ux2��ǋh�wsJ��J��vc4��N�n�m�+ܣG�]�7�qUiV�qwάC�糲�u�V�q��x�4S*[�z�U�$�Y�GV؅��^�b@��L-�vl"M+s��{�Co=z��֊�99o����f�k5p��,��ϳ]�۝u��.缘��w���Q��̆�� �BX�M�_vc<=�`�&��%qL��g�UAӇZF����e��gn��j�Љ��j�y��O8d�XZ�Vkx��Y���Vg9	����2g���#�~yrm��o�����vl#˝�C���x��r[���2N�Gl�������#M	Z�_]`ŕ��
h����[�+�ZhF��z��&ƻ�,��2�xA}�[9���,]�����O�����rzyw1�o/���Þ�@�XC���DUV��Z]��*��X���O�o��:��j��Oo�k�xUjs��2�Ʊj'Y��}|����%�����CO#��,�:�lX�;��s�绎wD�O
��W�3���>3Kd{�;t!�>��#��8��|��U\ŉOWe�[��:��ޚ�H!�m�������em���D��b�a�C��͝��ֹ�Sz^e(����v�/u;]]�١��z�g�'���E��wb��{������!٘�z&���%�+V_���<��u��_TO,�*A�u/z�y�8"5��]�r�
�*�f��x��Z��.�	]bP��w�=�ɝeD���}F
uZy�����,r�w� /�ԣW~�&�zfkN��Rwk�vR������Wl�y�K$�����J':co�N�t-����=�
�A�Td�f�+etN���g]�Q�X���+��l�v�y~���r��~��EtB�L+��g47���J䊺�)<��5����
e��xdvE�
��)��\�N^��ͯN�ךYR�i��K����5ޤ����U��D]����Uq�=��r�	0��F��p��f�M(w1��mc�O����%9[��̄���.O���}������E-y~���;�6woM��c���;���}�;P��lSv䀪�t��#MzV����iV>�8�ν��7�oBKj���nX�~S���X�v莗ǪL\N>
u���⺩�ObˮyDc�9���0����`)�!�`롮z���W�ϻVu��"��{=���=�utW�uk��������� ������ �i�Ff����b�w��0��@��~꧉U���<�����mbE�0��������J0�-�y<����<�Os&Xab�5�h��Ww[�a=�j��}�x'N��K��8�s�2��H&�i�{�ӛ�ҭ�[+�n��+ޢ�|/CRi��65��!�7ĭ\2��ں��VA�M����u'�!���oz��/�_��,���?u����!��j�#���D�Ѕ-���X�-�?w�3�{W��yZ[C�_�nKi�}Uy<���Zk5]��X��\ŉM>���߂y�cY]F;�үT�Σ�����r����ӹ�b����e>��*�st�{/Vtް����虌���=|�e��*�./JdT�4�"������0�coU4�L��h�s�w0<���s����=��N�r�*R5/�����m�5��Mo�T9��+e^>D���Q}ۜm-�6:���P7D�]�o,�k+n��7�9���Þ��z���c4�s���V�2�*�� }ϫ���J �}�S�;�s��%���ýz�dpx�2䪩G��� n�v��H�kC�M�ѧ]�/�����<�W�/��s�x7����u`q�V�Z���u�	�d*��n�wn!X�m�tV}n��esxݲR|�����D4����Ӎ��=�=�%���1D�wJ���8p�{w�⎋G@w���E]�G�K<���h��=��s���N��
�6�V s�.���]4>��,��������M{r�']��ΈM�;��;
l2P�WcW�,w�̭�-p�����c�E;�Ŕ7^+�H���↉	wd9�-@�*co�퉶F
E�`A|4�뷜���)�� �L�4��86�}a�}���_s
���in�X���u��3���9Z�ߛ�Q�evb��Gԏ�}r>�^r�;��_yt��o��N�G�x'�s�'5-��R��1�^��������9�^K�V��*o�L��8%wL�f���N;���z�0Gy�.�p��P�.%3h����彺���n3��~�\E ��1�d�^�\�Soz��:�V���C0���c��=�������R�5�%���[Qᶖ=}Y��J>�wCU��3]����R���!�5=�U>N�u�9�ג4�d^��>GU(��!�_�Ba�o��[���%�)�;��ZZ~*{��N��^��2�2��6˭��U;���z�*�k���FKN�j�u�\�V!��99YiTɻ˯&o��ou�75S�Nr5�"���]X��2�}��SJЁai�ڌ�	�N�A�����.Y���g�@샐~��=�fPu!÷gVE�N·�e'���/��l�`Fܳ��Nl�-w��}��zP�+ 1�z97W�o��%��+}��G�t�eHUR�N���is&�T'����Cb�,j�-�;6I����<)xe��<��/j�6�A�Ä��GT}�Ȅ��-̿Btf�<��P$.~wq�/�jSӝЂ;���y�a�~OH�c���}��VJ��5��B]��w��i8��±�}w���ճ������ޮБO�u�Yڎ�u�Q�;����6�i�X_F
�#�1mC���/����IQ��k���u��RǶ5ex�cz��Zâ��N��y�uT��
4�
u�ݫ�j���;�љ�o���0�t2Ϋꥱ��Z�����]�Qz�K�;@\�����	.�_>���Տ`�>�ݺ����SKyH�U���,�S(Wj�HJ�gc�A^��0�G">ٸ2�`^�_ѽ���tBc���s>�����v��'(k�{��3f;j�k��l'I�-�i���_6{�\�"եsM�G�u���8�B��S:�4�ӓ�o&z�.-;�|�%������R/%��+KG]D�)�A��9n]�YP�e�\���<�m�z��t��E�k����q�D�@�4}�\]s�f�o�?^���P�]~*&��S�,�j�����zT��i�!b{Ovv��#w�R^�N�-���j�0���ڬ�q�*���tZ���y���ʈ�'D��5<Ϫ{��k(�I�a������9%=QGe\��
M���3��S�a!^���XF�����h��6<�i�Vg�u�m����^�O�!B5>���7V��Q�v�D��l�9��D�^c���<� �ۜ4˒���\`h��t��X��)k�4�'ا)����\���wE�-
¾�BT�tʝ�P���y8����JW�6�+-
't�^B�NWߥ�仚�+9�-k���aK��9S�ް�)~���O�������84��]1��ӷik��l!��>Y�/w{ ��֝��Q;��25m9���j��v{O�||6Ii�b��Үѹʮ�Nu��k����\h�Ið�j,cqb�ۡ��ir�QK(�p��T㮄�fX�yGVs�`$��*-����Fs��9z�u+b����� �+=K0�X�Ƭ�����:�w<�#iLn�@�[����O� ���\Ϭ�R\����ҞË��E�=g��MsټN �v���'��_�m�����ih�2��8��gg� ����k�i��ۧ��z�:�B�)���[��n���D��|�mAoU[�q����\l�����k���}�������3�Si{�CZnC۝G�qn��&��W(�j�Jr�`�O�ш_.n���zy��RY��Wy�B�=�:�0��c9�J��EK�!ȭ��e��a������Vf�y��spc2��U��e�_v����?�R{�[��\���Rű��K�c;�a[塳�7�����]�I���ar^�7�mEw3���R�?n
O国�5��>�x�"�9�f�rW��/!Z���Qq7�+��9�a�VM�`#�����F�e�tQB�e���K�_Oj�#	�Mǌ=�z(J����X�;���1�����Տ�v���ìn��p��*�#�$.�;�|wDPG�_�O��������Ym�]��i��V�ᐽ���զ�^h���sJ�엞���UҰ!޽��`�s���)���.w�)][w�鮭v�:N+�q}�}X���{��ywZ+B�}¾IdQV�+��x������]ռ��<�U1��ok��[�F'C���Gɾ�p�ǹ�svr0ñ�6�]�g!���zapڿ	[�i<�1en�W䑭�y�UM��c�k��'+{��p�jkE��n���#m��^��Ǯ��R�6�|s��{����<����m���a�2I�#���Z]��Ix����2�Zv��!�#g�-g(�oR���oi�_��7w+X���"Q���'o�u�^g'�WwyF1e�ު[|�K���p�y���'�YS�Y�n�%u�~!�}��D�:�Ⲽ��a�ݐ^x�#�*�;n<p2��5�e�=f���^�N=�UeٰT�=]�}t>�a���.��Fa�0nۃ�=�|*0U�UͼI�΢�C9޹@pZ�sL��ݨ �.����[ճ�!N�������*�Gk>��>��!غ0u>bħ���כ3N1w�L�}�i�U��Zܧ~7�]�N��:�A���8������y��=�;�7j�'8ru��<��N+���mutGB�:�K�Hr[-nZ��[��9����7*w�w���}-5+�M��Yƫe�σ�ӎ	|;3�м�6�I��gB7W��~]�#O��Oag6�ڬn�m�]�ӣ8'&�*�n�={5� t�SP	�R�Z��	;�o��X�/:p��v#n^wI���l_s�{9M8�V9�"3EC���{$J]�![��7�㝪F6��\H�RS���N$�췵}�K�}	
��\-�vl"�JÜ���tD�u�1�'%Q���1,�������G-��w��}��5S�OB�0[D�yr��ͽ�5k�b�v��7nT]tBᕲ���)�>T�8^J�ct��]��er�.
/s8�1����ͫY=]����-;����Kofi��Qk���.z�w�2�����T�ᱛk��Qi�s.o*�k���)��z�D5 ̶����R��ȹ�r�4p����+�W���խ���z�d���e�M�/�����8Н� o#��x���@��B7�1�ܫ��������x����OfWW`�{ͰtVF��] ��c-4EK�橽���{ay�,�l=�: ҫ�z�B���9��/eE*ɥ���N�w.�	�x(qG�7�X�A���TH�f�Ů�Vw^�7�eaT��r�\CǱJ��}�q\U�p2�
���g�u踜����!���c:��f���x)�1��lΫ�G6KǀG���tb�^]9�:o��� Q[�tN-MD��t�~�L�"K���+���9A�P�/�`]s9��A�%5����+�S���+bS}E̘r��Vs����J�:7q&5#�,��RA_Fk�3�\�j�sw��v+�\�huժpc|�ދ	���	��>��2*]�Aw6]�7�O���Y��F;3//�=�i��r8 GƠ�c+"���h���r�9�y����Em�IE���Li:tv3��R�ݣ��n|������7�ޙ'X��ǨZ�F��D�Iq7F���W����E��4R�{��˧�{�+�%@�P	d�������Lu��
妶�Ò�8�c:����|+���@+:6���ܐ�f&��x-�!�Բ�ւ�F=��.;H}t;7�/�������9Ƿ�CA�]:E��n?n[�ʊZk2rYO*�.J�s[S�z����O�G�7q�A&����d�ki�`'�:�0�FN�y'k�3�1�3�w�!��\�b���m��hP�J�}�u���]�l�@[�o_$\���x�*sՒ����7&"�!լ��5'k�	��]�a�L��p-t�?��V��(�dv!���Ĳ�#r�}�pd8 \�
�	h�&�<�p�fjRq�#Ҕ����"��Χn�����kj�~�0�y(.]S�h������M=�%����|�7=ɟuŝ��I�g�T�f^� �5�����ɉ��ab��5LB�fq�u%��;/IZ��eeY�*��Q��[���{u���3��������k���}`�MS;E���SV��4�<���]��`X0y��U�G�����5��� �ı��7�k�Z�h�D\o�iV��V����+БgrY�*>��6:st5�b���v�pcfm%��6̎�n���;wx�ٚs��f0e�h�ym��4Y�J@hֽ�
ч�<�\l�t�˻�����Y�XR50�eX1��^���<<�'���	�(�u�n��*^ɥ֡z9��;�<�c'�}r
�W� �vc����q]��;��wxzq�ǂ02�w�^�x�޽�S��G� �cR_��Z�劊I�*��**
�s\��r��\Ƥ�4ƍ�nlTQlmFa�%E����5r�ws�ڋ�wv5��\�-�t��6�ܹX�-c��`�+�QPk��&�a5�)�)6�DF����ܝָV��1Q�Ӻ�V-ʹb����ssX���(��ē��f�꺗d=�y	��b+�睻�2vׂ�A�lF�J�8D��w�jN�Î�"Q�3[S%f�1$��ot-�ڃ�&�X�K;��KX��	.���8���X��c�u� �B�e�9�w��zw�<���aC��R�o�w3F�[b3��}(k���i�O�m�'�$e�
�S���O0�X�U��Y���:/
���N����mۅ�;i�J�d�s�1-vFc>�|ida��,��Kb�O�����nv�7��N��e�}�{�l�X�Eih��ۇ�O\ڥ�>3��.�@�?x>gՀ���)�v�z��#em���DF���d��c�EB�]�9� �W�YK3,PI��-��ݰ�#�eu�q�}*���@���
�]��nc�g=X�ΐ�a�P�_�o�����kiߏDum�� �݉��^�-Z�@֐����o_�t��g��o,cHm=�g+�-����,j���r��x�������}�'���e'��X�;	"LE����(n��Y��`�ݵ�
�(�r�����){����9-�fu���]-R�;�>��I�o�.��xa�(�s"�gx�:/�z�M~x�;�]�]���}}��;1�U�W��[���q��	�6���gR��]���j�����i�3Lk=�W�P��K�,�XF���������eͮ�S#���lf��p�eIn���T$l�HW�S�[�`39}z��Q�Cل�,��Sn�浐� ��%ӜUR��T.7L\�Ʈ��	]B���T�=�>2H7�t�a�r�C}�څnlPnܐ���]�rGO`�iu2���Nwz�k���v�"�#�p��X�aN
����NTl⇴��u�Yd�y/Lm���X��^g<v�4V0����*�n�9�qC7:ɼE���q<)��DS�4���֭<\����o��70�yvc�=�S�vu)��1�H�#�E�1��[�Jɞ�x<V}b%!Ɓ�;�����yc���oi�?��?��_��3���18�b�6��,�]��wqz6�z������Bħ��u�kq�c̭��3�N���9���K(�Q��:̻��}L�Ր@��l5�ˢRok~����,Vi���&��ey���	T@QY𷚀U���H�u�oLV����#�${t�6�E�7Z(��+���vqO2�#�OEn«X�'�E���W���au6��*ݨ����'֬T�6���V,3������������M>���ߓ�>Ʋ��)�pt��ss-Fe���#5��q� �d���(���;O�zy���	�q(RA�~���_n�؎r�fl�;�V�����ߔ%�%��)<=��{�Snn�(C���ع2��l`�|�JF��+�v��귵*H��;���at7�ag<���0��)�";�4�5�a�:�yr{�F�\Y�:�Q��,rƻ5����L�nn^�BFȻO���ج��o;����:��wή��]�iu�'���\C�§c9Rw��u?@��Խw�_l��W�/�ߜ�����U%���+ǚ���d\}irxGk3��{"��v�"�D&�Q��u�Ŕ�j��_(�j���]�C]j!S���BV�O(���x��]H��+�&�	��g��"$r���	��s�ܫ��U�Ż�M:;��Q�fd���+�:���<�=Yj�,=�F�h|�4N���h�������Y�&�큎 �t*p�"i�9���[a��6c���%��݈ٔ�mI�Bz�̏Nr����;t�K�!]������)�/���+_F�5ن�:�$�N8�;s�=z��\�����_����B4�b~�1?U���JK���lk�rcs�n�c�g(�ާ���vӮ��A��W�Ff�YXzɾ����:8%�Lx��{+"�be꾪[	=i�=��Z|��c��]�Ȟt;�׹���6��C�j��v!������O_Ok��7zj`�r��\S�G��%����2�Xp~}�^��Q�յ�?_m@�4�G���It���=�.�/s�v]��8���x�
�i�3b�h�-6Q�ݸ��N�o��{aVr޺\Dto�t��V)�*g[��%6��os�Y��z��&�[�Z�y�V64�к!P���u�]���z��B05<�\�Z�R���v�y�:p��y�G^�����IR�=:VJ�dj����A�9���mCj]h߰����S{@FoJ�f��ܣu,��ι�R%;v���]�]Cpj������|��ν���jN1e���@�q̢��o���z�$�'ދ�wp3����k��R����y�}|��<��I/��A���Mq�	�E���	�9�%���GuB!y���!/,kamvl"�J5kY�[+�|�(v���;.����'�#���Gn@�#����Ò�1IM�=��)�����1z��C�jA�p@T]tB���k�9[��+�3B���og3�N���ts	q�I�&�.�>���u�}^�]�"��
�&-�NV,�\�,��mX�f�������E�g,�u8c+;��+�X�����+�,{��6�z�߂�<�Y:z˯\=�������ar��=6��=�K�[��ŝ��v ��in��HBs<�߈G��K�拯y �Eih��]a�s�8�U�Vi����L1Ov�?eV�~ޮ�����1�V�����Xss؇���3�v�����6H4(e�n[�롍�o��9��s�
�=OP����j�kb���J�����ȗ��t˦̱}�������ɴu�P
��c���D������������n���]��Ӿ��͵����Y���nU��3��"fl�Ĵ��v;���d�Cys�-5���yr��M�}��,*v+z�����f�3X�#)��^�P�Zm��|��g[Ohw@��BQy���w��.V�2���DI[S+z���kv��������+#2��Lݰ�B��,w(�wD:���~�H��4U��O,sj����%�/5!U�Gc���[���|�ʧD�B��jV-��j�#�>W+��,=)z�櫨����gl\:|���YV�L�;)���{L��Į�u�i\<ֲd6�2��$y��Vuf��2]h���X}�S^]�,Guvl"9sA���;P�͊nܐ����xOZ���ƽP��ğ������DS죉�oB)q��8n��r�X}S�b���w�2¯OMO�;�dR�2�<�1e{9㴑���U�S�ۺ霮YK�W�w��)2�2;�ͭ��ds)���SnS��]D)k5���W�0{�<��u��	��$�  ݻ]3��,��[�u�tf�@$��4��sr�e�o��o�J0�U�P�z�Kl�L�0��ƌ��\m��_e��%̣�ҏnv��dv*q�6��h�y���YG����9�Q�"��ytN�a`w0��eN�9���'��J>�O���Co��Mz.���H|�{l��X	1���u����c��/�f��Fb2w~���5�sn3y�t�0�b|,�V:���Jz�:�[o�<��������\�0�F}Y]^�^qf�ɡ��tt�c�4�ѼОq�W��<���]n!��N�,�e�~�b5K��Aq2�X�B���� v�T�>�$�m��x1�f]�U��K+��GT���S�Im%{-؎��]�g����/�:5sm.�M=�Y��r�Dt`�|��R�+z��șҳr��t��**�W�v,�y�F���luw�� ���*h�[������}��"���|U։K��,k���k�7��N=��#��T9�ڪ��(���]ۚ����)C���c�fTdO���XY=-@ۥ��Yʜ�����e�.o�jǓ՞�ڳ��{�]�<Mhl�<O_m4�j	<ۑr�s/CHzݴ��{���~�*Q;f*���`��Ul�~�s�����@p=�?@�Jnd�+)wXW�9{�b��R�_��g}�E��Nn��l�By��i���-yp��eo&����7�dv(�$<�J�{�F���=0����]Kr�']���:�{���=Œ����#o;�8|3��l��v�K�GV�(sY��X��<�	�e��o�-�t�V��G,���h�����aMa}9�KD�6�ٓ�j�G�vu^��͊��Y/��O���w�o�B�-���c$��GP�]���-�i�Վ;���LV�S����G��y��Q��J�Xq+��
���.ǶQW����plEs��3�oO��a�/U�Rv~���~�9oօr�.Uᴼ�/��'
6O����8�z�]Qt�U3���֛���p���f�f"����	g�eu�q�D��.{E ��1ݺ��+H�%[PuJt���㏱�ÊFF��/3r8������\�ִ��;\�n��V��%v�+�0�E݀UE�
��X[���:�*o��Zf/�|��Mf��Wa�T��Ow���:���k=(���Ɛk�ڽU�5w6ʏ7 1�y�3k�q�}��X�
R�?^-j���S��x�g�d;.��Vm`��HO��ʂ{o�.ؖzȮ~[Ml1��N�o����
���Ŝke�ʠ�K�g{މh����r�%����i�*�yz�Y~{Hm=5ؽ�V��Ƈ��OQ��(�'9�ۺs�ނ>dT�;�B����Z��3}zd	<�;d��竟��Y��Gs��x��:��@�F��v���]�![��6xN�,��Dj��)�&�(�qʝ�j�d/5B���z�VF�wj��}��eWdw!'oq�N4�ˍ�]�����_GWLU��mg4��!~~[l�f�Hn��~x���o���;Sb�v�M:�:aq�>pݡ����/b�t�'WF��Vm��p�\h�I�����W���>�	#=��Nwp�b�Yʜ+�:�,
O(���+��!i�$6�i�.J;jl�������i�ܚ��c���.��ݦ���<�i����t���[�rdY5�$��K��c�,�$c�W��w�.�<X�ȼ���Zƙm��uF�Ϳ���"�YB+:����*��vL�PD����v�ߤ�b�8�.3`�}��G����elP~�#(Fn���Y�
X��e���z���.�l�C`��zd��1[���7ZG<ʻ�`���ho��������۠�2�YJ7Y�LEwO��]9�{�[̜���2���5u���E=Pb(�Ý3�f��-m��
׮�W!`Jz����5�}�2����2���۹)`�E3�Fp�������v��(o>aJY�"�S�o��q�(涯�t�͋݋n:]�~�\@�h��|c)��^�P�&ޡO�ߥg^���A!¬r���(K��mDW��,\}z����7R�%u!���މl�9g�������_wdzG_0=�c�.e!��m$��3K� �d��_z��#�NQ�]���LZ�9�|���nuH�N���� r�0	T
R7��ne��"�Y����{�����qF�r.�3�r��n;��摜���Y�qU l������8]+,�s7�v�b�f`Yb`.�qs�{(�<��E�L�����vY7��9M�@�t��kd+,wh��g~y�x�Kȅ��`�j�Ӈ�aH�� ��w,2����v��1��Ka�u�YN�\�k�� ����J�Y�Q(�Շ��8���X�`�>����i�B�x��I�7�I(��+G)��]���zb�8F_s`������[^�\�Op�8j�d!� ލ��:���-o��X�澀������i�E4a�Ȇm*���d�c��o<�n�ֽ���T���.�Ō�T�F���=���0�uˡ�i��|)�)fRy�Sh�Yr��y'�7�x,{����4���&�����P㬈gR㒣�Ƣ�CK'ޗ��G�yf�V��X7aJu�ͩ�8p���c����X|i�8�d����]UZS�x�mr��c�$�_ӧ�3.F�~�+z�r=�S��O��\��n�H�c)s���.ެ��:�on���j�\��M�;��%���A2"Lvd|�K*yt0n����8���,>Nf.�J���$�׹ˇ���x�gx:F��(>����r�Mn��v�J�]<���Nv�ֱo@Ӱ�����=b���`����е	��6�:�8��h��Ozi�ecƊ�Ͼ�l�B�+*-�d�	<;�Ԃ�66]`���fڵ��kӻ	��=ٰt�4�%C��O`��v'�.s��f�u��y7�2L=W�)�]��lJ��ܩ��ƀ V���Z�&B���p��sM��#�����&��-ewJ�0�&rf��YFt��?�r�G���
��kٵl��J�����y,ǯ�,���v��\�[�OFt�y�Rۥ���5�*���=�Zꛘ�;���-���;V2<�L�dGy�͡H�z�5�v��4.��Jwᜓsow;V;o���ճkV��Fա���r��_���Ӄ���9���+..����
����R�`��̗���x��t�QJ6�h���L�J8�!���C	�/{[��B��YӓN�z�3�=컈�gc�<6C��p�GH"�a���7������nS<�/y/(om�,��u3���S�����9;�Zܽ˗j��_���V�W��ݚK�|6��g���x�	�(q���0x�:��V���3�>.z��V�TVm'ج`y)�}ZV�gV�n��Aɹq^��K�jhn���z8Q2<�;�G,�b�R!���˛W�:�Z^9��3��δ�]Ü���r��f���D�-�G8�����#k�{&^�޹s����q�V�76�g^��<�iԖ�F���u*r{�o�pƷ@7m�by�<����ɧy�]�j%�i�hR����R����{����Ջ��ۢ�����m,:�>}�'8i�BWWY`k9{��F�P��:���s2���#�*��P�Mb)4l��\��N�t���N�c\��7.cd�.,]ݢ�r������û���nTl	9�Q�,�5]$-���+�wj��\�W-wv��Ѯ\�c\ܨۚ屺�Z-�c\.U˖�b���wk��sW5E�®j������nsk��b�6��n��6�����5��-���[�wv���ѹn[��Ȯm8m�h�]�cs�\�76�]����lk�\�pؒ(��1�͍r�������?;���<���9�Xv6��]D��Qu����LBe,V{d��#f.畍�y�������ɪ�c�	��s@x޾��wo��N���8�f·ʝ�c�^m�s��0��D�]S2��F��W�Q~5&D���z��>�0%�>�����Tvm���[z}e�>D�C5�_7�q4�||д���f�l�z꒢�d���b�{iѐ��Y����!K��rR�j!�`c:`���W�:��ې�Ot��#��2�����SP���E>;����U�T,9���]5G��G.�PP<e�"���0:�G;@i�|�����ˁ\��6�A����5Z<��A�4�]C���Ab�ު�~�%V��s'e�U<'7t6��ɛ��@5��_�'�K���z�x$ЕY�q��n=�p�<�}y{qގ���<���}j���?׸_��k�a~�rr�U����3�W��]o����;GE�JY9q�����Cx��F
_9����^�#~�'�n�T�P/����z�Ow���|������Ma�� >�@w�h#����J����5�z;�n(��y��^t>���=T��>'���/���)s<r)H��A��R�{�ss^�W<���N�F=7� /˯z�3�YMb�<�9�9��cj��t�e�O4ͫF����[��T�v�>�jl꺤��Ě�Gy��g<Y���5�c0;
�.P��μވ�j�N�L��MYVaMu��et�;��N��<29Ջ�}8�k�d��������|�/��	����OA��WF_��r7�ڤ�l���Jf/6�C���<si��!���w����7Ы/��7%j��'@����Sڽ���h`sמ�׹F�Y�x_��Bj#ܭ3�}%����J;��:!�y���(� jFt
�0$U.��ܫ]c�]���b�[s��X*�+��r�k�F�u㨟m;�az�K7q5(��:�w����w�!�Z���3H\����c�z[V���m���n�o��1ؗ�,��!w��cMtgp5g�K���:oH��_	D�U�d-/�&{��!���=]q/�23�i�=��o����%�%Z�W�B��Sq�W���J�tn�ӏ{��Ы�ւUJz�FOH�^S{�f<����P� <�M��[�%U���K�h��])��^�#��xG�LV{=��S�ik\w�Wtmd�M܁���o����ґE�߆σh�'���;Rc`�c>�9���σ�{\*�Vο\?}���ǣ�r|ʀs[�o�¡��{�yTO��)���89n��w��y��я5�������H8b7x�|��{��3����꧱��8F���m=J���Z)wQ��I��3�����gk�[��r�C��ۄ_r-�H�\�;*�}=k��ئ%Ok5�R�-�i�=�:n�{kEOGtu�O����Ӝ'0�u�v�=�{��^�f��D�W���X3�p>��Ѯ�3�\�c�Ne�fA�0�OM�)�r�}om�U��/TϹ�������;�C��g-������\c̺��9�f�A}P��U��Od�ym��ȭ��ro&U[ӓ��MS�!�K�7�q�����x�e��>'�\ʲ��\�%�)�P��K����q��=L�� e��$�u�n�އ}q���B���¸�{b&P�:�������޷��y�{}l��8�����f�^��y;,�>N[=-T<��q�[=���$���+�����8(^ގ�@0z��t��U+��zh*�O�`�P�Q���p��0�{�M�8��W^���(����1\?�?��'YZ�{��䑸��ի𡪓������C���3Jbf �:����@����o��:6�Q�DTf6��
;<�W�MG��Ĕ��3q��ЕU�ǈ��IQ��z��'Z4����m�;�&��.o�@MA#L�J�T@�Z]z L-7��_��ܣ����ëh,������)��?9V:�(;!ws9�s���e�iȾ��w{_�yry�ӗw'��WNİ��ٿ�������1�����m��u��N����w�%���yx��<�\q}�xö�����âᯁ���n�ݞ��f;l��il����6� ��^fn!UT�/�+��fu­��H9��c6��ϑ�����tdE�f��p�[�i��Y��ϙ/�׀��̐����HZ$i��z���G�������KK�p���xk��rBIu��䝚6����dT>����1?V�>���	N��m���Z��𹇷{$S[{~��M��W]�8K�L!����r�:���޿uǡ��S7�
˅-�^�9���r�J���k`������zYG֧n��x��P��tj�����S��k����	ю�����1'+�|�0����+	�q���o��6+���A/�W懦ea.9�ϣ]S�r�6��9�\���Y�;5�<x��Sukl���p�>
�����*��@�Ju��Cyq���6��N$�ˉ�<z���)�Ճ	�o޾�S��r1�O�ว!��a@uaWy�3�S��c�\n��F.1����:��������u�S�7���b�eq�R�4{�*�r����ާ\��ȹUg���hZ."������n�h2VP�3:��\�(���y���{��At�~�����v���}��7�oNsF�iq�le�x)㡃�v�����)���Ǒ&1bfk�1�8���z�eA��0d޽%b^���@s�RY19:�yY�Wؿj�zC�
�z��.4g����uR�/B��Ahn�s�-����sW�۔ӛ�����.��P���ì�L�3C�W��B�R9S<9�|�����}�~���9����{�8��=����T����~�3��R �5t	�%P*��to%b���.�7ɽ�g��_��Jw�}�S�{Jdx�D<w#.�Z3m�ͨ#�$<�@3�:��{$tNs9.�oK�������
��c���G ��%�Q>اv̋�UT�R%{P�m1�˹�����@ɀq9�qNu���W�ٶB�����Y�s�J�5��d�:��	���5��򦺍���혯�^ӣQ]�XP{��B	uU�J�.��ؤ5J�wG<�������n0
\=p+����I|v�E}+k0��)��ʅ���ylnkS�>�R���	�לFN<��7� �:`ahP�e���^3=ai���)�a����#V��u6�}�3o�=���qq޿\g��ޟB�@:7�t��G�k\�t�������.R4��u�1d-^�}b�9���BіU��f˫z_i;*�-TFA5�7u����t��m>��k�������~yaĖz'2�')�$0�����AA�Oi�M��>��P�ǿ.�� pu��˾��k��ұɲ�VS�]h��s����� `��i�ۅ��xc�8�g�=�b���������_���`����x��Q{����)�s���>���Y9d�=on�WD�z�fY�{Y�7�����8�=�k��K�����9���a{��v���}yH	��|����=��i�SZ��Ex�l���%EyP�.e1�z��'w�3ƌ�B���q��H�ePc�+Hs�+İ�f���+�Y�i�?R�N�1�U��5��<I�Q%q����7����{�Ty����Ë������=�~>�!���p�L�,gB���g�R<	=�:>�W.}�nc��;gַ�<�>�W���~��_��3���V�%��=���y���9�2��|
7�*�w]�#@�����ǜ�^d�4�1qS)9�/*�W��|0z9c��Y9����;�a{r��q��>�Ύ��kD�z\�q�@Σ l����>��(mv;�ǥ�hx�m���n�U��\���Q�1��ŮFu-��k���on$钎}�@}��[F�����]]������u���x��ۉ�����Y�}��*�H�t��!�ٰv��:O�R�+��B��Y/sk�V�3�hO�δ�ǒa|�W�ם�T�Iun�-��i��/��8���=������=5u/Zg�u�m-J���f���9�\��P0���k�������Iցr��q
��M��I\@B�tz"�ӕq�	���l�D*umШ�#�:=[
����=�n��n�Xϡ�߭�r���\GL��pvlTJ��P�P��~˅s7ٮ5V�[Vv��;������Tv;%2h��|�Pˇ�p�saҝ7,t��j�[�F`������k\�Xi����u^\/Dw;�1�Ĺ+�P;p���}G٪����o����v�4�\��X6�{���9��߯.�ޗ�]s�L�K�~��}�Αi��� _����#��	̅W��Y��>v�i���U��q��W����}0� �-�4�]�z����V/�68Bd«���uҝ�a�����w*A�S�ٰ=�:�/̏J�D9tƾ�O+G{��\cU�z�+'�D�e�V���7������V����:���ʫ�o�;���XW�@V�e�D[�l����o��yj}Ǉ�����ӄt��o��|�Y�Ӝ.�럪�5\�\S���-�e{K�������z)����Mg[=��jЏW�pǂ��������O���5E,����=F�rz�l�p#і�;��U�u���R�����h���Q9�[�^=����V#έ����"��~b]�^Qt�8m��#������KT<4������8j^�3X�Ѧ�/w���L@K*w���R�>pg@�x�qR��|�W����O�`�k�Hg��v�p���=�T�w�é�z����n�ſ��K<8���:�q"��H�T�j��P؅I�}�i������=.��{��g�%�8�!8m+w�}R͢ r�1�&
T ���A����=���.8ګƞ���ޞ�o v��+�?��M�u#n��7T\�" jj	d�P*����T6L�����7��׋��ZY�ݟ��u���G�9���'��n��u�f�UIB�����@��}�"��֟�}��zrU�T��u��P��ry9|K>��̖��ͲGMK�ާi����۪}�]ő�4ӳ�и�=��2V�tB��.���$�Ѵ��քǢxשA�W���ѪM�4@y�����wA�1��x=���C+����UC��2z|�0h���/T�q��?s�vn��fOX���'0ºu�n���Ѵ�
��Zu��-���|r�{^�������#>sANN���ێy���F���eB�K�Ea8]��{�0��x�~[��3�:�a�y5���3���Yq�Z�V�,W\�ge3�5̷v�\��e:ܴ�z��*�-Y��?ر�On;^�T9�aͺR]�ݤ�ծ�Y{�Ǉ�86��g��n��Ï�Ok���)͋x���j��75��ҹ}Ʀ�ЀQ�7�m�ߚ��K�UKI�5S(N�����yY'=8���E�c#�8����rju�gF��x:FGi<^}Ϯ�Ms {�N�a��#}��1�N��!��Gɱ9s���C��x*	��zO��ˌ(�*�W����
]6uC�\n������<j1�^Q� 6��u�z��O�2Ǡ,z�_D#��ɠ��U��A��:nU8˕v*���ê�����#3�.��Kn��Ğ�3��B�g���R�/|�t^�-߇V���/j��`���PՃ���ͺ�Ӵ�|�+���J6�UA���B�2����̈S��|��=U哄��8׾����7!�ײB��:�e�wl=ĭ� SRtJ`z�zz�v�qnu,�+ӝ����ӌ�;�.*�+�>�����NF���e�N���f��K���W�g���.u@����Z{6t.�N�1��m���a6۸��wl�,?�{��1ꋂ����jg��JQ��3 ��9l�t�Y�@,uGf�
�[z}e�D>Dzr{���Ҟ�M`���d�tot�=�ЂEV"r�6���b�i�s(�EkL��Dm�wCΕZͥ6����C�	M���=�^����D�{�\�J9��I���1Lu�n�r�;�˗B�n�ҭ�)��ύW2��J������]����u.&��#���R���ʮH��GY�^���L��<(=��!�K��^�ftQ���>c���K [�2���\��h�`����~�F�'�v:uK�������װܔQ�ӹ(Nz�[�3���4ќ��r�n�_����e��u�3�(-#���u�{�,�bo+������j���+E���{y]��-t�q�t��u#9���(�@5��R����+͈�w���V_��f�ٝ����H������xcГ��}�ڦ+��^���9��sUx�_�C��B��S�&Pꁓ����NY9y(	���Ё��p;�N�BsL�G:����>���� �^�������}��az��(]zk�팤�+�E�u>~�*7��ӳѳg��N����oJ����ʜ�ɔ�M�}5�;���6T���T�VNQF69kş����~έjk!��}�|�>�	���$�!q��z�H/�����ū�z|=o���w����L/}����9��������1��U��zϤ�x{bg@�QW��̔�i~��R�Rc�s�6������eKI��X��kM�C$r��ln/�5��A/O)��R�tw��A��h;���N�V���}G̬{�Mr��tȑ}iͻ��z�L�f���<�<0U�-��;�u%�6����Ӳ�m]�D�� �-��;tE)�n{|����ʷnTT@k�9��������)][�d��3�%y�l���0�n�bB��g �2.�m�ճB},1W�=ҡ���+8��ܑn�]9q*Y),U�ۆۛC�y���q� ���kg&��k�͒S�;c�Ąg�!�Н�Sx��|�k�Lv*�J�����Q���9��m5юǒ�=T�b��0W�wD����5�Ѓy�pF#��D�Hn`�:�VSTˊ�q��S���q6ފ�3!�4��ϔ�#�yt�:7$L��b�F���@�f��RB��G�h����!�y�z<�N�ԉ>ʸ%F^�5*i�]�}�E�,�zi�k��#V�����d_2�;���LO�
v���rX�����[��>:E���]�*!n��Ys�թi+�n5>�f%����{��e��x��=^B�^��H9�p��t�F1J�����y����3����;J�`�{p����P�RQ[}�=��$feO�zTUZ��S=�F���R��ۜyg�v?N�FoM�+��#���4\"��ۺw7�*9l��R�^X�{Bl����C��>�n�r���G��Kd���M>�M��Hu��:ˮ����i�S���v���`үD�J��Y�u���5�xt��EU�����I[�i���z�U3F���;���_�߈�\�d�>��>��[\��`t�M�<�MW�.mM��Yvyr3قyŜ�Q�+��M�9�iCC-n��O3]xs��&㦰7o'��獻Dvl{�`��Y��N�#|�iv �+�{��c���4\K[����&���W�z{ϳD�7���j=�8<�c��%�H=8-뙢PO�8�]�yP�Kq3�@��kޔ�d�����HŴ��p���s�\���������!�Y]��;k9<	�����J�$�[ۯ��:�偤�h�D�L�^u�[��]�2	���f}�w.�Ǫ�E�3{4",d�<pK�����,�=�j�PJ�\�s��Ӻ�:��-s�"�>���Gh���Ƿ��r�5ɱ�/�s��:�B���־�씦�U��%e�Μo�S�!7�Y�wVͻ᳞���Ǐ�^��	�й�����5I͍��ԧ�V�	�wM)�7{6b�7�ל�f����v$��*l4��n#q�=y.��"3�Cv�v��M�`S�՗˅�է_nO�Ɵw���[�z��vWɭ�H$Gv�wnUʊ�wv�۝+��*�5v\*79�H��r���\��3�-r�;��X�s�-ʃF�5ݻE�+��d�����nr��.Z�wv����sj5ȱī��sguwtt�-�KD\��ō�ZH6��I�˙��I4sT�s�ݦ�F0��Y�p��\��(�K�NqRT$X��W+��F78X��Z+�Y�RnX仓s\�t�u��ۛ��[����;�c9ۅ������Mn�拆�r㢉��A�	'�I��>�nY��s����.� �ek+wI�0[{�`�Թ�2�S<���͝�A��H�xK4œ5:TX����n�]ە��Q�$�L~��\���������,�)�v�Ϯ�י~�>�`�r�d�̭���xd .ٝF�@�s3�ϣ��X*�+�ܱ���aۇ��s�a��>�]^x��7n�ǡ\Η�@�`�@�����@(mv;�ǥ�hz��3X�k�N'6��\yi��&��++_:_��>3���a�����/���E��ɇBc=Q��˿� //WS%��g��ۜb%��&�UT�n8�+��H�?���Z}X���m�o6�Mn�Xwz���o�\����M��� y�#^��[��3�%��ٱX�yf�~D~�g�X�v,�opz���L9��RWtmd�&���~�j�[�8E}μ)˵���s�m�;�!{Z�)�w/��Sy+Gm��z#���bqNM��*��G�s"ddؤϜ������d%G��3��9�@��u�����qJp�����/.�ޗ�]sӬș�z�ڋ�l�ґ5�Q�J�p�y�^:�'��0��Na�u�zo�S���������S����$_��UZ�o�6��^ډ=�&�|I���K�A�y���2�����*���?_|l'H�P����U#�|^v(�ڼ����r�]��%M��Y+T[� ����X�W��DW���;;���7t���bc��뜎�̽�M^�%ӾGY����Uk���S�:̇�=��c�����8N`0���q^��qE2x:#��zUw/��me-x m��.:�G��Lk�Ȅ�s^��VQ�Eω��L�vc���^��k\��jC�/�;鿰�Q�P��e�[�l��ls�!x�e�/���x�c5d>�h+S�=g8u>�L��S-L]9���2�]@��vYtS-���8ϴ�]�
qs����ѯ�AUg@�W.����K�>�頪�?1�\9C�$��;N~+奍�t��A��N#,�3�i��K6�U|g@�{�\�n*g�?//`��:��Y�]ҋ�����Z���4��Փ�|[�P��K(��1�R���z�ai|�� \tvl���Ĺ�^c���Ȅ�F�p�Ԍ��v��uE�� ����JU�����[
k=I��dk�<헖z���k���'i9��������x˯33ʹ|'���+�z�c��U�=�[���4��.up���gx�vh�W	u�)�Ĳ��2_��Mי"g5e��ۧ't�^=׵�K
�_h���6#v�\�r��h)A+(j�Z��z0U���s��R���3��O�o�.	65�LΔ�[{���k��0��`�{ջ�L�WX������έ��ӗͪdCz���g%�L/:����x������UbDvφ��Ж{Ʋ2V��D+���_ܓ�F��\��!Ǡ�E��^��W�*B�> :ͷ������4׻&~_��X�1�m߂��wBc%�^��խJTkv��2�9� ��^��o�TwFO`���s-��Y��/}����4M��>���R��.�ٕ��7A��
rv�|�=C��]r��|l�T+��>=�)����O�<KN���I�0�Lw����UKI�T�3�e�י~z}'�:p9s+ƽx������N;����w����Zo�)���0��}p�:�<����\oz!��7c�ʝ7���)�~��L��n�h{�͞s:=�~��G�JC�(�®Do;�`z;l�;�����r�[��^�4�?-˦}���fP�:P��|n)HG�M�® �rا�\P�5�v��z)?����ş�v	g8�k*���'� �>5�.�{��c����Af^�D�S��w.e�f����o�U����D�s����|�+���}R��ĕ_��L/DQ�����Xg}{c��Pȗ}B-uy�"%Jgf�h&��a^�WR�x���k��N�ES��
t=��J���&�/<�U1��oڨ�rT2d����ƥt��DŰ�R���,�^�&u�-��YV9�ٍnϷ�@%4��U�=֔��-��u��o�B�%�=���!��������s������<ꑗ	ݰ�g	W��H�-zL�OM�c�^��>9.�z}��(�/O�����J����3�S#��H�V��7T>��tN���Q$e�=�8�t!GIͨ
NxW�i��Д��0��h�9���'�@{��C*���k#{��R���U:n6��� l�<�h\R�g=�,wf�c�[x��Y�F�^��q`��F��\�c�'��#�;l��̀����"_W�tkh�N>\�Ê����'/�|�%>�=���V�%��?|��P����~�F��$�6v�*%mfE�V"��ǳ����z��O8\o��C��]X�Vݰ4�}���.}μfz�>9>��ѭ;���Hϱu�^2��4�5��﷝ޕ�@tm��J�c�t2f�5��_�Þ�K��Ud7~x)�S�]z�����8n0�5y{p��T��I�s/fX��<A��WD�����z����e���~@���^�,�M[8'��Y9�t�������N�/L,��nY���e��OS�yG+E��u�ۺ]�%:Z�p�&l�6QH�!���pu-�2߱�%��%���f�A�Cl�.
��:�{���N��\�/��w��yX�����A�4�5�گ}ʸ����/�,��}v���@�[��&���\��*��"Jl�gf�c{{�D��_�GW5�x�8��p��̺��p�ˈ3����Ma�� >���د���W�m�7UG^f��>�5^�˦��;�����x�]q�E��sA�Mq���6]D5��G,B��9� �����7Ö��*�<�ssY�� ��N�1�U��5��t�����﶐6���b��>���͛�Vّ�9�ڦ�.�c���G����5Lo�V_nJ�<	=��i�LM��D�^j::�5�L�1qR�����5q�[���V�J;~}p���^u����>��s���2k�g� �3:q�`$�$�Nz�|)ĥ|0{�X�q�G�{jV��R-^^�����R�[�Y�u��=D�(�R Q���^�6��c�KjЬ���5�/R$�|5v�*:�8��n�I���p�;wq*h��@]�@�'�mK���\��N��!<�ؚ���g�����ݰ�%�f|6ۭ �w���OJ� �K�9�<v�+�f�uc]��{'i���}�¡�r�ro��p.��B5�*!�[�U[����Eu��F��X�y���״U�k�G&y��<؛�ٚ����x���e��*1��t���'M�No�E��ه�����/',�{�Y�ڌ6.&U[�����[��-��3S�})��#��18��>ḝ6��.� rXJw[7(�F�ۙq��if�^�T{�1��c�q��r��xj3^\$�U��̚7�_������P�u�ɨ78�V���]:^�nXہ���=���b�%a��\/Gs���✛� ��s�|}�^#;���}�|f�ސOW���'ߪ^�쌞�����o��}a���kp�7T�/�|>�*Oc����ݳ����s,�>��a]z���S���R ��F+[�����HnĬ��C�*���k�zs��X1��C���xVx��GV��n����%�$�E���_��ߞ��}dt��AR�-�	�h�CY|.1��Vu�*6�T�m�ҩr������{�K�W���Qp��uaTo*�]d[�l����o�琼j��?7����&���fFT�R�>q3�`��2�b�H�6�i������e��'-��5p��gX�ǯ��z���z�x�)�4������
��S��d�S��AU�'�0{\:C;�r�A�>�����l�ǉ\v�Mc0���J7�%T�&�$R9S<9����&[ٚ�O���ޡ�Y�	t��m�C1�u+$��+A\��*/pny{}o2Ng͛�H�Z.��:�KK���Y宐�ჩ�P���t���]u�7AP��ͺ�;iF��x[鎀T:9p���g �&��!��ϴ̎��Ž�"�O��V�;���մ��}G��+��n�Cᾩe����?�
;<�P�E��������b��n=��J�nS�p��W�����H˧v����Qsh��$i�txe�ʩ`Ή <���[Ӓ�1��.��ӽ�*��������|^�pۼ�]y�S3%��2=/�M̿����d��u1R^�`)���P��r{���,�m���k�]��/�V��ۗ5[��j�7�5�H��*��$.߆Պ�:��=��%a��D$���o$��ݓZ��o���Z���|"��RF�ќ�����t>W����/�K�W��v�XC+����ࢲ]z<Gf����:ﻝ3i� ���V|2�Tk��=p.am�'0¿��a���/C�g���X]�ј7�����}~�=���F'A���
v|��ێy���k�NP>��ʄ]LL���^q�c����qwI�F�z���XOt�����1=�{��ߧ�}����/�o����G��,~�˜�U���'��c���u�6'�4{!����5{�c����y����|m^����M���-�be���Q[v/6{�g@ooы�Z{�+��Xf �[�~u��*�̓u�.jQ�^��H��;'!����\u.�#�� �6���+�����ۏ�u�iH31�qLA)[�]]�5��`V_��w'������n��̓�	b�&tu�J���)H}7�W�U���w���m��)��aԿUaQٻ��0���7���r/[�*s�92���bgJS/���4{
� �5�U4��9�~�~��� +�Ф���\��8��kn�����>5�."�{��U_BlN1�g
#^Dأ�e�|j�'���
w��D�s�F:m�h=>�Y\�o�Q�G�*������A��M2}�v,��̯S͍�d��ˊ�Й�B�ˊ�����9N������N��3��@����NZ4q���� G�`1ҙ���+O�ߪ�W�B6�a��9v��-������S�ޓ3��0��	_�\F�x�6�u�NxW�Z{6t.T�#��m��8}B�7^����F�cr��J{�iBUkmZ���`�2*zql��,����A�Ovn`�h�'���׷QE�>�{��zC~w�ˣ�2B�;f*Vӣ!w��%O��g���p�ؔ=�z_����+�ҦK`�<Ш��ǮG?[�q�I|o��A��v]C��ӫ�&ы/�vi�����{��
��:{F)�!PW��{څF
�c��QM��Ii��ӵrgA�f�Q�	@���{p�F��f�B�]�Qu�1����gI����?f��f���5�V��Kx�M޹����c��4��Q:;˭��B+7>w<~�Dn��{n1�l����!�n�_���z�g:����}�gDP�u�Gz^Ӡ�Օ�o�=���iXj��p�����O��Ѹ�Bw����lbSQ����"���M��׿���,�py�2pm�^�2�*^�3������T���'���S�{�Lv$:(
3y�X�D��ԏ��5��s�rr�X��d�WS�8'��}�(	�[�B��^�[R����i�Ԏ������t濟^ዌy�Z|��+��	�9���R���ӊ�Y�F�p:s-�!�S���NuD;���O+�5�=|Ou��^4k�vĩǎ��%��e��%�W����=T^�
�*����A����cT��jk.�z"�<jJ�����]�nN�E���[�=�⋀���H/it�}�C/=�ᾟE5Lo�e�^���*�� ГN�=���k~�m��z��T�9��uȫ2�y*~/��YZ}��(�����Y#�<�����=�s���W��6
.:��:����1u3�Ͼ��X*⛵	�����Y�x��}�Gb�0��зYM�X�^���?b�>�<��W��]P�E<o�k"��e��n��i]{���A!��X����j�e��kp,�z�[Z�ƅ���si�"�7:�ŉt�5�+g���]{&�_8f�}Ϛ�w�� ��f���h��w��OW�1���]q9W]�����P@�F@�"�}5����b�l��s�?P�_.j��8+����0�x�'�u�*h�q�@]P$��}V��cL%�+�.3�������|��=��_��M�ۭ���&�UT�xW-�@ʽ>��%D��a]7*踊=�+&5���
�u�7	��\9`4&�M��7���M�vp���}��{|����z�r;���Q���5�.�Wtmd�&��۠5��j�Zy��i�'����Oz�Gt��h�Sck%���_�g�I�>����X{���%��H�5��3�sT>ԡ�+S�qY��>WC-u3f�H'����1��k���a9>����d�<"WC�"�Uu'�y���髷�F���L�=��)��VV��Y�}Bs+��=7�)�r-�(��>��޹ܻx� ���uJ�BT�Ͼ�4�����y�C=�'2��//����h����S+�/�mb��E"U�S Oc�#��2:"U1���������VQ�6OW��ኂޝ������:k��8�+�TW��MFLѸ���2G�0-p�
����aLm�wU���z�#]m�V|}���<}/��P���-�`��N����zw���.��Iר�V�.-Z�ԱQ��
���V!�q�Ȁ,nz��f"y��6�Bؕ�7zw�Y�Ӯ{�[��`�V���BL�C�B���lT귃K�ޤ����֝>�=Y��A[j���c�+�U���,#}*-�A��N�ғ�٦C�obٞ�|[>���;�ؘ�>�<�����P��9��͵9�{�n��p��ӡS�N)��+����j����H9�TxmѳS����t�=Z�L�ɻ{��K�6��/ǟG��$,�����+��r��>[��}�K����5�l�t� -g��6����5�v�� ���]t��xv�ӭ���[9t����`�L�*!�I���ٛG_�</��pX�͵�4����«�tC�r|4���<4뭽!r�̃[����dE�;Z7{X�l=�����b$}/��zӥ��2�]���]Q%�e�Y�C�����i�h���8d���f�Ӳ��=Z 9����yF�&#ohk����6�i���2��v�uZ�[s{V]��gg!Sv_J{�IC����z�-�ɀ����d�g��*=���f�S������kE�goy�����=ٜ;��膅�Ա��y�̛����Q�y��*����:�u�'�\�j�`��-�Hr�E����}k�а%��e������
�vr�Z�ӭs�p��e�ε/��H�G9�U���V{0��[޷r\|�YhCequ}̢����ݚ��^�JIW�u�0Lx���w'M��4�b�Z���C��׎;�k[kopI�he^�A������0��*��E/�P��F���sQ���j�.���)�hܷ�|�sz��w��a��p^$�H۫�d�,���r��*fg^Ihr7������c��{#1�y�5n �̅䛰�h��.B��L7c��$j���;���a`3�� �ܼ��K��b��o<�C\(<�1��lڳpF/��7���r��i�'cK$�#z�g��9I����.I[�X1[3գ��WX�L����rqN����p��]�M�����+��[�f���Df]$�<�ٺ_���7�c?���4?ŰZd12�+!�3�*��8�����Լ���Z�v�j�Ӎy�!���-���'�S�l���%sI��y��t皷����A�z'X�����M�:��(��Ֆ�j��@	�q��2��FC��^�x��L���[�A�����.�7/a�h��ɍ���r��/�2�Yn_0�<�s)�{ó�{��
�Or�4ִ�n`H�4,��Փ�[{݁5�h�U�NM�.��ݎ榲"�_R_b���S�>�ˇ�����}6���~��T:'C��|K���d��Ѯo.Z�k��8A#�_|RG�л���sK�����s]��Y$�Dwv#I����X�H�u��h��KJQ� �E��[��s���ˀa$�hs9��Dc��4N�%�i Lu�rH
.W'wE��Gww[�X�,F4��is��9�"776H�t�wH.�RMI���b�+��)�Gwe�iF �(�B�n��D���N�r�s\4�&gun��E�[�#\�S;��9�i�t�ꒋ P� B�w!����ݺMwtLHA)"A%x�k囇h�w��	�j{0u-�H���<BTc�RL��;a��t�\�C��Fk�]@"�-\o��Z��_j][���Ѓ�;�*�2�~��uaT�e�~�l��w���y�7��o}�ߌ�J�gM�B�z�Q��/$��c�&t;��_L_�JG)�[4����N�.��9l򵞹�܋�]ÇXT(���<�*����4Ϣ�H=_�'�_$��Ȫ��}���Uq�������(>����T�輌hs�����WQ�3���G�*�� �* �H�T�n�,U�^��Fe��>�yР�����{M��p��۷p���K6��ʾ3~)Ps���"L����3�����A�꼧�j�CXk�K���W���N�i6�Ԍ�whM�T\� ��#�rc�O&B:v6{��,�T
�ӌ��N�h�I:H�}�"O�pۼ�%י��OAV�U�η�/7����;���Iݐ �|9�
����zL�vh�V�[�'/�g�ϙ/��v�h�nfLoCZs�� �W���S�r:d��6�TJ�f��9�5y+F���]у#�]LT���/�}��p���f��9�@��5�������0���TD����/^J�k������+�ޱ8T��YX����{���x���h:(�t:Oq��U��v�c��-=��2�KN,���J�3xv�|���]�ĵ�&�HY�N�M�9C��k#]Z_S���tDCԙ]{�/vm��i`�uf�5,N��][W��ٳ��/{k/�v���v88�wt.:��`�~��>P+_���0��6+�������rV��|���g��{�i�u�#z�i�'A��:��g�BsCn9�z������ga����y4�:Z���k�뫸��������ﺪ������uLOz�_��d�2߅�v9����b��n#N���ex�ǧ���Xa�x?{��~�S\��N�ϛˎ�}�Ӯ��Q����^����)̩c��'\L��::�]�};PC���w��������z� ����hl���:G[�\n���k�\z,���2��҅�L�7�#�&��/���= ���:u��N q���
�t��E:��Ц��&�T�Y�O�=(mL�<�7���a�������/�?]�z#O�~���Dc��Cv�ҧ��t�J(q%i����9�W*��[W&������ʋtg��T�����J�s���{D-6�F_�ݰ�g	U�k*��ne��L��o� 8�U#�Vj�(~]�ȣ<V����J��F��=	�÷��9�߂)��5N�_�2к������V٨��v=wςSN���Nr|U�����8l+3IׯE��N���d�_�<�q�ܕ ��R�����q��b��H����^�T1Aס�f��if�8k���+yukt�t�1���Ω8}�g�M�.:��d��@��u9�^i���Д�H�/6�=�BNϸׅ46�<��q��Į'.����Q��X�6>����j�Ͳi��GjNx�尿�0=��`ek�Ͼ.|�^���
���&�Tӣt��Nق�]���{d���fhSЖ�#����o����]оJ�-����F� ����s��70��k���Ť�����E���z�.���^Tv�yl$����@*�����Fhe����x��fl��q�aI��G��B��QpT�9s�9�����V�����o;�>���tn<�7t6;q�զ���u&LʾX9Q�b�{�@8Y�������LeԬ'�����ۅ��xc�8�g7�����yW�s�3Y��Z�Y��9�~5�~ �}�+�9�X=�pG��NL^}W?mׇ��}�>nG�7�K�R��SW�ħy���3����<��)'2�3�%�B|gE)�y�NO�˝�v�g�םN}K���AS���M9�w^���p�Ʋ돬���aY�|gj��G�t�U�9�3gНl��-v�{�oW ĝ��A6�9�4��Hҝ�	z�/�d�'u�S�=�z�c�~��4��J�;�,�k�`��x��ݷ��tW��Ӷ�	�{Cs�����V\yME]K��
Xut|���s�/������������n�j��-�W]c���[ =��U:1H�{�ssN���w���ʲ�Zk.�z�<JQ�@�s.�s��G�A��te�*#kj�^�K�㌆_�c�o��ST�^�z��r��ԩv�#��M���?�}ᵱ3,�tECD}`��_�|S�(�W�%o�\�V�=������3����p����R��Ց_M�&!3��$t�0S�L�r�O�lJW��}�6�z_�{��gaaƼR#�����;�ax?T�j��0
D��Ml@(l�J��ο}���t{� �{Ԭx9��A~�cq:�&�㸜7�;wr��<�$y��/7�{|�X����+ٺ�c�|C	5H�IH���%��%L˩��$�.�8o���M/���%�ή�tq���ʆ�}�¡\G.�%7<�(���P߭�W�М���L{�r���i�mڙ�2^͝�=�����Q�+f��I*�<�y�F�@k�MlTbl홋���{Κ�H[��p�ޯJE;`l�;��8.�Sq���v߮�������v�/���	f��W�,xֈ!H#��e�rӰ�x:��@�ָ'��.7�7Ͼ�`݁��[{Z�M���*�/(s�R�XTyK����ʡ��3��y�g���3J�M��-�6�w��;�V;��}U�6���c�����,��T���Lo&v���`|����>��l�k�OP��끕�Ix|2)N��O�ώQ��U��6�+Յ��Ӗ�q�O}z�s��Y�yQ8Ry�^>�� ��3�Na�u�zI��ܶjy{�~�Fi-��رt���z���V��J�|�>s��y��g�c̺�'���
{���M~����1y����Ua��=���غ��s̎�Tƾ�o+G5�ñ��<j�di��o/����~�u�yY69���ѝ�wN�������ՅP�y�N�:��\n��$������a=O����T��>����I=Q2�A:��bQ�B٦W���y;,�:�e#�<<q���p�쑵E_����Tn?���kg��>��Q�`��τ�m~�/B����
�����nЕ3ͺ9��pq���r���p�Ц��~���F��J�3�@�$R/�;��V`Ɇ����XUø��w�c���^� ������;o+�Ί�p�}R��"*�1��몫ՙ�6n�-H�}9,��.�&�sډߥ.� �_�N�i6�Ԍ��v����=�ȹ���b���=|�o�H��L﫠�r�R�*��1+�^��~t5��R��<�(#�a�v�Q�p7Q�O7�g^Wu�e�V���o	����)���
�������+W�ە϶�{���1���i�U��<C���<�s;%�K�xBzwgZ9 :��0�A�P(9Z]xL-=�&����'�[(���w�V'�t��n���G4��3陓���'�l�6Cu®*V��3]�*�]nJe�,�~�������d_��Sƫ�<�׀]6���Ѿ�!u��*u�N{^J�G��3Em�
Գ���̓E�B2��&F�vh�r�k�#Q�P����]�0�ق���(��֞?#���+�����[<�s��~=�tM�,��?Ea���ȁs`�G�*�̝7>=��Փ>���]�����
�����2�r��V�df�?n��L�
���z�>����ʬsǃ(�+j�_��7S5���:fV�Sϣ]S���������M�{�>�>�u]\nr]I�8'�������V�̞5*����*��@�Z�F����P�fH��ˊ�����S�S��$�˙C�&tu�T�8%�|U �b�4*��/jz���޷�`8�N�+��w�'x�^5�\}|Ou�C��B�_�R���z勞M��u��p5��۩���ͻq.�2�큧�m� -�7�%�b�\���«:�~M�xyl?g7��&�u���k����E���g��&�+�dhԣ3w�to���]-�;ku�V/T���]�vK��l�����!u�ֵ�ۧ�̭8��7����ko�E�NvU�iÞ�ׅ\^��I�ge΅�MgMz���Ğ�3��CzͿ��*����}��+��B~^�/}�����厀[7h=>U��xo�Q��x���=�qiT�fz��ü�8*�6AL��2�"�z���J��jqC�!i���T��N퇾6oh[�>���r�Q6�@�Qt	�5P(9H�<V���ˊ�J���
�3�S#�5xd60���W���L3�Ҟ�93`��]�@�p��*�@ـ�@�u9�^i�ͭЩ�F0�/�6$�L���d��N.E�g0�I�N˪fB��G��\	d}4.)N��뜍�j=A8G��[#��v����.|�^f���Q*L�:IW�v�WҶ���:T��K��=�tmw���vi��_GoY_З]оJ�/�̰1���*��n��_��FL3վ�\5c
K���̸q=����}[�Dg<�=���p��
��`i~�f�[��t�m�nk��<ۧFf�a�9>t�0�Qx^�ƽWP�]V��@:7�����l�f,66P�89��2
��+�.�cK�y��#�*��[w ��e���o�$��Ie�Y^!)�8y:�����V�Ae}�Nz3��P����{���^wS9T�[0<V�'B�;��t�euB�-��96���G�*�5&Crt�QU�Yʧ3��Q�G�#*O�)�;���]J�p��y�����^��i፸Z�;�\��T�k��^��h���Z�~�
���3L��O��êN'�pdEt�'.3=v�mXS�M^����l�)��������)W��Ni��՞1��.��'2���������\�,�̻��i�O�]�;�z��"�s�D�i�d;����\cYu��|Ou�f��bΒ���:�����7�d���7N@}p2�1��
�*�������c|�/���ˡؔ﯄�V�ya�D�'4�����Qp9[T���ǔ�S�;��}�1��IԞp��xe5V�n�^�~�
}%_OOT΁��*e)��uȫ2�oؕ�>�5�ei��k��ksA���G�5���)�2�6|%�P@�Pg@����-)���N}�`��y[E�}1Q�T�I��{^�C��ѫ�:���x�'/�wh���o�P@�_`$@��Ϧ�,#|ۧ�����F��o�{�\48�ա��������7��q:eӨ��4Q�� .��DAgo��h�@v��qS-㇠鵁ɚ&��!?x���`3-��܉/	=���Ⱥ^̾�[}]�3x��,V�-��P?]�l��21��62	��c ����8n4떖S�N���ȱ���0��3�����8��V�A,F��yt�Qv�;�r3x����N�k�&Wf��-&��~f|7��.%��&�U:�s����W0z�&r���Hk$������L&uh�K�[�i��_����=�dEI�����M�W��K�}��4�t�k��5����a�ח��T���d���n�+qv�y������z��z���l��x:R(��6|�T��X����~�Y/'�F_�q}q�g�V���,��y�)7���m��������D�]8Լ8.��9��Rp���w!�u�Ƈ8�]�1��K}��s�C٦k����'�u��� f_�a�a�׉S*{����4���5��Ӏ��0ǭ�ﺩ^���fC͗�>�y�C<�	���_^���zvl%n=E��f�|}�Q�N�FW ;Tg�.���Tƾ��o+G{�ko�����"צ�5`{�3���S�&�h��GmEuP�=,l����&8R=��9�+&�lp���?�_��t�}dq�C� L�RK錊R��g��ںV� ���������
�ӊ�(K�,�o���K�d�wͩ�$���e�Y����٠�����s�R�^6�X�<z����J^k�Y�U�+�����k66=k�-�]��oN����ןnn�\��͍ڧ�[���hj'V�/��`�V;���|�k�Ȟ��+��t�?��H���C���{M��H��H=Pf6`������T�S3��b��n=H���F��;c�ء��B9ͫ��τ-�e��ᤞߌ���7S3'�ȗ���ه�aՙ'.�~*N�z9�G|��;p�N���?D�H� oV%;�%���bŀ}��m?80�@����5z���J]���O��u��x�F];�&*5�����-�M�guUߕ/�  4[�'�u�0��l�I�qqg4�s����=��i�@������T�G�욠�������O�$���'���3٢aj]ly�M���D�K\F��>�Qeϸ��B5�*�3����H]�j�GY�#ldY߆K,�A���^�tݓjg�Q�~�wF.NȸN\~F�"��> TG?S�q��'l�Jܼ��Փ�Ff�f������������!��Wt-c��n��s��7�������0��q��H����Ƽ�}]��'��w����'��^_�/5�ҵ�f��uaNϡ�����^��qXC� ��.���zDO��=d�u�!p���{%��<}!6ν��S�.�-t��Xh���`7r!}.r�rI���ݴ�N|�,�+7O(� [�eƟ!L�ͫ�Q��x���*�K�}�`j�f���&ic}�g0���F�s��Uk���<��zNw����Yĳ�D��^�9���|��1,q��9&>���)�����:X{�4X�ù�1�uL���G�u뒡4�c�W�O<�+W�&ŧ�:n��G{;���<���p#����x��[��d�j
K��gz���2vdbЫǎ�Z�`�^���f�ʶ��u�7(��[}#d�Vd�y�˞4�3�L��\^q��3��4�|�X��Rz�����+ڼP\�@�Ѳ̎�)-�e����k������+m�㚺�^d�T����Q�-Q���}�f<I_̊�'틆�H����;;+�A��������ʏ����f�%��sb��>�j�:2�a���-$ �VrW���n_(|Ϋ�c׾��Z��F���#����]F�o�mJ˙�X��ʇ	,�s˫k�.��15��]j�y���j8�'Ϊ|*Ŗ�uu
�<�0Ql�d�u�gnQw���g��I��c��{��	W�6��YXf�T�%"�"3�_�Gl�^"�ְ.�;��n�Um;Ɍv0�J�^�Y�s"��q��w���c"��@��jb�;8������p��Y�@��2�Gm`���֜�5m�̶�>�ʒAYL��r�%`�7Bs�������<�2Q��z�O4S}/��O���
�h�P����\T�
=)m��A��W��|$�)��ֺ�����M��8�s'�T�dq��d@��}6Rre�+���9���жUg՚��.�-k�n����>[���i��[���5c�hM�����v�Ke�i��a�ӑJ��*�]LX������nn�i�W8��H�I�k*K��#�#��������a�l��TX}��¨����l�3\+O]v[8��A_u�]Ә������ńi����ZX�~�Y �^*��{�9˥>e�����λZ�Y�u�He��CF#Ŋ�\����f8S,Nc.Ve�*�g�Q͏r�ΝO9��S62�����9�{�FZ���b	�NH�x��b�I���}ңԳژܓ<)bݳd��4,��y��{p�N���k.��p=��/�:�ŧ���w�4�ʐ�����^Y��O�_{��ip)�C��o���.�]����6�v�^�ejJu��ˉѐ���0W8s7/JH��j�t��jd��$]\��7,����0�q��sU�C�\&�M�_�WMj2���yq���5�ٚ�1[���+��ifc�&�'�ם�A�?K��ּ0	|�fm+�8F��5.�깃w|xo��B�1{�=�nn����<֋8i�\���@����wc��=��z�����Q1��% E��bF��BE�f%���&a����)0���ˠؖ��"IH�̗.Eː��틖��q�����Ȯt�"@ŤR��;rs��5	wp��HPN�I�1�s�r��h�q�r��!�&&%�ֹ�L��)����˝�I�����r�B3	����LQ9s� �s�3f� &����\��Δ	2c�黹���Jw\�I-����]�(@2���Fw]�30.[v`d���M0s��%�dMA �$L��ۈEr�`@��0b)�f#wWIL�J#K%��':�L���2!"wr;�i�:��b�#E�lDLFD��;��A����ί���%��]vw^�V{�N�s����}�R���&�C�Ѷ[
���R�v�'7	��dvV�]�V���wa2p��`m^�C�7�1c;&�Ǐ3Y�����%,s>��LWo��F�B���x��h�C�-D�K��[��sL7���8ת��Q�H���P���<)�Gg�F�ͪ��u>t�Q���s�/��1�ko�}��'\�\�::K��Qg��-4�g�5/v�&��x����?j�f�Ӵ�?��{�wZ�r;�H3�mU������c��[>�v�Xi����8�Y���T ����N�=.x<�Mg��]�:I����׶�xހ)�v/1��sNē�\Qa5�!�[�F8��z1�-����|�+����o'�o�ԍy����xy�&dz���n*eg��}�m�|Ԗ�|��Z^tǣn�{�z�����͜��Ʈ�8fp���v$�:`Hs�n���}�r��O��7�<5�>��ȼ���Q2��q�W#.���͂Ψ#����6~	TΉ���n:ЍV�f�w�l�l�ދ恝��a����'9��n�v��v̅32�}��$�y�Дu�fG�ba��m�-�t0��-�lm���^nM���w���&s��ཧ9sM0�C�Pڲ�u'w}:�\y]��!o�dي�i��Td��^b��0%��r{���xwQƺc�{/��Usw�p;����>���I�5o�B���>��쮌;�uu���x��Y�9�"[�����&�U4��L�����Vg�]W��[��͌�Sr��W���ݽdEGv��q�S%�,>�n<C~����~�po�X�w���l/9%Qpz�*w��I�}W�Xk5���%WEaaW|ݰ4�� �,�[r�N��rwD�ν'/�hn�9>
�Va����xW�}�~�^�wz}] �� �i�W����Vy�i��#�5��ƠNP�#+!X?�l{3�ce}&��a���+�����&ӫ�@T���8��Ƚ�b���o��4ϣ�H98O��2p����NL�wM�W�������]v<ֽ�1�Ҹ	:�=�sL�g���^<ˡh #+�~��ZԻ����Y�חP��򽃛h�\_�x5e0&;�"���D�l�:��>��c^���g����XuJ��������x�2�Ҫ�,��`eC���\��?R�N�F_<��F#��E{��+
���%��m�@�\�ƌ�:�/M�Q�Ƕe�ѥ�TyHE?|��})��� �����x�A�$�Q5����'NCN&��뮉�8��R��9� ���!ݹ�y��1v��v�����IN��׵a܏�:�7�w����������z��.pL���e�o�v�j�Ѿ��C��Wٲ{�]�5o��i��rƓ���z�C3>�σ;n,Օ?_�(�z���!����S<b�]o}ޚ�W���9��<�F���"��N��iA�-.�[�5�_�l�J7������ZSS<�EZ��{�7cd6=�
�{�ěU������#�Cʃ�n�^�,ڂ*�1��))o5��9�AM�˯W�Ͻ����5�8�W�]\�Hcn�Ix�'�N�}Mn#���l�M�wQ�1�O�NN�:�� ^�2|�/|&�vo�A&�\�/�σ&�u�\�?D��s�[�7�9�T���ܗ2N�$a���tn�ӗ0���	.�'�7\�ucQy���17Y޻�z7x�73���խ�j�rGK���K��T�Ϩ��5�-�.��鸷��W�s7ݣWQ�N>�h�j�����eC�>"��^�|nX돆υD���r�x���G{�%�ݺ�`t���<�v"��qNM�*�n�e���+\�z0���e`W-�k�ek�=?S�9��@�<�������ޥ��-t�y4�g���6�e׏�^X~�_�V�}��~���ɵe*�A�VlO� "��w������>��M�K�r�
�Q�"'����+���<4+�Tt{8>��Xm3k+Ev�6i6�ma��T��v]ggE7�b-gy�΄l�_A�͏�F�l>�%��5'��&��t�
0�\���9�s=��y�����ʆ&=omGU+�}ʟ9������ׅ�	�]�PlW;�6O;���n#Jɭpf�|za��W����O ;���<��Tƾ���r��D����m�]5�:�ud�<��_'��vt��t���*�~*���ι�����l˫g!a��q�WM^q<q�w�K<�5>�â���(t�{�}1q�#]�L�F�;���/GC�r<si�~βʣ�n[=�u.W�����5ă��l��u=\�sR_�UN�eB�T�3�s�IU�.�'��N#�<=���B9�ڸz��B؁�S�㎒z�΁�xkd����\󢲵ʚ0�}>F�e�^^^�B�'x9��'�Yۇ��p��۸~�o�E${~�Mѻz{��|1��f6�͠*�f�(��_^�q7�{��
�>;��f�x�Fp�{�}�$���&�V	qj�M���IGt���Ⱥ�Z{6alBN�>�3�Z>7坳3�j}����7���)��|�J�.�;�R��G�sGܧā�~Z���3٢a|��x$��u������~���Wz:m�M���鵕�k�ĽW!3油�XcY����$�}��Lw1̩)�\1��h�0�:d�zg�s�$�����^�5��n ���|�y�����K��=;5��ڙ�C�p��ޔ���v��49��=/�=�cw�̵���Y,���̕�k�Su�jW�����C\�忋l)��Ge��$�\�u��ޮ{����.���;"ӗ�
�!�4@�s�:7�P��Ԧ�!��7��6qң������.{^Lzw�1��wB�c��[,�w��|2�s�2z3��Uϩ�։;[E_��p��%u.��E�ﶸ`����k��е�f�ά)��CsCO��4�k���sF�S�O;���������ps*�XȒ�O���5�z��t̼)5����{j�f�
�����VI�t���Z|\�S�9G�"��@���:�����;��)x�ة'��j�o'1�p��gީѽ�p�1PΎ؊�G�)����`�� 'ז���>x�w�w���i��w��|�������	ε�c �M~]aI@W��Zw�jg��.�C;c&��aW W�;bS�Ϊu��SY�.Yt."��w{��ѰQ��=���6<�壋����p�����C���� �����ϼ�;�U��d���f�C'�}�=�	��8�zXv�GNgb�B�h'NK5�|������67mcZ+���{9 ���޶s���0�aJ6b ��z�|��l#�����\�:�YI���_��3�s��#��)q-Ӓ��S�P-��e�0qe�^b�K[�}�M��c<;��#�E���#� � ?U�t& ��;�3�d�9��z`���:Ԗ�}��!i�~Z/*�W�{]8m�z�S�^_���Z RF���=�����}������2���p��+�Ӈ��!�u�x�G�8X�F\S�F��,ڂ8��fU��tM��r�����Rr3Р�����N�1��m�79���'7�wlȸ�UR��u|$��f����5�g��>�w���N0a�{,�����,�d�7Q�+���%I�G�!ns�B7���N�}���k�s'h���&���6���uC{���,~͌�?}�#�YP��w���U��Kd�2K�gn����$�}W�Xj#5��]�d���`iuծcEޓ3yiΚ�$-�p7���@4��9>
��a�+�x�ݗ���w�S|y�Jwۋ�*$K3����L���`*/�s��U#���c�0�Z�Z����/��Da�O����Χ��Y��Ƿ���O�4�ǾM�s/fX���%��f��w�'	�; dਓ�	�Q�������::�yL殭���.~밞�Mz��>��LBa�%������7�������5���Q�����~�Xb��68ܱE=�R���1��!��4��9)��ͧ��o�n�X^��͝�5ϲlgG�:۔��ÝLU�o5�<gݻ�	ǒ�����p��Ԯ��L�.u~���6vς+⑙|.�X�7�{X�����:������@Lv+�E�>~�T�s�φi]���Ʋ돶1?`!�z�M���c�����6�����B��U�Q����`��
��\�ӹAꈧ|4m�b�@�Z��,����UK���r�?\�'�DI\h��+�/���ߖ�0�]�B)�o���NF����L�υ,��eG:£��2��J&e�`>�ROt�ES�G��H�`��8~�s'#3<��l���He��=���&��My���(�.�
�3�L���1�=~��ׯ�|�k)X~��ΰIN��߹��5�ö�'�fD�K6��ʠ΁���Wr<*�z���Ҷ����]��P����z �;��n�<w��ڸ��nh�����G�;n#����5�N��`�+�{
~��ڎ��_�5h{�����;ۭ��SԎT���+���7~��kT��� >��uO�;�	%���&�i�k�,GT��Əj��a`��h�~�q|D�Y�m��n����x�u�����u�� ϡZ�v[/�Nd7۹���|�1zna�S��,� t]�^�e� ���7�-C�#�Ù����c���&����G
W)�u�΅i\�T(��
ND�[�j��Lq%t�ٱR����|r��f�P��GO����M���Z��i�M	�_��)�Q���O��cg���|2):�J�ܵd�V^��oO�s���.;o����y8�&�p�s�q��Y�@Ʌ���������oT����4|%Әxy�]�!��{���AԼ4�f�qZy��Vs\�sq�53�VzZ���C�;��lK�
����9�r�)+����W��9S�>�\�s��'���ɵ��8�ζ�M�L��'	̳1�4^T+�Ua�<���) '����UȔJ�5���������E��3��x*�t/�5��^,����S��ˉ��Fv���Ua�*�qT��	=���Qs�k����/�x�:��;��'�B�ƫ(���O��C�&t+����.����{���t���Þ��U@����.��9l����Ч�v!9Zi�_I��,u@3�|���N@B.m��^���e*�?��S�/M�:b�}�1��t��jtuHy��ߜ��{�=Q�0�賽>d���>Θ*[�F�'V��_�����sd#	�gD]����
yQ��ɾ+<6g����C�h*(a�� x�!�B$�>ul��k���z�ϰ��8E�_p�hX���C�c�ܼ5�1��J��\�&��Z���� ?�VtI)���P�_��I�s�h�{E����p�Cv���^�
��%�ߋ��Y��L][�C*U�j���#$�ÑZ�Ĕ��t�|w!:4�rcK�w�uw�*Y'��"�u�	��*m)��H�%*�_@�L�	�����ۛ5<1����;���%F��i�B��.!'r2�ճ7�(_T��pH#�p��������8��{F�70�f@�zÌq������,�m��!���u�d_ʪ��\�f��B���^�U�W���~��9�O�Y��z�V�]ы�I�e��y�#Q�M�����Ѹ�|+t�r����Z�-R�T`ﺼWK�W,ev��ǾI]�X�:��nX���a��*u\A�v.�n��緽޻,ɷ�\	�ۊ��7E�{���z����uz}��f�ά)�9����n'���q���"s�F(ˑ{�	��q��P���s�+	�xy����"O�?V��������l��y|��[ڮ�r�5����X>>������+�Zn(�'�P7�&���[b�\o���T"���[��}��KwZ��R9�z�HKȽ�:����nlk�Q#y֥�ƭot}��1m;.^�����g�u�V,�]��7���#xP�{
\3�J!C8w9.)|m`�_���GLˌ9H|�n�{�ɹm������v�#���v�2�s�ʚ�ǡӭE���շ��c�ʝ�d�9L��x+���#������繬��+�;���>�=*��
%;L�|���N�^5�\}g��Y�=W#�=��.]���5�jd�q�7�3�&��Fp}�\��d?Sg���g�ca5�\i�ٹ�b&�[�����w=����f3MT��T��,��am�Az4�~�Kg=��}��M�h���f�~�^��(�q�OQ����
A@��"���k�w[gϤ�:k�{
Y�^9�'�$L�ilT�����F� ���R S�'@��a�F�(�ϡye�O���Sg��B�~�Ʃ��t�+�}�a���qN��g��j�d�	T�xU�����^�Mվ����[���R�N�1��m��nwIx�m?�~(J�mxʮ�����g�ͳlao��a�/j���>��ﲈ]ʸp9}e�9�d��۸���&�U4�}Q��lĒu��6��� C�ݥF���ܚ�Ʌ?nm��yI�i+�(�������ֵ���mkZ��U��m���Zֶݶ��m�⭭km�Z�����;kZ���*�ֶ��U��m���Zֶ��U��m��Vֵ�����m�mkZ�������*�ֶ��Vֵ����Vտ�kU��֭�km�mk[o�յ�m�j�ֶ������)����K��f/�9,����������0ʟ|��JB($�(QTH�@T	"AB������ 
"*,�  3�J�D�$DEJ�J��	RP���JT�B*TJ��D�����TUT����Q*�!J�%�Q���T�(�U IJ\������xӰ��Gh��n�R�k��j��n�Ht���%�;[G]��v�t�լWop�UK� J�[� ��+���٭�u��9�   Z`   ���   X�   f   ov������<vUsm�J�$*�UUF� ƣ�m�3��5�5ݷd�R�f�v�YN#UUۨ�%Ԧ9����kJ�;�&հeI
H9d
�V� s׳ր���]��m��'@`J�ڠ�VSUN�]Z�åu��alز�"kc-�����*�,!M7UIIV� �U��g6�S�Z����5X��ʪ�[kke��]k��,5�*���U-���7Y-���ҚmT��)ͨ�M� ��t+�'�P1ԗr�[����V�k�A���a�u�n�:s�����
V�;:Ll@��BB���*< f�L��v�v�հ]�ww]�jZ�j����ۭ]�9�m��Φ�m-Umk��C�WgZ���ɻw%*Uq�*ISx w=��:j���WSmf��Ssq�� u�f��3��1)�U]�t:,[k:�wf��\
��$*8�%� f��h�,�ۻkt�uw5s��UmJ,wa�:;�Z�訹wc�6����9��T����@�� 3�P�nGKN��˲��![nᎻ�e9p�]k��uR��rۮ��T�N�S���      �x��U)QCbh�0#&�b`��OhaJRJ� �hd� i�i��&�&	��0`��E?LF����#M ��M��~$�UJ���1  M� MHRF��d4@����z�f������$�C�/ޫ�h���Y�������V���+7ʱ�m�g��@ ���^~2BHHC�?蒤�H ��$�,��'�KI!!I�������?Ώ����xAQA$�	!!! p!� �$!����]��0 $�2���^~��0�?������$$$!����,-�X-���*!s�A���3�PO��<�-

*	~����������n�`Qy�fm�-�l&���gQ&�
�reeƊ�t�P�"��,��ZLK5�Y��R�f=b�:��R+j��E���i������Gk�ET7�����B��q���:�G�UelWeʽ�zܛ��M����2`�b�uۥb���i|�h;�(�4^RгuYI��ٴj�1��3e]�v?��]HeC������l�n͹�*K[`�%^=TZ$:ߋ�ܼ[=���$^nRM",�
�Ի/m�i�i���ֈ�r�/]<Y�M��I�?)�u�YxB8�o/>��Oagq�U�Ѻ����(3Q'1�`��V��e��xwS�)����5�W'`�
�[�6��\�Z��H�,�����/cH�R�l�3w$QV�� ͡f�J�ӛE�$6ij��w�M��� 귺�|w��hYD��L�E���9�����T�7*༣r��e��0↷>;S^ɉ�sB�B����U��0m�����h������/6﹋V�2���Vq%B����9�p��W�)�{��(=f����|3�b���:����PͰ4(�1^��iɱ�hV
"�J�cA����7ZUpX�g�9���1L�j��r [R��MԬӅ�7�iX���2�q]="۷���cx9�ub��K�H_Ìt�+q��Zj���mE��\��a�C��Y9��e��� �����r���[$,�!��a̙I;ʕ"����"�M�*��x�̤.�Ԙ������id�Ձi��GN��e�EZ�
��ˢ��O/��huz5����ݠ�5����)b�(�K�e���]l�v��F����'���'���L�K�u]�CbY%:p([f�T��hА��h�,�Gh�Z�5f!φ�%�k6�cs�J�%�PU�-m��`9R�D�tl��i*�f�eϮ�/
\O�;3��'H�/F�zp�JX���V�\'p;��ubx��0�5���7/n |��U8捌��V1FdPj'F��x�бa��V�J��*��A��-ٷ�U�ZBPR�V�qk2�u����;,��v~ۡC_�U��T�B5d$�G*k�v�<SRe�k�ʒ��	��y�Y�+.��ڒ��L�W��k� ]����:���/�&����;��T<,��t���6"YB���ɦ«�n[2�"�r�J�[�d�f�%�XS�s) �w��٫D���j�����8v��O�JZ��`�S��Gԃp�yw,ޫ��;"�%�0��FX8UkBɳ5n�2�)4�	�"��HU�]
�T�P!^ؽަw����Gb+�K���u��t�*�!�$�0��:W�H��6�H�p]�k���x�:��H#��쳴�iX�$�K�ʎ��ysL�p��4��AK՛hkѕ35^��
��_^�5^>����dR��n�����q�[tXwXL(�^�d��ͪuq���PGt�[�K0!CkL���IE;��p�[�i	h��9t�k
ݲ{P�7����1mo?�k{-�bP�RkN�Ln���zu� ^:)XC1�W���� ��ʎf�4F杧n2��^�i�Ԁ�0:�6�a�[n�74�z�Z��n2�j٘���*и��b��ʋ�m5��������`��,�v�܉;ǂ�]iR_g(Ew�N+I��^��S�z�]k�)�,]�G4�U��mS�����zs/k�XkHM]^��f�WLK�	t�f�f�]�w��	[V�Ws6�_5�n���ڽ��Iզ�סb�![D�ŠZYt��i�%2�@��t��)3w�E��M�q]�H�8ι�_ڪΫ�n��)E%*��J� �bx����kT�OFޓS��Z���nn�]��	| �۽Z���F���e]^SHI�vhL:�nk�z�1����L,����4e�˥�0�ܥ��|+XyP�[�F* ��8���	�n��V�Zɦ�C{5Y�ݸ!���Ѥ	�*gh�X�v�y)urࢷSMiQ�rMX&\{P�5z�y�����O5�T1���vU�8^��ƶt�ɔ�=��X'6�M
9�,u�ǃ�l�PH�qm ��T���M�[�AJ�^��7��dk)AV f|���bo�wa�YA�C��n�kJ��4��HbK2�e��+��� ��`v-t������}�
��50�=D"�d����	�x~*+��Kqp9"�n���і� ��k�i{|������'^7�(n0A/�Y�UV%ރ�s&:N^<�S�Z�2쨮�V�f���`�1B��R�C#�Dۭ&���K4�:�T�K6�gi��M���9Ef[̓e$@<I%`N�I��������-�V��Ŕ�b6E��o���d���>Ё�j�Q"�ܻ�@^ u�g3n���ŷw�ބ���d"����Z�F�"���-K7�@�RF�ԦO�%��.��E:��OlD1�yv76|�m+�[�F�.S���8!9�QF}a��`B��5+7�� n��Y�t���8n���+af*Ӵ����%�2����������(87l�9{��W�a�a�b�0�������</��ϏG��U�Ԏ����lj��A`*-P���lZK��]'�1� �D!��U46�⊞fDw ��ơx��VcAl.��41,7�����Iy�������)�=LX��t�GF��[;�U+	��RM�,=�ve�r��xn�k@daQ��`�m��.ע(]��AYH]襡�ecRY��FkJ�1E�oEk�PT{jm�/X��H9&$����K��.Eq�����ɹ�k-p�K�J��G�c,�N-D�ϗ��/�e]%D�q���;��	`Z7r�@UF�Y�op�j.�]��)��$p�t*x��R�e���h=DY�t�J�XAV�Z����ll�Y4�H���ﺬ=/z�7�pCR����cT�
����dfj��-6E��<&�"�oUd�u{��lV(� xG.���RU�ø����Z0K��GNn��r@C9:lkxq�2�NdT����lrU�1�̭����dY���]����,�k�z�fO�[��m�1�lL��Dd���۫�A�	��J ���<]0E^k`�Sgד7�����:^Y���\u{��o3q������ߝ�B����Z�V	��J�xI�?���w��2� k.<#^ҥ�����J�=�V�T4�(e-�Ĵ��0����r�`3oH�`a����e�X+i�@&�j=��Wq�}I����S&�²HҨ�9�q�I"V��h/�F��.�2�����ͭ��n�u�ur;��YEh	*�|q|�D�m�s �ukS(�Qڿ�[VѥpΪuJGY�2.��B[�b���7�;Q�4��(��[3]&ڨ��VQn��b�������\k��Pwu����,�#&�&��R�30H�`�{Y���*k԰��6Z�E����Q3unC7j�Xmn�Ae�jG2s����U�Ic����u�N|X͛v�Non<��ڬuw��Ԙ�nj2�]ҟ5�,kY��Xa�7�`�k9Ş�F�����Q�՛�q:����u�L�۫��B�'ux.�]�\*�)K��5l�Ĕ�Q7)���Q�XY?g���Ŗ���k�8-K��2�uB�,,g+	�nY[��` C�Ek1�سh��]KZ��U��X�t�Aw��!�H�4,�\"x�c���d0���զ�{�ըi��n�m��ODGmlp�*f�;6�f���(h�0e�j;��,]J(�nZ��$���+1�Y̊������O6k���3u�X�^�XM�%�V�T]��1��������UvAi�z��"BL�,R��}��ӹa;xsqٶ5�.�����t�5+�t�G6�T���Y��R�K+$,���ICGS�.=�#��R����A�)-D�]\Jc�̰�Եt+dT�r�X�TM��Q�*WyyX�d࣪���ܬ�ۼ�|I��X7"i�
(3P����{��0Eڰ�.�"$�ٚ���"#3ED�T���6�2j��E��j�5���ʨͅ��8�,e��G�-���4�&�WKjG�#���֦��؆��b��լ��~xB���eh�䛷j��&4T�`��]=����j�RR9,��v�V���M��M��W ��Nұ9`Pu�\;}��m��s=�R#R���� �|�m^%�P��^��kV���/��3��D�!
��gA����P��(B�æ���"�Ʋ�͘[��E�J}�6��-5a�Э��P�X��׵[�U�A:�ͺ@�bC�uyOZ�R���n���]��4��W'�����!(_ŃC�������-K��J�/��ëy�(�9h�@��h�&��u��ay��Iٓ��K��/9�w�h�:���?c?MT�����m�Q�$e�ڇ�|�v��T@MUC����VM�_U�A�}���"��          ���8Z��i���U�l͊ήPW�t                                                                           ?�  0                                                                                                                                                              `  �w������F�b��J��'oY�yeVӜ��3]اL��}����f�>�!is���纞���P��<�غ>���Q�6�f=n�a�v)S�{w.2*�哘�X��[�[�`s��6�wr�D�����W,(W]|70ܗ���k���D���[N�C��D�a�`���j��u��s$L���0��q���Y*�Ή��/��
�&6�o�t�
�V�D�jc{x��Ηz�TЫ(�J�C��<	�|C�p��u�n�˾zg��f�tn�tY=�P�X���[�u�<�v��xI`�� .-�{\U�*���n�!_�܈�u�A�'����ɸ�s�F��h����l���x�(��S�B�D��\�;����7v��)���;�%�4DbN˗)gwK}��3͂������2����ю� Z9>ЁhoS*gY���mCꥭ�|��][<1L��A=�&��`�[C!w���>(`ݥ�\4��ŵ�{7�pJ�I	�3iL�-dc�nեX�hƳ3��*�r�M��X/kT��]y/E[a���37��!�I��k6i{�r&i�H%Dn�f;@���/:tg6֥qD�����u�@Y�;�at�t��^B��b�N�U�`��J�ʽ�]��(7�uV�|�%�^���sЮ���b�*/��GyL�{��c�݇���ulrQP���eY����VX3ː����7r�QQ=���M	tt34B=�X�7�n�E�Er:v:ġ�T5Ǔ�s�<���[Q�$�V���"h���4N�˕����n�>/t�6�T�W�W,�o]s��=���*���Z@�\]x8J�i�sWƐW�&Ճ�>%��D,�JH6�T�_jx�W
�}�4��F�kZ�!Mݗ�V�;)u�)Z�rU�:�� ����m�t�wCx-�݆�3r���|4�ٴr���q3�u%�2�M��R�Y��e[����lI��-aU��i	�ah,�P�]ܑ�q��]��W�b�u�d�� 姱nGv+K5�Np"��,q�/�L�����<�;m�-ї05��Ӱ�c_ٕ��*�G!1����ss��4�"�`��X�OjF�Y-�9;*;��f�*�p�Gg%]a��:��J`�ɓ�\\I*h��:��Zo�YFgLDӺW#W��t��:�
�k]`u��3�2к	��%7�)wm���s���A�,�7h�Ez�Rы��6~M.�_z��1}�^@ӫZ�@�Ѽ˜.�	�N�#�SD&��R�W�`<2�Q=�����g��S�D9ZF&cGf��u�d{��L	n��k/�m,�0a��#P�X�É���q7��}y��XT,Y�w�n:�>ނ�P���[�BK/��0�<��^]B��9X;d	Lv��(�rUʇ^��X�:�'�e&�F쓺�I��>x��.��E.��;D���$]u�<v���m����W5��GN5���O)ד��=ధ����.,��N�$�kd�^|���"p͕�.��W$�v��R�kFU摗EV�ek��5d�
R�9�gA�1;S�
�bABN��Lu��P��'V�Wg�X�_4�Hg4��9��6쁜Cvv�����oPmгs>l�nY��l�bk�YoxiH��mI�,�C�Ќ}$F�����&�
WK�ӥ]�\4�G�A��X�Qv����pw��U�n�m�W^�˥�Qnxu^�K:���إ8-�һr��-j̹��^W~�K�>�~�*.W����(ޑ�Ó��bp�����ͫ4�|6�m�ԃY�q�����y�,7( ��|ˣ��R�6��8P�;<�nw�PROMv2��!���|ʝֲ���fQYQrl��Y�5V�����:3�2hmk,��;%��V>���!_&�!�v-s��@��u���YB�>ɻ�9Z���ݬ�*]L�>�A��Eu��,f��|y<��`�eb��I�2ﹻ�d��Ȟ�+8����*�-�y�w���b��w��p4SUH�Y�ۅ`�I%
�Y;�K��;Rζ.d����5D��lȯr���-���:OU����Pr��yj|�4֕ݫ [�+�IsV�x��.1gl�Vh *�X�+-%Gr'G���[P���Q�	��14��)SF�=�2�N&��E��׷�6��K���nÄ̴�{w�7�*\� '�q;�mP�v�Y3{��o���#J�F�����޼,��8���%M��[ѵ���K7]�eE[�U�b���%'G�YXs�}�w,Q�^���9$��tk\� 3��2�C����]،-��Ԉ�oIxN�/�E�K��6�m�!q����
��Y�"�ᒷ*T�t�� ��Eˤĩ�Y�֤�S�먲����k,v�ޱ9�i���:y[t�;�)\��@��S��6�=� m
�j9�ɇ;;���ϢD�'�α��h��g-�ts����2p~�N�7M�ݰ@چ�jFɘ+�Zf��ثo���4&\�&��ӎa�F�PN�oY��=�0e�Y�˥&eX�tP$�]ķ;�
��K�+U2��*̭�.B�J=��'3e� �qQ�+�U%��6��u�Y[r�E�v�1�r�`8�J@46�[T��Μч�*�3�+vn>:��m���	�ML=�.�
�r�s��<o�[�<lҹ�if��#]Cku6��A�B�$�UF.�;t�5��@N�C�9���@�A���1<�ee�97�0-��� �9�"4�`�I���nݴ��갡�a��d����7t�B@�es������1RiCg,o!g���՝�F����̐1��}�9_��;F_[�D���;���*\�@x�nHvm	��`�ws)�jPN�ND{n�.L�[�� f�'9�-�8n��%��� /Cg;s;aODu��u2�Q9��l����*H�mƥ�`�Oً�ΞcGSv��i�V�0�b�@!����,��a�ҍ�9+����k��d�������\.����R�����[0����Vw[�Þc�̑�&^���x����/�K�.,3R�%.�����q��oJ�(5j�C���"��-W_�[Y�-�s9,�m�m��)��B���6]��ô^�p!�
��y�0i��U՞��u6eM�)]�ֈ��-�9��]�2��h��fT�x}��-��'�9�^��Y�:F�&y�>�,���9�ye�w��JTY�@��T��p��]Q�����]�&�o�7��rp�c4ƛ�2�L�s��&2R��]�xNWy�%�j.���.��婩�J&��;~X����r�>}*ʦ�\����,���B�K�ȦEu`�B=�i��t��I4�+^�r����Z��r�P"�tۃs8�u�h)i*ɘ�:�*�ʳ���,w��Sx��mL�Ca&']��6�����`G��݇��� ү��7���H5���W��ʸ� wH����Y�]�!�\)��)�L��#0خ�`V"U���b�ո��~w2��z;ؓP
2:�`�z�)kt{H7�h�X��o ��uvwݠ�P�\/��'��Cn#:�0��A� B�i�`B�K�
z�'�3O�ĥl�t�r���u5G�f +�'�Út�	�~SB�I�w2Ŵ]��7+1�e&��q�τ޽���7&=l����1p���'0'eZ6�� m� 6��ޭ֧��n���U�U.����񟆌��A�y�wܨ�oDN+�0٘���;�r�.����j�vq��V�(�e�D��9K|�6��p�3с���9b�6�y;�/�Mik��%�S�vjl���"cx�fi����# ��d�ʻs!�N1�;�렠	h��d�,����ͭ����-�߂��O��j�v���lI��Ķ|������p㣒�p����vk��Q�\5 �$�_�5_T,J��QU���J��yVL���J�WY��߰C.^�=*��ͷ�k��W02�͂���:��[���M}������YT��4eY�*�JRJY�E+{cb�7Q��4K2���\x���^�xyX���d�`�Q��:���Y�\ƺ�v��y��T�)� �F�٨RG,�'d��x������Q��KMCv4�'�4�s�e�b���\Bnm��>�b�"���>�X�ٹ��^%;_K���Mz#2Ȩ;�*�v]M+E������Pm\;�v�Mr�"���E���L��R�Fu��s6P��P�Qm�h�+��jne��2i�ރ�\�� 2�}m��*n�Ӕ��B�I�., J�.��5ʐ�׭V��\��dճj�di}���2��˛��K�@w%���             ,��EnNO�ll)S-t� U���#����h�H�!K�Qw���c�*;�^��2s��A%�;������o   �@�@            ��7�_���'�>�����ƾL�I	!!�L^ݾ ��W,I	���>�~�I	~���~������!����g�=y^��`��Ջ4��I�s���@�y2���ɷ�:�H�ܭ��wq�0�G�0��3�a&U.r�bu0��鴞�
����.��>K��c+�+A��*ťyWd��c���1����J�n��8L\��0z]��EeG-RE�wJ�jm�۲'�����X���T.�/3^vX0��B�=wI)Q�W]�^�E��l��L�V>�	���Q�3)�kWijj,�R��c�
��P7*.����"���m����"��V�]�(��}z�7�se�y,w�B��:��u����ӻ�{A�=f���9�-\��B�v�Nf���9��L������'��;g����ɳ��:e9B�me�=����kqD�{*�gdlWm3�JQ�k��\6r�������4dx����.�IC�λ��6��!>�KE�m�k���^��5m�׶��hu�D�k�L��ft��eA|��L Г,�<�f��pl�����Q��3��@F{�ر��
�c�j�9��Wu;6���Vw��QP�� &9���y1e�K�e�s:Q���*�0GzR;�dlEȮ�.��S�DmJ��::�=hv S�pG]N���V�����9[+�h�),/�W����kVWi�qn��z�\�i++�L5���Na*9ڹ���� ��0��	)�>��;�La�U�3_Sf���S�:�d�PZ(��uH���J�_'!�P�wc:D������H^V���7w��Y�N𳍣2V��wn�e�Q�K3��td�J �n�Ԕv����3X����T��v���aU���� t��˵���]YlLT�l�f�7*۱���J�<=1m�I��Gu�}��V���D]������rPC���@f�>�z�x�f�p6N��b٭�)� �e��vmf��\3��Ѣ�E�7��T!OY�X�P����֌�@ep�����R��V=��h�@MZ�%�1Z�Di�x���+N�W<�n�YT��i�+��#�3/9k�-����M�ȗc�Q��F�XK�;9�т��¯f��p@_C�r���gP�s�Yd�ݔ�V71>Ob�+L׌��1:'
XD��m�8�]@���HlFuj̭�B3��w�+�:<�08@�Q<�JJ�e�y$�u9�3!t��`�Ҳ�ݹg�rVܝ�����Vl1n,|�.Y�6x�ig�.:WX�nьu'f�wW���i�׋6:����J6g8�@��^}�^�:�=۵��DM�Rh��t��a.<}�Fյ�p���%h�`���X`
��``KN�����:�ݝmvW�������A+�*2d��o�h1��H,��XM�W{ϛ=4h/��H#X+��]�mVK>��;�������v�׬0��m]�ñxv-�0V�i>eP��;��أ�U�O��cAC�%aYh�K!�����^���V��D�%�
�M�ڝ�z�Z���1nٜ��
��I�/W�)���[\i\f`�D��J��\�vE��[\^�a�Οu��9zn�1-ɛ�.L�ܡ���A�2�w[���
�Y�k:�X���L��k��}/
��mnf�K��L.��WC��b��m+��1�L�F`��nQJ��9whbn�HH�ʺ}|NIҵn��P�lS�ھK-�l�~̵s/&�7.:� ���i�z�� ��u7ih�pd.�r��zu��l��yb�">�x�˴�N�,Z�&�Wn���y�w$����a��/*P�i���Ϫ�ֵ�]м����]���S�T��ɴjCu\�+�G�n���Q�{K;2�f
YG��k����:CX%.v�j߂�A�(^W�+8@�\�rb�C���j��_>5Ơّ�� �6�GkuM7�/��vL���c�;��tm���S�����CXx�萴D���֘�:�%�iBk��6�I2���)�ө]�^v�L�f��@�"�,I�
�ʌ�K�)�n��3h+˧�(zv֮y����Nq
u�8n��]:t���S ��X&]j����Bc�7R�[��ݹ�La�*��P�ޥ���!i�ԑ{��;��v
h]�U}F�㵲ͧ�[r��B,Үc��[�3�1.�`Zu���&�bHU��Zp=�j�/5����ּҹ�T������R��g-��ύ��K0�K�ٍD����z��� n0p$��œ4��,����r�y�Zΰ�#p�nq�1K��X;%�t�RI��.�jBqQx1̲{��&H��.�^,Vnڲ��~*`����d(ͫ�3A��tF�_SS�mŰ��;jsYD�2��"���b��ٽ��R�![_Cp�JU��9�����5-����f��Q�ZwJ�P���4\�Z�v�����O��`�7��{ngZ�iU�$7���.�ⴕ]}D���Pŭ,,�7�b�l�׻bG�{�� e�F��O.�;z���"��j*�:�<�yv�eذ�;��E���7�����L]Jv*���{6����V٠S��3F�ޢ��4Vni�޽��T�D�Ԗ�2�mq��)�Vz;Y22엕��kn����v[�P�� 2Z�ʐ��bWm�H	�P	�v:ɜr���t/�4������d��LC�z94�g��%�z9ە,�ݧYj��V_q�cϚu�,��i�t6uY���
F�Tx@��YrvV^]����k���=qdv��a��	Iʎ}ҭ�X���8uJ,^�h�W#��,��uz񻣢<��K.Z�Z����A*V$I�YX�:v�R}�m��셹g���r���N3:X[η��ɗK��͡ `��z�2,U[Q�Y��\�㣺���ewJ��*ޑg6��	&����!�ct����:�`FȄ��X��:��הN�e �XV�Y�;�Cl��'���÷�ڒ�[�(3bQ����	��X�pK�m��m�ev�w�,���
��9qX�F����(ӹ���;ح�m���i��J]��sH���S���R��F��p����K�BվE����w��N����j��V��g>|3M����ʡ̋K�G4m٨��R�ZD)��gGD i_�Yd�.��y $	)�8�<���p�w �y�,Z�c���De�>�#e���v�޶�v�d�@ۖx�5t!:r�2�4X�E6�Y�L����Ԅ�+3:�ݛ�Yb �ܧZ+���˫��w���^�:u�v���D��Kh�m�o5f��yEc5mh����z5��IM��
�c�8aw*�ݕx�1յQb��tP�)�{�.q*�h���_jL�[��}ILp�=�f�2-�Le6��:���kn5���#�;7A��;�jُ^U:�KpA�aY�:�P%�v�o�X��V�J����}��pH!9F���J���Λ˃w�p�H^<:`<�4 ���K���J��1LO�3�6���ttp�܁��t�ʨs.�ԝ���� 8�F:��r�a�]@�h��ٳt+X!ε�`�w���GuV��ywxl+��1���f�{�!C%�ԩ�:[*�3{V��nuws���̔R"3{������B���.:φnXl!C&���4;��`�����YDkKY}�m!B�V����c����[
��d�u��i`�u�2K��6`�V�sl�$f_��V��=�P��o@��XU�:ʼ�i{H�6>��[4���{.�wA�;�P�hR�B��l7E@�i�EU��K9��#H.˖���o���[��Z��� �]�v�-�])�-�P �Ѯ��uR8�NT:P]v��6ڀP�������z"I���C�\�\���%�� �k��֘mw���\>��{;^L��<k��X#��HO�:�{3�C@D[�W3B����v�:Pl���ђ�v-�e��s9��̆�C�\��aoFf����;��Vb�M�5��.V*�m5J�t�^��$��&��S��Y�ڣH�Z�}� �Q�����X#�*Ɲv3��2VݒFqZ�,��uT�U�:�˸~[՘�)�p��/�q�(���5/[<�]H����̸'Ff�V���"vB3��������J�uN4�F�&4Jsm��H�l�鏰ewf;��K��Q�d�6h&��{�E(0����bν7��f�����L�Ylo���U�Z��yk�%Oy�V���E�>��nX�ǧ�B5fv��<5`(<�Xy�L���Kq]�9x�5�*XQ��G�亊k�i��5׃�����ZC���t]	�����a���p�N�s�y��gL`���Y��U��W*�b��15�~�xu��W ��zvȩ^A+����(;C�U���	qc���i(%D��^S�vΩ��Ӫ�$��j�/��ӻT�����M��j�m��L�si_�)��W�"HHHAXE��Pi$���!xHO�ŉC ���vJ�k���                     	��^��b�=��t��ݘ1�w�P<5��B-��a�qt�&�f�u�/5�A��v�V�-AV��W6t�l�Ŭ[NKpT��L&h�h�Y��n���Bֹ:�q�
�	=B�)c.�sw1�7�L�>�vB��p����c��>h�u.�����v�S��rp�U3F�-/�q#��ڰ��۸˽2�.Qg��C�l�w-�+!�i^�vl��ms���29���RzqRW�YV�����n������l��[�����s�2���B�:�3�±�u�V�Đjc�ї���t,P��FT�T�u��1�Er�}�)W�j�$�ݑ&]���F��З?�n���3Z��2g���,����zlPG��YS�ǂ�M`s�O�:U�w�듌/�Is&)��÷��u����3844�J�2����:ԡ�ե)%���Y��h�@�E̺��鉟��]��+�x��0��H�E��
E�$X��EX" ԥb�c% ��JAD�锢(�"RR,�,QH�X���,X�PXCuP��*ȲE"٧�)R()"�I��U��)"Ȳ����)"���Q@Y}PK���H��(�H�

DH�i"�"ńPDR)�C�(�dX�,D!d�L���"$���Nb��7��۳Y�o1[s�M��>�ԳIp������a��2� dLǪ=g�������f����'� ee�ش��<n���w�2�6ڟ�ڊtZn	!!|�mv�;'o�x�1��%���+��?r���Nc�5��`w�/A{^��o�;T���`��܇�����Nu��zV뗻�_*�Qܳ��n<&�����7�='�WA\�g�B�^QM.��Ī��V��96�/��\��mO��ի':/2S�M���7Zw���Ec{O��H�]sp�Lí#�35T���{WM^��K���.8��l��-L���N^M�֙սZP�?��z���~���	�~+�p�o�m�}�4�<y��c��1��C���=ˊFg[3�՚PoAq�{oa��A��-d���}��yxp3d�X�������vq��q�va�rJ)	:V{72���G�)�j����X����<b�u� ZSk*�>6O���%Z�&B�s���B���=~쫏 +e:њ/�)s�6�s��G��O{�;�V�q=q8��N��{�w={�!�x��eQ�*�m�g�ݽ�dv�����Na/����/��~�l��Ǹ6{kҹ%=\=^��L#T�nT^�^#^Em},���MF��/�L3�`�?FG�k���5y��C�̫Cٳy6N&�gb\�)�NF\����'�o������=�9�:���ʚ�Ό�GOP[���V��M  ����lP����Dݨ���s:�[r�i9�qd��}�[ʈ�QnMk��g|�#�]G��j�;Hbc5t�	hE�-ԋ�Lg�2���$LgX��3D���ù��X���Sl�D\Y��_���=tO�v��ob�^���
�����<�y���ru+������,��RW��4?z���!z$�L�����{����C�����' ����k�L���ݕ��ԭQ�K�K���%k�S��;Ӄ��~�����=U�،���F����x�g��޸[����S��^����Ѕ��=��8TD�Q<��͝36/d>�a�3�w��2���;Ǿ��K���su)��z1��Б�J��7Y�/"=¼�X��͍���}���Yt�G5{MZӿ薻^�h_]���z�n���nrc���ma���i���V}��{_O`�����3�"MBt�;钉P�4�K���j`s���g�9�Q�Nm��ܙ�kI���R��ߢ�9p�彟R/�9/ݺ�/w���c/��jx*�$�Rƞ�Rv�xec/9Or��������=�׷T�9���Gעf��o5zg��yV�£��FR�B�J^E߲��b�E��è����*�R�{4��p<Hh�-'s�{��n��V��M�[��e�Vv��uߖZOT�/�1�Z�K�I�쎋%�ڴ=ӷ�)9��u��ڳ��k�5=�_�I\Ù�:�z��X{�8uW�{;f�pr0<>���r_{�-��G��`����(i�R�#�����6��|M�w��!��+�]g;�z�Dn���a>���i�4���wu��{W^DQz��Ǿ�OJ\D[�K��2��&I��ށb]����I�B�)$5�B���9g[>��hr���q#�U�{�;�ޯG'q�Θ�sO_c7�1ɽ9�6�=�&��uԽq�L��k6�d�'g70��>����zz��_o�yi�����A8)j5��|�����ژ�r�ٮ���^o�zߖ�{V����Ģ� ڛΏ�X�ɯAC�[��2j袣���E�X#*���Kv�g�o2xp`7~;��>O>p\����đ��W�:��7M�/Z��/�g����iy���JS��-����x�[�6�+� �5��/v��#��<*�$�})��Q��骸��9��&���c��:Un,��jY�ԟM���좺֍�3�@k�k����Q}3�C�#�Kû@� #6v�{A���jWe\ziea�"ۏ�v��2X�|B[ǖ1�)��[ؕ���#����H����Y�oת&������p�z���~*�ļ�����'	=��$�:����|+��zmQa葓d1��/F���˘�4�Ժ�}(}���fQ���L��7fn�Q�0��oyŮ���x�_;�%8GLO,io��w�w2�O����5j:7��ZP�Tׇ-�٭y{̟n8���7���CnK��E�j���窼���$��C��?�.=�{Ƴ�3�Zں�N&�����8}��u�6#Gkx��ݽ��n-��Yz��Su�yt���i����}FD����
��I��1i]�t���8%Y�>3�x= ��Q���F�W�W���×�[tn��Lse�k;n�X�{�7]R�-�f��jŽX�c6��kt\2�l�a�Q�9��o���5�$b�I���7ׂ�fy�y��[���q̡t끵F|��'�MwGnj�9�#6�U�{�\��4�U�S�iL{Lp�G8#�p+𻋻�=E�-�n�|��
�^�^�N�y�}d�v�7Iy�^U���z0�[Q����îN�cΗ��Ͷ�W{��u�*�ϗ���&E�wu=b�&C����&��'<.���2Ξ���6vˆ�6{��~ޕ���;�={yJn���\։&��"�5�9=�\1o����FCQ5����y 4���!Ǵ���x�q���7���R���ƼS_Īev�n9}g%ŷ�7,
�U56���y�!ؘ���Fti�>(�r���,$���i�R���2����h2�H�yx6w�!A�f���9�tOd�Xb��2x���]��ޑ�U�[�wd����n4����ޞĭ�{���o��k�%��}Ȋׯ�x������fPܕ��돹���y�����Իe.��?9��罵������՝�s��n����Ee?�2�����Kx��"��>'ܺ��4���j���N������}܌i�ct�}g�'�,
�R'���}��8�#�Uoֳ
>V��� �'p�N��V�����jOӬ�z;Ζ����Uu9�\i^�~b�ubss�XB9^h5#ҷhtM�o۪ɞ�[̣����e�9�c��ɐ�1?��<u���;�Zy.����t�;�e�ܖIo�(�h����zY��Ij�^���URR�}�H�7F��ڹѩ��Y�Ipյ>��uj�.{.$z���2ۻ4�]���p��TkSh3�<~��<G����/�p�>�<����^<x�F':MS��NCa���
�t,��s2z���=��
��Rw�nt��o/&$�s6L>�>��.�:po9rs���r�_c���mT���0�~	cW���nv�K��!�3�s{S��y�d�
ˡxk���5�xY1��;�g~�}�t|�g*��Mt������%*���wr��{x���˓\��
�˲��d������Z�,�ڐ��H[��I����.��ASRa��LҤ��RH�f�p�d*��ݾ�M�c/���8�r)em�yK3��k�F+9S뷑,nE��x67o7�m�TN�1[����ٺ��Ƃ����qX��;nr�=7~�NE�E�O_��}3�����9l��s�����u:~������pݷ_'g��嵨M̹ƒf�����o>Y$h�pD�ۆ��'
y�{��]�e��`���n��1L���"oUfίeUՔ9o�/ñ������2iT�j�,>�����&Z~8�o�s��j�;���j��;b;�K�ɼ�fx\�#7�_��ץ,�������ןT�']�%}�=A�^���>����1�JHW��ﻸNq����y�p�f���+87D%0��_?�;�����jYy�E�`�
�^��l��'.��^�;�k+,ʽ4֥CiTfj�WJWu�C��op�w\�=Z��>d������Z���Ł�gCX��MbCkycT�7�����r���ssܶYwI��%ҡ�`��}wו�j%�һ�g�a�6W+�*VC�i����6��*985u"�(U��5�X�5���;+f�Aeg-5zjڂ+ӵ��Fu�%nb��o:���еՈ1�u�pd<��F��1&
ǝ��R��AA]�"��8�<�;���58���ku��ZkAA|�CB����J��;�cr�}��n�>��ҕ��̺�U���Fn.���F�L�Z%b	�]�F莾��'70WT1��4��;��*L�3&�nu�� ��I�k	"�pǪ����W,ev+6�GeK�n��S���慓�t�W���2�S0_t��VZ�2��H�6.�ɔ4k�5(�����|T������                      e�zש.fe*͒�=*���!�f��Fo[�mӢ�u�+��]��N��%v��r�$�\T�xpڈY��o�uو��.�y��ܴ�4Q���vU�K%i);�{��஢��3����ܰeA8���]$:������T�'����{U�$YAf�B�*�]��X��,�ofKKwkЫ� Eٕ��'���Iڲ���I
V�V����ۤs0.cP��.A��f|�n��ʸ/���A�D�Y�������,W�L���$�S��VX5����m����\ޕO
���D��S7�w'7*Ч�+��}gx��.�:Y4,�w3�F�tf�(�b�a˖�R����-凔N�p� �{�hodZ1�e>��c�E�6�ά���ٲi�g�yr������t�M� �Y��Mu&M�HvN��A>�RD-9q9^Y�� � ~�+��H(*��E�DH,Q
�:�2��bȠ����QUF��QT�E"���X�DRE'RaaXH�Ez�H�E�Ad�h@D�b�X),��,P4�]E�E�VEE���aJ�"�"�bAbȍ2̒ʐ�*�<���,��DR*�`
Z�e$)'�B,Je1��H��)!v�d �i�ŀ�PQTX-�8�ItaX)U��
 ����ޠS#j ŪQ!�5�c\�{�d����Zs�:��]���[���𝙀�w;7ul��h��]���M͸=[CNC$^�2�x�9���i2����䃞��W���Y�Z%/9�v� ��?~��ɪ������_da (W�,bM~��/������{��H����o:��{kn}�x�n��M~?h��P�+�������N���#���꾮�v��^k�Lb5z����̮p��5>H܉���ef�O��<��VR�����-�N�v��@�I{�Y��[�%7��1��f�-w�/յ��"N~�o��=����(�4�΅ߋ�l�9{��k�<�����v�ɉ���]�>�Y��V�\z�7}ߍ��?0ԥ���}o�~�&R\j�{e�J��X�uE�@kl{>�&�M��Z;�;GJ��q�+��R�c*<j�w��P�(��M{����x����B�<�T��p�+�[x� [�S�
at�P�ܮ&.�A�4����ÓSޔN>��͛k�E���ͺ,�>��y��^][���]�b���ζe�d�ZGֺ�4�f�~Ӹ���~�#���Y�g�O�4�U��FW�j'+*h�נ+٩Vi�l�';kӖ���w��)��i��N~�Z���1o/߼c�_��m;[[(�")�����\���U[u�?��į�Oz��vWc�Ù��O�~�����?4;�k�5�.��<�]��`��~.&��Y���s���9��O��=t���������Y�>��AjD����-쏩�W�9F���DC�L��ˁ��I�M����]cu�����)dm;��ᵹ7E�CH�Dq>�M��b��7:lA���Y�>���{�QW�#�S{��,�pv�.88�2��Bo��������f����Ϣ"����}���4Z۵u����n�^��B����n�/p���T����t�~���gQ���g��v�ztϪ\~�^[��u�#��U�f�l�����\�g�9'��.�ʙ �����<�˪�[�|<m�o���y���}��m�:T������)c�jkZ�֝�g�����<�6��M-	&���$p�^���x�7�ot>F`e�o>n���7ԏwS�\K�7�:5�aII����F��yɧ=Id��8��f㜾|��^�?������q���맱����9�L�a<��y&_2g�'{�	Ԇ
�i) ��!�4����$�K$��0�M��d<ɷ���w^��s�/�[�y�"�c�j����	ͧtr?�^nc�z�6��Y��p�d���mH�l�)��:c����{k*����,b��
ZΊ�B��!4��D�vMޝ���缾�.w��� q&\���u&���3\d�d�N��f��\'DY0�Q!��2�l�Jd�q�����X�w�q�.��C٠�'�6����z2��&/G�i�I�ڄ�y���u�s6����N�L�Xh�$���y�gv���v�I0����:�q/���9���Td�&�i�����v�)�i�'SE�,�K��@��-!d%���늷/���ݻ�w�����4�i�)B�2^�m2N�i�̆Y�$æ��a-��By��6�I/j	�:�����5oz��k>�,�4�.���^H\�q%$�)���L�m�f�L!���y%9d/��d�a���T�'-Zs����7�����`Y��<v�e�r� ��ؼ$���)�L���d�w�CIcr�m�3AԔ���� S�s;�9��Uj����π�I��fC��P�!�k��Ks�.�:�-��d��Mޠh���d�b���������G�����޷�k|��]4�i�$�Ra<b��`y!���
N2o~��!w����w'-"�����$Öv�횾��gZ竲d=ꆐ�IsU	t&K��2j��IImQ���]'Rq��9@d�{��$�9���J޷����z���s\�zE%۰=U�N���,�e��I�B����L!�.z�e�F�
۩t�d�L�d�&�-T^��:�w�6��P��?]��X;:��v(R��s5��y�P���|W�>��w{��C������}����Bb�իJ	@�سJ�1s<޳�d$��/���i����m�N'�v�R����BX�Ḃ.z��d:��8��P�$�/3GY6�k{���/�[X�u���<a�����L�d�{ےi��Q4ْ]	��USl�,���H[Td8ɟPN��(&�q�x^�[ٵ_��m����w~zq6�=�2��,&9F�<��N�u�0�7rM00r�P�B��P�Թ����݃�G��l���������2�I8�N$��q�I��N$�L$öM��8��МHd�2��B��F�&��n��s��F���y�r�Hm�0�q&�:��Rd���:d�i�	�<�$��L�Nwք�AdY����w���=׹�s��ClUd%2S$��d����'Y=��:���I:���M;a7�$�y�,:�4������֯}{�ߩ߉f���C�/TI�$�I����2y�!�Td�'�ƨ�P<���;I:ɋ�!<��w�ֽ��7���w���JL2zv�!cy��Y	su8� �ěI�`�A��P�I's$�Ad<��Gܪ7�׽�k~�a6���e��|^�,�oPq�u��nH^r����nPI�N&-P�d�\�C�0��Jr�z��滆�n��k����L���������@�!�\�Hq�_��u�9�Z�d7]aL�`^�N�i�ף���g߼߯}���=�y��K�V���𽂏�a��i_�h����Y�]��߯��*MǺ�;���w6=�ϴU�k�����s�4^3\VŅ$XZp�X(g*����!�y~�|>�	��s[�}�)$��e%>d.f���y�g-K!�P�!�m �M���N$��f�Y)$���&� wF3����k����W��'Y0�-A2��_0�$���!lWY%%0�.ԇ`�ԓI&�p߻y�!���Wk���o���)�I�ک�r�I&�]�Y	�CE�<�q��P0˲1]`j��II�����q����s����l�=m�=�ORa���/$�K��o%9d�dR]�UA��e�d�I&S�'m��C��K����4{��j��n��9�t�d=���'4��'Y55��K2cY���u/9R)0値��&���K�,�@��L��C��7�k����l��7�r� en�d��i<ɤ�C\�d딘�@�'/�z�@��ؚl�y2�m����	I�Hv����~��}����.���T�C�K�m'P�q�HO2q�	�V�8�Βg��o���``�a0�^�0˰7���s���w�[��g��I-z�H�L:�Y�&�u���l9�8��,'�I�i:ɶ�e��i �5�t���}�Z�k�t���$�Ҩ�I�<� q$�z�עi�Y6�,��:��Sک'X`�d�I|��<�.�8�5�S�_��3�{��&y�� ��S$�臐��Q�@�S%$�i��4�����'���5!�N0��I:�ݻ[����u�g��7� zeem��3����L�U�ǅNk~��y˭V�b$]�%����Vo����G\�_�z�o<�QK�i�2�P�S���痡����J�Ա)�]��uϔ
��cy�;�|If�'�;� u�,8�4���$99S�RCi.U@�`,�I8��t�A�M�H`� m'���u�g��V�o~w~�����z�$�K04�u�	�Y��*`�oy!/��B����&�q2z��I�o8�5mVx�{������Y��R*�y&!L�:�F�O���T�O0�qz �%��u$��m!d'ɳti�i�kܷ;�W;��gXϵ�W�)�ɖ��i�C��d=��`u&]���$5f�!:���&�v��hq�v�� o����s~�)���s�����RS&�=j��&�%�P�d�\�Ci'�(:��!/�:�y y�kMar��ԇY�'�%���7���k����{���fS	~T�&\ RO i&ۥ��R�Y�I�8f�<���q$�R��I��C��1�p���n۽{�;����O��Y-�X�$�Lnټ�d���"ɷ-D�I�)fCl%л䁹������ �~���;V���s�;'RJOb�2Hu�����Y6o��2\�3y+5$�QM�`q%ܦoRB�FS�M��yY1�e�{�{zs�_9���@�2�i$�a��6�[U8�Y��:�Ħd�d�y��Y�ͤ���~Q�r��T:�y1M��Ƌ��{��<^����뜮��	��Y ee!�	&�v�2ƪq'L�d넚��$�n$�qD�d�ɼ�[�m�����oٴ�T[�g��?,Ҵ�[��Ԯ�(����yJE.=q���,�
������\J��8����#ۉ�t�KVv]�>e�A�ݿ8��-z�Z���I�$ �@�[�9�s��	f�RM2���!��S!�LC�P�!�L6�[��$�2�2m���6��N�I��0��L�����o�{��Bm�����d����*���`u$��<�ufjC�0�i�XgTm �w5�3�u�So[��w���d�':ɶa����H_�%!0��Re�
�>�ԓe�`,K�4�l�JL�X_���ذ�߽�c>�7�x�I��d�	��I�l��I��]��u ��R�Q����8���Hm��I�S�5l��{�����CL�p�v�<��/�:�m:�N�M��2N�e'RM3���m��TE��U�`^�I�fuܖOr���<��פ�$���2y���2q��Pɪ q^��a8ɋ��|�c�	��%�D� �3{�Y	}Q�)���q�u�_^�u�W�6��$�2���ľ*d�jCA�N2m�&�XC��hCE�M���L�L��.n�!~�V=�Y�\_X׵�Sn�Y	�5"�Rm�4���b�e�A�'��i�̅�T��e���a-��Bx}T�G�
L������߲�%���< 5�W���}nr�=7;䪡�������ˑ�6��4ϰ����_��^WRqϻx߅�^Ť��r�NV �H3�
�I��j՗%Hu*ۚ���:j�'���!n.͎�/+q=�e�E�^�ү(=G;>���ð�;��a;��[ε� N���$I!{kV�9�w'5?�`���8)�#��[mq�Ѯ��^o6y+�^+�J]:Tڛ�=]����ƀ;���3�qOo�XF{ط7'b����]"�{��b:�~�}���Z���o��������ǻ��%,r�w�]��j1F<�WI�1l�w��9��2zq�<Fo�מ>��į�ṩ4�W*i�95 �ֻ|���5�*�b������'��)�^��_��U<=�7�E�q�ҹ��ۧG^�y���y����w�8z��Q�	K�ܑ
�㺭��m!�h\{�O{�:eOUßm�4Q�x��W��w@C���x�f�V{4g�4r�Y=(�ܭ�x,m�O-w�'��585ՙ��>*f�%k��>ic�N�/�V'5�u3׽��ɇ9���C�d�$`H�XP�Y"�
H)"�P�����U"*(�m�ţ���"z�*&3�u��%s�h�SBS���z����ۋ��Q�]R���߅A�ޟu{:d�eNF�?b�S�K�����C�"c!�G{��,�Gjڥ��Ng�O���7�̪x#���I���^��y�����u4�6�7�z��j�4S^ǿ1��z�������ʭ������?.J��{Q���rt����I9��Z�z�2�C�yՐ!GW��x�x�-��{p�ޜK'=
��[�Yt;�[;�a��|<a%�J�j��>���'m�c(�^�ۢˏ`��k�[NW�Wx�n83�o7si�l[�W��.�A'>��������'���/Y��(wj��z��cbXO8���g5��:hjd�����s:��N+�t%������Z[�Pt�<��@���e��/��nZ�]-��k��FPEw>���$�f�hf��� ����*��]�$�]]�Ư(E#�	;|�WZ��1��,Q�k#�` b�Z6c���z9�9��|''`]R|ۻ��8p'�]�xL�`�*#
�Yw�Q4�|��Ǫvz�Hx��g\���ƏaWMĤ|���1���.�hI^mrX;�{B=���)���|�Y�e�%�O�b���Y՘g;�Z��wL����밂��m@4��^�Co�`/Z�e��	��O���m,Di�]:�������t��"�����`�	8M�e���F��H֫��U5S�ٸ�)�2�o+2Q�0ӥ�AޛLWE��V�P=rd[�;���4���15k黗vt�{����4��vo=�m�����.�27w�vlJ���ʜ"��ZxlTd������z�~�                    �Gvzk����r�rK�d&J�zu�jw;�N��ѽ��
u�Z^%]��hth��M(у ?\�x�fuv<*lwK]����8��\T�l���o&(�	�z��w�w��wͭ����"v��ɬ\�A��q�k�cw"3�Ա��V����U�z�Pc��<���i�P�k������c��t��D�Q����jӡ�ap���V�YS0�D�������n
[�h:[�i�G�zb���hư�Iv�<���+�r��C�xA�R�h��:' ��y$'�n��m��f��iO��q�HA�����y��5���[֫~���m�h6�H楕�X�Xdw���2�Y,-�&$2��I�S�P��'`��J�y��Cz��r��+N�wT W)Y���W�巔pueь��FB]��o�A��6�wӢ����b/1����^�	����  ������$�M2| )4�0�� �,��U�)E�P�`S%�L"�TK$)�	)Y��!H|0���v������L�0�$��K��B�Y"ˠ �fM\�Bi�a,��
B�QL�I���)�j�S$��SiH�a��H�.S��B�Y
H���1H(M���.��Ad�@)�R�G�!f�L�t�)̤(I�T.�Iq�QH<�YH�t�$�d�0��n꯾�Ǿ�=�7�Z�d�6�^;7DJj�=�yk�9Z<��U-t����kslNn�?���}U���afO~�?{������c�7���_���o�==�z�������)�~�³J��썧4�r�܎�_�C�r8�l�9S���A����\��]�Zhf�g��@7螚���V���,~�U���w�q�,������/c��q�������X.�.žƆ�˞�Yި�q{�zB9��d��e���m� ��䟶������y��/T������u�~
E������[�I��u^�D��kg�~ĊHu72T�:�7ns�z�%@Fꍞj���N�ת�Z0X��j5[�Ҵ���p]4�m���S=[ܮ�,��<摹z�����}�2h�!&���Q��EYs�~��G?/�	������Xtm���Qyf��Q�Hnx����{�=��BGH���3P>�����vl�u��E����b����º��n7��3,u�w�aM}���PTpM��p�;_����{AOv��w:}ԛ��z
��K�(�W}2��N��^������6�-M���v�r���[¢%��u�����W�v��g���D��b�IK����o�/AX}7�t4̢��C� �_����$���{�n��!}̫"���z]����`��	��?s�##g4�I����#׻�Ϝڗ�s��6^+y΅�N�|.�Co�sO�i�=o�}p4�W^j��g>�Uw�~�˫�3N�0�{����kˁQ�w篷k,���h62f�O��,`�ѓ�������s!&��+oi=��ޝ����hE���S�������n詐8��ﾯ�����*{��/�d]�{g��kh�e2�z{�]瓻۫jq.�}��0+r��w���{��=��ϵ��[��P�v� 6����UY��S���g�d��
�1f�����G�n"��k�Eud9���Z~ύp�c���T�N��	���yn���[[&H���~���V�h��U��|A�Y�z_��u���Y�/b��مت0{#�4tG=6��JA{�m�V�y���v{7�a�}׾�)�Qw���o��Q�.q�Z񚽝��C�v ��{�㹘a�7}�w�Z��_���tF/>�^�����C��.�i\/�Q����ʍ�zٍ���'O����U�{��=�|:_(��6�<�%/Z�[��p�o���K��������	�&�6�,��磌�8�q��vRY�\��~�ھƎ��ѷ�oD�H�^�i�J�t^e�~+<�t�����1�^�l��9�>=|/F$���X����rI��9��F���]!k���P��9�2a��mR1 k�����{Ǳo��)��Gy/�ף�o���>w�$�s@��=�n�
�'�-����{^T{	S�-��4t�����I2����p�����Vm����<�i�'I��հ�m�V\#"���}��m�w$�؏�G�`{N���76�ȗOR��׷$f�c��)Nb�ӽ��:���Թ�c��t���[k���X4�^���s3�=ZZ
�4�.[e�+i�R���7y���VF^��F�5�{���Q�÷��g�]�պ�&b�:��Hv�ޮ���3>ؔ��}UU�|b���|�g�U��������M�z}�f�5%�{z=�<�N��A"h��M|�~�nec�n�Zх?`��W��oa��n[���k7ӳ�x��I�q�u����ϔ���5=�X����#^��x�)N��z�3���O̣o���^���h&��b���6��̫��ay�V�j7���39yڏ/�y8���d�*�9��-Ei���zb:����\R��La��x��M���{rU��9y��:�,zX�kW	�%�a��c�O��o�mŗ�
�19�u�ѧ�����QyŜ�*ϛ\�vR�\9�<k�e���'Q%��Ƃ�4gqE�� Ӄ���6y`��5��ѡ����^�@rֹ�Ɯ�p��]V$ �m�.�n>���:���Z�9C�cM˃"���U��_V,�)�Y���ZӱH��u���G�"�i&�aͲ!��������L�.�k�I̠���V]d��������T�c�9ی�ۉ
v�&�֯N{�ӣ��f�8#�=x����n����c�-l�wE�QS��j�2�nP;ۉ�﮻U��yvn6���Ej���
	�dࣺc��`�6O?���Oi��׏�ׄv��1m�����闹��9�����g���Ԧ�HlG���V�"�����t�a8F�{n���{B�l������3.if�D��W׬��<��x�s�k�4goQv��Z��8,%��07�^͚�EQ�������ذ�볜.�����q��qު$a�2V���,j4���}G����܄��Ѹg�sL~���ie��̲tE=���������|j�rw���jF����JN�B��Xd�.�$�%�s�K�o=� �6��G�`5���᪸��������x�/*�9�e��oބ�RpY-F}�o?7��E�>[����y��K�.�$�o���|E����]\b�{<%�1�Kvo>E	Ɨ,Ϻ��F�"T�uy��\>���#���Uv�lG�ـ����c^�T��ێ��_�U��(��U���c�^P�����[\Tc4+��ے.�5mԪ�+I��u�аnNl��n3;��i��wC�~2v!J�
��>��(�v��2RX����L���q�4�U �5±��j1鶚�����.cQ�X��H�t�GC��^t�S�[����귑�=�SAw�T��=t}��?�ο�J��>��ft���5��'���1}��.>^ʶ���i{g�ez�ǵ}��v�Ǘ�S����f�?t�S��6��C�jN�f}=�#x��מ��nфz��Aí��Ǵ�޻�o'�wO-�hx5gF<����?t}Լ�{¼�ߓ�>ԣj2�g��3��86ψ�ۄb��|���9�eo?={��Z��������WU�n}24/�q��;j�Sm�ն�[�}s���=�;ʦ�f-c����xS�������o)a\O-J*�[>t��*v�;��������T�nֻ*�"��z�u���s��=��/�GMȍZ�5�u���+#Pn�h.�oPOY�/gY`�L�;�W��q#�c�}U��X�"��L����g�c��8iˡNt/��	���O�ǫ�j-�_�dVԲ���*2��ɦ��$���8<^�'�«�eXT�ax�ԥ��:��j��8<◴������[.�ί�<}���]0q�w��+�4����Q��MQ���K�'�vnr���&���^JR��b���X�?S+ѦckE�����K��b��Q�ѹ"���/���ѻ�n�7����]<�q	��nm2�B�s}���>q-M���i�K��̯�S�
s�ȿlm׻;���
)��J�/�zX�p����W^b�
vW����u�!��.�U4�tMۜ9S���)G^�[�Iﬅg�RG��f��wn��W�|��u��}I���!��K�� �]�C�.0�Z���D��������=���o��Pv%;>]a
�_�4�Q�姄u�0�t�_�<���]X8̷^��p����`�[̢w8l��K�7/M�zo��A�z��1-C��P���T9@����ZC*����?�+�����A����+e��g�k��5�Ia��\�����.��76gEH� ���m���Hʷmi����(}I��B'o�����tE�2�$��%��	�O���?4,D;4�y?,�����Oq9Cs̑yԩ�1Ъ㖡�D,�1+�!����ofNGH�x�.=��0s�4+�*kqJ�P�������O,I�U�^u���	A��٨1��:}��7�vп[g؜m�׭>ݼ�~LO�z*�т^��CDq:��C;��G�uS˵���Xg��������Or�]>s6���s��E-�:v��48��բ譌�,ZiN��t��eh��$[�-�U����oI��+!�(�u��:݊Ƴݷ|����t�AT(�ۢ.�}���j���Aee���um䩗����3р��
���p��JZ2ԙn��8aٔ8aR�x��Ztnsuc6�&O�.9u@6��4�����V��h\�;LD���N�İ�>}9r��y0�S�R����B�I�C��qݮ%M�d�ze�\\{�l:��Tꌱu|[9GR�v8��t�]����yh��q�����I\v�w�J��,h��0ӛ��a�%_��s�C�5�
�Gta���Z��B""�QW}���=�����L�8B�f��`�E�N't�K�+�%n��0z'��]�\>C�ƚ*!W��ou�\���N�Va�Ad%oj7���?;�K�\ZUΘ���� �;�/6E\ �%+u��o�m�`���L�	�v{dRH                     Foyle�2���rIxoK�)�q#�9���]з�f�ԥG5oB�Չ���V3�>4�Y�M΅=�I��㼬�O^��v�m
*-{�9 ���u�\/s�+G�h��wH�Yf��]oO���Ƀ�;c����`!A/IAk����n��"��71�.پ�t�zYDZCL�V�.���Y߳B�cĨTή������ڵb���ҰK�J�Z����7:���W,�>ɄW;��q� Y�RF]�d�vq�]�-h�۠��箸�V��㽕�q����ł�U�1��㣳Gn�'�š�ifIB-Ś�P���)h����E̧,k����0���� �	M�4Q��_!� a���i�秎���ܝi���8_e�đNl�b�k`��3
Am�'��æAj��m�;��J[s�S⨅Nǽ�@�RsT�]��/�s*�g� � B��c6v&	��c�I)��2��]��S�	L��lԀ��!t0�'�;K2Y�-j�XJBS�Z��֢���Y�HS�(Y�%�2�))��J`�.�L)�JJB�2٠)${�r���-0��I)�SL�a,݁Hޅ)�!*�
!k�K�2a�˺J`������kT�P�Y&����[6K1T2��i�I��,��S
@, �*U�ien���n%4ɶ�uJݕ!UAHU�a"�ōP,�0��h�Z�˒QF���K*�KCwO��p�L�xj�s�V�v�N�%a��p��� >�׹��'�o��ܡ5y�5î���߯ `}-W8�-�\FM#�'q��P�"�퍺�|�c���#��P��Z�Y�c�z�����6�O�v!B��:@�R���l�᳅*����w�M��1.i��,���$:��c��T+�+�yGaܮ>� 2f-<�{���16����L{o��s�/�Wm�C���Vդ0�'1�u���&2��j��eq��������i.���cE�\p�=�-���:�0�
c9�}�iQ�U-���W���/z���s������ܼO�Æ�����!�=������5���9��4�Uz�ٝ�`�6�J�K�r��L�S
�������o������\���kX��#۠�x*�Z�֢����_�}��vV	���X����ż��dj�J�����������nQ:&�n���sy�JiSګ�ulCY����X�q9�e's�hf��f���9!0�Ǩ���ﾬ���W��u��(�g�UǏ�Zy�)8�k��[B�;���̑$�KVC��]�Ј�eD�@*V  �#��uK���΋��-Ů��&.0ŷƇ#�b(��M�ʔ϶vg����#���<<��t���_8n�
	�����Uq���]h�e����RP�^�evN�W��a�t�yѡ��ش���������$	JOǪĹ|���UC��J�[�W��^�S7�#S,v����\�~:f����#�6@:�hU�Ƭ�3��2�� }�e�}��ψY��O�$��¦�z��a�HA}�0)
o�\�����Ck~�P�v@1��5<�y��.�q�d�����P�]�1q���Q� ��{om��7��z�G*�^k�{�rX�#�L�e=�
�|�b��4o���{�U�P��}���`.xN�;�\f���v�-��[��u&D��Bw�dF_㇑�ORm��6����A��Y�v��.`��q���磌밦t��� u���5|tF�i� >��N����K�S4ֵ�7��V�I����D9��(I&�3������|��P��o�Xh:���e��|p�o����8f}5���
[�r�t:���J�M�m����B�����~��v���Ͼ�h��4�8�%�[u��,�=���KO���Gb�Z�FOI0B.�[��6���Ky�1s����B��v-C2;f8p�/X諪P)���fvNF��v��As�7�):���V�N�	
�O4�u�^z�zW�N��gJ�x|�B�,������)W�
�h���eP�Jeפ��9��(x�=�W���hKZ����*��HiqU$�m�^ݝ�A��cz�� ��
�"�
L�@Zv�	��|���{��r�GG�]�u�Ӭu,zs	0o���zXE�L�:V�9�o�;��{�{�:C:��%>�#8���Sp�Իڹ\jUŜ�L�Q��N|m�����_}_Q�����Eq�3�<ǹP0�3Y:����Fs�G��l ��o332EB�MPն<�WPJ�i/���Ý�������ng�3b�I:CLQ�T-�j����ґq�����<����:r���h����V_`�
a^Q�HWg�τYH'~J&�uy���j���A�t�z�e�]����"y��Z���rT�op�^��i�u8��R:S�[�na�l�(C���b˫�뫧�i'*��w�K�t�ͥp���l��ϊ�"�W4�;ڬ�����Z,�L�<���oOR��1t�u��T�4�';]��l*��ӄ��f!��t��*kL�����(�|��r��2A�t�3QJ�cþ�@��xl��j�u��S��b�o�B����fS_W8�Mt�`�7R�|䫫�@4�����a�Q!�lE8GNEu��.�}��.�Z��JB�������m�f��,-n=���O�}�Ufd��{�[��lQӪ�� )l]�x<P��n5��6������)�|���N@�
d`>9��4�h�`�.kqJlxcX�W�q�x�����3uv����t�D�P����F�9N��eb��5����H�m]
5js����T4j]�w/iI�����h���SÉp�o��_;��wHW��s��D��`:��yׂ_�Y�ړO��v\�-���&c�i~L����/�T��Pga�8��%�z���k���pz��>G��cե�L�n��g���̗����S�i�w��پg��P�+�y	Ȩ&*/_�Z�_��-������^P��Ƙ��	8��5�>_wMqĩ!��L�&g�3sIC��J��E��C��+��n?����W�����-Q���������f�9�9�Wb��_@�<oX��]kmx��!�+����#���)zD�CRV\���9��7�����Gf�AŊ�X淲ն4��̖#���gd>�O���8�4#]�h"���Y�6,տ_0���P�~������:��j�پ ��GRD��|~�롭K�]��5����#��P�e�z��W�'��zJ-Of�,�ye��\�6W�>��wJ�{t&�Z�a���~�Ua�k)�z�v3�_O��ƨa���t�7ǎ���kJ�՜m��'����};����)z����<Q�4�T��+���;��=4H�����ި��K�jg&x٠W�m�ٛۓ��3�[$QgNJ�j������wf]�j��g(�(9��7`F���}�J�f�t��~�P��v�e����p6ã3ό%Of;�})�+8.M�~�hV��T?���=�ٱj�g�	4��Zhmu"t�Gjfةy��l'�m��Zt�Iw�]��v���x�9��H�A��2y9)�� ���;r�CO�YiN�!��K�rn�j�%���������+�x]�;Lu�>������I�2������ɛ�?{��ln$Yߌ�{T�K���\��g����8�
���l��3ILA�a����^63K6��Y����ٲ}k#��r���;=4h%�V�5�Z{������o��EN����裔�xL�zo���JF�� ����'���}^hR����]�wh�66�_<#"�C@$M���yI+���s�{�yd�)�U���[=����FDǗܪ��MAg<hq�2�Z�&l�*�� �����\���p�	�lPl|ޓ�ճ2M'�J�ӱOf".����c��YK}L2�>5��#�E�nd��6�>\E������[�Z{#���c�m��uޱ��q�4�O(���ד�6�Ѵj��j�]�$�e.fn������º�r��n��T��$\H�~��d�ws\ZԎ�cBN�ւZ�;Ѷ[=ֵ����3:j������8���{�:LVC���!g_��,���	�w����{f����~��f�\��7t��]��2xQ��ˏ��
�9���Ξ�-3�p\t���+�Ӳ��/��H�o��CK��{4�[��l��1B�����l R�Շ��1ր���\��<����Ϡ��g
=�cܨC5�����<s�}I�65x�UW�����妭������\lU�c��`,��O��,y����۩wʙ�^˫w�'��t�5�����!8q����7%��������۸h���c�k����nz�f��1�[g��e�l��J��6�2xUq�ٵ�����xU�%�L�r��{#'8D'
�g���U��،�=����xA����)���y�O��G5>��xΕٯ��(�e�O ���6��zFcI3���A��C�r���b�� ����^^Q>��)8�~��_��˷ǎ�8hr��	���[=B�4wۖ����fflK� (a[B`���p��Hz򴭗�h�eL�V�4�yOt��!u���
W�"�2Eן|֙_nO
kb��Kӝ����bK���D ��Dd��f��
͚�~坂����X�Y��1�4���
��C��ۢFiZ� ՞m����C�W(vo��8�9�:d���8�d@t���܇�H��r�;jSb}r�\�X�ܙ�:�Q��I�C�:kB��"t�ch��g<�̸���X�󂕝���<+��z M�0��*��D��4�}^ʾރ�"�Kd�
Ӿ�t��ܡ��УD\�/Q>W-I���G��'�e����Gh +ɨīzj�>�՞;�n�D*���z�@U������~���h�6g3��
��M�^�C��K��e�����#�-���wcfHFq���HfA{m[U���T�"��Q	'<�+�����,��	�k���M�6�\�j?Cvmb����5
�mC�#��M�L�-£x��z�nk"�˹£��e����4��ō��P߄ʻ�t�L4Ǔк��6/?i��,y��Zt��<f.;�L~]3��5\q_$�xB���9=�u��!���X�t8��+���p�_V`��5Ҹײ��4�nz�s��G����F�G����;��S��S�e���jVuY��{���b��{I$��K\H�����t}/���O͝�3/��j�z��sT��������_%����Z{>�x�\���ÃX�7'^��Vz)k��hsV����FM�����\[�O�;fnNK������7�
�aѸ9j\8W;��n_�����޽͊�j��F�_/��"�ZaG�=��:��C�vw2�x�)0a�ދXiU��W2�me�,+���熰$M�[x�n4Z���#q�鋗��G�*ܭ#[�X�%,�].�y�Kun�⯦���&�r�a�+Usn�`Ǽ��<Zp�[\n'c|�ĝܗ���jH�]���ظr0-�aǚx�f�)�v=�¦Q�[��F[ɷ>�����v&��Χ�������<7���'K\�/c�y�{L��M�Jqw�B\>�T�dy�m��u"%�%�]��q�6���(����\3��\�o�I�D	cyY}�ݟ�8U����6K��]��6q=C���(�]�6����r�<b�Z���r�܎N{R��	��kI5�LW:�˪��5�l��0�:��ў�w��o[�\�.6��iqY�$�\�٭r�� jyc{2�����`���u�f�r����XU�(����G����>��-��M<����J��3/��=kU��c�v�m�7��$�a��EJ�!H�B�o�Ԩ&���/ٗ�*=jE�V�����            @  �       \n��^�� S:��j�*%S�iX䯧dʏT��ٮ�P�����՜5���S�ʛxD���]_d���t(�}��^���)Wo1(��R���)��6u�+�v��u��JŖoq���Y�Pg_i���͵6�8$N��N�iN]��9�V����Lx�Ma&*(!�P;��G���0�P�\��n���l���9k��mC� XW~R���*w	K?h��ՋGV:L�T�̵V��n+�]/WR q}w��B�ڝ�e: Yz�dZF�loUgJN��\�b�&��O,&0]c�\�w�������"�+����F.�Z��^Q�v8ͧ��p�9
/&9���T��w�
�s�|���u2kX:U�7F<��J.�D�:���sy{]ě]9�u�W�|�h'nU�c<lU�Ƹ<�e;OidK%j]E�}1�P�  !�
~�&>���H�b�,(e ���I
Tj�`UU	)$���id�KZ�Z��e�d)p�j���R�-SB�IH��IET�))+5 �(����V

C,+����D�������J�!LX9���i(��E) R��"4�*���,��"��Y�@�B���V5R�"S(@��VT��JhB���S)
K�,X,��"ABɛQ��IdEX,Qd�A�ZiD0�BȱM$�K�Je1@DH(�ILUt�%2] ����|�{�Y�L]�a����[�m�����*�HT�e����HC�\��e�ɟ�T^O_�d�!�Y����;��\����Z\x�������-�Uwd�4l��Dd�(�1|L��L/]c��̺��ѩ������c̓"<�f����w�`A�����f� �d:v�P��ր�׫�
�SN9�ע̺ʄ���\�qq`�5�k�vzIs�v5g�P������ Cv��gη6�s�f����<y���Ցo�޵�C����vؗZ���=5_"���}�d�������z���q�k�~�W���}k�M|g���K�p�̬��rw���1h����
_�;�[.aeG/�y�C׵�v��sa�Y5����4��F��N,2�t���\)��JU�Z1�#3�<nC����+:=#utP�M��/�F!��:TXk�S���nW{�k��(u**o��L��Ը+5j�}
\o�V�g����չl�κ7�2M�&���+�W��9�!o%�ʅm�>���\��GR�,�^��V���O�I�&H�����,0���N�o�Ӿ���´ ��Og���T� ۅ9��bh��U,���o+��C"���n���9��`���6gr�!0T,g��	q�y>#��YKZ�\R�~sS��VlΈ�*�&k�!��]CB��~:z����c�
0�PQ9��~���C�e~l����Cخ�.9hY��8���N�-'���r�"Gx�%P�j�i)Xz��7�1��Q?9��A#�����*iTK�s��/Q<�J�𝔭	|Z������\F+�rp�'��y���ET��
�
/���0�5aɃ:�K����eK���G�w�:� �T:Q��D!��WD�W�O��驕����n�k*m�>�_$.*�Ŋ��B+#|���T��HK�'���̗���l.����񒶎���m�����-�7Pf�}3�Re����V0s2C�{3�đ���}�F��NL�&F�qAGA�ϦU�CW>6����A��'Hx����hZ[�0��V[���ò��_���}�Q��6�S��Oh�};j���[G1a���ZKk�݂��Hi9�L8:�)�q΍W�0�＞�C��!�do�u�CYMҝ���W���Ö��C�Oo=4/��w����0����%ڝ��s�I
\�������I�;rLoW��۞��p] j�U�͙�$��!CRց�8��W��9.h�d�:6�py�1��r@�M�L���b㦂H�C��L��̣pyM���~~.�no��w(��&��s�$�,:��`�t��<�����y43�g�u*>���u�c���$f��#�U�*�<r��S��wwftHPe�t��(��شv�U�WaRڼv����uS�Kp�q�yk҅J�_���3�;&#�:gN�-�,'��F�f�Ya|L~R{�#�P��9�;q�{򵙧yԉ��2��E:�E�����GaX����7ӳ���U�ښ���Zj��p�@��D�P��Do�_���w��c���пc�.3��/�/E^���N�CDq+Y<zv'�=y6^d��#5x���NeX���0ͦ�`����X���ѫ�L����U,J!^��3�P�����0,�01�;c���uOŲۏ��4j�F����Q�pz���<��W=9�J�ۣ��jm�3�ԍz��ǽo��t�2^��x�svk�Z��d�DN�P����_��J�Tzu���%�~	���	�a�G��N���j�#9}��^,VÞo�J)��gc򘲗�28�s�wF���Q�6�iVD;��J���|��\o���=��;����8�+M�J��6u!�xN{-��_/�`�r:��YX��gY���m�B��w7n�P*�<�v8g#c+�Cj�`�ÙҒ�i�B���G�u�l�N�H(_%�9�jŁ��Ɠ�U�;��eOۇ�+�W�6͘��	aa�������~�f�߷lK�~s���{=r�_���]=��*`�B쬦�-,k .%� ��Ⱦ�*0�Q���;��Bu�p�S���2O>��6�p4T ���"]�xe��<�v+�(���'{2�Q�'��}�M��|������w���/��'cas1G�R�h���Hܰ(�с��<��t����z�OP6������^L㡙X�y�����_l @:�.���V������<阼[���a���{q�uTPܛA�]+B���T?���luu��nlb��	�N�(�5���hj�ʹ��E���/���@x��n����:��5�U�`U!�M�<zs�8�j\�^�ͺ�k3mf26m�\��˂�H��p�@,�}�*�v�n�p��YLsi8����Z(����x^.�e������}:�yzn����X�w;(sL���z�ӯ�y���������A�hE�x>,a[��d#�K�&ޓE!�Ş)���~�����/I�3�Z�-!5�m9�[P��aX�S��������'ܠ�a���4��F�2qa�1��K�������j'���|������;�P�E	$�&yX\��l��nzǷ�gt��Y|);�=�:8)페���Yֻ�ڹt���{|W��I�9.�V���/ ��1C�}��Řfx�K����$��&��{'��ݏ�7�4�:��Z�>����qcRւ-ܱ�3����ٰ{��Yv�K��i��8Xg���=��C1�Y�鵺F'��ם+��!�S��t�'bG���x�S�زb.q�ޯV{��6����F�K�T7O�H^�T�3��iZw�UY�_pnm߾����ݽ�M�T��Z��6���}���R�e���s�P�I�h]�)$S��@�6]VU�X�i8�ξ�V��'Ʀs�+2�baۉKF���V�y�ꛗ���Y��T������{$t ���Y����R��Nq�A�t��ZV�/��O�x��Z�U�j�� ش�9�=p$}w�좾9��!QFf�u�;z���#�[5�JAz�\�-��_���Aޜ���7O{)߀��h*=@F4�ߥfY"r�3W���+�ak]�V�v����8�ϧ"�~��Q9���:��g��5T��|#��#���\z�f����pQ�a��L�4�}�����X�/ƾ!�dw��w���Nf�nt^dOFK���zz�x�->�=��s�CAab^����ݙ����F��U�Qq�o��p�!x���V�ˠ���l�=:$ห�f{bZڱJ�-h0��/%��������_tƉ��.:��l�zE�) ���k�B h�[�Q��Ԯ|�.;��vA�oNYv�a�w(�5��J�8��#��!���+�7�h�@d̩�4��W:���î'���5��OyQ�G�u�ϳZ/�Zt�H}�u2y�2��;�p�i!ْ>�����㗑Tk�qeNboJg9J�xw���	���g�g�Ȓ[�]�3�)W�NX�
i���$^iz�5f6���i��7۫���E� ��!݄��x�,w&eK�E�*�@�o�U��z|[��[^J�5Mb����Ʈ�ܸ|
�U��N�Q�Aإ�f�d����Giƅ��0�zxx�V=%���P��g��{�>{;� C��XЅ!���C��ȷr��]������	t��}�z�"�Z��};)��h��:�5�1aAe��c}�x{�}6u�
cc҅tr�>圦�B��t�`�e�"W����^����zi�Yz9BCXkE�;W]v.�eh�i�ZwI1�m��i �e���f�&���k�[��{m>��7+���.+89�:oz�o�e�_���m�&rfc��,Ƒ/fq��,e�rEW[�4#�L�ڪ��W��3��j�����-/�w��L)Ƙ��	����1(]{/o9#�`���!�060�<If�b��m���[�k�����t�f�#�D]���Z8a�as�<)�b�iTD;�Ė���{_�/ �~���+�u^p�)�����w�.$K��^�fqi�yC��d݇�ݪ)�kv-c����Xh���Xz-=#�c�9T�W��x�"�Z��P�W��Jյx�����D"tj�_i�j$�++`+�XoW�q>8a��[Zz�Uq�;�q]�	�-/{7wa�VR6m�2װ�>0`������.h�q})l�����1l��`�D
�Lz��"$Ve5����}h��-.=�:�������JY.���,��#�`Qw����L(��ZHc �g	FP����o��H�׭x�G���C�ެ��`��pl���U�/,]�*S�$�p�[��ʰ�
��$ȏNn=كs��ɰڠ{v�877xo����'����b�����@�����7�wj�a|~M����ݙ<g*b�;���T�1V���?�9�q�.M�~t�
�_^[��l�w�7�����Va}�G���[i���)��kh����"���xb������>�H�A+H���#�u[ƒY�R���°�wa�w���Q������T��J�i������+v�̄R���<���9(vہ_����Y�M5E�|d\^(g���j~�%=׹���l�.�,0�T�9kj� m�h+�(��wtC[C�����`�����x�b�K��E	$���KT���뻶��s;a�8c������L�ધ�:������+O?`�����I�.�As*RWR��L���x�����|��0|?Z��������<m��F�gU�[-ԛYǉ$Eus6�hQ�a&��6��Q�̭G:�:Mr�fk���im��v!���6ֹ+��@2jV�<�hY�Y`��ZT���`���"ﶛ��uۮͣi���S.���&U�fS����+�i�8#�J�=���-�ts�6�h�Y9��l�vXHkB���`�lV���H߅� =z� �[�*��:BY���G�-��nQ�W|�]�f&Vs>��۶�r7p�9�k��eM�A���{t�i�v8�u�p�W.���C��6ɝ�m>b��h�Э���]dpjw��N��i�m�@�@Q*��q��n�p��ܜ�3Kpl���c�;l��E��qډ-Nm��w,�*� ZD�d٤NV����7Z�ǃ����8���3Gw,��K��A]�2fY[����Po,պ���J,=9�Fq���^Y�5w`^��-�x�ڏ�ɜܽ��#w��wsv�K�X3B@�+�Nַ�:�8��V���!���3_�$                      �r&o>�`j2�I}y`��_��h�^��Y^ꝲ�EZsJƶ���'8�wu`�Ի��@�:��J�]�ͳ�Cй�^�QJ�Kde9/���W�Qs��-�����h�����D�ݹ#J�+w�d�hF�w\��lt������S�Zͭ���V�)Z�h[�V���]�KZl|F�`mY��yM:s��S)uٗ6�7�; ��dU�H�Z�>�.�5Q��y���겯��t\%��'u�C]��Ƙ݂`�[�bԩ��Be��t�t�H@�y���sЖ�]�ΑJK�3P	�N$����m�Vvb���ɼ\�u5Q�sk���v��d;�f�r�ͱv����_[�j�ɕ����WZ��SW\��έh���*�Q�6�#{�eؽk)�mf��f���	�i�GX��\Օ>7ogJ��gg^�9�j#�O$ $  !�"�>����fb�0Ab�H"�U�"���B��R(���C"�X*��P��ň��
@DAK�3(��Cm"$X"��*���7LX�Tb�b�!��E�lʽ*1PEDb"���`�uT�Q��,UR҈�QKU
�UV"A �(��Y.��QH�U0�Rv�V]�UI*�b�VE�UU��V$2��1j��"�"�IH�DU�J�U���"#�F*�A����.篻�g��U�';e���/g[�s�L�*h)�
1�Z�#U�0]M�Ə�����?/x^���W,�% �+C�S0��n*��`d)�u]_x�.K���+W.�$L��i��8X�Jպ���4Fq��_�h��j\*�⡺-�}3�N��AG�:��8E�j/1]�qn�U��wyST8#�����ޫ���<��3�%�y�˾��u&t��T`"��yçA�z��W��e+P��,�x:~���C�ğ���t�,r�Tx���(�s�OI�H{�X�}���P�}t�Sa�0 h������,�L�����^���%^�)x���C�,/��B+:�A�uB#s�1���1�D�8��K���iA��ƾ2+6E�0y�'U�קּk�؏+ζV��]3;�aVr}��WGּ�R׹Cu����g�U*X.fBfV�~�y�kЭlY3�aXN��+��^J�Z�oϦ�'4n��p�Yk�ѧ%<� ���{^k�2k$t�,J=��G$�_ߚ�p~�����N�r��v+��<��g�ӯ_d,Tħ��������^������������i�pzW�l��S�ioU�Ρ��VB�M��W1xؘ��dC�ص�ҽ\e���}<E���#�=^�1����
6e�P����a�=KZG�^KqKXa�W���])z�7e/�sJ��m�g4p�� �ŵpLs��UGf۳G���$Ol�\�
H�elbW����"I�Xu.3G�'���S��U�Y;:*g�4E��:�<�)�!���d���TVc�6G����'.Eҳ��O�sD6
#A��==͎<�-tA��~��C��{W���ۇ��%�J�GN�����즩�|��� ��v)������<.��r������� jq�9���I�Ύ�k֊�� 3�]g�X�=�75}ފ�����֣������8�ͷ���M�;�ҙ����S,J�̽ն����K@:X����ƌ��I����'�~�:���ٚ�)lSuC�Xs�ug<�Kf����A=�oN�줬T�� �Y�e�S8.h��x�y�,�V��N�S�'6��p^�{��:�5S�j���B��}��x�)Iz��ǝv˝��⎘2�8{5��0����Ƀ��Ǫ����b�>���[/�J(�hqyZ}kIyᘴ���<h{O���7Z�Y1*v�`g�g��\�����Y�X��-�﷜65�&�d��.���	\Cz��H���u���P�=�^�w%�>�����o��zۭ*#���#1NET�e�f�����J���9�#�瓚Sʷj�?b�ᾧ��m�]S5�$�@W������x.v
Νѹ�/�V(ůNz�J�|�1�N�a��6��{ϯ����/ɕ�V�{�}��������wC���;����Hb&�Jޫ�	�%��h����yt~iY����	�m�������p?̳&N^]c�:9_�>���5>mu{�1�S�����"��|^(aQ�knm-�r�>�S���	jAx+tc���P�W���/��Z�.�oMD�][�f/oUud�����*d���Zo�;E�=K�A��*�2���(��ؑ.l9Tg#��/�<k_���2E��)=��(��Q��\n�X�1U��^� 4	n�{��;�},�����h�yy����������lt�c�F��I���!�ג��V�{r����r��%��=J�rxf�X�aO�d��g՜�ݟ�zr�k_/R�1l޲E�p���-��׍�7�Nn���N�t(_������)�"��YB�>KG �>q'��x�R��ͱ�;%	۞���W�	��?ynW��k)����ײ^���w%��R�^�0�/s�`�4�o���^�DG�o�*����Y��E��N�z�%�W��Z]4�8�1����+6]l9����;�=Eڟ�f>���ݥ�4��N��_��
|�<�m_�HT��r�Ă��V� m�v��w)Oo���.��ѯd<�2��>8{$���V�qϵ=6&�2�c7��칽���f�8��G��=�xx�ٛ��FE���n{�.�K�%v�gD���A��_yys�1C���>��默��c��_p͞�k�E��6�B�ack���=|�K��K�uɆ'��)�X�p֮#y"|5�h�CB��~:z���7���ܒM�40����$Y�(t�&�4t�������cv�ʯ*>�/m{76&ձ#i�Zl$+�4�[�3)��;�R�Z<W��G|2"����=͸��B���x,1W�[�Ww�J�������I�\��^Q�	�DT^��2఩��8@�_V�5�X�/Q��GH�i2�������m���#�(ͽKq�Ȇ�s3�u�@�nEѷ��
sR�c��� Hie����Y	]�YkN<Y�6��z�k�U|'���΀�=�?������s˃�G;�����d�i�_\[;�f�TnGf�xQ�H��^x�����!����/r�s�����
��Rc=k|��Y�-)HY���U�����^L̗cM��vOki�OKu��E�=�ͯ�S�E9���@��UJ��z���ߟ�������\a�+S9]1�5p�����y0��O>Tt|C��sU��5%�iaș����\ٟ;L+,NY�R�/��yp��Näx�|���qI��iC�{�$�<ToUט]�R�n	���
$�ޡ_th�|T9E=KZ,���▯��3�z�/'��M�������컻I�nݑA�ey�M��*:�h�thn�G����P�&^�&��x��tFOhU���ܧ�f����%�D�Ђ���3�n�:�=��M���g���c����͢g�o4D������eax��fֽ�L�Ke��!�y~|��N ����"�y�B��1�1�!Mi��f�(f��\+7?�\ɷ���m�7-����TB�	��Q$�J@�����z�y��_6�#���H�)Y�P�Ǫ독��PJ�q���\_���G϶l�'Ǌ4e�b���p�c��W��r��~~4�j��v�<�o	�xT�H�+�+�s˵�%�8tP���`�*Zܵ�I���!s%��-K�5�t��z�	��?��䷞j�s��j��<#�veF<�>�trע�T)�P�;j_W"��_zflH���.�6j[�V��y��R��9�*
�zu�oD�'���՘���G�$i;��ִ�,=�OJE�O�Y)�R�ͬ�5f�q}=����*�;�H�<'?��A�ŋ�C��+�z���;��ʺ��X����cqF)|+9�O���E�׬��./���%8Evŏ�M� �,�z�e����8[�x5��2�n�O�����+(ǌ���x��D\b�B�����}1!jg@��KW�d�v�=�?]z�	��w����YM�z<����/��3�]�� �	�H�-.�i��g���{\�v~��~����\a��3CK	8`7{����fl@����ל#Ƃ�Nz�J�|�Jյ�n��D{pC�IǙ{���>=k��OR�^�d{
�x��aG�i�#�~���F-�֕MY���^������b�Ĭ�h����F�Bz%\��&�:E�����~���[�}h�����M��;Ǆ�ᨎ�B1xKD�� RA�.��oE��=R�w���uV��$� P���X�u1�̌�[U�b��2Wב���6�|:�<|h��C��qB��|DjqW�.M���8W;7�]ɚ��"�Pm�Pf�6�}�&�"���p�҆1mT��Ur�m�U>3��#Ɩ�T��*��������r]rL�C_!Io#�o w �ګ��e-��UP]�//xR��ύW^�������,r�l �@���'����ݙ��ߤ�T'�f��B�>"�4�]B���6h�-(�e{�_^2��=����e����q�[�3�҄`xƘx�_^�G��ٻ��xK�ַT2.?T{���D���$���b��Z0�e���.wo�|T���Z����]�b�4�i3�L�Xxz��4����R����.{j׽��Dm��.=�5��I�~лֽS76*�(���0�XlNp�Z�Ԭ��7��dO�.7c!��==.n��}#K�/�sƆ(��n8~���)C���2G��w�F������Jg5#`�9�����->˕w���g�L��5�&��r�fZ�[�a����#9"{_��q�4(ڷ�w�y_��˶�!�J��m�R�,lc��w�WAή��/*C���`ݼ��Z�NvI��9%�Ŕ�]�EK��ƾ�M��n9h�ᮺ��{��|�<�nEx��?Uy3w:/#����>413(k}�(WK�k�4��7��ФO�}�3gV�\Ĵbv��-�����꡾��C�Z�������;sb�q�^!�KO�^�TX>\t�h\X��6J��'i����Ξ�r��{��h��xQHi��G�*ޔ}�x	OI�b�u���GԷ�OӽH
�՝X�a����,:�r���L�}�=�_Q�l_W�۹�z�����Ȱ������Y��!qV-5m�Edl>���Ɲd�ؘ�>��m+�ǭo��Ef��iJ�N�*���o���͓'-L���V��o:ya�Z�����?|�R�}Vzl�d��x١�|
���;�Y��K9^��];�����Z�������q�٭0�O��ސ�����zz!g����>�U}I٤#���*]��8Q��<�2'N�,���k���кӄ����v�'!��-4��c:fJ3UӠ��2��dd{�E��M�
��L�y�E��Uk�$e��B���"a�4��}���WW�em�w� �X�Ft �tܡ���P�N���vk"L�_N���YX���㛗'�Lz���X�%�K5
ù�O���@�B1��_n#���b�s�m}�����W���2�"V.+R��Q�7�M�5�^�F���%��9���+N�|��GQc6�Ҝ�!v�S�����w�1��B�IqA,�+:�\��:hf���i=huY��Ky�ӡ{l�:n�:��E(W58���2��y�?0C�{�z�m�4��v��ڱmV&�Zn��f[���q4i[�M�����FD�SJ�������+X"�({��S��R=�N)a��K�kGOe�V�j���bt8��t��i8ܴ��
���J"�˽呶�uF]��X��ƀ                     #5g���2׃}�N��w?1���2NkGP!wGCGI��r��Oƻ��X�֑��p%w�
�j����[De-_+�d\7\�Ly�����{W/�b
��o]�Z���8��&�?�g��خ���/�s��[5uy�����t�1�)%K0����<CT,ìY�ǦF�V:�Y2�-*�|N�zn���*��^��	kw-�"f���[���i2S�*�"��u-qi��چ���CP�c�`��ļن��sP��;E���<u�ncu��}�_�J��tΡF���K�~8�Y�R��mCR�����_+I�8cK/#ʕ���3��6��b�hT�6d�wkr2�n?��ui�S%�e8AT�|2αY�/h	��Ҍ�Zm�ӕ��ܚ3��,��EfTԥ'xAG����/oC���o,M5����!��0*����$�I9���9�s�����0��
�(�Qb���H��"�DT"i��J ��Ш��
�H�a(E�٥dX�(U-,X�b����QEEԦa7bV*�bɖB�QE(�IJ�X�����j�ETc��r�QTUX�ȰE"�(��j��1Eb�`�e5r�1b��Az�Y�m�"3-"*�TE�+P�
 ��6v4>=]g�rFD���Z�Hu�GEt��֔�3�wה�h�E<�d]�UPխC�z�/�b#I҇�(C<G���P��<k���SGO.o)L�������u�8w�����C�
z�Z�1e/��pײ{�o�gl+����
_H����2�e0-R����NW�9{��'��HO[�\z���Gb��v!3z���%�bK�;�If���-E��\|a��K7Xhx�-:��A[p�F@��&X/7'��w~5����wC,�5�v�j�I&�֤��vy��Ӑ�pa�H�8+򯚘���P����V���1�5*zC�!z�}�d]I�I-&�yiʣu��z#^T���?OWn܃oU��M���q���d�y�H�/����x�[d[�CR�;�͞�zG:�
�!�I
,]���p�;Y�*��|k�8������
�co��/c�0�U�����78���|t���E�e<
B���I���J�A�!�7�V�N��1�;e�}C�8Qeu#QA ��fؚ��~��sN��K�ڹ���쬕��e���{���s�X9MB���P�w}Y왱 8�.~9b��B���㔮��8j
��]����N���Q�sژ��P-`�8�9��^���L2�jw�j��pYG`���
������mZC��<����K�1����+�$���/�d5|��G�`]+��4X��.|cClVGa^������+�]���mt[N^˙ƨ��X�sp ����=K����l�f͇���C�{-��_���.1��*��uL���<C1P�f��΋�H8nc���>#Ɨ=9�o��������ҬCl͕3�j����tE�D�D��m����8��d{
�x,�ɧ�x��vΰ������7�X�֔��v*��P��Z�_]�"�kE���-`6���߰�f�6�"݁�+z\�faW��i�B��n�Ȩѻ/�o)'R���ˊ淎�`n��E(�zwQ��qf��9��%���c����'���Iq�xE/�n���U�- �����Z��qV��g�Y�k��/p3&$��ª�s%2��{�Z#��)
�Fg���wn�Q^K������F�`r}�4����R�/N��'�n�	`����"���C����yѡ��ՏJcL\?[&��:��_,�����ʻ^5�^]:���x|��̲52�/ce���;�in'G݆=Kl��}�Pڝ�t��Y\C�����n�l�����z=�z6nl�Jc�^�>ޯFN�Ĵ�P�|1��\N
�u���t�~��NJ�T�o�����󹩌�V����-霺��������w��E3I��=e��*ا|oH������$��}�<ԍi�`�� ����c�̎ơ���ר��:N��_���f�ʒ/��E2�/���}�v�ެo��֬�65w�NF);��;�y���f��	W}�P��.Tۙ�q��\c���v�D�����fV,��g��/z�zd�I��K�BXm�*,=�
N��Ύ
{c�B�א(4�~��oA�n���x�$��{5�B�9���~G���{N�j�{���z����g"F�ӛH1Ŋ����L5z�쉹�f��2<f-���.s�Z�����#M|GuJ��"���3rrֱ���v��p�&ek8Ŏ�D��:h(����kۃ�u�}���q
q[-N�7E��4���v�Sp
oِ����ژ@��@� �^P��P�h�@ן5����'���L�����N{��N)z�Y��~���4�RA��(��ώr��w�<�`�*�}�f�=�#�t���?}W�ĩ�;.1�GT�u�s�Bc �p� ֣�=lp��:,,f�*�< Vz��WT7�&#�f��ԣ��픝<զ�vSvȱ��c���0�6�Ǿ*�镵���<�����=.1F���*#�!���C�$��6�;ɫ+�f�6�,�S���=Q8�gH�C�R��%��y^��_��-)�0�^*�^�,#½2�ov:s�xkæ��3y1�w����P��8&�+��>y��_�Ɓ�����K�X��+��'K9]^��߹N�m���Y��;�O�鐿!c5�C�NWY+iH��l��S�q][�����'"�"���G��*҇��^˖t�����(Q�d�~��F6L�m[��b�4v��zִ�<�vc�����ȷYI�NcH���V����ɕ�Ԇ�n$B�a�v��]\޵מNW{&��d�$e[���ܞ��*S�|?\���LŌ[>���R�;���	ۧ�ȆV4G�C��yHSZCǴ��.�ۙ���v_%F��UC�n> ڿs���L�4.=��JCư�X�X��ͨz�a�Kn�����K�rK-Q/0-��t�T�����e$�4�C�q�O{s�7��ЖazIF],��G��E����K��92�&glK�|l�=�*2�̮�4^W�P<7Bon�X��6~z�Y+��ϹDߋ��d�8� z��lTZF���<$h�}��xr�H{�n��-��W~������K���+
�ئ9�����	��G�ᛙ=����+��5<h� ��.خ�k!�69}uIޮ�X�Kۻ͹��8][�B՘e���01�(tr�>��b���7:-�5F_/�#����G��᳇s[>�cbcp዗��NP��)�J��ck����8�w+��&������3�+�RBi\"\a��k�n�k��J��|L�Num>�2���2ޡ�=+vԢ��q����V��J�ౣ��\��S����+��=�fq��B!�*��"��U*�;-���Y���݁������}�~5~[q-�B��V�%�
��y�c��5��>Q����{F�GrZRˍj!L'�=�==��k讳�wo���.�oy�M�G[5�[5�(��L>�v�"���}��_���z@��2���g����ܸƞ�n0�ꙮ��_��ޒp��]�7W�K��L�SLv����>x��;p����g�d��J���e�A�q.5��Ñ}Y��c0�����wA�V�UO\�Zhƨ�7���A�5�SVq�P�T}y[�4f}es�f-i{ȸ��X_m��W^j%P/�hT ���-]aiV�/�,r���zټ8(;�b҇�#�!�L�~�{��YҬ����u�ny�)��Y�^��W  ?Da`j�K�qg6<s�U�{�~jg�V��H�,����m�0�yѡ��ՏJx���⯔>��#���M��3���s�t�
��h���q��i�ƦX��Ll�)��	��y��=(��^2������;��|1�M�G��CI���ɑ�M����Lybׄ��C�����c�]�&�wHr-,��moeۜ�(�QǭEe:��j4��'nX��'�6�vg`�*�V�j��|��38�#�zn�~��S|pp]�Z5�A��]�@�
�)٤jr�%T��G���>�*�{-ס������� ,E�)+=^��̗�3yk2��C�N�^�Ȧ�x�~�B1P<�{@6ٍ�O�M�ٳ;��iY�)�KI3P�GIj�^[}�}���O'�e}�I���$N�Z���I*,99�=�o�W�}�|�	��f�oԨ�G��Ͻ$���Ae}Ք�.s���4c��q�`Ũh�8��#��د��݇�}]O�Ӻ-}���� ��
�RgKO�>#��5�L2�s�Z�������?q�NwԮx^g�vwBE�:��r;`�bfV��s�X�tMlh��[�s�ۙs���Xp���[-LZ�ta�$ix��lj��j�W\(�\ά�y�m*� fs���(��Ao�-�a�8����z�\��j��=P�bҬ��r�ȪT�}��BJ�5ϫT��DnP�R�+�� f(�滈���g�y===������F�7�����$Uky��CB�zA���d�2j\�����V�_֫�<'�b����C��,z"���_k�q�^��<�Z�:V�z@�>�_;���L�[�/s���$��j!o������o3c�BWu��GR����$]��[d?�)��e�/�lQӉa��\6ޑ"�hZR��Vum��f�d�e1�����_Z�ս�K�pUt����M6��<���5��%��ڊ0]�,V=#ش���m���hۇ&+�~�3�L�>G�=���_��\�OUq��K���ޞ�l�w��b�b��f���0�c�na��aa�3�qm�tU�Qq���a�{����J���ʍ�����nzS�:$plgN$4w���w��j��'U����2�d�}N
[B�����q�z��m
�D9�z�
}�9�?`Nv�XU��jm�W�j�9��j�]86bm�7�5K����l~��ԏ�9�����i	zV@G�+�b�.��FK��F�g�����=����	�z��N$3���ٹ<)��
L�BXޞei�����;�I3�ٿ7�P��Xl�2��<"�R֑/݄�g����n�o�"w�Q��o�X�@��!/�!�Q���*o�l�79��lq�H�`��5��xV�z��#�b��;���������H�
<_����0���ch��r��1�#D�oέ��i>o�{�[z��u~��^W,{����1�6��۬�R����J�ɝ�&e���x����%�����G���;�S������R
���ʛS�f�ݷ��y�e�XMG�okiI���h�!�:�5�r��y1��E3���v�,��YU_־/��~�|�� �-+K��]�_�/)d@�Xu�I��ڬ��\�h���x��]`�D���Rx6��z�m���{{�n�mt:h�.|�)q�>2�qA��s�Մ*/lC$��Je��w�ʍ.�C�&e�O�/��f�j��1���RU��VbMV�;W����!�
|� ե/c���S��j�k8��%�5F�]��7�o^9�i��W,[�@�:�_Y��S��jI�~�'A��L�f��Ƶ��n�-�ϰ䓤X��$XЁh3a[�-�!7�]L�t�No
5�m���8�.�K`=��t/��w5oËv�Ʌbđ�T�^�Y����,�,Td���C�u+$`jn����5�_(�/wUE
0�Vs;x<gU��N`��|n�!8P�EL���{Ab��; �) �>$�����y�R�۸]�!� ���w.W�aQĂ7x]�u|��S�yё�r�;.��aէF��(((�|���C�`K�V���F�V�-~�=�����:�4     �I$              %�"��}�{q$i�z��+�K*��J[1۵2c��a�����,�{v�k�F��pQ�W.Gn��oV0l,}�;�$�.A�Mԩ�#����<1��<�ʢ93j��ks����P��&�@Ѽc���`��s������v��;��f���ק�5�j��o��C+��p�{w�e
5�|	�F�Q�[ؕB)l�Oum�9���-E(L�m�L�J޽�k�է��ô\."z�:�������-6���"�&GW%�U�^�\�Z��@�|_(�1�F=)����v�Q�n��eWe��,�V~�SUM�Q����]�[R!�f�Y֟G�$�F#Wa�#��@��$<��A�@����VHi9�+����Sx�#�K6����0]�<��V�����:�R%����"E�olԍ����}���AK��B �9����ނ �b��Tr��TL�v��1AAUe�P�b�*�DU�Rł�B��$l�饾�����QTU,��0�TAb�D�(���(łUv��"(!��i��X��b���ڪ%U*�Ec�QX������QB�II��J��CJ�f�b�UB�4�� �����AEb1SIC0X��*�V1R
��b ���y����f����j�cqnv�'ݕC�j��_E0�ܦ�F�R,��;"e�>��-2{ҵ�Y.�H����^�<��	B�|v֒Ǟ�ǯD�٭�O)�ܨ����d;%�x[������h�uӡ��؛��O�b�C�\}�᫏�g�i�Ҹ�H�.8O.3ٹ<|��W�3'$2y�U0y�^��U={.g�O�b�� �ÁdJ}kq۞���h�'� �̦��=���?_��S��-��1�k�!���Έ����������xИ�uQ�~߁Cཕ��kCƔ�����1�A��g<�c�r\o�᯲?��q�:���깛����4���ڔˣ8���Ғ���</Z�G%�W��w��؏}5B2�xj&z���J�P�AX �����%�<�{��Y��/&$���j�&]5Û�#��H��!C�����i]�^��-x�\H *��:P�$�YS�96ZǤ��F��]L���C��m�(��QRǒ�A����I������=^tY.[{��ɪ�߄��wL��7���{ʏ톓U�ۗK���A3Pp��%��7Q�����e������*]-��k����(5��G׷v�^���{cu�(�K�Ԥ�Y�.WT��_��LKϮ�������G�6��h�T��]2]F�O���џ�6�L�3h
>ղ�@��u���헝%{3'$= ���}���{��s��#)p(]� �[5�g��-��{�9ce�I��z�\S� ��Ƞ�\�ƀ��>O����fwq���yi�W��_�m��S�Cz�;����뷉$N�wl��w��}xxy�Z� :]A����
������ݣ���P���h�B�ݛ�<E�Lp�Vf�EK|z���S�{Oԝ�d�e�^�S���U5��� 0(S�崅�yys���}�̞6#7��j�%�K�-��,eHy�WX[�!�)ٮ�������������jn��i:%���	:�w �6���k:�W���(T�a��?�j�rd��{�9�-�M�|Oaw<UOL)�B���NK�,�v���5 	��!�x'�8�Rւ>�s�Z����,k�4���׊eS�ٓ�%Oi�F+wk��;C�L�C���]^v��ß�Nd�{w���g�B�����_,��A�g�3�˩D�{'Y�WM!ZyS�%�]*���'�,e<��-�G��Z�|Ҟ�_����ޮ�h"�(N�;�.��گѿI1$���ʽ��jB�j^eŞ�3��JCV�`�Zӵw�Y�ߏ�|�^d�-��4��*���<#��h������|.��]#���r6`�T*Ց����KN%��yo��"�д��ݞ��rnMじ�Ҫ0�a�j֞���d]�f�k�=�Da|߱2�#��<�J��n��x��ʟ�e6����t��]��2�㚳zn�=MI"�[wYDFyC�V������Jd4�����g7mڒ¤#%��!p���	;�{��<���M���@�߅c� L�K��9��Ύav"u4㩽3�o�>��~��`L���tu�ޡ-�w�R�y#�9���n��ױs�CKa������^�8���5�p�'�>����=k@�bU�p�,th�0�#��^�&E�~^�3¿����Bph~��+e���L���Eܽ�O���wI��|�1�1q�#:�#+�3�'��(}�&X�ĥ��LQ붥woMΈ�gĒf���R�V|t��慰c����/��Ӭ{�<�˔H�V���z*��p������C|�Ʃ{2N��t��C��͎69��_�5�~D׆5���8�
�Cֽ���ʮ���f�	:x��q�F�3�h��yj��FU�Q���Έ�/]NP=u����=�2��ZWc�V&��P�/q]yN���J`Ќ�:W"ޕ�0r��{��j$-ޒ�r&���E�p��keI�2��]�(x�}B}��,�k����D�Y�hɫ��&w'�n
A;�'��t��܆^�X�u˶+���Ȼ�thԭ�7��6�
�ձ*�.�ѯ�Y㶼z![�>�x{�j�-�i梟����=���>@�<��K��R�6p�kg�Q&��J����6dl��K-��|3c���P���R�q;��Β��x1���ә�N�O�q���J��{��o�	c�9�*Ha�͈�36�^u^�oI���k�C��|w�>��\��?�J��Z�j�EQ���o�sv+�}��-�7R�������~����WL����zl==��g���. ���ID֊=�e�5W�n�Ndc�ą�^�R��wr@�Ar��1,$��_s����<���|G�Q�w\4�l·�^՞�l* ��gD���9ϗ�{�+z�]�����F�NHGN�le���cS�f�\�[�
{$t�֠�i�:�	Y��n[Ѣ��3 -�{�����ǣP���"J���6�ĸ�7�~]b�L��\��{^8h,�c|x��V|�cpY�M��dv�[���iE  �s�n��w�
wei�L���ZZnS�7�L͝�"�����n-vA��o�r1J�!c�дGv�v�n���ܬ
c�1�ɼt���r��
L�� lKhK���{���$�s�W�����6k�����=cҞ>"���V���j]�l����.����t��R�竉�L�,n2�����������B�L�c9w;o��&;���H\��!�|`{U�u��ɻ���Ә�5�F�=-�u���=0ڤP����4aՋ�"�޴����f�ߨ||3�kh��~�����󹩌�ݔ�=��>Sl�L���֊�=���؁�h��;>5}�G=4���1�3�k�ѹ�ҷtd�&F$*�MrD�����W�#�x�.A��Yvԁ�����t�~=���w����<
��wp�&
z��C�X�U�7+�_bk�;To�/�h.���5����W����{\B޸��s��w6X�}��Ɂ���$M���s�8W,9������#�QB���ŭ;�z\gFLs��wavd#	4m=��yJ\�5��]V�����͏�AϏ�m�q�(dX]���6s�?i���Zm�Y~{uWft�,z��p�p�t���C�B��ĺpeU�;<����n\��!��m�bR�n�����8hbfV��WT�F����d陱�e�G��;o�PB�Ҋ��1`����HӾ��1���y��l���8�x7u��hã�<(�Mq�"��	g���oy��݆�џ@�`r&l���k�M|��^�U�1Hib*�@��\j�WzhX}�R����׽1��Kɚ(2���:s]q�̋.�n����O=�F�S-͖����0��螼��j�^eڼ���W��U/��o9�W
_�("��n��Bŏ�t���	`Q�Ս�:{a�WpK���}��/2�GN��9C�{�h|�]�ܖ��`6/��^�{TK7���֩+�u�,&�^
��@x�K�v�W.p|׼:�+���'�2��u�8<��h/(wc�Z�թ��b�3T��̞�F�vN���wU��05T�(�|����c�|����� �DSogw�1>�\i�ϫe��U�������
����^!�wx��=�l9tƏw���r�؈k��"ac#ǈ��
lfG*[���x�>�Xx����Fm%Pe��Fz<T�D���T^��P�S��;a��Q"Wș�yY�i[/�}2e�(��ץ�q������۟f�vVJ��t��\ad�c����2Cc,Qi$�Ӗ���a��U׏�Au�:8�t�(+5�v�@�1g#0F��lF$P͸1���$B����4Fq`s��A��;p0��Բj^�����#>�Z�[�}s+Q�3ܬס��I��(����kE�zgdZ�kc�w�Y[�O��S���{;V�h�S��>T���E.J1^kP�g��շ=ꊞ��5z����k�3'Vc���=4���Q�p:��	��ye�Ֆ/o.N��<�2*�v�iq�vJU��Nw�&��b�ї>�=)��\K/�U��wF`�ڔ�}�H��s���x����HZx�kb��_>���\R;v����|_�=瘯��f_�[�3���
X��X5f����[�����s}�cw��+��[�W�g�Ǻ6x=�c�u��:a�Y��~��Gح����@��Zb�#VL���G;/H���ن����Rlv}65�{]���N9�S������(�?VnlN)�?V�V�z7�c��~�R�蝓�.�g��\�9��}ʞE�6ڿ%�y�E���P�<�??c���6������C�]z����������:'�k+T�����u��%s��ּ��`�"l��e�@Wb�������[���9w�z>�{��2�'�rY��#���w|���$+��F�%��+dy��*Z�(�B�r�j�r�LȮ�,���^�'�j�o�Ptp������=ƹ��t�d�O���9�e)�Uy�Q=%`��ո�FN��y7��̳ͪ��ѣ-]�%6+�ק�"pȦf��D/<02�8��H+�-Ǯ�o+Q����Ә�XF�Aҋ� �%�m�s�})���V�pwP�Z�����d��u��%�%��M��6��꘶�i3��de);�B��2(����C���n�=�m���LK�F4e�kڍ1�dϺ������	�����m<�F�m)B2�V��gE =W�:P`�u�в�'�\&%w���yg��\r��5����X�n��d�o6��a5p��]�s�Œ��1S�U���2�b(���7��U�PM�[�n�wA�����Ω�k'wpkt��s�� ���C�%X��,o*�Ýʶ�+u��v[j<�Cڂ�K���4�)�m㊡��6m.�d���l09�xU!��y`Z�\s�2�"ZO.ev����3F���N��N$=��W��F��O�V)b�Ա6:L�`Z��Ӓ�Pf-8�\�N���%ef���wzLQW�ɭ��jg=�w9��^u�a�                      ����S;tJ[$��R��Ѹ��ra�]���YH9H���t�2��ݺ��Yk���X�Q�Q��=����4#��1[hfr.�Z������ ,PN��MtGq�ٳ��d�<^�{z;9a{�A�1�YQ7M����]�f�w�,�B���i:��ʛ�f�%E��n�lR{�pX��K�2����8�ॆ݅Lɘ��4,�IfRZ��I$�G�K�וƔ�'W�(ԥ�f�@l<�(Q��rZH��j��S8"r�����+�a�b\�&*�N �Q�wt�}yj��,�5�d�H%�D*e�H�@o7n��S���6SB?��|�ӪՊ�]*���-���Ma�8 z����:mFsn���Ux�N��83g=�������SgR*�Jx��Y�;����8Z��7΋�� �r�0l2� � W1;5���L�LgR�#��"-�X,AnҨ�*���X�V#)(DEQQ�C�X� ��VQ(椡U.Ш�aIJ�fh(`)���J(��̦3�
V6hb����RAV"��1��i�LUPQA]Q)XE��Q
�F((�b��(��IL�i��Ŋ��J2��X��H+b�����b�X*+"�h�"��M�H�U$X���"��}�7��\�u��f{���L+��-!֮x
�6��6�yR.�t@ͺw�ORO�OsbX۴V���_c&�':/v%;U�{۝�c�d��s.#�@g��g��z}R��M�B6���S�z�)��۽�>���*ǖig��4��U[=�Y�7us�����[���1ۆ�w{���Kp�1�i�����+�ҽ{]<�Qo�X�Ĳ�+5�GBNO�j���^��N������P﹤3)�sǇ&��N��L�ѷ~�U��4෍&�a�^�
ߧ���7��|/�C/���7~���>�-qg$�s�����.��R~<��-?[�o���Y�s0���V�j�tp���~��uۭ���̉r���('L#w]��gjb#@�r�H�%.'22�A:�Vݗ�3���I�6����.�B�t�j劌�]\Q?�h?�n����D1�����)���y�Cڭ�y��.n�.Yk٭:ّq�4�rɘi�/���м��ט��ߗ�7��}[�
n�v3��䪵�yL�*v��]��������� ��\�H�Bܠw���Qk��z�/L���v��W��������W���֝�YL�Ӹtfy�T]��{��H#��[\�^��6%�m�tA��u����{��sW�N�����c�	+��^z��6�+&�i��w�oqY���]lo��y�'
{�������m�r�*�fQ�WnZ����/���/�v�\
}j�']�-F���mݽЇ��Ԝ�����5��В��f�TG�e��I1(�i��{;���4���y͗֠$c����q;���0�;P���O+��9�.W<�kb��S�?�TgG:t����l��z�§{��u��<�U�L.&��9�JH�3���ta�����|'�$���Uq�ֵ7��܁�l����+͛����(Lڒ�忼���^���^;�旼k_y__�_.O��*���|+�t�ǷSgL�]�8�s�6'�h��^������q�ԜlKh�E�V��7S���d�Y���2��N��_)\(*9W7�im�ʴCQ��3��]9꭭.�X��s,o݇;�xFd�{~^
e���j�Q����|��͛�SA���w�\�[����������;��gZ���}�m��A99m�_
�J��D�����y""�R[e:/]\�Y�L�����O:5����a����_�����(�x�i��K��C��=�~�3q�R���5�{�}��57쳼&�8��㞮pP�xͬ�9j��/���d���;J�i�{x�mT��i�ߖ�~�ˡ�}ak\ߦ������I��~�a5�q��6��M=9��'�o��_v�ך�tL�	�=�g7�s�ڗ��U�n4{��,���G������S�>�j�1�?B�Y�Dm�5p4�	�ӳR�2�WP���â�juwy���'���+Y}�t���Q*ek2���ύ-[�SO��\�ⳍ�SU���zD�Oe	���+�3;z���MUۏ�w���� ����؂�gR8c�fм֚Σu��]�gI�Ie��ٱ3�U`=梞��|}1��}|~����Uԣ�O�&��%�I�z��V˝^�x
T�'X�J�Ц���u��xp�tr�Y�9����V�p�9IN-�Д�J�l��SF����>Ew�z�L����W��!��9�l'��֡w�~�������Ѥu.��z��/��s�_B��cW��e�>�k�_w�_�o�����jե����l��8�^+d��8�������N� ��D�YJ�ٹ�Dc��k��x_�7�����K~��_��U���-/m`UJ�;'p5佢���	��[�Y@������7�����Өmz�_��.��%��vk*(N��'���vǑ��r�����r�>֐�gt�A�77������Irs���S�/!���WGݵq� pC�H�]����;~c�&���|z�����S�c�
(�{z�7m'�|��B9�c~.�����g����,��ni�������g�sӹT�m���T��>�1�o���b1�mK6i���w��ly��}ݑqߧ�dZ�j�矏z1XT�4p�(8ZwM��z�v�2������t���"�~�|w��OT�\N������5f(�3��.���9�(�Z��Y9�TpݣB+8���Û�e�;�V��T=�냜 ����#��~+J����Z˺ƍ��y��
��"[D��jM{hu�5f�;��wH�|���D�Qj����8�1=ܫ�Ԗ��d��gh�[�����
Ï�A��+����~�;�ʖ���E?n���sF�)��n?Y\����^{){�O�~��=��*E��v{�����e�iW�P�c�tto��Mg&��0.c;���_;J}j�O3z�{���kH�����N�y��̝��u�.���n=h�[����3���$\a��i*3���2��&B7�}��kS|�g�����	�Q������DVZKݩ�k���{q=�x�H���"Gޘ�� ��\K�(�����K�ww�Wعi�!���ץ�S]K>�4�az&�~��$�}��&�*ŷo��x=��i,�Qg��kNe�ͣ��0��)6(����Z��\n���ٝH��5�M]��%H*�v��X���!P��}�)���X&�"���8Yʰ>���ǌh�5���>��f�ɋ�S������{����&){���kU�J�zׯ\r{�[�[�}�G���[�֓��2����-{��.���۫�5���u��HU��ݞ�pt�ٷ{ET�������K���xk��=�</Ԗ�[��O{w�R�����{���=�I�[KM�}{����{7g����E�4���p>�k�з���Z�%ز��}��ɿZq<q��g�=����{,�F�e�JG{s�
��;7��yŉ5��y-���Dإ����n�64��6��lz���Ő�w@V`����YŴl���7����R�l���޻2��⺂��0��C�[H����\�Z�՞��W��+7�c��?2��nI��vMh~z����J���~vs�kO�F+Ѡ�A���=����Z�O?c�ܜz�Z�P��؟.c)QE]2G�d��H4|�Wg��Ⱁ>�\.[�6����\��t�ԝ���S[>x��d�r5!y��{�}�z���(��z~�yeWBMj�7�<Wo��+�>^Qe���]G���||^M�d��:�E&tf�s���c��U���^g\ޒ��}�V�r�A��yn� a�yɛ��f$ʤZ�;p�JOoכ����	�O��w}�w�(%Xn����*�`6�kFݡK�*uL�$٣%X弓�Q�D��ܸ-i�О�p���qOz���������9	��U(�F��������Y�*�M�ybM���U>�2�j������}�k��\�>�c����N�K��4�#����=W뿥��]��8��F�!��|�����=��S�>����Qzt�oMU�m?c�f��`��T!�OMs�	�<�M�����S�<�3��'���z��s�i5���3�'n���=s�i�>����o�a.cٓ6M�����[Ւ��]���rq�w�>>){����R�[�}s+Q�'����)�#��S۽+j]�3�`�>��Wf�+s�����C�ܡ¹ϝ�Xv��o��333V^�V�Q��,��(5�Y��kuT�s@4q�a�s���a��Jq����@��p8�85.�w���Ntk�]��G��%D�ܛ�ͳ؁+E*�Au���~,nc�BS֨�J��U�=[ז��\n�8C��s��	4�X��q�<[��V	�@��$��f�܆aE�c+#F��"U����t��';ַ�8غ��m����DD������%�����ܰ�Ew���U�	����Ef5���0^�.�����E�㨂K��O.fR�!Ǧ��n��d�K"�ͱH⩼�WgߞX8\{�z��@i�
݀.�p̼��-���VkocO�D&�C�&s����l7d廛��ьh�!��LO(���W'A�# ��,�k�_�L�����&�m
�)�<o �����cL,��Ӷ��w�h7�򝛅� ��Lze<��ܫag>�$�U�"�2�a����1�G�S��c���� 8                      }|��=-�"�pX!���S��-���f5�ְu�}̨V6��x��z؏E�_�}���-��wƍ��hD�|�s��P'��1����b�(o�]s��o�؍�mMT䒠ά�y�EѬF�	�84�|M�J��R�;SF&�*Z<cλ+�`�x���7b�i�[K��b�r�K��hon�L4���R���k�EiH�C�,��!/>�L[t6�v� RT����ֶ�ٻ0.��Z'��H�F�#e����5�Ai��sK�t�Σ���U�&M�,���5Jt�
L"�ɭ���Z�ʃ6��ۼ�%g>�;\�9��	D��uX�g����ɼ�G9��mJ�Y	]����FĜQ\'j��&��V8@�bi�AՍZu*I-��c%6���s�Ǻ�aR�f�%�̡���*J[pmn�|����&Ud���F��!�Sh��
U`Y�K"�U�Tb#b��DUQEQA4P�iA"�E�T�EU�H���1�(�*�\�.��#"�����PH�0R,�Qb*�"*���U�n�*�E �ET�J`(�# �X�b+`�U�((�H�,�E"�EJK�fb�@QAb��DQA`�`*�)����aJ��I),�dFA@P��� �,H+lc�9�g9����<Ѽ��׋��<��fe�#et�9eu̔P�4��Vb�����7��}�����.�R��=�㖬e25���\�����T��:9��n�r�������ҥ������1�>��$��ǝ�ӟk�����E(8$^�A�w׮�r��S��;.��fC��^��i�~Xw=���֋�u7�(��f��˼ó���_jS3W��YZ�f�ȭ���B�m5�z}�]s����i�ՈL�Wy�.�{����{6�TT2��/��=-a�����I�s����=ۍcw���7����~��suO�/uN�M��ܝ�;G�Q���x��u�gr��fӉ�禹���ⶹ·���}�$�����n��5�����o5�h0{)zU`&���y^0�-�Q�_�����P�Vz�����G"�Sc�dD�JK#f��g:ۨ�6��i��@�m'��®3�w4|����{��菭v_'k���*�r��=�<k/��c��`*ɲ.�Ȟl�Ti�R�z�w���y.4z������V�y�}���o��G�kc�N�h�M�w]�.:�Ѝ?N{f��Λ$��&U��w{��hy�c^�Ҳ��\+Jn5Nten&ދ^�|�n��xz3�����^PN����e�e^d��it��=�js��9��j��^t�aj���|��9>��.��R��D�Q����N�P�Re���p?"�K��Xί,���e�vʼ���}aS�D�� �|t��<���i�&ԧ~�[�⓳��I��HM�Cu�l�3�%ֳ�7d�����U����,���ͥd��#�7�/�5s��/Al�(Q���*��8Pa�y��o��k.Ы�������l�"�?3�Z��Rj�d���������W�V%�]\�ɮ9���o]�g�'�y�]�خ����4��z�|������C��z���r>�]c�qOԩ��W�Z@�m|��������$e�W��˵�������\Um�F�?wOV]C����Nhf ��ᶷ�Ooӈ�gbZS7��¶�ٕr?���#�����r�NʦM����)o+|���l�4����7�p�R�t�k�B�{��J��v{o���b1�C�9��KS{�z��=�d�'��z_���a�j�2-��":�?o��ulF+D��F�_f��(e�d�e+��%����xo�V��ho�I�g��,>W{�l�mL9r���Ɲd��|zβnWt��zʹ|�I?����|�Y�]�#�en��d��z���3OD�׳J�S�v3}:�>ς���3���kfz�g(�#�K����*G�F���M~�k����3��&��#�����I�y��\A����/#��5��]��V��؜�.����	�$�;�Bx��،-�}�Y'�=�ů��:r�9�%n=�� 鳡MN�^�֒E���Χ�ã�ǚy�<�N�S�>������lS5UT�S�p��`kF���z��t�=�ȹ�_�h�ԓ��M���ļ	�x�=������r)TWܖ4\e�wj����d� �/�N�I'*%v�u�ᗱn��:|Z�ȷ!�ܒ$R�I��.�+�o�0��[M.u���lҩ�w��CFRu"�wg�#���Y�<cS�5~���+jq��/_sm��%;���V��؍(�[��,h�?l��ԝ���z+.Z�)�RH@k�>��3��eu��}s53ܻ�v�`b=�}�}�#���5�lT�`�[31�s�V��p���\MT8G#aZ�^����]v��w�r�86�rR0�V��k�]O];��v�[�۸��:(6�)���>n��{_���/�W)�B��%\l�<�2��o?n3'��R�`d/L�^��9^��L>g���/;����U����&^����U�劶E@��lY��6�si��&N,��x��V�<XP3G�t9����ԕ�c���wMST�����qL[t<���|��zyï]&�7{j<�vʹ�"]�8vQw�8x͝���u�����+�ߢ��i�wM�#�<���[���^~��ҳ������>��.ԧ�*�r�wqe��c���V�N�`=\�����F�Bw�2s+�nrYe��W<�sy�o��K��s�s~�3��5�}����j�Nb~#%���V;�@Ws��Or�}��f�g�c}�Lj���y�n�N������$���Ms�(��g���]�]�����y�I���w]�:��*g9m�py2�gd��XPp�ݷr��k��EK��}�VCތu$5�`��^e�]y8�rd<�%(���
sr=����uc��]�}ʁ��07�s:�,�D;b�mflW�G3$���v���U0����btBПQ�ۜ��Xr���4��ug�P��1��w-��������R���s�$�^*{B�����z�$��V�M;p|�ה陒TqC�0�_�Jڐ߰:���˔헔�mI2�F��j�V�{�H���:�;}�(�)Ʊ��.�Q���?��x�1XΉ)6t�Н!
��1-殻;�v�Ksp�y^,�Z�Ƀ�*v)<��o>�<獕�u��ܮ2׹)�`֭��T��vy���y8j�7�oM�^U�b��������l=���>䃞�ƽ��<��뮚��ɻ�Ms1��_���k0ۅ����S�Yw_�ܧ�AT^z�:�p��8sY��g "U����J"nN�5ם�<�֏+o�\�1���ue�ŉo�j�vAß �Ѷ��Wr���[J�s�lۚmN�B��?Vf&Y���J�?2�罞8���K��e��܎8�8���;;����{M-a��*�	I���M�̘F��:�<��s>�k�ږ^�.���� =�U'�!�z�]���P����� ���rKI9L���I*ʝ����_��a�}�$וs͗��&��1뇝
�<,�
9*۬�v�m��Ox�{ȕ����\��.�����8���o6梗z:ı��c~�~��}�*���uM�υK�^ntZS�t�?9�=�苚3{�&p����b�=��S��X�����u�����\�Ry{�IH�=L���t��1S g���:)f_J�h��؊��~�!�W�'���{˅�B:��y�t���m��K�qMsMqھ�cr�y����N���r�ƻ�녽��f�~|ޏ�ZE��(�j�_���uKYd��D�88�fw�R��}��ԏd�ݾHo�V'�c,͛4�j=�8�-�=���t!���{��$^�[��޴}vǰt�)�W���p?<I�+�"�nr�\�T��'\O��ԨM�y�����q�5�(W)� ������wV�����?l��ԝ���F.u'��Ƶ�k���k��G-�R<�D�j�~���z/y�(P�B��ƞ�vm���s��1��˞ל|R�$��m������KF�z�\sb���|J�ފ)�<����:�u5������7W�wk�5Q���'Qr=�+�I�#�{�83T+"�2�j%e1՛{0\��-�2I)5��A̢/1��W���a=�'Abqm�j�aB�@A%*��Q7�j�$_��;�ӹ=��+vf�	��=)��hWyg��7���oԽ�Ǖ*�;�,tKGn��ԝ�8.>����k0߾�rh=�i��U�4s}��ɦ�=��yӧ����sѮr{��$�u�1�w��X^�!(���G�.�w��輜�RvT�;S���N�.�-t�q��v��F����|/�]�O��oy¢��:(�c�)Y��x��O׃��kU{��dU:��o�l�H��=�&��v���y^�tGK�y}%���/Ll,��+��'���GG\(�}y��E�$}���=���>}�&V��c������P���M*EW�B�I		6�?�$���?�!D�$$$!�C�F̇�8X�\(-cVn�^B�k��\��Ld�D�J 	! 
B@T���P����I$#?���Ʊ�$�3%B�悠|H�HW��?0����e?*�3B��T?��P�I		~BE�:Bs5��}N~�x?���}A`�x:С�2`�}w���!k�.CA���(5����
(���֤��b����j\5�HHC������-�>�9_�$� ��	!!�MI!!�@���Ic���f��������\���?�%��`�����O�O�`>���4}ߺI		l?�C����>��Ĉ�ą�A�BĐ��Oԗ�	F��C�0��xC�`�HW����%�$CO�~(}0�CO���,� ���'��HHHA6}*v$����R�ﾄK�BBB��lKI'��x%K���*�`��M�\����������䐐���L�db��}S!�@������I��O����1
�1���S��}!��}s�ǉ�� �?�~���(�?�~Vu��ҏ��FQHHC�*Ft��?9���!��>����62\(���?:,N��
?��W��?g��.	�?�>��6��[�I���A�������	!!!��2 ������!����&͆aa���;���
U!�	!������������	�pR�j-��~O�J��o�وPH|� ~d2|�I$��2� �A'@���4H��6O�] IT0T�&�I���2`�|;t��4��@���	��$-$�eO�%�U���sr����� ��~��?��$>���n�~�O��I����~�����O���3����}P��>�|�X$?�T������ϸ'��}���B[��!���!�_����HHHC�?���|ߘ_�B���~��!�?���?�?�����������:O�����,|�~�ۮ��@�CPZ	��.1�K?u�|�~_��?o�2?�~G�����a�CD�п�~W�!��$$$!o��!���a�����6�}���b~�	���	�X}�(C�_nk�ق�P`��>�҄d	!!�d��������C�H}��?o�|�?A���	!!�O��$��&Ip������b9
$�`cV�����l��Ab �>�'�H~>>O|����H�
�7��