BZh91AY&SYW+��M߀@qg���#� ?���bE>�     /  <O�     �  @       4 h P   [(  �     }�G�iV��`*�h�R6�ŭ���)�Ʋ�̥kE[2UCl���
�F�TSfж�chKm)��d�$�k 4ͳa��PZEW�o*!P�xCU��B�Km%��U���X�A-E6�[f%�ؔR(SKKa���E�d�Zd��mUif��j�U���X�i��M �vαM����   =�G�O�k[�h�Z+m]��V��"�UV�Ov��������l�[�¸�j�g`=7f��OU�oJ٨-j6���F���ֽ�  z�yPuF�pfv�L�2]ԥ]��ݷ�{{�{aR�۽z�޻j��n��Ow;��=7<:wm�oW�=J^�k�-�V�3�+��M�P�*����X��ڛLm-J�RATg�  Y��T
�3�k��mmJ}��׻p�JT�C�!��t��zw����57��zR�[i��&G�(Ps��yJz�K^����TҨ���yv�׶�x5KS"���ikE"�N� ��|�zj�I����i�U����|���
5���꯻ʕ_kj�ov��+A�E}��T�,����4����[�y�!+�]�����)MO|���ցé��IKf*E��٥��o� Y�©���Ϻ���P��o/�}�_m=:R�g�n�i��SY�}��RT���}]g�M/����tԴ�����Q%S���{��֔���y�*�e^zRʰ�̊�#,�T��  ;�S��i�{�;y-��w���)�Uءw��=
P�w����Ji�]��u�kf�y���*����ooR�P�{��/XF�ݎq���UK^ޱ���J%Zf�Hj4��  O_R�VZ]�oNoekmM��t�Z�{W��Ҧڷ/m�Km*�ճ�ޏxP
���Uǯ,����/^ס�ty\����t�  ;ܽ����
[6�hcE��_   v> ���8h4��ptG0n� �m�]@�r :�7� :�=5�� ��ゴ��x&�I QP[dXڶ�ڷ�  wo 4q�� �� ,F(
ݥ��Fk�u@���飵V u�=^.�A����]]�Uno%Em�2�U��V�Q�[�  ;��� �8P�z��@==�j��K�� ��t 9�4\��(�=8 =�x ��  H  j`�J�&&`i�&#��ъR��1b `@�&��~J�� 4ɠ @@��	*��      d
��xj#eCA��h��	SS�	����ГF�� 4���_������Ҿ�}��ɛɻɺ���u� ]���N=�r;���ߑ����|n{|}
�����TT������ ��������i���?���}�UE���W�� *+�g�?�E}_������@��1��� xH � 	���G���H�����		�%x@%xJ�$������8B%x@ �!�p�1�8J� �$xB!xH����+�G��G�/^�!�@����Pġ�P�(p�8B!���$bP�
p�8B�$N'	�C�	�@� p�8@%��� bP� ��8H�!N�	S��"p�q�8@�%	� p�8N$xJ��<%xJ�� p�8H!���Dĩ�T� ��8H�!N��(p�< N	���P� �8H�!N!�E��)�EC���	LC�AG�����DN��$8@
p�T� #�C��/	U��'PN�$A8B�p�W��S�('�*�	@N �!D8@ p�D�)�C�	B!T8B�p�P� 	�PC���	A
$8J�p�������'	
� A8B��� �"��_	8�P�
#�S��' < 8@����*!�<%Q8H�p��/����X�	^�����	^	^	8H�!��p�8@!�	^'H�� p�8B!�	�!�P�(p�@!�����p�8J%x@a ��������AZ?_~Eڊ�*`��h�[R��7�
nLXA��R�;�� *��sv�	�:B�g�����z^���Bm��!Vp1�;!��p��=92L�
�g[��۽֬!�X��bp���q��k�H�m��x�'��<���wH����gn���}����4��a^�vN˲=��$�z!��ӹ�8g@��,�TbhS;D�ø9h�&t�=ñN�{0?�n�;��
tln�+YN��Ee�`�o]e+������j�5�
�䈇��>����V	�.A(��n(��ܙZ&!��$^�n��69��ĵW�+8:4� ����`3Mk�K3��"bZ8C6�P�p�uH*ű�r��+��ܳ��(q���ѭ�*�wkX�M�]���O8��Hh�ikl�o:����.lS�������i>A������i���YXXWB�-i�M^٤�5�h�Ś�x$�t܂`}���;���t
i�]i��#V�au	�����vd,%�6$)V�$��,<��������㰸�Z�=o]�ک��6w6���~��t�Y����5�
�ͬ<�vPn���Q;�i����@��I7,�s^��[p�6�n*Ӆ����nSE��]g�L}[�-���ͽ�p�tpv<�l5�SI�x.���yi�U\/l��+;9����\뎇�orO\�y���˲r/�Hz�%u��Oe˛���Ed��/`�ݵ���/qJhNeC][�X#�l��N��1P0ʩk��i��&�Sf^�V�#�鍘��#���r���}�R���Z���tFMW5�h����佣��\�c��Q_	�v}��N��xC�A��f���:b4����NLt��Y[\M鳾ج]v\f+n�뺞q齆�t�+�,�3v��c8�O3���{(S7+�&٫'�@�FwW�]��;nrͯ:d�7JtĦ��Ce$�����#@���᛭�}K}���'Uq*�����#�f�s����]y��Ẏ ��������t������]�9Ĕ�*�EM��I�q���W��TE��.M��p�;�v�u�Z靲�}Wq�)�b+#�"%��;��oϳ���o+�A�c΁G��0c��@ˠT�Z,@v�0�f�Ov< ��c�{	����:��g�5"�3�����W^\X���X�tQ��'QRݸ��q�%�ɫug�S����2�-W��7��2>�$i�L��씊4�V� v7����`�%=::l|b����ǻo�*����
�P8�wXYW;��E��"vt��X"�Z�a�T�t�>t7�sIs9�V�#��K-��8r���ph��{`��&5��׳'lÝ����-�.+��$�S�(���z0x�Z������9w�(w����5on@{"�^<=�[���!^_C'�S�gs�f]Lcݭ<�z�-&QL6'���I���F+t����7�u���Ɏg�ԍ0VY�y�<j��vPc��E���Y��U��}{�6+��eـ����y�/�9�j��&�� Ps��1[:MD�1%�{�t�x=��@���$���;!���gp��b��z�<.>���0t�旃Onr�08�p�&��Y#Iz7�NpRWږl=t�\���η���d�7��A2	d�@ɸ��Z�,N����3N86c8����6d�9&�KP�I{��35l!�Ձ˛t��؈����z�%>lַa]���R�s�>�+su!GJ�Ӗ���]���tu'/c�,���@�NG:Jͱ���j;zհ̼�;���Nm5:*�`_���{�;�10�sx5�����谆1l��0�SWji�
1�nOA���{c�k@�Ce_K�U�*9�Y����X�ل����.�Cۈq��m)E�Y���3N�lg#;��}G�%���Ź��>�k�F5Y���eyWcե��3y3v��\�y�o-�Q�^HJ��� ��ʅ׳� �MLF��`[���y�f�ðL�v�ø�k ���*����v����%�ۇ�K&��,�:0]y�o.���>���2���gdg����^�f�*-��n��^ ��]��xBxu���sj��>�J}N�
�ף5Yy�,�p�JF�`k���ܤ ���gB�]7�s��{�5��oh��.��rF�����^ң8q��84���{����lų
�7V
��]I�����p�n�XHsl�ǸɧHj=bl9h�wgk$<yt?�]���A�
i]�h�rɜ�s�d���-36�ɩk�q�C��K�U�̔Ҵ��Y�d��;0e��Lw1��R��>Ф��İ��ںeSj�N��2���h_>��nl8׫��4� �*���ʤ���<�ab�-k]��dk��ܹq/��N�*E�ؓ�E��S��.�����S�/�^ �#/{-�as��<{��q��`8D#)�wi�1�I�tI�j�r'K���;�!��tu��:<F;�67�s��s�驮j�n䭌�si��5ڢl�L��V����w�<Mv��
�yb8z9�XY�mUۆ�0ǣ_'T #(��q�k�d3�o�s�#��]=#n�ǎGY��/���  O^=��(��m�����ٶ'L�ά]��jA�������3���� �/��Gc�6� �&���u�N�H��w���j;���D�׎4X���ٗ�j�@绚xb#)dƴ�;ۛ�%�슢��9���β���c�-Z����u6�=Z����(�Ͷ΃�5E��l
[�Κ�T��cws�s��A�w5���Xf�דܢ�qa8Z˝n�m��RޅI��H��^:�Z���9N��;Gdg;r�
�ZGe���6o�M�Z���X��/����y� ��V�y��6N�d�a��� �`}���9���1�p!��;PD���z�7t<Ҳ���4꒪�۸n7v�����B �q�&wvZ�L%zr�w�L�`]@`�[��Eu^H��~�h춾ڠk�r�Ue���م��޹�Y7 /����-
l���rټyt;���˞���O|g%�P?tX���rQ3V��Z���H�4�7�r&�nkо6f�{Kզ�J�+�dl;Og�Z16L]�bZ:������A�U34�՝�Z|�J��<�S��v�@5�{v�Ѣu���Q�G����AVD� YG rf֍�R*�D��v��~ޯ�X>1���Օ*<O"�⺄λۋ7&�!Q�oޛf����ܷ�X("��avK&v�1��.*0z(������T���y�%��w����eWD�LkƉK�GR+{��S��.ǝ_Q�cŶ��\�Ex�]���2�K���D�ݻ�uV��Q���(p����ܛ��ww	g{v�6.�pv3x76�����t�OuL8s���^Ap����-�D2����/�Nn�4oe��v�r͛P�`٨����.�1��r��#:��I7s����E-_n-+4�Q �m��1^z�e���B͜.�W7��hր��s��ql���H��Gɮ$n���D�'CgoH�TM�CξXl��b���{��U��9e��
����s����(�U�x�gC�'�,٩aэ��t�ͻRn���I�Osh�'.��;���fg�,�{��u��F����ݗ�����iVd�Y����یe-��	���������3��tb��zG�o;�	�U�k��f���)p֎�T��[�L��6N|b�3�Q�Z���`�٤5�a�����=ӷ�]�����*3^�{�n	珱~n��ǐ?)ۺ�"WB�N;I��.���fۑ���(�9kwV"���eMp�\LWd���$��lH �6��e��ck=Z�Q����uX�R�Հ]5�t�};f�m�"�8
���B�
����N����"L�ܷ\�b�!��,�:;����S�(�8�D����u0���yl�!�

0�Z��ܛ�7�V6�7�`�
�f����ʫ߃��A{V�vo�]��htf�ޡtm�{z��zo@�%B�ȧ-����h�x/��Cq[�C�T�+�sn����+�V�.�u���tV�Yϐ�9��uu�xI2���rp]Ǎ^����*O,��d�#�Lȷ�;��ӝ�d!'q��_
�x�M����vO�j��$��U��4O1{�i�8��j�ض�8�=�����6;�q�hf=�����;�ˠ�Ac�跱(4r�ۺJ�Lܓ)f��\��MknU��� u#�X8\��|,#�/��UͨN��)*w]�𯈿N����>��ϸ�LZ�=���[��u#�)�/�Z�S,�U)I;�fp�_f�c��*�EJ��aT�ڶ����L��f�'v�qC��*�è�]���v�gl�Y�1;��qZ���� �p�ϯ^q��A���4U�eU�7I�a��J�"�ި�<1n��H�S��nT��7J}É���sy�GsͶ�١���;8��.���v�����Ӝ�v��׫e/��{
Y�*�d6zb�Lg93�K�!����L�+��̬lhS8@ ��i�=4�0��2�����U����;w~\�Ǝ���hj���t�b�$�7GқtLvj(��v��3��O':���6��y� C�pIp��e���r;c�ye#��No�r�ɽ0<�kp;b��'�R6Ah�H�o<�΀����e7�#�k��9�%콻�3�ݸ����Mod}�T������]��M���*��n�� z�oN{�A�ve"�D�WD\ջ��d�";M��kܥS�d�;�N*'09��pm�����P8���f�*`#
��η��Y׺n�7������]�.h�*f�����
6�0��0�`�7!-�WV�]wA҉��FR�����cs��"�]�a��]4��ô�� ��{�
��4L����}��0��F^�%!Q�포.��hnXz	H#P��N;��Ѕ�S���,����	C%n�ì���������&�`���K�|�r�+���JSu	��0�'�1a�����Arهw��Z����i�����ò�T�"���[�8�f�{���I��Ѽ�nLP4�,cL���HR��=9�4��1�v^Y�j�(�Z�)�>ݱ��}p�ޔ�C���vX�6f��{(������7yQ�S`�'i����Fs1��^���KY{�X����(oU�"P�
���睄�f����B�\Z�.#�v�	iW���8�P��ݜ������#�4�ӷ������# �!�v�əB���-e���U���Pu�d�����ww��H%�Kps3�P��n�i��3'Lc��y�t08p�\*�@��=u���Z��S����i��Lz��������u��w�lWx�.�J��F�Vdo,�;�uG��7�.b�rԁ]$�esF��0�]WX���Y�6�u��g(�.Җ��"�GL�n��:Km��ST.5��)��t<���&qk֬��g32��`=tY�f�웄.Q��th	�{7�����:�0���;�C5��V
�8��>8A�v9hm�HA��j�Mb�)�M�5s(=82�
���y�(�rj8�'�L���-E�H�u��rr����e|�8�D�e=*�\�T���sq�n�3�l��c��1��/TŻsb�]��Oa5Y@�:*[����,�:3�rkg``�ȣ��:���9��k�.�W��DHO)yL����ӷh�%	�p�����$���p��|�K,�ہ$ׄ3!�~ո���H:rK]�tyz!�.ø�r��5nwo�i���5�tJ�|�9�S:��A��Q%D�F���ߕ�G�J��Tڵ���(�j+��a��޸��nv�H��¸w��Auv��tR7��xˎ�>�퓎,��]�/$Ć�{��A	�/'-�L�x�M����&�i
)�|K�c�}8v���C_�[x�wm�6�:%i[`�f>���q�6��@����i�Ҟ�0������Ir�N�B��v��y5]˗5�we\�ΦA4�.cu�Ѝfgl��bq�j�V<�7������ӷ;���,*oƠ�c��� ��x��j��nSN�ֆ�
L�}5����gQ�`��r�R;P.^�KWK}�[��8�����QT������P����p�	�w���ٷ��L���ӓ��+���Ż�Sg#��dFe����4v�2��N�Į���͒]�6Dr�"<��揔�v%m=�t���.h�}���r)�z�B2�m�z�FM4���c��f��Û��M�}��ǳP=�o��8�ݫ-ǽf�8�QH��%�X�-엫Y�'b\hX��wd����G�^T:�'p�k�(�����(G;�=�g��!�Tb_M�	.*�I�%Ͼq�~R����^P}����&M�b#�j�ˢq6�V����/ַsYy���d��]c��Џ:vJ�p=T��cN��ך
b��'uf�@�J�{��9�-�3t���vw�6��jb<Sy�Ԭ%]��aK���׻q�1���]�m��j��#���t���n�y]19k�4���Ϻ��bƆ�K�8ށ.� K^n���:qͷC#�p��Y/\/	Mqѳ��U0D<ן�8�֢�u����|��$��lk��(�}?����d�sst�k8������i��w�[�|k���9t`�s��b^�dO��������0����h�,'��9ڐ���y]��+��X(Ozf۹6{���K��ֽ�8E���+�i�g��ף���%�=�|���f�:H9PS��	KN{�0����}ϦM���б�<qr3��|��!���A�*�i�ZaM]���%���)O����[�B��d�7���F�:�n0;�K�-�w\�[�g�9s��$�,���^ѕ��Tbw�+D��"�fvw�h���LZ99��s�p-���Eg��. N�%����d�o��9����1oZ��B��w���g�F�C��s����1��g*�PR|5v	��嶦6���:�2�����>�Cm	�l׎fE��nN�t^���l�0��q��{ھ:���2�$^";�e�'��t�5w`�yC��r����K�ܝ' ��{�[e;���O�x�
������Ӕ�rb�|G���?�r��p�������u:�c���0�|soN� �� k��D�U�9,
>�nj�9`x*^��d��M�Ih��b�ח��s{�3D�N� %ܓ{�jH@纞���H�� c�1��Ws��p���|�i� �@��ܯB2���qU������x���}�xb)Vc՘�Hn
�U�\s+S��xY��v	x���)�}�uĩ7��J��D���'�h<����tt̰xQ�S
5M���4�~iu����K���ϕ�I��iG}eL" ��U������Q]��[%����J�+;j��ҥ]��e61f�n����U��u4�2y\A#l��y�����+/��쬙�f���f�'>�$���_t�Kjҋqu�+�]��:	��ܝT��h������N�׳v�1g>��/#�u�������__�v,��%Pּ��b�p�h�ktn�(��t�a��R�����8��7"+.�$5�b_�矺M��p�8���䒾�6�\z[ƿE;��3!����x{nY&�
a{a����=G�[��[ʩ
�»7�O�h9K�q4��{mnt�%����&�8e˖�Ί�1��V��Rt�%�]޷M�2�
c1"�:\k���x/z	 �v�\��W�>Y�_N�i�/'�=�2Z|�9<��2ya�9�&��s:�b��l������j�1ؠn�5�|צ�����d��w�^�A�ٛ�e��'J�� 7t� ×=�nk��;����=@YWA���{gY�L�b,�8��뫗
�G����v�,�R ,��s/Ž���S}뙦,nTgXk��sRRi�*�[��g��T��j��H�͋`R��xw{Y֓��׮��es�d:^j�%�n�7a��09ۣ�|���^��Mi�p�l�6�e�X�Po����|�eY�����r:7�ٔ�i۔���gm^�կ�Md<��9v���Y	G�0�\�����Py]v.;���b�P�K�$2�<v����l��Z69�y	��u��yx,P���u)�]�D)�)g��}\��Yyee8��Tu�$[XrĎ�vZ�ٹ���RH��Y�n�:͵�5���sL杉��������N���X�֖M~� ��bi�>��o��6m9�S��L�a�Q�R�L�gmD�T0k�m	k�/,{�s���kk�}�����!�aj��������.���p�S�t�қ��/���z��UEW2��r��ŅiE��hȰ���JX���B#�S���}i`zмp�U�r8ag�� 4�PԲ��T�_XpU�����"�Y�	��v�Ҳ�\�!Ȣ���*���o���&J�Ԭ�|��C��V�F7}%\�$7�o��v�9��f�y�xbzM=U��]��m��@�`w������hƖ��$=��	�8��)=�7�� +[�21Ф
6���>���Hڷ�ަ�{�8��jyu�)c��օ7�,����Z'l�{FE�f[�����{�?_�����O�!nn��ת�ރ���m����z�ʹ�	���Mm�i�$�l����m
�Ya�ֲ�6�^M	�T��nc��J��������޳.'�Gm�;�ik�ê� �f�#��Ne^��9^(���DXٛr�=��:��	�B�*�2A�ˋFf��*����P��� n��P�%S�9��������U�Ee�1M�fo�z𣫆!�]���W��"�{Lu	�z(��M�B>�s��q��x:Ns��cd�|�{�6YQ�B�c�v�u�u�ٞ�>�Lt�3"N��l��w�c.��V���rr�]�6�ۑ�vvͬ�e�)��]�r�+3Of;���<�{�ќ����]���<X��Ѿ�!��e��1�i���6F���',l�&N��Z�WX�Fm"�\;Aҷ�G�)N�U�Cy<�M�����[�-F� ���>����m������2�=��q�0�i�޹�M�/�9ܵ�T�����G$L-�Ǔ.��M�e�������;,&�}��4�l]ٰ����+�Y���v��jحK"y��\�Ms�=ɂ��]g%�$�ߣ��g��Esmi؆F'���OB�	��`F��Tl���T�溍œ���d\�W�T�&sD��s+5�ʾ1��ƚ�Wu�DϮ��Vm�w�w��@Ս\T�p@����]���RoWQs�މt�q���t��l��a!�ٳ]��2�ԃB�%��m*��Gm��8^;�ptǚE�R�oeI8���I���p������n�g���^�NE�;RC�q�/s��tjSK&�3=����ڶ�kB#�m�%�˓��聓,[3c��>��tz�8�*3c��A��|%��G��*��|8�U�׫z�pr���j۽��<�.���s��	��1?b �.3@M�CԳ��ǆ:QY{������� ZF.jI��U��?aͽ
�f�GH�M+,ѐ<UJ�81��N��8v�Z��[�2����O~�򼽔p�F� u��߻A�g,�wʺ4֪ڇ�U�"�B��wo����D�7���\�b��r��v���WZ�=�%漼=���i�N\{�"jlE��L�l��{5�&���k�tD��9G����O����.��c<ѪK&kg9��Ax���47廑$��#����!�z���m�ǟ��w���*�����KR����ΣR>y��^�]�i1���������Ic�����4d6�
9�X�e)y�\��l��Y:0�X�K�ǈ2�p���fub)��;�/��ū�+�ѥQ�W�ǆ4�wu��R��� �lGh=�3N_uJt̋
�dD���	ڈ*	;���`�-�����8P����wzQ�5_QD^ J��=�,�QO0/�4s8�qz��y��mK�[<�;\��qQT�-
�Ў����
�$���V�+��R$�����79�l�.��E>@�gWĚ�M������뽹%F�������wP��խ�c��&�rd9���Bx|�Q�U���r��o|��KѹcD�pI��]���+]�W	ue��� b�y|�����j���r��D!���Թ�\Xk|8G�&
_M7C-��ֹ��1a���1��
�{��k��;+Dr� ��YÈ㗜I�9Q��P&��I�v�n��.�v�Mۧ�G�k����Mھ�₍I]���.��՗��'�Z�{n�Z�����X��I����&A�T��,�����+76��' ��#Bڗ����WdP��6hK�;�͔/]������R��b�h����L�Ba��}pܝݢ��W��T��Ƭ툩�1���XY�֍�:� ���4�7�繡�we٥�t{��JÔu���+�<]��J�|�����:4S��L;XRW��d� b�f���%\�u;}�3Bz�t�܁���M��*���5c܀�~'��T/�=U�y<����3%u��	���O*R�[�=�u��5�9��>�ؼ
Zf��ݽ���D3@�C�K�8�k-@2�i�kj֭�H]&ǲ&��~�I{8��M�t��Pv&�;z�ڨ�"��5F��=���b�:VE��7Ø� �k�Nn�x�U��.R��}�ʽ���;�1�L�#��p�.7����Yx�x�M
Vʾ�Ҧ�� D�z�;zN7��Ը�G���h���b�$;���X&ȻS
�Oan���gg;�{���>�e�����ĸ��+3�N�R=���k�Xe3N��t&�A���H�nn�=}���1{AC����w]��L�V��O�]옳%�W�O5z`��}�3@�a��1BSs3�����\�]��輘M}G�9�;G,H��%��uS.jfE���3�U��罸�gfi���}+8��M�3�L+�r�\1,�y�$�ްNꕠ��k����H^l<+�̺�-��\Z�~����u[2ۋߏ��Or2LחTU}�V�HE�W3"�nb�u]�c�S�L�0��9���@\>^4�x���6y:] �B������+�˧�뺘_[6u!V�w��.7��oR��k(����
G1�.���RQ�\�A��ؖnYn����z��ƺ�G��6:��l���m��x��b��ڮ�Kj���.�{��yO�G]�Y�ONi�I�U��Y:%t�X��tۦ��{�XX^���{ܲ+�mo����.�&���v��*t�
�{&��l�'Q�z����z��� ����0�M�o��h��2dk"�:�ݓ���i��T\�=�t	6��V��J�6w~���Ą������:�r�-�ȼn�]B�mZ��⫥��4�G@�a��
��¬����}&�(J��%��ٯ������� ��v�V��j֊�c�tg�b���W\���wJ��X]FsT|&T�P��������r{n9�$��|��c�C'
ɴMsͤ
��8^P��f�A�
T���W�7)cnh���?�փ��������PG�ONi���W �A;X!�*AjX���w�f��}B���]>�������/��R�[�������oЂ]q}���[+4-Q�E�pj�|V��¹�,϶%�l���ʽX�O�h��)8y�k�7zd���%^�@)�.X��hf�8�e�����Y���֡U���7�6��pN�s�]+Ӈ��x��Μ��d��A��"�3���C�W=���6�t�/^�Kqv�1gff��R��!*y�G���Y~ex���{����M�3�]8yq������xC`�m�E1�V�y%�����6]�r�ݓe7@�ۼ[b-�k�U��v���3��Qf��j��Kc�v	��mP
oQ}f���{��}�ӽ�o�d
��4��H�	��f�}{4�
rkFC���y]���XNh�8���M��ĩ*�C�荻b�^�2�����0�ڻ��;G�߮�&���F}����o�1��=��;���KD*�ɷ��
{53QUƯQ�v�Tz�9CA�+i��\�m�f�MSP������6c��d4�5f���t�W��(�7yU.�U�RX�_R�w4���X�v�:���v�t�(*[m`�'�7�Y�s��;���"$�]hyZ���:���=�-��h�]��[w��bS;�ܒY��F͡{�h�+�3�s|�ٗ�np%�S���;;��w�˞ �u>ﮯ����Z�X� ��2�+e��:����z�f�Ι�+��
M�&�9j`���u�8��k�'"�3�AkJ�Ne����7����ỺH�囗��=,`��&0��"j�,v'��ܠsը<�Cur�rs��P`�>r�ʢ1a\�C��p	iFܳ]rΝ��[Z�[�[P���'��2��6�M��
�J�Z��v�U5jb��Y�-�GgE�EL�d�tlfwPRC����!K/�b[�<��Q�Ӹ�"ҡ�pN
][\M̼Q]�uCKX��Cg1H�M�ҷ���J����(�Z*N�YJ<�޷��Y�(cz:�k�8f�]�}$�������:_Ju��/��vM;[4��V��PёP
t�\������.�c��gm��-���o��cF*����﹭z���mwE"�Tw�s6������#�J6ݲn��.�u�=�����.p�g{�u�r�zU�Zx@�,�_g��	��r�+B�}��{�z:�7��x����I�5�3�h���Tݗ�n�)��+�yz�:Z��nWG�0:f�&�D�9��Zt^���]0��#�s[�t�36囂F�R:Wѹ��@�$˲��ĚiV���)榫[���t#��Ti���p���eO��w{G�ڰ,��ċ�y@���$�y�t��Ac+��V:Q���0ۼrӘ8�%��'��s��m�3�x�u���b2r�,��ށ4p�>��3&��Orok��.�-rm
�f}Դg&V�ER�o���.d����J���G	�b$j����K(us���MtM�y�c��p6���g��{ljVh_�r�cs��{��.m�=�1��K�s�C�n��^,|����ڏu2�f�Qt���J�q�.d�H5I$�c%N�&�U��ǝ��OgGњ��1q:�u������(2̌�@bm��|�`4�gC`�LA��K6L�%0�BLH���?�d��qB�.�F$��� ��0rT���6�>���o䰼� �ډȓW$V��pa}�KYn#d��m(lL(�is��(~�����_�Xlʢ����(2�@U��o
����Y�(b���4�B�TP�
AB�L�n�)��m)>P4"%M�%��O[��o?Ъ���G�� "������f�_��c��>X3 �3����}^�~��=���~���Ω��^�[޳�S�_v�N�ھ�s ��;h�'B��y���4�����N}OlTcf�p[J�&��Q�I���=D��Y����1�GhY�>�� ��)d�Ш:]�zG;�!P�3
�3Nfщ�塈�NvOo\t=Z�<. U��z�p�����D�f��B3�]!O��(ނ���/m�kl��YHE��1]}�q�a�ھ͎a���wԗQ�m脢 ےX��%N$vPn�L�oN0����M8�"WKe��R˃z��+7���ݟ �:�B�vZ����>s�F��6P#Cg-T��1��u���ȝs��\<�I��up��y�2'n��7#�Wxd�ǻ���n�O����U�*�\���0W�w���:Z��/�ӛ~�)��g�ξ���ZO���>�n�^��|�1�A�β�̗"Z��m*���@��6u3þ2�B .b���{n�݈N.L����g5�����x ��Jc�M�/���zo�AD�(�:J�?"�m~=��iy� ҥ�XE u�rc�M�����#����M���|jќ\1�l�w�U���'&	V!L�����;X�w�������E{5��0�A[h�2l�v��&�H��/-���W���4r̚���<�鷇��z�Vx��Y��꺯��81����Ç8p��p�Ç8p���8 �8p#�8p��GÇ8p�ÇÅ�`k���s��b`�R�=ޜ�ԧ�s�#X���J�ط٭��� �r��}�b/�c�cu��g��{<[��/���u�=�r�=맑�Q�n�Ft��^+�+��B:�ѽO:�V*���z��e(dy�v��=�Gẍh����4w���)9`D��A�k�2�[q��6�W�{%	���EsE����ޝ[gB�s�}[U�3��®3�9F8��m:ǎQ�2(��4��N9n����L�g(��-n���}y,��R�T�%�]�pѝ�>��:*�w�PpL��D<���~ԸφL؞���me�������(�u��m*�ʤ~O��,���#��#�񨘝4\j�nI켜�=�t����Ӝ�8�;�x��𵻀|��������g'~��=H��s�a74g�ׂ���[WLOrE��$3�f7�76�S�IKw��]��N:Xɺ�kY.��6��"y���W�w�;=�<�9�\���
X0 ���9Ct]���j����
�2���m\�.r�ze�O��E��S���!:��.�@K�D�aMfmu�Vs�ۡ��b�e0w*�q�/�R�u@�;��	��>��n�K��%0�M�Ho�촙�{�_*6v��}b�S���,#<�i�c�58�O�y���&[��wu�٨�����|=�:��(Q�:�hႄ,h�Ç �Ç8p��8`�8p��p�Ç8p�Ç8p��8p�c�+�B�7��W�&�s2���h_���b~&��ɸ�$����]]������I��<��-��~��N!�4�g`Μ���%�Q��s��-p�$�����Z��kk�5��l\PMw�lZGi��TX3��͍m[ϼC����W���m��h�p��7ĩ�6r�d�^[���l���TDov������˶����eQ���� �k%"2	�� ����[�j9��h���g�.���b�7�<�"hT/Hy�b����hCݺǒ^�%�ww�CrEY{���������ED:�c�&�z�a��IG9�h`��]7�6KV�v]b��"zw�C��l�:����}f�ti��_�f�/v�N�YnN>������nZ�8�Kr��6�"ezܫ�3�̎�>��C}����KZ�,����>N�eoF�r�#�������jT�:3�ہʳ.���75L� Cž��w���aC�2��Ȫ����f����{�,Z�$m����[�,0��4)��]t�6{��/��r�f�z�̎�pŽ�v)ձ�V�V�s�A��KC0m�:7������W5	�"��[��$�������|D���%�?)o�"�gp��b�^0�> ��nIU���O_@>쉰��l��x
�����۬�,��ve���.g�dT�fċ��'�Z����TW�rk���lg4'���뇟aݹ��+�ӥR����8p�Ç8p�Ä8p�p��C�8p�c�p�Ç8p��8`埇�l���^�f[�ӗ��<��>������^��Q#���Ph�뜓ܷf:uB�)�-,a�{\[�
�s&�qa��J�K��~Ta�{AF�H�����[��x���K]�%<Tj�t~�4jq��d������3Njk��yNFMԭ�����l7�_o#�J�«T٠�-,��em<�(�PQ���q,��S��>*թ������1����݊�o$r�u�:b֑�[5;�f#�Xwq�N�%���=5�b�4�g,^�ͥ��޶�y�'��GI����kvZ���X
.�}��U����jn��Kym�j[���d�C���O9��	s�=���_�,�+���U��FnwQ�B�Z�j�/�J'���B�z(x�Am��=i�Շ,^ׯ���/��M�z�8���H����g/m�.1���U�f�.�+3��yTÃ��
�i�s�K��J�]Ncl6�lo@T�������~.�|�xz�9��ne^��%�b�2�u=;�ndR��ś�1AS̵����y�3�G�hd��&�6����,hS���퍻�xgzp�I�<u�ӤY���I�@>�:����
QY����n�N�X��	�*�4"弯���	���-��K#+jH]��^����5,��zC�<�\����ֶ���J�(=kx f��'8��N�5�:�O �r�k��'Z�Å4p��p�Ç8p���8p�Å�81Ç0�8p�Ç�Ç8p�*�T���P���<lZ�]���9�kOWw�rޙQ٪׆�KA����	�tN-v3�{5�p�B�ٓ��/vN��fhܑ�hn�NF) L�n��˕׌�OdC��JVe}G���ϻz����h����d�kv�`Jyg{F͘��W�q���%�s��J��GO;��3-���n��|S�y{�����f03 .��M�\�M�"��}��th���n��K�(��ִ6�"_^ֱC�+C/��ȓ8�]�r�z��!u�;1i��}�0)�۝����u.��\2�A��wۻy��������=�Q���v�N�j�c��EVஅ���_NI0�*� ]�#�����7����xUۜv^*�9u]7�êTP&t�;�Ƕ�?Q�:�a���5}��|N�ϥZk{��p�;�tt�_'7>�B�]R���F�	L�!��1#��;|_�����dws���yp	:�K7&5�=�W����曇��y��D���=3�l��He��dɺ{�����='_e�.�]�g�t�Ň��>���8<�;�7Cږ�3�D���zYZ���=J�\x���a+�\v���Θ}電`{#��s���r��*vU���"��L��]���X�����x����w/��u��F�u�� ���pe�OP���py����]��=�s7}ʸ�N
/��D�n��R�u)#xk��9�lc~9.L)�#9_�۔]]�ϳ�򞻲�j�3V!��XO��
-�,[\]�t�+ܢ!��lm4��&��`��\6��-f�n��
�u|�rl��&����r�?:�NA������<�=��w=�Vd�64'vҫE���5y*�m���=���'�ܹ6{/���o���e��þ�/����H2�yN��JVz�a���$m�U�(�Vz�(��
B���GF^��8��}�(����B�\PAg	�(gq�V �]ERŹy������w����������H���ȭ����L����yi�͓D�8���u>�=�;���u� ��щv�G�w�����6��7+�A�z���k2u����R�}�	�}�&�2Y��9�^G�Y9��ĕt1�3�fW�2Vhy�\R��ƹ�R���C��*-n	Ø�X��♪�/�x��wa��}����@�Wz�B�9���M��պ�yR!�!��s��,]�Pb�t��`-��+�c�\J�3lTS"K���3�Y�����˩L #��%Ƚ�n�rn�nm��n�VW)�v�D���YX�Ǹ)qr�c���NW>�Y�;N�PV��8b�ˑ:`\c��O�a֝L�r���1M�2Pǁ���n�vB$��������,�s����{#$n������b�k�4��}LH� �����ŀ�T�Wܝk{�7�X�x+Vv�Z�DR�{c �բ9����*��ӌs��]��u����%��=��n�Dt��備}��-�xFs�ӑ��k��Q݄����'��Mt��쬘��v0��t�l.��r	�w�{Ĕ�@��oE}�~�%��6��<==uz���6�V�Y�k�o���1v��U1+Y��qRv�]�����uf�A8�eg���h>�0�3��t�_(遘���3v ���� �����`�rñP>Bd��N2=����}G��M�>J��lkk���׳��e3���q���Du$�{l�����[2���$�����0�<��
���ڬ#��`�Vt��|�g��N��=�l�L#�a��q�,�q*��5 ��&J�iϔϵ_,�ŇQK�m1�R��X�&���vݠ�Ë 章U\[w�f{k�U{�YP��TS��k�bi9q���qq]�76+I��o/�Ý3��L�#yJq��;Z:f�shQ#NPB/v.�w�^��N�H��t�1�i�9�Wz�zQY·�i���]d�s��l�υ6��3i{}��9䳣��Y<�n��.�L�P]8�q�<Zݩ_�)�����r:�_:�5�;�:i���C�CM��W;n��m��� 1��uEnK1��㮻���ž��&ݧ�Aᦖ��5y�c�kk� ���P�N��h[�/����:j��3�ef�Ć���7��Dm���u�w ��c�ݖ��Ӡ��0&�#~�ŽW��NTIVP��ۀS�Vp�K&�"'<o�K��c��I��ww�^0̥��p�`�<�ꦽ2'�5o����U��zI��I,��}��Rǹ��(��X|@����b����㠉��rvTH�;pS���젭�*�����d�@�oE!�H����u������ ����;Ǡ9_f.�Ϣ��,���n*f+8(f��n�U І�Ľ�^񭚞Ǽ��J{�����\tE,R�s2��b��o���hg��F��S}�dJM��R6���嵜�f�>5nD>o�3;WwQ���b�7�]�}u���ˣ ��h��ܾ�_�#�S���0MpQ�C�U<ͺ��Scu9j$J�P^�Z�����c~��>������JjK�~^�=��x�M�$N%;��q�j=�zn�(]���wH��^٭!�A{��[4.x� ��x��;�1��vt�f����@g�d޽��W]]wb/=�&�q�3�� ��8˶�S����.Zl}���A�� �)jvl��4�W'g<�2L��;�L�]��(�Wnz8�j���g��vq�������e��<+c��c}<��ң�����f������_5g{�pA{�Sv��x,�z����]���ޤ4����`s�˛�r����p����ފa�jx��G��>(+9'L~ס�;�ۄv�{��mɪ�xY��>��=�N�u��:3���'�[��u�^��!Aӽ�2�s�i��K�ڀ���t*.D2��m��������S�;�ywf ��]�r2��#*����/���R�P}���hW���:�^T�������z�����S��'V�۩��K��;Nl��жح��S�S6�OWE�x�}||B�m�͠��6�}b�Z'l�]���غ�J����Q:RM�{r��5 ��8ݞ�k����p��h^������k`�nmՎG��d��v��6�+�)���/-����÷\3w0b�\Eތ)�U};z���=��
'Κp��$5�"�.Fʬټ;�l�fR��=�n)�e��pS �vr������2�^���f�P�G��9��\b[�������F@DH��f!aю��w�j��F63r�/j�/_�3-���Ο!6x���G���y$3"z���
s}PZ��F����#�29M<��	�s-�e\�[����Xg�G��wW-���.�6��Mfd�{����Y�!�%��������^dHL��M����wlm����+-P����+R��	d=[c���vή��yXq�����{!�J�����$��k�g{D9V{()M�8�8���]��m�٠�f�pn�^��+���'�6R�K=�I>~'��P�f����8��ް�f������˱��{/S�����S��ƺ1,�xT�1�&�Y��]��=E�AVd�f�kze�4�ط{��V�ϔyJ�Mn�1⥈���s/˳�ʾ|�콗B]��*D�Q���%!1%�Lyi���8�".f�%����qgp�E��m^!��|�"uI����WA�i�vz^gl�m��6Jv&Ù;i�去Wv�Wa���鹼0�)�m�s���f&�o�JS�k�ޘV���-��j9��kf��{���S�<S;�h��%_�:�!#^珔��/1��ML��}0(U�d��B��k�qX7Q�Y�S�,��\=��l�Pb�MD���R��ܰ���Uo��bzg��N��x96����`���&��T���NQYM��n0��eZ��nk�}�AS{�Y��nA oݢ��oca!K��໸�{�e�h^��;stzԜ2�����i5�>t�郂���]���Z���;w9����>۪���~�b��q�5�iNq������^�#��%��Q�����Y}��tJ�������;w��xEx�Ta�ݞi�$��I��T�M2_,�����g����0fo����g�}����+�����__��(~?�S�����rYg�j-�Qg%}��G�ٱ<�<;��L|=��p&f�şT��e��2�< �}w���/d����}餻ܰ^�ڱVe��Qi��Ds}b����9�{�ʴ�z{�T��-C�Z}�uJ�IEu͵Ծ�8��}���9l*Fv��]����hG2��{�v�	{\w�f�^��sOE������"j^NP E[��`�mL��]�.���ǝ��н�8��Nɕ�ҙW�8�O{R��c*���s7x�����V�;��35�b���u�f����J��Ǯ���]͐s���Dݖ�VKǋ �q
lU��jJ���{]�e>�uԱw8�Wq��"��΍�5���ۏ�;x�\�v_ \��fz�9�*�������n��x��S�-� j�v�G���dЊ��I�L׳i�T�n^�Ͱ�o�A��K�wg�����b�tQh�5R.�f�b����8#�o��O��`v�>GA��[ޖ�6�vO!��cn�PW�sX�vm���G�?d�g�D'���ݾ��������0����e��h�v!��k���-�U�Sm0��=	����V�ض�u	}-�(|�+�Z����듹۫�gi��6����t�Ҍ�F�����z[;���x=>7����5QZQ�ӮPs{�V̫�(`�_��Hm�Ѵ�MD؄�n��(79��� �PQQQ��D�U5�1��5�j�����UTi�D���>�:�M]ڊli��-�ص���&�UQAU1Z1Dьj��*�1,�i�N�:u�I��b�*��1("-����AM�QE�h�V4[gmTQ8�1UӧN�;�ƋM�#lڜi �h�)����`��b�`�*(�&$��N�:t��1U���(
�Mh���*�F*�a����cQDƵ��+5h�PUMV�
b	�F��6tV��Qr5���M)DA�AkUPkEm���H��(�"ŧC�(KcDPɣQQIRCZ43ENƢ��*��$������`�)M:���(�)h�:�*&��"�m5m���b�q�b"��"Cm&�TD�EQE�h��b
i����E1,�I0�'¤\׮'�œ�\��:��iT�q�P��,�LGs;A$f5OilV�{$59mm�f�C�t���n��iЗ��&�� M�Q��t2��ew��$G�ҡ��fӑ�OMn;�l}4v�8雬��~�r��(%������/oر��֒d}&��ʡ�yq.�r+zj�5�<.�䞉�2+uȻ�q[_����~;�ę8�k<E��T�tH�n꒸���W@�E~u�%yֺ���@݂M�x$ˇ��Vj�K��bI��F�CV���?$2�u���"�����L�<�q�����^�/ާ��+R�N��+���n���x��=	��>äNfM�%�E� WQ������C�g�L]y ��-����oǅc�q~���j(�d�þoٞoi�s3n�K�ko�78�c�SnLY���p+�"��i��7���2?=��sh��M4��<�h��5��v=ԑ����X��z���\P�}*g���OÞ�-�?u��տ{/UQ���^�/e����F�f��-�'���+�9�om��r��H���mJ�Y0֗v�0ތ)ԫ3 `�	ۋ����v���莌�������!���2sy��/�Y�}�����t��*�A����J#���mXUd�������~��s*�[�aW��ө�)R�}���H4�#��%��y\E̊�sڹ�
�_0���%��^�ݴ,s�^���[���g��w`$Q�Dx�<v
ʤg�ǅ\^��h��<�=�<SΨ،1u�l��̲o�A6D�O3h�^]�P-:f^���׮�k/}K}�%X΀�rj&f���@a� ɻ��ƑyG��{6i��<�s�Y�����	j}h�Ɉ��r��3G��\!���	L��%��iY�[WJ[[Ո7"	[�'�ge����x�.��[�l���x2[G��ͯ�߃�/o�(���φB����p�)u{תW��n��}���"�kO��α���$��� �/A�׼3ժ3n�����zW�Q�c�A��%���'���L�������~�o�)���{�j��Y�;7-7�=[�e�݊c\�m�;4�th�W�{m�+���0<ݷ�)�8u�v�gY��e8<sV�������##����� n��wF�\s�iR��v�ׅ�t磺�P�2��G�2x���v%Ƣ�c�*��V��7Ms��N��O���AP��ϑ�������bI��y��t����y���{�5����<=������:׶jRm���ˡ�c�Je�x+�e�j�۵Q���W�D���7�J�.S�x�"�V�,_[�*�9�)z<��S}�c�S��=:V�2O|�Iǈ@�[Ll^�B�������VEmw[p ͎��	��I^�z������ڷv��LJu����B��W����P>'���[�1&:��̧%�U���Y/�c�Uxױ��G��0��+���ޭ��uݲ���^�z����u�Nnй�[�O�j\�P�~��⍎���z�^��:^���{��w�-����_˷��2�������z���W�lX����u�v¼����69���Q3�^%��_�|_������l�+w9\�B��$��=\ui{&N;����վs{'D��]��&�]Q��R���@z�~�骙�^yB���g�����>��'���C^����x�M���QG�tœ��T`]i� �ܔ���A6� 'q����_�j(G_�Dh���w�/�&+��V��OVd�Hi�ÈzK���Z6i�j�� p����#��^/��������U��V2 W�ti'��z�z��q�NpXz��]=�#���]�_?|iV����{]JO��Ͻ�~����S��Ncs�M+�g73����@kw6,�NAݎ��Y|rL׷��sS�m��6�ph�>5���;!��� ������l���w������p7L����&z؈x�e$�q�x�v6��yA���s��|��o}��D��N��CN�Lu��=�*���3�W��f�i��ʺ�O���i�q8ϬKm�ތrt�m{�N��'��hl���y��3���\�ʦ��sw�|AXY9�oN��'��Z�x��i�G�+����s��uZ"�H���ę��y�r�P\-�,m��8=W����9ԋ���Ugm�4�5��bwp��]�%{��Vy��;U�I�a�)�XSѤ�6��YY�˥'@����)���m#�W^b�k�oD��Z�ۣ��k�>7jj��iQ���OP5���7vd�&�6��
e��J<�Zw{`d�ߛ��t2d��V�[�l�E�9�Z�>�/	��h��G��exsx/�����ۣE�p}1��!�5����_�tƂ:�a���"N���>��: ��{�XP�����#[c�K��y�{ܻ��笎�np��3�Ng�lP�ʃkލ��a,{oz��{<��N/��9�{��^��q��]Gi�}�Gr,��-Eo|{�1�� �.�>����TT�&�#e���I�}&��ʮ�ʽ��;��r��u�`/@��{��M�׻쩒�`����:4�w�	�<Y��x#^������ӆ�{r�@*���$\����V�}{�I�Be�0�"�ɫ�4�\��v��d�#'m��φy3�-�782,��[��Fu1�u��H�=�1o����Vϻ���C�E�\�w����E�N��`wq5���÷Xe��9Ƚ�A^ŷ<Ǜ0��Me�QW\�,*ӔF��ؒޠ��}%��٦�_w�f�Q��sn����y�j���G��q8��2�uu
��3� ¥���0^'R�I���MMvX�*�i�ba՛��;^�Ii�Pa�Cճ|�����]�eӮ�ڻ4��]�u��se���|�3LӪ��ݩ<j��~�>l�����O�F[�67aM�Ǫ�Ԡ����BB�94+��syݧk�uEzN�g-����s������{H��_]Jv=NeP���ڙ��M�Sۥ����7��;ޯS����Ѩ���F�K�����יJ��o-��&{���ԏ�Q��1����;�L�g�A�b�Z<8s�·�D�n�lj�U�F_�ܳ�2��K�����J����{�1�)�Qlχ$��q.w�i��OtyAZZ���o+�P�o�{�xP��VVA��G
��j��&�-�b,��绞��٬����� ��q�5�EӘ��oZD�
���%�)l���hX�0��^�{FF�����=^<������+7�Q6�����kR�4lo֥dC6��%tw��P�/���������]8�s�Bb�W^}Vl���q$m��{;q��ֽ
fp����>"��n��M��>�X;$Ӯ�۲�q���Z�.�b���/��5��z]^q�ڏ9�<�"����4�}V�Ո7"	[�$w����V��G��u+�(�O{��~3ƛf�m1�j:��1��4�%걪f��o7�U��OKtq69���;&I�U��{-t�F�8P�Ά�m�<t��d����n^�s���_2q�x��?��5'C}kwbu��}�����Ad�X~���xnڞ��&:����8o�{��>���=����H���І�U]t��D�hy��ϫ�G���3|�G�p/E�y���q���s]���3a��z{������E�PY+���ށ�>�q�g=G��r��Kn�R����Js/CL�\d�b�	���^�C^x�O;�,�5��{Y1����U��(jĳ_ez�-�|�̈j�Gw�^ �-����{	��Mŋ5=���[�j��_��<f���q���n���`˞�2.뇣V}�DBrC��oH��)pxLE֩� �>:ELU>�-��k`�)�F��-&:�0*� �8��(���}=ݷ�����C�(����辧B��UX��t�)lwV'nT�l���ŘU�}�q\wҿz���鵉zo��ʋ�2E˙���g���8�v{��n'�B/��R�`��k<�u|خ�
rQ���[�ȭ6	�%Ô7׽?k��9����5y��F�uL��p��M��/��đ2j���r.��^����B;|;�u��2.��KP�N�ܚ�͒k�_���m9��{�2����A�pf�N�
����Y(��t\��=�E�|�gc���%�[��g�{�H7�	�uz��H=�pl�J�r�c������.z� C�Ɏ�X��ti'y��>��留�	N� ��L���xü.��<p/������$��<Fǩ���QJI��=+Ґ>�{+��Ud���>�az��rL�0O#s�z�q�s*�}��9 ��yu���(�
l�3�P��[�庬�5I��M������l@�7&X6/y��73d��O��{�Q�;eo<���������^�p4�n��!�#�ʚFÛ�v��;���T��岵[��3"�����4vGi��p�'B7�����2�>]�"������[�tV��P��e��h��!�[��Fn�=�{ֱ�R�o��g��}}�-��8-v�0щY��j��mO0�����qT硭�~�>^ܥ�=���I�F�^�~6kOj��&yGHxRP����}�MWUL�=��7sއ�i���Ǭ�GΗC�W���-{�z��f�Y���5�3�7���c���;�V�LOiOa�.��X�*z���yх7�	MȨ�,.Ÿ����^x�����^��S��촨�o��=S1WL�g�����鷔��ǽ���l�9�i"{�9$�y�t�ڢ���m]��\�p�O�:�Y��GS��T5�w��J�G��f�WT[��R��>6�W4���5�TTEG��I�� ���{Zsj)��ye��ܹ��5�ﯣ'�%���=������m�n�� �I�gr�L�Wq\��j��DI�3���gn�����r;��3�_��.��4��NL{�R qY댫�����xm��<xz+��+�LI�p���1�����S�ќ�%�`�O �������]0H�F+7fe�����f�9�`�R��ܻn�_V8\�o�ӣاQ���),��6�ι�97w��Mh��解,�Ǣ6"	�ڧ���e��*��p�a���+�d��lrdm�c�.;0��i7�&|O���Ng1�p��'h���&��ڶ����U�D�i/s�L%�L���� ���r��"w��fkח��~�����Qi�U�;��+��@{�������x1EVUJ~L*��)Q�]�y����ݓ���g�n��οd�kl{����z	���IcD��7�����\�#�7;,5���?=��p��:�޲�eޭ���x��ۓ�ln�bV����qN=R޸���Az:g0:���O7'��O�y�5=���X�����'�Ր{jy�J��^1��kR��6O,��n���	�A��8#����G���7�vUٰ�_^P�A�m7�I�_�
�a�V�N�q��u��y=��1�j�)���U9���7�s\�:���0��S<��;�ģPes
�8}a;��4��.��l���xŕm�5�g�X�)n��';�<���{�p����&�Q*�``B7E^lI1i��'4�yui��.BF�O�Km�|Z7/_]\^��~۩Ol{|Z��kAF�~~~Ə����,-�\[�:�#�l	��ϱ�]� +��Um^ME����t�(���M��5Bb�z�����i��G@�%��i����T��1�v�rM�Ke�\�����U��Ŭ��5�:9&��7uU��L�ճ���rZ���;.غn��w��P�l�ί��XEEFgc	֗�����p�J�yh����9r������z�A��<�j�r�'�%�K���Ǿ��J��ܮ3]��G�U,�
��X�z EIqq�`�<�WОӬ�Mx�K�.�h�-�i���ky��D&�k�Z�:�嶶����m�B�}�77��3�+$
�|H��-VN�ia�wT�g�I.{����]�bٶ�pnSyH6��`&r�z���Q�����vΗ+�*�/r&�x يՋWC��P�1m�Z��;�JJ�^pe^�{3zwon���JГwA:j�}M�b;'J!��w�ֻI�`���p��ano�x �>�͞�W}䤰��;�٘�ۨ��k��4�u�!��\���T�,��,��'v:4�k\U�p,͝���.g�:�X]�N=.�Y��K�
T���Uy�=%y���=�o��.^g8�h��!.������&n���sN;���s�L�Z�oR��= �<��M�4��M�<�{�ml�^�*_��"��6����k�|ڹO�o�m6�_^��	�h�	����Kr���a�6+��2�%Ǵ�5W25��[�̭���>�w�����f[�o�k�+����=;��8��Ҩ�«_%��oE�ޔ�*���ՠ��עۻ�Jn���vm]i1m��JS݁��Hl��=�f�2e=�Ė�eA@�Dm���g)A��ge���G��-Y5ktgr�]�+�8���/.uv���Q����[/d3,��}6��>�M�7�U49����󣛰l��H&I�W�x���xp�Z���f��wvF\���5#�ؾ��gu��������!-5�u�ە
��-#�t]�̭���@r���%ůW;�xv^�8����g�'Qm�e���Lb���Ggi����WHv�4��BsA����!��PZ;����U���~}�%+��\���"dww�g�b�$buwtr	�}��Qu��)�G01����+	|t�=c�;�h����Q`��[;L֮;���w�CBgT�׿� �[ܴw;�"G�D�Yt����P�h�b�.r���X���,�U^R��J&xCk �X	$�A����b�&���֦*�=N(/-Tk�4�Ǉ����A؂i�3TS�C��/��M��� Ũ�����{N�A��61�#m����4PV�h"0^^Ll^LQPG�N:t�;���3��*`�j�i�#g��
�O����4�S`�+cf5jǇO�:��&�ADN+Q`-&�kY0i�I)*�bj�Zñ�<�kͨ���Q��j,&4�kXlMh5X�E&�a�������bb
��45�-�b�����*��m�*�.�TT�#Z����cSl����;N��M>S&!���AXlE4s��y�����5A�3N,I�0�2U�Eh�Qͪ��#�|���I3Fjb9�IM%>o<j*


Ѫmkc�ʒ$�J�	��&b�;\Ψ
|�kE�ꩢ�������o���m���a�)r� �q�H�&ݻ��ɥ���C@W���|�o�=͸�m�ѳ�qس��Ue}�M3������ӱ��&���c����MCI}�6"���%�)�ʥL0�^d.@�S-�!�lS�=c��l�okp�i�(��
W!Q��ȼ���ֈGt��?>q�n���	PS�1���?�Ҷ�L4b������r��A�ȶ�-��i2\-�E�iOԅ�r�)�}��%/j����%����E&��M��ȗ�Ȇ�����tu�fsc�,]5�bON0�ј�oV�^��;ǐPH"X,�	�|��g��3�d
�n�|��9G�y�!�	C$���e�j�����l�����0�>SȜ�)�i������SߛY�BrO=��9w���2H�Ə>�Ɩ;k��d��Ϫ_����y�w��`��Yz7%�L����,�%���=�J�z�3i��2)Q�����.O;q�.,5\�Q�n�4���ϟX 0�>��\0�r��gU����o��K����2�	}�k`�N�M`���*.�^�g
ؒd���s�dtb�b��B$�����ڜ�`2��[�;�?����IObL���F�@S��X�g���(bѳ)!7 �66�Ŷ��zt��G4`�vw󥢭�*0=b���ҥ':K��7�`gzi���(�E�f��OP�I^�yXղ� �}K_��3D���ɸ�'6�x��ѓ��;��<цus�)����^(����d�'�o�2D��ف'Xܑg�Iw>�Vw/B{������.>��I��cd߂�1���/��>yF�/�z�^��4k�{YDbh{Yʅ��a�^5���9B5�꺂�C�9��"�vx�M
�Wu=J�ك^���=��=zL9}�g:��N�3L��;$o<��W��C���[�sK�:�u���6H���nvF�`��k�G��P�&h�Wv,E��3��,ո3��|��{�g��R����k A�6� ���������!w^�^k�#��VE�
�WG*�b�o����iDß��7�\����T1P|{�d^�}]~͊�~/t/�Oӱ�ܷ:[vxG#���������E��׳f�c�gO������ȇ�z`��r^��..���gH��C�QVԌ��렜��%�����v?��*.��ft�m�C��7b�4\����Ų[�S]�Ʒ1���s��c���X�hR�*�
j򸶝�t��Ȱ��V��k�N7�����B1r�d
9]|��ӹ���V����n���L����p��\�`�p�8�.����s-<�0�&����X1P�r��:�:|����c�R]=�,�ޅ!%)�������[�vD����L���>��~!��L���	�뚶w��Z$*-���MH��F\�z4ᕏ�'��N�ZFE�UE8���3�2ؕ"�㓊�R]t��}����x�3������_K1=�a�ǩRe�/�r�^sa.�S����m��3.<���˥����+�=��Ȇ�n�8?�:�G��Az;YQ�P�+)6�ԕ1�.���8l��K�ͷ'X�7�b摵�zk��XV(*/�� :�s�c�&��,.��݋_kwxEfY�K	K%s�UmGr�ѧg����%�<켡�p@��'6m)1��E���?hAr�b�X�Χb�Қ�GLI�~⨰-t�)�'�ȁʤ+8eB� ��;"rp�)�	D����C������r}�#X����8�/ҹ���'E�yu�,%�q���;�퐮�R�ƀ�*��*�%h���l����^N��Xe�H�8��yΌ_�W���`��Y���c��o��gʼ��Ac��OC����\E��fI��K7Iܢ��,�{���:�^�9�NuB<d#��v!�6����W���yZy~�O����`����>�o�{Vn�6¶�W"`�k��Vճ����wrA��ɕ�W:Z�ܝ�R��/^{5�;�;˪�E�����ޗ�t8��[�V;'l�j&��٭;z>\ToU6��ߤ*e��oUwӠ~>0���s~��l㽋�۔ 3���$5�fZ���V3$v�U�8��dcl=�ǊN�m�Mx`0%����r�\�Z.��VEgNnuF̟V���=2�"{^��$q�/�,a  ��܍�MC�.s�<������=sd	� ,>�b�i=�F5+ʩkj�2>A�Yt+����Ű�q��~G��*�>K2���5�k>���q�j�`:�Ǻ<{�.`ᕚ#�q��Ȭ4);i�|#iҟ)�3�p�|"�t�n���[c;`AG���Ġ�S!7���#�O5t!>L�rgyU�0͜G��fzs�Os.עc�s ��q�^R-_���I�Jî� Í��@"/V�Sz~���nTk�^�m5p���tby=#�g��V���~^՗h�O��9�r��F��%軛�]s�4���ַZD�(��dRt��T���<���cJ9:�+L�@�x 8y(z�e���7n�@�W��UvLşC�b� 'j@�rT:VfvY�O�a(,it�\~!���U�����_ί��O�S�v�p|6e�=�{x��6b�� m�ȲT�˛Q��l+���VS=���7����[� |��+|7R�^�^M���g\�"*ū|jP�d���4Y�w���Y�q#�]��o<��#��>7Y
��ɚ#�m��Vf3�06��a@���փ}�}���1Y��jH)`88�J�}s�Hf�KUu��bnV�gz�>��֭�XA�|F�&���1&�"4��n��"wr;�]�ӵӉD��0�5h�,F�%�WO���n@�j!ddACh|����e�hmW8z�?�m���������(��RސPדo|cя�#X���1� ��`5�(`�	����E�{S��|�YbZ����SC�dnG$��/�
Fiq�9�,#l<�9!#�lxI��Z2�5�����Z22�?,{��Ԇ��(�%=�F0�'	��wk(zFI v칆�b�Z!BM�w��Z�
�\��H���C��@��᭹>OE�����+u���4�d���
�%�:��[C��(v�>쾜�r��3��N���	�dde9������[`\�3u��y�b�9���:֌�}�L%����b�Q�O��R(�ڡ�Ӵ`����6��*�#5ѕ����A�kb�3��P�f�ܮ�aG�1�[ռ�o��'xzX,�L������/5)�,l�k���+sPЄ%I���P��=���+���T�^8d�^iT�C�E�R��9�1�~8R��`rn_t�U�.W9��"�2ۉ������ۖ�<>����ۗVV�0%�9\N�V3�P�Q��.7��z4�U�y����Dd���Q���RŸv3F��fD�pܫ�5Y	�� u�7&r'�Yh ��{^��NI�vjM1�����<��S��D�:��)��XO��1��>�í喺9�;wN�.�7zC^qN�,�b�n��<�`���`W��Be�]�9K��)R�����ۣ���n`�"�B�n*vW ��	�$47Bvx7Vt�Q{T�I�M���-?$�:�/�Z�&�0oB!�P�Q��4�=�.�xG�#��5��-L��U��{����Җ纳o���G�zK�~�g�z����|�����	��i�C<�,�tyf������Zt�ͪ=|CƠZ�2��İ��1lF<�R�*n�Ǯ�'uk�v� �O��>û��o���S;���ζ�����Z�b���d�����ӎ�xѯ8ZF���Ht�#��4]c��k"fCR=�K�Z�C�B[קa��ʄu��@8y�`��4��
�-^O��4�3��ҡ��%�w��k�BA�+����9��x~��i��wH���u&$�q�osw,qn���]�֟G	�.�V��z�o�@����X|�ܻa�rW�2ǽ[$�~څ~������}T�w�˟RO\`�~V�sK�L�h�ڞ$�7�ܫU��[�("�uf�_v+�K�<9H�*g[�/~p�f�b���>w���C�֪!���L��n��	0�&��S,V��kkV�&���Qn��ƍ�qn��������떫یQ@�Io��ќ��|gj�7��A�݄b���8�������\Dp*Av�D�4��/��[v\s��w��X�ڠ�qG!,U���z�l��l�sK�X02FI�n�8��V�Vd�WgsW*��gdv��m��'����,q�%5��dA^����Wj��� �m���c����)�P��v����j���?B�=��Ru�Ȕ@�E�5���gY�i���+���w������
l~�qA����r>��pFz8�A���*,M'X��lC9�{	��6�qڝ��Æ?�B�: }��P0�b��\�Y},�7a�l �*L�2���躌�8�E2�]̇���e"���͗f�xa~є$JD�Ð��`_|��'��N�:�lh�My���ء��Q��y���!Şg�2$]ȬD��^E�!֚ւي+b��FxE�s�e�7\:U��WB��;E�W��\�O{Oܢ��i��r rt�q�v^D8W�M�J0��X9��3F�v��P�@���+D�}E�X�{u��E�Z��Sb�l��B�8� O���^��MJ�m0�/M��Y,̈6s���}B�,�V�گ�3����%#��0n���ގ�ȃسx�D�]��~�/M��8=\,Nm~K�;{j�cաym׼�gp�ַ;V����F�[j�%y:x!�e�}{U5� �ܳ�����M�]WD�r7���`�ŧ��ʇT�m��hZO�w ^es�PK�X����)5}���Q2�����;P^��T�@���J���o�`��di��@�	�u\>�^��@Y���5t_p�oȳ�7z`��Bu[j�V�����	ł�A;�,�O��ܻ�v	�|�"�9넶��ހ��0��'�K�I���+m؆Gl);�IZ���I�q�y�r��M�+�d���X��u^�*nz[-xi�Pw���lC�*>�e�}����r�>�`���E/�9�޼�)�oY�
9�zN��E����ak�A��l�/@��5��t�:b�7m��&N�:���os��r܊�������/��F�Kcz��!s�A�ʑ'J���mŧ�"�Ŋ�����԰�
��C�{�������i�9�>"u�8�xmn���,q���^�Nj��~�u�o�t�Wm�隨b�,�)YE�[Jq$>T�HM�x��Q��sz��<n��֝�*g��е�y<N��T�	�o@�O4���?))x�`�Tλ��0OIU\*��w���lj�s�e��'AK��$u�C� ��t��
��U��wy��?�Hc{r�7��T��V���W�P�@ �%u�|98�&ծL�vy��q��7�=<�	V;j�+I�fcN� �k�7�[yy�^��8�Ub���߀����.�A���fJtY��sǩ�Fx�eoX���~Sj�D���f���C�l��nV���fT0�t2�Cy-ht�#�):a�aK��L�S�P9j�6���]]m��*�[.���[�s!!2�	�	��Nʇ޲����ŧ�RRX��n��m���1y�ef��.�p� �mc�̇��rb�yu056��;B�	��Q��oofș���p�;��W�_���+a>�}�l1���d�ě�ɝ-G��<DXɇ���'�n��L�3v��K���{����'k���t?pC�^�����;������L����E]��j]k���i�*�K��h�9�C�-�N�נQ����\XxA�W=!�]o;G�Vdv�nc�#t~��py����?���3ڝ�B�+Ln�5���t�mGg�]�T�`�צ
�W�'n�m���@�ɲ�'c5��h27k(z�A�!Z�v�^����]��Ļ�=�L��[�O8��fh��T{��Ǭ{8;�sO�p�4Wd�+����{P�]{�j8I5:��t�3������U��|�-E�;��6�ì�Qs*�R�>�'�ޑ0Q��т����,��Yz̾Qӵ$��	֪*'�w�PﲟESa-.��/k�F�K5�1U��:�\F��3h���Y�^%(	�9��u�KE~���	?
�D�����Zf�Ň��ã��p��#[���'/2W�1x�Uܺ���5͆��g�N�z͛O^ǚO���(�P]������x�ꂽ�35҉ʍ����|�|�<�`��ɪњObWN0�z3���տ��P2pD�Yg#�:d����˾�ը9��B�ήjЂqC�K$�3M�`J4��ņ�++�+Ƶׯ����l����C.�e����"��.�FMdGc�O=�����Ju`.�L��Mm~������Q�|�0�V�-s��.��G�<�M��Mx\���GCo��̞��<EHPT�H�l׸q�	L�bxD{M�>�#L�j��y�\�C����C����W5C׾���,�B8��R�7���u�4�
���e!'\^r3L"7 ,��kr�A֌@C=��M�Q'8&H��
�ewY����Xֶ<H�#��;ϹW�?yċ��X��� 8��.���e���T�����g�DbR)����� ���4�iO�ƦI��H��A�l�� }��vD;�����u�|� ?U��<}lvd�N�ﰖ��"
A^�ZJ��8u�A���n[�Y�3>��g�h��!�R�S�ϛ:eaYl,�T����J���.���s�DC��.�d=�}���9"E����w�����ko�	,[7q��Bnw�)��RKYt�ɤ�H0ͻ���z�5*}�ז���8�%�
��� o�Nm��c{euGC�vK}'I�o>psT�5w�sX�;��{��⼻[�RQ�U����j���P)gw?z�|�:�)��������z�ZV��^��"��,Lx��$�ԛj�YԶ�����9T:�#�KrHt\B�խ�v�ї�����n�<w�?6@N{�>�iq�� ��J��{�m�[��ESEɺ�W@�K�
���m�U��������}Σǰ���[�<ѡ,f�b�<₁n;�	�^Ѳg1#L�s�\�v��j��"�[]{��d�V;Py��k��h+��<y�莌�������V�u���n�+�Mw81�`�۩uSC�U��ñ��Mg`�oA\�뜕�Jg�ڝ�vY��@�8=�|&��ʻ#��@歇�昚S�gw�|�{j�f�5�;�	�|v�]#W70��V�$��p�h*���0��|�F���|�:��wk��Q�$z=�=T�W����(����oC�̂gFk+j����nN:8Щ-:�A`Ҿ`�D����bS�Yx�w7(���{����Sb�yw'g︯_fγǅJֽ�e��K�6ۍ�"s�}W{����Vi�vV&� ��:<�Xv6�5�t��%
�s��R�E�9E�YVv����/kҚ��g����h9{I͹�|.�ʺ��1��h];!�{�9�f�a�r���-��OE��q��4i�@�LE-ƅl�XB�k��7���YË�K�|&�A{W)1�D��u�[�̩���d��1�vX&��Gr%Y0����v�=�P̧EϴC�c'J�k�]2d��gp_Ǘ�����y�r®굪/'�;�y�z�V���p��q?�x�
�^�Ή�W.��&��K|m�v�3U�N�\5N+B6���+�v��=if��`�EզyZ��]�@3
�`c@2�εj�{m�K�Î�n.���s_*9��eM۲�;!L���-��w�xY[!��q&�sT���I�4r�2ћ;_�Ό���o��L��D\�#���57Q���Vq-���� �w����=5}�EJ���[Ԕ��fp�876��U��#���CQad��5�����Җ<S9�7���\w���v��{�d���X�|�U�l��3O� ��nX|�]G�ݩL�4�un����N�2��G.z��p�����hG��[���>�b�t�]pZ�[X�9ۓf��ʄ���]wH[��8L�L���;Χx���V6|�T*׽Dغ- Z�q�-��zI
L&X$�d(�a�9DPņ��wLHأ?3���{Q5T�IWl3T�Ļ`���C�ITRUF>c��t:CDy�y��W����Ɣ֋l�풊��8�͞N� �Lp���ӯZ���#ՠ��I���4������j��h���<8t�t�٪����m�
b���ICL5R7�Zj�
1���ӣڊS���V�()��� �1<�Jb(�K�*�y��(
ii�-�AB�ER��C���J��O���P��P��T8�TPE�鈈��< �E5EU:��0�CD�D-h�T�UAˤ���F��h)
"cJU6�j�"j$�A�t�%�F������+��SK^ZP���]6�S*QLV�����ŋ���0S���[�h��W!2Nk��P���V,v�j��Ĭ��-����yl���m�����J:�W�����o��![��.Ba��P���I<&�Ʋ���Ao�,�j�	�d�G=��.��+������?����|s�	�|��q�Gi'1�`�������
w��*�lm���^�\�,=J�A���`XQ�ե:�[m�u6d��o��v'Q�g�-��w�J�vb6���a<����������BN�r��>�w��m�9�>S8�S*�]�[�\�����_���g�<x�tm�Y�X(������`����ca{QqwTK�3C=^��Z�#6׷PF+��
:X��gY�ٳl� [:y��`���_���6�Saܳ�c������]�mC�O�k;'�,�,�.�g/���2���V�v��3)+z�i��wL�O4	q�k��Cƣ����b8�2��9EpP��P��TXS,�U�l;������ew���䙻~��S������Bn��d���><O$�?��N�g�����a���1p��#i�O�UȢ���/ӑe�h^4� �h=8��7Z�a����#^�2��/���u��dkޕ�喗��,�wyv΋&S�	�́����o��_I*�c��/�L�D6��s
���o�v\�|���u��=n��E{�,+��\����n	���җa��MV�+�h_wyt|�1e�8o~��r���y�E�mA<d�7H��q�O����"h��|��u~��ȧfw�hMR�u�y�/$�j�fx�IJk6(����}�\]�ȜR±h� �k���"�ŦJ�g��N��R��n����V]
7㴘Q�\��=f�'�IcH�C		�ݚ;!��i���N>���xk��Tu8qg�>(���5"���m�|T�Z��St�|�S�֭+u����2�r���R�O�_~�ppD��`鹤@0�׺�soi�K�J�[�k�����wx�ξ�T&�س>�%�O!���qPKc\�;��p��d\�=�3��棩P�mC�0���EdA�U�/�\,��\;]�Θ8gq�j���[��1��'�C����]c*����ks�A�GK^���f�h�a@%]������F{C���,�)�$�bMߊM۵0�^AVi���Ӕ��lܖ+=�L�dZ����� ��˴��,�C���^�`����Jb��@��C˯�:P��kq�7H��)�/���pE�̤��/�+$!H���t�<~~�n}�� ;��[>�~Z��X��#�v�i���R;�(�U�T�9���씐:�bO�lg��ԛ�gPT)y�����t�V�7]x8]�@�4m�|�5�gyY��|���oOD{�����Nx��LU�!8W+�U����tu�<M��uR�iT�U����g�잶���*kiB��`��
��,�T��^UCer���a"Pg��B�[	�tm��O�;$�;e����D���
��8�D,G����0p�,�|�3s�d=�<3�ĥ���;�]g�F�7)�]�]�QE�s���ml�A��w�O�r�y�����.d���g��|8�`����]�M�־���1��Н ���9�5C�J���u�I{�����|��tt@�{�!'\ĲN�x��ݳ��ޱR���Փ�z\q²�3�%�{�b�5�k�51��"U���S��й��tS*����̹9�Sx_':�-�t��gB�]r��25	A�suVHLh�l�(qUeWC�b��$�G�;�5DJ�5���o68=��Ԅ �]�WGb�M��Yˋ�.�A���NH�d*�~�ym�Ǧ�SSٍ�`�#a�(e�)�di �8x܀���FA�bZˇ�}��Oma�`e3���dqj~��̾�{�0CR��{�}�U<�a��	�a�D,��+8Zj������b�
�U>��%L_��ˮF+�5z[hc���u.��7�t�ݷ!��d�h,�{���.w\�eވ�9�2Xc�ˆ��C�Wʚ��}x�Z�\og:J���OD�.�u�������d�Ҩ3����;�t7�Ƥ����Gy}�t��N�f��? Vj�y!Q����ڦ�9�J�O�lq�N�3<�ܳ,3��g1qֻ�vб/Y��3�����z�l�Ւ.�p���YZ��B��.6�f����t����y�ν��բ��h�K���B:+Sګ\��7fM�0�A!�'��{�N78t5~�ü0B��Qq��D&��2;[$�<�4�"dc�����vsx�vƶ�u�]��K�ġ!�rA^:���Zfj�X\Y���<yC�s�W2U�bˇ�$��pg�)$mgp��,؀Fx2Y�������6��U����X5 І��o�v�Nk���5V��6f�\��ӌjU��>M��Pd�-��%t�
���z�o�\�pB�TB};HS�Z��V'�TE���쐡�!0��;#��m~���(�I���V%Mv";�9�<ޥ,�`�&uȑ.�Ǟ��J������:/��'�O=��>x�Juk�S*H�k>ۿ}3�伌�A����u�-'�~X�n�8�&��nnc��$v���Ε(��"��/Uo�eWY�ۗ��iNj�[��9t��\����7W�3P@#�Xvfҙv�c��x�l=�t�O����YN4�]c���o9����!���3�Η��.p�]��Sk�����y�P(�S	�4F�|�u�n�0�/�;�uǺ�ɓv+�B�PE]��ĂX�X �>J���U𸝌"�b�_���Q.ϡ�ܴ\>�=�FuSm�9VI��30/F�pCQl�A�tq��^����a'�]Y��|�Ƽ553�+�'ٞ��ל��8����J���JAD߲�Y�S���[����21�Q�-�@!w/
�p{�*QizϾ�o�_n�ϋS�H�r��E1�d�5��I�b0i�ҟG�HNP�i��?]��|�]�>��������29ȰgF�b�G�e��nx�2F��֨f�4�F����i輇��Y��.��b���E�N֪3�`})�?0՟j�G��{6C���!�u�q٬7�N�B.C����*d-ȵ�\�$���⎏��?8��nlpAa~��6߲C�{Jqg(~�=�l��':��t�K�
�`��f�BN8 ��S�N��d=J�E�+��Ce�*O��,��t�g�^C��3Ee;�G���hٞ^��m�%@xk���,H����&1e�^�}�MZ��՗�bo�a�p;1e�6��ֳ�����cW�*J��WUG��14��C���[��c���a��ypC~�}=�q"�<E|u�M�u�ݛ��Xc h�(خL���G�D��	��9u. �ޝ�4����� ��Z��v��dR])Wk� _f=[,��	��iY�u ���x�?��WV �1-.o3��7��G��#�(abf�%c**چ�!?5���zYYRY6T�痌����1&7����%o���:�0����z|9�!�Q�ȳ���C� ��(����C�0�"(p�:�&=�0=�'�_��[%��R�N���&����W��?6���%Gs#^����귙\˵뉑\�QN-�(��v_���}�B~z�_B�7<�m�(N���FF҆@�U��8LR�)9Q!���>�:]�>;� @A�v!?n�l�jn�����O�@�[�%�x�i�I��Ͳ.��l\�n��r'��ew�a/	JC�%���G,�el�(����sE���l��F��aTrW<�f�'���]�	&�9�=�|oY��y��1��ܔ�D��-�����&��=ά�в^8�⨰��̤�U�;{^9�QɱGk�g+��&P\<���
��?�uH���i�j�Q+\u��\�0o*(e���d��^���n�/�dpˑe�*	dc�btZ� 8^�O]�'Hó�g���3���ŧ�����y� wn��=6�u�9h�<*�����O��n M(�=���wv+����� ۢ{̻!7��U���}pM���>���S�,p�%2H��h�t�T7�vi�;uՑ긑C!��*�3X������_�,W��7��,��A��`�4w�^Y��<#1�o���6�f�1rٳ���uP+c`BN0k���vN�K;|w,Z�p�o���ڃ�jf�zC6Y���E�]�q�;ku���v[QZ��BO�\E�1��m�
�#{go���w3�r��ci��L�3)�M��� �~�Pi��O���U�6����nL2nd���� ̨(pw��̛�矮�C�����x&��s�pЉ�74k`���TWeZ�`�~�Xxz�w��S�>��rw_ ��j��UK[P\�.{��TS��\ʢqv?q�&�bP�Amw8zz(�$Kzb�n(*�p~>>��#�ly��ږ潣���,���[vݑ��൱yʂ�B�ߕvл ���V��Ol����I�逐�D�:�k89���wH����R��0D�V^%:*;ѽ"���-j����/% �;U�,���8��v��74䨐��<����� p��^�锝g�ĲN���L�#I�<���2a:ӵ6�]�Z��m��YQ�|�/k!C!��Dk_��bq�B')C�dRt��z�]g���P����8�[�o���yNb쏡���=�]��؃�h�Q@��F࢔:pEqSBaca	�T�s��\r���t���C��F�d�H�7���PT�@ڛ6���K]���u��\D��]ʰ�;�0d����m廲��ع%�����	�@HH�J"� bX 	�'n�1�^�9��� �lxp�Ђ�li�IcbL�ʀ[u��.���ʮ��,ŧ棌ڈޘx�|#��g��]i�BO���&�!q�0F�W�f��56���h\^Dlsɧ��1)k���3�h�r�tB.f���z��`j�ߜ!�YLF;;Zˇ�t�����s��[�a�f�6���[�n������%�^�(�u,�]�q�t�A��`x>����=�3�_ݼ�Ũ�d�6��b��I���:�oܧӯ�#�����w���M�a��*OV]�<h]��/k�9�Q�8�p	���Y�0��8�<b� �b�fͣσ6vt6n�̏7�n#�X�o�|�_�����!�d�c��HrC���0=��S#vpeꙇ�����(d=O���2"��~�
c��a�|1��g�	��_������$��;�Х�Ŝ�8�c��u��䂫u��)i�5B�������bţ�GO��佟�u�C/��P_�{�FfHX�q4�ovPeK'�v��\W)SI�F@�����j{��׺�A�p����&����OI�.�{�^8)_n�
_�my�����BW�m��c9qz�;���'�ᦥ*�7\@���l�Ƈl�K�`�|���W�s\ZԠ��%d�����'���ٺ��h�0Q�R�@��sm�Tn���͛ǿ�w�nG/Xͱ�7��#��)@
�|��{s��~�o��j��W���=I�j+� �)6��(5H�ʄvG��UK�}SK�{��
l�8�X>�f3gvX�-`�a��"��ݲ|SͯЂqC�K$���+�i5�Gc�ܪ�n,m�s��}��i�Z��1��r'�P��>�xgd�*�N��D�VH�I�N᮫��	2�w�pX����rq�K��9�A�2l��m���ư�0RJ��㺕$���]�;)�hwY1]H˽w2�{��Eu�#����^vW=�gC�q���Λj.��e+z@�[r�fGb�2��-��='�YJ���y�K ��C�ܬ���Ԏ�w��؝5�%�O�Wh�Ӫh�����;z���J/� Y�X���\|��ׄ�/@ND��[��;�2"-� �v��ݛ_z�/�0%�&����I�^#&�o��C6_�$\C6���'Y6öF(�d�^�NGz��hU�:6������e�VJa�^#]k����Ɋ���4ヨ�(�>�(��^a\�&��yZ�������a}�d��g�㴒C�đ��LdT�V+=u�Þ3h���.���i܅���VzYGv��:k���*of��R�o�*
kH�y����o%�-����t����6��Y���7׆l����%����o��0ʃ�p#O���4��˷��S>�az��0�dz�X�@ Y���T�R$T^s���{�ߏ�������yÇ�6ڨ$�9Oa��
LL,sY#��A�߉{�cM5Y�{���pN4�=Є!�h�P��K1i���Z����5����^�>�vfۈg�oX���?�S��k�C�U?�fZ�h�oI.�T� �9~C��؞���\���~u�U)����{�B�����1��U��j+�BA���W6�#8�^͜eY���Y �;T��T�]m���{��8F����L*f�yQV�5A	��� ��@�T��z���6��Zf�[peh�����_5Kӫ�	��M��C����dY⼻C� ��E'[�V'��v�:c*6�\�E)�A_ϥ�F�vL=5�xSK;s�R���չ8<3��p��,�<;�k0J�ȞZ-���1�HеaU��:m��ȶ�]8ސC�X�H8��!�$��fk���i�ϫ8����1J!��4i2��c�E'�
�@�t�z�o�\W� D ��Z�T�s,އ���%on�P%�eHО��Ǝ*���R���=��u��a�rۑ21�±z��`�@���U��eB��o�����&�D�lGg�Ņ�&EC7Өh~�]m���j��mO�c�}�w�=�t�o>��nv�{��W�ê�Αf^���Fm�,,�[yJ��x-�]\C&L��2v3�/�<��������ɜ+oo��Zz�Cn�t���"{OT'-۪eDd�^ZL�ȥ���^�R��YG��A��oY��5w�C���]�}���Q���IL$��4�|z���!�B��1��B���jVx��-|�e�QR�T�	X{Vѥς�Z����)M�'u[}��He�}VEdѸ3������|h��<,/i91�۶#�X����;��\ͧ�)�8;�*<p�ǔaP�I�S�=<x���F��@���s�O�����$S�_2��(#��yXWj�.�e�\����3x���O��at�^5��qy���=ƅ�t��MW]Y=�}��vN����CiG�v����H�����^�_j{��M�av-���{蠯��:�̻$�*���mk��*����7�jq�@����YWe��n�P�(gK�B���
�}ѡ����OM||��Q�YN���ݷ�I�%[M�*���v�M<���`��1�6�"���mX]�-m��_P옥�&D���P^n�LV<�ھ�\�e�L<�Ml.\]5[;.��^jaun�N�:�-"��k,M�*��3�u�ݽ#B\�e�����:�X�ju _KkNF3��V}0,�p�\Gnm@RC)�L-� ��8�A��V4��i:�P~�t���x�2���N(�W�k���C0��� �_1XvD�a�+hl��\���f�} �k^��s�BCn������r_h\!�,�+��kNJ:��'Um�5K�(^�s����_^z�t^T��wH$C�H˽�K�h}��9�h������9�n�R왗W�>w��^H�,c��Zed�0�����4w��v���ޡ��>�4�
*�m��gopO���=�=v���)�)�ږ��s���FU�2�!�;�g.ެ�b\Y��Ņ��W��ӗa��_�Dފ��O��܃����=���{dqQ���p�޶א{t{����+[�W�����{��w��cW�'�S"u撕�:�z��s�<9ieY|b�"F..���S��}=j��4|�-ܺ�X;wjf�u���B,x�"�����v:4�*���Q�/��,z��"x�:b�j�%xd;��Y� �3x@�����2��씫�����̀����e��L��er�][����+�P����64w�<:{^�dpj��x
� �����b���w8b�����w�S���>��bӎ���ϥ3��^ ����{U0WS例p�l2:,M�Hk���ʙ���t�EAP�]�2�&޳Zrp�Wl�(�G*�M�����Y�T��t��ʷ9��*Ea1�|��Ox"":G���"��lN�@b���J���h(��͕��)*�<<>�N�ϩq��֩B�������ʓT�t����Ӥ�Bz�J�Q�.��Դ��FÃ��N�:v��"�"iJi��^]RSDKAA@�AT�Z
ZB���çN�N�^��E2��KCPSHҔ�(D�E4�-�SA@�#��	�)(�bZ6�44P%	E!E%ECCICE0�R�	A5 RЕK]6Jb$�(���h)b
��(h��e��<�$�)�h���()j�b)(~/��7������"���7�1`�GC��s���H<�e5�y렧TE���p���2�YT�k�]�FL�[��7Y,������J����E(R�� 1���,��t��f��߃$���ĨYB��L$�-yj�^x�7 ��0w��'�mЋTe�8Geg�H��u�,:ǎS;�9��F.���f�bN��kU�9������ɟX��8EGan�fP^ ��pVle�-0&4:�smv��(��8�X�hŮ�mؘ��ڷ��K�_����Bi�A.�9��B,1��,�z���l1�U%]CV�o�o�k@�p��2�Uc����;O�����,����!'l�=��.2;^������Q������jY����K7H;�XW��.�ٰ�ڑ��m����(�VYҙ�϶�J�-TT�ծc�z�!�mס�_W�nq���f�d<w@<��F]�Qq���≧N�0�['>�&hQO~�:5��!d��uN�Y�ׇ1{��vA�\0d;.������L�tͣ�m���Oi|kc����K)��A�}�c̕�"�;@ʨl��1�����oݵ����4�n�d��6�E�T9��g�!64��i����S��n�;��a�Ә�i�ޮ��acZb�����D+ԗe�<y�]��tZ���{�����(���]r��߮�[;��U=�D,0@�z�Ҷ�U�E}+A�!U��CP"��1W[�'q�����S�چ2���s�>�+6�P���/-Z��O���xO�^&k�����d|33�0`�B$h���(O3{� )X	���j��:"u��2*��P��z;lf L�=cռ51��>ݥ��b���,s�^������!�^�� �:9���	L��N�%�i�ޑK�4�֯��HB󨺅�Y����yk2M��hs�XW Í��qðϰwL�� /�:�7E2H�`���<��n}~���ܭU{��ߞ/�.,A�f���2�2е�I�`qi޻b����(���Q������5x�otT�����>��)i�R\p�'�`\ǲzBcGn�;JUYU��0�v5�MU|Ы^�b��v�j4�ܜK��w8Xɼ1�6C�ɋ��ճF���hM}H�=��ۈZR�/V���ں����0�('�8A�=�����]k7֞���A��god>i��I���U�Kn�v*Ϻ�	��S܌z!f85r�������x)~x?}����vm��ޛe`ʤ��x�}��}fy��,ƌXgc����ڏN�Sf_C���\	��8������P�s�%��y��Y�jv�
sK����`D�:OK�p���s��s���j��n���V���z>���wd�[�ɤS
ӛ��v�7[K$�T���n7`���u�'�8`���IR#{����x'`�N-��
��,CUO`{�طs�^�F�r�� =+62y�`Zy�t�{{w�ώ�m�o~\�cB��J#���Ā�4�C2���x 0����dX�ՅsP��[�2�G�q&80�Dy	�ϥ�\皾X	��}�X��OA!��h9[
�l]�_�jʽ�U�9��\�Z�I�[���o@�W�̎}0�=��O�큙#	z��NSZ�:�h��k�ݩ��0<7�#���Ԃ�^���9�j
z��22��S�=1:T]3XNa�+5{���nEK6��A���W�;TC�ͧ��V�S�`qm��{ p�t��s�Q����N�0�~ڊ��!)���j��Q�"XnK��iM'�8<2�Cb�V)�Z��� ��. q�b�N*���ĲO~H�2�����5-��
7h�n�_[�?��(>C,s�"r���;'�Q�4�5'��N���5]�9�cL׫�W��N�a�����+�^�C�g�����v����$} �O����7��F�F+yC�P�[.��+�,n�J���e�_ڥy�\1T�Ã��#�5FAi�o*���ݮ�X��{R�iY	�^�E�匤���:��[
����s���k\���H���Q��J �Ho7n�&5I&��*��������q�w�?y׭)��p��A���A�٭Vdٶ��n��ܰt�����M�چh��s���+9"v6��}^rW�$���u�43�q��Sˬ��)��Fj�r��m�_����F�T� �` `A 3 � �Ů����u�=k�q���mNf�[��W5߰�/�R5�=Λ�i�wn|ga�Ԅ-��0��c���� B�(tmvLd����0)�5�vzRr،y4�Ƣ�8�0LW�d�z�����0WRD�K�P�XC��C�k�k�S�W9�"���8������/����vlE\C�̧��S��tE�}�b �
z�3�Da�r�7�B6��\G�*f�<a(���/���.:��25`��F�	(�X>~1��/^�~�ͺ�ƥ����9\���ף�Pi���q�m�??$ ��~T9KOհD��_����^��  ��z}]����5�ڮ��eo��>�P͹�$��7.�coC]Җ��f�JUeWu,����K������HZ#X@{�b��|�؛ja �BZ��A�#8�C6q��ܗ�5��SB��z�e�D!L��[Ӽp�#$���¦nA7�m�Ȑ�[�jOAd<#Ӱ2taA��j�~O��M��R�J�z�Bu�N	MÜU���!��{<U%���e��m�Lɇd^�N�����dޙ���03O+י�(�vǲ�j�*E�3�YQ<����L=ӎ*�N�P�yy��}�JĄ�L�[�0�e�k�2c�պH&�\�<�O��/��oqd^)��5�!���wvf���o�o�ׯ� ��0 �Afd"P
A"`��P��� �����̝M��]�\vD�Ҩ�'���y�^�t�����Y�>�5"�FP����`�ߒV�yާڿu˿Zn�����4-Z�)�ߣ��H�hT:q��gd���c��5�L-�nurz�P׳e��3 �*L��hj	�g�Ȥ���b:l�6S��v��,�.Ŧ����2�᯦`\�e֦ʔ����*09�Ù���}5ώ��ڵ�BӠ�=�N��g@�l�s ��XChcȅ��)a��i�}"v��NU����$��Ic�W�㛫U���ς��GH���(����B��"n/Bz+��xq��qw�*�SwӢ��V�ε���!�ȵJ�e��\��`�Zz��6>^�c���4�s�>9�k�k�(��y�\�{�����h��6�=�2�����r69����l�Ut�Օ[��0�E��I�e�H'��k_��Fq�mbz��^�9�"]����|r0Q���;kt`� �0�y��n��XbK�v8�	�v:�����oU��+5��l��>0���{�E��9����]voMwm^w|�v[:d
�"{�Ow��U���4�q\6;ڝ���*��r��S0{f�w��B��Çʻ�*+Y?��x"���`��3ϵ��Y�:	Ӯ�bn�Q�<��,%\�����LX4��O�*[��ې�<΢��}_U}�U���#B� ,BA
�K	f    �ܸz#F���D8���(��a6\���wQ!�;�N�t��Tyv},�?emĻp톪���|'9�ⓞ�n	CÜDpz� 	�_|��ޫ9�΁�����;�,~�F�:[WFb�z4��>d.2�5tŵ�P��v�!���b�ᮼ���-����۲ݻ2�ß��t9GK*	�};PY����]�6�2�"���?B�ag�}E̿��U�>����}��*��W��)��	�ya�����T7#֧�i9�TQv�F:m;�$�;�^�(ӛ�(D��q|��pi�!QkhJe~/��c�%P����=k�<'h�}9vKo���T����k��0�Ʋ�i��=Ƃ�a�gt�N���Y'X��#)��7>!�ٱ]�A��:E���z.d؍me@�6Ϣ^�T ��@�nT>��r�ʥYY�ۃ �۝w�w�J��������� $+wVю���"��ۡF�҇���9���Z�su���Sk��t��M`w���� �-¸!�0�}=Sey}�3{��i��hM��{);M�=���+�B���p{�m�c��)��L+/kZb���`�[�N�+�X��^TVY����;���T�/U:�7]��+U7vT�e��Ë��;Q��z�A�a�ٹ�I�VC��r麷��%�[)m��1��D�G��_�"Q"H����V "P�@V��P���"Pz������x���)2�Z�Ы���Adi/N7 8��k�ãԫ '�j�|k,�{z0(��6����T��(S�4���S��)���<�=�	�TB��6�*���W�k�̽_p��� :���C��i&��E�N�e{*��)����z1��3�^;r�gk��$u��,9>���G���D	�����GjE�^�l�<���7m��Օ��4)l- 贋�M���2��W�歱�z%�,+��%M��;��x�g۵���Q�uZ���q�fP���Y���ަ|tR�`kt�P�
���A�al��=cь�B��QXr��B�b�h���`h%��R]���*��f�U�Ś�|�?}��g�'Hҡ,�g���z�U�}Bj}8���c�K6����å;A�6m=z��]"���Ь�htT�˪�mo��<A#��y��q��41�=���!6q���؞O��Fڪd��طī�z�Q��x�Չ1��2`p�H�����l)���A8�Q,��Fi��4�~�x��?X{Xc���RiQ	�nlѪ��f�����i>#%K3���Q��~|�Y�+|ρ�ꧡ�½�]��A���wR�xő@'}��6��S�S���8�E97�<L�X6X�f��q+�cP��Y�B^S0/㷿���k������Ƿ�>��R!R�T�h �@���DiEP�H�ǯoz����|����0�Xhr��Tm+��d��"r��`��3ݒy��%:Nƍ�g��k=�l���=#�����SA�5��d�>R뽎�8�&�?tssK{`��ͥch�W����w���>��U��E'+�R�-�a�@_͏��a�<��r!6�~r��N��H�N�j���ٶ��t�6� �2���>���T�x#qx��(�������Y���y�`�!���*ɨ��2�p�lv����g�N��)a�ɐ�mxH߽Q���//�d��SW��IDp��<�-SC�~5=B���ԊcFMc]����،�y�J|�(�f���u���^I�4�牿������r��p9�k�k�8��i�j�Ja�Ʋק"� �(�Q5���'R�O|g�e�{C�U6�\3.�
v�� :��R.\�͐��Xe0�I.ե���O#.7D�^����y�:�R�!�PH8��8��Q}1��/���{��}5 +«gם���!��u/>pЊ �����o.�{C�..��l%�!�5M+���<�SF�~|�;��l��4��3Ș���Ź��1�����9E�*J�C�b�d�5�"�I�S42﹪�H3�ݲ�ђ�g�o	��2|�Mm̰�	/p
��l�����KV�+3��+U�����c���mб.��
�����/�y�N������� H	D�1(��@� 4"��}�kd:�x~׿�58�nsú}�i�(oI.���a�E�����^q�nv���UO<Z�%�
���<�ڞ�*�}]��m�b���!-Id�ԑ�g���fE�2�-pʺ:8;)n�lY\�T���ɖ�|�5����%�M�C���P�|k;'1Abe`ˊi���^���ҽk�Y������r�HE��|�LbB9�Ϻi����.�����w�^F>��f|p�3륱\���:t�3��񜗧]-O❠>��MP�yڪ��
�m�՝��fbf���ɩ�I��Jt��TWe8��6���BΜo@��c[��RM�wV���7�o\��	��ʬ�1p�1這1^/1U�򑽛#i�+T��I��{�ux�����Sw�3^0D�z�РA��s�=YS��)=X�6Ⱥ�09�s@Ӹ;Tv8�w�OV׷	����O���!�׸r�tXQI���P�~i0� �yj�r��\��,�jx3�\�~љӂ����td|&�,glZ� ��:nw	�荮��V]7�u��<�[>1���v�ʕ�m�F�3��AX�e��:�n;���\�xv���>��[E[ވ�n��:��Gټ��4��뾥�'.
#�[|� 뗮m]�l�ީ
�A���c�"�Ao��w�AR�/S.Z���7JC�9���=����||{�s�{n�}��"��D�"�H0 ЂBK0`K30Q5ڶ�7�+�b7��v#c�|r�
����g��L�_��8����Pw(�Us��\��8�%k��VGb���Ti��ۀ�p�K0c���v>�<�z�QT#�������%�_����Գ�T�sQԨ	�k^�C��l9�`jEj� ����SE7�z�X��;w�$a��a <Fۛ�T�rs}�����me���&e��zc��x�4�c���^�g\$�\�T%cP�B1<��|a[78����3�x���e@A��MoA\�k���8N�v�LW�&�P��0!��c2R{��Ƕ�{m�HxnB��`u@nJ���Y�n2#��V%��Ek�"�)�P�ê6��
����ܯ+�xk�@��$�+�����#1c[/.2;���=-ީ��;��zf|�"*]l�y+�M�~�0Z����Y��
kQW*��5j]���.���O�܄.} �XdJ����Xg5�cռ4�{gjMXk��B���;wH��rīe�'3mL�o��4�(�f�!2��)Ղ��M@)�U��9��`{�B��5mY�z�n�Зj�b�.`n�GVAk{��݊�
�ª󱻷t��ݮ9y�zM_]�FV����9l��6���9�
�Z��/�M����n;�ܓ�Q���ip#�"2Lԗ!k�B���ރ�0S�j����TB�#"�Z�]B�}�}m��y��X"�v2�:�
2Wm�ړ8i�w}c��a�H�P[���uS{d�Y ��g�)�u��m�5-�;���ib�i���}�ݖ����vU�c�i%n�*Ժ���m<[���n���a�ʗ��O��p�F��^�'��Z�OLҠ�aJ��W�I���j_jV��u���ːy��>nP}|ʾm�U�c���wb�N�]�θX�tF�q��%�pκ�ˊyތ����~���;&��H7�?�<\;�a�EXor��{�.�ۺS�8�S�k2g��/*W��"R���8w|�q븶��2<Y����%_#���3����5�i��ՓLDj�k˼�"{�;�#����bm>�ݑ,B�Mz�Dv��n�X3���ƍa��x��äu/$ɹ���Ɗ횉l��.nr�:��d�ެ��v�6	��{|#� �3�I�\p�p��7�'��=��-܏8��~����U��5�<����[��u�n��L�V^��973~���nWld�E�䄎�/�v���w��@�۾�7/�M�t!3�3j�Л�V�ڝ�QwA����^��/,Y�52�9q�&���wG��k���cŇ;T�FS~n_�i���`Ȏ��N�%�r�B���Zw+�e?{���ˇ���� Mfݾ��i��u�-,��o���/�
_əhh2T��p�w_c�����5\�N��H52s�(n�Ĩ����kF����W>{)�,:C
).��s�'�}7=��.��������7D_�<�V�L�aXgb��2�s��>.�8�Rv1�����]j�l3�y���>FzL;R_9:�>G�பvL[��O(��U8�8��'������k����?}Ú�^%�fy����6{ei�+'"�v_@.�����Pz�!�'�Ɋ`kj$kX}���TE.�D�	2U��Pž���ӲFVcp�SS%����م�r��Y�g#)�����u�?X��ib�t�UMpfT��G�\UjG�Ri!،Gk�c���s*w>�����ۚ�	�ؗ�tct⛙���VeMGQ�{�Q����s�2g�؃�1/`�NV�P����Y&���o���Q��-֫�[�c�����*r�S�6�E��N��kD]�P��'�)x��Il�@Ý�~��6��\�P�K)�����6�vK]25���]�[���`AZ�9�{U݆�7������.]a��l��2�Z�f�2Rx�m�ʎw7�\N�e]�������3]+�p��)mH��br���z�����-���Q0DӐ.)��'����)��,1L�)3r���AQJPZ�)�������M)(�"B����z=%�
"B������j��b�3� �
�%�#�N�:��)�i((h"
JX� �������ӧN��ZZM���
*����"B��j�鎝:t���j��h��Bj��)�:JJ)
��)B�H�4�BTAM-D�t&��CTB�QM!KT!E4m�(����#mR4D��I�J��MII�4�@L�4ATRM:1,JSUT��RP푠+@b(X�>*���b���Ƞ�>�4U�/%0���{A^cݩP[/Q\�@���t�dӵ��X�C�9�\�wv�z����@�<���#$H��0�*��!H�z��|�{�����a�R/���GOhUfh�9����5��I��d�ctUYM9/���+��Z�>:�ϱ|��`��׆�]�,D&����4��Tr�?g��W#���ޥ-��<���E7a�v��V�A�A%ۇ9>+㞌��gn�Q�T$/�6�5gk�f?����{HE���a�n��Xdr��A]�c..k��5� �ʭy�@�ݍ����k;5md,������~%Q��-Gs��+�ܨ}�q�T�cq �?��;��V:>�U�g1S%���p��h����-l�)�	�L9�r^�ϩG-n�A�!y�G;�NmW�=T�}����]{���8Xj�G�oA��M�"�����Ó䫠ٰ�j[6#	�[qaa�xC��Gm,��g���
=��5ڠQ��T�.yd��&�=�)�;F�*�t��8������n���+׎�A�=A#�s�?��B�<ē�e�v3],&�v�xttN@1'�V4��!�X`CfC��Rh���y9U�����Ϧ��_&��B�EV���4������5�r��i��3ȳ�BĎ��*u���7��{���(��B�L\��o7���i#�_
�^�v~���#�ё���~!�;g6�'b�r\1Vgc���+��7r4��
%}s#�8֝�ce��$.[udqT/k���r�w�מ��z���׷}��>�b"D"D�T�F�RH)D(T*��y&g�7V��}ʇ4��h�vIa�;�#��F�y痱E'0-AN���9��C���X�3���u���)��Ҟ��͵IS7Y�L�,�`��(��ٴ��z���N�F�6=���n*ro]pIP"�֡��4KGO��r����M�8��щOҺq���-�g
��`����.�q�!�|6&����<B��0D�� $v�!�N��A8�Q,��*�y�}��w��z��5)]\�p�4W�+�Ơ��6|�Ȝ��������d�x��(�zl�g�PUݑ:�%�]<��H�IMM�;'���\:���8�&�3�A7"�0�j�?��#����W����83�a	\�q$Ѥ�E'=������F��T���!��~
7�%���<L5��D3�&�{t̸R���i�^:�NBn�����e ��P;��a>=���ɑ �7��?��dCJ�ΰr��wD��������/-Ha����"�}w�o��F�)�^���w�|���E���L�>��e��y쟍OP�u`Ԋb`͵����ϩGCG�����e�[�mL(m��[d�����_��	}�pi�7���X{�n��}�d�7��
B�^ׅ�&4�{K����ۄi$�E/`}{In���Ժ{����7�`U}���nXa��`b=��lr��g7��6:5���#2��w�3? � ����Z�@�H���Qb�	f`�	�����<�. ��)�kr
�j����%�+��ch{��0��,=n�<�n���bcK7.m�]�9Q�8dj�p]������,,+B������ݨ_�v܌��*V��9w2�,n�B2��qź%���v��&kK����A �9V|9i{z�)j���P9v޼�a}�4��[����w�L�v��]�O��w�ޠxF�^xbڦh�y:?��~h{�>u�
d8l[<>X:�m���{2�3E�%ڊ�d��jljOQ�;�Z/D`�%�}����K��~���I?�5����d_*�}]c7�۵{$P91j	d�̽��7zb�)v)1�gL5l+gW����/���ƒ�1�ߔ��DP��&򢭨j���mΗ�N��=��q�"P<�ĺ���P7�����d�C�����.�~C|���O�a��m��:�4�̳s�؊V��ۏd�'VvȞ���$�5=��]K�xD�LiheY���E�deT�\ٕ;w��Z_�����	'����2O`�N�$hZ���qv�dA�쿹���5��np����VK����\�4�R�]��jTy�;��Ft�=�ź3|��]�Ӳ�	��]��3��->m�(&,�k�75>2��;R٥��t$��S[�2�>L��k�̳PvP=�y�˔/���'4M�t��l��π�7��� a D D��L�R��~7,s�(�C�7U�� �;p5M*Sx��y��W�(��ӓhT<~��7כ�{�2>�|�������^��ʎ*���R���E�`sre<�o5Þ+�̱Uc�G�$xmc�.K
�  ��:�ZeC	���H��;I�P9+�[�P�1tfU𥃟�ĝ���S*�;P�Bxwf�Kʂ��B ���$��8��jEn����maBr�#���D���qh.S�Wc����#�HVp�
��g$�g�w:��K&�����̬�h��3U)�c�-���*	��B~a����BY���	���y�7��~̱[��jY�h�,9�� ��5�c�;N����X���-A��M�d�sCV����n��ʬ��|-/�����V��ʖeί�Y�@;�XQ1%ڸ˱�-���x�ج/��k�z��{��(��R�����\8s����:�^"E��ds���c���;�SH~��|�7��~�����IK���ƀ�xe[�����B.<̄�T^=���5 #̚���.�v��{,"��Y�0v紌 �Zt���a<��ZF���A�1gM߻X�Z�i����I^��=76�S|t{ˌ��y��ea#Oy�Υ��r�c�x�'�\��ʝbp��S��zq�*O�����9��Q�^��o�����7Tv�I>�xxy���H$@1�ff`A�n�ֳ�G&3�s��|�VHB�5�\e:n��u��x ����w4^`��BEWk]��[\+5xSv��je�FB�a�d��O Up��2Q�з�����)O�}����fv�s���i����bv���܄&��! �=���vг�x��O���5zg,��+ �,b�
֟vXi��L��{^��=ا��L��JuiI`���B���c�����uaE�n�w3�MRsR�$�[�Pt0j�0=�KC]�n����t��j�J��<�>�s׀��1��:A�8�����"՗5��3���:��'Z-9J��1�F�_Eݨ����K��}:��:���oe�nQ���2�L����xF@��۬uNP��m��b����^�Up�ZU��,ŧ�I�I�栜K�����;c�����$�"Ў�1�H�v]�^Ͳ��٢�aT��t�`l����֟1tPꑘ��a��('k� �׷��e�dN��9{gÜ�pS���=�\K`o�RZ�%�B=+^�A/��?6��P�ve�_�F~��b�`W������˱j�3t���.�.�Xo�H5����ݎ�ܬt��L���P�n���Nq"��$e[ʳK�����E��Z͡Sq�T�/y��,�a�����M����፪��I*?�O�E�V  �"H���xtfa]tB�����H`�0t!�H�\lz���E����VB���E���n����Ӣ���0�V�3�z�9�mpJ���ڨ:�^�W.yd�5v���N���L$疧�����9�p�r3^Zl<�22����	; �{C�q1����x��t���h���5��b��o[�����E��.�}�{ތ���k��5�1���z��y�n��b�앓���T��Ȳ��ui��L�C�KIe+��p�x�m<��y�mAOy|V�hړ�VO���PT���22�]T�Sн���)S7Y�A�
Y�1G$>�ٴ��d��
��`�T{��ù�	�	Gى�à���,�a�{%��½*��V6��#��M�aMK�K��%�R�=u>�g�#�k�`�{�m4�Ϟ��x(�ᅾ��R24P����A؞zar�����=�Ҹ�;Q�<j��yxᒹd�Jq�9L'f��_<Yr�ĸ�x@l���l��X����|�@�Juk�S)n�4i�=d/=:�MAƹ4c�A7�{�������R�j%�����;�l;�Y�@��"��y' �};�����Q���{�s��)(��y،:����7k��4a]��ϱ�����:�%�>��Ǜ��<J��Mk�V�BҳO��\�h�U�p읏QW����O�����0,`"�%�	��w��>7���Ϟ����,��3��$������WKu��F��T����t !�ZtAuk������l����C�m�9���rt�q�O�H%�yHA�YC1L�h4�K�&r�s8��)�s��l�:�DtK"�j曯9�s]���V�kO��)��+F�볆�\�O<����ʪ^���!�q"��D1�X�|���a�?��\��H�&U�z�NZT�J��sm$�&�y�t;3�0ti�}�1�m�"n�p,#A�T���zP��C�еR��P�wKK����
�9�F���v�q�/k���h!��D�����t�:��Z�i�{�y&'�t;����"9���i��
��w��:<�Z�+	ɕZ~��6"υ_J��i��`�Vl�aAۗt���w�f��Z]�H��E�sͼ-s�O(
��e�!n�e�ഈ�E�L[m9��>̳,ѽ��*q�j�e�cde����b�muga���o6𵈖bo��,v~�uW?WX�u��(H8�rb����ī�m�ݪ�j�=�'0mM�/J��?JQ�1��[��;�_�l�'�	�l���g��q��,�mwv�����NV�9�1���r�n��_%j���Sq���bY��nά�K[Wt.�dj�d=�Ur��wV]M� ��f �10 �` �K����{z���uǊ��0��Q^X;�����6hr�5�5��NH&�TU���q9�
��c��f�G>2�����������ơ�j���>�&-i�>����xޯ�me��J%Yq�p�~~�,����α��,)�\[gT\:�pF�PyoZ�f��ݒ�#^E)ܜ�Ւ�zc��},�'�SsS�&I��"UB%��ł��qw6�{"�ݔ��P�A�;*b�'&.�Msani�7�
{|�VA.Bq�f|z�&E�&)y��2
�`B15�W�f9U�Wp�uR���o'2�i�'��T��;YS�vT���{WE��z��7%^TRQ��ނ�����"qJXV(*/����S�I��׮���L(�p��e�βe�}���m'^S�]s��ҒƂ;P�rt�|�(d���C�㚤4c�::���3��F�U^�78��Z��ti+�0�GE�yL㘩dcB��mnnL��9���"٭��L`u-�&�@-T-_�J�e�W=�������Aڢ�^�^d���ߐq��¬��_�+�Z��,3*fu`2��������P�/{[��%��T�=�0�-�m�q�͗@�X�G��g�|kl�t�B��I�+����H���������N9L��|Ϟ��_\�j`��Ԅ@ie��VO8�c�۹;�[�U�.k�}	�JD�2���xG��Ĺ�/3|�M>���V��s�#�t�Yt��F.[6`�����]7�����ϐM�\���<&$��h\D��t��z`��ՙ�����k�.�]m��g��6fP�A}��xL"�¸Hz�������W��py��a@��w0�����1߂kk'��[Q�&P��\�Z���PUK�cetM�1�����q���);ت�ǶU�К ٪�&��#/qg�W�^���ò�J�!�DךE�S�����E<�1a}���9yaY���˺����&u�TsV��56R>A�.��Ty����	��T9זt�Wp��S�\�gn�>��x�2��C��`z��+�-��D&�d&U内'�*�l%�v�Ϫ������پ'�i��k�}�$��p��}^!��O4��%2�^%?ZRX&���z�)�i�ʦ٠�Ps�<�0���k��4<��>W�`��;z}�2���:Ǝ�����x�7�v߬���\�OɔSuy#I��z�K�/5�.�0lr��D✗�M u�J�ȁ���d����:�P���/�w��h�?y�S�= �7ײ�� �]Z����'�!��/�V�ղ�Y�
��E Q�aܾE�{z;�sB�_dDbs��S��Ϋ&��{RTvnx��ˉ�u���7��L�+��s];�)����� ����0 �13 X�`�a����羷_��ȦΘ�]�q���!���ZI� ��3cH���M��Qc�Q�ӽ�[CZݺ�ɇ�U��^��pJz������c����O�b��3m�#��B�,��#�Fǥ9�%��:rEo�Te�Z��R�Gs�Y�KӇ��[�؉j9�(��.w�!B�ã��ֹ�����UQke`)U�(zW9NPQt��q�\�=�l�[�K?	5FsݶQ�&���]ntc��5C:6���7��dQ�m��;\�%^X�X��}On�p�>�trgt=��f5qa��p�\���C:�^�W.yeۂm�� g_P�3���њ2��L�9^ǏD�Š����aAӒ;���M��A?=j�\�t��^&�u^o��[O����e>ݯ���
Fiq��˘�b����K��e�������8鉛`�ٷ���2�-����{=���4��%��%���K�{Ȥ��ON��0Α��UcߺS��w��+�a�a�@��N�R��O��^�6�5%L�geT�q�2b��w��_��G�t��i}`�h���}r�#�c���צ*]O�r���+`R"�g�Bn��0��HmX�ӡ�@?K�Q@&�ݾ1�8v&L_~�[��k�z���7�vw(�^�VX5��u��9w�Q;WjLǥ>r�����}�#ɐ��d�| ��W���?eݨz�Ǯ������CyA\cWL35S5�4��Y��s; ��snrG&��c@�Ҟ�j������;�� ��vD́�m֎V�J'ob8�����i���f�h� ҞoL�B�u�z2��7�׳�V��CV��G���+	(�,���e�8ޅt;�^��{�^���ܼ)�
Dз��GkdۢL�:�$ځ䵺.�;Y{WA%Y�u-g����[�k�o*�8wE�j�oFW0s0�[��z�|��&����!+�ל�xv�E�|zpz�mgi�y��7��YC���� �5�w��K�=�5���P��=�!&�]�8kr��=��\�W@ Kf�#s-l�=�s�nk3_5���;�B�S`�iFzW\0o��Ֆ�ٮ]0�l��:���+9�#z���qD���k"l�+�<�l���w�<{yb���t�!rߋ�W9J�q�k�O�r[��ww}���h{Y-��Ar���e����U�bvG��N�R�Σ�!2�vyX�vݔN��[�ܷw����2#j(Nn�@��mL��X�'�lWv�ވ��:XyV��8��q��0�: �S�p��%�܉��[��
��cz��j�E�p��v���y�{�Ά���{B[�ֽ�f.��R������v��v3�
��^�͗$s�H�8-��(bӽ]B/���Y��	Q�&@����11���]Q���`ΨV-�Ҩ�D�$��Mz1gA������Qk�{�iL�zb�d��}759r�U���$��M3����Y�{��VL�|JbZeܚi�&���~$��J�u��7u�0h��q�a0��k}�Q3&��
��U�U�|4%}ܧ�#Yu���-ߨ�4n�+��70�e8��6�%�d�s9p����2=��A��z72��R
%Ô��.��n��n���V��%���,�}F��vW��^b�@]o�.<$�S7U�e��G@=[�t��M[�]���f��2�0�˞OynZ�%�E��K坻��STc�+�7�;^���#n����'e��C��t)��������Ɔ
�R�.�b ����=�ohIv�lr��S��Mp�c�J�&:�^>�,����ǵuo_;��J�T���iE����C��w��h@��8��i��RM�����j�5.h^��t�G��'��8��H�����yw6�f��ޏi.(���u.�:���ݜ%��W�=N*��݂l������L ��.����.�72��)R1��`��1�={�y�|�@P�ATE�w�� ���z>N��&�ZJ
J�
B�iJB�h���Jb)�"�#�N�:u�%SSR�PT��m���h֨(�ӧN�P�D4SE0��3D�ڨ����*�:xt�ӧ`�]PSAT��j(�F�*
(���%6#���V�HU%@Q��J�Z�CB4R��:M:M-�K@P�):Ci4!4P1PkF�QtSDI@i�U�E%����4jH�IABhm��@�JV�AQD�U+K��+gU�HQEi�)��T%[[��H�M;ha%�oJLR|"���9��]���c�� G8	������Od�;ɯIe��r��muJ��.^�v�!+�۾{|{}�� bbD�B $�����g�b���|��);x!F�����%�Q^�;���`q�6�.��U��f��VU�n�)��[׻uoV�^���P2}�%��@$<�� ��U��O	�0�Z�ӳQ����b[R��=Q�<i,�Gب�P%RO\{��fxL&	�#�����
�fiv��	tėI��N�t�eA#I��Gd�;����c̛7{W����ٶ��ׇ�vi���RCmb�`d�'��$�E'+ n�J��0�A(���~��i�.�v-���ke������0G��Cq�q�����M��a����T6��r�H%�./#�2�ڛ��c��啜��u���!荂9��:ш+N{D��ګ��a�^-@�P��[�3<
O7��͞g�J��;Xe#�<(���:�����H�tf��鶫A'�^+y�_�g�7.��@.Rm��Nn��dS�D�[�V��>���ѵڥ�\⻇�{T��A�����lJaşYc�0��iʍyæ�&���@ǐ��p����=&C�z~��e�+Iu�&l�8�/hm)�rrwY�y��8�5�Jz6���h�ȯ]�W�&c[�ۍ�Kg羯�AIs�;5�,2�@����y� _:ҷ^5���u ����ۓu�P�V�һ�.w����&=$�+��v��3�.�v;Ճ��� |������4N��2�eCk��hGP;K���$H�.6�Ta�X)i�!!X���nT<AE��^�vz�m�x7z0Lf9�mH�G�C0��hEf��2�Z}��:��W����&'��zc	&�����!'�����<?r�R���wO�f_�����x}0��'�GΥ��W�.��8!;	�S�Zz�o
����k���� ңڼ�59L=o>21BA�Z�C\��ɴї5HZ�x�u���CVI^�g�b�o����z��ȇ�zaS7 �j`SН��p�X�e�"2�^�м�$s�`�'!d	e��QZ�_��*.ۆkA@��\c�3eKf�N]��Z���W�̚�dw=�A�=�QIՌF�+U�d�W����W����C�C^ˈ&�`��`�xu=A70�h���xFz8��r���_�F��2S��6������X��_J��g���}���ޏx��ЅÐ�=},�4����J�,�&+���cV�J��Gt4�F;�GM��|���؄��R/G`K*8�}�R�Ԅ��szTi��j�w�1 �Z��UJ̏{e+74�Լy���y�z��%[�6�XՍZ6������5�ɗնꫪb[�q5|$J�o)��ӯT�lCB�XƮ�M�/�8� �l]���}ӛ�/o�`�X��H�w][�^o��x�MB��>�A��.oJ�A&��۱��@-8�H���R�aX�E�:�:�s�c�-��k�E�jt�mw��E5-._29kC�x3]Qܣy��ۗ"��K�y@Axܰt�17n\��1jƱ�����r��ok�,��6���1'\⤰"�O2�zo��p/��ۅ�@��bI�$v)f���<s�-hecX�5 �� �\w�J�`�\�T���*:���{�@J�bG��-%������`K����r�as�ϲt�c�H)�'r�i���R�̛d\�������t^.aJ�]�B\5aqQoו,�:��,� �Qa^&$�kA�WR�kiW]���嵖t[�/�u���c��1e|��t���$���5>XEl��N{���W��jY9�����]�<'�������Pl9v�Z"�s�<1���`0&Be��3%'P�X�6���*����]袊!kn&~����������s�Y!
Dך�%�t=C���L�0A`���1�c"�HC/z�wr�d�Gd�=�5Բf�r����2���X�����똨s�>�)��*�a�6���W�b�@��w�~֢�Y�*Θ-Ek(	�us���zMG'�ON`d�͘���%�8>Ylu-�D�dG.�)İ�n���gf<3i���G!=�gV9�L��5v��9�5��:�P�2&S����<-��R��˳���Ɲ��˵b�d�v�������b��ԝW\��L�/1� �7t�վ��.��4²�
1�s�A�ƆHa�Pn�����W�^%:�?0]���Mμ#��XKwFd��{��~O�@��@H h���`������^���EcΎ���x�����P	L)�/�W��a=}h�a�&!0\��1ñ�"
�#{s}�.刚C�(y9]0�ʥY�'���f���)i�R_�9>1W����rܗ�q��G_n�E8R�Sr1���m����5W�*�{/I�pJ���BO��^�<vDD�>�*旅�r�2������D&��\��Ͱ-GNP��2�j;�M�]��kd��z��h�]�׹Z�����@`���ֿT��j�uQke~R�XR=+��PKܺ��Y��~�^���	��V�������r�pǢ�����T΍�1�{	/*��Ռ�%Rc�iG����JV��F�s��wd4Z���#���vu�wP&Y�k���C���W�ɝ=x�pFO�v���T�*�-��|�C�̌嫼�Y�"�%4;�S,ِΘg$ �5M5�������Y�'�Y҄
���:��f_9��D������(ɲ�+/7*ɛyemD"��FtK���"+#�`fV;�ܺ� 
�.N��+
��|��A�Z������t���F<$��,�8@"mv�f9��f����>�*�S���&C�X��OA!�qhf�􍈨udK<�$����|�go�Ϙ.GA��.Dx�P�=	�{9�C�}�����d�+����K�y���w�sF���"��m�CB�v~�O������X�/eT�9^�_��*f�;(2�,�`�a�R� �7�;�6�/�}�Tb�lb�O�:p6���0:ב�*��W���Jm�ݺm�
���J,�;�Xie�f��	=0�瘬�OߖZĘ��
��ؠ�?D��v�"31�muÊ���1����Q#\��? ��ebQ��b#����W)4��ܟQ>�dԞ�y������N�W���'�X����<b%9�.�L��Mmq�<��ȸu��0��yq����m�o���7o�=U~h�0R���J�|1���t�T���5^�N���v:b@s��3�_W�p!�����x-6��_�Lj���sN�S����R	v�������qXo���w�sg�㓅|�d�o.K.����:�";+�������0oO���<��h�M��U��ޮE�%�~Qi�E���u]a����jk���q����f�wSsr�	ON���|�T�ޖ�ռ�Ͽ�2�E��֜���G}fi����E�R(ց����])�ݟM5សy=�м�95�Hx���՜9�l�0��!'����2��(�n��*�,ٌ�8��H�>�d.M*�J!�;�#s��	�:՚��7�c`S�WC;l�v�"o�nA�������v�E�GS&h|JUA�wfwEÈ����� زbS,��}ǧ���>;A~Π��̂�.+��9���1��˵����m��jz5Ϲ�Dw��9�a\Z�b���nZ�{&a�ъ���P����ZE��樘8��Ӓ5��Y���<d<�a�Y�h���!�/}qw�jW؞g�u���G].jQI�C���lR�O�q쇣r�3!���=�L�VF�;�&�8���%NB����SHd-)v�}k/��XڰJPA�$�0����J�`�u�xB���OOX��>���{��pd�d����>{�2�Μ���:NI�1��r�0�ˋ��{�Nn��e�#'�vi72�%լ�v>5��sn���3����g��a���m0�KVy��QC�E�q��w�ǷPI.��X�s�ٍ����q,���+�gv[�
�SԷ	Ŗ�Zmˣ�ر���o2SW�rx.���W$i�cd�*�u}&һt��p���ܒ���-4�*�s�K�'�S�>O�`�rL,����a�� bo��f{`��S��y�b���G	��e���"z�:t�3�sg!S��yl�Y�"��v<wby
�K[�N���pg��6��Bd���t�H�yT�����{a<�H�s}�R�#�y��dx��p��2�_K1�b;�Re��#��}$��(+u����V�Y�}���H,=@ߣ���w�xa;�!#} ��~��AzcCS+:��?�#o*�Ė�ר���:�z)��A�i��#kǦ��b ��:�>� �)�y�=Q���1W��y��/0��2XJd�yj����7�ƭ��#�$L�yC �m������Ʈ��ǂI�W�,��=㦷�$닾*�
��̦�V��'��C�<aA�e{���0��	��o�lz��	��T� s�{8е~D�q�_�sߊ�^��*9���	���L*36fn�R�Ό���`�C����Q�0�R̶�u�u*7D��'F,�p#�!&$_yvS�t�c��|���%c�*�?ɽ�ו$���w(�>��"z]�^TsM�ƞ�K-u�2��ի��� �����-91w�W0;���{:-��׺�<^Tp*�%�~�*�K�z�Z8��3�Y�ת��t������A�$/���k�ICf bW��tj�ߛ������x�@ή������\�9_�Ufn��jx�'7Ўۣ�_-��m�������j%��B�-O����}ׅ�bM7͔�[=�fZ����BB!�pC#�Q����\�}Z�(`�>��O�Ϸf���Y+��lʭuꨲ�׆1��2]�G=y,��"k�7N���gG���g��+�U�c���?o����\=�Jd�cR��R���� ��A��B��G�=oM�~�Q/�0:6�S8"0��Ү�n�#=N��[�N�����k�p�.�8�+��nj���8�L����<󓽮{�U��4fp#e�YӚ�bS�*^�<9Q�B��Ed���<��Be}@�(�U�%No=��fn�:�RX�)*�؍�ǭ}Ǆ��o��!�x:A�`���ܕ4�m�Ra�����������d�`n�n����%c�!*���>5��3�ؗ��q������SO�Z�i�I��Ȥ酎U(���U��ۨ��0m{�E�u�);mp�ȥ����]��1e���RXH,h�P�~;JQ�=/µ�a��v{#]F%�B
��<�́2�7���"'��tq:5W�}�9E��\�(�	�M7b^+7��9�K��:�w_l���ӷ�Ko�Pp:��Z$V�+!F�V�n���Tr,L��;��g�޾�D�͋�����=��F�y�ո2ހ��w��ȱ3��|���FWE�*I��@`��ρ��6%:"L��t��J�/^��y�U�]�=��]�"��OF�2J:<y�J
��C�5�62�d�\I����G���Ȗ���\=��q����s6��|[��Kܺ����'k���tØO���'W�'mn�M��G�L�V���s��{������l�h�#6#��A;:�
;�	Ck��,?j��-{W�I�|���+���$�!�R��P	��F��S�hR3K���-�N����c�O�iS�v��\]��U}�[�"L��$�k��M27k;H=��- � �PŴS��"�ڲ��x�����gEo ����<1�cV{�Bs�^p�`��L�]�X���g��w����3E1�=�+r�\�r�R�8YT,>0�B�Ϗ�9U>�z��Ͷ���NBy���s~C����n2�!��7�H��<��SI�F@���4j���&:|�+ڊ�s-m�N�Ɲ��=O��p�	s�y��дg(�K�XQ1���z�����'K�	t5P`m�N7�5ӯ�����r��Rc�.�25L�y���+bYש�0�4��w?Xu9\�C��`j��;c�Ov���$�]1[G_�3~Z�6�j�ydn������K;�aN�x	�$���[Zi��D���<��K�y(���Ss��5�0�J�̷�j��prd��`��D�Oi`5l�U�j���|j��
*���E�½��e� sbT���杕�Խ1����<��S��D�V�E2�����#�y��.��.Ӑ�	ڸ�ed�T�� м�l3cLb�c]RC,0�����t�I˼��6���5���:���3�Q�m{6�F�q|��YvC4;8\�,���$e��Co��
\ڞ�ŧ�������ʨ{�Li:�J�]��nđ�@!荂9��u��˞��i��Us\��i(�4	��:�d�v�]����Y�R�Ϙ��y!��##��-�1�T��,�h�FY���jbl�ɚ�Hx�ZUe�k&Jr�1lm(�vևrj��"n�t,!�,�D= �nCi��GTbhy�[P��Z�_W<q j{=j�nCNP�y�#U�M$C�H�!ÞkV�K�L�XԴn-/!k:B5�H����.��s�P�;)8:��0�(o�TY�bVg��̟F�L�z�.ܙ=�o��O����c��^�xNH�=Y�(��I�^5�G��r��U����=O�
{SU��oV��m�u�)�E�;,�V�:/���r��h�UB�F{���|��D,�����/�楯�YB#ϕ���N�[YTfN�֭W3{hH�Y���ٓ�5t���2�g��w@�S�=�V�"=*bPf�uf�ι� >�/4�n .���%O���9�W6ѡ�hM�N�(0�&�Tn�:��!R^=��A���ʤR�˼H~�bZ�x�����'�\�~79�S���r>�C���}��V�1�Oh�/�}ҷ��� Jw�5�2\�]?Z�ծ߆��W�ه�ʋ��V�kx9���S�x3X�Juzq�1b7"��0h�}�7Q��G/���_z�;;�h�\����,"�Q��*.7m���X�-�v��K�rm�τ���������[��7��"Rk;-�&�<�������i��òA��*8浦ފ��5Va��!�勗`���T�6�Ǘ���W� ԍD"����M�+]w,M�(>ª��5Y�T֙��Fe�x��2�&��dɋBv�.�ɨ[x����7��ǗJ��|�s��*��g{��7˼7T�o����ub�x�\��v&�"����6��S���k�K��Q���>d�\4�1-�,��\��|)��"�E��Ԧm�&�s���3�ӗ���͓F����%�GD�u�D��]Qe���W�����М5dؾ3=n��.1�Q��D03�.�|�s�:� �g �=8j�Dr{q�jgCfs��Ӕ�"ǚY�4W2>K����yN��-ꌸ�����T{�b�;��z�h#]�{un4��i>1lH��<=�һ��^j/0n�WFU�z�O��=1��b�����������{����rk�Ǯ�����������jK���]Cx*7"�����Bۭ��H>F�GvT4�Zg�G��ʼ|�ɼ��o@�m<�"��\H���cCX#��1�����mJ3�!�vw`��w;uZ�]��Ⲥ9���>�e;�;Y�%T��u����1��Jw��$�"�)Y�z�pÐo���=� �4�ͨy����t�Ӧ5<��X�E���}X��	\�gM�y��w?v�ܣ�:L�үx������5�zeh�G�׊�tX=�8�%�i��<�(b����@����}ymj���Rʲus̰���V*=ͩ�*�7�4���8^.83��r��p���V�]��+wp�=,���
gr:���`֭W==�oZ<�[��N�떯Nc�R[�5��mX��9wr�#�,�򵯧�Idη��|z�=;w��9L|���d��r,E{a�/]�8t�!��{�vn^�n��gXɻ{F�>�"/Uᢱ�d�z���W��Ջ��a=�N�Lw��>˂��kI���-�e��B�)��ѡ�u[�e�}ClM��G��r�]�F.�̣`���M���#"3�9m"�"8�DH'6<<��^O���9{{�/���J�SIK@P���F���D�4$��=:t;#TP�AF����ɆAZZӭ�h�C�@SE4P44�:t�ӭv�����
�Ri��(+Jm�����:�4 ��t�ӧN�b�*����K`���[C�N��4�iH��5�]i�N�:t�]�`�1���I�M�&�5���ClAN��iM�����.�6��t�h5E%htӠ�Rh���44�Ta�jѡ�h1i֋U�ѠևE�K�hv�E:m��g��U[$(j��CBF�:���Chtt5M)0PU1h��t� -��M�T��%&���N�it�X��md�t�N����X64��G�% >ë��a��
���S�@�[@l�P���T5��׳em
ܦ�	�{wZ�Gg�(�%
E���.��s��ofe�ADJ)/ ?���{��p�V�z]I	������d\I� �-�M}��Tö���~̿B[#X�³a��-MGA������S�CPވ�kM��R�����N�=!�V�{��u�(��b�j��Ӭ����2��י��A�P!6JA#8ϛ�}�Y_.1*<�A����;~�kd�v��ڧ���z�T��!3�C���j��Y�A=�%�]8Ϡ�c�VT\9���U�����_c�̡��b��)CO,�g�FdY�/��R����y��J�0�����|������9��|L�:��-<H~,���ja����f�#�SsP~��=�)��#B���]��� �'#;�8c��+�ȟ���0�px<1��M���B��`��g�)L�=Qˮک���Ww��MWs!�4�@�Rnl�X���2r"��xp^0�	����q���cƣ�u��{��(k3_j�[�9�V=�m�u���sb�q{o�%�b������Aփ��u8�Wy~w�?��-��y�#��G�u+�%s�U���l%�y�a)���ݎ����Y �{d�xמ�w��\�x7�&��$���μ�GGv0W��F.Aó���V�_d����.&��d�)��E����Y��N��e�<�d,UsvF�}�d�%�V{H�xvZDe�5Jr��ؗs�kfd�|͗Q]����xf��s%��cq�������5"����k���QaV�y�߫�� +���+B���k˹8hӰ��D����ĸz�pXt�8���2`sm�hZO
ރwx�J/~����Ts6�1lvB�f��(�ggjY[�w�@��\-��8^�.`���N��X�T��5���%��bi�^�#`�F�,�x�s��@�g��1��&4?�a7��~*Y�u}���'��oQW�'��t���Q���݈F �Gdc�+T�O��&��X��a�H�W��6ꕥ��[J�-i�a����wH$=� �}�F`����s���c�0!�">e�E���uO�U��Hw`����ߪ���^���{ �t�43��.>�zu���Dk�h�[����:���tÃf����/bj1��*�_r���a�RˡF�Ty��^5��a�=8�*���;}L>1P��,�?�m��i�8�v�gӍA,��n!�FȔ��e=��l��l�1YW��oM��!��w$R�t��V��Ol��؜Q�0g�6ئZ�Y�	C��؃�8�{�v�/��FG�b�R��f�xmw-R�(޺*��oc��F5
�y��:_c��y�D1z�p{�^�h�S�u��Ý�_i��j�ܗ�.d�$3Bӛ�d��3���J�W����a_^>���[���;`}�}��0f�� EyT�^����1��RX&PT��ټz��	�����R���!.��e8X&�4۞]���.؊��	�)� ^%�.�y=-ݶ+�)N!�U�E�05�m�a,ʢ"�H��[��C	��t���"M�>�I�9\��b�P�������;��~���QUӘ�/NKe�!�k!C!���t� ���9}�w�iC�TqWL��1���t�lt>��a���$g��jxI%�{"���2��)�
x�nr�0��H����#b��-���w�Uz�C�W�m�Rh��(L�*m<)A_�B[��c��Wb��M������$+��a��ϧe�Mֺ���nռ��Kܽ�Q�&�Y��;!t� ���)����FN��1��1U�qo�k���:-�d�c~OO���h�����	�^�Ga��85�B/П
��vĵ��Y���ލ;/T��n�mۂo)��L����nD0͊i���ۣg�4���Ҳ��R~�c��@�}��e�^��$�c#v�����C��D�MCH/��ՙ{�Y�m�z�U����Vux��0����}��GC�m��xl��<J�z��a��c=��'#W�N�!�l���c�U�/2���X6ay*�`�T�l�ʅ��L4,�wt�4�S,��+pec���ο]���:���]ຜ��=�a�<��`��tۥ�I���[���U�e�Ώ>�uG�Lcוndn��L�]�X�B$^�=�\�m�Eo<�8M�$ղ�U�ZfP��>��Ub��U�Q��o׫ϓr����^4��J����N�z͛O�4����zG�X�+���6]����>�W$�v��V��:�c��ɭ��-���#v3�V�o���t��z�A��BD��M�r}w��[�^	_t�(Fu ^��$'9D�O~H�2�=�ƒ�T|1Q\�U%�%��>��	�ո��X�5{bqٺ��Xt�	Od�z�%:O��Juk�S$�����l��K�z&2ש��Mu�W�u�vL�	rh�#,�^ڞ��'%C��I9w��&9z�^��W�=s�����/X��!y�\�~�-������k���F`�?�E���iwO�eڬ	
�U�x0��]��:�M0�#�":�$kr�N�b��{�P�r�֗!��Q��Q���	�#�cb����k(R7�1q�C��.��(�n� ���G��/94pI�e!m��c����"{�㮃�Mz��/��`2�뛙�ά�m^��lսn{H�j��6�>y;N��CJ����{��〉��=�u����gf�c���¥�C���U�0Y�/IB:C_�Ho
)��Vc�}-:�՟��ŴKi�����۸N��o�����kn�5X�g�r�Cݱ��9���b���&��(��\�����CslΜ�aס�_Kׁ�b�]���Q)�}e��zAge��WA46Hts����k2َF�o������aPO�&05��U���k8Ў����a9�a^����1t˅��o?wf;�����b�Ԩ$y9N0>h��X�6�D��w:Dh&h�U'��d�7��\�"����wn��R1E'���A˰�O�:�]���m�$ψ�:�|���'�ƒ'�S4!�w��y<����5+5ɤQI�n�����4��,+v~�C��	���R�aJ�"����8M�/n�y�X`��rb���A�J3���8��[B}/N�0d��gɾ9���Tx/ytf�b�u>&�a^ڊ��wB	���	����亵���V��ZgP�/�?'�%if���L��)��hs��+�hN�~4B�nu��c�yN��J�*�
c4�D�>Zl�
�ٽ�eeq�]EÚ��3�\[93�܌W���G2���*؉N�g!���ڱq�����Y[��Z�o�k���D�u���tGt:i�b��;��ᾐ�n��%�t�ziŒ�4�qu�QKݴ�1�Q��}-�����J���)V��|x�+d���&�;�k�n�0����f�z�RĚ�~����F�sׁ���By��Q3�E�[#Ŝ@��0w l���Y�i�a���v��W�P"㖶�'�̕�Ȥ�q�H��/A�F;�	�  �cL9	��T���x�"��:�ˎأ6��\�-HrU>*Jz��ڻ�u�vcr'��b�@�.�!k���c�vdЛ�z�ʫ�G7uE(6��Q��D��̮xj���I�,y�a)�ݚ;!��EZ}p�p �N���0)N��[ k.z�\��h�p���IaKcX��XN��,?5�c���;u�J�ם�r-c�^��?1�0t�� �c^�ʹq�k��^�.��/k`��J�\�f�-��	�t��R#L�T��1.�-�Å�[72̶����:��|�DX��(9�����H��z`��+T��l�	@�`<h�Þ#��&�tmt�Ɋ���כ�í��6�F������z�3���P�,��j�1��~yR��%4&fH8srk��Ւ��"�������wH$9NmD�1��� �xcZ�9�ƒG"=��3����-���uL�<웭������n�(O2QH^��>��e]����O���TOS6��F:�#M�V
�l���W�;0�-��JȎ�&�a�:�4�L��=~�cj���k]� ����/��9�!�c/?��P�ҖAC,A���|#d�����כBq�����s�K$!A^iN��D��DGM\(%�q
�VD�+��Aw ��5y�_�r�3-��@Z��e^.���L�����7�m����{/�5,k���?�x����a�籞;����|��T!��{#F��\�[J�+��vP����y�i9��E�F9���+%��Dê5��`�D��v�^����<��S<'\RX&�%P�ث}l���֓�$�����/F��I+]E=��ޥ|4k�3�8k���I�g�2N�7E2����_8���P�����T���R�37؟�Ykb�}�X� u�5:�\��5'��n�cY�6z9��՘��˅�px�fq�A�����li�stt�AۡF��P�⮗������Ƅ���k�鷜�H6(��@k�w�w��&y �������WP��#Lv*���S1�{�{��m͋X�~�S�xJ[��R�zB�de����o�dΚ=�n�g���{����ےP}��6y�L�[W�q�Ņ'��<�
���=G�Ns;WxXV��ƴ��W2���/���{���Ԏ�}w��K'S�n�a�G�t���Y�����u�+�	��n�uazM�
\:eA6P�4/z���U��M| �wW���[�q�jS��9/R�R�0z����]�A��(<yO�I�mTm�h�=��_w!q�����;C�䫦͆�S��v�	�נSᚽ��z�r��lg���Eм�9�0er�S�{X�V�6�b=@�"�;<c��9��e�����wUljp��)/p�xVh�Į ç*˞$o����:�Fȏ�Q�k�Kw3���Ͼ��2G��y"�6���=���Hh�����o��ǖ����*�݉[Î�Y�U�HاR6YŎ���rhL��z������(]�]�?�f�2����zE��HZs�#6��ө��=�vj��Ⱦ������Ύɬˍ��{�� H[�D�ڠ{2@��3V�V���@�|�⍾�^���-;�^��m@��)J�3������Y�3��VQ��i�)��������\��)�v���	�I�+�H��yz�{r�s�P{�Ǒ�}�x$��Cr��!�"<|�.�C�˻v�:�F,�^:�@Ft�_gm�|�"_����}��e�B�<n�(�x;"�����0��y��:,���MaĲ�׶��*�A!��C��,�j��w[c)�6ܷ`��^����K%�ǶxRD� ��2�����p��Vh:r�x��I_��k�ge��3-���&�Pk<Y�r���Q8d6c��NG�����������GI����J�=��}�Q��Gd��䟽ع��"y�<��y��F�+�=��c�fF���U��"�&��^���Ȣ�E��c�{�Z?�ϣ۸ ��?�H�]*�d��FUU{ǒ�]��*H��a��Ɏ�f�������!��8���l�&
�ڳG���'hoTMl鶧*��˭\�����$#[���Ⱦ/�q��*�;��;K��a �v�/ś*8֊���t3��|��Ñ����:_<;I�RݹB��q��,�C;3vP�nH$Z<tQ�:)�;X��
»�j6��NnC��jm�e߫0�+]���O��-�] �ȉ�g�b<��-!5�M������s�ɬ����r`��Ĭ����l������	�z�d��Ȱ(z���(�[� �-t:�k`�W?��t��m�+70]k������+�`�b0ltL�Ö2��Y�sM[O/�w+B�&2Lli�W>Z�wf���g1����˓2/n2tV*�U�3�'
@�8����!.��yjE�}
�X���OC2sX�NL��&4f���3�<��V�%^Ɋ�ą���	�B]�'���k�����bȳ�K����x!dw1 -�МR:��,�P%(]��r+�Zb�v_q�;������N��mrr+$+G��5�K6t�*�^OB�u�˂8��2�+n��̉c`Hf���p{�iQ-��W��Y+g��ӟq���"��.=O���s�h!��.��ݸʎ�ӗL��i�����Jhi��r���A�����9��f��y�*�6u��hX[Fb�$����UY\��F��wO�c��,�ۼ�f��y��-�!��:\hGO*j��^�H�]�*V�v^���r"jEe��b�gj2�Lp�a�q#^�=՚iS�7UΫ��6n4I0�6������\���^4���v7pu����M��X������$�L�����v���� jI�f�8.ײl>�^h�^7��&��
�s�oQ�mǬsxy!s<c�����|:�ԋb֮Z��c(�����O�T�{/������/�t��h�[Z���_E����uϳ��U��ު��z�.�x����aW���3.�wi\�{Ө������H��y�j���[�f� ��	K���L�%7$��׏�^ї�Ɠ�I�C3�V� �+xu��*��_���EmA�s;އ�wo�� ����RP�Z���|�4%�z�o��=2v���)mܭ��nlQ�,X���N\E%{z�i_q���Jh�F�j�C��Cj��Uҹ�ʇ�Y�ʃ��	�+���ޭ�i2ޒ�"ݧ��坣/{�q����u���!=�XB�<2��.s0�����*h�4%9��|O{8*�གྷs��Ӹ�	T	�3�P�	���.�+"M{׼�-�6r�t�E���]Ӥ&+âY��:��&��`a��[,]>M������9};H��j�+.�'�է�dX�b��p��tl�r���x�x��IIyqY��wn�qK�N�&5��������y���~(�7�S)ԫ��܆��Z,�疴ѳ�l�\N��)�Fg9�ܩ)t�8m��*��$��Fc�xM�5%C:����i���,������nB�{Wu�`^�S�$���%�I5'gH��\+)_Ou�b�#ͷ��f����P��v�z��m*�n\�A3{�O�.f�l(��"�1�$�|�-�7)���od~ ����<짃���x�|Np���]��L�Ժ_�X�TV&�kX��w:���t��>�t�;�Uc��/�[��s�8�e��4=��)U�0>n �C�U�����뜏g�4�������|�`�n�`���;��0��$��5�F��Z9��r�>����V��d�O]�p�;�J�Mt�x��7��Y
M�t�s��ť�5�W�RO��O�oOi�4��_M���}����h�
�Y�Y���Qz��to>���^^��Yq����C�X�σ�w�\�^F��l�;�\/�L�)�}��5���Z�:6�"o��"x�Åw[qjf8�1�l���%?zCy_t��>�o��{f�*���X�>-b�#�n�6��i�<��<'����]]�sU;sHν/�2��牫sz�o)GR�A��c�۬v��>���2]�3��B��N�Z3t���klD%��g������q���_{"��Н�ȵf�]�_����R�5gUV�h;p⭍M����`8T�Cz����Μ�]gJ�*X�2vŽ�!��q���V�����.��9ي�|NU��L;=�b�) '^;6�\��)e���
��B�O������`��ڀ����CJi�C'�ӧJ��P4"��RAV�F�:]�.��+BĔ�jt��=:t��&ٶm����m�ZF�4h4:MB�b��&�:�ͰGN�:t�v��V%��bh��-��ДEKZWQ�&��h6�E-�ӧN���4��N	��̚h5LTV��#m��UP5A��i&fj((�"����4R^gTj�]V�l��-g[mPi���bڈ��
K��Ѥ�i�4��I���b�gE֘�C��5AX��Ql��-�kh���h4[EI�ti����Va�Z��Q��֩��PP�l�&���1i(�X�8�"��I��BV�!X�.��]��
�·�dtSAQV�1%�A �Q�R{+��;o=K�-g{!�'ܦ�������O�c�;��Oz���p��Ů��E,��.�s��[��:N�0�~����i^�_����Nt{�F�Pn����o0�ld��/I�9��:��KL��yS:�������1�r��2w�dv�4�%�G�0#|Ĭ0.6��֋��դ;Ƈ�7��v_*�2D�c��a�v
�4�6�᳚"�����)O_v���Fo4���C��$O�HJ%��tS�����n��;�y"����<�j�"o�5�ݢ����$�&�l:1M�sC+��^���藕��5�jƩ�<�{�1kQ[e�-44��Q���w����NI��֟fґsNge� ��&c���F,!5FG���>�������}�J������;W��ȫg��FP����ە��&��rEM�Ҏ���/��$%C��O%AIUA��F庑V�:�L�8���Aە�oy����%�G[h�m��)"Β���o����k�H��~�}�g�Z}�eC�-s�����N+);���vS���Gf\A �������m�3���W�nvl��evm2Ő�E�M����FU@��������b�˹���{�{�C\+c��=}G]��M�T������mӶ6�h ��{*6쑘�"���Q�y� m>��ܩP(t���&�<Tð��ʩ�x4��d�aN<������rh�y�mlQ��FY�ݜ��(}���kPs��]}}�_�/�����S���9S9�3�������<�ݐA��lEn�6�|i��o�XVw��-R�w�ʜ�Q��矨� �˨MEJި�����N���cژn�7��0<%�52t�=E�r���:N�2�-m���w�SF��[oF��D�n�<e���#16ϻ	��H��7�t���d��LڭW�����&�=�X;��>*B��F�`��̲�x�<X�M�����j�"/�AP�ӂ��"��V��C��l<���i.�vg<��E+��s\:#�kR�p�(�f���.we��D��ML��������2��'v�f^{�/.�Ռ���ݏ��/�I�:7��ȕ�=Inp�e`Kf�{����f�n�3:�QH�H���˛��*:��s�p%4�S*o40�R��8����۠H};l�����e�3�*bw=sl�n^�DX��>�c+&i��J�-U��ۊR�݄7iQGPz޺�sN�l�������0Ut��d^D���Vխ殥)�]Y1�܂�ₚ]&��G�$\ә���s�J�=��ѽ�m��l}9b���D-ݪ^��m@��)P	N�3���mDA��ŝV�ci��z��x��o߲�|��T��^�$v.�ܒ�tt�ulL�ml�
�����i����ėˍ�~��� �d�g��r�;4�L�QV*��r�����F�d���g��ɒ覟wj�'�{�n
�\��U1�:{ է����יm��c2;���͕H�۶���}�*{����`9�Xz6��ln���y�u�1W��k��rJ8�����}��1�i��gu>�~��%JC��<}7�h�f'*���Kt�zJ�R2@�`M����i�n��GC�������8+����=ު A<!�&���/���I�ؼtv*�y5/�u���tn���:�\����dj������C_u���+p�v;��e)KqBH!d�^�1ҡr�h�y�L�5���Nz���]m1v�\jܡ����{l��v�7ml���B�mj��Bl��`Y�q+i��[�$�).X�S�V��$�t��g�����~�vݾ;>8�W���gA�$�W�iyVk�ǃ߽�f�d�b���CÐb�rC�wuf����RՓkc4�=�@�1�w�����tQ�u �F�H/8/�0������l�u
٬�ҏ^�fzڛ���fZ#��a �4�X嶫���,L����E^Z}�Fo_7k�t�{hL��^,�1$	�
TA:e)��u"6Y@�<w0hS���Y|a��`�i�Q{}����8�ڟ*�]����Oe{�&�]���\!��y5���d'�e߂�GDb��hW�����i͜�M���!晋�o{�C�&���A�	�6֬x�f��	�5í�n�'�T�Rq��Y�n�vd���H\쐞߭�-��j3���+
HH�w_{�?�+�%�Cel��s>� G������o�|���:3>|.�>�I�^�+l�E���7�L���7_9ԏv����N]6�D��]�k��Q1N����6����^{T�Ġ��3�?f�SA&)���t]SЭ���!�푄po�[{Ô@:�^�����K�C�[γr��6ڬ�Ҟ�n�L�g���N(&ӑ�)P�+�������6�=�ێ�����@���mo~#$+2���׎]���J�ַ�}F��� �:]=�k�!���d��3+�V��5����B\n:m��9�[ˑ��5o3�<]�Xm��78��du0nHq !�5�������j�P��*�OP� �zL��l11�́�p��y���m��2N=������{������]� �G>��sk����EOӖ/T�s�v4l1��wl��1�ت��m�K�����9� ����'�%�v
���s=��&��R�m<��:�haeC�үd�.���3,���D���K��U"kh������t���w3K���Ɓ��"�y�)f���r3	�wB6A��y������{���F�&B����{a�wQ���Q1կKQL�jDn���>b�a������ܧқzc~!�7���X�'{����X� ,7Q���Hc�\�v�\|�����(^���@-��\V�5'5��ɘ�3��K�ͼW&�D��Ͳ-7�)�ݖ/*���n�,��o���KQ�1ί��s�ΎB=]�����W�jR�T����$���~����Y��Þ��]��xZ2�)듵s�sV�7%ce)��ݚ�Zg.����N"�oHnAH���))�Tm�i��(������<��lLqn�#�_���5���h=��mq#�RV<�Tɒx����t �E���7m���}���g)�;�k�8�O�ur�RҞkM`���p�r�)����n���ur�Sl0��,�Fj�ꃧ�[K6�f�h������|68tNJX�\_�f�H�i��Z�7�^�����l~!�9���엜�ۢ0����v�6�!�HB�WƼ�C�=%��ݢ��a�����ȸ��;#��K{�0&��8�y)�=�o�Ʊ⭭�d�h�蝳�2�uH���R�y���<c�H;�6�蘥[y7�6p���N�)}�'&�M�z�i\P�S�p�讬PԴ\�w����Y��mVۯy��{��*ʶ�sЁ|;	�	��=���}B�@�^<�vu˺��보m��S������ua$��(�����UZߥ�i�:$�:���p�#�Y�/��sA���ұ)�����e�7l����.+���1mtg��C��C�+��q��Y�¨;|9@х�Y��J�����<O�5�[>K�/T���GY^�y<�_O��}1��H!\ܒ��x⍎٦TʲC�^�>���=���%@���i���.��-`���R2ʹ�M�]1���y��3V���(oZ<m.
\��Y>��:��p(X�׎5��*�2��[ٝ������1�����aJ���d��s3p�<�>����2��'�d8�8![��ƪ���T9JIN���ߢ����H1�\E�őJ��[@R=΅H�S	� v.��s�4�KSU���x6�x���l-�1Y�~�t�t�"�:B<��H�h�=���&'_��^��e���f�M�2:����|1�E�\9dl���7B�a��Y�s����o{���3��YW1͙/�� ��5nf͗��f��]���]�Ի��{\�X���Gܕ4J��~
���7NlŒ�"�Z�3`N�:`|�|v��]�F���A��x�GsqhpŞT�3_S*c�K�鄰;�]�^�.o[��x�|���YQ&�xh��ei-�,�d�����՞AcBjjy�t�\�\끺kn��E8���M5=C�B��rב\�y�������54l�GfC�t������g'�+�χf6t׺U����ԷLP��T�,�lSTc�;�T�����a]0"<�Ƣ[����N��=��mT����_9����߶�xOC(��Q	m���0A�9�;n�|vN#ݻL=D�z/����Tqf�ys.��:|v��1���g���䖒���љ���kH�YZZ߆6��M@&4f�M@�������F�x���ˤ��0��ܣ}m�S�ً@̲F�Y���������O8GZ?Ro�;Xb^h���\2�Q�����]P�Y>5�JД�Ee*i�!�q����x�fR�ޟ{4?J��

�6�#�̾TEnVLT�Imvdڔ�u�[<�2j3lK������1a(�S��nE�{ڗ�\K�ߴ{�2=-5O�L�8{ ��Hv��O�����&��=����{A�'{7Ѫ�Dƹo�ǧm5+ɻ������ћ3�s�V��G�)�D׽��{��u��xN�U+����lk.D��� ����������B�Y�q��npd���>rw�T�z�GM<� y9D$"��JǊ�l�H��Y[̎j�xJ�H������ܷRfG�,�����]�K���˳7T�S�k�7��}#v	=��\е.2�[!��ϳ)�Ka��
���]���y#��7Tb�q>��Zaq-�O�sl���ܖ���lW��TU�lvgt�r�h.�C��q9S�;����Q�����L:gXɋ�x��|
��Dw�Ay�X��;5[��3F|s��yr�T3�2�<��%��"�lwL7�Jt:�8������5�%ӓڳ��F(������ON���\'�o�0��bWG����Sto�h�pF�y�)6V�5򛇩,�ǚ=��x-H���#z6F�Ӝ*���7��|�^Ж/a'�IY�O�PҮGdL5ރ����DX��&��_t���uAi��u���ծx�t`d��C=�Ye�^�����׫90K[���JqcU�`���B�[%��܆A8�h����Hh��VNԴ;���G7��W����Z� �{E�{5�E��!3��d�f���1�L�>X�;��r����iM�o,g�#��q#��1���үd�#c�ve��<	I	D�C�s�-|�2)��h�}���ưfq�n)�jg���zJF�]u�Kޠjw�_���k/9��}��M�i��=��>���3%>|�T?8�?V;N�%uy���~������4�(+�W[`���s{,�S�F�����u'��۝�/6�3�p9��%h�Q�|��K��g@ج��b�b����p�od��B0�������S�P��T2J�~yC��M�R��c���5��f��y�X�B���!����"6��t��:]�d�*�q)��-�o�$��jVG�B��e��79����=`O�x��"�h���F�P��w�N�g܂o�{��2m�� �,��]^ι5����4&��m6&�hA魫}~�/�'�|)-wϴ��ZN@�<���:�ⷠ�o��avi�38m=[�`����=�Zި��r�h��m�C�9I1�K���\)�q��t9���m��I��	��猿#\�_�� ��i�ߺ�� u�����o�g�_�wEf�He3MĲ�����!��\�)�k>�ȕ����W���t#����&�>��t�-WwU�bƾ3�� �M��!H���X��͊WR��B��z��F ����K��tqA��<	�\��A�AP�j��dp��=n[�{)w<�F��iH����*
tq�U�7�x�Po2n�dsk:�;��!v`&:@�·�#�JD���2e����S	�a��:-���
8uQA�W	C�ٓ3�cy�Yߙ̮�i.��%�bN�����|76U �����A:D'D�3F^�G��Orn�5�����e,C�v���6��5����]e�0OY,��$�nLq�7#�J��j;�ٹ&N��Li�N��7C�7t������rq����Q�sZ��!��5Y�;�w�lk�3�}�tN+ULJ��.;4_-��.gR���c��j(��2cC�pc����w8:���\��S.�a>��V�1֖%w"tqA̓{�72��3t�DY��]#c+�U�{�s��P���s���^w��������x�5_S  ռ�ol�^���^)􂠻��a;�^��AlCr�#Ya@�\���qn?�����U�	��*�8f�s��C�#kF����;��ٙ�O
�S4�*��n��e%_�H�@p�\ԥ>��H��P5'j��[�
��Ȗm�n�MޜἆöJܓ��$��-�[�u�&�Yy���{P�M����x0-�hW�Ś��E�%�ǻ�1�S����s�t� �hj(�5�{O�6�Ō��u1WZ]�Kc�a@�t	�^�9YzM)�<�������@p��}���$����Fy�s�Png<Z�9����KI�	�q�c��rmq.�w��3U�f�v7����5n@&^f.ͅ�{��L|��<��RV�=�����%��mda�֎�ʛ��4h�j�>Ӂ��ged�ś�N�J���-��$}Ѩ��8 Cg2���9s=��=���jM���;f������+H�Ζ�96n>m#a,t��,����}4���s=�/6C�)-��g���9�Z�6�]1�<{���	e6oHA�KB��6nq�5��m�6�{[X�F�Jk�q��@�B�SK$��+�0c�p�ՅFG=xf��'��s�q�Zǜ�:
.f�'�Ə�;םP��c\�aB���(������I��h_"x3!:5Q�+J�4���=�����̽��W8a��<���o��v�q���f��h	��8Nʻ�#Xikf+�x��^��!��b�:��e_mN�A��wdՌb��` ���16�h8~��,��B�a~IC E�!J~��z�y��9%���}�ƚ
���lE;�e���*�*��UU�����
���1[�{s����ULl`�N�5g5Z�kE�[:fM�RV�b5���_�:t�b�v(��3F6��ڴ�l%�EF�UD��M�������kE�P鎝:t���:�a��J)�F�[4DD��I��TE�lh* )���I��t�ӧN�S��.�馊4g��5�E!V��0MRQ@QLDELS[Rh���TPU&ڵlM������PA@����kTP�εm����mX�1DTX�Z����5�b*
-�EQAC�4�ґ4��gQ5�IE���ӊ6�4DP�Q�N��l*�""�Z��c��h��&���4�SCU$�LVɚ�d�UE;���A�"٧$LTM6ƙ�6v�5��h�b���ƵTZ�FƂI$�;9{���>�D�[%������x�}6	i'e���
�b������մW�g���E�-�s�6�_��T�慨X�)�D�%�廣�jh�A���uiV
&W�ԍ<w7C�������a7��)���V�,��H���'wM���@�g��ø�'��ܺ-��G�`�z�~��*�X����GGZ<���&���#)>�a����߀U2�G�iG
�q�N��C�T�&��W���>;B�
�l���=l��Yu����D�q�[D��͈�Y;����M~�ŎK2{�i
E@�a�5��
�];A��]�����<:����޺.�-1��v�.b��gB���[���)H�qհ�B��%*�M����*�w5ͣ��0�;a��4�A,B}�E�®��S��k����8fr�xB�߽�پ5��e4��f��O�PXg(q�'��6� Q�͕��l��p��Uo�:7��
UP�s������qh6
��AV.˯̋��������=._o�Z7ġ������o�Çvu�,���i_A��(��g-��3�h�z���{e�9���Up8x�sUA����n��b~��xh�:��۫ʣ�8���=ר�'$�7+���^���Q+R�J�J�g`}����od`a��P�s�.�!�l��
�R���k��ª��V�����;�8F<�V]��n���@N�ABS|,t�Ԏ������F_Ku�Ǚ<ےG]@$UW���]p�.$H�H60පr�W8�=�=s1�}�PFF۝3�ls�4�&@'WQ8g͘����-�r�X��SO�\��\q3O�(��2:��m����K���Zٝ����<�ȬbZA��`1��]8�s�_ъ}OWMOWb��^ErJ(����@a!�f��]eAl�z�)�YH�A�l ��6ut:�Ҕ���.�Uw��ҩ��l�~]}f{Q�v�h
�` �pߡ0��8�i�o�~���up����A×69J�==�7�7_y��pF��]v�砈��U3I�jq��5p���ҫ���:A�=!��6�l
�:�Sӫ5՗V����+��ͧ7��N�%`���A��0�=���eD��%b3yA*ϓтe�'a�/�?&�q� ������A���m�(����3��K��Y��j�ҲM���"1�/P�q��yN�6�}����o_c��ړ�8g�H�����~�K4��z8H�n$�â����43D xDX�� ͡�o�C���t���;uve��;�
" �� r�U�nw���\��Ҧ�le��@�J�	�`ח�W���8��%hO��5�%C� [�ǭ�#��t+�ɷ2K?����S6��T\�%�;=S/ks[���mgu��B٣���
�s adб������1 ������n����8e�i�}$Ʃӷ��O4�Р��K���t�Q��m�/�qi�@�$�:)YxI$��U��S�n�_6X�
Of��q��Nv����9/+�
�0u�݄M�t���).:+d5S�QmK
a�4����n>�JK�k�s�3*��U��R�2��m��xb��M�fn.��c�������	~
��tLr'&;�)"��
4��z�vބ��֓��n��!�ܳ��/�ܻk�M���%����6z���)}-�i��)��=�׷m��F�zw	� ���g3�,���ӫ�v�:��\<�L4��Sl�ĺ����IQ���lEu�:�e3r$�)I�>�\2�ڍ�A�}���t*-����{[�l�Fh�������;�V�s'��q/-<����
�g����F���vd���"!ծ��U�n���l�pv��c1l^�c�#���7�~���36�?��s8#{B�-ͻ��\�X�v���n܍x�E7E�{��6@�8k����+�]�-h�E��wz$c1C��C�#�&�v?&H�,p���W�&��v��&3���9B��h.��ɼF��fY|�$H)!�w��&�����[�D���6��10����lO��{�;�=�j�˦Inx,�Q�A ���M7�)WE��qC�J<�r^���ҝ��fqq��s�fe�'y{�)�vJ�l�/)H��3�΅=E�LKF�m2L��KV�#/N���A^o$�ѕJz���*íVŭlt�e
�,����C΃w�M��hyh"�b�G=u�T.�����:`oR�J�nN�+����aq;rb�BWJ=8�⇂���NY�l4�;�+�[m�<6��9�f�ק���`��r����K�n�y��o���xo�6�<�����B��3�:�]��P��]c�ڈ(u�P��y*RU6������n�V�L5#�-ۼ����?U3�
�r��b3o���I_��T�3�9�x�4����'��><$o�l���pE@tS������O�V����)�L��d'n�yʥ�3������&��aN��Ɍ�.Ψ*/K�Ù�Z�Ƿ0�^�ُ���{0Mq�����j2����a}��62�Yn��Ն�����94��j�F'԰��wd\~���W�c���[��ȵɿ�&?V���7L�3�tʟ��@�]EQBS����O���n������l\]q�o8�����#dnnt��χ+��v�y>�<�_�}�TϚ���]��!����-Xx#��W���2���Gb=E�Mvfʌ�̎��vE�����0O.��5؎����7�ѡ[��#3���v־�=/ǃ���lu�)��ܓ]����A��;G^Gy+Z�+���\(�h�'d�ǫx����[=:�R|,���R���G1Һ8�L�[$��/��$�5���J�,^������p�����V-�q�h�S-�����'@b�'�X���Fv*�v;Z�]?$��)��*�e7��G�f{ۛ��绢syK堾�yj@��!B�9�����&+�}�/��R)U{�!�ht���Ei��R.�l��ڻ�[s��^��9���g�p�9��"�k&6{�[�Ԡ�;iLK�=Y�j���i���+s���SZ���+�$췦��/j�6�h��ؙ Aٝ۹��մ���.aZ���b�oMV*6e���f��dI_d ��%O%�[iuө���
�ܶvh�,|���E��5���®%�&JW�θכd�:��'��}��C*,t?y�Guq'/;uL��B����e��R����t\�'g�w7f3�LMM
��;�ʯx`��H���f�UxGI4f���g��xE�J
�Av=�`<f��A�=_B�o���Ù'(\�z�+����k�of���vm����ɪ�ݞ�z������T��x*`�;C�4���� -���@��aYcj�v�{8��|)����K���ֳ,��	�e]���X51�; ��>�[Κ��˩��������U��)����.g��6uVI�^0r��R�Y�5��FLCt�3l�H��"nR�Ӵ��̆j�$dt�N�@�V8sW'�ng\ն�Lrf�͐N򺅝 �Pm��0?G��|����~�k�!l�k�i��u�z;[��<x���Lvx�I�2:��Ch�`I�*J�C2ic�,.�ͷ�{[���r�A���y�q�Ih�n
�ð�}f�ɩ��+f��l��AZ#n0��Z;��,��$o�"�h���iu�n��»�u޾%�,�B��	�U]�"&�Z���H8��%h6+x���P0�sq��O¶��8��CX8�ꧨL������$;,����"����K5�	�D�����Z
�9�@���p�=0��3����VCu��M�3������Ǧ��=PE�Y�TrOI߫ӧ`Yn��BM1���r���H�f�ĮԜy�p�'[��kb�k/�;i��n�2\��>>���ųP�H��җ�
������^��CM�(v�A�yY}6|g��EUǣ�HJ.����C����f��6��޽G]����5sh V�{���V^I.1ƛ%mӮ쬷��5)���%����n����]����
zH��#��'}ΒW�).:�[�2;;�lcVx��܅:�1���#����gS�`rQ��\F�-��8���ϛ��U�H�v�}=��\���y�F|r���W<��Ȝ�i��9���r6'$��3�w�O�0~��a��dս^���������f����۔N�V�w�I�g��E�Q]��e��#{�G�R��qK=[�������oAB��m=ԬJ�`��y�@�|(p��~?R��{L��'s�E�7#`e�j\u"�M��>΍�4t�b���W�ywp67+���U8q,}��:���������&H�qc�	�Pf�+�@��L�]���vf�Y
���\(b��V����e�w z��er��O��)qa8r�2M�cݶ�7\N���֊���7��b�bΆ{úzu�l�!jێ`�����'���.���Ȣŵ/�*>�!��g�e�f���[���̭�am��cNY.Ӌ%t��U�������u݋�!n��O����ֿ���N#A����$��N�e�r$-�}^_�Lj���:�Җ�]t�ܸ��Fv��k�ݡ�pȾ8C
$�����Oa��t ���}���e���#W��<+wp����o�!]v4��R.i�쳡S�;t��_2$�w��F�xs=���/����TLGj(rF�A�=r��ji�.�Ui�5ݻ-�݊�$����U�%�A��܂��� ��%Q�i�ݵ�tsE�`��D�w�>�n�j�$2CBS��G�����IYxJY��Dv]a�F����U��N�q��R���ݞN2�i�6 ��lm�~����H�ؐ��X%HY�#��C�)����>o�w��`�L)��]���%��;6A���Nj����	�`����L���C奷s��6�V�M����k��Pœ=ˢENN���k�a���<�?x\s�wq�I�j,�N��AAP�8l���]�\�YZ뭱�����)��fu-1a���>��.��3������ a�Cʍ�vk"+C�]��Zax9x���͋��W�=2s>{�\����������r�ɑ��&x���_,Z%F��CU���[3;Zo�T���^<�P(���EsX<o�;os�O��=��T�W�O�C��y�##dnN�R�al�ピ7����.t6x�.�#������2;ղ2mjg;̂4���w(��Kl�"ⶲ�ms����nY(,c��:@:(􆡮��;�#a���b'�2�n#k wa�m��ev�@�D�b{��`�#b����+�����K�O�^g]�q�gVM�W�t��[�X�"�W=jנ�@��b3�5M��?a�|fqv}�]���(Y{/RCGZ#��G���~O#���=޸IRڒ���1��vj�X%bY��,C�
iA�+��!���=�6e��c�Ww�:!�`U#�D�T��l��
���*�C�9���~��$���O36�=	��-}K�h��P��%�ޫ45����u���\����ˍM�c��(�t���Xe�����]_@�4mk�c���}�����ؽxMm���8����ǥ�����պ��S��=�s��B���G�9�U�-(8R�L��:���Z$	�9Mh�u�<�SCV5;���Վ: G��qZ`�Gv��-�5q�X��;��זI�)Ωv��:֚Ȭ�2m)J��hՙ\J ����6�vAm��V���s�8�Ἡ�o�c����[�X]&bz1�}Ǹ(��}�PG!�c��P�E�w��ee%WxȜ�EɄݽ����z Y; ����q��G3}�<m�uAc�X����U\��dY�&n�6G,��Z�\��gZ�웒Z�v$�ɩ���M�^¸J�������^�Xz��v�r���Ojs��oe��7��+���ؙ�}Q��)�[��o�7R.�Q���
;J��BX�����VI����,���d'��9&�R)�ʑ�SvX����a�A��'�币�E.� ���y�t���Fv5x�E��+�M��9�$[�/�-)L�y�j��;-^�EM]��b��K���M<�(���!W�2�J�c�tkc���
�P�<�4\-��c_���Mtt��	��7oiA��!qN��|���G�u1jB/z�R�Np:���L��/�vN��ΞL�Ldw�>�W�A���5v�"�phgY�ʇ�Y��fmr����d��k�WH>X�u�"���������Kօ�l�;a�7�iRWi'kDob�lӁ�;�}�
P.�}H�q�ኙZd�A(9�g�����*=޳�6ϥ*�۷�O]�&�� Jv�k
��|��xj�cM.��oz�.�S�������u��c6*�z/��)g}�Eۄ�����=U�Кz��bX�WV��!�D��(J�*�頥���ꘜ,<5	5�E����;�/{p���:�fV��/�4�v&���:��>�o��Ԝ�R���t������C�=2Ët�|VL�7����t^��*v1�J*���r�Cd�WQ�A�3yf|�����F!��zYz���1t�[�M;��mGej��׷��i���e�֌4lj]�$��ٕ���{R�g*vr��^���ڦ��h���� �kV�m�rR�%3c�wκ����4����K��j���o�0U��X�zO+I���M��;�CJ�J�c)�X����Y�oZ7�=ܔ:�u*�,�nP='"O��v҆d�/�9bT�p9N��ʙ3479n���u�Y��ͧ ��ꡉ�㡍�r�i������[Ѵ®���f���<=&=�N�X�'`�͚�w�]]��QGE�}'G�2ht#<�-V̲�'c]�׳)oT�Y/&t��VJ�\�`�9o���5g7A^a�RK�8�v�Y��P8�{u/w��"�e����O�$��KL>��A�\�U���mK��d�2��� $�$$QRQZ�SLlj֖`"*�k4�;=ϣ��ڈ�&v5Z��Em�)uX��MQmyf�*(�Z)
Lxt�ӧ�����mZ�6�-�RV��h*�*�ld���Z�EQh�\ն&�t�ӧN�UTS��QQ5$֌Z�q�UV�%�UEUle�C�cIV�Z�:t�ӯb��������E6������PŶ&)1�95Z�5��UET[.��b����KXu�"���l�4N�UV#�SE���b�"*5�
�4iֶktĳE@E�4�,V�4՛PLMh�h4�Uh5�����[m����(أTEQ6Ʃ����������m`��ckw�S3^mDű����5F�EU�UZ1Q��Qb50�Qc[uEEQ�TPI�V�CS���y��ￗ�+��Ω��ȳ�p�noqx�^��.����u�e���$��G�n��x����cn�yF�(�C�L�	��}�k����ίs�4Oԩ"�]�� Ué�����M��s[U9<��d��/S��BKy�m� �]@�21�E�g\t��ؑq�TfΑa'љ#��v:�O�i)�4�Xe��k['�Q��Ɩ�Ӟ:�瓆Ud�{��/����7����3���y�rJ(��	�$eos|�3�����](�&�>s���v��U�h�0r��&�ī��1�%�ڲ۹�lwLE%�#i�z8f��{��F�s�_D4WC�<V	'�ɽ�{�Z�v��Uz	�7=��w���.�?b=b+b�Fb�z��z���i �z�~�@�[>�pm���g�g��˚!�������3����8����}��d���#C�90�8j�aG3�FL���u"b0���ln��̲{��Y���br�ё$ְ;8Q�r�D�fY:�����Rv�n��(��)�{�W0S:}�F����"��ԧ�:7��LӔ�ۺV�F�}��,��d�}F|=��[9g��"�.��D�}������R�*m\�S��/N�s��i�!Ē�bu�+��5(~4h�?}_��!�,צj�bH8�F�����EcwFgt;��4pG�(ϵ[���`���ꧢ,���MjV/�6\[�t�r�/��3y����Oh2�TWk�xs�Y�]�=�JP�g{l~��vG/1:9\���T�!]H�7�%�gUQ���M<	�p��\1C�YV8��[d>ū�9�%�I/�V荳�ᮒV�T
H�ǺS�n��%�Dh�U1Jr��K^�Cn<��϶x)�GY�!����%�R��I��͕��{���w�>t�Fb2��]�A7����:�*��\i���"n�u�S��f������fF7���8oxఛ#�91�iJ;�ꭳѽ���i��k�9;Xk��I�u+��|l���}[ϰQm���m-g:�9귑�t���yP�ܢ�nϕ���a��A��L���J� N����-���2��M��:��)�U"����U����^��}MV��꭬�}�<F�#�<�O�T@'�hᨳ�0��,�J��˳%���UR�4Ok,��n�L�xy�z�L0��>��#��}����vs��ؗi�s��]a�pY�&��k�ދ��b��²��U�
���o�DJ�^f���3���!�*TO�uW�oK1���y	�C8�n:�VTu#@'�շ*3y�a��q6Nv�%�z{*�3T�$7�c?�H���!)���'��=Oz�
����R:,�' �:+g���t�,�M�Z<;�G�,���NW຺����êd5IK玊�y~�_2Ja��]sѰ�����-3�K��B�Ä=�gp>��k�=ȋ�k^S��T��;��S�qOʸ�KZ�W�h�/[3bb�^����J*��H+��%`��;��(cu�4=n�ջ\��,8�$@��D�{���!^�F~ɪ���y���#���%%��z�:[�ゾ�9���v��� �j�k��W{�"Y�L
g��h�A��!�e��3�W �2Z���F�dA��h@R���?7%���|�74ieB��r^Z�������]x� �b͜�+�����@����]��u��쨱\UY�H������s���S7{z���3զ�~���M�srW�������>o�%����gCd�^-x�w�.m^-��x���?P~��5ө�pE@�����*�O��6�Kc b�N������T���Xǅ*��l�b�)����n��n{��[oJ�3z�aE�ە@�x6�'Mp�%_>���lL/���魒�&�	��8�s�_�2���iwj��J1K�'vA���L"�jj�^���w˝匎�5C��Dn�Ma_U)��4%�Q5��^ݷ]N�?V����2p�gj2�����1dnH���g��s<��;BK��W�|�^hῃ���}��m:Clo3�����2#d���Zg�*w�	��'�i���"{���ԪX�1�b7 �S��t�1�皟J��&���:��_/�p�\��X��1{E��]����+C�a�	F�H�(ŶvC�t{(�����tC���i,B@�Z ��;��WΠ�Fք��]�D�s����q�\��l��q#��_�Ռgۜ���f���fX��^�z�jN�;�u2�J쨍�̲2�q@؛�������q<��汲�Y�e�}�!�(ưr_����95{ܖ�����+9�J��Q��M<���{7f�D���G>
A�������ع�hv��֑G�%�cJv=�9	�W9��h�*�c�,��F��L,K�cdw�*����f��g���3�|m�n�]ٓ�s"� �(G\���v�kWV��3^A�n�<[2i�#4hԼ���FS��n�U��k��'!�HtV�\Y�nE����bB�L�q49���*�$UP��{L.��&�_D��3sz���k���ax�%|�y���K�M��r�=�C��i����z_n�0Ȱ�Ќ�l�ݎ����Jk�.An���� 53Gi�׵�Y��O��pk^����"6WtLwZ�Վ@�IET�,��']��j�#g$�\�5�>�\3a��u�}:��-a��0n���rl˓|��In}�s��	*<�FHL3�̀F��������S+�D���eZ�y�*�o�q��Y�R׃� #�
�_s�hf2C_h��h=\��j��p�դs�w9���� ���o)���u;�+࠳�JQ��o�-l\��`x�$�o�qM�7�ꈩ��b��Ѻչ��s�U���%�=يd�6P�'p��-y8��V{ж܋��s�����ҽ���&ϢNO�Lb������8��K�����G�ǝ�j5��R:���/�:��� �p϶,؜����������}��d��'�/�Y����uoϾ���&���@B���b�Z9:s,��;��Q�g���Ⱦ���>��l[��>"�]��f��Ó�I�,[Z��<�fJz�؂� a�7�Ee�n�t���%z��6x f�e�9s/m
.����e]_na� ɵ*�]�'�*%��agA\Du3��kgT�Y�j��k4���܂�䌛�4gUW��O�i�'���e���1�)z�ƻ����'ml딕��x���T�IWN�M?k(�p�o�;�v��C�.F�
o��9���&��J�=
Z��>�7+#N6r���9b�Ur[�5
̵u˺�������6*'D�s^�T��լ#v1��W�Q���ܙ�/7���/���"C厂�Xf�Q�2f�G�,)?gXg��X��bX���B��v��qs���X�塤��7֎�N�wU��_\
%�Q8�A�^3;��@�$y3��pfWC{�F�:��k��U���r���X���ڪ4qk蜪>b�vm;����T7�#�91��-�ozs5j9�ϙ�{i�T�]���T0�l��`� }[�fQ���d!t�a;9}�]��8;�*�r�[���f����9�|�@x}W��O۟��0��#��2�� �� 8�R�] ���r�9"�\
Q��su �P�c�B4�T�8�؏��1�ϣ7��c��yRa�1�s���g!vh@�����䄧0dm�4	�uW��{�,�e�n�<�0VΫs=��ѣ��wY7��%I���N��o�\��ĊϩV��aJBQ/��z~�� a6��*���ި���7T{K3�\���d=� ��;�6D��&�#mP1o@�YO�4H�~͝���Ap(m��-:^T;�s<z���q��R�-~Q��\{�@��wS7}a|;6��p��Z}a�q^�u�vAo�Z���r�&���0��:ۘ����\��ۭF��'�/�.��;]	z
;�bֵ�"{E��s����P|{p�VE�)m�	���}yJ�\���UM5OU�+kT;4�C�'"�,K!�v����T-J:�6�V�F�6�!�������w�54�E[8!\���Evz�_�O������U)�����+�Hp�=�O�{,�M3��$FHhJ}��F��k��<5M���Gqٔ	��G"�sy�HÐƚWE���u��788�*e(A=\1��l�����w���+���t�7g���aNAԮ�5��l�'4��E��6Db�Cɣ����č4uZD�/ڌ�s6�Sn�]�e�j� Q��y�9Pٮ�ӓ��bif�m۸mB��9F��8' �/7~��'��r.�����,T:eOGY��uMBwn���9��i�n�$M��d�����x!΅,��ܑ���\��Β!*!lV�V{��#����j�
�S��f�c��w/E�Gc�3v����ox�QG v8N��xXO�^�f��
x���tb_wLgb�}_e=<��m�t��Y�_a<��;F�hI8c:d�-�
�u�;u�x`C��u�y���i�u��~�h�!�y�sg�E�6��2��׏[u��l��q���H����48��c� tQ�C]����R��r�ƨ��DY/9�Ϸ0�����O'�Xƞh�gb��ؼ���{_��BN��u�h���l̮~��k��9�WJv��)��q�C��\׋s��}���4lpU�F#���.u$:��4�ó3�u6��3&g�*�"vޘ��3�"���|la��rjV%Y1�;����ˆ�-�Ǻ�*,tN��B�;�j��ˉs!:(G\�<jYqm�;Kl7a���|IU�1኉�RFUFdn�θW
��<	�NE��k!�t*�^/#z�t�k-� s�@mH׹��%R���꾺u���:`6��319͋_�^C6���hJ{�=)+�6ɞ�쑻[��<(��OV\�砏@J�/m,�ź�����T�w�x�ŗ�����;/xsRV�x��Y5��\���Hq�$��}7$�� �f��OP��Iwdݞ�`�Ǜ�n8/l9	��r���%}�'+�us麵��X ,�Ǻ���6����l��Y�1�_�8��t(s�����ݎs�i�m�����~e��;6�n{�͖� ���[u�Ԃ`97�fWtLvv)�\��m�;x�����#���.�^X����]��]y��������ɍ-{S�&��f���{z���'OQ�1�T*��6�8�1�ހ�W��j��9��ƶ��Ǣ/uu
1�k�u9=�������gM�4S\"ۍzE��wh�.��(P�ݞ&{��ULw���;!�\�b7p���5��2N��t�g1����QJ��r��5���	u���l���h�Y���mT�4KǠ(�n:�R���otǳ,���C�_'+��+H�Id��ŵ��`=�0	�b5m�zu��瀅{�hL��ÄzM��3�O5{�P����A6D����a�������vTg����O�	������T@T_���!�̢��������ňB$!@`!	@�� %D	@��P %D �P��><!"b�`!U� �B��\� 1C  E �� 4J �H��H���w�b" �" �`� "�� �"�E8J
b(� """" ���D% ���As�<f Pd�(!�
	P&"@ �!�  ! ($ "	@e1��� rEW  @B��@   
��x⪰���� *��� 
�+"��b ��P %�v1��Ȁ�0  $30�,[�S+����7��X������L��?��[W�7����]����;����l|�A�+f`����߇���"�����Q_��H~�~��@~��?�}���E�������?��>^�X{?��_���ߟ��o��(
� �
� �0��  R��  P��
�$*���Ȫ�ʪ�*�#"�	*�+ HH�� 	( BȪ�0 !
�(@ ��������aUa! `Ub  �  �@ �UV�AP9��Ń�������(��� � )B�t�������~��ty�G�?wʪ�+�_�>����K������z�O�p�AUW��K��}�?X{H ���E����=��?�B�(����������.'���f�����8i�<|TQ_��G�~+���QEx��6�}��_�����������S�ª(��UE�������h?��?�П�����{�؟�`���UE�����!#�>�3�?#�}������UW�>���=􊢋2?��[��o����?��d�Mg׬���}f�A@��̟\�{�O      }4 �                           
 �ڶ�Y�Zƭ*��Ym�vwMm�͓ML�c1j���MLj��c��m�6󚫠��-L����5�VVam�j�fЖ�l���ֲ3c���_\����KjT����ee�Χ@����4b�m�[3`ݻ��fSa-��u�wH��h�KL����V2�mmR�[m5���L��Iժڷ�ԗk,٨�  7��w�5U�Y{uݯv�[];�w[��zwvҩ�+=n�ҁ�{n�jWM���n]5�Sy��[�N�;-۫M;Uu�eK�5J���U=�3��2QlY�Sml�  v>�hhhQ�(P��{xt�:(P�B�Cwz<=
(H��ؐ��].�
(V��7�����뺖Z�.5t���{M�yҎ{�t����5����&��ӫ��u�L������&eCie��U���ݎjc�   �{��SM"���׻^Ƅ���m��;�f�s�Ƿqv�9�1���f�޽����)�9�7j���Z�Ww]N�*�]]3�{zzg-[vԻlm��aweUk{��k6ov�m�����U-�   ��!U��7��=Q��WaM�lU�����z�{m�s�N�o]9��U�MN^���H�6���ǭ�vS^۪)h۵�X i��sF@]�;5m��2�*5�9�)�m�w|   �-��g4�tgY,AkV�t��%�s����Z��Ƃ�)���h��c*���=�u�M-�jB�Y)Dֆ�����lT��|   }ﾀeT>�Ӵ���]���UZ�I���Ѫ5S�b����GN�5E�m���Qn�� ���"tj��N��զ)G�B�sM�iV�   {��(�4Z_m\6��v0��wu��*�;�K;h�V�2Y֨�a2� �X `v�\ �,���wV��nM�J��ڕݜ�   � t��� ҭv9@ kmm  �� km`@�0  IaB��1�h s�� 4�mZ�l�k`����>ۍ�   ��  ]u  u�  h��� �  ��ph

;9��  ë(  ڦ��M�� h�:���Ͳ�ԁ,m�on�c�  6� 
 � 4w4� ѡP�  :� �� A�0� ;u� @���  3r�   �{@�)J� ���1JR�  )�15)ISM4`i�S��R�����4"���UCG� � �*DM�T��3S��_����1S�����罳w�]1ଆ�ў�d?&`��x�ٟg�}��}��V�|����cm�m�m����`����6�����6�����c�w���$@��W��0����*6��f�󠚷@��vN�9'c�����e��J0*�v�B����՗��e�*��
����5,� 2��h���0�}�}����[�e/TxpN����$��SF#v��&=�S��x�{�=�e�{�*�A�93�Uf����Ȩ՚Y졞�P���0nu4��oc���Ⱦ�9���:�1ź�.�1Ն��1���i[D;��2Տ��wj%�勝�^�e�]��F3����Y�q|��c�ޢ��r�HyΝ��!��C�u�q��Y9nu�a�no�ݲ�ۃ�	�&=��ٰŒsA!5���sf�Gu��� �M�XG�E7�C���;g^Nʰ���k����.>7�+�����$�9�F��v�Z�{"�ob�����e`���� �f��F��"b��*�F��giz���X�5 iw�"bd��M8��ưv��ݪv��-�����E��׆�w_\u��E�([��)�.�A{�)��1�;q">ۛ�5���X�N�bS�pe�6\���ܑ��LKr����A����"�w;7y��9%����a Y��H����M�^_����Փc�7Z1�/,vv�ؕ̊� �����<�]�>�I!{�9��-cku)���L�$� �]a���غo(��E��4�r�42���ńjE������Omq${��c���l���q��H�3�T�j4��lj�,�+[��t�zEk�1���9��"�
�xvߧn���f�Tv�!����L����4�~�79����K�hu��������XY��f��3~�W{8t���a����1���ˤ9�5��Y�_�+�����<gu%��7�w�>ԗe�6��ͽ�,�Y I�����f��Q��⛊0���j7z4� Zw�,�u�Nl����w#e��]�Vל��!�&�ҳc�o����`�`4B��B���{�,:�U�p�� �vOq�`�Q�R��wh�8f�D��d��\�0����frx�׃�n�U�[�t�E\��>9��m��=�h��Eo��֥OZ	gQ���i]�{
f�Y4,�X̧���ӕ�R�� �G�0j��F֧vvQgi=l\�����q�svYӁ67��n��)�y2(�(gHRL��ʝ��Kl�����U��4�J��z�oP@%7��-��J��th�a�u��ݚ9I�2��琞,>wbW� 띣�M΀����O|�w��v�ӽ�b����h�ԍ����2T�խp	h��=W&E�lպ�G�no]�wLK����>�MHm�)w���f��-s5�6��qx��\N<X����n� 
�c��J�o4��ӄ��y��)�����}�w�pj,L%W�=]�r�c��M#�����X`@���U����ޟt�rM��3Q֏nI&�ȉ��i�'n��e���<��	���'Ξxң��r�V�#��\�a<�#�3�pY�CdRXa�!j�|���/=#4񽣳�
���	�9�5�*#�]�3�s�H��hUK;�z0�n�1-�� �wt���+
��p}�O&��������t=����'��3�:�h��x��!��LӉudK����8ge˸�Y;��Y������b�ye+�l����݃s�<}�&�X��|oa���;;����+�C*&9KV�m�y>	t�zQg.��F�ukXy����R�=�v�Y�v��<���:c���z�qf���'�*7��]�*�)�e�|��^E�MB���,}&pT�v�ex����B=�ZW+�ՖK1�E�i�Y�ձW.ډ�N�<:����˻��sJcOD�FI,Ԓ��[,�rӋ�e���q��µ�;ی��@����d���3v����h"���F�+�@N�*b�F����<M����4ӊͽ���k�@�X�&��om,e�裖�o�HG��J[���B��]+y/%�i�@`�a�4����,ڱ��'�v�@�׋6M
�%Ʊ��%��� `kI+Ӂ%nMX��hk�6fP�u%E��2r��s{��; �َk$���)=�pڎ��C�nG������鼝ڠt�d�K:��e�Mx���.���76�݉��pr�V��6~9��Dw;�Z
���ge]��v�B�� ������:�}1�Qu��m�P�n4��f�RHޭ�sF��C֚�Ƶ��D�c!W�*:{e5���IU� �Qg GhSGu�,��X��&\qױj�6�B�dJmyU\�ٰ���t�ڈ�%;9�n�U�Y 1�W7ٻ�"j�C��9�o1\�[������9zDn�p�.�K����#cR�i�ZOq�ڏYܝ�A�Z��ru&����s��b�2��ig\E��t:l�/���0(�m�TW�q��!
�y�9�eVs���xo,�	 Dm��Ǣxֱ��w�5���Ϊ��a����^�F�s��{��v�����4��t�01���ڮ��N���q`�tD0 �p�L�=�[1�ћse����d#p�i�#G~߻6gm�piPA�px�f�Z��b��R�.���#{5>�سF���v1]�4��Wh���*]h*���|hʩd劉[7;�:4���sY�!�y��� 1R�wF<����.l0bb(�%sZ��8��5M��]�I���ú~s��JK�j��.���y����\�z����"�*6�wIJlT[���[�/M[O�;����c�>S���l�:��ָ�J�aހSN1&��:f���9��u��Cᣚ!�M㝔�@oԣ��ڇU,ս�Ol�5�;]Η���ݖ?V��ܜ�.Q�����u$tg!��	-�]����g:{-�*�^v����Ά�[z�Y �:�t�L�хt-�8�װ�gn�0aQ�E�Yݩ��L��ӡ&�h����7�2��oh�˕��Y�v�6-h>s�Z.�z2ul���Ι�n=$U���=t�wd
�@�Q;��q]����5��F�u����H���]sV<��]���99jƮg����
�V�]�s{pry�$=/C��'F�ݶ>�%��*����^,�aQ�L8��/Os٧HLn��jD������O\��^�_:V\�ޮ�z�Vl�w��`벙p�j�KL qT���r���3���'wY�;,U���g��(widyw�����8��;��ojᯐ9�r��U�M��t\�MX�#�n����b� }SˀJ7�1+��ŠÝiá�]�Z%�1�
�vv�
�}�:E��6�v��0�����n�0��)o����`I��@�� �l���u 1D5�P�1@6�"�N�:˵l:��k�Ѽ&v�X���WF�=հ����A�v�Ԩx�a0�aw{;w	�ѶH���b�Yq͎]���}�Lވ7.�mȈ�X���cPҺ���yh�cw[��o�p�]5n>���x݈��e��!;�3܀߫:k��)ӻobk�����ѓ���q����0g ����t �d+��i�y	17�|8��)��� �W��w����Oe����.v\�;�Cü_e�G
rG��g�]�Y�1>%��wV�W{�Jk���G�cjn�;��k*�\�3��7�I�Fv�UD�	��*�r��ݲ���C��pgq�uog�UO�5��Oy�Ǖ���u����4]�m��9]��׿Y��@��;#[#]\�z�6����!�[�{M[I��\�Y�B��j�BC[$<�
 �5�)D��y�U����+�s�g�l���Zyu�O�`��z;7.@]�z����ֺ^�wS&�����#s&64%Zھ�ۺN���s��7��{�z3�\�>��ޚ2��!���e����wtwN$\W���Ҧ&X�4��ԝ]y�.� ï��0Y7��8I���W�N
؋
Ur��ޅ눪�s{q�^����E�y�C7�HM�Y*ttv��-m���L:8��1ޠ7�P�fՍ}�o4Q�.%���k���똻��W��$3 kM�3��]Gm\�����<�8f���]8����]$��]�&&���E5+�p�8P�xtьڝ��ʟ���q�d�q\ֺ.κ(���ě���H�8�Z{Wa�v��V�\3nK���.��E�[�.]9m�aa@>��Q�$��&L��=�����ɇ)%1MGPVŨ�T��">"!���;sN;.�(*��+7�A��U�	@�[���cXY��8xB�M滚��q��v�0�v3��2j�9���1��eثp�v���,�9v�K����Uū����CΌ8��ey7w"z�p����F��%T˱66jV��z1'�m�� tQ�P)X��U"��7�;Xg����zCzz��\8{}���r�p�;�PԣU�w��f�:�� �� ���-�ە���J�^ڈ����Vw<��R.�ꛧA���H��bŃ:�Wr�,�NB���8��U4ڪZ��({O>��Y��Gc\�YɆv�*�Û��;�3�0`�M��d
�Y낇��'R�4���)�g|�����pL¸txn��ڍ�j]�7j��f	40"T�Lk���_u0���
��)sr��9�\�r9n��{��ɥ��9&v��� �3t�[V��Nq]E-Q���l�h1"��lm%���>+%qb�;�JD�m\���8��TJ�A����oF���.'g/���N@���з��Y%���{��ӫ��G�Y�*7r���]ݩs�&�K넡w;�Y�vr�**�<����%Z��N�J��΋������H�ۗx#�l��v
�#$��ri��5�U�׺�a����ݘ�����Q���tA��\�^���2N�R�\��!����`��tC�-�x63��c�w��W�(��J�J�79��׽��3��3s����ذ�4��x[��z.�(;q��Wa��p��3�;_�d����ո��%�2���s��7;vt��k��{d� ؓ���3�
��G7������N&`�p�$�#�Y��f�\�x!uӐR�g<X��j�xe;��
<��Z.���޷���wXBfݫ����D����!��:1�x�w�b�ډ��<�1�]�u������+�:76@�z�h�\���np��3zh���J��8Ouӿ1��畩W@.�i.3+�"O����E�&Q�͎i�I'v����0)8$�N�[��r�*��ǋ���7b%�SeE[�<#X�/b:���z3ѝ;�t��I�V�!�n	X�ٳn� �aL֬��	雹(7��@�Z6�'#kqӔ���
�����\+�w��I0p&���!��r}v����.M�������LF�k��3�''�e�Nq 6��y�[��)q*�w���]C���R���/'��w7y�!{;5 ��U2�T�����]��G2 ��'� ^r����no\?��}reHv(SӀ]�t��4ZqGX����bS.�˃흡�����~1���ݲe�FS�����/x�hs�_2�ø��|�ë�q=_@���	��j�Dr�7d��Dkub��N�����Y/v�t=$�=�$c�) �q��ܽ�1ʂ(e�;ɳs��Uو��܇�r�Nyr��i{U��|�b���F�s�vv�t���L@�;X�h{���szW��ވ�
/G�};z�H�ܼ�K�V��̓㫱<?O��*yugh5�0�%R��n�݊M�r�غ�8d��!�z�i޶}	,&n9��;GB񹳆�~h!�1H�A��׏QC����7��"�j��"�U��e�J٦�5j�en�ٽ�;//?{p-�ۛ������P�w���a7�����X��m�47�Hժ����F��P���,tv�Yl�rm{b�3׺�&�,���	�&9q���{�9v�<;{.�mG�D�F�3mX��Xe�����#ýޜ���-x1�p�'!o-�w�RZp�F��4���2)n�Ĺέ�C1<S����:��ɩ��`���
��A�GDw)�^l3�`�������u�cH1s@�0�|3�㭳ۻ�su:�oP��*.��j�4��zˮR0w�o3;3�Ky�0dі�3�gn�Q��K�-oi����0�{�[c��[t�>6����7���y�F�jJs��7�:�cCOIx�h�nh�(�/DJ��#y���E��zNμ1�����3h%��VC�a�3^q2<m`�L.��{ۺ4��-����uoڳzX�8�RmVs�]�5�4I�Ch#�<39vYV	��C���Xy�. W!�z�Wx�m�&��^�ݏӝ���d��ucp-���M�a/{��U)ݟv���>���w��ॎ�4^p��*�����*�|Gl�]#�oc��۫H�H+�2w�=p���s�M���G@���T�9�ޛ��nZT����}�5N�& Sn��cnk]Ons[�epk[+�J�F,��E�5n��o+H��I���<B{�m���=����q�.���nH�;ݹ��t�7.U�0��Z�wk㫹U��C��8F�,�fs&;ǆ\w�͒��ĳ�����'��������H<��Uܸv[�N��6�h�^k�9B�����rrx	�����x*�SP�{$�G�o9;�l�{ӊ�p�p�H��t�W֗%�Ć�$Rba��2��W8�5����m��C�:/���Ҙg���FA�Dz�����hut�����n�qF}5iuWP��c�	�k���ھ�6�K Nڼ7�ؒk.�̈́��P�I�'L��X)f�a0���v 8�û��4����1���t4;��U�I�:����C��Jp���:Ѥ�ԧ'�a��"��2w.Iٯtkg�U
*:���r��ͯ���7��q���*l����F��D���nY��SF?�����^C)���4��I)����N�Q���ujELnڱ�:�S���A�����􊦰��N��%��ꊲC�;c�9�N�C�f+�ܤ�oQ�,\�ŭ��}����-��81�l��'JgV̹4h<���#E)��깬x��7T�o$D|{sچe�[�4^���ڳ�?��|�<��.w=�݊����� J}�[�j�������z�}���G"�rOl1gmw�ߓ^���왕}����9��%&�{��Cj�Ѓ�Â����z��pn�e=;bU5e�g @=j�1��-�IN���T����#ڐ�	Vnv���L�h=��M=$|���Z+;�%D��݇xi�4���76(�25-�g"Fm'Y1)�k���
�9�k�.���E̗C4�q�#�͌H��5a���/�`��uhۍ�:���}�����Ԟl�V<�k�۠a�y�??S�����L�E�E�Iv���{A�Ѥ"̤�cje�\��c��]im;��5�2�#F�ų�xe��en�h�e��-��:MM�(��헰`�u2}�Ѯ�WY�<�v� Ip��O^K��$m�c37m�Y�U�@XI��r�j헣kj=�Y1f��	�\K�d�y<8S��칪ྻ�|CU��{]�l�6nJ��n�8Ƶ���)��Z��J�}��r��6��B���n'�i�N�R��z(�q��/OP���Y�Ӄ�<;ZV�[:f���ݦ�c�r{սڅ��ĵY'!s������@�E�h��4���+e+V�!��ѓ;.K��Y�B�	fh�^�i�x�^��R#��;n��j�?��z��׺T���sy�ڙEss!�$�-�e�׌M���pىb[N]���
�Ԍ�|;C��G=1�zUx;��j.֘�y���u/9�y'C�܆L����3�O۶������zw02?\������]]��F��%�3�zq���EJ��d��cΛ�8�1��e*ũ�Ƥ���#�\ad�\U�`��i�[�Q��V�
\��Z�<:�"t�2^͖Pv�[�\/{r6eܹI淒�`Q������;��i��&%��5�g7"#&�f[5{
⼰�n��e�X	,��!4���K/OC佸���B���|٤��fn�e��O2j'
����][L��U2,(+x���m��F*� �.���}\M���c7�J2��x�K�
�K�����#�0aW�D`�a���&l/�pT��Kާ=��Qk�{Z�{��΢Y�^7�U�J�n�M7��i��S�N�̨��p恆�
�rᮽt�H�������B���FS42h��vK�Э�Pu:�q���F��V����m��r�Ʒ"����n-=�ݺ�~OH��u��ݹk"�krn�U[�3[Տ��o;�N��d6�X��^l�]c1�/;�� s�L嵑�CӐ��f eL�{"t(���90�K�|󱭴i̥V�e%�(�V�3#%d�p�L̜0p�e�X�E���2�0h�	�td���a�Rw�'�ݍIj�kh�ۇ�ك�ꚪL'.--���kV�>�n����)Ϥ�[�0r��B5�j�T�8�*P��)�uzƩb�=i�o�Fwj�;�d�:(b]zz�*��fthr�il�MX$@�4�z�L���U�p�!�z�}:e<ݕҀÒ
�l�K���N�T�<�~v�9rv���hwr�rzd�H���<a�p���X���X0]�7��t��H�!!��P����~o#�#x����
��ή���\b�W&�j/���*��	���F�3���Q�s�ن���a��WH)l�z/2�<{�+1�NN���$\�W]WB7�����'I��e�kd��ky%J��d)���uW�{pt1ٞNV��:p��wz���5r4����^\8�1�%!�wZ/��bw|���+��?��<G�Yx���O�~-����Bf`���9I��!��y���x�\�s���HsR�9��E��S�<�"t2�IQ��K�0f�rӣOo���e<�5$Dw�x2i���b�wj&�0Q�ں�-a�D�ꓶ��v��"81C]�O�Sx����0�� 2T���oI�
�z��Ҳ	r#4=�8R����ۙ�]��4�r#��$�r�a���v�2q����^��%�)���� ��f�jz��K5@]fԴ��F�u��:�+i�߽�x�7�s5�i�hLI���f��؁�T>�+:G��b.	����tS}���W_f�I
�����B�5�hA���o�[���no��k�8�\�xR���xl��7�tw�6p��Z��.w�um.jz�4�`��m��:����O,h˞{��ˤ�tG�,@c�5�6�Sߞl��D!�@�Y�u�bDT�S(�&�:u������Qђ�ە�|��hU�q�G�,�(d]�'���jѕ �ͅS9�fc�H(fgb��ǆ@+.����_-KfQ�����ݪ�E��ed���M�yh��a[�rQsF�ۼ�F.������=�t����=�=ٮ�oA��ᡦ�.���]ૺ���J��L�#ֳ�u�Jj�v�}�s�j)M#��]{/��+1C�o�ɉ�;�
���1�O5l�wgϲ�f�3Č��ow���C[�K\�K^W�{ҹ��DV�ѷ,E�q[��5��A�jep҄.�]٥lhfM��T�ˆ�!�e:�Ӭ��"n�D��]o�ڵ��H"�n5	h�K`Y��|��p����ΉrWd���
�6��l���}��.x�ޕ������*�eN�z�a�u��\?:��}YI��$6P �ɓG>�щ�4��/�"zm=�+�ޅ��!���^��U�)�NSV��&�Nܩ����ͮ��a�`8ͥ�)"����7lD�8jee���D�ա� ;��Ȃ��OW�]&��C
����:���r�'a�q5�o�A
ٗ	ő"!j��lt(8�m�B���vl�O�b�{���Tt������:���Yƴ�٠<]����B���h��D@�&7"+%�1�Yo%�X�[�r��$<7D�C^X���q�v�`͔�6��̝Z�N��1� S)ۺ	q�Foв��q]�-Y�o,Q} ��������4��C;gs�Mn�e��sY�pG���,]e�]����<�7�-a�j޽���m�9�56�xz���[�y��\h]�P �Ra<E�������5� C�x��͵�#Q�+xv�;�C:�^��g ��G�]��T��Eށ�xV��`�n�\�w,T��g��SqH��G�v���/z4����{'������Fq��U�We�P*��4���A~laT���c�z�I�&�����x�J�)9���KI�(�FY���L<�X�
%����uy�M��t>��8���T�������GyDΪ�3 ����WFr'�4��eZ�����J+���F�a3�z����f\Yj�A��ŗ�t0�T/|�'���p��W{��<[w�H��f�wa�&[ui�{@��Wm��ܔM|4�b�(���Ӿf�f�Y&�����e�Z>r�ޕt��]'�(k�{�Ƿң���q��;��<���9
��c{C�h�Q�wΞӶޜ�E�����u�J�@��\�b2�����~��ׄ��߫�F����rwgDCB�$��|�ڮ�w���&vH4��zC����:xb��Z��V�j�-�*��Z��J0ύ���P���e�۷�����y0O��k\�
��h��0B�w��kqv�R���	��Y�%�8�M��[�,:e�� `�  �rq��e��/��5d�Z����c��$r�)�`YZnJ�=���5�>�S<�eu��:�*ec����� fU��Y�E<�7��-�=�x�������>�5��h!Y���k�Z���e���X�c��mB��[�}s����oG��/M�Z��h��!Sa��[�;Uͥ�Rk�[NCY:����hKR��[���lB��*/��V�*]*	��
N/Pzc��촟���}�t]bC���3��̍U�6_e#R�:�&�����o�zU�)���q	]ZD�P�q�6S��'e5[�Y�:�Uy�P�J�r�'2�{[CN:���RN�fR�t>�E�w rV��mdוd���Uc�k��љc����h9��fS�ì
��7�Lvns�(ب��2]f#��Q�ҥB���,��Вj��9�<��4���Of%6�;f.\�p��G9Q�iVwK�L�y�$�V�P.<R|��
�Y�iWu\�ѻj��7�����J���2�4���7�}(n��#s���΃]�]���ms�4(�-;E�95��Wp)��i|.�0��古Y[�1U�;܄8O�3�>5��I�� f"�DܵMC�۝�9⏸��q����25��-�P���bA��a�Jʂo�p<�"z'�Q��s|O)מ�uz�hC��ڌB�W����G���u��<�����Uu�sC���utU��Y��z�<�<#�m~�QXV^�):�1mݟbݨ�螦WZ�&;��9E�b#�i�v��L��(�	����ʈV�_���W�^�)[��o�/o�"r���OC`=��p�m��$z�V'���ݹ�(*i�p�2��E�V^-on�%����`�X5�[x����N����N�����������;��ʒ�Ӫ��6�b0�ٵ��'R���b�#��2�SRQ9k�iۺ���G{�4�r���~���VM�hy��;S!.�F7��t���<�n\zc/���'G�#�vm�w2�J�)h�U��˳��ݹ�^	AJ�:���)w�]�Uu ���֩O:�ڮ��+\�����q�#�r��l�}�1&�G:������;A�k�����7�գ }�R��3o��ۗ��LҚV�.��49@$7��rmO�7�]�Č�Ԃ�"^�[��z�u)��z�Okѣ�+�=�J�;영�>"-
ܫIl�e�y[�vE`�{��1E�a�&5Aφ&z�WK��
l�Q�7!�H��4t]�n�����T�Itܻ���z2�̱��?��p�<���P��gx �8_��'��8������vz�R��rr0Q��ۈ��>1�m<�B;�&"���r?Vr��Y�`j����a��JC.Y�Qv-�ΖS�qQ>�Փ���,�4�u�:]�����r���|�C��%R��Ѿ	�Ϫ]W��8�lA����4p&u���c+S��e�.fK����I��ؽ��q��9(bx���U���6��a�ˮH���5��w;=B7��]0'b[�L	�5�c�����
�%���ɸPL�q̖n_!\iK�|�+1��N���ȧ@Lc@j���m�1�̲pwk�Y*`{:�n�GL�����W2��b�qqc.V�W$]C�p��7ē�� ��u���/�e�U�@SZƍ*�A�̶vŚ�<M������[>��_a�ɯB���и���ۀ�nN`�L�6{�Iq�C�1u)�tJ=�"�y�6j�:z>�g>��9��e{�ǂ���a�y;�@9�K�&kT�h������Kإ�3��m�FuK�ЗS/��2�">�	��+6iK��L"�f�����J+�*��#�����R�J�05���Z��}��My���(���1��m2�$��ӛ��'v�j۷'�F�i�(��&�W�݈d�p;��Y�j〞<���L�	�nm�36W=X�َ�ŧ��P���	����� ����r�	����.��%V��*:�,�\˳Q|:��s�z�s�ˋR���TF.�Gt���:@��K��[�ڱ{����*� sgT۞�~��(�t��(���b�a5�	�����2s}����y^��ݕ{Vt�,���N�:f�����1��0^�K�TG&��H$諦f셊��e�Y1�˹n���ڌ.b[(m$�f嗷i�
4˕������s#���CО�Fk�i8��ޱ��j�.H�n�c�r���;��{�ӵ�-����V��e]�S�,>/E�fQ���21W�V�*��&V��������.�J����E�-Ew;U�ov����5�׬���mw=��ë�
���=B7�C�����}�p�ӑ�"2�*w<ʼۊ���ެ��U�۰�P�d�IqM5�e26+�����:�$:�c4�T$��"�����f�ꕏe�s*�.��������,<�TIM�U��su���;�Rĩ -�u�|�i�d��r��z"]3���j횝�����V`�.�p�'*����y�+-�[�/�3p���ƺW\��~�'��YD�re�T꯲Ud�]o��op=�Q�|�TK�8F}�Δ�n����j�5һqԗ�j��e5Ʌ)Dq+Vk��2ɚ�:"vN�CNDq���WZNX��%��_Tr���%�cQ���\�����Ͽ{������lcm����m�o>����g�3��u�s�K�n�O�,γfo�xnȕH�ٱ�رY�q<�P�Ɋ*T n-�L�w[��Ժ�zi�;%����b!�v��=y�o���Ū�k�*�e�j�90�y%ض�Kڜ���#1{WgM�&ʶ��b��6̮����l���-�f��A��.ܯ]a�֓'a��S[�9�T���Yw?�����5a�v�K�_��K��O� %��9�t�|�q��ܻ�XV�� ��}�[S��C���T�d���D�9�s�,��Ԓ�/u��A���JH��f�K.0*Wt��<V��*��pr�ewN��[n����sL��W[�y<�"G�S��॓��Ӊc�����q��4/w|��`�f�%ۡh� 7X�E���U��F�� 1�����@��-b��q�"��޸����	��c�*�íF�ל�J��Lo9�B�����QL1Zv�C�}<�D� �K��;��rm9X��M���l�V�*���)�lS]N;�Z$�\����t��-�p<�@e	�R����f�D�&�3M>�Y�u���Ą�f���҂���ٶ��2c�Z�W{‑����gR�;h4n���A%.c2p�<�a{޾D��A��s/�nDu��^���wR�k��fvYd�pǇh��Oo�QL�d�fjR-3\�����e"�@uv3z�cR�m�juz�	b ���1���}kS�V�@��twe��ɵs���:2V7���H@�7�w=�ѻ~�F���EZ�H�=��o�`Xǈ�>>j�^�PU�B<눅�;y��Q�V�/�����Ol0	�*1T��ن�wt��!�%n�Hֿ��9�Ls����r�+��8/7p�C��"�XI����7Zg<�^=�*<��T�k�����|)q����������v�6&E���<@eF�+�;�U&G84��&c�k�(�ӵ�r(�k^��碉��nZ��1��{�����
9��Z�J�a�6��ͩY9�
���:�!FZo�Q��]qmƚ���q�%\l�gD��Z�VS\ �2.�����yr ��F�������8G��Ƹۄ��������v?��x��9M8����{�:B�ٵ�2.�c�f��|q�V��2EV����v����5��L�鿖mZW�6�M��r%mT�n�٧o�$n�Kg]���*3̈fŒ�z_�Ol���}� �<�+8���:%�����=����0�L�E���/Q
Z�%Z����]�*���5����~@�Rg�@��~�x�Zӂ�rN�%/,OOA�=<�o�p��j���ӊ��*���,6+!�n��L��K&KsY;R�iU�ٿd����W�XQP���F�C�����7k-u[��w\��;i�l�H�È9�x�č��Fd(\�넔u^΄�z����x���βT��I��"��]3�=u:ig|��>�_W
E:;�9FG��?�	!/ѿZ��S�nٵn�h�j�WA	�Fv/5>�R���Ỳm�D�c�	�0��`�z鹺R��pk���탵�I����<���u�����ك�#�5�=����[r"�V���I��gs�)�6��>��F��w�@���f�Ӻ#�[.�<�����[��e5�;;4X�qNTf�.cm�.�-p��FKn'��&��}&�Űa��i�l�[�ҋ+��kfB��hd�t�t�}ٶ�N��p�L��\Z2k�x�on>�H�rz���I�qTZ�\�D��]@�)%B���!&ϩ<��@;�]��1>˱'������M�5�Y��{�w��F�~��ؗuen�^�v'7�1?.&����ʇ���l)�[3�v����M���|���k3���K�u��:P��=��`�7�pdӔż����4�9��"@R�|o�^L�\�7�6��9�À�X9ڰ\s���I{��n� ��nU/�Ю�������.�}���I���ek�p�]�u�V�dOyc�3�G��a6oh��s�?e��2J�[XW���B�"e�7202ek��]�7*���tⳅ~5<�
��]��{L�{F��ط������(Z����K	��u�j�e��ݰ��R�ָ��o}��+��9�p�a�1�kGR,[;�p���/k�J�9����j���'1lkTQa{�6�7f����J:�e�Ư*�jf s{nsS"W)r+sO%�[����#/�˓7��ｄ����9�f�%����-}�.O�%r%�ק%6���'K�Ӫ�VL���ӵ�=��;�uu}V<zA:ޭl��a�b�|
��t��h����;�7�����"ƎUu&����o.�U�C�"����%#敗r]12�Np�hEg�]��Ď�\v/#ԋ�HgIyS���5CJ�v��ȁ.)7����	�	b��y/��(+�f�4&�����׷���T+]�p�rĜ籹Vv�gg���ҕ̭�Ty��ݡ���c	��b!�N�9R����*����zij���-���5�:�*_�'��6��آ7��B>�:I���}��v9K�#[�s��r%���p�)�C�\�����zs-Rh��GN���#9�ڕ�N��u�J���;�=)87iQ�nۺ3���K���bϥ�ݟ,\o�"�q�OJ����9׽��k��H�j����&��d>]�[��C/l�"�P �^�ђ��G1jZ�ڋZ��aZ/��4�C��U·i�7����ӱ�����!��8����dɝ�5��}��vё����1�7���Y�n�����\oe��C�3���7NN�����
�r�[ϒ�^C��ք�@��W�cm�d+���s�l"֫͊Q�rԬ�A��q��=ZSR�,���0Щ�(V>W�傷�fř��IK��`�N�t�Y28��\�.yC"���FûŜH�_
��یu����w�5Ҧ,���k�v`_vB� 6�u�K�O+�5'��վ�t�uf��H7|��G�$�l��A.��4n��Os�¢{����Q�k}W)J,�Y�8>:���X��u�*)5��Ď�k���lu������g�G݇��)��3�A�rI�Z�x���,����U5��.}��:�X�c
%s�*J���΢�+g.'f�M����Y�򫨪A���_B����]r^�w!y���p�!�2��q�'���Le<rSHnj*��Iػ�,=� ��dͭ�:��1Qu�P�s��}y��Y�B�V>}�����j�$3�`����Px/+v�.����0Zı��f��؛a��b�in�~�·H}c�:-�Σtv���G�N��߀��ٷ�/Y$���-6d��~�gv໬�@�zlܓ+���C�[,�;W�nlk��JV���eP�;9��3�#b�2锆pљwSMbj���ե/)q�j�n���@������@��Ov^�|��7\���v�3�����V�aKٍ��� �;�;�@�r�]mL�VnV�^���}zhsh+)ǉ��\LՃTY*JRO���B���Y�!i;�5����X/'�m̓<��r��ɮ�9�{W��H���������d[���1z�҉�24ٚ>��rt33PЕdh�mR�j�6�ڳg�ں��a��[������&,�5Q_��l��_�mg�]�jK���<|�lඑ��▇4�m
F�������#{tT}0����V�h�*;��^�<��]��S�H`���r�duB6*�<�/6)�Fe8����3��,�r��/n��N�%sĚZJ�>�Whִ	ܳS���L�����Lw��k�eSB��ϻ`�A:����eG�xj��4H�S��������	Fan�K�/�K�b����R�2��dz�Ĳ�����]4�h��3r�s�N��H�ۼ�AN��-W:d���!yht�a�<�S����yn]�:�oU*2DU�j�j�[CjsM��t3���.��$idws/�1�m��K�*	Y��Ot[)Y�G�m�Շ�O�<+~[F�d>W����+��~$q#���1GH_Jۭ�*�|;�a9Oq
�؋�����]&�6'�v� _f��c���K;;z����vh/��.�ԆCO��Q��:���m֊ǋ���M��
Q:�M��9�BӲn��,K���.�`���*ab�W}�<���nޞ�����q`'Z]H�]���]=4����&gV��u>qCOط1oƹgrC�ܕ��΂��UWc݁k�:^��D���6w7VɛCW�X��b��C»
�O�{�+�	W�l�ͨ�i��]�p�Q�3���m�-��.���!@�O�Xcþ�����.�|�����
�g����6\��rk��Q��uqj>V_+��$�+����x���a��a�K�4�l�xMTd�ռ�����)��l�����hۗNeEێCѺ�;�Y���롕aZͤbo��߆�0&��ǘ�S�Ѻ0���,g	#�tc7���
�0'.��N�׋�����i�ވ�5/�ix����{��@���-s��zë3��p�j�*�]Ƴ^[/�J����C�[��˥y\�� �5�T��FS�Ls��L�׌��
܋��1��)к���
��y�\�ǒhD�> �.q��|��o/.]�[�ب�$le���x�'. �`4������.�C�䅇A����0U:�P����gº׳�A�٨{��9��x��|ʡk�4a�3r�.O�ck�ЩZJ�[V�� �pa�2�uN��+6����FI����7��ִ�o{���`5qgC��=֢_��=�n0W��t�sΫ���v�"ʃ�bE�$��.h��r<����Mx�zs����Q&H�&!I��'Z����F�}t��/앳�[\�a���f��\F�����t(V���4�� ��!�:�X�l��QSF��Y�ܮr�,�1�檍�pQ��ϸ��9P��Bv�q����=�e;�.�J2yB���\�C����{�}�=�i���iF�uh�"��v7(�]w�:0=/��@d!�x|�'�;�������aQO UW�ഓWS�W>�!�7W[-�V��<��3S����2�q*�[�@a���}0��%���u��oM֣��8|�ml������啭и��Ǆ���e�鶀ٶy"��km<�_m^�g�S�n<{]�=¸e�"O'cߤlp��uܦ���9*GD�	�����P��oU������<�p����e�VW½�"sc��x��W,�7}
���N�P[��*�%Iv2��ƹ��,�kSq�>ִ�|�\���0�=Q����P�l��ll�m,6��p(�)l��6��S��Ɋ�f�b(WSP��j�3+8ZE�$˭�W>~�N�.��F�C����{���Z�S�ɽ�ܖ�v��6�;}ɬs�Wq��o���zr�yov����4��L)tW�b�-P���x�0�nY���ϋ�k�1����v�5�"|_>����PXޭ�!793-��d�\�l1��e�ky�h%�[>X*g4S&���,�/e��뼭{��4����P1Z1��j���=i�>3B�A�`��Tq]	Rj�/����,gF6��Q;7D5\x����ٖ�~�đ����l%v+-=vq՛P	 ��.���P�%b���n�-<�Ui�-������pNW�Y��ܘ��8*f�n�yY��C���v�WqZ������=z�͌$���2�7�H��p��ڔx�9�S;pko��W�hc4779���4�kC�;G��I=�vG��s���P��<|���d�κ�s2�Т� �4�2x}�"�˥`Dx��)�N;+�P+�#�6�[��;%��)u*�sRoN��c�����d��|�x��c	`nn�"��Z&�K��e�7�ap�����[{؜��ׁs���ȃ%)�9�M��MS�n�7�R437��.
��)䠃��7�˳��Q3����̜�j���o���_K��R����`��V��x��3�ɐ��L�^��26 ���4�
#�ى�3�Q��ꑙ5��3N�pb�B,�E[�S+2$�"�g���w�8����{�n߫�qi=�X1�᣽�U���tm
j� ��Sm1�LլH��`�����˫R�M��5�4/�6W��DT-��W[����h��s��MeM͝O5�O{(�Ù���'.���c�y.�)v)��/�=�/����0��]���w�.����>t����Z�փ���Y[��tO8��!fUna���N��06lx��!>�`�c.똳t<���}���;�f�fvY�b�X,�Wa^�nG���}*00`�rG��"���/%��ɠ��g�N�����|��}v%J�1��c�&��V�k�{aFE�uv�&���0#���8�Qv �)�چ#��݅����n���5c�#���ñA�产���̐h�mA`cEV��N<\#-�we�76Y��ʇ%�{K`����aʦ*�LA����es����ϧBݻ�����"H�lb<SR)�r�t��"Y*I7^�;<��|C�kJ}��iZ�ʴ2�%:�W+;Yn���Q�u �Lv{L�{
�T�GVI��e��cX����؋���:��6� ��]�Iv򘗌M�F��ʹ�y8�fG*�����p��.��x�����Z6�&�Y�����+�Ñ�[Z�ހ.��폣ﾈ�>����;i�ʛN]�6ܚ����{�r�/����N��:���I�Qh��+fu���յ�2�	�6�t8�D]uغ�;Q�N�C�X�U��d�F�-2�{Zբ7gn�#4\s:�)�e�T�_r̈�}=a�%�����Y�\�cՀ< ���.���)E�lO��4���|Uom�ű����y@�s�����T栐O7�@wL�h=�A\����U��l!�,��@r�L���=��"9�3��19Q�=�w��@�|v�w`���$�|j���ޫzU]�H@�x�<,�h�z3�v7��BH��=ӵcO�u�S�%�]���-�/��fD�C�CO�s�������$�eKV�i��1�(�μr�)Y�W�OwDp�e@�]n�SV�Ku�5���e��C�r��TycF+�v� �;1���fV��&t
q���x�~돡瓆ӛ��d�P��.\=�����tI���I&>��+З�ٵ�� � �4�l�s��3��2��n�?��&!��O�	��Q�{�Ɍ,"���<h7�~Hs�����]V�;��A�5�pa�ݹa/2��Z`�婌:��ͣ�]�z�今��-;��:{ [:���|���<Ջ�L����X+�7}���3���/+���jE��V�	����`�J�Z�F=���̻�R�U(�*"9�L�D�F˓��ȫǜ��B�����MS�w"f��EP�Q��Ȣ".U\� �T�2" ���mȲ�s�QT�d�\̠�Ȩ��J�ATQ�(�VUDQ �G"��7.B�L�����Er(<BQȨ�¨��h\'9ra^%�ADG<��\�8G*���T�"8As�W ̃�Pr%,�,���VE���q%\���D��EJ$]:ʵ.s��J�:D��py(#�P\��5(*�(�3KQ�TjG��EM�Q*Fe���+A8A�ʈ�����DuB�̢���#A�)��*��WeZ!f>���7�Wq6=�w�]�ly�|{�7�]�.���x�ȹ5��	���YQ��'.c�J��n`��9���T'Ӝ��}���kI��G���A������G<&�q�o���ޫ/~�ܳ���=@p ֿ`��Q)��_%��ʵp�g�zXuB>z,)vE{R��Ǡ�F�q�t��T�O��y�ƛcNf�c�˹�=Uh����q6X���F�+�6���b�5o�/��'�[M���9�YRv�<}\ocϱ�C�N{��~5���Cj
6ߐ�Wh�~���������!<�D���������5��]��s�\�ugǕZ!;�{hv�֠���S:9-.���^�Ӵ������ ��_x���ϥ�64����g�+�w�;|�`orn��g�;f�i�Y�d����'EG�����W2��%�O�q�r{n`����&T��37��J&Ŏ-}���C.�q'��@�!W��]C�q���������	{��\��vƢ��
Y�e�{i�^��r֎t\ $�% �r��u�zw��K0��*�2��V�W�eI
i�����Xdlp�O^3��>�Y�6U�@� �r�$'�+�Z�Ã�R��֩�Sm�Ө��N8x�y�(�o��ۡ��2� ��7��<�Pl. Ю����f�1n^-i[]�5C��G�w�_�Ƿ	-��+�JY�{�_Nd�N@t���L4h8�Q�����	3�+���Ǵ���Y��Kޭf�go,�`��>�S[�����-�9<W<H'G-�?m�:�0�&� bfInwt���b��:_}���	�T���(�\.vd��M��%�S��N�#[�2&����T��+�aq4Y���2T3�j͌�9Pe��\r�p'd�lˈ�2\�&�'ږ��������m��q�U�A�yu�S_����!�R_��}��W��J~|:�w��}�R�I5���� p���E>P��"x���5`yE��ZSy�׫G�Y��V�p�4W����F���`X�M��{/s'� �ώ()��5�~�K�u��Ś4�pͻ�Z���|.9��-�'��l3_:�=��G�p�!.���>��fP�9��MƱM��dB���*!׾>�f�9y:�K�*���]���������J�_nb���}�Pn>����8�^���U�k���]Q0`9}� ��8s�S�l'e��j�{��5`�ގ;!��L��Is�@��R'r����H����}��V����=�P ��w����$lvg ]nGٞ!��:i�������NaΨ��R�V�v�m���ˀR&�6~�@�II����᲋X�e�Î��
wRޮ�,:N�W����tE>�
\��3W���k���Ww�%��A���[B6x
�ysz��v�s�M0���Kv4�9�9םG鸽U�υ]u��V#M�O�ZS�[L��t�ʯAhz�Ewb�)�d>i�g;̐,��Y)�:cuø3W���w&���N��m���Oh_uV؞�̄9�_�8;r2�a�o��=~��D�ƨ8�r#P�X�M�A}u�/E��\����n�ŕ5q�'�~�p�N�2�Zk!��a��j���]���>Ʋ�Wu''���	+�@(d�}�W���n�����J����Ѝ�u:;>L�0م�l���>=5�ޕ�(!s�"�J��X[�_�u3qN��Km�І�>��������j#�q>�"�1�n�FM}�I�?B���F���r(�1�?x�XK�b�R�.�9�=Tu�����Ԯ=6����>.
�ˀ��Oǅr3�h/��`�F�oX9�Ԥ[���u�q���Ü����U����H?���QJ��C�	��1��,���K�D)�hr�F|�.�.Ķ���C!��璮2��
�@)�s� 4!%0K;�h��[��0)Y(�\���7/ٞ���e������{�q�^�um��bC��b9J��Gѭ5sjwp��Y���$�b�C�Q�f���}�~��^�X�Hs���>��]�S�U=�\�ڷ}���V��%.t}\~>�"�����m�|/�)Ҏg�ry�8��uI�!�,hD�9m�oq���bՊV`�����忶B�+��g�_���6��v�1s�b�Ti�J*f��[�.�T��xim!V4��������e�&�l�N��Ldwa�0���Y*�|YU�ub��q��Hd5���Λ>�o���Lzʣ�`�ӴZ����[Ror3,�#.WQ[y��we�|�v����_ܯK�^�Xy9iA�&����]��/���f����@�sʶ u9�����YTXr6[`�$n�:�"��aJ�u�
�?n�
�,<�����g�C��4xS����fP�y+c���qC�0S���yfY�XG�+��Jq��%���1���c�U�<8,s�v]�u��>J����o:w�qP�s]̮����Y1��
�q6��� ����f�7� o�+�1P���'Td�1�X|>�����е�ص�Mj�ꭖk�YM���F�F��O>@rt����ɩ���+�ت�^�ԫIg9�z�չ�"�'�w_�8�6�Q���!�tl�=ԫ#�U�6
����1�Jj�mƩ��w2�A�YZGF�&/֥g44��gR���{ob�����3t���4Sj��Sjz8�ѕ-��pb���uu�xC_t1>--��Oꮔ�P��LLƜo��w� E*�#�:��B�#��߮��``#�nŎ@�2#��f̐��>��$0�6a7P3�ݱSp��U�.�Jܜ(b�%�8���O�n�AZc�^�p��)˖G��r�bk F :�UI�[Z!d�դ�c<�n��7\Mv���t��Ȋ�&Լ�k*\�K7_\$����Nd��O(%.����\��9�̾�1P��"��σۋ��o�oeC�����S��-��D���d��7}�j�`���Ǳ]�:��l߈���uD:�a�~�j@���A�Tt��mmeb��f���8z]̻U�=���2p��[���JLh�wՖ�p�K���j�P�TmѾ@ �F��0�fey
.{_�^��5�PQ�Eh�2���R�qaX�t!�'ζ}�O?����&�`nA�S7��Ý�wk!�{@���m�b�w�q�������<�X�d�wP���B��:v�/�K���3Q�ab�~X�}8���/��Q��:�z���V�-�*`Αȴ��e��Sީy��K���s�n���fr9SFb�$�*��L����;�֩���+;�X�*K7;a�21��T�"$�aml��]�Kj�`֖��\ɪ�c��Huؠ�M�>X_C��cv9za��n�	�
��s���-(}V|L��_XEK���{q�%w���7��tE�R����O��^�J;�����<���m��V�I���E+���t:aHC�R̅¶%�#]���s���6~RqƼ��d;V�+/�Ĳj��i@���_�m�^
ͮ��}���d�!�=�歷��İ�{�>kj��XS�-W@���K}�Q�������k���>o����n��gg �x���x�s��ΡL+��a���a��ӈ��gI�`Z��B��M��I��#�
�fL�Sk>ȉy�瓮���8I�
���E,��z`==���8+�&I��FEf��^�B�r��e5�w�ݠ �r�Y���h�{�)�Mm�Tλ�>5�(xSڱ��u�M~f�Hy��𕾅ֱ޴$��*֗Ӫ���<޵!�D�s3ӂTn"�(Oʨ<G��ׁ�;ǴU�m-�:��O�d�?eH.]�zW7i0,bn�Kؗ���F +�P�&qAN���y�����r����U����"�OEӅx��5hp*�~޸v��|�u(�*��D&�Q�������"�Eˌ��5"�i����4����JN�3�%�����iu"!�^����o�1�ꎣ7�S"���xE-�9�2X�W4`����Qj{:��NF�I���\Cc�nB�I�!��iMvD7�� �´��[[��d�ג��=G���Q��K�F͜W�FoR���d�­���]�;�~{M������̄�q��C�pn����Y�zH�b2�m��7]ÜB��+a;,GwƩ�9ݝ��9JJ\�����л�^'vʩ��G�j�:)O�@��w��[�hӔL)��9�J�뭊��_i��ՙ���VP8+�D�����j�-�Y�:���o;j�r�9wQ���/�*��B�,2��s�ј�ϡ����(l�b�M"xy�KD&��_�[�x��ع^�
WP�ṡ�����# 9���x�����Ei�TKd(�;��,���{�;y� �=^om��f5f�Y�㟲9õ;�̡֚�gEcVYq��i��tL�\�ǰ�N��@�y)Ϡ�BCe�:oԟ�S�������trɎ/�KB4��6`J���d/���0��u�p��c+�U������0�]�7|~�w�z	�ey�������=�s�"3og��6s
B��gHM�[i,1`:�ۛK,$�-���#`��$�!;Sψ��dg<�ηV{�����-C6<�tU���o�e��BF}Ǳ��Κ 5 G����m2'U�r�$�!Ms�s��Kv���>M��J�1> ~���MV
�U���Sr��w�E�z'��;�1���64=���	����s �����>O�(^��S�ɽ�s4m����J
t�H8�@�(�g�yW
��~'�#�D�H8hiE(.�!����]R��O�i�J]:����ҸFO�B.ļ�ћ��Iࡍ�Gx��;T��`Ҟ����7�*��H�%�?mf���u�����5Mo��e� �]U�t�h��^>,^�:��eT�O�{n�_Θ4C=5�>m���{���1���߅i��s R�S��d�t�^{]X:_�ʘ}vЬL/k�_��C��1I��v��dtx�\����8˼g.F�L ����C�k.+s۝6}P'r0|�tV�Ƚ����Tll��R�ލ���[���:�+�l�5TX`9��;>Mg�g�����8�d��gf�^2�\U�@��~>�(υ�|ǹeP	u�ׅ:������a\F��7Fv�$(�o	S���ҹma��i�V��a��4��ĉ�4�,>�/��H��{�L�e��ؓv�i�;_k�V�I�kWo�e��C�r��jS�O*T7fβ	�++6�p��I��`}1�.��1e�w]���θ�Ǵ ���{��ȷ�K���!�PV�X~�T:)��w(-�w�����n1C�1�	�`��,�+jLV�1�>],�"s8׷DdU��}�o���.~\.��(ة�}�WԽY^��!�}��M'	�m�\��p�-�Fu�����֮N+� 蟠^�Q�ې̩�t�o�}��C)��93̖���b�0�jP��w2�gѬ؞T��'�r {��`E^�Ԇm���6�79klxb��77��d��Ȫrx��1��c��Q~��/�L�Qq�"�;Į��y 4Ю{�6Q����GL8�#���Q�'i<lFČ�HK5b�{Ύ_�o�Q#"��V���h^ݬ�&C-�H��9t$JJ�M��:��/#�(ە*kbg��躮�(��ٚ�)Mn��#ګ=K �̯K�Ӥtyfq���_��hxX�5�I�ϭr�Z�oC�ܧ��jK6��g��Wy�������g��Ҝ��r�kr5.�?q��׹~��xW�����$�����x�>�1دQ�Ȏ�R>z,)vW�t��|y��-�J~��7�^'�W.���`W ��"�P��Ӗ�..���x�l��3X�{441r%��Q;щP}�dSV��+:lAfGr�1'W�)-.�C��4V�ƌX��rL8;�/m�D���X������̝H��9Z�:{��j|��i�r��Ea�G���T~`yŃl����8{�5�\Pua�gs5���׽��J9���k��1���?SF�L��\��	�X��Cj
6l��	���O��J�gJ޾^�L'.����l}q5����L�ֶ���d9�`��{M��y�$�#��mI�T}��ҋ����>����1/�ӛ��5\˜��S5V*w��ӟ;��r�ñ��C:���E\ߝg܁��7*�\�~�����Q���h�����͏��>� LI�<#�Z�E^���us;j`��<0���H[0��|�x���Q�#���L��N�M;ڀn:��7��JFɥ��p��܍y��v��me���F I��PT=Ρ큖C����w1�]Z���,�@"�1sW�2������%�/�l/�����̍Agi�ς=�s.%�h���h}�������-�9<W<H'G-�?m��0�����,��n��>ף=�%�GP�Ah�Rf.5;2d6��/:��u���=Q���q�,Ǽ[�0���W<�T�	h넝G�G2R3��N��p�g�!ؔb�v5�E�9wiޔwP�i̘�t�	N�nX��R�-Ov����\OP� �7	�M���<���a9�t.����_)�t�����S���4kk��)㓫��˻Z������K*uv�����h�;-(7�禥�����sx��,�@����+�w'5iZ�.5R�]����Mj�@�
87ٺ�.�����1� Թ�����OGB	���.�zp�����v՗z�6������_T�Fi��r�o�h�C1`'�{1���	�/����f��z�4�A�Wč��͝"����U]�pٶ1�"�����K���J�䉃�*�*�q6��V8m��9B�7u���حu�r�灧|����ć$+�a�i%]a�#�ŀ��olx�h��������4��Ց���o�}G�k5��WLq�����t�ݚ ��u]��jF{�*qH�ȷ=3���v�ٽ&����)��Y�%�Pd\��d�tE�)�b���!�#�J�Y�{�4OpOy��"DT�C��+v��o�=�瘜jA㕥�2`����Ǧ{ǔ���=�lP"�F��6���WD���=ʺ�ﰷ��^@��1�6��vAa�>Ϧq����mJ�kڦ4i�X;9b�Z%]�КP��d��2=�0�v�b�.�U4ԛΰ����!�s�e�?{ً95����yー���;Wc��(ʮ��8��0�7�Ϳ�f����H���Y�d����(oHE8
�Ix��=)����
gz{��h���_W��I���F�[1<W��CZ>�ݸ����雇Bf�t�t�!P��RuλR�X�Dv�e��"�Jn-k�C�>��j���7d.�w��eWװ�y:)�
�R+�u� o�`O^��F*U�]�C�jg��lr�٧���B_+�)u��^.����X��\�u]ҚN�;f�����F��|yڊk)�g^m�؍!�]�����ӓ��NRM�ޑd�N<ܖN����zLꟘ�l�L�}����k��;�^p )�x�F:ɷx:7`�,9��4q���G�Sgx&߂��Z:rgn�������j��.�9�`��sz+W3Ѿ�C���f�"�Z���/|n�>y�t�sf�T��Ҳ���G
�0��G��>p)�{����$X%�틬^�y%�wt�7*'9��f����jR}����q�����a��^�OP����9z�ys�[��aa�Pz����B]��#S�����Ƌh�s�-9bЦ�J�rmN��F�����
"���Ooh���X5�W9�u؛��\�{��ؔr�^dr�Nx�^)���.����-��;�1�ΰ�ei����E�+ݤ5�K=�����z�yyj�aK���N ���Q
.�x�/k�[g��F�ƻ��}��u�訙G�V*��.�+��_>��}w���\�����$�hEjib�Ђ"��Es�t�\������8B��%NE\�YUĐ��\8J�� I�EȎ
'%S�H�PTQEl�6yK�W�Z*mb���2���F��HDPsZr*"�$��2M�E�"�3�-Nq�DR�QTEDQU��FҒ�uH�p�ZUVIyB&W��$�J%���]��\5+�Y�$�٢ʮuUP\�K�*��� �Q�+��*r�Ԭ�(�2�D.RHL.G#25"��0��Z��R��aVJ�%�*9�9�,�$TE�1�UȥB�Q�L��Ūaem*A˜��$W3�F$L�:g�%N�s��DB�d���ǃ�f�U���<w^1��TS�a�kQKC/�v� d�4�i֖�#d���ʷB��̖�V�B�n����µ+����"��It!S��DX��o[=y���gg-Ωs��`�����R����&N��E	<C���(��_�n'��?{m��ݡ�>~��t����7��.i��<v���Ηq�	��0&1?_�9����	��iQ⶷'��ؤɟ��_�S>�
@
��__`	�v�s��}��n�v�|=���|L.�;9a�o^9w�
J�Sy�d�v�#�������7i��7���x����y�>&w����]^|z��nײ=پ\Q���q�11�N��7Q����ێ���=N����M�����	ӵ�O��I�!$� ����!�t�g�t��ǎCn;I�OS���~qҸr�?��>��������Ͼ�z�e�O�VmN���G�Ux|�W�U�C����ӿ!��w�{���
���t��	��۞F�'ݸ�<��z���I����y���������m��n;��I�ˎߓ����@�!�۾����V_��K�Վ�]8�z*~�t�0n���w����ѿ���M�v���x����������q���z>8�����se=N������y�����o�nӎ���{�mΣ}C����{���ck�8�vQ�D	��?|0Dz �1�}��>Qһ봁�vp���^;봝������n'����x������s�bw���:�o_���]���۪4|�}���UX�+�ƺg�H��1���:�x�-�G�O�~�@�A�?F'I���{��8����Ü�
��j����8�|���I���v��s��N��r�P��n�x��������p)�BO.so^}��wI����_����1���l���;]C�A��s�S�.��8�S�s�����p.��O��&�F����w�C��8t�]�]�O]�&wޣ�&����u���ޡ���7ۮ($�q'��a�&�br�Y�,F��ُ�zc똁0}�7����n>�z�S��o����޷�ݠ~HO�������ӎϗ�}���Wn�㉼w&���N�7׎��t���0��~�������puߟc9d{#�iȳϽy���L��B�S�ӟ����bw�Ü��q�ۉ�n�y�ӿ{m�c~w���|L*��_�����$�������;N���v���}v���C���N*N�o�O�X7�_9�hz7�����ރ��eۭ�]���e8n��aƺ�V��y�F���Bv:�#sƜ=�D�9Oen$��~a�^��3��.A�J�c:_cڵ|�w�M=;�ua��+��b��QߦKop_&�����#*���]j�ހv�.',����}���	�O��;����:L/�ߜ<v���.���m�aM���{�v�]�X>�������S��=���z��}��P��P�w�Y{q���A&^'�n#�䣾�P�R�k�>r�k�|�������e2��<����=&����|�q����|�����ζ� ��<M�5��x��T}���ʠ��*�V_Ӗm�"=�������1����B��+�Q5V*�������Ѹ���}ܷH$�qֹ���7�I�BO����㷉�<���;L=^�|;�ޏ��� t��ל�o];���y��߶�;��~;�����������i�9y*'�1����c�j������:w��aw��A�:q��8��ES�ܺL>F$뗏�����C��N��<���y�n�>�������쏔�l��6#φ��Y�u���|�~���|�n�ݻN/���'�o�����xv���ۉϛ��4��O\t�y�Ӿ�][q�:@�?G;To9z��i0��G�Aۿ��F��Us�S�TǦ>3l�L��N��/_�cL矾��aw��ߟ��!�aC�}�|q�v�s�n��&_S�n}��;w�k���y����N����_#n'^GIӷy�~#�n�<|x�T�?	��1�h_x[U{��8nW����q8���߽�ߓ�q����y�`��!븇��~�8�L.�C����o��ݡ��=�I�!&�	>s���ޡ���}/9��>��O���7OI�H�>��?|f*~ʽ�J��Lܾ�>���]����C��������۾�H���:wN����c�/�����sn�x�牾~��ަ���8��'��ǩێ=!�=���t����z�[���p}G�W���]Cۤ�k���;꟩���N�N'��������u�����V����a��ޏ�ݫ��N���c��=v�x����\�'������0��	��y�i�q�߯9�[x��'���͛�3�&�m�$/W.�;eGC�_���Q�x����;봘_{��ӵ�?�q�'q?�~��:L.�?8����!��G��~���|?|�:�	2���}�����;�������\�ޘ�?��/�D���o�3hi�څ^��r�v%�D!�5�5�BHj3�7�GkO^�0���ܔ&�W��=��U0w^�a�}�i�xm��&7)Ow�:�׺m��]AJK�˨j��Y��'��y��u��[-b��|v�u���ǐ��\R8no��/ꫳ{���A�N�<�7�������a��.��C���>'n:q+�����'�}q�W>F'~C�q>r?��N��~wo��޻�8���t�>�	��b ����Ŀ\�a���K���]F�C�����^�|@�'B뮱���M��n��c�¾�~Nx{�F��i���|�}v�u��C�;�����!r�븽�8��|x�g#�:�����G3!O���Z�!�s{�d������wΝ�ǉ�}C�����vQC���z?!�0�m����w���}v�s��N��?�����U?'��c�����t>��n+��]���I���Oo��T{��8̍FV%��c��p���S}w?]�N|�O�;��u���t�����x�Q�~s���]�@����7�`�v�O~p��z���Nw��8�]����O�~C�}]�R������6��4��ҏz��1��:C��V��e�<N�,t��'|q�����M���N�������t���<������������ۅ���{>y�)�v������1��=1S����/�gb�/���i���f�����=B�#f �T��{~C�wN�8�|��q!&�zܲ�|���:;v��N�|�ێ���o^�}�s�L+�~w�G���+�;Q~}�V�}��M�\|�L||{ܳ���D�\O��O�?z8�FL|& +o�����7��x�:��F'~~j�ǧw����x��|wg.�
�(�
=O�q0�c���n�����KUb��>��,�*+�~ȶ? ���sY�eI�}sSD��z(���b>郉����=v�����;@�O��?}���&��߼���\
o'�n'?X>�N�m��:N���w����3�����ٍj�5v\
����7�N1��1�1S�O�y܏�O�aN8�C�}��'����]{�$���8�yWz�8��?y�F:��/�v|�޶��ĝ��7�uݼv�n�����;\��~��ĝ�<�_����|��|:�6!�������!T��}�����.�w�9�o��8���P
o��8��~����N��޼���P�8�~�9�!���C����q�	�g���;L<��>�i��:H�xy�:���>į;�稞�v�Ֆk����:+cW�უ�k"�=���JZ�jB��)Α5jR*��ݝr�a;����hW�}w&.)�trJ�2��u�yRĽ�� ���kwk�9Fj�$z[��]�bf`fذ+r+T].�&�k�9>�K-�(�do+�r����E!�����v�I�|��G�t��Hn���;~N�۴���x��޺w���p�&��o���[��S;�������/#}��7��w��awn<N:*\�I�$\z�1���u�z�=�L}3;(�}�t���a���mӿ�&���en����}��Ѿ�����8;^��;��9�^G�n+�w����O]�{�_Ӵ��'����:W�o��Y^�Ӄ��}���وs���1_-�/�n��ڭ�>�R�]۵G� ��˸�*o�8��A� ��bw���y���S���������q����1һ������� �/���K��T��Ӣ�g=�ގ��s`N���ζ��v�o��z:v���=�I�BI���м�>�۾;H(z����t����M�q8���q\
o�8�}M���'��z���C�*~���T~]b=���~����z~������^tc�q������|C���o��?ˠ����@�y�ގ�N$��7�O�s�a_�w���7�$����v�:w��9(�;~t�r���ob�JQUdz8׫�o�e5����p)���=����1�{󾷩�<q�~N'����z�������;L*��y�]
��L?���;��7����i��[�|�� ~IS�k��B�yXƼ�tF��q>ȾM�(�莡;q]���e�I��^;봛�t���R�h8|N�ӟ�u��e~��ׅ{@���o��Җ>�0�{-��iW�oa]��U��q�.�
���<7T\`xX� ���P�s���U����q�R�Ͳu�El�Y�_ݗ�pϝ���kM՘O��W��Q֯���Hė�?7Үv��kQ�<�&�	gQ�vױ�W_��ḭ��m��jt���b��֫���80G=�x6�auo��� ��]t��W�&8�t>v�X�Æh����lzo��`}�.-�8�|�G
c��{�8���Q�ga�������]���$�3����.��^M�|�r��vA*b�ph��U��%8�+w��N��+��v U,}�p����9[��!�չ�u����M�2ҏWb�b�˽��|�r��9vDv 0e�sW�%����x��i�[Q~놮��R8S8�]­؜&�.�hc��
��Ү��x�k���n� 6��\�!���9N~�y��}G�������A3��k �*����#SIR�E��+�<�|8e/z_��VK]�b�.�|ԅ_j�����ќ�-O���Bd��Mҝ��WQ3��ˠ�QM�}n���O{&�O+}k�nk1��m����lȉs����w�-���Gƹ�?HY�B����o�Hy�*�`��Y�����Hv���I��â��g���PՀ�q�B~@���/�!7� v����ۀ��X�c!�DbO����u6���&�d������ *�n�=�����cNz�O��i��_�߰Nuv�e�|�6���I;�!3_:���d7���.Ȼtg�a�ź6+����q�a�"�Z�렫��l��|f�)s�.\�l�lB.ǎy�Z��q;5E��9)ń�ZΓ|�9:��`��}crQ�*Xk���7m<7c�Ǧǻ�t��<��f���{�L�������`k�v�2�^+�YF���f'�.w�ɸ�x0[��u�i)΢/�k!�oA���ձ�뵒�4	eù���O[:�l�2c��f|���l�����g�ʱ�*j��0�� {�u�V|��1~�!n�.N7=#��spF3�k���m�9r�_��wU��K8}�Z�	�'����-�e�U�T�q����~������{���ִ;Ո�f��9Ek�^���譺��-�f��|�j�γU�N�%�� �X|��|��1ݑ��Fue���@�:�i���=�c�2�r!N���;�.��u4#������ȗ2��Ӧ�׏>�|=���x�ۮ�:��L�b��|� �* �
�k}oǮ҇���������}^pf�bH�}�Hn���j)@[�
�>���4C s�*C���CuSm����������7�;V�iz'"�,���2�#�#
�N�ڹ_/��$�Su�p�O���h�6�;?8�s��;ބ:1L��s�����;2@ϵ�L�SZ�G<�L������j5�q\�%Fŋ������Q�e�\P��/Y��N��L6{{!7{2a�L
�P��t�Uc_�~:b�_Y:��y�;��)��)�������=��[���Y�T�������=宭yJ�ޛo�v��cqB�[�Ӈ���]�Z�<��/��h���@���h�H�����]:gU�S�������`�lǽ��$e�$;uP�w���2�W�ϣ�:�8�g��s��0�*�f�8�e�qӛa]��9�ˤ�A�v�c�֪�Aك��q�zw����ѫ�O�F��:�W���q���Sn�ڶ�%׏Ά/���4��X.���/+UA��u��]I�f�f�i]���}}%�ҀԽ�^�^����c@j� ��*3x��xqD��Z����=S5F�<������+1�z��ڼWgި�h�D�뺕�^D"�x�7nE��(}qV�*���T:zѻ@�)R�u42#�9ߦ�>u[���Ȇ��cX2�ʈ�Z�8hϷ�׎{+;�B<θ�v���C~QY�j��@z��=7���Cj��WY^Z<ﻒY���\mm*$�9�t��W�ꕍ��R��ԦVp�s�E�!�69@�#�t�k!��о�[�~�D�MjddW^�C�B�Ws��`�0Xh�V��3��ؙ��L�Nc_۷�e��Z�s}�D�!yw��,Tg2E]��xXy-|���,�v~�9v*w��}3���?eH��tz��(��Z����@ԭ�$��r�f�Wר���%�RV��|�.�祂Wع��x�L��y�Da�'(�F��%���fMv��j�Q�[��]�6Kիs|�=�U��WT�oE�+`ej��`Ye�%�Sѭ_$9b�E����<^�:��N���m�Fx��m}g�!����Q�
���6���N�dV�cX��v������y�dm���O:� �'�]�>�������r.�&��<F�k"�rH�!�hi��u�7�w!աH	.(�r���}�K�E#lS�bj�����0P�#Q�<��?�gRCC�ٴ���� vk���g�IqV=��2�K0w��ϝ ,�~y�Y�^�ߐ�/ 2>낎9S-�j�K�B�P�۔��wϹ�Us@���u+��4�����]��#���3�-�pz�}-3fT��D����f�qJNUu��w���ǒ�?�}iL?T
90�D���ʍ��!��z�S��	ax�JR��*�a�;�w����&\����{+o'>���4�7�Y%m���jF��64�,r��r�	��:n#�.AO0��s.�l������UnsR��){з�],凷�uĺ���9�r� �!0��,�Dt찚����^���C��}S��W��7�m�|T��iנµN��G\�Mz�V<�4�\�R���ڏ�糨�7ĉ�>�j5���J���ޤc�;m�Ng3*�3+ԗ%s���O@��Ɩ��P1�gg⽫E���Ot���{�~�ԽӲm��D�0�P�?�}�g�#�>~ݮ��Y�k���b�.��~����3y�l9�v��ú�	9��2j��<R{�+&Z~���[���c1�P/�{�
�Ô\`x_�}}/�P_1�P��,����~�nC�^;�@Ê���@=ύ��7垽��ͻ��{I4�l���=��C/�@K�E�=��s!ݙs���=�S��	:]|�x�*?�s󢫫���s����E^�T*�#��y���zp����^Cb1ڷ=�Y}'"F) s�O�M�g1:x:�Jx�2����C˴!ά�\Kb�+|�԰��)�g!I��G��8�/�;ܭ�fpv4��/��}h�]!!�ڭa�w��;9sćAu<	�P�����l��Ʀ�P���FU���p�j?�����TZ�R:`�vd�m_�.s[��É'�k�뮺�/��F��8@c���(��(�5.��o�\=�*���J'.���,K7K;��N@������C��%����~�]!Cƺ���㨄��ZyG��z}�M�o;1����ԺL�q�ەy�[.��:sg(�f�ua�N�.�7.
#�Y�p\�/���C�C���9�o6�X���1�;�L�ƀ�� ��z�1��"�ln���i.��2wf���K����rU�[	�RZ�r�8�1hR�׾�m�v�w;������9�q��W����<� �uX(���	�'�R)�h���X3ۨ��s����گo-!�8�dbO������L����^�N ��3�,�Ɂ��4�E�/
t4X��α�o��K���R'vD>*Қ�`�4&����k���I��Z3�b&MD�C95*a�7��@Q�Y/Ƃ�o�~s|����#5�J�4<; ���ӂC�]�7රMү��S���Oޅ�Cʘ��b2�n 
�y��A�^�le.�o�}�l����C���n��U�p�[����*�j�2q���c�]�o�36�@s��陨z�ڕbC�����Z׫�!>���^�c�Fh�{ޫ�����e�Ӄ��r��H�t�r��ZT�Qa�{�99��s�3ѝYC�X|,��ɥ~���q��o2��K��]S��q�Ћ�N�Y�ۑ�2�Иl}�Mu��g^�]���\H�=yA�WH�G%#��ڮ��wv�����S����{%�USҌ1�ꅺK�W�Ls��ԕ���9��\~�oV�����Ґ�i,g>�'VҪ��\/5�;S�]d']w}n򽋯�i�+�`o= q�\�8:""m��pg��5O���+�ʷY��"k�{H�=4SJ ��`h378U���T���v�-�ErH���.47���
WLAϨ��N�A��b��`0跀�U��w7����k��w���zq�l{<M٣2w�6t]������_O]K�gzs�5�۷0CW	����@�k�,�hv1i�^;.,��o���W銵�`Ŕxř8�GrPD��)�ev	�(G]o��-a��%u����a>V/���vJŮ�˞\V9���n�/%:r8o��A�@������&�qKl�Ly��HB�hؗ��L}����p�/b��[���������I<S�10 .�J�LZ�
�B%�|���;�ͬ��&U;ާb��# ��{=��sX�v�1w5��g˱mp��1݂�R�$��cHW�U�s��e�9�bK�A�y ׏�fɒ���Go<���n]�����:�S��
A����݌�%�����KP�_��%c0Q�����7c��Ob^�
�u��$2�gN󢼢;qUO��]+�GtNo�uT�U	��jU�kY7D�r�ʺi�]V��b�gm���e[T�GD�vlQת�|�z{V^��ښJ�ot�G���l{�ja��i�Mu���iǙ�r��:���so	�=01�L�!�6C�����o3m	�ƻ,j�Lڥ�����ؗ�쩱�V/�18mμ3}�s�w�y��!���
�g,��	��V6�\��!ݲC�����Z�V�}+�?V쮓&J8�U��L���U����� =���E�8���L<����'(*��J��97W?�����_�Ib܌�~�����#���%cA��1�h���H9頞�n����2�wS�b��[e�8�n���G���/l��*�����;��<l�3�)��k{���*�r5�yTl<�y�{��lU�I�^'Z~��o&|ҌA�6)^�w���-k�j�U�Ǝ��
�NWu'=KĂ�Ϝ�Q��H *�#���:�Y�Vk�g!f�̙Nj�N��
,�v�H�F��l�"%\�i�
�׻YB-o�
�NgCL+��ۏCs�x�%����h����٦3	�xW[��ɵ�C+� �.[�3�]��@��=��+ޤ���{	$�o7���Hbp:~���s�Ƨ��3;�뗎%��frr1v�����k��M`�Y�Rج���io��={.����%7ϯh�)�o�.�"�����&�e[2�����)�j�E\��ŋ���)��Ē���#�R��
,�:����F�G�Y�SsV���£�Y:�]��� �W2b����K
�Vf�}ﾣ����qS6V�ȒI˂�B(�PUx�s��J:��t�(E�fL���"9�sL"s��Z(�,�M)eh��#�B����gN� �qR�:V����ee9ǐ�!V-L���R�tS�8�
�S�$*�M'+q"dj.<�dHt-mdd�8��Np��A�J�i,$$�9	�)\�L�VFU���9��rd�<x��9\�0�I)��((��E'�.*K�����9�r�I��*1R�FV9qSP�QI��r�q���&9\9�4���\e�+C�ps�RQQm�I!��$I��94�Ց�HTX�#q%�:����$s0Բ-�K$̒��*�dR�JXr�QJ�VQ��!2L&�Ee��E�9uS�*��2R���U��dDu3
�R�

$�AVrΚ�s�3E:Z�t9b�d�UJ�E�Y��e��b��1��&t�T@;6;Bx���N�#��ֳ�������'�ٺ*�ٙ5'WԔ|��f2�u�GN�b�}
�睍��fx��!�������Ğ�* ����B�*��ܸ��ޙ��55���[����J��d�&����F�VgA��:�ϗ��ET�����3, ,7�p|�r�[��p�%���"���8�#����u�T?7u1p CYC����##˸Tk9T��5iHdSawP��/Q���!���67���F|�Ιϝd��m-���݌��F7��ϏL��b��2:{��Lg��v�
Xu��*�f{����=��wo��C}E*�\��C����A�]�x��Ћ���Ak"2J.�!]��nz���{R����\e�x(!�����j�Nu����/>�Pk�u��G��<��{��� \�+b��z���u�X>�Z@�ڼO:���]�~k�0a�S�`�C;�sͪY2o�.v�aC��\.�y�
��<^ϼ����yS�����r���Ӻ�6g��:<�=	%D������1��B�,gvs�%�Jy}�}�R��x7ƈz`6k�~�mm��Y"��ތ��v�D^u��/�u=���l��y��]��)���v���V���y����_=���!�K��e��1�|��KSI��8��e��BG��m�R8���ͩ]S�Wb��U(88nw-P�S9���\+��1i�t/�����36���4��Ġ��{w�hTEag!�B�,0"�ބ�|s�Y�v��H��L�g���vJq��a<���[����m\�S�L����_�Qa�ߞ[`ʝ�l���y��*pY�Y�V�*yD�`w_��a��O\b�|�L����b�_vw3������o,�:U�S��n�Z��<UQ\ྲྀ��eY#�y���P-�2���ǲ�z���߹�C��S+Jy��W]&,�Q��D)�uF�)������b�����E!�=���%oAbX��S'F.�9����,�r {��!w��o�-x���{�̸��ɋ��D<�]y<F�i������"P�'AN�c��o�:�(Ip�w[R4��,�H�R&l	`�u��j����S�!EƣfN�x؍��I��X+C�J�}�wzӓ^�Ɏ�����A�#讋_J�E��{����G��\qʔ�=w�
��&�)-į����=z=?C���Цc�j{:GG��gY�]Uxt�գm�4�S�+�@��WvY��96���ф V�;�7yiCjR��1����K�[�NϜJgk�%/V���=�I��f�����K�����L�S��jPa��{nu �]��]v�]j�[�6��QEn��%��]N��19Wք�舏�4�{x����v�L���_\&���%ә/~��&S� 9���g��� ������;Gr�S:�j�g��/-�m^XϧX�siә��%m�ñ��|i�n$|��{�%��N�1��w+&.���Okoj���ޗc� #�(1�H���1,{�a��u*�v��L<�bf.XU����߫���F���Z0�j�ey
.;,.k2(�K�iG��޹x� �q�-W�<�G'0�q;��"<��Nf��s��d9��f�Ҟ��]���ޓ��þ���vW<�O=�DyET�^�v������Yugl��fM�<cͰ��_��~��C�$8�FnT�q0�GԬ5C��d�z+�j佊dU�OT��ݷ�ɿ�p���T[�����uF\鬿�e��FR p��X���H\%j�xqд�a��FP�bRM�C��x|�n���:4�]e����ψ�)���V���c�$�=�PCc�u�ߍxeKT|]x��G�ı����]�e�jkzX����Ƣ��c�#�fqU��%���r�����kUc-��H̔*����`�u=��.! "\��R���Ʒ/%��(����j��G5�F�ʁM7��mC�lb��^!7X&�۴��3�S���N�E�/��+�/���X����D}}�>]��#A��6&�pQ3&@
f��b�8RC��u�1�[w����;��/Ay~!S�ˢ�Jx�{l"�~����FU�@�t|�H��C�R�LJw[���ۊy��;�2'�0���]:�n�5���"i��ġ�LJW5�@.����A�ԛ}�be1��f��u�s����m��vv���9(
��թ_���x��|�Pl�Kݓ�(鵪���/aƠ�62h��q����?x=�.���בs�|�y������B� >7�G]�Ǵ�^��J��;��}:kf��c�dH�I�}�����0,M��{�2UV�;{E���0L�I�����^13�E1��mv�c�~�A��Q�.7�FG�~��2���MR��Q�P� bh�G; �V����W0���z�]��B3F�͢Ә����(�Z�ݾ�ʬ۫�a��53��:��a�{�uZa;���f�z�)��2p�z���E����p�!�c�����\���}�.�������hzo��Sz�1�H-�	tv���B~3�-����j@UeLv� ��ڷ�m������z�"m}�.��Tū��s���e�}�c.L�s
n��fv-|uP'~�����x�K���$�������ߓR{Ғ/^��<��`��9a�ʮ�Qh���G�|v�V���޵>�X@[P�f�:�ڝYP���ՐZ�0lt�um�@9�֙4ޤ�8��r�)��2m?l�Йʩ���p� �ʢ�//�<�Ln�wPz�ц��s'U�΍4.\b�P*櫥�v]���8�hE�w����ȗ2��S���]Y���Za��IE(�O���c�[����* ��5.o�{1�c4�9O_�ס���I_\���<�)fVWN8d��md3�
�>���&X �
S5	uS����3[p�VM�ͥ�VT�\ԍr\7�Ѝ�S��924_��t-_���"�PFG�����;ffd�{g=�N1�C�����o ��y^�v��x��}T԰�	&Fm���ychl�ݴ�w������
$>�1�^�/�)�C`:ن��{{#y�9��q�ɣ"�[V�6h�ˁФ�=��9E}�/�[�K�z#����'Pf�@u��gS3J�CK}�{�ٓ,��O� ���޺�?�U���i���4�T�2=��#G�ڸ��͵k���U-�����\��#�B�@�>.�������D��N^)��5�r��]��H�6���;e����,�"�9����v�7����\l�����M���qU��a���VT5C��ͭ�ܴ	S���]�Zw4AsA�
cg��諭��B{$_�C"�K�2_��������4x��&��ǈ�Q��پCyeK[�g�ZTB�=�{V�v�eƣ�s�9�U'Nf��u���=��}LN�#�}�S��8���5K�¤wf��\#�zr"v��to®o��}�L;��]�)����$�bn�q��{=��ӛ[�q�Q�'�aGvs�%��N�hcYqY�z~TE�T���N/\���s�i���^����I���D�{�=�����蛞@�ɬ����]A�e�Ǳն�������1� ����T�nj� ::-\�Z:��ϸ\9�����n↔l�bt�{)u�V��+gL�5�����7F���Q-]D"tj$<�#i\��y�J�jgX!�/�Y�x+>�yЬ�g��`�C�2���".ۤ3L����\��o���d��8K�]a�d!�}��̘N[���8�s���Wd?_�ГWE�p�tO�a�Q���SP^o0��糂��g�繑Lg��%oF�R�vk���5����\� ���l,���\��:{n�æ�SR��%q�*] ��nkXb��Ț|�Ж%������:��c;Mz�v�vsXN�:�i��0dȥ���:�7��a�Dd��ϊT-���bڗܡ��n.��w\WI��7��:�f�a8�xv�����">�����e.K�R<�Eh�x��k��q�K�izI�UON�c��::��;C�n�\��;~�y�{R�Q|�Q�����I�0�4���!;l}7�H;��7�m��&�֊��tr��A�2+���cQ
��rb�:������~Kڵt��=DϽ��yE}��F���rώUW	�<���Q�|TGn�U޺	�
��~'#�����Ů�h�K�t��T��f��i[�K�2^�����J��v�H��u�I^o!��s:�V���l�H8YP�#{!�\"��6�,d�.n�3�쭼�v>�9��0K�en�������`q�o�f�#��s)Z�Q9�X��̻U��>��2H�Ҵ��x����	z%°W ���^�u�����S�M������)Ŗ��� ��;�y��u$�o�א���:!5xj*[+.��@!��z���s[[�1@:�����E_u���L?��;	�I:oH����a�3U�0?������~��m�xtT���b��Vb�w�u��>����/r�~�������9�Ǉ0��}�*z��������=�����䮉���%��'�t��p�����T����)�\h:�ܳ"�,�y)Ö����:�+�r�H�ٗ��Ҝ�����AVve4wOUW�U_f6�yQRf}�f�q:�<�qݶ;ae��q^�˷$@=�>7v��YΧ�4���q�Bn�3�x�;��A�73�b$���#C`N [�Om�TeΘ�����h����-��߯�ٕ�"���KB��u�n���8����fB��?9X��6#>v��o՗�zq՗N-(�'+��O�L��Վ��P�����5�*ة�J�԰���򞩖�ʂ�o3MYh�P����FHb�0&| �?�r�iR���+�_!�ab�x�����+�wUm�A�S��Fӟ���PTt0� ;���B��Hz�z%,+��ˎ�^K��Z�,ͳ~�o���/^�[����\\)��P�p�7K�c����ErpUx}�i�30�)8ȸ���N��)�ݠ>sr��ݫ�^>5�W�O������=S�̐��oQ�Zz�K��c�lԳ�7�4.;!G^E�=���(y���������j3�>�.�œ����>r%迆���[7��!�3�&��O��m\T�-����������@�PKϱ݆��6(�WY]�o^52'Pv�y;����P	G8�m&��S�]������w�����k=�{d.Wc@C���~�.�Z��Q�R��e�\H ��2ie8=~3���rp�*7S��Tv��^�C�9�H�mnjv����������g�[�6�}�0P�5:�˜�A���b>��!���S��0TF�pe#�fm�w��s��C>X<V*�^���{IÔ%�D=��'D{]Nt#c6e��8�C>�x�yB�{k47�{WW����y��o��6jwnp?! H�ϝH���^�s�' ᪽���7h�!?�v��uJ�1[	�b2!������[B��s�e�yv,Q*�^��b�J��(����	�5 U�9�N��l>ǵū3����B,��Sx�Y`+@q��kş� �D4'��S,0TXg���N:3��t]%C��RNӌ�:���_��*'�Q:&m����#O'������l���n⯞d��ɮ�k�(���m��pEi?q�*+�#j	iL#�u����ơ�������<�����\���w�'�aZ��2���C;�b)
�||I�E@���U!���!�3h�Vr�h��\:+�Y:�0�'����ls����.���$T*v��PYf��gw-ƭ^�_����#��"�YOr9b�wLjW,eté[���������N(;���v3���y��k������5�YJ��ݘTd�
`.���MX��ۗ56q��pV�c��h�9kN�ޅ���[ y��OrSO�W�}�U.����{�P3�;<��gS7a��3�߸��O>M�����H�[F�2:��M3��ZXe#s2�?�O�6dt�B��	�"��E�pS���[0�؀��F&�b���k� �{�b���+f���pT��	���/�[�G� ���S��D�u�T�m�����n9а��P� u�Đ�����w��<�U���i���4��#����=�)�Tf�C�傆7Q�%\dpl�r��y�1}����)ΰ^8���2��U�G]�s������qۙ�Kn���<��^]��Ɓz�O:�u��>v�9u�Ik��9u�!����;���׆�o®����^u`�sʘl�˭�[+�߱c�@x�'���;9���^�C>Q�8z��wa�;%����CYq[��:[V�7�zq��8pr��^R��,��:�Y{w� ]�#�9UՖ7<��D(����s����Sefw��u�Uޓ�����{�h�n4���W�u;xU�x�+�w�hp�Z=j�Z�b�F4d����T>q`����:`D�YRC`ä �@�Tא�7����O�M`ʋ��W]�T��a*��t��9h)p؅��֣�)6yC�
H�hҏU�N��@Q#��(R���M]�b��ji��-�f1�]I�ϴ�zmƅ���z�.�z�9+�[��}�&�8�Z���GJ�i���t�^(3��v��Fn�Wmb�2�8Ƽ2*��\ʺeS��%2)��
I��s�yY�����5��#���c�ь]S���O�Bv.�K���
��:���n�eT�v]	COWQ"�h[�o�uL;YE(��R���c1*q�z6fw<�m��͚l��{!�����pr%�ꙸ�rʺ|Fo�����g�2�1K�n���;�;�w��DMr$P���胒�W��j������M�Y�,�"��IՙH�%��h���Ó���,Օq�8�m�h��]������͌8�R����:��N�A�T՛ږ�O��5T���5��Q�
�N9f,��,M�BH����V�5��<G����=�����`Jh��8������'���:�2$7��X1bI-}���eʎ��&CtpˁQ�27#uq�\zͻ*.��6Ŷ��@����]�� 4C(�!�#W]CQ�Uv�/�87�Q�k7N��-5�q�㘰܇m��4�[�h�g�G���P_h�� n���Þ����I|��/��=l�����|�A��l�jṀ�*T[��k�1��dևg�M�����Rl�pvk�{� r��KQ9^�RWx���6�p�;)�rc7�Q�sHd�q�;�[+�罊��786��X�ˤ��w��׬��9,��ap�"�/��la�/&9�̏Fև��jC���o����(����Y�q%ta;��9�o�o
ʔ~�\H�u��)�n��E�iph�B[yz-f�Z�`�o+��))�����X���MF��Z�Ţ�����IL��+^�3]]*�,��E�+,=k@.b|�tN���s�'q�b��A�*·�=`tYGrӋ)oc�B޷$��^phg��%p�B|%�ۛ��Ml�ì�Tm%��gm���`���	���	�&ų��u�ȹe)Wt���z��L�������Cܙ�u�';Ě��Qɳ1b�-sXMqtˎ�O�D���~w�	�&��|g8�ۂh�����̝�{�I���(���Ʒ?\��c��x���\�gk����n^�T��֚T�����v��O)�C.�u���tޝ���aO��vUx�;��[&Ec��9���%gQ��^��d��y������5n�R��4�+r�v!�q`,FԚ�J�Cn�<�%�7�֙V"�{	K��-��X']vӨ�+Ա���P�=�2.8��cz{!KV:}��A44�� a79ǣ�T�\d��lTE�-v�N=����O޾w��w����p���1��4,�S!EX���"� �U%b�dHY"�t �$��:gU�)��D��)4�V�êI�ND�QUETb�B5�VQ%i"EY�hUE��B�	$!E���e	��T��h�I2Tm:�d���a��XB²�9Ef\�#L����f���%Qr���3K*�"�آmISi�j�V(��#�F�#�TdQQk(��)kU(�*�	�m*4��3fIY�S���fEUfȌ,J�R��2�I6���h�Lε��hf�m$�QT��R��f\-P�)�9�E�����4�9&�ˢ��M,���9H�L)U%FHUl��-4TE9�Z���XU�iҒ�:a��	EӡG39"Fi�E�fT%Zh `��H8:�v�(sl^6��{�rօ�W֍���'�A�\����BƘ�����s\�z;7�ӎ$3 |���5?������=��O������Ht����H�ђ41PW���V�)�Y�1]�ﳫ}ZjxZ<�"�Rzz���
��N�^>��⯍:��Cvh
�_�����sG�,_TUv��`��˔ë#��v~�N�aw�7�;�8�s��ei����"��N}9@��� I��r�2�e�VuD����-�ʴC幑Lg��*x;��X��w2�k4'J��E�����o�{ӹ�M�Pjt� �U�Z*C:k��Rj�s�$�S�u3��IG�yoVΛ}!���a^�����y�T��7�
L)�1�F̝�OKy
)1����;\��Ϧ�7�8���[=���Pq#"��эD���8��'�g���5���q���ϒ�,���wb�;X�#
}�\Q��wMT�GD]�C�g���7΢Av���p�+�P�q�Ԯj�\�ꯜ4�������e���y���'X(M.uA维��V��P�;�b���s��:ڼ���L����3��J���x>���Q�ʷ���k@_]�Qk�j�H�� >ɼŝ��ܚ�~b�u��R����ņ7x��(?����I��m�IY�t^�`�d5G�zV��:�MLN��!P�W�Lu�޸�̝ȣ&�*�g��Y:�㨸pw�5Dt��s3qDD}}ճ�7I �U�����7kԁ�G<ǠNe+ڥ�n��E�˵Q�>�͛꽋%UY�ob�����Y�u�k�r[�EXw�ƙ��c���y�~53+�)F�}����(_��)��NĆS�/|�Mc+y�
6Y_h�2���by�T�T)����m9�f��ƝT�۶��74�����B��w\��N�Iߍ��*�)����}0ȗ�g
�S��vV�}:��)^!N�v秦q�,T�X�}9������d,���n5��O�U��ʚ�rV��F��9���dſ���f�Z�ws���x��.�c��|<7)[���2�S25�%󝊿/v�o�}%����#jaɪHC���v�o�>r�#^Cb2�s�Pp�%�U4�73S�Z]q�;`B����3�-����ae@b����_%��.��EH�<k J.m���Y!D��޽wXS���}�%�0)���&�RC�]w�o���-�֥����r�g���V�/O<Hw���9�����)��F]D�T|�"��/R�E��������}�و���X6)�V���kN�dK]8ë��+>�Z��{"<y	��)��J�>Î��U�c��(V����u����3������ڶ��{�X�jE�p�Xp� �1�sr�`9%ǢٚJ��Z������Y WYg+���������r���j�*b�iOO��Y�N���@�����~PЅq$t�IWV����#3/|���)���Kkו�҆��s���T@�.rP���v�+� ��ɦ��%˦�I�pBj����9M{	g�n9�q�T:vd=�v�g�L]ߣW*���K�~i��,�Wm�}/�f椱�H��I�|ڨ�+i04= ��Ȓ1���EK�r�v���a%r�N�₝��a��8��{�!��5<���ق��7ވ��٪ݲ!�{J&�"��e�M��j�]X#��{qi5�\�Y�~�j�í-����p6�I��흄]I��_Q�V��͚�fq?zQ�C���΍]Nd�a��v{�� d���̞�p��9���
��ݵ�}�.�2!�,qh'
ܭ�r�^^#�#Y��:��1a3�:i-�}��xޟ��/��g��I3	n���a��yXx+���.S�|N����0��p���*�����ߢ$b���a8^r}�=1e�2��)��W#�\���=,�-� �ͧ���_���ܤ�5�%��o��^b�@A�v�|sk�y�Ke��I�����Ԅ����,{F�����t��n*�r|���%��w�Cc����}�R�O&��U&Y�^�菾���t��n�s	z:㦣:�|�4_�-���U� �nO?�˧#j�U6�WT��Vr'RW�U3F��͖���}�Ei�TdS�D��
��k}oǮ҇26�4b�}*϶y������0��a8��p�N�s(u�n�ݐM���(���rZ��L��B�1�Eg����|o��"R㵈��s���blS�v�:0h6_>u�-_M�C�z]lZ���;8��z���D�֡�L�VC��g�dw'fH�����v�����e�s�=��$�4{Hs��$ȕ���F���q"��u}\��6��lh{{"�vN�ݵ��?����1��=\�Q^H���_��hBx��A��Rc#�:���;n�n��%�Z�e�{����=��zL��?�'A�*�UޮV1E^X����dCL=Y���4�ͮ^T��b��	�b���#�J�ȿ�����! c�ݲ}f��V>����z�щ�r�[�%!xj����$�lA�"^�^]���n�_S �N�"��ّ�p�fW���� (z�# �����5,�Zi���k�z���-껱wǑ�g^ԨsN�e
YB,�UZOi� �M���r��b��}�V;���R�ou�1q�@��\�W�X��MC�t��:�Qڸ�̏�
hk���U�k�gﾏ�����]���vV��J�F<�0��sӓ��䪧1�M�/����x��B�ug �j��Nc� �/�4�g���Eu�͞��u�r��>uZ���Ʋ�_ D��:k�o	�w�z?}]����@p���z�VE��G�!<";9bՖ��y{�/�۬׶����%`פ�ć�hW���G]%0��O���\cܲ����;���-n��.r`��3h��k�l�#w��z2F���<T��
D�W�$�9�Er�2VP��˹B��$���}.�����N�;�<���o�}s,�	Fi���Ѥ��:aC(��l�Ĥ�V�S��;�Z̘[�t�s��;��V����"��NB�8��4���N/=�w�f�(�Nq�V�K.�V�*x8��#�5���Н�X�}Q�%m�G��o;����� y?��T5�W��2�FŦ�+*��0*�'�2�ں+����1�V��E��)�H]@q��BR?��<`��kx���q[��le{�IY�m�g�1o�Fm��ff<_pK؆kpX�P*��s���5�^�4Tvt�+���H��6�Y{P��8qS��W������W[�� u�j'���SX���*��A���{dW7*�W,�scv[�BE�dz��I�-�'������$g��xf�`�H�E��f-7p7�7
�!j��k�~y��ͯZ�)V� ��T�ku�-���SUճ��>���*vk�UW	�<��QGI��Dv�U޺��3�F{Si�B����5�<����4H�ȎV��sYR����i[�s%�^�n�{h]c�|�I;�J���h{��� ���r���C�G+ְ�5.�7��[W�2'X�sp�9�bV�O3�j�a���U�ਫ਼Z�^� n$}�/ᵒs�w�3���l��+�a�����,-B�d����b&y��/%����,�5B�ӻ"[������3���Ry<3�]{��������ͬ���ָ"��&�����F�
�n����uù�*� �Էs�N��x�k���x��veA���ׅg��zy1����g��7�ʨ
�.�wQ���{4��_"W3ӑ��k��N��<�Ϸ}�� jW��qTD�.�N��$Lq1��x�/�fzcP�;�Ƀ�:�!!���o��W]}��xnR����]r�O�,=/���GS�N��f��r��������״�|��Χ�6��'!��)��]��w����<�б�2^��1S�Z8�4>=��s�Ώf���V�>��X�Y�%����
�Q��7�!kX�&�y�G��g��'Wad��_�������>ծ�igAU7茦 B�. R��:��
$!q�fB��>r�#^Cb��A�ܤ]���i�(�P��/�XD�p�+��w�]S#�"�ة����AWg����9�J�7Il�)f+Р�!���3R��l�6uiyg�Ҏ;��i-�\=���[��O)�sm����<��c�)�o]�u<}N~�t��ܣ�;��it��(y���-��}(�oDU�2%���E�ۡ�~��^^*w�`9��)��}4*Òɜ��%�yW�_lB�#QSIKf^}/��9��Z���ړ�ڍl�g��r8��y՛G�����䋣	�/"[�b29�7ҷs1j=�9��q����OW�
���@]�qe�����6���6�Ί�]���ik�wum�z�*P׆g��^|嬫-W�uc���zwS"b�zw3�8x���������p�����o��e�958����20T��ݖ��:d��m��k#U��m7JYĮNVon,�s^��XB�epz�7�g�y��GI<�v��w�
� k����J�Y*7��1c�L,[�t��!�w����A��hu34ݬ��W3)r�S�Z�WSf؎5P݈˚�c3�}��W����.Q�d�>�sW�x�O˜��luחn�$�OP~��Q��X\�]��#}Mp�t���sO(��e�B�|�|ʏMH�+>> �^�gn����E) ���PF�xh=�^O[5}+G{T�IfoD�K�/kW^4+çʟ��Ƽ�Dݖ��*G�wW�Z��'�+���E��2r��Dy���1ξ�
�WjH���#�}v���Z�n{J}���؊"YyՈ浚z��gB;��]'��{��g���4=��\����^�C�����C��{u6�g8kr5���4��q7&��4_F�vc�rZꁸ�r�el���7a�7��$�"֎��fv�%q7+s�j��a6K������|Z�I�L��L��Z�o��M�s��nAJ�#�f����������J����݄8�#z
id�����˩���D���.F��R��Mz�X�Q�;x<��]�����E*v�ߋ+�$k�-˵\'^�9xCKw
�R��|��6�,`Q��x��w�3���G�������b�uv�WgHj4'���eO2��lS���ҟGi��Yjc�(9�Sr&o������8�����g%�K�.�c:}���b�Bg:
G��L�'�v�W�Y�;:ހ }^$�*��K��a\y5}3;s�yK�����%Ҫ��A�;կ(��v�jBKA�U��z�,JC;�ǌ���u$��m�<���_s�4T�D�뗘~�ƌu�/���{��z}�E3�m�dF��j�$��up���^���D�s���i�As�]�����ۙ��o�o��/����T�|�ã��u�{u�i�T��^�.�o]���8��;���f�l�����@=�+��	&�eM��-fkV⑊���^��2ϧv���'ڮ"����>�����)�35�=�I,�U�]^�K��rD����.wl,���niC+����ˊMV�Q�h�7�>v�3ZF�Gml�=�XS	�H;��h��9��s���]]cU���Bm�v_d@���ڙ�k����<�C�3e�C�vҲ5��p�Q�� ��ju�k���Π�x#gk;T@sǇw�ה��-�"˽����z6٫�InIbmG/��-j\��s�
�����آ�������>�ڼD���W�f�r�j���ՀY]����}������m7'x���#��Ѯ�Ѯ17���ou����/��q��� �	:���炿���}<���κI+��S|/���.���>�Ν�����k����qF������_�����������&A�6JT��1�a����Y�y�J�}���A�\�7�]Ȭ�!=;�O]�$N��E�y�<�NU��N^r[/vm7;p�2�%s�f�"\E�ΧV�_;t��YpQk%�/"^)Y�)RBr��5��Q��ϥ��/��U�Y]Y[�h;l�\4����+�N��.w-����^{��ji�{q;����ʹ��yu�/^6���t��c��q�a����zIe/r"�޷�|������wvM��������x%�[�w��M�+/�Tu?��ۆ��9���&��F7P��+G�S��^�2����ܵ�W`�׬�uZ� 0gV�o��$�,�{}'ARùd������'�+3(H�^��Yrؔ�{/z��L���L��cO�+��L�ߊ<�\�#)8��]V)���|C�aL�.�Iu�6�܉ e�*o�����|iq�ԗ �H�<��=)�� ����B�L����Kw��G��n��]�d��je����s�R"
�1�F���գ�k�$-�[u):&#{طU�&AX���htÜt.�ɓQ{(i��z�w���2�f�F����.Tꆾ�AG��n=���gڒkm4q&��ě���,��:C.�f �����%�u�ȓ�x�,��f�A�e�q�����]k�U�7C��\�]7(n����;�<<��+fv+�%�y�	�g��E<k�5y�Ё����@��K�vn`-_�M���fY�N�F����#Z%���J��'�q ���\���貺�dC���,��z����9�"��֡0N��*�)���s��	�e��~��nM@;`<�-{��)�.��ޏ�M�79�g/k����� �;[:����a�=^0��!�5�G�;�wu�<���S\�%��ӦK�L������C���}�y�v=�6/(�ݓon��&LWbU�t��I��@#������?ڷ��M�����z^3Lst����זc��\�y�w�sE�Yj@u%gw�q@�,���ߔW�7Kj���A�YC����f*��.�M�C�<���kh��v�Q)w���o!�����a`��1��R��{����ͯ��� D�|lD��e�A�����[�.s�,7�={	M��
hs����~�'3�eŰ��S�a�\&gH�f�ާ��1�tr�&p�ݮyy�Tۀ-D���x�mؓKD����Rb��,w;{��\2	��1�z
/�{c� �aIv��$s@:ӹ:���F;r���ɥ95������u��i6��H��a^:2aUh^�!Q's`�Ynt�r��5K�*_<��z�M@(��V���[�7��rjr>��!>ʣ����]WjX����y�Y��o��ԟ^h<���7�	�)���ۑTB>A^Z�7u�1����;�5�y�Ϝ��'5HY�Y���x�4�y�U��euo���5��%Ql��)�V֖A��>۸kK�+ӓxt��uls.G܃O��0��9��MĨK9b�&q�b�ʱ4�%J���6䠵��fmK*d�f�
���ע�㥲���7AV���]�ˠ���ojq_5l�øMt@g2�iFf��v�q���ʔ����8@�E�G�c��\���	��c��&�8sE"�8���c�N��
M��W]�g��n&��1�te��p6���I�������{�F �pS�e����Bo&��t1��l��v鉺Κx��ܚ}��.q�{�	�>��#���$�XQ�58�ʮ��e�UP��.��ڲ"�4M�$��
B�$bEa������S�²��BV[D�DSf����p�U*5dd���&u��]#��QJ�g:�e�VVA��-"����HEYPXF�"�RE6��L���D���Pl�I��,�+(��Vduf�a�B��24�V:(����Y�⤡)Aj��TjtV�d�M#�	��QB��-X��JΖ�s���R�J�VZt�b�i*�̤#3,�%��L0�E�ȱ4��iI�A����CP �J""ԫ�F��U����H��L�Zh��4�&I��2e��Ȩ��u"%��a��lH��u�QC-�\�i�2BTLΠ�1%�T�Nʑ0��rȤ�(к1"HJ�LCP�4���R�C�B�Q*�)I%�\�L�UY]uwU��S�LnlR����fW@٭LQ�]mêBB��;ζq7�m��6�L8��6A�Q9Gd e^�aQtEnI��}��}��8Z��qu���ӂ�44�����S���uoՕ����T��dm�dݠyJk�V�/Qnv�)����<;��YGc{�v�y=�-'s1ҧ �=:��
,d+-�=����5P�����Yg/Ʀ��K�.~����W<��*���ZǤIzZ��6q�}��������f�(��C-���7�j��/���Z�z��$sG�w��=�4ܙ�đ{�~]�$%^���q����s=A@�U��OVXa�#%'�Tev��S�h��y�姦�p��+�ZW�ܚ���@_�}�$h�!���V���n)*�Ew1-��֎�8޸��o�t���?1�j;E����k�h�zB�����1��S&[IDK�]��t�7;q��%e^�v�mg9��G�%H�I��Er�GQAM,�l�ȗ�9�eL�������ެ��v�`�)��̑���wu3�F�����Ҧ=	��G�[}r�����ʍnhW�>/�ȡ`l�.P�ӡu�DT5Ct�7��IJ��B�d>U�{��wRf�렳w�syf@c����dV��΍MN����B��*G����>�e�����Ѓ������՛G�����.�{��M��!aj��I�pt��5]h
*z�Bw'*�����֋�ϯTd�̧;�R��)�Tj�f��sRs}d*�5�c�˳9�L������ֳ1c1��6�2���y��n�!s�OT�����a���r�s���;ќQ��{���7���[�3���׏>*�g˞_��t˟�%�l�<$�*�8��o�m��aVMۖ��b뉣����h��Y_v}��11z���H۫;����A�9���.�+n&�����ᤉv�@.�d:��-���<�������W�q��=��T��枹^�C}Q��޼mx��_/y9�nv.���ϵ�k����:pG��cּ�k�d���ߘ��E;�D�,�?�s�p���9�;O�_Q��L�}@�YGe���TOq��Ib�/�̮���10R�!���>�+|ȄV�w���]>X���9�ݼ�g$�*� T1�e�={�TY{2��cV�C2��O�^�]� �}�'Bw\�-��6����Ӆ-� ��M�挽Ɯ5�g13e)\��6�&g����#M�Uł5�
��sZ�uɽ?s��5���4�>��ܚ.d��3��F�Y�n�Z�J�ɕa��pI�x�.q�c3��)�zh�����Y��\�]#�S%���Z�C�O0��y��ϟ��Z<�����wY�~�s���V�r��_FML�f@��am9�/v&�
k�� й'�}�u�u���{vSy튄%	l��f�G�؞͗�����w}�$���NF��U6̸v嘕�J��=Q �����-��N������Xk�vd�׻c�3ǹ0�6n�NE��+��bk⧲���[&��ұF���tY=�\v�udo.�oN�c�N!7�۾z'���
��5�|U�fmĦcuu�O������AT�B��C��o^�BaUv�M�����#��`�nv�p���WX�����<���e�*��Pk)�̞j�v9Z�M�����]���1��T��[��u��wt��s�`ۿ�{^�[�HX���+�훷]a&�l�)�V�C'-3c����q9Yk�MW=y�WU�(& �[Y2��0p�B�7&����9�-y�u/(�����{菾��X[��ގ�}����ڈ>C.�v]�O�]em�IϧT5[<5�u�.M;�����i2�O{���9����T����u AG��l���x9A�݄�77�!�}����DvK�B쎬�vk�SV�k�,�u[�dO;[-���Bm�v_g��SD=��n�:xWvl��jy��ۮr_]*����f�}7�����4�M�=ݨ��-{�����8���fV�P"YWt�Ֆ�|%'��p�s���\'5����'����R�~�%e���τ�Urz��$��3U��n�$�mrz��0{���q=��q�q�ۏK&�����z�#G癚h��=R�6mrwN8���?��9�m,���<�M�8tD$g���T�$tF�u�v�� �M*u�{~a��du�E��l�X��+β(UWw*��H�D�փ��zL����
��dH�&�Ew�tl�1qQ�	r弯{��-��"wvq�������Pn`dc�ۼ��)1�6�I��ɽ���}��A����G7�BB�9�(�n+�/�\o��\7PYy �g�
�n�X]Uy�/��}K��m�H��D�����-����4f������%d8����!ļ�S/w���Ƒ����w]ʀ�wh��ˮ!��Tak�H�akf��3�Us�<�� $�k�%e�x&�#S��l��Ov�6�3�j�Pٹ��)��^ݶ��9�YE�U=�����)o>���M���{�����z*&��f�'��ϻ�33�)G�G�o�p��_vЃ�]b-���O�C��u�Ma�\���/!U�~w��Bw�j�YT|Go�_s�O3�f�U���,��Y[sJ	��Qc!Yn]7��z}
���}�}�r���."N梶3�j�43��[���l��zD���Ux�a�v��n�T�S�mE(�����o��G�C�����F:�a���i؋��@Y�q7�ov�+qF��C�� =���FQ�{��jOd�}F�G��7���7��-z�%��+�dͣ+:1W7��׸���p1m|�)4�w�:=rս¦�4fP�����G_�L���h%]#��Q]�R��4E�ox�O���Җ:�ڢ��2�J
C�a �LH�!��TXo�}��f�YW��IB����p�k�����ZQRr�ʋ�%��nj�ɬ�W����b�\�!����o�gվ��W�~R?�w�����D��<���Z�[�S��d����^r�O�n1�����Q���X��{���N3�'�|��E���QSID�e�S�TW��'JlY:���ҵm����`�r<�zes�H�S��hu��T�I���fly��1[�6�]xʛ �r�U��{qG_�n#��+���Jx�י��g-��^�t�9���y�TG<EOWӇ�^+����]Y�7.��H�:�⽤��y�5k�'}��:z�o|��<�x��:^�͟�F��V��ĸn���n�Odo7q�x��g���OӼ�/#�	��{��	����Ff����7�c��il��7y�|ƦZƯ��M����������Y��:�`P��*@���oP��죯&_(2���Q��ө�e+�Վ��Q����g]�:.ӄz����Y}wˁ0k��v�o���=>�F��I�`�U����:Ƹ&	�P����:�;^&&��P�q�}�����gyo����}�2�ݸ�r��u����rrvQq�x�����m�k�{Rs��{�Ͷi��Q��xC�Y��[+җ�k�xEX�X�m�:N��j�\���l<~f��#^/
#�]���V�����.�1�.�bQHʡ���O���8kq6�S��^��<��5[;�T�b����W�|�Z-�\��wa�u|���nk���i�@���)={|jq��3��j�#�"z���ϊ���o�����r�q�q��ՈF8&�'w����F��T��r��.��8�a:��'%k=LL�8)iɶ���Nt�*uc��^@ު�G�̆oc�(���u�����;X��s؋ؗ�7	��v�D�y&ڰ'�m=�-��u��(���A�⒮�i#��˫�ٗ����Y
�(WA��{�m��yBҢ�Ҟ���ޜ�W�w���Y�Y���|�*�:�c����r�}��-u��,C��"��T������)�X��NE�Z[�K���'\�:�ԙ��)�CE�Њ)uk�-Y]A���f�N�#��n�{Jn����YvuB=���;��þN�f�{��]qɇ6n�NE�͸�+"��bk⧮�x��\wb+ΐ����^1q>��pq�Ͳ��yu���ϒwW\:���/o�SV����=c�Sc�W�k�&�YJ�Hy��g����"
�r8to.8$��c�-�ݸ�b�s��7b�L�D�q�����s���^���ػ���2����K��q�~�-�.wl<����������V�J���+g7�;[��I~�ڣ3ѷ���Or�fvkz�n����#{ֹ�4cVD�q��(�+�m�B�݋u�ص,�n*��KQ�ݮ��R�"�'���W��,�v�Csq��M���υ�wʒ��j�gz�gA�L�D��tj���ٳ�7��k��\-3q�T���a��F�)G�x��������/Z�g������ChI���tD��L6��Z��0�P�ɛ�p�M�{�w����9�U�{��bx�=]�[WP�q�C;�g�Y,�y�GXYu�^�m��&EL-"S{L(���vP��6l�X�5k���=O{	��χ<U|��}M���[�؆��L^x��{����2_rM6�guTV�0w�����+�nM����O�$����A֧�ļ�{w�{0��9A��<�x�jq���wΐ�%Q������<�56�R<�
�5D|G�I��Y���^��nv�1P���$�JxU��ᚧp�ۨz����_l|�wk#�
-dKf^K�+"%�R�I�੮70^n�<��M���Oeί�z�	O��ٺ�I9y�s��7=v��6�/>�z��Z/<�U��/(.�Ȉ�/�yiE�Ȇ��:	w�O6ų�ouTm^liq/.��������C/�/f<s}ٽ6z�09�u���;�*{K�F�>p����ko��<bq��q�zO׵uK;Sz�:��ң�S��^u����|S��44���x2�9N�3=i����;�1!�_S<7_ԩ��M��A����-λ�r����a��ߴ���^�~�_fd���$��S�y��t��Y����Jƛh�*K=�-�(W-f����,����������3%�V鎧�m�A����"m�BDV�쬹Wn�H7�8Ȱ*�F+C��sd}xc���f�z"Ff\�ҍޒ06�!�UUR7�k�A=���N�+o��N����8�ȅg�Z�81���lb��X�%ZUw8�_֤��<����V��Hլ{�Y���R)W�0��d��\:����{:�gk�������s=%Ę��d�t��{3~�'��m�x���UFL�{�l�#Sڽ��]��>�M7^�
w����Q3Lp��m�g_��u�+�ZW7&���|]���=j�Z,��!��|����1��V�w�q�q��ۤ�nVb]����rq#K�<�r/�{�Mr�s�ϠOk����Y/9r{�~��@��#6�g������=�}�}V�ߖ[�}���Ȗ̶�^+����yN����ʱ�/�/bͱH0o萕�H�Gk�N��ϕ2x���^+;˧]W]^i��[�y��dR�=R�r�+���B�#n���]�p�IC^WjYJ
7�R��	�U,�#z�8&S��4�o��5�[+ ��k*���]�V|�{��l�`��o�mIw%ٵ�WQ�6������x�vOCG%'���:V�ȕf����սΕ�BQ�-�H1���������$7�u�}ox��~�sn��g����</bɇ4�ًp93�s�iM�dx�\�v�o#�[���s/�ȹm��#�X܄�=�K��:��]���<�ʆ�WJL��"{�=��W��&=���
���Y7���vU<%�/gm��c��J0vv�[N�,@����&m7G��������C�+ʶ�OjO�ʳm�[��E��?��e��c�5�O[a�gQ����M��d�b����n��WF�OgmYx:{�a�����	0�1��.�9��\�j%����K+�f���&��u�wEL �IU������Wå�9:�1u�� 4�[�܏6�-=��ŝ��f��q'R�m��5��j#�+� 9%�ݜaY����|��BD����u,N�\ׯm0�
�^>���,���N>�媼���i���4�7��GZ�*�� | ����ZdW��gsҳ��t�>���P�7�v�[��&-	��HF�1�m��> ��u�@�w�j���n��@�أs�VEo	v�̍U�t����}�`~��&�K_�0�<)����;���x]�:L����A�/��a�ͮ@m�bB.���[3[f[���[J�Xo�'l�fխ),�bN�8�<u]��NHW(����v�s:U1`��[��o�P>Ėqv�u4�L��W4��ʚ�ՍSO2�m,U6�Y�
ݧ&�S��R��N�q�ȐS.r���il��E��=	���K��k�}��59�����o{�;%��lo)|���v��Eb����%gU��Shd����[u��������T5莑�b�ת���=z�=��Ddp�U*�qt,�i�����0�1�������Z��N|�M�;�&���gu�v�&�s)�O"�t�6`��+��p�zt��B��蹎D�5͢M��8��5�8�T��k&V��]�U��u�ʱڧ�^��ݬS���&�Fv�Q�d8wnJ�
���`=^+�SJ��0���1�Q3b��Kp���z�1&w�?33�է�hۋ�8br����-6�T�N����ό�}/��I���.*X�x�q��,���Qb�F۬:����l]7�)Y��uJ��xʣͱ�7��T!<�vO��:wz���/&�lw>���4�%<'����l���?��חV�v�� �7H�z��K4��r�<�i�,�����M���T�p���������+�mLK��˰h�3된�b�"���X1�'�$$C��I'5�����U�l��2f�̦�^�G|ƈ3!���y�C�"��N����(̡
�e&����*MH鳗3�U3�&ʐ�
+�iZ�%�a��ip�ʌ�եkQDK��Y,�B��H��6X�J%J'*�ԒZih�Ar�!
�LY�5.�У"IE"H�Ù�����h$Uȍb5�Uj%a!�4���4M �$���9�H��UKK��ZG�*�&�:aT�K9Eb�U����������E�J�Ȯt�es�R®hA�R�J�!�D+:jQb�����"���H�Läb!&\�0���E��H��FlI"���*R�6��9�5���C,J&����˙���hRBh��
.$�@\L�(��
��p�jW��U�Q��L0ÜSB�,�mB"dTUE�U"AG�DFd]��A�6-��Ɨf��g���} ��+�h�sr�.�����S�m��8���Qy���(Q��ho�.o\����;����;�:[UF�4��e
����*z�\KĂ��%�䆭�Y��o-(�$�i�s�V�@�on���r^�з�W���'^��Ӻ{�mt�F�w��>*���[���O�o*�n�|���Nag����v[��wX��ê2�6��1�&Z@h�6A"��o+qIEV�Yb��\��YQ,��v&���:�
2�m+:��W��%��75-��~��{Ѳ���~���XOs��l�L�l�@!���R+�(�d�J<���6q��v�QDv�l�V�V���+���oŚ�J���TvR���M��="�U4C߶]�ͥ�]n^�
�l���3%�\;���0+V���}�G8kr5����m&k��oN�ؔ�G�ۍS=@��$���I��;���JO�y�8�#�����&r&�\:�'Vt�7v�x�8����d��[3q��x�~����Ϗ���Ӯ���4iz�TH��T��I����N�}�� �-Dֺ��P�4��SU�f�����I�3 
�b�Ff�9B�R�1����,Y87��u5���PS�Wޞ�d3׎��D���|���W"�����!��2.2w�:H���w���gjZ�[ۡ�_�1�C ��H��2hza{��犷j`TJ)]ɳ����o;�ȗ��<�M�7l)�v&����4�Ní���\�ƮW�,�%Ʋ:�.��ٗ���ȕ����*z$�3�\,Ÿ�6k���Zz��'Օ�k�}qɇCf�$��sȕ�΄�VlVmƅ�S2��I4�S7=� ���m������7�!'uk\:M�ܷr0l�f{���t��E\�8��5Ɍ}��n)˗�|�O�9�x��I���k��O㝩����[=۵L�zY�/��_r��nil�OpR�} ؽy���<��ǵK��\a~͢�ˈ.wn������=��;��{�������f���y��Tce�r�w��&�7��<\�o�\�Sz���V�9�j01�e!�0ʶ���k26B��-;W\�2�&��6��t�������ѥ{�{U��<����tqbR���욲���'XC�A�^�J��V!� ����낇P�F�C�f��e�K&�U�%��}��ĩ��_U*�� ��t���E*p3�����-�C�����/>(����|N�Ӯ��I�-g�����]:��	g���}����C{��ϵ�pv=3Ԯ���\�#bt�鉂}������5R
��5q�`�4y��>�^�m{%�5�;�!*�QN"5=��E̚��eg]$�e��Wn&��
:�<%���*����]�����GT��{�G�'���$w��mZ}�v<QIWU`�A�Ʌl�q����HW�J��4�����7]�|H1m��HR����n5p&�DK�K~��6���LT!(��6��e�����tR%s�\�	*�l���du�Z�̸vdº"�4LH${G����{��W���G�>%;�h;l�ZI˧g�+�Rm9Z:w�[�9��#놳���7=�%�۹m�Ց���E��]E!�Nf����>]��;���s�ݹ~�j���_Q��]D,�3��_a�u"@���\�俰W�+|���1~É/o/Wn�ۘ�O%kX)��ն�R^�j�O�Lf%��ص�cK�������K�f��U��sL��ż#���kCU�����<e��S2I�/^u���sϥe�<Eɨ��Ѷv)����s�|��W]�Z>,���s��k���Q�9����5��X,�)58��N�w�^�g/3B�Ӯ=k��=��^uaU=Ȃ����#sK�y�u�E��*̶	�2��I�-�������������W�Fj��"�Wv���;<A>�/&�\�������qͪÝ�y!���Q`�-�;o�.��j�R(�#ŗ��g/|��v��O����]^�岤6��Y��u�z�QLe���nD楹ػԌ���~Djƈ�k��[��t���$���@Nnh�v�7��J\�����(v�d�q7&�����*�a�p�ʺʻ=|h�CE�pr����_$�9�]���W`��������%u��kkR�G��Ya��]Z�|%.�V�v9���s��-���˫�j�Y�ؽ7�n2|�]��GX��S�C���9�O����b{;��=�Jy���Ԇ:|E��&`�#p�ie��j�E�.لa�J��	w^����;��ܙ�K;$U��������l��r�E�jScx�xv�(���{�t�m�$4uJϗzO��M�-n�n#S&[I}/9v�}��9t,�|�S��p�m�����w��L�`?,�[�T
tc�S����7ҡ٦�5��n����t�&�1���BQ�+�h�dA)��tX%n<���E��τෝʛfZ��^BBo�P3·X���ێ�[���|z��<�i*g�\"������7�UV���nU�P6B������g�{�k���]h�,I�d.p����W<���/{1�.C<ݔfmĦn>��twl�����v�2���ka��VU)��z���=��a/|�޲m�&L>�[;�yEn2�X]D�I��{WS�Nq�,��Ȭ����}�B��C��rcT3���i�ԷU�W�����Q�%���ND��(�ݗ�&<����d�>DM��<��>7p1kaŀݾg7��,=��}�\�ͨ�Z=�{�:�n+]��7N)�p���=����S�=�k�AM�����d��zȼ��.��e��s��)����*S�9���TGh6��e�շӎ�gL���Ɠ�B�߭*�_�j
-�����g�}�6��o��T�^uՎ�r�"U����ӵ����v`;�S���ۆq�m��v�Mq�ڽ&asֲ��R\��Wg�
���ܙ�0+�j����g8ks\.���HL8S$�Պ]���՜��l̺�(LւNa�S|,$� �h�Y��t)�p�];��(VOU������p��h�-aC��jd�� D�ݬ�/�g8���Xܪ��&`NA�踪k~�j� ���M����5���N��^-�m���ߢ^��&�/�l)�`%9R�Y�X]�c�ؙ����'���GYE�l�Q/��VB
p��S�'+*��[q�Ͻ�%;��S6�ư�q_ܘw����bq�>�����S�[�6m��w�QJ����{g�r�k�'�'z����5f��w_�"U`xLa ��D^:�{F�KȨ�� 5�zq��-��M_JͲ��kinL�l���S�U#փ�G#̓ �����r!��b��)gt�5�1�U��Ψ�«�]r2r�73(N
�T���5����kj�׋}����K.Q���r<ƕ"o��;d�V�?����JN���'t�E=�6��/Tv�:L��
^#׼p�JG����:���D-�����n���e����S8 K��ě��I콴�����uO�
�r!{6�C/��v�<��j�~U��O*�ͭ ���Z��ȝqPu��-˭\�D��v4���`L5�ۙ	j��u�dP��[X���Suқ�׵N�����g����pr�,�"�����wt���%���F�����&�Bn�:r��uY�R��fw��^�1Ӏj�<���Z�굳ϟ>��QH%mf���|��VwUEv8ރ�ޞ������_D{��Z�F���N�i]�����+*M�kp֯�����A.��'�t(��Q��*�ب�Oo^�Q�n�g��E6D�I�����f���:�B"���,zdΔ3Ԇ�x,���)�Gw���µ��G�w`'/�e`ğQw�(|/չ�R�����/������g���.�kW_]f���#�8�=�`퉦��;�'�$%��mL�;�	{�ю� <��V����ʲS7R������%�y7���8ޢN@M(w�(��6����0S�hMBɎ7�	��0x�,�򊎜�4h�/L ��k#��Y-���36�����{&<�}��1î$7q=��\�)��	N�惿�7@�YQ�ae��Kc��j�F���lir�+��M=Q\K�]��e�f��]�6>yZ�vޓ��`v���_�\:��/T����yVbھ/s���߶��:9[����|﹵�g�q�x��es�L�1��)��mU��Š�ӻ-����g�K��;����{\�*���N[^zo?h�6M&��iZkc���*o�����*w#��*#q����r�W'[�(��_d��Y�l�Ko�<�js4,�e�4�����1Ynk4����;���$s����ԑ�����p�����k�%�5w�H@��ƙw��Y��[��;����;AP+>��YO-I�|b@S����Գpؤ���3Rð�t�ή��k�07���j{���a7�',��+l�u@*�ٱ�%E^�еQQ��oG$�����*V�0����43U�8��:�4A��]���?{_����;%���V�G]:������}��<��r�o�����k��#[g��\{�4T�PP#c�%�
�T�i�A-�g7G���⛱rO��5ٮ^2��srE^����ؚ�������@0'��]|�)�.gJƹG8޿��ܗ|5vh��0v^�G�ub9��Dܚ_@���OIk�-L����<ˉq���:�TGt�<��}U9��§Pc~BQ�-��꾴_)�cQ�7��8r�i w3����;P��sܥ�Si���lR����H��\G�����]�mE%]��I�ta6e��ȥh
�*z�����d�B�\�Qf뫕>�
�m�����xں���Zn9䪥���C��h��C]��z;^O����w�omr��ē�Z�S�z�syYI�{��������;��o��ۣu8�M.&�]��s�܁�޺(��JH�;�V�It3v����"�k�����La��+�m�>+`ߢ�~���@?��ߛ��9��p���f���GN��԰(XPp�gKS
qk�G�eYn�u]=�K�z7���oA������l[�ܭ�C���f�^i�ۀ]N긬}l��7u*�Q�T{w�^q�]���&�>����X|A�/�D9~sp�m���zQ-b�;�鑓��6g������~���K3y�NF�S+
#�Խ�*$q]�7 �N�oQ�R_3L���1�>�p����[�x��v{���{gz��n�����py �����T:�[��5;Y���p��&��i��{nC�	�3��֗m��ɯ�((���4�`W
���o��X���B��N��9O}BPf{�鷷�.d��@�&j4s��0�	I�͜�/�-������ե�"�,ü���Qfv�%sr���@_%ӟp-n������oF�/����D�\�<gSݗ�ΰ��*���D��q�9��Ty�0XĮ<f<�]y[�t�c�T�T4&g��}fmR�����t_�{��i�i�-�SΔ�ZEp�I�]ެ���]�r���RA�庍��*H%�7i�������s&!:�_Zx�}87��4VzN����=���͝��;_��l�<�gy��i+�%F�U4��BTL�.�8D%g};��z6/%� �G�o��\@�'յ�cS��`���l��4gD�C�EG�od�)�/L���\�=��L�x��C5��&��jY�F��2	��eH�h%���\e��"�9x�������b������0(=7l�F}Sgnn2�\I�H���y�!� VbI�F��[��u��p�&C�4�ԝ��[�(�}P��{Y��Bx5drD��!�����Tޞ�pOx&�V�Ƈ�͘Ȧ*��nJ[>�0�f�MIY/˵��4�|2,�E��xlu�n���I�r�7��!�zۭc+��I�̣��O{�G�Bŋab,&Lq�6�"u�N��ZIf��BR����Z9���.mt�Oa�X~�F��=:p�-�<z*7 � �V��]t�{j�^ǳ���u�a�HRo{��1�Y�����|.[X]��j���LQ�r�A��t:�&�w�9����1T�X3��4�+�V���R��ʆ��䟱Þ�<�J�y�D��yҺ���.����Y#愤��r�b9�=��޾��6ڡ&/-�{���X�S<tg�c�75qE�ƶ�y�ѣ���q�&w�n�2�u�fú��xj�ѬX�U���f���	�Wy��Z�.R#RPv+,,dެ;*P��t�����S�#Khf�it���& g=]����<F���i֙�o1��ՒmI��\V��s��o;��Y���*K�T&�YX��n��������:6T��K
+���`���L�x�rŻ7:�����8��GV2�O�;�Rlz�U�7I�{y`1^�@&��7Z+iv�9/�_z#l�N���oY]D� ϏT�Zm|/1����"z����;%���[�)
�yQ�/F�Vs�=+�/�K����sv�ה:�b��f�r{��W�wR�ȿ����l]	5G�EDS<+ngf���(hL��v����e��x9��a��E1#�5�����؛hE�{��RE'#��\,6*Q��=Y2���ej�U������e�1l��z{�D����,�]����.?��
l������X��o)cRA��v4ս�m���E����S��ZA�:U�`�z�f��z^6��36���p�\�U�KkU\���|��u��R	;m뛤kr�VF���-*Ė1��� m�Y8�3�#+�ٓVjS,p��n	(�(*�	Yۙ0�,��9D�R�:��.a��\��e�_?�.�Nf�t/|�Z��}�f�D}8�z��C��[� Q���_��φ`Ⴊ5i*	��S

*�20�2".QFj!ZIә!]�DRBAPG5t�i��p������]j���Q��ETQ�0� �AE��.E%B�h�Ȅ�(��H`� ��W( ��p�®�F��H
����g9p�
�L��"�E8�Y��".TQQA�j\�\" �s�QT�0��$!p���9RaΙF�jQdD�U	ʸ��I("!P+�UQAF��0H.�J�JU�\����(��5��vR�*�#�9Z4�hTr�TQXIL�J���R���E���
�PF�p�Q2�UԈN��.Tp�TY��Q�r#�h�\�dU�.YfD�eG""K�J����G2NG5
��-�Ad�˗L�:eY%�"9PL�'LʮB�( �!B�}m÷H���[L�kt���\�8g�׻ӭ��=��E�5�w^���*�ɏ����n����]�ٷq�R����*V!|�~�8�k#�
iC�nd���)	F�P���Ď�:�N#�t=r��G���/*��]�[Z�낋��ٗ�K�_��eL�����Oq5�'�G��}�"w(w:�Gk�]|�m��I9��;1��M�'�[��(}�NlnЗ���ƶ��(G�k�ya�Ǧ=��}^5��,B��	<����Q�{�5����<Q�MD���!����v8�n�ʽ��ŉz�q���i|���}���>l����1��q�Mkmy.o��hڣ�S��v�fS�ϊ�r����н��v]٣��NK�v�`����3�t�D�rcTtae�*���Nz$�X|Gb;]��"�֢�O{�c3���D���[sNȝPoBs[��m�+=ݴw��Eo,�	Q�]o^FI�ʉ�����	dO;Y����b1�h�H텔m#V>H�K��.�;��'��Z�����X�u�z�!(�Î��ͽVhaԦe%j��W���Y�wmn7+��"�:}��],�M7X��`U�a�r��{׎S�qL5�_�ﻶU=M��=��)�>x�c7�w	VW{�����!�~W�y|GZ�'���ˢ��}[u�e�ʉ��Mð���O�=<�N�������=���I/�d6�y�绬�eA�\8��,6���5���gn!RQRp��@Qaײoze�9[C���[�K�	9��DRdKd�����q�q���C�)	Nb��o�
<�ia$���;�;<�?��.$�M,�^s[�og�}}y�1%��藭���<�^S�nzG��W�|������-g�ٖ��²:qF��v_s��3�"NEu eߤq�As���z��S��$C�v`�Y�T���ř9U�Ow����ЗJ�y���5U5�Z3s/{SV����R�u�;\躌����Q�
�n9º�x&�.Lb��&�;qga��a�9m�ԑ��u��x�
vqs�Wlm��v�Җ��R[^&x�$�-f�-:]&�QYT���Z�t�K���ҵ�)�W����t'�z(�_N�麓���+��:��i���`�s��y����vt�='C�#���:^�!�c['Ox����=]\������/��]h�ί���ar�m$jևڥ̅B���ۇݴ�+\���k�*��S���͎�����'01Z0u�7��:Wq�sn7V�V�M:yA�q����s��i+�V��Yټ�+QG7���8��0Gc�+X�)^롒��������h�O��M�75-��~����+>(�߶_�Ї,)��ۚ�T��՛o����>).27嵌����a�a�e�zE�A�qjg���AUD�<��N�ʊ���Lف�����k��5�r!�}5�*I*g�v�5�sk�[䧏�/��E�Ya��݋�<�/W�=�~>q^H��c�թ ��%�2��[�n7���X�	,���>�ȸ�µ���7����@�;�r�v''$\��h��nM��it��Z�I�L��2bQ8�.��h������u�^���nv�0�VA�*�� ���E����Γ⽧Z4�h��Ϻ�h����~6��q��hk+�%��Oq��bx�e��~c�w���1��ʬ���7�{�s�͆�����\=[�K]R���S����5�6��4���f�6�Gd�n�
$�4J4��]r��
�1	sTM����]�	t��M��-�0n$%q��]���&�-��J�i�y�S��_4:�.�fZ�n5�!�J�T�HNA�P�L�0�ӻ���5��	�w�VA/�x�5N�5&�}*�Е.�g:K���Ƈ�y$b��\�ڴ`|{���֍�ĝ�.p����/zh���ټ�Օ�'��h���N3q;��)��]=����m��*�)Rnd��[���w
�Ǧ��'�,���jK�ŵ���:ܼ�9��0�N�+�n�n`Hq���ook���v�ʈ����4T��ҧnN���"��S��Q����jo4\���Y��*_�v��x�5�{��iKlw��J�ү3Wҟ\��q�ƽ��3RSZ(� ���#�p���t��Ӂn�B뎺u��tjv�477�܄�9�C��$UuQ��0�e�����I��]�#��^�B��՛�%��@D��9�sF��8�+_*��5�Q���V�fLUgV��"�c�r>��Y��^����k�ܙ�Ƨ����2�9]C�`]���XZ�褡ǀ�`��k:�Ώ)��/�Wfn^զ݈gқS��C��v��+���<9�\+Wɼ1��etfĂ�ky���
&8�� Y������T@?3q�I��;���vsn��,gS��£�Wz�>vW�2M�����,��D�礵W��ȵ��^N(���8��d���Vk���HR��D�������Ǫ�So�դ)|;���Q�)����{�i��l)�f6ka䚧h�����H�Ц{���ˌ����Qv�2�%╟K�C��X�:.9�e�IZQ/��m�R�ܗη/�_qW�&��ܒzӊ�}Z��ǯ��)5��K6�U�S�,�Z��_�]ݏݎ�v5�6\I����Gtz5��ޒ��<�=Kn9���h�58�4�y�ֹ�t�/n�꭭�e��hFV�μ�M��îP�
x���/�U���$����Ƃ�E<(-��wdv��M�ޭm��> +��H2�.�7�h�e�iz|}"�^����!�`Z��vۧ�WrN��$rb��rl�}� w3z;���Ρ�ȍ�ѥřJ��M�jro!��%B���_MF�'z~�&b�K��Wr����ml�Ϫ'�]��fyqG�ϟ�:��n�*�:�N���-uT%β��k���Yf!U�]�8�u��	����+#���O��ҋ��|]�h�i����W������-9��-�C��K�܁���"�+�H���7��dV����~ծةl�Z���ʪ��csѷ�O3��޺�ǽ'_�{B��v�� w�k^O�c��<�2S�=@U���+"�����5�z{�l��?Oj�ۗf���mc]�v�FM�-�u�4b�r���ޚ��{��]��gU%�rj ��d��K�;�+�]1�x3�_*�.y��E&E�͕��q�q��t�A|��!j�&�<�=���� 5�|̂7�2ridK�x���X�T��N�wϥ������1*�-T�}W֋����o��ǯ~a<*������j���Zw��s9Ai6�k�X�Z���フTF�::�jq.��f���y�ß	�<�ۮ�Y���,�6�b8$f�%D����P������od�����p��{9T�.:!���u[����SA�E1�s\�>.j�o}��W=�Ґ�!��]�	\����Jx�5�wt����w^����MYi�Ȗ�}+"��[�=�=j�ܘȠ�)����j�{IWok��#uN�q��+/����W���:v�_���Ƶ�!�!9���缰���aN�B������oB4c�v���z�E�;��\TK�On��Ϸ������SҜs)�����]��{h��r�����1�����s��V�- ��}O��ՕMŢ]nt����k�d�$���x$�׸=�}�c
k�_W��w1�/�E뜘7g��Ay�u��ۗ���:pyP�P9α��o,g�I��;��(��(%�:�nn8�]�<L㳶ﶎ�Z��Z���왘��hs�����;����g�5��Ί���ܛ2^�-;��c6�����(�w��L܀1{4�sgXo�R��k-d���˰�Y�dt�E6ė�)I�X�5�A	1�Ӏt7�=�``�����:���̅+��V^�7���s,h�ݍ�лk��D2^��t�I>d�J���.fV�:�sxp�<����8�ٵ^����nHi�$�ԋ}�X�jen�u�]���X��Y�s��
���Ib�v�pzV5ʅ>�}��"�j�\�.�QTr�?�'(!dLKW�n�j���.
��.ߐ�Ŗ�<�'�x�k��|�@��fH�X��T�T_�L�U"�����C�sLD�6숬��R�z(�F�.��l1�3��r�{2c՞� ̀��}[q�������gv0�{�<���i:�?�SY���=^��ɞ�X�n`�v��&LlT{��v���J����b��[E��q_���+dc^��}�,���`�����w��빣]��=]g��-#�P,�j	Ϧ��k'cq[��nN|�f˖�w�޹�ֹ�K\ѹǆg}�y_s�[j��3K������]M�!�����c��x�NA�����p.UW[��~�|Pͺ�h{��ax��h~ڹ=۩܎�\H��cv��׈?�����������"�FM@~>��Z��`Za� ��ۧD{G�*��h�&.F-���h��xT2����C��ym�MWr�`��,�%!j�q���S6e��S�^�2C�RXsWc�v�B�t�-S�1�\�elP�U�2�;�&����n�ow������WC����ˎ�쾛�������OD�C�!��x6d�t��<�o_�	��<:�z��2!U��	���!^�q� ٿ����6�ٌ��{�#:9�X�y��&�Iȋ�b/�ܥZ:���=!:^����ׇ ��z�#�7�3~���o��V�G��X��K��E�×~�mԱ��r�p��D����~�x/`��+���꧛5�7u뢢�E�D
��ʦ; �Q�V�>9v�իv�|��La~�t��Y�p焔yguT;#}��Q�{�����E FA dB���q}t�[ّ^��m���Fr}�Ҳ�ע������W�9��㟢#<���d�� �����_�wr݁^�'=�L�E���/��8��Y���u��~����`��U�W�C�Jq�i&={��}�u�����"�ײ3��G5pq?cb'�m�>�{�~�Gg�<*U�AA1��.�=��g��ʚW�M��������)ϲ;�*NBk=1����`z���װ�n��]�`�����rC�FW�ux����{��aח*ە8�vk3���d�r4.����K�vo�� �0��K��2]�J4�K�{[&t`YVݼ5/I�9��m��{ymGib��=�P� ��r���VSSV����vno;N2ckS�:q�*�Է�����^�}5�"���ܣ�/���Ͻ�r�8=~{����r�[�u�ޣ2^ϲ6f���ʑ*`��ˀ�v���o���QaUr��EMX�ם��#����S﹫��������$g��NA��HC�.�����
�{�ל?uk��>�`��{�a �|=�r2
����\ϭV���~��S`^�9N�>���£үj��'����{�n�߮��p؄k��dyЯp�	�al3�������ߠ9�?������}Ȱ�s�}U��'�������υ�`g˩��j������{}#��XZ�pK���D��ު��az���"#�AݺB���;�UZ��`��=7T_��~�y��&�����i��u����t���.�V����������?22�(��_�dw2�ğfL;v�;�$�㨣�yfMc��C�޿O��1O��e���۩���.��n���I����xZ���
	�dxw�㽙�����v�{!�����Eѕ`%
��* s'�F�����T�2�o�\��"�]|v��fm�ί��/��Í`*�#FPN���S$=9u����5e���I����!��_^>-]X����b��;S+��]��
�(�Z��&5��,��2��N�ZrR�wx�W��Q����㝆�n��iw$�
�|;��$㩝n����)�8yp˚;sw��'V��j宥1J{֥��Fgo;�9�K`����nrE��w�D6D�-o�&�]��>��o���W��K,3�Z1�g����q�*�O�7S�3�_`���	��t��u��pΛ�&Ռwօ
�0 �'#��8���3��&T`��u��M<ԝ^�������!NxZ�L�^N�\:�Vl�w���"vu�5���V5�T�OI�j��/jZ���a��ta���H嵇gP�'�����x���[c[�`��m���F@M���{OeoU����l ���(W�}k��?\�p��f{�}w�_�}s���z�f�w�l{j���珌��������6:�|�����3;g��n��3.P���3���;�ǩq�/��na�͖�0y;Fs�F�y H)�6/�`4ne��t7,�f*��Yj���n�pI��e�n*f�Dt�j�Y��x`L�Ò�����G2k��+e�Z�F��(F�6�wƤיp�o[��֤�e5;6�d��l\=ܵ�0����M�no�ɽ3@�k�6�N6ڤ���k�
R�v�؊�i��تÓzY;�L��|�V��%�[$q�gA�����f� 	��7'=��[���|�E��\�u�r���Dm�7�F1���D��8��ۤ��)�ԕӹٻnڻ:�*	�깝��9R�5	8�p�-�'��w�WfU��A�oa�Y9B�t2驮ę��]�,�X#����t�z�����0P�mE�2b�dΥR�ܢ��j�z�Ǜ��p�E��YH�m���B=!���vJN=9Js#4�E���4G7��=�A�4��)��2�&�����
jg7���31�2���!E^��*,RbSq�&����2����C;�jm�|�0�p��*Y-��S|��O�	��d��T�R��[���ޑP��r�R��	��1l�Rg'vv@W8܇n��Td�4~���O��CSl�C^u�s��_v�r�(f1 Ȉ�7V�)�O�4���]0-��������f�]��_atk��`�j��ׅ,7�*=�ټ��A.²i�Kծ�B@8�\EgYJ�Z��Bd�nU�Ҭ��5�\���i3L��sT�>��!k6�
Wr�.�c�t�\<��j>x��y��w��ˮS�`�Q������\7.��܀��,�|��Uw���\�]�JcW8EZ�P�o޹�ٔ�:q�:�Y��r*��%�x�y���c3����&�8�	��%.(���P�j��7����.�w�Ύ�*�ݬ�:�9��Ф��-:aT���0�)8���q2e�2�8��	,�U�Rt(���̮QDP���.dQEE+���ȃ�9A�9QIUQTU(".r ���DY$�QEDFaTF�AVE%5hd�UEB��¹Us�UTr��.I,�
*PND�W(ՙ��
*�2H#��TW
��Eʪ���*�B��
��G$��Z`��B��*
�r���*(��K��*�KY�U�\֐Es���iEʨ�EG��DUG"(��$̒�"�W+$�(��r�y[��EQ���������,�p(eE ��+�Uӡ˜�B̨񰊼a$�Ī(���AQfUjQ�16k@�*�
M�dUE\'V`am�E�`E]R#��FNrQ�*��UQS��Bd�)�Y�4�C�ʈ�����U���uutbJ��e�jZ+Cёv���y�f�kV�vYM!�b��cz��GWYu����&. ��b^X��ЪL�JLP]��8j�g�O�Բ�S�ܺ�ȿz���B�O�#c�R���,��X�ϢFHAt���r@��I2}��]�ʐfc��
����r���Z����Ld'��G?T�9�d�}ըk�'�`uU�u��g=�FX=�+��H��	�<F$+���Rd?+S��9��Z7�W�ٺ{���H�O p�w늸b��7q4@���60�4<y��z�T��{޹�F��4^j���
��O�q���%�_�fm�ȫUN��D����To���^z��-F�$6�da�T�9��H\{ƽa�^����̟l�ٛ�l���'C���n��&�����j�W�}�<���1�7ƙ�^�{������~�̟l�̜��mP�Q$��$/G��{>\u�����}[>˧ç��r��O�}�7!��!|Ϣ�c>�T^���+"Ew��r��=��)V��!H{A��A�����]{ç!c��N|�Ndzq;�ll'��~����ɘܜ�}Y�8����{o�u��;� 	�?m�B�����Go�㙞�+��LyQ[~��(�<�靐>Q��[�����Gw� I$Gsź��Ӈ�km�<� ����u z��P�j����ނ�6�Xj=�0����n�c��6�q�K�Mv_�XD@,��p��ȼR݋wړ���b��Ov^ù���t$��0�:9�ۛ�v?R���T�y$���f��u*X�!��Ƚ����䊋�oϧ�ŝ�l�^TW����,�����Cc�p�b�%�?i����S�p�
��P��x�f�����z���W��,�X߁�W:큟E�}���b���Y�FP���@Y��~c;��=JNqJs�n{�Uz���gg�iW'W-|G�ӛ��_��c��<tV���3���aU~�|�h�:�s1-N����Y�LdE�y5�W��gO���7�,tu�� �sS��U�J�R��j����9C�Й�9��B^���Tۦn��޾��}M�:Q��aͿg��y�E�R���	����}�*�_{f�?Y��u>R>�7d�T�9��o��,e�9y�ֵ�y蜯D�+s/)���O������1:� �:?�
���]/�;Ծ�顸��cX����Dw��8����@�����ۑ��Ι�VxUê���R���`�GW����^#��z�o=��3�W�;�Trf�c�����Wῲ�y���$%�+�S��^����fvD�5�/]�u��ԲǗ�'>�i�{pV`�P�ܹx+`�k[�d�{�:���*�X�U�Z��Պ�eĊ�sk��a�٥�ʹ�>�ܘ���v�n�a�0,
=��澹֓�bS@}�w�&0�ukJc���u�QѢ�+��.s��l�ߒ�FC^��G��,F|�����j1�ͯz�yJ�]��^�%������@*"�w^�����W��6��5���[�dT.��g�S��Z����zMףM�9�����]I� ��>15�!g�����dyw�g��kFN��v߷����{g�r�ho�>���y5��u�ʩ͎�\��ჺ��^ߐ���=>b/ގ��M߁�`1�f��A�Y��w~>��o�\WdGnt��m!�Ѡ<��,�՜.�(�+�G��=�w�.���$�����Q�`g�+��pJW�^�mWH^�䙃~�;5��%\|�Ut���9�}t�t�z�ʌ�2���H�Nׇ�l{/�ڸ����n����_��w!�Y�8�<�݂=�{n���W�nE�]��w,3>���z�"s�q�s��|o<'up�W[z׻[�
'�A�e�gba#�H\� dC�i�]Q�W�n�Sv���T���[��q�wYmϹE6;{�2�?c���ed���$�+�n�gy?��ֿQ��u�x�G���SV��H����N�����}� �`�zC.����yL	|j��3[s$60^�6�A����%/�0��'��쾛�#���K�f��oIJf�tFNfћ�:�̊j9$�7$V��m��>�$c�풍�+��Yh��!��Y>Ȭ�+��p�^��w�e���V'�~��l�� ��Kn������~�K�k���(����Jo�"���Hhu��~��s}���*��Haq�� ��;��T�y�R1��^�bj��#����(��թ[�?cb'�m�ǫ���d�W��'�1���:��q�]ݞ�>���z��P�I�"W�\��k��1^�dw�T�Mg����ǂ��O9��>�5[�oq����7�K�ؓN��S ��U�GD]3~���M���ϰ��O�zw{r�e}�gmUwZ�~Sf���>����>�L�C�ɞ��ʑj���R���f���e/v�7~�ڙ�W��Σ�>��Gt��{���C�\ϯ>~�L���^�NmԋU��H�d`��XbĔ�U�l�&A�K×_��a�.����1g�3�U�����S���פ![9h�Ey����>�����g}>�>Ƚ�O+�@�x���=�#����x>�̊9����骟X�_��a�~s�ӻ��/<t��AC�:��/��G��gE��vr���c�ꗳ�G��/���/2D��Ԑ���z�l�I�b��7�;�E���72w	K�Z:�G�)w��&������c;�t��e�H=�Κ�dP�<��ʷ���m<�oU��uYH����Y��[�����Z�w��ve�]1���q�s=�Ω�F9��ȯT��b5�W>vD<s^A�h����GS�:�/
�,�_��QC{O�⯺�i�����Z�F��3iۮY*��F��ݎ�㹖�;�SYNwox��)y�w�>�9���G�=�����b�IFz۩쌦 "�/��c��w�=����]���QW��ݏ|����>̇�z�ü'�۾�lף���w��2�"F �r <K�.M���v����I���}��{.گO=˯�z�h�~���|�F�d3����:�;g%V��>����)=�2�}*��a�r��x(�z��W��zu>�4����rd�1Z/{{{|��p7�vD,���2��X��١8j��wCe3�ReE{��x�F��{�����Y�u��⬐3}�����b��-�M"���62SCǘ�.�D����->'{V��T���%�G�hlD��Xޭ���⛪�RϤT�3���3~��a76����<�֣���Ňk�����������jG����(�w�6��
�L7*����H>����`���N���7B��Xz��w�;��sOnI�$�C��'�fwja�/Td�]�mY��5a�7�&��I
&�<ո��t����n�3�M���2GD��N�J�7�{���M�C�0�f�Ƀ�sWQ�2�o�z�+�m8�]�(n�\��=�R��WJ���>�~�7�E��a*��n<��a�^����2}.砏mP��x�/�@K��G�B��ץdI���K�O_��m}���\6�vDz!�E��}�4n=FRchm+�7�W-N��(${��Z3� ��ڏ,���y�׸t�,v@<iϜi����w㱎=��v>�͎��w�_?-��^��ނ�&�u�����h�����5�!�׈0-�H�G�إ/�ՠx���y�V7�>��xX���x=�N}]������|Nf�U�,���o�di�-�9��&oüX�=ffw�^ʔ�C}��l/;R�ٛ�Mm���� ��Yoӝ�Yyb�|�e7��z3�q�X��R��G����_���xx�.�~ŐO������D�ֺ�w�/s	n�����sU�8r��Q���:����{z�##}s��l?W�Ǳ�x���s	kY�д��=�=��)�BA�Jf�G�s�r�_���n��n�k�zL�G���Mlg�=���8�<O������X�<��Z +�Nf�%� 6�|�\W�/���/ߕ~�)h�?���ZYcc��[�6��^a�z�+o���}�Qx�y^�WS��7x�.�9��9�9P�-n�WO�c�3��6��yfao�c����|�Π�7fq�(t9{V�1��;;*�[��`�D��nV,��fa-���ƛ��ÿ�>�]~aq����#Av�}9A�3��
�5� a�^��O�Ц6s�?,P<����O�+>�yj�o�~�$�}���4��	�n��NӘb\�4*xF��*�\��4܏A�]�hTq�������=���}#��3�z�­� Н��c+��ٙ&��I�#�P���jo>Y~@��B��Dw��)����?W���o��Ļٚ�ݪ�W�Eo���}���U>����@��U��z���}��z��2���{�2�dBo�,fo��|D!��sH���y�kSs�{��6�װP��1��h���:z�{���nN5���{��:�:���o:�̵6j��s��&��{��8��98}�R��v�����}�Xdx��E�f0O�q(��7�랟i��:�w��O����l��ד�-۩܎�_�6W�@�m,J����F|ݞ���41�p,zb�N�����\�p����+Lv�M�V��4�p��R��yn��x]�����ڮ��4u8����>����%B�"���O�����+ڢ�<&'d���q�<A�z	���Q����2̲���@��«�ӕ�+#W.2ll9�u�!��u8|��p��8-�u��q���j|�s�Z��jІM�(o��F�<T�T��z�fZ��iT}�L�q�7 C["����|z�;�B��M��+�":t���D#�K��é̮�~�~Nׇ�lG���r�&�ï�+��m@�B~�zDiʮ<R���(�&�c�;�����=~�>�h��-ewi>�U�]E3;��alG����WƧZP��4��ÚQ�]S1�q��`:9�/�ւ�)^�E���]��;�^���\�/������r�0��C���p�Fc����򥜯��c�c��E!�o�"�"��p�^���deg��ۯ7���&?� ~��՜�Ф5,�*�F�j�<{�s1βG�𦇶���ߍǽ^������'Gg�bw��+ݞ� ���7�z{�w�&��y�cbe�bG�E?=�QC9�R�)�>�m���=�v'U�d����[�?����Uk~(?$x���K�k ��Bꍫ,)r�������\ۄ'�k{�?ۅ_nV['Fp�O�6&ݻ�A�z&���L߬m����n|	�L��nV@v�j=��O:�>�s.r��lO��'��2g��2�\*`�,��ۋ����D׽+��}�W'�y'ʯ�}&`US��}��Q�NN8���]J�kʍu0�=����&,X�j�v��&\B�X��WY��'�^G�5L�@����L}�Ik�Js�T�7l��M$
�T1��8:v���&VbjB5���4HBX8����F8�������Ϛ�g��uvC�\ϯ>~�L�헷�}�R;�^\��E@���{�;���K����{��<3��$y��d��f�b��}j�<v�{ݹ8���rO��v��V� r䨣�#�:�9��t���OdB�d7�?�ز=���F��^��+�&r�&�K�Y���G���?�2?!�V��?�V��x~t5h���3�(��͝nf�|�=:�׷��B�S�UZF�yl��ގ�W=�Y�1�V�,�
��^A�h�-�ϔu9��\X�7#|oNa�Y���>��<r7�e����=���h��ۮ���@�z,Q�xsٖ��Z�tJh���\�`�锽$�L{x{�'#]/z�G��>^�S���f�۩쌦 "�/
H戫�^��s�+Bõ��U���R���e�C�=~����w�=�[�~���ed�z*g�bz����Qڊ�(� �R���W>9w�W���xW�W5�y�4�����ީ`�����=�������4=ƽ�o����@�^��r%R���l9؆rφ߽jk>�{��}�h~C���#��?�Z^��c֓�b�o8DL�I����R(�'��Y7Z{���N������7K�d�����T���;�k��U)�I�o5rJu*��)5�n&!ג�U@1[��@�g]��K]a�sF����r�s��3�FΜ�5x�tu�E!��}$iy�ݱ"'(0�fR��%�BvR��b��}jLϑ}>���>�:�u��V߲}��x����{�G�~��b���p�K�ld���P���}�63�)����Q�i;Rg>���Ώz���l��[2}�Ȧ��D��Đ&��� ���ٯb���G�d7cݔ�7��C���.Ck=c=�Z�툟_�d�e��ۻt*�S ʄ�#޼�j��#�t�]ϴxz�n�_M����䩑�_�#��̱�C�^�?z�O�"^�K���N;V㦮wN�|�K|P�Tx:�
OD��yK�Nv3��߸�# �܇��1g�^�N,�AR�Wu��#����SK�g`�c�+F�Q�螾��u�9�����>ә��ݟF�56U	#�o5�[�WK�︫�׶�Gauּ9��i�;�UO΂�4���DӮ����̏o��D�������X��L�n�R����׃؏;�$l�7��L��l+�����=�c�J��өL�����Z�q��1���S�){�7�q����)e�CNS��C�߱�;�hv{�F�J��p?4�BC�l.R�f�\�HJc�^(U�ǀ:[ch����ĭ	rS=�D�X�@�٪ vp4�:>w�Q��m?��q�|��6��o5�"L#x��e�׺�;��n$n�'Oo@�i_B@_h���>�r@بn	ji�Sq r�O:�:£K� sP��v���8�V��d8'��W��[t��FK�փED��fLP[�X�st�k�/�;�}�����g�w���-mq����Qn�R�U��˽�d!�<;=Z���ѽ��' ��^��V��*m�[���4�_,Y�q�ݞzXƛ.�gn樿+�nm��]
�h�ܫP~���o����[���Y��t�eL�]��7��eۄ����AV�
+h����/ ��$g��V��7q 8�5n���^�S��v3�-�t��(�7C��s!��m�i�'ڂ30�̞
��+j�Q��gN>��xu�d�����)�o�9����R�h���2I-'K�(��{j��Rl1�I'f Sg�c�[n�����_jŭK�],����W�B\{����Ɋ��Ƶ�v��oM����E�5��wy��R�n�NĠ*�%����F��������|y<���;9�nWcxoڀ1&���:y}�f�ܯ��$�v��T��C_:��v)h���k�&���l��·6�1ǐ��sT�%��S��jq$x��5oZp�Cq��7z�!�V����򠋒��,�.�>N�폯�-L������6'|BjJ؍E������׸�|��w ����v<[Dm)
����9gkb�=!@��]J�\z�K�w&��O�:�o)H�u+u#���q�85�uX����iqg`��%(wi�,e�Ζ�s��Kq�s�Vm��>P��*�f?��ZXJT�P������>ˑpvөb����=�0�r�����Mvw.�oi�apm��^W:��Y�&x+Q�:U��0:�3�d����M/+Z�h�f�~ro����ӳO{*k�c�!GF���u�n5��?N�tK����<�Q=�.,����<�z����u�@+�2�R�\f���ƃ�5tzB�T���u�qf�V���z�ϝ@��Y�LR�*�݃ul��腫`B�J�S熶懎X�{%*-�ˎ�5VJ��Ѻ���v�����[F�j-���=�j=n>o�����޹��^}�d*ϸ��f:^H�B�Vj�țx@�Fj\Xg<7�k8��d»��P9`��j��&,�";|A�J��>�Ob�wdR"�}p���Z��lgk
�yϜid$.B��7g <�G�_�ot�^?�&�����o��90;[���7�n�;+Iw��#k�!b���S���&�wu��XB9T
;�RWN�*&�۩o�"vW|��r
�F��n�7|��<�~<�͜��w��{�8�Kv�Q�!�t �Q\�(�E�#���"�ԎȫDT)��\�"�W#P��G�S��)D9ZW"�ª'��&QDQQEPUU��QU�Z��$�
���lɦ�.TFt�#�$���ZΙTY��J�DȨ�HK�EAjB�"��#��9�B"���L.QG&QRI�Yi��.r�+�ɪ��G+�T�"��T"��UD\*4C�dQQd�
�5e2q�.EEUU
*�"�#�*���I,��9ȍ�eDTr"��iL�!�
�"�"(�L�"���\����AEp�W+���r��UDUEDh���Q�"��EG.UQEAT+��*MD�QJ�#�\�9yJU�}�������s5�Nf�F���n/���4�,�7�6��w�5��-�('
)��P�9}J���j���4��Ԥ�b]���
W#س,d�D�7�k��'�~������~cز	�n)�ٞ��󾭸�y��igG��F: ;�2�j�� �߮�۩�Z�W)��H��σ�?W��F�o�*Û�рv�7mE(я����E1����
s5<���嬿��t�C�y7��=&n��у�W{o��^<���+�;�W(�y�xȿf'(!p��
C��	z�rSn����:%xr����ѾY��N���E�}�0��x�Z��!۸y9A��&'��k�ݐ<Xѝ�]��w���ڻk9Fx_����.
�+���>o�~�$��N��ۚ�uAҙ�n�f$�l���AJ|T����>��쌏
H{����sB��~����i��FC���s�VxP����'z�f��y �x]&$�;Mڛ�Ym'����.Bk=c!���������?14W�����g(�j��L�:��U7�Q�B���t|.v�.a+dc^�>Ͻ�b;o_��j�:��`�G�[�[~=�bK��Ƒ��q;P�D״E�5�ӽ��E�q�$Q@vi!ulkǘ�H����h��m.�w�_g\���s��X��	��l�m��P�d����6�wW^�"��3�b��3��:��e^,7�z���\ݍ���y�;=Se(�3Mq������f�V�c�rDsgw�<�qW��$�sQ�S+�.����VE��خ�J�F���w^����^ޜ�>�|�P�^�;��?�t��_�{ֈ�@X�w�0c��Nϭ��g����N��ߐg�>\x����r�*�S��+��̿D�h���]���R\5�ҢǠ]{��׼2b�N�;���W|�p��c�.+��:n�hm�;����P�{ǋ��2�}U�'�O��� �`�q7��#��ׇ���W0_��9陊l������%XU4G��ڥ9�C�dUzv�j����X�u>U:�\zF'k����l�tWv�5�����t���ގÐN����;u���!�)C�9w���r�ߠ�^K9��܍���}�r��~����0�O{������`V�;t�D``"��)[�9v�ծ�Mt���ʸ��|d!��G�s�&�{�ӽ�xv�w�e��s�
����r�� +$Ua)�g��P;I���l�z>Yh��x�Exe��"���p��:;޹�F�P�.��Ϥ`�M��0�:�����3�^����=fA��������Ȭ�_�!��x":�x�{�����b*2�VulZnz�G�����;c��]f�=(��r["قܰ���N��T7d�V����*CǼo���E���n]��g��o<�QOW��*aʝ�\H�7�}������%Y��p�tt����=Ǩb|r��Yw#�
}7V����B�mT����)ؐ�E?=��29�R�)���8ث��ۉ���̧'��]״��O v+�
� j��7�lMP^Us���W���';��U�Gx�U!���O�UV�''Ë��>�qꌉT�(�?���h苊f�c#r�5~�<qe7���xz�"Z�I���ϡ�~�>�L�l������ʑj��$T�3��ҽ}�����Gj���ٯ4<���oc�G�Ϛ�g��uv�\ϯ>~�L�헷���u"�x�0��u�rgs�e�:����c%��w�2;)�����da�܇���g�3�4�v�}�v��3��䍋/`�vo
\�U-!	���'������Yl�G��Yt+�!?Qaf���q��9��ڊF*�Q�~���hϐ��섿�5h����.?�w*s�������Y�=��@���Z�����9e�U�q�ޑ�o��|��Cۚ�kEp��g�a�����z�ۑ[������}��aB�}������wJ{���gNUp�0<�T=(�7W�����W^_G]����W=���2�q�vo�X��Χ���̥���Fk>J[]yo��c��u��K���tRߺ탰�L�3�g+���x��X��Q�;ҩ-Ҳi��<��3�_�IgOq�+��j5��KKp	ڣ�����13�ovf���N������c�����K��ğfL>�z��λ��O�ǳ�N��f�!��̦ !��2y��US��~-Oi>|=����ʵ`���9��zG��7�S��c���*�����<�&	*b��߆E�k�����=N@
��5Q�9v�z^]W�{�s^-��>��doz���4��o��vl��^�H�Վ��X}��䌑�jϕ�
s5*���*�>�Z�ȯ{��)��^��j�D�[�ڸ���uV߹S��p7�LB��L�X�-����\�t��9���Rp;/��w-�����Q/=;�������$���W�)H?��n�����Pz�;��{����Y���!pVw�ԙ�O��z���l�1���>�\S�ED��ç9Q��,Uu\k�ܣ����}K��3�e6�Y��>bද���R=���̟C���ۡQ���^:uk.���)X>�U���ٺ&�o7-�ll%L�/ݑ���e��Լ�~�̟fF�je�c���X����Nw�� ��C�U�i�ȟV�˥ç#�����F��������������5Fi"������W�<��/v�l�a���n�+�g(�>F��y�t��z��ක�m�����յ���ݵdRN��'v�y���'R�䏘Tӷ�r��{/r�PkA&R��h�!������ 6��$�.+3F�s ��g6�����C+���Fh��v#�+FD���CY=}/.�ç!c��N}S���W�!R��o�w~���+gcc��+���+ɣՓ���np?!�5C*~���-����i2o�������7l���)���,��;�a��^c��Ih���n�r0;� T=��3>��mO��'r����`��lO[��M{*]��C���k~^v�oж�ޚ�}�<����~R�.>͊Z�U�@�Uv��S��AǙcW�|đ�j{��2����{r��b�&s5j׈����)E�r�w�h)�4 7U�w5F^���a�sN�9��^����O�ц8�0�"�Oi�pQ/;f�w�V��;=BA��9��A�|r�_���n�ǎ�oO��fh�]vPg��q�wX�\�9C�=�w�X9�#�E�C3��< W��HK�S���X��F+�d�puW޲w�R=�^Ʌ�0��tvz��������&'��s*�77�Uc�ߑ����ʨ���.
��({��o���2@���Og޻sL П�L�?�CQm��83h�4,kMr�7�8gL�1��n�Ƅ������ɗ8��s3�wj��5r��"��o��7���d�]�pG3���8�����5���4����-�Pj_H�)	���+�^HܽSH��r�!l��SW�B����E"�e�z�5IZ�d4���(sB�����{���_H�~�t��L�|���o����^�;�>I�hMS���Ym'���w��8��X�~� <:�Q����w�swq��ŏ�	ʊ����$ ��*^�Y;��\�\,�l���b|jmǤ]�Z͢�z�ǒSf����/����'�.�H��b`��jȚ��u��c�{.`�tf\�k�f��\��������3���.rz��X�^���/oNNA�]H��xq;P��;�,��>�ca���}�A��G��L�����w~A�T�Y����=���1��|Nd��GE?ƛ�V�^g�N薪�o�d��pߑ�ᇱg�]�������y���yq]�v�M�,��׽yG��`'�����ӑò��,z�^^����CӉ�����ݯ��`��tӝ����YW*�U8��W�l�KD�N���?�\%���t]�?E��2��="��^���ӑ3�5٩�*�����v[`�{A:�P��;u�"00<�9ۑD9�9w��K;�ogiy��3V)��\Ȫo��%뽅����g�Ȁ�C��JCw���d����]�n�-�wP
�VzL�2��^d�L��5�mK�Wy�U����s]���0j�|��vO���#�͖�e���squc��gp��v�0lHZ��aX���r}�D��=~������e���XD\#�Hf 2!�l
V�=8�W��4��C�w�腻qG{ra��t�z+��޹�r�ψ؊�2�r�0Il�Ei��Ș�j�����z2'�u����s"�2/�9�M�l/T��߻�2���<ꜾRH�@*G�ؽyiCmQ[���̵WALԷ~�d6f�J��+#��Ho��x"9����\kg�o�<�VxOxՑH	(�A/��$7FF�O��t1E�9�R����)Ñ������ֽW�/oݣ���;=w�Sp�U�.��4'h/*�V�xs��xӨ�M����ͺ��G{���T�wZ�2ٰǇ�Xg�p��U���nj�{>�: 3^���KT��R�qY豻&�C<�|[�]JW��T�s�yf\���y���2}�K�ٛ��ʑq
���R�޿W���:�U�Q�6�e��J�Խ���<7�����9#!�vz}�WaC�\ϯ��${b^�NA��Htu�]F]ߠor��X=��ul��}�";+�y���yp���g�3�U����Qk���>1�M�	ؖ�"����i��<�t��KRT^uu�m`������E��W=���Y��'=�\
���~Z^��&n��q,�ϲ;��@]������F㠆o���u:#�ԙ�������k�^s�s{`���7����#��װ���q+����0���V���ۙl�G�;l�{���Dx<u�_��{k���^�p�=��"�~��q~b�d#����/���Z=mc:,���ܜ��b�==���c�{��^x���FϾ�����Yal?^I:oH��Up���{q5�֊����Y�W��o�񇃗�Q�I�3q��/
������{/�~yjI���iۮ���@�z=���>�W�v`��َ3�q�XϽ��|�$�2a�{�ޮ~���o��N�Y��v�y��ܬ����q�|�]� `�B�n�v0�9�3�o2����T�>�\{ƽj��x�_O���>�H\j�������R���S1�P��mק��]xd_�y4[�pG�>�*�1t�CƯ;�!D�H~��߅c$d�-@��Nf^�Sa�7]�޵5h�_lkuX����_iw3'���K�:��>��s��{ vG�؇
�W�����١9�y�z��S���l�^�QiWz�|��N�{��|=�='���#}��=~���(1p��wD��<��A<�={����y|W>�S��-�Z�X�4�Sm������n#�̭z�o�^��%�T:��F�&��5n��4������tZW���b,�t{p��m2�a���^���ê�-����٫;��N��P�ɀ��b��M�H�ڛ\��5�c�A�l#��s[Re?;r�{ր�ϫe���ٓ��E[��R���0��S����&�F�>2��|=Bk��n�B���a9�#�bද����H�ϯ�2}��fD{�j�]�T�o��Y'7���V����!��s����=R&F����w�C�^�r��<ߦt���4Vﶱޙ=�nd�ڠ�x*�ӓ�D��^D].9�v3���6��/7!�=��*sc=��w�kw����o��1Jǣ�Nh��v��h�|1;P�O_K˯p�Ŏ��5~�=GrMi��Fz��ݙ��_��a�T�R~W�G:�nm{n�gi�?P�+ȸ�0&~�D�%!����|=�Ԏ؆s�3q��zv߰�W|�k����p0v�����L�T���z={��58��EX�+�[U�hQ=nfW5�O){�6=��[��)eq�tT��幵���{�q�ճ�B�eL���1^PYOi��9*�f�\��x�T��yp�/ڨ�-xL��Y:�(�7�f����ϱP �R�@^�r��Q�q�Ӭ���%��zE�UF<kE�Wd:�9�v_�M��(�R=QD���Fl^�M�y��n��}b(��d!��"1��y97RK����9�)"��3&�T��bټb�]�7��B���W#������O=`�=�9�2C���n۾�������hbpoq�F�x�u%��^�G��M��w�+RpR���@�3_D� ��+�v銣l�"��Ud]{��+"��ߵ,����������G���y9AC�p)��D��U#{�U�Y�'y�z���_W�ˊY~���Ȧ��;��_�]}s��o�H�����\!1>Q�4����c�e���{�>�}z�h{S��Y�-S���|�fH����]���ȝ��;WB���׍4{�:��&e:���5^vda��9��4.}	�=ZG�'�["��l�C����b��?��O�[y��}k<*��@40]~c�5O֦�[@��B��w��9�k=`wq�>�yՓ���a�įw+ۀ`�� =� ���A�� MO���yw�����/b�EqpK�����.�[���g2�c��
��OyK���װP�q;P�M{D\S]�9��������\��l�^ύq�כ�o�|��\���s�|��>��~�L�^͛���׀W;P�Q���c�����:�J�C�x3����f�a;�!�������������Ɔo�~��4������ff[����ZA�e:T�3���u'h�g>ݫ�]Cb�AZ��JPlLU���W%u�Im���zb0��s�G*7w:0RxJpk��z.�E�������t�n�1Jrvg��f��I��Wj���lr�ыŊ�)c��>����8~�BI;I1�M�-
�{8m����b���kT�zdD#Ӧ��"�.]%Z5�)��Z8�U��T��H�GRl�u�������[���d��coR�B]2�$�Kd�l���85�ݹ�\��;{O�
s&6<����\���Sv�,�E��Goe�k�n�tz,|��ApW���HtaӇ	j������� �%Y >m�_�!�۔��l�eObO�/5�U�Ge���S{)����35%�:�Z�r��rZ���G��QǴ6�\�7T�W�/rON�B/��s�+�$]3���K�7<�jۏ1��f�r_0��Rx[<f8��+�"��V�Jef���_;8��{�;m�N��rg\<=���ڷ�1���>}<.��ӒЖ�|{���ڧ������m��p7�X�ހ�WH�*PWfv�0R����K��F�2�f���m��vV���)f��q����U������b��#[]BkP���r���׎���:We���\�DK�?wMtvN����G��ځ���`ˀn��;�/����S�m�ט���	��|$aC:Q$f���a�xt�I���9G"�;�����UW��9��f��K��]�Wd�GB�^��d�*>�n�Xh��GNJ�Ҵ�\�{\"�`�[�9{@;ef���FiL׺񮙪+�y�]ԙN+�a����&���"��u�8��6�g%�)��$K@�yٿ�ý�����H���sbBuK��NsZr�dF��~g�[<:o9�ܷx��cp��o�7���m����	��c?��p���Ӳ���l)wz���VQKM�%pBk���*����U�B�QY-�z�g�6.��R#m.�]�$ܫx�@���J��J���\�^��o,o�7�.克[v�q���ݶ|�h�ur��sD}��>g\Us[t�	��\߮EZ9����\ ��|�K49��-�s��Z�`o%r��6r�_J���t�b��kl����JWPr��~�zk�4�˫���u"�����v�Q��y���G�!^{����֎kW��'HW3+���]���:z.$�٤B��p�D�֘0��B/��أ���CݗcRppm,�c@��*�W0ۭYBِD�	�����ǋiZ[;[!\;�Vಚ�Pɐi��`�y�d^Rב�m���r�knp�'�//Q��t�l45��4��ޚ�Ĳ+O-w2��3�O�4��c=�r/G��P1��Hg�Չ,�~�8t�zG5H�rz;�=D���|9^�5_Qˬ	r��}�` D ("��*���_�H��Pr�TRpJ.G+$�"��r�QȎE��ˑs�*��D]7�����r���"��Q�n9e�IG��֪ED˕Ur��Er"��Ƞ��S.4�ʢ9�QE\�2r�A2��9r����쫔E�UG9EAAETG$���UG9\�T\#3����9Q�� ���2�;+��.9�E�8E̹.U�dT\�� ��r�(�\"*���p�PU\����e�J��
9EUʠ�(*("�99@��"�9UU\�*�ENA�NA\��E\��A�G"�.�Tx����{>�tc�:P�y����5	��pad��Aj���;؟���^w�Ot���F`��9�au��N�Ԇo2 ����QG�����Vא�@С~�g��W��J!��y����xz��{;���V� ���e�G�H�������d`�^�u8����v�<����%~U��/9[�OH����U�ڮ�^�ò���V�z�NDw>U��2��	�Y2�ߒ�x�\�d��()��~�:�d�;�"�N�pȌ,�S���C���~��75�r�=�p��;�((�����q����_�ǲ��Ȳ#�ۤ3 �C��#4e�����Ό�,��5�ݸ�d<{�O�{+��W�;b;�2�?c��V�K�h£�MQ�3Cks��B���D��pM׼��ȯ�x�VSy��|�w�e��T']Ɉ�~��r�(�9Ek7�S����T̯U�3פo�Sa�W<����Y�bC`:�@ԣz�U,s�sR���>��<����uR�PW�TݙS�s��3�jԫܾٙ�0k�w;=�;P��`�׋Ç�����dz�¦�uA���D�T�\�,v����/�x��D�|�*��u��]&	�{ܼ�u�]5�YoVtm����%��Z��/'�z 9��1���&FF��p��2!3�#c9]�_�Vp�/�kLv�j��+�qs�� ��1
��_t��q�˒mcݚ��#șyy�%
�����V{k鐴�����}�T�y_�ˁ�,=Z�{덉�n�S ��B�M�6y�"=�c0����'vjW�5�cݔ���j�� ��O�#�Y�-���3���6f�~̩*`Y'�v`O˥o�<]�;��=�\��oݔ��G�C^���������g׏��=���n)�<qO�m��~�׍�X��>���N�#�VʯWh���PU22 �nCO�d&}s>�R��������xUϳ��RL
�Q�ۓ�{�� Ӑ���r�z�^}{~�WL���q��{G�\�j�Uݜg�YU�u~�#�Gi��Y�G#��c��>��շ�_��G��gE��:�y��(w�xٜש؊�L���S�����G{,���$�XDg��B���{�9�n��p_O�{��{��Dѩ�^��L�ڽ�¥���C�_���$���f��������]�;qx0��Q���]�އ��)\Z���=s-�I�d����`��]/z�G��>^�S��YfL?U����̮>�Y������ P(_�)\{U��|r����4G��6;�>����*��j�/�{7�K�H�*�%!͋{��'B�]C_^�k�G�iwOg u 7>O�-(���k)�X�4�vg����s���ڛy���O�3`8�������z�(Vt�SWE�Q3P�1q}�ʾ� ����P;+�iޢ���#���#�3�y%d���ꬾ��# w�� ��r"|��n�/.��_�y5���V�K�l:c|���՝�^���԰s|�߅c$d�Lϗ
s5�xVM�;�Y���j��M��%s�<�Nz�N9�߽��4����d�S��-@�JǬME�	��&��h�6�� ��[X�b���|�Y>�*G����{NzOC����A�������s��|`݊���=���}Y��줇�1p_5�=)�Z�z�����f}��E>��U���}�c5�k*�$I"x	�ԍ�°��?%��3��.j�a}�zԏG��3�Ma������{f��ݑ��R����pnRc *ٺf�o7-x	S# �vG�#�y�7�h�ۉ�|y�wW� ���72^Ϸ2p�mP�U*���ǆK輈+?#�^�{����!��8����ו=��������_�dG��������Z0� �v������^��ǽ�L���\�>���7�y�3gҝ{�>�^��y^M����^ۭ�!y���|����e��V�����:��M#)�L
�f'�+�Ř�C<mZN�7��8�_�b�w&��V�]�6nƮ4(_��h[,B����˕�fu_"6R����s�ufɇ�sf#�E@k�F��m�gC�p˧z��ʮ�]i����J�f��zK�K�\#}��^/��;~G��v�g�a���s���w�H�;Fw�U9���]���?A�͠���G`�wȽ��.��[��f�s^ڝ�������k~^v�{��=u��N���<�ֹ�u�Q�|}[A�`)ު��nA�fX6O�_^��G_��N���t��>ы.Gg<^Ψ�#�� ��ۊo�5�:s=@qJ} {�˿]FA�sN��~��g�ƽ�\�E�%���c=�=�����.=�#�E���c� �
s1>A���Y~� ����ߥ�ܨ1�I����#�:�o>����;��z���z僐��<v VxCȜ�����Ng�Ҽ����a@;�9h���US�R*����d}~�����J�_�\}s���Ԏ�Ë�
����ff��,�����P���������r
9�dVG��T���C�� do�bz�p�PQ^N���z���پS^���UǄ̷R�����2�5C�h\O����#��؋7�2�$=����B����/gL�Ы<*�� �υ�c T�jo>Ym'�
~�*9�S�#���jJ��a�rQ�ʣ#cX�O��P�s����F�U�C����)��ެ�x�U���Qݢ1y{���5Փ���yc�M�]͕M���R�c.RH������J��|9�!��noym�I]7�>~�U�oN���X��c�վ��fmպ���X���{7��\��E�x�	H1�u\��9�UFx�tГ�yfX��߰PϽ��I�˸�=b�R��;P�M{DWt�϶1\W��Y��բ���垿{�q�%���&�e�C�\����4W�f�>�k�,��kP���{<ua�q��1ȋ��Y^#˾+=&s�ٹ�N��>�K}�4C���-��u�D��s�M����f�O�W����#g����my����Ş���ߏ����U���}5���;QH�W����n������z(z�^E��Ax�z��=�#�m��tp����/"����`��4�~���G�]a��h��ÛIxc	p���t]�?E߯��
�=���5R����Fy����_��Y�B/N�p�,�nE�޽��E�Q}`Ryy�;����+�U�Q����k�_��������Z�D.ʤ``��T�|:���շٳ��[��}��Q����]��l-ۊy�ǹ0�{:v;�^���L�Q���meWӘE�K��Q�_��KI3:fŔ����ez�Aқч����\]�*gE�ł����jޛ�E���|c�]@w��Y�?L-]m��{a�p��E�Y{K�e
eF���dD�\EgT���4�.��B3kH ��5v�B!�Ǉ+��J�p��UaX���G��p`q���Uߎ[a�9�^���"�)��^���d8�4=pbE�)z*��f��0���r����f|����j%��)�٫�A}o�"��_� -�@�M�g��Ǽs�������}���8��HaD���$7FF���|�6��ϱ�7ۏϰ��9��}D���6�Q�2��;=w�Sn�5SB�bD�*����0��ȧ����1����c|�9}�u<~Mg�Ώy`�`5>�؛�n�`��^�_���u����zV�v�z���Ϸ)3W���}��*}9�{�2�w�=�������ٛ~̩�f��LR�s�C=�s����~�S�0v�_�M�������kݞ�������gב��<$�E�|��D���j/YQ��>���H�W�W:�0Bθkj@�#�c�
��0j�<i��5��ʼ�kwv�G/��+�&���Es{�>C�U�k���ӕ�=]/"��<�����O��rn�s7�칭�o��dF��׃�,ȣ�~��q���xuv}U��q���.��K/y[�٨+}o�ɋX�I�J��.ow�{��z�v���כ��hU�a�,^򱞥������
z�m����ɵ\Zo�P���顬�����ʮp�bL�pb㔁<���F�vd���é��)Hx�தL�ӶX�̾TZ�C���ݠ{��f���w�ǧ]���G{,�-~��Maw�u�!v|*��j�z&kc���v�QCI׺6}n��iTϔm9��/
����zF��xyjI��ޝ��Qhȧ�o�9}�f}�%Z���tHu�8�,g�=s-�I�d���	��\�����ڟOwI:�OK����:��l�ʩ>� .(y��+��*�cS�c9��{z�ü'��Y�?(����;���	W�2g�;�eD�aW� @s9>W�Su�Or��/޼��txG�G�4sqy��y�籏r�a���o�C2-�~���P&|�Q^|"�����x���C�43�Z�}�)*�w��M�k"+��=;	����}S�����T�3�Q3)O�K�������QƇE�#V�S�$&��xQ�ϭI��{�ϰߧ���H�d���_�Pb�	�i�6�!qtR>�}�JՌ9My���ړ8��9؁�Z���??z�gj�sDv_�ۋƛx�v(��o�Z�~�R��hH�XՔ�7�d?�*8�k=c�jG��5F�xի�Dg��J���?Վ�M�h�p���EZ�:�ݛ������o˦b���*Ɣ>v�ۍi�]�w�Ly�=�E�P�'���n��=�HF�*�R8��ٟu�Qr����ڲ7�۽��,���&��n�9���T����Ra���ک���M�B�`�O����o��rׁ���21�vG��ƍ�\���޼����n��MM����(��d�b%�d���Uci���l���ç;�M��}:C/�'��<h�n�=d{�9������Nǽ��G���"�
џ�h��ke���K#����!G��������~�j}�s6}:���lC>�^��W5˯f��^ۭ�vq"��X�l�'��Fg�k���d����㙛���=;��|+��׃�;�$o�h����߼`Tw)�7�Ł�=ϴ��{i��"=�~W�������O[���{*W�){�=u�r�>�e�'�Z��X/��e~{~��5�;2��x�~�F��wc����|ƃ^�i���	���w�CL��'5-��A�˄���d��Szkht�: ��O�,�W���w4��ު�5���Y���,����
�##}s��l?W�Ǳ�x�
�-�����O�r|p8���]�7�Dj������דy�=&t�=n{{�,���x�@����9A> (��`���������.��ͺ������(��J�e;�)�T�}�=.�e��o[,⑾�<xу)XA�7�����n��[����b�Gj���
<���䣚��OE����e�n�C��3�g\�+�e�5���HP��QKᕕ�\�����U��-J*�q����=�ɟH�mT窚�l3�����N}M�:u{��.��}JF��p�;�x�xU{��PQT����LO���4<�@^T1pP�~Y��-S�_�/���o(y�����ݹ�������UAR��n��I�ň�"��.
и8���"�a5�'�PZ��ު��`���g��Ι��g�_��h`�ld@4$?R��Ym'���~}%�ps�-�G�22xof�w�h���i8�{����o��˽��un��K� UB�*��t|.g����VNN��G��6��D5���̱��
�W�O��gA�`��N�3�*Z��c=Y�W�q��1�~9��i��ܖ��\���s��s�~�L�^͛��=,B3�{N��~����uY5�!��+�yqY�3��sҝW�Q��������q�p�7 _=�[ޥ֌��۩����:�l�'���W�B��ö��}��}U��j������j�oGX�=U�yq]�}=մ7 פp�x6���E���^���O�o�|f7kު�7�V���j����r��O�`��*,CU}�^�����t�;�0a�� �dPɋ�\�7#��S�[�;��̶d��ďF�Π%��qm*嚣�ƴvyml�EY�AƢr�ʕ���|k�z؈��Tzcݱ߫�+�)���\�~w���ڮ���;*�1��.��΁����%_�V������Q�@4f}��􂝯H�e����A:�P��;u�#�9�nd�9�k�͎=��
|����b��{��^K�������O?W��e��߅a�U!uKld	T�27���IK�@�Q�\
V��S�En�SǏra�!�gN������g>~�> �M�G�q_/A������zPȇ~W>9nV.y�^���G�^��ze\�]'����Z�[�D�g��F�b{!ݹy0���WE3R��FA�z��)�\S��B����žP{�{��kXDw�S��F��'�=V�\C���}^�5Mّ�S�s�1\���=^&-��D{Q�J߫���xa����c��dz�¦�Pj�]CphMF,�Yc�����-���W>8�{½>��ʓ���K����լ�>�ؗN��S�_}ٷ\��9�c�P媉�B�
�:޵c>ܦ�ZUsYR�!���I[�K�������6��1�m��m�o�1�m���cm�66������6��1�m����1���cm��`����m�o�1�m�1�m���cm��6��cl��`���m�o�1�m����cm�ݍ�cm�cl���d�Mgr+ƴe�n�A@��4 ��~��(
B*

 �`  @Q*P��QD� PE*)QPI!J ��
 �(�(��*B�� �e)!P�*HH� �	BJ)@�lQ��(Q*	HTP�UU[iJ�
�
(QJ(
Q=hJ�*!*T�!U(�UQP�G�$R�R*����U@HR��E*�٪	($R AB��PP*�UUT���64+�QIHx   mW��Wl�A�Ѧ�M,��h
����T�k�N�� MPc@Pj�U#UUT䦠Cm4��FʕURP�BH��"*��  ��%UUYJ
�M�D��4Ԯ�( ��r���4h��4sQ��=(��/x�: (�En�� �p��E QEp��B�TT����*�A�  =�DWVʨ(��1*�ZZ�B�A[zP(�50"�f *�0ґ@�������JEII%���  9@ �EUMd��UP��R6�[RJP,���5&u�v :���Q]#�l*���ֱM�(Ҥ��*P:R��#�  r�5��k�M�WH�:�m�9Ŷ� t�,�@�Ͳڭ*��m��ke4e��j�U�9��CF�-C C�ʧ]]	)F�+FDQ(�"IUC�  �e�WV�Z���%��۔�;c�hf5n���VWF�ΔUʶ�vWlv
֨�i��m�m��n*���֗sh*ۮ�#���Q�*�JUC�  ʞ��twX�V�JP	����Ѻ�L-�Tֶww���tYMWN��X0�lb�@5]:��j��4i�7N�.��dT�DH�%
��(�� �P m�׶�7qԠڦ�[k��6�h[V���ҕMg�Xն4��Ttu�.h�X�uݣ`�U�Z��ҦU��3]:h�R�x  1�Ц���J�^�m����
��w@P�S�t�T4������m�� &�R�.E
f�C+�(Ӹ�U*�J���P�!�  -O4�@R��m��׸��:i��kB�����F�R��2��+��e��Yn�l4j��cJ[k!���F�u;�*��� �~BfU)J� i��E<0R��F��20���@�y����20L�&S�A)R�`�M0�� U22i�`�$�SA�I�	��6�I�S;A�`�D�:D�V �Rܣ%��d�׺�����}��~��!$ I7�� H@�~�����! ����$�	&H$�g��$ IBB��l�!I����t�$��_��������6��W�ӧZ������TR�T�5p4Y;>�T��.���;�1�r��Jn���I#ƙ+��v�3�lݔ�AkՊ�N��4��Ӭ/Z���.` ��V��է	\k^���|wy,�	v�Hg"�Z���#1(��L]O���W-^]3G(���2�����Ut��[�Z��Խ�1%�Zm�ԝ�Yr=ۙWH2-���6��6�k]b@�y6�o���T�v� ��F�n)�������Gh�T\
f��*�ͪ[z7[5�y[PR�Kk�Wcŵ��se�m���`�-o[߬���nر��z��R�I,m�)k� v�{O��ދcX��Y�Q�m�hƪ9��PJ�U��N�f��H�*��H�3�1k�8�Q~3ek n�.�R
�Ғ&LO+p���]�z�wV%�MǹGlքʭD��@��oE�]5c#����N��(�Nx�
cr�n�Կ��"8�gf����ǖ#I���E&5�*���Ϯ�YÆ险�q�*�=�Wy�-ǣTF�[ ��t�T�t��
���2�CAޒ�2�=�� ���ۤ��SE���Q;�9Ff&���cF���ݢ{5��V�k
d��M�:��T�j�YT/1!��1�u}���hkh�M���r����D�ӎ�k$�[����r�'�2�eQ�nݧ{>���	��x�*�/�bF�X<�q�KR̸M�az^��ۡ�ᎃY{Mس.���Tz(A,�ֳFX��X��ą<��� �.%an�f�Vfm�cnk ueH�ۼw&P�m݆�� �?[PA��)�խ�1J̀Cۺһ�Tt.}@�Iuw�k�M�C\�yw��X)jO#b�Aw[�
�u����e����W�E%4]�A���$�I�p������!��n���P�9��գ�/Z�9i�DM������RKՊ�1a����QCk"�ҧ��
:���{Gw�[<:����0�;2J�8[�̴�2�׳�4+�X�
D�N^%ߤ��F::m����Xu��(��f��j��/v}��9n�>ŊD��q�w�o^8�+;
&��^K���wY ���u�ffF6�M�P��ǣ�X�]�eS���vL�"�DĶ��D%�գσ
�CT����V�N��ww��yV��f��[/uz��9T�PdT��X� d��`�^4��)�U����M!��uX+p]$�w�q��m�.��,� i�C5���'AX�̊Y�.7giS,�X���[J����T{l7l$��{|5�.���9�l�˵�6��W��,b���I#�cw1���d:����9op��r��74Xӻ���rA�Ɠv��zm�yiXڅS�Q��M� ��Ɨ@QJ�6I�j��{�X�L�MhF�*�4vRZI��H��2�L4�4�D�u���*��t�>�ֵ��/m���4�`�*[,IT�I��HʵR���]�d�+�$yF1��[�t���l�wmn�5:!\0Z�2��;2ԧ�� � k��x��۠�_Bh�J��nlQ]X:&�ڣA��I�j�c���CY2�\0Si�i ���W[.ZWe��r]��d�hͶ�BW��,�U�����ݭ6�-6A���w�/5e��m�skn@��ņ���]���'c���ϳ�lӚ��/qiq^Vۙt|��ֵEd��j/�������n�r��ܤ���X��PXen+�m0Ɇ��^'���g;Z�(��y�ʺ�(68����Ex+4^��ʣ%+e+�>���n�&&Uּ�4����|d]�8��Yܗ
m��M%�V�TW��^<E��L�.ܳ*tn�����	�h�j%z!\S�w���fnB-�lj^"�"�j����WBC�E�[�6�(fG���Z��-��j٬yB��˚s�wBwN�[2�B,�y��+؎\hд�鈥z�a]��y��6�;r�ȈwN�ݳ�Ŵ��N��e��'�dB���:���MA�#ջ�$�/$xH�,��c]�C�@���pbf��eY���g˰�lU�i���|�L�A�j����V����̛���P�-�0R+/5��V��t�
ˤ�Y���6���]�.^I@1K*ebВʋ�~n�3T7���-�o��n��f�X5d�Œ`{�Rф��c	�k�gh!C�-�rA]�>l�.�i�y2ܙ4�[{E�t�)0�,�»y*�=H&�<�e m�n�mm��͊��H�m�F�����w����2c�9��&V��\��!����5���K�a���A �����t��{����u��
+s
�Z�����9�2�uZ��ܽ�J�de�
8.�!,�b�^��k$�5vM��ЧG�GBCF��^��i�A$7E�a�Y�S�/w^b�Kİ�X�*��TD�����V�s)nq�ޚ/i0�x�H�QkL�����Z��*�Ч�4#t�Ze<���Z�;���̸$���8���JTN�5��Il�[�ܺe�Ѳբ��Y���jK�;�n�$��X��v[X���S
�%E����,N65ݙT�J�ZT�Ӽv�2����wZ �U�*=��t:�ϯ�Ѹ��x[�B��W;l�Ghfr��#�D`���5�eJ��xF�ٲj����Lw�-`�Vhf�R�t�g:��n����e����˨�sQۏB���JӔ-N]�+%�ksSCz�GB�rZ��a��j�.��ݭo��%�(YתRf��,3.-9v\̶�K��ͤ�na�	05�� ��-�v����(\�B�n�h�[����T1��ѫ`I��ٷ�)R+�u�'m)
%``��V�R�6�P�M���QwK.�Tr�e'g2�\��X��Pَ�P�H�V�iH�zۺN�������E�J�Uva�'�C���ӤU����5����6�����XM6�a�rń��F��sa�VڵjJn��^/�cp�Ktd��^
ɯt�Zݷ1�����LR�J�u]^ ��N٥��Йqn7h8�!��ؗ�%ż%���A�A�glXAm2-���G,�v��%��@,���YE��]^Z�%6	�hee]�T�+�N&�2�^f���{��a'�x�V;�h)L5wn��;E諚.U�8n�ʼ�7�12 �\�fMZ�Zd'5�H5*9�J��f��k5��Փ4���[#S۬!���F=��Mڰ^����u6�t�N�4�5Zo5�Y��;��lt�<�S&'��V���:B�6֚/Gk�S�w|����E;��[kr�V:��p�b�Uz����+��9�5A��@�Gr�'�&�V�(k����VՏ��ݨ��M�����i��I�g��X�{և$�����񹛸[�n�ҺL����	
sEX	�z��m�/w0�׮�\[��y��t�Uq]���o.�!������ڶ��6����l^�`�\
]϶�����{�8��i�ڮg����d��QuK:�&f55V�PH���j�бR�F��^YkD>(g����*�ve�5v3��X��%�2���`����¢QV	�HL6)=��L�ē���fSF��r�"r���xԭ���EL�	v��D���B�Όm��u(��eo®�����D'���n�X��G(��!`ֳ��x*��,k�T h�a;L+����b�0����m��M��6N��Z�� �fi.��ʅb�&�%����E�X���\�r<f��*�x�P�[��e&-'�h��韈���] lG���,{�	� ��0�"�[IЖ�3�\Ln6��,Tj�ӻZ�;B��I�Yy(nn�q¶[1-Ǜ�|��s�@�A��54^� L6nմ��b�&�=��n5[*�l��l�X�Q�̩��V����ܑ�%Yb���7o#]��j"�eh�4�Q�hSJ��^��J�I� ��*F�S�ё��]^v��+5�//��ͶS-E� �B޼YN�`�3=����c4�G&���ӗd��5��9EN�0��!�����4�n��	ֺ�-���Gt�;M�U�-\��k�E��[���&��i�X�5Չz��r4��)w0�oN�핍�T�����G76�@s��E*Th�XY�mv��m�Y��Q���Ұn�*`gf?��V�]���L�׍�̗[4��e�.�]4K�6�fN�X�}m���j�-f���Q=�5�	���٪��[5�>Cwoy�e�ɇ3i�٨���N��t(�H�[ԱWY�7�Ve,�w���V�
��Y��eY�Q�b� M�y)^aڛHi�@MM���4�,��{X�5���6��3fcTYN�GX��U�T�"ʽ��/m��H��ę�v�M��O`7m��#&�v�V�]ݸ��+-�Kɣ1Va�h�b�~.��ʭv t����y��h�x�]n�֕zVm�iJ2���^�Ǵ)�Ƣ�uҵƸU����T�0*ˣWA�$�,�D�YN�nefv9k8
Z=XN�fՊ�������N�"u���%)��vA��y�������[g����m�4S��4J u�W��xr6�rJ������aĶ�HV�C�.�$�C�P�M�ͥ�qM��m���R�d-7Kn-^�ՠ3+-�ON��װ�5˭�!�+PV�]!L��9���<��Ggf���۫�H�_*T�w>!�a��B�jT��`���O��f���݃`�Y�mʻ���݋/]+ܦ�ֹ�[�D��*��WvwMj.�����5�{���!VSݢ�|����a: ![�#j������֠O��L�N��ۭ���r-�B�$h�8�X9XY��7f�n�:a�`��P{�h2bug%��O�W`��t�j����q+f�U� ��ff�޶)� i�˵��{k*螲��j�^� �ΨȚ�m2�G��GSDM:�^)��ə0�yyR�;'4��wyd��iXN��z�Li+�h1�jhт۩d^re�U���vPu�L����1�*�3(���q )4��HF���Љ*�<t���T�haz�P$�"�(F ]�kr�p�yxU�$�୒��*���K���6֗Q���.�<�+en0c��:�V��A��u+��4��.�Z��c����^!�� Y�^ނ�n�S[&�HbM�ѻ��Q۫H��?������Y?-�K�],�r��vΉ�`�N�GS{��������;����jQ��ԩ^#�鴯A��A���EI�(�kM[�ɆL
�O��*Yݺ:��\�'����lѦAz2��N��U�1u��i�F0uմ�cܫmd�m1�{35%q�+`�!���Uvm�Pf=M�j��+^Ϟ[lP*�^��Osy!u$��u-釵��~��拷��cw��ŞƝb�����w&AX�	A�`�1lŹ�$ܳ��M�v�u���X�ٍ�v��Xu�I��`�+�Yj��H����;]c+N����]g�]`�-��ر�Ldӆ�ɘ�m�)�vǁn���hMYab�M�J
��R�Jp���If�^�N��%���4�2���Iv��z�틱Xh8�I�1�5��������ô�7�l���3�����W�xK�Z�,��qMZ0=���>W��D#k/;:��C�CJ{�o^"� Y�H���M`&Q�t5�֐һ,�+�up��]�K�6�gsR[2��$l��3k#��Ҳ�����% 3
��Z�%�c�хʹ����*2T�[	��-�t�]�*�ڌ%�U�*[	J�ʦxs�#��9c2J�ΚVԌ��AP̎�ٸ �/T6U��S�e<ˌS�Oa�[�	e�;����LIJ�D����8[����m��1���
���j�MbYi��z�]�� �[��G]��ộj��P��v����m��vn�����ۼB��7��j�T�W֕��l(
�CF偌����e��ca��D՜�0��wfC�)�	�SR��0�oIʻԚ�j��O.�A)С�9.��b��k����-l]�o-Ea������`̽yWIղa��`x���"oU��wx��"˫l[�,L�#�u�3Bܮ��M[�����ͥE��8+0�â&S�����|��ˬ�KiaBV��[�%�O"�u�L�4D)b�3T�b��%���X�Fޓ)ҋV
���6nʔ3)�us��*0�@��wD�Z4E��SE���cy��ʉ��S�O1�X@up���*�`ϖf\�+Tnj������-V꽭|���]c)�ַL�F1 tm�&�عX+`yZ�Yˢ�.o#�4Rw�gZ���7^��ۛ�-;G55��Y�S$��Īm[�E �s�a<m�����![c�iX�9�:tp:��#��R��,nku2�T,��4Z�7VT�̻�l7��Vr��{iZ���[C%��]MU�m�j���[ӧ	�t�z���s�6]���r�wv���"@B����Z����F���-xZVmZd��R*���Bղͥxٖ����ZY��#]Y]��	�]�0�׺�+*����.G3��v/)<���a�(徧wt*�s)�k��mM oŔfQM���-�kNC�`t�����J[GtT���Ѭ�� f���wq)W�(�b��̎c�l��h�)�DZ��)7�З�o�L�3C�sS�.��9f�:b{�U�3*�r�܆[�ġ�+6�)�¬�׮�JѪ����O��h�vAuf����^�[l�g���n5VIܺ2�˶h��\J�+#e	<��'e�+1_�!�%���JH�ͻT�ʟ)r�w�1wh�P��.���XVU��+^�v�6�9��0��Թ��J��fM��u�19��R�G$��8d�n#��fx�����@���`S�O��ȎX�ѩ�Q�_֥�ǋ\]�4��r�M(j;�p �@�2�`i)�����b&�$���盉�Z��[���د����T5&;ݡ�|�"7y:���&�qe�����ε��űn�94�K����]�
3�:�&:��*�6U�]d�6����vhZ�7qH��\�r��ϭ��wgN�{��WFVԽ�Y�fE*գL�-j�l�Y�Y���������[i��#X�:Y�2n4m�d���6����]�Ю(��Yiu�u��=�-�4l-ͫ�b��<U�o��q�.eE�E^����pH��%�t*>���6��ok%�#�g�Mv.pq��!��D6�^'6��C�}����M/)Uҏ)��ƗxV�)J��6k���'���Ȗ���f	�
7*^9zA���uKL�{5m:��5�.�����6i=v
x;f�պ�&�,�n�����koOdV�QIm�W2l՚�ښ(*qd3��2�d�e�h�+�V��CY����({���jާ�P�y�;�&6�Q]G�6{p���^�K��5�,�t��w�������k=���z�9���X�H�╳q��߷n��7�b��Gp���F?�׊U�Տ��+R�:-��)n�Ux����Q��ö�kt[�k���l�;����֕뷲 ���>��x^S��"�Ms��D��(��[��!�N��Q \��M�c@�eg^��-ܧ�8���F��h���ctY��n�(�Y�'�o8�&�6C93..Q-d-Ұ�&�I.�7��2�K������뒏�qA�~�B���U,fH#��])���|eG�M���� �ü���,&�4��`�̥B���!�0X����nYA6���7\Yw��ȳ+;�t��S�^���&ayI�<���)�e��H�ˬW�hõ+��\oj��:�k�R�	m"��U�����m<ͷP�/mc r7nݥ/�3/���QǳA�o#�]])V����YR��/�"Âb�{j�י)vLu�9]��R��΁h�|2�"�ʸHx�����M��c���R5�k�ko�zS��Z�!����pۨ3���e΂�!Ĝ|5��Z��c�.��;R]��[���-v�Q����溳�ة�ͽ���sa2�U��`42�')��ӷ���W!�4N���L�&�9]c��B�pq���f��uٚ+*v����ż�R��0)�PE�o[||$��;E�Ι[�C�������C���}�b����L��9F���gl���)af=I��1:���e����Ζ^Cr
��448\�e큚�,�-�Ы[�A������Y\�]aر5uh.9� 9N����m_Y[@\DOhW�^�v�bK9
�
^�Ge��PZ���p�ܗ����.L.�Ơx<;�K�s.�X1:�Mm=��d���Q�(��7�r�7v��mmw^�Ǜ�Sy�����6�5`�FI1IjX%��U.h]�Z��sA/L��U��S���3f�Լ�Ԫ��n�Ru�����r�i��֏p2�b��a��)��b�˖6��FMꥲ������c�*	������� n��;b�-�NsT�7�^��J8���x֞�,�BƞҢXV\Q�nP����]c�,DYu�`�]�l�˲v:��d�\�e�WN�6��ʻ6���X@&�#�ro7�^����V�Yu�Y\�ix�ܨf��9�jv�#��` "��tʍ]�{�񥜟aV. \]43Kc�u��VcNR��:ͳ���j���*���`L����j�/���F�&uq�C)$~*��u�r���;U�j�"���W�8�eJ����XZ��i�Ou�z��TƘ���G���{8����0��v��.hF����{*X1��{��:s.ӗmz^�����ܨ������,K`T�OF���B^v���w7:۷�2�Dy�����ށ��4PV�lI�=%˭� �K��ǅ���a t�-��� Tv�U*��{EYF��R�Z(��K�!�$*B���8�3�=����_+�.M�j���:��k6�YE��P�@5�+�Ho�����ag%φb�R�r� ��a\O�.�{��j�w=[̦:�F�|7�ז�.:��o�ȺF.к�V��X�5��Q��י���mrL�9F�ZVMI-�H���븗 �H�W[K��]v�J����W`c[�>�M��6�zW�|nwo3٦���4t�D�v���Жq�o^e���R& ����b�`t�i]1V�L
�	y���6��m�8U���T\�L��(��Ҳ��v�wi��wz���]�����Z�}���b�5�U�_f��Wx���%1�/皆)��nɮ���Cjk��� )צtF�����M�7f�����V�ǩ
���ݑ��o��3�p��f��h�	�\�j��9���u�)К6��htԴWf�G�Հq@K���d��m��c�5�=qєo74��*�V������M雫�$NGz���\����hٷ|k����%���ǷW��Za��4X(8��b�+Q�ϔ����^�C=�4L�"��x#}��]�*�-@Ȳ�ɵ�n�Վvr�� ��P�g-��F�ɋ�������c�qې�,��o���>I��H��w%f֜ä\y���$�)��}7S��]������SCP�;!��Փ+��3� �vWuni��D�w��a]�D�����Z�N=�ުw�0gS����)!�gI�Mi�v1���I*ˬ1E�z��\�u�"�!Sln����0a�����ٹ�.�J�{gCu��Z���\��hIV�|�Վp7�����|��p���We�nV%4���vQU��xk��bI�׼UFF�#�L蜒��*6�,��rb	��M@R�fh�\ΐ�]@�3�;;ulOM'����7�6�l��@fծpb�
��1�ھdڕl�89F���m�y�v@�Uf���<���zۻwL� ��
\5jy���5lf�F��L˷�ѵ��=�R��Jx����[t���U�h��Z4����w�;��5x��n�����f�{f�7�a�rm3�]��i��(s���oEv��;�nIu���q1\$@��^V8���d����o��5]K^���+�.U�wv�����L��m����+��`U}�m�d�U�b[ڳ�M+�C�r��(����_56�@:�����&�9���/�f�G2�+�����z��Ov^rv�.A����7�P����6��ju.�vw�CR�"R�U� �kޫU2��J�'�7��v�n;��I�#A�J�;��L��ˋI�9�ƿ8��Y���ҁ^N��9�A�[yո�]u��P��{w٦�}X ��d1]7��l�O^nWu�R���9�M�j�x9i-���fZ��ul��8�<��*��y��^�X/[b��*u�C��wx�tt�b�ǯ��ʳ��`��l�Ȅ7�n�	j��:{����+GX��&��3�1[���9�l���7H�V����ۺ&�,p�h���YJem�ҕh�(b}��^���+7Mu�U&����Β��F�˾)m*�Z���	�X�:��:Q/F6�V�v,��rX�R�T�F�#;��}�H졽�NbX��cU�N�#w"�!����t�7��.6�k����]�v�um�u��f�O�ΐ��TnŰ���hƃw&jBs���P��RD-�K��iK���`P�5�^�T�>X/2ea6��Ŗo�.�/��FEk�Nt���[Ʉ��	�]���H����l�wO
�}���:{3����Лo&RQ�9Gx��W&�<�R�P�Ud'�O-΋Bq(4����;/.䇝0;�f�C�H��T[3o������h��E�pBor���q��}kV��ò���Tsh�TKM:�r�5[�;Xڻ¹u�
f*�`Tst�v"���I�o�Ę�د ǃ3N��֦�캎q���<*��(stn����uȚo�ӹP_g�w�9Yb�3�g�[��"WY�tԻ[nؔ�w�Z]�R��n�q�� �.��/n�L�=h�>D5ċ��緪���n�a�Fd��������{ɶ��Wr�̒�տ�u"��)�F��a���d�d�B>������W1��E���
��t�9#��0�O�Uz�J�ɴ�wN�\��b7@̡���96V�gSSm�A����ܚ^�u�:	�{{�h�6tVw(�WUv�WtF���n�%׆�	�gW�j���*;$���o1�ٜ�5�<��]�A�"���Xe՞��|\7�&.w�:#-�����A�;�������?�(ӚI��u����D�;�vʭ�`{��J�і��Ҭo��\��Z[��6���+���d��fT��H��mrb��@�ʹ���X1���s�� }�[�뉥���3����4��W�\Zs��*�r���Qc�H#5E��9h�[��r�%�W�)s��8��iv�-�÷��X�9����N�AW^�"��5'շ���,@&Q��Y�9�ڮ�S�p�c��T�O�������;�hL��_>׏������[۹��6��Au-����є>9F'��rZ�W($o����>ʻ��2��������SyZn�s���V+�%�nع'��㙪��YG��ɬh�������{�f�Xzۢqvb���]a���v�}��G�s��z�]�f�=���<��r��"Qf�_13;2������dR�)����d�3� N�{c��;����q�@塰k�`��l��O �FԚ����,�ڙO��U�)_;r���L���ۓ��h�Ҷcn�U(h����G��u�ū�/gw�5wu��e��ueV�r"(_+�M�o���fk�%�����tt!�v�ա��J����F�Z�q:p�O�aYD'av��4�늃�\�\��}K;dΏ,Vb��mM��*p\6���ۖR��9aQ%��ɂ�R���z�5���N��	� n�L�˰/�G'1}�.�c f���e�Υ�ʡ�xo�9W1��N%�Ư]�Wy��;E��=��[}ii)��:��Kk����ta�沺�E�u׀5�7��a�i��ނ)����Yڞ�A�4���w�d34;�Ï8�7wC3|r�t��h��J�V��t�`����,�3-fT�Vz$.�N�����4��S���h]�}��<����ﳚ&)����Ne����k$��$v3WYn�
Vh*}|����%)j�v�|cn�h���XtG-��]��Y�$��Enc�s�]�<�Z�tH��3u�H�Y�����֙/�:̶I$�st�դu+�[4_ǩN�����R����M�z����'����������͌k��%d���OY����ۏkj�Z�q�:k2uo4��7v�r��r�Lx���Gm���]�M�X丼'��l���[�f0 �3��Q�B�5�3�YK����i*����4����n�"ao�M%T�x_�N�5�@vJ�VYR76�����l:�,�Ճ �[|x�sdgf�bT�8�u;}�cVhI��N��^��	l�(�%mB���kz�+pL*.�j���3FC�iŸ��W��`v��e��뫆���\�fc�
o>ά�^���M5Xtەi-����Sh��cjR�z�y�ϭ�:��]�X2��������T��z�j�0f��U�{k�;V��Z��)�aO.��Xȉ�Ϭ@�V��wò+���x9Ӛ�A���mT����7�F?c���k{U�ϓ�͆�jc���o-մv�N�N˝�i�[9���8Ƣ��t�\^C�&^���yMm|L��,�=��
o�0�:�9Y�J�ݥ�242;�WI�/b��7�,��k3-:#Ӳ�4n:[�z��O�LTӸn�k���M�[z*el�O_�X��u�|�C���
+��p;�94_0N��.���X�P�,�Ĳ,erTÑ�f�5�,�� �)Z�$NWR�`����Mm�u�3�q��2ޑ����$��������8ťwcvK�r�hcz2qf���5�4��\�q>2�Vs�M�m�gs��Ú7�PK�
�TR���g%��Y�W7r�z�^=��|�[�\s�����4"�[X�:_X���b4�B]а�oL|5i��J��6o39� ���H��4I��W�sr)��q��l�α�<u�홌�Ò^�:��,�C�A�$[v��g[}�V��DK�j�^ꅑp��� E2ސ��������#�I$�9�%�b�&II�
�[�Y���]
P��׍];L�	È��8uk��3��$�K�>p�#|��Z�`U��Y�8\�4<㐼:އݳ.�efn��z4��{���'��q�[X�s����=��eh�J<M0�����RJ:u0K�y(��cF�!պ�R�������:	<���R"�n*Z�4o�vu�:�ټ
p�������S�Z��1k�<����r5q�z��Y9��ѭ%P���������ڏ���s"���[`��Us�^>�C�U���o��R����8��m\��T)���I�,���;YgZ1˴��b�}ۉ`M#t���\�<��E�R�Cg_e�rY�K�F��[�a���Eྫྷ�X��]N�BR����=��_�@ �� H@���~<��{�������#�\�a���S�w{K/B'k�Fn�@[F�ӽM�32s�)�B��
4�Qg%�u�k7n /��۽���i���C�S�o&�}�(�/v}��v�n���/>J=��E��v�G$��M냸�ċ6��ǀ�V���}'a�E"�)�|�jB
�Q�r�@d�T�T�)ts��qK�h��*y/�*aw��؄؟^T���.ۗo�;̴ -K��vË)٣�wm�7/��S-�m93�vCj`XӃem�'�巚^����/��[��P]��G^r�_q��i>T��v_mY����!I^b���'����.�t�r'B����]@�3	� %��2�_\�IڻYn�E�*�e_�tڼXn�*���eV����k١�o�'mh�V�������t3��8ܧWyْ̬ڈ�.N�6ɨ�J�#BS]t�+) �v;��۴RC���tC��nqܵ�A�yĭÒ�e<�X�P_P�i/��.V���W�k7
hM�d�]G~�@�IC��+[�bٳ;T�E�ڻ/ť�49�X��3Â�Ŋ�±	6' C��S�d,�
fz�4f'�ԅ��f��6��t��b4�=SYD�@�kV�	a�}+r�Ì� \���aQ=3�,�Ùє������Y����il9����+���
B�+���Wt�J����Ô"�=�N���L�7ip:�a�:�a��y�붝�k�ҵ���84�\�gnb�v��|��;�`�� ����6��0l��+���뜑��2*;�w�2֨ƨ+3.Ϊ!EOL�z_r�;��NZ�Y�g5h��f�<-�����tST���S(dU����eb����]6��Ov��KAnZ$�١�g�wT��l��u�i�5.�AK��2R�*t��8etk&�\[I�:���r���&O����"�j��y�V��:>Wv�+ĝ{X�s�n��k������ub��(n�`��ygA�G�����D���Y2m����0�EGE��i���Hm��n\Տ����eGv��m6���<����J��h�V�e�8�V%�Ι���Ҏ���Y�#Ӷ�\m��m�4 V��>���^`REm`6����lv ����Σ�!]��v=�O5�l���̠����\����k#�8D�Q�Y&*���SA�6��k��P����-�u9����]ԮjSڝB��ܤ��·�]&c�S3-������hCa�*/�ĳ��[*06�!�t�]
���E><�K�j�*ev�t�s.+XUGr�۲�}Ǧ��4��̕Ŝ,gM"
���)�2���*i���n89ZB�5�I���ul�|�i�����~٦���J�Y�7�c�zʰq�L\���k��IT��i��X8��Mq�b�7}}PB��-��ΣPXU&�Y���{�B�%�����k]�˭�C]t�L΅����E��!+��M��E�SR��]�����LM��u�Vsb����>c�i�ͅ�Q��\F�*�3�@���jb��(��7�x,StY��hA9Gbe�
�뜳�d�J�y#z6t������'l�N��+��ma�8�hS�W�N�x�q΀[�)�\����.��WΣ�aw��u����2�k�u�����+`Ė_e�u�uj�ej���W���Al�!�δ�dq�t���=�MXէ �<���e�H�w�']�����Gu.�����pj��º�P먜Z8��V�ʻ�YA,�y|R��q������n���Gm�1L
��ɷ|��f�S1�Ʀ�Ψ�ytqԼ����]�=F����WM\��f��iKVGy�,^Z��ݕ��l>6Sq�n?���r��9�.�O�M����Q;v@�kA�tO��_E�:�����:��=t��L��΁�ۦ�7��G���S��onμ2�e¬ D�6cW�g�{�s�tx˕n[��9�r%�#��u01��d�O��ZU��	L8Q����Ypm��b�WR�g����Hf)�D_^v�:�,n���W@mn���*j�C�*�`1�����5O��:�.���;V���ˋT��[aW>)דh�
��@���V�rs�BrJ�v�)�����5%]����/uP�ܶΝ_iʜ;�����m%�k��\tVa�[�����a,�*ݛٗW.�z�]х�e�e76�aq�]DU�)�[](��*�+��L�\���`�����f�r�%Z�ō�>̝v1��<o��Y��0���� �6��_e�~Gc*ӷ!�9�N��v7ʎ��;�pf3r��=�Ϲ��$�����%�T�LB��V�E:��r�ó��׺�1�S�=D����ɺ�P�xΓW:� n�Yb�|$3%nP&�NW��arn#{ʐ�RF���bR�t3�.�Ȕg���邡�X5'���k�[����'��WG���K���u��Pv��Z]
.��]���Y��WիD��(�Y�Ihj��N�����jkh�ΐ#$�O������k��-�)�0������	R�Ӏ�qa|t<z{^4;�����wu�hF��ۭd�'�'N�׼H�������<�qL�͑�����Ӝ� ���ᅑ\:�6���X���n��.���P\�ǎ�#��5r����$��+&n�2�u�P��NQ�+�h���jBٰH	U�ͻ��N���f���_Eݏ�9����_#n�J������53{)\�����ཹ)�ϷK����f�)��G�#�����	];���^�2,07��.uN�E���t�;W(
;�]\kl�\a�6L�N��PI�];0)���p��D1��5�U��k�cA��	�)6X�Ĺ��;s�\��}Y��Z�z0\��Sk��4h��.���]n[�uA�sOS��OwY��j6z�n���-�q����:t�CC8Ze^��V�L�% p�Eڗf��K6��X�P�"]�*މ�r�AHt���IC��ӻ�,�{zK�C�ned�F�S�i�]R��Hu�!�J��(������j9n�b��^�s+����͈�9u5:�-kz�/e=wܦ��_	����e(-f�>,_R��qEaOk��Zu�|^�⛾�k�e�XE�k��x��V`W�ed�H�$y*V�ٔh�1]�E��p;�9��8���	<"�L��Hs���/���;��=���Т0kw��q�p�,mj��3)�0�	w�z�fCx��C1a�T�,�G+O
�F�m��|F�te)r�O�mc%*y׈t�z
�ہ�sj��M���i�� ��*� �dwPx^�J�sM�M,}�U�G-Dn]p�{.�\�}�t�`wFQ�i�SM�e��pm��7���Z�)+�f�ȋfUӻ>cA���jޭrMv��[�GΏ^���u�&����e�Ε{+/^�!m<�J���D��|�nF�C�NpK]��UN7Ζ�Z���GZ���7�qoG(h�g�7 93x����-�K6c�Յu��n�D�3J��Ju֜�p.Ws	��2�m��vI8���kt*t)�\&�)k��[[R]Z|v�f�.���w������	�-PЪ莫�["���Y�^�4��~������ξ-����Z���<|�a�=�ru��}�����1��4��Zu��3v�`�QX���9bP][{n��ے]����gH ��J����L��q�q�4�E���,Gkz��Y��)u`;�=�8FEN^��V�X:�2�V��k�>�gV�Cq���ܑ�(��6��<���Y�.Ӈr�L�d�N֕��D4���{iJQ��S�\��v�ьV���L�F��s��ZK>���r�蝨�rG9F����8�p�Y��Q��,)+U�88�C9�^��X�>t�:ⲹ���E�&�ΙceJL[��ڛF��=���>$�3a���Cxh+��㳲�@�v�:���0��]�1���a޲21E�ݬ{w�8�2�ŭH���\���]�����wif���Hi�XK9Z�`El! 3���=b��hb93�qT�ig_W1.�����`�S�]�R	hĹ�6��a8Ѭ�ގ^YV�S�5nFm+D�%p�2�N��$W؅�U���V�P�D)���~�t�	Z�s8h<�ݭ���V�6	
�l�:v�2�T7��Ar�J�ٖ�R7%-�U;;Q��w4ϜhaڰT	�[2
JS}��p���F��Mi��m�,�1Rj��N��/��[j�ʩ�i9R������[A�Z�s�^F�i�L����e�z����oC�*�dtH|�EC�36O�n�!�ݎܓ:S4n�:6�˺�H_gu�Au,'dߦM��+��-�[kU�����Q��0oCO�[��K�s30��sI��;��*덚=�O��
����e�X��(m=�C����V�(�O��/^�D�1��K����wck��+�m`�R����O B�Y��Y��J�g/t��.�����&D^�N�Q֌Ս�9�EU��u���W�F\8ՠ\�i��bTV^�hQ4��G^cѻL$��X�[���ah	I�Lq�K�ӫwSw%w�ZE�.��S���ky�grp��jvd�x���V�9d�
bVZ������=�colu`���eB���������C;�g&<�D�4�� JH��l����Ky��cya�o�%I��Hի�V�&�
M,H+��Yu�M!�Y}��t��W�V�sH���GP����j�w*Թ<�]��m�]�cM�-��Ꙕ��vus �r���1,Mr���ͥtb��P���l��N���,+�{f��T���@�1�yk�&lꖛ�������y��f�aihm���Eb��n�q�-α}2]bzj,u�����1�&m����2����%r�rh�@��]p�؅[��6.{y��yY�eF��gy��+6ђ�<e�J�b��Z����F廱�3I=���d9�P���Z(�z�H��P�]^�C�+&��D9�>/wJ���Whmq��WDt��䅎�5��9ہ峽%����x.�Ժ�� �b
�R,#LWK�o)M��H;cW
�NU��b������n(Рi�5���&���,��R�9Cn�:��Mi�AǍ��ڔ5!.g��0�PF���nt�������s�Z�o��a�O�����K�]��m_n�jӗ*IC{晬S���8�U�&iǯq;�'���\/�3�f2�<����w��jc�u�c��f���x�:��S�mv�{��8Yb��i=��Z*����JT�]
�CM]1{+��kG3�]�F�� �j[��k�6� ��[�a��]gg��f�n�oUK�d�j��2��
\bv:ǡ]䩡乊�㑥jr���`V)s�B�2�|3�;��]۹݃pRO��,b���	��,��\M�muE�q�F�>�s����ݛ������{0k'�Jm��1Ò�����kU+&�4�T��9ruս�-�MM�������u�Νu����0����3��K���|Ƒ$Z��w]�e�n�Tz�2(�S�gI��^�6����h����d�|���%G�T12����"�9��_eu-���u0֤�iV	A�A���
,,�QgeēF�^Z_!;�;��1vf�ܩϘ+)��^�1.϶)�cBHj�^n���N�:��S)��Gr�"���*�a�V0(�Z�c[Q8rw%	��Ft쮠�;P�͹ڛ�,*������{,���n�Fiԟd��Z���$e	\�n�<"��G�O5EwTά����[�w��;��R��ՓA�M��^u�1���7zjG�Ӑ�P�gqvp�\�>��ߛ���5v��m٤�\q�W���S	+��A�pXN�4y.���kt�(�m8�Գu��Cq�:d�����i�he�A��s6��k�ug����d�ʺe�/:IRmp`IҊ(�w8mN�Ԕ���;�@>���+K�2���Q���@�p�Yt�j=r��m��}�~��3K�Z��-�u5�gZYX�w��Mɸ�g`�r��h�AV�u��%eܰmR�� 9\t�jr�;w7�WMr�z}f>����kv�w��t��&�+��&�ɇ.�y��=p]Z��2-ܣ��LiL�L���
�Z�]����M����Lʳ�19��tm�p额�3:���s)����`O�e�ᒬ�����N��)�,m�Y\k��u���)*IO��,���0
�MYKV]��J2�ܽ�C���XE��^T��͎�U�X��.�#�,�,�wly+7��{҈��!�0���v�D��=��q��K�5���=/�|x�ob�M<3��q[WѱZ��P����t+\1Y*��,sC��2'�g-���=���zr��He�*�ЇlKq^En�9+�����2n���vR _����ڈu�gT��wG:���v1��˂���P�EԀ1S�ѳ.��V{Jq	.�>/�:���]-2X!���vUY58BD����J������J��,PwmM,
 �I�f�
����vtab��(��E�k��]�;����nQ��m���¹f��s@��/n��	=w��X���V�l.�?��"�[�1'��.���6��lv��P�i,�X=�#�TK�X�43{;E��W�z͓榬;�zU!g>�D���C4�OfwG�wQ�W5ut� 5$R���u
����s�nԙ�lr�@���q�&��o���R��sF�!#1K�an=�]�o .�^�e��� M��փ���p����\�	�TΤ6:h"�*]�E_���>�|�}�� M���Of~�UTk�ݾ~m��d���ƈ79��o�(��M�})F��t����Pc �4!,vV�z�I�YdG��#��N،����<.wu�˺���]��'atCA��׼���n�T홶��Щ���ESC9�T�qt�s�.��	�O���
��
��k.Q��V.⸾q�[�V+�.�/3�K�ς@�vr�9����7��v����x:��7����m���0�wcQ��N��_"�c*��m�X����cᶍ7C���Mt�x08��.�:�g��O��2Ҽ�^`LX�����%�y(���x^T�6Q;pl�Y82�d:�q܂��+�uf���`�}E�ti��}z^/��x7�,�ދ�GY7���2�@J5�ܲA���6���a��[�*-xˮu+]uĭe��A\��ٲ���6��1QU(&lb)��3EZ�#�g2����[wO�ˣ;t^���Q��h��3���K� �<Y���3W�y��>�"��T���x�z���պʼS.Q'{D�$_lmm��25s�%�w��������3y�YB�G��ƻ��+9Bu�t�t��V2�n��I����ָ��#�Q��9�ݯ4(�j̈́.&(G�Jٝ�TKr�\�*��ʑ�t6�2N�q�.c�nā�e�,��RA�]�3��$�-!Fu��S6G��~���^��;ZQ�-m�V���O�Z��QF�E(0�J��.[���m(�j�˔��S2�2��%Ģ�)��Z�TV�[e�s*"�Ycr孰�UUEb���q�+��J�j�emj*ܦ)1��nKm�r��e�0WV*ե�����b��cm+Cq�����X��f5D��Z�����U�r���1�,���j�bKK����$c��1EQ�*�4�Z[U�ڭ���DX-�6��D�f)F�V"�+`�nb��̥Z�KmJZr�2�ET)E��"řh�1,E�ˆf�fT��d���̘�Y�fTb��V�1�KmV(�En88��ڈ��ヂ��5C\��1(ƴ�jփl���[�-����)KD��l�*bTQU-,�E�b�r���r��6�[JYE����UEb1Q+2�Ƹ���*(�T�mW`bfQbXթVѴIZ����-TfZ���J�P�@}���^c�7��8d�����}ԍHU�敾�m�{�j�ϻ^*�֮2��ܙ0�8z��E�=Âxsf�J�6�ﻘ��!X�9_�Kq�o�ˡ�%tL:�J���hV�"Mrg�
�t�<�	�a+�7���6���wT/�傞\,J�}������:7F� �׮�5��v��U���n��&qV�7�}9L5�~�V����*�&B��0���"=�DҲ��;ק��|��'�<b�R��CG��=�t��ޘ)X{��8����伹N�~��&ӱ]�k�gC��p��ń0:�"��:�F�/�&h^d�E���7��K }�����eK��TlI�a��m�C��-[ɏ�| �9�Z��B�/��9y'��}}���X�ќ��:��wg�=������cs�cJj�Z�M�;{P�� �|�g��i��v��D���<T�;���=F�:�4`ܾ-��;/L��#^�e�}Ә[݋r�qo`��c�X�����R�g�HV��#�]�Vx��"X7-����;�Xz�	��uh�S;��!y�A�hꭩ��!�:�OA�ſq~�)zа����D��kif[����c�k�>N�z�<��H^�84vt��n��i��Ԫ��<R1���[�y����y�:檼M�&�lL��s�6l ���e�� �TɈ26s�͊�ov��k��t�iZ`S��һy��K��fo,8˲� ���}�>�n
�u_Vm6���w̦�NeYש8L�JW=Z;,�V+�f
��2�"�k��X�X&�0�jr��C�X�yv��oeͼwۈO�B�l��8h����x��xĖ�-TB����XYȦ����~~�;kɩ��%�5�6���v�X]H���A33�٫�����ٲ�}Q̾-e1��#�Z���v<��
�Y���%K�����˩���]sM]��Wz���z���W��NK��C��ü�oý�^�I�]z�C:t �vf�Vn����7}� ��5�JO˰P�z�҇=)r��S3Ǽ��O�����þ�u�zx;���:�݄ـ$���*�)^]���ܮEᲓY�t�(ە��.ެ��g�g�jۧ���~����q����	�µ��<3�Jx�;3��V���Im���J�:��{�����Sw1���5�JG�~�w|�K�r$Y�����_P72����PyVa�~�*���\`m�%a�*ܰ��%y�K�GKU�]ÏԼ�!����g��aYi����1䛔wx�[o��h���C�B�ǄT��{�@�٠<p�k��I'3@���v��d�l�D�wY��;��h"mZ�b�Y~`��#\�;
�l�6�.&pp�z��wVY� �(�t/43��ޞD�(��ȱO��)2Z��/�i��eؽ�b�2�{,��2��ս�I����{�꿷6����9�d�g�����LkL�� �{�ݱ�C�ґv���3CgN��3}C�Z"ӹ����2ӓ�fK\��6d�Vb^��T������l<v(6���b�ꗙ���=�N���n�z����+�MX���.�Bc�«mL��J�AB� ��΢�X����p�JB�es���Y�ǅ�w5x����qQ�{R���Uq�rɡ|*fg:!w�{ �7�'̬ԵO��B`.[��AcZ�{T�	y)�E�����B�^��r�f�^�K��#�<O�2N�7欱�Wr�0*�P� i=B�:so�3]�S����j�J��˘��9sW���G���!>��X���a�G}0�Ҷ��F�Rq�)s|����g�F�
9�X�L���^
zǻ���9��Y���ߖI[_g��.'/�Sӄ�w�a�޲a��D��h���A�y��?&{�:��hm���!QEO�)�b��)�E�*]���0S��Kլ�b<�1ir���ؕ���i;-IR��.šz`N��gu+�� ��J�%��|pGY1��|�n)��`p- v��4�HL�70�<!�a��r�ۨ�(.���eV�WG��6�M��Ѹ���G�O���o�?d8p	�P��#C�%�µ+�)�3G^s<axf>j�b�����T�]`�P�~��Fǽ�4�Cv�\��(�}���c��2L��#�6�_�ok��f��Ml�z�Xsz]%a�axe�$�G�����o;�{3%��˶4�\2*t���9�T�i��7�	�j��'����?j�t#D�S$��D��ʱ;�Vm��}c���~9�ȰeS�G<+�Q@��Wg��5��jrqqV\��8�a{�53^�����j)�����w^�ǩؤl�rݖ|w���@T���%JB�ŀ��[�=����R-/c���f8�!W+�jz~f���=T�:Y,�g̗%�<�};d��"�^��1k�Y��O)���Z��{�7�.i�bz\;�>���b�(t�Ғ��e.X��
�)K@���զ���ް�l��\�]ح�f`w/�Rޡ�|�y�ܬ��A��W���Pd��]�N�Un���OzT��Wl.i��T�g�nn�`�j���^��ʇ�VZ�!�}m]��-04k+sB��N^�yX#��:�f�XZ���f�o=���bW�q#�����P#MJ5b��*f��y�+ V�"7�	�;�)�;ʺ�/�foJ�elyXe���#�A5��["�\��԰�J���th��4�2���JMs�R�D�jJ�U������^T�������J���N�fJa���j��Q�����;Ze]��;�{{y�ݣ�kM0m.!�H�j�����;ip�e�zI�l��w���J9Nlޞ{w��6*�e��ĳD��Dl�0�G�t
s&� �z'��c�����:��v��u�wog�<P�����g�2� s�(��T�kȠ/yXs��=��������i{q��[mí)u�~iŚ��J���S	�A��@��H��P�B��g.G^5�Mޔ�W{�j�.�9�ܟ$�}�l-h5#e��ZH+/13�]:�������/,=r����>��O+=�tf|�(^|e[D�S�<��v�\�0H���N�O������x
S��]ȅ����E��23��J�{��9�(�W�	�7�e[�Z���ǹ�z�֎�Vh�c��&�2��9�tF�xy����p]�j�6�>�Z���Cu��T��W�aQ�����ǥ�3�2��\r��d���U��j�s�/�o��<�uocwP�v��3��Z+]���X׽�~h�iIs�H;o8Q+J�b�~��f�v.���
�������ۗf���nj5�����O�t�kmN=�>Sq��]������l�����Q+�Scf�����"#$��B�z�E#����j�$鄛��t�>;ZzX ���w�ͷ����'��ˏ��rQz_��K���|rq7��*�n�\�%���w�={����Ûn[�~���'m[�Ξs��z��]IK����]ƅ��D��f޹a��5'�xO{��d�"מ�mq�����1P��ͮa-�Lu�����;M(��g]�jZIAӛ��{�z�I���-��:<Xñ�	k[)ysglo,��utv{�F��'�y6_\�u';���gi��<X��XC��엫�|�S���7�j�Y7�^9�l�y9�`7��Gw,Ȉ�0K~�e�}b���+��K�ځ��ӱ��ό��\�|�͗+��L�l�]u�nqY�Ί�ȟ<8h_�=����v^�)y�\�9+����T�����p���9�g������zX<�к�Z����y�(�돥�:�1"b9�6ok��K!�.�۴�v (�کc�+����f`��@��F���BP-Ӿ䔏��Y�17e����:���<�w��Ďg��n��>�oˮ׭ج�{��z
0��=�S���w��(���=2?1=ޮ�tl׃s��������XOf����"w�n�1�r�B�N��G�Nvą��ϝ'�m��2�w��H�4�Ӈi�4��OC��������z�_�+����,��>���>�S+[��o��벜/}Tymp(x�H.�(|��՛P��}^��'~<d�&���{������L�d���w�P}�.>�~�(�/�2G���^o��$���cG�6��d��m��<j�	�gl�ۗ�~A�?u�n�x�3_���lby��WN̡�i��B�}l!Z#������n�uZ��V:z��b��E{�,o?r�(v�v�L���0\�F�ݛ���p���3=�8���t�\~�}�{��v�2x.��N��EU���_�H1�%�4�a��㺨\�N0;��Q�{��qUbz�2���J�Z��GcUu��޹E��;%g�zA���wP��{��u�Q乌I�Lm�\�w��Z��K�����қ���nƷf�n��+ �b���6�s����#�~��s
߼����
s>bL�2}rk�s��;�K;N��;\69L:�<�����h�δ���[֭t~��=�?oV[���;w�V��!6���O?_>;����@!�{��7=����!�s�k���r��{�L���<��͹�������>�����2 �vߋ���e��y�xډ{�o��%�d�w0:�Z�]:�S�͋���N�b� o˼ӎe�e����z�w��xI=�Ġ앬�����~�;0Ԝg����ep䡧.w콪~��|e1r��'���F��������f�^0^�@����ÏEI� ���/R��1r�}���^ಯ3�o��q�dO����D>��x���G��s��<��xkqt����m��L��Tx�b��C����}(R��{;�Й�]�ı���ؾ͍+|�ʈMpn�<"�d^\ۺ�J�+�5W�IR!a�"hD��^�V�3�Ki��;���I-�u]"ᰞ�B���!�8��R˩���6�c����7�)JNn4V�PW`{��Rk��Y�Tp�vk�k�{��O�)�������b'}Ԕ�J�":^-��CHķ�\_�d;��'�B��;}Υ�qP뙷�G��T��Ϥ��>~�����H�O��q�azY~3��n@���]���R�v+���e��-Թ�vw�I;|/�+2��ƞ�Wʼ�e��s:R\ߨ�2�V�����o�_ΧL��=����v����
��J���o�uoK\���]R�Z�
�������=�L�6q{����}�'���:l�+�C��+�|`�v;	s�[-_˛6<����&���kwm�s�ts�l7�|��������u�,�:#x��떇:�or{�S��c5�Ͻ�Dw����<����;�v�tB�\���*/�^��S����_���=�)<��/,ts6��W}2]���"Ƴ�_�|����:i{}���KZ�R�'c���pN��+�$W[K޷�^�͑��y�ʣ�-Ų�wVi㳝�9��\;#�0�f���*�a`�_��'J9�Z7�y�NϺ�����=�A��1�릯�Z�.��3
2L�o�;I���B#X��d��,���10\�5�枮�9�.7��̫���j۔k�����(iNT7�K�b�{�3�C��;���G�S!�).ͨ��J�R��_�z����]�i�Yޭ�߃CK�foDk���2��]�epyu�ȹ�LRV�����N��X���v�xt߸i7��T�Q��+�J�}���I߾m�o��׼!����<}�ŉ�0}��z�K�U�<za��~�f�����·�/t~�����mT$�_��{p��J�ǃ	l�o����k�Gj�c�:�ꔸ����E�~>�/��� ��Z�+��4�>8����x����&/��cm�u/ٲ=Ϧ�����o	�+��n�s��sq���S8��i�h�_����{����=]e����&3�� s�{Ut4}��/S��˦:���Htq����6�}-'m7v0���=3�[�Gp��_��~���o��yg�<��wR��w� ��']���7��/,(�[�����ΩJΌ�p��Kt�)��	βIٙu�h�Ř���4�`v�����ӡ\��7��\��#�N�pݒ����K z�mu*ܫ���+&��+�*��MN%7�/8Ӂ8��7���\�;r�݆�#�%s/+��ůk���
����,)t�V!�wFí*�u8�I'�b��o`�����$6x1M� =�6ѕ|���ۃr#��9����wܺ_]H�v\�(p�3K�E_#��oh�}8ô��^S����-�j_5x�p�OD�fq�cD��^�TZ��]������V��k�t/1Q�:j\:��d�oU�W���[�;��BE(>=5����m�s���s�̗զ�A�
�VFC�ϩ�ře�,}�u
���-R_fV`����՟:mes�4��rq$�5���d�s@9VA@�0GVZ#GV��{7�+��x.lm���4h�&*�@	<�wy7��Hd�ZR،.�8��WI��@!��0��+�rե\;v4������򆓆���������8.��V� mCU��g�����=�qX`�	L��++�=����ݻOfI�����.��=O���J�:�%kUz���-����J�l:��J���^�� bxMrⱫ�2�S�N��Ľ��o_ep-(b��gՏvr��<���u)t�an�7X`��ݡ��D����5R���6�)*�f���D�P�6ol�Ft����&L�ӭ
�5�bE?^���$�A;�"���d��O3�cwwIa`�=:�l�A��R�Cϖܑ��^$�霺+�e��;�qT(>4�Os����H�$��Ӷn��#U]��ͬ�h�oQy�k����7������z�S�7.^��<q��|�j�{e��)����@#[��h�
u�l��Xd���i�X��O3"]cV3��(�7A/��Z]>���!Uf��;��[����l�#DH��սhXQ[�;t�,j\s��gf���.v�[��s|�������Q�vl��{���Mv�+sq�N��9�[���e�7oN�pCN��"��*����d"�i�y���d����6HO9�m��cw�ȕcU<���J�×
�i�d�:Z��S�N�jf�P�g�E��:~)݌�7Y3��tu�E�۫�
'�`�vQ'q�Ԃ�W+{@sSZG>45V,�� ���7J�R�A9����M�
(ZM%���n��T�W!�+q"��I�.���X����.0t�hs��'V19H����QE�r��\�&qQІt2�u�Тo�.���9Mӣ���HTM�-�9�i��s��̏B7ݽ��*L0��)�)���Sg<���@�W���kVi-m�1��R�LyҬ828�S�$�aI#�;� 
E��w�9���4��~{\����>a�A�	�Ԡ�@�\�E��\lQQ�X��emhQ\��EY�p�Tr�E���csH��sRҪ
�2�¤T�1�j[erک��Q�e�.5�B"*�Q6؅iiW.0�pLQKk&V��\n4P\��D�T�Q`�J5�؎\I�f8�!�����P+R��ȫn[�-�R�QE��2�Fъ��3��dRT�*(Rж�q�吹��Ʒ�LK��b��r౔K��c�Z�*�Z%E*V��b!�l��h���fZʫhT+V�����0�DX8ىQeh�JP����(�ЭKl�m��\J���Kj6ʕ��b\[A�*�Vmj�e�b�T�X��(�ee`�l�hR�X,�iR£���F��b��1k�
��72V8�(��Vb�*Z-�a+�%���3TF�AbEY[F����!��ܢ���"9IA�&!�d�"ŭb1j� A@U
%��}c���:۹�ج|�2��ՠ�=��wyj��r�]�Q�ײ:"��v��|���5}�2dn���r]�k%�$N�|�ʹ��Nv�������,P:৫�-���ןol�w���֬&߰�{�'_�'<�����;�fW҈hܺ�O����W�~�lS�>�F��<�$���9���y׃�^��h�j; ߹5�lj�m׾��c��o�bw����j^v/ن��t���S窱���wm��%;%}���U��BY�>2�r�<��� ��N�2�{��=��s+�&��XxJ�Y�^����M�o^+ �t.1�����F�9*�rؐ�#>�t�vv4x\�ƌ�Hf|b��ɷ��j����=�P��'���F}C�R���
ܮ���ڻ����7��޼�\�Ͷ0k���ibO=8;���^q�o�wr^�vF����g���_mɷ�������g�&�+�k��e�е��Cl��Ĭ�8W��ʔ	X"2����r��v�����n����H5��\��k�7���P�>b�v�Ex���03F�9���
�9\bB�Zyj�VABQ�n��j��/6J�Fl,����՛¬�9w�/k��7��(�N����3�Kiw��x԰�]�����&=�v�0m��=�a���+TS3ñ���a��q��/M3��w��Zr�Ws�M�:�����=�7�R���$���+3Z��������(t�W�Nzn"�׫p?�����:qq�}�{�mڳ�����=Ϸd�۪�NIs�[,Sv�'Ɔp������9������̬�O��5	[��:n�6xq��v�b��Z����s�`���6�1+t�=6ZQ9L_�����6�m�&X��Z����M�g����߈�~Ïy�Mx=>kK}L88T��
�n�;�ی�T��y���E�������-�ǭ;̀-��ҲI^���w0:��n����bcT�]Ɵ	'�L��.����5���ǆW{$5�bI��tN��؝��+���|��\��[M5���3���M�x5i���Um0E���OQ�		Ɲg�\�{��z��8��-�u�E���r͵�[����s��{P\p�ϡ�ӱl��n�f_&��6���+T�K�TX��kZo2���I{�U�Fw1���X7���&�k�w푗O��:H�L\��$8�?<Ş��+`��������_q��U<�c���7�5��t�X��}�e�U���+�"Gh����,{�3�{b��L~�ۘ5�7����}3�a��!���%�>$Nb�؊ÔN�,(+�T:oޅҟ�O^i���s*\��3ͺ]E�_x��%.0���c=sƣޚoZ���v'F��Ϊb�lfۖK�t�����쯺ˬ�N���~��F����^����p�z�7����9Υ�3���N�^?33��6�d���sGMb���@��l��U��`g�}P�t�?
��|�P�bnSYr��|y�g��mY��{:��}O���,I�p&��V�z�&�/o��Ϳ�z#u��u�����ϗ�s�^��r_���¬͂��[~�8Q�7�ֵ���eC�']v���aP��w�h��V�<]d4�:׶��ཨ��-Tq��՟ ��y�^a�F2��E�Fa/��5��@��݇�u�4�9C80��#��ݔ�9z���Q�{�jC�X�����6{��p^N�c/6�읙�>�gh:!o����;ަ���a�r���>��n������X9�T��λ��t�7�4��Q�|�I�^~���5���o)d�_��x���9��K�ɒ�`t�=�W�c[�v�3������Ϋ�T��K�;,kq�Q�2����g�'��YV�����x�ل/K�w��>]w�\��)����E%��{���{%6X��_`r��9�|�H}X\�5�M�cgAw�LmdGz��>]&��[�����Lo�y$�@y��K�w�\7���ԯ��k�&�}�%t�7�d�<g�P�$��5݆�6�tk��$�&�o����~z/�Wx��i[���4�~��?}%C�>aPѿ��$��ߘq���sěI�*�xB��μ�'<>�$�l�z>�N�8��M>3��\����>�G~<����7ӿ��
�������d���<=� z�d�߻�OP�7�Aa=C~ӌ�J��vv�Ԟ2��v��2ty��$����d�o��!��n�����/�ޕK���|~���)C���;C��!<��z�2m�g��=C��A{��	<C�h>�N&�'��߸q�iP���2{�'��<d�:�G����c���⽳��)w�8`��G�WgF,�i��Hk�k�S��{�3��{=K��Z�҉�}�����"�;�A� �O{n@�M�
�]bFHu�"�%8�k�͈��V���EnT$���!kn{���r��.��� y|%lT�ms���^��-��ߡQ��?�D>����D����'I�m�x��CT8��N�}�2m�S��OP�'�ިM��C}d�i�x��y�6��u|�:낼<�씫п{:�@�[�q��?}���I�$��k$��`t}I�Rt�lє'��'�l'�*t��Y&xP�'Y6w�I��eMo�	��a��5���7]��Y��ʬx\�}����ɷ���l'o��u���m��Xz�whx���B�&2m<2��=C������'Z�l�J���u�O��3n�~m��y��#�#�~D~�����s��8��q�r� ����M��'Y>9��l'ɣ5�T��:�<ed��[�8ɴ�S'�m7�]�Λ���Ӯ���~�:ך����c�<��'�X����l����>�
����ϩ6��N�s |�'l���!6ϙ5�d+$�7�J�ԇal�
ɴ�����]/���5z߿}m�����:Nad�I��k�&�&:ϰ6ɷ�C���M�s�{�8��I�/��4��'ӝ��$�&���$�i�G5��'{����ix���Mե誹���@$����� ��hIĜf���N�{��,�l��xd��!�y��	����6��	��y�l�����Rq�2x�OXu����W������~u�}������:��(N{x��q+'FP>I��3XXM�z��Î$�g���
���҄?}������a�|��v�����>�}��y}��'�>@���m�d��;�x�zɩ�`,�ho�%J�k�m�d�+%I�2}�<�XM�z����Ĝd��7��&�gY�;���;�}����~�i��x��)�d��S>I�s!P��k��!�&��:d�I���T�&ݰ��=�je�l��~f�5Z>�«�!��߽�h�S鉝qʎ�<m�n���U��7}x�~5����j�l1YBS�\�[(t�O���fz�?/��γ���`�,d�]rw��J"��*�A�՘/��1֐7�5Jnw79�0�v\�v;��L��8�A�1ڻ�{�~=��w=�"j7|은����_�z��������M0����$Ĭ:��q�N�[�M$�
CS��T6��9�B��'�����i5>�$��&��,��� U_�!���3���G����Q�|ͧ'v2z�t�'o����O=� |�2q�߳����߸q�c�,�M��=�2x�l��a�7�*Ou�t�_~��x�~>����?4�K������a$��'o��MI�2N��2q��T�8ɤ�a��&ؾ}I<C�8o�8��1:7�d�+!�P������͟N�_�S�O�ON��i�M��P=d��'̚󼒽�����e���&�P�	�8��a�a:��SL�IĞ{�I�d�g���8��S�����ꗗꎕ��?͚,����g����J�s߰<a�O_Rx}`z��'G��c&�)<k'L�MXN�$�5�m�x�:Շm����C��A@����� ~?}��r�hH;?��{�K=�Db���Bi&����=f�O�߰�&�����8��O�Ry�����d���N�>k'L6��,��铉�,�$�*_ؾ�H��5����i{��o���9��$�
}�)6��Vro�	��C[�3L'?S��{a>��q�������|�8�5�VN0:>��VN�C�R���?}��������=��^I#G_��L��:g:��
I�o=d�V���,8ɴ�ѿ0�@�s'>�N0��2m�'���N�R|oY&�M�U����8��~7oC�sw�nx�M=~�J��N��)��'YLI8�����i�c��!�M�`k��d����$+'�k�9�&�:d��>v�����~��r�����4����>���s��d�����Y%a�!�i�&�XtZC�8��є��Mu���I���7����M�q�yd&n�0}���b��#�����xD6��Wvf���,.�����sWt#c)z���ɾۧ��u��f"��csLQW�[y�`h�V�:�5�;�7����j�B]Մ%K�x
aZ켌Q�Z�|�q�s�vR�ħ���v���Pǝ�R,71��Sn&�� 1�����������l'���M�!Y'����*
=��*M����>I�N&��O�m:5���	�w���'�`v��?X��
��t)�~m���C��Gӟ}��2v��N���q6��M=��!>f�57�E�m�d�(M{g�VN%d���6��k	�'Z�!�Y&�3l����X��~�%����	��o����9���$����4��	���d�;��I��'�:{9��d�s�$���T�&ݤ��%d�(�����ٽ�ߔ�� ?�{gN�k�?tɉ֬<�O=a�7�+�&�׻ɶI��;�s$�$�o0��0;�0+�x�����k��XN$�t����ꎩ�7�#�#�A[m��3�\��bJ�����O��M�;׸|d�'����vɦ�{Τ�ʇ_s'q�l�1�h)y̅C� O����>������u�t�u[���{�L�Ԝ��%ea=��$Y>{@��N0�{f���M�����M������'l;=�8�c*���,���P�~�	������~�{���|���i�Ԩ{�Xv��u�L'���/vI�{�,�=��k��N�S�d�!ֻ��q��I��SL�~�_���@D�z�}�ު�Hy���+�_r|��bs�p��iP�>�N�m�Ԭ;>�Xx��W�I�O�d���l�M=�t�e��'o�:I�ɮ��~���B>��&�����MngI_k�a�O�^}�$��h�xq���n�$�+!��2v��O}�xn��'��{��m�G��5���Me	��&�S����~D���ʗ+}��_����w���|�u�z�2z���5�z��6���&�q����L��w>�N$�+!�)�N2x���TN޾�IY6��FQ��?}bQ>=>�YO����Mr�*�Ք�nѠ	&rFƙ�1��t�������`�Mx��n��z'��o��sz�܋,�p«	�]j�,n�ׅ�R��g�Z��h1��D��(�_,�?�{��߮����J�ͮ��un[�I�-��G%��
�ͽs��]+��O��I8ʝj��,��J2q����=Cl�J��a6Ì>��&�N0��2q��,'s�Ì�d��'��$�$ҫ��B{����(yd�a��M��߇�Ɍ��VN�|�d<Ld�<�>a>B�Z��
I�z`m��R�삓l�J���!6Ì4o�8��8ù���>���G�O�͛�4I�"�������5ēo̟��d�2O]L���!հ�+'me���m�2�$��h�È,'�F��m&�X�y'9���HVN0���<枯������6�ߚ����$�%� ��ORw��I8�ɣ��VI�7�J�ԇe��+&�Xu-!�I�hˌ'�6���I���Ci6��޼��}�1�5������p<d��ol�vB�9�3��O�:d�}�~d�'a�b�m>d�T�$��o���a3�|�d���=Cl�ML,��f��V`~��?XW/�G�g~�B�������C��ydP�'>{C��a�O�M|��i;d铮Rq�d���\�O�L�꒰�C�o����2{O���B>����6��E�K�O�w��9ߪ�
��t�0�N0�:��6�$�k��6��i6���a�I���L'�s�I�OP<�2N&�=a�ww�a���x>�5�����-��t���vW7�� �>�״�'l�:�m��	�OY�~�q�I��d�}d��y6�q��9��q�o��N�>a�9d�t��~�X���qW�ڣ����3��� rN}���'^�$�RL��%I�+'S)6��'�XM�0י4���M���
퓤7<�'�&'o��N$�y�'A�S��ݛ}���z��g��H�~�:�$6��5��'��S���$���*V�_YO��:�I�OY<zu:��&����Ԛd�C߰��N�^_�P��y�<(���V�M���+����k���5 ��a�]E��7o'
�[X����
�u%a�23�[���C���.wz��/$���⁫�F�=�y){/���ް�&��M��\1�D�c��t�\���26{`�ˎ:?+���/���Ӻ��'I�)�&�X��B��O��7�*O:7�:d�a����$߶E����P�$��5݆�6�}���Wo>�������k+������#����20����������Y&'F�Ì� �9���OP���'��u�I8�����$߶Ol�Mu��{��W�_{����{zH��������0�4�>��3L���O	�y��'_wI<C�o�q��o�8ɴ�M�'�>I�*����N��x�m\�~fv�)��ywߜ�˙�܇�d�i�,'4�����6�wCI8����z�2m�~k$�2q��I�C߹���I�;7�d�T'<�@�'�Re֯�_��w���y�}������d�����c'lyI�Rt��k,����IY�I�Vt�q	׵C6�ɾ��=Cl�J����N!�����I�=��|η�-ߙ�<�y~���]}�k>��'n�NO��̜d��O]�d�:3Y%d���<jN�m��Bx�2q4e�a>aS�P�$ν08��Ma�I�T��{~�wߙ���0���q�f���>�>�����}�чf�2q���	��'�k$�$۬�IXz�(x���C̲'L�Me1�z��	�]�ϻ�}����u���~�������J��a�I�*k~d�d���~I8ò� ����N��䓏̚�M��%��Rz��Z2�m�N���d�l�ή���߳z�|��}�|1�|�I�Xz�2Ly����iX<�hd�9����a�\��ԛd�'|�@��N�;��Bm�2k��VI�.����m�k'��U����LS�N��� ��l��'ɬ,�ԟ'A�r&�&7�d�� 6���y�m�ԓ�|ϝ�v��'a��_�v+�?~5����'�W������lx�6��Oѵ߻ޗ�tnղ���/�N<+!I��P�Y�}�OOk���gmSЇY��� 6��i�M���W�a�(�B�ʆ��D�I�r����'A,�ޒ�]�R}��o=����ec̶�Nn��˹�=�+	�O:�T&��+'�,:��m'̢I�N'���}�I�jw��q���^`v�v��s>ɶOM}��a����/TLn�Uc��{]���^{�z��=a��RO��Nw��N!�oXJ�����%d�VN���M���a6��y�rq$�5���}d�wM����y��/e�?z{g+~;��~������2i'�����'�Y��8������6�F��T�'���䬝�I�2}�5:��d�;���p�� r|�S��(*>����w�����>�0�Ͱ�)�d�9Ld�'h�2�<Af�̐��jsXt�8�F��*T�=�aY>{@��&�=d�T�y�������5�{�:׹����9�2v���'�{����i����&%a��Ì8�t��2i&�R��B��OY��'i7՘�m'��]Y&����.�����_}����_i�~�N�92��	������N2��>2i�{���i��v{�q�bV� �Lz��8�h)Ns'�6��V�xB��>����na���W����N�T��}��<d���$���	��'ɬ��$��;a�&�5�';I�{�@��d��w������ �LN���>J~�c�z�_��}�����G�g︄Ç�<d�2I�'z�WI>d�|a;|I�h�a=g]�i��N�}���N$�O=�$�2q��]x�÷�7�e���緿1W��"���?	�d�VCP�0�'��8���OOu�D�M�5�'�d�iXN�$�L�l�ĩ�a��|d:I�Cۉ���{��Gy�˚�9����~���>�P�I�7��:I;CϹ�7����N2|���X0��oY%d�i>k&0�e��2q+6�<J��w��>��?�}Q�m �H�E��{q4ѳb���V��Z�6�Ē<���
�H5Z����k��νt�l|3wO=�{��Ѽ�<䒮��2Ѩ�H^���Nrz+�Qa�=eJ�۫2�;k4�["=Ks!mp�w�D�{KQ��n��|S	�#t� ��h���,y7x��o�2�ms���hTПrt�C7�ͣ�Ny�MˉZZӬW0ojp�4W;(���Sh�XV�\5�}cq^���c�܉j��%9|�#3�Lb�jP{�o\�;�pD��{j������kU��1�	Gp����t_Qh�q� Zɂ��V�� �b��H+D�K����2�x�.���Gud �I]�y6�Q�V�`��2�*�[W8dT�$.a�����r��,]J�Rԍu\�!Z2ޛ=��xn>˻�+�4u�̔��n����b��\1����������"^ I�np��I��e�u�S'\�q�9�TY8�3��ק�b�}��+%`3�����@�pe�{x.��i����E�<�+�l�٩�}���گ:�y�P�D�'n��.NV�^�
[�-�U��ڊ�}F꧗7�A|�w���T�z�N��2��;�5zFM�R�Ͱw9�k�Uu�B�[��U���6w�D|N.8^X�%6YY��c̗v>�&ՇcP�z��bE��3�ʓ8�A�0nv�oOD&�r߇QOv0)�q2'b�Y���p��R
�|�$h��+g��v�YZ�>����q_>)o$���霪#n�*
�E�w��!7ݛ���ٵ��j�M"v��s���}�!vV��K-V0�]衙+hUfc4�[�1�g�3)C�%Fp�"Mh��+"��Քg���v��[�(�e�<��OI�N��1]�̌2It@�I��v�}H�I��^w=B�7�ú�Z1i6sn����T�&a;C�6�����WgO�5����|$9W�\ d2-�pF�[ [;u3KB�h�7)ˌ�o:�hK2n��
����vb�v�����WJSL�&XJ���d�{+:�:Y��:�����U�9�U���3b�%+�S�z��5#��̺�A"�
Q��{�m1Ի����I��O�V(*y���W�*ٶhz�<��vYt���o�9�	�W �.�j����5��}�T��u��˫�qGf��W�5��T�R3%�/�cuh�N��ν�uz��ǃ�����Qp�;J��6F3�]����m	ŵl�R�E��:���Nd�U�ض�(���'��$�R/&Z�۹�@Ux�m�Q�僐ff��ZW�KB÷]@6]�wtt�0�qǘ���^V�{jh�k6�]C�u��8�u'E�vuq��t���RWo�}�87,��d+:���Z�M�H�D���+#�*āl�d�5���)��"y��֚�[w��8��r%�Mm����s-KR�k2�Ċ\�T�Z��qƥQ�Kr�c\�
�Ե�HڰPQS+l1�32��Ve�(��B��Y���U)r�#����LLDU�FTV
��=��ꕎf��uծ3�d-̅lB��KE�,q�n,bU̵\��oYC-�N`�\E*Vb&1�B� �4�����!�\b�X�(��AV"1
��V�AƥLql�+Y(�(�l�!V�oWET(�`��b*��V����+Im12�8X5���8��J�P�PUFEb�!m��m��"ez�10LES)Q���0rW)B�
�+"�Q�P[�cW-�κ��[E鐩�)KU���X,W3$��fe\e�Qq�*�WX,��)P�X�*դ2׫\��D�Ke+�"�^��Kim$���U��4V-h��)+�Bڈ�"��QX,Q�(�Ib��m�uL�X� D�=֝�4�궺V�MS�;+Ohؕ�{wP;R��ik"�ͱ׵�êo4��(*�j��{�Ҕ	��������-�g������~�@�}�]��R|ɴ�ѿp&�q�3L'v_��&�N�9�O�;�k$��q��d�����=J��M��=O_/o���g}]y��[�ܐ��2t����6�uC�����8�����E��6��ߘB�q��N}d�a�N2m�'��p�N�noY&�M��>��}�w�}��������g�{�+���v��T��c'�I=Cl��p8�d�߬6ɴ��H��'���rB�q�s'=��'L��s ��'l�ϻ��z���o���z���w|9$��O����i�z�+Y���*N �����N%J�|�i�^�|�$��ϲdߖC���!���H�}�$��`���_����7ҽo���Y<d�'}�q�'l:N�̄�4�ά+$�<�Y%ABd�ϐ�6����>I�N&��O�m:���i���O��e�Y�]~[.:f��*��=�>ܜ�ʗ�L뿞_;!�	��8}*��X-���z�Ξ�{�@3������2_�I{R�h��o�g�<����N�3r��+�)kYU7_c���뱭�2��+�!X$�����k��<����=Q����g��X\�����#.��؍�< �b�������wfz���6���ں�����rp=&��F�{�sg�2����7�x���CE���P�W���Ac��i@K�^x��G	R�-]͞$���ύ]
��6,L�sR/1���y�`�S2B��Vn��IW�˫�٩S=�)]���=1�G�R���exw��K�}Ͷ�n�M���������|���Tŉʈ�V�xt�}���kX�]�|�R�~��fA~ox�;�*Μd��T�G~<|��E��;�t5��֭P�`��,׭�>�v;ck&�����7�Li�-0����?�j���c��9V���/}_[�ួ�fۖ�~Α���v����҈�b��^3|���3M7�޻�h_+Db�Ûn[�s���$�ݒ5�#^���
��\�c������4�z��}l!Z7�6��S�Qҷo}�@$��w�9�����Vu���]N�ؠ�_6ly�=~�a���Q�ѽ�{h�m����y��,�Gh����;��U��u�y%k�N��_���w������׽Q�W����7���iݿ(/{�NU�t�v�S�޹�I�.vp�:�s�ˑ�T��e�r�T��'��2���ypV��@�_d��J�L`�&���PL�]�kå�3:���Ȼ����r�K�e�
��R�9V�g)0G�	N�yW��#���.����u�}���q�i\u�6i�ȹPnSu��t���j�Y�%�\��W�=*��I�ض���t��y;���'�)y}���{X&K&��������k��h�=d!��K�U���;�;��'o��>����D,�N,Џ�b�{O��{X����K-��d���{��삛��q@a��c��ɷ2��&W�O}VGTB?�f{��tq��k���v([m��V�/��>�t�vw�f�0k�<��hl/�ɷ�rǾ�E7�	�/�O&�$�����_a�E�Y���3Ӟ�3�/\��[\{Ɛ]((��G�]���j��u�]�����~��՗ho�<}�����>�*����.t��,��}+��.R���'��r~4.J��S���_ye��Vԑ�r�~�T߯|�o?Ws��l��o4fw�~^�a>4-�� �f��m`*d~wD�1T��ΙH���1e]��K���v��	�R��rfᛊ���].�j���۫���ꘒD����pJM�<�_=��o��/���m�X���&\Ǯ�o��Jj]}!���VJq��v�ξ�3�;�"�V�3��5
?�Wս��b�c�����S�|Ԟ�G�U������}Xvvb��<����5���sp�.�c�y���I�>/{p1:�4w >,HN�d#R9��[Is�|��X\ٰ<�M�e\�u';c`}K;����՚6�s붥=��sg���}�S���v?B.	��*���O�ib�C��Z׎z����˯}E��B�,P<��C��N�77�������g�7H��{Yfe���l<1�I'�'.u�����.|C�^��c;/�ێ�w�0å��QD��Ջ���
���I���W��	Τ��%�h�%a��6=��f�I�i�mKs#<��I�.��u���U�ݹ^���o�F֯6��V��<ܞ�]����$�[$/������};�}�(�<�R=�o���7��\���^������Ok���v��VO�]�,���=��>�^j�� �ydIR�`L@aQ�����%�mX�w���h
�]6�w����7[!�aef! QO�U�4�N�V�ȡ�咦͛��$w�
�l��Yf09�C+epVQa��j���o]&&_:�wĦ��~���������a�7�,{�3���æ�>�����c�c�ۖ�4 ڗ��M؄��_���N�>�"Ǡ�z���u��ܞ�s�{�Ύ���r��zN��)Ii�^��x���:22og`�w�	���u0U���I�y�`����l`�r�K�|:G�d�;�S�+8�>Q�2�/����y�ݬٗ�S�8Hy��sG��I��W�³>?vQ!�N:{�b���E�/�����8lg͇�+��G���=�j�]��n�sXp��H�gX�n����;�^��rbOM3��5��Mq���Q������ʾ��u�gZ;�,W�d����G��^9��o�d�����&��RΉ�$���]{ӽ��M��N��x�S��'����{�Ȱh<����xǬ��x&��ɑ���v�[�\��{y�U^/�ۦ�*	[�\�,b��5|�Z��Pw�6�oq"͌<7m|�� i��cn��{vl�&@Q�;y��[$��N��"�庌���m����n=��͚jJ�GI�������xlK�����턥�p?UW�v0�~����I&��y�v��Ry�W�J�$��r�L�vM`�&ű�2���1sGI�ڟT��k�y���[�)q��6C^$���C{��y�o&����=6�X��S]_��k�Fz��#@t��2�)�}T�a�W5���������շN�	���怽7�"߀�����療ב��y���n�ĩ\��|�FnxS"��[�M��Z�����j.$zz�����m�@��;&==ed�k7��c�ԯQݏ�<Z�[:d{k�6j�})h��R������?B�����^[�K��rg���j���E���_m1�ײnXu/��3='��_���D&Z�����|T�]a{����ح��p�ۍJ��)�'t�}G:�w<�0�-����՗@wg�x)��Z=����F��i�^@�V��.�� 6�b˛�b�K7�M��7�����]2R��[DL���4�����Y���U������4+OXz��{�f�G��ӶnJ�C�;jsKź�j��]���C���u��M�SK �[S�9D�-�UUUU���t*�a}y�\�����v�³��?|����X�:��;�W4h�[��n{�zw��p3���/{p�u�;@:;@��Gc���{��K���:Bs7�R8�g�x��N*���������gZ"��w�7{n�⯲+�%Ϻ�Aʹ.`	��.vv�ד�UH�\�e���{НR�l�m�K�"|��_)%��:�������:9�RW�V�CGR[j�g�<�ν�n	�E����ԟ�؝��[��.2#�oxg�����Xޮ�t���)͹bPvJ�x���S+�C%��nzܽ���X1�
oÞ�^�w'at��{�Óe���;('���}{<zQ�J~�Og��;�"��kF=���-��B�lϨ;��m�h�i${qf�����p���yp��-o�'8�ϠT�8\�zpF}^�OT�0MW�\��������2��S�� �z��Q�(͡��B��%<(���Y��*ʤ�)���xT�ݣ)U��r�o'��ǳ}��;tn�\.Дe��/2�WaD�dYr���N[Æ�ɖq�Ux1u����R�C`ˁ6���}��{]�ӓJ�l�~�����n��ޅҔ>G�]���j�X�Ϋ�(��h�B��^�m;gMd>�7��Gv@�����K�����S+.���wt�  �&�F����'{;�������l�����sk�z[`�r����WCy��6N���Ve|;Ɲ�T��ж9����=��dߤd��	���Ǯ5:sR{���_;Vv���^���N�{�%x��hշ~�fK}����猯�N�����[��Yޡ�R�^���Bz��~gD3%����e��sf���6q�����o`}B(�̮��y����\��|}>�9_X���C�}{֭t~ϋ�=�k9�q&�ޥ��}�y��*�����;2��B�3�}���O'|$�w+9�j�jC\�Q_xڋͦ�=ˇ��:�K��q�TT/brfߪY�T�F}�\���$�D��u��(���S֯P�6���^����@ �[S�'�0�3�+�Mh�t�y�c�y���F6��#���z��oH=����7�����E7<qEF�;���k�v�u>�6��˜�#{���F�o�}U�Uv��ی�n3���������~σ��eI�%�N�CY�Iίk������;�u.��)y�{<�]���ndxe?HV	'����|�^x���Gy�me�9�xW4s�/{�l�vn=�)�lF�INS$/��>'�}�)�p^�w��Ԟ���9�4vPR��J��c��\ވ��}�Ұ��r�[�w�Y{~�fr��x����4��V@xt��JP�x�Ҳ��/W�%gg�R����t��<����c-�mH:�� ��s��d�V���KB�9�B����1#^KW�M��t��N����w����cS�b��0m�n��>#�d��efW�Ɲ�9���0繿J5���N�t3����\���I��U�^w�iY�0�i}NR��@ᮿ���[������Γ�|�~�MU�8�=�9�g+;�;��K�L9���˗�E~�4yt>*��ns��>�677'�"�G��n`�+���ZN�Z�y��`#2�bf�T��E7�&�0a�rp��7��r��F��)�#f����{�V���޼���6�R~�꯾����{4H"����K
����S'_�e�\ٰ<Ğ�&�/kn�Nފ��ޓ0l��������`%��zՅ�����I��ײj����<�p����s��H�Q�:!��p�+��Ti�h �lc�������?V̃37~��<��\��tE�����ٜ�^E��;s@�)s��t��N����x��	+$��v�	���;��>�m9ݲ�sd�Æ�}I��Z��=v5���|ew�Hk��s�i�_x��{�<3<���[d�=x�ʺk�����w��#]$u��7A��0�L�c�"���x@�a��wN��%։����� DM{���.��˿Z�R��t���Шk�X���)�vw��d�y�ӝ�XN����7OM��L.b��7�}�1�2[�ރ����_a�f�P}��������^$�M�	"�ܾ�2��9��j͊���\��l�tx��i|���H��B蘱�����R�R�g^�aӝR�B�G֯���`�_�{�(/���5tONG�{tZ���y�N5�r�xlovj�j�n��� A9}Ff	k�#�Hk5��� ��@3*�F\Z��w)�q<�nS�틯:�#� �x`�o.\�6��������ح�,;���*�ތ���f�CO6�nR�
��4ؒ�RSG ��*��b�p}����n��r�[nmkjC"��U r��h�4ͭ0�hEI�����u�O}}�����;�H)�a{���	����G%\{{�.�zHY����On�:��9m�O��e���i�v�s�+S�c��R[l�+Y������Yp�q�c8♑3q�,ǍÙ�ϓ M����]I`:͝r�+���=*���T�0�_K��e5�J4Ł�65y\i�z7����w�#K6:�2�����md3{B����X��Z�y�N)+������U8e���OL�wծl����k�q�����r�D.�!�q�L_)�^��nheq=]^�h�Y��2��p�r¡���ʻ�n���A�d�����lAYTR�em�w*i���!ٺXB����u4���.��KC�Q`빃j�R��}��]�.����m�C�O�G.�uc,�-�Z&ݤ���'¬ms��x.gg4�a�tY�w�M�u��3d5,�{�k����J�-�!`:m���i4��x�5��up%�墙F�%��$��i�K.��#AvL}�]Gg"D��#K�����#g�:R�fF�]���`��sp�벘vͳח%��&Iǔ�y��p�̂�uZݽQ�)M��M���u�s���W���FFE��r3�����C��IӇl��H[�L���2�j�ɼM%��ǝ��ы��S��M<p�R�o |4$:��ބ��9�Tn�:
��:d{}{z�����0��*��q��eԣNޙ�6�b���U��/5�+�:�n;��I2�ň����p6p�7�]oc2cx�X���ڜEm�"ok����?��Qvpb��*a��Wy7�
)"Ų�ӕ�z�w.!M8����Z}y;j�;�	qf�	1N\��=�w�X}��p=ΰ�И�sˑp�{�ħlUn0n�;.��	���3�@���nH��f�$�Y�6V,m_	��?��Q��Vp峝��y���gc�Д	��N�!�����\�H!]�Μ�����Z4�}yX7(�m]*�2�;õ��[��ɿ�J�h���&�[���};��hsA����9�b;4���h�
\�9+'+���Jga��NR5[�;�+g�P�&-��5T-�\!:���ī1���ʚ2l��%#�[�D�ɛ�9|�:��Ē��c�5���>TEV2�AQ���Eb-�X�,S�E�`�b1H���"1`�\e��,�DQEQN���M-�b��P��2���W��*�AbȌ�*V
�,�=XTN�Fڢ �,�,R�Ykd���Vui����*1C,�Q@U���
(�H�"#am:@��l,�ʋ�,�Lj�H�,���*cF��*�(*"�QA�DcmdEEƠ����+TE�R�R((#:j��#�dX��1Q�!�*�*�Db��DV"��UA`((���Pr�AH���"AQ����E�T*�Tb�ŋ	�Qe(�����"�cZ�r�EQUD1��DU`�*��ŀ��*��QTE��*���5�O��<��($�En�%h%g�������[i%y��h�듏�x)��.;G�r��t]LZ�=�q�� �.?�������}ɧ=VS���G��<�P}�.>�~�.3�ǹ���V���Ƒ`Y�z����Oәۮ|q�ʉ����}}�ǫdm��Կ`#7=&�FĮ{�q��N��G��G�藯����Y��(v�X�r�K��%�j� �,C�q}��.U�>�9���׏֬��4�/T�����8lg�������*{Pw��YNڷ6�<jOo�����;G�;u;Ke����'��Nfz�U8f�l��rg0=��.M��|�L�GZ>ߏ�v<;�x��g�W{gH��[�ڕ�j�lߞ9�����Ǔ�$�K;_:"��S�뙷zق�������޶\��̝�X��*�w\.u�����CM�2�o��2��ύA�!}�����J�����~
O3*�:9��fW�܎���Θ��{�sj��`v	N�@k<ON����;�f�;�Ћ>>��R���Ld���;M�X�.�_�����u !��tb�_cŧ]�R����w�����srV]Ww��Z�JP{��-�yL�'5y��m��ӻǼ6EJu�:�M�&���� u�N��P[8��Mgu7�5����C�m;�aG��ﾯ������^���V�����`�6P��ߵ�5�{*�4>�_���e{��[GI�~f	��9�Ҙ���~�.C��beGd���U��7&Ri���������nMz��Di�un[$/��>�t�ͼ����j�u���Az���@}C��px���'�n?�8l�zpF}���F��~�A��S��LX\��Y�z�M���C��
���oc9���\��F���:lWST��L�<WQ6�}��}���M�P������ �<6��]�p:�S����K@?>9	�������:�D�����')l+���	�.���:o��z^^�EηTX򭰸Y��G��ԋ��y܎�.�����:r�)�����x��P��/�gG�sR�h���Up=~�ێ$�﨟9\����2�t�^����=ѯ>~�sj�k�/_����oC�����f-�R��4S����TؔR������1���ަ3�o�`A�'�<P_�Q\�����*�S͂�,�ʈ��[�Kld�4�);��ާc�4��̩��g-��g1��4JT	��9������
�$��.|{��--w[-_˛7��I��e����{ǐ��kٺz�:�/�E��/Q���k�s�{֯���x�^�,i+�~9�=��x���a)o���	ܳ(J!o(Ϭ!үy;�;�{�(�u}�o�gby���S��z�z��w�x|�5�O>�A��_q@(�?6�]���Z^�'��pb��~rW�
�eW�Y�3P~�pY��mԐ�ֽT�o���3�kj9q����&ܺ�(��vKZ������9f�.}W[(gf��2����%Xr�����Y�jd�\&����n�z�WW�X�*�k'~���
o��^������n���wI*LA���6b�,#��,E�� #a��J�0ߒKR����^�PR&���>w���|�;�n>=v��o��oC/"�Zڶȧ�#��e`�����e.�;���Dɾ��J� �����	�� �]:��*�8�6�ͱ�T!�;�.]�-�yqڢ	�fi�2�'��'W�o�@oE�E��=  < �Φ3\���U�
+����b�u�']v�w�����"t26c��꯾�ᥪ�s�|y����҇ˏ���}��x���[K�N�4�,�n�K���=��6v��|/}W¸X���,:���͓����㥉3R��� 7s��_%)�WF�TYR����h�^pp�s��sG�Ū�`'���=�B�C��k~*�ua��f-�r�*n����Uߝ���Xη�w��)�����Vv���]N�K]��j�\ٰęGR��3�~�h�{|�ZN�.ݒ�I�3`�cr���3�d�:Y��hu��o1��]��=d6M)Y[
z:y��N�q�tBŊ<���w=��	\������837o��<�q���<��~J<A����<�Ol��δ#�{�^7�<��2���~�W���.������f�nbWs�ܑ�\����oj�{Y�s�3�z�L
\b.�RG��5,���B�*�$1*��>^��wr�����y2͉M�(o���#d�N�K#�p��ize���X`��b�#UwM�}�up;3��%�7�E��X3�&�6s$�@�ǝ�%��t.��1!��q��E�ʼ9zx��nO����}_fW �I�zT�4�?��I�|���d^܂�q��ޗ;��e�M@��~gɽ��`�ֺrإ^����:���h�I�X��/�����t{���ח����tm���pr�}�)�m��#ݰ��;����)Ϯ5�=��(m���-��Lzs�����Ú���oS"���N�g'屿K5��ߠ�[���P}(.>��R�=/��#}ڝv�B�{�U=�%��� �밻�'�_\u���={ ͷ/��_�t��xx��_�w���׶b\���������	�հ�h�^v�pm���>��/
����d���|s�I�b��ՙ_wg�yN6����?�>���i�� ��<���:�05'�ӏ�÷���|c���-��7R����$kٸC���Þ�4�����=3�Y�tt�=�o�v"����]����b���n��,�w���a�B<n)�beP��A<,nY��#qݖM<���@	|��e�B�
#@̩��$���M��މ&N��x�8���A.p�)'z�Zy�*�-ò���"՗u���	��\g�$ǖ�j'�����8�ގ���䜺�Յ͟;s�'B��7�@���������~�X�\�.l���Gy��s�/z�''�̝�}�u���Gu{�nz)m����'��.��l�D 7�5���t�׼��nk2cj^M:���u�s��r�~]���{X�]�����4�Ԟ��؝���i��i{|��~.k�}���U�dO{��lK����4�ʺz���V��+2�Gk6����wc��_�dx�$=�~�����N���G^�*�<�ғ�ͭm]R�A�7&��{�c���b����S�e柲�/�v<�9�䳛��DL|{|�����}�I��G�͇�\�zwj�>��>��}ڣ�{�����!cόU��t��{������)+Q��{���NQ�d�1[ ��� �����T:o��J��^�{���>/�� y���讈4v����oGQ��"9��f fec��/�s~^�r�e��HR���ԮD�nn��4��]f�c�gJ�M���ʚ�'5�i]N�7�e����]�Z�;�c�r�,o�3M�p�����<}�u�=�8CH��ɷ�dl(�U}�U}U��cn��)�M�B������<N�8��xӰ�]������4/.�1Kp=�`����sg6ܰ�_�l�fɾ`^?Z���`���U�X��y����ۭ{y|)�c�8Fl=q�ј����W����i��ֽNL)ߖ̩��z�Z�Ί�`S|��;&B��|d�r���~��2��o3��S�S~fpm����"`��x�k_e���c:eѫ�=s�&�N�e���6��/��Ǟ��M�ǂ�q��G��Z�4�\��֦
��S�G~�����z����B�`$t��5�Rζ����g�Os�0�]��F\�@�<D�\�e
2�$ʳ�-ۛ�{��s�~P-��?)c�s�3Ǿ�������d���4OD�8G���T�'wOsۏd�^��©^j���2�L�0s�A�(_�9S����*�i�����ǲ�(��=��1��KR���m/��f��^�M[A�����.ǎIJ׆	,NZe���o<ڗ��Z~������i��S�Y�BR��aƒ]�[]�^ ĥn�D�c��i��$̰CU��-�r@�Y�]�JƙԷ��Cɐܾ
�=0Q
KC�<%Zs0�����R�:����X���q�{m���&�h���4ڑ9����蝹_ӹ�yۭ��Yh��H�n���N�>�Ð��Z��t���0ӗl���n�X$a1�7��n�����eҫ+0g�;�1�:8)�u(g�|�CB�ަGj��ޗE⓻mh�ɖ��6����MOP։��;#�ʱ3�k�<+ڢ�3wב�ж�z�y�ǚg`�̑����r�gK}P:�<F/�h��=~��>&�z��+ ݖ�j���.sG�\�t�b�'���v�Za�Xذ.����4'�w�����z�x�D]ES�%����j��g��T�J��8�T� cnË����H��e��nm�υ��E�q���v���R��-֌vM_
�:&y�33�r�O.j��8�4oݥ9We��B�kV��ܠ�m��Yi���׀��O*�)0k�pq���C�w
�1��m�m�Y�%='����6��ژ�P����!kMX�G�5�o'�B#É�T6�����#u�=��و��%�j�I����12���]���5���$G5�2K�CId���1�2�T�G�G*�xXO��L����?	�rh*�^׆�i�?[ ��؈Hlޝ~�AK�t�nЦ���Į�۳+��Õ6��G4�K`��7�ۣ��`M�҅Hv(�5a	Fyp�q��j?��ﾯ��CH�/��35V�����r���	���q�N�g���`-6%�&�:Qz�s,��M�]�꽒$��t��,&��o&�+�k[�5s�Z�F\�k_�3ރrF�O�_��̧��Est���^J���5���^��/}R}R�ֽS/Ńb�%LB�h��ΝܯmMֻg�w�U�S��{Z$��#�k��9M�k�tt��d1������"�t�nH]aZ�I�����:����B%'�ZHP�k��}N�˪��gVjƓ�����+w�����ޢ���{�h�z�J��C9�a4�<�R|��r �P�s��jP���i�G��e�	�V�}7 4lȘ7􆞥�,���ч���l�����/p�w�r��e8���د����Z;�؆r�%��*����d<0��@0<��4�±���w�r]q���d�e�6_P(_�����"�Acs�9�,�^k�h�Wu�7�|̈́�h�RҒע$/U��<�R�Mk?m�ו���|8*����p�]�=�f��C4{���V��X� KXl�N�O�s���i�Τ8]���p���־]u�Mm���,���]էo|Zþ��cMx�S}x�T9d����d�@��v�;��j�u�3+L��@�m��E�	��f��(#�ҥd/$���ͺ'����7o���w��}�$2s�1Ķ��ßL�Z1n�yJ-�+�)iY^l��`��q+$���ܨ:�F􋛳K�iD.z�0.���P���oP;-�Z0�f�,�����WA�6��`�A��6R�мҟ{EB�W�2���QT��Ьd���FF�G��K���ZKf���QI��	̥u��[N��%����,�~L��yzhNɘ���ٮ#�߷�@�E�7/��da����0�Ϫ����!xW[em���u(�s�i��yfH,2�w�3<(k��ǧo������5��"ŕ�E��fX�y�{�'���\� ȸ��xl��W+�R������n#ǠGg�eN�wbyݠhj�W�u2�L��:�)��ּ*K�~�3�]8g��H{`��&�~:��|{z���9���'�bρ�C��F��,��u�l���R�\�O/�{�e_�q�����A�,s򙐿*��衽Gˇs�L7�H_k��X��K����$�Y\��R��t��vtZ:R�3y�a�ȃ�l��:0J�FǇ@H��UҼW��b"v�1-a�u���]O�/�|�ֺQ�ʶo7� ����I+��|)of�p�'S�7U�(g=�)�jo�����&i��i�unt �}�"��苼�tbc���U}�g
��@Y�u�ٻӅWbc3�j6݂E��D]�v�j�W }0�9�i좋1�.����N�J �r��ov���[����a�)�����[�\kP�5���,+�+X�AP��Ϣ̗J�;R�j�f�Z��.�-�
���iw�!�G�6�圆S��=ZeM�ᓲb���Z9�JP:[���֩y��m���Үr�:>&�<�:&��um�4k�|{ ��#�뷢�7�����+���s�^��H�خ��N���m+Q[�n苐�1^U�6 ��"r��M���&闐�tĤ����Q_;�ViP�b�G(�:ef�/�E������eY�gM�ޤQ6�a�~�p�������%nN�dm������9?�����=�p�͛�mZ�������9K1���,�X5!!S���F�t!v(��w�[����'��A�z{�)��6܂�7P�Y`�Y�Ք�NƳ%�l�y����\�YoD�]��4�y�s	��/h�=&vv��#�l<�<؛׍�}�A,u���\�7����N�����ٽ�� �SwPl�f|��3#+����y3H���*��VG��\�I�X�M�wG��U�W|u�	�u`�cH%�8f����,5��S3kd'u���ng%#[��i\w�NX�|,�ݫ�t��.�vf���`�f��� ��=ݻ^&���sm6�)E��hd����2	/X����W:�P(e�Ǣ]ދ%�@fko@̠�ŔZ�����5��FC�	K=�Sq�K(�ţ%C��e<3�!�-w�7u��&'I�Xr�!�����W���B����Y������gY6M<�/{R��f��Ϗ<�����=O'(�(u\}��S_n�a��Š���3�jDR�E-R֑�q{C��rX��b_�w+u��BK��G��T��3R�23��I�T6���ʁkl-.�|]m�w}WK r��fƶJas��f��͜��������dmj�fx�AM���^�W���z������;F:��u�X����)�e:����a�n5ӕsLQ.�7���˨�<.Hpv�n'��NK�c�*��R���wx�Cr�j��VG�2s���3L�HI�^�s"��?��#��Q��u'>�ҟl��_�Ѐ)�ؑ�N�U�B�/���VUJ�[�����J��ҩ;�k��ZП['�i�K4��K��V+��.���*P�3�p!�4zV>D$���V���H�.�=�{�w>"K8 ؜�u��K7��q���KP=��Al뇂|d��ZYZZ�=�=�i�f�R�v�X���J���N�P� ���8���Eʽ5���oj�o[���kC���9 H�~���"	���H�*�j��*��DU�����*� ���c�T�E�(�,��YDQX3���X�"*(#U�EQ�X��QdPU�b�[E����*�E�ʑX��E�������4c���QATb*���b �R��b���DEQH���0��r�
�Y����eTr��Q�2c**�1X��F(���**�-�F1hƕQ�Kl.9��T*[eKF֫4�S�Qf9i��U`�h([W-��DX)im�T�[�DQ��[UPm�����c
̫�r��	mRb,*"�KKs2"�"�B�X��ʕ�QE�s
+R��1,F���[Q[���8�c�2�UE��j��n�{����1�z+�ζ+�D�m�k{��i����moʧj���.rB�ܙ@ݠIz��dd�)5�9��UUWկ��9��K?�6&�)��vf:��׾7ozR%��ȫ��II�X$�t��׽ĺ��ȳ"|U���8�ۺ*_Y��h����u�sz_%��b�M�����m���zYc���rS�t�X�l��Լ�9U��N���N[�<2���"�Ve�7�]fPOP���
�������E�y��S����������X��X4׾��`�ü�*��VE<�J���=�����/K��:q�x�	��0�3b��C�f�JK|d^u����-�$N�v{�ť�=�ژ�w^�ܪ�<w�X�33�w1i�(^��.��^[>*ʇ�U��ć�ݱ��t����r��J�
�7�E��|��R���ܻC�2uU�]�ji�\�ohz=G���I`|bKGJ~`s����D�V	�����Bar��G$���>뻪J�}ݍ��ۃ)A��
��Z+�߯�a��r$pl���ө_RJBh�)�k!v�a�'��g��s�H���)�Ɇ�Z�4��0q-j ���:�*9N\տt�%��L;پ��K����T>@�>�K!UYL��ݝQQ�rdU����
R�k�+yl�=hD
���*�ѡ;sS\�V�\�&HЇ_QL��TO(�O"��L��^�Q^�T���f5�s�V�î�0p3W:�;s4�&�1�dl%磌���ڙ�w�B'��}�����Os�0�]2��%�Q� ��1�cki����y�aZ{��&ܙ��J��~�sxsǨ��B�9�J����Y�=l��&�h�)H�8��gf�V[]$Ik��B�5cV}�er��`�e^ �B��9S����`�s��f�Mۭ�W��7^��E2Z�X!��3ud/�k��g�A��=0?v<s�%+^��-ν��{���0��lw)�yv��$��"���q���=�q=�QY{��&a��o��q�� ����ޗ���n�t��6�e�Ѻ�͞h�˪^U.W:�N)v��ܮ-��PU���od��/�=�T� OU{�޷�	�D[��u���6k��ZVxo�����l��3زt���P|�en.L鏪G^ǈ�^/RϵX�n�p�Wb߇]%xb���g�|���AO�e9����`W����Pm��\�Zs��Y7n�<||q&�k���4㬭�׸Y��7�-�f��J�:��:� ͻ'R�{B�=Y6\/�t1��3�K���}�ϱnS{"��IS��
��R�����&�S��c ;f�̫���&�.����ݒ��H����<����m�`��4�f<Z%�j��i��H���qvl��L���f�:�i4��z�}YƝYE��2�]�)��������V�o�=s� u�
��<Z蕇�ť[�x_
���Ʉ��y�3�x%֍�k�&��Oȸ�N�:2���㚪��>/���H�=)�Қ�i8�߼�H��4�\��w��-'m4G��c�U���Xʆee�B֚�y��m(+��ͻp��i�f�u�x��w"������s�5�9'[��à��|&R=b]���f�6\D�������d}��]�#iA{ق��o�l�3�ل���Qv�ed����G��4M��v�u3w���y
���COX[�A��j�R������ֽ��B2�f�ۙ�7C�L�q���ގ�>ܤzR�$�k~���+/���\:תe��a�F�v��~��[޴����O�+$��M�	of��!��.���{�.OΑ�\[]��_�	�O�N�9��s�_x�ڮ>��4��P��(Gt�5��,�\e��9��EL�:���5����z�ީ��EXN(^}*�&�4��9�TC6;	��EO&�i�������8���f�35� ]�+tѫ�bΨ�x�%�w�l�0�vhy&�Vd~�)V�>e���h�2so{��Ŷ�r��2�(sV�/�Ŗ�R���+'�k���w��E=������^��ڹxx����O�E�T���꯾=ɯ�����_՞���Ι�z`���4w�"`�S�](�5f�7�#�8F+����׷�i����O@�����j��qxK�s�!ƃ�,rO��]�1�%�|���-�h�.=^���}�t�p��iY��T>k �S7���f������/�5�M�/%o+{�X<�D^^ޮ�.[9� �����g�HC�z��
u�S6|i��^2#e�.�7��%;�.k���E���C&ɝ�qn���j+V�qe-"�2<��8/EB�vy'f��d���Kn��w3�T;�d��u^&}�VZ0�l�ŀR�Bԡ�P��z7����1Sی�WW^�EN9���v��f:���K�8�>���쬴x��MC5ʉ]z��˽�Utq%;W*E�+�k�iX��֌/� �o!��; ��陙2a#��Co�<�D���1J^F�+��U30_]����l��jj��W7�ڟ;�5t�6]������3�ߖ�D�4��@��ԋ
���A3,g<�=�K�`S.vփ"���n��`�)�v�N�OA(s	G�i��j�J��&���y+���s�����ꊏ-�v��yݥ��;]G��~�gi[���m�X�`�c��l�c9׵�o��h��B^�ĭ��V8�D��.ݧ�SEh}6l:BB��w�D��7Y\�:|C`��Ҳ�vr��W�������܈����ǁ���x�7Pֳ�
�l�_a�K�/~�L�ηJg��5���Oͯ~����>'�=��o�������ߴZ��������>8t��䮗Eחl��B�3��SX`�{An����^�)��2��"E^G��p�	�L6l�Y�Q9��o�����1�Yo��n���c�zR�3y�nVD��`���:1Cؙva���gR���8o���X�t2�
�����e��Ŝd�ޕI>_/w�����b�2�vg>�a�_f�,z�7�!0�+P0�����ٱ�����u�poK�7�G��%]��`����{�t*��zf,�U9.�c��L>�Uxi�*�9nx�ٵmT���&�v{;a�����;�.�o�wu�'��1,�Au@�-�{�Y�Rƛ�mH{ŉ�ּ�U4d��{�j��g�n[3>u�8ǈ��e��lط�"'ف1���r���w�XdD�cjY����n��w:�n׳�)f:�kǌ=���p��זϊ����b�w*U���/�a�c?��<�{w�v�VK�8\Z8��H�w��OJ��`T<�6���b˓N��^tM�����:�]a�:��iT�uq�ޕ8+Kx�ݩ�ŗ�6���:K�G-u"-i�pP]ݴ#o9T�i`2�M�rO�����-W�E�蝳}�����[�į �W��8���Υ�aY.��<G�N˜7�gx��&k&���a�ͣ��X��������	ę
~I���w�Q���U��/���s��=2WyO��hr@���L��x���|�YK��H��u�(J`J���$W�����=��C�Àl�g�a�֨�4�6֦
��u�Tx���f�k�r�=���Ł��5]Rs8�[���<��(]�)	v�x������;|[�J��G��:��0mA��7�\����qt0��������L�ne���}^�5}[�uw�c�-D�g:С5X�j�χ���gI��������9S1Q�w�ۙ]�Ezׄ�I�kݍQ�� 
�%��Z��\1T�3ï9�2j�TV��Īn���>��?e��W�'y��6�h����p�I/���ʥ墓X�1��=f����D����h���A&��
��7b�Ԑ�S�����#e�F��6xmC�ʥ�u��R�p�$s��6�N�����U ѹ�n":\����?c��[,�ݕ�'�*WZaqf�pɧ��ˬdL��K�P�|J��3�r�B�[če�6��f�i^,�����ו�\���P�q��U{ϱV��'�KỊ�v"�r�b���C������}��������z����wE>�Mht#Dؓ��9!o�ק�lٮ�3�y�������,����&{�g/�[�Ιo�PC���߼lv5X�V��݋~ZF	̶ݭ����_����nq�X�0C�]��%֜e��M����l���i8z��M����[�c��F=�i�W�̪gRȡ�b��u�JK���};�R�{!��&��"qM��W�3ח��q��[���}��}U�q`�ZU�vM�R#�vL$��e��2���Z�X�/V�ܽ��q�F����E�^:WJ.#H��R����i��e^�:���Vx�,�)BLfzT�NU����+�s�O5Q�q��js*��t����ƽ�5eϺ!�U2�*�]f�ʵFR�R�1L���Fd��Q�'[���)��e#�.��a3Pz�2'ʲ�u�K�� H�ܙ���\���XY��ل������;+:Kg0L�x޿)k�1*�Jv�)sg���/#eC	q~z�4��#E�H�!�f�ּ*=��HeN�Z�W���f�q<ZNg�(�t��~�tۨ%P-�.���m���g'��rq�P��7=�fG:�2���"ŀ��Zz9��D���Q��M��p�_F�w�s.�@$�V����i٨�ۓ�{2�_��N}U��iS����-���}�H�J%uLưPP��������S�T�u�
�~/G�m�椔ozv�o˴��n�!Gʘ���A���s�ZI�]軇�{�.O>�{ls�b[��{���Z�)[�TϸJ���$�E�b����B��k���u�^}w��au���ů�~��}��Ԟ��EpR(^}*�&����pJ��Q�a4�1znu����x��[ui�|�{6�.鑙�0R���fD����Q>j�Ns����e�{��Y3{�5=�!v�)����r��w��\��c�,W���13���;^$D#��J��w)�/+H�/�g�X}�3�e�{���C7�oݕ�_H,l�~��C�%�����d���Ll��xv&���m5��u<�?�����^��-̳G�<V�?s���˝wd{>޶�&ɝ�@ź�>֢��R���+�&G��u���bÓ�!5�¨�g����l��a�j�y�Is����3�Yh�m����Km
sapyl#/^B<�:�wp�cs����#f��*��Kv��m����툩V�;u�r� �5͡z褴�h�f+0��*��ӎ1�i��yI4N��a�=>�P��޲8ӈ"�H��e�劂p�/�X8v�Erߐ$�d����,�)��A����W�u���W���
B��ig�T-/c����:�=��N5����G�������C�tӻ�B��t���ژ*���4�ъ{����x��p�y�	�g������^�_d���h�ٯi4l�E�US3>��!]u�V�8��9(��9�..�_i��j�T�s���V�w�vhm���E�+�� ������K�b�s��n�5�41�|ޚ�u�0wog�۩Zc�V$7T�����]u2�33�Ҟ�N:�2�{�΍����#5J�~/¦g��:nK�7�O\Ň�t#Y\�R��x�b�����mV��fU�]5�y�F!c[�����|e[Z|dW�Ԩ}.���l�	mZT�W�^�־�5�J��˯>�����{e&�6<\W|e�9!�t`Pé	c}7Dl�#��J��ŏVXD*���������0�����0RV�2*Ù�r�����w��I�Fs�kg�z��}�l�KϵS�Oτ��n��|%f�����{k��u��y�2Pc��5}�u��z��v�<�6A<y��{|lF�8%�W|�xb.�".���ǆ�(�zӍҘ9��_e-k
r� �H�u�$�+3���"�q�4�o������*���m��K����ݹ��lF�����*����[��T��f��ô(˕�(��U����Y[ý�m�:ݞ�^�I�^���0:]��	z�$l��ҽ�[��6�ʤ{/���[�d��\^w�D�_��n���=k�{6��u���h�����Wg�	{2!�V`LvI��@���3���*�Xj
�^X�*�]�p;��f`ws� �/VM���{�E ���2����u9K�FM5g��Oj�&��(U����<�ϝ��r���YVcB½1ή��Ø+w�MՊ�I�Yd�줰>2�Z=)���z� u5�X҉W���Ѱ����tF�'*X��]@{���(f���!�P:������/�R+GO��@���%;�o-��.?#�/D���O��>��z��;�߾�9�9��ZlK46¢<IԸKb�-u��lm�5~�}�<���L��~{��z��,1�o����y�P�W2��T���ޏ�yצ���番�C]���cw5�3���oN�d��==r���_��������@5s6a'\(uU�#��S�}mgVkrk�C^��G�_���œ����+�ޣH����+n`�[%��C���F�N"v.i�1��,_vK5�ך����;m�B��3+A�>&э��Pkݎ|�'U�nQ�Ӥ�
�,U���]O�^6�w0)�T�������[�5���t-����X��t�R���kהiӳ0n��h�9p�3���O�wkz��t*�k&��dr%��	V5�Zȏt9X폹
��Vѭy-�G�S�O��C������'[�^��ҽ��������0\u��ԑ5��@6+�ޜ�)6�D���vo`��ߖ��AV�mv�}$Y3��l��Xomq�{b�躝Ngu�> %���z��^RP#h#}ݝ��#�kcvaM�R�����w*��ÐCd��D~���|7&�NymH�K��ý���c$F#}S�ۊ޳v�����k�/%E)f�[�YX����XF6Dle��|6�(�$�]\Η�~uw������.�*��e�Z������R��|��[nN����:"�&P0�e�-)�3��=/���[.�H�%θ�ܱ\���6�"w����������2��*}�k��w9�v����S��'[9�䷮(��|�R�1m�!wM�!���x�7�c��-�kuǎ��JuN���`��(�wT�����H	b��@�o~��ޘ���d�I��keK�H꼶4F�:�/jY�טF�}�tl�ԫv-¡�hn�����0�鍺�C&��γӻA�15��"���>�8�򗽓��m��e��gD�\�N��p�,�Yo�硘+n2؊�⻣�zf�&��h�dۘ�q�B�VTkhڽf>�l�Zli7.�n�3��]�`9X���X�}�Z'���ஔY�zi%�	Uy�D����JP��#k)���Ze��^v��A�G&fs4�[�FͲm,�B��p����i���|j��(�Z�+yCVi��`+�|l���N��'�]�ꎴ���h"�1U�ՖS����M��sh��e�X�0nZ��R�h, k��D��P!�E}ڸM9O��+�;�%�i���vF�P��v!�i��s/��Z����1��m�J�1�2� �{Y��é�>AP�����I�z�^E-�4&P�:����ڸR"������֧����B�ũ'<e歜����ݼ�M�S-����TO�r�,|��u�D��l҇4h��.�;i��s�+t1�⾢��U����!�&.�w�>XÛ@��SxK�3����eib$�yn鋋=/Ƭ�[ ��n2�]��)�b���)-�,���-d�w����2��/',�L�'e-��%�6�SQ��*���.�����Q�c�*�K}�Y�	kJQ��J��n��l�h]���<{�V�z���I��I��X���h���[DQ�a\L�(�*�[E��f)�Z�ZZ�
�mQE��X�Z�Z�30�Kj�ˈ���0Z�EV*2�"�"�*�,)��b�TUE�J��D3ŉ[�\�V"��Qm+��8ج�DTX�D[EC-b��5ڊ��DT�"+�J5"��UV#,*�c*J���Uư��«U1�V�UY2�3�c���qF)�TZ�q��d�+���#b0�ʂȰ[[Z�r�. ��h"��Q�dphb�m��Y��a�ɖ�J����*lD+Q���TE��
.[�X�l�#YZ�Ƴpq�Q�Q�b2�b��lYiCQV+l�"�6�r�V�&VɖR��1�em��C-�iH��� AI=���O����6�V������7��٦k�H�/���'^ �qY�2V]��1��N���ƶsl�BP��M�q�ﾪ�����trQ\�D� h�P"�Y�P|��3I�_���A�B���*b�zS�5r`LUz���'�����j�VK�9t:�F�%����5�s�^��ϱ6��{��;��
�C�Z��;����cv',�eC`L��D�Ģ�+�o��'��3<�N����1�8�=����|��2$F�J^V��<�E���/*�5�
l+�+�T�wY�xڷ��t ;��������já&Ĕ�|����u�͚鴰y���~�T2G.�p�>�+��鞤5��7�F=���[���z�8��R��v<ű�7\ٮ���^Չqv�!�ۘ�ܮ�ǆ卋�M���ɻl�Z����\��'���۹g{~j$4�(��"�T:����wp�θ�6�8�;��b�=�0C����Ll�6<�Mt�����f�r���S�*��7�H���z����vH�n�J+~�B!qjާY�(�~~�]F���8��S"��d��L�I�v�+���ݢ�s=/��Э}R�Ϳe8����#8��Xz����R�j��ݼ�M-]�z*��v��a���-6+�攅�o���Q�m�V�&��]�m]<��s��v�2nnr�\���^Jg���e�ta]�1�#p�����ROޯe���?���K����;�U&���3�x2��B��+՗��_wk���dq���&:�o�0\ZW�*��v#/%�hd�o��AM�)�v�AY�S��nq��_\�@���bL�&�<������r�J𻭮���o��^�ˍA�}[�9�+�t�m�q�>;E>��Ѳ�5�i��t9t���J�L����yj�#<y����{z.^�<a�t����0|���ʽ���%U3��^�c�.=6��K�Z!���;&�޲�G��玼�9q�,�S��*b��A���C�"�MB�E�=~���^wJ��d�:#���{T;5�2�~2���G�ȡ����,�:<�y��aQ�%�w�痒�yf�f��o+=��2(_*�'>�.�'�ֹ!\5�k�ծ=�g���WvC���V�9պ���P>��ˠ>�+�CF��0nCOR���ڵs1
q����T����,��f���/}���(j\Ab��9��o��D]Nq���n�j�Sh��b��I�w���t��� �~}��x A�U���_n�\��~�:%�X�ĳ/V�5@7F�#X�@��p3��[�Z���I��ʖ���H���Ԛ�z��`�ˈ�{Y�ݠ�{2���-�s�W���+E���[3�g�݀`ǋFP��D�:|W�/ ��S=�갽���^��� @󒷈|�޶�kZ�<�ws�jԃ���]],2�[61i���Lxy�]�5.�&zs����F|�÷.��J���ɝ��vF�8��\Z-� �j}w�Y�>����,�W
�j�V�`C��N��J�0I.wV穝ϫ-m�Qs�ڜ�ʢ�C���.e��9X����h�g=iifs������j�V2u��;�n��83Wy��Dh��V7>���R��]ACo弢W�F)�mY����y�G���t2�볇��3�m�0C�W��6
�"�UBX��!-��9��:�C޿)f�1)q���w,�ڽ��(d��"ĳCmݣ[ԋ�+���ќ�	h;B�:؟�R\ń<��󸋇}Unc��y�����X"j�$7T���rP��e�L�w^'�I�o�wJ���K����)�J���3�G*ύ�w����6�:��{���;YK855���۝ۧ�Z�{��d��g�X0{M���g�5`�O؏���^`��|����32.t����`�x��$��:�� ��GV4�/C���x��(���k
w.5�f�?�Sw�Ix�xǶ�k�������,o޼�&����r��n�8=)r5��)�; .�Z|dW���.ɖHg��x�p�[ެ������H��K
�I��T,�)5��=�r� �e�9!�w��瞃�D�}��p׆{ɝ;;.��D��F�������^�՛�H���K8��^����zlSo�{���$נ���s-�t&i���k�GK�K�j�gßC��Ǭ���;��HYQ�(%.��n������;�ia^�E�r��et�j���C<���.J�w�z	��u^�^����h�u2���ڄ�bO_i^���{����_����b�5����C��5#������;k�}�ۆv^��:�Μ�x��3����vnQf^���`��ֳc�n��.U�v+�y^X�^��ǎ�6����Z|��*�ډ��1/3��ţ�5�/�^���	���3�/ �*O)WPs��9��˅���f����C`���2��S{��q�c��Y�C}J'��M�����,����&��!���Y���]��s�ˤ1T��l"�%y;|�N��ySǔ���©��;�%^��h�ռý4]��J�=6-��:�SI���w^Y���WL��.|a�%��u|���� p��qf@��d�fb��^`�KA�񊒷�so���Q��|*�{7�������:�-����rρ�C��T�P�P�W���4^2�t]���{#����4�f_�Ki�z����;�ߥk|6
�(���Q4�|qY�5�b�ə:�o��p��5��**J�FeB2}�`ɵ�Ys���.�	��:�x�n���'�����=�<	L]�P��c�ś����z��N�u��4~��G��x��z�n�t�s|���)��6f�k�"I@�=���^lV|=L�%�7�B��\s��ӧ�����/r�Y�F�?z65��羗C��hC%��lzS\L/��5��Pf��ړ&Df�6S�-y���cǚT�l�',*i%�"����I�t�c7�����V	�zEe��GS�嫏wU%�r�"D`;%/+yv}޴Y�e���z�=l:�%�5r������Pz�S-U�þ37�o�V�6$�I艿<�zא}�ܛS��.�,����1XjVX���Ȇ{h\\7+q2ό���4m�x���N�|��o�f;�WɃ��$�^�ڭ��jyE*Η쀵��Z�ztc̭d�L2�G�ޮ~�Й��v��+��Է&C�&�7������!̃z^��N�i ՌS�wH��;�	�u�t!�&�e 溰0����m��y����O��%lU�6��~�諭\���3۽*��oZW�����ۘ�ܮ�ǀܱ�g�E�즖_l̒Ɣ�M�Q���]%�Ջ�OUk[ۦk(zet�*�e�װ��\�;P�θ�1݇�n���{�����T�'φ@��g�C�\3hx���U��
u�X�dо"=|bӘ2-�)�V����>I����r�@�?&2&j�WJ-#H�V/Z���[��uڽ8�W���o�_�MH���X&��'X��I��2���2���V�kƃ8>Tk�#W�W�6���Ȫ��!á�u[,Źq����5�V7��-�̛v
�O�U��{�J\��X����#yX�0V
��Յ��M:蘭���r��iM�@�L߻�t�]�k����F��Ϲ҈�!����d���(�\k��v����*.�+O��S}��v]
cC��fU�sr%uLưP_!^�c�.=6��������y�{&���ڥv_�Pߖ	*bp}2�,��Z49�-+�P��wx��R�$�l�ٍ�N]�癖to��v�v4Ժ�u�D��pb]yԵ����ep��8�=vQ�:}��q���j��u�*O|��|�8:����z��B��<������+�ѫ�z�[j���=�޷tkX�����(&�I�h7���mwt��t�t9��q����,��7=.�m�����{� []T˅��.��J|�P��(Kyi!_k5ǜ�rsm���}�����w>��Cf��G���FZ�B�V�8$4��Ƒ����xl�Z�sO��|��'�'ʴ���1���}�͗@|��nuM�hّ0d)�,��ϳ�����zt=�j~,!J�ם�ֺS^�U\L��Kȵ��<�J|�;}�q��:2�g��'��������}vl��p�f�	YɊ��^����w���}+h+\5������r��+�|ۮ��iM^kO	����� ���
Xe�|�����M�o��:�4`ܾ-��,K]���q�0M�;��[��eG���%�b�5GG]M���2��H�.�ձZx��"X7-����=�C��\��=L�Fx����|3��������R��ZP�0V�p��e�+K1�NP�(g��ux�5$����i�[d{�)\�Uh�v�8�Te�T4��(m���Jǝ��Fg�5��ç��h%���=&���n�c�E��TM��|�����\��F�����ewQ���n���mW����Q<��77S�����ڳ�ܹ;�,�Q���g�Z�Z��%��$ܹ����nr��;u�k�5�tb�M���9r��7q݌��n&�����ޒ����y�����Ɲ
��#�:�t~�$��eRǺ��{<�<#�t)T�0��|��3��AC��K46�wh�$X�\\Y�̼�V{o���oד�͓�7��v!�/�k~.&ld�7r��\"j�h
�\٠���ή���Y:�{:�5��o��ٷԦz\#Z�X{>�3�G*Ϗ�3��	�(�:�s�y�+=�W�^��-6�jR��쪇�:�(s�=)r�؏�L���u��dW�Ԩ|�ߍ��ӞN��szJ�O�	$�i2����}v+�uȽ��Y�c�E�q�.�}��:o��}K�	�a{��2�th����	�
���GE��OˇQ��\O}}*���ϛ~����o��T��`���5�����w�^RV�*at)���U.�,t���~d��m��T��r�nɰ�nX�nJ�,)�Qd\�}���U�ji��1�uv&XԔ�b�� W��Ǻtf޹�=�4��`=�I���Ҽ[��6����c���ə�wS�y�uWqWF�i�^\G;7�����F�%tO�՗�:me[�7܌lνn5ئ231�ًr��M����q+�8nR�U�Yӥ��;n軽$(cl�t-N��j������RA�s� ,3�pg.fp&<��]��UW�������޹e�U��T/K�h�|%\�����Lu�8�<G&��������6c�@Ƕ��Ӭ�k�7F̜j��U�KVXdU��p�b��l�ws�a~Wgf��G|�L+�5�ͧ�&�wr������j�Ϫ���*�&��(/�R���b|y}�7mw�����������;T�V��q�W����N�����$�yyoW������ѯ5p1����Ե@\���{`uze���CO����2TjZ?:l��RI�^�س/�mx�e�'y��9�;��f��G�|�������:��egz��\��T̰2\�E9S˂��G��`��|՟=�<p���"�^�H�V�n7��-��@@Y}�R)�P���X��7S˂��,��7\�4j�=���.�ML��"юWk����W���Y0��4MD��{o�(tY�P|��3I�_���;�bw�����؊���豪/=Rl��o-�˞���9�`��Jk����x�M��Y�<�!3.�1S�qJ˯5��w��}@��7>j�kr۫��+��b�c]!�y�yN8lT�>GU �esM�v�eoS>�76o��:��� ]�E���:�㽒#��8�Ѐ��y*osn5�jN��ne�s�ݛ�+���J~��ּ痟�J�g���Ƀ��wc�>������L��$��#����?���9ܝk/c�v�mꦶ�Ma��t��6�`䔈�7%/'uA������S'�B`}���	ft���mxu��j�ޡ㺤X7��V�ՇB4M�L��n�	m{�
�.gz�:�w�N�J��X����s�r��x��m�u<�\�����Ծ=b���Ǣ�ۮ�ّgޫv�D��m�%xd��y�Oƺ�@T�Hk(��R����n����f���"��c�̦���{����(L�M
�--{	��v#��ի������kiV�Bڃ�s�s\=~^gf*�E����&x��u���u���k��.�sc&�8e4f�I�<陁ܼ��oW�2&s��c�Q�+--g�ޞ���NK��3�ޚ�z��خi�y��,o��;��T�\w��o,*
�j
�x��zr��A����EC�/�T�{�����0����y,kC�o��AM���j���j;����h�hR�v�=�Uv��.��ʳc�1�6�"�
��W��!��).�)�N�� �I����p�s6�R���-6�n#������6���(���u��w%�u��6��L�
��άU��-V�Ps��m��Y�Չ��̳�*�_:��L�W}ʂ��� Pu����F"/�w��R���TwJ�D�J�7+;dflj��cS:�Suj�Q�;x�]Nm��
���	f�n]��wD5y�n��j�<�Vu�?g�f���Z�3s�+b��o
L���j�:d=(��Z���Ҿܛt�.���r�v�)t�Ά�q��-�7>bB�ɚ� ޞ�Fp��C���u-��v���iǑ�7�R�hT�C��#l�Oj�Qf�f唈�qލ+�d��%��j�P<\���f�}y�ԅ=�}����cenX���V�3���Y"�1��U9�*͊B�i�ͣ����)\$�WbWh�Vt�
�a�z�ehu�m���7����	��g3u�L�1fwU��B���.$�U��Uc�VowZ�zY�ӵ!����셥PK�|���l��;���NF�@�g��7�'�"�("g%�B���k,tA�H�L4�y$�r��u$��|Z��
�T���0$�Qb�W0�S��:e�<j�A+�AN����냻�
�a�!��en��M+uھ7(k-hr�k4���tVG���.�|����lT덠�<�� �ˡVPqS�M��Cmw���)�&=�f
�R���*uk֜���X�����ZL�������!�Z����t3�}!���R��M�&�D�:�h�����ɖN����7���~��u���oN�Q7��p�JAfoq���`�ymĶ�-��rc�����l�oR���
�e4��W8��y��k�\f��7fV��� ��`N�D,�.�)��F�e���w�r�ob<\�Ѧ:���+AgǏm���ۘ_r�U�"jJ�E���wz4J�B=<�KQ��}v*t�4��8Ǣ]�l=�v�Z���ml��|�������m*4���*�\�w�	w1i���k��.t��Gy���5!/-�bL����7���:�J�ő`ou�\:beinnu�O���뇓� �+	�Z����p��.�T��VĘb
�����U�=���vq� ��۵�Gv���e�6ܵ[����(���|����q��-���ò�.�3$�>s�7��q��Y!a�;���+�E�#&l|�s�0�\�v]ɓU���,Ba� �}�78@y´Z�!4�ʕ���Ϟv6a��2�!%B�V��|PxR�����w�N�d\r�pt�s|%��p���W�C;K�W_!Z�4^�AH�*�gG�&�FJ�G�srWs���Nr1�qrQ�؍Ayf�!Xr]���^{���N�ֵ�t��2�3I+��1����Pm(�X���aX�bd\A�[ef[�P�Rc!X��PV2`�*�2T�*bb[b���\jZ��X*���#��P��j"���b
j-E�U1(��+�eH��X(�LqP�LTTH��j�j���X�
a�QJ�dU�$���+P�6���3,�V[k��c
��H�6��UB��B���1�p`VVB�1k
2cdɕb�LV��J��kKAe���@��q�U�R��\�f[��fJșk"ʗUCi�c��br�R[��2�J��q�s3IPq1�k�VbUk1+d�E��q��@���آ�X���X,aPīi��0E����[ejUb�2��j,���LC-*UH�1r�b���*��w�z/��]p��y��ZvRK�{���I0%�Z���r�v�-�j��㏶8�q���Z.Vᕜ�M8������Fndj\����w������������W{3`���XY��d���Qu@�+�w��9[�%�����&�੖��Y�y��(CH!��/m����q��%����yh��D�i�X��Y^����5��p��S!�s�*Û�d��IdǅVCf\R��6�]��Yג4���쭂��֔�á�o��1
�z���s��27�M��xsiR�cg�U�D�{�9	��Ջ̵1�ƺ,2�~2��҅bJ�\�B_�-$��|�����c4^�5x�˸k6�Pg��O+�����ʶ��͡�ܽGO[�'���/U^soXnd��46�Wy_ԧ-Ϫ�B�?nz-�L�ޖ)s܆��dL�N�̏ӹ�O����F�U�Pwv#ذ�9BX�2ץS\/��K�~;�r�jgy֓�+��=���ۗ�Du��O;��K�+} ���| ���D�=
�~2���c=�����$c�{�o�7�]���3���s���ٍ,kZ��֛��ÃV���z��,3��~!�S
�9��A�����)���M�Kr�FQ�a+D��m�w�0%��pz�g��Jtq^z�G�$�:�����P�L�@u8X=�aO���9�[0pݥYov*�s�)��pTjj��<��R�tP���)0����꯫�خ�{��g �~�H��/c�>��ΗC&ɝ�qn�)Ec��\^ff[#}���q�}{����Hh�)`��\`8<���}�l��aΔ;�g�K�չ�g|!�=����M�ʒ�>�4x�
^�,�5 �+D�}�2ӭ,�ws�>u,{P��ޒU��Yz����W�;�~��e(����z|�t�E�LP�[�%~tb���F�ޜw�T��;׏xқ��k�.���Н�f�Z�X:=�U�K]RǺ��Mv,��\:�3��)��W�Gr�|a�Y�H,2,K45�#�ԋW
��[�����'�^�/w��<�<��=hA�6�62s��Kg)B:��������B��/'wr��i-kt���C/%�SҡiԬ<��"9V|`�38߾��6l��2ꗐ��T�+��͂�*Ҕ�\�=}R�0zR�,kv#�S0vQ�>2+�E��NfV��>ݚf�Mx��!�HCΖ�R���a��uH��Mf�r� �ɕ�]Hi�󼕤��Y��U�83W_O��<�cM���v�sz�SN��Պ,q�F�D�G.]�b�Y6�,�+x���E�K����)0eo'�o��
+	}yv]z�ew�x�٫;��#˱k�� \��.���&ۉ�������޲�7��G{/*|xxg�C���!P�T���S�����I��i�W�.X�Zy���ӣ�)(7jW�1��Rkp	-72�����L.�1��[��Qio�zV�k+��V�N�֙��d���hr�r*�»Qd3\�}����U�*r��אognM��o?X�
�����tw��#��4�}0�jE�'���5��sl5�ʰ�Q6f�x�e򓞛�}���|�����B����s���<�}}j�^�,ym��0oR�s�/�DJ�=�>K�t��ˎ�RyM�	CFx���K��}r��0Քنf��|�]�q���
˧@�^�a�[j%	5�9��ѵ�L��r�����7]NǣJT��Œk�z��;f��(�^4�
��2�7�]燅�����>��g:$��Q3�Ǵ��'P��r�킆j��u@ꠗ����/�5y뗱���[����4�8�ᲄ��6���w��J��`�7U�c��V��x	7��5��ΏY�G��>�����u�K�|ͥ�8ਊ�"��:��N��"B�4WY�j��(��6�l�����f���M�p�v���"t�:����s����X�7�"��-�@�x�2Q�3ym�x�Q�r��
��&�����ѽ{����I�<���:�*9N\����=�L�o����y�
iW�o8�1w��&���F�Ў K�yB�K�,qf�7sW���q{B�|�5�~��H�e5w[�)�9�{m𒫭���i +�J�+6+>�x�&y��t��i�h�z��	z<�mlYK��������|;�NO
���H�JM+���K�>���!e�����R�\^�,�ǉeKv�N��v<s拉k��',*i%��"�������i�ְ�Ob���ۜ�m�v'�K���.�f_.�9%"<�%/+yvw�$΂�ƛ"�Ul�_��Oz�FY0��V:�T�k���fo�
�L&�ЍbCL�`t�}OڮP���V�����"})!�2��j9w���"3�c�ܭ�<�\U��{�v���,ܹ�}K_��Un�)|x�;͞Wۥ`�,�Q���K?!�d�Hu/gU��ɤ���W��)>e;�[�Z�ʥ�w̚��z�z��%�+�S:�E��� 6�Դ6]'B�JqUN�os G��]U����J�vb�:o�ܜ)�6�9&J�e�����5���^ޮ�қ�uՕQtx�g�d�~y�[��JrA��b��z����b<��*�v�fc9�̒�����-��׈;ø�ٻ��ĩܐ/%&r��FwC��*�p�ӥ�M���G��q�����.m5A��L!l�*~�~\���IͿ;½;�w���0;������Nm�3�x'���x��xg���+-Edq�.V!I���VN��s�%�ݪ��-����|)Ďy��,�m�-���5Rmq���*pxѠz�hɏt�a����\��CC��ԥҡ�/r�Z[���fδe���՞}#������}yx�]1�ӊ�<��#,u�<N��\C����f
��,��7�0��ODstV�G�s7��;W��gݕ'��
e��G���χ:Qq��qv޺>�2j�9�[p�N�=uY8��Oˏj��-A=P���fş �i�I�s��T�i��p�u�UQ�^}����T: �c�~�p�^��_��Y��d��Q�&Tœ���5�:E�Ol��Qק�S|�Z�x�˶]��\�y�="meL�_�2������P��(G�m�k��e�Q�����3w@n�Ӫ���Sξͬ����yY������(X��&B��\�ZjJgX��f��t�-�uY�=�)j����+��n������w��O{0ʉlF)V�bjW�"�WaQ¡8��Ob�P�*�^�i�$�{ja��f�Q:nV��et�W|�8G�{uܛ�%(kYa��f��w.r�^��[bG8vtF�	�X3ڐ� 
���[e�=�o�4�g��t���'��s��\���r4��׼�q��s�}�+4Y�Gw��=k#\/�����~��u��sJܐ����ݝ����ͱb�y�`ᘙ����ѹ��f���MU�zӿb�6^�����zzn�s��*�S�q����|���-J6���ۇ�J����B�<>)�ەm�Z���Z��w�zdGݗ�9TG���P�6L�Zd6���	���T7�wq��5�X�����qT.�+¬�|t���rَ������	���7��j���S�3��>�ݹ�&]�-�ف>3�q�C��`�Z%�s�)��V�e���(}$y�׫K�2y�Ӹl���W�9[?_���Yh�:T1/R���p��3�+S����yh�a��V�5��g@��h�5lL����Jzf3�>�5���Mq�eUq�/��^�y������k�2kݷL���o�}J+��%�y���XdJ(o���k�,�.+��s��5[dSb�蝣�V6ooDt�WԻռ��"fܛ�4u������'/��[�r�T�kW��t�����T�T��&���9�:�e홂q��I�{l���iGw9՞Z�]��7�Y �;�i�[|T��n	�H�]�zj}���YN��]9���׆�V��\Ж�"D�.�3�j��ח�*�|g_o)�ZZJ�yB���:�)��֕�;��!�#�:|2L�72���N�=+��癭���e>�EA����}K��)��딡��K���؏�fx�jZ�nJ�-��1{���Y�Vj2����&�#Z\V
N.�a��r�)5�:La>������$���y�U�Q�Vt`P��ѱ�:�!P�[�xg��V`a���ߎ�z�߻��z�i��
JÕ�.�;%&�d����w|�yL����������ȝ�s[�툽�|��im.�c�ng)[Z�ӫ�Kņ긋*���":�Cӳ���+������E�3U}�篼�߻�x��<c�d�{p�.O[Ҽ9n�B�ʭ�/�Wy�I�O]���-kԽ�0T���[Vx��U�e��l�Ǳ�'�\�7�#��Z�y�Ӷ77(��n՘���,r��/��qؠ��y{�n��YD�f��$�|�4��X�(�x�D��Fd�5�<jNy��.�U��q�̖���\ė��
oki�Mڰ��Y�ч�-���=}�m<�Mn��{]��vY�Mqt���#�.p���h�Et}���*ļ�kF��a��$��	ۗ;��M���RN){�aw�a�4�Փe�6���xT9⨷U��U�y���to4����T��m�x|�M��V��|T��F{��D�Vn��<��m`U����O%��go#w� <�. M o�iE`��&-���,kXm��T���k
K�������%ϻ��U�`�3'R$}�H��;�߄��a��Wr�0��,d�a��q���˥7K�#�I����o'��qx/�⣂����z��&#c&�5g�y����q�h�%Vt��2��ީ�H��n�"�����
9�X�L���Fe�	��h�B��0���I)��w���zɆ��h���"M8������춳֕׼�\��k��E
�:Q~]y�;�п,Tŷ鱗9<*"����Z툏;k�f�
0������k6�Z���Mf��E��LJ��~���	(M\�PؙI*�"�������zG��w�޴o��){�C���5�zU%����l��x�n��uԶd��5b}*gY������U�<��-���m���eC��+&AWD�Ƭ5Vqh�W��ڊ`x3{����p���.�KۿK��Z�{$��k�V������:�m�J�˶ݎ��M��(���w�P��0.�y��Q�,EP&�9!Gm��U��ȒǾ�7d�w\����.C�LY�.�},��B4M�i�k�䣼�F�x;�gfZ@_���l��f�{h�=�,{}W��kֽj4����h����m>����	9~xn,�Np�ݺ�-��J�ȗ��sƜ��3���L]iN�A�fU����`����C�����7m��4顫�3cޥʭ՘*�Ԭ�
�<�����&�����uV�gݔ�c>۰��s0o��B=��Ϙ\�j���I�-���N����|��Q�*{�0����S:ɡ��\��;�	8�31ܼ�5-��Y�mZ;=��z�l䞶��ԋհ�#)@)e��2�����N$s�T�`�p�����5Rmq��o)XU��>��ו�9u4��`���M���Bk��
7�����*�����cZ��w3H��p&���6�V�(بԴ�l�G�Ҡ>K�d��{�٘++�4�j����^�x�E��$�L^N����+oeN�zAL�e����h��J#`�0�G෮���Ϊ�K�im���[ϱQ��eT�L��ZP>���艸�_W^�p�@�#�@��+z>���4"�� ��Zf|x��m*�(oe%��y�v�$�|�N�wKe���K��[��H�m��6˽�H��2$٫�Q#b7�c��s+*�枮3Pc'<��	�e����c�x��׳Q�	k��\�.T�w�:�Ve䓙��sH{ʄ���M����~8Ӌ5xd��Q�����Z���iz*�7���qda>�r��/ϯl.SΑ��D�R�%W?�	kA�r�w����xN�Ǧ=)��r�AU_Ŀ�M�*���}��R�Z2�/��m��ٳg����q�����GP��Uͼ&��»��>[x.�Bǟ�=�Fg��$ �G�Hu����n�i߯����v���z�t�v�pzD5αZ�Mp�2���]�_��뻱5�#�IY�D�W�I��~�~s8f&ugL'M�͸p�f��Yg³}ed���-fr���Ro��Ym�g]��;�ؠ>��qAc^�i9��r^mi�ڇujA�� �Ey����d��G{��Ხ=���x��zf.��n2�M�;��y{ϭ�'����zZ���j �%me."�2<�]ȯ8U���n[3��w�t��'S_����|˗N��4�2��.����1fi��z�N��Gf�Y��Z�1V��L�Ռc߅.����N���vc�m�z5�G�I��R�M�F�Y��M���ד1�����������pO�g
`v&擗�u�V���-�������jv���]��	�=�nm�����YY������p>���bEe���ܒ��w��wJ�Vth���v�5�R��+���2�Y�tV���X�*=���sI��@�㨠;8^�QK�7��R�=�����!��<����3N�z\u,^2��[uݰ�Kn7j��2���Xp��b�]��:bv��u\�����w7y1�,�v��J:{�L�9��x�W����!�XhW���b��j��P���~�Y�5�*Qk-Bl�̭�V���[�8�&i�r������k#�p]��Z���;nt���<�*�����:�hn.�$�WD՛{�X�]�(�Y���-��W�v.X������:�n�N����d�y��V�cH
��4�QM�:��e+��%L�)�WC�w�c�r��*��M\�eQSz���j��:{�+��:&�0�5*w�� ����t���r�|X���q�rƅ�`s���y��W�G]��^O�����>(�o*gv-|�+{�n��޴k��J�����Lo�ݮ�:U -�ӌz�P+K��L1��匭6�{*qW6�!+o�a��QkMF�U���Z���ԟ���w�L�MS2�x�n��䅆6C�`��2��̻bl{%Zj�ε�'}y]q%:��"K��y�)!5�}Ζ��
h��7�\��㺦&le�9o�vU�p5�5��a���m^�!��̀&a�R�P���s�&�DI�9PB�vU�O3��r����D�;Vu�WG�3 ���d��]�����K�+2QS47���O�h!a�\K׽EN�\uu��$��Z�u`�"�����Юe��M���h���M�fF�p����L��Cj�;�o��K\�D�O�v��S�ȡ�F�n�)wN]Mo�Tp�1ᴘp�"��[�{RnAK(��"wr��{���IH�%��6v�����qi��l�G�'k��(�s��DZ��y�b�O-�4A���V�h���V���m�$U�b(�2�CY�ZL����7k�v�V�h��:����h&F�!T���nu�������s�k3�V�a&0cxOaw@	Ϲ�#��P�lي���^j&Vtv(rRG�'�=l��)JeF��*�l��KH��5�t�`4���M9�Æ��J�&�oJ�$M"U�����ɴs+��5��e�w"�a���wl>��-e���+��R¼93X�L��.iO-S�Dm����C���\p5������;���p,��*PEc*U�!���G4dx�"'�aw]>%Q�$Mř�É��z�}u�tY���*�AqYU*� cd�L@��1��1& ,+,���c*�IPE�VJʒV�JLeaS�mJ2E����AIY�+E�m�,�,Pm�bC
Z��P�UVe�QD�d�!X`���Ē�h��r��J��%b�T[�\��+��[��R�2�-E
�"ƴ�[�TZ°���Y+d��+"�ʆe���[J��VJ�d��b�"�c@̰�+
��Ԩ,���S-F�����1
�q*b`����e��.e�al�`(9`5�[�U�.[��%C2��1�pF�C2�U	SVc\�V�#��'﨏�A
�Q��n�5m�J��p\kMպ���{�"����^g�(P�!�N�%��c�;���+3��r�^^���rG3(�l�1�L9��O���х�U��@�9z�/�D��&Zb��5zD���g��ǽ=��Ǘo�M�Ea��+g�Kb�Ge���{Ϫ��υ*Ba���o׋{2��d��~<��^"�3�<�o!��;�g����崚6
�"�U\b�a�㽫��	��5D)�\Ұ�55{�:�W��K^0�Y�l����k�~e�r�ܯ�D�5ǭAA3/�0�S���Ynmh2&rs�7�z��b�:\"$I���괫Օo�y�W7h�K�ڕA3/�Ҙ��I�a�Nf�����d��o-����v�W��W�C��Y��8��!��WK��L���r�8=)r���L�����җvs�ӧr��w�Wj�����FA�(������q��.����a^ܘ;�=���.���)���}/:��(��ȇx����HjΌ
v�˳�H�GZE��]{L�K=�dǵ��w�r�z��g`޴�`ޘ)+r�a��II������wıND�e��6��bӷLSC/v�eC�C��\t�7�cD^^+k���Q�ҋHKk���q��ky��}o*SMGJ��K����u~e����+�YO�ڜ[N�MLjc��5L�&,�	�0-��_p�[��7�� �� A/�j� ���=��]��JQ��9�v�K���֪�|&o�%���V��+�j^����p��od��g���;Q��x������=�X]C<���y�L�ý׍u2�L&�=�I'�Ey��5sE��>l�Oʠ�4�"���cí1���+�Y��
Ƿ��$n��Ъ2}]������i����Ndȇ	Y�1ҩ+�y�Q�
_=���3�ԫU�5}��c*F��6@��as���,�'6\#|.;:ᗁ1�,g�/%�R�k$tW5��<:?w2k��������.��̇�RޯE����%՛��m+]),��B���$M�s/}�3n����ɡlWo:���iE`�� r�����k���uN�7ٓ�_�Zƻ�:��[j
�fe*�e��5��D�}�P�SR3�N�7�C�ð.�w�{�8�����W�ٯ���*#%`��lO)W���Q�r�=p�xl����o��WC]ź�����.@��_y�_�U�N@��N�;���!��sS>�C���9��s�>�W���+gj[��Y����l��G���6������\y�|L�^3ˬ���S�y���V�Բ�q##"��W���f�	̤=j�0ߣ�`(�s-nc�ڃ�֍�"�e�E�˴��G�ˑ�	�Agh�QZ>�V��}�jL<X�����j6{WܛqX�ԥu��'�����`{�L70�5Α&�_��ټ�;CK�����jzz�&[}�?g��A�/�$��o�Od8p	�P��H��I���Z����罅;Q;���WҐU~W��v��A��*d���8$�k�$�9K
�I&�2D¦���޶��j;�}[ZE]m�`�-�{�����z]$�0�*�$�G��,E�+���׵��&����A޴��^4��]pT�k�P�>�}��}��&�4����Ob�=P�t�Qc���G�uo"u��ٳ^�K,�?:���:u	���y����/�#�����'��W�~�h���g�[�K$z�B�o0��.�V�:��W�0V{E����ۂ�����n��O��i���:�k��k{ue�5R8�d�ɔ��2 ����=�.�7_��a������ە�1�vX�f��Dұ=.�m��b�n�~S��r�6!~>���Z��c�WG��t��r�O��^��"�W����V6uM;V�Zk��l@is�$��r���tߎ�7�Jw#��nuT.�zb��ՅѬ0�y|�F٠α._��^���v{�9�w�OG�U��\��h@RK:n�n��&{�|sq�fK���J�C�W]9{|�noGc':��*a6��7�d�9w#��Q�P�
ZZ6�JZ�����8��1R%�M�E�S�O5Rmq���r/);��C/xt4�L+l5����e�B��A�����CeT��y'�*_��e���K�0mS	��"8]p�~].r����H��v��@I�$F�uO=%)�ޜL~�r�h��Xp�$2V>/ǋ�'a"�����<�ޯ	2��<tK4O4�>��0��8��D��'��;���~��D�h�9��=k���˘; ��6��:Q.K٦ϵ����i-}GmJ
Vڰ�2���p�J]aߚqf�d�������Q��Iy��:�����d�es|���G�]J���{�Ar}����a�6��\/�]��	K��7�q�ûf�ݮ90��~�'�PCk�i!��&�r��)�S�\.���ך��>��!���5�'{�<�j�TڇnU�P�+��R|���D/�ݞ��se��^2�.���Ӄ����B�qό���=KK'MY�Gz���<%���-���^]~��M1H^�I2�|iJ2��C�=�f�V��ї�&����Z�q���Q��@���f9}���us�zB�Aε��g-
�Э�T��^��cg|��y�=����	�	���)�H��K�L�n�/v* ��dMF��IɃO?W�(�<C���>��p���f&t�-���T��䠿fe���̾�����p}�CU�����]���?o`>���{1��kZ��ZosnsLI�2�5��yf��T�g���V�%�ˆ�Ŧ�8=��D|e�U�w��/x7���:X#-oB�#�Y�sP��,#	dc�C�D.�q�;�K�1�l����;�������y��%�³;='mN5����E��FG�Ҫ$}Hjt9 �Z%�s�)����[W΃��l�Uy�1Ա�S���-�24?���3�H��G�����#���ss�5��Y����h�>jr�����Bl���VW-����7�k�</�-�=����Y��6(�/�X9�9(���%�y�϶)טU��ô�u
=OU��Ş���ꂞ�GD��|�P\]��k;�gβ���"g';�}=|ױz �j/D����k���κY��˽Q:���Z^P�e�[�0K�k^=~<��2:�p��>�rX�)���RL0�mR����F����e�t�+Xwv&�� �[NgaS�[�ݐ��
���]XH$�P�lAC��u�5wG�ޭ�4`ÓG[W���H1%�V̚�V��+�P!�>ǀE�G=�זs&ZBݍ4�m�s^�+�~nK���9�^�ܽ7�w���t!f�WK��L�uJP�ޔ�݈�F����w���~:�N�-����.ɖK6�F������.��c���Ok3ԟ
YJ����o`�.�?{yO�2���՝��neه�h�;�ge�7]}�����F���5a��5��0RW��s1��RkF}%���ѿ	]h��>������ݭ������|,A��?	sߵV��+7��Ab���ߤ�5�z:Z����i�=��eq����O��S;��)}�h�rӖ�g�m�E֪����}��
iL��W*�&��+^̜�=1,��7ּ�^��f
�8��mY㶤^�}׆}�zfl��^C�Z���ތ���x���Gݱ�������,�ۦ�����XZ��S�o�6�����-,w�М�3^\6�Gw1i�j�&ˆ���b�����Lt�,g��a0�9L�J��C��^��,]:�q��W���|���s2}�-��P�n]�"X�/����<����-��;�Sp�1.�8����KQ=7G����o4�+Wز7`��2=x6��� 6� }s�$�����Ӓ�8Χ�����V�����^Ւ3��V^�34���Z{,)��Y�Ix�h��vӻ�ܶ�P9-v�+����v�?Un�l۳��I�D�W|��V��L �oWoAcZ�m�Ϣ��~�W�_7K�ȝ��(~�,}Y��]����M�OZ�����9�;�=�諹����'�v�TF�.J`%�DW���QNT����=�b5��+���/k�ǣXO#�~�����~�\���].�"�����
9��i��O!�=�����v��vd^}���Q��}D���g��ߖxO[9�zɆ��D�:D�q}a
-[*�}w+.{º�ۭ�,�4�t�B�?|*L���~2��H�6��< ��^�!o��U�O����ͭp��(��g��3��Mfuz,TɁ�˱�"T�l�',C�٢�J�H��i���n�P{ԏ����dR�g�űOv�Û��+��axe�$�G�uB��A�D\݁��-�ZU���d�[G�]/*�5��k�|{�şoK����	�z��s(\��Nn�{s+aۡp���D�Ҷٳ]�\��4��O髆�*�\�7��jDޮ��kjۊ���lN]�[�U�{p���.�ԇ%�7�+�N�w[	\Ɔ`���/Vs���QJZ�lkD>�")�}�v����ɝA͆*�ȫ&KrSg��佷��[|���� W
$
mnT7 {�jc3%c4i�ٹ�����憉Y(I;ĵU���=Љ�c���`R�v��`�m%xd���L��=�.�eI�����~��c���1�cb� Zo��Y�ݶ{����Vs%�w=�n��	��y)& ��o@{��|���;1��\D�aŁ��dM)���Pf���!�o��o�̤�.H��5:pUi�X)֕`c�j�T���0�����<���Eڏ�nOl޵W(~����[��VZ�`�"��)z�ʗ�b`��S�5"L	�ju��}��==�e��?9x��r髆�7��ឥ�L�U���y���.�<o-+b��{�������δ��H�7lH�3��t��2��]���Zjiq�#���b���fa��M'<�l'w��<��#I���;_]=Xخ=�-.�'�h��ie�{I�C.�sd�v�j����F,��>S����z׾��F^}sbǆ��t��k8�||�*z��M=�^J
�}��z����&\�~�p�^��_�4�nyzBz/C�u��7%�xQ�U������WM�_-�17�xX�W� ��G��4�T��>���^��j�4p+ɮ�,�p�����O�jڳ�	�q;�t�Kd��b<1�FLQ+(ax��`�v%O�e�@6M���s���	/�D�f��ԉû|Q�W]>����h��J��P��w_�������k*e��e�:Ӿ��i��/'r��׵�Š֭"}A_s��/���].Z<���L/p��G��ԇ�R��>�S������'�Ͼ����i�9(C�*����hK�w��|�%�;���ɮ-0��%��V!VE�p���#�o+{��9�6$4�,������C\����p�53(Rŝ~���M�q��o�@��1�TO�O0S�,U�9�-3��:lnm�,�����qg�����a{'�>�!g�Y�����P(_�<�z������?WR��Z�<�6}�(�����[~��9�=\t��G�/+��[X=�_e�U����PBޅ��Z���|%rݼ֠�U�ٷMiԪ$t��#ʅ܋8*,�yiq,�rٙ���:�����V</��F�MBl��O=L�}Yh�=5qe-�C��%@y4Z͓�sJW�����b�m�Œ�M�g���m�Ეdhg���K�EV��k�J��Vz�^A����S#���Z7��b
�f�:�z�V� �k~�t�cv��X��*�@����m����P6��T�i>����}�0ދS�S*,w�<u��e�4LA��o4���8��͌�_�v=^a3�Ӫ�=����n���Z��-E=h���f|�o ��7�c<p
�\N������.o �P.���@�X�y%o��n�W[en)�өEyd��<�g��D��⼠C��V���w�T�n�6�QJG����υ̿��a��<CC��6�"f���<nesY���C��6�S�Y�/˅ꚉ�ݠkW$����yB��3�ҙ�p�k§�ǽNb�.��3�ۛ�����KU��7��x���t!f�V)s\�g��#��>�FY7ts=uVMv
��&z�>��u������u1i�2+�r�óс�r:�{�\n�J��w�֊!ŧ�b�gч;���|������ȃ�oW�5gF(a�.�9�f�/n]1�*7���ᬯ>�{رH���K��~Y�ޥ�e�J|�B)˶�%&�d���uP�lNG|�<��3{�fY�����N~�8;uV��*���X���W�Ԭ��o��H-�������VM՘��ܻ�o�y{ML5�*�)1�S��g�}�޹�]j�2�}0��~��yW��e.���ە��:��"��R����B�Tx%(Suī�'����/_"6vU�%�L�2�h��KxB�"p�7���M�A�ӳ��'yy�-vnk:E���P�A�Ҵ�+��$f�V!��%8�i,QOn���ݙ����XKP���,���Pސ�ΣV�[�R�P���.�1C�07�ˣ]í5�i�`��;f=�֭�Fb���x���t�tj�2��Vr���ea��e�W�������L} �d�^C�iH�473-T7�egV z�ݻ�j��j+�7�eag���oUѕgj�,�Q�0+�"��t�DO"�ō�o7@!���+%�f�FD8��6@[�΁ڧ+'*��na�h#P=��d֢�|�Y2�=���b��#y*�O�n�O�y��^4�M�c���Qo��\?	�
�b��&���:�v^d;��qYԥ�U�'�ݮ���4���RgQ��5���jyua�Ǩ�����pKϩ9`���ڝ��C";}�
/K8��LtwV03ݰ5/Wѯ"��v4�bWQ�CK2V��&M��R�(��H��+ykS�5d��D��4��k��2��36�f�C��Rĭ�L�^�K`���ջ9ff\��<��%+��+]�Ӵu�N5����X��Hp`g�b�n�sH����) $W�����G
����[����tډ[�f���&A����d�2^V�T�h���˾{Z������iM��u��(���a��"kACP��y�	F�ϲAdY!E��y�
Y��Z���\���ݢ^���H�4,I���V��н	�8��V���WQ�]�T��l�r�Yܫ(,	'����3��������3(Ѵ2'*�|{AN�O���vC��EE��)[˩���N�������#�ܜ%�P۽y��)�Z��n�[RȎF��kլ\c�">�RmM>�mq�Yh�����lSo����r�3��{Q��v�߬<�M�Ri���6u��b�ј �欬ˡ|��V>hl���ݖ�T�lۺB�ܳ�A�s+~�ˮ�C��xfB6����,ZŴ3Yz6���Oo�
ҁ7�å��xe�0@6p�u_a�M�Ki��07x5N��������T��	2�:�ξW��R[Vݎ�҈�7���)-�y�����	�������aI`���w�mك)Y�V	H�n/��;�����a5��v�|n̳ֆ��r롸���C�V�Y�"�{�˙��-]K�_�Us�7r��6:�W�+J�T\�s��r��ؽkX�X��Q�Sx.��/*�M#�6��8,3���f���f��e^��c�0���mc�3����t8jD�rh����q6�����:�d�G`�N)�$9�[|7�n⭚�)f;g��t"�s/q�8q��d.B3�tT�ݬ]��IwFf�$`��~,��W��$S�,�$�%��WLF3���Z�����Jł�mRZUU )�Rbbc
�J��([hѕ\Ti&*��H�F���*Ƞ���)m�aX�ڲ�*AE���J�*�mUQ!m�E��B�(�XV�ė,����2��kY*,
E�*
E��e@U� ���X�E+
��q��*
`�\��DAd��,X��,V��XE1%`�%jʅ�ŀ���nf8��TRJ"ڵV��(KF�T�JQ�ܰY�#�ܸ�-�Z�Z��R����d����H��.Y*T�Z�0����LJ���Y+�A���c*������j���ƪ�[XҶ�XT"�	 � ��*	s��X߹��%���;iI%=���f��L(�C)fv�T��Ao�/k�qハWtHV�ά�iS+�K�}Ͷ�n���)f6t�����Sır��{{�w
�7�N��VՃ�mH������j�s�0�9νf���Ϻ��Ӄ�<Gݱ���Z1�Y2!�0;i+���X\u�	�ʞ�7�7��ca�\ ܶf;��O�j�&˄m]a���P���VZ[JfJ���NA�uis��}6D�y�6��*ء����b���.��̇�RޯE^F�Ey�&��i�ŭ��f�e�ym�N�)�yyZXi�*���,�¡&��Ǵ��d�9O�v
啙�{BERj�-�pi��ڱ�g1�5�z���/>�����ȑ���M�e������p����s�n��\gp��QI�:��0R�/ ����
r�)�z��v{������oM*Y�у�o��q��mB�X�H�v���$�^��q�:�d��;�(�y:=�^n��0�~Qo�y�K#�y�x	�o�<'���l�y���dئ��x|.�r{t�t�w=@���;-���xR�����/��1m�{!�0(va�ZX��v�;���[2���l�L����hT���������7B��)��
�wx�'��r �.��5�$�׸�O�E�)S�MA��v�����T.��^t�͎r��%:$gZ:>�r-Y�V�˜{�'c]s3�+��	��볼L�e&�I2У9�(c���?U2:��D;C5�����Y�A��*d��e���%+^P��zx�>s������{v��d��Du�K�E&��caȧ��k�t�0��v��y���B�~gN_�����"���0����M�<{�!�&�����*j����0�/9 wW�t	�'�tvzv�;���U�@u� ����ץm�f�V��3����^{lcR��S�f;^`�>���a[מ�ǹiS���=����f��J�ۯ	[b��J��Ip�aF�*��������Ɖ����\��G�,lX�i�9m,o���M^G���||q���nr�y���bK{���S1+3}��ە�A�nË��4ȚS3��mP&�=��k���y�G�M��|���-X��_=���0��t���^	楽[���Ma�n���~�lE�N�֦{lnVZj��)����L�|U��}|)ď�R$��#�d[��{$�U�u���ͮ:#5��L�y].C�Mlԝ�J��������J^��R.����ߏ�7�x���qw�@�yE��Ax�R���=I���m���g����D\k����p"U\8�7G����W�R��V�nr���25�&�k)#R�Ԥ�3h0���y��!FCfA���;�Y@� �f�vK�.p��aG��JI���U/��u)���|��9��J�x�*�%�;	�P����=ZB%����[�x<�vY��	��QߞT�T�3�e����5=>=$��u�IU��k����A�aIt&}Nd��+�=Z9NB�s�Z��B2��;���N���R"y��d�M�.n�1�^I(d[A2/yP{�eͧ�R�ֽ�L�iŚ�2T�(����f�oA<e��{V�A��h�H���B��p���.O>�z,D���U��Eq�b���◝����P�L�P��	o-$+Y�J��\e��p�mf�σt�QRV}����CU�}뛾��^�^Q�qC�][D�z�(aەDCa�4%��I��˹���A�g�M�$��z-Q羓e���J��j�-0lHi�Y����Y���8�����n�݃��{�덣��z׭i��vz.k��,rX�~s8f&udx���ۅ��@�z������{y�K�8}[�φk���KT
���<���X}�ǳX&ֵ���Q���sg�����N��&p-*�O8 ��-)굣Z��b�t�P�*�j*��q{��ǵ�-w]�Z.�lyf;���4`�eN�zG9Ri�TI�^�X�M]�m�Y�39,�Kz�GS�8�=�� �8|��}2Ĭ�|Jh8�;��4D��y�X�+G�i].V=*������k�F5c��6+5(l��>�~wNz^�=$]�`׷s�0��/f�q-e�p>;*5ڄ����*��K�o��-7R�ߐ��zd�!s�>`Z.uE�*���oP;-gn_����,���hr����v�x�ǒ�t�B�f��x&yAZY���(|K�9׎�����'J�0*�ԎK礽��]����?y!�J�Cl)ɥ�Qt�Fg(K^��Bt�g�V�ʪt���>UP̽�O]�F��I(f����l�,�SW�R���d��[��j]��f�Z���v��!Flz�k�ċ��2,�����'A��-ͭ2&rs�7����K<S�%����̼^�9j�$J�]�t�P���̼�t��B<ҙXw����/��"��
�[OE�4'�wƼzX:t#YQ,���B���:�(z�+L��f��龍�K8��^�p�3<{������"�G.\;�e����B�qWI�ֺ��^��p��fc�\����Z��٦w�M�s=�R��ܬ�f�ň���F�m�j��*�}�c�SՂꨞ�~~�,t���9�ww�)���;�>�<��s�5�����Dvl.�En�JѼћ��>4���zF
����V�b2�A�ʋwsϝ;�v�ҙ�W�{e&�I���+"�˷�B��w�v�˳�H���F��!>�	��xk�#<�Լ}�X/j�e��EloL��P���c$�֌KGJU�[�gv����Ԣ|U���8�ۺ:��,��z��J��j�z]$�
�X`���n�sU�=�Z��+qI�٨�.b5嶑G`�co���g�e���<��ڶ�CLC���3�(*�6t
������đ�)��7gk&:�Yl����7�O��hp�,hƤM���U���哱��f�i�^��:�Μc�s�cuz-;csr�9�)+񒗝a]�n�3C-o�}ϲ���"�Ux�㼘Ϸ-����Z|��3���YS�Ŏ��Kq�{x67��i�\�f%y�B�E��|���fC��-���(G��q��~�vT�Y��җ>7F9J�%��ڪ���W¡&�u�X҈I� r��Zr��l[f�[Sn�Ct2L�/r\�����/�a��D����ɴ�[a�bt�t��;:o�u�e3N�s�U&k��2�wBe��'��/�6-4�C�F����f-��|�qd�����f26��=�g��=^nl�)u6�X'i�h5��5�}�S��9�̔����p2�ٴ��u�M�R�0Ze-ɲ��vr��[�V�Q�le{�|oPmY�uA0��TF�K�`��DW���TpS�53��T�qt4�ud���2}9�96��,do<l��t�G]Ra�4�P�����}cO�
�U�=���;΢��+��7T}n���v<G8�,����z��zɆYN�����]�_o
��������5������<>�0k�
^y�(_��Z���p��o,��o4J���ok�\��`�^J�J�gk�س���Mf��E�2`bU:$�k�f��F4��>�Dx^y6;�3֒Yґ~X*WV+m�=�b��i�87��L��W3���F�1���K���_v�3���[K�]��I&w��V*P�gXf��g�L�=�b���lқ�ƕr4�i��t��.��|��2�޽�w�Q>v�Ow�y�n)�,{pz�!*A�Ѧ4����zn�y��1���w�Q���oc�pE��,�d��X�;�ץ��:�C�����Ŝ�-��Ҭ�8��P�=���֠���P��r�Y��[=�(iӧ�3Mg����݈���B�O���u�[R��=c�nK��sZ�Y@���"f�A�XD�1}��\��ovͰx��6n�u�+e*�uܱ-��Y\�Pt��i�Xցث��T�<r)��f_+��b�'5�9kNw`���U**XL�k��H�owxc[ڌ=��2%�	u9x:��xnW�,�`�"iOJ�uc	�W����!�}O��F��;\J�C)y`.s|���D�z< ��@�^	�_�?��ׯ����.U�7�5>:��YS[d#��;-!�Pq������GR$�������n1~�=vT��6�`~���k��ky`�P�
�\����7�I�*0�����Ku%V_mOHɮ�E�=�P���#,d��C�[��'ɉ��J�x�-5���l����n=�Bk;t�=ɁZ+cƖ�,�zY!�o{*w��
e������ �ՙ��A�x�4z�b���ύ��z���y�9�W��螮3Py9�LP�����t3����m=�S)gw8���OY�m���(��3�A2*����2���p�^��_�|Ӌ5y�
��k|�c�v�
9[~cX�L�׺�쫡ΑiX�P�˸zǺ���y�= dM��j��ɏ�]�s�w<u��@j��!)@x\�E�b���ZHP�k��u�X���rʗF��~���{��h���CvG�Ӽ4׭-�Fc�R��Q�nX:��yǂ*��.�e�����
U2ѕ���2aƓ�X��;Yo2�÷R�T`��m���
�X[V��Mi��LH�5��U����)1bO��:��Z`�Z�z�g�����0�NaȦbꃺ]�b��m�Hi�&}�J�!���WyX��m״����.�����Q��.�_�o.%f�R/�{��-0d)�.�O�x��A�鷞_ef���q�gw�z����MX�3��^;ȸt��zX��*��0p�L���#��7�h+���|9�U>�`T���/��K��=�m���,��[�,k�m'��j9�Ƌ�z�m�-�.]8O�Y1����i�m��X���>��%\x=�/���U��ۈ{]�pu~�|Ⱦ��P�M�;z�b�➁q�F;D�B��"q�;�ˬ�_b��]w��!9����ۮ=��ϧKPɲ�uh�gU�0�髋(�4�<�NZ�_�v;xǦ��|���)X��`�
��V�e���Rǌ�X}�����<|��1��)C)9����i.o�\�C����asQ+�Y7���N��zP�.���^�P���J��t���ZX�>:�U�WU�+�����M^�u(�>�i�y������3Z�ۊ|f�^!��b���8����2c��ǐ3��[�j�=�JG&�c�V%
H�-�,�:�Nk�>�e Ȩ���'n�5_���rGû�bs��]�{M�&��Gc
n�;f����z��_ۑ9���2��*^]{Qn��X�.U�����fg;�[N���6����K[�����i�X��}�{��0ײ�+%}.�:y(��e��)��N��K�i�Sί�'��o'������Xt�dy�ne;\p�A� �eD��5�ke����Ӽ�U9/���A�����K��n�~
fx��u1i*�<.\;�e�ȢH���\R�I��r��ۼ��q�z��ǟ+q{픚��0Q�+"�v�zCVt`Pö&]�p�#G5� fN�l�+�Ò�_��tun2��C�Y�����>ޘ)+r�a��	)5��f&��h���yMպFloD�FϦ�*
���/�w��ej�g�f��_o�.��br����T[�g��V��3�n,�;�c�wxUj��N�*�P�n[���qUWI|f�����t���Iuޣ�^�A���f<U��͞��]U���}1��&��eɂzq5���v�;���/Lj6:���]��>��dC�����I_�(WY���|덝���z�ӵ6���͔@���;�P
_t��@�8�+E1@ k��T�ho�x{�f턦Э���g��<h"�2��y��g*/C�Wʝ�I.��m`��\�{���0�+��Ԭ[ܳ��`=��*�[�	 �-[���T�Pn�r�v���2ǈ��w���A������-,����.����5�رސfq�W����-��W�D�Դc/�gQj,�q_��d'�?(Y�/'����p.�[��vN[.��(+�E����$�z?0�^ :����(�:�>�c��F���7�޹��钱�ء�_����*��Iy/�euYyJ���fN�H��By{����HbC���v�E�ݞ�����a϶
�Y0��
��A.I�%�L�\^�x��iRm�Gw�z�Bo�V?#�# �dз��V}�<��-#��@��`�K��ܩ#��^oA+�p��>���}R\����w�v<E�޳��o�=��I^���o�o��g��^^{�'���g8�#W��G�g�OR`���b!X�R׭�e߫��X��}��U>��3p�5�I��#�x�w6+w�y��K~�������ٻU�{Dx�{[X�wP�Q�e��}ґ~XJ�*Ꙡvע��k��H����D2�v3�<K�b�&�����HfC �-f���Snw	��h��k�%�u;<t�\e.4e$je;En�6;c��z����:�Z���:r�X���XŜ���gq�b�2���'��f���b!;u���J�ۮ!��j��<]����������q�^�T��{T}������P��)CR�Me�3F��m��R��&��R�Ո��]�}��H�щ=NVB�W���69�Ùr������ hmVf�-�S&=����F�Xu�tU��wݸ�@��h7zӾ�#��0.�ز	$b�kh��yd'Ƥ��� �˘�n�S��e=ܴP+h���)WU�<7j���ѶD�$C[.�5�D�r�f|��a�h�殜OK�/"v�7|!`�����
ϰJ�k,V�����<
AC��X�=��Wr)i}��;En�s�ά͜L�AjS��5��\y�:�􇨳��9�*�����0��ͭakR䓣u�R�r���Ts>˵@EwՑw�-�Yh^@ECf�����8�ڽ�F�����U�CmI�i�G�2�U�A<�8i�<;Cm7�r˗CY[�����������[)ו�%���vv�l>�
式�b�%��|w�JPg�[+l�����⚊��L̸����V�.�y�����F�yL�������*��Ty�E����ՠ��V�:K�Y�d����`��9���)�i����$�qw���S�m�o^�*�iy���($mD��g�iJ��s3��r&�u^u:�tԔ��)b�;��ݵ�l�w��x�m�x��K�Y}2�|Q�*\6��7RRl�j̞O���;1݁RU��]��N�,}�L�4�d��Y�m���d�y�)�8����QH9̩-�X%�>-�Z0eZW��8�͆��D��*�p�">¨���x�\�E���U�FÝg+R��O(��}�!0�ν4վ�����5
�Kf��m ��@e8�Hw6z�5b�t���ee-gt�-Z��37g-ޭ�:�1Q.�ɔ���<z�+���*����gqZ�9%�|t=����E�uڀG� ;9D��I��f�O�96�7{��y]Aٰ�uW:V�)�tb��{ÝN�}��r�Xոr���&��s��)�p���ۈx{�(X{��[�%�:��כ�FՆ%���a��+MH���qr�法���̥ƌ���Ȁ�ǯ�jN>�ȰUs!EV�������k+f�q`���"5���{����o�l�8�S��R���X9��2�l�+��蓴�v�Խ���uc�1��U���%s���/vфA%(�v�x��4u.��Aݍ���8c�;X�#^�`r�[�S����$I�c�
3��W���'���!xd����*�脅�D�κ�VV��W���H����jbU" �⸌���U�+U�[J �V���ņ&T��U���F�TckeU.ZbfJT�b�J"��XVX��Db�,YD(�"��((#���(-q�P�(�X�(���,b�T�*2���#ʩR�Q������`Ғ�B��F*�*�V�(��T����eQ�mQ�J���#"�Z�$X�(�[YhR��%VU�q[�"1J�T�b ��Q���b[TDU�0�&[X�6�)6�Z�"��(��Ek(������UTX��+b�V
+l�LL�U1��eDTC,����`��	e���F,�-�Q���+r�B�1�Kh��ֵ��*�`w�=��|�����/�_0V9Y�	ˆ(�eXw�͚��u9.��$�i��3�:���&�^<�\��К�����j6#u��䝫���ե�?}�����������t��I������R���R�p�K�{�i�+V/���8U=~]���VL&�Ѝ!L��t�}o*�ϻּ��·�����?he.=���=�Ç+�����r�����_ϮE�v�8{�1��=~����ms�z���t���K��;�V����@�*YCX�E�� Zly�id�[=��Mc�Ӳu��^ْ�|ό�jiv�I�%�d�lc���� {vX���R&����;k�;��I;�kˎbc8�b�W	�\��|*�f$֕�c�o�����N�L�^]���_g��x_<����0ȻW�y�ܬ��Bi�6��V2�7�8��)ts��G�d��5����/�)�l�u;�U&����i��VZ�-i�͂:��J���f��yj���z�OG(�7-���c�S3gZ1��X�	{]��X��	��\�G�����#t�Z�kk���p���ED�q]ɘ+ �x��e��K$1o{*w��@�w�#B�~i*��]�<�
I�e�ۻ������1�M�3)�ͩ�A���9��/��e�c�2�����ߖT��҂�ɸ�'�Z%�n�+������@\3,��{K=u���p��+��*�^�A}d*�僭���ÙKp,��*hΰ��[9��,�(EP&�s�^�ԳZn�6|L��^F�\Y��]���ɫ�)^����r2s�Z���]�/vt���>|N��P߸�ty�o��5ΔJ�S1�"��Ys��l���o�~�;$�[j���g��^o˽�yLt�
8TłxPvZ�#����Ú^�����@_�
��-���q7�;�j�u7e�e{W��\�E�b����B��\��u�^[��q��PV��9߲w31�k5�՚�������*�'����(aؑ�%	�+��W��ao��W���-�nh��w5��a`��l�����!�pi�!O�oK'o�f�5�q�n�nl�QRC���@偯ݮ����_fz-�O��c�}
�13����2��"e�uk�D�fY�W�w>Tj���xg�	x߇�����O��?WR�x�i��7/R	�� l�!͘�L
m�oqk��me%L�S�{-���h��Ȋ����վp8+[�.w]��;m��}6L�[�u[ͺ��J��K�����܈mj����f�̏$��	���l��q���"�Wr��m�k�sn�6�+��9Z\���u�� ��N���J�)���"�tLAm¦��8����Y���,�Wsͫ2_f�zZe��. �Qe-����.:��Ɛ�&�;dɑ�[����&�8U=�M�fc��w�,=C&˝տg��ϫ-^�Qh���>�9g��c�ܝ��'�↩C�
��`�T-eifXws�>u,x����}~��+Ge�Jrqꗾgdt_�Y
���2���2.���5�F(�M�a������o!�M	�����_P��A]LOt�)���G�
�8�������T���l�,�SW��Qd}r��c�d�҄}��n��] ����T�{�ԋ��qm��wf��v�.��Ww��n���������ɦ��kL���o+��L��	"xK�}�����e����n{�=^��.O�93�л�})�Ӆ�Xt�zfq�}=o|p�z�D��5��^~4�4��{�֮�jg��C�zR�/[��x{�.�-"B��~~�၀>���Wko��O3.G.k�J��[�ׂ�>W��r/l��`�0Qq\A��]�RGÔ0�y^�e���ӋzS�V|`�F�!�P캭L��Y�ޥ�邒�*N]�o�l0����Ls|�����qjϞ�~��[�H���ZӖ���(�*,֠l=�F�w�'��N��ad|�ѷ]ۂa�AMK���
�F�9��K�Ƴ��������f�Pôe�G6��N	��5
ܨ�kG��/�^a��Ŷ�e�a%	�(���D޴t�ݗl�KޢF��g/���.�}�����f-K�f�q��P2�;�7B��%�*��0�*��Y�wz��ѳ�50�|yT���-��X��v^͕��vAv��;��<z>�MX{p�;�=�q ��G�罇p�}����7_o%/��R���C��w-Ϋ?����P�Ӏ=�ɻcuC��_��<7Bc�ӊ�=dn�w��Io'��^.��"����A�r٘�ŧ�B�/w���6.�yZ�zQ羛�;�lڣ�Um��L�Y�63��8�;�����ޡ-3瞃��˧o�x5�t�ꡄzVm�ԩ=Zm�U�T�}|*l�%�����_�[�y�o~"��Ǜ�O�������^K�;hD�)����)W].�h�r$kn�U,�7F���8;PzR=x�y��٤��2�'��d	��x05����#]�|3�º��r����p_#�m��~{�ϭ�U���ib����|9�2��wh���1�M�7�������k���3n���q�M�xN9�2nzq���~]M��&���i�1��w[[z���2�O���t���ؔ^���z���B��Zlls6��[���73����%7�n��7%,�i�hb�xN*���v�r//f#�Ĉ��tr_Z�"�t�VG&M�)���e1�����c�~��OK~Y�=l�}=d��b������T���& �"O���(H��V�=�v=�)y����ʯyz~�4ۅ[��@-�9���:���t��l�H��I��#�|Ϸ6,����Y�3�:�0:��EoUX�j~���8�=��1�V�07brɂ������%�,vA�>{����iV;�K�t	����\pq�{s<�_���`씈�6$���?}޴�7�O%�=�l��E�N󟗳�N���j�}m��oK��K&��,Hi�z"s�*���aʂ�j9��g]��Y�_��L��;O�G���uaCP����y����c�<F/�o�,�C���v=v��}qbs���\�;ۮ�x{(�R��J(u/`�z�_���ʗ]O�!J��V�HUڿ��X�;U誇Rȡя� >��A�vN��i׻�k�J4�S8�aG]�T�V�-tJǡ��`.s��;�	4;O���]�O)5Uh�2�T��bmjҭ�=���U��{��cB��A�I��oλ�$D��<��lp�j<��vm���Ѱ�3��j�L�WO�A���ܟL�vHr�H��{�w1	��.���y�	���sL��-���A�����o���Q���O0wap���OɃ��{�󱲔gŊ�K�F��^z����Y[n�72������o�`h�p�i�Y6�N�<�6��њ�X&T<�� t���̙����~[|׼���C'%>�`񳧒��T3};��Kaς{}��kɔ�\�G��'T��t=�;�Y^�G@���y��W<i`Յ���`����m�7��Y-����^��0�P7��ԏ��4O�M�8��T�ޞ��U��~ðhi�٨&�"&d���9�q�����r�ŝ��t�8:Q+�f5�PL���<	�6��K�Z����K�$�t6�W��XhM�4��^�z�W>��[Ȏ%�^�~��ˇ��u�h�F}�|ܬ(��9A�j�S˅�v���BZ�p\�E�#�I�Y�i.�-w�['`w=�٠=wٙ�����KSx]o#�O�5���|;��m�z� ��nU�&���Ư�xC��I��z�2��n#�����X��g��Ι�z`�a�F���Z`�S�Z:Y:�|EU�����^��ۯhXyVO�;����ӷqT ��"y�p���y�������e{n�V`V����ݏ��
�k�N�d�c�)_�b����Ҧ ���̾��#�I����u�\*�:`��p���ұ�7{D�����1�7�;{�����bk%5��Ϯ.��g���{��%��*��0W���R��	����}<��ҳ��GM�;3�A���+���<��=�V��}Vj������,N{3թ��V�ԧ�����z`WZ����疲��eB�Z��(���1_L�c]��A����u�<���TG��n2��/u?�n�v��XG�v�5ډ��0U�]]渻Kx޷V>8����K��-?h~A�6\��gs��FM\T�w�����[�ϻ$���� R�+���+G[ �
e��,��r�Υ��k�����<t�z(���Q��ԏ*�%�+�G��2l�4��V�㎸<��'[�N~�y�3<Wfxh�_C�1�E�A���i�Y\}��Qq�$�;�!X���ϋ9��R�K*lh�z�u$������z���3��"QC|�Z�u"�<\[A3,g@/rmA���
2�}��h����?T<�9��z��b�Aڸ���h��@mu2�L�8l�w�N]�]Kˊ�ʞ[U���/T�g_��}�n�U�Y(G�R��_St��jqк5F�\�(Ϛə�����eǇ4*��i� Fd�R���+�D��b��/K2n�Qq-ו;vN�:y�}u�:@�k'-��8� XD�Bޙr�q��D��vqPn��]�x�^\��9�g��Ӓz�!`�� ��Y��Tqs۳^��w�v5�Ė�Z�
̿�\�zR�,n�~S3ǃR͍�xB���`p��(C� ����Y7��Z�$A쥅X�������r/����0Qq\A��˷��Hj΁޷Az2�M����x`�}���e�Ep�iv]u�3~Y��޵oK�9P��Z�93*�%�ykj�Dmoz���t�ʞ�#�^�Z6}5P!������(��>�\�n���cb�#�W�)���_K5�GKU��w�l�}��?�*�����3�1dѳ�Uz�z��ٵ|��e��	��	"A��+'"�
G�罆�
��䬵�Wn�0I���9F���9R���?��0xv^���6t�{#7�=�iݽ�,��L��e���7$[uύ�pU=Y��j��_��b�7-���b��/�y�#�U{e�����{%�$Y��U��_�D������z�/�Ү���E��;��a�̆BJ�b����,�S���Z������y�hf���5�Y&�Vow���1CRD��ǘW�����ͦ��.��p/SYgVV];�(iv��sWؑ�e�8C�7���:K�4�
쳙"q�)��f���Ia�o�'�\�c74ۉӮ�)N�:#3�q��Mf��J��U��Iq�rɫ�P���l���a�cGmZ�$�۴����we����,kXm��V#d��-Lt�Eh�O} K�F��puK�˷.t����4���y=H��;��C���
�Y0��TF�K�`�[�!�י�#b���G�<k�O�ϯ�⣕%�^
z���&����V}�<���)�v�,¬)��*Q�[|��G��%1vP��yc�3���^S�=�Nǈ� ~�0A�����}O-@��CdJ͟YDϽ)h�������A����=�0k2�|�/ˤ�W�����ѷ��$�Y��ˮ?c8q�T2�GJM&�
�X��g�����}��o��r]��xH}�^lQ���/U��6��->��'�,���(���'˖;(d��ng��;��-�g�_'=�b�;}�IF���lR#�ؒ�����<����}T�<s=�Ħ�D5p)�=���Jo�`���@/�şoK��K&�:�lHi�z"s�*�쥈<��v���Y����et�<n�Zy=�{�s�<E���[�7�Bh��l�{5�h��7 ���6�WSjb�STT�`�;��/������3N�����s��Ms�N��L���gT�yw,=�8�ٯ���$�蜤dm�ޥ0�S�W���eK�S��,�üp}p6�x�}�gK'��=^��FU���l�����Õ���j���&���n`g�nWbcn��� Z|�4�i2���^�g��k�V��:kM�����Inᄺ�^v���q`۰��3^޻g�5���*����ȹ���K��oٴ<h�s+��^2�`.�0����N	�OIi�Z�W�Л�}gI3�e������~L�"�Nr��Q�B�R�E��^z�ؤ��c�)o�9�TԎy�q,�T"�M����Z\f��E*��`^4�d9y"��ڮ�i.c�T�l˾���J��C7�v#2P�|��j��*5�L�z�F}�fgg
������;�Η>�x�xK�d��z�f
�\��3��w[]�;<Ơ�*��>���*�t;;�Y�K4M}ΔF����kz�<�2j�螭�9}���؂�:os��_�\��z���=u���hu��k�>�)�vQn�#�>m���o��忿�$���$ I: H@�D$$�H� I*���	O��n����6@��$�� H@���!H��Y��u���r�	'����O��������B���D	O�� ���$ I<��C����~D	N���_������~�t��!I���~��)��	O�@��$��B�����aB��y��ig�^�1 H@�c�}��	'������������?���	O�c����$ I?���D��������g�����	'���&������$ I5���t@��$���vN�/�~���?#�LPVI��xr_݀���A���y�d/�������p-�� P @       M����R�      T�4h*�R �    T��UH=F��@4    L$(Ԛ       4d���`F�b0L�`TQ&�ɦ�0De��Ѡ��D��;�7�D)��Far��ɉ���:�"2F��~k�0�"�\�{<�~��W�/�y�:�G��ߤ?�;K$Yi`��AS
9��ϭ׬�!ܩB�n�KP��*=^m�^��OY_��ͬM��$M�( � $�� 
H R@R@Rd�% ��%%%%   ��R@ � @ 	(���j�ȷM�妑���bSFԼ���8o_O��]�Ł 1DQ/�6XV]طb���	&xL��,Y��5�1�A2b1�����)�	@Z!'�4�$�ـ����a��I����bŤ�nb�ٴ#�|#E��-�8`am��
D\%ú
o�^u�;i���~S��1K3=4߱ӻFzkx��#5�1�W��;;|{��qlg��|�O�˧��.�}��tpi��
�<��oN�x$O��Ds�ËmD����a�0�����ъ�/B�b��/_Æ�P Z�F1 Z� �b�a0VD�1�$�@LN��.�JR�P`���R�	�`V&$ Z�ĂR�� Z�j�8_����x%UIo�Ma�*��#�9!�n0��ED�[F@�%!8 ��BG������v�mػ��������k�����K� C��?5���	*�2c�NN$���!۔=�ElԡjuTk��X�7)�2`�hy�xɋ��Ss�Dl�@��^��E�y%j�\�k���6߯~|�7Y9�a���r�l����m��m���� ��06%I�hd�������:e�D�'cC&�lP�N�F��XC$�f� ��P�T�Eo15a��{�;#�wn��h�mkAQ9�;M���N�5zB	�
!fii ���U���9B�D�U [ۄ�G�����i�[xF��0�0������߮m��m��m��p#�VR����u-��U�;T.|��Y7A�omS]/E�R*(@O��	�Öv&�w�EŁƪ�ѹ��	;Y��N�Q�q2f�]\.�Y@�b��P]B^�� r��Џ/�{wx�m��m��l���b�{P�Ә���"��,����U"��@T�YD����hh���R�÷bBlX&n�UU��qǴ�P.D���q2bf�����gOG��!��m-��������DDT�gWK�Wc~�6�m��m�ޱ�����T��Y�~;Cg�����ѽ �n�*/̾��l�ŀB�f�����* ��1sV*�Q�;V�x@�{J�Z�b��L���W�D 4�=�3F�ѓ�o�K6T�6�m��m��t�"�<}�({;�$�@IM�Q�`�Ѹ�d��y^ ,���b���ae��C���6��*���"���C-�+$[��P��ډ�T�`�@31	�2"�G�`�!�����m��m�ث��)ج������@{��q{L�SP����"�9Q[؁"h"f�lٺ��t����,��� ��4!Aq@BQ�9ձ}d�Y����>5m�I��)���m��m���F�ϱ����cwY[�1jf���[�x���Ks�0:*�qo��s�S��'g|��T*��uU���H�V�n�O/#�h&��$ɐ�-H:"���E�J�
>*o+�j�m��m��m��y�E�g�����A��Je����/6�TF;r�nkZEK0�fv����Jj-������Q,l:�����2�����ԡW��j����ܱ�T���/i�m��m��m��n�o�st���lI�yxӁ��3s�o��6d�3��n,�Y�j=��I&�ª�p\r�ݏ��s$��b�=��v�����@���F#��ղ[j�±"A�����G�<�b?ib���&13�̙o�5�4]��&��3��f�`�˒�X�[X4��a��C0�5�g&"cca���<5ΪSE3����Ŋ����ZU-��*����J�iT���m5S
U-*���RҩVER��ZU-*�K)h�ZZYKKJ��R��hgL�I��50��Jڣ�5}Ř:��6�[��y�&hĘ�#�ϻ"-����Z��^Lt��w�m��G&?z1�CI58���Ubm&�N���%5у�Di��uq��#���ά�L1�[�价�{c	r���56�;o�bH?r�^�9�O����0�x<a�M�W󅐶���;��}���;��O��_�X��N�/�e?�=Oo�,����I/���?���pzO%���Z=6���I$n�7����I�>��2Ml�4���$}��MZQ0�V�c3����=����d������+Y�վonS�.��19K�g�����eh�*�,��ft��I�'�Hb�N&���e��鉖Nl7�1�5z߷Vh�����M�6�my�d~čԘ��H�$cE�%)�sc�{I�����oМ��F��Vg��i�M���,s�$k��~f�N̿u̟��ݬ}����\}[�F߿~ILD�j�L
��;�̝m�<�������-�}�؛v��<������a��{[�Y��l��ڨ�OYϹ���g�I��?��p�z� ���(�r���|R���������eU��~�Â0�ċ{5�$�+'�$��O��R�}�G��-�;�\�4��l���߇&тG�}	��H�m��-�T����nSs�]q`#X�1&���wfH�z	�Ѿ9U���cK��.�I��V%F�M����R[�q��\����N�#���0���y��zos�N��	5K�z�b�����2>3G�=_���O��t��l��^1��i��4$z}���m0���Y_7{�X'��{gS�Ǻ��h��c��l�/K��?	��:v;ohJ�z�q0����$q���A��F�"��~��Gޝ:���|��莾�L��{��7l8U��3)������_O�C�7��h���9�Tn�r8�j��~�v�|9r�8&\Zv�^�����+�����L^q��s��4:bx75XqS۹���:�Ƽ�������eL�<6�{�Th�<���X���:���bX�T�I��_�\�H�_���=��O_t;����N�St��o^XM�u�c	?N3��y�ל��Gl[+�1K�VH���9�w��w$S�	\�� 