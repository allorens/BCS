BZh91AY&SY������_�py����߰����  a>�    �   �h      �8E$ HE  (PR�( UUPG�{�$UTT*�\� }@��T�c�W�{�׽��]��)��;Ol�2��=o{���+�^�ǶtBps�G�9�	�� {g�ѯA�@�P*{����@42^κ(t�` ������4�c*�e-h��yǎ�c�=8V���Sރ�Yvװ��;�cH���s����ֺ�N�L����m�o��j}�T�� ��|��O�w����&9\um�6�`b�������x*���ε;����˱���흇��{jSp3�۰=;�ݗf��  �$�'���΍i&�f�z��]om�j��]�ǏV�ۅ\C�GrAU=�s���޵�{���˞����ݎ�;��xU  /Jgw+�M��=;����r�ץ�Wov��+�lt7��=�ӧY�*��n]�hn��x=]�2nƋ�wm�lг3�\>(         (                 %S�c�)U�	�#i�4���C��"J�h� `&  S�%PMT��4   � d4i �*�2�#L�L��b0�LSU�2h�����=���ȞL)‪J���	��0# ��4d��G��u�ṛ�W9�ÎMU����k]:��<v6͚ls�#�?;36��1��m����?��������6o�wf�:}�7���������p��n�Ƶ,7�#t�l٦r���ڝp�pP��6͛�؞�AUUURC�&B�A���c�|6���_{��?nޏ���:�|:qxS1�X��:~?vD�)�d����+��#Qe	��a:'Ds�,\���D�9�1�JOK(J#,�$���'E��$�(f�,��'�@�1�cǏLx�x�f(�"I�$�U0��b�87	Bo":�ĝ0�擂p���'`��f(IH�RH49Q�#�0�&�1L�I�BP�\���f��&k1%��ęl�Ĕ�N�%�yʲd����fI6��9S��a�ٌɄ����t������ԔÖ�H�36a8�h��I�'�Ç�� H,b8'~���Yf��	��ZI�4N��K��.{1̄��Ʀ�t�sQҰ���Q��҄��Y���ChYUT�#ؓ�D_��I%�1��N�CW0��4Dٌ:$��c����1�DIcS1�Do�	�����9&ۘB��G�q� �L�I��b�������d�h��DY�e����&���ӦX���,�L9�&))F��0��Yq�cJ$b>��T�";�	�w�0�@���YҖc�(I�� ��d�`��&C1�v>���$1DȗDBP�Փ�d�A4D�va0±��8�Ĉ��a�CH�S-%3S�D��I�G>�(g	�4�K#�YDGD��pG,��zvK��͓ӈ�<��IFxNGb#>G#DM��e?C��<�*!�D��Tӥq'���p�$�i�X��N�|^�6���־�tߛ�8?Gf��F��w�Ĉ�r{��"?Q��L0�f8��4�"f�a��&Dò�Qgi$D�f0M3Y��b �&3��t9� ~�bHH"�R��dĔLG��n>D�ي�bH��������"/f$��1�'x�%�{1�1tk�	����&>��s&8#Q"Xq">��"��p~N�Gb�a��62cDJ�"#��H�&$v>L(J�D�*a
�/II(��Dr�$�@"7�gX�DN��pH�f�����"SC�P�\�H�I��"H�b�H�h��:p�ID�M4v�Sr8&�I�9��9�fDwbd���,K K�$�c�"��܉J��4� Iyf��?tK�ĢaY ��N�Q��t�n��M�#���O�	�!??BI�S��&v�Sp�ב:&�=؞�?,M�P��Ju!4ŉ�8&Dt��r!ؔçN��"5�H��_G�?5��ȚkșDr:"Iޱ2"9#�L���`��Jt�X�&'�%��Dy	�kQ6Q<�!ȔMb�3~�D����
��1f$�%�BpD��(��v&Ĳ��'�7�12I�'*�R�KX�4DZ��,����割J�Ľ����ԔxB1�؝(k�)��x�s&<x��pK#Y�����Ǘ3�#������S�1)"J��Ç�:'^D�	�bQ8p_�+y�����^���%B�<(��B��0��93�̦���Y�s�f,~�G�3�,��!��fm�yI�a��35	�r+�DG���2"ٜ8Ęr�fj:%=����$�c��F?Bh��'Kɖ�"���fg��L���JbH�3��y��O͞L��N*��������lfD�Y������qɞ��(����vbz#Q�D�;��	�f�8Y�",N�Du���D��-D�cW��(�>�1<({�k1)1�B_��D�":@��K1(��I�ф�$��ϑ'�Gj'�DE�$Mn&j"$D���Bu��7��#��M2c�Q\�(DN�2"cQ)���ٔ��91�`��'��DGa4��Ѽ�N�ñ�=+�O(~�DN��D��'����D�L�Q�ߣ�*&��h��&D�3y��`��~��,D�Wf'��:v�8k1=8r��Dr��`�f�8;&�����8&�M�gN ��BP�̲E ��H!��,N1��$%�?�.D��%�ϡ�t��&�;P�i3�PID�ID��"t����ML(���'D�dĖ@���@�|�Y�LY%	Q(F�a,Eٍ"�gK�:h�LƉ��I)f��tJ,HD��bp���%�H��]�%:%<��8�N��6I�I�_����'��O�&#�T��	�����J%lĿQ�N�+>��1�&��93�%ٛ8%32I�K� I�=���L�N�vgN�Y1:QYY�Y�N�f�&z#زJH�q"8a)�ز�72��޳:Y$��ؙ9��33)&�re$�ӱ??1��X��Nrfja�}p�5�(�^AQ�S)���i"�Q�`�32h�̦&\a#�GDJٔ�2�Ή|�$y�|��'&��������JP��3�q= ~~�L��G�����LOj-��K2c���'�9��M�p����DX�'��Lj%:4��%VĿQ�Z�D�ȝߣ�]B$��^�&��r'
v'�8���NK�r*��RN�M�8s>��{�`��:'~�i&�&Ήfv"(I�>BɁ�9��X�G����Ga$ϓFa�"?"\�M���pGa&8#�D~��8��"b����t����bVxu�W/���Aߙ�H`� ��)�8�	�;��C�)GX��i�iјN��
"�N%���Hji�܈��Ң�D�t�ޱ��� �4I����N'R�b$���aќ���T�RW��d��-���p��8COR+�OJ*;1BMD�&@��Y��4�{w�c�Q=ɉ/�		�1N1����7̘��DD!��G���b�8�&D%�@�y0�M;�ښkɜ'3��nc�9�N�_�����[��Р�:��&O��Y�p"�_�?0�����j)��w=)����������_y�\*�v�voa���g_Hչ�x��Y�YD>ֺs���t������㞶u�S����]?b�C��O��`��Vb�Y�'[9�b�V�����2������7���լ����:n��_C�8�R��),�k�Y�&u�t���B�[���'وߗp����н�<�O=]�[��G��Q\�gn.*v˾��u'�i�C;G�������ǿ���w�3�U��e�؍��$�~U�'�p�:�uu�����Qޓ�2����������v!��ʤt��^��|C{��ȶ��]�f����c���v2��k+e������s[��'�?f��~)F3Ͽf�X���h��ϟ�>���)'u�����7�c<���g�wn��:e~����m5#T_3j3�/3���}͖+���Q0x����ΣE�\>��J;
]*):СN�e;���3Ӿ����ܖgN�ۜ�t�Ϫ���.��=9^���oN���p���Ct�}Ǹ^��h�t��{J%��y�m��KYrԗ��3�;�XN��Xk5��|ɢ���\kڄ��u{z��+�����.ܴ`��q�:����|g���'�5|�̨kAՑ�)>H|aL�y7��$�}6�74HEF�.|��r�R� H������^
+~�pիcr�w#ܸd��K�(��w��!.sI���p��̼�{���ݸ�S������g��I����=��ͅk���
�1�L�oC�ӑf���~�ф�D��a�&<���,�E�I���L��j�ѹ�$~�=�>��7�~�s11��	����޾��͋F�V��\���g�ۛ��S����DO��.{�}�2�F}->*^w5��m}]����Y��o����K��.�N�gL�Gl�o��r��4N�w>$TB�c1�
�X���VU�9��K�n�.���ճ���2��m�~��l�l�D�.�2;�v�#�[ӓ��[�0����&�7b�v���Z~���'���[��z��z�&�=[�S�[��[�1���s�#o��c��>l��w�k��]u�n�6N���s�܎�9u��ӳI:�5�%�è�[Ǒ�`cI�#I�qF�=��0�g6av������g:u���ٛ&����WN�M�[��מ=�|N!QşY���������Ǽ'��$�y�(��{	].�l�����غi'rڈX�aÓ�H5^Ӫ�cŸ<a�ZNs�#5��Jw3�b7l�I�����#Tf/{-�q�Ŋ��&|f{��ߎ�V����Ñ�{�	�-���΍���ok�r��b�J���t�'�fDop�_uf8���Hކ���Y�s�p�/�s�ufI#_]�	���Y{���a̺�5�Na��4�Q!�$����vZ�W��a�f��+2��t�!ɆG��!{��{��W'�.�b3ݜ0�W�>�\'�b8��9�(?)����{�z��Sai�v|���*�Q�`Y�2Ά
I�}�\�6��ace{���[e� 7,��5��A���J��os�����w�	�c��n'>w�w��֙7����N=��ݘ���3�:��ow/ۣ��:W|Q%����Gϧ_{�z��k�;׬�-0���N�����Oe�z�R�Qa{-l�h�z���}խ�w�F�t㾇�ȊҎ��1۟��c��7��q,��*3g���{$�v�+#bo{��ƫ�ڄf'�]��u{\z2"]�7wh9Y}�V��ݙ����t��/����6�Gwf�_�D�}|����S}�VK�~ͯA��^v�O����˻����N���5����sQ���J��;��w�����3^ܽ��v<�G�������>��FX�c�^k�z�i�l�㕼o�޷�Lw�e�Vo}ˏ]E�;�g�غ�/���z�v�5�ne*�[)���8�r��^U��˕�z��h�a��l��ie����=>~g�=�s�0Үh�?��+��Լ�%���\0b�T�V"�ئ�z�~Λ&[�Ĳ�0�9|������G��s<A�e'�n��ω�������u�;=�;{��Ζ|]�_:^fD��^�;�~�u��X=��.�]-�[%��/l�����s�OEOӵ�9�=�e�Z�F��V�ss��C�Hc�=��ڝ��l�����T�w�����+k�}��(�7�K{l��c�e��9ijV�T��G��&|V�ެ���b�jJ>Pf�a{NW[���7�"�~��h�k�Ț�n%�N�628�5u�ڟ�L��,|��̆���~�l�ه���wz�{d�)3������י��"6��s9|��d�r���IL_;���ihoOz�
�9Ӈ�6SM��Oֈ�`����dj����w�;�Z���]�^*�S�MŌD���G.V�eWiKs�d�S�s8Q��������&^��<����.=��s�gb�16�K�<���0���cŶ�s�6 R8:�
>�^�44�'/]���2g՝�?-��K��5c���.N�O{�>�̊���<s�`9=`����:S��BZЉt�z�B"ߏ��t�g�B��]g�)�ҏTG�c邊�j��hU۞'n?3J=�3Ik�W�qN�
��{����z�`���淥�{��d�h=ٗl;\C��}�k�`�F��-|T�I��ra�p�q���
}�d3�wp(Z铯{q{-�]f�:��q�L:�����{�.�=7��r=��<��/L���{��v���3���ݯ>鄅��~��[s�˺L�o���]UK]�t���s�m�[��{��*;������wL=N��f��hR77�[�||􈲥�w���w�d�]��[�v^s-�W����l�r�A�m3l�X|fu�i���NU$NT�Ѯ�vr'_\�{>���"d�%N�����=�k��;���n{J��3ۦDǲ��Z�D�d�n\�w*��)�z��m������b������+c�B���	�+~�B�̠�RE���&�Ϫaߛ�cy��<�:�O�N���U�{����/PFg�]£G]/uk�{㎘F�\�'[ޢ��1����Vw^6�f���u�=`Sw��~#�����T����S}�����EC�vt����<�Ks�r�p�u�� ����fZ;.L]�{��Wo�����rbK��{��� �$�Z�M`zw�{W1�P�?y~)���#��n"r'|W��K��WO�b����k�;��!����Ϗ��naa�_���&&�5�v}O�'�~|_�|�o�i=���c������A�� F���/O��s���o�:���雿u�^��Ԯ�`�~���}��ӣۇ�.�p�kS-<�81�{Z`._Uq
d5�m�Z���l�F�5v����3�ˍ1X�]���k3�e�aJ�6��7Y}�6���-6Ԏ�bJB۠a���I����&��5q�
�Q@�1C3�Qh�����_[C���ץ��� �cp��y���U �
��(� 1��h4W�3ý���<4G_�����������熬X�5���$I(�HYeڒ�)��s�\+���wO؃>�p��9��PH2dM�Ӊ$ |.$
�2��Q32<�-z�v	�s0�1����b �ƞ7���6��
�RXLF\�U����{��J�hX�RI��2G !�x�QG�Y:S���sm�JH�]��aⲉB4�i���}^�p�2{3L��z�~�c��W5ͺ���b �]�7Vs��AZIŎ��L-q��!���P�{���:\LQ��^ٺE�Xx]�<�)�B�) EfH��n�/\1��A�[A�xͰ����:�F ��㈾0Y��
'P����N���sL�gc.�{�L�,_#h¤l%��2I���U٦��O����-Yv%cb���j
cĄ2$��d��J�kǯJ���l։0�rQM]i� �k4�a�����]�F�S&[lޗGK�'ݝ�LzޝSX���҉l�In��A�3��c�V:j-��ŝ/1o��:\���)�C�p�JǴՖ�a�٭���e=A�?Fۅw�f�H��F�^�����*�E�I`H�ԏ��U���;1xɡ��h�Z��j7�smèR���6Z��%%�4�`�W��	
!�JZ�+Ig������j�b_X�]��4b�F��=r�Jț,��Ch�uY0F}ojZ���Ʒ�v��)-���zX�[J���.@H�� �9�B��}&����qD��*��ʑK��\"p�dH�E:]�*$�@�x�P�YU{#����b��]�f�&w��Q��*��BJ%0�DQ�9[I�َ&V���6J��'MRb�%��VZ-�E�;d����au��`���>�C.CK�5�@�y�&�T��B։�/0�����m��N�DK���HxYMr4��G}f��.�#B�O�W����z��B�68k$��k����C���OҵJ2�ك����hK pZa��%4�f5��/�}zη����O��:C�y�T$�����0�`���x�˷��.�z���qn������w���y{i�6��}���}��3�_�������YUW[V�XUUŕU�^*�Ux��V����z��*�.����*��^+*��*��*��*����~�� }�����[[ݥW��VUuUU�u�UmZUVեUn����[VUU�UUTUUŕ�*�U�U�ZU[XUUX^|�|����Uo5�UmZUx��V�V�UuUUU��U[���[V�^*�U�U��U]EUmZU^��U�ڷ�i���o�`�"f �B��i}��}���<*��ʪ��*�Ux�J�jʪ�����
��]�ڮ���U��W�����������
�ڴ��U��ۛ6ԭh��V�[jmM�����O/?[{1�6h��*T~�������������{���v{��0�h�&�D�4��:'
4I8iG	 M B��8P��Ȅ�M,�$�4M8&��Q�X�&,K:H�D��A$�( AJ,D�4D�8@�$	"IP�p8p�
8 �	d	"H�"""jF�$ �(B���tD��M4M4L:&�(LD��0�D�L�tN�"@��: �&"igN �$��XR^<���^yWL;lg/ߘ���9��?��OIen�*L��0�Qh����i�
��$b���7��np�;	�se��/4If���jla�D�j	$q��3��JQ�"N9m�/&6��B�Xp�.�ʖZ��l�2��3���y��X�Z�_����A�L�A��P�[�K�4��Z�z��BY��C�u�۞���X3��ƭΖ��C��^��j��jh�a��7���x�G��*���>EUa�ܭ\��4aphCF����E�p��Tj!$#m$"�g@�
��R�Z\��3i�Hd${:y0�<��䈒2� �qH�i9`���a4T=q.B��iu֛�M�U���	\m�5�hM�,��l���c�l�R���k~.�^Ld)�:�mJ��l(�T\n�W�ijʸ�6���4+���]�[[�2�eB�$Q�a���;��V�-lȭ ��6�2�ZΙ�`��k�߷|�9�n�n��������s�߮l!�����9�s��̈́www|�9�s����(�4��<i�"i��b%	F�t�0xG�O�^m�h��I5=���5*�a��3 ���l�/nm�0�	��C�W8��($���<��]�KQ�ғ��Y�cƝ��Bo��f���
�?�D3���г�I��_�Pߢ�>�RsA��ݥ��&r��:*~<��uJ�-���䇢o!�C�֊��������&S��Mf�@�Xa�V���tn��}ό�a'b#<�90���ԥ���[�>4M0�:"P�i�M�왑&T��k3`0O�G$�d=�u��^Oоǎv��?p@�Oڥ���&��R�=vB��2��5��x�2(����K]�@�?B�4�pY�d�=���@�$`��Lm�*��]�b��|I�N�,S�D�f���=�'%�aHZ���.��2�1z%���i�J,��0�4M0�:"P�i�M<8x�M~�j]j̮�^�4�-&pN�AxR<�K���e��G�s�p���4��(>]eL��Y�xf֭�B���M40Ĝ�XSM&;(4�)K����ӱP�lR������YJd�Tǆ�f�.�<C�ba�8`rB$�o~���_G�t�,M0D�4���a�u�^m��[���
ȝ&����(����5�~C`ܼ?i��c�[Qպ��MÐ���SA��B�|�܄�*����R��6�d2����̗&�Zצ�̛�%���o�vd5�4�ؓ�N"Ti�F^Qjy痽��C�7���a�"&�X�(J4Ӧ���'Q���KO�(�-v0AH��zܐ>μ�{hȐ�:�[,㇑�a��`�S�LJE�mdΦK�BjX˥!�nini|օ���b��G��t޵㈓еk��5
!���f�[-�\3Z�ˋ78zG�����d~=A���K#o��$�����cF�6$�V�E4~�g�,I�A�y�,�.���.��)��`DW��L���&�cq�j��+zH�h ��(����I�Iw�˚lS1DEz0`�%92d�T�-���P]I��0�f��?�M0�(J4Ӧ�b]���{�F$R$���Sd0�OBs�D�=���>s'�����}�vf\p������9#���-��ݞ%���5ɣ�CS�:i�x��a���䀴"e$h0���
<(�y@�`g�.�|Xd6{�r�<0�<$G�w
5���9)��=ۓ�)��m��4����%	F�t�,Ng�(�j!.x��0 �E0r��S!��-��SG�@I��Ҙ�'�*y�VC�8����f9�oG��rQ�d7�sr~C�8^Z�-�����)���!0^���?�İ��vD��MA53I(��	,h��$���Bg�Ӷq8�Qz�y�LᤵZ�[���xD�����M:h�',�~�+t�m6I~��h����,����(t�|k1���H���1�r��c�ʔ��d�<0=��߃���0��N��1�P������\Tjo�u9�үP��+��=�p�.t�nl�(�C�o P-�L��r��m�uמy�'J�4�X��ABS$�syS
�y������e22�F1�4ĕJ5�燌���k+qH��4���22fNTT-�TM4��e���P]����ȡ��-b��mGcTҵ����~�a n9����j�S	����O����.�ѓ�0�W�m:a;?3;��d5;C�a���KO ѣ��3�{�Fi?_�*����d���8�)��q*�cm5O�<4O)�L�,T�b0�U�i��u�4ÂpD�(�N�%��Æ��N�Es���82~T�C<y��Y."��e��u�k�TN%�h��2D9����3�y��8�.Qٙe0�.���D�&�`eh.M��	 ��J��N��i�l����v��a�RL&�i�G^LK,1��]�aN�� �[]��>Z�<|��WO�%4J�D��	;��,�LG��ʹ����ӧ���)6�M�Sű��Ŵ��V�N֫uV��o)�Ħ���[�����ʷU���WV�S��o6��ZU�^&�kR�n-�L�XaV�jl�M���m*��&v��ڭ�i�r���ZUi�*��m2�YL�)e4�NV�M�ͪԯ0�Zk�*ة�aj�g������|_�2�������ʭ--Z[��mV��f�o+�U��O�i�m�X�ij�m>M��Ui�m�X��|�:�m]K���lRm6�ax�W[ꭗq<R�oT�[M�Z��}�}Ҕᇦ�SE)�DOJZ>��OK����7K�ε�϶uS�k��9:,|'�ޫ�c�T�=Y~�(i����n<�aD!�F��_!�ν{�J#�寁F� ��A$���`�%�10"���$�!D��b�(�F�����I�K�l�%t��p��o�3c�����uJI@�[<B&גdɛ	�$F�$^}b}m�b�y���K�s���� |���z�rf}��;�g�ʺ��d>!��?�3wwwߣ=�{���33ww�;�{�������۵B�����9�r�h�4���Z����<��-���ͼ���Z�y2�b��D��D�j���!"t�����?""����3c��v�M�V�IӶpΓt�I���m��!�g ��`�0DD����j y�}�� {!�`��z��44�h�����m�Xc1�aqD�
����ٛ<��JR�H2C�����Da'l�d��Г�����k�4���DD�ؐ���'�	�������	��i!`����X��	�st8���a>��lЌ!Ԟ��Ɛ�Ѳ���?��fZ��(�H q�MBF��Q����G�N��Sͭ�|���aka�󭺳���{�o�V������I>Ї��R�M�Y"I"�I�{��@�H�����$d�DO~7g���T��aw��!�� b�� s/&ffɢ��C�[ r	?F�y$�,�*!P�iA�M�1'cҙTCI��v��,=ld��9,��pM�C�[�
h�P6$�a�<%&���}	�&�'��i�O�#NA$�i���!I������`+N'��BP���B��������aؔO�N	�D@�Ύ����3��Q�_L#r�a�JM����<�έŭ�-�����6��b�SS��D%�Q�a��1k#��S-q��8�%e5Y15e6�bØ�S����i��(�i;	���T�`���2��㘛��ʋ\1�� w���BWCKVm�rji�m�t�ɫ�q�.��&f�f���=<,����2�ZI?��@)���~;	?L4{�h�5C��v'��DD�!�� Ұdf���҈��"�=F�0��D�dQI�Æ�# �i�d� ���kkE��C�O�"{ �a�{�=�L"ɣ�� ���t���BQ��F��l�`�I�V��i��ddt�'���<���ۢoBۮ����M�$��=�K-�����6%hO~��o\���	����u�_(��"XC`&�$l��'���u��ip�Z:�m�<�ozf�al�l6�^y���o���Tbgz���{����O���F�r�����$�M��a��L�z!�2"#_65016�؞Y�'`��d�v��n�<ۘ��`���SZ��'�2~�]�K ��~���e?W�d�>Tc�覤D��%��&�)L4�Ϙ���bJr�Q\��C�b�DD��ύ�Ժ͚B�
&�	�0pƂ�6U`��>k�O�Y�D�d��!�d8~pЌ�A@XQ60܉�%7o�\W�N"
ZtDOd@��Z�|4 s��LB��Hn0DI1�"�FI� L"�VU	I����D2m�ϟ>yo�m�R����+e�ym��zSx��3c��*��"{���RQ��}[��x2�с�&��Pm��"'&�C�Ĝ5d�|��D7r\�!�O%)�r�{R���ܒ��)z:!�&�,�?=��W'�<6�`�O̐dL��"F"'���նئc���pYtOu�l�!�ȦO�޶���S�'�'�$�0�(���Q7���?M!�!�����1��C	a�X2~��
l�,2&�g���DL��������$`x��2J�Ad=<|k^�PDFC��D��ODdSRbf&a���S����?-o��[y���l-l2�^y���yUB��s9k��]2bb,����"� :m�*�"0㐲T��7�C_�d9���tD@�af�O �hCέ��C���bz!�ܙ'�"~4�鎜s2���Z8�֒�l�C�'�
B)����Y!D$��7?{�}�-�R�KGP� �0��3�R>��$�^�-1���+߇	�>+�?C��x2��Ne��\]C`$S�3i:&����6PX蘁."�DK�k��D@d�=3$�� �l��	7���bO�? �&�Y��P�O߹�sPm����)���R'�6LA��ZNuEV%�"A����!���B�IL��ϝq��|�o6���-l2�^y���j��W��Y�2�3Z,FAή�6jӀ��P��T��2Щab�eU�3#$���)B�|�2��"P�G���2��˕7`�b!�I��+.���-�̹�qJ�vlc�[Hݕ���ɡ&�;8��!��*�[�Z�X��s3Dt�6�"���P2|�4'Re('�D�X�Te �=�XM�=�y���W5��ǂΨ�~F���8�-(j	?��9�m3@}�dD�2n쇡w,u�\m�;��&1Г�g>�ng�b)�X$�KVH����ziِ�j�J!�P<����$5�%O�%�ђx&$�K�RH�n	xR��yۄ�"���c�3�o˾� ���+�|�Mf�����ŀ,��O�ZRla1��&�hC�d�CPgD�12��"���)�j2ٶ�e��-��^ZԵ���y��[s?'_kK�MW\|UTC��ZU�1{�2,���O�"ȧ�I=�=;J2M��5�!��[ ����-$�E�̔����ÿ���������ġ��&'D������hy���$`X_p�M��Z�4���)OU)�Ѩe09�)bPO�d�������cj�e�.���]aZl�ۀ�5'S�C�Si�&�6p��:��n$�Y�'�lA��-�/��!��3e!S�>���>��6 � {��"�̶�N%����0bZJ�#E���[�u��<�jZ�el��o=8R�Ԣ/�U3�UD�ɝZ'�;�d�!xΫ_�}6h=H~K	^�T�x�e3�&&S,%	A �{��Hv2X-�$��(���D`bC�CZ��D���5��sB"!���
�b��.:�\��
)��q�O>��O���JQ6��=)DLm@�4�0|$j%���%��&��(Ob_�m��h0�ܖ���αp5�I�8Zh3�[�`���feύ�ޔ'�&*�D�y��[�u��<��k`�٣�Ç��NpJ�r�r�jf�d֯��f���`��p���!�$�S��
zl�h�> �7��	�e �i�4䘙�DS-���{O�9���-��Q��3r9���8w�蜂�����0����,Ei��/��3�'0�$�
P)�a�����HSÓ$��LA&�!翚�Ô����a��2w	�	�d>�v�ga���)�'!����l� ñ����F��Ƙ���*�u��Kyx�-�-�<�y]N���iK���6Ҳ�S*�*�I��6Z���Ɠm*֭�VꖟS�y6�i�v�yL-^M��uKm�-�[��t���0�-YR�j��kU�^qV���)u9%VM���Ų�-�Z�%��kU��T�VZ�J�酣�{TMЦ�����)��7SJ�KU�[aKN�eV��^&�i��۬[
S�|O��?+�:�����?6�g�-n����W��qV�-]M�4�en1��^]Ojv�Ofg�VV����}���O��J~OϪp��N���ֱ3n/�:���wU��҉�N=*av8zQB��O���_�OP���_�R��%�$˘�;���y���#J8�1���<n�IRل�Ȳ�ӀnQ�&���ǐ��ݵr�Ch�DQZ�J�_b�=P�o���o�m:H��Z��YT�o�c�j�F�z��j��F���H,$�XI�$��"�!F���L2)<�^�KW���m@�]��#F��(�G���^���{Hi�C��K�4/��ȑ�g�Pg.kch1����fA�V�j�͑��!��c�G��&���i-�	�М"�P�i��A��ы%n�4���1�T�$BDd��OIU:��D�cP������'��V^�ʭjx5'X�'��`�b���
,�3�6w'{�a`�D�-���r^|z����ѽ�ܣ!H�˲H������iPI ���dj���$���\�w,
����D*R\��!!��	,,�X���A�eH[XQ72֩��xd.1���L&p4<���5fj���$�m�:&$!��ȸ�7%�]�ʠ�&��ѽ7���kH&�XI���%��XQ4�jV�i���+0��-	e�#m�� �"
&qD�Ҥ� �_������ U��{�����_�{��=�{ww33�U��www=�U}�����|pD�0DM,肵�kam2�ͼ�c;�VqQDʳP.��S�MX4c�"<d�(#&Ʊ)5Ocyc��7��P�Z�
SZ�/���ַVз�[vL��y�]�l֓X�bp ��gJ�12H����@4h�
(� ���4)>����R��hԴ��·gM7
t4&aϕ��Ѱ��*\��L|����z���z�lPP�}��k�a����������a!�Ůe,F���[�B7(��n%�&��9�S!SA���W�t�Z2.e�1�J:��J�m~}��̦\a%f��=)��C���e��|�ϝm��-jZ�[L��o���>0Z����$�I
? �ʇ���f�9L���ME7O4T0Z�2���_>f!�T.)Ox�q���2�嚇��g���3�cIp��X��exm���̨����~�L�P���]Fdت��Cߔ�k����s�����:�6����)��_!���}]�1)�6	UX&��`�Y�L���S<ۏ�:�O|�-l-�^y���rL�S0��"�2VE#��ZUTCㅘj3��}L"ܦT�eJ�%�u.6��� �$�����5?tSS8R��)֩���MJ��x�L�"`�Kt0K�$�d2AN��!�y5�X"P�	�;N�[�a��m�K�`�y3�L�Y���U�h��}9��0��Mvg�L:Im�a�?6r{߿\��q�$�8rl��N�TT4�k|��y��x�֥�����6��q��p�>���Z��32��;��R�!��!�Roblc���<ڀ�&�e@J�:0�!�gt|'�f����;��Z��&c�8�Gb�쓹�b�t�A�7=>|-:r�=~�pj��s���~��IG/j}Na�0Cg�{��C<&�p��!?0��q��#p�^h�clCJm����ϟ-�ϝm��-jZ�[L��'�����;D�(�J��"C��`���n��ݳ&'5m\%E Ke_<�^aP�KU�WR�m���L�4�e��7�F#	�\�l&�*��lm�,�F�0+���Kl%Di�I$�@p�Fa��Hmr�& �jd,��p5 LB	�?�l�0K�[N~��3SN���	�G!L������fj��ޜ1S�z����RPG��a%���>����������hD�����kF�qn�4a�{M߁e��r!�~}L5��fǥ0C��w3�Im����0k)����ן�ԙ}]�bfzb5
(���e�|��sU�`�ì�:��|��ζ�ǖ�-l-�^y��㘹�78��0�L��6����5�&A< }L��~0�|W�-��є��H��%�����5(w�NC��Ϯd�nN�Ҙk���a���Е�!�h�p�7>�����+�iѥŞ�B�0Ї��Xh>�뿵u��^I	�A�p�F��r7y��2�Ql�N'	��13�\&�0�&m�4m)5��'l�TL��Z;M��y�ϟ:����O(�ӂ%���M�}55��UQqX�a�p����o��8��`'�)��}j�(w�Da�g�m/�E�~��J	=�����F�oС��V����������)c�|\�H�:՗���rO��'
`~խm�w��9�9����t`R���8��k���sK�f(ɟ|�|���+:�JSe�������7!)�D�Bf�`N��N�3�L����n�u��<��kam2�ͼ�Z�*Q�TzY�1,U��2�ܪ�Ҫ��z%����L��a��I�\0w)��p��~�~"}愈�3e��_dS�_�a�VƼ�&�uU,T-�})���c,0����a����~.Y����>�xldB�>���&�u0�����a�� ���g ���	A>����f�p!�>��!�t�rL�;��l�m�|��_:�Oy򖳇�:"X�4�	����ʩ���VrY���	U
�#:�iҨ0�9�#�"�T�dn�ͱl��fIo��x������E&�i�H��,�Bk���4֔�[k���� �\B,�f��m� $�Y����aeY�D�A�[��Z�����8`Y������Rcs�UQ�P��亏:��bz'QOJP�x
,�ٮ���B�O����0؃�|&�u0������)a�w�a��l; u��"2��<ɇ�Lz[\~>����A8+�d��W!�]獽��0�N���ѿg������Ӂ��L�d@��"w���2Th�l�2�g�KI�
u��:믝m��<�K[+a��lx}�ML�_Eo�U�9"�)F�"��D(��g���`�!$�D��}�!�nb܆M�3,�:ʍ���Ǿ���v}��O},�`R��MQ�oG�=>J�>��v5�x���a�4�6��I�����ܵB%l(�a,pڎ�����j{��ߌ���ٯ~�ۖ��m�p��n�����	d�D�a�?[P���'C��}}H���h�+�W'O��O�$��וo+��v���M)m�Ͳ��YOe�-RM���V�Z�3�&�[�6�>]L���m/-*�y6��+W�i���ۊ��c�W��j�*}Sj���l^�m�M�]mV�eX-��&֚�U��-��mV�`��ڭ=NSe��[M-R���FI�e�%9%iJ�jU�S�16�R�­�ZV�ix�[�Z�>�/����_�>/����j�>5񺟖ź�n�m�yk��x�*���jujS����ٜ��S�S+WV_�=3�k��v{X�{W����|^�}��}3������4Ħɴ�J�p�0�4����iKai)�������M}��v��7��s�3��@`��OC���;n�f����)��⸝�jD��2. �=H�H�s�3R��Uq$�Q~Bw:�sCXR]"w�ҏ��8��{h֍(���O�q���@Pnvx��w�\����!�ȡQ
.S����;k��9٫w�zp�&�r�g2p<����׮�~�n����UW=������Usۻ���zU�n����!g�xO[���疥�����6�׹���O�O61E������~7d��gt��4�oO4օy��dK�0�A����d�������Ѷ|VB(�f+D��]��L�c�o(�KM�m���..����1�hk
0����m��'-�h���å�m�N�2��)�i��ks<���^��v��5\M��]y�믛i��>R���io6��êW#��%X��������j[��D0<?	�0���|iȗT[��0�\Z(VV����>�h�b~L�Ѱ�-?@��l��P��<�e�4�|��C.����^Q��uK��I�P����F�}7>����2S�C�Zl�w&��:O��_,g9�g*aF�N��q��݈�6��ۭ�[κ���<�Ե��[���P;z@o��X�IRV68$$Z���anb�2��'JEy��s�kE�!��QE�l���ԮU㨚td	���+���:���A!����Ԉ��1�*6#��5l�Bxl-8�%����t���I ���)�He�[q͜�O�nM�{�����26���f	��"�Ss�ðcδ�I%���MS�;�GT|�jfg>�p�\L��z�E��8wԙ���m��y�s�=T�3;����ѷ�~:h�å�N�Ml�(s����2f��c[t���Y�4�U���l�/&�.�r��ݖ����@����N>|�6�ǞZ��V�Ky��ӧ_.���������j�k�9`�3PǦes�I�-��3��O�8{��ō���d�O��2�n7=:�}&�wI�-��!�d_��rp3b��؛g�R>����]�v��jV-��ķ4���USge8x�Ҕ3�ӧ�%1������?pa�N*"~��~=9�XyN	���m�û?�4�Zi�V�]|�OyjZ�Y�><>BP�8�1>&�`���&ffe'�0�S��'�3JO�I���a��4����q7�SJZ]cr�����*a��I���D��|K	�O2eh٦BP\{6���4D�ӝ밦aN�-wI�0�ҕZ�T����EM�A���0},���*����5gs	4�~�����CD�'f��2Ɗ|'O�u󮺶�x��Z���[O6��T��v����ʪ�>��N��Uߩ�Z0�S��;6d�l�M(�� �j- !%��Id"�u���-M�O�}8~A�Y�JS4�3�18���!�K[�I�h��>8vh?�x8�Ũl>;U<����Օ�N��CF>���86�J���y<6l��t��ّ��/�'��ai|�<�u�ʹ���kel-��ynܧ���bj�⼫��QYd	��P���p��L��M�U�H�+5��H6Hk,..�����-s3fs.��c3�[n�Y�mGٻFٰB�VXK����� H�Hs=�e3�ѮuYn&6�{?'�A<�XkB�@�<�7�_�eʳ[8	=:a�Ozh�e����:lL�r|h��	B�*d0�_NCBŏ��6rO	����Jd��KӺ�ORX'Ӈa�¥C���֞X�����ZTb>�9���&m��]lYa	�~E/+v�m���Ne2�wT������4�[���V�Oy/-l���xp��ޘ=�EDQiJ��b�ѭ(ۛ�Uu��˖{�UD�����xv:���OND�v�g�6�&z�L3P�JP����g�߆���A����05����)k1�t&&���Ո������m�x
\ ͟X�8�fʙ:�TJ��7��`/�2Jy�����B��l�u:n��V��-���um����������fzW��e_�9¹}�Q=������y'd�a�)ovai�Ў:[!L��������Ȋ0��P�J=�Kto��?0m�Z�(e��f��Ҥ��O�����,�mE��.�Z�u�Ӕ�^�m(t:d���揼CYLMj�)�!��|�L�0����T�|q�u��N�f�,�&���ف���D�#,ĩșf�~�y��[��[�]~i��%��l����o-�wQ�V�8�� ����
i��T��I$����G!���˓�O�×�j~?�K�4_*���-e���-��ِ�d=0�$�0����N'09/�d�v�ޟe��<?L��?CG0���yإVO���d��C~^��y����T�i�*'����3�o�zf�#?2㸙�;[�q�Γ��|�]��Z|�L���r���q�&�T[*�՗�U��Se��-V��s6�]N�ǜU�]M����y1i����1o*ܩ�u+q\[�[��t���*�e�i���6�Zxҭ6ʰ^S�M��M&֬�V�ش��kU��&�[2�Jդ�ՃOL2��=)����ZQ�'���ԥ��y�L�*�
�i���x�OK��z_Ok��ҧ����>�����>c����3n�֮<�&�i���۵3ի�6��6���;3�[�������~��X��:Z;C��_I�Ui��s<yl��Zm>OWo��/�Տ�|R�p~0K��i�$����%���x\@�9�6z�"%붺qBͿ.�0��*6��h���R������$VS�ѝ#CMƮ,Xn֍�Sx��h��uӊ�Ha��,'l�EK]���-���]r�cf@Z�e>Ok����)ۗ��+R��3P��h�N&�d6�P-y����=�4�C&6S�es�T�!8t�L2<��x阡�(i��	8R1�4�U2��		N�^�o��a��U�mĪř0���+�4ŭ���s2$��'��(�Z]J	�Zk�6YB�q��q��H˴9��)֌�D�0�eV�qLp�hH5�]�1�<!�Ht�.I���X��ѧjҁ�׈+�.���Nf�s���:Ă��[���$P�D���{n%��B���I&�[-I��am�e�ȱ\a��"9���:K��bd宜��(��LQ N��;�18Bp7B�|��em,.�����Met�۩��-B�����0aPDטdiP%��0��$ۇ���y�dd��$�ob�-͡D����ޞH,&CMP��0�(K<E����CM�f�$�@���8TGK���}�{=^���^��G|X�(�Z��&�fk��n�g�������2�$V]�TH�#��Ą6P�W 씂�SKS-&��%URF�\&&�q�{!�dq��s�����z<��������G�Wsۻ����ʫ�����p��V�u�]y��<�^Z�[+y����=ߓq�k��AD9���-m��]jy�q�����l�+A���L�V0�0�TJ�:-���a����(XB��[�)��3��)X������zPd�a�4Jƌ�I$�@�8��J0��-�#E��i�GF��?��sggʖA7
N�q�����D��ǇM������PQWSA�����)�A>4j��y��ܦ��4r]�53���M�Yh�L&R�]����V�31�R�p�.oMx�$�'?����΋of�a����ߑL<�TM�MϏ�r>��MD��Fb;��Kmo>u�ŝD�<x�㇄���왜��wY�v�qu�UD)��Zd�&s�K0�6��ɔ��es?��>ɪe�Ś'�JX~�����7a>��Y�V�>J�`(
)~0��<�(y�i�D���cm)Z��%����Z���5�=� ��0�L�1p��8�q�p�(�ne�î52% O��m��N/��F��V�][m:y伵��V�m��猯/�ۧ<���⪢6��!��J�+[���O��0?L9pM�����ЇK$�����~6p���08�(`;���U1�����Lr�s2xl�٨z~<2N��)�~��\s�"r%}NN�:p�u��5���e��PןCpD�Do˨������H�1�u��TҞ[�|믛i��%��el���yn���;-�N�p�n�3A}$�H >LI�S��Ɲmg�-&c.���t=��i�0�E�0���)4$�qO9��7�`��" �{�ߩ:=���s���t�d,83IFb2�a�j/2�55,K��v"�l@�Vj�;�j('��0?D���@�Ǵ̦_b���-e���+@���L0Җ�o�:�ʹ���ϙ[+y��[�3;��m���q&�%��d�*�)~�b�kP�uR�M��6�oH�b.�;Q<6��$B�H��Eit�́;o[^���T#��/�q��Y�LN�k����&���� ��D���ap�.�uӆ	>$�H 1��m�$c-���jj�!�Q�\������?O�aa������ ��2i������8�������n	��)���У=�Z�4�x�d��!�|L�����9i�>�Ѡ`P��z&�0���ƯɈ�)��;i���,�T�ƞ�X���^�_�W�_�$����P��S/a���Q(�9{PDd���^�M%5|Ucb���o)���n����<�^y�+eo4��v���LnmUQ
zd2�>��6�a�o����N�t���kG�0F{�{�́�~�#S�I��¼�Z댮�8�Kµϓ1�c�3�I%��<����2�Mj75Y���� ��F�bim��#d��!M�p=W�0�4	�|�������r�j#�k�N8�'�������j����7�����8���i����$��8xN�'��NU�8�PQE1�f�UQ'�{�wP�f�NB�f�D>5��>W%��C���%NC\4zU�L:hם����=��m��o��S�a[�u�f�76v'g����ɇ���YL2��I5�vn(n(�tL=,�~��;�~�f��R��nM~C�]�t�D憙<��iK�9���h4�!�����f�D����0�4�,頉'�8xN�+v��R1Uə��J8�O��O�u'�b���7?%w�}qJ�L�93Xb'?uf�ӧ�=/��f���y�4��ֲ�k���J�p�Z^ViEC�	����!�s)m�Jg��Ҡ�/�є���s,B�}vIhq�Ɋ���i�>��JI�ф�yF�L�jyj[����gMH(�x��,K;��"��x���C�����W���U#dS5��r:���e��
	"������b8"ی�6(2͍��R�8��j�b���Yn�u���	���}3���$�A�3B��ʜ\M�$P.���Pn�b
Xrr	'=����S�z�up�0[���%C��	��Wi>���7K0��:v"�7�仗���-�-��E:0DC�}C�~��f`ښz�N�s1�Zn))1,�δ�L�]�e�d�*1&��속H���)v~��j��dw��:v6��vԬ8|n0Ó���&�?%��bLaR��mm��]un�K:h"@�G�<%�d�v$���k�d}�RyR��� #E.�as&��y�UD?'e�>�"r���[C��?x}� �}�ʧ�Ӳa�l�p飄M�>�(h9<��p϶uﶔ�տ���Rz"x~fqe��Jm�WJ;�aq����)�|���)FaL6?�
h,))L0I����QL�EJT��q�Xq�|��%����-�6��S�<�O<�h�&tK,�:%%QD� �$	�N'D��LD�MH��,LΉ�ag
舐"pK��$I AJ8h����� �pK�KǏ2ɖR�Oy/)�4J$�$DDK$DJ AZֵ-�������y�y��0�0L�LLD��$�pA�8��"l���i⍼�^R�a+E���������3��F��\W�Ue�{<����7+�v�ۥ�Y3:���:v�rZ�b3j���AZŧ��x�X �J�������v�{�[][�3O�	�u�rG��z�к|��lw0@��i�������<C:��(�.�-�kX��:�%GWA�!���gOɳ���{��s�}xی�X&"���sۻ����*������{ޟ*��������򫻞���}��Ox�Ɖ��gMIy��V�o6������I>�������4�xl�L��2nna��?�.��ӳ��3.l��B��T�߻�	���p1 ��X؊D�����Y��l+Y�xS��?B���4`�R��}-�*[�i�d�:�:�6|���`0�:��L7'�!��)އ�i��E<���&9|���vJ��D�#IL��4��|뤳��$�~<p�%�w�a�h,��I$=�A$��Ӈ�B-TQ�f:�u�}�%']L�L�1qABt1x߆��Ɂ��E��� nf��e�Jp�n��6n���#%4R�#�a�a�KO�b}�;��>w(���MsvpD�lK�Qm{F'�w�c�4n}�E(l�~�-�mÞ-%��C��I��)�m��uכi��%�Z�[ͼ�Eh/6(%D���P��h�2��!Q8���0�0��X�\A�D�2��Ԯ�$4#�	x�$�<�#A������S\�9ͫcu�iH�m�	n�$�H \x�qF�v��+pt�Ҵo�?	��(`�<�����wG,�4l>$K�0tm�H'>#�Y�8�3A���\=���B��3+1,%��֔Li��pѲ�"'D�?A�!��^C3�&�5|w��-�3��zR�C�M����)������\ֵ�ygK�=���Xu�\�v��5��)ʪ���>����!v�.[�!�Sɞ�-l2�6�^u�Y�DH(O<%��9��ǜ����y�UFa�i��)CG�e1ٙ�����Q�i�i�a���M�N'Xt>)�07;�h9#��3qP��f�I}1=����C ��0�6�Lk����D�)�eS5����>�zn��!�Ƨv�ԨyJK�B�̡�����[��fe5�p��=
F]�:��>qNi�4�,�B@�Bx��,N�=�-o�g��a1	ֳi̼�AM�i�مꪢ:&��xpÅ�.��ɣ��h�M����(`lN��N�����5#><FG�HP_4���l� ܈�	�%�ˈ��R���p^sn�{
}�S�>6{�hL<�e2��4=9䧧G�\�"���?|��F�n!���|���)���C��TF�a�T�>y։gM D�<p���I�69z(�8�0}⪢����~��e3���=�x�%��)��%ǔ�RKz�;Li������R�zd=��v�!��R�K}�1�Nu8�jܹ���FB7
�vn2�K�D`a���L��a��ٰ�������>����ì��kr��C�	���v���Q1.V�a�<�ξ|�6tMDJ��t��#�S3�k��^c%�HDʦB�@d�&�P�Ѷ"����$�M`�V�J�0<LϠE��覔	
k)���L��AjB�����e�c����� �(4#]p�U��$�H 0��"G�"\PH�'�8�������8�\7�qĶ�*"�ng��
h�Aյ9��	u%̊8{��6"i���{�3)�I�2|��S�nD8'?5��y%E6�7)�F�F"T�=��`]p�Ͷ��qP�)P��[�����!�I�N������/�S����<��^m��yO<�<p���I�L�&I�T�g����]��.����UU��f��G�f(�?�R���r�}�~��7G��K"N�aF��[vp���ɟ���a��%�z��3�??CE��'��LN��{�tSܸ�Y�+Yr� �����M���Z�$ݺ��aY�o!���=,����f�C�:�ч�:���xa���oD�p�d���L3��Ԛ`��-�u�:�ŝD�����&2��(��"r��j��!�ă�zaĹLS�D7g�ð����	�����;9#p=��Xh�Ji�)���?J&&K,t�MM�
���-�ַ3~zS>GL2������F��ae�)>9<���=O�-h��?�N�:,+�G^w�����p�����{g�4��m��~MΉ�H�Bx�����U&Z�Q��W��]����W&�ՔXST�3|UTCE��?>�$����#�m/�92�/�����W��.�Vs��׬��ك����~������������M��N�l9��1RNĨ�[�-�579?M�M��`��Ʒ��('��e�)����F��a��c�,�ϒ8nl��M�l�h`��"h&��YD�d��(�(�% ��&X�tN"`�&�h��u��N�$�bY�#�ig
���BtM8QbQ$�H�$�"a�D�0A$�$ A��8AHHD�IDDD�(D�A<x�G�<p��Ş<`�&�&�h�`�&	�tC�4���ΔrHA���,�4�:"Ao<���<������3,��:vGm|�z�.�y�>�����b-S��OS$��G��\����`��.y:A8 ��җ�[���uPN����jm"u�DRAMo�����_\�=[C3�9�&Yq�
�ݐx0�Mc�@��rđK}�W����J��&�[$a+6�
5�Ւ��5�$`9p�&���#Kl�<���2��@޷T �
����Ϸ))D0yC��H���p�`�2�ĸ�%�&-\R4(�D���]U��'������H�5�R��z`���V\�:D�3h±o��N��}��I���Igf ���p�%��8�f�]�Wִ2�U�U��ΙB�f�C�N�h�!@�Tn'��YEّa$3Q���wF��qbQ�<�/�UR�������Ӂ���c��Zd���A9L9�V0�v؍�oo��Vs���6.���{ު`�@��O���U~ �\�G� �t\�K��C\��f��|6��Ŭ-���]v�%���B�f9f�T���d�A��eLcHx�Ɯa)�(��qF0�U�C8Sp�7.����-֨ы|�t��3�ݚUAN�l�=���VG`ă�,� ��A8�r����QDT�ɛ,�m�-c-��M�cqa�І�g{���JĉB�)�֦�%H��!X�'ap��3!�N-<��"f�J�j^����{��*��������R������{��yWwsۻ�����<Q��<i�Y�4I(O<"4Q���xMH!	�`$�=�|�I����Up�lK1��������U�pS�ym����Y���k�D��S!��$B��EU��+l���I*D!�|2&Q�$R4��:�v��ú&q*JXt��p���\��LԣCp������y���S�"5y�g�eG�R:L�vz&���^�r��y�O��C�
�=�C�❖f'ʹ���fd������!�{L5|�8���*Qg�i2�um�ִk32b��F�Ɂ�`a����ލʰ�F���㬼��M�$M(����$3���L�+4�A�+UN*J�u�2^�uD�&R`�)id��fe�pRu����Xhن��}���ƴX�9�mhM�d��n'�S�U����I���&O��u���� ��5�	��)�K,"_D��{���}�l��|{%��c���H�������~�ƲE�3���iku�V�][�:�t������ٜUZ��Ϊ� ��ZxyN�sה������t��ݝ2TѠON�SC�^.�&��t�H����DvF��Ya�ᙘY��s
~)��'�
0��a�&`�}i�b���p�a�<\;:J}N������.�����No��'а�ɡ���31�&]m����&3�i�JV�m�l�����yמa�eo:������C���L�CnZm�x��ʫ����aJ'���/�P�:3�*}��`�I �99a�̺�Em�E��:h�ç����)Db~8s����j{������N�L�P��v�if\vS5ơ��0A���018/��K" �,�6'a)���e�#7K��D�aaK���a����Q2�;5�L-%�l��,0��eo��q�DJ4�NO^�������ə��)I�4䦻��x��Eצ������v�eӼ��B]|�Ȧ0�p�UȤP���-.�M�s!ͳu6�ZF$�k[�
	�J�4��ĒO#`�#nH�*�m֎`�ƻ ��?4����NCh|�X�:����ge>��U�!��=�`�)���ն��zdA�a)v�����'x�V1��IEd<�QE����<[M�DO���A;����!k%(B���$m�9�
T�ff�Z�2x0��<:a�)/#��z_�㱆�e�θ�?���	�%Q�<i���8]\���mR�~UX�����y��ܙ�)y��-I4��0�s5W����b���*""�6"\'��`��""3oFҁa�X"'&����A�Q=<U��>�]4�m���F8��2Ο�>�O�0>�2��癶p����(z"&�����h��D��؊)�S�>�.Ee��ۍ��^y�έǝy�a�][�q��r�r�n�1�Frk�*�DC�0֡�=Kn�	�<JZjz~)�ga�	�2a�	��N~����6p�т&�1�)��4|�rU��-�Ԡ��?#��.�=�DN)���>�*(!�g�(���C����Uw�B~����=�2�֙��ޙ�y�,%1م�	S�<o��gD�(����ϕ�>u���N-�KZ�un<��0~0�h�z~=;9�i[ڨ���CΪ�Da���@�|�~�[����h�Q�9J'�T���3q����������_N��Χ��e�j�0%�Lm�jK0�R�dp����Xk�Ҙ~c����p���d��;?Z�����8%�>0�JQN��"�L5�ɓL�������4���%=m=a
e�Dw�%�}�ɯ
c��Y�
<�*^�C�5g�S���SM��ZY<&�0M(ҍ8i�O?�W2h�m��I��"�H�Lu�29�[^ӏ�cL'h�If\�`�(�h�M㐲2�m�\fK�[V������u���h�;[���k�tL�M�	A&c���N�sv�,��}�Q�0��}�yQΔ߇��]�2	��V}����/�N�����|)Y�&6okM�D�KU�URRc+KId�)�=&R��w�-i5=9Zu^��<�v)D��\T��T�m����Is�)K��G>���:�J���,I-���m���#��R�D̝P���
^�o���Êqǜy����Y�h�F�i�OxäQئby����:�T4l;M�°� �e�{P�h��
��S5F�i�#$���wܷvZ�&��=�4%���:a�ѓF	��h���Nfb�'�J!�S���KcOK�5*f���u�3��Od���t����\N0��p�*$�)+�3�h��>��`�~���~��75a��ͭ�k-םy�y���%�X�0�:%%$�8@�$	"YB'	�K:&���"&��D�,�0�'M8P�A�""'l�8s�	E �@�%$&0K A�/))x��L��R���%� M BD�DN!�����[+Z�Z�y��S�M�0N�`�&�`�`�Y҄�,DN��Y�i&%�$��$�I|�X�'��9U{�q���w�_97rMO�R;��:sm�6=R���Y�Ӯ�c6�)X�2U���_��j��<�>�d^���`�Lx�&�\hy��zч�������J�TJVW��s�	��c��ô,H�{���]�t�E1�PĞ%�wp{����n��C>��L��T&{۹bX�U���؈��������{��yWwsۻ����qWwwۻ���{���n�㻾���,��N��i���(ӆ�4�I�U���?	��cMk����Y�����m)Jaq�&�J^R�Oq��9��c�Y����+,��Y�=<8a�(��ȝ��j��Z�q�´�V�6�h���y,Ç�CM'�g!�t�wx����`�M&	�aL83��m�=V��?t߫���-�=)y���DoI�j!��L�amv����<�)v��>S-���i���q�^y�X~4~=?�5+�������������6��O:��XX'�������?S��!�f�#��K��)��n'���kno�:��k�����+�F?���ӱ�KQ.��<�4��rrK	[4n�b.�q0D�{
{97+F��a,���";�f	MI䩔����<���5�T���D�m
c	�|�-Ƙq�_4���[�:��:ì��V�[�e��+)�LʗXdC�x���Sf`���^u�Vd�*���b!�jǌ�6�D\��dB��i���ˠ\��i)9F8��qC<I$��1��!�r҉e�CT�H$�6
�5E-n�Sge<������3r����jnXR��l�揶x}��)}P��L�w�>n1�R�SsO��۱���J[���9��)}vcΒ���	JYeP�M%����d��3����"0��=)���_	�y����=��x�Q����}Ea�'D��M<`�"1��D���}�%brI�g	Xbrr�UX�a�Z���țS�E<���C��l��N�D;����-m���	���?Ey��`���|���u3�R��!�|�e)J��8����b�K�4V��G�y+D3(��L���Z���--�S5��]6||a����)�h�+���������q�Yq����x�4D�J4᧍<a�Gq�mr�uUb!|�����\�|��5�n	'ᇦMOaD�,/JlK�p��<��
�G>^X�~�V��q��ȩ�:�3,1�᧘9C�*y+���o�������	퀡���7&	���������B~!��v�ju�a����)(�[a�_>[K<xM<`�"P�i�Ox�_��=M�˶��Ϊ�DO����?:&��VaM�D�ݮ�&�A��1�ZB
�(&#+�`��y̱=��Ғ�x���{S4q+�a�s�4~�`�?C5��N�E>��>0מ$jv:'ߡ�Kpނ�[/m�%-	�.I�0��pÉT0v�`�GĖYE�a��'���	�%	F�4�ǌ2g�TLAS�3�s�92il��0��3u�j�����LA�R鳜��iRU�t��{0z��K��>�a�J�T��`�$�7���V?�l�+�{��e���6)��j����ҬY��`7��6��U���t�r6�Bf�b"z�h�� <B^lp ��K�e�74妌1d�QN쥉�A�`1�K�	�gwG~�%4t¡���J��i/C��S��i+_kcp��*����N�%n����f��KNF�{�a�j��֖&��Spڥ��9��_+���0��A�Sf>1������u��f�I�P�]q�^q׋�i����Na��z�UŸdv������R�͛	��e&0�3X`�L��7��I�0�	���f.�Қ<�M��6g����Jq��%ݭ���6ѸJ��5�L�4��ɋ뀙�.���Yv}�.:p�����!�u���a�	��0Y����D�g��'������	k|����%�/4�N��V���O&�%p�0�G`ʘ���-��{��G�a����.8&�R��<И?|d�ʵ��!�&���a���D��_GFe�ɽ|z�%�!��miMfK	��y�O"�/%��I�\<�Y�T�%�1�L���u���A�'�(�4S�D�Yg�l��'�WZ��N���OcM��=חi��#0��2�KoǖtD�ig����4�`�BQ��OON����jh�S�kZ�1��u�i���O1�D���ѯM�DK���~>������D����	��U�"@�L�\�oAb:3���d���6��ldY�C���Q�%)D���;�ͷ��3��N�^�I���t���8�SG�<�*t�S����US<p����4�j"<�ˍ-����[Ω強���So4�keǘi�0�)/2��$�e�b�b%	�&�"&��D�,�0�'J��I B���� DN	�X��'HA^Q/a/2a�R�Oy)xM BDJ4M�H��ykel��&������g��xD��0L0��MN&X�t�
K(N�f�IgD`����$�J$�>A	�x)>M�{ q��J&8Q�����ԫ�gd�aJ$�S��q�\��ot�VЁ��$y{/%4��:u<�d��S����ETŘ�����Z�Q�<��h�i�U�r�����8���k�:����a�����r��%d������Q)>t���N^u�\�-�f����v;Rh�L"���N�E���A
AQ�� �B9�y���8*�	dJ#1Ln�@1Yi�HM��e��\"��N(�1K>8n+<5��u�e��T��t��gs����d/�z�	%#��g�ɉ�3�n�ǆ[Ĥl偝�Y�c����Ɨ�\En>�0]�p`Y�gT��b�b;ZI#�+q�F�.0f����J=�ͻ��߳V�<���F�U��)��>յ*�'�x�AlG�Z*~�ڱU �\���T����vv���t����Ov.����>my�V���#䬥,2���P_�u:�_��x��YS٦�&����|˲Wms���F��j�]�6R��]��m��lR��m;CM}��bJ8	
"��n��X�h�:��h�t�H!TY"�y�3 ~38��D)5����H�	v����,�L�]�d����@�ȵ�Ջ�QSE���N���:A?���DҘH8���k\eab�Iĉ��DW8V���o;�ܿۙ�ř�_�����.fe�1���{�\���g��{��W33=��}�Ŗyn����V��<�0�.����oϟ�>��h�Wci�Z�2���0��|�D8�$�J0��G���.���,	� -�Xi�	�]n�I��p����Yn�b�EF�9i�$�xA9�ACajUq-W.��a�Mk�/�ç��R�b���/��M4�*J��a�5!��pK|3L�B�~�S�ަkQdD��;��č�b�K0�0�;30��fyٞG�Jy-5���v�:��(�����Q�a"�4Z&�<4lA�G��x�F�+����7�A'K,O	���a�]qkq����fb��$-洲�S9��MC��������t��u��-��t\�6'=ː�姲I>dX �䠍�>�Ή�#�Y�t��t�qa�B2y���n��'$�l�a��<W�r���g'��_X���7JdmK��i��̶��xk���~7���Dy���)�a�B|T�䟊p�����by�I�
(�N�&�,O�0L�y�Yuŭ��u5�(����fff%'f3)�CL%�5���[}�|S��mn��D�\���8p'>�}~J8-$	��umG@�N8i֩���(�Q̛�=T�bɳ�{=���k�֩3P�4'NCg�����<4[��thN��i�l��?z���34�r����=0�Zy�V�Ky��[�-ŸD�(ӆ�x�v�v`�&��GI$�D�5�"�%!`8;��|��c0#-:�(�	n ]�5��k�����ɩ�	������3�舖�:�y�aߋSV�Ե��Ҫ�w��!��:�u���I�"^0��gFR��/����"lߪ��xS�d>�&���<N���0�~4�?�0�%	F�t���h>�,��$ѐ��z��ٖ���f��"��e�T���k�A!<eb`�T��l,ќ��ֲ��P���	�Ό(�$8��r��F�-�����))��lIN#4�I�JA0�'\�Ƹ��ŗ�57�N�$��e��֧Y�^�U5o4�]�m�'Dd+4��>�!��_"O9�MN�>?E2L�|��2�Wɔ�Q�u:j2ꝦH�k~�㽑��⟋���e��٦�K$&���%�ޏxfP�B�1徙�Lbr<��>m�����0�%	F�t�ǌ;xf�G>�fon��ʫ7��<�ɣ�'�%p�|���mCIT̰��>�V�"'�O�s��a�rhLM��������B���z~�a�^�|f�8hM�O~:Ҳ�oY�i�2�.�m\?t�:'�R>��M��]3'|����;Lb3�O���x�p�����lч����g��mky帷y��u֜Z�t�=k-���14�s0X�LΪ�D�G!�K)��^�(�����k39�nٔ�e�o��n:�1�ʈ}}ð�q	������ُ٭MŒ3<i��ŕ���rYD�ڜ����𛆍>p�ֵnf������u��--����{G��M	��vw�)âhO@�8{t%�Ѽ�C$�x(���(	p�d�G�Ɩۏ�6���-Ÿ��<î�t���46�N*��B&�5W�)tY|��Ow������M����<4{77<�����E1�a�3bl�!4�Ja����vvS3���2�8'�����a����9��c��ߋ�2O��5�vC�frq�-e)��M�,�#މ�KF��;�S�a��S8iS���u��q��[�x����M:a��ˈ��&j<�����R1�$�(O#�p�Ñ�A`1]g� �,��t���u0��l����{"�=r���]Y,�X_WV�M�J�2B��$�E̩|%����Cd��-�+����çL;&he>��\���`�=6�/a���ya�l���j~4f-6'�ᛚ4}�����화ˇ��'�Ha磆	�55)�ĵ7X�*���iK�1�a��ᆞQL�}��
e��M�b�A��-3�������y%������҄:t�:x��X�<a�	����Ξ��7�f))V�1�8��𒉨���SH�O\�%ܭ�Wjg�b�[�n����Y�6l�4"'�F��R�=T�Y�O/�(���2p�(pNz/=ks��J�LJ�	�"�D�Ѝ�e��p�����`�1�&*���a��IK�HL��A[���̩�\��Xu,C�L��b�[����p�tO&��(�4MK0�OZ�[Ͳ���)+2�� I���,K���4D��Dӂ`�%%���YbY�DH,j!��	H~H��"'�L� �J^<�^S&Tʒ��ǏG�z�I$����&�D!B$yl����������)��4�&��&`�&�0L0�,�"$	�4K$K�4��� �$�Q�@� �	���Ȯ���gf�WO�3��pi&��p��[��6���s�;�+�g&Isݽ>�s��4��D��<��>/7'sk@3�Q��H �>#�E���I�� �wv�J��I�/M��NK�u��Јo{<1����R�BŊ�on�3�+���j���7FD�[o�̽6�[=B�6f�;�1&HMfH<WB��+XI�3��� ��y��*뺇��i��_w��,�o3f�[}�r;}�1ZH��{3���ޞ@���s��*E�b7<��^�=�9�����Bތp�����Ov8�G4�d�&뜲9�vf2���㙙��}�{��|�fe�=�{����33/��{����s9�r�w[k[�������[�<a��l�����b��M�R�,r�ئ�cvJQ<
P쟶�Ѹ�����ۈmP�T�#Is7UU�kI�DDI�̋�4Dl"X�G�"@2	g��W�<7��%��':���V�y�6&Ζa�z&'"5֚i��Kmo6��y��ż��:�N�n%y��T�T��333�������U�C��A�����Y�>�<��HaRpȟb$����~�xQ5��g&��{?Myco���)� y�ׇx"&p�83�rvt��	���I�xp:`x�0�N{�n�"t1D8d{�m�T��Z�����δ�-��<��,�%i�O3�b"���y���'��0�c�5��Z�\>�z�e�e��ݕ�Ӊh��ȝZ	/4�Z�"��63QΚ����{0�u63�Į�)E��V��I'�Xt4�6�.؍pCbgi��h��6ٵ�$^� ��;���=_�kFxR��=��8{'�����ϸp�v�8&�����.eɳ�s�1>ɳQ�?L8&��,=6�b'����2?A(�8:|�1��u��WYV�Y5
��x�x�P�4'�{���o>Lʙ��9)�����L(�L<h�xD�ǋ<%	F�t��ӧ��dSI(�$�R)�!u@�T3IuE@чV#���c�L���i�Ұ�l�p��'����zs�뢂!�+�	a�S�e��ɍ����g�q��t�|P�pG58�&.ff�]&
�O�z��{��� ��=���XN�q.÷����q�
K5%虎�m����[�e��uո��qkmo0��ӫ[��SUQҪ�O!����G��z�,�{7�8'��^CÛ��;�ТxF���-e�Fq4
!rGd�0�P�%5��D �O��ba�Ǟ�qײp�f��ѐ���9L�^�L�r��1���仪����'Ƀzu-;-��x�<&���L<x��P�i�Mӧ���}joZ��K�UX��)��}V~0;8~d�}��b_{Uuk�E��sM��K��N����~5�'�Ӫi*[��������ӌ&�5��4'�MC��0���*�ܞ�wm��+�C��4O'D�ϩ��hB�=*�=��	�JNq5>�N�����ξ[�y����0�:��_�-�u�X���a@�DD̢�l6�!1mɭC�v#К[l$��_h�z�5�Bҥ.�Y�X��M)����9t��f���U�O�� x����EV>v�B����cM�Ắ�	�
y7��}������a�D=8nqSA�&�������3@��l3�,�ϕ}����x�"NB�R�]�քˮ��@� ��ݟ6�ix������5m�5�jN��S�}4�ѐ���%�Yy��:��-m�l<î����h��$�ό��%i$��!�U�m��j=L9��:�z��˓٨p9"����K��3�jQzN>˩-�s���UR�2�"n��",S�5#�F��Gσ�6jM�����3��f`����ħ��'���3����L:���|�-m�l<î��xzt�g��(�uN��Z�CV�-�IYUF*Ŗ��8Q��c(��E�f�q�ڵF�N������ٳ�(r�%8v&4�]�'[�fS)�y�E���'�d��6��d@�͢�J"��u��FB�l �I�fpA�.���!����CF�lÊ�B����V-e_vj�L7o��Y[a�7�͸�.L��í����yo8��\Z�Z�y�]iכ[������Zm. �iIγh��a� I!�\�e�#Hx�%K�:��c|�q���gX���F���TP�Ae&=nNH!���5*.�PNa��絷a�t�y����;���(d?�0�NKi�l���q6�I�����h�6C!N�p�8�����`÷�K��������3�߷��.���}[�=�M)e{"��R�F͛7���??>w�g���ߑ��Y˔�8p���0l값K�dw��&�dsrJ����{��DBȑdYE�h�"h�E�[DD�����hЋ"h�!�Dh�,F�",D"�M��&�dDH�����b-�DZ&E�B-�h��E��E�2-�h�DE�,F�E��Y,�E�H�$YDF�B"�[DD�`�"E�,B"ȑdiD�"��M�DY-�DD�h��	hY�m-�A�
D��mH�[I$�md�Y"[H�$KI2��BY&��ZD�--��%�im"[Gn	m$�D�Ķ�-�D���Ki�D��L�M,�iiKi4���M#H��id�dɒ�Kil�-�&X�$��[H��im"e��m&�I��im"dK$Ki4�m&�L�d�Id�l�Ki-����IibY%�K$��%�%�"Y"ZD�Id��L��Im$�Id�,�-$�Ii$��Y5�Y$�-��I,��$ɒY$�-$��[H�E�K"�L�dZD��-���d�,�$I-��#I-"ZBY&K&Im&�I,I$��-�K%�d�dZd�-�K4�"Im$�iĉm-����&Y$��Id�[I-�I%���%�Ĵ���Ki%�%�idɥ�K$K$Kim$�H�H�Y-���Lt�Y&�H�-�HI�ZD��-�H�I��Ȗ�im"ZM-&�&M,�,�$��KH��Id�[I-������m$��[I-�L��,��4�!,�Ki����HK$��4�2%�[I���[H��&[I�i�M-���E���HK$%��Y&��i��$Ki4�"X�,�4��Y!,�K$��&�I����d�,���I%���I��,�Ki4���m&�m!,���im!-��-��M-�%��F�Kd�i4��Y"[I-�&Y"Y"X�[Ki$ɉ��im,H��ibM2�D�(�(�K8��F�L�4�ɶ�p�f��I&œ4���F�f�f�&�Ѵ�$�d�!�6q�7��&k&$�$" 1� ��7��5v�Ӂף�h�dHYX�m�H�$YF�4Y��DE��Dt��Ѭ�BȈ��&�h�mE�h�&烘s�4Y-�Y烘rE���,�D�h�8��""�H�",��"Gq��m,��D�q��M���bˎ��-�E��YF�dH�$H��ѤH��E�Y�"�$Y-�"�"�4�D�\3�"�"�$iD��"�"�$DkDE�m"E�D[F��H�$Y,����"Ț,���ș�dH�&�4[E��0�(�����h�dL�dL�"h�",������E�"�!d[F�H�$[D�!"Ѣ-�h��",�h�D�dL�"dY"Ȅkh�D�m�di�Ț,�dM�4Dkh�,���4H���#B,�h�dDY,Y�"Ț,���&�""F�;�ۂ�[DE�4H�4E�mЈ�"5�mDE�d$YE�-�m	D�dH�,���DF�",�,�
"5�"E�m!DF���DB�E����h�,��DF���"!2",�F�"ȑ"ȑh�,�"�"E�b,���dH��"-�"�#Z"�hZ5�H�h�"ȑm5���$M�"�$X��dH��"�D�m,��dH�G�3p�D�"�"-�D�mD�h�m���"�4D""Ȉ�DYE��-�"ȑb$[D�h�"E�DYDE�����&�h�-�"�,F���dYE�4[DE�i��[D"�&�h�,��YE�h�k"E�DYE�"ȑdH�: �E�mD�""����"�Dh�"�!2$Z$[D�"�"ȲD� �dME�,��h���4[D�m���h��DM��D�d-�"E��H�9�n	D��"ȑm"ȑmD�h�dsZ",���� �D�DD�"F�H�$-&D��"ȑdH�dH�h�"!h�h[E�H�$,��-E���$!F��MD�DDE��Y"E��Y�DE�HX���S<m�\��^�ۖv�;��3�������33(�ƴl�Z7[oGǖ^������;��^?���s���՟�=�����}~��?���$�����ў���7F�w�N��xy�����w�ɝ�����zsн-Ϡ���^N7y�o�/������I��������yf͛7�g���8��w�S?�-���������o�X͛7��&H��[��~l���캿 �z�#�N��,���6��F��$����+���Zu|$��+��c6l�������*$������n[�ۆg����m���y�r�5��>����,�8�͝���0�pn>Nݻ����{?z�׏/���n��u�文��o����gM����7���6���ٹܸl�3m��0x�1�6ٰ�lft�u>�ӝ�#��p��'���������ޟg�y7F�����m�͘;#7#aD��6Hfۈfڌr��A�|[��4�,�ۿ~W���7��fE�m���ٷ�yo7v8?�x:����o��C���{�lٳq��ӹ���߃m�;�����m����#����nǠy��t7��� |�~v�������l��g����K-�s�On��ӏf>��<~7��~7��|f͛Տ��#^~��h�q�q�������o���=���g�z���l�u}8͛7�=��s-����g��>7�v|�N��}�ۓͺ�:;<��C:r����ˆ6�v�ǭ���nUs�]M��w�ccl�lF�G��z۝��|��-���[����ۜc�����c��q��q�a7+s��n��s���+�w���~�6l�lv7������x�Onۯ��f��n����GӞ��6���Ǵ����@�F���g��&s��V{�_���p=��<����dm���r|��o��c{|�x�Cf͛���g�dM���~ݷ��f�7���=���?SQ�{�|OVyg��g-��w��'{=}�ߔӻl���������tJ�88c�^M�ܜ>ts��X����o��<m	0y�?3�C�7��Q���1��I���f��[o6ޞۦq�q�&z�f�o�����y�޶�7��=.�ߞ���~L|�Nݝ�l��|5o�~�6���bf`����Ź�xr=l�w�3����n��;OK���z�St�S����v|;v�������?��|�Z~��nr4m���������H�
�^��