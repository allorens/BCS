BZh91AY&SY;�x[݁߀`q���"� ����bEW�           ��T�)U
�(�$�)*U(IB�I(R�A$�J)E�^�"IT�+l�UE-������"�kMz�RU	H]Q4iRYT�Y���P���P%!21&��()J(	�%JJB�M��"���j�E�  I� �J�SBfptE]���D!U*ж R�J�%R�J���R���"m��
�m�(��SF6v�
+� h  ��RH@�tg���|���K��eX4wm�`4-T���m0wa��p �k��SaKP
d�SUY�a@҉U���I(�>RH  ��}$�<;���m,�\r���%w'��J�k��*��=��uE�5ίw=�
U)��ǩ(R������(�s�x�B�5M��dV���T�)ϒR ��ﻘ�)J��Ov�:i�S���OM)S{m�h=)@��h��z��T�
R�s�B��ҩ��{ʠ]�*�;�ׅR�*�t�{(R
���$�S`¥J%E�|�� g�R�*���q�)T�P����R��{�צ�J�t��=R�/�ޡUEޯNx���(s�w�T����YH4iy�� �jt��J�(HG�$�  �ް{>t	*�����
(P������*��̘�I[�P���wT+����T(J.�u@T�Yv��*�B�oFt�J ��JPփZ�[$
4k��R ��[j]SnK��U:a�p� �B�d��(U%g.t�R��j�"%R�D�m�@Tn��Z�E�7*�%M6:�� �{m�UM��X-R�|�� ;��o� `}��ޏp un� 5�� 2��M{�����  ]n ��� :��bJF��x�T��  7ݮ��H�. �:��r� ,� �;p �,uC��!� wnop= <J"�f�#e��RUli��H �{�| �����
��� 4��{� �O[� t�  ��N��� �{� ��@��IUB3:*�䤀s� �W� :qv�M v���s����� {ǽ��on@�k\ �0 �     � Q@  L%)R�M M0 &hD����F'�i��4F&A����d�*  �    T�"dU%F&4 ` 	�S�)HF�P@�  �  ��RIM2h�	=�7��lI�3OP�'�������p�o?�����?�z�룷�j�3$\�|����^s>��?�P@U�?0 ����_�,����,�G�?���G�>*���PV��T�I>h�T U�d~�����
��������l?k ��>1�b�ضŶ-�m�l[b�6�� �-�b��-�[ض���l`�ض��-�m�l#ضŶlؖŶ�m�[Ķ)l��`�-�� �	lB��b��-2�1m�[��`�Ŷ1�l��K`��-�[�S �!Lض�-�[�l�,b�#-�l؅�m�[��l[`ŶlB؅�b[�-�[�l�%�b��)�[�lB؅�b�-�L-�S�!lB��b�-�[ �[ �ض�-�[ �	l�!lB��`�-�[����-�[�!l��Kb�1m�[�!lB؅�m�`��-�F[�!l��bSش�-�[�!l�ib��%�`�-�S`�-�[��m�[ �,m�-�l`�-�l[`Ŷ-�alŶ�m�lb��6�-�l���4�-�lb� ���-1m�lBض��lbF�`��-�m�[�!lm�b��6Ŷ-�m�lb��6Ƙ�2��-�l`�-�l[`��F�b�ؖ�-�l[`��1�l[b�-�[ؖŶ4��4Ķ-�m�l[`� �-�)��i�l[b�ضĶ-�-�lKbF[ضŶ%�m�lb��6���m�0-�LضĶ-�m�l`�ضŶS�0`� �lb�ؑ��m�l`Ŷl����l[`�-�[-�6�-��شŶ-�m�l[`� ��m��# ��m�l[b�ضŶ����m�l�%�m�[ �l#��m�[�!l��
`[�
[�!l�F!lإ�`��-�[�-���!lB�%�m�`��-�[�!lR�[�؁lR��Jd`��-���l����؃l�[`��6���m�[�61m�[Zb SB�
�V� ��`�[؀�V� �V؀� �*6� �(����@�%�T-�-�@-��lm�	lQ`+l)�-��6�� %� -���-��lE`0���� �V؂�[`�l@` [[`([�Kb�l@`�[[`�[[`�lm����"��V؀F �b�lm���� �U�(���*��V�[X�V�"�[`+l b�lQm���@-��lP`��Rت�[b [؈�@�� -��lQ)�6� �
�P-�l ` [[`+l`�[ m��`�B�(�Vت�ب� ��تF��P�(%�T-��l`�lb�LT�(�1 -���@-�%�`��-�)��i�l`Ŷ�m�l�S�4Ŷ�b���m�l)�[
`�l[`��-�m�l�[`Ŷ�-�lضŶ�m���-1b�ضŶ-�`F6Ŷ-�b[ �-�m�l`F�`��6Ŷ-�m�lKd`�ضŶ�m�l[bŶ1�lb���m�l`�ؑ��m�l`�-�[�6����m�lb[ �%�m�l[`FŶ-�m�l[b[�6���m��0m�l`���m�l[b[#�6Ŷ%�m�l[b��6��i�-�m�l[`��S���Ty�~������Ez{���s��.��C��[T艣<$���^�fI�*�wVe��-� �%�vV:,l�fLA�����ÓYă��R/�j�<�.a�Di�FE�r�U�w�k<%`e�f��'M����#�������h٤�^Q*��PǴ`�0�7��1��r+s|���큘�Wq���v�Vw_�/��p��{x�	�!4fਜ਼TC�i�T�i�c�˗Vj��i��F�I.���sk{YP;�ͥvږ���*�:����<��7^���
16:������6X�P�U�Vv��2��z���7Zqr
�Ie'�5��ds٤��I�X$+6laP{,�͗��	���3��;ϩ�]��)b����7{SZ
�=zf�!�i,˛�n�ܼT�:T{KF7,��c��U���7�+(����i�%��^����L�<�(�l�[�6��&�B�N�nݴ��E�5��G�Tƫ����r�m̭�Q�4f�0��R�
��� ���X4E4�ݬ�z�e��N\2m����QpI����7�`�u�G3�JB�]��n�l���`2��j��G2�������4�O^⭀GHl��Z��_�˪�jH�1*JES�+nXB�A�����G���R3�i��7A�Yx�a��T6.���e8�׷�m��5�@nc�^����l���l9db�VOLef�ͩ��Ǌ%�!��լ�v�M3���dV��n�C�,�[(�i��B|�����i�v�Nң��$��#	Y[0��#.ٽ�Y��f6J�KҬ�Q������/Jؼ�.�:W���K*�0�V3h*@��hE�����y: ���c<�m�
k7)��5:�Xjl8�5�R�S�7���8�K¬(�ƶ�[QJ���ǈ��u$�R'��vDZ����ئ+�к4L<����ܴvx�����fO1H����d�7/\���He*��lQզ�*�ՊR�aЕ�b�;j6�.[���ҷp(�E�ؐ������CP`�r��+5��7qZ�̠i䦚�BT�đ޻�F�R�`Ӈ*)�wj�[�"m訔�DɊ��\�32U�Ê��M �+��M<i��^`ɏ�&�e�;��[���S�Q䧓E��6�;��37n�5$&�n���Ռ�g��Ɇ�B���v�hua��9�r��;�)�e��|!É{dڻԬElp�KU��I���l�a��4���{ �ܻ��N�w0�- ���c��d�7BU�y&jP�&S9������7IB�36nԷ�V����d� 7��3!�cINZ�v�<��YV�èL�XSf�-Y�X�H�ػD�8)ږ)(��M�.���We�P���Ul8��k�-�Ȧ�5�n=�Tb�)��U������)j�ȇ��7Ls&�RcmM����E�,�,KI-���~^hn�o\�A[*����"�^H%SsV^oUU�*v-�zM2�5x�j�:O*{�����pB�\;C�v��	��+c��Ԫ�$U�/ֽh�Or{eER�j���AYVU^]��ݪ�"ìAT˳��i�^S ċ�K��X�f��7��@�:�1�U�Y�h��/ZI��ۼC\ܰ�ҩXT7n�EfQ[T��r��#p��;LH�,蹷*m�	�,%R���Ǹ�n��D���>i�'2��ʓB�D0R��j<�a��n��N]&���Q�� o�Fm�f5)�4�dRM�qZ�F�T9 l�F�\�6]���i�Q�ԭ�wcv�qm��i(�p�+SVc	=�+����2�F4����m�mFne�zנ��%���3�T�e�U�W��Q��vЬ�����ufK{�.L����mU�1����@[�Dؚv%�1���#��k&9��V�.�hÎ�;����(J7y���1�4Y�z]����Mn����Q�]oqe���QY1ل�Gn��� �VX@���4�Vcjז�ao.Ǉ��hm\�ΥY��&$71UAR�ƪy^�(!Be��N)�"�8�#p=�<Vk�H�t�����Y��C����5[�pD-�ziYTQ�������/D]QzN�Y��܇%E �0�b��EЦ��b���XxTPCuj�i��Xޛ�⥶Ա��.[�r��%�л���{J��m*��@ZVђ�2�y���ݻ��Om��@�b��$��h��[\�Bi2\�	�[N�w�Z�1�{	��޳��X2�TM蕳#�j�S6nd4��c&8��oZʊ�e:,
P"wN�v�VC�si��n,æ^Ö�`�	S૑G�˔Z.�iÔd����n�;�n1&��r��ҵּu� .�<֓urV�nnMFU���<��fPI��Ȳ�'���y�$�J-b�U��GfZE��-.�1X���6�V���f֚��U��	ܔk�tjKu�ٺh�n�uO�,9�/7�=���oR�x-9��6��k��;`��*�>wbR{�y���R㬕,fSz�,.��7��:S/M�˫64T�4�YNT�-�-�-j-hyB��Ӷ$;e�gԮ���
�SY�Y�Um)N�YxB9E�Z˔Ֆ���_�Ǖ�t]52�nTAAt(ؘ��FJ��1�iǙhD�5#u��S$�V3w�Nc�6���\���Ƙ��hf��6�XUf���ô] ��X���4k���5�UnGjV4�*b٬���0��w�x��`;��<�]Y�2I2�L6t��n�"5�ӱx؆�LZ�y�p!Nk����R��Lq�fV��6����	�:�inҙjK��љ�ܛ��e��Y-�RQGA�";$��%�]g��fCwx1�����):	����ƚV7}��Y�Z����!�r�;ۑ$Z��P�0k� e�V��7�����	J۷���Փ{L�Đ�Y�F�b�xEb�$fn���t+�U&�iջ�nXJ,�s�i	h!j�a�1K��V(�����(�ǘ	ݬ:1QV��љ�,����i�7/v�˭�t����%`�1�ě��ӱ���t��o%�N�ХkQ����zv�<��ʭ	�<�)G3J�8���xΚ�E6���÷v�,�Ԗ4���l����%<��&��&L�5G	�Y�F���D΄4H�P�9J�u�zbV0*����=�Q�8��[7�ڧ�k#}Eo�"�ͣWnJ9�Z�� �)�*�YfeMng�[r�ƭ��I�+�PSI�n�Iy2�I���m];�P v�i�	/[�S]cM�xP�.�ٌ�	�{nn�-X�f-�&{4]lz)l�fS��UG/5�ڼ�3�x�]f����ЗQ+7��H�;A�4���+RkmL�M.ˬ"[v��#Tk&ɺ�0����U)/!�7r�i�n��vóm�X"S�V�p�I�M���t�#]Jsi����z���Gkm�������Ғ]c�ݗi�v
��2�i=�5n�nJv/d�E�勥��E��C6�x�%�u]8#�Cc��~�V��W�SMܓN�Y�Y{Q�KY�0�;�U`�B)�%��J��kn�z��Zl�1j-�'j�wN��������)z6�&�kkl70�<t���X����d��S.�]��fܐїv�Y;
��ՠH�i����l������!^�*j�X&Ex�f�۳�.�ݑ����T�{���֚�Ñ�30���^S5h�@c�6����ݧ��M�KMd̤W��Z�@�]�(%,x+�mZ��۠�(�D�,df��d�RP��ge����ب���&2�����*��e�Ў�f;oF���ֽ�+`S�N�jAJ2*�D�tD!���۬��$Q\˗�&��A�i!q���z�\�6�ә�X��d�hF@ܤ�m-Ņhi��R!X�.�M���۷���h��KO*�"i.R�PMn��$+d��!�K�Z���o	�VjŦ�^��F�V��T8���#G,�~;�:6ͼb�
� ���6M}[μf)�q�q{���h�M
Muck2�f�Bfȅ���#k2�("��)J��G&2���<��a��5t��fe�4JNT�,V�&l`@���Їv�*D�rm�Af����{��8�wHfj��:����MF/�9�Ve�v��!�,�J��V��h*h�v[;X�]`ݤV�څ��a��n5�1l�hȐ��5��F�ȋ�[��5���Omҹ��j�r4������C2Ae৾
Y��f��ћ{4j6��B�����x�aQ;�R]�FK��^S��pG�å�ƭ��"t6qP֡���M�N�wF�jٔ�m�;��V��M��uLڙ���7��t�X�X���v�h�"��`3��hP;��e+���v�e���.�~PnD*�V��d�ٔi��Z��ȷkNɘe>�u��ئ��#X'��W��(�P�˽�n���&B"���Էx��l,\u��,YC��m�-mش�	� S[&3��"܃<T�1��92��v�eX�wj[���,�2��Va�l�r5��aG\@=���G�ҽ������lń��\jP��
����"Wz�Z:� �:lcWccKUj;2����K�yCo\Z�B�j�Y�[R��qQ��җnǻsjM��e�B�ڴؔ���A3P skof,cX4��=mS�h��3$��[��fRvM��V'V�f��i�Y�YM^�m��B��\���[V�*;:oI��2�V`JJYNU�p$�7��ȅÚ[�w/%$���x���
Ҵg���=*j�W�������`��l{{*k���ڙ��i�r�X�(Cf��ͪ[�i[y+D�rhT��j��:�+*:z%���z�,���`�O@�d<v���V�MV�B����bο\EICT�
H���I�dx^9�]A=2��Ą�`�d'$W��DSf얳n�t�K�
H�Q!*�/4��&���c�q㣍Q�e�Y���cZn �ٔ���T�k'\xd�I��6ٶ�ɋe�A'Q�K��e��戞���ʶ�ET%�9�fVU�y�յ��J��7+YD^;�#�����T�P�M�W�r�[��u�n�ڷ��#k]�6�E+�3Ξi	�,PVʫ��f6f��RX��F��asXZ-R�m�L���XTV�xa*b7NmR�yp��r(X;��-n����ӔkL���i,8��	d����6�{����M;( iK�yGB�b˧l�f�	h6��;~r����6��ҡX5YK�sK� :�[e�CQ͘��2(��[����&��F�������{ B�6�5�wSl5P����V�\)bD��2lU��T��Jٵ3h�f�ȡֱ������V"XN��Xbq�88!�MіmP�r���VeV��)�Xc7�4͍n8�(K�̽��n�e��̨�f���]�i�	���Y��ͱ@5M�e����ǡ�{T旓��a:q-���ŝ��r@S�d�1����\4��TF�V*T�+UJbf�hV���Xh@�[S^���d��%�n��.�x[�7��cW��m!M+)L��/%�ʹ)�/31�����Q�1�v����rJ"�=�ot1��˹�+nar2�*��JP'V*�9� ������z�lA�-�.�J��ƕ��w-��d���0\q"*c+U�tnC���M�iSn�br�Z�z�d5yW�#����D0F,��P,[L��~�C�5��ʕ{���csV�U h<,a�Y�ښ����`���ni�Xe,�M���R+8kI�裻)�gj�
�UL$R��[��E�& cc2��vEP�[+�N0�j$�6��"�ϰN7L�j
�̧�2�S3v޺U���� !&xc�
��Mn�Z�XB��Q�j�*R&���y+(֩�JҮJդu<=��5�Dp�^�&����9KZ���iR�H<�Z��4��][.&oN�]Ǘ78�c=	Ì���n&4v����idLfl��S�)H��i��Ξr����v�D���U�P�{L ut���<F�%�j��-ĴB7{t��"���U����m4�r�]�H�Q$�'��i dDo��3�C!�]Y���i�&�#4�I%��c=��4,��a�T,�^���N�4S��E܈'Uj1^,�V�(	�iV��r���X���R��-����3't�$���V����;�3�dG�je�[h�W�� ����kV��⚠=k-.OT�A<�\�Tm6��4�qg)iR�h�ה��C\[I������OZ4yL]��Q+iEX�V��*I&����DY�]�eð��FΫ���Ia�e���{	�Cl����(3b�ޑ��Q���,W�5@�U#Yh�FɈ�8���Zl���x�#�sH��<�F�o�ċ/
U���[͟-I]U��U��mD����UKR�OR��D�Wj-�Yj�(�(�k�RU�uvG��u.HI$u$�*���)dY�!��(i3NC/L�H��LKRV���Zc�:�ԔJ%i�f:����P5�l��T�шj�K��Q;�C8�-��a�%2h\8H��9��$8��aT.��V%Y�)t����7@avF��hr;
�iK[K��H���Nj Ǽ�iT|��(���G�C%����ȕ��,Kn*J���h�y[�9H�I�İ�	��Cܑ�ĸ��0-�l�N�d��E���ITK�L\�F��*��e,
ڣ�m�-��Y4;j�r*��F�JT82�$��MX$��A`��H ��Q�R�9�*ɍ*Y���3a8U�H�(&b1)K1(�%_Dͤ�E�=Uh�mV�P�������$2Q$ޗe#|cE#��ݜ���U�щ�Tx�����6u�E#,�ӄ�J-��4�#K�٥���9��q,��RԈ))IR�V+�*�ū-=Q���N��	�o��� ����$޻�r��x��u��o}� ���������:����Ci�껹gy�5��s��j�t�Ӕw(&���]qp�P��s�w�8��G=闕��X��d��倞S/��>u�0�k��jW3UY�q����5%i�)�Jg;����¤$��Ȇ�jt�<ټ-�v�no_���r(7�ճmZ�캕�������AV�ڶ�c[����<;%5��r���Х�c
q&�JG�.��5oss��>���#|d�l�8-�2,(wMɨ�/�Hv,uڌ�Gj��-]���<�󁘻_`��!F���ә�S�*�x0x�R�Xޖ)s�e�8w9t7���y�ڢ�vu] �<6�Ҳk����{�5{�����$�@m�}�ꚽ'�:LW-(ܥ��a�׈��{]���}6��t�t2�_�*J<{VU��Mm���<t��7��C���;��̻;\%�
��݉�s�rl����8o�`����sN�Rǒ�Tv��Z��k��䝆Z�=:	�U�>���\-X��j���صc�L<�s���;�lXkOul}s��k]P���7;7�����O�	U�vV�=O^]�OmE8ګ���}Nf�5�5����Z-����(�jirZ�ʰ�Ti(�g�5�7oJ�h5fn"u�ea�����<�r�B�Z�
��1>�:��ˠa����]7O��bu��V;ԷBu��2��)!dtz�!j;���Yͷ�X�G+�}�����GGh<sdJYЦ�=�M�bh�hbyA���;���4�'f ��̂�p���Ǻ9��!�u�QG[��7U7�v���]q���]""���ξ�dEwzU0�Y]dZΏ���,�xԫ^T�2T�n��|ݜ-��{�㋞�{���i���fU4O;T�H}(hE�H5�3t%uK��t�N8��L�6��!��]SP�2�o�=7!�/6��z��>��N�!V��ˋn��(q��D�|�Y;C�4/���O��`~{Y���Uhz;�_N8t`t���:�*�ܨ:��B.yǰ�oy�t�]͡�Qu}xNh��ňjW!*������C�˖��GM��4P�z��]���wȅr[��f�.6��f��(d�bHd�ז\�y�U��l:�u����+�R�z.7(AI�9|�֢�;.-)�8�9dҽ�}�ٻ�������gE�a#�q�<h[��ʷ%�\��!�/��N!$�&��J��P/d�l��Wuq����X��5��m��:�QDu��H,�C{*�>���oHk��R�--�{G�LZٲ�JXa���Ucٗ32�'�r��I��ά���n��S�eP�7��k%q�Ȣ�2�sq��{�Щ�W�n��
��7Y�hl���
ζk�)�έ��N�U��E�8%�hے���\go�:/nWX�6�	���ܜ��P=���Ek%ey0����.A	zy�k' ���Fڊ]9�MWY˿��\��ٔ��at%���/7x�w��u-̫ݿ-	�IŻG
������6������Y����$uh�� <�^��U�6W8�6�H3�L��C��QmUwY/3�%eދ��F�3�nwv�RciD���Β�����Y2���њ�Kp;���k3�X����N �4�EP����%Ïy��=V2J�m��s
����u���S�N���}�X����a���U�k�)/�\,��t����B�I�<�&�%9��M��uK9]��͖*���ܤ�nԫ�*j{�b�h�%���yl�[���9�Y��j5�:�:i�v��Zq9x"�yS��<g���>y'� ���iYeMoZ��c\��{[w��/�L�r�جl5�c�s�vQ{��ʢ�.�a欤�p�ETp�Q]t��3�a�VWq��.�o���ܬ}V�ҳY	&{9(�2�y��	������:�b��)�7vƃ��^n�U�W9��ḎB����s���u%
MN������x}���M�zZ���(�켋t��v��K����zQb�7��و� .�x���p]��J�5q��{�
6�L5��w�jG;h����)j��F51|�� %�Bٚk�<2�̺�c5��]�X�p��{�cl2������	$^�B�+p�gC�f�S(��$f[܏B|o:��1H�t2����ٚl;\�Q���a�.�\�%�]݋S"c�'&6������J��T]�bMw�w@���V>�[Έ���r2R0��D��\Z+�����d��n� �͕�}hn1Sb�a}ݐ�ci{궏�ff��jt��.�)Ś�*0㧇�r�hbf����K�
�v�v�k�P@���emN=F- &9B�i��T��f�ֱT��v�v��V�^Y��*u��)(q-���2�ٻ�UGK)7V�[sVe��=̌�%V�Y�/��tވj3j�d�ӕElSm�����J�+���K���w�l]��gKVZ�������]���\���tk�_�!��u��殼z{��Ѭ��;��{j�%sGk��t}]��"�ek�Z���������(�c�򯋲�UW�m���#	nཕW_Z������6R[��7�V����jw��	�r���V�aFƻ鄁��]&b����"��k9͛���]%)��>a�Vc	n1Zs'��F41Ka�i(��6�Ӷ���F��#�����]
�]I�Du6��wVt��{{��X�d5Xۖ�\k����*u�q<�����h_\�C=մ_R��&�ή|��*kp��_2J�6��w��Vv�wl^�2����v�%oQ��1�@R��[���qr�P4��D';,���n��8����zJ\<��uy���c�V]�X�u�ib��ػƺ=���,X��@��x�Qo=�[34tݐ\O
�q����F���mݧ¹��`#��o�boWQ4�[xȀ���;� s{����������� ͆@ډ|�}9�:�9Z+9�o,<ܵ�(�y��j��v�	̅�y��IY�N9{�+�K�PC��E��0HP�<^+����u1�AMx��4LҴ������e=kN�{)�T���2��7�v\$WYD�e�us�g�S'�4rtT�ICR��K>�����A(op�u���zۏ�����ֻ��v�@� ��)�/.�-�U9D�+�]\֤a��#n����Ö|�2+$�d7�w'w�����ƞ�|9�5�]̸k�)���ְƜ�-Q=W��P��Ǝ�J�o����c���E��E��v���1s]�K4'o��֍�����t���42׆\��)��֛r"][f"� a�"]���Ys���%�8:��ݮ����DgU��$K4�=[��yv�Z2^�ƀ�a��sFN�a�`�e��֫D�-́k����V;�
UZ��=����v��2����i*,*M��q���oZ:�Eމx��<g`���0qȰ`&�����m�uyW�Үi��Mt7�MYA�c�B�g�����\�����H�0t��(��<�-$�#wj7���r8����w6�n��`�EEݧL����R��F�Ӗږ����������̋�	�~ކn�]���������L�0�!C���¡s+8n���(�s�
�Κ�9O^��#4�h5���z�ty�X����1��=ݜ�ե���f�f�2`����YG:��ravH�ѹ��Q"¾<o1���WRKz��a�3��ķu�Lv;j��@c��ʇ/Nhm�\�o�1���G�ԗӺy�Ϗ����z�-ܠ�@�ۓ�ڲR��e)oPQ7w�n�0��dQhө�6_�ë���l_�w�ꏔ��Ct�I��|_=���ݢ���S�ek�{������Vӝ\�:/M�#
�ii�'Yq�Nu<E��]�f.!��^���<��8�=	a챨�ONx[�zM�"��u44�Y��Fe�N8�u-�y��Cq�ks��OE�+a�Y�����q�ް�C�Ik��`��^sں��Eך	e�rN��Vi�nR��g�Wf�!ϛ}�K�P	Â�֌<1�o�\�+�\�gIn�d��.̆Y)]��^����r������Yڇ;1e�W��[�7���n����N��7��tk��=[1�{��-�[���=�h7��K�L�Tph+���R_\�&l�|���4 �[��4q�®���Wd�[k{Dّ�d>`�Xיg�	�ޓ���9�oz�(VR\�V5�x��]B�t�K�m�D=�%�S/9`�7y]�N����oPO����IJ�1�;qrT;s�<�Y�S�� ��5 �p�2u�H��a��98��wa�To�rr�N��S���v�]�d��b�ꦗ;%���xWvaܤ�[W��%��p�ϞL;�DI��RJćWע��5�t�����t��p�ؼsO�,��o*�{a'Ab�����v�L������1TO7Ir�T���r�7Nv��M3l'���̆�jl����u4���ii�ՙJYއr>��"�}�^�NT�����������Q�K���܇�^;Rv�M��>��[Y�9���\U��
��֐�kg8+�o.U��+�4�/��X��N�t�Eo��U�Koi��m�͝grH�\w�������l w����Բ�Ƒ篑0uSu��f�;���DV��gXG�r�c�q]I���np���{�)S-�^����q�9�m��@��fjf[Ts�L��dצ�y�Z��\z%�$S�i'��iWn�6u�h���<f��z�����_-��V
��1[&67W$�1��-��j���\X*�@���}���޸k��Hn���leu���5�t&�ur�}�M��jF.(�8ƺ���n��o-=9,���q>�dxĢ�ɚ,�"G�gR��^ˆ�z��v�r*�k��2N�ݝB��#1��:u
��nfd��`XA*%N�a�}ϝ\\�Q��;5�ڔ�Xٱ.����f�����q��q�hT6.U��ʚs�t���KSչ��O]�յ��R��Fuf��q^\J��.v�7�T��4��U���.Z��'���%���\�5����j�s7R��|�G�	��Χ�
���]y�ȅ�G�3�-}7vɹUӑ�;�
��`��Z�U�1��k$�������Q����j�:�
eRu}�s3�P����op�ǐ��h���èw]mƂ/�W��nq�NYN��ड़��5�k�u����X�a��kwVtѩ0���(��|-���u��{� X{Ro���n꫱X�K�����t�/x���m�.����A�G(�%x�aG:!��JH���4q�j�����yÜ�`�˻���(@ދ���-ހ�:N\��v��������_Q�8�w�[!M�kY��\�ѓ�W$�]�>ͥ	��PS����O7��s:�=�H\�0�;xE��ĹP���m����ѥQmاaf��iF�=�\�q��/7q�F����D�48a�ޔ]�r�ӄZuV4j��{��td��\�U����Jw���^s|��	M��[�^h���;u4Fj�DJvk�x.�	&�^�`�γC�J備�d�ӥ�&�CshM���T�*�������̧��;�Q��#�����2�=�7Mu��xw8%\YW��_�/�m��XkP3�4*ץ�t���C�<���U��c�̚H�e�V^�"l�خ\:Bj����ޫu�h���=xr��k� �wu���^\�������w!�gk&`<{V�BR�L�yw.���#��Ǿu}�����U�+쳥�V_Q��ۻՎ���{*Kf6���5����Iy����Wp�͋��erwPWh�Is�}��2�{/N�ά�}ϣ�ܔ�g'��6���:�ΝB�b:����\�;x�{p*����IWNY�:�V7�R�f��p%Og׆.���#�'�zC�a ��,ȉ�$;;���)����ߞT�jH+���� �y7. �{V��<��&��x#��"&J�*{�}�{!�V_��'Oi\�D<��$��L��jdWr�;��r�B�^y�@7Q��D�!�(�D�ѐ �K�=��ʮN�C�a�����4Р ë~��qD��\�I���:D9t�N�7��n
\���_wh������n*�R �|�d;�.B�J{73T!�/'��J�b'�����y;*�ߔ��\�g����p��Q��?���DPT;��	�������>(
?�����?���%~oͪ<~����<+\��d�JJs�ѹlk{��U�w
�J�/f]��]cg*��w�l9���։HeS�ռ[삍�����Nh���<���;zfi�X�T���r��ห�eˌ�;��%Te�wr��Vb���S�\1	�M��f_mؐP�f�P;M���w.�61V�cdѹ��I,h�ڰ�GA��lrMKy4��v��y��ҡ�e�62nwT3�9R�f�֩�W[WK��J�ϗv=2Ř��q[�%���젫Tpel�oq��4Q��"!-F��9���5�j7���pbJuҢ�'Iy̬ZrL�@fG�<(W:-�x�ک��v\핝;�u�����-��Q�2��1�]V<��\˃v�/k���,�ӍձSnYe=4�M;��8)R��>���AQpA5��ˌfSoŵՉ+Lq�GU�ޔ��t߆��T]k���s`�&�V�r�9�{��Z�+
B�wR9/�H|���>=��b�ɿ+��M�����v�O�սμ��  ˱:����f��UWWUA�ݷ���윍g!$�R�H��ˮ=(l�Imt9��QR�i^Ӻr-l&ȉQ�8J��Ԗ�u}�;w�Nk�᳗޽z��ǎ>8�8��i�q�x��8�;q�q�q�N8㏎8㍸�8��q�8�q�q�t�8��8㎜q�q�|q�qӎ8�8��m�q��q�8�8��8�q�8�>8��8�8��8�q�t�8��8㎜q�>>>>:pq�q�q�q��q�8�N8�8�q�q�t�8��=��{}��O)�~�sD�.�N�*�v婷KU��.9���\�i��x��
���Dqs�z�	P�s�pZ��t��;uxb���J��=w˭ҥ�EY��ڎl�I㒅N���(��A�Tu����ܷ/(���I�t�	�*ҝ��Ӵr�/:�H]�2sb
��sj�#�N���WJs;�$��{+�0�<ōۛ���0���=9mR~���	KZʡ6�p�씈CGUg:�Cm��x곧�S����^v��%!��s�5�C%VN�B�>h�U�w�WUԷ%������^�d���M��gO32�!W����d���(X�[�P�Dx(�)xf�g��-=�_i��O1�]=�s2��������4�y֜i`;U�o�Z�ff���Τe�;����/�y���5lM�������{��d�_Z��W�9���u�6m���{�Ҷ�K�.(�>���ȭ����E�*��%20Q]��L�ꔫZ�ʾ
:1�P�k�]7z؁�P�i�y���͕8�Tmm ;h��'ʺ�-��	Ƣ�d��I�y�h\��j=B�[S�
k�(�6V��m��(�LĒ�Ɋr�{8Wp����7_����8��Ǯ8��q�q��q�N8�q�qǮ8�8�q�q�q�t�q�q�z�q�q�q�8�8�8��8�8���8�8�8�8�q�q�qێ8ێ1�q�8㍸���q�q�x�8�8�8��8�8�8��N�:|t�4�8�<q�8�8�=pq�q�q�q�q���q�8��eW�w���$�T�+����y޷]b��p�7��3���sb�����q�ut9��Q��/s���Mu+Sb
>��9��se�J��ISY�.r.�Go���+���:��H0��%�%^Դ�lz⼫��v�\���+�`fV�U�6&�� �<�^�j���U��4̋]��P�p�xyD8�.��3�-�j��'u��xVR�C1�z��/s����M�UY�
���s���͡��"-s���׭������/\�b�5�7���L�\kB6�.n�ذ%�Ɗ�6����z˹{{Z�&"ctR�M�$���(7�p�b�@k"����.N0*�_;�Wݮ��xx�Os
Ȳ��{\\�Viv���r�H�ѠB������ �ڕvh8n� H�{U�%B��e*�V��+s� Blt�sۆ0�ݧw� �<�Z�ǽ`�gQ\!S6�䆹y�8pԅI/�eu�a�.G� ��ѳ׼i]�{�)*B��^�[�]p�n.y����We.�`����,�fVq��z%��cT��X"[o['ë�ܥ�mr��qX�aƲ�gmii�J�3;%�
�����2�tzU1��4sLޕ5앆c��!*�5���J����w���L�N�t��x��8��q�qǎ8ӎ8��8��:q�q�q�88�8�<qƜq�|q�qӎ8�n8�8��i�q�x�q�q�z�4�8�<q�8�q���8�8�8��8�6�8��4�c�8�q�q���q�q���8�8�t��n8�8��q��q��q�8�6�8��q�8�8�\q�w����xe;]=�ץd�!(���Q�cEX����-ȭqd��\2.rk����`��w�u�J��Ѽt��7s#�1���i��KALǊ��]��v�d��NN\�x�ޜ�ų�n��S#z>����)՞g2��H��ƧP|pV�#��xU<�e:c�Yhˆ^]wwluܤ�cq��՜`�BA3�xwv�[{ε("�ݼ�b}+gc�Pu]��\ŗB���Ӯ��V�nX����p�s��(^ �Jr�;�f:S�Mv�f�"6��_4�h�:�Be�Fgt���=��E0ޛ:AR�_RĞ� ��`]�ޑR]g�)7�@���]�:�e��N�9�^Z ں�{��'N�f�������Y>����A�{x��I��X��V �0t����6���r��;��u蜥u�l��.ִ�z��>V���j�qV����A^.��g�T��;r��W\��͏��vF�E��3UÅq%e��K�li`�×�����+:��@W8�\����n�3ҷ�Z=�_l%N�ٵt�[��w`�$�:*."���ʊR�D��;w�W���*��vwn�}Z�][s�(�u��t��i:�]�YjN�}c����:z�/�����]���ùQK�]^�oR��]�YT��#C�-s:��ٳR�w��zmSn�x�W=m�1=]��ˁ5��݇/��T����r�E�p-��w5@��;�f�t\�����V�e:8C-j���$Tz��gu�m�b���uq��7���tYA�]l���Oj��"��[���.�AU�4oK���OT��u�A��|�l��R�	����lG�i⎳��p.�T���2���!�����фO/WK��*.o�X�[�3jy�j�um�SvN�M#��; ��Kz*�2�i]8��"�ح���#tε6WWm�9��ev����F��ŀ���k��f�c�W�hh�p�wB��a���V�W;Q�G�]��V��hH�ξx#��>��w �r�/��>+I���:���.{��Č�/���Z:�gJS�W�3�f=Y^�zoт����*�-a�r���%���$�o2Gf�%�hVA�G�O'�@�{��GC;N�ڮ�/������T�n��e'9l��^7�d*qu� j�ջ�]��n�q/i��E�j�k�u�2Sc���4��B,#�7PaT��mK�w�2�r���ͯ;������f�Z��V��qo�fl�I�yl]���Y{���
���i�h=�xy���eS�,\�._:!�!J����u��m���YIeS�:��Gvr��!qUk���jҒ�eR�U1tU�G�,s�	���W��]�hW:���z��KM�
�W���i�sj��:
fG�_uV
�M{��Wf�����*���4 �Q�m����^� ��% =V��<��f�w��Cy�Bצ�+��y����U{���Xn0E�چ��c��R�H�����Xd�L�
�*熮�W8����E:P����F9��Z  �'.�5�P1� >��j������z��}9<.�4�.�`�̛^���z61'�krY��'�NN��Ƶ
��WeR8%e�T5�b��*�4��J�,���7�v�:T��J�+�o^kBjY�1�ʘw�;���ᒸ�b��4�&������7Jh��[ƽ��8�Vj�={Є��ۖw<X���s�����f�ͰR�����U���a���ꪄd���w�yj9].<j��g7�kAL�*�M����)V��˗0Zee��w]_u�4�՚�xz|���%X������o�k�X����&���JE��	�ƕ�t�V-����5.��V���:UUV\�3lDKt��v��B��.Sԙx�v������^�� �3B�O���
N<6����\sfv0�vr;4���g-ʗ�y��!殨�=/��s{r�����!ux4)�EvP��,�}z�S���X�s5��DPu�%M�I;v�qB�r�څ� �K��shxz���}]�uw=X��kb����N�\'`�������,&��-J-�G�ssQ�����
���r����U+ɪ�IV�:N1_�v�r�;J��Nik��d⨏x�)b3�M�D�"kv����b$p���j�x�31�<���b��J����^��v(��MJ��ʔu���rF﫡]C�PY��T!!��=�r���)2�<��mb��V<Ӈ���>�u��;�Rdm*u��:�9M;�I��~���Ө,vG>�+��� e]1*��$�N���(Zإ0(+����{�s��ܸ�p���5Nz�.����W����)��5=(N.��*�p��"��N��ZU��uRU�������wP����&` �+��"�U�c���p�����y�lbU;]�]�S�si�1lxt���b��{(cWd�6w؄dc転�*���vh��t�E�Vu:�9mK�ʜH�\_�����{�c�h�-�u@N�$�k��r�y�*�MLѷn�f tu��۽����j����N��M����E7!���F1�/yۮׁ�:"Mn��xkg_5��<U�+��Ȳ������3��;�;S-j�nWM`�AYRU�%�7{U�*4qK8#��Q,�A]�>:%x ^��_YD���w����ڵ�LN�X�6,����Mt�R�ctg�	����j�˥� ��>�4c'f<5�v;�=�y�:pȥ��0nV�v��y4�β{j�U��=�;kb��48h��|˰l�����'�ɘ7I�^ͳ�51ww�`�����kd�������о���o�M��ۺ����y��)�h[��/to�g��<3��a]��uGQ��j:�S�n���(_L��v�N�N��Ub�ӈ�:cb$����&�[r��Bcy�Q2*�s�.�x�b�K]�T�q1X�r��tι^�ʶV���M����hL�Nk��i���#�WsT!tè��u(����P6�u��3������[R�c��=�ys��(�-�rD��hg���C�+z�k����:�w�V7�\N�W���
ݖ�����P�oNs�Y�SO�٠դ��NޟZ�3�Hl�������,�9�� ��fԅ�is}H�T]�<�����X�u^��]573�.�o�Y�%�+C�R���fa̐����u�#�,ܘ��|i>��q١�t�;f�vb��;�d|i��U��t{w_�>�f��4<Vh$1������^9j�=s_Q�=�)ي۽�%���gwW��4�ݤ8V�ӱ�R�h����	ݥ���pj��ɋw-ӫ̉��K�&�x��j^�a"n�{��}Z�����\EpF�	t"ؐ�[�Wk����<�v��<��d��P襣������m��`Q��w��V��b�K����B�������k���*̦�T97������R�Uӏ�q�vT0":��]�͝$�(o��hW3a]�>�1�� a�Uz2�7oC�S��!;�f����K �V�ҕt��
�2��M)�b�:rt��-�/G\}t^ۃyj�ԧ[�]�8��Ub��b��i��
�b��q�9rG`�
�v[�t���sv�[T/�Rü�GZ.5ʶ�aE�|^.�,ҳ���S��b�f�l���ɋ�����/jY��`z{��S�ݤ�=��R��%�x� ;y��j�w`�[/TW�nB͓�c�9��6�b�����c� copu�!���aL��L��r�{�I�ӽ��[0��C�\�or�ʾ���TI'8���y�7��f ����0�yZ]����s��F�7������;{e��8�{iEfR�Z�o��ոd�;�M	�n�E���s�<�E�-\!s䌶��SV�>*�3B�[�8���R�0��^8�h�88@rԳo�>�.`��\a�Ρ�����[j���U��Y���u�����e`�.f/7+@۱,��#��`e<ɸ����x�e]���RU'����:qf/.���4mK˾��I���u�����
6�C-Dp�r搨��LA��Mr�ժ���Y����41e�=*�<0Ő���UG޷`���iY�[�"�Dg?f�rf��;*��Թ2ռ7��vpW%O�<t�1��������w�u�
�l�Ę':$�WV�^%A����kJ�};(�	t�,�zoj�^M��FIm&��7r�=���H�5��$P�kJF��S�3xqv�fk���oV�5��n�+���n��f���2�t΢�i6{\�/2��t8�鷰ӝ�x��1ĵݗW�\+é��CC���T�Ǘ����~�������Q�v �[�S�FDU�C�>b�mpi�V�:-2N�v_R�K^��Q����*��<:�%-J�O��s"�l�[��o+��W���19{w�+:��lL��..��M�5�;���?�� ��2��ߣ�G���⿤��~~��_�_�BbM�J)	Q?EG�R�.�UL&��2 ��.���|D00�I��p� ��e E�M��t �H$��1djDAE�Aa�Y��`��1R� m�R�-B#��)���"�8Z�4�0��Q�%���&�a(cT�
M|\s��FH i	�H�
�D�N1�`�!�P�&�!��
$��I�u8�P�p��i��X$�� ��I$Jr"��"�g�%�!�E|D��Q1&cp�L�����H��] �H?%0OR��F����TO��,?���;����B��L��
c��\�6���utYƆ� ڧ4%os&���Iv�9�\�_J�#'�9:����� �y�$�ҩ�<9^ٮ��1�u������'qۼ�c�-��%�;ŝvh���w��֕.�t3e���8h�{[8ımp����[;����5�n�7[�y�<�c�j�# kij�_r:t�X�6!2=V�F���U[��Ǝ8���3��������]Q������$���k �>��¢�칺@s�];��j���&)�\+o� e�
]�c����3��켫~��R���\�fn��w�AO��[��L��v�K�s�3+�ڡSuy0�U��1�m��Y�>�ݮw��\��I�r�Åc����7�Z	�Jjb�w-���b��l� �l�	3r��a�͞7�as�I��X۝�9�0<�Ǖt��e�R�˝�n��f��8��c�1�ܘ�,Ps����ٹqD�Yw��ɢ���u�2�A>��ݸ�[���1�d��6�\%uE�r�(�ョd�h�b@gM��ֹJ�H��'���ΔuGE�t*�N��́#mN/�w�Ȼ2�̰I4JE�q�lF�b�6"P"*�J$�¢����)��Rap/�(�"�S��Qa�"14\(����j"$	ϊA��i�XP>h'(�Z�D���H��J�iӅCe��B�2C��,�Z1�`2�_2��$)РRPI#�"T�'F�T��ĵE2�%�H%�"F4�d8R	3 pE!BeH��"�N}
L�d3!0��� j6'��Um��(\�Fbe�K��d���(ϤdC)1>��JT�$$-I��i�XP>P����MDD�8
A��	HX%B#O�.��(�%��)	e?�L��.CEDL8\A�F�-����"hN6Cm�SqC$-I!	���eP��(�>re4 -"J�4[��LH�M�/�"L��a����Q��h	1����i'Љ)�� r!7>A2�I�̑#P�ّ 4ʢ�4�"�K�#��H��7
uJE�AbQ���ʍ ���T�MBYM9�#�`RB��ċ�肤k��@�E�z#���p��q�������iN�ɷYG�@���Bmӷo�=}q�qǯ^�|q�N�7�!�P$��jTg8��&]��:es��
�$$a$�56��8��q�q�z��㎚t�f�j1���I�vZuf,�_s��^jdF�l։�6�Ԍ���ӎ8���=q�q�z��㎝6���!�K!0��l���&�Q&��V�P};��5�bw'NF�A�+n�{����;�:Cmy�q�o0���v�Ou���{��o=�kT��5q����I�Vog��׳&�n�7���u�uy{�'-���{��2{���l3��u��KG��R��Rr|�	����E�RY!/���n��>��㯌�K����w㳫�k�y{w]�M�o<��WBGu{ׯC9���yz۷T �9|����Y���]t�R��5v��zi�ݱ��{�����>z�w��v���[tj���I�g���SJd|��7���r�om������^�O��%�Ȳ|ݽ+�u�j��j3U�G5֞�=�k5�����f��{�k���\���X�6��i�5�k�������ޗŝ����M��%,Ӂ�$��G@�� ��x�D���6�ۻR��/R(��mo-J=����i�9��޲(G�|�w�������{ɾ|�M��.'#.2�L��AA>�R)	H��%6O�D!�8Xn�QB�?RAg&O�[��L���)<3���vSm�<f�#z�r-�{�)p`��uV[������ӊ^�t��(�]c���mͳ!� J@��j"�P�"d%,O� �[�$P3�Ț
|\BA2�$A 6��I#m�q�������R&�O���\F0Le2	$'$���%�&1�`��a�f���|��/{����Kٔ��	B�*�,U\��܏�|9��_?wu��~��<V2��߭n�Cf�u��nN7�W��=�{"��GR�`�F䁷sSO�^���rB��խ�t4mF�z�dҏ'k�����	RE2*f7Z(�w�["��\����[T�@�Hۥb�#�oΉ�U��is�2ͦ�M�QQ��[��ES�Ũoj�,�
�X�·V���7>�A�qQ��u���2��IڣyH�*��&���K��6��_�Y�:�X�ҟo�z��/���[I!i}����d4{a���JJ�Y��EP��ɕ�Q�,�Ti��[��� ���*�� ��gl���y��U�/3J'8S%�y�17��jN�}x���KJ&`�K�V+I1{|h-E�Y:���j�ҧ���	C��]T���X�;��f���ge�'.�L82�$;��Ֆ8��@;��A���ۡ-c�+����
�
\Ol��w���3��\��!ٚ��)�+�!`��N�R�N��J�x8�ϒv�v�é��`�툰�Գ�j��T|�qbrZ�\�������Hs-x��*�������6�6^ܨ!��Fߙ�&{
� �p�g����/���[b�d��T��Yg�2�٫���F�c4 \X�xThE����K��Ⱦ#���I>-o]�X7��>L�N����8f+��뿩/n'��!0�U�yM����^���U)�^�oV>^�oeK�~V>�e���X=��h��V&4Z�U,v؋���ǈT
�)+i���M�z�����,Ԇ�=
������5m�D*Z�! vP�I��Ա��I�哳s��j��7��fmE�u��Ǖ� �	����1�I���i0N�AP��˽�W4� ƫބ�o�Cv��%��21Z�L��[�&�ड�$���m�.�}��[�$�i��ۢ�#i���-��) QH6ʔ�gr�C^��{��G�z��,r����w��jʛ��R.oM�9�Gk-+\�\h�zL��\�V*Q�w6_�O��0B�.�P��>z��zV
4�x��͟�κ�7�X�F}����/�&��f9�b�t���XԀ���������0�X��_���羯����,���`={Y�3�ij�U�(�li1A�'l�ٴ31��ǟSC�X;��!�d��e���w�^h��
�s�朅�(2:�i���X���k�֗|VL�D��Qד]�"�6M��wU��;��F����3��0t1�Fly�Jc#�4k��)���+���ָx�O�#�ؑ��̃(�����`8�SL��Z���͢������'vdib����E�ʁ���T�����k��E��L��`*����ړx��
d��bL�1�Qy(�^��[��{-V�hg���KD��yz�5�^ �#V�/f�-\�s诱>�ukew!*��N��A�}�^.@4�f"����}��r)��M��WV�H��⺌���C����}k�����|d��;\�	�՞�>��&͎�+5v؀hv�]Ie5��I%�s�F#��Q���WDte\���%��{k2�\��7+;��7��T�WX��<�=�}K6�r���]�p�3'�[X��rT=�3Mq\��a�z�M5VW\L� ~ ���6��4���uJ=G��K˜��>��ªC�0�H�CS�I�U޽�/[����M%*�lώ��٧����@�^Q��5��'%��Q��xI�k[�Ζ�T�*�ϗ.�b�� �*4e��>��7A�19���!#m�!��ؑ%�ևGi6�I}�$Ḅ)��B�ϓl�A VzF߲�Q0�W���^R��Qݴ5[�ge�	B�-
}�+`Y��׸���̼]ؾ|D&�/ϗ�IV�cĐQO��q�\09���ĭ;5km[˵
�T��lC*��=�הVgW�L��@k+�����������M�����xkK-vb�k�C�wek�>,�ň���s�*��6�b��֢���q�B��e�_����q���Le���g+LY;�Ä��8��"������l4����Sk�����u�m��;~�$����e�����w��N�aRK6�9�g���5K���y�%n�ס�^S�&��Jr��)/@���4�*�d<�U�:�p=q�J�n2w��8���ݧ�*����
��K�ψNѠᷮ���k��H��N����}i������Y	"��4��F��;=ָJD�R2���l�xA�H93CD��r���	���U�U�CpNM�fOR�9A}AWф��,��:�ֳ�m��2�p�CV�%��G���}����zJbjZ�C͜�msF>$id�S����D`���/Y�5�KkZA����2K"	��g�w��z�O�=�jZ��[˲���kM�׀Ό':3a�wBN����:�;�
ʗ����Ji)U�F��n�(��\�LȜ�&P�#��@
*���*���75�yh��ݼ��N�/��m���tR}��ǣ�q46�N�$��D��r�m;kv�t��a�`��թ)m���]­pj]\y�&,5�4�0Бs��m�m��k��nRT1J �m�>�vI�!�7���a7>�3�k�����f.�,�]��X���ԭ怜sc�v�;3����T���2[�+S�%��hF�l(�����{�!U��V�Iu�
��&�����,snpa=|3��غ�w[���u�*mj��0��7�m�,����{'w7��̋�'#cKyz�t$L�-O��n6Ck;k�ʻ���#.�S�<�fI�]#'�����KQ)n������2u9��\�g�胰�a�k�&m�b T67wR��XC31��LɎ�FMbFJ����6�����= �CM8��u���,�qbԶ�R�B"�e��߲���ʍ��~�N�����]�{����Ǵ�������Y"J6cix�`��8NbL��8힄ńc�
�k��vX4�ݬY��Y�]�*d�5-׽�	iq�#`����zc��R����~�����}�H�W��g�����c�mEo�kR۩���(eۭ;,�PU%~��/i-�����U�3O��0ۥGK�֣/�)�{o��.����UU��U��Qe��i���P۶C6^��r�r�P�ٽ��`���:��ֵ�V;	������>�u�P~>�>�u��U�>�Я�cJu�mU�M�/N��u%Ѹ.9��ֽ��C��9P\|��K�������xy7wy5�ݤ�@����u��lG8�� �����\WK)�v[�S�3�S��H��[8<
p/XZ�Jg�n����Nb�-f׺my�Ţp��yջ�x0�4�$|�oK �U^}�t�uz���n&˕Y-�'L �M���ݔ��1ESl����>kk�nK��4푉�ҲO�:�؊.�X�0%le��6�l��!i}ݕ�����]�5�Nm�
i�S�Y��,�R�|[on��[bh��4��MB����UUIXsV�8�l�砣ٲ#�L���) df�V�1��R�R�D��6w4� ����z�F@##�>�Q��l��:�/qp����`$�f9�%�ٴٓ�����;�|���ZֶX��!,�����L� 2�������ӒH��Q`^ί���B� B���d�k��Yk�!^șU��j�ܯ����S��;oZ��X�m�vEk�{��Y�ض�D��H2�*$N\"y��s�k*����|K�m0�v�냯��3�|4%pz�j�\��\z�s���u��I��*�^���x��Hѭ��{�f9|�vsV�V����ͿA"E��TrZ�����W�CE��
K4�\����3ȼ$�0�Yqx���c�d-�
hd�/2��*�"���5�P�E��eĢm�E��3�HLnI�؅�H+گC�*d����Z�d��֤��O6�6N�37su1��l�L�n�n��(Ic���p7�T����;�Y�r�U�9��/ײ���UW�ϩ)T!l�۹٧�4�VZ�+a�޴�MI�U[��;�T��il�ɨ���k;z��KR)�3��v�!�)]��hL�!Z��U5;贵�q���ǐh�� �$�%��!�����4�hn���I�ܭA���"���"خ�W��m��/�E�*�uL���ͼ�L��� �쉨-o��,n!l�1��p!��[3w��ý5X�g\��]�}zi`o�������*�ν�5�*��Vӭ��J�e�0��H ��O�� $�J@/.붭˚��a�0��6۷���G�3o�VT�;���g�p����:�����ȉ5�sK��w��Ha{�x�|@>>�!w3.�ɪa��њ����=ٶ[�HU� ��:�q�ݻ��m\>;ǰݝSa�ۻw`o���v�E�$���턝�)�[0L|���a��i���';WaFO�.��?4�ef3h_��Y^6�����>���8�������E ³f+�Z�]k0dR�zQ2|�z�`²��l��"ӪeP�� ���K�������85ue���c�zO��66^�9�N=fZ�JK�Ղp�`תh6G�2��{�7!�P��G5�\*L� ̓��!u�t_���tA �,����7����y�k��m%m.�z^�}ϬnĤ4�s�mV4o��Z *f񇤪�-�s%6�L�nAeŭ��^�ZS�G�O��1o`�����.A��|-Q�w���0�i
>%c!o�5���X7�W���ӧ?`��1�j���)��N�TZr7U�j�K`�0i���Y�UXٸP:��I�*���E�7��㜸��T�� z��v
*bLl�r�>�V��i�ᯰԩ��!Ц�o�'�X-Mχ��n2�S~̴
Ė�-��aQ`�M�3Z7�v�ԏ�e�y��T�v�V'�7ͳ��	
A�}F������+���T<<<��L����>�^p��/�{%}���˦�75�[	�*��/��E:[��ocң&�)�zi�@�(ۥ:F��l=B9���6e���Ͼ{�/\�����<>��J[ke��O�?���up��HvǦj�;���d�E���GI�t)��W+X�}y5Z��r������}�H�O�;��j�$���B��n6S�	mNS�z#�}��~�}�Q$Q��"�*���X�-�W��sE�/+u�uy	�3�jI�|E|���|Oҥ�"�,(����v�jɘ�֓$��[�M�����槎|�r��y_es}�����kٿ��������ޕ�&�N����]�]�__���l�c�N/��5�jI���g;ȴ`� ܓ�#kh3�vpF���|��{�{�&��;�E��l��/?ZU�8��aP�P���Wf��*f��u��Q����9�,.ב"�TLtҌS���R�:T2��:	�m;I���{tK�v�巁��"�$��W�t"֕H5q�'e(:�wX2��{�9�y�Vo[�z���.tr�KX��K�����ƛ�D��Y���t,^�U��7Y{:����\�N}�)�#��\� �r�\k"pʏ)p�D��6�H����7��Jż�aޮ�K]��A����b�Y0`�v��z���f�Ls�N8����"T���֛�����Ds$�\�r�m$ZU#`z�.V�B�|z�..]fQ�<�ڳc�J�`
��s*��#���:�����w���ma�(S3�[{1j�����z���kym`jn��4�d�R�]5
C�Fm���ګ�ɂ�ҶC�#��e)gl�����t�|�H9;�x���m�޾��Vp�[U���0:�.���ַr�v����پ,V{yE[V��#ڂo�5v@)g]�P4rL��ɏ7��>`�����*ͳ]]��$�\�G5+QF�jf�2l8X5��
7V�\�����0&U'�B�@)����ڹ{.�,i���2rGT�m�9RH���x����}�u��B�K��C3+�䀏UZ��a��6UN�d�׏ț%����&)@ƭ%s��언���l�D,��e���^���Y,<��mu��T�U8Ԉ?5ĊL��E2�M~�_��r��_\g��<�e��-O���3Յ�w}��褪��$'����[�㕗���\��x��7eg\�iRUs��mG]w��������K�Q��r�L��c��:%{!��@���k�pcg6��N�rt뫏�*_t�A`�f��µ<��������4v�ю�n*����oҩ��^wW!���Bq!�L�]��퓳����t�gm'ܹ��7g9SP,m�{[�pS|Ǘ1�����af�3!��v��n�ު�k���u�[�^&�j�ޚ¬�YL<��E)+Դ3F�&�/,J�/�+��N��\�]7��nWc���^��B`O�X��އ�sW��aŌj�f�:�_3����{L3.7��J�Y�U�3�5�~ D�����2���Y�1⋤ʻc�,�(�D\+w����ڔ�tf�4�6s9���iːh���!��ஹ���Ev�r����e�odz6��������t��a���^V����lQ'\v>4p�Շ�*VoZ|�Ϊ@�v�ť�Aބ���x����#�%β,�;kg"C��j�77D\)�*��3��W$([��c�yH���ܾO� 76��.�U�y_G;�����P���[���;ﵵZ��z�փ�Z���o��5|a#�����m	K���۾�z��EȅUM�}}}}v�_\q�z�����>�v�폞$MJ�T���HFY'}03%9љ$�J�$���@�;�Fu��۷�o���qǯ<}}}v�n�4I!�#�g���'9�Iߚ��/�o/mÀs��+r[P I.����r0��Ǐ���������=z�����n�<����-�p���~�dw�d_��G��%��~t����]}Z|Ŷ�m���������|�sY+�@�p{�Жh)~m��!9��6���;�:{V�[X��#���6��^�ke��Џ�����Z-�i�f3�J;9��&թ�Nsn+{gyI��l"Rp%ed<�XvM��m�$��NlݺA&�7)���t��^}|�֑�Okr�~�=-�����q�9!h��N��j')�k&��ϙ�ֹ7��A^����/j�L���C����O�ז�����?5�侕��}>{����n�[c&��y"RD�H$�D @ d��|[�c���y:��N^Tbv��@�m\�����ǳ/��O�a��}wy���g/w7\�<�&�F�hh)���<��ݸD%� &S�6����{����sL�4�y����v��E���@k"Y��[/b���b�m�^��x`o	n�Hބ�\
��[�^H�4\Q����&{$!@��y�^����2G�������_!��{��6���C>�-R�0tx1����Lzȧ�=��B�s=(7.�oh��0J}�0��7�f��<ɝ�~S�ޛh
����>����`��R�� ��J��y��'��zmꝥ���1t�o{�^���D��<�R0qP�V�UZ%���	�v��;�������8������A'�	 "A?	����ˇ�����٩�.4�1O˔����@����P�1��l�Des�?���N7Z���4�;��� Ǟp��D�t���O�����J~�wO�0����mbH��ƸsF=����;�+T7]6�l:�!����ip���_[÷���M*�|u s.�r���U��jJ1<=h��-ƓF�O>i�<<=yyR�T�=Ԕ�Y��fx����� t�~��"� -"�t;��y7O��97�w���=�����1�ׁ]�4�4ǂЬ����:�A}�����f�P�~���;�_�u�nd�D���g���N,姥M���w�b]�[c�G	�Uv(2�����f̛V�<�CmL6���J�]e��s$�[r%��k�\6�jAM�6#��E�!����R�Ju#�ff���P� �~���0b��n��|�{�}W2�&]|>{}���]��C�kga]��|�^�:c���<@�Y��fx	���Z�LK���x ,�S�2qIxɇ�W#�j�cK`5�@F�vhp k�Z���R��v2�l���V18xp�6ǅ܊��j�~G^b��g����ue�������h!���}03n��KV
��R;�
X���	�C���mH�2k��y��7� S@YIQi	ͺj	�����=�[el\Z5ڻ��Y��!���Ɇ�Gc�	�n��7JAc}J.T;&I�ft���~�W���r��vY��"]���8����c#�<��+��͂�
:wD�����7uG����ĸcA��# վ�s�ǐ����:�~�( ڳ����Aud��V~��2��U�����c�q�pb�����~�A[��
���`��W�/���Ѫ���)��~T�Gn[��vcO�b9=��4���g5���������>�{�
��B��w>��%xy���ZꞫ�K+�|����� ./q[sM��ё���`ʽ|P���,(��_Y�k�����z��9�GO�� Ɏ�u�3;:�b�u���{�+�ҧ9�F0�aճe���m���Ղ���<.�f��0T�UR]��N�3g��vzQWs����A}�buNtpH��]�ڜ��}X�Ʉp�',�Ɍ�Dq�\�Gvh3�	YP�T���>>>
t辜꺫�T����]Fk[[۽9�!u��q�*m�t�-�V��xA��3L掏����|���h]���̆�%���ds�2"{}���J:W8�4[mҞ�і�m�8����v_W�x~c��>�t=K	E�͡�z��.�d�wd�i�i���)�N^]Lj��5��A��|w���h���߻��1A�邔��]x|9?����{4�X��Y��<�T�g���|5�M��Ⱥ�09��<�oP��pq0��f�/�A�U�u�b}V���j9�^o���i�ω�fV�W�ڙ�j����	�{��a#��#r�mͷӰ�\�J�^0֬p8KͿT� ��ҏs&���Síz�
mi/N�3�b���B�Eޮ��� x0t��~n�_�F0�9�+�D���
3��\�=2PXv�kC�]��*�\D����xx&Ըa���3�����vn��Ioi��m��׿��������Sٴ�
�S��k�`t�:��`��������R�]��'�PZ&��~}"Y�3�>;�K���l�x����W��=��oE1���GKKG�H�'�B�(Դ�Aӳ�佡���	І���+��|��t���ge��6�����u�ɭ�m�5	+�g6�S�kL���hW��)X��	��O�}�z�Ѳ}W�Rm���Z�q�{��9��b��ۡ���"
q�Bz7�ogp�=�s�ü�e������y�Bj�JHx&f2a7����������D	���&w�a��c(��ge@8-Ơڠ�w��\���	��ZW�Uh5j˻y��g3�ޫܟ
ʼ�q���f,��,ZY�]77m=U���'_%���L�<Mc��t]�cߥ�mH����;����
�R���g�ɜl� ��N{�*x��1L�<-�s�v_9�Տ��#��������~Wd$Ӵ['���Tq����3y�78��L�b��|5^|�:�F�����ӭO�%0�,[Lê�h=�y��w�I�:�7��MQ˨]��kf>��}k�@~hy{ˀP��L����$����k����)����U�����������=����R�z�w�b�?��DscX���c�`�]�t�x|���
�):/)���Sr~�1�n��@�S�C�mxw��6�3�O_<��s��1m����jD����)2�E�]p��4�-^�Җ�A/O&�ڟN�i�}�1������h��4�֘x���1a��^�B׊��{.�{��X��ٰ_4	ܻ���)�4�j8�sOe%G�Y&d��^R�Q��Zλ3�c���n����/U(����A//�*��pY|s�,���P������Yʩ���$88"F��v���c
J�b��o���-��z�����滙&s���3�v�ϑR@1�a?���@F����b֙�AN��o
�=<^cj�3+��ԯ�Q]�	t�K��G�S�c�P�c��IU�/�9h	\t{�.��v:�L����'�h��=R/�Le��p.���έ9ܸ �� �	X5��ݿy℟ &@-i�b��L\MŏB����;�g{����p6�/��D���ng@4.�E�&��� j��ΟQ��5���w�6��"�}A;u�͐�d�Ól'���Iׂ"<�,����`SX+u����=0��}�Ҋ��X|�>���EN�r�wsk���6S	�됅R]�ͻl7���YV���{�����i��(S!���O\�DǠ��z�g8�ga�;u���ͨ�]��	|on�9A�6q>50��7Y�H��q"�$�T�<��x�����n�O5��F5�5���9(f��$Bb�:�1n����80c�M<&��3g�M���� "��W͜�5���e���_ l~	Ō1-���uler�U�q�=���n�!G���<���J��;XQ��r���,`3��'VN�7��h��/�[Vw�[rT�"��t^rV�Y 6^]@��S h:M���K���B�uF�z9^wMǹ��3��6"���;y�jM۹B�W^�й�������<<+��¶iK�}�xe.3�'X[{X!��/�̓ߜħ��Kq�wS����|r����~Q,0��7�l`���{���1��x\?3�`���k����Tt�.�Ȯ�r���L��s���櫳qx̶��.pY�����y]yr��=��@Ht�s6ȸ�Et Z�zt��}SL5�C���"!wFI��x_�������G��-���~P��D1�ݯ��۷�&m����*m5exj)�2�1����^<J�=- 0b�D?�������Q����_������]�m�9I��Ky�5�8�3�����G��x^EÂ5�O�LxN�)���J�R��U��>��nu [�z�>D�~��/�u>#a��'���?�'��~-��!�dl0m�6��ť�q��˳���buw����A�ơ7�-z��ϴ��ώO'#�Jh g��J�H�,�z�@>m�u���� ��D8���Dc;A
<!���0wVHlp ��V�"S�*�gwc_'h�O��ܫ+� ��xg���.S �>��e�[Қ��Vޚ����G��>۩޽~a����Y�3�o��	. Eg
JA�i�P�g��G��܏e��#[&��[
X
��a�?A/5dM{C,�s�������$❮)J��R�f8�p�hei�ǋF��Z�U1Ӕ�<��f�����d����4F��)�4���oy�0^òxK�<4{�p\���l�bHFk�9Wi�mӶ���=Z7���6�C�;����������g����l[�bOg�wē�=�>[1���ĴGd�<��p5���	��\�pY~���l�j���{6�G=#9����� X~/wC\7&ͨ�uע��x�om�ѐ�b��K���}'������A�똨u��r҉nG�ن $�h��w�!��+C�K8|�y�(��?���lIV�atʹL��p�����[W ��w�5�KnVtwxO���X�`�oB��p�w>o�b"�G6�>�0��Gr��v�!���S�6�r����%�|�a�o�8����X~p+$y{��5�})��e��f?O�9��Jl��b���QY�S�c��>��$�|w����cc;s��B>��&����ܳ�{�����S���ܟ��xsg&��bu�����(�������e�T� �}����T|�3,�5m�)O��+�U�"��h���	�qU�#��{r� ��&4�GF]��x�߀�l��<ǆ�� ��)�-.���B��h�V{��	�{`5����Å�p�nB��f�h[6K��F�'�oWo���
8�����FWMz�d})�єI�������� J�]�}�k�>��K�3.�n	f�噅з]ڹ���6���*v..�6�o�mW_|+0�_{����A��>1�4�QM1� ���л�`��>0�L)�G1��ejWj�\�根J.��������uh���z�穲���[7�ɓ�x1�>��<�@�4����� p23e���;�A��;Ou��3t��%�7��P���5�c�_���Y ]�����~7�[q��)h�/3�=���r�΍�%xR ��؝r����I���ȸ�t�`ח�G��>'a��m�Q���^h��ή�6�xl\��	j�
��=��o_� ��#��bg�,�s�@�bs���|�����9:W�`����ׄ���c���<5nA�=�c(Z4;���ߘS_RCh�ۼ�Cv�5w��1HR�1�C]
���^� wr��E�{AM��)�nA�֮}7�Z�Z���b+)�����������xa�LSz��)��-���Y�9z�����2|��O5����&	4�S�fL*����vh�Q:;�i����qv����̥e<:��8������o�Ӭ�,S-�Μ��W-$�z:�W�[1�d�5D��M���T�o8��uz��@���#>�>R��Z�ѻ��n2+�'���k<�z�w�)�jl��)BTp-Xv�Y�Ѣ�hv�W5��M�����I��,�a�np����F=Ö���V+��S�ݜ���۷�k��jv���۽�Qv��ݬ�{yv���W��9y��4i�)cJ�0P�9�3���>|B�0��*��:�J��b���e��K&�5�n���70b�\`{�[C{�XO�HR&U�%K�{3���ʕ�2o��}۰;�	<�3i��v��y7c���T	�l��6�Cv�0�g��5gw�,�� ǃ��A̪`sl����}����@Y�g=���O�C�.0��dԦٍ�u�֐WI����"�^l)>=���� XQu��W��xk3��7|L����}��8����^�p�T{�!]�0����b�����f��� �V\`C�W���?�����Sk�n��}�=?l����j�V�9G'�\�����U#(l^"M�
�$l�oP�^>h���B���C��w�$� �lǘ��:�OeG���W�-ް:��io3;"�P��*Ƀ'����	�x�П��߮=�c*y>�x��!��5��X�_��N�S��+5�-gWx	�gfxL;���ā�i����9+��!mc�9N�=�<:A�f<�?��f×]�X�s��I_x�0�������G2f����2�?{����o4_�l�xP1ݚ�7�c�r��X�V��bS�s�˵R�i)0E���S,�}_���z��9C*���0D2�꽯�"��4�Σ:E�ݶ��9\m���!���3��s*'�hA���&�Ә���967I�w ޻��es\����� )��hh\˫�'���I��n��)��<�#�Zxt��p?��b����|�xe)�u�Nt)����A�S�QG�v�d+�6g�Vpl�6ԁ,X^�@��L�ў�	?��O��Sk�=�8�3�$�W���8r����|@�/�y{��g�Wh
0
O���:<<�Ab%���+�&��^7�����\c���axd��˧�
����� ^������\&���fP��+�h�����&�<4H} "���+\����P��^6l��rᰣ켘-K��.�
^!�8�@P-�B�o4ÀK:�pXt��'�FT�;'�+��`/���e�-��1�Uw���׈gy���w{�,'i�e�T��-�g�|�痄�N�]	�� ���53���|����HQ���^Q@����@�!��� ?��5|G؞����5��Ty�w��+'��
�^nn�\�:q/�JJ�"/�؅��!��@)'=Xa�FVSm�noM��L.:`K gg����+�%�� X�n�X�2�mH3A���>5o�dH2�T�M|��C0�~�~}Ӯ+�n-�>�Z��a8fo={J[����dl`f?ٯ�Μ
�
N�����z90[4��f��;��v��OL�\9�#z���I�d<*�e��BD.�Ohݷ������n�d�-�]��{�N�#tTΊ���/L��Ï$j�j�ٹ��!K
��,����`{[�^����)#���� �%�;&�.ȼ�V`�n�ݗ:���:�Je�˻ו��O���X!��fj��o1r�}���ے��W���M�����x��{n�vR�i��U5'�CB�4k�oSqIg)�[V�5b�ڍ���1\u~���6T�i�t/!Bv2{8Jt�e)]���v�.�7n+.λ���1X~�,���:�=���8�ks��э�ǳW>�fY�!�Ҭ�6��O8��{{�m�<���S���t��R�
��5�/J����[����ͮ�j�ʎ�B�޽�r�1�Z�����C���1wb׃mډi�Wx3!<.a'������kݻ�� J.��S�}�J�d�oR�G��)���;1�.T�t�]O����N��%M�)��n
���;�gI����z6=�,�����3E��rޅ7n^��Wh:�*\5���K|���t��U�D5\IU��X��J�vX!�\��.U��T�ċ�@��"��LN��C�I&;J�R����vBb�g��hq���Ф�[�B�R£N�n8o��(��d�\�D\umNcဓ�8'� ȕ2�,��eBsh�������i�>9|�%$����D9�;0�/k�]7fn229Y:gt���t�D`�y,����,)�GH�b���Dh'�����\�[������8^��JG9�Ys�o
#7^4�5�e���
�m0$u;��9IiŨ�K�5�5x�{:�LK�(V�eT��`O��`yQ�;ҵL4lKv�U��p]��W�X9�z0����)L�J�h�ټ�%�g>*���bUqΒj��it-��d���Еux<��.�G�*V�ˤ���~(��gf��m�㔮g8�4*�D�N9�����s;����׵���G�[rdn��,M�;��Sؠ��k.U��s.SW�jR)rX]FNFW#�I�Fٓ

	�w�+��4�N�jl����&n�7������t$�r��D�;y9����ݎ���o���@v��=d��:J9���c; 7�ȩ!�,MH�x��X7^i��Z"��GS�,���%V��c�r\�U���E��,�}����ೆ�]��lŤ㽸�e��ky�B���s��%>��fa����꙱��:�ٛ�+��)S�+�]$T�VJ]��v�S�꾎rX��_]�~�������~п2����l�����D�HAK��Ξ��B�J� ��p����]8����Ǯ4��������ǎ>��v���wj_L�В�ۂw�J��ɫ��yh�������I���^>�x���o������8�㏯�ݻm.��@��%2|[�񓜯�b��ܜ��n$	$!ĸnHO�������m�___\qǯ_]�v��B]S(���r9	�|ZE���z�JI%$��jĒ������p���8p�~mP�Bs���!$��9N%yݔ$}���Xs�p���N�$D��9;��(�B(��âH$�����ӄR8K�RW���s�$GK����#��_�$�p�q���6\���8���D	85����8����q~���8C��v�'8�$����e���c)6D-A��p�$E2R���1� 1��h��ʅ�Bۍ���Al�U�r'e՝�l�n��������t���h�Ԟ��uI�f��!�v�\B�5�1�l;�	��
�`�S�����7 j4�$ƾm��,�$�B@a��I��i� P�PfD�iH��J6B-$�F9S�AA�SPB��&)EI���a�"e��d"�M6�q��~U��A-�4�SC@�44������͑����f�׹ܛ
�Θ3G��F�2)�:���L��6cU���Nq SM~A����DA{wS�������W�{���:���(4@�o�����sz�Ntʂ��k ��`�bk ����%۟-@���ϻ�h5�r����t�T��& 0�v+���#c�x��t�~D{�L���Q|�#��r�،u��d� ��9[�����%�ue��{�G�֞�]�؝�m��~���vDI� ��$riQw��������W<����0n����S�5� z����pm��O�� [9�'�x��	}��$���+v}��k�#9r�٭�^�-�l�p1MV�?�nG�]q��w)�i���?X01��S�y�,d�(�&ˇ�=��{� ��2� ;c��6�z��	�8�%�l� q71P��󻪯��U��Mkm���x�pb�C�B� '�V|e��������n�g�W_����|L՝/M�~��˝�{�5t�_ܥ��m{�VQ��@^?1��]}�w�ϐ��3叛��8	�%�H�v��4z�N�:>� M��Q��º6q��z-�i�5�C�&���t��X�����僩��7I��f`&_.�s�����3��\��!�:W�^�S�Z�Te�rc����BB���0ğ��wU>G��	���d�z�k�t�;)^:��]�A�jJ���qk� g��빼�QknP�����сA\�*�-�Ui�����u����=v=��	���5�6����r�u�2{��Z6*3�^���{����Wޮ3�D{�U����/8�x���9%�ە r{�N���ï���t��ݕ�}M� O�f{��i�P�P
�fi<�/�XqM��/M�}"z���^� "�֪;��� J*�����܀�m�-6��ּ'o0�koM�ܞ��Fǁ78��S37Zay����7�Z�}�m�>_A���j��Sۧ���K�|�|
�k�D�S�޴�x��7�~N����zk�Y3��7��e�÷n@ƭ~�?P��l�_�e&��W�>G�������#tf��I���7���,��S4F��f@�[�v�Li�#|���( ���0��]h�u_�(����;cs��@�e��LU(��������ʁ�HƆ�jP��P���so�S�z�WU�3����?w�(|P������!Y�	}K�H��t��#��i�P��f��ր�e֩��d�gbxW!8w�z��@kY�jzҵ�Uܠ�Pw�c�1�H��ph��8B�ݢh5��a����wkkF�&�)G�*�V�"5r���q���Q��`fa�!���/�xfn����I"�ޡ��y�X4��B<�X�j��b����n������6�	��6ɨ:QmJ��;�L2�f������z���ХAX��(�T�R�����O���ht��Ȣ�j�h]?�AU9ձ���gt�m�!�����G�Dn(�����e^�{i÷�{a�1P�)���c`N��o�mݣ'���%��~�3���7�r��b�H����-T��K;l�X�Ϻ�7���8{-�ڭv�U�G-n���Bi�\���/&��eO]��s�~��!e�{������T�g{w��;[{h��
�\�ߦ�t����r�Ã���<���CG;x��BW��ߘ���?ޤK����xχH�I䘤���P����ʟ��+tǛ�Fz���"�*�C}����������^9`F<vlτ��oC	8���,:M9�Mc�-�2�%Y5�{��x�z�fժ7;a��D3x��������>����E��0��*��C�Y��΂��v��]��x�32L�u�Z�� �4��?���֖4u�����7�Ey�ϲ�^��].����_����s�/at$�/~�
�G+�`Y>� ��5�:�"q��J��Z��8'j�?8DFg-��CD0D�}���<�3��.�u�����՝]�#��_b�Ab��aHƧ�T���HQ!?�;���b�G�����}�^#sF+�jh�/�YL]��l&3����}w2w���
���)�w����~���
hhPXY�qQѼ���{6)��H�cy�������/����lq��X���F�A3�};�
,KfN8��>6�ץ۟&�3\���m��zX���k��� �oPg�;�u��D.���b	G׬�e�dü��q11�����rC��l�]'H8+�H���]����)��vy�;�����t��8S�����M4Ǔ�8Tދw�y>���3oԘ<�#͎���C_=��P�Gw=��j��+^��T?Yg��_Xza����퉿O���S�8�����pض��Fn�A�(��L��ٳ��1ퟤυ;Ň�pG5��g�>�"'=}�y4jԉ����s���k�3�����<��-�4c1�[�dH���c�\�wtJOBE+1�=�F �c�ݯGl@V��#�
��?r�n�2�i�Ƕ�������i:�N4��G����������.��O�c�D�Q���̓�Ĭ�v�����64G`;��{��
�N��ظuF���c�C�]_�Xv9�Muw>:�e�[�j~1�m�tZѲ��̲�6����t�L9W�2��[�7�3����p��V;Rc���2�]�1��|=���f�P$�^�V��JS�̋��������]v"����]�6wfC.*��{[Rn�>^��c\n�����_�����hhUi��E
���A�����MP��qi�6�4b��;XU7�E�{�cJ�T-36��`��Ȫ�4^���{��P�OO�G�v-��p����u��O���[{;�y<�}=}��{C��n�_��=��v���f�������h���)�o4���\�/ͮXGR��%k��콡TW���(���t<A3�s㸀�&)YD1�?�@B��|<��t�{�����7v��{Z� Cz��J���-�`�j�%%��*����^z����.-�@�`ƫv�<7]��:�����i�C�~�}l���Oa�,,�-��w)�P��V�s_���?�X���`�eS��Q.9�uC������C�$�%z�k:F�$�a��i�P�Mn��7���@��R�ә'{[��Az���:gk��C�u��	���� �o5ST�=u5W^���{����
�a ��/��elI�a!�g�8�σ��H�x�S��e�⠗m�3�^!�׸E�P���p�q��P�/�|增{d3`N"xE��u�r>�uw=�{r{��z[�Jtk�|�aZN��A�����Y�kW���OVbX*,3��{�ެ�NI�������,�T�K/zؕ�u�d������W��(X�BslF�����y���uk�l,�[ty���P�5�"�>��q̬;�ٳ���t/�7s�z��7��8*��ột3�/��ki{�������T
hh�d߽���Ή��г�5v����9����y���G\ځ,�#X�v�(8�_�
Z��c�|�� O�<���@������'��
{a0
��P�+K3��ki�=�=S;/qa�w9R�X�ex.��>�u���CE/x��Z��O�p��`��;!�UpXOI��d'�\�l�������/����[��T|:x�_�"�ڍ��O�2��!�ws�^�J�����$�8(}Ͱ���\"�vi7�8����^�-Cv���TSr~�1�@4��ב�/A�6�57)�Ύ�8���"s(�(�V�0�wq1Gp-C�%��p�s
�Y�^�j��wBeC��a����	h#�8)�=g�{�_��W�Z��B��_����*A���Zw�G��t�n����b�r(C�TX᧜����^�c�P�\>��!��S2�c��Z�]@Ĕ�Q�/k�_?P�-���s6����$�Tsڍl�p���5��Las�����=#�����{����(:!�\4ݻ�Nz��3gHسSZ�ng��˹/$vxQ�aMGT��}Ii[��˳�s�NL6;'&�T�e�w'J�n�Պ<ۖ���p �4fu!�N▮*wm[�73����X^��v�}(����@���B�DE}�;7�y�>t�vYt;���+�/c�CNBTJ�	�%��6C6���Ds�a3��HY��	S�����oy�v|�)�k�r]���P!h�eF��ֿLCpPrJN���rfDg����"�p�=�gݱ�HWn�
s��TJR�!h�mg^}.Q�*wP���ŧonC�L���������/����`B/[��O\�+Q����*$Ӧ<�Z�o��nZ 3�ۦ�|��U��+B����WU�������I�[fi�l��F�Z�ݾ�ϱ3^����Tƥ�y�f��ޱb�s�@���٫��?}�=?'���4O�ӣ�PҬ��rc�����Q�y��3���fRf�+(��3�!��{ϧ��?fp�ѱهt�����%�����1<�`wJa�^�]B�����G�g������]דg]>{SG�o�"�+p7���V@B�z�y:�c��\�;]P�y_��������~�E�.��e�h��olw,\:g�dt�$�LS��ʧ��2����r��C�L6�߼��VJ�n���v%�C��}W�Z]q�T�YmثfʓjYӖH��$�Q��rݐ�wt#G��=o1��A�o�fZM���Ӳ[���/�Mg�b'm�0b����W���`��P{���i"��9�/��?��H����Jhh����o/��f}�G�8�U���ǁ��C�9f|%��)2�=s��n��A��v�I;���]&��Ĵ��>h�?7��x`i�z�zF�c�����cu\ݖWk�o_(~�Sb����1�w�$ȫu�Ťg����/ص����wRZ�Z�<�lOomᆜm�xZ��.��z��q�UR�l��S�l�p�"���v|d+;kSq淖�vjO"�Sul��1��Tz-�%~���7 ��������f��-�͏�l��~��&��.��n�j;��x����^:����ŝ����q>U�����G�4�4Wz~�յ���w�Z�K!4���(H8G�����ήm�̭�='x�}ɨB�}m�\�8S�a����G� sԽ[ұ��thB���ݶ�.Dnv�[��;��᝸0P͚��V�I�W���!a[�.؏�}S˵�PR�5��[p7}B�B��ӌ9��e͋�χ��6
���!e�^�~�i���0C{��d(��9��,�u�1^����7rX�X�ǫb������-��H��٥k"��AU���V1�#�^�,W�G)�W�e���/��e5�����	ãc���ò�'K�g^�ܺ=�vt����)�wUk62A�< q�EhiPi��DSw����=��Ծ5��]��d�ʭڷ1��b���̐��y&��C`7]B�tl��3.T�ɞ�����e��އ�H#<�����ܧ1��-z/d�fё�{��̎���uh��"%�Ȉ�>쀦� ��z�[���4�`O*�m��d�b�.��'������1���Џ�W�mqy���ֹ(��M��7'�%��r݅����_��眂e��Ƚk&<ŕ�b�kA���"���Os�c��-�J�sU$H�C�whvx��#�m�W^]I�jJ1=��pc�xy��C��'A�a�O{�/O2��wm�u���st��|���i��S�� #u�(@��|>� G��y�Dke
��q�}�ܮ����b[w:D��k������sώ�%>�pb,�=�_�摻v9w��9�=m#G�����9>ɕ��n�y
�cx��s�UR2�-�F7Z�h�����x�S�@���!���G���K�d�Ԋ�1%��m��v��g<�Ԁ��iJa8:���{)N��A��_d	�2��
�t馡���#哞��y �!���n�_2?<��\�8�I�p[�J�;saS>}�Ts����	|*���~vgҦ\ʰ~{�2-oeU��<G�(#�����P�Q�ipy���R^�`f�*��(�^��+s��܍'?�/C&���e�Vj��zu��{��_�� �C@#M ���;}ɽ{ـ�|us�O�:��΅A ��O��E��u���O�`d��Ӳ�39�O�U2x�1�;6}-�IC�ʝ�%,�`SV�+0d&<e�[���J��k7N��W�cw�J�����yO�ٖ�EF�����84�2�Z���­����j�����O{�ד�Ȱ�p������QM�?��!�R��W�Pc����$�<�P�zy�f�k���;�C�@:�C��E���\�A�涠7!������~��g�d���̋B�W����ۺ�w���#��_c�1_Y	�=PyY�Z�|o��}=��w�m�/��^u��۹�׶ލ��9J#x>�Ut�5����v�*�C���OOA��0/���4rߎ�{.vֶP�a�SH���~;�,��9��=�G(��qk��0q�~?V������`y{�F�Se\�f(�����X�J��|�4S���~��	��1�~���YB��X�����}��kC;s]ֶWF��G�.�9�k�n��M��J��g��n���iɧ�Q�/��6�x	����F}��o�n��`��`i7�;j��r�iᕪ�y1�J�wt�Fvu´i��%��;��*�ܕ]8F�w|��]*�+�J�Z�/��e��;H��7�,�c�P���N����`,6��(rD�d����|:����+���ޗx�K����:gq�o�ˠ�u��6dci�����lǤ���s3t:��e����Um��e�Ӫ�:��aۈ%�)�^�\s�#��2iR��CN�^V	�r��Y]X��Mv�mA'n����<{ǲی ����]����JB���J�ٵL��<ౡ�MA-��t5.W҅e���Y����:�vQn�S^^%���Y׃@ft[1�Wn]���;���K��������dpX�Edٴ)��m)��D ��}]�S�"��3����\�@Mͼ��{g3\�@�0�kOU��|4uȚ�,-��Rх!J�(���|&��M2ŋ��݉�xQ�]�j4��V�\o;��6�����=�0�L���(h��l0�-1��W-z�n�m핌�;�܇X���w�{��d��mue뭘kR��n��Rt��.j`�vV��Z�FX*7����݈|=��K��ب>�y��1Z����kKo/���8W'�alTA!J����kK(����T5:��B��%8��E��^+k�G@�BDU�g�=�T�w���0�B��С���ޖ�M�y��$?rD�CF�Y쏴�|?|v�O�W˴E���Ӊ���ʏ�P������1�h�^��W��4΍y�]��Ѓ��}�c���z�[��NQ a�a��Er��������\���+���C��ݚ{mN�&uA�|uu=�p��AtcU8�c�%بW]T��ջ�X��9����z��0�b�0�u3(#��7�z�����,��Z�9Eܑ�n�}$�����X=ԪLf$�g�k:"��#��{�e:|3�c��F���&����X
VZ�t4��V�Q��t��fu��������׶��C�#J�	�vP���WC���F�ǂ;t�q+�E��N1��:�_v�*��s�o��m���#�[�da$�s�{�ެ�ϵ�IY	\����+�ۭim�=�kCx��6�@[]Q	�`�]��E��wS�oq�>0:%�Yر�M�δk���G�uݽL��I��p���QY�\BK��A�Z�Y�rpf�o�-�tK���p�oB�)ݭ��i�Ȯ��V��<�w�ʘ�fΜ54����2��Y���6H[R'��w���v�Ni�q�����n �we�.SjM)�z9j��9�{2��7f��L��xZ�%M�nfk��Z�&j��ɨhZ
���E7(�'Ҵ�k�`s�S�u�;�Z:_۪���D B����z����q�}}q��}}v��e�	!$��"I��^�8��y�%��pq$$�!�~w�z��㷏\m�q��q����n�y%�wHpq�?���qGG��N9H��#��>���Ǐ\q��q��8���}���8�ԗ��GEs������OŸ\!r"R���I[K��������JpR?�; {ap�s�m�	�c�;��~��)\������;�~l��כ洈���G����' P'')��NN�r���8���i:�jq���O��I������8�S���]���P�pS��'q�-���#����S�u���s�t�͉)
ΰ98�8�ֱ8����2s�Js~�P�9_-����Ýd9�97��>�nOo��V�����Þ��Y��*y�O+��}���ҋQ44*��� "�߾�w��߿7����m	�>|O-̴z��B���aUfQxj�{���2�*����Owj����Y3���y�J��ߘ?Hx權uu��$�igZa��7L�G2V��~u}��[��?<1/ A^�!�1�8v�c��\���U�oP�|Ç��}2��Go�9�)��PXv������V��+�>ɦ�\���7wu˞ف��yQ��Ϯ�Ȱ��i�S��dk%�Jz���fq�@Y��A	��پmn�}y��=��K�3U�Ql�ϝ�ή`T�'�yC2ׯ#hyef���yw����/�j41��=��x@��ʃU��Vw��H�T^�$�
��IJ]�����l������=��1��I��+^�d	JZ�cNdQxj܄���.�F5VmZ�aԁg��"�IY�������Mm�T������i�T֖W��xyT�W"eH���m6������ȉ�������L�ԃ.�AP*�K=�vq����u^ئ~-�s�v�r�{n�j�����]i�oe*�P�c�fԃ	Өp��(o,�y&6M�]F�\�ue�yj���T�%����E<�ޓ5����j��-B㗱��*Ы�I���N�Ԁ������}����mE]�}"2*[�������33�U��9,� �_�� ���
"	DU��o�+����u�l>���-)	���P�{ye
F3�@�����gi��i��qЉz�{O}���A�|CE(Ɨ�'���'���0�^�]B�<��
�1Y^Tm()��Kم�a\uQx�p_y��Q�u_VTc��1�=@�b����\�y���wus
l����ֆ�3���a�i�%��p��n�6�`�G7	<���_*�O��)�5+��Uݘ�]�y��à���,]D�K$v}ϖ���������ܮ�3�~{������m��͢�{۽��.�^uƽ*^؏s�h&�h�����|���94�-r��CzA�
�6_x��q��z�������c�9�I?�q����zH�� ���s/zq�+��d�e�3Z��8	�,g�7���)��BOr��T��[�5x�^o������Y�o[�G�/4iiD�[�(�U�~�4�_�����¤zu�9m[r$�v<y�v����C�8�7 `<���_�M���!���mg��}a��E���>��Q����Ŵ�N�t�e�9cpL�_�=v��u���"ٗ&}������%���	�R���5t�5urvb�1<YRc�y�v]E��C�q%������t�U��y�5)z�.u1\�W
λ��� ����V�
hhG��{�.r|�~���^){�������,�ir^�[N�Y.��3%�@���zr�G���I�.�������������oi�l$���Y��>4@r��w��!tV��{����)}ģ^��
�A:-�G��\U��!��)e�C�t;T�����À���٩�]Z]&s��Jv�g������T_�f����x4�U�ұ����d��sd��t[m�YL�Y������}�RN�uv�"8A�|�{=�d4G�~1霋a�C�>ԄsU�g�sU�O?r�a�F3�i�<K`�衖ȩl�5�<�K!X!}_�P� '�Ǡ���/� ���ʽpB�4�~�T+'X!6�����9s7��+6��xR��a�>�t�~�a^��!
��//ѭ��1)��1bU�]�^��OE>��m���� �9�Ǡ'����Cu��Xt����-��V�槃�Y��Z��9�y��冱���<�l|�9�`Bm�����Wl�"��^^��j�����[HܟO2������7H!�K��t3U��_����h}j�ˌE�����O�f�6�~��4�軈B�Dz0�3��ɏ��f]�ߣXYv��u)s7�vG�7�j�b�(�79RB�i�}2�e۩��)c�,����c�-�f�����a��Xc��q�4�_���f�\ד�|�o���i���G�?�����W�;̸���ړ�%D����P�[:^jԎn�\���!/D��/��;:V�.T�Y-gNj���<���!y��C�Cn����d�s��2y���ʦ_7,CU'T�&'��Zz�K�k�A�{�4|��_G�������4���R3��E��s�mP�׽S� ��~�����a# �A�A�³ܑt�C�zd��"�rRHT]�i�u2*��t=��E���3L�w��M!=qǆ|J5��
^��#>��ǆ��:�0Z$���nX$�%:چdҔ3QU���o�R���֜�p�H�f���ηI�5�fz���}m�7�=ɑ�� $���x˲mj�-�5��:
o���m��4>ջ=�o�J<��7�LB�C�Hc�m��kr���R���ӨjG�����Ӿ��a�<��L�"���r��<�l����}A��7q���&���}FԚ;>��~�Pu�%�Ms'>�`����B���|�|pb�k��71�3�I��'�{DL�ߋ�+��3/������d��O%��:1�ݒN�5�m$;,��"vs��s���������'���.�o{a���x=)�{�ݻ{}�-�9O&�R��\����A����d���$���҃���i��E$@�'w<��֘�gv�&��P����=N��ؚ���{g��]
E��s�[���=Yr� ,W�2����l��~u��w*��)�-��r-��c{=!������[3m���k�hᢞ�{C�ɏ���s(���2+������y��v���������ik�ƪ��GF+n�>�Ȉ9�D�����Rz}��m��'�b-#k����<�n�V�al�ĉ�}^.�/���S>;��w��'}fQw�=Z��{Й\?>���Uv�lB�=��s�9�2:RB�+^K��C�k����5��
љ%8�	u&R(=0:TZ�6�zwO&S�]k		ױ���$� A�8r�#˧n1�� �� ����$�G^i�,���N+-��Г�XP�Hnu������f!�Las�۞c��3�ՙկj��#i���omK�H8z�x�(��)�^�@����Lv�C�%��������܂���ޑ� �-\���Y&�]�G�\���:wI���ȘΞ��'�x5�.���3N����ȱ5�%e$S_��p�x�}�dT��}�n�s�Q�W� C�@�D��t�4��zInE������o���\v�>ӂR�v��FkQ�,�}�*���"SV�+��;7�5�^ϰ	��4�SCJ�4<�x{ވ�Y& �g;��A@��ּ��=�@>}s���BB�`Q;�3V���,/FG6��;����cS������I���	^ğx;�
׼��Uj��6.�u3C8�v���5+�~��3%��0gv|}o����{�t7~v\��C��{����'�bv� N�-*r����+���ƭe^JV8|ض0�>��v|(p�yt�A�[��Y��=��^j���Ke�>�Zс��_u
���w_8��ZfR���U���c��,S���F8&��gg�-��l}�6��0���)�5G.�v#g1������Slb�$5d�h��¬k����S�8M¶���3��3��1,��q�M����aϙ�6����V�d���e�fz�K���.b9��^+��-��t�<LR~o�S��)�ج��ay=�:b�[V�{���VP�}��]5�HU�X-��߃�ʏ���"̉T�'���1���_.er��)~[�Z�G{��,yĴ��Ƽ�����>/���x�@�U8+�WU��U��;b��d�S���.N�#�T~�)�+7���l��z_�i:y��.��$���2�
!�7qHV�C��E����ջ}f��|�2mc�h��b�݂Ў�i�[���vw�]��{�yy�Wa>�v� SCJ4�����A��r�ث�?�J�"�m4����+$�z�a��19JS�kk�6�GI�
m�O�G�O?��.���֪�����n���>T��0��O��k��Tv�����s5�P㵃T�n�ȈkQv��a����9/R�:�GUH�b�l������4�4t�����-�l�7�y�H�^(��\��G��=������,��O�'-�nEmq,�)����$���>�L}�������a���ߺ����D��:�����,�ݾ��G���}kO�)�UJg+����H���O���wS��+;s����yp�2�yC�>���@����-�S���Q��epx0����sM�}�QU�S92��m=�<%RE��ᴺ�%�{Lh��٩	x蝹KL��=0Ύ��*6P���U2��[=v�y��ښ�x[{�9����̈́��p�;�P\�~^���x�K�g˄��J�#{��x�ϒ�
n������E�*�=w����x0��_D��(�1���<'В�s�	���C�>�7�X�as	y��q��Aq^��:��int6�k�.-�Uۿ3�7��A�rs��9��3�QQ��"���o>�m-�>�/�5.�E�μ�_E5ԛ~������2�Ulc!=V%Ve���Oa	�:ok�6�z<��[L&ݮ1֨nk�^��x���L�����(����iZhi�q��{h�JJ�;}~c��}��)J�5����Q��*}�0P��G�̓�R�UϮ��7f������Mk��<��A���y���p�k_��s�R�yP��󅻁�!j7x�Nr�4�a��w7k��ظ˸1���'��3Z`Z¨�����߶1����G1�lh�@�wf��p��5�WAi����T_9�n�ZGiyH�0�L3�^�c�8X��Y���������H���|b[+p��]���毤�zt���1<=z$�d����&�r9gc;F<6Y�x�jA1y��'/&V����!C�2y���>|��vP5����dAa�Þ� �WB��Y���p�_`�/^��t0[��Mv^�K��8v^�}��=��d�Yh}>A���d0 V�"W�L��p���Gː^A�9��b���m�'4��./�c��û��;���><T�&S�zQ|`��Z�[^kWUU{�F�v��C�_P�1)�vd�;0'��o4�t)�I�.��!��I�IR�3�z��p��뽕q�2�5R�e�K�����,@����,+:v���W{��ӽj��|حE������	�ٱ�ʲ�dR�{�Ϋ=�N��C$�Q�w�{(V���ht�ˋ[�W�kv\-�ve���V���G�H��д��
��`y���U��[����t� q�$w�\��?��*�
~�|�1F�t�5�^�yǅ3��g���٣a��"Ғ�܁���7x�.�k+�E�Pק���!c�,2j�x5w)��;�:l�ʲ8��s�����cW��&,k|�5v������/<�l�q�u5���H������l�%���ųl�=+\d<���n���H��+枩��������<˃�xf�-'h"��f-�����:~�I�� �N5Qp�Ol���<�x���1�ET��jӋ���&�b��-���9�{�~�R9z:{�]����M���l�Ø)J��d�ͣ���}��[M��=\�	���<����@���+�Dw�n�L{׹3����S{X? ��@�,dD5�C*1��_�V9/-���JL��n��i��FS���) UV/�#Vm�����H
/��3�����ò��m r��yjU�\���ժ�-	�u[�C	}8�9��7̟Ϲ,x�)�ꝃf�oP��w��+Md�O>������<�M.�eᐦ:�%j<�bٸ]�z��ɚ�;�jJ]��ײ��`��ֺѬڀ��,lH���m�]�����c�o]�q;�7]�W
�5]:��9Y;�TEu�ss9<��=����ڕ|��  ���
hi$�$Mg����{�u��`�ɇ���tٺ���ZM�.F8`�}l��'�0����� 佪W&�E��C��wP��$��[�.�I�T;=�Pũ���f@�÷�y�m9:�bc`��O��֪l�z����՗�P'+�P-+`&�L�J�r�S�ڭ�{S/T�T���`��������3VWJ`�禓�J��t��1h�d��Q�wZ|/R�%��V�R�<y�E�VENϻ|��v�/�n��|���w��pƅ�e������$�;w�"-�c�<6�@f<Ğ��߼����>�o���\W�s�m��ۍw+K|�DdP�����ot�`]m���W�Η��@`���<���{��"5䕭����I�M�JE�>����PT��p��<"q�]�tS�b�<�P{�\�<{�\�W�|�/��YY>|�>f������P�x�r5̿E�ռ55��応�i���+F�ӂ�Z�`S_D����)F3g-�LO?wB`�Ы��[�]�:�
����j��ƪ�5\ϔ���ԩ�K��Gf؉?��P��o3B�5Uj�0�LP�cۭx'F�2����/��nEI���cGf%�[L���v�]�ג.ʁx�:k��1m=S�o[�,�,��p�لm��h QVt�fE���@�C.�M6G\�݃-`��j���t��㽺��;��2�&���C�.�IM|��sh�ҳe5�8r�s��O�lw���dZ�Ў�f��ja���2+���ǖ�@�b��gy���|/�� �����;�y�<SWE};���Β�j^-���ֳ(���;����������C'��f/�a��X7�ei����̜�]�2]�e����N���n3c��ǘ��V��4f��8i�m}�0�8o1ʥ|z�6#����C�,�֝�q�+țsl���^b�B|�-H�ܦC}��b��i��\�w�49Ȳ43 a��`XL��`͚1<�����e_!Okﯘ<��a�ܱ���#Ͼ����7T��r`��S�Q�ӣGXb�G�V�[n����*����s�o���t�Q�R��*W9YzŮ���+�3R��v9���ݜ�?MS	3�w�lWD5l��}x��lh��Y�J�t�
33V!AL��h�(U]�n�bVyuwR@l�i�%R����t�v�\�XW[R��m��]:Z�Xb<�jP��M�*'
���D�	Th���Q�W���v�E�f��)�hw<��ʮ�q�yN^M�y��n�n)�5�y/��]r�wPٱ��Q��ۘ�+w�>���wp�7^�6�m�y1*
�b�*��!��\y�a2c�;ΆVZ�1Lͣ���ʳ��&��/���=�Zᗙo�%�R悪s��	�u�;�Е.��V��K�}}�v���>=�m�����Tw�󺼉�x��f�³,� !J�{��㏷Y�V�{��gTj��}`^Gr�!x�hy�g.=�wg�e'��2����o5�>��jf�����뫼��*@������f`���2v��=Η͓����:4+*�T�{һ-��EJ�+�.�N���w6�K��������r�k����JG1+��
䀪��H[Nw��[��t�+tp2�f��)LƾӨ2�ta�C��nK[��z-D�/���-���MԩJ���Ƅ�)h;��u���JU;�	�P���NI'�����\J�Ɍ*6xq�0Zؼ���\�u!�eeI�/��n���t�[�ެ�J+\m�� \�ܲ*_AW��]��������\��gS�B;����(_fj�Ֆ�;M_>�&�;ogTc;r�qX�H'�Om	#��v����TB1$�$dd�Pry!N;z�Ǎ�x��q��N8�o��ݻh���';��wC�GpI�BP�!��N�Io��__[x��|q�z��6���۶����PHBd�!9���a�p�~�*�>;���8$��u��1$$���_^<m��q�N8�ׯ�8��ݻj�$�$#.��"����
��
8��C�))(#��(�_�Q|v�Bt�DGQ�m8�+O�e�ީ�ptGƜ%��ݣ�7hS�'>���	L�qIq�\DQ�]9'}�\r�s����r�m���G;ls��$�8�rrI. ���p\����RqI^�{�nW�u�P������b��(�r+��ŔQ�u9y�q�I~>>��W���o��C�8���.22�E$�M�Q-H��2O͒���AI$�,�P���E���9[��lN�i�n��{�	�Ng>۶��x��Y6�c�f��R��9,sE%���8 ��S�S!P� 1�d"K��0�	�ARRL8�)$����`��D"�!RS�)"I�TaNI`�0��E���"&I|i#nKm2S�~���������������|��e���t"/�Z�1�d����ʝ����-�]����2r==*�l�~����a7��4'�^��P^�"�[#����.~��z�Y��o3�P�h��8��w)����o˃@v���H���,��7	<���<SWo�U}W8�h����tS� �4哸mvji���r#�hNPfj���a*D�c�eU.���3�/E^[$��y�"�.��-}Й?P幄2�}��765"5�c��c�D9��+��R��	�i��B쮥W�F�:��n��gU$�q�����O�/�pck�Ƴ�A^��+��p��P�C�6v�
���WO�g�W�k�>{�/��P&�[5����緮[ѽ�72{�P4|�`h�Z����잡�u�X�ϧ�JV��y�g4vG��1Z$�r��#���Q��a���P5��U�G����q�<�l�zZ��V�P���]9��+�ݘ�g�J|z��4,�!V�������`] ������W�-_�~x��6|f���U�ne�E��Շ���^Bנ�,���8y�����F��AF.�,5����x#{o�FG ��fY��h��ff�3���2�������L����d6���#o��eҾ�$���>ؽ@�|,�����n��h�t留����cGE��w�^L�[���#�q
st��+{7}ˆ��w\�<������������y銴���<3�_�)��l����&����Ԅ�wե�f�/�E��=0ΩO��}�)����'�瘭z�G��4�r�n�wӌ9��ew�,i���c�?%��!���wh"m��z��7��C�h!�=��%���l9T{x�<�{i�sg<c��q��[�1A�%�H�E�{����>;�!�2F�" $�}�;r5�_qcK-�D��V��9G�'�臨�ym�<�����i8:Ǌ��0
�$T,v��(M�Բ���;)�nt���1<������C�����q�"NE�����	��ơ=�$Fzm�}���+��������+���k�}�p{����:�e��EuwR`�=�OA�<��¸tx�V��K���S�j5I$t��1��}p#�E(-��C�Q|籺@�7�m ��	�0��O5r���b��/��"0|5h�4ϱ=N�Y�3;B�2x�Z����˷�]�s�ov�H��c/]c�A�y�[���;��_���.����ڐ���	>�LL�>��3����HOr�����_X�11�kP�{7WL�kz���N%�m�����rG��̧)È���`����u�'<ϽE�'�WQ��W�5O�7�9��Vws���������]�9&���]�&�cK5c]H��%stz�FX^��@S�4���M.��s�a�{����K��$R{����� �"}гR'���	}l��n/�t�[�]vO_k�q��~����~������W� ����4 V���TL�����s����e�C�&}�g)8��:��PJ�&����A ��O��?$�<ǂ�e�b���P&;i�	���C$69�S^l����d����;������ �tU��Pg��1C%�Y�6A���}1��=C�Z~�dz̈́���Pܟ�����p�� ~��W���Nm<.��bOdV}��-� �E���gͼێC&]q��Ժ���1{��_���l�G��,��λ���X��<1F��_E�F��X�f9���A����i�]:w}�;��qF���w�M�T:�����:/�:�>�8eh��[z�ʍW�|�#'^33��"�-{�����tt�C;�c�R{���r���W�
�|�xjܜjnF�h �x_]9�8N�x~׏1�li��&���1<�~�T:������:�|r-��N7����|Ȩ���÷Y�K�����o�<{J���X���o�i�r���ұ�F�j󋋶q�ygEsۆ���O�#�� ��$,W+��Ļ�W]]�Ĥ2�:-w'�5��vܻ�ޕ����]����Pf�m��[,R�m�l�n������<��&۴�g�.o�W�'!�5MF�>��$�W7c(ˁ�<�;��^s^�e�:6P�y�1U�`��\�G��|(��C~�B>��� Pܩ<�E7s�1���m��LV���;�ݾcth�۞�/��P�u/�t���Ųb���aƽ*D���'|rQyfxlȉ����L�ݥ�}��.�ʾ���ɤq�"F||s���Q@:�R��Z�*�a���g��_ޮo���>��]a�8`�'�+�p���
9�D�/�$L�kq�C6�4�j�۲(ц��q@g��t$��/>.;ì�N��J����(=�o�=z뽁eb'���n�|�k�
%g��
�@�揹W6�4�p@�bq�)�5�%�ϝ��	�'��i=�L�OG�a֜��� `<��$D�c��Lh���;6iΤ�J�ׯ%��P1�LvC����E>�jx��C���WTTK��`<����(:v}��$!v������ݸ�.��ھ��������쯦9I�P�>�<:Ğ�D���ӏ�L�(n՘>V�T�b�h4ح���p��Y�D�\��c�؍Ѭ���ȅk�î':�uk\��+��'�ͭ��e�E�ތ���P�a��/�V�+�.�f��:�:�焾��¯t|��2���΋����=v�m�����߫��y����YaǕl�ѹ�����b	9&c�nm޾&��IݛÇK�ïӎ�����U�B��^iw�Le����r��q�.���2���D2In�����ٜh[^(�o��z��$���͜a>��e[��f��8�y��o%�����C�ל|n42|���<֌nW�\���	�Ǡ-����1�u_Yu�IL�� űaw耏G�k�oF4����������Ú�������p���/��﹀W��4Q�T�!E�wW��Ӎ��ax��J�2�ic����L�F��⨨���mὴ�S��ᮢ��@���o64��e�`�I�d>��H��K�Ótn��<TG�mO@0
�h���6��6�a�7ë��B5�Le���K�
}9�3:�k���Iq �{��۔�o�7'M��Ɣ:j�O�3@F솏(`鱓��J�\�uT��s��6�I�g�����9�P�������澯y���߱�`���Pg_����E���oz�Г\/t����������g>��+k�د|��q_���9��u����<�rm�]'7F-+Z����ԫSz��.�yE��vg~9�6��t��b���̫�w��:�lz�{ژ��A3k��@$H$�O���I.�Sx��3�rnXb����٫�]�wt��x�ݠ�^��#hVi��Wy(�ڔ�����g���O�p�q� yj/��e�c�,޸�a�^�D�鶉�+]��7�<��.�N��V�s��dN��Nrnݹ�T
=�0J���H��W>.Z݁�<�Pᗮ�P��*���u�0���n< "�}�h�b��>�0�1�߃������xmk�t�wLS��R<xe�`�$�N|�8EC2O����CT>��?�|a�tG�����׵�y���ݯv5'��y���@����XhǮB���p��Q~�����8�9}������_-C�>ɞQ�C���wP8���F6��"�C��뀎��3%7���k���[�E_�
I���p��RB.}T:)�*����+�0r��@_D��'���Ƽ���9kr�[7��=�|�hZ�OUZ%xu��Ä\����\cC�\i�c��l��k����y<�'��~��u��B�t|`+�ퟞ����#�G3�s�=Y�37w�\��Bմ��/o_I���	�{�S��H����涿A��-��'%��y�(�da䥅�
�S�J�g��"0	��'�_v����D��j��#4"���F�־�fpU4,��1>=�3-�Xog:����^�$Ԃ��&^�z�T��U���M����X�9��u��ʛz�gt�����ĪU�^8���o߫���^o7��-�M��v�p����x�o��	����:�O2�e9漱�I�j���#�b��΃�ݭ|}����g{)��n���]��K��Ϡ �kp��6�3L0�)��q���s�|��C�'��P���*\9Y�=U��˛=OԎn���	t8�v��P&8P���m�u縐��I�^��dOc^�����D��?�5���k&;�*Ƙj���Wf�]����y'���yUH�-�@�`������̟���P[qE����B��kUU����zO �ݯ~\�R���寠���d����u_���;A�I�$���jh|̀x��pm��o���^�E�y>�iOA�c����0���/Erzu������蘬|��Hf��r�
bS��ɵ(f��U}���r��	ˉ��]�UN'�����B������0ߗs��w[W�)=vǇ��]�rKK��!���E��w=E�it��`%pk�`��8 �"��s�:_;�����v��3j5զ]��,uwPJ{\I�����t��R&K����f�ȡ�̄6�QO�2�}�3:e��8/c7�xw-ev1)����\�>+h��)r�;K&��r�n91,��"X�F/l�ɖ��x���HR�����
�� o舚�ݥ��l�]�kX01�<��x�g� ���S��DS�;�rʭ�~�Rn��C9�mk�#^��c���(8�@���0J��9��:�����GW�؅����i�U�����4\GV�_�+��ҘKX@��9��|��3�tށ�;)�"*!��\�t��3�a��0�ިM�/��K�s���C{������F�0�������/sp�ӸV�7���ǜ;pe�}%�4�0#vz��y���kfvg�k��W#w+8u̮	���G�~�x%���4yY���1A�tђӹRy�ynOӋ��O���\u��^�h,�$�t��=�sPo�����A檋�o�=۞"kz�Y��S!��������<���K�|�z�����D�ɤ��}Q!��㑱ͥ�^S��{��H�dDu,��Z�p�ۜN.��RaW�Ktߺ�XO�F6���\0d���+`��싍r�)uabE)loC
e���35�1%8���uΓ�t����:h�5� �u��6?�R99Gr��'擣��vt��a���]����@�yusY��Q�[].���%َ9�e�lSƻ��$X�����tHƾi���t/kH9[c���'z��Z}-a�T.v�deR#WC���9�|���R�%U������c0h�r�~���ɻtJ�CNo��dծ��6�1{J��Zuu`�Ћ�iË�� |JT+��*x��3;�df=[8�I�3�,��	�P]�����<��'�3�z���L�Ȍ
A7�[q��(,�m��o��,�S�JX���oe��㗲l��峇�b�Ņ���80.u"���w>�+�P�-埚3.qu�u�b�e�����͝}��F�vf'I��0J���WlF'�R�oL�\�8���1�23M��鸮xjY�y�: O�n5�g�Z��)�a�t/yy�c^n�뭔r#{f���=R)�T
m�!���x%+>l[
��w�ݙj�6%�ٓ��,N�Z8[q9�C��{eپ�f��v��n�}�+��YB�1��=Z��K�����{�����V�vg���i�!�	o�1<�~�Ø���1cw'��2�zu�xf��=Fc�/l��SۼHq�Ǒ���S�l(ǯ��<�G%1��r��.Vm\��i�m/��S]�I&�A�z��Qo�F��P��~�"c{�y�x5�ٌ�vW?�}�ͫˑO�C�$�R����r�U������v�J�GJ��HfZeG�����2�}H�v=�T���ෛ}S�N�PF�$��Z�J���n�W�o�j;�uj�ޫ�x�pr��C5����L�`�����=��ǟ�պ�[%ǜ��r+���0w\�~��)��r����預8���B��s��]�"�8���w	l�3�jW�Z��A�Ң��_��2�'ԥ�X�YC�f]t	Wu�4�pr�����+�$�Ly�>|J+˯��Zw��v
�M�����(�u�� M.�;qlsE�э[wϙ�9��B`e�G���lT&D�N�x�`UGk�r^���t�������fSӞnG�=���� ��t<�o܌����)E6��_�m1���Cs�eݛrn�%�{s����MQ�"K�n�8�f���DΪkNuTG˒�&��]�u7z2#ɡ��Z���"�۠��׏KJB�F�7��+�����#��0?'�Q��M��s�ڧ�o;`�1�e[i�l}�A!IR̛��"*q����C�j[�/jvqr|�Y7C�xi���"<�w=B+ٲ��`�%�^�)�/R���d��Ud��u�z��斒q|�bw��/V��7��8�7ӌ9�w,���G蝘�h_5U?�b�������3f_=���`���ɹT��]U�Z��ھt��pkafw;��5��kE1|Y����˚�l��wc��Cu�N�ܠ;�he����.�j۹݊麻�S9k���v"ewt���-����.̆���*W�;f:��3�V#N4'u������\,
�oG~)��4W7�sef���e/e��}�u�����;���������Pk�ɺn�;��mb�o�N3G�Gv^z���~�%5B^�*��Ԟ[��K+g
W��3�W�)���+�K4U��r�w���t�+���o���ɨM՜�o,q9�3�����%v�H� 
fVd]��>ϱ}��'3>�E:�OFwU2��p��wS-���٦aZ:p�q�;�n�
4w2<,f,l���)O��ܶ�&��WTþ�#a�}�ʾ��r�j�9���g+A�&���A$w.���K{q,2q��AA��M�&걜뫻1Cw�:��y+U�y��d��>��s����:���]��޼'�+��L.��g-��L��s9��������#�:m�T�����,J4̸���vD��Ԇ���1q��OzZ���5�h��_n�y�]�h�y-m��Ȃ�Ƹ��)�R8�C�����y�HЫ�V,˦��մ,�| A��a7Gv�d(⤲}[E9�.
̢L����!��x)Ԧ+>z����� �t%;xa�(�ʥ�,0ί���I�t��tx-�Ǌ�	��� �E�E7Q���Ewc�c��JG�x�����qCb�)�l㝚�_Y�OYR�w�����/�*�-�\��Ay�����a�9����47��ަ/��
f(�ܾx���Y�7)d�ΰ]��]�r��{}��;�sd�O��ը��%�c�����Tj�+�Uɗ��Y��֝�GlK4��w�Vv@�^���ѻ�]�Ax�����.���Z:���7@�&WRhJH+��3�D� j�P _;��B��8b������g;v�ŷ��yT/�:<���F��վ�j�v�_I�5w�3%�p;O��ݺ�4�Un�=�l�}/H���:e_#K/�{,����¤�¾����{QU��Qq�on�We�wB����,��u��5�����JY� È�_u��e�*5�v�ÝC$�����׎���)�Q�"ܚ7�:�ͻ]vn��r�{ ���9�Y�s{dY&@t��z���"e7u�1A�ы�MY�R�r��5�X�l�1���o2nܸ����Z�����hu�*��| ɣA��i��7�VM�x�xR�Vh죪�ݾ�#�������wr�U�[󒨪�꫑��'e�r���rU5��Wuu�!\��j����_NJ�d�Y��i��v�j������9����i9#�q�'��;����~-��Tq��׭�x�8��z���{��}��}��ƒ�:"�II)8��ώ�}�S�䨤�$�:�����O=q�8�^���O�;v�v�yN�.�I^���.I9��RH�U��ׯ_Zx��q�n8������۷l��D��A�������`��ڳ��L콫^V��C�Q�ݸ��s�y�/篾�^�oח�w+'ִN��BI'�tD��%�AD$w�v��~}z��M���C�g?���n�� ��]/n��O��G6���Iwwְ��]����Ϻ��9�9}j�+���t�����>�\w��>�сAA�m��������@ ���u.���^8�=:K�{�1��ޒܽޫ��Omtb�,9�gu�Ԙ[S]��;��k�u9�9W"����<�a���7xK]�v��d�����
�$�!e��.�@����KnG�y	�Fx73�m2|�s�籭�6t�w�S�l�⑔��p���������1�-��^�����ܔ2'B�8}�: bx�?;��i���\�Vy��򂕤���?��9�|��bdr��wn�qU5��<wx`�vO̓�xO�t�n�S�1�v�ȸ~�y�(�Q�h��Nk��Tf*6&%��o�z�T��2�S�g��˨�]a�������ן#Ιi�.�oI��&�>m���8��"9�zc�y��@����-��:O\�&��v���8�^e�X7wM�F���_����񿋌�,������ i�b���z	���A璮g`�ƺ�Fp��J��5)a�/�����^��^��v!��ܟ�~�.��#/�΃:�Zvq�%<�ߦ*v�9�Lh��g���ye�r�:ߨ}#6��9��mB�t@:vO��_[ʻm�s\���F:R���I�i��Q�����>�S:ҟ-���lc �0 W���}B��D>�gGG����[Nk�B�	��k!�f�\Xc ���%�Me�*��
�ϭǝ�y	�ݱۖ.�x
�]Uq�d��$ ��A4�b��[���Q>ʨcw;N9-d��e��}���	�N�Z�v�l��c����[O���j�s:�7���ԨW֟��hi���s�3�����Ҟ��䷜0`��cb~9=������Ҝ�iOA�F<3�`���I���o��93�
�V���x����,�P)�] �3&��À�E���-r�]�d�m�z���۝�w�H�?�g�׍���o˸8���ߨN�V��84^4ꭈ��/2n,�B�o����W/�-L��+��I�솭��S?Q�ǖ�]	8l���&�PיuF#sx�8�d�{$����
����q��g�.�B�Xv��j�Q��:osҫ��"l�PnԏSw��������Pw��%�[8x���U��..ްJ��>�����ԈmmO6d�^�4�p	���[�G� ���DG�� ��~n��=I�5rX��gB���	�84h�ߪ79��{_`T:O������w��I��zk�gwP�����F�0/�}ƚ�����ʹc���:�~`�����A��+�9����:�O�`��R���GO�z��^�g+<<�����s���0�<�c^91O,��꺚fr����#�'X��Y�m�mU��
���7x���m��F����/l�S�v��rV�v�^�mV
��K<�����4�.����a��&������K,�B�.˻���ǹqڬ��bR�Lԋm���'s9��j�������44�CC���Cu�'HK��Tm6�"����͚(՛��ewvYc$ylJi�V�|�<UU\�RSi�ޣ�w���g=�W�V�>Ab����߬>�52����M}��Boa�'���4��oC�=�-}Q�懼�{C��dE�ĸ�!Y�#��q�۝�>{�컻	��}*|���%�I���W�1�#�����kH�/N�3����aoW}���]�l:2����b�st�H�AD��椌�{��'���s�����+�Z�E��*���K�g������D;_�v�RaLs�A!��k�K�+aH-#{�[�U\���ȱ�\5�!��=!۸&��C	�����$����E�:��i��l�2���.���cO��x�cCX���ߝ5<= �sˁ������,�͖`TSXX�E���,������$-z�K�A����v�,����3�@��}B�?y<>F��s�m'�N띯��r���I�����i�[�������������Mlv��
������s�9�%w�|���<��y3e�>c9H��nA�ֲ�J��F/�l�º�+;-�5�W�$Ƀ�ZU���2�m-��Rёt�]�*YupHwY}U��+��H��q��e�f%��-�S�95O�U�ŉ�0�O'V�`v/@�im��ޚ�¬�����M(1�iN;� 쬧�7��ҷP��o"�.��G�o0��?��r��V�v�2�hb�5���z��~���W�֎� ���͜�&�,�
�<��dK>3��UXo� ~��ۙ��벼-U�e�-�4u�����|}�����^xb�	��\�}���v�$��u�-�Z�]���j��[�(�C��\hx�c?��@����{�P�c�X�nX��]I��ķ'�1M������绘筏@�
�߈��5�w��*��+}� ��Q��TW?3��{�� ���E7�Ak�t��k�SO�a���2x�՝�J$t��MP��P|��'��Rޚ�<��X��L�,G8��v�{�j��qW�fhKi%�������>�f���Mm����]�ԡ�[����^� �y����;S�û��K�S	��8F�����~S�nW�=B�צv�=���z�]�s�&{��*񧤝#�~lz���*#}�V�#`��v�h�����[_V�=��z�v����ܪ�-�{4�#��뼌�q�->[r$�v3��������Xy����pE~۶tݲ�l��f��4Xl[�ر{��fazف�.����	�����)a.��Kd6�����#>�b|�[��1]��m�=1�K�<�Z���F���ݨ�5,���_]��i��:z>��Fb���|���q��88�Yo��ܧ�����)��Ì�_���i$D1�&�t<���8�O���D������uzW��]A1}E᭑�2Cd�l�f�O^K�������Tǲ���D��At��kp4@����;��d�tbҎ��Uj�|�w[A�2t�7��#����A�Ь���Q��z��|錈�������w�����+��5n��q��O�~vsީ�wc�R���+���Ǫiu�e���[��}���˜VWu��[$1fX]���7]8�,��c�G5�`t2t�=x[TuNltv��1/	�S�)�{i����n(1pXp����{�{;�v�W����lW}al9'w݌���*%�:�����)�g��+��k�1CX{�=@z"髞(<s�Ø�;܀D��;<�	�=�1)���Suwus[X��q����A�+5�'��Z+s��L�ݙ�ﵣá�2�Ve@l*�@�o����.�t��(���a�V�&��N"q�7c�mw�>0��`���̡�1ˁ�+���rܞ�Q|���� �{ٮ�.�v�6q��)8b�|S��ww�]u���52

�Nm�p0�ow�u�S�k�}�Ӓ]}�؟i���|	�>W�Յ����sG���J����賺�cpkf��8��ijy�=�V����pk�x��7-���<�`��y�a"�Iv)tnW���������|!�\/ˠ���b�5�f'�N��/<4ݒ�Kϼ<�}w%���� 8u���/uq �SI����"y}�2����Ԃb�A���/��m+��\Mk�DT:�+$]�E<KUJM\/��F�f�U��ݨ�/��|���C�Ҍ�����.߬���u����Fy�{1A[����y����{�}U��\��A�沄d0 |z'}R��%�!�\!��bĎ�-�ؗ��K�>_@�rW=1vFi�y!bR[S�t���?���8M<Ў��W��u�� �hhZ��W�5-u���lLe�s�_n�ZP��Z��k�������aԁ�$="�++�%���_�����mQ�:��G��"/6Rz�]�Y�}VM���=���ᝲ�%�9h���6CW�0&)}<'+t}�bX�JR#y�>��-��L6�f{�/@���+�# ����}~�SPuRNưŅ�(���,�γ�����F�Tz�^�7��m��K����3�8����ld<<ţ]��'�\t����2ꑏ�����\9./i#OJ��x�Q�V 8��K��x�����ЮuX�8��;҆rE��x�To�C&��h����@rn�s#��=��r���+�Ζm�&ݷ8�t2���o{EۓN^��AZ��!�Ű�W��xxUW�T�Ͽ.U������W$��8J骩�VZ�F���S)�ʬ�R��v�i�p�Z��/��:�xl��Í��cq��z���tORijdr1��\?q�i�h��n�n]b��g��ޏ��P�~��pD
�l�=F�5�1=������Ņ�շ3.Kwߔ����ȏ��?4k��}�y��Ǘ��|ׁ�艇Az���=^=�n�NbT��S�wU��U1ݻ�5����!k����2��dNq�::�Q�Ć�^!ې�%�"�i�ȱ[�K'U�P#I�:��i�nO��4���6��/A���	Y~p�,ڙ����В�\��''�ͦ�q��7��G'��y�Dw8�*�H�<;���C��q��ͣ���׎�3�2��p���o����2hq�)�j]I��%�o���k>���0i-w������oP�:׈��s�v��S��&���=�$�3��:OM������c�V%����ŏ��BH� w�q������>ag��f7PX&���@�*A�+�����|$�~m���8�o���g�k@�c���`~!��學�Ĺ �z�CZ�� �I^�;�,�y>ʙo��Ɉ�E��f>ƕ��2Z�Pm�[(��F踯�frn_,٨�@T�5�~'�:ze����2���괶���ρ�)��Č5���u�3W+�ܺ���|�G������u��7�y���X˫�bX��A;�[�p:=��Y]SI�}�#�S5�`��q�h�(�� ����k<�3xpɄ�$�z���� �(�m�;yj� !��
���g+�0J��x;O-�Գ���g:��l��$v�_Y~.Z�V����L��=;�c��ݯ���Z���yז|��8���x����������U��^�F&y5��f���~�[AW�2���Ű�O���l|s[�o[=�ͫ��I�B�}c�bdg�].r��f�O>`H��6X�B��g��k�������zn[����Ve&n������#V��k�O�BB��iq��*��ƺaW���yN���jq@�k�J�ŷ�n��.�� ���=�<�-��$8���_+�`sEl,��ˮK�ն�1���fL��o��s�(����o�qb:���9��A��p7�8V�l������U������C\{O�x>�i}�N&���7*�O��1M�3�J��=p����'i#[��ae�m��p����09�mH�W<�H�w�=���_tU��T\�q]�@�\��v,;��]���ܫAmŉ{F��A�(�Yo�?��>�R��0v���*�Ͷ�˦o|���ǵ7ZH1U�>L8ঔ��Ӓ�&�ȱMgb-^����X9�p���[�;�r��j؝y�J��p=��{���u�$W߇���� j{�3�[��
`�v������!/-,=Lw�L�tL�q�Z]J��[����oeQ�h��lG���?s��7�K0l�)i�:�h-��<��!�2����������b�yL45��X�����L��v�=�c�1�1�
�Aޫh��6[��F2�;�Yl:}6'7��	�t�
�F?����"Az���y�5_�As��Q�7��IU�K��wǐ+��K��W�/��f02������i���V����1�jd��v���y���$�\�F5���ǖn��O��s��/�ʲCd�l�ٰ��B���|�q�k+�G7x��N��;����$��_�e�0[�5��Wo����	��B5Ip��RIZ%_�8����>��>�=�-3>�
b������B�Q�OG�` -����81���a��3���չP�j�tK��3�{�nt
xf��++��D�XB�X_�LUצz-�W�hT����j�ѽcQ5�Fx2j����9qA�z��xOS�B@��p&E�;��P˲�C��>����v�pu؛����Z��XW8:ww9�جJ�5��K��bM�M�>fb�Jd>�tȋ�u���Ye[�en7f�p.�4�η�;s/����`�gSt�W�r7��h�7�.k��2���{�yy�9��G��?P)��vN�.��C5����8��%�:�܄�T:>5�~y�B\i+z�+��vU%.3�1� V@BjO�� kлG.��wwUO��xY�~���pY�o�)d��!���~�1�~|ü���ǅ����H�0	��1�6ʔ�I�/u�E󞷻�+�&�}�#��v�����<�*��.�rӖhVu��[��o V<&�?�/1�4��c�p�`Dv�}��%��TTf�Λ6f�����L�8�Ѷ�ٷ�a��������q3�V�,aQ���:�^L���H��QAU�����>y�͏4���b�����"��J[ҧ��A��Q5AJ�ʯexm���X"¶��<Z�C,F��l��~�׏7f\�f�q!�eRAd����v�D1L�îs���z3wu�}\�~+�W�_�݃0�'��X��G�a&z�j�]��.E��Y|�؇N��nb�}MC���! �n�n�F�7w7�Թ��V�G_^�0r�����=ו���#�zW���;�Ǌ�o}��΋�l�a�a��׫uX4��s6�)T�|�켃�r��ˌ��ݓ�i��{�����ګ�a�e��'.�����7Y9ku��`�ts1ꅾ^��ѕ:�!�:F�8w6�� ���۫i��g5w}�塺�u��+�d,��ð���5���d�B�U���N�9E	�;w)>�s5䀎ȍCSRFwZ�k(Y\^PE�:�hYn3�n��.�0#d7:�8rw:�a��jY;62_<F�w�#���xtc��P����5,�ggt��s�U��ʂ����mP�K�j믺�r9"�'�����R�k�pB��M���QC|�Ap`M.ܡo<N��:�K7�Zq��x�2*�2�,	1h˧�C���@��,�F�Ǭ�KZ�b�ὫC`�'y��.�s�Ǧ�����3.�<--�i��[�z��."8�"����9.ڬ<ۨ]�N=K���o�M[���k�9tRh�S���2�����S��u����o����+����է��۩�T�g@��6I�.`���U�\B��#	�ݔ�_S���mZ�\�8���[��u�=Sf�[��p�2�,K��0�맸"�ڝ^��x�����;,u��bt)N�MRZv�I����b���q�Sv�v�[a�:�d�!���u�2�<����8f����+J�$�t�D[Y|N^�_1:����:�vn�nT�^cǫ�{s'\tp��ɤ�r>MbVY��/�՜����eoc���s��>!m@��+5]ۮ3z��̻M庵E����
�B����4.����cJ���m���X���{z�r�L���Xg�D1>˸�y#��)���F��c�V��U:�w��m�ޫdqO�X�r�����d��mu�n�Z��r�H�����e]w:���;(����,:R�WVw����A>�4om�މ��gR��uh+��P�fiQ�mQ��p;;��ųS���;�c�lq��z�Ayr��nѷD���d�}�x��R����<�ݖ�Vp�{�eX+%6o0@j<;;�1�ܝz���ۂ��1;�L�[҂T	6Uk��+VbH$,X�㫹K���Z���y���շJBrՄ	�`���c�N��s��ֻ�n�F���΀�j���S��e9us(&edǭ��΋[%�̾[�����B��(8+Xq����i�4޺�5�&4vd�gx${��V���7���#��]�3�4���;'7y�����9��`Hg߾���_i@�i:;����BD��|՗^��~w�c�;x��qێ=z��^:t黌W%~�n�.:�Q�K�^����I"Hm�����N�=q�v�^�}^:t����Oi*��R G���͎��m��wF��������;x�8�z�����ӧM�p�?5����h�#��.;+2lT�:˫�]��|�ͻ��)&ŗ�=�_��/�n�;��wߪĤ�}W{PBY�|ui�w۽�w�'v��;�hABW���N�+�9��n���g=l��8�;���j��6�|�ߞ�A����É�_�w���A_L�}���y�E��ʷ��ο.�A<E��-�&_�d*h }TW�UGĳ��%Dc�����`�ˍ4�&6p���!�)Y�,sM;
K�DU�4a
�X=o��3_M�xsf��a�y��1l��awPm޺������>_�r6�
(3(��Aҍ�R6�1ȃ%}b-��L�TIG!6c)�QE2�-�1dn6�r������H�bAF@�4�f"�p@B,8���DB���J"�R0��Db,E%���� ���s{��Q}3�v Ĉ��]϶f�\����ܻ�2�17�j�&��ޮF�R�<V2��Nˤ�2�y�^څ�@�U{!�|̷�vG4lp�}l�k7h�:|Z|��AH�y}F-ԍ�)�����qB��pЮCĐ˒2�I\�� Z��C����7��L��
�v��;���R�{���wF%7O�*�e�f��I�=y���Cu��B:b�4V���r�Q���3�0�C�B������c��E�u\�U
�z�Vc�&�]ʹ��.��&\����3
�Q�1�������Ă��pV�T뜗f����ڂd�����lTz;TH���t:�i�V7bx�@s�Q���g�q�ӡA�˟�*����k`;���E�9=�����72.��{���.RJC9vu``��a�k�7��/s�,OdnXʫ��9r5�u��꣜bE*��eh��zC��Xg�E;f��՟�;|w���A�^vX���V�˧��$S�WX3���%v���j'���������\h��@õ}F�+��-��Σcb�s�3���v�ο�>�\~���ص:StWF�J/�q�S)�8�WO����`wXe���y_6h����oe߻#��U�x�|O@�q��g�r���t�=Fv����È�f,�n��`Z��`�GW�ߗ%Y}G{{��S�~ 3�k��K0�u�֤	�q�[5����xva���.`����T�wdg'xkr�4���q{��VӁ��9�B��46���`�e��*)�����ot5Qtٍ����W!'����al�t�w��7�gC��y�
%u۵�:�����]�E��i�ϔh��0p��1SYY��2qd�`���Ej����X�޻\���D��SM��~U�6�Ցy͐�Pj�	[�;-��V�'��2za� M�uo����R�!#m6\;�,O�'ۮJ_�u��p���sz����Tuw)h�w����\��d�qݝ�n|�۹�����vLt�О�򌽶Pݷ��3�kd̹�և��������0�j�l/�Q�4���6�^���қ�x��-��{��+9��{�n. �uȼU���{huJ'���z��i�>#���:I�A�?���4J��A��}���=��,c��9�v��ߗ��K%M�u���K��˪�� ����t�P�n=��S�ß7K�@�:t0��o'�}��䣒��Wl�I.�?yb�Ǹ��Ϟ�a]<����]�9,��1����"�n�
J7O�����9_�<�H�FP���h�AM��k���v>!*ղ,\�9��ٹ5ǯ�+�������X�m('m�wgot��h�^a��b�~���v@�垻+��؝cy�gkf)ǁaXm(!R�w73����n7i�ǝy���ہ�cR��v�&zR܊�ޓu[�ꏎٕ���
�L܌�Wm�����t��y��%��^o/cL6$�_P4�/�+ON�Hǖ��dl��.�r.���k��9y[��8l�YP5Es\+���3�Y�<8'N�&Cf;S/@i���wϥXK�p]z�����.��E�7|�B
56%v���X2���c�a����|1�t	׻�
yA��u�Wq���9��-��ɖ�џm=�e;t�u�vQ�V���D7��̛=gB���8�Q���bQoU�gg���f���}�5�5��H-�����
O1�����x|�w�ˬ��ҫl ������̺��z��zЗ�z���^q�9�ԓl�h���; �k^����ƙi�|�酵څEM�J���q{��Γ3.��`P��˺�so�[�e�+�޹��^rg���4p�nF401���*8�'��҂��Hu���+�G2}sN�Paê7\7wftF\^�#�5��2�����nJK�q�3!kݾ��O���EkM�k��4Sd���pZ��uӚ6��q�R]]��t��y��nN�eBb�"#����+�ψR+7��~��p<U��+]��5�
�ה�2��nh�}���1^C��P)����'��`��5Mڬ{��cכ�20�>-��{��z��������Uk�qSmw*u�lN�,�P�t�.�wM�q�q�4��m���~0�f'#��-�������k�]1�|�ٸ��`Ka��l�>*�FtƼ��C��j%�
�|�VG�2�?�o��1&-�����У����`�I�u�zL�Ia�I9t:Օ)V��d+4�w��Q%fb�ۣ��r�u���HEY�޹�������
�����?۽�_���)A��}:Z�gJs��A��^ڑ�h�vV��D�L?����ƫ���]���t*�����6=.f���@݇j�T.o�%B�Z�V��`�mI�q���nzʃ4�eed���4%=�)�#e�����̘��!@�y���vg�\��a$��CJ��c���\�F�؍�s��O�?Q� �u��)�<��Ck�D0�l����u�D�!��#V��#��t�z^(YX"c�<�*��,�h��x�\]��/׫d%��
(��[�C�(M�e28Z�=�o�5L��&a����n͞�KQ�R��"�����n8�`Y7�58m�nx���D�t_�7���e�dz��w����S�h��fݸ[Qh�,�U�ےNI,���=ö�wPk��8�ѾWjK�O����#�����/+��fܜ�OJ��='���:�u�VY��]��y+c�s��/�ѯO24�|$
l+�^��ydf��X��e�ȅ�s]�U����X��:�iA:���/#���Ȁ��^G�ۡRC��p��^]�J���l���c����E<�gS�!L"�KpĆ�b].�����[n��O�����j@���s�2�^��i�!��ʯw��{&VVT�u�r!�"����ݸ["��`�-��vD���x�}<�JCgDˬ�pY�X�kα�;X��y�Ʌ����|X+F�Vg�����M��!��G������&n/i��A:(O{�,���kͨS�{�G�������OYq�v�#����t��MaZ��dC���3�ad�TO�|OD��xn��r���T�$���O��7���L�{�Ý�"�;.�����w��&��Xl;F;Xd����9�J�B�iRd1ɩ�(��� �ן�ǣ6�<�uI+=��\0�j���Z�|Ih�r̠v/I�fbDoT�Pe��K0O93�7�3��tb���h)�(����� �R
�(�x�:��v��D,�d�y���1s�"��`ǻ���O$4��D�ח3e����!0�SqN�u��w����n=���i��@�J��]�*P\���Gvmη�cN�k�@Ѳ���RVV v��7���M\U8ޡ�Up�������U��W|7�w/���-YՇvoRb�`븇u8�r��g�*��X}}=j�i��j���>F]��V������-��MO�.������"@é�ip�/y��4�[�}/Bc;�=�Iqbw�;��n�R��ٙ�蚍���T�d�ۆU���},���v���ޠ����duJf;R�t0��SH���.��,��s&��M[?��l��$@��MkؗŒb����%�8h����M${�t��۾���4��`@����c�>l���֊���^+�i�J�����$��ٖ�~���!	����%ٮj;�6��B��#R�ic����� ��UX(��g����X��#y�6��f
�d��f�:k�xڟl鮳�]��u����eu�O3<N��������G���/�ۮF�w]0N��t����N�4A���B���Z�5��*g �� �4Î�"/Ӝ��b{�;%w�F\4���0Te��������*�tIS�V*C{h�w����ӅR�(;/DX���+4�F�0�H-"@ ��y0�ol+e��Md�����|g[��J��Q��4������K)aj��7f4�[@X=�iɽJ�1�B����Ə����`�0
s[p�:� =w��4;������M�u��R`�~�
`z�h�/0\��zR�:���-����Eumr�[Pdw��k&���eG6;�����&\;���\>]Ȁ�ڹ�_-,c�9 �:$٠�sR�wW���*���f^n��E���,���h�m<�\�(�)�"���(Ch�8�N��Cw�S��g�q �wP��T-�T���i)nɖ��g��R�8&�ݭص��^�46-��-c^Pt5W*�����~�u��kff�g8�Y^����Wr�ͮ��~ �8�wlÓ��&���n��3	�=��N=�v��\-�"�z[V�x{�ɹ�T'�7e��Z��y�"�Z1w(�Nv��`n(��M��K��}s�g�w'��<[&�E�v�����3��^����gx�������J�����/�*3:� i��c�ۭt.x�in�7q�ظpB�(�K�w��b׎褅n���|Ɣ�Z���]�Ko�}�n��pRoَ��oM��S㔯̦��srP� #H���="b�uЛ�3��6�I�}��yy// >��xv���4��B�+-���2�*��O4�vQ���- �/*��h���S��Qꋥ����B����Iǧ���W;�ǕEܹspummK������;��z�y�6��:�xvϮH���S]/a�$e�Y��NtI�Od�b�=a�`{��O���%����zU}ή����R���h��k��y'mlO��tR�x��N�m}��8�,ȹͽ������CSVQ��xx�3TAR#�'�z�����z��VO�P`����[{z {����
(+EX��Wo�������,E8���S�'/�t��YoSV�;�Uy��F&�V��"��{$�^�c��
�^1��kG�T�L�������2��3�Y�~�qk��c�t�oӰ��j塽;��k{�$w��M�uӺ46��C8zp9��^k�v�sQ�QYF�ӵ��9+ź� Ql]�Kӭ~Q�.�Q�CB�Z*�7a�Sٝ�^��M��4g��ܰ��h���R�������鯥e�4ZL�R�$�;2�N%�rp�@�8�q�������bS�o�����Ґ�Ӣh-3�4��9ˀ��wZ!�u�4.�Vqg�������z��8y����详ES���[��0C�W��!�N��uL�����l7�'E��]�>j��=R]��7�NRӍ(�>��m.c0~ �'}y�ܓ��>=n��w0:�Y��
�R+��YX����k��`�'o���6i�M7hs��we�"���� +��j����ʆ�>wf/�ɼ��i�ISevn[�s"E���o�C��QK2���n�+�� �C���.�c=>�J[kd��O�ݟG���:�&{Lø�N�æ�ɇ��#��M�޶��#R�Ӝ�e2��]25��E��Bk�"������)F���G�J������GC[p�54L��d�\�Y�ȍ�(0��TF���`��bG��bx��z+�v\YMl�S5�C�L������{s�3�����Rs�b��H�l�e3hց����}e�C2�f���Z���ܞ�J�J�2��#K_r"������+2�ϩ�/aQ��wD���g;Y3����g.��NB��J�齴��X/6!;w,�q]�EYv�j�����p
6ic�����mmg.L�J@�˾�ԛƠ�2�Z����u9z�5�t����Ę7�ǁ�Ͳ���t����{YY�vS�{J\������]i�HZ������w!ci�uwX����,r�y���΍g6��bJgPpp�L�l.V&S[`h�t�=�i`j���f��漜����]��R�;X�xT��ox��.��U}��jۛ5�V+8K*0��Z;׹�5<X��2���|��떅*��Yq��wx�+��ZGvI0��(0C�hXQ��W+�)G�7�s&ő�vjOw	�0���ǯ�<YA�swj�mP��\9w��#f�Y��N��L�o�E�\�V���f����(���`�Lu��'=v��hC�ٴ���fh�gMd�[���n'4��jշG6΂]fT�&{�L{[;9]If��v�8�4}�	iY�x���9�4lX����[�
��F^�=�9t/�f��rxA�4�1���(K�R�5�&x�zs�5�5З�ue���E��fT�wIW&pf���Mev��϶m �]����e�S����̕z����"P��y�\�U�2
���-�g�Bt��Ɖl���\Vٱs�͌=4S�:4��ջȪ�_	��k��`����ѧ��)�ք8X�̝9f�/+��z��
��V���jU{[l�_M�>�E�x��c�ѐ�=�.ݬ;�8vs��淫F$��q��d�6�Kҝ�n;FQy��܁�l��������ځ�k:j�w�5�Q֗�)+��_eY�[��i�h3��1�������kt_�+TT8�5�ʻ�ЎT��ڴd{� ��S����wgF`\J�V�۬�Gu��d˹�R�Z����2J�U�nJ2��/����t��Df�ð��_y�׶_X��su��}[��F[˭u}]ޕY�±5��2
:�}�;���+z�ᾡi��)-�;��6K�����mn�v\��q�)Ǖ���oo.���T���<%��*�p3^��q�84W>}�5�ŵ]��xE]޳%�K]m�l$ZXX�;��&<X�ݎ]7nCn�p�X��m>����:��&7L3���{����f�r�^��VVL��O9uo{Ɋ6����Vs+��sC�܇!��,�q)�+H�}pf�7:�[*$�t���n�{�a�@��W
[���I�Ս�Y�{ߜ��˹d+wZ��{�
��1d$	q���!�5�E�j�z����}}q���ׯ_G׎�:l<��8�v�gU���B����)������q�qǎ=z��}v�Ӧ�$� {R�<�N��z{����$��~��~��8�8���z�>�t��g��Q@�Z*���;�������(�d>���ʃ��i}.�}��@ܞRjv$Y $^�*��R/���?��j��u��8�%���_7V�|]���h��wϚ��:��D�:��Ф���[��J�˼��/�ayvgXww��{��w�sn#�����N��du�ypW�Gӫ�Յdu��ۼ����oƫ����L컎�<������<���l��|�駮�ϛu�E�S�'���r��[�)�}�v,;bnu�R�l�M�]�;%	�@�(w��y�����JF⫹��g��� ����gmQ�Z�y�?��vuD���[���شN��B�ZE�;9J��5���Й�q�y�o:�OAns`5gT��/{�p6�.�2� �+�>�O:���{����8��b��knrb���Ψ��*����>�W&�C}rӜ
������df��9�9�DhZ�"/�b�M*��]�y��j�0�dͺ6�l�T�e�� 4PΏp�k�7Ч�O��WCp��"uɼ/�o��k+��-��G�ڊE������m�!>����`�ϸ�A�E�kY�x�̧j>����o�q�W+n�Tөl��OmO���&������7���m�6p�*c��1��˪�n�i��=�9S�����h�Z2oDo_G#~Nn�_T��r]no%���m(��k�E�Ȍr7N�az�z�*����h�=D�S�yqhvY2�gu���9ɺ3{�ء�����2z��7/�0	�������3ls���ζ�L+�2��z�����kA�t��p���*���������<����X�O�e�� Q������B]��4�����W_��M�֭��י�zW�2�4��@�Dt��c{g�aH�PmlN���G1��}�i�pN���ک�g��=]ϳ�ـu��0�#aD?9;��F�\�M��΄aM�����۫^|S{=����M^�q�s�L����Ǣ3��8V�$�>��|������w���{ � ��L�R�����?� ]�D����֨���΢X�Q��P
{_���gf��E����@2`amμ��NR�qv2@��LPOo����Q�L��9���z���-�I�E'o2�~�X�sΞ0�:vA���.ҙ����=ڿE�H��fg���/#JR�uUW�q�nɼ�8iI��3�z�\�ƀ��H4^�������ף��/���o1�+xA;�t��j�4��YK^\�5o>��@j�]��G��$bh���>*6�6S�����7�8-K^����eeM��iא�N�����+�g��4T�� �i��!u�#��'j���F嚺F�U��#������XK=|��L��fm�ʮ�M�Ϊ=]���IԎwf�6�W������Ԍ�٥Rf�����:��	Ά�U���#]Yܧ>ݓe\4fFvf����@Ү��X��}rܽ��ŉ��Ȋ��O^�;��"wl�����5�B��.�t�U��:�[�sO�Ac�[g5����/sN����";��z����*�z����߱�	�'Y��1�d%H�<���8O�7)M�Ym܍k��	uu(6�c5ڼ��=�z*H�b���ٱؾZw��Nߊ�D����ל��9�6I1�����S:�N�֥gn�F8�	b��}�:�·k��Ɍ��z��x���ٽ��œ��C��������'_ޞpK}����#���Y�s=��)��&�a���S#m����t���8����o�ΐ�`V�k���}[j
M��wFk�QӺ�g<J�۪+ʹT卦C�����7c+��mF��_F�;���nH�=&�1ޝ�9Pj��5�Z"v�]��Q��(Z�γ�.�=�ۓgt���g�ޔ4폦��1�Ժ�
pʝWJ8h��9k�v1�6*����Dc�B��6���Q�Z��;w÷�.^�+!\³8T�E���\d�����rW�x��λ��,~���� ��;��j��H�4�`��Ŏrq�*�}�LvWQ��!�7�LM�k]jq�6��� �n�ig����}�v +��a�SB.���h����,���d�H�H+rX���8���,�������[�Jf��ݒFKޣ�.�<���� ��.�:��haaC l�˻uD�h3x�/os�jy���W��"|�_	 �܆/����PS��|�����i��;,�Z
i�u�z�׶�r�2Tv����RL�T}��ʺ�tj�SIqtv���n�b:�W+̷�hNu c3jpԸf;n��n�ꅽ�</���?`t+~��"�,󄑇pë!Y��#���I���ٯw.�IU����~�yC_w]B�����ߑ˚	;�8��a�&�~]��z{������]�H�4vp>��l�Y��	�+�ef���b&:��苶��I����,	�ڥ�0���%��}��ܮ<Nr[��|�P#����C��	xd�0Nh��=5�jl�s�ń#��Š��{q�(1��Y���2�}������x{�y�e��i�.�����}
/���,����#<U��H g&�'��K5Ɲ��1I���Z��GTx�ꊞ Ũ����/w��Bt+�{��%k��2�SR�~�[�k��KTy���d?v��x�8Vz�� y_�yw4v��"��L������r�?���@ސp�PP�����ͫ��W��j��.�iU�h�����to�Ã�x1C��:���C��\B71<D�;�r�e>5��2N׶L%*�-4&q���{���5��T٬�Ld���b��ޭ2�z�'�,��mԍ��wQ�oR�D*�s��t�( S:�9�h��t�/	�)�`Qd0K���5yv#��&:!a��9���2W[��]�x� ��bjM�ݢ�k=�DD���O���F0�u$�7};��8�\;��#=J�>������i�ϯ3���Td��da���i�'b��T�2gfnvk��h�1%6M�)O�ju3Lnp�8�T�Ӌ$Oɗ�e�^;�wh���g�{�
uq����W���a<����K�&ժy��CX��&���U�,��M���{<�7���Sw�aN ��3����ϗ��a�p������Nvl�{b3x浲4��(��25D���g)��s�w5^�u"������6P��W��?W^/��߻�f�E�PFH�m7�e��(����:awq�~*{Ϸr6��i�岑��c�E�V����$����t��{�9 ]q�iRK�h������M]w�˼$���󞌍G�RZ�A�.��\�؟W6k-m�f@�-]�[+U^U,;{A���|�\{�?���6aH��h������Rm*���I�ǻGu���~�)y��=��|֡��y��w[�w�<�C�t��R�t��'Ķ��8�L� �<{�G�p-)u�m5��$�f������pҸ��w%sC����W_����x���By���7���)y�&z|>�E|���&r;%�;*4�bY�j<�Ѯ��r��]�W@�˽�F��:7�W�d���gq2���ܟFjܔӔ)���K�սI�s� �*�����Wx�xI�� Ɏ��������4�ͮ��u�='7����x%,�֝ݪ;�QG�p��Ot'+u^p����?��� Z<��X����w$|��s0�Ĺ&���Wk y��K,`�ֹqWxoa�_�/�M��wm��}0��ח��������o���8��i4�!��;�@��,��m�}���E�5"�V�۳J�j���f�}P���Oc���3�p^�h9]�#}yJ��;����&3u�7�`���wZ�<^E���܆�`�9��\�Z�c�huʹM�E�wN;I�ت�y���sC��9�>|:�^I�;���l��tl�n%��mG��Z�;��O'�Y��Y�:�xt�BH�hG2E�:��������_o)ow��4C�؅��θ�dN�e*��=�3F�n�����<^�W:��T���[8����G(�� Rod�GZ����%*��X�LS��l����;����y���S��|�G���Щ�=C�R��!߯�Yܛ�x���`1"�{Ͳ�<Q��1������0F���1�*��X.���⤵���b��7'iY�<*�G,��no�Ǩ���:�n�Sz��r���ci�O.u�
4���bKJ�Z�_d���w�2m����
��y�����s�WFK]�=;Y�mn���!}��%w9�C~�||||G��w2��+O��N7�����e>�5��\k���_6η6i��芝y��ư��-H^��;}� ���M��qt��e������Eb��7��[Ę)gCP���2#�dli�{=>���n(*I>��]�0�N>����w�=�Ӌ5�Fy��,�z�v ��>���_Fƭ{
ݔ+]��f7f�쓯L���W���(�`�ȿ3���1�@���=�ݭבX�Y�wFE-�D��qB}����+vJ��^�r�+�89R��	 �SX:V� VWk���}�M������=��*q�<P>`�P���s���%^hX(��v�P�f�E��13�
�$�3O������b�'*U�'�p� a�U�b����ɢ���͛lĥbe7���W�E���!_�&�����D˧�Z��w��vО�&��qm�ʆS��}u����Q�����_��@b�.��F����Q���ٝK�'[�	��)K`�ѣ�X��2q�����L'�(�E�Q��q㳓�I��:ZE�!� ]M�Qk���7�T)�E��f��e]ng9]10ƍf_FV�љ�� F�G(ݱ�f�X)��� ||����M��}>�]����3�ꉸ��nu6%KǠ���>�q�A��G2�y�E����I� �pm�E��n�KĶ��`������!`gƦ�{�]у۞{%���������{#rߤȑn;���y�q&m"�z���k�I���m��v�ܖ׽�z�R�嗕��u݃�]���k)ˀ�:\�"���'���_o��_�}M�^u�����i9���X
�[��.dG�;|��#J�����+T�*�� T�&mģs��Yl����q����#�g�]�<zM�L�1��ymv{t��sy^�k��6K0�,��ޛٞ�T&'-���7Y�Z��xwye����&{�x-�2w٠���g�u��=
XV
45�y�s�}>!mJ���P�0t���|=���#�j��#��.����coU���X�ҭ|��TȖ�T
J���EKC�j�8`�qa�p{I+�a�-t���j�}�,�XF���M�>�>
5uѩ��Ȯ���,�7r5�TU>�^7KH{��I_�`F	[��'y�׶������;�|Օ��`�$ϒppIN�^�/��DEh�������X̼.0��EZT0c����F><� ��֣i��O�g��Í*4�X
�^1Ndo7�e�Z�=�H����>���O�p���9l�c���'v�Y�n��>1O����ϯ��@5�K������	9aj���n�v��V�#m>��⡓n��?�S�)���P��"���+�{��n���G{��7��O.�W���j��歟}5�(���y3C�����:U��#-�a������K*�8q�A#�B9uW�n�i��'�5�2�t���Ӯ�:�Od�����uOg�=��=�c�w$�ǘX����j��p�G�s��$+�>�vЄ;��Z7d�r�\^�m㫙�)��Z�R�n�Ბ�>nm>��|Ge��7���p!�|��Wm��Ǚ�q@�ƺ�sfg.��s����y�S/{��yd�@�e��pP��ވi�6�]�n��d��њ'���kn���2S�Fe¸](.ԫ�b��ݴ-�'��[��̺��ߴ�����-]5'I�8�t��zv���2�(�ѭr�(#�=��6�v�C���55e��.;���q�7Ň��e�\J��̼���ƴ쳪em��1n���)\2Ĺ��5#5I[��n੺$��&�J��	K�O1V�]�Jij�c��B��ri�$8T��q�����=�p(�츉ޝ{Y�=ϺGb�<0Y����n6�������+;�<�7Ǯ�˞�t1�3�R�tV��Q����X��������ZU��U�{�=�r�F��;yg�4����Z�
����OR�!�3�<;s�nv����gbnی��OoI�74�[d�(�;�%pgWqy
�mǹtw����S6��,��n�P���Bh�c�ݫ5.چZ��^�+=Y���w/**���Θ1��v�kL�¬U:�/*5���oF6�]:��-˅����"���Y�о�k��%���"�V'u[<�ӗ�(_>�<�c���r�̱�kr�ܔ{�V�Qɯ�T�P�KK)9��E�P�a�sN3X*�C����fɯ��saVo:8$��A�k���h���/1����8��{t9"W�"���*��Wb��'6���n�G2C�R��|4�fx����֔�G�_'}':���c��Z�0�.A�'#%$6tj�I7^����_`�WK�ȬIF,)�I�)�{�H�H��[T�ѩ2���3w{�2��~M��X	o���s*a�%�t7�����|�vy;ݔ�#��fǥl�����L�2:ϕ��4~Z*Ǆ?d3��98��Z�,��n��_b�M���t�yΕطϮ�<���ä�Zh�X�ɶf��^t��%��}�E����D���y�s�qa��B�m��j�N�iY4	lRkr�&��T6�^�͹͓�Wf,Ŏl�:�P=+;1;�SNI`��:5���퀮�L+*m��p\.��&S� k�1\�-1tac�MfN-�;�ו�`)̩X:��۱f��##z���%Z�}�M�zT#�|I�fU�j!�N���z�c�͓�R�u��pgc|�:7X�a4�wUUΣTۅe��)3:s�6�h���s��a$�Jp.�t�$9z𞉨��3E�:Μ/Z���ӧH��D���i!\���o���<���AmᶋΝ1\�Z�dGM�wv�S�H&0d\�̏L"�����EŎ�R�,���g+K�d�Qj�����K_<Ujj�stأS�H�]I�Sp�._Wp9y���2�A7�p7Ȥ�WU�@�1N
�e��df��jӓ�i����Ż�v�`�֤�z���]�fp���9���Z�����܄}�@.;�<�$��#Q	�*\RU2Dy�S~T�
����^<�z��8�ǯ^�a�ۧN��)4�9,��?=n���w��n�.H��tY��λ�|��w��x����8�<q�ׯ��v�Ӧ��}n�W��vecoׯn����#�[�J�D�R�N�>�v;x�8�z�����t��J�<����]��G}+��΍#����lw[�t���e�n�m�k;��c���6�X�l��w�֬��������_N��+/�j>�vg�[8��;�Yw����;�ε-3���ok�..��m�fgi���^<n��m�fwG�`����I=�M�jˣ�������-8�������g��K:����t�ӳ�,��ζՐqǾ�~h���zvc��{Aq�W��Z�Y�����e��m'�v}{]�};���Y��v�:(�*ҭj�[Zʷ��.;�E#��>�@Ā�Ap B'���Q0�I�!�@��Q� ��X���1�08����b�GB�ڈ�xKl�U԰��O�7�.�\����)��)�Q3��[��q�ym��Ul����W��xF�\n�*�,�1H�)E>��Ri6�1��ɐ0�!��[2�,�$
�>!��D�[�����!� �P5QD�,��
�)	�|�)�@��5�F�p�Đ������y^T-�]�J�K�_X�1��l1g3�&t���u�]�Ҝ�7U������2I�+6P!���qb�f���&'�W��"Փ�9S��:Ku�c��뼄�:����uNi��k^5-n�x���r�ڞQݕ|d*g�g�0�I�%�&F��}Dq#mLR��JǍ�vPL��������ބ*�F���Hę����\'V5 A��\�.�J�������*wQY=�ݺ%�N���S�4���@����c?���R G\�Mq��K���6=u�������6���s����/`�gBj���W�"Ÿۢ��*�U�lBӘxj�_�டm�wg���Q�x��]1]�5���"��!��VANL�{J�'�KVJ׋pq|~����G��::&L�������<3D_�W�}�<%8��F���v�}�;�4��\���;�v,c8��ͧ�nْKGG��<ِ���q��{�G5В5ڎc)�9��sߪv-ΰ��fj���wg"7Ҍ�m�}�w]�ZkVұ�dWu7vK�kfe2s
�$�/��䫵)c9}*G�u�S�V�Z��3v���ܻ���D%�-�j���4�MKA��|�6�J}c7��8Wu�Ͳ.���`F!��ӻ�����Uo�O�>V�*ܘ����x�i�8��RW��;��O���1��a�����3@�g��׋(V0쎠/����T_�]��>F�n��j�F�U� �Uۼ���ѫtI-4�4�1u*<��͟K]?H���~��߈��ozۄ7SC���9�_BE��>L(l#�����l�n�ƓQ��w�F���[�J��_wM��[vǻ����,E�;�Er���n�#��Fs��p����G���^?s��#�	ڹ�}���[S���<ռ�$�"Ni���G:(xC�w;��Pu�`Ot��uEyWW�+L���L_<�
���Y�у�΁�L��6���j�w�giɠ]�TC��ft�֭�ǀ2�,��{'�7l�x����/ou���I�Ү35�-ՂQ6_i6)��43��H�D��!�8<�^��Ƿ�.H�y�U\��a��[ �YLI;��
:Z�Í��mX�yY}�9�:�*�(�fR˖�|!�~q2����	w��g4�Ԝ�fA+oj`��Hv��V*�LYTA�=],���7�Q�dl3���Gz|�7��x

�J�}`��xh.]w{Tv��G�sX$����:'�;U"�����L�Dƿ�&����uϺ���u�{��U(�R�$t&�֍�v�<+Zp���{�N�35�]�e�������"ñ��,8��[F*ur����-`Ϩ.��Rj-�{��S�����e�\�c�2�L��x��U^����V7Y����8&a��r��,�KznsNX��z���d�(G���%z�=Ô�s��6F73P���fg(W������x��̊��ӹo�,���{|��&�fp7͛Q�сEb=E����wpc=��_r�d�
gF��2QΎ� %^���p6	&��lE�Q���� ~��	˃��g��6�H�M+�3�������9��[���מ�	?)��=���u�]�y��xRj<˃r��/:���!���B���j��YUUt������HFY�C������nNL����=g8!i>�|ܹ�z������(Ǖ/��m�]��s�7[˒�U�ݍ�R���:Fn�G���̛�9��J����1	�沯=<�n�o��N�O�3�6@m�yd���B!t�	�oUs�S����[;�+�f�(�xun��@gl�fǘk�
}Ƥ�]�ϽS�����n��|m�(���mMu�[Zf�[}��=9���k�4�nA��Ċ���5]�7;�y����.IӉv�u��!��~�'�[Z(�tM��os¼�b�>W%CL�H+��1��.�7$�K7��T3�� �6:���ܴ`�̟S�Q;��b��iyS7qӎ�{�׳iD�y�����-E�����> �	<�)�>����w���*̶3�Nܫí9�a�3w�omI�}v�N;�=ܪ�2�C�\���b��^"oԽ��M�3S�V�4�yjni��`ަ�@��W�j.�MT>�m*[��T���G�����4#��[wQ.��?g�-�+st���{DlN�*P�S{�4mܯ�pm.2��N���-V�;�+�Nq��;p�PN��tn�>�� ��b�@������0]����<���j�99���˻����z��ݔ�j�g&�ސ)���4vFm/~�||||G������c��~wW��/A%ͩ:w�c�05l�=��,�jg��NE��h\W�q��i�~���f�@��d����P�]�;���N��z5t����ż ��:���c��ߴ����c�an-�y��Ky�[P�vI��Z����_m��dhWǨ�n��kl�'���&�f���{٤�tύ��_+[��1�q�8!���0��h^�}�3Y�<:�ؔ�+Y��0��PT���䧊s>�1e���j�aL7l��|EZ��귲F�ZӪ��m<��v�{0.�z�O���쒥��giGs�kȽ�j�rL��Vo�� ��$�ow%S�b+Wlm��
�S�Gb�5g��O�%������}٠��H��rn�Z$�VdY�ċZ#�ϰ�]d�hx<�b�mX����/��.f|�l$*�O�㵮��m4�k�x��g����<���ɏ��.��ةSQI�i����n>��)2��Ē#����_ۗ`,����Z)���V��:���a�o(��uMyYs�v�8�=���"H�̨Ĉ���Obc]oc��.�}ؒ*Z�a�;rE�	{�;B�̝�j�W:1��w;��������r|c1��.�,l�Xa?Ų�(�ؕ>ꍯd1��L�Թ��hg�1uQ4��/{ŅT����
�'Q` VR��s��X.��]4X����|��J�'��Q�jk�ǀ���O���j�}�������om�%E	�o�vY{GT@{����j��C����]	#\��T����EO&ۛ�i�\�^AU�����t{�����i�2�I��n����+'!�-��XBٟ-���o�(g���S��*���8�F=��n�)��gw�s� �J�r��������~�r:#����x��}+w��{��|=��]��6$x�k[1�m�u�pWr�7�y�r]l�Dj��>�P$�e��2Qǐn��/��-8	b���-n�^`\۶N���0w�7�^A��eBI�M���F�w������jH�xr����7��\Y����}��iub��E^|�r�f[��1i��ϣTur(}�l+B�^��.�p����(�l��ytr�6�NٖC�t��O��,s
�aо;j�e�l3����h����� �A��K~,�b�DH�����@G`0%��.w��S��g<Ouz�v�j�Kܥe;D�ve\�3�<����'˲�r)OH1���PXJg�n��%��3�OU)Փ��c|��qc��d�uֿD?]�V�/n4�g� �"��_e�N�:>�>2��2��=c*"��#��vf�f����u�K�y$+����:5�Y�5��5������I#�j�����sHUo���/w��*�r���;x�y�:"�G%G!ʠ�E�|ޖ���q3�����;��
�<���/�g�2v���:�j9�檃qh�Ӎ�v�V���<�m�&v[A�-�S1R�s���ȸ�SĴ@��w=\��f��MT�`���l�}+c������'T�Jv�#�遻Þ�����(�B��ݱm�n�����~��[�5����c�ӝ+�T�]K�7jhH�1tw.	u~'X��K��2u²*�[�5z8�G�=��:��I䡝����1~��e-JT/����x������Y�����9�/�����1�`������}�L��K�-"y<r���誠�>�ا�9��T^(����J���S:=Z����6�|���l�rO����]=�$�^^6�����9g��A��g'飻ry�oq7x^H�A�(t��ct�������uǸ��㔠��:q�;
a�VM��U����ݼ�9�-/�:��`���coi���=+����U��{�gn�9V^�f%�P���a����� ������}�8�r�ε�j���.�TT��x���ޣ6_�X���]}F�����[��W#�t��q8�e��7�TO@6��������s��q%!�ޭ����|<�9TMC�84cX��㯯��!7��}�F��H*J�.g���I��̈�&���t��,-3�v�u~�!%�2sum�샶��v��L�g�Ɔ�����-�����uN�r��&�wk����'#l��V�EY0f0o�G>�k2���ܶW1s*U��ob ���PC������(���:WΖ�.K���Z�0<2`\tpTŭ����e�u |�Ɓ-dB�wgj�+�;���y�o7��ԍ\j�̼�̬gSV딷���.Y/KP7%̺�W��V7�a�"H���{[/J�����DU�\���]���{b��B�O���Gy�i�ѭ@�C��T�;�K�%3D��㏇�HNqu��+R���/-H��R�8ី���ZY�������8��n���:���B�*�#s�۹4�㨐z���H�D]٢_5ݚ���<�T�v�P8Ö��X_�J=�˥�7rX6p��n��/]\��QS-��޷�qܲDs��H��zx��U���a���FfɊ};��ŋOS�R���f�HY��`���U�,**�m=f]G^�#�ۣݦ�u��=]C��A6W��D1���n�v>��Ç.�{Fo^0����܃���*�4��	JN��Q�KJ���1��b���~Q��g�)�<^�s�[���T�0�-���-�;�4�o��}��$]\�+_J<�<�\�&�1��F
�X�ڽ݃���4pG+O��>�_x?���f�807�1��Dr�͌��[Y�>쏥5���{%������Y�������yE��2j�y�����ȝ�J��a�w�.�dD(��h��)�ԽUX��.�s�f�d��.�`�!��Gt8�.2�
2��1�;(iS���u6�34P��	xo0^|������<�aϣ�ܟb�H��|��ZݱV��X�L[M�ӭ��t�r[��;�A�v`�������9���Yf�wI�fԧm��Q6�e�bT��}��~�Q�w�Y�-ͧ���H
=�j�助��w���#QlX�F�9�`��2��H��n(2ҳ5?���Z��*�wm!ī�ܱ�ٳ�鱭8�"�Y�a9�(�,Ԇ�?�u�;Z�}4G)��o!��G!\���6��`xcx3֫��h��������9�C���+(D����]5����;[������������P�emU�zߦ��qΪDr���guP>�:��y޸,�c�W8xL�̢h���/u�wu�TZ��z�T�/1�3C�@z�������b�ǫE�׼W[�{$K	Onc���G>f�`]�W����a�paY�\���ZTHCSu�M�9ʫ���y���n�tخ|�k�}�L��K��.fή�a�}��%1ʗnEW�WQ˻�����R�6��e�8;�礪�nU�u0�R�"����{;�����V�D�զ���]������^���%�Էp����o���Wv�ga�&��WY��=c�	��tT����I�����y���}3*���|}J�b'�렝�n6:>��
[}�����t6�)�@��e���9�*�2ѷ�X]]owc��PX���^�5� 
_��\1S��F�	�&J�}�;yv���m�1�%`��r7���ˍo����rm���r����>�k=�_c����;5�v�`��6��In���d�o���rZ���N�Y]�������45��8+�8G��q���0��E�ݾ���5�5V��'���A���^�oiWI��.�%�l��n�.3r�`�w�[sz��&.aݗ��{q��Q˺�	��� �:�{�2�`�.�XΒ)sx�:*�Wkf�
H�fm4vN3̃,٫�;J/����ɪ���T�ȋ�)�x\I@���/�m�VH�Ǧ���ۺ&|˗��%g&���m���uֻ�cM��n���p:��TӼ���j��5�F�\.e�ԹǺ���ZL)���c��mX�擎�Q����ľ�YZ>7��%{4��!e֘�d�{�11ѡ��'ZDe[*�hɷ��$��]Cr<�N�Z}�&߮+�<�g9%��.�;;�z�Do�olӍֺUȆ�VN��/l�ջ�I�\�y��x�[�tW��+j<u���x��6��XWy���.�Jk�`>]� ���:���l{�t,#s7dT�k���2�^@bw)x�����x�/����էG�I�-��C�W4�ں�p�����'֮�:�n�Ы��WTRCWʝ������LP�C�!���p��(h���nvr=t����v͡��<�l�v�֥�V�n�[�o��]�)>ãD�-f܄�̮'���c�)Wt�VW�t]�,Ԙ���|�
沋�i��%,�S��5�!�ye&��"����:�N���K��̧{��vfY��d�j|4gm�ܡ[��X������j�K�$+��L��;���3���i���3��(E������u��3}����M���b�B�|y�d��5�]�it�z���23VQ��`��<��!��z��]myݳ|]�7dXQ�yhK�U!(�����;x�v��q�z�����:t�MB����.ADM�.�F����sZ苙��~m��߽�߽�����8�8��ׯ���t���r���[��w���+f�����������k_l�������T|}x������8�8��ׯ���t����	U!L^"B��I;�gE�kk�I���׽���ݗY�r\T\u���s�9OD��9,����?]X�̜E};{Y�յ���~��8��6�r��e}U4�,��ם}l����P��V��׉\tW��p�gm��R~��I�RU����AD�{q��99~l��u��n���R�=�INW������u�ˢ���͵���������-#� �D2����ժ]��ꛟ��p��0���]dHY�.�/�Ź�C�]��\�EwH�C��S��d�ZsW�rLc�g�����^�]�UQUCŋ���}?���_r�����N���]ϳ��뎱��Q�`꯶=6�t{l<U2�j^\��z[1��t���]�^ع��w�-�"'�Bxtu�1�OM%\z۶;�vz��6��"���al��b�S���&��z7�����mwMwe��q�fR,ȥ(�x���y�l��R"3�B����V�.�i��Ⱦ�IڷsU�ު��#]
�$m3��p�CM���>�o\R>��u7���>�׋{����/�ͽ�Aq5^S���v�n�~a@o���r�y��nÅ��ïϡ�^l�������H�j2X�,C��̴��Kncqj`�͹���~�'�7`�����(�Z�*�
;LX0�����T�1�3 �!�|�IP�1���$���FwM=l��xa�/3��j7hcIu��8z��a�.�]��mu���2�܎��P=���Ә.fC��|�#�M�on�*��Ùg�)ؘ��u-}������G ����t(BU�]�񩷨� '������o��W_��*����̭��i�J����o�#j���)@{�U�s5N+���+P̄�zo�jo�ЛKv��8o�L��ܿ��0�z��&����E���p���R^��,����qd���zR[m��</Cbl����S�r�u6u��f`F���U�=�������;܍���<M_� ��ޕ�Rq�Q1�i>�[4��5���ܹ�S�ϗӴ��t0������Y������sq���C���8(�?v�Ի�v�$�,��K�*4�̔s��L�t�8���z����<~�V�c�;���h�y�1v+%���F���1�����8����aO��2��H���x<u���پ�F�u�
/�(� �xE�����7!�]�nd���T�~'[ʳTI!����o<���^��n[!��~`[��]��(�a��,� �o%��5����p걳��]�H<���jׇ0.{�!J압lf^������G�ʈ1 (�;�e�����6��Y�����K[]��ݔM��1ј�R��֫���K��Bum�Y�r�NK��T� ����=�uw������;ͭӵ8M�J����qr+��c�rF�Ġ3ƾ��=n�li�]�D�X�,���Y�b�IHV+Kݸ��������ͽ!ϛ�j�N�l����$���]��,��M�9��x���ĸb�6m�(��T\��M��^}�4^�ȱ��eu�]�\oY�2���0^��x�:�gTo�|�ی".��SQ��SWM+;��[*���"Nmo�s:X�
�����/?wLMI7���u6��n��VAO#N��DO��H�o\�?�ƽ�6��wvk)z�`sU�D�U��&=0��=ެ�+�{���M��V[(-�j�j�9�bhN-:)�T?I��U���uw_o��ǻ�x�ʹ�e���w�X�v���jx�O���@+�������8c���r��GLl�A���R���uHe2����^�Y1�h��N��䙷�uU�J�DW�6$^Wws�U7B��Bj�h�8��a�V�G���2n�*6ɗ�[K&�Х��p����jÙ�zĽ�L�qs���9�7+�?�}��"��Bag:楲�?(�"��u�����]���];���wU>�8��c7���w{�4�oڤ�)%�Ye>N��0�.:Z=�_�o9x����m淓Q��Km�����`̸Dvw�l�dϵå�컮Oo���h�J;c5���8{\�+�F��q���=yL��l�ɸ��=.*�vF�P�O#!�)�ol�s�t�y������K\u�i{eԭ�#��!��/.g��N�Cc4�=ҹ�O/PEF꧚Mmw�)�����f�w��ƿ�i���ˁG>��G�s;S�^I�
��І�=��_>Tl��֭��98�V��c�u�w͚D��cjۡ���S's۴d�g�;O�p&GPg�5��CSɋj��3	�ͯ�-k��1���?) �P�sbT�3��p �%����an^��ڬ������-C���Z1��|/t�>�!�δ��pSJ�X�r�p�m_c��đ�'2c�~ٽj�3^��Jv��y�@b�����_�<���5151��{�W��u��v�>��I �#�]o�����}J{�!x��1��VKk�G����:[�7E�՜#ʃ��x���c+��vk��!ڦJ�p��`h&��j�#��@���9 +�{��X�]��\De^޽��pf5�Y�C�.��S#�)�q��t���;��mT.��2j����9\����{k��:��[C���K�R�y7���!q<G �\dw*�&V���@��xK�s���#�;���~nq�Ni]�;6=L5�x]��#�uS��:�ߌH��Wwz�P�m=�uG&�Zb��
�Si�c����G�#d]����!�G9VV�Ѽ�ܬG�
�B�\�0�]\��T��_�O��L����[��	iT��:K��c��_pF�(���eokɰp��K⹧�p�V�2�����'�)�� �_�7cδϢ9�8@�BL,d��{W���;��;)R�H��2��0q�3�<#܋�{c�;5�e�w�ҐV��*��}����Hi�Z�֬چ�Fw5wW*��^���E6�o���F2���u�B%��8n���R� }K}o]tgl�3�-�ُ���2ND��3(�b��KvU)�X�>�y��o�x{�]�\�Է_~d�RմQ5Jo�+onX�o���qQ�|����@˳\�@=Yl,��H������Rď{�=�Pn�6Q�+��Z*�r�S�^�D��b�jg5���2,^�+�
A �I�	8��׮�	婳d�n�pa�Pσ�e��ʄMr�]z=�p���d�ä�f��7Ui)ӛI��gm�ק�e�: p���O�jdTz���6�kR{�Tŝ�t�(j��7�$\R�o[Ƕ���z�5ü�7����lH��JV4����l]�6B�R�!#m+nD�yP��9مϨv9��,C�J~���s�<U�=�way���gR�]�������{�q U�j쇶�U�V��+����@������CLwP�\�<Uk�vW$��q�K=�<�"�Q�%����D~qK�j�������xo4^��B>�.^�=ӵ�TP"Af��;�Ɯ��T���U������E���l�%5EK	��Ut��2�ʺ�o3��ͮYY(1\������+Yg3*�+��Ȼ�i�����5Vi��5�42��L�����B�j6W]ύ�ߓ�j��>4�1� 8l�&l�{&��c�1��D�Y;�{&o����S����HJ�[�$��ն�����f���� ��Z��F0�f��[���*�0L����5�f�`��$�ν�9������[!#�#�ο���]Ut4�GPhܱ��a5������}ܱ!�_dt3�q�_�;{SU����H����n��w����Q��y۪�=Zm�n��ē���Es����k�R���H�b��/}*L	ff,uviD�_TzP;U���m�y��[s�;���;�¨i`w���e �{(j��t��A.!�Ode���M��c���4�fD�B}Q�D�;�)J���5W�{t���C{� .�ݾ3H@�93�+/���g
�u�,������xaq�VnA<�G.����^�z~�d<E��t�S
�#��ΣZ[%�d�������#�'��c�-E���g�o������ͮͺ��h��U['E6��v�؆m^���2�<�p�4MY��(Ku�s�]��N8t����wx�fB����[M-2�ݢ��q�ٺ���h+T���m�R��S,�]�ʫJfu~�� ����5U=N-��y�p�A�U?�.�C�jR6ה����;-�Pe����`��Ly�:���l��g[˻��Oq����x�1<�D��_�k��&m�h0Cj8�
�~P;2vCd�CwLLDb�s{��ko2
6t�CRY���#�]��e4� ��+^�9��ݤ����GK���{9�C�0�IJ���>6s=q��o8U~�}}�Q��냉p�D�ջ�z���X�u3��vA6d2m�����f�X㙭�MG)B�D�3��:�m�'��x����=ƽ>� <�3 n����+a�S�;q�4��+�<GHw�0���ުry؞AY�iW�D3W8��c=\�X��k��j���t�2"3���F@��\OA֊���'F���^���.}]9��#���q���M>�쌹m�� �W��YYyY5K���mdE(]	�h����������rt�Ca�ei˸������:�vq��q �O�������AD[@�pR��u5Hn|������澁���l0V�PP�Q��0����n�|������7������&�s3x���n�_����΂H�����ßh����|���`M]�:ƽ�R_g���V\����N��2z�ƻ?���N�#-�0���q��3]�1s�GP��3����>\�A�lJ�q�}����*��M���X�F�a�ܹ��[UI{�kǈEY;���\�l�h��7df���@��;;k�p�t��T���#*�9l�����hܧ�-P�S�_OJ��7����Y,oe�t�J�L��"�{��(KS���q�mF��\�(j7��r��uX�B)O�����昽��sr1C�>��8Au���z��d���y\MS�pN9�+�4�U>^4Nna9.|���٣���k���z[�.��]TF܍�~��+���T!7|݇�J��AP��>_w}=�m�.��c=#���z9�`Լ��&���f��X�t2�u/H�yB���~�j����V.�%�Ǫ���T-�77��e�����w�����٘"�b��6պ�e���"�d�\i�'�:>=�t^�H-R�[lЗ�)W87P�<Jޕ�V��������o7��(⓫c����v��,?q�!��V��'���Swi{蚼ݦ!98�p��ǔ�z}�]��[�f��s���T�'��l���R^��mh��8��K�l���k����bO�o�\ �CY��D�/T�%KoڥWw���� �y��`��������+LVϞ�#��O�AF���5d���� l���C���^ʬOBCЙ�
�Q5���7d�����vU��3,�%Q�a!Q�fh�E����:Yx��q��)�g4hB]b��\�Q��=��&�[����x�$�|�M26Z�v4𹢻�d��\�n��e��mI�ܭ�t��6�{oZ_�`��8R��R"}�k���e������c2�3lB;{��l�>�(->h��'-�����+Z�G�����z_��G� @k�@�����J"�����W�� �j:7^#C1�(�V2�A###cX�D"  �0A���E# � ��R!X�E"�D2 ��R�T"�DB(�B!���B!�0@�EB!�"P�A"H1@�5M�D ���B D !�BF�D ���B���B D !`��B�D"���B �D ��Q��B �D 	�B
(D"!��B
F(�D"!�B"�D ��$B(�E"D ��B �(D ���B(�D !b!�$BD 	��B*D"!�����5H
D ��$B" D"!�B�(E�F
AR(%E H!@�RP(B �A� ��B* U""��B �A�"�� B �A��b݂* 6� �� ���B �A* � B �]"�"�� B
 A���"��B�@d v+dA�@d A
A�"A�D ��$B ��U(S �*D"�F �`��d�FA��B��d`F7v�b*FFF 1
D � �����B �d`��P�D"�(����,d ��1��F
��T���S��wN.UW�&���5�n}�ޠ � �$b
��bgB���|����??7�����k����?`���?�4t����J��������~�PW�?x~����x��"��T@��G����,������'�����X� ����=�a?�촋_�֜���?�N�~���>�D����Ta B"@��"!�����"
XA���$H @"���"�QwR�uN�uJWT�w\�����H"�� ��B"�'�H(�QT@d �Q�S���몒��N���		�		�B0P�D"�BD P��"�@""�A" ����B	�"@��P�� @DBDB @"ABD �Q ,D"�A �",Q �T5g�J������?� P�QQ$�R@@I�O�}����??�	����p����@h?m���y�����/�V���?���G��*�
��֟��<���A U�* *��?�;���"����@p?�%�x�����}i<>�D�q���x�Ҩ �>�����C��}��������������?g�~!�z�>�� ��84 �*��!����
�`<�x~;CA"~��������h?Y�<΁�w���J���rH����% ~����,?ۋ��>��ZDE�A��f�D[���9����HR�?�b��L���0	��� � ���fO� ąw�|�T@(��
�R	
���UU*EU
�EUQHPH��*J %*�*���)D�BIT�I%"� (�"�)B*P*R�$�!
���*EB�R*TEQD�	 �%T��B�P%*%@����J��Q*%*@�U**J�QP�%��(�(��*()%R(���Q*��T%!R@� �
ERUF`�)J*�8  �յ�SDe`}9P���&����9ۑ �ՅjU[c&S@��i�kl�(´���3I ��g]٠��U$IU*
�RZ�   Y�Hz�$V�E�@�y�΀���T)�/z+�()"!@tL�E�!�J�i������cFJ��WTa��'Z��5cmAF�&���4����@�"�U�%$��  v�	[SL�̪Z�
��6�m+i��Z��$Ŕ��̡����L+h�Ц�Z��j������J��ťh�(�
UHT�UT*E7  ��HCj�Sj�+M5j����u�T�c�r6��Z���h�+"���[t��Q\�H�\�R*IH) ����   3� f�h��Ҷ�TT�K��P��֬��̌�Z�Z,��ZʘZwAv�Km��(�$RIR@"T�I�  g56�*�����Nr�� ��j*Q�m�m��dij�֍�m;`h��ʆ�Ί�֎�aZ� ����$P�����   ���l�u� 8r�* �n � 9�c�  A�P )��ҝhwc����]֮ h�1Ѻ���$�@����  M�( W:�� 3�g@ pa�@�� S�,�A�Fp� �jܮ���C:VN�9\ 4�vt����	H��  l�@P[����.���A�p�ʔ�SZ��t, ���((�Q��)J�P�+�;f�Z㦚� 9��$)J$)
!DT/   Xⵦ��Ұ�N���A]N��t(�s�  ]���:N�5�@7!�� `�t  uo "��DƪU#@24Ѧ�S�0��� �a *x&H@ �JR�  ��T�MF�F@��)5T� �3Rz#d@��	Z)�����r��!�� B��ؤod��8�1��"��{Ժ��j�ֶ�{Z�����[Z���������j�ֶ�mUV�������u�^�)���[Q��Id	.�ݩ[kL(6](���fi��"�U���^�܁(�.�^@�%r�d��6�y���K�SF]�B�F�iHf��V1�sv�ю�(I�ԬW{e+	�­�t͔o,��1&�l������3wi�ɩMxKŦXbdܧ�U�/%�"P�v���{m�����[��2XMՙ�e+nl��!�pSզ��U賛	kkvl
"{Y4��]�s�P1��C�:��j�TR�O�6�4b�a��.��Ҝ���U�E�n%��A���/1l��K0�y8�b�%Ǹ�!���vE*�a�GU����m܆�r�J�w������!HՒ���Cʽ����Kv`sAS+"�JhlA�6VN!�S0�K�f��v*&�M�Iݬlnm�ЕXY�2@���f��'6^V�i����ܕu���M�q"]&����ɪ�TkhT
�	�v�0�m��b������u1ѐh��.t�bk���L�b�֎����2�V�I`v��i�Ԫz�f���J�r�7qn�uk4\�Ӆ���]'�B�ܣm��b��%���
�*3��H������c�!�k-�[�ެ�!�LD��\��j��k�IJ ����鼅:af���^��i�C]��Lڴ� n�̉���3n��xK,c`9Aᒎ���@��WH�Ի:�T���׌�(�f6�-��9pP ���c�iZ4�s[V�v�;��Z��\8���n�f*1�R�D��5�13Y�jI�5e@LW��w�VOׇrӂ�B�ۓ+6�"�&P��f�q����D�V2��H�"ѡ� l�K��6��,�-󩔑�D�	�=��"X�J6�v
4�r��
�
��q �W�iބ��(ջ��B�]%�؎�p ۢ�k%{��
]��7X���L��5�ƪ
oD��y��4��f�i&Շ5)W���9u����t��.m�څl�k-�X4�T�k�iܱsD��2a��ۢ(O��-��4(V+�շ�}�K��F�(�e�AK�Co�%�!@*T�����Yyd�-��Y��%>�a�4fƦ�Y0�T�r��m�U�����[�.��Bk�8㌼v���l�h���Ϝ�˻`����%�u���W��ZZ��.&��B��m�n�q�@,���))<�0�iZ�õ�+cP2�,�mLq�d�f�V4�ɛ6Q�]%��4%�������M��e�@����u�; F�0I6�&�z��fJe-���Ā�B�������l�P�δ����j���Y�	ledц'��ɬ�0#	^��l��R���Л`7XcŔ+Yx��C5���G-KU1:�+��u8����"6�½��n�*0�KԬ���X��yn��`�����fV",cq l�"�Q#h��Lf����-A �U ��4��3e�" �����r��*.�9��U�v�B.��4&�fif�E#y&�1K�ց��
,\�)�ol���+W)̫Y��{5�	5��ۭO6��˭o[�Ö~"1=���Ւ�-�),(�����V2��������L�y�f�!ۓ�h����X�+��e��x�F�f�V�Xwz�$;�p�#C5�����(���[��ӭ���Y�UJL��R▄��vUeɗ):���77fe@V6��ef�6ٛ�Z
MQSUYz)���r��T��- �:��bX"#j�b�x�Zb�Tk5���M�Gt=��x�vvA��;L'�B�5iGZ�ix%��ZN�X�bLn�G ́��4�
��0�f�Yj�v�D�Ce�7@�f�EM��U�� ��H�U�R=ʄ�z�<���{<�S��i� S���T�h]퇙x�.V�逎�Q��B�		*l�5]�m��WF�n"�ւ�
��)b�z���hG[ZT��d�X�Մ�B��ɶ+���i�;ŷp�jL���pٶ�Cs�	{�n��k���ɔ0��0!g��$�K^��5��h@o��OOɰ�1[r
 -�)���
�qm��F�Ts1V�j*	�� �MXgY-+�J�T%�U��]v���TE�bj�ȍ�.Ɣ�b�l�H�J�b�����)£j��j;��u)�QP����Pj-�R�����w�����%��L��ɯU{�0�Z���hndʸ�@��r��i�wgJ�p��i�hV��"�1"l�m��)�-�S���p���ҳi.hf�8��F��Z�i���#,-ҁ�qb�Ru+a���b�n�bhn�ʻ�{2�aeB����" �Cb��e�+]�SF�y5)2]��M�x� �*'#ƌ�z�հ)Mw�rQS^Jlf�ҥ�i+�֭�Z����U����a�v4m����>N�>�陰5L��X�����waw+ci���Z����B�,��o��v�7�
][�ݝ'h����Ux�=
�S):ǡr��!�X��&���x2SL�܉cJ�7���ʗ��S�4õ��W����"l	���ۍ����n�e��e`2��$�! ���nkC����;���)m�4D��)h��� ��Cy41dGI�����Sp�g���S��{�6S��++rܼ� j��tȰ-�{[`ܤ���n��Z֥3l��1bn��:�Z��cR���cwV�1�j���:Y��6Q��j��N�n��?Q.�O@;4Y�C�.�$&����^��X�][�J�D��= ɗ�{��Ⱥ	Ćn��!���e�Y�Em9Vщ|����e�TC <2i���m`R���˗Z��4$j�E�Tꞛ[�v8�T.���X Uq4E��Ȍ;C����}���Z
kQ ��/�ջu1��ei:�!�s(�d�n0��F��k�X�-�)W�6�h�-@��²��@�pm\�i�k,Z�q��$�����w20�sCǲ�yf���U�.�e'�&ҷE^�Yd�MMn����o�,�6@/R�m�BշR�	�;�#8��[��e3wz�qjj�������T��[]φ�1Y�	w&�G0JL���V�?<�	I�D�*�F��w7b��c2Z�1U���S{6��V��i;�q��3'�ݟfa֯m��zYUd���fm�]欬N]=�q�˹[ ����R�������@T���R�m7��CI62��0�]6*�6��#p�Zw
)���
�Z�YV�c���z�!�-IB�u0b����t�v���z*�F��F�B֥�/�R�.�W�1fB���Hhk]�]k�V6�SJ�
����%���wa;������G����K@��v]��.靬WqY�n�0F�Bi�fQ9W�x���7�KU��#��xq=�p�JĆB�K�̒��i�-��\J�[����d�Q6�+YQ�*Jn�!�>x�� ���KA�v�iHҼ�Q�v��ĴS��U��f��n��XA�osnh0�2��42��J��ͻ�7u�d�i��ye,
�]".���kk���42evAe�5Xiҗ,�`	V�ᮊ���ݩV�8��a���jCyQĔ#�{&
n`k��5mT���uoe0r��u,VVYn�t��U�Fe�J�L�U�bڃAJWu++u�ԮP� hy*�L���,�zn��e����Fe�E�ܺa�W�v���i#xV"��T��Z�ܐkԡ��hr�7X�f �v~�Y��Hd�w��n�r�
����;wэ���D?JN����ŋ3*�Q�]���e�BѢ�e���3$���V�]l�.E�]�ɍ�y�����R�$���i��J�DB��� �t\��+���F��qhZp'@�%���51in�j�XE�q�Y�0��CkH�(Ѻ*ĳ�m�+^沑/ehe��kS�Ы�e\Ȧ�rRu!�ӕf��
6p����ҫ��B�y�n����S��n^�h FE^f�K4^��i��b
D��I�ܽ����R�-��΢�E��I��zɮK�Y�23o]_�m��M˷�ڧV��E�o�S�xO��a
���+zq�NY�$#.bNMB)I�������ޕF��&��0�����;bwo4�-��)O�USշ�^M��E�!X!,��XUM�]`9��L7v�@V�l.kP�Or�2���7P縉r��J�֐Y�vP	<��1��<�l��@�lM�X�lecs[�"��az���'U��7�-8,
�uz��ӳ�#��Z�u�Q��MUU��y��.������d��M�h�cl��<�p���h�ct5����]C��.��)SQ��7�ɂ��"ĺS�.ц�S�WPՈ�q��2�4����=9X��t��o�7��D�B��tUKK�ͦ�'uny���cn3%cT���~� �4"&����UcM��/HٻZ�_l��W�pǴ%��+*Z�;�N��#T˔��Z��t�2�6l����׵n��J�JS9���XGj��0�0b��	3W0U�(�U�Q;����:��X��Y���'{Sr1%
<�WWh��=@�˨̙�X)c3�[U�KTE�%�-�kpm�yor�x�XM���R`U5P2Y��S���q�:[�pC*P*���3<��*�X6	n!���]ۀ�#4�H�M4��b���.�!� E�LT2Q�Pљ�^`�*B,�cn�I`�6�џ`�t��+E+u(��]�f�j�`h)�c.�D#��6,m4j-��x��JQ;����Fč������gU[�C��ۇ��#�4�*rk�eɷ���Á��+�|�ѻV9L�s"ik7�J8]��]��aR�u��e��V-�ɶ����	-�[����Rc�i���F��
�Q�:EDB݉
n�L(�r�c#�u�$9FU��hZ����DԎ"N��4^�n�J���;u{Kz�N��D�xǕ�X�r�����O��[*:��eeB��Ԯ�k`�ѽ��#',�e�xUm�w*T��x~?;;tѓ"�d��Y���g&ڦҳ��)��D^�5f����ĥ���V8���<�ouXf�᭸�-��Q��mA��TV�Y�X��nQagJ���/^A�7�n�I��"b�A�Y˗.�5�`nH�k#�%G.�����W�N�i5�T;&dwZl�Z�Ť�q�ӂ�T��ױ`ɬ�Z�k�"���^
��m��.:�[y�.���r��S�m٨%lx�+n�NlT͹�)�Zlҽ�Ûv��vU���v6fFMaN�4��Uy�4թ�����kA�M���UkJ���Zm��7`���u����A75���jMغ����%��V�9�ʭ�Q�v�U�+"3r�M����j��8ޭ�(VkL��	Q���[(}�@j�e
M[ٻR��Yg��1��3v�jIسz�AQ��Wt���5*H��W�ek8otl�ڲ�R�æ��[7)�`������9��Cut�Eac�[B�@�v�����ʔ�����gN�bP����t(���nO������
PdodUzE�%@�v֤�|n�a�V�FR-b�DY)U�dg�24�*��S)�z-�#b�1)E���7���%��!�&)`�����rK�v8���F2�0���L�MĔ��XN���l̳$d*�	c�JU��v�Ђ�9	6�K��k$�ۼ��*����gpEfe�C����3hQZ��/�65=��Ҫ�7�c"��b�m[qУ���0���E�@���w�V�Ww�6(Т�u���	�n�N�<՘�ۼ��r���*�;��Kkq�r�M-#5n�b��bk���I���X&i�PD����50:�dԲ�,�QۘI&��2Y�)�{h�ki�j��
[�"%)@�+ZG���֨Ez7�Y�w칐3�m;�umT`��F�:��gF� ;W���4�ب�3�I�j�*�g84T�I�bv�#�2���¦�[�Zf��+�o�o4GGK��j`�Ma�m�]Ġ7oj�'J�,TU	/a��+�hlV��+&ԏ.���4�I\B��\ĕ%f�+W4�\"���\��緍@�d��aŀf*�jV�f�)��MJã1-�95,R���K�Rk��P�Î�B6�����8aÏ����q�y�`��	7��I�u�� p�Q��,[ĩ �yn�4�I��<.\��6�0 ܚӍ���Mң�%Ӓ��5xӶ��a��1�\�`�	ճo\J4c�iҵe��'^ivޤ2�&\����p݇\��Q�u`����K�]L	b���E]�X�k���M �lG�}(��sr�h����:�wR���ո��ڵhh����t��6�j��M4aP%jA�#�n�`\��Up}�G$�[�1�0e�^��[R�����[FP�ܓ,mhW�֫M�'Ṍc�	��Zx��	*Y٥Q8��8-XܖCN�]Ԑ�ւY�=��6�G��`�2+4�{g~��^ّ�.M��j1���̐�4���Ϙ���/@��S��w��_-r��	[CY���|) �[*G�B)�Y�  ڔ"4m��Lb�˷Dv��[���c3i��&=U î�q��]����K�q��	�ˡ�$i�SZ��<���KQ�BfV�b�Ri�,]�z�uu+P%�	xԸB�6����3s���`-�[H�ϛaFE���{nioBԦ�&��w�]�PU�e�*�I)To)j��'Z��#&�jz%�X[{{��/�GQZ钳m�No��N�,%B�k�-[�ob���U��.��4Ӕ�Ë]�G��3{�G\��:�I������-reݮ���X@wM�޻�O91�[�g�v5ҷ�+������n�3��u�����Or����z|��p\�]s{A�]4�^��󓺻y(��`�Yӻ�\)┭��Q���G�������c�d��kg�7C}�{ׅ��� 93oc�&)=����iV�����E�q��W���ч8��b�����)�|G�r�cY��Yكs�)@�W1�4�b��;�B캳�o)6���Z.�E���pB��,BwM��GW)B�X%�RN�u$н�M䓨�n��W>���&��e���C�=o`�]9�r�4�L�6/gcFx/"���,��&�~�h�6�{9�)�wWI��y��.4Q	���MlwG8�y����E-�M?oHc�s�6We'RB�5`tǌ���s�>W��l�(0.v���h��!�$nL7���<�������e�ـ.�'�o��)�	����(+����7/��X�0^�om�@p�64���|�k��j.4n�Z<[]���`<U+E,�f��u�g��N*� v���ۀu�6rZ����E����!�p��p���A�T��߻
J�mB�AH��7z�a���`Ҹ_]l�������;L�}�U��b�^ܑ�g����9�"	����QKi�H
�}݆������7�%*�]eG(NY'������\3�l����B�������;x��YL�����:�ם95,����Yؓ�wz�V�Lp�q�,n����;a�^�M�LM��}���i4�Ʈ��9�Ʉ`M����e��ګr�Vx�|�nJ��U�O:w<H�V��;�R=��n���N;6n-��\ڧ\�����r��}��Ȏ�F�XR�j0/g���n,�좖ֈfG���e�u2�鹔������m%�8e�c� �k ��֛;y6�ӂ����_I'|�d[�|3K��pZh�����h��IǗs���:��>�ګm2�\��u�;ka��~�=�e_@~�T{���H���1�=tUk<���[ǲ)�X�
Z	���c�zlK�a�� �����M��dh�֛�W\�o�L�}��SW����6h��G))��7:]Щ�N8nX:E��uIs^�>���)h]M��c��v�}{���]_	L�ԩ]��i�U�;����x���r����޴Зuv�C�7y��k ��1�`����%��Ƈ^n.5�U�h37��T$砉�л�&�(����v��e@sV6ӣ'�6�n�g��}}��Z�o�5�]a>��=���B��h ��+s�]�Y�Ub[}���*l%\�=բ�p�c����x��
��3��X�|�����>[�eD�b�0�Foc|7�%m�J�ooOA�CDвt�h��y�We����ERoc\޺�����Y�ʓ/�A��Y��wW6��{m����j�s�Y���"��x�U,N��T,����k;k�q����p�����I�J	���*�Y��P�`�2�Ix5p��^rv����r����̥��?5Fq9ҕ�����U�5%u<���KT4��H]��Q�r�g����c�5^]m�o�<�m��K�dN�F�Qwa��.�N+���{�d�;�歰��#ؠ�RS�5z� �g3�N�]�;��[��\��im,�F�c/D�*.N�OU�d���uud�HNԚ��G>)�X���H�������M�j%]\�7��
��Qffh�Ԩb���I.����.�N�/�)�a}�*��E��5��\Tx��*�3��hS)l\�d;��u��S��"R�Y��k��MtXk"4r��>l� ��#%��!J�;�J=n��n�^bb�%	���N����N���]h�T�1]=�%1Z�r�@�u��n���0�<廤�8�x#e��2��__'S��2�\��r�F�P.�<nM���	����%�S��~��������!���鲬px`�*r�F��*ɏKc�5�U�L��XV����e�(wf��,�]ns42�QG��;�&s8�8�<�@��YZ��6]D����	]�ڃ�fek_^㝀�P��i��t���-r��yܶa՘:�r����p"^�%��Uς�F�V�v�O�����PgA��I���΋x���Q簐k�5�:�A�0-;z�zda#Q�}n;r�{�{�w�}��ܳy���rv
:��f�Yق���:)Җd���B��]$܀�(�#!���[w�wʠ���e�c��ɮ���]��;��k 4GqΒg����,ϖ�%+U4
{�D�ӂշ�G7�G����e��9gZ�7R�N�_�*�Ұ�(ଆΌ���<�Y�=:v��g-�K5H�S��҇wΐ�>��2�J�2'p��p�Y�Xv�t���x��A������Ă&��{ô�ĂP魋"�.� d�*�gIڪ�ܡT�FM�_mf�X��Ww��v�h��)�%vqf�i�sQJ������sH6�oP�@�˘v��y`������n�!��8L�*��83�J47��u��h��x���WJ��ؐ[���Lu4�S(��N-q�fެ����u�g���"�s(��:繍ù�ù[�,Zఒ��X]�	����],	AR^i<��̓,o,��`��r��t���x�F�x�K"�����#ay�8s�n����}aMZk��j<���)RV���)�%׫>ŝ/tǧ����v�1��}}�;,*��O���s7�+A�pwS�G
.�鷚6��bn��M�h���w��䭦m��O!�BoڍY�\�CM�.��b����k1��UH{��hĒ���W�^��z�t������u��7�}���[�t�L��(��G�s��ZTu���_ҷ:��v��OyL������*Z̵��="����w���{�MQ��X�l̒����.��B��Ι#�r�%� �1E�%��Ł��.�
��vQnvS�ہev�l,�`�樼@�*H�X5��U���$�BMv���%T�̘@s���.PD�ĞL�&*�w,�t��W��G�%���v@�b�oCx+Z�.�{�!�wYۆ 0T�@�Jos����r]j������4��ۦ���Zr�r������Z9�(���g!&A���Mq��&��܄�P�a�:�w9�Tu9���8��}xoS���4�F$�l�f�Sy[t�I�;�K�d��vu!#�5��TW%�f���r���F�wGi�Nc�9��I.�r�X�t��OGDڋtRP��KR�/kI��w�=�zPϚHÏ�Y1dU�f�N�/��3n��{��Ϣ���Rxr�+�n��os\���Z!b�9��`�oMC^(2����V2,��Uc���B��l��ȟ�;�I��W)`�:�ߺd>�F�v��X�1�s3-	ԛ��pǷ�S졦v��f�r.b����㩣:��Է�#�8�^��.��
�[��
Q4 �Z:m[t�3G�Dґ���0ї�3��j[]%�.��S��ۿ�����zDS�o�[P'���;�q��˹y9t�]#��EzE���u+%՝�h�7���9�`Dh��.�G���oWܫ+�;B�b	.���J��v>��c�Y�Y�vd�y�"Z}�e-���W��9��7��_�D�q���F�2b+-�;.��K��ފ�R�R��b�Wns��e6��w����L44%}u,��׬�֫hɓ��jĺ\���]�4�6�]�6��������|�Q�뙯Qa���5֙ֆ��ë.�"�g��˖�1�g�9ZR�ݼ�`]WgY�,c��-[��,�b��]ʼ��{6�:<����hG�K���4��	z����,՝d�]��RT���Bu�C�ӧ��t�M&ˬs�j���h9�	*�fRCPN�rUX�ɭ��8�9HGJm���7�fk��scX�v�T��.��V��-�#)k��r�P�kj�Ґ�o�����#<6��/&�/\;�O��뫟s�ʈH�p�[l�;�채�&k'U��;(�Yƶ��Q����\ż�p�+��[=�P̭�sPww&�^��ZRU�A6���V�pY4׺p�xu��Ջ��;��jr؍�]�׎ϫ�@�U���Ǐ�!�J��t��KwNw}}���)Lx�NLS�uڈ4��G^M��&#eF�ؾy˅������x�V�Z4��(e�OZy�l;��,k�]�'<�R�&�SR�����'v&��|�M�f��Z�݁�RS���^c�/�_L�,R��8u_k՛O�&#���g^�X��r겸�ŗ����Y�lT�u�q�sT@m+����S(�i�ݳ����������m���K�U
=g��iLm?�Z#}5y[�ף*�-����1u��-��y��ky�JS�	��[���\Z�T�S�x)�M&|0h��}!c����S�o��8�1Z��)ս㜑��=ܛ��1N������a�o�t¸u���h@�ss�ޫ?t{W��l���QޚkX�G�<cUe(�:�n��f��|{u�ՠ��SwL�QL�����c�&%2�'H�<KiJ������Dg�[�CY0Wf�y�o;�t����ӫ�Xd�sp�֒MsQ�9��;N�uڷ�jh���\�)S(֌��isWs���;YbN�͢⫗LW#���{m�S{H��\8��8z�J�ڡ���[�2���T'��T�Pvp�CCt��̼gq�X����E�z�L������q���ea��j
����8z�h�����-�,=Wj�޹��T��wSn�n
ş%��
��V
N��_.R4ζ����r'k�h ���л���[n�ʝ���V�=\�S-�.��`�K��ġ�m��~��;rhG�}��/��� �P[(�5|=k9�`���Tx^��M��%=�E�q�N��W�f�I����U���9וg��z�*A�<�w�-�̭|�A�*Ub�AS��nQspeiu,�/������qQN�Ԯ8�:������57V�Y��ւy�[{՛�U�� �WO��U��.ԣȠ�OY��亿��n��}q^�<Ep۹(�n���*px�!�Mk9�[*�ZŽ��Z�n-�Ժ��	鋞0��bߣ�,��ռktQ7V�����9A�io���M��J}��f���<AO-���������].�	���4ƫ��j`�lkVg.�SfW�`A�e�Mͨ�j�ҡ��s:�b�Ђ�[7 ����f��M^��([f�y#k9VVJȫa�:�p:�z��U����dޣ��0�E�I��'S�w�gP��=�C���`ǫ+��T���#�li#U�V�8����M��3�	1JX_��G�X��nCNAV �w����;�9q:��
�OjQ!���-����]����A��
a�%'�PRm-װu���_�lO��=o �4��E�&��T÷�Zr�>�&�<�r\�%J5XE�4�u�9|��ϒ��R���*X�)y�v�\����g ���:���sa�}ԩG�A�"��.KW:�-�d�h&�_t��������kT�yKuH��Ub�ݏ�S�9�Оj��[��n)��*��]�c���?vu[y���jK'��*��I�>��4$�	�t�9r6�ݜ�}���2e[G�P�M��si�S��w��J8MU54`���v���8�-�3��.
Z.VV��a\Pu��*�mw<�-��>����ǂ�!
\"�^�õ�2�����,K��!�/-�K�b�$9a���| �RW�t�/�`��Q]!�O���s��bJ�[ Drˁ�ŕ���Q��Y];q��ubȧ�ab�&��ĥ�К��I�d>/$��w	e���sF�|w�7��G�U�xij[�b2آgy��4�"�i9�0��X�t�ꗣ���t��G�ېu���ת�՗�҃��щ>+���y ��0�]XFu��HШ4����r|��-���ܨ�+�Q�4�6� ����%[�OX}x ���V�p#�KN�\^`t[y��uqMgu:�y�S���wS\�u����d�	�-�������CF�C��Uӭ2<ʊ�AM?�t}גƈ��b�ӕ�b�ԔF��z�/��G,������*��.]&~l]���ʗZQ�}V�J��$P���ڲ1VO!�J�\�/`/��w͍��Yn��]cb�FU=�WR9��	.��n�m4�	��3J�F 5ۅ蠭�|Dͷ`���O�/~;W++�'��ݣIFަv��t�=��t����]�v}+s^w:�����@tb�Ԯ�Ϻ�ъ���L�}�U�^�e����io�ѳ��c;W&����h�5:��~K����;w#D��Q�@+:�gf��^6���f-���3�-Û9��nZ��Z\]��� .³�%�h>�e�|b��Z���W9���q��a�s)v��-�g{�����q��c�SM̗X�>��ˉ�(��[���u\��q|OƎa�[�v ����.#E���v#ͫ+Wu�t�Ll	[��v��h=�e7Cn�n���o��>��y�t��;��e��[a`K�����R��q�*xZ�-�7����m�]P� S�U�:F6��e����3�Ȭk9	4[5}�@$�Z9�˲5]�=z�}9S�b�IɎՎ��+ݭa�˱of��8��<��SgsY��)�v��_`���=��b���=]4��׬��{3�12�\������|X�]
f�##��}Y�9��}��RR<m��gRg������H���d�L�m��׎�������Oj���'9��hum��§f����@�a�v�u>��e�����@��U6﻾n�,�ͭ����gs��{�w�~���� ��?���{���>���K͞��p��wy��u�^������3]����;hX��XT�b�x_aS�8���X^��޽� �፱9���6U
��&�n�٬�U�$��1���)���L#n̜{;f�S-��kS��!ڏ{7z����M�ݻz��:ɩ�7��{Y6��S"!m���m�m�ur��ڥ�
�� ��x��ݺ�h=����Ios����i����%��%>Z�<�rA�"�c��4{)��%C���%|���Ⱦ�1Ո�^�!�W����Y�U��8��;�Q$�����Z�6׻"V����[�a%�:�]�l!�M�춫�j�1�u�����eA�S`�]���L�;�!]��鉦�-~���_oU��S�vSc�v��wb�&���Ѧ�mѥ��[��	u���J�,&�R��i�s���:`�t�p�ʺ���[���nA1��(��,��c�.�=kB�[ nm�+�ukKB��f�x7Unk�I���f�#l=Z�(��7n�E�;��a�G^+&;�n�v+<�U�+XZ4;%R��Y���h��W!Y�L��5R�����Oq��g"}������SK��2��f�;��.]��r�-�u]b���ŕ�,B��
�|3'*Q�o��^�i��n� ȧ����Is�ڂȍz�{ue����F8-ߎ�Z�++^c� �\m��x�.
�+�����V���;�o�Nuk�xE1��M�[yp�-��Bw�h'!a3���Yz�ie<7MV�I��Ⱥy�!�`iw�ZJ�r�uǉ�e��Y6��[�P�.�FE3(R4�}Y(K�׮�J�H���Gk{7	eS������v�{z�˚h���:/�����M=�F`�Ov�'���3-=����[
�lX�B� �����n�}�YQ����C�RSd��"f�X-�d�
�P�Gz(���Â¤Mm1�'mJõ>E_ ����jY���Č�.�q$���Jz]c���<Scsw7N�F�ڼ2I��۬lsR��(���b�5؆�}0Nhӷy�2�c2�(;�I��p}��>����V@�B��8b��[��`b�Lg��}� T!MDwX�:S�S+SR��Ƌjģ��^V�BVW|��١��h�ܵ�QBjbA�;.ܦ�����e�7�h�鈲����u{v�,���(�ɚ�m���Q���#	q�t��7�.��#7ݬʵ|�nn�i��+l�+��]�'U<�n��.	\+2:h�h�����ӬPǓ����[I�A�99���������o�hۣ�]�-KNEʾtҔ��!�k�%�p�nq�c[w���']mGj9��v�w)�6���m�`��WT�ݝ�v-�k��0���Cܚ[8�5��إ`yWy�r�veep�:<��×D+�(��-p��C��^��Z=)TF�{(q�o����F�^�]B�T��弦"h�w5��J��#a�<�i��/j4q��+Sf�],�+��ki}�]�m9%�����+�Yso�
���ٌY���N���_bh���	��ȭ| �3�oT�[��g�i@�����RP��a�����KD���=גkX>om��`�����n�����}�u1�k�70ú�hh�ʹ
Ra����vu����z�(�v=<9�ջ�o^�u\�oAޘ�K%���x[z(�S����$q�
��i�)�]��޴��Q��M�WN���9��8�
C���]�����Ѯ�	��*���$*-os��qm��l�4�p�d�쭾G�W��^����^�l	�J��V6�3�.m
p�+�Vձ2��ŠE�䦪�cB'��3t��y�(m:[��v�a�Y�]g ���w�E�5X�yqvQ�얲�v7Z�'S��(%�yX���v�o1v'ř�6�y���.�PH�5>�t�l�U3Wg 5�,���FV�Y죮�ݖ��wHXʊ�`T��&Ҝ��L�J�-�93�Y�L�.su�˼�=��}�o�'Z��dVr��pȯ�ˮ�m�f.(^m��[ (��e���뛶���[ݰ��5�a�t������\��ⷶ�Y�AoLem�8�y�^�)�֞3�q�`k�Kr�\�,�P�ֹْ�[]܊ߥ�y4p�ǂ�$�K���jIR�!�[�}c^1��m��jڴn+�W3�*�=Lep��ꈏ�m��i�
3�Wm|�q�ɕvS��M�?���X�0(��F�������Lk�z��T���sG�b��!��Y}���Р�Ჲ-9�K�Z6��q͠�u";���������E���}9��$�̊�-�憎�Q�
h&@8US,�������9���*�E�q�+w�cp=P4��S(� EUǗY˱?�mwuܡ�/7u1:���@Э�ۓ*��1Q}Fw4I���W!��a^��>3��N�)j���Pø��\3Q�ð
�ھ�ȾS�=m9F�^��<(�X�R뮝�3L��ͥ����w"���_,�rd爵�+8+���[񭇋�=��,"&��ι]ۿe���iwR4'Moܭ�8�<tP
��땐�.��1n: iZ^q�٢g���E��j#R�k���G3[B�gDwp}��+�j/hu���]�)v�bOrN�1�����$(�/��#u��I��D��v�>B��0wv���nd�
w�mG]36�]ÇQ��xg5�1M;�A���4�e-A�"��N�aϨ87`+�AqF�j��vWv���>�Mo�q%��gd+i�g<��h�Gp�&Qs�ѣ\�4flK�S6�@!-�Ŷ� K&�C�H�.Z-c�dxUY�kc���������.�C"$�q"J��І�kz�����T�b�-8�y�X/��9酎�pY��INr�����L�S�Le��j��MTIJ4��8&�p=KoHUsvbsK\Swn�̀��H�[����1��A��ňC�r���ư���+)WVT����TR���E$���͔���L��Y�-�\��l���*%c�w��\��eL�T�+���&ݕj�ݹrIY*i���AOm�oSE�S��`���W�ij�HSh�:� u|{A눥��Y�����"><��Q˾��ǧr�ڛ�y�2�֕�`Tn�mN�rEc�JIt�罹�6�ow�w��Ь�H:��X��n.译�qӔڛ1��.�m�x�������۽�];�9{�_a��9�hr���]7�>�tJ8$�v�q��6q��	��	�����.����sC����
f�2�<�˭���yx7 �r6�7Ք�_Z��r�r���G)�
ghx��.ЭlS�{�=/��0�A�2���GM隕j-a��a��5�us���c���/^\Q�3��.�N9y�:��c���*�������Q���9i�X^��IVVӻÀ$�٭��o���m�Ʌ����g�di^qa�?s�����o�}Ę���������{�0��%�k 3l�A�1ti�����[l1vuv:�v�봩�ˮ�TX�6�(�ή
��mѝ��'��ʂ�5nT�fӼ�fcB�+@,vbn�}�����b:Z�*���Õt��k�l'es�Mr��\���	�B�W�b��f�ņ��`�H���v<p��@����⮨�U�3!Agoj#�����0v̘.���\�Npf��oJuoU���
�Օlh��Ż�n��v>��BU.��!̴��k��]Pu�ݮ��D���c���3>���;�ͅUR`�|�鉱E&���V2���n�L�K�V]z�tn��c�.ᶇn�ǖ������Ы�)T�η�Yz�$�p{�nZ��M�X���MF�t~��e���Ȥp���uގ��t�\�N�3�DS�c2������{S�n�n6�Ѫ>U��ӳ�p�+#W͛�!ز�Ɯ��C��\����l`}"F���]�Ԋ�Skr.�2n>�46�m!]�j�s�-	d �è	�"���yK> �l��o3Ҹ�J�9�V�ji(٠u
���F3E!��U>딫RR��3��4�QX(n�лt��,7���������	�Fs^*z�a�}9�㈥��z���� t8��@��|���s�"�Lo��17"{WV��Jۮ2��֐�G�;-�����]�YD[�h�Ύ��z�ԭ�x]ȫl�����U15�HnӼ�h��㎮���JG�[����H���.���>���iMˍ�u��;_2���\�u�M�뮣J�֨�ΟlKhn��<ކx�Q��Vsg��[�5�!]���ܛ;�9�zA���82������$�.��
���L���-4���0�Br�9
���Z�B+�k\qZ�ܧ�w����*,siST��-B��:1�yQVM�	ќ�RܬQ:��!�y��Q�����{��*1=��m�S-ޅ7R�m����P���X�'���U�T���9���P�[�j�7qu��T�m�B^&+�aV��s���69u4�8+.�pY������\*N-n�aK6;v���Yڏ j.��]ћ���MS������@�ޚ/9�X�#�Y�`W(�ۙ�'��<F�^�I��*De��J�Y��6 �P3[V�Q�t����������f�6��1X2VWK��Y�.��ro.|��yyA�X`�T��WP��ח�(�Ҽ"�@6"��������',����j˘G.���R�7QU��:B�V^�k����ฎ�����@I��7.�+�1�
��M��]f��dm���m����E�v���n�j��N&�EGUmY7}8嬇��Z�B4�4��[�M�|q�6�t�#>F�;�22�}��U��s����1ޗ(p�xБ_:�h�[�_d��1ul��)���ᅎ�๦X���z�Σ��p=��'2�|%<�.qv,QxWi��+o���d7�ɮ��:�*+�f=��5�J����;&`�����*�6�G�J$�hK9l��H��z�E�X�k��;q47����c�kg=�ZD7��$ܗ��fAFr��t�es�|�����ea2L�@�s��7�j�f��˥z6cg�đ�����{���}���Be�]/~�.\k+:�^(�4����S��@�v��\g!L��IQ���=#������T�:�zaDqXq��P��(\�w����BOMI����N���^����Ug�Yg
*m������n�h���ln�bt�ؽ��	�#-D�GHkf���n�6-�L}����A[d=��[��Ҩŀ��5��Z��Z\��
MMY�&��8h`ö�޻nJ���m��md�oජ��7�%躒�-=X�fq��`�+�m%��� ��}q��F�!-����<���{�J���)�U�i`�=�Pi.����쥼�\�5�V�noُ*�)�EN�bI��ϵ�n=�ae�rށ;%��G.ŝcn��kr���g�6�mA�lX�f�!��˔-N��rʾ����5��yK���X��|-�WemA�I�#�������{/#�@'gȠ�v� ��6:����l�ǯ���B�IwhCp]��+��n>����Z�`0:��݉3@ �|hJ��f�F�'y-�TCqS<A͓vb����j{���:5��B`ʄ5���mge9Q�Z�?-j����A�ܮ]]d�dogc�[Ғy������S�ԞN=v�u|�M;�E�j�q�B�5E�R�h0fMr�Vu(xt��o�((t��V��w�0���{��2�F'i�ط���.��ض��')�iF�J�w��*�mk�.�Rx��=��/6�6�M��r-�AWiR�u��B閍�'���QSf�\�È5WWb*���Yݻaq���+��%s�Kj��5+G�V���`w^��2�@�=�`��|#��H�����8q����	�T�yw�쁩�Mt�Mug`�d�9/�]o�'p��J����P�U�:�|���[�A=�6�RX���ȉӧ�b�ٽ���+Y|��-F^�ۖl��(q�(�<p
�J�'��ݵ	��yZ#\��Aوڎ�V�p���r�tAN4�t>��j�����͘���Ի���B��7,f^QN����6r5�%Z�lA9�F1�}`����j���x]���kT�SP͹�����̢��ŴjT
X��FJ��*
��U�*אF�[���ooGX��w}� [C�۠ά��BH�;���6���i�3�\�d`U�����6J�6kV��*&����.W��u��k"ݿ���֠��;xE'O()���wJ�����P�%ԕ�-VP��Mm�_Y�FSy��xs������Jo[�6�fvÝa��Z�P��kf��ݑ��ՏqU�54��PY���f���d)v/Hs��
�^�h�׌+�:U�r.�H9z�&țye^�S9	�VuN���FDF�\˖���/ZA�Ú�Q�HpL�W[G��-�\o"vȓF���1�,=�+���$������M�Z֍9�P�͞AX�>���M���5��h��Æ\�$UlW9NV�o�E��ۡ�E����A�&e	[�e�Z�Fsjۈ�{h���(���8m��u�y�) �JK;9���a޻W{Ӓ]}�,#Ů馥䒶���%�K�)�,��loKo*̖7��;-S���ty`�b���t�%f�2��<8�9Ʋ�0�9{4� ]sƉ;�9T%�Ƹ�+H�\��(�U�"*����fޚ�ْ�v��3���Q ����霑s�3�}Ѯ��^e֊��/�$]e�$������&j<�u��ݻ�	��[4��u�P�4w��E����F�U�Y�9bc�S��s��VL�3�z
Z�W�XyF�Lq쎁]��I΍=y�j��O���������k�l1��}=�/pI9�u �oj�Y�F �sR+M�ݪ��R}Z2ҕi��z@|�c�їk\�B��kJ�|��s�os(��4�����z��OE��&X�G�]Z-ή�o�k+�:v,�+i4��y׆�-v�~ӱj�|��ol� �[���I��(�P�b�Q]�ۢ"�VD*��Z�fe�QA3u0ʻ�,�#�|����[Ni3��VX��mh�:m8�V^uk���Wʆ�)����&_�)�e_	�dY|�J99ܻ@����\��!q�{zc���I���[5�=�31�WRՖ�d1�A��FvI�h<�AXç!G).�јܧ���7:ܻ��Ū�D�3;�^�C-��3)�7��zV�%�a���Q\��kN�LV%�A��4�V�QG[��wٷ�,+&���Э�˃vC�,��9W;n�s6�`��JBN��l�K,���C5:�{�͵�p�XȺ����������̧
fPy}$��:��]{�hTF`O���8㕮����+�S�+���ڸ]���u�t�8� b���Kb��r��b�P���v�}(��,/��ch9]ʺ(�).�ԕ�4��إppu^�5���� [ͨ����AS��Z�a��m*ʋs��3��賁�v.	/To9o@�)�X�o{�_8NMy�&p�H<U)� �ht���S+k�YǇO׳����wwt��� �]Av�w.7 ��Γv��)wX.ݎ���75�w9�M�Wt�ۚ+����t�s[�˹�������v����v��wf.�wD�l	��s��1�]��wgv����tێ��� ���&HA˃���k�n�λ�5��I��wv�ȹ�\���7+��IQ��sn�W9�;��X�;��;�DfQ�;��p����ݤ��s��]N�GwQ�p�L�:k��G+���.�����D�F���W8k�����ҹ&awuˑ���$̹����A9]Gv�u��Z$�f
Q�b�jN����E$���9ۦ�1&M�Df���2H\���q�>7ޜ����VP�H�W+�C��������4N��n��r{�x�Ps]եntv��$I��ٳx'[���⃱�_}yy�6o�}r��5V.1��`�A�ֳVԺ��5$hT������<������ ��\'��X�.�T³}b��WV��G1���x����8d�K���I�sqW;���\Ń�	A:��5д��^��l���\k��&��ggk��$.�c"��9UכR��11\l-t�,BL��Y��"�zN+�l5U���7!���突wg�Rձy,����UX}a'\�=�i�-�l���NE�"��E�6n�m�P�������#\q�����F�2g��������]Q��{z/���NI1�V���C&ٌwK,�c��l���ۺ���W�I/�m2H��I������>�|��I����P0@�!�ڬm�/�y��nOTtDtt�Q^���L�@����l*$,�H�ۥ�vf��w�Õ�>���]һ�E�~}�C���Ԧx�GW�Γ ����2x�,�4b�Q=�J�p��4r�s��C��{HG8&�3bۇ�;:eBQ��&A����č���V'�[BL����� %�^
�u�ö�:�!X�q���p�Dm-�Ԏi��fˏ�g�k�����ܷ�(�/��Z�7�L8f]`y؎I�w���B��of���nX�ܷ���6�����(�s���YW;��+d�{�M�49Y3�w���	C8Z�K�s���8��:�`�T�@���G��UC��M�-���%��2"�4
#E�2nR�������"�7b:,�>4���v4�ȑ�y�19#a��m'L�TMz ah@[�� �C�V�w<�2,�A�+��W�SKa��� :1V�*�ȓǈ'��Aؑ	�TX�]�<���b��T���%n�׭X���e��0�u�A�� ��x�ߚ������|{�G�m��=��SВ�j�ݙ�������j��jS��m�:�u�ׇO���8<�Y�%�l�䯆�5-��w3Ϭ�X���L+b��冓��c�(�nX1�����G �<A= 䅹
twPQe�웬bc�qP� vF��G���eE�loS�5:&��u��'��#ne��e��}���7�g:"1���Á���(p�d�΍ˠ�Q���X�4DtN���L�&nvƷ�c��{U]Q����D��wg�1U����5��o�xrJ� �0�弎bs�pЪ+�Q�&�mm��r���A��:c6�4E2���z�ڲ��ݴ�6����j�u�,��-hc��fD@�tX�͕̅��Q���;D�lmHm�*�3x���bڲ��%��W�E��W�Qy7Aux�m9�oK����9\�4��q����f��}�yg�z��eў{,�����+O1!�1�C��u���@�급P�jH^��������P�dw��t�����^J��pu~��p�5�O�%��Kھ�7�7�vqhs�1�Da��@ЎQE�ܷ=M_����,WL�g��`�Y�M��L�f"�K���r��
��L��H�y�.5�A�S�>�hW\��8���T>��-8|t��~��d��pL�yif�7*Y�a�-@��J����ѳQ}8�+�����c��1�5�P����`h4%D�	F�S>�Bu�r��%T��x3�����ܮe����l9�̺�6��q }��{�1w��
�K���=�[��_����v��9p��[��+��F��pR|��ִ{T�A"<y�Bal3�FM�W=ۺ]�&�5�P�p��7��c�C69��C��Wy�'�t��Ԉ�1��V荜{����������K�8s P���%��3G$� [�X��@u���Y��}���Ǩ��Ĩ�m	���0�+����n��Ȯ�$��i:��B��S�+����uL�XdA<A.#7F_g`ʎ���5���9���T��{�
�ק���8*vt�9t׿9&�it;�,NN�j۴�bN�/~>��"��pOKȫ99���J��(d���r�.ʟa�q�{G����a��D�/�θQ�"��9ǌ�)���Xt#��o��}�<Pz �_��}k�{^Ot��znuD��c*H��@ŗ�wd.��$�"��q^̽�H`ݑz����F׽�ue��MI�=��h���pXߪ�s�.�"�Q�scf�|dc&ũpz�T0�紆�l�{��
�W����PNxˍP�ϳ}��Ŗo io�x�����^��ڧ�i��7�3�z�����{T��+��Z��ƅ�v�-��3o������=�;����KwbH̞�;���l� ��q��#%IQדE��+�)��p�k�ҹċ��Ur�����o��i�}�4r����+_������
�i,����:�x\{L�բ����Z+x7��A��T9wZVDdC�򎈎���&���yF�>�/����1��X��:�F)���tOl_�u#�//���L+RI�0x�1��YJ$�Bq����r��z��%C���h��u��vs���v%}���v2�!���֓���sP~�}ad#XF�N)w����������v"��Eb�����N�W7o;���Y���u[�9�����N��>JoT3%m>�4��ǰܰv��`�[��"Tc+��ow.w`6�Υ�z̭�ў�$��m���B�\�(!�P�'d��ٗ����؃	�.��d7��Z^	nہ���07#H��F:�qF:f:H�ˌ�WE�Y�����b>U���Y�?s��N\5P��Q	��q.�\-u�Xm���ج��c�`�X2H�ѥLP�[k%��%�\��ۮ�y���	o<�9�a��-6�|�g�	��χ��Q�2��{H֪�k�e3^�[��=s�����M$����y��^�J��h,��ga�SG/���3΃�Vy�Tl�w][�֎c�1J垮x�w�x�Mfr��a�wѭ�.a��F�	��&�k\�G�\��r|���Pא���&�'�]X��xH6�(�\��~I���i`�S�FT`}12�fMk=�Z�`r����T2z�`޹����%�De����X�9ફ�'\�=�w�s�x�X(b�v�^Ȩ{xS̈�K0J"_�*�/�^�ve?/YDȾW��4��CTss���wء�
����[/�#�F�J΂�=ˁ��gK��з m���nzOkcFQ�O�Fڂ���][�g�;��v�t_a���/�e_vF
e"�1k	���}��wDal.�V���тA<���[��^n=�i��u�հ�X��6��*���f��Y��b��<�Le�Ϻ���Xc�tDiP��P�$��d�������eɘ�4����Ku�y�.�v+6�އ��ϙ˚ ��鄢�����}B�VL��E�8��B�z#P���MD�"_����N�p�����'o=f�S:	:�K T=��P����ӕՎ���J��2��MN��8.C���	������*�0v#Ic���w�����L��f7�E����*�P���6�iF󓰲8��:�`ʗ�S�nB�%=���КN��N�>04�>�Ϧ��"@�u�M�]~����7]��؋hʅ��㛌�]x�G��ϻ`F�� �^2N��j aj�d-ΡO�����)v�r�K�寳;��\��u3Hi>�w�>�t�AM�_�H¨����9��
��u�ㅥx�C��ׇ�Xk$\�״�<.���6L�v�Z��S�B��>+e�ʗѵ(�r���y��&�Y�=0����]BMr��*rN���������Pg²�m�h�[i{L]N�	0��E�1�}b�i�F+&�.<�y S����3/�Mm��Ҭ���b��թrk�X���Sam��َɥ��JJZ�wH��Z���gu��c���n�F�3�v��wjTj��H�wI�3���ݵ:����R.�G�Y�������K#��@I����"�r�������V��ܺ��s�r��E�}.O{�܎��SF��Qeާ�59&
$#;a��#(iWF\v䴆$n��R���"6�O��c2���8b]�.:�+J���~�-��oJ©'�9��5&㨈�|��A;ˣ��tGvEF�z��a�&9�tI���ɨ	����o��8��^-���%�ܙ�X�O=��qh��v<��1!�1���V�� �#G
����r�b�e�Ju�s�8�ϖ����;b��a��5[Q� �����gJ�G���fVsz�뜉��!��:k���d*�r�p�-�n�^ބs���D8�� ����M��}��O|
KkL�.S޵4B����0�A�.6�j��P�|>َ�_��>�r{���4L{�q��*���*��Z7�U;����g��-@��J���%����,�v�*�6t�ƪ���ڇ܌c���>]�|�����{Ҕ��+Gs���Yg��cAT%�V���i�=�l��>�u�GӬ�#��U����fb.��/;ά����x�ah�y��~SOd�ZB���t����[�G6����$"��N����FX ���}{�k;��R��A(Ի�J�n�U��S"�q"=�q_l�/��!s�w /�ʀ�^LpO���� 8!���t�x�]�['<��ա��W�`��ϼZ��<!��c��1~M�u4D�����~�$A�FMŶn����j�uB���f7����r�j����s�!au�ׂun(۪�'� ��DFlh�N��;��@p�V���_Y���<j`P�Ì� c
E:7�F�Ta�y�t����T��mXdUJ�aø���w�RUTQd��nY%�=����d�֚G�&�D��HΦ�_FQ�U���~k��½y�>�.7�
]�_�l<�쾧�ﺷ�݇cJ�ܩ�X�{���ThS��N���/��n�Ve=�Ç�m�vc�I��ݹ��=�q��Z_��-�M�!���\7걟s�.�"�Aᘃsc������w��zE���%{�Y0��-��1<�����꽶ָ��ӭ�F���9{��W�3׏��c���K�ڍ7�JK�҉�U����	�q�T����@�k�3����s�����Z$��O�w��~țVd\��-0�1�B��L��S�Qn�v�N�J�.ZM!�U�����C����i���q�EQ+��wS��T��� ݽw�M�F�����6;:s�8Q{A��S�r9�9�}݄���-M����L�ѝ�6Mmў��C�*$����ɢ��°Mb�pȗƺ�+�d���O�i���:X��[�x�C@V�?{J+_	M/i��Ϊ�z�CW� �$3��d
f�t-����_E>m���û��.���
(I�EW��]]�|���7P������L�ԭʓ�|��������~`vo��//��vraZ�O)��َ 2�L�����F�]]��'%�@���\;}�&!��J=�ƹ$un�廫P���$Rz	�u0�JA_���Z7��`��@{/�ix�m�ȋ�[��U�B5�S�:%UB��͸G!ǝ�Z���"�$c�zL<SF�9�G���U�N�G<嫇1DPM߄�)�ҦW���\�M���|��}Z������(T-�42Qy�RQ\���t����j�>�돜��X�5|������|�~fiD�L;?�k�e3L��PDO�^Z1}kzpl���KC�Wn��"rVT?�f哰𩣗\<�9�~1��B6l��unĕ��Cۼ�Xh�@E�s��խ�U��kdh�Fc�	�ܔ:i�>G��g]p���6�8�S��P�މ�la�d�A,r��F=��j=Vt���).E4;+�Ǫ��]b�k����v��ڽʔkf�ձ��d:�k�j�����і�ȜXjl��;��NIs�F�N���]�� ��D\���r|��[�nc��D�ԄE��N�lF��c�U�����=�c�0>�f�m	3��Y��b c���Ѣ�6�i�A�P�LPlj��ꖫ&�߶W��v>�w{g�~���1I�������2wK�31*�"��Ft3UsY)K0hd"f�_7�]Q������&wތ�~���_?.�KM�F��_�}fDF������6�$H�D� z��yH�s<w}�>l�ko��ӟ
Ӟ�jڪ�C���9sD A0w>5��E��SS���`��u��&���E��K��۠�-S=+��V�Q��%�/���+>�=#y���1MD֞!��)E�2�k����%��ä#��ՆoЦ�1��TpJ`���.Q�;��̺q{$��a�܋���.��Ez�p�k]�9��W���I�d4�a��MN����ܫ�P����c���eh�[�N��S|�!��g�U����A���8� Vɋ����f���7�F�N8v��o�.�lt�]����v�'zR�v�c�*��6M�r?y��׎�|����v��Qs��>Ǹ;��&u�l�hW޴g:<mT\f�L����!��f`{yB<(����mkm�bSη���՛ɐ�1��q�`귨�,W]]2��S{�S�</r�][D3�3	�U�ܞo"��u�Y���a�7�d�M�5ǯt��r���y���]M�)!�f!q�n�J�K��jK9[��9N�����K%��[�>��k�ю-��8�n��˨���ü�D6�A�+^��t_b�`D��e��Q���!e��MPVa��^(�Vw4v�C7���))�_���  �)s̥��j�k�*Y`f��9�!���4�����A��_U�wn��ĩe՝|
]���q��r�
�θú��kHFe��0.w�x��n=��ؔZ��U���"���S���X#�r�v"q�tCӺ��B�5�H��K�oK����mЦݎ"�����z�	��8�i�fed�D3�c8�QU�ʜ�>��U��gr\�Uc�w=z���j�3�s%�	p���M�Ϝ����J��2����ٰ-ɣu���n��!m>T�OD5*��|e쥺~H�ʾ)##Y{�9SF��k����=Ʋ}������
���"�U�}9׎�vl *do<�2�J�3�[���k=>F�yL�F�r���A4��sü�!�ˌ���0g�!a�^�wHe��i��&��^�ﷇ3M��{��;jfeJy�i��ة���񚯨�נ�r��eSai�$|�_��ŭy�XV�S��\լ`��:ͻ�I<U�ǵ>8���O1����7�����U���R�u}m�WACW���k��������9cE�WIs��ԧ:�t�C���I��_v�������t��=\U��;J�gF+�h���r���s{�:�y�\
Fw�қ�-z��ζ�*���ug_Q��,�`��?��=\AQa�b�7N�i,ڹ���Σ�>v��1�M+)�0)�)�a�Pm�b���F�R�Fb0C�L3:��;�&�ׇE��;��;�����ob�y����6A�re�vy]��b��rq�2��H^�W)�h��"�&�u-�|3��Cq؛g����F=�GQ}X�n*Vs�ol�A�|;�,����]�k9�̬������1�t{��*3�+�7wH$И�g��62
ӽ|����z�|��'Klg��a�⮓�̺mm�y�2+t2�_6èoS�8b��IV���Ddw�;�ӊ�V�A!j�U��f�*ч�,�j���h�BT<��u�����V��*�8U�����>����#@` őX����hf��_bB�nmXYa��P��7��`'k��Μ�z��S3x�2�%Q�D�;��U���wq!�u$n�i�Ȋۣ�$����N� cD;�q0�2D�\�	A��k�s@˗d1D�	�mˉ#���܎"G.d�ˎ�6Www\��d ���#��fYsww0��]��Wwjq�`�DD�DM1J@D����: L��wews������E˧w\�w!�3��nNۑd�"���A���뫄eΒ��S��$�v&r���F.�w;����ݻ�������$�W)$�`]��L�4lIL˺�	JcD�N��Lr� �wn)�2�wk��;�1�&��!BP�)0�F�q19��˕�\3��eAL�B�|(E'�;>�E1�K=0gs�Y֏C��J5�[��Y��u�����a�et=�<O2m��NZ�9$�A��0Nȭ��RW���ԁ6���<	��^�ߚ�߫��^�?�פW��^-����cs|+޻�J�so��:������y��_m��[��uzZ@��_�e�>�"O�����}� }����]}.vL��|*P�`I���|�<��W>�x����կM�ۻ���~W���Z7���5޻n.U��U�[����5wv�����|k��[��oJ��_�x���-��?������PHRf��z�OclQ���#�b��߫��6���ϋ�~��;|Y�*� ���D��r �=�"�� aϠz��_޻z_K|{zZM͸m��׍����D� O�L28� |G��_1���膣��}Z�~l�W�iO��d"O�<�"I��N�$�#��|-�@Y�~Ni���	"M�zN��{�=��r�|>u�*�\�o��ט{�\�7�ߞ{W����^�=��W��S��2$�NU�;_vQ���bO�����T2+����$��#�|��� Eǳcޣ�G���r����x�|5��a���kţ���[_��x���m��ln>��`��@D{�����l{�@D���o��7W��`�ε���� ��������_�}]ס��r���˯��o�/z����>�|^
�>G�z2�M����}�@r���(�#��o?�޸�z�{�$� f�lF�­���<[�Ä|,���,����k�����_>yoM����������{���_j�i����K�oﺿ�7�n�ڽ�����s|}�ۗg�<�F5^�3�< �H�k&��u�43&bN�����f��$B�,� |��>��A'ޕs~�>I�����#H����ߜ�gȁ'�@D_�{�/KF������ƿ����u��K}�����޷�x�~���qW�A���V�����
�:w��##;�7��>����t=d��G�����@��GC>�"��}�ޢ � �����|���7���}��I'��܊#�}FH�#�EG���#�d��qG�>G�.�Y��"O����߾����9\����Ex�U������lno׿<��opA����Y��=� ;�sdxHgގ��� |@�<�����	>gރ�^�,�7�oo��}�yW�����^���ſ�p��-	�[�2bU�
űs�kAkGR:����h%�~�Xm�F�m�r3�yr� 0ttܶ�X+�6T�6=��;�G*G�YCts$v![��T��W�9��6��N]���+�|�!9Tk6��N�a���[A`=ppL|�u����ٱ�>����S��yzpHWޒ@���>�U��E�M���#ނ�������`�+��<F�u������Ž�WϞj��Ƥ�F��@da���\��@��,}�Ӏ �$|}� �{�ݓ;�*n1�ᓜ�����{O�z��Ǽ,�q��  �Dy�>�U>��(�`� 
>����y� �s�Hdy�>��x>��A���d#�z�ﾙ����u�݊'�1�~��>D��H�C�4�&���{��[�޷��x��w��*�\�5�w�_��U��}^�����W5�TQ��B�����>��A Q�S���>��>�|�����g�G�3z*�ߡ��4"Ű��d�Y�F����#�d���0��0�}��)�8�>|Ȓ7�u_���yޖ����s����\�_^v�ޛ������/KF�oE�}c�0�P#(�/�Q�$��&��ʪ&��{	>Gރ�
=dQ��d�O���Y Ax�ȉ��P�=:G�D8}G���.�ޣ�@	>��DG�?�F��+���W��u�����|���I�YV�6�o��Le/����}$Q�>M��#�$��Yg��$����}[ A%�Ͻ;�PH��>�L��~>��Ȍd�^@��=D_�
^�x���s��^�z^-��zo������|-KȨ�Z�U�h���|4�毛�x���^+�n�����|W�x@��H�<	� rj���D��T�D#� ��+`y�$�,�>� "�o������I Y��,�Y�� ����)N��%�9/�@���q��<���>����������G�ȅ��I���zH�>���J����̏`t���QG�6��|>#��|^+�������_[���֟]�G�Y_5�&���W��?3�6G�� �#ﾟ>��q�I���(�|��:�^->�_=_����ۛ��k�z_}�z�ɏ@�:}�_H�<	���ۯ{ˁ����ވ�y�"����0���;EK𼼭X��dT��>��ğ�#����'�i�o��9 Y 	φ�>�zk����w���o���ο�^-���Ž>��W�}W�ן�\��~5�t Di���˯a���}԰g���k5!�b�����ZŃ��t�s�e*'e�v�d9R�����0ez�u��񒆷B��.V���w�5��;p��K�,ZM�Qre�Na��6�����8����ל�P���T��oW
��`ym2��PVm�Sa����2N�7a��uNBqn_as��9���ϟ=W�Ϳ�z꾾z�7�ܿ���z}_�<�齶����]{k�\5����z[���_�{����\���._��^������}������׾�i��"&�]J���`Vrط�.�`�|<7 {G�<�>��A��U�$3�ޒ ���,�z	�<`uY�|[�����;_���r��:�^�ޛ�鯟�zU��;o����y�ž7��{�@�l>g��F+��6-}�g��m!Q_{>}�I��>g�'�O��#: I���>�t8��x���+�����[�\��z�o��~|�_[��-�{^�8����� I d}"6�zI>��F{��Y}�2}���>�e����]X>{�&�}�" � ���DE|#���(�����h�}���DQ��>����W��" �I Z����� �=;�����|}7���~^�y��-�q�O��#ȉ#���Y�0�K��}E�G|�d}��G�����}�� ���\׊�.om}n��]�x��s��_z���o{�o�z\����[�}�zom�#�<�C�#��A������	>$�E�#�G�#�$����?(8���蟠����k��|�G�RH@�$����+��_�ƾ��^r�oׯ;��o�y�������_˛����o����r�v���^���R#У6~�y���}�>��ڇO��w�j�iux0y�A��|�,���Do�8I��||����a�>gfg�L�	>dI��8��#�$I��n�-�^]�����ݯ~��2����}�8��Im�mҷQn�b�;bS_ 0�#��F�>�8D	#��
�zI>���@� � �}�2s�}� D>u�a'�=�x�GO�DK��(���,�"�@O��� }xH��ȒOæ��������a�=� I>�"�>��qG�>�0U:���$�`n�Ũ��I#��뺵�2E � �t Uu殷���d�`��4`7��6�֗��������i�[t#m�<X7���O�V����8�vd�ޝI�Ӈp<W�}C׸�Q���ݔ�Ȇ�����ͱMu^�����b�{\��S�J��/l�}f���foN��v�j&�8���JV:铴��z�-�nD�����U�R�s��������j.D�IΛ�Yh`cA$c	�٣~�3�a���\���9j��DQM-��sy�)��r��Z�Jsz��R#�( (֜E��i;\<�v!��/��kH=����ٕ�ku�2���Dsq<O<�a3�鏝r���(�i�c�K��3�k�ժ�J�*�|��v�z�T-���ɳ����NY;SG,C ���}#f˞��t�XM%գ��^Ҹ_�^=���uH�;��F{W�K��PH�	�.Vy�JO*�*1p�/�h��ܥ��VK���OVMV��=�K(�\���LW8}2�r�Г�ȳ5Gt��Y�ȧ��f�+DK�+�e�W�8���s�c%>�}�UU��9�k�q���BM���C���E�NF�s4D�}���,R�`��Dό�,\�w�_�L
�h��^Tm3���@����������g��x*���}fcdqf:%A/{i�D���6��m�5�Ia>�Jk@�L��%�;�u��շ'�\�DtAJ2'��C�r���}6e]d熡E��06OX�Y�ǫhM��b��>6��+7�G�V�:���W����N��\C0��B�O���T��eN�+`�[��,*}o%�C
8wbwԻ@j\�NϮwmk�6V�A��88��ǜ*e�H`W��{�M5��!b�j�P{]�{��ѻ���� �&�Ξ����(�\�A(�Z�z�]�Fw,F��tu��{��t��_�dl��Bb�d[���T�<��Q�^���g9.�x��Նnۇ�;:eE�r���R��F�m���)l�=D�e��w9*ds����^���6�iF�e��d��ǹyԇ��#�?S��F�����'�D�2`"L��>�����2a.�9Ӊ��6��t�t!Tn�!��GE��>�'"PPAj��t�%D���΃!mgX��f�%i��w���β'&�!e5�f�4&�I�S�N��M�_Č*�����9��D�eʮ�S�&�7������0�u��K0o�&S�fͺ��]���u-U��gY�tY��{��a�_��o(�W��C��Q~m�<��4���&<��:۾��u����kn�z�ʬy��g{U��p�\���:)x}�O���g�vݳnb�z���k��؆�@��h���PUc���a�W�Q��eE�loS��N��#y��v$ǐk�_�st�HWݏ��m>�;��]C�.��5���V]2��y^@��^J�WJ���b��( ����|1�z"W�v��Qp�3;�2^���#|V���~9#��U�/*8�_+ʆ$��`�����rH�/:�B]ŻӨ坩x}<kX5�L�51�O����
�C袎̔Y�ˠ�� :��",M���r����&���=t�NsDGE�{^�����j�#�=Aݟg��Ls��2�t6fs^WU�H�K�]�ʙ���E�]8��/��eyk�F���v�$*���|N+�����e0����:��{!�"#y�88�d3��f�v�cU�r�D����W�r�/tx'R:l�׷2L)I<k 3Ր��!è�ܷ
Z�o�8�A�]��W�.o��_nz�f�>v�<���
��-z#k���B�r3��#�Q����KC���f��9^�2σ㤞e`
����]{Y�.y��,�vz���f�M?.7[��!p{ܞ�(���O�P����`h5�J��!�Qu2�ӶggGp�sv#oWy �q��g�k�hq�@�RtN�_��')�f�uR��J2����Q8ԫ��]�LNvFP��<]���'IFs�%�a�M��P	<.�Z=�N�+==��rC ^���m��I�%�!ܳ�5};���cZ�Ov+]���{��Ɩ�?�R�ͫa�f2����������.$[[��W��ֹ��:Om��p�b��XT�H�A�ڃ���f�:��,;��G���'��;6�����㽢*��  R���T����7qdW�9B9�E��
�u��GK�Q��&�M�8��My\��@{5�3uΧd�CՉyX���� �p�4���.��Z�50(rN��p��1d+3NPm���)W�9�@΋�Ϲ"+_��4�c�7�R�*�rs���	+�1���E�v��b�蝙�$���hk@��>Wl�,��y]��
�b����i_*��$��[��{�Sc��P���C���9b���=�F�?j$�`��s+�e=��iw<�\�t8��Cv[&H�e��W���<fa�ZN��ڦk���N�I��\����[��v�3[����Jϩ�x�3QS�+�Z{Ĝ\k��uL��>�ȿs i��<n�>X
�)����	����̖����L�F�%��D�*��<���9����5�~�}LZ��?e�Vff�|�L��,��f���r�����ɢ�����9�#8S�����2\[�]uLr�q��ߩ��D�����	������3��
�$h�.�Y�\0�l_Gf:ʉ������nd�,c=~�q5��+m+Y|�g$9��h_8(s.��˜s,Æm��3��|��)���v�6"Η�p�����3p%�t��{k�'�f��������#䞍;3���Y{�~���k�����r�4��Ąq��w��r���n!F�:I�E}D{Ms�Wq�V���R�u�P�4��\Q��_)Wk��m��A[���//��vraZ�O)�Ć�	ޝ�6�d�o�13��܊�D�7--�7�{"�R]5�#���z��<\��{�	"�m�*�&���bd���#�qBؑ|�K�-�p2"���i�n�l�7{s��.5}��G@�e��>�h�Z�1���O�x\��������p］��������ؗl-��t��ޯ�Dt��U��\�Gv�@hD��-��I�ָy�^�C�;��X!��[��;�s�i�<%�Η��?�r��ʭ(�i�v:t�^3=P�����5�	���H�o/N�]E��f哰��M�b�r��y�Tl�s9�T�i�.qdM�����*¨�큇:�,��=��.b����y�s<ť'�Z+3���CVYg�K����pV�W3��eUns���/o/��@�bb���k�Г�#�<S�I}L��+��b�u�bqĬTv���3Z��U��Ⱁh�*���<˳� �9�oo<��%9�hj,`�¶���'u#���ӄ��T�a��JSo:�godB��ج���S;:�׎)&!�|�鬴�����Ԭ��{���W��4�>7FD�Q�nb ez�rp����%NDe�f��T�����F���ꡯ)��q	�:�����Wx�X(b���-�k�駆������8��4�Īܷ'�v�8���&r�,J���N���Ǣg�c�p�=�����Z��ഺ|�}{9��n��m&�V��=D��&V���[�G\��p��A�ۓ�랈���J(D�z�헸$�e�oq����xZ�F�P2�X�tMd"sm�n�T�B�㋧f��]ی�����ɻ��xK@{�ur�C:G��
2�k����%�����כV�
q�xOUe'�keԸ�t���EFɛ��كDF� ��a%"b8�)*�TwZ��~=��Oe�ٓ�r{J6/gj���UA�>��u�u�ʕ� �TO>0&cg�Ma�D�:�&��)��A�m�7��[�玴�#�eO�ND8���I�>�B:F�6f��u]o6o5��S9���aa�E�Ӷs����9A7ZM�ռ~�2Q�tWE��"��1�,��������_xM�>��˛&��GlGװY����T��Ŕ�pm@)��n���+�WQJ��&���N��髉|�I���k�Gi8�9��Pj������B���B��ܒ�m�[(p��2	��y�-㛙P�'W\`�Vv��������m��3�������C���q��8�,��
8L�v�)�u#A�F�T]�I�K��i�n/�rl��leC��ح���]Rk��Pےu��	����#��D�����۞�e�n׌^�˖�z��W앱�WAjN�c�(��9�� s�8�1�.�twsC�B=Ca�5����Uc����+񩇅�l�?9���ԡ��c��+�v-�#L�:���n�1����n�-�>����E�W��+6ii\_�ᅇ�LXN�9�sDGE�׫��]ƫ��P��A��k+3��`��x}��ʸ|�b%!EDl$�����2oЋ:�q��#�O�%1�".�Vו�#�ine�K�}P������j�������B�do:��d3����F�ƫj8��$'`ز�i�X��Ad1�^���0���/j����xnY���C�Q~n[�-W�v2�	��{��*׹j�D>�X(��u��X(W
���b�_)�jh�`l:g׌:G����Б�srR8՛�^��4ȶ(ͻ,��E�.��v�$
Y�v�TWvF�NB|�vB�l��XT�s�7�% ���F�c�g*��8g�@ax�K�D�n��5�^
!�3ѻ2���*������� ���K�Ɣ]�Ɗ�&`���T�#s��~I�沂u�]YIR���}�R�	�Y��X ��Z�͗@c��C��p���DYȏ]E��)uK5m��a2.g!���5קh�-a�Jm�-&)��"6�'��f��ɬ��!|��P�W\�r��cy��ŕz�`�!�7�д�En)٨(��&h��Q��'���a��V+�r�ܤ���6���:�sJ=��5��aZ xn��K�4�tiF���m������'Ďw&J�΅F�r���5kf㹼��9�.����ǳ�/vji	[�+z!���6�.��E�}�s�.��C�J6r�v&�.��z�{wt���#�E�m�\�o���:������ۼ��7r���N�VRHƨ�Ѓ��u/#�5��9U�j���Y���� �Cb������"�T�l�{4�  |Dc���R�-}(ʇ]�����}�ܧ�����'>��0��۽��k�ַ��B�t�[-a-�g72��p����	�h`^[�9�h����;!e1]B�	+x����,��®�ם�ҩY}��\d9���Gf���!\5})��d�Gυ�2��L˫U�+U\�(�Za)W\�����Cs��	����ݺƴ����%�FT��Ü�L�̡)R�t�� ��l��B�4cN��r����fa�Ӯ�z*c��Z�\�M��/1Q���ȁ��}�^�Χb;��5�3��ѵ׏��/��=���,��[�y�Rd�����y���(�zfޕ��=Ii���q;6s�v
ڃYsrv�;��R���[��W�5E9�V��ؖ�]�ɃE�5j�dԡ���[Z�{�i��гV�d��1��C�-)Z��u]�W&ԲQ|��Nby��t���)�cs���d��N_Ŗ�r��D����F���{���c�Fa�w�#0*ex{����vn�f�03���C҅ۂ�Y�B��]Oq�D���=�J's�P;��]�t�7b4���f�Fn��%�t��ĸT�ܢF�lR�-��=���;v�>�S�;x6���mGE[���-����!�/)vG������W[�Cm�a��2���r�X��Ip�J��nsU����m�|��^1mu����+��.�N
tf�ߔ}�+�ˠlK�;�� <�X�-��N�mf9��m�m�}&���:�[,k�M"-9-4w�3�u?�.�2/K�VqT��}���,Sk5Iڷ�z��,��(�֪�:d�unou䧶�,*��j��|��''_q���5��9%)p������Fu�Wwn�{�dAhVwa"Y���<�\���0)#$o�d�.�h&%,!wt��(�dFr�R ���b2S(�(a,�(�I�K3&�CM"����uɈ��;���I&��;\Ɔm��$��'.;���2F�2$�)wn�.��"J;�h��a(�nWb�q�;�Y�4hQ$��"7.LaD��v�Hs�D�q.�afs���a�A���D�2H�$	wn�L�""�]5�wNr�D0I����
]�4�M�6S	B&H%L0K����Jhc��is�롂e�(�B��w`&&1B�L�.Yd��$��`��� a���ϧ�����={������S1`WX������p�������X�@���2gl*�RiV�bn�bS�$<��6�$Vt4�O�ꯪ�'�}�\�d�'�8���!GDG?��U�<%4����Z7�S��!���5L�c$v_N�v��UsgKl�P1�Q���v�<�F�(�#A�BTMz�Y��5+{Sr�\��QX�,M�;n���	�;���4x']�ה� �JX�z�݁s��!J��y
�B衋��b������a�M�u4D����pĮ����y5e��D�0����C#b��� �G́qD,.��ʩ�ִ*��9y���p�����n�bDn���W�p�4����ևqБ��u
"bw�+�F���vi�"��*�S��������$Ek�q�k�Ճ��kֳ�<~���_�,Ǝ�{;��̛�,8d��',�����5�.&8՜���o��Hu�)R�hq�H����-��+�
��7�.udbr\JE;6�"���"��b#��,��7t���NI���
��{z�o1�3V:�E���I�!�{T�w��D�`|�d{ ���֧�Ñ:t.S��������^"e�-�=�#�����^��`��zy|8E�̘�@��*�"��W��MAq����7+Z��ʺ�3�E�z�a�3��v��|ZW1�6ܝ������� ��$t��*����C����E�ͮ�}R�J���}��W�m����x����b�kV�Q�#bǶ �M����S\����۪dv>���5"s]JͨC%��f��p��%���t�f�|��`�2����������p���eG�]],�o�ި�s�z,dwF���l?&)��;*�1��΀W7Gt���8ˁ��5k2����F����M�4j��iEk�)��1���F?W�)O�6ڷ�v�w1]�B��c^�w�=�Hg,=�_:�=��u�dFD(�6�}B��W@^�8�ڗ�q�~�����d}�T�Q�\IdPī��>�2;�kᶽs�A�������؁���Խ׳.�\�,d-�z�\7��&!�Д�WF{\�:��pr�wV�mt[���۫����17&HcD�Bd��6`s�"�Bؑ|�K��D^����i��پ˧�\�ݣy'��M�"�Wv⍉�P�$v��<�h�!��G�;cʽ��(�2q�,Y���XW���.w:?D؊i߅4�)�柙���@��Ⱥg��\���8�����u2/b���ô >�0�xy�A�F�.��o���YL|B_=<�4�[W�xDV/���v7Hn��v�r�1����2ȧ��U�3Zb�����R�*��e��usoѴ��"6T�E��b9]��vΨ���u�T <=�xB�㋵�f�I���s�	�臎%��{	��W(��҉��v:k����%�s�gw�EX�3�0�3{-��B�Ά`����*h�� ��A�+1���Kٽzj� L��!�ǉZ*6�V^U2�k�3����z��*��a�_!�o)����c�9w,�(�$Yb*Y�C�&2�s���YG��^b�˘�q����[�kwgt[�v�F�]�XB�c�3q~}10�{N1���R�dܵ�;����(>ɪO`�l��\ N@����=��t��+�`�bw�w
�*��n'fS��C�<���s�d:j5�ߟw8f5��Y�(�P?{���<�Y��x*!���d+G��{id�s�j���Iy`<�I������,��:l��]~�=[ssD A*�wfz��|0U�����*3<�0/��B8�d�=c�
���B.m���-S=+�%;0;u{q-��us����"�����9Wz��x��g�YFTM{�����g�uW_��>�������в�;�����O�����U�J<��7�Nz��}�u���l��6�'0[��ӆ�sY�-�e�j�(J��YOX{��v8���v���o��l�u*U�GF���]�[y~|��6��ǻ�Mk����kfu�*����k5(;-��EFE�b��{�Ji�*P�2J���\�^2��*' T5h,w*�*��>U�BP����䩚��/�7�b,^��O��N�!�;�.,!��όI;�hG_:�$,�x�ufCP�s�����=nx�s����GE��>�'"R�T�tȄ���4�5���8 <B�'e+{��^��DhwyZ%��9I��oέ�
9�	]vK���PL��S�k%��[P�Fln�3"�b��T��q��+����]�<���WK���B��Ie%�W9$����vx���ʎb��q^�����)N"��tO0�ɀ�+x���%�TWvc�.��%t���5C�����?O�w��*�v�.W_�ޑ��_��Ok�b�Ab�����	23O�����h����`-,���0שN8�r�Qe�(5עc���z�;3swa�tLy!�ح��m�F�"6���Q��
`>����1�5l��B�5�kԛ7[��F��WA�%F�����9�#���z�w�G1��wn��Ytsڭ�����$�m�9Lk���⭽x�.a�sk+A�s<��}㝷�I۷�E�U��v�ct<�*�r��Na>�����Ɓ��RO}]�)`j���nĶ�%e޻�6霢&��)�QR�짛��RwnE+4�#���S����YO��3����������/s�]&j&�a���'����yUPdߡut�ok��{\o�򶢧�����u�>wn���'�b>��T��Ɗ�E�P�PL��\�C:�;���s9�.�ɑWP5�C�%�ol6�dgUF�y1�+��3�ة��.��Ɔ@g�!P4#�C�P�7Y�6q����g�#��5����5(�qu� 뢼5�(WT�����s��<�>��=����o+JK�6��U�W�s�f�y��W㤞e`i�U���o���2Xj�oo{z^ߨ���E˖p��e��J���	۰�� �r���ϡ*'g�Nh��]�nE��|,��Կl�5��j\���|�w��7��e9�r�$���r���6+�Sv�T6o�_�e�5�s�a��(b�\'IFC�!(�9Xa7Pw���$�ʡ�n�Ɇ7��' DF���1�7H��q酰��;#b�]mC�Z+è�_����wΦ�;}DF����qbkn�jD{k�W�p�4��y���d��O�{u��]<�}"��v�{A���0�奏ZN(V��;v(���1ܻ�R��v�W�
�]�.H�]�P
{�ռ|zɝQ]v�y����t���`����M�Oge��������M��<�~�}X�4V5G�(ܩ7r�V\K��p�\����ӿ�� �=A��aC��Q�Tk�N�w�d�^g�䈭`�4�v:�x���ʎ�G ����1�B7S�,6��ߜ2T�y�d�`���.��sˉ�����C��$��H����M�#��Ղ��Vo8*U_y��Ht��sDW1u$P}1�b�覞P�r�d�����h��H&*݋�F-F�^�8`��I�!��S5�?}٦���[t���ϻ�ٳ�~����{�{`�az+*�,T7�`l�{a`���q�9��GW1��i�����olw�/�!����]��Ö��n�/����|���L�>������{�!M����Ƿ���#$ླྀn�=��� ����Ep��XxG��:\��Zc��{��/}�hW�=�˷(w���V����S�-���^��>]Ԍ�>��e���K���o>&��f�,9���d%xsڄ�r��e�w��r����ȅ���1�9Sz)��{�,:9��57
'Fq`�7WC|G�W���e_�������V�\��U {T�-�K�3S_Qm�O�N9�*U����]s8u�7I8'%Vq�U�o���ngx��~=U=V1�h��F�>���/��n�j�Ɗ��"�mV��{/B\D*F`ںJu��:gt7C��<{��¹�/�.3����m���� an�{�5���c	�c��h�L�=�N씢\6���W�i�rH�����T��赱���´9&�#XN�"��C��vAJ��㈲��:��[��dE�-���' pع�'������^�y���'"���H��vA�{4lR��Y�z��<�����"v���<u�95eO;�Q	���ӱV<�i�X�)Y�x�F�1U`L��Ǜ+Xں�Rj[�M6��f�_9�6�8�O1>�s��>QY�
��x>W$���n�כ�T��&��j��A�9���Jj��f哰𩣖!��g��9���m���i��d헭�eOz�t�r�r7�a�^��9�d+�w}����($m�N3�)O���ǟ+o3;�ʻ�vC=�9>u�u�,
���8������`bbuŚ�gcP�)띛99\�K�����Ug��I���-X����곱 �,뼭^����mO]�uۭ(2��ݟg)އ�i�-�;[M\M�w��
��Oq;1��#��/<��S�����FI6�\U��/�M���
��a�P޵A��2���4�ו�k��;ڮg�oB�}K�f'b�,�I]����j��vhS�:`�|�470���+.V��{(�+#V6[�Q8��)t �fG�i��d򨩱�Դ'X�/�}_UW�S����P�07v���*i�9.����ٱ���޵�J2'��
��[(z�K�t;���Q7�ciFI�o*�������~�~��sC 0�qc����5�8}�p�}Es��[����եᲰ��B!-�nZ�{��8"ɫ�f�<ݤ3V��*`I��3����#}0�(�Q�C����{HG&��8�N���Y�U��G���a��u)��&�O�)9��U�	C9v��
{Z������y�{�lqY����v�K�A<�'��dF�zf��u������"�yEؽ�af��Ĵ��
�<w��݈�T�Ԝ�qJ-W��t�%D�u�=!�Y�d��ק\����2Ρ��V�zW8�aȊM֓n��
9�	ZpR��װo��8#�;n�C�7x����(6�<qZY�e&|��1UF�9��#b͸2_C�V��b���@��,��Q�|��������9�z���k��Qm�'�&�/"�n��x<xZ�P�k��X��qع�ɡE�]�t]>N������B�<z-�Ŕ�/F9���q�0Q���m����!0j
ty<��Q��ϋV2e��ER�l�ۣ����)`
���%�£�WY?�'�:��Vu�OS-\��$�h�f�N��7�xxxm�ڋh@�������U��S���m���;Z�/6\���l����xWR���^�*潱��3��;~��@����jB�20�E��8�X�G3DR�ՌśND���Ǵle�=�}�W�� �$#:�	��yUp�"#�O��c2�U�/���Μ�	ɽ^��9h�����}�LZT��{���~ǵ�	���ݰ	�3ʹ��7u�hRM"v �n�L���~���-��b/�;S<��z�<�oX�^�y;0�9�ݻ s
��jV��W��X^ίM��2�����Z�.�f�\�m]]}fs�2��LŰ9�˚=���5P�}.ђ�
��[��۩{8�r�ו<�q��gk��A�������T�u2�J��v�L��k���څ=O\�NU�0�_����{p����B���tW��@L%g�!R [b'�'B�ș�ڞۃ�[h��1��o�Rtޛ){Q��\�䣵�w�����>�u9^�Ld�n'�<���;�v�4��G�條íWU�;X
革�~��;�������7��U/6��W�s��F��s���|a��ˬ�2��
��>ÊT��������w�b@fT͆VZW��B��{�{���bz��;�=�WB]�S���ͧ�2��ד�z���A����:>f��o�*�[W;��1����j�_r��~�z�V�9�J��g�a\��p�T��>f�L���A}"�aW�sV��p�&c�sN����8u�}��i��w�t���|���ۃ���J��'>��\�D���R���ɹa���1�A1#�ۚ�x�L,���k5"棸�m �Ksݴ�p����o5�3�SI��ʛ�(s�Ɩ׊=ˈ����N�{�0��^�#��󮱉�甧S��b�>'�>���[o1��VJ�`�BmeJÕ��VV��yA&5�{.z������*k��CnTfh��w�Ba%��v;n�ߝ(���9X�M�W�<�����-�3�0�q�[%OV+ď��o��c����x��Xqnuzm.�Ft�U9��P�|��Rs��݌���LU��Q���g>�GO1ȃ��WEg�W+C��Y&�Ї�4{�Y��68�5*J\N��X����N�',Y�j���Q�2����Ϥ0h�\� u���Z���M;̊���Zwk�����O0!��+�f�|:��ګ�Ў�{hwqY�KAR��2�����=Vjöz�A�p7�^��Y���OH�x΀�e�9�J�Mͺ��u�����ݚE�m��0���B��b;��P��+1�Ҩ�����2��|�ě��q���rΡ��5�ܲjf}�x(.���W�j�8^�اO1��1�m�rvd�;䣐`N��6��g]Y������ZEQI�j�]�vewf%��3F8���/�u�W��T�st��z����s���$k^X�N�޺k5N�z2��h���SQ���A䳻ږ��wQ��J���p��x�d��p璍F`����슍������������Hʙӥh:Zݶ{W�s�aC�m��ZhT���<�4V����h���ۓns���Y�9�E^�B�;Gz����r �eh���M�7�4~�ubF�KE_Mt~d���z��N�D��PG6�e`�ܩK-Zﶞ�ZT̸*oo�@�f�kO�Sڛв䇮�I�#�����/���U%�:�S$�\!�˲�k����n�{I�QIZ�\9� %�a�I]5��k�MoX�s����ch!Sr�[R	��-=s�ft�Z��ڕ��*�9���W�҆���fr�� c��Tz�U��������jf���3i��5���Ӳ)<"����;�;~�0��7p |:ƓK�T�o|��o��q<����U��Qᓰ�oA���1��'&��1�իnCr���,E�2v��u:���j�G��n��8L�ƺ<��ޮ�`Y Y���)�L+�Y`#!�G��8f�R���Qj\���Gm|$s]����{e�?Pއ����y1��Q��vӊ�C�k�y^��om�p��u}�_S��ti���<X�[�"`�pI�L�y�5��;3���9��+��r�E�ǥ=��ƱUo	�k+]�uƷq��gw,N�*g�yP	�Pj7���%��Hǂ�c+H�o!wm-��K�����o��҃�x�b�{�X���8�Rc�.�n_ch�q�"�{\"���iqͽ����$��83*K���V��uG�]Y�7�����XآsU�uē՚�m�w8��Q���I�P�.�����e"rQ���`Q׉r�e<�ʻ��oL��r9��LƝw	�*u��n���V��,��we��f��v����L�m���&
��U�d��a�4�J�Q.��ż��0)yƕ�vRd��-$*F������W����8	�����U�{��ڦz�Ӕ�/�KJlq�w]D�y�x ����+���uU�U�f�]���o���<A��|�{nF$�E�!&jc;��M��
ɑ3(B3I4�Jd� ��"c�BJ��$!
L�2L�Bd�$�"ntH��
H�la�F!��JJ4f2��*!2�Ć�c,IR�	0e)IYΑQ�b�bK#
 u $b��2�fPH�s��L�D�BB���h�	�30�
L�FFL��%9�H;����w4C���DE�(	$�a�E$��0ғh�D̤F2��P��
 $#p������_"y�Cz��S����uft�WA�Q[ӷj}e�Ef�b���d�d���K\T��jQ���<<=[\ecJiɜ���G4�%�m���c[=~g��+�cUK��J����o��	��:X�;=V���)��/�}����\OH���|2�U9W`���8���jC|������F���~�����Ņ}��,�P}��9�y��;��0�_�)Q�;�b���o�؇m��`��V�#{.�Xz�و���"4@q�RU1��%�B촱��5��kE�H�4�#]�ԣ\�h�L�����
B|w�M�����6�aW
�s%�o����L�U����>�N����j�I�6���{(�rF����u����ͣ�7�ĹQxt�FǊ�1�(�L7h\sټ�X��U�R�zs�%�i�Ų�0�$�Snk����B��Ȗ�..-��ɡ;�41��W�Mx,�f�c]�7Z�T�/¸��$ۋ�L�S�]M��#(�)W.�~�����;�3��F�K��+�ѣv�v���ܫ�O������7tgI��:���7�O�b �'��K(:�G+�LL�Tgr��[�M���G�2��3'����ۼZ{<{��9�����x =�moCk-�Ȍ����o���۞�,Κ]�uxba�<B7}Bp%u�cr����F���P�����t.��]�]b��;s�٫��q;֩�񣡍N����#"Es	OOX�;A;ɻ��s(C�9����Xo!=�f�k��������r���ֽ�<�藴�� ��x�ۇC�i�K7m����:���:W1b���o�6���?i�������m�r�6�U�D��FK��%��C�����tۆ��3�����d��C>dr�{7͵&*����A}��*�d!7ȧ6m��i��U��T�{`��*Lgvdk�'�F�+���z:��k\Om�F�\�H1�J�=[p�r�����yW����;܃��4-y���˕TM���]�^��h'M�܇A{��E/o>��H�bT��P�<����b�Ak�Y56�`�ޚjE�>�Y	N1����C���3ua�q��륙W���WE`ZڝO����;!��L��'%��.=��7v�l�D� F�,�Գ(��W���X�h���@ԧZ���þ�Y,ܶ�UX�JR�B-m��ʄ,򘟽�xxx_b��=T�6c�9v����[����l�S�Na��O��u8�v�9uљpX��A���l��}��riYw���I���Y��)�,i�z)��[w����T�̿��ar�<��ٶ_�\�B�₼�V����.Ձ���|{<�}���\$�T�$̺���j��a�v���S�E�H*&(H�nz���j�D�Vw�m.Jf�aRq���@߼[�����Hl$�c�jr��b|\GW�-���^d,y�ޡ�(�'Ur�طi��`s�mB��qO)Nߛ��w�v���o�]��q�X�@�'��仺�RY�6�r������=p�{���',5�w�s���ʓ�s����U�T���nr7�h�_>v�1~��vy�޾nCx���~��Ō��������6D]�1�
2{؇H�Bw�1p�}�7b���EH�Qeۨn���^�jx�^Z�l<�`���*㣙L.r�\q��U`��y�D�áfo6�`�k�~ un��'�]7BN�l�����c\`��wl�KH֖����'�nrT "L׎���P���RN��v�uk�����荒S̈�uv��w�6���:nK�|�zo���GHu]�R;;ʞѝ�������픽���o��q=0�W1�S/��AGJ�n�+1�x�9����Fz����>W�i���Vw!R�Q�^/� ����E&C����E�����l�]v�ܕ�Y4��r��c
����{{������2�EǪ�񶠥�+�EK�ʷۉ����A�)&W8�O�;/u�br"5��946+�S��{qT'�e^��q�B��=Q8o�x<��� ����'/$���<�jV��_M�¡˚kr,��WD��xT�s�S�y��A9s�t�ђ�-s�s1�q���՜�A�z�!qU�j��I�`�1�X�&(O;sP_����0;�)�7�O�`a9�f�$���)M�|
���X���p���>ő����j	-�lq�
�֒ҶU�ڇ�ϫ�PI�����X��+4�-,b�Yty��L��"$y�9����x�s��ޱ��_J6�	O��gj<v��S�ܗ}m�.�-�w�:�h�LP�Vhڽ���e,R�z�W/)�pU1)����wu�v���U�}�sG�e���#W�Ɛk�|�<~s���L8����k���U`����3y*F
W�;�(�6�n��ڛy^��s�YZ��^XI�oaΦ!Nmf��)���:3�z��u@�P{$]ꚛ8�]����wӱi�KNr�'>@O!gz��H��-^K��v�9jv�ŵ�^�K�,�JsT2��[�����z�7*�����m������M�rcUK�h@�7t�ɼ�S�z7-&Dsw�!���������9���\OL.�u��K�a,�zN�}�7:����q+�������}`B�W��lwd���է��]��:�h�m*c�	��T(щ4k�����o�XJu�yn�7��Kf�VB�s�F�=�|ZPy=�%�P�bV֬c#�V[�ě�Q�sy��aS�L� ꚰ�t�ȍ�R��B��z�}��X���Z�4�z��R�gL�`YF�}��w1�;�����l�e��(eNV�|	x��^ 6��v������_�I�Q�,L�����"��H�w���g(�u��)���ڌi�놅��)�J�4�]�d�r�s`�	�ᩈ����&��g^�}U�}���ۇm�u�97��ۀ'�k�����C��ڨV���g��M5���!:�h��@цҎ��V>.ÌF�z(4��ܗ��;_�+=wQ��r�rK��� �m乼ɯcr3���6��X�����~�O)�_��B�&�tv�s����瓊�f�VU4����lk
*PU��� ��㽹�^��)V��~�>����Y���%3zOc3�����{�w[��:�%������"fu�g��}�j��]����kiOf�=6����?1���fnn�!���s��47yo�̯L��7��z��u�.���5���1E�L��i����|�\��{v������x��c�+g�d~ٮC�]���}+N�� _.4:_1p����z��z���~�C��J�f�s����e[a��1�2�o.ne����vp��J���0�=�JC�f��uu������Q�s����f�<8�4Ec/ubq�{���Y]ǥٗEO��k��	�����9dv�#��8ۥ%�)T«�z{�y��]�Y2�r��/��4<��H��u�1�:ʙ�����˂���TK���}_W�Us���M9��a*a��	��%T2=6���:��}�zj�)b3'a�{���'Qq�E^1����x�(=�yR����蠨ql���H�1-c�#�I���w!P\J� ����C�^~�����/���b�q���EO�:���;��/r:(�@f����{�r�O��$�I������i��m��T��s��afE���ft
�\�ӣ͈A�Ԥ-��@riYw�烌�I�ӕ�}r��qj���OM��s�>�@閟���L��w����y��یe�L؎��9\ƹjq!�Vs��ՠ{pc_�&��������Uݭo5`�B�T�/k�����}�]�cX�~�nz����]���Mb�
l���5���n��2n��Ht4؍���C<��:�im�^��&d.YΙU��P��ml˝��S���m�kA�������������׌�l���B�;܌|�EN�w9�S^f���8����"�n���ݬ���K�����7��q^ E��3�'F���\��̹B��	��Ddr�'mY������Չ�~�$��j�Qw��k�{���O����
��;��o�3�����oX��1��]j�t��i>w�r�ck���X�G��Iv��{�M���'1��d�z��|�L�<[���\�U�qsj�u�Cc�1L'y.�Zwn.�ީs����O��|���svc�KGT�c�v�9C�cͶ�o�>ߩk�����^��jڽ�I��鼙v��|WM��C�!gSkaخ'�C�3TI��
T��]�]��o=z�.����݌a�zVpm=�9Xr�Vƈx�"��2�CD�͹�ʘ\�RY�I冋[�,�|r���c
W�tY�ќv��f7����o݁��:��-�w	wYV�q1�A���_qL�<�fZr�I���~�s�!>:�M��73��wA�α�7�A�[�H�'�C)U�;`N�f�`|����$�Q�4�i�ۭfT����b�@6��i�h��dtWc3�X���m_X��z��3OJ��Y�r���Y�/�(V�Lk�B��M����wpaX7��Wc�{+r�h�(a���W�W����Jv�.�D���3��ה�.��E�=3s�����1�ĎK1�ܺ�"�V�lVM�Ѭ�/A���9��\�+�����h	]�2���RU��-JM:b/���my���rL�-�v
�!1By�f�~�Uod�o����fW)�8Mm�?Jܜw�g,i)�XM�v
��b����]�@�X/��[㩾93׌�BVeKǷ�'.�o9�L(~k{x#�V?)Y���c���I�_#�DBa�vM�ųo(	Xr�s�YZ�&z�w�8�����V.��(�Y+����Nkπ�.ީ���]�_�]� !^�xx3+}�N:��T�'8s|���X����S�[Y��}bߡ<6���eZ@��i,5��X�����Ϳ7�K���rm9V�/6�P�}�.(�.'�E��%�d!7˛���X��W�kc����Q36�0r�y&�ީ���r�7zpȟ]��Υ{�%�WVt�ُ9up|��4�W�{A�v>�w�q�·&a֫�$�ǽat��PByL=��(�V���3h=��-݇�N,!N�WC����w�C{dV��#��B��/�����B߹��+7@��Lvԡ�v���N�%�:O��Zd��k]�e���]�A�6�	R#DΦ�	����*1'|��X�k	٘�	��!���{�Uo0w!ׂ�)�?����v��w���C�,(p+_�S�x�F)���͌�LއT����/r�� �$��`���+��Ή�m���İ��V��4�u�9��m����)*�˽�y�j�OU��^�U����`��a��Ұ>.ÌF�z)�9�2�
��S�M�N�^��f�؆z�hJY5�H��Is��o��8c]��',������E&�9א��؜��c`���0�&���^Œ3^+IT��fkɱ�c����*��hf�V��=,{��>~>�7��VϷ�^��)���:3h�7v;�� ؜�C��\��T��zA}6�.߳�nr��{����}4��c�l'�
N?�C���o�MnL4��C�7/���T#9t� �փQ�p������ٷ��s	Y#�s�X{cJ�oS�Y�@�|�{J�uq��^�O)�;z�0!2."�S��}m_�YO^垾�u���j�Y��̫�G��7F�1m�k	H��q�,
WT���SJIlccwhf�TҊ)ޡ�RfA�Ѯ���{�\�A�nW!Ȥ�`ʎ�7�!��Ez�}t`�˥�ޑ��+"����\��EѮ���6�y�R���MՉ-5��l̡\C���4���kkd����*;=�kV>��wy���Vs��YH�t }V���[����oM$�$	��[������IwR�k�wKZG��6��P�n��`��xw�nK����v��Iw2�B����}�ϔ}Ҝ�NP�(±��z�:i�y�����Z�s�ڣ�P�V�,�ǯ��ŷ]JB���j�X�<@�.��[��)�mJ�3V(Pկx`�j���z�뉍�5���k��Թ���&�*�:��w����u9So�WP���딴:�Y��[Fb�r�;oLF��vSD�_K��[o��j�.�bq�aQu7�.ܙ�ܷ�ݓ�o�����Ǟ���8�2b�΋��[�x�F�R����]��t��}���Zq�M����n�\�2�M˛�We�c�[���wn��t��k�n�m䘉�
�˽���˽�p��Z�W��`��b����C����\C�Č�Y�+����/PN�]�
��*߰�8h�k�:�)��K�e�-�2*�<���Φz��u�a<�.Js`��=[nL�NX��^!j�tU4%�ѕ��4��L=C����/�14,�2ڄ&5דn��<K�x瘕k�`嗨
r���	o�|-6�gN�wB�i��nz���Y\~̰�wj
)�W{ڨ�A�R̫�����1�X:l�=�ė_X�ONT{kwci�=H]4Uv)˾�oV�6r�8��oz}�e����W �˜��$��fk�\�\�����հ�-�R�����.��k�9P�k�M�|)�W@�����cO;�s��B�we!��L4�д��]uH)�x�c48�.���T�(á��Y��I�.bs��|��
�/��6���)��R���5MxA1�Mu��㷷0(��c��8Ww9��sh�L�)^�5��u�m��ިX��w��+]�۠	�W��;��^$�f�T��.��h��� 0�|�[�2�Rn݄���_q�l�ݙN�T؃������3�.��	sC�\�f���^�FG48>ǹ��ӡ�Y��8���1�쾮V8�p*��c;��.�ly�+�V�jH����u�EsUl���T1ʜ�ڧ�M�;s|�wX�Bm����VT��rl�KlX�����֐�e07YVCx�
���qg`I%�A�X�f�C7�����h��D�{�h (
�(|*�Ii$i2e� ���4�1zr21��JlJY1�"%h�$�LB3�F�sv)���(�Mƒ��	)baI��L���&7wae -,i1�W9��$H��ґ J")�4���0�B�����6#�!�� Ɉ�1&L@'-�l7wF���"#bƊ4���"FlR����ɨH�I�Y@�ˡ �1������&̘b��c$s�0�Bhwp�&��,�dRfd�F"L$ș˄�D"d�H���DSQ1�&Hň������A� �߯�ϯ�����߷�E��:�m�ɻ��N���*��ܼ��6h�G��+�V��$��:I�<w�V��=�
�$օ?����r�6�ʇ�n��Gg�cc���=c��̞�.�j�]�Sؑ�l0Lu��^iW)�&M��G������a'���^�{_f:���3�U���Ne�T��:7.vv=��|��K�/О���oX�9�/s�M�<��W[�����4�MZ����鴽S>C�Ξ�Bx�f�t���m�����Z��S��Z�1��T�ʀ�}YO��Ng$=�ge�)����6��}�^��ꅝ�Cά]����:(ʦ;�-�Cs��rՐk�}��X��5U{�.���i�����r�V��=�AiA��n�����,r&v���vEM�V֡�gW����r�GFE �7&3{M��U�Q�D�P`�l���qB�U��ot�g5�)����v
s��޵v�ߖ�4<S�6Vϯ�ri_��m����s��޻���Qi%on�b�Z�r��<����>�C�~��w��Lb�ml(��ڜcn,a��<�Ǝ�{�J[=dV�]w'JKf�yI.\���i��Voop�r�t�So+92_ ��дǚ��e��]:aEeN��=�xN���v���1��[%�x��}4%ne��>�
�.sM�.�WZ�ebޏJ�G��y�����]���x���V��}�X�}��`r�����dV4��ɹo�������(w��3�[9�����l��j��{��~��&����mU�u6�Q�6#Z��k']������am�#�r�ɰ[M����%b���������������yʥo`�-<�f�e���V�WU\]����+Z����39������qy�#��W�Ϝ��8��g1�{���{�v���Nc�79@O3��B/�5�t'���y�ga�R��>�>�^+���{e�T���!�Ppr8^ �L-�uJ�mv��y��X��X�=��G*����:��֑�=�J�i!7ޖ*r��!7��6�}r���Π��w��yUj�w��c7~ļ��y[Gr,��Z��Y��G�s�<q䇝(뙽�;Fd���s;.��;M��h���`;�Ou.����k�*����"GG�"W�\���8�)��ڙq�;��l��].l�0��i��i����}p�d�غ��]L����a�ww�v��L�W]-^�wx�YoJ��i�Wˁ܅^\J����1ݩ�9�7�wBa������޴Z����z�7�\DNo&o.�������c�� �'ťBc��sȡ	wX
-��c:�eL�ӝgz�ʅ�j�f�����뺶�za�xc|G{�g3�Q�ƅ�o���n3��2�<�ao�/����L��~G��\K;�҉/Wm��qu�Rne�(:�9�)�4:
�`j�5�7{ ���^<�a������3�]3�&]��5�V%1BD��l���ne,�>�t���7�w��Fs�a%S^X�lk
+=�X�`�|=��7�]�z�`�r�U���$<��ϖR:x��w��|������F�^�wXh�l�b��m��[6�9^�u��@闍U��� ��2���H*)��O���I���ݍrA��aX<���7�8�0]ۘ�����(i-N��mJw��Qz+y+�ܧI;�r���Gjs��J�Vu>��+NQ���j�\��)9�.�D׵���D��lc�e���ڦHW�^}c+�g:u�3����k���>�Ay?�SSjq�W�b�f�}�K��=�\t�g�.��,ng��/]�/�vV<X��i1�jp!V-�S�b9Y��vs�	���\k�s!6�%�m���cO&m��q��v��~�-�)����:�,����{%v2�ss���ϬBΦ���G����<����݋3U��r%�K�dwVC��݇����>�⫭�.�><�Ɍ֣P�'���\�L%S��R��$��k��YEe�]lZA��T�շ۳�
��O�D�d�NR�<.n孷YZ�E��UQ77�Z�~�3�[g)�$���Dm��w�M179�9�ܛv�\�0l���1	�~.�ny��^��ӪrT���At��T���(b!J��Z��]7�
�&����vb4zK�
e�_��D:�Ջ&C��ٻjα@��H�՜2.Af�����>�]	�@����[�jI�fk4�x��Δ��;i<���l"H�;X�۶i�_jeK絵|3�`z���N����O�sqN���h1u�5o���]t�����,����8���*ۙ��&���gt*	s�m�v1��V
�č�P����Պt��Û١�_Qƾ>�Mw�?��^z�Ww5׾5_S\�6,�.��e�bФS	��M�/����Hr�5���3}�#���{���E;���"nn��hМ�kT�V�mZ]��9Z���K��wAjQg�J^�9Οv�M���<�j�c��-�]�]��I�Ȏ{4y2/<����ʒ���9X�]-}��|�\���(c����7�|���L�x��Y��zߦ�ŵ��n1|��K�.�����=�V�l�c�4�����>��fҵ���Ⱦ5��p}X�NB���.RZ�LE\���ة[�*�Wo����c�����L>�J����-Q�r.,+��]������ ��~i.�KO�v.�\+���|��fzw���Q�P�z��2K��N����]�ښ̀7��l�Iq�h�]�N�-G�UF��kJW�.<���i$�Ѯ�t������ln[�*��]p+�!��滥��<7�����ά�υ���nb9Є����������Ny`ѭu��ꯖ3y	czb������A����6��,n�܄���7��br�1\�A0
۷�Rꢮ��f��dW�'�ƻ5������r�W���w�*�ם	����$n+ǲkS��u�����4-�g����9o3h��L�&ws^�d�~�f�uk�+f�aW&���[�����v���r��ߪ��W�oc E2�M�鏯�3s�F��Tc���	"11�vx;�B������|�3Jo�����#�����gt�uoS��b����m��&f�lk
�k'��&z;g>vc�f�at�ؤ�:���k�}�V�Tׅ�Pm����k�K��]�2e�x�>��O����E�B�۷��{c^MeZ�oK�)�r��,{�j)|���g��[�{�����lOc9�So�^�O.uo�eiI�Z�kë̠��%yd����y�+�}����9[�́�s�;Yw�l���θ�>����Їl^�݁Ҽb��k���aT��|Y�m��t9($���^�gq�h4"�5��fd���NfD��b
N#"����,�����/g�V��:3%q�=�nl$��8LW��'/ϴ�؅rsznr��=X�_>v��$!|�}�E�l<�{���L�>�^+��۽�Ua���W�]Rfd�Hc�,}x��sqYC��!��^kz����X�=�!\�ƪ�}0�^i�^y��>��"9�ެ�/�ny����녝M��b���E�&Y�iW��
!��hg���SԢ��W;�+a�����OlB���
��5�J�@����^.><H*�|0A��&9И�v)Y=ʹ_c�0���9���<��ER�I��6y����HP�S�y�o�.��}��F��O��2u�kplPT�7A�9����};:����K�c}�l/d�~N<w����vU�����H=������$y̾�t�\���~R�n��$Bٙ��Tܦl��*o����v^"�����vg�~��P���@�_��<e��?�7�;z�m|�݃�#9?)����]���VmZΘ^H��V��,��S�d�ۭ���F��f�1"�t���
�q-��-ј�V
�.�@��wl��Xs
����M�����{*T7�&O]�e�<�y��]�=Z�}_RMKu���uד�̚��zꔓ-ƻ*�bG:s�8�eL�����&�������&�1d�9㰒���)��쩷��:ɾ.�'e�;��[$Hz�������Ȏ>S��>GO9�qw��Ϻ�Չ&��3_M�Y�T�{�?��~�s,�m��X|�+&z}�_N���z2��=;��Mǟ���>~�N��>��r9�����]��~z�&��1^��� {��P_bu���70=�aL�
6�n��`c̝oau��(l����Y\��8��"�q���_�6�^o����<�MɳO�B����Sn�rՕ{�vv]�/�!	˛��6�ľ}p����=�S�R�0o&1���>��c��(r�dwP�uB�sv���H����Ố�A��*��\'พ� �
Y0�X�*(I�Ւ%��}T$���q�-l��)&�;�GdE�7����g#6�Ш+-2U�v�k�9�y��v��ǐEB����P�J��Ͱ��5wV!Hj����%ث��k'TϓۻV��a����1#��i9�7��dď,q��N�Xw;�?��w�ɟq�b��９�Z��|w!W��Lh�{���OHøZ��;�%�����M���4���]�^��N�+�:^�F�]^�,���-'#�;����������V]���z�:�\�)*�yu���1�`$�K��b6!��������\�K�����#I���Ylt��X�Je�]V�dE�x�+TЕ�419��T�-�-k�uXz�x�"UJS1��c�>��)L��xfl�j��i���W֯=}+��
*�5Wr0dm!�Y�9B��̾|5�*oX�Μ�5��kn���w��@��4�����uB�7U��]��[@�y9���u^|L��Z]��Jo��Q��[͖���i�O˺�k�z^߱1��9��[����Kj����_-]'`���2z�`��"��yZ�]G|�������<��3��;AO�6���=�\j�ί�������V)�m������vuݤѤQo.|�\5빻œM\ ��XNf���o(ә��F�Sx#We��Û�uf������7d7�򝂺�zhD�o9���^��0gS�W-��9��l�/)���z�������R{!�ȳqy��s��	�����!ˍ�����v7��B'6p�OD1]�'��<�LS�eا������=BP}X�aB���csd�P��L��;[�*�N`�7�g�f�϶�{�C[.��V�Y�;P�k+R+�w�:�=��\���YA�����m�4����]�����#DP���Ԣa.zvg�9�t���K���ư�=/凭&w!P\J:(�n�֤�Ӹ��3%���1ܮ�ȨI�V֭c:����t��asO-ҋ�4�˷��U��#���0�+[��u�o���޶εy<��c�2������1r�SC���6Kڵ�Y޾�\�H���dɺ�yu:��H*5Ŵ�8�*"t��F�)�Е��No�-�UL���v�V5	��dܱ�Yv�e�+�Lқs]u���>�~w��R�}y�p�ۺ�E�H���$�a�dy�N��!��;��:�Qܵ���bwC��]�)d����pKN�;C0������zr�sU�9���i8�q���5��i�u����]�Ԛ�!�.�N̲"��+%";�@{��j�ޅ�q���&��p�o)�w�����[Y����-��g-�a���0բ�*�!�*!X����aJ���8ȱ����N�]�h?�c c��B�V�>窶C��A�5ՙ��uY�i*�̒W^�#gn�v�*"��`��<o{"����sڑ(��8��J�r�*�k�$�� �/��Y�ٌc���*}n�]vc�yDK����m<䋖�*��g8��ԑ����zk:@��E�5�"�Ә�yp7�+h�3�ᖮ�LM�]�[8Vu^�LǓp��StP�̘�=�'n˱��y��!��I�3�&e�GIݙ��eY�\��h�Y����ƞ�΋U���. ������D�	�ӝ]�^}�M��Jad�D	�<s\;iV3���h���9+�;=���ї��Z�M�0��Z�ϩ9l	�\���xm��֌�`���T�C6�@gB�@�]a����]̫��eD&9�ܺ����4�&k�w5N�{����ԎgZ;�8�Ѕ^�����'u8 y����=���E-C�_,a�+�.����h���5Ƴ���֋XoAƜ��Ri.����5�)�MV=����7��!^[�6�v�|+�Q��ӻ�P�.Z�׀�u����jZ\1��)��d��jǺ
�h�e6���զq���1�l�r��8��6rI��Z��s:�X�ˑT�r���4�\FoU�{,%m���xB���O�L�;�� x��&�m��h�T�qn���2i�����ttC2���]�Y��m!�a/M\Vkf��;�V:Ă�I�Wo1�	�d���l5g^�n��B�%��k���0�ϲH.j Ϋ<���YI�.S�� &�Et�.��$}��i�ܳ��!}-�.��q�=�-���*Ƶ�����;�G}&�wu�K,5x�����i�k�<�ұ��z�gp]b�t:ט�vs�0��SfR��b`�s��j��m����\�nQ3N�8K�v��Z�B�00(��%wa�b�ܥ�|�=�N>{���ej!��=���B�|�Aa
�W�{z7�;Q.$��jr9��`V�֞���r��;��j��v������10�'�Mg��-��]�ػ)��#C"VN9��/7���X���T�+ZE�b�u�]�܄��F*�VEjH�b�'b�;E�������>PR� �@Me�a�k(����)#���|��+i)���c6�%�08k3�������D���{D)��C�VG�����*��TY���a�fM��@��p��׸���X�ut�ʎ�c5֚n��7��
n�����o=��wg'����K�f�ծ�K/V���.�orT{�W����6�,�s���P���I1B�]��iA$�aDH�C3�d�����AI��̚"c2w]�3r�A&,�f1�D�&���u�%��7u�"De&�X4$��&BIf$#LFDQ	]�5��"��%"�	����L�@�!���RR�2�0i!# �ȍ)eA(��fP
4$r�$�CL��I2L���d��&%�2&9rK
h��ɚ"DU�Dca(&3��"����B ����E�D�	"���f1J�]��I�%$�$b���&�$$s��W{&���v��4��Mr��.�����Y��Wa�"�G8�U��}�4�cY����h����M@�1;{���k����ۍ��9&e�1�A�P�����|6�L9�YQ���zUʝ���e/g5���2{sh���6��NW���1���sՃ�2��<{މߺ{�nD���g%���i�G7���iw��|�����e�"��8z8�/IW�#	.�z��b�)�R��qbޙZl�7g�M�骑�r]��֋�F���y���ܭ'T<r��Ërz����|��C{1��m���91tv�s�RelU�p��-�^�K�c��&	Ϭ9������#6;�b��V�Ɓ���xv-��	��%�m��Pƶz�V{��0��G��''�|�]�d=�U��ߔ!|�s�m��K��!gPml9�{��(N跽��ё�VN����`t�[����a������������T�_KZw��3���ƈ+�	��c�إfc�������!��&+��LN��⪙9�^ 	9]�ٻQQ���Y)2(�Y۹,��|��r�[k%z��M�R����7ۯ;�� ���D���jOc<�⃍;���5[��>��akb���ՈE�YP9ظoe$�Ȫ,�Nm�u'��Mۧ�M;��9CQ�5ݣh��}S���
����1�K�,c��sȨK�c�<�i�U�-o�."ֶ�u,q��T�8���L_wϽ1�_>��ֲ�H(��9��b櫭�7eޥ�3&����yL�z�k��Ԯ�5CI��~�6����V�GUc;�}��sH8|]����v'��O�K���_��_7c�5�{�p~Rz�vd�W6�gt*	uM�.�lk��O�9��e�:�/�j�Br"卂�l��{�o&�,���ߒU+R��'m[؇��z�����g��bƺ1�k�-�Y�/'O�R:x�홍�ͻ��wZ�JNa���98�jv����>'��+K��UY��Ҟ��#��[~�[������[�̬�������|��=P��^H��56m˜��H̼٘����L4��kz�L�
6�n����Ǚ;a�;��|⒁LMh��V�^�idߖ_l�[�����A>��
��nŋY��<��,�G�{����{\/��O:��Ѭ��0P�Y�U�!P�ǶK�y��𭝽$]�7]�Ԩ��-#peg3b��8�Z�l�턕����b,w����WQeM����c%��Ԡ���\k��	��%�m��o�ky�K��M�k�;�o��:	��.Lc�S����_aC���=M��>�k�g�6o�����I�v{�S�5zI�U0���ʽ��Y��Û����u��}7@�p,y��I6�u)���_��%����ʀ�J���t�E���]��S�X�j��ʽm��ޕ�-�ۇm��Z��Do���*+6/e�������@��ӧ��,%�vxk���PuI_��t�LQ���ق�>R�f�K/f�k��`�ո{����S�S0���4�Z.(�[=���̊������]}���J���vb4oGkxУ׹#躜N�Q6TFN��F�Z�%nN'��
��5��!����F�f:��j�(R`�|�#@)�4:���+rsҞMb��k������9m]_g�U�Kef���[�݋YM���I|z�u�2��z���	]vd�!� E��pky�������~ު�U����?k��v:�푎�n�o�_Fk�>i��Nقo���b�
���Ǘ#R�Y�no����ٜ,�Ϸ+yYv����f[c7�P�9۔%����OfB�:'�H}"8�r�w1������V�\�ؘqB�i9�X�����]@�x���:gmoM\���;��H�k�Kl[��5�n���&5��\���v�w�v���R���r+o��w�[3~�1�dG1OU��Zm'�ƹ{�5�j����?6c�{�XW���a�CƔ�Ëj��sWQ�.?U�(�Q˝�g�u�wJ�ߚ-w�~���L�90NXp~}R���:}������:sɹUQ]��1�+ܧR�<��]��~��pznuN��^�;��z��Ɵ����/YNoͷ�->�Bά]��W�Eʐ��G��׷|�9��vh�`
OV�����#Z�Y~K�m=�X���B���o'r��@�J�[0���f��L>R��I�k��3�[���q�c,9 ��fbl�ygR���(n�O�[Po���J�w� ���hE�)�B��=,���t"]F��ٙ]	�V{��t3\��u*Çy�+� d�~b:���W��%?��I}�t��d�ıŵ���G$V�l���g�����v��BAϷ�Ί�o8��Z�P���o��3��=�����ԁ6���]45L%潁 �ծl���C�K����A^.,E��F춞��f�7�A}Ӯ�Ü�7�RّN� �^N<�8˭��]E0�9��a�3�T:�w�����i�cT{<�N���5����˒���i9���'�N�'w��lk
��#�;s��L�}��*3q���%x}T9�j�śT�b�zOL�c���;^jsX�wz#�k�+�HW�q�[���Y��ZOr%���~|���ϡ�ba�<�;�T����۱��o����w�v���mux�*�}BV���έ���2��-ZBr�:O�oP�Y�>���淼V#�v�9V������F�)*7z7I*vT=p�����y�۽�կ\�ZwMU���8����S����r��\��>�33z�K�T�57+7FC��2�9Ի7V��#��$��:\�El6nd���z���O@��k�'�ڜ�[*ѝ�hk�ywH}]/�3��K�%t���%�1�e[΀�a�tQ;�Edc�nT�ӭ���k��-�(��fv�{�#��HG?>9o.`���%�m������=�G�U�5b% �2���ߑ�׫�C%u����[����}p��6�O��Qb��ْ�����sUۼUr?za�	���JZ[��0�[Ҷ�i�N_�c�2*�����J����nzK.cD�T�U1��
Vf;���kWG
�G.{e�d�r�,5�):n��Kܤ�/4�Lr��sȏT�i(u�N��)�f�8d��J��ǂ�Ɋ�vT��2p���V���^�om[s�If7�x��eޥ��a�g\˜L¡�v��D�F;{7σ������>��J_e��@��U�\�/���Tt�D9=��:�y
2(���ŗ|�x#s7��'�;�PK�h$�v[ /�V'��T>S��m2WIn�k�`��v���2ħ�^Œs�a%SAc
Frf��=j���v֭�Y�i+8�!�\�]�1�y}�cEF��zoTI�1Ḻ��'3Pt@EJ+���=���=uhݮ��ݢ���[��@��cm��k��0���4ب�(�g�鬄���3����n-LH���(��]3]��JZ��.n���>�f8J�t�K̡���ϒ9�gr��D8?�;ӄ����S��h��P|O|.�ͼ�Xqu��{5'|��H��α�s+cZ~������k��!�j�{Or���H��s��գI^����*���	�>��m������<�����0٬e����g��6��b���J���ƺ_1bo��]���M�Edqq����z��З�ɜ~�8���P�P]��r�|���So�:��j��Y�㣹d4km8y�Kc�W��]>9A}�P�_Y�VyIR}�H��z�{k�Z&���I.r���|��-\OH���ba*���Go!��'^9��*j�ԞX�[`=+j�-�ۿ�T��}�����=�7��9�{oN�g����7��q�45��/]RV�kܯ��n���n�Y:�،n�v��6_#��*w[��Tۡ��n�-A���G��,�Ƶ��u{�5�6%J�C����:�;��yv �>9[�IAu�x�}���6�/lmlý��E,37��&UK�E��iv�M\�u�B��`88gv�}��+�&d������YWm���o���Hz�{��9����I^k�9l��wn�� ���]1}�,j�]7��I�f�q�f"�.����,j���&ԇ�Jk�2��}���
�4%nM{��A.r��.��x�2�hV7�e����4k�V		�*)�V��uC=��z)ҽ`*IcO��oen.���T�5S^y��&ƻ*n��aV�yt��<�m�Y{So��B����2���S��5e^��]�/x��O��:��l�F�y�L4TT.sِ��{�ʵcz^�cZ{.z�9�n�.,oW&����������ZSp����
���Zm'�ƹ{��\���X���Gp�8LS�y9~ױ�p�Nr�M�P��W�������0\�OC���Q~�a�8���6���;�s ����{:}li�Ap�O*�H]t�ǚ&ԣ������
b�[�)�����Cb�Ƒi�z+��.WE��1�8����q�b���8v�D@s��R���ζ��\��X�����W����n�+%�u�u.���JQW*Wӣ�B��W^,{���VPa>��im�y�֪ƶz�\OL.�cU0�_��t��։�l����oP�B�崵�i��ά]������6�_/>�-�Fg�C��L��FkK��)QK[�Xk-�{^m=���c���n�=2�N�D�:
��P� �:��wId��ƻ��o��"C�Ņ3�f�t�1rc7��}�s �������B]�U�ژ
�Q�^ӕʽT����Bpwo/�.��'��RF�HO��sel�텮�c{���	�J.�_:Ȝ�L��y���z(9�5�ك���鏯�3s�X�̺[W���y'�&� oe��Po��o���v
�)�4��׺
� �}H>�H��
ͣ��&��\�ɠ1���:���$�כc]��k,s�:#u����\�/�Q�=x6�ofX��hb�ΫW��hz�
)��Nȓ���S�����ES��Kv��lW��c�Y����/V�}x�[��2�$��a���B�e���ewZ�R�NT�l^ν7�vuhwYh�=���䗦�q�|�hϥ�S��D�]rt�K�rڠ�!��Yr����7䋘1��;s{fu�uv!J��e-��s����i�ϑ����4��ឫt0�Kp����Ѻ�9��N�n����A���{^ş�M`0~c߆��}g�m�~K��׬�蚗vK�i��q�&'o�<�
�k���,\˲��éZ^5�'N�=ŻQ��n���΁R��Z�|�o.95�[��{ܼͳV��7�||����87C��'{�h���*�j�τ��~<��ꁚֳby�g|��{-��1��KNѲw`q�i�cU����>:�ӱN ��Jgp��r=(=��E�L&峒�c���c]aؤW��W��o����|I�f�gS��3%�쮤8u����q�����#��}>�躚�>�Vc����h�EĿ,a�,�q�O#1�& �Q��3�iL��n���M�c�MGA�}��Y��m�7_j#��x��� ޕ��;�@s�j�=��׼�VLM߻��x���ɹS���6n:f��<ȳ�ڑo�J���i	f���<��'�ܠ_�=5�s�77���Z��mx	�OxTz39�9%z�Mް���F���7�l�*F��ᬺ�#�bD���ժr�X��o���ȗ8k};T��l#�ԟF�sc.��)U���	y��t�C��z�N���O���S:��w�&��9�xc.�xp�nޛ�K���tN���Ƕ��hI|;Nˠz7@�Ǔ���u���z+�K8uh,�vŹ|�_�d�5R��^�Ů�*U9�\������E��nc�g>�Wu�
	�e6֖�6h]Mc����)>�W�2u��YB���O�6��Z�)os�Z��n��zL�
��8 ��,]�P ]/m�Ѥ���%^��}62V �%�i0onvMEb:��Û��Gy��Ԩo��O;2V�e8E�E�Wl4��	��)ub�×����miRԭf��v���s���>���<�_pvn�+e<�V5KQ�.��R?&3�K�Z�8�e�g.���˶��0`�f��2v��;R����/O![��{�ȫ���dR��^�g+&Zs�Z��bK�,W!�]��(N��Wm>_,��z�k�=+΍1Y�j�0��;K�T��T��:�hL����7�G]+nͪ��&���e�|{xg
6ax"���Pϯ7}��I�ܭ��Ը�0�gv�)`�fXv�{����D^e��)%�PL@���9��7�d��|�Y���\x�\�HX��;�p�us{B�2��#�d�/Cu̕��r�u"	���]\��`�\bE$��w�8�Д)��M�qB��s����:i���֕e�L޳��m�C�fs�C�|ރa:n��c�S6��:�
�j)F��.�� 4�����S(�>�#E[���l�a(M��ۀ���������6[����ZԨhʼ���͠Ł%������❠�
ή���t�
�%�*N�YHo�.wq9j'OAf8.rv5i��pwN��!O��ƍ4[�4�[X�k{���t ����2�Kv:�k^P� 5�h%u�5�#�JŅ:��N����ŐL[JzP�)A��J��>����U�-C��5�Q�m^RW�j�M��S=��܁�u V̏�	�X��e�Y7#�N�CY��:��J_��
^i{�{J�I��ܜ�b�7^���6��iWn��|�O�ZY����smLR�B�!6Fl�$ 쩽y`*� �\⏨����5�qNSӾt/,+Hۚ,�
$<HT��u�e�YB�o���������X]0c!K�4�����e<G�$��	.^�b��ܼͨC�x�d���YU*���2kX�
}Y!:���જ'�Ӄ����bUuzX���[B�|���Rs˹�z]�*q�DR�e�f���z˭ĕ��\�wݕݪ<��R7&�A�fmڬX�{iQ��Ș�ZOZ�B�����+((�]�Ƥѫ��w��آ6���ݳ�;'�DP��
NbY>��	'ȁ1L��		�[�1L�o�5�j@�b�A!4��&�Ay�DO;�03 B1��L� �n�3"x�C7H�˘،A�)L�RL�2m2)�##1L$�d�2d(�F<��7��/;nF4��2��B�)EA�F��DeݷIDQA��;�-	��ݍ��RF�d���4gu⼁��ٷ��2�*D�%d�!� ot��I#2�"��0lP��&��Q9ѻ���;���۔�S#��X���u2��)��D����.�H���2h�GwT�@)ݸJd�Liy�*������^5�j=�2�\�~;�Ï���ۉQh�w�g�MV$q<�b����96�F�*�	�itzVV>�J|�d�Mө˫�Ŋ���~�5tX滌ty]��g�&���9P꩔L�>�RGjQ����qk}��/8S_��ܡP�{��coqH��Lh�؏\����\ΝBZ\L{cHU<; 	���N���${(J9عG�Ҫ#���nԎݵHTwrd�e��s'DY�(fD��#��S�b��$����u��}d��G)B��^�y�*��^��c��"�_:�b�dc˂��������U��0�M�@�Ց2�ŗ�~��~;�[�y��(<�K��%<���_��N<�o�����v�B�t�V�.f�� �PnX���i�.��w�zZ�S=���Np�&ˆwJ�VTm��b���m�L-��~�	��e3����D����{�y�m+�A�����58�
������.5-�|�c6ܦw}k|b���Xw{�y�=�T�^w��s� _��`u��;��
ɭ��9'�ci�7�Z�����ۜ�MX����}��S2GT�%��3bd�5�Rf��d�јvT�I���t��^H1��� �-�#������|��0'�f���6�2yS>?VN��q
�p*v�6%�f�b��B���E7΁�/q.��jh�� �]o���ru�/i�Mu����/��wk�[��T��0nLO;���/m0�&�/���C&>	;����VZ[�^�	�]��T���$�#�ٝQԌ�2:���΍�?R�2���ܚ����ћO�!�w*ٸuɍ��nOgN�N��Cَϔ�tĹ"�س}U�=S���XS�/��Zg�ӳ�=��axOm���-[.�>ƺ�� ���2�����7Q�y��e�,g�*!L�sWr����]�s_�D����`~R�D�3�3�����F㥽�m	����D����jν����p�.�g�Y��j������ۯO��X��<ʼ�ђ|+��jz/��Ђx؄�M0�>x��ܩ3����ܵ���TqFg�b[�[�=жhq/��`�u��j}d��PH�;%�#�|��(�W�J���z�V]iW�[�r���,�6s�`�ܕ�1����&���<ϑ����wg�YM�J�S�\6�Q���F��:�F����$.��d/��t٩chd�q�
��u�W���G�L��4.��Ӿ*#�WQ׺�ǹĹ=��t��1�f�=�N�z��ur�!��8��w{"׍e@ٷ:��u+�I�kp��ߟWN����h�s_�<���9
^MT=}~��p�U�F����C"�YҦeu�y5.h_N���/�CB�[��$r;���3/�u��B	Y�-uq2�S��֤������3�x?Jk�pJ~XNL\?Ln���n.=�r��+6<�E��3`x��J�}�*˞/������V��t�Typ��ᚗV�/�.��]��f���:+ry���yTq9ٍ߄H�"��T���b��
�6�&F&�n�.ql9v|%ݽ)țO|A����q�k���Z7���T,�[0�d�d�&���������gT�{�����|y ��kxͮQ�r�:�e��/�G�,GB�Iܙ�L����)num߷oV��;��2��a��鯼e��s����7-���ꇶy{O����� �d��q����$���y����Et���إ:�L�ޜ��:j;��x��x�9_7�/���üu�4zt/O�9Yv��?lK�/�ĝPg �{I
Oq�tk�o4ɰ%��O�'��I��* �A{���:�t^^�DS�(�/(�|�� o(3~=�ru��c�Ucu_Ovދ9���ce�
�0k�Qw�sX0��h��uU�s��9� �@h�(d�Y�!�s���*;�0/f�f��c�n�(v�Eh��f�nͩ��1[Fa[3�cvN�8>�t�Mdh)��ݢ�y�!:������v�ƞ\��Y�8]�%��=O�b20y�*&襛�U� !�]�ss�$��b��j�k��SӖ/@QK�i����ś`��z)��l�sx[,��<���L���<=�Ol��H�Bʄϵ���=�o=�x�){f��{�£���Cr��nϙ.�/ ��d�����}�$v���\���et���h�vs�
Y;�]�{���U&+{�k����Qp��D�ӓ&��G�n�M��E��1�(��c��x_��Uc��I����-����2�̭�Ȟ�/э��%Ƣ�Ũ��*� ��`WջP�>��gN�]3��=!��|mh3.|X�@����fɻ��w*�n5�����|�|�MA��u|�=2;����2�nޘQЕIG�}=U�E{�x�~3;�\sLk7�bw��c>�k�����p��˲<|:jf��d��(�R94/*�o��� ���l�	����+Y�5�m�Q��l���)�q�����f�Ā5������x�ϣ:(���8)t��_x���ꀾ�u����M��Н�{^���KMwzN>�b�w�B��7��Z|tI/O�]#�ץ��� +��W6�;i�s�8��y#<d�uY��5�r������޿{O�a�+8y�W�	#vkO8�Yf���u��u��j�*8g%:�ޫ�ea�Q��Ү�vU�q�
ށ�Y��rۼ�����U�����`&�7؅(N%�7�������[)���A�t�>�K�SD���f��Ó�%ό>�ʝ7t���1�T�¡L����C�\an�_�K��u������S+�6=C�����r��u��j_�(�f~��u�LB+��mm�G¥���E��ٛ\\�ۣ~P�侜��@v{$^s�a�a���HzW�p	�ܠ ���h	���,\�7=$�Gl
yEQqO=Q5��M�L�;���x�C�jW�dK=�F�$��F76!f�˄ϓ��Ύ���p_��paQ��u�:�1e�Wq������S��P��H���ǻ��bkn���]�<Gy��6Ay҅Bs������#�{i���o���OC���+�`�v_�e�{k^��8N���L��DVv&�B=��Q�G�jG
�ڤ;�Y-�����˖s�{�{P�)�Ѫ(�*�-릍}d��b�=�vr�|��(�k���/0����л�R|5g�F͙��E�hU��҅�c��
5�3;@��#Ƈ{�׼j����<����Q*��U����/�[꺏_k��{�ɨ~��g5#٭��z�:E�6,�뽦�K��ާ^{�וj�s�FD2oo�����-k"ʩX�[V<Yu��F�+��5�L�7��5�CQ^k^��+r��~�"�Rt*�H���h6�����Zm#Ri����;(�kb�����^�;�HZ�".� ����[m����9�v�K��U��(>o2J�����v���R&����w��9�����Y��*�R��_���oam���aC�4�g�$���{��/M�hS�c=��ӡLd���NTi�]*#ll�g՟vpT���ߣb����o�����ޯbr땝����0��W�f7~!� gT39���$��.oz�_jz��&��8��V�I�b39��uYs�¢<�)i��d�ј� ��Zii� v�mx� �;}U!���v?f�H�O��N�p햴1�=���yHݩ�N�;M��P��5���ټ:b��Z�zz�7�ۡ�*�i��<�of�rco��c'�z�tuL����Ņ1x�߲��%:����S�V��g=�_�n�g���<rި�ij�v2|'�GAz:�R3)E]+��L��9��`��LT)���w/	��{�G�u��z1���~u�uU�9%L�u��Xbf\�NS�u�%��@�Pd��[ (9:�U�_^����}\,��g�}�wDr	���M���ݓ��	�pQ{U�
���Q�@z���N�!}'�_X��_^���_o>��\/��~��"m�WO�C/k�E���{�D��tE�k�U��ovj��A5��Rۢ�빎Vk��F3�m^���B�SzL�ѹQKx���T��S���iۘX�|�v���Lc��9�`� _b��p��[�v�*��K67�����2��%5�81�%N�Σ��ް���5�W�S�U�rI��I� =��_#�|�1���>�Oxo��N�E�6��<��-������:�G%mLW�2^�}&���^	� "g���\�^Y��Jwe#��o*c_ۻT���%�m�����hY�]8jX�������ɏ�E[}��������Â=���ؽ⽵uq��L\{�'&��<W��TcB��:v,�;v/9��B�&ة��>�l���������S$��{��\_���m�V��>��@�.f])u%E�쎌��o��6n�'ޣ0�	��;��E��鍽�I�����T�G�7��SL4��(�j�p���{�¾��J�,G2�*�e��])�xe3ᮭpܟ��EdO+\�K�٣^Z�p֭��=�;�~X6��h�����<=�7e�_&���G��PҌ]�O���4]llO(��~<�Y�����;�Z�Q쿟e���:.�I:���F�6�1~�c%u�	=����S7��s��gkǔ�G�Ga�l�P�`����t���o)^׼3$�Ty{Q~[ܭ��Z*=gV�V')��B�m4V�����No5ˁ� m����z�9��nө�v\��tON4le���]��w�&�����[����_N�Ov���uw&ī���T-:�<�\]sf���N�I�_����K��𯔵��){Ҹ����lx^8k���,�C}P�(+�׵t��r�}9�r��8�<j4�%��� �s�iL��u�~*"{�x[�'�_6��H��|yO��&�85����|k�:�a�G�n)�H�dn��+�C��/���aJ�9I@7vO+vj��6Q���㶞����&��m���.s2�#� � �_����lf;=0h��{bmk��/{����u�l��-�9��5��Q*et���Od��x^������q,V��k�S�t�p��A���F�n^�͹�2]���sT��4TVnD��Qp�Ҷ��ܩ���5PS��P�v����W��[�U&*7��E��y�����Q����^Í�"��޳>ث�Ga����`�~_����3����]R|���c��P�#y��n��ZEK�6��s�P3�;�1��1�	�x�#�/2xX�]]p�B��fi�F�~��-׳GM�we�hq�~T9d�7(eF���od�x��������Ȅ{	�{-�徼�� ��#J�[%�'ol�*����l��3��.�P�\�;�QH��E�L���n9�v��e�)��q~���#�g����E�Rs��9�k=���"�����vP�v���.�Z`RW[�R聉�xr�4V��J�Z����9i�&��z���߽^�-��	��ƳcI�ۈ�����>�|�9L�+������n&���Uu��w	�^.�j���k \G&���ݨ̿�y�}/�p\ob8s�y��O�c�D�O�_�g�ҝG¾]#�kŁ�<z�f���<�q��Q~�^��8���j�����6nyx�6O�����,T)���t�;_zP{�� ��L+m6u^8[��ƀ���V�aXt2�M�Çݕ,�Q�N�3H;<.�餥���Gw���B>Mw^�b����@5���W{@ܨ�\���ׇ��:I�c Qz����P�tk=	�6�AS�R��{;Y{J��{Waz侜�����ޢ=\��td��$��� �@��6H��޾��\�r���#>;��+_�$�-ӱ�6���9;_?:��t���i	f���=�<Bt{7�&�K�:���mm^��Y�E����/�n�:ۍ��>�5���uT�]�74��F���{��)ċ,�z��e|$�_l�P�q�X,j�ܩ����#�q�'wti�WOpVt����;����H�n]�2�o��Ȏ��ˎ\��۠��1�o@�5��6�}�7�Kk�����|n�![�ܑ���}y?<�e��-vn*����,�xs
������ԯlDKj�@/���x4��Q\�q�U;yq�^��+.��rJ�d��ϫ*�}=]P��R�$��P��3�4j!�J�g�ԮK6ڻ��7� ������bP���:�9�1��}�*�(�tѯ�ɏ�X���w"K�2��{�J��n�j�}^��_:4��8�ʑ���_s�dV8�cZ�3��G�c�5��y^T�Y>��l���YV_�w�z����V��s@9/�x/g:C*5�s4�H:pܱ�����J�$�Q�֯R��|k��U�ʎ��J~1}��p�&�ʆ?�L�oX5>�'�A��uf��-�s�3�c���M��I�'��U���q��������3��t���>���6Ͽn����l����{ԙ���}���~�gT3b�kb\��N'H�Ы����;��Υ&S�ń=�E��	��q���쥥
'w"�Y&:����P�@��cPݩ�z�U����}��ei�����^��{p�hcOZџ7�R6�t��I�*ꎤe�ht��8ft�� �t	wȸs86�Ǖ
����������|T;�X�Ɇ���T��;"��L�~�+�?�(�cg��ӂ����޼)��$uͫѣ��}%ꫮ�1
����t�mC���M����,P�]��(��z��n^~a2/����y0z4/�N��&�,�N�8�}�+�/�DW3��_h��.��,m�c$c���
U����A�ʲ��Mİn�Y�{�(K��:�g�:w! k�uh��ݗ#&E�&^V��u9����\5�8Am �õ(����L����1�-@�������k�l��"��Pd�0�ۇ[Ԕ��&�]�\�P�f���ۧ�-��W�r�P������t�� �4���(jƫ:ƞ����t���4�˯ED�u�]9.�����]�A�4������>�΀��:������Y�z���Q���W7e�l��z�
3;��p���M�}�^7�m�l]Y�u����I�j�I�z�
�_v��n����ya@�k�7M6 k���ZZ'M��Օ�j��ɽ]��u�)_R�V�+U�d����Rw�f���z�Ll�Tv3NQ/��Qu�r�J>��Ý��#�NgF���Y*�g������W�J�(+���7�év:i�sx�'7_
zgn��������˅��V�#�";���c�c�s����(f5����6S�ػ�Z �:��Ȧs/(��Mo�-5gd{�h���0.}�9_1����|^vgRGV*�Q��`'gUa1-�d�;�Rײ�c��5Ty��k��ч��eC}�U����]Ӧ ��O��W�wOJ,�}}GCz@�&uq�Xؑ��j�r�-��n�6�K�U&v)�7�맽jXo�;�
V77�ķ���w���J�led�:��rz�Y���]i����ߓ��Wd��X��rۥ��:�ci�XCS[��_@��U3]��M�S��Y�+"[��u�1�@(�wwmnY�-�8%GYW�u��T]n�V��2�5=���������!`��
�(�s��7@�Vuwxm�{�A�K��nU��4����Da%
���*UԼE�ӹ}�I�����YM)Z��'�쬦��ެ�i;2��[2K�O@֍}ٯ���R5��ڍ�]Y��Qpy��ax.s'h'@e:����ˎܨ�oF�9��M_��/y-�0�����at�<�x*�������WS��ϸ�6W	y�YpLr+��� WA�L(gVy|�#נ^_!���z��[7�W5շ�}�b��W7Y!D��V���7\6�4��׻�A�]��k{�'�JWf�G��u2���L��J�k~�|U�����z-��n���T�jĥwvu�5�������9u���� �=	K.4��#ӣnG��aNZ�Ĵ��*��[�S��'�k�ړ���Y�Tu]t���i;��[N+6�)N6U�k%'�lևV����wt��]�m؝������Gׇ`X�>��;)P��C �W�0G72KιA�4`�R��Y*y�6��Ơ�3,RD&4la0��Ky��w�sr�ecRlj1��t���&$��6�ԓ)$�%�E��W)#Jy���FJ�Q�K$E�v"2h��ŮsE&2h�b�F�b'"Q#��!1Q㍌���St�SQ�+�ƌ�<����&��feH;�#m��QIc��Ih(1F6"���㑨��Cb����sEo����^:C@h�L�#D�E�rC$˻���-�`���.Ah�&h�H�Is��=}z���y}'����$s����6}b����F��Su;��Y�z:@,����^�F�j��aԆD���7ݠ�Χb�r�,dn�3�/��g=1_)��WJ�>�N���K=���9V����l�>Ʀ3/D�l��|E=߳b����}�ώ�|똒w��Wr��{�G��y�i�9;_?:���_T�sw���ܭ��|G|{R�ЂW�OI���������X�o���y\3����>�5/S��a ֓���%��R��F��D	'�_L������2��%�����-U|�=������3sO�;����O7>�p��MM}�I� 7�4j�>V4����*��{$T�]�m�M�4i��q� �p9xΩ�Q�[S�̗�0��xi�)er"�G�|�D�����{��׋�^��C���j;Ӭ�k�@c���ƅ���t�ߡ�o����{��vS�ǜ�Oxؗr��Ox�m]G\F���p��g�sR-��.8*����ޭ����ð�|�L=�^��
]>'�:Ez���5<��sC\��xr)$���%�j)֕n5�,-���|�"3H�݀����c4�I�x�z*<�
��}����6�mǢ�'�x7jΜX�6�h�y7*�k�ޛ�5��8�I�o3�]��hBG=��W�֦�(d>�}~���D>�w��^V�\T=3+9�"�T�2��w�b}o籼:p��#h��x���5���1��Rs�#��Ú����syHD�MM;�Ozo��(<�Ǔc|�ԇ���9�ã��Qԭ/���ww��u�t�:�@��EF�����Lgl�����+Ey��v뗤�˙�(�(߫#d>0b��z�k��>wţ�x��ǐ�:��йGq��s��[�}>GF��'oY3Տ��j�<��];��T)�Ɋ]#zk�Y���}{�x�m�l��n/i)s̆g.r�Fq{��Ej�����ډ��^�t"x�~Q�R�%/zW9�c�</5��g=��/(�_��*C�#��<�Ys�ɗ}�I<@�s�d���EOs�>��P���X�~�S�%�m��Ӡ��t���ȳ_q7��c Oǹ ���3@�x��w�zG��y�ͲnT��OoW�=�����]��ʈuU�W4��q >��=������Ģ���\=}��6��l��*o:�6\�ϡϗ�����*TʮII�Q�Ol���˪��٦���*�N����/p���M��zK6�|�q�`s���3����{�{C&�&�tuy�z�.�4�<"Z~ȇu+SP\����ܐ���/u�x/bDr�ZdU6pf��#�SZ܍���r�+�%l��zp�Z�G�t��ЙUd��h]:�7ҧgY���π���Jކ�bټ��\'\Av����[���OV�<��$_���8�,핿z{�{���U&7����r�c���K6�����}�)5�MA?yJ��W!���%���t�_G������֒�n��놈��Uo�B�Ld�� �>�^5�8�c�2v�LvW�}�I�x�=���7w�@%�Q�sy'�O�v�MǛA���C�M�r�V���wQ'��l=4}�J�ӧG�;�O@	������%�M���Q���q�'��rcY�z�|�V3��#��Ä�>�����D���뉞���?�%��l�>���&q�6z_n�f^uc>f�N5�CP����Yvb���?�lZ>�O#�P�CٯW�T��Y�O:l�bq�N�J�J+�L����.lÍy���6N�b�</�2���v�(=��E�L,�C"��S4���'|(��M���pZ�1M�T�tt���=(ήN��%,o\Eu!æzXC���5Ur�Sͽ�3j���n";*��������x�q�O(3`�Q��qǖ�b���L�a2nLޑ�H�`��,���g+ +���eAҢ41�������,i-LF:%�W3xa�r�ᵕ�z�s�^(�gL9O@��%�)�ݷ]y@:؋v'VP"p'�v�c/�5-����ڡ��F�7}(-��� ��Ջ+�ރh�����u���/�<���z��G:�a�=� �# ˡ~���ʓ��+��{����p��xn��Q5=պx�g|v#����R=P�W_sHK=[��z��~�]��G�
��'���[�ٗo>�y@@�9Рv����]�.���ɻ'�P|ߦD��u:c������I��@�����$=� d�;�(R��}��ܩQ����/h�KT�ј���Yi{�t��(��uB��)����Dfv&�#��U���Q�ڑ�sQ�5>��&Vw��W4�x�2]�,w:��.qUk�h֙%飔�Ob���f�^��tl�)z��N�%n�+�h�߫��T�w��}Θ\q�^�P5�D��_E���{3_+���}�5�&m;��G�{�������]V�s����\sR=������ �{=~P�|���骝t-��7</Ч�O�����ʎ�2��Dw8ZͼI���*���s5��x{�1{�����I���3�c���M��_B�d����
�\p�Է�K^g�gM����Qwu ���n֛�,����[{��*Aw�]R�B�Sgk��|�.b�
,)8�Ѥ�&�������r���B�i9��&��u���C��ή^(��Mj�2�X��)%Alpc3��E㡂1�}��N�Iv��띺����ua�o[��o�W��K󜓙�j�O	�>8���ұ�}���Ju�*q���N{rS�6����N�V=��Z+ϲ���6N�A��*⎤��_.�;Z�>�Kz��L�����R�P�y ���)9a�'Z۞�ho��n��'J��AَڋΟN׵��wo���|\#�ƽ2���-P�����yP��],a�X7�O���2��c��_�Eg
r_LS�2�b�KZ��J�5��~7d��m�9oTw��ղ�.e�{�=7�s�<ȣ����D��x�.Q�r,T�N[u�lKv�����h��+���!��ڟe��ޝB������c,w���2L�@_�{*ȋ�X�o��X��9��9f�lW�A��F�F>k0���Pp����R��}�@�Q@�'Z�Gx��1ۗ@_J�h�S��5�qf�'"��r�;�	������TCT�L�S�3�z3������`��#��/�޽��/,�x�4���Twv��}8?����r��S�i��F̗�y5��/0W��\N��s/��'�7:�
�Dc�x�|{�n��+Ƽ_{B��\E 	]�l���!���Qf��r�*�wV.U�4�]��]�9����҃�9�v��.���V�5��t�8-n��KJd�K�
��},�]+xBN�upG1��ٺP��nwH9�pj3]=��E�q;��W�sO������Q��T�w�Y(������cBȮ���g�q.��{n�&ˑ���60��;fĻ�������uZb���Qnz�Lg%2�ޔ�o�����gH��a1��Hj�����?li��6Q����sܫ����A���؋��A�јg�{/�V��u7~��p�I>�A�{ހ�VW�)Θ��d��Z3E�5+jy�A�Z��6�V|��7��>ǫ¼흶���`!�����1�3�"��)n��S>�q2㠲��ր'���"�r�A�cݒ�φ=yZ<�|��W/I�����ǖcg-��l��c�6�?�%���MG�@�<�Q��Y���;�\.uˇ�|+ϖ#���o=�{ꍘ�.&�f�Z.~$�_�,)���J��;�a_��x�{��h�{�Oj���g�1s���=[�pr���1��%�=z���B'����:�L��+����������3�ّ�NyǾė�dlz�<S�yQ�e�32�x�$���t�_=�4�w��Kz�k�j�[�&w��`�e�ج�f�BYNW��͇wz�Wl.J����U�YE~������/2U�J�;�=���2�Ň����zq��5�U-� �olh�8������Ӌ�P�j�8����d��R�lN
`�ٓ:����ήon�eEO����4<v��6s�:��䳜D�c T� ì�]r+�9͛�Ŋ�N%��/�{�_N���^�kkQm�2��WQ�)s\@�A#g�����y�}���t2oū�1�U�_o:�7��l��s��y��3�T�陓�r��[bg����,tm{���63'B��l^@<ʋ�*:���h�Cr��n�2\t�u�����������p�8HmZ�k&H݌�.'�BY�+ޞ�^Ƥu}��Rb���F�+4bͯS�*v2��,՞K1�O�W1�.�Т޴�X
�|�=�*Z�Ӟ�?lU��wUU�=�L�m��m/z��������A�hl̀������
���;��.&������.}g�����]�[��3�uhT��Ǯ�b̻�b�%�o�sA���C�O�D��ٹG>S�0����v+V�h��X�"��s�o�q���;�Z0���&�1��=I����Q�ב��l����~�`�\���|H��	��ix�9����z���I�d
��������	��1��a��
�p�sd� %u:-aU�"*Wa�@�r;��*jn�l�O4�y�m���wQ���.F����q��w��n���$���uk=����k���},pN����H�y�*S�#	v�R�G�k�� ��}M[}gM�{��M�͵��Ν�JŰ���5�pG�?r�XxQ��Fk�f����܏>��$�j����g3*Wj��Iw��_���D(���r�OC7��D�.�?+�v	�����6Y��E��(SPv��k��q�Z�W�)�ʖP�4xv ή�wM%,o(�0�G��_9�������zyՋ��D�>�x����s�Z;�8�
"��ߣ�A�Ǝ*�^[�nn�*䊾�-L�f�����|�K�����jޢ=QΩ�nOq gN�o���si����Κr�]�
�q�x��v��狀�OL��9;V���Ү+�K��������^
�.D�q�G�S d��s�
����Ń�y�t������Γ���HdLg^��rq�Mw���QF窠�D�L��s�5�S�,��}�%_%l����]��|>5�mo��T���8߉�9E�QΝB�R�5�$v�	B3�Z>G�Ҽx9�Y������U���آ���ᾪB��ɒ�,=��}�*�/��4kL��S=5�'R7�6;{�*_�T�0�3�S��FǦ�ݩw�s�B�u���$�v��x;9C�+���#������3�ݽ�Y�e9�w�oDh�t-��F(e\����������Ś�R��8��EЃwvx�˦,s�P�5�2�
���K����g���tN�wX�!��Fx��o���w*F��4.i��㌊��P�fg`!�}��=M_{�^�/�.���vZ9��pu���WQ٭,7�@�.�pY�H��2����(�	�ƨ��BX���C̃d#�����Ǫ���e}^���.�dw8Z��Ę[��]�R�
w��8͌��X�ߦ�V�y�%R_�1��V�	O�𜘼�o.8\j[���WF�;-ƃ���m��dT����ӻ�{[�~�,<Ϥ����PuC7Y5�t䟕����s4/�ɡ�nI~[ڨד�Ckw�Ĵ۝�&�{~���a��Fc��8��KM)��n(��}��;�u��2��m!�j<y{ӭ�辶�u��=kC{�#:�I:T�Ӗ+�R��q�J��'��� �8��3�j<Z�Q{#Kw*ٿ�����ޭnO;�>ˤ�Y1�}��u�M?N?�p	�|��ι��K[�q�3}��p�K=��I��Gye�[�v3���gE�s����<k`��}��R�P1�r&!?����7-�:p7�����t�e�/�3�4?�б� �:�z���V�1K�&�̯l�3�]v<�c�:��Q��x�;1�;��u�}��Z�6�`T�K[n�L�j��/�ɤ�,a����U�\��!�<���'5�1kη[b�uUc�%p�&f^�"���m-P��9sy����ku�uT�u��,���d�{������z���
�NU����4f�����Z3��fm�>8�B�R��i;W�@�5̊��/�='1;�e�R�=�6�`'_��r4w>\8���l͎&���P�;�\�jkL��@Z��袄et�q^���/S�-��(l���Q�ݴѦ��]�����s�`�rV��\;�ס�h�^ә�Sr8�˃�ANb�U�Y�5��+��Q���H�zu��7 y���eNmd
�uے�^�n�F�C�١��1xt�j��Mv���b��{���;��97s�}��b���d�����} �n��kB��I܁�����?��������~u2K�?��S��=��G�Y��MMS����/��cΡa�n�Se�$��z���:n^�`��ح�T�0�o`Zh �g����V�/����>��:���XNe�f�}�:/��s:&��%�ݥ��Mu��{	��ɀ&�����ֲ.'��>o��/�ѿoκ�`�f� 2������d ����48۷tƁ�h]���,���].s���P���A.���RK�Θ��Xڷ]C@mt��_�^*u�������/��X���hC�w�<!]�dT����R��V��5Q�ԼԻ4��$$��ל8iݱ��K�G��Sxa��S��Pe6�b�cX�Ϋ7τ #�%�ͱ�&�n"�91`L�ԩ�@�(Šv�<��90u�Ap�ZKծ�&|3����O�庐>ٸ똳N�NV���N�-����K��ۮ�Q���	�o�J�����(֝��Y�����]ZIUӋ�wu��[C"E���V�i��ۈen��``v%+b�Z�y,�j���ʾ�ж�:�غ>�xJ5����;�_�n�V.nV��\��JI����N���st�7{�Aai�����qK�}Q��-'n�11WYAB�5qj9��e���&λ�RI�ҝN�tNP_sю�w��){;+fݶ�^��}�W����+�9�~��L���]p�!I��d�����[�B�9hp֒�m�l+�ر��f�`V�R�<��ƹ��P�����.��� k��X{7���{���x��4z������Eg&��{#u���`��$�'m�&�5l�1��m�w�R�k^[�9��e�����ü]-�qN�n6+TTtf�Ӹ-[�U�jJjvI͍��V�E� �or2�P��*|C2���n�8}1�|��1!}��S�#HNg,�,����[�E�;��٭҂��M�+0Lyg9��K�_��]�=ego3\ʼ=���>�n���ۇp�r�w��H��U�Wn��I0D ���u���G��+V�.�w�U�[{b�� ��v�wtF���G���Ên"9�	��<�����7%� �j񛝉�D����ښw:�̔
�z�	��L|�ӽ��|�+�W�\�V%d/��u"l��g6�Z��������R��[B���"�եk����*�SwۈS�5j���c��������B�S���!����5|,Q�TB�
�z�۬�n���I�.{�Eb[��ʱ˵-I]�W��j�ec�.����9}\��R�>Uۘ�4�ђ��s�`�Nc�]69�����r���E�O �A��5��r,d���4���*���\bΦ_�8ɊӔEfn�wQ3��v_q�2fK:'v��\.�rc�i�;��e˽{f�5�E���tHβ��$�mzgP�m�F�um,��hWY���/8bh)�Q�w�A���*�7g����{zR^l���s�و+Ya��8c�+4��0��Ϲ�J��c8��u��Nۼ�K
]e�LV��u �ż��u+m�o��z��^�Ґ}o�X/$7�<��]��Q�D�hi.__T�TJ�j�k�����g�H���3�ԅ�{x�t��r��+:n ���/�K�0��WM��3�]'r����ˡz ����[��i#��H�,��˻��2�y�r�TS����LTWwUr����t���*4��yx����M����W+������f�k�\��)+�;:��tj]���[�s%�v�ܺ3��.�nt�wqE�!�s]�.Eˡ�Ü�Yw\��\7wl��V����Weu:Qlr�7w�]:�v�s��뮧�n[���r�MNu;�4t�W��h�\�9͹�.�U�;\�X�`�ӷu"�2���wqs�9�Qk��]9���7wV5\��wD�<nk��n:�NnPQ��s�5��x���S�w];�Ѿ�_}�����vh�K�wG�KX$����ܮkW"�^gM�[Y����N�u۱���;��(T�r���]Q�w]�NN�e[�d�����3�6�%�G@�9.�@,�Z����.:�e���r�6���O3�q��l�H�?��I�2��8{1_.��5������(����r����2r�z��N��=���O�װ׺w���w �0�¾S�E%/zn�P鯻��>}ѹp����ά������������}P����0�yO�:L:<H)D���E|�Ӫ�,�x���{{�O`���μ.5�>;�hx�[Z�s�P��f������@�܀�Tq��ruM��W��+��ٗ ��Q��&�{���z}��ME���uU�TsJ\��@��'���\�V��SY�P��<��aȽ£�y�q��76�n�2�WV�w��O��ty>�br>��?S�I=�-�5`T�����T^�Q��Mn^���\���N�J��X�E9ӗ�E9�*�FMN��!�|1P_ON2�';�zϾ�5#�7��Lz��^��ci_d2��2��;t�G�@�R��a�Q��{}^���weyAʒ*(���?X�ћ��e[.�r��2��#���^�4��囻���om{�9k'C��|�G2p�2WuX�N����9���Wu�c���3!�ҥ8��ΦK��7t�a�e���c,���Vfۗ�����w'��NF�&���3�2�{��\�hx6��
�-�:f�nX*\/�qj:FN� T�e	��u|���.�N�<j��Oh�ʷ֏���y�=>�!���C�M�(ek�Z=D�(�ӕ���ɷf;^q��>�q�j��E���l�]ep�Iv}ɍf��L-�<�
�v��w,�dI�^^���vc#~/"�}>ng��'J���&/_T;�+Y�Yź���^��}�L����l	sE��o�x[�G\͋�pm����<C���a������Bv,ְ�
���W;4e曞��γ�y��Ӵl��xU���F��3��<{
��N{�8�Nޅ��v�*Ӏ7�j�����)���+��T�Q�N���Ҍ��Jgt��E#۠�6��>��?/�������S�4;�?�X������qθ<'�tv��<xi'��@gb�Q,�m�_���;�qm�S<5���D��e�/����5��Dz��S�O��L�{-w����y�.�	�=r�O��� γ ��+]�������;�̋8��n���F`7E�p,~����V�^��j�wGR��APeYeŉ�B�ݙv���mn�XI�d�έ�]ub|I%C���Z׼ϯ���=�q���u��ç%Z��1sΙ����R�m�8�T��w��S�;��olP-/���zF��J��N�Y+P��'rwr��#�~���'TeE� ���I���c9΅`�{�\���Wq������r�]M��<�-i-�8�\P�O$x�;pH?�e
]8Ϭ5D^�HsȜ����[sz�*ج����u7���5s�P�9Jh�̑�BP���MG�Ң[|1Ѷ&k���ݳ坒��Op۩)��!]ܙ.ٖ8���U@Q��Q�IzjR�|���e��*�v%z��-��^P�W��L_w*F��ʾ�L.8ȯc��
5�3:�(fR??kX}���^��hs���5�/��=��T����߹����L�?�N�7�t\�b;�SO~���H�&g��A¾�s�hz|:��=J{���x�*+Օz�?��Y��
&*w#)GRr�HQI�U���eq���$�}Q3�j�z|:M��?��<+yq��
8�12;�v�Inf�q57n�^���g7Ϗ1G����{�x�+��zެ��.���^�8,i��ݭ�v�:K@>�+S޸�O&�칡~8�-}����D%q!���<.~�J틪����t�2ա�:9�I���jʊ�!��>T�Gm�}��}�6��	A:�]K����[�+������ؚݔgSw'h)F��Dǯ-:κsC���^�J����=f>6��N����J�ڽ=x5���P��l���5��u4���Y���(�;�����G�6�y �ykr��4��kC�ޭ�T���t���H�O��R����EӺ. �Q�FwD#�7�zgF��-P��[�����c6{գ��{�(m>Zښ�qo=�Qs&�ѳ�I�p
T:�3�1%����\g���؇�Y�6�OSؼ���0>���C�-�.(^�:��b���韢�Jf8�*Q�1�r.�S�i��0�qè^��ة�Z��eB��v(����;]�Q>��ݸ�S�0IO�I����оS\c�G,k��4��ť�o�7�`ܥ�,9|�.�g�Y��j�|�B�R��i �@�<f�&l�������M^��M�"��[�ܹW�ϫ�nt�������X5N�Wܒjj#L��{���(�GEM�{���1%��V�D#�|�0��{t����h�͵��r�z9X�S|3|�}\�lyg���؛.mL<�=�G&����Kg���=⽏�q��H����J5͠1�Q;�K}�_&j�����B^���d,j�]7���6I�6'\���Ox�U(�֐��k3hum�M�pW(j��]�e�{�:+�Yַ�,���<�h��ѐP�	'�`��w�gG�S3�k���=��[{�m՞���圮ҺH�IG���w��َ:}�� �=�yC�c��ᠨeV�`�Ϡkx�lk2�(ېf�ޡ|T�MΗ�Ezr��c�B_T�*���.7�`|�_��f�N������v)~>-���C���@�I�7<{Rt,?�.ˋ��h3_?J�ẅ���Tٷ�I�{��z!ZxB���V��L��ߣ�/@��mF	����z�����7�9A���c�ZB��k	̿��;!i]��p�{0�f ��p��/Ա�3�['+�@��4��GD�c;g�ߖ����i�ǂ~ԯ{�gߩ���o��9Y#�c�f�>P�rAI�E��� \f�����q��s��F�Nn�)��>��vFtL�a�ň�tF�Q2ơ3��L����8�2�U�PכE����왢;�O޵9��(��NQ�_�wN�7�j`�0:�|���J�fc�燭���<����G��{!_>��6���z:t[x�9P�T<��/��z��ф��8��¬���k��ƴ����u3�?]��n�P���n�-��9q�����|j#�:���ڃ^
<�$h+��l�7"�&����8���LrwB0�TVk������:������j"�DeD:�૚R��쫷��q1�3f�<��T�z!���-˓��o��Ցu��p*n��|�Y���u�1���3�9�97�ʝ�r�q����_�2u��T4x�����o�`�K�7,ө&��iK9]���n$J�=׳�J�_v����t(wk7�ȼ��X��Q����;y�v�dS x��3z�6y��Lv{�:�7�w���=��9��5��g�p��;fo=��%�[����l�%%��R^�|H#��S�,z3�{�GV�����1��76:bX�y%])�5����W��Ѩْ;j*�2���4u��cR:}�qR��ˮڢ�z7���]Ɇ�_7.��Qp��k���pNQ�=�����V�3����}OE�7�V</��!Q�)����{�Br4w�(}�
��}`ΐ�k;E.�=�4|Ǽ���fĚN�q��e��G����TG�����4���C�M�(ek�H���$��W����Z���nG�3J��U�w�:�Z���f�,�+�YZ/RO�K�ɖ[�X�\�_����Oa��eQ[{�-#͵��=�O������H�=���R��ɬ�
͓��Oa^Wѻc���^��j����ꎎ�2.NO1�Ɲ�����'�jkg�ڼ�8^���J�����u�w��G�۬��aB��E@>1����8��V���j���EJ]6���k6�����]6e�E��4�}���3�lV���.Kkɖ�i���,8)T����`p�S&���hֻ�:�|����)wZ�u���״��(F�ޚ��y36l��V��4�*w�wV�X��b"Of�*_�k�=P����ͦ�ۥ����zb���qA��(�-b�@����k�n^e�j���L���H1�[���K�뇊;+�u�鸞�����Qt���/��[Usr
t���ƜLi���$��V�{�ٸ��_Ny���G�����)�����Un���a̚�I�?Lq!�!�Q��zрZ�lM�nШ�gp������E��=T�����=�	���;��9Ιqa�*L��|� q�P���ưu����q�V�9P�N.�k�Q���9���|�_�w�Q�35A-'�_t��)�}��df���S���<�f��O��2�x���b�z#�:�Q�4kfH��s�4n�?TV3y�ٷN:yu)����ڑ��t�wK%�2�����s���]�F�L���j=���>�F؎��z.�C��o}���]E���]sL����P*��{��'���̮�ݷ]e̛q ���M���Y�ȿ<:�j���������?O	�ǍM���c��h�v��@�c���=��/�o�5r�ڰ���=ՎD/r��*.-����;<HkHcgf�#�R�N;�^�e:�{J5h��N�v�q!ҧу���Q�b�n�n(C{v�g�}�ֳwP�i6�����.P�r��T�ƻ�ە�`K����k&��N�����i�TB��>5㬯�ԣ�3e?��1�r~�����Z\w%�o��1���f�?t���L���&/�i��3vY0wpa'�#&w|��}kx?�]P+��f�nS9�{[�~�!�ܛ�a�	�
�x��3z:���m�tl��k@��z�Z�]�����ڱ�7��Q��KMѲu@1�q{��A�t��f��d�f�7КĴ���8n}��ޝnWSL=��De|�բ�����k�7���!�f�ٳs)�'�5�A��Re�zi���^-B�������ٴ�1�P�8\wn�ǟ�/rN9��i�9مjQ��@L�2Z���3��Y�����k�����,�����MW�N�i�퍏Pg�p�*;/�ղ�d��D�2
�b����u2���X���w-�yUS���k=���v<~u�}�x�C�k�W�w2�@;�2:A���ҾS[��<&c�Pp���s��@�D����u�h���zY��[�(�~��}�5�8��.��&���x�+(c��lij�V�J_A\���F�=��y��7��ҵ+zG�(0e��t����_��E+N#�����Y��mE2T̫��(����j=�����X�t�]������g�9m��������JťJٝ:���{)$�,˶�z�������Ԋ-WuJ��?��MY�b�ܹ*7�W���]�3c��m`�;�Q�))ƚ��E��'w���{Si�{���Ũ�<-\�2��
���|�Z��P�;����V4No݊��B�z����8Az����N|}((��aW�y�#_x���5[�q���Y(���Ћ[��靜�c��Qj>��yXkf�5,m}&�f��֝駞ci�F��3�����p�}�~=�:l�K���;�`>t��1�f��@{��iwS�ƛ�F}�P¢��'�NVEe=�3�)�k�����To��5���+/�����6n!��=Bj�v#ذ���x�-��O-ؓ4�����}Q�.��Vw'�n1�M��έ!mω��j��O���7N.��=t�1�4��G4�����z���e�d\O&3�}�`ۈו��F�F8������Fg�b�?]�"����Q�Z�:5�4.;C#���t�`�!���S�ӓ�6V]EzT�ezr��]�z�8��踢4������ي]#����vU�t=�e~G�F!����L��n1\�Q隹��=*J�ꂃ]�lDӷ�Pre�vM�ځ���ʍ��P��J���L�*�ތ��CE̒c��O3k:���s�oW׭9�#��}��P�����{;=��Kw�aWn���`���q����ú����=+opl��<�������u^�Ӹg���T����P�V����`�s#P����9yo�MJ~�z����fkj�ߡ֐�ʕ�D.��g�^��P�k�Cn�pg�_�O$U:��L�g]o_����^��|r���փ�kߏ�_���uo����税���W&�d�����|�o����&�{��Y�ON{��{�${>uU�+͏)䳳s?t��\i	�s=:I9xD�����-d	�¯qGV��e���>�>Zcz0�В}A����Z�m~�km�h�9O��5�Bt�a�2�ߊ��*:�{i���s2ЅjUEמ�����s�%��`.j�����GI#�>�8�G,ʹ�K���ڕ8a7��]Rr<��R1P��Pܸw�Qp��D��M�0�#���^b$3^�K�z�3N�Of.~�mXb�w����C����*T/��k�d�T�eP��TF��O=�K��9���5�ǲ�Z��/G����?*�o�����Y��}�[=jR�k��,D>�O����]������+Q*�����I!![.��s�oQ���9��8��ǹ��.�!��U��}ǐ����6t- eb�Jt�6Q����Z��=]��y�J�۳�K0���Z��:��%�+6�	�3{��̣k�e�\�:�ϟ.��q�y�����H�X�f�{}��n�68� ��f�U2խO{3u�t.�:Y�u�e�Mޘ��ՏYBZI!�@��Ŏ�������-������vt��`�G.��hl��		e.�h��^�<ի��9M!����Y������[�#.��6�����X��UM��[ܶ��[4��4�,>Yi�W*��o��Պ�G���]^Ք�S�&�ֲ1|Zۣz�E}ݱ��Ӡi�a9��Z���^bg*��iu����<��UtR��F*�v�z��V���A�郹(��D�f]iw6̋��@�ĵWX[�%��Z�vl����:Gha᡽x�o0e�L)R,�n��D�b�=�E2������sj�H���Bސ1T���egU���b�*u���=����\�:�$�(�
��r��E.},�P��Yy�+C��L�v[CH����1	Ġ2a���Z�B4�4�kw����Ղ���+�1��*'�R��^<�-rm�`;p�n��C���:U�:�9�\�v�[�e�y��:w��([7�������
5[I���J$@iAՋ�̷�d�T���1�l�K{%2G-�9|�zѺ���UV��7XZ���.x
篓��AZ���.ù��EǱ̣�X�l�������Ù�����>�xƘ��)2���.Yfh[��s)�V�NlBk]>���Ӽ�[c���<�l�z���8)�͊�e��*٬��{È�[��nd�z�nEqtuq��`���Ru0�ɓ�n��Wo7�uk'4<���a�uP��ۜ�*4l?�to^�w֭eBs��X��<�����%�\����iN�U��4:�Z��gw�0�;�����U���fM����פ��4���9��kLоǥ�Ii�	���+����][ 34E���+�"y��(���X�E'�ra�w#KD A|�Jٙ�K��rj�j�6�͇�����lQ[!Y������F�0Y����7�8=��R���l�F�m4'r�\�qf�����J���G�=���f\\YY[78h�29�喦�܇CG�tE�'3]CY�����2�}g,n]u���F�,m�P��mb�A,�c���3
��[�g]�	e��Y���R��h�V�z�;3Wu��{�}C�Vc!�u�K)ٜ��^��V�����N:赔�De�]{�z�]s��nv�6a�N�^�,�,� �Q]ǖ��Ǉ��`d�˨VYLpގJƮ捤����$�m&rM�A"X8*mIk4^��d4.whow�Á���e��.�t����U~O����t�76�Ԝ�r���ѩ��.k���)\ܰk&�\Ӽ�ɞv9n�y���tC��;�����\�9]ܹܮsn�y˗]�n'U˛�G76.�x��.��1�����]ۻ���ۚ���;��������s9��,�u���;�\vػ���wr��Ƹ�*���t�u��]�s]$9�wq�:'u.:t�Ÿ�n�w9�r!+��v8�u�����˥dB�t��t���\��ˡnww+9���Τ���w.\:Ww;����w��q��L®��M8�$�v�s��n]�r�7K������I��NN����\�ηw]��]�b"��;n[��@�܂]ܮ���k�]͹wqK�]�W.W
��T����#��	N�Opw�TY��j�>��ӵa���z�t���ݢ�c$�-�w�'\v���$�|isd��3��[s�U�rG�Q�
�
$�&͍g=u���ԓ�wK��ĘZ$s��]URU�N��f�D���]�#뇪�������
��H�$o�z�(��חnox]���1�N^�5[�N�"�����ʏ:�3V���k:v�*���)�����~�+��뉗&��M7[����s��0.%�ls���Ӌ��.���g`_����[V2R���s����)�����;�Z��bN�(f�5 V�LKm6v�����+���lA$�^�f���}Q������˰���xk�);p�V/�%�����θ=7ִu�#�Fǫג�9v1���V����/툀F���$�>�3�Y����M�}%��ǚ��[�����r���a����c>���ߓ�t
�A�˸�V��o�߲R���Wt�;�c�����=�g��7v�x���p���t�����K5i���0;� �8&�|T^5��Y�wVQ�}��5
U���y��ܻ���s�x����9N��B�'�<j#H�����*��?��f���Վ��yS,F����.̟��#�� �s��ŝ�;0B����^�n*��=�?
�*^\�+�ÿ`5x�� +��skzÎi�G@5dT��O�̈́{q��r���0@�A��]g�	�\� JXJx�(֠�0��Fl���W���̀�K�o�F�w:c��{E����Q�E�\��*�)�_l��'�q��ux�,i����'�z��p��ҫ�������Hwt�[0���v4��P8����}ہI�ɍ7��紮Y&����Nb��6��w��?W���#�,r�t��㌊�Gz/����|�/P�.�'�~N�co�(����k���5�=�ѯ�Q���u�i��4��J��i=2��Z��(ְ&�T�q��JO�̃ś^(b��O��������꺎B*�yx��}s)���z�Ի���=�߿R	��e3q���O�g����Ԧ���ݳ�a���o��k��v��h��_%޸7ε��)��c��;�/��9'2�õ�i��8bsE��)8�&���������=���s��N���o^-}���D���Hr
��	��{��8�.ꍨX���o��7"<y �7��+�SL=��G�\>�����s�-#c�m9���]ˑ�>$�Q%�_A�P��Џ@�5��Xڏ@(�������sL�_�Tn��
�j'����\%����n�UVE7�����7�l��n�[Ԕ�Bܻ;��:�w2��.�ە}�8���6���s�x�s)S�YvIyM������+Z|w_��-,����v'��G��d�)e-�V��[���J-�7H�m�V�ح�|���D�Z�}��u:	:Nf;!L��RMo��\g�ӳ�ԉ�����E�Rά���O=��7����C��y[.�O������Q<L�T����u2�ө=���]Na���}����/���~u�}�G��j���uLñ�R�@{>3�@� gpw�0,�q����<��ё�[˻�L9E�+����g�֌�6�	����u]P���f����k\d}$ݽ�Tc��L�w$�"9�Xd>�{�#�F���p]�e��g���6�)�2 ��/C!��f����-_����2�d�-FGa���W׸Tuom4i���.��c�m����4�]�l�bEt��Ϊ�j1+�1����&���¥/O�����eGWv�"�S��z�5�чh�Qz���+F4(��Xkd"���2l;�c˚�U���if`�ۯl{�}�퉤�<��b�ۅ�i�pOތd��Y���'��^��ǃҚ��U��9���yK�;F۝�%CG�5<��9g���k���O�}��J��=�K�Y_�-v]��+7�Q���Y���cof~xsp!�A��c^��{�c�:��uu�7봑mu�V�xkugf:kؽ�����'`�V�X�4��*6q��U�cW�q�jr#3�����&+Hb��pqve���)�Ħ��2��>rYcD�3������9�L��97�x�6�Ɇz�+���u`7ܞ��d9ɷ鱮�!p��gV4\ú�7g���;&�m���9��"�;Q\ ��{L\rKY��c;g�ߖ��1���.�Qͅ��A��]Ƶ�pe���Pgm&��#������ǐ5�dRٗ����e����ZY|h��4�<��\G<�}>GF��Ӥ�1��3�~�7��U��B�K�^SW�xK�r���?��:����'�l������2��[$��t�:�cNn'$3���G�y�p'π�~ڗ](oX�LX���y%�o��C��������qnD:<L_f�a�ƽv7E���~ށ-#a�S<5�w_���{�x\C�/�\y��*-�ƣ�:�q���N�,�%�%���W��`& z����lB��L@{+���ߥ����|�7$_��h�DM�v���\_�'/#�rD��}�N΀��#�{�2y�Pc����;��w���=�nV���j�8�������3��Έƥq^䔞��� e�kB��Oac��/J�£�S2�ނ�ݟm�z^Qć$V�F��F kۺꟻtL}�3:�7��{�mЍ�|b�/�Y"��avb� j�ns����:췻Lb��k3�������ki�yo��Ƒk��,Ϸw^&"�:,9���Cz�of�g����j�W.��>�x����OC���2�rI�Q2Gm@�AD��(O���f�nQj���+��OQ����j���{�n��:b��Т�]���s�=�6m[,�-�ɣa��	���O��*�zX�oW��T�Gy��[,=�P�j1Ũ�wFN�G���]KO�y�9��.g{��u��i���1p�Q뫮�V��sA���C�M�r�\�h���{�a�\�o�'���4}�_+O�Gx�>��Tz�+��jI���C�q��P_��\�8�)v�O^_�s��}>D�����
��P��||:���Go�ڢs=U�yW���4�x����/�Q�G���3V�7���X�@���6��|�C�5�}~��=�f���n��h�޸5�o�l�|��{/��4ǟy-(Q9���C��"����o�ξ/���G��=P���l/E4�ۇKC��Zc��qGI:9�����{��w�S��̵b��������x����}p�0��W��h�/1"HL���6����:k#�h��KB���xB��C��ũQڻ�Iѣ)Um���k����҇A���U���J�[���^�5T�:�=U�ʭ�@�»�@�Y.�S�w�n�P���Z���lꄑX��q�Lo��],�i�Ƌ�Ԝ]B�~~� ��c O��P���L��n+��{����K���@v�f��J��L�V��/m�炏R��O��� oJ��H�PT=Ƒ�<��wz�j>���^S\�5��0�G��ap܏��tG�Ү=p~�3�Xb
�S$�nA�c�ҍ�;��ns1Y���z�M�X5)={Wq��w��|��V�AʇUL�_O$x���@�2Aג����u������3۞��{&�$�6�9^�Hu�����,�>�k���
j�B��)�Q2GjBf��T{�+��~��-�3��}�NV&;۪G��HSmi.ٖ;Q�:w�X�?J�+���ݭ��d���I�,�(Q=���-�*����T{��wJGc�����t���5��kʭێq�{�D�	단暞���0�~Z��#�Z6:�����uZvu���UCdFc���r.�`l��H����}���z�:Q�eX;:]����Խ�ر����S~L,�Q;����=I8���]�<�N3�<I���R
�S?��sy?�Ǐ�z��������~҅��Z�!�2mА�}ò�f����#{����z�{ï���#$��)��[/E�n��(�j�3��^����� �]y��q�s^J���wa�s�������so��)Wy��3X�o+~�=r�]��l�9��Z���'9\��D�s�+�ё�?\�u��2ϳb'��Q�:¯~ɂET2�(�0���Z�{~�3�#nv(���K�c���dϱ;D��S�p/���[�ÏӃ�ϲ��;-��8s�~���N��31� �a�.KMB��}���ǐ��ZܯSL=��G�T3�=:5.{̍�':&K���eHw�N�t��ٜQԌ�5�#�7�ze���ǐ
�F����8橐r�W��nF�Q��Դ�pۉ~�٫����' ���Jgvb�kx��Ҹ̎M	��P�|��������g�nI�Ϫ\V˱��<{I��t�`0�k9�br�]^n�x$�ɥӆa:g�?:�>����W:�a��k����
��c�ÃK���>�9;�*�c/y`��=�Z,��ў��a6ڃ����9ʖg/�flנc�i?zk6� v8�/��/ǜ��H��hq��[œ���=�;��|3'=R�n�ݵۤ��L����5H�0[Z�B=�޸�1̨�£��4vkA�N����˥�f~C�v!�N�ot��c�T&�ǡO�Hx�um�,0Vu*�f�LS�u[�,��!{�YH�&�����e�(C���or�3C���p�sMo*d��_�J�y�j�fU�@��o7�i�aV�Y���
}�&L�h���[���R��l�p<�r�:��䭩��fOl���X^R���x���s���,��;���͛*��.�2Qm�z9X
1�D(֬5�crM�=;��p��~d��:Zs���Y�T�m�&��)����u��T�_8���ܸ+�ԇ����A?(���;!���//������h���&/�أ�:��(��U���ʾ�s��{��+-����]���{$�)cIXf�y����`���k\]��1��k��.��O.�����{�=sx�;7��/SP/�<J�M�_k����lL�;�|O��ò�>�73�#Y9�\ ��״��KYɌ푝�cge�*�ܰ�wѰ�z��~��)�~��s�}'��7e|gmB���|�@zj<z�@Rg�HS��D���'}������?�Tn���Σ�m����踫��k��L��2�b�H��񕲨g:����ԿQ���tx�n!�l����=7�"��,�ղA�X�t���Nȑ9�3�>�|��z��S�2ov]l���c�,_�5���r���y^�c<��G$�S$\�u�l�ʏ^N��
 ^���lh�P��A���".�^,��N��w__03��zX7���/��#�8��G|��r;.����U��gjJ�����8�o��w�Q����u�s���pV�k��O���7%ΙŕLuw5e��x&�>˿�)��_S,o.�#"{�x>��G�r���|k�:�e ,������[T��,�E�� y�1�r g��1�v7Q5=�z/�֞�nH�ˌ��8p�z];��#3��Z�Oj�B��Jzj8�����-�6K�`2F.�	[q[m�*_�.���t�+��q�s`�Έ�t��_rJO�{g"	'�hR{���{�]q���Y�,Ѥ\S�ٷ2��n�q=a�sT�3-}�$v��ӌ�)���`x�x�b~�ݿV�%[�)���W�T�]�T�osE���p<�r���
 (�i������^�?0����e����+�teڭ��ixǗ��^wrHoy��[,=P�k�qjz��z���W�o�²xɸF;�O��R������p�^���f�Zn#��f_�^�g6�����
/Tap��}��xtZ���I��w1�R��=�|j<u����z�x}��>
����2��;�8?���*9��>��� 0����<w�Z�`:;�=W>�K/���JExW`ћ�F�[��=��X��o��N��Yn2�7P �f�%��>����.RS�s������
��}���Y�Jg����^@N��R� �ލ���J��Yu��&��F�2�r�tI��e�����"7��.��' �W!"�wi�&>�Y��O���Mg���2��V3^s~S��G\���Q
mw�|Zn6�����ѱ2�츆t	��;<��Λ;�N�=��i�{���l��3��al�}!z�0�*�q��݅���J�Q	�gj=(v׏T �����M6v�-n+��T���g�����v��OĜ�3˅)����7�#�F���_U���D�>y,<�u\�~s�G�锣ʽ���� �q���:I�f2��P��S������l�=��sk���w&q�y:kw@�S������\9��I�� oJ�N?�=ơ�̮�Q5�L��~�U.�g���:Q����s�wO�3�x�E�Dy�\{�	f���<�@��w(�s\�X;��vj��++�jVl�K��Z:�'�w��+����j-���꩔L�>��l1��5�5��@s
h�c�0�|�f�Փ�7�U]r:��p���Y�.}��su�Q�T�C���{��䞬�./��.a���$��Ǭϙ���ث��b%wy���������������?�Vֵ��խ�km���kZ���ֵ��[Z���j�ֶ��kZ����km�5����Zֵ���[Z���������5mk[o�յ�m�Z�ֶ�kkZ�}ڶ����j�ֶ��Vֵ��M[Z���umk[o�kZ��Vֵ��յ�m��b��L���.* <�� � ���fO� Ē��=*�! ��T�"����2��*$*$J�)ADT���T(R$�(U	JR"R�TP
������D�κm��HR�J�[4ED�s��P�kD�T��hE*٫[m���)N��R������kEH�T��(Q���j���u�"D�V�Z�MS6J"UJI*�IH�$P%	�UmfH�*kUAZ�"V���Em�7@�lj%
�	UC�IS�  ���;��e�yp��6���Ek�B��f��Uu�t����Sx�.7��ܽ�������;w��UU�����;���k�A��A�U ZR�M2�"�U�  �}Ks��)�펏i�:��u��ͩ>Qw��Ǣ�(��(�qEQE��Ɗ(��(�����J�(��}kǢ�QE���@ ���x 
P�P�i���:�D�ZV�e�7�  �Wz�US���Ԙz���˕V�ʺ�{^ݻ����WM"���K�=y�U=�=�ͫ�]v���^�S�K�vf���^�=�Ul���IT �V�)��  �k�w�]<�v��{���B�1�m�������W�۫m0�;���{��ǽ��7�pm���F��^Þ�t;ũmWm����ws{{��^��K�k��jQ6������R���T���$J�j�    Y�h�k�8����=�[[��G�z�^����w�n=*�۶�m�����m�U�=��]��X��vݲw��z�����m�缵�ol��uۍ���yz�{��r�oj��owM���
I*R�H�a��B(|  ��O���m��޷{=Vٮ�]���ۦ�h�s�=Q�ow��8xwwd�{��J�����޺y�벛�ݽ��BӬ�����Խ���wmz헵�b��{�kM��=5*f�MTJ4�+G�  �|�v�w6Y���O[��w�{���w�{u���]���];�yC z�{m��/u���Oe;=���{�w��ޭ�����!�4�������۸�n�W���C^ڂ�D@>   w�{5mN�������F���]�����Vި��TZ�v�̼�;����]s�9w{X�[��M�UJ7{�����^��y[ٻު=��shݽ���^��yu���yC��[U�b���e] >   ��澵7���V���{om�;�k�{�'K�]��w�4��{͝��n�t��C���׶��-軳ۭwq]{��U�w��������;vO[;y�^��r���ݗ�y�vj��f�����҅o�  �{����=\z���׶�y���5���p{w�=�{{����w�I��ײ�;���{�]�{�V�n���L�����N��oM�w�{Ͷ]�۷����v�'�RT��d ��a%D��� �oL�UU4�� 4 �~%*��A�!���	�UT� i(�
�z�0�	�?/������p�W��Ve��ax[��pn�������35����HINg��BH@�y �		�!$ I?�BH@�i	!H�B!!��w������?�~�~�_/�e��V:{B���;�gn�+G�fQv�c��p�ܭ��l(�p�U�ǒ�խ�x*�,��wwa���J�5���Q�L��x^ZZ]\.ۉl�6�F��F��6�j�a+YC��Ղ՘䎒�vʦMsHFc�f(s'd��b�Fa��2��1���#�涷
[K2�
T�p=�r7+EF�d$�Jx3e�5ܘ�&*˃
�[x�Q;
��l�;o(�V��G�Yt�ַml׀F��Єm��Z�-�\�U��Cv4�ö�&n�7��0cQ�Ya��X]핡]�iK�%ӎ���$���\7�2�V�v򖗇æ=5�v�n�L�o,�5q��x1f&˫J��m�n�Dm�Mޚ��k]@]��-e$�/RӢ:Ϡ5��4Reh�m��d��qf@�Kڴ��Cl����Ԭ��#)��H�F��ڂ���R{��o^f��+#Qf*Ya۫��f�jȢ��+��:�-�۷"�Rh���ىn-Ғx�T��܊An�?k���k_bc]7��"̲M֭i��zh�̬� G�٢�!	s)�F���JYf�R�ܾ��a� �\T���!�NVm��s���մ�ͦ����y��
fp5�P(/ST�؞ɫv�C�e*y��GPn^��i�2�u���f�
�OVh���\t�n`!q�!Ѝ�XQ�I��I����JxEb�\#2�R�3��b[�&��&1-S��q��X9l��xQY�a�����\Z�t��\��WN��K��P^�#�@�&�Ōff�,���박��n�B�R��!��2�֚�h�@����d� ��	*��u����͌�U��n�ٳ(�R�d�@X�i�sD�s^�V��;tp�:�u�Z6��H�ZtX!ioH�8iY��t�@��I�(�6��~����%eE�2<'R(��1���F�ַ��h�QJ�{��W$uueIb���ukC;��ieA$� �8�br���٩,�)�0�T�B-���Q5	���H�5S۫�>�mb�&�l�-�P��e��vҳ�z��bn�قf��,t�[��U����V�Ĉ� 	`�[�m�lƥ��
2؏jԳ��lۧmԦ�tS�˒�Y��f�-�b��6��I\l�%��NJz�ͭۥ��ǄaF�ꄔ5K1��[�[,���(,1Y�w�3]9�_�*���{{� Hhƶ:?��R�	*.�e�Tv�JÇZ��E>�Awf3{�q��A�J��k(��w�V��S!XY-���4<#:��ѕ[k.�kbc�,����E;�#p�*9���.&�6�U��wr͇jU���C$���jS	p�M�f�
�X�R#)\i]�^жݰ�n��/	�$��IT��桐���:"-��%aƐ�U�l$E�j^�7�M)i��u	�7��*e1j��M�[a޺�:��ᥰn�pA%GH�M�%��ѡyr:��˒��1�/+%aM2.���f[O)�����ŠcwZ سkr�=OR3]h�'W6�h��J�0!��hh�.�nP�
��E��G1�ݬ�_+vE�MǙ��ֶh	%=(뻗��v�J��?�5�C6x�����G"�����`�h-Ď
	��&b�l^&�D�v�S���z�pC�!yd���0��#������n`�z�I��W�g�Y�$vqd����Y��-"�JZ�����p����Ь�WB�c7񌽪�ia�JښZ$�defe9uXu�WKV:dH6�mG��i�)�9�E�1b̅�����T��<d�}5��rRַ[sF�|��,64�*=ѯ]��=��f�ٶi5�������(��xZ�nA5J�!Ve����Yg��bX���z����Ɲ��J� ��ÈT�t�S�j�����Z;f�%��*�˥sm�+)������6�F@��Em��F�a5�(�����zqԒ����^'���(��O��Ժ��k	�.�B�D5���U�[��aH��o��%J���`$BMQ��d�{�6a����,N���(��a��D:u`m cL��vֹ�\�LT�Ʊ���)���kt�u{L���0m�!��Z��6��AI;հ)K������f:+_�@9Z,��Xݔ�<`S�p$o)֩6�u�[�KkDn�
켰PL�vH�P9ak�wE����b+襶Aֶ�����Bv�U&n����N٭VjִS�c�Ķ)Q�%��S!3���h;�� ŮL�F8d�G�Tِ�[����*��.�ٵ&YE����-;����<Xa4��)Q�\�2����R!�(��
�7����:�q��oȋ�)�,��%^c�4Avt�e^e�5(���2���3kp6oe���ec�ɷN�ZذH^�����0�2�<�"��١�t &������/XH|N	.��*�N��1�U�%��M�);�{Z���
ʐJ�]X�&ݺ�v��VT"Vƥ��:���'���u��3�E�wy�RQFRZ���:Z���m��,��u�Z7+*KOE@.�
I-V����lPՒJ�(!��/l��)�b�՗A0�SkL�k�l�]L����	[F�f�n⦒�A��wL��.ZW̵oU�&��dD��#������sn�Jb�/b�F�k@�;�\��iM�#wn,G�OK���&Y�IX���+ˌ3j:2�M�A��І�Z��7��Sr�*�63p��=�쩹A4�$�KT�bN���aе�*k�or�Ӛ7j�l�X��˶¢޸U^�D�x�1���͕�(����ԥ�l��̡�c�tV�F��ZM,D�E6��ˬ!eI��"��dMS��Yм����n�<-�%yYt�Ă���)��n�^p���ͬw��8��`�`ɲ�H��o6��D{C��D`Q�H4쬫6�������]1�*[9�A�Vt�j����e<p����e��1���q[A�%Pme�5�<�n��-&Շo �ҷ�m-�L!F��^%n��k������W!f)AF��v��xD�݅*��;גqKI���ӎ�hjW��k-���RKi�o���hGV�(㻩w
�hjQ�z�m�(�j�OF*�����r���ٖ�1tqlw ���Zl�%��U�c;��e��� w���kє�Z��;ĭR��N����kq�!�4��(a�*A���-`�2Š�����.���t6��E���!<��R쥴"7l81�Z�`���	en��f����6J;$�4��a�*3uZ�zk2�n�vC�Tښ��0��C2�܄�2�-��t�s#U�E$�����cY���ǦJ.�^M����-m��)U�i���Me���V��ߖ-�,5���(˖���r�W	�+P�V7N4���� į4�6���-�I��"�ڪ�sQ̃u�)!�_-�%Y�ն]�2Y�,:��U���� �sp&��Թzw�IEoA���c҃i��Ɵ��aI���{c�,Ճ*��م�N���i�S)@6���:��d�/f�R#�Л"�	Ft��3�K��wo[��c����^ ࢯGA*?5m�b��2��,�`*�m��V�Wb�Y�k���&��<@R; z1�j|��Y�1�@h�KP��q�Y�f`��ܽg#����d�bl��R��>L
��6�
��ZE��j��6*�1����)��ey[��E5��[�*�L�/kUMyyþa�y��f�g���uYh�\jA�p	d����8�ƅ1� ;tp���*
���"4�g  /U+a���\��m�X���1�Úo
��6X�K��P�St�ʁ�qF`N%�L�E�e�bע���ͣ,РZZ$�x�H`)!* ^J�*�'eU�Y9-�h��wu�,��m�F�Q�ĄCM�×0Җ-e���V����3)�/2Շ���1f8�X�q
T4S2�����@��%�����ݰ�
"&��&���L�)�����T05F��2�j-<ժ��r�ng�X�Π9�U��.6�w s*�becw�]���N�Y0�mY7���n��T-JG����ܤZ���P�2� ^�kq�F�l�9�e�9��l��D���������0�Ô姛E��i$�ջ�N�0*���-�4-H�x�z�`ZeDP�X��Ht��6hG[2ZCh8/5B��f���e��۵D�hV��rq�-O�k�-Y��n���8�yu�����%\oZ٫ՠ��V�\1^��;�"J
�� �����6l��jQ8�8�ͼٕe �6���U��4�:��i��Dd�J��^*�)�+e[؂�'�uӛ	?T�%�25��ͥ�n�͓+Z53bI�AԷ��F�C�HMDd��Ĕb�v���[���wv���y�w�檖*�F��J[.�0�����-'dC-95]�u�#�-S��aO2���xۚ�l�wY��nQ��He�O�4���5]��f^ �"��V��t̰�k~9�y�bCx���.U��,���l�b׃%��ײ�E��([pV�L�	�-����)#ixU�5��w		���)r�H�J�k˹��u��?����m,7V$�h�btHܣ��),�Z�Z�Z�i�Usi�lLK�z�ڶ\4�j202����%n�WŴ�]n�����*���h.���j;���ɲ�ck�*	h��-;��QQ��Ղ�n�dk� �R�*U����&�1wR�o]X��,�z)�-�?b�p��X;���e	BY���1w�s
Yh���ZP����`h�3a�Lm������tT9�n��[��V�BPbdRJ���Ѭ�g��n�Z���wz2�n�y0�DN�T�ں%�^Los�+��k�rQT2��VtcYJ)jM$��-Am`��P�t5����DN�:+ҟ'v��o��*Ԡɘ�л�]�3�ce���X.6���Ŋ{Y>GC.ct��+�J������v'&��f*�n�6�ue�-j�e�4bUm���Rw2I761�{j�����@!��C2�!v�$�.�C�Vl��MբO�d6Ue�; ��+A�W����*ڀ�c�VF ���b$ɘ4sr�0섅2;�L�NӸ�x�P/2ej*�f9�[qk���X��b���1OU������X!�j�a���en\�Z��DV�X�Z�%0��#7͗OU�WZ���s
X���a�mJ�X~�MrκCX�jGĬ`���AbF۴HЪ�i��Y�k�����D�j΀*��T�;v�Kt�+�BͰ�+V�m8m�Q:F���7yҩX�����3J[rӛ7M=��-h��11�qѷ0��
�����f���i	�gě�n����V=ln�H+���bUڦ�l.^�;MS������sCˆ����!3hYj��4�v�yv�Un�
P�gi�[���k@�H*6u��Ց���Mb�%֧������ {M�CKN�X�:	���4#-�D+46�fF� .-r�V^M��oQX����KpŢ=�^=��-�����*`�u�o+VC�*݅�AA,֕Ae�ce6w�.�eI�`��M��e�@v=m(k5� �i�hݶ� 0nG3����V�4��"�CF<�r*�Fn��Vn��_J�։
��crL(���*�вC�k*i�aZ7�`�h��(^�J��*�.c� �WI%2�E岀z�WtQJ%*5��B����YZ~��t`;H9M1��YX3%# �!8C �*{gH��Z��]��j���맶qЬ�alK[���tv�Rx�9��
2�n� �+��VV q['g2 �%f,�;r<'�ڴ�C`C����a�)+���rң�QaO+e�Z��ـS4i)S6��Y�R\N��`�#���]�� t��vI���I��ѹ���:�E�{5#z5;^�^�)k���X#��ݺa�G�U�z-ͱC3&$�ҭI�Q�F㖥l�)|�$3W�n��<r[��t	0�x�a)	�ٔ%��֢�9����	X �x�.�g⊕��.�.^�䖄�\X5m�ǚh�ZނL�&������λ�)�Ҥ����%Y�j�dY�&&Ž�؅���m2�1R,������D�A�7�m�4m����KO]&z"9T�M	�&�fL?mcb�x)d20b�����_3J^=��F��e�M�{�f�^M�뙴���!������qT3�[z��Z�H�,r�5a$���,�Lں�W�k�3@]kӘ��[I�Ŗ-���*� #t�Ӹ�0���cӪDJmfP�̽ԫ`
�u�����ƥm�N�ɡ���N5�N	X�!rXe"(�I�l�E"31��	�n���.؎%�	�&�B�)F\��<kU�`b��CA6��FX�wV��t[�`hm�-}�J��컑����o^Ɔ��A<b��e^l 7i�R�?k�,�f��i�V�=�����(�ҹ�1DK!��tD��j��w.�9�j��e],^+��@�D��(���f8�Zc�qPą�Yr�:	D��I��V�yP��s&Syhԩ{Rk�������,�� m�j�ff�9���Unen����X*U�4���sY��M:I
bVZ��ǆa��{h�ڈ_�n���4��Ij�mf��N4tk�q4�ښn�aɥ���ز���ЯJv�e}t���&�J���++���␼�E���l[i���R�1 �SϤ��r�1���P�j�Guf��Dgb��y��-v:�{�sN��V'a���m�[�>ە]�F�9֢��]mq�"�)��c���{ˎ������9��2����95SwL*f"�� (���8��\�ꁰ;t-T���jy��yYW�
�%y4eN!���W+s��p�Y���$7//|%tӨ7Ъ��L{m���G^�]!$I	�����c�iy�C}/H��X��!c�u���Q��N�n���A�"D�}�T�-63)��ޗ\��P��e�*<��*��Ɏ::�zÆ������NNA���`���˛a�\!+�WL��jwf��ǅ2�Wt�Ŋ�ٙ{P��S����X�,)1���7TZ���`Éf��Q-��(� Px��x�!����
�NP%S��i��JV%�t*�k�d��J����&�w.���YCc�+���Ε��۷|6N�1�Wj��K��wdA�w,7�M��']�(N�u}C���/I�0^b�&֮f��Z�������JOȯt�}��z2�wC�Qrǆ;�]a�vCǹ���mQ�: `Osa�r�1�t�\sH�#N��(3�n�>綺-�C���b�7�&c�o��L��Fc�kw d�0���z�����]���U�Z�4��N����&6[{��7����.��UNxv��q��HQ5�γ� e�/h]e�}8H+{+E�HE�
,т�d�-e�K��Ux.]��i*:��F���x��Ә�+��ب�D�vga)�+4��W]F��"�͓1^��S�x,�(P��ˏ��ͥ�D���|/�9�n����lK�1�9����Σ֥;\:TV�R�sN�VLu�n�ǒ� c}�4�=����b���mL��,C#�����8�IJ��nk���7c��Z�'�cr[�WwpMV�����|���=(�PX:�)ή�KŐ�/��8�y�Y���@�X��ǅJ��iR����Ϊ��[��[�)|uR��Nvy�.�}Hwq2K����j�5�n�w����kwӀ��lC]F(d��_[��ZXE[(��`�Xv��s(&��D.��K뿸Z^��;[�!!9�,�e��匡S
��0�,E��#j}��p<^!�0`�i��tM7!}��9��s�c�X�Y��z.��[�H;T����ubY��&�&_[�1ڡݳb\Fe�S4�5����g��؊,d����rV$��Fau Ŧb���:P�|���s�P��5Wy�U�42^8�١V�M�á��45��j�5η*e<!�;r�]�+6�YYH��v��T�����ts�nMz�*ıWCє{bo�RًF�ֵ2�r���L�h�hhϠ}]�U:�N�}��^T��j/v�	�!�dv�E�=�-�iWq���)�Xa��{��F$�.[���6&�ʾ��U�E�.�mf����T��d;�*g5ͱ��G��nk�R��:��6�:����z�
�z/����"��v����X�T�3�e�2HY�٭	ej^�{u{�)�1���B�A��J#F�5ha��j�+��V���� aƴ���5`vcΫ��dX��OZ�vY&ҳ���`O��]���GI�
{f�=�P֖�'u�۸mZV:�'���Xw�dc��B���,��ڳ�w;�a����5@1ÁK����]f�̳N����E�͟8�v�Lo��)ۧ��,NI�d:+)=*#U�-����qu��֬t}F^��9uh�]-`f�I��_a{W�)�0.�f<_[|�RFՊW|�{rL����T4"�:-�^N���;Q��N��S���ݻFb\|��=p�V�]��ܧ�>d7�m��&TS�}B��[���3��r���8Y'IZ{�՗i�{h��ͽ��F����N�`����ɾ��¥,� ��.�ys%N��pU�@�oL�aq�1���'�p	j��:M��P���)B���=�jm���U�b﷚��ؗ�Z��Y�/k�����D��Q3��KHUñ�b�P堻�m�]��z���1���:����jq�I�CF��FC{��-	�(���GW�{���Yಽ~LJ<��G�`X��b�,�=V*�Jn�>�6�pW��a�&k��w�p,����:�c2`P)�%�NBumpW�0E�ym��O�<����p���w2_r!&�A��|���,�-�`�Ҵo ��m�AM�h,!���rsv�2ih|��̺��î�����ؼ���x�C��|-��D��A-�<l]�q�M��:�ʓ��0��}n�]Z�^G�V���R��d�V�u��1q��b����wf�k"���o����C#�]�畑M�-ZlgRFLE��k�md��+9�%b�;S�C[��|�wJ+1��n:�/:3�9q'ŲJ�B���������ΫɐU��D�
��;��x���%����噁�r�fd�ӮB>ߦuJ7���T�����orT�;�l�Q��|u;��K�k�Km���f��bgf+����>�4�<)Ӷ��$�lAN,\�E��C����*�YtE��'-B�aYXoYMV��JO�9m��v�#�̅�����U�n��0f��y�A�;�%��:o4����F�tU6��Yy.E�+.�@fo,MS�;��N�1�3QTh�g-bކ��,�Ɲݶ�uu`�o����v�jWn� v���2�&@���e��L�{���N�ŗ�����픤YV�Ѓ&��Z����
t_>�0v��ܷ@0]mX��n��S���W[�Pp:��>��<�g�RN�uW�N���,��8(�֧W�*̣��8_TKgUۢ:�]y����d�:q�|�S��CSN8���R�vM�/V� q������X��6�v:!�w\��Z�E��Q|N�.���%�����d�U��ۣ��TvA ����/��O���'Y�Eq�H�
�P9x�u{m)ePGb*8���<�¶��}��cKC^�}�=Smu��:m�;�!+66��B��X�)�W!�B��gȳW��v�����-�I.G�ǀ�ض7�/�w���1*K\ffR��r!�#�V.�TnPx2��i��y0�I��XGsھ�s���^��r��$�E�^[��/�[�	{�.[v��dl��Ö��-��ɴ�ޗjW�%�F�^ޖX��斻���t将�X-�Pm�Z/%$��)m=@gt�XRf��R�u�����w�`^�Ig�+3�A{�*yD���t��RUvD��0_-Y�Ӊ�:��e%��q��ӻ���+��B����ДA{�]WQ�4��J����e] �֖��yV�f>����~/�:�Y�WR��nN����c��Zܮ�H��ɖa��ޮ�b߷��:�wU�q8{8���V���+P���^�ޱ%�$�rC���,oN�ɕm�<ˇyN�x�DJ�:Ĕ�Y%,��(�G���Y�WCXF���C5��rEZ����50J�e���S6�V�54E�<"���ҝb1.̗A�zn��*x��dyv1�� ��WʳD���}�m]�+')4k{�c"��5W}��wu<��t(�؀;m��D+B��r�̅0r��p� ���ET�W(��rlj���/^��B��T��{c\�bg����m�ְ���׶�j��@�^��I8���t`�E:�U�G6���v�.[q
�zN��p�]#N�:�x��������(���?�Hb7�sF��
���"v��8������m�Zu3�*#�%;���Ծ�yj(җ-�j]�M��3�p��"�S-?����҂'m[�Y��\����{����is�t8�����IR�6�h�n����PN���f��{�3��!��λ7y�;!���]�!]�47b��/n`(h[3o(�{t���@C\U��Vf���)B<�x>z���t�緹�����
����a�n�q�uaRe�yEȷ�k�CE�ۖ�g</��m�	W�*x.ѣ^ѾwFy7d�sP�l���A-yjgp�Kwʉ���N�Ҟ����ꀍ/;g0�sԫ�ȓӇ�j�B��IE���R��݊)Yn���\����0ȱd���c�aC���nj�5�OL��E��G*3Q>d�BJ|�ΏZ�ݺ��l8��&����Ɔ���=gme,�z���G�l�l�pO���kY��w~�.C5��n`X�o��GJ�ݏd�c7^+��rI;E����ԝ�b�VM���tU�<�H{rx:�Ȧ�ո�� ��@���K馓x��7m�2p�.�`�D�ϧpxӬ�f���!�����÷oN5�,e\��Z�}�:�<� ��+��f��YO~V�oK�X��\�_saq��r��3�3-u+�G�m�s�:�c�rF���z.�����ӳ+h�6��yIs�'R�{D��#��|�Y"�ձ�/�\w�r�F��V���M|qCj�M�������qc|��8Ȕ>�����tU����f.X�DP�PO-uY�7��q�m*!1�L�_Y��&�� �f�ֳ@�P�P�֯m<���W%�hǙ�v>v�"�h�/3c�hq|n<c���L�S �[�*ݳww�7�s.�h�G����Ւ��1��70�"h;W9�F����s&<N�-Jٗwҝ�5���۶Q�Dy�
Wp"]:��s�]��9,`r�!����/[����|���4�С�{+thU2�%�}�;0Nn��� o��LZx�D:�:}x*��hd�ӹ�&�r��P���4�D�Pn�Y����1!H6:�澾w�ya`$�V+�#y,�\�ƍG�[�>0 ��ɸ�I��L�N�].�ږ�B<���2>bWnp]���1Z� %�e�K��ݥd!�¶�!��z!��m�"z�h�d^<gm��"�U6��WDygj�
y���}�� q�_b�c�p��5�H���z
U�fܺ��<�4��[�A���7B��#�w-�\Fou��I�[�Tj�1.YN]�aѾX���"R���v��^8���ُK/qY�����g���`�6��ە�9�?6G^賜��On�t����єP�S����=�̧Z:v!ɴVLK�=x�NQl��9s��<�e3�T1�����[6�w+������Р ��w�|�+���K:]��>�g�y����``�a�Ng�Kuu�"�!��Km���:�5��F.7s�Y�Q�A8IF�黋�F$\�q���t9#�3�Cg\�@D�.Ũc�kJ&i�|������&P�uj�#�~b�4�X9,(�Su�f���@�ܣ������]��s��N-����g��[P����;�~�e
5��{��]N�M�-i�-����\�z���+h��+�2fia�]hWo��v\��Qu]����n�0��v`�Vlƶṟ���A�Y\�ΰ֎���(����&��s��*�^<�XxN�s@�"{v�i�/3��6;�U����r}�/O;��(�Ij�x��ϖv)��^��;���k��0{(�V��3��g1J�vV�\���҉+5͔ݟ���ʻŽ6�zA!�t���[�e�R���Ȓ�Y�C�jʌ��9b%��z�[Vč^�|6�/m�NV�&�O��@�D�Q��t�3^:���Y�Y۝Y���,8U�V���ra��-�c�q��˨�\����!;W;�rN�Z��wb��F}i��U�;��:_3�ƨf��ޖ�R�2�D�t*m%tljO�s�(č������0[]�>�e�N�I$r���:wW]"�7�#s4%�]j�E]�a=1u��GA����6S/��y����u��+z����s�6J;�+6����p��m�Z�b�7�	�+O��u�:��6�y�d�q�Ю�-G��E�!ܸ�(i���iز@&/���&&/�SF�NVvX�E�o���8�u0Im(�eN��.WwJ���N{Kb蟬\�m���82
�n�)�[v8��E,ҨX��*��ή��/qS�C�K��2w/��ķ*�0f��yMI�S!���u-X%��tl;�ʎZ������r�Ob��Z��XҵǝB�fR����;"�X��[RLa�֫3�0�Z6�=2cL��3@;J�t+#�50m�x���v����z^���ה�y-n�	\e*{&P]Cʲ���i�eZ=n�p�>�p#�ݙY4����9�W62g('
�ֳ�T��c�OV߶W���=~C׃OC�-��cFV�x��"ۃH�y=�A��kx;��VdI=7o�,)�g\u�q����dsC�L�Gd�|�l�O2]�)�S
�I�N���@Z�h�����u�[G^�\]��~b<��n�3zs�ǡh9۴������5	�v�,.��y�gᐋ��^�ae�5=�н�Z�pvҹ&�2��)�ҏB�k]T�2���!���I^^��x���Y�"�������`���L��9�>z��C{1�v\#��y�5����v�!�o���lJ� �<)}�,łW82<95U�2r=����ү):uv�qٸ�Xb��h�7���-�B|̠M;B�@{�&��v��yD�ki�9�N�Y�l^�Y�������V��e���m!�����ө�G7;B�ŋ�����{;`ڴ�`>�k-v7W��x)�E�p�&�A��Թ�OӧT��I��T���(&ۙݠ��wǪ��b���e����f��6�m�E���2C�4=%��/Q��������yT�Ơ׍�D`�gG6�Vʳ{�;+��PW>�ǘ٥@*s�Oz�P��S���s�ǹ ҰI�A��Ժ�&�3c����@$$?�$�	'�>�o�������n{￷�i�+�M��kQ�^��@��7*]5h5@m��a";̽u���_|��R�Rj{r۩3D;[�fD$�ٝ���A�A��ꭐ�L�z��$*�A�ێک�Es�7sk$H��ͬo1p�	��7��\�9�Ԝ��.�`�x�՚����q�ڂ'+�è�b�sV���ۖ�ɝ3
��2�򻷝C�A7�����u�]�M젬��z.85ޜ�u$���ű�h.�z����ڨ��5�մ���!lc/v�Á�z���@��z_HFB�K�n���ɡ��75|حF^Ư�����%Y�)�(�UʸTW6ю�E23t#è$�:��ke�n�w���9�W�,0o�!�y 0p��.���5���X�l,����B��tr��N)]�(V8��]����*����=�ˌ۽���o�fٲ�V�s$n��.6V���`����ڏ]Laځ�H�wmΛ��"(�ZU�5tlXӆ�Sc�UK�K�TVs&?�w$#�l��rRZ�ӈ.M}���M�X6�,��lk��Y�2*SP�.�t8@��_!d�0˴.���b�Q�۱��då*��3ѼR�ߎ�#�N\�h�s����ՎF�jiyZ�S�����ŜM�9��}�����
�Z��\kp��-��&V:�j2m\0�rv��t֪iL"�=�h�����F�[�gC�Ks$U���� K�[ɛ�t�9�_�vx5L��,��]u��S,
6s^9h����/A����v�3>��}��˹$ұ�7V�ׇ(nj�F����Fd���W+��`w`�����f��]���(���z]閲��e��u�M�Ɇ5��Qm��Hd:�FB͜���V�^rD���
�U˭�3��G�ɖѷۙ�-��Z���S��XZ+b�t�o>QT��"�H;u��pFL���`^�>k���e[�Ò*f�'q̊1öW)	��v0�;B��Ʃm<��k�1��4d��DI��=$/}fi�m���Z�-2�ah�Fp�ɔ.�#Hj�2
ާ���J��u�b��^��d�']�3F���X�Xle��wu-�>[�SK]%���T���qC���2<l����'�:��}LWM,X�k��7{V��4-�NUoS_mJ�gP@;�]��(��ɔ,�r`��(��,�Hā$���u�%k�rZ�A��Ñ��7K+��b��Ι]D�]������4
ӛ�z���i��3�Jݴ�����r��QQ}(�4@��z�|�(�
L�9Ӹ۾UݭvK�]� �
aSZ&���
�ť;��ɲQ\�+g38Ԃ�q 7�]�yԹ&�"�5n��W^E�v3q#q-�%��a<}�F�
�b���Tq?�믬�.�G����`Bf��{`X����"�t��]�.�-4-� �:�{JF^ݫя�^
��a�y�Ll�`��E�����s�����1}L�K��5�YGk�9ʇ���'{z�&�#>���nئ�dx�P�g�uV���%wvBWIuͤ9
�ʓV`��œgS�U�$y���4j2��Ȯ��-��nF3>|�Hu]�_v�n�9��gf���J+�y�"�ij[q�5э����.q�ϸ����F�:^ 铦]h��]YsAz\�b!�s�m�K�؝Xձeř`C��o�*�F�}»WV�E펙2�G���-��&K���Vw(M�%��ֵ�ͻz�4��Y]�+--��Nˋf�X�̻�~#if��P��+�"T9[i��r+�t��WwVA��1��k �r�Y��le��t�l]�?"�m�f��YX�/��wn�}�*��5��v��!&vb�n�T�J�tl7��N�X�;��9Ӑ�1���F�7�w��ɂ�b+�1��B�<z�=��P�����ѽ�q���V�B'��.�!l6�/����^f��w���QH��t�9�4.�1_��A���ޠ��ۅ�U2�/{R�,8q��kN�Ņ�f��*�݅\6���R�6�a5�u��������ac�_�9���4�N��v1�������Sn���MՓ�6��8�)n&�ܗ#,){n�(���غWN]ٿ7�9�֌��"j��^h�#����Q�{@���
�m�%��2�=É9�٫�-�L.�7x�`<ְ��"���D[&d�߸�tޖ�r�7�kr��A_q��UB�Hs/xf��I��E�N][�P�j�0@�Q��V2Sҳ:�T��d�n�����YE��e���I���JK��mmֹٕ�j��S������5�Ja�m%A���C����
��C�J�ONo(��2�u"65��.caض����Y�v��X�J1.x����zX��;QYz�*����	����Sp�?46��1c���Z����:��t�F�T��@�e�0szYUɝ��82^���z���]p�q�H<�N��G���\�ل�	"ޜOxg<�;X�m�;C���7Ok���9���y��aqt�
(�eu�o��9O#�9?������nm*4����5x6KNd�j1�E���d�帆K���t��C���n�3��H�fs��cU&[��v�P���9g�6�4�+-Ρ�ˇ^WlR���s����#�V;��j+�s[!��<�c�������N')���qY���A����8(خv�{�"B���oYp����Y�|�8���Vmt�q*�V�1*�t�A[�������.�,�N�s�� e �*�Ïk�>��6&N�2����_u�ɻz_"�]�M����]o+V�W#=�� ��l-p��AD��7�0�#��!ބi�)���)r*�9�j�R�fN��x@��s���6��mS���{Av[���[�RyؑM��Ƿ't�s{@�m�h��1��V�>5����v�_Z����-;�Z�,t�"�Ko��mSWYW���΂�݊H"�#�w}�D������l���k�:D=������\i�*�y�GYl�j{I6�[�sr�m��Ξn&$z�a�2�-�YS�M��J+�h�-���ͦ�.��!-�&���I�.>�NY\gJįV.8���0?	�y��ơK��ܸR�%�����fMFZu��=1^����n�����z`t�����Z��x����o_(�������m�0���Z�wCy��%��H�	ٻt��Q���NZxu�wH�|�z��G���[�*�0Ƈ�(�c"�W"r�}��'�F���v;pG����r��6sU·�Wl�偕K6�^����t��ǚw��Hq$�ZV]�e���9��\�KL��z��9f8��b�4�#F�e(*:�B�{dV���ɜ���ڤ]�����|"��L�p*�ʟJv���ώCإ8f�@�r mxqN���\M+y�^�eY|�u<j xW0�o*U�>��"s׺�m:!:�;X��]���9��K��ѻ����P�HW	�u�����C��L�[�]��#9�r[@b6�a�[�D�v���0�[�1=�hQ�?7Qp�P��u��޳c�O��Q�w�GG�Wso����2Q}Ba�C����_\ށ����QT�2�q�H�ޒ�q�m�L�.���7����'6�3�XH�l�^1�:>w�����!�X%JF;_M�ۂ�Jӆ��BM�u�ډ�&,��N�E��CMfHj�H�^��v���;�p�.��
����-�ᯣ�5d��`{�K9Yݽ�Gzl��lb�@]�ȹ��9N[ݔ�X�^�hd];�F�ڛ��	�N�x��R��ڦ�e
����XJp�X�({v��Z_v6Bj'73u����f��t��Ԭ�\�@ [�e��<o;517��Dk�ø
��aG$"��n-��ޥ i�р��P���YW��ŗ ��N�����W]]sb�֊ś/2���R��6��u2 d>���çc(������u�X�g`Q����2o#���5�٪>�[�$�*�1�UE�6*�a^�#I�6���]��˥̔釄a�i�V�96u�5�ZM��ŵq�Q%��N�o�52��ѝ|�CS�릾��+�P6�b�R��nE9�q�]��8���{�l�Tϛc.G�n���t�Xr���DGR�rsʻ`�&�p��v����-d=������ͭ��Ɂ��ɩ��o('�`�����'�����wI��b*���4��h�[����+	gc�gn���5n͞��8���[.+r��A�5��+^P�,e�%�+hn��fW�Z�7Ǵ`Z%�E��%@b��9�>�S�r� �$�u*^ w���X:�u��]�\6��T���ZZʠ���+�����Δ�r����UЅv�\`����!r�۫�8l.�{��Ѕ��ý|�������ݨ����hf�^n��Hz}�#�o�pmʕ:f�f��*��[�B!(u�$�y���U��1z��ʊ��O`��.�\9��%1۰Jn�5bnE��c����O���k�&������mf`�x�S�%�r���[�#�Kn�\�$�7��$^F�e���%f^��ջH�C.�e��/9˛��w;I�)km��ņ�k��!��ŋ����Ip#}c%�(Z��櫱V!J���c�b��wo{�WIf���Jľ�TY�G�˯�&p��.^b��!��Z�3��P� �mT]mM�qs�����@RtP��z�陳>��T����jf��(#rU����\��n�b�@�א�ʱ�/*�M�vu:}FZ<�W	�i���ھ7S��J�#x�F��>n��'��pc��Vfa�ySO<��-.�kw����8Pp^���W[$��jޔ���8�@�pW98�!�3�dq�}WO��\�R��U-��0R���7��zx\��.l�O�:uH�W8�+L�/o�L }��C�B�]H#��|�L�������ǽS��oR��հa�������}AoR[T�E��ʉ�;&xz��=+��$�K���k�V�Ic�yu<���:�k0�d��� ���:D�˫�VN��5\��Z�6�Vq*�.1��)»�wm:US�q�-�B*)J��U�Ƙ�Dp��"�h*akC�a�\����a�<"{fM�,��r]�	�u��JӮ#e�C� 8�[=��z��]:Vi��\[�Ai��=��������m,u�1ΙZ٧���r��ߥ��"���l7�֟\`V;̹W����\�u��PS�8�υ]dݬ|����;��E?��*�Y{n�eЧk
ƕU�����Op�/ MS�E���eK#`�����@�]�F(�εV�q�����œ�;u�����4�:�X�y��/3�ut[L�)�I�	Ԑ�}H��OjZ�kG.�o����R��su�zY(��V#�a���w�<.���El���9b�Fl�qߨ�<.���Y�Y8�1��¯c�b��H�o�<]EV�7Ax��s9s[����M�u+z�3�x�(r�؜��J��b��1��x(�n���[\c�(m���>�p+�z��>Ts#�-���un+JEa�l��4�g���q���$�dھw�*��돛��F��^�ݵ��+�,F��(o0.�F<�t��9�^zM���!��]�3CM�]|�5+L�}r��
V�k0#�.mz=��z��<��m��'r�k}ے댵'��u�(���-H�������C�)��ץp�Yn� �9��.���� �I��d��!4,G�X�>�+7Z$�i��3�d�ss��:��'um�7��%���=�t����9�!��Ю��t�X;�X\���Y(A�i� ��'s���kH������]W>ڊ캜.'�V2˺uHZ ��eZF���XR#����6��0S\߅����P���+�	���"��9�{�2[�k\�^�w�E;��O'@F�޼�Kd ��S��LWwR�Nbj�:����)iԱʭ�w­��/p������{"ݓ����D��9դ�x�Np��}�ffd�}:��KV�1nc��sF����ؼ�X��g����#0�}}W����]��gvkQ>�L�8� ���v	2ܧC�Q՜��V�J�r����]�UEt]#MKl셝v�*-@S�31Wc՗�pή�%���YX��9`��Z��-g�mh�oƧ�`a�����N��/W$M_7�M$�[ݸyUՌ�i1x�@q%:�L�M�L|�e3T��s�ׯ�DL����G�9�7\�N���ܙ�5��MG��qJ����޲��.�� ̸�3+)� �y��(2�Jz`�W���V�ڵh�ڎq��j��Ss�e��]�2ؗ�^Y8EQ�/�8�^ݢ�aB%[Z�;��n��r�W��Av�W'��dt�jQq�@��\io�$�|HZP]�͸9>&&�9V�w��<��}� �b�h���R,a�]Ië(Xs�Dq�i���ό��D�V5��\�Lq���n.�Io¶�s�irژ�݋�$���J4��RD�C�8��|����f�U>8v����6Zj�ұʴ$��Y��k�57�D���!����Ū)G�7kj[ɛ�)��[}SU�O�PPeއ�����X��JÁ�37n}g#psolSƩSz�5q�7�uӗt��v@����V`�֜{�����v�gh T���)���w9Ճ�uӵ�'h���hY��[+pS������{{ j<;a8��\�g|�$V����ko�Ӳ�����w/c�/0�����
�E�c#e`����%b֎�ڔ��X�ۙ�䄐�$ܜ��ys��>9�5������`���X��	���(�2������J�+Jw!ǒt�jQ�7��br���b�3r�
�!�S{+\�=�hp��h�x�%�i��)QY��Mm0���Ƨ�9�5��R��Ҫ����J��e�=2��W۔�+�׽-p�~.��ǲ������-�%1�qmʺk�[x�m��\��p�Ũ�#����R�l�	����&��ֹA����7/��N�*E��C/��*�(��%�;�-TwHt�B��n]ɴ+N]�w-��Ut�L4���V��׿\�+z� ��n�W��S��-c�6��J��ۅA��[�xClMZ{QY'�i8(�0�MR.$��aD��/;���Za�v�϶�j}WR]��a���a���}�\M�W�o�J߂�G�~AYT�ԃK	�R�Ө���W��y;%��<�V&_E�
�?r�=��	��L����a)t���u�ڦ�'%�{�_uK���np��]�W��1�E���hB�5ln.�Q:�=��Je:L�<àS�d��G.���:y�8����Scq�LjM{��z&a%Ny!��Ck#l��*-ԋ
�E�p���yM$���w�m,8�I�����e��o=��gjsh�|P/-�nf�jќ��	�t�ي�Ɯ{�V�n�щ�U��6�����{ڭug>̒�4��Rn���s�}R�N����>ד�<(�QZ�O��k�l�����+\b%��ffKJT���J�F���cV��e�QV����V�b	J�E���khQ��[F�-�KeiK)�T��T�X�ԥ�ZQ��T�QUE��h�A2̶��R�j�cj�"�D�EPJԭ�����E����cD�+)Km����*�m��"��B��p��ѣ(�[F�R�2̴�����1E�B�V���*�Ԉ��U�[Qej1�EbV��R�1�ERҙh�F��+b�X�l[*4lm�
��UL����A���-�Uk\��X�mD�%J���U[m[T���X�YUQTkLnJ"[eQJc�����E�jլ[R��m��1�B�(�D�[hլmR��Q����Z��X�$R��Z������pd���VX�ѻU):e�� c�sF�X}V"�Hmo}���P�u�l��S[hb���x���}�ǋ��/�]�s��>X�=Hc�u�(gx���M3~���7;N^M-��'䂗�ob��	�`�/F	}�V	,����~�k�m9K�����[�W
}Y��[>����y�E3S��M湺s�C%�:�Ն�s3kirU�5cn��5/��X�ׁ�f '��IҊNF�)g7v;t��Zw[cU�J��t(w�n�ȏ:o�yJu_�HmM�A��o�r�ڡ2\�1�2�Ɔ���Qy}
?g
���u^&	#� ������u�9����'��I��ce�G��.�hv;%�]t/zx�P�z�ŭ��Z�:{��ڍW?u����D��ތ�9��h�۫�
��F�7�h]���5)�)�n�]*��X�{���:���Z�u�Qv\��V#�TF_�.�pOzyvtG��L�c�L٪[��pa	�u_2CY�B�^s���#l��[�ӏ3G��w]�s��������!�º�#M�����i�Y�>}�k���.�S���$�����$1��"�����즠�콚ɾ!�޳����SY)�,+���1��|be������O-)�v.��Y��Bn�ܪ�:ʋ���E�A`m=X/8�W���{ʹ��ub�Z�W+x+��ۢ캁�r�\�'UK���L_5�����1��t��Ep�Q��+���|�6�\8��޿�r�:tQ���d{�4jyi������;��poo�EUt供gW�����3���jѾ}���ap��J�8���u�����w10	�G����V��*�3o�'��NG���܈���PYv������Pb�'v�<}�g�νY�a�<nb��v��<cX�%oMJ�aO�պ��m���L&�5�1�Y��|f�ǅ`�&b���>0��g��yۨ阮,��)T�l�$q�'���U'e�D%"��d��c��D4k�{�[(%}c:���o��֬��{��9 &3�	��'
�8�{��O �e3��V�=���ͼ��� .���"v
;lb����6W�^x�����ͭ}K8��c�b�/��oRIީ�m#M1�X�#2��s�6u��u�"zb�:�\��h�͇�7:JM^A[�Ā�$�=�OYwv���� �0��T/4����|x�Zೕc�v��v���acB�ţ�f�<X��,�fzU�b=�5�ډ2�wI'P��ݎ?�e+��^WV�td�8�O��Cq�z��/��G�"C��'���� _�)���
�y���y�a�<A�"Bv��9t��]<ݸKv����^mW��J�Z��LTNrwҌo���`G�6�5j�9�3�-��r��J̨HM��^/�҉�����Pު����m�;i��S�d]���=���Sߋ/֝K-�5��ZNwVu]�Zv"��&"�<��M'��|��y��W���p�]f�#YW�,�ˍs{��v?��\��g�sšJ�)S޸L.��v�V����۾]��׍�p�X�wz�r�����#��}`g8i�w](���{^S�+�.��R:��X��8Y�5�A�l���5���V�J{}e��ޗm;;c.h��7<��4_�����dYn�����0��o�d�����o)�&���W�J�Kwr�d�W��N���;�8�����Ј��3�dh��X,S��'�Y��S��wV45�b�M^��j���ڷGe�z �4�3�Ԟ����	�vV	݄x>,Қ��M��e[>^�a�´̡Իvg^9[[�S�ǥL�m�źz�CȀ�	�4IZ�hF�ܐ*��S�Z^�9s�K��>��:����LR��q��V�pS�r�RPN�͞ݺ�����o�}�^�zV���`�q���	*�'Φ3yT�r���
� �Guۮt�����̙�3xz�5	��7��x��)`�w�iJ��c�¾ͳq�(zk�K�+���-ˋ���=/Y˘җ@�h5��t�WR��g�޼C%�B��B���qb�
�������u�j�]�J��3u[rw��I�au�/s%�V��R���aV���>��+�����OA٪�5�����mĬ�W��a~W�a� ��az杷(��8*�Ō}�&ΰ��h��yf�o��+
����s{@6��B�ħ�;ĕ����))�
�y�����>͝� �w�<.�,��\0B���L����E����0��lHF*L�%�E�Ȫ���3X�Ҭ��7�F���kz�42۽�w&��;�U�͕Ҧ�k�n֮�S����%2��)1|�ՁLr|����Y�º�f�����������e������l��X��c>'O`�e�ӣN�����"���b��]VhZ�m�����x�@���+�t�s�jN�>!��W�	�y�^�2��}�iV��MK�<�L>C����:෪SN����I���4���YM��Ŋ-��b/�Щ떇8�h��J��&�Nc�և�f�d���G;�u�ҭ�/6�*���7f�NC3W��8R��r�C_��voO���n��[�
V�'�P�ݱ���[9)#3T�n�3��N�ր3%*������z�ݐ��E�Q���'��^�/��PS�z���x�c���=0%o�ud���]����A�Ulz�fJv��t�ӏ���E�n?�<�v�`W����;�ҝ��|��ވ�{X�+�Ж�O^�*ߢ�Ѱ��2wHY*���(B�S9������f�V3뿂�jkmi�_�蘤8��Zhś�T��KI���M<���y��2���I��Uc�N(��
��k��P̘��-�N�; ,��ܛ�2�����m9꼮^����fy=��{��E��-h0ƛg�uM��Ͼ�����?ED媍N���*-��i9<�/�f#�f0�����=��O`:�o�ڴ�n�U�-�Ozu��7-K����(T{��og�EW����#���n�o�����<�gOt��ZͅR���I���z��d�:k��fP��YR�ޱP![8㐱<{��As�%ML����f8|��=�'wZ�Q��Z ��	�B�j ��Lڻ�Q����{��2�����
�7���`M�ԝP����oM��7�����x�Ԓ���	I�s���po��f۾���:�"+{�*�d��e��=X�-k7�7��s����@�44�^��4Ϣ��$7�A�uѮ��w�ꝓ+Lw�u�	�pS��Н�B��G��{���3��|�jx���we����/TЬ�e�O�k�L��D4��
u���f��Ǎ���bL];sQƀ�"Z�chO�u��Vn��[[�W�����u.
N�4�E�R�}�rX�C���ƍ$-\����j�Jco+[mN�)v�[��gt��Z���gw����7�`�p����Vϭ�\3qf>4�v1�WMP�2�-i��&�laoLR���>���~앂�k每��Yͦ��"�g����6���xg�X]�F�l�-����ʕ��8UI��e+��{U ש]�z�5}ɨN��0�Ѯxq�F�Ȭ�jk�<�ubcy�ήܹXj���7&y�u��/��`��j��o�wj�g\P�]�����Ҕ����pB�ŝ���N^��^�\Z����u>lwg��Q<ͩEm�Z����
�y��x�l9��^��GTjcU)�ڵnʼ�OwkKؼڢ�>���O�}��ځBQK�02�{��3)ǐ��X�}9�I7-I�y���4]E���y��ubE�gq�S���¡btS�w��,ۄ���¨p�=Rm��K���8i��fi{��hW�E��ա��h_f���R�;is����{>����/����Zr�$פ�UjRE)������<q2�k����{���J�d[�x�u{���R�S�Ŗ�����r���%ف^%�XO�����w�+�ؽT�X��	�K�Ԟ��_+��fߟa�輬�ju8*�R%7��j�=��6�3@d}�1sZ�}�q�<�v��Y�n��J�;$DVOh���9�Amrk������������w�z�Kd��O���b�N�g]�<��m�A��)��}Ao��Y-3�x�z�|Bt<6����V��g*s���S��^��D�'�oMJ�aMU7[G�ü8*繵չk@��Mj�6Շ/m�[��5��h��T�m-�~���S�U�w��-�����T.�Њ��p�*!7����#�>�����É�RM͔6��d�+�5���Vb9��ҊNqz�p�&vm{�fVJ嶲Ce�5�j��t��予�z+���kڴ�n���L��v�6�r]����z�����zk�)rC��,����iߙ�Ǹ���"�.�C���v�����B�����m��3f�G�1�MM�+��+1��1�;�l�d��q���+Κc�����6�[i��c8w�ˏ7E�lT�ۖ�n����ӴTƃ�<���{XvE��y���s|��er���� �ghN���ś3^����X�T�Qb��ֺűL<~~r6|ڊ��B�{�hU��e^jy�z��j��,
���D��㘳�Y}��1��+�[�yu��;,)77|������[l4��4.Z�X�!�6q��������3�j���3��rQ��{���^'UK��LLz�!P�.O�B/�Jɶqhlw�us5��rI��.�����Q:�=�W	��ZЦu���Qn2�Cu2�͓��c�ۋf�c���!��6�����[~K��"�t��˦3�|��\����:�Yi�{g��1�t`[�c�dk�✩�Y��&�/�Ie@�u펬�����X�z�10L�+g�ֳZN�t��fy������;����'գ'u���)ޠ�e��b�=�9�WDU,�Ф=Iu�t*�_^[�Bۖ��7���,��ۼqf��L�{����[���A߶sV1a�Y�{u��ut|�3o��ϧ
�)�TQ�]��7�6j/ic����#�wW�|��_ʃZ;)��˾I�]��;U��f8d�'����3I���=�^6���xn��#�xeM�8W��Q�O"a@��t'\��7Ycp	�C�-s��n�U�uQ����̼Ӂ���8)����������dao��F=��Ѯ�iC��Q�z3fz��V����L]=`=݁;�EG�Ţ��6q���^���v�p���+EEQLމ�����3a�����Ƃv�o<ڍyƽ���Vg*�3B����{�\������������:�ZШ��wޮy�# ��I��kw���9v�� z��岴�ߝ��i�Y�n�n9���z�D�����cov�����OW��1J�Q|�婄�ƶ�팇�(���;Sr�j�qM��w��M��^']D�3���H�Nb}��;,V��Y=z��jH5o^(M��7(�@j�s��M�O�/��{����C�Vh�J��	@�>9���K1d��ǽ��̽�i�	o��a�7,h�I�'lQ�<���E����ف������}�,nv�lSB���Z�R�Hހ%��I}ln摥w*g�"������j�vCd>�XYӑ��[a5BA�u�PB̾ߌ�7�tO�G	���y�,�Ҳ�Xv�j馷�sVA.�Ꮦ-��A�KH�<��$LSl�:�n�n�wVmwj�B6�f͵Ӧ��YaQ�\{e���ġDn �l�>!8woE߶�F�[IE3��X�T<�ۚs&<���6��׃qJ�$]ĝo9*��l���՛���F�˩i��ήFm��./g�<�.����i����ufPew#4I˺0�;�5�>洝��Kw���y�}��F�i*T�v#��wz�#��;}p sD i��X�k�ۛ\�=�kR9����zeلr��j�ΥܰQ�wH2Z��r㎏WN?q�Ԩ畇&���֩�2����[6/3y�}�qW[&��75fp�cJ��C�������u�v���+��$n@��[I�ҫ]�9C���;�v��i*�1�;�� ��4L�]d���)��Z��Z�l����(n��V:#ty09��R�XIR�5$Kʈ���%	ԡ�������xNfe��o�ҔMlo��csa��*]�%��P�eJy
�V9w<��3���r�����f�2��M�Ɋ[����A|���o��F*ɂ�f4j�����+Ʌ1G��BL�n1Z/߇�4�]Ee��1~x���r�=Kk1Xm��{�IRw�f��u)7R��`�������x�e٫�v�5�̃f�d�lx�V�|�}w��n�\;�l�VD�.0��0�<�Щ����;�x��"x���0I�u�������˧�cۘ/r�{���N:����>��b�j���:�8�^��-tf�G*�p�ܬ�3 ϱq��v3���\�7zf��u.D����*y%�t�v�A�Ԋ�ԷAmkW׬`:�Zy�X���\�6�8�b��îO~.K��_i�wq�T�������nԎ���ř�-�v�^`���[��f���k��1�)���hSy��|���*@�е���7H��Z��ۋ)�-Ё\\󽳐�\J��җ՘�(7����u��4���"��)�G�
Sz�仙��cnT�<nW�ZGe0�c�)�K;���e����w\��WL����׼�y.��Z_N�qKn-��G7���5�i�����i�J�TMU�P%��T�GS�*��l�)��gT=
�ݔC��i���Ǽ�Ǒ�8U���>��\��F�Q"�":�����(�쌥����c��B�+O�;�[�gM|y�1��j��B:��J�x-�p���hk�9�:ɫr���-F�P�Z��=�=-W:k�A`�]��LެA	S���G����YZ�-�|r�JU�E���
Yh�#F�m���+E
�(��J��m�h�[-J�pF.FX�F҈Ѣ%��P��jbW-UQ���
��iDeB�[iY[��
[V-J��b��b�h�2,�["%��%��ʭ�+-�e��Z�(#mJ��RڃD�(��m��h�"�Զ��"Q�����X(�Ԣ����iV��J�Q��ƈemQc[-)cV�J�R��e��X�R���(�ڋYUUDX�R�5���E�m���T*�rщiQJ�J�*6յD����bZUUmeAb5�U����"�6ܶA�-b	kT��V
�E��T�T��TZՌ*Х(թm-��9k`�!V8�W*�-���ڑ�[k-�PEe�UiDQ�ƭ����[a\s���ݽ��깚�{)[yw�кg��yX+�^��*p���q&����_�*�f�����9��lL�"���aO�ݼ��c�[ۖ�9��ך|����}��D`�߶���W걳/�Sn�A�ҷ%ĩ�+��;���O�o/z：�{gT�B�*��ljnW&'#�ؽ�ۓ�ei�F��^�VD:o"��V9�VVbl�=Uٕ}	M�Soj3ǜ�]쭗�Z��;�*�sk����������ڲv�2;�RS�6�V	݄��f�
k�6�q�l��������]�i�ɸ�j[>ژ��X�/%1B��'K�G}�	�W+6�{}&c��������\ڸTW����^'tв�GX[Yq��3��ܒ��f^�{��cYV.�ޡ{��7��A��6��4V�7'V���D8k�j�M͓�
�e��[e�ףy��XФ�h�t�\��=����۳'Y�Z��5�����*�t�;��Ol:s����͓m��Z�j@�V.g��GpYyz􀃎�-�=�T��9_����7��6�M1���B��8-�l%/��IO������ʸ�m��U_IC��x��S$���Y��$��2����q��]ݱQ��=u�����}� �]ˇu%gi�f��v�[y��o^�r���@����
�{�)��8����i;�?p�R��Y[�ͪ؛<�RW٥m�y)�>�?iQ0���]����D����:mL���q�M�܊o��+2�����^��t�R{�j[�ʷ�xA����� :�/�M��y~zm��nV^;m��gL������2qץå�=|�\-
i=hzwy�&}�o��e��$kȆy�;�2��E��+��疴)��T�a]h�^����k��5��|��6�p��޴�n���冤~�o�=U=x��F7�W={��5o4��[,�;m
��ɚ���[2��w������L�o�+n��_vǛ�qjb8��:F#=�p����n���1z��sY�������`�sz��B�jy�ۭ�t���y��/��"{E	)۹���e���4�T�+lG���<��Ԣ����"�����+}%�-����8v����VW;ʫl{@���*X��yy^ѻ�ݱ������n9�^�]{��b�f�g�E��'f*�tչA� ��m��������wR�x�V�·���5/��}u�W�sz��B*58Y��ל� 9�ʗu��ܥ���Y�a�h��t�u��q+�����
����A��/v<򰧍	יGbћʮa��X�l
�_%;���ɞ���>���;Wb[ñ�r�O�\�1�2�ǅl�q��~���Y�Du�1�á�rk��ކ/dO�JQ��|Z��'������l��m+�o�Ćg&�,Y*��%�v ݡU��tV�d�9%�����̙�7�5����%+�}±1�T�9'Nz*�O!W�����g_�vZ�p�u4t�SؽwZ��{^Jh�Õ=���d�z�!^�����-�彇q��)U[K!�ܬS�*�ĵ�õʃ�������Hu=<��	���$�+��I�N%N}d+'o��I�����c�1���eLI�����ݪ�0G�z�vkyP:��L�����'�w��c�=�Jɤ��I�ze�I�8�é��o�,8�l��8�|=�4zf8|�ܸ�om��'�mP<m��0������x�ڣ�&w+q��fˈ��=H�m��B�����m��c��LǏ�E�~>��HD��[�g�jN9P��kv�xb�l@\u�K,�غ'��:U�����d5mU�{\m>�-h7���u��u�i.������!P?!�o<a1��s�������i��{�ē�o�2La�C��B�m���d�Q�m���B({�B��s]q���kʹ�z��>��y��M�m�n���p��6��Og}�I4������O9;��&0�C���$�'���+&�XyhG�{�F��U����hZ����vr��6�{a�N}d=7�d�O����d0:����o|�hN��:��i������=I����,��zv=�캫����ݽ�V�Y$SO�s���T�eIP6�L�J0�d������:��i%~d5�8�ԟ;a�y�4�l�d�������s��O�G�+�7���j���ѩ�g� {޴;���*I�j�%I�VO2���d�������5���J�d5k'J�a�7��I6����N0�js��|��˭�bjg����E{�Y�]��CL�Þ~���u���}䘕$���Jɿ��I�M2u����i��N0�~��J���>��Qz'�u����?��i���+��蘜��2q���d8��7�AI������$�ןy%2N�7�,��`xe'6���~��'OP��'�<�xn�i?t3wM��;��moވ�{چ�v�+*�xu�T��0�'X�$�M2��o�AI�O��0���o�y&?2N�Ȥ��a�$�`�7nk�9͝�{�s9S��G�D#�d���i��1��.��$�!���PY&'��a�N%Bs�~Iğ2��� |ɦOf���I1߹����Ļ�l_��������_�z��Ї�i8Μ��M�<���x��I��&��/��a'�8���N����sT�'�8~�O�q�Z��,�4���/>q_㋽1%M�>���9�������c�+�
�B���{m�z�l�i����n2�<��M�B.=�GL�>�y�F��>��1����rY�5��?�dqo0�`˝C.��i��fM�**�X�|��[�_h��Y:����mb*6mF_Q[��Q��G��=�}�TM�0�'���O��=Or�2O���:��O��C�N �{���d��y��N!������~g�|ì�t�o]x�u2~��E3ײ�:~��h��{��=L�?2|���$��_��q'�>eB|���іq�|ʞ{C�,�'���'Y=?Rm'u�9��:�z��ΐo]g����a�h�yG�L�	:��~;�8�Ԛv����:���yϼ$���(m������!�<d�{��I�:��P�$��Xd�V��݇��٩�͞��Ǯ=B<�{����Ed��u�I��3'Rq���;� q'Ι9�'XN���$ĝH{-2�i��VP�N'�S&��s�/)ռ���e��Z�>�=�`�"LC�`y���6�ߨ~9����a�î�LI��2u&�0����I�O�w���I���}�LIԇ�ΡY6��������|���l�����ވ����>�=�'S�������C��2
d�'}����
���f������u&���'���N'�����C&����k�]�������b���"=�G��DVM����8�I:�$�I�����'�P�'_̇����I�>�CHa����$����p�gY?0��֜{����qT�U/�ޑ=��@�N���𘂄�n�!Y6��ɔ$�M��,':���RN3�I���h�a�R|�e!�	���sF��s�{W��������O̞�������l=y�	�<d��?x$��쒥a>�:²m+'�P8�L���q�I��ía8���I_������Z$�u��f�n)�=�{��B�=d���:�H�܂��� �ӝ���N�	ԟNg�$ĩ'��aY4�@��'4��)���f�9���+�<�G��l\�~��Ig�/v�I3��y��n�k��第�*��"����σ#ugN�u�#}u��ȫyq��I�O/��TS�N�]ܪ;]��8���81�p�c�%�;�%>�����Q���8�q�0:jF!Ԧ�ƽ��)F�C�l�gvriB�m�$��$�z��Y%J�S{Ì:�9�=��N �9�2~Af�� ��'�����$�N_�&%a:�ُ�!�"	X�́����rE��zm&�'|�4��yힿ$�C����βz��ﳬ��a����$�����8���s�2|���}�
O�yϲ�c���K�d�,*�y��R��*_vL|I4�vȤ��̰�i??'�(N2'��Oq�����'P�zΰ�B��[è,�����q+!�،�=�G�N�|�U?��f�ۮU/��i��;�^�1��[��1���6Ȥ������䟞�0�O�i�x�ԜI�&��N �ϼ$��Xk��`�����P$囃pX�Q�b��_�cޠVC�]���4�'���4ɶOC}�~�1�߻����I�{�"���OY�Y�I�T����	��>g�8����䏇��@7]_^�gLn��I��k;\��&�m��4�RO�~5�:�Ĭ���p�'Y4�'Ǽ�2i&��;�	4����&�I:���!�4��Vq�|�<`�@�t|�8&:�uS�sj�]��P���
C�N!�M�g�ϰ&�uM���	���'�&�w:�ԛt����'XI�9�	?0>��Ĭ�$�˓�FP���b<�׬>�ZѴ���D'�Vt������d�V��&�u��Y�>��I�=3�;�$��3�u���Ӑ8��I?s�'XI�O�#�ǽ����j�����ٮ���I��3�Hi:�*I�:ϼ��o��d�V��M��'��sY!Y8�����Y'X~�aԛx�~;�$C�#�a:kjV�_՟XNw��H�m:w��&0�!��T�Aa�-!�4���2��m'�(u�$�k2m+��8ɶN�!���
��{��B=���ߨuWb:6��V�7bks+Ss3������p�r64M���(��`I��m6�>a��Y�O�*]a�.���� <�oaM��m���Ҏ�����eI�%֩�4⇓3if�S�]f��ñՐվwiepƘ�9�2�Ym,t�����#���ػ��_�ֆ�����_�`�X�����=����k���I�����1	�:�I���6��:��d�I���g�'�P�&���@�M���~�v�ƭ����3O�z#G���O#ޑt}����d&��'������{�{䘂��ݜB�m+'�(a�M��A���{�}�{�{r�v��}�\e�j�UWֵ��!�=)�|=�{C�d0>a�9���O�m㿲N���I��w���{�?x
I�=���IPP�z��m+'�P8�L�|}��2���Zܯ�4�U�{�=���������$���֬��>v��<��N�N�2u�����&�Y�(N��'sو��y�yQ�<G���WUR醴9�w��%d�VN�'��d��zya4ɤ����&�������}N0��CG7���M��0�)Nw �ğ �ӝ��CL�]�p5�W)�����w������>d�I���XM�o$Y6�@�e'4������m����_�N!��`~N�z����Ē�������H�LX���=�d.��4�y���?]�
2m*�X~d������u'�s>�L�d��o$Y6�@�,8��O�Ɍ���x���I����N����z=� ���+k��f1�G��{����}�k����N�2u!�9��d�V��,4�����&2{�����u�E'���ì������8����h�����z�[`w�����ĳ�_}��}�f�|��t��a�����3Ӛ�Ԝed=�ܟ$�&���s�̚d��~�l�>��&�O[�R`��'�ǣ�=��|>�k�f~�٫�Z�|׹��s�°�	��q<d�'��!��A}��$��X{�a���|���N��+!���:��M:I���>@�OG���p�F{��!B=�<�S!�������_���^�io��5�J����A�-�K�s�h�f��t��)�>�Λ��c����nl��X���� ��*��nhz?yN�ƻ,�癋�b���<�s�^R�wE��RS�r6o$��R�&���~��&��;����^����_}�w��5߿k����6��?��:�m�<=������N��{?P>C��J���Bm�o)��zϹ��d�'ݧY:��h�;�}�p:���WѶ�z�7'�k�~��	������OX|�d>Ld�+6�i
��è)&k��A@�?Xm'8�=9������]���z������O����*7rk���+wu���s���5��<I�l�=�I��i�y�>𘓉e��VM��C,���'Z�4��La�n���N��<�a��d�T��B�q�����~���1�	���+�\�0{�C��}3#��'uj~~d�w�q��=���Laԇ��i+&�Xyi���g�.2M!������maěe`k�5��t=��J�����nZ�Ǽǽ�ǚ>�C���n�Ld��0�M�a?�V��Ogu��bI�{�{��l���B�m����d�zad�a�k_}�?,c�����#2��^e�Ϣ���}}I��C��8���Ձ�P��Ӷ:w�4�O>a�>�r��'���N!��{䘂��t��h,?{�!�_�u���v� ��{}��{���hu��i�{a�N}d=��2q'��s,�C������H���u=d�S��M�Ě9߼�u��˕��9��v��v�R��zD@���M2��(I�N�N2i�!ֲN&��$�̇��N u&����d0���N�z���y�q=d�=�{MS�4`�r�?v���'�"�}��Y'P�?d�*I��*M2�T�d��O�<��@�~C氛a��:��2Mk'J�a����'RM����ߵ���u~���~s�׽=d���r�C? ����d��~���u�/����IY7����N2i���������z��q���|��d�����.�)����X\�W��u�IbU���p��ɖ�4�b�3�;�x�GU���gq��D,MhA\6�5[�+L)R�to�_�ؼ��L=	��C�dl�]��dN�՗�<۹��s3��.�}��j�oml]�eY������~~�믹�z���f���J���ް�N�����Y8���s�2|����R~d�����$�ןy%2N��H�o��Rq�i=~O��8��s�[����u���߹���$�M$����HkW�������Y%O7�:�����8�L�~�p��L�w���&2{�����;�y"��y�~��<�6S7��ӿ{�{�v@�M?���!�C���d�R}���/��|�P����$����'�5���'i������&�߼�I�ָ���v���s�9�uZ�J�R��c���|}�#��E[0�N�Hx��O����:��>�i8��ԓ�8���N����~9�:�ĨOO���N2kT�����o�s麪�JR��${�=�﶐�{��9lǓ�	�zȤ��'���u�|��Ohu'�ݡ�'Y?2|�Y:��}�6��o,�x�=c���w�{��{����ޝ���ޞ�x�����:ɽR|{܁�&�i�;�xI��_��q'�>g�'��'Sܳ���T���Y'���N �z�i8�����k�nzy�k�ߛ��{���]	�'�:g0�z�m���d��	�9�8�Ԛv��l�@�O�����O���Y<a�r�~O8��Ld�C��� �L����|���f{������w��c&Ұ;9I��I�T��B�u����I:��3'Rq����9�>t����:�u=3���u!�4���=".$�#�C�b2�o�ر����O��kG�o��l��'|��x�4��8ɴ�ԛI�N}C��d�d�=�t�bO{̝I��'�r�|��w���I��Nw�$ĝHk]y��~9�x�73G��}��w�w�\�Y4�ö���:�+	��O���x�6��:ɷ�!�Zd�'P��HVN0����i&2s�u&�����w	8��og���y�r����CrJ�/5�Ӌc���
��#ޭ��{(E;3ysi������7M�0	2���b� �}9W`J�ِl�R8�v]v�H�[\k:msή��{iέ�>5��<�Lܿ��s��BK�HKiʽy��>Ƿ<Ϡp��?�� >��gy�et79߽=�!��c�" ���>��h,<���N��)&�q<��i�	�ze2u��zo08�ğ;C��0��:Ý�x�c&�g/�>9��5�|���{�n�M3�M��ߴ���'Ns�d�C��}�1	�ݜB�m+'�(I��g�	�N���m�'�{a��?2��8��O���o�������j�{���߽���C�'4��O~@�7��=d�_����z���d�C���*V�Ӭ+&ҲT$�&��ǖ��O?Xu�'s~���{������Ϲ��w5��{��
��d;5�:��M<a��0�ì��i��I����(x��9�!�>d��?x	Ԟ�g�$ĩ&�0��}@�d�&�;�}��6��5�eV���J���=����#��D^C+�������$�Xxoxq�Y'?rx��)y܂�>Ag��R|���W�G���d9���A�|1}����	֫���w��}�}��H�m���OY4�����	���ힿ$�C�����d���d�+O��Y%|�2u'R��AC��%a��'�<�k���}�߷����vz�c'N��$��o�vE&��e�XI��?yBq��>N�x��6���d�޳�&��=���D�x��{1����>�}[�U_m�;t��Z������/ϔ,mO �j��|O�r՞��T�|��N�����{3�3=�&�E��<�}�ߋ��f�R���r��}�Z����*Y~�f����m�+{V�M��;��3-u�>�������=�ۅ�<���c1ʗN�q�t�,:�SR5��w��T�Qc��U���6��k���g+��l�{����D�j7�X��\WG/�Vgq��{J�B�#lk��*Q�+v�)��%b�P1����q�n�BFZ�N�qS�b���J�9wF�4�e�\�ԨY���n5�|�Tv�R�w@
=W����OVd/\3�I4A㎮��n��/��U��< F����KE)ٷ�A��U��j�sOJauk%���E�$����`���Ve�S���r����̬8�����A�:j��tW+�]�@�S��IT"*j�}t�%�`���¸@�*h��^�!ee˗c�um���q.պ�k+KY���.��ew	%dGC�;�x�6�mCb/$ӛ `�m���r௶�B�m��֖����
�W�b�=Je۶�õ��u��<d��*�7zV�)T�CJ+��*lDfjN���oH4���Ki�[��c�F�M��A�4�\����k�=�[+��7gv������"�C_es��4Y$T~�ݍ�)t��g��7Y5�L��%Q僸�XH��j�S:421g�r\z�A���a����S���}�S�� EtW(uݘ�+��+�ݕ���b}O�Å%�:���׺�=�gM�nX؇JV�2�hך^S�t셮W�9/U��Gr��1�R�J�
���/�Ů�2��.���:�̏N���eI[dd��WQeu0�ũ#����q���wSs��I;���}��Q�	��.wp��ڔ��'������O�WZ�o,�>��@Q�0��s2�.���͋x/N��}l�Nwu ����V�4�1�Ԩ����k-,�K�:��F�i=;�&#Z&�`V,=jC�FƠv><��I�R�U)��c�F��|�f�Sy42�x-�4�	h�	�p	����Ki���n�!��q�/
�[]w��i��ڰ�F�;ݎ�Ƶ��YdP��bGW].}�.;A���SwA��wU�2���x�
8�X���ԗ��
3�X�+ "�7[A$vGs+up<��Њ�4��f9X��ݔ�!΂e��h;a����	\�G���㬫��H�3m.8�+�V^�R���ŵ}��I���:�*��i40X3-�bx�z�i��}�z�.QJ}��YZ�^��J�v,{LaKH[*���������1�'T7��>�Oo>nWbw���铅Ni�;n�$�xOm��2���[��;�g=��l��Y���������l�rT�6j��>�T� ���f�}/fb�t���\�vke��5$����ɖ+i{��d2�&(��}�}������g&�n�جu���-�9����{��s{;.�$��1��u��q���淦��FNDw6�EN���"i\��,Ѯ���zgR2��t���PG�0�YV�&��f��^���y2�+��i��H�J?jV��f���-Rֈ�ikYZ�ir��5PX-KKF�m���ԕ*,F�FZ�Vԭ*���-kiH�mQ����XZ���[�Z�R��*�²�ڡZ�U�ʩR�l�R�Z�6������FҖ�իb���ڕ�kR���JUUKh���Z�5Z�R�mQjֶ�JT��m֖��c-[QiB���2Ѫ��*�cK*�Ԫ�-jҕ�լ���ѵ�F#h6�YP�eJնU�,����*%mh�mR֭m-���PF((��
����R�����V��kD[IiE��Q�Fڨ�H��0kj**�eZ ()[F�D��EjX��Q)KIYP����e��KTJ�ZR�j��+
�h�,J�ʨԵ��V,e[k(�hV��ֈե�ch�DJ(�*���iV���x�����W=�`��j���`��L[�N�͈}�@Sc���\�Py�jط�>��ǻK�S5���S��D{��'��_d�'B6�c�^k��:U+���6��E7�~���4���Ν7ϵ,v��K�[��[�z)����
X�z
|���W����E��|Y��)�<��U\����]�U����_5kT���/����Pd�,8\�H�[+_N��k�X��ZN_���M
v��v�v!Z�@������^�ָK��c��n-�Hy�b��XA�jd��g�W�t���mN���U�7�H��Cz̙DX����f�l&=�d��jy�k�󞀻���jw)-��#�S8���H�,l��})�:��u)�|�mˉ�l)�y��SmXr�IV%K�S���.ٳ8��ԛ��y�sm�U�mb�+f�:����A�B�5��taܢ��3LI��E�����ot�ձ�Ϧ�^�u��SW���W}྽���wb����t%���Uܞ�;p���ܓ�+Q�op.8/�k��ޡc�I`w��!���j�
ֽ�<m�dY�z�Ѩ<Ҭm�ͮ7�����z�+�'R��1;�q�Z�Ak�Ήb���5�r4���r��c�O������ވ[��;��g)�Բ�Uߢ=�z=7ć`t����k�����F.1�_�U�sU]�I{������M�!1vB��J���յ�\�`���ñ�0py^������A�]�ټ:�s�-{�{�:�k�z�/K�>\�������<͔WN�er�v�Ź��^쮪��|��;�4U�C:+}����fZ��:^�
fѽg-����K�e���M'\Te�`�-�Uw��m�kEl�7����^OSټp���Ĭͭ3xrz����u���HW��^)�*��T:�9�Q���9V��>|����j��gq�T'{ us��C��עz��̋�f#�PB�v��|��Y��^.ˡ�|�a:�\�Z�Y1915|�2^lcʺJ���~Z��i���+|=����W����H�"�]Mo�r���t��n���Qfu�:�aT��?{H�\�U[B�K��U_�[V�66���oֆ���g�Px**+ -���ңB��MJ��8�E�#�ھN�o3��@�HO�VZ>���h��܅B�UΘ�������FX�ч3QXf��\�F�<�0�n��B�s�=-��ʌ�y]tWB�����z=�fyV������v���+��וR�ȅ:�>Y��n���9�6qF�$q8^��U�%7�M�1>�8L�F�S
�fF��q۞��!/�Ǟ{h'�w��sLb~�Շrx��Y�5қx]�fy�q��0k���n9Z��=�3�3�C��p�:�]�jWO��\�Og��p�Ļz�7�כ�v�_���,��=���ϴk���vL�ۇ���Wr�|�aS�M�"<����U��umw�;?OS^��F�SӢ�~���
����j�s�n�-ˋ���:�Ǖ��ۯb���^,H��"C��/�;%��WR;���[��Ί���ޗ��u��z.;S���������N'�-��L)V��|�-<-܁
��KlΨY'��6q;Uy�!�{������fb�N������²po'LUM���x쀤�tG��`8�t�я���)��*����ȍ|F����rM�����M�M�s�N��.K)Q��V�:�,h��!��hqjlJ��Y�%
K�&B�p}ox��X|�EfZG� ��
�_n�p��b}�k����꯾�'�M�$G�%������j�4����*�!p��r��ቚ�G�e�v634�K�n�T�u�Z�+��4��B-e���i�P]�V���,i��c�u�Wk�U��^+��5�B�OKO��ó�Y��Źַiu�+[Xn��֏aL!��`r茙4z���y�o8o�G�8��:}:���o۪�5���}��M�)��|f�Y]*���)gb�`*ˑ"�S�:�1��u<�;s/ͻ��_o��&k#����Yw%ѹ��	i쵝������ӽP��iNҧ.�*o ��8I[3k9�7��9!���旹]�T�2��y,�9�T� �t�����,�;؝�u5p�U�U/�;}�������_�3���	�sjÕ�,��q���8�پvo����9�a�h�����	_'n�ٌ�=ɨ��`އb*����F.�>Z�q;t3�@�������b=n�F�c��Kd�CoKN��uv�7y�k�R��1�Ǜ'V�� �Jea9�]�v��57�k��;���x�����ʗ�v�g���ԈR�,x)��m$�.w]��\���=ک��{�����}�[���R~�nw1��k�+��qv�3rg�`��?tk��Y��)T��8׏E��Zsܰ��VBJh������)�z�:����y�+f\^ȧ�rRڏ�g�%�M�����6Q[}~�8,GX����n��w���>��꽋j&�ޝ��2�]y�.�Y��=$��j�C�G2�֍�r~�[Н��*�����g=�'eI�����W��;k���x�ow^ug��7Q'�.ө���B���>w�[ˇ�f���Žŧ��8Nq-~��a���@k�qԸdE�YkB���0r:�f�؝�kB[&����utF/���^��N�=PW	��$A���ւ���S��Q��U����c��[sm
|X���!�A�GC����h�cz#R-9�7'��ͻ������0#Ć���������}G�{W��{b~{c��/��u�70��1�իf��-J0����נ�{�g��d�>۫E��KU� ���&B�T;{�]��븼�<wO����7]�[��l�0T��}8�8z���nѭ굷�:�M���˞B�-��Ц���{_z=�{������3�Ta|3�%��,�S��}{��u[�L�,��@��M�JҺ�[���Z8?�Onz�:ᙺ��)������n������l��֫r9�v1�,SҶ�;"-��A�.��J�X�svdMݸ��S�ы1�����s�&����E۪�@-�����]�WUܧv���A<m��;/��}���;��]K���*㳧-���n���|���z������q��˙��Mw�W,��"k��m��w�z��v1wP/�/�sԶ������\���\�b6���kr��|3�,�ɹ�(V�v�9mu�Q^��Z�e�օz�{�K7��l�X�QWI}��ݸ$ͪA����)�	�;�9ˊ�ȅ�m��D��S$�������Y��;q�]v��[��Ov���EcqQ|����4MLh�����ۜw��2,��xg+k�	�F�Od���Vuvl�q��؁}~ WV!ľIU��}��kjoJ"�y7�޻��'*.��mt��/evՑ�	ގbM9�]� �e�2�a��پK�����m-�9��]w^~_|>  6��������ż�U7�r��;��*;"��L���L�cr�q����:c��h�OB��|�e��R�Y*��	 'Mާn�-�l�&��\-
n=V$�3���qm�6ӳŃ�f��6
��v���7���d��{|�]��og[�Ӓl��t�v�����pŨK�X��0��萵юuë#ѧ���VE��{G%Z��~mڰ�`i�Z��=��8[�'��>+f����v����� �R�8�[��K��s��w&���1�b��%����������.��%m|:�d�Z;�����q�z�tc����c�>�:�sQ+���7/����j��o{����ޅt\�:��.�F��V|~�P��;v���'����R)��\��we�X��O&��Ţ�lߣ<<�}){ذ"���f�(����#*�r���ھ��gt�K��]�س~��+" ۹=X��ΧN��!�:�W��S��1� �͗�8,�ݖ�@MTƸ=���*���Ψ����W2�^|��uLX���잉�D����z#�f����T�����Gu�Fܮ�d��Gn:�pecA;X
=Z���G�;��'�����y0�ҎHZ�Vz�[��QS��S��9y,R�׍S����r����9ͩ���3l�s�)�������g'[��-{���}���ξ�䛖��9ًlu=~���PK��	���w�KnK�����^Z�D����O{)�������6,�b�&�~됟gF�9뒡�Z�|�腁�O���=
�6�.:qI����I�7:�+��*"z*��Fhc��?�v�9���~t��~z�3)����kO�u��(���NX�N�\��}�4�5�h�]��ǄZ^����LS.�s�v9�;��8X���!�j0���Ry�]J���Ib9<��e���74��F�x�����"����yˮ��}|�\t���UǸ��yJ�M���V���^�zy�9���ʳ��k:��m�_>Ի�pt�AQC��J8��S1"
�HWi�R���(�����נQ��:V���|����V����^E�z�E*Pf��":o;�W}[l^$������=����Ujގ߸��#�w�u�)�T幸U��c���0�n6�n�����z�K���ɍ��Y
m�f^	XC��)��G��Z�z��[�G5ܳR����ݗX��ڨ�@w6�9Q^NE'�����4b@���Dkuٙ!��CF���;u��J�7sޫ���DL~�r���W>;��(%�v#� ݴ�=����
�+�޼���S�#��W���-�a�޼듗]�!��vE��i7΀��;ۉ�N�S���"{�r�'@<Hw����s/2l��s�z�؀-B�t��"�_�1����C�-:�^F�B�Bxa![���m���^������	gz�+u��u;���D�n��4�thxp`�%�(����ђWw���z�*/�J�D��L�������T�(NV�6V���׻N1���F��Z��V�p��E�y����b�S$b-���1
s��*������۬��t��Ѯ�YR1�nF��Q.�0C*1F聠�mvL�(�z����%�\�L���0�-*}���K��}`�L�
����n��`�\1s���*}�tUv�R^X#���p���4�/�������y�573��izN�ʃ���{�H��ވ�z=��FV�5�JS�0���,�F.	�#�����w��Z�N"��^�_�/B4bќ��9e�\	y䜎��Ýv��Vl�kjB�4b�	�	2%��+��*[K��hᘐmǏg�V��he����*-��s��5�~�,�x���J#`�Y �d�i���[��?�}�+�/�?�U,,���9ˢ�eqx;0n,sU��ͪC�&�����mQ
�w5}�6.E� p��4���a�q��e�:c��;.�!y�F_�XC�Uq���/��ozI�h�m"�Q3׷|]�=@�B飂����M�	@uLv�7K+;��)�r7�#��/x�\�?B������4��].Z<�7����Y��U�2����p�	���GtS}f���a���C�}�=��%qں����b��U�ܾ���s�m���1OT�.;oY�aQP)8���s�4:4xĕ���E��R��j�9�i+L��jS�ai{�̌z�=߲�
ue��A��<��E�xc�)v��Tl�f�έ����A�C�j��FW�r����No@4[/�-gb]t^��EkJb�0w;a�]�O%bRػ8B���в�4M��j��;ܹ�N68�۫��\5��Y�3��w�L<2c�B�ˮŀ��� �ݙF��O�˼O@'����M6;�FE'�<����Vm�U.Rz�Ѩ	�`���a�H�Ѱ���]*�M9��YU�g`��F�Mulo��UE[S��M"}�&���~�yT����D����N��ي�a�iw^�6�1�w�R��t���x$�ҵ ���Y��mMy
	���P����Iu��Sy�Vq�S���L�&�y{<יv�.)J��jws�Y[լ:��r�ٍ\�gή�ў�b �K;��NC�fS�A�5S��}�����K�M:;�k�7,�虡�뺙��ǣ��m!xo��>�㋦���N���^l�9���9O��'��DN� �����Ia;�H�/��<B���'����!xѕL�(>2/\��렅���{������̇K�U��5��(��t�S�%����Vu��N����Ҟ�[+�s�p�x�X�@�J���$�i�Ӗ�ɠ��u7fiM|&��'A7&6���}3�`Cl3�� ^�?owD���@Xk���Ũ���[3�y]��tlNͱ�J6�vR���m�46��'�Y�'}��Oio(2�wO�ǘm�=A���
j�;������Su��c���>�h.���V/Vҳ��H�׻]���:��~
�0�r�{�y:�(h��|�>ۙ+����
�d�u#ܮ�wogw^�;)��Qo�>�y��q�|d�[�w�`�Y�tm��:v��whr����#P��T�;��Uݪ���嘴:Sm͍&pl��ɕp�'���e�5k\NvԦ�O�{Zw�����X�m�voa��G��B�^���,�^^5OlΔ(�*M���ȡ��;,����A����U��F�0��&��ծ���.e#@^m�/1��1�(���`��f�:DnN��Ȉ\�3���� }.�������uc�v�gkvY��rħR�������aL�S����k��J/�����N��7b�M]cx�����/�T�w�(Ngv+đQΊG�؊�rR�ùqkI�~W������C��WZo4�k:���6�Ҝq-7:	%�]���l��N�v�3���.���;""������ք`��tajI*����pd�ڸi�J�$=�o���֔���A\���_P}��J{�j��唲Hy(<�Ǹ�y��J]Ą���q/�C�ui�Epɳ��Q9��T�a�gciX.��Eu6��6��t )V�6u�q̾���l�r�`ޜ�7��h{�x�L*q��Nv�5�gn¢��R��0��K���sN�n;K#����4���[��ڇ�b��Sʓ�����^�QF�J��
6��kE"Ԫ��h""��Aj(����Z+[eV�EJ��h�PKJ��ԭ��T�(��хjU�X��Z%kYR��-(����� [+Z��kZ�ʍ��+QV+[*V�Z�kU�J�%l����YDj
��Z%V�H��5Q[e`�[e��R��#mdb��(TmP�KZ(�ȱ���R�VҖ�F,Z�
��V-�+cj5U�Ym�cj�V�Q�RҠ�Im+�H��,�b)YQ�m�V
�EH҂�hڠ�[b�(��-iD�e[jUU
��kDjTJ��X
,Z��+��Z�R�J%B�6�V-Z����Ƞ(�V-V
�`��-[X%JԌEѡR�
��ڊ�)�PZ°�R�U�*T�խ+bF�PX@��V���X�BU_�7����o�kY�<��x�z�#�'t�]m�aya{��!�(�	b�y`���@�
R�3�J�"��Ү��5�=�����58��ö��U�{U��l��N��q1{��7�Y�q�5�nX2ٍkh{��yq��zrѾF0;ۦ/L�62t6E�m`wΨFZ�h���ї���%�O{N���}���kL�Ӟc7�����	�f�JB��P76S&�ip�݌�����!�7���D��S];�r��yq�^q��`Q�B=CI<dPy�/k�ũF���0�k=�K�s�;�낹g��D/��-=���OrC℡�面�L�����8�s��10��.��8���[d1P��ũu��>����A��4Ş��W�c���z:��K7�[�N��dF�L��6V��Q�Z�(�3��9�����72����\�׎��{{�,��P0g��GG���`�jT�S�=y�xW]7+�S��Y�
�*�����W˭�'S�ऍ����$�137�^TK�)��:�<����S���ޗ�!l�.n1�p[��M�g:z���C�v�@�|i�t���P�^.K����}khR3�0(W,�Ǜ���;ߤ�ܪr��F��D���,#;�ò��9+S�q0F�pP[�\�45�c,6*�gd�}6��c����9Lq�������Ɉk�]H�-R�S]�@�ᛀS�X6w]Bv���>7{�d�PE��7��r���j�'�^��g��
vΌ�,V�:?�w �� {�t����iw�P���7��
����)-ƞ*W�kD�/T�Ey��1ЦV����~sm:����\���[G�y�}�u��cy-K����gn�Wk�c	���{��A:�S��ŧ@h�n�e-�]^�KbWyٔ�s�o9�#H�*O��;�X��g�݈���@����ү�a����E��U�|���'��ے�m�C�x�6vj������V�����pX���>����yf	�a>}�'�}\�7�9���7����a^b�������٠�vl!�Ĭ� 9
LQ�mt��~��=^��"U/=�¯v;�y�sϳkye��=�ã��Y[7z��uGɚ��]��:/H���⺐��gy��n���S��s�r(4�_Vc��=lPA03�Z�6�Mkw�5mЎ��ŕśU��N���t��h���n���uaq2o]��#��1�ڭ�n�aq3:�=](Vx$���2�ÿ"�i��P�9�د!���dz�m�\�������,k��ӡ�r�������z�9�o�H2�f'�:Tz4U��5���)��h�}-��E��f�{x!�FJq�b]���G4LJ�uyR=	rP�z�t=���5�O�X�o}n���R!�dw��Edr�rz1(��Dz=��a^�����G������&x)s!lL�H�b�XV�z�쉷0�O�\���efG'dU�r��	ڬv|���irL	=,��lEJ���K���\�~[D,���ٗ��mgB��}/e^	<����BZ�E�<�X0�|���(Pr�٣��L�^w5?!�,�E��N�7_��W��r9vo��p�l ���+&Ô�4�YNO�Mz�i�WZ"�ܼo@�]��_��cS3��3��Vz��9�E1pG2x���#�t]fvޥL�{F��<��㳣C�rc�XThl�7�C�n�)��k����[5�[K\��r��$�$d>�yh��K���9��	�g2J��=�D�y���Et~R���#�.��{���fH����Z��x�
�e��*�e���^o@�-��W&.Ս;v��]������ �S�Z-1Of:�%𭲪Wz�Ҟ�����tG�h��ؚr��HL]�۰��w��<yMK>}d��fࣀ9�p'���@���4�ﶯN��t��Sf��m���p%��$��.�i_ɭ�oe��V��:;�[r���A�b@�^�{�z�ܝ�c�j:�K=��72Ժԋ����6�L�"O�Ҳ��� ��7��%56�U&�iRLN�p;\p�+}hs�:bK�'�k���-Z�5G����־�={������"��]eF3~	��K]"o����؉cG
�d�{Kɝ�?L���Yy�[�d�^�o>�F����y�l"+�X���aL�m�ct��ѡ��r�0�(M\{�ٳy�2{�X6���g .��x���S��t��\��!�l�#ޥ��}*J�����պ�g|�&	B�R���SV�,��F�ԉ`o�slN�9S���ū��TK �Z��S�W�q���.5�B�V���Ug�~���J&�a�͠�Ƞ�,G�*H��Aԃ�Vl����+�4b���	,�I'}v�^|z=��̃�ז�cI�i�=�a����ek�P�ytYq�lN��T,�u���b��=���ƚ-!�����tSV���`9���GS��#coaS��P�Ug黾��\���ª�>������t�ک��z�=o�*�ܺ���#�ͫ�@��s�E�͵۫^+�]���l���ĵ壜��5ڠ95��zP{Ӑ�)����Rx���,����L�������҂���՘�}���!���k,i��z[����Ps��E��m;�,��YW�]8��߲��a3�R���������lT˫�}�9m<�S�6�ǡǥk�@�v�����ȶ5��H�g��W�qvΓ�E_p+�z"=��Ă]R�
�@�\�j&�I���<MD����T�a�(l!V�]����5��������ϳ�P�����J�.mÿb���!�ts:�o�^���ͭ͡^��������kd{����ʈ�P�;'��gб�+�0צ���<6���S};|.�ɼO1��t�KV�4��1��OF�K]��CO:�ι�ȿM
S�0���y�λ7sz�����W��3�Uǟ�[k��i��=�]�q�gI�ph79�k���Ë��oc�ٗ!����Wb/gڔ;׳H�:"rl7�e����ӌ��(���S�ō{x.�o-�Ǐ��x(�,�Xڳ��<*ʦ���:���w��<|#�Dx5t�u�CFU���:�\؄��"��������%�O�8�AJ!+z�S8���Jfu�6��g8as�Q��c����i���c�߲��x.),g��Z#ܾO8%�_^y�g{%����2ҬO�)��,_.!K�E�>��C�A�������g�t]�Rob_Vv�0:�l:��eD�ܻAV�w�٤Ź5������Ȍ֋pX<���r��ћ�U��[��aE/��3���x�Z�ooT���V�J�=�^�shR���t��9Maeh��W�������J
������F̮R�{��}�}�+�hΧ��m���L�qS"DL��.S�jQ1�<�''iA�÷��{2�A)���j},e���D�ꈴ���ؐ,��vfU�_�Թ�[�3�3���v[r��e֒�ww���N[|�[+WԈ��̠m���R��(T=yQ.�����u۲�M�/f�x���w+9�+&��W*��a��i_Ԧ��P�]���qƖ���&������3�,�<�5�k�~
]��ZE��6�e�� ��'�B�é��i>�=��<:<�H���V�cx��)(��PE.�f;=U.)����sm:���8d�GY܋v]�F_D({Z�ss��ǹ�o��5
�=���pI���4�ځp��v.�4W��,M���N�;�f�%{fε E�c��zOD�~���g�۱W�g@�]��f��tI,Vp��D�ײR�����r/�p.��P\���9.��٤E�����.�oJ��.*�W�R�@].9�N��y�/��}VXc�R��/�h���ԓ�'E������`�;'wwXe��Ʌ���)4Y-����+��S����ʾ�ƕßa�@lCDg!��y9��u4�;�Ա��,���f�4�j�ϳ
�:L� �I�G�M����0�Wj�Y�3o�3��C@O��T�*Oz䮮,�}�W�}���'5�s�d��f��g���^�w��R�ON�Zie��j]F��� )�2{k����w-����BG��++���g,+��1��[aW�l��Pi��1��'n{v��:gi�zqwU�"`�((F�_��0�_t5�N�.V|P�~�l{n%e�Q�]=29��o��;G��Qq2��S�&+��+�x$���C/�;E�ӑ���T��^#�u��t�S��9U�'I�1y1��V�^Hv%�$?��u�]���픟p������o��o�k�6�}��k�I������O$�%�s�L�*J�eAr�]�Y0U��V�	�k:��ZFweh�վY�6!�*4�*G\>��~�0|SW`�A̧JG�X���DF�j	e\�a$\)�CV��p�'��_��xoW�S�*<�Q�H|{6󻂓��~��ly+9��鎯Z���K�9����-Gm]1A�Ȧ,<��Ⱥvݹ��[ʶ��P�&�G�.x��І�U��g���܊9	�=%��ςʼ|�.��z�f�~1�!�_xR)�]�~=��}WլtX��	K��$˓z�n3v@�1۱���F�aSP;�Nn��Aۺz�.Ս���JO��:��W�:�;���0�?y��Kh.9�ǒ{ݖ6�%���B�?z=興X����<�z?y[D��"6̥�E&�e��坛�I=�aC�P3wl�R�mnU����|\�
ގ�F��w!�$���z˥����K�e��f�ȃV���xhԏw��.Iɤ�&���e?���P��@ʄ�&����L<��j^u��맯+x/R�&��T�N��NO�:׹�u�Oz\>�!��%�:3����Әf�̴�@�K˳��Aiŝ�n�L��!�vq�/�z?`Z�x����cG
�9�Ecͺ��r�l�Wb�-����N̼�}�뀠�w�Ġ��ho��xz%n��;�[\:uB[ra͊��{��A�1����d��w��
������f�Lu�tS�X�ʧ�:}댘�˞j��s�X3�S�%|+�(_��r끲�et�H�[%D=�!7W]Z"6
>���5ff�
���3]��!ُ��P�!�y}F�F�/h�pm��k������#^y�ym+!<���B�ֆ>��ڐ��C;�f�$�'�D8�W����܊Y9����z�U���m�[t$2�����0fK�K��~
n��k���KkP�=y�+\�-r�ӝu*9;�ڼNc������!�'��䷢���zT)Ս�}S�J<��sSO��*�M�Y�Ƿ�~�ꯪ���~��N��g�*�5����b��+�������B���eǊɜ�Gs��엙J^����]�7a�� ��Z�BX�[e�Wq�#p�)���GS����sy��������ް���9�U� 	{PP��F�W�W��K�w���lK��^GϢ�(��߽St�ͨ��N�P���rF%��̼����P&U5��u���U�;~<�����Mg%Gy�w�kAɕ�r�C��I�Bx���OWT�a�(o����0]u:���*n�����N��Xx�DN�¦��.<v�U��b6;��t�ON�_��ɞ��FL-/r����ԽPN�;Lȸ��^N%i7΀ڂ��a��,����XN�v��
�y��'9���neO��Zn;��È���X���]���p!�㝁���\�˨qܧ7�_^M���j����E��xvl�+&X������mg�́vGır�&��V�ii���>w����ˈ���^D%f��\��K+��ǥd|LO���̅[X9�1��������f�2	]<�-q2;Fը�hǎP�pI�R/m.���˔�{P����Q�h`�ey^d���L�--��c&۸��,��|T R<{����Z�0S���w���8QR&�P���΄wv���Z����X�G�y�ʚ����[6�Ͻ�z"=p���ƺR�����;�:�f���1�����_�A)
����mNJvi$m�ǳ���s�q����c�Xact�NŹavz��h�y��W�����A��*RJ�u���WͪWYiܜ�!)A�ҩ�c��zVQn�]���!�(Js;E�]�ӹ���x��1��40��-*yo�l�+Ⱦ,\B�\�G�	�m����ļ4����f�*'��{V�V�'��c~���Ȏ��\�*��l�m.�,98���a����SM���燺��û2��ԌP�H{FK�P�B\�e`�o�oX�]�B�T�vR�j�x�˹�.�C�"C����Ŧ ��ʉu�2<l:�<�dɌ��e�y��$�t�^�W-r�{�r"0D�#�g��t{�����kn���)��r��;X���ܷ��ν�!�h��R���P�"�]1��;�p��`
[�tH�����F�^�V�>�n?K�t��d��ۖ�N3�|q8�a��:���)�D?�
O"-�og��qok��^$��=�m�E�K��8��4s�ήy7&�:�R�!��mSY�Yj�Z�hf�Ys�hm]`�6̧D����39��8�Î�C�t�O�1�k����M
�Y �v(
�G�g4;���ϩ��^j	��If��0׃�X7z�K���z.�3tJ-�O�0��9W%��\ݖ�yGSU�q=�#p�%��ݔFS櫦f�0�Λ��R��r�WHm]f�w0�ץz6��қ��X��84K�z��}%�I�rz�w�*zJ!�I$��T{dZ�53����o)����̣|���lήvo%�u���4�Џ0�VI��x�Ѳ6 ��\6��]�Tź'E�G5Y�|M.#�1P�Z'�5zA���~:���w/NukWn-˷)�廭�h�o�mCnEa���I��х��o�1;t���|�,�<��m�p��W%֡�v�>b��O&���Y�9s]P�'}�)��'BgV>L�]jv�.R��Z��}�h2'+`;�^��d�i�������jSpuZ�2U��4����giC���C��x@	U�-��#��\�#���C��u���Q���_F
�[t�^�*���zWH�l,P�s�Jڿ���O�,��p���I0k����Yr�և:�2����ոZ����*l���^M����:Ofuf��>Q=h���z&����8�[JݛCgB󍱳T�O���ATʻ�����.�4Sܟ|���k��q�n�S{�u9���="}���I�xKwwGk��P�xaݒj��9r�k�J�k�uץߤ�Y��C��<ÁǓ��"̾����q 7.����-�|,�i杁f�r��dW OsQ�r͜�����}�ۻ]z�3}�R��Ns��<��!W����`w[R���}o��T���3N�زh�\�d�K����#{NZ�PX]�f���P��{l��wZ����e���KBcC(���ե\Ͷ���>vᲰ���u�� 	�مm3��&[����6�j+�.G�Q>�R�ĵtv�9�  ��i���o��S�y0Q��IZCԱLj͖���`�.WTO�8�N4)Jђ��gu����-��J��*"t���,jR3�p��
�@���wH�^d����:���:d�7���^괦����'N��f�Ӧ�H�ܫd��A�J��wv+(�{{;K�8C/�tu+�(��P�eLe�yv �!��|��7N^���J�^�I�s#����
�;�q�+���e1��긷��6Ԙ�f�樳���{�q9t��mV.s�����9�\�,�ۉ��4u㣢�o�9[�^�$�eC�ͥj⌡cQ���t�/���s Ro``[u,J���`�Z������z�Tup�*��uj�X�%�y�}=U��GE�mT{��+{�ʝ1�wf5c]=�+Ύ(�vƗ��臮f�I�h��R�[Z�
[J")hT�Pm�FX�m���PZRщKXVRձ��-
��[b�m,V
�[URU-+iZ�-)jR� ,ʖ* ��J�J"Z����aUY�lV���(��#iQR�Y5*T,E`��)QEKV�ҋYb�����F5+-�hU���`VU�*UVŊ�eb�QE����T�m��EQ�ETXԠ�-mB�j"�T��,�����eE�l����eeZ�mRYh[J(*��lV֖4Z�ij�V�AV�*Tj6؅V�EIU�QA�dX�Z�4Dkb�F���ѭ-U�F�c���EX5PE*հX�Z�kҰU�R��(֪(�U+J��Z�#m*4�)Z�DQQ���Z���U
[F�mѪ�%iZ�Ң*T-��J%��U���,��b%�F[X�Z����U%-��*ZRР�)DTE��`��H�����J�(��PU�(�VTPU�Th[eQ�b**�Z���Z�l�h�H���*1�DYU���*"��|M�>�`�t6�it���(en�z�c��;p�����3sKݣΘi�נL5a6��N�	������ ������ވ�DfK�i���Z#��CUO�,ue��å�v�$�%,A����ET�m۹n�6e�gU��~�[�ؐw���P�:�IA���,���c��KӅ������{D�N�M�Q'��q�uR3Ў��H�#�̈�@�K��v�"�k�[�.g�]�ջ���	~n�䲖���x�s�q7�nt��&��cD�_T*����e����@����l�i�u��V�L�����e��a~jtu�=Y9ꚊY#��]F��hĠ�5���+�ۧuc��]& @+[�j\������E<2�W��c��p?5xv�U��d�O�����i�JK�AB���p��1/��N��.��7�ݱ�E�5�3�YF�M_n=xV��M�L�o�3�_����g�@ߖ�f�|a�.��f���Z��ת�d�g�[B5�8_X\�&��-Lt�V��͎'�H��]fv":UP�
��ܯb��L��Λ�Pu�����ڿ�aC�"'�&���N�Q�e)J���uԖM�h�FW&Z;r��y2�.��"���k��{U�����>ȯ����|�\d���V��T�w���o\Z2Y����谂z��ըD�o	���k+F�ɵ.�������8�N�Vv�,���Osx��x������8�;��������*��w�t�T�W�QV��H�V�f�oP���Q{�2��0I����]0̱t�S�j{2�����a�.�ծk���r.�xo<�]��l���.|�u�[ w.�sۯ9���Lk6���}[���1'5�B�f/KTg]�s��EaO?Z�g�o�پ�}&iH�%�U2:��!��6%�5�CB�rc�Y�F�nE�⡶2]�9a~}�|�?GՑZ.�I5�H�7�s�&�2�	z.Yٱ����9�g��v�g?b,N�=4�����H��F��;RK�a��<3fP��U����G\̢Y~|��������6�a�艜$�D����^Bt�W�+�ya)���RG�]
t3j���k*c��q�;~�,h5��p���Y���3�wYKŚ�?Na��2���SE�]�s��%�r�תcu�����աp�����싉w1w�p
����o��;��p��E���������甠���W��O �(<Ŝ����,j�����(9��i�[ăA5���_`�cn��*ؽ%B��3F�-Um+�F��n끜����nv�v�wف�w_K�3��������з��f��s}\/1���7W�َC�wl�|�p�n��%4#�5>#.<���}�R�Cy��(�1�ɨj������G��v�O;��+���������r���0=^�px��f:�bK�Xg��T!1d��3�� �M^��e�\�Ӈ"��R��]L�*B�NH�.�9�İ�5n�f�+�{0C�Z�yof1�8��S2�4<l�J]*�����{��rg�;kc�i;g=� �g�KC=}+�C̮�����VQ�a3L	o�T�Ĩ�^����3;�<.�rCO�����-��s���\>̢��Y4_����}��ߜ�A�cE1���0�]v%"���aǭ�:������|�a�=���ӻ�*Kou<8��P��G�B�{x��(ElЄoey�q��R��)��J�I���ŝ�5ܵ5�x	���`��0��5�s�U�1Փ )��'C~sW-��b�f�;H�lQ�	��1�LpA�����T;���1�'Euo�iOjOz�s��ZhuEC+�K���ɤ��h�ValJ���8T�Kf���6D�މ�5%q�Vw]-���=��{x �@�C����^>�̢ؖ��b�h�.�>uqu�@K�٦�{xN���+XElj��[�;+�ԓ�v,��]q��ѻ����{�YٛU�� 6�����sk�V�セ"�V�)�{o���R�ȹߢ=與��oq�btpH��1q�:"�u\�I���	ĭ&��P]�Z�6a���M��*�)�Ϸ���u(���XFz�o��c"̈a7����ہl�CM�4-5w��
��F��w�{1H~`H�;���U�]�%=/�F?�k<́c��'�T�3/-mJ��e�+۷���LZ�`���ƻ��.>c'Cd\V�+( ��(��,ҬYiڻ��uw�v"���9�F���C��xE#�g������"�i��{M�w�kl��w��%�lC���Ȧ�`r��l)�3��g(�!����W6���w�>yَ�;�G<��Je��:��|XE�X�=�Z{}n�]/.G��t\$��e$��b����ύ��Ui+��%�����6"����O��6���B�w<L��n�S�uJ��L�X*���uD4�+���y`�J,��g'xy1ԯSZ'{b��U����+m�D�R���P�Hz��Jf:�W�U'���pw�d�n��<3Ĝ��7X�q��L��:�"�����t�.z]��EV���
�F��D�
���Ȓ(	[�k�w�dֳ�;�\�~n���SZ\J����Ǭr��p����Ǒ���RW]�'�mл��t1�m`'��j����j`]�q�]��#�����>����v����fZ��w@�h%�.
b�v�;�sۄ�M�͞�VOOoE�Y�}���D���ޫ��8�y�Z�KDЃ�X<ND���;�D�.t�9m�M,�դ�Ä��P�W��֎�
]��XG5�y^w �>�-��[6��9K��Ǌd��[���!��y��'�p��넄��	@uO�Bq46-�1������ޭq�4�ۻ��杳�S�����[>����Y�(����o=���CMԲ��7�� ��*^��!������c�G-�>�@Tp�m�2_��V#<�b$�A@�>�5x(�0zz�����&�s��9�Gחr.�l�}�����\U��^���'�g>��^�=>v{j/{И�%�^�!�ͨ��"���s��x�'�^��ji��.X���V��ʾm�g���*��-�VR㥊�D[Ɍ�ڝ�Ǝ�;i���
l�O3�٫�G�ۏ���{�BxP
%����k}�R�o���x�1��X7K[:�z�wn�ƸA�RO䲘�#��x���=�\�P��뤎J{N�؃�!yys�y�Ss8z
놊�{��|�m�VT�"�Q�Lש�k����}�p.�؊�Odв��)��u���T�^f��1�;�)���.p��UnBF��:��{����R��o����D�Qd��も�8z�;���WF�j.�~h���vH��ۆ���7��yk�Yx%g"��J��>Ih���z� p����F!�Di�s�mS%x�Iy�&����"C~�@�v��� ��~ltK�Hu|���F�8/n�]��4��9ی�E�.Ց6�)�|'��O* ���O$��	=]��33먏zV	�i�-UʌN��s��0�g�}��^M�h��s�}�BZ���E�F��t	%i{ӭɪ�ɝ��^�����p�Q�~�R��)tƭ�s\=I���6�tW 0���O/��I�ú��^7�zZh��3�hP�X��c��Ԯ���c3�����C�b�w��B�������	�du��$N�<ML�*ȇhg�ڰtû��/݂x�{^r��ԅ�>h��n�RͭXzg��{�Fٟ/-�%�B9Q�������
�x#~��~�عF�ʣAF̨�# T'#'�p�ɒ|6��Yk�E�S.�H7��'K>�J�/��ų�ޝ~�fz�8��[�p^�����t�!���u�"����2c8��p���cQS��k�9Ϻ��N�U�w�K9�U_�z��n�P�?o4V���Qp�M�][y3(��u7�ұ��R��0]_O��BZ��Bʲ2I��'���3�}ڳ�q���%D��
0�|�J /�W�k��+e��'��w��W���=�U�nDR`��U�+P�G��Vk��-��)�`}d��fࣁ�[�۲��dB��쭜ە�n�(_��S�i��녌G�ES�G�A��I�kFc�cG�w��ֹ�v�=�p�la��/��\0�<�Lo�,`��V�x��6.��x�����z�/�u9Y���țlz��ˊ�0�~�)����,�9���x�8< ߕ����(��>�5F�79�v�@=5L7��y�ۧ�0Jp�f#l�R��\]A|�NH�S%K�9M~�R6���O���zk��(X�ꙵb=�\�qw�/��h�����z�dbY��b�ܾW&������P�C��������5�!\9�C��z������Tfr٤��!�# h�S��q*���(=��C�\���p��:�e��Σ��I#���V��wB]� ��d��N��+��gΪE5h-���<^$x�i
���Z�6���{{�a�����6s&��Ru<,ו>Y��'Y�s���ַp�?��]ʆ��D)zFΤpZ'ޡ���W��={�v�Κ%_^�<8r|��:
�`T=��h��:v�ԅѸ���W��oM��vTHv�"}}�]��}U�������TN����b�]L
NJ&�Xqe�P�oej\_���gX��C&�P��*�<9��T�OT�,�+�۬��p�ـ�!YЩU1Փ *<B�;;�P�=^��j�t��7�ϱ�ȱ�VS�c����w,E9��wಒB��i�u)��|X�mwPB��z����7{�h?#�΢r2��*j8;�TG0��b��\v����ֲ���"s�cs���{�~͝w����f�fE�tT�'}·��������M5;]Wl]��|�{��*�ֶ��^��o�H:��Z���gx���*QR�o#�b��R��͹;`w
E���͜�]��ħ���F0;k<3`��z3|�N�Rv�����N��~�� ���z��BUgc�\�U,��ǥd|T���k/�Gװ53�uv�3=��c���K���S�C�#�8�f�!�9��LZ��w� {��%!'��9�+��<Ϊݞ[�O2�ɩ�R�7[H;T��g���C"���T�mKb�������#MZ���N0��[�ѝ��Aѥb�Wd��S�[ä�-Y��4�c��S*�q�x52&�]V0e�G��S������޻�];sO�+�u�9p|�)d�a V�=?Ug�J�;Y���vK�-r���K�lr�0[����vC�JmY�{R�`�Uќ�~�z#׭�zv���g�����ft���t �%S��.b�=�Zz���/.B,SQ;ڞK�˼O�M�юg(�!�q1�NY�Qɸ�75�.�i_g�k3�a�m�V,	N�J�Z'��@,s73<$C�TeX"r�X�QX#�1��Y�d)f���Vj����}���ݹ�)H�eB�`���FmPx��R��Q/z{VE�u݊�sP��5���	�ܭ���Z�9�"X�̠Y�0J:�LJ�r�jk.j�nb�IU\��Dh~���=����/���x��^<�Ȍ2bxP���P{夷�3.��sqm�y+"�Pmq;���8P����5��G�(V�q�t�۬��3�����z���=�^��hK�U�Gq��(W����焎�S������R�%	��y{x���8�զ���[����4E#��Ic]M��Yz�Y�)ȟWuO�F�x�6��1�;�}R�"OC�@hB���VQ��
��k75���2X�6��g�'5��Ac|^�Ŝ��:��ى���>�R
�}����6��fn�����S��#����w'�,�������K���w�:��Vt�iF�:t
B�q�{9I���+�_E�aL�X��� �b_"mY�E<�j�T�qu��4�Z��ɞ�}���ꪞvnzi>Ψ�?��C�^jq'9��Q�.�_���ҧח��(lL0��L�
�s<��"z����sj���羲E���+��kXl�X7�+U��{Q僅��̘�6�6���_bØ��:~�RV��١�\V�ŉ5kVE�ڍ���r��*��zv�hx��:s�c�m\�C|)jPy���o�j���߱�b6\��,e�w
Og�Q �Vn�_#�o�^��*�O{	��LO��
�Ȳ�ɞ�Jwldt�Zvl��H#k�`��<��f�2��||z�g��,J��Y��V�KG��=^ 8Y���r���N=��%��j�i�����Ӟ��P�9:��Γ��KS>Eh���藸�mS7:����V���ξ�̹����j}6�>��P�f���MV&.�8��.I�$����શ�N�;�5IR�Y���8p&�"�"�鶌�����&s���BZ���E�<�_��:�p^��嫟I�]��ۛ�gO�P��Q��,�������{�!÷O���w�8 aǱp�3�LRӔ�]���P�m#p�W�56���(\4(��hR�󕹈i��7�kJ��.ⱌ��^�)���4)bZ�z̲�03��5,��2�}�	ж��K�5(�t���H��GOc������Ք����%�ё^�3���6c�����n��CGUۧM�a�pV�ƫ�VIr�r1��E�p�R���j��i�
gd�N�H4' ��R���=������QS�N�;%ةO.�
��P4���H���6������:���q�L�٪X\��&�<ٴ��t{�i�#����Sp���5u�u��rAib�~�|uu���egU7}�Ү�9m�;�8:mAK��s#��*Q$游\�萔��o�c��3�S���3�m��s�ʺ;�&�V�w�A�Ո�]V�����b�wG�YHL�讴� ��}��nL���[�6���sz��rAo/��k���H�ާW�k���Z�n���X�]�X��I����N�@tb����ܣ}��KSM\���`#�|��}/���ᢎZ݈��>f�<���nlȹf:v�p'�Q�yصo�mI7v,�rpx���!�%'ou����[�|՜��_������W�N�ܡ���·��i�D�o)y6c�oml�Em����Б*��>�ݼ򖧍$�>s.M�g"^���̽�gk�Q��6���ܠ��n�.�]-���}��Y	�J궷A�3^�Mi��bH\}�/2oSu:���ֻ�v��T�iȻ���_Iy��9n&�4�0�Q�:PG���=���KN���{��|�&�v��u�̉�ʝ``��Et�֔/��	1�p��I*[I@"/f�/k,�V�'��j
�n@K�:�����h]�R��M���/"��َ�Bi�WoX�o	A��*6�����)����6:�f�p|Q�f��ȴJ��V:� ��xx�j]	WX(��g��\4��
�$�	ɊR9�Pw,���Y�S|�����;�Vkr�RJ4m�ۥ���k�\m��u,;yh�Lo0��Uk���1���,���[��̧�Sձ��hS�!{6�Ѓ��Q��]�լ}�Ĥ��Oz+�[�U��"�VM�6Y��Ħ�i���Q�s�k��=:��ol�>��1j��(5dA�wSjGk%c�!��+���Xr��kA�n��uz�CsDU������۽�|k���(c���Er�-w��m�;���n��Z�����(���ocKg1�s��,s~����G
�jX|�jf�Qf�|���7�v����~���W����"Ƭ��陱�9��r��Q���s�u!R/�Lz�]f����+��S��=�R5���H<3y�ߺ��{ \�<=�ER����u���v��d��v��G�\��GXw1J�u\Sl%�s�Y��]�gDn��z��@Ď�v�r�Jܓ�2!��:�[x�����O]���xn�"�ڊ�j$���d�#(�E��0�)j V��Y-�U0Z�J�V�QaQeJ�ՕJѶ�ƕ�EF�b �ڃ-
ZT-hU�**�֭��T���kQE[l���QR��5ҲZTj"��ՌUQR�ciU�
����[QjVKF�EA�YX-����hQF��cR��iT��(��m��-�A�B�#KD�X"[J�-�X�0��(�+Q�Q�E(���V�m
�X4��ER�������*�YZ1Ab�¥-��J�1aR�H-B��
$X�-����TPR����b��Z��+m+dQcV�H��ձA���2E�Z1��*
��PYm�*��%�����Y(�,����"(*�ժ���ڊ"������?"0/<Q�76d���u)c��5�&f@/:���{�N��m�#��d����t�C��7�ݑ�.-Gq�3�IF���Ey��Ս�	�>��&��_�P���,c��Ԧ1'5�BȆf/Ke�ۮ���#l���%"�5SyK�x	~��H�}I��!��"��bX�kj���W���p��m�R��c�,��ؿM��l1����V��J�D��Q��b�o�*��׍
�Yٰ���R3p<�}9��wf➭$��X�
�@�N@��I��^O.��ڒXP��s�6eͩaT:�����1�ΣB(l���Q�X�L4@��P�����U��ʜ0�D��4;3o)�+�Ԥ�l΋�bٿa�/�V�w��7���yMKY"�ٸ(�u�?q\}[C#�K�s�zU��e�����I�x��1g�WAÃ��!�)�%��[�NQ�;UT�wO9@��-;��ÕZ���a9���Lj1g<8*�7��b�]��~�z
����Jh�/V�ƖN���}��.X��T�{�Y����ǎ<r�GUi��kr�k�ww��Lp�R�f+N[uåe`�a�$d�\�==C�1���.��ھ��n�w��%�=�:��a�cv��^y΂�f\i�"�C�خ��ͼ�G�mZ¤��n)�"�H�욱����-��K�G3G]Et�,t.���u�b�V%!s=�8�&�JAP/��Ur㽭�I���� �f�Ͼ����6E;�(��R�/e��\<�e���|%��Ƽ3#�ƥQЪ����ڶ�{q�uY���pb�[��Jo�}\J����!����yK�C	{��L���!��`�gN����o{5�� ��!��.�ʖұ�P���x��s(�w1�m1(v쎤�1j}WsZ�e���c���<;�Y7��Qag� ̴�	r��)�@�,[�R6u�f)܋�fR�z3���:�<�<5�͈˓
�9�P6'R�%�ŠPP��hKC{���<�hS����g�W��ٙl�C��s�%ي�]�7	��y9!Y����t=�4�<'e^��|
���5���'��;:[��T�aa����R�u�I����-qy��r������X��O҃�gٝD+�u�SH�~N%i�6�Ub��*\ϭ^++i�Upw�m�����ٔ^�K�<��w��3�'E�ן�<<�A]��G:Ykw6߱̈�
%���ʻ��TY���HQ��ʴ{րn;���#w�y-మogV:�+���Dq�n�tӅ�p}��E��]Ji��l���Fi2����$�Wmc�G6�m^����`Gvif`���-�+k����X�H�Er�U��p��"�mޞ{�R�V�V�nRq� ٧y��5ݲh�C^<�a�e_X�gR줒*+;�W���r�$5K�B�?G;�6�!�ՏNBt��+qpu1�{gh��tFu�z�X<q^��r.	��,\��I��=��g����*�T�8��5�jb|EAm�~��ǯ{�mn�Hq��s����\�fVipޜ�ɋQ^`X;��Ǯ�ZX49]l��ڄ�W��x�.�|�~��:�s��)q�n@��/JxWas�!�-�G�n��6���sL(s�N�t���t �U>,g��i_��A�o���aV�����Q��Q�N���*��"�#��%_bqE�qa渱+�ŏ���S-p����)��}��;a��������x�q|����TC���*����&҈ZwSl��-����̬ͣǚ�X9�f������2�ϔ�g��Ed��fT"��Z�$�m�������s�B��
v[r��Ok�DM�̠Y��*x#1ا;�Sm�;�w���S�J���X{aUpv_)��!��v�̈�& G���'Pŕ��Q�l^*�^;kBt��s�-��RO�*kQ�O5Ԡv���辳�}P
�;ҡ�oZ]B�+��R[��p6�e`���םT�OF��;i��.e��Nu%;�nQUj�ז]M��O+
���U��V3^����֏��<���W�,nm�}�{̜0ѱߢd�W�t�9�wyMh�
]��P�"��n��@m�b��i��n����$�yKJ��v��b5~�P�Ե7�Ď�%8�,����hl2w��)�"�
�i�=k��gי���֫DB������v�/n��s{������N��Q��^	O�� 8�!����n�e/�C|�9u(;��~��g��q�粍k�b��G�"{r�D�FŅa��uz-KϨ�{�̣q�8]�:@�5O� Vj�k��6�'˴��Ľ�߹��f��~�<n�� ED'���9�7�U�޽��A@�Y�*�{�n�6nu�qz9Q3g�E���Z9�*�1�)��|�;=Љ~{M���p�>U,�%��피[^Y^f����
	^���!�4'�-K���k}��s7�g�"��`��P>�{�x�S��.!�zl�m�V#���%�Ei=�3�ac��
��c�(�3�[�0�b��F�a��ͺ��d]r��E��RVI-���_S���twH����]sV1{��SX���H����%6�"�+�m̅:��v�#vfq"O�[�/R a�)���}g�gs��`�#���:e]r����kz��kQ�R�E��m�Ù�A
�������\=��0(󻭡`�ػ�H��[���[]�=��ξ�٣�=�1���/�@Ǡ|+�ܬ<�J�gC�0Y؂x��q=4�+GO���č�0ݟ.�|6>�����M#�:�i��1�9�9�z맕	 ]hq��$�%���Lf�����I�o*��vJ���ZeE1h]P��H�2n3G�s�}�BZ�9��	ʺG�x��=�,��>{�Wcp�鉎w=%���J]1�b�T'�!=<�fz-qR�����Jon���SI6xwyY7��'�u�����hK��Tƭ�5�B`�aܘ �X�^&F��o��IQV�����X�#�M/}Ut���e5�`�w�+X���[�i͏��=<���T<zJ�6:P�tEaO9V����Y�R�W�Ccd��y��gJ��[���|�hs,+�@�N@��I��^O.ᡓ�z��C���KN�{J�r�f�2��:+k�;jǼ�c\�U�6#�@
�rRyW�*p��g�Ml��ڹ����`v�S�U1��f-Ô]��*����7�#�������,|�n�se��N�����	��[P@4�1���fh�#W7wQ�µR�q�6�ֹ��>���3��,��Ჸ>r��預�I�\�Ğ�0������\���e�jo^���y;�T�:��C�c����J�<���ol�+�ܤ�&�q-��}�a��S-e L�ܱI�U�Y�x5h\/�0z�yk�ML�<wu�žW��9t�,,:,`���C�^F�P�R|�%�/	��߼��.��(z��m]�]V��J�Kr>n�d3L%|�Sۥu�{7�0�1�����nT�5�	���7I�{%�o��so��I�u�}x �]�C0�Zi�ѽ�[z,XB+��.���x
攰�=]���vI�繳C�i"E�ɷ�����#-��C�/zs�׆d�ơЪį�c^X�ˮ(b���E��P}�T�M+�}6��+�lE����'�e�s3�[DeL�a�܉�FN�7�ZGXH����'qJsϬ�*-��cx�}y+5�]�V����/��eyڢvu(�0�����u<L:���/Xp2Nק0���SS΋�S#3�`x�v��9��6'R�]WPP�e	�7�E�0?J
u�1M���Vb��T�}��a�1��^�F\V�&2<�J>�Uyh��������P�����׉�^�׌��=��U�W�f��;k��9a���ό���-�B��wr�0?n���R���tR+��pM��YG�vSDp�/-|�:��-��`��z�s/,:�xa�0Td�v��W*�n��J�N�@��i�̥�S���z<��,��YL(s,ha��ܱ�B1�I�V�)�_z��rc�f�)�)�pu�zxX�Ә䇪l1Ќ�N�5���vG��X/eOJ���b��Y�!��m�Fi��Jzy}o�����`���ן��]v�H؆�����S��E��K�ج��6��#�k�t}=�+�Zn;��D!��^ovQ�i��Q$�D��!��㕁�]�H�f,4�YڀX���S�����6��mV^ݜН,�[�nV�xA��`nG��7�U�ߟ�9f��٣O¨���_�3�u�03����˭���t�������:%�o�N��t㕚\7�<�b�W��L��1�FQ����Ng{z�	pw�չ��/6[&vP}
����:��1�{����)�F�� �bo^���u��l��&���]A��
�����PĴ����q��ac����ۯx�o�r��u;;�W���8��#�`����R�Ⱥ��0�^�Qg�qo蹮<2�C���!��RÔh
wyZ��7X�o�q�4
����ݕJ_!u��,*Vf׫�hjxFX�4xTrΞ�!]���.�5}�0S����E�|��s�"wi"	��vrOz��2�Γ	����XN�w^���|�v.�/&j��w�ȏT�ϓ=2p
�+�:Mq|�US=��h�<!2�����s�6�,͜[��X�72���S�f��`��<��2��),�_$=�.̗�Z6����m�R?�!�̺��w���V���VY�x�\�"oݹ��`�R��U{�^�%�����om��z;]D����(F
�t��ª���88dy��x������x���7m47u�Ξ����I� ��ʉq�t�_�����U��
]��ZEºcfT˛%![o%�AO��NV�N�8 ���<D�a�����.y/w�B�_�u�7�y3��;��Z5��U:�YcP�s�児�
�Z<3�Fxk����KFd`�n�z��/ɐ�Kd�����r������JB;������p��P!�a��5�Τ�c�7Ԛ�}tD-y��^v�-;�䨓Z�T��
Nq'9��^חr.�p��4�S�Y=����FO(�����g�Sy�qFQ��	�-� �O)h9�x��T��Ֆ*� ��I�Yꔦ��,��dw{����%۷�I7];�4����pf��;P�)�o/��bX�"Y��mA�i���|�Y9W7ٝ�Os�d+�u�����w<9�/���0���0��br�Y��?��v>Qb�&�����T�۔%�b��R���M��٠��k��(`���Y�j7N4�m�?X�,���^߳�ۼ�٩җ^�����C�,-K����]o� �g,.�́M�Ef�f���㕼��~��j���,�Pi����[�E��8y3�a����w*d;�'��NF�ѩܫ����Sӑ���D[�=�u���n|���RKG����x�ڮ%g�y=�VN�#������h�Zr	Cx�l�r�:O�o�S)��#ܒ�ų/:I�;���C�0��-�z��f)���l�5X����O$��]���P׷�o_35��·~�tX,�!�"�-�Z�/,��ӓ��]���[3�鶴fft��f�M�tSҁ!�IM]��ו�P�����
]1������B�*�����/(�O�RR9 1Op��I'�u��(NW�Ж1���R���Z|e<�S�^�Ђ�2��u0�͕���lXsq,o��H�rx���#�ׄ!�o�s:r�i}�dnݎ]�ܤ�h�;"fԫ�>KT��2B�o��gT���TN�Fs���ou�m� k�ʹ�BἋ�Z/�6��x�P��{ó��t��M�G�ܝO-�DM絽�k7�n���U�7cc��p(S�,������;�i��d���z�Tc��D�y�^F�J�*z-V�7�g\���gq����,\�t�����ME�q�(���ҽet�ľ8���8�e��a�s��z�9,�G��pC�Q�(E'3�\�U�3���}D�����U��zн��@/+s��S3mػ6��Z����o�Ø�q�Y�}5x`/5����"�´�g�n�ݗbzoۗ]�W��2R7Jr�����9���;EE���A��L��N�uߜ:	�%�.��Q/����(`���xQ�6�="byIp�\��s�+�}ҵ��J�r*׷�+H�36.��ħ"��+�`ͣ�8a�'΢����s����M:�V�ot庥�i�����9<�*�X��!�l�9�n�t���XnNQeM�E�nY��Ѵ���\)p'��"E�1Kd��#�S뇞F[yK���b�½m��K8V� ��԰���ݮ��s���YȪP8U�DױKsϬ�^yQ��R���|%�Mz"]ޫ�shd|9jWI�ki�JQ�D�cEf�����BS����\�}�ؤ��:]��h�Q0T��p\3&}rUӕ}l��ݼn�Cpڤ~�h\�mҗwWD��P��`LXq:yhM7�AT8�UgD��W���T��R�iS�^���}hz�KFk��[�x�n�J�@�A,TG�+4��(m�
�I��V��@32��J��+_N���-�ˊ���FGA�[͛��к�6�S���|�5���Q�z.	�EC*�[�2�y�X���iq�P�]y|�}�M���;��wܹ.碂��6�d���(�7��P@�\J�n+4&�߃�i�`�ϵ"�A)�b<������=���Zk��ZNo����X��E+�i�K�F�����<�W^��Y秩4�K[�ExN��[{n��-�;�3\�oe�rX�g`y��ֵ�2��m�j	7�LȆ�j]�5��M�3:���]��^oto�E4�6�k��wL�g"��6f�b����JVcr��u)��U��M���e�J�����L����{(f�w*�M�2�=��IڹlsrerI�٬�\Ok߲VG1t�6��jޛ:��f���+9W���g����4��s�*T��l����
żÅ��γ�ԃ���n˯�Ca�Z�� ڲ^œ�%j��P�o�5��i`9QvF�"���@��[ǧ�j��u�����"	&>+�
t�@<ݡ�x6�r���I�PZN��ԫ�`�#����ޕ�T8]��kJ���E��]YWK����[#G�s�u����U��s���gL����{^{ ��&�7u��18p�(~��J�-�����2Na�z!�ý���X��G��0z_v��B�SR��X�8wqU���BiB�t77K�7���D'�En�k���<��+��^���0�0�AI�Et�#�8geJ��X��j��!ぅ�u7	L`vyR++��A��B�b2l�zM�[����w!v�WN-�;YiR�n�������>�
��.q<��ڔF,�퀸�v���S�]3R)=y�}ؑP.Bi]Ҫ�>�y���[6��ή��/�~�B��<��;:&:s�Yg�w���Z�Hp��2�h̋_���q,��q���
�0T�)��4�Y�e���u�{E�7}׭�vu��9:��q��(�Z7.ղ�!��"�PŘn���3S�~���a�Y՝��wB�6���\e�ö�|)@�4��ue��ij��nN��L'�n�p��:������E&ܾ��=V1�B���5,�������w�^t�N�Y[\0�`ũ8������Z���[9���f)�E��F��,h�e_�Q��u)��k�=8g�},o�rg���Љ�eM��]�7�wttƩ�ۺ:��^�sJ����ߤ�~>̓|vt����`�+�C}~���Z�۹���'��(Ԫ"0XѩZb�F��mEB�U�E�ڀ����N"�(����(�E�+aX�X��֮5�DJ�Uc+Q�b�e�DYm�&!��R�Q�+YƪV,b��XR��EQPZ�k�f�Im�X,�$X*�#*[h�-��l�"�**�R�
"�T*����b�R�AA����1L��D*�TAX�Kh�[b""��Z�F"[,�j��TU�J����!Z�BV)b�("�PU�+��1
�(�[��Z��ʑUJ�eF
�X�#&�QPTV(��*��m����,[YJ+"��"T�PV"%kjֵb�YQj�U��s2+X)�
"+.%�%kUX(���mF+-l+m�AZX[F�Zʪ #cYV�R*���JѴ(����PQ��A��;?h�-<���t`� �'��W�`�r�m�{ےh�O�%}ec�
�F�d��n�V{�&�M���cmu���1K��ݵY���ߡ�4QBzx����z�TuĪ�qt>��|�@�;4&f!�2���ъ�qT_���ˮ��x���J#`�Y��A�i��v�L���u�n2���/ȯ)�%������Ϟ��n$5�w���.�x�*���xR�P�<*"��o/m^�}o`vˎ�aj�u<5f���K�-ܻ6�"�[{fd�IgB����@M�����/]m	q� l�O��O�8�)��Srr��#Q0��I�=��cR��7��<]���~Gv\ՇJ���TC�)��\4��J�.m����[ ����v`��j�Y�={�~��^��'��o�^��lȸ���C�Z��'z�wu�(2�\Y;i��>R�!����i��ִ���z+~o�L|�K�n��e[o���TL�{��[8�|��6!�ՏNBt��+����=�D9�w�l{��Z�=���^�=�M�^�� ��Vߔ9f�=�4Ъ(gñ_�c�ߨ�/�5Pɹ�Qf�YYw���WPP�ɕmQ|���썻�X���t]���E�C~���M��\����d����*��5��7�w�{WC����%��9ӯF�L���/����R�+T2ngOFwB&yvo;��Q�Z��>�N�k
����]Ը��g�0�_��اx�.H�K�>��P;/�f��CA~�r���"闲����Iv����󼮄��pw
���s/ct��bܰ�8��iq�M���o^�#ס���Vg�q��X���+z�uKL<�_5�Һ�1�y�R�UD�2��������0�~�Q��Զ�m*�aC�Wؚ(��!
�5�na���ҹe�����i��^tC�A����='��X�n�Z=>i
֗h7�5�ר�;=����l$r��Rxյ�"<�|'�o��}�u
R3��PP�ˆ��*�EWy�ݽ��_�����˫�'�sz�g�v[r��Oj��"v��>D�(�q���������s}��^�~���%l\���Kj���S��<w{�	k�~��=ȣ��Φ!�կ���)��
�H��(T.�.61��a����^,EּxPޢ��s�;{������uˆ:�&x�$��.��؍{J��/&�f�I^�%c�Qu�~ܽm���+���W�F�ۘYo��}[��<A�Y%��\�v>��2��w�F�Z8�����gc��</7�=f��{�.g.(cpt�Hȣ��[�5�,��Ge̋um���: ��ht�60���)l��(����Ω�r�=�8;�:Pq�&�ũ�5�U3�t���RP�T�=�v�2���e�y5rT�����v\��9��:�Z2u���e,����(o�g.*Pmudt�{���{��t�jv��tI��`�u
y9�t��#�{^]ȸG���zY5*2U�2�8ێ��&�Ĕ��ۉ���c#�i�~:0>�@N�� ��V���|k��J	D<��fv�~ޓ������4ϰ�����aoK01�9�1��C0�����Y��9����NT�;��<�V�9*��Ƭ���}B|*�}N��5���r[�������M	E�>�#r)�Ӟk���cW�R�\�\u+}n�����;��Be!�{L����$=Y2��oi��c{-�Ү�g�I��3��$�{�z��m���5�oc�������Ya�Ћ���(f�:Ө rf�S�Pц�9�Yz�=�=�)Ӫs)+�´��=���*���^��=Hq�f���-���{`��'�9��n<`��ٽ'(4�����Mon���h7E����{�SOKN��V¶�4'�<�cxf�礑�Y�p5�`���նzŮ��}�7\��s�Z�au�s�Ѯ0fDm�tK�ӒoK���}J�8���3s��O7����� X����w:��r��r�]��!Z��#�����v�yX�yR+!�7;̹�x���<C�]��
���C�S���]|uo��R|�@2��^���1=��׊�ڮ6�e1v� T=�@W) 	�l�Y]�e��Fk`�3����O3�}d�^a^4���eγ}�(�~��
���~� =①��J���!ܣ���kӥ�rS8�G���֏�c0�N:�p���F���Qȿ'P�����$�s�;Ĺ������
�Y�{3.{���X��Qq���It7��@����	�e;���&Ib:ݵ��NekK3�G=���9-yV﮲�V.�G1�cyX�L4@�N% ;�8Y���tn���O��]�r�B�Q=�����1��{1h���:X�kz�*�dK����о��Z1ʤ��s�1ۤ3�ۧ�K^���w⟍+��q���ݎ�\́��i��w�)+�p,.�D�Ŵ�v�8s<���{Z�⒒ᄺ�^c~���?a��Q�� ^��n
��ꆾk�%\�M�5f�aT�����N�U��l��/w��j��0�͐h��7�42������c�a��/h��,5�{kA
n�� �X�vp�OSz�L\ƞ3�Э��:1�.�Z��@`9:H�.v��N|�����t��6�����	�&��7K�Z������cIus�l�t�e�C�)vn:o:���Z"�tp�rx+��Wt��3��-��Ҳ�o��"�܌�r�+;!�}���*�F�?K��T	����d������#-��y�9�a���X郂TѤss��]r�,?�,�����^�(��)a�D>�ɍ"��WK����D�`nr2�3\&w��{TfuYG�������^�a�+���(=��C�<���UF^h}*�fQv����P���Y��Y3���P� G�=&s�bM$F�k5ssV�S��s�vE�\cP���e�\Fc�,�����S�����9���.�V��J�SO/9�	���k�e�;ʷ��axv]FB��e�abLdy�R1"�L,Tn#$^nL�=�}e���:��MO�����M�	@uLv|g�8<���BSM�R��k���9��L��ր� ^��n�橽(`��}���jl1Ќ��q+H�d�3{���Ҹ�>Wշi��2���M;�����U�]<f��U$�
L�ϱV���Z����9B��!x/�^αK�ԹrhVbwÛy�q�h[jk璹���ۇ y�T(t]����t�r��R))�7)���1�il�׀e.&0c��7�*����nv���vG�|����Ŵ�[uP��=��%U��Rft�]^Ox��[[%_'���;1�^,��&�8�q+I�r�6��<'ǐ��5��᷊������mGV�2�j���o�<�4ZJ*-v�1a;���Q�:�Xxc�r����qp�X�j�����G�����A+������(<��>%�r�&y��q�o�ص� ;3ʐC�:$Q,c�=�'k���o}\wץ��eVzC�_�ؗ��اx�����+4�s���\M:Y��ص^�]�F���H�4�B�i{��������:�^y���"��=Ț�5o"�κUZï�9R���_o��~j�R;HCS��N�p23�nt ʗŇ3N�T��ʽ�F����V��qϩ��t��{�0�}��mv}J�!@���C�aqE�S��ZC��%^����PE�"��f�>������='���f�g��n���_�&6���9^�G{ŉc�J�M����Q��f��`��a�ݹ�),�_+��멭������(j���)l�:&��h�����V��]�ԅ�8�6���7�����c�Ӱ�Ȼ6o��wh9��
>��1u�]��y8��	q��ou��d�Q�cW7k��1$R�Y݌�l��n����8�W���"o:nvRW��K�ꆲ�V˫�'�sX2�3j���z#4���G�4���Jďu>N���i$���O`�L����X�dx�R���_�P��W-}��e�^[�tE�ӳ�6�_Q�O-=��!A"xd��O�ɱB�v2�.61��a����U�y��t.Oav\,ͅ�`��WR���!�x2s�	�`
U�GAh��M�iu�%
��:k�θH3�kg5�e'�}�-ue�FA��bAK�҄�(�~��V�F�!�P�]`����"c�Z��P�4�����>�z�q��z�P-9�' `b����8^GH�C�w��)Q�	�s��j�xZ��GYnh_VVUNʕs�� �[���@����v�nf�$�s^�S@WO��c"''����4��:0>�@N�� ��򖃑�w��fSK�mv���j�}��/�+�4Ӱ\��q&��ٖP��x�t��ŉ��%�MB`~�͚���=��M};�ˍ;�ӍbF�^�]a�����=˅���4ز����یz�#��$`�V���Ι��xvN(�ˢ.;�h�Q���9A�N��vƤo"�i���s/H}PѺ#^4�a�כ,i�('o=�m����F��\�=m��sg`��*�=�m[հup�����"T��U- �tu��8�C�������-�Z��:<�nX�T���k��_�x�3�Ixa.z�=5��a�Ŧ�J�s�wwf=���y#R����i��cz�1�蕗�q2ofpR73<.c23nU��5C@~� ���0ml�i��V|%���˘,���=V�����r���A�3vo�Z,��*U�ih<O��'?
Ρ�P�9�z��t�b�*
E[���fȟ���Q&��W`�L�R�8+�yg�t�~[D*���E�[�2�u㥵:ӣ3�ʜj[V̪:���0�|����]E���ԺcV���e0&����iW�C�j��y\.�Nx���m�D�"w�'+�	c�� �0�z͜�6f��}Ֆ�e!��Mpб����tv����b�FG9<���S�n��{���gK��S��D�)ELh��c�Y��E��r-4&�LT� e�J(�l�ǹ�o/������C�㓄.� w�j朁�OUc�atT�\' F@��a�O.��U��t��r#��юjm���C�LK�S˵�X5^(�<��[�Z*7g�9n͏�ZO8���Ex���b|H�X{�܏�� (�E���sOZi�:���ek7)�Y�2�5�Sر�Vm �Xm�U�*��E˫orv�T�vL��:���Y�N�� Å��x^�ESBp��ãQ�胼��> /Bq( �vR&K�fײ{��3z'J�ڳ]]R��yt߅��ًF��Ōw��"��n���j�J�p���r�"}���E���a1���D���N�ćy�8�	�r���	��E�6��Y�}����|7O����h!߯#j��	l�EJ����z�OR����#a���Tl]���Aȧ�N>ž�K7��Li�l��+��N�2n�qn�?eԂӠ&��E�'C TNO}J���b=�[uò�ބʪڙsks7��͍�\���%�e@��L�x��n�Q>�h�ay�-��nt���3�-I��U���o%�QyJ�멃��Lk��p8TE�D�,<��C�yQ���gOv����ةn�]���Vl�ɑϪ�<l&i�K"C���򥴬zRz�sX�5�ѹ��k;1���הs�5��B�~�,���9(�0� �2'HK������^۔0�i����x��D�v�rʧ|zA2p���z��ݞzM�-�f�1z��sUs+q�g���yꗇq��jjG�c�2�[<;iЬ�-�u�v�
ԻJ�]b�nt�gyJ���������R���[���>�LM��֜�mH=ٓ�0���O��oKv�h�'����S�9(�X�Z��2���Í��Ͼ�����|��TA��k�P[Ҥ�΅=��9����w-�LP�c#�i�+O��j\O��o,$i>\�y��k�@ySZM�U���U�����,:;���}1@U�R�H�ō�zZ$�2z���;�uSۀ]=P�:�{����lW'�<�v/t�E<IL��Qu�?4j��`LMEm�(��L%ޞ_[�=xo�`��	��Y��k���=I��R�ِ��p2Wu7�Uo�ϡc�Q�!�J�6�Dc�a�A���/�a�LL�f���{��z�����vp<p�������Ňq�,��f�q�w�svCE���zs�1���p��.�^�qP��'���<K0lkι�jD���"z��Ϊn��ײ���Jg��7�\��zC��~�b^�b��.u]�Vi�������	�[�U�6{]F�@�Y�U4k׳C�f�ʈ���wc2u��?�.�ϼ�b��^05��p��c`�y.�w�m�eh�(�md;2>˦-�O*��v�����ʆ�3�L�5�f��W��w�]X�t����O��mt��ۃa�0�-R�b%Z)��`�bwK�˾gi���m�U�l�����G��ռ��r���$%Z����Y�(kL�$m�EU��4��jy6���u	�IZ\rme���,r�e)�*&�u�\��UX�f�L.�G��U���^Vi":��L�mQ��@:�p�
f�Vt��/L������c���� 2�jq����B�Q��ىb�v�,dUٻպ��1)�٦:��BX�;�����LґDE��p�R�|�uʾ�]O	�N�l=�P宄lt��(u��V��9�r���cD�sF&�
��ޘ�m����خk��r{]�KMl�i֣��'ܩ)1�\��}[��O���,}6��V�O-T6Z��A�,=��i�bG�`�B�V<c9�G3iS(ho��gJ��T�`W'���l�2u����.ӽ7�C��3Fn5�'c�|1@̑b��>\���IY0���T���֐r	o�V��W\�6DV�+�疰oe��g^�����=۷el�
� �q�R;�4A�&vm�@�䂮�敖e�X����7j��N?7 �����!���nŻ6�zJ��k�����r(:�(X�d���v�\q��C^��:�ȟ�;���6��ͬD߶g�5,a��)�$u�)��W�/�=�q&ǀ����hY%�*r���iTzue� 8h������)��OCd�$��Ȏ��!m
 eCM
�&'�:L�J�¥
�[&���Ӫp=�Χj<����B�f�Wp�}pR��O����JT��5Was��R�4�s$I�5�<��z��D�m�m�Λj�:[;y_r�����F����W�ьs�d� e0���Ks�����<����5�!*K.�:���Z�[.���-�@�-�pݣ2ιwj�L���xWV%.�u�k��������g�(¬n�=����c��[�3d��oDiMy1�T���i���k�e]pTPfo(�}[�w9Z�����%; Ɲ�|���$����vKA�"1J��&z^�W|ge\R�EN��qTM:Jk���h�/�wv��/�R��e���t�Aq�|LR�f�ZS�Mo6�Q�ӂ��qR�Fq��ݚ�:��K����w\j�X�Ҝ@r�X�x: VY�v:Һ����o�#��L�.�u���J�5�.p7���{�.�rt�vJy�,��ë�QAu����ͼ]�j����ę���a.���6j�Qx�:���t���]V�K�M��`��:Bs��u��U�څ:�mnuX����:f�e�õ4�X�ݡS��ȼ�"��ʹ�Yʶ�ծ��������ю�s)�g��ѽK� B=_��������QU�����b��J�V���EUm��e�a(���*)S-��ڶ��f*��6����U��%EU��[c`�QS)��a���)�Pb �m��� Ŋ"ahb���EU�YB�\��(9C2��E��6�.f
�2���fUUf&8�X�EF+l��ffH�h"�B�h1*6��UdZ�[q��AV�2��QE���Qc�H�8�m��""j�UPTQ�fU�R�h�����8��U�F�,(��P��EB�Y1\E���ֵ�Z�T2¢3��Q�Q��m�h�m�h�&4�TYmƠ��(��TlADELlD2�Z�[b����\s3��!�����*1A��Ĳ�E��Em�ne�Ʊ֖Ŗܴ1l�嘬��3��h�Qj��*.\Lʦab-l�����.91���V���R�4�
��e�[J��Sˑƨ��ek�S�2���9As?{��_�ĕҀJ�rɒ�wb47��[uEI�#�O5��� ��tzwj�Y��sk�z_q��.��RL⬆�ɪgo(d��>ʌ��S����|`w�(8�@����΄�2���E�,u����wŞ[cH�jw����Q
��*��"�!@��%�S�����{;��q���A�a<=����(8='��3q3��Wb6&Ofo���e���Y=�}�-s�&�c�(᜜X9�g���l�􋌣Ȏ����ޭ�m7���׺���\���s1�b��y8���-쉵t�N����"7���5OJ%s�6�{ѩ�xr�0LL��B��P���c��g�ʫ���pE�n�]4�	�/���x��u.z�q�:����WԎ��J��?��>j���������"��]� 3j7�)R�:(V�V�2}�p�lJ�|���F�&�n�1(U�:s{F#Շ�Sy�7��~Jm�P�^����na��uw#fH�)�����p���^49�-o�9:ai{�Ջ�ӫ�����%q��3�k�	�F��g��G��)�q�g�O1�R���|��D��W�JJ��H�'�}2�
*�L��[�Sf�*EI(!k2��Ը��Ǯ�fь,�[�v�-�S�G��ޘ;�چ�Һ^��YKy����Z8�!�����u�Z��I��.첬�o�Sz���z����{�����ո���,�4��<�b$��+�<�Wz�ce{
��E�'9=��v��l�7��G"'O|�}x�>�]���|��=����~ S��o�[��x�mf��S�\ͱ\ܭVr�VW�%E���������:X�z�yVb4����x�Һ�#VLf�tu�=Y�׽7��R�Q(4;W!����j�/��+o��k�wO�짚_v�x�5����Sc0�}\/��ƬY9��Ɠ�|��WO�X(��6%-��Dh��¡W����v�{��Ӂ��]:c�z��q(�`^7�X�h� �e�����bZtӔ �Y��+K�2�øE�ӑ���rgEJ�(�9�P�gI7O.���j����B~�2���P��E_P�,vQ� �m�"oPs=]�Yo�~�riݺα�w������6��z"�lk��/.�˅I�c#�Nɡ}60E�4�v�7��WU�0�}s#�Mn������D(P�_5�R�QOvxߜ�VN-��UXܫV��!��N�1�cg��*�(�֣�7f��ҟDq٨H�m���Rd�M��B�ܳ��W��(s��VK�~��2��r��k9V��]}z�i(Ҧ�Y�\���-:5���^�g\��z��6B�m�s�˚�m$�4�hy�޹
�<7�+��byf@��$ �p�tiW�xi�37��9��x�Z�{K��Hj�9�1Xv�g�=s�	^wO�UX4���$�E�Gx7X�L�Ү��Z�$�*&(�ɯ�W�+�u�$3�J^��D&��V� �D���H� G.�|-nG���no,D �nxD�΍�40u�vhln�f�22�o��# Rs�Ğ���&�u����ZZ�h��~�ORI�����઄P�x��p����U��
ġ�}9�� ����T* >rR쫋�<UdK�]e
�޼���ɐ���hǕ=�ŵO;��-f�,�S�pms�++	�s�"q��H��n/�E�׉C���i��]}��R)���h;�y����r�uFi�E����'��!����t�ɝ�3-< R�ޏ+G���
��twL��:!�Ɇ3S��DշLt�=�~��
������x$L{�[�/y#��t�'�ҙ�Q9<�ɆtS�D���+=�<��&j��-W���S���R���m.������LEٹ��a�`-<`��u��l�m�\��3�q��gL��snּ�C9*-�	�NW\z�f����3ƍl5f��b��9ͺ]o�=7���N #(U��3i����eN��oqr.��撚)wS�5������/|Q�Z1�՞(:�Զ�"��OML@O�#-���wv*�~gt�ܙ���nT��r��sި�&hx��#+�T1̨6/��Q�Xod�z�� KV��KOs˛��H-�e��
��!�L��L�$D4+���;Ԫ�l��2��ǲ
Wj�;�m�2�5d!V�܆���j����9+:�DY��pX�8׮w>�1d�y}��}���o�g���`w-���ui�u��zi��S���e�O��6�O,�]j]�TE�p��E_�Cg�ê�^wZz���.�!y�K�t��~���X��^M�$�4	��J��L�Uqv2�
b�I�ZP{ӊ���'Lpa��Gӻ7�+Ct�OL�E��!����RI��'�(�u�LvP�gwѠ�[�s��tZ���)u����V�3ޞ�IxO0z����Gp���KZ���ϵ�g���2��(�IvuL����
�����vh1pyk�P�O�k%�4{�{:=rZږ�>G{�u�l�cniv�l,����n%�n�� ��&�����9�#�J�Z����[�,���� ��x4��Mr@��+��9Y�9]�%x������=x������;�`_pGn�G`
�#s���t��OI�S[�Ze��LvriL-.�3#���Z߶��N��nvp89xëa:lozѰ{����g��àA�}���ҋ/r�Ь��=���Z���&��Rs��9�ph�l�u�Җ�1봤9��W+�����+�~�O �,Y�H|��l��yاX���؀��f=���x�3�wL����Z}�zpL�z�����C�11�.3e�:Pj]P���6���j-���.(W6j���9Cqɖ3��g(�aJ���^����<��p�O|]b��ۻZ�����Y�c�y��sSѝ|c��Q��;�[k�A��
���Pҏ�����'���KK�;�M����X�R�z'ח	��\KKS	q|���sa��=����7�TFت��"��~�Ռ|�E�L�7��xz�٨�N�Q��qSv5��GgMb��k9P�665���ڙ1 ��ޯE����*�s��P�
�kc�g��ѽOO���+<N_�S3
��eCה��aԹ��K�{����z�^��yf�>�/�]7a<����/�26aa�53<����
�Q3��r���nsu��7]�����s� 5=���^���WǄ�u躣�}q�A���gjݘ,_S}��(h&ekĤ{�Yt�LZ|�������J����Vq�Y���t�Y�o��k]�SkΞ�ņx!�;l CR�O�s��X���:�a���r�*���JCĩУ����r�՟t^<��x����c���5�J�Ʌ�ò�.�\��V�x�Mw��N���SM�/`Jؾ��<땖C�²8g��{F�\&�4���˷9P;X�3�)L�`����%�_���ŧ@hb���+(�42l'v:S4�T�5��x����"�Qw����,\Gs�MjqPS�P59C	�r4��k���η]�O37�-y}f���Mߦ�.��fƌ���Ki�"�c�� ��lgJ�Wh��^�]-U���o
�ʿ	�(x:3������x�y�>����N�~��A膵��j7N'::��Vz��zn*�
Fr�y�p���C����0������w0^�-]�cR�߯��y9�J��[aUw��1A������`�}%�8���]'9xh�t4y|�z����Whqr���c�)�ˈ����L�0��b!�a�c��о�u����IZ�f!k)M�%���RY�:��P[Fޑ][-���.!�'nӅ�'&:��6M�����8⬽T9l$�ߚY]��򏍝�4��c5��Ž�I�х���o���h�F��-C�i\�
}Gr����Xp��qwk��C�'C�tq@��	������t�؛��f�!�G^	t����v�V˹��J�(�x��~���L�W�u
�r�Fǥ	�M�e���3��(;��<�lk�J�32���;���eц*	A���L�Z].������m�Ok�ۤv�1�>c�VJ���y�y	���E��@��'ǰP��+d��K��������5��b���Sʐ�WR|�E÷O�<���gGo���D�!�a
|<��p���]���
��=��tƦgF�V�����b��E1a�1̞$�qM8��)�UNR�|�H���hs�b�h�ɡ���W�+�u�D�y�K�D&��=����KKI�`�zwj�@�~�t�\0!cn/PJ�Cō���T<�P����L��=��K
�uA�F��x��yw�Ic����ve�6P�.���_پ�h���gC���^�=a����Oo
��Q>�޼�U�s���+�ya)����2ч�+h^���J�4�.Va@��lܧp���
ܬ��6e�w�0��#�ے�z�i�re:+4X��5"�U�d�Ã�ی\�h�8�3}�fN�(����h�C+'H6@�s۫۝�)�p�L#9���`�tf�;�|�UEl�=3��"��HLA���Ջ߼�0����K�(\x�y��q���)��f�
83�B�R7X��BZ��26*Tc(85k�N<�7�X���/�6}�^({jal19�$��*��h�ޫFl��%��Y�U��jwq�S(��n��;kk����>˺�G�eZ���Ȱ"w����g��򉮖ȿd�`���Ꚋ�s����6Đ二fR�]�y��R�6{+P��&���]h5랁5�ٌE�S�b}C����Z��>�ԏ��S%^\�ϫ���|�{�����d#C�UӸ��XjP��j�U�ךq�k�G%s�|9����t��x�f�6dr'ýB�C�676g$���x/�V�k��.����3+�Ra���p�Dp��G���Z �����C��'����ɧ�XcMG�bԹ���7�y��|�����w�֨x�/k��͜WYVݭ�COJ��"}\&��g�=J��j6=�<f���9� 7�^�ʏ�*�q苍�w�z���P��X2��ݝ���/_.�F�w1s0�C��0��C}�OP�Y�#V�WeNV����5�1,�ϝ��g���zG4�.��M���N�aqV;�n��r��>���!R���gfoq]����T����&ŏx�]wb��Ν���ԌJ멙����2�2֥b���j�mw�
�}����/C��(e�L�"±B��֒��J��r����k*����۩�v�W���c��orT�e����B@��k��HW���<���Gp��o�����Nd���I]�Z�sq��^n����2p��8TՏ�����8�C��k7����c,�&cԒ�W{y�{��a��U�S�hl�U�}l�w��^Q�����o��^|��ݹ�=}Xm>��_��/(P�;��[k���tF���H��3��3�E� �G���m��G�.CojD���~�����ze�!Em`|�D^�����q'�����/%�a{=����Oc���Y�z����^��6�{�<\�������F�-8��������1r)�X��%�~�/Jxn�"=@��P��{�mMٮ�6��k��-,��uJ\�~[�g_��������ܪ�]�R��)�=x���ܯns�CwD��\�2-4�rɑH>�s�j��ۯ6�T��Ȫ��˗�,Mi�~UK6E���M!P�xi�[�jd,����9��.��	B-��'nk�4�]�)*Sr���%o],S�Ǧ��=��*a�L<��S�<���+��ĺ+K7��!�	��j]!oD�=�N�a]���t�ǣ�w:���q�U����p�I-3���UV��[�&�c�p�Ŝ�3��ۊƪw;�?x�2�f��?z�-"��傔=c%٘*��O��辔.k�/���6v?R�q}�GB����\�>��")u��<M-�t�e
��*�ȳ�R�ߥ��^wf��p����\�Y4!�_+�;�\��zX"/� G�h8M|(�t+}��`k<Y^��8iۗA\y9��{nv{ٚg����ѐ������3���|��E�V�nu�r>��޾����))(��\"қfDT���R�(Ob�&��겏����]�f+��+�y<���q�{�죨�Be���W���\�:�Z0N�t��tX̚�� ��5m���^������Ϳ���_7����p�1�%�6'X�؝P�-󄫒�Yץ���iwV����]ȸӀ�w��Ϧ�&�.��f4X}����i��7�d��~m�(��b݈��f��^�ݙƷB�OӺ�=W%-�{�$X9U��v��!��(t��
A�P������6/�Z���w��bf'�\n�p:���[���jt��F�̲�X2rHr�veS[����+bѳb7`t��RF%����]�o[��`�ܳ�v�%��ye��n��$zӝ���_h�Yn8PV������u1�s-v<����"5*�7�V��+5<�yƊT�i���lr�����*z�#=t�8���2L^�kΜ������&
�y�F��f�͟Kt,����¦RG0U��k.�����xoT�W�C%���d\�K�u�X���$c�c�M�7`ꗘ�[�+� �3�ʅ� �!�ի0.Y����v��w���ҩ���X����!ʆ�$���Z��+����ɘ�J3;�����n�9����.��e���zр�N��U�Է��x''�U�[�kk W��_ʂ� ˬ�	���f^]b�9�����0\����Qu��2V�Gx�W�қY��5��f)�bV9;5��,���'����͵�x��Q<�Uzpz}X*/ݒm��*f=�Ir+z_u���Zk߽���nf��w�ޒ	�	�گ:(HD3�Ү��jn�v��4n�(K��
���+bط4�%8b��cl+���Q�x��֓�����gWc�-�rmP�<�O�7'�ʋHjŊ:�=9] ��'d�G�JK�/k�v�]LfZ�q�0K��s�ti�N��x���j@��h�&ڀ�7�z!eh��EuM�4U�@ʗ�i��`���iT���ŪU�gwi����W;��j��.HG#ҥ�<��P�@�:Ri��xp�J�/��懆�YhZ����"�s=2a24�9��m"��j��5tt��T-ɘ�f.6%#��S-���8�:j��t�qح;�Aئ޹38�6f��9�"�߁iV��m\u"�Q�7�����u���pƣ����-.f��\��ٕuc-�1۩��Y���^�v6T����([��p���s�n���,�p�S�&]�Ǳ̵�F5��	Y�f�E��!ڕ�ٺ�;5�`��X���d�c�d;g�N�/[˒�z�^��B=�ɭ���ǭi��������ɇW�tλ�4�v0�rھx���V��x��[�C�]*��P�R(L�NݫX����X;v@(;�"W���gEpסk:k�^q㦣�X���xq��Qw�,�So:�Z��c����|m2���p��f���[�Y�PW��w�;$V�(�H�Ud���9wQ	N�gEں7Z>�<9�N���9^5��d`/s:�����{Qsnȥ���Y�;��5�+��a21l.�h\�*�ùN��z�6���QG���=�p�=��\������f#eP�Q"���QV5�Ym��J��L����X�LKF4W�`ZT�f	W�Ub�(����jUr��E��qQLj9KmA6�ʪ��-�F��Q���baK�J�\Le�q���l��b���Z�ƙjѶ���-r����-X#��R�

��2�ʊ�R`���Z���V֫�ƥ--��B���[J�\ɂ+�-S3*�KJ�T,�eVڵ3%E�k��.a����b��ơkJ�[�D�b�2�c��q�H�V�#r��.+R�[a������B�*�(��"#��b�ѴZ�-k�B�A+E�G*Qm-5�(��P��fF��TD�U����R�he+�q3+lD�h�J���B�
V9fe�[%[h������J"[m��*#��KkY[e���Qq)Z-cn[Q\�D-(�KG1���[maYZ�.X%�bdŵqU-���-�cakj�1��ܲTĪ�fU��ԶʣPEq+R٘a���Q$}B��Q$�+>ͼ�Sa�9KYĩ[��iۃ��r��T����!l��3O�|���P�Ռ�S.��KgK��eB�'9p������2�]��M #�ה��)�Z�%<��CaA�5\���2�������̎�7Z��Nc��\�T�t�~���Y^{M��V�ٝd���z������
��藺"h�Qg%�w���=�q��V���\͌E�-�b/�)VӐ�W��V/�昍�7��1`ۻ�H���.�gȘ�B�������+w����Z�P�\^���mߌ�`����]��^ub:nDΊf���5��g�@�,w�|b>1L77���,Z�.�)-x��-����u6@�r˝�A���B�����0��-�E���5��W`���r�H2�eA�t8f�]I�B@����("r�JE`�Tי�>����xS�`���C$���&�����ei���"_9�0r+�t^s̠E�`�Kǌ�˭��N�9���yXI�����B|�E÷O���h؆6�(9H�@�u�Ȑ�[vj�W�M��[�$�ؘ���Zn:U1�\��^�n]��ylX�:Ȧ/��0��RYӜ@���evb�P#����8�tzƬ}�`�:���O����L�g�cs���������U�uc��5�o�f�8gH
��.�h��9��.��uZ�נL4�#�]!`��3Z:�wd�ϕ�z�tԽ�uouo*�<OޙB���7¢b�����c��U��g��������4r�nr�t%���nEpp^Q'Y#����S(m:�Yٱ{��e�g�Z�u�!c��)W��P>��8]T}�h���AXZ�ё.��<���-��h{o��qVcƺ���\c�(� �rRyW��<Q+	eݪc��ZMnm��ݜ�m�ojP�j7��F����������+ݛ��ڷ4sd:�D�7��PΙN��ƫp�Th��!�dŢ��aD-t��{Hvjݿb��{JG�t�8'�&bq��Aj�������c~�cum+u��zJ���<JE=�q�-���p(*=�kJ�s��+�d���2�k<S�PjDpV�$�&c�V$�}��~��9�Ȋ���5y�[9��=�F��c*�(Z1��Y�h��!}R�᛹i��GFbz;�������ٌ}/zX�7;Ԯ��B�Q�U~��P������T
����yfP�>�x�k[�0w��+�sv'�*����Y��&��Zzp)�U�۝��R����W����5A�Wx1 s��܎Зmb��pHʊ�����w�I�]s�if�}&.��yo�$���0-����);k)n-���Ų���#�N�C
_d<ʞ���,(�t���2%�D<��c5��0� ��"�vު!�Ի!�����h�`�j�.�.<5	��w��L�n�MҪI�r7cC0cX]HRu��j�SV�[\lg9�z�}w�tcY�f���ЙdV����c��~槮��ғV��Ϩ(E[4%�6] 6�m�^��F:��K��^���Y֧�nX�'��u뮹L��Bpsq��"8�K�GO���ɬ&���٪��*8Qq4�جp2v;t[�״5�:���,u`��)$6�?�S=yw���Ѕ�w�CW�Sԫ7gb��"�M�,EQN5���vGS�ؽq"�u�p�݂u�5�ǽF�՝6�sΜ��}/1��I���	ĭ7���2
�f��
,��n��fV����Ɔe�G=�7Þ�#dCެ����0�v��yD:X�AF6�¬nu�t9*ZbF�9z�͜�A\��+�����3`A����J~J����/�H��AZv����>���fR�I�v��T�
5r��J�T�S:�_
#Ħv]�xIŔ���KH�=�սN)�5&5�t��J�IJ	]	��Z	.����o.��&%��:&��l�G��S�æ<t{�t��iG���}��-߫��Bf�A
���+���s��!\�n9�Ό�#'*���v�^9T���l�0��+4�oNy����,����T������!���{�:���J\�:����o�{�v��ݬr��L��r�������P� Gxo�<�>��oL�J�ĸ=����T�<Z�tNw5;���}}��,����U���Y�?.��ŽZC�T�M�G���T�X�R�z'׉�/K�LW(��rNU�f�:<����l�$�%㼒P���!ت��#��o$���"<���<<���y
���]���S�n9�w<l�!E�2Bb�ىh�eO��\ׂ�u\X�Ś����ڜ˹�, �ןI0�`W��:��3�({~ʇ�2,�:�<��׾�֘젱f�Y���CY���
���v��=,����'�g;鮡0F��Xx��u^�wY��W�>�nkG\.Όe
�J�؇Y`!p� "c�&U�SS����*���7Ϧ�z�O�o:H�ŗWȽ�t�o�y�:A�&� �Ö\(V��H��!M�m�VOv�٦�����@Q:�'��}x�Y�e��)�k۾i���'a��٦L����o�}�{�_[��(�],�g]򻾼{|�4w���;�:48�3l�������0ƹ������fQ=��MS�f��C�>_�*h�[�9��v�̌P��W�@L�r9:B�s�,ݬrޭ��0cdjUه@W$�q�X�����N� �;�_�+!~ݔIѝ�p�w�;�����r�h���F	e܋�p/�geO�.&�.��Y聬�:B3u=Q��"��9e�U\�n�$\���x>�Ձ�炰NܭV`9����Ŋ�}��*i젴;州�H��i�u��V�L�ݫڮ~�,�/=���c�jy�����i�5��`)���W�Xl�w��g��4�����3K�����������n��ȥX7W�;g ~j���<�Z�����i�視�� �_[����\����t�d>�t����n����C�tg3�Y�4���Յl�o��˙�L�P;�t�t�Y��7e3r_w�zGNdI@^oW�8��n�VϨ���i�,(�$�~YN�����}d�]>�L[1�<�yr���u5�0�s���7�M�Om��N;��v�Ms�5:�@����Zc;QWE
5��tV~1R��O�ܩQe���J�-���0V�R�s����ӕ�\���q���
5��YO��˭���t*�3鰲�y.�j���*#�Y���=�|"nWZ��Q�Ďna�+6{�i�AɆ6	i0l$�L�L��C��ė��L����8�v֪B)��#���	
�Oi߹"�����(f�����Q1��,1��s����J��oh�Aʕ�ܺan��C�o�ȷn�Ǖ���G���VM�H���՝�;7#��gf��8E
s�5���:����K}���<;Fuܷ<�Ⱗ��Dr�똝���r���A�I�k�<!ʰD;C8ؗ��kj��k�	~�Ǯ�E�.����y[U�w̌KO�Ⱦ}���x!�d�[�F��yh��Ꭸ�cqrڳ�J\��ŝ5��6.kOM8�� j E��+�Yw<�%��a�t��T"�b�A�ֆ�{lh��	�<gk��~�y�W6�`�."np�I��O���\42f�>Q+	e݊�0mWL1�z{#OKK�O*1,�^���ci��{Z�!�XN�:1��H�*R3�ns��H귞���N��n\�!�	�fуr�ÿl��d\K�����A�E{\�!�9B޲+��"���/��i�@=�VS/@�[�b��\�+u�Vʼ�n�
x���q�u;��z5�֍&�E������oso{nw�髅�Pj�GM��-Rí�#��ϴ��m��o�A5t@��7z�[�ڛ��纜���|�da����-���O����᢭Ł�g!�Sn��+3���0v�������Q\^�a:�,^X�������� ?��>��U����T�#���z���e�����������"ΑX��/eWW*��[ b-�ǩ��"C�gU���M^^�aۿg1�Ƥ�5S�;�0�m�̔b����%d��wHZ=f�U~�5=�-��a��6�j�m��:�"��O����ki��3��GB��tWk����4Rb����eft��t`\��\��r��X�ϧ��v�8us5�~�,�x�5��[�,�~�ݷ��bh�a� ����`W[��T��imq��2�[�FcN�0����V�Oe]��E.[m蒞�~�;�lԢ6W

V�F�SJ픪x;�<�q�Pj�x�,������B˵-7�Bp��@��F%WS3(WE]��`+�:��{Z'x����]��׎O���K���#���_Jac�q$,ƢVu3.���V�2|�j�nep��)�+�cb�t�`v�`�n�^vt
��i���c�(��/���h���U�H�q�r �z9s��)[�({n [��W��םxv�6"�e��RX������%QV`�Y;��"�_f����%�	%ϓ�S<�;�ÿ́:�)�tg���"�m:����w���!��=����t&q�^+�E빼̈́=]5�J�DSw}(�[��P��@l	¦��>�v��Vx�q�l4���w.�rnl���AE�.U�ދ�������7z�Kvp<p�寰�5�*���-Vdi�p{���}��R�
f�n��eP>x�����׋��tF󉃾X��7�7��9j@���p>��d����qC�~~{�m�j
�,�d|LO���-�O�;��#�{��%��k/�����W0b���:�������Ǭ�*�ئ�
��o�\���إn����myE�\��/ճ{�����D;b�Sv�+=�bM���z\�#��<��ݨ�0@~�19ި!��P/ا�7�R��c:]FMS��n�]�OrF��BhoW;�/5�D�NÜn��T�8�1�+��}�Q49R�!�O���KN>��N�`��;�^·yۭ��:��RQۙ�Lߦg�e��UFU�C�<�M���p9N�2�^�1�sY�
�����g9��{����`X�x��ʠ*����T�6�%��c�W�z�K��<I��'s;p�V�&����S���Sx�&W[7�Kte�ЬW7\��{�I��+�R������k�D�Y݊�����by��+<O�Z�ܫe�dtxjuR�ArB�f�3(;�R��v���ިA2���/[ň��r�mOX�/{�qi�-_:D>ۺ����<�zR���.gҒ�POc�N����7�NڞR��<A|��į�R�a��`���Bx�����Ġ��Ӫ)�<�[�yx֒J�J�ʟ_r���GN��)M�8 ��'�R��ڭƛ��3b���C!B�)j��[,į����|׀�gF0�ӫ�s���Ԯ��٬N�v�)Xx��b6�z$�����[P�2Y��밒�+����:'Q�DԈ��6	�r�K��xYkIܤ�k�F ø��ܗ�%�|��ے{@��C�M�X���BOk��k���-b]�uN˹���H��O�.a���e����������QJy��d!��r�ߣڬ�v+
�e��ͬrЅl�P���߅iİk���������Q�V�F7fsC��k�� �P��"��n�Ntu��:���t��B�E��J������Km��I͸�G��p�ױ:J�'#/���8����#d^����Cm����D��ugZ�Tr�`]��v�meb{H��R�s(k�f��;.��Nt�]�*�͐n|{��F��̙L�9��f`��5dt}��e����^Ur��:��v��:�Q��	c���V��"��+���vp �%[t�l���w��p��Ӊ��j�k��;G8'[œ=���
��/�7����
�v�GK��,n<�9�'.ҳ���t%=�>ñ���E��%a�ˁs��xx����S�R�^��|*�����u2V]Ű�}���Zw �aEi4��Z����O�u����WY�xu��9t���Dp�,���\��N�#���^5X�Zl$�`�I��*�uG�Cqf˺V��A�w>�&�u���Z��kh�Qko��V�f��@H�9�z�uԫTc�s����B��Z:�/ʕe,v?5h|��μ�qK.���͎����^𮹖6���~�ɹ7���<C;օʽ|&��;
]1�\�ڨ�9�w.�^C�b�5��mn��e*͆�2:���&��B+C��lK�e5�0�j�<�y��u��n�s<�D�X��\��Lt��X+�����$Z[]L�G�YbƸ�qA39��{ݺ�@1�"+���]S8Z��W�n�'�}�Y�[ţL�u�} +�s�˖0wT� ��gYBQ<��"%�<����AK�g�Q�n�7�.��;w�6SK5T�Ӯݽv��NhNއ4�2�J�� C�C�m2�����	
�W��ΙXé8��e]%�/�ƹ���R�rw���ΨS�"q-�qPe�p��[�܆�>�H�k(��۲M�G�r�+�lǊJ��"�2�[R��"�z<�ƃ���-��V�딺�nk�P����Κ�땨.Թ���-ջ���=V���x^.�A*7�v�\�p7�`�C<+*:��Y�P�y��uFM�<!��$f*�6������v!5IӦ�޺fxǰ#��yw�R�'[���]L�#)�0��p�Jݾ��:������t6�H�%�g)��S��+��R^���;��!X)��2E')W:��H��/iB��q��+-�|����gi����{��&��8 *��ij��aU�!�,�n�~|y⚆�2�����d���S5Y�8_Z����Uۧ1���k:��KT��xe���Sz�.i�d� ��T(�q�+�ƈ |�m�Z]��76oV;���^��u�q4�.�4�=ҳ����jE��w��q��;�*6`�,�;��R%��n�q�尢�P_�滄e��{w�q�()Ԝ�1�[�hT��X�iv��kl�c����A5Pڭ��'�bրi �w������Vl���"7rv��;��v�%2�@� .l/ޖ����[����u.�kaE�a�2��h���Yak����ᨬl�.��O-ܣ����[II�h��
`��};rJE>��"�;�ך:a壁=�w�"%��q����1C�[����jjԹ�/*��Bz������\�7�Ƥ������&�f�ݗA:�F�[
��+�"Vһ{���(�`Wk�n oq
m��O$�����\4�x���n�wl|)'�
�:�mo,̤�&��Ճ�o3Gmm58A�,�9����a�ٜuԺ8�B�V�NV�C����j;*��X4�?e�ooT[��+cԢǠǆon�wF�ʾȖG�J��IЭ#j�q�@�����홦M1�Y�����#�k��O���ׅc�됩���fU�#���(�뢠Ըᵁa}"H���p��b0����'�G��>�1K��1�zcfw�˞�젟�.	_]�g>��2k�����J\��\�۬�Շ:k+����P�久r�8��S�o
OiM�eni[D�����M�9�t{1*��k@t��N� �V�ՖGe+��,�ނ������-�.4�)�ͼ1gv�s~�Rr�-U�9<s����&!�]�eÝ����*�Um�)�"T��4��̬�G�ĕu�s��A����Q1�	�Z�D��Z%Nݕ�,�
��7��� <`I!id���֒�eAT�6+.e�em(+V�Qƣ-�T��pj�-,[[i�0*V�Z�,�ֱ�p�\l�X�Lh"*��+�Q+DmD��Lh�+�VR��iqE�[U�Z�c3)%ʋj��Q�E���d�ZU�[in&&+pk\�pʴQ��\��f5��.1.L��-��ĦXZ-��m��m�+[j����qU�2�r��X�Qknpm�"���-QmT��p��E�PR�\�R�
5+Ls��r�*V�bS3m���ƙUb�mQ���L�KYl\d��fe)E�0V�ٌ�LAJ�-pL�\D�2�%� Ԗ5�6a�cEj��(T�"�ʭ�2֍�JƣjR��
���E���+���*�[Z	q�+bQ�l2̩���[�[b6��aAG)Ls-�崪Zcqj�����U��-�F"(�J��V���eeU���̰�1�M���g��ֵ�4��ܘq�����3�I�ܤӋTJ急���Vg"b�HI=ަ6:����^�$Z�/gd���>���\�v�Q��T�$@�����7��,�K��5�s�jꐉ���|��B���gW-Yٸ�Ga~䨃[�؛s�	Ġs�2��U�C&l����K�3n�"�o���y�+�*{R��T9EH�����J������1��e���ofV����K">�{�(_�U�76�C�^����/�񥮑7�i%�5s�3W���-�p���G�ͺ�^�o�X�r��.F���#���nx�(��)텘^\X������M�<|�Y��Lv���.X����'�%U� 5kG��9~�l6:au��|��pl�4��aQm����|,h��q'(��\\���/�����F�Kewwe���L��=5�c�I�&�Lڟ2'���g
�b���X;kS�e���-T��k*�r۹0(=R��F)A��C�N�����+zZ�a�`��=�s��<�rڹ;u���rDo+�����j1KrY[]R1�\>�[�~����a��T9)�
�IcWĠz�����+����P/��xr�lNj\��s��TO*RjŻ�Ӿ�D�̙m�{hXU1�zK2fo�<��:�4]�z�b����L����x�#L��X_���ב��������pc�	�Ę�����ײ)���R��L�h ̰� �S�ґw��g��o:�[[�ݻͫ���cr��-�\u-ح\�U���.��Ԣ6WP\)=
�Ѭ��Z��Y�h�G�/<&mR�*V���U������X�ۈ�Hė&fЮ.�P&U֥���Ք�N���q�0��,�\�=ڵ����aa���X�sqP��$����s�U�1Ҵ���'J��}�+s�$��W	�����xe\Z}8U�8k��g��**5	�+MX�{��Q�Cx�Rr�w���i�`b���^l���	��̈rT���@���AΫ�^�A�}�i��#$�z)�l��o*�3ѬNÈ��$��sz8<��_[�g����n�R�ԛٝ����	ClՏJ�!��>x��2'�yX�}����(�7j_O"���S;x��=��>�n��C�_:�5f"��t=�B��-��DeL��QN��{;���c��ݺF=�X�Kώ�Ϥ���Ӟc&-Ey�7��=�f����s>�KD��l`W�<OZll5s�
�K�e��!��������p�L��YS0,uZ��!$��/mq����3��q�&��-d�Dތ2&��+4�$�}jjlV!s}px3�����JM�Tv��k��YG���M�W`��v��;3q���֚C�ܻ���������!܊n�9Y�ۓlo��Ҟ/Kms<ů�6+v-��ڶܣ�E�a���tΖ�N�D�vXΗQ�������0�)�Hѫ<�4�ѹ��7��z�F��;Eܙ� �>�Y=�ȣ~[d1	���]-9��6.��5�tdl��C��X��88���YRx��e�f�g��TȎ%p>�U��x�=��Ѱ���.u'��*�Q������;2�g�u#��|�P���f`1�`#�朗w8f{��5��R��TNf�M���;�|TkϤ��S#�'G�=[��Wz3�a��$����L��Dhӓ�u����8(_�7x/<�,����Z�����*S�<"���~��o=S8	z{�v����p�.Ό�(W����:�g ��f�tB�	��ɽ�{���%"��U�b�Z�����m�Y������0ƽ*tZ�nrn��T��ku� pp�!�
�_���j|����*׎�>̌WuO������:-��VC
�N�ؐ�X0t��xqY
�*MwȭM�N�������������4h�AU��WYV:��N�es��v�]�p�e:&�_J�^���@���T��-�b��Vn�̮xd�.aV�Q,�Σճs��ӇQ-���m���QLp}d鿢�\p)l��
�P�ܦ�yԙ,u�,�V�D��~U�V��]�����;Sr�{P�T5!&㜍5�O.�!`�{��,���qW�z[
jɞ��k/٫�k���q�j#��Ki�"��R�r9��^םq6���~PsMAs�-N�>�˫�:/Ԯ���뎟�B���l��'f�ޖ �^ZՑx��t�pl�|�,�9��X�Ȟ���K�W�d���Vz��
�qt7�´����_����0�����U�t����vb{}F��_yr�#~��cM�f8u+������r�w�9w�]sKʾ���n���S+YU�hnҮ����J3ԕ����
���ã����W=I^E,���
�8���%Ö����C�x�r���O�q��<�@*�h��V:J�+�"f����ǹ��Z0�>��m�`�M��S]{��Zm&��OT�J��]����K*D�;{Y���8�I_�B=�m�,d�f�L�=�G"dV9�Cg�EB��[B��.L줽=�wKV�h��N՚�x�o�e�)�R�t��i����NV�+��k,d}�y��6J�GV�#�bn,]M��X�����[\��`C���\^#�|j�cC�r�\L��+M e��5b���	���]��Ⱥ�]I�/@X��2;���9zu�bc]]:,_���&�T\�u�F^�[��U��z�ʈ�[�n�|S���MXO	)k�!ް��C��ac�)����<Ĝ��Fu����S~�H�{�]�u�<%�_0�_%�:�C��;ﳍ�yMmX:a�u�w�NvSf��tz�	y�zjl_���pXКe1S�e�Jei(T��z��m��Ts�ᵛ��fƔ{'�>דq�n)��e��,u�T�_��# W�����.ᡓ$��
�Y�2�nX�9{\{]������:�,u�$j��b�8(����#�8a�*��t�r&V%N7o�"��*�`�1L���6X�kz�*�`\�i7΀��;ۉ�Y�"�|�w�6�%K��k���V�{U_!�6�C㔠����ϋ�ߐ싉w1w���_ ��ڹ���{�)�m�ͼ���F�`������U��X�S�<J;9��U���D��+޶��=Vho	����р(�[cǞ�^��_�b+b���\�S���O�J������;���֊�cu������TY}��2�b�_��=����|��NUin��W����qMH#��Cp�lzXĊ���p��H�1�
@��ݐ�5�l�� v+���0�;�Qt�w�uM��QS`��W.p�kWf�_	%�}Z�1}�L3�"C�l9�mv<�~�fR6ϥ.z��h'i�y�0�$'6mNu�W;�(��ԤM��b(����c!��v�1�t�%���c��lƸ���&���-��-@�� ���E�y�Ә��B�ֆC�+zZ,73`�7:M%./
ܬ��f�uZ�Z��h<^#��qX.�Ϫ[K�q�1�<G����wPq`�jO=�B+n~��'e���a�ΩCvk���(�3���N�w�����R.���s(��G�!�j��8vz�vC���=Wsˠnu(��W�f����~��|�U�����=zע��^<����:�"�����(M1�����fe
���L���^��j��]nZ�$�|XZ�N��	Ս���/����I|j%u�̸��ъ���&��;y���H�C�/�M�:��:18��/ņ5�Ȇ�&6�i�a`3�\q�k��{��w}}{�^�����W�SfG@tT
N%i���h�����WB�k���J� c17i^�&��ʵr��<{��;�٤��+���cӉdZMM���V=w�j�Li����4W�����|�ע�-��tњ�1�=�v�7��r�+�Ǌ��G�rG��Yݝ����7�q���+�ܥ�#wl��3Y�Cm4xm�C��L��Ѭ̈P�;�A��V�<+�+}Y���{W�5s�����ۑ=f�zjv�C�g"���V)�.��@q��&.\ϭk�|�\��'k��n'x����^�%gcX\��K*�����3����}��Dכ�l�|V��o�����P�����N,�E����v6�*
�o����쥖*�-�*{Pcò��y�y[��ޏ�o�}�!܊l�}��^�U,�Pia	���]A,�������v�຃WB�w���y/[�N�.�j^�(v��N)��\��]�?A7ԽlUZ1ѡ�T&�ɫ<�6��b�},"�a�d��͗�ν@��)��}�������L�N�[����ʪg�"��*���Nj�����^�1�\�efm5H��<4C�3���6\���
����6:%["�X���Q��_�ڲvu�ʟG���)�Sz��Or*m�LHW�(��9Ϋ�˶lH��]���u�N,�=��Bg���a���e*H�.:��ͺ*���&|Ar����j^'}xf�4�GK�Ş�B��
��b�v���ړ�*$naТ�fQyWRA��dp�b��z��.[�6��r�s7;���2s����٩�v�ot���ֻw���������ȇM�R5�9W��
ʝr�����;����g�dS�ae�d��՚���;��?o��*�q	��t�f"�Z��w�m�A�S^��l)�1��^)��9z����X��H)[��$��g
"�5h�HWm5|��Į�ޡ�'����ΑEOp���z�֘�dao�_�����Vc�[(%|��w�n�ؽ�.������<'�����������F�,�cF: ��Wk�0Ho2�b5kD��u�ۃn��3۰s��_;?OS^�T�mT����_���qs
<�٦����)J�c��[��<��h�F�yͩ���ʗ�|���v�r�9\]��ԁ��b������i��&�[owg/P�앯[����	J9pI����yX�P�d�n�yU�#��2�+C�*�c��;Y�*dJ3߷
Xޖ��پ��r�+S�]�\ջsw��	��
oZ�'"��ZU�w�z���'������gJ�ހ\�$r�s�`u�����]�V�]��*V��\H��ັ���aǠ���]�3	�5nΆu��\��}��u�f��Rn:�;�MQ|f���kS����j��L������U�+R�[�zm�ov�aT8vT�D�q���9��-7��w�7/��F�߲����"�_���~��z��C�D��<j��*�e��Oz�7�-yr�{B���^}4���r�^N1�ݸ�m!�N��9]X�>̝o\�w����R�<fG�v�sx�R4�x���l^�/��Ƶ��O-=��""�w�����F�[��A�QUv5�<ZW\M��=�X���\5�*+���%��*oO��ⷦ�V�
x^��{�����^�=�mG�f��Kg��>�8�)LD=��ηj�s�o���܌f����˳�g�z��ֺQ��,�M�y�ӸGkF����0z��R#�敹x�Ȭ�g@�%w��{����u�`v:58m��Lm���m¹��L���AD܍˷�v���I:��2���z6�>wS8�Ԏ�(l��˵����.�0j�lp�(�3Zz���}������������,}���j�]sN�Zg�3n�i�P��X��5������/����=��lz�� ��~�u=K=�.���o(����h�s�����|w���n�!��"C���򇦻R�WS��7.!���޽���C����z���8����l��,{+"�TU�QS��b����R�\\�;}7wݝ��f_�u��{�왵I��r�����g}��q�;Yn?(��.j/O�{V�M���rN�
M����[7R�e��K�>�Iv�1�#o�쏍���ٜƞ�bf�m�&��xo���+���g[|i���+�U�41�lOM>w�E�f�J̎��Jl�[#,����Ҟ�Ŗ(޴�]u;Q�:{Ц�i��'�wv��n�FZ����'bm�!c���9m?.x̝��y}W��tڍ[e�畧lE��=}��镶z���v��w�5O��t֬�ޏ{����	!I��BH@�섐�$�$�	'�!$ I?����$�bB���$��!$ I?䄐�$�섐�$��B��$�	%!$ I?BB��HIO�!$ I?����$��B��HIO�BH@�|BH@�ي
�2���@I��N�������>������     � $    @
         
   l�.�Q��ZT�v̩� ��J��!Z����f�\.�F��n�,�	��;w
kVT(-V�y�� �2��j��ڵ2B�k6��kQ6�j*F�f�B���mlF��e�kCKm������m�}�zT�$m>�  �v��ػWX�.��N�m�z::Z��B��{��]+�����\:�u�q�v�{�^�ͦgZ�Z
��)۶�Uv� =������U��t�=��h %�=Gg�Tm�6a���H��٠�{���`���({իl��W�8lk[6�  m` @  ��  
C`�  ��p�@@ {{�   =��`��v޺;Zwn���pݷ������swwuV�.�j�lm�T6����]�� ��@���i@=n�eph��e�)��]1@�hn'A�uݣ�"���wu�ö�݀U��[���*���֭M)����  �c�{�˪n�PJmV4�`=���W�����g(9�[E��]��m��@5!��p�;$�b��:�T�eo  x i�c�i:`��������;�Z�6 �ji F�ؗmB�WH�lj�M���Z��  �HKjK ki0P����ٵ��+��s���m�Aq[@�5���Ҷ����o   �"����� �I�fIE�RH��3�)Q۱�"DwT�ؖcV�*�o   3ʞ�XZZ��7Q:5�@;��Œ0�ۚ5���������t�l�b�;ְ	��̳� ��L�3l3��A�B����)��r���
Y���V�9�JϟT    ��&�R��0F� d224  �{M�)T�тh�0CCCCCCL"���QT���     �~��U 4      ���i��#F(dL�4��z�I�P�J�P��F� �L��9�N�<���S���3�9W<��Hg�o|딾��ޅs��ʴ��[�TAL0��`5=H
 �Y���.  ��qU*�� ��)Ue?_|�	��`�#�HR��TAL��HH���TAK������Z�=��sᐈ�) �������@�g��=5�;t�e�P(P��pٵ���JX�����]�Ȯ�5�wkܼ���r;�p��M"��{�'�.�aS�˪ː'��ĺA�P��E�J��b�+x�]!�7�������}����t�C��:�Ac�lԸ.��@�p�wc�kl��Y�%����9��]̧4t1N��j�%A�vt�{�]�a����D��\�U.��E��`���!Q0}`O�70�b[���ݡ���eD�,�^]�a����p���ѝq�$��U��H�wT�\kco�9�݄Ș5n��kb�t����Y,lwh��L凷�nu���-{��֌�$9Q�����mg*�j�k���S&٭�����n-�4n3��3���8�(w46m�z4o�dX.�.u����؏'ENogf���������)�wY#��8	ˉ�N��Μ����m�I����I�ww�-�Au��Nĕ����o
;ȑ�n�g��G��W59Ocu���ȉ8,�;�����j�v)|_ni:&I��f�&ʡ��pUI�}E�lQoV���L]'�D���]���s�A������]��&�{B[ws���N���х�.�#���к�aL*b=�$ 4<]l���&�=_Y�p�����tR8:�]p�^�����A�,=�m��&n��]�X��u)��:e���Z��,,m�!�V�"�;I�N�㼴<�/Ў�o�&1��W��wV3��6��N]�R���,ոƚ�ľ�{��:�*����Hx9`j����fwf��ͫt�����`3x�I�o!�z�C�C�on�;�|r�
L��J]�X���?Sojn���>��O��Z�	5ົZ�|��^��t�(����r�o2��{�OX�x�^���j�����7�\P���u��a�ۻOż�2�z.F�;N�s�<��\�1`Z��Yڻ�`Qע�LЛ	.h�p��ٸ�KF��>�)И���t��g�����h�G HHğj�ǝ�$_�٧���,�p�s����3m<�K�.x�/+��f�D^��a�=m �ǚ��"�'�Nk�%@k����#"�O����"A�5vԨoS�.w'V����9�ŧ4�$��N���Ů�7�x��f�wa���������u��{v�ڧc��Hh��+b�5݃y'X50&�ծ��R+7hz�����O%9�á`��,�8�fH��e-�C���|n�d[;r��m���;�p��H��D�pһ^7��7d�3O%�j���
�p#��g @�X��A�j Wn�ۋod�7Tl�v�y���p��h\�KGI�c��7z��;ePop���J޴Q�a��m5o���,n�|�Zk��)�[2шkT7��'G�h�i}p��Υ�0�<�B�%!8��G>lQ���FD�>�.�s瓮�%ct���]�,<;v�Ky0�ۅA�����Uy-�!4S���k���Hk�	�ń�sq}},�хna�&�L����yŌ����ԥ�΋�8�I��k*^g%���gN(aqt��@my��;�A�ڳR�Ɍ�p�oG>�2xr8�97�[{��ߎ�Rγf5��.-mv7����Αv ޑ϶]`�e���&E��j�^v�_{� ���3߆�ݎ��Mm����)�:�
�$x��<��wU�2�{8�s���c��{_\�t8�� ,L����A��͛�4}��h�9��	G�v�ܰ��P��{�EVv��ʂ�j�����xlL�fqIM2]�beŜQA�yXͼ4��5E�8��`��x����v��w�q���kΠ�i�&��pN.�˥͓�EZfv�@N,��R�]����ܷ�9r��7���Y��3��g�/I���u��n�I ����*A�ű���l�]}���\�J�`6[{t���4�,��v�7���8��� sH��oS�{qH��S����^�&8�㑠ȝ�ɕ�h0�x��Z%��{5��	Vh̛�wSG>���u�k87���cv�{�u���	��5�4�t��Y����4��|�Y�������;q��$�r��st�&�W��5���W<���Y�(RI��c�_P�����8��0�7���ƥ�� �н�ӇRг�]��]��ؐw��vy���60�GÚ��I��.��rS@�-�:=��E�h��E����9|�zrQ��K	���n���e��h�;أ��-ցX ��u����ki=m�s�cKQ��ޕ�����Gcٹv8������e�֊�BjQ��>��nË�n�]��ӗ�7����Qc�D�k&�:��� �\��D]�]�~�1L�ulX3�b'ru[й��81��B�����q��^��r�q���6�'�������9c��ga��4��B���u��`�0�^+�#���s��zI4v�f�f��)PJwc�i�{
:.ҳo
]z�����;Z+H-�g�m>/;pf�!W�j\�����
��Esc�n��t�R�f^��j���K2W��7v�(�FłC�-K9�%��u����+nv6�<�Ń����
ɑ���u�h��1��0ÛGuw���h�7�x�l7zUPVn��s����4��r�R���rrD��O-�\}�m�4��}F��f<��#�zŦr0fj�!�a3u.si�ٽ�M�`:��a�9���Lt�2�ޑ��́E0�8_^6��q:c�
=��/s�����k\�7��с�}���v�QB��v���"h�47�0�'_fM��:1i�]���d�.7�2����}�θ�T����h���a���L��g=ˏ����t���q-q����#��<���Q�wIp0�*�%\�����Ӱ�ȇ�r�
E�*�d�=ۻ�ȱn,Ú�����n�[;��y�;h�:��4ym�9ci�t� ���5����`�n���n��$�u��B�f�^S�ɸ�d�M0w]�gwt�w:H�H�R�������`?LX��ou���&��~�񇷞�@o/���7Q �Î�WxM��,k�vH���M�-�3���L���]9�N��qr{u����7�z�-�ͩ�c��hN�2�]I���=��6{8��s�ޱa�5�ܽi��xكb�	�\��^�ǔ�v��\�dX;�g�^wEW����nY�C����sf⅝�)���rpB���49uN%�t[�.xc�w&<yHh�T˜� �Y����u��3դ��9lͷB�$[S{��yC�����c�H�ݥ��o �S&��f� �'aW%�5�̓vi˅!���RR�3X[{r%�	�Pr�����*&ٱ�7
+`wu�;�nM|���N7��`W-сsP����F�Vcp��&7MVl�ɣ��{�o7w|2��A��"�&i2��;{J��x[�e\�'Ԝ������4㔮��(�q����Y���A$����`��ŵ͙
Y7zH;F��/o���7mB�[��y:��$���Wƌ�[��u>���a�.�N���(��yx���I8]X���^����(�����5Q�������hSF�� :�uA����]�2kE��z������n��Lp�d���f\G�+.���w�Q��^q�k���X��4vk��#U�iZsN%4r2��ߔ�Mp�i�.
�`�κ�I�l|2"�Iѵ=s��04�y�x^�k�7Md|3v�;�`�v��e������[���=w=��b��㜚��7��aPn�N�(�Ǭ�mָ<�8�z�rv��p���u\3�C3�&�s���Q�:��.�(���EJOV�"b��Q�s�GG56b�x��mqq�ˎ��[:�޳H_om)mΜ�c�E;p�Ti5�ˎ7xlT���o5�Jk�WpF��;���@֊�r�/i3�Vh�qm7�_\H�@��U�Y�;9��.�-F���"��V\e���j\I/������[��n$ط�.�yc3cɺ��E��v܌w���4mء0>�Blî�F��`�wocA"�&\�q=��I5b'�놜Ћ=�ktr�P@1;����ģ�(W5o7a2�N����`�23e4)=�^S���G7�dO��/Z]֢������M���>b���k�v�)��Ʉ��*N	���BW�� ����ή�m��oCtc��sV��^��xU�1�_6n#pv���.�n9vq��,����E��Ƕ]�N�����;��k^G,�˵����"k6M�Nv���9q�5�����ׂ�q��i�@�M��Hv��N��J� {ăL��5g2�u|,M]I�!�1���ћ�4�f���FL����d�j�OV�fW���-IQ�U�MJ0��.���y�S5��8�J�.�h�a5��ˀ�jB��B��o.�	����er-��:d�lJU�����U�ɏ({�yx�u1�Ւ4 ��n���\T� dȶIϸ������SAjj���w��I�a�ՋON۴:b���U"ՓNE[��X��
�yq�[;9ogl6��ͭ���T�Z��{�ת����iZɄ�(��f^�h��4�`&�e�p5���7yS�+�|�kZe�О����2%Y�qw9w�&��܍�ut�� I��pn�a٨�q��w�p�zwpZ��w�_lN�{�(z����F�S����8{wNw�h�{�m�C=���`F��
�!���f:�����ظ�N��$��7�M�V]W%Lz#�/�xsZ<��.�k�U��"eۣ�*>�hW�K����2����Q87���������������Fr��0�*V������0¶��ƙp����rt#�7�]XS�W}����W.Ψ*;����"Y�e��&mb�N7^9ֹaƫ)�..C����ʆ���R�.<��l�����|Wu��F�6W;�K%'�}2nj9�M��k��YG)&62z�k1�[�+���:Z�&E�.!�Y��E����Ӳ�����90�1g|I���od�`���oF���@{;���{5.8{sw�j���?��ko�R�6y,�� �[�ْ�=q,B�M���R�:�`�֩�&������t:��Î��#��
��͹��m�Mْ�,�V^吢Y�Gi܌*��q��R�(s{�+�m�����z������xݰ�:�R�����_M����:@k,�k�>:\Y����28So�93U�����d�'�3�T7t`(Y�N��W��<�̙k�{WXܮb�(K~T�زh���f���zL�SLD�=��s+c�fB��HS׌���k)|�\-;��@ d�a0��w�ţ{�꿿A��5����on1.��/җ+Җ�闚
�� �ES�BA��\�E�Y.����{��s�̽� \��r�T�p%��6�P�ܠ�.�,��iKp�jgŢH�c�Ǿ�������y�gT������rd˼.�b��K�^zqu��X��W�9�=��9�k6�t^�i���=�\6܃9F��.�.��o�G4t-�{M��{
��;(V�]���ۣյm�L͗0��&�����u�J)��ǜD9��Sp��l���R��;N-����������-�$q����}���ޙ��ߒf��/���	-��^��<uyjD�ImI�i����)�vn�u�	6Ĝ�4�*5�γ\7���ˎ��}��-(�8+T�1���a�:�{<[��V{
&��f��{�ujˣ��䢴�V�6E�Hm�F\�V�k���Z;Wt�VCh�8�����u-N	������@wE&�����N���@VT�Z�3u0[��͗]�f���� ;�^�j1[Y�Y�K4��ð�j�KA+�2�;��7[�k�ۦ.u!xA(����qVd���3]��gdh�yQ���_,�٘�Ѻ�\]��g`Q%ҏ�4y�T��k9]��M��Q�;:v��H�F�J�er�ܘj��*}Ħ�tkw�!���Q%��غ�ξ=0/$�>��wϓ~�(�-�9u{�ɖcQ��{=�<܂gyQ28�n�ǄI�c�i�Caf�������EV1���Q؅hwVu}5sQd�Y��Z�!��"nk@꾳ׅ�q��cr�'�����k�w��,��u�)ϯ��9����������g��ͿJ�
��i���R�l�Cn�.�\�h��i�뾜�L$����~�Қ��¶2�/:F0��8���X�X�@!���(R��O:� ��վV�]-Č�ܔ:��L�Th�~��j�|�2�b5#�+`v흾#����į�EJa�}W'f��P_Q׃₽q!�v��<�!��y`����%u[S\��tr+��tR��xw��+7.�ۮI�2��
�J�O���-Yx�S�(&:��#��=X@./jޭh�<��^�v�5\�i)|�ą6�nЀP������ҧ�����EMT��%BZ�a'ۧ���t3!\h�Lf7_��	Ʈ��0�wy�X1fֽt�<ы�n*C���6r��j�H�ٔ�b����[��O�x@�+Y���cD�Ͻ�\o]�������Tm���HW_H�O!A�h{:�1����8u���zq���N�;�ڦ֤ޢXь�Ί��"|�x�5�T��;J6�yK]��b��8����f�V��+z�<4m^���wuL�3�ˣ�u�(o{�7��w*s -7S��� �@�w(8�C�i�9Sj:JVh��R:�����vÆ)sip�-^<wқ�V����T՗+�ɦ���a�X�V��a�M-�W�$f��9�hו�*ѧ��Y�t�pU�aH
��c%��tC����C���r/J�+}����F�g^Ty��3E��w�^y��H��}z��ݲ	n�%Ĵ���ڻ���8�j��q7؞�jl[2����iʳcU���8��s�Fv\r���2�3\��X�ƹ>�;�T�h�ı��>�����Eb�bu-i�f��2����<r�u�����]�[������|�đJ�H��D�@V��RK�c-�vIw��^b�C �R��澢�WY)�X��t�l#_^]%u����IL�%���e�{+/d=kt0�hU�Ub��Ur���VH��÷����* ���r>$�++����ͺ[[�t-|z���!3V�>�lU[2�����Ӳ̫�u[y�v[<�:�����p��F┏+<�z�+���oN�.���&�-�@_�`��kgZαQ@$����SI.��>���J����5��B�R����a���x�����,�R�5ƀ56z\���p��cq��E��bJ�T�I�Az�=7�Ǭܠ�-{F��R��Q�>>9� +�ݑ{���8L�z{��f��5���R�˘*�73�'��L���$*�r�Y��(�KK}��O4�T�Y�'e���:8�#5'��:zg��u� ���F�uw��w�f3��:�`�s%E�{���BEcŬ���}/���zu_��X��g�����Ť�'�Kx����r&[ HsTwv+��!�9��>K��B�1tQ�W-��!T򆌽��A�:���kK�:�8%��݀$��ip��CuR��C��Z7J��`եT
��%�UNub-u�.��a��]�H*mHU�k��=ݧi��� �]e�}�^
*����r=c��ndQ��;�.�	q3�.��u,8ւ�&Y��,,�t H�Y�7r]�A���9�`�O����V�얦�+ڮ0}z�Z#�2sy+)��S��N픸�*��L���v�6Z��ۊpE0�l���}�>:�0vXGO ��\'>/g4�
r�g�IM>[�{ۛ�H]�2{�$��� �xGz���=�D�nջ�hwj���t��=N9������T�P�	�k�*<�ކ-�/����Hps۠NAl��dX4I�<7B�O��ب=:�T&|z���PL��1Tz��]/;��x�k/�r��;�Ք^r4�Z�SWA�(��rE:�7�e�j�1����A��E|�I�U+��c��ռ���1u��a��pێ�P��Ϋ4���g�9���9��Q4���/')#X��v��5�RL7�re㪀�,��;*�����<�\m��\��G��V�)�h��ňA�T�e��i�2Gp�}��G6p�{��8e մIG��Y��״��	���$�Mm�Jߧ�K�w����:�����嬚栮gPd=
��Y��׾V9d�� �c�c�i=2��p͟of�V�d�r8O��I�u��.�o��.�
��7m��k�'o2eՎ�x{2T�=˔�����K��M�Y}���褜;��h�&%y�:�\Xs�t��J�_F$��V�i;X ��������C�o���P��t �9���P� b+x�s�{`���2���7����v4a����|O��3���%�-��F�/�ۆ����rq�^<A��k�{��)�Ў�c�)�/�/e��S3f�`�ʘ%͔����6�x�LC�G�5���ޭu�/��rfdx)��A���\k\Iщ6���
H��b7���-R��6�o�M{
���Li]�O�t[�Z �:�IWy�s.^��x����9��('��Ĺ��v�ca�&�W���&M&w���qQ�>��]��s@�M�.�U�npX��o`���7����yܺ���w�ڷ^^�T����cs2�`j�]��������v���D������F&�Һ}���y��(|��e'���5{�e@�vjW�}i�9T�uxc�6��WR��T�1ٌ(̶tR�B/\s�V�0��z��X�%Ty�>�����ٱ��d�R������z����Pb���_g%"<�����`mɭ=t�Xh97��{Qd^:���D���2Sy� }�@<t>	��"��1Az,� �%�+�o,���Y;=O�{�����1�R>�������Ǜ$𠬷��y���X��vkW��h�Bm��Z��v�>�]]���E��y!�dQ�쫹���Z[��G��o����>%�x$:y��1�]��j��XC6f����=�zZ=���B�~�b�g����8,��\��sC��r
��-G�A�&>o�����=&k��N��ǹw34a�=���ޓ�A�@9��V�C��`'����#4ܞ5�Į�qm/U-��m���V��^�+��,�c)s���ttR8��zaȻ�c�xZN���ĺ�אS�˽����j(�xR�F3�b2+<���&UZ�����ݻ���%��q��w���=��%1�(>m�K���P�aC��[-Nj!g��j���UjS������Q�j�QA�
�Qс��P�q�v6Pi̾l>BL% �R�>\��f�=Y�#���C@.��#S�*�xU怷H�x�Gd��y�^���L�nlxD��8��7Z{SS@�)s��n�.��V�^�Nv�Se=ه����9s.���8Χn(IGr��z�8��z�S�'��hG-8�+�R�5�n=G�[�"�jK�*U���t��9�r��54����rf���ʋ��*vAo:���Kn	!�#���$�7$�w)(lJ�t���!�y/�,�XK�Ɔ��D�D�JmEA�kp��k��x^^�bжm�-����#�"Д�y�eGRU�.M؎�;�,J=��N�g!w�{$<�f[�J�gL���F	� ���ٯ��E0[u�V�-�CG�����P���`s�E�4s��r_y����L�ؖ{F���e�!�*��Jr,��n��� ���R��50:�MfcF��=k�^�Fm߫�s����鿷ys)��,5�ƾ�Dݱ!���� ��Π�ֹ2�� ��cK������?�@��^�n*��ۡDu�ަL�͒�Pܪom���rs.�tp���3���af�H
8�(���m:��F��.R��
۴�Ա�����u��l��4̬w��#���X�Ź�����؋���Z�8�ɉzD�xf�9�[u��BFP9��NUH�"V?��<���Kߥ^��&N�J���n 	oA�@Z�3fM`b`kS�yn�
�!��+u��th��׬�Mͥ�(���n�78�1��ǆ����w�����ot�-��{� rs�Oob��>P�$A������9�{�Ec���-ݜ}�y�՞���Z2n�Ly����v�~��@��e �8�����Nk��L<����4�?:[��w�ut�C��*Y����:���)T��p�����s4lH����Ȟ��4b07;ɲ5M��:F���dl}�ܞp������A�{�,x���:��>ν؁7ѫ�6�����:8���_7.`�گ��)y��ID{t7.���.ƫ��Q�>��Л�s)h��Q� M���t���6�Y�q%|��������!��=y�n�e�0����t.�2q�#C�N��vnpsJ8P�yf�CT}ϫ��]�:�{+�ެu��0����/m,� c�8o�lzL�qdO�(B
�h&�x�.�xOs��6@HYGw	�sM��`��؃���R���Qv޷}(e�"�{YF� �S�\��^]���[t*�X���s{oX�1ʗjԗF��gN��C�J���"Fķ	�[�d��*os�]�Ly��*�ƕ����%7�D��&Σt�gFPt�@����'l�.�8�m��fb@#��fN*��2��:�o3�V��O�ޝ�-to�ޤ"�ztˡ�~�	�I�S�z���4�Ns#��H8w�����1�\�kA�7�$|+������xq�/C�V�d����Wkv7#V�ۛ(r%Y[l��J�k���[�-r���S�r�ѻf��MF@wT�<���RX���q�'�Q�)p��f�'�%��Υ����M�`����{��.Vx%B�Lh��wVYy�������8V*��)wYr�	<�E���z*v6�G��o�K*�4�&7��X����٫�"Hup�=�V����Z�fhѩ�8�u��]B�s֕9}Jf���)ne8rdi��C�*�$-mt��B�4�#S��p��������؋�
�u��
�1�H��f���m�c5�{;�����g'-�D;��c�>�u�	���n:L1�V�9Ο|�2�6�E]�z�;)���0�.���SM�Vע]�>��Zx��|S��A��y{b���i��i<�
��?M�W=�	���R{���G��ҷz�ɤm��������Qy�Jf�>���b��˚:[
Eh����c˕���"���|����F9�h�wh�Ѥt��4!� �Ţ�/Ց-���2`l��X�!Ĳhழ�}��#X ܐ�lw{$v�!�S;�C���/��MrX���'��P�J;��,���N�=����gk|�J�O^봺������;���e�����F�z�g_
D_Z�����oXV�T%m1�rnG�B^�8���Ѽn�����5�xO�%��[Ӌ�:?e�|���S,p&N,7�f��X
xm7�D��G$Pz]��N�܅��.G�a�1>�o+�:s�g���A�Iv�����iKhTT�Ny�X�l�0}.:2;^h��S���;ܽ��"�g
>�e;߰e}��p�,�~�pe~���;��}�y+A�;�L�k �N����|F��m��0�T[���/,Iُ-�j���W3E�۩tp��9�|��Bl��:ZMx��(�l�Sr��z��Z�f��N���P�4Q��.��b�-.�'�wT�F�"rA��"P9��{;(~Y�T�nT�6=Jw����5��W.�.#����|55h�w��|��A.YM ����7�^�L9qwf�����`�"Hy�U<7�H/�;c��Z��=Ox��"�f�|o��@�hn��Sj �����2��o���:e�yqSD�>��	f�ѷbY]�uj���s{2_X�׋�<ň��ܗ-bC�GI��o<|0�KZ��)-u�,0����U�{��7ȊpbҾ����#u�� -�C�qv'!C:�u.�]�,�Вvp�>��/�|���:����{��#;��ix�M�J�FO��eR�Mc4��t<��<���'H4�}s�3n���-ɵ��|�I
.��}�z>,�=��u���X�u޲vW�R���t,��@rc�����@� �6'c��$]<�Cʯ{��+��0�x��v�m�U�KP�\�Hw:>��ܴf�v�}d䅃e�M0ηvWu�����}/�� 8�.ӫ��ugg�W7�4H�.��a���D�ׯA)�N���c�:q���객q���;m���e�81��uְ:Y�=�ǐa_}�&� �OqS()�w��`T�]>�J]��
g��gp��R��pf�lo���>,�^{s�d[��-񁴎��m�WS1z'o���I{PEf���h#�6$�T@��囜+�v�BOw����&͸+p�>����xX�xT���;�M&(�U
�ӷ��������wD�	��j�!>�o�<εE�(^�|�;}XZ�|7݅�F3�A2d��Ca�;�����>�vNnJ�S��=�5:�{d��c�D�#L��|`G�$�"����~�� /��t,�y<#;.�>�pC�-f�F�d�Zu{uw���|+8\���{�َ�V*3%�t&�@3ob��V?����gH�؞��k��SKPW��������*�v�����[\���Zdw2��6�Bx3���6#���NU��WG�55g��dw¡Q��s6�Z���E�)�}���+.�c+�R�Ӯ�nS�K���9M���Z�"�P�FnS�y��].Q�4�72�Vs���P��E�!��fM�R�L%��1���wyeU7{d�'Ǩ|{GVK9��BT��S��[�w�jΣ�L��A�'�>י���m��iDv;�`�`)0v�;q��s��g�Cښ�\xv�
S.�=��f���`gr�z�/(	�����¼;�i�)oa)���h=w
1z{����#[ l�u)N�W��Sߣkj5���e_8�/&v�ڊ*s�D,#�}$v�a�)dp6���˰�dK���ݳ|Дe���Xdӳ+�`�ON]�8�G�������d��n1�[�Q��[�}K@����W$��[5ā�$,C���s����{ۏ|�Dהq��{�v�́�A�.�\��°I�7����]��w+��<ՙ�'ܻ�(`�/J8�5J����]��ի�1E�|F�<'�!]0N�������P<;e4t�P����M�Ε�O��tش��-�v���z��(�)��X7/Iꢷt�%���W7�|�e�׬�Rr�"���4��7|B��V��#ÂNŭU�(>���njY41�:��n{�LL�c�>�Sc:q�=ケ���{��g��¬ZO�t�7��?;� ����T�CCe�5��;1*n��׎�KL�k��xn�V�w��)z`Ƀ�-�R�N��Ȫb)���(�k�i{��܃�Z߈bG0�UX�s���s�T������R�5�W)�m����&<�]ك|_�*���9@5��H�s���j�5�.���,`%�+��T-H7��qoLs`�Ϩ��@�PD{ޭ@����n�\DY�s�@^�xUO�A�X�'}�uP�暽h��̑=�j�S�1��H��p���*�!����Y]�oh:��I��O;��İfح�ZJ���F�]������od[���|�8��eݞ�,	ˋ�:��4�սj�6�lXu��'Y�b$Mly)]wJ.�|:�v��5�ku;6t�q��_9�n7޴&��ӿ��>�nw�v9���/�Nf`�!�6�7j=���xiu}بk��7��r����cE�h>�H���-42`���/��k�k�>IuLE��{�|���q'�.j�UYݪ�&m�)���W]���>��-{<�ٶm]7.J��LT��O4�]��c�"�2s�;^R���^)h��np�Pznܝ���:J��啫���T�2���齸�v�jfOr8�~�S3�n�1{ʹ�p%�n��o�Ү��.r�u 4Ȍk�J���M̕9���[�w^�άWB�lƛs�3w
�_v��&#�"=�5�z���)��U�=�GX#u}�
�r�S�P����hÇ�v��7�l�k�'��
լ������os�@&(�X����t�x:� �i����-j�!n�)��)�Ey�¼	��zT1��.���NP͵�%e�����Xh�۽��8L�����u�Oo	���dPJ�nM]9���m�ƣx:�:�,�U�*����-�����9�#ai訪���+�|��$s�m�/ ��|s���W6�W��B�A������� �9Ҫ�<'�� ]��o\�����D�ʰ��֗h8Z�E���f��Sl�F�Ýc{9q�5�iAYj����̜�qԘ޵B�h��(Ԝ3������<���-J�}�y%䲷�Ù���$�̧uڠ$ڂ��W*�Aә�S�.�x���EmEN-8;�"m��5�IE,�*����p`��ӹ�Y��Lֱ��:��2��;uQ��`ގ��u�v����i،��Wٙ�3AhqY���4���k&��ŨN��a
kL^Z���C�<�\���G���3/tL�ƌ���Ҷ!EOLJ_]����Jj�q�p!�r�H�f���V��N���t�3�`U��xN5#]����.{G6Oq4����fw��W}��k��~'�!A�'���eZ���k}딵%+MeJ�Y����RR����kQ�����\ڻ��AS�+2q����C�囡T��c1��1%{�� a]]/�;�nmMo7�Q!ېK�/�m�>fR H,���mB ���z�=Q�8��,ݛ�+��Z�yH.�aA��$� bE��	���ί��Y����"�}&�̖����mHe���7�ӼzM����Hӂ�e��hv��j�wRaN�bד���<���wW��J����ܓΫ����w9S��h��L���ND�۾�`���:q{k~��ũߞ]�M�5�;}y����W�{ڒZ.�'�
�@W ��e� ������Z��@�̰�e��xCx����U|-f��6�hP�er��{��:��6})�:ި���r�u�C��c|3�����d���:���Wv��:����k]��Yܱ��F�X����|wx�<s��Sō"�79��+����Cf�o��$�z���+�ߎ:��]o�}�޻�,�s��V�=�Vnc�K���-j�Ֆ�j:���4*\sɆV��KK�Q�sQ�����W��cij-��������[�L�Ҷ�����P��e3r���\s)\¨�m*ֶ�[A��ͳ6�Sp�[Eh�*Qm��5�[Z[k
#�l�qrbefft�ꂙ�-��)m[c�V=9�������%�w�kKVfC�JQ]�\���`����;��(�2[�m��eZZ��W0ŕ31�6��mZ[Yr���.9AF��&[-lܦ-G��iE��[&V�3�+R�ce�X��k[m-��ŵ��mTic.���rڴ�e�qE�[QM���Z���b-��m9
�����J��-�Rhu���h���Atu�2܉�wN�X�^TM�2��Y���V��:u�^���BU�������2?��,�/��~���IV��e:syI�}��W�v'��J��(
p�VX�?K�}��C+�j疯{���uƣ�ׂ��b�BS�ϨuVت����\�^�%}=�V�ܬ�rQa��ޓ2Wk9,`�u+�,��ņ���Uz�/���W5�v�A�T"��u�~y�?X�����yf��T��ai�쭒�TnCԮe�����v�܈���*
jĸ�P�uv�x��G��	�v7��k�ۀ狖:���DT��©/M�A`���ב�5��v|d��qf|o<���L��xmhW����`x�\��+�2��c���\=ב��x+�f^�I��O[7}�ռ��~�:G;�u{qzGǸ���ë,�Zͻ�TN��g�����W�+��e��$�YC3ߖ�P)�����f�;M�C��	����� Ǽrd�:��s��eF� wN��FL[�m�yW�2���l�I�b1�p��z�[z"&ٸ�t̟��sg NM�%�j���>9|�С��2��^11{>�;���k�HU�%=R��+�L�PW�����2��oX�����ő�'��M.��蝊�t�A�J��+>�Sc<+ʮɔ�;����-�&V�{����L��ex�E��~���u�O��;+����P����6ұ%�v�XB��P���i��ɝY���t���͋�pA�gp/�W`g���j���*Pl0|(݇/��(���+��'	�~~ `7�ֽ3�Ś�>��Ǝ;��Z���Ϩ,%��{/1.'izNI�Ńu_X��ć8뿥ܖ]XQ�wT�f�+��'�s#\���a9E۬ʇ�ƗC6ܱ���L�&
���n���ww��%"7_S�%��%�e�2V�}���U%��*XU�b��P̎���xUu�V_7il2��e���YE��혲�є�Pt�?؇`�?c��9��J=�y$�CD�����6oO1:)S9Z7N��Xn��Z�G�w�2-�k�]��\�uX�gX�����:��߉�������x����tchS~K��� ���� v"?"��X���i�K��h���
b�]ōr����j��K}/Z��`��V���`���D�P���ɻ���~���V/��~�K(!<2�A���ן>"��wJWd�ºyZna�]�n�Q�rá���X���b��EA��>���vgtq�_H,��߲ތ>��GW}����u��J��ϧ���uTm7/+����Z4z� pV_�&�����!��>�ٶ�z3U���,~R#�tP�}�]{�̻�y��xl����2���w��}":��""�4|����c�׭`UUy��"��?�V{��&�$��䏧�����#����B��wY^e<������d���@���)��\j��y���>��4��Z8�Q��o�5؅ Έ]gS��������j�ǹ�1����/1�59�ގ�2r�U�y��o��.a0�M��` �����h��I�H{�ɔ��`w����*���+�\�ML0(+.E�j�}'���^���<�ThVT���?",:=aT0���)���W��$�o<{�:���7�ޞ��d^rR�+��ټ�������/;��-��ZC��t���8���s���nY�Ȣ���뭺�N�"����(���i��֛�oo��x�uQ���]e3���>B���T����)ގ
����`U7�<`�(:֨�d5�����g`]�3f�q�6^�Ϳ�g`ud��t�(�Kuw�w[kԆKO͙�������ތ;^�{�T?�+h˃��)��������uq�#D��*��}�6�#H�v������yr�������ٺ<�8��]�&Q ��W���`�1�^Q�� :�!R��'��~�C`�#<�:�Y���rf<����NԻ�����3KưkR�-�'��k��R��A�}��*�Iل+�vΆ�m���{6�%(�P�P 8����Z*o�^�Z<7���8V���?����dj�/�v�_Ͱ~��f��m��=u�l6��C�'�����Wxrr
�{f��Y,w\����������|ge���e87�2������d(��BZ�C�w�-p��=��;�4�Q����BP������׃o�����֕�źL"���Ĺ�����`��� H��|e��;	���~�:�{��^�ַ���_8���:��]���U��݅2�P9c���_�����yl�J��:x�cڠ�0�	��W^�n��.���m�hH�ރ���9Z�!]f,��fJ�%��u+��LP~�]׮�%�Wh(�E!߮Vz�K�tg	�bK�4Ⱦ�N���S�m-/w����e�,U��_b�v�\���+�*
jık�ey�jYTٛ��K�'���@����j9��i�y�/�-��\��tޢ-$�����u�� q�J��oK�D��]G\ǚ��9�"�y�9(�2D�oA1r�ōgt@int��z���ӿ/�)g�ykNV6d����B,�uv�Y�<���+6�R��˛�bQ��d���׃��Y�9/:��}=�v���~�I�$O���pB��De�WW��"ǯh5:%��s=��]�}^~|�W�~���ױ^R�c�t#��Tt�P����α�&�e��V
��ںۖ��
~,�Y�(r�u`�1軑r�_���a�]��|�>%X��8�ϮS�r�������Y���,�dk����*P����~�G��̤E6=tʮ���%�V��m���C4UM����B�K�'���?
�0e��z��j��l�,���Cu��,bdp�S]]��Z�\}�m�������.7���jq-ԧ/���T�6�*��|(�v�7�~���$��-���t�b{JL{J�����xGI^��}:�ˍD2[�[��P5��G�֎�y�rW-��M��z6-�mE�T��l���a�N&��.t���\���;	/cr+lp����}���Pf�`h㽑d�_�h&��(�Y�����Z��pW���z��ј���L����u<��]�u{���}yǙ����������_yJ����Lɂ����7�CIF�^�b�}R���]�2S���U%��6o+�ͱ�r����_�Hȗy!��`��;kA"Q�_X:q^˙n���EC���6���m�q���n��t���A.��cE]�ў�����
A`����O��~�J�dʀ0���6��_]�d�e�Z[��H#\����D��s�+��
���GS�k~w�Z�����wȺ�q���l���/mz���({=1�ϫ�X�#B����/8�*�i�oO�f��U��e�~��:���T��y���U�˫��W��i��w�����+���x��)��Q�N+�DX����R�״E,
�F׫���%�_ժ�����ﰓ'q�����/���Ǹ,iq�
�$r��+������&�ۊ�/�Z1���n�ˀ��b8���{�+��O�ܾ�~u{��z}��&�]F���*{j��˼�m���1WBS��h�+ӭh��?t�v������.��h���FU[�x_ޡ��U,Y4׶{]��L�8?pS��+r��]:�vt.�UV+��/6��=M�/H���6��~�5K��7>X3��]m	)��� C��8��^{���ȩ
Te��	�PU}aT0���*��
���vwVH�gH������}TC�����`'�J��)ҩ[.wKn�t�v�F��F�v}u�ܲ+��E����"�S��D��{�� ��h�����W�G��Uf ^T5c�U�"�<���T�p��pSVE�C	�q3b�$f�|���U""�V�X�q��lfYt*Xp�]C�x`�|�(��"�V�wZt;�*N�H�K����)W�Ś/2�&<,��(�WX�	5.��I��G��{Q_���څ��)��'p$]Fx�i�*)j�$�	�֧7�-�+���)7�l�ïP�φ|a�����ї(�*�7=WY\=�.���z�y0�[�*9T �T�V�}�k�=����vĥ��p+����{��^�G�
��T���#.T7��=ck�	�]mi�{�+��7.�B�[B���79zfU\Ь��B>P�ə�>���,��m��������!� &F�.��wo�����\���O��s����=�D�q���Ϋۨ��� �];7��0��#,�.�g�-���(���h�~��ұ3�����qz(:
(�{�� ?�wƅI#�t�±��z�7}F��I��c4>�Q���S�������N����?S���b�W���*�#!U���{��+�K'��51�t[����e���fa����w��Y�}-?se�Sǯ
��n6VoX��71�+{z<�(d�]^o;GXD[Gi�e�x[���`
�������v:���?���b���T�7G&Ƌ2C��K�wpWO�|]4â���nsH{�� ���5���]K5=��~�b�����XH��l�r�$,���V�z����u�!�ciԯ�ۧ�F��c�^e�K��|<GٕV��ԁ�,�>$X��d�X��x,ӡ����ދ��2>JumS�!�ҷB��ܕ�!�n�ɡ`=pP��]�^w�J4�ѫ,z���C|�P�;���Q��W��0u�~DT�<�n��1r������_;�7�f�(z� ���׃6f:���u�~����>��u����^e.Ռ� �)�qџ���7���������D��K\H���|�
��x�W��YP����>�s��t��~�{�V��L3mT���9[��R�r���bb�ߑԞ����N^غ��dv[�(����i��y��+u���}.��|?��ʣ����YJ���ե_:�ְo�x�%�Gj=La�co,Ye��:i��e�c(�ޠ޹��7�S��0�rD�OZqA�5=�e���`8� �>N��2֐Y�����/w��#;ۃZ����ے�}�����LZ���qG�m4�BWw=���,u��������S��ICt�gfn��;p��FR���6��:o�i�駲 M�i�1,�9o�]�pT[�ݺv���>+X��C~���^])Ώ�ٞʬ{H�Zr�Nv'g,�C��1��l3���A����e�w
=tkѸ����V"V����F����CU��`_� [X�GȾ�#-���=ǈ5��Oc���'�6-|�������xS��oHf�vR� ��Be�>�$J���v��^(�>����n��P�����7��TQbs\�Z��삇qb��L<;7���^i�v�'c;�]��.�^qG���a�G����n��by�*�b��}s�3-M�̻]b�k4�ۈ���YS�wo 3�U�}~�ǒY�ѳ���"����ڟ���5�/MYə���e���^����:���#�R�%�	.�谛vr�u�n�;����͵ȭ��x��mJB� ������^ aj
��;ςdZ��yY��V+a7�. ���[�k�5fS�i�gZF+k*�eT
߭��u��;N_#V�7)��K8m캽'�r�IIV&�wF����]d�{7q����4�-����������'�U��!��Y�Q�g,���,r
; �mM����ݺ1�v�A6n�lՂZxƹC2�}׎��/_�ƟR\hu������h��,՜�w͠�mV)9��9:�m��R(�ݾs-֧�����{��}���qvJ��lX�� 6a?qs�XY�B��U�����f<G�T��e#8i$ב��sin(9t2��27���Փo(z����\+�u|m�����G]gb�L�W}^"�ڢ��c�x֫q>�M��܋�j�}Fc���c�hSz*�,��U-{��V��4Ե���{W��A�]L��hP��n�L�WmhT�Ij���-Z�˅��ܦ�m�#5�[[j4ej�K�Ĩ���X�mJq���+�pJ���Q�WmoW1�Kbnarܶ��.R�\e�"c[u��A��7(�˙Gq��m
�%LA�6�V�f\L�r��iZ�kKF�ؕ���ىG)Th��JX�j+�X�J�̭V��բ%�51��Q�,�e��&�UQQ+X�lm�)�an8��i\��m�����L��+F���i�m�"�iF�ѨѥTj�ƨ��G#�K[ˑ�����D�8�cJT�ib��JֹqLZ�\̴���Yj�U��Ѷ���r%�t����s��i�}o=U��2��"U7+U����Ћ�G��go3]����U��al�~�kZ_��=�9�%��x��i���i����I����_�r$��x ���$�W�i�����n��?�{_�~�{%��~��t�\qbMFF֛� }���,'��n| d,_
��AWAn~ή�9]Zg�߽�;?d��D(G�R��C�y�R_ΕXe��G�复z-��t�����㦍���f}سX7S�c�W_<O����yę������`�:�c�T$?:���/iѫ�oT�-[���;��>�T�Wi>�N����CL��m���x��S}~�Y;.>m�$*k#��}r��������U{%���R��i��xn� ��G�h.Rt��P4'ֈ�)�)��?Q�{j�J������C���I�9��?g /�S�pxu��#<q\?L�4Q�t��Qf׳�EŪ6���͕���f��s7��sWQ:�ӈ)1���c���g�R.jz�����|2���l���ݣ�7��7��*E�1�t�>3��ܴh�C�Z�e�l��@��ɜr��{x�i���Qyv��֮�t@\n�8~�ߺϲ�Ed�WBΉ��ό.�^�R��(}n
w��Ϭ��,�o^-	{vN�����6�����~����{=1��,���G�7O_t�ah��W�*�v<`dE��e{+l�U.y/)}×_L����G�ag���]�.�h5���̡o�ѝgG�$���n��޷����X�cB��t4Feܠ;�ۺ�b���Mmvq��lJg�O������像^xt~-��+>Y�����x���X8�)y��Ɯ�}��m�y�C�w]^�b��,r�nx{�.Ļ�\�n�Hj��,z�u���>?a�������Sن����uܹ�Du�x*]
U�_�]��*��`�0]?\�"����Z~�_��t��EeF*]��Q�>�>�ZE���{�J��+�����Ff������}밼ށ��]ҲKǖu�'f2j4�r#Y�::�֐"����v�5(�C�������鯧���r{)��|�q�����˲�eRxקF�ŕ�f�+G�+�"�[��(���Ȼ��~�R���W/w�rt�ԯ����Z�ʬρ���ʝ��X��1��ZI<@?zJ��4�}�*�$Ix:�d����ϖx���.;��;i���3�~�S�xQ�6�_���F������u�C�/����ok�D�}캡%�m�0�<���R��?a�������ɇ-���Z�\�Q��k޹l���p�Du��[��u����+��ܼr���MN9�jz��dz���2�!�����c߳>5�����c|f���:��Jq����#�Cdnq��N�6?X��\�^~�.�����߷���u�~�m|����_���|� �ܧ�����-e�o	���Ԛ�V^YsF20�����6FuE��"�T��2�xE��Vw?���`�y�5vQ�y=]S_���7��&gp�R�W�Z� �pjo$�"����8��7T�	`}��+l�$�XD��ֆ����=G�ҥC�w4Y�6�c�I�W�sܕ�@���󁇴����4E^�ԫ�i�$��u;�{/>���E��^�D?B�㐪��!��9/%��X:v�������g�w��tEW?��B�UPSl�2�Q����=w��R��wZ�]v��%��T9p�O�Z������q�/>����6%	>�*�*���=X���.��䱃mԯ�����:��w)����e���
��W�X���Ia|ɂ����u��Tܗ���EF�	.��D�v�	��]�:e|�����~��B�O�`���+�.��M��EUHT�G[���+�m6#}�Y�A�<d����N���U�k�H�諸5��*�Y�وF���O�G����㈱��U��&��@���"���QV�8��\ޙCYͷ���Ճ��-`�^�M�����'Ft��=|���o^BV��Y�͏��2=�^H�ü�K�ɕ�;D�P�z����s������tQ����*�M�< �)����sϥ����yf
k�^�����P�j��-g�ڨ¿W��E�\T0Y�����K^7�kו���X��r����3�G��XUen
b:E��׷v$͏*�e�h�u���_�U�����6���a�嬽}u���)WS��}G�{c��V����T����2��Kd�^�A�;�)��&�����~{�B�=����ֿ�zN�����,�y���e'I�y��f�=E\���PJ䱁2�
Ǭ_�
�LV�l'@�����>�(��յ����#���T�C�x����N�(6/E��<�ؿx^?6C~�����,ѱ�m�/���u�
ۦ����\��Tcft���>��Wi_��Eq��e��mPks<u���K�k��w�U}����T�;�7[��Mn��+ݢ�.C��]E$n��C�4	�K��>�~X�:'v�ݻ�������z�x���w�ђ'.�1H(���k=�"�k{��y�`N��&f�}]:�֋����n�9oH�Z�_�)�Y.������:"_�CL��m�c��}�wn�ͽ��Bۓ��DO�IbU��_U�U��6��`͙)��}�{ơU=E���z���m�@�D,����4D��!��u^��D�N��6O�4�7�c�;�u�\�5FZ����������2�u�+*1���6UM~sЙ�>�c�f��f��j�u���ΗX��O��]�k���$��8��W��hǒ_�LVP�E���u�w�����7�/�h����˩U�{{�u��lϽ�D��B�p��D���[<OɳgM���h�{*܅_��C 8�'|iY�eW�|bE1��O<�d��h��y��BU�0!gn�]G��i`�>��e�^��Y����J?I}N�z��V�n���y��8����*�Ȯ.�@��q���<M�g�D�*W�<�\����ؽ�~%�����Ɋ7^�?/{���ev�>�*܌��szf�z]��g%�{�����^.N��s�Yݶ#��>܂P����N�������ꖍ������C��;������/#*����U.�.��SY�'Ul���~4Վf^���*��_�:�[�I֞��^&�H荫��5@3bU�j�|5g�|~�l��,*�j��Ǿ\O�B�hۡ|��j��V�ߩ]�:«�U#����n��̨,�H]n1���xkr�3���P���Ͻ}��Y��O��`9������/���;���dQv+� ~��Z2���N�hCx�C�~�LN��~����3s�U���U� ��ˬ(��,ώ
�r)ɞ�K�۔*�5~w+ ��_�i��=V��Z��>P\_HX�R<.Uҿx�G���<�g�ƨf���X�HUyU�u�1g_yX��y������wF�]�ݨ&�V�f��<~��y��ՙ[�h�Py���m�e�/�T �l[�̲R��5�ˌƼQ�{fL0t��+�a�TX��C�MW�ﲖʞ����J}nM'�-��q�Q_C����f��wx�S���r};����,�^�{s*������D����%�Ҽ�ML���j����%��?O/s�f���φ�7�V�(������fo������Fڏ�I�צx�O��
���}�����G�����h�0~^���&��/8���˙f�A�_�ph��΋�enS���x�2�v��f�MѪ!�D*�.m
˞hmН�q	n�v{�$|5�Ӻ_@�����O㓱/��L��DoY�Ϳ�qE5�,�q�x����b�Y�������`$9j�߲g�L�-Pڟ�����1{�.�B����ٟ}-�x*���!z*�)�z�]}x��w�J<�������mܮZG!�%��A�7����c���CT[�Q2Ż��&�]`�T��z�o��vc��e��u+�v���MJ�k:��\��9�''^<����z�y�CH��:����TW$z���ʅ��8�&ނz�V��W[ �,�Ĺl����,���S5������rk�&S���ؚ3�Y�C?�}_UWn��=�h��9�)��w<�2?���S�ק�L�ВƲ`�/���4���^/���d�^>wO��>��F��x��,�:�.DE���;����^ؠ=Z*Ȗ�J}*±�xH�钍`���%����T���UG��v]P�b�r A
���g���B�z���O�SY���<��%͑��쬃����u�+��Ћ(�x#.�����״"�x���Ĥ����ϰi1^��A^��v��Xa�, :�*'�r����r����6����Kz����0��	����?s��o��!Nǽ9^`��0����jʬ6�l8+���c�*�\�W����Ws�sn���m^��y���)V�b������xS�w^橨��Y\�w(�`�	�}�o��{r����H"��\1c��#,���� ����+>^��la:���^���ʊS�}P���og�UE��8�����U�s�6�\�#�A��#||{e���;`���P�9�r�'�bC;&N�ܯ�'�5 i����������u�!����(Д]����(*��v:��� �b�(UJb�w�ueg�^��I�������~����Dz�*|!�v�K�:T����u�y�bJ)�`$UP���Ə�������,�]L��Ii�E�95r��ؿ���]�����}�Y�0ڠ�!�㿺yP1t�r�I�o�Oӓ�oU��go����_]י0CL����<��S���9G�	��"J��%X�n��@�=#`;��͇֝.X+�?Hi,���+n�
�P�X��K���꼴���C뭛�_^�޹�|����Y*��^��1��V~d�� x�
³>�s�2�T���R
z�e`q�m������̓R:N��� rc�6�Vi;����������e|h|�.�+|}�Xt�Rt^`Vo�L@^��0�>����a�/(�G��°��~�0+1'� (�`T��@Ć[��'�O-��y��}����)
ô���i!��d�'�$�*,�J�2|�;̂�{�o_a���Ă�l���T�����|ʟ"�~�����rϙ1���!���7~�����(ڂ���h���N]�/�{iS��N��%3b�/A��x,[Y�]m4�
�rƂL.R�z��V�Evbxn�J���c׮�C$S��vp�;$��71L�!�+n�t��Y��i�]V`;gh��:#>��G&cݜ�U��k	�YrC����k��o4������ӱ���ޚ` ��~�G�Nx^����7yIy����0���X���}Aav�J*pr6��7�{�C��Jkm�f�U5�4��Vmjz}���ۂ�0C]��2��n�܎)�}(
;E�ۙ/r�m��D�b-��k�{*>���X�����J��vJ�I�����djs�΂�W#��\�d�n�K��^kf�ۄ�'�a)>ȭ��R�S�I���k�N��͞ e��==4�<}5l�Mu`�\��b;y����6��B^i�;ٱj�ʬ}�v�ø���/jwIֽ��t/A�ɜ74q�`����G�=;���żt�cw�xE^��6�mm)��{<����x<�Ѥ�iN��3��<w���ڐ^�QZ/�E���Q2�K2�kW}g���\*���hɼ��/r��ϥ�p�	�7E�x�M��QUxW�3u���H�3�Wb[��RӪk�/���b8��|U\�G7p��M�ٳKYM��C�M����5z^s��/�����qVQ�����N�,�zc'��m���V)���9SpK)^e3aE7�trE�F��aj�k�A��e��sec۫�b+�Ľ4�r6��`�H{�7î��CG-�oU��5=ꯧ{o��{mٹ�FFB��LHs��ҕ��&��vnXի�oo\>��a�V{��5F^�Q�iӻ��L���w����
@��)e��w��W ����&���{�RR�Tþ˭�{�)��=B�W	�%vVP�����ب[V�+2����eˬ[�<�'^T��l�yyr�{��̥gb����r[��]���:��NP�lN�Cmja-{10q���#xW�P�PvF�Jn�v&��Ɏ!L�6l�;h@���$�Mw�~w����������|hX��V֞8��[iJ6����3��V��[jTZ�J[U��5�eJ���QLr8-��օ��6�Z"�e��ml-*��4��q�,�A-��j����UZ�L*W)J�V�Ҕq�V�F�m���nS1�5�����bckm���c,V�)��j��Uj�j�31G,kV�֖�-��V���mB�"�Զ�Q�J[[-`���Q�j*���QF�fcqDq�\Ụ��֖�s331��Zֵr�`�0�e��Xڎ[�W)M�qU(�kZ5(�ikD�6��Q-��ڶ�mV����B�:P�Kۿ��w�]���$�Tە���c�cv\��Ф���k�4ȶ����o��������=��Q�Aez��PR����d�1�4�0��9�B�[g�5���3�J���wζ)<@��L��T��Y>�Ê�Iՠ�q�'������xo�~�߿~���������8��c~9�I
�y�靲T��Lu�!��Lg��g2Në5��+:d���̕:��&�����񿼻�}����~����}HV3�����Y}܇�����f ~�R�J���T醤=����ɉ:�b,5�O�d��Aa�/�μ�yח�����o}���w���Ì*wI��g�u嚀��7�!�^�3�!X=Xs)�i��OIĨ�}�!��&8ϭ
A�I�(���݆05G��:��"�;�?� ��U���&"��*x�w�MH,�2�g������R
t�Ɉ
)�<a��d��bx��=�(Ì+��S�,��̕�9���yz3z�w��s�_��)=I�e�����l�X~T+:�&$|ξ��
,������^�,8�����8�����/�\Cĕ����~w�xo�w����{��x�3�N�܇�s ��
�C~��Ag���*J��S�Y�Ϭ3�B��:���I �uMa�:@Qg[d��f$���}�T������y�s�����ߵ���Ă�凨k:�Ɉvr�"�XT����:H,*r�Xz¦�@��g���j��%E=@�����B���������y�S���z�����~߃�v��t����S�O�=}C)���k��ğ�����V�uE�S�RbACԙl�~N�٩!����%@QO���]�ϸ��>���{������*v��=�|~���
���g}ag�J�:6������T���C��B�:�@Ԃ�������-���e�TE{��T7�����mW�|�b;���s)�ֺۆ��t:a{�\FE4�q���)	��q՜mEzi�\��6��g9&��d3u!��jf�N2-�R�V�0��f�jt���!��﷾{���l=a���$7�Lg����j����@뾰��2u�ÿ����&0�i�a�i��J��w�����g�L�!Xc�;�g�{ï�s������:H(yLf��1E�,J��b�T�l��,�q�0<��O���LE"�
§�Y��ä��Sg�7�(��H/���ݷ��~��׾{���v������8�P:��R)
�:a��Aed�ԝ���>�QH)��}u��H9{���t��1�Rb�g�e��'��޾�_9Ǿ�￾�ߓIR
}������u>�!R&~�&��T?ZT
��Vw<�bv��9a�Vö��)���W���}����ydѓ�T������]9g-��k�N?����M�6���Ă�_���1E�&'��d�bA�C�V�H)�?QI��%a������O�;:����2i�}s���+3�|y�̿�n�Ϻ�ϸ���� ����CS�J���T�
��_��!P�<�3�� ��Z1�����
kf'|� ԃ��~N0�O6�I��r��9�{�6�߿������*}�~h$�}E�흦$���O̚�����bt�Rv}C�H=�:���0�R�{��I�!��5�P����q*����ԚN��W_
��T�v��c���� jVz�;�&�(�i�2j|�J���0��2bx��1 ����3�%@��0S�
��_i
�2z�s�K�O�|g��^���߽�/�k�W{��R;a��ֲ~�)��2|ʂ��Hs,8�w��X��q�!�
)�OY�a��H;a���a��H~��d"��,�y�6�`��_*�믿z�C�J�����!�Aea�Tw��?0�[E�ͤ~�rMN$��*? V���!_>��q:H(u<��kɌ�I�9�v}�uq�����a�,��w�H���d�Y��Z���-�y �s3HK�k7��㬻Ҳ��ˡ+h�+3�ۧܜǘ��`c�қweΫ�MZ��+� Zݒm�;ӿj��拓B��韟;��N�j/I �N0�,�z�x{a�>B��hv_rt�Xc�p���YQa{��Xy��5 �2i�5��T������g��v{����O�s�����n�T�uCXt��X�H,���^XqH)�����,M����}C��A@�S�ʪLH,3�,����r�H>��&HOw������뾻��^CR�Hq	��~Hz�2q�󔓉<f���$���q����V~d����$1*����E]���3>�_]|hC���>BT�& T��_�Ì*\�!�J�2^�0�!�J����E ����[�!X~g�SY�'�H/]�d��%T.��:������~��}���<@�>��ă큿]aY�1 ��Xx��T��ë�MH)?c�V,�z�����Vu�v}a�Aa�ܢ�}@Ău;����w���������V��g���t�\ar�g̕�i�`T���e �Cͤ���I� �����!R
z2|���I-�|������w�s����߾��98�P1>;ܜT� �e��T���=�ă�����a��T��-���J��ɉ�N!�bAN�;<�:���5�{�d�5 �[Ϯ����z�}�������ɩ��2�@�'��.�Hs)��8�jAa��c>g�c'S�1 ����;�
A��Qa�8°��(x���11 ��J�~�߿��s:�HH,��2N��V>!��Or��钧*�������8�A�'��g��=�5 ����_�H)���1 �w�������}�~����Y+z���iH)<B�:�퓤�ü���� ~��X_h�W�:a��y?Y5��T���1��n�=���߽�:a��U���u�/Wx>��NW�v�r0y�w6{�CW��P�~6��8Gb���ve��N�(�*��q�j�K�3�[RvTq�(�Aew`�ǚ���t�:���n�C56�9���Z���!N�?wߜ����	�����.��*)30��,��w@�c�d1 �y��⤨
wl�2�IY�%H>��9=���T?Ph|*�������Bg��X��6�O�h��
��~��������
È~q����S����_̟e1%O(��:�&�ԅ���R
xw@�q�!�:<�H)�z�O�ys��9��~�߹��v�R�]�=a��Vw>�bIY��s��P�o^�ӏh�^��Y7{�|a��Ne&!Y���W�����*oW�Y������<���I�W�����<����t�Ld� �~O���R
d󬇬� ��咱g��9�t�RT+�w�퓤te�w@Ę�a�/�Y1�0����ٝ�\���{���� k?2T>���_8ã�5!�`+�!Xce;?P1 ����?=$�*,�ى�'�0X{���Lg�Q��R�b��%@s�o}޽�����z��;�����&2����0*A���ɬ<aRt�H,�'��@QN W~��jAO��}�+'�}f��;L`uˌ���2}�U\ ��b������M���k�?����vO���*!m ��z�3TR
|��d:H(uL�0��W��C�+=��$�<M�C^�P1��8ə�!_ٽ�繟���9�w�����̡�ﰚ�2T�UU �9��H>ӽ�k3��m�$k��������X|�H,�l�풱g�PԂ����]Ϗ~���ݽy��x�z��Ɉ
/���S�P1�J�\����L8°:�ư+8�QH�����w�����7�3��a��ۤ���N�I�TX{���߹�s]����?oЩ����m1 �@�3��{��I�r�SY�9�b,�2�"��*AH6��Ma�
���1 ��nPPS��8�@�=�޳�����ӹ��n��'��=�ʵ
;���Au�;�0�E�S��K�#��DmwL���}�fͽ{���Ƭ��N��8�/�2��	�&�[؉�2�C%	jP����ѿ������[s���?~�=r��x�+�&�2'�c+%x�̧��S��,>f�l:����P����Y�1�����R�E�$���a�a���z��~��}���9�3�P�%~����(���^��1���c=d�>���°��O���VVJ�3�b�AOXz[1�Ƥ4���!Xq��οs$ԂΑ���h��}�Ͼ��)�
(SXz�H/Y`gVJś��|ä���
��û�5�O��c��Xc�)�LaXVOY���}����Q����������ǀ~He��w�Cr��:N���AHd�2x��|�w�LN�8��y�Rt��L>���l���T��݆"��*|�~C���ޮ~��s�u՚Ɍ5�~��Ă����t�����Y��!��aY<�rB�F��|d�1�sl1�2W�N��Z)<@��L��T��Y>�Ê�I���:8y���>��)��MM@QH/ܿ���
��a��_{��AB�ӜΙ�%@QN��Rc�1���x��s$�cVk'_nY�%G�sϞ��7?}�>����T����,5��P;K�!Xz�&	 ����8� (����&��1�ق�}�V.��;a�AC��(c7�&$�i���>�����s�.������ ���:�a�
���c���Y�
/��o����ۼ�{y��>���@{h_����{{�%,m��ٯ
�luEb��Sυ-ϻC����*^�z�n��Z1����ڸ ?x�z� ����x|~�� (TЮ������j�i���VY4�qV����y��'_m4HW���r�p�xU��x<th��Ю��U�OՄ��T��c.X4�0�9L�[[]Ӓ��[iU��X�Jȭ1A;Q�������E����J����.��"�PE�V%�y��������0�G����J3C�+����B�DSf�*U�^'�~�������A=�Y��7txCmۣA;��;2K��4�|�}t_�:�o��z+{���K������ի(?R�oF��\?w��[�Ev2)��ԑFV?g���U�P�p6A�Ue}�V���Yp�*P�ˡ�"�U����6�F�*��
r�vm�/���?~�{x﷡��?`�`���ou��[qExO*?Y�u�,J+;]�ߥ�f/�ْ^��N��/�C;�y�N,��Q�W^�AwB�e�f���aA0ie+)��w�^�8�ds�n�^+�/�Sw�w�`ߞU�B^![e�Q_NnQ�'ƃ>�'�����<��ˋ��B�W�a�ꨀcʄ|��C�D*��{^�D�Vz�����ؓI����em�lY��'�6�IBb\�v��)+�8;�:�:�l�S�޽'k�l�(�oD��&�^�o��
s��*#���SI�����i���_��~�9逬Ϋi�KϞ���+���\2
v�ZD%ʓ��#6;���(w���Y��h�eY��,�A^R�n^��Mu?I���梯v[�b����qF��7�`:[Ͳ2�����=`�4�L��L�����~�����p<0A�9dx����`���ߤ�P�[[�0�SO�{J�z�|^n}��tWRϬ�]b�h�h$B!w����P�]�9!�W�+�c��C��?:R�;�TC���/E[f���~{/5&�"Բ��D��e���|!���.2X͵Aӗ��זs��S���9�>'$$ax*��>3��}�ׄ�r_�a�Wx��cNu�[_B�T��+(���W�ju:%���%��¢]~�z
I�]_
�_��hr�>b���L�|�X�>��:�}'
�����Ęn��!��wz�<���tH�S)����V�����(�μ0��/�k�G0MgB�V�*4�oq�ZY{,�z�0�����*����lV!�5߀� ����2��~�D(P���KB=��Ci�$i�(ӽGGp�jO|�x��c:�(�w�XU%�U��#߳������~��Βa�ߎ���K���|�m��,]��e^��/!�����y���v�e�����}�I��z�!Y�!�oP�a�t\d�t'ޑ�x�e.�.�b�ǜ�����|����zJ>�CC4w��͞��P��YpQ�6��5�+������v\�(�巠�1(�#�RF{�f��,��r�x�l�V��ᵃnY�>�Д�^���:b]$:�K�~�L�Az<r*��ղ`��yqL�ڨ�-�LBf�Y,J^�^���ΰ��0rX��
�c��J���Xv(U:�P��:��{O҈�J����RX�&[��^:xwE��Ǫ,�us�+��u'�"p&�17�W�����Zpp姽z�&�F��M��O}�5�A��^�BbU9ԥ�����9���л�W�+Yv�	g��ӗ�o��}��|+/r�ֽ'�)�'�rZ~�ܳ���7��ɷ�g��e,�����G��S�U��tg-���;��PWm_��:�ϥ�b�Pi�s��EyD,�tq��}���Wr_S�Vx�>wT��Ԉ'�)�ڇ����{'�Y�6��̡6ұt<���ɂ�6D���ЁTGXF�}���=�u���4���y�r��R�@T0V��y!��Օ��ӧu5ї��$z�:�ΜW�;�ox�x�E`-�tW��L__��+��SO��WJKU�]&Ȃ�c٩/z�1�#U���c�ղ�Ք��j��S΍�p�fz��T.�^W��Icj�;bTv;�����3�~���
�����B�#��2F������י����#�WU��5C�!�\2��o�
�������;5v�G�5*��xy��$�r_���Pc"�NU˦d{-��j���l5�u^^�k���v�Í��m�l�z���&�W�=z�)M��GPt3v㙪]\l۾:ٓ�}�UW�Ļ�=��K��<�e�ڷ}�o멐�� ��PA*���9���}Ϙ�D�:��x�=+��y��~0Q�S�Q8K�A�
ҴnƟzI��J�`�Ugz�P��#��O>s����8;
�k�$c�Ns�ev\e�������8�a�gC��U�(��@V�EH�a��%�9O�'�VK�s-UWU�au��u,W�\]�3�~�x�z�a�����a��:��r���i��Qf�**�l����VPx�w��W�Y���thIj��C�Y�03�������:���N�u{�����#�#-ߠ3>�bW�,�ь��h�z���E6��	u,݊���1[�W�Ef�yoD*���r��>t���z��:�.��}e�+=b����X�k�3�����z]�B��VLk�) ���Ӛ+:��Wf�;�Ӯ{
�9(S��LA��h3i2�lWm��j$Q�)I�o��K��@�����Ї>��I�3�w��.k���q�k�r�ff�.eYܣJB-���L*ǭ��,�]��Z��[��r(0,Xp<uܵ�mn��34D�T|�m������mM�͇J5�C�|�m��;G5f��$��n��y�Y͗=�I`C�Z���)Et�$��V����]6�Κ�l�{jpgw�s	2t`B5�wf-;/L�5|Ft���c^�����CP*sU�&u�{yR(٣�+�~����7x&���U6�e�ˤ��1�L�w2���uT��,r����9%݅Pn�G�{�y�楓�]��n�>�j<�^4��r��� ���M��k�K��O��I��-�9}��t��c�Σz� �{KvP����-�.t��V�fA2Ԋi�u��ן�2�f��ATx`p��nѮ)���⺁|���&_Q�yf� F�f�W��m1ۮu��1����"4����θ�O�����?>.˕�yF����+e<�X�Ml���V�2�4�!Vsl��7����0|vmffS��W��L�c\��U�d�M�m�w1f�k"n�����+*:�pZI�'O�������~>~�c��e��v���"b玗SP�b5� ��$�^η2���ې51��W�*�H����o�Qː���a�i����JL�8zs��)���0�Lo'��˓�33È<��tz z��ܚ�MdD)�7���A�O�7bΓ}O����7�i��������6�m��g���6$gC��"��3�yZ�����K�;j�*�N��3Qww��!���)��gi�<��<����T�<gq6k���g�N|�I�4�X�����	�:'q�h�E��sۢJ%�`�����c#5�����G�`�=j &���F�-�J{,!�'+;>)K;�V�оW)�Q���$���e��0`�]<vC��6�o���k�� `8  ���Dp����D������Pjf\��f6R���ƫ���6�Ef[m2؋mp��Tb��������f*V6����i�P�Aau.�Lqh���p������B�B���b"�s*��5�1[ne����ZZʪ"�E3\\H�V%neͲ�����.�T���TnaS"��w��E���Z�6�Z
)�[m,�8��n�G6�DDL�����m�Cp��\µ�5�ۙ1Ƹ��SS-b�Yb�F�ar��ъF--J�֫3pܰ��ݢ��c�ۂ��%Bʕn��.\�#n7�4�vԘѵ���T2 ���fAW�IF�-�j�����DC��ˮi���x�O��ԏ�^��yzi�t>I��6ԝ�p,�~�������ѹ�NN�b�(mBJ?YK!Aזv
���z���,��/Q����+��;�7�M��С�+��U|���w׌("���R����)��?I\O�}�:>�VƄ~�N_�;�ڰo�<B�[��6�q�GP[�Θ3|�()�nz�[�;x���i�VV�B-X1�x!��5]�e��{ލK���7+=�3�X�wo+�?#�c#U�b�}�^~��ƍ׮�����{� TF\(g��U�+�������罙���5d]uM�w�'d��5C�5��+��Hee<>4�p�5�u��J����l��>�J2�*T=G|֊?`=]V=c�K���P�:�ݹ�]��ט�]9�}�A�]����??2�
�b�~F���z+�baSz[�ڜ�+k�]R��㟯?X�x=��=���K�x*������o9o�*�P�;ElΛ����vk���j���+�<��o�xK�&o�L�>T/T�5cP��P�[.w��.32�zcT�h�J�X���v�#,�t�o���9�����vp��������&w��P��UA��>��o�ĥ���y�2��5�{µ�����K/,d�� h�>�*�c.�u�MCՒ�:�X�b���&Z��7�ixj���W�KW��g��F��u�2�&���5x6�c�7J�tAqd�}Ѽ?\�a(V4�^^\��.ݮ��1W�������Mn�9G�/�J����zد�T�(����=�0WҬ|�z�F��+<Vo�H��3��5>�n��+UBx"*_Ac@W%�_K1�وJEz!ۃ����v*��Q��5�+6˴:��}�+��dY�x�w�
������M���/hr�~��ۤ�{�4�g��ו��:�#��K�W�q�S�TU��6�����ɖ�݋�/`��}^>�I���:u�={��<�+�RX�d=�D>���EZ

�]��R#�*���#!+hfx@�
��~b�|t�Ɍ�:�~��ذTy����vRv�x<�]�����ܱu���/�S3���c�c��f5:k:�P�T㯍u�WO�س|�N"���N���� �<�����>?�­p������Q��Vq��U�\���kއ~W�)�W�Ϡ�e��4﮹����j��o�E��Q\�P����(�+�K<U|���ӲP��K�
�s�C��K��}��6�;X�(Uz�+M���e}�4���G�ҧ/�y�8���#���Wz���AA�z*�9w_q�e�}Z2�,��(���j�4����t�;5&����;��PWm_��:��,�����k�����4�<��&K�tj����S�+�R �Q��9���{6o���^�C6ӱ�ǝ�|ɂ��ȕb�}Z�TG_�v��WC�u=# (O���Z��^zꜼV:��Bʆ
jǀU�gֱ�d���;����׾#@R�u���2��2�]TVڷH|�=��\�	-Pb��F��w
�����<�����ЪՌل�7i��t�ѡ�|U	�&b1�36�(v�CjW/�D�d4��縋W�M���-޹gi�!ǋ���ȹ��������I9u��.#0@~���0]��>�lS�2��їeݏDА!���{zm�a���{��_h�B�0ؗJ�(
,�����t�T�6��[������H�~�A����yy���8��\�N������񋠯r�W��ʸ���e}��=�Pvǁe�G��©h�#�'ߋ�J?#��L��7�*4i�F�RV�ϕ[�}��R��}ޣ�*�j���i�'��#�on7�W����C���)��;�o��y
ݎ�U��rl�����wWPV���A�R�|@�����oU��]���F�$`���;���Y�y���j{�7�3o���us۝.d)�2*�r�����:��|�e���D#TP�)S�g��\,R7�$�?�_������Yrz��][\��"Ϩ�O������8';W;�Q'�]b��5� ��ܞÄ��-P��{��g�*�Q�䣺5z�l�zɳ�u�ۜm��Q	:P�ÚeT��R�-�SD²��jX߿����U��G!_��%`x�]/\�A����w���}t���n温E$��33����n���*V��q[#/��<~Fez��*�m�
�y���ܓ� ?J��b��cr@mZ��/��0=ʩ�|+
W�$u�@F�e^ E��_�.�Y�Q��X�E}u%B�����4P�4�S*¦���c�XtVv�ͿK�� Y��S٘�wO)�qs��`;X�U�x�}E�y�`�so�Q���Zm�Qr��C�o�>>��h��@r��q�4A���Ur�{^h�<,'D�?x�����֞#ӌ����:���D*�v��Q��&��k�������3�%
��:�_�#�Ddm/i+yT�+�ʳ'���zħ^�.�b����zˇ�3��e
��>;;��i����[�h���t]J�`�p��F�H��:!	yz�7׵���-9�Z�<��.�Y�"������e>�d=q=닇�%7�\�����{��)� �+�����GL:B�W�������P����vn���P?ʚ}`�W[��}~"W�-�� ��/��?b��a����{�������xQFh[=wǊ�9dx��Ș?��'O~|2�=珊�柕����=M
��_Ƒo�/E{��9��˛������V�!���y����~?O~?:R�TEUC-#O�.Ry���V��%a�i�<*[?�|ev/`^�/������~��Py�w>����*���`�}[.S���V-�U;��g\�'U5Nq����W���F��u�2�"X��T���׺��=���;mc4zg��R��+O0���,�
'���T�_�H��c��ok����ZQ`'��PSV%�G��WҕSWLлJ�>7�G�Y� ��>�X�}�W%�_K�>-�o�4Db��u6[��xN� dfXT<����T�Ls0� 3e��Q0[2��}�2�q�������{��-J�A����O��$׺�x�x5�Q���߻�[��|�}�o��2�W �/�-񣰙g�x$6�.�2-[WT�8|�#|o�y�$�]_��'���c?eܗ��i
��!�����J���N�.�i�1�ݮ�8 U��c�@(+��d����U�n�j\��)�O`��!��G�:���f�߸�X7ǝ��C%���߳��D먊�h���y�G�oX��g�ő�� ok;���w�h=Cpy�9��_�|��R��8+�j�̮�t���ܛL���[�מ�Q��z��l׆U��:�x�"���?;%W%��@���y*�ܤf�m��
�B�PVa�յ�e��y�q��+	��5o_E� ��֝�)Pb����v����=�]�h�t�r�}=�������/(3r��;�����}A`%��`�+����f�k��=vpY}�箭\ Ը�R|r���I�n����B�R�uj�M?x��9.,�D5g��H��Fp��A���q�]ȧ8�n�(�p͙�:r�%^^��Qh�Nl_������l�������z3��K�-ӣV���1w.��/������q��M~�9�J��j��ӱ�ǥ�|ɂ��%X�n��@�uJuV��-�[��9C_(/�V����玵�UT��+B�������.�ǺL�m�g��F�� "ĳ�4�(�J���빖�q�2�+��"��x�����W����F�HF`��튣C�T��m]I|:�1N��P/8��mٵb���/�`�iVP��%���_�U}��2Ѱr���~�Dl`��Q3�͇�(?����2q�ǝ�m!�e���� NN]&q������]Y��{��h��a��Ɇ���%*y{�/�P�ɅVo��a��������|>���������@���~����/-��z� ~�Y{�Me�a��	z����_p��0W�}o��f�&#���͜*���QϘƳV�t�P��Wk�>�p���
�MtWЂ#��Zn4Zݜ�S�:o8�I�)��S��[͡"�*�,J���M���"���I������Mn��T�^��Ы�@s����r�`�\V)���R��V<�h/l�pɧ�'�E~�/�J�}+�ӏ�2/`�s��&m8�N�^�>RvS7=�<2��Q�T��Uz�H]�-�^������_T»�/srx�?6�ר{�0������&X�G�~��g�ۆ٩����|�XT}a�Gs�(�r�+��̒�z�1�L��b���]O{Ƴj��_X�];X	���J�%�<�u�f�O�y�K��n�\"�c��Q���EO��D@~ꭺ�N����������«7��'�~�����	���V���>���W�"+�r���x�-���^�Hҋ>��M�e�K�a���?Ykb#�h�ͼ�?\�#�-��Dߟ��/0�s�LPx�@�r^|����T�}{Ka{^@_��{(�}{n9��opv�h�Lg8@\�:�NU��Q�[��lol�h�^U�vlY]���k���	�ھg�F'}�Wb�q(�C������̶��ε$��~����*:O��į�)3N�C���%z��<��9q�4F^<T7�GOMh��:OAM_��f*&�)#-�gƵV���5Z�j��Iぇ��Ξ��|�V���e`vb'��坚���s�t_y�Z�9k�>�^.�S��[g�J�wd$�?]z�WO�g㐱X6C7%���������ޤ=~��nZ��=b�]7�z>�*V���Xvz����D���~���/8�����W�a��,��^2��$ �߰+���~^�����x���a^n�m,��F�����w<�Ѧ��2�8,z�=_������Z�bu��{�|C�.N��G|���Q��
������UP��=C(uJ�����׻�r�R�\�hOz0B�uҹ��{�B�`q�2è�C����ptfb����6�q>��vWy����x*��b�����`w"\��^����,�nGZ�gg�D{R�CՕ�Tdn*w��X���W��{]��Gr0i���2b���o�n�Ǫ�ވ����{R�L�v;�ae�aպA	f�a���7�Ç��m�O��dγ�ݲ��;*�{����G���;�	D@��uDE<2{^r�kǂ�P���]TJk�K�Mښ����+����Jf.ޘ�jկ��h��N-}���|)!�k����9��Ѯ��1wQ���F�P��4x�Zt\�P+x���ܱI}�#�l��"��v{r�\yJ�]��KV��;V8;���v�lU*ZN�����0*j�s��w�Bػ/�KkZr	��Yy6Ų9��xD}�3�c4�$%"���N�Ӛ��Ғ���V]�z���4��GmܬCQڕ,ּ����H�<Z�����[y��â�szMz{ޕp��C.�:pn�cTP��ցƨ�%\L��W�F��p�T*X_Gh�M�v��E�{���
㡌+a{�ߓ�M���t���Yި�ݦ�B�v���Y�|�L�Yj_G]I;�D���ԨK� 
=��E��
X�֨e���}����X�����Հ�Ǣ�=N�[�&M��i��}�u�.�}3n@�	�J�=�D4
`����F��Ag��l�/�ח�i~CÞ
�CD-Y��e�O���rS��w\���8t=v��ڡoa����:Å�#�a�]J��Nb�4�G;@SI����rK�c0p<���Co��֘�uf�&*��;�5g6�#�ʅF��0LGk����T78���Z��l��]G й����Η�ȥ ��;�KB�ڱ}�,���΀�Մ�ݰQ�9�p�\��WZ:�=]׊P}�K�{�j���n���t�����V�D�F<�,·-M���ؓu�vc	����
wt·)*����`rK�!l�^�?�2Cw�� k��g���Z��i*��	Х+�䜛�Gim%������i�qhΦ|Ȥ��o4�����lں	�uGZM�`w��U���{��}�=��1eQ-�maQJ��J�ZYZ)�pT���LfW*�zp�X��Z�m®��֎��ш�����-Qq.�5�a�1mƹ[r�)�A��h-V���f9��+
�m*����Q��U]�+�qV+�[AJ�EK]m2�X�%����)s4�tj����mK(6�s)jV��nP��lCeV�LD��V��\\DT�����8�X;�.7w%�2�ŘԱ���Lrڊ*cL��,VZ�AEU������)imb�Kh�[[lCJ]J"�[���m��*T��lTQLۛj3v���L�53��kR�m���+T�"�"*,V.ndCZ�XR�g�wޘ��1��r��G����,g���ճ.�ʍ�`�*S�:e\):Xn��O߾���v���Ϩ����g�n�}��XņB5���\��K=�*=�K�n3�@���՝�>&Ö&
ƞ�,ӠU�*�X^Ӻ��m�
{���jd�}?��\���(	PW|��G��Wҧ;��s�.P�]t����@�n��c:�V*^���R_��_K���ǩ�{��F�ނ(��2O�D=����e���o��b�)�4�|�N��"�Z�+�}R�'������Vc?eܗ�t�/ib��w:�#�rN4�m�Va�-��zеC�{��.��T��3RC3G�L̢*}�`������^�C��G�/h����׼�xT�����?p�2���a��%���e�"�Vf��<�/�I�٧��%���_QyH�lz�=F�����CWo��?g�ݎK{���a����PnV�f��T���:[{�-Kw�,m��`f�+��l߬VN�BbNO�g�n��ڇnwY�9h�����d\��s�l�bk��d��Y���u�� >�{ן����=���������z�,:Y��T]�XdN�Bw�/{P�M�:�:ƫ
���P���]�Ճo�?i�Q���'���߈�;}���;�*1a����r��Ȍ���Wp�hq�Q?3�}�ϗ��}�%����Xc�g]0#�����p觳Wso��_�@o�'����]���ྐྵyb�2[��^};�0�yL-��K�����]FW�m�RXFǥ܄?�g����_����e�H��W[/��Tb*�m��B���n���,up�����^S���A��s�y��z���{kI����Uʆ߮�尮�{�d�����ۓ���^�wu�����lU���(��٩,Q�V�,��g�K}Ag���A����$Ka���z�`P>^��e��-�\��]�� ���:��x��"��?E�أ�Z��aK̠mK��:�Uڱ�*��QKvmc����ob4T\\t��'[��`�,lD����J�����f?������3,]1G��i\���>�M�y�����z·8?4���y6O���g���J�0W|+�X�<�g�D7�_^�y��n.��a^��������ك�e���Vש+��~�e߷�Ak�+Q�z�maAgo�R.����fܮ���?Cԫ>W��ے��y�mY����!�r��m�6i���U�J_��J$�<���&n��%���P�_V����P�e��l22g��f�����z{7�Q���fT=�� �(m1wv���	]P�X��	��h�&wk���+>��z�*#m��t.��E@�
wvErRoR	���A|���3�R�x���)e�/��a���i�݉h�=ݜ�����P��o��?u*�*R�/i৒�D;�g����GR��������KR�"��wn�yg����@;�e����uoM�
pF�;[���1i��g�������.t����I/Y��w��7\J��yA;|�~��_|*�v�7P��b/��܄Q@��[uB�舌�����ZC6�V���I���g��fQ�`�V����E���}g����U�1��e���aK���o���O)eXtZ����:�,:G��9un�Ǒ��yI�Ϯf�F��}\xl��<�	��9t�����⿞[���y��۾髽�^�0�?y�v�3�!��p+��S�����~yC�Y��w�F��� ��,mb��7L��c��r����uՕ戔��'����^�H���b}�F]�a�Y7��O�[�`ϴ�+�<C��?:�	�3|��F�f*�k#e�eK����({�%�Y��g��B�*��uL��^�rg��k?
�C��<�΂7t#��N~O�I+}��!��㮼F����t=�"���J�QذQ��"<G|��%뉎W]a�����{�~x��@
�YV��k< �U�geԺS��V�5���F1[�W*�K�kt,���[��N�|V���7���ĞwD�3Y��4�� �k�B���v�z����z��i�粣�e�3�S�;��iWj[��[�c����v;Qu��Ug��d<����W����*���\���eu��/D+�z�^
�'�����'�z�c��a�#��/�1���1G'�~�d���8�s��vrS��M-?yw)�>�2�ևr�u�l�B���Йmv?z|34/�� 0�<~^nI
������'j�UP}pm�����X!�cO�N���[�!;�F�����+�b����}���ܜ��(	PS�؏edz'ϫҽ�⿍^���quu�cv,`��*Y\�*���C+��z�\M}�7��b�z��O�Q�0�X��}{R��uKH�ƅA=�?+�C�ؐ>�DV��T(�ۨ���0�if{�S}W.�ְ&-j����̳t��-`)�՜�}5_�;�F[VXU7���,ev��=���j앏a�k��FE�<|¯ۮ�����3OM���y�8�r.�؟8��z�h�Ի��>��q���Ԡ���U-f��� U
���U�Ė!�7^�Z���9\�P��b��.9^��A�YpQ]�KG����6762���Lo���WP��B�ꂁ�r�_5�>�g+X�����dh����"o��W�����Q4��Fr��a�g?,߸іe%b]lӏ��0
����_���>�f��[���bHT�NnX��g�9(���tm!^����<��� Jb��άv�ʄ�*��p2sn3��į}��_Tv6�*��|(�*x<��n'�]�,~�������3���_�Cn���K�p_���vճ�XT��35$�a��eX��wق�뿥ܗ��Ճ:�uN�ל��]z�>��U�f�*!�э.�m�c�K�d���g͑*�9�-/$y�a�7��� �`[����|�_�1��ǷeGʺ;��d}��E�4��(9�q�n�w��{m+����G�?*�$����X�o:I5ߠ��L�е)�[Tt�O�>|4����n����+�w(fit�x�USw(z��B����~��UYB���W��~̯^N���칖��Q�-HӤ���(g3߰��ȼ�X��,�a,b��~��*
�7���v&��o�!����������D7�Ŝ;��?R(�+�o�W�Y_�����Mm?01�{?dY�7��l���O
�R�3�rc��d���~���K��d��+�
�,z<�e�+�x��g�m`{�1����������L���:J���ǫs����M�^W��Ў��^]к����~��^�<~f�AMB�Yr�M�_�gXu�B̻�y��x�b�ؔ�l��Z�҂C�o#�:�������g��!�*�uZo�=V���2/`#)��o��|+/WےB��/w�ɵYo��y��>�=H�N�N�&��/1� g*Nn�궿�T.����Jos{ӟ:����|����-K��&�צu�qe?�:�s��_W�(ߦ���ߴB�E�inW1�N���L�Wu�e��9��K��mrq��Z�w>��~5� ?xS���ul�����z��xs���EF�eA-��O��tz­�0]?\�A�a_�F̒��'�o,m��/Nok����H^�k3�[���w��9���|[�!/>����G,qa�t�f2ұ��{��\�F���a"�?T��^���z����>�G{s��0���^x[j����zeaU�RxD8�k:1�8qO�e��'����1HZ���-W1T>���%�R�>̃g<a�H��ʓ��\�x�'7S:�A;t�y�sL�D<^��ݘ��eg�F*��'B���)6uIŋb�=��p��xYxI�,��l���Ot�]<Ѿo�p/�]����'��K��
��d�Jf���q�ƀ�"�����T��'�<9@�S�~W�UJ�*l���mσyE(Gf�^'$�C7_�<���<�o�WF�&�o
0�tZ�0lW�&�g�_�j��N#�t�`�n���wd<���[��l{.z�B������
3��bg�����-W��V��[��N>��K��E�3����#8��T�I�joE{��čs��O�,�o�ȏ���~��΂wVW�s���'�X���R����Zé`��)0��i�ם�L�^	%O�!�mqv)��ƻ��[�Iy��k��.,NX�[a��z�����+�]�˓��|�̝u"�-:!h#�����`�]D��X�x�ñ:�!��s�U;�A+�a)���W�i-a`OA�ї+i�٫�E�yKz�b��؍��Gv%l�-=ž:\�,p�v�V�ӜW���_�^^�����8��:CK���AX��!:$���D
�5+�cN������ِ+�V�U�G����[����м�]o�"�S᪺̄���9���=��WN�KٶF䓈�\L�4��G
�kAw��nC�x�~}Ͻ4���x�lcv*3y:*Q�&��͚ɾ�d�����;�!RSj}�����*�X��b����^O=�ޓ82�H�Wl�V�e��M9صپ�(\��>QѯH/+���m�>ĥw��c��m�%Vv9�\��,{M�_��^X�ߘ2���G$��PE3T~/�z����X�.)/A���M��<��<]u3%��j1�#�h���/�6���0��m�rJ��gF\O�E^H6�Fα����yֆ���K�_)��0��fM"��}D��8_��,l̹��;�|���\������7�ٶ�>�E�dS����j�C3��W�7S�{>&�X��ld���̗)��Y��n��ui��u@m�o[��0*��9� ��)^[@�Z�ཛྷ����8�*���NQ�A�,P7�M��s�"�����iɝ��=!���W�}x����oK�c�����8�']ҵ�o4^g>�(ּ�<Ż7�+�đI~HNw=��� ^�,M��w:V��?M�76�v���VX��	,b_����-��g��۳%�9w�)��4�� ş����*Q̺D�"�S�+�8�M8s��ڨ]����dg�P]/��r@j���3M<�JJ󮂵��\.^�N3����iX����#,�b���g��y�,�ɤ���K�)�o�=��y@gr��(�/��H+*�3�8�b�&p��E�Q���OL� �O��t�[�*5�m���7�`�����qgu�Ao��	����"[�o��{��CɭU���\�f=?זa��N��`����p���s���Hr�=�74���@������t��^;;h�M78��|��R@�uI������m>!'�ף 6�����T��l�@�L�	q�+���i�s���k*_�x���s�sWjX�R�G��g���a�'.���۬S��k��<���bJ�K-�K�����TM'y��X���o��M���n��,�� �Y(_I�i�����'U���*�K�n"�7��J�s����9���b�N�żl�^�yu���:��Titl�"�]к�378�E�v�ѣ��^��E�1�y��qC�y�'��}d^곔���z��D*��_��ƶ����ŉ`��]i���+'Sw�1�\U�����N"ÅG��ԪlU�j���t@\�s�N��`9�9d��VHC���zx:;������N�H�|�}4xR�K��V�>�-)aHw�R�}b�2	n����-����6�s�-���w�z[/-�U|nT��&�֋5�C����Y�q����G-��� b�F�Q��.mF��֥J`�es%�T�cj8+Z����1�p�5�&�`�Z�aR��Up�*�*:�mQ�UM�++V"���(ۮ*�#j2�f�n�.��QJ��V֛������6�r�Fm���-����U�LB�h9h�Q��&�F��PEMk
�m���Sۙm�h�5*U���e�LlQ�ܥ˙Y����Z�e�8�B���b�Jj.ڍ�Z
*1J�Tk1�j�6��(�0V#�8kG-h�V�
�ZTr�DMj���A�ȸ��E�Wn���V�2�PDc�֛�b������W/�t�;�/��K\a���9�;|�z�V�9wA,ز{lf��I�`��o7^D�c?�=��O�@\��MY6<2�7�W�x�;���z�n�O{�����J�7�޽��|�Wo�f����~��.k[��d2`�hц崭U�9��G�
A�!�k�����p_Z�v����؅�������P�p6���=wY�묛蟪�
�$��~b��e����Y!{�C>a�Xe.�X.���ҝ����'���e�3E^�=�RR�����`�+ҬseuR����ō^�i3�P�9��^�=� ΪS�;֍��Z5��^#ϱ�����S+{���݌/8B���n��3.��9��#5���y��-��Sz�琸C9��*�)\����}�b���PM�iӴN�[���o����{��hג=�t���\&�[]�N��z�wDX
M'6��9��n�n���ﾫi{���<w�W��:r{���jIt����1{�T���x�tyB�m�t�_����v�{��O<Or����`Ls�=�O^yV�Ҁ���P� �`��j(}��-��?q��"�Au�ǲțw��e�����m��Ἄ�rv��}D �z���\	�?tR���q,��a{Z�m��u+ۍf����	�7ЋV#�2����[�O�]��5�Z��+�I,�����*?�g����[�屹х���Ƅ����>1��ԥ��:rL���x���F��-:(P��u ���=޷��^�B3&�TUg;��Y��� ���YMCb�9|~�ą����=��J>��享��ld�:��N�nL�8h�M ����Z�6T4�4��	X�ݭ�;�W�����G�g5u�#Wc�DS]N��);	ބ���C�d�gY�&u�P�:
B�UI���j���)�����8^����2�.�>�ή�w���@5�r�pw۸�f=ۛ��e�̙ѕ��dm�/
�\��i��W���?d�-����x��i%67�>-����� -tZ�0lW�&�v�Ng/�s^����ely[��/�k��xp���W��2�{�gmR�O��}�m6;��Ǘ��}�	Ҧ�rR:Ki*ІE�;B²c��N�f*��6�W��A�(h�9��_������ۙ_�W��7P/���o_�͖3r�%�9F�������V�������X�D��~�T��f�JmsІj��Kܚî�--�h�qen��CX.t(<X8Z�F�'�v�	^����W�e�}�<kO���O�@v��t�v|���{���{�[�Y~�{�D��ǚ��%�!�@���X��y�'/{zj�=�#����G$ʕp�]Q��.���B��5����Yy8Ԛ��x"��>���է�������4lr�LB4I0+���uW��J�yќ�j�jn�:�:�w,��;���ﮬ�QN���K)���E��̶V�{~/���{��<H�h�(�]p]D�½��f=��+z���m��r����)��Wu�q�㭭��L�ʻ�J������@3|F\�TS�g��V�r�A��va�{�u��\����,�F:�My�H�O�u�}`��������I8Yy�Ej�5�uՄD���#�:��ګ܅���4K���־0߯����Y8�#��o򪾡�w���*�^y5X��=F{��~�܇�fƴ���Iu�;k`�[o�_�;#H�-����sr�+�NN�s=�����,{O�h���Ｊ�	��z��nd��;�{���'3TXWCG��������$n�Ord�QO����\�_0�J溺��K���h������cϤ��]�4^I(Ϛ�V�n��]����7wQ��kZ/�v>�'f��2��G=n�u�=������5̿J�o��K��~J:�����A��u������U�3]>��&��s��-J�W���S�q�D	��R�ߘ5W�9��)ʘ�Yq����E��ԱbcB��a��߮�7�T�g��JK��]�:���ieQ�q��c�'b�MM�i�rp�����9��Da���M��/�,.�)��UT)�y���J�JyWW)�����A�o��^�mH�yiG4���y�7��K�����S���Iyka�n�/[rz�S��a�c�t���痻b~x.Q��{��K�z0|�Y�����ֺF�z眅��NOxdC��J���%_h�{w��.�b�
�6���r��\ױ�����+��t����r�]ʷ���5���!�:0��jo{�'�ך�M]j�cO&FnF�f����ё���9�����+�A�M	���m��o�9LW]�K��ֈ�\���
����zu;\q���B_��1	v��uZ0�V(+��t@���.T�����pr���Ƥۀ��G\jL9I���|J7�V�n����#s�BV��#����������s�W�����-�ȴyK�-�e���y�;������
n���C��z+/��<VM���/_H��o��;3�8�ac�ؠ�E�A�T4,������4��S��HN��D+׼Լ�X���\�!@��9\��rb��v�-zD2)��Q>�f~���^3{�N�<���Ԗ�t=�Zg8�5G�lz{Y��Mӎ3�x���@��Y)벽ܧ���K+�/*+��^�&f�3��$FU�,e>��s�^��ڶ�kL��E��:NH���*�{�3g)\C���O>[mⷫ]41��b��;O�|�C/�w8�~��X,g�1k�v������7lMz�{O$�1�����D���s؊�<6m��dD��T5۩���Na���ְ݉��Y�9�w9��U7��~���e���~�ww�u	��*��āR��w{�
��sM������	��tX����N�T�W��
f��W<�A]�q��v���Fk;m{�ڏ�si�tŉ��:�h�L��/����������ٖ'��Q���������������e���*.�q�R��<�kǷ��E��Q�R��]�U���s#��J0���Fxv>�a��o�:�Z1�W�kd"���H�aKe����!�:�<w�}�����H���z�����!#D�W@����m�Vӑ�!1u8؝z��Yܳ$y�����c�M�=�bxSW</��T���>���WG(G�]pg0yF��x:T�+����&��$j����R�4�}0XsZ��d�Pd�N�:��{�Jt��Tb}?k5�{r�6�o�U,�J�Yp�y-�ͺ�ɗfJy��tܹ��A��D��Q�݋K�a�+7���A��=h�!��~N�	U�o*t�JI�iwp��~?P}�xܬ݌�
�XGeh����KҖ�����m.W{��1�����5�.,��<։u���U�t���p�����m��'JR�l�UV�,����d�j?UIP�k�Me�ly�w�-�Օq�QK�D
rؼ���I�u���\`ڡI�&'=��l�{��(���������j�0�}�G�e�3v���٥�#=`�u��9e�o�Jz�c��ͥ"^W;{M�f"|�I�:���;p�U���ۂ򀓈}����տ:>A�uyP�缈�Ati�u>���?h�\�$�5P��m�C��s�ɷ�͵uE�3wY�Q?wa��ί���H��{����k[���}.B����B,9��pͺ/�ꎹ�Çޙ�/�2<�3�8L���|ԝU��^�#�0���^Ï�ӳ���e-~n-~�	�����F9Lg�z���Ϋ�G
�S4�w��T��x[#���v���T���.�+��OL/�}�c�Zd�at����]Dg���ѭ.]#�~^P[����1�@���!�̿a�3�D�����DM��H%��`�G#�}�{>�`��A�G{<hT�N�:�ϴ1�P������qf<��~r�z�q��U��;�E6�y�ګ܆�����v��V�����.���&�5��)w�M�mZ��c^������B���&��R][G����@h�y��q��*6:�ʶ��~�x�!���u��*���wF��"z�β��K�6���c���>��;{ʎ(}���P=��M=�W�S��iqngVgd�[����'D�:d/N'w��^�����־���q��7�Y������v�9��	F:��ͦ�4Nݨ���x����;�Ny�R�;�1�d�d �ˌ��=����o�Ȣh2���t-��=����7��z�\�v�H��wG	���v\���8>Rt�M��jmrB�j*��2�7OUF��N4z^,��I���;�V���� <��B2�d�פ���d��� k��k�vI�Z�T�6��^���-E�ꇉt�T�v�y�F�7F3��`�!3�^M�����r3˞��ܸz�5�p_L�^�f=S��N���dy�T�(�S�T^�ObS53�-�]�.Ş��ϐ<�{���6��-e�����K^��`i|���.�5���x��ђ�y:�f3��p�b�T�����wu%���w�5���bf�]}���zv���	�lor��ul�:������D#�1������y#�78�+�Nvs�f30f�OT5��#u�-��dI��ϗ��U�"뫡]�y	��ѥ���f�J�C��ו�N��j�dd�y�\9�$�~��	+�`���kK_$��)�(C�j���DC��5$�c��5��<]�W��ٰ�7;D��W����8���T`�ˋ����A�W�.��V_t�C8�,���nk�U����ze^,JzR��iwQ��3e�Ǚ׭�e질58o��W����'v����U�Lh~H�Lk��<}�S��*ouA�9HɌ\�Oe�op��Zx��}�$�d�Z%�]n��I��ޢE�6Ⲱ-��q�i��H��`Ξ��)���z�TX��*�ަ+��ln�a�ܸj�˝�X%K.@�Ɯ8�K}�������Kٸ�J�V5(�:˃YNڠ�1�p�����9K����r�u��*8�� �)�U#1����,��:R��QQ����Ebe�*�"ZQ-��V,jQ�ۉ�U6��7l��Z�-B���VE��EL�m�-��i���P�\j��6�DUa�Q��Z�fT�TLjf�������%�2�-0�-�-�ī.%f;J;j+pQA�+UT[m�3-B� ��ؘffQ0��m�ʸ�R�H���cr�e��eX���6�neX���.]�f6ц�jS�\h��&�S�QWzɓ���WS�̘�[m�77J�(��Gs28؍�\j�4�17.��a��fS�壯XJ��Ꚙ=%U�Z��q���*�PE�6�(^�
�ZV�e�6�ݱ�#Z��^�]�"�[���f������TUF�fYD|���}�eǩ	�y�]�c)��Ҋ�ޗ��tbom�z�����c�WE��C�������=#����3�]����r��8��i�c�F�؎�oH�{݀};���\*rO���㦫�����<ߣ~r�ר!�Xcϴx��j~�N��5�͊S�r3{Rpx:�>�`�u�ؼF�U#;���?+��]vϷǞ�b�%��Z�՞R����:d�f�{���y��#T�Lx(��pޯ`MR�^�w����Lk/W���8���Y�~w��y�k��k�Fv��C�3Y���Ӣ��7r��dƺw(}}C$xӖ���U�%N�]N끞�»�4l��e?jVFL�6I�ǂ�|x�h��9�Z#��:@�RDޡ��*�^���R�d��;�zb�}^��Oͧ�I]7����^9�d����A3�C1:�6�=�n���<\�'��u�W�'�U��UK�ڪ��$p�=��g�#g>�2Y�~��~�q�8e{�N�ʛb��ԏ*�>&$<�~���nN�K��v}3�*W����?p�E���e�h\���&�d��tY���)y:�5+T��k����=1�}X8�g�*����^�}��v�3h�!�xݳ��QѮ�="�U�ep.q��]��o<�a����U�Ƨ��g��`]�=����/������n1���5����HR��=�P��y��r#�lR^(,�x�/݌�M~���k�o�!�����}�U3B���ě��߶d)�;|u��ܒ��R���:��M�>�ww�d�*�;�P�Ԟ���!9��5ڎ<E��ںK��&�I�M�o9�(މ��Ȝ��cz�>�(�&�t莐���ݸ��爦�M��䣦�=�� Z짽���M���brŶV�(���&�~���X���ϩ_�1��^	ċ��ph�]�����nN�5.���F�@�G�C�I��zT��x�i�S�CG�H���MG�����y$h�殽���m����)9�����v�g&���|}W��?k�+�9j{oJ��\h��xW�b���{�FQ���l�7v��\q�g��J�貈~cv���D�wE�Y^F���@O�N~xk�A�m�Ϳ/]@6}ޑ��d�ޏA�98���5��\~Iv"�~��N4��)xz����,���:�ﵷ%����OO3wlp�I�i�mۼ騜C��^M�Ze��QZ���w5u
O:<����.��&]3S�0uC��F��q�e������.�0dF�Px�\�c_Qo����P;�������1zj���w��ihW��U��˲�ٓܙ�9�͖�t�JCɪa}�޸�%]̾����7���OO���5��<t.m覭�7���<t�7dP�������~�KYx#�Duk�k$�?z ���r���rߡ��Z�~�}�o�k`���I(��&�@�!a�Cʽ�T�����s/�m��'/ݭ�����44�, ��8��������=#L��0w�kj@Z�� �V���/۷��Lf{��2j�]kEE�	c�DS���d�
D:�j*g�ѻ��/�U��3�B�XR5v��w
媱z�{w��o��� Nk���p���4>��s��~	�u��FH������Vk�DJ|�Wh����&�d�SIT)K��<�,Y�#:;��{
Y���>Wx��=? �x�^��7Y�
�������'[d��������:v�6��S^Qr�S�5"B�Y�i�S��=��_��O��1�.[CG<~��x���ݺ�>�{���e@[SQy���^��/��Y�G�(.L�9��zl~|�h�i���r��G�j����۷/c���u�7�h�4R�X�.�����5o�i�k�9)�Q�3�	V�-�h�N�O݋���4�G�}�m߽LS���y�,`H��3�>;n0�o��\c��u�y�Ƅ��X���J�{�e��L�NK����'�=�o�ɴǂ��}j�_y�P�K����2f�����j��{e�;�)�ݏ�3Ւ a]<ʙ��u#�tp�>��xad��ǋxu]r-��,ϯ)�w�W%"�-Le�
b	�$Nv�Y��e\��Zz�q��>������{�������Mb�t�S�, �p��K}U�{�.)ժ��_�>���m̖��&�5 ?4�[��wAG[����]���p7���Ɂ_@�����6�}�5�6�[s[?@����c���d���J�u:;u��s�T7�#���}��1�q�\�~Y]2j���w4��"}��q��_>���R<� �bŭ�C}���K܉JY=ZEw�0Ǟ^�)òj�ɫ��Z�n���Ld,o�b��"��]��W33�P��L�q)b��7�m�{q�uMz�F�F��u��[$�M����Goԍ��
CU�d�5��	�.�ɲ�4`wz䅬�Z�Noj��Ux�(z��N�ޙ�h/�?e:���2�U&N)�%�����nN�+�&>c����-�z�����ƛ2e�6g�(j>��W���I�p����Z�ޡ]�=�����l���"���m�ӻ��
�����(h�I˲"W�4���.S�������{�5$A�,�)OQ�]M<��ܙ�B�w��7��o���[�T��u���Il}�ޑw`Te�u�~���}�����l��N��ޒ ��������e_��^�Yy��nE�LH�de��D����bS���Nu`�U3I�u���Ҷr�Q�����8��|��ǝ_�r���q�	[�7���/�W�;�-HZ�d(J�k"�w4�!�A�M5���{�A�(s�MƊ�'��L�����~��'6\��d�>LL83�>B.��gg��������ktl�?ևZ��*�@��6�b�p��R�Yu�}JO�z�B�Bv�Nzg��0���w�t�JJ�:0�vE��}_}�c��9~V0O��c����u����c&���t�������p��7c�d}�ۿ��47;����w�s�T񇁰+ޏ~>9;�#\�5�/��ܹ��~�G�yk�.�U����օ��<���_V���\�f�^a�ϟ>�RP�h���`�}��	}x��o���Q�~X��v'�R�����<{��R�&�4�u��{�^;��a�{M\������>n*���7��6�DG�;Q�����O4.G��_{g����z#������	��bwS��g5��o��N)�m��<��GyR���/��>�'נ�mKI��o3�-6�]%:v(����]]��w�M������)�F�J���iT��^}@^���U!�ۙE�qhǵ�k�.�H;��9��:=����>��n��XI�DZ��i��AX�Ts�������\�78i8X�����5+�G)���P?vae�F�%
�W�Ϲ�S��鮧|��ɹNs�5:�7�
9�<1�sL���B��X��/w���t��D�UϠ��<��.M�0� ��A�{v������c��>��Sw+QoV���`�g:>����ᇱ�����1��ݴ9��"���ܞ�N�C��Q����ϕ^+~�U�f�/�1���rK���&�/&_�:���X�g���c�~�;j��f/w��?
�vk�����:�V�k��r����ߚ+�n�{u�)׬"U���d�:��'����F,�����wL��֎o<�i�ݑ�~1�Z��)��w��!��ʆѭ(���X(T�t�Uŏ['.܉��$�Ҭa���4o�?��^]��o+�bx�F���go4L*jf�t�!g���_#���@�Cêz'�뻉x�ރ۾I�z��5����(x?���jG��r{,�v����fE�4����$Ͷv����ϯU	��w�gl�a�콞�d0�rű�)k{-����R�o>3��^�\����U�Ӫ�t�)ܩ~|�Q7�}(M^6Ķ��Ɋ�U^[R�}=}蚤3����-<��Ig���3������Wy��I�!�U.:�����p�~͘��g��o7�I>{�79�_8ں��x5��Ud�����~�.��?QO��[wS�����j:[ld �z$�%��wb���[�]���1��ř�h�i�s�)���E��Tj�ԎF}�{O��.��;V��R[d�������v�o}�h<��J_CE�q�N�v�Ng:{3'J�V�6�՛g���9n{b�e���KW��{"������.Ʈ*)��ו��RV%�q�olE�4��k��̎�a0�4'9�����1w۔x]@1�t��V�^�2��YL�]}Wn�W{|���l����T���<(���	���F���&�1W:�ߕ:F��~���03�a��R���cr ]�<h�5�cy||�h�B�yݣ7�qF�˗��|^�JU��Go�R�w#��N�S�k��8�� n�K��!ݨ,m��6��W�w<<�*�� S�X�1���}rm6�b�|�>��06�'��l�#������Y�鶖��%�A��-	N���"Y�v:���S)�̥�1p�P�Aa*�����^̖�^���L;��M�?d����zTbK���v��
�ke��eL{y��]�EH^A{�j��8���	6��bSX��}���e�En)�I�>�K)J��C����jK������=^'u�Xv��v��Ʌ��Et�us\7Ҟ5��z���^ǁ�T>�Y�˭�ϒ'gP%(�5��y�yt6&�yr��}�d(��t�f�K�`r�$���ܝ�F{��H]����s�0�|��ǩ��{�U�U��5�x��Pf�����v�h�����!�O(��Լ��ևki�)�K+C��N;q�������G%�g.ܝ�a_�k8U���0B���6����{�C5v2�*��Z�w�S�6]�>K}�A $0��:��G�xo����R��a�U�N���P\֕��[���a��T[���Ev(q���%���$�[㗗�2�[J�M�ZcH�۵�+�+�Xw����Rm7[� Tpd1-0n���{��1���V�ku��3�9cJ�Y[��	�)��������������0�Ub��ݥ�F"0Qƪ�bTU5*e�c����R�*!l(�6�q��Er��*"ۮE�u�j̵�X�mij� �b5�[�6o�fڔk�1DUjS�Fӧw1M�X`ݸ[LۺY�V+�eVh�kJ��F��-j;]��w53iUG��v�R=R�U��QDX��G-ޛ�i��lnZ��v��DGRŉ�J�DfSz޶�ٖ۹��T��J�W�� ��6�:��L�+[k�em��b � ��t�2؈[A��fTm��kbb�iY�LA��r�0�"9�Q)�c:h���\�3R��(����+B���dEF+��ݕ��ˊ%V�ř�˷��γ1[
e%īY�J���ܝ4����*eK�7M3iE)aE�a��1i��Gw&*��Q�h.0S�3sR�X"�S�}�;󾵫�,H���2�h��ɪ�z�K11Z/���P�[�m�|u�'��>�`��Nrg����Ϸ�(��q�Wȫ1e��Þ�0�&R\���rw��Nt�c1�}�G�ek�f�v�6�>�F̈́`���?��0�þk����K-{k��pt����H�B�:��m��	y�R�տn.^�<J~�El�!���������+�_f�v���e/Df{�M\����%��)����-��B^���r�<�O�x�,��w�~��(���w��lxP~�6�n���OF�)kNy�)a��ڻ̾�\��KJ��1�ގ>��@Ѵ��{�зoŪ0#��fk�����̼���!��!}Ї�Ǯ2j!��<�]s��c!����޳�����4�4jd��cW�wJ0F߻���~:�_<,r�V�n%.�s{c)���p���J���Ψ�f�\�ox3w�H=��X\v���>����bX���@�e{��8�Aoya�N��u��C���U�~��X.�6���HjQ�,KG�/y�j��xK�ؓQ�*}��;��CU,�HA�}2=��,�&0�rG��'e���s�	��v��zN��2���ޒ
�f̀�J4=�bV#+Ӳ�+���6����t}Zǜ�f^��r���у�
�Z����^�jIՃPc����%��g��������:��ؤl�9y������U��ۏ�+�T���]�����y�N/������(�P�cB��S�`�Ku�6��ed-N���j3;�΍�x&��uߘ*�g{�gloPG|s���\>��̥bE�譎4��=l��m��*:1��i�	Ap������=���|�^͛�	�]ɔ�1�OS� �E� �pkO$*b���G9$����M;�\�"���imū�y���'���ۛ�C�ܑ&���
������K���ދ+�����'
��9��]����ԟ;~D[DZ#����2s�y<�1�N�so:�ڒ���Y�Dl��C�E��"4v�lo?oQ��E,a��0�Nw���-��᪃y~����(��������`�̝u !�.ܯ0��ͫ�7�Rs���2GGJ��~'|��@�;���ˉ�H�5D�;��(��vFLg�'��W���jd�x�N9�Y��*�5�[�xOn���n�r�`�d��Y���1tO�®'~e���0�=׾g���A��;u����ζ�#F�X������q�2�,tԫ���GE�'�h����;��L
۾��K^,�v�d,��S\��s����-�=��� Y��%�Jˮ�^�)��"�(���|��e�^p,���7�8k����.�<�yz6u��Id/;�Z�^��/8胶=�jC���`��8x��9��Nk�.<�MN�cݓ_��
^���B�N۰\���ȼ���X�w~�ٽ}Y��IG���̃�d6���2���ӓ���>�g����_:O>԰O9��G�i�)��zv3=�F���$w"ذ�KGh�))~��?zto��z�ɡ����I�ے��E�U��b�(6m��/� ���S�^�\1��}�F',alռ��eKMG'�)��z�������_�GS�4h֝?V�W{z�ԉ!�N�m����u��+�I��Sˬ�8���d��,{z$�+=C����U1ul��Üc��5�\:���"�a=���|m���Y�\�������F�=nD[~�X�#a�y!�"�<_���]������9I? ��|�^ߤ����X�@�GvP��^���HyЧ�dw��D�`Õ�}��oe�Op!�7�J�L_�c�t�Eq��|=�ع�J��=��=�ݸ���q�e�'iW�Z��u�/��;�Q�V}�^&���7�b�vDs�*����D�y8�6&!��Ƕ4|H;#�7�w�+�zԒu����U*��zY�B>]Z�P׉P5�]��o��$�<��ʟ�j���ۤ]Ք�<�|eRt���NL�)��'�RTC
�h���j���Ooed<k}4�ܰ���-�n��hyw^�]vT+�� �<ë�|i?����1�>�G���ه������^t�ֲَ����sf��Π���Ot5�M�r��nn��nkI�J����/�L��Z�:T�b
��hf�so��L���{�1ٹ���Z�d�N�f���8��s�7��+�������b�4���k��D���ApޭjÈdy����{�cމso�t�!�@�j�����aXn�ɥ"�޳��蛘2�����BA�J�W��՗%x�Kj{0_I��ɫ'"Eg���X�xS��3�
�ہs'�z)~�(���Úd�c�y�����Y��ּ�F�$w����$����`���wj����Ln*�t�R�F��~u�k!oP�=�Ƹt��&���ٞ�s˳�J�*��w���"�3b�qa���1�{�\��^b�Oe-�u���Věe=��f�����L2U�K8X�ם��v������g1y���;���z<7������Ӹ{ӥޯN{��B�ȋ8�?v�)V���m���ƴj~]�s<��_"�����G(�C��%/&8�����e�����]�j���F\G��O��r�Q�������\���K�l�3���c�(�oyۛ�Mޜ�V��@���q21�~xf(��϶�~��<��1�%���,��C#=73�H���\�R,�}3�f��&m�cy>�����>~��kp�[�Hy����G�I��?br��˾�e���J��!^��@���q"�5  4�ږ~^4�{}��ȇmH���d֦���w��6gHW`�r��:�7m�I�x��C�=�-ˍ~���f�%�Ҧ�76���T��]�[PN͚Zz��ܺ}Q�|�(�Y�C2���MP�k�X�/��}�rg����g����D��y��#��lw�,쓩��7j��tT�����B{���m��n�d8w7t��g�Z83.q�9ǉj7e�Z4_W���߆cѾ��X�L��O�rW>��>�~�DB�3��7����d\4��=z^��xve�����1mǅ��C�l-/[��^^~���o��Ϗ�3ܱ �������2U��Y��x��]t�o�T��qKm��َP����O1k;�d�ek�I�	�zk=������rk�����_$�gt�y��/������듒�s�d���ٹ�غkZ@fP��J�1�*�PnZ�&S�룖�Wf��5�w,�z�Yۗ�\��ް%�i��d�%m���i	w����&�=4k���P�2�v��E�/[���uS��^^bM�9>�Ͻ�<�RMv/��])V3�	���Frˌ��cϤⷎ�5[r\��}J��Q��ӛ"�zn�q�k�"��c��19`���b����(�� ��}�2&pƳYx'.L�FG��y�J6�U!�B
��ؖ/#�!:$�����b�rګ��^��Pb��t�M�����K9�,(�:N������%@�����zS�:x[N�{*�)U��-�Lӄ<#�\g��R��н���ߴS�_�K��_ٓv��A�@�_���X�*]�zVoTnk��w>�x��ek���lnj��dG�?t��5G�� w�(�`o�ʥ,��^˺S����m�ﶼ�z�7��%�#�E��K�]%�u/�t��\��G�n�/��[�J���t{��<{�/0���̻�A���VL�j��E��zu��(81灱^�z|NN9�3Zl(�Ih-������y�^��yhF��n�����̝4���l�q��*�t)���	�y�������S�=E���X���,/�xW^WN�oH��{~���?/d���-I5ک[G��wggJ�=䚡�!>��S@�4�ڏX�Z�2��(���V�bS���]O���Q����Z��WX:g%.y7�\��S�t#m�!�^�ɩa�K�����9&��o��A�:
����E�`7��x��vo.��8x����IQ���n�ʿ��l+���̢�s��RO�4�z�giO�%���z���@%p�މ�X�[0f�2��nM�w�[�Dn�gG�ۡ��LF���}{9NU�*ʧ�Bx]s���]�Zȯ�����7�n�G���j�.�TM8�!���v=�w9�ٛJ���86�>�&8�İ�c���%�kib���:�B8�ޜ�9����O5��?T���u�/�ɜ[�#t���c���+�R��N%�w(�ː,��,��^�9�s��Ưm�D7�Xv�h��9H2�+�w������X��_��H�r�>�f���C�ɇ:�#��.z��}��ϐF`������K��^z��h`t��tS���e[T�d�|��뮥�R���3����w�g]e�)v[�Ws�Xf/��i�"#�z�����ir�ڶ�WHqou��Z[�ܥ��k�2��+j����ѴW
�5k�f���v2{^�����8y��ݚ�{8F�hbLW�ofɍ���u~a֍�Z���G�ޔ��3�o^��lѳ�!�/��Ő�[�7�Ґ}aأ�M�/W�����v��;3�s�y�� ���O�{�g�7H�z��VX��(��㠋7��� �m���)ul����FX��"%{�'[��E�L3q��eY-R� ��靃�#O����嫽�$��`
D��jֽozC�q�$`���n\�vj�%�9�;�������藳�ih�)c����{f��7ݒ�d1]޽��x�y�w� �� �ty�6�&����ŬZ��
�ҫ�q�(��zE&�z�"�c8�������]�����oo,`�� ��p}t4,(%��2���2���w܎t[���5Ϡ˱VB�¢<$���?�y�荵Ǩ�EVB�#����6�ٲg�l$�qy�s�����ۼޒ���ѻEst�.Ɔ*˧����-8�.1J��>]��򥯗J}�VQ�\�B33>�Œ���F�5d|onݠuX�����$]�^�Lk���9��J���iؔ�"M ��,�H�veIq�ϲ��yI��}�p0�^.���5ݲb\��0}�����b�Pȵ)P�;J*��l7)���r�72+2�J�*��f`cV2�*��Spܹh��.�Җ{a�CPD��f"�."̶*��^��W.�Fc.m�5&��[����SJ��b(8%SRĭ�pƘ��2���,lb,r�D@w0�w3s\�*��-�\�u�����3s\Gi3+KL��-������̫X��s)�Ҷ��น*T+�]��-���u��0V�ڕ�F��QE�c0T\B��3w)�r�j��2�-\����J��ٙ\�05�-�5�����q��W�E�3���r�:ш��"�ձV��Rܶ*.]��CR�����,R���4�7�]�[TM�6�m(5��rՊ�(�\IӻeQY�Y���&�U�e�L�
F3,��S��KJ4n2�rcUS.3R�ؔ�ܻ��sj�+Y*�F��-V�ZR��[+7MkQW[��n([X�zi��i-�3��_��Z��|���O1g�y�o-p9���R�+B|�t6�,�;����F�M��2���FxT���k��; �{���Ȝ��8��9�S���=�WQr�Et.�n9�[��8�&��0`��4����_z�;�����#¯�p�����=M��7��.Б���24<��]�ǏS�9��=6G<�*'�Alf��; ѧ�-�zў|W.����o����^`E��J����ꠧ�Nޥ/zd��/.�z���!4q�F��/��Oͧb��ڵ4���5c]�ӈ�OM�˫b~�`7�^�{A��A�E��
���z�M6BCg��ZG��_�ϝ1N����wh%���FTǡ��彽獟�u>ʆY�����iή
�@�]^�'�ڱ���W��G��cO��uЏ;��×�Je4�ot���y��5ձ]��� T�ٝr�-:�ј�;�g�l����ȭ�A��������)Vv�����/<#Sh����Ll/�7�WX�u�ƫދ�gl�jx<�0����f',p,Z��t)�wn�ɑ_\��C-p�^N$\G�4�˘��v�m��^���6)޼��ĳ�!~'+���X\����<�V�����E������'u����b�����!q�U5W�p^���3�<�/��+0�������^U��6���_���ſu�U�.8=�kN��nw�����GF�<��ʤ9�v[��M��^N�q�#D�R�
Oa���<"����ɏNz��}�Ҏ�dA���<���s��z��Ct.�˄CZ��-u.���Ve֜p�F�����b�vR��W��lew^n �K�˦>�-vEK��2�j�+7��iiNt�)�M9���u�T�.H"�;ެ�߭ p%|��Gk��f�!�~.�<�.v������]��v�o����w���#��7�[@�X3�y2B�MXӝ��q{�^�e�WΗ�\G�����^�{��=�.{����:+B��3�H8��N�ҟZ�|����[��y}�MV�9,�!<ۘ�֭���F���퍝~�_#������hm��;���4W�,�hz�m���8cY����׬��v�/���U��^��E�Aw��/#��-z��s/�����ߦ���:����+��������F��j�E\��]�Hp��a�q��t��ծ"yຕG	�5P���C*^����ʲ����:�e0^��R�\t�vd��	�M�ob'�d2P������˝�I{��X	o�ߝ@�B���������Ьn�1(��l9��J4�ꔱN6��b�`|�7,����P|������y�SFe2A��C��kM�Q�n���:{��z���csP�����%�X1w�"�^�c&�J����^�z�8��s���j��2�/a^�q�&m2�M�Tz�p�"��涺v�ǵ��wyHK8�{�ɣ�˴F�7=v����WuZ４g�8�Ӣ���>�b�T�k{8CO���wv���AϯE�:���?���~�A�&���}��Ԏ�i��x](~�Y�S�����U�A��B��}�Y�κ-՞sV��8��n	����p�-�*.-��,���^B�`��688�ST��̅��kYh��:S={��������'�Q�O('j>��gZM��پ=�J�=~T��v=��0�֖�SA�;ש�T��v�;��g�#�z8zf_��N }|�bO�
8}Z�a�4p�
C8u�x�a5g�w��{��RC�s`��I�q?\F���	�tN)nǭ�g����u`�,p�8N���w�E�r�I(����gg!gnNl+Ε{�p�y4���8���(��a�ӎC�VV�@fĢ�:O��W���Q�$��o9ۧ�N*�����k{�ŏ��z��b}����e[��h��.�oN�Y�yǶ���G�3�6u��X���߇j��J��y���zX@����[H�@��O9��Q�q�kyG�Ի��q����ou���xT��g<�x������V�Ȕ��)V�C[:���)�%;��#��1p��xmw|�N��6	Nb���N���*?O{�Z��;
�S�6�F9ӕzz��}�k��gNrL�3w�z�D��5�V�k���p�-��ݞ���u����{�J�Nļ6�s�%2���O�L��%���B
�O"g��H�wb���M(���bpl/E�����L�u=��y9/A���S2p[�d�Lz6_�8o
�nM\�s��r{c}ky��~��9�)������;�����X���
g�4�v����F�ϛ���}���mт��{,+�@^5%��0ir��y_�������t6V�u,�e�r�6;�o~�$7����C�w^׺�v��#-�#�$�b�T;�[��1���8_��ZO�"w���!�N7�ˢ8�#���#5�Њ\��1#s��sލ������efNM�;U>���N�Vmukj ,��s��L�I��IU�~���7v�K+E�ɻ��W`�ϱ1��� 8���{Su#ح�8�׾�]��ﰤ�����抵f,�9��Q��Ú�8��Y.g�N6j������x��eK/2��jʊ'�T�7���|m���EM�rĠ��Vuh����F0(7�d���qC�ߌϯ����`ԧm��O��7ſOL ɭŋ�:��Z�^�gI�O���3�r��k����v��|�X��;E�N�q�Yk}$��g:a��O>�Ƥ��a��� ��{GPЕ4��1��W����do:۠ګ2N�^��gj]t��w�ԕ6�$�wRA]b��+�A�,Cm�±Y���O�kX�6����1s]E�c6ݾ�:ծ��Q�C1�=y�8�/���Oftjd�s9�x���V��Ia}�[֗| �,�zl�h��1�]���7W^����C�lV"1���{�"�ڻT���ZFZ�D"�Ms�Q՟@�o,�4��(�:��O6GoGv9�~�,.tZe�β£�����?Ge�ܳ��
�BX�-HCU,�(:����9u�fM�w���`C��!q��6�WG^���F�$-�Y�O����:��f2A^�î�1��"��F���?^�3�ْ{-��<7� J��!���ٲ�i�)�2އ��7Z�N9��;���z=��g���זL.v|��vuP87<GGu�גٹ+=H8���a;̛f�˘��}y�iױl�& ��{�+�T1:�_)�)�Os9ֽԥ����0�g��z�ҜM�gT�x���J��6���q�܇7���;㭗;	g9�����Ì�|ץ(i��?ѧ�הS������[��z4�E�zy�Nf�Mm?�1g�J�t�/E��|G�"4����~�&~��W��X�;V�_��p���W}<h'�eŹ�qՒ�5m������"��̒W}>w�����a�+$a��%�VwF��N��2s��@��a��^���#��*���gdI;SFE��`>d\��֝
C�{���i['����J�o[᷁7�n! ֥�A�<O�/}��;�P��ަs7��P�J��R�+��n��9���>��&��n�:~���Kg.D:�(`�SӢ��C�嬲�o�٪��Ʋ�Xe[ޓ�ˈ�j���L�L�{��O+y�>��ojg�Q�W��M5����n�D�,�}���"��<�����NG����@aǵ���%(@��jg�⻿rY�v)��Gwg/�D���x�ĮF�Df��oI���W�M�U4�;T������诂���{����u��t����7���V�-�~�/ű�Э�u_��zzG�ᚳ��K�%�qګ�%Z��}�Ƹ'�'AW/^���y5����M���l�g�>��ɲL��<�jπ�[�D�"��er��G�l�Wfh=�ȥ�*aw�{���`�ļ��r�ח�8��_��r���YA!��r&��X#��������x@~����P��X��mJ|�mJ���y8r�Kc�-�l�i�F������<k��2��z� ��MK����ה��%��U`H����*�F�rt��o7ަKc�ʡ[�)5Ir��wz��y~=CZ�.���T�n�z-�ʴ����7]�.��E�˾�$�G�n���T_Gy�XBi%�ﮍ�`t{*+�jx�'��˃{i��n��4�͙	)�QU�c�؎��<��)R��w[DN�)k�w�A�=�I-� )��{��A&�����,��Ft�X�:�r���։�F�eA(m�񀬅s�L�Ժf���*[������+�}ᆁ�X@M�cq�A=lw�$����:�y��.�8�R6��:Qn�},�-�QQ��2WYn!G�V�5���<Ϻ!REV�F���j��ui�q9�d�Sҝ֢o��gF�@���	�Y�G��]��4ۄn`�+�1ެ�	���#��z��G�����F�����,�3+wQ�����4y����(|��1��Ϩ��{t���qB�]�bRٺA�;]�$�J�hd:%���\�̭��]Czq�u'��k/.pÛK���2̶�]�[���]� (X�'i�Ԧ�&v�+)�I��֋&��~?f4ujN�so2���l�r��*��
s�2j�ʽ?k���m��C�\��n[Ļwq|�敤�Pݦ�+)P�b<scG|M�y�#�͈WC�+&f�t���]��/B��4��ݮ�^j}��؊6V@IYYI��6�Ύ��Ev�L�s�@c}xEq���õ���b� [�������n^d�R5��c��r���4�7t���Y,R�%���YW�F�Z[7* ��&��/��gj0�X���]4���5��&�`ڕwu�/���bW��+6.�֦ye<�<�I����0͸�P�c��ֽP����a�g(��Cb���=7���o\�趎 ޭ�;hڔ�3"T��MS�¯TY��m�����R��/��Z�uG�nKS�d#|�Wd�a�3m�>U�A�i��\	��-�3b�e�uBs���9�<r�>J����"�K<��K��1�	�Lk+Œ�r;ܩ.S쮗������ۃ8.F���e&�n^D��	n�͋������
Z�*��~��Q����m�-������"!X�)���Ģ���M�\\���2�-m��V���Z%e��۷m���Q�T��l\n%�j6�孥�)��m�T�p�n!��+(ʶ�������յ�l�K���6墌�]f*k�ZZRڥV���U֩Z��*L�W\E��ʭ�Ww(Zc�.V��F�Μsb���B�ʘ[-���5��ʮk�e��P̨�S��i��`���r.Ss2\�1�.���q]e�ʍ��R۸\J�s(aU\�2㹤�m+��E.�u�R��E�ƈ��%ۃ�յ���t����,���V��*�Q�H���I[.�[��)m�����|�7�=���z�κ�ʙ�_j��}�������wZ��	�B��U���dP,}]�9�sIǺ�6Eo��$�6x�ʏ��a�劯LI�V�g�m�N�H�������Pҵ��8���s�&N�u������T�p����ľ�h��
��s�{�wz8�
��/y���:/6;0ن��b�A᧽���ܾ���� GFB��\��8P�߶���j�b�;�ߊ�9⏱��s���F���=��x�h��/D6H���O��g7�feiwZ��E�{	�����'�m�:N9��uF�z��sq�S��ʵ��qV���.x7^�����X�f{�~�U�%�[�'g�vI��Ҟ$;M���P=��!����Z>N�yAj�C-iR����{kmOW
㥎g�	�7#Z�&gm���y�U:�uX��Y�6��ԃyI�Z���R���+�	Z��Dgjގa��6�k;u�˺�'�En��ns�����hyU�ҝ��Ь��+{>ի���ަi�~o���M��ֱ���
��HU��3��|�����*��%�.?dOa�I6�.����ߓ�W�����}�Xu�9g��<����E�E�cZ��x{�]Kp5��+ޛ;@�����{���4�9ce�!롷58cH��wZ�+.�6�Yw�Ҏ��]����6��H�����o��T��~��U�4ŅΈi��;�yhƪ�!����2��g��^�;���Z���\vo�xW����`���l8�;sLa�'���~�hl~7�n�˛i��ʏLJM(,�Ng���yhP	}��Ӻkm��S�5��3&r�.m,P%A��Lй7��kU������N��!!WN���W���ޝ���D�L�0{2N�<�2g�/��U2=[u����G:���Sf������V�����桷G�Z^�;g��8���6qd��5E��� ��ˣ4@4��DW�'k�v�%�'�;UU�p�7�z;:�m��P��md�kE�]�g>|�(T4�~�y6s�?8*�ٯ|��Ny�b��*w����I���i�=��ٽ���p_��?�m��xl����8����>��3|���o�<,
p�"3�>�Ki,�G{}��=y�fdE䒈�;��F��{�8=�w��w�iz'u���v;'`ɮ�F�t����7��%�[�p�4�!�6��\��=yZe��j���e'�z���4�b��j������٤�k���c�M��3�'��[7&ۖNZm��\��|5������P�jXߍ�f�6�l� ����5��
C�z��?e-��z�.PҠ[��Xǉ$�.#R�/fqU����F���T�����V����s�ߺps��x�����7e_	�x|�h^��,�:�ByޯxC���D�� �W!�U���s�kwH�%_�_o7Q����Oi�z��\�j��7��us��X�ʓc���z>����e�F��C�X�xy�k��]�����=G��q�7�?;�Bi�Z����'�o�F�פ��������~#y�|Фf�8b�Pw��?;(�/;�ҕ�P��^���kPՍa���ƪ��!ڗ�U��B�ʫ��2ھ'TY��`i«Q���;v�Ί�#VVjgu���X�V(6�q֧��%�_F��![�U�[�6(k�2�3����z8��_W
����Z�,�kp����T��W,���-�7�{w/T����s#b/����u����2'U{(L|s�f�#�L�m�t�؈�^�r���o\�Ս�rjPW��#�"��\Y�M�=�O����5�|����q4��'�Ҥ�q`���;�<t|�^�b��o����V}��ב�ԫ�I�VJ���E�D=[��ȰH^�Z��S�H�]�*D��W�q�ם��}!�^���xq���Szo˪��
�����W��D�(3w=ۋ� ϕr�m]?^]c�B��x��]zq��z&��悔3:NK{�Wڳ�ڹ[�(^T/����4�}�u2�ӆl�tp�H⳱�J�ʗ����4K�c�Wn_
�q��'d��#��m�;��QPŜ	�'O�X���>s�� ��g`�J4n�g�t ^�{fN�Cpk�s�Z�r=�c!��Ut��箊Cf0l[~��2�xz���a�����I=>]>����/s��qC��r�5�� P̓�2M�Lfy?c��?n���Mu
O���m6�pN�=����U!�Vx��{�.c,+t��g��j��૩/lOvDRCL��~�CRA~�:���>�&�I�<,WB/����,[�'-��s}B��e��U]�o�I.|�Cx��.��|dz�V�����F\M��1w;~����~a��ਸ{vX^���}a�����x�{�5xN�Z���;3��|� �%�8��xݘjw�;V�Ϥo���;���mv�OC*K�z��aR'Nf�a3κX���'ő�;�=|*�$��0��x�Ɯ���+wý��1�X�xWk~��Vr}Î�"��#�HjTs�1+X���ys����'g���><�)�y���#{ �?~�E���i�G������i�}Ѹ�y�R�3NU�iw?��{X��FX˔D+f{����\U��Q~g�3{�ϯY&S��J�"�����bb�s�,?qV�h\1z���X�.��y�
ow�\«ԣ���S������{�*�#�.ݣ|yO{4?P����Z�o��p�39�[�KnkE	yI��ѳa�'��{~���U�U���d������^��W. ouԻ��J^���U��t�_!�zRg_����+_3\jVk����8�����SQIJ�($�S�+K��x�md�v��\�|U����;�����u'�µ�`JB�(u]]��Z�]��l�����Z���p�X������t��U�}���꟬m:TXd0|*�9zo�s���tp��*��Ϲńנ���;/�v��w�He]|������gi�/�|��x���=c��03�]��%�WV#.�U*u�����F�C��Tj�>�?�K��rXύ�Kρ������`�_R�c��%y8���/�@v"�ْ�1}���U%�V:�Kj+͔p����ڊ���������DS���W*k�Q��ꧻ3լ�*�D��T��j9������]�x2�c٩/�j�w�������F��MU�Ue������pY;YB�lz�V��
��>r�^{ݭ)]���R6¦3��r�o�}c��|�Zb��2%�R���B�^Ks��s$F�,;Y.p��{.�R`�]�b�!d���.̻r�VlY��!���^�74��'[mꬷ��oBz�\��II�׊�M��`|�u��T�J��&c��g�z�.�U��� z2[���7�_;{c�:��ޤd�5,+˺f�0��a]����Q~��~��B��
˹�7K���]�K�ѣz�ma;wB�BE�ʽ��^^?2!�U����Ey�6W7j��5�j�w���/��٦+�Oj������}�1�J�fj����2�y���.;U|�����L�*�3��c-���g{N~ҩ{�|��
<����˴���٫�)��f��C�]�~�V}�̷AW�mX�g�����^f�*\�x1�;(�/4�w^���,z��u�<�.��Q�尯�?l�/�t���˗;��#�ﾪP��o��?X�T�R�\C���k�w�g܆粰R~��_G#�G�zȨB(�~���"�S��hɒꕎh�"��x i̽5�?9۲1� 'iU�� -�C]�mk�y��']��l��̛����BR�zO�e΍6��2���� Ƥ�\v�VT/]�c���\%:Dժ3y��9	7��k�ĺ�����V��>��6���^`���u��ֹ��z�}uɑ��%V���Z�Y�%�2��c�f��L>䟱�����Y�(	��\����j�uJ�V޴EvB�{N� ~8��lӳ��?����5�����㶬�y�F���Bvo&�6*��������Kv�f�=+떫B�;>Y��T�o�u���$!��/���2~�ܓ�+��u�2r����k���U�7!�c+j]�/����=��]?m��B�b�ڠ�[��3��g�%�uYJ�_�v;�t��������h�Cac��Ou�#x|kG��9x��e��=�hG��Y;b�aqxo���P���`є/����g걯��,���
<i�?S�r>����!�B��BBI%R�A+(x�DAO/����)�C�(�������<�Ο������ߊ~�	��U�b(�	HLh;BÐ@<?���?}d�K���DAO^�&�9��}9�m���D��L��J�K[�T� eU�����|4�*_=$�pH30�agba�j" �޻>�����(C���)�������uȌ�E��4����u�慗ҵ!�l������,t�
�" �_<i�~��I ��\|H@yv°.U�o�v�l�%��^���P�;ku�}�C����8�p;�Jw�B�" ��	�L2�6�xտe�KTUA=T�*��L$��4*R���+^���<�����5n7�S�~���7���T��	��p7�f�Ⴟ�qo��P����J� �5����)��*3A�������9t�,V�D�iG!���˧i���O��'�Ø{4ߪ�/�������Srr�	���d_�Ә�X2�=�M��j*�
T' �""
}�;�R�<��E�fy� �̋%v�C̾ڈ���no��� �R@��2� PR1mE�� :���`0���akRRa�.��ص[އ�#R%(�x��*'ơ�(���
�w�����"
a��~��ޛ���}z�ק@��Τ�v�R�G����g��w��㧡��O OY�+�ujd�g���)��a�r��"=>��A;��-�&%O��?#=��!�vA��ߊ� �+*C��@��uS�H����w�������ƅܳ�ÓdS����bo��%u�e�D�1i���>�� l��-N
�=�`�lR*�����=[���y�1��ڪ"
v/Q�w.ip���-b\(�m�h���$Ԑ�� g�L�?���)��0