BZh91AY&SYa��ߔpy����߰����  a9>�   �     ` �TFڔ r    �P�       P�  ��ET�����9J/j|�H � �( }h�@( ����p  COv�Μ����}�>_mTۧM�ۦN���g�}��N�{:��<uǎ�2��ٕow�h=�V�ۻX�%��%#f̧��m����f]�٩� �{��{����@p ��� ���ڱ����wXv��YM���V�j�}�o�Z2}��ڶ��֫G���r���q�Ǚ�=��_kl6�'�7��j�U�9����w;��vgJ��t��|�w=Ă�wbE��E:4$N ��� ��;L�c���E*��9�k{71��ƽ5�{��"P�B�1�t�g���AܥT���EP3@�4�M��h�|�� xX�x  �i��������&�iհ�-��̣4�F���^�R%�C|��)��$:[+Zt3��G���K�4|G ��Ǽ z*G�pSZSրWM�;�`��[-��Қѣ �m�U|K��:h��S�m��J�	��[V�jM2M�                        %OD�JUC#�Q�ɐ �4��L5< RT�LF�@bh`��JR��i `M121 F�hbh`�S�$	R���FA�0�!Ie@��b4 ��ɣH�3$BdjR��A��!�� 1������ȴ�-��f��~p��|����~};��{�E@s���tX������ �_�>�A >�uC6���������1h?�����TP��yUE .!���|�2l
/��* nH���Ա�.�P'��X�̊������A__�����_)��w|?g����Ey��[�W' �0���y,�͛����36u+z�oi���r���i��y'���M��	&��PL��3�k�
�dvIbK����Y���$�%��͡��dב2�OY��B��<�N�܉�F�J#"w��D��g�B�+�͑8�]jP��{G�e�n����!�N���g4�wU�
ȔGQ0j"o^jR"'y���w�VA�D��JD�N	�e&�:�+���N�DO_�nId�D���g�D����9�u�#���:t�۔��">�Zuꕱ-ܤN��������D��"s̯�΢#��Å�D�r�D�MJD�r�:�"-�Ã}��O�%�Ng%pM���6���핪ӹH��R'q���u0�ߥi���e����5)����5�jR%����QnV�:})�r�&��D�e'M�+U�r�})���f:�s���ND�2���$�L�%�ܔ�x� ���=+fd���x��;%��U��ZGӢ{�T�=֫Ǎ�gNIcS�ȍM�ؕC��2'�2�׃��	���V�-V��j�D��Q͉�%%�X�g]/q̕�2_��ę7D샸�{���Ok�d�ԫ�^UpLN���,sS�9uI��'���q���;"5<rOO	~j��!㬃����J��GI�A��$;�rM`�ɜ3&f�����yTn�!�C���M���*��)����`�Ю�$�u����\��K��Ҥ4�ZK�,ږw%��^��<i+I.I.��YQ�}IWrV����"z��si�5��k�]g;J�6(gp�e"H�t=Fu����P^��I
�c'%p�i"MC<!G��!�ZW�&��b/�Q�!G���}Z7�lb@�!H�*.�u=DLD_{Y�Nkw)2ȏ�N/}�8�<읳��qd��$p�x�;El*ʉ'v�ɘ��Ҩ�I���&��/�8K{GtsVB	.���N�Τt�5���O'a��i��;�n�����qC�ZOUI�,�ܗe;�M�ܝO>�{10y�&k�$��=�O2O$<�<��-��'���s����d��-�!!��捖MFMD8�RD����[�Wahm�	HZC�{��l��)*�,K����a.�]�<%'��":����D�i:��ؙ�J'R	��E���)�":��Q�L״���&���8P��Ĕ�2�p���|N�n���t|C�����ȑ:�2$���IBs`t�d�Fl�:����DO=%�d��ig��,�a	�0���&��%�DK����ؕi0��8Qq"'v�N�:�9�"#Ӆ�0H�4��H�;�L'"x�Ȟ7�M!R�:����:��Rp0D�a��I�f��i+�+�DKRt��}:��(uh"v�")<�7��:��:P����y�4��p��Ĉ��'D���d3Xn�'x�1�f�&�P��%���x�)�x�����XU�tݤH�x�<bz���t��:#�IG�8<!fj�z�n$N�z�����0�DÉI6aK#!�YCQ�9<&�`�&�㻝6��)��a$���pF�9�3�n��lnlM�E�Nx��7&ȉ�K�N2��f�*�<�G�(��׍Ƨ®!h=��&g�8=�>j$Ʀ�Mt�QRi6��R&y=Gh��erǻ+�����i��q��K�4|��F����vPLj��k��D%��4�GDB�^�]�_�/�|n˪����;.�6�ra������M�ʞ�S�ȕ�K<3��j#؝�S�nڜ���M��ǽ;榓��&�xGq0Oy��(�0��"#؈���,�.���D�SH�,鷕(G�yS[5�7u,G�֥Tji��� ��Lv���H��po�D�S�"a�M�ޒ",N�A<=�D��&Z�'cSdD�%;�B3��0�I&���<#�DG��#%�U�M�i]DN����TD���!b�%��J�TDo*'��R�2i��Oi8��<5;mN�Y�#*��wʈ�DOM��W �"pX�.�Q�jp��a��9�wʝ�������H�}-�O#2���ڜ&D�P�z�Լ(���.�>�D{�h�Q�pe�9���"�����b��6%�l��0K,�Ce���&"�P6tW�0jxk*�GU����#ʨ���>��C�<$�U$K����x��(u�5�x`��`�����9�=`�Z,vu<�b\�{��ʐ�C�D���ԃ��!нb��F���}���<DYF۩��l��N�js�%�D����ȉ�JG�DG�Dy�vp�Į5(�H��R����ga7F1*[�\�\�\�c39�E����b�B�T�:�<��E�}�}�}��� D�h�4z�=m�����8Ԅ�!�k�׸ױ�u�u�" n��uUn���{Q�}ꋕ)�D�G���̈����㈱Ї�е�	�'���!�L�'lM����w+�M�'���3�8�eY�+�-q��4��d(Hz|�����>�+q���I+[Gq�,Yed���5z�U��x�q��Q\X�1Z*�G�����t^R9~*�f��)�<-#�z��N����+J9E3w��8^��X�x�pg��4A:.���G���H���W#��M�+�𣏕��|h�r9��35���H��e7ȰW#���{ML+����W5Ү;����z䈝d�!�#�H�Y^/&�Ա\��r%�&nR&>��J�$��D�%"L.���G�rWK�:})���gDG&�
#����">�C�MMf���n�"u�D[���+N�JD�\�	���6���핪ӹH��R'q���u*poҴ�ep��Q��D�r���Mf���n�"u�D[���+I�ԤK����{)8��v��iܤK}):'����u0�e�����eX�jV��I<W$��C����T:E��2Vd�D��'#C	�		�6͎Z�|�7�WNI���HnDJ�~��/"C�����!�A� �� ��Ql��j#ɱ6�R,�3]/q̕�2,�.ɓ�NH;��u���d��N듯��&<���窒�5<#�T�'���A׎�N��;s���Uu���Y$I�Xz�:Ld'rA��\G$j{���s%fO/�=h�hބ��N�0�G�i � � �\RO�'ԓ�+��rWZ�z�$�$�$�$�҂�v%]i`���@Ǝ�[Q$�Iu$���5ؕ�%o�ZvIG��;G0���Xh	d�=F���!2z	�8L)�}���'5�;֥��rp�U�:!F2"&�J=��3.}�f[o���&�����g܌6Nl����|8L����F��=�i���Z�kWV��PumR?�#��Ï����\�=|��_�f k4�Diq������@]�tO,�1,�[�
5ն�J|�ӛ�$��#Ǐ]wVI���%3)�:n
ab���TQ�Q6x�D	J����h$`�l�]��
Ξ0�%��11���Σ�O��e�p��͜,��n��,rEKmSg�
%�F(���8�*�:Q׬�����������t:fi��(�
���+
0��[���;��Ėwq�����!��Хd��*8f��^5��U+�~�vn|�/M�/5�U�#zۢ�^�Zt���d�7+�p�ҷx$]JGs(�����A�Kl��y���v�<B��j�zn��͛�	v���u˺�ĝe"�7��Q��u#
EQ�}�.[їh��Ŝ(�ô^ʮ�:��d��E�{�L�46��>ۡi��f���Αz�-U[���6�N�ʪ:I?k�:i/�R���0�|���s���Ms�۳+�]�tzi�g�8l�IC2��l�6XxNk�K�]������-�wNr�a�م�fb���V�2pj�p���E{�'��������rr4p��>��:@ �+(+Z�b�K6x�iY��9x�#v��K	���mF.C����Tل�\jL�¯9�v6�N����mL��F���ad
ָ*(ɯh�$��W��s��Ӆ���[���Th�$
�FΕ|��g]Q�>��xp�N�,7m���!����h�e3P��iE�<t��0��Nh�Q�n�)��m�v@���d�,�l���^㭷�J&c͏�Я���rf��&�/f�(��3]~k�~~>���Y�����G_?��I8@kE�qP�O�2�ףXac8f'��zEE�5aB��[VVIҍp��2a$�m��4p�3kP�Q��(�G�����Okt>D��;�uaG�:_GXQ���B�E�>0������x�*�9�}u��ۤ���9Q��D�>Y�-���c���J8|,�҈�l�l��_��S[>����k8�υx� �ʧ��a��φw��� WM����Lu'��yc�uyngN����#)0�Q �9��5A
)Wi��]Z� �>h�O��g��A�Λ=HQ���	8Qq��@]Q���¼,�F�6�jW��,�᏷�OP<����e1u�� ��8h�ϲ9����P���Hb�Y����v@a&>Yy��:���!��^S���=ӯؖ�AUFɽ�x�d�	�LM��u�O�9q�/Wv���y��8GZ���Fr��cv�����O�����]wX�wf�ׂ�p��!T�s �A���s�~����H�{���]O���,���@�^d�.�+�~uS�z���^p�ϕ�G�B���0��0�m�?n�4P$��¾^�|�������v��M�g�@�$is1���"�����*zV�,�[��>�,,�����eN|@�*��q�ǈd�%G����IFϰ����rO��)����FI�XYZ��:�\h��4p��&Ʈ�	�����;�Ӗ�04�%�%K��
(�E��Ӭ���Y�'����6h�.��S�J6h�g�Q��d��nS����s3��Tb�+#���櫚=�F�X���x��h�6B�^�h�O�F��h��a&^s�D�GK<]GĞa2 �F���k(ɡ�0��kf�t|l�[*֭]p��y����1X�㦏J�J��n�ƃ��3e6l�&�>���XY�GCP��i�Qˣ�k��Z�D��,��ٲl���V��H��=��]6YR8t�bK8t�x�[��ş�|����E��8h���(᪏�����l�%�ܵ�+���G�^��e�M:~ b�Gk涝4j�ȍ���f�V��[�g���Tv׎�=}�H�f�hY�i���i�ĝ4aG�m��gI4e��m�NΘt�:Q��`��1o�|���w�'m�4e�Ğ&����9��)4Y�e��XO���^�t���\9vce������>6c�J�tI��}���6O_;��Tj��w�.�^>��}[_l|q�.���0��va�UTyZ�W�^U��l)�9OU*�;N�6���}+F"p�\U�G�Z��
,k~tɁ$�'�SF��2�kB�K ���4f9��$i��<�d�$�S�g�y����{)�e_8p�NU<9�B�<l�g�>6x�&6Q�y�Oƪ�L?_���(�I'����%\����G��:p颉���2�0�Ǝ�h�f�o���� oj��F�,�Z$��g
4Y�Ǝ��Ƶ]{��䯪�o���ֶh�N�=AYD�4Y�F��#<�Q�I0D�Xx㧥�I��Nu׮��l����|x��K(�יTnݒ]�I(��{&�V�ke��zI�͊H�Q��	o8�0�Wv���'g	�r?�I<t��a7o�)���Xs���(ћ5�8a̾���?&��N�>'�S��]�K��:YG%�b��3�q�ۜ��qٸ���6Q�O��U�K�&Y̧ƏW�MYZx�Ea��ʅ��GVe�5���۪�����x����Ƿ�7Z6Yg	4a�ɪl�F��3�Jus�m��l�Sަh%Z������gV�tRf��z��f�p��h��w<4�J��e/],ä �id�6a��4��m����zQ�<u�p�y{}Zz��l�J�$�g@���k#���<Q��Ͼ�2�3������էO���ePH�ʙT�8r�� ]$a� �Tx�|��_S�ü�ӧ�3�ny��T����O�^��eܣ��N�p�ƍ�0��7��n9�\h��v{����vn� -5-]W2�Z	Ⱥ"�TYFZ��8hZ&�W�:�c�}>�!� 
K�6p�}�aˬ�zr�A��V�ca������#�f�8˹Gw4�Q�Q�ϵ̾?X�F���fR��ӭ?���C�z�K$�Ν����άl��H�~�gv���={7��ꞽ|�����%�ˈj n�k�9�&��|ř�lf�cx��g��ld�[9���k�+N8wq��vI��G�����/d78Ъ'J0��d���Zt�F��Qǭ6ܺ����8�M�6x��m��|Џ��t�F� ,n���f�U5��كVX̝���{�P��B�����Q%f�t���2,��(h�y�&d3�U'ω+�#�`;��2V���p�Ҏ�\tن6@R<IG=���p�T	4l���4y�|6"ID�W|��K.6ݸI�����QuVUc��$�Fe�AQ�K4YD���<��UǏQ:޺�5�T�D�Q�����F�>4m[d���I�4p�����ͽ6�Ҍ�V�nV�Xju6s�	Ə��es�`Y������S�O�U�4I�&���r�/�=5-�	P��Z�uֽuΪ��lO��'���ѯg�ߞ�}��������{��e{C�{Mf��~��2d��K����t[u�v��gJw[���J�5�(���H�1֤k���\xe}+v3I�����W���u�d���k޳��1u�C��c��N�KsL�J���ɰ��ǈq�1.�fy��38�ᡑ��m�ު��놈T���.er���٘�z����د���F�І��l}u�D��u�3v�;�����B��CF8AvjF�.Ia���f]q��g�����tcmH���	!vV2��.�u��9�6�R�m�"�$r$�{���h_z��JK$z�:�p�wX���m�Fz�4q����.Ad�UlJ�)��m1s�K;�t�?�'�,;r�8�)$��Fj����7�&G��W�EF���A��+R05�X;�
eFSnn�W�R�#�f�A�D�M���ާOH�uX��r�#%^s�]kD"[
���7���-�M���[JI�:ړ:�A�lГx�3Y��sن�ˌ(��+n�a0�&Q
2í�z�Y���4]O)��g,8O,P�5+S9v�=׉[!�GZ$���5<WOSH�����vۛnʒ�YU^���f/�V�$���3�(VjVD���v�9N�����:�7���6]k2r�2��BӔ�8R�J�T��V���s8"�uh�ͻLN�3#6.`['1�+�	���f���k�x�d9���u;q�G0�0��ĥz�W;���F�;�O;�����x�f��a��L�F8w�����H��ex�߭lB�uу�/A>�-�M\��:%����p'�8
o��y���AsrY�q	���e���g�oz��XRo	�u+��H:��5�J#Իq��6��ky:#���!]Hu�1B"��z�깙���hT�aƃ�8�� y��|~h]�R�T'�ԇP�`䞹����2k�}��Z:��a+jyף��J������{�EU<�w�=�p =��x:#�]���q���������}��M\4~��!�*�U���������U��U򶪯U�U_-*�v�*��iU_,UU�UUTUUTU^*�UU�Ҫ�WjҪ�EUW���U��W��Uv��H������Wj�*��V��-*��*��*��*��*����$D��K	M!�=N�	R�KI@j2X�D$B���r@ bD(P��(W!B��J�UEUUEUW������j���*�v��U⭪�UmUz�*��iU_,UU�UW<�j���V�U�*���U_-*��iUx��[U^������U�[U^��T�*�������U|�*�努��:֤5�D� kAH� m�,IJ�D @��B"PP D�"P���B$JiM�7j��b��,UUŊ���*�努����[z��U�U��W��U^*�Uګ�[U^����Uv��V�b�Z\U�*��*��*��iUx��iU_"���Uv���U*��U⫵W���]��v�j��ր�A&�aR4%%!J9��Bά"hH�)�+A@>HT5�B�7/wϾ�︪�U⭪�U]��Uv��V�W�UqUUU\b���U_-*��mUx��[U^�����U궪�Uڭ���Z��b��"����W��V�U�*��mb߮�j��[UU�Ҫ��UU�Ҫ�V�4�5�`BдP�@�
�������(�@4�Z3�R�)j�)
)P��#��d�䉐�z�P��Щ�F�hF� rV��V �NӴ&H�FDBg8���@��R��R�B{�w���⪊ A������?���8�C��~c�|��|M���ÇO�x�C�DDN���8AD�8"xD���0���6 ��AĲ"X�"pD��xL �xD�<&	�0DD��Dᲄ�!B&Έ��'� ��A,؈�:`���6��:pK<Q�D��D����(A�6""`�"'����x��6t�`�%	BQM �!�,�$(D�8$gD��Ǐ1'H ��"'O�"`�8'�	 � �� �;�~���@,5�D~�����u���v�;KڕL]G;;q�[fն흆X&�f��r훶��~7�離*c_����f �APeXL̑,�`[�f��e�-v�X� �Z&ߓ��k��v
�c3]��ke�B3GvN���װ�\��-B�C2�R2ʋ6�s��l�`	����s�!�g�m�֐8s����gf^�⁦
F&9�K�i�=���mB�f5������ʞm�lե���V[�1�$!n��]oIYm�|po�s`JG8���ޥ�����1̺:�߆�m=�m�r"^��6Kqe��������ηF��vy��c}ͳ͡[X-��l�z�-$e��h]G�������Lk[���m���SMkٽ~�f��S%&�Fʪ��cE��Z��iPis��x)e�I�;Ki��;�Sh�K4�M�-�����Hb��m옥�1��Ǽ��[
*&�SR]#�8Y�웿Yb0B�r�w��Cm��4��b�	��gm�f,�u"�Xi����ͦ��b�o�]�y�:$2T�"����={\�v���֝�@��]?!v�ƃ��SVfi���(x��<b	�ka�)lлM��&�����ZͰn��k&Ge�L��ec�eR��c.��\�%#,�����$�e�GUJ�f5�F}�_Euv���m��m���۞��C.��`�-�k]�6:��ݱss-6�G��v)lI�)��csh[P�Z���%����f��vn��l��U����{1����nS��Ŷ&�ڷ(�mh`&�v��B�ɽn��͘u�lcKcm�۵�&j�[F����m5�l��g:��z�3���P]K4�6�+� �n�5��)�ap�=U_W�$(]�H��k�FQ��=-�К�ƥ�LA����u�VX捌G!�TKun���M/K[�VbUf�Z�a~�5��ކ�c]j��&��5���6�Y����m���ō�Ø78Wn2�,; �`�mpCmֆ�^�Z�#�WPl�m���<F�ikc̃��]�&uƻ�GpmF��f�5e!�J#�WV���+�Q��
r$茕M��8��]�761����Cɫ��6����3`�h��1���H�e�+ t�$bYsv�Y��e6�w(��q/7^�2�5�A�8Ի
͛nGV�x�����iu����
��]�8�eh����Ʊ[���$�q4�{���lMu+��tRY�6�8�#1W2�l81��V�]I�Z�8�ɬ�rJ���6un)�Fzٞ�yj��\�I��kP���e��4en�q��֭5�⥷L��Wޙ��z�V��n�Z��fͮ��B�Yt]��_o[���ݲk�-�`m�JB��0�Y�X�3v���e��6�̒�WYrZ�����[��qWE��Z]��ͤ�%�5�fV�f���AGe��s>���=�6ͥ1�-�3f���Y/�<F�&!��lѮ[0A�%������hj�İ։eě0L\�e���С)e�bۍ����7-��0њZ07M�7ﷻw�-W,.�Tk�[-��&l�&��zm.�hin�l�����1"�)�����W��Z6[� �+(Djj:�0J��]����iKk]X�%����ݻˍi�;�*p�9G\���㥚�U�GVXHB%���4i���E������$�T���Ҕ�MM(�m1H4��Ks�u�lų��
\�jBm��m�5�Ymae�9�V44ڶ�HZ]�ı�����4�;6F�(3e,Y���͓9VUk�ɋt��ꪲ�5B�n�����45�&�QU�ig׽�+�$]��ޯ���6��m�5��og:���g���g\���t��۝����Y�S-�C%�z±�Z�u��q���pJk2��Y��EX�d�;i���)���]��m�
��਺3��!����K5uֺb��Ț�%hJ+�{�~~�EUW��{�߀ִX��؊��1U���������������{�ߍhѡb��b*��*��������A����I4�J4�Ş<{�����0pѠ���z���D��a+͉���!fX��KH�-ƍ!H���1��:a-�Y�"��Ja]n��E��mK�F��]{U�@������.���CI�"�k���Zg�Ys�-�AV�P�]&���ji��-p6���؆�霥+��uly�v��0�uf���b�1�^�R��&��&K�,Y�H���-��lW+�!*9tyXMjԺLE�\��V�v��h7XoN��}v��bh��L�er�VQ��1�����W%�T��1hl�h;���7Z�d5p]�P�7[���+hqnq�Sh��z�ֹ
�K��f�D�3s6��c�`)*2�A�u]��ٖU���噐�`T#�ZCE�u����f���` �����nF�>㻕B���Xڬ�54�7b�ey���L�g/J�34<���-I�wdwAo����IU�m��:F�õugr����B�	Z�Chj�{84ߑ�=D���7���/�A�����ae>�E'��:�IL|�m�3�&ccd��u�	L�r�i�Iβ�g)�.(,�7#)J�m���ɦ�/��g�nttt<��[m�Dp�b�yi��<{���Y���$����!'p�$�O�����&	���a�<t�r�����d��C<��ܧ�I$�^7���A������2Lᘭ/�dw�qيI��F��@����@?!X����߈4�$kM$�E��J�Y%�P +�	!�,&��nP�[WD�`ݕn���"�p�Ӓ_IPC}a��6��u�NX���N�`GH��p�XLK�p��y��f���B��;,M�|tDLf	G��x�c�Ep�rK!:���ʕ�%*�z!�d�{�H�:9dȕ��@�
"��9�%���\TB))NE��N�@��"DΣ�m�EJ�Klyz��e8�<ҕ^s{r���j�;KȢ3;��p�h��g ��:�K'��i+�t'�.P=\ � m1A��D�#��-�h���8�ѠeᤘIet��<`�0J<&C�K;�_n�e���2�!���gcm?t;cQ��cO�
T�l�6,�f�<e��d(D���-�IN���)b��J��u�;�<�z"8<k9cR�*�3�V�p��:4�e7�I����|��m�n}�|��tz}��W~�ĘzvA�h.��,h���g����S�^��E�x���9�QN*\�!bg��,��0���D�0���a,�se��;vm)A
��(�T�Q�h\���ާNLߚ\{����a�����RFL��p�I#*�/���.r����b�N�[�si�<T��h[4�sqq�X��p���S]�(�W�����nmX�]u�4�Ƒ}�������9��P��\��u'JJ�v+<-��S�9��p^���B��)�'��:V�-J<t�H&�D���%p����U$�6�M��½��Fx�4zR��e�)W�9O���CGU��ʂƯ4~��N3:���#<�KNKvժ����GM͛n���]-�'y1<��Fzy�Ȇ� v��|�(��0��0���0L��0�:Y�1�m��^m�V�&�Q��}���Q�2��Z�ȋ)^]GWFZO�夒�BY��x�s��C��;/��䍍���)Qv��E&�[�N��8{��A赝Md-�5�e|�cm����uo��G� ��ڤp�A^�|�˒L╋���\t8x�,�g��'DD�0N����NΊY<��6��J�V&�p�0�����I	 �UR�J%E7��y8Ȫ3�&c����O
 |u���x�����QB#:���KHRgd�LDqP��cl���z"��yW�!O}�ʧ��ͻc��h�IA8�9��漏��3�ߒa�`v��������-�1b&��	b$�u�"d��/�>�z�N�h���A�b��2Fad�Iҏ'DD�0N���x�f�����cav�f��US���9��y���+�)qa�"፦�%|~qPB�D������*�f�4Z5*�������8�t�JX�R�cHa&J jI<3���e�vu��
a|�^Y}��]y��6�g(�@K�:�N��L��0���J�:u�<I�K���A����Z1�gZ�3Œi&x�DD�0N���x�g%���ɐ�Зe��bY^��HaÀ�	��1+�����!��Z�d�Iv�~�\C6��P�[y�	wX��m<�٩�^�����­@�̩��������Ё4�s��f]����q�C-8����ٽ�b�m�:1�f��,�`�`�w��oI��%8tnꪉ��yڇ�\>�5��R�gMT��=�G�8JBh�A#�A���H����20�e
��u00UD��I������JD��Bq�D6�ƪ��F�^������n�EM�4R�93��Y
HϭW&ڱ�튖�XD�R�=.	��oXn8b	��g<l�tDL�xL0���u�Oo�]1��X��USp�8s�T��9��'B񄥢���}b+!����_���ܙ����:�P50�0�ޱ:Lc��`ъ�X���GL"x��0��1�o����/��h��:��sRډl:s�w�oZ{����Qr��V�ux:^h��1�h�TQ����Z:Wm�a�?�<��Ռ����!��N	�z�U����c�4��M�������,�zC4��G���,�4}6��z=<BӰ�fxra�vo��F�g2�<j|�)�>O����Q���D�i��(����> �j��Z<��H]���<A����G��4v=<A�<=� ���<>�F�"�����#G������z?L"�zA�M4�,���4vx�m�=:Bњa�ƺi3��C$�����n7=�����z=$�tzY�Oh�A�����ޑ��FA����
4�C�ɤ>��#�`��G��DO�H�A��8�	�HU��O���'����>�$Dnx��a�0�zC4��F�H�H��z���z=<A�a�4���!�CF���#���.鎉��44�!@��������H�ӟ��",�;�8jF������b7TR����j���ʬ�Qů%Zb�'��eV�h��=��h�Br��D4���f��D�Z��W˚�;�� �0�[a�Z�'�o�cZ���	N,��bY��)��в���]l�d,6��_sѭ_mؚ�"h�'�Z��&jV�˪�}�\�g@U�A��芪+�B��9A�������+F���t8Q�l���Xq�T����s�����"�����5�̙�������|��*�ݿ֌̬��ϾϾ�}��+��wv�h]�c��{���{�������陟j�:C,��6a���0L���OD���ߢ�Z6��$���B��9�6}%f̭7o�ga\:�7?���$�ٸy�"a�|"��60ݎ�=8@Q`Z$�y樋�����;c�Z�Q��rI�&��L>�Fۖ �M�C�NqӞ�AJ,^?6�KdRz,��#|�|F���:4!Bs!��<&�4�<���#�$���!�^�N�D쑳/���7��n��Nyp��u�T�*!BV�tb>�+;�n�x�"�9|(m���|2Rg��B��zIu�}i��6I_]O6��T�3t��||YӦ0�g�ƞ���N�>9�R�vBHI	��̘h��i����q;��6�b�H]�<��kF2m`m�';QQ�S�~q;őR�~4���2�ѳ��:�	yd�"�iD4C����}[��ɹ@<^�Q��K�C,h�zH����/D�'�!8��˗m��Ot����nTE���K�L�G�m3x/ѓ�Q�V%�7�Ӳ�*��4�&f�w�Yn�D�D��.�cm�l�&dl�n	�ӭ3��3�HýR�0���T޴�D���Q����xr`P�4��Bj�!����|Y'ĝ(O�â"`�'�|"C<@�
{��a�F5NSg��5Z�浕6��s`'�q@����Ͼ.YF�ǍU@(�	4C!8�*'���N�I	!$!�7��}�k�s��Y��¯�oLa\��6��hE�+����Z������,��fZ�K_Aڬ�����uJF��	�(Y�V����
�ȼ��V.��3W���{C-j�6�E��_>��+��&��7�Gc*���pZ�c�#Drɢd��=a�;��G{5��ɀpA�!�t�;=O1�A]CT��lJK��xh!�� d�뺴i���12L��N���Y
��7;�p�;�)A9�G:R ����S�6�]�Gxt�boӡ�^��$��$mѾ��h���u�%ÈL C�&8t!1:$<5���\�i�$���� R��F&y40���I��1V[�?o_Il��������8�Ђ�w�
!�~�ȑ$�}�A����u�A� c
$f"W93�J%�`I��|I��|i�g�:x���GÂ�@�el<�#���$����3���� ��臤�Pa*x���G��,ѤK ih<0���4�d��)�{�W.�`���'�b��"R<��D�4z�plp����J��!�<�m�A$�L�]o�Y�; �`�.�p�ܔ$�m͑�@��+2��gB~~�4��쓻y}�[u�,ь���#XbhP4��Pዱ�WQGda',9˯U�h�
L`8$8 �S�C�nD��� +�$��1�4��\��&a�y�L�1�C�y%9c���aܦ�8 �h�l�>,�����tDLǃ�N�A����!�P��S���wi��~���@�a?\�d��L�j��D&I�;_�p|�p>5f���0a��F��ø�Lw0761LI�N���	�ƹq�� O"�!p�#���OJ?t�@����p�fk��/���A�$�lbA��zI�8`�-.wq7�C���OV���Қg��<_��6/9y�K4����0��������}#��&.�>nyo����4c��&ď$&8���<$29'�7�0��� a����M�YjN&���p�s&Q0z}��e�a}þ�3� �=hW��y]�x800�؍K�d��J9��*�CY�tk���a�&~?��<t���:t��I�ۡ�aP^��e��<����������@�a�bdH8��>��0o�y3�7���2D�ԣ���Cx\=(�18��~O�Y�Ge9�}�: �p�B[�����n2��n8i& �H#���p��79�}�D�dN���؃��t����'s�nvC����;��� �dF��lGr.�(e,P��t`RY�[d��#%=2&%A0�g9�����n����UIn����7(��(_yA�|��i4�z[d`���=�4h#Dh�L9-'F��nBv�c���(�#7��"L)��)��!��'��6$1�!.&A�$�G�D�,�OiQ��k\rK�!���Y�?â"`�<a��M 鄋j�K�=�|��q֥��#�nܖ�2@V+"�>�B^Ag�c�K�Q���� ��ݢ6�D6C��mF�m��	 �ȇP���s�ߋo�r��ſ��z�~|O�R���ݒ��黲�d���Fޙ��U�}ܬ=�l�f} '����`��^L�,��f�7g�%�0�ªp��&�{��qV�bSd�L�8 �!pK�/	���Y���Ө� �%4L7\ �:������*K�#TH��S�`pK�N~�%Eӿ7U2Ci�wvL�F$�z �!�_���ʖ˲�2�C� ��Qۆ���]��/�M�D��!#5r� g4o8<���R@a�S<�Ai4��u�p�&�M h���z!&Lcf=!�"�I����Ý$7�(\��D&<�/��X\�U)٥T(�I4w�8w�搣��3N��CQ��V��C�9�e����d0�,�Ϗ����0DO<<>!��L��M��HCd��<���@�o��@���.0���]E��&t��c �B=9W��<; x!�~���6xŖU ��0�#\"ț��\*HAၥ���:���Jh���8�l�hP��|��-��mߣk����	CA�G,�|yP�`V"���9�!��]��qd�6�7M������\Y�s=&{���^֜��{�����J�âV"~L�'I��VAr��@p`45#Z�J�J)J9J�!��\YY<\_xq�HGUAki�0e�I��4��Ǐ<x�Ӧ�t�K�}2�n*I8�r+���t�r�$���>�?Rkl�)�u6י���
\���_hΑ.�>�Q���w�,��Δ�#Ƞ��2��n"&�#�URae)
����q��	����&D�v�Yxu�w2��
�Gd*���$$!	@���)m��N�J::��N%�b�@I�O�x�8�Q�>%��E ���\8�7`�Mv���1)9c7֓xx0-3��"B���Ւ����D�Ї�C�����6�M��9��6�5~����4��J�_4�0`J�T3���!xb($��x���	���:"&���C>(���w�K�5I�0��H�r��	 �	@���٤/2�{O74?d���F�(�R���8���6�˜s�&3��>|�[Ke�p�u1!lz�d������a�ǳsN�qoGhߗ�%�ta=N�-FJ�U�gC" $am����d%� �G,xuqA�X@µ뷧���O�DY���e4O��N��D�@X��lG�be����{���Ë�ή/}��H�+o�#���,a�i<p����y݌M�=�i؃bG6K��{�:.�������@�@���!x����wR1
�Ad:���bi�3O�p����>'�֑��0֑���:F�G�NK�4l�4zI��f����ޏ����0��!X�G�Hc�f�٪�����.�#�=��G��pg�T|B�g�2��>G�јiFh��x�Oig�4d�Oi�?���|=>#Ft�(��?��ГO���4z=�������A��Hєi�A��#[v?A�3[��4�8A��;�f���>�!�A��n4�4z<4��#K �ɡ=4�4��GG��h׍ ��4�8=�!xzYp��Gᣟ␋�;|�G��ES�*�O�)��"F�f��cѨ4�����=/���Ƒm�6i=$�zF��#G��������Af�c89�E�Gm]��5v�E�Bt9�?Q�B�s�W���W�7n�1�a��n��I�v!b�|큛�!8�N'��r%#��3
���MHG�,��*�1B&��Č� uwG/G��EB:c�"�vED:Wc�)9�+-�����w<�v�͡��B��Q�;��\��f80�I�j���]Dk����\�F�#�c(o*`�v��U� ���W9ܥV��u吵[W
}ʀ�*�:����͖�3W��.dMo���ɳ������sk�A�����B�c�{�n��-�F¸S�U������Vb�j�g�Ԍ5�ɛWwF$L�pđ�T)�kb��\��r:�>oM�C�rϞIwU{B��#I���cr�qB�	��%�kK���e�rՅ�&��L%��X��X[)��y�]i/�}a䊞n��m��Msº�"�<5��`f5Q��Y��YGM����ď��FmY,�B��ڳ��ժ�!��� ��g}����7www{���L��R�{�{������}��g��-���y��}�iW�{��������{��v��G��{۽�wvf��ѣ!�afp��舘"x��јi�V�x��0��7U�*kl��9-ͻd��\4��H�ɥ�[ �fɺ�4-������-Q�����1ֺ݄���Z�L�
TR���2�]$d˵�"[l��f�;k_���/��.��5�f7`�<����W�We��+v�R��rC�ޞ�6z��8 ��u�6��W9�5���kU�c;KMq4u�����J	R[q�sL���Zy���[[��&��D����h������m,iV��KkM�-�v]���6�i�6�&ל5I���%�=YE���.Ś�ö�)pk��<�GKy
͹�����p�5�y��,�R0��m>����.a����LWv�XKILM�%�)��eЬq�(Sl��a���si7d�����|c�1!��8}��t�B�eE���[�,;��q�7�Sx�H���l[	����;�yp-Y���.����t���E�7��{�����,^�0���	��Q�3��>��'ïE�Qf��>cI�a	�8����;�j���ù�A鋀c;��tz������H$`B\Rj%5��d�(7,��2!~���n�wn��wh���4���)6�Q��7'w��Ѱ�{�A��t�ÛW*���05$�rx �Aԛ;��1�-��D�s�1�S����EH�"�hA��~˚y�2�v{��{A�9�g�p�����C�o�wa.�xX�E�Ss�ϰ�|7�>$Lce06 � ��(���q����s�/B<`�0��O��:"&���C!���<�L}��ݱX���$6�Ϭc� ��ٰ<L4�q"gt��uE���F����Ŝ ��EP�>�	K�`�*V}��r��I�?|8o�O��
W�nIG��$h�H��a��<�#�x�1V�!2J���iP�h��
8��GF�ᭌgW*G�]���)��	����{�#��8�}���FK��~�3��/Q5��{�y���8Y2"a:��D<���H3}8t
r�2[�%���B�"F�Dj����'RJ�0X�D!�HZ� hh;چ�K<�ål��A�H�,�	><p���O:x��<3�A>ʲ	�U�y(b)VT�^l�b�C�:���~�.�1�aE ����QD�fHo���xx�'}��i	��Q�R�Ba��J�X�%"Q�+�e�a����v��R�L��Ѻ9�9�a�*x``C�n�v��f!��yq'���2����KN�Y���Y�Bo	qQQɑ����������"�I-q��ıL�x#ĥc�W�qTWr���=��8L�!04CJpg%�J'��t�I��]#jH���u��b�"Ƒ4h� ��*�c�ws�ge!���t����A'�r��te�4�!�%4�,�E�-��f3K$������4�㧏	��C!���3��ww.��*U�YdA��茖���ʯ=8d��G��=vPT`I'O�VI;z����K��Rf��l�F�5-49�v��YqA���$c �O!��u30��x%4�G� {��@�$j2���8��SD`V��&)�4�M�M�\��I1�ba�5�Ƹ�
D"���o�-8�PC�8��!��
����vD�F/	m��$r2<$�㌮4���GFbP�f��0�z���S�}3Á��"-9It�nBm��I�6LŏI���#I���H`Q|x���p������"x��x��
>�+�:U}K�Ϥ'*�"���4�bl>�������c9l���W7-�M��ٛd	c��^1�c���7�����道�VM�N.˥i�;u�ea�5�fs�v�cʺg��\�%1M.K.�]�������fooQ��=�]ʿX{޳�@��p�Rx��<�}G��R4����`�·v��;�j���R�hcA�|�!�	�~p�s�N�7(��}����1�'r��&�8�nJ��bS�����s�2g H32s(�!-����o�퐙N���8���fwr����ƒ0���옡��IUE���d<۩�gc"z ����� �$8rby��4B��q4qU'h�~jդ�p`Q���g�0-v�Dtg�ܟO�(��0ba0A��\L����\ɉ�R�Q��6�e+)I�!~8g�G���r�����]H�|J���:j��4��
	0��Q�M<p���DLǄ�C�ǈw�:���˰�v	^���1�A���s읖�H@��	�#�a*����Z�8T��j>���B`Ãp�}$G��!����9�)���! ꅤ�m�+��X02�@�A�T�R��Aɬ�	x �� ��
;��U\��J�FyA��j�?(!5�>M�X@I.h��7�ws�>���KB[���tN�a�s'x����]�(��
iD%�"fp@��B�/�`<��K.�=��I�CQ�Gtk�2��/�m��e�=9`lFɱ�%�p���^~�Kl�ko��g�� i� �6%����ç�&���C!��={�$�uɗr��K4��c�!ף���R�[�~�)�ݹs  @��Ng�ϭ��C}S��.�ė��{#�p8%=a��A��h��!B���x�
�ڄd�9�FBltJ%t�$��"$��~��e��.���u�?~�vjj�j&����u�.��Ȅ�&�6 �X9�FiѠ��\�l�	K�I޷��7�P��P���A$l�3�m��O�G�gO�nHH��(��}w���k������s4CpC����A��gY�<����E"Fp-3��	CG>$$b8l#�D��!��q*��ۙ��upd�Q�&�8||Y��:x��h�F���mߨ��i4��"���Å^���1�A���4Jd���q�\P�`_#&��������=��g�l�j,�I����j�\J�k(���;@�H7���ը��(�������'�U!��Qn�i�R��F�'6�0kC���B��t��d��hU&_�ڱ�G��U���%c��A� d2��Bj$��8XZ��y��0�jy5(J�IC��'�(�Y�%)������>?R�.��&�!q�gZ8j�D5D	:3�(��O������0DOa^���W9n�1��P^��e�!8��)�Q����X��=�]�/�����.�Mde�[a���>��d�P(�}y,W=��g9��ci˿e^h3��vu�,wӍ霷.��S�[!���������"v�af�|>��"q/���hb�����%�z9t�H�� �c���;��M�rō��o�n<b0[D�&p��Y+�-|�4I=m��*] �l��)��a��؈�!�|O�墇���b'��T�:8\p�d>;&q.b�38R{�_�D���$���n�x뚊�%�Lh��NζS�qy�X	�H��r�YXHC�B-3��F�� @���"�z�|�H"-�0,��M�b�HǧQ(�4�k�JX0,h�J��d%j<I�Ȉ��[c~D
�Ō�FYGO�i�`��<$0�>*�+UA�\��nI��Ӿ�=Ǐ�ٻ֎��c�q&��H{�(��A�2�aH@�gC�w�>[D�NT�B`A��C��К�m��cI:�]����b�clpIG��K�o���ǙД(���l)��������DIṁĚH$b��bE�<�J8�Tg���>��0�t���b����.��L� A����v]��[�wrl���9wO�\9�[G%4xixi`F�aK�I��`���>��m'Q�i07I��y�fp�y�{�#cCbr���-����<<�4�ǛTU�F�KF�	�c�a�nI%��x&�4����?��������(zL=6^��Ӥh�~M��`z6il94���#G���m�z=<A�Xpvg�Z.��&;0�ڻ\O�G�D�s� �9��L����p:�����>��3����5��<C�#G��z84��4~4�Ƒ����eC�M"M$��24z3G����=�h�4��јl7�Hѐp�A���Fi�|3��,ip�#� t6x���#�H���{��M#�ӄ@������H��da�4��H4~�H�i��B����
4�?�h��_�����G���X��a �9���t�4a����dB���};/�`�a==,���F�[�I��vi==a�G�����H���SzC��D�Q>�~"zO�D�~9I����A]��V;�_� ��[�V�4�"w?fй���PvS}�:�wM��ӯ!���H&�V�,��ԵL�N�޿-&li��.��,Q�]�1ir򌮹�ݻ5GF@�D�Wd85�0upŞ:E���^=�#������UU��Be�����]`936�-��t��Q���Y�o'F7�'�$���O3��|6m띄3�˸ҧ������Ͼ����{����������陙y��}�iU_,���������f}�mUz�~���������g�qV�W������!��6a�8i��i㧏0��:tfa�EÒ۱�1�c��A_�	Ԛ�S;L95�$����w��S�68*4��܃fn�I�9cAcd���g[Å �!/2:I7H��no�fy���`�p��'ȨGK�]�"����N��tn��$��a%�/A���.����ӄ82i��6%'F��I#�#�(���a`��A���&�Ǽ4<�]`fe��.�t��>h�"^:b$1��J�C)5v>rI��s��6L`���M��;��;�j�ԧ&������ �;��{�ULi7��Ò<w��,CT�4R�B������PQ�>(�E�t��Śi㧏0��:tf&N�'P��\��%�!�t�1�d�A!ED�O�蹢��]y�{��<O���M��)pt衟.B%�!f��#��ҡ���&}GK��a�$��x�x��fb��P�џ-�����Jl#�i�م#���<y�ߋ�a�gc����ˁ�>��'�t�	0������(�\9פ'S'���A����f��wq6Y���:�I��)�8�x�M$���p��(���$ns�h�s�*z6Os4rK�6c�D����6x�^x�nDS
��!Q���0�:AK
R�����g$Tpfp�J:|p���M<t���h�FzQx���ې�F����Z���tg����Td�A��b��ֲ6��s����8���Ց�mѾMkfw�H2 ��̻s�$�H$�!^��͟%����k�)^����!��֤'��F�C�/���[{�h���3
2���]��-�Im��:A���P:����,�=1w>�>�� 3[�O+�Px)��<�O3/Fe�N��f���Ӥ�t���b��[p[Q8� ir�R�
��HN�IH�1A,,gv��$�q�рȯ����8p�2	q��pp�^h$!м>���NJ����)QX�x���T��J!E���KJ�j���e+9t�+"z��b8HH�b4���ғd�y�� i���g��C<%��D8��"����F�G.�uJ��#$la,�L�n~!��(�8n�O}Us L#G�O���$\	$gǉ0��Y��i�O0��:tf���۩S5̎0��s�<���L �u�1��ɤ�16cst�96Sb;��#�I(if�T)��;���ˉ&��Z�����;E#�V6��a���\E/�>�H��d3�G�"�6"t�Zӈ�t`�E�dU��k�ȍ�ӹ�&�Ѷ^�߈&�h��T,�����ݫ���Yߖ�(4rZ;^���L#��Gpz�/��|_�J�ã�E���e��0����1��Na�(�.Gh��82�$�K4�f�i��4��<3�Fa>8�El�l>�	!$$�A;��̖Z�=m�,6v�V��yq���;9�����D�����T(�h�����|6K8P�/|w�5=�w���a�É2O	��GQ���P�NtH'��Oe�ť+���I%�MAQn�U�.�p�CCCG`mJ��ʑgtm��AC-&��D+ 5h�5Zl�1�54A��Py1�T��l"����׉H�a�h�1LuJ�ϰ�?�X����WˉXʊ�UT�C�w(����o�>��(~�E{g�v���0�8�qq�""Q%c(��|I�K0��O�4�N�x�ӣ0걐���*�~�I	!$�	��{�k�rri8d��$��7�č	��<�n�.�˞�(h�~�M<Ņ���!���X6��C�!@�>>9�J*R����H��������g���vA��M����L;9�ĽxH�J�qH�h�+����~e6F����94�uN��`Цo'���Ӊד�GG&ΟBx`nK��n8�m����@����	ҳ8��n�ۅ9�����'�EG�f��8J��8�PI8t�	8t�f�i��4��<3�Fa2\A�}��α���S�o1�����|p�d��&��DT�ZF1��b׾ �	 ��@�ڷ���j�K�*�_�taU��9&���f�ݣ{���;���1aT���@��[�uq�:�Է�p9�2��ɞg��G��v��ʚ's�5y��z�U��]:�1L@����	8�ϋ0��só��xqte�r��%��4��!5�ȞR���΢�c<��gI(���,��,�0�4A�����3�̔�~��Sck8�C2�QG��8���O�,R@1������_#������%���Gެ!4�>
��t�&�M��:૬2�����������]��T��?ap��8�4q���%<9K��t�
!��D��aAA��O�4���>0�M<i��xgN��:&��7��ď<��u'p�vWX����:]���I	!$�gX㟷
n��Gz��X�]�7�O&��� ����Ҫ�Ri&uw���{��ב�6�����+E���T�h��qp���T�{�66���-,8;E��Rh� �����nq�;��0��7L�'����E
Z_O߈I:��&fj���M�Fj!a�#���h�2�J>#�_��U"�*3!��f�Vs�ݙe�aᛎ��x�F����Ó�d�8t�<Q�'K4�O�4�Ox�4h#b��Z��R�"L�O����L ����� �7:C����r�ac+i����1u#I=0�Fi6Q�c8�����j��_��ê�3�fQ!�qa���0� �q���&�h�A$��������;ZZ[)l�hvt~?C��2�|i�V��8���D�ȅ���|x8g���>8F�Μ�A�#�?q�w�2(b"Z�~p%
�	�<<��s1���!��Stۨ��P�xX���wГ�q3�4CdӰb��b���IN�x����Y��a��x�ǌ00c�s�Pi�HIz$$FyH��5*��⥰���Ͻ�BHH�@�%b��R8ab&BA� �4a�&=��DN���SaK��1�I-�܈Yd�:��Ω��D!��Z�l,gF�$�DQ����,�a=^�H�E�3���c��P�Fa-�G��ӈ��B	��|�ֲ��X|z|y�ϰ��V�p��N���/��y6�t0gE�'U�/�^F"���[�NI�籸u[�G�xN����۟/B��:5#��
:B��3��pt}�A?"G���tz=:F��Q�1�= �za:Y=6[�������qm�3����f�v֌{j���{#�;�u� ��B�3�ѭ,��!h�z3��4��<?��4�����v=��4�F�#O���zG��Ύ4�4�4zQ=�a���Ѣ~�~8O��|Ǆ>C�	<84��ViA���:�ӄ94�4�4�4��Ӧ����|CH����4~�I:3O�<i?Y�Y�i�>G���"�~?G����&~)��~!?�� �Z?.A>U>�&|:�h֎FY�i��C����zt�6H�Hc����4�3G�m7��l7��=����,e�>��U>O�>��D�(�r���~�w���t�����V�"���(�d&�#V�	�	��-r綬��%�.u�����%E�N�U�5��H��x���EK��V5,쩅R���˪>�O)Nr��UŲr=��@������K����o+y����b�I�VU4�[� �.F��:��esבcR��'/V����2:d2㾒r/�M�YX�C��D�,��J�YT��m���g�;sD��=�Ͼ�ڦ+5SGW�vU�R=W�]�[��H-�S�٦[̤�ds��'�j�����$�f�k2�8�N�e�D�*(�1���r���ƙ)v%���������_�]_���z+��Xm����u��ݮ>�z����b��廈q*J$�Q��Ů���b�4�0Ӓ$�W_fq��d��#n��/mUz�_����fff�3︫j�Պ���o333��}�[U^�K��������f}��]��V�s{�f�:t��(�'K:Y��i��4��ó�:5,EU;�vGWwu�K�����-vfճL��,��B��@���%.�{O1ذ�È�+6M�6+CZ�9v%����XcMf��lۍ{;b�>���	=A!��hu�5,����p�UhJF묥n��G�V:m��a+l �������f��K���m������Z]��V]]5aTt.�,��lJnX&��\`�����+n�0�΄� 	m�"_K�����Dt�1��I*�K�����ir��Ҷn�J��2�h�V�F�[�2��K�P�*k1�jj@��]]��o8��b��6�t�]\Ԣc�X�k�is,&��6���,�	N{����,u�m5�u���h��1��X �fe��Ri5��G��BHI0�s��O_2�E5�	Ro�[��9�̂G3�\��؛�'j�k����<n�8���#�P�Z�WR)��Ɨs*���b���=��+��U�D�lZw�[�^�˿Q�M6�A�<7�W���\>:��4&q��7��Ӈf��0�~E��Naò�����0|-Co�T5� �������q�[*D<�/�����\|iI��(ca(�Ơ3r�c��Y�6���t�����cc�C �*x���r�͛�Yim��l����)�3�?���a�тyO�d����4I�H<Y�pp�H0��I0���>0�M<i��0c��6�?2n�����|�2-(�Մ��L �S!Ju���å�c�)]8G�X�g��5�q.d�j�Qã_����2!ů������D.Y���қk&N	��^�$p��#��;�AĘ�]�ppC��>L�C} ��Q
���8M-�#�N�Q��@�ޘd���F;&Ȕx�t�fÆ�U�#�R�/R)&3���gNHR,�$ �H(�GI><af�i��4��`�+���p��&hjw����L �^ȲFOp�����;4_#�8Y���Yt�(P�VrH	H����}I�5��] ��2��<�4�2���»"�#-Rg�і���݁�gg�4q�����ޜ�4x��,�1�/A�}����1��T2�������x�@�n��Q0B5a�:%��4I�8{!QpQp,��yٸ�'�Q
jģ�\_#�  $��(ҏ�:t��a��x�O`a�,︩�-���Kj���BHI	&JI�y�{��pRt��+�]GGX~��bJ�����K�T�K��:�t�W�"�1̶��U5X���uR4��2�Z;�DE�Vs���x���=�t.p�OQ��3ʓ��Q�C��ype��>��Bd@�L��p��|q	�⃈��qc8�/P�%W��ۣ�80�dP2�-�-F�Qkg�GzJCLEYGO�,��4�ƚp��`�E�t�x����
���ݶ��<{?m�]�,���8��hL���m�3d�jϣ�e�$�K�>�<f�])N�N�����i�᭥�qv���P+�p��N�n�&H�$���vN�x��>��x�)�E�{��y��o�_��!>bw\�Ӵ�k���p��X�f�F���ɳ���rn�JY.��g���gǐL�fo��>�xsp��ߕR��Ө����J�Ъ�vY��iAю{�H��}֔��'�e����)�n	O;�6�+��8��#}�k��&V��U+��QC3�|o���]*u�8*Q(�G��q@�������!�e)GQ��ʪ�y�3W2xYfVR<>�Z�
�:b8ǁTAx�@U�4M��.D tNS��Z���K\��N�0����4faG�>>,�O�4�Oi�0e�:󔈉�:���
E�O����L �����>�����	@߇�
�~�eӒ��M7&y���(?����J�tꤜu�;!+�tx��g�83)�7��LW��q��'�ќX_8g��z�j�~%J��p�#���˨��Wӫ��'wB} �T�,�o>ݚt<s�]t�V���咎{"�������t𓛳,̧���3����x��:��8�e#�ҕ���#0g�؈h��z�Zb�P�((�Ŗx�4�ƚx�fe���34��jT��~��I	!$�	������H�QH��B�:�I��:2>��\Pe�DA��(��ўL�:@2Q�$�{�U1U�Ѷ����|Z9G9��$�o�:8N��{*��6�LF,yuY�̀���]�ǆ�>^>E��պF6��\M3���8�Q%������@�3�.#�6�6�����&���u0|�C���f�Q���4��M4�0��YJ�t/�А�m�~�e�[e����Z6�֩pe����G��*���~9a��Rf��_#պi�c=ۯ{�njT�C�A��nI5�Ȍ�,�d������g�qX4PX����d�%Þ;M�&��T��#bv���9�oOA�Z4GK)Ã=]m�}=�z���o4�e��>�����R-�D{ȡpg�47��7	�v�:�_*�����.����t( �Δt��4��>0�M<i��00��S�F2
>������_D�6�T��H�3�|�g�����ޡhc\E�\Mr.b[\�z�Ļ��{}}6[BH$�"nh��we^^j�.�� �p��rXN^^Ĥ�y\��7Jb�vE�����i����c�H��+��Cl��;{UZz�gC�4)�$��:�^����Ƥ��ER�:����ܬa�A*������c&��S�m�T�M���y�Ƒ<�������C�8��/ �?$���P�#��à��?z��Κ�݌��yRa�xp'�����L<�såo���7��ɰ�b��b;��c>Dي��9�$��Q��c;D��Q^��:8w�~�����|�껺�lcw�G�I<����|�}���>4;7
��)OW�a�;�eL�T+D�:���x��t�Oa�i��4�3,�$�(����ِ�� ��]�ɂ��z�DA���TY�Y�߼PH�<���>1Z),f��(��ը��t�_�1�0������JGV�E��X�*-��0��4�w!p�!3���g���W�wa�#~��R��M���F��W�c��%�{_]-Xpcg$�	��������#��F`pd���."�ϖRh"���(�DQH�*G��(�L$���Q&�3��ǆ%���<X�$b"tD�DL�6P�!B �"Q^�6%���'��0L<`�&	�`�'�bl��a㥈""X��:�<�ؖ"lDO$0M�%	�6&��bY�"P��<"'�ckMm餚i��l�㧎�<t��pCblM�%�BQbYL�L �!��!�>>,���<p�ӇǏ�� �D؈���8'(AA<x<@�@ϯ��N}�5;��5ԑ��E��$��jr앆۬�}��5Om�xJ4�!᫼�x/o���ZE*u��ۼ(���o����F��t�ٗUv���/�]+�h�9�б��b��֬��h�o��A�ڬ�������e�lRcrv���dg^p�n�J�tkM�u���6CSEM�
�J�j�^=7k{zr��^+K��oo333��}�Wj�����������}���Ux�.�����ffgs�Uګ�iw�����C
0Å(��L0�4�ƚx��?�~] �	 ��@���z�IJ(��՚ut��A�A!NgiJ,�:p�٤�u0��G������D8���9�,;+�ܟ�GQJ�#��Hϣ|���Y��*��K�i�j�aj���4���g�8G�4vΌ:3�m���Y�YF(2�Ǻ��*s�]�y���0>Ç���+��"M'$�0��/�������xA�e,�4Q(��l�aq+ � $��Y�(���i��4�ӳ��;!��ޒ����2X��	�ȩ��}�HI	&I�����HXM['��ހ�ש9C�:<d��q�a��(���g$Q�c.�"�lK~�B�[u���g�)Gq�C�8j��/p�:r���,u���PJ��D(d�|{\̾�����&}���j���P�G�3l;QĴ���>�
��ϗ��t�s��-�����ICߝǇ3/�(R	��NiGN�0�L4�Oi�0fY�3�0��m��LQ��Q���}��>��h�f;�b��pZ�/A	j���	 �	/\�h|kp�,Ț��*�#
���5�ux��f߰PҮ�6U�n��j��MVIGuF�ś���L���t'�W	�b��Ҭ�L���D�{1ޕ�~tilp�9�M�7Q��;9����D�s�)��0�I�d8�j3ݝx&�oO/���,��kn�N�aE����O�M��L.k�]Ç�'�3��^"4��J��g
4�p�K��6�<���DB����+
�
+���O���xo뼗y,��Ŝ�i�X�]D���üm��E��P��*;�3���$���$��$�Ҍ<i��a��x�Oa�0������Y�ʈ�96�Y׸I	!$�f8S��q�dN��.f�6#�8�8��J:.-b�I^�㈍6�)E#�.�Å�$̸"e�#��"Lm��d"��V�$��,�
��<D��n�
A��<�w�n�7Ϣ>��E��g�ܦT������r�xA��xW��	!&��*x�,�����%"_H�:����/Bh������;��$>$��GǏY�i��>=;;;�	_#�&.GH���GS�HI	!$����##(0��0�@Y��*W�z'�ְm��(>DzG���8���K�m/��몉��9�*�ʖ��!�J%��3�Yl4(���g�a�ƪ����J�`y0֧���h(:��"��8V��߾���~�{&2���j%dIH}�{�VXϼ>$�Bh�~��>8���tc�)�E��2�,�'(ӧ�,��M4�0�a�Ǒ9z�eM`�.��6M����$$��DZ>��s�<R�`΃(lC����<R��B:��x�E��>�ƒ����%�UW��2��9�+������W!ţ��a�ը��H�m�3AG� z�h�K��:�#���o��PT֣��|��-b�zp<x� m�;~V��}^,�:P��HE�n#QA�<GMG-1�3�,���|i�a��x�G0��k��U�����)h��a߶�ۢj����R�B*�2�P�`�&͗m��ɫ�O>�A$A%���_&�l��v�h����^�c�XpvV�!�f��8����8�����i�c�Ļ�+-�oյ��1k���w�r�[}Bѕ vŹ�9��V��꫽���C�!�1OpH�'�A�m�II_�A#?���='�z�Go�����)i���kP$�(�(�^�P�{ �x����]۩E�Sf���%���ԞPû��q4��L
GV��J��CY�,�i|b$�&�n�'=�"������Y��D���3$��<<�b����/���x��(8jcr�x��15g����A��p��a�i��4��v'd:;��1F����5��<g!fNo�DDB �8^P��y}ebm��W �-�(�Q��mǩ�c@�~�!�Ff���w�ʙl����F!U{���A�|j��i��GʐҴI���C4J)b����zή�KTY�#���8>Xp�Ρ&��a�WYn��1pֱI�ߏ���T������7۞�(h�H�֞,G���we|i�tI�o�Q18�s�xⓁ�INp4���4�Oi�0fY�xEb��[E���$$��)�oJG H��X�ֳ��AC}j�N"�⎃$��	�����Q�5�x�p���8|i�a�2���O�m�X���j�C�:>�W�w��1�VB8q���1qa�Q�C��F2W�xp!���Rs�%"������bIdKrR0�ȅR1t����R�PZ��6#��*�3�p�GO0�4�Oi�0fY�&�ANf���C��1:fɵg��{m����I	!$�g�)���L����S��f�Qh��D��Z$iEdXp����֥�\���سd�w��EJ��3Q3����r�!e�|:Xa���i���o��(��,\
8����hҖ"τ�k���<��B]�]�6¿x���3I��|�($��!�h�a��t�~o�}3]�Z�<J/�.Xu�DD�'M$�&���E3����DD�<P� ���	�"'���,�A�DJ(��؉��x�&0�0L�xDHpDK<'�"A6""xL�6��,D؈�0�(N	�6&�<Y(D؈��'����:%	�"|i��,��B�(�I4�� �<�&�&B��"XlD�:	��,���t�N�hi�4��<x���s���,�AA>�Ais慠2��gw7����Wg!xij�P�U��唙F
n�
!��iSjY�n2��H���%=x7qd�>v�E]�X�f�鎢֚�r���{eX�A��"���Y��*V�+X�,�]U��Z�Tv�uu��R�f��#������
ͽ�Yt������̻\6����U�*�����r��|U�\�Q,��"c�>9,}烸⤍�cJ$ݑN�r�$c�ß[��I,[�E��l�k�ﾙEqPk��%��2V���Q��#�ֶ���OU���E�V�d��UJ��)$��,�$���\��]�\������S/����e�;�A��Mc&ֺ �ܶ��ް���Y�o����앤G��6�Esoi7m/վ�g��ܚ㶙֚R�v��4��-���ե{m�#l�lFc�t�M��B�>
o��}���v�n��7��ffgs�Ux��[w����333;�}j��]�۽���Y������U^*�V��o�ц��$�e:i��a��x�Oa�;!���	l>���ƭw]���k4Y�g��Z]�kp��t�r:�4�����\V[,���ōd93���v�k��Gg��������m1N��mS<Mh����I}|^v���8�lI��)#l7`�vF# k�Mq�-�j�-�S�Ʒ)MH\:�7K+/����r�����v�itv]�{M=�9��Zٹ�ش��"�.Q*#h9��af��5]vbSqGW����T��lYl
9їF��kd��������s��m�̟7��Ks0�6���&0Q�G^K7�tq1. 9	����Q��1+�[4:'lb�tT�c1�1����)���m���{zfVn��פ�G#REڒ.����$���`�fv36�AP:`���gٔ0U���Ы�F�PN�U��=i�L�ɓ`N��M�5y}�OkT�D�نq�T�Ķ�P�U~���7&V��Z6�egM����+��ޅ��RNFԻK�-`�UJ�-���xg���8%*D7���o���	>-m�1�}ҌA����EP��@����_&
)k	b��0����z����	X�u֑�,$�<��!3T���L"�8x�*}�Qʋe�72Dr��Ξ�N�AД�W�
��1h����!]�\T�6��N�xP� ��OQ���,�M4�0�0!b��kgƑi�� ��Y�3`�#�1i�8�D̬��߳IDB ���R5E*G�^����#ŏ���A�%��(����٠[K��/"���n�4�E�/��1Z7��PQ����N���
+��a&,Vr!R!i��p=��H�c��3�Jd*5X+���>���ю=(��Mk�#WO�}�F�X�L�J2��b�y(>-pd:���ʠ�d��$���<|a�f�4�ƚx��g�&-�(K��HI	&߸H����g�uj���5�����pj:�iY��b0�c)Z�>km<GC���6������|?#xњ�Q�t�I�u�;��M�!|���$�[v��A�6݃</�È�\��)_t8z��$9(�β!�7|̈�H����q�oa���1J<�)4��I�$��I:YG��a��t�Oi��0fZ��UQ0�\)��n"��	-��a$$��p���g��!�>���$�#��ozx>PO��?5��$H���4�Tf$!%1U'|�.x�aɐ��h��#����}zF�u�>&��q6v��p8bZj5�����#�3�����EMr�L�-y8��ɘ	��]�ۇ����3K�p��cc�R�g��Gk��3QH�t�Գ�m�|C�ז��8I��|x��Nt�Oi�������SQ��Wٹ/L�C�O,&kY�h����*	��xB�Jm��p1-]O�A$A%������ο����w��«Xp;,9F��uCt:�sw�+�}�ߊ4�o!�;3P쳎��8Ԫ��V؂�p��:�6Og2�p�{.��U]T�K�jZte�8~�w�`W�(ኔ���6YH����G����eKm��p���3��[�(���� {���cV1�]�p����G�$ �}�$��cg��]$R����J:E&[L7�j�^�����F����\Qwc>�������Nx4��cm�ն�]� �p �4���,����G�Kx`�p�&�Y㦘|i�4�0�0!~�K�e "A�7)�I�DcnJ�h�ue�)!������\B����
K�'Vt��WCI�}��Tbbn��v�ACv$J"��|�(:��x��K1����	|:yp�i197���/N"	^'=�j�0���UZ�wz�W��/!qF	��:tk|6���\2�g�=��^���y�~8��u��|�I��Ψ��J�N��G��$�K<|x��N�i��4�L���>���n��D]�*y��!u�������BHI0�O���L8u}ã\�v��\^K��.�����N�D��q�1��1���E#�n��y��8y���	�(#M��Ӵ�U\���v���������%�� �-x�Q���B����F�u-��lvHt�Vw��J Fݢ?4�E�;t�+� Ѹ�A{@���:�2�<Y'�,��L>4醚x�Ot��Ag��LS� Ye���}琒BI��.=	�( �[]%D��=4�_��*����a)QU�S���7{��ݖ���r���?g�UD���3���n�T���\�,8�2LӤ�Q�y|B)b�+T�%g�PU�MR8�����ڐ�Q��鎑F,��$Ίf�y����<�i�
8W<ã��#<��i
#��s����j�d"B	�Y'I4���t�M<i��:`����C�F4�T�\�!*?Q�)�gEVDJ�W`� b���G�Y�
R���	b��v������!$$��?��~Kk)���Ѯ����>�ж�QΗf��1V:�Kƻh�Պgu0��IR�P������#Ӫ�M8�����@�g�R�}u	���0�-��9�ư���26�ΣJVèR���ĔꔩSþ����q7�����p���I3�ţ�p��՘-	�u�p�p�����X3 ��	$a��p�>���*A��������E������p:tŧ�l�>"���"*i��������Z{$�2�2W�+'�5R�e� �0��Ő�)WH$�-b<`���H�Q��$醟|i��4�0�0����3	&���D$�C�
Q<�.|i���>!��҃|��\Uw�6CŖb��*NaVj A�,�J�>p��� 9���5D�8�i��k:�yh�އ���2�K{��g3U��y�����<$�Ohy��Dy�u��n=GT��+��Km��$��Q��p*ۆw%B��
1�K:x��K4�F�Q��D؈��'�D�"lD�<P�""x���,� � � ��Q��ı�'D�&&`�&	�`�&	�$0<'�"CM���<&�!BX��<"`�'A:tN	�6Y�� ��b'DLg�D�"lN��e�'�:p��hpӆ�I��A�Q�ɤ����D��lJ����N�0O �����>>0�舘t��8YB!��x<ьek�7��|�����e�+���`��W]����9l���XC[F-#j%�&&Y�vI��W�X�ۘˮ�\�@�(�ڭ���De��Y9��l�J�Ư�wx�L��K3wV�t8H�:�)�%gY�}����z��,j�~�'.��ٜ�5Z3.�{	��R�᤽�����n�����s/�疕W��U�{���������R��V�m��}����}�*��mU�����������R��V�����u�ӣ:t���(�M0�N�a��4�N��-�~�ǯ�DAD�y���F��¿a�?r>===bҕ��&�.���H<Z��Z�J�1=�q��������v���K[(X["�I��p��vp_�G�Ӎ��i��=�y_/χ�|��d�g���7����Ki�#c'��N	{�rg���r��H��8�h����C���ؑ�3�loC�8jQ�R/�M���Q��Y�K$�F�x�Ɲ4�Oi���[}��� 8���R�Y���1ݪ�͸�MvO}�BHI0�O�_L7y�b�:|�A�}���N~�~НPiR�W��%Q�I�dP��<�(G����i6!�����1��|���i@�$c����ѿ���?f�Y���h�9��X�=n��˲t�e���P'�	Bh�_v�I��b<�sԖ���e�PHI��8I��(����t�<i��:tfm��s�""!�&F6J�D�r��v��Q&I�q��u^c7َ��υ��/�E�]��m�����X��P-y͸�X�I�Ix��k�����A��)��M���tD�>��]إj����(���������'&��(�v�A�A���h��Z^��-Vh�is��SN�8��$+A�2����or�T���tnd����E����t�l�4#��g���GϓGY�K�}�+��ыC3�U�\��:��I���xg����Dc���)�5q��=��ȥ��y�G`�p)1�c=" � Ll��>'��=v��k�|�cc���%��+h����G0맑�s���^��#�6ƍ�2Q�'�,�M$�G�<a�M,�ƚxçB0+'(���	xԡ��K~�h�mӪ.�}DDB8�)>d�o��x�����;ͼ(��,9MmQOG�<G����M��O�(�&ŤqG���P��z��5Z��I��1B�W:�H]>X�à�"w$b�=���Fr˴����zuVu�!���Dds�v�^֏�F�9#�G��n�j>��|Xx!���ن���l�7��O���I�Q#>(�Ğ(ӧO�4Ӧ�i�M<aӣ0�mӖ�!�H̢j�@��v��I��m�ũ�g����q���+@u�׌\F#ӿ'1�}��P������<I'�P/Xy�W�-���u�Qz��d��w	�s��:?g�~���k�2�ۖ������1�N�3���h��8����Tj]01}�$F{~:����C��C�{����t��<Q���t�L<i��:t#B�o�pV����ۍ�V��	 �D�G"	c���#����"
\���ִ�%��E̊���S����E�<.��ޝ�)��`E�c>:#m��<�E����)�$v��J|zg��i08{������Q��3�kkaǦ�K�-2)�k��J�X{{��qu�Hyt��c��'U1<��A�$�Nx�:x��N�i��4�N���[�&�q��c��]�V�P�� q�~o��4z��fV�S�#LT�)�[�t'�_xS4�)��$�P��b�X6*����I����%	���b*<�O.�9�f���[1�sT��f��u��Zk�)��ꆰ�ֵ���^����đJ��[lCyE�]0&�Ъ{A{x��jQR�bEJ_N�����`1d�LT�ㄜO�Z�5���J��z~�8���|���h������p�K��R�e6��g	�p�5h�%G�8�\���F�<��l�.��]ESTt"Ǩ�(1_�� �s���am�|�)k'r	-$k]�d��f���d��!r�D��к�텘2�a&aӧ�t�L<i��:tgH�ܿ=��dm���I	!$ì.L�b̠�qCci��C>�Q�8.n��ߨe�I5PU��Z>F+4������V�s<�!�N���%H���:h�b�\͙�I�����NOA��9s+�-���;�Iۑ")��h����\O��G;��:���3�8R�E�D�K�_�ÑɄR��2�$�M(�O|i�M0�0�ѝ"�㱎�k��9Å�uy0��y6���=��I	!$��w�HG�"�a���Ss|���J ��`b!E�B=4�4yo�0'���;2M�q:�>7���[%�ۤ:�R1-��^'�z�>]V�:���@ڳ�t>9��G'p����o_�V?�>�.��-��D�uI��h�g��u[�.#��D4���<I�L(�����:i�>>=;<<�t9}�ӭ$m������I�Ixk$��Ht��~��(}��^r�C���G��`s/��� �G�#�]%��Mb?��2dr'�)<��4�t�t������8�5�;e��V�^��b%
F��~S���&goę�1�(fDll�q-E.���A��c����$؏D��q;�x��t�Q�����ᄞGW��O��Z:)�d��|o����Æ�6A��0N� �D؈��0��D��,� � �`�d,�bX���tO&`�xD�0L�`����<'��"t�b"""x��D�ıb"xDD�:$6tN2tM�p�""X��� �D؈�0N�	����(�Ɣi&�i�֭mht��"Y�(K�Cǎ:tD�<P�$b"'����������>8YG�� �'��xk�%�5c(��7h����N��y�=�+�[v\)e��U��k#�Xá/��%����ǒ�W�x����]!�m���ct����ц2"��QУ�Q�q=��X��%�W(@j�)�(~�d��0%O����3�{��i�7��U6�+�S�b�Q[Ɲ*4�8��Cz�ү�vM�}�����) �0��{Y[EP����=A6��r����~:���MJTZ��._���ao]�YzQ|U,��>�C�i�a�ɴ0�*�a	�^B���_Nj�v8�eκ�Ꮃ��T����t/.C�������߰ϫ~qb_n���ߴ<�����VVP��ś��I��P8�,���Zt/\hCJ�;;].�-1lLv���n/$�������{ig��Ǵ��H6P�ˠƛm+WlL��d��K���i��,��BQ�%��@�a�����U�����ǻ���ګ��{�陙���}U궪�{�ߌ���ϳ誫�W{���ffff}�EU_-*�����0�afaGN�4�M:i�4��:3��~e�OB�����q��iPی0AҸeڭm���0�@Z�N�J�#2�m��ʖ�0X\:��!�I�D�u��&j���SF�K�,Д�bʶTv��m��I�gKqvCS�2[����s��-WGez�:��q�Yua̌i\��L�ְ��ưm�)b:��u��,��١SU���f�]:Ԛ���B-���#]�7`��)5�&�R�R��kY�:�*��0c`�l�l�!֓J:�:l��m�qA��L�e�#�;Y	q��#iMf�w&�/-��U#)Y@ՌiT�I��Eu��-uh��� �$v��fѪƣF��k4�M-���r���������3m�����s��̤��dm��%&�!W6\��[!�lZH�ڐI�Ix~��}��#��������{bu]i��
�(����q�C+���&��.��iSʄ��{��V6�uF�w��C\ê����x�Vh�u�����k]]6Xu�� 5`�y�ۣ�͞ݪK�k�K��W~��~�~�����x</���j�"f��
dD(�֓��TDCnQ-�5|tr�,-O"r�\<c������^��m�o�F������R˶i]���zު=Ihw�Рd}��*IvI�I�a5n�p������ξ�߆բ�F���I��Q��<a��4��i����.�Ü��R���E�����.�U��A#h�p�Xp]���ʹ�B��o�E�߾?!�<��LY\Qq�	�B<s�7k���ģ F((����>G��$�8b_���&xo0~�~L+�I,c!B�p�;'��b�{�_V#Z�����hb=e}�%��t�|�)�#Ǽo��wXf��$NC�Y��0�0�Ӧ�Y�M<aӣ:Y%瑬!�p*���"�.�o��l���}�7�_#�F��`՚�R��[��Oup��2M���D��}4t)B�{4��ſ{�PoG�LF�Q1D�o4���&qۺ��]����<Z��������� ��6��^<� \�t>Q+�O�qZ8�5�G,o���q��C�i�6��^7��%x�`IC4�'I0���K<i�M4����ӳ��<:(�H��`��ccch�4}�Y�agÇ�h�@�!?e�	�a�8�D������8���6�a�B����88�-/���Zb�Y5#E���'����nv��d�b�3���E&�UUa�!�<Jc�ؚ9w8D�[ѯkz0x�"��݊u��Ch�(��Y'I,��M,�4Ӈ�4�N��d�o;2L\��eG�T$PU*��J�3T�6�Si��~o�'�~��L�m��5sZk��їw�(�u����g����~��,�Gn���_�$��N�q�*��9�n�`��U�����8���A��ë6T#UUȴU�&�(��\nE}F�<��H��J}:吹�I?}>Z0Z��w��?[�cfY�t"$S�I����<�.��F�Q�{�>���6�+�n\(�8��<Y�e�[�{��ӇBC/!���B:H|q}�,��QK�(�$cl���G!�N0��B�Z��.�Z����_�����4ݐݲI$�+W�Q#V��>�|�R��8�T?�K�Qad�Ĝ$ҏ4��Ɲ4Ӈ��ǧg��xtQ�U�����D��9��<�Qp�u�s�Sw����t����qH��&2P�Vj#��J�I��@w���axB�^����: ���W7=��e�l�\p���D��,ս�px\�|����)��y5 �q�b�52Q��,�^AH8�n�{�
�#�A���A̍��gUi����Pj4��R�|zf��#�D���K$��ƚY�M:i�i����<�:�H"b�K�P*f.��>�(��C��2I�vϯL<x�4z�i�Ő���`L4�|9Pt�����Ԝ(��u���� ����izBR�*EƓ#��z:Q(���C�#�o��ea�Ŋ�u�Bhd�*QAt���A����F�.J����O�_a���Z^���ǍK��#˨���FI�OaGN�,�4�Śi����*�C�Lge+爢���������M�?vL#�V�V߂��H�G�W�?b�N2��BA�8t$�L�u4u�����`L8���}��2�m�!}M�!�Q�Y�.[����C������#�w���s.Sﴂ�s;���\���u^$�+1]���ӡk�o�V�.�gE��#0�%�x�㦖i��4��4�N��d�M��ˉ�G\�r�H'f�H�T�VlT�h\ �*R��,8*�L�A��$Cuꔋ����k��$	����JC/�X�=�����[3y����Tq�"���0���ggt���RYS/���oF���Z�ݭ�B��8���P�1������FUX�ӁR�*h���ypT9��E�4����m1�$�i�-�pl�F�K���G�>Rp)GF��j= �êE�팰�'�?̢�K"�~ZE$7�7��[ߴá�1�^���:p���}�����Ӻ�h�h�F�?�qA�w�ក?X��u��3"0%��aݕ۽o�>"<ó��s<�[�~2)GQ
��yp�Yc$�Ot��O�4�N�i㆚xçFt�K�9�h�{�(���N���p�;2;{��Zh�usb"DDGf�B<xэ�Q+��Ԝ�uI��>J�x��	����0����[9�a�g}���YUݔ�~�U�0�*���<�qB��?L��e�|��U�>N��~�a�E�l��yq|��hk�5'�ĘZ�C�K8p�8pæ�,���A�"&	҄�D����0O�p��X� ��b["lK8"tN�xO`�&	�`�&	�"& �<t�e�0DDD�B	�QBl؈�=�"'������:l����$DDD�JD�"lDN��'D釄��l�CĞ ��4�mj�և� i�
,؉E��<x��L�"%���&�||a��NA������x<xf�i�-I>����G	}Tg�,��1��;$F,�lIZ�R��Ōmy<��ge��W�4�{�A#.�۪.��5|���
�S�����]�l5&T��{1-�-,kM9�����w�Wn��ƍm��	�#�"R��wt��ײ�(����]�ڷ*$)��/Cr�нA��$�&��(�[+�Ўf�׸ �)�ٷ�-�̱FaZL+��Hm���$��T����e�ww����ҫ��{~3333>�U|���{�ߵ�����Ȫ��W{���ffff}�*���W{���C,��(��K4�N�i㆚xçFt�O{X��O�E\/�'�%�e��1p�gC�D`�4�J��D�}m���s˻F����m�Я{�Z|8�TR#�E�����,G�"K��m��B�G݅�'<��ުGʑ(������e/�q��T�\��h�F���Ӑ�f�0��C0�%�x�OY��t�OY��:tgL$�8��Fϟ������s��~:����a�f��P��8猢S�q �ŷ/ӡF��.� c����LF���8������i��W�4�����.�)jXj:`|��w�rC�p<4�yR8��QC�t�PZ�H�^e�6�Z*X�$�eLHah�u+:��B�H����p�Ox���,�M:i��,���h���l?IX�ԁ�q�-��"C�(*��B�@�u=Jn:��y߰�Ïah��E��`��Ժ�ec����=�UPMΦS��WJz��Gu��x7g�U��+��*Y�Z]/ [�e�w�q��嗩��0q��★<o��QЪ��2�b�DÛ�"x^�Yo�h+�ު�|w�ʊ�5D2�)�}�;�=^/��~�
����J�Z�6��D�BE)�޸y���Zj�	K<@�.���r�IF�R��Ӂ1q]�����i��]�����ہ`|]7���lx�0.�Oa�`�i�
�l���HI�1)	���j��upT5~7�./��(2�����F`a:Y'�,���Y��t�OY��<<ò���5����ӟ:�=o7�`͝M���6NOx����t��<=�s���;�+�nUӺ�{N���-��S!��w�5k7n*I���ʑh�x��Ӷӏ6��Wp���OOB�̩�����]���gٝ�s?�(\��?]�Bn��G&@��[m���f#�h_F�tl��='��3��(�$ߊ���0��l$YԟHj|Fa�|3c�8�6�t�O�4�M4��Ɲ4�Ɯ4��ad�9�����8�B�䉣�x��x���~�<��l1�C���,��ʑ�p���û؈n(���_<D��;5
&%�Y��%RR����T�~B�C�'�y{<A�|t��7��`�����p�+������Q��:8e���^L��&���j�I��Q��{��0W��vJ�����p-}!Ã,�NiF�Y��:i��8i���7_8�����}r�$&.[B1k�$�Gx 0^=�㭳��t�ʖ�J�+��&b�- V�滑х1N�~���D�A���4�)H7	Yg�)�G��j �#/jC�z��,"F���SO���>�O��xw��$��y��F�4��t��q��������A	a��CM��(=�0>���è����(�	>(�ǋ4�M4�<t��Y%z��z�H�K��j�7��)h����BH����4�^D�#3ԓJ�ݒm���"L��YY�n�$�c�����t���o�]��fE1�c)�%]%Ӹ��i�^�8ʣW���ebo����f_ruuu�C1�h���Ҹ����+��Kk{��8�kgsf��q���MR4�R�,��;@���
KX`H��n�-w�q������رC�|�d+���j�2S
Wxf����༈�\�)��ȔB�����h�y�<|���)�:C-[GTpk�Y�P�� 1�>q1�D&I�C��*��e:�����g�Q#��Z���ώa�w�z9�x��
��,��t�gǌ<i��)���؝�5-�e��h�i���:&��3��3A�h���xhᾂ?zI�$N6�n5LF����?���ѥ��������><+\%Y��,��#_t�yKX��Q!	��Q"�
����n�[�p�sUL!�&։�$��y G��ga�z�G���ϋ4�Q
:�l� ��.s����E��P0оR	:�� ��~U�(~��C�D�$:|Y��<x�ƐtӦ��73�=W0��K�WJI2��]�)P$�*}ꪤ���m����D��-G����4ZA��q4p�鄦����>�p����A��l\�^�D�-�����ڲbmR�|$�s��"#�a�},��G��x8b(��A&����z}��"�z=7�އf����7�R��o6�&{���T0�9����I��]��R|H�8I�'�,��x��t��Y#�3;3^�C�D�v�����~���>����D�i�<�����8�uҥ�IW�6�1�{��=�B�������PㄇI3Z��⃄�XJ9�2ϗ���DDA��/��B>��u}D-%2����j���4�(��t�NM�zg�s�$�:��|������(b�+䨪��aP?K����������fˣE�0�@�yR7M�����c~6�UL$P�� �G(&�&�#�L	�$�b �&�&"	���&	�b"&�&"&�&	�`I���	�`	�`�&	�&�`��9!L`$�`� ��$���� �H$�"H��	�����H��"ab	"d����&"$��"H�Y�� ��	������ ���Y""a�"&"&"H�$��""b"H�0 �
	��4`��3C$DDID��D�0IDDD��D�D�A�B�DAD1$D,D�$A�B��DD�1I��DID�DD�0�A,DLDLK��"$���"� �!`�""H���"%�!e��b"X�""%���"%��b �"$��$�"H�$�bH�%���"%��b"X�""X�"%���""HY"""H�� �""XX�b�"%��b"XYb" �"�%��`5��A,DD�D��DD�AD�DD�D�I���A1LDL,DD�KI�D�D�D��L�1�K�ID��DID�@@D�ADD�d��L��DB�D�DD��$,$ADIA$,I�L,�0DLD LDLA�I11I�,�A11LD�1LDL��LDA0б�IL�	$2C$!$2BA$2A$D$2C$D@A1$C$!0B@kX	�R@���� `	�1XH�� eD��5�jЄ)��!��2$!(@�0���m�M�D���&�``H�� `HT�� dI�1R�� eF `XBU�� LT�� `��`eH��``H���BP eX@��@��`aP `B�`dE��`dB�� eF��� aXF@��`eHXF@�dXR��``XQ�� a����� d��``FT��`Y ��`% $ !@��H	@  B�	��`!BA !RA %R`$C#"�b %F@`! !F !	�a�dBRR� !�a�!I ���A�V!�ea�!HBXda!�!�!��%Hda�!���T�VBXaReea�!�� ��V�!�!�!�!�!��FXadHRV``a���@�HeaHH`1#!�!��XbaH�!�!��Hb�H 2�e�!��!��a�RXb�a�Hbb�e�!��H`�H`�HR!��Xb!�e�d�"b!�a!�b!��!��Xba�e�"a�e�d�d�d� �Xba�a!�e�!��!�bHba�b�a�e�!��X`�H� ��H`�Xba�e�%�d�e�d�!�b�b�!�`�H"�	�$�%� �"	  &`�`H�`�& ��`�&�	 �	 �	 �&�`I $� �	� &�	� �	� � �HH �H"	 �$2Ă$� & ��`H ��`�	 "	�a���	��H��"	� &�:�`�&�`�	� H� � �� �  ��`�&� �H�`�	� �"`I ��`�H	 H &�`�H �H�b	��&�`"�"	��&��$�f�� ���H�	�`H d�d��HH $��	  $��H $��H��1 f �H`d��HH	 �"	 X 	 �	�$��H Y &H �H`f���`��f	�& �`.0$�303A0 L0A�D0�L!0L4D@B�Lq�"`�Ba��&��&����&
�a	�`����;���a�o��]��S��=O�w���UQY�"��|��j^�������w��|����׃P���>�ϯ����ߥ���־����_�0�=��ێ��owΜ�����kb��;={M������?��vSt���o[?�v{ @�_o��� ���8�'�QG����(�����@���vߕ������#�Zɂ�����o��������|��F����Q@�Q?����~�T/	�����O����o
�ƙ>����I����ٴ��?s����O�����7�m���ѽ�"):�����u��* {4hDCB��t���H@�J(v0��"	����6��ϵCn}��&k}G�����'�w	��L�4B�0"�P  �@D
������A�|�=����ǵ����y������zC������"G��/����|��* b|\�������?�z@����z'��~��b��tl����G���~,p�+�~�6�I?���� >�v{_��{���9?���� ~π�@ݮ�u���g���I�����q��Xh�߀*����Q@����++�?���ր�6���~C^��;�~��u�)�~Q��
;��|�ǃ�4���&��P `�~�t��\#�r�=�����?�1����e��l>�u:�cI��}Bu'B~��T ������}�����y�U �8���� o��۸�o��a~S�ݟ������;<O���K�N�	��/�~�友��o��v7��HS�0������������UE =Ƿd��l�,��~���Q@���|�����:��W�=��=�}�m���_�(�1��f�7�w7؃qv�?S����$�O���=���d=޷G��q�]�nï]�CuTP����p�8#d�q>)�=����: ��3��z��<:zO뤟���`��4���#�N=���H�
?��~}�4q�X�0S�?G�|χJ (��ޛ&z������O<ܘ�)�y�����}$|��!���;�'?��?�.�p� $��
