BZh91AY&SY����8߀`q���"� ����b?~�     ��2�iH 
֨�6��V���2
QQ*�F h��Ѧ��m�d�lց[Q��fQF�[M��V	D�VϨ;���yzə��ڤd(�m�U�+@d���-�-��E�M�Z[j�X�M4f5��[m��٥[4�U�ڥXm���R@QKd�"������T{6*իfڨ��0��6ԩJ�l �%��ƭ��)QE	li��j1�U�**����[i-m0U2�R�1��-��V�Q�:vHJk*L� �f���E�����wҁ�h���;TpZ�2�UU�e݆�lcN�̶u���UNCQK�[g]SER���{4�ť	�ݥ����  ׆�@:��t[p��)� ���wI���T�q�j���:��  R������t���
޵����z����i&�jYdh��  w3� :����=g=q�J�0��=�P�oy�=PN���� 8���v���x��)ucg���E�W��J��y�V��DkkYLƖ̒   ��� � ��|�OB�x^{ǭ�;�k�}>W���U�=�A@{����$W�{�
PU�;� )Bp�� {c�_q�R�CN��5�H����1��I   㧉R�����WC��@9Y�U nn蠪P�q.�
��4\S֊ʷA��J�ݱ�B��N ��y�!K�6�E��R�&�T� ���tH��p
�m���)M�ڪ
 WwK�(P�ޝ�u��f 
G:��  �9�����N�M�*�[a�H͔�
���W� w � 5�F��׮��=���P��UpSPSZ<n ���pu��J �f�� ��  \I*�T�V�)DV� k�
�8�t�9v�� nK ��ۡ�
��� 7pۀ 3v\ (;sn���w@S���IE��R�E�Z�MI�� ;�� m�p ��: Gà� v��@:pp*����t4Ӹ �40 4�ٳd�aU!���Q�F�  ��Ǽh p�  n���W:� (;� ̦@81���( 	��t+��   �   �*R��	�&��1JJ�  �    '����j� 0   &�0�O��%J�р�  F����h"�z&542Mh�1��$�5L4�ɦ��h�@h�&O??G��/>���i��J��̅�4�Z횯aE�]�Ď�.�f�M�
���ꪪ�﾿�Z ���DT�_� U����	���������_�|�� U��5U^��`W���$��)��������3(~���?��?S"~L��L��0�dN��8�<d2�`N1�xʼ`^2�f�
�a2L��8�W�+�U�xe8�<eN0�*q�xʜ`0�S��^2���T��<d0�'fW�#��*q�xʜa_,��&A��xʜeN0�S���S�+�D�(tȜaN2'S���T����aN2��	݁8Ȝa0�C�q�8ȜdN2��	�8ȜdN0�0d2'�� �+��3 q�8�d0�0�����(q�<���	��
q�8�xa8ʜaN2��(q�x�<a2����a2P�aC�	�T�@�*�xʼ`C��v8¼`^0�P�(xa8�L��D��ʢq�T�*	�E�D2�Q2 �`x� �A���@�"��8 �  �#�A��'@N0�a8�"q��	� 8�(L�'TN0��d8�
q��")�S���^0�=�U�"���Ȁ�e|0"=�2�<exȨ��"v ���U0<`P0C�	��(q�8�we8�<aN0'C�	�8��a2�C�v����"q�8�����q�8��S���� q�8��ex�d2C�vN0��x |���/��_����}�q����3�7��a�@�4�B��S�i��wK��N��ͬTGw�"�0Q{CZ�d��n=A(�4+��L�>W�!t�:*��V�oSY��;�8��l�opb�|UjV5�b��R�x��6�����[�)&�=�]2i�4k�-u�{�\8����S�j����ol%|�!Rśņ��%�$�j��*[��`�3NVg�t�1�+ �P��{�^
Յ,����4S��e�t�̒�".�Pشː�V@�X5#R�;�-1P�r�^�IR��-#��6�7BD[�IdZt�/#��
V���i;�YV��P1V9�dB�	Eq��LZ�C��V)����.�TH��5R�F��y�*f�:�BP˫��;�����L���"pbXu^њ!Y����/�k6��a4�x��C��8J�fF�㊝9�ɷblj�r�c4ˤ('��S�$8�4]�K$������i=��w&M!Z�:�.{0�3`�~�Ƶk��[ۀF�YKsd�"۴),y�I�u����m
�h; �N,f��2kA�m�`��x.V�0�w-��D�tζ&K7�I�8�H�Ȭ�z�;E�)6#oG���V�&�4�C�v�쬙%!h�!cݻ�)��n��9�F%���ڊd����S�:HԶ'�AP�W��Y`x�˳(�=��ӂ���I*-�Zj�8@,cS��*�o6���0�&7En b_�\ʼ�Ƞ�f��OJaYr9�
3�ZX��(X��CD����Ap^�μ�{�m򍱃v�W�ZN��n���P���!��P֔�NGD��,�bYz��	�g ^�0:x�#n�"�:�Mկ����¬��󷹚f�x<!�J�K@R�fә!��
s��KG7�[w*�G;cp%�(���b֩nT4�b׋K�G�[���~����0:T�dU�OL��a0�g5�HB4�pm�HMU�١1���:B�qKa�M��(��Xjf30�U�h&c�T�p�8�Ec����w���טe�Ĥ�)6��܍5S�ɓI�g���À��Z�5NL�����x��X5R��r�+�����K���Ul/P��d�c0n,L��N���]Œ�	K8V�.����;ắB��3��$�WZt��W�%�J\U��"�V�t��D�z���3nbr�.�̆ڙ��OJ�X�	�2q�nC��,�y�Oh�i���FV��C]X�c�!rnY��ٮFa��.� ��P�{slʖ�J�y.�����ɴ�����y�[�Z�mfҤ�9n���D�l,�2���Q��n�*�^j���R֨���}�Hz��i�w��;�m��,4�*a@t���;=�RB��c�Vy5ɮ,�ƻQ�h�3Qj{|���)�ܴo|�;aGH�xM�����mY�+I�6\��-"5�2e,�J�2׮��,û��K��b&�CɆOƨ�{�d�9N�p��i"�̓	'8O���y�4�ۤ��]Z%��ؚ��SE�<�s5�#4�M�W�#ĪV��}��#U٣2'#�҂�n����˘bl��� �^*��*��%M�̰�Q���L*G��w�ZRN����W�w6� �*�6b�X�T�2n�]�w7^T�E�y%��GS+B݇0D*���n�pa�,������dw�L�S��j�a�BQSt�J���*��A��E�x�!3 �&pk�lRڹs]:��Y�.�C{��U6���[�Y��Y�6���ڹ���K��e�Z4
�
��!@E&Ӣ��IHD���1�b�A%	�h�M5	�B�YY��-��:�tk��а�d&�2��5(��r���c�V�N!�g7r�͚��+X��cܦ�cԫ9�C1�^� ���F����YV6[Z[�L�y��7�l%�n���yl�
8�H�;Z2��U��e�R� �ԧ�vNe�=���`Я�7��c�C�fb�dgoZ�z픵;5���i�sC�"kl#z���)A,�ɴ�wj8���t�A�ڛp"��/-��Z�+j�X���Ub^��o��ɢ��ږ2��mIze9�Kp��b�5����{�1Ćݲ���?3��t�(ا��z�+,�֊*����p�L7lvmnL�(ͭn��)r��v�#"��5A�D��c��m��`@kk!�_��n"-�nJ�S���m�(��h(��SV�(Ħ0���m'���:�Xܣ�1��L��dl�Vu;Y��Ķ�3-���VԔtcM�45�t4=�H��ӯ3r�ǲ�P�:6��ʇ$L#�k6��@lɶ�-�P�m2�p����1�[���0�K�n���0�`����%MlfnU�mBKOc@	C#�H�ut��J���ZZ���A&S�Ks2n��r�تh�n%�GS�ź�C�q��!l���	c��d�/ ܂n�v�E��Z�����G���B�ˁR��/V7F*;K3(
¢�+t'�"�t��&k�*e/FV��ыj��T�9<c������[��Ԯа��,l9z!�(:Y��an��!��2Z:�B
�da�EV3��Y` o)�P�e~ƕ����1KFQ�m��M*���Yt��,hUu|V�ń�F%3L��p�V
٨V��<H��C(b��Y�eqV1��v��Diu��u+SW���(VZ8¬�U�7� 5�����ǥ�4Vf�i��v���K c3,��&h�g��ݟ�{�0]K0P�vƱ���6��f��9���%�����7�ؓ6���.�d��V�iehW�˥q�\u���s��k[['͘&��Q.�v\-!��!�o!�B����ۭ8��Zk.3)1���Y@3��q l��MG��(b/ յ,knX,喜(��"Z�1�`�ge��IJ�ȱ�N��e�6LT�o�*Yo{��n��T���x�/��4h��0J[7Me�U� ۻ�&�͆��V��q9/v�͌�%LѺ�@+ ��ڕ�Sp8�^;��+v�x��rA�O ����}wO.�(Ҋ����j�+a�3L�E����Zb�[V&Pe�LG���Z~����4��i���4��ae��Ma�淬�ۼ.�b`�Д1 qa����A���Ӊ�Y�ě���ɶ�]V�%�-�E��Q�q��%xb������7�ebW��%>�N��ZG>mpKL��ڌ��T�,�8^�0�+�d�&���cA-��D�jګ�!ʎ��4𼷙(��IF1���
�6<��X�N�VX��`cA;��ˠNmD(���픶-pr�u`�Si�z�2�6���Tʍ8�Y�6�ѓKɉk�Z��k[\�ùk�?+e���j�]2�&�7cpg��J6���v7 ��i�5&�h���,[4R� ��P�͋�/>ѻ܁�LP���Ke�N঄:�'jI�-�Ƶ��a:�p�8pmec���fmXZ3��N<�0j#<m�&oKOT�b0�.CB�J�*�i�M�8��HAY�#��bޥ����b���ܷ��� �j���ej��IX&�
Ŷ���9�~W�����m��3E=ĝ!�^�i�^!���1��*aˤiV��ԥ_��9!ǵ����`:�ZP��j٩�*�6����ܩ�K<�xS��e7D-�ȃ���q�o^�kR�6͂k�'t��4��LE�x22�[5"A
{nך��gH��]��/m�(��@J�ѥ �EP����۲��ɚ�R�;��9%9�����t�3�s,��B�x�&PO\�TL�W�4��tr�bMswF��V�/-��C�uّ֭abAj˴Zx�Ňp�W������'O��`�%�z����u�!R옆�z�0yK�-��YY���^ID���K�XS۵n�i)���"�fh���V��ͨԢ^�/e�f
��Uz$lòш�ˢ��	\�np��P��hu5���̧H`�0Pܓ6�@؃��*-U�U[+l���C��H]+����rVVk<Mm�ǘ3e-��ԁ�L�[i�UW��g�%�%�2�J*0�V$']�&�b��J�S@i����Q:��VVE�A2O]�H��hʖ�b�6r*#1Q�3Vj�j��iMh�%�]k���!��z.
q��,�=���op�m�vƆ�N�
�.��E�1�7Ng@ծ�fܡcڰl&*-��ڄ��M�ݜ��
cX;2$@��&J���mZ��Z���z�ZTHK��dʎ���²�f���F�5e�P�i��H��f��-�o(�0� -|�-pyě�6l������ل�X�E��������Q�1��m_,|�T����(�1�G��W��)�yM���=/����t��%�!�	��.`��s����2Q��˭��f~t�5Z��Šv��I�C�XЮ�+�˦�<�3Ø�5nY7�����	rY1��	��;x0nie���\�wmJ� �;�PH��U���8e�(nDJh�ڢ�Aa�0oeil�Vs@�d���ݣz�`�����iǴ
i�[L��ZkVSA%,���`���,Y�*�l��#y&�Se��I���3):r�h66�tnT���	2�;r\�/3"¤����QژҰ�G*-,�ֳ4�X�� �f�)��[Q�(�� ��^F�BFJ�2�(����"����KTii#Aw+2٠l
z���[è4Z�D5*�U���f��9Y�-(��j��å�Y[5j���h�t�I�����kJ5����I)�FPY�X���h�f^ ���)����Bfh6��H�&TFdw��M�Rƚ�Ys4�&��1�*���O.0^4ZR��s0n7	Z�L���5M��f�5���q���G$Ԡ��U���G]����4��ٳ��h<ڻ:�Kn�z�"��ܼupeT�I����d#*�˻Y��t��HC]�Є�1E���w��06����NMP�͓Z�л��ucGC�qn� ��m��9��aLB($q�I�o������޻w��/S���cLH�n��h,Z��� oq�mP���%G�ޱ�?�T���V�YoD&?�걢�r<��B�e��NY7tF�����V3��� ��kF�G7*泮�A��5�7/mҵx���j=�XSk[ی:i���f��L�ai�׺�V����R��� �G���
��&�M����][p����������[�;��*'j��8�-os6�r�w� �3wR� ^kxT�;��n�6�1�I�E�!V��j���� =�Э��p+s&���m1�m�sh&��f��[ǽ�,gi9�Yt���6��J	�i�X��W��e� [2����)һk�YJ�OP��^T�b�5m;#A`gN��$��fu��w�c�Z��[vr��b��D��J�M����D���P�<6�ǌ�2\�V42���ۼ�a��G`'mڮ޴5kw�|iX�1dZ�'zr�j`ܖ)�6�޹R�^��������]k�+3<�D� �Am��nnޝch�!M�Gɘs�*fВ�W%�L����iɤ�ɖe9�+(����F�|�u`�=���_>��j�4�{-�v���zMC��������m��]�Q"=]bŁm8Nӱ�v�MBm�۬v������#�m1�kt$֠��l�B6��÷{�V�x�-@�`F$�{i*�e�5S�����^F��YE���n8����S5�{4�,5�ˁ��l� Y��kbJ��y�8��m�~�
7ut�=oqƋ֞����㬷��4_^Ɗ�(i��X�6D,�H�N)F�zq��	��L�i\�e�H��ݣ]�z�ʺ�rX�u+�T[��j�6'M�j"Uଇ�lc��Gv6�!�U�X.nB#��y'�e���fG�q��2�V5H�&
��!��w����I��$��S�u��A�T��ڱV�f<gI͍�I'�,�ò֪H�	y�*M��Hf����v�t��,v̛�n5ab�2�l^E���1#f��̶L�V����H�(ˣY�q)ne�Xe�c:*CJ�
ܺwa�Ok*�C���Ո�8���уu��U�I��d�2 ��R]��I��f��5b�Tۘ�N�:˨nB��̣샑��+VMuy&����Pô��"kED�X!�lbpf����6ܙ@f`���դ��X%0ֵ��Ǚ���{U���i��ya94ݻS1��.
�W�A��#A�ZSL^L}.��d�C\��o���qK��[m�Nc���T�ӥBa:��ۡ|8�V�����mUj�]]]}OQ*���"ݑ�W^���w�&���HCڸ�K˴����%� �ϝhg8F%}�� �8M��'����;��b<�#�r���[���M�S��{�El�d�9N�*���t�*ٷE�,f^�YQk{lv �1���DcS&�e��9�w� ��aJ�t�5�R�n<Z�䂎I�H�y'��j�r�1��yhk�a���p*͠R��*�J�+bT��&�ٚ��^�owE>h1�1��Ǖ���yݠ�/^�s�����4�3�"����=fm�9x_�҉�[Q�I(��[���6���g듩��I��D6�Ђq<D���*.��a!��*��d�"�y*ɱP2}����V쨬|�pXi͖Z&zFɼ��文�谽4�'ipF�!e��I�^�eI����J�HYa��U���L���3�sY5��P�N�л8E��3(7=tڹV h5�G�З_�8uZM��"�%���L�&�I�*KE@��4�<@�P>���#	��3���$AD�O/3��@#Z�[���'k��Ȥ��=F�AF����g{"3qB+`"Y� &	BgH�*�*ik:�����!Y�F
H��d�K�`���bxMG�ԏ���ɼ@��������O����?�<�e��|1��"��ҀS܉ۻ]2�Fb�1Dz�kFAPe�h.8F���Z����&Wh#�k��>����Nf�.���W�nGQ��gX\ٴlQIK��&��n�toT)Ι�����c�����L��M�#H�XLu�Av���F��A	�:ٮ�j����9^���S�%�K���6<�HT�+'gf��/q�'� ��ۥҝf��l4�맶�f�n�uoQ�J��i�/EA����|9g�a������vI�F���\6�R�1��v�[�	¹�ղ�]&J
����<5G���NZ�v���;���fi�[����áb�HS�h,�t����Ո�o���R�_mt�������=w̗��h���fґ�Zٌ�_X��:6s��rVa�LN�C/�_-$0뢋�	u�������nXb�c.'���ӧ�u@���4�|��qΫcjѸ�kv� ��.6��ٽX�G\�.'��6���0�ԥ�7kcsi&����5�˺�� e�yv�v�v��/gG��$z�3.�ë��`����E(��[��)��iV:3'm�*3yQ�����(�E'x;)�;v�.PBӇpK�tK��层���MMe��u8��P#Ԥ��7����pC��Ә��s�[A!f���X��W/�S�x��[�6"�B=� �i�ʸ"G(j��u��"�}�[�Xq�Kir�t�|��J�5��]�f�|!׆���E�M�ط�P����	�	�Y�8]C��>�j�E֗d#���업�ȃ�W��S��cw�!+mL����'/56�Sb�d*�c�6k�'ir����nmht��-�-	�VXJ��{�Ǆ'ɡ"�Jħ�+,��+�)�gYۃ�\4v9"Ip�2����wh�E�y�UDqɔ���xfu��Txq��g�
�;N�Y�k�0�x�;��pR�Xx����X}Jnee�7s�Z=�KA[S[�mű�s����
�8
B�[j.Vm�nn�:�]\�˅�˗q
�Hێ�z���P܆#Q�n��Pv�to��wX���9Qf��xn�t�H ��3���P�5�m vS�wY�:XT��r�7��le��ٞ�"j�&=`�y`����ކQ�աꃫ�,��;!�7�G:\�8>��bG*�z�e ��[�}�c���k'	�kImôhNo;���s���)�'��f����,�_d�/�+���c�ۣ���`Z��흗E���sBY\���;�RJC�+M�h�1k�OY��@���gZ���s+RSn��J�]h��di�O&��bR
�����,ae�B�h�"��s*Y�*�J.LÉ�|�ӝQ�S�����&�nor��(�8��R��.��g5@G���t�u1�l��t�R������z��wݔʺ�W�{ ��e�~b���y;l�dPK$�:wp����Gg�M�\uۘYN���ot�Vt��� ��f�67�WoU�^T�y\�xw-�EX�s]F׊������븱��fTӶ�-;���
:GG�Q#(eme�k��\Y|Ĝ(V�	���VS�7<��b�S{)�`�u�[V	VyYA�+s��{�6d�j�4(�E����=uy�>���n��@�� Il��G�C�3(�B�ߥ����k�j<�Z+��'�Γ9�^��5�P�.p͎m�7�`JKsS�g�c��Z�^�i$`q�᎒�<�^V^vn{���,j�ʗ9L]�pg-ʺ��Rhʘ=w�`�a�y��4M��6��:7m0/i��[�� �niq�� [vEp'�c��7��zP�S�w����wD�>�sqh�8�@��`��[��2ۡbT8s�x�S|�t�HEʄu�\ƛh����հj��o{w4(^]B��Y}�<��3������^=�s6�{wƟ �#6���n�g�LÑ�|;�[��F�;3q�{���͟u�\�$��[�-�=�o�+{��4%=���qniB�������6��]IJ<�B��pX��I����Y���Y�#<�&�F�����/U��y���f��3kw�T@t/*JeT?+�8ݖ/sV-�ה�	���Amڗ�Y6.cl#;BV��mV��7c�S���
�B���k/��[b�}m�5�4���Gw+W,;0*�wQʗ�����+�Ý/���T��Д��fd{��������r5Ց�}����{�㤫�#x�b����N��j�Wqwp�B�A,�����s�FF��ƙ�Y{Hȡ��ī4Kp�ǢSd^�L�\q[��zi���R�1�3�`��RK�����e�W;!7�ٗ��-+�����8)-�s%��WV��zs��)�;�^�]���ل�E�a�H�	�4X�;��c�-`�����F04r�����ES�N�w� *+��˞��n�9m�Q�D���)�`���fdv2�}-�6��g�U�x��8#'PA�-�L;��:z�wS�tŬ�{�WA]7z�bq�K��Y�U&`�:{���r/fIKy�bbS�r�Np�T�����X��T�`(+���� �)�N�f.
#�09ۈ��jdn����ҁ�K��R����9nK�L�fntG�J������$�A[���E�CDzc����z2.1��|�e�7w�wK�D�WdU�[��\�sv.(iC&�k���at�3d�n��	nc[�qY哐|�+���ҊW��8kk�-%2dgƌwV)��v���1w!fu�*,�ܶ͡�Qk�������t�dyIk��4����%'`
��|����hѻr�ġ���o#�ܹ�uξ�o��Ȩ�'"\�v�hJ�m�O�%�+:K����l�+6Lh��m\�"mW:y�H�R	��B�yK�x�%s7&�"�e��$�ٻ�6�A�9o��Θ��GP����^�y�u�d�[si-(V�l-��Z�L�=IT�A;�L���lo7-�{�f#�����O�rk��Vms�$�4�.
Ӄ��AQ}�P��ߒ����n��Y�@�a)��ul�w��^d�����ȕC_
7��ؿ�L�r�:�v�'A�׮�7[vo��5)tmڸw7�Z�p����^�q�Г�nM�c%y��|�p肼�Ӥ���UwwE��0�9o�f@�>*�u�t�GC�vp}�e/g�ݣ� C�b���D�|+�MB���6,[U�y-��YA��o��+���n1/caisF�e΅�B4��܉.Tx��﹢HG|��_#Cy�U�^rZ&1�5��Uz�?���VK�G���t7���M�|�3�Jwwo�և0\��p���}4���qt�I��rZ15���nw2_�1�s0Z����N8�J�I�[K��=�����4F����l���R�sF�z�J���b��h����z��֡��=��|�r�3�[0a�,
�QfS{S@uo7�EP+̐��S�Lާ{#v,e���%�n9�Cq�[���耂w7ufU�2�&��U:�����fYn'p6���Z)di��Wn����n]��*k��,蚳m��H�w�i�H��>��Vŏd|iQ�N�*���m�X�|GQǳ��q/5Tk�lB���c�Z�fM��DNM��pV�M[h]e;�BK'��A%�	����j�C�ܮK_,��;g� ����pM�MɅ���5Y��#��U�Xt�����`7����3c�	�5�_>�����!ضbE���n���:���R��o���̇���R$:���%GJg6	1��*M�cƜ� 슭��1��Ck��7N�k����Z2)/tk�[פ�nl�',��\��C�L�{�l[�%��֖fU�Ř�������m�S����M	��떞^>�6rK��}��2�.�B���Uj")���i�{,g���ƃ�m�S�Z�|$�[Em
��Ҷ����K�nP���f$�QV9�D𘳫�]@sy���^���v�K�W��F�m۹O}(��gl`�r���� �CJ�Lڳ�J���(���w����	�cF�&����պ�V|ze0C��fšm\z�S�N�Ql�y�uS7(�B6-�u�N(����묗!T
+2���ZQ�!���o��/��}�Ń[y�'`XMF�b�@Ь�7��fv �<�J�R�P�X�S�L�;�&Y�������:���7�9�z��+�X���`Fn���[�`����w��9���Qu��Dd�"R:�[�funy��R=��Ļ�������a�˘9N���=,͡��5��v锥���:3����l�b��g�)�j#-�s�%n�glǄ�`�0]���-z��:�����Zy�e:�L�3b�۵���uf�ug!;j6�WVv����
7o�o9R�n��i��^����n��`�t�`��5X�����k��r�sZ`K}A��<�.gE�ms���)�]�����]m�ܚT�%��o���y�Bs�uM���v�Ca��}}@Diݶnάy�^�3��]=�.�<k�1Mgo=*u	V-H��̺[Q�ݧ��+U��!�9�,H�6����δ�O)f�lI\٨4kغf�٫��4�>��ݸ�x�[���*_�3-�J��[ݮ���<aF;G]�v��N��o�>'� Zw_���{*kϡ��z��d=��CS�rgj��Š��|��U(o;������� cb�}�W;�NZl;v�&j��6��v4�c"�6,u54����k괽|��h��&�Z��%RMwv�g[�G[�4`�P�^oC~~͒��ko��R����̮p"��V�6km�b�ƻ &�7]�Cd̎d�׫kd�6C�����L�Z��z~��bj�\x퇤=2eڽ�3�a6r�\x�hs��r?����K)�7W
�t��8�R�]c!��|�q�5z#�j���K8�V���VT��A�x*䰻�sB��PV�HI�g�����<e��m:o/��h'�/{V\����AV(�+z'N5}�]�,t)w�v|��XIVB�%Ӎ�]Hc��\����Q�DI����V��R��]�]�dqbÊ`���m:��0�����\�#ܵ�Z9Z�W-����w"�������PY�D<�ѵ|�4�^�zL���аܹr[QN���j�X���ю9)��o�|�-��5�j7K�ʦH�~A�Оn�"Wo�^�T����>B��.m���wV���Wc����V��5Y�]Z�B\��yt�8;/��:�3A92�v̞�yS����v�8��=�F��wJXt�0�����_z��`Z����1[����7b���nل��,ہW-��8������ܚj����D�J��N{�ãnJUfi��[�u���5l�giD��S�C�����G872V������K��4�5���=��U���Ł��v�!�;c�*�G����4d���Ŝ��˖��׵����m���[|��|oyujӒ�l���[�nΣ�P]^����XZs1��x�_VA3m��$w�|ցg{��,GH�7Y>/whhѿV��z��}SF��j�ɼ]t�m�.[�<�*`���4q|l�f*�ZHf�;�%��]A�z�9|�6��!�
�ۣJ޾靬j�gxܨ�9*�u�[f>-�_=7m�V�CIL��vvL(�V�\(���k�j ,Es,�JD�����N�m�
�;Y���ꫭ�����m@���0��VM��M&���$��0�RP�oNG� ��c��h��c���j��u�Om�š˒�Z��b܁=��\P�7\�;��z�������i۴c�	�1s��G{��衒�HWJ�68�2y�E�Zb�Ŭ�S�\��tޚHf�����]����C4\Ĵ���f�:��frXq�
��sg$F]A4Dg4�J����(5��|ID�q-Uwt��v� ��7�F��!���:*�)��$u^��:��ܜ_�(o
��jRWc�RW@'����ͷܙ���r��an����"��k*��k�|g78>�b��J�]rw'�� �eHpT���UjY')ɳ�h���}=��n[�:��Xg��s��J-A��\�|vH�V��e,Fnޞ�Л��
Ͷ���7��q�h>��qK�X����W)d��꽙R��8��8e�y݄��U���.�w�i����՛�c��˙id�v��2:9m.?J�Q'ws���2��o�Q�����,J�y��&��-{��7���ҭ��`�ȵ��ٳv��$�M���޾O�hjw!��؂{f��m�R#iƑIv.���#�B�m2���i�R�*4�-�]-�$w����$�S,K�jp�^lKTO+X;:��/]�f�+�@�$�mBy�//���*����7Ƕ��]�3`�|P��[���a׍���<�����1�e���z��쮍@�p]4�����x��}Ǔ�L�s�M�X�j�Vܖ�s���t�|�\�� jx˦�d^��3�v�V�C�R�p���N��B)�1o�N��ݹgO6b��i�:�q�ђ�Ry�!ݞ=��ۯg�޽���ǵ��Or��HҞ�t�l��p �'R��4iܦ�97xOpP��|{�׼���
S@����[įi�;�^s���W�|Hw�<�lv��u-��Mz��/y70�DE~ߡ�wa ���/����'���)�x����}�N��dO���K�ꌓj�r��[(a�C����`��*�akub��X7\o&�i���%YW��f�N�6�$j<!���^4p3�Bt2`y�Vk
e0�m�^(�8��z���g ׃*p�fn:L͗@�Z�u�wv��:p�l��D]���/�mv��֛� �h��R)���O�upԹX����X�]�%2%��z��tKF�];S)�ɫIm���S~�θ�����^KV���EL(���'lÊT0��*�"�K�V5�����`��7���&�JH�y���Ґ��:
��s%M=��x��B`�m�t,���X!�|���&t�5�&�|Ft���ϳ,:�+w�X����*Ǔ�.��;�@�6q�ӵ�ĩ#g-<��Vj��voS;�n�a2S��_Ig�������8^�(��Fm���XbʃZyfZ͖�и�9o�L1�P�������mf��X�G+u!6F�cnVA��NR��j�)����{+���u�������w5���Wt�s&Χ�MZ�$+�q�[��Mi�Xrի�l1S�0&�ι�-��jT��9
ܷl���V�W�7�ɚ�u��۬��\`�C��7�e��/1��-4�d��V�.CL^j���\�1��6i;��ϝj��H*� N�`�B���\owsU7�+ݰ�#�a#
�6���W!C�X�{�,��V�̃]��l�ǥ����Q�"���QK^��T���s5���;<V��\ok+���X�wE�kD�z�m]�.N�Zu
Ш,��h�hTY��LX��|�-��.M�`�:֪�aâ����Յk���=[�S	�AM5���|�U:�=)��1ne���p5�[%<��t��U���.�2�f�Ib���Fn�L]����m[�^��i�ܭ�N�9#(T���ɓ�3*m�l���j�b��2Y
�׷gR����g6>5�n�5�s�r�3�i��s�>�nh #�� �h��wI��a�Qn�ֱe:���*00X��y�Ħe�H�YZ�P��s�Ǫ�Է����9Y��4&`�e=���v��|2i� ��v�N���Y��o���B��V-�
��Pbx�A1�ae��Zr� �vf�U�ܘ��3r����N�nL ��\�KJ�P�l쌌�C���Y�k"�`��+ݚn�N�|a;��
)�d�ʹiL��/�F&����_caV������
�JٍS���5�ۨI�fc�@˻��<�,�f�ͫܩ�)��{¬�O�u1 =(4#��i�;gw��]���z����b���©��H�ۛ�w���ф�O����4��V�Κ�N��+���^�C�:�U�v���z�F��58��|��^��N������빼a=\�v\ټf�M��9(�R���J���zeJnF�m�2j�ug7:y������%��ܫ�9e��y����qU�-�Ld�3⬤b��d�il���MUҾ��xe���XԀ�����D�5�������*�{�Է�;ԏo+e�䗉��H��Q�.�q ;�ى�"�Ȼ^@6�W�͚BM��頻D�P�:ӏ�'b:��&	���[[�U���=f&^��!OGƝ���,+%����(��}�I]S^Q�MY�ʻu-���� 2`���ɕ�.�N�ס��(m⮻4�[�y�J\�;CS:�n��*:�A�]�r�eG{���r[W��oN"�tH�A�<�g�\p���r�[��ugj����d���N��`J�Q,KB��پ�����%��g�c���%Ivo> �v5���4��^<��W����}Ӳ�.@�]kJ���M;2�;������̫��b���.�+��;��(Լz�M�ʹ|7y3�+S��C/�׏V��pAS2�7A�ʡխ�.WJ�K{ ucj��I�{Ȧ�P�p�ʉ�:(�b�X)�6�qJ� �8�s�1`ܢ�ݼZ��Y`������u�ǻ�dVf���t���g�c	鍃|�-��@#gY"ڛ#8�2�2K��0�x5���q�D�S�N��JkE��Gr��(��u[�,�s"�j�ڴ��Z�V8L��Lw-(����늁5!���Da�Z�PE;�2:�p��N�'mp�8��J�r�*�$�3vFZ��7�SF���Mұ�a�w�;�^�b0�
��p���J�ĺ�r�Df�K���	lخ)�UjZ���GN��:6���ޡ�f*ı�X!.]q�)�4c�k 0F�:��+�X]�D3��z��Ƹ�:��4�<��]�6�,yN+��lb���s����,��7��o�aFv�כY\"ůk��;re
��6c�u��5�0���V�+����U�F7�:�%��'F�="��;%�t0��f���]V��ۓ+&b/��v��FU˸zfj���q�im]�ɑ���ۘ�U���t�Eǌ���L��B��F��f
��=!�N^��j����;t�6A���(j���6��,�d�3\n-�Z���rT����ɠz9
�t"!)wGD�ƹlM;�L����,[�ʑsvs��S���헰��e7s��z���}���Y�)o8Gz�����X(L�kHAu��7�ǃ�Zu�z˺�R�����L��`mݾy�TJ���@��d�rg�ƌ�C o.��L4ՙ�Qe�3VP�E����i���#�UB
@�.U�7���@Ӈ5%5�����Ur�:F��.ͬ�BL����t�u\HY��}��ۑmX�
�wMf#G6�D�=r�D}+{�f*��(��$�;-�;%7�]s�8a�J�כ���C���	�-�hޛ��U3�7��XhP�&�0��ܨ�i�W�7��\H����3�`"�lj�yZ)�R�5�j����+��V��d�ث�$ҍ`�([lus�D� :�M���0��F�X�Z�<�RZ�b��̉�3��$֛��ٻ�Q���ĳ/705(m1խ��T.
�M�bAm=65<٫n��W�C9�h�)ZN��ܽr���7Ӹ����rX�H(�֛�e2mZ�<.��F�{��2�b�,�85zu�ӹc]���I���2��1���ԕ�����n�8���jP�8��;3u�Y!yX�wڭ�2 �3��{LδU��R�d�a_ �BP�L�^ٻ76;�bu"�wܵ�HbJ��Xd��o��v\q���IZ(�����#�N��_i_.,���:�ƴ��7��x
���J�OMᇊ���G�〢8o96;Ux�h.����n��I�E���؎;��:�[W5��e�o�'���������]��z>���"�nPQ�/�-���BA�n�9U�[��DjO
Ǵ[�ʖ�����P9�T8����.$��b���1��o��*�����y�<�]Y�i8f�7����Ɲ-�	\�)��ss^^r�z5��V��p�wԁ�P�^V�{:��wvh}db��'�훽�n�o	��$�P,�:��Ksoѱ뚸1��c���ߥu
�HMi�H YZh{b�[j�RvSGd#��f�/9�����+9r����e؍�j�J��ب�6���c�,�m��C)Iw$�/��	���pVE�2ng2ξ����ʼNށ� �,�B��ݪ.�V�8�{�.���u�u4�j�U�����z��Cp���=�3
����qMs*|�CkK��R�mr�1L]�������'������ܣC�e������hp�#��B�W>�C�&X@O��:e��L����۬A����tu���g�;:�M�D�����>��\-tv9��J^4S�ee���	3��ŚސY$=��9rG��@���yT{�5��gF�^�IuBI�;�2��P���zt�1&�T�8�m�����T8n���{�3���Li���ۗ�t�gS��a�܋Ұ��Y�u����P�+��j�J��9�ۇ)��vD���:�7\��̱��0K��ZXW+y�ldu���ۧ���7���F~;`���V�r6��.t��Z�,��9��	�ғ���<�ޕ1����"f���A0$��n�8����q��!�.i(РV���*���R.RM�S������a�����%�R�������Q���H�7�vSG-�̎ɼ<����2����B�ַ�CC95]�sh�t�Jt��.��4N�'z�A2�{�u`X�_-���sf.�	b�]%����'���OC��rt�,b�ϻ�9�ڊ'f�9��iޝ��h�)m:�._6��-�j�_�1y���"����8 ���ڏ.����{��rnNz�����������yp�MIs/D���ޏ\���a�����+�p	֮�:+U�F�Ϊ|No|�4���b�6��lv��b�Q��,���i֬�8u OI�pk=Ӊ�PY��/r	w�VU�."
���z3D��&������zN���ZFvO#�~���`{uҡT�q��8�Kkv�	6����t���yY`������ZWJ�e�hUsT�{�����-�.T����c;�O9gĥ��e�v�%��1��&T4Ვ�,�"��Yط`[a�y��SB�AtA�o��]p�Y�^}Q�I��>ݨ�
��.,�l;:���-�*d�Z�/3U���P�'0�e���tV����V,Z��0_���4l��c䣁Ybث��M*���U�1�2y��Cb�+[BKIN�֌��n,��oNMy�����Ú��`�ҕ�F�JF�#� 6���[P�Q��[�CR�͂�A���E��±P��/�����H�]��mA3�R�<%�<��{ʔZ����q�����{0�D��:۵ç(w럻sx�C�@���C%I�ж�v����Y�y�����&�܆���V+V����gk��wAY�8;��::=�y��U���ikfX���Q�up�s�])g0R�J/F���t��3n�y9:�va9�wv�R���8�ܸ���2_2t�w�sWc76���oS*��Ko2 +�و5sn�|��_}wD��9P	q�V���1�Y�S�0ɶeX�5�QS��7�9�q*%�gA�,P[n=n�:�om��Jz���t�oSZq��LTB�l_��&��,d�絍�.��Wn]R�!Ge;ۧvEK�Q�z�;0����z���v+)��VJ��A�;��ɽW ��;�Rl����Y����[�F���I'Iz�Y��B�^uc�wǥ.}�P��y5UX5t�`)׷B㦰':J�sE���
�n��d*�j%N��r���ҭc����jA����������k�j��g�Z�tRc62��:�e-�]�R�C�s�Q+�w�j���N[&Õ��]m���u�V.�ū̩�2F�7�n�Q�0��T��ĆX�t_m��׻9�(�,���Q�]��_�c�ҳ�\�j�
���o��*q0G	�G̭�7lV�
���̪Ӯ�h�r�C�<�Q�|5��p�W��p�-�l����Zg^�黯NZ���S�i�rV�M�(��m!�t��tV��,=�ͧl�Ƅ�Qj��*w������V�]�;��hׯu�&��0^��HgNDuc���eS�J��9�h������oڶ>�J�U��w�Z��8�v �,�i��p4R�G6���s���=�ǫ>�ٕ��C[�;`���*Ee2&־w�d���(� ���9�$w�M��Q��l�L����d���Hi�@(fZ����.�┨�Ja�Y���rVǼ֩��WQ����T����^�:0;$H�0WN�<�a��}�\fŰ�H�/��Z4��{�����{�d凪>R:|U�~Ob/4��e���/u6���sM�%��p�Zsn�\m֯$Hr�͵,a]�����9@�{�)��5\킨(�J�S;=���ЪZe�Ѣ��v��hoAZ��9�J��OL/� �7ՓtT�[�mjn�c�aيfྜྷ�,��i��gn�h�������,�u-i�Vh�jkNy�l[Ô[S�N�L	0�}�ju�4��ml�{k&m����sm�������:���s.S�Y�;���OT�p�.�6��WY��Q��r'���K2�����n7�Y��9w�s#�X�խ������v�{-���/Q2i]��K���Y.����~�Y�*�t����Sy��>�[o�������A�-r`�`8p̏�\xJ)�R���2��U�R�٣�3�h��{-�k99xB�J�b�DQ��Y���YtFCd4�w+B�:��k�@ �	t{7;�6rL<��Qzn"��Fܱٖ:I�ҙ�$�-t�!��>�neLeb<�SY�cWL�_@�2Һ�ԠOJ��W���W��fb�U���b���e��\YiNL�*��"Z=d~�E#1_-]Kp�
"l��ܭ�ҠydU�f�P*�
�� �z8m��;f<2�C|]�{��Wsf�A1�|* �ۏ�>�PNڱ�]*�k[�-��j�R;|�q�Ҝ%Wi�1�Em��S���Z��*�92s��Ή��
�[��9��'�����NZʡ�I��	�9+{�t�]�*�+5��wj���gq;]��a7�[��������\�a�8X\�a�l=�i��1���[FĒ~����#�e���5iP5T��T�n��X&���W�t
#@Z-���9j]�R�����l���c�.��F�]��Y4��d*�at	k������E�1]q(��Y��;��ub�ݩDՒ��[�Wu���r���=��ޘy�f�8�::�V�W�f��=64^pU!��C����n� E�`��;���O� U��??��������_�?C�?{��~�՟���W����}��O�����{�=���Ϗ�~��'_�f8�(�I#�1�$�	�J��a�l*�)q&���EQ&�Q�4�-7$t|c�i�d+H��H�ӂH�&��R�&���!0�!�e	�&[?��	�M�_���X�u�li�ӫ�o*|m�d.	� v>�X��F��"�{ 7���-��0E;�������#��V�΋9�u{��$��<�'�l7�L��W��z���Ͱ�����n��p=�V
���FlլSt�
4�օJ������V���͚al�k�=��"$�
��I��gN-QK�faˬ�]�YX����2���'kD�30J���ؘ��N&��L�p�B�8��@�'{�VN�v+��v�nN�ɥy`�
G@�&��+��)e9��L���nk��;���Z�yn�k�7"����[a8.*c��;j��邶�o,N��y��h��F�+2{9�V�q_Vټز��f����H�:]ww�Y@�(,���֚��]J�'ٍZ�3G�ݡ|3t������N<Y�̼�y�d�V�O9��ҍ��ttМĥ���C%n���G�u����j'���n���Xe��:u���B�ò�M5���+�fݙ���ϸ����r74A�c�m�-�*��|u%���-4hH�o��U�^d�(Q���~�.��e��.��5�d��7�'@������>�H���µ��AsC�ђ�&��}��h��J��w�cUv�2f!E��c9$�LV��"��{d�7؆%-�Og)�;\��b[�;�����.�V�����"��
q#�b
�6�sthBp�RH"����e�BH�BHRˁ8�$�C�6"G)�da����8�A��/�"&FC��d����[�$YE��'��a��%�$a�&�$�T��q(�D���L$��#���Sp��'�����Ip�8(�߹v�P�P�҇|e�*

t������F�j�$)*�b��&����8�AUk-)�Z��D�1D��H�MkCMPP�[&���#A���

�*��h�bH�h�:ii���(JJ[UP�]d5HV�TAAD��QD�U5kM!AUT�ETX���EM)U[glPk�!AED�����f���"�֪�"
�&�b���A��52��BT�DQTS[:��B�$��`��$�*h�)���b)����J�H���*'Y�f�"���{T2 �H�f"�i���.��w�i�çP���M[o/���!+	z�dK=b͋�ű��Er9G0�S!Js�X��8��΍��SC�;�].Q
��F[�B�B�m��m�A�CaB$	i~h����/��s��������+;�b='r��.�Fv��E�l^j�^w�,�����\�%�'��|�.����m �w Q�4 ��m�z枌��spK�M�Y�NĎ�\��o���;i�8�,I��.ǒhb]�5��u簌��z��*��>��p�m�{v	6��2��V���7���G��ѳD��18A��<��l�m��Ȧ:��ev�sټOI�m�g�5�{��0��A��y��/��L�����Ng��}'��u��룴	�P:^K����a�����G�;��,�<�.��U�s9z���ݩ=0��o�ŷ�y��u��<=�?o��'���D���թ�WS��*m3�4`��v�Ǻ��l�A��d��9\ԗk����/*W�
^�ֹs>u1}�
��T�t�|K�����������S=�*�mi��B\,��B��F����F�ͳ�s7�k��F�����ܵ����Lg9S��]�s=nK���N�����*k�Y����Λ�Е�;K�fY�	�a�C]��bbb(��oup�u`͵Q�9w\�u-���[��/���}׾�����s��M�[^iW'ގ��O�#�s���Nu�󴌙�V�T��1g�*�c�:�r&9Ȯ���dv�p����7S�j�bw	�x0;�1�(��Ű~�W�o��^v�pm�sUo�}'v@}�WTi.���ޯ	�����yW5�~p&n����:���9\'EQ3�=��Û�.@�HΞ�J�o��֫�y3�^�������ӽ��T��hsd�F?�x��A�==�=�b�O4�W��3��m�w��P:I�v�T'��)5G��}�Vg��߫ވ�.W�n���v�r�<�y��	5O�s��=4��1��	����4���1g��2�+�=z|�$�0Ma�Lx����t�y�
�$c�f�gs7 ����IZT�C��72��o'�/<����ɳ'CW�!�֟��b�5{|���O����?-�]��m���s�r�{ YR]F�4E�}l�ܸ�Y�� u�"��Nu�k�S8k�{�T(t�y�K
hw7aS7���.Yh���S��q0�e�y#zs�^t�yd�^��o�L�G`�d�묃:X m��nD��:ݻ�.�~���mL]�v�O���o���CK���0�yC�!��͎����꺏.���}�O�i�/Z�ݮ��ܽ������r��c$����g��L��fR�]7u�;�e�jT�����������|�g����|�gI���3��5�F�yƒ�ݜ;h�:����O7v�۞O�.����{�_�l���������O�T�N��C�jup�r+I���|.�h�>��2p�-ћ���&3t3j����J��Oy�)<������j�'���\�p�4����w�l?<�/�"����ڴϻ$��"�1���Ǭ����w\�g��� �"C��kk�w�.|&�f�;����h��-c^A�j��"jv�"���\A,�Z͝��i;&1���U�8��Y�n��i�I_}�~)�5������혛�[������&i�LR��8p^ڿfK4(�1��{y��r����dC��_i�u�Ϳ��вީ6[^���t2��y�O5��uV�'�8\�8�8�q��^��I?o�,�w6��Y�A9������gL�mu2)�9��\�]nk6p��(a#�Q� ��;n�K��|=N�!����X��W�s�춱��Č�;�$>�>bA��j�O�?zOm�)zU��z{�Fꖧ�o����n)��n����n�hq�\A&���n��t�a�h��Gt����M9"�C︉xM�f�n�$q�28��%*}(R����5�j�������H��ν]�=^g%7�����x��o���|{'1��}����k~ߟ�ݛr�}u�^W)��fy�a�U�1%7�Gem��%�\&޸)�������������5�מP������>����Y����>���&��]�~�����7I}pf�3R�%�o��{܌��yd�9����'A���c�p�Iv 9C$m^�D\y������3�����G��j��1{�|[�@������������y��q汇tה[�����P��嫶YJ��o/i�cƌ̐c��<�Э53U�Js:ALE�7�C������!��K@n��l]��r��:y���xss�Wq���t���\}�p��cC/�d�^T�o��7Z�S�i������O���*I	�Q��hD&e!��F���x����{ۣtv_e��(9ir$�f*�,^[�$�H��Q~�m�/�|���u���V�#�2<�:ݎ޾^�.�7�y��U&\�>o5�}�,tA�vNDշ�_F�D�w%͇����;�t��;��#O�d�s,�T;^��.�Y����3d�9��ث�"$�Ћ��i�}��2	�������>���ԋ,y�m�E�ԫ3ʲg���O�oMFF��kp�Y����m�꠬��^�v���ƀ�v{rg��"��@�;!�����hq��o�� �U��3]�2Z\��[�ZZ<�z���\�8m��@݂O0"�kE^7i̪�m�͝>��,ggē 6֊�9y��Ó�66� �Tt9р����6���F�9�'���28���=�����E���xx���`��ә�sf�9B���}��Ćz��ŗ��9��J���ܭ�2��Rݎ��g��*Fu�OOzQ�f�)�VR)��|�g���S�a:���z��i��:%I���1t�[sT��������,��=��CU��b�����&1�(�9�'�͜��.�M��}�v$�;D�H:]����o��o��i�~~�����S0'ّ���j(�d��s~>)M^�谴�6ژ���o����^�V��B���#�|��m{<�ޏ�jzM������?{�O'po�NFg
����_N�ާ!��˱��k���1�ǀL�~y=5w�x�k==��uHj�J��K��>����5�i*O���ٖ!����jW��N;^��_I���~{W2�X�T
�C����q�v�����,]�}|��mb�R]qʩJ��Y$Un C�u뫁�NMz�%',�}�^�c4����it�+{��^�']zt�Y��9<C-߯"t�]1ᱣ�UAx}ܸ��q#(_M���'��V��5gs<_k���vi�CP�N(�7|�'�=���x��>Q�)^R`��n���[�y+=D�iw�`j����E�:#���ذP���+ɯ��)V
��a�Kܯn�AuN���^՞�����,�23�,v���<��r�>��^��u���Z�{���5�����"����4I�B�diN�`��9�^�����'���g�o���7��������%eR�Gy���-w)Y��z����u3�/>��xɞ^�����Q�]ly�����i��nf{�]�4n�����2`�m�N:	&�+q��pk\p��{vX����uXtü@�::���^�=�y��[>>N��:�P��>�c�����Z�j��ꕴ*�y�t��\�}8v��]�}�:x��h����N���~�>��oG���nr;\ץdV2�o��;*��M�1���1���շ�^����e�2���T����חX�'�M�8~�_��5R	����+�ߛ�ݛ1R��9�h����K�R����
^��Wd��d���*U��@&��<��U�y93�8��yO�T�T�I(c���q��K��^��F���^��/[�ޒ�!?9q��l����?v_V��!�	�A0�F����G3i%�ZEy+m�����]�m��P�b������l�f�X׍=�>��\��wS�
��������z�;nkЃz{U̢;g���\Hܣ�D�5�r-������,�W�I��S��A���=�#n���Twr���Uz�e��JM���\�p�r���ֱ�pu;<FY���&	ǧ`�^���Z�{�y�c���99(����Ak��Gy�V����M��{/�].�!����<0U_'�̌�H5�a��7U��P���m`��5����7��Iy��C���Wp��D;6�H����Ök۾%��p��U���z�m�ĿX�� ��/��ޑ3��4���8�.wK�����I��\���Y��|�����e�ԇ>����v���f;�[h�Ӳ�I�7A���\���]q�������Xu�[�`�00\$7^�mY�vI6�x�m�q�:��d���{ӆ���ù�Ь�0��^�zDXݷ6�<m� և4�^�5��K�N���x<�;G�6��]h�W��l6�1�>�L]�\ꎱ�����o8͌ʻ��I\�˦�i]�ǆ����&>lI׮X���&�Y�<�����h��V��z�i��u-�t���T���>B�f�G�ۋQ{�z+��
#jM=ٯX��:"ڎ��Z��rW-c�^���9[��\Co���G��g�S;�[��h�'����<x]��r߮��y��ԭR���vvM2j�9]�z��� #e4�S�7��=M"���/��9{f̱�qt@q{^�Ӻ/m1ӵǺ��9T�|�����Q����uI�w�w��傽<Ě��^��V�x��cv���C���
{���[��}��oX�ږ)W�XZ�:��7M���&J��6{Bl��ث�<٭�}��[>�n�d3�: `k��&�n�9 �c��j%�9��/���9��G i�`�[�8X�]{�}]q�y�P3rl�4����|�ު���M������[��G�6:�{������0=FK��=�\|3��./�_d�I��ӛp*%��!�a�m���n��v�Ψ�í�~'�A����5nW�OzV�M7�}w|!�<�tjwq�V��.�,�^��� ,��}}˰I;w6��B;`�aJ��so�B�~�w�]��O�%��ձX��r��Sx6�ڛ�f���ܟ=���`�G3����Ñ��+�K�G!��E�5��H�e�\U��vi暆��0EȂD��v[H=_U����xx
��LYr�-w2���{�o2�]���
����1�x=�=V
"�j������l����=�u���{��l�{2��m�l��[Π+�{װ�I��cS�ӏ�>����U��&��W>��[�����8�X�/�Wq���"�wG_I�/ u���O��3�Z]Y�G�������G��j������x���ߡ�b�d��^��w�߹�f:��.���)�����^�v�R����B2p��Q�$�i�o�/m%^5p>������*o��TOm��5��7��{l���5��L�P�f �µ{�;(��N>1���c?E�M��*�u,|��.�HיZ[��'��`sL�H�B/��O7�}���+v�n�oV>x�x������?���~?.~<}����o���������#�<ONW	�h�4Iv��Ԗ�����=��B,{M^�0�ӝz��"R���2)��)�in��tya˶�2��
{����J�6�X�T��LT��B�):6�w�&�Ls�WYݏ�U�P򤱍OQ��oEE��]� �bq��g�����g[�^@/�ac�V���� �L�l�Hgn=���=\�M+7
t��ݫ���mE(Z6��B]wh�St���b�ܢ�|�*�t+�n4J�c��{7u6�e�GAX�j���JÒ"�ie�/������ɶ�B	<*����R�M�W�~���LM�-ͤ�]�#�sF4C���r��v7&(�iX��5���"�1��ஶ���Gz;��Y��!�M����f;x�d�A���6޺�]OL�-�w���4&\o'J�غ2ACK�WQ�&�Z�G��9}�Ew�z�7�]k��@�3�Ս�t�e��(����B'��-�}�;eh�D�FX�7��3W
�6�iԢ�o2Z'h���E��w��Ԓ��:`�j�yܑ'���a�	c�UvD<�gL&LΦ��u(��Ҷ6����juZV�V�� 4����n�v�!���`�q���.R;���w�3yR�hgEǚ�ƹ�<�]'�Hf��r*V�*=�U�]�aH�Y:��7�ږ�2s�{o6p�+4�6�]='!����dI���o���AYg(���8��7;;�f�\��J�[��.M�d��t�P��f=���Oh�nVP�;(6[�����F��mxK�-�������DN�I��Oe�o.t[/Y�v�A4o:>���S�+m��VL�j�.Z�i*���Q�R���I�31"n�Ňk�vW����F����e�H����C�ƺuzV�\g�ZUg��w87+r��f4�p�G��yr�ӷjLLIsX�����:[�Ǝɛ(1�|�f`ņJi.�O�Jد3E�c T���6��i����d$�^���Ѭ)��}���껩1����K"O��U7s�l�"5���-�)Ζ��m=�-;�jn_eݴ�&��v�z��#�F�k}��*ҋfg]!f#q�(z���,�/w�r�ռ����Eo4��TGs�r�Ӛ���nN'j�%a׵�E]���j蝼j^����(�Ȏ�+%伛v7�����є��eo�ɏ�%m��*�7��m��te����wlM�)�o=2j9\m��F�3�& ��9O�\6���b���S��Nn��Ŋ��C�%.���^%]E|��jfМ��Yլl�/�찜�7�.�}Y�%���J"H��݋3�X�
�kB�9%��ک3t^e��j��ZtU�{J&k��n�j�'��/��o�WxW�J�H�К�U�P�����Έ�V����;�#7+58[<2�ݣ�(�j��NкyMb��va{�y�x�翿~���oU�ǀ�����gDĒQ�&(����k��*�&�����"�h�IAALQ1ET�4TI4UUUTUQ4i�4Fɠ��j*���f �h���m�Z�DTP�Ѳ
���b��T4v���h�����U=gD�bw[l�EEm��ū8h���Dh��b���N��6v�����tY��SLEP�&�� �ثY���ΰ����Q��]��MU=N�1�ۥ����"��4�cU���clƪ��cm[h�3���)�[lX��[u�E���`���m���j6��ŋQUf�IbLu�&���*��讬Z� �kTUcmcc:�Qgm`+j+i��GE]mE��L���ŵ�'6��%�Ri�������u�j�Q��k��c>��n��烷�s�|^}1����RQ@	���`'O6łX�LR�ϰ[�V��	�����pcѷ�Ȯ�W����VE�͖���3g��LbtI���v�����Hz��D��P��O�؊�����;���2�
�3��Oèkn��F�1�{�5�����7p�4P����WA
��h��Y�j��Y�k� E���3�c�_��3��?x|�1��^�*~�}ȋl��m�2� ��0L�֖�ܧl{��!)�s�������q>4��ΑN�ŴKȋ�O
�X�+�C�;�����O���W.||5�n7���CMsؕӌ(�f=[ռ�|w�����������dޡ�a���e�dE��*� �'��i�|Vf�BR��.�����b*��Y��@��M�:���Κ�W�K�����?�I���K��`���u�r�L�ڕ&��F��P|��T:��kۧ�j"N��Y��bϞ͖hS2�} 3}�guI��NV7H�Kk�sQ1��[]�gBO8�{�����v`��a�0ly���Bm�����)�Se�t?��K@�p/yo>��̋�:��x�d-xt{�o8~�l�e����r9�Ƹ�eϢ�曬v��~_�/� ��p��֧�bT�ŵ���se�{ps,i0���z,�OІ��ƃ7~3�S7���@�R�C|��VUg]4��ΐ©�yл1�}��xWn[�����	��$�=�MtV\;@QA�\/��3c"���ׂ�z��cgz�����t��ܯ�Lq"Ƽ(�����F�ˍOo�_:��	c����]NK�����Us�7`���1���n}�f�z#2
��p[�~h���U�}�}�n��W=y�����VbS�1�ם�_�������r����܅[G�ųy��
��3T��w��*6�,ke���mC'��4��a'�9�aŜ�LW5x�rŨ;�6i�Ȅ��K�6�VF�h0δBghkLL,u~��d�wPny;�^�$�ov->���Ci��S��=-�~�M�[!At�m�j��!�m��@}c�a�^�5�Wu�%�͝���L��N��V�5�����s�������kM�R���R@?�<��,"���mz�7S�Us"U�~��#��㙘_�߻|X���r�PH�3׳gV@�t�9�� ��,3���|Ǧ����i��ѵ'6����jFO�xa��C$�m��m�T\9�~���(ށ���CK����]����'�s�S�ӻ:|sϡ�e�`����*��+�i��tޟ7��޹V�TB���&���hL��$m��If����9r��Q��_S����������V�*K����5�r�q"{뿗�"y��H�t�ʯ[mf+��ҷC�]�v�S�8��І��9Iݍ�+������	s94�!5֤<ݬ�}�����Y*:�9�}9�P���~�{����O�9_��Gq�����7:d�����"��'���OcS{H��ͳС��h��N7����qp�2��v�׽��F�,`&)��!%%���t�����Y��j��cͬ&p�6S��6�0!�BuSy�d	eC��0P\%q�X��7GR�ָ�$f�7�,�xع��ib��j���j�ׁ�U�q���3m0��dŚ�-���@��x(=��«�%s�P�r�̈́���چ�Ԟ]٣ۨ�:6�(�g�����r���;)R�i�������/�5"�<v8��Uk��M��a ��^��p��;��1&{ʯ���ͭ�kb�=����-��9��Ȥ^8�t�{*	{k
��J��.͗L�9. ƓSM�ܝ�3�~^�,?����H���0o��캎�0�u*�����gv�t�1n�jQ���_{�1d�'�{�A�.�����#m��%�'V;����r�xW5M����Y�������ڳ���v�rb�lk�[9yחx@������H���½s���|�2�{C�v�g�Y�E/%�Զ�NT��F<�܀���ܩ�r�ݎ�"�T#�����Mn�Ri��X�p�7���֪wthd`u@N�}��R��ŵ��_f�8X ��o�q�E`��˄i��N�Ӵ1�89�$��J��["�z�y���-��6�0^΄C�����H�e�A�ʼ:n%����	��Yp�w6�70n��c1]Ws���ME�����"�8���� ��B�ך�i�M�鋇U�L��RO�0��i7f�;�D`��!��Eǭ�ױ���jQ�m���Z�eK.�$��������]��
���E�0m���ygo/`��>0��9�����6��{��o|d&K�1�
NwIifܺ�3X3��7F�f�A�Kcu���o"������!�$:��7�<��Bb��ή��L����*�oݤo*o[r�RXt���FNc־��z��;Ǥ8���*`����Vgw&Gc,��[u���׉��ޘ�%�2�d�g�tS*IRaA�/�P{���Z\d�l���{ﾘUV�ݸ2��$�r��Xj�h�����Ȣ��E�7E2��P�^0i�3x6�����yE�z�x����7g+z_pbf�^���z �x��w�iC����^�r-?/>y�Aoҡ��'�����'1��U���/��x]��|����#��}n�2���1l9"��3��]c�:��t;��y;)��}7��0J��ث�k��c|UE�i����S���w����nӛ-B�v�w6��>]�*��Q]���Kvd҃N�]5!�m��1�~�S�w���
��.��t�׹�^����rTz�.vU���{����r9�S�;����|�+�F�^��8u��; Sj�uQkejUny�1\���sv�Y��x����]Ӗｋ��.?|�'hs�N����'�������<h�*��g�����Z�Q�U�����n��.b�§ģ�o�3�x�K1��ɀ�぀�4B�g���o���\>E�ڒ�~uo3嗢������!�J�E����C��v�1^�lZ��!��D��ż*���s1L�Gg_��)/j��X����Q�p��5��M3�X��|z	Ŝ��������?7�d?'}T�׻���Q�������5g�*N�_��ws����,%t��;yS^fj�-K%����/�y-31B����>?���Ә���q��*����V�ڣ�M�Jr�ń���`��T���@������|��W��K�?|����
�.�ء㱆�t��Z�n��p�ԗIZ��4��t�
=�V�oYľ!|08E�=���K�x�g}>�Ȃl�y�^�L�^s'	�d�#��T��#�񹩝>z�������j�Mwсp��B�j���̸��j.,r8k���L��:�\;de#j]vR
��6P��n����@�ʝ�ݛg���7&��9q�d�38�{�4'�^j���{z�Kk��j�.�ҙ��X��5X'S133�n#dM��ۊ�������j9��f�}a�m��v�?D�I�9�N�@��IRkk�%��.7����h3�X�D�C��mi���צc>��`���]��Q��E'+�R���9��a�jy�R<�mMw��Z�=G�d0�a��y�t�bc�l��<�^Ω��Y��\b�ɹ?�d4���H��۷9�H�����=�.�C�=��xrS?rΫ�Swju����_jܤ����v:E���۩�1�"�����$:8�ՅHlg��0~�����c�O:o5�*�"�Hy����sR�2��I�^#&�ls��2r�A��;Z�  <ǂ��d�Cc�����_kݦ�����2wz�Br��v��D�^/�^����ʜtyn�~�� t� �7�m:�yg;w5h둡c9ML���<k�}�;U�;I86��0�- ��@��1`%���^�S��jօU��������������`���v�4����y@w:�P�4]�2�[޺��t�WFm�k_t�8��~ć���ʵKO����e{j./�����^���-��g���}������؁
9�]7��G����B���̷Sj�[.����k=��Vc%��uv�8��W����6a]�T�V%0��{`�����2�&?)�(�{�E����gjV�9�}ޝ�V\ta�s��`��"(��WC�D'3��ڻh����f��J���]���{g���3x7��=�θ8-+��k�?\wk9�
�b?��q�4w�0Z�*��U���o��x<!�vĽ�5s����loxoq��U��^�;+��	,���W(5��=f�2�dgO<��`���	?������F��fj�����=o,J���m�`��׆O^�YW�5��c���5h\x3ϩ�����[E�M����BP�\m	�3�wN�"�̛lg=y�e�~&):�F�+�@&��`)�˅r�a�ݲT�^��E�������1��7�R�p�;f�p����h~��=�1)͂�Q��+1�����W��ө��l�[�9��7"��oHA�'�0v!���v��{��#��&L<�l�`v-y�^S�l�)���H�t��_��ϝ��O��x ��X�!?C�9��o_)m�Cd��@���6�CY�<�Sl��ϭ������8�55�N���!��@A�ןC���B��K�vi�7�����|���UХam ���b<��^RRO��m2>)"hn5���O索���Em{.����	^��^�b��5"�x8⏁*�]�UN0E�Á��N�ze�|��74�<ֱ��4�������-���#0�bL-�	^�d>A�I�+,w���B�R⭥�3�^�RY�Au�Nv*5��8���xn]Yo�����������3��]�]S��C�ݵ�z�t]']gx��8N�yMr3���x�kx��{��7�O<nwZ�!�}�MR>6��PX��m��BՅ��Xe�\�9/LB�����fbU�*�������'���`�f!���9oF����m��P6�ָ����m��6�v����<��ۧ�g���������c��Lh�{`?FC��(K��1o4I32�h�d����~�Z�r��ba���&e�ސt;>�Ø�������&��X�,��V���4�I���5�;����%�����Pi�e��ze�ok`38�c�[ٙ�A�t��J+w��>K����z����ƛ�D<��_�W!F��b�E��z_�J�Ư� �g�᪲�Ow5�4!"9�)��D��`j�j뜩l`+J���0�*������oN�sV�s-��k/��7��}QM+࿇0G�D.G>v~��gI�!5�d&M�m}Y�m}��l�:����o'2��_wM�X��2��_����?�0��:�0�x\�Ҹ},�3{�����zl㟐JK�	*�o���xOm��g�8�L�|�0Ny���w�<�[R,��n�ךGE��.������S��X�l���Ff�r�$)���l���m��r�ُj\�c�S����+�����wIf0s��C�r�|�(��:.��t3�U�y�9X1�pU��t`�b�n;�d���oG���߾��|ʅ
%;��>}�X����^$3�7���3�� �%�u�� �I)L^��=��}ml�a���kC���KЊ�c�X���K	.��1���a*����dQu�q�:�E��\�����,�\���M��}=y���1��fDT3��:nɀ���;㴡�Q�]/G"��_��Ib�9o{��e��yT���;mr�Л��!�{a��֘B5����tf-�m���3���uzYΩ�s�l#�E(�s�N�R�}@�w8C�}9��T�cq��A�C�s��_k��;4ڬuQke~R�[ï�B�+�n��ݫ)�	AOr��4�n�ht[��� �ß���}���񣸀���;%ަrg��AM�k���U�B~���>�z��^;��w7����f~ǴB.ך���W(d�m|7�z���t6���ݐͲ;$��/�C������B�;0y.���&��|0]�婕�]��/��S�<(�|���<I�ә6�؃�O����$�6�-Ǧ�by5�\BBUn��\�/cL9��{Zy��!�zQx�Y�fY��I`i)��AyǛm������L˴�O1�����JcN�Et�0��F=�5 .&��������Z�m��?h��ʲ`c��<�ڬ w;r��Ҧ��=4d��ͣp�;�u�HE����X���R��VP��:���[I��ͼ�A����3�Ʊ���f*�&����몪��o{��Cg7S�i�p�yd��E��<4����<��?NT7$�jJ���Yӏ��~��\������-�a�@v��l�z�o
��)�=�Ŵ/>��O
�$�ڥx������fHl�y���W�j�,(2j��{�pw���ø\+�p�_��e+�˶��i.Q[�g[7�	��[�u�����?y#4��*Mw���9��t�On�us\���}�/����
�^Q<��C�	��ƐD�ݓ�v��?9�N�@�]���c?d�MZ����7�<.��T5���V��������2lƔ�mLpe}�e��q>�h�E'+<�"�� S�}؜�լ�x�����+�[u�㵿�a���D&�m
���<�^��0�,�n�]'��Nj�U�̡ڟ��Sz�8��CQiK��p����=���L�ׇ/���_x�3��\�q�|��ǫ7��nB���x^��^���Tk�)��v��ga6y��������N˵�螬�ͫ�w�GS�R�ޔϓc]�zRr�16�{���Gc<vr�@w�P�=G�
�*/���~��������Ǐ<}��o��Ǐ����Nn��a;�E���9jƉύ��C�����#�W�u:����j�2�"�G�W�rJ)�N^��!BS$:H��Ky���ܳ/m��5�F�y{�����������ut(�L-t����,�(V����75]@wI{V2�Խۇ��nAi>/HX�n�v[et�<P��2`%R�v�Ŗ�v�jy�pd���X죖��d&��sdZ�ZQs�E֎䐘�h��gm�t�,��	�\��:�����������յ�����>hΡ��/)ďv߶[�}��kgl�cE2��#F�\���n���0 �Ѽ賵���h��#zë�7%����8�.ʊ��ն:-ͺ.��aR&��a:gj��"o�:0�]��6���<sb��r���Ǭ�s.��y��h�`�	�"�嬳!��M�}f����׵3eh�=��5�N�i0S�my�bf�զ:\��m���D����i@�m޻�ܧ�H�2��ͽ���Ρ�;r3RM�(�G�����6��!�0�����Z#��/ ���X��A<���Tv�_�w���Vn#;ov����8aG��oQ�8n��m+6bDv^t�=�Z��6�*S���T�^J���
��7's��y���7#
�M*�S��0�M�ݵ��kD�f�<@a���;��$��,�z�mI�2�0e��~�kҬ��8����V��&2��u�eܵ�X�P�����9,�zM�ڂ�Q�3�xXZZ���ʟ�[����nU�]�%�Ps��R�1m�}+'���S��������Sc�A^�#3��\�܍�E�k���ީh��+](l��-Yir��t8��4-�t�L͇7�O=A��7����h�g�)��%hS�=ۖ�=��Ů��9{�L2���V��c�qM��8��cÝ�x��1�v<J^=���#&�j�ӭ�X�$��f���f`,�v�ilA�yn���`�w]J��a�c+a�$��l���j:ܮx��4���S��qY
��<gg'ӳ��Lv��t�N�/�(���CR-蛧H����vΜK�ި\��+��k��6�a�ݾ;Մ�y�f)��g+%L��*3)6�ʾ��F�q�v�d��;N�2��#�Mqq���팼)ʸ��z�كN�uq06�/L�MKu��C�l	p��ݚ�,K�]���@��۫�R;s�d��L��滗y�`�aƺ��Q_���`�òZkL����ؠ�\��b��;hq�¬s��F�.(a��QI�IZ�d�c(/�KnS�H�%�'�kQ�縇Xa9���Y�սC��Ӵvu���df��˛-�!b��3�DE^.�S&�4��I�V�=f�Õ�J��{uН���1���]7�
������,�V3V��5kܲ���6o��|x&h�j)�&���X��b��1��1�h��6j���I���Y�qQTbɛF�3ƞ�WEZ��*u�V؊���[���TE����T�D[��ӥ�CE^�D�v,Uv؛fcm�mF'Z�EZ�5kئh��Fk��(("������u4�3IU5Q���*�"��Q���Z�Tlb���$�PD�MU��N�-u ���`�&h���������]mDTIE�z�������� ���`�cX���u���%���j"���� ������`��H���h�(��mui�	)��͝j�z�Q�b�ۮ�]lAD�RQ��GV(�Z�������z�[��j���8����(���"�(��*

)��b� �j&� ��(��*������"&�����UE�a*����	d`�M���~E����2+�'O�^w�Nu�^����k�2�c�m�\��2,�6T7"�lu"�p;�܎�H8fK`k�ˤyP�o@����J�]��e��l�	�ъ*�T������#)&$�I��x{��u���Th��츠��'�[�����t�C�е~Q)�Qx�Z�X���������t�v��\*lMu@M}]f��[�}��� �+��$:l@=N×��4���O�;��9�a\Z� ��`y;:E�9�B����s�\l7���Oa�F<3ǼDv��Ai���lN��J��A����P�1%ٽ�%��4�"�i��Om=�w>iv�@�%h��\���a�c�^�|`q��������G�[3�vOc�C���kw�9[�o7�S2��Xb�9ب���h�e�lִ��O6E;�d!��["�A=v3�w�'f�CJ�{�C�p��,P�qB� ɨ%r�RFq��gP�Ο�]�X1��|
�l9s#1��dYn����f7�X����V5oB	�� ��@�U�c=��Ơ2���y�1���3q�x�+��f^@��DIq�&']�F�m���A�y�c�1I��4��J�RaLY��JK�gۡN�����y���8�$AoBBvk����nK�	ң��OЙ'�9�N�Ҷ�k�i��㵻������B�J��q��;
h9�oG�����A�ݒ�a�z��=�+')�[4܎��`KX�e�����3\�{�!G��Wt�|픡m��\�+j���4�v����Im� ���:_+5#/��{v�kV��=ӽX�V�t��!�υj|M��ܤk�
���*
u���B�나ǔ��!����?~�TV�
EB�
�]�z��Ü<�Sw	f�KW̠&-�m�)=y"h1e��-��{m�!?VԂ!��2f^
��޲;����ujC��44���t��w���^�������+���D4�^"�4f�j{�����{��DnS�K3���N���kk�l��aUe�~��MxnRy��K�CxHO��7!����c�Yi�:5]���́[56��Y�y�:]6bN���*��ʏ���@/v���v��`�kc��5�{���_�z�<`|�>|���hZ��V��������zf�ZE���ь�*9k7q��\�v'[Z��s���gCc�D��e�m{��xsP:��v_g"K)��
L��ݾն�%���nj]׋�g&;ׇ�D&�� ���vI�q�C[Fȷ��KS�W#�3J�Z�.��2�u虗i�:"��G���ևt���^�V/*�v\mEO<�i1����^nS��L� ̋!�='��9Nm�#.�H:"�s�<1���7�gOS_�ɐ��'�L�������t*���^۽�6M��_A��T7܍y��-�h��8�?
m���^�dV��9K�qqŢ$Z6�e�4R�+#�TcA��;%��r�a�A%���5}�rC���K۲M�SlR믅��		)=���Zz������2F�J����;�z�r�� � �"�n�:2�.�tz���f��C-<�G���  JʉB����������9�|y��6��Ί�?����v瓊���2�cV�!k��2���R탍r���G7V�����p�-oN�������Ali�0Y�?;V)�J�j[��������S�۬�]�_W粒�]n,�C�EB�b����TQ~�?y	�eǶ��B������sܝ�ec/:X�c\�p��T�]���z����z��y-�:A��ڞ�Kp[��Μƣ|1�)�Y�;���wL���I�
V�,�J��p�Q	�k�fl�;x��sW���8`��W�1���tOcH�B���;"��ʥC�Yw��Cu��vU��ũ�����\�_ �������7Oa�F��P���LPbӁ̓�8ӏ�6U*�����Fؚ�ӏS�j�܄Ao ���ߏ�M �==[R��1lo���vJ�/1
����C��g^�f~�����c�)ܲ(~k(W��ì7G�2���M��KS+��-��_[���nN��e�]x�%��{
�}w	��d.�48s	��Q��㿈�ﾻ�c~����q��}3��o��+�c���A��o{k4�&��|l�θZ�G�~�c";�g���L��uֹ��*�L��1����Z��aݬH���rY�� 4ԫ�XhN[�T$-9|�\\�L��H�W:��Q��+
{X�v,i�_���^��^��U)@hQ
 J >��ϳ�)�^rv���f�Z�I��Q��|dzq虞j�ܖc^1a������3b;M��=�7���_��Հ���E�IM��Z½�J���zLy��Š%��h�b�WX�c��yF�>Dn�Y�g�݅��С�ht�=�ָ�Mi�v3],�4Ϸk;I�$=- ��Nԙ�^��3F�u���r���0��g��~�<ן���W���=�ǽ��CZwp�0W�X6��p��u���5��b��p�{6��)i�5B�������<yK�*~���ۅs˶�Z��*�����j�7%�l$rC�E��cռ*�� `qm����@�ċY�g�G�m?d�aE	QCҊ�,q�5���t�
 ��Ve'埯?~��6��<lE�Y�+�Z�����W��@8�A8%�~#4�ǥ*Mw��Ʈ{gN��u(�{p�S6HQ��� `t��)ٲ�&=� ��y۞��^�]"�PJ|�5�E�)��L���m���𹗟b��ty�(f��*Y��������.�{��O�"��^��t��%uUj����~��"3���6�b�x�FL��^����Å�\!((%�K5y���]0�lZ���M�(b�g���"��,����^�H���l����:2^3�Y2ڔ9Ft<=�5�/�޹WW@돫�K�Yo=��L�[�Wn�G�!��"�J�J���<���rcZ��J�m�}%�h�:�����c�?�|������;Q�;7'E^O��edF�O�4���[�F)m�a���p'�^�����M^j�������;p���ۣ�v֣����h�m-��ޤ8���E�H�R�䣹�'�{�u b��*1��!�;���z�
���
;b+�[�9��&/3"u��"�3mY�zRr؊�����/��1�j���E�����:[
Z�'uf)޶����v���y�OC��v�5��L:�/�^������6�/1�c�󜭕E;?�,����E���p�+�'n^�>��"��T����	�t�^:i��^���I�Zs4���ij��2��h�ΞA���u��>�t��{�92���^)��{@����;�P{s�F�n���^X7��xg�d�]����/�~��~U�����4�|e��o��I�L[e9�<�#R�v@�ٴ8��؈pμ����-BNܔ� ��˴��Z��E<"��HF0Ǿ�c���E�vLm����ۜE��M\���حlNPqE�b���$g�6s]8�ΞAzw�0����N���q,�q�!8X���J��xJ4��5\�ug�9<�L�p��Vnub�Ba���y�4�+�sP��ɝ7 �y�5kr�ԕrAʦ=xVۍ7}jd���︜u�U����۞��Kƹ��W���9�R��☤n�,�z�!��F�����6��{�� "U(AR�A������o_�����HG�F�����&�G(ם�>�-��0�{N!��k���c�t+�,Uk�&�����s~�okͫ���|��a�q�&'��j�d���� ����F�,�g���0��B-��Xk%�8մ����_�~���������P~�^t���q}bj�GL��4�	�mz�hY��T���8�}�Ы�8މF4�t���2ۇn�آ3�]���U�/it<��N�ԩQe�e1C�J}	@�����xa n@AֱB~w&8$�E�.�/D��"�8n!��Pݓ=q�e�y�k/b摴vk�������v-�������p�������m:����^��溍
7㴘Q�\����I�ҒƼ��0L���ls49p�d��Dl�}vM��[� &��=ά�lq��qd�,�k^WZ��m,sP�b�j�ٺj�㳽��y>8x��}n���0&1�9�Gi�j�J�a�J����y��;m�J̹�����q��>��'�bi�V�9���(�|d@|Nh	�v[@v�a�|����D6�l6y�kB��a����?NE`6��91�PŲJh�1��=lY��ftԩ<m���@52+a.M���y�8��59�n�Rf6n�>g-��*a�L��*X�R��0���ݙ[�9t�}�Gt{�S��k�ۏ��g�!��¥(�H�ЂĂ 3 ���#��^7�^=�R�ըc�g�%Ӥ�76��0��Ɂ������~A��|\��rv�;����l3寔XA1%ڸ˱עf]���8:��ևz����Si��U�}��綠,�C�:`�Q�V�̋!�= ��T��l��˓�ϡ����3�D{�����xjq��B/�UE��^�cM�Z��/�+��r5�v�"'x���{j9��|?�񯫝�?Ņ��+�<�Vgh�R�ڔ��a�����꛼���3�����O��t����uٶ3�?����h>F����&�<d�?���M'&��s��xjZ�6��Oޔr����zǫxi������I��!7���؈��a5F�5���a����	Lo�bS����3�dR��ǡ���o��!Ŵ�9�eMs]�㗺�Y\��08s��hv�{�e'X���:��ʒT�7=s���O=.`Th樻�չ�Zf˲d3l�X"��tv4�O��.�o%�ʥY��Kza����sኝ<;�rQ��Fu]��Y�п����U��e�̎u��l������i��&�RO
�Rs�q���C�v�Ԫ 4��=g8��8�Y���4V��2-�WW���\�@a�y�� 5Ħ��5�9J
]+��y�n���>}n�=z�={��*0�
���M �"%(P�	�y�{�����W-ȬN��!��w���pN͍q>BKt8MۘhQ��(➗���[j�����d��C�1�ՇwϚ��q���������ڔ]X�:rE=�{n���5h��Ni����V[��S��t;���ť���0>H����/�s���WW�=s5�"p�}�m͈ʭ`�B�)����>�7r͵����3��G�IHb��"���z�l�Nɋ�=;���6�Ā�:�o�gӎ}a��1ۆc�,3���p�`�w%�2i����m��t�e��s�|چO۰�Gd��e��C��v���-�Y�m������u㪮�<�,}�����g!�>����t�A�����A!�qh9>s�\p6(��y��l� _E��"*�p��~0��������{{�i�k^ۼ�۞�N� ����v�Q���������
^��qt��ڡO������c��t�`�]�/L��� v����=d�d7��m�a�PY6�5$v��l�z[��%��8��a�{�w+ŵ�
,e'�����3I��O��+/n`�wi=�ɧ��J5��J��Ųս؎%�A\�.v��N	�"��<@����oy���Xbfs��P��u��R��8��L�bW�nb����g���gj9��)7�i~<o>�x7^���D�ZU�D�R!((D&B���R���P�@���:��v����m΂wҐ�r�s�ϫ�����ԟ����(1�|��Ű'�1�ޭ�z��KW(m3�9���#!(,2}	:vA����'�bY'���e	Jj����F��M���>�� Χg�@���N2��)ٲ��%��֐D�3�����;�䮑L�y��3�ey<�.��s!��^|��U���	٭�BRͰ�`����.�{��O�.��;�EQJ��[KOk�x��2�F��\Ø���o��"� ����M�1��r9��UUk2ӆy�D�WJڣ��3!C/-���Qi��.u�ˢY��@~�q6����G��۷笆�]W^�Wuޙi�[W4���\�~�(�R��^��砟�H��
#�wD��+����V������;[������Sq��e-x��y�s��Y��-ݛb�l6 ����.m������(C��Th���_�C��v��(�è1�e�c�O�l�����/�2�n���M��吚<�;d�!�png�!1i����'a��i����$���҈_��>T}�+e�,���3!ɿ�4��jW��(d�[>�,��Z'�xn��'܏>�/�`�uХ#��(C���l��ᖷ�t�
�i���s��w!p;�[��|�Z�4��׍���n���kQ�����^�{��:�u���x�x�z<���������*� � �(!0�R I(�0o�{.k{��IO��t���R~�h$,re04>(�?�ؽ�`����7>d��:zd�J�(�h��BFk���>;�|�����,+��Z���K���DL$�ZY��X��Q������p���W���f��]��dG =�Z�*�-?P�)&0y������csh�:���{�b^�}Gu�p�AŗA�%PC$��>l[+qL��vu��xĠ%���x���{V��< ��H��{`�p�Ȭj�'ֿa��q���P��N�7���׏�l��7����1l��BÞC|���i����*\�e���F�,����[��_�P�R�XSw\[gT\:���K3�sR�,�_���w<+��O�7�N�Ť��\z�aֹ�:�SR��F����I�ߣgO�"��oD�#|"�	!�d�f2b%��ͫ����;Xm��d�b9�n#`Ir{�w��z�o$m�$JF�e��ރ�Rͯ��5��9�ȗ+��r���jGeIO\b�H�9�b摧by�;�?>�O��������{��ޟw�����{���O������N98�:�y7�ݻ��A��Zӻ5��b�~U�U��.�*p�b�M��I�Ư*Xol�J����t����{��km�Q�'Aw]�Q�#ںoAT"�AU���q]�T��B�4\!)ӣF���#�Q�h�����J�ֺvrUc<�tnبoad��_6�񀻗K)N5�	3sw+2E��!Å��]u���-��w<*8a��Z��6S
u� �FdV�P�of�^G��m����|��R��n�y�ȹ���jYnC�40�d��j�dE���Z-�(�ĪQq!�tM�a��L�s�<*`�J�Y\N��.�]�s�I�V�7�5�qZ������
��������OLn�t��LU�;d���ܬ}h��{�dgnʲ�q{w��$����4�i���Y�8�S�t�X�+gE}u%����vKܬ��BN�8���wV��]�%H�;+':��M�M�D�ҩ��X��K����%e[���eu��,Ff��m�t�Z�3�/Ts��H���`NKX�V)A�Yqb�V�O�C�e��^T���u���ZrS����g7����mJ�u�5=��6K@>&n3�9�!#��Z�����yOPX���^ga:��w2����I�k�6��`2�\S�R��P��T}�$/��"t�Gec�Y�F�܇x5{���A�lT�G7�zȆe2��Ȑ���β�9[![��f����LU2�N8�;�+r��*�MV��٦�ޗ5��p��vPpf58헥�)AC��@?���c՞��7��UpV��p�r��m���'��n�EP'�a��f��['%'V/9��S������!.�i:r�q��*^d3� �rfviP��{�3 ��*���*��y��;*�C�L2�*�kV�+��ȕv�"�D��'%��^K���4�Ή@���|y������ue䍻�s-J2�����
�6��+���8����|�����KPM�G�׹L��ٕxC��J��׺P�$�� L�W	���鴰\�H�u��n%ż�'jPe�uvd�x�bzb��ܸW����+�����qij�l6��݃��*+=��2b���Ϧ���-���6�m_%�J;�P����pL�,Tt�Ml�_P;7�κZ"�ьpR=Cm��m!��wn��Їa��q�[��t4<����TF����t��b��G^�5�U8��<��Z��;W���9� /om[�]��v%�F8-v!�� \{ǈ�:���7$o�5��q��*,^Ccd�r$J����)��c�����%�����5��1�Ո����@n��^i}�c��VM�*9!f������̴],-��}ǰ@B�e��S.���N]���ڒɔo ��CV����@�YsU��ټy���xڏj��޽5�32ֵ
<�j�Kض(̓J��z�v�jh���:���6�[IQu��3h�SDT[b��H����1EQTժb)��"�lRQu�T�Ah��*֢����U�5ծ�4褣N�&����:��]F�b�5U)0M]n�b*n�*�&%)")�)�����*����&Z*���AEI�"�DEUEQMDPE1OQ�	*f)"��.�6�1AUAQmPSJU4D�Q�IM1TQMQD@�IAT�QEAQT�T�EDAMST�MPD�PT�1TRKA]��LIUQESTEE�YUTLD�Vɢj��JJ*�)����
���ZhJ���"��&JJ)""
�(���jR�����þ��^����;ڿn�
L����j�`���2𝛕�vMPr���Z�Set�<�-��=!k:
ǎ�e������)bAB�JT�iA`�F�JD~=���ϯ��y����|k��±��\�/%��ȒrS	>9+�Z�\��iIcH�CWn��d�D�:v��ڊ��[��1o@w�,��>˱��n��خu~5t,ى:��RX���Rj~Yir�u��!sj晻����1�1\0g��`����9=#�hv��D�q˯m�Hnԝ����[v��YN�A)���G0��'Z��aߧ�0p8G������N˲�VQ�N����Mrȍ�ұ�2Һ���5�~�Ӵ	�`9��7��̃"]���	��&Ϊ{z"o��֎r�u�[�#O�OK�NlwK7O�ܢ&$�q�c�LC�:"��1eyiiWq�M�#+�t �u�3�E�hZ����K�
:�N�f�Ȳ(�	^*<��L����:�e�����l�\�,���23�
�{.3�3%'�zǦ�n�4��$<�_A�%r~��OK-�q�w'���/1{�,��\:��g����w7�1���j�Ɇ���JBש��l8��#)�[bٽḴ7/-��8��^ޜa>���5�L��&��װT�q� j�e�8��р�^�A蹏̨��H����u����{� F��i`WۙAw�r���_�c��D�H��\�ˏo�Ѯ,UPzaU�Y�'	 7Y�Ylh}� J{]X_d����e�'�5�M4�`�&�D�j�b�����i����s{=���B#2�J�*�H	0)BP)*ҡB�}�W�;|~w�T�߁�	-����ё)�uȢ��z�o4��Ё�d�|Q�ͺ�.S�V��f��5�b}�^�Pi:y���Lm�Ju`�,P���FNc־��z��xڴ�4@Ջf���o)
I��	��~�pFv��wL��ĲN�<�H�`���97e�n/��1�g�V�g�u���1	�=	r�ݍ"U�zL>��(�ac�J.�s���l�Z��<�v��oCw�!?|�����x�a{�|��>���`&��4(��P�⮗�ר���f(Z/��j�����a��p�;X[��H5��z{#�_h�L#�ϧ16̨�4�^�_k���w�"���K���}�t	r@-!=8x܀��a�tz<�ֿ&�I����\����.j��Z��̪�=+��%�]S�#`\'k�;!t­��Lv����\Eb<n\�Yn����7�0�^�nMӗ�I�����gӎLG6��,Ǽb�;D�����������h!�`0=�<��|Ocj�Pݐͳ�(�_�Ǥ��Š�b�|�Ϻ1�
����������o99ma��f���)z*�L���A�NHlBpl��~��iϟ��a���;N��������`�:�r̶K�Ho�ZK�����/�c��gB4�I���Eջ����a	���vK��a�4��f���UU�|� R3������D(4��H8����/g��n�<y>=�^a�OP$3)��?��Xh�J�x/��7�1q D����KBTn�0v��C�E�I�]��V\5�)�g28� ���dK<x�--(d�����zC�+nc���/7M�!���m�;�S4/~�ï������}s�����)��(S�a�|>��/_�I�v-������mV�;����]S^�k�)S7f��ɶ	�9!�"��M<#�)�08��&���VsV�#����O�󽿣��	�'b�܄&�eMBњOr�q��ǫz����tq[ŷ�kS��=����K��x>��F�1W5?O����I�\f�_�*M}�o�@g�ۣr�����4l~��~f�!@����n���KH"}f{���Jt�<�%9�L ��0=����6�M�����}���M{9�Ly�f��D�Lpe=����.����*N�MݚN�Q���t�Kg�s{�!�<�>`���?�/�ڏ���+���X��
k��M6�qS"�&�z���'�K��ZGW�M7��������~q�J�0�y���Z�@�zI�/r���r�a���6��s�������//s��8){#ZlՌ��ۥ��G
�ܚ�(>e7u�3��w���@�j�m�Y�\ާ����Cm_-ƌ;3ޝe��M-2�l-Ȯ���@�X%D��E)&P(�	ahB�+���_{2�AX�Eı��sL��\�xev��'zn�����y�����8�4�X�
��;F:D�5"��3mXzRr�16�j����m����O.�Զ"�X��/��Ow2��O�O�~��������s\��}Bը�è1�e�c�O��#rn�P��v+�'��}���_�~����`�^�~<`�]�=h�6�����]�}حοu��MxpvT�#���� �@�%�|��-^�$�C�*�����|�c��^��`�H�q�j{WV�~<k�M�u ��m�����_�v-'`��:"���x5�%�q.9�Z7N�ka�z3�g����jq��gt�2��m�$�W��~��D`���U�Z~��RE�����g�M�sڷ��!h����h牨����i��,����Fq�z�l�#μr��R��X1�Ldj�n�9���q��<��=0x��"��ڠ��]�G�j3�L�$��KUs�s��s3��{d2������0.��q�7���c��ƨ�E��e��a�S�����>N�g��6���A8���_�
\��]9��k�5t}[�s�n����+eÑ�3�͜�w�1�*uwV)��İJ*ZՅ�a��oh�A��;�DJ�V �u���R�7��k��~u=�Z�Z)�*g1��˾�V+D!S�]Ʀ�=;׾���������V�)i(B��
E��JTh`� ���9V�w��o<��J�(�DC�۳�S_xxT��|�	���܊|�5k��m�[5�}=����9��=��No��J��]�6q���Ы�� �Ƒ�q��B��FP�h���l����R˗bɇl��&@�LP�]����<�,�"���2}�-�*�_lTM�k`Ћ;X�*` ���1��P��RS��d]ax��\�6��s��-\
�7{x�[xG
`�^p�`S�pn��K�~��hQ���Ux�yj9r�ե%�H�ch�I�<�j9��T0���H��XAa�Ǡl|{ʧ:����l��.�*�E�V��]�-d��ڔ�����N�-T{p�5�p��t���"�Ƅ�m�db�R%���B�9��Y'3��W.
�@\�,�%�T�bu�s�w��@`�y�ǈ��p؜��FI��^č�f�[���5�W��@�~�׾0�:L�sh=���pȗx�ov�x���V���3��'%���n���bK�{��z̻Ls�����y�C��0����9�?v!���+�ݛ
rL}1E/��Y�7��W]�t���oQ�NL�B��u;m]|�(/gLWh�<3'�b�4����t��T�|{+rwR�ㄣ�Ѽ�N"w�9+� ��%���uy9��-j�#w͚���Җt�IΰN!N��{����U���<�%2/ǻן�>��<|{���o��@��]�y�ۜ�9;�L�=�C�x�C�G�c�p�6��bט���g�(l^Q6���f|d!\LfJOb�/�u�ܐ��� ��Mc��J�M�q}���Guy���[=��^�tS��C�a}����Oųq��́ͩM��o/�_���P4�A�ʑ+R�������s{�BcH�0Za�s�o3�< ��y�r�aj��-E	U,��!)��2*�
ObQ�`��T1U�g�H(������y��01u�Әwss$�xc
��{����������%�j���FNc�m�'׷��a�0;�i�P�5������ƀD��ק��):�t5�IRa��"#�T���;����xmt�>\�=xk�HN͗��sЗ!���B���ݑE��R����E��,��o�{U6�j�E̹m����B
��GM��M݆D�iC��a��C=�x��ݬ�Էv#.��E��)�{߇�<��h+����Ć?u�L|"ۨmMS������a�&�nic�E�7�(�}�\�M$��VrY��bH8Щ��Y6в~G�~�v��xxJ��Mb�L�5¯�N.�C��+^r��[��U��6�P&�<˄�We Z��L��q��]�W3���n�{ϯ>�Gn��v�߻�~`�eVe�H�H�H��:]S�7��ĭa��1��5��ȯ��2��;�U�t;���4��8x܀�,�y��Tvx�ΧΌ��:���&曺����Ԫ����s�Pu�^¸�w,�C��?H�\��<���k�>�1HEۻ79k���;���*�+�(�}��}8�<L�5�f8�A�b���e�m�����-�|�G��(x/�Y~�$^��Ѵ���7d3od"����C�g.�]�vߣ�mOhn�~���-�P���:%�<������ߧc5��ɁA��v����{���\������s(��89↏���Fyh��kt�be_������2O�Qx�D>m���N8En�!�w��O�d4�L�B̖�����E��z��t��X|a������AN�fʋ�dd�*�չ:L��	����93�\9:�m�a�W�M�MA#�6->�ռ*��O^v\���Tw,����p΄�Ϣ�W���J��1����Mk��ɪњOr�q������~�����2��\�ٍ߅��Zv�]?7?m�>�Kq��5l�*1W3s��h&%�t�K'�T���CǛ��������nq�E�;�ׄ��c%��k��puF�Z�)heØ'�ӕ,P���6�5x�������F��(-�r����p��p�	G1�"/	���y�4��P����]������	���Z��Ϗ�]���so�_�V��(ZS��ռ�6fb-����֦t��{w�H02TIvl���H�iH�����'����Z���s]Q�ֹ�4��R)��T���q���m}C��Ǚ6c��N�|����m�v�ܴH��a��b'�j�E>���g��R��0�c�����a�G�9�f��gs���z�J�Hj^̔Ԟ��j�	�/�`q�Ok<�A/���i����`k���p�nYGM��������$Ȗ<�:�i��Us]�2���5�����>;�/��.g^��-T�e�e[;8\�����О�\��H�4�+���'-������)��RщSV�v��$O���әx.!�`�ySF:/Bz�k�еaD�LcYk����%�^qm�Os,�^�^UY6�t�v��̂���?���ӞU�k_-��P]��P{m��/2�����1,I��	��P8cߋ���3�އ���ygj���X�N�LF�`��2�_�V��O -Ρėm�v->�HO���ʹKOհD��w��a����^�&lokb�y[��(�5��}ԯ��/��;!pyY�����+ܥ����Ն�X�re�A�Ζ��!�h���lc�}�����jr�өZ:���;1
Nl\�u�]X�̻��fGϋrŝ�3��౶�����y��n�yy��xz�庋N���wf|Z�e�&/��n~&}r�3E�]����F�P��i�m���<2��V�7z&�9�}�E!n��&z�����=����j���ml.�pm�b�%��PH�3�Y��݋L�����]F�d����a���K��N�&��Ȳm�ڧ�B}i.�vp�v_��N�fUCtr����lEuk=lv>5�m�5��\؉.2����M�2:�[�B�������gCt5E61 hR�*�
j�q�uEê��3���A�k�L$���<�О�X2�+x�N�t�MNa2N��9�Q�j��I8��l�	�hU�o@�DcC��k�U]ީ�J��cr!��Fܻ��L4�R���LU�H��t��L gӾ[����3�Qq�3��qWvM��T��Y؄��`!�>�,�v��ʒ��W�3����.&�kQ0v�?���|3�|U�	�<�v����9;�(vt���KA�}�I=5j�e�i0�3Թ��Z���{W;ʵ�����;ܯ����P�}��viP�����[��n/��\��H���2u��zfMeT�����������:"��D��
�	t'������^��W���EB��<�9x���x�m��6+j�8Cy7�ޤp6�'�˲,�{�'Sߺ	�I�bT&�3f;�!��-��hW2�i��1 H�G�n�K@.z#�����"�!�>����׳��;��V0��[��u�$��}j�=�x��`�C�t���sL	�zzG6��4�U�����<��Hvs����^*	�F6y\Qm�=�/W�!(��9n����j��u�f޶ns���i�T;@�&��@�~����њMKsP=�/a���([d1ʦ�/W&�3i)C�F0���us��̀��cK�����c�^&e��zcm��-���8���t�5�����������H��H����m�29��f3"�x��	VS�1�&�O��&�Eju��l� tE��5�L��M�bO�~B<����S�Vov1�^A!垤�)
�?5�}���V�@e��*�S��q��������>�(~�h����)��iNwV�˃��4S5Z��g�4�^t7���cve@,��*<����skb��M���,iJ��BYBTޝ�փ�����76��%6_���U�B�ؔr����z�*���������C�}k�ڶ�p���q:�^����|;�P~BS^��RX&�	*b2s���^^�_�ޟ�������}��Oo��������{��u�$N�'��.���է���	��t��$����w6�ecw(S4�oO���S�/j�C/#t��{Q����d)[4�^ٚb')�Gw�)�A�]�����WK �����Kz��T�]y��-�9���*4���A�U^DZ��;(uZo�����(MÍ�Z���f^Y�;�!.�a����L�cA�D�p��y	Yȼ�¯�:u�_7�d�G0�XŹ��eӔ��h�x�#�4����㺷6Y��@��c�9�T�d�f�v6���^J�F�@E�3�w���J���wn���{C1�v���^���{Z1PΗ��֪^�]-��*HT텃�Vt�q�dw��Υ�:��&jC��R��vi�]�)�Y��%�P�i�pB��V *΍�;�V��,��9�p�U�sG_k�^�!��P�1��'J����5Z�a��7#w��{�`���p �ӝnq��y����ОM�5��:�M^�$+�BY�T[�x����̙:m�R���x��{�f�RҖ�jd�{R�U���)�Y��$��3���I���t�Nʳg�W#���MS��%��湐�T�v�d��Ve�,�C[T����*7�M=���W��W8�'f���WDw���੓	��ձ�x�am��8�Y�tBbkt��2Q�ªS��r:�ǽ���Q۲*�+���7u�jS��٭���/N�s���[�u�%�܇��nhT�0��j�"������j�K8��ƷI8)M]{wvJ�����:To�ӆw-�70�!��N��w�l�Oi�HQg�G�����˶�����=��CHb�e�x#��ol�H^� �r��0�9N�ʭrڻU|s����K3yõ��1��\j����;Η-X҈�Nw�%��0���΁����i��X�������:%"{�&B憪��HÆ��i��]�{�l䳵��aҳ2�X��$�=��Í6�gM��j�ab�[�-������[������\��$����j	V6���	z+Yӄ�Y3�_�t��Qud�*�b5�^�[��b�mû�c��`�q�t�}����e�]���0���38bۘڧg1P�*�37$X�]�"P�-֚���y�`�>���A��v��=rwL�v��/��1��GQG���5͙�x���i�6��L�K6yo�&���"�4�3�}�O�;g�ؗ
�zf
YSxp���V$�s�]6��En�p�3��ʹc�v�3y���X�L�1fu�t�6r�߆���3&8Ve.�89m�΅ͻZ���=M��H��`[H;��v.W:���P-vZl��XE�5J��KK��K�+�F�1�rZ�����?j�"��9ʷĘU��zV�.i��rݺR>
�_o!zY���<���}��ǭ�2M�-�q��@c���z���zu��f;�k�����3bD�$��E|iJ��ei*�����������B������%:�TSAI%D�Q3��PR�EČ�-%1)LAE1LU�DZb)����0RL�u�f��UTT=l4�UPP�EI5$N�Ĵ5BR�1%$M��P%Q�j�$�*��
(�2M|�3Lu�LF�[*d�&�������$��F��clLMDSUCKE%DDI2v�U!@RQLS%1!Ժ��bj�ii�����
�����()(���
K��
��)b��h�H�(B��ij��J���CAMQJQT�BS4��Q4PD�ӧBU%MUST�E�	$~��?Oe�{L�D���Ē �p�	���W�s�oq��]�m��u�ǽXt�y��f��A��*��sn����B���{�:�㬫0�Mo����[�
vC���5?� �)2J%'�d��b4̉Ĕ$�����y��hnds8��nZY��v�O����[@�D>C��c@"{z{�Ru��K$�tVy��$��&g��{�r�}Ɗ�q��-;���NF�Gܨ�=�XWuy�{]Z��%<T��Z�M����M��/-�oT7P0i�k�@� џ�8`|Ǫ1�������
�z��;�5���0◰�R����rPX����Rq.�;@��!�{���鏃���K�N�WV�u�]n��^�dKVл%Q�����+���j sO�Ӈ�n�d@�#�^��}�Rm���W�NcR��sBrb����B�a���~A/r���ܳm{��?B���ַ��f��j��0e���7�a�:i��mǯn�6�I�����1��3͠F�A��Ӏ�sxc��'4���LܔX(��	��
hyO�MY����][��و��^��Ir�~�+ߩ���7�i�Y�
��:Dg2j����%�,#5�F�"T�=��k���b���C���T�����<��Pt=��P�mط
_DT>�ȖxAid1�d=�K߈�7���}���e�hG��D���c�nj&���ى���$ �-�ٽbM<4tƭ��B��Qzfsy��ɫn3y��&Gh��MP�f��tӕzu��q�ș�j���Z����D�u��k�eS8��7ئ��\ �`��_S��E���.o?�� �����=��u8���{����4����WA
�����O��xi�с�Cd�ŵ���N�p��[���ssS�/[�8��)S6��(2��m�d�H}�l�|i��-މbw9��5�w�I�~�d:����)�.==
q��<cϷH�֯� ɯ��+�vu�zk#��sZ/���Q/�4�][�����DCέ�C�mЂq@��I���`������v����7m�,49Y_)J�b@�
$�g���a3��c@#3��^�Om�-�2Ү�@�Ὃ9κ�S��%�y%I����<͏P�:<��a��a)f���O�Q��²Ļyֳ=U��х.2�ăԨ�.�
���-�a�@���0��낿W�>?��'+�u�$r'(4-��ώIjo&��a��&�z���'�Lz+yH�@d�	=�8�,�gx�ts�o*�=ρ;L*5���'#bX���Kwb�j>�(�R��^���3t�mו¯u��+��ˣs�y��=���}�
�0���~4'�W:�jE1�d�5��'-�����;��&ݘ��n�C�޶.z�@�oT�$�7V�m��F�ޓ[���O�D��gmu�oK1k/�.an��ͪ	]'�gi:�D7��Г��̚��n�����/���v��I+�gee��¥7�&;��T�ȂWoRˌ[�i�sU1��8Ț ��0��:��[}���w�Yc$N������>��:��|�]���i�jL:�6��	�J��h�o.k�A.�V�4�e����A�ރ�A�P|��5�<�Mk�r�����t���æ�z͓�9'3L+�@���q�.�k��A�ɔ�h|Qx>~3`��S#n��%���M���n�?!=!27�A���s�A1%�x˱i��üxFeDy��["]�!8;�<ҺQ���p�wft�l&��)���q��`�fY�h���6�5{��i�ִ�ⅺe<�L	��b����+c�|�^
"��'^B1�y�-�{��ϫ�n�����
Ê!-@��͐�Һ��G$f����(��RΖN2��l�����a8�!'���½r	�Ȭj����a��ۓU�#OݳZ���α@���k��c�W����[���\�a�!��9���l_�Ƹ�n�����y;�ۅn��c���uk�I@J��d�P�&+!�\k<�M�Y��p���*�fou��۶T;p��md��{�Js`�BՉT�z؝�a��аt�y��׽�6�^B�J'c^��x��Q6!+���yλ&��-�+��[	I�etl��@[j�{WM���&ݮ��jWm��&*S*��D9\z�S�P��K$���%�Vb���U�ێ����
�4s��y��yܮ��0�!έ�<���� 	�7nNe�CRo�|H�A�� ���s�Gu*L��`&*ۤRzH���3ȷ.}B�^f<��|������#��� �~��a�nɂ���2�(�͉�a��MCkD1�PP�<m�u���Z����|���8Z�9���Q�FD��L%yd�yk-5��+�$�ZN_:U����;P�|�٣w�1��Zn�= l|{ʧ:������w�7\T��ݕl�;�{o��S.*��`�t�����o�+���Z	�@����Ѕ���0���nG��Z��k;r�󐦤4�VJ�l�W=����Q�$-�:��a߹�
��;�s5�f��3���/�.�d >'ʝ�e��E�5J���ê��a�i��&����xaz ��s3��`�J�!�՘'{Z�|��~`�朡9.�:�wK7Iܢ����e�����szx\c6��mר����HP܂�l�����3DawhO�,F��#��a�e������qi�Wy{p�?j��'D[*ok�`3g�q�Yq Fd��/X�ۏm z��׉�2h�>�6]�H�1��0�]g���$�#h9"jg�\�h�;�8kH@������r�G�7���]S7zs<����*������CG�4�v����RL��\{R�{��3���u����D��!�L,�p���� s$u8\[��2��"���vC�d> .��D��4�wSL`ŴѴ�uD�C�Q�.��Ǉ�wޡ�g����=?��&,;���K�k��ɒ�e��u���{5KQR�[��^���,�����ޜa�Gծ���t�<�~�"�q�[�>�{�^�b�P�9�Gl��NԷ5�%6Y2*�
Or�P����|i��}h�ւ%黜S\9�Bv,���i�S�Lx"$vW�i�y��	���1�Ov
��5IP��`�����'B{����\��&e+I�E���,F8yOֿm�z}�2K�cō4���x���؃^�og�w�7� �C��ʆ�0y����sЗ!�{D��.��[�2�e�	�����d�s�o9`�5)���ʼ�i��y���$������N��|{��S�w�^h�����vP�^&�8�����Y�O̓�$j���^N%� ��,#�`鵳�s��,��/C-n^_�����}ً`Y;B�F^�Gs�Ur��1�� �q��B��v�h|�b.2�3�n�h�)�G���s^��m=2Z�%�#ҵ��/j�A��m�8����	����ڝ����(f������ɛy,k��u�LW��>��~ s�H8Rt�St��dj�������)!�F����f�|'.�;�b._gRd��S,TA��K�gVP���3U2N�y��&K�歮\��ɪ��N{���KN��������K�'�v�����6<���(����mn)��?Y�I���O;����q��ꌳui�!��r��!�{c��2fK2�:,3��`�0����	�<�m3��݀���"���p�"�׶���t�Ws���^I�wRQ^�-l[�;��}9aC�p������H���^�˨vU1�u�:�g��L���!�qhq2�~.�۰鮯��L|�3������Sy�[�����]s���p/6�*�ǽ=#�����_O�}P|7��H+�_,��`�
�����=���=��p+kdF�i����S�O�m�RTͶ0��d�ԑ�Y���oC(A���ӥ2�q�	/�z�\����a��2��� ���_����T����Sg`��L���w�ֶ#����K�;�e�S�ʊ��*#EE�[�f���Cέ�C��>�B	��4�Jy
h�y����m�둚c~��5߃}���~��A�z�9Q�G���U��$�)+ǥ�����bS����)��&�}���ȸu��٩��m8����ޔ���r�Aqn!�t�)no}��Uw<�S�V;�%�����[熡����}w&XX�T2:�Yؚ[�i���4s��~�)��ڷ��ɥ�[���Չ����*��(=������Z�a��쵌�{��2����8��{?����4�8��_�vl�w;��O�b����E*[E�5]����h�m��bfKn��cn�=��'��nO5:���M���-?,<�_yF�8]4�^
�'����E��f�~A�,:H�C�LlK.~��n��\�c�����%�H���o]���m����ǳ��8��∡�}�"~]�B�ј�|�ƻ=)9n�H��9�w����S��zFM���'`��3��08���;c����~}�2)]�f�\or,�k��l
�Yk����5\�_l?�uq��B����~��|'�џ��>V��1z.�tyG{"�VPuKi'�s4»�=��:�Cˆ/	���7��7�9\��hʼ0j�6��3��k�Dŧ۝�����A���u�L�v��]�qr�0e�y��n6�ޣ��/M��{��ԑ?
���X�����^�m�<;��3,�4P�K����F]��MM��K�]�n��M增;3�*��L���*K�cZ{W>���֜0��@��(1n�jG�ԉ�w���F�}�׷��4ʢ:B��T���k��B�`7|š"��C�M�7��g|x	h�.X䋡�ˏP�}D��6^�ą�b�͛�w����������[!-���ꉄ�J���W!1]�Y����sܝav�U˥epC�!����s{��]��i`o�+g�f�2��-���c �$s+�.z�:�k�a��⪣��u���ՠ�2�(@�Z�	e^H��{bpTv��ޢ�����a��x�k�v�&����J�:�f�Ν�ML�z�A�=��_��ҩ0��.���z�Yp}��M���E�K[��7i���W�}�砳�D_��z���&I�9�Nl�B�ʤ�]��0�ȶ��I6�N�TeN�E�L҆��i���v�ٹ�=ԩ2�0m�mi�7 �;)>Kc�5Qȧk��=_%��1�8|~.�#��%��Pݒ��f�WV�:��	�qE��E���ƹ�9d�ZB��f�}\d�f�j��ڙ.ίP�X��aXi�L��UX��XPk2�˹��U�|{ｴ�����7!���ǣc��U9� >c����Cr1�1�o�x96�ԌJ�d�,ts*#��XI{���Z	�@����Ѕ�������-�VCm����Ô��7#��T�\�V��eҹ����P�\P��:��aߤtP��^��?u�|=����~܃P͑2m�nS����
�9ZW����,򟟽2�J�h��|�6����9��HOW<��;�ub����
�4fň<�f����H]��bG�g�Pɛ���;*j��\*�]�&�7:Q˼wɨ��b�,*Fn]r6���[׎{f�����J��M���H�~G����-_�~�ղ��@v�a�@�T�����;N�5-�^=�o3Ԝ�j�Z���L�g(���1�� ��� �������#�۔X}���]��V�(���iV��u���i��-���~|����ϴF�yO�*6��f3"���>fpC)
���]��QHgC�I�c��tM�>���yᯂ�!��ϾR*�G\�~�Mͽ�"t�.�H<�� �U �9�M�[��t�ê���X@��?��'�
{�WL�j^��iގ�6�jWFL5�j2��W�]
V���5�q�\�C�ئ{[�1���M���6-,�����q�F��s�-�A��M��L�t�.��r���ǩ���h�0)r�ɞ�O����4(���*`$;'�6{��������Ί�`[Lc��
`)R���l���!�ѳ���}Ǆ�o��=!Ŵy:A�0O���v���e'U�y�$�}�S9m���-Z��(��IRaAs�@�7�ӇDd�����P��O�u�'������p�C�lE�"2CT��e��N$~�7r�N�����֫�ާPc�u��n�r����>��=V{�X�>
�z��]�C�sd��+�}���O���H5�Y�ܢڂ����uoh�ț�Cq&��ely�z�)�+N�u����U�q:ۮ{s�z��a�����Iu��)�r�匹�-�w�p�Ђ�li���N��j�v��+�%�f�m-����F��?7y(,hj��̘C�k����n�����M�U[������|c�_���t�����YΪ���zY�|^�9��oc?c�m�>���6qh�a��c��ֿFĶ��-L�R�XW��\�
�^��@Wϸ	�h�S��)j��vz����;!l��W�0���4u|`x�n=nt�+U&7�Q��7�A�vQ����^�t9L��-�f4Xgc>0����4�	I���=��n~�n�f�N�s��U�vgܳ��^=:䳃�	����nZ=�!���xA����Se���U���B�w�g�g��y�*��v�����Hz����'��j�[�F�T?P�馉�����Gn����.�ӻ������Cj/�wP֑�������ﮇ»�䂂�_ˋ��FN	>m5,KbysZ�u�#�Zx?�&���usS��ɜm5䩀h�2�*&�&H�����~/�>�O����}�o��������OOO\߯�
��gxb|nh�rk˴�5�w�E�}3���mCk�����V���Ñ�����5�5��q�Uq��~�\�:/�\\�7��i��,M3���ck�R��v�y�(�7wQ�^�9���v����=�3O3��!H��.�a�epT�FF�n=�y[����1��IU�:�Gze��������h�*T|+�8Hft�Ky�dҚ��R\��0���f Z*�fo�s��c)u��*;} �^�Z��2�,ǧP�|.���ovV*�`Ch>���V���1�V�1�q}���**�F�z�hWd[�_P��W����n��|)SR�n�Fő��^nr�	���yP։ٕ���K^R�sOa�*Eb|c���h��E�:�_�OݗV�S�r;����6v0:��r��7���y����Ya��tr���Wx��ʳ(<�������4p�{ύ��N�&e)1��%gD�C_S�91�n��t	��0�赅�ű�m�Y�⭵N��݊]�I�o ��ç�.=�YK�ʣ�:��M�b�C�ㆸ��#���^\�m���u��Tf�<����f���N��o^]^��R�t�AC3�i���20��cdE�qhX����ā���P�H	�\�XMu;c@5�N���T�_�*[�t���"SV-�8E�)s�[�S�k���]� w]�[ԋ�u5���o�*nw>�PF�c�&wfǠL���u�SU�0 ��%�\�p�;4�|hV��	�_%/Wmu��me��t���v�n�Ͽ0���x��W\�L�/�9�n��#k���6+cp��f����Q<5h��:�ɮ�S���1T�W6��Kv�ͭhV��ݗ)�0n�Jo�>���vu�0h�cs���n:�M�c���,n�]`�wG��c��q��i����Q�����<����5�	��^楩�6o2���}1ƌ�/ke+�y�4����v;�˧'ѲWqo���x��ē\V�<��˯�������A"5����W�A�?M�/xC�9����G�]ꓡ}|`�j�59�|ήbmθ�Y�g_7Js�l-�S��^�J�Fڅ���bi�𸯠�Y}�I�E]���sx:
S�m��/E�WJ�c���z7\*蔥�K2��}�:�1g�N{��b�ّmFԹ�.i�Ѭ5J����3��֬� v���t��>�f��"�u��Ī-!�d�=G\��t����OX��ͫ�ޔb�x���-�qj��a2�M`)�v��.>��F�;�e�u;����$��kN�tF�gwR 6�N�&t� ��:�-�m"m�rFK��w}\ߖؘ����.1�d<Ӭ�������
�.tx����d�U�'c��ێ�.����S .�v�a���o��ok	��.����X��V�
��[X�ᅝ���L}����^}���}��ؾ;vh)*�f)����+��)�(
��J
��F��bZbii(�J
���|Ji(�d�
��4�SALBR�HQT4,HP��:]DDĴ�T�	AQ	ED�KKKIB�HP�Pu!H�(��e�!���ZҚ4���("�WN��
�`"�h����%�����5�
�hNѤ(�頪J{l�DSKCIE)MT�KH��!@���	ZJRPP��RA%D�H4RPR�4AHPĚĥU vؙhS��=OR�:���[��H�C�����vqN�5N/�z�踷�KLv@���"$O3+�p�F5��u��f.		�a�[u�P�G��"38��Z�c�#�M��-���3��o��Sl�N�z@�"Se�5�8�c\�u��G<v�~�Y��l�
�1�[ռ�o������%��@$<�[+̅��s@(V��wr�Yζ��	@}Q,K�Fi��J�]�v>5s�:y��A���Mf�	�y������L�I��7Y�I���)�|rJsat�eI~���$�w/*���?������v�n�Cz1��ܼr]��}%�_s�4��QX�ct�Q�[e�5c5��<�A�1��j~�{Y��5��g�q;E���ra���E��kdڟG���<�s�z�H5n��$t(�����5zs>f�|�������������_�	�L����]9���<�F���^Y#YK�GbzmE�[*�76�2�{�s�s��xwj��v���{��t�A�%�A�ƽ=Xmڜ�j\|�}���=F>����a��m�\��U	�]�N�d�x��!�]��~}Gu������ ��w�;D��F�ױǧնW4����W�;v�������y����.RSc%p[�at�����
��zm��p�����wh��Ҹ�A�����"/9;I9���2(�"v�
J�5��=@xM�ؾ��8u-�C�ӕ��-�Y-����r/��)��
�%dL	W`"=�}�V�2�U}��ƈ�f�4l]w�b���']�i/��:~�C0�s�tRN�3L(qhk��sP/��j����̲���s8q��^k1�Э���D��V'dkq���>;�B(��Yv�j]�qr�3��/R��a̯s&�/�&�s|�^
"]��h\sLL$���m�wO�fY�h��%ځSl�1����l4�xU��y���	�=i�W=�d�e|��Q�P�/ϥn�5�b�����7�Vl���r;H}Z��{ޘUه��,���I;l�m�-؝�����;�����"~�ӆ�K��\�q�	��:	�8�)#XW�Z��ZT״[������Q~�+ض.��2�\�[آݐrX��}~�c�1I��4)X�I�5.�ƯuEë|g3:�Ў2�F:ꈰ���Ѳʹ&	v��v�7қ���2N��9+�Q�$��#g[��{�.����c�u�4R η�����5�~�h�9�s�0���+	�S�b�i�swR�m[n�ǩ�C��Ӿ[��F4���B`���ga�i�)�|��Ĩ���.r`�����LU�`n���k��<`�N\��r�LʝRc�2��̯i��ǧ�}�SY>g��b�|�5n�]�2�5:� -�� 5�p�^�B�;�_R,��1�`їx�u�B��k�"��fT��[��㋟-�ƫ~���N��;ؿ���������lo��\�l��V��{�E>]��I����t"�5��E��m��jX+a�)<��)=ZRX�GjJxwf��|y���`�}q{�K���~��Ȥn�����Uе`(��.�TXPY�̩T��O�����\0g����Mɳ˴[���8�,v\,ke#�О��hv��~Q+\u��\�9/LB���'[�������2����_i~|���c��E�;.�hv�a�GR�m?Mk��ӴMKsO4V fm���C�gg��B9׾V
�a�@xy��h�omü����5ߠ�,+�ėdf�D�Nh��7��U���ۥ׊�v��E�s�g/�O���[p{�����5��C��C8�ӂ�����˹�x���Pi�e�|tE��tM�1����`0&@B,��bG�ᄯY+nr�
��Jsk�k�c�9��Hxj��]*�����4���M]1p�E3ǰAaBj���X�����'���=�H��M�ƣs�-mCJ��.}�A��ˡJң���8�E�T9�8��0�Î���5�������M�d�gطd"����.�B���.�zD����&p�=�$��A��w[�NE��)�0���/)�p3e�3-�j�>��@��>��y��-�r�i�ɥ��S��\��D�T���M�Mv������cG������p��?�h>Fg��_��#�~cb�ȋF�'�G(_C����f[�Y�n����܀�LѲ���>B|��		���ا������\�V"���9+}���9i~��o&b�[��[㼆�] �S ���ƀD��k�ɼv�3��0�h��g��/K�tS*IRaO�|��z�־�H0͓��s�ݚ��<V�n*���
��6��E�i;�yN�h�R���tS*z����KԑQ�B�_�2t�����:�)6̽cY��Nx4-�`2�ʇ�ʮ��,ŧ�I�5Iw栜K����:M8�؈ܻݽ��8����M��'�ښNl�`Z�t��J�.���R������n�C��:��{�C_k��x�L;��Aí~�٦�~���Z����A/r� �i͛T�TUX�'c�A]�S�s�:����{������VeRc턵Z׃�''S6��zH����%�3�@��>��v
>����(���jj�+L��{� �e;Kf�X��1'X���L͘L�y�
7���ҘPO{;J��|��T5QӉ:�Y�v�Ϝf��ΆΙ�О�n��z�ڋebT�/%Ĝ�:�<�`u���s.� �>�����)���6o��p�7�G}�uhz��ܾ<2�=�?� 9�Vc��H����'�x�<���Z��1^��ύ~�A�$��yu���T�su��k{�<�z1:8M3�X��OA!�qhONŴS�����g�-Xzt�OQq����u�ml��->��%�uE���H��7t�4P����R�W�0��6q>��s�a�f�|��;"�쉟�B��a�����<�����r"�5%L�xeTM�L�x���\.��$����AזN'��V�z�����,9/1q�����	_�b�=�Jly�Y�}n�q�!V��6�xb�{�g{��-U��g�>6qq���k:+y���5Jƌ/�w���%[ �'�K$���e	J�=w�;ڽ�}���|w�"�d����d����[�.i�rʬ��X���47����<����>9�No�t�~����NmF�VǍ�t4{�VR�9���b�E��y��b��R;%��%�OuI��Rr�@��m�Lay�cD���8�8�]�>~���=t!6И��;��I��T�H�M��Z~X�A.��yǟm��qq\��B�X�ؓ{��Y�h���c�W��o��N����D[�v��2�[|�it�{H�x'��y��q���j�7l�l�}�4�F�t:�Cn��6�(���V�R����OG*WӨ*Z���&F/��V�1�k����������s�a��_ݓL'z���+kO��`��˟+��;���s�����3:�ȯ4���2��ղ�d�C���x�Z!������F�˽S�W/��ي���ZqQ�����}�(�Z딜��2m�����P����"wQ�ǂ�(����^e �72"/�����w=y���i���Á}e���O�l�i ��OP�n����73���V��VM��0������=N�הm��h?Q�I���i�- �1n�����
��2"%;m҃�����ڇ=����c`k��ó`]�r8oR,�ˈUyo���gS�~�[��X9��XU.��q�T�2Ƌ|c��/��a�^�����������v��U�ږ���ڱ�2l�M�������C`����I�xC�������o�7�ӥ{ߡ�ۓ*o^��(=]�~�8A(A���d���{ȶ]�-�?4�׬#$����,���=֢��2S���B��e�a���i�	�Fq�G�v>5��sn�Ϝz�^�c�0K���|���On�ˊ���G-B��O"�'n=~G}���|�1�ڗTy%�aM���b�YR_E�1�sj\"9n��M�w75��q���8�*��Sn�v!���r�=��l��Jě�f8{��2�M[4�J�^E��yA�*�z�Du�O-���-b�1��IѮ���bj�`�����#���Ox�=y�e�`����*��.�ƯuEî��e�b�S��O�ggs�1Jא�ޏl)f���r]�vBnmЙ'�1)ՔhZ�*�qx.m�
��dM��>��#}
/j�h�g�$Ƙt���!��˷��� &(1����6v/��)��>�!X�j�jvm���B�~�!?T�#�Gd	e]����+;�q5��Y.����M�k���<�Ʋ��#i.�.�Y�뇶���ב�!���/)��F��$��F�[ꎍ�B�4�U��-@�I�ҒƂ;P�GɤK�k�`!|x}�&Ja�!�ǤZ�o'�9�]M�s�MH���)��.��QaAgO2�S�4���P��N�K��0��7�mac=�����P������
%k��]+��T�o�|Dm���٤Uz����]�{q&k����
�0{�gsH��\��-�Ø�29x'�{a���A��8Y;M��q��r�,�@���>ul4���O���&��_��__��OA����G鞧�
�cK�53Q�_>��p��-�Z7
���d�[�_:�B��gƳkB�T�hR�XY#Nŏ��ę����G�o+�B��F��T9��个[�Ӝ�l�U��is���-���Zk�8����t��q I�6���C�VBh���9q��9;��v����3.�tE���eyA�%�����H��a��?z{�j�X3	WT-���E�,�E�(�$?%��;R��C�m�{`38�P{.;l�M;��D6e+�ۺ���Sn����{k���A��B9�H��t�P�:)��̙��uwu��!:�����'	���Z�ږ֠9t����dBˡJң�z-��z���1V']��Ԟ�}�['iD=��&������b�d�NԷ5?)�ɐ�U�B��nY1�&o�������̄5-�׬z����v@�2n�I|���W�n����L�Lhي
�%n�Y�Cb��!��c����T.�g1����;�al� �� ��;�LhO4�0V��[&�W��Qu�̢Y'X�ʀIRaO�|ᮢ O�_Z �a��Δ��]7�ENw^K1�I�_Qw��]0�ީP��U�P�F9f`��=3��c*��aQ���ޗ��f�^������]泂v�8�����1i�����ߛ��w�0��_.U��]v�Y�v�>���O2+�[��硼m�dj/��E*xY��߻����οma,Vd����h�aQ_g@3M�rYLe0�!�0 �/��[+�;3���Z���A�%5�o��6���zg^���cwS�gNA��\��(hs���S�y��>��:��u`���t�%I�V��hԍ�j���⓵��ܾ�9���5��á��#X)a�����;4ںd�2�*��zW?>;U��x%�ʚ���O���K�pZB��m��l��!�\9�����_4wnt��`�o�ȃ5������u.b�§�J}8��'��'�<�}<�Ip�	��|��y���YM��g�_+�"�w&ǥ�C6�Y(�_�Ǥ�qhIy� tE�j��g�]�,(���`��]���;;Ts�R��N�k�L�9�l��$?pF��S����k����0���0�9x�ޡ]�-����<�!帽��{8;�kH��L�^����WAP]Éuꉾ��V.ۼZ6�ǰ��_���U�������)y�����2���Н�2��;��	̵����k�`�
ݠ��8�����o�T>xhq������U��دwwn.e��F)4f��wCaׁ�5IZщOҌ�
=�Bޭ�z��'�"X[�y�a��¼~��?���3�_��3���@�=#��y���,�q�n���C\�L�H� �2d����l��gN{o!{�ǹ#�St
�rؕ���4���<oqoU�b�F-�N�@J}���m��e�'0���ld�n��]˧�W�cΙ��]scQ�d�Y��u��B�~�

���0�qDĲOa#4�ĥI�߭��?
{w�\gf�T\�b��f��u��DpW�p��W�A��z�)�|bS��S*IRkk;\�����xf�q�8��tN��y2��
�c�v�.�M��q#��$��'+<�"�-�Ûe����5�̩��h�k���8���-�O�����k��;Q�;��Qs�!��6��1i�V��V�ف�����k0?Y}�C5�<��a'�?HdH�G��J>�����(:�Q����s^��-�h�;F]���~��]���_{�ܾ8���z"(���t!w)��'�S��\��}m��~g�Z�"nm�;�|����*����ROx��y��?]}%�ިH~�B���
_Q��e�6n���˛$�d��]M���v��D�^c�^��V٠+���_P�n��aK�=����=��d��B-��C�bz����j��vRpHNf�W���LW5�1�b���9[��e���֎�����ߢe1A�E���?�z��4�������Ρ�f��q�b�=���{�|��o����������o��x�=^�W�5�����'A���H�ऊsϵ�2�;NK�|ECz���hKRiǪ�F�}�:=k�p��D���׉��kF=��:���9�:*[�t�s�v�6��q�����حY������;{]H�4�v����*�+W���:s(S�|�p�]8SKx���B&ԚИ`��c$E����7��d�Or���Z�q�j����d��R�"�3�u���+վ���\j%�s�E5�;�O�إ��|p8q��; �9��ϲ���Y5ע�0F:��i�Z\�cke�ы3�o,��4��`�/ O�;[��S��g_e�T���
ۆ7o3ho����d�o�]袶�@�<׳+��F��f�a���Cb�<0MZC�i9�,]ݣ�&mqu�2�GJ���wJ�[��}b,.�T�3�tZx�u���&	��	����]�ѯB
�_t=x޹�ٽ�ۈg��!�c�{A)X��MGXsv�[f��(#0�BW`��*&����v����ή����������6����^Liܙ`��16�V'n%��{5 .�\4]�]����뫋� �;2�Ãvf�����*�P�4��X�Z���],���8K*�;Nш�<��I�F4�e˴�C��;����LiqE��i�]Ӹ�BM�72u����,Y)�)C:�
�cK��Q��Ԍw�xv3.������U�����,��0����`�&E\���ܼ'*C;[��4jT���vk��;�o2Y�B.��o**�f䕸HP�s�j�E��&�� ��k�_[�+K����i�l?{T�NO��7E��Y��#���(Elt���:�����\s� BetUX�u۽S������v
r˵�z�4�AL��>'���8Ԭ���gc�)l�٧zF }�p���]^Nb��sb�֜o�r�M�c�s�����C����n�o[w����M���~0��|ks���[�f�%����S��z�W.*����7���'��ˮ7,�F��K*���ڼ�&�{�ȥ��-n�wr��h{�wBh�X2�NY�Y�c��Y�a\rE��ŋr���b.�,"�A�%v��:{����O���0ZtM�ŻC,c{�up�UҌ��(��Vո��Ǎ>�{���gS:�i4�֬���%��z���%�1��꼤�JkV[Λ��
��>�H@��٘�<L���<�ʎn�;���ꭣ���:�
\�)�&QMs�hJn]jѷu�LY4c����A�Co�ҹ�u�L\[W���
�VJ�#���yu/l���&#\l��C0Lb{�Z&�4��^M���������|Ul�Lt�oN][��K1J�A��@wNN�i,������%�ݴ�G\��7���	�X�Ǽ�t����dѹ�핢�-ာ5��5���ѽ�f��c�T�i��t<yI�ʺx���xzn�x�ýO��ק����HO{  x
�'�GBPPД1L=��BP����B1(P�5EABMA-��%-!B�+{�b��X�h��"JB��l�֗T���JJF��(
& Ӥ(���JA��M+��ZJiJ���`4EHkAJ큠J�)4�)І�G���������j���j�Д���4��@Ql�(�T�K@���Ӥ(�)B�
 ��҆�ZU)I�a߫�Xi��M��@�mF߅Υ�7k}�
,�˵Ͳ�c{��5�ffWn��	�+�us�BY �q�����Pd�:gU�N�Ǽvp�lY�?˄h��L4�a�ȑ/�Ă8�6���đ2$��j���������f�SD�d'*� ��k���;򯔴�C`�?�2��o�?�_X�v׻���i�M�~	3cvJ�O^_�������e�m��=y��I�&E;�A�xCV����\�]F�ڙL|����s���]Аq^ �-^+$�Hŕx���ŕ�&,y����|r��r��E�w��v<�x03T�V5i��X�'X�%ӌ��|jQp��3�e�b�K�5�C�e?Ѭ0zB�<S�^]�Ʊm���OЃ,{&):o^#"�)L%�vN3a�׋2�4�^L]�E��qD=��D&�
Y�'lr]�Od��nt�?x9�N�hZ����]څ����ɲ�iq�ѳ�$nE�.�o@Om��C-�v�ٹ��*S.-�m�Լ�ӛl\��So H�z	@����|���A�z��B`���=��)�țYuL����n��AvX�Qz�T�"� c�|1sH���zw�~yp�Ѓ����\�ޔT��h�Ӌ�_���w/čS�$���U rW<�ʄ��),Qن�.�A[����^׻&ve2�G~S���jqY�Ҧ�h#��j�ݕ�����b\��>5�e�=�X�0_,ԧ7����zkڹ���^Al�<�R2�6��F����bU��b~���|����d�Y{ U��*��s�0[�t�X`��Z�t�b�<��W�\�1��?��g��Mu����K����,ts*!^�ل��}j�^h�Y��tf2�E�cw�2���,ZD�tm��Bը��8.���A/V���\۽�sGކ��uW��c�\�Zþ�XC�a(G��k�P���קe�m{��c�H'��k]��̆<��eOu�ܝ��N�(��-K��׋�g��D�����!���]`L������r�/�][�qv��ڹ�̀�Q�~��U�H���ϫ�����@���S�z܇c�ḃ{פZ�j�5ص�Wf�Ȳ�z!��@A�v�"�Pou�6�����*�{�e�3����G�~lP����s���o1�fB!ᯜ����C��6�e�j1p��DY�4�Cst�^D��l�X.S�w4���cW\�KcPT��xaU�B����%�u���}�~�5�0�銇�Y����Bk��أ.��nf�!5���Y�R�w7�x�:���k�˂�^b�b�L�J�,|<��>BygF>CNאi:yy�o7��G[�
mȸj���ևu��u�,܃�5�BD�2��b����o+����e���4��W����W��{ߤ���Z�X�����p�4�TFB�p�*�:Kc��7z�e��-�����G�/���|�˳�����>7H-�
��8�=�L)K���GŴ���.��3��V�8=k�<'�[�	-�:A�'}-Gs��艪�ѻ���XC��.^�t��%�u��L�R�w����=��z��$fÙ��3��T�ʭ���R�1��"U_Qo;OdQt��*�]ctS%�0��0i�S�m{u�
W$'fU��������K�[("u	����УgiC��*��f+��zq�}�rU)೑�y|����a�6���݀w]Zu��&�-[B�Re�YΫSR�,�\Еf^^E� �r��z4�zp��W��a�ã��ֿFĶ����Ԫ��
�3��ѹ��8bi#�VS����{W���E�~��
��'������4w��*{�UX{�!Kn���k�W1�S���}���9w7�}�	�y�(�y�W0����b��V޻T_|=C�>�VKH��u��V��NI/�Ǥ�- �� �b��!��üԘ��!�\��P� ��^�SJr�5�\�	��vq��i�C��� �=.ŴS�g��J�l��l��Ro�`�� �����m�J�$\sm�;���;<o�ݾ�4:�	Ltz�|�u���G�5K��ni�P�ٽ\H�0є�n���k��:��O���h�HhZ+_o �i��
el;ݥ�[Z��w?���_g:m�y��V�E�/��ש2��`~�l���ǳ�;�i�*�Kx*� ��@Ύf��5�a��c�:_�V����R�3T3�'�0���?������K�ܙƭIS6�DW7V�{+xw[���V�0֠I�C6q=b�O�$������Hh�~t�NL!(@˳�K?��+�6%{�݅ܯ^�#(2j��4�ģ8��z��x/B��$`�ajm]FG��խ���{P��̂:y�����=�f�\���w���It	��=Լw�1r��nk�@��vn�LƐD�I�?D�I�9�NoڤS*IRkk����e0�̼q�>���^�6���ɳ }	�Od�}�`�I>9�NV7H�j��K�gV�Fޥkd��z|�>�E���1�nb�0b#�vKR{�ޘk���]ZR�<��_ݾ0�����7�\�O�[���	���I�u�L$���Y�|�Ƽ9�~�}W(�މ_z��uc�e�i�e��I�jF�������,Ht�$X��?��Ѕܣ_��<=t�����|ӯ��	�M�p5����1�&w�c�+.�8�j f�Fg��i4Ⱦ�gQ�:x���o2�S�f��X���(R����B��#�S.���[��Q�z�t�q�c�pU%Ƚ�@�:�"7d�xx%��!�OJ�p`6��Vi���읈�i\��N��:J84�]��n��B���M��ƻ��I�Z���j�Ʀ ɪ��h}GEC��ߘf`����zr\�Yn���Χ�6��T-'�Â|e����@��H/��6�;i�h�+fE�B�u_kB`�C������t�=;_hv�Ge'����P�����F+���جm���9\����{��,�x�oѐ/��$�b�7s�P&�a�:���d%X�o}Oq���\(m=���p�ʹY^���`|e���'����bs;��=M]�s[3��[�E���S4�W����
���r2�>cM��r����'�p|�ջ?y/��Oݸ�^q������W�m�����b�\O�t�]{f�/ΞKӽ�q��럤?�����%�ٗ��x��9�\�LcͶi��Z��	�� K$��>��q?��G�>��O9�q�$�A��^�sa�lᐆHT��\_�㝱F2m�����2��L&T&�Ŭ�E�5�u��y��d�>S�Y���]Kl�C�Ol�8AoB�,�S	;n@����Ιb��[������Ū��+��aD��͛7����J�������J����J��<� J�v�+6a>�>�r��Jܺ�iA.��κl���VOgڰg����ӶQ�q+t��.���c<r>w�Uu؇)q�t�¹���}�/��}|7�Ji�r�n*K9w"��_�/<�+��q�~��1�Ǘ�'�e#n]�6�@r�4"�s����C:����\�6�IB����l0�ǖ�n���i�:/���~;��Pn��n��l�Ms��B�P��R���E��	��cw�+� �T_��?�Wm�"%J�.[g��#K2�ӎ�KT�6w��XV0�%s�P.R{	O����T0L���;!����$���k����o`C�`��1 �/��]@�qvJ��gG2�S�{mf[a��VU��N�Z}�F�o(p�	p��1n���qR��`k.���Q+\W.��`�%�����f�uJ'���lms�������n�z��69�6���vYCr���u*�w<�)��zP�ݫ)ב��M~�Cƽ�g�yX+���2G�sC����]s"?|���9��R��p��bUk
F$�P�.�\���D[��r��yw������u7Y�^�f6�f��|�_Yy`�u�c���;ّl�;dw�`�I��=���yxn�3�����N�=jF���}7gǇ���熩qr�^ �ӹwl���*#�Q�6-��ɾ����n(7Н�K�6�Un��z�r�ި	�ل'�����S�oc	i�4��0��o&+�.��<Xt��L��s�
M�'eLuQ.ŝ9��ps��Z��͜��������H��/]Qx��7gӍC2W�K�W!
��4�e�n��z�9�9I<N�Q}��.ǈt9��, �8���/sP'�r���jR�A���J�o�`�r�OB��[N��$\�C��+������?4# Ϧ��*�Y$�:kxr��3�&��7p���3H�勨>3�����d9P�P��`!W��A�RDF���G��wZ�r�����{�qXCq �$�H�J;���+��?�u�F�5m�S�`�|���2o$�7|���(c	R�2I'��2)�F�	Ύ�w�Tgr�E�^�"���y���ᦏn�"�7w/uyۃ�g��c������ɍ;�Ѝ�>������*��NE!gvj��i���,���ca�(`��mdAU���Y:J0�lQ��=W77;��{Wٝ@-^4��롽7��ޘ��C�Q�z�"1�Qk�_ߺ����w���YCy��f���u�=BeZ�Bιk(��a1�U݋&���e$�kV�&��BG�ۻ�������l�2�w��"=�3o$zP�j:�H�O��U�ui����t�0?���������{ۚ�5�8�B�����&���+�����jK��j)S��졶���`�8�q����.�
�Yuߺ.���)d��[�g���9CyNP&:A�:Clo6�e�zqXɆ��9��i�+���\���#,��6A�������7�K��1�롛W�o�^�L<�z�;��:��p�xV�F�y'
s�=��9"$qcӭ�A��Tތ�}�8��������.,�rs0�n)w�o(�k�� �(w:/o�!m�3������]��vj�7�N�d��*�����7#ͫ�rm4b�h���������$�T�֜�W,�e�����re~�h6��M,�q���wbx��>E��PSJ�z�x�d�sNd
T�Uv�}�ƃ\�d�L��Z�÷N=���
�L�A#*���۽T��6rKA�f�u7+H1���N9"
���ˤ6�i�WJ�J�����߱�F3G�S��ocKU.��2��,��#=����F�K3陵.!������w;����޸�
�kE��V28d�kr�;�дR���
�:�!�Iќ4Rݬ�:�,��;�I�ȅ����6r�N�)���y��� ��gj.���᷊�֛1��(S��(�Z@��ob��|-����m[{�Ғ�ܸ�cӾ^�y'u�go9����͟aԨ�3��x�p��o�~���N��tr�:�}��j����Æm�����	�mkdzGe)͗�!��r:�au������Իq���6�ԭ�5�^y#�w.��]�����r~�CD�b+7�k6�P=N��L\��J�\���R�1@�5#,m0|��ʆ�g�cu�qV�kH]��=";�p��`�Vo�; ���)��vy��{��s�6�O�W�`:�_Yn���q��UŎۧ��r�)��_{���3�@��@�]�WT_$�w�r�_T��.+.�N�����/Z�FGSƇp1 `�f�T��\��M��=��\�����m���yH� �#O4r��j�t5�@o-{1	Hܑp�9��On��#�=��X�v���#\]N�S��m���y`Nz���:�2�A�on��wA�_;�����1H��s3]��WK2 ��7H��m������Џ>}fv擧�څ�MA�l.�r�Mѽ{�>���ia�ϳ{ݷ9�K�4��b�#��"�ܮBK�
�R5[��cЦb:��$���Y՜r��F����q9����%^Y��!�Z�A#�z�Z�Ȏ��~������Z����"�&p0+�b:�E�F�b��*�J2(����{j��.hXm����71j[��/SL�Р��	|6��ن���,��1`ikp=����!�'H'��3�=ڑ�n�vd"�$����`7z.�F���2˳�l�mwC����Ô���*B$�ml����_�##����Q��sjw2��1��(IjM�_�
�i��jK5��z{�@0�j��B�ݴs��7�Oc:Df{�)6����+��.�(g�<Sޅ��2f�IS��g�4�Cpf���{g}EDP�ʯw.Tw)�n���:�]�1[5�l���`��1P5�`W>v��� �d�ڶG����x�G�����{���g�����_�����u��f�e^�j����7{^*��,��&*O�=�t��Ɵ��vӐ��c1ͱ�x�J��Q<��(�m#�q���˚�S�M3z�7�!�-�SfYK���nׇ������V�-����wٖp��J�}�+�yN���)�Wͳ�#�Ll�aqV�IcU����]|ŏ`B�Xiܦ�K��c�t��|��(-�c�&r߰�Ǻ�e�nVs�����f�������e9�d�_��ε�n��6���w��|�n�w�3�m+{U52`�4oE`���;���kI'�9��>��,�{y�ށu�ނ	ƕ�i�	�h�t9h��)�Ќd��IwC�i�o<ZWmѡ�j�(�pdI�lZvq$��o�'ZdB=㬝��ju�[S�̼�1C;y,L�w{CIՋ��̴z�%��Z��b��T')AQ�m��R�ɖ���f�p?:X���a蔹/�Iђuk�	xa�ϰ���6��@+W��ڗ3J���Ӎ�u��f�Y4dw'H�ݕ�Reǜשzs%��zWX��m�fS���IF��ɦ�m���=n�o����5`\$GTk���M9���E_^^�h��e��P�|�2��E��u��pdH"֍w�a�E�rUە�״���:2=%���v��fP��S<� +F��;�K9w}�Eu&��l�21g3)�޼}��:ymoIƵ�X;Y��pr��E%�o�g8q���"P�+��0MMZ 2��E�!fX�9�|82�݆+i
�Z!�M��b��KH���짏��W�&��c�CX����2�M���� �xh�՗�z,+���jQ+U�_X���p�֯%Ѝ�gw��t�[��C�<��B���^c���3��
+��A��6�nsZ�<͹���:Ŏڼ��+X=S�X]��5�q
JW`ޡ]�fG:k�ciM��hh,:�����+���3)�o��co!Sf�!�2Z�z/!2�w�]�2��|s"<ʃ=ջ}�MH)�b�s9���������:��7�����Ո�:[6� I��k��J��v�'K�s�	����U�b����T�	fj���M����+(���3���Z�&	|Ml�G�PkqnK���I�3gI)�\�/��b�j��ۻz��,��ճ;F�Z�a�������s3��Ŕ����W�_)�|�k0���;���勜��(l�e�h��r�&��ך��@�Z��M��k�6�u7U�:CUN5���s��`�)��p�j�����snL�k#V�L����k2��}�c̙h��5��a�e�6�qT�n�ExV�o��+Y���sC.���QFs�ٌ �k�Jo��+����귾��XWàt��qW.�gYu'� ��ǆ�bz�H+�n��8̶4�5��|��,T���Qeaݘ�C՛�wj�}nBF�����Z����[(D��$�&��
CHRRZK`�bhuB�C�4-�ѧJ���lhM��$JCAH��ӡt�Q����4�CB�&$4���MhJX�(I�K�ֱhM)@Q�)kJ�S@%��&�m�iMB��*��ĥ:U:Zl��Q)�m��tWC�&�-(�:v�F�6�l!�)MBi)5IJP�((B��Jt���Ri;=>|������lx�y��r�价�-��Y�� �I��TD�w@�����ī��ǖ�0�y� �u�t����Ŕ� �a�4���fm�6���hoKu�s@Cz<��W#/�r%��6�dFD�nڻ�~W��[����,���v,4l1�8���_Dx�,ds�����B��W����`<�$O8K���i�� d�W���S;x�Nԋ�$��»�ã2�;x	$I%��kC�3�Z�,H����7�2�'D����3��]u���C�q�d�y0}�𠧦kj"�[]Oz������	G��Mz&;-��"��C����;�]�ؚ�a�;� +�~<tM���z�#oQ�qbU~Bc�C�v�{�s��������,Þ��Q�ͻ��7V����K1!��=��k���y[���@e�D�,PG�ǹ'IO �w����i�;/X��	_g٫��+�x@��=Ғ����L�IM���N���$Y�k�-�Jk7��n��٘���&pK[6BեT�a��f�|Y��趜m�x�(�w�wn���m�%��q����t �
��^#+1�Rc<��a�j�X��QQCN��)���눡�Pb}���U{���i��s��w��dgt���:�2w%0�{��c �J[(�-��r�Rҥf�n)���p�^�s��/Dj��W'́�5l�s�׎'�Ek�Iչ�`_gb���[���^�W���<��V�`r��ȃ)��}��մL�
Fu��m��d��".:��v���cۮ[˷����P�o?�o4>ށ�߰��ݗo1�����v�����'�(��9�"�e'��0:�:2ɱ;o6������ce�:�n�ةQ����[\vr�Lt�����_��b��eb�S�9����Eϝx�g� ��&��a=^�����d�~�� x�����~QA�����#���7���;���@;���(H�oqU���f�{�l�HdS�;R�B��%�������.����$�kg��Ջ��A%�
�R6)́��c�O��Hעz'���%�[�[����R��qU���
E+�t
K�M�7j�o5{.Y��luD�a��i�AhE��6=}�r�Q�3˺�+~����SM��>��ӓ�>���G4X�k�g[��'u̼J��N,T�Ƶ�lsT��%j��»�YˋN�S;�:.��h�	˼�Ցb�C�Nv�zD���#�%^	i��ju��@��t��*����R�i���9׊�[����B�P]�Pd��z��9�B�����ƈ��&��� 腓�ӥ�n�
�)W�'���U�܃͏scK�����J���zk�NJ���"�t��hy�Vqp�
��(�e0ˑ�sdcWl�l����p2������@u����ڤ^���)+{lܵCjt�igg/���|�uf��rA<��^'��x� ��n8nۘ|���
�^�FUm=�c"2��8��*�$�K�v<��n��� ���c;�n�5�>�T�U�w�3Hlԓ���5�(���s{�	mp�k�L���dZ��T�⡧4�I�'L2�J��4���ؖg�CUk�w�ʦ�]�Z}A�����L�vH�4��� e�x�O;^C2&H*�}�BDB�������C��҇V��b�WY�3%�eIj�j�?=�Y�����ݳmc%��P���V�l��=�ʻNV�ә��X�.�hq���׮붆]�I�3��9����f@w���w�'K@�<m>x���QX8y'=U7w�u���}@����x�����ۭ�ç��V�mdV�[uW�.�t�kl1��HA�t6�i�|��]B/�]ëfc��MM�yG���l����K $��G����t`�gH�\�O"4Eĺ�ᑵ�y��y@�>��H�Dxi�s��ث� ��4�C�=�pwp���7�3��qYKؐ{��蚺�fd����	TF{��	𼥊����Qg��
M�t�;s�+�����8��J�D�ꌋ�)ez�� jU����k�"�weu?x����g+�a߄Z�j1p�a(����8D�����<���F��y~ݑ)��v�~�wЅ$c�/��gaN��5����]���\qPM$T�&����r�O�2="�$������sr��N1��y:��Pv	6��JۥJD�ml5;���~o�~�����A���IQ����ޞLᆷ��6n+aw;�`D��o2�лQ����S�x$�g�2��$Mh�j��ڒ��a'#�$�6)r��L���t9��/1r��G7��<��[]����^���l�cD5���%������r�u� Ys��A�qMP�/rV�\Hmt��o>�<a��z�����%����*���ڿS�q� �{��v%<w���M�]�H����#B��U��Ǿ��v��`�S\y�x����؄�͓�s��r���V��L�է�]��s�v%㛰�-���7�u��@v�T�c'B�9d����.F�{nI:iXU��ޖ��h�r7�8�����涟fq�5l�u�T=�T�V��ѓ��l�6ǈa��L^��3L�s׀�5Rl�V�]:}��� m�*&H�����4۞�2{�k����s7�]��A�:����ó-�ݽ�A<�`We'���F1�q�2�����SX.��f-L�f��v��A�Y��h��}�z��氵������Ǩ��x��8�r	C�ɨ��ޱ"���<f��v���㎮��j�.X��e~����xɑ�
���G�W{ʸ�sv��	���ڜ��N�*z�߬�Ì��7��{es�F��2ħ����hl�Y�L�Iف����{�mr��h��.���j�c����&��ZJ�ܺ���יO��1\9�(��9O�?Q����c-M�9����T
�?
ŉ<
{|/��@mݼ%��H� �qIZ0�\����7V�Y�~=�t1����jȡr�#���B�Ѝ�:Ki�n�YD�����k�y�M��\("�WäBP:؈|g�RVJ�ɒIT��(�<3�ų �e"i�]��*\��<u��\Z7g��T���*�G)z�كՄ?u=�m�v������6�&�T�p���gs�׎'�Ek��o��7�43���k��^$X�x�#�﫤0Y�qܭ��EDk�ڦ��=y��D�z���oI+��WI��f�7��N�d�Iv��9�V����rd��6�ǒ�(��T�2.FR}��;dm����Y�ξ�r�����|#X���F�����>�S�Lt��!��^�q��|���_ӬO��t��C��i��E[��]��J��z���z�xx��q�dh��g��3m�[n�uL�hv��%M��%�W�J��xo�u"�^�vAZ���F��i��:nwQ�f@��ˈ��*T��	�mu�Js���s�w�0T�x*u�J����0�K�mI�}����>�)���QV�>_P���d����}؏��7��Gtk�1�%���)���[��zC�C�	P0#�^x��n���O�Qe��◸�/��x�A�Jv)�;PA�
�~Itg���nb��ٗӋs���whsĮ*�!ȴ����b��5X� �P�&˲w��כ������}�333Eb�)!<��^*�PH�{6��2�i��p��3}̯$�4���sd�\d�(,�AM,���'s'�4��S馦{�Ү�Kl�Eo��ƈW>��7��{Z5��I#����U�	��Ik���V�>��x��'B�0���;KjF���j�j��l�j��-�39�YMS���V4��E�B���2�T��g�`Ea��c�6j(����ٽ��Om�$���8d��}�A�!l�8i�G���#��]}y<�J�'�2`Ǚ4m��o&�K}�JP	�Չ�ײgCG�����ø2d����?'���k���R{���{z�s
�\�n/���y���/V�T��v�R��Z��a�1&�:��������J��ͧG�&IyĮ�X�ql�(���3<Ի^����T���-�[X9�ݽk\��Zѳ��H��䞉���̊��Ê�PK�v;���j���܉T:����j��\�
���鍝��U$�ɣ�H��+�}����hnq#^7���5P�$f;�p��7��j��W¹�Y���5�V�v�j������0@�y���[ v�G�s�Sӣ��k�2G촂-�>�Oȟ��;�N"��s_�e;b/�%�0�4�v�,���+��� ���}3[�%����!�/#��UF��2��yu{уD���j_�.���zV)A�o��~�&�(����%�Y�����hU�=�u����8H�� �*Ȑ����庣��imk�y��r5;��kEc�U<�w��#"�*�m��A�)��˧@��TV����bv�t��� �?hF�lQ�[��w4�̄k�X�BC�ǹ ����f	�n�w\�d,���1o�<�����j<��2I��-Fs�2���m;��p�m�5G�h[F�+�"�>�ِ����u�
�ǡO"�ԃX��؁9�Q/ө�p7�<��-Z4#Kq
�:;;�J(�8֑�{]��ڥ {2zi暇���d���|ɆJ�a��ˋ�=�65S(J�QS�$� �kr�`�"�$��_��� ��t����"�G_n���%mҥ)�5���j������ގ�f�}_m�p�A$� ���qGG�Ԛ��u�W��J���+yߦG��4wA�H�Y���J�O�O��A�]>���g��*�.�r���K���Ǳ�
����J��﹐��0G�f'Ϫ�b}%h3�|p�\����6�vU�R�{�̒kT�{Φ�(!� 0��э<�)G�[��P���.ok1T�P}���=Ԕ���6z��}����
_��_~�NL�9�������)�PZ��'����$wF��z�l1�Cp,}^ȷޤ�^�S��/��zf�r����ԫ�%��]��a���rr���u�E���>��xH��g\]�J5��;�yU��]�׎���1���Wa�{{ZA9:���r�n�d)v�fT�X�V�)��n�P2,��@�F+�\U-�O��n9�g7Ǣv�z6�cW�P�#mq�d��%��]:m�e�1�*o3�fF��hv��:�x4�2��p���y7�H�'ė��;���������c�������r:#�YjKbj{F�G�	 Wmx��7��[sM�7���`�������x�g��!(w%����дd0Q��>f���0�ݨ� d+�!.�������߿V��޸%F��,����X�m�Ӭ�؞0`��o$�Z2�B�v�@��3V���ȷ�-ϴ h,���j��ww2d��ݡ�#���7 �z�O%CВ��*�Y���5�^(]�ٕ�i�v ���2D#}�"@�7>.�yl�$��U\a�r[]j<6z���F3��[S�G��Eqm��r�TBc�Op�� 'w�V׃��/?��j�[���Lj�΃������z�c������{���w������z�^�W����}k
�E�k18�6cO��4F��v
�9+�	̠��3X��i��No���t8n���ۙ��z�V|�tZ;�MK;Y��cn`��6�s�w����'m�OF*�:�*I y�m&�V��]�I�:���#DP�RWtL�=��Ɨm�м�ڟR�m,W�A����$��[,
��1z&b�r5Ķ�S�yfY�d��FMΩ�+�H���ŷ���������͑����,V�Q�;�L�w�̩sGu&EQ�1�*pc�=���(�%}ęg�����f���ڂ�»�K{����!챩E��{X1�vq�ԣ9}�r��x�~!��Ƞ��BE�Ǹ=�Eu��"�M��� 	�c���Ԅj�2��{��)4b߰�m�'�3	�b���u�E����,�S��3���zM���kT���ͮ�On��m���E� �L��Y�f�p�+�\�"�(�r���n�l�J��O�vn�ޖ�9��ZJ�S��D����q��+(^4�m�2t�&^�����v�;#D0x������3����i�q�^XkX3Z|%�gSj�ڕ�"���c�h���({�V�C�=)��3|&�Fz
�ŏ^˺�J�:\쾕�iE՛o�R��l�!V-���(��\�)L�k�������i�T�T��yͤn�=F��!��r9i�)�\VJbJ�H.��xԸ	o��E��<'_W"�>�bV ۈ�4�� B������M��zf֮���.�8�t�5��n�Q�];k����/_#MA�J��ώ�\�@;-�1{ �U���'��:���*a�Zї3P�ϔ7[�Nu*3���@nm�o�ڳ�
���u�5v�q-�/IX��ҥ^ܨQ�v���
�,>KlB�޾�G�e-;8l�d�tQ-�*�C�-ډ��8"�V���}��Uu[�m��'Z��j�Vn��==7�0�>�ҩ�/;��I��i9Q8���tS�C��E�v���P4�#�C�&a�En�x%ge]�(�:�q�)���wq�.��H�Jxq6������i��s�p� ��s�8�
58��n�e��x_F9=���u��,g:=LT���B���������T���c���˖�S�!�ύ�`�F�g)�/�:u
��`iJ}f��G:}WY%8^JZp�. ��J�����l���5֙v
��U�������nwp�2�)]�LI\�\.Á+� ��/x�*Ww;]e�V��|[0q�I�4S���6en	�YUl�k1̉�PoiJ|��1Ö�t]S��>��_���p�ޢ�J��u�����b�����`��o����V�ڡ�Sk{G(��;0�x}��	�14Q�j��0L�%lk-�
\��R���xf�;�ō��o����i+N��(v�P�-�()�
P�C@蠠hh
J)v�T4���Um�l�:u�c@PKat	N�ZR��i�I�446ɤ(A����4�ց�����4(i�l4�hSN�ih�Bh].��
V����(j����4i��ii)J�5�ґR��q+taДRP���P4%%R�SMR��$@44�PP)l.���bi����Jh
Z��)�(~�}w�{<��P0�"���Q��j����|ԮҬ�*!1��#5����\�܊��W74(ۀ�ճ2'��|��Tp=�.p��k��]�.�P���22o�QȔa��_�18"!�PE2�*Fm)$���Tn#]x4I+j�n��}X`ɱ*�ITs�= ��[�"H�r1g[`0�� ?��(��iic0�Y|#e����9(�bU�'vA��0�t7�����>����Hl�y���!�3̙�GZ���]��
�qsc�E���^��RAQ�{3{7s�m�	Po)�knH�4�Z;װo*�9v��S�a:6�1��w{��}ǥ�s�1���c=�B�}�9!7�^������br�ɓ���������j~3�Ϯ��0ά؍Ĩn���g�BJj��:բ�{2P���g�Z;)ا��gp�t?$���&�wnpm�esdw�zx<���fnG=+0r-����b��,��D~3��\��}���s��W�FO�'���I$q��St�a�fn\��606woN��0�!�c�w3�z�.2u��AM($�-=�^>�mVf'��J��s}��;�aݱA|)�g�N,[֕Jh+���U�N��I��j�׍�p9;���ըvN ��;@uN�Z�=y�� �%�*@T���������<�%r�*vZ��b�'z��m��J�ʹ]��c��[���"�4�C]����w�85�PW";��X��ji2������!�[;�=5裍Ѽۙ��Tq[��[<��"�Њ��� v.�Ԍ9�����Zr� �vi���V�)�
J@�}���v[��[���{)�h�C28�C�bU��wC��_Go]��l�'�Q8d6cǶ��!p��C����ΛZ�J��	"�;o�=Z��irM�kZ���]��|,h3:%����U5*��{	�}��1C��t��v)�\��
�%��v< ]����13SD�14�������^�a��q�EW�U��Ѭ��G���`����sP�]ݳ��O��8�p�!�pQ�GvH�4��S�j�Ak�f�K9��]��/ٵ�\��,���A�=�a�a�t�E���a�ӑ�������ott�uo�eW�c��Lt��g�A�t3��q�U���O�i���W{��G��f�d�����Q������rm��t^@�t`�ة�$�a��,c�5+�����t���L�YԹ���v4��{��	U�$r��� ���6���{]("���]�l�P�%����5���7܏�ť2��7����=V�W�c���߾r�g��'���8Ē��2:���n� �fC(��0�+��"G�[�/��<�������w�
oO4{�Z��ni�� 2�����xlFMv�D��fga#�����	p����P\me�f��v����{:���U�z	G��z�M��#RY@E�荪��q)��3��F��>��� ���s#8A\X��"գ^�]t�����b;�۷�s��x:N�zM<����4�&����PE���Yg�<��tuwu�n�9�ϛ�F��TQR䚠�kr�u�ȼ(�(U�0�����:Z���O�6؈����$G$�n�)6v�j�7r�!�Qh���Y���/n��G��6Ԫ�/ u�T�\l6�!o>�3oవ0��8�;W;�e��)�R�tH���=ؔ�����}ߘ�Y�b��.��J�m�	L��}"V� �U���'��G�7,���KU����yIn�tr��c8:Nu`�
Z]1��E�N�@�=��}���d3}J�%�Veo<il�\;3�ЈL����l����`�r�K4v��Ǘ ��F����2��!��6��ْ�� 쭧�Q��zz��/[_����f�nɽ��l$���#;U_;k�h��wZ���wܭ��p�9��u+򮃴6GSto�G�"�M=��;]�vi��"9�Qݟm���HOӕ�2Gtl���`��,����ӽ�ͤh� �P�֫ь�F`����@�"}Ŏ�bz��g��v��3���U|�̻P�E�<*4#/��љm��1B����ݫ���y�f댃*-��� _4!��ϮW<��27�1 ��bZ^coB�i�}�t���V	��ה����8;���>����p�7TL�t���f�����`NҖ����]m������:����M��Yyo�	�;����]�	x��!V{y%^�eW�}���s"����̇�q��<����6`z��8�&Wo�M�N�sK�O!^8���q�S0@��J������-�~Ng�u���LE�>!n��e�m_\�T��f�{f�����dZ�l�w�L�=�"�"�KS�a�6�v��X����m����,��:O�J�Ɖ�����?S�|��INbغ[�S�Ѝ OO��IU �wj�4��/2���<Y�5�H�h
�!nQ���78��J�J��"s;��1��g��cIl��5 �y>k�[N��[S)��۳�(!�
l�Q���y���j�y������_�l)�;pY"5n�Alu�ao3<�⫚8ǆ{!ώ�8��`�u�F`x�l0����fF����n�t�<n���u�SGfҥ�k�/��ē�>6���nw����O5K�p�]����1�$���d�]2g���丢f �O�"�)>��������9Y�:����8<�5�'۝J�-����sk��<�������$��y¦U�3��A}�9!d���>�G��M�󩕃����:�*�|��<aHZ/�u}vt:}�gV{�؍ѧ�膡�;<������n@ْd���x�T�-����s�`���<<�����ݗݶ�)L��(j�>���.�Sr�l�G3E{~�Boq��Լ@���6c[�Xvsn��G⡼ҞT�v7��p�����H����teK�3���k��MN�:$�1�[��(�ط��g@�!0�M��U��k-S,髬~��1�yX@�qw\wy��Ee-ysc%��:;Gn��ô$�s�y�����+�=�������-�GZFm�L���y�cD�=��o{�ꏜ�s��w2�ѡ:�Y^E>��*���n�Q�m�VՖ�O9��x#f�υ	��7!d��j�/kF�Q0��x�X�'f�jl§ѐ{_�srgsۙBU���O���EH�nظ+�upy���/AF��Y���U"-%Tn]:���dyՆ�}.���Y	��?ow��;�μ��U��Y	�I_��m� �\M��n�B���ų�-���:,�#�:����Z��ir��ֶH�#����x��¯&s7�Ua���Ǆ�p*�l��t��v)�Z��Iw.�7�����DI{¥(��2o�(c[�^$���ڌ.�'Y.Ȩ�� Ò\��j]�ۋ��=�q�.gԟ1���+����+�=����;�O �=Ε�sxmvA�g���j����n����.�u�%�S4[�3��|�3��=����
�=s����eg_����I��U�h�0r�J�郷Xy��;_VV�>���/��x���8q�C6|ހ��كpңO+#
�V�����[e��$��Ux�ǻhf�m�`�0๻}e�NZ��B���f�.M��rF��r|3N��3���d��;fGPcK
�z�~�o�r~����!���$3;3�֟F����t,����F�q�Kw�ޕ��I��/� 31p�y��ꊿjC?b}VL���!�w$�#O4r�LA�jو�UV������r�A�=�5WU��	׮��%QC�Xs�.�Z�xM�����n� ������OA(��OP���#"�%w�y�=����$�<u��˷S�~=�=�f�=p*%̌,�A]�4��-Z8X!a�h�m�|y��i�:�I�G�נ�=�=4�� y9>>�I��Zya�v�w�C�y���7���@'C�Xs$v��wr�^�� �:�W#b���f�|�G���]�L,/Xq`�Ys����{���7�p�В��:��{I/+v��';�{�4]�jg@���C���g�Kۅf�K_Io^M�6gdP#+�^�6��.�\[����i�庞̛J��T���{�Zs���Y8�Ц/�)�n��7a#a�$�7J�$|~��U�̉w>�7F?ޓ,�U�~׃FPt�}lm�Ta~�+L-�R���	���pK����>�Rj�u���A	e��.�]��WbUG@�3l�C�eɓ-���:@�<{��u!C�l��e�սCfJ�fΙM�ld�h����yö"M�*���4n���`�l��a����Ƭ�׮�=�%^��淧qPW����Y!v��_�Jy��;z[�j��[����A�l���طYn.�W5�R��N�HO�ㆲ��c�6}�p���-�i�W���}�n����5L抌�?*�h��ŎH&+�׽[mW6�q���]A��k����Ψߣ/�%LK�9+*��>Z�W��z���-��I+���m���
�Ύi�V�+��$w`���_��qy`��T��[V�t�${�Ou�9�^�5�y�j1ҘgVvv�n���xc�ҲJ�����l�K4��Ҳ{��R�sc����:��s1d�"��$�x��\�*1�:*<��_3�b<��zJvj�n����;P�^�^N,�6�9�C�'dDH�ɦ�Ԏ�x�g���R2h����D�qӗ[��>l�����v�+�!.Ƽ����,�2�Y�`Tz��cr;��$�4��70����A]HϨ����+n�j��+z�c1�u�؛Uz6WC�y�m,Sr�XD�.�܂<���_�%L%��.��X���;k���6��g�$�6Dj�b/m��t����%<�z!�[Y����d��Na�M���k�3�<.rou	!G���8���|�Tl�5�ta����4���Rnχu��m�0�����@�����K��O����@�#pek�5�="�����o���eX�+d���Y ��e��ͭ�K���&�D��>6�M0q�����cw��C�ڛb0$]��.�Q��v���n���ܽ	���:�N�,ĻA��tV�޺��0��QdE��Pi��}���7�Q�r����� ��5�:	��9��'���&���6�s�:���2Ȕ,�ݏCV�5���ނ�'��ٷP���4㾭����|h�����޿lʞ��y-�MB����q��l9�{�3�6���+�	�q��knH��T����o)ʘ��F٭�FD���������6h�p�-�o$,�n��G���ڡ3�L_/B�$p�X�6d���+�Ch�g>сxVkލģwF�m1��:�<:�V��B)! ��n�*�)�� �v��=�a�&9�nO�F)�[gsљd<��4U�#�h�>T6l�}rԄ�T��|Ւc��A����U�B%J���Ԑ�+�2	���n��$6�w8��V��w�'Y���z
�-��s!M�Qq��W���
O��ߵ��� C�vdl����F�й�頁��s�j�M���s�n��(u�7cF����Zzy��N�̞V�"��@)���T���}����{|G�����{���w���������������&\k$��o�YY_:�=:��٬���}g�o�	�
��r�z�W3�cU��s���Ww�]c�}�=*s��5�s�b��s3$��9xM�r Ym���E!;�K�Xq̕������*c9�Vg`��]��z9��!�\Uk��q1V:�$���5eLc:��g]��u�0h�2��h+PS�"�+,�J�ä?��8<�:����c�w����Ge����/t'�c�4��+���ѰG-s.Wa��܀ˋ;nm*=�ո)et����]�-���Q�Vf������e�	Q��D�L�Y��C��wz�kk!LwgXr�H�zc�w��=�o�f%B���u�HN�Gxn���T�l3���Ë�X�*Z�v^�@�wr�N|(�j�7�U�/��Ҽ�Y��^�x�&+���B��G�P�n�z9>T�u�Q�;���r�h�'�9��ZM��˽t�<�52�8o��΢��ξ��O5(�*�`)w�R����ƛ[o��U����s
Y��!i 7�V���#Gm�W�f�.�C�p�֊��ɍe�c�I�}9�Y�aK��U`�ȴZ��%:��l�n����ྴ̽��V�(9�6�I�W0�#*�x�Nȟd4�jR�q���L�9��a���*_5��r�i��	Fֶh�Y����4�ǧa�hc�>�D0��v󺽡�#�Y�ysZ�zU�;3o\4�jspa���'�Yw;1��Q�5��p��JpX��f%36'���xɂ�������z�͍�*<[�2�r����J�-��ó������.���M���X��&D���r����b�R�s��0 ���L���l�1�QuX)�u�Yo8����9��z�}�ȁwqÇA�]�m\�������#5w�X���D�tU������'�_aZ����]�Y�X���hK%p]��.�}ܯ�w����3B*�N��]�"�NV+9��J��{+��<vVg=�5˨Y��MA�@,�_ܩu��ǆ�;�Dt���ai�n�!�
�U�����+����u�R���I@��]P�1����Ov�u-ƺ]�ֽp�T����N���}����)�;�w7F��N�����i���2Cj���3ym*׷��������nk	n%���KR��gd
�o���Q8ܹ�g�Ե���9ջu�����fP�̦�Ja��t�<�8l�c�	�IK���S�gm��tĻY=��"!Q�1�<"�u3�2�Z��靟 8l�3s�[:�W�`Y0EܤS��P�E������X����c|&m�(�U�b竐�5C��;���}o_VD�
h>��n��eP&�:ށfd�z�ؗ�+ƹW:�Ҍ�|�S��c��zok(�
��zNq�[:�P�ֆ)���Y6'�{{7Ws7Ԋ�g��	��
SF$)4!�(*�������1T��DhhGA%R�EPP�44�T�BRPLP�&�4�%[)�)(�Zh)(hMihB�
(���J�ZP]�Z6�BU��QIIN����4AT��c&��)�
���	�JF'�4%�5KD@PP8�M1SHP45l�h�)JF���(��61T4P�t`tj� �`�(����tib��I�
��"���x�o>����͟����8��5��x�um���^V;�Y��Q�o��]�î�*u������Q��a��N�A�����ss��C�_��߸�J�J�j�]:�b���Uw|j��r�z�q_e	�e��n�)hn\F��	���p��a�m��fC�S��Nn`E��͞ʭ���7�ƙA����%Ei����Z�����Nˍ�ٺ缨���m��n3�r9Lt�tLv�3\��¹ G����'1�+����֧^�N>\�]���1@C��ȍ�]N�9T$��z��EִOYɼ˾�����U#/i��!�o@pQ~���ii����K�Ǽ0t��H��V�wQ�Ô2F�m�7;๻p�G<��;u��h],樽�'	��}�^��d>;fGPc�g��d��/\c�a���{j'hXi�z]�w���z8N�q�KA�^��/zu��
&�m���x4}��Ń��T�U�{�3,���D��#�y��ѝ�������Cs�`��I���|�L���U�8.�K���rXzY
�1vv�!:kB�'Y��Ր���!#:Tv*�Kѩ���Xdߪ⬬ǫ\��P�OeM��vV4yNO�\�o[����;H�B�� �ښ��-�x��/�����<�1yE��h��B�Y�%�W�^����#�vGVTh��J�y��1[��j�ӂ+(ϵ[��g�^�P��iҹ�:X��vq1����}��Cgs��;��R�8�@���%��g+�a߃1�3q��,+r��w
��ٔ��,�VJ<(��yU�c�4�&���r�a�+3d�\�{��a��#�G��F�l���I].))I�{��N�r�e�U���5�G��DffXR���o�v6�Ht$���>�V�ȫ5.��������Z[uԎ� �2 t�D�6̮��:�eq�|n�n}��o����h���ÎW�����+$?κ��g�v%G9�V�.��[eBӜ̷t{6N^F�"W'�[��K�l��G�V��*8��n�b��2��"#���x#x�W��%��HU�>���������՚�9���k�Y��>Xsqѩ[�˩ںF�7�>m��.xӉ�B�h,�&U�k	�+��=�ɍ�	��^f�xz"�֭�;�y�ڥ��Ԯ\�v�N��!��s1d���X�i�C-�������,�n��>���[�.������z��f�;�`��m��c'G^�5�q/C�ףVu��yB��mq�aWA�#���*�"7f��/y�H��*�=��c��rF�*��h'��/xt7�{.�9C;�Ze��J�=U���C
��C�_Tc%9� m�4L�#���x�{Lΐ�����ǻ��
��+~���
�F^#c�ve�E2�k5�v�mg!ݝy\:�A<�q/�^w���p��,ۿ�*7u���^Z�F�g5a��&"v�~�	"���#+K�M�kA�x��A+<.u���i�l«�sgz(���닐0�[�@WQ��v5�,��9�h�j�ѓ}�75Gi�0���'�}zW�"i
�o$�ѕP���bٹc����c�n��ut�qj���YhW�r�ՄO�HnAO�B4O%@�x ����\������3ų3;H|��e1�j��Dc�~�b6��y�X�̥Wu-�)�r��<�u�Ƒ*�*�j<k��S�S�(n�V�瘬I{U8i`[�.�p���#�����҈�|�zB�1m@~�yu�./9b�7�w�!�G؉�����&��g���pv˾�+\1����ѧ�/n�O�C ��i�W���oD�tg�$����]�W���*��-�[,'y��XW:Ȩ��{M�װ��d�H��T������?O�[�Aۂ�Y������_i�8�F��)��xO QZ�GU��x��[�����aD�wid�+��p�c!�Y�[6��V�qE�^�N�]&����(��S�چ�5��Q�zcgUtʞ���,%�
&�����t\w��h�v�[�#Ɠ����q���n`�J�����8ٷ��;�]Ǯjt���Pd-���=��4s9�ټ��#��-��gR?�w_����W���=�k޸�}t��ϫ���0"ά��a���i���a>ڵ�\,��t�'�:�bN�b��?�O3ੰ��EaW��ۦo�Hfy*]^ټ�~�qwD>���By��S�K�`=���iR%�Qb]�Y���)^WVTN3ȰU������+V�2�v_�#�̔9f��G��9�`g�R�fm��OL�F�>;�>o�z���<�Z�̵Qkp%O��;��ir̙wz�cw{��)r�<���F+�MuNW�}�M+�/"�R��ȭ�j�я�D�r��{q�JAW d�I#mؙ�f��Q�1��`���;]Oy-��qA\z�P�r�}�����9!�H��"ZQzi��:,���9��VG�G�$\Ӛ5y1��0x@հ�=����g�m�n���w;Y�[z�r�ȣ*��v�}��w��/��UxF�c���MWSjy�+xѬ/�ް{�Kq&���I$���q�u#K�@"��括��f{��l�Wȳ��!�lm23{��	!�x�ɐO.�pϛ1�6��k'E�*]�k�m�	
��!��;i�դ��8�����~v���>W�ܐ���} K-�<��B���A��gMOW��rך�*0������b�7��w8�"<k�e���<��:�1���M��O�r'=�+����;�}���#R2���0#4��pQ~��W�כּ�+3p�x�*�����U�Ճu�H��e��`�#s&���M>����)�Y�?�ܮ#f�O��x�ʯ)�oA��d֭�R»4�#�-��fZ��bT��q�ݴvUޣ��b�����/�6lyC�{������%��m�RV�e�g��
p���{�����{����r�_�m������L���t.����� �@����k���*8���0gv̎�ǝ�f�E�mdL�]��^&m����#�hЋH��t����#y�ω-E���e�R�c7z^M��z
 {xJ|jѽәd9�����d�����NDQ�_���]6-�F��
1�E�nlfb�GU.H:t$[�X6_7P}�����op�YFF�u��PI���(��ݎƥs��]vx�ݷ�Ӈ٤�_M�Iv1=q�s8Y�W/�SRy������T���lƠv�������W�J3G�נ�
�]�i昵W/rݩ�=yݏ�S��$:4k�6�h�[!��m�zR���rMA��8�^�S]����ɉ�[�u���(�B�!��G�؈���Q�I��Og����X��;��|����*���֥�=��v䋥[�2�U��z���MY��O�c���¹�s���ѯ<uF���]�r���P�B^2�޹H�k���̖*�V�c�ӊ��π��c�#�{�j�J���n�4�Aj��r��ds����3x���j�R3At��ݣ���Y8�O8ڢ�eW)�l��ݳW��������p�\ VK�\�u����,f��9�u�����Ju�(W)j]�K�e7)��`�V��}�r]����7J6+��v��͓��w8%Fw)*�d�����axm�9��c2	G ��cu��m?d��;�3�0���ԕ�Y�5[@��Vt�6GSt�l�]�2q�FNv:��W�.��l�F65Ü��*�҈]���\��� �׻��0��Q���Q�+�&|Ah���f͵Ɓ2E�hb�jFgf�h���骻��g�޶Ab<;n�s�����<*5x����z�ɉ6U��x|�����h�3�	/������� ^B`=$����g���"���糟r�c٘Hy��*"t�i��#���;��G�ua���T����a�eh(-R.�n�L\�,]���b�&m���H�i�eg��{�"e�d<�ݫٜ�Ƌ�A�tJd8��toG�0�x[kV�Z�|�9.��n'�Vr3��>�V��5�J)��9��rGv��*�|�|�G��R��?P�3bc�.'�Y�.������.Ƴ��X�MB��m*;^S���4z*���0q�Q�%ё��B�4��eT.���N��|�	 [���o�5m���++��.]$F�"{Kr
OB;939y.z�Gtݖ����X�n�mU���&�]x�2a(�[|k;z�^��A���m�;#׽�0r�2I*����ө���P��'���U��0)��~�˨���;F�wZ���Gl���"�Bб���_K�aNe(ʺTE�]�Y[x��v3�z�BJV4q<QZ��up(�E�>:ێvn�"�R�����/0��9
2 ����Y;�^'3�h�=d�D�`6��I-��|�̯���_{�_��FΪ2����K��jW���F�b��Oy�[�mN�q�st�do�r8Ƭ��0�۽��x����3��6�:7��{L�7�V��gQy�t�[*Y�3@Ux�dt�`�AB�1Ȭ�t�y�|���ѯ�o�v�r�����67�J���rB	z���#g*J8u�����a��Εܥ��y��UHS�F�Sg�
	ont�9;���r��9D�O�؎�� o3��Gy4�22Bŭw����f��c>)������?�c����G]M�ŏ�D�Ja��yy�DC��K�rl����H�'�n���O��Z`�z)λ
� �d��Z���b:Ē/��]7�o��{��,
�'܋Ee%�Og�wr��6Fܜ�OGh�ɹ�0��8�bN�Dעzz��d�I	��G���x�#3w#|��St�e� .���|ɐ��#x��*�z�4)�d�{����������g{�Q��4�E*�B:��Ո6�p��v�A��.�ot����ATR�:F����W�V�j��LE	1C6:9�g^!��u;Y��j:�G��6�h7A<T��J��.���U��|�Cj�̛�;�|0h���L���<;�$9q-�I��	½���ў�,��kѡ˺���8W~�V����Z�M��
L�{bȶ���~�[�tB�z�ɱ��u�C�Z����Yޘ. �}j�.��.�q��I	�FfiM34�g��s]B+nj��p-h�$�ލ�����X����i���������l�m�6 ۅ��t��.V}F7&��ƽ��E^�ǉ֣�S���an��r7�=	�g�������~`^����O��{ s ��,Eg����ӯ݃���3���tT�Out�#y��<�V�U=�čȃLt�wLFd^K�w��7�a��W�6m�雾9wF�H��4:
�e�hOI����&j��}���ܸR�����~��llڍe��M��l����&:A�3����f��r}��>�SH�i�C\3�uJVs{<�w+}3[L�u�������舘�7q�4��m�$(����Rjѱ�c2�y<H��(�Μj؉j�Z��~����mP�3ᡅ��v�Dշ��fw�2(p�
���^������O���	<&��m�7s߇��tn��z��������ݲ9 U�� �"����̿�PO��";���z��v!(�00,��̫0,ȳ
�B� �2,ʳ
̋2,�3�@��2��3(�2�ȳ�L�2�ȳ�0,��3"�!̫0,ȳ�2�³�+!̋2���"�2,��*̃L�0�ȳ̣02,��(� C"̣0,�ʳ�0,�����3 *�2,��(̋2,�10,ȳ̫2�³
̫2���=�{� =2,�3*̋0,ʳ̋0�Ȱ�0,����@��C*fDH�� �� ��ʠ��Ȉ���@�@@� �Q �D �D � �z��C� !� !� !� !�(� �@ �  �UV@�� ª�*� ��2��� ʪ�*�n��*�2�2��� ʪ�  L(�̋2�:2�ȳ̫2�ȳ (̫���Y�fU�`Y�f�VeY�aӁf &�V`Y�	�f�d�o�`��x���@Q�EQ&D&O��7���<���=M�C�o���1�׼�6�/��m�~�������=s�|��o��@_�~���������xU|{H U���?�>H�����S�C�~�?�( ��ӏ�����:Iw�y����� �О����>��,W����,B�B���1(D�!2 �H� �@��ȠJ���  (H �*�#
�� �� �����*�$ �)*�*� � R�!Q��`����_Gޟ�(�"�"-@+B�~�� ���Ͽ������ð>��'��� *���?��v����O���	���~ �v;���w?C�
 *��ԟ���ߡ=H��( ��!���?hz��'c�PW��?��H�� 3�~��������'�`����};�c�=�?a��v o������?o� U��}��y��������~o^����I���?�y� *�����3��pPW����}|��)?��������?~�~��{z�=z	<���@^��/��L��`>�0t��x�'�/�T�G�����
�+����Ͽ���>�����(+$�k&��� }��0
 ��d��HOϟ��l2M5(�J٪��lX�ق�l�i��H6�͔$���[4����j�Zm�%RUm�[�gl�cQB�T���*+m$�H�KZVѵRʛ2--�P�pm��ԩC!mZ�ѳ��[mG��l�F�X�&���V�e�*m��d�X�͡�j�SX�)��VD���P��Z҄�k#UiH�U���a(�Y����1V���iF��KCl-�e��k6�f�́���ݬ�#E��єRժZ2�-���,�[Sme�x  �s^kO�uz��:��\��u]�7n��ޕ{��i�^��5���׮��*�j�4=��t��뻭��U׽��k:ݵ9u������t��y�v�kW�@���h�-�SYm�lV�Ӂ_   ءBC����h�;�p�Q�͛Y([2>|{}hP�4(t4=�I�СB��p:���U�;���n��k]�ݔ�������w����n�Ji�.�w{�==Sݻ��s�k�=�����[@���[mbK���  ;�κ}=j�+����櫽�R�p;�޽�(C,�[ӥomokT�S��G�ޯ]�w���V��u���wy��{2�v�����ڏqw��:�g��m�6��:�v�����   �'��A��q��z�ݚ=kp��{�z[U{q��"�3V�[�^���v�s�׶��:��ٜ����ev��C�U���At�êY�13M���+u����K4�   7=U�V��5�WZ[�p P�F��gY��3� �2�b�o��(�z�8
�rˉPi[�mh�5m��-��4�m��  ;��]V���᪣��]N����0��l��������B@G%�v��k^�K�Ir����U���El���b(�m���m���+I�  {;QGۢ�ѐ}Á��pv Pɛ�p(u������X���dzz�À ���
z u=ƀ Ԯj534�SZ6&�kRV��� ǀ �w�  >�z��z�����r�= .���n�נa� {w��zz �bf�� y���@zk�Z1[f����ٕafYS� �J}  u����@uX ��Þ�� �z�Ǡ:zx1��e0 �<ޮ ��L�@)�^�  ���RIV��*���  ,��� 
��  w#  kѽ�0 
�=�([���= h{�q�� +�S�  W�� ��` t���R�(���1JR�� A�)���� 4 E?i)Q@ h �� �#5  OT���UI� 5??���6�~�~����z���m>2ʽy�6��__^��]�)�Ю[�_���{��o{~�?=����խ����������j����m�km�M�ڵ�Z�[mm~��?�*�o����^��SQD�bV�3FV
 ���#��}J��5nڧZ����h���:�4����旳UJa�eU�{l��0����l�(b}���X��Ct5��
��k��D	%�11��-q-YJ��s1�x�eָ��H�C�c�F�\���JȢ
��J�X�(�뺽Y|l�]m��[���(������4�%P���K�W�@.�*� �r�T�1<vu���ߒù2Ĕ���jN�9E�)@	�6�`�&Y�b�-!o��<\��:���4h7�M��WQZٍ븒���fY�x�ҭ�H���ʴ��Faq��fJ�^ږcʺ�!R;��Xs@�z��(,27Vw3yKeaVjv�2ыv�W���]���	�NKa"��S�{kT���M�Z��ir�X�����^�'Uڵp�ܬ�YG��҃z�F�.�Z!to6S�U��4HڵsfB���JͶ��{Zv Y�L�6\rb%6���(T�D�$������N!������$�VJF�f�.֝��t�b*$2�Kc�i����bؘ4 ʔ�҅�m� �7,��:!��5j�e^�G$͎�����,]7�PQd��I�(	�*��ҖX9a���7M����Y5��k`��F�P�)B��E��t��V�Cך��VOY��k@��N,Sn��ݘ�8h^��b��4Uȋ����@��+)�C�,y�k&��":CZu �m��n'.�ݠ�#@+���:]*�F�V���h�J/~���]ʺp�
V0��w�@E�N�ܨ~���oV+�8��9�͜��=���7�R�-l�Խ�A�
�ޛ��R��$�rf^| ŃS���۬�4ڋ]��aF��[zpXv�D�l�$3��D��j��'h*�=�-Q��R����*���Y(�)V˳��[w���R��K�d�j$��>���7WE2/v7��
ූ,�`f�w4GCͩy�a�\��U� ��*�0m�v}2�����d��� X�b��ke�?ZB�*�nvWi�w�@t%��i����ah��&��ga��{�j����bM���OHR�YG�W ������+`��Ӓ\ܼ�v�F�Z��ch�qM"��{XL�^,�`/�VJ��,�\܎�b�Lf�WN�7�D���gw.�ݧ��b����RD��:u"&\㭩M�Wp���3��
�4H��"�S�iSG�>��[7m,�ZVb� �cl`��xf5�G(;�5:Е@("K�(��Y8��2B�0lI��F)-�P�n�'	G.+v���I�g8�ͫ��R�g�2K[t��]!H��v%�#ldm��Y�C��r*R�4+��rf���;���=!��aP[�*�^�,X��Y(�R�D�F*��ܼY����f�������)
����(�͹�N\��3eT��H�Ɠ�W�L�f���L3Z�CZj�E�0K�I
�)P�E�Ehwf��H�v]gq�o�H!Yt\z۠�θR��n`�������-b;��摸N�=�tE)�`�5r�j�+��]�&��R��b
r:U����P�����&i
���Y�eh���%a5Rj�0�j��G$�l�T�>j�/���;�im�c�Ye�wʂpd۽NZ�+Te��2�鋱��Cpcyr��4���+��-�f�;��9�����T�����ZX�̂�i��V	���\�����d!(�-�,݆�,�͈ԤiS�R�:d�C`��0ޕq��� ώV�XF� ��Y���_rX+(Ӯ���|��5��˲�Ӓ�2�F25�,8	:+(I�+Y���ݜ���
[&R{B��\��˗[�5� �y�ivn��j�c�w��jKyr�2��l�ʥ����h�n���*�̖F�vS��q��6�e����5-A�P6�������en<2*�V����6�U�z{�*nU�3H��u�}kF�enĤ#^,�^�0ʨʄ#y���-�v4H���-�j!6�#u�\����le�G�Y�Y�$*�c`�V�Kx��0˔��`f��0v���  �%b���WP[se1� �Ce7w 7�Ld���ٹ����8f�j��l;�L7��bF7
�KR������;��.��N��5�P�(7�u�(=sq�f)�
N�aQ�-u^�m�h�J����jb������`F�:�Zw"-��j�ʼ��U�g>�u����*�	��.a-�pŁq`��H��V���w��aƶ�`
yzȲa��fl�#�B�M�wXJr�3�4��*"�&�fM%ˬD�m\�;m�y	ba�id2��ݼ���Ha,'i��"��\�/Ӥ��X�*7��㵨�s�%����7�[Nj:RW�����ӱG�����#�%�N��f�U5N�өWP��zS2 B�>_e��oH�l%F���0�U��Ɛq-�	M�*�a�˱I���M�$0GWYڟY�U��C�Ǹ�n�k����1ʟ"�*W���X�� �l+=���ƥ��g^��"�h*+7%
�hõu�p\��1)��с1Bq��첄�ڻ�t
A6�V%x�'��k&���dl4�����eeͲqؠ�؉
75)�`Ji�/)݀�nS�n��.Q�7V��
3aOr��B�ܠ\�����GQ�#q
�V�9B��HD�P�&ZGuM��Axw	��[� ��Q�ӵ��j��ȓ8$Q�6�2V�6�B:4��"7쉺0��/hKgeGFf<H��5X������ZEb�Gh�7��#8!�N�E�x�#�'N��挴�]\��mV��,��j�C#�j�^�莆F�
jSt���,b�%N�ف^C��<*dʊ�jئMŕ��b2�ժz���v%�(�PaU˩��VϬNP23���skn�jHC����M�p�<�ѧ3솳&6q�j=vӧ
�)�9��ֆ��{)�wu�3-Jʀ��L��k���2��A�s�ֲ��x���T5�$�:7ֲ�hU43���l�M�%H�iGs� ��N���.�tV;nf�u���m�23�aa���:�+]�Y��ȱ��ʕ��ڧ`�s2 +H���Im&,�u���@6�d���dh��c����`�X�0l;J��:aL�m�i��&$�I��v�edf�Vw5���6(����k��S@"Y!����y�I��#.��74��c�w(�����ZP���h{HoAJf����w! ^����b�Xq��*-e��ț���;75�
HdY�9���1�C�e���ŹVSٹ3	��#8Y�X'je�UeT֑�Q7�:[�v��ē�5xqmI%�݁�Aed�R�!Y��j�ɦ��BowR_`�.��b.�:آ�y%e�y$����Ŷ�j�VR�p=E��Rd�Dt�)�P!�R��-��/6�)c5T2n\�����
�����m0^�b	[&3P�N"4hE<�j�yx���/�rl�ZrE�ǧV�W��|��օ@,%=#���z���|*�nk�f�b�X� ��)Ra��cPP)�p�oq[zI���ȝ��vɏ`
��+R����Q�Ք�f�.�k��%ۀ̳��#��tκ�r�@&<J;o.����V�:�A(�l��$�Y��淊����At��b`�7l㭂l�/qK�%�J^���� �crf��+�7�^bKj�b3Y	ȃJ�M1Gt+GU�l����A�̹�ETbFl@�<��X[ŗ��ѫ��ih4�
6Jz\9n�&=�`!4�
�KL�fK� ��ۺamn!A�ސ>\����K*�[a[�׋B� �Nw�!ۚ�⫉�)wJ�[sC�"ZW����ks(�ur�1J��leB��G��Z��[FV\�`B4�u/lU�hݖ�B+���;Z��fn5[s&��AoT$ʱgo&�N�1��,�dAm�{�:T3�(;���6Y��ԧ�!i�Fdr�+`v٩R`��H��K5��I{3OWf ,�,+��w��^��o1dv懈ث;v�\�q���@6Y�#�t���F<jlʵL�Զ�h�AF77
�?KP�[�ȹ�x[@<sD�R!��E�Zu��QW�br˦M[e^���`��`�bG*f6�9p�Cr��V ��ܭ/39��n�XZ"�iQvP�iRV��<;�3(ٍ۩��\�V쬌ؼur�f�+t��~H���V:��n�p*���2<�%�!7��	lEZ@������ �u)32��T7V�ᱪ�(vg;-��]o^�F���
x���Մ�w$��X���m��Xq�ܸ�i�7V1�����u&���!�ۙ�Rm�BV �]��6rk�%-QP��&�1²i�."c �b�IAR��6��<�,�[��[Pдe���҆�i��I��0 \G��#+�����u0��T��Y��+u�5̺շ�(u,&�46f�zo^fދ�u �E��Y7Z.�@�y���v� �n3�q@�=��Rhb�cE�wV5�W"1;;5޹�����Wn���p��Mʂ̧Q]Y���K���a�W3+oHBr��\+F; �n�D3D�`g�æ���-��f;i���b�Ѓn2͝��n	N��.��6�X�&B&
�D��h���v��hd���Mȩӭq�1$ĈS�S�ckk�kӖM�7>�i� �äE��ԅ�B���ͺ;l=�>Ÿs$4�A�È��b&q�IԢT4^�ܾ��ֺ�����9P���SU�6�Ưi$��׳67f�2�'[
�T���q՚���a�7v����^#m%�en�ؕ�P�F�+]�t	��bfBk^��XɄ��h���mRջ]}V����F����:�VL���aU�XE5Dh&8�lG{�J&���c9G�ʙp:�Ti.�z�$'9e����Y�X~j�K�n����t���Vu�Q˷a7�d�՛*f]]�]Ei���]����k��]g ����-QS�ЙUn�PQn��X3��`Vm�P�H��Q:Ž�E�V��7u�p*��h�9�8�&X�KJ�^�Pi̵+dǻ��ܕ+-VO�ܫ$�!��a��Q57
f-�(P��y.1E	�3��S80� דU�%�V+f9>7��C):���yv�j�o8�ShV�Î+�MY��d�R����ɚ�vf���fFlP�Qn&e5t.i�Y�B�fV��(�Ia�&�*�#���"`U�Mc����j��n�H�kn�]�j�B �˦��'�����R���[b�(���,R�m�Xrh��K^6���, v�hSu�Af��S\�4�m�2��.��2��DY�JbE���j�q�ָs�״�zK=�4��Qi���u���Tn�ʺdR������M6 �����>�4Aʰr�c ��
/]j,j�兌xq�ZGɭ��J��I�aCl��.���N�����Yx-]+`��ܭ��*4������ĭ�RYR�Fi�F⩭�ZM�ر.V$d��i�h���Jn`���0e�y@���#ki���v�3[�1Z����p<�j�2B:�ɸ��B�v�Kx�Ï%9;H�la:�Cp���Yr\*�uYoX�`��[�������+f�Y�ՠ�"���e|�ʑ�7�lĪAL��6��@M��*��n8��Ѩk2�+љLXA=��m���m��[@�@S�Ue\�ĸw��h���� �Q���*��MXU�^��\�]�u�Nb�KVw�%$�������6T��z�8���3n�R���f�H���t�4k�ȅ�q̇��v�4���C�5OXxT*B�$h�wz2fn���U�рA2f<����um��U�-b�V5Xv˫{Z(H�����a��a�Mf��n�W[��1<?Y�6i% $�n�YX^��]�EҨ�Mn��1X����I�3)�@��iEV�j��('k^C�Z۲3&�t*h�3fCCN$�%'GXߋU��6���צQ��Q}d�E��GcU:��	Ou�ܕk2�;n�Q���r�%+��I��,7��Bw�B�͔C��_Y�0�$̀��������n�-Z2�����.,j���4q6��d��tM�3]�y5��c&�<xkf���4�( 4�OOF�,v�A�ơ�xt����h��4�՜1�WJcw��
���n��F�`��&�A2���ٸ�C�
�M ��F�Iպ���w�x�谕��,t�s1�;�4.b�� �آ��@���:��x�(��e͠����;@�Zܻ
Gc1�w'�*�t��K���.�p����V�F!�GH�5��;�5v�s2���CqG%���d���1���m�Q�a�-�����2�J:6�v�a1X� �UŴ"{�� ��'Q�uq�] �f�Y��6rS�*(��2�������w���@ګ��-�0��1�6�Ґ����a2��/73H��؊�+*X�AN��4UM4IY(ȕ�Jf�;IY���Q�U�v�q�ƨ�*�q�;۬[����mܑPNF���'rxhQ�a�(Qys3䍍Z⨮�9�34��v6���))$���t\�����x�M�w)�AT��V��o([�r
�y#ٗ��)�N:�3,MxkѳE���a�i]���.;$*�Їo aU�a4�\Cp�=W�)����ZV*4��d	�2���:ы(�Rf�1���T�e�/7� �����м� 㛷B��C4�i��h��F�K*�!�cv�4s�����3�c��d*Jʄΐۗ
櫂B0�7�»&�a�bf�.˼/cn����R�m^O�:��Y���y*8�&�뚤����m��Bo�h�r���>s ���ڴ)Z)*Y�����.�έ����T]�΍��	�N���.�-��:�tvdl1]FN���T!�M.;#�"�d7�nev�k�!c�ٔ�_L��=�)�I7�Jwf�
*>��vI�Ĉ���&���Y�,^�.�c���n��;�t�wΕ�& m\��EgQ�˃q��#�ŵ9����z\.�c닞C2`�����4_@�lp�a�9劚ڷQ�N��la�� w ��M�}L0���hj�R�-dIRzС��e�5`U���&�:��!�-�x�݀rѻB�o8xj�ι�����K��UΩa�����o�u3J�������ϠU�_3��
�%l
�<�&MJ�㸐mT�)N����/���v]@'z�ܲ7[ޠ�c��\{���*�Ԙ�+��m�~O�>Ӗ6a�	�$��e�X3֋�w����Бp!)�tWX�v:a[�uN�Iv�,kK����m˭��F���2�"w7ox��-�_	r8�{�ݎ�N�@M��
������$�E.�
t0�9Cq^5��rj�:�Tp�R�-�/����Z�$�NtgW��f�sy��ή���[W5�Y���}�"�x�Yq+�h�Cv��"U�wr��(�i�ib�/��dkhvu�6�k�e;�>'�;��w�C��EPz˽ׅ�-|��h�����X�Kwʞ�W:Z�8:Wa�xo���e�P��&�qy);Һ���Yy#��'�ťH+*�0:��4e�˧:����v�*z����'�;;{9����0}z�-�^��ʰ���ռ�a�U�����l�����s;[�th�"�fȕ,��7}�h��w[vll��
1]8sp��6�v��t�+]J�fbO-�;h3�nZ�Q(�5tg0���h~�kYƍ�)pbꗺ�R�V	���e\�E�
<��8���+�Σ-:�G�û�iQ���o�8����j}���1�<�
Q�ײu�$�]8�B_q�[黎�A\�$�����2�%��U��3��u/xg�7N���é+K~HJE�-���	5S�rk�{S#���ɩ��i&i#��kF���9�r��d�P�X�E�ꚅy�]LT�zq�Hu0����WQ\U�X�f���汷�a���\�k/��/X��x��Ӷ!ت� M^|jN'e�̠!Ř'A������h����Yja�)�R���<�e˽٪6�Z0nrF��4Ρ�`�6^^\j;��5���\uYD-,�z��J�v������a��%�.�(��dXF-�m�a1�q�aop�W ��et�#�:;m�&]I�JȎ��-�
�N�*��ir r��5�>�:�IyI��UZ��vk�!9R���.{f�oT��l���ED��[wWkRr�kĎ>����g8�ը:Ŧڽ�3VpY{.�.��׳A�Qǒ��HvKo4v��nbz.�'hlR��n,
)[���/��ɷcS̰�״ƃ����c�Os�NQ���k�=[0.�4pt�<�x�3�k�H]7RlqЭ�W]
Jl�W�wfE��4_��sA��^��k!�E�[I�t{.���-�Ѻ&�f�V��p�.h�q��C���f"���4�\��#�ܴ�Wj�����+`t��j��l�7z������9fij�����=��Y���.�����9�c�3')J')�UC/&hU{s'=�ˬ��1��D�iu�ѵ�>y�gY�1��
�F�.R�pj�n��7)�+k��s�]��T��kkv*R��x�v�� �r�]�;6Q2�L��V�A�o
23]���>ܦ�u�z)Xd�N��WY�X8�F�]̦\߷�U�*���Z�Jn�\D\�{�ފ�c��B}�̋�
.�[�a�y�SՔ�k���ucd�hon\V���HN��Y���j��d��+ur�g%kkK<jJ�v�KK���A�X��BJb�R�b����/�ذA[�l;�Q���h�5�(v���ή1=S>}A��Ϗ�b�씸�{�������ԓ�B ��3+���iRӉ��ӕj�S;�v�*����9�%�-����B�}�.R^�mod�N�	�xD��T�g�L���Dc醳�*^V*ݫ�o���K'QW YN�f��+�}����ˇ%��skXLz�Z8H� �V2�x�Z�XyeЧH�S�"̮�M�ɥ��y�V�1�`8�v�ռ��H�W`%CV��*f=��r�n� k�5'Z�ɺȔJK��b}�Wr�Vv�r@#�}�3��9��Mu�@�o��1X�k3pZ��洉�f7;s�4T��]Y}��IGɍ�Y�9]I�FJ��>,7]M;�S�ց��>�}*�uM�Fq�����{����y��*������HwV�C�/3��H��{0v��6���r��[n^nJy��aN���d���f�K!t�j]e���(�nb�.�~$<!V��e�U�WN�qP֍*�b�1���4=3r5\#^t�;3Ay��^r�ʴ���aer6s*�x�A�2��C4�u�G*MǷ5٬4��3�e� +�-Ш»��Y�W`�qQ�<r�*��Zr�ՌP�)k0�8c��]�Tuoe$%9�ja��X�Ώ�-MZ��h���pק��H77�3(�� ��ܸ�E3[/����&�-�&J�N�5콥���@��-]����!ZXkhTN�)��I�fH�j��еJ��aq�����!v#0m1��b�Y}Xe�/K{��

s��w��܌"ER�&7��	p����*s�N����>��T���> B;	iڵή���s�Q�K:Э�z��8�֟S�ruMb�.�W�]p�ld�g+�g@kPv�\��\�V�Ӧ��P�#0�0ɒ��7�wafr�r�f\Bd�y�.�m�E�gGb�4����F��0]��8�7x�32Χ�V�I����&�͒Zf�9�q�����5em�굪<�g�ռ��]��Om��a&�EN�̌%r��]z���4��[����.nL�9��B�Lӣ�P�· 40b̾�F�*OI,���<X�+v����SN�(���q��3{Y��-
�m��F)��M�!�K���ZlP��_oJ\��f���n���Ւ�_c����z54�K�W��R�ʔ�
�|��:b�Ҵ_�G���\��Jȯ��˧�Ww�5���}~��T�[�C,3f7>��*�s�O@S&wS��NM�e,4�@��(��L}�V [�;�NŐ���γk��-c̚B��v��B9��I(��6�'ca����f��PSz�@��;4ݼ�)t�`��Vt���kR�|����>��;GnQ�
�)�|`�E�)��<��Y����'�_�e@�5p�uaMsE��vq�GU��0��X�v��6Cǀ�Q�/�̽�ZZi�t�uHt�D޼����k���r����d˝�q>��YM���+�]����2�ehܾT_�x]"�v��OUЅ�i����6��NA�v�ޥ�a�,vӖ���D�T�)Ò�Bu��sB<q	��s�ǒ���]�6 �0ܷ*)Q+������m^����/��F��u_;�B��lR�T����{,�eF��X�����{��&�!fn��ʰi�Y:��s(fM=e%��������%�2�jLb�-��6����#A�" (���S2s6&��!�h�.Z�F��������`�U�Â�1KA�������':���l��ܜU�G���vc�7)ظ�%�S+���Vq���~8��]��"���oJ�Ԝ��[�Y]�}�i��;�q��q��j��̛\��By��[|�[e!��J֜�X-r���T�љ(
�]b��e�_�畹�����Ȇuh�v�v��<�KL���sK���3�hs�������_N��%ob���znϚ�"�gR�Վ��q��s5��Ay���(�ư�KOV�Ro�W;1�=�(ԭ�{�l�+����+jJ�!��+�λ=��q����]4����R<R|��o��c�Y')k��]'��]<C���\�l���|ޢ�m���w:��^T݌ʸ�.���c-�W��%�۝��p���;N5ty\q��'f_.�j�Y��R�����EΔ; ����2@�6-�Q����:�`�Kv���YȭӉ�u��Ζ[St��]n�����AyHNዤ��B��J*��=�ʝ��n.��T�	Kl�Oo�ҽi�km2o��}%�88Z]\��ʓt�\�r� �©�Ì4������ݨq.���r��*����v��x7i!�*'�:�8�=FV�3����C��o������=�K�T聋����֒���Fp����vV�^56�ՠ�<�By�X(L��ϕ(�=ce5�z��Ce�V�TT2}��������s�=�R_<�/d2X�ؐט�ͳ�8���e�5�Z%%ɒ�fJ�H�ۉ�4tfG#�j�]n����E��8A�*C��7nV,n�Xw�g�+g��Z���)L=-�82ue<^��@��f��]4�ۢ�iͰ��S�q�u�*h ���ٚE0�����֫�S�'a�x�z8.����u�F�a͹���p�VlY�>�-Ί��%ǥ��(��K�H;G�<۔��Z��[/v$�+
M�s��s6�U�v� ��ʭ7�0���ɂ��s��m�1#����tоζ�qMY3����jF,�b�$�[[������0��>qj�6�µr�I�?���'V)�L��h�f[�sb�ۣfN�9�3zg��R[�j=�z�[.�����Qjۖ�Sl%v�ن�ɶ�g=� �of�!J͗�)Wk;7�CM�R�#Pt��Q���w�I�xo�-�#	2�X��!�V&�:�ξ��J��V�^�A��6P6��.f�R�y�ܬ���;�a��t�To����|^�s��$��6��ӾV��oi���S��0\�'�tW�Rб���9W��wP#gv�4�Vxy;n�}�Mv�sXk�;
��*8�}�n��:����P�+�v�K�,���������|��K�-������a�s��U��%�p<Won�W]�139���8N)E�ܫ��U� ���o�-��ho3p&�����-]�6���jl�{�!�,��Q,旓U�Jt7}مf�$qMx���Z�a�r�oi�E��y�N�r���vJ� ]$(68�V�����NV��;D#e�l�Y��\������u��l*����B�r=I]d��O�������r�r�����|&#Ǖ�S��0A�Y�Z�M2J�4��Qj�}P�.qe�"���Fr�A��빷J@y*�Ӵ�[��sQ��hU¢��Dt�ћ��2�&ec/��r�B�
_N"�_���*�U�R
���8�p�h�\=�2�c���C0k�J�³�����4>&�f����h5@�wo�	x@��f�R0:q�@K	4��'9��s��;�S�oR�hPC��u�j�q�Z;+tJ1]^h���-���'
�{MY��o}�|�y�"�U��a�͕B]	1���EP*��gvV�[W}zk`���O�[���&���T}D��Z����t��k�\�n�GBX�X�cm�{ݝ+j.慠�H�̩+7@: �tMZ�M[�⧙�������36�<cs7���z��F�F���Z)�G4����g}s�X�+(ݵ��V;A[�Aap�3Jj�:a���+.s�X3 �ϛ�r�ۖ47�v��T�{x�b�!��%�ު���8����'��L�`Z1�8���5z{�>��!�(2�.��gx�;��[��V�@|82*�Ufg^N�*S9&����n*<�]+���+81-��;N�af]3d�<v��kw��C�c n���[K�j�Eʶ*Mqn)M�kt�r]�E��E��
��g��Y�y�R�״C<��)<��J�|�̮s���:��2#�V��V��A�1����|��u��,̄*O'�u4N�Օ�7S�"�k��vP���6;+eum34I�qkݚp�'�Ѩ�Ysh�S������2U�[���ݑ�����W��a��n�{��뱘O�,�4�q�˺�-ż��s��\B���|�ʃ3��-�FIN^]����4/$闔����Ye=vC�FY����Y�w Y&#�y}��[N��(�j%wӶ]���%w�8GY	��,��H	;J>�"H�L�c^- or�e�C{����V���$.���6�W�p���쏤�jF����U���]s�77T��B��i�&�N�]�/�t�h:춤��N,�p��s�I�Z�����6V��U�*䌺�.R�*�;��*�r�CD�X��W+��_e���T��������ͧۢ,�M�����eD�ijܮ���&��u�W�jWn���E�'Ж\�&��X7���>a=�Ű�{�U0��2�"gL���+������3��!@�_5%���Er���e3�����*v�E4�9��UBz����;}%�sl]]$A<k��*Y���.��9��
���`�s��5]`U��yN��*�q���y���Ki\a���S�����1v%P9]}j��Un.�;������{�y�YE��oehj�M{B^Zb�aa Z�8����ՊyX��nv�� 5&=%�8\ѓ��(>N���r�粥u��A;+�7*��5�mѼ���ʊj��5�bb8�$�-��\�<���K�F��¶<��u}$t�)��t�:���y%�g)���{��kmm���;m�km�����������&�or���5��]���;ARm�h���5���g*"�c���Ǫ�gq�Ri�D7ӊ�a�u5�]u�H�II�G8s�X�Q�.+��F<l店[֫,*��Є�_MF�[n���72��g=�ve��-��*�|.�x�b�P�g<�zo�r�rn-m�a#>�C���]��5CP:�T*��V4Zƭ��o�;����u�ƨ�Y: �3��[�p���]k�.gf����v2oT���J�J,]��[)1��ʌ
�칛Ҟ��#{ݸ����u���(I��"5�m�Ϗ^[薁�]�6�\�� i�ٚv�<L|$����n3������y��W{�2D��d��q�v��h�,��R��:�b�h..���r(_��8ܻ�L�PQ�;1p�wte#�Yf���K��ȠH��q�ٷ���t�M���vĮ�;�ީ͛&�e�Q���*�
���tX'`��_�7�h�μ�h��E�Dt-�7''�� 3$��B�N�ne���Z�m�{�K�t⩜�f�P�2��$؜�ʂ�Y��a�n�Jq����sR�����pCn�.^�\	ͫ�W%1���)F���JAO��`��u����Y���*�l�'u�X c�ԛ���Z˺*�,�O�t7Gf#u2N��աiv�h�t6��=Ŭ�ζs���o;2��ݘ���R��z�k��w�E��3���t�ٙp�!Uu�n��ƥ�������
K*7H���r�Q�(�LSPZ����^I8T�`b�O`����O8�5��*�
�d�X�r�l���³h�����2�3�aL��L����E+q,-r�@a)P����X/�Q�ӻM}����u2��WB+`F�����
�����4� ǁ��I�y7�5a�C���] �Di��@v�zܦ��S�M��Wj���jV�Q��mAx�F��F������Omܠ&���v8���80h�e�giA�p
��*��5�h���oeDj%xM���vr�wN5���+40T4���c�b@��`�� � ���^��^V�_�.����:�3g	��@���:���t����*���]Y��X̥���*�,�)CYi�@����o�pS�czN,d=ؐ���0p�/��qή�!I��ک�:�y�ׅpպ�YeC�5Gyr���m�"!�uơ���zy�yO�e4�ݰd��A���םF��M�!1�]݅)N�v5�XO��2f�݃�]&��:�
��1]���v�%}���w�e[�sa�A=��p���]7$'�v���H��a��:𭕗��naK���:��;�f����%�)DlL��9m %1�Ysn�^]��v�2VVJ�%l(T��2�����
Uܩ�B�e��_�	8�B9$��6P�4kQ��aD.S��Ӝe\v�1#�m��ܣVr4z�}�e���C�����.3�+��*��+\Bs2�YΘ�H��}ր+OqU�8K6��ɛ\��%�ĸ��R[�>V;��E�I)v���}��bb�)̨��Hpw�z:ʊ�J��ONa	]��~���m8�b���`�L��h}���#X~n�#�E]����1tT`|�z1�խ�سٕ\B����Zr����,vUŎ�����wc��0dez�l���������U �XQ���f�_
Y@�7wVQ�4�|4.��ډ<���d�0՝�a�ЮV��<��3�@�̒��ڮM���7AGQB3e���2��l��/WP� ,{MX�Jpۇ$�Vn�e�4�"��G`
�����"�>D��I�����4@ڼR�e']�)AR4p�(���AΈ�U��6�����)��M֕I�(�y��FS�d�.���u6�ѭ�r5�@wT/3-���hF��7�\�$���bK��%d�0*��=ޤ��N;Y��[�pʚ��:d�0vr�Qj�^.��V�@�0�7:��p���k�T�9f��Vړ,��7Iv+qfNE��֔l���Ԥ��4����q�pq���o[�G9�9$����VK�`P���Z�ə�o�_U��\�)i�8cMN�I�X���mtc�pP��:�,c�fy�R��Ð�6`���Vk��V��ݑ�*ʭ����v|�64v�H�@�[�G�]�gi�о��U��r�*��j�
�*�+�[��P���M�j��v�e�U:E.[�΢�nqv+�DF�c�kt4vܤ.�O�N�etW�S�]%�n�fa�9լ�����]��/Vqm�on<O!�VJ�\��V��$qwyx�L�%�*�{u8�B�
r�W'igwZ;����\�+�H
����3�ZH�hH��.>�	��AGC� L2�kU
�)�8K��9�Q�i�a�In�Y*�u���j��6���Z���/�=��M>��x�.z�{��mt�a+���F`��5KQ)��ͦ�;��ֽ���Ńdk�ݑJU�f�/��TX�%���5pZ۲H,�ƒ�-�vuq�G4�U�9�"g�a�K:�,�AS��[�x��g�z�(z��L4��l�l}��hP#>i̲k����bL{[MjǉYeL�.t�#Mt,��0_m�.��(nZ�̄��7��7>���9C�<��
�KoYG%�+�kJ+E�� R�8mG�֬���r�y���\�AA+�&p��k]�+��{q�ھ��%�Nۭ8�]��x��:_"jW8iL��U���x�B�Pێ����[B�P _=�T��}�r<N! Q�"kkn'x�P�G�"m�D^�κ�Ƭ@d_:(:�6S��j8���]�#Qa�u�(��T3���r�ʏB��4����N7�x���ʔ�V'Z�COSO関ڝ��]�N�@'6ç���s]H#hʋf�x��\w �a�[o��e^6ӕ��X�r
�j�9�����k�{f��4�r�(�AM���c�z�� fl��L���T&�I$�}&<�R��-:[�8SS�_�P{�늡�q�d̲�+b�x������$+f_�׵�v�Y=T�9�3��6�t�1�(��6)T}�.ă]����0-�i�WJU��I�첖5R^���$*�k�)F[�U-�3U�k l�`;T�z�Wº�x7����a�w�**ۣ<�`ô��_]�#g-ŵ]�]%BM�y8JL�C�vٕ�X�|l���̲i
�R̩׀��;W^a&�a%8Awxc��MT1e��rȢ��n�i�Ư��Ԭ�Ԓs��/�|�>&��wE�O��pC(V9y�̫<��+w)<O�����s��GU�I�:�+��/���؏TL��:p"ʫ�s��4ӱv��q#�S���(F�o~�:n,"����8�Q�[ɗ� }RY�P��ت����[�qW}Qّ����s���Z�;�ܭ)s��������G9tY:��F��M]og2b:~�f�M�{�ցJ���kۢ�h�m��@e�&
�$�ǭb������8�Un��@I7o���m�[�͝�R����;��-[�zk$�X����2t���1��v�Ŭ���.x��P�����'b�f;��fu&饷�@T)���H3�e��n����V�'��	��m�l��3抝r��cP��<^`ӟ:��ݼX���a�,3��:)r�iuQ�O9�|��q��z�;��(��ݼ��\?������3�&恫�3���c�"��0Z��\�3{C^��s`]�t~?%49U�g]2�7&��:�{�Yy`_'� � �@f����HC�nGۡ|��gd��{��\k�T�<�j�ykX�s��
�� ���lۙ%JB�����s-���o
�q'�F+i�u�]�����v�k)�˭L�1lUo-Ϡ�0��C���bE�S�U�w���WE�+��5�y�0J��y4�������sN�!���QP,f��Nql�bѳ-\x�
�6l���v�Ol����_$�ʓ`��k5�p���m���Jnn-+���=+�Tڭc+�!O���d�;ui!��p�fc�/��i��B�!:��ٍK�|!e��X]�)��"Krbp��(nX=R�Ӛ�E�o"Aa����g4���\�����(�|�9�Lм���\M��w��B�L�� ��˫���<Ɯ�,&U�/���V��&k�)��=��x�}X�f-�,hm.�z��Y�nr��5�g7��5� wO�*-W8
f�p�|BF��+��-�N�;��U��V_e��L=��޺�K\�*^E0�l�S^����G��ٽ������֕7�B��� �qW�#K�j1�N�p�֐ܽΜ���h�V�2Hw�]ۏ�6�Ia�ffT& +�ʸ�G�Բ��W�+����쬺��?��n��妹M�w��|�ݻ*ܦT�M٨>����p�?����۠r��fp��=#	("<N�)eY���s#%L���%
}�Y�]e[�uHe����G�Ջ�yK�!�H��ӹ8���/YtJ"J��h\�X�7�샤�jAElke�b�S���ɸ��$�M;����c��Aڭ65�7R�1��Me,���
��v�˱j�j����ꑞ�MꦹS89PAi��mv�����hs��9a@���0.���Z�f��൅���L]�U�ùz�]�QW<���I��䫚�B��Հ��Pܓ�s���pn7�`]fZO�����U�Nm.�*v}����^5(Wf`H΍-���๛:2��Ⱥ��-crB^㙛�o����6�Xr�9w���,���ڲqbV^�a��6m%B�:-�u����Ξw�V@@�:(l)h�����]W>�i�@�S�9�6K�cv�ӫZì(��LVf�.;D̛
��P���w�+ ���0(/n�F!��te#�EL2�7WM�����.[���Sv㮭Qs�jWKA��G*��qB��;^RI��K�����lg+ΐQ�󒈡b*O[���9-���n�'B�;�Cq�Az8��3�=jA�&�ԙT��Z�q�h���m������QN��:�~�
��`���6���	��N��B�n�^��@+`;Պ���.(�-2uA2Q��)�޻��f.���Ӓ�+�H@��R�T����/��	��J�W�w��O�����SLbRf�+w��;����[�p^r��ڵKS�c�{��E��N�Z���� ��2�dUAY9m�vk� �	�PV!)mh:%J�y�)����� 5gREz�6����8���\�]�$3u�P��[�z��0^=���� �\ ĕ6���8�F��j�wY����: R��~ɜ�I�t6�vBw��Q�����tL�f7�D|zg$�5�ɘJ�ĴԺ���(�aم>�ܘF.WA��wR���7W
�PXo���/^�a�Gq�2��7�dW��X%��+�v��=:O�!�S2�,��%� R�7S�k���N�]��$����*2��䩼�@ba�81��4:�7�e^���5"K�Y6�﬎�/��Y�j� ܕ�>q�s)����K�f	9M}V�0�c������Xo.e��h<�fD[C�7��`�j�p��Y�&9<L��\@H�J9�,�c��ŭ�vO��JX��@��(����m;�l����!@ܥ1��\F�T��!O�p��J�nZX8��c���hES��Ep��)J�yB���gF親kn��%\i�em�֍��T�+��8c*���-Ǯ�(&��!�ݱ׮�Б��a��X�I��f�x��t�U�������E>�Q9sN�F�g,����Dd=��Ko:f}�z�pdד��Pك�dŹ�I'%�kw�-dh�`˦�&-=W��)�A�R�^n��kL�t[܁���b���,�@�]�t>h��F��勢�����s3�N8�w*<�H�F1�tk���b�@2XLԻ�%�A��[}ʞ�I���G4�M�������P�j��T4��`�k�ϳCoQ�o��D����Cy2����X��A-pӨR�m�ȵ�e���8j��������)Z�o. ��h�%b�D��گ�0�/��Ҥ�\B�2��lD�5k+���lR�pU�����Iq�A�oX`��ngkh<�*|�mI�i糃���7
��j�;t��3�m��pP�4��t���Lj�lYx�������R�;q�1iӠd��j�΅m��̡ XǨ��FС�N�"����uq����s��d�b�b?'��&z�fޤ6i�r󑹊�͕���L:��m\jY(��͖~!���'����� o��P���Ĩ�I[�b%�t2���ź���T\��x4��d2�ٛh0�07.nB�}Fum��ШV���P�7���XB���]����OF�˭���@���F�]��S:V�4���V�f�AM#�Ƙ��n��K��e+iҮ�:�]`lԴC;���+O.�]�-�UA�w����i t�����+� �[=w��/sA�ocB�i>���j��<ྀ	��N��F�ڝ�#�e-ur�YS�n�{e�՜�ue��^��l�x]ֹ����pXo�έ�$0������Bi7����VZ�r� ��R�($5��i��䤧���:����n8;\���R�}�{W����R�Wvj��y�2.��й�9�s��4���q��A`k(�ۗ�Y7��ՔQ�,�6E%Y8��9P��Z�*U63r�)^N� �w�h��L����X�庝M�oM��N�ql4�H,�5(m;����NSr���v�9�Qn�CF�h��.���aO?�}��}U�}���ޯiNGW��0�!�q�#FoB^��[çb__|�N�M�˙5.	j�Q�Fv��j��H(��Wr��:K@�ƋgП[}������V���2
n�|ifZ�߂��7�*�MB�X[�B�I[�3[���X���e_�w��nd�W�E&����;t�i�]�R���WY�,�/=�n��u�L�~���e@Pr'�FZ�٢g=}D�w7��oh�lRҒx~S�ۣ�� �d��{��;�C�(���j �Ȕj&��h�'Tg����,*�
�m��^T�B�P�ͼ�J��h��2��lX��6H�,���Us{��-����/n�>��%����;k!l�1�
�����lgR�B>p��m�e�7�}1�WZ0I6�����nin�����ݹM���c1�2f�{��[GE�\%�v��Xڦ�]�>}��u���ϊ�ml�&�4LɋP.mݨ�Ke�9wEgE�S۔���"�����8BR櫸*��{��/d7ziN<��. u���d��1�QňN4� "7�ҭ��f�d3�G#�#{���@: \v�_a���I2f��{Dz���D�fm�h�������N���J�|�m�p�d�I'Z���į����k��K[���/,�b��5�)�ޠ�ڶ����"��d���in�}�j�!��t�����A5v~{����w��wk�ŉ�nnwWh��L���1]�V#Q$\�D�5&'v�E�j9�����ww��B	\�r�.sa78@[��ō��l��wn�Bc�ɻ�1-IFff�r��Nm�"���1��e�]
�L��D�ݦC$��\���1�d�)!@"n��,QK����wvɓ3Q��ؗv��Z (ܮQd�D�1�PNQ�1]8P;���	���#&D�wu˔��;� �2wtF�F�I�X9�6("���;�w]ݷ �Qh#UҸi$�D;�&e�c���Ҁ�%"��$�_w�?���X��C$�`a}tkZ��Tq:�df�췉�� ���'���*���(p�����z:Ӄ���g^��f؇w���_��n��Bj�9L�N��
{;.��BP� A�y��S/_��gOxI�нqi�W�>�y uD;��m�����zUu���ҴїV�t;�o����n�
d|�[�ݺ�И�K�vD�D}�w�ƫ^��{�$�1���,Mn��̢�;W�Ù��/�W�N૝��F,5�Fq�_N�[=�DI���߹�n{c����މ60��ݦn%�ÙUB�S��Buv���>G�5]�.뱏A}ڒO��2$8�Bl��t!��|�3#"�uM��U�鿛��3o�k��뎋�ټ���c�J�������`�ePX�5���L��$HW��OS�#y.��R�usl��D݄-��}1�u#'Ұ#�� [�7a{}g4�l��OMA*v	��#+�O�铟P�p��F.%�cl��p���'I@_��B��F���6乭fQͺ�z������xKM[��2�ƈC:u��6��l5$���fiZ�lP���ml�ϯ�d����d�ىֱ���FY�ѽ�\�MG�E)=��U; )ӣ�M47����F���8�_K�R�/c	N�X��q��[:7*R�c�ve	Z�v�];�����n^��
�x�{I�{)�o$��$'&V��Jp�F�x�;�zy�m�����e�g�0�*%� w ��8��n�`m":��#����s�щ�ڿ��҆�;��7pt�g�Θ�3Wh'+��]�ƔN���� j���ĵ]Fx���b�PF��V�9t����M��f剁�qw����t%��2���=��q"�����E��tn�R=iW�-h�m�UH;'.4=8�fLulknT93pl� 4\0	�U)3��;�ы�{^mT��v����-�3jåp�S-�8Pp���mTH��̚7�{�`O`�a�4�*�WN�()��G`�5���N'��N���z�WVj�;-��U��I�q���&�J�:�e���8o��.as�ϞG#�2b��\;�S���zpN��cb7e�q�CΟddjt��~���X��S��rD[ͪ,ۼ����� ��{��Cd�Bn�<�8_ݶ����e�fs�n���sC4����',��<**���h\:N`5,�>��V���x������d[ܩ ���v������7���K@psW7�Pä�gF^�@ȵb/�o�5�G������!6{��=��g�N��̵X�q��,V��B�����TNgJ���q����hC.Q]��j��W-��r��7:�)��3e��Renf��ҷ���ďԭ��b�]�׍{��pT��%dZ�!�`�K����?n�k^Uz��'�0D�'��"�ow$�/��Wm����/�fۨ�zjN���0c���%؛rN[2��sl<s���%���&%_+�.�6X�7ܶT�_oA���D9���PB�o��<��1(��(��žC�eJ7�(�N���ä3!�u�P���3"8(=N����i'����pe �$Qه���K�o8H��,`�yM��#ۘ�p��aT	�#���wo0L��[���'�a@��U��ʾF��_b}q7-�p����?N.�o��MF=#I'0Ҫbj�SQ� �L���ط�ë]z���xs&s�;r�B.����%Yw��%���k�o���Ѓ�)�W5)& !3�*1�aZ����Sb7�@����~�����l�1��7�����p�/���.��$wU�zƼ�=���s
��VrwJ2�$0��1wK�q�ԇ~�h�ޒ	m��},�Mk�Ahgi*T��Gu�'����Gu3ٴ�V
��f�������f��35��H�ͺ�K�rs�2TY�9v�\GN����^;��֨�[�7dR�izQܼ�+
��*ے�Y���؆G]k���,��D�S��b���/Eg�$��I|VM�gd��zʐh�U��ok��M���iMߥ�<N٨X
f��4����ތ�
ʽ�l�u������,'��RQ�?j��6��O����p2�X�uLE���f����B,����+)OZ[�Ռ��+oj�t��	�@؞#uWJx���iV
�sWx��0�����ʸ�@����F �	i����]��^����GKTdx�YYU��{ĢX�hRD�|��峋(��������,���\&���n�;5���8r�.�%���;����=ů�jۑ���z�t�,�MC\�2�ȧM���/6�F.4�:hC�Wv�Y��^g�(����"��p�@�m:��.�,�K���P��G_��Yg8�%�{Y i-�y=�Cq<�qՇ�h
�~�U��JB�C#b�S-ތ�q0�c��V�S���k�+ {��̥k켣��@�ay�?`�4�[.�Y����E�x{7l��7�S���c\7@v�{�#mU|��h��m#�*�Ǯ�]���j�CGe�����z�e�Hgo��^�P�/9�J8޳G{n	�j�sf���D��e�q�f��}͒8ŵ���\(5z���p��۳��kP��'��ǉ-��!�]Yj�o�������B���h[�WV!Ԯ��6u>��Vl�*Mт$�3`�V{2�f�)�#)*"ۚFiL�"~��8�rE�U�=�9�/g\�W���U�`��<!��F.����m�Ϡ�H�As"�u/�T̊�2Q�S�s+a��q��suTvHrq�к�P��,;/��\��Cj�8LZ%\3_D¥Q��	>�Q���I�2�P���
�A^�GG"���i܏����hxX�k�;��y�^f���r�eS�yҍ�F~�9�a�ee�É����n+���s�KV�!����X$�$l�
&K{ԥ�p��΁��ɡ����������+ynz�q��U�&2�l1�&�������ۻ�� ��H���n��ˮ����^�pG��uFT�����V��>'���.��m:��$�cn�+�/��eoVF�.If�TQ�v�'�Ө�:kz̜'�ͭ0?T�?T�Nv���Ʋ�T��u:�uOi����(�=����9Lh�}ν��[@N�Ua
�|;O��0</�5�6xe��x�f����7��;M�Ab�yH;kDU��l����V&tveli��s��#���Y+*	y:���ߚ�m�t�#��$N��gzKjY"�Z!�	�ٝ"���^$v:�ʯ@�ôOT�e�p�^�Y	p"E6�^��wȪ��;�e��%+K(�a"�\2�Vc��I۞�u���TN��|/�`wg�c�V{��/���#�N���j�M�:]?R�ŏ���he��'KFx�+�Α�ƠhP
5�]����D!��lw=rV�p��,���6b�Z�7"r�u��J�ipz:�iq�3,�þ����5O�W%wUw�,��"{�-.9�e����y�Y6���l5�@bI@,1}��[���lZ7���C�}Qn�2��zg��Z�#̌:��?e9�!T
��j�y3�f�'Ra��c��O/��d�1�H�;<���3�+������p졸�wq���6�mپ�3�k��(�hw�g�{Gg��gV�:�7]1����Wh�MZ��&zv룓+d`"Im:����0Y��~H��"bVӣqґ�ϒ���ֆ��K�&��������Z(�s�X~��E�B��T��L@	����[8F�����"0eov���@�1Bk��mTH��̚7�n���
��Q%j�:�P}��R�+�5�Y���":�� ,p�Չ��n*D�Ǆonh�n���^r�X;'gJ+t������U�#�`C��N����V[�)���f�M�P�J%���qa���JM�P��nqqTv 2�wg�u��x�֜<���ވ�j�buw��3�;�E�ó���ެ��v{��W�	'U���ɯ���	�ٿ��+�4���ӧR���gVԔ��*��v�r�&/vPzdXc���q��Fk��S��b˦0�ހ���޷{��V�,.�^��*��7Yl��v� v�b�gY��Y��T�����,%M�!�U�<����w,��x�]��s��U����� 6�u����+�+E�ufJ��q�����v���0U��8/"�i�>&����u���W��ewPk��Ϛ�>�|睙�U�0Y���x�OO��N���������Z�L�ؙХ3�7��O�T���-�n�	1_bu������G�����QCWA�ق���i�H�z�/v�K0´4���f5�q�V�l}k�Hf9������q��'3>ʑe�+ӈ=ԅ1�0��@2�vc��+��t�p�r��)��F��u�y��^�������%�>���l��i6�a6��7b�|�mSi��z]#�:���b���Y����C3:v>u��n��X�W1�k٬��M��Af����Z*�����>JV��8k��YucE>G���0�I�Nut�<�ֻ%c���"C�-����8�ɡ��f��t��+bPSҡ��n�i��'KBBV�Ȯ�@�5g[uÉ�s m:�&���� ?x|�s�lj�}����j�8�gJ6�Q3�O���9��ϋ��Su�3B
S$�7�H� Bg�z${kr�^<�(p�����OQϭѴ�8C\�%T�$?��ҊU=7���dd>ۿp�gc)��=Kʴ �\3M]H�M��懮�v����0������T���9�BP&x�w$=RV�{�1}�@�)`���OM�gF������
e��oi�9q��3%�7���r�o�1W�����,�uN.�%�h��<�/�SX�K�I�C]V�z5!de��ߗK�yS��]V'bx��p���2L`��l�G[���3hַ�9q���X�d�&��q��]A�^��u�ж��������U(����nT=��\�͚�{���p�q5F�{�<U4�d��y5_o}�8؊�9�`�d�u�Wk�܎g���F�y_g/�Ւ�࿪v��͙@-F��S,wM��X�w=�z4��r�㮜���g9՞�C�3��=[��^K��VeK.u�)�f�[��)f��xVw�>�\��e�E���E���Z)�+�.f$�C�b��ՒUq�[��g�8����n��s5.��e�.�g����EG\�I+�;T��2���9��/Bߝ�k3�� Ӣ���"�iPEdiuaf�_Qj!�r��\m�GbYp:��B���=]�"��n0h�����*>Ґ����ح�>���Q�o2�\���q���Y m?���M�Ό�<�fÀ�f�~����n�l�R��:C�>�8�ׄ.R܈�=�N�wi;>��C�m���9���@�c����<�ʼ)�ǗT��(C���ʹ]�ʜ�e�O���L��n
�c��y[~�"����R�DC/2&��>�n���8�Fo,2�j�|@r���F3�b���)�f0�H�s!>LO%�}mH�tVi�Z�����`�a}��&$��uΡ����e��*9���C�����W��� mk��cCJ��8n8S.����n��ߑM+�Wt���HA��?TrT�zoNe��o����X��ma�����sE��j�\@�vЏZ��kRڗMO"�Rr�*�����Q�����Q]E��ܰ4�jŇg�œ� ����t��J���z�E���־�;�ixQ崦���1��>�F9q�~ٱP=g��'tWH2��>�n�4\�s�UͻPʰ�{n���/�i�w`�3��	�7��$떯��#�P��W(qB�	Wɣ��,a��g185W�X�֨q�X�e�>c�Α�gyɮt�f�CNpF�N�D.t�q(���.����, �k����o�'����ޝ�:�.w�3�rSG���̯!Q8�g�s���tf���l�iD� �Z�ϴ�n�7���n�$c
pe�NQ���������j�3�C�u:�d'V;��#d^03�������S�����*���<6�0<.�� ����(*N�	�6v�R
�s�����nsW����~[,�ی#���ʠ���<j#mP	dG��}e"E�K.��q뽉��Y#��w��e�5��|�J��p��J�,8sW��G�mg r��0{T�&QJ9��@}R[���|���pً�Z�7"r�u�d���N�NK���=�*Q�����s}��s�ۄ�Rc�08�Ù�5�[��2�ƈC:u� R*Ǻ=����eu�3y���8��ce�����e���Al���./�î �?e9�!P"I�!J��jO�U"���Q�� Hq���;<��:#�:%�\{(js�H���HfoZf �S��;k]a������v�QYĝ�c��}��<��Z5�X,;Ϲ--���Vd,�Dmn�ѕ� +����\�S����J�P��+(ĉ��w��[��0�cA�\�廄V�V�3��4s�y�9rĲ��K�y-:/��H�튬��'��]�.:�Ղ�'NN��e����g*4�l�`�7>sZ&C��v�GK�Vd�o�<s��Cץ[1h��=}p�scd�l���s�!u�I�/��o
���S�A�*�+��g����!�YQ؜$� ���-�G>r�R6E�@���&;	�1�<<&���辨h@7;B}l�*�Td�(�ٽi�mѬF�DNn��r�6��\�M��u����$Ƚ��}�f
T��<�8|(�LX�Waߡ�{��C���;2����A@23}\������
�Lq��:�e1{t���Bq.�N��A�:�&RݑЬ������̻��!P0����ӏ��b*��9ٕ�]g[��v�Ni��C8�=���$Z����͜z���MX�bW3��pX�M�ҩL"�Q3I�ja�+�j�BZspu��jF�)[9m]g+ݸݖ�.��־\�2I-QN�Y��s�&�E��k3is��-R�oh��ҏ�s	�z��Ɂ�<��NY�XO�veryt��z*:�"����mJ�*)Ґ�!&�o�Gy��O6�Q��ՎID�o,�%��w�P�lI_�<�v���h�Sy�O��i�m]�Kr4��1�b�8T�.��gIp嶯�DֶW�\1�6�so��oS�����bV��|%ηF�j*ұJ�����z;�D�r;���1���YR��U�7Q$�py{���M�ʾr��*R����"1+��-*X��=M�*kY�M�U��<������ݪ��=�"�w}�tk�u�<+�*RR�����3�h��Y���UjU�;{�x��	+*SB�����,md�����}��O!/YV;k�u�j5��:)��N�/D�a��,�2H��<M�.�i�=w!�Z��`�T��]�ZXbs�f���ҩ�޹9)w|M�����$�,LR���ݖ�����G@����(>%��;Y���0��9��)��@�T'��bՊH飶\fT*� ����xV:Ҹu�2�e�!�7 �tbb�q_�I���I�q�8L�F,b�PL+7 ��(�i�4u��­���kz]J����]3\�<x�.EC%��ʷ.P��͜,r�Dyq��,�O--E0z����4�V��Vm�9DJ�E��..
��%��*e۴�pCL���[��+Z5�D�>6d�)��1b޷K��BUs��YA�Qi^i�ؓ4�짚�J!�_9*�	�{�J��~�/���&�?uCu�n<�����H��oz�#6s��\�(�0�J,TF�X��62Q���a"��u4Ė��s�Djda�(��뤉En]4Y0�X&������]c"`�E���"LTb�$��\ۤ]܁�(�M" `�2�e��$HI�h���c&�3��c*&ЖL3$d&�d�H.�B�$����i�$n�ؠ�1�U�v�"�ˑ�����А&�"��w4T���-ûth2]�b�"d��(������ΩQ�eDJwp�L�ܢ"�H��u%ݸDA�2	fh�s���cD�@d�!�$��wu���bf�C��!sv��s��1S�a2�ܷO7��
e���F7�4A6�6���aR¶gZ��ĩ<执����	��R�X,�"1m̋z�Gg��ݞQ��T��b>�>��X���C�"E��^�^"�|W�z���v�������������u��m������[�{m�z�KO޽�����ѼmʎD_�����1��Dd>�p>3� �{7ߟ/�?{��W�����o��������/?7Ͽ-~7�n�߿z�ϫ�hޗ��v�u��c{k��j-��W��:�m�ε����/�տ�~ߞ��M�|kĄF���@ }�,[��:�.�������_�'�}׊�Z~u}���Տ��o~_~��~7���o�>������w���yW-��\ޯ�_�ϝoJ�+�����Ǎz��m�|_W���^��5 }%��"4G��Dz�/{#�Oz���ڻ�\<�������H��b$y�uzo���7����[ڿV�_�~��_�zW5~|�y��[�^?x�����5�r�}|�[�o�so������x���w��������m�k�����~��{�}⟯_/>��D/�_��?�;z^ˏz���O?|����ſ�߽��޼���x�����[��V���ϟ}_�~�+ţ�<؊��+��}�y������?��ϾW���;'�5h��Y�(����o�6�3�i��=��=�����D�Ř�|LX��O}}h��ە|_�]{m�x��ܮ�UxUX� ����}�TG���Q�1cy������Ͻ�뵻y��y�G� ��#�>c��LE�>�>(�ת,�>ճ�7�ڽ��b�TO���>��Af4F��ץ���~�o���w�W���9�k���:�_�zX���x�f�d����zݚ�������x������r��y�ן��xޗ����׮���r]�gxWw�Q��>�$DF>�>�_~yzo�ܷ�/>��_�z���v�_��^��޷ﾯM�^7��W�u�Ѿ+��r���h7��^-��[�j���߅R�
�ZDUW���W���!��Z�`���}�>�DG���}G����o��^b����/_�����ߊ����������s^��w�z��7�o��׋}o-�]���]��|[��6�p���e���E�"$}9�.�9Vgq��K-uM׸��@!�
O�{�����>�����^6������m�޷�|�����_[w��o>�^������}W�������/K�����m߿�[�<m��^����{W>��o^|������xF{��h��(��7n䘩1��^��,v�rE'�iVy�`���]2+qr��� n��{�[ĸ	�h;5�ĥtQ�\ܭN���+z�1V��Y��yK�V��vq15�?'ϭI&kﺝd�)%l\�P�r�� ����,P�E9��{�LW�/�_����׮�����~��|�6��o�����ߋE�~�w�U��[w���Ͼsr�׋�����}��M�}k��z���~-���;�+Ưn�����%mk8h>)}�=T3;�=T=p���>���_�*��˛|-���������o=�^5�~����������<�|[�߭�|�E{m�^���/m��.����������H�K�o�H�C�>��#��W�o�r�-���+���ם�*���k��y{{m��+�����z{m�x׿���KO]���������r�v)������o����;4|{��Nވ�� ��*��Qd[���#���޵��߯�齯KF���_��^>+ſ.�*"��m��;cr��9������vN�^I7�����o|��G��}����"0G�(�ڷ�u�T���u�v����}��>C��=��X�>��7�_���/Ž���x����}Z��(|v�|y��xo0���������ٚt�nm����]��ܴW/�:�7�� ��P��C��
�W�B�e��̹K�W�D} }b(}#н�""�}�}��տ�����z�ur������ʿ��~��:���ϭ�V�W7/�y�ֹo���>u��㗦�*���|�ď����#�<���_�nf�|�1z�ߟ/��o��^�毾���ok��_�w�{���}W��_���^-����o��ߊ��Ͼz[ڹo�����*�����������U�\�/�|��~>6�H�,��A}�$|.�`��=�~�@^�����z���7��Z|���zo�ܫ�77���߾k���7��{��ޖ������}W箵��o�{��ޗ�G���_��Z����������_X\�b>���P�]S:��zj�P}��S�^]���N���ᙓ��{���'��h�����{�~�ŧ�z�����o�no�_�5�~/���7����-�\�>�sʌ�1FC~���f>�>�>��$��"�}Pc4�q@���^��(�sY�k��m����������r�������~7���W��[�|^5������/KF����޼�������o�U�_��ߚ��>�m�~��U}\�ͻ�����
�>����-�\ZU�J��w� {71YT�<�A�B�AZ����|#�*�6ҙb�bLխ�V
�mlZW!�(,�;�۬��sR-�5��SՒ�����V���0�ݲܨ�b�C1��;�GqcʴN�X�;��S���gadM��ʗ��.��ג��n����I@Ȣ��x��@��~uk�|y����޾�s~��^?�?+��+�F�m������_�zk��?�^-�x�W����?z�7�}o�+�~-����}o���כ���\��]���n&�6�z��鵢�}�>�"<����~�����y�����x�|�����/?����-<���|���6�=���M�noֿ/�-�]�m�o���^#�>�""���>�>c�����x�U/7֤b�}�����D��=SC�B#���^/�:��W�￞���Z}��&#�������y;,�7���Ǽ�jn�3r�V���}��_�x�����_�����6�"<"�H��>��v�~�V>�����_��O�������m�����x��m�y�ֹ�������v�ץ��yoM��w[�����X�[p��{�祾}���:�_|�񾯭x���~z�{\�}�8F{����D��n��a��n��x����}��sƿ���X������J��oֿ;�=v�m��U���צ޾�5�~y�+�so�>u���}�_��ە|w�=4h�۟�;E�zk�\ ���L}B>������{`]��bO��Q�iz�>�H�a���Nçf�f�d����j�7�zo��Ƹk��?��b��[��������W����צ�/om�k�����r���~z������}O�xE��}�\n[��y�O��#>�&߭���>uz[��ݷ�}�>��5�����_���ֹ��{���׍�x������׋Ƽ|nx�~w_W�x�����?��7�||[�������} }^?}>��X6������I�|���_|���ߟz��x�������}m������W._�>���m�oJ������5��:�~6�y�~^��sn������U��wW�u����.���)8y?ϙ+�HD�p��]}�X���=���k���������|_�F��o^���/j��~�|��7չ��y��X�/w�߾��U���7�y���-�_:�ޛw��G�}��\���b����cu�T\h���">��oM7-���z[���k�\?��T[�����{�o�}k�ڼ��������Z}y��W�zo��^/��|����\����U����_�z�_���U�t���ubJ����Nm#x���˻z�d>s��'���{J=kz�{��O-U��)��K(K{(�w��+�yu�9�S�I�:�v�pu7@����e#��]c���P_��n��C�N�a��S�u��_507��憸�(�pf>SVM����׾�>�������|���KC�k��^��\���>���צ�m�^�o����s����-�]�����E�[���~�V���ֹ}���׍�x���<ѿ�|^�C4�-3Rn�T�=�l̪>��} �>uz_�i��o祼���z^����k�w^�����h����n������m�ν��o������U�r��������zm�}W}����j+������Qk�[�OC�3Ѣ#F�����{�?zom��o���w煣�wu�_^��6�_��^-�ί�_�v��Z�������������o���/m~/�+ƿ�����7չ��������Z|��?o�/bN8�V�j.4}����}�{��ߟ��x�����|�U��x��r���;��<����+�wW��ƍ��[��x׵���|_���y��o_�k������+��l��~z�׽�7/&�~�t}��>���DO���կC_������7�_�O}o�>�������_�翾�ƹ�__��?ݯJ�h~��o|���[�\���~���7���qW��om���~����w��߿/��}R�W�lv/t;�S�� >�>��+�*�����[�¾��ԇ�)
�ʪ���_W�{�����o=z��y~����~_?�І�_!�,��B�u�:�bvR�����a8�Ň02p;��?W�Xd�l�2�\0��T��u:�cuc�H%��]v̚�㡸�$�:� �a��QW5��P_�a1��23�V��%8ݧ��q
@�Zmү�Ky<;{*xݖJ@�@i��|/�{��[{����/6m�X�kRX�T��!���źb:��;"r��e�'���Y����۰d��qt.��z��yo;=��ZR�:�/����7�.IV��*�hU[�̈́l3Wg�;9#a�0�O4�5(�r�Hmk;Y6vaU!;��\º�7}��)�f��8�[�A�5�U���z~:��.e����tƉ=�|)\Â\y�;I��2F��o	�V8{�!4��=�i������c:'+G@�c��ٙw-��[�1�)w��Ƨ���)[��F��F�o�G9�84BO:�Y�?X6ۚ�|���%L�mz��1�y�u���=�q�z;��1��ˋ�@��������<��G=��y0��B:$�= @��ZH����N�#:"���گ�w���ʩ(#(���/8���z]�`�y������q�E��J��ۊ���Y�[�FՋ"���Rx�L��9�1˵Dv��"b�1�M��.;���c��~H��&"Vӣ<R;z�C�M��9�ﻜ��Ϥ8OMF�uJnxP���*�I���L@	�=11@��b�gev˾r�չ^ah?'�`��~?{����%���{� /Zm-Lr<�"K��y3W�{$C���QS�~��{l^F�-5�.$�ь}?95��Qx��DK��*oW���)Ȟ�y���*Ϫ��RXU���a��s��W��A�F�_���Fjt�Z�`�C�#8�[^yW�': �^�ÿ\�j/��!�4J��VBz�u���o�"��iJ��<O]�|�Lo{r����q3'۹M����TJ�۠��`V�޼�T�M�X�:�Ζ�َum��Me�u��9c�K��3�D��.t
t��1��EÂ��f��d��A�� �
���7��h_n:�\���kO�U��F �Ap�T��)�pg��_(�6ޞ1�5�/��|�ՙ��7}m��X�G�U胾�:{�Y;##�j�����MS�h����E�R��=�qV����+�rV�ir�Q�nv֗Nb7�̸
��Y1���˞�s䝃U�t6:i�(���@T�l6E�)���{�q�|�ґU�u�b��������ۖ�Ȧ��1zm�y��9�X�"ns�t%ҠAFϜDe@(A^�Q���q\i���^�t�d9����݄@G&YΧ�	J�܅���'�$�|e?�Hc��n��,X��B���5�y�lQv��NF�1��T����|�PS���[�F��h`�rɽ�û��s=�mK���3F���0�C�BiL�< �>0R���Y����{+V7,��<�����\k�N�9g6s�������G9"z�q�%����/W��ad�m���Bl���^�����T,�"T3����f�W(
�M��:\�cj���`�'��d�:�38�� 嘄��`���v2�u��q��Ӌ%�-��7�.l��TL��%�5҃Ē/x�V6G�S_]JԬ�����.��9��j��	�Q9/���2����ls�tn!9�\6�y�U�?���EdS�[�N�ޕ����|R���x(��_��W��y!�&7�Q����#\��y=wYcfr�m8�ݴ-QM��R �a����:F����~Λ�PW-j��,��v��9������5��&\7:4�����u ���c���X[�漳
��{g�_��cb�'���˚=J� rrp6ꘋ����R�t��K��?��9B���DVSFqp���G+��ˉ뫌�zI}t �&|Њ���oEׇ�AW|��	�=7�޽�0̛l�0f�I�Nv�u{aF��m^����7��1��Tz�S�wFo@����Υ�{�h�A/��J3�����E���a�s���g���n�n�Y��Pn+ɞ�;�r���z��|]
��ex]@3�	%�϶�V�4�K��������~^ZŹ&C+�YΆ�(:z��k���l���⊏��Ґ�S,}R���:�L9ｃ�7t��썉�Tr�eY��]S��{�^W�Q����iqm�;F���.��L��e�2�����kӐK�5yͽ�2��)3��Uz{�K�}���q4���y����ZeY���2����D1��=���	�=F�[C�=|���7�諭���p��g';G(1����[m��M�Άl�c~b &�Ϩ_����d\��[1�;َ�F��D�qGQ���OG9��y��n����U���Lq =�x\�ȧ=N���{�em���!�a�Wj���D���a��N@���f`�������s�ah�p-Z�~�
}b���B]����<+8�B곣�b�_�*Xx{����R�{ʄ�J��:+u���7��si΢�CI6}\���5�}4.+�C�K>?^�>��rՖtOV��e1��:v9]�}�eN���J8�?�\���z��Dh�)��O�|=�T�;6�r�����X�b�O�=�%c2������Q;@�Zl�����1�{�׆-%eF��\['���`�	����61��健�[V,;?	�����MAɱѫrb��j0(O#2g��soA����+��Z�n�U���΀tle���]��+&pB�s����.j����
~u7\2⺗ �|�O����̯!FOV���A�W�{nz���v�MZ�Z�
��-l�}�ݙܻ�.�&4UNB�� a('Y@�l�u��d��S��گ9f�gJVuo���SQ��*�>X�ʙ�me��V��.`� ��#$.��6�a��g�	�W�yF�oE{�63`[;����Ͼ�����ݸ��z:B8L`�;>8���7�v��q��2R�b1��=Y��U�Ë����1j��H���4c����z�xn���
�6�s�}���נ��x�5�� =����掏]���ykʅ����"��b�'�V�#1:*��tX2�%�j��>3ȑV皞طLG\���dN/�ۍ�p�_-�m�]�xܡ&z�8�9K��P
5�bwp�9xTF��Yc�l�ĵLn}9Z:�Xn/3s��ǽ�_nwMes��Y�.:�0��:�=/�r|cD!����ǎ�9��D����nB�V���
���t5w��[��n�5�l��q��E�p�ޱ���V�=.X��.J"O��債��.QGF@?3IO59�#:"�:�����Ӭd�d�]ϯ`e��b�-� a����t���b�g\y{F}1ݟv�����W�2��uT]�.�D�۷4���r���Hi�r���K��h��M>5�qgQ	v�3^�)W�NX\�h���G��`����}�wD��Z�L��(B!�w�qӸ0�v2�_[Z{UI���d��X��m�T���_���^/o�*�V]_P�bs;���{X'YoPS\qt��s��n�|�>ޠ��C�E*,�}\(F�>d��j7�}�F���P�\�����71QѨ�J�ɨM��:`�&V�F-'xYS4�룵�z�Q{�跄6aP_��9�����O�g۠9Ùb�3�U��Wn�����`c��袥��"��
�{����.BN�ȇ��O%@��Cz)��Ԃht����6\|���\	�
�<8*�V��(;�f�9�ێ�ݦg�v�Tp��v)HY�X0Ŷ���^�-���FX8��5bA\ѯ`_YG�� |��J��1������Xm���U��O��=Y�k�S0�g�ܙ��5?dM�M���q}kT�IT�o '�˻�=��*@Ϲ�.MwE�-�SNJ��q��`~B9�{^��t=�r�\����f�[��S7]1%�@2��y����Y|c6��p��f��4C���وv�z��t��u�I�,OPJ��n&�l��CG�z=�gG9>9ߍ�ۖʖ��J��;u�-�Ì�bl��]8�:ʀ xW�s�]��S�T}��\k�Hg��a���B��~;��h��8s��mʹ�.n�k���+5�X��_K���h���E����b�°�&�ׂqq�t�#�%�@�c��>����=���?*}KGpu��v�-��c��a�Յ��{/��3�症��O$�oA/.Ɛ'G,������ө؉l2��cu�5YU����w+� �RxD�IR��k��gD�c{7kf���Wi�*N�3����&/n��Ǜ�yڸ�qRL�w�j;tC��ð�:��@@�r�[����E�Ñ��teֻ�	0��2�I|c�ǖ{�I&�c�p!j˕}���lQ9rfPq��t���k�x᷁ѥz�*��S�&��
�Oe�o���.Q�\;O'Rl�݉����Z��
B�*�4C�nT�=�&IW{��R�>�!N�Xf�F�pg�|��u�R�R�
�л0�gF�3�ae�`���h�9�D��kM�4k��v��N�P�ٛv�>�[[CdҜ]�ء����U/7�dRYS�\�n\.f���n๻#I�IyV�3�s����E�nN�e"#�c�OBTՔ�k�e��'' ��3�D��	y�PݽYg��l-=a��ڬ3Yo��[��N�^��I�i����V�ƺ��?�2������#^a�Q똂�I���L�)�Z��*g����L�>�t�.�9:��@�8h��'�.l��������m�V�V3��-M��]Q@�S>��y
m�# ���!�+���=+ҁ�[|4CKϳ�X%δ4l��
V�1���Jm@ �\�7`V��ӛC��Wβ�<"�%n��+�d�җ^:�p�4l�J��x��LA)��T�ֻ	^K�r��)/�����sw�r�H�0=�v{V���P�y%P���MV����%�Ըp\�������&9�r}Бp�/�!�˭�r]�E��!�ŵ�W��T&K�z�9k��msq�ҷÎ��L �.�:��<-)�ҦQ�S�<��/u�)�K���7h�u�-h.H���X�\��Y���;t|��54Ty�m]@���h�ܻ5�)l?es92���.U��|hk�֕#�QPn5̦)���py[�9�N}�i��FYׇ�^��=ZT�`��Sj�����4ó_`Et�+��q�4u�|�͎3�.3nm$]��z6�%4O1��N21]��U����y��[l�R�\&�[z��4<��"�q��wʔ�(a�Nڶ#��e��G�k�\�*��,V_$萃?���2e�O�ɣ�Jug��5;su/s��H8�Z5;yt��(m���R�Q�;�F������'���Fast�ni�Ep�V"}'��o�������0���3m�v$��{�Ԕ����*]�#���u川;�E��:(��$D���w��MGnVLs��@�cpYgv�{w�Q�s�\����w��& ���O&�.4�ٓO aA�ޱ6�v(���/9N�����{@&�� W� O�PH�,�,�0Xb�I�%�J��,�XP�BL�L�݊III0�M�'wB�F��D� ��" �.��Db# !9�c1L�JbBȖJE���I1�1D�	�@JH����\�	b0�&S4�ܢ�"Y�]�D�#2"�f��.�a0wt@�D(�f"4�p���"),�H`���w]N�q),�)wn��1���DP�D�I���D��J�)0݌����"��0�S��`��t4� �B%	�]۴d#��3$�wW(�d�dd��� �H0�L3$�U��
��37�T�{��H����K�3�.J��K�'���snHcx;�U�pQk��}�r��J�$������W����9��S��a
W�^��H��C��Ę��!!�uT�y�^�����ZS(�ю��mgc��pd���SF3�r0�1���J�X�(�����`�ZH̫�<�]k�*���	ſe��x��'�1AWO��:4�� �uHMB�*k� _�7�i��M^֖r;�c��8��V��~�5��}\�$q����y6��@f��2J�g)�9\���o�]��g03���;v�m��%��&6��[�p��b๶K�� �æc��Y��'/1�(�\�!��L>��Kʼ�4��"�7[�h{��mD��;�&$Ou�)ⱍ���b'c�.;غD�81���9�1��^�lu�^4!����0�"��������ȣ�A���.���U?��a9g[�m�.�[.��u���~ٻ�p�.Ǹ��>�-�;�u���uLE�-t�ϥ�MBs+��D`D�c��	>����3��o,8yS1�0_۳��Ҧ��I�F(v�3��ٝ�,��X�]���z}CKz�mPT�̛αS 5��^{H6u�|s^s9W���K�Z�&��N�nN��i�p�C%G�x;E,����n��%dÉ	�&c�Cr��@1��Y�����<���>�)
�+a)n% 	��V�}�of���D}��VރWWX|T�ۊʭ6ЖpiV�2f���f�Q�p_�k�7���y�9�]���ឤ��̝�� �"���� ������Q>B[G��L�P
�MCQ�S,�wM����\��Jy��K+UI4#*�f�zl4!��(]��4�+W!ǥi��<�/2$���]E��֞�IȪ��q�N�4��q�4j?w�*>Ґ�,}=�@����|�q�g�'��a=Mt;��G�����|h+a������m[��N����zCnq��{.�Y���O�Z����(�@-7z�m�suL��赥n�{)��g���ژ���O�����v6}�W�$�q��2c�n�ˇ4�ȳv���������E*0EzQy�d/���#Je�F3�b���)�f2���f,FҚY���m���U2��M�3!�rG��5�:�"z&3�s�xn^�/��Q��A�e�ޞ���HU��mOEN�;��n��b�˰Z�`l�2�O���];]9_�H�2�]
�Պ�o33Q�x<��Qe��Ҿ�aoH;�e9�H��\k�(�N��GcQ����e��)�q��bXR����x�0�;Q�oQ�97�*f�MǢ�fe���w��J5bP w�}��L��3�d�t��<h8��j�d�Ҿ��ﾇ��9z�86T���~��T�y�2��e�w�ކ��жq��:���/؎'��_^��Z��=BcFS�;�#S�c��WF�c !Q�K���Xv~ظ1��fy���d�Dnk�e�'E��r�6�T�2GL:�b�g6&r3����g%r���r��EW��)���ղ|p�c�C�ꕾn>�Õ�w�����^�JOV�����"Z�KCߡf塋�J����X6k�,�ʃ(ÁdENQ���d��m *7�c!�+�"�dX �p���I�z��xo��bI�aF�V���B�>(W�sXn�P_�W]�i��͎��fÙ��ф���W�L�q�*�t���6�t�Yd��.	�0x�϶T�h�6T���U�w��F�}_Yl�h�S�-��.�1�9_MV�F�g��n�TO��0�}rv�s����e��ɍf�F��q*�]�ONF��Yx�1q-S�9Z:��bn�֨�N�5Zs[�UC4t��u
�eb��
5#Bu*z{�r�p0G�Y�[w��%�DV:H� ���kby3��Uۧ���d����k[f�X	d
3�]�S����0����uFt'�Y��21R6˨�.�:q����i5Xz-����v��<�G'
�b�[����[8��՛�.��@^��ڊh9<Z�p�%pݽ��>�菾⯱�d�(��  p�O31�#�D-��r���˾���M�:�Z�g&��s�AA�w��&�mdKc���;��m�ǅ�����t��v�{���0s[5�Ӄѳ]��F%;������,��x
�-&�)�P���b�_8v�����Z��1TӸ#E4ա�]"b�5�n�n�t�f:��#PvHUt�.(���م�X�� �G-�&�J�b�Z5%P��j� �p�&R�5(���r%e�w�j�[a�r.���8���\S��l��6�l����Ud�����aIc�����ۗ4�e��&��Y���;�L?5�������ww��]����:��N�e��Նҍ��P&�r��qxg�`�����F���9�5u��z���&.�桾��9��b�r��j�
�_^��9n�t������� �w+�U����A�VB\������}P��,�2��0����g�����BP�ߊU�x���g1��-��M�z���~X
�q*��������	���+v�nӦ��W'�i_A.h�M\4:U��7W���L��ZW|�J	r��-��[�mu��o9�%��p�L͡�r�i�d�w�5ҡo�#菾�7];x2�b�	5�/�/�w�\�Y�{� ��5�ɮ跕��d�DQd��W6�V��`=���.��.������q]1	ٗ\�'�L�Qn�c����8vxj3��h�M��?W�6�`W�3 �+ugC�_Llu�c��,���pܶQAs�W[Y��CUQ��b��q�G���A��\¸4��2�.2�LP5��lDk�y3٪na���2FE,��㴚�}�q����$�*-|S`���h^�.l7B;wV�z�'8HK�0\7�эdY�aX"M�R�:���<R���J�S+@�}V�B�Sf�Q�p�|�b}q7��Tzߡݯy�	��5��	�G��� F2W`���r�>aF�S��=�n��8�ظ����E�b+����`���?L)n��NW˲��zi�l8����wm���b�-��[ĵ�Lms�tS1��%xBڜ�@�w��gfQ��9�H����&f���
�0Ċ�i���Zo�N�;s¤�+���h�u�f��P$�۬MRI�4��;�_!�F�+o��]��VZ �TD5��G!7/bNG�(��ޓ�[�c���/+����$ʴ�s��&�mN]��hl�,�':C,�5��X�Z[{ҮH6�3s��/�+=U+��l���#��>�θM����F���f���jhk]"l42<��p�Hз!�\⧦��4��ܝ���]�o��>��wB�e��[,u���Dk��ke�цl	�?TK�� e1��Sk�k�����;cDdܱ�ꘋ���5�Ń��i�vЧXx�t��v<fN7��\��W6�ʞ^[��j]K{��#��_�RoуJ���.vge/��������u���WGp(È',��~t�X"}�p�MQ{�u�\��"1�W�n�:���349Sy��߈�O��׃�GZ_�:	}_���H}8J�i�b9�����k�:�8R��rtFcn��6��w����ixS��q�>v:���%cw�lUV��%��NM|�S�r�����]���4j?w�*>�JC�q:Wq�b13�պz�n_�Ǳ��A���p���[m��I�����_|� M�b�^�Aґkل�ױz��Fբ�/��2ˉ���3��Vr~���~���������4��Y���FnE��6o��'�����4�r���z��&��YX���Ͳ����#�B,�OYf��XAIܭ�0��՚�B(�srZ9��c]�[�wq^���������iأ��#M�*�yG�a�[]���_U}_}����M�dܑ�xtƈ���Wj���D��c��0�iϓ�#j۲1�"6{�r�-l	��ind E�J�&R��iL�E�_b���)�f3�oe#]��.�D��5 �1b>�+R�>��#��=��ux�^��s���?f�����'C�ܻ��س�86�d⁫Cg��-��X��ΓgO�ed[�!�V�Ю4~QX��|]��o1�ћ��'�!����䩒�`kυ}�L'PDpD�!i��&hE�lƜQ�9-Ք�)����1�j�v�����]����7,.M��c�����]UH3<��]nn�:G	Ït�>���kV��Rw����3V�����W��8�>����\6�gX�ܱч�t�]u.'��L��w��)�zb���W2���Y�"r��p�i��y���K�[�4����S�3B�=�����@Tn5��ڪ�������)q�uת���sٶ�~.
?#ۈ�����W��ݧ��`xOx��;R�Ns�G-gֲx�+RÏ���cTx��5�4��R�6�5�J��Y��k�.���F��*1�!�c��C'���B�^Qy�ÖӅ\�X�X�әr���r07��J�Օ�8��Cx�kgP��&�Bv���}�h��(��e%�B`uu�o:d����}�W�U�\��ں0@��dy�w�T�܈�_n����_��S���%+�?XD%��8!K��[���Tj۝K���8��$HؾS�G��[��	����˪�ĝ66'����e�1n�uNv���NL�ifz�����L(�J�/
�?0�Cf�Cӕ���Uf��Ң�5�A&y(�#�[K�x]KTx�qAeou���<}�]�F�s��Ha��l�Եh\6�0M�.K�C60﮼���@�H��f�喙��l��R��hu\�t��k3K��:z��?eC�B|<_҈:(U�]��TuOrݮ+EJ��+k��6���r��Q�,y{�1ZP�N���n�鸁,�1�G�����S�3���v�+�⸦M�Wf�=7����\���ա�]"b�`D�� ߾x�$@f;"�#1�\�[����[�N��!�)�Q��h��BW�ј͈J�ɤ�p/>�E�B���R�)�j/WY��(�Q�D��	9?I�qS���V�Ok�ڨ�K'�4o��ݿI��~�$՝/���!������$���6`�r���� �4�XO#�P��^�*��|�}�� U��[�DR�X9%�j��u�H�.�����F����%������F���lY9V#���:=�7H Y�m� �$9=O2U�t�gOlh��}UU�Iƶ�L����1D��;#
1�n>o��Y�YQ��'���T�i�ɩ����`d�	�����l�vU��*�j�XU���
r�k~ݔ����/�F�t]���h�0`i����#5�ê��*p��Q;����
�����U�S9�����n��6��� 7��:����3�,�^o~����O 	S�>F���ӥA��H&�+F\���\�
��\Oe"8s�����o��5_ӹ�S֠��N{�*Q�z�ܙS�A�Jy+�Y�R�`��Ps>s��x��w�e�ً����ND�ǮxJ�z�V��ޢM"|9��r'�T|�0�:�\it���eaֆ����u��WA�dc"ߗ�1�t��~+�@�W�s�*f5��*`���ʽҦg`V�nZ�O���p��0�{�{g�Vx���Ę��2�f;�K��َUf���75W�N�c.\����4c#\�;p�84�T(�QϠ}��]�YRC:�Ę��^"7��.S�X�K�� ��+Ly�y/����R�I�`,*������}08'+�F�"�^٣�i��<�'/�{Z�.R��c�*ߒ�Q8eݖ���	
��M.�M��Ԋ���s6qSz�u5���0E���~����"6��|���5yȐ!a��5�O�$�Q��t���uÉ�����Bj�S�V�X:M�uE�����A�����?g��ƾ��:H���/k�����\ù���s5����"�H'Ib� ��>����ow��uZa5������*��F��J������f&N���?�>$:�CJ)T��5�uK�x ��jC�s���l���_�U,Ԣ��"��0�=�4[1��Ƴ�AXhd3��ǜ�<�!��lu���`a������k����CN��B,2�`ѱ�:�
'b�v�;���J���u;��w�Nʲ��ݝֆ��ed�|ꘅ�C5�X�t�bFu�7J�� �{���z������z�H�����)#u3#��)��ݵl@�p
�M�0~P�g�s��U{�Q���gݫ�nY�}�ܡ��:Gn*"Ʌ<�G#fb/��jL�(�F5q��2�z�8}S���R["k>��z\@��9�Ä��d���|��H�i�XO]�*����c� ���}�}%t�9'�D�%殙���+��A݆��}u��Z{�㉮̄�S�MNk>����`�P_�*�|Z;15j��u[�l�ZpBmm��!tW���F��'��6u�<��܀�ɚD�"�+m�N�[Ќ�d��K8a��;}k��b���n��̐.�7�)L�{zf�q�p��]-��n}�2�he�]�0b�O$a`w������\ԣ���wAv��D�ސ��lJ5�� ̈�w�/�d|�3��]Ͷ���!�kx�
a;�a�tf�UjVQ�+~V	�{j	���Zl����ַҝa��zef��Me�C}�o�A�w2؆e�{�#H���=ҕ>.����� Wb��̕d՜F��4�㥧��˳�QipC���r�JAvnJ��L-y�쫺��C����l�W�P-;f�2���-^0�9t�e	%q�^S"�[���x�T�c����ơ��r��e��h�
һ�u��k�Q,�S [�ɰ�dW�����+���/\�Ҿ��Q����ْ�;�ev �0�H�2�*��=,fɴن1>�6-��:��M@5T!=H��F��J��}]���&�� �u�-�����e��k����G�t7xG�ֺF��D��<�Y�aۂf���X�صyVy��8���)�^�F��tE{B]�˷+9+J�	�]��Ҹ�v�6�F��Z�]�hv�b3@g[C�̱dhншLE�5S�!�qkU��A`�8���8K�Ev��E�:g�w��A1����5x��Vc/Qu�D�n�Ӗ�������r�{2���b�W-�u>ʗ}��y"ɨ�gH�X�/�h����rj��E���vp*�TR�]�&,]�®(9E��;i���tЃ4�	V�m�����;���mj�x�ϒ�c�,ai�j3�E�����ab�(�~���Sܨ�d%/�Lݵ7�љm'ۇ.�wC.����fͬ�ﶧd瑈�&,U�A��+>N�d7+�\'�G�n�uI<�O�ᇸ�:���E��YO��`iSZ�������'��%{һE���8@�I:7���ϖ�mμ����q6�����t͜��3�
ߍ0[ɯ�9V⁭���>�Ay9F��\���S�$���xX&��9K�LfX��:����������F�v��}�n1�@̠��@������z�[J�BW�$ .u����u�*=ʣ�Y��N�vvn��M*;�p�C������׈��]}.�e��#���Nش�K6�۳��\���UӮ��ܕ9�Y���o�qb��1�J1���ڝYJ�q�)�*�����/���Cf��I�|'%��u��cQ��vm�w�rAS ���f)0Ha�g�h�&��N�5pۑ�ӮuaH�+��ؔ
��4n��LX��M���Yw�J��P	s�����7�#�J��x�r3�<�,�3;6��������u�f��E�  @��  %$l�`H0Y69��#�;���bd�
N�I;���ز���Hܺ%�!�Wdl�c�a+��#\�$� �8`��M `��60�QD�c$!�\�K3 ��E
0$�(d��	��i��Dh� Ib���HBl�BɆcH�JC�0�%0f!I@A`D��(���H�	,��dISLM�B�DD�)��
�Xl���"�HM%B#M
K Ȍ��	����b2"*�DL$�(M0J���L��I2A����LfcI���S$�Y4a���R�!`P��P��t��y�f�wT�y�P"�ͧyk�9NVJ��g�P�Z�t�x�q��G6p�a�K�[)`�Ǵ�Ʈq-i���_}UU[7�l��*'7��?��4{*xF�u��}���_b�ep�
���^�_1Ǜќm?i�l�|�>�UDބ�O�8�������e?8=��Yt�������/�i���쥎�E7�����N���G��Gd2�����:ku���MΎ����Q�V�S�s���,Z�g]&ʂ|������؆8O�y�����)�m�@דܴjn�q�衴�締�����~� �:F �yW�1��Wj���M\M���#v�����ys|����.Jp��'�:�)H#�T�"bR�����_��Êtف��-:V)���q��7Kp��jo���0E6�\C�fEB�(�ʧ�H#�M�Un,6�l�����gubͦm@�~�[H ܵe����Jb~��R�P�-E�:M�,�(h�-�m]x�v�s�����i�m������T�Q�S%�2�������� �Zg�c[ۇ��epoSs5<n)�.�c���Bѩ�6���@�@B��`iy�[V,z�à/�k��1J4��dSz��Gg�6
�{��&vڵ'
\E�G-��:&���ޥK�1��*�d�eU���U%;�D#����;:D�8����%�-�sHT�W�0�j�W�*N�:�op��6NE6i:"�+!�K_zr�3�e��(su�~���""5K]����I+�����a\WV�/���cܜ����@tX�?cճ �L'��0[�ar*�k48Grg/�5�P/�����J߆]S��0���7�G��{�[`�j����吆��:lC�ެ�ѥ�-�i�������B6�{���a���0�K���l�`S*��8u:�cuc���aneN��E@�Y�����eAP��.4�nOj�su���W*�d5i���Sgr�}�}�v��b:����������Q�wk��Y�-�%�����5C�	6"ҝ�m_��K���6�ɶ��f�,6�ۚ�~��X���dV��tz<��"��J�qt�柘Y���������=f\�'"��j2Q���(�q�N��tu���^-Q�]��ou��s���Vj���
X{��7[�2Dp���p�m`�JGO366R?\Bڬg")���s�D�������h`|��Ga�:xc?^���B��r�?� ׍v�Sܷ9>de7�w�W��X垊*����%�W��]E�Q�4�����7NZ��篍�՝��苘���Z���u�̨Q�(�$]+�'�C�����S���%�-��uG8�s��'����͠����>�Ό�--�#�
���,���$��W�UW�<>�F�a8��)���Jj��oJ�']��cwL~�F<�N��k$���W[h^�q[7����0�nB5�T�����ˤLXc&�u�\<wF1ә2�U��Q��Y-���]1�r�Yô�I_�V�j6�*�&�M��:`� ��Y�~�j��J�S}Ԋ�r�?*H]�G��v�Of�b�n�w��ژ��'�4Fɛ�i���j�6����a�IU��u3�
c��#0��v?[�k�,�w�x�\O��3f�P������ڈ�Zήw��èTO�g|B�t��3^Á�9�I�[�ydYY&��2;,���[t�#S��;�k�G��'0��B ����c�Ti5�h��}���`���#�`��r���`�0�B2γ8�s1q�i}��De�H����i��N3��}5\��CN]gs��J�`i)�f"< Us�ȸ�w��읈䫄_<��Krb�h�͗w�:�
A1�^�t�t��ek�o��CF�f\�&��e�ۿ������o0pz�a\b�{J@��Z��]�Ź���9ue��K3�-��F��Bs�^����i8݃l��a���u���]��׼��P:��3nZ�j����:M@�^��������/��kr�����˧Jj�2�Χa�1.�At�������}���~�Ԃ����צԢ�g����Z:���_0�<�?�G����I���M^raeR�mn̜��i�Ee7K5zUC��-� �<�>���s 	t~}��H��1�Nǟ����P�`#�ڸ}�q��P�'��(@�H|n�hC���D�۹SnK�u���{��t����1�ˡ����ʴ.���дBWl�v:�Ic�+U(����pA�@T|L=-!?p�O�&廎]>;�7\8��s mC�BA�B�� �^'�:y]\��㧣�쿡4�����=�j�}����:�Β9����lN�� �������\��V(��=��q���x�N��´����`R~{�z�&f�NIJ�eX�8�������>$?��Ҿ)T��x�^:�|f���v��kΗ��Y��z�3�z��s�<*LT6��6��k�
�#K�qD������,�� �KҤv���H�/�T�? ������e�N�8>�wRDl��}��rgx�������Җ�V��j�X��]���jS���J�8)���'�U�L*7�rC��=G�S�6�j�E�V�hh?#�q�{et��>{��ݕlՔ5KXN!�v��(H\�+@=��]>ɫ���c� Gu8jwk���zЮ�Gʑځg�~�">�>����:�S=��K��u��dw[.VK�:�"�Z�3]�,X:k��(uTȆ�]�cYY�!4��ݷ���D=c���-���Z+�����"Ϯ��$Ϛ�;A.�KOp�e�&�j�M��U��zLt����*����h��g��5�̙�s�[��o�ϥ������72��xo���~SC���K[� ����'�TO��G�j\]��Y�3�U{���}�Ɋ㜦P8�=�T���n����:j C�
:P���b%֗�[���T��w�0�EU��iu�j!������¬7*�摝�׏o]6i*j�ޠ�2jf=��2&����n��Ou؎Ȅ[��&�r�n�vJ�o��ab���F���q�j�9�PـS��ѭP�L�ٖ8�:�C��TG9��c��{�#e����gd1����g+�`�9J@�J~
a���"�mX�9I����;�F�7�s�*�:7v�V2�Y�D���fY��HR��"6�s�1��xW
�g���(��N�Y�x�1S,܉@�e͠M���tY�;�2J�U	�����!��*� ���e�I����:�J��U�~�ꇔ��t/]�Cg��b��M��oUiN�7+Om�w.��=G*�吻\��W=�o
��ṋ�32�q���J��/N�*�����Or���F��+gQ�s"�u�26G�����A�1��:���,����N-u�����������������<�ca�6QrΓgK:��7Xs^5g�w�oՎ�#�~Rw#��Z�C韶9*d�fX��_`�A�w I�}�>��%����e��;պr�a��ݸB+S�c!�WF�c !M�KȀ��L��U�x�;J�K#�ڤ6��)K��E�-���Me��]k���z%v�]��XpW��F��O=�Pۃ���n��=	��u֚�}�'�3�Ι�U�w���A<�H?s~@��:M�����r�H;J_v����ʨ��ڵ)Z���ޱ&{��Z(ÈOy\9�l9ũ�b���]��.�
�|� �.ى��40w=��X1]jNOF�|�*SaKon%vm�{��vX�ǜ���p�)�2譀����넮4�U���K�����6��;,��V'�.S��k��:쨱���Nf��G����pEu_��IM����T�q��9�2Ř`cC���ϼ���D9�kdo۔9@���U1�uǫ0��7��'�&����y��Em����OWrs�*�k!t$����Y�p�f�J`k}_}�G���M������oX<�K��iAU�R��ۇ���m�L�ʩ�6*�FS��3Z���N�B����T�TII�I[�I�q-�|.�W^�N�ő�W����J�;�}�A�Ƥ��3F*C�3т�ݔ�x�'������k�ڇ��C��PS�wLzE}���P��G��q׵	׹9z�9W؟u�Ҹf�nB}���P������#gMN��e�Ct7Rp3�f�;��k���4�����T&���>�r[�k�֌�T0?}aM�V>LvV�ru��u.sɾ�z�śB�3���w�4��I��c�3���s�f��8����znVkNLl�X1�r�@f`��{�rG}�l���T�eN-uq��f�2���� ��pڮ�z��C�i<��vn��c�,�]�V{��{�"���nhFuAn�U��������@Tr��gCO\y�} 4 �)��ұ� �QS�7��C�,���6�����K���Y��H-T�{/i�[�[�JT���s���9Ivvm``���̧�ܫ,^C����SM��zLV�}�D}�MXZ�۫�~M�ܬ|����J�+�^ȕsaζ��u^
H�)�Y츚�x�q3��m`�|Z��}<~S/Y���sy�������z6���n�P%dhHUE�qs�6;c
��HWO$9\ͩ�!�'<��E��B?W$���ò��z�\�DN�j���TalW��{�lb�@ml���:�+iľ�W�{g*�0y�:��/�6�X�*`d��p!R50L�����<�E�Lz��ݖ�}KO�����@l�P~�}'��"��q59p�um�t��՚p�����p�[ж�On�B�O�������3�����Ҋ��]��:.��4Zq��{�}����D\{���bH�˃���K>��b*����U����.�絉��u�V�q��_[cH
�+b.��vv��2�R.!���P��P��!_v.9_ri\C7�٭bрb����}W�υ�fj*��.��N��tU��]+�D#ޖ�������Vvr$��5
V��)z��$���2Y�,:ۈ�n��ʺz�F�}�}]�a�D���\z>�k9U���iC7�[�7!ES#z����+��ב���}}�qS����G����H�!u@�6�Պ�<�~�\��y�1S�Yԟ�{�y��أr��
�a����lՇ�ZD^����?�X��6)��^��5љ<��o�j9&%7�ȟ���l�[�q��^��<����
@j���fvgM�r�q)��p5��tF1��	�K���Y����¦g������F�c��/�k�=x�m|�Sǐ�V�d�Mvޑ��p����ʾ/�:[�O.u�2�%�D��Bd�vjS�r�<p��gD����ƻ��:_b����_p���z]Z�pߩ'zL��� 8���/{�Y��:���G1�E\� �p�v*�����Mڝ�p�tL.����æ���o9}�gj�A����F>��N��w+q�nqk�҄�K�q��j���o�%��7��g��,RӢE�͛\(}�u$�������"���ꗨE0������I��Y<{N�=�W8�$��	�ި6VP4�I���o��2�K���u��J��uΌV6�. |xŝKl	X��+�uob�U�j$����#c��Tϗ-�{��}_Wǥv72��큸Fg�v�����5v㱶���/e��+0WV[���$S��:b}��K�+�:�KMAI��8kn��DŚ�Wf�j����S�xӇ)�_�?���=g�RH��Y<Əy�]�%4�!����T�Pj��q�V�ʇ(eAq��|=`H�j���9��g-��je�릥u(4z�Ŧ�Բ�	�{Y�B�|4}9�.$\��^���mM���p�u�>;\��o�A�
ᛉT������sXSY��r���o(�V�=�o��[kE�C}SQ�0��ȘN��%��jq��y>q8�6$&
U.One��{[�:5=w�����6�_w\�Eӛ��A��L�U�!�޷�gʻ_}������]�˞��qS3��v���fWG60���'[;p޹�^}��uC3�ԯ��S�m�ozUPޱ1����J�u�S��2��}w��Ay3Kq$ﲆ<0V��[�x���^�y�IvJ^�~xp�(�\R�1�b��a�]��_��^�u��l��\�Oe���V(��XC��K�Zc�U�ģ�'�cf��T8V�D�V�X7����ᘑ�mX�/���GE��@h�S2��U��u-������df9ʺu���5��&֧�}�G�����hඹ�9�3xJ��On�x�x� ͂������
u7)�ܤඓ�ݨwi鼧0�!0X������h^D&����C|�-��-�,]D1��l�U�-�D ]�۹�X�@�R���oLW4����E;�MX�gs�=�i�Ќ��:��j����%fU>\��p��������;����,..��M���m�u��(a��Pl4��F��3�d<^��)��,�8�A�Ql�xK2;��3Tv���MJ�Hřǳ����=��@��#��#��Jy��L]�f�z36��e���-gnK�*ݹS��4�ChE$Y�Ι`qn�+f,��n�~�҂ E�x�݋D�s�/M��+�-$�=�f��2z���z�Ús{B�������7*lcLT�ۅ��.���.5KI*�RD3t�vUk��z[	3�^^�� pV�*�C:���ɲ1��T!���M�HK�����EmF��W-Ʋ�9y)�GH���������,�X�.���S�>�+�j�V6n>Ҟ�h�"�a���2�۟v�l��T)� di�ҔK�CtF���f�h��&6e�����BbN��ݗ�+�U�t#�
�Gz�S�w�e�3}�m�.d�صv.�]��bA�:�ŉ������i��)gtK���<�g\��W�})0��ӝ]��^�>�ڇ%fqQ�}�v`�@�ܸv݆�Q�������V�
Uھ2�ҕֲ���/R�C֡�7P����̓r�J3�����^kƍŸ���<52�'���A���+���U���K��7�S)`���v��K���mNj��<�Z��g+1�_��gQ�����Ln����L�o�� �5�i��'s�X�qB6Џ�v�0�+z�33���mY2�Z��3�$��������>Ιz���\D2���nY"b�gR�̽�{9�h1Sc.�zکxw\1�^=�I��m�V�Uw0C5�Rw\ﻥj���8��IlC;����\���$I�|70�m��"�g�X`�(mrR<�M`W�ޗ�eGW��sa�g[�	�0��V�9���÷p�!����mۏaJ�\���k�� ��*v^K���]�vX4%�vL{y��˟`X�^.��U��Z�:�6lM��z�{hh�����c!Q<B��6�_F�훵z�C [Z�\�(1vw$���%N��-Ƹ�1qV��gB�0�C:��.�˳�m�j�#�3�����,K�̷ҁ�
P>�)�3DQ�PJR��hd�$�d���
�LcFJD���Je�� bHQI�$M)DFC�H"����d3,f2P"���e��F �LL�4�0��	4PR�`�A1H�H�!$��$HH	c$��1!&i(f�D���D��1�,lH���e���4%,J)��d�1`�&�K&�1$Q��Iɤ�DbĐ��CE�3L��@ e% X�(4%��F$���4B�d�c �$��Ĕ��()#w������z4
��}# �����֟2*�2�3
b]�t� ��N�W+�s/6�&�^gR�L�NG4n	�u���R�+���&QN[ �D��ێk#]����sa���ҮN_gq�B}W]�9p��n���N[N�L�c!֮������j��bo[r�4)��7o��=X����ʓ���¢o�f�&��Koo�]�m�dgn�*�!�4��ͭ�A�PM�Q�@򨞞��	^�j�b���)��/�\��2���+f�i���p���=����D>�PRĩ\io1�W�֣���vz^ƴ����1���
{{od�!�!'��E�©
D��*���ְkZ0��?��Z�,w���U���y��'���$�Ҵem<�c�~B����B}{����6�x�W�R����#^)H��{Dk��$7���w�8���!}щ��P���o�[c5�3�!/����!1wlosQ'TB�0_l���⨌\w�IC/��hl&�y�j��;��,���%���Wv��c]f1�G�����@լ���y\�g[�I��ϵ/���ԏ�{e2���m��)A�j�v�kv\�pÊ�e-�E�"��Va�iVV�比�;F�U�y��N[X��;]º�EC˘��}_67�����'�ŗP*�7<�j�������9M�}ujuO�D�w77YS;C*'X�x��-g�'��f���i���<����Jm�t��Qmc�"�ˆ���n5�S��Ș�:E����OfWӋ]opa��m���/��ֈ��s�o)ֵÚ���s�k�u�t�-u�n�+�fu�ʼ��Z۹�������p��^���_����'�k��nUQ��̋�Cj��#e��F�gR3�V������2�w�z�7�\s��}���ۙ���r����N�a������m��ð(ؾHTt��ϥ���ݙ����ó������6_/^�9�����㪾�P��\,��r��ٵp��ȴg�#hD{��V��k(?U�k�F҂�.s��T���W�D�CPqnˆ��i������H���|�q4i�Yvx�%w����xy��J/[�BS,��`X�B�w6#R�u���Wu��|t��)C5�n� [��x�gK��]|�8b8����*�ny�y��q9W� �dJ�I�{e�䗚BO�*f��x�֟H�E/.��Jjz.Y�ǔ-��:v1����}O4۱�.s�|�ʯ�S�Z�ۍp�_��m6��kE�`v�ȧ�o�q��b�uR��7�0/_<WE�KzjO/�5ٮ3i��R�[y�� <�U|�
z$k��!�Q��աz�1>!��
�n7�3l�1V"���ǜ95=S�H�
p��Gw�d�P��0,�\r��IcV#��{��C#	������P�D.����S˷c��d�\_j|3c'R���
&Z|�|�l;��&�Ҏ�@<�XZ�RD�hݘn��$�n��)����52����bj!7�\dk�'�فkf����Ol���.I~��xOw��Zk��7��̇����P�UF�!��ha�z&4dQ��ƨހ�W:��{2�y���{_nV;�r�k�:���8�\\"#)�ͫlsb�TMoU�.+���So�X/";SYy�>����=*�54�n��r��s�?Yb�gD��~���s8��h��Sxt�5���bZ��~��'�4����O�-C[]k�U5>K��S�Gj�U�Y4�S���e�y$��C:��	��K]n'��+H��\ܭ-o*g9t�l.;��\��ŶR��|=�==3g^_��_C��_;F�3��{|Y���z��/�S�WO��������a�qe42%���[��*�syU�;Ŝ9ġ�붓O_R����3�*alW4�r����Q�gj��Ǘ*z��oὸ�;/�$��S�`^ծ��.��lW֡�m�/V�7��{���+݇�]�$���ց�9ʁ�h�T�2�)][ˌp�^8[P�{q<q�r+��3\��d�7�#7@L��"����)i	;q���Tr��e+\w+�B�qfH�Czr�R�:c�}0T
z��RC��f=�<��Zgd�o\WFMs�;}���6-.����KE�MgN�uمkl)���Ջ\|SJٽK�	�z���+g��ܚյnpor�Q]7�.%�۟"�F>;\��o�P���R��Q܈��M̪�Z��zl���q9[��柆���~���]Nn��j�h�Ӯ�9YB]������h��ɻ��ۺ�Q6�ؒDm��[�J�y觬�=���i9�r�qL%�%F.��X�U3�XWk�7[�-����E�@[��@�D41s�V�nH%�'T���m���ru�t�T�L5�.1¸cl��u��8B��P�
\*Hp�s�=��J�Ü�um}��mT��
O���w�ݢ�-�3�,��dL%�-m@�Q������Ȧ���򶲭+�'���dQ�pڅ5)N�'�Q��ֱ��~�������{/U-;���6�"�ѽ�� �r�}�oj.Sti�/�D�]�=Eb��|[�N�:�s�U��P�총��lc�]'[��:���!wJ�9bn�xyvnr��fq��������]x\O��3*M��[zW^k{�"��qac՚�=ä�Е�UD��P���F�F4��So�owTݽG�O-:�dA�l�����v����ė��҂�+b0����nqj��NcSݯvd�U�M.-<�7�B�rGV�=8��F�-l����y6������j����=z��� P�::3��Z!U���V7���[xVP��q[ŉ2]TT�����&�n�c+�3N����p�c�i���g�b�B�i|��Uͅ�e,�yO�%��Z��?1�n���{��7���N8)k�]�P�fJ����\ٮ; 1���~^�Dk���s�����?��O���ǵ�Ν��ݞWsecn�\�Ƌ}������9_9J��}�|	�N3����y#ƪcZ(c��9Չ�_�[I�՜�h����9d;ݩ	�\���ȍ�{Rx��=c�H�b[5���X�1qʎM+e�w�'�U���ϔo�(�8t���� �F���O.ھ��Z;Is�3N�]hb��w�{�*��c���c��T�y��|:�
ܚ��{W�n�B_ag@Z*�����mT��9�m�>���Ddr?[Qۯ��6I����5j�q�=Bs)��T�ߒu�\9��1�yU����&�l7��U<��~�h#��}�U켿�[ܛ{�_\bq�f�_Cܪ�Wf�Jؙܬ7�N�p�B��86�gW�ok�/v���i�^3�7�_:�U��J���b�v˕+�^u����4K�4�5�Y�l+V9��ZE���8o{��I,[~��3�p桾��#k���wab�6���ͼ��u�f#��dt�X�<���v:=�	r5!�VE�>h���.F3��)�q��o�JN�ha�2Aף2���ʦ�*Jc�0����-6"M���4�4O��9��~2��?E'�L�u��&:=j��הt��ݣ��e6�GZ�(����W5bk&��܊m������L^�ʤ�v��/��u|-f��Ǫ�e���9*W���E�k/���}��ToT�1�Q���9X��2�{f��>7v��`^G�H�LJ{���Yx�m|�{fڨ;V�G�.U�9��9��
���PF�#;��t]D��4�~�vk�ڈy��N�,��y���gP��Pو_'0W�h��fB9Չ��to�����t�H�ͽ�	(�,�q͌E��
c�Jb▊�j�u}��(R)��sY[|�o�3}�>pT&�)�3��R��O.�۔ }*�v�j��A��.Ӎ��7�����B�'�v<�u�x�0�xL�Jg�ϻ���ҥλ[wl����N�y�r�߅s�}ث�OZqx|��(a�-2cD�����~�m��͉O�X��k�(w2Gm�}b�96r�x�X�bAv�ٮWn�r���X\��{uH�9)p�������"�s�㾐��I](�@oK�o���tje�}S\�I��pF�#�΂�J5/5�S������ÕA��<���)��{sf8S_6�mCYTU��ddvS��\�R�2C����pf*��ykގ��X���s��};�.�^�(ݬ:%Ÿ� �ۆ���'*/ھ#��[�쇼,QLdn������.$����9����v��xfWت&�*$��n��Ò�ػZ�|�qeԮ�ldK�֚޸�YVr��ʂ�`�5�p0F�|��w<��''�z���#
b�9��æ��v��ުγ��to ��f><�tV�^ԝ��p��+��+�P�\6�\K����Sκo3'w-�ㆢyP�m� ���΢OuD�2�)*W�����Yx�n�')����F�BWQ��J�1����ʾ��]uR��)<ќ���5,AEN2��lM`�W2mͭ��i/{�E�`���j��ep�S�#�b#-7/���1��8;��	�v����-�5���I���Lv�)sj�^uw�ի�"��S�byV���EƬ��)�x��q����7N��;x��Rҷ�7��������E-:{��E��Iw�k;��`��*��9��t����i�t�98ͧ��C�g�B�ﻦ �`���Ue��FI�}�aX+{y��:�w\Ҹf�,��D&�T9fQ
c�$�j�]�T���uI��=����6���j9�V��;A[7
Qo.au��nn�k��Z�`~�
o֍�3�kM7=��.�����&����6c����[z�ez�t^%j��W�qq���Su<}�j�����!����5B�.�%����F�#����_T�Ë^��~ܠ�j�q7}2]����Mg�����Oj��f�X�o�b6�]�V6*Me]k�����nj�);S/n!'�F�Osi]����)��(.:��'���p���R���x���_g�s�yy��$s@� ���^��*��8����Xr
� t��*ӑ���ۄ��c��g1ץ�����	<D�P�x*ᩃ\[o�d�R�6M���(���J�83���q���j�V���I7�Z7��B�W+t*Ay7��� � �P,�@^��m�X��l�L�-.n��Ίn�uN���D�߆Fl�IP��¢�&T�A�-��]��:�G ��v��
bf���e�p����=S��2���4�90W]T!��1$��*W�����:�Sl���g�9�>���y��c�"�ʄNI��u��M[�p�^6����T
<��������nT��pE�y�s����/��.on5�Z�,眶��B�O|�J�dV	 �>���Ҋ��E�]p��ܷƋ}����5�7�9J$ �c���*.i���N�v#��7�̄s�#��V���o�TE�5�Ti����g��{ld��{�/�����nus�.7��6_�Ǝ�˃2\ۮ�A�#��7�Q�Pg�� h{���7<�"�6��Cڽ��KnZ{�Xn1�p�'�̀S���
�N��k���4q��s��e�F�m��z�U���HinaUi.r-���|����Y!����ԫOQJ
��)ǣ��hW�T�*nqƨ�B��83f�aW��qK2�d=�{G#Ȝ9�ր��y�ltMf�"R�H��:֋㻆��o|�N�I��mc�-����^Zã��Q�n\�W�XNck9�%���W�9f�`=�g|��� H�3W ��{|X�;D��f�k&H��h�u<�]<�R��{6�1���j�z8ܱ�L���F�,�:qm1[��\+'��U�(U��wh���\���R�soM��� A�̢���f�ol}Kv�[��lB
�9�/n�kg!إ2�[�Z�))��՝]�,���y��k�6�ƕ�����R���!s�*������^,�� �ڱ�E���lm�ߊt�����\�"ޱ���j&�ި��+��� �
d�.VJ�;VqJo/��:�T�uH�ǂ�ۢH���8S�/a�ރ(���eL��]lD�t��0�(�˸ے�)��VJ}3����mC��Z��@&�'��KrY���|�������rH��~L=3��������+3B���R�]�,D�o�ʾ�k�+l��ܢ/:���`�F��WG�X���Z{���j�h�� �Jy��G]����Ձn�4�44�u\h�q�%7cU\��*��/����`�Ѕe��=��a�.a����c�,����4�M��:*cu(雜���^W�B�醓�ȩC�7��]�7�b��Z�ү��}��"����xi�֙]�+;�����ӹ|�yz����6P�`�J�]ή��!�xd��&h�Qr�s�v�cSg���ۓh(�"��3m��T��Bl�=�f�.?��n���93#����n�W"����8:��ͨ	�Z"��U�-a:m��`�Pk�AbX�Yp;ȨR鳳��6�x�����ʅ��ZP*�w'S �7Z�+[��v:+�ټ�p�R�?�0� ��wZ
��ҏ,��.��Vwt��������3*B�b蹶�1]�P�r��ِ��tkFV���:Z�+j�(Cf�
܎�+�!}l�:l�)���dΫR��V����e�Ϝ]�WR��h�$�D.5�gne�e �7��D���� Ѡ�s�h�k��:A+�	�S��{�}Z�����I!���A�.�9<b�k�7.�-7j��h�t� �iH8"T�;aSP kzJ�G����9�cnۓY�sLR��siV�î�K�/��x�]<}�ԧb��r�M�N�j(#W�q�N�G5��|<�ʽ�dT�7�]�,Ei5��4�=�:v��ұ��gi���K�����nS����ѕ*ъ��6�eз��Q�jm62�r�h9n���p>9��̜]=;�"��������azEs�B��9-rӹ�$]9�a�7#��y+3��O��`���8�卓�y����z�������<{��&`f$�P@�̳a�F	E�����RA"`�d4��Dl��@�b4�E$��"d"�f�E�M1$03
!3&��P!�1�f�&�,�$�"P�f���HQh��
E0�KI��Q$j�0�&D�`3*%,�f2	I Њ,B	d�&1�!�b����4��I��,�JL%�4`��	MbM	�X���1,�(
iQ@bQ�LȢ��	�
��J)KI�I�%2lFK%FJ �~���@Xg� �n��\F`}��Qj���[�H�lPr�ܒv�lV=Ը��R�+r��^m�7D9"�Iq����%��`��kz�U59���q���dO!�ka���J1hbu�.�x-V���YѪ�\$���E�V���ux��o�����t���)/��8뀱�OfTO-���r��9}q��5����˴c��dF}��):Q���^�}�_L�m��X2�TLe��L�g!�k2:�4�����_F���ݧ�z��޿_uͯ8�p��j�J�.K�A.,���Wϳ%��M�f�����sΨ�ï��1��.��t���}���県��_%���0�;¡���So�%�m����:|�<�{�W������+��ޥj9m�-n�Q�Ҹ�ط_6�\��AY���e�x�A�:������2f��m}'uuQ[��GSy�[�p����͵$�Z9��]���\�)D�q�OǠ��01$��t]D���O/�y��d������"4XDP���"o����u�hBjPD�c�O�]q�u��!�H��+��;����j-sC��T������JLz(����$�u/��Z�p�KzFc��t�\���i�bo,����2I��dk��lzjU�a��6r�0�W��A�S��ݡ�6{�>G:�>4[�cjhj(=��9n^����W�Q�B�*
Z+᫞b9���7�-�L�-+�,�D˄�v��x��E|�D.��@�J����Z�|}�8��R��Ø�u1qϜ�ɾ�����(���sY|��B��^�h��-��V֚n$�|�T�rLMD&�\+�rA<k��g=�R�_Jn��˛���A���w���KuM�IԬp���n�����)���_.3(Uk��D���ojgT���^�w=�ܬw�_^�,�LOw�g2[Ђ�W���{�/���ӮS�K����Q+v���P��q9��Z��pJ�J��m�Y�s��ôo�.���_M�O�B��S�DE�k�A�����zx���ϥ���o}�:�2��s�TW(xx��6�%&�P��JZ����PJ�
�etx�ۏIu9@�gE]�PM#�Go3�g�O���(�ź�>��
����̕z�DpGk. ;�����ի/Mi����bu���l|�Ѿ\����K�#�H�����^��lԦb��I��r�g����}�S�	���[·1Cz�3���)lY^9�_���m;k�8մ~���eHij�-��e�������h��f�>�\U���8��r��-~=t�-�F8k:&.���+y��W�5n�E�����{��Ls� �!�!.���-3�v�������pd�?��[=^q��JU���>
($�IK��
z��z��gk~��G}�yxo�>�
�jqx�nQ�D)��������+q����4����vW���4'��֤�=�I��Y@+�h>�r�L�]�iG>pN�!c�|�>E���k�4���x��n�w=�q�;�9�\	.8�� Ul=s�k��;�����ꚎI��.]����9��(Ԃ��1:�Ș���n@+aՕ��9�j�V��y{�S�>'��B�,�v���7ٕjʍ��B��˪����-��l;��싍tEޓ.�՛BPn����ӝ��J��ș����m��p7)�Gl��i!'�<��gjx�����oy�S��V���?u����p�]|�N�[��l�M��h6����+�Q:�h���C�B�{Ξo��^7;S�29�����������إ�L[;{o��2:�ܸ�:Ͷ�r�]�N8Oj����;E����sI�fp��ՓKN���捸��u��%��$��#z��$R��eD����I�nu����fTM�TD�c;Tw�m;�L�`�[�'Y���Z����$�ԟA�Wh�t}j�r��ʉ*^�3j�b���О���G��_��a[�~��[U����.A�Q���uBW�i��a���Ə���Nr�E�s=�^�<��P+)�;%��<�s�}5u��[0��s�=C�n��+Κ'��y�ㆳz����ޯ����A��}�7��-�X�nsm��w8{�=Q<��jOo�p��=i�-�iT@���>�hP�Y��I�M0�W��n�-���X��o�D�.#�5�ۘ�<"��k��QLdq�ov9��)n�!�3fgʞ��lEuu�#�~���ww�,�ߕ�/��nl�w�BŶv�֒�u�)��kr4;1՗Y/Ŧ���4���G�O�=�+,��-g;`z��TUr��5ݳ>":�����GՖ��ā���S�#=�$#j 5��o5��Tb}��m&+Vw���'����p�o�{���$�p噎!Lw�O�A<�j'W=�k��M,��c�)�����P�a��<�M��,�,��h���5˶��8�ڨ������|�'�Y2�O��o����c�Q�P�Cd�ܕ�=��3�p��ʥ���I�5�N[���U4���������dO!��Σ�ͪ�������7���v�$��%�b�=���jځ��V�4F=��%�A���86P�9�39���S�m���n<��<�^'�F�f5�wW9g�s�6�ʨ��
��b�
R3D�ڒ�e����iڙz�fu[�gGMQ�m�v0�S��6�f��a��}C��o/�1޽uPuͧ���9X��<ռ9<�M��(�T�L������o���j�?g�������0��r����I^�5��E�α+/nF�D�`�Z�ɋ�+���� ��"̭79,s���J��
�n���^AKd$Ր��
p�;�fH	��u�k�Ml������=ȵ���ʄ�0��F�a�*崫�-H�����('-�I����h�U��Q�7���}�o:b��U!k(?z]��.��Gew��#��=Ru�mt���-��p�6ި��
����s�7̶'H�k�zLy����%^�/�6��D�Q�i��p�_��m|�z
==3�����G��Zn��ek�6W 䯻�cI%tYoN�ZyqͭcbB���ͲjeE�1��ӈ������u[~���\��`}�"�
�؟z�Wf��\1���d����)|��,��5,�!�#�K����ae\�ˈ�M4��f�,�=�P�ʇL�!qK h���ȼdl��Hm���-����sÛ��|r���7��m�!J�����Y��5:�"��	X���NDM�Mn�L�����&)7��Z�g^ۙ����>��\*Hp�q���������~�jOnN�L�J��žq&�;��>K�I@�wZ.��șC��B���%�Vn8W�RyYن]�B++������&�7k�����՛��4;F�J��ek{��}Y�O�����3���+{&Z��^���/�("i!(F�P�N�w��Snx]-��UOY
����D}v�[��7�UdS��ϋ2Ớ�I;ޫ��gv֟U?+��f+F��Sޟ\�����oK���3x;���淍'�eh��	�&K��'�k����_;F��~+�=��ez!����"jޓ�̾��z�{TW��θ���Q�v���Y�蘙�ح������-�Jݜpʉ���K�����c�l(t�ܮݸ���<Ti˚�`�7ey��������G���C�-����@�?z�b�)�7�d�a��J��=Ce����vw.��㩗��Ur� ��5=�'"�����s��
u�˗c�y3��k^߫sT5'P6&HG:�+sˁ$8�����5������1��0�_O�S�OΓ�|����N�Usr��X�%>4[��o�8��n�*9j����{2s��d�S����v�Bks�>Y��;yh�7V�^)YD��m`�J��-	m��9ޠo�w[d|�&�Y�D�AiX�1m|qܿi\DS2��s4�Wvr�٪����7e˾7�h��F9!�k���s8i�3���<��3��@��{8	�DuQ��Df��Y�˸&���=����[y(Va�C6����ӊ�#:3��A���S���B*b-iʍM�e�p�	!��뜷.�%�2��)E�q������.ڿ�����)k�n0JwU�Fm��^�fl�Te�l�c�"aM�N�,?W��B.��uW8���d�a]��J9�U5�Ʀ�q�ϵ�EnT}R�
ڨ��%��C�tNg��d��9�g�^�t�{�~^ �[_YA��z,��s5�֣R�#q����QZ?ror^��N9�r7���*�U�I��l��L�{t ��n3/�O*$�2�TLe��!L�Ž	�m�a���؝1��st�z�e>d�j�߃9��0Gvy������9/jm��Q��|���'r�8�U=3o���%�t�"�ΆC㺶W��`�Eq�Aj7���f-9�vߗw{�æ�M��;w����Q,��X	�f[ ��}'N`�SI��W��sY]ZԤz����r��$��`5�f=���c��a��?�)�D�
�s��-كPs��s�ƚ|��Ŭ�C��q��_e�j�=!y�m������fڎ>���y�>^+>h���oi���sPu��l�X�ʺ��[PL�q�R��Kun����i���z�N��_Vu*� ��: �l���S�FEX��}=�w��p�X�p�-���B�[��~��)�*b�����C�^z��7۽/��������v}�mC�sRz�.;�ڪ� ���P�_'%���fB9��Po��F��c(8����u��n;��d�|�څ �����?=�:��@Y���]-������bs9ն�س|��v!P��r�|�ـ{�`'��˳�̝�2�j��kPr�KONW���p�q\J�'�C`:\fw�5��B|�K�;��|���5�?-Q��o�y�͸�pLF�"b9�i��ϳ#2o���w��s���3�ҔڍU��'U)m@��z��4EMj�����|�3���9+	�L	nh�\r�+s&��N�B
.�V��>!-���I�u��)ŧ#&�Lة}��8��5��N�K��O���
�E�q*��L��%�.��P�o��s��:�>��[�qO2�M=�v8��ͱ(o>�s�}G�,r�u�39���f{7���&��׉��r�'�N���c�g��.l5:�����J/ت��q���-��Ȟ�y��*5c�Ě������[Qr�d��_vЇ>�K�N�Kt_&��']��k+��Q0�=U�-6:��3��L�?s��~��4Մ���)�'�囧]g+�1��Q�nu2�;�8��0�+�n�[zV�l,齳�XK�j���He�Z������p�1:W[��m-Kz''���B��k;��E�	�S�r���Α�ֶa�g��ˈ�e�8[�^N��`]�F$Į�5[7�C�����Pi.WEԷ��O ����֠�i��j(����q�O8�B��0j��j�(Г��6{�n7>�仜ż��&OZn>�O6������_���UD���1wSg᧋e�\���z�g�ݎ��Y2�1.�����իܥ*��v��m\��e�Ӏ���q�glVԓJ	�6睷�%�'@p411H7�hH�8�Տ�oM*�:.��u.x�]Ԓ"��SJ��;���l����j�����^�Ž�t�"/�y�*����Ū#k�A���.�Tc;��U�.����췋6��$�l9�H�s��gA�����9�9�g]:��옎���n,oN��q�ԙ5����J�u�:�R\u�eI�/��k��%#�.k6��h�U��:P��%�(��h��v9�w������=߂��7a�0� �U�ӷ����.��G�� ���A��n�q3s��$ G5��w*w����uXk����y���p�WC��v�8��W`�6"ٱn�#�[��z`:;�'׫��o���]mbl]l�Ն�i�D=��T�l��ScВD����"��
�L�ԫ@�;a�*���K���2��R��5���u��\�)�s6���&�F��-]�s��B�3/}�+���W�b�~��W����C�ڍbb�pU�]�ċb���e&�5¸���Y��c!�C(㭱wF��r.x�׻�LٝV�Ҩ��v�0�[;9�Ы�8��O1w��(��8ws	��A��}V|wB"Ft���}\���\׌�9J��@#�B_F��+�œ���a�F��]�CW3�:}fj٬5�&．��B��,M!sĦT��N��ʾ���MZT���[@�2e�9C�Y��-�Li�W���*�%�j���B�et�W'���%��4���k0��1'K%
��M��+9$/��Sm9�KZ蕎[9q�x�xt%K�Ku����aL�����}M���"]���r� ۜe[{���xԕ����YOJΐ1o�syw)d9�D�V��%�YJ��u0u�0T}*f�mIu3��[�	b��
&w��.03R�
�_c�,v&�
�T�Q���W"�f
e�	�)	��*�뫧���r�}�d�uv�(�\�flI1�j�Tnb��$���T��u���c��KN����FG��#Cq�=��h�>8薹�㯭Ͱ+�{��>�N��%u�����[ImI�;$��0��l�əЅ��]}DBe�����ƅ��4�.�VS��tb�B�^΃!:z\��i��\ѻ[�:�Ӕ�2��:���շݫJ���*5ֵ��#V�����&�\�+v���R.�M�m�,�X�;L-I}|ﭙ�22��w:�`
�ZwҜ�l�m*孑}�]Ѕ:O�,=ƹӝ�����9Smu��	дKŶ�*��;k�KvI�l�������M�!#�XR�k��%Zz)8<�޼��,�����Lƣ��������묦����ENՑsJ��֦�kr�Wa��Ty��ֻǙ���3xa*L]�J��wY4��� 
� ԂRP�Y*	2c&a�lJ��� �I�a/�F�Nk�b�FiNV�r��Ėe���&ѝ��F2cE��*"B@������(�"�!�R1c&Ƣ�H`�BC)2bH�����	A�����#""�IFɮ\�t�QA-�$QD�A�ѱ�b���X��(�PgunlWwF���1P*D�I	��Q�їw,�61;�����黻A�1$EA��#Asw���mt�*�Z�o~��i�U���SۛzbvB;y0B:�����w��9�cgm:�:�f��`�&]E(K}I�)�M"���W�{k�[�ׁQC�	��L�"�Ғ�����{�.�TmQ������׹��|r��|�h+g!J������-�޼�Q����`�c�N}7�5��2����b�q�d6�;'B�H��[�2���7�%k*���h���?-)w?�On-�aQ(���#T+�2_��mCyU��"c����Uχ��Qy�qj��w�ȃ�}���������C+�yU�Щ�0/�|3M���Äb�y�=Uַl5���ഗ8ܤ��ۄ�5���S�m;F먜���@'I0#�s3�Q߼�8����T��W�/�}�M����!<��]�FU��*�o,ɪ;�\s�J�!,g:����*^|��i�p�+�:[O[�ܖػ�D��uV�ӭ���fAѪ���P�z�T��1������xW����	������k���ݕGR�l�{�pQJ�#Ev���W/�Sk$c��˱�WC.\�7FjV��[�r���	ҋ�td��[��&̙��f���9�-$���F����gPZNm�'>��ۂMX�i<�$ދ��O:�Sl��DׁY_4Fg��ߍXOk����7��T�s�N����Nc�f5��{f�����(0=������z����36l}�j���^�a&���[oB�yة-�C��}0Td+���� V*Z7�m=�X���u��2���Tr�ې�f��r���Ad�i��;�RV*��
��6�ɪ`����Ȟ�ׁP�.��{��y���4�On>��L�QD��2ToL=����P]��9Z�V����z`B�elgq{#�����ǂ;�󍰵�}˶�;��h�͑��$�˗r�6��Y��̸�pD�
@1�2`t�[���Z�҅�Wo`�ۺo�]�%�kz���M,jk��k�r5���nC��6�U�=T%�m�,�U�o�u_F*θ���sP��O*�ٽc��̋��2.ᾛ��mo%p�X��s�!6S��y9���>=�3E9x��<�WY��&ڙ�;��j�X�2��YL��֝�.Kgk�p�Fm*g���Բ�A�:��z8@D�O9P⺏��pWM=��t�-L�&ܢ�S���ug�^v��B�igi}g.�عtX����8v{\��{��yh��5:ܧ̼�I�5�k��of,�[8�cLZ�I�qV�t�p�fQ}03'�K+�<�\Gj��iڙl_�ޮȱ�(� ��Z�}�-ڵz�.��1wPU�{����DIo�0�����q&�L:�\�*�ۥ�I7ف�/r����5M�/^�V&�㊎m{�u��#y�{ؚ�j�����o%��n7{�G2)���ƑXr�-����t��NWDin��W&�_��ۃ{=C�9�������k0�KFT�ݸ���fJ��[��������ۃi;{�jw���S�G)H?VԊ����%�n�-����vC�q9.T��۶��9S=$J7�P�߻� ��KE�άO�}�i���nF\ȭe8da5z��m�� �q1�t�z5s��9��ě�{��>X��hadL��u�G��5R(���V�k�FYWr:l�O<J·lE���e�9Ƹ������u�9�T<r[�X����4T�ys�{F��!���2%:΢Eԛ�9ո8�
�u�3->�����iJ���9f�6�Q2������)7�N��F�=�<����f��V�]�(z�ng�Zi��{Ϝ��8jӀ�%J���ό:f���{��A�o(�V�=�����ymjn����M6�]�N�!J�\����Ac�A��lQ�W'nN���n�7V�F��p�����6�k�����/*��q�*�&y1�(Mk��S���@�ꗙS���S��+��+�vj�8��y� U�ܯ{�.l9���[|�/ؾ�=�;\��U��u�9
�+�)�''�Ùz.�ת��nm}�f�̨��~
7]rb�g*i���-uM��\:���M����[�{7B�PyEXqS4}���#x��+[�D�ʣ��p��~�����#�%TQ��}��Q�Է��v��S ��I]��o؝+�b��5��}r��i�5<-S0:��t����J�e5�Y+'�^� Ef�W�����k�q�:�Fʲ֨z�)L"z ��{�)<�ܹ�6���8짳~��K��R�t�*F�V��S8
)ޫ'2��=S�LC#}f_l���SJ�0�s� M�.�t�̙f[����f�R\��0��!�]BJ�`oiU����[��f�,ͣ�*���j�<�Y-�����O��ࢢ�t��][ұ�}�e�Oo�onb��pd�8�n8Y�<㈥��LwϤ�0b�jJ]�ب��.�mB9s�t��5>�
�jqyM�nQ�D)ﻧ���]���'�4��K�"m�=/�~�����g�W�7�`{��M��r̢���D��t�j:q]�]�	ނ��	]�Q<��|u�>9\��o�A�
ᛉ��	���v���N&�K��.���ے����N��?��ө����0S��r�/lg ���N���'�1�l����|"�9��R��O/
�_[��?Qȣ�����k���]��v|-m@�����Fv{}�Rų{��=�b跣#���)�q�N�k�*-����UDj�u[�/��c3�"�Z���lg��Kw3�͕��:���r3�����kw�*[O/6�#�-�� h�>��64��X^J�]�\�#��E�v�|�H�l�M�g-����f	�S�}��IV��o�JT
6��ٗ�����S�-��=�l���3ieAW�~׭жr��"I�͝o"��r~]���/m'�k��ٵѺ�c2�=�u��ɹ��K�=W�/���Fz��-��e6ż�f���=��ҹ�7�z�7
&���h̢�Gr��ʉ*`Q�|�6�6.7��`��T�x�yh����D�w�=�η�#=k�w�|���}RC�[��h�DV�~��?>�@�y�~���(ީ�q��5��H�:�*�Z�Ɖ��2�y��ߛ��h{�y���=o�%��oz��@l� >Q��L<|�_>v9~�ҳ��R�F�Խ��סgC�[pm*�P��s튙-��W9Qۭ����p�������r�-�\rƻ5�mC�r��SpI}��Pŭ��E�OD�q�%&kZ(o5��uF&١�I��:yu�Rי��x�J972^�(��s��jb�y����Z�\v�4�D7sYܑ̅|�N�7��:�QZ����18;Y�.�M r�o;E����vJŞ�����N5����Ol����P�e){P���<:�O�fĪNoe^N�L�f�0M����[�`����*��10�B��:]�ǻm�G:�"�2��L�m����y�:ew�J���������5��YJ����@�e�|�|�.1¸�R�_T᪨�-�Lt؞�ȻJ��:��	p���M5��l%�5��m�z����ԵZ�����7�y���h���䞚J-��ޒ{����tg��5ٿ�Ε4"v$J{��}pΆI~�sѳ��Xp(���ަ=}�x<1z��5�GzS�U���Tz�$v���-HP����uT*%��.�M����m`�:l.� ���u^�񙈁��5�]�4.��+}�o����}<*2����P���X��]ߓVg��9/��`�����K򓞺�]8���R�$��(i.�=0��<^��I�,�ܮ��}Q�a�i�x���~>���q���q���+���L�{~�C��Y���m�ϭ%S����S=�V�O����<����7��������>u�oJ��Bӳ�侣e��R/���U��Wup�u���.���� ALҝ���v�vS�Z�N����2���x5IR�X��{�Sy�!�l�J�"H��oq��;'�r�f��9���k[td �q�g5� �Φ�k�W:�<�%V묂��ytx�b)+&��;$�BO�x��2�����q����#��7#�E����q��i������o�B�8���^�rx�(��X$l���T��W��$\D���dB�יO�����Y�Y��{ޮ��t�������Ku��ǥx��f�Q�~Wkmq�"�cǫ�~Z�rZ�z6k�{Ӕ��~�8������SNd���sP}$L�\�����ƥ��Nr�W��t|�ƣ|�M���>�ߏ��~��y��~rA�K1�|�Sr�Q򁽽�~���+�Ez�<;B��q�F�n!y_�����O�A���XC�d�E��tv1�UH{7��<�"*��C�@�`��Hк�K��T��?T�_���o�h���z�G]G�eG�����ViN�.�2J����1Q�ތ�u�7��Lu���C~��o}A��E{�F�F���ұ��X}`�'�,\B�T�Œ�d��;��s�z}�J�8\v�߇�]��"|��_S�ͬi�أ�����edo��p��b�eH��d�|�pwjQ~���ܟ�;~�����W$,P�F���V�v��;ck΁� ̨m�̛C����;�������#��oEw9�]m�J����&7f���(Z��]u!�nL�uu�ε9p�Xwz�m5],�ܧ���`��>�3�h��I�ݣ�{�V�G���N7Q�NG;�=p�s�������ӷ���<t;GNt��[��_����͟}S8�㑳>����92�Y>���+��,U�pz�t/�;��j���E�j;��=5W���ˣ�;�&Xۊ������ٟ �:�<�O���޺��KUI?�ڠ�Z�xg�������b����z"Β�(^<|/��7��2��>�#O����z��z}�ݧv]���d��/��t�PK��*��r�q2pn��U1qS)���%JWBx�ע��@q(���%��##ׇ�;S��gG{�rQ��Y%Q�p������yw���8P�)O�_Or�s�-q$��K�x}��#�{>�P��UHۇTðl�J@SRX��9��'l��ޫ5�g}�V5��~Ws�ZD3~+J��F���޲6���3NdiA���w�t�B�
6���N��oᲑcv!��u�C�K��c���.���~����W����&^�O:m�ui��|t���;��AjhdRt�{`9���T���~a���>�d�w<�R���r�6��p :�r�Y���e�2�TXQ�/���u:2��0p��m�/Rt�W)��Z��)���Fwl���^�]���M�K1Wq�$�M�嶋��\��i�'����<�snfa�P�͎,�I�&��݄�G�*����TW�k�c�Y��}^�qY-t�BTǯ���+� �L��'6�v����:1�+��<� z�@�~��iK'��d>#�1��z��Y?z�5� ��~���#�ʊנ9����]�o�W�_���y47�� �)�*���alW�t�U>�Z#gvs�����S�Ӹ|�>��YP�?]����ߪ`痷,\qy3�,k�v� d�x��S�c�[�vn{�d�ў���������m��d:��ϛ�R�{�*��^�fp�������������
�<K���ꁳ��S�t]O�����`W۞y�~����V?U��
���ys҉����_��Zc��N�1��?�b�kL� y`�����t�^~����B$�{�moNo�H������l��VT�>%+3=0���R7���P��
�d�]��S�L�/K���xyez��Y��p��eHۋ�I�_I^5�P�(ϑ�Ey��d��ͭ������>�7w#���s����yNDW�x,���Q+>R�'�e�����Ŧ��|�����ct��(]�
�@I�Z2
�ɉb�g���,�[���Z�*w=���#�Z�Vu`�&�.ݱЮ��\#&� MXEMqG-�;f��;aI���8!�	�A��c� �%��f���nuqɑ2���z�nfR-<�"�V^��x!<$�Nn��*d��n���,����Xv�Y2r7fo ������G��RT����8�\�i8_k.C��P���U����t�ƭJ�q��w�PDh��#��: hsջ��J��右]�17��kv�N�h��8�,����/�zY?<t��j-�Q��3h�W�v�9�c*�t�$D�y��m�7�B�L�m9L�!�w>z�n��ƯmP�Qff�`a�o��y�/��yj�ȴ���r��n��+9ZP����w�1��"zV�Wr�FTT�:�V�FA�X����s���A�ë���Ɣ�Wٲ��G:��ʳ@���Z�qA�
u_��=V0�1���٫�/�η`ǃ4�E�R
�$I�m��(���-�eh�z��͗�b�r��"]�e��3@z�Km�Ѭ�$Ud�{"���m�u)�ܧ��rwC��}lr��z�7��2�/[޾m��������!��_eA��rm�+�W�7C���Uj��cuR��"+���Dŕ�J�ނ�άr챧�<�6�q�����<�t��̼GV�l�DT��C��>3W���K�vE��\���H�^��I�#��Z�����L�m'�n��k���X�.Wlfn�����{r�@7�U��r+��:8�aҗ,i���t�h!xo�[�T��匉���6-�ٸ5n�n�s�b����{7�x5�e��%���y�e�ڑ���n�_� ���Y9�Ri�:�3F]:	����wmj�X�3���1��Nt���wp�HYL��^`5)�Cc�&C!��{�{dw�41GXK���qV�}z[�&��]V@��}���#��fE��n���� � TK�9�C�IL�4s.���dћ[�J�p���.j�fa�\�&��eadŘ��+��=g�ͭOH]�P�2]�'Y�]g	�^3�Jw[.�c��M��;J=u;C[&��=aw]���9[��3���n؄��R��]K8�T�WM�B9]Wl9V�v+�4��*�rH>Z���!Y�bU�w��|k1,����Εa��F��_!QY���]i*�Q�3�e�' OA��t�n+��4�QH��ᷘ�\\���T�5�}o��#2���T0WmY�5\��1k�4.�i���Zˮ��9�v��/[]��ۊS-��(檊>u�U��G[��Y�oZA�B�NS�:�j�'Tm�������U�3�����ӆ�E¹�#4�v�/P��F���7R�n�pc�H\�ϳ-�Q^�����Hs�-Ƀ��L���*V����[���P�st�����UܟR����H�����*���M�"J.�2q�wI�Q�(��D5"��uɻ�dIF+����ڹnnsH Ƥ�wv ��d����nZ���A��r���vK��n�ّ���뻫�-"TF�E.�$ѷ6+�]݈���m;�QNur�K��wb(��%�9&ܮN�ws�\�H�d�-�n��\��4E�EȊ,�suݴ6+���N�9��k�˚�w'r�*9��[wuΘ�E]ݢ�p�.��\�p�r���s��utыst�ӝb���1X���\���8�1��Er��s������~���[%b�)e��T�Es:��YY�m����������Q�-�+�(:��;��2)�v��9��X�||.Sرl��Q{U����jxR�,�Subo�n�ǼG���=�Y��ڮl��lF���EY��g��V|����@���+Ō��[�^�!7�Z1=��{�a�������g�'�w܀�]ه�rxӂ�A�-��8�9���W�ւ�;c>��[���]o��oC�3Ӥ�{�M�:uP̖j�<LOҽ]Fx�}���w���8RӾ�Qo�7~�x�j��o�{�ԉyӡ�~��@�g�&�ϦU�27���_W��R��Z�|j}8�k}���jPr�3Ѵ|�ƣ��W�7ޤ�'���2��)d�������0'i�@��9�W�)�b�^�#�s�����\{�uTT=��h߽��do\ɮ��x�U_��z� ��%5�'���#a��i�V����#���{p���0��>��*��l�H��ײ޵iD�����B:K�0��6�;��i�qI���Ǯ;n�x/O��F�P^��5�{%.y��.�g�z3עżʜ7���pf�N�VW��s����`
�s��u�n/��(l��f����w��=��N�zC����M�+~�$�[�x�笮�dl	LE��irÝP��.P�;2�Ƞ����-��Y�h�E$SB��r�8l*X���47����WA��y�� Ӆٛ6s�(@��6�2�N�;$`��!���^��"<���̩q�N��f��T;���qS/ĭ�[�q˹�M{���� z!���q�ܜwQ��>M�!{mG$�EωCn"e�=P��^b;̙ޕ#�\��]�5mη�YP>�@w}^&ץ�������q��:3�$�I=U���}�,
����	�ɟ1�>u3�1���_���>�q�/N{���^w@�}�k�ʧ V߷�=*<��E� �2��R>*��B̩f麱7�~2>�G��Ͻ�Y�O�v:�B�vHڭ�w�ʔN�zc�.O�B,���$�vRS��u눯{8H���ע��x�..��K����SkmC�0������������:�p.K4���Pf	��q6zW��f�Q�ͿyǱH�.�y9jɓމ�O���#ӕ�{ޞJ�=�#�=T�ә.k�@�I-��HI_��m{��f��r��U��G�9�g�Ѩ�O��ȏL�x���Z����%�S��X��G*iMMi�`��w6yr�5S�#�/�®����}���#Q���Fߧȟ�����e�-{ �9���:������մ�l���P�m��LL|lX�	f헁�d���^�%ʷJt5��_[/-���.i��W27#Ď�u=�|;$��q�����.=$N�a��1��de�n�]�7��L��8�(v�����C��0s{�:�h���e8mo�3Cb�Ը�%O���R=~����7�����ߨ�m���ɕ4�����u&:����5��з�����s���7��GUl+����;����j}�O z���.#�� �O�T2a���պo�R��jW���\����wx�E�w�9N� ��72��r�����x�C�Յw2/#e���gv��O������v�k�맚N�}�O���w���N7Q�N}��>��вrN\}��ӷ2��F�UA�:��{F\�C%�B���K�����~8*9}��|�9dB��7��g@��E_���^�[=}	zuGx���~�2���Q�qR�yNDl�hu�yz����O�u}��t>eT�X�N�,��@�`S>�1�s,�,�R���ē�w��e�q�Xy���F8���4z�O��o=�����,��~�Ra���#�����~^�H��=��e�T�����3�fjY{k���pZ9�@[����qȜ�
(�rd�Fa�S>��l��b����mn��VG�9*���m]+4FW-��v�ܭږ�m�W�FG �f�:NU��ju�}cǫ�¹���7�۠�"2��R�RW"{��;L��V�%>�;��P��m\lq��ҸaΝ�d��K]�jZN��h�U���u�}a+���AI��IW$��U�l����n%���!zG��}��������`�)��t��{Ķ77�+l��`�z}��걨�S򸛉��#�\���#O_��Yq�fî��˅��ng��ܤ_1��.��j�/ōߙ�GZ�9K��c#ӝm����%��9��}� �~�4�7Fi!�#ЦN��S���D�I^SBⓥ��χ�o����^>��2�O1�P���[C�=���J�D�\��3�'��}/��n�Z鴥�8�;���U�ޅ8M���Ω��-g�b��������|�F�?]�5�OP2?EC�r���~��M�)jK��OL䰚�6��~}hg�����ަ�&���eH4�Ī�pvp/b��qt��x����]t�
;��}^�"�ߒ�����'�*!��Q��=uW��lqy3���D��X����]P�v�K��{�;�<=u���ԩ�<w��q�n���q���E/��*�߯x��w0{��ե�R�]��3�99�&|��r��*|Nb�����s/��gӨ�=�����&F�1�:��ޠ�ئ�vF�m�|�!ՍW7]�;(m�8V!��.���r\��/,�˼LC�\Q��~]�FL�Lz�����z�B�h��Rs���U*�i.���^��R�9D�p����Y���-����t���($�/<�ߙ^i�@��ݳ0�O�b����T��4��;~2��z/��{]f�-�s��>���G��Hw���B�eO%.��<4g��^�F�� �~�uw���~�t��K��Q|!�<S�/���9툿W��������p��*���0~([�J��\D�p�No;��J�,����*G���>�i��H�{�������^"r�+�U�	<�q��[�5n���j���Rѕ>�<�늙�����n�M�w�9�w�x�9��\{U��8����9�v�$�7���=���U��&����l����|s���	����{�h���z�������Ԙzܩ��}Ngo��F�� x7�FA�^s�	F�Zy�-'�t�H���װw��q7�{���>�Q��h���`1�,�1v�e�u��^�q+��&2'����3���?/_�������m���z�i��e\!�pzH/��f�}�;4<_=���]su>\z�����5گQ~s��x׀��y������`���=h
��3!9� 0��Y�x҄��+yH*����kyp�����ɤ��
��5~���B��H���U��sٕxԠ��p�R�>��4rof3V�*�h�Ղ�Ӑ1 se�#WW�ho]�Ve� ��,6vlE�x�W\7�
���'�������&��?R���x���������{����^&�ǽ����
��%���=�`ϒ�ͭ幨q��.E��N%i��V�����{p���1�>�W��K�;a�m�m?zw�w!Ҫ'���6|ωU2c�6t>��i�t�q=��Lz���|�^Y��X@���Ş��1
��y:k�6q��{�ɷ���TM�s�6����h��r�sW[ oy�b�����ݿs����{�u�e��W9��}�Ԇ�̋�,��z?r�N��Z�n�r������n��KBP���U)�8�WN&���2���9�	h�g�.�I���/3�������\��}]*���@w}^&�^���ߢ�q���q���B��$�6���2��T���1=5�N�gC��Ύ��jb��	sz�Vq�x��D{���^wQwԎ䞃������u��(����Q��$�2����Ԫ^9�̩f麱7�~;��c&���s�!w���Go8�'Ǎ{����0�\�iP,��vRS��Q>��{8HQ�n18�'����ʞ͠7|-���U�2�C��Y���z���wd�J�qZ�w'CC��`��&j�\m�u��$�JV3����1�����G8��S�+�Ҏnut��]��q��*�ܢ�خ����k�u��.��^҄���ǰ�]�=:�1�He.�����Omy��Tt��i	�n�C�rY�D*3 nx���J�{�tow����������.�=u�~X�9��=��!��{�Gze�d�)sP}$t磱��}����ݪ/�6o<����V�u��F�m?[g��x��߽z�x���Ih�Upf���:�3Z �AoHd�O*B��y���#Q���F�~�"|p�s�� :�<�P�ܻ��a{333c�U.d��g��Pfc�:ld�{ƅ�V:\o�����{�UTc�M��(e�c�n��ϕm��-�>�ހ�6*�̓_#�z�L>���TK[z3�u�7�wS|��1�<~�N;l97���3���G]{ʂ���z|���/��T��Ĩ�xN�q^��t�����~��Ӻ���v^
���c=�#��C�Vo��p��b�eH�,�߁��F��s箥��~�����t�>��sIӑ�+����c��q8�G59�O[�.�7 �6��^N��0$7Dz�k�~���_E��=)J���֗3�o�����QN|�~u���5+W��6�ez�=�f;m�E[gR�J�ϑ��Z�I;,d]jңkD�oR��i�r䙏��6�q�V�����S*�f��Z���Vهmh�ǳ{�V�,�z����YZ�Н�4!�)jZ�ջ,9nR��碢�;X	��Xݏ��o�8�v�Ơ�����ih�MIӷ<2	�*}GEԺS���K�p�O��箽���O�Kɻ���Og����\�欨VL�l����Xp���7�u�����4���f�U)��Χ=�۵'"����K����1U���]��� yz�'�:��=3>���=�=r����-p�|�?}�^���O���P�޶=����F�I@Ágʡ���lϏ-�Þ�Ԭr���H󺨔}O�q7>w�9��9����j�n��`�*�R �W����kޫ���ԏ��᮸��|�U�G"����z�!��Z_�þ�=�#n=4��8ߕ��ܜ�Ē��㧣�
>�2�'���:�o���X����n5�AdK��c���#�@��ulp��{s�+�R�ٯ�fxQ��:�d"H�cˠm?I�dTO*�qc둷�5l1�~���>�>�^����~(��8�g�5����e��&�)��/G����������=F���Q�=^��弋{�>����+��:�>����4
���AE�� �|n����=H[�w��\��߸�
�n�Q�jJ}��0�aV��S8K��u�买�ҙ�\��.g,_��6�pM���	����(�"��$�$�3��O��C��D�ƶ��d�aN1g-�䛪w`(���YQ>6�)��輸":��k|�귄�n��.��t�\v�����_�{ή��H��~�� =����.�-jm��jvޕ������=Ҵ�z���ۅ�����ޠ=F��u��t7�/&r��}������X�|���ȳa���co�T��9�/��m�{M{�7��[�=у&*��ܸ]�^^0�j�������Y���W)|�Cy�[�)��[���L
��<��T���Ι��5�{����!����~�걽���cj�t���PfA�,md֛�t�i�|Fx�ME�~��5��'��}�~��}�)��=�/VT��R�0���}2���w�z�!�_>=Ҷ�^�5z����q�Ss�~�,�Z'+�B�w,�Ƥ�b����_N{��\�\�sr���F{��J�Y�����q�{NF�G��uG���μ}9\�6J�Tx�x_{�ޘ��s��J��I�P�c�2�>�K2�З�߸�zG���%�Q�W��ﯢ槮L{k�ܐ��A�+��<j�`B+�{���c]o�}�Rq>������&��%E�6'��+u���[��	.#7V�k�&X{��Gq���й���J56�Lb�l��'X��\��ehVRɕ',�RJKw4el�}�Q�Q[x�_q��J��h9[\�fΙ&���:]krȱk5	k����æ����
�2j��=y;!�"�i�Q9�UxñrY�P@H<�#�J�`�K_�����	���W��ծ`ti�!�N+C�=�\N{�z�Q4̖P�<LLD�WQ������{^*��״�$��tg�����#�ǟ����D��N�M�{ޭ��뉯�ϦU�26zHV/.��9�x�k�T3�o�}^��^D%p�n;��u�j�E�ҁ�� 7�h�ɔY<*|����&���n��e��|���O�"�%��Sf��}��\{#�wtn��4n=�P��Vח�8-ͱ~�M�W�ޖ���멓�Ǐ�����S��R��}^�����<��v�d>�W���`�5+
~����q�3�k�e#�3���U@Ɇ�ᵡ�����:�;��_mޏ|ܥ����J�<�ƑS���󠜽�U���u���l�N���9���Q~�G�X�}�����M��ј�[��~�lg��}�;�/�43O�g��̩p���pf�0̨?9�
����6rtd��r���[g�S8�Y����vE��Srq�F��M��нS�z��ġ����"�'�^�����?^f>N���;+vS�".�+t]Z��eWP�5�J%G.�F-O���]��
c�i�b�f�s��ihfh��<y)�
��B�i�_'M�C1�.���.m�ى�G���W4���
���PL��ճ`�sw��[��=���o�D;�A�SRPm��b��*��٥t�1F��û�|p�����-���˜�
*��֠�Ux	�K+z\�W�K���%�M,�� m�{D򯝋�ܻ�]���Kr�60�����m��Ăġ�Q�/�����]1���	���[�f;�o�ywҶ���(��
�S�U�4��ݹ�AiJ�-�O�{��R3:�,�k;HVN�ێ�P�{n�l�������ÛH\O��=�4&a{�}���t��ыr����y6�h��]�N�{����طt���D8v�۬=�J�=w+��蹗�V���,h�3��d�W�P��T���#LB�[��N��%�b�PD�[�&� �X/��8!�r��D�2�s���x�،�x;�a�a�(�곔L���������W�����N�)���1S��8�qΏ�e��x%G/���ӳ��6]"B���!��Tm�'*�p>4eh��sk��������;Io�,�k��
�ժY�n���֪��\��>��va��Φ��u��h!Z�`�{o\]�-�]GhġEgfr�M\�Uc�F�Q�{��8Y��B]�d��۬���j�F�S����}b���o�G[Z��xr8�4��z_�]q8oh`�n2FF�X��[�c�"����`��ژ�ں8:�7�+��*Z�pgl��қ��e��8S��] I���Yw}8X�Y��ؼG7L��pܫ:n%E�ft�A������%��)�`j��%��ͳ��Ns>h曩y�.�7#GmK�&MɈ�n��=&��)bLv�wuQ�zU��g�Y����������I����I�ͣ�-j&�N�p3��|��q��db+w�j��(���P���ǋq�l#{�Xh��p7��+��Q�P�㧮�,Z��v�q�@��}�)����^�w�.��;7e^�Ɩ5>ŵ�q؅����G�#I��&�8��Nӓj�#�I�j��M�[ZiЁ��[s��fl���G�+ӗʡ�tv�>��T�n����Pp��м�F��Pb��ֶP��-��}��tQ�At�����-�ҡG�oV,��w@l���펎��[H��Iv[W�Wb�on�Ver���XE�,]�G�:�{@0,T$���ZŮ)N�s}�w	���S�aQ���g����e⤭��;r����̸렶8��bR�i�E�ژ	�$�1�r���eͤ�\W����\��뺆F3��^�`|oT��U˧hh:D�w������ؽ�Mu��E[WpD���5�P��φ�BS��Z�U��ק���Su�O"Q$�q��1Q����p�����c��W1'+��N9���qu��˺㘹b.����b��s��,�K�0�nG*�F��u�s\���N��.cW$ӻ��ܱ���Q\ۻ�-�X�(�F�.U�nmr��wW��s&��%Fƹw]���9����;��;��mnnT]έ�W��F�\9���79�h �55ʹr�n\�L��[�����r-r����v@�Ȃ�sX)+3H��q*�W
�n�Y*e�\����N�\��ӛ�\�J���y��^����*<��np��lʌ`�8"`d  ���bW�6�]��	�F�Y撏,�H��
��ܖ�^�;;Ȯ@e�����>�ۮ��u����@z=>'������q��}^W��Cs�[KX��h�����[�'䎏��I�Jt���ϔ����K����z|
���=���׫�I��^�P>�M\b�5U��nN�{��|O���@��3�i�-c~+�2���n�O?W��P��@��&�%7�2FE<�~��_���ݟ�w���|��*��AH�Ge%9�Q>�3��G9�s���O���?^�������*:z�����t��.K5���Qa����lo1�}�Q(zZ��U�lש��x�k7���n"}�dC��#���Hq9�I�%��� r���d��ק<}�^y�..:��8�A��H��1��h�m����������߽z�x�t��	�Q�H��m����'Q����zH���
��SG�hR�n7��m�+�~�"|p�s��(��	���(���F}@z=5�B��A��;�Ղ��=�B�.7��>7�R={��vw�k���wt*3<h�v�@�F�GO��5�z�L>�>�-m���^�}���6�WLy�?i�㺍(k��.�Pv��-ibDl�թ��!�� H���K2��H�7��A��|���{q�ݖ��A�9m�u�`ǲ�='bZ�p��zd4�"�L,!��%j�7jfi�Ùr�'�\3�����S��"�u���<P�{B嶔��86��{����> �G�k��g�	���kP݌U���.�p}ʛ���+�(��,|F�zt�y��8_ݷ�ᐽU�s�ޡ�K>�^��~ڱ,ʑ�Y9��&�u)+���6�[�Q�s���Ez�����t�����m��ϝU{���9��Sy��f��U��1v?^kf��[v9�}䮈-[�-d�>���e����Ǳ����3���ޜPf�����gSZ��>�o&X�jN����<�S�:/�C�sfXC�нO��������u���=SyáH�a?Gl�e{��j�J˓��=C8�bI�;n�/8��;�F4��<s˳��v;9>�G��Ԇ�{���^�<��q�]�(ݖI�3�,eL�r~��a��z�J��Y�������?~��>G=��_��[�9<��������1���S��x��Q{Y~���יZ��'��+�뉿����!zG��F��|n=��mêa��V���*��N������< ˟}%!up1�2�C걨�?+���z�8\���#O^{�F�HO�;�+F��p@��;�-��y^y�;s`ch����t��YY�(v\e�Y�^���rE��L���\k�����zi,�6WpJ�R���Ƙ�֡�j���T!W�ڰi�ʒ�V}WV|�LeG�X C�6g\�+�l�B�gvv��m^�nf���ڒe(�l�$?��C>��D����X�#���8�~��dG�:�/f�Lq~�N��~ �N��\�uLȨ�2YRa��u2W�и��x��>����j�ގb����Ws��ز�!��VYϠ�q��&.�uP��=bf����}^�u��M�ܳ�o{2;9��Wm�jWF{Ey��B�+�	��>�,~�@����Y= ��z�lyǫ�B3���y����
@g�W����w\{���_�G�����}�_���j�x�X_L���WZ��7�a��F{s��c��u�5�R�g�?@��<����N�?]���@z�����{r����ڰxK��$�Wg��p�T���,���cgG�++�n"�>'�oK��Q�&}�=�)x����r�u��^��ᙰ��g\�~��C9��<rsbg��i���(躕_���U07<�<<�k��5�37M��$��{A�;ǽ�U���^���:mN홇��	�,\VMi��t��n<�ԠN]{����t} y���#>��_��]{ǲ�!�}�ѫ*xݟ������m{��/��}��?��dn���I���M<G���
p��w�*e���WFjK֫L�%X�+w>��ᰥ!Z�'me!R�'�KXf�X`8[V@��4�J��\�5h��;�������ti�}���C�Ể�ۮo*f��˗�^w��c{eD�z��R��~�����#�P�anȿ�Jn{o���^�<���Fu�$�#!R��l�##d���*+�K>���ps_ށfg8�n�O���Y��Ǽ�+μ8��T��6}GL��phI��o�
P$��e!*�]L�>��7�X����r;�<_�Ig��
P�.��S*x�p��g8�����&��6:[,>�?����,�����y��V�04��D�w~��J���}�4������Ǫ��b䲠 �� ���I���;�΅ޅƴA�_�7o�������2|��D���<o��_?R�n3޸:n#��`�r�����uV�fN?����]-M�k�/G�F��Z�/������D��C&��V�{=q4�}2����@��A��/�Tb�,�U[�=��WQ���#׉\{����u�ڿQ�~� }�> g�u�W�ꜙL���ٗ�"�.�E����%#㳂�uh���x���R��?uǳ�y�Ѹ{+�ѿ{�{վ�%lV�{�=�qT}��|T�h�b��>7Ŀ\-��k���O��y�~�F&�`�����W���J�P+��t���3��-ud��]+��5�Jc�OU�6���O�Ew5gm��z���`�s1j�*��(�#�h����.b܍\3��%�]�:���j��i���f�U��+*tV��'0��s¦)q�z3�����J�)��u�5����Q�a�7�q�*�d�V6�;���t_ԝq=�wS��p����{st���@��G���##}����V
�u�w��b}��f?�����
�Q~Ж��Ĥ����^Ӛ�����WV���l[�wᎫ��3��/��V7�yu!{�R1Nf���Eި]3�����ۜ�F{��V����Y��`
�M��Srr�j��M����rOy�0i�H��y�
ꆉA���FUG�L����y�������z������ǼVW����N^���IC�`��G���qcK��3��>S��K�����>�y�/Os���q��߳ۯ6Rl��DW����a�P��O�s#��t���s�z��m��2�К�tnr��y������z0��F�/G��ȏuz��q��9���F��%��� aK����S0��ִ��U㉯W��r��н��y�Q���'M���;�\�k�D*3X˞��w�S���y���M^y������5��*�S�,C!�W��zxi7�I�P�9���Cz>�E�aW�*e��2�M�D�w(���E�[��\�5��mfv̻���1�=]뻘Nϰ��V��o�;و��&&q�k����-��Ek^�%#�c',a=���fd��;]e!\�:�T�omI��P�f�t�&:]�NGU�E� N�b���Ē�uG�g�}$L��c���a�b8��c�?[g=3�}�=�����@�%��I��W���)���$/� ����t��ׅ����g��7�F�my_�����n{���1X.j�<�hg���s`{�4���Pfaz�V�x���K��/J���{ ���b�1�AȢ��{��f������b�}fI�Y=a���a��koF}����W�6x��F��|����^~���#��t/羠�n=������.;�Rt��a���0��
�d�,J��W4�~��������a+��q�m���U�_zG�s�9cC���N�H��l��%.o�A�N,�O��>�����RFIzN����~��Ks�W;�=o�8^Ps�=�߳��M��އ<�����
�ⲫM��J72�Wы���L���̮]64kت�sG�l��F߾�u�:*�to��t�̱�O�T����t<�6e��4��6��5Q�Gw}yw��<{D��^��O�Fo|�Q����qe��pe��C�t���?!���خ���k4�'	��BVM�6��0�r��=.��]tU���h����2���$8��������$N�ww��^=F����o�]pܰ��(�� ��<~�4Y�����rL:�ia�5�v��]�ŗ3���,��+=OWo!����h��O_b)e�6���U��>A��W���S�G�^�Y^�<��1�.ʔn�$���FU1�Qq�^�����v9e�yq�z�
�^��=�����sѾ�\{�Ǹ�ӓ�_��H�J���s�~�s�{o���GeF@�j��L�(yw�>�TI�a�/H��� ��G�T��Tï-�����w����S��&� ����x�t�[顈���q7>��C7ⴧ�z�\wEh~�Aw���|Ez=5�k�AE@���1-�c�����3��R�(��l�>�g`������[�t"0#�O�|��ﾆ+>��O�j���W�и��x�3��mi�ӕ*�w�f�2uP(�Ez��xa���>�d��ƪU�������|F�&��;#�_�2㼮!ҿ�[��n���6ܠ���Ǿ���M׉����ƁO�r|�����^��	?Y���;��jf�����[�>���_uG������utn��u�W���Վ�̃ʐ��=��\z5��x��ax����)V鸊��#�K�q�{p�!?]�����*bsMȜ�EUԷ��_��q_��;�+���-r�>��}+q�b
ʺ;(����dz{��hi�]�*�`���C����3[�)���%��L�����M�I��$�5f�f]���8��jWlPF����K�5��BA���G_Rܕ�]%꣝��79`�CeTM~���ɜ�s�QX[gC������>'�}�/��m�yɟi�e�����{��[��,��i�y��W�׼n<q��h�����~�:��*����y�N[���k�O8��S���̬�����z�ʹ�*d����|�Y5��Nןc6�����uu�R��c�����}�x�DS�;�����YS����R�3
�.p-S��p魞k}Cv�}.e�}֨>"}��"����^Y^�<D�p��eHڞ����MG���vy����i	��t�Ⱦ!��6��3�WtCoa�}e3o�x���\{�r+μ:�<�g�Ul��Ô��g�7��=_)@��2����C�����-]n)��<�{N���nɴ�G�F�ו�W�#���'��{�p�>3���liAʌ�& )^3c�����U�R������9{�<ծ/�'�4y{}m�uG����fQ,� $��H�=+�w��F�6�^K�)��������=��c���g�pt�}��D�K8���|'����{W*�������j�@I�5.�F��VSe�9N𥶎�)�>o�΋a��sw$����!�œ] -q�w�7԰>g����/8Vd�Q���!��e����~�=k}�e�j�r��Z��s�#f���䨮�q��u����Y�X���ؓ�-��]�j���{��,.yQ�^���f�]�kY#�~t����D�>���{ՠ_����ʛzQ������z�zC���T��ԧ�j������5m���J���}�h~�z{&'�W���U.�&Qd���D#`��7+�l��K���Q�Ux��ex�2��y,˪��7�t�!�xe�]dy֑qW����,~X=mv�T�������s��y�c*I�"Ś���r�r��}�7�}��ֹ�d��rO���D�%T�j�և'�poԝq=R
��S��_���g�+��zϽ������N;�`���z,\<ʜ:�ߌ��@�����>�'�4����v:o�Ϣ�+A��;��7����3�{Լ^B�X�9]H^�T���,���K�w�Vj��֜i��EiLg�*��T��+#Mx_bnȸU)�9�WN&������)��"���}W
.�o��{�]�N��	[��#���Vʀ��pFL���)��u�щV;1Kō��v��r�2M8�����mWȓ%����_�U����_���>�rܸ�c ����Od̾�.�.�|SJ�Z�-�P�gL)G��g-��;-h�^��G��ɰ�u��IG&eG,�c�6�Fe�2I���巗�}�lF�h.��ޣ8L��� ��:*��Y���/Gd����l�eec��x�D�������+璨����6���hU�{L�i3�s(�A�,\EJ���Y+G�T�mշu.]uˁ%�<�����z���Qg��y�{��|.J4��*��AH�{>|o�*���{�vy]��Vϣ޺�r�|$tO��FB�י[�z�������Өw䲀��l�e��,��y�ƪ}���\M���>�f�Q���\Mϼ���y������z��L�?Zp�A��&�n��=Nϑ s�=$L�����C��oZ5p����G�s��v��D�ؒ��)o������fP������f�L�Ѹ5?���I/ԅ\E*h���)~;�f1{��v�3<ƹ=.wЭ��R{p�}ӜO�� �sL�H��Ff�u`��=�Bq��|�>=����{{�V\���>������y������@u>�$�Ћ'�L>�>�-m�֯�td>��ml/p����~~�����c>o�t-�:�x����h�}���[&ylM+���p��O�1���v���W�+��q�{~�^Gz��,�^�߶�Z�F�}U�N��u����;��b�M�Е��G�e�.Iԫ)��%�7
�ǫ�ޘv�Lu�̕*>�3?H5z׸����Rq��efRC%���cZ��w�ϵ76��F�_�
u�����&�?�iEk`���tZ�#�Hk!]<=*���׍�(Γ���^��"�BmH6��n�q`S�m���������i�/i������`ߢR�R�W��(U�+ rb����m�-v���Oۼ+����E�N��< '��ySJa;gnf��������ɴR�l�B��.�a�˵�s��(ӊZr4�	�q��77%K�����Z��3�,7`�Hب��[�:dL���&ˠ#�>�����Ĝ�h].��u�F�-�J�[1�k���Z%!��J<�L�ԍe�����!���ih������a�˜H��_d:��sS�\�w�i�s��9U�0�ï�1����j����q�p��/���(��U����+����K�ޖ%hAʶ���z��X��i ����l2�-�έ���[����ͬ��R��f��j6�a��&Μ3�µȢ\�\Ba��F��l�	�aokĭ��_γ��k��s��i##q�ؔ܀Zm�p�Mub�N���f�'�FU��j�\[��6�:�/
=.�Y!.�[3M�ɲ��0�I�)av��A�k,]Y`�].I��6�"K�#����786�!v���;�Rn�]K>IQ�)�� ��ǭ��lGAڝ��y۳/J����@�wg~ƕ����Q�uu�S�e��s_Qb۱o��3����z�#G�)am;䵵�ӷ.��ѧ��2���Q�w�������'j���9���������P���Ԁ�Nب���o;hD��L��`HtsI�.�N�R�W]0�Ψi���&��Jm&w:���zV����4q����5�6���Ҭ�~[&R���e5HLN���1�}J>Z_>�ź�X��79V���.�s;9A���d�uN����(�x�CNAus6w>���hR��"֜��ӥ�l��ԣ/��p�,d��4���jk9�u��Zd(˵IGh�׮��mQ�)=�.�d6���G���V�;����|bd1�ޜ�A��9O��Cgjv�&7��v�����G�XM]���2�t���H�e�it#��8+�����s1U�7�ZB�}]D>& ���nwYI��}s"�Y\�TL��H=F�ʖs�����c�;��ޣ�J��*��k'�\Yb��r���hk�T9�a�#x�B(H���O7z�����(���
O.E��\n�R �i���=���%�t��㍪٨�JU��]�!F���4�W6Dt�B�� �EPB�q�tq�0��HSR󓥚�n�я�l��,윒r�)����O���[���i}3r�;���]�ٮ�닖+��v�\���WMrMr���ưnm��sDj�]4��wTgw4Cw[�r�7wW8X�Ĺ\����v��5��p�Qb�F(�r����F���R\\K��r�sh�
��ֹWi9�������D�Q��V�k��Q\�E\��i���7N�\�h�!�(�W.#�(�
#N�]ݤú�M�q�Nt�D��J�c�]�;�,��s\�J�h��"�]u�,�R��F5�*�MJw\��$hĦ���ܺ�2RQI��۽���=��׿���YWX=�q%�L) �2[��3.=��ܰ����n��+�X��9�W�ƌK��˄�Eth)�0,��Ip,[?���Q�YM��^��!t���wᎪ���u�󩃮3ђ; �o����'a���m*EK6�r˖�&>V��,/Ж�SZ\�[�C}�[��� !m/l=�����>�7��q�z���9o��>�@m��!����ed�8^>�g�՝){���;Y>�}��X9^�x�SW����ʝ7��O��c(�ē�jC&�ޙ�0׭��U+h��R
h/}���E�S�G�^�Y�z���9�\�;e�z���o-㺵<)�ھ-M�Vy�}S=�t�����������O���P��c�T��W�(��uMOMt�˶��8*j=ĜA�T+��^/b]���W��q>w�8�#�{7��q�U#Ldvf���s��	�B|D� s擄!��1Ų�Ϫƣ/ʢTO�i��<W��K��Ob�����qd_�������d��(!_O���끿�K�cu��n5�AS����t��]um�^#�ӊ׎�Oi7����ު�Nd�J���D�%yM��x��i���S�����E~T}��E�ԻJvG1.�oGma��μ� v��Cx#�\v��3'�k��mE4�E����cY{ �,�W,���r�;L/��'2Mj�e$wU[�� ��K����a*n
R���b3L\	�!���9�N�����{�A���^���F�ʼg�V|s���K���MB2����^��c�+)3����v���R|���)t�%L{��G����M׉�}�>}�ƁO�r)d�����D��:�ξDM���:�=;պr�W�^o\>7�?m�g����=� ����}&������z됪\&\��S���pw���w��7����ӹYQ���9��P�3k�i]�!f�{��/������yt=�&s��9,+:�W��R�����~7�m��:v���#�ﳚ�MO�Ly��&^������7���G�gI���goΩ�[G��c| *�T�����a�~��z��<׫�Y�c{;ר�����Y;�fT	�,g��kn���1(5�_r���|��EJ�9f���'o�F}߯����:���>�����eO��R�p�"}wٻ��#.����g�=3�z�@7�ƨB�-��Ss����:���r�9�����UlU��k
'��>��Q%D�F���H>Gk��,�uP�W����/s}q�)�����ۍ��գ߲�Ck �,�b�Z�(D�V��1Gis1dgT��}X$�G*v�*o�v��r酢�����60g�#a:���#�d��G4*7�9g
ܫys����*�����t����Z�"�˧&D��)v�:�:�boB�G�`㷽J7��R7�_�')�d�	=�2����C���[��WE��n�O7^�+����y}㕏��ZQdg�����(��{U��3��
9
@�.��1Ų�������
*�XÕ�N� $�'��~2=���{�a�������fQ,�( $��Iǳ��y�F��r�:°W����gC�~�ȟy���:���\M�pt�z�Q5�2Y@@os9*�meD�3#P�>�c�;��7�l�}��F�ֲG������>������h�\M
�t�F��i����驕 �Di#Һ�E��Е���3Q����~� }�x׀�������֔�9����(Ϩ2��'@%"8��K��W��z�"��~�g������W�i@ި7[������t�>�{��U�G**�a�6����i�t�����({�r6��Ow��ǖ��=�yݢ��g�A>��3��w�rKa�
���>L5ckC��8�����]߼�-�u~�s����;n�x/O���s��h���Xws6t2s8�/;�j�QKi;>�+�X�揦<}=��; �o z]7^�>O5B�x���9^'|�@S�N�\��X7��� ��ၐ���NV�S�2R�*0_bo���zʓj*���H,}�Κp������YA�����J�U��hԭqg;1�p�s��W���K�r!u�Dny߆C�����{Լ^|�V7���
#s*Fm��TO�}����9@�q�%���5L{b��M�ϼJ�,i�!©M��wQ��!7H)ܷ����5N�w$�)����{S�2'�=�S�]��%'�p�T+�U#q].���@w��W��������KQ��Q�}U7�
="ϡ�Ey\oc�B�:rN����x�=�g����)���З7�VU%"�GeK�Un�>�g'��z��ӑ�O�VEy�yg�s�B=�Q��$�p�bJ��p+j+�����Ww�]U�O��V&���p��G���IgW��=�ߌ>�rQCĕ�e��pʪ
2�fC�>��VҊ��� "�gнu�{8H>~����V�ޡ���HN��N��ʷ�;Ӯ~N�d��]�+����2�^��~'�݆j5���\Mϼ�s��{}�C��zH��oѾoEeU�>�2�W��zd�� �.H�n�-n��j:ј�O���L�x���_X�yeds��.��� �9�f�̒ѳRٳ�D�/ԅ\R���
_����{�@���̯Aw�.�+�����vC�({N��HI^!T��^�S2V��\o[�B&\�[��
�{�zPou�|M�a�ɽ�t�_���(���j���r�&�%����/gw�VU�vUk��Fj����-�/�I�����}��MЖ�*�ӎJ�e��\���' U��h����8�*�>nR�~���I���/�.{ƅ�c���$ۅ}G�W�o�ctg����HW�+�1i�Y��}|�:���:}fIA��f��}�:.mC�����_�쥂����W�K��u1���C߮�_�}A��{��\y��ʐj#�Ĩ�(�o�� D�#}��J������ǥN�ߢ�����~.;oo�zg�^�C5�������D�W,�6���sY�\��O�PW�r��$���}i0�XY[��{iׂuU�'>��9��E�����w#ڸ_c��;�5���y9'.:|��/����x�+��Q�.F/;�_
ؠ��9wվY�Id���n|��>�O"�=�q�z���ɝ�'N�L��O�>��K��)n�t�4��vwW�yp�t} 46�D{��|�}�)����֣�3�l�|�� �c�rnj�=y=[u^*�g.�j9m�y�t�"�9��9`�c�S��W�VEz���Ʈʔh2OnNm*@˞���/��K��>�<�Y���&�����,g޽�>g����L{I���.���v$,"��_�'�ͬA��z�Ik=�գJ��"�_�-�n�N�U�4��v�����l�!�*�Xa��y�����1A9��Hk'D�w��7�+7����:�3Mt�2H;Y�������͹G�[N�~c�[8"6`�m��Ha�xK��V~~�!%Q�P$�Q뮚l�uQ>*���i��sپ���跑2�7*�n��^r�zOzE�=U�X6O�H��,	ׁ����o��#/�Q%��'a�jM&/=�]t{�����鳜}�4�{�Fwޚfîʀ[>�'�n�/ō�fu3h������M��������O�~�j�VOqg�,'��X���O|��l&n�u1%yM	�����%���ڛ3��+��ǷʤgB�2����N2^G�F@�n�j�'��3ۑ�Gm������U{�Ǿ���7�d�t�BU����+������|���*���]���L.�>��;c�K�BG�w**WV�ȭ�x��o\>7��~󚢾{�׽^O�|�s=Us�x�{��^��ە ��V�q���]z�M�l�>GT�0Z(�刺k��n:�g\Ƴ��O���G�LN{�ܱq��3���DaaF�����O��_�����yo�{������M{�d{ފ^/c�w_�^�q��Nlχ�ӡ�ENQ�*�����{�e�jb����@�ث4��WV��:��C ����K��AB�c��e�|�4x=8�����u�'yX�Ϯ�,����qԼ�&��iuHݩԎ���Ӣps�(2	���a���^2��[EVf�R�R�
�Au�N��� �����F6 I� q�: 9������uO��gӬ�����Y�=yS�Nf���m3��I��U���ѓ��c�^��qS�Yi�Q������}���K�7OG�ԅ�ʞ=X��ɭ�M��mG�+�f7*a�E*�z��ڎ5B�싌R����xydW�V�dS=�vWg�.2Q�`��eH��΁�yq�rs�-�3�M�L�VW��o�x���h�zӑ� �r��ő~��}�8��P(���z����*�qS-φZ�,�sB_�wYΪ֛�mv�hÓ��̆V�G�K=~�p� �2��liAʌ�$)^3c�������W5�搹���ٗ���%��Оz��w�i����v�T�;%� �����ߣr��~kK�5��$z�ܧw�gB�~�>�<oi��.&�3޸:o�W�&��,�%�.�*3�|�9�8'Tx@{��bb|���WO��11�\��3��D�<p2{��hh{}7�>���κ���J79�ڗ�},�}�X�9�/��R��Į��y�������z�>�����/d�X�Jk��n�H�Aۥ�x�of�1�od�xd��ovR#��;�^��������n�j5C��`di�T5��;4�G�xR�S�+����jU�+*�Xs�"�	��g>P�
hjq�`��wg.�w����4��1\"G�>�^��)�qom��g;����1�K�'ƪs�[ŴTo�I+x�F��*���fS��߱�u[�;���_Ql�G�{ޠ;�P��>��Q���A�C�zp;��i�qZ��-��z�{&$��uW�s�GVe�*7�~�F2!���F��.��^پ>�8xx�a򁵡�Ǿ6��9��fkW4�)�#�^N����=�U�þ^�,�~�ޔ��`���z,[̩�zY;��Tɉ�5~GWz���Eo�J�����7��*�������d:�_xϽ=��X�9�ԅ�������3���M�>�����pf=��UⲫM���+#M0bn�RSrT;��ӱcy�A�=���{���vo�������=qs��6�^zadE~�F���9�L��>�s��]m媼���>�ŴNya��_�*|�3{�hW�Ӓt]�$�L��<�L�L\G[�.n�� y�e�;�[��u�4O�~�U�o=C���z}Ⲽ�<���G��7�� �`@�,��ݕ��M���s��]��>�~�q���ý�1������d�w�P��*��<߶�EFٚ�vS��VN��3���5<�H\��E���.��{�b�"��"��U�b���u�X�˗���ٲ]�d�΃����l�+GJŒ��u���I^!ԅr�ㆎ������U�5ceǕ���	C`}�T
���P�a%J:�� �@-(���9	�D����.|�z1{k̭��=�'�0�/D�/�"�9�ZP��|t�!��1���9��^/u��G_�D����!�9��=��RLҩ�1�YN�Y����ܩ�|E9����" nj���끿�KG۱�j7��j6���o��##�b~�B��P�a���}��U�>����#�_� �%�]���:e�F���M�K�7�v�`h{�K'�[�D�+�?+��z|��7�}l�!zt������Y�>�;�vrVm���g�ƣ��5��~����~������߬ѿ���;��lq�'!OPɇ�c{E�Z0�߯,�w��5>Rc�J�ތ��K��K����wB��:�x��w����A�y#�fQ�#���tj���%�\�����T�������~.;oo����C�P񥑾���B����6.��<���*�i��̩ω����0���TEL�'J��_m��ϝU{��9�\��R��}�>�;�=~��
ID�b�,�:���ꊈ�a-�4��|����(�͵_����,Pע�tn�|:�f�N!^�y��B1���p�)R��P�l��
&:@�ܗqTH���N�t����kn��%&	��j��I�װ<�x�v���rX���vM�����Nm՞wψ�oTK2�M�t�/�X���Ep+=!y��>��3�3'��SL/��yC��/^�zo&t/�	b��	EO��N�1�'�NeD�{swg�R���S�2�w���n�����^��j�y���Z����c6�i��&�LNc�[�t{o�ŏT�x�u�/8��<���"�ǩ�Ͻ����J�s�.��mw��Tw+�כ������{�:b>�3�BI�;]u\RYbx�ף#}�w7��z���xmCv��u��1��)�`��ơI��O�C�2��n�|n��|��W����_����
s'�Ѻ�Y��dg�UL;�%" ����u�lt�[顈��TL^���$S���{��{��vO�Nx�-��=�-_}#���_$��>��2n�/ō�g��ȯ[��$��]/ux,��l�zs��<w	��\�ό��s%��T�w�����e��U��WX�=�-Et��4%�\w�>��+���������ώA��%�x�d
�v�&��:��Z�nGcnn��EX�,p%ي���7�d��y	T:�j�1CuR9)�����������_������o��[ko���խ���mZ��m��m��mZ�Ŷڵ����mZ��m��m���mZ����V���[m�[o���j����m�km��mZ�u�ڵ����j����m�km�m�km�M�ڵ����mZ���mZ���mZ���խ���(+$�k$xi5`^W{0
 ��d��H��z(Q@
 
� 
  PP�%T*"�)()*�I(@QJJ(� �IE(P R�P�D%I$�)P�4�%IT��DR��TW��TJIT�J�H*�H�ITR
����E�
�Z�U** �*��� �H$��UP���**��D�H� ��$*�@�BP�$�Q�TEE)
�(QH�UR�4��H��  ,\�]ڶ�;rݶ�;ێ��m�2���g[��Kn�sY��m����h���p(趵FI�U��U�YQ�gC#�Ut�H-$H����O   m]J��z�؜����lݫs��3��:�Q�E{ P 4\�Oz(��(��pwhѢ��@n��tQEQF�t (�Eht�(��sE$Q J(RP�E0  �ƀ�G*/yN������l�L��@sjT��;�4֮ٱҀ:��[:H:�]��wY�;`km��$P��D�I%�  �QUD�`ʠ�6�1�]��Q`�.����wR��wm�ڗm�'LM��k]:�nʲ��K��k�b��ݮ��9�JU@�R �M��   ��[l�mU�v���n�]P�qp�"�mk�㖻����eYԪ�wn�w֛���K�ۉE;��5�:�B��n�i�C�S�N�ƻWwwYWr�Q))!E��x  �x�[Z�wr�nan��*�]��cUZV�j��6�Ctv�wN�ih�qW+�Eέ�\��v���;�몱��];����:��:v���ڭv�ծ���Ҁ���!!/   c��f�5۶�w���Н�)�w%m�յke-]ve1�[[mj��;��Ym�v�us)\�p���tm[L��T���'J��t�Λ*�v��Gf��   6�oY�*6��+[jں]u�:�-ۍڮmv3���Ԯ���Uv6��Y�Ws�]n��l�4�4�vi�B�]��w]ٻn#m��N:�%�MZ�V�.�"$JD������R�  t�ۜ�����6���C�ݻ�5t���wk����Wl�ۣ���K:���h��6�흵n#e�j5V��Y��v���t��j�����i���u���E��%�FP�W� �G��^�黡�8UvkZ�	[MV�Κ�][��n�GkM�Wm��C�DF��[���[����gR��;gv�]ݍ5�XS��G*�n���w����fU)H  )�)J*	�414�i���`"��	R�  �~I�UT�b  ))�*�� d�O�~?:����1��������o�ݜ��pX��}w�����������:��* ����
�+�E?�W��* ��AQeE7��9�������ֿ~֎��6��ιVvV1�5��Y��R��)��vЫ��!��  ��ڽ��S �����ق�e����u4\�A�nضE�W�UmZ���/6���0��>w��4^f�`�C4n���B̼��W�u�Doγ�^6s�E�9�wMZ>��ثo,�C4�\�)5�dn̹z���Eauvs^ޕ>.�k!�74����f7W�,�=��4�@�ܫ�nby/Y����i9���.�(��e��t��;Cs&�6ٗ[r�����ʺ4�"�z��C��i�4l��B-��Z�lT�jV�^l�i��Cv�Jћ+l�k3i�+�P���u�1��}˪�kv���i�4V�'���c��ƙt2
Ԃt����D�c � ;��԰i_#w/l�Q鼹M�ۃ�E�����l*Ӛkm]3V�D̂9���U�M�V�m;���)�ZP5�]�[w���z��+8��t/p�IifX	��]�2cՌ��]fh:e�i9QH�^YG�:Y b��"�:�gQ��T1���Xv�^B��Si�t�MZԶ������ڰ)j���̗����Jy3c-l�Q-��{5:�Q���u���
��#��gaZ����ZQ�%f5):���\Tս�%0f�Ugb�b�o1�ƽ����{M�Rծ�ԃ�^�J�čZ��ͻ�$�4�X�Mt(A���4��p�k@K�X��E4�q�mR	u=��;9[������,�46A'oln��-]�8E�t%���-1O�U륗z��U�*⫉�гoran���U�l�3�3D�B�dl�ne'�h����^Zۖ&��,�$	�!�%�DZ2<{�Vm`jh�� Y4h��Q�ź�'n�[,��H+zL�.夎��C��0��x�<�xC)Y�S�7�g]��n��+t�Ֆ�H�U���1점���-�F����aO��-�:�ՠHM�ۧ�F�^�R�4qr���&�ҵ�k+]�ɘ��K�d���I����a��D'�1o}��X��Cp�ay>TA����D5xEK3M8��˙.�XB����k�ժ�\���Y�� ���u������!+]	$ڻ��Z���K6��*��qec��
�1B�^�J˻g^̺cH˥pb�%*��#R�iP2��T�B�MW6�ףQ�*�Ѥic�W1�p:s�$�e�\赃+7$��j�՘��ڊ�ոq�����yn���vl+��.��(U�io%������� 66�-�p�s.�u����v��Vg��k	G�m%,Q���f64�n�Y�Z�n�j��X+�eI �p�Eyj�9yte{����E��cb�w�����ku	����yI�f�6	�>���$n^�"�]Hn����Sj6��/�7)�2�IQ-4lk��H�sU�ˡ[������.4.$�l�]ɒ�-
q��$�A��pZх؊�ө��`J )��/@��"?f�DA�í�U��D��l+õ[X�X�H4�0RC^�B��͠�5J�̆�.��ZY��ز��k.���N�VJ�[M�m��P��@��ɂ��3�,ª�^ hs����ӻ�$�|:ӻՙ.=���â��%CH@�4�K*�ҽ��ȯ(�dg׎��/d����!��dqSQC�$��(�v�.�hd�Ǻ�ƪ�b�CU�ZEyL��t�8E|��A;(1�r�`
7��	(�	KC;�7GඣET7�te�J��ޑ+r�!A��q@�T�+c[�����!�D�wwQ0]B�T��w-^TŐe��o ��Kb)X��`��e�y��|& ���*2�)hO4����-�I��Æ�sZ�il30$/��1�Y�Z�VL�.J8&��b�n��s(�����5]k{�grI/e�4]2"��IY���ėvC�iR���
����M�,YN�ީ���RښM��᠂��f��(a±խ	��fPŰ��vq����&<�K.�ǋ^�:J��F��c�'ʀiv��m��-SN�T����M���J٢���q)��#�^���ܚ�"��r���S-M����_5u��w�U�a-+0��S�G�؍����ɳ��5>9��Q��[�BM��u��̂�J�	��-8ퟚnң�����@�o&��)���L��A����
�ڏU��M��%L��kr�X�.m����K'(��Z*�'n�h@�����75�q,CsDF��dt4��M�W�@Y��&$YV���XH++ Ք��X��Bhݐ��Y5en�N�i��)��Ť�w3���*2�B�k��P���5�X�aгs^^Q%�Mͷ��7�WKA���M�Y� ��<�x��̘��DB;��f�j�G-�*�^.!Q"���<6��>�"ȅ�+kQ�نb�ᙗxki]Y�o���u�-{���Pu�N�Zͻ��jOXs~@V��髥�U2�,`ͺ�Pa�x��@�G��ИX����Z�Tެɻfŝ�V����K�Ʊ���;�� c��0�^ڽՒ����F�iP��̇0�G,N[,�%�m���T�vN\�yb�a�B�CwK�.%��0�fA$�45W�t��6�%�+u�պ��U�m�՗a`�@�M�m ����,E}�cH���͓=��6.�C��VY��h�ƞ�&�̤�f�Ug (�Z�<�e؛�a)��r-v7�5������)��q�jq�in9l|M�]ٓn�dV�݌�ɥ�i��J��pO��sH�l�܂�<�suPjH��L��.�J6�S	md��2��ťd��5�s!���Jt�CqT�l�⬌IM��ɋ4ֆB*�X�h���z���ew.�4p[H+b��kk�;(��䁠5�s+���A�4�m����wg�����	n�����oiY�Y�,'I�L�^S�Wm�f�rۊͰn�����@�#�x"��-�vk�g���ݛ�CR���5h��f�+T�%i��ilnAuj�ī�y�[;x�VXQ�w�G֫c��Z���tT�)m= k�:բ�Ҋ�cV�]�q����ܳ		˦�y�!�����]+�$n�us\˰K��p�[����gUF��ql�S��cn��i��\1Vnѻ�$'��*��4YN��=Ma�֘7{��S��zpS{{�2L�M ��dT�:l˼�vhm;���c�b�f�n�n%mh  �<����zJ��
�Z�J�Z0��������e�˛hU���R:��aJ8ł3"ݺJ���8o4Բ�����9�d�����,��Q�t!��&"�!�����P;QV��4��9��L�g\����V���13���(iʳV��-n���t�h�,�t�EY5{V&[��Lc� �5l@2��MK��ݛb�Q5z(���7hn��x	&�j���6���f�D����=�+��V^��֥�Xh�����*�a=���vw��$`-���c,���&S��=�ݧ�۔�����s��Y\骼�y* l����wK�ޏ��uֱ�n��ꑲ2[��-��҅��Ve��Y�{���D�q��sK��0k��P�ol۸�pU��I�k2;o7I'��N�Q���X�����[r�4����E��Պ%m86B�FY�I��7ww)؇e�#[L���5��V��|��+H���X-ڨ�)��M���L۰Eh�ݕ�"(iJͨ T	jKd���V�Kvǘ%ɃjƲbI\S��e]�I�R#��� �SW[�"+ki;�,���Ƃ���4vA�*]�����(9��e6��ZT����lhy�u����f�ͭ)|eӶ����l԰R�+W%�΃�z�k���*�m�|�yV^�a=}}[o��^&YZ�*K>ҩ��XGʳ0�Q�V�{�,4�ߝ
'r,��'i[WvlD-mI۵|��G8�O����O����$P�U5��
��wuެ�ƥBƴ6Ύ@c��/�kIK�qN���D�M��A���@ek�A��
ދ]M��7]F�x����L��`�i�|�����!�\�$�\�@�{�vl]%��X,e٫������|P&�=ŉ���I�+�(hK��І'�&m97o!�ɰ!��1�V�|�໫�7��oZjԸc���x� �[�Y\�n����D��7��h�N�}y۫:��\z�SD�t+Ze�	k�Nf�e�v�����E��,手T�T�R�ij�܁L�ѽT3��LX	a� Se���q��˼y������������
]\�H.�9+.��[
$%Y�F�L����A�U���
�S0�[�0-Gr�HVØoo�#%+w�81m0��,p�<�M���(%�oh�{�[L��o@�{t.����2���4�/��x�3Q��4t�3n8�YV�Ў�,D�I欦6��;����j�i�i��oyP��9��X���&f�0�ek3f��j��k�[1�L<d	*�SUK�t!ɧ3k��f�H�餂%i+#W�.0�V�w���7j���WZ/f� U�j��ne6_�����z��[������jm
�9�z�m�XY�zS���<��1/�Zq��؛��yX���M&��6��M۳�]�j�^ª��n�e1pݪ�	\(Ǵ6֔�j��f��D�IZ�fh��f�Tn�06��%m�n֌�O��ϲ�.�h�W��s4����"�^��*0����^V�v--��߰"B��b�W+F5Z̕0�i��������/@o�OB�Z�u�Mm+E�|�j�qc�Ya�W]�$�p&gd��jӦ�ĶK[!�&ʽ�8653+35���̔��&M.���2Z��fY{Flۣ2�����4�i�F�&��Ke`GC���0�J+7MB��� �ۑ�yC�����6�2�R�`����xn�Sw�X'(�ֶ,����4�o0���`8ƝM�4v���wC�Ql�X(bMۮ�t��*�ՖH�1�9��y31`cX��,]�G��l�Wj���*��ch��q��X���u���&���˽b��g$�+�ݫh�$9����%�hҭԎ�4���M��j�%��:ʂ�+J����b� �.�8C���K�M�a*z@5�t`햓������r�0��e�L"�;��5[/Qz
�h�0V���[�>�aA�vD�VqJю��Z��tɴ�jS����w��/�s�M��|�V=O�hf*)�e]�ۀ�KS&��.U�×tٵ�0�tܖ3�$WM��q	n��J������uv�^^B��R���ɦ�{c*(�>d���n�lv��]Gn3�[V��#m=�X��CZ�D��?0.��
orR�0e��0��	N�ݥ�f����x�I��T�LF�Gq�6n����o�tkt�w��Be��P�ml�7��ͥ%����;x�Q-ۡe�զ���K]n+�������okAYYh�Ys#�spk�N^��ѹ�d"����p�.3���|�v=�+��.�;�k�`-�
d���/Ch��*�����b��2���fޝ�躺b�{��,���m�B����:�U:x7N&	��\zL�8"]��NJf٢Fn����K+v��2��`b��x&��V�/�% X WV��#݈�W�+���B�PL�=� �]�O"������J���װn�[c2�T����-8n�	Y�yA*���9���;;���n�8s0��K+�ͭ@�P���H���@�H	������mEt,f���HIRhU�DsiC�J�3/)X�x�/��&ɛ��d�+J��7�pQ �M���_[��Z[tm��I���g2�,Ř�
i0�]0��Uҭ�n����%V�u��T:%A�t�OVh�^����-������Z�ゖv�쵦Ȼ�#��d
��`���*f;�b�q����7[��/e��bn�l�Yj�����3"œb�I�F��t��#E�դWS��i|{�]��6��(�e����n54��:0S�	Dᗑ!IP�YZ�P��rݱy������k%}�s�z�8h����y�����%f�f��˦�x�Ͱ�ћ�l�kcj6^Y.�e�ob�4�լVQ�F�DCY,h�&M�n�,��ඉ�v�͂ޓd|-IE��ـ�?Z�GB֖�)�SI��q�>�0�����P{ݹ`,Ra��nnhSY�S���k����&��5�:)�t�f(��y{x%&%����#nݸʆ���K1ј��-��XU����3F��ۚ��uw��p������vSꬣ���]mԥ�j�QO�d�L&-#q9X^^�-�nn�-m۴���7CQ��0}�,�Q���nh%f��8vy�+k�fm&�I�"V�֍�Z����ۊ2�4��ۖ� ʵ��,Ě�%��N���a�D}/2�T�[�X�4i��e8,[�v���:,"/�=�m�mm%g��z��~����W�&01���fM	 �h���x�(�P��I@�@v��D���Pv�'�eJJ��x�2VԚ�R��B�D��Kp+2V��yB��b�.f�^�8���9m�iJ����&��&�r:,LŊ�;�>�F���FZ���꫚v��yE��x ]-��G�}/�+]c�k&f�Mn�r+3n�/p��{�l��1a׻P��r�C��vK3���k��n��T�kwx�#��
o.�eh6�Z�l�J�.˼NZh�j�f]�1���J���F���@�U�E%v/�!�P'y��"�g�6J��n�*�^f�9,Qt�R:��@�Zkt]�1��άi�y���XQ�rL�0��6�yս��a�y[ٱM�t�g]�ø,Mo�2�.��+x��/�p��ܫ�2m\Ŏ�}�����,�:��|��1��Ւ��1u7`{��2L��[˨�WK>6zp�Ig[�3��|�u,�c����<�o�om�1.�yofտ],0Uv����r馺��BcyW��]β�uKd����̷�UƄr�Z[�&^Y��,,��N�ט؏�(,�uN�R�q�����z��^Q������n�L9[���t$�V��/�8*-E�V�+v�[b����#ۭ`S-�
��7)\�F��E��'C-6�d���|��y�X�z���c�J��2]�><5�{Z�Ū},�� Jux�Wn����L�@�'9�"�������b�3>Wz���#Ò���V[HQ�u��5�M�0U�w]m(�o-�͡D>��}�P۬�q�0��:L;��sMK|`qtnl\�6��o]���w���]�H�͑��{]�:�)�+<����n;��َ /�y6���%d�1S�oЩ�ڙ�+iO���N���}b��gd�;��{��"�s�ڼk�d�I]Ѽ���!Z(M%c�
^�{��Q�-MZ�&:�N�]�S�#@�����6�y��@�y��fc���Do+x\<pqg�K2\}����5ѾP���yѢ�*��l�����������;%CA�ȇ�� m����k��W�TF m�.���x�r���.��]J���h]�.�l��߁��*m���*�<�Z��W6V-�����թ�>|��Ey{>�^sW)�+B��pvI��H�ɵ�ܭ�,s�ԭ�\3�[wa�î�gNR��y�P��+R"�*�Sm
M��X՛{p����^���:������ή�e>�H��V��JJRb���=n�X�O)յgDKM�8I���w�hmaǊ��Z�wS��evHl�\��.p�\_,o[U�bһ�R�Ni��f5y���h�nG�K��#b��-��/�J�̭k:gX��s�̞WlU�A��#&�`;�5�dD�n����RP���[J��F����:�Ք��'����mՅ��2�i�w`1��D
Ц��C��KD����YsdRz�KU֟N�0AYpݘ�� �^�5��t:3+�(�P������D*�,u��&���		�o��:�;��쥬�rKg�H:��=f���*7;҆V㞧�VX΍Ň�C���Ҋ�]���k˵+�G2�BM��Q7��u��x�ZJO�����V��4o��G%}B�H���V���2�p�Ig�g1»�O)֭�'����x���!9x��_k �Vn�e��D���J�kl���>4�%��L�]�E�0튣J����@�����w�'�,M=��e�ҭ�Bp�=��Ѭۛ��&��n��\�b�C�Z*��I�W�oU��®7��c2��Oo:�0������A��3Nj���nWK��8o���N�vj
�r�C^v�ڋ��ėIMb��yFH%:�,AB��B�4ƃ�Ue�5*!Žv�
�i��l��-g�i��YO��T�T{+�陸�v���Z�&�QX�l6`Q�J㙒�޴/���J����]����v���e���0���:�ɈU�O���w�n��6�^�lԱD��v�b���ɵ6\����(tǪ�0Ȕ~����f����M[����gˮ���MW�Mz%b�L�w���;�=���#Ʈ��J)v�R8s�)	�mI6ҽBP9�Z]!c	p�Ꙏ�)�{ݱ��5Z.\�@��eJ�t�w8�ʇo]�R����%g�?,�׼��g���u����6���[ݝ¡3���rayL��Y�C�@:�����k���wi���D:���`<��ua��[unѻ/m�4�ź@Ȫ_$�u�1�l�jZ�5��%�]e:�y�����6��ঽ���N�/+������i�,�y^��ͼ���hH���Ȃ@Є�k�<x���d�ALF`�j�dZ��] 5�0��Ы���!C��xwiӑfH��.�GZ;U3pea���f��|�ޱH�I�[� }�md�{�b�7֌�y����r�*!4���fl���'/R�-ULf�F���H��X��X0Ke��~�utw�L�1VMf�T�9�e"�R�ݾ�ۙt�*Ԟsz���]+N_[Ws�ŭ��^�֍3wf��NM��ojz��>R�Y�(�zrs�0��v�`�7��Q��L{l�p�h-���ئ�Ž]�
�9�S�w�d�P
��[��� C;�,\{t�[����	��u�R�1��^��}B��I�U^�=�f
MN��4�u�������n#��×ˠPI7���pR=�m'�)��e�ƹ��d��6h]ȴ��u沱�E��ݲ5n3x���U�n�7NJV�:(�i��Y�j��c�t��.hM�#�Pe\ڇ�$f�Hɕa&Ú��fu޾��w�΍j鮳����tm�R�^ �許�p�jm1�ҥH����A���`��B
\��v%C���@`�\o��ҡ�o3��>�I�+3yQ��gN�5��s��Z72�4�nS�IZ�E��6���-�[x�g00�	A]�SoC�.F�)l�0N�`l��ۍ�+Rt$I*�N<4V4N������4��T=C�&�S�_.9H
�����ə}�hWV;����T �}���#3�K��
+QG��Z'e�]Sh��QV��h!QL��Sմt'�
zu޵��\�I�s�3�}ҵ��;~��c�7����8�ғkRY�EN��7J#�I�.��ȋ��6��1,n�
\T����ٻ�P͜�J��������&nE]�*�][���R���D�K�9���9C�qD��P4Gt��\ۺ��&�uv��4U�N�����b���]-K5��ו˺ҭ��>[�D=tz��Y� ���!�\d�R�u&�0�-���t�8�v�9\I"��hX%�В�y��f���ep�p��(3�YBV��A�(0u�x�b{�lгD�[��데�x�L� ��0M�rAsr��a��/M2����:��x�y^��f�x�l)�ژ����E^���p3),ꆅkH����n�֛�b�bΌ;�;ʲ�7��B'�[Ŋ+B�w��pX�g��&�S{�0��08i���t���u�.�Ӧ�ݗ#=�2%�l�Q�{m�Jv���f���>��5�p��F�f�����sQ ׷c*J���z�'V�=��&8)gB������ʕkJ�2�T����ڬu�����q���i�@t#-��c28 ���8��2�N������J�źt�g8f���W�@2������PƊ5�p6�NP�3�b��4��7���j�\D���f��k�!�R��J��Rs���j�g]���R�!Nh��wΠ�)o�WWS�� "y�X�5u�kŮ��枾υ�\��2;�!wF;rZ�چ�4;����Ҧ��%��[|��j̬D���~��r��?H�����P�C�y�o��t�O�M��o���7������a���lWdfs��7�U�?Cw:�5���s���w��.�i��Jf>dM��n&�%f-mX���<{\�g;��l8�ѭP�Pv�Dom��[[�I��7��Zw�JI���]J6j�@����y�N#{�.�S�n�$�˫��D�:�e�\���dı�,޳b�,�9��$��dԧzc�*�eb��x�Q+b7�C�Ѭ��M8D]���\8���Z��Q�+v�s����i�"Ԧ+�8��1��F����A,���JTf,뙻L嶵7��4�`���S3sD��T�S�l%鷂��y*Z��C��a,�I�Y�U;p�U�aW���czj�oi�=�W9fX��t3C�o�0%1Ǵ.�t7�iӖ��T��s�.�U��E�D�*]^��to��ꎥ��`Lt��u�oVMκ�Y�7ީ�����Ts�<�I&����Ig���&J<ﶖ�q�(t�2Ȏ�w��M����O�ݲ3�8v�k�W�[#���_e'��;��'![��,�ړ)s�8yIYEf�fu��v�M����H��T��q���%��
��gH�����b��Ik�E_r]��&�Ԁ4ˏ'jҩ�͈1��`�sl�Xz
���3ub�)v�3؟p��׷)��vw:iX���	eJ:V:��ڽ����s��	o*Vum�kL|z���u�t�d�o�.t5�u}"J�2��s�Y��W��|7t�T�J����Ք���v)��2�t�C��yW`�S' "Y��/{/IU�mM�i�)�wr�k�;]+�C7��o�?Fm-��"^����I���z!�*J�,��H"BSf;���P^y�L��QzJ��m�g�R3�bf�^.͕��x���i}�B�(鮺�zA7�%IS��`��դ�G6�L8%�'�L� �ed��+cT��Wqf����җ�y�j_v]乔Y�a�R��U�b��rQv���A9���̠]_L�����K�x�0��U�S�e#� HqS�����[1���V���8[���6Ҿ�k�����m���:���;�p1s� 쩝oq�3E�agF���Gd�5� fPp���� �Jh{�aY\R�_��0͝)�Y�]���Zu�Cw�%�qn�=ᾞ��o&��_��ǶV�z`A.�"V�IAt�Q<Kzo��|��끚9�6��Z����##/4���ZL3���fCJK��w�T'^Ѷ��,:�����w�w���gi�&fVd#y�F��P?��Q��_d��7m��7ғ�"����#�A�#6��1��h��p�<�E��B���E�7)"j����of"/'`� �C dnը�N�w���wJ�ӫ_N�씘`闢�C�5�Z�Ď��<=�hE�ռw`]*�!����&.���K�C*������	�|�&b���������Q� �УX�Y�V[Fe�]���z!��SvUMW$��q����ڡ2����b�n*�[��Y��l�=O˰j+#ud,�����l:Kw��!��J�X�y�����zx;�$�H"��6��:^�Q��-�2S,O�����GS-:Ҥc�L��3Z�d��\O�+��Q8���g���A��B���o��nvH�g��=u30 �m⹣k�_#kK;;D��ǎV�pBsܐ�}Wv�%r��^�'W���`R�r�/*�r���b��&W\)���Uʃ��C5eIV�9�|"S��/T0q7������㕋c���i8"#z�ɕ8��|U��������'���!��`_O����N��KV&���bM��N��+-�OJd�^����:�]Y.��E�w���}�d�KN�( �fvNf�,���������C%�Vz�Ք� ��ر˶�=�wݖ-I}89�zbӍq�^��4S����Q$��}�@y/h=I�6#[QS#Vcg��Ɇ�ae��U���Zg]_P!�I;5���f*]w�g�j�;���㕰B�)��#��vw[��4c�#)^|U��Z�e���N�Ү�8�{����$�	{�Z���zT�i�om����#�-�.�(q �����82����l�#[�;-��c U�m��c�2����cR�'}��}�3��)v�<۠�*av�R��H�i6��9��ֱ�8�Ȩ^��JU����GJ����*�!6�̊�왽��\�#���5+(^�Y4�u���,=�l�D0��EL�O���4j�Wڨ��A,��Ll�˹3�X���v����i�p�[������gr���-?>{uGK9Zq���\�����b���s�Yw�5�Z�=!Ѡ������q42�bt�ː��Mh��P9	0as���2l�����]�Sh��t���B��KT�!y�duc���{R��y��>.#�ٶ�.G��+��3v_&�W�Tu5���H�Y��%��]7!u�[ɛE��͡V,�����������Y�f��Q���:��5�д�����7��*<x�S.�r�.�F6�d�ձ���7sy*�/f$�bӋ�.��w�\n��(�P�vvQ�v���(������Ձ	�`��SRN��b8l%<��Q�C��o�Յ��[r�pVu���O-��NQ��o3Irg4:��!�Ս�
�`7��wf:9	�i��gnp�d~G��;sHc�nU͋p�?`|i��d.��}W�6q[0Æ[��CtAN��oh+i:�|����f�Kh�-s{x{7��=����)��� ��F����7enwS|\&'�27���RG��ۋ*B���#K's���t�5���g�[f@����e�+V�$��\T����W���l�B�6d��*�s��:B�f��ƌ��V!Ő������ .���+���O�Q\f�c7�ʖzhIAWG��x���o�`�<g0i0��E�HWe���{i���`�-;���U37ye#�6b�2����O�j�J��ƙ�J@�IX�\]Vv��Mbӡ��j���q�Tq�܇Z�0t��c��8;��=�3Y��6�˹�yM��:��R���Q���/2�N�S���=ƶp|fv�ۦ��L�S���-�姤�9�2MS�۩q�����Z�A#�e��op�=�l�se��{�]o`4��w�
|��^թ���R�vL�r��]���h[w�d^�˵Hrd�]���}�=lW�o[��|�\�w��������ߪ�������]����7����-X�
�}}M�];���
�`�DS(^�7l����7:�JAخW����v鳜8�fk�{;��3�ު�L)hJ�H�.M��绪�ġ70*�K X�Av5]�t�ڻ� OJιtq�Y�G��u��;����3��
ƞ��7�7��	�e;�޽�=IV�\���3N�R��7&s7��������%�MWWwJ���@�Kt�
���.�
ȧ(o嚌�rr�Et���7-�C�z�f,*�c�^�iY
��g��nܝ6ZDR�Z&fut���ۉ�(�rh�so/j����Y�]+.���I�ѷDmު{{ؐJ�1�6Sq))���&�R\��2E�!�O78-}��v���5ibg7�o�7țO����T�5��s�P�#�Cvй�ͪ�X$ޏc֑]@�
������r_T���"�J�}��T{j\v�#w%�Ovdu�|���w#Bܡ��pT�]�fGӯ	仚�{;'��(��y]�'�[�YYƶ��7B�3�R�L>�- Mn�>Tf`@�;�,�yMV�i6��U���%����q�:zni�95R��7%�VZ��ℵ[��0��6��b��Ѩ`��9��|��*��,�ZC�gR;�E]�I�t�L�ܛ�t��$k��<�VH�y횫D��i_��M+{�B_
o��;����-�B�L���_KM��َ�w���{�B`z8��Ɠ2�2��c�$.��lAD90���+Hؘ�S���g���B�m�gd5&�оǯ$;�IFԂ����	��m��.��O��ât&u�n����Q�ۭ.���dY��p��{KamH�_.\~��̙���Ǟm$������ ˸b	c�Q����K�Z��q\�� !;u7�q�l�|#�ՌqE�Œ�3�6S�@�����"ej���h��]�L���H�2�@>چM�f��d=�8� ��IgaNS\�C��ͳ�n���j�	q��m�cOi�����u���5h��ﷻ:� ��^�N�gkA�ҾR랪橪��M7��i�쿍څN�)
&,T�o+was(����<�Νƥu�/@� �f򓚍@C��8o]��D�O�n3&}�V�ݙu�����r�s
��z���N�޾<���\���z*B�n�菊���j���p��3"���t�Y6���r�Ï3Z��(��7iv����0L��&��ܭ��8����
���O�Kv[9R�l93!݀2�䌚�.}gjr ]:�ǖ�J�9ۊ�#Ѷm�|� ;0n�8��^C`�k	�"v������!�Ed�w�mJ��Y�*�[V�xnF��j���]R�=�F�t��9�Nan�����&���.���W��E>�В�i��v>�X,G�jP�J.ݾڷZ��u0��<�0�!u�7+ov�6���N���L^>eڸ���X���f�T�+Ox���]�"�ewx��Gu9�b8e+jK��掽)�<F����b�zt�5����9ʕ�W-�y���v���!
�y�Z��@���q|d��
��y��멞�Y8e5�k�i��L�A�eż��S-�j�u�Q��{Cٷ��L�9.\�yf��)/�R��ع FhU��<Z���Q;��[�ݤ�e><5�5+,-Vd4ftW����,��on�ooVD����3Q�ޖ�v>�F���j9J���O��;.�WTB�p����H�G�N�o(0�8mκQ]tB�����%\ߊ��}F�P��1�`0���k3D*����Y[r��ѷ��Et��b���
�/@��w�ތ����Q�>�V�!W��)�û��:W�lůKWJ7�S�t]t����������2�����uJg�r����ͽ�G�]�k���Nn�C�� �t:,T� �{�kzU��Z��f�I`$f���\ا�6�'�x��d�쬆�o����-}]Vg<ז�s�K��=�B����o%���lO⠙Z��*����ņ���y�VaC�g\��n��v�5�m&v����'r���I_�r�*��Y/�LK�EoL��:Tx��s��p�N�&�S�)�-&��u*�ن
�+�&o��g/&�����{�9�6����_���؎����B����]:VS&��M{��۸�X��q毁�b��%�]�B.P�g���4A�5�.��uuD�����uf�f[˾�3vXz���0�)���(��u��~Ɲ:,�{ȝ�к�\oc1�j;�𶣧��Q��J��6��ˏ}��p.��s
F��Ge���ioq|y��a�ˊ-�JÇo3��A��%Sr����S�؍����b�ܚD�+�,���TlԽ�QF
]@|��Aqv�4���@�]� ��L�]Fʭ[����w�� ��������@GY��!���i��u����Yw�:�c��2N�
�7mZķo�.���mc5��a˔�p�DL7���%����d�x�����걐&/ �c	]ؾ�K���:��er�N��W��
Է*ә��c(��C/JR���FgY*�#w��*���ݝO���(I��c�c �N��u�)>�V��8\R�Z�׺U7DQ��7vۤ]����͞u�K��L�kQ3o/N,'y2�{z9WF,.�4����]��*���l]�r<���x��Z�{/�%C�2dm��;0�=�	b��EZ����o���bnk�kN[�2T���2c�][1��v�L����e	�`��]��m��C�fI������MM����zy�uئgvIÐ��P�t�Ouo�X��Gt�a���Jږ�����anj�G*��p���i�ƒ/r��*QWf��6[g��{l'�f�m��`��ԹSy����0��=��$P!Xb
�L�����	(��:Ⱦ�8I��y���h���f�m��wU�b�k`i(���ヮmԼ�DҡK&kc�����τ���Wp�}>i��v�U�PX/r��}f��wP�P��$���35Y7��t�����w1�+��El����m6��"Qi���Vka%�3�0�3��*d�I�T;�L����W��H�u�vi<�B�ڙ��QQ���i�����x0)�b��&jo!���;s)ݪ'�Jv氥�1�M��Pa����|�q:e1V>�Ȩj6�*�o"�y�
u9�����ဥqY!N��\�h��x1�)<���s2����צT�$��}��Wt���D�]�{���-��Y]�޾�)>�u�WE�el���u+�Y&�Ǧ�V
`Ш��L��`��/�ܐ*��O���^S<�L�@�2�`/�Pb�L¸J���ON�Ҵ5ϛ5�驅P[�OAX`d����A���u�um��:�Ѯ*��K���&��c�+z��e���p´j�vsKy)ۢ"�nRj������X���Պ��jO�:6ud���fM�h���*���Z�6}��Y�]+T�%�X��gw5�EX�Cp�R����T:��M��7��!�n
ÙYNn���
f�D�?e��<�*���p��_p�`���;(�	ݏ�g#i��u��ڳ�o�U�r��VB,���<�v��,�`��d+�Q:�7���fd���ʺ\�d5ڧf�\�F��v���$�!*�_׏yU�c/V��X\ۢ��A���x	���LJ���Y�n���<�z{���ݱ׌P����+GA�18�����xù�g#z�̽��>�`�*��:�{R�28H��-���H��pҺ��p��U�a�r	�G,��t�fU�pn_
j_P���&�H�;��,�"*Y���]G0|m��,��v3HZ�r��`˂m�4_U�s*�}��#���s�o0��D�]]&iݫ��?e�`r����`��»�!4�����d8�sXc�s"��Kf#R���0��)�km�;F̜/v`�1�E�K7ᰠN�V��եyy�P�[(w*�3e1{t�q1���(%ͮ=�M�>�7��d��cF�K�T�-T���2�V�#n�Na�jN�J���5���A�Wb�8&f��<b�A��Pm�5�j�'P��U�%`}�SV��k��OB�q�G\��uj�ZV���w �I�f�qu1�v�����$InV��7뻮L&��esB�5�GK)��{Wwφ�4*/��X١����H��xݽ3�m�n�2i7��)ᮉ�G�β�+x���y��@l����jcܼiq���kFq�֤jVf�Oε�v�w�����c��UoT1�����[�[�F���n����y�F�X��I���5�Rٗ��N��7S�΋�݇+�,XC�V[�jqL����R��9}�t�ev�\1:�#�[#6�L�ܕ'M�u�kC*gA�u��F���#�Z�����,�'mM�l��m�'l{at�YDS��T���ʺ��+Y�!K@��zN��fY�Ov�-Śsd�g���y�o׳����}�i���LY�೛�VJ٦��c#]���[!�}�����uG�F�3D�d:k#�q)}���^�ƆMZ�N˽�����Y�Tt6������W��{�y"��A[{ֈt�p�B�ƫosx�/b�e������׍��n|1&/O9սld��������{�;�i��̲StU9�^�w�*{8/��7z9��49MC*�)E(j[tpi�,���3�>R�t�De0j��ۂop�V6�K��pS�8,�WiSד����������!?���P�ܤ��w`v!A�:r:ق��a��5��wd�eYU,]b��˵���o+����wB)�<b�;�u��7C{oo�h�e��83%	�X���#�I�X���y��3zF�S7g���"ͮ���X�@�ҁB�����Z��`�9ܺ2u'��]�V*��M�s0��tȄ�n7X�6�̩�y����:�J�3R�
�p���7��E^�D_3��Q�.B��a��[/'G�� X�FU����{}���f� ������ ����=��nK1DF.sH�Vk�u�J���]>�Zb4Vgo$�RC M�b�.�[7t8�5&�Ķv�CoZ	�u�GK ����}��v���i�����t�˥�JV���q�c�͙f�o[��1��6��V�(���fUѦD1὎�m���.������(���)�k7�B���r�����V �NJS��茜7Rn��,�r�U��F櫾�I!�T.H�b�&�%Q�i���i�쳥e�9���T��5x�2��Z�v��[����֖�4+c?9�܏��k wِ���5�k�9Z�>��C�@��J%<�︌\@��pb�a<��uj�YM�*���ygf�\i�+�93:l�3`fc'o{���X�͏9&�u���+�'��E�K�M͉m3.�pN)���I����ƛ�p`�C�dq��z�&n���_������^��,�G0�kDC�K�ӚlrR�Uۼ0�r�H��w��,��Ǵ�K�/S߆��N����hqϓ��^�I]@6�B`Z���<:J���}Π8��
��ЙJ�<�m����ݎ�M�s���b���/jJױ�[�j��u�J1�Y�-�Qya�F���$z5E��{jHs9���f�k�^�]���3B�Y������M��UŒ�%�̘�L�q���*�-4tv�)�k�2�l%o�@���QI�C�e�y�Ǩ�G���4E�]��%��.}k�d����T7�����95��n�d�)FП��6f�ES�Md�]í�|�t��k�dC]ۋ$�aGz6�5�:�Y�9�\��K��tQ ʹ��X&�C9ܬ�6�d3���������B���g�喪l�����%�(���MvT�p�7�Ww-�ﲻV�s����#��ݫ��]]�6��1S�43&B��=�o6��0�0.+8N�Vxs����-Ã��W�}
Q|����R@��E����/��SAsI\1�zd�(�V3(X�
�s��wR�׮P�q�ۘt�"�:�K��1(�\3*R��1��F��5�)K����n��>�� �$jT�7de�܊b`�ʾ�}�8r��/�j��έ]`q�޸��������ڼDVw|twb�T��5f�R!Q����ȶ�c��A�X�������9J�׃d��,"�����om�H���q'�~0Hn��>k�m�HprCsFaݖ��R-�KYy�:F�������K9�gS7f�ȑ�qp���"���q%ln�`{��w�2�+ ���e�������i�;q+�G��#�V�b��j�6����"�ut]d]5���T��y)������0��J��*k�B��V��ˉk�9\$u9|wY��'V�W{��3�*�]їu���c4��m���Z3k$���
�	r��v�HR���L������r����[S�e4�{�U
�23�U��-J��R�<��
���{�K���Í��>��A���孑Y�9ǩ�5X@��,,T�̊�Ľ�X�xx:�V`-�r�5�����Xŋ�b������S�V��9:�
B��m�G�l�CE��7V��+��Wb�r���J�\�C������VΦS��)�;Wi_S%1or�������##6�՛�,U՛�9QiZ���`�wGAՉ����w{�)��^��^�zA�� ��1>�1-)�ї�n�p�V���zqt	�z[����
���F�ʝ���K��ʰ�9k�;�I�u��l�E ZJ���`�)d7�e��YX\_M{��+S�9m�s�[����_8`O�@�ߧ�}���>���ޗ�sy�����X�	uf���n`���q��/vbX�ʱQ���f�)B�5�d�\��'+���'7w�~0�N��������DY�%�A=���or)�+��� ��#��݋pl�E9��suu��W5}�:'%�j
x�F�7]�����Κ�ˍVXݖf�n�����{v��kĩ���̦���Ǳ���:�|rV����� �(� �(k�}(���)�7�gK'�����8h��X/.Zݤx[�e���Xn�k5ܹ�'��򮋭�.׹�Ҙ<]�vw������:r�5�]���]�.e&ZS,��o�t:᷃��y}1(ktBOX�WP�|�\R`x�N1����u]V�@V �;,�X�蕗�h�Ht+�$V@c�'�5�Mp��Ҿ$S�x2N;�A���Ղ����=ξ��Z�a�X
�t����n'ˣ1.�����M��u���u�l����Pь]�����X;n�(Dk̮O[�i�7O��U����3k��=x�������c�X��m�`Hxn:���h4q:�mh\7���"��M�Y]i���=<�2�@6�o@�%'�=�'���>1F3���Tdc��/r�H��]pDB����KZK/6��3
�L]<�����*��5�mj�Ä����k�t�P���}���=�V�Nre���<�������i	�f��(������(�
 �+,Ė���s0��+,
���i�,̉"H����r�,̢��*',(�,Ŭ�����2� �*��3�0 �$�*�0�"���$�"�����+2���j
"
,��0�*j��	*��30�̪���,$�	�2�3*2�#(��$��¢s3,��#�	�0�30��,��22����*�02 ���i̲��*�p���Ɯ�2� �*f��"���f�rɢ�3
*���31��,����3+,g3�*rȬ̲1�0������ �0�ɚ����#
�"j�(�j2Ƞ���h�0�'***I���
"���������"&b��*�J�#&�&����&��0ƚ��'*(� 	�T I���g�LQc�/v��wpܦ3����Siu�v/�:�IlUҜ�E%�t�V�R3����_]�f�Xgד��;����s�Z����zf�ߺ&9ѭ�����4I���!v�����ao��^�ovC��]@��Nz�u�ug�b��JI�0˭��P���ϝ�$+��%�z����r��Ώ�>���(d�Ρ>����֨����i�.
~��:��"]�X�ɪlj������ܨ.��UN!��u�Z�qwK	{Ȩ�3ɋߧ�" �8ރ��W����+\���,!�!�<CֲU5��Ϭ�_T��������px#"6����U���6�{�68a��&? �9�����c.���۸f�{m@O�c�H,<q����JI˕ש7[G��@8�g��~60c��p�5�G�m:\�z}W6_]��l����F�X1��ڶ\��.^3��Tf���v�ҷ�>��o�mmR��]q�n��:�^q���z���OS�~5g�ߏ�����e8��������o'(z����;���������7��e��=t%u�K�_j1@{Je�����9C�9�������B��]{�ނ�V�e�'�I�e�X�YA|<"�y��w�Bc��]��Y5�j�)8%�.�U���cs�K�؆�P
]@���H+0��iP�X�] Z����i�l%e�'h>�Z��R���kf��7�����>���q�j�8я�+N���,��w�� ���X��c��fU/��J��r�(����� 4� �]�]����ݳ�|�ZG���$�Ɛ�u���CҦ�=�Ay���Z�عȟ�_w����r�y�����(������.���1Q���Nlq��1:��S��z�9�5]f�F�g�9�d�sYk/�D�� kW%�˩��e�9�[�M�����6*uʭSɑ��a��|lY�%��3�՛:�� �ܱ1��=&���w|k���.�3���J�<��ןJ����K\s�����ZGʐ����ls�>lx�ۼN
$��kӕ���*J�EҜУ$���I�R^��i~��'�����b<#��Px���ѰY���gb��m�ⶑz;����0UW��<���Ow��<��b"��0`�u�D�S���S����eC��{۞0�QP���[~�My����-0o�95%�
	�V5�tGWm�лJ�ߺ���T�g��8N�{[�k�7���jЍX���`ռ���I�tKo���袘�,r��y�x<+��n����\-a΂4��n��!"���:Σӥlyz�zӼ��].�f�ψL�
��[7��Dw.W]��Õ#��};&-� Q�[��'�h�a|Ԙن]����v���!ٿh�0�OT$���^���Vw�	��^���{E|����aI���=Y�F^�[LᾯuU%xf�����2��|^ƨ�����^����T��)Q���缤ow/��{��	��_��/:���$�Ϲ��3,S���q=T�����~�Ӣ�����|�X�AC��,j_�P�^
�4=�5?|�|k�2�o�rw���y�o��M��#�}�Q�
��~qz|��RKG��aP���E֟���t���H�*k�ԋ�baq=����N�_]��b��=��c͸,;��ڧq��� WG�gz��]WjF>4&+�H�<���	C��8���K4;�Qh%�0z��yd�k��&���}Y��N����ץ�{�r���]#�?G�9�!2�����|	���n���ۈdp4Y*P��~�S8�Sk��C�e��'9���OE=Yٶ:3	�����������O��0���7���ޡa�[�*�P04<}��P���B��VR�s��F�pi�}+��_���M�N�4�E��Ά�g�%ǝ:FQ<)����儐�-�N�R�j�.���ЛS�v��|�惇--&/{+�f���7�35��j6�Ju�n��[����~\��Ww��J�o�{:�'g$��#�ec�1�\~��}}�Y��H��I��*�K��v�܆���u�W1��=/t��ر�q�$͜ʟjɃ��i9�Uxg�!:�	�p��]Q[�GY>:)eR\=��C>����������5���U"�B�`۔H�|�O�A�g�L�pS������J)�5*z�tA�O�nҼ���q�cL��)�\�Qf4N�2O�Q9��6����h��9$��'�=M�XB��|'�m�{¶�[]�Xxx���
g��ױ�3�����������'�O�/ ��>Zz�6�ݳ��%=����Lg����j���R�vl��i�\�5tP��ml��KV�i�0�%�p��V�:�����{k��R��[$�����7���ݨz���n�w���+L�yD� 7�&+�Y�����3���m��"k��ү�ϱ��I��fX~���=5dBD�e�:�J3��V�\]#l��
S�]�n=b`�]��{�^�}u��`ӳM�m�*�MP���<w&��޺����_hb�O
�j�O;��Y)^\���SCW��xa���ʵ��l�4	�n�f�1۵^� ���O֦�f
�\\6�ҹu�7~W�j�������H+rA�v�!wd�ģ��d�ޜUe�[g6(S�Uň�8dwՓ��E��9L]9q�X�b�DIq�m2��<^|x# #�Q]X�L+㎝Rzj�:ў��O}ܱ�J�W�p�%\���{��v	F��
;'�\�*Wrl�q���T���&��N��~w�������9�ɣ��+x�~�p�ɯ=���
�Gi�<��ߵ�����$œ9'��!}�a���t���撚�
#	�}k�,�t}��]ޝs�>������j�2%07d!��=:��y����D�68'�U=��=/��}��x%[�r.�L�'���>U��$�&<�~��X�;�����f)21)���ro!:z�ׁ�M�ֵ�/nϪ�{��G�g�<��}Лq�u��ϐΧ�u�篱�����g�dj��9�3U����32t-��7�j�C��m.^��=s)�Z&W���|�K(�������q쇸�j�τ)�K����y�����ڪש��O�62�E qmz^Jj*���#�=�u>�N�y�rĝ��M*�j�ږ���E�X����+[���S���+�s,2Zp�{���O�4��r���i�z�p�0���l��̹Q��i>e��E�{�x�}S�j���)Î�>Z^�z܁=���_���{cR����~��0^�C�^��2�I�����^C�6ЊV���kޝpf>kޟSf���ٮ�x'=o�Ǒǹ𖼸
>"��{Yj�o=��~�z���;g��<�,�3j�j�k�=�~���׳b�ц<YO�-���8[�!Bx���5�ٖ�������,}�,�}���@�vϋv2u�\�B�Igtr{-ִ{k�f��'%6H{�8]���d����Y�gG0�
�V0y<�Z�{�o�;��A�}�q��G����f�X�Ja�,��0l�e�v�XZ�|߽:�Y�
SU���@ss�j�Ί_�L��׳��rk=�I*�<�jz"����#�b��܅���L�9�>���E���.�>b��h�;xuv��H��v��Q4A�J�+���WL�r���I�\��m.�=�-�O�Xv�S�`���U���E�<@�2A�)�5�Z�VN�BL�h�wgz�2W���n`�q<1���V)}˱���XAf�U)�*v9�FWb�؃H��Q�f.���`�"&�7�9�O}��=��bd|WZ�n�]7�I!���U�����&\O	�5��)��뿳�q��D����m�����=݉�3�n�_sL/��t����aƆ���gIs��ͽ�Eg��H��gz�f�O;�7��s���H��S��J���FS���4�H��{�5�3�'��A�����˘�tt����f*�N�˞�u�z�x���Vy֮p��%�\�"�籗�L��n=�{e��=�vӟ	x��0ޜvfQ�݆�]�e��Oݻ<*��a�o���Mǖ�o�ۙ��Ö3��+���LV��
�_��ZT�3v�kw������:;�s^c�F_iɿ�j�^�c�|+޻�E.k��i���{Mq\}�|�e���=�N>��hm��7�[��;X�ϚuG�f6��Lz���*�1�TwGǬ�\�X��a
�UW�:aǏ�y�����䩢�v��4ɏ���E�:i�V.�� f*}�L\��hC��oR�Nm��LsgfҼ��uʽ�����'{h�ⲻ�Dx�j�ĳz�[s	̈́ڮ���)��&�a�ְI�0N=�#��h'+OU�-�3w������{�{U���C�@g��;
��;Ϸ���R{/Y��mI��	�Q#�Zb�x� .B9����}=�ן���'9���{���K��=<��������!�.}�����珶`�1�7u����/��φ���������n�?<ڬ�[�y<=ŭ�����̽����o%���{��~	ɨL��v)K}q{VW�x4cZ<#eJjMu�>���݄�#�0�~�Y���h��q�EBT���RF�:֒��홃�y�l7A������r�0��w��f�����Eo�.�3�bw�g�?�S�p�$N-j�G�u#�[��*�_:L����n���3��l��]r[�]<��).�aY(�֡����;�v�8�k�ѫ*e�N7ꜟ��:�ƃ�gޮ΂��{�_�x+�FG����d��i��H	C�7e���a�.�^��$�Ε��-V��jC撢ͺ�J`��\�����v%i�Gx%f-������\費I�o5E�_1����%1˦�c�Ĥ���~�����ޯe���:~���}O1q�`�����i�\e�:�P��������G�m��(f~Y<^��'I��qf�&i����k��'��~rN�^~B��M�I���9�]��ڸ��[֧��h���(w�e�w:&{���A�������W�]������������ນ:���l��,M2�́�iA��vt�����ͭ�g��"�u����m��T���ynd�>�̚D�Kõ�^�t���K˚��Dvݑ[ŋ\#���k�?[t2��cȷ��}�m�dm�2s�ɒbϦrA�w�(ol��?$��x���zTL�=�����ח73��ȵdȔ��(k<z�z����y��PT�2�,v��v�ϥ[�r.�SW�`�1!xL%t�KÛ��_ȦHRM�����h_[����7l��-M��|�TxG|+�u���/5���wCj�m�<��39�7hY�n�b�j��B�$5�D�C��E�+�'%�B:b���
%��撜���(���ܞٗZ$�IM�TJ�D8�ߞټ����k<�o�c�|[����Ƈ�v���MӫE�O��K�?t�~h���*o�\w�vn?wBly�Y'��k�f0W?>�D2��u�sꛓ__MU2��~�1��S��9�s �b�.�"�C�����̕�<b�~��O��_M���C�w���n[�s�����&6�n��.������{Y<�����=��ez��ܩÍ��󍓉>��˯�j����Ⱦ���e}�M�'��X0w�6-�Љ�w�����;u>�+�#Lny�/\T��}��q�˒KҼ�X�rN�u�{�=������!����q�cQ�v�{��:R:5�V�ǰv>K÷�)�=RB�����m��q���*�!lwc�~zd4g�����Q��m���Z���~W�c^����ʰv5U����c�����~�����qmi����B��]-w>v�w����n�,���r'ʴ����.IQḖ�z�ʻJ���WV�M�V(%�KU����	yu�.�YkkmJ�k�'�]EN����0g�],�tv��U��}x�wu��;���Iur��hs�]s�.c�U4��AL�.��X�eu�ڠ��h��L�Ϝ��d� �J'6�v�NQ�ѡ�L�X�ȗư?�g}lƎQ�,���[P4h��-��luX��v6�,��J+{��o��q��v�²�����lSV1�*�i3�Yc�9�Q�����o6��VL�%�ڛ�j2���Q�*��]�oF�֔&3F��ʻ
�%a����
��2�_;֘7���gqb�˹/� ��:2������7�т��N
N�p��o!������}��g9%��t���edm��/���[v	gVt匭���{�vF��O:ѽ�U�:��ә�m�r�f_Iz��קO#Ҝ|e5�nj/"/G_��]�AS��OV)0��Ὢ�Zv�*�Y����R�]���awe���<%�ĥO*�ze�,�պ5�bv@�.�)�Ό�c~}��ܧt�+�h;V�΂��KFZP�<��b����� �&
���=�ղӗ���j�&�n�r�qf�_���o���vN��if��m�RU�m1{)�)�s@��/���n���93���@��ޡ�n�0K��lVn���sr�[�Yf�Gu���Bv]Z�Ɓ��*Z��GY!"n��0��FP�>���V��[��c�SW��-��A9"V�'�]l�R���R^T���g"�b�E��� �j`�s�ϲH�ݷ�T4�gG��m��Z���%N�an�ySB���ev�	Y��+���}���FX�xr�\c��M0*u��vYܜD�����
$�&�W�Gm�l��5��d���i(�'Z�}=N��,��F�W�}��|�8:�C��qW��^�޷P��iҥ�����:8��c�٥V�	��&Ƞ�1mwmN*ɏ��otu4��]Dv���X�j�塴�X\en���NH0�V5�lV��5�vf�*�SV��� �D�9+[�+�؛��uen�͉^��tT֦�:�z��e�C���#*n��i�;֫dO/�V"��SƅB�'&�9��y�>��q�}]+7j�,9z�ZA�.[�Q
�P�F�*&���Yv��������dpƔ�H9�J�5��/j/��*Y�֖G�ub�9u��&smD��F�4�Ru��s*�ܝA=��%�J����{(�TȞ�v2�Mub8vEY��n���&N'0:r\L�M���X^L��
��4�,�j�i��ӝ+3���Y�m>��'^K��!嗒���Wk(���v�WC�˷[��{����׻W	3�&@z����¨û��|g��g��W���DKT��4��PLdbӘ`LRQT�DDdR�f`�dT�fe%I��TUTUYfXQNMT�9RSTQQ	5MY��Y��a�E%-�DdQQSD�eT�A�6&E�9%�NXU5dّU-fe�e�d��MFa�TPU�d�DQAT�T�4�PSTSMY�TPP�$ә``AXN�e9SfVTddU1D��Y�4��$VfE5�ef�SY�f�9fXS�ca�TPD�U34YcX�PDřFfDTTKfV9QEfDULe���QA�1Ef5@QUMU%4f�Va�	CURMAR�L%4�D̅LEEEDIVa�UDTĕA%BMdMLVa�Se1UQXDQ34��H��Nm�쳈�&�[}l(�b`#���>�Χ-;{Wɾ7-l�����b�Չ�E�yLZ�2�ھᷢ�ݞ���P�QƓ��m��{���s���";n�����u�����)S;L1��͎����=@g��y�{-����K�J"�=��R�g���y����B�/�>\g�:n �ٹ�\��3�����37������ձ=�H�B�Y������A���ג�}P{P���-�[�-z�-��O���4M|5�7Nu����L|�rO����4v�v��z1<����v��͋�NM������{-}n��c���7�j]9��l��k���KrV��a��eo��5��묯EG��3""d�u�(�ץ�aw�+�#�s~��=W�9�K�<��ߕ��aƺ�K����pV����-7���
�5�f{��Ɍ}��#.[ã�k��.��f��7�ӽ��m�+<�M��N�5I张�{���s��7���/��D��%ߍ�~j�y�H�2�%����.nmAoK�t�d��X�v3:JC�f]�Lu�U��ĸ �̒�/���Iy�תݻ�=d���r�x�Ѳ��O�룢T}�ܷ(��>"Ӆ�ٗ��s��ԋ;�O5�\*�N^My�.y��a�^��\~&��A{w���c���`�s�
]��P²��/Iً}׺����v�c	PZm��{�5��Ph�#&u���_K����'������8���fgi��z���e��L�a��(S��RLW�[w��^�7��t�,��s�8�:l���[P���iC������m�dyw��b�h���/K�M��c�9Dwz��F�����S29S�m�9��t���]]�;ֱ����VB�t�>���������[��`x}{dV�b�����]m���0�S<�����N��e����jD�nnkŏ9'��h��0�s�(9����ѯ{���`~��v���+��L��,Ӹz-��Z�	�)��h��Y�uӭ{�z�(e���=2-����غ���}��EQ��:c��%�Oį�����[�Ey$����ǹv6�J -��n�E�ӱ3�����S��R��Z��E�	�#Ϥ���V��C�p��eS.XV�Z̛#�7l_vn�$�H�绑��O��V);Wi��Y�z�M¨k�qwe,B4k6��VG]��t��f�K|���\�Cтs��;Je�4��%�-���83��~���G2��c�M�pt�����}wyo>��v>��8|�c���&5w3w(��k�f�-t��{rm>���<��{fUwt?j;��l�U�1JV�p�R�Čik7�r�>ߟ_G��'{{gq�G�쫛㗙�׺f�<���>Mא����k�˳b��;»�S�k_9.����L�ۏ�}ٛU�
�ؿ�z*qg8�#��O۹�����گES(�Z)��Yit��
�ϯ�a?���s����xz?9'y�?!H���o��á�ea�T�N=��'����)x�p���x�S���M��b�Lk�������l��k��d��:�/L��M2�ɲ���JS��̧������S��Y�2�}f�e�Mͪ�cג^�g�=z렫M� ,�AY�@mKvǗ)x-
Q��χ$�T�k�ҥJ����9����WGDy%<�������nE���M��r�����a�䎺�ۯHm�J�u]�GQ���y��J���$�5�ꒉ�˦�%Olw-%sz���=R��;�Y�{T�#��_o,q}C������X�b��E	a�|�L���~�9��w�94_�vEolW>��ײ��HV}ޛ���ca�7���=-nז���K�\���J�_V;���~m󷻶|`��ս���b���nZ�"����OM��d��Vo'dj^�7F��3��h[����>-�b�K�D�-����Y�ؓ�w1\ �|��	�8vX��@q��(⯇�����C�û�{�ry���������FH��M8bY��S��W�z���G���A��(7/��t��	C俍�������\��߸����X���:��w)��w!���~j�ӿNՌ�������u���u_�����&A���r
W#����w!Ѿh<�p�9��(|��μ��%���.]���H�y/#��'!{������%<�=��S�P�����b���������C��.௽�{�pp�z9#�o��q�=w�>C�}���|�K�{޽��O��<�/��>�w��5�<;=�?rA��r~������W�?F���~��}ޏg�y4���%���t/pr�ޞGR�Of���w�|� 9/���u�!���}=�+�g����b��!����1��jOW���Z�+�j�4a�Z�?���.>��D�I�}�_���\V�!�T�
���㯆��v<�����cɞ���D�
��B��' &�������]��O.G����{n�e�u�U�r2���oX��r�����?}�߽����C�Hsx>Y�~��b��%�:u��|����<����d���}��7/#'���p���<��{�������G��3�g����]�η�^����߶}/r�����+�ѯ�\��Ǹ?Y�w=�|���2w#��u��)_z�9/ ����C�G��D`�`}���\�5&N�^���gy�}��~������>�:�?��{?w��v~��=���'%䛃�b�G�w�R�������)���z������Y��:9��u��u��9������?C��y�)��'�G/�y'foO$�ܻ�ßZW��y�r?G���������w44����B6�Y�︁�巣������6��g�}��O��W?h7.�$7�p��`}ϴ�K�9�^��z���[��{y��w?K�δ�+�~��.C�%?A��
N��_k�Ú�?s\��}�������!�>���W�y��M��^]~�n]�Jvփ�w/<��9����u�{}/r���}�[��z��4.�z�zL�䟿{�k���s�����}�}�u�����(g�2_`��;�p�xh�~�q��O��������Sy�܏W�z��O%�G�����O�<9އ�Ծ����u��s�7�Y���}�����˿=����]��J�;�C�P:}ϡ�y.@}��p�ܾG�br�]���re����Ò�[��`�o��_0^s��io��'��?D��[/�~����?OR�4���<�ӝ�)]��ع#���%�2\�p���x~�w/���4��%���}�%���q�컩�7�o{���~�O<é7+����|��x���)�iNA��J�����]>���~���X���y���)��s��!y�+-�5f���{\�vt�ny�-��=j�ZVU֬���� �{�-�w��	��WA(�W:�IDkJ߬R�o������5VO��¯<+V�S��U��!�O�����y¶��Z)B$�Ģ/aۗ�Y�3����&���4���Ar��>G����}��?��ҕ�z���u�\���sz9'$u;枡�&��A�{��_��(|�����p��ޗ;�}}LW�}���WGHYHg~����{�2�}k��y��G����&��S����^��>�}�=���}����>|ގAJ�����;����4���2NϹ�����ܿ��}����f{/�{������w���^�b�w{/#�b}+��u�'R�S���9/P�O���OR�k�h_ ��AJ�z���q��?X~��G�f���~1W����m?b��j�xs�?+�|�.��_��X�w��=kr>�#��N�܏���~�����K�K�-{�z��zއ�0���@_����Q��fo�Ò��߇��)Ͼ�y&�����=��z>����!ט>Y/�w:�}�SѬw+�d~��nG���O��
����?��@6����!+?`W�L������������������~�=��������<���X�/PC���M��O'����c�_##�7 �����,8�+����[����,������w/ѓӿt���9?�y'��h仼��|��9'�����.�|�5֗%��{.���w�~��ɨ:|v�ZQ���~}�O�}�'���B��Z�7/ђ?y��9.�'�~hL������b���ގK��}��}i_/��}iw#���Z\���=.�沈�Ѵ���Z[~�r�<�y���~���N�Ի�kB��_�7�~����r�2C~�䜗�p|s�)������q����o����ƾ��ǈ��[���pL��l��m����}��$�S�a� ���'�r]�A�5#�;��`}?�~�>�����޴K�yy>�2[��%�~b��\��o�ܵ���ֱ=*ܒ/��;T��U����y/��t��BR`)+m�[-��F�c(����N���p�-s��i�iy�����O��Xv3�q��A(�7%�`��0=�G+�]zn�'�n�&�>�U�sm��k�_3�*����cl���� WR�'Q���H�z��}�2W�ޱr
���pP�f/��^GN�W�w��>��;���h>�����փ� �ᥟ�r�ߠ��+�wv/�k�*{_������׷��/�{�z^G%���w�~����zi]���Z\���~�%�d������F#�G��|�}�������3lW�+�$�n�%����_C����J�n��GR�#�oK�O =7�/#�}���`<�����?;�K���=�Ò�.@�~?|�7�����k�gz�e�߃����u��&��s�	^��{�Ҽ���GP�W}���]��{悓�>AO[���ΰ)C������_~��g�J�;����'?m������sX>K���GG�Gr��W��^A��Е�z���y�\��{ǒrW4~�pP�撃p�=愪�_�_�^տ��D�>����rLֵ�շ�ϐ��z�����Z^]�~u��d��{���w)��w��.��ﴇ��{����!rrǛ�ɥr?;ގK�(L�}z�:���s�-����~�P~�q�s{Ҕ�K����~���\�߸���C��?bnW�����w)���y<��7�{�<�����rG��kM���{z�޹���}�Uw_|.��w.� xoz{�r�'��)<��:ג�������#����G��7+�����w#�xy�䛇�u����~��=���ݞs�~���O���� �N�����w�<�s��w�>C�}���@{/���޽��`�d�������GN�ܯ���~�<�~�u�W}��}�߽g�}��=��h�u.�����>��Wg�t��N�oG#�^����;���;���}��ǭ� =�۽���|����K�]��߱�W��a�i`���0󸲊��GV�ڴ7��E!}mz/�^g5Ñ�qW�t�A�Y���@4\9>�鎷^7���h
7��u{�����.��N��trf�Jz�s��' ș�yR$qvb��O)P��ME�]�o�}?���}�9�&~�����W]+��u���w9I��}�`}/ �����������#�9'[���Ԏ��ϴ�]����K�w{��w+�����rpSxJ�Me�}_�쿪��u���M��X���]�Z�r?A�Ԝ���=��n^FBt�y��w.�#���w'$�7�G/�y'i���y�'���"O��ޟ��v����>��~���W���+�Ѯ�9�����y'��bI��N�R�����؜�����zMù�����^w���t�K�>Ƌ����ׅ�r����~}��Ç���~�g�w%�{���y�%|����y	��O#%����C���jG�w���_�>���;���|�~������k߳���n����?}���t�@}9޽����/:�=���w����x�B�?��K�H����w'��=�r�:4b�I�ލ�t���w����}�û�G������~�~b��5��]���o��r=w�[��K�s�'��'Q�;�?GR���o�� �u�A��2^�>������wko��n�a�7 G�~�H�W�>���n�]���ܼ��a��W�o�u/�=���!��9�/#��I�|�)�:����)]����cio�eo������Q �>�aC��?�`C�~��_������,��t}支e����ܛ��I�]����]��f���u/�S�~�yu��������>{��i���z��}�󾴹�sp�?NK��_e���?b;��?>����y.���%n_�o�t�G#�t�;����ϼ�����5�9�������� 9{��oz�{/O;��W�t�.FH��Z_��;5��}�����NK�O�h;���w'�}�>�K�}�~��v�q�?��5������Fs{'A�[��Zo2�e$+[�� t�$��v��o���È��ܜo��5�o�/���Ma&�{r �Gf��8����!l8��4��q���O9Wl4�=\���Uޚ����ى�j�ɬE����Rˮ����}�(������߾�w+��=��;��u��u.�7�J��d��sBP�.�a�]����r�W}>�iy�!�5��\>!��?}�����ҫ'�n~��z7��{�����>ސ�:�pv���#��ÐR����pR��w��w�4%��|����^��K�r���H�y/#�ߣ���}��\�wߝ���|g�>��/����u&�wޏ'�}�����?K�+�h_ �>�G �|�~��w�|��;���7�C�|�����/ =�}��h�<3z.��}���~�޽�թ~�q�X�w����G��z��y����R�hy����V���^��'����W��ߺ9.� z;��}�;��=��vn{s��g���f����C�߀���>���Hty������X���z��J�>X��?���A�]�K�}��7/#'���p��[���W���k�o��ɍf{�.{��x��0�>�$����~��sK�_,��������!�� |�K���;��L��X����V���
_���w�#�Vua�~����|YOݥ��U�]|o���~�w'y����=��G�>_K���/л�5֗$�S�`y9/$��<���22W�9�pR?F�����Ҟ���gn��/��^I��Ue����W��ra�r:7��y'�����/$�3zy'���_9��|����Z]���K��	��'%���3�+���������������%��W��u��p����+��o��r�2C�������}�2^I�����K�=�C�p�/o>����z�ZL��?o��!���;���^��wIf�����^x�|��|������pъ��ԟF�~��%�ܦ����^y��ϴ�п�����{�����p�V�������+����!Vif˭7��j-�g�*���P���F�BQ{3��%!W��'Qܧ����0*�U�ĪZ��"z��.�X��ûF���}��\�w0-������ͥ/r�2\�E\��Փ��%��Xh�/fs��յ�P�-4��I�ϥ�b�zܳ�^@~��w��y�<�^y�L��'���(��>A��
Oـ}��zt`�C��O�������S{փ��`����K�_o\�/r}!њ��ߗ����;��{������z��:����]��J�7և �t���%�d���}��zш�_c��zNY��~i7&_K�;��rW�po�x漿~��������)�ݟi��~6hq��G�@��OR�4�δ �^u�J�7֗#$u��%�2_���%��~�a��!��q�>�~�7������������_y�}�+�z����9#���<����nh�.���|�P~��)�|Ҝ��z�z?J������]���~����.��^~ì�����}u�l�:��=����}�:���z�/r�}�+p�'^��J�d����:�]�OP�
��IA�|���愡�����Џ������}�����v]���������{�b�#�����y)��=�Kܜ�Ͼ��R���\���?>oG �r�x��B{�i���Q�y���$}�|S�s�}K��ߝ�y��\H�^s�.]��t���wy.�X����:{��]�~{�G��{�ry׺C��]�w��/�rN�w��R�B�c���E�LTxߛ��՟���k�Ru.�$���<��_z�J�/}b��>K��X�w��=�܏���O�nG��?K�yν��R������7U���0o'���B7~$��W]K��}���2S��A䜗��|���/_w��|����%�.�X��!�rw+�d~��nG���'�w���*4ul:��U~�-t����|���~��w��[����;�G%߸�g�ѹy.�a��C�.u������K�M�ӬS��/#�c�_##������0P�i+�+��Ò������	�Q3����\J� ̕�"j��&k����k쭧��7n2I�.�G�;�PFD~sN����W��ln=-�y���3TkM!9Ө;��[lʜ�ҶI(��Kϰ*�{L29EՃ8̺�!s^���{c	=���gc��9��eNOn�����$۾Yuv5�ח�F�mR�3�t� B��ϔ'�oMNַ��ݫ����!V:ɭU�}ʎko%:#+H��[�q&�Y ]��j[Y2��;��<Տk4�'"�iqbYo�wk�	+%g�;pGj?���>�S�ެ���]�D���L���6���5�Ҏ�Ov�����LY/Q���HZ�K���=����<�o.��Z�pZr5�ȼ閭�stE�ej�a���K_=�8�m�It6��Ż��63[eC1\���[��L��6P�Z|��u�p�q;Ö(#w����2�V��7��ÎeC�s�R6ܾD�����`��wSP�vR�����{U.���@lW�K�r�{q�׭w"���\e��K1�[�'����2��I}�&:���V��W�	�;����,��w������1��:�Z�ȰpѾ��%�y��y�U�^ul�5�Y.�n�5�s�vФb��F��Et�X��H���1�Y��P�ރ�j�l-En�4Ǝ��fN���-�mnR���Ů��޺L�G�>ce&�|k-V��:��{���r�����ɸ3�9����v��a�u��0�{շ���(���4)grS�7�
zіr�FN���.l��k�Bi�Z���˲�}���$2�i����+�!bv�2�/ �oU���[f�Y$q��\��Cq���K4\n^���ϑ/پ��e�S*N���]��驄o����tWv074���:mg�3�@��yD
���S���6��bSn`�z�F;^p�M�2vЈb�vJ;!H�Ww�d�N��&��{�����Ÿ����3��/�o��-�E �#�՝�&0Јețrh� �o_Pl��j�N��.�.��u4����L���]X�}a˶�<l>Πt^T��3�WwR�Љ'V���l�]����� }�(�`+cxK�F ��lySs�؂p�k2�@�퇣,^�Kx2���j9ڍ}��@�mՌ�=�P"d��<z���J	��uz�w3L��Ļ���6\ۤ��4��.�\ύb���"�n�*m4���b��z3+[o�Xg�X���Q�Q=��!6�Vf��
�P�M���?/�̻��Β0�gJ8f��tg-��X�i��;��KP��n��էOm(qCvy�P;=�;�yPwi�[��:�Abf:�PTw���! �f6e�¶���i�R�֬v�.��.EW9��f!hC��c��0p9E̼���ގ�g'���LHm7���+=-:������]�	�I��I�c��y�G)�������yW{�SX�k�^u�w��E��EfLN`eIKDT�RQ�DAL�TEAT�T�XEQAQ��1dfQTFa�S+5f1I3DTQNfQ�eDERRMTE-D�PD�E%UE�QTMICAIE5IE�Pd9DEEUTDa.Q6a�ET�JRD��T�E��FRLAT�AMUE�c,ED��PUQ�E�PU%QEfdHDLLQIT�4EL�E@R�UD�DTAM35TADE2TTf8U�cPS��&A��)�1M5TQT4��SFf!Q4LRLQ4�IALT5I�MDR��E,DIHDDP�QDA5_w�g�N�V�RV�2mA�Gf	Ǉ ��=H9��M9+��)t�E��lW�n��f%�ל+�������_Z�����k���Y���DG�~��H����Po�&C�������w �5���y'f}����G�|��9'�����.�|��.K����2_��}������f~�5��ލ#?}����m��}���?�=��׽k �^FHu���r�2w�	���c�q]��ގK��}��}i_/��}iw#�����9����5�^wμ��u�_w��qrO%8��d�C��X'�~�q�������#�����ܻ���ߺ����{�d�������?�������/?���k�Ầ��ov��������}�0���a�]����\��O�a�2AI���9/##$~�q������ߴ��~b��Z%ܼ��ßiL������Pc�;s�璞��q���~�?��埿D�a�ȯ��y�B�;]o��`���.��c~|�Ӻ�{�����E�݇_?����9)�u3��C��uN�둞�E�=Β�;��e�m��Z�dJ`n�CY��6-+�]ύ����o6s*
����[��EQ�2��+�&��s�ر��^[��y���7�'l�<�˕��^��Kvm���-��~v���r9��v����Lt+�u�+D�
m��t.�-���.�t'��`�~�b^7�	�v������^\r�ޱX��!W�m1^4X�򒕈/�ϕ�r`��^��5�#X��6�&L�N�Y�Ҽ���%s7zܜ��c}��!�__�\�覯����,�E5Rq�@[��$�K��^S<���n�v����������M9�h���n����M�mS�验�]-�)/Ӯ�[��-�G�jo��L�!���I����������H��Ï���Sȱ5�ࡘ��jY�$w��۾��_/r&�����{�syٱm{C:��,�Oa���9vwc=e�T�\2����Ŝ�/#����������Ǭ_�.�e��ێ�9�w����p���;��`^���xG�$�rՋ5%.��z8�܏=�����e����fq�5
���'s����ʻw��&��ou�9���E�#��k��d���_ce=2y�_x��.�_�|���93[a�o=3��tw�vM������Wyi�|��Nz��.�3�~���_�7��yp�Dvò7����D��=�ه�u+���fZ|�^t�'μ�����_}2LY��Sn�R����z����N`h��yX�:V��s��3)��w]5&��<��_��)�׽GN��A�:���&����ͬp�R�"��A�KL�w���(�N��7�{��^�6sI���[��/0t�%�x��b��#y!r�)N�K���W����JwfIR���w'諭���Ƥ�g���7�N��g�]�'�7>��;^CzL�	�jɑOo^��
��R]*����r��t\h����u�{{�Z� ������`���u9;��fh�7��zܽc�v9_j�53r$u4�=%��;G�㪖�q�1J��k�Q����>�g�u߱���Dsk=2����̀�����;����׽��l�rRq0�����zڶ��8��2�5��s��E}�Y��e��������S�x��`~�9�Ǡ����on����t"�v\��+��܁{��<��[��ޚ��{ɏ���q�tr�:s��v9=���{�S�y鸝�[
�ъ��s���3�=��{�n�q2y��f�8�/l+_ I��A{��;����ֹ��Y98�33�������q�ͯ����z��S����5���䱾�ݛ�������y��Q�(�/)L��3�9f��,�-+����"��ﲘhM����Ȍp(qS�8~O��Ȑ͏;E�qcR�+f�^�%OAŢrG��A�ܠ����&Fʎ�G�Sd�ƥ{g�XCd��vң�꯾���k��ꓷ{x}���N�'��m-o�Gl��m
���DnY�QO�'+��B׻LK���s��9�	�:S�G7ㅋ᳸{�̑�Ǐ�����
������M�e�3�,s������V��f'�<���B��T9���:��0g��u�>Ωޝ����gH.�đލ�V�:���:��`�ϐ�����:{]{7�{"8��aS4�(�!t��Ժ�Z�眓��+�fϽA��B���~y��C���&sQ=ɝ�g���z;覩��h��x�:�o{�'�ot�ak���������n>fH��-�� ��2�D�<�pB���6��噻�����J|�{7��Kv���n�[Vܾt��W[�,�����f�G�H�b�{ݪ`���|9�y黠w-��w2�c��GzV�O�)�!�k5?i�n�a\�����f��t\v9b��Z�Dt"��r̒3�A��ݬ+�7���մ
5��}o)&w��<�K��������pV1;8��s��ǭ�cV4�Z�o��=���u���}�Y�TYظw�����-{�����#��3�S�v�&k�''x�K��̿}��9�ul�W�Ye�LN�f�<���eܘp�D��dh��zZ��U�>H�'���v�����Cy[鏯�h��t5ks�Wv��k��m����N,ϛ�s#�j]�u��ಥ3���#��y���U�}���SE�]�!O\B�Ptx�?t^~B��v�7A�*{og�ݍ�秔�q}U"�5al�:N�\~�N>���m<rvVlވR��3v�_JG/�E]qUkW/�m��L�&�o<�U����n�eI�O���St�mz���󳣋Ȫ������:�XW�=j����wy�~�����6^<}��Du���b�8�s����3���OX:���p�^�u!d�ߘ(�<�O9��t�M����}n���G��Ћ��u�S҄?S�P���֏z�#���Θم7��-����U���%���N��̱����<�U��*҆���_r[�7ٝ5ֿ�bQq��6�.�R��d�2\�[@>��%�MTM-WȭD��Մ��V������en>���vd���gC�O>���	k��o�E�&D����ۜۢ��G���3����oKV���Z�]��}���'��U���%�&�wNw����X��Se���_���4�݄�r<��c��dh&�wp����[�'�\]���h�b��_�}wyo�'�t%-}��6lW�{�큰�w�����q��������Lu��c;8�7��ݞ~~���x�)�zs��_��5�䀧�����1|��U�ő��������|��/r&���ʙ��Ol�b���K��fL��无~��%��ky��e�d/z/�ř�2�9����g����[���j7��ǅGf��'��@z
�aw�À^������M1�خ��2�9GE�(����M���h󽕟E¾���N�uE���Fœ�{�*�$ф@L�˼���9ư�l ������dW��e�+��+S0�����*�o��}f��
���k�q�3ۧ����M]ߊ��-{u�Z�t��2�D�Jq��e�uZ�
@�\t��Aܯ+t�Z^n�MV��9}i�������v��jc��{�/g�|�毚����g��Ul�;ݍ����o���Ky�ɞ����l���>zgJ;������ed�3�����wN;ת[e�s}8˙�[˜/�tB�,y�1{��/f�w���!�ܞ��[X�Nw9�\�/�%�O�'L�u�n�$���\�H����B9���~srS���-�3���Yݍ���wnz�F��{�	�\DW���}h[��}]�>qʸ��{��^Y��w	M�c��9��M_L�Z����V���67��-5`�Z���R����[����l �~96*�xL�ò�=���9RX�~���<}#}��^���wB{�Jr���~(t����}6�{��5$����Fyx�~��M�A��'��L�N����瞜��G݅o�-Q����ǤR�69�n]�|6�Y�Q�0�y�#t�ף0��p�;��3A�ӛ���8R�����;�66��t'VG�w�-Nsdʧ�CJ��&�7c@K\Hz����<�vǴ2�2v��gI���7&s��E�6m_�T����w6u$��W�_W����Ƨs���r��Wg�إ��(�r��ދ_�����x�o�8�ң�9ϸ&d�l<��9��g6m����}R��S�.qz�l�M3s�y���~�3�^�~�my}�hVą?'�a��k���ff��tO=�7��>�����}���ۓ:�W�m�^�_&��q��o��������)΁ɝ7�Թ�txǁe<��g�8P�0?ܸٞ�{���1��/�	�W9��s�`�s�<�R;Y��{<��O<Z��z!U���m���o�L���'؇��$��]�Y�Ns��m�X>0_�cT9�������Ӻ�O{-�C(&AxT�f���ϝ�P7FzY��0X��~�w2������e�	Mכ8�95�E������<�V	������`�{Ev_�<8�|b�U���q�Y�;k}�Zb:���y��CQ�v��d�&�5Ҭ\%[����/�|�"ؽ���}VY{���XV��	�p4f)��Ek �#��r���#f.��n��z���v�+��mB���|>�᝻�������s^	k݀:�p9�lA�'F���ιD�}o�{������A�g�4rC���$���-�8/�952�xL�zH�k��}��	�L����VxR�=)^ݤ�4܉�a��{3��P�s�y�%۝�����_h�t�!�X��c�v��	����0Z�[K��:���9ڝ����cco��}ȧ�4g�k����L~[��>��L�w��Ż��;}
��Ξ�[7�s^|+<�ٸ��ڤ��ȷb����}���?���^��3���W�oWwX�/n�o_�#_,nu䝼��[��Ƹ{��X�+�����ߟ����"�!ېJЋG`��kP{5���A��p���)�zs�zyC���a�5O�)���}�MO���d�TQp��-��gIӨw��ʿ+n:�����ݍh�A�ϗ5 � �ouc�6V�W[�Zgmi7\���hHK�v�q\]�9���H�f�����h�w(�/z�-2|i���wr�,ɻ�_hb*kp=��iB���(������Sh|���iw�5[up��
w�������K�^�]�ο�kT��>1��d��}������i�Ѫ��sPL��ݽ����W3��L�Gq��<_�&|�5˳�<��T�=ծG��Iy��t�>ީ@L;`;"��b�8�s��wl?����~�v������^~�;��5}2LY��H<�"��S�����evvN| ��Ͻ>���[Ǿ��t����qȵdȔ�����d^7;����sK{�`�����V�}߻�R���ϥ��op8+����y���6$����v�2��5�������=�4�݄����^��koE� " X\Z��:8�+��C[Rt�������b���-�v�d&���g�|��i<'7���Á���W݂sʹ���qv��O٥^'��3z���_z�/{_�\��A�zs�����ÍvyO��Ru�9��[��=�Seڋl�J�+T���/�Z˕���V+Q�egf���<:��
YO�,�S�Җ�
[t�V�ZvXy�V���T�-۬��3j=`+����4%�C�U�ڇ�O�6�t[EY�L5�U�j���ĩ]��dө���F�<��ݚ8P���I��l�A��o/��ܹt�/�Ӂ�,A���Y���tEh��3�+͈sEMϦ�na�ܨÇs"���t�=ڻ�S�:�N뗀���z�[�>�L��Ev����ps��N�S�P�q���9�ÚE|��5,��T�m����N޸#wFd�[�p@�����Ғ�>48�q�i`�7E��-EvͰ&��r��ь��#V-�<v�x�3��:�n�K��{�g-D���IS�ǳ�1O��\��ɘ�+�\�ƺ�NcSq���Ge� q2}yٝ4d�љM;����.������Mُ�']n��lZ%n�-�*��v��S\$"�1�k3v��;���љ�� �R��O���X-ѭ�j{Ñ��nw%St��ރ$`��w�:�j_��ko���X5�d��S�hSf'W�]Jk�>��]k.����4�gq��(n���h�����1���޴b43d:�yIh�9�K��E�)V�@�u���L(�n�1���yOZ��}X�����^�o��$�(�E�f[�6�,3��Y&t�L���d�����t�.�+~�i�pئ��D&6 �]y�<�U�8�Z_�ݨ[�t��:���0���jf�ںѧ/N�՗��ɱ��"��йCy]���5ڲc��P^�C�� �����V��L(���2Iz�\�i�e���m���8���L��Jvn���T_HB����L��=��ո�	��Nxn��\�@���(r���af=��,�1��P�cF՛�<�i�xp��c�K�+=t��Q˾�vN�/������=Pڭ}�-9���Y�#���q������r�a���r��`�>q7�p����:��:-���j���6���,��o��>����Ά�tW}2���X6mK��2�o9&���r!װ�ҴL���j��<���eZf`����q�:
1v�K����POcƕP��R1[�<�{Ys�V��ؕV:WW �͖��k���������w59�uoU�M25�.���?M4�Ζ�Z(Q�w0�(��P��)C���K��/�ح�R��jE��[C�^e/���+5���k7q��Oe�TW3r�R��ܮzpu3���W�� �/��-��T\B��7]+�ӷx�i_){l��}7u��:O]]I���`�'b�ɻ�n�Kk6�֨����XNd<���hj���KoL�O���d`᧱�o���if@y�;�G)���
֏:���~��SS�Ae�T�RTUDM$ITY�S9D!��T�A1TCATMUMTS0�UU�Va�f`PQTKBUIT�UPDET�4D�faUM9DJU+IMU�MQEQ	D�KTEM��A��5ACE&YT���A@P��Př�Q5UP��@QL�QE-Q514�QT�LQ6�0ELDE5DDQPMIT�ELU5EE%0Y�UYUT�5MY8CE4QU��E�DQI�H�UTUPECU2URAMR�D�D4�AUL՘��@PRTCES1VfUT�UMPDd�DE�M4�cU%�5�d�5DUYAY%%��5�VNPSM`�D%6a�`a�DD�&NEfd�H#�O�$�A4FW<n�Z������|��:���@�ҖP�����Wj�}%�w[C7�a�ȯ�o�n�iڶ4ٌ�˷3;���_}��U�[�AW�{���N������/r/������������o��W�	�7��[s�O�Wx��c�S~�ފ�Y��edsv���z8������{�X�����4g��5��k�/\A�O�\��N�>�ME{�q�FnO|��F��!H��6�z���b�
��囵M�N3����z}��'U\����S\�Gl��Ъؾ�;}�z�E(��׊d�����=�'yz�i�~{���ŋc���u0���N���v��u�i��%��.2��9��e�ދ&of�Gm��Ť��=/���4���{�=�ޱ�C�@c&?M�������s�s��Q1��p�G�-�;"�L7�t�(t��-�6����&uu��o�2R��O��˔�<ԇ`v"��x��~����B���|��社��.����<�}�|��ssޢ����>����,M��U��`�E"�j��v�U��[ŤeR�P�5���Čz�_l�5Ą�L ���9ͭ��]�K�ϟQ+WV�]�vt�.��es��ӊ�o�2Ϋ�s��������1�_,|s��� �M��K�忇�W5�z:)�`��45�7��X�/O�z�iZ��z�-Jy>��#�e���95	��e�ú�9�=��s��)*=�^�.}���g�Л󒜶7��]��hv~�mC�ݔ���u���Ŧ�ݕ�R�ٙ�<;�L�u�w���s�N�o�^���sӓu�sw�y���r�f/{��(�r��ދ\{�y$�{p��낱N%���Q�����KSG�^�9s'O�m�����0^��t�D%�wʷW��x���I={���?l+~���&�h��
~6��4Ğ�m=��a���#y��������{��Ƿ&wԊ�4�Tߩ�ટ,�)�V�i�<=����Kɗ��κ�f������1U�ܳWg�y���Fr�P��C��
zd*x��@�=s��[���W�ʹ�J!H�O����GVu����gX})bv#+��`:U����V�������7T�������5�����@䛙�dK��`�0[AoqZ�]��q���:q&�:�!��<�Ι�镡����L0I�]����ip{�~o<�m� >��S�E5��������
�k��M�{�7�q�&v�'5"~�������|�=o�k���=`m��/� (s��ˮ?3�g	�Jj�=�t�Ǒ�뵷�\�s��De�dW�x�g���./�����ϳĥxqd��|���M�����<�L�V}3���v"��n��s݇:w4.�AGi�xۮ�_Q~�w�s^K^���E�Sb��u�2��h�}�����e��߳*
���=���d�#�e����W�.$�Yl��~�/TKy��-��0r>�)�h[�����X�v��K���}]�	���׽���Ls�Pv�D�/:D�'�� �「��%�.������B|يܣ�<���U�ʄ㽳��c�Q�ZB*j��q���މH�#��^3%�t6��.^�=|�P�"��lV9��L�.����] �E\Ft�y��4��)zR�^����с�C3}�e�y����tnSW�lMV���VA��A�B^��-d_n��tZ��5�z֤�Cw�_q��\z�۫�*�rt4�fS]�ʖ�A�7�U�I��ʑ�-�����U}UM���=1��c?���j����3�'��G��f�x�B�',frWg��瓉O�x�3������ ��8� n=����=��rî�Z�]ܴ���c��v���P�c��p��/��0��9�߆r����[���d$�+`ۘ]��ro�,��|i��]m޳s)�=��\_yˋIFg�z��׉���(�T���E]m
�k��u�W�I��flӗ���5��:���ݮ�{ٟ=3���:8��� ��<~�/x����	�"�G6ߘ/��ƭ�]�9':�>�;"��b�<��f�^����l{�6�/P��:��y���<��K���<�h�3h���[<ѝ�9:�ٿP��"�~Uk�\��%�v�r-Y2'��2UP�ݴ�u����r"k8�uӮ��o�k�5/�y�W-�����^Y��ֳ/�J�l!!M�
6
��S��f�ZėK��u� 8���=�=V�R;�J��!q>���9��'�P{�k���]K�<��|��+	��K�f����un��$�d�����5f�j��*�ɡ]L(
ͺ�v]�&���z�_�>���1'w1|;}�����5��*{-[�����[���,�=�{�� y|���11a�������u��D�	���Qл������{c�L����{׽�ϱ�h7��t���E?ȭ������L��ݖ#柄f{��j��T~W�x�˙�/����ӑN��A��ݾ�v��˂�n��L[c3�?-��j�py=��2y���לx��!�e���{�
0���v᳾��JXW�]X��{4��~n^�4zf5������3�q�X��3g(��h>���Y~��=y���TRߺd����|����{�H��/?!H����T�i��Qp����<b���IR$�˝e��R��Ｏ5��H����[eT���y�}�ީ��T7���禘���s�7���v���6�zQT�F����O>��N�Z>�O{���q;%T�{�f:��wn�҆��!@{P��%��]nc�6u�l)7$<7�-��<5^�����(U!�G��KN�9��F�z�R,�s�U�-e֧S"� v�(歋��4������������c2u������{�7ӌ���E����Y��Ƴ�!D��ܾ�����#8��t�]m�������Y9���&*Wٛde�ǁB+k�n��[��ϥ�@u��a��>#��/��b'|�^g��{����M����{�t�婩z&�5�'�VS��r��6iۼ�"ڞ�쏳��I�djv:��K��MB`��5��Oe�{�g�A��-�ߧA�ػ��9���2E?�0.��¿�?6��;���&�~�n���нW�+՛X{���ҽ*�l�E �c>r˭�a:P��:	�K��/��s�M�k���kN�E�O��S7w=e��P�t�%�

e��cZ� 3(�ͬ
uju��PM��������&g*�4ϕK��Z~<6n9�Ls��X9u���Y��K���z�x�=M����11�L��r:�?X
=�����uT�ϗ�C�8�vS�:�JZ�?�[}:����������jb���j��R��p�ݣ2�����%#Y��q,��n3����϶��bX,�O67m���v���2��Op���Vz#��I����
���)�-�"79�
F������\q�)5�\=R���U}��Wl��sˤmk���hb���B%�γ��c%u�C���]�������"�ݩ�{N,ǜ�z�*�u~���Aں_��h��ȟs�^^j�@�Bc��|)�u��n�F�z�,*��X����W��M[��$�z	�MX��C�j�aB��i<�Kx�Ԝ��H�7�ϕudl�Ywp�Q��P{td5�M���.u���ΜfǺ���1�{1�{[��v�ZP6��(�[P˥\]�D��Ғ����M�	�FOwd9��7�U��{��Wc�=�f�+�;48�4��rL%�K+��Oɛ��TYP�p���K�����=�e�����zL��T-Reъ%@����W:�c������[��ݦ/ǟ�n�%� ��5?}-!}�?{��=ug��g2y
�a�lt�$�_nQ;�)�魶��,�46�.R��X璽z��"��W�-p�/��0T3�#Y��/�ڏ6K�����}ٵkK�:P�k}�!~��.�+�5)I��Ć�rʯq	�8WU/ Aʗ��U�YȨ{z�舻�t��jC�v����4̀q��Yo8L)n��7i^q#@h���!�!Ü�>��t���Xo-Փ���sOe7��wBApR�Wv��W"��m���4������2��Jُ�2��w�j]�R���O'0o��Y$�d������)>�K[�ݵ����]Q�^/��vΛ>T�ٔ��URʆ�I���Q&{��~���z�ߥ�?��>��Ą��<�C`pS�J��5�̦w��|ߴX�)ܞ본I/���u����2ODN_�	ݞX��T�.!��,���c�1�'6�ͽ|�}�x�Z��Y��|�;F�3Ԭw�
y1ׄ��o_�^).�KE��&d�J��k��N�v8綺���ȬE<����L�wz����rӇ1*OE� �����w��[�MfK�tL�x}���@��E9v3�^����U�[IVL��ט�6�ɬ���e�JJ��*�,�0�������J��0[����6�R"�,���5��-�|���gh��]V�u*�,z�4:�8����J��"ꩋ٦��eى�y�)��%�`.�m�ߣ7��L�f�]AV��:髫�(���i���zz�Y^w��{��[9s�QhO!���=]��|n:ɗG�J��3Px��$G5P�mW1��
���[|���8���=��V.�wsb�R�B��mi��燎V5Ŭ�,��|�����Rꪐ�&u��v��:�D	�U�qH�Ŧ�J��Bvs-��Z����s��^eJ\:Șwv��Ӡ�T�3�ZĬ�KE�#?�}U_W��>���{�?jx��z�����	�X�n�vU�f��<w�<h��Du�Ԡ�{o5�u�ߑ�igR��ɵ�w��֛�a�kt��1D�*x)��eYQ����N�ۼ�c��R}Η%�V��o��h>ʎ{��R�X_|T>�nT�<r�z��i]o-�zw^;�T�xX�b�����uH}n�k��j�;ȝ������"��k���6o��s��Q�=���4��#e�^�53��3��G�o�m���/|�Dp/~��$�&��O�i=K�u@N�২�I���Y4��S�>Y��H��4�V��Wd��䍻����:�.���;����,|৩t�sW�}��Q˩˔�^��^��{��,v��ӱ^�J�|W<\*?e��)=�*�W�;X:a:V�u�����u̜vL�~�#��啦ڿ({�ͻ�{��@kU����=�ҿ�V�܅���iy7��9�b����vl�J�]���2&Fm[�y~2Qk�3Ĉ�ӞD۬��TQ���@��f4��zi�hV,���Z<5J

t;�b�V	�d���.^�̰܎VfJ8����9�-K˙i��SY�[D��W��T�� ]ެ��H*t6f��9��]�a�k��v�T7,tԥЛ!���� ,e��du����2�=1��k?W�W��y������lW����P^(��8K����*�� ^BP(O z����[}�cs���l����3��~��ȣ�ѓ�=���6�`��C�P��A��꣭�p����ٚiuTf���~,�S�S�x��xw.//(V��U;��sj�#��^Q����`�����-'�E3�Z0�=��Y��`U������b���F$���r��1~�l�wٙ.v�]=~�e_�jj�:�^���㼼��]D�NL�mŠK�9���F������=�Fq��f�H�4��w��o~�=r���q�&Y�{�ޕ]&�Bd˱���绋�Cfy{����5���z��v
fvSJp��F��x�%fs.�'�	�zvyt(�~��u�0���&zZ���@�5��#�o�����Cg�IeUyb;��G��k��Ү�~�J�7�zb�pO"aEF��5���E����X:�u��w^_d��=t*���}�F+����}%\A�3�`�8"��o熑��-�����x�K�}.ls.�[�fw&�"f���R ��KQ��7��>��۲����Tk��=X����tW
B���o3����(��9H}�o�<$�b���ס;�:�۹b�S�F�w����m%��DEu]���[:�cn���oY*L�n�Z�OyU���Ν�y�#n\q-V��bybr���X�L�]�F�j͊�͖����+5�j!K{gn�u�L�6��[�@'�	��CoV-k��Դؔop��M�>ޓt��
�:v��l��w����t:�k��}�dʶeh�68`=���xL�rN�C,��N���������Ҳm�\�	�)w]�Z����y%�Sbe�ޡ�D�`;�=��w�Y�@�z�Ow&��*q"���.��2��7msR:�9��f��oN��]��v��$�k�����'�lv檹�o�Zy��I�d����JRb�{�J{��VۺnJ���ts/r�f.7YJ|�$.��z|��Y�uݮ��q���)2�v����DE�hY�����i��bl-�"��6�=r�YcT�Oi�d`p�Nm��ND��������xj�A�HdU8�U�
��q�[��=Ў�G�kr냡�����	mѫG%���'��B{�t.�;��n�}���	w�ؕ�\�7	�q������ю�U��.��������\i�p�]�S(Vs��fH�.pvqC+�n�{��;�`Fs0#��pK/o �i��2��X&TʾH!��2�u�x��o9�g�P-a��,���űĆSNk\t;�ZY�ٷ\&�f�M�R$yvU�(��,�eL�ܖ�bӴ��pqZ�um��.e����n���ǳ����T�����t|�:��w[�{�nEՓ��m�Sn��t�4Z!��Z��X1
9��a�:� .q�1����,Z˻ƣ�7���k�[�:En�O�O[7�s��W$��={������
�u�PGk`����`jV�n�n��t��Gj+Wf��FAS���\{�[�"4U�U"P��հ����1�B��;F�3Nie��x�H������Ȱt����2b}�wS�6g����� �vR��.\��䮝E�`
mH�S����i����ҍ\��Z�k�v�k�mԚ�.ڢ�)��V%0V2���@��j[��33�A�#�U���6m���,���hD�3�cф�q�\�W�!9��Ó����j�]4���:Vl�WR[�p�  �eMw��n�)�_ThlѠi�I5��`E]�
���Hr�RͰi�=�7ܗZ�&I��սF聀��/��=A��e�=�cn�k�J�Sd��{#���aF�r��ѥt�jB��_��u hi�הm[�6W;G'@�X7���<��w^��%�R��N'R�@_G�V�Ձ˩D�*G6v��kW-�Խd�Vn"�]Z�xgC�)�a����`��GG�Ŋ�uUs�Y�C44�eMQ3�@DED���SLe�1��%5Q�4��1MQT�LE�PEE1U&fAL�DL3�PfSE�$P�S`Nf%AQ9�U�M,�A3AQM4D�KQD�5T�TE���TE$TDUECMQA�QD�UEAKDQ5L�UT�T��4AU4T�TU�QE�TQ1�E1D�QATSEPEDHә�E5L�ESTRDS��A-%S%DAIEPAcITMUAM4L�ME4E%�DQ1TT���&D%QEL�I��4EᘑDDTQSPљ�TI1U5%UDMT�M5T�4SC1���0> 
��Pn��2ú ���dy�y�:6�7T˅�I�4��d:��Cdr]��0%�>�0����`��&��	�^u7�  Y��\2�o?�k�u����u�ⶑ{ܺW��US�e�)Ę;�]m8��]�W˂3+99��fM��{֍��1t<��>��<^�Ut���p!Jj{.�n.�e��7���y�������O�*�4ϕK�I�
Ksǃ�O��:,O|=i[��rc�ŭ��L���$�2����Lu2������`(wV{i^��6���U��p�.l�cW���2ɜY�k��w
>8�<���ڷX}���-_RW�s��~��1Τ�z�R?	ַYD���Y�*�q����9���F�ࢇƑ�s��h����B�����C��� ; j�KlT��3�1���nvC�qM��C7�C�	�GU"/��90�\W��D�b���1��-?(I{Td5�M����bg����2�BEu;l����6�pz�P�ҡ�d��8�tEh���c�7�'�kk�<��`��X���w�ML�����bq�>�x�҈�ij\�Kb�.��2ڦs梛[|f�ub�܆OJ�±s��Z��ޥ`2�V��Ȇ�"K<�w���=��`6uC)�+�`:���Se�������V���cm���1Ou��e�sr���Y`�-�fMJ���ؒU�|����ǃ�z�#"h֟��)��٤�j}`��G��õo��)��dg��S׮���&xم��t�:��������:Xr�Og
�`=Z�n�b�IQ4�\��2<�C���!�?x{�N��L�}<��u�� ظI_09G���^�us`�ȅ��c>�5�X�X�塞��U���˙]ç��pc�W! �Յ�\���7� ������u�އ!~�u��qf$Ɂ����V�֖n�;��k�.�oF�e`z"J��":̥墓J��'�g!����/�w�6�yL�ڒ7j<��ݒ<
nϩ<H<������U(,�{R����(���<+%ٷXJ��[*fѨ7�	�+�tJ��d����-	6ٳ]6�5�R��Y��yM���q������c�P��]������{�J��L�|�Un�xM�o0�jL���ď)�{:pczx���z�ǹ�-��c�P����@=��`���v��OV��z�8՜�sz��^WS�ok0�v�c�S�P���`�C��r�f:�����Ynv5��j)��B��LA�1�iu``jyHe�j`Ts8���L���g���º�::{�&��CX�1�!.u�*��D�C�w����oU��c�|-����������g
��+�oejc�,���.>��ᔲ�Y��VcCq��Ͱkͦ���K�w����H�9��X�Q�R���V�.^�X�6;�G�!%|�ٙ���:��_��R'��^Z�y��t:S6���U)4��B��R���-0s�ӉMH��'�q��=9�J���ϧۺ�<ԛ\tFkZ�.��^��x��>���ȡ��)�g%$C��pE�r0��s�䯊ӹZ3�y!}������ˣ�%G��P��=����z���͐��~�*&�랖͝����u�(y�X�a�N��)�L�<|'���>����YW��<�;�kQ�,�G:�z�\Ձ�k�|N����ʼ'��&`쬙ܩ?C��}��H��� �=�P������X�<Ju-_���mSצ��G�l6����gs{hx����
���4�K)�/�P����N�'"�ˌ���6���^�æ8�=k�ow��8�������P�f��w�+�}�9�T�������ߑ�[)���
kΡ��M��OQ��uD3�:ɠ�����^�gv�ѯ;冉�[I��G9Y&n�@��[o4nܮ�dmjW���O�6��A.��E��w��ك�+�N��^�Jeҟ�e��X�elO�{�S�@Wt.u��By����1�u��E*�E�<�wt香٭=렩g-
�n�B���_����s��s��伇�7:�-:�.�t����(�5��OR���颈�iƲcj�l�~��"�/Un+>{=zL������g��B��J�gk�'Ǝ�WK��1q"c)�Ȟ{�2ϽH�ʸ}+>�[+���f�� �~!�CӳӉt�[C����
��n�)�oZ���l`u�މ�	�?��m?��Χ��I���J>�r�
ɩ�|�MOo3	)<wK�l�����l*��&=�p$JV�!#���67����Z�W/϶��۴�*���S�f������eOk���["��+����L�>�S(��m%C;W�}�6��WZmb�l+�Ո�iN�K�0��ù����]>���3���3;��<�vN����}Ơ�B��`��q�<J)>��a�.mCa:���W����sՁ��t��)�S��ޙ��\��q�_�T"H��7��+������u)O5`0�V,��V��Y�yE��k^�HV�j����5����1Qf/�4����e����:���!0��C̋�Q�Sb<�>�����M���A���M��h���*��nc[3;�<e��B��D�+��Q��w�t�>���YL�]���5]���J*]��Ҡ��޵�cu���謶��6䎓��z����uw�5j�7��_�}��<�R�[z�
��L��]htHvҠt�T>��^X�b�&����i8yo����g���w�{)�9��89xx̉i��
q�*%��E�T�_t�a��mI��9wew�(g����ܫ�̩�B��	���H���E{�n���0'2���i���V,�PmI��	�Z��Iy(?�9��ђ�:�$a��0�p�.��+�,� "�׫k��^(6�po3�]Wr�-�o!���pk��V��oo�����0K���J��HG���kL��¸�{������[�!}ZȿW|��f?%���x`@]}���gÙ,�K5�yT��F���gj�Ef�>��%7�7���:}�Y>���$y��5�V������
\Gv{i^��Xx�p���x�9ȧ&6�K�rӢo���6�h��(f(��ױ�c�%��?�1a酿���7��p��G#w�Ρ�� �32ߥ�8\OU������g�Y�(���ܫo��^� <D��}���P���9�:�]�����E�Y(2����E\H�G
,`��X|+�ю<T������*=ck?��0�K\�9�� P�8ܘ�}�m`��8^���)�sz�5$��ʹ�P���k$�ғˑ���̉�S��OL��V[U2�S3p�`諸�s_9J�P�?l"��r�u
�.���S���i�e^���O���Ė�J~`-���.K���s�+ȣ�m�KVP������K9����K�,w׬S�̫C> �-V�/��x�E�JJ���OW{�+>os��*w��ek�H�gk�o%j͉�`~aV2�X	����KG8��t�97�e+x��/W�d���+��z-?-t����㞨Z��ˣa��"ΐ����|:�jO�I�IH��[S�C�OE6�/P�y�G8�L�ug��g3��L(L6NSٝ�7W@-�oH�5��$��ۈPmnq�;�q���*� ��iʊ��b��'\�9�&���q<ܽѶc�H���D�U���������-]�,��.XbU:�O6��~�}N>�h���;��¾�uUc���2���M*5VP�=y�x�7|� v<݉�Ļѱ<��e#;R����#��D7]��}���<��/*�5�"�j�]jZN���kSv�ՍZ�Wn��*��1]�.[�n��%���{�zƈ���N��̡`�\d�u��v��Y����qk�;�U����5�:8��oq��Fwu]5O�26�n�#��;7�W�^^� �������̓�r�;*�ΰxކ�wEfI{��������/�H{�<����6��\�iS1�)�d�:Y>A�;.���8^����{�?P�
���C�y9��Xxz
��Q@h��<���Sڬ辱��!��>Z]Dn�z�!kޙ4��ۮ��zbe����oժ��zVJ��|�'U���m}��n����|�k}�#�z���]�{+0]��Hd�S�P��@��+-���p����l����^s�׃���v:�F
�)J&��06ʑ|!%�fmg�g�ɦ���^=kP�/����m;�x�R#H��>��zb-�}�ܪ5n
�"�)r�������igWӜ�>.���3Z��^�G:6puB�h��a��P[�ʵ:{�j�w�a�]T��fo�e�����>7g�.�(�*�@Q�R�=�=�z�'v7��# �#�$�'��}L�NTE�jX.w��g��ǽdі{}3��Ii�z��\̓9��&t�> �	iv���o��X���>���9�zz���@�1/q���,�k\���2���f���
�s�Б7��D��U����s/;�LI��4#��񾮟Ū��:�Vr��s��Ӿ��Cw,��p�-���4I��C�6v�鋖��m ����G�����X7ijlA������ߤ�[��W'i���s��f4����W���?,���@}����	c�5�ɏ#�7�k��]hx�wR԰�~�xs�.�[�Z��<��@��O�t�gQ�B{7�B3��W>g"k��ݙ}��=��g�P��)˄D(O|�UP�f��N�ŀ%�V�\[Wv�����������CL����vɋ�p��KN�pS���vC(va�4\�+�g�:'��F�xN����+~�+�
Lv3>�*���h�\�����_R9t巃���ɒ�������{��㚬e�9��՞C�Pĳ�����,,ꄝջN(���c<�z)v���}3S!�m#��U��^T�g��?��0�~!7YSۋv������E�;�@����kNz�� *_����,���ͤ����%�N=����_I��vлʢ=5�2��r��ܭ�`L����r��M�tU�߁�pֹ.�Ց���x�ۙ���0�iV�3�˳b:���۝�y]#e��F�|�1�}��[��rу��趥>��/Ow	k��H&�Vs�]���tڄW*�Ҝ�wV̂��Z�9Pv�՝Y�\�T\��5�c#82*�;e�vV/нt��\��~v嬎���K䂎�9�_u���7҆[��`�e�=Kv���}���k?��~��
W���*�?���i�]e�f/�S�}N!�o�~\^^*<Bp?b�e�8�����*���C��T7W����Rm#|\چӭ�-�:v�g�+��nc��ݱ�L7�n�k�����_]��.�X:��M�|']J�wN��貫�{�γ�5����P� 65��E�k���X�b�sa��V�R�[�b���������7�}������^�3���*d��Ҡok���u2�3;)�3��3��\57$�o��}dq����Lӟ�����d��x&{�P#��B�5�.�����>]��<r@�?7f����6�P@>hG)!�󫒸�T+�����y/�˻������oU�n;��V=Uu ����%x	�]d�):�3�8.,C��:jصw�ײ���=��P���/�x_5)�pvf;��ϻ�
�_	.N$������(w���\�C~��tn��:SġyU�7��f����̗��ˎ�C�(����O f=���p[��#(o��߼��g�����:c+�ay���V6�6��1>���W�����X�mu�@N�g'<���P^ڽ̼;p���6��ph��v`nw7��sr��3��)Q��ڪ�i�R7�!}\�{���#9������}��
�;P���q�n��iu�x>���50�U.&)�R&r�����o�f���c�gɟ������$'<���Y��&}�TzV��f\COlW�EY�����~���\/j��yr��|p=�(�P�Q�8�u�ӺU�L�Mb�sll�39����e�#ۅ(���-L˧�k�z�:�c���Κ�<�kuv�}�Lk���n��FeުuL��6�r�(�|��Nzt��]v��˼M�"��S�S��n��ok)�,�Ih�~`*ؼ {h��ev#㙗[J�������X���P��⇺��C�U��BuB��J�������H��Ս�]���`Z��9)��h�)������׌Ұ��C}�0�Z�襁T�������9�/���}Xf��ԯ\#:r���E�?�B�/�]whGH`���E�=���rd�mm��k�X��b���M�K�=�v���8��\��y3�ܺ&>���fZI�����<)���۶.5³��3;���ȼ�����w��k�5ΐ1c"���+9��Jf�Ggc����Ʋ�ec�f��q�ʼ��:�/q�Xl��e��[��X��0����0ኍ:���n�WHX����l�8�&����3v���i�G,O�^q�Z���5��/v�CHccu����7R+�]-Ŧ[��(�ڸ(Q7[k�
�=X��C�E�]��8��5�S��_�L��sY%ҋr��om�-�m�qCE]�kgc��N�C��^�b�z��O�\'�[�|z���)l<��Y������#܁q#Yf���*,ڳY�V�&��L�N��(�dg:z(�v]M�o����WYH�Vj9-�rG��7��5��S8�+���Յ�]`�$h�&�I��ygQ�m���c�y�QW����)��-�qn-�w�R����
�ˎv+�M�kF:<���_r-��/�mgd�Z���/��l��%]M�&�l.K,7/J'f�8�
W�-ĺ�
�G�Ѻ�%CpR����.].���I��!].�5e�k���m�ա�����V�S�Gf
�4.�1�voC�z��'�%�y�h/��R6%^ {%�Pw���-�&6��t�c�̮�Ie�,:�����c"q:������-�.m�z��ג�J�ϱh����p�xNd��P�'n�3TwOKJ�wuI�%v/�u��{5���k��:���[��u_ p@�AV$h�:�]p5��]�-�dv��v0�0e�yr�ݼ�t�������Gsz]��?E䢫�k���LN�D*��3�"��ps��k�GnG�T�1�N�`�õ��L=��ޫ=6��X�i	ek�*\c��:ؒ���{�pB�������C��22��1Jtf��>���F�`N[oDp�wiF�`�����G\�.f`��
�� h��j)�x^��JCj��+���7�,VvG�9&�
C���Ʈ�]��,�6$M+���g��a�Dwɉ����2� �
��Ǯ=�6��R�J.���^���#}�.����8%��*@�v,��r-�1z�o2*u�{����y�'�7�}�X	i��^�N�X�
��b�����<n2����ֻF���;.�S$�<w�'���:�fS@d���2�u`�u٣p:��䫟r�R���wQ.��;K�C,��'[�3p�&�E�N��l$3�',������M��7S��GS�Xiu�"�9��L;)i2���C0ʻ���+n�ä"Y4g:��&���xo#-�X��|;�6���tL�{
'�1����AC:�,=O��i:�O���/9�k6�l�s��y.�"��p)g;=�������]�D����j�wK���#o�cK�\�k�u�	�]�t}���՚�Uc�h�
 @?	 �1ELTQUUDESTDTUSL�T��UTAM4UQDR�SE1QEIM�dCU�T�EI4$U0Q0QUE54�Q1�UERKRQ$�DQ�D�5UEQ��A$MUAT�U3TTUIL�SIEE%MUUD��$QTN�5LPQULD�QST�ER�MHEKTUfc5PE$1ERIMTIA%SMTQ0TD�QAEA�E1U&fT�3LU0��VY5ESED4PM%�UT�PSTQCUCT��TQED�DATUM4T1QEQ0TTfe4�DDCA,�QE1T̓EMQEASDQRRf0RMEQRU
| > ������0���%
�{����'$4�;v�j���(J�pxa�)yh��.�T�v��yG������(��ص�|f܉^���	%|F���܆��q��lJ����V�kx<t���\J���M9�����L�f��I/�-#�Wِ�/��.��fC�dvDzz��yt�51��P㼍+��2���%])�E�V���*7ϵ��gEJFdQ���gt���I@wS<�:�09GԞ$w�P�S)�3�� ����^��㯒p���ו��:����Qf4N��2ODM��t��+LH�t�yy:�f��S~��������eO;1jE=�(ឧ�Y�E��y_o��nީ��Ϲ;sͩ���s�f$�-���ө�%p��a�X�x�x�X߾�� �����P�.�s�<z.�QfE�]��tUkWuP�^�C��ހ�{\DhtI�x\�7s/Ʒ/�k{�:=��>�'c��
�T:Zd�"�u�[�pu��|!%.��z{�����v����9S�8��[����T�F�}H}u�S.�Ŗ��;��07RBU�{6F"�G��歚Aȵm��s�'�ƈ���&��Έ�PF�Q��/�̮�߰��4|e�٠^kL*.仔�Eo�I-ʸ�r��л������e��8m�V:�9��8�t���R����&u�9}e}�ވ���'e7 ΍����<��ad�� 6�֔�o���u��Rmq��kV%�,�p���U�ЬGiz�I���z{��������,�qӪzjb�y!G�����u�e���Ʒ�EB~ݼ��3�m��İ���U�C�w��gq33>�h���z��:뜦]�uV��⪯t�/>����n�:c�sR��!���R�}.j�굦p�C��w������ޟo�^M�p���xG(���ּtF��GĴ�{�T~5o���{ٞ��夭{:��&v�[��ܶx�]��.��`���#�"��-4����Y���G�S\��='�ig�:�3��q�4p#e��l� V)x�hLw��6�c7����=͇��VsԺ�0Jo/���0����Dۂ��(F4�f�ɠ�g�m�[G�{�8|���j�m9�۔�VJ�����Ry��N{U�tD�g��zŪ�^�I���ח^��Rӗ���_�{�>��1��]����j�{2���[˕{U����G����ɸj v�o뎹� ��u��E���nm��kx*p�7�z&Ν��� {Hf�R�l8��pE�4��λwq3w���t����wY�:��&#�2�o.4�W�d�3OS4��,K=���]"�m.�P�nsu�����zD��!�;�ɏD�A��3�X˦}��p���0�XC���챺
s���k���)'��6��� ���&&���m��u<�:��6��*�k�t=����H�FY3�^сD$F`�40z9�ԥ{k�pl���� �5,�5�7��6ڛ�5�7�q�a�]�o��)˳b:�3���rr��/ʏ�U�")��2;޼��vL��sY�S��V4����;M��/K1juC�N!�o������xb� t�y��!���׆��we��B�,j��*�{u*`��~Y��������4���)�!5/F�3(<7�}[u(�k���v"vF���&(�y���(s��)ݚ��J{����<\��
������<\[A3-��־a�j��Ԗ^����[~{뎙e���x	��*�*@:$7w@�6���^̃�"��Rb髶�g\}q����RN~�i�v��ܞi���/	��&]���G1WWE��l�78�}�<s�o�p��B�7�[��$�9���,���6�[��-.�}U��Jz:�ҷ_t�"��n�����qK��\�cH�gL�.�we@ƃ�6Q�n_���6��6u�Eߏ)b���[J�$7=]�7dy�ʴs):��ɠ����w�C�m���4#�9�����WQ�����n� g����&��-��7wK �t�E�!:����N��2t�EIy(1*��C�0��󩗪���7.+Ƙ������Ѱ~�V.��W�)l�����t�Iw�T!%�+%h�E���{*?s�hݙ[�DN�&%�T��H���&W���x��:��[��)�W5q-��w~���m�ͦ�V5�`�G��C�;�j_P�@�<Nm��r�m�c��-O$�����XEw�u+��C\�Sۄ���OM9^��;܄ܺ=*��^8{l7�3���O�G���u'CUq���/���|q�|,�WpU��B�-_�gJ%"�g}�}<��|\��J�R�!���P�R�ٜ-�����=��j�P���+��L�7��V<�i�m��U:�I������S����5�}��߰����s���{���Bڇ^_�#
�e��Ғ���Ih�~`l> ^�#�D��x��˻�Lw���_Ldp��7�Y�S���xy#Rdla���3�F��=�0����x��;7 G9��O�yהx԰����Jb�I[r�p-�j�nKPf{W7��F��y\�.86��k-9�CBgE�GN]��wd��;�q0��\���I��o�)��t�<�`�|3��}�w���A,J���W~��z���.��M�9��z�#����3����P��+�<ho���Ը%�C\�/���wN���;���*}��q�Sk�^�G�5�}o8�}~��.��2��4)���7�{������:��2��L�a�_��WK��������N��������p@ٿ�{�{�4u)w��f����Pi�B����q���>��*�V��B��ö��ٙ=�4G�;�e��q�L��F�Riz��J�#�fC�_>�j�qfp���>ǵ�ܷ�˟n&8m���u��Y2���IW�)���\ExU���齡n��ݯO+3��K��ʶ�d����O;ʋ+�L����T����8�\/�󶹩u���g*_����Z�&����A�d�:Y>A�3��Pv��}��Z���C �ރ������%��1ז��?c�k�c�D��-��>�O,��0���=�˭bm]7�����J��$�[�-b����O���:6ފ	�Z���8�������ߕ�:�м�ߌ�Ρ�-�;˯.�ѧ:_=Ԭ&wbik��t�8zH��xT�V��u�R���l��>��RՒ�8�����1sg#���X���+�"^�x��ܒ�]<[��h�z�}j���	��E�(��9�휓�o��ˆN
_H��JK<d�]��K%��P{|D�t�>��/����v���ٺ�xtv�+#P��~���XUf�L�=�,r���A5g��I{�#]�ǁ�f�e��������q3c��1z�XF�\��,��OqCoq�J��-�[o�V��U�+u#�q+}jw��]I��Df�����i���J��M����;j�H��I]�Ӥ����";~�pg��k�p�Ԟ]�8�����t�s�6���r�*�����K���U�}L͜���s�g>�{޿]��\f��X��kV���ё��� �����:<4�hx*m=�D�1AV�2��67�'Ϥ{�o|���<�;�ޝ��uBi�I�(�U3��&Em��v�9��h��#�>�\<w����l����|�W�ʖ���u-K=w�t�%����7�Y-I2�䔈��F��y�g9_���
^��yQ����kί��q=n�Ъx���ʆ��2�����#��Lߋ}��Xe�[D����6.4/0�x�'����q�@������Y��Gh2FC��Vrȓ��-�/
'�1�m���u��3g�b��g�P�Z	�S���Pϵ�ꭿN��mꡙ1�'�p�`;��_��K,�vrS�˕f"���=F�
v$D.HlAU.F<fc�t�M��4-�)8�bNPO}��Z�����<�J���L෵A>�48���K��璖j�O{��="��=k'�p�6�	'��ݭTtCj��p!HXU����>�����d��X����?%;W��C���i���AεA~�x^qp���=�^C껼0�|���I9r��n��S^�||��I��1��̵��J?Ki�V=.l�|�v��wN&��#d����l�Ѯ�2J�.�����n�r����V�Ä���j��
_|���ݻ�QX�`�,���U^&҃��e�r������}{�NP��ʏ���V�W����G��e��t�+�:V"��b��i�]e�f!mN�}N!�o/�e��,�c`�����mno^�l���2���S>���/���[2�=��+ ��a@��	��?�x�}��qA�`�MS�.�ݘ��lR�Ѵh6��n���7���WK
!<ゆ�+���$tZ�q���*�����I��;�j�^́�3]5��X���˔H�vQB�jj�ef��C��n[�5�/��R{��TN��{��k��5:u��6-���*��>S���W'��_���v�����2+��2��Q�M���j�d�%{teOl+cdh�nw���;��"65|ҭ�]tXF��T1;�����u��E�o�/z�P�)�^xu5��Ō���{��ν��T��D�"T ��^����Szw�t�j�ȩ).����Utۄx��G�ry�q�92]�t����@�7,���ʤ�������5�AI�B��vy���ɡ���*�OcU-q�>�l	~�vc��R�8�{Ⱥm:Z<�w�>����AH �P��]9\�$Wo���u�Y��P��P~ ğV��_�{[~�˷ts���1�ө�F���dvR�-{s�d�z��T�߇7��.2��{�#V��"+|�7e֌�8�Ҁ��	�Z6}+P����^Ww��f�7�}m�O����3��g6��p ����tGS~�6�)c���;�u�gBEb�Ǽ����J0{Z~�:3�d�x����T$��MX/ؘ�^׻�t�/=Or
���ݺ�K`����'Jr��R�#�Jcޣq�z5+��Cݒ�_V��9YN���G[D��=�U�_��7fG۔���8��(���t7/2�N�ڭݢy�}1ff�=w�z�I}:]ԅ�b���LR�t�\v����m���r���0��-�{�Xv6�J��\�c�l�~����5��w���o���<j�.����(��E�ߥeK[� Ⱦ:�ʃ�e�~���.'�zȻ�2��f�]^�|�V-PA�&����|O��OR���a���]:��|�F�M�{��=�E�ڊg����)�6�u�a��h�_ۈ��,��%���`� ���{��N��7{��vT�r�s�K.y���jϚ�@�'�`��`R�/q�	$f���/;O��ƀ�Gy^*��3�'c7�_Ӎw+�hw��4�`J��YzHJ�����R�{��];�t5���}9QO׮�y9A<|9�2FL���;�Z���oL���}@�Y�U�S,X��ʙƚ�^��{�����}��Sՙ�o�i轧�:MŽo(�%���4:R$�#��qgۜ|����0OK�W�Pkt��fo]�NĊE��y�|{�fXP���#_t���du/���7��ϼZ��3qA۪��^Y���2��;��8FWBe>����d5�MvG���xQk+��t���'�v'�Kzn·'
x��eftL��ZBJ�z�n܁�	h�DY��5�}�^�I.�#�_^,����7�]�ܹ1*]�u�E�=�D�e��|�L�ZCK�n�hq	Ղx\(L����E����Zl�/�k�-_��v&�z�3|ok`֋�8;���\�^`�r�,��ă��UT�*z�Q�k+܄;�+q=FT�;��~ݥyݜr���Z�<J<_"c��'�&�'^۳�mp�E'yj���8kы�TϓC۞Y(,������Op�^_�(����3ԭ�)9闤ҩ4ܓe4���"E�Ϸ��OUf��v�K=qy�a���Zb����(��[�>?Cy=��[�_�UPwjg�~\0hu����p�|�ᒒᄿ���{����m�`�j�<%ݣ\�=:{9�B��'v��3� ߻�}m��E���ڳe����Bx�99��Z6\��wnFtiUy��������3�qd���٘����� �z����*����q��:<�Q���:�j"Ԃ�}�c�%];4�Fޚ�+��CS�'|]I��c5�w�������� � ^{��3�w���]D.�G�0x���R��f�N�~���W븱��1�}E{�J����m4��s�F�H��[�8�b.�.��-jG��xF���+�9��W��u<��cb�{���Zfΐ��w=|I� T�*σ̓1�0��qU�����ׅ�V��X`���ˤ���j�z�-���q���pek�S{xښ����܃w�A��{�u"���J޸���ӗ�R^��W�����cU��m�Z���P�r`#�C�:V�ݼ�f��
�6r�Euՠ�J��2�;����.j��u���U�\[6jX�K4�U�S��lq����ڍ��w��5A{��G�f�9|�^$Y��_>g�-0zҮpt�u*e╭K�f���(��q�	o9�����ۗ�Ũ{A8P�`��3Ee�RämE�ft[��v't��А�b�gT�BB�̜7���V�W��s��1&ɕ2�'��$����R#Y�4���sE)�C:��7.�n�y�)B�w��B �Y�K\яr�>y���n�C�o�e�ڔ�T@S���]��k�����]��j����znhO0ev����t�zt�'יx�U�,��Kd�Le��Ti�b�j��߰���a�s��Djч �P��[�k��H6Q��e*:	mv�N�Y���o#�z�w�>������\*N���Ȥ(v��k.d\��ʍ���2�so0�R���uZ�A=]��]g*�W#���7���k��T$T��]�g3���'�u�[�����T�ބZs&^��lf�F1C_b�(l�5�t�]7���b��(X�R�e�Wus[�JѳlU۹���|�	��[Cf���˒6eni˛&`7���x�p�Fh�/n���[	���n>�U�%0��sf���V�p��*C�.yZ"ȥZ���1��)�|(�<�D�7�X2�P�J��ե��m=WH������pv��a�[H��Z|r�A�3R�Lf��K���+id� z�!�ieР��#oxk|������ju�+rVҧ֩m���}�(�n���:��SvmTkF�հyG��4�Jf�:3C�{f��֓)L�k�j�X�Te��9��G�`5˨AbkO:�a|s�* {�Fɂ�V�3H��h|���+d�p,�M�P���bg)L� �p��rUӥX%_i`�gK����,���ww[�+oX2�-)o=
�2=�ݻ��a���{0�B��]{��yr`)�3rkYƝN4d�Q��qn�x�T�*M�P���cV��
[�{%���1�JX��c�ޓ�*K\
ҥO���rvO�Ǻ�==\=���$��]���2�eҲ+��.B����5"�%f%@'��-�����+�9��⭾&}��D����9r̅�UԵ$c���ݻ���2��_��Oeㅹ��T��w".���v(���#̰��ն�c{)�)��$�O{�и9m�r�U���wU�"�{^G����*�o��X±s픷��SzN$�Y��q�6�q��<>����3���D�0AUEUET�AMUD4%QQTTD�TMIDQ1R�EII3D�Ȋ*���*�H�h���b�"���)�h&*��*��&�"*����*��j�&�L��J()��b�������������"Z�d��d�"((�������(�JZ
R���������jfJ
�
���ZX����H����������
��"� )����J(�#��������(�r2�& *"���	���&**)���(���
��")"
j�f��J�0Ȫ!���*((&��������30�h���0*&"�������$���2¢*")���**�#Y�ITԕ�3fa�UDP�c�A5���E�:�f�f�f4C5C4LMLSD�TUj2f���(H���S�LL�T�A4�QLγ"����#�@ʯ6�ܢO-�QV����J��xU��D�{}M�4f��ewB�J:y����-�9uF�^`)�Nr����m�S��	!)��bDZ���f���	#��T;�y�J��L��:ч�\�b��dǲf�͙�m1����\�n�b��Dl��k�+�8�M{�������;���A�B5T�<����y��@�z�� yP��˱֭�]$���LƬ
	�[||jws��W��x��^�2����{�:���i���Ω�xL���xXi�o�wE�+wJ�b�����H��<}F�h��ج4�jW�%WuU��P�`��U@�<,�Jb�������ܔ�̿y���z�+cu�3 ����N��෴s�����X��v얻Wm���lj.z��}Z�%%��%>�!>邩y�g 1S��y���s7;�	��s	:�D���
�9Bm������r����>�1���m � r������6̽�� �@;w 8�ŝ�0�+s�T�T�W��Wy'���Y7�A�=I�7:��y��a����WZ�a춖E�jP�����ܭ������r��e��g��$� ^'��`sj���3Nrj���]f���nT%M��t�(/�v�r���ӕ]��������k�y�J��`����\���V&��8n�0L!e[{o�PB`��ƭ83+Fwf5K�rZk ;��ؔ�vSK"/����rc�j^���u���|/%����χ���Z.V�3�Z��Ux�C\��c����w���o�Yd5C�|�;x�Fjq*��'�����=B�?Gշ;��y��'֜�5Eӻ"�v�z���i�*����-����j�K1:��b{h��d�F�u\̈�)����.�vi��^*<P����z�Q��{�b�.�b^{J(��z'½��Lͫ�o��c���-o��{�I�DP-����"��������6UA��η����j^G�Yjs�ׄ��-`0�Wbq�d{�<hk�Z�$X�
��	���R��v��>�&�w�2�
�}0��͊|.s�>�3��Z�]"J��J��(i�g&�\��P>�e��B��<�T�5B4��Gw������2]��j͂X�4�~�s�f�����OK{��6���,��
�xvz%͞M�xk�*�O`j��8P���қ������ӏm�wD��!}��WNW,H>���I^�e�ds����`k��-w$T��aUd�b&���U��H�(M�2���Ea���䢋B8L5����S���.���0践�vS�v���I�7����k��I�Y{x���j�;[�w�Y�z�fE2E��@���ʏycwʻN,�[�?��48q��G�a\��'G��6-�v!�1#�tl�;)]3�]�3�z�}܌�})���̯d����~�I�U����0q�.�`q�LJ�YS���|YG衛a��ӂ��V;R���
���+^�KZ%�7�Hk�
N �@9~u�^�g�ġ��Tβ}�(n(���T{;��AK^��xᯮ��:/��<l��,��=wt���`�����+�=����O9����;��;���-�xf���/��(����MCv�R�k�uy����v�<���ۖt�ۦ���ˈme�G�
L�*Z����0���W���N^��k%�Ƞ�ް�^��bXϧ�xa.��R�`U��vRj-�{JtS���	E���~�ݿ,����>���{�C�؃#��P��]=zS����˖L�a���r�ٚz�2�#�U�����K��競3�Y�A�U��ĤW�ux����x׃��l�y䟼��
$z]�Tf�*M�g�N�n!�x���W��C���3��}��[�&�f�X4���J��K�g�#�z�� ��k"���Qvq;ٳ�o,h�6����uk�cw^9,&.l�|���>�-��i�6�������{�0j�$m�tN^�n���[/JY�"Jq|���Y�)ud�Ő�+��RJڔ��H)#�;��͸N��|��NZr�2�z��.�L]���#0G��a�٨}8������GB�S��k���H�~�Q� 5�N)P��\����ׄ�P��hq9��Dǝ�9޹��5Lߌp�ϲ^��v�+�ɾwD�#���R�(3�]��d�/�u˗ҴL}{�8�)��{Sjye��.6&
���#C�&��%���u-e#��p�>��XT��G5s���<=Xt��R,��1!� rʬ�L��K�E��R��^~W����=�� }�(�ڜ�ū7�<� \�^`�D�\��_��uT�'hǁ��nS���U�b�T��90{���2���L��)�k�J�LƉNd��������Y^L�����y��6��tM�\&{+�;��V�@ub��P���@h����2��խowvP�`��z���|͝W�P�%��[�5/��l=V����z�ЧJ���*t�J\$���ߩ���[-���l�r��)j��Wj�L�W:λ�ŴR���}�l�]X�Y��6�rU�m��ۏ��q�l���c,���tDu9�,�lY�����u�2,�2F8��^S�6iu)�	m�k�44e]kSF%[:'�'l�C�cu�����nV���:�j����]�4lZI�I�z�Ѯ9ǔ��-�	O��t���uJ�wW[�q�XF8��
�2�ӭ*��m�y'����{'���e��ƛF���$�L��xt���ץ)�,v=��T��-��7|q9=�ȯ�U�y��!m�C}�]���N$l=5"W��B<N�0�M���x���g��_xa��vx�8�I�BW��Qt��V5��@x�t��ᛂu�&P����	�y�'%�6����u�c5Π�tZ�*���!�C��o�i�� Z"_��>뮳B�y��;o]̍�O[{�
3n�ʐ�y�Tx��6M�Q�0�(P�Ю�U=�DlyH�="y�͈d�m�Oyb�'��$9V��m�u@�;�UI������k�j����\a�g�u��ߢP�E�NNVu{��A�]KW0Poԁ�i.
��4��^����+y��|�P�&�K]�N��L�X"��1&x�.�U�`��W�����t7����O���P�`J]��A��Z�7Z�3�xax��{Gy��+�SWng	~�Ὓq
���4��t�Ga�jQT3sn�6YA�����E:E�C0ɽ�'��ː�]X�C�����7Z:�eΝ��MlC/$��z�jR���{��cV6�ss�[>8���wP�:�4Ϗ:�0��p��+�ի����\\�qwK	{Ȩ�=��8�����#Q�iPd�����\�w�����ܖP��/I>���¼з=,Q��]�u����9)͏�ˀ�X8a���`y1�JT���	�..�W��<�e���鍲�$��髃#�#����e����rP�Þʃk-b5��-�]�/ԗBq?w���:�wx�+�ͥ�qyi���\�fHث���_��0����{Tq?aC[��t��٤��K����1z�,��X6sS�V�3�˳�#�z�����L��TJ=�������["ì��Uu�����a�+�F(}�m�U��N��ez�������vI365~ou�{uA�v�z(�����Ic>����U�]lʤ��T��ճǛ�UѾ���wy0��fӞ�8�α.��b���4p�2+U�RDsB	y�����i5�ǩ�,4���߼c�p7�pvN(2�iVҮ�/���_|.��Ff��vf⮭�Ez��`��}�ҿ]J�[��H��+��w�Y]��\qJ�C���������[Do��D�Zņ�;�yca���Ҟ'y.���CEɣ��,eHd����fjm������6��K4�\�RQ8�g �r�<��ߓ�{*ru�{#�7�g�
�כ4^�����G9��>�˪�0S��Ų�y:��j�`�bb���xJ�Ph�_��/�[�qx�^a��ݽ̽�EG@��Ƣ^�.��S=�Q(zl�hX�xk�����L�.��;*a�/���w4S�>x��?"YEEk��J��� ��o%zu���XE:Y�Ȏ�{ޗ�n6���{s(h뷵 �Z:3�bS0����ő�J靊�i��aE�t7w�9�<����ke����i���lQkC�O�Wp��T�$"���h������Ƣ�N�>V����f��IM m)YX�S��sPZ�̖�����y���}��Е��Z0�g�z�ѝ�
���0�Aꄐ��zV�����ux��}(�;��)��ׇs�k9AK5Z�8�����\�z���ϝ����$bk���1ݮ���ޞ�;ݖt��0]�V`��R�#�ݰ}�6T�b�	1��!XT����^��	L�:U�fI4���췷t�JѭU��j<�
d�ϯ�d%���3��X<E�Z�?iWc���K:V�{Z\��t�T,]��jw�o;�U�&b+cn�C���-����MB�ӠR��.=�O5;PW�A�;�龺F��l�}�
ëИ�Ic>�Ixa/��T��u�!BFc�os�>��z��;�6���;�tOk�:�_�G��T+��S˽)��KG�}m˝ZĲ!�u�~��0U�IA���5��ԡ'X�\Ok�2��g��uRX���_�yPU$�s�k獿w��>���rFcJJ������6���;��Αs��V0��­un\�n�7�����0$��|�+��mS8�Sk�K����E?^�G���}�(s�e�[Z�����t'�=����J����u(P��\�����ץ�^�hq����� ɋqo6�:z��M;ܧ�&[+��0����TI����(8�8�|5ڧu{nMxl����'Ш�d�D���S?\��:��ֶ�e�fXP��Ĺ'T��^!����I���;kȋ,�}=E��,�>�͸3+�=*Z�>1!����Bu`���K�E����y(��wz�HS�|��w6}���XpwEUH*���H�(,����]Ҡ�X�r�p����Rmu�7�V�/��1;���<���b�T�jH�B�m(hSV�eh+x�%��|�܅��>y��ћ�i��]]�$�;����/��h�u�90����\GE�_v-��*�����S�.�vH��M���2�p�ߝ@���V�Kϻ���w��k�R+��%x&cD��2Hδ�ŏ�"�C�n���={ �}�t��n�����D=�<�P�m���ܩ��V7�7�b�q��o�=(N�R�¢�@��ؔ�H����9�-+��g%���=y�a���Zc+��M�3o'NoT�����W�﩯l�>[-�Y�V�X����K��WU3�\P����vǯ�9W�h� m���k�u+�m?���fz�ޛ�l.�]�Ѽ��wU�Z?Eٻ�u��$aV��׊�k�7��m�ǫ�$�����X��m{�U���3i��&��d��E���;��liJI�K��W��=e8�xT�A7І�x@�yZdf��D�x��\��b�u_������f�_� t���M]Xى@x�qӪOM�6r��~��E�p�)V�y�7�ϭ�>Sg!�7`�ty�*��UqUή]�/g@;�DK�]y��)�u�7�:����#���z�6�Ɋ�f��9�J+�\a_P�ů����!u�;����&P���'ǡt�w2�Y�Tl8�ڨ�����KЍn�kp��RB�����J/2.�wA��;u��+ҝȪt%e���+��s+ԝ�ܶ��@Ո�۴�@�F��bΎ���~|�-�MB-�{�6=Ѳ:�{9(�H�,Ǧbb �ߦT���zׅG=%l2�����Ao#�Jf4y��EC�9�����B3����~���]KW�˔���̠�L���	�a��P*���X���}׺��{��n�ŉ3��	�w�;+>t�u�,P�g�P�Z|&\#��5��u�*�}�:���2~I
�j*R��bP���A� ����֨�H��i�>+oIk4�Y�3w�:i�s���:u;�!A�6"���]>�WrP؋�ྩ1�wU7�6��z�-��Փ�z����0�
�{U��'WԊ�D5������..s�x�R�d��M]���C��������\Sؠ=��v�"|w��P��0�ׇ��7�^�nf���q���Zg������H�����{-��dZ��`u������i����&}��N�7��Y��w� �_�{ͥ(߯L�oo�H�Ǫ3C �s;�FKީu��-���VO{[F�����;����XJJ_w����r���f[��ލ�g�x�ob�.KP>�.�{�i]*]k+!n��9ʛ��.�U&�1mu������(�<�oAu#�3�Bҭ�;%����$�N�������Uv�4*朝��b�_SK���t���)�X*�Xp�u�")&#���Lv:U�w�/>D4�γ��vef�)=��\z���Pi� ��&o����c9��fƭz"\T��$�D��� (0��l�,K���;3d3���c�� '^��\jnS ��2�	vX(u2ҺC���
��"���3����"sb��=K���V�K��$���&��%��uBE���ʸ�M�n�MK��D��8�� *�+Yf�"�"�L�M�]���b�,]/uD8˺΢Y�7��oz�:"�fY����|V�F�YȺ��|AF�Q�	�4���sj�����ud��.�{��C#+n;��p"�sɨU�msъ�W�(������ES�B/0��f��)|M���,��=x�����|�2ݷ\�$f�#V�8��m��S5N΢7�͙ݢ��f�����'����If�a6嵗�α�2�P��H]]�� Q�z`�2�8�D<M.�9��V˙#N`�%L�����ё|�U�ܴ�'%bQ��-���$���Ƴ�����7�f�ê��Y���cX�P�nӵ�eD9gL�w���9Lc�,$��k<P��Moj�˹�9�7,Q�1<��Vs�]z.���b���K��x�7p�T�f�	s7�#�����.�&�\3[��"L�<�}��Ncb���G2�E�����P�9���Z����;w�G��cW�5u/eK��F̢���sYb(��g7Q͙+�٫e����@��Ŝ�4˔����c�:U�&h�WX�h4e�tT��kIŤޘo"(nՓt c] 񻼨�s��.�H��=Pf�Z�:Ϻ�1�ic��U#�W(3�CE�R\�F��y�-��xv�\��ya�|��ց����0�S6�8���>:�K'P�%n�د0�`�K�\Rk��j>9pX4�Eu8�[�1�R�9J5wf��c�#|uE��]_�J>)��8�}�^Ő�ى���`b��wcP��ѹ������=���DUiX�勗���f������K�{K�S%��7{_9�X��5k'd�����2�p�Xv�,�[v��V��ێ�ǩH�n�m
*(M!�z���Y����`�Wh�$>��ƯS�����_Su���X�`TON[Q]�y�ͨ�J�Jԙ���'��S�;P�yb<�Q�<iM�>[h8����pbᕬĮ����`)m�͎v�}�i�1�(��8����J|�{��a��H��zӛ�i)YĖM�����}�1M�4q,	[���p�:�wWp���ࣰ\W:�Z\���Rcf�6��������CV:X֛�/����]�N�6�M�˂kY�:�;��]���ߊ�#�Ȩ������3�j&������f)3j�*"����"s2��(�j�ol��*u�k�"����՚ֲ32+,�e�ՌAL�3	��"��5��MfkYZ�*�(�h�Y�TK4�T�UAT�.UYaEEMf�&E�
b)��)��VUSFAQVa�Y%LT5T�Ȥ��0���h�*�)�(�
i�Ք��TV�Ċ��dј�E$�UZ��V5A$AE��"(�*���Ֆ�EU��h���&(����VUM14DUUQQ4�U��VT�D�YF����(��a�PEfFFEVNS&fUa�EE�kTTMDPQfaLٙTELDUDM$T�Aj�XE!��QCLYe�j5h�+,�hԺ"$���\��30�32(33Z2�bfF%QME������S5�M3ݜ6Z�������s�)�Ȥlٰ���5�&��S]a���c���t�P�)n-�t��lǛ;_��qX�U�h�t:�,0Ej1@s��.�K1a��U��驞z�*�*r8�������Q�tbXϧȪ�G���ڸx�sDH�ew�hr�{�,S�v�>:�.W4�Ъ�W��(�q!�:=�)%�����k����K���z�<�f��z�uԥ<�&W���f}8��Q�kB_��W��"���L�}�
�����c�3CH?P�~Nm�YC'<���k-].&l�fՕ��7���y�y�� g&�uCLͺ䤛�F�Yh�[ZGN�tϧ�g�*��wkf��ݓN�[t�6�Cx�Iu�b���R����b8��Ix��Ve�E���\D��?Fj=�=J�σ�+��x��yȲHC]�WNW,	��y�	�4pE��dʆ��T����9�]:�Fn��8:����!h����ѿ�dvR�gb��fw���伭���js�GȜ
�ylo�o�@�K�R��9e֌q�LJ�^��
a��y�Q�	����� ����J-%�;�H���N:�W��Pɗ�n�J�ә	i]>��fZz.��&y	rWq}0==�sx�����X���#�Z���˘Uώ�0J��|��$5�Uǜ��xB`,����X��1��谝�R���ٵ�sU�����UC��UR���0P_�@�5v�د����~�lF`F��0��N{��	-z��s���ǟ��Iꄐ�y=5�z�=�y��E��\�l=�d�[^�GA����{i��N���J�����9�(���_*$哬.����c��@�Nb�շ��������Xr�:�K`o�M���J�w�,X[��^����}��}/��b�o�a�~��Yo�ŉ�
ý	���UL��j�A-�`�/'��$}X��*�ٚP�g��4տ|��.�ϗO=Xc�u�dyEB��T�ۡJ�}�W�
5�7�zQW�}H��7��l�ؑ��{J/:��瞮�φ�`���Y�hv;Qݓ6��b��[��S�j}[^2�T2�Qz��6'Ԍ�m�5�X�h[��똣C�����V��c���<:|��5�X��-���x��g�mx	z���~Z���d���Uc������93 ���*_ǈ`�W:�(sы�3�56�/T:�&rUF���7��>{Ǩ�x��L���A�i�(��$Q�ѯx���	�Ь�M�~�����فڡ�[`�޾9��k�!�e �äI���(�3m������WYԎT�CW/1pՔ��ٛS`���"7�[e��u��x��f+㖔����/��o��5.��i��;��V�y���&≾t�?q}�
/ν�ݚ/�9b�{�qo�Q��2Q�,��,k�+ר1�N)�ˆ͉���))4��du'��m�^u�3��No@�=b�g��.	Ⱥ�Ş��Y,1*��a��𜥅�IR�K8�t��r����N�h�)�m2)&oW��N�]"�tUT���bLr�T�Y.��Cx���-i{ۭk8�>����yh����
�R�p�Ӄ����&��Mh�tOd]��h+}.O;���a��tNw����;+qJ�/tg�!y�<�b�(�C�^.Zv���[݆{sw��Fwl�l�=J�x��j�/l[��I^>K��U��N��צ������wjnW�d���ͬ����\�ɾg�j<}�L>�2��CUfK@y%IyF���R¿g;�mq-��u9v1�ZN��=�tZ��ٲ3"��ٵ�Wz�N~S`�>t��P[�ih��NQ׫�$ྲྀf��×=NP��׆y��.�jY�Vf�Z��6	c��vE碾�x̊�s��������S�Y,&�Ԍ�ZU�aӈ�%��M5���{׭gD�kp��V/@7�|n����Q�VV|T�����5��H������c������*�fب�/v��QևR�&�*IV;T���j0z눨�K<����u�q#=5"V&���u��ԛ\lj�.t�^�r�{_s�x���k��OAx��*�a�G]4-P�U��M'�C3��hɍ�yM���R��sx��k��+��^��Y�ty�(V����!�G:����Y�D��}�̥��Su�tϲ}�(��s��b]oe`p�.Ŀ#�QD�JQ�\a �.�����9�k���6�q��
�ɬ���PD��2����s�\�ޒ���Ϲ�Ao#�|y�Ͳ��W���îo��P
��l�;��O�%��X��t�gW��es�2�V0Py$ɘ*<3޺�^[t�OK{�����ڪڅ�(y�	k��'e`t�u-\/�1&{¡���t�J��p�toNc��D�B맒B���rI�1o�(y��ϟYyy��)^xp#E��f�{���Eߛ��_P��[��"b 8_z��O�V����v{�@��-�.� 
.v��#�{���A��ud;����Έ�_R6Y@uk�!�Y)��\\;��EL�G
�倨����^�A�O�U���-�v��	��(��ڢ���2�=|��h<-G�8K��k�sse��6����6Q��0ǎ-᧷�o T�t{NYO������@�λ����.�[�z��*����&C��o����!O=�^�S�u�}��R��e�n,,�ΘN�75B��>���h�ШnLJW�i�;lzvK߉]������>��!�=�=��z^��	^:V�gM]�
�����i5Ҥ��/�T���;�W�o�B�m'G>^Zd�}xgH�{q�]�5!ȿR
�}yO��9�^�Xp�č���VW�����P�����S2�H�F��V���W�7�t'ß(�����_��R��U)��@X`��b���6˦+%7[�C:'�73�m^�
�'�����l֝w:�dhtp/O��}U��Q��Tb�:�;��y׊d�l` �:._�y篃��N43�]����q�[I��W#h�2���{��z�m?{���#Pi6U�2)�>�J/L}r� a����șb������X�G��zI��9���"�	�n��T���S,�9�^����o�4uO;�� ��1��-$\*�W��(W\/,[1w���&�F��_��kHs�8v����{P6�v4�\0QUZ��d�t��7���/�գX#�M�J��;�EH�f��V�C�:�/�Ҋ�wL��Jiз5��36�\��]�R��0N�(3�ݽ|��ꊴ���/����e�?�7Rʖ�'N��X�{Ge��;&�Ǎ�L�1ü�d�����A� �5��z�5�B��vz%͞M�=�.���4���q�*s����:����7�zb�p	�K(I5�q��iWi��������,%��8��k��]��>ޘ(�/%�}^pZ:0Kꘑ��!�ʳ�t��w�Un�m�S���RT{����_��ܬ�UW	.N$��,�с�N��ġ��R�>1�w�g]���U����Y���
���<}u��*�Z�B��R�g���~���b��W�53ӟtW����=>��|�\��%�Y��}m��Y)�BHW�ޒ8������O�3�pwK��ڋ�p~;T��ʴd/��Mc>񺩚��[�b9uY���Q�������.:`m�"_��a��,>�؆	Y�1�+�y���"�aI��7�mT>�=y�Ý��cxD�/>��W��r�ף�G�QxX��
ý	���3�Ixa;�У��2��oy�-ֆ�҆��\���Iġ߫�{B:���G����y�q�������˛%ry�;sKkE��n�u�ܡA���Z�Q�y{�M��kuh�i��m��bÃ~K6ȣI��U3Ư֞2Wb,�/�(���eD��%�q�����jYW�l/H�H�K�-Ѷ��{HX��rs;�q�:1��\�FCoG��W��6a�IC�t[5��ԥ�L͈5�{J��
����çW��s�"{�	�Ց�@�m��;��ݹ�=�78И�M�g�N�o%j�x.%��+B$w�5��ζi��A�F�I���lQ���?&l?OMQeB/����T��%/�W�Ws�9����3)�s<s¡j��tu�,���S�S���K�|��ڍ�\~O�I�t�gvhq�9��̗2����d�&&'�Q'��P��gN��z�gc�6q���D?}��R�ټ�C~��;�*Zۗ�|z`�},�=iL��,���uz^>0-����"2q��ū���ҥ���bCN,�����`�{�A[�I(0V޹~��d=�vI����:�W���M�oO�����/|\P�3�`�r�V_(�� W��7��2Vy�g�LH{yUT<��|}�H3B�2��9i����<���咺uP��Fe���\�q�H�;�2O��9�ӯlF쭥�|��dOƜ�O�<Y�U뗙¬I�h��\[K�����e��KL��t}t����Ӭ�Y�J�&��Q�iו��{gp���t%�R�����ua���F!7��=��/��]O/r��w5��[˵g-�-�*���ח%�@��a7��'-.I��*���zS��&M�c��~��B ���w�
�v��m�x:꒼2}IK>��xVYU�bݦ��#�鍤��u��<��P�p�؝Vzjg�n<i������w�ѯ<�kq^���m�N����Tt�P�����^��'=�zB���r�{�=�ç�tp�8���z#Ӵ<�;:=�������\a'>��f���9P�)���[��]��-{c��͋����I��)�R�&�qZ.�4:�8��=�<r]1�.��wy�������J(�p���<3�J3����V��6`J�tꞚ�x�w�����e;�'����G&w�,�	ﻓ�'.��*<P�7B��hUΐQ!� ��N�\}�Κe�	o���S|.^�3_Ϛ�;�������@-#�TW��s�_D�oy�p{�6<�*��V��t����Nkw��łf��P�Kٸ*�K���tk� 1�I�u��ħ�L�V(.#o��s+���ֽ�X���-��d˙LwZv&w;�י�v�.D��r|+�`��f��Af�Y�Vm�:힋����Ӕ�Wc�k��d����%�^��v`�P��*��뼲�w���V�o���.YEu��ΏzsoȇfƘ�'so�f���eJt�p˗�*vw�s��4rus��KlYݑ̋�%]Z�(ڢꥻ��(yv�K@w�;)�c�"��1&{n�yp�=K�%_���{�����<�!(K����z��R�X��ݫ�A�>���n�F]f�zVyz�?S���1=������D�bޢa�"DBݓBp]k>��o��C~{���d��j�F9�I���9:�/<�����L��DN��,��h?m��=L�l�q]�^=�3dl�ǜ]�����]hwJ�k��=��Ç����N����E�p�&�5����s��z���K�1Y��=���Ww��}��i��[�m+�[%�j�F17*v�3\���aF�~��F���ꗕ�O�>0�#)���ot߽�ˮ_E��)jy�1G���⏞f���{�&'<����v��"Ғ��E���NUg�S3Ӱ{nv߰Td�Y��u����kN�hM���G׹9C޿*>(=6�Qۡ�v:��"���
��C�st7��l�8��/��ꄹc}7��yyqx��
�p̪K��S�v!�(�e�;�����o�6��]ڊϻOp�L�����(Nɜ� #U��~g9kQ�={�ޯqQ��i�	�#�z��v��R��\�_�ӺA'}/��sk�����Ηi�ԼLqX�7\���[f���q�
;dl�,ovT8K/-|dJM[ޱ�|6�꧵N�tܣ
���}N.h`�hg\�g��\s崚5[�5�D�,��D�жf�z s ��1��x��Ԙ��j���x����jMӻYy��/��|�#��Eb�31ݗ���`w���0�d�+�=�e��WRL�ۯ`��y�l�P��%@�Ӫ���e�f!�N�M�A����Z?S�������,+��3��d����U��w�3�{���;�!��K�R��
g�;=���<��]�};��[[�8�ݘ�<�V�As+��B��LP�}<�e�"���4�	���v�3�g'����M<]E��:Yu��EIy(1.����ġ�Uq�h�:��VÇo;��*	��+s7﨎C��ooù�u
�*N%�������(LJ�f�]?*3.g��>�X�Q#�q��#�>�ͼ/B�P����/k��9A��V5�X�^�ξ���.�z:k;Y�bL�e�g�@�k*���g�M�8�<|f�����{ۗ�}�kzuб��k״7.}� �!������o��7�'�3���P}�ܡ���cgɷ��>j�];/�&7)C�C��Ϙ���10Q��|����2�qf%�l����k��v���m��Xˡ3, e��6^�"�n�;�̱F�J��(��N���/4�4��Njx+�,9,��=�Q��?�.�Em���?��[��
*�<�Uc��;7K�J�m�5��)�E�м�+C�n��3�/7������e݄��vp.�����+Yy@�W�Һ���P��|3�RoAj��n+�Ӧ��&������"��n��q�Q��c��h�L��Q���q�7uzi��loE�
�������!��V���]djk���n���ch��
t�}���=0멎�aβ&d��\S��}�����}GTO,_�h��ߨr䐼6�½@�[�7� �g��Eo!;��1�y'�Q�1Mw�DJ���(�W	mJ�F��Xk*��F� vK�2�5t�|[��5���p��[=���Ol�l	*Ѵ�bv���d�a�6�_%B��k�'��{�ճZn�.^fg)V6�ou�&�csv��O(��jFV�Ѭ���q�]}[�
f�r��B7���r�J�d��3/� �b���v�d��_�]�Y�ȩJ������5�����y8�QH��j��v�d������i8X��E�oY�<I�邸E��&JP��r"��Y)�ܮ���u�=�k"���ڸ�3�oz)�B"�Uj��oR?>���MG�P��� �	Y3##Dj�s,:��P��z0�9x�%S����f�1u�d�cʒ�,yJm���P�S�E�[�P	@����\�@^>����ځ�X��ݪ�aR���Ǯ�8#$�F�K��z�;�<�Su����ҍa8w5����!+d���<��uH�Q�Σ�]$���s��r�;f!��2���
�W("�pu�}��g��6�iE�����k�Y��h;��([b�o��D�����"30����\3�`�����kշ� ���`�����mb9*�YȊ�Wt�lP���co8�v�"�q�l';9�9B��ǒ�i�	�<�dwoj����4�S����T��䣙���{DG�J@j�.uY�g��7�M�Q=�$�e�V�9�Q�j\��8�8IC+�٤ڑ��o���l��f=��N��Y%ʕ��#Rଢ଼4ޜ�����Y7��l�Ü2rn�U���Y9�u����N��,(A�l�S+#�y�4�ZF�Ɵ�Q�2e���l�Lf��ڻ /j�m����߽�<r��;��#'��,��W^��>�x���M��f�54�C����3�d� �R���o: 2�-�aݶQ��_4�$��[�5�V^X^��m_L�=l�p�xޗ�*����(�"+��UQ5AݔEju�J!�e�dSM��XMUUSQY�fj5��
j#3$���̲(�5��*�rb31�h�&(�X�5S$�fefVc�EY�eaY�XYa�A8XUDY�Yf`fFXDSfefd�SMFAXF0�QAANфDTANFUNFa�f6aQ��f$YV��QDU�Yf4T�fT剙��fY�a��d呆ea�ff��YFa�fQFF9�5��%S�U9�XU�fYe4QYdY�c���eS�dVY��f9RYQ��U��eeaFfPa$I��M��E��UY�Y�a��a��%a4efe�d�eVa�Y�����faVa�NfY9�ad5�QQffN9UX`�9feD�4dfeE���a�Ee��XőE��9�XfYQ���eM��9�K��fk^^�F��.9ʸ;Π�M�z͚�c=B�7��f��*ɽ�Ih��x�=}�Ձ�m�s�nպ�}`&��-���Ʌsm�8TC.�|�ج������8/	T�U�C���^��H�^���l�q�aA�����q���;���;c�%U�f�r��ob%f�D��E�HmvԺ=�K�c�L����U�u~�A�c>Z��mL��?S�j�Qx���q�.��Qͻ�3�6��^�޳ig;�vR�+�8�N]À.�z�ơ׀_�#=�x��8s=��e�{{��^|�� �eJϮ��6>�5	=���҈I�'瞮���Y��&�����bPS�E�A��h̺�/���%Q�8؞�n�O���14���"��Ӓ���l���]�t
�X%��D珧ȭ>k�����{����P#�y=�lM��ѝ~�OG�9ꅪBe��ҠE�x�	<�zŎhb�L���o-]�篔S�y��o��w3�mG[�:⡤s��<eʖ��&s>�D�d�;�O�_Oe*������e�QoIJ�Rr��P04<~��Ƽ���|ejqO,��pٹ����B�M�$d4�7�=���W|L���AX���i
��|:�gYz�D�
짔����5�׼�p>�^�����vQ�~3����4�7H�r�w\L	�Le7�w��ws�{f�ov��,&���gU	 <S-_MM�*��L)�J�����_�����#+8?fK�] C;{�9��>E�`�,��j Ļ,(�`�<'%�0J2��X�s0����˙��k$�U�#�g��E'T�XY���"�t���\�^�Ǎ���Wg����{��C��W�Ą���<���qͪ��^e3���]ґ���	����DL���pM[�ل�Ӎ�u�nu�:�ZG
�R���+���o�V�A���g!I<Zy�F��:gJ���
>{�fbz��сJݺ��"��I^O	�ƺ�6����E����ܾ�kP���q��m���4�d�3ݢ���Ö�s�2�"�)S��9����ՐU2���g��]�kW�â��˱����F��ǫ�*�y�I+��\�{��Q�6Zؕ�C,�0l�"Wb�	5���.)�}�$�4����=e��ݜӔ�D=\V��;D;���)\V�t��)Ď�5"V&�Ջ���T�
Qn��1��l�M�;�f��^gM�}����=�N0���M��u����R�lꎱ�ӆ�љas�#����S�\��%Wk�I%��1o��X՛)�qt��g�m]8��Ӽ\��%�M���tY�7���=��͢gT1����������0���|W�p�XK\�������K��{.K=��6�v�� �����QU�D��U��*��{@]8�����E��YXz��� ��S3g*0�=�8&^���L�WGL��<҈�օ�V:�{�'�u�9��q��B����\�=�|���������b���F,0vV?fe�kZs����>ԁ�KRKi�M�>à���߆q�8�J�=�4�޵�i�Na�I�}��������R`�=/��"�N�kR���@�޲vW|�� b��];[X=;q�M�5tz|��&��S��*���U -��%v�1R�G�;5N��;�Ϳ$�f}�a�.Ӣp8-�>�vD)�6"�����ա)(z������>m�w�Y���눾���c���&�R�&V���8M"�z�o#�IS�gD��=r�\X���&q�Rc�]҆%�

��7uX,�>��CX)�z�'N�;�rsY�6}U3��ü��P�y(d�r�>ސ���������
f����i�/M��83~��Л|�o���*�ݳ��ʜ�ug�� +ݎ���+wԻ�(�)�����o�'�-#
��sH��<ğr�@F_��ݲ��ԝ�vn�i�Վp��a����;�V;42�蔵�/s3R��a����-r�ST�6.�._�-𕖱�G�m5�ǭ�T&�G�J>���"D{}�����þ�,�������^���
�ؘ��{�r	/ER�<Y�{�/�^, ��j�۫
�2'�Og<�}���_va��A�N�`\�C�Y�p�禽;Hbt:�����%�_F���_���ٚW���Xx�)�r��f�Y����Ҕdhtp/D��^��Þ��a�k�����{�"[5;e�/�Ҋ+m}�.uC`'=��hg\�g��\UX��jN��l���m�.D8�wp�Wdr�4��S�Ӯ�!<�%�0�Ws��!U�At�L&��֘�������66���H���2+)��4�wa�Ynz��(d�+ޯՄ�m�I�=<⾕�8���N�DH����5������˱B���ҝ7�V	^V��y����klv�n���75�{z��ϞK�7�<�X6tZ�D��hS=��D������e�.�K�;�G���ː�熼�w���������ٖK:
$�u\kӕ�l9�`{�%9��m	V/�Z���+��hv47bc٩��K����P�|w�G;f��4��q�-_^�Vh,��'��`�Q�e�Y�\�x�z�x'uGz+;;�jC��3^)yO�ۧ��a"�,�L�Oԙ�j��;J��Q!S5G�ǆ�r�ئV`�R����]fG0QR^JK���GF},C�]�|���y{��O�꾅G��'Z���ݨ׏Exۇ�m"��Y��U).N$��,�џ8���UL����ֻ�{�ܛk�{֍���
�b���V¸�s�誫\+C�0U/��u�ݗ������e:���z�]𺮴l�j�ӣʥ�LpU%�Y�V�h;7��y^"9�"W���$�]����z�;�����^׺��C�83U�C��5Ð�)���u��Sns��d�2�{�٦�	�o���||���0n�hX�&x�^u��<�;'�`���z�en�4�����7��32ڙ^>�{Y��#|�����~({��Җ�^&�<{Q����G/H>̗ ޕ�]f��&�u�E)˸qt�Հơׂ���W^�:K{��䒲���9����Z|���������Gp3��b�K�=]U��Cˍk��lΕ�����>����A,J5u���\^�6:s~�"{B�Y�=j�s��0�6lݤ�x�C��0zi�l��i����u�zH��1P29s�W���6�;�w
qͬ)�ꅌaH�pV���k�����ԷK��W%��S5�Ow�%Ѭ�9�Ic�y����U'��1�.�̧���H�#����S�53U��m��w+Y��TF�y&��TϮ���mS8�m/:�|���u^�I'o9jn�o�tb�Z� �x瀨Z�2��iP"��7UΦ9�ּ̽a���Hۖ�n>��yV�0r��x	z�׿KC�_9��Fd���O&re�4Mt�;�����K�o�o:��NdPqLf��v���Ƽ�z��ej��K[x&\6e�o�|�n�w�{��zj#p_��`@nb�x4�v��C�_��]a��Jqd���9=��Ѣ<�'�j9S���DΊ������%])��WI3j�Ȧ}�Ŭ9�U ��i`B�U�<|���Nv�=t7H(n���}��<���JW���4.��)����j{��c�3{}<��i<���&�qn�A�l��K'�<�&}�U��nT����CS�z9W�魵'&_nS#�1ppz͇�)�|�;DKO��Ċ�=���9�/>���C��sU��"m��-=<{�Y�כv!Ͻ�֘��qC��뒷��vT:x��ؾ27����RY�[����z�T3:�^O	oZ=����b�=�a��>h�Xq�}��;J��Gu����y$|��%]�3h���#�vyO(��W�t�V�R՛M�p0�pܛ��zkO���Nu6"/�Jzq�d��o�4����R�#)E�L=I:��]ʜ�E�81 do�̖�ޙ�ڞ����� �z�J���.�|25鲉zH��,�����[�{��V�l��+�倹�[������N^�3�F���T&�Yj��j�M�{�htOV}x�6����#���)yTˋ�,��r��znJ��s���vX:�m��G��K���*�3Z�˨z����=��A��'���[��voG����^���^)��`{�f���}h�}3�L6���c�Q��h��<N�ĸ��ӫe�[8+��_��v��v����~��q37�FL�a�{/���y1Q�6N���4L�rG��w�֣
ӄ�8�ԃ�z[��y��3����b�z��C�}{��·��%G���sǩ `Υ�S1���78���sm�%���b�˔�� Ut8��eCp�"�[~���3YS~�����uJ���%/�P%����Ι�f&�T��r��y��'�{����w�	�_L#WUC �o����|�����/�2Eh\�Z8�r#,į���[�E��d��͜����M�'��n�T�Iʺf��#[/��f>�L��Z�z��|Rv@˷��}87�ϒ�޽�;+z�[Ƀ��k}7S�t��F�{���L�0���gZMr gfs�԰��d�[��t٥ӊ�o����֏+����K��-:'�{D��K�!A�6"�}�B��j^�~�:�]�&xI��� �^(�>���`�^y%Y�b�
��oj�tD�l�Ī�= ��-pN{��R1ib�n+>G�׿gRc�]�~ѩ^�<������Y:eon=WO(f5֧o���>i���l�p�<��;�T9��]3�ͻ�o���P��k��,=���v�� �m���qU���Փ���i�[G��F��si:8���F���c<���-ܙ���JO�o�^��{�
�ؘ���:�D��\#�E��׋�[�*�k�<��p��wS�TM2���>���3Ѩ��d�z�����ԬZ�C����Ϻ��Q��{��\�[� D���s������@[S�S�x����TZ;j�dhtp/E�eu��=va���-��G��>�R�]X�^��eRiE�6ф9�|��42q��K�]�&i�Ϻ�׬��L�Em_�<^�c���Uq���Q���e[C"��%c떰��X ������f�{7���Fk����ةP�|exlЭ��e�z��ƪ>"I���=+`=�Գ&�#�����C:dkrFj�i}Wh�ّ	:��ޔ�iw۴��\���r���[.r�Sr�
�-��59n[ӽ����?mLj�S�R�{�D7���t��|���r�gE�>�*�B�谍qr��3��/A�� ��ͽ��J���X�x�?lI���;<���!(�.%@��U@Uu��S3Gy:�uyo����tXc�qE�Ƅ�l��\Qq�>�3�L���8C��E���p5��۔�����v�>� l��I����ЎP���w���Z�5���;�y�Ek��U���Hn߹���=6q������!%M�nS�e�g��T�����8*τ�!�&$a;K��԰�'��X����>(�e+�dW�-�P�f��܌���0UR�K�Rs1���.�]�k��
�����<���l҃�u�gҵP!��{�����<Y��X����SWug||�����Q
ʿ7�s-��vﯾ�z}��O�ʥϓ�[��eq��r����1�;�rsp��+VJ[v#[U�v�`����^��GA�#D�W�\�C(�'�b���z�n��[��谱�/�S���=�(�ޚ��x�F϶�!�f�O�+�4��Y�6���%��	%mӁSwZ�'(�p:��30�OnK(�\�(�c8Ԑ��\����:mE��SL6Booբ���!�a��}��[�I�q�G�M��6=��c"t�Ke=�f>�k4-}E��L���T\�1B�u-zc�X{7}��7���eNC���CeA�-L�ڙ^>.S��F����&�%����!Jmh�n�̷Gx�
��/�u+af�ݔ�����=��_P~؁�A�R���Q|ם��ɻ��8�-����ҝUW�(���nP�]�=���:��Qѯߧ�G���?���'���Pu^�P
�8�r��R�.�Qz�"F��Bb��ؐ����׻��[��#pgk�n!�x���n��k(V 4��x�QZ:5���罚�O��{ ���*�Z������~�t�?G�9�P�K�GP*X<C�\Ը���%�G"�פ�޻���i����*�(�ץ�^�-!�y�����g���g���Y�s�pU�B�vwV�}H��N"L3s�
����ZƻT��c^	^�A�=�ܩknZ�d��n�m��O����7F�;4�c�I�԰�v�!�-�������9�]P�u�w��w]�b��˻�q��ӎw?.��rv3�%�)�J�/nٿ�����ˤX�UQ����E�R\���Av;+�y��F�%uon�g�r�/p��ݫ��d�������	��.��N��r(��vU�`h�9��Іd(D�,��}��k!YWI줴v�K��(�W�����j�3�fU�9�Q�h\m�6'r��Ұ� ��U.��8����n���f�ޭJ���@��_e����3���[�Y�'MVVwhwh��)aCn����R�Z�ӵ0�,�&�m��,u���A���4�ּ�\bO�+���]qS� ���8��㻔�Z�Q�,';*b�Vٗ/3e��(:��nng���yM3c��n_��ý9j,�r؃�b��|S�zmm��h���۬�^\֐u��$��6&�\X���i�V���Y�3��@\ܓ�V!�c �ۨVͺ�ίif��Qм�e����nPk;Yl�9����vތ^H0���5ݪ�L�oEW��*�ji��a���"��̩�K[�B���(���ntUb�f��ݳ��+7������e-�8��"�Ʒa'�^	7.>7��@S(�g�9魡ShU�\5k9Nk(X�p�kv��`��e���x�^9%���M�g/��X�k$����]��,���+Wo�J&�^�`��'����;/Oʰ���B���G�����Ꭶm�r����S����\s����l|�!c�Ź�Tm
��|�fU���c)M\s�,���yj�c�����%t\��Ox��T���t��k����o8\`�5�8#�����m�ˮ8���2��I�"ƪn37���Of�.�Gq�'�\��A��pP�:8��Kz9��g݉��3g"u�Pn[��!,�V.�w��1F�s�`xzt�GKy���Ch�Z� �ev�M.ՋY+]bf�`*Vp���,��Ѹ'�;f�7cܛk#�d�%re�*����݂�c���h��;l+[yP&
j�A�j�qO��3�A�PvP�|IMYz �V�;oU�F��=N�k�)>X�t*@`�g�6Ԛ-Xh�i�n�s ��ۨl�
]�oa��mvMĠr��:��n�S�ǲ�T2b������z�s�3�ݠ�Ț5s��ըJ�52.u[ע�@��\|��(���n>`����Ɔ�Q�4y	��Kfe�꾁9�)T�鳳5Pܧ�v�����߇t&ܝ�B�_�G�>T���h��h�x���Yn��X�fd��	�[[H��^�.�iȏ`'S�[�H���p'z]ES	��0�ז��C�o�(�;�_�Id<��7�¯6wwl�&�I���}��וh�����9z��4����N[!JS$h�u��m^�K��z�����s�
*H�@�.�E�o^<D;P�fP��s�G\�C����n�J�3C]ҋN�OL��9{p�kl6�8l�+�i.с�x�/�)����w����E�^��ݧ!'��3'`į���>���i�2l������20��2�*"�
s32������*���2��*310����+2��,�,ʋ&�2���3#� Ȫ((��ʰ�"�ʲ��� ���1��*� �# Ƭ�����0��r3&�22�,&`�"�3,0��"����3�33'�
�0)31*�#%�3���� *�3�0�1̠��)��2���1�ɳ" �b�2��3(�3&h�����2��**�,�k0�"0�22��&+",�*�2&���f�*�r*�"�3(���̲2L����̳*b"(�̬����*�(����*�0�Ȱ�(�2rb&�(�3	�������ʲ*��,�##"�̈0�����2��`��
k,����	��A�H�ƛ>�^x=j�gy��k�Iͥ�;�sXͭ����� �8��\[�[d�[�9\
�	�T�^q��`�v(���}C�7�m~�^�ۢF�6���ۤ�,
b�J㛃�л�̦U;�|��-Mɼ��^�=�{���J���>pS$�����3��Py���3����UۣKxw{ݫ�8#0�8RO+P��鞵k�k�=�ѳ1=J�O2��8a:�c�W�Ͻ�v�Y�H^��g�7��ͻ綺�=�����y�c&���t��˙%��˙y��%&�d��#ܸ@!�1�ݙ-����B��9�"�:.�.�`uJ���~�O=}C�^}79�ǝq}�k�~�ٲ��V=\�U9���>�z< �-��VlQfI=���T~�7�P�/�ڿ��a�|�"������g��砸�7��6�Q;�a��h��=�w�6�,��#��&Rmqߣ5�O({����i��u�B��͠�T�����wڞ��@�:ꧦ���'e��a�]�t���=U�������^��YPx��n�b�Hc1K���Pc̨�k����u����Ǎ˭�
g��"��ެ��c2��MW������Lde�{�~�w!4xֽ�ih���w�*��z鎑�����
Y�ښS\+��<��f:a��ӡպhL���7S��KC���Y,���޸��v���&�⩓"��;�rR	��#k�;э�}s`E%I��Q�w�Ej�Ý&��3�q���ޖ�4��������w�X&T"�z�L�|����~�̵�n�j�L5�ԁ�ΔI&c���s�>v�~�C������^"�/��ķ��]S�}��\ʘ(6����躤-�-]��ځ-e��X6.�@�{=���$��T�V({����
��(F�'��$(k5�&��jP�����Œ<m��ػuP� �E�^��2ī0����D��yC�����؈p��.ǹ��%�N�c�~�S�Л���7|Fgt�T���*����p[ڬ:�#e���^g�M>%'�+���g=ո��{%����CvPĳ����pagS��\/z��v������<d��6l�3�uY�j��Y�����p���P��j������N�>�2���{��������n�����}������J?Ki�w�0be�Iѿ^�(���^��ϥq�#�$��X��=ۢ�zX�T}=͍�(:�{�+@g���n]kw��z������t�����o�0�ʗV��Z�b�펥l�V�A�_y�В��䠾��W�����|x]�[���!-�;R�{QXV5��.i��ӧ�a����r&�M:0҃���]9W¢�wzҽ�Ga��֕��6�^<��o�Ż�����{M��a�M�`Z��-�Ù��/���h�އ��6p=5讖�	o���U�J��t�)^���a�)�����uZY��:�.X��M���^\^}x��}9��UՑ�6�7�ώq�.ک���!b�.�eRn�JɹF�T7�s���Ɔv�ݯ�.G�JF9�#y�\��ݦx�Vk�҈��D�����&�`t=*mx	�R��)����	���:�zk)Wo�654�h�Qc��+�f!�"��~����刚Ѫ��|���2t8�{r������y�k-].%Oy_j�:K������g�� �U��9R%�wY`����jg�t�����y<C����-f�^��iB�k-;����z�����UqɱS��G�)/���WJ�u�b�p	�K+�"�]��댒Ϝ�/V=�����Fw���Yu��EIy(?}^GFK����
��;��Y�Y����2�ñ^��������r2�;�
JE[�r�=8�{S�գ+4��3\91d��@���L��ZaԝlX6^t��	+�*:�-^gQ�dj,�G����ݙ'J����1n'�K���
:��U�ju�C����8]Ӧ���R�uY۳�uk�6�,�5w���+6��z�bpf@�N� ���ȝ)�P���^������(��@���A���o� ��Y���;sF���4�J��S���J��0@�?e��Y�֍�M@^g�K(p����<2�ay��c����Gg�̾0����,�Z�K�Bs��t���;܄ܺ�~��y�x�\׺x�S���j��h5O�oZ?����NR>8ǔs�E��5��2�-ZV2��bJD�7����sw[^�[A��8��(�����g
~�����G�Fԫ6l�V���vGڤ]���v`~6��.�S�vΥ�pP�(0s��QX~���{�����nw��@����'�5�٥8�[��Z*�a�:�E�'�-���[��;��؏�jQX�K����93w��ϒ��޷��(k�:]��b��H����h�.�Ql?zD��U����ɓ�1���</�t�x����C��`N5ܧ�Qu.I����,
U��JqxM�Ó���9�6.��{���>�{R�p��ʊ~�t� �x��	�GSJ�x�����/%��P��l�s=嶘]�]u�!�Fgd!�R�z�VmЋ Wz�0�f����,!}j�e��x�)˃�i+qT��p5��3�Ȑ7�7����{�r�m>�
ƫ��j�<;6����c��x�Z�9u�В�]�u�n-$l�!
��=��n7������S.��WK��V4�7���OVx	��L�a���[Rl���N�D[�(��L �2/�P�xnq�v���2zXׂW�Px��]=�ฎ��x�5�]��	�+Jt�`�},�5ғK�U2:���nC|_��]fWzVE��D��Lث��M�=�g:>X,�')aC�K��t�^+�\Ex
�kW�E3�-Y4E�h����4�-��������W7e_O *�>�_�����<mYt��^^�K�Ǹ���� Pe�~�Rw6��S�/+tTi�a4�3��+��w�ٵ��8TT�����,w%��y��\��wF�h,������ܩ��+]@Qױ�7񘞥҉3��Y�2߉x|U�sY���0���c�8�J{ۘ���<�Jϝ@|P{�ϲo���l޾�y�ʣ�#�&[۶Qf���KWX��V�:��.T>y�pX�]X���}���C�B�Q��{a�U7W�N�#����]�@�� �o>��T�MhƉ�5%WI}��k��&
�\�ic�T���n#�M�f��R/wJ&����aH$(w4�����;�>����(�L����쬵J�kIݧ.ѝ��q�hݜ�N��N��Ƹ�6��Q�%p��H�E���˕'���Z�ٳ��M��W�\��J�����>�z���{|��'�/��R��!5Գ�X��+�L���Q�Z���H1�fit�0d5�+j�:��6��޺ɗe⮠��A�ԛ���#�yX�~�r܍��O�ж|��:���3g*2e�Oz�j���e��"Tx��v�nv,�^���=5����":�v;ܞ4���ܝh���xؗ[�N�f����`��Խ�����ݤt��h�6�D0�A/�u �ޖ�c�֞�=2s�*ɚ��c��8��wh�쏚�9@����n��7�;�T��1�����nÛo�(u��#�M��z�!̏v��I�ǰ����	�`�9���{.e`��j��t]R�p��C�v�ny$��E�bߡ��{k�蒆��mC�Y�X�b]��u�g�L�B��*���U -��Y�|��W��7���7�yЇӬ���j���/��4M�=F�|��'���mw;�U�R�z֧+R��oV��vzSu�-؅T�$�8b�
����O�v�����{��YLk#��Idmp�����;�!fjԽd�Y���(
ˡ۷�Lwʥ#n��6�����.}���i2u7��sӗN��mp�8��ңu���ٖ��H�Y�
��W92#�-��t��w����K�9H�1,�k���Ռ{ٜ�fN��!�x��d���..yJ}Z�1�ڬ��̀�0��xV��إ��Ί.�o	ӫo��p�/��B��W���۸f�{m@r:��f<裒̣6/�=��[�������>���kVz�#�Nq�ܘo�=��si:>^�1H�U��������ӫ=>��#,���y��+y\�k��e#��<*�6�GI�޵6l��[���f�`���J�S2�H��hg�Q�������G��ԡ�0��l��x�zr��ExL�6��]�(i�];��V���S�x��yx�������q	<Gp����f�:����ɢ������f%���QM�0��Ψo�繡�D?un��n?=��V-���;�zM%R�hG�0t{�$���+�9rM���zT���Z�d��9�}<t����ʀ�r�>�Pd(��@4�h�Q.S�Lō"��?:�sNZ�d[$�z���\�e}����	��Ѕ��"W��@��(��â��Ե�y�Sv�/+=���;sW��*��p��!ǁp���M򻽊��\&�:4W.��CƄ���Ɔ�:��E. ��o��Gאkv��1!�zuY�^��';�R�b���]�7/�&N�uN�4 *mr]{ұY�#�����o$:h�@�h�s���x �3}t�óN��3�q�:{���=<�V��`;WAK�Y��*��'��qJ��ɠ��T3�=�l��b9�>�w���Z�(}�ܿC�3ĳ�{;ʒ���7w}M��p�'ýK
�ԜS�Br��*J��.�s$���I�y�h��������ͥ�=��C�4ǏA1#�>���T8V��G�y�O�Y�`��f+�	.T!	�t"��{�Ϻ�y�m�`ṋ$D�S���S>�$a�YG>�j����K�n�Μ��׌�g0�M���6�^��������t&f�/?�*�.^ Uaמ�rs��\�ui�cՎ��q��&�T$��]�Aҷ�_P���.�,�j�ץ�k��@�$��xΥ��ۮ����{��_�������C1o�֞��Q�^�o�C-��^�=�[�tk��OU�����B,v�9�P�P`Z�����\��q��]-��+������s�t}~	��c=)/%�=J�V٠��ݔ����.��,c^ie�ۇZb�tʛ��RE����I�Z���S�Y�y��!=��+%f��n2����V��1�H^�W$�5R�U
{yzF9.MRt�ͺ����J��\S��w�p����;��U�n�V�Tl��M�k��;�/�:�A�j�Cݴ��Zi���2�_^z���%����f�P�>�ғ9owez��v�{]�FP�Y�)�j�3��e�aܛ�ۑ�q<ޣO<5�{ m��]rG8���{HǓ���o/8�r�f�x*#M�&	;b�*�0�e��T��l'%��rhw��x��K����E?^�G����xKR�e��T�zg�zlm�y�Y}T�X����C�4�ڕ���-!9��G�z)��}<��0�!㊫�t��|�Y(�h��$�g/�Xr��qA�:�TqL�-f�~2�ڬ�U�{+��S�L�e��gs��2�ٿ�
��K4�t���S#�|��܆���Z��=(�|�MRJ�}#�����1��6���s�r�:%�J�R/Ԯ"�ͤ}*�zV$�_���!�wk�Շ{���r�xI��Y#����_<n�m�O�������yb��r��s�W^|���'u���g=k�s�7�59d�&cD��2ODM����_ݞX��>�bfu�g��÷�:������D��-ar#�V���m\����Xw��t�ᛧyVIV놘�h�J��R���J��ob��ӊo�,n�qw!ґUz���+���ރ�,�c7��2��]�k#R��ىv��n���AcO����$�,�v�f����Ũy���C=��[{�<�4����{Q�=Oj��${����T�-�9��ûR�U�gU�Y�ד>�P^��|��)��zV|�​� G�f���=�k��'��j��88:�G�%�d�K���^���R�7Eg�7]�g�[��В��àM�����{��{�=�ap�y�+�U.X��[��������{znh����5�ǧ�E����$���Uy�����">�砋�wcW��z�9y<��3����# ziĮT"�������ֵE*��X�a�ͣ2�cչ:�y���PR�rǽ�:uH=7�};(�<��pS��^�н�}��1��7�2?)w���;<�::eq�Uq
�9�
$;9<uV�fn	֌>��Ǎ˭�:��^oI��ek�e��&*<W#d��u(�k�$���u �ޖ�`uZ��:u��G��c�y�ܷ���-|֪�o`�o ��%��;�
�tu^Sڧ�����W�PTA_��* ���TA_�W������
��D�(* �� ����AQ���
��Wh* � ����* ��AQ�
�+��TA_���
��W�AQ|AQ��d�Md�_	�W�~�Ae�����v@������w>�|�P)UH�AAT�� ��J��	UR��*AQ*�� �UKvUP�>�ID�) *�J�
�� R����)Q��l���D��R�J�*�(%	
�)TBJ�(*�DR�JP]�:��. w@i�P��U�
i���gs�Wq�,[��Z�Vj�4%-�e�T��"U (���j(R���I���R�[H��6M��-,���i�d-�Xh�EU6�d�*�
I]����  wL        #�    �  ��[AD�k4��v`*�F�QbF��%Q*�\ qTJ����X�4�F6aZ��VڒU�XiF�TR��01U-Z�%m�rm�5[UH *ER�  ��)U5l�9�ikL̢�m�vsX 6aDPDH�"٦
J�%
n    »jB�mU6�%i�fT��3P$�f��K
T���  f�%�f0�!)$3j�P
�C ,P�[d�T\ �J� �j̨e�P6�Ѝ,�6XS�3fԅ!P�T	���ZTY��cQ�k fl�C�Ef`C &`46�P֩�n s"��)�A�cM*ZI61B�El6������Z P���JJ����4 ��h�0�{FR�5#&&20�4ha20& �")�T�HѦ��mM�� di�yO$"��	U*h�i�� �L���CP��L&�i��4d�2A�hi$4ҥP� �L   �	��~ ?������[���?;Š
�NF
���gkT�x��/|?��K�2IC���X�@I�I"�O�@�$o���������<I$ԑB��撤DB�KE��U:�D!��2�o�fq��������a�]����[Ɲya��ҨU
uw�O�,/ě�_�?���rKEltv�9��uO���E��[��$�!��M�"����T��4��4�*i���e��Y���a�f �ܑ�x.�i
:����뎱���E4��RfTR�;b���X��&�2��̓k>�J��$�'7�isYd���d̏�CFc�K(��v��ҝ�W�����&�������*f� dʕ2��9���v,�H���{,�� 3*�@=�6���	B��8��%c.��rb�b��V�	4��^�6�F�㧨��堯k��ڎ��u0	�jL�Qj9z�������ڛ�C@��w2`�N�c#�����V��4N��#���4*t��R��X�R㠚8�^��[����[�+D����JWhL�gr�W.�#xԛðԦ৔N��N��2Y�c�)[�-V�Q�*U�ܤ�J&G)�0�6�IWG6��ܲ���m�Q�+7p��&��{v��XKN���0�,�$�|(w��n�w/Vh@9�����rvq�/?��4�eh4;f����<�SE�$.�k���RKC)��HR�C0��1TPq�!�7w-]��&���rをP��y��h;���;͌L�q=v�Ҳ6Ls�c�$�dr��D�w$��j���Y�h �t�	xgٻm�[ykT��j�JV^��.���j��z�˱Iíi���I������0���`��Z
V^Pv�Z�U��ͭ�� Em�Q����7v�W����of�R�偉��b���� �c8T��!�X����'�5r����*!�^�׻mmϒ^<�Sw�-1)�;�[�8�@d?(�c	ڼ�(P'�KݽH��Q�	�S��b�o:)�~$�a�8��sv�[�LH����AK�E��헴��z3HS1=�<&�*f��.ېw�#o�x�ڃ�YWD�/(��6�j���uhIG�i�e�̓mI�rd�X�
j������yf�1�&V�d8$��snQ/n�-;;LѠ�ŵ6���.��ֵV���kI��L�onV˵)6q�!�UHj`q��U��]�J����ͨ�\?2�b�f�KA�HRb��72�<ۙA���^�X���Vf�4��V������^�ı[#s%]ht��'C/um�K�R����,g /l�7L#):ykvԨH �xM��Xo����Ol�yU0(��D�SJ&��<Z���ٔ���e,�t²I�����)�e1��dSN�����:���V�U��^G��%!9�V��Pk�(V��-�30�/`]�m򘴚[-���R����$�ʘ"��=V�t�Oz��h�5{�mE ��V[�vT�Wivw�����1oV_ �ո�TQU���@u�����BG(��n����!�[p�5wqJ������w���G�,�&�L�N�:d�Jި��33($��[��-��Xv��fYw`-[�loD�ɔ!�x������ۧ�I��X��R]��I�hRq��X�����Pӕ3ktT�_,�ƭ�zpA�,$�V�EMk@�:�M2ZD^�C.X���Mjd	�ڢ���X��Υ�S�.�Iܬ�Y6=����n]3�ȅhn*ѕ,�v� W�����?,��A`VdT��S(j�̼�{�p�B�%��M)Kk*�Fj��kM�Xh�'ۃE�<go*4�v�;Z/RE�aު�t7Xف��B�r��l��T"����uͱ�!L�;v����a]�:䬈����A��n9K2��څ�+m��ˤ����)������W�)քA���љ����ISbR��n͗F���7���?+nnB/b��rQ��¯���ӫ�JL-��a�2��=)k�� ��lduv�Ź)^F�Bt����ݕM�ـ�#@�2�l�kJ4����*y���E*��,��;j�4�d�q���/QI �;f�:o*�$4B��hTh]]�cqd�Z���\��z��9y.�*g��){x�5$i�D,X��+���_�8!���i�FM"���I4aj���,_j*�����K�BٱzS,Y���u(U�q�˨��u-��P��Ml�c:�K"���z�k6Ӏ�i�E��x�Y���Lə�]�2@���e�)�5��l:�uu�bVZ@�Hnd�i�L�,��*�[岥�ԕ`7�޸���Q,@̤�nR(`�Y�id,��/kA!ꭡ�<�
j�6��ͻyF�V��[�n,�B��ۏn�Kah��²��5�*�ah��-�b��Ê���N���z1�JȻ�1��i�:nB(�JMXLn8&m��P�	�R`�(f�R�)�"n 2��cCnfko�cmz���1��Kp4�T�AlF�T�Q����xM�K�/6i��¤ƅ(%J��������*�f�^�iCh<+.$���wv�MLYv�2�Г�D�R2��O7����$6�š���]1������i�Bl�3܏,�4��VZ�L@��tS�	M�ߎQ�6���Mk��Ĩ$��n��a���+�QYb�oo72fÍ����y76�7�˭:����C�	�H�P*�֮�B��֔�$b�*kcJkܕ���Ƞ(�N�84��v��r�B���mgn�E�$��jܔ	oiP�-fGm�`ۚŬ�)SLc�rΡ��t��7B��Ӂ����s6�C�f氫
Q��ㅵE	-S�tq�.�J�HZ컰70	P�2Q�c5$�V۹�`L;&�:�m��a�	'wm��b�RP'hBՍ�fK�Ib˷J���/in㔭�ar��6ۼ��܏oH��7��ZIF�֔��ݔ�P��̒[sz�j��M���7[KV���^ѫ��������-hGX�����_U��K[d�ԉZ읅�[�r��3b�&9�%�Qum=jڲE�u��?&��B�p&ɬ8ma��M7n�Y�'�ᄲ.������٫os���1�M��6X�s,ش��n���7�P��@:�z��һ4�l��uԼB��s~����E��� �ka�y� sl�C��/ul=��B*U0�ys1�T��涮jJhYjU�ɨWMl������%�yo�Zˡm�˫���b�,:SHz�U���QD�%�ۖ���BAaD%�f�RËt�Aek�h%&�-��CA.�]�,`�i�јi������KTlXm@����h˽�TͫOL`����ܳ�PU�-U�-ު��J?C��0]j�f�b:�Ҁ̔�)
��dI��[����(�,�&����(�([��*S㌩��+#���-���.]���k�Z�\���l�J�@�h�,IYJ�`��V�lڡ-�z)ӎ��X�
T�+@z���F�(�}w�8ԭxV���@�d )zغ�����1h\��	�w�V]\6�66���+6�h��(A��?"�4�܇Ii�4�^d�j,���B[wy4�J�Û-�ɮ��N��	d�v�ژ�I[�6�j���i��n��V�]A�hm�1�~?Hp騈u5���kn��:����v�0�R��{��Ր �ۄ<[m^�f�ހ��n�s�d��i��;�+�n8fK��z��%�֩��{F��Oݗ�aI8�n1�TFj&��2���j-oriXiU*T7'�3[��bΊxq�v��O��|��7�3Eۡ��!g��m^R�a٭��v��b�/kd����Hc��u����LͰE�Y�4VTvV���%B�v��۫��n[�Hl�b��+4�to�#Bb�R�2��˽��t�z(1��B5��Wu�1P��љ�)��U��pk���"�mTRd�v��P��E�L�ۗKNfd��JL�d'r�L�e��)�QS�)�͢�Pȴ�KW�0U7I]e^[�8�|�]��LT�m�ѳ0MTU;"��4ѻ��j�*�[J�҆�v1S��$�
��Wb���lR���{{G^��bL��V#.�2ܬ5D�32���F�a���v��#�hu�zs�t*m-�R��"@W5
�"�o*�����f�� ��e���0U��[�[�Ұ�Ml�ռ������&�p�"�YC��%;k-ak7�]�Z�77Lw�}xg��W�I�	6�(:����q�-˼y�J-��ë`;#�����
�w�D���qb�K"�R���_話�O�so���T�e7',�Рa�4C�ub��/����w6����ٗ+FRn�;Nٮ����m.ۗ��S6�
���!55]s5uOhM��c����Î��8o.��O��'Z�u��9�bI)\鯄b�f���`@�{k��6ܶv�p��R�XQH�z9�w��lѬ\��i7I�r���ɬ
�^�q��H��:vNW
ʾ�XJn.2n�!��q�1���n�������0�T��)sJ�Wk���mER����]beԠ�sU�L$��'�fnaX8��`��Lm�} �9יK�oa;ú�
�B��Q�3�Q�]���`XՀ���N:T����|��G\(X����f�qKL�4b���`�Ȕ�c��vUۍ��9��1.@8�,oٻB] μ�z��)X��vhG�k�%]� ���dۆ�y�
��v�бJ5 ��@dҜ2	W(���HZ9�lx�.�y���vᭋ�-��e'�{h��H��S���Xa�-v˶�_|��L�qeϏuJ��,��X~7��w�\	�e�K�x0�w}��t�e��+8��N��5�N��t���WQc7�����]����^��w��mw �m�7�3�t�\��Se��	��W6=�}��}���S8V�flbod��3�0��w:�)S`k��L7�p��)V��uH�Xw����6�6���#�)�PꜟeE+5�r�mvք؝��1b�;*En;O��X���5��zy�8���[R�	9#w�ݛz!Y�X�v`#52��<��ͥJ��C�su�C���Z�*�h}�lF��m^d8Q��]���q��6�>�/��-qm�f�c���WoWqu8dy�V����}u��,]+�"u=�Nп�3������>cnuћ�P̝��-���&��t��s�;)�e���j��h�1َE
���YŴ%�N������G�\��(��Ş� E�s�HN�l����`�
�q=�HP̬]�hv��-�*�	�W�1���|���:{��ͳh��dS��9���*�s\��WC;uAf�"�G�ۧkhc��+�
�+ܺ��v#@�@�I'm~Y�3uesQ���*tN\��֮��n������i5�e���|m*M��4f_�<4~��/�c�I|���v����l.�y�����؛��ڕ�[��Zm�Biwm��/�|������+^�;޶!ӳ{U��k��}�Lg4�}
j��]r�V%���t�]�Y>xp�ݷn;}���+�����o�*��]�0T�F*,\D����s�q��@u��90�x�e�5�C�����#�����n,�6�����D�����K�V�H�oM�B�t����u�sp�y�&d���icK"����b\���&�娞�� ������ܸݘ�Le�e]�ug~�@gm��������Dfp�s�u�j���|Yu�w>��w-:�(o1BJ�̭C[u��L�|
η1���΁��L�u��8Ǵ�	tK���x���̻zGR�js�S{O������x}��|�Lv�ї�h��2�k�4�n��đ4J耲r�ۙ�@�2��`��V�=��NU�O�J'���7�gK�r�����ݮ�9�M��H�)����ur���3��L��,]��C��2���ͤ���`���6P��]����ED(5�ttWf%��0�Я\utz[�1���F��R3�k��c��W1�ݫg��v��g�wٸK��2IA�ꓭ��u�C����9���V�ܦ�[y�Y5r��O����uX��I� wU� ���o[Ѣ�U�]f���;�r鈫��v��V���Է�T�0V�j�	�tr�[����h.xUN͛5S���q[N�v�}��v6Xس��H�Os1n�}����E@�����m@3��[��2���Qވs-���}0m���4���t�����bH�0+�
{�Ѹm]�cQ�ڰ��,Pp�Uy��\G{�f�ko���p㕌��ޏ4]v��m�[�;:�𔜎�=�D�V9���B/HAn�Fo-s��-,QsB�n�u���7�gDD��ݜ���8�`���l�eJ���>��B�3��*��x�2���J��n�u
b�ZF��j�ց�.��aJ��ۖ*� ���ӗ��[']���@�+2^Ѵ�x�ZLҌ�NV�&jwq2�T�w�`�r�yZ�/���y-��'���`fN�n�d�ޛQY��AB2zqm.��ٝ����%:�gZ!ʳ�n��0]]�(���ŞĆ�W��5J]�> �p���E����d�6t��ɣB�.�#��Y��u�V�;e1�r�.��<slbF��f;䶊���D&Dޠ7���^i�>�/6T;�1b�m�:sB�콅@vgF"�Z���D�a�EQ�Z���L��X�e%�!s��u��F�N&Gl��&b���EV�ϖ[z쪛����b���r���ހ�N�k.ҷݏ.�#��T�X6S�����{8u�Ёwr��8�QcL��2�
��U�{�G٭`���]ݧ���ib	S�	��v�����I�)f]j��Q�B�,}	�i�m�O�,�������5�tm�\�F��9�ؠ��֬�)��H)]pǭE=;��f�YǗ3=��*p%m��P�WlQޙ�.�E�/6��U�a2�5],;(��&�Q�!!�C3��OtA�i��XY;���4�a,�T��ަ"-��x�E�fm�TP�1�t�ٳ���9!#�����������s]��ւ�j��0u^n�9����#̝ݘ��8|���ǌ�W*����hu�#��cTɭmn0Tڲ;T�{;VQf���@=jS�eΛ-�{������-����X�3�Ml��ifޥ���ms-�9Òk�2v�+�%"㤁�*P�{ZeT��'6Cf&�t*݃Nh��S��K�صsDuFM�&v�T�x�Qߛ�[��۵X0�ܕ�u����4���t.�)�����Uv3 ���.�7�	��e���;;�9��p5u�e'J�8X�*�����d��r�2�շ1ɭ-��rι�z���{�����I�wӬʶq�{���v2&_Z�	�7�Sr�z�Rt���> �a�-��q��S-�1(kw�n6hJqN��.�E1�bz�'w����T<��f�s[5� �l���v�}�]=���:����pPFl�@����G/�Y]��G���4ĢMp�M��D6eF�U��]��x��1�,�w2�N*���.�C����t��Z�V���wH�*YMm����)��Cf��_.v�Rf�����M��O�creC���l���>]_wm��������쥗�4�.�Wn�v><\�Qf�܎��w�b�qW�څ��Y��r���y����۩Y%m�|�r�͈�s3�r���%���Tt�GV�v�r�`5�Ry]e�*+���ށ�09+R�#S�8��M���ʙ��9�%*��r��W��'e�R���N��]#�9R��ܲZ�p�"��mm����6�W@�L`t�8�Yh�4��]s�ݲ�
�Ti�S+E�S�n�'w���ن��Y#n�%����׊����_c�-�JS4�`���{f��<o�x�c5�]1�&v����Z��k�%l��QZ:��xXMn\T�6b
�� �qH�yظ#�u�z�v�d�7�U�،�T���& ���{ogP��fՏ�<����Y��ME9;p�h���m4�t��L�W�8�O�\�*8�G$�H�]7�$�I%x��K��|�N����;��N��cC�_ׂ��O|�Y밾{��i�cpN��$}���@h�B��Q�������Q�K�p]��rJă��N���	��,�ͭ$��/����l�,@����D�lq�L
DЋy݊LQ�R� 7>��X`]��j%���"e&�Y�kc7~�ݴ�)�t�h�2�aѽw�˧cY�6��{�|�/)U�W9d���Zpb����B��t�A�%q�~��-$P�J��M��ٱ�v�K��o�I!V�M0�x�I!ygrC�L��!~'_��� >�'��n�<�L�C���ƵrͽN�^���o�J����ty�t�yK���D�xxۖ��H��;.�6ݺ�}Pv^�Kfы�,�V�<	[2����,�M8��X�@�*VF��W���Ԃ���Wpv�⹞yr��Q^I�+�Ozګl��j����+^f1�ތ��&'ڭ$8H0��3��͖rl�[���[�t$:�m5�^�����(�j�$F��e�PV^��Y�ȕY"[c��T��f���t��@i��һ1�ڎ%��-��H\}����KlΙB������t�}�,�${v��Eg��m2�N݄�LKJ�ݑU�`�Lv��h�Z��gr�	ĆK��0�Ń,5�Nwū)	B�Έ�3�p��q��m;s�2�\Y�lgXZ�e��Z�SO�mN��v���	7cUb��Y��Г)ɕ{KrȤk��1pp	�s�fg=�`2ͧ��Yf��&-JՍƇ�,�m�w!����cU��V�i�L�4]c�"�4��W�c�#	���x�J۲��[X��o�m��3�&���9�N�!���k4x�זl�S�RaPMd��<�$M���}�Ds�I�Ǻ0ihb]�:͞���G��Y4��������-t�b����68��M=��lo\C��J�0n�[�ub{M��jE�}�0�Ae�y^��ēJk[ֆ�wj�����[��d����@
���u�*�Ӣ}�:��.�Q���R��\��(�ߑ�Wz�%Ss�+/��1Tt�[,<�� ��鋾(���բ��� ��ᛶ�Ӽ�O6B�.���Z�Iۑ�jj�9>vo��ˍL��6�a�dF�}#6-�J�I�'��m�aҐ�%�I(=k�6�C-�I�eۇ���j�H���)�.Tw�MVfR�{2�D�O[�;B�g0��@J�Πk-���h�+6���k4l��].e�_ ��Yv���C�,�u�.<0�=YjS;Ul�����4�ʘ���(0՚�Z#�WN�;�-���!�`ulyJ]GY�q���z
��.��1���)��[]��cu�8؆����|p����Uos��6�O �q�!k���ྵ�;=�L�������c�MKWg!�Y���ȃB�m��u�Vb�W�ݓ���eh̬�}K"��V
\T"�
X�Q��;em<3oOL�)f���K��>6�|�z�SBwg�v%�dN���1�!��Viú]�TG)�>@�=L������N��X�dW��C[`�)�T�H��P�����v�)\)�6�%�x3;u�V��\�Qc���m�[��z�5S���yYs�"�A�o\0ؘ�������06��]!B<���8��vfn;�Y�'g�R���M�k��}2��ۄ0q�;	�n��Ln�|�]-��3���v��Nh�
-F���뗶�9�%��:�A��q'�:8q$���F[���� *�Z��r���7�A]����S�:\�C��0+4�F�e�
����*�wWc�VS�[׻Y�K.��Oh��uC&�:Ɔ��5ls/M��Ε>�xwT�]{BV'�4ډ8�9W�@Gvl���T..y������&�p�²Ԩc��lWM���Ƹ�b�h�p��/p��[��鞷̻+P̩�����-e )��v�
m�9�q[�2�� ��=Y&��i�g/�Tn��4�A%���R�+�D�KZ�v�:Sfe�e�
�u�k+�4�R��2m^l�Ѡ[�3�k&-6D�N��f�w۹u���1��J�|���)zӖx)��]u�f�擥�sw]��v�m:tu9�#�v��Oc�o:-�������/�G����=��c���p1�Q��K*�	W��;xB���n�2,p����$Н}�$��w/z���u��قH�@�^�(���;q�*�;�
��Jr3B_d�/N���]�Z�꺒a9 8���c�d�}�Ϻ��Z�v��!���Z��T�\�bY��e�����H�K�ʚ�mY����?1����E��a+���U���"���].^�b���v� Ms�p������K��zq���(��{�L��w����t�i����yd�ސ�n �hv�@�"����̇����sK����H�qJ�$B��Ur��@ݣ����WT���ݬ1b�ΗE�ͻ����!�,�v�lW-z��V��\ɒ�w�+#�.�+
�]�hw�y�|M�o���Jܽ�xf��E�e*R�h�u�R�7��jú�Ev;o�]-T-Ws��"xr\���L��[�O����z蓫\,7�+D�3	wD��q=��V��2�l�U�r�����Y��ӆ�j�������� �ܜ�kZ�{{v�8�f�:��q{�ėI�k�AGƅk��`v����u��LOz�Щ�V]=����5���7���K3B�o�NСE�S����sP��R�Е>�D	y@��Z�Q6%�����;��m�$����Cy9�/�����Z�WR�%�_���[�n�W�ML���.�<a:P%@��G�7sQ�ȭ�U�U��T��,�s����2�bދ�ɍ���I>ƨ$�[mWuWS�p�9�fc4j�=s_��t2��j1OLC��q}<��T61�X2��z�:�@鼨��os2���p���	>�;Y(.����5a����@×�_;��j�r�b]4�.8) ����.W.4ڂ�:}�� � t�����*�e�7�-9L�Y�*o��WBɜ���m�wc�0]��e��å��qr�<뻧�Ԃ�5*����a;��4vS�ssl��z��i��tS8o���q6C�έ@�Ŝ3����j���5�f��D�UjI���5�Ĕz�\��#�y\C�7����]�;�3��q� ̇�Gp�[����4�0�vb������Y����n�+x+KAX���Qm�S�l��-Uډ���m�5��]� ڗƑ���OYF�p6-�y�PVd'4�����q�',|��<n���HM�u��5w�jN���v��8���u��[|p[}���+�wH�>��٩�j�d�F��RK����qq�9rr{��e�W�$Ć�uG�iJ��e)�:�YW]u��5�Fg��ós�����Q|���wNU�j��(�7͵��5�[)Y�I�ouL,;;�Hr%����|��L)J�٪Y�I��bF!�}j��+s��+'A;�U�uH�JgwP��WעVYr&�kmla��kl��\lܫ!�,�`ͩ���i��Y�i�י֘K�Kr�g�����V������Pu��r�h�.���f��T9V�{*}J�0��ub�(�:�t�Ss�y�7M=8u�ζ�OLE�f�1��y��9���y-9Gl��9��z�+��!�[���Uf.��K.��w���%��u�A.|���t�� s���y��k�M��l��^�S�7�{�@�7;��}ۯ�'9��j9�wL.�|
�Z�=z��Ӈ���e��$��|��f�ޣ������]�ΠY�xW3X�6����&������>�w)���Ev�u��`4,��^ �n���L4���b��J��GG	;IPihf))+l<�G�\h3&qh���W���n�(yhp��NٖՎ�s�������A`�x-�����Rega
�Ԓ�#wU�#�ջ�����Jl����4U�jsL�Jh���-��f5��b�n�eI;�9��;�!�����S�����%�+��X�V�!f\�"4�;W��O���ٯ��61��9����c[x �l��C5���S�y�� /�%*�v�r��J���F�"��+/5��Y2��BlȎ�w��<���6^�7ю醓��P�!&��*!ܫo������ճHo�u�0Y���얺�5]�ø�Ƿ{��5󱯋5׳��f�%��z-�[����Z�0l|��E���
���$�e#��7��^[�4�Y�']���N�j�=�+(����x�g*�lI`�nn�8�n���3]4�O��<��5Q���ך���q�Z�Z�����I  ����7ޯx)T=����*����1�g38+�A�oH�:,YF�98�*A��:YC���wWw�]ҩX��+���im+���7oJ�BƊ�ˋ�oi�Y Φ�,�]\,"/�w)@N��>å�`���Z��m�I'm���ñ7��J|f����3k"�כ�k�\���i�^�[�G{��h� _j]�)�7mJ6����8�4*�����<�ݣcΚ��oH�1ɔ��7���aq�HU�{{���g5��TʼfҘ�Pg8]*ٝ]H�_h[��ۇ�����&ж��q�7z��0��5�@f�w��pZ8�#�:&8��:�v�E>�\��5n�jm�֎� d�lW]ы����Wj�Ժ��lJܹ|��+1$��wǏ)��Eυ-,��\{���>��
c�9�����9���5�ƺq�fN1gi{K*�+�(e���Tm["�+B�mZ-�fRf�TX���Db�
**1�m+(�kJ���(���������m�:hb6Ȱ�kea��6V�(@�
���PJ	��P+"�,U�#Q1+�ZʊH��*�
 �DAb�b�Q`"M����S�[�ʪ���K `��Vġ�euň�'p֣K�ɍ��x��A�U����+G�G�.ruj�M]?���j�^p��V�v�|���ռ�Ek�Oq�jc4��,��]ϼC��o6�YR�"b_t[��'�h���9���7�
��*n0��G45�RV��!�>މ�{�D�j�_-%=	�9�MX)3��+gz\O#��(cz��a�*��Q�i�9��g$�����3p��dKْ77�j�e6�F9DP�5yk�5���|�)â��2��۽=�+�GJz[��1ޞ�7�`�	TZ��>O&g�}������m�Ŝ Osa�Uڭu�d�N��{��}���ŧ�]�V�(�gL:͉Yg5���ZզuYN@��Q�B���p
_����=��r��1�����b:w��Ԭ�<��N��tm��j�(s�y.7�D�[i����ׯ��	��p��}�}���虽��P��Zٰ�N�v@����iF��&���,{�6!~�� �dS��G�kG7�8묚~�Må�F�1X�N���vC��2*�W�I>L���s}B�m"S.�͹���ֻCdP��ň���4�&"�M��/��<P�`��0��v"Qz8Z΀�W1�Մ�>g���"�t�FFn���N����l[K9Omr�\�rteg�F����X�$2��/��P�:���f.V4�ӣQ}5w�zu+�m]^�d;}��&� 쉸MyAUt�KZ��-��1�w;0�4*�G�tn��"m�nU<\}�k�n�#��h#�0j5��J�Ľ��4\m�����]��vR�*h��.��B�j���e�*91'��;_�P�O�z;���*����9χ�`�=��o$���6}���;(��"��a8C�h�S���1��g*g7��\�J�'��#���Ԗ�!�<���v'WuS�vmi7�8p{b0�o�:ڏ�8�.g�[ѫ*�J�TBU��s�w��D�֓}�>��%H�b�n��b�6S�['6��t:���2�k��tX'��o\}�*����C��<�VƐc��e�������uf��Q�sQ�(��^���-����/��L	�r�	9�Fv�)WF�1(��ˠ�䑃Lb3�ݜ��q)�jr�6�fq�)���[��i,#*e��X�:yN'�������(�`���#�;�����t��kB	=�;������gw;�Y��]SM7|�5rX�x���'���Ě��N$߻2����R��Mݛ�Zn��Ӛ�)�w��Ѓ;��IӈI;lƽ�0v��LXf���#8]Yy��n���|1�9ot7Bkt������x�Į�襵�N�@�� K��Wv���Iu���굳�r��u�<�g3�Z���oQ՝��$��iȀ��Lʙ��jo	Z��:�W8��5w9a�z�z0W�J����4�?�D`^*�}�:��ќ~�C�
>�����MXn�TO
�����Ko	.�ƺ�
�b��N��p�����ʻ	��o�ɛ�>jb���2c�j��te[��.��Wujۯ�
���v���O�8�2�5�.C��
��ym�,I#�з�s��4�pѡ���<i�PxQX1J��5J�ִ�u��@QN|�M��t�(.��O)�WwY7n?&L~}���꧝�ux��؜M����aO��<�K,����*T��e���U깇)g���#� (�n���(K$�z �+��H��W�^S뎮�б���i���me7�kW%M _w'�+*-ϹT][Ȟ�r<�G[i\օ�&����U��Z��8��tD�蘥t+�T܎��Ј��Pͭ�mխ�x�ydgӂz�����\�N�^KXX���.�����#^qQ\����`��n9^Q>j�y.�es�gteF��i�4Q�aUf�]/��<>�g6�g��i�E{���t���I��^?1��|�љX�4ɫG���3ޖ�
A
>*�V�ׇ͏�l�f������1{G?M�w��+������S�e-������p���/RZY�w���w�i�y0��O�i���:S�{'����Jk��RoN�c̿R��d�B�x@���@8-�FG�_$O�Ŭ>�c$uHP�Rɸ�FE��C�PTMo�G��Y��+��7H�p褶��.n��9�9��=�y:
fOMb��o��s:��9�O���&ͽ1ĨuJr��l���86���/:�I��QIo��0o-�z�>X�ߒ�;F�8��������/�"���r�3����Ïp=]9�q>�χ
=��U� P�\Q���5�>˓���n��ሷz�P�q�%8�1u�"z/gν �H���U͌���ǢM�=�:�����=�_O�@�4�̅G�Օq~rܫ1�`v��v�zW��<x��������M[��{��7�q�}wع:軐�B1��>�J��P�Y#�w}7<LrOx����o�jP��޳R��A��?[?����|��w���C�k�������w$@�XȾ�3]9*��qx1rc�C�o�Ƭ)ʰ`�CE���`���J����;��2<GQ��g���j�1�7Ps�NB�vw�� 寳���tו��ui��,:����k��@u*ި�ï�l�Q��1��2�{	<]󫭚��q���O�Lu��W�+�����_be@��e��P'��no=02\T[�F^ϯ�#«#-�
����7�Ս��'�Wt/S��B��ں�0/�V��IVd�[�EAE�N�����iM�u�`8Ȩ�LN�9,���j��կz��W��B�߬T��96���ԀRo�w���Y ��^S��ΧӲ:,+v,T��R������L��cC�PU*�w|5�Uz\�@qPw(�ɜ6s1��2���X���Aa�t~\l*&���Q��9@�I3���'��a��@�]��Y�j��F��>�%������;�"S����Nϸ�?���*6z�0kB��a�WN�2]+��/w}Zbr*�&�T���z�(.�,�m�Q#�����t�X^�f�i�f�)�]m�ᜟI��j��f���5z��,�<����O�b�%F��Ҥ	a;ns�! P�P(t�6��ڛ�8����@`9����U�{C#q����fפAS�=��<=#�����(��W
�0<5&�Sv�c5��@H�$9�Y�.��.OC́@����faE,�܌�j��&#M�gP�cy[�)P�4�nI����H�fZ��y���_gkW�䧢�C2x���V�KL�n�Ehq��\g�}y��g�h��}��P�P��n��ᡙc�D֍��[e�o�d:t6�P)P�V{uӲ��~���]���X�O'3ޖ"�:@����d������~�ɧ;�Ӝ�k���>*k�Uת?p�o>�^S��u�Nׅu��%J���i)(���aJ�u�Rk}7l��2�sQ�]���@(�o��#"�v��#�fw��|JbA��3��ξ1��������wb�:����\V{#�[��p�*@P`�w���:&�U�K�r�Kg�tb������Xl��ˆ_�^��V��+&!f�!=�<��م-Ϥ
�f 9
)pw��Pu^1N��&�����ۺpQ�p!���j}Q
R!؞�#�DS��ܸ�>�o�����Rh8kB�i���~��Ht�����%��L ���5^��侺X��K�tT�˃��bj���+R�6j��4zl@����G��?pK�W,|S�ݛy�Յq�PU�v��^N� �Y]/���T�K8j��7JL�ݑW,@�
0l��&%x���Z�~�FNt;�J���z��M��)�ې�	<�ǻz��j�Ƽ���U�����-�3�\���y�{9©h�܍��Uɝtmw<������p��1>c�Fĳi���/��b�rZ�]�I��¹u�ԧ]�lH�v���${sX�0�YW�n�ˢ�@'ݪm����ĕ��R���}ơ;c�-�d�bٳ�G'j�ȣ��Jٌs��ܨ M�^�:�wۖ��d-�����ݰ3+����g�8)%2��؇$�ًS��k5�����v�2�}�tY���0&�Ї�aE�2ݭ-��A`�f�v�[θ�4#��3��o��ݚ�X�wO�;W��: ��7\ʴ���b[b�u[E���*a�<��`]�p>ѯ�gf<�1]3�X��I5��*�t�w���,�amg�lw*�D=�{�&&*Xu��v�ܭuh!��'�T[�8LC��V+� ������d�
2͔���K��VÙ|6Z�I��-��ǿ_�o���l~��	�tش��on�դ9��Wj(.�U+� �R�!���W{�g����7�,c4�W#�EѹBb��g�z��' �_1u����+�^9ȵ��/��r�s�R��T�z��q�7.0nu��%-
a�@�^1yp�E��e(3s�fЙk��(v��P0m�������^oz���Y���5B��$Žx.�E��,f� }"&�O���dwqZI�VQ�(��+@�{�����v=���p�]-�7)�]��B��άdazN* 4斩��o�����)vY�^�>id���o1��h��b�wӀ	�4�|�9��nӭ�Y���Q>mN��G������h����aw�P�������[C�D4,��Ǭ؂Pj�ws��y۹�[�w�wy�B������Y�Iu��?�/�#U�*)X�(#U��Z�U��R/v��Z�����°�(�1
�J�+*
V�e
E�P�Q�XcbH墰�V��*
,XE�PZ�� �TQ%�U�R�"��6��!�"�s(f4(,�������#"�[+(��X�@m�[`)�� ��T��|������������y"s�c8�[�����lw���o��FMegw+2ґ(�_0��ߣ�D2pO��`�f���tk0��LuE(����û�yC��Ӱ7p+�^��G;���}��n3�vM�1��h�ȷ9��C������4L� 8p}ZhM�����r_OE���X��бc����#k�RS ���;��y�w"�� ĩ0�˃a׶��<��ޓd����X�׬�z�c�}7R()��.�aWV)�q���i���Jm�p��P�&�����VT_&tR��b��ΫQy[4�#Ǆ�W�pS���^��1�N�����K$�y��/�-V��W����W�I�8|TLI��Y�fZu�Ҹ����:()���'��A���'
���08{��+):�����E��v�G;�qwn
�\Y���hj��u����W�Qr��S8.��_T2T{�n-��T��fN�-��m�`��_[ٲv�'dޯ֯<(�4]������_hT,A�;�J��ibn�������|�S��]e{����G���F��f{���Cb:O\�d;U��/(��P��ּ���&��B��j��Oq�l\�S�b�h����StI#��'w�Z+++U+���Dx������� ͻ�z/������xia�?`�.���WV�G����^��W��pLrH��1^���T��ڰ�|�t����֠)N�1�A�7�0(\ї�����Fv�I�<c �,-$�!MW�b�T;ο\��A��dn*�0"�2�4�o204k�E�F�K�G��X���j��R�Cj����6���3����fG�S*�]Z�+7��9]�Ut�U���TŢC��
���̼o�������K(�G�����YnuXz;x>Y��'V)=m��pw��:�>�/�U:��<p��4}���X�D_�ğN6�3�"q�3�s�W4m�G���&����+�a�7������=�W#��=��'bpH1&}S�،!3��j�x�F��q���劬u�֍f{�[�u����m:6�b"�z=�h	���ΐ�	ʁ])N.�b�n\^��m�VX� S��i1�j���?���p�����u3|��1P%U(`~5iV�υ�~U�V�j��v��Z��,wr�|i
�l�#�i#��1NE0z&S[Pu#�*��B�W��Ԋ��"�I�����>e��a�;�Ƥ�$�ъ'�TR�W����./'��J�
Q��F��nz�^�,���
)���ۍ(�y���=4Nr�;���?
݉�Ç�Ó�fN�����*�c��Z���6�5V]p�|r���s����.�P��߶�o�x|m�"����p����Z`Lg]����	
P�vC�A�8����ex���cA璻�2a�pb��F�@�)b6ꂧ����W󠨎o�;�!�ş�O�t�*�qnu`����B�2�5�*�te�Y��J�{���P�aWB��{MH�
��3E22!�{�1X�ZZ��Q�r���ب��V��Ӂ@)L�X߮Ư0�s���c�x�
��.U� &w%ŧ^�B+�t(��p��*�̗�`tD��C��H���('^��R�;G��i�5wkQX2����
����*&��A��<��N�ױG6�]c��B�N�uq�,}�~*�`T+F��az*}������7�4��[}x�׫~�#=C%��y�4�L�݀Ɂ&��5kG�SE1n��8%K65>38�9�hJھ�ߌ!Wچ�ΛU~�X7Z��LJBM���Po(c�c~�b
T(xmסϺ�r&f�Ѷ߻rg�M�C[AF�]Z�x���A�b�}����Hu�yubL�F=�#T�r�pVk9�}��+Dƒ�Q��g7�Ed�H�:�:�NF��D�S�}�?;z�׌fuq9}���_�~���vL\t
���Gt����X�)5�=�
��"&�נA�#�����Ð����M�޲��Áq]*��;�E� *B� ��(
���RKV�js�7�(��1���22�9W<#a�iR7�����
��2
�S�B�ў�&
�oMǒ��&�)QJ.���ZK��u\�`M�z��@�0�vub�_�S��n�.m��;w�>�<;hK�&7U�p64ٰ�*�EjZ��$��&�����Ϫ��Vg�,r�ݼY�a�Q�W��wT�͆_ұ�*uK��I�I$�+�a����S��g���u���&��\�W
�8x��E������J6<>�5[����2�k;�{Q)���R�}-PB�M�N�ғ�AEQ�=΅	��5=�).zb�@Qâ�n�IVR�՝ᶅ�d�E��wQ�|�A[b��ӯ<�K}.���H�`�˧euK�>�1��~�m�� ����,l�5=�f�4�~�hJ��7+�f6��p3$���*�e�:�kxÐ�M�6�{���5aO*���tjX�"j^绸�/���5������ò�.��sY��f_]52�S55�yӪтĠ�k�����)G�m�8:���x�c��E-�=u^SZ��N;�3V*9YX7�M%Հ������Of�W�/~v/xi9z�S�%@_o��CȎ��%�n�2C"�I����+8O�R/>���Y�EK�5�a�����?vԺ@������g�\K�}A^сNv.3��V��ou&�&6�xH��A���*��*%U��^M��������>�DZ�X
��T��v�]I���Z�������l�h�n|��}�D�0�|�Ƕ	�Λ*�m���{JMF��R�S� ����}Jv*dA���F���/��!��Ȫ�����9@��d�M`�8��i���Ϙ��"&�.g�<�Hu[ڱR�����c�z/'�:�&o%ǥH��s��!R:��)�Rm��t�x�b���i1κ�Xs����uY�!��:(��
�&�j3�p�y��"�w_p�&����a+��@��Oyhz玷��ՆLsT=��L�_ے��R����2�MH݊z��ǲ ʮ#�����Ш)����X�j�υ�~U��]����m�s5aWn����
�l�#���G�x��������'�U-U��;�}��ٛ¶��e1�C��e�<�ؽܩ1�z�S�#>�%�py���Ժ0(;�b�X��M�m
����P��T�w��`b��}��C��7����r!�[]C��	S�b�;[HgqOy�u��Vb^|/��E
v5�+�#j ("7PnL{-ЯѠvp��A������Lu�u�>�����I�+� �] �)j��r�) \#.�#i)FxɊ�H�f�}}"b�.�*�>kx(aȠ�aA�dl\yf�Q�\R�kd�k"%e���l8�2h��'��W^�"�׳��c!Ъ�<���%��z�mYK_ 6r�Bus�຾ythk�;�b7�&ޥr���"j/3��>��"Jt �C�S0恟M�ܕ�ߪ�fP�D�c��m��ډ��T�	ݠ�`�t����U�R�c&z+fo��C�� ��0*=��8�c(��Yb��#�G�2BsQk4��B"R;��tpAZ4��u�\[���j����p=<,!U�5�4^-���*���׃�u�Z�k=��ݿdˋ�Dpˠ�k!�P`��];�Vaӈ��Yz'�Q�3��B��l[א�� �q��Tٰ�9�̋j�:�Eȡ;\�eH�T��t4>^6>�����}y�[�-�� S�8<�x:�&j�yU��>�fmllԔ��"��Z�[*���_#G�&��+��`�|�}硃
%Ւ+y�[��oVt�pc�S�����T1�)ԗ�;�����~�:l{��
Ƨ�"������hc�tN�_dw.]}�~�� Mr�*ȸ�q�฻5��*â�a�J��T����,X��L�h&��dynW�PR2�c��6���7pb����)���b>d}�u>�"���z3�?A��{zr0@JTp�3y�.<v[�������x��Es�R�\�}Պ}�s�����-����
���aW�����\~�Q|����;)'��NX���=>���(�i��g@��u��󹾙�Uoe���f��yP7�#˧:}�)�&d(nY�1�9T�"����\Z���TB�]�*����6��ʧY��M�FX1�{�-�f:c�xӅ��m*��,e<�]+,�Yˡ<�9<�-{Ք8$&��,ֹ��<M����k��n!'��Vۿ��n��������3CK%a�Z��2��H�v��O��޻��:���^c�A�c��s�m;4�����w�(�JOw��X\�C����]�v��j\ 6*U��Z��t��Ԁ2u*C����m�`.�PҦ��v�mq��'<�i�I��=9� ^�.�܊��2�*���M��	-	�ơA�u�W�p^|3�?���Pn+�\/�]bU�{:�	C����Ŵ��@0U�
�	�H	��enr.������ۉ����j��ެ����:� %ʃ+:����ڻ6;���4b���AP�:��͵���Y+��w����5� pu�5��Ik��]�e}}�}NS]j���֬��W6�}r�� ��̈]��`4Q��և�:�8�Օ,�sW\��Û[��@�|�
��n�N����֋<��sA�k����,V�/��oq./�N�oGNh�V(��X:�^��=��*�@%".V ������R.����:j]@/��z��oH�Ex���L<6WX3)��B�oS|9����7p��5�\��GM�-L�;�u����ʹy�Q57����`>�N��./����o+��WC���W�x>��'+|�A�$4����c5���f8���_W'Ff��v�җ]9���]�5�"�����n�%^oe�PF�ٜynӈ,��j�Q��÷,��}ۏ�	�)���_̣c0��S�����=�n�j�Q��V��#����=U�^r��Zb[�Vr�[9\�v�֙A��(�ʞ�ZD�P���z^L�`�6�b9�#��P}(��X��<~�m��D��:�32��ȭr-`59��4�]G��ws�I����rv^��&���V�8{*�Gr)g������@��@��a�e�V�EcEU�Q���d���Z� 1 (,D��"�b1b0�
(����
����X
EEV,bedc"���VH��k`����V[EdlLJ�X��E�J��T�12�b�X�`�aUq���Ȉ�
�DBЫ��
�(1�F"UJ�j*!ZŊ���(�T�b �X*�PU��-,"(�R(�D��Oxj��῍�}3˞M�����q,�rX�z'�zL]уp�_LB�m�T;��< ����W�#��똌�ܥ���a_���@����� �2+�U��=��qR⸧F���J("wǑ��t:,�*NB���[���Y*���P����f`L9�l\�W���)��P��ý�*TWN��#:Nϯ�"DX%�-L�ك�Q���>�@����Ă���Ϭ��mH)<��H
)�:݆�'̩����������tnɌ񒸆��}��|��}���A@Qd�*A��0ڡY�%H,�>� (�5:��l*Atu`f�=a�u˶H(q�3�%@_��i+�O�|5�������7�1�2u��,+VN{c��ϙ=���Yղ,5��/��a�:�4�R�T�'H
,�Փ8ʓ�*A��S�:�^����|�{��'l1 �v!�u��XV8��bA`x�E��O�+��i�1E��좐R�at�gG���R
N����<��믾��٤�8��*A`x��P�
Ahz�0�,1 �qXz��AM�LH(g��l��m:՚H)���T��:�f�ֻ���}������T���;@��s�i��W�N�;�c<d��ѫuE ��
��*i}�+U
�݁���1E'�<aXa���fn4�R9����7����4�ͅ�G��S'x��T˴8�q�����µ�k�V�^����܎�H�u����Z�t�c�p&��������w�����l8����a�����L���uj����e ��Ng0�m�aX}���Xp��U �!X��ݓ<�+_s딢r����<Ă����� (�`c'PѺLH6ɚ�E�N0��I���v�E�0��6�'����Xm��a��Y��E���u�����Hv�
Ѵ��!^��5H,���IӉ=J�A`}��L
A��'ɦ}a�x��qYX�(�5��������ν�o6��*AM _,��|}a��l��%@S���gvLN�.�1�0�
���s�:H,�w̓tyd�O�R}����3��uמ��~���{t�R
���@QC��La� �a��6¤���d�>eE�WI7�4�Y�'_k�!Xv³^����ι߿n�L� �l����}�1 �8���!P뗌�:H):�cSR&�S�
�wC̱bϓ�Ɍ�8�f�d�'[��ם{��s�Qa�>��I���Ϩ�V��Ă�|=ɶM (�'G�M$�}C����0�e �0+=I�!������u�^�����y���"��`|Z���{a��
�Y���a4����*$�ZAݟ2bo�6�I���c6�P7h�� �����g��^g�o|�>�{�}o�u��a�
�QLH,����i���)�X��*-#�!Xz���A`h��zϐ���1��V��,=N���0�����7�5���xIY�J��TP�J��a����&���!Xx½j��T�����H
�L9C/�R��u�Y�t�P�%f0�c"}�^�ɱ{Xޯ��(Veaٌ:�j�~�p���H�˰i��ڬ]c�%p��v��G�sk�,}VJ�\�)j�L�n]ero���[ꃰ�}@Պm4���y������;H,�'��� ���ŜM��*O����,Ă°�)P*Ag|�g�P+:�CI��_SL���]}�4�Y�wo<�ߺ�{�}&j�{��t4æe��.$z�n>0*ACL>q��d���7��� ���RbAa����+&��H>��&HNl�_r�u׿oz�4�<Hx���$�@��i&�q���;d�3��z�OXl�i'��!�nϷ�������o'Y�1!�fXv¦��bAՆ��0�
��T>IY�K��!�x��'YdR8��:��6����ZAg+T:�e��>}~�]}����� ������aY�Ă��@�V&!�J�Y:��4�R�9%b�'�1;@�8�f�O�i ��{�S�
�q�~�{��������Q@��8���2T��5�R��H;�ީ4°�)5��YRf�Β
AO�8���}Re�q1�9N������o��'�!��'���,��� ��xyN�|¤V�Y�J�2T�IP�4��w^��0���I�t�Y���o��w߿u���	�N�>��H,�M�H6����z�i ���1�3�c'C*Aa��a ��yE��m�a��(z����4�P�%yz�3��~��s���1 ��Y;�0�a���$=���gL������P�v�H9d���Y��CR1��^P1 ��T�ɣ�o��}��{���_���X���
NЬ���ԝ$�!���u�1 �u��i ��G�M3�J�G�1��=jC�H9N�0����{��r�M*�a+e��F���;O#N���s�aםiغZ�}�,�G7���M�xpp�o�+*c�c�v���Wڢ2�v�k�=���W�~x������y����b�h�@QHa��5��Me:�|�ë�j�P:J�U%@S��a$���ɉvq�n�L;aP5�1 ��J�\�ֻ|�����>�I�)�H)=Chg��a�<q��LH)^�1��ܢ�5I��5�M$)
0�P�;ꁌ�8�0����l��}�޷�����
A��5�tö�d�q%g��� (�P�cX ����{�*j��I�'hVm��.�R
AO9d��A�9�{�=���}|E���c'L�����T����Xv���X�i�<M$�
�T|�iE��,1>@�* �'S�L<aR|��߿[�k^u߼��4�*9C}`VMwf$=��]���{���$z���ސY5�1��X,7i�&3��>Xi ��+6�*֝a�y�u���{��1 �ĕ��$���a�'HT�ͤ�wH
)�u���;Me#�!Xm4}f�2v���5�2W���P���yW]�z�;�����,� ����a�R��6�!��Ն"�Xk�H(%�0�a]�X�V{��P�<�=�+V��'3�B���t>���|���=Hwh}�&3l��E��AHY��jA�1z�c
�Y���
)�ْ|ʐY���풱g׳�$�K���j��_y��}�& (���'��T��(f�i��V�q�
ͲTR(�`T*J���8��!Xi��5�
AM�N�@Qa׏�^���u�>�^Ì�gIR(L��C��t�Y�Jϕ%I�TR
����
A��i��*�&$m��
�zɇ.�
AO����|4�m0��ߪTTW'qUv�׻7��J-�e�iݟ�<�]�uǜC�6��t;���j���{�i�ݠ�{�+�olT��/��K�"��W����]�ﯟ�R+
�ɤ�O�vc+%v�̧- ������a�B���Y��x"�Y�,*AI���0������s�.���y��� �ĕS��E�y����t��'3��wL+
���^�1����*�Ad����Hj_p�a�6�ηdĂ�'}i��=o��ϾϢ��(�m+'���,Ւ�g�S�H)<����,���wq��T��y`bA��m&0�+'���
�I�_X3�5�^ʽy�^�p�[��gt�a�t{c�AHyl�'� (��V�Ö�H:�k�i��XbA~-���IY�
�AC�ה4�X�/�s���3�󾷿�~�,�&0�
�����& (�t�H)u�VK吩��톞2v�ù�g������օ �5�d�2���z�T��s��u��<�~���7��
Aeg���A~���$=Ir���Oq��/��e��x��?���י���E�I��C��9	NG�:��P�~�hh�3��T<ܐf����e7�nhŅ.:��܃:v�	`�њ�S�IX�2�H�s�r';�^���!�F�0jN�������H����HEx�5j�L�L�/ث��x
Ř�#(^]��Oq�!x&�*c�*�a�g�-)�I��X�d���W�B����*�p%V�n��^�:\�֧LuŔ���ո�$ Uq����=��Z�����v]�����Y��O�?�\�#��L�;��LϚmcd<Un}t:`FÇj��Ѳ:+S�����j55Bc��*B���W����Da�_��N��g��S��MQ��77y]'.v�����|^s�1{�km�(bdF�i�O�C@�U�=<��TE��v���؞NϢ>�*�2��)!����tqw)�Y�%�2O�BF�+mX��ɰ�Ԥ	�ݷ=H�<`�/���U]L�\3��+ >��t��U�/�3V�v�&�Zc�.���}-_�E+��W+�7�̴2�����l���zA����$Ȩ����AG�_K��S)��XF�N+0�E���9,܋kiZWa�s`�]�����p� �����zr���&� 誝���#n�Lc�/�W�<<��\S��[���Q}#���>�-4$5B�թd,)�pO�ڛZ��J?]g�c5�
�C�3Y��k��FWq�m5`�N&�P�څ>�1탷4>ѓѐ$��-�}��#T
��Z�UG�4~c۪��]���w��6>���-U�,pX�����#r�:t`��}Y��qt���ci��
�;3�������O��:�(���V_$p����c�z�хc��^�R/�1�3G@Y��-rM����R�Q@Ȫk�"�O��Q�\w��y���J�B��k�f�_�}4�P�͌��ߨd��;�7��e�s�o%6������p�u���nd�~y��7Qo�XDŘ���j
��%��(6�w�z���5�g��<C	�K1B��ь�*1p47��[�N*n�5H����G3�$nf�}� ��\VTd���J�#� 8�ݮ��:'�B��y&& �0ֲgt�|]vX�:�l�"�(P�J@���V�� ��!`�<�[If��]B�ҋ���pt�2&�Q��t�y��=ju��tN��m����e�l,o�p_i�G۞�j�2VKB��zzLz"Ԇ�p�"���g<pGi�+ѳ��uh��xS5�<A�{�V��٭�Lg��|���y&>��[��ƹ�i��~ (����pSE��r�=�%��jx�S7�悝�;�M����G��O�}J����gy��`��U+�WQy��TĺwDDQ����E���B�MX���8kE���*�x�8,v�Vw���'�<ìW���x�	��3�����E�(;2��!y:����]ZT�3���N��-a�w�:�+%Λ�a*T]���i}�l��8�r��
�x{�Mq)_�BF�����ŕ,pv���7�|��T��2�mz�إ�7Tvn�PS�\� ����-���w!��ϺeG�l�>���_�r)I��B�,�R�[T+<�\Ƨ�μ=B�}���V�j��{����N���t!�FLCS~s��@�B2�t�}�A�9���7��J�*>*&x�Ǧ <4 ��`�ꆃ�;-h���&���1^�="`W�WN���N�C��ma,�;Z�3&|K�)��Ç��ފ��
=T���<?s3+xJ�%���z�aA׍~�i�,c:�R65�*g¦cT&u��l����W�Q�U��B�d��'x���d*i�(�uk ��e�R�ۍ���juv��w�z���i��T�vR�b�w�!kZ��k+[.>Yaq�:f�6R�R��Hn�vNˡ��mS��c�A����؞��y�*>R��WNA���ԫ�����ȽFwq�˵Q����Ӿ��ц��n�}3�R�yW�+�|�ﵤo��M���6�.�_�}�Vׄ����My^�j�G����It.�b���_V�����[�ɜ�Z]W���T��H��k 1s�p	����b�y�90s��t���o�n��RA�Յ�xӜ���5�E�����?@�ĜOݽ�2��箚;f����ʒ�2p�&a�^Pe�t��v�̽A���xA�&n�8Y9띅*��������_[}�K��Ը��{�e���@�U�{�F||���X�4^m�^.ed<�ċ5��&+�D���ۗ�=�t:����������G�U��j����Z�՚WZ�TC-z�ܝ{��1�G��ۡζ�����N��Tݗ.�XkN�#���K �]r�2�z��	+(,�"������Xw�L��i�:��{j�� �U�\�ֳ�2#m�����p	�{Y8q��n[�Z0��'�@%��	�i�gm+=�þ���d}K3����A��ZΙ5�ho<���KW�I��,����+2�v�|�tKA|����[��'��!�� ���F���okB9E�))�g!1-��,��:p6����P!�u�}rC�l�=��"���6(�E��gT]/V�S�;&fpȢ!3���2p�%���s�1�7/ksisNc�[i<�:���n�.`�#٥��:�)�N���R����T��RR�y��Jd|�tv�Z���Մ˪t���A��q�F�P���aq����+�[P�~�s�g�輥y��V�sz&_e�N6-�O�,�(\p�)�f�H����sɛ�xHo�t/ ����ܩ�V�Ӏ��
� ��Bܕm��틼OM�a�B����&6��Xn�gc��:�#��l59T[�+��ǯ�p�!�Av�>���kA�e�KJ����v�;!���ml�G��Ԕ���9�!��['�3�3D����w)8!����s� �p��(r�����vl��W1���gqc��v�7�Ҳ�7h���Ѧ=�nj���.�����jVD�ZXja���7PV�`�p��yme[��^���S� F�Ye�r���=�+D���պ\�Rv;�w�{�z��A�{�}���筘��	�}��2�TOC:�!��+�&1t��^wwB�I��ܝ������x`��5�{��{n�^�}���I�
��,*�IU++ ��$��*�mETVE�B�"��dZجl�cF)�AT@QTm%V ��EPUF��2PƢ�R�R# cCT
Ԃ�QE)l"��j,Y�T+UPR1�
cF,b�
�cP���
�DcYeHe̪�%a��4��QJ��J-b-j�-,*KK���V�Q�h[V
%c�2��*4���Y*E+(J�$��-�Z�T�!Z�V�m����"�em��D����������e�y��=\��Z����������!b�U"r"�m��׀��%1��Љ)ϟH�:6�����s�@Kt�ܴ��viYA @R�P�/��4S�X�P��uc}h�{��yē]w�M� >�=v�t	�pxT	{���t��j��*�X��S���hظd��"/���B	���o��`�s��E[�p�]�p�|��-P�5jC�uӻ�z�\\�S�	����g.kT+�+8߱}��z��n엜xW�菗�t�Y?�b�k�o��Eh���7qʞȭ�k)CT06+yP5��X<k-*��#¬	b���M���f����ey���
'��7j HRDl�!7��'���$�����_e{No���h|7�����?��?�����ƌpt�.��D�IA�1��L�vMp՞���|t(��F�^�� ��ՇʝǕ:㗛cy�ا8�2c��.򝽲%�\l��kܚ�S���w�Y)��L��;.B�C��\u �±�c�i)DR�Tڽ�狡��#d\��P$9�P�B�Y��r���\�<Ӎ�̀��>R'�]Q�*f��ҡC� #62TZV�18�r��sX(��+'ưQ�m�ȐҰ�4��՛�n���<Y��,�s���B=B�֭���:�\���:n9�w��v]
R���X4"'P�])H�����ј���ua֔꽱O([4��m(�6걊9��+��y�.��;��_u
�+v/�|���k(*�V�P*����n�H���Ed���Jr�W$@�
6&�@�
#���*cG����\�j,�#P�����V�T��Պ�����dP�^Kf���LR��7�kY�\~�9DL�&��t�ZRMGv�އ	�)�;��]�v�YCXd]��
�"���b��IB�"g�3O���4�x�����|�Ӷo#�ų��H
?J��J׃�ߟ�ߗ��i|�2`I���`�Ck�"\Che��Ż͒Sp�(Ph��.���*y����b�
�I�S��+FȈB ��tk����+�)H�􍎧K'$���T<:�5���Є�]F�&��G�J�x8-����]�-I^����0��r�`�2b���d��ET*���q˭F�|���2�"���Y���H+l]���7�/)�6�ӯ���\��� 刡=>���O�72ؓ��-{��	���WAjw�1K�s�LJB���Z�:���˓pz��7)*�\>j&x��a�@����F��Z����!P�!�Hꠉ�Yw������oxԗ5_]���Rp�R���<��k=���EK٪R�Y��D%j����j0'V����k9$�#nv�E{c�X��	*E)2jX���&���w���&����NI��>���L����V�� ����Ο=�������j��i�4���e#cg�¾m����.��]T���p�n��4k��0MDG)̂�6(l����7�\P�Ã�ޏC�~�eE��Ȕ�cjN.m�2�R*6��r1K���7 �ӱQjGA��l��Z��6b<z=X+��G�º�"���F>F�䓑1��S��nmN��fH��h[�S8)2���-�ӻ:C^gz��b��蝎9O��9�~y�b��sww���T���.5�����a� A�K�u^q��DD�kh����m��}=�6PȪ��*�U���o�1�A��7����N��7Kjrw�R]$��/6��@�|E�h��ŭCCh�����'?<������S�|P0�И9"`8;>Ʃ)� I�N�_k�"8�%���ʆ��cY��s�ls\�N\T"*U���Eq��]���>J\T�+�T�x]�I��=<��K�ې��]��]r��C8}w-�X�OK�S��dڊ4�*���ą��ӫ�X�t�x�W*���J�·�<ޮW=�_H" ��`P�jmO����X��Lh�<`&I����kG^/���
:�����ӁU
6�V
2��;q�Y�9�НP���cL��:���b�n+�L��:k�^>��e��/��f�t?Jo���P�*��~��Gܩ�=i�^�s}��kG���Q��~=�3[�C����W�8����IKmm\�e�.o�"=M�V u��`*�V2FC�\�[YN��:N��8�
ӕ�\ie��s31��֨�ξT��Ub�M?��{����%Ut|6F@�9{F&Čق>��r�\�ѕ�<>V�$-g�ěۣz��ӣC�V�Te+�iUp�G��y�Ӻ�Ҿ�6��H��>�]6!Ep�E���*H�ѣK��|�gc�_P��h}�J~��r=J|��dW���§�I[��B�25D�r:)�QB=q�L-�״������#;����
����#*&��E�,�Å�������/���Ach�P��$wLl��2�Ҥ����u���v�%��\��P8WP�5��
6@���CJ�4;UXB���ƹG ����G��Kꀣ�oo�âԅJGl�<���t�b��X�
����څ
)H���@t$V�CUd��C��6�|�B���X�ʢ�E��t4�%��Y����æ�"���XĨ��˘�j�0���rYSQ�NN^o~x{��O7�I�폠!�~a�T�˃���V*�ѳ�|�"5b\`+��"�"�yEگfU8�"��V�PT��m�}��W���Q\l�}�\z"Ԇ�T ����fd�M���-�������Q�2W�\���T\����eH�t6�旝�c��j��q�.�~Ջ�V����F8�䀣R��X���u�{���
 i���B�O��B�L��46�L*E<�d��
���y�`~5�	�����?�a05R�_2��� �s: T�P`T��#�~��B���旞�er���yf�C�j�/P�ď��^�g��ȶ�k�����(@*\_I�2<!ˁ���.��\~���+��1Bm	1^_��+,]����L��J���6�DoLŻ�^�n��O'$�vϺ%�ҥ��@����[����Ł���wt��{���ެ\U;��J�{.®�s�2��wWE{�#�&rR�ΚX����LFW���UˁFF9�IXp� {�тv*$(��oJ�x�H.�>���J�ȈjyϹ�9�T�'{j���יĵ��ĉS[*d8=ެ����t�81��Z�q���w������4�R���H�)w���:�P�uf���ה�K��uC`���C���GM����jېk����h�Úu=!��hО��	��٤�=�D����N���;<���� ��4:$�@�D}(}��]{R����y��օ5V] O�LS���J�fTTx���^Tk���Ј��0&�򸜌r��|�� ����x�:ӛ�����z?0}�Y� g��}���������(�fk�ƹc���pn�{�̧ǎ�V�Z���`���2�s��I���ӝ�-�~ x Xx�=>��@#j��N�4}��mxOVU��צ_n�j-�!�f�ߤ8w7ӱ5¼��"��V��.z=gT�+��ke��;.����g�lp��|���U�㉓>A,?���ׂ�ϴӜ���5�E<�QǆM��'�ϢM�6lL=�����e%iO�2�c�N\>9Ī��֗�N��GōE��B�b�����+�"�ܾ�D(e��
wz���dU]�90��6H�G3[E8�	���*�*5���-*���9t�����7����ê�د\���
w[fŉ��q�.I��XQ��$�>��D9��`y}������a�R�]>>�-�W{3����%3��3���\2*.�+�Wv_J*&/�Lsv0����[^���[co3�CO���s6�9��8"<����⦃�%�������U�w��I<��z�G�]��ˊ7X��O�tl	� �����eC2]�V��Z�R����t�ۡn�y"p��{�=Ƶ|~�R8���ʕ3�#��b�W���,�<��H'�nE乞�p�
rԛ�h��C�#����Iq{k�8z�k�*�ukT�T�8�>'�
���I{�z���j��U��
;j��֚��*)X�|k.����l��re��d
��ؽ�S��s�΂�Q]q^���@��2iNk�%ޡ�s��S��1SF~_�s
��+07�����K�Z��qY~az}*r+�#U�t�р�P�d�ֶ�B�-^6���6+���3D@�p'!WC�
;dlX��>ǚ����(5�·v�l��N�-��]C�
�S�m��7�t��68k'!���� nf׋sL!D���s���^��\����2&��e���BxdD����-V��cL��-�-)����
ʕw;TnP�YoWgt�G�Lń)��]9$6�z�}��)]�����;���JX����Psi+�u�.�(�� ��
���GE����՚��m�w,Ѡ6�X'h�	ɫ#�+�܄�PI�o?�!�=�.�8����l�J��Ⴕ��c��M��u\1)J
����:�S�� �]��4[���n����{�pR`��J�=P;=	�Æ��6��ٍ5	�e����4R�F`�Y���ٗ`�]�y!nR�(գV)��+k�O><��1�fq{�C�����3�r�w=�_q��5-m�X�������[����vG�#�u�\}��֘��e<��˼��kx�+����|B�w�ս�+�3�^g7έn������^���T�T3�`/�C��rə�'c2�^���|2�M�ڽ����3�m�箆*�/l �Pc=�60XS���]t�{3�5�����=F����p��AhhxK����ҋ����5�wç�o!A��1��� +*f��է���o��@�e!���r�B�ho&�x�ï�ۣ�y_Z̻�o�APAXu�����p�����in>}C63�9�/{:�^:�;kwS��l!���u0��-�o2��O�o�-l��H��^�zN9(�hU�V��3�r�X)��rñ0ZՍ3����M,]�L�r��;F6�vY[�jtl����ե嬺}��Ie���d�� ��ݺ���S7hU��I$s�â'4A�I)����JUgoL�'%�9ݐ�PTTJ�֦&0�E�V,m-��l��Z��Z��V��2��(���QQZԶ�m�[ij�4�lj�-e\s*�[PF��d1k-�-+U��R�E�T��)D��1jQ�me�)DjQ(і���6д,Q���֖�b�.9n&�4#T����f0ѕ*��mZԠ�"Z�Ѭ�*�3.em-iQ���J�hcUF��
�UJ����ѣh�)Dk��m"�B��PDT��)hƵ�h�K�rіƩAh��ۉb�S,��D�m�m��6V�V�U�m*X��F�aU��m-�j�j�R�R�FղڥAZT��-q����[[�Xe̙�УYm���r�e��s(�jZTeh�hѣFF�1[A�TI��@�6��2Mه/o��QQC��i�|nH�ȣ�B�+�0_iF����}����I��Uy�V��p)H)J5�E��4�?ʰ�����R�>g?����`��X(���a#g���c��ۼ��*|��9/<�H�b<X�����(G�f��Sz�*0��tLU��V����BE��7���;;�5��BT{`���\�mڋ����p@�"S��-�ɽ�Ie�]���G�W��B�ab������Q/eEe�;�[*-�e�=��Aˁ4&�kdv���*=jr�pD	�6����u���)�+��84|��Z>n-�#R���YR"���O��NF����u{l�Ĭ:1��D
R�hn=��Ul�|��n��B��}�\hu� ��9z�͵c`�K�@O�M,�zѵF.������u�*[>{mn�u�㰛�sv'l��/��j�Y�M!�{{ZP��a�(��ܭ�<�dś�T.���"ծ��My'b��H��u ����5��(9&��-}~�d]	��IE�4�Y=����)[C�l������(3Cy��y;1�	�ox���.�$l5����g�(��>���I���l+�i�9��gρ��u���	#Ô�
et�H�*b��i�7=~aMt�������>s)O@BA���pc��;��[�s�c��\�E�R,T�S)Pp����@���ch������@Ɂ����ڛ����%�"��Y�ǫ�2;g#м���x*����
���{��\�ƛ;�_z���]�y{<�xY�yN��g7��n��Ź!��:�w\����Q������gCe*6n��-3��@�Y��-��-ɣ/Ηb�qo��L���'�xY�+b�/9��2Ef7ؖ*=����ӗ+f�k�`ktΤ(�bnWn�`���q���{��\���y 1�>"�����Ǣ=�=��=�I���,�eʁ�i��}@[j���)���:�l�ùɭ�.�\�[1����\8�=$G�:W���Ċº2oK�\��=9R*˿5�{*;g����g�ZVd0y�Ԣ����|�L�V	jO�A^��jK�͠4��e�?�W��uF�[/���֤(2DX
B�^���u��d�ZrB٧8�<� ����3��\$u*��r�Q]�,�w��7q|�/����`�����B���wuj�5�?o��{�'��X+�pu��M�M�/֪sJr�`r&u#z�� �S.g������]Z��ls\�����������Z��33����<���&�;��!��JeZ�{@��믘�f�ou�a-�卡ՙ7�:<�Y���lImQ�!<8^����J���{�Z�Is��!�F���4&DFFU���Z�:�x��	Q|���xڭ`�V,:��Uҭ�3kj��j/��TZ�#�mX�B��G���b�MhX��%�n���[�r��sUG�oa��j���X;�����E, h:=�G��{=��?$�:���=�喸+,u<T
�F}�q�:���P��⹋���]���f��]]>�|��3�E�Y�hO�(�U�n��#meu�>�~Y���8������8cĉ���-�\�^ɯP�"�Fgf��t�~�b�`c�ظpF�#��6�>w-*����/{[�e��G�+���J���ޡB�6.�[�3F��U��3�^����	�C�A�:]�)�7��tڰΣo�2���r���fWs	����y����}���Yt"���s1��q8�?��}��|�x�T} �j���M��R���EA����x�e{�Z�z���P�}3�������tc��.ڷ?�NG�����i��Z3����d��L��z\��A��Ar�n���{g1��2�O+zE���;���o�R���<v�}z�^���y����o�\)
���kb����F���\N���%1 �����T��W��d	��GB��	N������Kr"kl
 ר\����#�����4޺3�޶�{a�!Fت]J&6�fIȱ��Ј�$_JS@�w_=�<S~�ѐ:Ϯ���ڋ�^���R�zVnfx����^�(��Ϫ����T�ݕM�l�!��Z4�k��F�ux}G_z���-��i�wNU�ưǻv��f�:��`�a�tc��Q),�Jˏ�o���;@��׮�m�wy>�����x.t���;��$^n�~���+�KO�rM �����d�����3�lCr����׸J��)E!�y��H14$^I���"6K�Fʊ�F�EI�o�(@�N\yr�֪���D�[��x��k/G%s�q����r;} ��"�PJ�l����;6-s|�B
��gC+f��,��4�r�m���D�p����<:@�6�i�_vI ��]K�����mf7�Vֳ�4i		��I��G�E[t_3S[/;�w+d}֚�����lRޭ=�;�|�89�Nv�ۤ�'F�ຢ^�'��t���y�4,���{��ݡ-�|�?G�6�ѷfB���0�����ա��m��"?3Q�c/
�봊��:�|���f����fd��v�Y{�xl�A��%~{�:����FHzjC��W�ʡa%����s�o	'{�`��t�9D�Y�|�X��A�
���iIP�A��񀩏�J����c�#���^O�5=�(i��f���3:(��B�n�e_s����l*OF;"�pu7�r���h��LI��qf�8��mQ�5O=ր�r�����?PY�s�N�+��ò�����sS]��:�U}�;�Z�E���b�����9�����|��Wu����~��l��]8�`]\�f�ZէM`�[��g���z�ݡX��K)!��A@yw��)��$��{��6n�������a92D�VVu��*���%�W��.��ٷ�r��>����=m~��0��"�W寭�!R)��_��wW��������,�̚�u����+۝�\����yT��4��â���ė�#��s����Ћ@���F�8�W�m�b��i�����Ғ�$`�6`Fi*#*\�d���x�//�V�Iکe�PS��Yl*gt��v�k�!��x�IQ�gnd�������q5�-7Ð"�	��ƴ���Z.���M��)U띤+���(�B�tU�|�����̵���f<��=F���1v���i�[���*:.�yg�ͫ-5�s0��)/v��7ɛc�}�$N�%���4���G �/�d�����nr�cWa_L�jW�/o)�#�w��\��\��{�:�t�&��,�Y{xDU�Mgqٔ��!�iڌ�H���J�o���<�2����a�ĵ���k��r���g���N}Pt�G�!즂����L�ϲ]5ŧ}�t3t��U��}K��^3�㑳X�-�
��I�V�~��y���5ӣo.���~�N���O���o9D�eVQv����V줬�`�̅� Y�wS��\J�Y5Y|�]��͔�:�� fԸf�[�x�\�d�/j�5�	Ădq�9�۹���^7�y�,��[��S��\(�������\�Ү�W}�+��k�-��qP}:
b��\Ѷ-�{]�'�x��I
�K��!�E=�}����
m�Jt��6X��AU��8�BJ컊Bn�j<��aˮv'4��\���Aتr�vE��<�k�j8,j&��n�^9DLTSUm���zls�Zfb��K�{x��2�̚u�1������œ\�Kt�i�x����u	0�k-��s��Х#��ܪy���JTݾ�����.�P�,���F.n���_�{&o�W:n���f׹�=rSAoy����@���i�Gn�[�Ug�zzmR����֋K�5z'�틾�ݝ���m	"@F�Wu/~��й�[���9�hi�zf�(ʢ,L<�#��ӳ��������8s�D��3�G����sxt3�l�6��=:��Ċ�;/�VC󞏃5�Xf�þ��Y�2�[��As#7��XM򷚥�[��V`/�[���{��axꍈ�/#�ٍ����(+Q���7{r
�Z��ؽ���Nm#��k�+�\�C�:�����%�$�P9�Y��-�&hr���4�ޣI,����MP��*�5�5dʡ���l!���D�{]P��۴�j���^74봝�gp���ДlYWA-� ��Vέ���gQ��`�+���4��Er8y�3b[B���lϋ?\��ІlC��X��z�T�KM�����a���Е�]�H��Y2Z�8�E��HX�YLVYI&uV��ٜ>,�=���M*n�oI�"�bb�MG�$�O�<!�]���%��t󝅕x)ָ�b�
<0�33L��쵁���\�S1b��|�,����`��ɐ:�%���N�������C�o*s�u;��i�t���!8�����0�n�9���9d�.�L���zS��т��݅�+��x�E�c@ܩr�*a7����{��n���sYN����h��p��&9qk7����ߍ��z��թ�=�x�KKo���I@T�AZNW]�PV^��-�C!�r�-�/g9,Ì��>G,wb{�+7@��[���}҆��V�T�(������zˁ�?*�{y��r������*�%�4��P]&�ܥ�>�����7Nn�T7��
!�����۫�vV�����>��2��>�94����R���GL*��L����B��m��R���+P��eJ���e�0�p��(���)m�-���e̊-nY�QUm�G1q�6+�-�DQ�V�,m(�,�!1H��8�(Qkq(��QbV�Z�"�h�lD�DQ0�m����hTFҰEQQE�.d0F҈cQD��-�Am
�1�Q�l�X�*Q
��e�j��Ler��U�P��#R�QV��Z�k�T����Z�F
 �EPV9�bŒڢ��
��D����[l-��TDX�m��b喳X�@PT�2�DE��b�ʓb+X�+�b����]���^��FJ����n�b\M��Fl`9H��LA��Ѣ�
�72���	�[�a˽�b������9 �'RH�� �]�Y�1��r/zͩ;ș>�Ҽ�u�oa%7�9�p�C��3��$	�3���-�yjޤ��4%�5Bh���	cb.X�j*{Rf(;�;u��d55��ʡa%~|�Pr��%�/��AS�'C�lJ��+(�t��]:�ogf�^�@Hpv�WL�Gl����uz+ձQ��,�3�t��yG�ĎJ�N����
��ke�Ԋ)f��w�k(v�S~=; _��%��M���Q|ŵ���t�c�^�eA�V+񡴼�==�ө��&�Ջ���"�2�*�ᛪs�Ιӵ�����0���Ƀ�Tӄ��}>91�Mui�+�N���h˼�F�����&����]Hg[i�X�0~RO)ꖛ3yt���5τ�����;lڞ�3�ˁ�v����۴ݪ	��r45X�5�]l)���%�d���G���B�7&�S��{��LA�Q��)|u�VX]���p�e��j�<�)Rt5�Ջ)ٜ};��x!���m��3�^�
�Ü�7�����^�u&��p������V9��u����<��}BrY��<X����J6,������;8l�2�IJ��n`죏J�Y�k��}�!=��t�ZwP�,��<�4r8�X��T+:w��C���rCt�7]�y���:o7T�N�}��A�u�"�C%G��5�K8�H�}[��.Ǖo`L��9��~�U�i;;�N�-�C��-EV�:C�:YQ�N-�N�6�܄�P�J�dNͼ���=�S��×����e��J��8v-��[��z�9ODڄ�9۽��]!#��������K���>8j�Ԭ?o.t�T����gT�GW�����5a�Tem��p����R:9:~�<�?k΅o�D�a*�������cp���c-��z�y��r�n�p�T�"ȭ��~1lrq��P����W�}K��3N��V;�^�w=�b݉HU�YB
�7�W��Þ��Do��yGm��6�8�[퇏 �ɚ�2ص+��uk\�F�������y"��N�qə7@�^���-���$��8[�P�)�+�J�Rl��}U_W���ͩ���ϒ#��Б�:w�:E�.Ϟ[I�k3�oRͬ)�I�ܝ�2܇Ca���x�b\p�*G�u�>Hz	=zg�`�GYKBW.4�Y�4m�BM���a�k���c��&�ԇ ��|XI=c�];s8Y:��� g����Q5�4�W��c(��(0�OL��dkU5oۥX�C�;)o����^H��/v�B��Nz��X^3s��c͝Z�)�%�^Ѧ<{qD��S��Tsvؼ�7�u�7]Fh��1�z�Ʈn����(��z$g�f�j��e�z�;3��Eʄ�4^��[��*V���V�
��]1u%󷽬-k�d7}
��N󛺒�}��W�;����M�ղ-����/X�J���UP�Zƍ�K�OF*�+��y���]��<ͼ:�R{�m�S���;-��˳�l���N�ԯ�ϔ��V���ԑ!};�WU�U#�UT6ڬ���ތѶ��F��Y�����;0���j'+�k��v�g����V��LJN^IΓ�m"G�w�^k!q�Heٲ�mBMb{�ejl��P��nF�$FNI{F���K�U�ƩFuz���CN�;������5J�v=tkn"���#�o:��p��C�۴֧��-(F��w��>���A�}N�[�����T��KK�,@uqu�u��x�7��so��A�{�v�7x��˔L�I�K*[+�!$G�H���5\5����|ڃNk^^e�ܤ6ƕ4Lo6���!����t�ˇ)[<��,�OV�� �+�M�#��jU+���+l��O�XP�+��"fA���ҫ����{x�6c���q���.�&�::��hK�ZTn*�96���_i�������t��n�p�!-֑@�:KW
�/(��f��c\ގB���婮��vt�4�h�7Hg���m�}��W7�ݣJ��}�&IG�ZI#
<�ݡQ�^�*]���k��_e`�f�h�X-���:��S�]v�b�����G��I��Z�=t�w�s�1��u����T����:f�����F8�8vs���´��LW4y4B8:�l��yQX1i�G �5x���e���Gx��B�i��!���R�s+��޳6�-�/���%�Ψ�R�Z�a���jd�kq$���F��蛵�M��{$_7�W��.�B�3��G)�Yc�8O%Y��ow=+i�ٌ���~J��7ڊ�ud��jF���l�I��=C�H�-�w�	��\�]�|v��OgY 
����޽�O-��3`{�OZu�r���!�g!��+eNv/��0�9V/U
��� ��Ed�9�k0�L���}�O9�ŧ��P�\so�hOWJ\��������Z��yf����C{��ԓ�ύ��u90��Z�Y�}J��lg�W�3
_�e\N�Q�}_�ײ��ʈs�/��[	^�F��]�O�no���C��ҩ�t���iq��'��v�M�#20�8�4�����p[�\�݃��TM�0[�i4�!L>�����9v��$U�ᝄ3V���22C�R����	+|�v�WZ۬����`��z#��#TVU���CF!n��^͐sr�%�+hb�#p�h��Ѕ��QL{�d�7�u�;K�ī��`; qv����+�#����Y;قWn�2�Պ{���q'2�U��t|ݪ�L#"&��V�R9���g��\��Gtj;�ա��ɗi��C�5��u%}��=]Dv�S�vBܭ�^n�=��[���o�)>/G��kf�[����{�R/���=�,ߖ�*��^@�zy� ��	������CW�i��I���%���`�ԘB��y��e�-ɻ�u���RkV�;��(WL]NhK��o����r8˞Y�;!R)�Ѭ���\�L<�9Rz裚��+�gƶ���M�e>�)*
�]#k^/m�J�|%^ۮ���;yG���ыZ�f2��T��ܵK��&�3���U'p����Ǜ���#��w3;���*�,��O(���	9�FF�SI{*�B"I�֝����U�r��U6���c8���������8V�� F��FS�J�L^��K1n'	3lH�n=�x�f���y{��sʸ5�{p���EGT)��4��EN̒����Iv5Z*�]�bI�TOm�R�y(^�Ҧ�zފ;�`�{��[A��˹9ݦ��t\A�>�X>ܓ��{�A�t�l3B]+�ns�՚YZ*;i��NԶ@F��1�L�-e�Ρ[CV8�F2%f����)<Z�)�Z�vM�y�(R �H��wojh-��Gөa^�:��7�����i�7��=�j��}��A���&��ѣ�jkTJL�J�p��q�x��qo-�ۊ����8/,����nۛyC��n�II�/�*�Ӑ�w�ru	]�wsV�rn�����V֞C��*�2F#�]���[�{љ�t��jڰnew�N!uv�-C+@#���+�pN&9v�Z#|t��u��ސ\���4T"�Dzt�O�ҷj�bW�gm`u���ՔhQi��r��qM@9�a�'R���>�S�fw�c	+N���иU�Ŷ�I�|*U��N�A��lQ��j�s6�8���}2�*�n��deEM��n�_d��X2A\"���;���Z�)�ם}��E`�k�ݝw�9��9�X��]I��H@�)��GH�)����U�m*K���{����V=#5f����&�
XU]N���cx;����w��6��y�hu�N��SÔ���2p���SxA�:�HN��T���n��[������21�U!�,!�]�BĮ��v��{٩"�%��Mu��t�
�]J�޻�AQ@×\���R���U�r69�Rv���*��z���ꂛ��hJ��mW�Y���ǅ�����Ѐ��s�R�1�ګO�Z��7!����L��gZ�=���ͺ�ў�C��N��T�VPC�LM�o���*q�D����m�J�_	Z��X�_ۘ���D�e6��=[L���6��J�*jC�KJ�YMKR�n�ؖnU�C_�[��4>��j�)���J���QCsU"��`�U1�8Ib��K{�{�s�)��ӆ6��M�:s��G�P��������*�c#���"���TĕKj�"(�

���PH��,DQ�
�QX�[TDH�QE[h�"�����dY����"(�ŋ#b�Qb�1BҨ�b1@�EEUF
1*AU�b�F�UX�X��(������U`���-mR(����Ub""�(��E�T��F(��(�"*�b�D*1�A� *�`����F*���DUF(1UUEDE�����)EU
$ATPB"��Ub1QDE���
�� ��*m]�[��n.��vNQ��*<�:�ENw���,*�������'E������6j��]+�3p�絕�[���·�_X��{mn��2���4��:�D�z��Wʽ����Xvy�e�6�H69�S$����g�/�����5%��ͳ)|Z`����J�7�V4��aԳS��[� �����f-S����\���V!��ҝ/���p΀X���H{���n���0��o�B�w�@ɺ�̚����01�7��U���`؅!l��%re����Se��Q�����������Y�ן�j�Cr�o(Ts�`Q�z�&s�or�Ke�"y�51�}:(��ϩ[�W�a ���`�9���MN�`c17k&�X|�Y(�yV�%G=���U�7}g�:}����[]����&}%�LѦ=�{���i{�w�1V�aI�G��՘����y���SwO9�e�XEq�]�j��� aj�x��1a�JUz�-�����W-�E4��zJ���uP�m����ڱ<� w/�5]�2�H���.Q�}�#����e}��O�qgM���]D��"���:N�:��mG�UȽ뤊�$�>��!�ݑhoƷ֩��4.i�p0��3�Z=�<�-�y��Z�st�w3r�@�D̎�R;�װ*�lj�i�'�ֳ^ ��7����M�S� ����3��u�oA�UXd�t����t	&U</�άU)64�Z�V���V ��p�:�$���I}�:��AH��S�C�ap�Ym���-\t�_8���9���:t��mi�=.��Uu� �BxG8�sc:�hy��׶w��Y��޳���T��;6�L����o5�X:�0�B�V#yWX����h�z��x�=�/ue.����f��B=>��:y���J,ps���xQ��s;.�0ALU��K(d��{=;:��K	�!>vg_u�;�*P����*<f)q�Jr��G@���_�g_r�2�9����_m.�	>��lq\ō�)�����E��oNE:�8��>��N��[��XW���q��y�M���`�ز��Zg��d�w�����ތ�5��l�˴�x��K�x�V��V�5ک���[�J�3�7�A�����`��@���G%�N��#}��)�eU��Ktw<gyU&'���"x`�[0
7Il�]��i�I2��'G��%Y5pGq�������4�?;δ��[�5�I��h���5�%\V��s6�w����}�p���ð��_LU}y|�d�[Z��[7�1s�)�h1W����8�j�f����4�ù>�YQ�swpD�G�[:���b+T���������$��l+74��W��z�)
�T�53O1�T��.�(`�̬�4�>*���Y�����Z���=�/�ud��U��n��vдմ�ʣ4�	�Z����2δ�7��]l�)�oa�N'c+A��73�h�%�z{�}���;k�2���s.-u�#}�Lg�Sx.ܼ�"zN�{�*��ax��؋2����ܸ�+��jJ'-�v]*�Y��eж��/x`���]�O��S��'�ν
��|�C����)��V��@����Lp����,?vP-�i�ۿ=�n7��ːw�3�L^����:��3��L��&Ae����(�ga6�z�e�b��r$҆vF��|����FF���HO�`���b����)��O�z{[c�e��J��'�w�d���#�-�i������&͵Ua%o�!E�4�;��m�T����^���q����on����(0�Xi��h�G ��Y"�Uc�XD�Uaeia�5���
���뵛�4.&�	)���ro.ItLH�޼-Wlo@���\W7Qͥ���x���羙�&֘ƕ�cO�M��"�Oo��O{�Mq�5����bY���^Ś�W%n��v�U��S�Đ�x:��՛a��i�[�w��IԔ��؅�!l_�ơK!�I��̱��eN�����wX
.v��-Ц�I�Ý]f(�s�#��F$z�R8<-��3����Z�&�����-=ս�v���BT�O�yJ�x�V����'�]��'�8l��~Eme=vK+-�����h5�;-%�I�}�����*��]�b^�TA�����ֹ�#���z���������_`�T�P���c_:����wm�	#9�Q6k��	#�9W6�V�F��z[z�W��r�TMe�}�S�Uͧ��"��=]::�ȉ����W��tmd�xt� q���XU��ߖ� L�h�m^Rz4զ��¨�{�*p�Uԙw�TWܥ#�]�{D�����_	�_p�W٠��A�8���&1�iݧ���b�^m|��u{P����z-\}XYOxk�Ƕ�YC�]Z��Q�`���5<4���|k�v������e�3}#����p�a��K>�.�ȱ\��W��h�ZΕ��;�2Eez�V-�W��j�gpsT�0��JJ������ǉ�X�UfnK���#��Ⱦ���Uo[z%������jWX�3���T�ӂ6���-�M:�/9΄�S��t��IB'L�Gu�ܢ���lA<}���T)vG �T�vy�CQԲhe]ŝ7םK��&����3R	#��e� ƽbVa�s��U�a,J��U�ʅ$V�u�k���Jj��̋����E�ױ3���5(�L�c�`�l��#��"T�~�C��o:���*���7��*��-M���J��}Z�T'�u���[�˚��Ҩ��SF������nv��+*Y2���嗀[k]�6�'o�����8���ƞ����C��wG���.O�%��K��갍	T��m�F_]c�[��F�޷�-MJ�i��f,��q�m&x�����{ݽ�h���P�Yv�E�m���,OW:�6Z"g���qn%3�_kL�Iz�nΕ�����YB���fx�����F�1���u8r��<����v.F,��q�Q_w,��yz�RR �(w�6A8łX�e�hd��T0����s�5�����ca[&���^�N(�λ7ɶs^j����#��X��V�ڈ�V&MM9yK�ͬiX���T��۽7Fb�8{�'EŚo�aۺs�sipv��7�]�)�NH}Jزlc��2���6R���孽���Z"��vV�70j&=E��d���I��U8b�Kmϓ5T޽.�Xk�vt��LM�y"�J��)�K��{����Z3��.c�o��}_���X�g埞�0\��M)� �]ץ�r%د�p^2�W�]��9۠7�c탱�Q�5��.4FAC���x���t�.F_aw�i2��{@:��� �O�kU&3P�`�A���]�76�e���Ft����Z+z���X�u�#��l\\�}��T޵2rHѲ�!���L�7-L>ۆX�0����k6=u�/w����E��w!��t�_6ۃ�ėo�n�*��t@��#�������-���i�q]�a7(e����b�h.�X�F��j���kIˠ*������m���s&sGn5��KV�9���|��^�{�O�Gq���T4WrU�	[Ɛ�uo1��*�v���]�@�L��@Ov���P��mMW�s8�wlSDD�cO�4vYz��y`>HV�ɗ�r���#��j���ȎԎ�@���J�sl�NԳ�:�1R�s/�]V�
M\l��G
Mf�gr��4Oc}q,t&t���ѽKy*C�^�Q]6��kUD�M�OC8�vN����=���	�s�]�9'W��k��ӌs跎B�n�r ݮ�E�8��7�h��x�[�cv��Gc�V�.�C��<����jpǀ'��*oK�uuE��h[Q�kle+�������7	�tʼ�l��,�^�����\��\�5@}�u�;�o(JH%�+p]����]�(��I+�ogfے���ֻdC0��ث�ɬ��ea��i��8V=��t�WC}��P��2s��0�/�_XW{�k���r��.�K{��a���z0�G+�:L���͔K9�>�bIG��䚆m_!�c.�R��uz���kȺ�j�l6�I���B�-|krV��AV�E�&���9�t�����0�����t�VJh��}{��o߹�S�
1PF((���*��QQ-�Q��1�bň�"�TdDDTPb��Z�EUADX�X�"*�*��jŉR����EX��*+PUb�(�b�����PX��X����1�[(*�+��TE�**�X��1E��QT` ���,�QAPEDT�b��PQAEEA�
0EPm%�U��""1��� ����U���F"�Qb*��+F1A��VC����\�jȜ��I�;s %�@�t�:���6�;��z[٪v�'k/��e�L:=;>��b�4î�`��ZYJ�1'���C�*�3}&��t�˾���/L-O*)�a�}�۵�E{v*W4�����WF�������#Z�xw����>Z;��pz8J�{��wB*eW&]ڻ�Oj'�-�R�����y�r���ɓ&���D�6RPB�ˌ�-�e�أ&OI)f�"W&�C|i�\�;�-byD�u�F�������هI�4�)�>��m�ֳ����E!/i�l�u?[Iǝ�^�w��S2��͝D>��T��{F����T���3�ˑxܫ���]��7k}��Z���w�N�8�R�ʼ���ǓjK��Bx�A�@6�M����h�㛅��J����5J7*F��[k��^�f{\́�Ob�{�v�4꼫}l��Ss�4����8P�N�N�v���7m��)ʐn�7�D��[Ҧ�苊�gC
���K�B��~�5�J����U���]�{_(ld����4�2����.��(�oI;r��F��1}P*�k`)'��7������s�4��S�Y��3��#W�y�޴��MG��Yc�ߊ�&�V>t��x���y0o�C2�6��]�l�L�=K�J�#����������i�n��~`����%�^h�]b�9uú�3l��j Z�T_]ۜ�f�%N�IG;b�������vq{X�]�lLz�۝�iܠ���0��}0��)g5L��pM�7��C���z`��L�=�!vz�q��-WZҭ<�%�B	����'$3U
������qud�ǅ��*��7$��V��lRꅋY.��4�U[-��5flX��M,;+t��i1�9�[����jPI��s/��I�~a�u�n�R���w���Js�MV�oo,{H���_T�Yx-5��	ݗ=�9t��d�,[٦�՜n��K/��TK�*r��P��5oDa��t�J�����X`�^�a=؞��OY��-��sĹ�N�9��79�t�s��z_W@L΁�Ve�I�5(�u��˔kJN1"���9�xt��N���.j ¶�d֞q�U����UVcOp���&�-C�ۧ����t����o��]��hBq;��E�<�����l��/���s�iN�'��a�T�m�vP�NB���du��b�e���ލb2t"��L�cj�7�|��+gl�1�-�`��I��\��q֕tZ-ٵ�+�&��C�pɻ[�<Z�7 �����jZ[HX7�f�0U���4ˠ�A���7��)\�a�#v�*�U�H���!�1��q���q*���&fT�\W��X�p�PDf3�][`���tV��K�2�VHt��I$��v��/��;:?T����Kܗ(��j�y�*�	+�!<שs!���cG9b�Ī�m�����V-��W<v	w:�0������4�A�^s�wyJ:9�����fNRrz�9��rþ��+V{�q��i�y�����nr��*��f��B��y��]r���3ܕ��Qn�Q6�/:�[C�X����T��YqH�[V�E�cop�����.�=�c�ֶ��-N�;�dnT��m����qDkt3*�k�t�\��cj,�^�a�IС�R,mβ���ʞ��V��0�5g����&W��1��ە�����ѩ;�K�G>#/�S\��Bx�7o��I�9kt�d�t2��<�h�����Wt\%��Ⰷ�{t�9]t����Dq�:�4%f=+��>ac��3"RvqG�k��u���x ��s��D���^��X1Ӿ^+��Z^�Rm:�5o@+��n�Ȭ��P�X���Am�N���oJwP�]ӱ�O�8��ӣ�1�d�,7̗��>�r���z�@me�o=礽�lB�0�U6��(�ԧ8o����o�߇	u�V�^�{���I�v���z��Kz5.��>��,�=�X�řbi��q���^;ʲ���1�4��Rݻ΋��vH������%7'��m�]2���Y8��BUb�%�<���޾��R��o���j�i������WR�Q��78�_S��w�'s;�K�5����㹾�E`f	�Q�{\���T�}��5E�#��F�K6�lq�>�nyQ�_��/OX�3�g����ညȅTy�6^ܯG
C&�*W]&ps�y�;|�˷yO����Iu3�圱[9�������)$ �>��eзzv��EG%����H�H�6V�d�z����x������o��YJ��B������'���u�����$��:k��o�-��{9}��f�\�ANt <8�vt���8mZ��+���nq�e��.�{g]���R��s���f��Ted,�6�r�����T�!�"�kK��C����TU�2)Զ�rC\��/ݧ�L/�M?�M�2�$���W�d`��R�ZzP`p��Wa^J��:�ώ�Nr�>wi��("��#]&z��3�U/lc���W��	��R�-OVcN>�O�gOT���B�>����fBv�	�=��^j4�.}+º����eh�V�oQ)��I�{�_����i�8��/m�Y*a\�P�H�־g1ݵ���xe�FԶM:��Q�3�u\��tj�1��=���{��H�)=�\��s0�:6 8�=}}g���]���:��No$���z�Xq|�3�:�I1�&4�>t��JwE�9�|i���np���;�>.D�N2�4�����������X	�R�uEmM�E�A\Z� �mV-�Z���B�gY���=KQ���������Z6��hj�q�p3�Dk��+T�T*C^וU���^4L��%�UcG0�F���U�/]+���uUkZ���Fp|�.衡�2X�f��]��:2��N���^�,#�q������M�Ⱦ��"�9[��]��23���e�jj�e,�V�5�d/O�s�o��c������9�i�-�h��Xp҉��zvGG˒Z�{�vt���z�U�&��r�'+�l���WgKc�ކ��9�+ Y�;��NaՍ����s�M����R#YP)�\��xU�����9Ǥo�-�V�3��*g�{KZ�R�3�����<䞨b.�#�<-����1�^��9mz�L������r���t���O�w,�H�_#�)}����'�;��R���e=�����\��F�[ٖ��=ym
�Z��k���'jd>����pZ7�ݷ�Ӆ&��;�v��j�����y[$����&$��6V�H(q����{��sa���<�B��ޟhP�xC��yFM�N��Mc��w�G��
y-��B��ۜ�$,\�f\d.��d��;�s{�r���p��ϝ�4y�Q�3Y��h�����l���Y�=�U�N�l�'_T=c�H�.���搌����m��i��,�����ݽTs@������s���M
��z�j9Ox)�vb�{O����J�W��Vw�	�"2^]R�tm,��*B��+�
�+K].�e���E��k�޽���¯�epH{'�iբ���#8����Jو��I2�������:���R�H�r��.#��\��B!��At(Z#� J�*P����|�R��9W7*���ü����L1'%c��3_l�,B��b:���ΜҰ	:��2�4�N��±���Y�4R���Gnb	�֦�4a�[��<Ppu�Ci�o,p��V	��Z�݅�������;o#�d��z�;��X��R�;�*8b���K���'ciNɄ�BoN�V�t��ɫvB[:Wi�آ����aљ;^��e2���Ja���a��v��Q[ɞ����&�_(yT�yۨ懘�Qr\KT�f�Մo}��:tD�Iv��7�`@�^n��&���э�]L�4���ˤ�с���f�1ە����b�Wep�*R�,d���
�˽8he��]c���oa�t����+��S
wn�3X�5�{���e�.W��.��!~��o���v�}�tl,Cj�6ɘ��UI��Ky�Z.<���G����)�fp��22��(D:::F9W�4�Y-��a,��u{g��BHNe�� ���>Kf��P�	T�wf=��TC�F�ee:��c�|yu�8��,!�$N�(�F�.�J.',���M�
J޼޼���}��ޔPPEAAUUUX�TEJ�*ED����1PPU`�X��,��UQPV""[*�,Nڂ�-�iF1�(�*�#F�5*�e+���� ��R��%����ET��B�(�Z�b�%�X(��*LqU�V��5�DE��-����X����ھ5��m�Wr��IÕң�[��u�N�^�Ƹ�\��_7�~e-�jl��H���8M,����.&��R��"xq�J�Ȭ��{}�h�zI�'6���{P���m�7��0�ى������dᴶ�a7hv<\y��y�.k`a��S����j�jw�����܍HI�K�S���p7�MN<�ͺ����ܚ�{Cg 흵AĶ�Ь	��웯D�O�����c�m>���o�m�&Ў�ba^�˹'u �FBɚ]W���g��iw�y2�_5���}^��Y��q3!}�o��`�:�v��ļp/����F��Vť�~ON�zh4��#h�ņ�8U�P�s�Y�˛L�WpE�Wo��)Ն�S,�7���]��>���rc�z\��	�|f�;��=��2�i	/lR���Ұ�48�28e�2uom�no5Z\d����t%&�'��U�_�\�投�~}O�1�m.��C*����p��!! Λ�p��o���^u=:n�?D�mt'�J�b*��J��n�x�jI��U����;����:ӯ>3��{��y<�-�k��lbЭb�1^'w�����K�j͞�,�tX��GpJv���~���؝[|�r����"���Z��+1uSSK���	�_ ��9���W�Q�%�v�%"���
���L������9�	���^T���q΋77j��'R�����pn.Y�@k���f�>���9��Y��A�w`�=c������8��P��]I�9s>e�u���3}������c8��[�N�#q/����e>*�v���ggc6�F�����#�/�k^�'z�W3��Xن6�D��+i�95��d�'$Q�4jo�2�7q$���E'��N��}R�̈=A�C�ҝK���۰LG;XʚYCFȁҌ�|-�*V�NIۋx�or!N��tƇ� �ԧ8�F��F�X1��A��ޝ�\\�y�"y�mK��߰�s�l�&�:͸��buո�{'�on��6]=�T��DGi�s�p�ztJ�A�|�&2u3�.\ܡ��6�\���q�dC�υJ�+�]��G_��F�N�W�.��^ia<~�G�d��t��k�$Ԇ5�?vyk���e�s�'h�2����K)�����T�Fb�G�:�����#�h<}�lF$�^Y|���3"�j�{6�zrվ��*R�D�@c�)�U&ڎ}��s������8H��b�S��X=��Λ�w�Cޣ;q��W=��.��E�}�:2���m�ޢE�80�}�˝��`��:aoH�[]����[\�5��Cs�p1/�2�r_7�ۺ�gt\/�S���ɉc�ޕ�q��xt�\�K��z��/�oo_'��U�8unQ̞�T@�����&��Ɖ�&jN�T.n��b�+�^ٷy�ɑ݃�.��#U	̝���[-�k,Z$�l|#�[� ܰ�B_5[��*�k:���d �;���1k$�Mƒ癋�CɵcC�Z�z%R��zq�+u��m[�[�F�Ì[��f�q��-c�T��fu�WT��d��m�j�E��������f�p�Z-�C<sC����$[Y��ڶ��X.wn'!o7v���O=\�V��z����K��y�y�|�]ڳJ�I~�Ԅ��=��=x�1B*^?(�Jƫ�ʎ^G��i(�f�+��!%�` ��P.e�S��k3pb-�\V�}��~g�}�,����hR��u�;�CD�U����ȣ!��3�����5$�Z��:_�ab�1qe	]6��Y�3Ϲ�Ss"�s�}�dk�#�K��>�5家`�]��6KYux�U����L���i��X�*@����g� Z}���	�C��R/9�d�J��T�M�E7>$H��uG�L����Ә{��.v�O��B⌬1-$�ц��bO�u�W��&���T�VaY�PBX�-y`��6��~ع�{��jl;��/i⟖҇IT���y��X�-4�^�;�����g/H�8i��7��Q�y��t�W����֡�v�ZRO��[�����o�˙����[5���m��ʹ��Ɨ'�F����y�g�+u�oy���c��$s�j;�S��1��-�u&5�N�����o��ѥ%鼚�z���aZ���� Џ���T��R����|�t���(���s��s՝��9�2�=����o�������*<���=mq�w	�U�C��;}��R��ؾŇ��ӻrD:{s�谽�Ʃ||��b�/w�KY�*t�o�2�6�I:)\�_Jv|�B��Vؼ��y]y֔��^�ǅd���ͺ�X�2��}y������\�We3h��8����lֻ�YԚhd��r��:���{�C	�R&�eJZ�Vwc��gW�����G)H�h�s;�.��j���H��4@;��龊���&g2M�MT�������:9J�2�̇x���4�v9I�%��4u�v,��s4wND�y4ˬZ6����8�F�2DF���=�Wd˪Wا8l�rS*˒�
e�D{��Qk-�����yk�M�h�+�S�nԪE�B��	�Y�w�p)M}�9�߹d�Y���W�O)��r�(c�U��Ùfr\�C.�U��k��*7��b5%I˒��,ͩ\��+w.�㖳��
��)���oXIw�fWi��.P=ly�!l͝�7���wB��S��7*_�mi�"�E��eLV���WR�y���D�7Փv�V1BSӪ�~r��H��t��LW=�K=�lD�
������ֱV���MK���H&O�0v#au��Hlq�-��5�;=a9@����F�9T�[w��ri�Y�8a&�<#���u���y��79��RA�2��F���'*9T���d��Ή�h�cB�CP��x�1�3j�$m?t�;�*�IU�Ug�J��a�;��j���.���,�?,�-5Ϸ�WC��Ɔt3�7�uhsǕyn��L��|�2Ըٮ�@G��=`ml��/��U1�r]��P�M�kD<΂���zC+&��CzP�=�+�m���p,l�7s����d��&��֘��u�c��{p�	����n�����B���n�����8��x�%h���N'���흵\wv�E�1n֧`���%	�J|��Μ�6:���9��p���V>t�_�P�:g�<��y#��^`�Ǽ�bxv��=�3F�DH�!�}Q<gMeM��-*��)���㕼d��	,M�n\�����/��p�t��m=�ƒ� #��3�
1\������o/�t�<ʻ�
�hЙ ή�vZ�X��9
#�[�˔�jt�j�]�W��8Rwѵ��&���o��}a���5v��N��3)����x�p��w8���DP�3^vL� �o���4�5;s����m�u���׸�C��s�t?6xgU=HOs��qr��7��k5R���̾fv�C`��_P�ͺ{sC���]�G6S���n�|������Az;��q�����sN]_J{�z_viλ�٭W2����$.�b5&��yݝ�@{I��Sl�Mԏ�F��]���.�6�mEvi�)h�r]�s�[�h�3���rލ��.�m�И���蕏+��cWS� ��O�x{�Ll7�!���f�b���;��
��Ɩ;[�ϴ�ܷ+�eu�����>x������K;U-�j��-�][Z�+yu ����0d�����~x܄!��w�L�&T�R��"Op%(�]u^�6	�7��M��(�T��p^�9F�.ެ�i��l��v%�����[�H�=�Y0\b��MW��E��\G��4= �1֘��b]
��%z.%�*�1����wJ�Q�+G*�\��q���Ž�}�+�Y��*��]���o�+��k���VP!|��2\o�Te�ׯϠ[��'uD0�¹v,��78h�!�{GVT�|��1fWd�F�`M
ҩA�L�[(�Jewi��q+�gf��GS�J�&72p��CEl�;-�MI܏ +�M�%��}w,oZ�[v$U.M�N�,�d%�vWL]/	
ޢg7�z�N��z�Z�b�t�NK&d�Mn���FM�y]m
l�,L�79�/iM��iS�]����鑮�Z(�����(�3>=�gL�p7}.N�;\�e�W�AqU�[���V|4(�zL�R�U"�lAU�e+T��j��Z����un4b1aR��V�[A�B�Z�+b��C-2�E+D�*TX��E���ech�Ҫ�T��L˄QX��-)��*)�F����fJV��b�2�P�Y��\J�TdƲ,1+VE*E	iAJ��J�k-1���*�R4E�R��tVN�X�}cu&�`b��w�[��ۥ;�W�7l-ު7��ea]Ī
�����;4,��Z%&�3G��R�9����`@r܊j�Ui+�LA��l@���Y��j�{BV7��9үp�Y����9��)�ϛ�M	�^o����`����h�R�J��a��ug^����g���;[������C�f��G��:����S���V�Û�8�Դht��
��K���4.s��2���2���j���EM���I��N$#!Э�r�4#�Z�<�ܵ6K���qe�/9.}Zh\�E�<�j�'�缱�(������ń64X���Iw/>Pz&�a�Ǒh��4�6��:8�����ѽ`�3���촩��J�uvK�L�Rt���C��P�un���n���}�q�*u���VI�;���S�#4R#b>��>��o�4z��;�Fta�
�sL��zYcU�S[�V	�eh��Ė��of��t�$����2!�6�ܧ��a'vV�T)/:Jpw�ЌҞ��ґ���"��������*��
��7�Ow$��9��B�"��[;�9J�Ij;�R<����Mm�"��r�Byvsv��o#�[�ek���L�����%3N[��݋Y9�a+�NX�Efr���kK�>�EEz�����W4���,�eK��j=���'o��{9�<�u������gu'ۓK��.���*�8�m�R�]��y��Ѭ��TT֜-Ǚ�l1"T�3�-�M���YX�W:}�jr8�nr{)�n�:����H�-L�+�P�y��U@�a���w|v������O����)�fS��󇱥ڡ���C,vyg&��x��|�#�zӽB�����kf�DR��cf�"�1(�]�x�/��S�Y���TLkx���~�51p]OMl�+��b�/�j�b�wě�ك�&B�kGS�b����uJ�=Kz�6G{�F����Gxa�p��mt����m-��檼�s��6�����4�<Q��Bn��K��S��kb��3��]71�u�VrH`�EB�&�9&�rv>�~b���8�Rla3���+*ky>N�r6C���i �s!��t�gܔ�ku�
u\�19XkC���=c6c��Hf���|AK��Ǔ�^���wr'9r&��!r�3�gA���6�"^�rZ�[a�i�d��ƻ5�����>đ*qg����
Lz=1+�ǄTDOPq�U_o9d�ۤQׇ�t:W~*h�*$<���۩�	���J���[�_ez
iop��S��9�]��B���¶����t��8-8��t戌9�Zp3��׈_i���E�W^���d�v�"��'^RRj�����D2��`eH��뫥��փ����À�љ�ؚ�δi�X�
o�2ӛ�JT�b@��!l���_u�M���V�8q�3�5���FN����y��aQ�qT���S�=����;����g�G�:�x���-��:ٮ���dm�$��s2�xe�ʠ�}�덕wX�JT�nrZ7�t�h�;��F@���������uvVr\��s�
_\��m�n�T�ȫ��D���$:�9g��t�7a���&^���k�PZ��E���栎��a�j���
��?s5|���Ct�'���ʹ��Y����؋�4I	��������ٳ�u�����.��z{�(+ ���w��e.(
%NvrՅ��� ��A��{�t#����EI8�fe�V{��$�*�t� �:�}���ɞ�*��!�;��-���ԫ�(3�"{����Fk�-�'�v�9�W����V.u����7ie�GP���Q�HL�^ԟd��w�Q<�X�:Ghyem�	��W��v�=�W�p�]�z�f��	]_'Y�үWhlcz�[����W�/ F7�S۸�6�~3�6���N45�zvS)ž�
o����Ҽ�r|�au�{�Ŏ$����Ew����BN� �F���G	.X�:qN:|~ږȕ�����d������)vG�5q]��nn�1�2y�J��➎������>V����(�bU��::Cq�nƜ��O��V���!z�ӢVFE�aV��U�]����{NJK��+i�\l���sI�|���Iu�UY=sv��+u��n�.'>�����J�n\3���Wn��OM���=�d�+�v�I*z�E�Wk��uc��uo`�Dګnȵ{�����Z�[t��u>�b���¦0�)b�o��/˅�9��6����0#P��k�&��tՖ�������P��^e��g1�&�]�.`��;����]�^��d�;s�9AJѐcс�G\A��l�g�n����&%��n�xD�:Dh� ��]/E�
m%J�V��Fyt�2�Q��=L��ޏ��⤝8��l_Ab8l�>��k)}��rf����鼫��"���~���+�^�2WV<-�u�vR�ě>��	;@��h�f[�����g����).:G�G�0�X�KS*�H�Ft<T%*lI<!�Y5�]�9��"��f-�SA"�3p��R��i�d�<Hls�+TNSm`lp{�u�td4�,��j�T-ҫ�:��s;x(��-]X���x����~Z^*��]�f]�}�A���u[	��Q�.x�L�б���/>����5��;O�l����/��\e%����)k�.da,TR�E�t��l�Vʜ�����j��4:�7�M�����A��-�XÍl��$���[�'�?z+�1+1������=������d��c-��݁һ@ƒ1�/�7���S5�q���\ο��m�ƝY{ԑ���;hH��𭗈���L-�������V)�jӦ*�Y�>Ε5NU^W[ר�;�A�C9��w�'F�.�w_)�o�mu�i]����6s=��*W�|`w�:2�{|�xm��)_�89�{o)����_.x��Mܳxi�KT��UجU)cfww<g�j�(`}�X�RDd�w]b�����&7�*4.�[Z';���WZ�k�'h�T��Kb�1�*Kb��lxv�nж�\'Vf3;V�.p)������n��}�Q���S���O�+W��Q>�j��D���gU�8'[��?B_��*|�5pHڮѴDܢ�}�=����SySM�|����л���uoS���N+�l�T�ub�8Fjֵ�/ݓ[Ɯ�Y�S�p�H�^-�k*|�e��m�X��7�{��M	T�VM��Wf^�6�3:a������e��΀���m1|:
��ԣ��&W1����+tץ�qB���Y�M�~�~���DLDW����t�#Y�B�rf��r��o� b��q��w�=���5oi�N��I!C�̄!z���$!g���	CX#�	T4�h���g"W�U)$^�۬��L�x� @�QC�����hq���4%����쐁����Kd6e���8O�G��C�_Fp�x*�����^���{&�i��
�ЕCRV}Lf�u0դ$!�'W�צ�<縋C�IC�T�B����%TZK���X<#��i�����.���|�K�����Y�!g!g�V���s����R���.'.�^���c�wu$�J�OP�����U�v6F���2Jυ�	j��O��a!VxV�1�n��y�� � @�[�����V}�^����jŨ�b�:��o!l�&T�u��M�}��Ix��T֗�<�߮F���O�{#��B�/��z�1��EK	C�T�ҵ���2�$�ܺl�{~�ۍZf�2I��ӹ�p���&����g�^��te����jow��7G*�V~�)Tz�m|�<�L�tSє�����.W#���=���IN���IҬZNˌ4{ف�h͌Yky��qe2o�UR�u˪��&i���pH�-*L�&L����à5�ÄN��K�Or��L����T��֏թ�3�}n~�0��:�:qxz���8��0���}
%o��
O�߲=����Gd|6�d�D����K�s�t鮼�̏S|_�ٱ�~�͔�C��ۤJ�$N��xI�8��`c̭K���>�7k{�i�N��_Y�Lp2�%]OT�f
���z�.�<aϿV�4��4������j�)���;0�1�!pu�0���aF�dL]K3�[0ljΐ!w���ŉ��Ǯ1�"�HB���w��;�vW��sWo�$!2v9&�FF�8�dc��-&jLu^Ӻ�b��I�%�N�nd���H�
����