BZh91AY&SY;�BNڭ_�`q���"� ����bJ��        ��)T�AQ*�
AB�%@%BHQRUH�R�UP��R��"R!J�(*D���H"���%QR�D(@�@RA�!DR��(�$T���T���T%"�
��R!JI	����*�  ,%))��D��S��*�UU�gT"D��d*J��3��H���\lTEES; ���'st�RUR$@ATE�èPU$<   �-+�*��F�V�
�FV�IQH��$V�Ul@mZhYC*��� �R�����Pm���)T�[���R�   �*��V���1` ��X� �`(6SU��&h
A2�������+m�mT�UI"@J�JH�   ,�*R��f+ h
�P u���+�� ���J�sr��@]W8�IJ���@+��w  �`�AE �$D
\  �p�K���UR�p����(R��C��

�\�P�p� Uښ̹� uJ.U�U �Np@�J���*B@	B8   �˕@(Uv-�(��s��$�����*�]'7� s��R�(�V�tԠZ�� P�ȹä�H��4�UE*�P�@�T *���   e�@J\�v�� �K�J 
��N�R�&�v��R����viV��

�,�JP��ƕAJ�`@`��)TJ	T�BHp  e�( )0�a�����+�MS�2` f�� 3%�0 Z�� �  f�(
	) U.   ��P06� 0��@�,��iX 40�P
Eh�����J�a���b����
H��A�  	��eX  �` �`�X 
&�3+ h���h )` mF h�b�� )(�*D��  8P�  Z (�b�R�51� �  MA�jX 0`4(  ��  T   ��R�@�@    "�ф���F��P�4ɦL��B�T����I�A�<ԏ$ѡ�hښO"�� ��(�  � L 5�13OP     	J4����  @2w���"�H��	l�����Dq&���(@��w�<���~~��@Xs�?�
�*�� @U� *��{?���5O�( �A�Z����WU w4*yP����og=�ӹ�?�a?�2x��`3~d?������|g���������=e�������e�/X�`:��C��X����	��L'X�`:�u��Y����!�C��Yz�u��=d3���Y����!���X��`z�u��XN��e�������Y�e�/Y:����`:�u��e�=a�/X�d:��^�����d:��^�`:��^�u���d:�u��`3	��Y�e�!��a��^����X�d:�f:�a:��C��`?0���/X����=d�'Y������`:��^�����oz�u��/Yzߘ����X����Yz�u���^�����a��C��[0�`:�u��	������S��X����/�=e�X����1��񇬝a�Xz�u��'X�`:��:�u���C���`:�u��/�N�a:�u���u���S�'Y~�u�� u������u���Y�e�!���#�s �U:���D��TL��������dT� �X:�)ѐ��=a�(YQ:��N�����"�d� q�C��=e�"'X:� 'Yz�Uz�	��
u�0���	�N��u�S���`�"XEzu����:ʡ��(u�C���e��	���u���`D�"'Y��=dD� �e � �YD:ȡ�AN�(u�G��aP�"�X����S��=d� 'YA<e@�*�YD:ȡ���u�����^� fN� u�C� �a�*'XD:�	�@N�"u���a��XO:�!�0�u�C�`P�*�XQ�
�`@��e� dG�������z��XU�+��Y :ʏY�('XP?2�����Y^��a�'Xz����\�e�/Yz��^����/Y:��^�u���d�Yz������Xz�u��Xz��N������̽a��^����Y�����`:��C��=p�e�!�^�u��!�C��e�/Y�e�'�������/X�d:�u��!���fe:�u��!��X�a:�u��!�C�Y|z�������Yz�������^����Xz�����N�����`�Y:��N�u���d����4��w�0U��{��j�c��lC�Fx@��ifppU7���]�Fdecñ�v���L���Y�Ĕ������Ɓ@��qۘeA�S�j��r��w�1d/5X���B+6H4���q����7�U��5xyYZ`
���3���Q�]h"^]A��R�LA� ��p��AX�ފ�[���j����nQʙf�1;�ьu0�i�p�ۥzA9C,
�i�����XK6�-��F�)��hͧS/|��c�zM1(9J�{�v��km���IzSSʖsKT���M�f٭X���*k����+F �F��,�,h��%�a�{lShz�.�mǯE�����kD s�ajlQP�3a�v�-^�J��.��3����@��J�Y�2��j*Y P��\�.�	{o/�@jӚʛ�Y%�r�����͚�H��m����3>��m�Ch*�h���YB��n�Iy��l�)���N(��P��S3�C09����؝Z���4��yG\Iݒ�;�;F��oV6�I.A�A��wml͊������/5�䅁I�o!�m�����@��6�Z����ӳ%�ɕ-R{@ҕ*������~i�`��tn,��y��d�
�Fm�W`���ЙWL%B�L���jZ���-�Yf�{2���mӧU[�{�\ߕ]\j�'���U����ID�{dm`���ُR�i%f����29�����@���X�J�c��B)��b�@`�A�'�6���sA�td��_�z��]<H�)��jD1#B遅�5iw��h{!��bk4�Э�KaVK�#1�h��*���Z�M�Ek@XJof'Y+4G�-L�r������!`���AaϞ��S��(l�j��7�����J�gi�ܑ�]*Ue@C"�i	-�cE��;Z��X�ՙjC"�(·2��iJ�7�Q�J��tk�N����0+1`�0Ln�̃�����[�&h�� �E�;�"�N��ǑH��*�d�l���@ĮB�l�%^`�m�ZTn�^�M1�77-^��Zd�����A(���E�B�+q��o7�v �CC#�'�xr,w+4.��,�f�hD�j�^��Q��L��P�����k5�L^�n���mkV���ܩ�-#4˻L���7$�>RH��z)����.���ș2�����qf$٨O[%�۶#����!���*�V\�fR�B �f���2]Or�_�J�G����x�����ڕ�����E4�J�9�b!C0�Ʈ�i�,Q�:�p���d�-4�ub.��H����р\)қ�m��p��ZZ�����Ւ�Cif�fb�b�Ҋ�	�wrnG���L�
��*nMʹAI��\�b=��p૙����%+N2�TVi�C\Ia�F^�tɹ[Z�^�L:� )�pP�����ލ�_���m���Fr��X�3iՌ��{�m��5H�M�t�ԩ%܋I�X�Y9L+L�ow0U�@�q�9#�}nm�دJ�S�*��+�;��!AV�0�W-�Z� ��7E^�6��,�FTǘ+���B�>Q��3U!x��?]�Ia�K+Z4�[��ͬRn3B#
��>��mYӚ%G�5]Ǖt��w-���<t��fYܩ�\�r�ե-C�gҚ�Р�<�N��6��J�n�fe$ѕ�u��͕4��$ڹ)ڨE���55{�M�b�Q3���J��Q6�V��,�H�R���Kr[R�})mKJ�,��V��h_I8��YWL0�k�d_+�w��:��,�.�K�L��)ʒ��M�j�)�ӊ������݉v��g)m�zՆ��bKI�P+B���4I@̘6�� �,[�.�8LL� {��J�^���jlh	Z�j+P
5wZ30ٙ��C�)m�2�=�p7\ߖ�t�l6M�OD2�d���c�a����hHџ,i��YL�5���]k�Y����b�ŉ˸Lf�yh��K@b����!)YX��TD̹VP�W�-�� ����B]�B�Ko%8�FZ����jCt�-��Z��vn���^��Em��M'1Vjnb��r˵�(!lnn�����2޺"R3M�D%a'�,7�sn���uw�8�e�lE6+d	�v��� ��=+#�4e50�e��L+6��p_�vX��"ލ�ܣ��31���b⩣���&��iP�,4�U�(�O��ѻ���NVӡd�W���^QMj	:M5?]� H�Pb��J��[�h��o$�tZiU�1�Z��{g#�ַFj��NF�Q�h��1���CYU����I���зv�U�"�`��x�X21q^ �K��`�ND
&���6�R�q�x��R�	��:��^�w����)<4��jB�.͊+�˙nTY**1-��3��l�w�ʢ�q����e֨s1��'u�<p�,1��`�VǴ�
�SQ"���w35 ���P�WN��WKWVko{#����I�w`HX!�b���f�;`�ff�Io(��(�`�*�am����^��V�r'�ނK�Ȫj�F��y[]�Je��9W����{%fT����t���z�E�2϶��X�S���6ȵ�&��%"�I���J,M1�6���Y�Z�Y�N�P!��3V�*�]�����*D�`횙�җS^��t͙xvT{Bj�I��{,Lk*���Hb�Y�Y2�/��ɴ66���u�����2�������v�L S��h��1�r���,gʣ��@�;�V�:�l�ق:Jnj�mw(LW[n˭�N"6�Ո�wUt�
 �Ku�D����N�$��M�h�T�)ˎ�2�3 J�x`���Ұ��������e�ܥ����E⫭���A׷�ucZE�H^#`�wak��i�XV*A
�/j@K܄�t�t��0Єއ�e-`��(kYt�è�>;-֣F�wO����V�y��՜���t]���2�SI!HĒЪ��qeL7C)�׸��FAUt0d[B8�nۼ��YM�b����0��f������I���ص����,���&َ�X�1��K�9���wܰ��r[B���"��,8�ݕ�]��X�-�+L��f�������m� ��rIXs(�	S6�X�eM��n��&+����-�HV�]ط��j�ɥ�%>��lɒb̤�Y�N0�Yt��[��Uí)i=�m�̊����ǭ�i��#6:�p~ۼ$��?J�AM�:���{���6�`ܤm\(�[d^����LX�l�R�;q�H�˅�D�ѕ�[��L����y�A:�gi�pm ��I`CmǷN=��c�opl"֧��Q�vU�o`Ԗ��XR��DTژ�wA�mP�C@{��M�˻t�!(4wwYG.����(h�Sӻ�84HNЅ�OK�vkj��KD�Z� sh�x^��f��� 
�L��ZEw�w��
r�h$S��3wt�M�j!"WQc�72��˨��Ł�pAn�b��#�Tޢ��p;��b45S
A���6�C5K�59�\ ���=ll��<YW��l�1��4e���!���>�ҥ�Iv+0=�8�v���4�gᬣ����y'	 �eP��U/����s!���+[����AYj�7E&h-��a@�6d���N�J�[A��yQ����(�HD	3	kq�D�e3��yu.,��e�	y�ZMF�;�GZn�ͅ�%:ͥ�%��������ՐV���ǋ�r�N�	�%���7j+�nKVrD�f�1=1ScA�3򔝔pB.P�KY�U��p\Ƣa��%����Y���-�V�"�?M��"Bb�ue:�{e1�S5w/
��:�>@�;7zc���L&h�����eWq����-���_���K]��fcC'��lT6���Ji7���J� ���YD#n��)e!�����u�/fE(��+l���Z(��6�K͠7�-4� ��)���ڴ��U��C)���^���J�Orؘqh8wE醥*�F���F�����,S�w�cq�w�j��:�3`Ѭ�v��;������'�J{B�MJu�&�gJwu��
�������	��N�ȲK�#-�vHU��9�@��t�QT�h~kf�m,��$�%�Y��.��qk��LO�wd�PŶ75�e���u����(��y+XSUj�R ��3P;D�"H^�h��[���u�CP�l�A��<GMd�XU�t�����gѫ��'�{0�m��܄�5~�觊�-l��s�ZpkQ�w[71*a޽y��Z���������z�ά�
�ekz��k7-���.��{���{-حu��I��v�ՋgeJ;�P�ST�8���WG5���V���2�;2����4�P�q;,�`�q
���j�'Y��t��2��hO�:^���zX�{5���[�; Ցmi�pU�҄���*5�&E��7�˩t�mh82էp%r���]V�MS�t��V �V#�Cu\œkS�ݐ��^��J�8�ɔ@���Ҫ=�Fd/����2�\�0a�Ò�Y�PY��j�В�R�K��8Î�*�r�E֚��x��P�b�ِ���i*�&��y�#��Nm;ţ�%�Vl+ �J�]�i�t�ٕ{�],�1C5lY/��K6����Q-U�2�ڸ�5����(lY�)+�9e�Ȧ�y]��4�07��j�1-#5b�71���-��bo^��������í��S֤"܈�ٳ+5�f�먒T�@����9�=��Du�Q��&o@'?ΠwGniT�cM�mk��~yv�jՓRkݱ�+1�NV�5y/ ���,[�lJ��(U��zN�"b#F�PJ�^�*KXa�7)�(�۽j�B���J��4a�K��QVM�#��gi���ݢ�4�{�c#�G+6R��S6�^���Hp%�0m�mn F�M��T�V)����X�2��*�f�~��+eFv�SpVB�Kz���&����<VR�D��J����[vM5Nu��2՚�4�G�iP��M��%G����F^�hR��i�X�K�fԣ-�q�`��jd�J4�4�k�I+(^�d�2�3VS�5��� O`Ul�fU�r%�@ss�A�]
ү+\R�PW�.Ս��ٓ
�02���?-�r���[K1�@������^�iM�WvI3J�dTVU�����Lč#���x����,^���W�e�v�L�Rԫ@{�@�3��h5��R�\m�P�*h[ʅe�� �ZWkv����-L�H�RӲ�GlS"���Â�3-%Kk&h��:Ba̧����d�!*�f34VV�W �c]DڄSp�5l^4�$ೕ3+1:V���Ry�V3Kb:�X����l��1)K\����dڔ+t���Z�b.�;���͊���[N2�i��wF�Ȩ�{Z�Ya���a���:�ꎐE��4��sR��j�n-5n�[D�/4Q�Ei�LV������B��I����;V\͠�K�{��b{Z�Z�ڤ�1ɡ�QB¼Ii�t͊�pe�r��&�Ig�V�+5��nI�Ӏr���9��ǎ�l:����or���\L���k�[�Df��I�!�ia*���d� pn��LRB6�U7ķ2�6�o"�Q7,�7kSX�� �f�;�b�I5q� 4E�rRW4��魭���e�r�ێF��f�&��h=�ݫ��d9��  &�
�X��i,����F&Ȱ*Y
�Xv2��n��r,�����M2$�I����D �K-�*X@�El֚�M����f�1yz�һi+WOS�.��E`U�cGZ���X4�#4�V���Y��ʂ�R�f�NC.�z��r2��lVF��/605����e,��@K��f:v��,~ڛ?Aж���*����!�%�ڗu9�׭G�)E����8�Xn�����H<B���%ʢI66$��n)(��5�Zo)J�¬
8�˟�ڽ?��E �˖ �)3Z)Rb���!Ն,Eu.R�1�'xO%�b�T�Xj ���R}z�p��}3��:��G?c�L�*�޶�^Ï[�̚�L�����B%�";�ص��9�4]�m h�.$��4p��.�P4�}���ҍ+z�%��FV�je��J�i^�w���6�N��g=�o����������ƒ7PV�z�13�f<��D� ���,��Rb����`������FXQ��ȣ�ٷ�����{��݊��\�a�(�Zȥ6�)��U78��p}~5�̼��؊���:ʰIF���&o��KG:Ƕ7�i�9�y]��
�_4���lG0.r��:�1NƐxZJ��gN�w�zwI�l�an:��(�.��n.7�_Sژi���#�ӴMA>u��Tb��{J�+'A���Ł;���៟��{ц�V�r��-|�4��b9�b雜�TE|��V+ƅI��Bٵ���<��'i0^�F/�㿔6��ęYc��'��^�ak{��z]��v�6��f�.���[�y4H���S8���dZ�xV7��KvJh�ĝ�&�R4.�Py�)�e��#[����Be&��ɘg��jy�)�y��T�[��h����K�X]���ժ_4�/g�G�*_{�@s=��_OC���bL��'�������R��e}}��"�tuj�}�-���+`�߶}��ȅr�%:Q��v�[�.B���ɣI��8�y/N����ƨ�\��7��������8m� w�"�cPŨ8���h^�ا�*�Z6�Y�/�V���jX�C����6��^�J0���'�`�w��0�����'OrӺ�qd�R?q�W��^x)z�ө��6�fִO�p�9ǜܟ'��_�T��e�_
�W-d��^���ǯE��4�R���w_�����~te�jkOX</F��Re��[,~���s����N�2J�6��9�w|3v�XU�V��:5$�������tB99�ڑ��˼����7w-�}MpYB��Xyt�𙐭U�PH1��	D]���OR�7ENӽ6ۆ3\���	iD��\k"�0�n��HN�w�����!$X����|iԚT2���۽,D��O$�XjU҃Q@냰���25%�˫"uj�|���F���[�n���P��-^�3;��9�����z�'���r�2�47o"�"��m#Ëfh`L�7��7/��B�:II����nX��:�����r*���g�4�v�h�c%��<��D'V�8ҁWNy�}'K��ʸ���wq	/�Ñ1o:�br�Y�#s9!�`�z�4�Z6�k�N��9�tV�W0�fr�DªVU���#(u�����۝�ۃp�@����"���|�'�9K����wD7�U]_2�++�:�R�s{uw*g
JP���BU��H�As��\�t0��3v����N��gjZ������9f,��A^�,�#ڱvh�=����i��Hr��lڼL�hV�;-V���G-�DZz[�r���JˈU��h���+�X�m�h���]ͽ4�핺of��uA���S�}ǼrR�����h���p��A�s�:22��t�+n�R�-M!���ۥ@�a ���iZ��efm2�]5�mZq]�#��8�%3]�0����.q��3��9E��$���mw%� �X:���W<o�6rNc~xkLa|M���y,�/���8ۜ,�V8sg[5��D�P3*�u&��d��`��������#9 �;k�a�B]1=Ǳ�5��*jB��Z[P0K�ݩƭGPfr�+���cü�g8� ���d9׳w	����[�Ԍť��2��ʻ���IqLnPՐ�s�<�5��g�W���d@uؤ:n�և���c{1;dD�f�y8�s�*ˣκr���Y�G+8�%F5�n��C��brx�u�X�wn֒�a��]�A�;uf,`�ʀ��[v-�q��ؒ��o{;�@�����wCC�����u�_����.�U�x��̖�cŘԳN���K-��C��_c	��6����9�2U���*3H��~�_�q
Ԗ�l�4�K���oi�g6^Er���3�;xU�B���0�&򡲎�HM�O5b}�E>;���J5v7��/t+j6�����U��P���i���hG#\5+��u	��}X�Y�;a�Q�	N�o3*f���_<=[�����.�bۣ���<$f�.����[v��۩��C�C�He*�[B=��vu�s�T�����su
ս%W=���:0�S ��c���[f�)\�(�2�L�R���P(�ق.ղ�V*�^)_d����P��� (ե���O6G�]��Ǻ��II�N7 3�2����4���ׯA���R�����ek�R�dU��x��V:*�a�`Q�;;�7��s� U��*�f�G�D����IJ�.ޥo�Vby`�k!���v��t����́4�+3�C��:���K^<�7Aղk����X�����Z�x$�ɝQ\iCO��t���Mt�	�T�k1����n���
�'��4�b��7����!���6.vv;��q����;z:���ׇ��:��sz�/�;u>��w�������'L�s���T�������s&t��$��%5Ƙ"݂p���`�[7n�Z����\Sr¦��8J�8G-�����6e%|�^�o#��o^�
��_%��K�ۭ@1��~��(���sX<�*�JP�z3��"gC�p[e��@tBy$�Lj槥,]EG򘢮�n�m��$azJ���}�v���"�:��yC�S�E���j�ڤ{��w���mk�^$śEt��#{���:x�
�ܙ*u����|��٥�B-M�y��-���;ǹ��񅜑X�q��8nv����7�LU�������-���%5^|�*���W0N�d������G3�宝W[�Wm;Y}JG���A��F�Y4]��u�Ç{����۸���u�Z��u��A�K�qIi�FP��V&���j
j�Qɓ�wg0�?����T��S�\)jgoI�VR�vа� CR�O��4sK�^NE�O��0^�pbl��gb���W�����\����A+=AhW}MG}A�`)���|�
N�k��m�ձq��9����>]7��d�J�� �=V�p8z*��(;��ӗ(�wK9��P�|;����+��<P�ȃr���y�&T�)�:�k9qm@�缕�[�Qe 7�g]^�)E�P�ws�*Zw
��F�:]�1�L�k/�F���6k�e���;.v��;$���Xr����Y�
ʱM�k���p-�F�v����n�<ܞ��a���3�52h뵓�6�P��������N��To;]�&<u�6zjY�̓�B� b�ltֳk�p%�~̭mw:t|��-֐� :�Q�M*�_	ռ8�>%^Y�իn�4H��3-YO,�e�Ο�R��k�l���F���l�TJ�;��E�o6=r��^λ���E����J5u�@6�Z^��#�8r<c��a���b�f$tr³%�,x���cflM.�s{;mc����(ҕ��.�Ԏ�+�ω��0o*�5�)�=Ԯ���|��P��X��\���M�����aJ^WZ�5Ԯ-��2n��]��|y�-U�.�� Z�[�<��L�b�Փ2^6��k�m5t-}�����r�3k2�U����ٛ�DMԢB���ԦΘ�[�u�^A�5�(�� ,��x�B���z����t{a��o)	����]��+�P;�؈����'Y+y����p�Bȵ����_ۺYl��W��K/&�	�|=nثM�a�gJ��r�vR�'
o�oE��u�ĕ��CM0�6��ް��B�.;�.l�mK3�MBV1���6Wr{awY-w�#��O��R0�m��6�����ej�/=��G��������Q�a7�E{E+���B�,���� ��/8m��b���L�I6�I`-=�f�S���}���~^�guM����R�u��V�msL���5o(wa��MY{�v���5r#�ݙ��<�s�_HVE�me^�oi���k����7�]�=|�˾�z�PS[��&@(i�qb:�����Պ�j-9b�\8����H?7�ʭ�2Cx�hv��1�X��S���n���9�����H� �k���cs^�v���vcJL��t�5�e�n��l.+����3)K#Pj,�hV��{t��"�0�"���̴UF�,]bL���R��R��7�ۑR��@�^��}fg_���JU�N�ɴ�ٮ��>ĉ�fq�������Pۭ����ͼU��X��yt�,��v�{:��+դ�XS�T1��R�_tCX���9+bC���*K"�|Mp1�ӭ�Jou�3:YsZ�#�l�f��{�|%9��.uIGE_7>㴵uD����f�nKޗw����afzW{�xe�3/* ��H�_�{#����sh�\�V��O<��qS�Ed�/r���T����\�u�[��� W.���ī��;f�X�t��\���EoP4�g'c�G7�j�u��pE�k)J�u�l|��V�WvM��yX��S�7�q����֗�7t�$έCk>(`;����;�y�q�S[��[a���:���|Viy�BW��d�ٹ�n�S]/grL1]0��u�n>�� K��"7auϷ���ǲ�:{��qfv����*����-ӷ�N�/W,d��z� ],�<���KV��44,��mmc�7��"��ᒔ����I1����f+u�jr��e�+p� k14�Dr#i`����+n:�ϳ����ݧw���W�
rQ��"��j��m#�`e���'.���}P����)!�i㉉��w��/���:�](�����p��7u)��A���ﺋ�16�n�͆W9D�=��%�u��J�,o�K�A�G�:�i�4Ѯ�\��on�-\;�z@��pL�Ǣ��`�Խ)_6+��W]'?"�]Y)�;�7:8wVڧil�F�X�P�4-]�e�Dк}|E���6����'z��ˬ�#���0�V�K�i��.�
�
ٚ�a[X���Nv����s���i�5�k;�S��9,���Jۘ�q�>x%��s+H�(P�!2�2�F�����jI˺�k��*�4X�B�}1��$eL�ڛƯU���������9F-E(�L�Z�c�6^Q���:K-�o+y��7�;a.n�rI�N�K��g��ҧSB�󭹎�[�;;��ڝ�u�e
V�� ����9r������3�%q��me�A&M/U��;e
�M�� �Pһ�h��w��]/�Xu�7��e�}��TM#��y��6�Rv�`>�õ��g];7���,�������^�u�����c�͕'�w��%��q�.��'�#s�׼� ���WuJ�׹J��6/q�z�԰�t�.�kc�d�$��
�*;��C�h��뫖&oR]Q�Uf���-vu�6 �S����=�	��ه5uР�	�Cwp�#|5%fX����6�$���b].�ckwN0`���]j�}	�����ڹ��բ*�%�]\��I��*�\�����DWY���.��j�*j��3o$��k�\ar�8�lZp�9,j�<4T��vc�t��fL�89�ݦc{:�N��驠!�芣`�u*<t�zN�;BN�:�B��nD��ҍ[KI����9n��U�측�7t�͝���[�5�b�ðl��z5��ցE\�XxL�k�]/��4�K�Ӈo+g�	����@i����WK����o	v�.5����IS�*j��t��b�N��+.9H��嫿e�ٺ���P�>��̍�����(�,%`��6���j�s�0�6,�:�;�S�ە �����SSrF2�*b��,����r��F�!Y��y�q��+L.d�/�Q�xh2L��.��wq.
�+q]{HKj��Z'��L��-[�����vi5�AI�U�l����)n�\7"�5MnTW���-�Sp�j�u������=�EJ���je�;t�A:��Y]��jU���7�}�T��}�+^F2�£���)��_0�J�gQm��L��	Ԣ�K�W�Ƹ�nX� ((��0��sn^My:��.t�.]�r�vk�53s+q^����+r�%��
^�:u�0';��k#u�T���g8��+U*�%�׭՛�ă��Κ���5e�me����U�a\�%MV^�;�9w܈��-��r*ʗ�jV��Ώ9��L�h���9*�P����
i�p��'������k+���]3��m��?|�]arTƊ�zGt���sע������KmX�#���zU]ü�xmYw����'� 6��w�*�̽,����h>Mv%y<q��94Bs��ɼ�Q=[R�Y�et�����=y�@�Umm��f.�����-�����B�������c�Fk��t�V;�=��{�%��\����N.�s���wZ.�s������+ �{�;�%p��-Q�5rsF�-�l%ڤ�K�U��2n�S�6�����\4�eڼ�Y�z���1:N���aS��9C��v�]��J3�v�8M��ʦ��gt��O,oK0�:����rӮ}�]}�;��2ޱ
���z�d��5Pڛ�(�5�F:�vP���o4��9�up���e�� �z~�T��S|�;��6�!�����h��T��hN��N�J�՞@����m�]0W�^�ʺf�W[齉T�٭�]PI[���d��i��B�vҶ�\[��y���y�=���N���R�����m��;�7+�&��݋���]�3_I��u涻�F��[�[��cלa���K�<kt&��[bѬ��d>u�Y��y���4n��p��	���f��t�m�J��4v��\��<�6K�a��.5���e�d��څ�}�`�W���C��;y��O��˹7{=�� q�O�Se��d�&

��`^��HF	C�f� ��2֐�=�1D[��h�t��٦�����u�c�NW���s����Ln���&��ךtK����4k+dRSȹ���Ϛ+w�Ttzm�������ԕ��CiW�E�u�<�IHww5�"�wpy��wwsh������٘A`D�;w;f���Q�2����Z�0�&��Л�F"��@�/�s���Ȝ�R��@�##���}\�P:�0e�J�f�I���\�aS
��y8*�:���R� M� ~B�!4ѭg�����-�DФPي�
��*D*�A�ti �S����w�J�B�Q�J ���ͬ��Z��]���TE�7��A`�,���4""�͹tC�-@����z�0e
�*.hl2��Q�� v��]sw˕�i��&�+Ty{L�UAQ��w�Q�t�T��^Y^0돕S�}�
��B�5�� VJ� ��p�����Q��0k�q�Ml?��]��#��C�R�t�������a���\�rS�EѤ���6�&0��*��Ud������" 8%e�P�6�	��p(�[i�Y(�L*�Ci�$uY�j��=�G��d�t����e�z�H��F�.�y(���g��m��x[����(�*?���q	����mmm�/E��eH��(���7Z1�;��Kl��|km�TN��I̓#�;
��\�0K�p��QS*�W�oL�Ѕ8S�o���X<�/R����h�E�7f������"�v+�7es�� %�G���Ώ�m�07�o�ݶ�]�{t�F�Pㅛ{8�����.�s����O����a=�1�t��2���QC�m<����WI���]AB��VQ�W���ܺ�E���Ty�v^|�Ď.϶���t�A��XfS����)�Թ{S2;��'HI��tpR쑍�\{q&Ѯ�8u�I�}���HGv��k�Q(3�NS�P?�):�3{۷
w�[� w���87% 0�ڠ�Lorp�:A�?i� ���ʬ�_�qV!��Ln��r�R����Z��p~��YNN��D�S�6�T���B���}/��I�.>sZ|)����@�5�]�"�j]�n���+�}ԭ@���u�Ƒgz�a�:n�\�[;V�M]�O9ᠯ��	�ʌ��oNz��H��mM쬮�|�Rb�*�l|�Ⴌ��`�)ˮ�ugd%3B���L�����̅ȑ���G�jɧ�w!,��3KS�=ڼ�S(�U��wR�݄���L���uܬ�j����A�f�f��ك����w=ܻ��nLܖ��H�G�eÐ�uZJE$c�X���\�{�p'}�X�W�����>��ׯ�����_________^����������~?__Y���������>�������>�}x�������/���߼�ϼ�����|�C'=�]p�]�E�]6uon��dˬ9��\�ֳ�� "v�gd���Huۍ�1��\�պ��k �|{>�{�*F�N�j�7�Z/��[���i��B%W�w֣{���s:��i�+ve���o3��2�Uq�\�՗ps��e-@�#'U��m	&+{�s"���t��̂e��ԓrb���TGM����[�&�%q�;,�ƱpL�WN�"f�"�K�\/�#����z�Y$b��ݾ����e
��ZE��������^<{�8aB�9�&��Q�mX�᥃�����,M�|c��Ҭ���{���5{e�'x�Gv�*�+pQO��.:S��'
Վa嵙W*b�CF���\�nWfpKU���Ya�Ǎ���$�
D��\g>������\`��V�Q#�{�/3� [�)ru�sČ���Y:k�Ś��Jwqq���{��ܠ���Okb��H�����馝�wS�W����ZB�,�AX��Jw[(���kj�$�}�$��Ʈp�{�����E��V���q>�X�}r{\e`V_hZ�f���|P�b`�#6a۫/\�� ���ͅk�Vx���u��'��7-7}�v�*�q�X��m�S-ϴ]d-��;�q�U�YfBY+�4>�D��ݴ������:1���1�sc�1�c1�c8p���1��1�l}}}}}}}}z�ϯ����}�����~�l�>�N]sC����D1u��iv�vD��>ȸu���,'�)wn��������&R� �Փ �qr�r�gl��锚$�Y�3�U��Vv�R��QL�I�)������r������ws��.Tk7{�U�+V��Щ�w��d�U���3�`�W"��+j�v�yEWVضOe�݅:�EAT9^	���!��4W%X/�m���]��Cy�6GTժ����/j�vZ���	���C�1��B
q���łT�5ΝONh�W�GJ�tM'�o>aM���0��gt�X�b�#-d�O�xL}�@l���u�T���}9���rܩ[��[�h`��3�V�b4e�S�;UgC�+��X!���v*N�\�-R��ʹO���c���aQ��yS�NM�Eן���n'�$f�٨ݛ��'[�$]��Eq�V�6�
�%�D�2���9G�[iu�3k�`<t�9��u��x[����v�o.��:ƻ{mR�T���I-�-g9\�ԮSwIrVGI���5�PD��(U��u0f��2�Xٵ2ӝ���kU��)o��ϟ>~��|�}����=�߮x�z������������}}}}>��������____�8p�1�c�1�c��1�c������������������x~�/?w|���A�ʑfI�L����n1�]�Fu�+s��@�j1�eʲ֭�[+#����;Ư��N�h��u����]�uҨ�4��W��G:�3:彺��X�U�	�v����.�lne@��i���jRd�.5YuwA�F�)�y����c�ΆJ{\�+m�vinQlg��Lp��(�;8����L����ˣCf��V�q�t���>�^�V��e�m!�nM���
���m����O�/�����ˡ6nN�8Y/�Ā5}�x�$���o�,��Dm�G����͔�
m�������X&ê���b	:�����������e�!�d}��d޺�5�i��J�Z�S�!�	�ʾ��о���ŏ�G�dn��4�[�r��t��Y3�,uGa�5.�=n㩱����.f�	�V�6��aX1έ��e���.������|����q" �h��y���l����;�#2���c7�#5#K[���Mˈ)�K�e�����Ge�ՍRZ��W�>�Ba�w��u�2����6ѵN��	�`J�菖��}��z͸�k����e.+j���w+J��˙�Vp�25�I61ʃܽ�'�5���t�fe��.�߇����|���}}}z�ϯ������������}}}}||~�_������������׏��������w��}�_��}�w�kN�lZA��@��Tޕ�$F\5q���u�tƮ
>���,����d�.μ	�aV9�H{���Ӓ��G����U�:r����[��������k��ŵ}|xw��z ����\u���#ww����4�f���D�^%{g;�L����]����Wv�Jl���;�&�ՅI���*�[.)	W�yn�.�JZ�
�N�]!��GV�2:\�� ;�Yw�̛w�q�4�թ�&�u��htU^�j�|�_V���e۳�&�/]���-u}s��ͺb�r)G���%f0-�����ݎ^�]�ӳY���w9���P���sz.x�
�wN����m�J��q��}���;��,ce�w�|g.��1�	�`_^w�ͥ%<ice:���W#�T�w2�ᚶ�swwIV$�䢻�P�HlzDa��/9�G7��醜�7:\uպ�]>�UM=ő�ǔ��(��&�u�E�Ș��T���NزV�Xv[z���污�z�v�R^�wOa@���2��v�]Z@�����F��C�%R.�j��3
����Z߬�]�L©tN�؀c�Z�b���,����Z����K�ӷ��s���q�RM���&��{GM�ڌh뷦�.���t��Z]#�)��ŝ�t7�￿G~_{wߜ-}�_����������������}}}}}}}}z������������rp�1�c�0c�1�c���}�w��K,����X���*ţ@��ag�WdR=�I���5n��ˉ������M �Y�VIז��-x+j�op����S�������ـԀe�`nƍ��Xj�Cz;R���ΗP�Q���du=2�h���8Y��R J!�8��3�5ĺ������9�9j"����-\/L�SB�Ϗ5��S:Ŭ
:�ݎf*#����V�z��Y\���D�.h�g1h��ˠe�����#&R����!�gnX��	��ʢJ��ІU���ܗ�H��[Ζmsf�H��rڳtC���F�4���7gM�k��Z�+�	��{U>Et��"�t���o�E4qn������Z���
:�wBKJ1���vЦ3ɮ�	&�Q�{��^<����3�?iN�k����m�e2��	ø1vL��s�$ъ��<i��ܘ;5�t@uF��	�s�b�o:Fm91�ڕ��
�a����K5U3�"Z9/����==n~�ȋ���9��)ۊ:�n�ED����Jz�	[Z�*���;N����(��c�%��	���&�(Fӹ���ŝ� �Ob36�ZPppt�t��-r�rG���k4�x�����.e+�EVV]WڊcN*�����q�xIu�{pg3���|�fe��g���X���,���e˺�q���εY�tw�qG32F��?o����z����������������������������~��?\������������ϯ�������______^���;�=�����������p�;���U����A��̻x�1���OM�5����x�#��؇Τ$�u�8�[�Y,ڛ�ە�͢��>��R̲nd�h'�-�dU�n���E��j*�-�=Yպ�@Y[N��T���@�gWdd2��Ӹ3 숞v��ɪ9	�[�%,�L��7�i�Q�N}���F�⭮�!g]k�run��R��,u#��6^��������DZw{�n�u7���G���j�+���$e�z�s;��]`�x#����;��X�]�ȡ�.�*�*T�{�vΐ��V��I��T�>:N������(=A�U�41Ӵ:�@���I�9Ҝ��ެyk(�<v���M4p�9lNۄu_ru��\ueيqJ����^Iˡl9��t��
����I���vKw����F]���N�Ƅ�sn���3��K�W�(n�t�au�;F���v�ؼ��u�Q��*����V�[�o&������"������&�T�.�g�$�(rH䤵V/ߪ�Nm�ս����W�I��[J�xAwk0���[����!�F��e��i\�]\۽j�H�[�hb�9��֊ζ��.t(�qbm�*�`�m����� ����[����l��^�m������n�����"�^dW3-m�SDja7G�g���q���oT4\���)�@Y�Gr�47�5�f��ڛD�0��c�	���		�j�,r�//�ڧ��߽��ݼ�9�񞾽}}}}}}}}}}}}~>�����_______�������Ϭc�1�cٌc�:1�g��}�̥ ���n݀�Ƌˈ�8���T��Uo`�XZ��,��y�
o��S�&Z���i<V���Gn�}�{y*9W�d���� 
���Gun��2��:!��O>�����Э�)�.��jWs)�!��˾ Wd�<��j�;7)����cSɹʞ�Z�P㦫�D�-��N��:>�:\�;^��v�u�7�W3"܅�ͩe�x��O)��WP3r���1gb�L����}7+�e�۴QdGz"KfUU\�q�l��*��׺�-R�
�VN����+yI'��-V�R�3���a���t�m�}Xn�[e�.�Xj]Q����Ht�6��S����5N-��{W��*/��B����i7F�ġt���f.�� WG�2��_[�������IW�9mD��i�}�ϥ����B��l��U �5�V��v���T)K�/���-�R��Y�O���HT��S$"�d�.\��S9}�]r�s��[k"w�r�N����;����gCt�)��X���}��*S.��<aQ�[f��e:����3xZ�jN��b}��V�-KY��R�kev~��kZ�{���!]G��]yb>˝��ج�$��E�F�]�:�pE�t��4,8�դtJ���Z !�u;�M��ՑR�w?~���=w�IK7�S��M��X�(�:V��w�r\�L�Of�-�w4����7��=������z?_����������1�c��6c�1�����Ƀ�1�c�1�p�1�rc���|��[�7�S�6����N�@��/24��N�{%Du��<)d����S�����g�k����6�86��kcЌ�{���3��y٩U~}�=�M�ֲHSG�L���U��� M��]+(!R�7�5��}j7�HU�����c;�h ���aK��/j�|�Κ���tBeiYb�[iJ��[��TƐ��_�+] I��u#wՑ�S�Ɍ�{m'�r��W��)��������j4�ݳ�[lRː�����h���>��j������q�5��伽�'f
��%�E=�T5��(�^L�r�>%O6�@���NqC�����N�#�Mf�[]�o�Sh���ܩ.����.��`w�8uW <���%K�]a�ȵ��j��8����W����d.�QW}�pp1Ų�FJd�4v��+�u��t�v���������Q֭W��o�agV�J۰��C+J3�-[+�t�8�7f���˲�HrKɝ��.�5�s�P������'7�ԧh�1�%�!�:�۔X�ZͥM��/e�����V�c�ݢ��q������{1:g��J�@�ݣr�cg��R1������m^��i.��Ս��b+�y�&Z�i�����3��߿�jE��*ׁY�UM�2K�yko���Xq��w]VgkJ�5�m^��]\��W>j�Ӻo$x�J�3���mg絘\QWn�)];s��kT6-��8�B\K�LV��@6��V8hrz��9���)J����*��3�1�	�DgTQ���ˬ{ܡ��{��/�G��E�P�
N��cY��6��Ύǟu*�ޢvD����WjZ�=��kk �:w�"2�P��9_1���[�Z��z�|�q5��̬�p�{F��k��u^�2�"�_J�q����V�X�z��c��o�'������
���5n"?n(U���%�����rY2�d��/]���c��uo#���e�;��bU�B7(����r�ʱU�;�`\�a;C�vur�UN�d�B������^� ����%T+"�Rz��3@�k6YԌ��',�E;�4��M�s��7,�K�;=���Ż��J� w�!-��	Q��v������r�v�' ��6]j��q�w%�<�U�
��j�O�-�+��V��WW��C"t.������S�^�b��km9YPLT:�E���B-c<�I����sJ�uj+u�(٭��LI�V�wy�*;'n�H��ێ�T������6'K�=����Ɍ�dc����+�����@���f���p���-��OF���F����Lh$z��=@�Di�V�ZR�� )K�T�_��˟�x�ZO�Q�ۻ��-��^ֽe�_��  ��KDLn�B�:@j*�T`"V�l�`"b4D�J��` �\b���Kv�MfS�:���j�O�[y���oy]H�m|�=��P�Îu���0*)]'�d���iP�֡��G
�Q�h�2�����$}[�E��{��w�P�O�s�5�.�}r ��k� �����]��d휆�K�c�l��n�'C(��/I��w_ɦ�ɻ�m迹,ݛ\�p�FG���;�ކjS;����N_(�̭���e��$�ɺ��vW7`���a�̓{w>�H�̒MS�:n��<�e^55u*ej�w�)��uu��C���
�\n�u��u��u���.�WAaZ649kb��m�v�3�N'Pఅvu[���jR��D�y6*�%+.�t�g��۷|�m��Vd�#��/��ҰS����HN�x������7�#�/�cEJ��tw���gK��Y['[�P���.��a�!?d�j��	����B�D+M6g.9�;m,K��$�҆v�֙!�7��6�� ��7l>��)}�.�G�\ג�45�4���z��v";����>Ssu6��dp���7�;�M�Wfu{`�0��-���yx��.%�_'JֻO����9JN�Yt��G$wY�p��}�_.���D̝׊�i�,�w�� ��G�h�ɗs��S"Nn�B�t����;�,	�\�����m�j�/��S?�Mh	��Ŋx� JF���L4*$�j�R��)1'MjP���O�Q@���sϼ/�����~�@U:
�A��1P[D_0nd6�Th5��S�1���ׯ���ħ�uIDGy�Um�b'IF�#Z�m��Dm��Q&��9''C�(�*���ׯ_�:��E%P�΍cc�5T7��c+LEkl��������c�m#&���ۜ�ME55M�C��d�����Q9��ׯ��ƛ�4MMAh�Ls��W��Q���nW5D[;X��\�sh��Zѫ[|�|��s�������6qO���ű�ܰS͸5h�\�5b�8֎{8����,W.nnd+[Y�g\�9�h���_���O�z��|?�vк��c\�s�lIˆ�Ĺ��U͢�lmn\Nw�9O��X�s��	8V1�u�G-(rh9�Uͣ���"4�E�rxp�m\�z�������~�c�+`
1b+�9ns����˟5�B���+��qܹm8�7.p�mr���grӢ9���G�)�)P%�ߨ%H�DA�=z�����煭�#�p+sV�&��Ü.��9�r���48a�[߉�x���&�8nq�l�[bc�8[p��s.�8s�sSE�m�s[c���s��b#�ʣj�3�E���ocw��|�b��I���Ȩ�k���9�y����P�?U^O� j�B���e��N6|�������z�	��#���혅�;zX�\/�t�)�')�1(X��,�#E��W�~�O��ri��u���埶��Sث��w�8��_:*����K����+h�s�5�`�t�Ɂ�"����p��a���n�7{�R��&'�s�3���������O�j-����#>�Y�u�]>WwoBK�:�P��;sd���.�w1��a���.<�h�3}��v	���g4G�wcqi�����G�Eo�8�U�:�>��h������y��J����կ4xɗ�}�Ι���/˔��d��9ha��+���94��q�Zz'o.�� �0}�L���v�;�$��y�>�ǥ�t;��g�u
��Nsjn����O;(�d]�A�����Xy;�oc݌�{��!�Zc�|�-rt�ύ���n|�5��{X���ힳ��wM�1�dN]��#�A���c���B���W뇶��1�e��jO?E�����{�m=W@���WAt�����R`�bKʵ�!{o��h6Ec��A��1V��>nxYB����Pޢ�Ӹ�&�޼�����mun�ՙ
� �o)�ȩN���bf��E=��u�|�j���;�P>.��:v7/�_�UNS�{;H�w��ڟ/�m| �޼�~��~[��4�s�8h��~�����3�^�鎊���usWϳ�L}~��o�]X��|�} ���~I�W܋}�@���ޮ�::�����yU���)S���WnJo7x��zw���g(����ц�F�t�\l��4��42�}a`�p�zi��akzu%��TY鉳uri��zY����אS�{�9��.Zܛ������6���TC�k���O��H.�7��qm���r����~&� ?�`�޺���}���_��Ce��ͦ�����t�sr(�8[��c�C;��t��5��ܖ��y`{~FÝ��W��#����֓��<xH��X.w�����z�G�<�=[�x�U�+w�Y��(w�g����»Z�J~[�U=������������{䞾��7�WƟ�u��|Ы�{
��=�l>���Z"�0.��E[[A��E�J�v���|�����@�5f;�]N��ro�.�EfU�|����*}���̢ݫ��Fk��f��	u/�ӑ�]%���'Na�	��0mq��;��9:8%٨ϗ�R�y'��s��o�S��^P{Gu��Nך�����Ԃ�P�L�����/_�5+�����q�z#,3o����vĂ~~Ǌ����Y���ϧ:k��l�^�k���mh.:�h�}��=�{*K�z��շ�د>C����}��=��ٟ��u����[V��t�.���ع_��Ej�ݽ�lj>y��|��$u{�:F���׽���uQBM7N�x�z����|���Z����_]�r����C�k�[\/{���V�@�3vcq���Y��'e�r|���r��a�E�����y�ş4��P}��7��b��fx�U~�ګ~�V��We���I.N�Y.i����yi�t���g�*��縫�7��c���A�{�]�kպ=�^�A�X=T�jS��{S� f�"��j:L���3)��W�-�ex��O�<���B�,�pS'qF�VT�&/�ޗ9�;yT�c�B� �?E�W�6�M��Zg�ܱ�YA]7�`�v��to���E�[�/�﮳��u�پ��Os���f��!^��WsVm�+w�M���1����@��f��ov�kx�(hk��~�~�S�ό𥙵6�Y6��&�rgw�{��q���&�w��s��Ab�����x�&�����.�7oҒ���GC�z��1���Z����+|fvf�"{�
��ג��n�ِp���d�m��m�c�M	�4d����gs.@~"+��7��û[�߯0q$н���㥈���=Z�N(շ9����8�)�"əÏP��{���di�h9�,��z�'Iʛs�;�tLߠ�N�׽��E�h}��;�7ig�u����O�Z�4��t�����X���w���~�>3����ptک�^��ɱʿo0쳻}|q����;��\��q�%���ٔ^�Y~Sp9t+��.�Geg��{�E�Q0g�k_��5=�+�H_��ޣ���q�_�3�ۍ�ݰ���tZ��� q4&z |�����.z.�֘+:��ʘ��aH_��=�l����nt�dހĞ��n�h��A$��l�s6Ծ�r/q�������^Dw�������\:�Cwuh�]Y�<�4Ar+Y���9iSF����ђ���j�w�݋����G#���=-ވ?mDܐ7@J���^u���,V"�PI(V!O��g�a��p�Q�}|��wُ޹�$⾏į+���w��[���SAu�3����9fi���{od\^�~Wd�->���0��X=^��j�-�O:ʾ)zsN�Ɲ=-A��y��#<ߧ�Gh�~�,�P�c;�����>x�k�;n���E�y��v�����T����W|���������+��3�ګ��yb0���mU�=�{}'�s��&*�����y��j�ͼ�'��Ջ�>��mj-tM?MH�z��c���GmvI��Ͱ���Szy\����j�u.;޶#�;���15mp([���w�i�]������4F������@�
[ڽ�V�x�ү}h��{�iu
<�v�﷚\=��%���
=��~�s�}������p��Vo�j��|��wR|lo[;�����\�׍�N��8{E�4��9�Eb�<t��+����x�\��"-�O%�m�;�dō�J�\:N9��e7��q�����t���i>kBU���x_m���Na�9������:���z�G�z�*G�^��}Y�͓y��e�5x�� �W�]��P�Ki��6�ޱ�'h��&����l�ՎV�pTJ�^�lzE'?:����(��b�m���M��ǘ�٬�������z����|�1�-W��!u����o�W��߹:����^E�}���Rh�rzo�,��T�Pt/�ק*�������)������<޿h�0g�Op�p�kKu��a��!��=�נv�mPu�v��g��{bw�C�(kj3�=-�n���U�ϟe
b�݁���n@�v��.�5��k���v=C>�|���N����¯�_���B�.���D�v�5\l��
�J�="ś���y�׋xк}��g ���byJo�\�Ef�}��WO��g��w�Z�(VK�g�2��;>�l�6rw+v�&Lo�{���N�X��=�Oߺ��+�������_>��{�V���v�6��Zl,�؁U���w�=��e�N�<�Ӌv�W�*k�&3\P��]E(�L޹�V0@V2�g��*�,����p=��T�,�	g`��'q5�1ͥ�s��S�d�/!���S��I_�
�B}���ت��������s6&Y򠊺߇yo���]�}�h{<��FK�
���|�ᣞ*�yd��s��s*�ۼ@����V�� lQ7�f2ݛ�oM^��K4�{O������N�1����Q�w���l���Nf e��w��+�����z��מƘl n�5�s�j�gy�+����^�'�w��U�r�#3�1�Oa��O�u��̚�p�ݟ>��7�<��&=�^2s�37oMP��s%�ḷ�[�g�e�1�����z*Ψ��Y��n{{��]Ԟ���tPW�c�M�}���y�?Vu�v\�@zz|�h���#8+�&�t�;��Z��q~ۮj�4�|N㴑~���'��g�!����u�%�s8P�g �����;�q�'��,��s�s��Ҫ�����^���I<n'��&��A���	��Q��3�;�7Oc��a�	y��׹�b�b
���D���4|x���`<}߼�SJ��cjv�nh,�-E��v�O!Kx������s����߱��]��("-`����]G�`�k������`��ë�˭�T@V�ΧO��x��cSP6zqVY\�^	���:��^u^�<=�u#�����e4��;�Z��P�=��;:=����W&��[�|�U���b�g��z�~�B�τ=�]�T>\q�y�^�R�^�}���,𧷖�x?yL{��6��](�k��@���
��F�3ʦ�:��8��?jQ��==7B˥�x]/���I=�|궟�5wK���Xh�)�����و�ޤ�<��z���Rr��v_����jm�qx'S��b�W�(��[gϕ�76�C��]�����*�ߦ���"��7������+��0���7k���U������9��/Ha�v���t�T�g��v�+�^�lh��D�>O�Q':pI�s=���?/F�Ǎ���X}�%���N�S������z���O�*k{����+h։��OC�	O��u�.���/��v�F��mR��/껯�錆+=���vϟp�G��Y��:�ނ����+�����oVTU�^i�}s�j%yTR�k���k�:2Csu"BJ�x��yR-8�)�s��;��s8�E���F݄��y]���p��!Ũ�}��W˶Vwa����6ˆ匽�^�yB�7qT�R�����u�M���O�����}�b5^����Tq�oZ>ֽ�C�=��^���Yw�(ΑZvi���'��\{�����;�5��[�W���xH�[�	s��Mٻ������=إs��|*A;�p	�ۉ�ڎ�i�M�Y��ͮ"��P~v�@D5�Ɍ��^�=�'H�~a���9v��?Q�>��~�6/�O����b]�5�q��*OH�,5�0������8T��8�Co����fc���_��1�b���1�ܯ<�4fR^urf3`��^������͵��怮���[^;����P�ˋC�����+L�̗�;�*o�'�t���S�����u=�u*�4 �;��^2<��1�/z�̙�TjL�x�ͬ�V�cH��b�S���i��oR��@/}
�/�ez�����z{z$�xu�Tq�Җ߼�i��{�~����7���-�&j��J���m��$�K�d����B�/I�q��g�P��g<b8 �9m��t�S�UX��ǃ�n����.N@YU{x��λ�Ġ�ǥ�`V��u�!�`��
�[.̈́��G5�>�>bY�<�WP�ߩ�]&��-h�h�}m�����ϒ��Y�>�A\���Ӎx�4�$=�3���~�f��c�W������{M}�Z|��}TGe
^�x�%柞2�S���}�9�+����[T���U����!��W+>Id�6e{Y�L�ٽ��������7���y�]-:��F�������y'�j�4����uSO���zK�Ν+��#��y�YY�<����oC��ȸ����O�:���ߖL��ʨWv�]��\��ã�~S�Z\�7�S�����Y��]����V`��}ت,�i�w��<k��[^�f�p�$Q�Nٺ�H�,;��h�pc��t�p�FEPku�w�?%���W���ogT́���nw�����H�וV�ە/��6V��"s��<�ʧ�����n�wPm��·�b;��o���� \ݨP��Kg���}�����CV�}t��o1\����L���6e%�M�����w<CAS ��;��zl�_Q�w1���\Ks�d>�mP���s�J�vqm;�����;�/�:�r��T�H]\�>�poS�4���J�5F镵Ƚ"��É��-��%>t^F�^K�j��OmU�S���=��I���-d5����y5�B�����u,��@hs],�콶�G2�o	���*�d��(֜��,=Kw����O5���C��x�T!t
/$���N
�[��)W�8�.���9V�1���]���A��ut�reg')��No`"NL�2��$��L�s�n��8é�f����>=���0�k�2��V��������+�5��.Ʀo7�:"'1L�M=p5�$�}�jNlh���ر�s8yw��E���<9s|o�7�+ʘ]�J�!t�����3K�V�h^LYk&�|��d��A��*cY\�\޾�amu��꺍ҭ��ggo���L׸�<����dy� ;t:�ˢ��T�=2VS�,F�WY��ʃt���. ,���ܸ��V�-*�
޵�k)�B  ;6���2�+�E�{�8���unKۋ3�K�V���ul�	cv6�<�0�F���\�*���e�guΉ��r���w����K�|�^�8{���(���@v�i)���}��VWL�x3p�X�,ºJ�������W�4��XC�[��B��wL�|�bdE�;*�o1��^諢��!(���<���[mS��SX:�"]=ï���׋Z۔�O`<p�D�r�,<�>����;��H�u�f�4WI���jٳ]h�!I�K/�4Ѓ	���tt	|��2�Θ,خ�(��>U��a�Y�Π;���&bX�M�g6�W22�'y���ǵ�*j�gb�؀΃��}OLS��6�u+koT�G��x�޺�y�6�2*t�*%>��W:;N��Wpp�g���c)�e:e7<Y:�������£�W�]�t]a��V:�������=��<֩H���$��o����$�0�B�������%�|���.��:������qͽ�3/UuMLY�8it�ڧ����0�0Q9i��ъ��ԧ#;�6s7KlvՉQ�L-�V��o@[��f��W}W��r["Z���a�.��oJ-�1$���R��u�͜Ȑu����9l���]������d�f�
�fb��ʭ�c�b'��q˻|����vN����v����6�Ű�����]��T,��S"Ѱr�v4�5��_=#��ūw�z:�F�WNP*����dk�t���K]���Ư�k����B�-mۥ]Y�5��uk���DchF�o3\��C�T�Q�xx��ɽSEۺC/X����x�hӎ���b_��ל�.m�;>c�h�m�#�j��m�V���l|y��y�_y�D�?9g��'r�3r�͋Iǯ���ǯ���qGc[/.p�&"�gF�:5�4V�pŭTG:|��m|���bM�G�mFή9�������ב�����*�UUZ��9��A�8�h��lmm�EE�{b����U�U���T|������||&��-��sW�����4W2c[9����lF���f���ij"��h킟�U:�������m�P�Fˏ��(�Ngns�5DQ��nrԑZ�m�5�ڠ����||O��'�5\�uc���UQr-V��ܬ��Ӣ���kj�Z�Z�LE��m�&�~=z��>m'����q��lj#���&��-j-��E�h�M؊uZ5��DU��[j�����7��'?_������s���ov9�4ƌɌU��8򤉂�m�DIA���O6cZ���_�_�+F+��M9��3�~r���\֟xh�������\ƙ��k�8���F~�h�\9DD�1mF
��c���Sو*&4b�����#H Q��P�T�����G����uv0��-B�t�]f�g�eaS��#=P�1�sC�a%=t���������z���N�vNpǆ��F6���0���5E��b�;�f���zq�UR���5EU��������{�`%���Pvud��s�M��H��O��/�����3�*˽ٜ���������JǇǆ�k��m��q�{�D]za�n"��[��A��L�F�d�/�5SWL�'�o��;������m�����w����?�o��?h�h~8���PP=�W6ä%�2'���4�w0�_G��~Ѵq�������3ճk���}/�ga��x�	����C�<��^��o�_������蹭�����pa�9�,���] KuYE�Ʃ�xil#��C66`nFT@N,u��d�)V��P�1C�s�g�:޻���|��ɀ+`K^�S�nz+ρmkzچl;*����+�3�w�	��{��y��a�U���dt��� ��2c[�uA����Qi��"��V7�� M�F<#��&��W��Vd��O��9� OkO��*Y>��ދ��v�/R�j��B̸�O�%@�뭜E���}{���s�>���ĵA�|,��.CsO��MwHӹʥ���]!��R�ӄS6tE5�B��p[j��PZ�A��nlhĄ���x��N�q:r�t��9�w��n�U.���,PC^H��"����
�1�?Q�1�N��gwG:�[´��w�.���W\�fu\G�V"�I���l��M��w�J
i�[r���������\�c�on:*Sm����0��v�h�5�5]"៹��/)�ةϘ�Kw���fb#n&eZ+P������  ��ݤ<Q׶�C�f��*�����Ǔ���΋����紩���t6:�E7�i�,6����z��觽*�:��`������`���G��<�(�J�k��wy�{��/,��3LcJ|�3�n��� ��
b)l�4V��I1aD&���s^c�;���=k�c��q����f�wd.KP����[�5��t�l8���n(�h�.,t�AC�B�ʋ�U���Z�o�[��c�@v�p+�GLVC61���a�`2i]�y��Ӂ���x~��ߨ������+��,��~*����Q�8*��u�����N����5���ӹv����(�<� n{W�)]C<�v?&~<��4^��ߟ�O�*��P
�[��(�u{�h�?���� S@����n�G΃i�-.���L�F;�������|p�\1R*�4e��h�=Nb<IH�]�	�@o>��Et,z�A�:�E'ҲD�0F�����n�à���CK>wM��`����QJ`T�R��N��(<�Y�n��`��u��݋_^Mh~���{l�C+l:�@�M��[��SUy	[��ٕ.�W��]��>e(�>?4V�z�oKf*�k��Ʃ���V�̕:���_,���r3Vm���
���A��ϲ���{r!�a�`�a�8�Ȝ�v5zu=��6^ch.e�K"�탻B�Ҭן5Լ��~�yB������"�!��wK���cz�\�P���'�ܳ)�aZ�튞mx��Q��J���s.ԶMҸ��P2�\T�cw_E��[��(u�W��]�m�5����<B�i�2� ��}�1A�1Z��9���f>���\�w>�yc��qT=�f�mI��~a�e���1�L���.Cv>4'��$�,��N\�PT���nM&<%)��MIn/�#�ɑ���s=y)Z����m\=�۶��}7,X`�uc���$���vDԟCE��G�K�?���5��Z�ae,Y�3�'5�� \vx��jBW��̻]��+x<��0�#^ڽ39���2&��;�	ȵ�2�R[�V�N�<��yƲ���nm휕%��ż!(7���3 ˟>�2�K+�d���rV7<���jU��ZW��:	��Y���`�-���L�P3��.���Hx�ր�d<����z�1�R�?A��tgB�������d�G�Էs� ��ƪK?�_:�u���@v��~��������XM��D�l�F�;f�m�	��3ݴ�ٴ-.�M��V;ܫ�M�"dq_�lӉL��m�+rp�!��
W0�C�=�"���夈�Q#pi|�m�KVZ�mP�bՅ��wY+T���?�;8R�r�wHr��s��_(�m۷�u|7���7�m��7Gx�lmd:#��Ս1#K=���U��r�ꂉgok��ȉ� aq3���q�ܫ�/���ѿ���<W�i�E����: ����q0���gN���L=o�?B�.��+��~zt~�,�&��E��������La�&�6�"�M���r���$^�U��j��Wf��݆�k�xku��@FA��q���z����kkc�ɢh�y�+
��7��UZ�2�YZz�m��=�3i>C@�8�D<��z iw����*{ĸ�p.��T�O�k���T�~��/Z��ל{��ɨ]��tY�:�0���(UYQ"��=C������!�{� ����Sq���k{T�����q��jSwi�e��.�H�~Uu�(�� W�|hnFP�	�{�Ȭ�����[W۹G��)j� :d�矢S��p*��n�H������ʷڰ27�
��T�����ڝ���������؍N��tA`6�@M�&��i�.+�<[�و��˟��k�X�|6wi�����������	�����}ho&m~�2%��RX{����J�N��u��N7�][�{��t��yyL���jy�W�F��5���NZYZ^L:�]�j�Rru��Nol��m�BM�>O(�e�9�e��0b�V��-��<�P�����H��˫r6��V��X��_}J^����.٢wj�=\X�S��U�H���j��? <�ݕ�K�.�����p�h��u~h�X��oXz�m������g[��8�!E�Ln�D;kM��V�k��2���Jc�F�\3o3���g��̣��B^y�P��֘ΚfQ��^��k�����]�.�־/s�M8��ф��
�.i۬�,]�593������( *����E�Hw�������7�/A�Zs%W���h�^�^�rY���^��\�����?��I�|�j��]��Xn�������]���gHx�t�lj؀,�Ǥh�q��z�p,3��7&ay�$.��.���r�9��bP�h�&�q��1ٲ�{2ô��kz�D�D���AR��\��U�Z��y!�Wǎ�MU������T�/��/҄X^O�������l���ɧ!<Dݗ�1�og!2�����7]�g�z�T��BƫU]�/�r݁�k�����{(�*���e_4{_Sc�O3k�Eem�:�Jط�7����e��ب|�brE�C�.ժ����PڵE�cܒ����?S�^ƆL�`m������ִz�ڨ
��zȀ�"E=����w�[�gR?�a���0t@���R�Z��1F:�pP�͞�j^���kz��X�.(EXo)4:Iw�U�u0e�iku�S��ާ��IK�0����k]�$��A���d]Kv1Q�-��|A����',�d:�ބ��,��z�h��}�d��9R��e���x8�ØE'\�� ��al����Sx�`����^��N���k欚����qn�1����ƶ0��FG���ƨ<��ec����j�m��5�,���B[�������K|�h"I�b@O��վ���'�4x�7�e�s4^�v��<�yW��χ�>5[����༩���b�}"Y	�In�7*��O@���`\+�5R��P�`����̇�s��;<iW+���3���y�y�ڽ�6!@�A.��;ǡ��5�l�-������l��M������:����O�l���z댧iO~*<X��s>�邍oi~wv�~.�#[�(��NU��&�;���O*��t)�Yҁ7ܨ��g��Bֿ���zpu�F�����@�lK@��݇o�)�w_v!���8k�-zˬz/>�2��`��n7<���ƫ]!��V����_�<we�ڨ��z7�jgٙ�g���T&������㣀�V	{�Ρ�^ 4�z�ų*�'K�lM���wv�=��z_�e�����++�(:R!�:0��+rY���O�ۦq��U��0�5��U�����.we[��t��V���U�ŪMP̲
�w �O�Q��mo�@zo;� ?V�n+�1��Bl�;�!{�sz�`n9o�}�t��0��Z3.�Q����r�ݘ�Э�����V��K���W��3`C@> ��f�hLٙ�2��fɘxh�f�v��7�nKPsl���^]�s�>.���7ΫE4Վ��eχڷ� �o\U(���[\�S�Z���/��䳖l���
�W�VC�nP��P{2.�%�Tu�gz�ԫ��ި��;'��=8��}�+!0�W�B�	�������pyM��HP��@��D9��@�Mb�g��P�}5Р7�[͇��FU�1�c �RuemxV�6��o��.�n��V�2������g�g���F6K:��>j��nS��1���x�'���Ƚ��'�v�����<d_�j	��k�"1M<6�:CxNlW��[F7���<���U*�c���֧[�O�1�p�JkS׉�0�9��:��i���ެCUǣ��6�8�l���,3�p#
�1�C�˨d�-��x3V��T�E���ӻ��y��u�s2��x�L��
}� yc��n�;��.����
d��r��}�S{�5�?w]v�E����
FC���<��\��L�7G6ג��*?8mp']��<� �kצ]�gf�u�i�	�X��V<�{FE`�&I��&�k�i�}aBԳz��@c�9|�f��Y��uC��c,j���l�f�b���s� SO:;�
|r������璵M���}P[{�š�v�ק06�gp<k5���[�:��ϹP+�h`�m�QT��!�����狲�s y;�M�m[���V&DYZ �۔�UW�=1.�G�d� �w`9�[&as���M��Ra�P9�	����/�R��5�a�^����_ �Ψv�!����h���j��Nn��H��,=^�P�J@�ȋ��ٵ}t�/�2w�لY�̌d	�gN��D�ǎ@x�xH����sL�Е:�J�c'���v�#�����Z��}z5Rf4!۰tP��������+z��2>:*Ȏ�g�WM��U��O
^fƴ6�ZF�O���i�x�H�j�T����ޓ����4����|"Q/y�uV�1T�̋.]��z��r98���Ck{�q��Sl@&m�=t��ܼQ<i�1s��u�)xa	�Mp�L>��Bk�8r3�_Z�@f�}c�� !}��H��6��W[G�������B�ֈ���@w�Ȑ`��;L���t����B�~��>
Y��j�=4JOJFF+�o�sr.���}V��7�뙝�}�zwƗw���?^ǿK�o�������)���k!Z��i��\�n|T�հ�Z���W�-w�	�B�S�8O�e�a$X�?x��P?
����X�ݠ��8����<m���
��OR��x�u½o
љ�K<��nC���.$U�j�V9Op����삲�6�sU�ާ��j@x�{=��B��}�&+��.�ɫ0v	@,�.nj�hm��(X������OK�`6��M��ﮯ꫺����;�M4�XAE�7��T�e�
�d\�H��yS�$��!�� �c^���iʩ�Y7�-�W[��Mq�]s�l��K��\��K���>�Mܢ[PW'�	�V��+P�X��<��!m~��3}.��>˷5I���4zɐ�W8��5���ͧ������(V�kT�0��4m�
�<ЅC��t�S	���_�dN��n����#|J�@:w%�U�n�UXH7�����ոX�R�?ީg��[ 9۞��-pa���6bWLCnRW����5=�x9!��hw�U=��t�	(�'c�i�*F����m�]��|_���0N�{�g����}JC��h��s��X˵m�@�-�^�^f�K����>sn����3a��]��P3&[m:�Xrz�4�ӬzO3,z�6^��|��}L��1>$
�P�nu1�ޘ��Uڦ̫���śօ�b�
7"��(tIz�̍�C���5���K�=#E�U�b��3�ly��qeU\n�i]��<3\{��ZD�Ij�Tc3a���;o�l���[hq�lb�l�_�U��Q,j��t���,=x�a��qج�����''���n�}3���c ��i4���"�9b�4�;���je�;zf=ڄZS9�$gN.����lt�i�#�U�;���ޕ�o�<��Hs��w����rQ�����立�~�;)�O?U/\8gN�J�Q��^�^9�*Ӓ�O~�H����������m:CoE�\�.�3�	K�M=��G�F�<9�OK������j���'�Z���ȏn�_��
Q>�_Oկ1�=;�2�[�Z�{��c�W4�z���ק���K���Ʃ�{�"ߠKw�.oi�S`Ģ�f�˺@�P���=o�C&��d��ڦ۔�m�fJrE�e��v�V�/�S5�R̫J�j�8�0G��h��=�I�|�fӬ��|*-=hSՍ��:f�k5��!�ZNf�ï�Rщ��,�5��.�Y pk��s�%�{��^�qi��T/}\e��M��G�w�X��P��i�ˠ"��n���|�K�|v~��/��p"We� ��;�v-x�g��$K�5bj{W�.�^�r���,��Բ�5o@{��Yּ1�M~�M[P�7�8X��v����׻B�'U2Uά3�;b�c(:�ɀIH�������(/��v���^�NR�:u��s�P%�nz�����:a�{]c�B)��%�ݶF����<��GJ��ʸ]�-��S��9�O{D�Ț4��dM��׏��ǲ���+!%jKvݥo��&�c��l� )�Nvr h��r݅���/GE:��M� YV)��<S9�6(b�iwoj��1�P)�&�.�+w�ԧ����Xl��WP����p��P�7�X�Я�/v�ut�g��ͥ�ݹl�G��B��E-�@���tv�Wf���Ea�U��)��E�H�@H�u���N����aVq�\4�wZ=nt�6�e������}��u�D�
��lP�ϕ�L1XōБ^T�Wu�n�����"�F�^�o��n�!Q�#dK�E�첉8�A�[T�݋Y���.�t^[��y�6���F�4Цc�e$�.e֧�_vn��ӡ�p�|���r�1Hm���R��M�:Xgm,��vHL�H��,�;(m5%L��<�ˬ��-�W�k�pY�V65����0k���("]et5������C)��C)�9 �t�k��;%cC���-sWc��}Xqv��`����:�0_�Suܨ�B�o�����ɰ����bp]J���aV�Ƨ�y��;�V.�x�3g�#`�Zh�����r���,wY�I��"��3������hm!��
a���5O��7��3���ޝ��\�:�n"�^ث�C�pNη�����J�[���h�Y,�y��3#|^��.�G��ѕ:�6r�ԧ��WI���Vue&�ju��e P�ڸh�3y��^��d�	)�]�OW��ԍ������_f�;9q���v�P�9 �JqP�[$��J�\����v���G'w��v�(L*^޸��ItZSr��#:j����+{3��S��ٕ�Y����.�,�Frȃu*�%�J�Y��W��eaw_v7���������N΁��*�∅F��f�7W}�gg.�����n���u���}�PX�٩{���K���p��Kם�t��C{��������7��c�tz>�u�������	n�.�i�3(=��-������0v�Z�;ʾCv�@|��|�jrʍ�H�OI������4�AW˫�)���bf�7u����7nfbrK��[{+�M��&�W,ʍ]�%�U�Ǹ�L�����&���u
�f�"��Y��d*�:8� �fKx��u�֩�C�0�\.l(j��V;J�ݳ���Wob�(��e�M�z9>']����,ژ�7�q����v"����-^�w����u
u�[���q��.�Z1!�z�������aa���+e
�{�֥߬Y�.}PeU�*_���`�z{I\>���".u��1we�1�B���Gpj�����܂���	>�g���p���}��V��=�t���]8>��C@�p��=[]���3)c�.��n+M�6+FQ��w[��9ԢS1���K#�HV�Wչ�k����u7:uk��p����:N�j��hQx/xm3�VQ��튍2�2h�U)F�E��2���e�"�����P�t�)tbs���3@��)c�l�B�	B�Z0����߳@�?�5�˝����lSUI-6�Qvx�->sGƽ��kZ~�L�<���������墈��xh���qQiŶ���mE��CTD�վ��=~=||"d�)�&
���4PO6����NjcX*��fu�֎����^�������G���t���'�4Q�,j��Z�%��7/6�IIg�������tTUI�=���b"�-D��"��گ$�O����~��(
b�(#�����c%Q�MLDV��(���b��<�6�m�Tsb?�Ϗ���/1��-hi�(���(�������T�Fؓ�DLMM<���'0o�'������<�$�\�֜�E1��p�TE���M+bv����d����>��>�>Q�3�m�X�����D_3����LIF�y��("��"F�*"���s6�1���j&*�+�ǻU�'�����"�o~�N��5c]&��p`!]5�m�ю��ڹ��N&v����K����-�]���t�;ݶ����f&W@��(���-���b��!�||<!�>��{�n*$c ��z����|Ot��cL��ܨ��g�խ�=��{	������3����뭶��{���P���}�[�|Z�:�=�@cW�P5+�l��u�W3uw�<��&C��t*��"�G��u�"��G��u���b�����lqg�wђ.[��r�v��0��+��������߷�CJ��-W�S����%�}�kv}%Z�z�e�ݻ'�����P׌�zK6��KW�ŵhȊ2)��<�Z���N��;�}�Q������tV�F�z`/wvB�7���	�\�{f���3�)�u��j����hX�;�e��V�ܢ��ӹ�z[EWn��8����*y���GS����t��\r9��<$�|��?�`�}�;�<�\���w�]����Y�̦�q��	B��y1���6��l���0�j�f��Y�wԎ����f����;^�F6K9��1-I�w��ېhs�kn�L��<��m:�v�X�	�:WkoGDJh��qw�;PýS�N��F��w\�P��J��O��ypv�4�U�Pg���\�Cb�]/�ެ��
'א�젥;��<��>0`
�7	���"��/7M�=�5=v����b�w���	�m�Y����#��,�gZ�4�d�i�rMؠ�)([����e��b���10u*2o4S܆��5���?��Ҥ���Fd��|��'
�|�2���N6��ƿ;�i�iS�P�'�u��Cf��Z��\��\v���iA�M��z�Nl�S.~§�!Y�*�9����ۥ�.ri��k9�x��go��t6=�V�Cل�<z��}*n)��Ph�Z��$B�hi��監fU+������R��cmLd^�<��b4.��O8����YFK%���	�o�V�}m��{�}w��p�~�&�Z�C�~m�e4��t�B�w*2�7b�Q�п��Ƙ�vo���:>}Y�ɭn��,B�5`ڙƊ�����{��Ne�z6Kz}}�V���r�J��=:�cg�3��{g�LIr�Y��v9��,`�3�<��L!��}�4�:�f��kx���C�ֲ
t���5��|���>�dw|u�4�?y�t���r�Cʘ�4�N	��u���K�0:c#1V�;����8�Ş�� ���Rjur���^��sb#�Y!����fowp�벚\NOc����$���-��goz��63�����11L���]�]x&�AB�`��wc������������V��+eq�0A��3�>mrʁ[���Z�W=���vN{��.�2��Ğ�N᧊ѩn�=%v�J����[�\�*�V�.T�ޭ�t{�aG��b��ň����e1s;�s.y���;���Ϝ/�����N�bt���?�jRL2�t����f��>��|*ME�������*�Kt�6o��]�U���$�w�3����M�Я��3e�P�'b��K�j��=��ScV	��@����&�;�圌#���5��Ё)�u�]a��B�1�̤i�^U�W�[zcj����T;�>�vj�@��1~�q,��S{5+��&!��k�c�S[_�����Xf�3�^u*�۾˹ww��Au���|��Ҫe�p.�^~|����9;��b������q}GO��-w1���@�5��c��/�CϵI��酎U)��*�Ӑq��ͱ��^�V7a�y6��6���t!� �Z'�]��҄��@Md�y�L.p�9;�|b)8���ͥ�=�3������t1�\,��BL���"��b�����}C&�mAo&$Gr�/POb�������;��]v��j�nj���"b�;�k�T�И��M����e����Z����{w7R�ֱ��GE%ܶ3Р���(m�2��Ɔ���>h� ����g����+�������k/Uv���8�k�:yr�]����|�����}4d���A�v�\��w�/�Zĺ]c\h�O2+�.݌�@��v�㲐2��Xo{s�Y9IK{=�7P� ohf�l�1����;��7]��Ώ�.�����|������߇�o�14�K�4��;*�7кi�9MغKE��?��<Lkqj�c���35���C�W�uS).���n�G�
����4��F�Ƒ����m���1> �g}j!�\��lV�Dr���v�cZ�t�	Lڛ#L�K�׺t��v�J�sͳ��"۹��-��4I���0F�#~��߫�|�~(W߫#$���<�r�KC*�����-�i����^~�� &�p��3ū6�e�s@"��4e.�x�,��C�K8��g�7��ѓ�hp���n�'���sD��/�=�ck��L;d���
�����Y����/�|c����~+�o#�q��7��c�z;Sb�S^���8�&d�TKY���a>[��N�^����H��g�t=eY����ݼ��)�u�\m󩶼t�,m�a'j�R�mk]�S�����EX���L�"q�nޣ��O������\��gf	�����Gb��|]���-eE[��?[v��/62_0���e�v�A���ہ~+��_|�ɋ�,}acTp�V:OI�����݅6N��un}ւ��[�h�_����+�y�eIH;�>�7�BVuj	S�����V��/z�Q��E�Z�+�7��R��@lZ��QnP�.\�Z��v����(X�޴��W�bVgp�^��Y�;�Y��G;n����uǓ�����z�g��� �X��9F���yh��߾�7�����������YXU4ֆaV���ec�
���E�z�k��a8��>�0���1�/���E�U+��S-���v2�zrđ������s�P<�PX��\�� ��j��^���^�!�H��M�b�M@/9yw�qЩN���6���Rx�##�[($v�������Z���j^;�ry�	��sm��ܫ*K��S�j.�P��~��n\���w��,n�Q-k�ݶ}��=E���)=�vhj�2�E�/���R�)�������3vF�'���D��j=����s}/�����Y�}�y�j{w�d��y�(LZ��a�i�(��ݱԓ����,}Kd�L�Sf�e����:)Co�*p3�׈�� 1��T��ċ3��P��/~��}t���������o�T��&\ߎ6��c��Z�`�ڢn�\�ã}��F�:��6-x��yb��\��xQ���,�XZ�J���Ͻ�;z��3�D3/'�-��x��C��ey���>}bYӖ�},�1������z=�CY~6��҇�+R"��������ь�WP�>�7��|�u������Y�^�sNj@TjI������m|+�ʳ��֢���˨	�Ӫ��;��\�]�5�us
�֔&�����*�&� �tvޭ�z���Y���y�8��F��vY=���4��9dK*�ғF7u���_�>Ul�0̌�́�����_>�����ޛ��R��-����V)v��!�XLX�7%�oM�ע��Yz�+9��E�����>{#�G�)�#B�#.�e�)���G�X$��egT0�� oܶ�mhaF����T>Dþ��ŏ�eS�:?F�~�hs��Q|O�ň��kGP�����L���Ҝn1͋���{���9�i�zT�8�������Sŷ��cd:Q�>�,��S�Y�YDh~�z��=�TN����le�3*=��Ǘa�^;,qwCw��K�m�
l��	3�c�v�e+��{�㸷�D!A��f�����3���L��
�l�f�|��Jr.7��d `��	����v���^f}wmU3;����5�X�OX��8ބ���_������m ��q��G4�,s��B�>s���+�Ҽ���S|6�(�n/m��ń�3�㮔�Q��`s<�Ti�)�ܭ�*ç7t�����k�<I�9�'���Z�aW�\{�0Ю�&\g���a��x���D���GQa�s�H�0�"9D`�e�S�n2�8@g,�9�/���a��:Sz���Kg��)"��c.�oF���J^�5��f ˻keD�u�e
yd�i�ܖ�S��(X��-�5ҧf�.�	�nš�h}��0E��{�D�K:�ƙ�{�z��76�Y��0Ҋ��r�۪��S�|�f�I4�5�އ8��C�Y��L�����y�~���>�.�?�� f��	��	��O{�w������}�s���w���b��<�`�W���ʡ�w����(Hxk��.���,L�%���Y2q����:�,	r���q�m�3[�L�����$#�*^v�O�����������S�?0�lf�q��>�灅���T�f5�׆|~�t�u:����[}�������{jR"gf|�����o-��ϗ������3o ���� ��Ϟ�Ǘ��Oe�꿕�[��>�����<Y(k��)���T��Z�8ݙ��d0��m2:��eEѣ~�kߪ}�;&�޸��d�xS��Xd�x�8��ŵ�%K��-=C;1��Вǰ�B��ʂWB��V4�U~��tM��PH;�Wy�:��Vi��$����٩x�C)���`d�^�R�om�,[�,���vk��|ǟyޛ]ًe��ݫ���������@�)l��rú!2�US"��G�(��aEE�mH�3Z*�Gnp&�y��n�~!9"��e���@vD����]0ҪSwd�g��)�n�ӍΚ�}ƛ��7^Ww��NP�5/>ov��� �:w�������U'���U�L�?Nj����������\�:h(cݛ7�Z��X��]/��&�T���W;�oh�j`�=��2�ʂ��
ޣ����\���7���{���<��?�,�2́0��̌���������<���FХ�^����5��iK��#���@M�Ω��T��x�)Ӽ��!��*�8���9��K�D�iIN��P�	���ğ����ivP�>�ѿ�|^�u�5;D&�Ļ��/�ʻ.�kG��7i��<��%�����`3�pj^9��Bm6*e�re{��;���a�zCxjS��������#(��^͠�43.�^���si*�&Y�,Rmg�׹{��!��}�b�y�2�������C��d:�F��P��ʆI��1^�K�mȗM���\�F���&}m"��|��������h�;�>��R��B�͙���~�$2��a0�(�{kcؤl�~�a�w��X�?������E�j�r��V��f���W@�~��[1�WR�=g��5��R����ݟ`�ܮ�rU�[u賜S�N>ѓ�V�����W��j[?œ��(c�o��q1m��)����[XA̙Yd�׿'e��4��4�v�Y�˷�s3f�-)�l8��~O}X�-a0̫���uC����Xt��H`�t?�]�����U�����.�;k���\5b�+V��Ego�d�)���]t����͢:����V&=�6e˺�\&��Xlه�f2��c\�T'W��勛����܁��t��������<�o��r�˅s�9Û����� ̩�8VaY�f &M{�ުL��۫2�4c6��8�o/W��p�m���z�:X�YU,��<5��t�$#�9��˻[.�aB��z0����۞#�B�4ԈOr���Q��y1j"Y6ߒڦ��[B�EC�:S��E�sXԪ�����d*��X��u*T�J=��7P煏]Йs�yO�l��[+U�'���|Q��i����G�i�O�
aڛ}̞3��6�Rr\o���������&�3�ckd�~��|��Vni�7����T��l#�SO��a����	�iΐͩ8H�����s;9kM�kX���/���ڤkG����" =��ь"T.z�!�������+L���
ڙ��f��/v�s��s����1��;A������]d���z/��'W��e���ſL?S:8�H��j��o����2k(�d�9�B�Xm�� ��0^U��}</>���̰��2}�`��_ �����G�L���DF�6�����g�dL�Nw���_E�f�������>��`\0d_�%ƣ2=��i�=�%8�H���nHkz�
�7Î}�R��D�mҶ��z�G�^��|����96��*2��M��Ov�P���3ݶr�v�p���̜ۨ���{g}g�&�[Xa/�,�b���qVwS�9^�u�8`�}�q��m*��d%���.�����W�}���2�ʓ�
L�L��(�u7 ��{�ƫ�霾`���͒F�v��>[�\y��̰u6��fn���4bY�oC�z9��7<jQ���3���U(����_=zC�P���:i6�1v�f^Fgp�,�զ<�m�|�ܘ
�M^sΞ�<���Ƴa���J�}��q;۝��+0xrծ��軇h�VOq�<�N���*A�v����js��EtmT���x�42�q�~@F�a�"} (�z�W�K��Gh�f�r������CTۻ������-^N��]qZ�Å�n��&}������Cyi`�§��C)z#tmBd����S�R�k��K4;�0�;U�)��C�wmK�`c9����^PS�L�Κ��pK�P�m6D����ճ[+���]6��ܟ�T�qw���52�n��zz�+�R�Y�b��:�uݬ�q������ž�fOΰ>D�+�^=�ݡ^�s����%��]����>��b����V>w�o\��*�-�Aڅ�\��z��S*�0T�eY�{F�f,C���=#�xyY'���������j¥�vm������M^���ܔk\�Q�����HrŹ!�T�Z���÷�V�M��/*�rm3U�t)�_!��>6
�w����ޭ��MՊ�8�A�m>���u����V��v59w���2îI�o�5g�C5}4��`  ���B��-r�-�t��$�/�DV5�^�ޕ������Xݑ�t��`�%���Wn�r��4�l�������6�]�2wHF�X}C�*3���Ծ�2|fu�7ծ����L���G�P��2�,�@v6�c���jFk��'�Z��<��[Bmfc�NL lʺ<�>�t��@�.A��,�۔_f�+�s�x��cp�>��Z)�Ҡ,���L�K;hp,>j�ܹ�.&n��A�R��(S�2w���ګS6*�GeMFVȍ�hrU戦�r���ሗӤ��l�M�e�)�*xŕ�ˀ�%�؝wN̡�`N&��K�v7��6:���! �7 ��4`�F��>"F8^�-�ݗ+-g7YR�c\b�.���IDC���/��H������AS��)��B�����;nwp��BSh؛;9�����
R���\�8q��,������t�8.2'���^���:3�1�k)���Xu��_;�P8��Z=%����db��Bh��irX�b5�fS��A3x*d�7����;x��0q��n�9KV/n*�2�j�v��Z(+��A�TWn^��	s�������ݎ�� �/L�j���۱B��z����S��(�׋�7d���᧡����M®���a�M�v�������v����R�o$�+n��b�߀�zB�%-�V;�عj뵹lV�jL�9�Br%i�u>����*j�ٰ����e��l�L�kxW�!utP�i�70�f7�jp��K�c�;s,��!r��l�{`Y��v��r
Fΰr7�M[#��ݹ���y�Gԣ=�Ѭ;Ox��{V����9#��gMx�j�[`�v��G,�ibڙO�JZ_b�.=��cl�\�7}�:�ծW[���z�;7�JW�_p������j�0Wt��x:=Ŧ
Y��Må��v�@�;.�m��:�C�^%I�#6�.��=6(LP����x��;�bv���5ޑ�i^�!�s�L܍T�y
��k��]OuL�y��c[YE]/y�x�p��cP�]��v�;˩S�-=͎�G�S켝1a�FJ�|�[wR�����y]��_P�MA�uw���rhѪ��ېl��xpv�	�sP�v�︀l�'���� (U?�Vf�E�)'3x_������x�'��y�^�o�6��Oe��x�b �K�An��,�m��]�nB��Vʫ�?zh���xsjmcmE�����&"	+X�����m��Sǯ����< ����* ��&�j�`�U��Q�&"�-�5���<z����}�|؎Z��"(֢	���
�����AI\�51Q4ӟ����T���֘*��&�N�1QLynY/�UD�TQE4ǯׯ׭�IE|�b��J�"������e����o�ܳ5���x������&�"<���M%$F�ǌDTI?BqCG�~�?_�M2�US4U�IUQ5DELDP}��f�����>�K���IQR[{p���4�8���|ڒ?3���||�O�E|��_ Ʒ�;C�Uϼ9QEAQ1�� ��)���&���ݣZ��lEL�|�p��Q�����"�"b����Z&��&+Y�_~y|�睿
��Gm�^q_�]A���T h��%� ЗnfB`�n�g%������dG1f=�eI("c{��C�P��*�
�L �
L7�x7���{��A�m��Ϟ���ױ�E�!��aC� -���&���h�Z�н���r�ث��	�O��N� )�h	�[y�����׆�8�)�
���V鵂z��F���ݪ�1���QlZ�a�>0^wj�	`]�]��DBO��̴hWr�.��mT�zz��kLs��o8�	Ia#�֢����η������q����2�҂}�RDݬ��\m[yrҬn�F=xZ��$�֑�-��`���!� �`<h���/y�L��[�ե�v�J��Y4ɦcO�6y8���8��_��qt(%�]�p���C���]�9-��ܺ:�I�Q�S�V�ӱ~a6�Ƚ�i؁c��=a���j��}dym�&W�����Ue�xCo2�zr�G�#!��	�х���O^�lqv�ՙ�Z� ��@��Y�[s�E��½�9X�G`�R��}�`��/�(c�k�M{�S�����Fc�#v{�g4�e�wS6��ͳ�Ȇ��#�۸�Exqˆ^l�q�o����~���GV�����Ocv`X*f��?t��^��M8Y��W�9���Gv�T�SC_��1Z�G���}8�h3ƻ���sgESW1�|:˿o�ƍz�Q[�1.9�Q?�m����ػ�&cY	r`��J���|w�'2=�
��W�}U�}}_}2�L�"�!2�L����<�=ˊ��\�������4��U;t��;����[H�2l]�E��)��4�%�Z�^�ꮻt����c��25n�b�r%��U��U�œ�ow\���o��F�Tۖ�3��sk(y�3Ev�5���xR����\��M�T���`-]�q�]�xz��=l�Gn�����@�1׬~k`_�T�z�]7�R��)��O(J+�j�����5�����oA���UUXv��.�b<D�m��/�CΩ\��/QϙM= �+�,��h�2�5헳��뫿�O���ʈ^�[p���%��!�ռ1�S�����3�r�����Kc�Е�W'��9�[��A(��_��F���:�^��O�~�~ׂ@O�fK�y�nLjo.P%�-uKv80����0���u��P����>�C��ߢ�bW�N9xV�|x�T���Z�/,�c:i�nj�ݕZ�o����P��z;�"8
6����i��jk��r-��Hyc��]7{�kR~B`cGF�O��ϭ��;!򺦽�[�e`��Œ�Ԡ��?g�q��h��₱X�J���������҇φ~���6Х��&�dBpk�]q\5�U��N����R,
��,�6#R�17JGsq����ü�4�U�����W	�(Yڵ��uL���9��CW$���1U�Zi�q[��vw,Zl��u�	;��F�K�"�l��
+��&�Ps ��ʬ��20
�Ͼ���������md�s�O��W�@\��{ʥ:�av�{!�9�n�9�6����������ك:s܆h9�Z5I�?E�v�ة�p�=,7�l�z\+Ȭ�v�Y7��ؑ�3���<�ت��SO�y�9ӯ�|�]e{�~4=��N���1�|P���bۖ��ie��F���|G2��O,�q�C�}V�:�z��i��+����n�=s�j��'^@{�Llt�b3�����y7���LtS�V�MG�kf�+ׁ�N���S6��]��T_�X;�ʧ&�¾(�z���&��v��b]~��Y,�Q�L.����FS�*�}ZA��M��j�l�*�:��ԧ�*��s��Ja᱃u�55 �s� >z:�XQ�	�lZ���2ץ�I�9�K��g׆g�	\�L�稂-����t����kg��[O��x��0~�S�59��̆U���g.Nr���]��7)��V3�&�kI7&^���Hg�0��H��j㙻/�S
Ǌ�l:��qeR�Y�eg��������6sHV��©o46v�� � �K_��sk�_�:k�t��O5��c���۬�����>y���:���Y�u��B�Ɯf�RR���]<�}������m7��6���\�Ld��oK��'�˄)+U����uGN}��>��~�����2�2 L
�(̀"3(!�������l��4�3� 7�y���R��3�$������tke�دC�w>�1�5�7W��"YW5���:e�1���s#~��i�5����{��2k �%���}h;s;ڷ�/�����9�>����B�Xr`΋�	�S���Ȯ�%�p;<О�l�����i�!T�]���<��3?�h?R�I`j�C<t[5�y�:n��q�9�i�)4�9F��O�� �䪬i=��VXC�֐����{.� l2��G�![���I颃�ʞ!���v��e��ݳ*{�~j�$�j�]3����T4������W�A',�+p�웻��3k���kky[�&����uN6�E�=x#H�o�+�8�wЪ�����Ͼ����{��2�0�^��a11l�z088�f|���+���fעZ1�|��i�5����ɇҮz�
�^j�P�O!�e��=Kո��w����i�,a���A�4	�-�n�r������܅�LԻ��7���;��wΡ7�)��*}���z���Pr"�}c&^�cĶ�d/����EF�Ud���*�w��=j��Hy��WH#����)��n9����U�&u�N�b]֝bN�Q��rJ�׭��Hξ���4k��wT���L���5t��]�\��c�_R�
��[��x?��}U�����\���,�	0��y� o7� ���ob��6��c.i���g�}�<�����~���l[�?�s����Nt�E�Nݽ�ήJƦZ�����<��̑��M㋿bچ��@�~[�;�֞"��,}���[v��gdf9�c�LY"}�2[ɷ�f~K�q��@vfP�s^����|jj|�������&yUq=]x�C�;Y!�f4V)2�����2��*}��f�m�;ƭ?n��@X�'w^������)����h�L��K�e�C5��L��S-���&ӱ��7!�tW�2�sj���*%�-@A�}a��m�0o8�yO9��oV:�M���R�PjK�:󳝏K��kn�R�jz3� �&�	����M+4�^����`�V.&���8�n8��起��\i1��%��%�!1�������O6y��3'E�d�Ǯj������t�2����j5(R����E`�������q�h/^.�����n7�Cf�u�@E��Uʞ��e�:�����׮i�Mɘi��rqD�5��<Ϯe�,/�ؗnWmg.��z|�I�o3Q���,:���_d	ʖ*`�q���� ��}�W5���Ͻ����Ɗ�����9���e���=\�0��a�]����d���JH�+�y91�{]x�<�_Q��Ld��+V�kP�:7�!L��:�I@�_��dD�@�VeD�@fAY�F`<�������>p���R�)]�t�P'0P0e�;MA�5�W3�t�v�U�jU�؈¾�4��Ι�c�=�P��0�L�4�V��Y%>�<���$]˴�cǴƀ�D��^����2T��4sN]�n���
b�7�}Ʀ��M�#�g�e#�|�8�ر�o��;feS�Dq�پ\����e�a쾆�ℌ�Sn���0��v�A�['l���D�-W�٩J��br���N؇)���I���	��WB��ڱ��g��.��Z(8l��V�����y�n]v�=N!:���`i��x�L\�wl1~"S킧[�e8��z5uD<�vnN���qfü�/���C�{� �xZ����L���\�lSeu�"�35���nʎ�30����]��h��Ƕ��-t�Ny���h�a�T�$�$��y06����]j/�&�5������|j.,����*]��s�5�@{�s�>�u)�7�t+3�T�]������LsjP���*� zux���$~:89
�y�\�-�q=������[R��j��s8��#��;أ��v�r,X���F��1��Ljۙ�&_0������� ��|7�8��C��WZ鹜eڍ�@��zN����p��F5�ufZ޹+!�ՙ\ޛ㵽��N�������W^�7���}��~׼�G9�s�����P&EfT	�Ba@�A/0 x7�����ݢ�7
f�a+�ߏJ(E�r{���.�J����3�b4F@�gZ�箢y���|�\�t�ͭ=���sJ��T�P!��g�[�Tsr��%� E�R2���d<��fY��N���3 �\ax�y�K��/-���-{�Sm���B�j=^v��bgZ��˵͵�N���l��B�L��@��p�G�)�*z��^�='��ͮ��&}M5�-�ȊG%#t��*n��0_�EJ��7,;kϝٲ�n�a0��FE�����8>}Z?;×��> �
��.c���1�����&��媼9DJvOA��
Ԉϡ@b��D�p�k�|��ְ7�j�Y�e5՚X����s�l�韇Wye�������0o����v�y
�K���-����~�o��,�{�Ӷ�k��v��8Ƞ�ja>s�YZ�K���)�����Ru�P�d"৯MG�}QL�9Mz�����̞�Q-����"��{�cnl/Q}{���f*�����Pڦ"5�1��a+5�y�۽�\M2m�[~�m�������X�s����\������.:���-r"�Ͷp��o�o�؃C�Ŗ��ƥ����I�y"P�M�ݶ��Cs�������q6��#�;�z8$9٫��S��C��������Ͼ��ϗ�o/~[�����L �)2L 3 ���o7���(��Y�bxo�9�.�����~��&�[#�s�ǡ�	�?^e��XgbDм�����s�ȦĢ�銸��y��Dy��5���o>opg�Q�.�y���7��V�����u��t�:�	�����,�a�\�r\
 �z�{kiz����MC'�oX�K=t��R�uHf�[�R|�8Rb�����l	P֐���7P�{�_Ph�Xw���w�Þ��չjqϥ�42��M;6㍿=���BWψ�ϊ1�Fz5�*�\3�]��/+�����`��30��q֝�NÛ�网t�.z�-� G>E��7���L��G_�ϛ���ED2���N=�̮��^l�i$�����ӄ��B��8*����Γ�抽4.�:����gYӧ�t/�r<(��<�gy	��*�ߟ�`?����c�6�n�9ha���=�":��#W6�����hc7�y,�U��q�L�d-s�������V���U�	4�@ϕdV�뛳�g����Fu�꬘^�C�hjz8i��Le={�Ff��sb_���g3�%� A�5)z�j:�8�d�}��ɏv��&��X�9��7����\�*�^({S�O_Z� /$?dA\/��N�L!��9)=�+%��u���Ms��!�̉җ��b��դun�/y!)�ˡ����M(��=�o���m��v\r<|]������*��,�#0�@�ȣ2������|�����_���K�$>6ȸf�2/g�7zq���]�����-�<s˾�T��Kn2}�ry`އt-�L@Ҥ��d^�?�=P͖�qg4�fנKF �),���&<��ۘگ��w�C� �c�j&S��r��{�(�2��5bᬞDmL^FW(A���>�mp[o0r4j��5�Sn��w�#S�:~�~�C�:��W����CaA(V�W4��� ��YDD�g3��(�z��髆Ͼ�S>�b����E�DF�=� '��hi�<T[�����oF�nWpi-���kj�ts.{�ؤ�~K��^)�qw�K�r³a��{ol����N�h��+^?I�[�_�ʗ.�����R;�Jl�ʼ���*�|���*�����,9G��BggcƬ����vq�9dxl�+�6�3D�o=ٞO}�m�s����]�hYB9�X֥2��7�y�L�,qt��m\�ש~y�`�f<�:e0��ľ+��LVT�x��nFR��{���%SJ	N�N���|��l8M���_���e���'�2��Uź��=�R�)�f�4�sWz�lU�p�.s�Ҷ�5�7*w�5 �a��S�Y�!p`A��傅q!�\��C�&s�\�j57{z�ͨ�QZw�vp��k�m���)���b$���P�~4�2��D�:�C%w��o�A�DI�`P�&	�BeP�P�Q>~�VwQC..5s�R�,���-����<y�|��,�Z�LF���)�\{x���8ƺ1�fNq��B�aV���Ƨ����YRXH�*u�3ok��.�iu����'c@�`��[+o\5Z�����FIoO�s���2��^�j�Mi����v����2hw�v�M��.,Kr�}�XPZ�\�sH�S�O���x�-u�y�\���lK�u�h�j�E,�
\�uoW���"G����όd|pS��c�>z8���M��`��}�W�E��ߧ_�}�z�4��h�q@���P"��8\P�������拸v���/�Ξ�<�M�e��k<й	$q�`���s�:]�1o��Q���T_�8�ز����Pv1=<w���_E�a��.�2� c\=xf��"橷p�9]C	هl,��~gML����f_BɰJ�;F�D Zъm~2ޗ�!4O	���cެi��!�����޷��޴�z]*�km�U����6��Z����P��wl�.�)��H*͋���0��ǀ��\�醇�����;F�vl�w�s�}ٷ(COX�B�@��H����LV�'J��쬘ٻn��Sѓ��Da�m-��\����Rκ�-��i�)E��l�E����^�&�-����*5;s��WS5��m=o�����`���ՇZ��[
�tT�P7RS�+�(<�,�VөkvK�nv�]Y�%ug{���}�2�`>}��{L�}�R��^g&�'Y]��Wݢ�%\�(�!φp�����wue\ĵ�뤠)�8���d���&h��y���-RU�ܡP_mb���l�B�زK�/]�����(�I%��>�08f	eeG�҈��hk7F�u���[�sj[z�t�T_�{ ���ݡ��uH[�/e(͘8|�/w��3hLm�}܊RtŻr7�$�r�></n��f���w�M:�
:�pVbhE�J�4��˾��qp[�5F�6U��[���b٬�%(�m��ԍ[�2|�X�]6���GΌ��s����c��(�8aPGl�j��"X���°�P�Zk)�*���۽S;W�4�ۑ��#7���k��U��y���Wn����)t�
�Uۑ~n��m�of�mlj�#�%_l���N�}>��ۋE�S��I܋�X��D�t�ga�{�\��KcliQ��"�;���<ͽ�t;�{��)��q��0�:�ҞA{,�)�K��q&���2�q��C�x2b|�ޚz�]]�R�)�Ɩ� ���e�_緲�l/օ����LҬ-jv��;�0�w��=
�FK�IV/����k2f+U6��k5��7�Ɲ��]���4�����0��W���}�F�4V�+�\lC:�����r���Q9���^�	���fk\����}�ڣ�v��
B9\?n�p�f���r�h1c�%\u)8FX젬�*t=F��ײqe���T�!խ�����mm���Ιհ׿D��F��Cytͱ�w�Z]�s�j�r��-��5���i���Yr_�͸�+���u%vk���n��/���J�tv�ƳV��N�f����3���t����)�I�Yxpf�<g���7������Kn�c�X�Knva띆X\���V�L�¤�
;�s��oP�[���^�gT�CW��P���0X��w
�W �XJ����P�uUҦ��;��8�ֹL�[� ~��c"<�ëBne-�����K2��[�]��`*�e�^���}{ڪWO�� 7^+#���b��:6��a�	�5^��e%y3h���L�.1 Q;���\κG_)��[���{V��h�ꕚ�1����BΩ��]��O9�%YC/3���Y�� ��T���f�����9�N���b�ꃸ���؅cΜ��@u��3�
��ᢄ��G��N�x�]oU+K@��/�AJ�>R�T�S^�G���)��� ;�J�h��� 	�HI4��AiWq[�o1:$L���P�T:uVڪd�`��R��ګ��j�.l��EE~��DM��������|||�PRL�rh����SQST��o�SDTLW�s���>>�ϼ�S3Qٙj
*����/l��5}��Qͨ��bZ}~=}||�g�h(���Ɔ
���wLUU<���l�h�QS6'�z�����F�S�9��"*�����3�h���X`��j*5Q�؝?�Ϗ����
h�)�j�%�����������h��������x�i�E�F��PUEA�U�mT<٠حDk]��ѯ��Q�EKYϯ�����R�QAF�b6̛�����)"�)�N�����b��Ϗ�����Z"��^ؚ��o�K�>mEW&��Qm󁦨�Z(�j����hִj�����9�Z�M"��1ED������y)�h��&jj^n�Ͼ�4(
�U0v�1+���+�܋TT�y1[56������5Q,����Z̮�I}]x�����*��<+nn`�k��/��_����T	�ʸ^|������?��
E�& 	�a��	�P Fh�O銦(P��WX0���zkge���p[F�8����=�2��Ys��M�E�h%�fD^N�j̬�2�V�^4?	x�ր��d����f/˨]������_�$�`����/p�)f��H�D��>�<+}�Y�F�*���*]��tٞ�	��g��1����vNCU��澾�[�e��^�E'Ƴ�͵�k�X�;@�zDux�	��z^��kBw��s{_ �R�<ޑ׈͈���҈��m�7�Q��@�;��y�҆�fn�o�V/M8x�}�R���[o7��0��5�j�(�����B�ЩCw�3ч�����.�b�����(}Fs����~e���B0p}1-}�)��vy�U��5ӱY��E�I�OVٳ��M	�ك[b��� ��!����oI�ck�zy>m��l7ƨNƲ.����=wLݧ�}鉿5�i��H��
#>�߆ԯ������F)-V�WP�&�Tk*�no�,�=�u�����Q�S�����2�)��,�h`���i\2����ә���ֹ �@{nҴ�7����o������D�w-�׷7��^�m���z<�ͨ�:��x���kF�b��,�#�]�uu����lM�k��G��}�L�)�������ړ�>;*��՗7�=��X�/rݴ�r.�ٛ����{��U�U�D&A	�`@o7��f y������I+�7�S5���^��}Co�m�D�
�O>g1�9��Z]�Y��É�q���G0�X���-�����h��N�ڥ�������+�O\�ڪ]��VݹWs����!�=��[Ǩ�<�5���Ƃy�xVt�x���	���i��Y�u[z���r����7&O�v����2g���G�u%+�Mu�F��M@��[�� Ũ�K&�g5����{����!�wsŵ�X��͈}�*L�PuƇ�?�
Wdy������:�<,~;��;�:�^�����{(�u�b����)�7�m���\;.��o���cP�R�>��-�v�J���e6Mݒ�l4�`�L�q@ɕ�Wz?Z�Vnm�����\��T��)��ï_o�iX�xN���oO�֔�����V���F6���_�E'���`f�75ym+�W(�Hl�c���ae��V3��{r=	r4����v�P;��+=�K?�t#�[($v��ݭq��i�"]Ї��G���K��.��d�����OK�T&M��$�y=��y�6�L>37��뫿od�+:�JU����͵�vtU����7\&�҄Š�ԝ=c���M�++;D}+�kJm�;���/��,�Yی&/T�a8��Z����Z��t���]�9�s��kvnvH��B������ت�.x�2_���~����{Ͼ�۟���#02�0�2
L
�*Ȁn5����_G����U�����}�i�F��W��iz���)����k��Z`^���yiR"���rr=ZcY��u�I�2��|xO��^X����ϻ�j�v��[� ����s�/�Tsj�g�^��U�,̯CB$@�D3b�{yn�Ku�za�]���
e�ly)��5�p��sN��3�4��7<jQ��<g7Ί��)��)�����>�ΝM��V*�ԁ�a�����W2�lh(��6٭������K7=3��@�6賳��m��m��t��h�]'���SMX���h����U��u���.��V:��y���=�>�]�x2��>W�<��"u���)�^�ŵz��mY�i�(rGq�k1#Kլ��4��%��K�!ޤ��ߚ�*b��=��Hʈ��^k�4��L��Ģ��L���ͮ�C��=Y��@��Yk�A3�iTG�
����l[���OǢZ��:�7���������uߜ�w����mc]2磑I��ݡ�E[��YR�wcM�oj��Ŧb����3���`� �W�������O3�hu���^�˜�g̲�7��u�i�-�b�u�)k��n������V�\n��95����H�t�i��ogf;���b�\j]��ks6�0�1�x�w���Ow�;���~��{�����|��P��Y�d �E�A��S�� {�f�%�(n���s��At� V�2j��;�M�F$��N�ʨ�W=/7��w�n:��Ɏ�4�'�t����?�CG��f��u펪6��)�?`*}�7�[��B�c�_�����U��w���O�%�a|@�Mu��h��yҘO��KqxC}��YI=,�Z׹Jm�T�qBsC>����%�Jm�Lݏ��Z/���͒:��3t�"�*�l�\����X(�x��1�;>V4O �����	��#M#���>�>�!K�VV�Z�razP�hV�8U>�po"������:��oO��cFU�Ⱥ�_g��ߖ��HR7��e��ޯX�E`��L�Zp��63����h��7�7����N/��7��_V���ݣ�O��_P��I�{����������<�_���U#N=#k��9���dھ�����^�ٮ�k�td9�F��#ゝ]�U��=J�d�*���B����c�T�S��Цeʫ���r�;μ3��G�*T�v�W����;c��pk���g��������xSs��u
��9�ۨK谞͕t⥙G_Q���&ԣЫr��O�|�ܭekmP[I���i�Z v/�Ȏmf����MI��n`F�^�˾������"�uAg{MǼ�{chS�f�4�5~�����ns�>o�1����ȁ0�2�0�L�� 
�  ��D�_'�v_�}�h@�� /�K�|: �W�0%��6Ξ�L>���d��0vE@ɨ��X�JҧV��-������<�;H��P�H�<�l"F���4}�ЭD�o�Lc���_���w��l��~3���j�]�mǟ,WL��^!)���M��VX�|��1\�<�0�{..��<�0s�/�Е���)4� �x�2u�7T�z9�v)�>u¼�g�	�	�s���ݭ�u����v ��j
��ʽ��-+�9�JD�}vX��s��_@g1�nW���|�]�/�9z�����Q~���`��9"��e����kd^�2�g:ǈn&cr�z2������3M�rq�6�/@���g��*]��tۗ4$���w�Ӊ�2�	��p����I��%�A)Z����@���2"!>��vq&��¥Mmfnl�k� �l3�ht0�g�e�k{	�J�.�� �]ndn=y(��-��t3sd���C,��֕�<R�qP�y�
f��]S�"Zz�T��@0������A�hL
��E�w���M��إ���a����x�J�e^d�"Kx
�9���mj�rP�n��LWV��۷��8���C���C��7�yB6�M'��G	�{�_S�Ϥf�4tѻH�V�v�;���*�Տ'u��1���������U>�f�P��f&P&DfD�?�{��=��_�����o���|�`��t�/-�"3��MCsR���ةO��`'9���-Z����Mr� Wp�d "��t{%\�\~������I��dCn�'��M��p�M3��^vH���e�E�����`���5�[kC;�g�>�e�a�>
0�|d��>,����&�e���A�� �j��Yz�Ҷ�y��+�E:Ԉ�!�>O�@&
��\�c��H{�ѕw���ܡ[q��Jy~Ր6;���[�4H*m8o��?��Cr�(G�=��~O�^xu]�׶S�����\&�wm��ڹB>g�~dU���~M~e��R�2�[��7쿺�f��:��J�UV���j��l���b��6>�^�lm��9`K��������kt�=�#��5�����Zȸ�R��̸Sl^Gw��f�q��9�Wq�ܚ�,r�"m����*L��(p��,�l[�=n���N`��M���Y梩�v��^n:%e:�
��Ϟ�8��9�]"�it�=�N45�.�y�	0��ƠT;nf���HּE�%8X��%�ƭ����iH*�=Ҧ��%���y�{0�
|���غ�ŷ!��u}];�}����uW�P颺8�蝷��Z���<o��k�ۍs�P��,-9��
iNov�6>?K�4`��������<>�x ��U�T�� &A	�e���?������<����o��<���(G��R���&&�P������W1�^�ç�L�¹1B2�ά���׽ѻ��|�!��\&h��`�
�j�9��ߌw��j�Ҭ��nE�qѥ���n'�&u���aM����xd�/�]���D�T�s�/H��wε�`!�K�?N�ġ��Q5	T�'��{�}���~�X��w��>g�/�Þoxwߡ�[�O�ӓw���@
����ϊ�jz�?b�H(3���������;P�/i�;� �\L�t�ǞUW5{�We[�ak����kg�Ls��6���?"N��`
��	_�5�yERa\=a��T��I�����z�=�
q���g�l�l�1l��`���7��=�����ۣ�}�k��i�~A��w�-�OC��-�a�z��h�.(�X������v�{[
ͥ�w;c���kt����x��\3^� �ǻ{g�3�w��z�AM�l3aXPaϽ�"���A�P�Ά��泍`-�ȉ�8�DL[r{�N���S�y�Tn{De�`s��+�>M�c~�ًi�
�� g�P~K��J�Q��R��X嗾;�]��'��|��ͫ{.��WpXѴ@e�s�=�⏼+�;-k}s��&���	�]u�6���\�]X�e'��ov�Wʺ�����f���6�����Sr�ʋ5Ҥ��q�*��YD�T��Q�P�C{�0������ൗh�el�Ԇ�q��4:<ڢa�^@{2$FAOR�n-��p6b�x�݉ƫt�*z��ne-u�aеPJD�V��w��nH��.��T�w�P!�_4��=�s�Ulڸ������	���s$�?������e_-��=�M>�+/·�	m�b�ݴ55_��;y��洼�Ήк�T�ѩ�u�xMmCv{[�I�֟u��X�W�.�-�a3y.ڨ�A�nh��e:{:e��yx�[L:AĂ�=Jq�V�H�锟s�O�7�ٯ�fP�����z��mLB��3/�Ӹ���]�w���)֡�{ �f0��l�'��)�?E����.��^��o�����R���g�R����qO�+��@�*��}�3�>�?a��U�A��a'���͕oaj��u���E�����J�	Lz�Zu��H���S6�ױ�L�̬!Fn��Ug[��PEB���kL�I�`��aӊP��<x����V�_=	���G���f��t�3�x�m�*��P���+~�Re��^8�	��cu�_),'��:������L�}[��m�EX�v1���s��ˢ7f |r���5`�|�CB��m�%�Sr��+p�ͼX�Jp��ِbǥwm�EU
+�,
_��#Ϭev�Λ�7;��c�6`���Q$�0��n�3RM	�n��x�X{J��]�X"T+�7s��`�Ç(�[|����mF�M���"L�2ȓ	HL+2��<&R�J��!�,����Z����^�b�O�#'����U������߱@j9#[8Ŵ��x���j�@�L�y�[G�d��0�O�5��%�<�l:��]��y��A�����s��~�*9,�av�~���d��v��������AqZ�^��
M��S����7I(�̉!9o��������� o�?��>�	zP8zR_����pT���#���da��/���c/ousc�e{�Z�#�hq2�o��*��;���?hP3�K
^�������n.���v5��l�ѹ��b�B�ℌފwc��
���Y�K-Y;k^�L�F��zs�1�TSt��XH�"SE�Bm�~�S����}Dn�򨾊2_vV��� X����v �'��;ى��?��g�v�\��,�[�9j26�l��5y;��V6<!���Cϭٗ<���������� PE-�kÞP�)��s��h`U�v�=�n�Z�1�"��>J�3��t^L�yO��j�@L��f~�F�N��-�L�ݳ��<Ե�w��k�U�ݎ�kxKO�,�[�E�"�?�%����R3k|�v�iLʹ�Z(��JD\���f�V�LTH�sN���J�j�o�Ãm�I����
oi�W܏fM鐉�X���ʌJ��>}�|�����7��_����@"L L0� A ����������}ۖY��s�Xv����*�3d�sm���m���[PkjT�8p#�&њ�V�Y�w��ۡ,�����Ws��N��>Q͒�=����z�q*��+�3ǋ�S��㻰/��t�&~��ߪe�M�2��}�����E=��s.��F㠘_���Nz:�֘��1\b�6�V�h�>��ƽ\)�K�]q����L1�������L&��9�l:}mZ*s���2��֭�dtB��ٲ�ᡣ�vC�x���CF,�����|��G���Ա���7}-�7����S�����"��i�T�h�F_x��<v�ϋ݇�5���9�;�(�4���`��oNm.�P U �J�?_�T�>����OI�"\\�9m!۝��^_c�H��`P��CFJ��;P�m^L-5}R����X�lۙ������=>@��z�.&�Cw#<��D��3�R���k������������P�f�9���[C�3��H�F��qA�˭�X��͛�[Z��WZ�#֏�u	�Ub�ξ�Q`�b����v��6o���8֤��;��<���'N�%�/��=9���W �ò�m�[
w�ocg�]]W�'f`e�z��+hR�N����u�ڨ	ٺE�stNu��z� � ��K�֞oH����[+�<ѽ�1n����;D�)^�PbB�Ur��y:�m�JI7���yt��`4�,��"V6�.�Rmo_'@.e��JO $�deh�!���f>6���{t,	ʟPqwZywWmܰp��Lp�}&Ȯ�*���L�ޤ�)���B�mi�U�ôKۘ��yA]�Z�	�p��cHY�tKr����PLe�S�t��`��	� e+ܻv�U�}��]s^9V�dq,+&���4#:�Yyӌ�͔���u�;�d��%������t�������K6阳y3Tg-�+���aףi_']]�N� ��4,�y�ܺ�\�����JS�BÙ>�&�gs i�.�Y�*�=�wc�8y㱜ޥ1)"cO�	i]�J���U���']XCiS�E��@�9Odx�Ve�kF<�P�P��R�,�;���(�遻���eMo��Z��޷V�]�(uj��������7�y2�%ߕb�Em.�fX��E��[7X�Y<��U��*v)#��Տ6j�wW*H:��^u�Y;5��-�z�	u�FN�e�4����՝t�Gv#�me���	wt8�צ����x���9r����m��ᦷLxh�(�V?lt�� wt�:7[d
� �����A6�����s�ZI�ƭ�'��C�h�y��8�� d��	���Qؗ�o�܀�ch���.���r�B6�̘��诡⭛����B��qHe^Sd�X<�r���<i���t�[�kU�ݔ�� ��,�9F.�g�M���t]j�3m�����՜1��Esmt���j�����N�[��ˤY��U.n
2歫B��4��Tk��qq���u7]S��Gɽ1Im���(f��//+�[u�+qp��tYk��?��6e�̦��t���ƈ�Ywu�(w�?nu��bSgC�������D[�X���[5;y�b'�f�Y4�C:�@�r���D�򬤯j�
��/ �S[��H���:��m�uwu��HB�7��0f��e�[x0��9:�������
7j$K�"�/Yr��mV/�ylR\ ��k��.뒬TF�����@΢z�bӖ�phӔ�b��ס�@��\���ti�B���9�n��x�)v������u�O_3����\��d��V	%�(���-�o-0����KX��;�/k*ga}�틹ͨvn<GZ2��nbfvB�ZT�+�q��2�G�4�R���m�cG�q޾ꈛ�э�SCH�O:��b�&JH�5-9j�Ī�@(~��@
���(
"�������+�1CT_c?v�
j'ZZg?������J!���|�;����`34���rZJ
y&&���<z�����<�v#��>�̛�1��5��
�� ���iqh��������KF)"]�TSG����S���*
����)v�r�N�1P��x�?�̑P>߹���&+cT�[�)Ȧ�J�����o����F'?�������$y�sh(�H�B�i�.j�Aݩ"?C�kl���|�9~�z���ETM.�yr�%�s��cT�Q@h)4kE�t�q�ے|�jƖ!�����||om��"�AØ:��xM��F��4%Dsj�$�j"/�?a���p���0QE�DA�������U;&����1���44�[j(��o#H�N�M�O�f�����th4��4EkAZj΢�-oM����{������}��,�	�.J�}���tl+BVԀP}:#�]��_	÷���������(L�2��	2�ȓ{�������MQ����a�<	ח��"���5�������շ�`�/2�3]N��v�<T[�8��.���5*����,I8a3�����S*�c�/&�-\�eN�E��S43�M\unIv]�CKT�&�[2�A,��]�U����kk�� ;���
g��)��b*e�],����VO��ε���ju�)��&�M���{OL��}`d;#MpTS[p����T�%��n���N��o�싐�*�q���q@<)E�M��*�V0��W9/�6���bԔ6��3�A9�!c;1��9�,�e�h�RU�a�q��x�'�iP�VnF���C#�Ũ�[fk���7B���`ѻ��*xc�g��p��h��j��oLrY���h�g�vf�vqu\D�i^Kv�T��	0QV��P�w�=.�U-��Ӣ�K&��mT�諺�Y���J��A#)�c�B)��0w���g����`��|���e�A�?x�Cc��KF.��I��^i2wz!
CJ��[�����[>� �擐�����Dd�6�\|x$<k�Ւ���7��<u���М{0�/�}��BĨ�\Qs��K�}\~W]3�깿)���p�}ۖ���x/ՠ�+ʼ'���=]a�4o��!n�qd}7k7�<�:���}����mq�a�5�U��WE� KA��~s�~}�o����?�$�
L	5	0$��	Lȿ�����;�~��y�c�y�dO�t��pbN�Ƶ�2���C�˰Q^7L� gp������7uu�ż����dH��nh\{�⡭��ho����1�;��^� [���K��;���=�w�oI(p����u����� ��!��`ۥG�v����.�	�l�a6����|�_3�v�I����~<�3�N�Z�:M��S��}�'C��8/)��b�*m%�o�c�e�Ү��կ�Y�Ҩ�iĜeǙ�Ļ�6(�y��fD�2��z��N&�}n�\e���/���_��׳I�0m��"[g��n� ��80�r#�f*O��K�2�%ЖJ|@^��ΪWn��s�c���gxz�&ҪD�U�)�?���uC��g��.��ҙ��G-��v:� �%��by���hs̵�}�Lu��Oַho7�/.�!V�`Z�U6_"�Iۅ�Oށ��?&q!��i�8Ũf�P���������X��J�wP˾�f��~_wq.h�R�"����[�ķ=��&q�2��K�灆6�<��Jzƻ���������U9��m���=Зe�wK�i�)�W�1�^�	槽s��V�{����̩gI�{ܲ��sW]i���1�8����)�O�t{�����j���֚�����j��+q��+��ê�|�]v�Fr�w.r���-������Nt�mS�콈3Q�$i$C��_��e�	��`��^��[�RSt��ww�M����{����]59'ƞ�,F~i��.���?W�C��T6��\]�Xy�1���ڪSi|*Su��mJ8�Q�>�o���¨A�m�U��.��
�'����n'�_pJzu�]"{�q^&�s� [���[kQv���3�~�Ϻ��;���Uk��hR�p�#S���J�W�9Y����}��9�Ѩ]sf��LǊ���u�}�f��ؽX�$p,����ֽ�L��y:�UmszGr�q��H�k��N7�#,�h�U�w���uK͋a���y�9�k[�!Ƹ	���}q�Mp��C�rqD�k\�^b�+,��vSf���ۥ*ށ4!�h0��B��v���3'X��4c��ɪY�ċ���ٸs�Z�]������o�f�5E����;>?dG�
0��r�fV�O���i;>���o#�� M�H���cꮽ|���wr�#��AQL���L>��xl���>c%�>�raf"*5_a�3Զ�0��̋ʀ��a����?'A����YT۸y�u'ە0�S�k�i2'�Y3��*���s�̗yb�1�������tQ��Ho9W��Ho@����֪��}��<�Y��Wpj�-�|�յ���|D��
a�kgJ���r�ewG��#���.�.9�f�n�h���t��~�/���d�&&& `y��d�"m)���3�[H�3�9��E14=j���Ȅ��l�%t+U���Օ���{^������X!6>'�)�C�j��ri>�ʫk���m��d)a-��f ��l�Qȶ��M�]��ZT��nP+���j���G��<�[ ׹���40�<�z��~���Z�h.��w/|�m��M����*�'谚;���q��}�GP�>���tK-���w}���t�.u��S�U)���^7-3�HQm���0#^""�<�DVZx���_��R6�V��μE���P�h�y�:�8���p���O�iG6�����44����i�FM(78$f�WL���� /����������>.�s�7�9D��K���G2�dn:Ol}����B��#IZ�����B~\�<(�?��Q�R�{���;����� � �͍�]�(�Tsv(���N2��[��{7z�b�$L���U<{#�ޡ�Pi�K�:hhmk�gM5��6��J����13�&y
�ԋIAO��9N�^��˴����ZU�Q�t]gy���(|;��8�;��W�X���ۈ�J࿩��� Ͼ�/o����+���V�#�����ES�gn�
N[X�Q�lVg���
l�؏7��yg"�q�Aܲo6�ƔK�r'����6P��k=�b8zM������Tgiܭ�7b�q�~������$��25S-��f�)m�wa]N�{��<�}�Ϋ���Tq�G??ݶ�:L��4�@�>]��PK��<�6m����߱tj��S���,��?H���z���&GP٪ �9��:�H��=
/]�%䓋��7�{����;=�[!.
�>�6�dfW�n���m�x���j�.�:{7��R�_�O~~���̘>%��P�|���	���`l��̗�<�f�P�i0�-����3�˱L7/�ϱ�n�?��@[�������h�z]U�k�1��:�0�F'՝^�g�|�h�U�8�<b3��Bϸ}�Y����������<l���@�`U�4�*`ryP$�m�Tͧ���w�66��C����ɶ�YT=��%
���L�P�Ƈ܃6-P��&\U��~[u�*;)bk���t%�T^�a�z�t&Z�^S�-�M�Sx�`/&�����#�_����o�����mc��@�A��1�⎗ҥW��)���B����P�s��͉�cxLmQ��[���Y��|G��a��3`�����S�F,�'ݴ�s7��c1��'�`6Id�S�u�O�T���Y�ع.�oZ�M(8\��Qh�y�CÁa����n�JԵ��@ g*��U�:Ϋ/o��1t��Zb��:��Ԭ�|��w+��XڂTqv���3:�e��>��t��WBo�����33zX!�h��������ߟ~��
�C|7���4c�s߮���2i�.����f�D���sV>�=N����B�иq���#�d��/���n5�'�E�֒S�5�c&*y_.��9���:�~ʂ��#%�dy~UR����ڑ�?m~\)����t^f�#�.9�έ�=�
[O@���V@aٱͩ��Ϯ�3�4�\��Y�`��dDs4y���A��w����Х���\n��=���4(oAN2�]C�����u���r�v0yIY�E�d�m�5��Xh�v`' ������:�ܥJ�W�����د����	�SK�<2��W�����W�a����慾u`\;�5MگMk.�^�.�����'!��r�ч�<!A�+�fצ~|�j����t�*m���L����)�6H��Ѧ����)m9���)g�0آY���4c4�JO�!�u]mG�B^�����ҥ=O��j�]��L�çu�eU�(;���kL�E��U0�4�`�~vIu�;F�diL_�����wR��O:��Eڸ(nX�J�:F��)!�����{���N��B*�A<w��@zΉJ�}v��J���X7��qP�S1�M�n�{�*[N�R�J+�*��W�ځ:8$v��!��+��y��w�����W ���r��[�jm>����"C�iy��/S��`x{ �:����㹐>�4���5�=[���0�h��YcUc
jLCϻ}s�A�5Bv�zz�nDB�S9ُ0
EP0��L��	��7\Jn�1��Iͭ��U���0ӑ��)-��P���c��8ޑA�pv,�~�vYŹ�zd��J|��d�6��݋�e��(]?+�q��{��q- =��1��o�CE���Pu��M����ѐ)��:�˟�>�U���ߝ��q"�TM��D}�U���[Ǔќk��5����媭�'�u^Zޤ�L�n/�*Su��7���X���CX���gq��xM�_�:������>�����&�jP��u�%�gH��f��4��]<ħ�a�ScQp��f�iW ���|��w���[���4����]���UhЪ�Te�͈O�*;�aPXv!S�v�/6�e�ql^���n��=�{�F�>0fd��3�����+����a���`S�{�"ȖTE��<z2;���{�����"�x�yѭ?
�b�ќ���c�w�xQ��2�@�o �/�(��u`W��OTP�pk��^�]+��i=�%��@�`�����������]=f�Mc�O)%ݝ����
w��E�W��b'j�j�ω�����������\�*_u��+i�j5h�:��"��>��M~���K���D�.O�U�w�#g�r�7Ţ4���5���]��l��爾FXo��n�WlX����S#Ys0qnϥƳp�Ye��v�:"+D�by�t�y�E�[A0-�x��Vr�&Uۡ���]ô�)��t���'��� ��t����67�jX�R]�����h��I����"^��c��A�q�y�(A�"FO�M���B�'�����C�l�Y��}Eg��ϭm FA/[L �zj���	�Jh�2mt+�W��f/��T�7�~��޴�+�'�a80Z�%b?ށ�n'�ҡM�n�b�ӦZ29���x���h�ww�pk�Х:���Y��ٕ�h�l�d�$��tL>�s�ʾ�[MmٱKO(�镌0tAl�5L��b)�8�z�K����l2�5K"C�}5"�D�]�M�3��a�SZUѻ�	�rr ��(˖����q2�u{櫓G�Ղo�v�{�&�6��d^���/Y�7un�F�`�ʺ��.{�=\�_��=���Ơ��n��(׽Vz�����5�}}�@�]��*�ƓWY���_�>�6
���>bvrD]+Iƶ�N���$���б��vA}c�������z�L���dN�JTx��\(ʱԺ�A{E�Ve�Nw����+��@v��c�h`�e.�3 �}s6��x{�vfq3o�F����}p7�(iy��K*�����ȉ �]�`�w�˭̍ǎ���z��x����S��9�V�%~\�_�}��@�O����rڽ��%�l.�j�	�=�Bb��-1Y�-\4�VӻB�dL��ϻ���I|��~f���FX��g8#���&J$�V�[�*�W6�L�iW��A�A����C�J�*;΋_x�xas�RJ+kT�,��ݑ�X�lu^���0��g�lQ��~j䳿5ֆw�xg�#��I�̺n)[���Yt�
FF����#ʰ���>H���{O�O��L��\���}�;nv�Q�G*�x�f�x>���o���[�"�����f�:2����m��-��H�>Ҫr���*g_v�]�f�!��ƴ��/B�xa S���ςV�w����.��9z&�r�f�kT4S��:ݬ94j�t�)��}�eѮ9���N��F�@ծ�Ŀ��QL6|�H��BkM�#�U�s�#���y�\��-��WNÓ�DX�{/^&��wzx`d
k����o7����"������n�[o�Dl�����n�$É��ѝ+8���C����%�WPyB�����	ۛ5� ��f���+�*fv��w���)����ӵaR���xm�؛Χt3ZF���v&wi)�9���)��^SI)���a2hO<=�sv�eia,��!��{�2n"Y6�+=ٍ��E(�xb���C�v�J��~�z��\Z��t��`k@vGW��Ez{�2��˦ә����b|��u�������I�=D@f��ۜ�wfo0m33!�Ǧ�QjY������cZ~��*��x��{dU�
��c7k�\���yv_m��6u��go[��O�4.��f���1)֧��X�>��6��
�OF��/dM�@ܫ�a��5O��1�P�`����d:���:���nUV::�l��U��!q~L�IF�ZL	��)u�a������GP���B]7"y��:GN��|Q����B˳U|�,n+���s>�hE6WF;�3`iP�ь$B���޻X�h)�[W��ݹ�&��
t�T	�RXag�խ�]<��y�����A"�����W���FiC>k�T�M䞆=��q������,%�1��/P��u͔�gO���Ջk�D����0md��0�eݙ�5�!տP��21P�z��B�Le=q��w�{�͕��s�c�5�-U�r�G?gQ�=�.f����u!x\�����j��cI��<g��bx�S��P]�ٶ�v��tI��&��Z:��L���s*�KewXx+b�?#�zNDk��[&�ǎ,��>ܢ ��g{juFB�1��SP�V���6��8.��>g��[QP�.�>���B��o&��Ѹk�l���_Y�j���+h�=R����´
���:�F�\9���_
y��� �`�r��������P����s��x��i��Z���.����Dz+��;%AK
�`�����u[��u���t�0m'�ߎ͆]gz��ͧt�N�T�ޮ���Tc�k�5A�z*F�/�'o�Mg!�­56kKm���9҂��2ob;A�Q��W��m^�Os[յw�҈�;g:�or�"�f���<�>�oO.e�1�|��nM��b0n�+�m'�e�ne�(�V�m��g*�С>�i'�d��t��t�3-�\��Q�=�E7\m��t�p4Z��`{+�˳ّA��+���`;�=�Hu�Skw^2�� �so�\-3��;W>a;���:�6(!����Z>�W��t�+3�J��h������iwe����7E�s"L3P8��XSê���G��R�d��q�5�:���UKr���[��v���t��Fi8�_m��ƒ�0H�+`x�����/l^�Z�'M�IA��7?
gh�,�8��Q��J�bɴ4�B�H	FnIB���s01.7z�"$�4��n��N����5���Jp�)s�fb����U��k@9տ��|U���3%�c���]o�,V�H��>�T����,ؗ(p+�[��LR�'����K7"���A	֠b���Yװol��WI��Ms�b0�`������hS
ݘEtޮ�[�͜jI�]a�{n��Y{˰�h�D0OjWXyM��8t�cr
=קc}�r�I�Ǆuk��>��f��"wU��WJb�Wa�-����GLW���ۚ�����yY����I�^��vBT�u�d�V_2;ݜR�y��^�%�h��	�H���V��jf���)Whܥ9b���غ��9Y�Q�\K���]���T�n*A���gn�G�nؼ��1Y˫��SX���i��kvG���(a
�HS"b�w֨��*]jVU,o[�V�uqu�N
ŝjt-��Ko&m��wK���9��F��8;ܧP7�h��[�P�.���Z{�]*k8R��x*9`�S$��k�y
��Y<��[��z�m��Nk�t�-_��fƻ�k��r�8�,r�����T�t���L'mو�e̝&v�������%t���WQlT���F-mr��V��S��:\�.�}�Zb�|㢋����b����@�{�I�o�T,��Yd�L��zho��=��z��UP�|8�DY��@�j�%R��(�%b�䩶lяYv	%J.��XS���f)#�b�S�tZ_��Jh'�	E��mS%T %A�����Z����T��g��	�(����N�;����݉���}||O-m�E���v�DU0ϗ9�j/�9Ȣ����"/���DRMQ<~?�Ϗ��F�)�%`�����8UZ5EUwb9b���("�nc���9bj��������TX�󙊋��j4���T�cZ�lgQ	[f���s�
?������S�U0D:14�Pyh��"�M��,���o�D�M3��ׯ����Q��Dskkj*��Y���j�tָ�U�IQIׯ^�>:������r5D�DU�0SI<��4�MKSDU$��.Ep؝A�j?_�����d���bR"`�����#c�:���h�~�T�j����lu�r�C��ׯ���٩����&��(5������y�`�� �f	��61E���11M���Q$AUU�͒*5�gUU5{����y�8aQ�v��U|��u�����6�o	�S�:��))\�pQ�n�ά�02��)���su:VR���ˡE�bp�!%I��������t�r����>��噷�<G�����i���Htɽ"ݚ֧ۧ�74ַl���RƇ�7���d�Y}wC��#��	��X?\Y;�F�V�sΓ�<�L[r{���%�M�^�u&�w6:fB�+��1����1U!�E;�6Bu�=�ӪX����N	�1'��Ϥ�أ�Fm��T��v����ΨA� L�l�5M�y۔SzX�aS���֜�PJѻV���B�#M�B_���Xռ�A���Jn��a��f�a-}�s�2������k�v�wk�ds�Rփ>6K:��Q-T���yR:�:ki��&%��I��ݡ�E91������)�m�%ơ�jH�نF�F7���m~�)�H.Y�U*�-kd�/P�ɶ���!d������3o7V-VױG3(P�e�|ǆng)Ɵ)�e�70�F��/@�h!���s�mt��o�T����8�,�n�8T�g���ۓ~�Ɋ�8�ysaW�R퉎�?}��}�5�w�m`�r������������_���g�{�Ͱ
��TD8��"��y>��&wy%k��O��>��w����w�^��ƝJ`;|��Ř��v[Z�_���׎黍�o�]=�S��k��Y�JP�\�W����zIG�X!̽�1����t�tMf��i�S��2$�D	�(�:�2o��Ջn�;�/`^��y������v���%�4�g�X��yO"ʑ�`��h�j��F��/L���߄�[>��y���RRp���J���֥�9�z"?_�=�-]ʌ�3ل�Tu{�f��X8���}y�۵����H����6l��C�0��m'�b_�̸��ޱ��EX�	I���{]�Ľ7B۳M�;��jC�i�m�ޑ���h������*/����t�X�x0h�0ܚ����_d
�7�|�_Z�RY��UHF=Ba�=����v�dO�>�A�<�78�"3fU�aޮ��X>�J��:U_;�`����i+`�ZP8x��t>󥿛W|<�����?N���x�(]
W�xW��o���b�����������H�fM�i&m�=����8��ڔuܭ�ކ��-��p�H���"^�Fc��ێX���@�A���6�w���e���x͓�����+���Y�������������S,'ՄJh�2h��r��𦯎��s2���6����D�>S/�.���3�v'�i��U�v���󰟽��!��k|InM�j���Ub���^k�w�ܢ�����[̟|dܿGN��M��ŉ,hf`���NFXث��M+u�d�내U<7#؁35��P�����8��lϐ������E�U�_�����z<��y�,]�-��R��K2ŭ�}{feϞ�o!ޚ�L�`��Q`'�M�z�h*� >�s0�3<d���<�6�+�A�:�S,���M�U�0���`U�:���^hne��\���֚2�=-m���4��hegdHй���h�a�T�'W��э�0r<)afw��鼮E��^�O�;1DB	��$�Lx?vH�P������O�a(�s�+�Ѭb1�%�\ֳ��qU��7+_CD���e�ǔ��^1�b�Cs�;d����(��\���9�J����l[M4��Ml�̓7(T��c��G�#ŝU������]V1M�_�����)�	�����(4������ç���΂_[�!z@�*1���\>�l�����jU3z��A�h�Yӻ�N�!���'����YMXw��w� �y��$0̱���L0j��Y���1Eɷ+wC�M�6�b�m1�M2;����w�!ߺ��n�_��Oyh@�2.^ˬ��y��~�frOH��]��a���%8>@�X�;:U��VP�����y˲��A=�B�4�1d�f��[�Y�k���i���nޮY�T���;���R��zEKQb��/;���R��U9�X6?��laK��3��{�۱W�vva��>�IǺ�e]�[}�l���[��N���xx���0��}M�m���

��"���]��m�$�C��m�S�ء�ރ�������k�h|R2ZxT��V$�\߷�z�U}t��KC���.[r��[3^<<<�q�z�e����}�?Q�J�����&A�t��jG������Uǲ�VVov����_{1�2|L\�T�|9[������2e��J,�Ű�n�x�f4����=N6_�3���(�+�q|Ǔ�n�o�)��5�z�c���6{+W���H6�w��p�%�vOQ�W��&|U��ʩ1+#Eo]Q3���A��կ9v�\ү�p�J�[�Y��k�u"�jD���x�d����$wOs��V6��],8�v`-,�6w"�."�:qOs�u�=.�VA����ԢDs짘Kl#x�,}|3j�$��[^�O���i���9Imc��l�9 >�%��Y�B�"П�Оo��G�>��:�֊T(���B'�I��s9�x���p�3�J|�(IM��K�����A��Х�v�%Z�OXf��%��4�7{(�]�����Uvke��lk9��YP��p�0:u6z3�7X�.��M�?���z=W\H���	�_��`gw�<oI��u�8gfqL"�e������|ܣօd����+ܫ�9ݼx�Ce���ѱ�DVmM�Ǯ:gۧ���u4�@�'��VO{5�s�tڻN�;�۱�+�i�vBXf�@|1ۥe�<��O��Y�5��I�F7�ͼ�}�㞵a�hmP�+���-���\����OU�������5ä`�S��9�2�}ð�6��ͅ�OͨT���-��˾޶��c.9�8ٟ5��B���d��[�xVg�7�chWO���N�gOv�@HF���,ڊ� ���rڬJ�c��S�ϧ��SQ3���f뷚���[62�yMl�z�_���M���Hd��p�o�3@*�5�Wf�'X��I<�\�ެ;����d[>�Ȏ�=X����	�ܲ����d�v��{�o�I�ت�m�r��|�@CaR�5>3�Gn�hvg瑏~Y܊��ޕ�/O)�m�jUa�|�/6�	DB�	�ۦlѬ�|�3EÎ1��4s6/7���u�a]������!�t���i
WǛ����v�.A\\��9m�����i� C/���:��]�I:=z�n�r�4�ǝ�gI��G�����<>��j1q+�՟P��H��!���W�+D_u��MgAB��CYc��_����*�n��FG���8ޛ^Ww<��}W�st���K������.+"3������f���{?,��[��W���A����P�����L:��=}1"(�ma�:�3���<l���rQ8B�tH~�k���k��c�D�TY$��V�{Ʌ�׷XI��
��N�-E J��=�1^����]Q{槌ά���,]H�׳�R����+�ӛ��g#5��S�v�S��D��R���r�v n���"����SG���DB�L_uE/l�g�����ܘ��:���q����:��5����[`]���"V{�m�OEu�ԓ�հ�9�U�#͌`���5����>��	�<�*2^����wr&R��L���t�ݸ'��cA�mù��^��|��S�!�0�n�J��&k��z+/X!����Uu������uh���&���mh�*�:�ujW0���_)S?~C���*բ�1@*ܜB��eb4�H�7�����챖�u�M�ǲN+��\�-�ġ�Z�}\p���}_}q/t��f�ys�fŨ�g��8�7x���:D�=��>V/O�+i�9w;���h!��0]��~U�6n��U3��1C�>��h���9�/e��ys�Ҍ�e�.�C���q���W}=�"�z� �y󑙗��6�v"�o���J��2�[@O�#����q��S>{�����-��&��Y�m�ydoM�'�w$b�zo���<�@>��1N쩞�8�Uu�x��گ��Iv���M�X
�����A�ڈ���r�c0��eY���c=����x��&#<n�F�mCh�7O�V��Wq�M��5 ��7��ە��;j]!��W��b�%�s2�&{ŋ��n5�,�9:�*8�q.�c���r�V��r���]�ʮ��������>sQ�^����ok��Zzb�	��s�F�N�����8!��ev\f�Mu݃�dv�6^�����9\�a�s�z3Ϲ�����h/�hs��pu���J�b�&�)x�9�9����nu�kq�u|tYk���pCf�t]qjH���*p�a�^wn�ⷎ����iEwY�D�n�B����{޲I�v��:dƣȕ��+|� m=�ǜ��@}�>�Ժ�,�5M������݂cu�LwI���W�k��v8�~�_�b���KI/��/�I�ޝ��쒬
w���z����[���O`}��xrK{������J~�X������\���P�-8X����f?�n�x�O�R�>Q~���d��]�s���t��Dk��vLʺ��Q���1��b�_��i�Wu*qT��_;Ы�q#��[>/�-��T�hq-e�gB�سѹ�k�]u���R���Y�O2�Jݠr�S������,7Y2]�M8�'�/l��}�g�xO�h�Z6�	���T�`�X
^��T�Vp4}��[ty��b�BN��~�S� �y`SU ��.�̋T��Uk	��}�LKM�e��b[v@g3 r1kz@�og�P�Kid��,U�W��I��fg�!{��<�`L�C�,����yWYܸ�	�mtd������;"ƴ;��ژw�m-޺Mm�݊�D���BU��H*���h�F��������;�R�ԯX9�vNZ򓜯ۨ�{j�B�n6R���� {t��㳪����`���W��o�ֽݗ����ww������>�[�\_]�螄��~IOU]��;�L�X�����u��?T�m*[䃻2��Uː��W¯��C��/��7I�C�t�I��ӓ+{�أ�kT�]t��ާ�5���ޑp�s��n\r�no��CO1���ٷ��6��!#���zc��,��:瞋����d�gVi�{S�� =Zǣ�_���X��^�:\3�z<���[
�i�c������� "�Ȉ���X�war�̈��6��@8Տ�q����cufV��gL�7��y֏6;0W��i�(�VJ���i0Md�����w
%�LEr�&:(�l�n0e!�sO�'p���ż�s1-�,׳�o{�Nkt��a���ж�j������f�2Qe��X �X�XfBf�������ݮ�o^�j����6r��W�a�O��[��� �z����F�T~��Aa}q�r.>Ux�h{��)l�<{i�)�ʧNc�
���@�_My�hUxUK��K�u/,U�Ω��)�.�&����䷋�N�uƖ2�H�»�wV+�U�`��z�x��	������w)�W9X
�U�"C��ˆ�-b
�zYX����Hx�^S�e���j�֞j}�磲"i]�`��7^F+B�JoNV�f�r�G�os�\k�3�ӸDSkV�\t�L,��O�}M $�E��@��;��K��]es��=ѓL�}�{�T�U��t�?M"���Obxu\�U��&�y�:�םG��o7~��Ss�}T2\�}2!�,7�qK@�����=�Q�4|z}'3��%l�U�C��O�к
�r�2��l�jf��N��M����$I�iܟ6��+��]�4��f���Os���v>���cw��lڌ���Od�iG�O/+in�N*�<��Ҳ�� ��n���|��7�8�>vGz}GiW���@��SC�j�)�2V�Lق���՗em�r�GݍN�h�t��Әw(����*�-�1 �:#�<��E��}F����ׯ�X�q[��[q��4�����Y��P�/7Z��,�`�X�M��Y�+��m�E��uu`�V]��N�1���k�bS���p°���n�;�*tq������Z��`F�ZJ�����@$h�s�m�P��ii9wa�6�F�F������"�ܚ8�땣�V���ϸ:��4�z�s�kz�����N��YO�_s�3�o�Z����F�kgp�t*��u�o�~;N���}�2Ͳ_S��u�h�i%GnV�*
!�\W{�8��r���s\#wՖ����&2s�ţ-�X<��c�.ą��Nm�yف�{�_khP�>�gh��]O2���>��X�]uw�B7)�(X�I:��K��L��%������nl\�q�y)�8Ⱦ���q��<s�� �5�=��UG�*Eb7L<'J�:,�b���2�S�']jmmN����(oM/�m�Um|�)P���'vȳ��a���@�kq�mݥ�:�������4�͗;b�Q�����"�
x�qއ]�nu����S) W���j��5G����2���!"��9u�AB�v����*d5�<nh[�.�,{�r>`��ݥ�m�h͌�}gL�7L�&�3�h�
I
=`8X)*�u���b���wk7��&Ǌ���5��@���s3��[�B��YL0S��7�������M���䒮����|6�N���������JXe��_d,e&���Û�&ݑ/7������,m��w�c*T���8�I��4�=XULÝX@C�����v��vWSٝE�X�*{���ְQ�כ�(n�eJ���YU�)1�YJ͔ޜ�F�q�#�K5t��KH���u�|�뻵���M�d��lŘ���N��e��4@v�<s{�n^:������ͦ��o�f�&,���2K�����X֮���r���fɽxJ�E��v ��t��yw��U�iˊ%�m�]κ�8�_l��ɧ7:�:dp��]��w:����X؃R΋TY���K���޴���7�j�q�)����/ALǀqu.�0�X�'V��Z~�K��f9X�t*�Y�_ɭ�J�_��j�#��0J�k��b��V�+��fwM��V���Gs��Y�#��� T�M�]׹��[���<m2��[��Z��<���$�ו�]�J}��5��,�6�lJy+:�ty�q�l"�X�^nA�RQ������w5tq��Y�^�u��6g&�.���S�ُ��.Q꼷�B���%Ohh���܆,B�ܽ�6�Xg*F�>����5W	2�u:EP�����u��#f�QBP�<,oV�m	�sU�.z1��^i�oB��pr��z���53����o���G�Yޤ �}�NX�RHaq�)TP�M]��:1��71�a��lST����������_
��m��~�3E���홈�ъ-*�*�!�����j9��=z��MD�F�D�QATDD�Dl"
*Jc��NMQ�h�z������h�QTA�QV�{s�����������b�j#Z���$��?�*��cmlh��cb4��9��1�14h1DEEm���cZ-���T~?�����ڱUT�w�xQ�6
1�c�9ڊ���Z�����ڲ�[D���������h�ӱ��h�+C�Z+�AST�����l�q���?�Ϗ���H_��5��-QUT��٪;�Nf�6Ʃ���ш+c�<�������(򿶖�[FLK�������LKT�����h�[nlA����E4[�F*k_g�Ss&7�h)*���g�t�-���A��aدY/�L�5ٵy8p��W`|o�';�o.ރ��rOk����й�m��A��clLX����}�.�"t��n��d>������Q}��n�X��=�l�J�{��+���Q��	��f����o��{����1;{�ܹ�`�9O��nw��v��1ov<������[L�Y)R�:�!��^��묞>���X����#��vWs��������Z-\d[#�������fe��	�F�>�FlX�a�8�s�i/ܩ ״��K���su�yok��M�@��d��� y�u�k��&5!�{�[Z�
�q���z��GS�z �a�ֱ�eb�<��)�R)Y��΁cK(l/��\M�99.0t%#`�f��aخb&���=r��!�jW�7[P�q�va�����f�å^�RnP�Ԯ� �n��-�]����a�Ց�˳��m���2��};�ܩ	 k�J�&�ܪ�x¼����V���w�N#��zᖆ�+F,FriK����I�U��j�u����� 3�������.�G�{��?(j(��,*�yT��)��\gM�ėk�7].�y�QڕaҢ�m���!k���3y��`��:l�ɞ����06�����q��U����z���F��]^��
 vz�.�r5W��/cu�u����Wj�Գ����l��=޶��Ii�����<���Ǫ�}� N���;�ЩL�]�]�9����ar)�4J ���F�s[���X�nS�J��P���a�0�*�n�wo�srw(��Y�:a�}��Bީ��x̋)���ķv��wL4M�t��*�]�/Λ�HEΠ6C�p�m��D�>ƍ�=�Mֽ��S&=���\�Yٮ��yL[��:��;א���A�RQ��_��.�f�u���kn���ȣ��ӝ���t_F�vP��i&����9�b���=+a�^�׋9�����cC�[1/�����o1�~��!��.vŎ1����H��"�Qj���̩�f��<&��d�v�g.�kƋ�4�v�G�C_g����C���{ƿ5����V�He�
q�#3TfT����K{��C�o�|���D�P�K��K<\�T����B�y�_�豗f�Z�MZ����I�̇qZ����>��pfM�)\B%�W�L���c��3\�c3Uӡ��w�z�?E��t=N�l�(i�1�Yș�]@ *4�d�i}��H���n����_��[t
_�lm4H��^�Y!+v�T�@����.��?ԯ�Fi"��m�K���9�
Q���_kPO^P���R˕;��v���w�`/������Tk�;��3�5U��yH�>�����!f��PEeVKU�dU���b�H�&�[^��i��ˏ6�12�E-��W�Y�|�&�4�9�椤��*o���Ů6��c���*�9M��p%_8����	�
��ܵ���n���n2�I�1 ��0ko?�����-�!�(�QA�v�D`�}�:!�G��$�j˖�>b��/+v�X��2:�?�w_Hi�D��q�ۼ�V2\�I��w:0=Iì�k�wJ�~.W+nܔ�K��l��[��U�&��bb��a}���/M�3��(�.����rT����~V����j���!O�[-��Omy���VyH�f!u��}T;�09�[�[��s��]{���fvt���t�?m�])����w:1->������]7��^��㟕m���Ax��:�����~4��
��vf[��-����ojT�[���h����uL#z�S����]�w�;sx��r��ɲ�s��^��zro#��kg(g�c�h�!�$��ҟ#L�hU�'Vg"Gk�mg�%g4����ì�-��w�����.O8�n��q>�;�h/��^��_ec�����?���s�� �0�]�<F����/����~e�u���mU�e�5�Z	��nV�Ci���Yv#j�x8jw�g�]gu���]�&�:������5y�� �+�5u2�U�u�j6��^R\�SǛq��ɉ�UvzE`z&�!xyNV�fU]U#3��i�~,;�y;��������Ώؿ�?��Ʃ�jj���n�!aVkwgl�NٞW�ǹ��[��J����©�k� �A Tv2�~��m��h�����nJ޴��bݥW4i�[.��{Vr\�E�bhҔ!��:z��k/y�oH����`M٢�7��U��*���1w��g�?)=#}{��s9��O��ǭ9���A��]hw[�wC7w	/��m�t
�����˹�K���N����G,?.�I{E}�Q�gE�]�vEP�
+	�]�ͮ����m
�C��{�ΦyV�W�]�%� ��qWI#�d��ϗ	Ճ}3���R���ݳ���Zen�Z�Vok��^o�/F�;O�mT�z����:�9�Q��.���ԧ��/+h����פˬ/B%�c2;;ڻl�[sD��R�� W�ޡ��+�/��Z��y@�����kq�N��xu�ϦR�V����w��_Y����ъhïr�Y���^��ge�ٍ��w��t���BvH̀���<���z5O�ur�F����;��!-+��.�]!u�r����}v���>K ����t<��0}����׹2�W��̑�˨�ĵ�fPm��u��s��i�v=��8Ւ]7�t��խO��w��N��������d�� �1��rf᚞M�y5)�vqֳ��*M���6/�1�a; s���cy���u�9O�]��	�W^|�t6�9��kf�6n������\~?=��a<�[�Gn�
j}�i���ث	�i
sڲoN�ЀL�����)H��bL�]_k�j:�W����~�P���ʯU4�������p]�����	�)p�@r�u���[:��R�8��mbInc�����U`�8����W���\�-�u#hz���S]����D�/T��L�%�o9X�8�Bu�k8�~L�Q�5���.��6Z���z�~+�M�MR��TH糷H��T�Bj�o3K���槱�M�����M0�n�+�EU������nY9'�����A�o�u��<�YP�&�5j���J��=QX��S�gn��!����Q���l�|5.�X9��~*�u�Xͦ��{LC<�n�s%胚sb�+�kFm��8(֫P/��j]>mo�����"���p��g�Kܓ�JR��E�r�g��i�'N������~s�e�C���u�~� ����nw�D,.����u�����[,ܥgy�&O��N�.��U��]:�Brv��:��季�<#�	���=�����&"�گ�JF��F�u�B���	y�q{�SO��lӦ��"���w�-��a����㭛��!�9��]Y�Xz"�e���9��Sop)�++v�q���+��?� �4��G��/N���U��Uۋ��|�-�mB��)Ɏ�.���ϒ5��F]e��[���.z���{Bv��$MD;����f�!j�
�Qm��������ً�<�xl�C3��T��P�}"�e�{��)��u�c�6I�������Q7�qa̻�~LḌ��a`?��1���n�U��ӛY�ч\�͡��i��x���#��1�z$����%ߧ+�����˕b諸ȼx��9:������ou���C����ݶcG\��+*���g}�w�YS#���S��{z!j�Ō�$qC;�f7�V���W�K2����s=@מ�T���(�U*�nEa����S.T�~��gՇ�/�=�y�;�#x�?��g�ڱ��t����iuY1����]x�&x���p�gٞ����~A��n���M�?0t��g����vk:��s6<��{�ၘUS���ͪ�o�[-���\���~��#WsJyb��,��z�;��ӽ�p��������mzC�n��!lnzX'���?�9/]�@	�){wȬ��BwA�� �򩴲��Ҭ����qe?i�"�ȬT�����7k$���f����9u�U�ZF�����h��w9�+:�w�+�ZU���:'r���	[6*�� 
|��5Y|Z�@Gm�j�KB��Y9�Ț1>[}!��j�h7:�n#�v��9��"RɁ����w����"ݝ���^cӭ��+�]ߪ�<`��B���oC�H��*v����t�����q��-
��TB�p�����ڍwU�����=D_+��#�Q���;��Q�u Qݳ�8���J�3+sr�a�]N������ƻ �Q0y.����C�Jù/��D�S��ߢm{�JM��;�t��q��/>lLu��R}�AZ�P�R�Kl����� Ea���6�71���L�02��0�y�dIޯ����R�l����)�M���]������k�!<2��M9jf�l�5P�:�[Gz�	��y��M��3�v�z�t�IjUw�A6ʳp�q��3��ӓ���;P���ϊ���,�&���y�<�/ �q^a�ݞT���|:���Ю��5c��<jDI�Q��ۃ*�0�]Y6��M�r�����kN��N�#Fm5�=I~���f�����T8qc\��Xj������f*c��L�%�{�a�p����]�����0ְ+��7�`[:r���W��k��p@��vɓ{On�z�a�%�@nU!���L��J�񱱆�L��q��Rg=���������q��~��+�-��?nLj�s+|�=U{����7D�p�9��]�s7�i���u>�df�RϡX;�p�.�g+��ҟ��HeG�ױ��M�%$od�]�򧺶1�u��	��̎�<���߽��5�)��r������m�UۯK���J�*7�����4:m�1���2�F�5��U���.��(�a֑� .�	���j��lȸ� ��oV��ˋ��^��g�t̲��oVhzFc��P�Z��0���3��z�s0��S��@:��a.���]^���g�Q7�'Q�����"��d�m㘯�Z���|y���u�f�d3�)щ�����;ݓ'�x>�Eg�Y)zoM(n챼����Án"���J���`$ۛ�)���8�e��+._(�����4c=��_.�ٮ�G�@6�mc9{S���jʺ맏�v�vK�$Ju��s�N�LnR���c�үo�)M�U:s=}ĳ�z��[��^sڏ[
�����je�O4f����ox{\�l�ϮT?o�u􀬜�:�������Z�V]XT��������3z�pmPR73��)�^�F�����!MnM�`�a�CV�7�Z87S3;l����Vؙ9zg�TE��t�+�RON�.�z�����$Xޒ��v�M�M�:`{���W��mW�n�\�;N������W����Ûs-�(�1}^ሑ~�]n)S��l3�o@P��@��UkW�U��OY��{�s���^:�sz~KkĬoV� �Z�2Uk�ݪ���2��U�SH6����G`e^�Z��o8�Mn g�rV�Œ%��ޖ�1��,��.�ٖ�{�9ZY^Ht�IzXg_���KliT���q���6X4�̣{e]�l����ws�]�q WT8L����{x�W��ӉXJ���������-���ɨ��}�^��ȺSC�YZ���K�ǀ��tf��OQl��ҷ�l����a�Z��i�\�v!]nNĦi`eju[x��v��N��O������N�O�H�n�����6�J�wY;1Νsf�]��+z�$�s1l���<�;�t��01���"�:���F;^v�u����IF=����fmP�URpYe��6�
��F%��*&��u���;+���D�J����r��3�� ��h>�;`B��+pӐ���������{��3���=<�9;X�k��M��������f�p�a���A{Ve����l���!��;�*�E��6���>h��M���0Z��v��)�!/�UgH]�V8��*�E��@n4V�s_b��R&��{�K ����&��/��H2�,���>3;w%!jf���,������<�Y��rC�q��|�����i�C�ɹ�6�p��w�w�n�5e���?rQ�#}Cm� �S�_ZpVBu��
c�o&�+�Pde\����w7�ãæ)��Β̶LZ�i�gB��Reӽ|%ʙJ��v�"	�ɥ���کXz�R�o����U�p|���Fq�hq�}��[���\��nX��~���vj�72.J?ӥ�1��e��gG<�n!����Xj����1h�nqYӃA�Y�[*�[��R]�'����ͮ�M�u�6��{[�����]���צ��k��IoM�B�(*m�������6��z.S
�����V��`��D۬���i,�<�.J��2�Mg*�:&�P��%r4�f����&�F�db��/M4���R��!OHK��)u\���#��(T�S�˦f�����M^8웑�]���sBM�,"�'s�H�yT�AJ���f�_���*������ͤ$�ێ�v���0��cˡ�)��;v!���fw0bhͱ8���c�-�Ǻ���DU��>�W�-B�u$2>���.�є�\� �=��;�e.���YX��f ��vTW_^u'�k� khꮑTU�$.�+�l����Zp<Jt'_`�Q��.�"ua��.	Գ�IHɗG!m͓2�us&��"��(5�(*�]�f�kz�
�\�V�*Z��e�����]t��gAl}4������U>�����w>����c2X5�dN�Op^;Mr8���u��
�o�ݍ�V�R�u��X[�a��=�kMk�Z��Vޠ���ƕ���� ��C�6d��i���umv��R�ƭ9O[����@eAt?CK��5��r����8�ZE��E���㦭+�g_~H���m�9:V��"���;�XTw��mt�$�I�0��n��/�����e�?���������#6���FA%b��X�N>m���@m��*�S})�u' _t��y�UM�)�n�Kh�i*P�f�G��9qKC5��o�;����B�/4�TQ�� v�Wv���P2�h*�nN�V����nU�r�+A���8h�"�r�J�� IP�qڤ�e2�]��1PX8I=,S�-��@~�¿��5�*'Mj��l�m�o'�P��-�x����>墪���~��4�U��]r+AF�&փHU;�9��i�:��>����� �i(k�l4b��CG64�M�(m����NګA�E?��������Ȫm��"ѱ��B��UN�V��QF?\�hĚ��g������("=�(?NƢ�T�z.�r��t�g���l֍2E�k�Z��1&ϯ�����D^}�9��Q��1:��o��nG*�V�;b�
v�	�[PD���ׯ���1��`�R��63��o6���ŷ-�U���9G�mN�ճ?_�����y�j,cb����U�g�6��PD֐��ZEh�h7��o�������|6)�1:kZ6�lִh��T����֊��h��t:h�m�HPК�b���m��1cF�j"
�9�*� �h��ꂪ��(���jV*�*t)��]f���<��M<So{����\����n�5r�%�D�qt�]tG�T	Ƨ^�ῖ�Z0��o��3���7@b�
!C���P�KT� �����W�M4ރ?��د���IgT"秙�Q�u�6)˽�E�rl�n���}���iu=����\����s�����8}��R����={:�Y��=.{�qf�_�;(��!J+��g�2غu�M��&d��V�j�s�ݺ5��VL�\gM6�s׎��N�-M����:"Tݛ���oMU��2�#S�k�+w$k�9~'�}Gq�;�%9��ͬ<��Tg��[���uN��a�]�����ӽ��b,?����[7_��,g��ι>t:P�h�p�vL�Ȭj}��,ה��-�[[��6��j�r֞�F*�2���Ό�WJ�=��[��$�����9o���N���ܐ2K,�Sz٣�:��6)x�P�X�ɛo�����E����4qc�s�y~[��#U2J�z�R�>�>\V)��/6�4�gL�)�/e�n95`y�H8�M�|O��:L��4�g[י����<j;��7�w�V��4  h P�}�
S��wX�.�	�y�����m�G��Y����wQ���s���Dw=�౔�@v�M�]�<6w5�pd x�9�X�kV �P;����U�*����aiU�<<:���l�3�Lf捈��N���$c�K+��e�;չj���uE���d��h�g{'���f<A�u@%yE�F�n���7>��!6������ˌ�Ri4,ܦ�[��޺v3��gq�D	�n��+�d׎�Iv
؅��}3+�+�z����鷀��p=�s(I ��������Vd�[�޷��,f�˨z�ێ՝����ϞX`�^�Ue�W(�����Ox���s���B�]W/'j��� Dy`��!�ϡq�\lR���U��bA�Q�P+��z�jgYUf`�^md���n�[3�����7��3:�̍����M� h����U��M1־J���v�l����C���A��T2;<�n���:m�s��I�`t�{#0�%eZ�v�8�љM�����y�?�ش`N�C6�x�ߩ-��a.�P�(��/�����y�Z4�??ng )a�c�л�C:��#��܄����Y�c'w�c+~�+��o$��Z��S;�Y�w;����Yٰ�绑�z�M�T��b1%kt�ι-M��E���T���"��4CN�i���4�����fV�ud��{7���!�28ay������J FQQƟn�M���\�٥qۮD���0+`P��V7Nmv��}�Te�-�v����jV��6t˾�1���6z�dǨ6^�j��������b���wv2�tY���Me�����I���� Yg�%�jC&8��x,�����5;�z�x��44��֥�@b�C٩�t�mx$��I��Ӑ�械G]�x��L�_�ڪ���]祺=���b8�i �׶5��a�_(�팮!�Κ��j��%*Y� WU�8�E�.��ڼ�:PJ�W?^vf�Q^K���޾u�5e�H�:�j�r��������|��r���'0�p���{n�_��p`+�@�v[c�{L��%��Xw�����W+�%��'��"��jxEmz3�b-?���K;��׾S�ri��=���v�]�b6C��@���b�x�NgVf�s��.�Qypգ����f_�=�����,���J�R�9]���ӓ7�Oq���]�v�����d귆�A}��c����o���u�4�My�)݃.���/,j11�vP�~���g��'ѫ{�#�z_G'�m�5\ѷՃ��f$%ɗu����`�2Α��u����1�]�x��]��FN�@�g���a�����G,����\�o@�縰:l�<��+W�#f�8�u����A�PyV����?{*Ȩi&!�k�غ ���n�D�ɽ�Z��'�6ȸ��-x��>�����L��}K]��[r%X��bѳ6�6�M\�S6&V�	f�<�ثm��<��@��
+N���MM�X���Qɶ�F�_2��=X´Z����
� mx�����H�;u�KE��\���{Se�d�ǟ]���^����5^���y^�k��RV�����b7t3xl�r�ݠQ�S����R��SL�]�=Օי&��uۮ�:�tĠ�w��\�l�������Eg#�����=ۓ]"����c n�[�� u��}앙�#8�]��N��oƯ�bOu�̍�ʤߦ�~��.���^��^�߸�AE^�^��J���.���)cٝ*�=�\7uf���䂔��d0Œ��-�VH�{���Jh��u�{��X�@�F�k)�!n��!����_��un�jĆ���΃���_BuR�(x����;���.dZ�u�O����?C84v�U��q���!�]�W���v��U��hK�B�q]�4S��E�z����u�/	i��x�$dsW��Ի}����+tg��V��G9�b;D>N5�{�މ��Sr�IL�+�Wtx_sa�E�7�e�^T��bl��Nuy8�.�IgW���\�Ӱe��,wa�b.g�7{c"��:�S��a�D�O�GeW����WÖ_�\eAn�}�{bs�k�J�S�Df�
=F!�Ɇ��O�U��c)�7	��ٵL�OQ�yb�"""䬢g7���{����g[:4v��ٰ��`���Mf���+�w瘪護y\��`�n@B�s��~g��5�na��Vߒ����Pw�]p�r��գ��9�D�e~�c���yљ����#P܋����]�ؐ���3�]yg;�k7\u�R��n�f�tcx��m��:��U���x������B�zEtUH����z��j��j��ȩJ��;X/Z`P��j۔>�������p�X++Ws��ʅ6��ԣ2^���tp����w1�ZC}֚'�A���?Xc#��%���U���S�ym�!��Y��� L���`�G(��
�!�2���/|�&y߬�6E "2�͎+%��ϭ(�g�Zy!�=̢|��7'�V8R�������n��p��SvDK�\�����ޑ�^Jٽ�RЭ@9���0��nWV�Z��{%�Ϟ��������O(�~J��hq������2�-����cwy���r���w�LzZ��7D�R��:>�m[��^�ZR���u$E�U�س}����W�E[��e���1}5r�4W
�QDEûl+�w��j﹚m,�O	r�K�����Y��9^D��m��q3TH�M�t���DY�(��$6.D�,�+WVG��Gq���N���´��8�!�t���L�fbP�]l5�07eo_9H���p'bbwy�b��c��m�K�!k# �o:�E�� �k7��C�*�z<��m9{Լݶ�B�y�Y3�qC�� 0ED~����:@4ެ�`�LU�}ٰ���b*.�+��|/�=���A}�-쏵�QwvR��@��n��T�nW:�f=��P���׬�3���]��N��Զr�C��!�o��{h��s>���pV��4�ހj[۷�{��{|�����k����{Gȼu���� Fә���Se⊭]Z+���qZ=�r}���sSp�9�I$�JȽ��t�����]e�g����M�YB�/?<m�M�8����6��}R���'���i�~y5�M��0a��Pqa����rO]oi�h���j���]�)�߃<*y�8wu9"�R�^�˘b�t
F�����K�`Z�؁�\q�L�͈�3n�,����y�����QX��6v���M9}�j#d���.�[�����K��<��m�s�W�~�7�XN.�]t.Ϻr�l���\ʝ��l�9�gZ3DaS�m�8����b�|�&c�co�{�M8T��{���"v(G�57XmUX�+����E�~�3�����٩�\�9�c�����WI����z���:|���M_]J�m�u.�e<a�6�c��X�κ���^��I�Ε�m͓�f�	u���ᮥ������������r��}�Ř����d���è�2�/�׼*{{7M��lկ����6�{�Z̟wOf�]2�w�W�̻�@�{KZ4ڽ�T�'�^�F�%��"od��]�Nuh3�����Ͽl}3�.�0�w�e��O��l�N�+�G�v�lr�4���V�7i�؇
xa;�5W����,���Ɋ�T$u�-�[y0�[9,��.n�f$8�c55��n���<Mǔ���Q�V�� ��_3"�h�qU;}�7n*����p�Y�u,��Z�2�.]�Y�!�<�o˭�f�f�S����w"ĪB���#�x�}�v�G�!;$g@jx��[y���$�/X՚��c��֓`d��{պ��A0-r.Щ�v��W��߸#7X�T�3:�ز�'�!�r�};�)*��R��u�������*_-_e��͐i�7M�����o{NHX�����k�z�5�	�}m6��gv�2�A����(�Q��%Ob"�q��n�G�Y���{v��.�D����}�]L�YOy�8p��x�X*q"���u@�k��+�Zɜ����4޳.����%^���.t������;��o-돞$ƈ�m̫������@P�)2�(^6�n�z����wf`�h!ʸt��v�ݖļ����ߺ_1���t���b�󳩧WgOc�o8�i�6�@�l�̻	�}�!1-��V�C4V�W��wz#��Z�8��	k���瑦�H�m22N����������6>UF�c���� ������4����R�`��v�1��/�3%#{�q&���f�B��������� �,�%Ʈ���+�8��m�K>�y�*$��޷ޫIEa���]	e�!5�#��g��� ӗs|7y�"��i 8����̳a��T���z���=)�ik��}ms����.o5%��8��*����Q�o�Y"�^�Bǡ+�sF��ڙ��k�LD�m��7vm�6�� ��PK���u4��[z�'�TM�^��Cg�3�w�ݗ�2 �o�N+��(~:9�A�\e���g���P��l�`��u�t�3��2�יL:y=FU��uol�������cz���.�''�ƺ�~뷞!�׌�̰y?�~2�vL�����ՌԻ2�ȻჇ3�уk1P=�Y��Xk��9��I����}����N��v��՟���vsroOP�xK����.�T��N��V�S��UV���z�����'�:k���]�l�H��Y3��+_J��eU>.����3'KS�R��/K^GMl/P�ɱ�X1��qÖ33D�dOa�A�F0W��Ȝ��v��E��6-i�k^3���qa���2��[�Zr��J_m�7O\n7Oi��6��޾z�L�H�ca��@dW$�?[��r�o��[hhJ�n+�m�x;\FQ�i�l5�xŭ�`|��l�oޛ�,�D;w/R�EK��%��n�-��rCh��e[�)ta�Z�Z.�6���ƍ����c�H�^��Ww�Ȭ!<�C8Ϣ����8Z��^�>y�=�)bw�?y��F�19�^��K���hq�X�V�����(�gV�6�;#	ʡx�x��c��<�Q�~�\�Z� h�F(��mr������^Z�%��f����N����6;�s����2��M(�c�`$5E-)��gb���^!V�� �˿�o�eۇE������#�ي�.�B�ؼq�[�nK�������;]w�rWR=�F,�\w!O�QwyX*A��^6���P-�[�q�W~�˛ф'=�F�øB�8M�*�R����Q�g-p�U��i�+�k�Q�l��Z�=������;-���W+�a�S{��:�dz����+��vt
y�rRX����������B��s6����,_Aʘ�j�;�G��������V�	pn�U�95\gS��:��{���F�k�qK�[5u��2��N�����1�n꧵��tw�ԕ��&��� ��slV�y�2U����v��=�|(�[ץLO��aM]����W�ے���S��U��p�l�@��m]1�\��ԟ>�˼ӵ�:�����i��h�t���TX�����sg]w>�[	4�'�K�� E87��_$�6�L�܌κc�Y����ގ���A=T�Y����y]�����}�G����L!;�Ef��o8Vc[Ճ2��v��rM�D�Z�z���tmǪ^ы)c�ܨ˕��d���n�������9���gn*�V�����Nv�+r,Og:��Z��'+�;�^�;��:��w���;�s��>��MQI%})Jb�)���ۚM A��е�ϧ���c��e�>͞;,۞��W�Z��7q�;GmvR�����S�'R�]1�vJW�^�f��%��۵�.�<���<��̂��W*.:�A8$gi�S�_����O�q��᳘_u�R����]�O��5��s&Ⳕ!�٬wt��`�[�lr(�o����D����|��1o"�}6u��]��yV��&��7�G��1}��лF�
㝈=K�����[�8&k�4��y2RyR�Sx��5K9���ZcJKm�b�#�0OVF&�&֫Ɲ�݇�Gd'��q��)e��)��W&;�+sF��7g>]��J��Zz������:��[��T����t�_���ĚѧM�9�k������ӬS0��7�kX�4TQ����c�)L���Y�r��N�O"��5gK.�	�Vb(�X�R�j�'Ksfq|mb)wt��P���:��m����M8^DA��LiV'H�ꤰ������s{���%��s23�a��*�V���I��X��	��;u�S3Y�J�ra��g�3ΌwF4�o9�S�i�C}�ҳ�V��c�C�Y�w��]m�S(!y1M.��D�����:�zu^�4&~n�nJ�}+���V�>���-�V@����󫉡��[Z��TF�W�xy���*���Q��Il�5�t���V�����.c?�r��V3E��~?_��(��h<�F�����s��*󜹠�H�&��N�:�s�$���ׯ��/�C�{p�4�4m��Q�Ѡ��ڊf�[c�\4V���Bg�����<���4�STh��F#m��5F�+��tV���A?���������k�Zճ���E�g:�kRRlmZ�&�װr�9ƀ��
5�1L��ׯ���:\���v�ֹb��X�%��{i劒&�����O�������"
t��T��Ʈk"��TDci��F�#0SN�'�5�����<����M�����j��Ɵo��[}�J8A��cAEi-�5�gF	ϯ�����%>m�6�.`�TLTl[AE��m�����^��9�-j��5PF&�w9�+c4�a�5������4�0��"��
�\����(�Ϗ5�7 �o���)���sҮ���(d���^�w���8n
wʺf�x��[I�f��H`����I���Św�]�ۻ�'{�Tg
��V��|���c�����
#�u,�۾ۮ�xF���9Ҳ��4j�j����/|�ڹ��"�V�$w�Ƥ����V;�&��ݲ��|�����p����nM�)��3i�;ۯpF��Q]�|�����QG���n��tJ�_;����@����#"|�U>c�a�L.2.6%3Z��=t�9��U��@�{���k5�s0���g�as���~7��[���'���L���ј�#;/xN�9�������ǣ�r�@w�cϞ�X���Gj(F�i��[�WvL\��zx���Z�yv	���w�ǜk��|=�Iժx[��g9֭���i%CWf���07��3FC�0΢�gQ� ���3x��b�_�����	���B��;��9��撬��|*�| ��s�^6 �ٶ�#q���1��o�z�]��/�V|��C	��J_E`f��nJ�zj����-뺻*�m"�S��}e#�v�<;�������z��܋\^���\�RN�i����ڬ�o�,�s��\���=w����~�l6kN�e�Yx�W(wv�3{'��
L��uf�`���ʽ͖�n�v�tЁ�M��M�|��=��]U��!q�������/}gv�wy�&�d�΃f�m#U�r��e����GLL�`ˌF��u�:H؆�О�>�\��{U�=3�m�5T��}6�t7Y�̮Mڠ	 glU�ϽNnFG�&��G��*��3��n�B,M��3w31�e�!�A;�n��O��}�:�eqK�⬐��e��\Z�m���Z��DW�Y]�������1Ȋ8є�W��G(0��C;ϑ�ƪh�oL�;�C�J�ܯKh4���VLp<�q\Zw)[��n"���g��5yDs�mݵ�m:׷���w�-��Ʋnj�a���l���;{mݤv�:N�(�Qe�W��}������&�ܾ6����if�BW{�w���g&mB:���:�Ƭ��F���fp�/Ĵ�V�Є��};�zy8ˉfZ0+���h,��;]q��V]v����	�om
/��36��qIG�n��� �������S8������&plĺ��TkSP��;�j�J_�SE�(�ɗ��Cޘz��m���8`����^�`Z�$�1��CH�^Y��0)Eu��7��ͳ5]�[O���i������͐f �~k��EbH��}����5���h�mQ�o���e�z2S� F�Mʀ\c�&�NԎ=����>�p���7��2.&�d��x�wR�N6X�~þ�!a�����5�/}�m�꓊q�&6�5	O�q�m��Y��ȼ	��҆44v�|$�ku^w�g��-.|���+���M��=9�RCl3�5wL"��w����u	�u��l�vCɖ��_����T���Zi��x;�uxѐS�ֿ����n��}����[U=~��Ea	�ⶁW9Z��G�[�0����[ج,��Δ0��I5�}Fv��>��N�J����&����1�K�Kg:M�c��޷>��UeW/��Ʉ�32�RÍ�JZ�L3\@CT^w\
��"`��}�� :��1��#H���xR��Soԙ�N}�Fl�u��d�"�i�ku����?\���ﰬE�oS�s�y��_v��N�K9�We��]�vu:AK����j2jp�|G.�b�\�V���x��=����"�w�m�Ut`�iM~����P�u�8������b����N��f�8�����d�]�t��\Ԋ�)��,��ݳj#�<̴��W�w}���n�j��v6��畊�K�RY΋߳ǮE�0��[��i�kv6l���+}�U�r���J}*��\�.q��ؘ`�*�{h����ܳsH��N�C���)�*AO]U�P�'�흆�&Ew+d���mfЊt*:sM����^ ��v�3�Dm�gU����r�����ƽ���O�`�[ڨ4}����ŷ��}�א�7�$g�vf�6���^{���ba2�=�;�<2~�?%`�gFU���{�f�>Hi=>�E��]H���Pm�k7{Mt����#vqu��Ĝ$�?Xc;��^q�2}�p�4:1g�����J��-�j�U5�?</�xm{�i���'䇚�Cz��I^LB�*�0��=v'{}3z1����e�@f�Bs�k����)��{sO�t��e�Lv�P��џ�m'�����]}����7�A���Е�Ҿ����{ib]��OS�����#� ��gr)��#��;mm�.�ʝX�_�ꂻ0��c1�I�D��<]��a��[98@�6y�ڧf��Ѥ>K��'��U>gv5�ϴ��ϧ�5���}u"�k�\f���f��ٝ�U�/Uw��ͨ7pxou�u�.4�}uވU���.0�F,�~J���.+.2V��;�R�g�C�Y;�,��I��S�ZdE�3��2�l�o�S�Tm�+qv��n�a�|^nF��b�ٵYIw�l+�6��p$��x��eV���<e�O�(˸�'�����K,���5s�v��^Aݙ�p�N2��9�"&��1K��E��8��|�y�y[�
ob���^��}���
&��4B��y (�.�#LVzU�iգvV����AT�4L	�m0G*�n�*as%�l���,��}��+�2d!��v�F�7v������G�6�Z�;��;+ل7��Q�I"�OH׈'i�K�ǳ$�5/��v�$l�/ԍv��ٳq`�޾��N+�Ox�U���VE������g%�/�.�Csj�q�������f>�X��bmG.��#ɳ��Yv&oBi�]��m>�.�������Y;/���V�$R��"�� �GZ��c3<�| �x���GԷn��q�$�l>�أv��lܼ;��{�+nT�pS��J�����A��	���x�e��<�+�g1u��39�^0��3�����.V�-��Ն$ױ͆�A럑w~n��sq}��t�t�)<�Y�G�W@����u̱4,44�sq<9LOi�%��*8b��/�K�sS����V�f���ڦ���q�p�43>:�zxU� u��A�l#�P�656�x� ��.�zj�����ie�C���,�N5�1yOx/5Ga�d9S�f\�*��f��5\)�
gWi�����%��E�	��q���j�;��x�[\:=����ی����v!� �jN(�������JT�2@)z��cڽ����Q��\�=�Ѻަ�^j2�<��Q�3�ѻ	e��D������e�F�6�?;�ҕ.�����෎Dx��W�po<
�W:q�K��NX 6�T�T�u�L�ŀ*	�R����%c��n�9�R�&7�>�7p�v^�]x�x�j�_Wtux
�m]f�&��Nt�;�9���G���y��� �*�8���&�Y��{�sO�6)��W�����q--�z�[�	�ec,��+l��-�ϛc��[�gh2t�^t��|�#J�6shA���CS�O.����pY"��-9&Ы戜��֫2֐�S头 ��n?��U���2�ռb��+��T�k�T��`uv�K16�U�A]�[.��+���pق e����f%LƬ�\w��\N���	M<9oA�>�\w�
7��!�|��g�C-�� 	���%�^~hj�w[b!D��j*���`��*:�h�q�5�wy�R�����Za�\��.Tz�>g#���c"":�D��{�������(��u2g;�a�"�f�+6/�Z���7.��E�����G���*�đ �����6N�ƌ����Y����XdE�b�i��n�yų�Kڙ�歮s�7��	*��e>�x��9��S�{��Df��;eeG�����p�6��t{�j;h]tڄ��+���
]�knŎ�b�4� z9C$��gK��쬩W��u=;/�:!��[�����v&���w�l�� �\ݕk'���_uҫzp(I�R��F��]�7#̷���%珆�w^^�0�j�2�UM9zLP䆒�akz��i�W��h/��Cx�ؚ����>���P������DV�l�Ԯ'5[P��γ?S��O��<��d�)��\O�5�ɨZ�U�ꧻ\��gҵ��S��ZW́[ǚV�ܯa�x;EP�}7!'VAok񫹨�9�Q|ޜ۝�ݧ�h�ج�V�y��T}N�6^��ܟp���LׅlѤv��Hn��S��wY*��3��8Ԋ�)�{��8�L^�̦k�)�Ր-��pӽ͒�Ē����楂�'0�d� �*P��~���F6�(yr\.X[z�*<J��!D(.:���K���dޞib�0�|j\��W�&6�E�ܑ���j�(�ws;�"(�$ϻ9ݙG+C�΀�ϕ�>��e7���7���R`��ȳ~7����u,�v��(���J58pýB��;
$�b������n�f�(��������6��lX˹��N}8�齼q�v܆́aw�Qãq+y��ծ�ս{��z�;��B���֩{i���ݜR($W꯫�f����"�'_P%5O-�-M��~�m�(��Ð�(�ۢ���}�����ۅ�Vz}F�3��A�{��-�ȿO�#���i��u�F�GNA�11��F-�߳w���#�^z��KU3���05ջM�'���P��b�t�[�`nf:�z�D����cL��j��L��|���w��À����S���!��#T<V�����ۄ��Os,	Q���r��9�kL�L;gK�ћx�jU>��"�.�,��(ˤ��}|�nwm�l���l�4�GwZi�o�WڝQ�ַ��,���;�����f�]�F�s��
�Ī1�8��L�Z�K+�K���9ԛc��ޛ��5F탩o�Ü�W�d�nI�*�	^UYX��<κ��6.��7\�n����~ր*�D	���o�n���H�4jVf�f� >��`�SFft^^��t�vgz�&�f��to�������s������m��YiJ�*�ɸ���0�sm��e�jN�W1(G���kZk���4�LN����]r}�Ǟ���}�:���2�T�M"�����W�������GSr�����EY�5���|���n�V�
���C�D�]}QqdGR�o�T%�i�� =w5rok+�n�V#fI��/�:�84C(�^|Y>(�x��s�څ�}q�))����L3B���7}���Dv�t��P�v|Z��B�Gc3���Y�!vLAD@���p�=m��J8i�4�ϯ`��<�����q�;6��7��Ln��*��|�'w�_b�^�%C�v�W��ye�m�;�t�g��wt�����s����h�V�+��.RT�~7G��ۇ7����E�@�2�-#&�d��p�'����(+��_�{7��g-̘̙���!���ZΏE�=!�[�vӾ0à6C��VL���X1�Sp ᣍ"������[]�|�7�6��$��hl1���ձ�-��v�e�>��{|ϡ���Yh����EG��|O���P��oe��	 ��~�o���&	��!��਎�9AR� DR� AO%0�) �|e@L ��T L �s�����@�  �".�  �  @�@ � >� @2* @0�" HR�  HR��+ @2 +B�L � � 1 �M"@ �+HH�Є� 2�!LHS" B0 �HD0���L(!3 �H�Ȁ�
 � �x�(�4140��00	34!"���M+LL L�4�"J�0�$�@�L(l��IX@�G���md
��g�A��3�o%U&UTJE"���������}Z{x������n?�@��g��{��Ж���L~�5��* ��=O��(������
�P�~��(@��J_4���j� ����g���Cm��ܚ{�Q7`wt��V��E�B�)�P!�H!D ��	�	I �	�	d@�!B�	�
)V dBX@�B�F%�@���@��(@) hAA
P )�@
 �T �@
A��%q �D" R @ �0 H�$�$�$H�(�D$",�(��$!#
B$A �Ȅ0�$�JH$� A"�C
(@�! B���@0���)B�
 D�I(K"J�	"@�����Ƿ˧b} U�� @*�B���-��ˏ�	��0�ӥ�E n,v���_1=xO�v�G��`�u `rC�;w��4�W�� ��C�C���-�c|\��,��K�d7
��`�~o�Q��;��� k�N>��PW�h�@gۜ�;��;��{ �
O�h{�A�( ������
� � �40I���,lX4Oe��m���p�v�ӎ@��I�SUI��4�@�zP\>�.��&��
���8h,�aEE�~?�5�����sO�b��L������x�� � ���fO� Ď7|�ҩBBEE*�R�P���Th1D��R�J�B�h�U*��EB$�BA	%JkR�jD��J��
�b	5f��l���[D)��4kV��t��Q�fQ TM�֫3X�mQ3J��J[jR�e����m���Y���0mm,V[(��J��:�����k[	�����J������-f&�Z����٠���Vb�ͩV��
��6#j��
�R���+jĬ�f͕KP+J�Zafm2ٮ   ��v+E��nfv��۹�jӵ��ݻt�γ�5�gF�8ꫥ]�,u��vr�ڂ�p��JW]gs�ݧN��Gr��l.�*KIgGn�r�N�i9jP"�Z�J2J�j�   �qz�B�CB�	-]7
(P�CCJ�Ck�^�	��"����Oxz/vhkm����*�Cm��Mk�ܻf�wNU��ce��v���w]�T�m�6ƧN٥�]ʪ�(�m�U����V�5�<   ;vޡɫme���\�*���8m:��v�k[i�ˢ��9�j���V:;���Vڝ��v�u�]wS�s�Ɗ9է[���ݠl����vj��N�u�Ԧ��[eDM�   ����lԮ]��ҩ��v����K���7����)ݪ�4j���U
��n)�6��;�A!�nut���L��f���3]��D7�  �{TT�����:%B�gn�n�]ӝ��s�˷v�h���ҵ�[Rm�V�����;��ۺ�q@Q�n܋Bګ�$vŖ��afֵ���j�  #x�E�U�gf �u͝�-h�+UV����ٝ� l���P9��'Pgl�7[wI(�f�����S�衭���km�4%��-`5����x  �+ �P��h.��J�k��  ssp �k�p  �C��˸� k  n�p vҴ�!f�@em��m]ǀ  �  �0P 	�p  �ܹ�  FР v� ��0  �+�� ��� (d`  f���IFٳRZ֨��  <  wV�: r��  ��p  6t8 5V  ,��  ܘ  �a� �m��m�lXʳ0F�m�����   �<4Ly�  �� �5�` ����
 -up  �wkp�ݬ` �w[� ;D����R�(0� )�IIR �d���ģ��<�@���R�~�  ��jU5Q� I��&*�� �R�M�[��WÃB��2ԓ��DD:=h�;]�L�
}kCҁ�����W�_�z��|���cm� m�����`�6�����m��c1�@��ظ���
��6XRZ�*�0i�1���"�X��O+oT���)B��:q�V�f��J�]�ê���$I�ո�֝`���i n<��V�'�z�&5u���3�'�c��'�Z�W�����+ul��Mn�2�TFV9�M<��r�`Ȟf�0ELڨ�n�4707�6�Y8��e;2J�Dڔx��clXI$��.�	�<�x.m&��xр��Q��a��NA���3�=�FŤfX�w�b��m��TN�E+!��d��q�'��0'����/�.'�8��肬�������O2YY�V`M`�n�R�=�0�vaFr���q���ij�8����`X��a�B�Q��[��i�u*զ5�0���q�V�\3�i`�iu���JčӨJ��z(�7���հ��T�����:��V�P��TkVRԅ�K]Ll`ŭl
4���pVM��Ip^&`++"r�E�N�A0�֥������]���%D&�!�5��s[�nc�{-�y�ٵ6�K6�%��yI�ڒ#y�V��Y�.�� �X"c+6����fk�V�(�����B�z��j��Z�=f�Y��Ԭ�)ʌ���*�cY	�d�ˑh�V�j��mc�����u ���7\�"�v�$c�plӉ��R���_ZU�m55�tְoFFr�"�X l�R�F�Ue��%��x�(`c�F�oĂ�B���{[P;�9�V�R�����"�9)����t���A�H�A�5����Q9a��NA�S�V�h膱LۺJ�"�����nh ��1V`���F�D��ϐ���6��P �X�������7؋إ��>X�Xi�V�V�܈��M*�h�Գ�{+5k)<�RU�sj7��ِ����(Eq�Keսm�
r�Lϰ��.�;x���
L�)e\�
�;�i�1��n��1���R�j�ݛxP*�j�8v:BZ��T��w
+VҒ��uim^慵��u��L��:��/���1B���)Tv��R�y$�r��1����`c�E-ܘoY*�ᷙ���-���k�6�1�:��7-I�጗��n�3�D[�YMJ"M��%P,3��
U��![X�)a#�[��ZEah;�:[&]��KI����!��r�2�Q�X��L8Z��]�e2��J��v9�w,0�H�=D��Gr��{�ٹ�C��!
u���O*�c�ޫ�q����+f=AV��SpY�S��e=WX)X���Xu�*�wa�!�S!3�%�͕z��&��me&�VF����U�P!�,a�ܬ��b*߮�u����GL��)	0�\�{�ܫ�ֶUdgVenj��V�0Ĳ�M�Ss$��;��+h:���H�h 5*<�3	q벋��$�l�n�aj2`N�$ר����t!rZ��j�i�ǎ��<�<Jx��6bsn�l�;�Ŋ�tI�k�,|�Z6\)H�y@��ؼn���H���^:	��!�E-��v!c��ƝǤ�	t����2�;���mV��5+��`����!���X�4m�q��*8�ֶ\�U�	�2+��Գeb��d[:DhE)����t�i�hVJR6�����l��SZF]G���N��p�+�)�KwqT���T6���m"&�F���k�r�)�vb�%�i]�A6�襁�4vV<�,��e�U?�n�Ⱥ�o_0i�m�F��׼l�ܛ�J��H��cY��4ו�ZU�k�b�1eێ�A&2�fA�Nƌlb�,���	jS�`���n�l���om˦����F*ݢy�������i�ɢ�[���:�*L�ZWq�Tr�i:�u�u�v�b��[Q:x� �Cj��y�l&����2"R��p&[����E0j-O"B�,�0�ZuR%�6��Q�k%z%�Jk��(f�ʋ+H5�� U�wQ�h�'���nA�gImPK�{�\���Æ����.��u���ڄP��b��� �LV�t��y�d���ca�#�R��՚����ȟ.��~�]j8kcjӑ�&,�Mx,vm���
��J���'l��KB	b�,m����Ȗm,��kf8u3U���Md�LWVLSCzH.�qe�ƍv �6-�B��t�ط%n�eW���5��CR�(��[v�5A�IJ�̒�ۻ{��X
j�+�"�D��2a����h���kq�Q�uڽ(ێ2	�Œ@mV�W��]�بh�%�0� cm�����z�� �l�:$�����];B�j��R���#c�i
C!��h�S؃̱1]Me�� ˨`jެ�\��d;j��6�����7ġ+��Eݫ ���4+�L�[&$�p�.����L;����_{�3l s���Z�dj�dw,��V@��d���y9R�	�� �e:R��ūX�w.�e��VSU0���e�v�X�d�A�5l�0dFc�D�ʲ�Ӭ#���D��X�j����!di��z��8$)���*�R�R�Z*;t^[r���fEK�������fY��l��q�31�a3@F�aR6�0X�5V��㬒�%ֳx�)�J%�Y��l�D�1��M�j*��eƵ��U�K(ˠF0���,pˣ[�#��f#��,ཻ�Б�勈��*h����N�Iʷ1�fV����K�&��i���a�m��CXf��A�(7�K�z���Gr�˽q��QmFT�V>�����Y�Y4�*L��qX����<o`��zV]�2U�i�W�X�fcߜ&�
�$.d���ћ`ې�!���:�^�4�Ő�H؋&h;ld��Q��ndj	j�ա-3����V��Ҵ�*čL�a�l�ȭ������8PkRśtVZ"��Z���׎]�T�nc����f���Iibpb�Ǹ5��i�gM6��qP��)I���nX�/ffŧTM�2E��ǭ��	-��XL*T�}������ض�1f��K�eh��ޜ��^8k5N��u�ķGlZ��%g�j�:b�����pk2��7�=X�PH����J�lۥ�e�7���}.�۶U�r���Y��CY��0����XFCXԛ�'xED��s�Ф�Wzkf�mh����"��Tn�]5r+׌�?�ą�
[zl�U�,4��X�l�K�����kn���֫Wz,�8�H+в�*��n'HзH\�
/����-
�α��,U��Y-i@�L��
��ŷ�Się�GPtؼ���R��*��㱃N`/X�f�����2��}�P̙Q��f*zAP�bJ��`���*��x������ a�
��[������,LOw��p6�xY��ZM��E�u�!s
�	O/i26�,���f-�]�KE�*��]2�:�a��ٱv�)�t+�«r�N��*^��m��C�i�[��<�S��l`��x�Csq���*��`� ��&�LiV��\����
�`�fwv>
���[
e�V����ѯ�9Gikb�j�C�CM
5ж1ґ��3�	C/sIZ����X[cV�Gʶ��DPYq��7�m����
kh����@�/d"�EPHd���J���x��&�FV��hM,R$�� te'�-�7,Y*Ls7l�
����6j��EX�i�tĒ�[*ʬ��
	E�T�ו���X����d�s6]I�5��M�B�`�u�8��;��ՊTŨ��An�ٹP�-�,�y�oB�%�{�7AWM �����-ۉ����%�EV�;�b���NKk'̌�]Ǥ�ޅ*���⽴�tԂi&��b-F���Br�멒�K�����`S��X�@�/(А �c�B�fP�M:v�Ʃb�x�l�)��[7�u�Rʖ� 
�tL���@�'OV76�((�r� [�Z�hhì����R�&�f����cG�B�2]dX�U�	Em9tq��>J��Z>`e�)^'�I�2�7�6b���?�����tc��u}l=y!�ǻR2і̧WEB�9��n��¢�$"v��E�"��i������P�է�3LN�$V$A9u�:��Hn�/����EY͒�ڐB�f�%\�*l�b*�x�Q�Ҧa*1�b���D�ĩ�Գ�4�R�!DT�Q]���B�i�����L�w���NVY�����l�˸�ڌV�h&�J�ޝ�6�֞]�ڌ��Ǚ�L����OjR�+p퐬����Ӡ E=Vl[�XN���lY�D�	������b�{VѱV��#n L�[AU�%�W��y�u2͈黫9���eT��j�నn��*�KQ�{��ڲۧ0�u#��V;�e,Ub��x�n��]�<jJdB�;�Q�ٳe��4]�YSwG�b6�3�P���-�lcN;L��S�32�9,Kʙ��ոP����9V�]�)b8�$T�!v�W�Y㲮�E�1�2�'3e��\1�͏͋I-R��Ȁ�'�ɻ��)��f÷A��䰊�R��L^����\�B�����T]��Z�A%�KM�)�E�~H�M�؀±+��e\�l��8�1�Sv�5i�]Hd/nu��@��n�eL�*�蟊w���BM�E��m�V�B��{r�,j�����O
:%d�����-���%z0T��˫�5 �,FI��0Q3qPF���_f�Q,��m��G/�Xc�F��y��F�ِl3�'G1;�]9�v����:���Ӕ��eⳙqb�D��#o1ڹO1����S��Sy{�����]]0Jt0Ӎm��ANa��1j����'ZE�F��}�1��-���*�MnF-C�-C%e�:�+FSBx��FMf�Pӻ�.�Rɻr�2�$j%b�k7L:IIBM�HI��f�,� ^��q!���2�����0n(�Ƥ�Y�w��-�E�j�-жɹZ�
/t�X��ј%%
#�	]�*ư�gKW����1���G.�X�h�-�PM�s,E�][��ڔt,�3.Is��z�_j� �P-ѓ>8brT��RX��{3>kZ�]D�F����`�ɹ��!p\c��f�4n�K�쀻IY�y��i�E��̽ѨJx��,T@�XsZ�Q�"�e�V�麂�#p�.���nA�1x�I��T;�Hx����dV�zR2^�ڣ��2��ؤ�C*\��Z�z����M�י� �A��eZ:�\�e�ܰљ6�U*�v���k5�_�QYպ���ޡ�*�7-]5 �LJQZ�Ĕud)h�(^�@�wb��Fݳ�Yd��F�uA٠���ƪ�x���z�+�N���23�.�AZ��`�`�ʍf�ڽT,J���9�Q��a�F��X�WSr�Ԡ�N�ldۘ+�t����j V݃YƩ\;�Bfa8ĬE�̺dwt����`ZeZ҆�y��d
�	-G�SǓf,4�ݬ��+d�x��#�U�8�^
Unǃ^�[CX,�=�V�3fnd� [u3�T���w�u���(��\qX�	���y��լ��Gj�r��M0p�%���l��{zi���6����!QMK.����R����ͦj#V�z3D��S��U-�b���i[�a �CI���4k���A>��mu2���RW�����L���T���sUm��h�i�8έa��Z��jp��n)�ʛt�܂a�ʸ�4��l7V��2��f]��252C�kQE�c�4��#F0p�E�ҩ��,��MN� �W)dI�v|�+�%t����A�����Hur�sh�`Z�^�t+\��!�L�4�e���j��,L ��,�R1���*\$�NJ�;��2�e�.��O�!20%d�4HNYuU7*-j��^�Sv�q�;V�
G�i9�2���+e՛��֬f�eӸ�խ��9��Z�����Ԗ����j�Z�Y�+d@<nY��!eъؽ8*��U]Ʃ�ݕ5$+ߢ6kE�X�G�U�JhаU!mS���j,��ו
DV^�.�F{���F�G�Ɯ*ٲl`b�ZT���Tqݧj���3w��`c�w.�B�}kJ8��R=�x��aŊ�5��m����S�ڧa^K�+Vm7x�2�̵vr�**�d���Qed�!e��h%m�Sq��Yi�&ύ�Ҷ�=iMWt�G@0����h�$���DR2�]���Ǻ6eԷi��B�$�ֺ�@Tn[@Ʋ��ͱ1`���Zc��`c����ŰâXx��m7��D��C�)���7�*Z.�`�^BD�1]
��ZXU�`R=��b�s,wH���mȨR&]��@ߍvr4
�r�6)�l*4�Qԁڴ�qb�fh� �Vu�i��D3K쫴��;)]̨.��sq���Q������$N���Q�X�rԗ6�F����C[N��ٖd�O���m��q�0��8�)$w�w��"��F�4�	Q�t��Z�̖�]i����=�zM鵱1�����B��dm��˔�VAR�$bW����J�*��wQC��+�@���#�S�r+��-j�aN�Pt�5���x���uwV����	�@�&�Vk.��n�RW�-�\7��v㵵hf캵J����vZ���v`02C҈�gO��N}1Jؘ�[I}bF3�*6턙�k,0h���9����r����̥u�
Um��$�1,��gvL%\)@�JO`b<�#�gf|nˊ+��W��ȳa��3�n�{X�Yn��Q�j�ˢ��
V3t1|5�5�w����/�u`tL��I��q���:-�Hs�3�� ��L@�*ͧYkL�!V�ʜU�=�w#�;����Y�8��$����-��o�a�'F��KG�\����e��ѩ�m`�q+Q&��J�fJWe��r$и�맚f����U+�%�
��1�5k�bmpt�s�oy�V� �����E�5szO+]�D�ΗpY�{~�5j��c��L�kֵ�A�l�CwIֈ�,1��و�P�^6���w���v|�]p$^�h���v�����n�\��:tǜ��	TAÚ��F�v�n��d5C��m4�q��d`}�\'��nV.85.��V<�F��c@N1�G�����[v�Xw���﨩�S
��qt��8+B�0XP�#�3ȳgq[km��CV�\���f��;�Z�9�LY@f�b���pf�SB��*f��|��v�Y��,^n+۽*��8����>c�Η�'G�-:��w-q\kZ����4����v�w3�>s�k��q��m,�QƲa��lm��\��Hk��jU=�%F��o�J���3P�B�[]ˣ�U�s:�c]q<�kMx��. )2�����Nu;/b�V���48��g�b������Sv���YG
���<6�(�i��u)�.��)or�H.u�[�(�Xe�S3n]'�:�ݶ)e�&n Y���+���yE[�(��j�w$|o�G�uy��VƵ�g��$n�J�ru��ܶ�n���)�!D�˾�á��ռ�cV���vG���bǳz�.0V-��]s+{����+t 70���>��uY5.�f3�7,m&�n��Wt��^��eКE��J6:�'��3�*2z�Nf֐eN%�t�F�Bd8Nz9�2�#h5�϶�{&��`�5;sad����a��b��'FM����P�PC��}G��h��]�(eԠ�e�9t ^u%31�NY[�L���d�H!/i��XD9)]�2`��&n N3اe����\�^$�hc�:��9�u��'�lLJ;.��*bC����s��tu��#vGwd]��5%Z�g��`��3��wa[/GZ�U�f�}u�|	v�� /R�r�|_VT�y,�EWյ~���x�f�JV�7Wͼ��>������6���n60�V�r�ل�D,x�q�6�[��:r*C��﫨G���4�!c]u��n�	���׉d��
8�kBve�T\�������;U�2n���I��/�>޻C3-�����#MCR�)[|dqS"<��ł3r첐j�ۜ,u<�cF�N�&���\\��F�u�5ݓ&LR�5���Z�Y��4�T�_G��(�z��K���G��u��J�°���F>4.�+6�vH�ۆj������F[ȷF0v�v�.�:�_LYٌ�h�V ��0��jO.��3G_ґ�QAv՟{�c��T�H2U�i}=�vu�Õ�X�g�:�T$7Љ���b�4rֵϭ�$�/�3��sk������Cw���m�)W1cJ+��z�!����i뽣t'T^��F���::�ē�g�`[�B�@�H��7Ư��ۍ�{٧ts�S�����Z�)�a�utM��9�'pt�
�z܋fݒ���m>B��L�'��=K��2���AW�gn�[�|6�bi<v�1Vc"E��P�a�N�*�hW&��:��oN���S�SE����^a:���L�f+�հ����"0�DL��k�IS�F�/]�2���e�9�N��9+��$���˛т8�b*t9��j�sz�IY�݄!�	�]h6�SA6����.��"�c���%]u��U�N���y(��[��.Hrs%�rԚ/5�I��Z��6���W���.����+<�n�BgV��#�F�u
��{��
lcU��|�����|*��7-[�Gjl�4Rp���W�zn`�9 W5��Q;q���և�ٜ��6�7��|����d����e��F�SG�)wIU�f���
�14�.�cWZ2,�b��^�\�:�|40X���vb�P"��J�����T��5�r;���s�2�m��;%�cQ�=`��;�,�L�
�n#1uL]��\h�5q�KX*�^�6[VR,����7-���Ӱ���T�²�;���33=%�y���@�l��4�.lGzA#m��b�t]5P�ܱO�W��HE�So����7�r���x�6���U$�Io�u��I+5����J=&�®�ʣ+c��(����Q��G`Uˍ�35�Lx�d��Rea&v��	|�ec��cUGִ��<���G�vu]�ǳ(�mR��X���Hm����9�]��_�i3�hj��QH�ܡ��DCan�̥��n�h�X�nh?x!�3���y�� 4�YY�Jw��M�R�%�ӹR[R�7�٫�YEJdM�����ayEW����A�ϻ,�dm��V��c����� ��W�3HW���^�w+7Wc�O&RjZ�n�R����f�8�W07��`��-�v����`�7��KrW��C
�9�̤�4z1�G�^�_>=x�h͗����iz�6�2'kA\	���l���`�(fd��6�e�T��v͜ƅ��1 ��.`��q�ԫ�I;SI&P���)��\*���0WA�#=k��FT#3��7��� ���:��4��Ҕ��Ļ�Bݗ[���o_ -[��m�����+�ĕP�S��=����s��f�)C}�u��y���]e�l���u��|��qvFf�W�c��e�i��w�����dn���Jb�����k�xq�����A9��o�S�]{5dl|7�I�kZ���=�cp͋V�J���Q�X1=f��3yܺ�u��@X7��|�"e���'�I��:��*6y�z]o8+���󊦸S��='[�K����Dܕ0>��)S��feÌz;\���0]k�Oj�����	�	�XE :�|��Y�x�}�WN�����{x�3WB�]��ine!�7�h�r7����$k��R�����I�����sH��uu<}�0.��u��D����r����X9�-��6��Z�W#�䥝���펧eJ*�NJ��ˏH��%��{��[�iF.{�9�i�yM5kt؂��Ր9np�ek����t?��m������(s����][H��v��K�v���R�ͽ���B�-���2�!��b�Ornp3�Z���q�Ӱ����Z�lr��^�7�(s�4�c�vȈ����&ma8R�]_u)��շ\�k�.J
p��Zo2q/*���XuU�Su�m�Z�|O+<ƻp�#�]���0�ˇն��o�y���Y�����%����v�f�Z�@��hn�5]��6sOq���Z5��q�E���L�*�Q#;tm�p��(�v��l��,�L�oO[v��k$��·��Yʱ5�BǷbZz�mA�#�[45��C���w�G^�5�6�j�{��W5���ow��ȩ��`RAի�$�{�]&7�=�%ۡ���i�;R}���ު��F`xu��,#�ȴ,��wqVA�����P�7V�V�p;܉�ୱt���n�wI�����E5����N�_1ȉ���;Gl�E���
�2�er���C�e�������K(,r���O5k;+:�Qm�.S�+7���zJDWVs�����yc�����*M86Z'�ztX�
/��~�;�����"Ν�i`���B�շ!=�7F�f�E;�!��s�Л}n̳θ(`��`������,�@�EnT΀�$��n�Z���d��Mmŋ/yf��(b��K�Y�٤��Tz�V�vT�_օl)�1L����)Zm�YW׺�VrX!�Xݧ#ʜr(+#�܇���Q�r�]J$�g`��U��j����d�K��Xc�����+-n��|��������{Ώ;���Q��2�CV+x)��͖�"��׀��2�ح�����ݼ8��G��7-�9 H��Lx��.��-���uv�$�ɲ2��q�dw��@�����XH�{K�P��B���m
x��ⓦ��++��3YDr�#hHol`P���s.(r�TO����G�B<'s������*�sH�`�r/�WU���*�m���t2K7/yŖ)g,Us�Ho���ݭ���a�޶gA ����X��J
�Ѩi�i4�J'�����:.%LE(�x<�7!��M�5gh����	EG���m�m�u�����,\�nbĊ���՜�=x3�=I��f��8d�Z.��F������Q1��6)E��1&\zj$A���+K
�µr@�]s�`_�t�kv���i�f�0�W;��x��΂��4(ԷD\Ԟ��b�_\	v!�]�fT�NtI�%�;|�s��CYW�YAU�������PyG��kX����d��j�R++'ƆM�-f�6��n���z���L�y��Xv��x���Ύ�SJ�knPV�����^.�)+fa��`�V��\���=�: (-ץ��E:�e۔��#n���T��g�{�ҙ{�y\��y��bv��U9ǸB�KC�IDtV��⮜딇��=H�w���3����P�`t;�=��E
��l2�ۼ����"Pǩ�9�ޜ̆D��yJʠE��gK}m�<�VFE�mL�Pt��X��mݪ�z
�5l]u>0�wOzF�j�޳SU;$�;���v�1�(L�s������{���{������s�D{���4�)���"�*�{$��ew:���ŭ���*[��m>ŐSARܽ�9�U4fmٕ*;����*G(���]qc����%N0SV���-H\�:-v�������ۣ�W ��[*n`��)X�������r�F�*��6e̚Ⱦ�u��,�5,WW���}hv9�ƻ�y�r\�Fн�I�r�7+���f��8җ���.JCXqơζ�ShE����l�|�N�,�B��RО�me�d�E�)-Rv�ʸyN,N�T�I{}x����T��9���g,aе��V��NSγ��a��9.2�g�im��K']����8fo,���[�̝�������0��t^��^K=1���=�ge&$�uz%
��N����-�Oc�=�K�|1n��Tқȯ"�Д}���N��&�l���XU:��ψ�ݧ-U��i�e�ˆ)raj�����*�o�-�l���uyu��kB]�ٙ�ui@�r}���Xb�!nBe�sUɗC��)�.����a�(��C���4���ي�Wi���85�u��scPIp���)���^*��,u���΂����	�+����KP+K{3G[��VV�.�i��6�6�����q�[N��r�q;8D1���3��M��.�T<4gGC{Dj1��e��j�Y����*��'��q\b�[���� �۝tP�f�%�*F�����ܒq�{��cO<�..ˠl%N��/9�����ȼ�7�eɜҠl}E��ע63�ͤb2�f,sA��<`�b���K��ڭ�S������r���ֹR���v���0ʸ�澴�u�*��D��[2����X�o��?#)�Uӡy]�S�77JY�����Ȳ.��ܜ�:�`y\�S�$��6�=4eCf�^YT��enu>;tl�
�!@�1v�B��f�∔�٘2���Գi��<C|��0�k�*`�wد��B�r�N1ɩ`R�hgZg�����p��΢޹mh�65[���"J]�4�٫��~ow`,C����g5�M�30 Л[g9����C�=;��C�5���a�s!��;݂�Gl��ʵY� ^.f�7���T�mc<�vE������ffT+�\_0*��+��6���j:NB˃�u{"ެK�Ms���;�um��UC�ew*S�(Z�x�Ԯ�%s畖#xQ�pv��V�(u-�򊉦��eh[ڱ��5��š����m�5k��$��5�-=�.��'��c��@��"�Zǻ{�=�#�!s�l����F���G���I�hVo��{ne��s���׶�q��nCuċ��j�&��U��U��Tƌ���?��F�r�J�\�x�p��D�{�<�!5dV�O��n�e^�26@Xwkfq��-��f}�.�.,��p60�ۚ7���&�8.tLʝ�%j��"�(�r��=x�5�����ۛ�����Zr���T �yp6(R�a���\*���V�t�9</��wH�v��&�������3��B�'1�GUc�e��B�1;"�L�,�곑�L�mGha=�m[��Բ�m|�:��
Ѳ�d��z8�u1��J��[�oV��NoVD#j�%�������{����O/�lB���-���2c�a�^�.���n���G_�����HR���MQ]��E��ܬ�8�����ָ�qެ��$��t۬��}���em�9�����̎����$�W�Ύ���J3��y�BO�gz"�7�F����X��!κg��ݘ�v��Bq�+�G�Sצ��E�qAJ6bջJa�{kѹb�ͥ0�C*���\_�����H�S���:�۬c��ȋs[���!��(�Tvv��q6@H�#3��p��C
Jl�-wf����M�n�LlBfn�ɥMk�ɤS'p��=Ik>���4��=*h�u����5C��m�m:"lֻm�ϱ�*�˱
j@9��,�p����gScb�gn�nut.�+��T�K�.�Z�fJC�&̈́r��;qo+�%
Pd���w����bmT }��8�4�ns���}�*ћ����Cݡ	/V#ɰn��ճ/N�8q.+�Փ�̦S�d��JQb��/����b��0�CsB��.��+-�����l���ǧ��� }����0c��0cn����������<�$�/��us�����gY�|v�w�jƽڄs�n]����򝉦t���-����՘oP��f+;�Q7J��a�;7�c2�^kX5+�0�Mڔ���0vH�Z4H����֚bƣ��c�Ë0*J��ə�7�j��u�
:ڴTvr+�u�0ǣ-�ڮ�/p��m3�M��*T�7â��N\��L�̡�Dә�2��+{M�֡���%��N�,)��F��Q"^>�$=�h�I�'j�+.IB��f��E(@�7{5�n�ښ����V�0�Dï�R�A������Mۻ_";(�����:y�vc��2o���l5f��'GȾ���6�}C�)�|�]��n��o_f�#S�3����1a7��L.�qP���Nޝ��>ElA���q�T�hht�32���6�@�1�mr������b����-��t�ߤ���(j�����4R����FU�Eԣ���S�]>�1Attݞfq�mvw��!�_`}��yG\̮'�4�Z�s].pĊ�j���_yaJ�:�c��q�����v7H���7�&M�"���aPlEK4�	B�v��4Z����Jsq����9�\���:��qm��8�#�9����Yr����qԭ���w+k�<!�%�5�BXst�v�SV��5w�F-O�]���VڎX�|,"4sD�o�Ŝ�Z`�٘��Z�Ť��$̩�)��KUu��74!TцnG��t�t�ǯ-g7��+�@I5 ��)��,!��o��ma�����G���JW�������87~W���I6-�у%sI`������[�!Vm>L-��Qkd��q���.u�����[@����uP���-<�E�Rܤ�ʊfY5CNlWM{4`VEY��#uy�O#��a�(s��53sk�G�l��a���:ij����/����OT舅c��_
Ѱ� F���g��ŠP��]u��cX��NT6k.�
إp��0c���$��o��^e5ɈG���j�Je;o���u���[_#����R'1d� ��9��}\B�\4����A-l�٪��m��(�%����'Q��/&h��6��tGd�z$�i�{��ƴk6�R��
u3�����I"�D�0,A�I/{�I{f�vC.��P=}��5Q}�q����£��0��o��9�M��+:�wB��x��,���BT8�aJH���Ew	�REXu��]�dx���΢4|��{�X�"�9�:�Κu����o�KWf7��X�|9�9��P�D�;�.\�Zܫ�'�[X�X��P:�������,h�S�{Yt���2t]f8�!FP@)�d�o(��r�d���PK�Z�n�.[�sx�v	�Y\ˬ�x�[olb0�]��;���7X�(=�G�"��/W=x�e�K�)�>�h։��ƃE�ٔ�&{X�������T����-u�f&�G�����6D~8�y ��E2뷶b�k�X!j��_N�b��.���swE�h�۵.�&�S76���v�����qk��r�prt�G�Ӻ�p!�%�:j��H�Z�q��[���62���`�c�6�:����ud��|�M˲Q�o�p�(�=���L��Zʱ�E񼾰�oQ�aj8O�ws��<FΜ���C��̳��'���*�r�h��f5�8_oJ�23��	��
��bX�ڼ�Z��#��5�Y&�����eB�ݜ�;$���5���oIӟy�p�Z�2��A��/��	 ˅Z��r��,�!h�j�h<��o�o��|:jņ�X�`���J>�[s �Q�[3b����ٻw���u�y�	,�Iff������U�$�;��x�v�З�\���������z5���)�a\6��"���-�~�J��o�:���@�	|��z6T�s޹uDs�5*���Ev�����M�/N�N��S���D��;�vAʣa�)%��@����a�)��vӾyW0�ǡ��:.��W�eJ7&�=2�<Ի��4�C�Yx��SG2!Ի���%}��	m<��]pޠ"��E{c��vt�j�Ԗn<��h����Y[�[���-)�Q����=��W��ˠ�)�&.t�5�YӚm9��t��
��I���7]��#Y+�;֘�3$ ƻL�ա4P�i�ۮ�-�μ]Bmý�݇�{�êT���]#�k���5�J[2kk�`�K�κs#�m���lô��K[�2�R�L����;G\�g6�݀�DW�Ř�� ]4�!BA�un�yH��2ڹ�%�N���]T�g,�kK�[ʹ��Y6�1si�FM��lrnk�Q�↘��·:c��A�[�Ν�h�yQB�u�i.���}���2�	�c[`��R�B` ꅽ�<̧����k�kA[J\�Yj�w���6��*}���\�N�l�W�%n��N֨9��V�:��B�4�4=�'}��P�SrP�'�J�Ӝ�s���yfo%ٮ<զ����s��v��u�z]�ֵ�}Gt�ja	�䍸��ĳ3�n���m�c�=-�tl>&�6��|we�)E�We�݁+��i���wSj|xn�
V��td3{P�a�]��	r�m�5�'�\���#.vl�6%�}�A/++wt#���uȣLO��.Cң�4�`�.��S�EE�l�kjS�T�z��&�b�wX��1>���W[3�b�mvɶ[YEC�.�LO����/��V=+�-�h��u�gC8'6���/Ih@w��$�Ky��Ìvr��EY�˩�Oj+Wm[h�BWd/���]���yZ{3�MZ�S���Zy�>YNHXD�5�	�`�xu*t�	B��w�нF�lT��["\�� ��۽�<0�CT�t�!�B�ƛ1��3`�^8%&�7L���v��{+L�}�lL�`���B�:��,<��]�?u^(�vj�!�X{�9���]�5�L���1�}cf�RZ`r�]�����)I��0^�K�5�\ޠ��l�p��1�8ЮE���6�9FњL2�K8��eXZ��xNC�� gm)wS �c9�-u����u�S2��(u�obD\��ɸ���Q��P4����ѱe�U�i���.�\{1+i�������У��E^�N�/�q��TۋCEZr9�_Wk��V����<QS*uc7y�Fq��Zn�� `�"�:^G,޽3�v�NI��=��n���VvD:ޅ��t�D[@�j���r鑴��A\�'�mNUf�k�]Cg;E^�j$C�iٷ��]��u'��`�X�C�12*�g%ˋڋ��ӳ��O.��\1�d�S������v֛��aK��n��뺻s�f�ᘍ��-�� �����Y�`Ԙs���Y� ��
i�_u��q9���J��y�2͗�Fg�+l��l[F�Mm�
_�1g1��^H���q�f:�a�(΂ΊH]V�E��HI`y����7Y� �Y����n�e
��r��Z��x��=ҷo]���uX�q\��1H�ֵwXT���)��,�Yr�G�����\k�`�KX��p���>�ރSi��\����ԝ^��.M>�"��w�EC��una[�,���2�UePAԃN��)b�aȬ-�et���ˡ3��@4�n�/-���D�IMt��V�M�y�v����:��k��K�ACb�h����e�1e�,�%}{ZbYAv�W��N��ҟv������]���P�i��ܰ�n[H��Vo� wkW-�g�ʲ�H[+	֚�T���c��(�E��T(�$��gk�h�"ʜ���2g��y[�I���Y���:����(�w�B��a��Q�H8��Y�g��
z�`��b̬�x���Э�f(�,|�R펕w[g��{���G762����L��)s�v$P��[S_d(�X����
K��q�=v�ȶ��H5YZgw>ଂ�A�Y�%u]N��H*�}
iY2�r�[�wI��rto��x���v�ŵ$���څ:�b��iiE�r�����������j)�-Y��2��J��&;Q������k�]3�������6�f�-Ov���8��ո>"lZ)ë�w��Q?-���:T@�P�]��2REf��dg!]n��b�n�r댗@�%tк�-Y+_�-��S,���Be����4xF�J��Zw��,+L2�\{Z�;M���*_H�\y-.m�η�u��C.�ɨn�K�-��_^v.��M6d�џ5��;=�����tq}��N�ͭ�\%���2��i��Wes��f���%��&��{�%�:��q[�6��Ә7� Z�1m'k��[�����qu�)sit��P8Drr�q�ȡ��m�Qp��g�r�j�΀ԛK>��M<2��#_\[��h�_ 2}�͗JZ����0���.o-u���R�Ws��_a��%UR��pn����wK�\��V�v�W�!��:��c�vX�Qr��q�٫; ;��S��(��ݽw6Y�B[�K���P8mv�WdS5��s�2u.���^�.U�|�ۺ6��2�4Ü���Y�r�sM��>;���.�T��p��n�Y{9J]�7�K�<{i���ȊD47yv�]/�E+�*�d���YW.��t"�W����s
�:YOE�.�m^d�rXƮQ��:v�b�W��80�D9�{b9D��k��s]H�s�o��61!2S�.�(��A�5}|�W`���WMP���I56V+��t+c'T�wb�.�s�/yw�"]YJ3�]����n;#o���N�Wn`���v=��7���۸[u\(n����<�]�o:��ü�w��i�U�a��N�m��#V��S�t�����t��5�,e��ڗ
#Izy�J�V��f|ҖpY��;dcI�0U_�O�9*R�����.���m�I(�5����ؾ�N��L&�귔;Awmw5h[־*����.3X�1yt=y܂��hK��8(M���3��u�y���+���4�h݀$��K��]\��2�c;o���)�����ƜyVue��!aTْ���z�X�W�6����>h�=��]��j�t�a���wN�a,T�^�Ҷ�@S��W*�3AG��K1rV�"
�'sNaB�KX�
I{V�^���%j��U��5�2���Az�L�6���4�
楳}u�^�������A��'p��厝oW��ʛ�O�R�� p�w�$ڮ<�����W��<C�i�5;B�� l�r*=��xð�'pP�|��U����/��\JQv<��w) 	YGr�Lv�\GW*CiZ�3Eڪ���`�ɐ;��)�e��3te-�W*;"�w�Xl�)��-�5ݾ�U�P�T���+	'����q�����ꮖ�g��p��И ��#���wf��C��T]Z)7�7� e��+z��N�Md,X�me>�x8�;WՉ�s�]�y���wc��HUaT#V���4�!فCpj�j������d���R��Xm�j�vt�(CYf�n�X\ٙ���󫅉Z��R �:��լ��,3�@����r�_
{��x��Ԃ*'8�+�SO6�T{�t@�,�֍=2h��湥���N���o6�N�p�{t5J��%D��IiFt���%c�r�R������W
������t�[yM�G%c����(F�5h����Z<���m��P���Ő֖k\UcE�/L׏6�� ��1�]�5&ݼ.�vĉ;�ֱ�Tn]�J�|$�/7hg>e��q�8u�yOV+6�]Y[x�m�bM�D��
I��C�'[�����Q�d���y���i�+����.SΖ*a�b���(�'�z����wa��'W�7ĸ��i��L`x���}M�̓�r�T���N��t��Y)j����fd)�7Q.*n���{��5t*�Ԃm�����1[q����g0yX��u3�(��v
�V2�"�G���lqKv�k��;�ֳv��u�i��ĕ:��ӛԻP5������L�-M�.�Q����u�/Q,N7}��H>Ok ��K���+��S<�ݰ�SܝۗY!�`��
]�U�{Ѥ�w�M���L��rr�kR����$�p�ӗ7G3��4�ՙ6�-�B���ڧ���N"	SVq��
Dt�Slh�pB���'XeD*�L��b����l��}����Tk�
���5����Mc�[���휎�*��$vt� !�[�t��w9m�Fh��Nĉ�zdQ�Ȋ��#A�g��CFl2t�ZpP(�7,]�H���Fƽ��J�F6�C�K�Lp]>¶Vڦ3�����Ā]v���b�[�NFaU���Շȭa�C��i;��u��h��Rj��HC�����4f����Q[}&�_9�cH񺑙vB4����s�FI�8t��L����w<\��!5P>��ǂR��5��tl:7��� �nV)�h0o��f������V�u��$8�����z�G��X��.@�ބ�p�6�sڲRq��6Y7Gk�P�<ӡ���<�)�oWf���ټ���2^��ڴ7*�/��U=�Z��<�S���0l�Ў��t4��ʠ��^�츢�b�.���U���+n���TG7%� oQ����c��FW7vpv�.P�:�MPԠ��m���v��XXI-J
�cܾ�V�B9��6��E�6;%�0�,��#F��'�q�/߱jݰ��]��)Vc�WS%}�*jJc��p�6����M��E&�|�`FC�b���zkIUX+���Y.	�ց�i�@��Ґt��w��Xz�.�HM�7ֶ�LcUљ�^�4�f:�ԥ�L��T�cY�e��9�t��gU|;�.����|>}� �/� �Zw
�yV5�R�Hq��9��WY�DVl�yC$��@�Y�OZ�����N�M'~�eT�IQp�3��i��/�\ڜq���+��՗���z̭l��FX(�N�`�Id��f�9Ұ�)�Ѧ���dkvrohc"��<���iМ�$jDs�%�j�yk)1�;��-T�SǤ��G���%*LV����m�4(_;�����X�R�ȴ���0�7n�ff�r��7"��V��[�z����osf�n[P���l���*��\0����t�7�X��'32�1PΖ��}��k�����J�0WZ�u�b�ag�Q7i��.o>Db�]-�˘ѱ�{(�o&z��u6uґ���at�u��Xts2൱�Ŭ��d9utf�A������|M)�b�9Vc�pgn7+�&�sJm��_p�/N_<�b���'*��L�����_��Wq+:���љ�3���al��ս��p7��:��gS��Pj�鲯j�6���sX)v�w�u^�pV��h7�73!ǋ@��q�FWQ�X���34Nܖ�S�,R�St]�Wi3
bG��h]Y���.�5�u�&��|�Fw��N��e��\A�,�U��p}M�/e���ϡ�+$5�c��m$����6�?*�e2pNys~/4��'�Y�͍W>=W*���Y��~���YF����:���r�S�'��]+�]Ўp�̼�"�+��E�Ԣ(���be+N"�UU\�&r� ��(�[�Nw<�"��W,���hM�;���XG*�*��r�L�꣮x,�v��T\����s��MIK%�T�EeW�dAQ�͑��-�IU����R��M�"
�Y����*ă�YQQ�QZkAD�Nl8�0���XQ�H��In��t�3�i��Ȃ.螬R3�qs=�6���H�C�;�
�㻅��B!ZD�(�VEȯ]ȳ@���k�K����B�wu�8�IY�JnqÜ<�RBID�6�'\2t.XQQ$$��^[�v����qg��r�Ԫ�J�Q�*��]�Mκ$�8y���2��V���"�Ôz%�+�3�Pr
��b2�4�d�]g%(�S
H���2�rwk�-G]���G�
�\�кVI� �h�E R }Y���>�s7��Y�/�֗lVr=7�d�K��אX&ޫƸ�+0�u`-��T(k탷n��O]*[0h��i>�UV��s��-�� +,��	�_ ����-��1��jt�F�����S���cV�'��:^Vp��r������a��+��������^��g�j­ W<����bU�.��s�v(��af�w 陱, KR�[FX���T^Wʮq���CL�Lu�{��9�u]����K�ǻ�$`3
1D�m�ǔl�� �8=·��
Hu��.��y!͹��Y��nW
xxq����;��0�[����X�{1����C��{�[�#����E�}'�Kn�<�jѡ�a�<#��c�!��(	�<)6y���:��_h��M����ox�����F����l�6{�|�������e lt��юY69��l�q�Qo.��L�W12U{���	�j&�N����+��F3�\����8���t��ZT^��r���x� ?w��,��	�� H@�}T���w	G��˼��%tOM�j�V���\e�r�H�<������.ϼ웋>��Fت���p]�s+�6/;�Mf��*G�����Sʧ�������:@-���:�������zϣUق�ޮ�%��,i�Vf��s���~%os��wo������e�0���u�+���>�ݒ��nL+J�_'i��[��x7^��N�AYva�:
��R}�X۞���3������ѱ̄{M�r�`^z�Ϻ��!肥�]D��n��~�!��议�Ͷ�b"��X~���϶P�V�E����\Oq���Kv�Ȏ�f�ɘ����Z�gu���QpK�덡����7D֏In�]u�Ѓ힜���@�� 1���L�M��}�;<�1��C����,�Uʎ�H��B��Uwn�s��x�b[oM��tד��s����wk ��tD"T��޵��^:x��)��*y6���Dū�����Fu7׋�[�y�ږ~K�8��Q����=�]�"��:��G��kl�	����nS㾍ͭhW���+��U	S71p����jP�l���%��yJ:룞�>8�f�����3:mh��}���X�R�F�Y(\!�TCj���}_k�VQ����j��B�y��� �ܵ��쨋��<;�A�ڄ ���a��_��y^��V��p��cq3���\�p��h��ܪv�j�}_^��aL���H6i+��P��	�iם��`e�=n���#d�ԔhZ�$�av5���z�u:(���uy*&P���T��Fe�����]�R���*�<3d\	��p�VėK��]�n),n�w�ː����J=O/Y��A���u�N�T�"���L ��u������.AuѺ5u:{��@�g�{C��,e�}=�X~�gJ>@K&�	��VϪ׺)U��xo�z�<9����b���~y�B&"}�k�Eנz����x/�e���-�_��󨝞�ZY�J�f���E�����������L8�?f4��y���Ձ�lϰ{��(F"�+
uP�x�����%��p.�+�@D=���<�LHUv�?d5��Aaq����=����5���&kۃє�㚻�o}��I ⧸�_[�bɍb���K/J���MN� ��ٰ���\�����Z�P�Q�@y�+���,���R�u��Dn>�y�s��36�W*pw@�Z�f�t⣤ ��/�x� ]:J�?��ʏq�_�v�e�:�,M��oǷ�y�6l���܊�8P7�>���tGAh��㑪A^�R�R��D�Y�4�sk�KIr.,����]n���h���²!�&��H<����䐅�s}�3/��R7�"�G,Á.b;��neS�PN�e/*�{�Qs�� J[K��A=���ѩ\�OIZ���T� �"Ւ4���ΗP�Ho<���S٤{�uqyM�.��3\�Z,���s^���1�WJ=
�\�d��+V�݉N�`�ӭQ��ɳ�Ns�q�lw؂����Ry0�鲏��gKa�:A����ԅ�P��ex�8����;پLyy��
�<��}Yq��wB��wZ��g9�p͑j�;)UlO¶�y�������aB�c7�R��D6�¦otu��oy�{��K�{�Cl��	hx)^<��Z|�n��w�\C!=�<�,�bmƆY�iGOn6��WM��2�p��V����0�9�Ęb�h:7��a;E����[���.{[<�!���<�sZ��N���̟��6r�L`����!�dG9sjK疱��+����q�F���`m�*�?uK�(n�X=sf�н��"%��;����9�+�Yn��Mv��1�՞Lp�R;��o:Ѐ**|c>w:6Ἶ���*,ڎg��I��K<U�DY�UBF�E����n2e�W�lȌ�.�-�n�S0�0[���׷�P�����}�.D1�����,�H�/�񼜏ƭ����x�8(�;�θ�kّ�[�?�9���Ed���Z�FR�b׺Tߐ�9��e���c�n����8�U+A;�%k������1��ǰ�Os'q���\cΣw�&5�#�������������%���f��B��n_X���pҏ.�E�nB�d'�H���cY�+C}�  ��L%�V[�o_^�}���w��n*Gp���������u*s;��T���P�s�����(�� B����C�T����U��]S�Y��78n�a����:���g��Rg#O�&��'�שC�)� ��l*^�9I�t��X��9��=�x�0�tFK���j��=�|�k�_�n`r�C�=�Lp�D�-.��z�mj��Y��ٞ(m�f�)�n�`��G�=�dX3��k���uX/x���n�jD,����G�v����.x*_>׌�5����)�����n�9��rsi��5ǎ��8p�@p�X��w"��1��%ԶGO,G0�3���m'm-�]�({��v����"�Vl��H���v*����=���忹�^���:���H�<����_cV�͍����Lb����p�V��Q�t4P^^�C������o����V:ϳ�=�"��j#)�����Yq�9=�Cn!=�� ���u��uuK��Q�E}!9uU�����8j1���0�@��{l@jto>��Dc
u�Ǽ��tX#�tV�J��
wYsW��}�B*�Tcs�eڬ��J-&^�dʐ��E4&�t��Ox	����L�n�6q�֫ۊ9/��Nw�윐���9�:�,>�l�U�.Γ/7N=Y%=�/ib]���e�ג�� �Ăr�]�3x���e��:�Fw1��=���Τ�ՑU��!S���mHb+��@g�q�^�ד��ݾ�68�}�!��f�����É�x:�w�E��l8�� �g4K�s{���|����8��G�����_W���؎���`0�4�M�
�z�a(�g�NoL�2��
(ݶ�%�3��}�b���+J�{Q�٤c����蚉r$v�Bk7�[h�Qz�y�'u�X�6�S#�G/���������[/O*�p�Fn(�g�X4F���mǗ=���7���*��}�Љ�[�.&�#����#�M��a�R��m��ceOe��Ͻ��Ҕ:�hht�Ϭ�Z=-WoGX���q��/7:c3 3;!ʎ��8�:V:��c��$o?]t1b�zӧ���]��R;�'�%.늞S+w���/��]Y�i3f'HY����5���I�rE��`���J�Ø
gt�"{	dʮޮ|F�=ޢ��E}_7�\8��U��7��0 �<!q��
��G��j�S����<����<�hյ"�ӕ��Ҩ�Md�kz��a�w�����Ǔ1���N�z�ƨ�ދs��w��[��WT���oK���h(�C���Ad<�-�L�l���"-E�p޺;WyHc��"�D^&QB��u�ng�Ȱ�	B����|�S���^�.Z���*f�.���ՐC9@T-�%Q���4pl�@�����[�w�#��vk�'��댨��.P�5�cP{�D���0ڑ&7��
�%��F�gT���.�ggc���o�N$+����t�� ?w]0�)�Ȩs���s���U����r�*����W�ow����<�!�/M�J�V��?�����.��y�Ev��)��<۵�ڃ���6̊��5�t�d
���Y֖=�>Y�8i���}�83UГӼJ�Oj쀝�X��#���^��N}�b�?����n��?����O
�sk([`�(s=90�͐�W�~Y_|����eq�ct�7����e6�`��e��w�����n��`z��4BsN�L�/#�$*-��T��ol�\c*�,�p�<eË��o73�޵�h��i��3� \�\e�K��xp���D�0�c��� `�¾����ٺ�4�qv�hr��+ H��})P�̪ȍ��+{P���B�`('O:0ꆍ�\�P k��5h!U�5����]����st:u��8�!-�f�v`"v+x3E�w�GZs)�ȗ��-Vt\����r�d�R��I{Ъ�\:�1��*�ª�7�𾓬�5ͭ��eٱkm�w(�w:k���v&�K��qrΉ�9��9>�BN�$uG��@�8?9��%�:(�����-(�L#Z�{ϻ)j���[���}SԬNz��%DmBOr� �'�B�+܁7M��.���g�az���Xu�k�x��Y�-�.cDp�{�Y�~�D�3ޥ\�]��+��XZY}X�y���1��+C�ݯx�9�s��f�f#���5ji���ͯz;�N��l����t^���	��b�7r��4>B�ul��59����B,`�"w�CtsZ#� ��P�U߹=��y��k��t��G����y�>�
��6���N���kw<!�18ST2��LI��,v�M�7���wJ�E����Ǒ�9�J�}O��6�8?���pt!)��w]7�a��P	�dzl:�����/���~��x�7�h�K�T��p6�	�fx�>ݿ���9�1���82�r��7<D���o�����f��q�#\�G�b����]��v���[0^�&��Q-���@��T��4'YN�cV�Yv/���|ъ[��vt|��Cw��u3~�k�;ALTE�%Y�t,���h���d١n�wZO\%��s�4�#t5�7N^��\�p��LHj�^L�ʜ�s�*�TN�	iWW����ެ��rl�=<���ǜ�W��1��;��֎J����W�`�0�b�y�E'�ɖ!^̈ʎ�i���ܰZs��i��T�ݩ�dvg��ϴ��Xz6��m7�|��'��uҨ��\R�3�O,��]!��ᙌ�\�d����c��Ou ������<��)��/���p�,71u�B2l�\�R��r�,���:�0�6t|����(S�~��[zVptq�)�<oՙن�N���RQ˫��o�����ѵ�N�1��8���˒��*\�#���Ƭ�55�θb#�!�9�q�*a���t,��jƳ�Ὦ*s\�.�2lDt��7���-cx��f�1��Df�]ąZgڳ�!�{��X�SC����퍦g�f��b�����>*������3ƅs��Ƈ�xE>�n�{�UYn�w�o_Nfw��ŀ:���ջ� �c�L��WהB��['B���}̜��;���NC+X��|N����5ۓ Z��IV���u�wwr=Xp<�D�)���K��o��؏3ˤ��k�W��c�7r2M�V�olv�袣;p�͸�Pٮ5z�y�8w9�ם8.�jz�pѣ�Q0�Z��Ri�[`2E�r�jP�]�.a�'Ӱ�mr�VH�����j@h�Ϊ��ԲVі#�(1�y_%�Oz��K�bU.��yl���X4��\�3���z�gs8�<�f��� �5.Z0�Z�cw\^�}�L��c0�E�
��g~�@Ou��1�ۈ��J�y��m{�C���\�;ד�ȼQ����>�~�m[���
���Q#�Bt.77��<�Gޗǩ��V]ʸ4�1�ҭ|�\�!��	����7��@��\�C> ��G�_�9�t㽬�N�n��W{NC�/���)�-ۯ����h��Vb��/���~7K����,����0nd�����8	ƥoNi�\:�i��(h�}��vGk�KJo�S=+�>6L��5{����f�
����Ƶ:̅�
����O��͈�����.�;&��]D�1m��zK�Zd�f3��8[<��P�p����y2�����B2���γ�s��oݧ��_0n�����j��ۏ9%�֟g��9�������%\ L��.��h��U�8;�`}��2.v��N��.P��4}#}:��i�Q,���V.�0ǡ��D>Y�x!$�z���즥 ��2�C����ua+ޫ�er{��w �ҙ(K�H�u&DH=������(�hvd�R�Ec�-n��Iʷ�-摸x�Y�]5�b����#��lt4ɕo)^w��ԯS��w2ı]7�!�%��m��t�1Y�Ḁ���i0�ۥQd��#+���U��bѤ��J���:�ܹ��w$ja���l��q��xv˭֝��w�	ݦc�|��q��;�;rX�Ԡ/x����L/����
��q� ��b��*��ԷyV�2��Q�AL��'��4�kja�e��xv�/1o$�GP��邡����s;@:D�Sm��ظ���`��v;����-�2���vҳ��0J���X|$�Ҫ�DڵWKa*N�K�x���g�5�W��h���;���𝻗�7�Z��#�&K(Zr�Fc\�Xm��3s���	��$�0QS���j'�d��tm��9���u�YG��j&�wn%�G��k��ɉ�YW[�j�Fe���8VG�opНe=QiV�-����}w�X�p3wb�ƴ�j�;��<V���y�]�Y�X�{���t��^9r�DnQ��a�3�Cg�ܻ��+�tf#C��]��Ⱦwȋ�jma�5h6#���&�Ÿ�8�m��߰�U��rdt���ą�n���W\7q�\��uǶ^�J��Z%H�'�\��9��}����Az�O�0{��.�:�vmSvٜ�.�sO�YspH�{��kOf%ccUv/u.�����>�!���n;R��;XF�L��q��t_e)!�e=����S݃f�=T��J�$q��H.������ �ϭ&��ۼ�7;$��: �5-��VM���7ϋ�����֓��9�$"��I�#PN8��Szf	RX�{��1(�e(�(^�$a� Zu���L����n	���V��ֹ�o =pp
*�	�Y�/U[�eAgH/4^6���̱�}���Iǘ}����:�{a]sK�,��GE���)ENU��6�W�cS��%��K�{,��
������A�WdF�JB�or�
̲]�)a���X���U;é�S��{v���q�xz��ě�f�&Gf��Y�>�U�N���-b���y�b��E�5Z��+ b�>���=֞g�2rCWMKP3m��H#p������4R��ͼ�p_1�p�im���f����7��k��M|�I$�^dV^�����C����,e��Z=���d�9��93~N#]Ps��|z|�u�Q|bGBǺ��]\�1B:c�wJ7���zӢ�A4c��v�U2B}�l�ϜgV�$C@�}s���S�ٺ�;�%�e�t�Z�}9���X��@`��y��!1'�׽-�0"-<ﳦ����u�����xn:��3��5���X��ˮ���s�9<sL�����8L����w�t��5���=wW>F����ޓ:��9^��V�����H%Z��#B�r��QH�)S(��<��Z���9��hh�r!��ִ$��Z�!J5P�-T虊��R���iQ��xkS)PM3wiX��J�ʢӞTC�q�'"�^z�-KVgE"��;�W���J�y�bә�f�T]��kwny��=E�k��h��T��뺭"<1Δz˪����'\ݹ�tѧ��N!����9	�橞C�w3�̽�s:gEK���=jb�iU;0�Ȫ'P�]4�2���	AdDk���G���k9�1�wt�**�HE�\�u��:{�UKʂ�A()PNNn��B2����]Kʊ՗���wJ�9�Bp��QA���Ri!W���Ks�4w[����]E2�J�(�5(/P�����"
��!�+�d,�9\�:��T'0ts<�"rJ"�S�G�MeAE&r�u%�hB�rI�T�QG0�5�Ȩ�\(�w�����˦�M�ܬ�-B�w2����"2B#�C�D�H#�?/�.s���ܝ;#W����_�-Rl�"`)2�������e8��7q'ٝV埅b��%�
����RAG-L�w-޹��N3��x�]�ǔ��>y�o��)�S�l���]ɿ��������ט��'�|���������9}��$���t�>_@��ZI�� !=�?B>��1��"
��*'���6�ծ�ξ�W� B(�$��A:�� #��k��>>�<�ô�?�y��>�������9��@�B����{O�0|q�����:���yq��ӓ{:w�!��Dp�o�Џ� #��s�n��34�{a,,��}"4Dp��Y��u�X�]�����w���S!'?{���&�Bt�+�z���Sr�:���9����N����?'?]�~weۓ~B�o!��Į�x�����۹���{��>����ݶ��",}$G�#H�:����ɿ�w���ߺ)�\~O��ߐ��<}�����=>s�����<�N���~���SHN�C��o
�M&����_����#�x�;y@��.�ߏ����E����컯U`c�>����P}�W���n?!��{+nC�i����;y������<~�ϗxL/���ǌ�����G������~OE�׀�$��~��Ǘ~w�9>��O~�_����m^����V���/�`�A�?x�HyL/�����U��HS�A�4�'�nO�A�	i��=��}B;{?�|�^�prS^��|o.'��0��ｷ���w*o�pxW�q�\ ^"+���@�=���t3�C�|D�'�����I���'!������?������0�o����i�L/��{���[r�~NM����C�����q|�<x I�!'����_��x�" ������g}���=�v������rs����ߟ�.�o^~~��i�U����󴇎��7>�z������&�O^?��]�7��^�~��®�P{O	��&��~���!�(Ddq�A|G�Aɿe���Q�<1_�Z�|��D|DA�nW�`����}����ad�v��ɹ�I�?~������v�z�{C�s�������xM!>��'>��}��SO�����yL.�>�>1�>��C4>΄���d7{����~��M��w?�v�C߿�~C������;ӿ!����~�yL*��>o�}x�zL/�=o�=�Į�M;y�~���&���v�g�7�<!�5Ĉ����#�"��G�-OE^��j�d�lV尺%�+`��̫��F\Ω�f:����Ԩ�CP�zd��=�6�H�m�1�o$#���+uχ�:���l'kr�i�7�ʣ*�wp}��ujo����ut�w�k�գ��ԟN����+p`�)T
)d� *�ة�b��W=+���89h~?�ǈ���a}����H}w+���ܘ_�=��ߞ������w�>��9>����_}������r�������]�|��O�s��}����>a��D���g�H�y@eY׾������O���X?�
\{M�!�y�ɽ|�yޮL}C�����7��|}v��|�c�]������c�|d����|�4l*�=#0ז������}C����NM���⌾]�';�xO>m��NӼy������HI�Տ����ӏ;��	��O�=w�����?&�){��;~g{v����i��!">E�u~��ؽ\o�[�������?z����1!�4��{���0���97�ù7à��&�~'*a~�,��G����	$<�����w��_g���^>��~C�L} xW�-��r�}Ƨ�����mn��\zW&�~���O}M?�ǿ��zM!!������&<�������x�!�*	ӏ���ގw�i$>����_����>�8��yǤ9�\|bG��������&�˳��b�}�<S���ܟ��|�P����!�>���߭���������
xM�	<�����oI�!:O_�v<��&��o|xq�'��>�����C�s��ԅ�|E}iW,�&l��ٟ����������on������zw>��>8��}����S��t{y7��s��~��&����~�<3���>����ǤI�ϯ�|o.��Mɤ/_�x�P�b>#�[�k�?nU�I����BIG�����O��ǏPrn@���v����>�X�������zղ����ILxF>�#��c�6�����*���7�ü!���S||�}�'���Y�ޛu��{��v��]*��~��xC�$����_���r|w��<��ϫx������}C�*�	�yv>��?&���E�&����?��8|�$�P��c�7�;����}c�>�(G�J=��-�w�^�}����]��I.���>_��v?''�O;�F���?��'���]��z���?��OV?;���q���q �������$�м�|u`�����#�NPb�
��:O�!���ힺ坒fg�3�����s��n:׵�u~������9#�4j����/J�v!J��y�'J#v��"�!X������[Y��䉔��k�<q�ځ6 ����o���&J�,L2n��X�س��G!cNo5Z�O����.�����<�������>|SH{C�s��}��];H~������w�	�!|��OaׇۂC������O)��_G�ϔ߾A��+�� ��D@�|��5g�V����'�0�yC�����n= ~Iǽ�<;ÿ�ɹ4����v��]���~���P�_���ؓ�I��B����w�C��<���㷷�^;�)��>��#�(`� ��!��c�B��c#��]�j����������w�k�o��xOG�W!���<���0��{>}������ I{߾�������'��߀���¨y?~��S��� ~��9T=�ǌDDp����Xf_�����gcט[]�O��}B ��#�b*�Dp�ϫþ;^on}�����C�����H>�yT¨��w��I�<8��y�?@xC���?|���yL.�":'���"8DH��<��^�4�aɚ]�3u��`�¾#�*��*����W�2k��o�׋
ԓzO��y}�ro�O�pxq�_�����q>�����yC�i�>�;���EӴ��c�^?}�� |��1���A���F�;=52�7}w�Ԍ��0}DBG�>��b%0���{M<���9�8���I��~-�0�����>>\rԝ��xw��nq��xC÷�J�'&�!@���<>�Y���| ��Z��o���އy]����"D�!�h��LE���$������7�'����I��pH|��᝼}��|[������=/)�\��;�a~���C�}H�S>�`����"}���1����2>[���c�A�H�H-~G�=!ɿ{����������޸�����m�~�H��@c��F~M�����ӵ����:���ӧ��z����$�<��yT©��߿g窊�v�Ǧ=t�mr^��C�(}>�o���������|���'���ȧ�rS����~<
�����C��߼��$x?�~��&�����s�ۓ~O[�q�Ӵ��	�u��xt������7����ؗ[��DH�!�?o�<���.�zy7�/�?8�} I��A�}�����!��~����7����}e7��o������*��'<��yL/�oA��x<����"!�=kj������%��� b�V���R��b�����0����1�on8��/�[�Ǻ�r�v��	aо�.��8ۗ�x�'9Ȟ�|��$2�=��/$z6�v�׽W�;SG�S8�hK5�j�.'zZU!;ic/r��ʢ���}��L>��~�{}&�~:���һ�r���<�s�?;w��sﭾ��]�3�>�q�&���}������7�|������O_��o�n�z;������1�=؃�QX"'3��ڱ䲎�/i0����_?���;�a"�d>��9��'�;�'��<��9L/�=���O�{C��u�?P����d""�"<>�����)�؏S�P�տ�5�@�:��-]�r��(�̘`�n�lb� #:��TLk<P�.u�7�ݿ��J\�!�*o'SCH�kN���P���2:��f͔W�.Z#���"�u륊�ŮWP�fö'*�Qq�0L7
�;6nTGU`�K%mb0D�,���Ũ�v�w3���F���ݤ&�|4��i�u�3��t�f)�(�㐝V���ٯ���Z��|B�/u��]�Ӯ�pT��c0��.pP���f������<�R���)U��]�p�I�;�%��J��K�;`V؆����t�D{Bc��y�1 �iں��|�|�/��/%��lK��L�_s����=���*�j��<��;>Ƈ�f�l�hln�/��ke�u��b�ɳ��z]q�����ݵڭ:�Q���^������I~�
	}��u���uJKm�&Bϸ�[����Tp��ˁv��݅-\�]��݂��:	Yĩ'��X��kVrqh<�i/��sݧ�w��ܛ�۝��k��@|�a�_mA�J��-��W-|��p�i�k&Ѽ���z����N�#T5.ޝ�a����F������l���`0�cA�M�@���Ҵ�ܶ�<Y;��ft�Vc���
�Aΐ��Ga�ƊF��\j�����͹�u�,w�����oT�eGx�/��2ep���8�ltk��㌽5��걑T�ÛV���k!>q]���M��pS9�x�R��x(4�|���t޹�F�gR���O�%�5ǲ�q�_������;C�6��K|�֤8�0m��7+��z��]��w�'�vṻ��{�/�n��p%�6 iy tڰ/�����jԤM�y{X͊�vծ��R��Hk��m���Du��|��*-�+�$O:,�8|�7y]ڷ(d����Ґ�}�m�/���V����`3h�=+(���OGD��]�6w5x� ߝ�<*������:Aё�H�&��l��z
�j����Y���g��F�8�U���jy˾�6�����|���J:ۖ��8�1C���u��<'Ð��,��۝W,�g�͂�����������2�vbJ�,цC����r���bnR��P��q��qVy��g>UynfEQ��
\�P����:� ��{�#h�N1���űb�]�[kCtgahէ�DP��q�����fS�vv�BGf䋖��:��A����z����z�\ ��a�^^㶵�o�P���?��2�I�޿�F��U4�z�������G�_#��*BǺ���Ceg��g�{\�^��@���x7{'H�Z�s �;�u�� >|�̸@������8j�dW�܁����4�Y�J�����`�+��!Y��{�g�<Y�B�1�ī[I�ߠ\��G��lOg`��e�;��L譭(�0���� ���N��#��iW3�cY�F��R����+�ct�x���'�K{�3R"�2§��fI�O��=%�y�}QW�����i{O]w:bj3i���KG0�+��;�.'��$��J�41l*i�3��& Fi骤��-�C~���pr��2K;qvַ�g��%��؝Fs;\��u��K���*��1�U��}�˹����q��6���a��gf�bQ�{�e��2�1ۿ:�M��jO �LBR���qR�`�Hb{�l�Jz������K�����9�#����=r�z�#�d\]�U��C�sԵ��8�z����g�Z�Dp������<<Fٽ)��Dœ�|J%X�)$U3q,�(�mW��1�o�������
ɬ����/Ry֣!��Y����揷-��R'x�� wOt|�����2�*i��1�E2	|�����Q��#ᏻ��}��q#�\�b��a����Ī(-�y�pC>s9�c�"b��r@�Ƕ���.�����!�0���&b�a\����s��7�ʮ���JR�І!���Ef�v�Dt����@K�H�}7_e}rɉ��+���i�6�1"��[39��M9�[���[fFt�,`��%c5���T�@r�H|ϱ�W�^Ş�j6{m�٠-y���C�0Ȅ+��#2-�,@�:a,v�M��B͗�q�c�������Y��~�FǾ9M���ͯ�2Y��� ��=�����/�&lD`��՘�澻x�u�rb��N[�GU��4��f�A��w��dө�cs'�o(�jI1�E��k`�f�Z��!9u�/&�*�b��9���6�\D�{O�=�"���]�m�����jպ3�ƒ�z��2� *�}J�"���ү����{8P���Ӻ��j^���s�>�C�w��?���ޛj!�R,�����~�CyU�j^"puDk�߸R��{	�ڈ���Z&���f�辶g'�g�fw�	�n�R�	��옧�Q|��B�8�p��έv֤��UԻ�$����T�lWw�s��YR�!O�p�Ϯlc���:���7{��N6\���ZhM.��P�Ӊ��J�+��c(~����|�;�vF�Cq��9T�c>��W�:��F̔���?X���{#=IS�Q��~�(�r����X/�ڰo���ϝ�-U��X������
W��h�G��qכ�"sܤ���J�}�< �Ǿ\������Di��ӌ�Ӟ�6ǻ
�as�J��W�����rqU!��p�_E��T%Hp��S��d8�l��Į�k�;G:��W�}:p��t�-��ﺅtXP���dI:Σ�L1w��Rο��Lk<��W�^h�%�؏n�w1zn]����D�g��E�.1້,���!�:���ytnl�if�A�N��={��m&*�r�7��tC��T�>C�e�au<'�񙆼3
�图[�=+�;:8znӡ�x[f���u疄�e u7���;"L������YhQ��ǯ�Έ͵��V��xR*���;�0�<8s�j�h�	�b(tM	������v��+=-r�zM������:�~N���zL��J�����`�TL�ߛ����6I�ى�"�v׬dhg�9��E�G�b��,�Gy^���{�S2.ԣ���è�K7�J���s	��h !�Z�����7!o�7s�Aw�y!���9��.�%Z����Љn���wY��̟S;�'Gf���q�ͦ�v��#����)tY=� ��>����}��� x��r��qh�Fŏ?���:�,��m_o[�c�DW�u:��D=�����o��~/�ُ��տT�d�an��-ҷ\ ��o�狀_	{���W{�o7Np��t�x9;�@ݘ�n��M��Z+��8t��]iʛG��?\���O�Hh��D}�����H� >sh��u�&Y|#6���IE l���K������=䅿^��
�n�θS�p��K�BP���ن;3�_n�nP�q���l�b����u�&{iR�=K=���N��n��i�2ƣq�4:�\貆k��Ct���ޔ<}�燒��:�l"��eD�̷�V� Q!�2����E���f-W�)��G��r���T�"z�I�ń1u�&�,��ɍ��)Y@왇�]I�O˦�d"��S"�=��p���F&�R���v)����#[����>�6N�۔����kG��]�-%]���:Uw�{d��3G)�5�����99S!�f���"&F��Eba������{L��V����Cw7	�7
�]7���!t�����K�»^6D�td뤥���],t�����_��1��� �`1��y#e640f�]�������;�]#����a�K�����F���߶�F�j�^h۲��ט��{c[�N��tj��{c���磌�Ӟ���c!��}!��Y����h=��ƈ�wDW���$\)��R
�w���ߞ>ס�sȻW�p��H^��}M�18���/(�o.*-�A�)���w/�6�c[U�FҊ�m#�x�Ƚ嬩���*B]o1���*z�Ach�#�ca�9��q�H�,�����Y�1�Px*���5�xW�J��M��,}���.�=P������GG�5�n%�G�韮b����#������6��}�q�9���2fx�����i
U�����t��y�9>X�ϯ������@�wSͷYr�W٥K���f/y�0.T4ͳ"��Di�.@�2�Z�x��m�>�:܏;5u��������Ѫ���`�y=�޿��ݎ���6=6�m/���$Qy�y^��FR���UꙵNP~D����V��̼*�����OM%t0foٽŧ��g�b�hi�YOnį��Y8�����LHZ[?l&�����ŕ&M�� ���Y��y��]���*шf�|F��sv����=�Yv~a̶�N�f���r���Uzs�4�6��kN�w,�ք�.��u%yl�hJX�r"��(྇"Ɇ6F��Ne�OWb3&T��f��6�ۚ`��d�S�{2v1mԀG�/8rz�+��Wn	�Kf󬒻Xqc�����ڱ��f��YL˳p��V�ewMu�+��.�ON��)-$�$h��*�һu�L��nT���-o5�	�%
�Yo�5I/叩a�'v��y���rJ�_7v���L���ۘ�Kˋ ]�A�Գ�u��e��7��^Ǯ��\o��s��i������K��2�-�.���|�{V@Ƴ���8�Z��NF�hp�4����.�P�-ѕ��
�:�U��f�<fW�v����� �b�3���,'g>�3�Y��^IYq;qc9b���D���A{wa}�E��*eܤ�X�/4�-+y�hItaf�=�c�wP�׽@����Au�,|_b@\�˚�n}��:<��7:�+�ʎװ���J��/Nbn��ͽ���D�7�X��e�G�!�qeZMv���<�}�K$m�Ϩ��7�DYZF
�a�JVťԹûqu4)��[�i)�X��XOo���2G8YRc&��_p�I�y�Tq|8]3�77�R*�8������k�R��=��=�+�i�q¬С����*������w�e����N�e�5���R�d��^1-��I[�p���%�{-�t�W]��b�>�a6ɱkS��J�*	���EK#n��WY�P���b� ��es�/��/Yp��.��f���X�V�
,۾j��y1��YJ�,�F]a����T�׉���mL��k^��E,4��D��uL��^����Y]5���}]*A��J[0<�[�v�=:���YzK�KaT�f��9�u�a_V��۔U�E"��5Wn�>�
�zJǝ��VƘ�Hœ
b�5�t��8�*Wח�^|$]W��!��,+ʒWo.�++{�F(�6.>Q��&i�(RҲ]��K�q�LĐ$���=!>X*ڼG3M�;f8�H���Odz^��Ǫ F�gvAS��K����qM��S�L�=���:V&6���;*�w40��#���*�#6���\�X?^��w�T�9��v\���虮n�e@��%٨�W{3?�y�@���H���I~��a���?�ڻ/VAv:��۸�'�[7N�u6�R���E��N(�<�y6�N�XY��h�W:1Xaq&�7��[*��;��>L^:����Gɧh�L���V�خ�z�W;Luũ��G'VcSXe)w�*��+�M����;����h�����zM�g����ֶ�LQm�b.���}��m��K';Wr�XH��e�;�͝��Fa���+î�u�XQAQ����别2���&��D�"	ZA�=�:Hh�Q!�d���vPQ���uc���Ȃ����R�Rq��D��exaEĐ�4<R"���S3%RL�TT������"�W9��9܈��9D;���P���qӮ:ub�Y����9Ą���$R��D����IeQ*��#����t��e9�(uayzJ܇'S��<��S�-�H�OBJYR�YD����'GR�2Ql��5��"���N*l�*�T�YT\���Ԝ����t؄YQ��VNU��P*ʠ���.(��$��,J����y�D��E��\#��Iʊҵ٢EJ�iaWC�=k=��֕�����I�s'"ʬ�[�F���#�ݮ�RmP�ܼ�x���I;��ܝ�B�������e�E�x�=u���C��u�ō��WA�|��; ��%�ں*i�8"�F�À��|Ʃ�r�䠜u]��t8ᛣ�r�� >5폮.�-'��ך�d_��yVT���g��Mg�9�\J�����òVo������ض�Ua��Ҹ��(:�U��W�{�2V9��h[�����:2�]6fd���F��)����>��v����C7;�w)��bo��( ��� D��wy���|,���继\�V��4k�|~�ԝ�u99���Ӓ���m�f��E��탽�)���{�	:|�)ﮅ	>Bȅ�f��k���:X�ncDp��aW�<��N�Mݫ�f���	��vɆ�&�0a�]���W��NCN�h��C��-~U:g&�3��s��l�v[�w�����خ�<.:��Ȁשv����|MG���ڴz�����
A
��1s��Y��T���u�5,��T��Dۮ�oʟ����^^G��}�X}�7��H�����,C�Rw�]��� �$���>=�Vrϵ�g8���GgYS������V�r��۹
S2��`�n�uIgc��L!�>�Xv��#�����1ü����2mV�+ܻW�7�ɵG{��8ۘ#�Ô���b2Y��N�A����@ֳ� ES��7�ܷ��hմ_T�ye8�%w_Ϸ7r����W���"i(��#�{�NUɣ����{�����G[w2
r�w��}_}UI�~>c�ci���z�X��bx�*�I�5�W5���K�Ο�ys�2����S��c��1)���Y4�]�+uMs�.����x�NuJ�W����4�ޕJ�a�1�S��e�sR.�)��D*� .̥�^J�Z"�'f�O*�u|�ـ;��p�x�K�=E	�[;`��~kr��=�{r�����s���D\J�ŌgC�_��>܍e�%�0��aC6��U��D'x�����!��1��O�J��=u���>F.����V�M�a-��[XՅ\;M��qc��cT�7	�3��ЕZ�����@�_�f�`��o���S�4���_0���:�}�$w�B�uÄ�~Cp�7(EC���V�w�­�.�0�^M��wX��&"s*�~�8���..���f����j�H^�e�%5�-ZQQ@�W73{���q���^8�R,	qu�y@?����)����
���G��+�d�$ٯb���&zL�{G6껇Q��+�b�y��"��ϱg�NCp�}_}��^\�W����n�0e�Jde�7Ȭ^��/Y���-���r׈t����<�lf��c�w0�һq>x�s��6�)o.�T�����ǧw��)���h<d��S��S��I�|����*�x�Ǧ�R���(BQ��{�w?�ﾏ�37u��/����g���e�� ���"�,Ȉ�}!t� ,;lLLR�4���Τ��7G6����� n,]11�'�ئ-��fϗ�l< ]{� N��P�}�说�٩
[wR���xE����'B��� ��y�����o�j�:���W��#%l/̽V�����������s���k���x�5�i��O���`׽�����^ߜ�q��>��E)r�ϔ���D ���*_�;(e��3F�Q�X3����CU_B�]$���`uݼS����ʞ̚��1mC��m]tb�\p5�O��u	�'`���
S�ϭ�Y����T@�YH@��r|��z��>D�d��|��y�2�nj���]��!y
e]�3���{��m�w�+殸E���W%ؙ��f��<�훀��K�޼��9G����5z�pc+����O�u�w�yC����Y�tL/��F�~��^̾Y���8 _�o�SvWJ��ʙ�g)W��X,<)��(u1b������p��/8��-`��j;��=�8*tsz��З	�U�t6��"T%N�os�������4A|��A35q�<�C}Y���V)������7GU���O���=p窦&�u���7&�j ^s�m`�ƹ�C2w��8���n��| �=�P?M0S�t�^������g4���xT�n�1������C;�^�;�^����s� \�-}�o��X*{Թ�<�܍ו5\ �O�SC�D�S!��d��ؽQ�XԽ�g:G7�3~y�+�� ���!������@�-�<�>�֏I���ʞz��ԧ��6��u8�}��T�#��*�=2t��(�;f�f��\�j�����w�r�h��$����6��a��/+A��4E[�"*HϹ�e�h*���6�R��`8��	���8��V����p�9�f��Ϥ�����iaD�,y�{W�哴"|�5u�4���}_gW�������
�J�������
�TJ+-&,VNNy��ohO��^G��Z�u�*�`U��&�[18Pu�d�Oa�su�s��5/cVj��0��?T�� �����Z:Oݕ7f��N���q��ߨS층����C�J(<'���9�N�u!���N����;P���}�֗�"0x����?t��839�I�l�t����_i��cJ.]�;.�֤u�a͒[,����;u\֛����8���l�Q�����4$�4�B=xܜn�_/�:G�Q]�幺� MS5��PlK�����˸w�
jXN��٪���'u�6�,~�|>�h���;P����� W�%���u}Pp�˧�m΍0t�����<I�&��Y������C����OXT�����l�s�������2��c��=;+��9���e��/��,����H���ҭ,�Y�
V~�{������6�S1�[;}D��8o��r�{63�q��b����8?�K�Y���L��c�fIV����P��1l��
2�����{u�<m��k<i�*��U�L�`�x #�{Εg(��8A�C���X_ʕp�`�ʲ{�2ꉪ���@��+T���ֆ�Z�R���Ә~���ۇ��B�K���E7u_�7E 	H � ^Ϣ:���z+�=B1,i����* _�u�r�#����S	��!M��ddݹ3��90�9���'��Q��аG7S�qX�L���i��¢�N]�]��5��]:�D����!��/����<t�I������:�nb�Pr��vONfmt��h
��r��1W4�V�*����赜���FQ���>7��z�!l�L���e��.�0C#ebj�� ���
:y�M��iii����W ���֬��P�&	t����\���!�Jnlɒp(�*�ҥp���_}_U�������%���Sk�M=��D�"�����GB�+Ž�+��(	�/:����y�o8VĈA�����5!��1`L7_D�L�f_蜨[yZ>�rH�;[n$�0rMd��q�k��j�FK�ႛ�QZP�R�ST1�'?5#�T,v��p="�{vn�'�������~�7�CHT2���۹B��X�#��aGT�_�a��ydWF=�su���N�{O��F�G5����x�5� �u;�����1�S������Vw���{�]:Q�x9I!���4[�[��/
�Qx;2����>U[W�O�;���r���k��v-|��s����;�E/��ٔ�����TU�*-�1X�W�!��o+v2����JnA�͐O�:�	�X��8��<Ql�b��U�.�c:J�_e�c�P�ך֊k&D^⤋�0�c��N���^�z:�ȌA����<�od��{-��1�3&)�H�6OgQ�}QvS<�jwLh�U}q|����n��8�NMP��a�$��Pcg*uI"f�gd�MF뤬Ҏ٬Q@�K������L�~���l"M� [/v�z;����	4p��ԉ��Кp�0���q#5T�-�����˹`�{3+!OmE�.����G		��%������}��.w�q����Q�&� ĕ�xA�׵	�������B)�;Bq��U7����T�Ү�$����#�ר��M�����*��u�u��}ޜ�ds�Hb��wT*_:��J�O�nT#��_�C��H�%۪�A'��ߊ�b�#%Y���0�8Ѻ��SOOf�ɸ�:5�˝���ۃ(�L9tɎ��F�T��t;6J�w�c��`8��Q��k�;ݴ(9�c�g����7�B"Z���} =7��l1��yx�$Ÿ�S~�g�+��R�4������*ڶr
�b�R8 VP�~� �B�`ء����<2q� �i����Gג�+j5�D�:>}D�a'fͶ��|�(��B�a�K��vq���O`��o�o�E�)䡦f�҃��s�`3��G'6�SƳ�g�>�)�ر�T� *p��@����c0����TF��f���o!�:U���4߶ܷ�79�V�jS���}��p����2�V�t���C�Mj���B��{C��ub�	��d	R����p����{xU�f�Q�s�1n�ϲ{�������\[�NZ��V��MT�hM�Jt��٦�T�|ވ3	P0�E�E\��:���*:SU͉L��<�T��0e���6�ڳ3�J��X���Ad���	NW}��<E�mͳ������SKgy藨H6*����6��:��݉��h��.F;?PϬ����!1�z�V=�z�5`	v�^�g0+�S8��P��
pO�X��pay/oҎ�a�k���N��{�~�1�p8��Ι<�a�܆����7�G��Ӯ%����t�]ε�",8&ł�*����:~�T��Mp�����YN���9[�7�_F��8�o!�g����Qh�O>k4�%�B0�⯹@�L��)m�Ƚ�E%9ͨ��fA=�0�-��?\u�!�K�Ǥ���?T� Mg�m!��d65��m��](M�{~�s�ޫ�P��2ի�8�U�}��^ET�+�J�0"�X�WN�.��D���ފ�2�z���	��qn
9JdStɮ�
�]T�D�xT��u�缋��K�^O�/��������V����K�"4��#��8�x��-���+:���z���B-���Q���t���M_���.OD��8�Q[R��];�Hs�-k�:^I�77�{	����L]�d�K};�2v��\��	\k�^�i]��%�<wsZ�����ӄk��W%�����rw]^�a�#��RhƟ[.��\o��m�U%���S���}V�������۞�VsZ#�����!q˛�"�#>v��ey�8�YBXrg�(/)����Ev�ՕͥTgbkE����P{@L'o��6��u�-ՎEሱ�ǃ�����ք�tƍ�ݮ������+�j�1p�bø(�*!�'�ܹh�X��B"���1n��޿,���ģ�[����eLhш�A��2-��'�5�1�<���#�J^cNE���>�D��Y�9��54S���ݡ����c�f>�L�qʪ���m��,cBN�a	�asv�.���kZ�6�Y�r�Z5KY�!�X�b�xkV���n����_ �_\Qضw�4�
z`��EvKD �����ٱ��*��VN9���A���1ͅGS˚k�l[Dt���I��m��Uv�:|*
�;���us���o&_�1#Q�խ?�]<���ZT�{jgO���qM=*'��-��Q}��!���U��M��mP��w���0ڑ6ni�e��r�[z��:X�=�H�D;�9MWG��1��
R.��U�CSn��[���_^��C�c�次|%��i��,��h[�,kB��(Ҙ�h��8պɆe�V��Y���^.4Yiw��Uݔ�)7���6t���3��N�� Ԝ����RuZ�z+ͽ;Ff޴���uqV
�˖�sk�ݸ�_� �_�u<�/k���w���!q����Q��K���cʆ,�U� .�F���ۣ{��z�r�@F��,-���	�}��NR*5���b�*���s�n�$㹋[ȅ�F8� j6`�;*����5(W��^����=���eW��EpMa�[j�^��X^㙽��{Yy��YΩ�a0���WH�=f8BR�����\*"g.ڷ��u�r*�68���ߧ���r~D	KjR=�1?d�Rɉ�[Q#c1;���}:���ݚQ�e���Tl}���W��R(�h��T�}���o�rպ�o	��Tq���������iˎ�v�K���CoX�.8�)�@>�5C�lP
��g�B׆��E{�iq�u=qz>��|��nǵשphi
�ОO�.%�y����	�k�&�ժyu����ps���$?D�C�H�/o+�'kf���3Q� �S�x�kY�3��.}=�����o�}��n��9޼�l��$Ն=CE�V�\��\����3�}��S��ߨ>ͱ;n��Ko�5+��A�o�Y�iC�����LF����U�vRy�N��
��Y{Cky���F�3�[Ӫ��I'nf���d_4�a���Z�6�ԫ�e0U���ө˻��W%��$w8>�⮧l�m��\(&�]��}�:{�r0�mK�Z
|Ojt�űJ����9K3~F���y+Ň.�r�\���x2�[S*־�l�SX���%�f�g�����0-�I5�Y1R2�cU]L(����Yŕst���&��X��tK{�����evqy�#x����H�ٰ�tr����6,U�<Ų�]�s�y�n/]���C%�fE��j� ����r�N�����+�3�G�gV��u�I�S̔��ǚ��\�J�����"<�
c�V�畄��q�\�;V����� �����x���(�V���i|�K/PQ��av�ҍ
���nͻ@UHl���j��r�+pD꩎�VP%IK��H��Xz�r�����N+��]��G:� �1���Pv�e�r�[�N�{��1��]f�h�	�0e��sjP�i�rn>�!U��w��Ѱftw+&�%E�$:��u��d|�>���ֻ��F^W��WX�Ȳ9����K:���S������U/�@��@ť\b�e��(�h�����x�c�\��.9��j��=�]��݅�n��dFi�2"��ہ��{��:^.��Td�S��U���IJ��_b���c#�<Ȏ
ĉGY�r�땱bXS�ÉV=�N���,E���*�z���ݱYcrc;�x��u�/( v���	,`�X��J&��kZ�w�!����!��P��~wJ���7���{��������+��$N�#|���; �ڊM�&@���Ω5mxk5�k�^�LM����.-�6`t#��`�k��0��cd�Z���N��NT�T�nT4mu�gl�5���q�mҌ-ᕈ��_vt����,��;�C7�K�ݭVf�Y�@�3Mծ�>bhf�[�8U�u����ԩ��8�]Ŭޛ�Nڨ�0�Z��E�kkn�r
]��{y�ʃb�K0R�;[8�$�{�5e��c��*Ɂ�AR�Cn� �m��nae�
�vӚ��x�/[�T������'�c��쬬B�cw����!k�[��Z�09���fr��Eo�e1m�9��O1.�G/�t���=E��W��r!��v�va|�[��D�jf��;�B!"U���b�WY{��TcG�vX��j��}����U(���*f�Y@u;gkeL�w!"a���BI���,��V����IĐද���Ɩ@����C��2��+��r��*�屲j��.�w�m=�\�ۻ��y�@��#��Nr��Lv3;���}v�,��Aj'��N��TCY2���Ύ��MG�绮w��uK
���i��F�.DZ䇄�#�9��7��#��t4�7!��В2�{��"�wTu���=�C�#RC���u�I����]ʂ�Ը�TQ�L��"D�r��dng��f��.�	E�U%J��9���)#��i�ʄ�Y楗L�6�I9��T��*��wW����(�"̩RPH:���%�-,��Q�d��J��e$��4���Z:��ZQ�eBEJC�^��,�t����(�"I!C'@�e�,Sd�X��+B�����H�Lȋ����FwX�)U�Ae�Ib.�u�p�C'O�BBSB�JXT*E,��)�YUY��Mb�j�EJ�r's��.�RWP�F�V���TJ�ʫ3�rMRTMʫ+(��0�B�������s�$�(�$�ь�8Gn���3��Ox���㌜����Lټ���kjwhڦ#$n��GV���45rS�V`毹��#�磌���f���g�^��@�J�7�"����5 n��r^ʥ\"���/ʘU������N_j�%N�R���[#����.���r�5u�{��1�V��#jf9���:��n��:���WL��v�vA|@��DS�;U�s[�Cr!�`ێyh��+�.��T��	ɻ��r�(���M����C� ߎg\�U;w�;<��A����!���#��e�e���饭p�+�@fK�,	���&��+ Ą���D������nX���搸&���[�ִ-���q��@E
��e�Hu��B�ﰡ�
X�5���U��zoDdX�@<����h	��|a`r��.;�])D���$�'�x��j��m:��Gʗk���K~�1������F�H�SrɅxEz"�]�B�L��x4��2�r��*���C����],EGȼ:
n��e��D�q/�ɐ��l��EQ���^ًF�<{n5�3,L1�s�}4�y(A(������Р�uA��j�Y�t������j7r����mt>�2�� B�8I�v�Ē2)`;3P��d"�I�����vI��>�5mw%*)ûs���H�S^����+ػ~}7U-bbv���w�$�v+�U��[��6�]���cI��lbPNf.n�k�U���5���ڔY���!����+e��W������>�+��׎4�){�?!��.35��<ǠT�nm�q��>��a�Hj�tdА�0T�u�[Y xkv��B�C6l��3o��Sڅ���(:�����t�f3q��b�x,:��V�Y��Z� <�M@� u��r��k�CuLZ|C�ʭ�O��ʻ��nټm��N������\'.vZ21��u	��V|h�;u�!������s7��y�h9�me� �ֈ.2t	(S V��bRFt=��E7��_�h����f����Bh�&=�~�TҜ��tr��Vo��{,z�
�1O%���:��BU�_*��p�x�c�2���Y{Ys�(�$Կ��U���E��k�.# 1x��%�7��W�ܡ�^����S�7�6W��L5g�kv��%�
uP����,'O�f)��Ub�Br�\s��YT���%���]k��Jvl����� �¯�&}�޴㚍٩C�{KH�Z�ֻ�{���q�m���S\���am��GeD�2�Oկ�K~�۲aԴ)Od�	*ɖ��Sm�+��6ժ�����q��f'm��6Z����[��v���n�����v��y�B��t��;
�4>�^���޻8i��_�EE��V��U�l������,��b�B���[��NM�FKo�����������~�~׺�&ۍ��q���za*�	T��:��|p�9�Iv��v���;Z�r�鯔��n;�㌘�H��ܲ�`H�sl���6�j�hp�/��s�C뮌M_t�n9��b�v2���щ�}*���3�}qW��.������|��S�75&a(������3�J�P�V�<+D���X΋y'��s/��vI�鮠�^Xa����e[����� �X����6����3����f����X{���
����^6�p�O`,�:���h�y��H[W�'%�4�;4t�^��O�L��+�.�➣��8T+�_��U��[
����}���36������5�j��S�z����7�V�g'�t�V�z�'\��>��7ud\�o1F:�Te���������EPx*z��W���P�ښ��Kky�0f��X�sYՍg�Ph��Ig����xwv9,������x�ck����|k�L���/j��iw���uL];��QXy]��y%C?6M��5�.��-e5��;��՜��������/�?L�r�p^t�./:�\�ⱎ�Z_F����-}<E6�i�ɱHr�R^�r�oS�)����v6�����UqTY|���(3Mc��'o6���Ng�{��ˆ3�y�*�w��u��L��0:��J׳�P�8>���9��]Z��{r
��(;p����$zO{͋�t=S�.w��s�sK=�}��7[z���Y-����c�1����q�Rx'��A��I�����cw4���R^�y�g�zC���}WS����n>���>�W�5k�쩧_�Ӌ��L��v�*���Eߙ��B�\�ypfXL �9,}W�	}hiť*L=a5�S�H��p���Ɋ`ĭɣ�;��>J&[��l��:�a�7��5����&�3�٦�4��1���wܡ8g�q�U�=>��;�������Vsg=�_�a��v���9�}!�f�|is
ݨ��
���o�^����<6v*�Z�:
��θ��ή!V�BTa�mV�x�(�Z���x�W��n���<J.����%sv���tV:��U��W=�p�x`uF��#�������`��>��5���ޠ�51O������@0�!J�4��>}4��0_>��!G��q`3��o]�]%��j>nY��u�r�¬Y����H�N3��e��}�y���r�x�Q=-�6⮦�8�y,/[H����|��ާ����O�m���+�z��أ�/m;,P����!���w��I�^�f�y�[�V����8qv�=�і���F�H��~J��;�e6/�Or��M_k��0-Cr�xۇ��īӝ�����]%��c�ꞌ���K��k�=�<�z+��γ����ʎ�y�����"%ʃ�n�����ڥTO0�S{*{��彭)sZl��K�s��=����O��+�N�>q�_c��ay�l[�7�.��٤����B���Ȓ�\2����򷲦���[[KM\x	��瞍ʹ�'`~G���Ğ�n�y_���(W�T��A�������w�T�z�]3��վZ�u�s��ڸ�.�.���c�T�B���*L�3ch����R{L��F�\ٕ����؇H#��9'kx�o����}�V֜����s��tg���X���$L��/�	޹��v�q����oc�O\fN�m�Sy�c��(�U�j�F�<V�ӄ�LK�y6�L��~^�6�d��H����7��m��:��V�dR�b��������!4F� �$�}�
��ϏM�3(s��j��&j
��n��Ժ����n+��w�v;��A�2��Y_Z��y���P�PڇΪw]�m��ԓ�����etSq0��_`�}y�����¥��n�v�����[����1��S[Y�)��X@WQ�Ѯ��w׏j5�--ųf[7b�9�MC�ʷz�����w3���|�9�d[�ܮ6�v��E��ժ�W�������y�C~��I����!������:Գ�e�$��{��4�&�8Ǯ.�GG]<y�}����=��Wc�ŝ~7Ղ�)-5�J[��u�ܾ"�X���Vgz���PC=^��N눿Cqy]s��0���o]�7ܪ̈́U�fQ����:�q�Y�if�>��s�Etq�]�S1�A�4)���OSq�]���u�9䈙��*��Ņ8w�}�}G��ަ����+��:�Jnq��j5(�sb����v����mkbb�r���>���d��aw�@��Xų�pT��r����.7=y���[�oiMv_��}obU|k��J��O���w����������S��:�G���zO.Ȇ�\��H�����Eĥ���
��`�!j�-�Ng�������z3I�L7M�	_�a*�бLUM#;�՜ؽ6�S���	%��O%�q�6�=!�s��}�2�r�s.Qڵ����^�3O/V��_T��D����@]�q��B��:��y����܀��'n�%|�;:WN�Aq�Ca��&"�Z���ˊc��S��^Ǿ�el��"�ax����ŗ��zt�8��wu����ie[��iw�7ǵɋ��\^��H�i�p��U����W��jY�}�m"�3�/���d�|�-.-���-љ�{��v�X�f��L�ٌ������rL�c���$-���\���,Uz��A����S����ɔ=�Iy�М1#����/����Ә	��0\�:/7_�������w��p�NԻT�/"�چ�L۸��	��,�����P޼	�*�K�����gmk�f19�����K��z����;��]|���}�'TO޸9�Ou:[:�|�Z�|���mr��/a޹�5�C7;��u�Ӌxl���G
q��*;(㺈�ɿb�Լ���:�;ɒ��ؼS�ݞC���.sz��ս�ܭ�=EC�p�����]K��$0vt`�>��(cR�>�L������=�ϏXt�n��S��7���r�^�5N�WQ�F�w0�Ա��ֺx��ʈn;�lJ�[Ƴ�*{��O໺1?�O��������5�^Ǽ�S���Ujn:�m��JH7z�����N���BN%A�':&)�W+�!$��i\8}�o��N�,�0Uf�fs��`Ak��Ga%í5���_l��4�5�r���)�7]��b�d�Xwѻ��m�K���3��v^��2lq`�+칞b���$�|73�N�K�0 J���D�euI��;�޾Hk[wݰ�#Q�9�Ln�N���܅�HY���
[N��ꖄ*�S�	���K�nJ�<�� ��Գ�Ƕ-�o*:�y!H���U9a�p9��\�L�jG޾WƳ.Қ;9*"zc>j���.�k��SN�qⵘk�V�Z���o�a�n�\�}�Ok]�=*��u���݈�LD���!^E1p���}{O,Z9ɗo�n u���9�u�C�]�}*��KY}ffA���E(�M!y�Ҫ�,O���)a�ŎkVLoPU���mC�M=��
̛4�7_gn��̾�����z�3C|��^Ҽ+
�w��	���==B�ݸl#e4�[�n�J(ۈW����/�o�ʼ�W�����u7u�Y�i�n6�2����;P�*[�x�ʂ㲠�z�������ő�"�q�j�/T×��i<hq�ފaf�N�\��"���{��ݼ�%�r�7��c����OX�h���Gͮ��^���>䯙�M��<x�K|�i�椙R�/i]����0� �i��Tԅ;�B�ް5Wh�z_x���^���919�U�:�^d��%�On�� k'?��F�ܲ��s��L���o;�z h�(��ճ��׋A�k}���^��%�:�г��U���庁S�磌����5u��������߭�:�71�Ӽj܍{�������{�I�c�,��xW�K�|'����u����*��ީQ�ަ��OX����������ß���`&;lT�|*�%}���>u5�Q���չ�-�o�w9��`�8��V�U�U
:�$�=���=Ȯ�7�;ӋOV&zp�:T�������qmJZ)q��а��3���#���;��H^Vk�醱*������x�)�9]2�5"9,::�9`GQ�YL���aa�]����%�(�}�y���Un��JQ�;XZ(��nl������b6P���p?One��!Vw0�5n-2F�j�k�*�oY�h���7�����ʈ�vŏaV}�ARLU��ȿ�D����_>��[�1?�nq-1�pi�ٵ����zq`9�����4���������u�Y�)�[�WhU>D�ҕʌq:�jO.�a���@h��Ṇ����<��O�hۭV��oC΂�*W
5��Ĥ�cc�9�"H�a�ց�*q�I 4w��w\$ jw����]�R�(�ȝН��+��a��~�����`U�̢5��v��d��ȷXJٗm�,6����}�͝d7���I��"2�Y��K����<��]ήI��i�3�e����`�(���%7y['7F��
� ���Ϥ�M�ª��H��[�KqwI�N��ͨ�qUۛ��'�Zׅ���Lj�	�N^���+㻀�n�Y�����HcŤ��EZ�n�����cy���`}�U�q��eh�f�U����5�F<Jѥ���Z��݉���4�����\�e�9@��Ec�ʾU��o����ri�I�;��C�Nk}K��$jfvi+P�Gh��,^u]˭���㸥Z#��_��ţ]%�*4I�Ճ&d��e*#f�X�X�!\����p���!c��f��2t4<�]��g	��+[��e,��}EI�RUc!FF��ާ��ͼ����'v¦q�f��L�-dA��2V�x�a�w��Yy�j��'s�f��,��ĩ�}I�y��ʽ5�.�LE�M���3�����7a�jԪ�H�%���H����P���㵹i��?���\�������Sj ��"�իb���S{y�Y�_^��(R ��)@s��2S����E�W���T�w�Q5U��ֻDGV��\�Kneq�(�A\{$�ޯ���L�*�ˡ�e��=s�5y��\&������ԛ�|��;]+]�(�nA��-3�ǭc��s,ƫ:�ƘĹ��tl
�L���Ѓm��R�d����L;z���u��U�I�$G[��^�u���J�V�J��+:L��,���]�N)q�@&@yְ���l�YQ���61��oi��f��t��}6�2�0l�H��^o�< $�k�Iˮ�]�VTۦ5�{u�Mิ}�J':����쫁��L��:����`ײd�p�S�<3n�1�A�Eͣ���U�r�7k�.$��������0��g,f3�
��,(���M�{��pS6���n�H�Hvf虭�r�ふ�;��Y����>��	YP"{���
�6�ž���e�k���p�;M����I"/{;8��w)xx��E\�P�t���,�M��X���qr�����N�l<&�X7�V���M��IV��z��_,�=�C���!}Ft��4�s���zB�0�:2 ��2 �U�����UxQ� A��7�}Q엇�蘮_nΕ�.�sy4��.����Yi�338O��6��e\�0�
Ci�b����(�2���pջn�������]���E�����ܵj�ľ;�`��W���<�S���_t�w��g�����v���j�\`˂dv�+s�ZW;E`�Ƙ.��k4��\m�id�U�Z���Wػ�r�}�_��z���)^zE�u,4�6-��b���Ј�Q2�\��م](�,52֖��LBʬؖQ��(���MZ�e�IeeV��I&qD��#֓��d�V�deUis)6s%�r�]���h[L"�32��0�H*d�bI�£��F�Q"JDTh]l�MG$����YI%h�0��R�����T�!!FfRWZI��(D��r4���%JCN��ԣ0�ԮefiH��FEbZ!��X%��Zde*�:�DHA(e��笔�l�B�6Y-8f�T��ˑ��AmR��F�C2��HU*�T�j�YV�Zb��EU2��Q,K�!�	H�\�*X��TH��ͧ"�uKQQQ9�ȥ�id�Y��d�fj�dE�U"�IP�B'D��H���$��DRH��@���Rg�K�4 2�yu:�+�*Y"ԯ�Mځĕ�h.7��v�;]�ܺ]�+��0�2��� �m�͋{/��~����n�j�ln�do��2J�Ƣz�up�sW�ގߋ���_zm��B�co+)�U����]%�C�v�o*k�ko��;츴.2�x�ypjf>�T{m��q�9�a�Pb��V��������]�k��BȜ�;d��̒�%�<���\�Z��q���ʌ�R�������f;��ۡ�s�߻n^�����M��[gDb�U�����P�>��%���oa(���W���T�>���W�A6���_��h�N4�9�X/
ʏ$�8n!V�N.ڙ�q���O�֫��>�
muAO�|/�%��v#�v�fg��i��.HOPm��V��k��3�{�{�t�)�酴�:��*[�f��&��tM^��ҭ�4�G8}��v�R�q7СS��-�zs-`��>-Hc���)Ĝ���Z瘻��MB��q�r�q�^|M��zˬQ��9ZV��鷤f�vG�J��$��z)j�@�Y-/K�u����nɝ�l��KtcJ�S�y^pQ�uv.�ذ�}�-��]k�M����op��|
�1���@N����hu��X�H����wfw���G�}�}�gKu��6Þ5Q6��� �v`3���y;�އ���7z�k2
`Jy]8h�������!^}�V���.���(����[��vk��\l��n�E)f.������2�&�ݲziV�j�ZBs�:�V�e��	'3��7E<�P���*�������S������J[�d>K��鯵f􅨆�B�
f��X�]�\m&��ҩ���{��y�}����mk�q<��jze�Cl�|ԸN�5s�:��0�Fnd�+,w���M�>�bڥ�a�-���b��KYW�^(�6��ws�5s./pe|���`�Yx��)u/k�Y�Y������hl����F�F�m��7y��b.qX�j-p{7���O.�����*��Bӈ��+����ߛ����Ya.7cjS���ME�MJ|��D�7]�|�~�7ʀ^i٫P�L{�|pMmR��H^�PEw�cA�n�Ak���ae�*�j�A��$ԡw%v�Vf���=ݱ�.��Nn�:d��pqj��Uo�M��2�=T��TYvR�g+!z�s�ky��ojA�������}U_}�<�{�'�:㞳����]|�T<��!�ڈJ�kW����9F�.�K�w-��W5{�a�m�Y_>P5<{˵}��|���0v-��|�>{YK�c�O���p\fWҠ��|��J�ϝ�����Fi{����IXhhŋ�/"�Fg:�ޱ�I`�ڏ��{잛�l��w{���h��qW_�f�jnP�{���-�m�xa/�Y�������8Va������N3�@��N���ϯɤ��ȥ(��P�s��V�}��G�)��lNUӁ�1�;�=N�<C�!��n�R�b�=�B����Iu�_w\�v74h�}.3V�s�èo����}���X�܂��o�&��㠜��f�*/�Xg9��[Q�EW<����J��z^��Ǚ�g�3]0t���J,�'/��t7��K���ϗ+K��ƫ�@semI�A{�}9��]��ŪA�8�w\�ss@Sd�/e����z��d��Wǉ�U������yt1Gh˜�Ńt#��>u&�/��\��Y.´{NU��WL.K-���s[�8F-LN�
��o%�i��N�zL������p1����|>+͹۪���+�nʇ#��	`�����1�^+w߁U}J%��ɓ�է{3��=mj:��t�X�\ʆ�eD>r���8�ޮ��'#Y�NE��V�����I���N)�/K_{��ُ�5k~�+n�Zc�㈞�,nz�ײg329�9�����R���-)�pl�s�=�c�o����8��e=����U*=��?ey�q�)�鏝Y�V㖊��Zw�4ֺ�ߣ��.nt��SKq�l��-?��z��*.+Z�<��/��P5<�M6���ܱ�"�c"Î�<\4c��s��u<��*;*%A�蟩�W)�>|�52k/��:st&�����Қn��[q�Wã��K�)p�jÛ)�F�N�yy��=y��)�u_�4���8�S�����FB�&��2��kܽSwm���WM�J_u�{�\F8���#M�*��\Dl�A�,>����s�Ve;�d9�R���x s�_޿e���v��r1�9i�V P������W,���zP��CPE�m:��p�yKh)q�dV&u��*�(7T��N��v��bf=�S�cD[�V��4�*>�Z)^B]F�G�}��w�����_^�na��2Ի��W6�pI�R)؛�x���	�}�<9���&о+�w���;�u�}N���mF�ܼ�����53����o��Y�Ό������6!�K���8��vZ=�W ��N�>Oн����BYn
ظm��f�]Qy��ޜX�W��KO ���Yt��W�c]g#�(�L\n���w��.ӱ�LVy��y��4�^z�OoB�7�zr.3��n�����m�9���/�wqd��A����<��Eb��c_V��|��|1���j���n���荪���4�ۗ�ਭ��Ӌ��M�Խ�԰���^;��C5��˖�6Q�Ո�u� �z�V�y[do~��8�h���uN�<���댝0�����{T��[<����w�?v�7L���*-�XŲ�/N�t��WCF{�<�5�7{��*-+7��D�7H���ȶ`�=�a���^�`��̸�ĺ��4�B���{P[�rJ��F��bwr�L:\���\�B�M׷ /d��;��*��%�N�^%�PؖV]���z��������77;�:ǣ�>�+jV6�ծ�5�~��5��=׍�|�
�]ƥA�s���5�w^Y�q��7��^�y�Q^���q��S\�8�[7��kl����,6�^�
��ݭ���:Z����[�pJ���hm9n��J�1�j�Zv_^�T�t��*K��
�\��R��;I�T7�[�f�V�v�V��ɾ�et�Ƈ��}2Yj�a>�����NU�J:��O�����t^�b���7c:��b�F2���,�����}ۢX�wH�$�>w��*ѝzm�'Ҫ_&z���LR�b����-�T�mb�zM�3&O6|�Z��^wD���m�tBN����U�5L��lʽ)n���2�4J�望=J/RP.Nw^O��e\wN6��S��+�:��1��d�k��������c����8��W�65h8�%v���:��
���]�f���3��z*NL�xe���|C�F�V7�V�}׈(.�Du�L�.`ô���aS�SP�(<���*�֪K�����*�s��d�'���j#���2�9=��W�6�%��X�G{.VQ��tC��cǙwͻ���Ju�{����������N��i��Q�~��D�g��TE��F'�����c�o���B��Y�އ�|{g�6X�K9�v��W+]��(|
�Խ��P�\ؓy����`��b�w��C3|�m5�v�./8�ϮqX�8^Nis|�tЎ��ܫ�A���rw/b������sװ�o\f�P܉M���5���T�g<F�3)�[Qes�sasz�>����j#^�:�l��zt�#�y�/'_N�Qr��s��ξ���sW�Os�ɮ������nK��bG{�VWx?AO8+h��pbR�|�d��\��@��c��/:6�)["��p�|o�],3ɳa,�P��ۥ�I����:[�/W��ު���y�KuvT��ơ���b�P�oþ�*�wnLʹ�M��Ysi��X���gX��:_ո���}7�8��[�r��3����m����Uįͮ�>=�i^�Wo�ȳ�Y�zܤ��Jb��=<;z��Fɂ����J��G�'ww�Z��v�#C7c�����^�}��'n�{�݌���&���Υq�{z�|���B�#xs=p�T�Ā�.���[�XG����x�o.�7�Q�w��Ρw:�s��[���w�˺�Y�з��OL�ួ���侴�.��Wd�,̀�cy�M�;��>�����7�f�U]ڗ��@�X'm�x��1��jɍ���13�l�.�?Ob��oV���yES�JL��	{�y���ŀ�؜�]�B�m��S�7��q7�o�p[�Ofo��������I�+�.�`�5,1�x�l�Z�ML8��|�mG46a�T�Cx2��E�eWQoUc}u�Z�[KM�#�=�{Ժ�}Y3����ss��XzvǦ��xf�I�<�W��nL��tc�K���c#����^��!�&��T�zv�=���v���s�<���{ES�vDO+�Y��u㖊�֝�M5⛮~�w3݋�i�e�m��r����j�wP/��^.�1{��9R˞�괻+��0���}b�����#ki���Ԅ��inWb�
��gͷ���Ï��o���&0 ����]k��G*N�2M�78��08hu�_s��:� E֓����S�#쳒�]�Go=�-e���T&v�>�[Uru�1a'}�lOﾯ���W�{32O�ϝ��y�l��/�ö�@��t�6�� \������t���NW��Skx�|(,X�Ttu�Ia.����bg����f�*�6�\;{4�J��v���%�n�8�*�%P:)���t7sڱ.��ߪ�I��it��]=�j���
\��E��wyѵ�q5�`L�����b6X�򾞙�v���2�s	wMB�n������RMNmT뗭Ps�!q��'f�a��\ҷ2�y��s��dOvO��ͪ9J0�l��Ű��<	K4�ʶ�a�ŏl+Ц�z��BD�O��yʵ!�'�UDsP���8[G����G{�U�O�G��*ҫ2� ׎�4��wV��8�|�N���a�
�h+�o�^p��Aچ)��MJ���}���A����B�.)�;P�4��-�@ɶ�!姞~%���*8����,Kr<�ɑrG�f�z:N�>Yy:���*RK,��B����L�m�[�Ou�*���������9Y][�����Z��;9�t��&GX�J���y���Cr�
b���an�22�N��d�����}_|1���K��P����u���bzuF}Y֢��x���0�gKyS�A}G�ή��5(�_�I~��W�x��6������2���w�۫NrJp�+@�k���;���[߽��4	��d���/jꝿ1�Mޗ��,o��+��ӡ��nB}���s���2X]�ب�,[��ϝ�*��θݗ��&��v��S]�p�>���*���Q\z�Y7������=�;������*�V��[��[q���_�B�n0��Ț�Õ\is��e�c���k-����L��=&��g��YU�o�Y`B����A�T}��X�k�w�K�E�y��,J���߽�~�����|�.lp>�S�l�uNV@��G%S�!>���19W�=G%qv�x����˗z%9�Y��K���b��v&)J1MC]pad�p2��َ>��3����� ie?�OM�`�5�3-��r-���D�Z����Y��<���FKY;lU�����M���.m�h����h�W��~n��@㏌���dt=-s�L�5��?�.�&�X��6&���� ��j�ϴ��q��,Y�Տ�m63v�J����*��V�_�03�:���of��Ҝ̰H��2<强TH��Gn��Ǧ��*b�j�j@�SM�\ڀ\<S��W�t�bV1`���o�����R��r�*�8��s��l^��ea�и7&��V-ZqJQ:�t�oW,TH��I�m�v��^�? ��֒�ҁ�n��J�.�=KV�1�٣7�k��Y�[!���sj�KŊ�g�b}�~��x�ŋ������"�:<5���6K����}VZ�4*���w)*�v��)S�ʼ����m�n�*K�ob���S�eN��+\�j�q�;�wuT�N�����X��8Vd�YUz���R���kV��p�n�#6��}��hB,mn�z n��.�iv�μ��ٹ\�`d2]�'$�P��lFMj����b���A_�T+��Rv_vU�-��x���l����A��֡NmeM]�off�?�)ie�j8��痝u���������-OIx)<�Z6����Ӭ��͝Ž\�Ĵ������Xh[�@��.��Z5��rű���n��sa-b
��$@��s�^�b�W��hq�$�iw,�,4��������a��TѰ����Kl���&2��.�����D��e]��3^��(��^�4���&�QrV"R̲wT+ <���Do��nڢ���)���ս$�������cI�*��,���.��Og>����4&i]�\�\�V�ɵ!��"�ňb�.%1V˖�M]w�A��D�rT�j�Zc9,����[��׵��81� �3L:�2�B�Cq,���S;�4�Y!N�f�m*�VҲ�Lt���+�"#ug�]�,} Y׫9	��/�׷����n�E���EAέ�SSC�s�9��鏂���k)�2�Z�)��!A{ʛ'�eL³�h�w�u�`m���� ��r��n���)����v�9���s��I�(p�:�յ�J\$u���+�9�R�e���m>+�mKU�Е�`Ȳ:�!O����\�=w���c�v�]���n�r�YgD,Y\wiN����Q��c�ڰ�� ��d}���2WtV�T�1^-���l@j��;�rIO����(�dyT���"P�8�[�s�,&{���� P5&��8�nU�Nn��lm5�]�K�����A�PK�a����b�Borڲ/ǥ���T	�}Ł����Kl�Q���"E�^f0ft�O����|��j+�����!/�ڱ5vr��XTp���J{�8��rsc��39���"�I֧�W�\�OCo�����]�0�c��EL����%�v����]˛�n�%�P�&-^v�\DH�1jD�kg6dTa�	"U�@��QiYf���:�F����i��V��\�ʸY&jXeBD��"p�!]:E�Ue�(#9gH�&j*���L�A$�sMITN�f��R��Ј�*��ȩ-K�YЮ�gH�
3jad]3	��T�/<�ΚRA�#��;�,ȓ�X��M+H��.��U刅dJR�����A*��
#�C�XK���˚��ը��)�E9#��
���K��[��mML��	N��R�$�kʸ�z.[3e�L�DF�IHP��$)[D¬ª��9t*
��	��*i��Uʢ�2�������Q��)�)�]�ۗ�mE�S�1���%�,D��[�9�����j��K
��!\v����P��
�7���]��-�O���ﾠ�0�A�����W�+x13_��݈��a��f�W���w�)L���e��^L�}�a\�Pt��a�|C�1�5L��[�u!U7�'b�:���L�W�y��>c1㚍y1�AWڤ:��5�Ӡ��IHaXzS�Ӯ]�l��yiK����V�8���۵�\W�Qܰo�O u�r��{9�۸�����ʃ��ǝ�iw�}Kf��\��G��Ϥײ3���F��v��5�5�������v�1�b]G�˫�]S�6��ݮ5���N��k�_M|��cs~./8�ѕ��=L%���)Q���o�=��
X�n;ݦ����`J�ݍi�z��m7�?^ճHLߧ��{���kM�}I�:���+"j��0'�)�������xo�����D�!�h(�jw�y.ȇo�J�5t��U�iT��K�WE!��r.�����%���.���޿PQ*�����C������
�wҀ�Z��Y��`�8��ۇDw=�7��A{��\��˾�N�=�PZu�-�)���^�U��g�Ce��ެ�N���|��8� .�ot�I���u�M~���4+k�)p�����ڄ�U�¢�R��|�䮯�>`sJ��%��5ʱ�g6�����=�~v�K���B�o�*-��wKߏ{�]� lT�7V�C�)=�.������q��:JٶVK�G,���`s룝��:��y��b�[��78�-}_@o4,��:�u|8�!�k����VV�癣�w�p7�!�K��9�w����v&)K0�Ef�$��9I�>ݧ��l�n+��{rk�Ovf�0�U5�P�AO!`ꧻ�t��e-���pQk(����)��9�y�ATjb�����\�I��;��N[�1�ɮa�0�������)v��.V3�ޟ\ŋ�<;�Y��3Q�<��ڕpہ��.`%a�߯�\y���U�;�j� ���`���٬�A�`5p�n�N8|�w�r������7��8��Z���+�q�F��?&D�݇a��Q��#I�LPG������(�Q���J��u�'yѱl:X��:��0���>��V[u�Я�~{�E
&����6��Fn�����ꑮ��*	u.b��U�m[�)�N�s����	I�rm֭[��/+�b�F��PWR�i-�z��k:���}�R���ӳ�]?�,[Kc}�WR��珆C��qڜ�X�C�t^Bɠ<̿�\�yS��mK���ٴy�R�<����y6��I��[*lX4�-���Ep֨p��f�{f�mKs��+�"�r����Zu��oth�6�s��[�o�w�+����2�y>�N�`O��P+~�1t����T��+WU5*��q�et`-+�?x��f���9�Y�%E�ՎQ�N�r/`�d~����6���]z�ꓹ{�?{�vo���KqB����C�3g�S�k-�9{W݁���^>�V�i���k���L7M�q�U�a��юW����[�Q��uA�NI��Շ��r��J_u���nd�:J��_�=;���ʱ��bv+�hI`�j'�~]�]�a4��aN��:FH�S�7z���k�c�m��,�|�5��p2�2��]��"�蝂ƶn��:����Wz�C9և�	%B�Az�4����yG�us�9�< D.��o9�]L�F���#i������z�ZA�o-�'K�{C��Ħ7���E��͚9k��c|�s��n^eE��L�+u !�۟������}��O聘��Ŭ�n�Ĭg��2�n,�a�`<|�s.��A��y���\y*y�n��7�PӇ�
nq11�}�����rSޙ���޿uf9���z���%;�B�.��j!��aX���w]����)o ��ss׆z�^*f��f1A�:����!�+Z�T�X3�+��pm�ВO޵�9� {ڇ��믭k��'+���֨?WR���x�42U��jEeTl��|�殅��X�?`ݳ�ߨ.:qC�u/m?R�)�z�i���2��=�5K<�?���]�pm%�v��ܞË��^�]S�-�l�^��-�򴐤���>܈w�M��}���7e�@��H"���VMzG���s��8���5J��^&��c&�v�>������3�=���1���.���ϲy�Z�jx�-Άޣ<�����RR��^f��X���zZ��f�7d��XL}�*RFj�%�C�h����=����.z�b�Y�!tf}zHtF>����Oٛ�x�J���6{��:	�;��<[�NlՋ�fv��юR7�ݴpDnN�ŃuW*���QYLJ�H.����%�����G��Y������Ԗ�Y:���r�9c鿊i[��_B����{7YY�1܂=�}�a�w����I��������L��IP��������6/nP�*.�#_7,����]�e�bywA��` L���(n�dq�q�7��p����\x���HB���+]��ؗ N�e�@��F�m�g��x��.���Oԥ��˶�,����#9��85����N�q,�U�oPT���>P]�{�n��)B��c��J5�X��Z�Jx��Z�8��F����*�RCj"i�%�{{)���{�t9����O���<&��f�ی��X��ޘ=Wd]F��i�-���Ҽ��~��U��j��P���˷�+���m5�h�NU_f�k�K�%u�zyJq�8��pǔ�����eA�u9�͟��
u���� E��D��jh4�dUᮞ6�֕��a�_vV;g7�y�x�N�{����5�E�Z����;]���1AIz��T.���|������1�'�u��H�٨�!������ì̔��ք ���t�vr��7+��a&��yUv#/�N�舯Mު˦�����62l����oUC�駸6���E@�Vq�0��\��J���k���q�n(��^T^�*!b}��[����Ya)�Xױ�;7q���y<�i:�H�}[)Ŝu�Y|���;P�����܆�~S݄LU��f����|{�=_�5*'Z�ˢκ��5cS���%��N3�vJ�b���,�Xg
���ap�
�U���;�{��n)TP�&{KU�{��zʽ�X�{ �%�P�����G{Fw.��<�����gլF��ΒH~�wm/Sp���}[뒰W���	/�����꠳��4��X!�;w)���غU�M���
�_;v&)J=p�4��OkK:]mgn�bU�|� >̰���$�S=���:���t��WW$�+ޫ�+������ɤҷ&�=�
�y�M�8j�U�P��4<o/�i�KV>/���k��!Y:���h�w�s���j��T�s���u�-��y��,�E��Q�Z�dū��s�LG�;6���{�8R�#a���=õ#Ӣ�g*g��u';��$ş��K�P*��u��O2%2с��pg��yһ(+�:[ä�#��I��Ʌ���o`�n��K��K*/���~�X�U�m��ʍ>�R�d��}y���=`�4½���f�U�*��g���q3;��i�Wv�\��A��aP��Yy���eE�;
�k�k��]u�E�㯪����;��Jq<�o�O(���ʈ.J�L�2�[W{s��^��JM��K�|���7��;�{��C3k�Z���	u�p�2ϱ��@�l�9��t_E~s���_?�/\��B��M����̛u�ri�n�u�g�rp�W�j�6��x�����:0s���]���M^�w�W�ظ�d^e=����wZؔ'��ҠֵVyW�_0
ѯ��AF>�Z�]^�ɧ�z��Mk�M\֥Ak�:�쨉Pbw����ł2jf�ӧ�F�^%H����ި|���-��?��w��یP��tvFT���9l S�7>�('r��ˋ������ޓ��Zث]��ݫ�.ăF�1Þ�D�����x��}{hƑ��	}��Cu�A���:�^j߁��8�+��`�#��ss���,�Pj��=����.�dUܡ1�/H7����R?.G�+z��/d�4z�Wj�b�of�i�z�%��k�r�t���o=�=N!r�y�Ȍ/ȗ���us!�O]���1t¾�E�s{�^8��\c�ت��g���ݞKB���Fk��VLʾ~&��E������ZV>u4���΋�L������;Å{�Ӡ�������̰�6^ۺ9��p�v����i���:����T����f�U��lA&��Z1(��Mxy��3N������-t%ơ0�%�e��_]4�u8��쬌��fq�x�{ӽAR�-�5��aX��u� mv�B�]�kǥ�Z���Uyf�(��e.�:�+��|-���p媝�;������zL�G�V�,g���[�ژ/�
�y��La�����jYy����&�y���׹[f���]��)�M�Խ�ԍM�Lp�U�u�|���QU���u�E�yA��r����raxrC�VW,�qJ:2+�t;-��6�[5��T筨vٔ�+�2���v�\4��`gh�����j����_c��&L�D��B��!k�C�{�Ϟt��^kyr���?{`ϼ���m:�ʎ.6�3�B:�N�}�r�����h/�_4�x��|�u�Y��u|�B�nJ��ݸ H��"�*�6ك�t�VW;�*5���[�ޥ4�~w��>{�u86,��vt���\�\>.w����:a�>�>�����l��h�c�Q��Eq3��dM2u�rq�P�쨗%Ao�8l�<���I�o���W�����kUr�K��&s*9�Sv̈́�0�T::�#�����o�}}���ҡyD#ĩ���x����w�Z��e�4Ԣ��B����*���r����z�:�.�u��3���s����n-u�I�j�
炛���Ӈ��4�Ǩ�,��B˷�{�6�T��e�w
��?J�`rYݒvpK*�c|�҄�䣱]����_b{��zBP��C�*����t��es����Z�J9�Xxӗevs�SÄK�u�����/T��l���y�S+�&QX44!Oy+�����1��u�|j��Mܱ.���㵃NZ�԰o&�Q� +�fn.���^�r�ѻ��pbp����]cBu6�}cx����2�K�:�ow�S#j��΍�pJ����6G�Y+&�,�3v^y�7�x�ﺊ�M�pt��mȸ����zo���V��N°�f�m�孼{Z��Nb�v�>�����G��oѲ6�Ip{�)�V-�A�صJ�*��ʌOLd,G�Nb{,��L8����qq�����;0�#tR�����M8�żWY��c�'�7�����Q����������zi�����p\^q�(I�Ud��o 5�M���q��Kʋԅ%���'�MvT5�9\8כҷ��>�ġ	����U����N�B��ަ���w;{�eF9.��{9,��(վW��1:�Y�K�|����{���u�ިq��3$�3��gS�N�ެ�:�߲
�e����:�4��j��9�s�y�ylo%c��c[P書�a+�0���}�I���묾�����Itp�X̂u �EyќᎳj
 B��>(V�[�-D{]Ċ�6�qTu�@��8�e�Wf��Qc�i��&x����h�"�;�`3�rު�ہ����^��U�Bf��b�'d�s��M���L�������j��ҳGϷ��]��l����K��+(氳���]XM/�p��84vB̼��m0�*��N���8�y;�>�]1u����)�U�j2BT8j�+q��+q��j�b���'�a���e,��MG2� Y7�_C[է*d�/���CY
QVAW(q�y�ӥ6�asEFWdGG���>�ӉAmo7ՓX�`��b5�&c��3�����t�v,,��z�)4-=�I*g�����eL�S�F)�K�ޗg���b�	O��+p����b�|���Uu �����7�g}k�]�K!ͫؒ8���[����r������T�y�,�yY@b����v��L�|GTf%�mɯa���e�j�˭���IL׺��}�ƛ�w�Zژ m�[{�3e�/��ؑ��w:�����D�׹�Iξ��+��]X��k
	�ѡ��.��i�Vu����X����JV��l-3�Uz�9����x�<�7���{�;�t����;��%�c2:���z���F0�בF���X�W]v�U���xջ����g9ge��a�f.��*��|�ӹ�)��){���$ݼF���c�*�iU�!h��QOE�D��A�4�ܯd�`|���+:;�ԫ���$֓s_p�N�9��>7�>Ǹ����Om���aub�������H}�p\7����}U1{X�����Z	��Pef"�_4IG9ܶx���%I*2���Q��2���i開��5t�\r�V��N|\;pF�J�L�ZU�f�"zPF�5C)��}{U˕��eg58:��:�QI7�Z��d�P��B���a�7�'q1�f��٤i]`U�a�v�(n��&:��utx=)���NQ�����6�'C��[v>�v��x�th�Р�N��WR�zT�����\hk�N�w�<e\~�S˲���-X��)'�p�YhY��9vj���&F���Pu:���emu����]f ���Y������j]��r�kA�{i���ӱYzk�u���1�
�!,��^��Y��i�K��H�M�v��r��]�p\$u��K�N�]R�EfL��u2���se�����A[��H��VZ	�kmԎm���{�n��[���ö]�gG��S�`HC�(e���.U�4�6�Kb�3BU���K*�(�1����w���A�Bx//xe<�C����'p��W] �G�a�ҹ�>U���>jS���ί�rI��A|���Z*5�U�]����BoY*�m�$fbs�WIW��x���[ �\A|k%G'l74�w�ï�\�湲�&�5"��h�`�(�����4v��eJ,-�1S���;^w�6��� ����><��">�Ͳ$戬KS(�P��HKD�I�Zb2(�b!�rP.$%U����$aF�șZ$�f Uȋ3��iU�$D*DΊ6�H�!T��Dj��Y�\�	,�*T-6��v�V��Up�5,0�E
()5+Q#f�$��NEp���;.�i�+�\��,�t���Iq*T�0�dY�e��	DFq (4(�HE�.f,�p�)JH
�.�	R((��D�G*��IjQȡ�Q�Z�!�.��VJ�mT�S��9WNh��d�*��m$�YUI�2Ī*�
H**��*���ML@L�XUq �Ϯ�tL�t)�.��xL��ɧ,��E�j'��@�����ֺ�1�ou�Ц<�L��u؉˝�J-p��e��/�auC��R(�׹�pe]2n�r���Ż�õ���d��J�u������u_ɥQ�5���1N�d�+�BRI�G
�:Ѱ�;�j��#x�wf���>�W�4V�n�%�1[���"�TnS���Kv�;|���N����r�Oj��,'0�s�)[��bڄ*�]�����I���Y�ݸ���nMDb{�\����	�݊�۩Û�;�	y�Jz�#Sk����	f�=������ �r�m>Y�����	�����G=�*��jȂi�Z�L,���f�^Z�e�ggy���l�ozݬ�^w7T�IuT���
Gc�˃�=���]��D���^��$z������ݛ�������n>Gk�n��eC�7�q��W�[��NWW���ю1�Q7Ԣ���-���� ��}j�*�&��:��p=�"��w4qv���]K��-/��o�Z�-�64�B��t���;(6$��NX�`cb��/���v�;9`i	�G�u3� �)�D�l����)}�Q�W�m������p(�Gwm.�`vNq�Np{ \P�&�n����ov���!!��<m,��Z�Y�XTg���ڒ_Ql��[�rs�I��ZYS�|�l�W<��`�{Y=�oo�/mT�f�� �E�����'%�}X�;����Ͷ�Od�~�W!�u����:����DN��u�-U"���4�&q�˨�_��Ӵ{<�J�����-1�b����0�L�Y=���Ǎ�iOԳ���j	�#\.�ƶ�<�G	^(TNW��%��J��(�Ĕ3XȾk.1t�{54�5�v�����+�����kf���=��(Ƶ�����~s���*��	�Cw�k�}���,��4��N9#ev0��0��"zd-w
]��+�gqd�o(�G����b'��"݊Eơ��&+������1�
î��6�s�\�&-�ޗ�C�MT���|S�V��[�AK+�Kk�a��o>٬Bt<�.��������I1U�j#P�+�i��4�D�y{�����YemqJ|)��f�eYcӳ�7��؉����^���7���dc;��(#����Un��F>��y����;���y:��ʷ�3!��.�uu�<����m�}$��Ey�����8r���c�����4*��R�ps�E:���v�`��(f�N1SZ���X�o]]����k�g�����\S�u�b����0�ר��y�Q�&�w�޺�\[�\w���Eb��c~}B�f�5f�������)�����v���_>-�;�U�WQs�Q����KƑzp�P����Ց��ڥeW��x�sUӿC�Q	`ݳv6��s8��]N�%46x,�s�����>���V�sba�7��Yt���Y�*=cV��(vS�c���9�܎C�����o�^L�}�d8����י�\�K����,�o�h�����#dMN����tj�1��~;7\�Ox�_[���ڨ^��;��B���7�Z=��W�;���=�g����K�|�o�e:�Ts�T��-��p&)��ԯ[0�O=�����]^w�F]��y!��s1�E{���P�~�S�Yyd77�(�qFG�t�߲Z>ݘh�~�eqF�)������Ǭ�K@�WC���-�n`��Ȱ�,������Y%s�W��&	X�q�[�cWV��/6<�T�����+�K��$=���_#Sts�]д��2k3y��A���ĥM��T���(�6������3��y�	.;���;1BZ��q^�V��O�~;�:*/��E��^��I�
geL�.|�nnV�~��	�)��r�����>�bW��+���%���iw��"��9 \y����10�.��vL���Y�i>�N#� �^��|2�/ZȏU+��m?L�O�h=�lϤ�}8-1�	�.�o|�j�(�M�{n#)IVѸ�s�ݚi���UY,\C�׈~���T�r��?#�@�E�{�|-\ƈ�@'Ѽ�x3�sbr���n�w���Z^�U�xh�V)�s'�}��6b�I�}᥻����c�t�g>>�DTG���\��g�p{M����k�n8�&j6��Ӭ|�=�}�;ӗcw{h�C�UE��Ͻ�Q�(���}�i���2�=Z����1�񽥽wo���1���~�\{~Nk|@�'S��ݻq^�Qè���s�6���3�4cWY�Q�wԼ�VVǲ�{gEi�#==��f��.3���@��y��:�ݶx��碻�؟f�@b1�n�Y���Q�Q�]���t��3���@�}R=���"޺�=��]pڴ�w������*�*3����N�ݚ�&خ���>���9n*;d^�\zn�l����i)uL�{r��s({ڗT�2�� j�Y��"����!�ݾ��k�:ջ��X�qʈuS��sb6m�۳X�-D�L9�_u]ъd %/e��sy�D�j�;ѩP�1���rNa=3��WL\dγ��&���^ң����T<,����ξ�&�����3��{/�����b��6���`Wz��)�%���O<�~
�t:����3����.�^��F��ŭ�_��uj�F䳾�(�\Q`O�����'/`e`�;9�]�Ng��;��ͼ�+��q�<V�����z��B�ղ�3Pz@J�*�y��j_�ۼ�-{M��eG=���i��1ޅ:��H�W�w#�+�X϶b[*�L����%�>��}�1�*��|N�Xr��>	�(��A�}����˨�"�:.�8o`�^��j�ua�'��F{�b_��({n*�11O��s�Z;�X�Ct����*�>�`�+����\�U�[��+���ِE�Y���=�2�__���>��i~=�a���^I��O�^�˲�w�yHf~Hx>۴�}X w��1^��I>x͆:�h�Q~��_iz}G�A�����+aW{\��튅��4{�t��UX=��"��9�/hς��7>fֆ�X��>�;[Z�����Й32�jJ�sa�vL��{ٴ�O�	ۭ� 21�%�j]�gj�(��6�i+�d��˰{M�+0�*���׮��&i�'9ͻ��v�Vأ�n�[�!KN���7�JӔ����ԬKڡɤ��O9���պ�5�&C��F���{,;�Ww���L_��EOw��yen��xT���=_�J�s���;�Y�[�B}�{gt���:ρ��uz���V� dyS���mX��{l�>�u˗��ԭ�T�_9+bs:��>���مw/K
3f��k�7�����x��>�}ӡ)Q��碾y���k
|�C����H�I�:�*���ه�g��޹_I���<��r��ɏ1w���i�;s�J�M�!���RrK:M�;=EV+�w�L���&E[S�����g�V��:�Z��?o;������}Q�iy��Z)����������7޸u;�=�tr�D��d������,�F�������s�i��~-Y���\o<��(�P��J���Q�kѕ�Q:��l�[�wz��S�E}r�~9�,~��!���p{}��{�8ۿTz�G��+�UPW+k[�v�V}���T�S)�M�^/s��ø��Zd{Θ��D��Hih{$z&���%-�Vea�KB�Ge	���!��zۊ��V@h��mCT��4�R&>�����5ME��]ppfa�ù]%�D��<<���x��P�I�fy�P{�������z71>��Z��O�}8Ƴ0A��e9tl�	ur'*`�;�W3���â�p0u�qd�Ң�yǕn�.W.r�L����7'�v�+����/n��{���W�w"������sd��̣#���Z;�a���_
�09�U�&���Zl%���R�F��x�V F{,���T����Ϧ��E�"��9���ϴ�K������Ø}�5�xTz�U2�>��� ���*-�zJ95ț�6[�%�Ey�{g�Z������2+T�`,er�9������@���c��w@Ty�zK�7�>
&�i�ٞE��<����~��ekc��:N����1��VK�\\{΄������57a���C�)����7���釗9�����O5�� %^�M�ψ?DoM����܋�{�����M��_b����6�V�{B6]y#�pVؚ���X��0׋��_q'�˂עg�;=w���k�8:�xЃk�Pп{Eh����ȟP��vX��ۅy>W*�yV��o}P'r�.��_�������}~��u���3��\w�V����n8�=UHz=��>��탗A�{�<�\�{,ףf_L\k��7�G���x���\v=��}�u�ym�o糤�f�0��*=쭫��ޚ�/=��8��5��Y[�e�_L�x�/^�WF�b�����3��W��5�OSƬ���~ǩ�����3"Wr`�:����9�Ϭ��]5�yͻ��J����.�Y�@4��V�I�<��={Rl$&��ѫκ��Ar���L	�縱q�:��ϑ|�CP�x��9�;��P�x�=��Qi�xe��_��Z��?r��7o�M�U�(� W�e�ڨ^�=O���G��g�Q�l�)��̿E���e���U�s��w��(�ۚ�b��-��mCF�{�<�a�}B��b�O�����޷�k��g}�q^lw���z�-Ue�^����s �d�h�h�x{��_���_�'�f�~_���F>5�����sސ�g#}���n��ޯ�I�0y��U@h?w.�{���E߻��o�ԙ�J���_�r�x�r=�Q���u��̹ Ty����ݪ���YE��;[��.K�F�}���zS:0�Zw>�Kԇ�3��A����O� +�{.��Π[�1G�x�;_l�|��H�,�+�$D�K��S62�1?SU�o\�wd	c*;��,c�׍���Mj�~>�cø����=���g���	<&�93�z��_�[�竤֗��q�ᢹX�+׎w�kѾ�w���Y����ϷU �G��g�����Ĕr�������ݨw�^�|_/�`����{n�Vq���*�(z�_��E�X:"W݇��N3����3�M=,��}�f�S
�:��G�iN��d�X+�v��f*��D[՗���]\@働�l�PH9-)\���l��S]sB�����N)�qWN�er�Jآ����=��Y�[P_.�M^f_�+��22#���Q�;��@x+�%�� ��,^�z�;�<n�SmկU�k� 4��W���=�7��M��G���3�'S�ݙQ[���t��Ӄ�'�=n]K�i<����������dc�x�"1ϸ�6������c��H�TM{z�}�.���0cW�k�Wy������8E�~�C+&����}�@��G�b3��C�>㾹ѯ{rGP��UG��V+ᗭH�X[�G�y�l��s	�~;�+�/��n2g�<�tc��{M��Gݗ$T����j����O��vW�[w��^J�P�$PJv"j]�a���L��U�~W�k���T���Q�K�<S/�=��Uj��,�G�@S�(�tXM�<�u�%�p�$�^y�^�Ӿ١��yy\{�6s���|^��_�}
r�/4��*@Z�#f/D�=�W{&�!Z}�"�Nq6xw�{��V��o���=�|��0�z���r|(���Ս�yZ[w�X�e�����D⬆W����<V�\��=�\��6��Y�ʊ�|-[ކ_�ytV+F�7H;Z��=�g�
j�b�V���-+���#y}c��GhD��Y10���C\���l̅��i
x�7�Jݦ��;��]QQ�˱:̖$���8�8h���'s`�ӊk���GL���/����L�6�Fk�:���b�ޮ�J���L?}��nn��}��bǛ���~�yff��ܶq�Qޮ���gb�@�X�+�&+��p.z�s��� =7�c>�մt?��L</6u�ў�L�g�TU��6=�գ�΀��� ޺m߮Q33�e����O����B��6&U�ɼ�F]Y�>����~Vj�Vٿ'�QϚ����&��//���rn|7�omo	��:V	�.������<'ѳ�f���噐ڙ�L(�8��~�V�C�4v#�Ė^����m_�*�����t_�W��.xg�2wK��tV��\���µ�����}�3���ׂ�u'*��g�;���<yr����DW��gnv���{��Zu�3����Ul���^�f}38z�9f����m;�1��?|�Eh����M�h��J�[�^�W��3<��Jև��9��
�z�������'лվ)?R	�Hh���p�2#vK;s<0��=_b�����Gw���ۺ�=\��\�� N�Dd΍����N}����~�\o^�|��c�Ok�����_U�������׿�_Z,s#���d����ܲf� UY����Q�%�+QB�]�+��6��qvd*�aB	��Y�7�R��2����#/:�����\毈�]9����º���ӫw���r�\�oQl&&�_�i�on[�5��Ҙ>j	�m�i�c����q6��f�0�=�+Y�rˑ��j���gV�.-dh��;�f�	˗w8c�m[�2�g �3:��C#����jV��1� ���em�v,#ʄ�r�zR��m`���-��w�b�7�[��]aĸ��[�W��
�h\�ҡ1�F��XnM�q�!{��X�'sT�w��Į�-�wQ���iZ�]S������>���:��%�]{�wP�C��I+49��Tw�'q�ٺq�xtw˵�����v��ӧNEkU;3t��f�"v�+J��v�BF8��Ld�X��H�}C
��X3f�+��&1Rh�B���h�]Ϻ�g6[��7rwM���孮����R�t�����U����}��ˮQB�����\���h)!*�ŉ���8��Lnȥ�ݳ�:"s�q�a��#�y2%��n���R�5{g��7d�ǲ�}�xlŸ]uҧ���9���pצ(��.û�t��"�k���"�en�j����ġ�M�K��\�P��2�eu]��.�u����=G�t�=i�R����.�V��I`,�t��dYSIj�wY���*�s뗖��7}ڀ����!{m*�r�A�k���#t	��#����9�r<܍�������`8��/]��,���,#)rU�lc);d��Φ
n��D�����̤�\��x���8�0��KZl(H0���\a�U��n+6bm�-�Q��k.���Nc�eK
SF��*d�X�&�yB�5�.���q5���ߺp�#E�eJ�=�g7v�:Зx����Y�5���2Pֲ�kNw�7���\���;5��u��R������eeM�ϔ��S�Ƃ����Z�����eAPLI�8
ONu�B�8窺p��iC\U��}EV�s��43�7xǱ��$A��܃k�v@qvfT�/�V9�Wwv!���ρ:tB.�$Z�5[c�M+�o�T��"��T��p�z��i`"�����]\bb�/.�A�b�e��,�'���v�J�"��Q�[W0@�	��'q�aP��c;(^!=�W78X���;R�����Pʽw_I�Ukh��kX�tEY� �M�x�4��f!����T��=��r=�k�����8?�{oRu`ӄ!�K�x�uw���v_L�{3L�lr�.ܖEt��q'E�RW�4�M(�˾�]܉и��S�}n*���[3]+ǃW�L�Ŝ$�F�]	B3ndꏣ�B�
V6��t&n�l)�>5���k�yۊm�3!+.l�q�����D�C��Az��:d�D�qOW��z��㪀���$�
f����ڭ9W=�u�) ̹D�U�J�IQ%���[�K�y�AˤEd��)D�9�M:Q®�J$��Y�QeTe��(妅�N����E�t��$�q�%���M "���gH�MVU(�ҫ�BU�2 �#**�*��#��9IW(�i�r��$�7]��fg �8�F���Q:��֚��!�I���bIV�6��E&U�h��$0��*< ���*��T*#��ZJ�B�J��RB#LR"*�k*Ĥ��w�UW4�T
1*�V�$��P\L���Y,��pZ ���DŔdQBK�8XI	�S*��K����ue%�_t�z�e�Wўйi�/�)O�-�8v�y��t�gn$�����b�,e�\\����Y�0tJ.��:K�V����R��t�m��ϰ�?K�h��8��Q�Qe{d	E�b1]���WG=P	���1<���#�s�c�^�=�����.9�O��C��ǭP��MD��{ӛ|=��e~^�vo�*@[uR=_L�Q7W���aS{�B�?:b�}�=������6���Fm��2Vx�?�eD�7qU!
��Xp���fw]Ƈ�`�S��{��n�A�{��׹7>�>����y����~�R7ޯ��i��6H	��)�_A}^�G0dw�N����o�Wo�Ш�⨯G������\{���]7�t����"&��Z��_���F`G�Q���҅���{�|��ωxjb������s���}$���t��ץI��h���jaP�^(N=���S��/n��^���;>��B��u�s���;�����
��'r�L��;ګ�,D/t��蛞g�r�m��z�O�I��:��Ud�ԟTt{΄�G�5w\Vy���b���PY�vY? U������m�V�f׸�zx��`	J�~����1]Q���1�l�k"���*�/�:��s�V+�է�T��ЬI��j�CX�uHhÿ��~�Wg���Ѫ�j�K ޮ���j؃�����}e�c������Q�yѥ���4F���:���z��t�Pfv���;���xvt��=Ncg�ig`|�ɳ��z��BO��GL;=��y�Zt?����A���Wq������� {v��lߋ+�����A��߼��ȟP��e����^�FFxg\�y��W����<��k9���x�l{�	�<Wq��<[X w1b����ܿm�6[xK�t��:���FL꘸���2=�O���w���4-z��?��l����rϏ���s�`l�Dٰ_��`L\�����L��ꃸ�����μ�o��q����J��Mt_{ۗ�X��u�+��L�D��⩁?T� U�S/#j�z�S��L��h����U�Ǟ���
�w0��î%R#a�>��z��% ��j
n@ȵ+��mCE�6���=Z�yޕ��u_�=9Sg}õo��_��!NQe�͒�{7dz��@�����sӷ�US����g{�����Q�ґP}�y����e��d9�'�2Hh�-���̓<zέ���p�~�#��<�϶}�O��=^�GӼJ9��#K��Yn���q��잻83J�"�B������t�Y#x9�j�u消���:���|�Q-�U��h+����%6�vX�oEBmճ���������n���;M.l��7�̜�je��tI��u��8�]W7oO�AZ/q��جi���R9���%��;���j��/�ڋ�L�Jy�}+N�/}�z���]T��雉~��V13�}�ϞzY�J;�c���@�Al驇�^&&)��:φ�-Dr�%�o�~;�L���M���Ӊq���}���Ǯ�
�@�D�y70�r�L;��t�����:�4�ӲL�E�����kN!d{��}�g��@n�?`�5�p�|���9�0�3k�g&�+���c���$�wB��L��\j=����j�|E��'���m�{�8|�(�}>����2�=�e��2�ڲ��O��3�o�7j��i�}3||ū�G�9�� �iO۷q�GG��d���&�,�'�ia��W�?O��a�+�'´������ڌO R��zx��#yb���tP<�L��wU�W��h7C�pǣ;E{�D�uL�^�Mib�&w�����P��Sd��}㸸�M��w�3����������1��%�rV�0�w�3��FL�'��Ƽ�p��]�ގ=�7����*��WhhϽ��ȇ�)��&�Sq5	��ÿ��ZU"C�^g��ʳ6OoF�s�-�����Dѽ����
���V�:�߳��ߌ���`N�3t#5�v��#!���+=�z�n1���1��#�ԥ��堄��Ts�J��&=��u.|�ٜ�:7.�@���b�8�+>�6`��}tO?&����kg�v��P�'v��^�q���~�c��*b�Uz���
wg�[7E���q�U]�� �~��H�Ny��2z��R�8yV�#my\{ /Sg7�<W�}/����ᐧ(���2gg��c���_�I�Hp`7��v���Kgt�����m�Ȏ~�o�~�j/���ο���y�η܈O���)��l�A����A+�a�.W�i�N��QS�<���N{;�B���^O��{�p��/wfA�f�g�O���T���}^�Y9����#����Dg�r����|wi��!���{"7.0T}n�nĪOd�M��Ӕp?܎�Y>>�˘��9�O��W�t�_�#��)�q�/�� ������5��YD�EUx-ό�csd���ՙ9q�r�!�5̟a\U�Q���6n=�@y36=��&��;�]W��+��Ǯn��{�u����^�ٓ���g�>�d�F�=Q�wvs'����Uh�@yF��l�d�|b��fcx����d׉G�t졟�6�~��tV��?���`OЕ�#�"��@ȏ*s�^��}WF�lI�1!��1��cDY��k�c
��%���F������/�>۝y�kA)o�˖��l�ޔr�G|��޴[�jgbŵ���'.�F��M�o_:�p�:��i�=f��(��h+���nr����M e�屃���aWѪj&������`�om�0��=��G�Kz�[���U^'�}Y�~�����0�]�_��X�m����d���8_�����Ew�Iêf���}��7�@�'4O�P�o��S۩�����7��sǻ_�qyhp�-���g�I�YL��勞�?g?,�D�Co�����Nϰ�#q�,k^�aQާ���ˍ�p���9�(��+3a�ޣ��G��ʯG�]Ȼ��;�FL�1���_s��:����W���V�79�SJG��S!��ZWj��.
G�O����?T����"�ͩc�o��dJ�3�>�9Zo�o��削u�ӗ�����Y�������0��F���H�D�exW���i���y���B~/�˚�î{��1�En��;�8�5ѦCs�=����}+԰���l�I���us~�̈́�,��񡎕4|}ԁy�<'�~�d���5����@of��4+����GN���}�ۜsۇw��m��0��=�*�u��{'�J=�����Yn���Cţ��z.�̽��@��ə�hS��7���j���y�Gf�QA�������ˉU��ˡ�����H-��Uى�����CHOt0���9��ܻ��em����s�����|����s�Eϱ�ױ��r�+r�Jt�m�5r�T�:��\�{R�g1�r3�z/ӈ���9�>�P��G��W~:}:Ϥ��P��+޺�(�
�}PZy+��R�G�d�D�pW���}r����ހ^�V*�^71~��9��#^�T��ۙ^�\�������9s�{"r��N�v|6J�:���SD�Q·�W�Fo����h}�E�s���X�+
��+���=1����0�g�{�<�F� RO�����lIv}�f޶sx�!��d\>�'��{n���Eh��e~�ǵ�R�6�~Ou���}�xV����eϒ��\�k�z���+���	��=�ǽ3�4�,^Y�r�B��1>7�~���Q�n7�oS�zX���Y�����ǫ~��7��+��e=�7�GqSf�u;�_��Ū�Хb��A�U`U5��:�;}!9��>;pׯ��{]���t�{��tt��z��ý��fϷ�I�9�NN�L	��X��gY�ɟ"�Pw��:2!�י��g�Ox��X��gvzAF�k��������,�ES$R*v*�<��M�mL/�A�y5?E��O��M�1V~�V��s8>`�2��7���SRi�A
�Z��� �Q\76u3eK�-1�X{�/���&�)&r��E���� �8����]Rn�V����rg}�!���D��SݤGlO\5�,	}|8jQm�5�Q�!W��6Pӳ�;|c�`�ǻ��{�`s�A�S��v{�=rf�57 e�^.��o������.;��+�Ѯ1D$�ǲ zR7�8��v�~�_�gЪ�.��no�x�Q��5~�^��yE�>ђ��ُ"�%qW�ZG>�zB)��~�r.=�Ix6Hl�GWB�ˉN�}Ԟ���}�������Xml������t��o�ģq�H��3�dߪ�Q��0�wK��y ��@���鉏mZ�&)�x�+w���z���R�Lg��O�;�M��y�ź�:^g�:���^�Ĩ���y���b������{c+�^�m�#A*qN]�w�=�~�}V}�l�	��@8�T ����&g�鹇�9���t��/O�,� $Е�5�����E}yb��*��q�:�!�P���EG���\O��vA��y�P�V�p��&�B䏜����}S&kj=�_Cy�������L$_��+��8|�(�􀰤���L������H��^�wߛ�p�����1��`5Px	�W�d'5� dr�q��۷~��ң��/q��RN�#;ȚU�l�YQGh��M
�J���#�i����o=i��b�
���}�G9�+ƹ���n��nz�v��El	ɽZ`wI�5�	��hoc
������{Ϭ���C����|3�b,(��\�t��u��*K%%�
��Ň"kE1\�Zxc߬s���=r]�&��r%�;(]���%��q�F�nzXjy�}~�
����S�s[)�W����}������38R���0s�Z�X�ɭ,^L>��ی�l���-����T_ejӅ�;��/e��YEOtSd��j�F+�/��p�ۅ�J�n�2���oz����L?G�y߸���^����S��!��P��)��a�����Wz᝿Nח��b��oY�V7a�yq����9�ˇ�u�;�\�����*c�NQg�ޠ)��Pfz;\aj���>�0�]��U�
<�^��k�������/���>�^��U�Ywy�=�*+��"�t��W5��x��>�1L��%SD�d��w6XU���[f3�
�9�c��簦��8���3��.�nz�����	��F��޲��w�	EO3q�¾�R�Y�݉�z�H��_�;�����{�F��n��f�\x������R&'�}^ӐKGw K*��u\�IT4L�?$%u��t�Ҧ��A��d{נ;�fA�����Og� =5~�>����~c�,�R�V݄$f�I��OKw������/�B�3]�wi� �qJC�I�f��ݝ�O�D"�˽�����w���*�z�/5/[�
�ɛ�z\�����Z;7��`R��2-�e�X2�H[Y�m��h훛���×���^�x_�����=�.� �=�*/��r�ɟ�l1�~z�f|�S�b��7��7�o�ݥ&�Oi����+㟬�����*U`��I����6N�VGD�g���Y�����=���u����_�Dr̸x�]צ2<�N��ުc��R�n��}�jF���o�(��|x���7��FN�Ӭ�rX��ӎ�_��~�Loe9jћ�{�3Jn���ϻ��U����@��D�B:va��W��q�5�����yщ�(�.>f�\v���V����|O���Az�	��Z.#�Ew�Ië*��o�^׊���/q����{����7�6��Ľ7��?Z
���C�G��A�Igzg�{�}��wc���5�>��j3=��>�.�cm�_��o�����\o��ǜ7�l�+>}@S�X�2,E,�{-�ڽ�Ar�1 ע��7�p�&S���g�ғ��y߸�?��%�Uj�W���3��+��g�jX�/��<}��>"��>E���,z��hz�83Ч�����rt�n�2��_-��9�҂ы�*{��0'�j�柄ѵ��2�o,�OQ�R�l��Ջx�#�*�-�#m�D���v
�SQ�����t��:ZS�+��u��w��O4���{�t�hc�R�̢e�d����*�c��n��'Z}|Uʷ�CzGE���O�~_~G�D�S� -����l�o
�϶XO;օ���}����{�:��z�>=��2}��Cm��-2��U!
�^�� ���˩�������=kslWj�Fׯ��~�RG#��@������N�{¡=2<��${7�)��Lk�0z���_�Ұ]�>�W�0��J�;Y�9��R�M�G�1N��t<|���>�yTy��y^��p\�����g����Ȃ^K£��+�>�g�K�w��XC=����z�q泥ح �M�DT�?ț�6����ZdW��|{>�2�ޫ��nb���ĩ��:��*%(�^�w�O_t��(�g(
�l�O��D����ʇ���]�O�I�tݦ=\��`����c�����w{��y��hW�ۮ����,�+�	Xo���=1�茭��ͯq��O*����N`�x�WD��@V<����O�{/J��v`��<��=�h�ܙ�v��ڇ��3�P����Ӿ�w��9�{]ۭ���Q��u0�Z�X�[⏝Aңݝt/��Z/�h���xW���곇�Ӡ��CnÖ�g��V���WL���=u�yӳ�B�Q� ��O�s��Hy ��a��i�\B�Μ��Υ��&���N{5����6����n7D:W������W��
j�٥�q����9�v��V>���9ʞ┺E�~�ϲ��-����E-{4���~yp��H�Bɸ{����uI1�鎯F6B����ud��!�m��5f����H9k6_VP���@Ġ�9AKjF�<��]ؙ���x72@�+ZO�n�gV�b��ZK�bz�8cP�~ǛG����ɨ�O�ğ
�bJ�:rn&:`�qjCS:ed}�r�S��@��)�>�qA���=��K�B�`���E���tl���꽜�+"���� /���H.��L���k�.7�j��GX��Ϡ����nԔ�6+�%�a&��f$e����f��7�ksW#}���j�I�y6��U�ջ�	c+��LΗs����V%��t)�X���,%�2s���%(.��8��tE��_2i���W���.v��&�)��;��ZZv�9	j����r��5ǽ�r���o,��@S}���z�Һ�μ!Tꦵ��̢��6gS������ɱ*��lJ�N�W6�9���V��
�n�R���>�i��z����G��6��s�w`PNY��*A��.�$Nb��Rv��v����,�Ә��V��{�Ѡ�-��ޫh��c�]$7��u���8v�9ad;�Xƻ5���,&���7��S��������e,@U�.讽/���Z��=jM�w>ǃc�g]K�QD�3e��G[�q`k �)I��9�;1�$M�Λ���|k~T��q�b�e�S.�ܙǵ��A���
n��XqR�ۑ`F�xv�ࢬ���#\�ێ��aR��񕃻��Wr��C0��ڳ��o����k�8�4���ڕ'OQػ\׆��R�8��7P0Ƀ�	0�ų��x�'����[�>�rbq�����ti2��%y:v��A:�Rv!Y\���b��4�0��]�q^3�:�vm��mIh>�m���"��C33��aL��5M'R���ܔ4��ժ£�v*&��_
E�&V[$�N���+��ǖAN{�ñ�{�)�U&mC����oZ��%+��B(�m
�v�+Y]���S��Ӭ�sod�Nc��X����l'K�n��b(���=P���*�'���ac������P�Sӛ�� &1��R�������r�܌wM[�?���>�.�wn	$���C���\0)�H���mv�i�we3���E����qT�;�Xx���&WM��������Y�y��U�9�^�d ����<�e�7�>�b4�_Ui/� ��;)"�J�:J�����6��Ub�L��T=n�D\��AsM(]'P�UaW(BY����7:y�JX&uX�H�*&UH�*$�(��u�0�� ����(��
�]��E*��ET�&��TYDD�0�9S�W=nN\�2*ndr�

��*�h�y\�r*��9��
��#�m]�� �:J�i��*#�A�e�!9Ud!�E�Qt��(��s��2r�9AAr�\�Q�B"�ML
��rnI��8r
3M�'Be��ES�g+ZUr�]]w�.kr�c��G,Ȉ����ċ�L�Hr6AU�Y$P�U��.D.;�t�'VTG.�N9%��"tB�]ܪtBrDT��vQp�ԣ�;PJ���Q��D�I#RΌH��;�e���mCX.5�V�s(Y�}O�����7�u��c�Ĝ��De�iU��Ї��@�1	:N����ꥬ�?,>��7�@��@j�w�*��~�l�j����F�]���7!��޾}S|�x�����}qTì�����k���}�G��g��m?�}��Mm���qY7�N=EުR�F/C�'�Q��l�-�f��`M�x�y3��L��ꃿ�O�tJ̻�(/`�U�����q^��m�/��7�ʏ�/lL�E3Ҫ�Sȁ~)��1�안�A���Uʲ�֖w;���ӀjU���-�z���] �|����ޡ뛂PLÁ�� �x8P��Wk���_�k�s�^yq�ɍ��=�Ȭ���7���]��E}�_��!Ue�^��% ��z;ڭ/f��3U��q#����M�@�H��4j%qW�ZG>��"���D訿[��Ϥ�[(�\�k4�>�>U�.Ϡ�~;u��7����l��TWs����'8�}�<^ړ�xֹ�}��oS$�>gz&&��&i�x��>��p2�Kև�2��ʤl��љ[�����,���y�L�����fA�s^��*%��7P�'�����m�\�wAb�u#�-��.WMK+o��n���h�p�F+YC*�=����*
v*i3js�ԬY��� X��������;ֲ��5�{/eXF\����1���q�jr67&�wd{P��z�rU�%��>�r�v�����.���Yƫ�>y�����e��qmJ��!vw1�dr��%�}�'V�A�;s�&��@�\_yߍ�Lϑ��'*�V釞��{��2a�ўɿU�m�S�U�Y:07BX�:��~�<����^�"�Ĕr�}^�W��N��w�y��w0jI=�Jz���>�>�f����y�������'�ǻݙ؁s�|�(�vb�c���\��^�j+�S>�}(e���<;98�̩.���ǘ7�G��<}ٕw|inv��}���<�H�l�T�}��(a���&����7�F�o�,��O R��zxu���|���{{�Ϣ�qW���=�s��:��c+���������w�#�p��+^�{:}�����G�����޺П��F.!�l�vOlUC��R���:��4W{��9P.}��vp���W{��Gyz��{�y��φ�uv�����P��a�JF�>���V-��Ι�?.λ_����_�L�%�����\<����i��u�����J�.!NQe�G�@S\�O��6w�.��%�9���j�s��zd4_{���6s}#�q��K�q�_��S��Q���;��h�l-P[t_f�*	,fGں�R���a��9%�W��u���E�)9��*�j����L��ץ��ᾭI^���o�ZfwX��tY2��R8�2(���ǜ�wm�k�X��5�S��wN��4�ֺӄ.�}��~�v�n
��T�T�h��c��B�a��C�?Sf.�:�x�?^��o��}�n����r|0�h�A��ْ.	�d2�ml�*x�
چ�<')b�ɞ�����u�����s� c_g� ��t����3f
n*�1O��t���]Ԯ}���ח΍{^�
��l1�S��qR�Q�V ��p@��x�_t��n&@|k��W>�y0'*眢�^:��>G�>�0��rb�.=�W�<�ps`~�X��(�����f9<���c�+��ArP������s�p<>�����r�P�#��N{�����P��K���绹��5�=���\֏qϢn|6�kG����,i��,{���֪���<o܌�1�A���[ѹ}ڪ�P윟!��l�C�'�zrO�=?�vN���u��f�i�)_�<H���^z������r�@�W_���&����G{̉�=q����y��,,٭:��50��ϩ�u"`��O<Z�@z�����D� ��-
����WqȏT�:����ja�.�0ߤ9��}�{�]]���a�	Һ�.��}*M��5���*o�o���G�Mlv죋y_����������\��E�h�S����`M洱Ƴ�{�i���Gm��mܼ(-/�C��N���v��{7�~�?R�v���PCs�t¹��~�ǩ�!��6�q�X�xY���g��6����W��a��.�HW�P��Lꛌ>����cn��N����q�m{��-����i=�I"=9�'iy[�u���͏��7޸���)�a>^�fBq'~���_Y~3����a�D���{kyX��u��2�����ۊ��SȊ��-�ږ=~^�=�O�ё��F��o�����R�ꪽ�d$}�>�q�\{!��v��E -������g�S�aM���}{=]}�n����P��v�C^�l���5�_�<����nn	P̐�}+԰��s�2}��������~Vuz6��G��Hиu�H�{�H��E��H������i��6H	�
�m���-��n[��	�wpL{Ŵ�+�u��>��V{�� {#r�U��$Gx���{�i��d�឵DLR�ӹ��9�L�+�f=���s�>��+(�x�G��zY��#���ԉ�ٺco��ꋕ�E}�wǰ2�������������Zvw��<�J~|�X�����t{����\.�}���Ez;\��颳�Y9��]�2b��p��v gZ���$a�'&A�U�ڜ�5�6&4}�0�a��ی�;\�(c1\:��}�Λ�q����[�H�y���(00�x,Ws�ʆD�u�����y]q�W�j�,�I�h[������o�@W�w^���>Gzr���n�q���u�rX�֬�׫wվCu~�xn�U�9�צ�� =��� %a��O���m�n�w�^��V��O��RN�)�����{A�� z=���dCUS�/�u9=~�݊碴_����#��w���?TD,;���g,t�Ԓ�C�1����J`	�X��^���P8�gz�?`�y'N���϶2�=�e *Vm��j/�S>�����|�tx���Y�����ǫb=넏����'$����;�'ǸjT8zǣ{h�qϧ'�nMiw�;��!9�����C^�q��~-��d�ꫯu��X7M�4�>����J%������"�X�u�ɟ"�9���Ӵ:qH��A�����u��O���wz��l{+�n!ի����ό,�tU3rm7�Sb����)��.��;�W����'�|�!@��X��v��z�^��*�/_�=��Ꚃx�Á룣�⸌���7-�q�]�x}};�VF�y�� �M��D��H;޿_�)�,�7%]�v�Aׁ7�W��6��3�����c*腋��A'ye^��>��N��n~�]c�]ݩ�[Ο��s��M��%�S�Vub\�C���.���|���u�c��K:�����^+[٦��=��Z�0S��)f�+WZ&�Ə)�҈�����]��}�r�1Ϣ�����`�h�mCF�x��5^����uϠX�߳�#���w��x�{S����/t��$j>0S;t��D>G0�϶_�<J��{�|};ģ�}��z�۾w}�]������z#�,��Ϥ��q>f�����3�t�82����율��~���������wi��z� w�pf+ޫ� _���7P��LO��mg�w���aHp���J�Mz:����
��Y(_���p���s�z���My�R���}9P��L?G!�Ԫ% �f��5>=l�O�
EVu1��	b���?PY�Uv7�}=�E���\��W>��ofd�z�qW71_��y��p��k�O@~���ڇ�M�_�S3����7�TzIG.����׽�.e���J�h��*�zo��C.1֏a����Ǻf� �g/l{Y�����YPn�|���W9�]�9��Ez3�Η�L�ZW�9(m���^MiW�O�i�Fzz8�6��w�ɑ����U����kǒ���RF�k�_�l�<�z}#��c*2kK3�7�{^�>��pd��
Ȭ.��B%n�:��B�VWh�����{��b�UD����},�:Ю�?���4�V�>!l}�L<��X����7��鸹bմӝ��J\��;����׎��庌�δd��5Ջ�4����[����&�/ �7�noň��K]"N��זۃj�mpJ�J^"ߣ�H���+�����y���Q�{��9���z���c7��*Mz꟎e�������c�#�DmD.���s�3����uv�����H,}Lܛ	Ly�`���q��ը��=}�
��G	�^*'�\<�ν�>�Je������Tũ�,�_��z)UVnߪ�i�\�g�n̆E/\
�.|��]V8����=)�#Ǹ�o��w`E���ɥx�{+s�B�p�uPG�d͞�̑��]4M��w>�a<Uº��a�ﳊ��U�s6�\�b������4������Ic>ىl�<ت�0Ox�!��k���X�'je��otr��'���Pl�S��HҮ#\Q~�n}��n�R&)��/�0���QY~���ۼĽ���(*�z�>��U����L�V �g� ���^7�%E4{"d�����^���T�l�pKw#��~�ToKg�ǰ�v��ϣ����z}@O\*@_?e�n�R��GA����O{V�Z�;�lpی�#��d��Q��V*?Q���<�:����;js��MTwl��g#����_ �/ub��Z��m�u�c�'9����w��ؒ]b��Eܡ�Gm����-PӁ�@�B�����AOt5+U�Q�Rp8��R��S1&s��cb<*������ksE,�]�;R���҉�џ����o������c��Ǫ9fd4�T�`�X�>��5������G{��UZ+�M��,�9?�����;�����Zn5��f���yUw�1vU,[Q��ټ�<���>�7g��T���V*�=�/�	�7����C��+�X��f��^р�>�.�������_F:�-{+̜~w�ʪCG}�o_z'��z��K"��rR;W����]�M�ع�fd�>� o�H���@(Y7�k� ��-X%�h��\)T�b2Ƕ��*۔�r�1&��p*λ�y3�n0�f�e��j}~ӿw�����1��O��Ï����e�^�l�5�A�y���`��So�p�&S��|�+��w�{N|�/Ţ���q��_�p3������U�Ưey{�
f�Hn*�SȊ��"�ͩc�^�=�ݗ5W
..����c�Hz�>G�\�Tz�T�alC�tB rت��l�V{�=1�}��н���c�z3��|(\y���z%#�����������*���=��HC~��w�^�.�;�qт#�A����A$���-cc��·k)� =.ϵa�h.�B�s����^X�t}{JP��P%�ڈ��ߋ]���^e�Ք�N������b��Y�^�t3hG
f��))��{��k�w܏KZqvH{.�U�1
=�`�2�7J�.w�E�~�?����.�󼤏�^��{�H������~���x�3%�ki�/=�<��[4+�;���>�a��ި�u��>��VG�z w��!�؛�vƝ������\�H�gQE��0|6ԑ,��_���^\�.=��U�����k��5W���g�ܳ;�/F��*߲�H��L4z��c�=Dz��ZdTk���^�pȷ�,�ˏC~�[�}�Y�71��=��T�\�G�פ�*�~�ض���[4���O��g؁�*wu9�ފ�{��ڲX�s��2<���!��� �� %a���m����q��a߻�)^����H�a_Wt�[�gѪX3[L)_��!����rz��/�Eh�!'�\��;�V��M]�fv��ZB����U
�j�ޗ��q��j݁�Ӟ!z��鿽~����hG��zJ
�}>Zo���ٷ3��rxU�T++�j0����f�>��X��7Q�|��#�8����^�R.����<n���&̓�T��2kK�ɝ�Ʋ�{z�.����Gw`�o��AAݤ{t��*mrH������P�ʴTг{��V�v4N�S�����Q���*L�ٯ���E�V�M�	�\�k;m�.�.�\��3��
��NC�#%[���Qe֔Ô���wx�����x���VNS�n<��+�D����4V�ݓ�mW��w�qgIl�6L�(�2gY�ɟ"���cVϱ�ʫ\{=B�ԙ�s�w=��ګW��g�{����6�����5<��#���^�{���=w��u�\}�1�gk�,a��ў�-���Ü� �)��;#ފ���Ptj�g֍��;-l#��E@�S��h���Pѧ���=>�����ߝ���LoNQG��^ת�^e^Z��ְ1�>�|�d�_����[P�x�EtC�ZG=��w�pt��"{���sk�{�B�H��L�\@�!�p`�;*das�s>��3e��J��;Y�=ެ��_k��u�R���TO'0��]?S�r@�8�x��""f����>��`1t�)G�l�~˪������ʩۘ�>�~�ȟN@W�e��s^�ʉh�M�=��MV�q�c���i]z�u���x�{�X����Q~�[=�/N���{����Vlyt�7Ɩ�������ݥ&�����|0lG+�9����<����/E_G���o�������{t���L��gU�=�lӔU��2�,�g�[�U����$Gz��.����y�v�❱��VR�ޡZ%�d��E�ؽ�,Q"�,Z��Y�
��:�ҍ�3(��n*36
�b9�ֳR:ʔ�gC��c��t�\˗��x�[�G+t���J����C�S"�L��N�S�����L��NW�N�z�IN� �`K���ುr�׵7h��'��e��֚��N�{J	X��ޗ����\��Q��Z�O(���P	�3�\w4�ڝyc�<-�71pܽ��7nvI��b��i�uN����;���F�f�5T]2q��~���TD���8��<�+P�]��u+x� ���ȱ�t5mHR��)Gׂ�r����ӜB3�Z�p͐=:��v�6�U�U�q���mH>��OKFE���zv�K�ҕugc:0]L��;o=��aq�e*�UЇLg��S#�j��� ��wՎS�A֩q�r-���m
ޥK��s#�^�&��z����TQ�O5��[�| �w��V���5�a�u�.�u��v��:��їJ��C��f�[���c3;+�b샙�.�������u���&�yDݞ��OFeW`J�ٖx%@m0F�"�͗@��.���\dn~췲r��d��!�Q89e�gqA,��Nݘ�8������g=dF�&�&�V�çh��@jdS��ĩA������(\���"�1����nm��"%5���n�Gme':!c��c��R�p�9Zn���+�����7I����'j��v�!��c��\��9�L[KP�3B�(���	>�u�o�J�f�zY�P�'Nή"6�i�����PgNI�5�����wj�2�J�#�q���M��ö�.yԢV:Q��J^�l�nb�C�F)�6�e吸6�����Z�Ҳθ�ź�����z�l�2���%tBNxh-��3r�Uq鹊�	rt�dk��g*��1+�4k��Oo�=��;����aՈ8X2c[̋�o�:�Ku3����ɼ.�n��Y�z_)*��@�4�T��(_e�i�d�J���N�9}�#���rX�ۺ�(�h�:\6GM�\���3 ��{e���+�F(Yf��BT��*�;�mZs��s�C۷�b�j8J���X���I.s4A�Vҋ(,��D��zr�J\!ZH�'
��"�s���cCi���l�34��̢�N�&�wv]e�Y�aU���j�e�1v����*J�v=_^��-�)<����h�ҼvC꬙�>���3
�܍��;Ir�����.�u�˥�a���˽��%0��\j�Dk/���s�i�N.3�J������{P��q��J:�J�<H��J���a����UԦ���R��mvq(j�Օ�w6½��z�B�ሪv/�u��Y�9�<L�K����a�[.���39w�����u	҄�iΦ�EzJ��#�_q�e�"�[{��ع�9^b|�\�����$�A�	D�M!T
K�J.k=p��"�J��$�$\"��z��'
����*'2(�W�9�.%r�z!$$)�����۪*rtn�.�k��]R*�A���"��dȝrvUy�#��2�a�jӞTbT;�N�*L!������z;�sJ9Q���P�Z�#��[����	S՜��zb��w:I'�NN̉i��۳�L.{�;�Na�R�'	%$�TAk�O$�G<�p�+����=u���ș�Q�]\��*���*����wsn�O7StU��HI�����*'UOVh.{���ĕ*��Q����*s��AUNN�.�:�B���Е!Gt9S�30�J�\��AJȰȮ�tu��`\�Y�Á��TBlKbT̐�D�]��3dNiP�2+�v�thW3s-��3�-ì绸{�Nh�ä��Q�,��Eɚr��=���~���||��p*r�n��-�ft��\Z��Тm�/�X���uLvv���ҔTxb�wV���ä:uY:�fX��Ƿ+�Q�7����Mez|����f���P��熧T|F�1��UEWX�}��j3�C��4z���F��rg�t�{�zp:����Ǻf��&��#ə�6��g9W� #��}�糃f�},�{v������N���\2R��r�<=*����#==Ł��G�>s0�vZ���K;�j�@�g���)�G_�ݒ�d=�O���U1�gKNx�Y�'��!2�e�6g�}����$\=u�{c�\:��;�(�	�l�vOL��(���B��[k��.���3��fz��"6�]�~>�>G\G��G_��lp�!(+{B���e�q��U��z{ø�Q�*��D�x	��\z���&X^'��8�>����Z߽����Z��r���k���z�K
����*�(��X����孚���Y�ٽ��=�������{�7��gнy�鹦\ .
�9L���W�,y���O�n�U�_"C>��D���9�pW������F������9^��F�Kd@A��H��{Ǚ��x��9;1^��G7���;%*�Y<ܒ�:�;�ܖ;E�5�8�j�n�ޚ�lk����j��i�1��@U�P��돛��u*�n�5rn[i�ЗI�s��Ff��`�~��Vsv������R`냭v�}�%�J[�Ӟ/!^��*�|�x��(�y���=�E�*ǌO�8<ڤLL���d�o����V9�*��gĤwr�����z�_�A��g�z�]�n�nR����yTc�x�8�ϣ0LMyVѸҙ�����yU��l��{l �#�v�]�9���[U����vz�o���Uh�g�l!��m�/ղkK��7���b��s��7�<��� �x&���;t��K�>b�;h
~��"������6�;����cL�ic��2�}:��O�^&ۥ�n���M�{��<W�V�E���ߤ�����x�D�~y;�ד���}�-I��
9��q>p�@{��#�#ӎ�_��=7�p��t��=���HGn'j^W���<��/ձu����վ�}��U�S�׈�/m���H+��-
��Z/�=�r=Rp�kb�V������Nn7�����ʎ��U�w��uH�ی<���7����hu��_2<�R�nT	�{Bޟy�u��6Վ�~��}7Xu���L���f�X�k��9�o�����f�U=ѾoM"������""�v�Q35�tS�Uο�KW�`u��WD�������c,���͝~t���8?�9ܵ�;��w�j'<$:�nO��Z���])Vs�K�gm|gQY�^H�95(�`@z(�pb�k����;��A��Z�5WQ}���*�ǡ=���uN�̈́]Sb���&S��|�:̄�O;��$���}�\��8w=����S�n"R���Yy����nT��⩁G��ϑl�=|M_y{MT�����9G[ў�ҙё��q�����_�=��c�\S�pT���z�[ 5}����<ʲg���׹␿v��{�q��A�y�}�{}�#o��8�5�1-%�{I��:9~qG#�v�,z%*Xs�R>��j�yi�RG=���X*�n�_��x�;��J���ﯲ�ݽJ/Ǯ}� {�7�R��]O�݃ǚm�[�^��tq���(s5K��ߣ�֡x��+d�ϴ���W�j��s�w �p���/
�\G���}/��=�uw�{OA�7�=��?�Yl��� u=�D�*��g�t��z��E��"��xv�[9x׼3�]8���U+Hz�70��zPP�|�}%ѹ���9P��6�;����=M/O�p+=qv��X
��
q�3ﲸw�4O�����	�顾�l�*<�����O�잨����fGD��$�Ӆgt��S鼈D�����bu�G8�'��p] ���筇A�+��nFh�;^f���z�fГ���1nv�
1ff�2N�fM��ǔzs��FD��]z�Q��c���B�m�ei�����P�O�;P�=PtJ��M������\o�<��^ JW���j�|G�S����H�hN
�y�<t��O�]6��팙0����֣ �Q첽ꇇLyFmV����� �V�^��
<���箂��G5��ӷ��x-����,�J�3M��y[p�'����7�OO�m�:U��C�tJV�b���i�z>t��/!�o�ǲx�<l�C�2kK���L\k���q��{=O|Y;ۓ^��]³��-�x�;��7�c����l�ogIl�6lU0&�X�ɝf�I�Q��{s�[��ގ��U{ǆ��s�w#�O��Z���zƺW��e#4�K����Ks�H�_��g���F�&c�6S,~��	h��>櫂Nq��P���p�~ܥ{�������
�ܯY��4^{�<�?Sg>����F�����汿xT30��dfj��`^,���ޛ% �o�2=Q-�Gأj/��>���GFp;��|��Wi���ǕC�n۹�>���!�)���T(��9�����%qOrI�2�w���.
�V$�7�T�[�ׁV�?\%o��غ��Ie-�M�.����:G3�;��� =ݚQ������Y���F�weLE��ӱ��7&�{��VV$ۛ׋}cv�P���^��K7LJ�'t���
B���PL*��I5�O�S�ş��L~��~��ʩ�B��9 \y����TC�LӞ��<V8�4�ԭs5���{o��	��1����}8�{2TE�� TJ�h驇�^&<�:qC����b��G��C�>�r�'�[�_���.pG���@��5^G��ܫ�T��W��X\�/F�mn��9�=���\uxh��X-��N����=�fE��
�DT���,垍Bm_���D���@��.�{� �i�ɏtf׸�q|L��P�i����j�|E��yf������o�E<{����Ћ�%�� ��N�q����ʮ7X�L��Xx���F�5�e��#�췌�>�^v@�s<}��o�����n"}���1�5�^O�i�r7��J����j��{�ʽ�kE�N�~���'��A���#~X�*��g�_���9�ueSY5���XRV:���Ozpސ3}�!m�[d��|�̧s�}��r��S�)��'0���i�@����������#�:k*x{&w��L�/t�����s�������Whh���R
��N�ɗNK���o[��+��Ԭ�|��s�em���:�1{{�!��S����B�S�bO{M���Mf(؝������Q<]-6jYX���Wl �4\n�#MS�^!W�fT[S�i��@�����D�݂cY�X��ܼ�3���zM�l�� &��L�d�Ĥ���i����[.;9�2I�z&�>�9��Ԩjt+�G*�^z@�Fx�C[���S٠Ѷ��=���SE=\��N_�e�um*Y��>�ᓛu�%#��t����^�(��L�ٸ*@[2G���Q�Ǚ܍����4��I�\9y���%���y�s/�a���=�⋓�bZ6`��d��{Ǚ�F]��}P��X�~;���^��l��ح
��]w��m"�7���fA��f�g�O��0P{��<�X ����mv���>�c�~�Zp�[;��z�n�>�Wㇽ��q�����{�M�uog|N��\����6�.�Ӫ<K�L�������}[F�4�ǻ��Q�¼/�U~9΀��� b���_ek��z��8��W(���޲ə�l���m�/ղkK��7���ʄî~�d�+�`�}�5�ϝ-��9�o��G�<z�c�K���n|6�kC��������ߘ���;�;ߖA��F�sZ�����z�������O�z�G��򍛏~����:�����6�z���Zk�]��O�&���$��S�nY���Ij�{��ƑvyV�n�I6�F(����q�Z����0����ʽ�|�%�d�:��a,�[Ç��\�lro)��ݎ��on�Y}ˣ݇R�>�v6�"�T3&)�2���6�+�:��Ȝ�!wv`�Hf�{A�}\���s���r�G�j�_��tſ0)q�8���C��^�t����=�/�l���CٳZoz@�q��&�[ r�W���H+�,�(_�����Ew��hM��矩b{�����UFᬭ��㮳{�]�H�ی�`R�Y���������('�עg�ٳ��֨p��om&Ş��>�U~ɝ��@L�GL��z��=��_f�>#X��޶{5�Ac=x�	�}	b������a�JJc~}7��KK��\���3!�V�����]m�������]��l�����Gc��mڨ�欲��uL�J��Sjy_\���vF�s���g$�[֤{v�GyZ�=������9�O��ί���SA��q.�A�m�H��{@4�A==����Jڿ$@��{�^
�瞾/�?;c;�)ȍ����~���9�p�4�nfg��YN<�:[J9r�`c�T�;�����l�J�l��u�l���z��V�\���>l���׵���� ��7�'ޛ�@^ٔda}^ÐKGw��J��{�mp+Z��uЭ϶��nM�Y�\�^�j>�H\I]�Z��*y�LcV���cD�,���fr�Z�,;6o6tҳ2��q�z.t�/��RĄ�˹�^`y�e^NQ�T��LR8U���0&�l,l�oEIS]oK"P>�uҶK��'vr����z�I=�`/|�,���UzH^����]$8�=�r~;�>%�K�n<Y;����z�V*��{�B}v}�:�I��?e�n��F˨h�M���=�+L��\�G��$�4�/����]	���x����:S�� z�� �ωV{��=�9P��+t�ގ˗nz���;�֏�T�gJki��h�6v=���A)Ͼ~�MQy zʟO��p�ͯK������]�K�^�����\o���3��	_��>j�|EǺ����{n���Z-��ӱVc�]�#~��=���K��:vaY߱�G��ڭ:��}��*1[�-zs�/*���g��exfiM��O>Eg�����-~x g?m�D�b�쭸W�VoK}7�@ڈ�v��s��_�C��<���+����>��	\$o��\~����#��6lER�ɭ.�g}1k����})\N*�f��/+ћ=h�O���8�y�^G�ejJ%������S�x��~�5Y�P�M��Wӎ�*�N�}�;�9�c��:1�י�e{�ëW�{�g��&YRm��*b"�'d�9b"?/O��J{�Y�ZWw�*�5<���&��ؒb�Oc�
kq�'.	�@��N�f�3���&o%��ޔ����I\�E�������z�ںBa�jNm��α�����"&�u��d�����+ԕٽ3O����.�-Ls����c><�z3��M��ޯ.Pc�^���4�7U~�n�ng��H�Q�>'�o��P&)����J�u�P�y���?Sg#}�}@`��o�=b��p��9��]��^UC��d7 p'h��Kv�����\6o��>�����ݎjzn�k{�je�+Ok��{oף#�>��I0[;qJ�T>G 0���Ut����*g���wlǝ�Yw�W=IDN�(�#K���dT[�r@���6`�ƨ��=�,ۃ���ǫF�s=\��y��4ﾀtg�޶<OO�=��霟N �=��5~�\���_�u��WN�<������;�;����i1�e*7��ǰ3��,k~��r=Ҿ�s�z���
�;�	�t�3����������a�:�5��}W�ᢾ�b������� {����w'\��x�_o��c�˔�#��O�\��]�g�y�P�������&j6���w^�US�)?}�QX��j��ܷ}ux�}"Yݙ��뢍�	(��>����3��߮r�o�/Ǥ�}U��{Ɋ�3��[^�l��S�o��c-=�Y��ez�t��͒�Y��;��ؖ'[R�DO��𢋚�ͭ3� �u�E��7yb~HR��ï@�p�ѳ����'C4�G8���/0��s����'�3�,��F�!�s�	@��z�M9�3�t�8����̨�����7rI�7>�Co��c.2�B���+�^�U�*29���ڬ�^
����4�X��)e{=<ǽI�,W��<c��>��VES#�O�T�ѵ��'w�|]cƲ�l{(��̾7���T�nu6HO]y�ep��{1��V�pKf����'�\�٬�����k�UF#_g]1��=3��U"7w��s�g=��Whh%�h���(�G3[{{W嵞�?A��V���`Jnj]�a�*-��"y�����s})���$��*��/�:�e;z:���>s�Y�z@��+�,	�n�TEϓ��47�Y��Q��9@�N����V�̗�}�8����Zk�V��:r�>ϣL�ٲ��U#��D�Kg\���}1.���%��v��h�E�_
�?[f2;Щ3��k����Y��,i�������E��9//*���э#�B:��6XU��hR�KŇ��ϧ΍X����S7�1>�"�u,^��������lww���*����}KN|KGwØ������!��7��߾}����>I�-����v0co�`�6�����m�������m���cm��1���1����cm�͌���0co����m��`�6��cm�1�������l`�6�����m���cm�`�6��c1��c1����
�2�τ.x�(���������>�����t��$BP�TTT�UH��"J��*���)D�D����R�RTIH�*�����UT$�*�-�Q=���$*%UB�
*�"kR�*���(�C@hRJ���R(��(UTѕ$й�UD*�TT���*D	JDT)@�U
$(U)P�EJ
U	(��t�E$U*�T��P�v�HB(�  �u@mD�I�YjS%֐(MX&� �j40 ���M��B����i$�An  ܸ
�����( ض���
)F껔�����R��.=(���Rg^�ҊRJ�K�V�(����
^�E(��^�z�X ҅("U��P��   �Q]mZ -��J�[ �F��F�@ %l�A�j�A������AIPJ!��p  `��i  ���ԍ�+V�Z�2�c!D�´m�lkMj����j� �f��i���i@����@����   �mj�,�
ʊ������+eb�cP�(
U�d�B�l�k0�[f&Hfj�C#D��B%V̪TEG  ����V��c5T�&��� �`ʢJf� k@�ckS �D-V�J*څQ��ڪ�Y�S)�lKa�єʹB��DBIM�  �W�Ҭ0 ������eZ���4
�E�R�4�L�V��L
jکmUV�6ɪʪ�
0d����P!\  -��T4`�kE Ʊ����1�MDA�5��5j�����S[f¦*�c$��֩UFh`�j�+a(h4�T
��C� w1��h	l�XkT[0��Vћe�j��-+0 XKH�ժl���+Yf�J���jMV�-m�Kl�PJ��(�� ��B��FH la@i�� �lY�����m�l �kS(���U��E��    ��eIR�` � L  �~CR�M �  �0�xjm ���i� � )� �HQ�b`�����&J��OHhȓ�Dژ�����J���� 2h     bֳ��`�`0_i*B��A�� �hR$I�E��z^�_�PTA�bX䊊 �?X4� (
*�T�A�������g����0�#�1舢)0j*
�;Dj�$FA-D@���m{�g��˺��""�9Pk�R��7�5s�����i�B�����$��/�_�?B�I�pA.	�m4I�Z$�Q�*�Qe�B�"��Ʃ�ehP��j��ec���w�V�.�{ow)kK��«l�W�C|�S��H��{iE�wf��(�CsR��@�|Pd���Z�0��x��Q���R�!�ڠ�b��`,��(�;vLnG��ؕ��&��.z�T�P�D��t`��Rx��#�&nU�I&kM�s�S�a�{N웏(���$l-��8�2�#km+E*tD�	�
v~Z����2��"�ȣ��%C+lĮf����.���ݤ�/Wc���ѡ�ĵI�TD��umO�Rߣ��5I�Z�夫h��]�1� 	�F�N+�0�DT��i�Eqc��
T�*��D�`�qR�N�$J�nKx��p��n��Q;:��`�&�[�U�(�2`���U-<[Y%ݍM��q[����*¶��F��H��7��$ׯPlF�5(	5�2J�a��6�6F����N���阱��㩵��"ƃ����M�Cݘ�w��
L¥���FR{J��4�KYW��D�e��ZӰ�«)�yRۧDd�&&q��)�eKw1�͢�3&�KEH$.峑� j�ڋu!>T!r��P������,YYc
!Չ0:.[ĶPi�@�� �H��L�*k����bU�e����mX�M5��𝸶Vfan�����+[:�c,������ʂV�Sͷq�����T���̻�lZE9�c95��E�9���V��wmX��m*�;���`w�6擮�)��8jLB���g%Ջ�0�J����T{ـ?��y)|`�YsT/�ӯ7u�*���r0�R�5w�&⡈�sA#O�Y��cumR�y���v���AiuLi5)��w6�ܽ�� �Aa��CS&�Vm �V%၄H:M'��x�-[Մʂ!n�>����W-�!�#ڷ@@�Ml�V!�`�E	.=ĵ�/Y�B�+U7�4�K�r�Sn�6�2�wR�L���0٦�^�Q��ne�)h��I���]Y�2=Tu�ɹ�B�!���V�uu��' ��P�D*��.��$R͂�f	ٴ�@v��FoI��S�b��WebN�f����Oj@�#6��;�Y�6�������M&TL-^�pi�t]�pĭP �P+@E�Y��b!�����C���o�uy�m]��S`q��`V�r�1b�J��)B�њ3qf�@f�Z�v�x�����S�(�X�E���A��h͂�#.���dJ���H͎f�nmn5J�%�_�kF��`�wI����mK�#u�x�*���Wb	XF����l���a�Bb"�ICt�̣N��-�f��ǳd�N�J�v��3��K�f�&E0VGv�<�m)cR{rd˱����+�Z�p��'>�t��Z��Chء)���-30*����6�ח�o���;iJD����)�A��~ʱ�A��w	��V����ʘ���8�nΚ��^\%���h����5z�y1��Ŏ���1h�jmZ�˗z��e�3B�x:Ұbi��<�l�W�Kj���@f�%ٽϰi[*��bH�e�d��1�`�s3r5Af�p*���I�P-�ލ�<ܶ������P�V�aQ�b;˱�H#��4�ڛ���Z�J���*��HmE�n�3���oQ/D�,���Eۧ2E�L�[QI���Õ��[%m���o>Al6��wB�mZx�gsfʼ*�˚�J�+Ykb��f��H�Cn����TW*쉐�Ij���ʱ2���Xܦ����g�t��we��C�f�úƔ���GEЋc���Be�)$K�CE���ZܥfͿ�P�v�e�Pie�v(e�u7TAU�4�5�Y���G�p�
f���K"mmem�X����d�Z�:<e]A����m��ѕ�W4�23p���߀4�e�ܽq�vC
�M5���U�U�j,�D�b;�;W�q��^�T$ywv�/dT�VD�!�P���(����qKX4��`��6�WrQ��(�ӛ�L�p�R���� ��z�.�x�%e��(6fU�DtcU��8%�44�`�ۅm�nRSr�E�Uֳ֠D	��u5�8u�:��t��袶��+L�e�)�f�A����w��$�ڙC*1b7(<�$lK>�Su%����έ*�2�4��TPŇ@� :�aṂRQE*\
�|�!���ԫ������eB�3fT���IL�˛#a�5&�%=eE-4Ԙڐ��R	����N���T�R4�;�����b��G-�'j薲�iT�Wp�X�]�52�-�P�j�ʘ3�'H���M�l�P��]m�[�n&U0��j�G�bQ��e̢���hRI�1��ɔ�p�1f6�v���ɪZ��*�]�M��� ���M�D������e��M�[x������dQ�*{5���ҭ��jz��(ހ#4��F9CD�"��;�����ڑc�Б`F[�������E,�Z���H�)��Yr����
��j֗�df����M��@a4��Դ=/.ge�x��u���2�c@�)�J����l��~r�nĭurCA��_ۊ<f�FU�Ƌ�WX��KY�4\�Y�w�_�m�b���SJlԤ�r����9^�ֲ��� ɹ���1�IYVP�����E-w6���&[`W�`+�,`�d��E�&�Y�Bk�[FL��l��+@8�K��C20ݜ�[e��ՐJ!���f֖�h�C
��A�"X@K�e(� u�dE��Vpm�/U6]�Z��fdq�h��E*��&��u�K?k���F.��S��{YO�PU���6�Z�d������M��#��0�N�yn ��b`Y�-�6��nh:��y���3%��(]L��Jz1-{n[2�_\Ɣ�B�(jT����Fܻ:����цZ�N	G��p�45u�HL�))��UcRsN�MKM:J\C��Ñ��Ě�p�&^U� 7�mͳ $�nK#pʕ1�0�(+�J�s0�V:�k%�+U&-�9��A�zQ*(��Gpa���,ٛ���0�lc
�Y賾��>�յ�M�X?��H��K$VF�,,7E��[t�n8%>h^�X;�w�*��hdNHᱣ):	��zPj�юju�j���4f�ij�E���Z�Ij���wA�J`���	&kQ�^�gn�An;��iq���d"�-c�q"_^,oK�GY �{��5��-���(�c,*ܨ)������[`�4�g��Q塘�	�Xe�6� 0˭͑�"���w�.hٸL��e�6���n��eڍ�"��0"z�7,Z�ul<ƣF	[�Y�YʳnT�*�h�t�w2m��-�a��/�E��ʐ�(�w%�itS�Qm�����n�[x�l�-�6i쳨�b��1�H�`��Av�1�:��+MMi����ZX��%�ȭSsV��3W�P����kr��a�f�ŏk/�2�ڼ��J"�X�m�ɪ��w5^֭��2PSv�"�d=������Zڑ,ʵzr�8t:U�b�v�+Pܠ�5��O��l(�u�Ӧ�^&��`��7,��EP�I? �mݻPڤD"�h��3���5�X����Mݦ+I��/e�����-���MbR;�f��y,�yJ��K
���&�0E�0�Z	��޼���Fk�ӧ�dṱ�VnlOr�s0��M�`������YmݚMPB\-�l�o��-72#h-�Z���(ޚd;ǧ���b�Mx]Mj�t#���6Em�7%bj��p�x*`ܦ����UGZ轵(�e�6WWw���N��j�lM4v��nt���"U��"C�0���Ne�1I��	ǎ�q�[4k��6�4E�� ;�x����B
mm.��t�cy��$p7I���/rD�54�ʛ>�pF�ܣ���j�������X���6��)��代�>�%�@^9L���� �ע�47r�ZNY�P��褦�z5d+-��db���ōc�Dʙ���,t���"����%�j��v][rX͔��A-!�f'u
9x��Ө �Uݭ8���M�v�B�V"uF��YH-�]d{F9gr��jmIO4��-�f^��zșv�G Mз�e����SX�l-�(�,=��&��œl �UW,S��v�� �E&��U̽(�OJJ��k���N�m�X��Z��4�N��ځ*�t����nd�9Ot<[��9ZM�fc�p�MecB��+!Z*h�	.*(ͺy�F�)$A���z�4ͫ���$�t	���N+���PZ�,�fZ�sghX�Će2΁�u�`2�V����o7N�͉�ri���f�X�1s�N^����h35�Õ5���1mj�ͣv���SZ��0˖!�gM-��J��Xr!YX.��[�u�9f����b�m-eJ�F
9��N�N�"���D�٬G���7����Q�2�̩�0
��fd���5�_\�Er�v��7�)YClژ���B�͢+)�.jh���ol��
��vA�H�W��!6k���7#��ɀ}����>QEK�z�Rb���+i��hڬ� n�%�w7)�R�w�b-��Ӣ�;�&S�iԴiW��Q1.�bu�|݉�a`ب���6.�[�p��N���2�֭�dQ=�3r�������t8��Ӊ���	9R�jf�w�-�!4���rv��cK��� �s��F���AKf⾗���jfJ�Y�2Xy�3i��jh�(�Czj��Z�[�O.�8e�I�hTPͺ�� ި�n[a�jh'(*U��2��{th�Է#��V�x���&V=�anՑq�h=ZpMj���
C�GJ��2Ri)ub�4�l+����e8��%Z����fJ��m&�WFm,�� �D�V�r���n��$�u��j<ÚK�P:s1Ըu�@e3*��eRR�+ ��?^ۑ���e�NPH9K.��9XO��s Ip�)A�����V2���yA�̰�[�T�n�XΚ�t���)�M:�,��IZ�����	�R����UA2�df�]i6̤+1Ӛ΍�V�h� ��h�i��c 7V&F�}g����n&�i����$6�7OV��j�����ػF�κ��ؔ��T����)5`���F['ᙥ�#U�.TԳ�;�5�X�Tl��*�^4�Ԧ���8�����a�Ӕ�]k����$��7G W�=���n�C�VV8�[w�^kʽF��X�Lz��0<���݊L���ԦC���ۅ�;*i�f"^��A�=�۔�H�|�ziAc��ݔ)Y��Rf@�ߛ�{�a�ݶm�ab��R��H�ڨ]n]5}��Q^��1�B������iQ���zc���wYK^!������Mj�n#Phϐ���x�4�F��5&E�;{���8�\[��t��u��e k)i]	B��gT�eѺ۶FQ!_w>��X��.̷,u��Z���`���0F\u�!&��Ӭpķ"��A�沯H�6ЋU�*��N��@l���#Ee]��3sX�%��q�T/}�-���=���(k&��Z��~��Q�_����/�ѦԌ����$��$Cpƒ|���#��� �^f֩��G.���䒸䕎<��΂h�xV�ٔҠ]�^��0���B\̤��I$��6&r�g����]0��Wed��ti��=Em��e�x+b��}��z�Rk'%����:í��*�0��-3j���[R��ކ����y��|�I�Pǡ�sQ����������a�wlM���&�y�{�����-���uq��;D|�"���3�&F¡���`��H��<- �fV,;Q��*����Vc�yl`Q��sy�>�;R��*Ӌ5�mN�����HF��v����=�0�3zu�}����˽��4��:
21Ҳ�;\��&�(8~]�]KP�6�o��ޒ���N
��=�hٻ��Mӷ�vt�Rѻ�K��E`��L� y�M����u�W���V�-!Eh��A���5����8
5�8�q7W�퀝^�qq޻��S�es�HSwluc�L�1b�PЩ�Ve�\1v�7םP�L�w)+�1D����wN�ٜ*�Y<գ��*̔�����=�`�@%Xn�ض�w ڜ�wu��h��kj��%C�7޷8#l8Z������k���d2���WG"Ac'f���WQԄy8�z�q#�+����O��t�8��'��:3�8��uj����ˬY��$a�b2�G�;dX2��siT�Y�4����s�vR<;��dMY�m�wK��q i��bY�o.-�-Jy�v��OK�dܸ�۠p�6�$gQ[;T��m���|�l�kNF^qT�L��N�ɝW�Ī�Z�:G�l�W4��ClZ��Y{����ڳV�&;`I��|&�N��="�)��rvpٸ�����JXh椾.AEh�w�F)#{>�n^��� }Ѫڲ����aP�)���օ�v8.L�u�5��蛐���fݖ�bɓS`��H��,N��S[��6�i�\!�g3�ɳ�eVe�[dΈݧ���:*߮�g(������f�Yb��o+*uB�bHo�غ��sV	ө���o:n�jvn�Z��iu
�+oi��H˘3��Ҧ���ZEaͮ����;o6'*�jn�|3�vP���qϭ���V^�|l�\G4r|-�P�hG�kK���f�����,�βi�0i�\^�� 5yy�s]�G�O(�J��Q1���U���^rJ� Uj����t��3b1��T+�T7���ĖasO�DY[o�[׮����fQ�[V�r�tkX�k㇙��ҭ�\T�j�����vf�Xi��w�X��]A��u�9�[Լ�s�*�c�,�z	��Y�[�%���`f�/gk��]h+:�;^�	��z�+IuqB�A�,w:T��*J�T��u���s�]A����ò&�wY6���*gmR[w�E2�٧H-��!R�2�=��b[� ��L��n��
��W8�'[�R�osm� ���:��ܾ�r�j�Z+&Q�4��*.��$Cl�
�;��\�7a��YZ�mu�s����J����
4j�q�-��/z]��l���F�[G*v�2}ǘ��8��<����4,sV�.��Vژv�o�d>�f٦�c��DV�t�Պ�3�/F������Ϧ^� ��+���ݮ����ɪ�	���Dw#2�k���.v�Bv��qН��d��+H��/���]p�{�%C�*;�.\�]�;���D��n��W�:���5�k�fY�3CE� `���ݬ�C��8%K�>}z����u�t�m-�N���BtCv1]�-�:S�e`u
��ʲ���V���J�l��-+Nf���G�qkC��u_&�,�۵�iO��m̤w��3:D�.��kU�1����nor�K�iPk=�/�o��PN�@�����eC�W74B�co�:ދkT�j+�;U��{G��ӮH�ok9j[�fhX���)ݹV�g2��fސ�t �Ǌҳ8�}N��n�Ê���	��r͌� ��ɂ�6��nP@od�V6��F4=�Oc�>�w���v��Qb�(v7N���܁_p��ķ\��M4�M�=���&�
��SwWk�=o��n"QwB�o&XV���螝�w��uj���+PH���X]b��iS�m��ϴIl�K�H$�@�-U�9�.T��i�1
:7�U�<ǙBGӮ+kL�P�ro��Ώb�f)YiDNގ7[ӯ����N��tzQu�9�����P3.�M�0�w@�X���:e��7���Zj�.	^ΈB>S_RF�w���B�v����Ң�8ȁ7�n�(om�*���٩����[�K��vM6'�\yc����﷙�#�)��Q:�jv�R�A$α�����b�:۬���2�i�;��Y]Mu��*�Z;r���P�&����O����O���qؙO�U�]�ǜ:��}6�3'J�QBw��k3����0�#I;���e�4�f�5�P;]���I�+J��N�U�����ie-�ӛp¶ܮ�ʄs��w�_kGc�(�J��^�r�3�+E�6��<z�zU�N�-�4;^�pƤ���/^<X˸ƴ����OuU��]ͤr!팏��ʇk�*dY��&���]���ނ���H��F���V;]74��Ŏlov�!�qi��2�wLЍS�|34�8.�SL�sy��WGR��f�ȭ%��C�����Ω�1��������us8�H�����s�V�溯&c��Qqb�k�7\v�xn�ة���	���z8�F�^�nu��-���K�6®)�����C�������0�ލTHOebʹ��"<N¥	�DlՊw�6��
�V.�|V*<:�D���mV����]�a�8L��;�$���(6�5ҍ�/(�e�!d�wv��[h��f��xzYy����:|��S|���q
��v-�����!/v�=RT��I.m[V�#���gncT��`��})J%�4�.g3�,�5��2�`&Ś�{X��7����&3m�Iֳ�#�������-��_V>�=����J�'�/�'M��N���Y@�h����t�!�أcegKn�W��gt��ԃ~T/��}�/5[��nt)�z���R�[_]B�@t]�s__L%OGK)���!�<��"`r�>������p`�S�/�u�g�P2Ty��RՊ�OJ��汹���(�}�<�󒫍c�b�2c���>�[]�B4��j���J��T0_�e�6�����vjB:�ӕ�k�:��R�ك���s*6�l�*�L]t@̰e�f��Y,�ŀ�������*B��I�"�ă��3l���������5�i=Q�p��S���ڌ;c]�u���������.��v6��ړa.�(Tbvn�Α�{t��ף�yX�|�c~�'l�A����呜��G:H���J�k�t���kU�W�H��1g5p���bO�b����w=��[��xY�i����s��(j���,��p(��j���^��Z�f�אnQ��]�n�z�U��֓\��v��n�%�ɑ���� �@���d��a�^r#��gY���t���o��z����w#B���G�w[7�\Ҁ�{e�Qiɫ�[��9��p�3Z+)�z��s�'��·r=�rI�F2z>Q���t���"���A[���}���c��36�E|p�nFDeU����N=vX4�SŔ��%��v?�:3��ַ�1�!�u�n�ښ	[9��{p6��lԈ��r���Єx(�5���*x�WJ���4eo	h�4�`�g!9-a���A�)���MW�+n���>M2�6Q�ʋ_i)�k�䗍�u2��Pn��;��̕���h��ܰ�Y�;�x��(bS�͊�>�ֈf�پ�r��������@f{��Sp�+P.���\�M�)is&��=�et��y��`G�j��aBwt��-�邋���IuY|��Z2���(Ђ؝�Pm�VF̐X��U1#%�4Gn<��)��m�F���jb��̑M];�S���Ե4��ܫ�uZ�t���� ��Ln�Z�U��Y�����'C��{W�,$,�IY�<����;%`��9(=�!b��jX�����kzԤ��˩�v�N��F�k����;S~7�C�*Nf3�pb�A7X�}����i��Ev5��૕��s��㚞v��'��nnR{�[�j":���w2�|û�����|w6��b�^�2�'k%������W�ټHI�3�V�Ȼ�6+c���凝��Y<.t��OU�ru8�����O�{&1��n�+��낼���ݻ`RX��opu9=�*a�Y�jsB�π�l���˷N;�\\��~��Ƿll,�\Wօjʇ��T�ӑ������^*�/L���+���p��"^dv{'\0��Z���Wj����2�t�fA[R�̕�,z�e��*��G]I�0��0�p�"z����p=;�o/�������	��$t8�;�#$VC��5t�}��@rs&g0+�6�*T�҇juJ���[�i���m��uzr�Z��˿����YK�{VL�r��-��W��
���x�a�=�&-�;G۱}�����e�*qC\sJʱA>��#k�`Aء�/��A]�}���h�W�u��l��ݝ����&>�g{�_-�6r�ظh`:�/��1L��u����V)ђP��R�A��������ڶ�G ��.l��{`^��[�2{Q�6�R�W�4�v�G�WL��ܛx�[�wuk2�jH�v��ƥ�������F���YytWb����Q˼�_.�@�M���Lx��-;��m��A�e�ƬviD���s������oUt�mtW���ئ��[�E�db4��t|�{o�sP1.l��X�V�F��(K������hxj�v���L8�R3'7�U��u^9{��3F�V���/&U��\��Sc2�,<���5C�Z��NgV�s;��k�q��X���(�o,��;������ �V�K`ك)˸��/�����؋��Wh�ky^�T]'Db��j-�5�Dou���.�9���N�̸����)j��`[.�z�%�:�\�guռu�6n�{.�jg�8L�R����r����Ȇ�Q}@r�Ʃî��䷶Z����z��S㪥���V̝K��N1w��.[�"̲��S3GSws�p䰇-,۟r?u;Ugg��B�Go$��+�q����xF��Ә+��*�|_P�h����ކ1����x��S)�l�j�2oj�	Sb%[s�8a'����������>�-��`�i^8z��XPv�n����SX�o��aA�5O0\�r!یJ�MՖ�Ih(YH��\��W_v�f�B�,�q�M�f۱��G�Wײ �>p��h�s�ו°�M��E��6NWǊ���s�.�'֑�U��ӂ�F��MsV�c�W#�.�f.����ړ�}v��M�8��7z������"��� L�K��k)-�7���y�&�f�s���I�)i:�f�m�gn���W�᭝����'
�8TC���glf:Pذ��ë�ZU�G��xD��cF
�feteh��r�G�˸�a�3�:�
1��HP�|�>����]�K���;Ow-��=*�xn�I�^�,�E<�ϏR�{$å��
���Q�c��+�C�Y�5P����Nb��訓��������,X9`رC��w9�YM��moh"� ��!���ؽQ�2;��� ��r;[�~+�[�����Ǵ�cejQ����G��֞��׆*p�,���U�Jӥ����*+�w�SB.ն3w�p�:�;-3�G0t�N��,铬���
Pe5ۓL���t��#e��Ô�<����֊�xpo���W�jE�u��Q8��㹮踶b�vZI��G1Z{�ʢ�|�U���I��,�Z�*�DSbt�\��ͱ�V��Y{���	ݍ�a��5��̡�m��ȷj�����6J�����u���ws�������V9f�̕�r���v��ck�s�S-�r��WA�c�hU���$�K.�M�L�.��:gm�(���1��PQ�J�i嵟v�İ㳔y_Ja3"{o;��mfV�}�a
��H����Kod�o�S��K�E�����ׂ>P��β3�f`%:��%�^�&�ܢ�ۭ ���Xݢ�
`�QH��nnIr�9"�8]���]A��k�;{WED��Z��+oM�a.,c-�k�[�r0��ZG�oR:��3jqB�M�TF�=i]����4x���$ ����1��V���9 ��O4��O�]{]M�c4�}Qv���H^l�@����ɭ�h�j��ˀV��0���.4��D.��ਢ�FTO�A>���Z�����4z�z�}�F��0:$��<{��`i;J�N�U��m��lS�.�ε��݁e���eZ��udw�����K�fLG�`oa�N�����uI���OE_�;�unS�TBi��5�;�v�i�����Zt۔l��¸
ŗcw��F�PTi���h��h������gZ�o^�|&��.�,Í�++r��KU�-�t�)ΣQh��G����3KK��y*�%7|;cA�J�kw��y#�:�D��4.�*����v�}�	V!Z�2h����������_�$�W���Is���Gi��i�pv�4��/�t��7N��W6���Z�Jb�38�`N<rf�ܥ�p��Y���@S�2ť\�1�8IûMY�[4�	K*�Qؐw
Cj��˫�Itg�+�lŝ/�Ww��f��Ms�:򐬬�9�ɏc�Ć�K�P��ׂ�zll�%X�a����d���MP�&)ZKzN7�L	e�t�#�>�a,�20��a��&�e�kv�bAc�-P
��݅���jҕ��
�sO���S0�}����V�x�lt{!]���X���%%�D�)V���_f�����3H$�Z�^89�Փ�r��r٥9Z��8b��jS�hP)ۗS�^u3�e�ܫ�g�s�9���X�WX�ΛF�ŏx��̑��V�}f�00��Zgl�q���[�Sk��صZ��FI}B��`���M,Ǹ%�8h�iޓW���`���w����<yb�\�
C��&���{2l�S���Ǡb(}��&�:�On�l�V�,5$�]��]�͉��։��Dx�$�S`=��^�h=Ļ�|ڮ���h�y2��,���դ�k���	C��c�y�kY���i������c��@�.=��N2똑t��A����.h�\m��nѷ�{�e�&�yBR���6�hq��QݎE
{ENf-PC/�l��w��|�:êE�>���[	�j#1v�
YՏ���Zp��$����h�+�;fA*ZmWq�+��
�E�(���[�SR{:Ѯ�[�ҟNU7�c:`�� Q��ډhem
��и,��k�����in⹩+��N���
�r�*q$;����c��I�Q;�ԓ��Y55.�=ֱ^؝�pð�<�w&J�b�_K0��3�*{K���6��K)mS��L5�����> ���H��I�/�P�f�]s��Cw^5�7�)G�{�-P��p�R�)6��� t��� ��ۙ� �U;Rv��TݎQ��2ee��˅��{X'U�n쳗ek�4����S�⡱^���
��S�C-�D�0���m�xQϜ)���Y����Pu;�����N�y���0����iL��[N�+�<;�3ui��]������fVŬ�]֐�9g���<��W:ђ���4;QUW�[S����q��=0�;]ά�l�؍ko�GO9�&o�i���de��+��6�DKq������.�����wø&�^D�m:)�Y�M�R���峳s�[�zs�5�l!1S�䮝�g�ns���$��FoU�].�6!Z(͏�v�:�]1vV�EXR��hZ�[6�8�y��P� EC>���iD��]�h18�.H�ǔ^���ں�@7`���bHcٍ��!��ӊ��{�mJYش
�ܻw�0�KM��𣽻	���ɥ�,�|�īGq����|D"Nv�6uǶ5>r������i��� ��
�O��-�e�u����U��RcNm)� c�W^��]�p.�]HP�x:�(��sA�[�c�XK�Y�ZTW#$����YsuK��ۓ��r�9U��Y�w���N
�딫we�{ϋ�+*�m
;C6�2=���g�+�֍�b�ǜ�J���V
��jS�u��֧�F3���Tk��Z�(v/Q�宨*ѤU:�ڳ�R��i9���$��>�R�7�5�r^Y����K�С�F�*�N
\���t�),ZI�y}�$�!��>r���iR�ϛ��V�Y8�Ѣn��gEutLU�8�2���&��7�Xs;x\���Z;�Z5�`�X[���o)
�ג@Z�W1�5D��7�
씲�>'#Ы]p���3�SW��!��rN���S�u#H��׷�*o\�$nG\���D�cT�
��L���r���\p5�k;�1�>��V��Na=ث$�ބݩ�}N�ő�ĝu�%���<��31J��a�S�2^���yҲ�G��^�����1�N!��&���f���
e�՟F2U�_uB��ֆ�����si+�vx�qL	H��C֥��בovq�`$���b�D��a}��J�q���9�Q޺vz3��Ղ�+�!��ٰ�m��\ۧ6�K���	�'Q����<З�2b����k��9�
��D��tV�ϐ��&�_��N4{��˄��L��I��I��wmY���}.Vv��ЩcZ6�p��L�3�}o�]�gzz��%u�3��-�k-6��Q�Nw(��/�*�fm��1��bݢNt�jHp����v�6�r�Z�vb8IW�-�h�L���4wqmY���m�ǁ�4�"u���Lu�������ILfS�O���V<S&��w��q��3�b�H'1ʞu���i�z��<d�Ii�ekT��P>�"i)J�f�דP͸z�����S��:���R·[��|���\��Fs9��D����L�*��z��9�lC�-c���: �f+��d�Ƣ�4�fE�p�Н�{���']2̴�[q��'�Jچ�����ky��8g�
H�
׼P_�{L�G���U�����(14�[�ܼ�sS�3CGz����F�d�bn��F�O����ʵ&���&�OAw\Q˻��:��
��KB�m<՝V��knjFw]�)�&�Z,wV�����}W����T��[�Gx7�J���V�L\��re$���
Yx0�u���C �����2:��q�N�)�Nن���N�^4�d�}��0YDiЂr�ɹ�c�}5�%d���ؕ�]�)��2Vj�(U��v�����5�iv��vrO��͢K���-#ev[
�c��@V�e31FEb70)�4�+.����c�zN@i���P�:68��h9�%�"U�+L��w�]*�v�_]]��̄�)�ei�Ԍ_MG�)&8���Q���67�h雪f��`�VK�̕�`��,��j�#�=}|�A��k�e�dBksٺu���a}�u��lBHe3�R�׻W��Ҭ�H��1Ɛ��u��q�s�,Iyܭ�<�hCN��w|8�96��K\�-yH���r%�i��ۗ �w	嗣~
�]�l�Si ���uBb5�V5�� �m������W�jƻ�s�{'q��}O�����ic�eqJ�Wg'.�7˹��ty^eX�e5z������3�y��{���d.�3f3�J���}����=�Ho5Zi�p���Y�v�M�+6�E�9nT��]�d]��-�Y�����Ô͖��w:uZV�P�g5��<
�{�.
��<Yhhg�	�E��Ek�{�7�S'T���-��c�mi.ٙ�Cʺ��������:|V��qD{a��]A��QCFn�^��vr����/�}iZ9y[M*֞�f���]N8�珮�8��%
y2=Uw�;&��ô�o'i`p��-��ʽ��F���7hE���A�C���F���C}����R�ր�]X����3+�ܾͷ��"�	p���ks��Rh:��+��FLf�f�GM�ԅ!����\�}B�,G/�f"o��P����!PU��{�X��(�+&���t�T�@7l V�+��I�5�Ӱ>%<;;|��A]���}�S�.%����l�Q��G-+�}B*�}d�GA76뙅�9*iy�<�k{{~]�V�W\�_2��$Nmmи�VK��ЙC5b�ҧ�ۨ��1y���v	�(+I�j��Հ�Ĝ�[99����I陚L�I�f���VBc���ھ�;y��2gDj�[\�6jn��.������ZZq�]=��S�!�Ň���w!��ϻ����<����s��Xk�ML�>�P�_.
�q<��]7
5;��u��¬�X�ҙ���ٵ4�r�WQ�L�;���Z��.�'b�V���sX����{\{v����:���2��Nq�t[�t�.�\��j, #�F��B���!2S�u���V���]$&wJ��n�෫7x�%�:�v�ɍR��1�{����`
͙��K$�i�Q��_%�ڻrV��]i��H��t� ���Z��.z6ԑ�T(&�YD��g41�*��T~�Z���K:)+5��.�m�	X��Sc��J�jnnA\��w^�+�]�>����//o��}�E:�\簠��nX�PR�*�\;7k��Ac;x���}�;f��o�临��f��+@��︺�9�hA��qo��΢f�Lλ�yJ�����g^�%���>b;s&����ܻ{;+$da���v��k*m'��6�Յ|�=�s�M\�d�E_,�{^�d��6v�YeX���iX��nb�Fn8�M��2���-M5n�ȝ��3,����_��w>�G�8�t7�)F�7�¹���!j��<�V=<�ݎ�J5���rm�o>S	��&uД�V����e���ul-�k��[���kn�^3J��W�f��R�^�3�Q���$X뫡o�y:o)��R��g!Y�����iS}oD�R�1�B��c�O^m�K:���l�t�g+�X���uI�1���e�C%5�ګ�h��Jh���飬urt��IJ��';��h�Ehfi[�옷uk4����C�y������U��3�t��*ԛ(^���jə�\8]C$�IF�L���T�_*�u�n�����-��6��*$*�wMPa�ï�)
+l�W��]�Y�1|	)[������uH�Taɴq�*��.�,M�e%��|��]f�,nts"����D
v�Q��Rgf�A�K�lU�ۻֈ�˞�w�RZP��_%Z�	�N��f�M��� ���'����i�vM~���� �>��l�@�
t���5�s�.g-Ra�V�t�[� 3�k�@E��b�{���Z'zLH�QIv�][n�L�c3�l/o��LΩ����,���������ڰ���/.
�žB�/��Z��wQJ�1հ�ʈ��}c��<�k�*�+�A��R�^
��]��ި�wm�5ё����M��|+"�7��'¶n9ȋc��
��i�46�F��E�H���f�I�<�&��Yƻ -a�@��J�6̣v�BQ;s��:���w"�Rd��33��ѦLWǬ<����i���B7nX�Ǎi��L�����2�n��soB��"M+;�d�\+��ڵ���\үp�\�����og:<��芛}���6v��ke��We�E*=m�m-{�k����1ˆ�s��wh_@� *qÎ�`�V\�͠򳯩$�C��F�� �/.4ki�������Ej�ЩV ӗe*}�۽ɑʕ^�jWXc2�]�o��9��X5�9=\������<�7H�HYzh�@�p g)/3*�!=�L��ԎaZ���}B�Τ{d�#�=w%�G	��I��͈��ju��L�modi��/��XP���v��_Q�9���p�S���9��j��̜���(�6��S>?�������˻���v\���NQQr�9C���S�j�Ep#�H���bHwt�Ԣ�"�ݖE©�PG�$��E.��RkI��x<nET|2��Q$�3��W�7wrN�sg�L�<���wp�6�*:s�rBs
M�W��!��UC�Q�<�=�eAQUZ�żVG
x��r�Ի"eʠ�\J�V%L�R��M�.���Bjs*5�:�ʬ�UUDED*ˑTE��j˅P�i����*��"�S�&�UYҊ��κ�K)P�9U˔ZԒ�*5C
"" �QݡE�(���5��#�#0.�9>��������ן_�_he���x7�L�+iU����@Sʼ��!�Ϟ�E\��B3t,���Wn�N�{���wIڔS�9��Oy�OMz��B��+�m��ەS�-\��OֽJf��Z��Ӆ��JB�Šc����Si�k"ݛt�,g�oW�^�'���2��@�F��V�"��us� �U~��ks�`o�T�ҙ"F�zRI�����'y\#����a�TН[dǀ�U�o���g^����A<'����P�	Nd���t�*z'r�5f��1��oK�!�at᪣j�J���b*L���[�`][��h6��w��	ۤ3]�Sǐ�3;��j�c]e"i�v�y�Smr����h5G�"N�mds��8�W>{c��hg3��{�|鬵-�B�x��~3�{��77SH�AYA`LҒë�za�J�a�ư����U�nU����K�����=�����:�,��>��Hf[�Y���ۭde��7Ρs�;bgM��q�m�y٧-�%��|܈]_n%�u{���J]�KQ��1��Bb�5�\y�[�����u��0׭u�+օNF q���o�"���v���ͪ�.��OzT��.�~IS�Cd\�P��C����(0d�M��Ofu�D���j�T�\}t��`鵆=�����Kӯw������]�>]5l}1/]K�T��sOUG3�1��NqZ,�Q�vWT��N���7����_gH���s���D��Ρ1��^,��Bt|i��*���e#7�s�	"6��r/� �p�7��F���>6��X|������s��	���G����/�5�t\ꋾo\����"sYLH�DσL�!2
�v�G8�5�����ak�a�c5։Z'���m֪ٶ䮃�7�q��`à�����[��ꏺ�(7y�ֶ���W,�pu��6N	Ϛ�}���6J�ɵ�Jc���':wNl��>C��$}IP�s�`l"�9����N-�n�N]�3:��L��3SK�����n���OE��R��pi՗GD�k�ʚ��}�.Sk9EFwLs��#B�ZgB���<i\,���R���)�r��CL�_���֞T�����Љ�p�`�X�S[�����Ɗ�%y@��κ��i��Qn���=�ԗtZ�~�I�q�ᷠ��3w+E�oYW�a�˭�Y��}�5%���_�K�+y7�Cb�Y5�3�k��T�u��*V��1z�rS�-f�IdR���.}�C�a��P�w�X�T��F��]�q���u���Ӻt�R0{��K<�Oh�ͭt��.�c�c{�9��k��c\�j�fv��l���_��8H/l��]2�띧X�hg���K��^hP���Q�Ku]"�,v��J-����ij�[]b���q�$���$o_n
ndɤP��m�����۷V�NF^b��gV΅��t1��H���V��6�Y�Q�d�3��3b9N��X�g�O_��g�=G��$[H����eף�P-9�WSa^n�M�+'�ja��bu(<#��)�b08�����ݻýLɕ1L�\W�����J;���!#i
]�����X�Ri��#�o�X�hZ`�=�׾�nhfɛ��'�v�@:�R��ŀ�<W���N�o9\��uXys��h�j�5�ڗ�0���}��^�ioJ.T��8;�|J@�}R�(�|�\�{ٳ{yE�%m���Bt�ܞ��%�=��ĸ��ò^��
�s��!�,ԏ ���őA��lN��U�U䔸���b�H�b#�a1��GB��{�T5�rt���d�݇�ҡ�w�Z���^�*���ݭ��5Z��g �v:�N�=��	`������k�1�n(�9�{R���]�+#�9�:wKS�Q�3݋��Q${�>�������V�Z��q;$�鞩ׯ�������*����^z�_x<����Ov`�e��g�w�>�u�昿\L��P8�S����u:"*Kآ�Uf�IJ.^7~�qf_t�D��^��=^�� F[�W�|������[�un��䴌��hh�r��c���f9\s�iE�V�Wu�v׃��i�[R�\r;�^�W5*}�*���f�s��!Cvk9�;ڄ�x�a�V�Y2��L��}S�+��B�rl�F���D����������_S]���KT?:�2� 45Ў7&p��APhl���"�����I�B"z%�&Rfa �G/=bm���U�=���Չ^2m�ن��/�+9�^�4���1��Ń��u˳�cYkI���N*͜��.��n��gg����I0i�a}ʢ׶i�{P�yYٵ��'i��:�e��ZWNN[���Fb��	d!��υ�W��@���Z#j�jwB���<��O9��S��#�[Y�џ.w���;�hf����uY�����w��a�%�YSꞟt15I�\�8.n��T��#�6��8s�i��5�����X������{Ϧa�|�� ��"w��\d�X'3�\�ǳMLծ=��yn��Fd��Ė�+b߭�y�&k�"�d�}�6}M�H�sw��%��-��*_.��t��t���#*{+d^�#����]��ǭl��K=����F.�B��5L��xc]�f�x�=j]�]���c}�c爡u�����hǙmtZ�B�=F|oiŞ��:�:��Sr�T.Nf�;z�X��Ee�����e�*�."��:+$J=���E,�W4�*���M�핋:����MT���x[�Z0�	�Km�'���aҬϱ.��"9ݮ��樳��r�b�E�>
�
r�uꚻ���̢�&���ؓ���+��4n���Mμr�:�b⤭�R�m����.�C���>ħy���nw�]1iM�hi�[t!ms����HJ���u��Q���^�BU���q�����Gs�}�oS��+hSf#x$-�d�`�z�ήs-.wIx�Or܎��u��>����ա�+�A�І��u1�����I��Yutg�[�Txf�R4���S	;*ꡧ��,NMc�q�y�l�b��U��-i�~�HSQ�`��hܒ��]�#�t�_�&�Z��r���"�:�vm	��7Zޕp÷T����z^#qu~��/x������h��]lgk4��t��,y�<ع�kΉ��s<�`�:��^(>���={WO�iĺv�9�ռ��F��d��j|a�w=���{u��=ޮN[]l�u_��Z����wvk}|z�r���I)�\&�(�G5�F۟.[���/�jz�<tх�q�Y�Ǽ�DK�;�j�M�w�)���b����T�5��K��c!IݰU�T��3n��s���Z4��ǡ�άKKYW��J4�$�tr��.w�r�w���u�Y�ϻV�K�U�Y>i�[���Z"='�r�y�X]�S}������gM�p�u��"V#"��������FG5��s4����g%J�)��h�Q}���k��?u`�f9zu��i�X�ˍ�.�a��u�k�:��G@6��jQ>�D�6�U�4���k��:o%���r���B��+}7�����*�*v�qP_k2!� �uq��8j�q�W]�S5=���* ܱ
+/�*�IZ���**q�%9��u����y*6v�{w��t�V���y?�w�/��*�kv���nd�:�5����7�QfA5�]��m��寝�)�7&�q��2t�9$�
�~��eE+0՗@��B&�j���Js�٫�*Nv�ޅ���q+��o�7Q�|L$4/�/�V,ܜ,���V��N��2�:�X�l4�P�P;э�e۵ӯ��iM��,06�׳y�V�*��זvCwwx�"r'��U�aVr+r�#�HW3V�u�+a�]kw`��Tm��9�U�]Kj̆d�s#�n�j�BJgs��������Gj��T�lD�l�FG����5m�sO���ae���6�Ve_0oW>Æ�l�WT9n|\���1x��nO'�:f�N��[7�V��;�`;�Ä��V�~-j��q���.�s�(�|�+�kq�^����_{�	eg&�Al<r�՗S��k������:;7=yƭd8h��rL$�+�J���L��oW%�]���EQ˻��.�\�;�e�ߕ��n���\�ù�f��ßNw֥�kl,C�#����K��$,�E���F�wX�:�i�F������W���w��o�ɾ׽�GE!��y8�,�U���svH�bը�S�j�<t;��)�+hk<\�V%0��\^{"��^�,���ޤB�!��|�i�r�p�Y��	��� �}o-�W��M��b�9�a��f��Ֆ4b^���Zb���j-\�-p���5R�f���#�c�e,[R#=�6���ޥv��5��R�j���1)�j�ΪPó|oo#j��BX0�hʱ���![B��3��j;�	����[�#�N�q��/�*.��%~��ԧx)}�+�N��S�}��H�N+o�����W���E��F���k���Ї1>�|/7���MV�m���_b����I����lV`z�ۊ�,�͇��H:��kZ��/UF�Q�W]0:��	A�YgGQ�G:����T�\���T�㒰��#/��bѱR��Ey[�nj���TF��'۽�k�#�M���
E��7�E�{��v����!��Әx��Ic��\(�̻���Ь_b��v��8�Wt�+V�R���*��dkdLzHګ��U�S����l����5ܟܾ�]��M���Bi���C�o����Rox�N�����[�o���ou����=�2;\qR�;�����}�+��NrAG�N��y���$�J=k_R�_\߬ڃ����֜T�yת��&�uj鱉:J�{�k��}��K��)�Y�@��6*�ܾ�Q&��j9V��s�Ί=���S��Z��X,ԫ�n�^R��:�D	�(yLú���"�+w1D�o�c�sF�B��iőC16[+�x:�\�}��AȽ=�\��X�q�F./�
<_"}��luY�٨WT
�.X"�� �LƮ��k]1Ԯ��u4��ܮ �i��!�/;P�B��ᐍm�����Rg1\z�mP�:��p5�!`��ΛQ�����3]����5��PFTETX�k��mp�k��9F~����ҫ����|��*�t)���:�lZU��EZ`��˗R�V��I=�n�B�A�J�h��f�˼UY��a6N8�TI�f�U?5J�*��&��9�	��cn�7m�ܣk�)�w������.�i?�7��KW�VPP�|v��/D�A�U�i��WO+Z�Y
���0�V�^��#]��l��t��L���j�$�D�4�
z
ʈ2�\*_�6u�,d�O�����&�*VQ�� :è�kM�����t��Y��j�ּU��H�e5o]�PF� �.�6�PL{K�7cB+`@qVZ�!
f
�,9�^�n��7��\z�Am؀Yӳf%����йL�scUrюSW�^�(�3��Wq�N��,K� ���
�Ij�	����*��T��e�yºwf\���@���u�&q4��!vL��}�+�,\Z.���:��Y�8.�E�kw{v�X�F&�{�rQ-dgXQLsbwIq��h�,�42�Slw�S3nNo'n����E��<�%��y�����tQ��]Z�5p-ͺ�M36	��s�Y�f����*v���;῾�rA �I>�)�Tj�r�$������'<�h���J�z$Tr�G0"L*�BF���0�0��"s*T�9TD�ls<뻉ݕs���93�E̐�5<����Lꂡr���D&��U�.L�ul����g#�,��
I�w:g���W��D�&繢�*u�)�)���g+#rv�sps�Q���PHIs5K���Z�P�r�qJT2�$�Nt�$�T��ECk�a-e�Y�19Pj���2�,&dG]��D�s<Ȣ�P����U�%k��NKu��h�5�$I����Ii\���=]J����u�Ô%hbH{��T�tr+�9
�te{������a��N^�DA#��4	P�����s����z:8E��� ��;9�������͜k�ņ�n�����ԵS�3v?�.����r>u������pJ�Q��5���i=�p��k�5���ְ�K�ӽq*9l��M���YKy�'�l�����wM段��H���+��\y#&�lMv�uV�k\]���P;7��}�M�P8|*���fY��3#s��j�^ q�K=��>���mc���^��l�����Y�cC�CQ	ح�}�q;�����U���S�"��\��2-yZ����-_��,3��g�y�k9#�:C��muCx�AH�ȅ�V�z'�+�߻#�3pN_Sc��w��U����$%45�5ޕ���d�.ݮ���dPP��}`�$w"e7P�|+�F�*��.ԇ5V�?�����b6��)�*��d�����v��r��r��X:%W�U���J�T.8N��`4�x}K߱?�7�ثYd���>����&[����Ҝ��c�,n}���<X�M��/*��O�gv3���ݾB���vgk����{3�����{�^ȯT��T|��O��]=Sm&�����߷��,�݇��i�`r���L�����7j"�nf�J��U9|����q�z�{(��ĪGa+�mǷ��T�@��c[2q��]�kG-M�������[)-R�ֱ���w;���G[��jJ�M�=/��)<�ξ���!llP��4Ħv�u�;x9-W������n��BY{�sq�#d�`��hGi�n�_s�����=<�N��\�o�[}�l��-���,\oF�Ww*6�'{sy��K��V�V�?4�1S�'}��S�߬���ݛ�3B�	g�+�kP�^�
��/j�;r1s��W����t�j�����������BL�{�����_���B�:��㚤��eO>�;!��}�V�S2���O_-Y�R�"�=W�������w�Z��}|l�>t�NNS�gyȑT�9U���R�Eg�ǕGgE�s����P$	���s�u�跕�5O;��y�.�����R8�c�1��+���5s4J.�R{�yN�6��ub�t�#Bo�[��V�r�5tj�6[n]4x�Y��H� �螠n�4ܨr�\pط��(������c��,>.%�/�US�/�f�j㩮o������x�׮%4W:�҃(T��5�670̾����}
�Ws�Xŋ��;R9L�N�k͆���^��Χ#�C���z�&_N��Э�p�����i[�7�W��j�q'!d�Ʈ��5���UDF1��`V>�7����[�l�.ml��\�Y쬨Sl�}�GV����d[�[��A��3uY�5�<y�n|�n��/y��d�.���<vu=�G�6��v�\�S��t�q�|x���W)K�zI�bk�X���B���rmak�L�j��x��ٰ�[���F��=����,�J��Ԕ��z�.:�$G-���u���J�$)U��wڶ`�xn	ks!;Q���.Æ��Do��G���& @��酗^}S���S�����oi�շ��_�N���]����7��?��0x�-��������ǀ7�vU�"�>��H�1⚼*�kwg�9���o�o�����o���c�}q��;zv�����o������6;Տ�� �>��,��|/� y�� E���}�*�8k�W�$<޾�@��M�ӷ�l�o��~�����\zM�.���u����>@~v������o�ީ��g*S�{���v���w��7�ӏ��vߜy>�M�n:���ON�<F����������]��|q�?����z��oN$�߾���x�������װ=�o���\~�����nq���~@�x�>-��wｔ��o�{�|M?����ӼA���2 '̀��O�k��ޔ��� �8�?c�)߬{Wm�<Q���ϐo�����l~v�x�.7�g���o���zv���|vӿx���}�����m��K��K���dQ��<8�`>�v����M�8=X����>�~�ޏ���ۨ?}�o����ɷ�g�'���F�ر�\È����K��[��yL����7�xC�>m��}M���6S}N��}vӻo�?&��ǃ������9;���8'���������?6?Y�6���[�����g�p̾Y��C �hA��®�-�/y�)�=eeg�ߨ���<�C�n���i?���{��^+!M��9���J�/9����W����<�켊�,2F{��r�y��"�bNL����||��� >�y[���������z��h�x���oɿ;oS����۝��ɾ��+���W�����|#�h��v������
pwߜoN��(oHyv���`��o����ߝ������D
<=g��������>�G_U�{�����N7������~v<�޸�����<��{oN����~2�;��{L}C�Y1�mL��po�XH-[�u��(�t~lL�vm3���z�����k�kGH��Kk�l��2��k��m��{�X�ɏ=!ɲ��v�����{H�kb)��i���r����{�~�����X<�o�<����{p|w���&ݏ�zw�c���}p��c��������xP��}� �����5�������*�Lx#�|(���S��tG��@���c���������|N��ޝ����Ӿ���q��'>��}p���Cu�Z�wR�L�q$�#�}����@���Ǎ��o'}�����)������o��1�����P=�����>ϧi�>[;�fOf�)^����^��yBq��.�>B��c�`����@{@���Ͽ��7��m�?���~py��o.��\o?�yڹyk�����G� ��^�0���o�N�y������]��ފ> {M�ɼ��ƽ�7��Ϯ7�� ��>��/ꯈ��!�N�%�����������<&? w�c��]���l}v���������`�FޫM`��[֋�C87���T��ݍ�s��XV�2�Y�.�įZ�on1�
5���aiњ�i������<M��o7�c{u������]V�h�����%ox[����V_a��Ƶ������VU��')����ٗ�s��s:CsV>��U��u����t����|B����l;Ӄ�p��x?&����S�����"�~>}�`P���[o�<~��������`��O��޽{=�~�WW�|��}�I���(���E@�϶�������~v��N��|p��o��>|�>�U���c�������pt�%��+"�H��N���moVR�)���o?��]�&��>;P�x<���]��oɏ�=F9��6]������]�'�����wϜ������������u;�x|>5X���>�B���6�VHyw�>8�q��7�O.91�7��cs��|{�dN��ނ��#�i��w��K��'ou����@���x?}�������d1���˽;��X�_���0yC�~폨onӷ�@��m�7�o��Ì%�%��~ϕ|�{Ҿ���>�{r�A����<�?8��~��'��P��߻o�zq�cӏ.�ެ��� P��y� �E9���~��W}s����ߏ��8?�C��h�}���}O�|�< ��������N�܇����ć����
pq�`����aO�`����\wʥ�� ��?[��E6����۷����}p}d�}��㿓�����>&��Cz��?!�����@��G�>��y�+W8��8��g���Ǥ��H��~���&�y����Cշ�o�����7�ɾ��������A���?'�ޝ����6ޝ�_ޣ�.>���r��O���4O���|�+�=��뷏?x\c�;o����m�������c�)�?������>�"�JA�UK�����}��n�un��溑�����]�X3�>誇N�[Z �kü�γZ��Bm-ؒmR�)�o�p����.����'S�p�xS�ヂ
<��%j�M�s�����;t=DKv�r�j-\�9�;s�ս/�-]��s�e�#�JD�u�[&�]!����6�ߓ{v����c}px�=������ {���7����������z���QDL��\�yx>�>D"=��o����]�ސ�~�?!����o���~M��˷�@|@��ǟ��6<_�G#��ڟ���&7�1|>>�ɷ�]�?��n���P<~��yL|���ǟ���������m� {v�����=��t+��wt�r����t����z�yw����m��S�������������һ���7�'o~��6��lG��#{���}�-N��{��o��c�)�v7��vސߐ�v<;��ﭷ����ۍ���o�]t�2<Ͻ$%@��vfޫCiN�V�9�]s��٫�\{�d{�b|���i�˷��m�������l|v<pO���|��o���zBN�cb<d<6�:�(�	Uv�����_xBo�܇�����!�~��c�8\yO�7���4�;z<FߓN�������m�1�7������v<�<��7��������~"��X����､��X�~���So���Ss�ʔC�q�-T�+H�֊�چ >>�g�´�۷��Vj�𯇽�ޒ_�q���!��o�ձ���v���<~��������I����_8]�!��������<�~}���ߏ><1'*�s^�Ӓ��>�`Y����X��7�o�����������?;}��gߝ��7��<��v	�M�߽�bp�H}�|E|�u_UN�5/��z4�y++*�-��E�_词[vϫ���L+�W�y`��4`nЕ�/����g4"[��q곙���Mq�*�ܕ�>�Z���+/�������9"*���[��K��a1%��3;��;_-��C���_�<π��>���W�^��;|M�oA��7�o�������=�����zq�Ǆ��x�������?�ߤx@�\n�3�˺_g/����$A ~ެ����������v�M��A���1��c��o�}q��~O^P#�����Q��ûN���?}N�3��z��7�;�~����?�B�=l{C۱��;yǯ��oI�����m���m���`�zq���<|�>&?'��z�:��w���۟���"O���_@y�&�SH��E���	���J�	�%�(��������Ǵ�]���x��~�������<^N������ۉ�{H�#�����<~�������~M��ݏ�o��C��o���y����>�{M��`xq�����}�" _=����uDi�����+��Y��{�{�����d��ɼ����=��!�����SS��on$=o�����.ޑC.���k>�H�3��۵���L�{���L�x�o������7���6��.�n����>;{C���z�0$	��O��@ڨq?�|%u�)Z�~}o�P˃㷊2��ӷ�?��c����=��������o��˽'����z��7�����<�s�>>��׿W�߿׿����4���e�����6�h�ޫo5�������8<����}q�ѿ!��N	�S��|����t2������_���<�Nσ>��܋���������}q����M�i��Ğ���8=&���v���>��|0�y� �6xi�������YA���Q�c������9C���φ�0~T�N���Vqw��w|ZN{�O��ŵ���F9CP�w�	/yQ ֑{\D`׼������C6����ܔ�hޮ���1-Z������>G�?���s��\��|M�78�����8�����ߋ�����Nz� O��k$q����&#6�]��W�x���z���������܇���|v;�ǵv��A���.� �]�Gｱ��q}�����|��o��O���i��8S��U�Z��{�}�:}��Ǐ��Ǵ���}X��}M�ߓ��c�o������x>}��H�����x|#�8`�{��jn����y�V��������ݏi���?��ۜ}L�>q��o-�	������zv��/�m���w�]��?G��v>�����Y@�V+�K[��O�A�|>���c��P��ho�α�����;o.<tc�׻nv������o����ߠ��S�|��Ŷ�z�~���=x������[��{z;�#�@�\>��4C�����ǇnMϓ�(o�~����n7��?�5��m���[|Wm���7�o��y=F�]�Q�ϯ��}<?_�|���׼o���V7�?X���>;�G��8���m��y?{�bpw�=��������Hxv�_��7�?�o���k�ʻS��i_��[*��ȏ��� ݿQ��������M������S��ie6��m⫔V�mVA1��zC�c�N�{v���s�ߏ_}~������{ǟ��������6�� |M��yM�7�o)�>�-�����oO���q�N��x>�����������;)��xk�%}�+�j���G*��y�O��`xa��U���Wg�m���� -�K6~��Wz�)�T�o�6k�:���/2�MRa_���B����hmeY����F=��?�>�<I�G6GסI`'�,c�����ޅ�Տ�kB\B�m���C�j�̎76P��$Y{'TR�\c��y���_W�1)=�މ�_�]w�h�T�Gi��݄�m@x��dV�*۾��ZV�F)�����R+�8���x��lĨfn�|�t�y���|�����k���m��G9�P+i�ZEFjGe�̧�K�S:�u�Fvz����#�yE!�au�-�]�:��2�jG%+x�*xm_��d���������*�'wr�֫�j9P�s��7��Cc��0��;�V٢���ϰ�	��ó�N+[V"i�j&�OqmN,U֭qPX�fD<,p�5���q2�	Z�����.+��v�}Ј,JhӮ�ĵE���l���୰C���2��jnR¯d1m�Ex6����_�Aj��1�o�g�2�h��*����ɏ_m%I����a�7�տ%t��V"Y���8�]��2��7.G!���`���sރT�]�7��K�>x٨�t�ކ�i��=�2)L��W^��n��w2��Nt�;��_V S`�Wg-6���\�9���R���W��`�f�@h��J�_Y�e�hT��WoF>c���Wl��bj���-8�%W�nf�,u�x��t����_�L_�B�̭�������,댝V�9-�md��7��31̻��#F��6{N��JN����[v,��T�����1Tߜ@*|Ӧ^eu�=;Gd4# Au�r�묏�����OH+4m������j��5���j�F�dr���K��߅����wT4t��U=�w�q��9l�l4I�f��w��@.﫪97WX�&�=C�H�CΞ�<��+���5�	��۬;{�8�p��N��udya���yC�i��R�gd�&=�kt���Ň|6�/�mQ�x���"���Qtyt��̈��ȝ�s�=�2���W".@��(��թ;ͩ/0	g"f]�{I�tL0�.��y\�+�MT���ύ�cy�[������9+ƞ4��ܙֵ���E۷r���2XkUK�t�����*�Y�`���9%$��}!�ݾ���-��,
�&�>ZJ����6�GJ&�����]&C�a� (���o�U꺔�ى$����gY;�呥���J�2����I��[�x����.�K)G����ul��m�ot��i�RJon챵��ҥVz{F�T�)�4��6����Ģ	5lȳ2X�����:�
�!�X"���#j��u
�P�fДOX���]WV+QB���h�	�:m���wn� �����Jh��,Pz�ݔ�b)�ǁA�˒7q���$���̱R�
�J�W*�,�0�U�h�v7���k�U������G�/���)C~�Q/dN�BJ��̔vGlm� �� �y����r� ��,�
I<��YB�[��Zt%�zel�vn��ֆu�x�ȵ�ι�x�b�����ݤ�K\�;z����yRWd8��ˤ�nxzt]W���T���9[)\�,ܤ�����N��s��;�wtv��o	[\�U��Com��e��Xm�鲏_"�u�ש��ױ�o��W�W<h�0]��3bȗ���,��*�\�!%U[W��~���Q��>3 �2g���t2wΔj�����\t���\�KC��Ue�B-e]�vp�$p��v�9��݈�](4�ۻI�kRws�4B;�jT�ET���IJ����EU�*�E�wr/ZL(��)������WC�2Η�L�÷]�\�W\'"�ʹT�Ir3ܲ�y��GaI+E�E���[����"�a#�ȸN���I�']ď�R+R%���:���ӥfr��[T-�q4s�:f��"<�*�.�9�0�U(�#�T�CSL���4��-�Y�dW�xTY%vDD9&`�E\rO����W3+�w"�(*�<]�"�<W �,\�OA�Oa�N:�XE�r(͵�wBPFj�����EQ�\�<G?_?�����߮�_�o2�S����Z�q���.��� �Յp]ͫ�'E�op2�ܕ����_��=�֤�d�Wۃ��&lS��S��ho��֏���������Ǌ*sX��Q�|�N���5#J�b�J��fv�Vo\�o�w<�%�Ә�~����W�KC/�C5����KY��`-*��휾��ъ�
��:+ѮEB;5�o�=\�(C��m����X�4�Z��;��:~�������-�O\���	��7=U�O۩�����/��r8I{tr�Z��'F�֧���`��]�Ӝ�ؙ��y��mRJ��=����Om��Yk��!�o+���>�\�	�څYZD��k����Z�Ћ�b�:���!e��Gt�n����Uy�ȍJ�q
��+3��ޮ/�OU��}j}/*�_S8���R��]c�K�i�����r��Q�^Y��z�5m�3�_�qΕr��ݷB���H�m:7*�n�!�	;)#D)��-H n�,��̵k�]	3�pAf#�J��V.�Q�d6��ݥ.�>��ͫ��ڵ��ؚ���_��{��|��1'!AW�O��_Q��V�i�X�6H]���/L6inD{B���lϡ><'����s�jl�kj��qt��İ�bfWZ&zf�j�K�����*�z��Z��7�Q4��à>u\��������,���݄��	�qp�ԩ����N�S�Mb��9�l˦��q��D�=ג�&Ft������>U4�j&�����:�!5�k&z�[k+τ
�t"�ܦ��f}x���"Hu��C�M�7\�-�S�e�_Tt��\2ofN�Ce3�w����M�����'|�gr��3���ʣ��V*�R��3������7�����/:��J�.���]CcL�%���4w���n��D��$tMm{J�T�C+o�K묏�;�",1,C�Ol��t�
u�&�5)��|�ݶ�J�:���ܟg��vva*H�X���Uu�VB�<Ef��O*#F%�K�����gF�K�.������\�\�:�������ӭL�.�i}uZ��E	���a�m��u-f�|5zl`f��jkg���	�1Vu�.C�y>�2�ގ�Ǒ�r8�d�d��W�9yhwn!;
k���2��4�B�LNwD�/��hiT{=�Ǎ,dss�/V[ҫ�<�>�b�<��������J�45�q��*p)�.qo5)C���c��ǡ��R��S9�B]��,��1�Z�;/�kUkFqt����@����qPZcC��ʝ��}�n�7���Tgiw�9kJ�_k\�E���.g���η�F�H�G��dO�����9ꝛG�������k��������:j|ի�|M���9s��8XxЃ8��;�/&p�>���9�^�7ȒQ����_����uF�YMQ��a݂֚~��̈́���V=��r
Û�ԝuV�>�a򨛠�ҩ����9����f���Hv���n�^.�;nWn�]1���{����>M���2�t��S�|���o���QV���Pr��Bj~�~�'/�&�t5�f��� �W^����^Hl\��uTL�P���_���ݸќ�j��O���[֕����U��qn���2-�S"�=B1�	KZ�v�Y��ܖ�uA�t�ޢ�{T^بR�lGi�t�b]X���E�nM�^G]��53��3ь��;:hr����4"9P��뜧դ`pQq�c��F�oi�>
w�_N�CrC|��z��_�����k����z��xv|�
U���/$4���P��}�V���ū�V?Dr�םYy"-�r�!Ԡg�D$%3���'=y��.�Y�2��VgP��a�h	]ԛ�"c�h��cuz�T�������r�yw�T�Ήo\ٙ�G��hl��C庨��R�0[�A�bT���K��R�E�2�et]Kǣt�N��gp.�mGY&�uИ�l(������-���я s���N���꣭�ފ�f�?F	HNq�{��+ŵU��}Q7��ߘ�(HլW���^W��e��x��p���o�ˀ�OY��(&!����v��((����_Yc�j�"�z�Zڒ仇��u'�nV����|po<{9��A�5x�F�Z�|�7�
�w=��1WmO9L���X�m�9^|wXT��	M�OФ<��|���[��d���x�#c��AKQ&0t�&�������9u��2i���	��N��U&���Ou�+�_x��t\�M�br�c���gQ��d�{}/2xÃ9*���ϔ��6�3�ݰ�n�� r����\\ܬ��9���yݩ�y�N�6����da��[��y[�1����m���V��8(���CvJ9���TY.�}�Wyl���b�wէ,�~��B;��AhD�Б�g�]�q���D�?gGK��{�R�ն��;�̉��OW`M>�<�e����������uv�o�.��]9޾���:���OyP�A
L���JWm[S�>�~+餤V�V'�jf�����"�\ev����	m%�.�M���+C2#r�u@�[�r���=�����J�D��w�}7A�sHi��R�M>�L⡏$�["��iƱ4��)%<���A�z�8�Ι��av�,Mq��W��Z�Cg���$&#��-3�X��#/#�x�=����=���W�3�� ��������-՗��ka�*�]�sZ��
��p��0����C�nv�2���l��V;�y�r��rqq�u5*rr�X���S	��[)e�3*������U-!r��l�&q@��!�B�y�V͎ꭨV��=��MGFn����=>뀟"�� #�	�\�����M����W8u���b`��՗��D��O���	��������u]F�̽�x�7�Kk9�j�Q�ػ�3�N�du���;�ם����=��qu�t^�.S&���Mt�M�B.db"�i�J 솓75���^��t�xd�Y�JZ��|���Ob�*��󻥶j�)�oO[U�{�fC��"�j�z�՛T�EN�ӹ���y��	{��K�y��˛�b�|p����d�*_��]��:���x�u������N�,�Z^v���j$���]K�N췛�X[퐐� �;�[=Q(�}���;#ckҘ�2��bĎȅ�>Fmyϭ�3�h#zrZ�w�(�����R��6�qt1YK�<�j8AM��v{x���~}�bw�������!>��@��ǡ	T	�q�1�q/���-�Qk�a<�Tf���A'd��R;�2fa	~�V�IU��+e����H���l�X�-drН`�y�U�g9T����"��K�9c�L%�^pt���fk
t����p��;�.�q��p��S~M�[0P��nv��L���r]��lG˲��f-����N�p#\�F��N���jMmf�Q���V�VV._ �����IΤ���A�7�5@`��QR����iPz�8 m'�Io8�<�"�bq�������U]�
j!�y����8��X�7eT�%�fCC5�U򫬥G�	���[�o�L�f���d7n��@k�͇�܆����F+�S�*"8�엓u5ى9�S�c2)ޛ�s�K1CwX���2B��O2R�B�����j�J�Ü�u"�����y���b�ԔKmzy��{%�*�ҞN��p�O��)
��ͤ�C陶I��Kw;���fKKc��?8� F9�ȮG��x���%���k���V��x�}�:F��aHq����эv�4�ի��9Y���V�b�m�f�KC����C�y=J��o>+GCL�w,l=X1�s�m殨̹�k�4;'e�ɝ�J��+��Y�IX��K%�;�)`Ӯ������I՗�q���M�.�9����Ӝ�j�S��n����}[j6���f�<�P�$A���]���F�za�OV-GgϞqx���
^���m1a�%9��<��p���{���j��tg��}Ʈ�j@�2�'}��[s)7��W���[b��T����3�� �dNl�wE'٭>�j����f��qliɞqX�ڟX�D��KI>�M�ս��x���Ȩ4��VX��*�O���J���ԟ%��l����z �3��ľ&<՗G�j�E_H2N]�jf&�ROZ���s��`�0�8[ɾh��[�ٹ�#�ڊʎ�V���҄�e��b��3OqR�	Ӡ�u�xo;N���g��I����Vr��3}�/��H�o�e �2��+\�����|^�YBQs���S�6����:Gh�d���3�uܡ9C�C�N�Q��3�{���7l��9���a�����4�R��+i1C3����]ʰ�+
��9Q��nyr��������8ow��˳)��{.�?_U���VM�3=��c�ka�9��.�+fߟ9�"��P��#T�@�x<��v
;�Z��ӟ��]�g��_ޝsU�IWdy.�N{X_^z��di���4��iS�]D^M��9�o8M:c�!y�X��[q\��(�>z������l�}�[�Ί��$�^��]�lj���K[�ż�,?�4"3i������gkڢ��׎{�-.���Lr�o&�7�P�"7l���Z�[����,�'����{o�&va�'9HJ�hi�#ML�Ux��8��s�q4�˭�M��0[��0-�'�pļ���OL鉾�
��0���
��.���!�Ti����q��{�y}S�Y���3�z�=��
h��I�P;֐=�kT��z��}�\�v<9�iǣ׳:��1Q���Q�2k���]o8���F�E#�81�-pyPj��9��1�R�ʕi��@i.�z��� |^K��7ME�����]v�Zǆ_%�������!�v_ƫy�<굺�'V�㾮=�:[sY�w3�	
��y�]X�Sk�2_�&Y��f�v/d�nnVuX��ݜ=�kd/^u�C�&:�X�3N'��_K�GR�0Rs�}���Qs�ͭ����XW�o�%�}W�:�t��T��M�"L㫇Y��mebR�?�ݭ�FNi��Բ�e���/�DPӻ�K����3h>Z�K��z�{���ǹwr���-��hyz��Ş�B��.U�-@�2-+/��kB�K��Wu$#hnb�]�(hQ�ι�u3.�]��%�ϝ�ԯ�qC���3!3s��0����Y�ڠr�	�i��R"�ͦ6;�+v�+�g_`k���o�1+��y��n�ɱ�*kw=@Ve��0"��g�|�t�����[]f�7�e��JC9�.�TR����zZ�r(�, �rG��ul�U/3(WbBλQl27���2���e�ST6�ot!�)��rʴ�ve%v�B�������[4}���rJ�YF&"�R=4$6��gT���!�]^`��A�B.�E��뿛�9i���5� <�Gp��5(����:~շl��a��
ޓ���+Se<W`�d*	�X	���F�GV��c�h)wd
�-�:3 ��L�N�J�N���o-�j�*;L�G5�1Ջ6���Y9Iؕp�>�W�	\�m���3e��k������"�����+�J��U�Vd�K0���[
�(4���g����$5Ձ{��-��q��,]�y��pB�*<y{]�V�2��3�h�y����>��#;�漗��kRab��Wi�`��[��v�*2ۖ"bC�C��X�JX�l7`e��,��e�Vh?/QY9 \̝�6�3z<��9��_A§K��C�"�����>:��l\�%�,\q��ï����&�9�F��u��T�2F�[�鲏L��,���/���z���	{8LV���r\vb:±Y�"�BS*�/����RwL�A�n9�d$�Ri9�s/0��!2(+�*�ՁQ^(N��4
� �$�q�7u�5��N9RT�T\�:WIRH�<2�Ww	$9�ܗD' ��9wQ$���8z�.nN苣YDr*�s �\�)�):��uC�t�wL洓��U�]az�wB1qU�*+�by	�K+u���:��W)˖��xH���P�f�E���d�e����\�z��VL��ЯD�^t�j�""

L�Zy8Q{�� �U��w.[�^��"��;����sù�p�9�T���U�躹�z���ē��=­r=dQ9Ve�ۗ�3*�![�s/PŊ�rT("��ԎFd��Q�{tC�2]�']r�ʽ�ķv����)͑fTTu4�"�FmW�`�=]�sM1�S��Yo�L����|w�v!�{7G,��Fڽ����x:��"GJ�[V��Wܿ��{��ɢ�b�{�8�V*8O�8���K����Tn��Eo0���u�W�f1R��t�U48v{TĶ��wPC���N#��&��j҉b��N���^:�R�fN��ܴ9L^s4����B�Ƴs3n[�]�NE�b��3y��Pq4y�i��*�W-WS�[6��>��Fb4�G(c��'e;Uػw�Һ,_c/9۴֫XT�NV�,.E*�`ޞ�Zܒ낟�is|͹���ց�z�e�fl�w�\� 0`S|���'�gA1{{)wg�����].�C��;u���9q�LՌ\̱P�Ҟ�"_+�sifߵ@��9v���U���Ѝ�v$8I�3��T�k���)n_+u3�j���NC\���NT��f�9��]lT�1��j�a�VU��U3�!Ly��}�3&1��}Ӯɵn���fG�bcJC���lR9�
�.����&��4����Ί�\�gB��g�m�[�/��ò󝗎��X�ִ��Τ��v�9}��xx�}�]6�+W*��S�O'v��K�E���;l�s �O�)�s�}@�VR��p��=SʠP�E ���V�Bٗ-��>�V�W#������d,'�Cq(	R�>B�5�+p��a5X���=�C�P���"xv����L��ݞ4!wT��C�栩��F�Fo�:j�D
�C��Ysݖ,�D�n�ӷk���h�9�3C��;Y�T8�
�W4'��􂁉��>�*���5礷e�x�֪U*F�����U"����W��$1v婉�nCV�_Z��p�⫍r�q�Z��-I�J�.�#���lE��\`ݔf��E��Pf�t���`��Z��SiIE�35����d��ґ�C�T,��,,��qf����k�m���}}�����g$�.����aUN���aX�_]F f��;F%@����^m��J��]�!=�ѫ��Y���xW˵������unTѭbxۆW�\Eޡ�+��3�o��f���{;���<��U�=U�����C����R�4���y3X�7�S�]S�Y�����-�8Xҍ{T�E���G�
�"���a�c�b8ֹ��Y�bCO��ۊ�M7��Vl�J]�<b�Y�x�9��ts:���y�{w;�z>�6��5Ӧ��!�ζD�[���Q,��1zY�Fz�Gz��uzÌ2����f�`�:�?��t1����*_M��J�@}A�Po҈!i���S���j�wW"N�4`�U^�Z+
Ε^��/j�3Ј�Zʾ��Ֆub�jfH�{��C�U�I�Oβ����]���¡�u⁺��R-G�6咁a���M"D�T)����F̨r��23pf;Ր]�PGU�-kzQ�0�3:i�f)�dO�eAf�m7�f]5��υO�C���LZ�=C����1F���]P��i���
� T�fk�מL4�Edk�<͋�ܽ��d�*p���u����ƗM%%4�v�(��u>����Zq��z�Lm�ޞ���F)WY7�qv\���ֽm8�[yG�dIb�yBSd"�-q�f�Wd3"8]aY3g8:��A�=�ܕ���%���9�>�P��,��t�+Ǯʇ� ��0Z�6ԓ�״����X��5yk�T�V8 �Yu��Ň�E�L{����l�k]��<�4S�ȃ��Q
��������*gƞ�FǞ�D̋�lw������8b�U��0p���f�ę2��t�C�CzY{�������X�hʭ����0�N���.�sT�
�ej�p�]5� �HO��`iX��1���Y�W�':Qa)e�֕#6�<mP�!9�#�Sٽ4��s��&���1�d26�׮;��j�ן+e�-f��v�.h�k�ՊԶ�6�Ύ\�}�GQ,p�%��4tk!�K�-����kY��{4?"s�g.��|k=��P�����&�+�-���a�R��^q�e�����t�ʼ��w��}���:��ν�G�S�G��&�D~�u.VP�xUrVT�e�sC0/+������Z���(��k{��O�	��ݯC�@լz�b���sh�6��㶇5�:r����N����_{����Ụ���F����q8``��؋�t�b�@�����_["�\e��R{�D#ŇD�uq�;<cC�$*Rt���gFICυ9��m'��"��/�w����W�^��q������Z�0��L�U�V����}��������H'���`��3%`���B���	FbA�C:6`��:apL!1�cB�Q.�����d���qQw�����w�AC�G)h�i3�ϗ�0�-X��fʞ�"$9h�"���ݤ�����R��Ѧȩ!y,���EW�J23&��c2QV�tzt�X�3q��a(ȗ�e�YK"��o�Y0e��f25�%R�?�My-�G�	�ٝ}���\;+
<h��Ƞ�+�+v�!��-zgRb��m�o^�T�ko*W E���uqF�]i��x�dڻæ�T�;��y�^H�I8y�hh�(8I���Y�r+�[�1bU�5G��9>la�3���)�;��wsΣ�6����Ʀʙ'�^º+��N�uhS�P�<K��`V��RI5Aɶia�����f⬮�L��ڼ�!]����1�G�8ZAu.�_x{��9��U����g	�ܩ$v�hŐ�Nǧ�#��p�
���f�N��Ə;�B4�ěL�ƭ�6�D.�ȱ�_i�u�3R���4���R�q�<����V\CpȐ�N�B!�`7;<_����ˇ�.Vq�v}k���N�%S��S'ѱ��c"$^�Cq�Ȍ���<aE8e�Jx�e[ާ��R�����
�V�P�;MU�b}j�,��VX��9Dײ��ӗ�-y�M�{w;T�l���t<(�cz#�p*�p�iI(ȴ'b+ҤA��։l&��;��7|/���#��Y����d�W�וa,J��7�-ċ�*fKL���w[ٷ� [IxIj�jƋ�l(@���z��'񮡺k�+��z�F<c"`��5�:ڜ��Wc��C�w��E�e��d�RC�or�O4�mSElEY�&A--4Pg���2�e@F}�U�6d���Ï0k�ī&��ݫv��ug�׀��
h��Σ�����So�8蹽�(lU���gV;w��fj�z\�,�m,Ԋ���y����� �C��	Ǘ�OT��
�`�n�E�r,�>�1!��"��������Uq/
=�ۢ�E��e��Ϩ�+:UD�NY�Q�� �F��`���4I��IR������p�<u��k�l��dS�LY��q�}�̡ȩx(�V-��e�����ε���]���^,H��y�M�ґ�!ǺՅqƜRΠ��U���މ�g:o/o��y�"��3s�F���Bܲ��\F�
+|���,�GUb��2��r���qQŃ���e쭺T�*E�T��qu<�>'�c�k�g3
�}H��E[Ջ�)+(�(�^'MoO�G��U*�>7L�D��]��wM��X�F;�z�G�zx��F���iK.�'�W�Pf�@�#ŀ6���1����%��'�gN��U1�hc��Z��GZ��Q֢Y�@b��C�;v35ɼˮ�������p����"ٚ���}��My�s����2�N͊�6�?��M����Q�U������
���}gYB��q�Zm��wy�l�
�F+������O�N���;�.�waĺ�ͻ.�w1��h��2�4�uq�M�2�X\��)r��͚v�����N��{�k���^�?g	Q%O7*x�!�3�Tp�6T�L��i����J�us��'�i)"y �bh+hR�f�)����{(���Gg8a��[��1n4�����c⁠>�Y&�j��u'^�*��-8�|��}��3�����v�TU��}K%#��.�
�P��/�_zQ����x'Ľ*��|�FZ�sd�Z��z��3� �CX�2
."|��3O��!��ZP�e�5[E��;w�R�P�3]ԍb2�Aǖ�����ʋ��0u�p�.�\�>g���25#�qg��N䢆E�If�މ	C�1�A����+��{wrƭ=6�rH��el�|.�y\Ez��u:=�Y�\S�D'���ŏnO_K�E�<���v�0p���S0`�(���w��&o6��r��%{�s?d�N0�9涸�S�x+����Pº&�A�7Ԅ��B⑛⩅3pф^d���������cBz�q�A��FM�4�2w'<���R�㝙e�#����
�Օ��XX��qVfP�!X��ׯ��W+�;l=�m��d������^���՗\����=���j���0+�f��P�Tν�2�Y�ћ97l�
�x�&�x]��Wz���~��o<���üHc�ȰC��(�9���ٿ8��"7���̘:��f{IPe߂%�3�p�X���>�?l8�[�|xg�ty/c��&�e+���Ȗ^��G��N�><���V�+�[���J?*۫׼\��u��6�;5%:��r!��ѝ���R�vL�������5`�Y���#���L���|��z��b�g/M��_*B��,&�#g1�>f�e�z2ߜ��Ӈ_��T�P�D�Ɉ�o��B3@WR1R��#n�/j��*J����]���r�T�bS�L��HT\�BF�R��[./�ݏ;����=��|)��z��0dVHS��mHE��1	Ը��LD�d��i�I��#0E#��c��%N8@�����p��a"���a�hM�Y�yV/����R�����s" ��H��l��4l�R�������	���٭���5Z������#L���;�e��L��[�v����O]؞ۥ��ya��ݙ����� fj��F���g�L^��1�^/	H�E��.e�!௻����������4�
b��ȳƚ�Yԃoh�)��f5��@�/7vhfF���4�Se�Z�P�^�3�ï)gy��\��֫��j������zv4�3/��5k�^T�>�c�6��A.wŔy�Pɾ�å�`�T/�%����b����	�V���2R1�:S�=���[�|;s�r�l˪M��k�!�m
�O�����[�j���1�+�3�5�Y�o��k��盻���a7^0S4e'ȪW�C�o����ұp���C��>��&l���t�����P�3}#�O�TM�_�,�1-��x�g���]]����-my�ft����U�2ᘠ��͡��Q�C��k��ܠ���Z��JE�����t���Y7j��w8G��g�өa+�=[�g��Gw�s-=T��t�e�g����2�h���<�V�Z*��ԕ��Rk^"�.j�g�J+����YO^ve�/�:"*���(��۳�kH��A$��\3��Ѭ�E��cp��!'	�ԧR�rT�⣙�#}xn���& �fJؾ��J��&^d�5&F4w�;�0��gv��$<:�(\���N���U5�9M��_8��b�6������ 駧C�õ�Q�x$g��K,��B�`�[�R�׵��C���;������&�7G�nا��?��,�֕��	���Á�+�)��6�p�ϧg*�G��j��L1}κR3{�EBX��ޘ�P˖7s�7:=w�R@��d�(j26u{(��/J*��ц��0�.[J_r��:�q �Scvnh�d_,!9�f�8��2����@-�9q��M��22i9t�ӡmV��u�����iB���
ܮ�|�.V�S�����ߗ%�G%ܡ�T�N����֞V-�yQ�w[Ρ�����c�3"�:�λ�W-�z���}�}�}�&"�@��S��v�NvvN��vEVJ��"(n{Z�\��;>T�Z��R�CGN�y���6��`q��H���V�
��E.�F��Fyi�!َ��נs�5��&W ��.�t۬�Z�P�:ڷ�����\!A�y,_Tw�L�>����H��w)4V�iݨ(mD;f_(qep�j����
�#f�]N��f����mi�����
��h=����^GBwrv��&:"g*o������W���Y�j��\=H\�E.�Yv��H���Ӱ��%צ�PL����'\�O���&�/ᣬ�r��)n���sJ���F�Uҙا;��><8��z��񎃕�0��02bM����Z��v�)�L�4%��:�k��5�r�J^��L�a�Ⱥ���[]з������ޕ�|K��;HhU��+��1�Ij�����vg|c5�ub�G!;p��EQS��U ��e}�.è1�U$�
ޫUb7u� �ﴜ��jI���:oN�ׇ%+uC|q$��_s�9��o4nuw�����;�}�U_t�a��ޓd;ۑ꒵*�/�*�M��'�f.zښ����r�]2���G)W-ǝ}���e���.W	�@}��^�td(+.�Nޣ2M��s�u`�|Gw�o6D��u1�6I&�JXku�\(wM�r(�tGP*$�C�s�%Đ���73ĵ2�\,�9b�^�{ �D�=���Gw0���s��w�)��EW�$��ȜJ���r�0���9������N�;J�Y�);���y;�j��;(Ot�II,�nx�+��9�Ii�/:ݫ���u$�Gws��ˮ���������4���t+��"tGtwnN{��Osݨa̬�Z��h��]�y..���u�t�/%�p�u�C�:��jZ����y�������=��j��7w<E�r=D��"'*Y�".�뙻��SZ�����'��OP�winK�9�z��N:��):�ȋ�r*����tJ�-	C�˲���[�gI4WWS(��.�$�2�l�ww�9Ԑ� �rs
��=��p�.������a����Jd�^�t�Gv��R��Iwww(4�&��N��^���GƉ? h� �7��o���U����U�عR�Э������c�l�v����̡��+��̎f\�8�������0��6 �0��鞡@m�y8����Р"3�-ċ�u3�*��o)l�׽�˰�
QhC.�x�J�,F�h�V�B��X/���5�m������ؓ}]q����7�(�)��豋���χ��J�&���@;���e�(�)T������+�rW����x��4�xRD]7n����)aVt�~�%���r�0(���\M�/=3y��Y�u�4TNM�$�%r����4��B��*@�uS�[�,�~���Li���䀜یXw�Ǌ�`CFN	�6G#�)C=1g�[��(ˁdfR.u���W�X`D�b2�x����MdiHŅ�b�� u9����<����u�׫��*�4�����z pʬ�\Er,�U��|�v��{���Õ����.�CQs�}Co�V�H�S�`u5x����|�#<��c?l/r��Y����Veotth8�=�]#�����E�9�K�5ٮU΅-�1;k��eޝc9�m��1 ���:.�R���s��w��ރ���Wml�3K�F��$7[ϏE�o���ix�$Qr�t����W�� �{�C�4��8~���mqE�3�t�B(�u
�ER,>P%����ѳ�L1�V�S���/���Y�,�Y��Җ]�O�b��@�%�dک�!�x:ۉ������Y��3וNۛ�!�ζD�e󥐴�0fץ���"\3Ú���i�}����0ϗ�ςG���q{ʔ��GɃN��c\�c�y�R���tC���b���.����	�V:|jA��j�|��)���7�&�K��D@O*&��	�=�R��2��f��#C2$�N5*^��ޥa���8{�� 5ˁt���m���6��'S##�N!K:�Ӧ�5=B��`����Fa�d8yPh��S��F�c5���{���:�tb�V�e��� ���Qq��Y�}P`�qd3Ւ��RV�jgn��u|���~����Y�],�sHE��!
s�<��t�(��A��muʕ�0�(t5q:�����FU��j����x�;˾�BPoG^�:��1j�е
��o��>\�d�V���^g��ygF�}E�1�܃0ܮ� �3�f�L�C�����깙�&5j���ܿx�{�/;�N2�#�.�
�Գ��Xy�ÍR9oê�(�.8�Q#;*r��+ݜz�+�Ju/a���{�=��V~��%��a�k({a�xoK.:��݈��T��M��F�~��r×p����&�u�K��{T��I�P#$S�����^�˙Uٚy�)����Ҙ�\�6B5涸ޮW�r�l�N�8g�/�wV�ש9ұknOeZ�^c�����Ft3o�"�PΨ͊*Fl;�xڡ#[�1�2w:�8N�UYB#
b�I��� �]6x�9�'ezu�x|��O?yc�V��g�3�g��C�V������s|'ȱ��[���Kϕ�j��N�������N�}�n�ݴ3b�DůH�	
�J�7�����G���Ga��r���0~׫י�%�P�ȍ󀈑��)A�'��"�t�a�5х����z�+ujr�������C�x*X��HV��1��Z���q��3���6��?,�p���f)Y+�[�����'{��#�y8!>��v<\����z�y��jhe|��3p"����[>&��oo�'2���V�jq�qVwN�vN��q]��Sv����������M���H�����|j�<8B�Pt;�����������Yz�wf���Bư�lGL���l(E��f'��'�����1R�0c���gi�օD��#���<`�d�R���$�K&� G�&cf�w���/o�W;��Q1B��!�^h��RT�tO���C��U�и�w��;6�]������.��{�w���/�����=�4tI�F�R��n(]�KkM<�.�T�&�QfZ�Yԃi���Z`��r5�<T[s[s�Q�B��^l��M��)g76E,�[�W���#e���m���2�ԗ�޻g�'W\4@E�z�l!�Ş�8t4��"�UiҚݥ;�	�+.���y�V����\��nI�DyʔF�6ݣ��L�)�d��nǬ�Nh�e�o��A��ѓ<Q�nQ�nTB��eP�l�~����ҘF���=�<$��W\c� :�u����N��q<��]�fQ@�Ȧk�T�E;u���sd|�p�GGaُ�-�v��,�ڧ���GoK}ڱ]�,��_b}w�d��2n�,���2����  �;isei��d�m*�g�����,����������=|R�g������n|��\o���"�C� P+��ʙ_��B�,�%Õ�2z�msz���Cw/��G��gG���Z�^��FE��̵4tY�j�,�Q���h�4`��=>��8?�^�����R��M^��[Ʌ[O� 8O���kVu!��oכYd�D*�Z4/�Ұ`˵|Z�XKF�W��J$n���5v�{mg.�Ί��P���"���X��UF����B^���M���n�)��遠����DT�T�b+a��0�E��F�4YF�D���S�;���-�RLLp)��H���8����a��`��r&�#H���c��Z�St�r(�2X,�e2ܸ��l��6:p�YPCC'K^���SNsه��fr�Z��=��CŸb�*z]D�	�5�Q�*����@id���>Gx�������6����k�Ɂ���6/���܈��#�f��Pܡ���s$�z3�fpԻw�9�U��W+���`M|��Y]�&�ϸ��+���x����^!;Ո��!���k������M����;���l無"^H@�	�_>=�@��+��%�x;�6<V����[e��!�S���6�K��'N�A�MdiH�!�b���3i��x�ͼ[�d�c��>���hW�z��g�ѭ�<n\��q��R�0�
+.Ok޼� �:+��og:�Z���B�1E�t_K�G*�[�ՙwJ%��a*�*�͝6m�Kk�+c�(�
��G��P (��X���\�75iR�ӈF��p�)d�'�i�V���1�$Z��x�P/L��g_\k�V��s���:�kI,D2��������mM��`�dH��s��%�"�>K_��{K��Z,��)�upt1��Crr��P"����Mɗ�uͅ+3��J���ltB�gm���7�\j�����N�F�d���f+���N�Z�GQ:!ҔDBzA���VЮ�aq0�?-b� �ä
���2*�ZD5�Z�7�ݯz�~��I������6�u�\����3�m��l� �㫮�QҮ\�������[�����QncܮTr��y)����]�WNb6:U�N]���}� �7�]ʌ��7P�?Y�j�H�X:P�����ާ*itKN�Ƽ���k۹9tb�W������
�^��|yp}�Q�r*7*�ӱJ����Ukw�ɳWS"��3yPP���0F�q\�/�ݲ�tT��2�g("K�ht��3g+�Y��껴!	|�k�\�D�zw#�4�u��e��}��H�ƥ�D�Xg+0,nJ(X8Q&�Yb�ІCooy.�F�;�jl�KʜdFS�pg#�Ȩ���?�YA���g.iv���d��_Q�Vn�"���\2�D�N���8E��0`����Z/.��QO��k*R��llCzYv�Jp�-l�Y-�趦�X_�/%�K`�1���y�Z�!��ݦ���t���E�YF����<X��v���w0kw�����B<�̑ƥ�@�].8���j��*g�y,(��=&�m`�:�EH.�]K�3R�{��W�{X+v��s�`N��Y�Kh*. .�h
[���3�@�\I1��k��Oi	_C�Pu⳴��9]��ͦ���j����r�9ilvoRK���� eV&��y��>�\mP�s�.ej�R6&��*�xG��+'��Ά�[u����x�S���F�q�2d��@x��Z,�yx:����PWJ���8or��5��񷛋�>~�<]�V��g�p�}�l�;j�W	>^�T'�o/����sHp�;,���Z��Z26�
D��j�0 �T��F1�����<��eJ"��t�1�ȡ�&!5B3�ԌP��#<Q��Ӭ�bO�jA4�ʈ��5!DP��a�9�f%۠M  �ifc�Z3h��ƙɧ�zQ��&+gƲtւ�K�YVI2�PPH�BF�m��qv���H!0%g��ʮ�d]@�a�lq4��)��j��V�,�x�fK�	������^L�}0ba���HBg����F�od�X'�)'nG�=y�{�����)u^E�i���MH3��#���c��bf'ϼ��si��)S�Nv������J�x:��3$/%�)��vR9��Ncɼ-ڔ�#b�괺�8vj�0让�j���p��5,�K-�Jb����sw�<7�q� �AA�N�=\�c�֪����x�'urmì\��3��3y(a
Qj���XE��YmR;a�$!����DR���m�Fr�[v#���6X#.1@�Q��ŝ�u��<=5T^��P+*;w���X/� qgX�4���%#|�N�=����aӯ��q�;�I�|�A��uhz��P%��x�~<N٦4m_.���{\|���\ҕ��*��G鞈�㈞�:D,�68�T��\��։�é���N�s���RS01^�����RwT���m����o��B�)�K��*/1��ɨ�+ë�x���a��73���e����E��TAg�AF��juv�s��F�����o���y�r��O�*̦�J�L*o_����#����~��pC�:O��"3Z1�yR��9c�-Dʑ��Xs(o�ьo�%�=-ڴ�THb���BX�d t���E8��XЪ�5�0���]���)#�\{xvQV�V�����݅���򮤶�ӡ[��\�}(��֒U�q%Ƿ��h��Q��J8hb��'7jwX�����fM���V�S�#��An^cķ�̵��˦qd�__V�רּ}�U���׽���B��PPa��S7&q�:,e.TUS��������/Sy��4T��]�'��T����{ �xZ;x��Y�<�l�{��S��YyQ�Q���V�0[��f���1K*������\t*��?���ꯏ(=�.#��)��p��g����r�Q�� �C����E�*����B ͩ��4�{e5t��6BeL��τ��x��j�?T�ѾJ_sq$e�E��Pf�t���F�4�r���=�q�G�u>��T�1=ZJّn9�<��qfЯ8���FT3bvh��N�ˈnen�����O��)�f������4v;���k��k�a�!�H���X�����;��w����L,N�q�(f�Wl�EVN��b@�x�mQ��H�b2Vwt�U��.),gU��؆lj�qc\���D���iK��_˲�)�� ����Q� �G�2v�t��v�S���g&���ۜ���$^�\��g9���b΃��xX�\$+,�U�C֢�[k��b}�7]龉m����N�rЩ�T�����%��!�4�]���'Łv�V�٬#���S9.6Xt��;��Ɣo��r�����}w708us�kJ�ņn����	pLc��m�/5R{�V5{l�A�-����j����������&�	W���K�gv<�ދ�c��Jr��g�`#�h��E�C��{��~[�-Z"�l�����͡j,��˫浰�*f|�{,���v(�i�ի���gO6�9N�[y���:p�\mՆ�M�ը﶑�i���e+Y@�)ks>�y
�'s�\�^hk�16󱽧�~ȵ��7t�,I�M�֓�m�%P��oz��h�ۢ�ep\�ʇ�%r�T6q��[q��{ܹ���q�+4��E�Fo%�}'F�,�t�Wm��j�R�ޒ����T��8��oa���f�
K3v���G�l+չL�wj[����m�&;�V!�̊�t�wu�w��-[�����1���\��ܚy���q���v��;v��K�YsX{����s)B%57�=�w�y}�{m*a8��U�+H#	�u�v�M�a~t�U���-�OÒ5��xLF�
.bUdr\4p�AguZ�]��\K<�X�R+�++	لT�K/A�Á8��t��o�	���ҝ��#�_�MWn��D��oGx(+�)*�c2bwҺ�qV����W���.��]�wnяȉ7v��Ԇ��+g#E�f�v-�e�PT._ )�\�>�<�6+��f���j�ֆ�Ui�t9�e0%�n���v)�Jc����Z�i�Y���]{�o/�X�Xc�i�9�f�.%��l�TzY�0�͹[0�)�=�5eA���*] �����w;�:���T�����5vL���p�n�2*��t5�A�p���>���Y��y؏�󫬋�(�+i ��ޚK���o��+�A�����SE<�v��r�b}O������ھWP�)��S��T�dv�Q^S�&m�G�f�^5��1���7VU���t"�X=�c�k�ޕa�"-�Vg%��\U
�}�3�Xi�� �<�v�uԻ7WM�ݢAo�l_Gw�<�Z��}�����]=�,~�j|.^��͂]���3���n89kHJpZ�<t�I����,ԗ{�&b!��a23ogM��)�5�՝��j�PC����K��[ʶ
hq]���uN��MH�Oh�)��������u��y���.�TsB�e���*{��H-�,�*�9-5��-��2unH�*�u�9㫎��Ўy�;�U$��D�*\*�2���+#�/�J�ʈ����Y�ud�����=hZ��Ju��'�ft�#J�wB�v�s���Qqqp㒎��9^���sW<"aE��;��D�A
�Ki�4#�Ep�]]=]`T��i�	NIAR�e��y��S�!W=�UȄ�{���	SMH��2N��IEsf\���L�]Zs�@�M�t��w)�h�hX��Mu�UE]��uHSd��D�$��I3��D�u���t&�&r���U�I#B��Iˤ��r���<G�����*`���v�ӷh��:;�|����y =��a�����v>���}�h
ĐΑ�K�'�U}W�zy������F�h8y��­�ӳN:_ey��
8k��^K�����K8�4�w\Κ��t/�R��.h�,���3���nRZ'���=^���}ٙ}���-+��
	Pq��#b8K�"��%��Ƭt5��������Skw���UiF8F
�D@4'dm�+�]KI�oQ�t<<eB�c'+���n���_�F�GH�
A�P46D���b���od,=7����wk�o1L#/Uq9!�'��L�Q��(�W���+&7�u]�!��ܬk��k�կ ��5��^旄0P^R���0B."�fOV^i��n�\>�Ϫ�]%��T
�����E���1~�(�4$�]�ve����v��o�d��G���HuҬ���}�]���V"5���ڵc�V"�.���pl�i-�Uf_�MU)��Kʜ/`F>�|�ʜ�8�P�Gx^ҫ����[��F�{�ү�%�;}�����{g4"v��Ɋq��0L�@V�4.�������}o�wOp/7��
�l�k����#!�C�ZW>� �
��ʧ4�u��|�%_cH��/U_9���UW�Q(%�n��K�H �c�:�,񿔫�o�elM�gN��H��f�1&���������:
43��P�,�r�Q�Y���Ul¨���/��]�w��+��U�;P�8C�����}]���H�A�lؖ�q��e �W�SV_���jv ��U�Cҙ�\�jaq�^.�l��sڤ:��l୞8:<�]���U����Mmq�*����t�	�pϩ4tka���Í\mwX��a���׻�t��Yӥ����d�i�ʹ����D&�<���4���F%�%{��+�c�]G���e=x"�>�\)_|��_�q�0��uɴ�Lٸ�؛9)E��x���7�4�,��$F�FD�R0�A
��0<�垛'��N��O_�����|)��>��tI���]A�3��|��Kf�;[�G>�XT#�QE0&z#(T����6#��3��#���`�W;!/CJa�\Oڴ�QxmN���|1��؃^݇t7��2�*y�Z��K�yU��X%o�c��kN
�3
:*^�݇y���Hb��5�����"^fܙ��\0�GñN#�=�A��e��9�mq�E��WE�*��k��!��N��YYp���G���n�+������3'57N��8��aD��?SA��b���m/b���uP�D�	OGsǳ��O�t�/�6OM׸"���6�ϕ*p� O�sD\l.��v��9���*l��Ir�H�҈�^L�S$'�rhNl�bcؠL��J�K�/-7��W/�]VpS�Z�1(5C*�TV��u����Nw,�E1���9����S:������ŅXZ�l�G�Kb����g��t��aVr�C۞;~��T�C���#�p1GDqg��ܢl��qumڄ�����8[bQ��Os���nI����f�_��ב71$��е��5$#b켍�7��.z�l��������Ôt
!d
(�º9j�����Z�!����N3�jZOa�YF�PTOY��-y���	�=:nt8��+)u���V�e8L�@�eO�
lrڦh�wL*�ɞ��x{�ҥgSBfe�R���j����PJd��vْӫ��0�֙Y���D�V7f�"��1�tr5��s;ˏ]���vr���gkNڌQ��R1*aC<����ᴍ��Y�54B,�) ��wk��s�(\�Z�P�C6z�T@�C9{n��s����2$n�q�\�̋�w�Q����4��
��a.��":5ጳ�K�x������x��F7����/�8��*�,9f�b��(]L�%r�X��T�aBĶ�=�&w�ٯ��Jx��gϤ81MK��(U3p��>��`t�QT���n��|bOoOP[8@ǥDG��@���\�u���{ �xZ=x�2��0���J�",��`ٓ�*vQ��8��
3��A�k.{16م�]���k�'7�;䥟i�uQ��Ժ��g��Q�9f�B����W��kY!vo��nj��JL7�* �x�F�F�:b�xa��w��:�.���ڟ&��=}���	zr�h^�ʬT~�d)�O���2��_P�� 1;��V�۾R�v��p���VҷoY��fC�l�u)]vab����wn���cf�xO\T�E�\�e�A���5��%�bOW��3֊Yڗl�6�K0Z�AaF��!�g8�3}��J [��f�)c���&���gfg/���Z���ޤ�~�k��]�΀򧼱Pg�d��;�٣CxO��eiZG\�i_l�Ƌ{ED��c�Qu��K��L�B����U�3�P�>&A��Q'�0N���I�ZBt��z!��,��,ٵR���Ǝ��x< td��������b��#�C��؎7�qō�L��Dy\mt��x��=K}��+�]���5H���x6t�^�eף�<\��T�5Hz�u�&�3��%�K��!׻i�uIo(�J0jq����q�
t�Y�E����k����GD�'o�V�8Ͻ�1�j]�WhngMR�0�Qߥ�b:"<X�>����p�b��@�l���,��ԥ�!K�eצx��`�t� ��R!cB�!��1�^�<yZz���K��II������!1s#��P6QD�Ң+҅P����B�5r4�GA����u\t�@�bݢ(�����0`��)F���1N�"��	ӷ�r���u�C��ޢ�37��K"�jXK]KY�c0�>L��>9��I��Ö����5�^z��%�h��`"�EN�;�m�v��o<�g�+�Xޯ�,K�9�'��^rCv�Ht�ܧ~���^vra��P���8U3qq�*xĊT���(N5���(����t���%��ꦮ���=`�C4p��뤠�Z���k=B��]O���aAwG�����$]���ݫ�|O�i��Dv�#>&��A�#Y���K5�\x�'o�FqN�=u,�DoR�������c��߹5&��N��[K���;�˄a;%�*�e�M�:ӷ"}�,��5\�-s�S�F��*A��<:�ݟ!�[�/~˥���eod}��7\��G"եI:Z��j�>��Kf�OD_C6ۤY���Q�AѼ�Y$�U�T��K:\�'<p\�B�H�BW����qc��gbm��񌶭�2�;K��`dD��\�@�9�2�6�Q�b�˚|$����t���I�k�\m�=/	\k��1 ߕw���pBt��eo_�,V*g�����M/nܼ��1^�w�cv}�uN�Cu�R�TK"��u[r�wxe�,��yO{3Vx�oo(g����%�y'n�q��l��r���W�������QwĻĲ����o�;�������1X��2,ۥ̜wu�/�,�x��N�;�M�hvl}$��5+�to�������:�����w �'���d4)Z�իT|�p���5�W"qБS�;��8��N�t���F�Be�8d��T����DWn6��u�H�vMO��}�4�\�e�Ԉ�vY���dtJ2`�|x[����:-�S��{��>�C��1��XN��	j֋����%��B�,Jy��i=s�n8���E�_.����b�U�-�;5<�c$�B&�K���]�䷡Dp��n�3������|,�,)*p�'���qb�n��JnTmaf�)�.vd���#�Kɛ���E���gQ����km�o<핾��֘��ew��u�.�iȲ�o)�W ܽ�`ޚ�Oz�
����s|�2��U�D��P"��@�l�p��.T��76E���FҴ��6y��w�:����yO�����T5�j�&�3��Ś���������@�6��SY׸����Je,��u�����k���t�i�$��Q=����uXj�Bf�WK�՛bR핻���Vv��ؒ����G�Q�x��Ρ�a��<q� _Mt��X�,�;nR1�:�����
}�����2e�T�y�ޛp���gTI��<Y�r�[����ʨX���	�+�4{����u�3QT��L%�q���"t�Y�����[�nҫ���gG�
����i�
�X�88��r��>�C���wV���JS�qb!8�UHܩ��<k��^��]�+��(��	u������	v����$ҡ� .��lc�d���^Z��?��J����',�\�3���Ѿ�Y�|x�:�k�����S�lnZ�.���/���r\���l�.]q�5��XJR���0��(�t���"A�g)6�1���>��X���"+��`�t�+����!2�B+a�x�*Dhؗ[[S�ر7)T�h��@`�3���P(�/�ʓ椙kMW�x_mzH�,�
���`հ�pB%�9:�n�v�[��q���+4�n�����.�x
x�-��2�6���u�8[�GP�(�{����o��<6�8��u'�Z58u<�"��o��\�Z��]{u�YJ)�,MK�Dp��gL�q���ܧ+�^v�=U<'�	<6	O��)È�ёf^��;�"�^��̀zl%?.�e��;�w�s�t�F�)֥�3��)��^e���E�"�GG=�8`�YNs�"��� ��5t�;!p�P�:#3U��w{��B7X��\f�."�=���K�u�^ p��$o��"�R���7F@o�i�ΐ��^Mw�?@��g�,L?�ih�j��ӝ�=��uI|���5>ne!ʌv�Xw����1�u���B�t$�q;
�%��k�Pc՝|LO��x�`u�Ϲ�9�Q��ǃa��\9��Xt@q�,����-��,��u2+ٳƒ�TU��&3�l�-�A��bPt ��`?z�Բ���T��=�ȕ5�nv��Y=���!/g.5F^�q���ȰeF����4rܑ���4�F��������H�k��Y�5V+)�o�ay��MB�_m����s~Wm<&��$����_S�2������̹SiU��k��Ѥd^T��/��H79<��0�j�M�n�v�T�G�>���Iɮ�:��ȴ&Y�`>��07�F������b|��Hp޼~�7�s��|p�;�	9���+����P]ԝw����ϑ��ι'��g��3<7�8.�K#���pĉ��a�%x�	Bh1uA`=)�%�X�R�E�^8��^Nd��a�
�]CB<�H"��2�7v�='N/gU��G!��7荸Ɏ1*Q�3c"J� ��k�fA�p��N��s���f�+���̈�u�d���E�tv�!20�*C%Dts���J���*�U��������D/�}),3��u��1�ɹ�˺z���^�h08��D�P���������\AU
��R�����D�Ek�s|���'9�XY��,�����w=
����g�a�"�n)�Y�*�%��u�3������+i�zG�e۔]8B^�o������N*�۳3��f��x���p��FN�w9��]gD�	�D+�,��!�
�5`�F�Ф֛���k�I�C�+�iS[v;3�t�ND���pi7[�{��r ࿚|F8�� ˻��j%��˫d=ʳ���P�Y�EtiS�)@f��--2g$2��
MԈ�Պ��)(RU-�#71Z�(oK�I�&����&V 4�;��5�-�� @���5��Z�Lv�g�o6p�J�|ʷ���9�����,�[s�Z�.�b��s���B���L�wf�3�E�����î�%m�*�$�Y���%��K�f�����n���# ���&�}��M�#��s����Cb��ڡK:��u�l�Yvi�[�^N������X��\�!U�n��k�V@q�yoa
R�wAevFXھa�Z��DZ�K2�i��s��t!6��]<���Nn�N9�붑�'y��rr��\2
���gJб�Xn��hm[�7A����QZEB{��]�EV�N�D��=v�wڝ�WK��P�ww�ᝌ���M��(vm�-<�}���e���S��bqN�W��ڔ5;u����\B��`o*��%N�UgpN�S{�`^�z�B8f(�}Y�cf���&��i���\�f�f�mv<�~S��i^��hd�hU�2&�+�׷�E +)e�u�1^��Ȩ3�U���l��$e��VK�9�^���I,\;b�y�)�	ȱ���QVN7V(�*B�H`V�C
�/!�E+�C�nְ�0�Hj����M�S}�*����r��
Rw6b�mSå2-Q4��a5w�%0M�̲8�5�f��Yʑ%�`M�a���Xn^�6]J����.���!t{����ꣳ�u�����HUz�u�|�(�7��ҙ����#��[J��Whҍɔ��n)s`8��.�ue��\+�b&3Lw4N{Ab��Z����J�R���sikJ�����{�gc��ftò��n<�B��d&�rڔ.VA���M�#���1b�3�4bW���ȲVnV�ݞ�H��\��bCzЄ�8b����{G�uo�c����|�u�%Ov����D��
�yWZ��C�7����xS�ʭ�Ѭ���]KT*P1v)9�k7w�,>�4"��N��[ݩ+r�sjU�$��il�:N��������A{R��n�0�n�k�
�*$������Bz�=d�;~�����|�����X��ڔi]�2�97P�Yhҋ@JΙ˃��u���ք�Z!�j�AjV�vbD&��I
�vY�IR�L�"���BU*B�̪��΀�)��ATk8Z�iY��մ̙$�)*+J�dFKY��Fr2NҶ�I:pN*%Dt�CQ%����,�Q�Z!�$Y2��AF��YSU��*Ȫ�+9I�Jò�R��QJ��ēB4�J�R�2ʚI�B%9V`S"Qg+6gN(��J�����sD�26�D(�&���$�J-:TkTJ����I#4�:Z�ɋ(�:r9��؊��9��I�!�j�
$�bId4�W)i�ًmD-�+:5��2eˠ�nL@ޘh���-p^�:�k8�v���՝���k.������jL��*75�kI.1|��'Vf�:qy:R��e!I�`�c��#�S06���"�C6��g��i��,,/o1d.jn�l�R����s���t̑��O�<�3�@����{�3o[}�7y��U�qG��$dEy��7�BP5x�2�6�5�<U��`��ǡ9���ϲ�X�
�Hځ�ح�&���Э�J9T3cV�Q���n��,j�#�R[	T����V�lz�EG¸T�mVK[����A��.�\5q!��σӃ�ٖ].X=*�
�s�kp/�E�&2&8��Ǿ���.�e#����vÔF�;L�Ǳ�ȱ�5(|m�,s�92��i�Χ�z��g�Y�0z%��j��gE��ٹ�nA"S99*�j�K�[���DP��t��0Ģ�B��4B�@ˌ�ւ��*�^�Nm�^J�M��u��zD;�D=$%."�]0�b)�0B�v���8X� ��瀕�oˁ�k�sϲ�F������Y�ͮ�2
��"꺚�f��gW^��`���+T/�rB��W-�pK�K��sy۽���+�5s��|�����V�,g�as�$D�-9*{3�6"Sȩ4
'6Y�屗7i��3$UD�e��@߳%np�
]Dӑe�e,�ƨZn�vO1I�IYˉ���wF�6��Ȩ���Fl�qk�K�!�-�E�����:�앑M�h�)$G��K��5^)�o�"�3��Ś�ܥ�+:���&�>b�ۄ~x�dڻå�w:hע8�^�'�[�GW�R0����˹�������G6��8r�p�
��g@�4p\�k����܅���ZN�ҭ̈�$�~�.����:{*Z��K�O)T��@GhC��Պ�����L�bT��e"��VG`��3y:E�G�����;�F��^DK����r��	�0�/b��3
)�=�\m�Ǖ3�����4՞�Ls���O����B	�"�hq�{n�ϰ�K>?(|(dB*��Y�[�m��4�Υf�g2�l4�;;���T��
&v$�w���b�wB�zi*R�V�T�jâ����wP�Դ}�a��gZ���A�/E?�T����}��Zus�ǩ=̓o!���8�s���sgp�WS�8#����:��]tF�P5����ZU�8�#�ӣ���"@�3�ןJq"��0h	b��(.�3��1`��TK�8�x���+Eh����!=�MK���R1�jZ07^�l��r(����/�{(�(�0o��>��I�eI�jA�֛"�"\m��v���[�
Ńԏ�|�3^Kg��O��/�Q��8�hȳ5�b��<�N�e��\�:�pCcg�S7��˪dP�@�p��ҧ��I�'��toVn����7�<V
C��r ��)��z!9e�}N����Y��R;h>�Q7�w�/m�S�2a�1f��s���#6�"���k,q(XA���2����Y�oef<�u�
�u9�[�������eC6'f��oc]<�ƓSV�e�x��|<K��s냹_����hwg;fSٕ�"��ϊyꘛ��;�H��n��X:�$4�����$�R<�/FiA�[��$�TT������w����A���-��*��՚$��3~���7#q��'Z�Eۥ^[GH���-N|R���*�,�X��%��B�F��5�Q��`�X��[����[2?$&j��
4�@�#A�|�T��ձuŸ�rʽ�B͞+6x�	h��⓷�6�'�W��D x�:I��0K?Y��y���^r��C�e���r]һb܍(�����,��aO�2��^��F�273��f��*R�P�bʨ،4���_L���с@>���3����lÎ4�9�/%\C�|)����X87�aP���h]i�]It $*���(�s*�Z���s�6|�pM\"σ�>��`�J�P0���(�BzQ��y+{N��p�\��po�PR�n�3ѳT�9��d:�\BU����q��^�����ҷk�#0ڱKɂ��3�"6�,�1AJ"^�3yP� ���Ԃ��9 �&�}Ј�,��3�_L8��a��x:҂��ǆlO�ߛ5uhM��]j��J������N�c��.:��73�_n��}r-X>ZK����ĽK�Q�3�Tt����Lr|R��gX
_k���J��U��ۛ)��4oA�Z�55_A"���]v��;��S[�R��D��|�SBqʈ���E����C�Rω���b6��+O�ﻹ�J���N.p�M]r�;smΗ�8؃��TF�pDW`m�e孄�Ў�7%S���,�����a;%]*�6D�(�{q�nvj]�*�@�n�6X#&� t�t���eӔ]�#%��R�b
P�U���Ve����$���X"��H@	�I��N)~޾�s�Γx�G�⨱q�(&ݳ9R�
���,�8�H�ҸРC���t����%يv��K�@R޶mG��Hȇ�,�(�<r!v�R8CB2�}{�ɭP�Y����4��n��r��
�ْd<^��!<	Q��9t�uG7��]B$l��x���#�'pz��0����2~�`���܈d"7ؽ"6����%c]��%��)�ɇV�+��MX<&��.X=�_RYς��gr��`�i���Ib�Yw���\t�T�'��i�tL�������ʐ�����v���3�c�Vb^�'b���u�.�*����G�ͽ��d��ٹ�#����S��v�jG��i��{;t=Ρk���RuI;{�Ι�A�j�+]Nc�0�>g�.�t���l�����;���0X��}J�=0t�feJ1���#n��%��j��Nևu˃��F�Wz��ӪS�X�.�g���@�B`��4�^���i1]*�\6��%;U�)�v
g�n�Y$���#؄������L���|�X:|�8x'��2��Խ��<����a�&�����%O�d��9h���^L�S%<�����{���Yׇ|��
ՏR5^�I�\dɣ��d��>�.�9�p(�����U]Jޮjaf��ˢ���%����,�ު:��V�S(@p�͎.9V^R��TX}�Q��z�c3+v+�:Ԓ4_O`L�Ek8�ԠEx�b|F(�R��'pD��=Է�e-�;��.�E��æ�bt׳��<Y�#Oo�
�V�ec�9��t𜳮i>F���4�j���Jp�����+��c=3ś����W��om�ù@7U�>rA�h$�!��;�tt��Y�eL|�[�9҈��{;|��T�/k'�jD��d��A�*R� �*����7��u��6�T�Ֆo)���Mw`'B�"
q�w7��]3o���s��nC�3����'p�m[���{�d�"0�#j�F�TB:G�<�����w�)�mƂ����T�8E��F�����N�^�b��"�V�u�(�{E�V�\r����O�NI�[��\n\ۆr���C;���#')���&�uk<���E��<b��
3�AHh�	'�J�Z�'��}z���xn�3e����}з�b�V���̋���< �:�k�p�o��J�[5~����o6�2�)�Ɇ��T���X3��n$]u3��*Y�#K��0D(�3�-CD��Q>���6h����V]N���~�U�]��i.㴬)X�UC+u�;�Z�(�@����Q��$�A+!��$��Ra�tr�[���r�b�D�q����JE�3�B��:�p!W��O`�/\�/�N��(I���%��!��7�I�ʺ�)�]A�<}R�A�G;��a�<�S�Ti/W7��0ճ�t�aw^U�/����S+�;���}r�A���o���hᬤ�tQ�[%oc�ם'1�4S͗5`6e����M�*j�syro��R%�7&�|�52>���rtg����_��(<萫ݏ@%����S�^�]AC+6�.�cN��p�0%C�4�S�,�H����.���"�t��2plio}��ٷ[���ʕЁx��5���>�V2��+:CڞOzŃ�11����i��U��V��`F�mB*�Yq�r,���Z�Zz�;���k��2�o�{��y��h�[-��^�.!��6�����g����l��r�g'�,@��CƲ����\�ۚ�؎8��V9g�e���gf�Zķ�����y�`�u�ǨJ}x G]G�厶鬞\7$��&ܾ҄ekՋ�X�yZC�nz�D�����ߩhg��2�.�:�fE<Ec��A�ƝB,UN�e�4�Er�"��M0k>�^%{�/�>'��	�r)2��7�����u��p��0LYu3�C٤"z��BBh/r�Ƚ;���J����^S%Z��;M%)���|�Eu��h4�lb wK��k��A�-b����FmaRl2��)������/<4t�wwc����Ŗ�ަ#(��c7�kt=�N�ƯOk�V$��G�oN��t+��D��gYD__T�ȇ����!<H+�Z~è:�À*��.T�L�V���P�L`0�&�B'M�Ƽ��O
uf�@	{Ȃ��u�\�;��L��<f+ʃ"D,�,؎��+�tOޞ�����;,����ۭ�J@�3LD�؉�e� ��+���X:RP[�P*���J��=�m%��ܭ��^F�>s�hM�ʡ4�,;�,��VG�j>uWl ���3·���^z���Ʃ[��6Y&C�.�M
t�r�U<jey�6g��2��Y���P#�FR��-�Y�oK.�;%�*�{/bx`U�s�m�S�ȼ�S��h8D�uLؘ�%�2E:@�7��f�������$4W��w��_��E�:9�_���N`puڝџ#���_/�x��פ��^8�Ob�����P�&��kT��%�Ԣ�lhIR2�Q�ʄ�Nx�����H�����,�0%�K�*��ͪ&��י�'˧%´���w�4b�R�¯�i�����!�@�..��;�Hw�Ў�~����y;��ج����ٗ�éK7�9��ڛ�'J6�vsf���j�Y�]��3/�pޏ��`�o��t��3AǺ}�#">�P��\�,�����T��u&��J=Ś(��g����ZХ��+�s<&$��*��B�LD�9�L��n���N>�. �x~*����j��R[�A����V��#��3vwj�R�n� �|%DS[��|yxE��+8�X���+!�٩u�N�KqV��"Hv��5�ታ�d���������=�T�H���֓�b4�c���bg�g��Ơ��Ii6ڬ%;Z.����v�8Ȭ�oT��T� ��^K��fb����%��p�!X��B���T�L&�l�x���(�JC��;~�&xE8$F1"C��R�@�b��Y��:S	O,��^+��R��E��0�8uJ�ds$SU���wKɛj`�1�W/�e��+^�α(���t����r*�Q̉:fJ*���.�h"�;��~o�ߟA��F�P��+T�r��mf�Ri���W.�RT�&�m>]���(�W8�١d�;��b���#��;�\V�&��Q57.���6DM���~ܭ�2`7M��cv�L�9Na(f;.8�a%����Պ<��T��,��Wy�O�X��X��J�<ٕsP�ᎏu�m�Sӌ����-̧}�5���Q�ݮ��wT�Q�g*��U����q�Pc���]#]#ĥ�z�����s7����y�da�V	�Uw'P�X�
sI���4!�3Y}ֱ�u��uE�s:���ݭ��Ȝ���ʊ7y�]�wA��6j@V΋��	o�{�X�1�-��7�;W}ғ�U�k+�Y�9����kEN[�mJX^u-Fl�x�&�h�2u�H"u���Űb���ۛ5�n���OB��ȹӋ���/;"#��S忶��k�^�Ώj@Y�go4�m�5�β�n��8�ux�as�] �[s��:�Җf'p�Pt�k��^>s�ʅp�i�T�����D�oI@H�u�syȣ�$@��K�qBp[,c޽�х�{���ä�[�a�6��f��ZGol�{����P�K��$w/��#o��ev9�u��Z�uk6bVé�K�ۏ����^�{R�n�3&c�J=�K�x`��
�A��$f'<.�Z3`ډ�)��^U"гb-$l8.9�WJ��Y@ �$S�ofM=��Vj�K5�)n��/,dvq��e����[k!^��b�
Lm�`����2�^լ[Dmf1бv�IG;.�%��J� ��{1|�J��7Nc�Uud�-Ҹ��B��T1̬�T��˹o�CIX����7wg钑�WL���[�S��X(��6�"���4��P#��Y@��˸��sum�F�_c{)En�r�)�,�⫬�ĸ�R:�a͹�Pa��H��3qhՏm:7�B{�:5��6�AW�Ƚ(^��&%���9\&ռ�5�f�C���˃�ۖp��rR��5�OUpxg`q���ZX50�6�"��F6h�*���Y*�_�;Y�쮭C]��u��7i���|Y:kf*n��nm����qy6�����qN��>:m^h�ݼt�'5�:���FjR���Q�#��yv 3lK�S�@n�2't�n�خ�I���*7�m�]�^<M�&k-�=�Z�AK�>�6ᾔ�g���܅8�Ӣ�p��|y�޿���6<.��9̀�Q�i	�Յ�E���5m$ȲQa�Y���1��UGN&AEˊhJFZ�ҋ�gJK#��(k(Ŵ��$R��UH���SU�aQ��.	�hVd�d��t�9BgJ����\-F�ؓ&�k4�J�2�TɑP���&��LV�e�A�
HeTVBe��u�N�N&E�")9v���#�jUa$Qj��i@h]P�A�i�eRa��*(�2*��$��U�5H�ġ ګH�IET���	�BK%	-:l�,�Y$��Z[�_=����	Y�^�������r�.�|�`f�]-sh/�����'#�2�;�&�l!������K&R޵In�Z���J���k	�A�V�Q^�"j$�Er������ag����xN��yܓmwA]&�(��جW��&�x�8j��j�$\&b����L�SjmWkۖ'��j�q1S���m�4�Pɿt�0Ou,�0����Դ=���P���E)��1�*t���nѱ�Zs�� 9��&�SGK�	���U�KZu6�,z����k��O��뢃%�0o���
u�n���W��T�r�RQq����\B0���"���dv�5eR'�ڳ���[�yb�1{zC�L5�	G�b#��DoE���6���k�{ҎSW����q�p�ud"�m� �X��$;f* :�chq�6�#%�˳dm����qbk7G���=�Tx�� 8:�8I�D���Ðrfd�с�Z��i�	��ء*F�C�ne�^��E��3���l�S<`�Z�"�0T�猉x�uÐ�ړ�5���쫜ø�����K�i�]w�}B�����Sb)�'�34��R��Y|�[���/�f=�{t��x_��1�]�#���Ï]:��R�u�\�c����ĉ�<�)ː��å��F�q�!	��@�@Pa�q��9Ҧ��[uk/5��0�*-xp�M r�]C��
[�rbd=����M��ɽ`�x͆�g�;6e�ʀ��UB60Jӣ��/.T��y<�\��/-�"̰�K.�������	�ʨ߅:Ժ���q��4�r6��������TI���4Q�� �G�`Ϛ��b#NV�8j�
��O7;A�Mg57*xX6E���֢�Lٮs�,-�Fm�*�R�a�ؖ=�<�kgN��'
�/�4'�8yB�D6;�����A�N,�����S�~��%V�h7X�v~��4ƭK+a��zE����[lߊ��Etd�n-���n�;�{\�F?m
�@�4�b��'M�J�E�iB4t�涸��9p�3�H�U�����}��T#�k����l�b]P�z�#��q�Q|@Ȑ�5q魊U�v<�P�����fH垘0��t�kF�2�{����W���/k��*��+W�;�p>�A#�MX7vr�t\��I�Q���eCV�M:�k-wJ˓v�݁Y2-F<�Y:�nTݑ%9qk��JQ�b�mۦ^�-Pf�0�I5�Ttǧ�m��㗬��Oa�¦�cH�Om� \e9�F�ؽ,��-�-`\)����+����^{s}�s��gC�r'����J���qF��o�����5�U.�:�����3eN�4G�p��g��%P��Ju҈�a@-6�j�����J��i>�AXLB�C2�.%��E\<]<,IV�xu��,f	KcKaڴ��K��b���X��[!\�GMS����U�~d"�y\4<(��s;_t (�a�<f)PdH����Z!9�kAO�
u�߃����Va�N�P�ƭⳌ�.Aq=�`�E�H\e��L ���^R�:]�YR�AqROx�񽏻�Ŧ����m*��,�t�j��:在��`���^C��3i�ˡ�yM-��[8j�D�J,dYD�qe׹M
P�͆�Kʐ�\���H<u�2e�^&�����w��������z��sjW@cD��J�4͖�P:�Y5l���IlY.�-������Y�F>]\Pz�غg#C0��uQ��Cy[�<���X�#=�&�{���Y�l��2����4.����Qf�oS.0M��Q�
U�6��L��R)⺹��tt�]���%�8r�!��M�S0`�@��t��~ޗ[��p��r��ҙ�p�i��Aꭘ�r7��g<�kX��$T }!3#j��!��z�`C����F�m�� �i�.���(����~����H�蛾�j;!�$�;��l26�l���(�V͇XMY>�^^t��>Z/@����c�[/|���s�Ruş�����<V�T}Q���3:p�\�Ui �����9�M8@7��(m\,�G�S���PWO��pE����u���Q�ɔro�Y��V<�M��0zD���	ݬ��Y�������GK�2���z���ԯ�#�`��b��c��)B�TQ�#Q�%>�?	��/�M{4ɘ�w�y8e"<R�f�	�����3�W�A��-&Ѭ&;Z8��4*�g�:v�,��7�[��7�:��D@K#��M��x��Y��$=�ӌ�՜��N�S�xm���.�����4�裲Ft����9�}��^WTV�sK�i�t�e����b�X�!���5�r��)I~�3�ׇ8`�FY��)�(O��q�x��,v����R���`��C����0�D�c�.1AtÉ�����VfV���5K=R����9�[�<�8kC���ؘb��((%kUDC�0��gm��}N�y$����/��!;��?^��1��A�\:yX���V{�X)�<���{-\"0�˹W�n����2�ce�&�P�Bx�W�G�^��
�����W=����Έ;�A^�]eƩ���}^��5Z�5��q;J*b�q>����D�Pî,�k�6ܣO�Wxt�hN�Κ4"8�U�Er��y���rHy�o���4�h�C�7�Y��e�ZETe,0�"W7ڜr�U�W�0�dS����*Ͻ�4t!\xO��$k�ӝ/���bW^��f�!��<DfF�2��(�]��K�i���l}�����͙�
Rh��go*)W$�A�&l=�.�q�&-�xwX�#�]:�ӥt��:��8r��L���i*�*�q�Y�lk|)_j�,�V\=\�l��k���� U��wC8��Q�|s���[��Z�U�Na��79�Yχvb�z�qN�k��(Q% p��n���S���E�725w��v�o7�%U��4):�8�n�,�!$�<v�T@uGhu2zp���p�w����qY��ބ7T��s��Q�<{�ʬȞ�`�O�K	k�p�K��ՙ'����d[�p2"�()ćJ��^�*��X:_(���uʫM�%�bzz`p�r��P��Wr�_˩�0k�-�\AmK�©D�on�{���,Bn	�:a����E�k�M4VBa�I�:��MLR��r�z��W^�*L=�b��%z|5����Q�Rf�/��xA��J���LX:bw0`��؊�fE���$5�46x�&o"���e�e�����E<���{���*/"��e8�4�iŔlߚU&2,h�-l��Di�(����7S�]^>Y��\���5�-��yŸջH͹E�z
b���?>8ǹ;O9m�Ann�q,���wû���+
�9�֚QG��2�%
��g��fV���e�O[[�v��XD`�wV	���-����Y�>Y3����3���l����i�d�guwgl�r���`�]W����,tq����gJF7�9�v)q���׮��_^:ލ�~�6�<��a��<PO�po��#��S5�B��,��y�9���Ԁ�r��͆#�_��;�D:31�-Ӣ�\B6']3n�J4�H'������XC�Kfp��	�%O0J ��)q#nz�#��q����Ʊ��qWi�6t�y��Җ]�tO����u	AQ��Q0p���Bj׽���F��.����*�nuPz��C4��x)M3ס�b4�J9&�����s���v
C�x*·H��<f�5��сA�M�Y�P����{��֩���]�ȓ�3�xcЂ�`���<K�-<(С=ۢy`����j�@,.�V9�Ut���oƲ�̂����#0Z��J�RK�i��8 a����+Ќw]>���|�W���YVk��"+�u��Ы���:�{OfgJ�ͼ����+�0 ��m�3]�.����w�|c�IѴ�DgTȌ�'W�r�@��������/�� ;x#恨��9S��t{�zs�������G��B��x_]h��@�,�QU��0~�]�����j�'w����/v�bY�7.T��d��G���$G�,Ȇ����3C#!eAf�V��ی��1JQ�r1i'��]tm����\H�&���J�,�>�0d8�����BW�	8���~�D�f�����/T�sLF!s�<��t�((H�<*;"�U������z������|��c�G賗R$nK(=�,������Z��s��NW>�[6�T�sN2�a��.�
��
��6.�5�;�������
���Ӧwx��^�r=eGdJ�p�N7�L��~�@�������j�X�S�u`��5=�Q�i�4�2�V��pʩ�Q8it���"����5g���!'>��Xi5�C�JÌ��btף��T��.�u�\��֋ &t����*㖛�Ļ|����"Ns�=�J;ڤ:{�mċ�����n�P��&�p+=��{�9�;Ԗ�9���Ml>����p�\��Ā�5�
��c����O�4����qɧ���8��"^�f��������\$���X�@���$\�Ͻ�[[����3��m6:7�.܃��y�!7z��]����'cM�1Y�jXu5A]z�	�xo�J^ٚ����xҹX���V���@����#�%|e�n���l,xFu���c�z�"���N��@�$L�\dX��)ȒZc���ŭ�y�����p��ȣS���k1o�7B"�3,���W4��u�P`����F������`%��7�2R�/ObZ�L�p�Č�1R�0g҄�^�D'0++^�M������:���Ou�9�0�j�D=b�x�bWL8��h�TI���׋��>�6�(e]iS��*R�{�h٢�
	K�2D8h������燦�=��\��j ������1��Q���eY�l��qa���m��	Eın�U¨��{D�i�]QZ�O�e�p�����
	Qoy�����-h��{ǆ���z+��#�ݐ=�V}{.��U�,�횥aƢ{���lX�S�I�'�f���#��/�SJ�u��w�^�'�w�D�lW��[��'�k�� � KDǙ\Jy��O]���p���][��3C7��ܣY�$���;���z�s����s���*W C��1@\p���G��:�hk�cff��hJ5�颎���Uv��u]�$���Q�z!jIY-�)�������H�+`ZyY�[�؏+�B4�飂��<h[�m]�,�����1])<���)m�<���{h�S�����`�AP�>EPڷpf߃�>��狄��m���	�V�x�y=�#z���h��!�e�{����D�
י�^��,�=rx�;��y����6�"ε4h�16����)�z��@��t��J���&_-��wJ8ޢ�Κ���F��3�h�k���< �R�].TD�Ǎ�D����I�Y��O��j���XK�ʥ̰hsU$_��e��cbG�ӭ֣j@�3��*T���,FY$�^Q�'҅FF�
KG�����{o;϶�����z��֖�r��e#@�e�g��9(��ˈ��}.��_]�-���֯�����
��sl������+u��ñM����),��z.���ھ�B�ut©��ЮR<�z\t�hQ�"�8�O����Y7:a&�S���{�Ի�J��].鷵*�|YMNQ�N�����pN�Yw���1M����{�;�6K�E�X�^�<.����Y.T+���o�+5�0�S�`�n,$�����y�{8p)s�J샫r�ӜbHv��%4Uܮõ4<�ݖ�yQe���$7������H��Ao�v��!�sRW���ө::z�o�n�f�0������)� �
�b�=���c�ܼe�,�&g�(Ya���˥���|/9�+5#}y!֕_X��N���1-�Z�yr�4Y_�Y{5;�1��EF��NT[Y����dW�Ρ����rD��\6�G��;�:�{��z�5��j�dn���Հ��ث]b�l�G�8�RS�pq���x���֬����%�y�����}7�Ǳ�U��άX�g���R�\�b][�%u����(+X\�=�B@0u1c8s�@���wg[��T�����}��
#��ui�.��I�֗|�M!�5R�*�\6���P����wժ�V�B���V�ur^ۧ�����u�v[��,+"�gk���pd�-!xr�)������Pl�I�qD͌��tJ�U���fTՅqм����x��������k����d�����yN�e)�&��BiiI0wM�3A�e����u�Ԛ�7�jY��5�[yF���֋[���I�����J�Ռʐ�X7a<E[[$��ʖE?p�9��Ң�F�m�N���uh�D��R�M��:B�b�{���3J��oʇh��kbi2N] !ZaL�˲3u����o.����)�B1�Ȩ�F.+��Ӛ�vY�]��Y[+��R�\�
Ŷ��yzzoÇ�,���hQw
�-��k2����,<�� 46��� i�Z�v��u�GD�g�hr$j#�g#��8$+��sH�w�{	!,�O�.�	I����m���5m���oJ��^�.�/W�j]��(�Y�kTq`}�F{����u���{�r��[8:S&�3m���.������nD�h��HN�;1[b�S9�v����]�/�{Ҥ�b�Ȱ�!	2U)+	,�M��%D��j��C����EIXrKK)�S�S&��"�RHC���QđB3��V¢L�dt�&�APQTJ��8�hEb�BvQDv���:��K�'-C��t�$�\.U�ETΒDE*Ӕ�Vr��v��q8Phē��	�����ed��(��0���r�$�f�$�Si���EQ�ԄÂ���B�6��X%�(��Zr�(����Qb��38�*(� UM	1P�J�-T)4T�4J0�H�8Y��ȸJ=#��H$���i�^Vƈ۹���ewD�Qq�4�HFW=YV��!y[rQIv_&����9����ԝG{5L��̀+4�WK k�A��~6o�N�F�FT#f̞@�e�]�����2�2���4dY�}Pa��!����3y���dlu�_,��ٙ�z+|��z̳�A�W2��,�e�A��o�A[I��,[6�8�Lo����՝6�J�^�����M�����8՝H����.��PGjZ<�������S�X�%���=]A��4F��_�ب^�N(,��atb���HD�t�sU�~�u��|6��xз,���\E��ER�+�Y:-�k�*.��^K�FQg���u��A�2Lb���}.!��f��,ىXYYК�Wv��4��,=�45O����U
�@؈�6��lGmC{���fĊwjs��W��W�� ],��\b�@�7Q&�8�VnV�ìy��]�Q�!WX��o��5�:���d3m�\vyD�����'K��.�-�G�܎��$)��/�M�:j�v�zL��y&��-�Nݩ��p�v�P�%L-i��Eeu�Ĝ?<��=2�� S!;��[��L���I@K�q��w��)
t�y�" ��
�����e�s�9���p���*TZ{җj���g#�Rv�B��+Q0@��#�����*�K�|�5�U�_��¼i{���0�q&0��*�b��5���*���{4�c�Ѿ�[ٺ�{�ZK��X��d6&�hOD3=p����j�c!�fK8a��͕�����C��.~,�I�OO�*P��{!d�8��^Nd�Vk�В��z=�s�ďC�0b`h(��q�f(A�VLY�i/J�~[]+a򫢲l�֭(�]V��%-D�b`�E�rFY�t<tW�K�^�H���$�gG(j��QU�fF�>\�D�N�E�g*-�-�Oo/t�y�dp�s:p�9u"F䢅�'
$�{8]��*�y���ƬE��v��n�u!-��l���}qԋ0t%�lj�\]{�^[:!7i/oI�5ai�<=�~ٛNt�`��ڦ`�yN�:w��ey�O|-�6�}�۶p�M��V�9��+T'?m]�@��B���'��s�b��@,Wz�ܵ�.��0d{�Whډ����;�v�֐�+����S��S��Mά�3��O(G��T��m�Y�}�]ҝ�"߶v"�3oU2�5,�3a��2�x�j��Nx�n��g�K;_:��ҟ�d�4'�Тt׮8����+f�9�`a>����k�8ѽ��g)�j�����FO7�"Ǝ�X�}l8�օ/��*�kwu�3��iJy��~]�؞-L<�'�����Â}K�(�tsn����79������Z"ù��Qj:[��'W�^
j��+L>��%8a�R+�>�&��#=�`�(�/W�����HW9��t��3�$���N�e]�y�xx�r��z�Z��Q����e��L�F�FtWR1Aӳq�t)�t�����{N+�������V�5�f%9�k&���e���Y�"P�rQ���ok�U��")��(T�"�D��U�(E��$Hj\���=��]��/\��F�MM���$�e��,w%�-[;6A8�/l�y���$sA��9v�Z�ҫ�{0z�.��`}��u+"�:�;]���1��*�4��O�:��-X嬔�&�h�|A\���5'V��r�|����0�bt���\hߩ��b}B\@�$Q��Q||K�vv��y�u��k�}~�$���+�K^H�����Ҽ��êzָ��_Um��p(���Y�P9O��-�UQ�T�NY`�i����M¹U�`����ɲ�K(�nl�ov�E(�od�Y[8k��S�DNf}��)�\��4gQ�b��\Y���Kp�<U콮�A���V�>�/F�jK=a@ߵ�Lz�B>��6��SOp)���17���z�;��T��1\�1K�f�]�ՠ�u1�)-ypsˉ銠���t>���YA�Vt��O�Ú�;���C�����^:)j���7@�ѓ�𔟟YႯz�ް�.ש%'t��+�^��1@�eN?J�����ϵ��x�I>Je�i�]�6=-}=~���e�jh�E��TAg�F;`�^��"�j�ܬO�7n����S�$R�������6*X�һ����V�-T�		�o�W��w����g�K�q��Qhp���]��l�V�ݙN3��'�z�C���عI��&e��]ʠ�����\�G�:7*�ڵfE��`�J6�<N��Y��q�6�p{�8J#�k�ΪT�+���\�	t�R�%���*��3�zdO'�z�J]���Y@���:��b.��
�Z�P��zs ���r�����.�M�]s;z]q��'ޫ�=W���to��A�b�U���aueܭ��K�t,�dI�=&(�kM��g�1ٳ.Tg����: ����ܥ�Y�!ܒ�:F.#<2,�ك9��"����f�PNF	����%W���S�q�C`YS�Q&��h8������Lkk�<�x����Y�jm\�1�8j�E��@L׺���zb��Z��4�#�s#��7um5�*�AA`m�;s:h���J8%�2Hґ�
�α��Ni�Ro���V*I��;Y��w�ږ�hW�z��eC6'f�o	�n\6Yq�"ʵ<T��(˄���a%q�^|8s:.�d��I�w(x�j=F�C���[�Uo��n�o���l'�A>E������/:tef|7�V _5�P����:X[@��ʾCv����؂f}f�yr���7�?�W�.v�V�d�{�s�9�5(�K{��3%r}���:��&�]\ݏ}��|7�>�ʧ��맡�!�"����&��\3�x�J�+n�Z�n)�Å�.^V�qhy�AtxhǮ�Ч��R���/X�������O�N�{f[�ˎZd�{ӝƹe^�>Y��R�]��x�d��#��t�'�S�����ܥԶ8f==[Aة�scT���28�y���W���/��D�Ǿ}{��g�z����f�
B��x?�3���n%�q�ʕl��|l7�g��y�����O��>������'��B�uad��
Ύ&�us�΂�]g����i�� W^��D2��!T9�=��Eĸ�X`���ʥG���������	#Y�8(��zQ��Ч�o`,����*�s'�{�"��2������g��� ��MEtY�47�R�y�i���dx��l�f���um���^�w|R�UFua�Q�
Aq�D��и�3^}P`�d3�N��5�e�c�9\D���n���REp�l�����9�T��n�i��{`W$��,���.�y4�֑��F��PՍ��9�cv�\=�t�F8{�NX�u4�KT��o�n%��U�O������b������S}�ı��[3����ԭvl>>"*:.��Q�ݰ�S�F��O�%�2,�K4Z��.yb󮪔��-�%ӹUԅ�։��<��s-N�u��e�Ζ\+�Q��S�Է�!��gs�B4K؛�Zt�l���f�ę(�:@�Fj��j��ҫ��3�K��AN��[\;9X[]c�`Xuڝ�#G�f��_	j�v,���Ϊ�
��z`:��q�ͻ��A)f�r7��R�ӺGM��>�Gv��As��ۼ>�|�^�,q!^.4�����:�7�H��y2 M����G�f��/hOQ��.e�j�R6�:5��%�Ò��.s�Msru����3�uX�Qfzd��t�+A*�$��N>��W����lu���m&�[K����9`T�HE�@Db��l;�tup�yx?��3���lX�Wh��X�Z7�����t���|�e%�`(��wO���V lA�����R�\���j����r�lh�vrgIo�ޡ��f�`�}�*%v������{_wS�=W}QJ�s[�Κ��q��ot��"v��]����"��dN��+���h�8�3�&=������m�*����{���b:q��=|\�<%W�A����l�;G5X�b�"�Y���42�p	� .]0m\�1R�0]����������QB�Tfy�'j��u�l��"�	�3�Ue��kiZ����>/3@G	��=58)�5�4k�QBVMq�xq�z��>z�l#DC-��=���LJy$"so�Y�q��68$l:���j��{v8�$��6h��TK�E	�,�jA����9�7�/�V���N���<�gY�����*�C�h43e��.�����"�̥�I���Iѥ��̙Br�^�ٝ�z$2�"����|Y�s���5玽�`+�:t㮞�Q��jg!XXܚ4"�C��4�$v)D���o_�I��:���_}9�\����&�A��둎h�_6���`n����8|G`h�/.1}[]��W�E�v����'�n����po(��6�m�et�4_V5�����og65J���QA��{T���s�{M�"�幹���N�N����8�^lXqT�Jℯ|��yp�r�zfԫ����rr}��5����<=�]�a{��<,�\xU˫`�B��nvxۙGD�E��F�z�7f_�r㾗��]<�Jʙ���B�V��wuL��W�9�ߏntY�ƫ�ON1ԍ�2����P�O�Q��$�q�1]j��f]�Ժ�\��yW��t�����//�xVbZ5�8-\cD"J*������7xr��P�t��O�Z�#�Ѩ�����l������A@q�t� dB��mB�\��[ �D�]AKW_�٤ U�P� q��B���ꔧ�&���V�8�4/Ux��<NR�o��0��с�_�V8?������p���Ld�۷�PZ�ƨW`\�}���h��=4��j�JD�,��f�L�7�MҍȢ�l�b���e2r�(4dY��KYpi���ZR�$��;����"�v��{�V%����/�y���o���3��}�h��/�INU�ioq�;0�SpB�6��8�{ѳ\�.�F=�D!��+p�8�#rf����Y�D�kT'�m֮�X�MI������P}]}��i(���/�y%
�mɛ!L��p�J�sW9ee4�`���`�w��T�u�O>�ۄ��N�b!q��]!B��@�@L�p:"�8�-�FdduIt�$���4�b������Hx��Ԋ�.w#��T0lP���7�F�֧�4������ͦ�7���UL��i'�z����Ժ�]�����)�6k��7�����OV�UJi�̧~�ʷ�����|�w�[����i\��s357=y�|��S9|�L�޵��M���>�r��nUQΈ�3w�Ks����S'�z���X�u�
���̮>�8n�[=�}��R�G����M`��cWJ�?<[�Ajڧ}�{p�t�!�ik���}l�� �Zqh�Vw��ߋ�֯k���ûy��1�LV\�����XcI��fֈ*um_�N嬧�pnL�4�R̈�ug?^�]:���F�[:n���{�K9�Y�ՙ9��/��Zd��x��jLN��ṧ�V��/>Z��:�t<�1�Nut&&��u�;W}���>�}�v^�Wځ+��8�g*肘��w�[!�m������*T�29Vp8�+9o?� M c.���p1��j�%�b�EV�(����	1IǊïe�wWu�e��&�e�'�����U�F���W�C]�.�.0v,FZ�Щzp,Qݒ��v�7x�a���vȸӮf�;S�ʻ��l������y\����4�����,n�k�X���T딲2%V�ƶ�8iU�t��w"�tV�����LXy�CY����5��\����ۂ'�gm!MTF=a��K�6>�8C�Auce������}X���w�3M����`W�҆[�B���]룕�T�C[LV�%n�=D^�>}�e�sb
���L�7W���:�\���j-�>��Y32�gf�x���r�y�ZT4M*�ʖd���wf�xnN/3qm����lՓ �Kuy���
h�7)މ+PX���z�Iݎ�d���X��2����1t�V�޽ܶ ���Hvb�6�!,]o-�F��z�t�rUOj]ʾXJ������&*�Z]N�O+���"��Gu�%��v�0^u«;4�ݙ0Mw��+�QC2���b��ڝ��>i�N�N%t���@v���Ͷ��WH�."���2c��gQW�{{�
�q[Fd�]��I㫕	�w�F�����P�N��w�ͅp|ڛ�ՍU�)(����QA�C����2�l�BkV"K�Ȗ�w*�a�,�r�-�I�Xf��ʶeiv�ȋu:��Z�
�)t�R�li�vJZ�л��_r!�6�r"�Zc���:)���7�j���E��O�U|���B��!��z�<aF�z;Xl�5��-�*ح��S�[�ĔM�]�}OT�SWֶ�fCה��x����O�fD�Y�9e�*�%�bt�>��w�{��K�s��ܹrVPw��A>��Avđ�/������F�ͤ���I��ڏ�RS\��YZ�`w���W�.�$���_ov`뿠Ƈ*�b-u��������\�I����mL-��Χ�4q2��2�����>��u�n�ė^.�f�wT"����ɧx����� ���� V�D++-��%&tR�8�U�l����b ���#�"�Й�T�eʎ�;�w\�E�"�Y�:��w;�N�-X]��/S�we��*�4�\(��Q��"9��U�J3"�wf9��ͅvQ:������DpԦ'L�郓YK�w]��u
7q�D�AVL�wG&9'r"��s��s��� ���%Q�p��xBTQZ�.zĮ܄���T��J�B�Z�l�G9fd�9�)j]��r�9J�Qfv��燙Z�����]��T�ER��:�"��az�åWi�xS�A�,m�k��!4w`�{'�%+������Oױ��U��R�=M^ެ};���Җ���s$�do���Iϊ����ԡ@�Ѕ�h"�X��Y��.��#abO^oG<�' �rPk����|,L��!of�h&�]:�[ηʮ�!��b#���8%}�A���+��v+��Kۘ�Zt�l�wE���
��2���ħ�8�y܏*�Pe�35Ӓԍ��t�֠s���#nI���͝;�{|���}�^3���sYV�`��i��\r1��s5�gR��E�t�K��xo|��b��`��!�};���͝ꖳ&��]�;(%N�Ǒ\�)����"=�a{�ք3`Z���=N�RB�sԅ�m�.]ү��%�M���j=Ώ��ǲ��w7;���v�q�T�˒���QΖ����9v�b��d��Uۭ��c�G���R�L16KoR~>���wp����a)���w@��q�=}�%�Դֺ�]ܬu�U�ڝ: �I��\�^Ыgerʘ��G����}�Ua���_)�y�5���3��QL�P=)�L>3�u���k5`����#�љ�+kzU�ŪVy`��.yl�:��M�f�K����xs3Z��[��^�ut#є'�'*w�3�Z�s6��s�7)4�8��1��8a���G�W�Bf�;K��wKm^�8�Uv+ѩ@��e!*�Ӣ4�ӽ*i�y�Z|y]�����ΰ��fa) ���Q�Ȕ#���r\��뜩��N,Ԃ�bɔ`M�����4-�R�⠓�'g�_b��s��B3�2�8؜�-P�©@�#��0<.S�sit��a��+0�@��Q�t%]5��f�!�y�+�N���(��L�w��/��qp1T����W�!=&�f��lu��-:+�����^l�3g	��U�0r����<�j�JP���}�r�\������;U:'�aT�N�yLqm�x����ɠ:Z;�[.뻃��
���e�0=xz�# �W|���%���s���*��S��,1���QI�Ʊ\����K4]ur�ʋ�Y�d�`��X�bFz��\��:Y�(5��Mi���vf�ګ�[��qf'
e��\��fo<d^[<{�ނ��f��i4�<]�ڱN��v5��R�$v�-���Ȩ1O
����4�Y�`ni�粆ȹء1�E-�g��-*k�c��h�.ě�(�w)�~�0����_���=�Q����T����*z��~����f�sC��d�7�T�Y7f�L[��9^^b�~;=�'zq�����}8!&iy�S��GEX����u���G�T_*����"��4 `x��|��6����9�|=�q�TT	�}WjbўG�����Q�����9ڣ�_4PW*G�3�M��6�4Ǽvml�)g6q�g���.��(p�E���k�f�]�s�M�������2���	�`���Zm-�P��S�N���>,�v���Y{\����9�3�QIe���͊v����=2�j3��tTq_���Rx��,[���1�#�)30�����s��Mkc���A���}�A�5���:2j秖��Q:rm>�9���m��a[8�����C�Z�a��\�n��5��Xk�S��H�2���s��Ԯ�so����]����Ѻ�i�]v�9r1\ԧ��LП�V�znP���+��k`k�@��#��V��ԍ'	���n,O��3�>�[�ӧ�#��l\�K�3�7�|�ܓ��v7{q��7.�v�5yI,�ok���Q�i	N{�N���4�vE�N��+�^.��v��%m�R��v\o����m�^Vt���`J˲�:��"r{ �����:))�� .}��]bX�kS(�[w�l�7ӕkr���X��*S�����8�T���t�S<�� j��v8���N�YQ���ݝ�5}ڑQK_��n��R+������z�Πb�->��U����w����/�,�K��&��]��V̶
�5��/_���S_l��#тu��Ǟ%���&�7E1{_e���#ܱ
��?w|~yZ���cܩ��wt�I�V?M�ws��i�;��x@HJ�gѦ�{'��4�-��{�n��O2Z&PhN�QC�A�" |+Ɯ�P�泃Y���~�R,D&/����2fD ��b��w�r�U���]]O����W+��]��ݦ�㰲{���'����Z2��b�jm�
�V�֣���C˾�ظr[���V�7j��J@�h^;�M;*>�=���\��i8��ӌ+C0��\P̮������4B��N�+=��Nw��p����R���vj��u8�.Ĺ�wU�����U˾�)e��*X{��Ri@K�8	���oVN���bJuw4�w9j�zmڿ,U4�kb�E���zxs��#{����Q]oݬ��<�)y�dW��len�r+#pw��gL>Jf{�^.�FoW�s���u�ێ�k�L�˕��Mn�*d�<����~���'�hz�(�V���՗���G�C��j������~�~5���fz��PNY��L�~�2�?���s���Nu:���6r�7�\�Fj�fq��i��%ysCD��F���T�YS0�=�]�=�J���N�ܔ��(��^��١YۋZG%+y+�N�ֽ�7�	�FR"���&R�C�b���Ux�N�u�Q�XO2�Ԣ��30�B�(�h`��p�o�x�vԱ��q���Zz�,�ÂP6T5�i�K�U�C�}1.̹0�v�ZY,��y�^i��0����҃w�r7V�S����%+f���b��m�+rɕ��͙�;��|�Wn>.G��u����OX�k���=��l��olXP�9hpHQ��}�,�S���<!4G,����9}V!pJ�}�4?;��;+�o����Ah5e���ՙR�vNR�1������)K
���#�Es�mAJ� мv"�vs(�7������d��4V��!4�V�_
дf�����1���JmG>ȝ���/����z�9s�z��Yx����_j�P���>
��y]�\ϱ�$3֙�\ts��t8S���uM�nb�[�k%��l\�L��F���zeZ��먥(�/rqRG�z�d�m
z�q�mm-��z���6�[t��>��bX��NE��T4��r��
��n|��S�	�����Be������]a�����)1`�K�oZewLU�򻎄��
��˩0w4v�b�06;��œ��b���2��ю��ā��	!��Jm�ǫp܃��v��W���gp��>�۝1�k���xLغ;V�S�k�O�a��۽Ǯ�_wB���K�]�ǜ�w�
n[ꤙ�^iQ�QyL��y�E�H[7�h���]V,���:V��eܱ��A�)�*V�W��Hi��P��D<��jDZ�쮀 ^���_S��#�C�N	B�45�5r���VPHlt��:*�HƮ;��rޤ`�	ϋ\(s&L�!2��nq8�n�k]���4�>N.��u����)OqPe��X]�s5{�c>��՛1�SAe53�}�%��#ʥP��:E�lH���Y�֗	��53�D��U���i�n��������^� �����y��+'����egV��Ɔ�=.���F����MѹS8(��`G�ܵ�w*w��I��A�9�N�u���4bx؍�fr���0�7���7/;�kf����:3��VXUf�LV�D����f� �S�K�=��B��+3�{�m��\��_t</nM>�w�\ʒ�Q�	'�Dy�u�����y5��]��7�+��n�u�"��%�u����2i��
��0�U:3В�,_b�>s���K��I�ۇ(.����3�o�vf�V�=q\��J����)-ޑ�eDL�q[8���X��b�;��>�N��{��ɭT�LT�x�:�w١�F6֮�N�?n��u�oL�4�f��m���K��V�s��q����vQ�yϫ�l����3�7Ow����y��=����T|_y
�DvX<��[�I�}N��R�k�0�q��u(ԂXha�j;L1
v1�#���l����0wU��L��U�U���qû��[�*����w֧�#�D}��S��Wܜ�\��е��cw3y���0o5yS�V��s���
S���I�k���L�J:�ޅ���h�DՃ���K>�W�x65�����~dG�8��ݗS��%V��'L	�T����"BP;��!�X��W(�w/t7�ucD�sv'LOG��@\p�pX�4�W3S��ݤӪJ����R��<5עjv����+���*���n��H˨�Թl#P�6i*���c���qp1T���Ѹ������q=i�w��%���7/�_E�S��ݾF)�	^B�L#�rf������м�̵���KVŻ�lVs�7��9BP��K���v��̋����o�{�l¦!���N�����N��st!l����f�:���5��c��Bǽ��-CY�e��-"ƽ�u`�}K�
u��/�9�վ��8�u5�n��r;���ц���;����b��د�W���x�C�
JI$�I���"(�YC��A�x%D�P��L>%(Ɩ(�*n̡lO.kV/����T5
*�*;c����q��ݟ	�)�?���Y��_}Q�]��Z�y�@DQ�A�|���p��������j�i\��bT�X��s�e�c��Mٵ1��fp
,�P�R�WɶZ""�?zk�;��n��}�2�Q�8UEP�FD���6�r���@���� ��r���5���]���@�;=H��@<����� �q������H|�~�@9�]&��)z�i�Z�JwWF��N���$s��ʯ�1J� �?,DEf������=���� )� FTCFZI��B�/��E�k����8�M���ǡA��A�A���߉Ķ����d�{��sK���[C������_Ef^���a
"�7�h�FUx�7�?���o�L��68R��@(�����|�t�=��Np>����<7�r�<{}G���9"�<�Y3>�WP���f�y�s�!�R��OA��AQ��DE}��3����P����2kP�s2.ظ��?
�
�8ՒB0}�V��O�����0�r�s"�����
�LV���C�d!wT��@F�)D�"�-�B��?� ��<�'#Ө�	�� �{�>ls�����>���ׁ����?a������F|N�@�8�շk�i�<D<t�ǎ� ���(� ����'=iJW�����"�4_���ͩ�}S�i�c����9�s������1tȎ�P��بBV�������yz6�/�@hG��q����3��������}�D޳��i�tt$��vX�fCѐP�6�� j�Ü��u�s.���`�AQ�`�Ct3����]{�QD��v':@�[v�����f.dB�W��*��y	�|J��r;pr���)��A��