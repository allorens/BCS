BZh91AY&SY�a}o_�py����߰����  aU��

%EE��� �@
�@RP
���@T@�                �    }$�U% UJ�(  a�@�M�<
HD� ��E(E
>����^����g�ݖ��w	��V��v�Vi�!�k�5¹��4�  �ޫ�/,4����B�p�=�{9�Z�V��[Rn�P�-kR��'z���J�Ѷ�J�p�6Vj2��p�    yZo���@�ß]5��݆Tnݦu�)h�ݹ�<��vƔ�Z(풐��v��h9   L���}`U:э���z��cm���,Rsm�Q���%A���π%S�|�o�@*��b$}�)����g�mO+���c��� ���:���;�����U0z8�Ȣ �e8���ُcs�s�.v��3n�9[
�@�L A������"�� j����q��[}ۘ�4m���N�5��ϔR�@�U
횦�}��3w9ʉ{g_v�ް����[��5��	G t/(+�4�B�:�4([KA흏Z�3�W]�OGsu�{פ6��qRV'� ٧mZ66�k������$�h6{�ۧm��m
���                            US���J�JMi�4`M4�M0��*T�a0&h0���0C`D�*�OT�       ��R!*��10	��` ��ɣ T�"Rz�4�5<SѦ��4h#M46�A� *���(�� �0�  ��~r[�\�߇]uι�f��o����=<�zu����{z~f6<O�-�����3a᱆f���l??����m���c��u�o����~����\����K��}[Ja����6�,��}W�+�����6f��f��>�o�۬����?�����\���������G�?N��������ˋ[�2��ٛR�������f��M0�L��aq���[9WZ��-kmN<M���|�I�a�I��I��cq'���$�Od�I�x�i2��RI��q&7��|�~bI�E�q$�mkR�Җ�ͭkZ�<J��Jַ�I+��Zē�La$�%�I>m}�$�i�<L�K�I$ט�|�/14�%�6�K��I'��'���I��'�6�Y��Rq1c������[,-���ַw�l-��3�t�O��0�I}�$My�$�1'����$����0���IX���	/�$|�O|�eȵ�kiM�+[JZֽ��E����J�eq�Uũ,l�KZe~�q&��$�0�����ո��ղ��iZ�[�u�uL-0���a�|�q$���}0�ԙZa'4���I����I��OS,1a$�Z[M:�V���q�,��u�J�3	�K�x�&�O�c�I�&��&�IƤm�Za=I>�Iǩ�Od�Ɠ��Z���V��.�:��J��n�I��I'7'�=Od�s�U�����iZ��&�\L���O��$�)�yěI��	0��$��ĒMI<z�ǒI���ĉ��L�c�x��ͺ�ֵZ�ZV�M��V�56��<e2�?��I�ba'���$��	$�I$ƒI7$�1�I&x�yX���'�N�+v�R����ڒ����n-$�ˉ��2�M$�c�I$̒|��	$�N"c��-kZp㮭L2�����%&$�I~�I>�I��	$���q�LI��o��x�ϱ#od����RI���I=ifx▶Z��-k^&-kZҶ���I��{ͧ�W�<I$�JqkK6��ձs�:�ɵ����I>I�&��i>�I%�I9�L$�y$�rq�I�q$���)�I�RI��}�$�I�Ӊ=�OSԟX�����r|�I��I<�2�ԟI��O�I$�3�?I&^e$�)q��~�I$��O�Z�ͭl-n��Z����ɵ6�I��>�]Q�<�i��1��iMůSk���͝m��L�kO���'�/���L���I̧���]{��Ӯ����K8�L��I=K��z�%�$�V>q�IoI���b�$��ğ%�$�)<�0�x���$��I�esz�+�I$��8�"�<I&��8�ܞ$������q�|�K�&�K���s-�%�<I$݌$�K�I$�~�O�.bL���x�[��1پLn�L��̥z�^�	_'N��̻q���Z�qzJ��v-+[��K[��ܭkkS.����Է��np����jZ�/S�t��-�ZTͭ������Kksn[Ic���;ik��־͸��2Mz�Ĝ}c	��I+x�'�M�}�����Jqu8�6�6�akv,�Z�4ݯ36�����eŹ��i�a�Jԕ�;�Z�f�i{e����u}L۫e�M��V�gN6��9[)��n3SkZ�;R�q�16����N8��[�[���㍭x�Z�ɵ��q6���ͺ��v��y�M�m��ka��+-�_&���ˋ]M���1j[�8akZ�:Z�[1-�+��ֽ�L���ZĞ�a���%�I;�+N۱�[e�a��-kamrml%�m��1�$�cI8�ē��ORm��ԛ�$�&S�bI'&�6����ORI�a�q3$�$�I>�$�,��I2Ռ/��L}�$�y'NN<I�1'�%�S�<Ϟy�qm���ix�-kem+x�e{�$�1��a��Ia��cI+I%�$�j�Ioz��I7��z�Yē	����K8�I��$����I'�M��1��Zē䱉$��$��I5c	$M��I�K����ֽNV��l쵧
Z�R�6�e��8�$�X�Ē�i�4�ēԘ�'���OW�en-�Z�[\�-l2�fmkZ��fԶ��mjZַ����s$�$縓ē�bq�y����y2��kqnre�56뮻����3+^��㖴�˜�K���ska���gL�{���[��n6�N�[��ۋ]��ër-���'+e+�͖��jt�^�V����6�k3K,�M������پ�����]���1թKM�kZ�1�	>I��8�60�I��\ZV�-EM�kZ����[+��[�Z��ͺ�����kZۉe��5�խ�K*����[��۽�gt�M��S�n0�4ݧKS�s+kF0�R�i��h�v�-�\��M1�����z�.�j[�ey�ik�۬K�L����ؓԼĜ�x����4�mjj�gm'ji|���u�-��m����+[.ŭl�=[�-�Kkm���,�t�&ֵ3+ekmw;R���6êj��ڹ�,RYZ�e�Ҹ���J�<K+bnkL���+Z�ͭkf*ek[�0��6����4�������}�-����-bI���M>K�M4�V-�[u4��3n�����V�s;a�-x�0�Ykk[+��֦��jJ_cԓk8�|����K8�$�2[k��Z�ٵi+Z�z�e�nt��m��Krf��\vil-��-3�$�[`�I︒I7��x�fe'����$��Ʊ$��>�I��m�O�&>ǉ$�k[��J�ٵ����&ֶ��m&RjL���1>I&�y��_fei��m-kmz��/U�i2�~�L$��$�Od�4��d��<�$�c��a'��$���6�m�	$�؞m�L���N$߯|�bIn-��ڲ�����Zֶ��,�$�I5�q=Os�I+e�I'�r�I�/t�e��K�c����m��a$�I8���=I&_I&SI�I��ǘ�$�I�'��I$�N/޼L$�I&^qx��'$ˏ|I9>x�6��&���bIZ����-ŭ�v�a����d�R6�e�fZ�O��֙i�[�[K��c���+-ij�e���m���m-l�+iki��Ke-��[���g�*�G�q�-ԵŶ�2�t�nV�.�Nvx�S.�I�JeKM��K\m���8ʰ�6��f��̥�qF��\�[�:Zm��֫un�Gm�����Qŷe:[L�nZ[Kw�6�.�-7Iu<�ZX^��붛z��%�I���$����rV�mku{�[��.6�8J����LT�Q���sƗ�㮵���mlu��Nm+-ȵ��t�um6�t�l��e+.%.�L�ki��m��Ws�4��ӫV�ske�Ͳ����L��4�-K��,4��ִ�ٲ�f�%ki�OT��N���;��.2��_fԷ\n�m����k����vmIZ�m����ٵ8�U4�י�+[k�w	[��i+_&��N���ַ9=[�]�e���mn8�M���Z�ɷXT��3OF1R9�������\������>s͟_W�yߝ��8xK�Gҏ�Ǆ�����Q���$|I�T�QFf;:��v2<��w����z�����nVVtUo��\�S�����t�+����K5��/�M6�aD�QG8YF�4���#Nb�S�M(�eI��(������dr���8Q�p��Z8p�Q���O�_��Ӥ�a�Ҍ$����s �ޅ��&�t���Ƕ�Y�;ۘ1��>k��/���7���*̭Z(�^eZ:���26�6�[����H�(��G���'���L�׮�5�y�TW��(����6ap,�l�Ĩm�Fun�J1�ۏPZ����Ý�_���Rm��X��3̠�C��`��.v2�N~lI�wO�vtDk������蔓���i��K*�Δ}8�Ov�ۤ���;Ӳ��U�2C����uk�)�x)=O��{0h"�ve���&�-%�F�nSI����r�wķy'w7
-mh�Ec2�h�؏�����a�!T�:zru�H�^Jwj��雄�`c��e�	f�Ε�4�nt��2N�&->=��N��+�HT&�Xd�Go3���Nf�'u.�gӷ���;m����3�'�dՎ]��os2>�/h�ܡ��x��Wq�rw�`�[��HW �f7���a�c�ϙ�M?f癨̑�C�D����{݊�[���*���C��옇�j*V�RSj]o����ʹ�&�n�Vi26i�N�d9��|���wT2������s�Rw�.�q��ٵ���#{{ze%��>X�_}�4���Ñ�����np׳
���[�B
��0�ʵl��,�t�,����CYޛ�c��l�eJ��y�3�D|~ߟK7�<}u���3��G��ܷ��I$���oI�D���
�0��|k���+��=�E����7N�x�)�=�8�'qL>�I�Y92����2���6vK�+�p�3 1���.������N@���!(􁛢^����/�L��|O�Ʋ{0m阯X���p�4�Ѷ����+���9ז�n����s[��f�I'��W=�Q��ǆ��k�3�������]�y�K��o�[|]cgO����Ow���<�� ��{[��g�����ENl5�YH���Z;���Ӟg>p����xG}ξ�=>������ K��Y(���ܻ�νϡ�E�>͞s�f�#�Oo��uξ�t����i���fw�e�� >�>���߲lE�t�I{��7�;��$�s>�x����w;���wwtn�7�qs+W��v�6�7��p�v=y�;U�yl*��ӄe'�6Z.iU�fpM������:�A����x��q��Nd�F{��6^��L�S������g�s� �uv`�>ۯ6������u��v�*I���z�g�mF��Ωuy�x=��{��sw����'g 1u���6��J|x�'c�A�柰.�yd�|K�8iͦ�3n�މUێi$��!���v�YSQ�h��k7���,��aR��b1[�a&�-o��<#3�%��+���KΙ�׼�x��fo��F"�3/I9�=�u���6��i��D�}o;݇k�;~Ӟ23��"�L{}I��x��6p���d�&������@�QR7�8aj:|p�l�p{:�*?<~,�גs�5�'ɤy�6�E���1񦈂O��I�2�z�[6�A�<-���<y�����/���	�-�-,�R2�^>��o0"���RPݐ�ʧ����M��G*b��tDhE�ZHg��	!�c��z��VN��^��wGo�rL/����.��'cG=rק���=����u�U�:3;*��R��/]Û�����ӏ��/m2���Kz�lW��Dt�z|^�޿��2�f��M��ᰩc�}+�w+!'}-p��y��Ṧn1_^nS��\l����:\�z�����V��v������S���s:a��u�:�y���V��=>�[�_L&�ۿ|~ﻕ�}\�`��	�ϊ?`�©�7��	SM���n��dҋ)u�	�bg����8�7�tosN�y��n�f�]ы���):P�6��9�kjEbȄH�&���oOM$��ws�.?,|����z
��R/k'ks���Q����Em��p�y�|iXޞ�iU���閼:|zsY�Qf�lW�4�p����t���2"�:|zI&��{�@�XIGل2t�Ӈ�|n��㧦�2�8||a:����=8iF�8d�ON�~)z���c$�N}���zaW����t�=о���V|��ҟ;�Qg��3y��V^�;pL$��^2��mR��������m�ׯ�1O���="�:��ٖ��$�ۙiE�>޴4\ɶ��"f��ҷ�O�{�
k�_O�===���	�_�Ǳ't�}�$��n8���p�{���I4��(�>}��	��T��(��n���dx����M]A�o�c$S�c����tw� �y{|rV�z����{}Q��f�h�/��#I�~:�ݺZ��6�5��ϧeݨA�g5�+ޏ����=�!��N�{�]��z��nf��I_92��_�gY=X����oˏ�t��Փ$�y���a���
x�����_</Fzk��=p���zzfp3n[}��:za�eO\d�}�ݰ��NhQyN����9��������9�[)J��^�����=��)c[(W��,���7�t�y����aَq��և�N������.��K����W�f?(�m�'CD ��2��[vb����>���F}c�Ҏo�-�x[�M)�f�vb����B�;���Jkd^!��'�$�޹��_w��n�C�!9�Nez'�i������&ܺsJÄ�=�:��,��`Xz�D饘���xv7���{X���9�����Y��4/puvM�?��x��e���J/%Xеy�N%��2iÇ^Ir��N��v6�z�Nl9��M.`�Tm$Ncfo�$��OIҊ4���LO[ǹ�x��>1����ߵ�K,�p��,�puS�/��.󈳆Y�����ӆ^a3�8:_|� #�y�>2���8��&w\>�Eu�r.L�C�*|7��mc����DDj'�Ԋ0%�%5��P_`_ln6���+;QM�=����ֆ.�l��sj�י�����ٸ�;k/���|T���\�������ǽn4���H�qtyw�g�ᇱ�#i�ICS���#L���2'����M»vǮ����p����v�>]��oB�[����ϳ���	o�������l��r6�J�<�T�Y�x���}okG�����z�'M!I��غ[�V�f�o���N��4|Qx��e6��s�V21;�?k��Sl$^�(��&IÆo�4��W7˽�_>��6W�Q�^ЗPTӚv�I��^�6"Yg�f��O�����0jH�D��U�C��+�OO�*�A,{{@&>�0�W�-����T�
C1op_,½O��CRS��{w���wO��,�
���,}hӸV>�����w}w�|�Y�p�;��L�O���*{��ޮ2<��n�b�pѩX�t�p�
���7׍�y�[m�s�O<��e���]�l?=�a�H|���|��#�h��$"�ߏ�F;o����B�:�XV�@��V��j*�[yZAny���a�Q=(��A��(Y/��JȫGV_�Z�����G~U��_�4����kT�k����'�O\}��k(-��m=hb:='�T��ǂ#��z��������F?/o�I+��[Q��a^$��&"+���x�-]�x�j/��T�9�5���M2�G�E7ۏ=_�+�r�&q���&���%xi'�F����b���rW���e��+���>>4�{����9�n�O�z��j��?k3�Ԩ�u��y�t$:����c�On5��.��^�,Gq�եw5Ε��g��,=(�=�jۗ^@�|�w���Ҋ��>ziݥ��M>z��>��n�|8Q��:��cJ8zt�^agJ�#�������������?�x������7_l�������?7ݿ���$�����?����4��齻3)\JBMţ-2�u�g/v���?a�N�%o�t�*Ѳ�f�g��HKd�'O��W����x	[���������`�|?�&pnrX���.y����3Jl��E��S�c�n���k��'gm���6�s9?w{�q�ݙ��(�i��,��n����r���g�u:��<�n��y�^̭�$c���f�u�'�[�w9��vݥLWS�SiMǫ�Xnw����Fyp�t��]���|�ޚ����ty�"��^EE�	�c��&�i�lՓ3�J.#n��j��;��w��q��Z�v��z��s�\tI߹	���W]g�r��ٙ�7�<��z���P�`���̛�/)��?Җw��K&].1�򜇨������i�yY�ٴ��� ��OzyQ�*�g���;i���d��'
�Vm&��xI9�
#���׻����� �ii-,��F8p�IY�4ְi
X[,�Qmo1��L�L��m�'b<^)]\�8�z��x�ԑ)�H�Խ�:�ٍ厼#Jf��N-#s&��*�f�ɤ�4\=<:� �Q����P�.C�V�kʸ��k���s����� �G-w{��/�گ{c�-��[�%ҙ�铈밞w*�N�^��g��0|��<��ݽ�{���VG�r1!x��⺉Wb\'^��u��F����� p�����s����<䉈��\������Ə�M{��-��Ԍ�fa��D�2����;�JJ��[!�9ל9_{�N��J�)���s���+�z�{*#��TbB�H�iF�Md����Äv������0������ٳ��f7{i����\L�1g�-&$�TjT��k�K��̷延��'.�����X�_>�a��u$�%����
��\5$��wˉ-����nůf��H��,R9���nY$�"� ���J�<�G���0)����y,��k��+�c��z�f��9shu�sF�f�5%EE�Id��;eq��烸Uo0�{K̑������i�Ww��u��3L0���3��[L��ai9��o1�K�:��g�%N�;%��{��蘾I��
[5�C'5��^I9d�u����{:�5߯������)�Ӟ���#�-��03��Џ:�=���	a�<�#���P��&^_�s�u�:���x��}�8U�9<!S�T8��L�M�s�3d��s��E+<\F���xwӞ<i���~?��ື�<�fm���_?R����6o�����Ϸ���������������~��$��m�9�MF��������,�ʓT�~����3�Ի������W�U���򪫘����X�j�݊��U�U[�ʪ�W�Un�ڪ�W�U�U,�}*�ʪ�X���b���s�ګʪ�W�UnUU���W�U��Xg��f嚁����n-��Xf��r�9�Hjej�n[7,�j�rB*b$T�	����o�������n���u\�UV�ʫ�2��U�U�U���5W�r�j�5_UU�����yUY���UW+ɺ�U�U�U��j�ﾳ��UY������b�����U�^0�3ŶQ��Q��c�n�ܛ96KnM�l�nMLάc���[�*��yU}Uf�*�ܪU���ʪ�*��^UU\�UUr�UUJ���W,U*��^�{UZ��UU�U[�*��Y��}�UUR��u�U�U��UW%Y���~���cǈ�ܳR����:�(�j-mw�w�ݙZ�il���g-�d�Im�n%��GZ�չ6��9l娭UB��E5m�u�Ufy�����)���j՗w]9�M՛�|��߫�7�3a��[����?��?���?33��}�������������&'Oi2�I'�$�i'/4�|�&�N2�ֵ�l�kq�u�Y���$�I�M���iM$�I�)$�$�iǮ8�6�a$�I&I�2�����ۋqjK�ZҒL��$�$�e$�$�ׯ^�I&RI�I&Yem4��jR�Z-iZ�R�J����KZR��Y��֕��V�M-եKZ�R�u+u��k[+uia�q�\qŭM-'�RI&�L'�<I��K[�)Kt���m2Z,��K[em-k[k[��jp�G�C�bf��`x��;�^�֤瞹��#�=m�ז3lekn1��)8�9���ۈ�z�s$��m0��/�n;FT�S����tv��q�"�،�Z��P��g�����L��e�h������R���K�d��[��B�K�eE(�μܭ:9�L�
N0.+qv�:���	۴*Bf7.8n�n˧�i7�^MϞ�^+1��sN\��I�cYL��}�ۮI5�r�S8��G8����[e�W��{c�]r�Ζz2ݖ�2f���d���DC]KQvlS1F���k;�ˇ�ոj5tדq�أFo���;9ߎƝŚ�M���ȗ�ck
vYm������A�-G��GO�+ʹc=�Up���W<�X��'m���MN�8��pNw��b�'�����&h�JF՗d�[��)xkRc&�È��9e�-c����Bc�\�n;uL&�.�du��Veb���,�cu]�m�X������ϟэ��v#*4��ذ��)g�6����i��\����S���v���SZ��"m��nפx�ϣ��9�l݉zcq=�p]���k8��Kl�i�a�r�2�C@�;�S�w	�W��ـ�j�/$M��a5����3�8r'h��el�H�%��و�����F���<[�ln&.c!�2g�s��8L��8���Kp s������X����h8]�1��%�X���W5yd�9xqAk�ރ�e�mq�Ƕ��^óZ�׋�Ӎ�95(\dD�|�Oo��X�8�Sq���釫�k(���&�z�B0^������76{Ys��
bVl�qu�\Ee� ��p�X�/~p!ĥ�����%�зnN�%��8���<�[��k*�@�ts��
]l=�#�7:���Y6�m.Z��Eg ��m�(\�z�;Gh��>ߥg����Aȷ��p���\��Cز ��Qq&������7��'d-εm��q���9;F��b�o	�`z�rq�N��}a��mn�Ž��ŤF-ң��<�g�hs7[	���5Y:�s҃���8hTA�tPP>��L�j\����$%o+,5�v�r��q%�q����U7
l&�&,t��^1͝���xxz{�i:w:gӍfv���>S���h������{�m�ku��Q���"/c���;:ش���[�YL��
vv�܆�qې��9�ۚ���g,�"�\R4�˕A�r\�eLj6��D�Aö�ۂ���,��)qr�X�|n�kb>�c�v�����s2���m;D�vY���&��r��p�[�rf�A�b���g�D8N�-ͳ#�����8�h��۴Y}IX��N���)��*����<)�clEҼL��u�ܭ�n,MH,%t��k��㧀l�+V��g/X�3��yܾ�k�+�p�E���Du�WR��m�Sqr)�;� �?�=��{���{��9���=~~�����{U\�9��3�����{�{޻���{�ޫZ�B8�6�μ�k[�8��an��ַV��ť�����+��tySX����ʶ�I�3�m�%2K�Za�)a�n3M�I�����b�jL%&F�FҎ�G@��rx�t�s������a�ik�ܖ��\�V[�̐�Uh���Ww�{���X�����:���Cz�8,��R:K�kk@kx�1����M	�3w�{4LsK����n�+������v�bPq;�O�J��w����LAG62*]�h���s~�k{K�M�j�eT�,���VY�3�r��x��u�ZL��V�<c`�)�7;��Ʀ���Vi�;zp�t�y)��5�B5O{w4F���l�g�nQyA+9mLI�rdԈ"�TN�k!	�M��|���ږ�5�b1)�Gaf� }-<i��MI-�SPڣi�	-V��'��]m�sJyNe��u3�v���`�qE����GRj%ԩ�MIb��}��_�!A�H}�~|�>|����2�b�̖�u��Ջ��k�-����;t���J���\)��RIC1xK�'T�&S���Z�&k���Z�yn8�-����Z�Zַ�Җ����j���`������
n|�3��Od��[o|s�<�/��S�0�)�ޞ$c'��xt����/%I��eR�)-��*ڄ��d� �w�<��8��p�-d�ѥɽL��*[M�J�L��P�@����D���ʗ��|8W�K�I������f:�m�l���{M�/+F�kd���Ӽ0'�O�cS��7ߤc��e���|L������m'��I8�>��D�D蘦����DUx�	ZY,�gU^��%|ǆ�Ǘ����LxRAb��M�^s���5�@�@�	0`�^����s*�歈�ѽ�.Yz:�	�$�ğO׍ (�m���$���v��4�<�^t������t�y�J�j��Κ�:�&q)y�������_r\�hb�.�tT������^V*�I`�f*1��$�^����e�c7��#*m$RR���N-�^q�Z�[����խkqim)i,�˂a�Ԧn��0�s�&�����O�?)�ye���QǛ�w�y�S0���F�ɚ�McT�����iW��ȖJ��S���,��M&#-)Fb�u��a��+�I�RMA�5�^�YS����^=)�nNx�!�!�����x���>/�|��gߪ��}�X<�Hxcs�a��i�9J~���y�3��z�E��9S2�z"c�ن����Ϟi$�m��OS�&�q$�L(" ��b�XI������B-��ۻ����G=;���2i-�V\ɭom��Ưb=,�
1���7(HݦfeF�I*Wx��1�{{{�!q*]����!	��LT��<-9l���u&)�I��Lڤ��nm�NY�����t��z�A[$.�U*�<���#Ї� ���Y�⻉��ߨ˥"^R؅7c�I����3'J^hO����Q8c�>5"FE�ޞ
xuN6���TMc)L&<���vg��m$�G���9�>|1M����8��GD���.���$���܂nc�Bp���ߝX��s�ȩ�Nz<�ߎ	�~�����Z�e�,�	��a�2�yG�:(����y�	��~��ʱ�+/�B�e-���y�mŭKuն����n-��Ya��!i"��LN�L�mN[�7�UQ<���3�� �;ojVۂ�0��1����m�q<��0���i����L��,"|�)�������<&�y�総9�����!��?+�^~Io��Lʉ]u�H�T��yk���أ��<7A�>1�:^B�~FB5�8��(x^t@���(���K�N�fgQ��m�V��q��e���Z�Zַډi,��c)��*q4�D��U��O�g:'��|!9����4��C�����nb�nt��f}s7��37(�X�	�a��s>��<��σ���(@wz�H��9u,Ҋ���K�\�:֌���z:a�ʋiL�E2��l���ģ����Fq0�{6��13)�����r0������:"x�v8����;��֚k�89[M.��!�[,J�un<��8��Yn��ַV��Ŷ�ZeL2���kE�c�}��I窨N}�>��8�羲��t��!��NQ�^�;��==)���?oIO�m]\Yw1��p�\Ւ�=���y-Y��9&z��֖�駵m���ZcF��e�n�<z7�n�!q$�B"�[6��!3>���ɂ�����u-��2�Ts%�����mڽT�Jk~�.����w�����t`�̘�gƗ���y����3aJZ�l��F�)�c�-֖��8��Yn��ַV�[u��*1������֋�Ȉ(c$�\���i);UXB�<�IE S�*�'�1��̞��lkiI&�f��2��k��A��>E#D$��W�Nw��i8�D}��Cf7M�ى��\�.UT?]��LH�HHH���p7���HP��@0���D�U$��2�4��-v�9�6��/��'ߔ�7�!l$�K(�YG�F��a�
ylF�Ҹ�#���F��&�sƫ36������)$�(�1���ۦڈ�l3L��^o��c�T��� �[K�3q�����ؚGa�m(#ܼz�J~��E1�P��#M5�%1��Hwɸ�m8��g�C�tܼ�1�����~���$K���1א�t䮤f-�v�ރ0�HÕBI��1�@"�r�XCsfm�n0�n�t���y��{�l��p�|E	xT�F�s����u�]m��H�q4��>��1��[�g���&��;��T��~���p���/���B..�G}�lw��s����=0`�|���S���K�z'����Ie�3�����w���(^I��<�[m�R#�)JfwS=k�<�r&��wN���/C��Ӯv1��8)�0|��N�A.�����h�][ؼ�K�=�}_O���?�F S��a���4�Qxʪ���F��o5Xo	Tm�fg(E�ʒ�i��>p�0N��y��d'�p��i�Lң,ƎR�۪��|�����|�Z|O�W�U<�'��/1�Ϙ�ט�u?)�1�m���K��ʷ��<�'������y>y^yZy����]u\qV�щ��y>yR��y>O�W�畗�c�+̼É�ͱ�^c�+���1�+��������\O��]O�kW���akbީ���Zi>y^N������Uǔ�ʏ'��x��S/0�O�/&^W�O+�>V�W����؟+�fg����|���y�e�y6°�O�W�W�V�y�'�+�+/<ǛVӤ��m�y�[
�p�/&^�򩇘�t�{���x���^yQI�^R���e����>J�W��<��)���>V�y�6����|�y�������o>aL��mj���b�<��V�W���/3����e<yT�ʼ�y^N�����U�V�'䰟��e�|��j�z��_&S/)+J��W�����q�y꼹���/[kҷ��̷�nuV䓠M"Y���	�������N�N�.#��a�+x�#e�����(3r��d���Vi$��c�����	��~Z=����.����D͉��(�d���*�V��=���rK$g�|_u��yj⊄�>0u�H��a��)z�>ݑ��I�#�O�:Mm)�;a��ԙ޶
X�.����u��$�K5s-no��.�/���o�U��}�u�׾�~k�w��]�{ڷ���{����w�{����s�����z�%��u�]M�Ӯ�q��N$�N��%M4�+Q8�U*�D�4�6�oJ�8��`�����;L��J�R:�zjp�15��G�#�n���q��x�x�<���fӍ�6����s�γ{q���q�C�r������{����y�Ǘ|�7�;�8���&���1���"F:SIFa�C��âr���Y����R��������:H�rǍ�>.[vaH�JG~�Y�{55�G"[DA6����ku[<gn:-�m����Y���u����˓���l�|=t���9��nm#�x|�>�v����x�7���c�<��><��:<9���Y)
>H<�{z��{M�X�i�xx9��3�<+c��:�՞n	�� s�ˋ� %/�Ⱦ�d�ɃA���m�Cל�U��x��o/o��:��O6>��N��Ԧ^wl�%(�K11�[<�_>|덭Ӯ8뮸�<�Ͱ�T�L:xvܷ-�|[�u)Q
�Uy��s�D<�:M���g����s�����[S�o��zt�鷑��ݬ�7�o��Q�M��_�KI�%5K4�����q�S�hJ�k-k��=�\%i���ﶚ��E���zZ�{B������ۑ���D<��m�sGK���#̕�gߪM����p�#��t{�ql~M�y-�M�M�7��q�;㈖�}8;��Dgn����j����cM��)�"ҍ&��a4�qJ9qB�!��0`�����3��yq�f��v��m�7������x^_O���k���C�bv�v·1�t��n5;Yۣ��}sn���q�Zv���̤Z�d�p3.��c"�]��t:���!�m�\֛��.�ON�c�v�s�ݶ<�xOSm0��a�|�κ��,�][k[�[���l(�4�4�W]�1D����A�a4�j�xE�b)���Α�����y����As��n+zv�:���+�Y
��<��wgNG����_��Nx�G-�K�T���OY�;���tZ�t��+���n ��c��WssT��%J�y)_�,��`��}ѕI�j*�"�
�dHR�ڤ�[�{��1c��p�Cݢ���s�E"�!��!)�	9��N�vGqG��b-P�E#05i�4�Ih�<���D��ӈ`b)P0�R"R�o~��珴�i֘s[lG�ͽ[zM�o���GRv�qsqJ2�q(�U�Q���ɤQC�#�G��%W��)�rfF؈C,D6�b-���2���b�8:�Q�J��e#I9�#	�T8hC�~���_79��4�O�7}m���:G�Sul�n-�ӧ1ӛ�<�"��T�pT!�L��j"*"9Z�L��+]�s��:�j\`vX�_�,AԻ/y4r%���2�F0>|������'��ӧˬyM�� < ��xz��m�x����n]m���|v��)�>�����9�i�;��8},<�q������v�r{p��7�Kg���K38�jII�(���y�^uo���\y��mkuku�^m��N��N��M	��fȥDg�6��6𜰻�t�q��m�Ǥ�H��s"�|�ޛ�+
�a)�Iz%(w
�r$b5�=&�͖�N�;�4��9ǜ眐'%���%����m��|�s�OoM����|psC���n(���L�L�lTA��wJd�k�4��v��w��ݸ7��������8g-�֘�YJM��\J5��mՎ�n3��\n,�'m1�#q&�%�JɈ��a�ucݶ��w
s*���<��5��F��v�u�f�Y̳��v���0}�Xy�6�������O:�ۧN��c��}8�f�q<,�lu��������(�f�|�\{���{y>t�q�u����8C���Rp����H���~/w8�T��[J$�Č��e���<�;)K��~��K1�!��:��j:�n���V��]|�ź��Z�Z�m֞a$���a�z���y
�j��ψ�������(�7�l���'�-���ե��ˍF�R�$j�E<HƇ�s|��O9:|k��KT��H�L.:Rﵪ����l��IǦ&c����$�I��Ov�[j���X�O��vC��;M�G��y[xGo����
s�x ����=y��vt�� � �R'2�'i��m�f&�N�y����F"b+ޙ�d�%�j%���#��IF���H�`��t���9��_���É��|��:��"Xr�%��L#;�No)���w[=��ӏi�g��p��Kl����\���x�)�4ޓ�xys$o��p�u�-��3�ӜS��ĳ�H;؜���T��o���4pI"�b0�u!�ÿL�IRY��!��TC0�&�Ĕ���i����y�뮾y�κ�ַV�[u��I*i�i�w��Ntd�%���	+ȋ�2r%��!�T����7?Ð�{���"�8k��w9�<��MF�ޑ��]�������<��uQ��\Q���I��l${�ߩ����l"��e]�hY�������w�g;��UQ���KI&`�'��;>S�yNN-��N�����XfQ2�n��k�&#~{׆+9W1��^OKo{Y�U��M���G��{N.u����ޞ�=kg��RN��(6��%*���U_����G��H���ǂk,�2L��4�yְ���J}����qLᑔ�����ҟUUV��:f%OE���g�zNi���ƙ��v�u��އ�o���x���ül G,��-�_��09�s�8.����a1+�Q�Q�L)+��0e,�34�q0�M_�5�`۴��&�%uHZp��m�ϟ:�<��][k[�[����%)SM2b��蔿/��o��É��2�d�?:.4�񳊳L5j��V���Z�+z������qd�c1<�q��8�:��;y3�!:�"݊���<E�';�~�_~=떛LQ	܉ ��!ӫ#sH�
�%�y$��I�ڌH�:���6����K�SA��6{����	��F�/�@g@����A�����v��t�w�\qc���;�a�Ι�˓s���d��ryyy^w�����t�[>��Y�é>mP�7��ĳ1�����8J."a�K���jk�Í�0�d����x��N�ռ=�>�x]-�Q+�*4�ۊG%&�R;Ϸ�V0|��s�����l�9�\\;�m�u�õv��8���΍,q7��n#�<��S~���On����T������3��޺�{�ǧ6�x�Ɉu�#|RS�QD�׵�«��d�Q;o����-܈�vIm�f[��kS=�zQ�"O�Rc�F�T�i�����W�<M����ē1�n�5T��Ug���L<J6�a1I���|��uמx��y��խ��i�	)��a��3ʯ�����N����E�<��;u����ι�7����q9���`jOD�QL������&!��s�g�ks��'8���aB��'����Q�Qi�u��g0y.D���nOV.��prt��n�4=����ڹs�Wu|�� ��7�����RMJ�����v%����j���J+�=#.%)}��uX�T�ݏ'��f�3�����D�	K	v&8�5Jj�
�Ҥ���D.r�G?l���aN.3X�cN���w�����6j��Y��l[�t�IO9��L|=/<��=օG��nO�|y��ם��n����ׄ����yyݺ�G���:<Z�5<���㛍����Y�=�9�'�>��,n����T9O}ʪ�!�"���T�aڕ�*�_-n��_:믞y�כZ�[���O0J��L��±�UJH��4'��(�A�M�%8D�!8sw��C�xS�8	�#�F������)O1�;xNgͶ5h���L����bK-�������n*�� ��i��Ϛ�cn�d�[�ƶ�&쏯gӺ��\�5'�Y-&�R�0J5�j���ٙ��!���l;cS]ț�.�:W�@�Xز�yR�<����>�����7�ۈ�}{��w��Å�2c��yxD���զOA7��xt�-��.�ޑ���Y'��7��y-��^~�˗s�yo9�<'ֱ��q�m���D��z܄��6�R��eQm�m���
S��g	L���5�f�NG�����s���[��!���i)[.����-�]y�Z�y��ն�n���-4�-;�0��K��1���i�Qx�N ��q�?��>���{΁�S�S2��*�QTt�(�zB&�n>9��<,�֋������9�]��-�זY�P(	eĞP\��em��YLB;�
Fc�;�i)|���b!iu-�ڡ2����eQI���Tb�vXv�>���0n8�FTE%ICje&&	%�G҉�Φ��d�F�=9舟y�����>Ŝ���>\�:w��sY�,����:O]�1�D�A��7�|Ϩ�޵[m�������2�v�ĳӾ��7ƙޞS�VxG��}:��������|'z�X��T_��N1x��n�
�Č�&3�U���q4��O�W�+�e�W�����������Ն��UǕ�故�^y�'�4ǘy�'�<é���ǞW�y�6�:�:���'��|���y����1���<�i��|�Lm�y>O������e�<��y8yN%��.����Ŧ�ոǘW�W�W�W�W�W����^eOL��L��y�u?>S���ɴ��L��&�*S�e�y4ʼ�'���|��8����y>O��Ǟc������*�*������>W����y�S�1����j��1O+�[
�p����y4򼜴�O�+�+�e1I���*%>O��L�:�y[S�y4�'�V�S��|��y>M��M6�	yO'�:�6�<�<�6�>Na�����\|��>�Ҵ���͸ד畖��i�y9yT򼝼�W�e_'䲟��>L|�=qZL��e2�R�S�a�y9yO'�+μǓ�������ۙg*��q�&��L��$�c�"�r�V�5~�?h��f�����X�1§P����SO;Jo�#8J�P���CJ1&�;+����tK��NkI��mx��yx�!��@z\�OkdO�	r=<nq��\[C�"��0X�D=BbՔ�W���LbČ$�թ�FT^�)�!��o���@�	cf��A����mCm�f'!r���Nx�cg��d>yeۏZk���\`��8ح�jU�
(�T��ga��AXl��d1�������"�"1 ��c"&�N�訶3=�0��Y�"�t]��!u �n1���*�^����/q�ߵm���L�������+$�"�!#�!K���M��P��2->o�#��U���	-�]r!n��j,��B��zE��ӳغ'�<}�ӯ�xukNBx�����
㓶�A�m�g!4��̳I�G����|���>�!)AL�
^�Ҥ���:ܼxc�<c7=8�[4�]=˵��f�c���q�rqd�*5>�IP,'�p��6Fa>��y��Ҩ��Mm�+�-�c��{�&2uݽڑ�1M�1GH�c���n;]=^`�78�ŜkW'�g�b1��&�9��� >�����ߗ��}��}��w{�{�������{���{������^�?�k��w�㽮����o�ֵ�O̴�:뮧u�yky���Ví�����t�:~��yY��3c-l��]!��E�����挥F6ػ!�w8���>���%ɍ�����ă��KDi�݌�A�Ce�Zݍ%K���+�k\�Xi������'����:��<�CF��g36�Uh��WY�3�#EF�WU㋧-֐��bVrƑ��)y[$]�����'�� �DI$�5�XG�T�K&�%�Y���$J�;CEv����6�[��$����VmI.���N��/��u��݌��=�]m��{5�M�[s���#��$Ok�t�FZ�Mb�\�+�	9y� ��Vbr'�ߑ��N�>�V�y�!J��1��P�e��[#&��ْM�7zp�f.���F�/�F�y�]ɦw�����I����I\�L�u(����Q=i�[�R�jh�F�JJ�LC_zf��UV��S����tMkumN'��6�x��XK)I1
��K$�&`�E=�64��]6ǧ���}B���0JT�#UĘ%��ݸ��Y-٤���a]������4�u(Β{i�gÛ�ԫ��_=�uߌ��h�JL2���i�dO�y�������N<�xQ��s�Q�vjJ�}<m�7�zŷ���+xGI�D�<���#È'/����H��E4�I5m1yk_�b��Mji��M���+�Q)y�N���|h�>�+�����m֊ ����ϻ���O�����./!��9by�����qn���<����qթ��i�	SJi�Zw����=l�5�Ze2I0j%��%3�S蘇P�<���"NG�7��qm�}7��鷇�5�^�4�Y��H蛽�å����WH��;-�J�44�d�v1�]{�g�77�d��Ǥ�湷��M�A��&!�Q����%*��S�u0�Q�9���:����A	Rb;�O�o�\�3�����NPN{����奕��+�HM�!��?t��C�&AHe�̰��f�Z�:�QJ)/��҉�Q��:q�/N:D�5�i��o�ë;G�䇚�ϰ�t�9X����
:�&�]�n>����q=y�Ǎۘ�[lIc㥸ޭ��W_:�uPm.D�|�N���[��y���y�V�[u��%M)�1ӵ5�ۊ�t����]ࢄ���"�İ���K~m����Xe/���]:�z{N���q='�g��$���m�	�ۙ;"Q�L����j"R|�|ꑄ��y�1�}�|eֳ'����]�S4W�X���KE7Y�^j(�h���ܳ��+c��2��e���iu���G�I�q���R�v)�z��:''<*��'��K�ߖP������:	N���B�-��NӔ}1C��+�����\y��֓�u7�n�&���t��δ����vj���m��Q����6�i���K�*$�1P�i�_6믞q�y�Z�m�u�:ۭ<�.<8������7��ucI*�U,IJ�y�܎{R�#�<�w�+��cr6��T$�$��Ln��_Gx��-���#8M8�B�QD���ro��˿`,�q;{�d�b�Mɋt�$vӧ?'�!��=1eOFT�\ID���JQ�b�����w��M����_�oi̖v��&�=�p�o/9ǽg���8y�I$����ۍFs�����ie0I-�Q���_v�SX���j)I�J�#V�b*�*�1�L�XS�RF	2��NLE��n%��55ڪ�Ff#l�J�&K1�2��Jy�>�SS���(�N���>[�8��<���o<�)��i��Ht�:|r��}���\�d��b2�,R���J�pR.{����S�a�"�"��<B�cޖ�|N�^�j���j�w+]4��c]���l�Q푱�vt��R!�� ���M~N۱ <.�p��L��n*O�ӹ��fl�����	�D���3)�KYi/7WCt㌊��D��i�Hӭ��)�Tu'�&�	w��e�祣�I��I*�c��}'ã��"K=MF_u�a���%�P��ʪ��uQ�8I�1qY�8�i�e�C��1��a3���L.8���OԚ���~s�Z���,�$��&w�Zb֙ќ7����b[G�}�I㤛a�}3�z2�N}S\0I0{S���絛��F[`�I&�q��wq�0<>O���1n�,��g��Bɳ1�̤=���thPJ?�$���F��MƦ]���e=;����yl��Ϝqż��-o8��:�m֞`�4�,��|����q31Pl{$�?,�9ݾ�)��n�*��x�p�(�jw�Rfv�r'�U�N���Tt�LC��%�q���J+������yFګ���<	<򞈘�S�e�W+�I>|�gO�(c�Ӊ�ǣN1�$�����(|�g � @���!�4��l�����͟��,]�=_����LY�ư�fɈ�����������18����1�9ez&)l��h�O��]�}$�'5�C�L�)î��i��m�뮤�n��Gu��%M4�,��}\ǤcJ�S�(�C﷟����i	>ȲJ�RJ$��v�0�	-�L:l�Ka�>�k�3�b ��.�I��Sn��ISN�g��&�OWɚ��Jp_׷����K�-r�jj,�י�Zr����e��F0I�Jp���b��I�:��3S�����J��L7�j�u�-%�GI$�M�kÃ��Л��#�1�r�� t>8��1����Q���I�>���_�ˆR���4�`�H��%��iǝ[��8��y疷�y弳�����N��I��a$���/9:��I袜A9x�?�'�FM����v4�c�I<�:�c-\�>t��OӖF���k�f�-\�aT�n6�m��D���9�<?��Ӷ�=����8�ä�m�����U�c=��c���f�,�`�.i2�,e�̺��$�aO�����7���"0I�̸��9��R�N&l�&�؁�Tǝ���I>m+T��S5���K�>���bf1�c獒`uy^]��S��d�&4�ͭ�ϟ>q�Z�yky�^[�i֞`�4�:{��ҟKjnX���Z�L��6�D�|s�~z�-�2�2���^[�<B9�#��g��_:M_��Л�/$��{u����cI�n\�ν�/kt��m��C�$8@ Ih5�T�{5�r���j��H`�����9��ݍj)
j�d��I�iCB�D�T��0Xe��!D��
+ɏA�{�*��]�K��O;��;!��Iy��d�1�M;���D�ά��O��p�<��|�I%�ʡ�-�Y��A��P>�4����!��Ϩ;�l�Z��53��yL�x��,�\Wfe�z2��][�I��n�cg	h��rg-����I�a���Y�4ޏ"I|Ɔj%���S�6�pt�]v�M0�FO��iq�l�;��mjaAڃ�ey�7����}M.;n#�6�S�3�d���QwS5?T�Z���^y��-�V�8��y��yo<u�Zy���L�t��N�,�4x��(�K��}^J��&cd��S�LMy��7��Ƣ�$�c��ZN�1�h�����1��ڛ��S��&��K�g�G�x�SS2����&�����ú�����$���a��_B^��)��\$���^A�� �u�J�B$)���Ҩ-�@�l�������	%�z��!�>jfr��v�I*��	��8`����y�����fg�zoɩ�^T����8���N��Wβ�^S�������ǞW�W���'�+�+�8ǚy�y[NEy<O�W�y�2�:�<���<�u^yO6�y�:�u=q\q^y^yL��<�:����4�:�6�'�+�+o+�+�+�)�����O�[>R���L����]W��-ڝ+�+�0��<Ǟ��ںy^yO')�}3�<�<��Ω��6�x��z�>T���~'���|������3��>Z����5SW�W�W��3�)O<�<�����'�)������y�y>y[mZq�<��y�a,'*S������,��<�)�<��m0��9yD��'L+ɔ�O���1���zg*���T�\y^Kɷ�s3�y2�'���i,��y>O�W\W�WXu������c�ϘK*��>y�<�8����e>O�W���f<�'�+��|�S���)�|O�-���v��ԯ�$�NT�)Xy^�Ҽ�=Sǘ��y:M��'_L��1\��Ω��>�V&A���̌P<^s�]<�P�8�/��_���0�5��@��-"Y1�Gߓ�~xg���"/�`�)����^?!����e��2/\����N΅���)q�RxnT�ՂW��̚��P�M��}z��Q���z�/Oz|_��A�}D�y�P�����a�e{��u>��1��iT(;6�����׽������{�����Z���{���Uv�ϻ�k_k��sW�U�_{�{{ޡ�[y�ykq�yo<���-玴�O0R�i����eJ�ɩ��&v��u���&]ffmě%/jg_���{�賐�h�,�0�2�I�R�Z���f:Q.q�FxA����t0'���浺�+v#�ND�牮�(aԁ�[L�24�C���i�����Sm�T`������d�jχ�����O�CB<��.n���ef>/����˽��Ap�����W�+Ͼ�b�ޭ%�6�1��>�5kn%s������p�-�b[O�UKѶZfLQ�iku���y���μ��:ӭ-���L��JbbS�s��d��)�t�X��73<���>a�[JJR�#�q��!�/�sjJR�����[RԤ�ˈ���2���SUN=qM�/z7�c��\�y��$�V���᎟��B�������s�uJJR�V�fX�%���t�e)J��K��aT����e�b|bJR��4��^g��J�QA�~�5�!��-nL9>}I�"Y[�J�RjghA=�i�����K'�PB�r"�^T���b5m��RCs3����R��<��>u��:�<�����[�˭-���L�=����0�=H���	��D�*���o)PR��P�/�1�#$IG��e��9�q`�ߚ�vz�jݴ��7I�	�3��[w�?6oS�t�5ŐIa��	 �"L�]�Dۑ�p����M�Q�/6ס��E��,�q.��K��Bj#���cZi�NA���?f�"�#�����Q�\���8�b�a��,�£u�J���m)J]bw1�k�2��x���7	i)Kq)���RuSZ<ӱ���yIJTq��UQ�ϙc�Rza�
���u)JX5��Ǳ3�4��DDL��:����8x�<y��<�BO4h|�t@A@H|̥+�>/��ӡ�C�Nu�"#�{�$��K��(�j�3��ҘD��r:�ʉW�I�L儥-0��j:�z�mֻ�:�4|��4���:�<��מy��em-���L����3�ߕ(�N��g���yyyLu1�yq��3*R;��*���&L�����M�^�G6��3y8�tG[$�>֣/3�ʆ�I'�g��t.Pt��������xD �h4>r0�D���f��H*2j~uD��G��'�Yss&�㉍���9g>���YgYKI%��}M����u�/���7�����v���L�����M�3�4�&tq�y�|�<�ַV��-o<[+i�!Ӧ:~��ǟFI8�KY�QA ��X��yD���	�8��a���s�bqW��C�RI}(�}c2�ΰ���0�p��w��e����9Υ꩚�������I��9x�-�"0C�~��Y'󱬛B�0�:�l��YXO�q�� �U<�@訙��J73؇�UŶ�ԭ��\�fZS#�DCs�|�59��C��N���e�Ǔȸv�I]��l4�s�n%�R�L�Ե�ξ��w/�IQ-6�	�i��q1�a��%ĩ���&�8㮤�N��u�I�||(B:c���%a$8�Ȋ���袂!������c1�N��*<��K�/�}�Jgp�|�֛�����c�����r�T�����FO�b���Py�h���~~` bQXC�I�il�k�����==�?��Cp��87'S����yJ��[r0��n�3>g�N#�I�!�ԕW�i,9�*��+�Tד���=q���0�wu5Q�\aMaL$��u~��?����س��C� �7���5}L6�E�u��y�κ�疵�����y��[.0R�i�O����V�L���^G����yybB,�XNqW��`G�E�ؗ���j#���o�^�u��$j�OS��S�T]�f4�k�ۖ�I�nzѭ���y�
DE�	 ����`yz��9��\y0Vs(u�BT��a����3�J�E��e����ذ�Y���m�cCy��p�6ﾪ'޿K�x�+�@�N1р������bR��Zq�RH�s)�>�
1��I;�O��)���)��e5?[H�N��Y}�T��f[������M|$�
z"����f��x�/>�OvS=��[m��5U�1�Li)>�MY���t��}��S�R�c[L���y?V&���Xj6�ғѹ�����7��v��<�-�-U�ǋ����m��G[�i&{�Z�{��NY���X��Gu���2��<�w�i��-�m��|�	&8����c/r.�&~�f_)�[6��u��uמy庵���Ų�[`�4t�O}�>��BH��ı���^�PD?��)�!����qt�b��q��k{���II�S2��/�;n;Q��X|��}8�T��%���)Q��i�La���Y�Ǚ��xj9�Ҫ�ҙ�6�fm��//xy������?�Ͽ�䰰H:k�©f?�������{��O6B��e/���fR�}��v=
>q�/y�~�ե���W�?R�Q��MFW�a�o�b���"�qI=��^�Y�S9�c9u��L2�Iu��8�o�uמyםZ���<���l)*i�V4̜��e2JL��n4�8��N�*�؉��8�|��D̽�q=��]o�����[�x皳�,�����ד���|��>yi$�]�F�q�j3u�"i)/;�{���dp4�L�q�Ɓ�J���+�ʙ�p��[f�k�O��K�5K�Iĭ��	�̥��L�T�(����m�2�I1�L����fe�'�`�q��#�*k1�aje����4���ST�M4�V�s�)۽�m���֘��e���뮼�μ��n���il���a��陜)Q���μ�{�QAy������J�8�Ox�ç�����A�x�:�?�c|?#_�w<2[T%��`���v��ʫq�¸�r��3�v%Ź1�[LS��kL��8��U���4��6��Jq-�e<몌�%),a��be]}��x��A�V3�(
4x`QG�sy)��f�7��I8'��;xy��w��u�XI�Î���P���r�;m)(���6�ۧ�#x՝>|�n����I��ORL��I$���I�2�|�o�O�x���I6ٶ�i��O�I>M0�e&�OSI'�$�I�"M�|�q�;I$�$�(�ORe��q8�q��0��0�L�����$�"I4�I�z��I$�I'�&Y|�+q+[
R�YkJ���k[+y�<�^y�<t��ml-=q4�i$��Q|�RZֶ�K�q�q�yמ)疒M�׉<I�a4�i6��o<�]y�aԼ�0������kqŭ�Yng��oƓ�⻭��W�Dq$+���(L6�)�ՍI��6g��)iKޑU��y>��oNB��J)�U�HtBu)�BH,����n�=��J6C��K��e�;��ŽU��gq2zN��%-ʝ�|ӭ�x�\�8��rqRQ�8y$H6*M�حrd�nKv�nI&�B�4�q�a
>'BKB�
�$&n�l���DJHR7^�#_52:��Ч���v�qb���Uv%�W��6KB+vY�hɃ5I�l<�E�0�J�SQ
g���l(9){���N0Iy�K4��fR�����
W=�p� ��E��ܫ��e624�I	{��m��`f����h޵�K.�h.:�i�:�R��&�3�N�DL�2(��67߳:O���W�>q4n65��e��V��w��ln�F��2tkh��;;�e]��F�<��%���=ds'�� �V�z�?enV�י.��`D�v��7Invy�����d΃Q���s.�U	/i|絁o7V�/B.��N{'��vSɗ��h��tvi�ݭd�<�)gȲ��h��K���X�]yT��Ĺ�7����}����g��~����k���ֳ�w����{�U��=�u�g�Ɲu�Zq�\q�]u�RI�]uӬ�ǅ ��ҝ;�ﳟb����֫l�mR�rɸ����ɆS�:��=�x��1��m��`u��YN���O[�	�u�O<=��=��e��5'���`3�C�@cp���ݵXΐU[1s]aul�T�\Z�m��\�q�:�������
�n�b�s�xmA#V�ی�X��X�XL���t@w�'P�<ם�x�K9���3����\%#�T�<N7F�;I�M�C�⮞х���m�qp����un�;��� �I3x����Vk4���K�9��cO!��a��v���e�1�m��	��EʈZBm�l��dCj�e�|x���	.��ْ� H8�6��cU/SL&�%Eb�S	t9�'Rb�ˡ0RUԑ���5T��zKo��v�r6JN�*#<��G�6��s���e3<K�N�JO�V�#5��i����O%���&��ӌC_q�'Q��:����i��Znfp��u;n1��F�<㏣O�)ޘI0u�V�ϒ�k{�*�����<y�z3���3C�O��(Y��㎞���i#1���y,M��{Sz�A����,����ͱ��:��.��m<�$�u�����Ə�|�u�^[�<��]|�μ��n�o<�Ki��4�N���~~�4��;
("{<y�������!�4d��2�b�S[�ggx����m��)����7�4�u�����\e�y3��N��)��|������詩b�S��Ӄ�X�q#�y��u�5�ǯK�����������)�H��f�q�|*v��e��-�R2	NF����0��%�B>qi����Lծ�KL�'�Ja�#M=�#]����I'�ڎ�$��}3X��[s����q�|뮼���ֵ�����-��RT�L5¦'u3I�? )�l��QA���d�dɦ�#;��T��6��GI)�����T}��?{醜IHRT�6�5���~�=�����"!�K�x�!�OӚ�.k�2T�
����&ͥ��Ö6ffl��٥D��fZˁ$����to:?Ѽ��e��s��״����/L5��S[�������GYӷnn�]n$���IK陗0�K���0�U�g��� ���Ç�Ͽ�Z�(Un?!$���e6�r9��z|��|����uԝI'u�YL���!ӥ:<:���y��QAI*R��W9X�1�z���mC)2|:)�|'I����A�g��5b٥�hnx��w���o��~���r4�f0u&�r94�MTLB)��QL��UW�����j���4�aq1�Rj�U�93�fp1|s.�T��j� �$��?p�:(��x�3Z����k��y����>��%�>�顔�=��f�����R�mE$��J�2�e�ƣg��y�6��κ뮤�I8����e��<e�<���z�����i5okl���L"4��2���q��r�Y�ҝ4:U��z�C�S����A�xȧ�`��mr��j��C����<�5s-A=�=��E�@Ć0�J8�mw՜�&�@n{�������ێ�r��}PD.�=Vc��c�4��)��ݪ�H%�'��O��4X�k���ֺ1�,{:��ZŨP��h):D�h:�ce!BWA�6�m�qk�2�l�;�ԧ�b**:�a,�JHے�=�98���N�<�	Ip&*1��T�5Zi���aϦk��$꣓9M�Zr2���aέ�-��t��߃O	U����I���)��Sϫ�5�R�g��n�^T��c����u0�̭�j*����aɌDJN�2��ү��2�Miyv�%���v������Z��SH˓�Re�Drar���Mk��J�����k�xm��L�}LMUZZ��Kq�mku�uԝI'u�YL�����;d�aFx(��-:o�:q�a�FR���*�5SX��`5m�ʜm�3��R&a�B�Q�w�:G�h��M���c�!8_s��y�C��~�O��}�DD7<�j)��~�0����X�Si�,¬��c�b[l�W�����MK�a�a'^a���������bi�Ż&<ʒyi�f��|�[0�-�X�MZZmN��o�[�[�8㮤�'u�YL����:t�OOO�Z��)^r��:�ǅ�����'�����^��I��p�{O�u�{�i�gU����υ�E��!F/*_��<�<:A!����A����-�k�8y�\ˢ�a�RBmZc���W����`^w�=3L��GsM|���a'�ja�O=�MUF�|�I�"��:��s���n=�_>�3���T�v�'��^�l>_�9���2�OL$�71o���KJcl���ǝ|��y�uמZ�yk[�[�<��i�)M4�������f1Z�e2JN��%�͹�T�jo��WϦvң�ˬ4�����)!��.��P���X�W8!��D�MT��Ă�L6Ca��0o�1ɕ1D��ss����K�|=>�)'��䝉�:�q���U0����UX��ʝ���JN"5*�13136�N��m�b�)�JRW%�|�F�c�M�;RO�R���0�۱z���9q%ECL;rfs����ۭ��\q�N��$�u�Y[M0�)��ӐĹ1ʨ��'�f'��g��&�y3V^d�D2G����v)��Et"�\��-l�bPC��L��l��"yJjc�ٱ[$읲K��A�{i��Y8Oi�qH4���Q����[�ϟ���1T	���I�k�6���:��Y�^���ܬ�tZ2,�Q��q��g�fS�-�dpn�$��g�8,�X$�Rr��c]��g�w<a�sH�Y�n��=��T"��LĮ4��]8�m�ՒRO�T4���H�l���&���������_���!�$'��>����ک���Up�T���5�f>\��<J�JJ���<���>�1�T�}3�#
I��>����1�*������M\c����÷
6��Rc)O�I^��U ��pP������J����t�x��0��|�n��:�I�\I$뮲�e�Ǆ:t�Hm/>Nr��p3�vE��3�]ܫ^+ʔKo�ӣ�Ñ;K�N����LS9O��URڎ,�a�2��<�	���+�D�	�Y�\�L�%�)6��7�M���a);E1g��U��QU�'�;ZgL�"q3JuN�#	�c/uL$��h�CGܦ#57S�XO	Z�D �Fl�i�@��^% �ψ�֚b��	$�\Ʀs�}�f&���i�q)RK�F^Xa�S
��^YI��Ӧ�i�wS<qƘ��d�m�ۍ��N��I�I'�&�I$i$�0�	0�i&V��R�Z�Zֶ�[�q��I$�I'̢I�M$���ORI$�L�I��6�q��>I&�I>D�z�)6�I8�ƘM0��0�L��e&I&�x�'�Ϟ>I$�I-l-m4�,��V�)K,��kaJZҵ����8��S�N��N��댢N$��Qee���ki��q�q�yם<uԒI8�$�$�4����-kKμ�0yy/%��V�����a��N�9�'�
|q`f8���?,=y�/y )#Rʥ��-��=����p��wٔ��=�MoF����H(��b9T�N�3�@�7� A���KA�p��}l7�#�Ţ Z؏�q�:I�I]bt®'�3�����GYi�	��0Ո�yRh��F�<!6�ɕA
k�`cg�t���d�D�$����q�[�C>��Z�x�w�w���]���;^w�ֵ�w�������y��Z�u��ګ�s��{�k8|���6ێ��u']qԒuך[M0�)�����I��);ED~k:�V)�.��K):�Cn�֜Ki>���Te��kb����}qȊIȄ���̜�4�m�
JI�{ߜ�i+)����B:�qf^2�L�lS�y������1� �B��N�7)��)mJIؕ%���f|���e�R}���&j�����+��-L�&b#O6��\�m�hz>�ey�d��.(��N�뭥Ǟ[�8�μ����u�ky�[M0�)���"�sRA��^3�&S$���٪�ދ�&�Y`(���������c�C�C�N��H!����o-�o�n���Ku�j�J06�L�
���ξ��q�J;7UU�,���"�YL�eϮf�>��k�<��Ң���a�0�K0��0��Wl�ʪ�)��x�Zj4��RS1�S���K�u?ffU�y^��cn%'��e�y��q��TTT&;��\��kM6�J2�X�	�ao�*0�4�֗ζ�n8�μ����u�ky�[M0�)���_q�
#Z�<��]�i�I|.9��g�O!q�;�X��Q�iy<��~;��e��#��#܂�m��� ���#Y�lt	 �}���U�oJ����_y0ߙ����a��Ǐ�o��g�x������t$ֻioC�hz1�Ԯ��rË�s�/���{|fz�"|���<)e6�[m/ã��h��)�;SII���T�Bd��M|���M�ɝ����m��m�K	E�b]�oX�-���3?jW����aJJKD_�UU4����jW��U��fv�IJ�����S�ZJN��rԚ���&��*�&�[����D��>!�>������f�rYK�%���)ޝM��;{7G�;�D��C,#�� ��8�_D�5�V#�E�����]|��q���張��<���im4��S�ٙ�j��EIZ�S)�RuӋ�ڵ�M$>u����F���R�O|�R���$�%���MF�V�eE�s�1/����x�p��f���kL�357*���ܯV%�uii'��8��|�p����>t�\V�$�,��mZ:]v���|��.R���eǓ���'�>a�������	��>w��Kl>��O:'�p�c��c��R����Z�9)Jsu��S4�m޴��|�Ϟu��>yo-o<��-ky��M)JSM.�h�����g���2<Q�)���ӧ�~���d���%Sʪ�����O��i&�GX�=�X[�i�c����:�?�����=?�!?��=k򖨦�n�������4c��v���hBi����4�_K-;��ʒ��T�����T���.8ʘa&�u�R�9��7B�yϹ��$��g�< {Ģ袔���)9�?s	�+ϒ�1�H!D�?�w1O���	����u8�n��u']q�RN���i�)Ji�}�Ϧ4���8�S(�����ۗ358�MR��S�����%p����a�ͩ��)�99y���x�}�m.2ʛ]qJ���Kj Fs-���P�r������ē�'���	gI�o>�ç7n���z�����W�g�ڣjb�K	%.�g����f�3�6�Y��\�S�9mԔ��np�zg̥��bg�8�zc��4j+*Lש4�mGˌ�i,Q)��ᚙ��i�K�6��|��|��yky�^yk[�<��iJR�i���fU*��&R̎FXX�
=��$�PT�T�h�[��N�+q��(tL<�%瓑<t嵵��sC��Xm��Qi%u�n�)�����#���$�m�g�s�~�ȼ~�iOn��5߾��1��.�:.�՜V�E,��-"a�(�qa�Hhw�֪+����H�u+�w��$�|8c�'?�:^�JZ�yl���&�s2������u�IKmj0Ӿ�e�<��:F�ʛ}S=Ƙ|��G�a.�.�'���0�Ÿ��2��*2JRԌm�F%�G�l��)Z[4ɽK��b�iϙ�5��EF�\J��-D���;�۟����.Pϋ��9#��ȃ/L2r�\($��J��D���3��v�r�%�V��"�ۘ��X��nW��1��iʜi�8��u�y張��<���[m4�)M4�J�2G��3��e3	J]�\K�*�,ks4�)pK��Me���*��J]L&"R�ձX�Ti�n�Uky�b���;鄺��>|�M���U�DJ��4��λ�>�\p{雍ęJR�z0�&c.·3��At�Ť�HXR
�f�H�l���`����(A����3>��;Ħ1��NQ<���!�~�m`b����o7�f��!��D	�4㌸�f#*R�Kَ��R�i��b<���Z�y���[�[�:��Z�y��JR��N�4�JL�����s�:r�c�ӣ���[#/�&=1�A2A7������#'����n0�R��ì:��'1�(S˟�3X�E�^CZRp�.H�=~�r��+�j��4�B#�0��"�(���*�s�q���f5ٚ�ͨ�)�S-6��"=1�S���WU\SN9I�7JIv>`�C:���R�#M�k�>��Q��K|ڞ[�q��<����u疵���m���!ӧ���|y��y��*r�9V`��^	�>r����di��>+�I$�y�Y�&-��)��fS;�C���2~o�1;'2r=Eqg^�BH1�����r����ࢌ��D��,�8�o���UO*���3E;1����R���=���3��Z��/Ge�q9�e5�cL6`�\��4�)J��<�8��?�K�"�`�a�=�h��:3��&[L���&��[n:���yi�I'	��$�I6�����z�M4�i�<I�-kuiq��Z�q�V��խ���RI��鉄����I$�i0�q�I6�$�&�O��I�m��m$�i��Dm��$�I8�$�$�M�I<x�OI$�I�L��,���JRҕ���l0��jZ�Z���<�*Y��%��e�2�8�oSL"O�a2��l���q�yמy�^y�I&I�I�i0�m+Rִ���e�#�%�a�<��-kqiq�#|�/U�n���;=����N+�W՘y�^�Bqc�A���E5����C%>'�Ϋ9(�q�;yt�H*�!��:٥M�\���B��E۳'�]su��=�R�������va,�����N���d�j0�(�N�pV�1�vn�1I6"���6Ɛ`��(�\��!�a���0��*i���!�m�f J�fq�N��zv]hb9�\���|�32@`�	=m�Ȥ& �Fra6`��.�7S�`�(���&�/V��#��a=�c"F�R-`�3ď1�Kq���s��f����	����x㸘�Ȇȍ̸�i�x�/`I���%�bQ��d�&H��.����m��F�mtu���)���&�J+`���v��KKeӁ��(���N�{�t��gt6T���
z}����uu4UC�a0�L�B�<[��T�2���+�0�Y��񻸿OwU4Dp��h��r�7nBnk�hڍ6I4��$�Q��p������%HK��˄(�X�J���i�š�rgkT]�h$�m�����s�l�6�mXag{�>w���i+t��`�
�Gs��y܄��v+��3�N ��\�{$h�^�n�|��`������H�N�$��\��b������~���\�:�3���w����W9λ��=�w��UV���]�s�Ye�^:�N6ۮ�����u疵���L�JSM����;VH;BB�1t�����?}qcֹ�.Փ��7N�un����8�S��vf��X�KvDV$��X�-.(�©�vU�ݷm�
d�e=t�ø�q\�Ku<q�ٶ��Ǎ��W�n76_:$y�n�(m��=���ט�sΔ��^�=s�� �c�m'�9M�}J�)l'n��)k�汮Β8x�T�v�Q��k�����9���1�=�tM����N�����t{��vx:i����X�d5��j���ny\��L�w�h{v�ef��v�����7��Ŧ��bɱ6�!F.E"�$Řo4�MK��*(�7��O���I_��u�>#N�%�GBg�A=$�%螒h��e^U���3�%��8�].P�K�Q#ʑX�EbKa�G�$�6͖��h�>���<>�0��Tz-L1���%�i�Q����R�ci6��t���x�����_m�\��`�\ϾUq����1o�SUR�55[u(�_���z6��fS1���U�:��a+�L���y��^�� +�+9�����>ԈDD�Im�6�E$&?��Y��6��ѝg:�d��^~>��|e�L��Wɚ*����wU[G�qO�|�\q��-��y�ky��*R��ч���RcM'�S5�rqx�!m�P^p�/׸|���O	Ώ�
nS�<��;�����M�i)H���L2���P���.i��ڙ��)�ĭ�b4�����(�.\��2���q��r��][�-�2�:b6�Υ�л��0�{�?��wn'��V{Vn���Kn�ñz�O~/��xa�|:"iip�p���c5�fw�ĸ���;LJuK0�`a��uX±��Um�%���M0��u�y�Z�yמZַ�[m2�)M:y���'�(A⼹,f��^	穈������뙮"���~a�e��>q�`��%����x�bX�k�A��>@?����`#���8;8$e)-I�XS�3��FB�h�|��u��|��S9)󑇙��Ħq�JZ���U'�:�����J�S��p҉K�-��M9��6��QY�Xu̵�?WӉ�Tc���qhӉ��ˌ�����Ͱ�ku�-��Z�yמyխ��L�JSMEM�q	�1f��xw���OϾI.��~|~,�q�V�%�c����-�,�s5S>��Х�i6���R����z!�Э�TvH�NX�&b;�q嶺��URU�	2��.�ɨ��e���3-"_S�9㑩�^n)��?MWR�y�y�?#�Ta:���;F�F���k8��S�u��QN�0ԧ/Gϕ%{��Q+�M����y�|�V�ky�^y強�[m2�!�7>}��5"�*��݂7���;<�ʜ�����7�oj���mL���; �U-�1��w~�;�q�h�vDz7d��=|��&�ݹ�y[�6��?~E�_:��2����9d���vnc���3~1KĴ(Rj�1tL2k9�fѥ��7Ԏln����~��4��%����T�l�_Ǒ�=�{��'= ��P�a��N�x�����,���0�0����1���fkmǦ�r�L1�眙�q�n9p�^a*{�SRfS���t| ��0<8��4J�w���Jխ��ɭ����.D��i�I�qU>f��k�j]��lu��/4�ڂ���B��l�~M��A}�C�
4��!�2�L�3�����uja��q�\u�Z�[�-�y������LB�N��dY�0� �bQ-�Tor�L�\��s��sUM�^�����7�dڨ���40�`c�S�4�3�5!~�|�I[^Iy��N���z�X��o/W��m���)QM�������g����1��(ɾ����T�C�-��HKlrfi�IGE���Ny��������E`����OE~��܂wG�Tq����!�=�{39m��+I��"^�O�;$zQm:ڝa�Xqպ�-պ��yמyo<��m�T�)�������q�<�U��s�~?��D��Z� �=�G�c����a�8=�vX�M�����;ҹ3��c����☎��v��ù�Uɬ��j�FNc]5>��~0_S���'\�#٩��rfx��n2�$�+NSL_�>�"�S*a�u��n0aĦ%�w	»(�*h�bk}N6�{i�Q���'ng��+1xM0K�U��}?v�5��y|��.��Gy�kJeL-�X[�:�-պ��yמyo<��m�T�)���T��W�>ֽ{�U�'
���z�ə�$�*L��ǌJs�늍�e�7�� 3���GF��z��g�r6ٕ��Ҷֳw�]�R���i��Xr)�
%��C=}�Θ���
�rb7T��*�9�Uq��m���L�m�窬�Ka��Չ��ʤ����)}�ۯ��WѶfdK�<��;���s�5�Sd����a�u�_%H�����!���<(���y��%�s�m�	0Ӌq�Ϟq�[�u��<��y�[L��)���.{�?�Sl5r��J�n+1�y
�L��rC��&&E��0��C�,Ë`QR�j@�v8�s��������?Uc��ˢ�l��P@�t�g�.9�u'���J�e�a$��~Ԡ�Jҗ��:Oc��'�Yufb�1Z�|
��7��`*��P�⤠�-��e�wq�;��#Bb	iXqV12�4�˩RaM<�#�LLc/O�7���3��*K���ò�q)	��P(���$i�𰕡��	��D���f��w3����rQ�'39�q�Mbt��2�;�g-:��`�B��7�!$f�Z�w��95
�Tku:r��%2�a�:�)vB��s����Gb�)��pP��ŗ'4x���JO���F��\f.�>�}U�g���%矏�q��8���]|�μ��y���e�)M4�W�+5S)�a�?>*��q�Ϋ��H �^�n��Xe��[o�2ˋ���q:b>��̟2�q�P����<+�R��/��)���#���F7��{�y������Ӧy�O�Ť+)�^+VN%��ZJ�bt�.�j]�e'��}?s��9�|_9����������`q3>������x�j[Jj"�"(Gyjf���-�a�jfeJq�0���O�e֜q��4�ORI$M��$�I��=D�z�M$�ӊZ��Zַ\m���.��I4�z�I=L���I$�$�M��'q�q8�I$�i2�$���KSk[�-kq��J�-��I4�O�I�I$�L$���I$�Iuiem4�L���JR�-kR�e�����Z���[0���%�^e�Zi�����m+-l�kR�Z��κ�q�y瓦uԙI=I�ORd�֕��V��iq���KE�/<�,��O<��ugc-�<��+ �G�=s z��B"RϦ��g`{o�j�^�g��[����o�WW�]��3玑]�\ٞZ6!�FZ�|c��w͞$�Ѥy���5��kܭl���"�SoK)Sy'K�B�g���͓0��j�)�qx������뀄	CW/hA�/�\ma��ӧ�h������Ӣ[���N�Js\"�I%�쌒/�D>	�&��-�@IRh�q��͵��7_��y�<�W��W9λ��=�w��UV���]�s����qUV���]�s�̲�<���<��<�<��yo4��aJSM�V�33$��M�:{��k��^0�g	�,��ĸ�����S���O˹_����
�|؛��L1�T�;��r����.p�d���؟�~��>�f�V�晍E�mbSқ�*�G��o/ԉ~␦���yĳ�7�:K��N���V+4��!]o�e��aP��=��f�+?&&�Կ��fza�r*0�J�vTی�y��q�[�uמyמyo<��[L��)�Oy�=$H�|%,����ϊ�%�˹�*~��h��ӱ�}L=i�FG�� ���K��:���%r$!�ӕ�����#%�K>E�>z{�-�9X0K1��nf�OL�r<qD����f9���b&8�2�0t�9wI\�P����B���I�-Ư�s3X��x���G��0����B#@���<[��ߧ2\���~np��ч���0�&Ҍ���:��8�-ź��<��<��u�t�!t�g��ו$ J[���II-�	4jR䘂A*ʐ;��Ŵ�7��T"�RB���s�w�:��nXfao1��U�rƹ|���e �{pc�b���V�*��n}�`��Dp���H�v_{��(��՚�M��:��*�"u��B��M��1�.1'^���]�?zBh[5CěEZ[|�|p{�`���Ɓ>[���v�f��s�q�ף�c�=)��ENf�Y��ܙÐ�'���*��Qܹ�\�\��#��*t��UV²��j:��3��cϓ��F�}m[��$�)�]��I�O����S
nO���u�W�Q�
e�|$�X��B�9
����r�m�
�k�gK�����������>�%$CB���4`Cã�s: ���C�@�0|[I�]���hn:�2��Y|�8��[��o:��-�y���
R�i�ǧ�(�s�����^(���@�y�%��TO�w��w��E����t#���*����`�J������`��SP�ѣ�@�F ���S�1��l���b�|���|�G�v'Q�S(��٨LK4�0R|}�٥��1�cW0Փ��Q�n�'^����e�����B���zM7�������氩�UR��l�Џ�^{���x}S��a1_��X���iy��l��qkqn�����<��q��,)Ji���e�LL�R�933$�">O~z6둛�qR�[u�/��tA;Ω����'�#S�C��<�"l�w�V�����ƜRI}��0�ƹ���N��q?��C9�5\q���j��l5-HB�酼��ءO��Q���6�{1S��:�.�L�3+JRS,��`����J����j49� >#� K��U�A����VN�X�'�>-��>�e��mkq��m��N8��:��[u���!ӧ��Y>���U���i��fk��0�D���/ѕ�����v[{�+��"[,cn�sw����UT�_'<p�H�������G���x	�ל�9��y~�걭�2^t(�"/Id����!2�'�Rn����ш�tӑ���ɺ�cX�kIm�K�f1G��ۙ�%�3���ˮ�*jX���5M�7�|u���Jmז�kin8�嶷]Z�y�[�6�Ki��4ӑ�f�Y�Ve�D5*��a-�DJ30�1q�D�e��ʸ�<x�ĸY�Q��w�zi^�n�<���e�a�ʡ�ö9����ϵ�"�!��72U-�u�UA�m��y���[�e�(�����c&��#���U���2�P���h��a��x��ʢ$Lq +b��'�5�cz�62RJ4#�b���%S�f�Yo
Jfϓ�Y4�OS�n^���1W��̴M���YǢ#�^ӧ��
^fs�����Ѹ�l=�Jw�MJ���ͼJ�c�N�R�-�ݧ�Yvw{��n)$�����zZ`�x�)�|������X�g4�����)8q��
�#|(�9��B�Ȩ~���ެ�زG��:�����,���:�<���[�y���<��e�)M4֙��?i�]�UA6��C�2O|
w�S�J�MF'v�]��a��E��Ҁi3��֖��>���|<%2��7 �W��W��|�1�N}��U35��>l���^fi.���]W�<~����B>��g���g��yMP��i!6���!U�	i��If;yȬ�;��C�s	��<��4�S��r�TE�w�L�t��-}3�b3>�8��R��}5V�L{ϙ|��Ϛy�|���[�Z�[�0�Ki��4�{;�bR��1<��̒�q�����GU	��U��';�����$�Ӭ��`*\9y�O�����g	�܇�����?c��xs�q|=���=�X�5Y�DRِ�a.�5Ӕg�ܜ�l�=��zP�@��A�Ʋ���-4mq�Ly����E�"��g�:4�����?Q�-?hȥg0n�ﴜ�|����G���4_�1(���˾O،4�P[�2�|�<���[�Z�y��Ki�!t���V<��8��ު��b�w8��I�9z�\�|����?���>��}p�1N �K		�f��ڷp�.u ����)�Î"��n0��z�X����6�m8aU�&ڄ��Iu>�щ�R0�OW��=��0��8��E:ʡ���L���4��OE��D�*4}=�����a���g,�6�qQ9������'��q���ֶ��$I"I$�i<L��OYI��i�I�Ēm:�8��iN�kin-jZ�ZI0�I=L$�I=N$�I&ͧq�iI$�I�M����Om��e4ÄD��I&ZI'�$�$�i$��z�$��L��|�2��_$�OZa�-m�l0�Z�akJ[Yka����u�[M<�^I6�D���&�O]q��6��<�ǔ��-k[�,���V�֗�K�J��\m����kJ��[KZ�yמ:�瓤"YKC�^���Q�.��0�L�����oU���ĈLN�K�w��I��*�� ���ˢGK�-��Qߥ��-X�b��/
��2�`��'��>��>��$���V��4�%��K��f���S���5n�Ƌ��옉 ��h�tኂ�Q�mïFɆ	�y[_����yW)���8�RDL��=tR:6Q����W���2۴ۇ���a��H|���a��E�#+e��T��D�Ҧ�������~N�� �#{�GS ��2�)IF��%T2Q"c�4Z?����)�UM�{���p"L�g5!e	�����~�]�v��������E�����3�(m�L�1��m2(�k��q�9��7n�c�f���_A^ce��M�����]�]="�{Ȟ%�X�jf��톨�v�yp��nّ�?���G��rf^^Kmql�iq�+۩�Z�kc1�W7&���\�G�΋{s�it��rQM[I�~��;����E��x޼^���@y���z�m/��}��J����u�4�/�u�x��(�:��3�@��hP����yܣ
=R?�d��.e��yz��J�q֫�yH1�yi%� `��h�	�������x�g�_��+�5���?���*�\�:�����;�����:����q�����s��9��,�뮦Sm��i8�M��N������B���=��O�&f�m֌y�X��Ѱ�br�B�ېlG6bde�~�L���'
��n;y��s��Cu��i��Rűҝ��t;��冨���-p[9�/M�7A;�����i�+��{q���U�kC�> ���!v�]H��\�l�Մ�����3P��
R,g�&Yu$�&)5IV���	���c���/�����%��E�9>��H7�ma�ek<�{T�v��n�2�;UY��%��E�M�\j�q)]�����m8�zѳ��=�t�r�+wm�w�ٹ�����xn�]� _+�N����B��ɪ�#�=����]oճF�Ӕ_
�'�҉,�LkX�Zd���ҫ �$�#�_`x@���nޏLEP�d"���)������|44t~baN�s�oXF��i�L̮-��CS����a|�&�a.ny��V%�7	�{�n1靺��վ�~וU����C�������<��#Q���V<�#��T�*nD��O:ۉO~Oϯ!��Yn�\��F�D�꿔�T�5��_�����|i��1�bd�92�Rf��uU��-4�ŭ�ێ8��[��n-kuo�K�-�XR��M�F�P�L�G��W̪�yχq��H4�=[�-�����SǕ��c�I��f�5��d��+ކ-1��&#�mܹ��f����g��'	��c�eE=�&{$���l*�*S)|y�!]�E�J��	�1����a�K�3��a:�Zf�S�q���>0ͷ�r�d�^^�SU�������F�/8㭸�[Kuխŭn���JK)S,���'�x�7���U��>��3���Yn?t�U|�)gH<�Tr�a1�z�&S;K�V[p˱%(�E��G��G�|H��$1H����7���QHN�˜�Q���G$�O�����P�Fm9�Λ��M4������Λ�$���_9�s�À�?T�|�+O<e���}�L�"7^�[�c�8m�ѸJ;	e���κێ8��[��n-kuo<��RYJ�e7M�Nj���r�s�32K����;��Ϯf�󑥭L0KQ�Ӕ�_`�t���߳C�0������Yj�+V�2�,�����C�����C��9Dy�+O�ӡOx<��D�F���n&:�_8�b_+������n����`�bh��y)�噽�\s���淲v���/�7O9���#ϼ��F�nx{�A
a1��'l-��qn�ێ8���]Z�Z���y/4���2��~ ���U��̅�_��Y�2���b�i6F���Y9�'c��5�b��q�R�����&L���u���E�4�2M��Frͭ�0ۣ��,V�,�Y/
�{ߞ*���1��ɪ'"*}:~3fb؋N{)�fb����S�u��^�����-���&�H\@��l0�r$ԧ�a��9�stafݭۻ�,<��aEH&	'�}�0`��j|�$��6��.2���#L#O95��Lw���3���bg1׾G�։TJ��Y�4���N�Y��<t��aM�f�i��I>�Ů0��s�g{�$���N|��^S�>��xc���N'�;��+�D2�2g[l�Rͥ��r�n.�v��v1��Hϯ�/!���L}�n�)q��+Ѩ�&S���e�]i�>qm���q�n8����ukqk[�y�Ғ�T�.\Re3>���33$��J��UNRC�ߟ��Mw#'�&���u<N��"R�W������~�<?�N 4s�.m'R�=KY�8�m蜳-9jf6��~��ߟύ���F�%�
c��,>P4m�QL��%:83��xN~2ˏ�pi�Cy�m�]r-1qڌL�������(�y��5^���V��2��,-���ϛq����mkZ�[��JK)S,��đ��6�VV9����Z���M�.LUM�ffIw�j�:�'lG7u:����)y����2|�>yq��Xi1�w�X��SiL�a�ILZ�>	���
7ԑ�ё|F8ݱ��H�%�C�7JR���}�*|)�&i��!������0�����;�#掱�R9Ķ�<D�^>�\�n�.�SˤO[7����mC���Z���ǳ0���>q���u�Zm��L�M$���_.<$�8���=ޢ��j=�.d�R�b�7-��TY�����m���������a���ü��Jt��*��֒�K�a���ʛ J�7�A�熇�.���3�����ݔ��U*�Q������A��y�z�Q=�m��B�� �0��熌c �o �����))s�hxlH��[MG���v�c�j9(z�3�|��ӫu�>q�ojf�����JaJ!桧Yi��[�8�[+uն��n��SIK)S,�S��+s�TǴ���*v��a7���I;iK|n�<.c	�.*���Qf+v鱆���|/W�ٷ[����mqM�#��H��hyn��L�-��\ˏ|UA<<~y�������w�k�F�W?v���D��^2��`ǩ��ޓ[%�جy�����,�q��LHS����\��'�)1�LE!a48�BJ����&�Ԓ�;��������c�צ��*�4�h�2�T��}t�/M���Tј�%��4�Gg|��a8�f1�Of0��.2��B~�5O2�$���G��cm��Lq�����&r�^�<�Q�P3�Aar�� ��iWDH&�M���<~]$��ވ����Y������	&)*f*xef]��e������+�k53ٙ��qӋ����Ϝy�qken��ֵ�ռ��i)e*e��قf��̒��!O�1���~��O�D�I��9��L����^�-�G#�[x�T�v�%C�����6��..)2��>a�N���$��:br�pK�L����Y2J�/�X����2B���$��E�H�W~��n�8�;k��J�G��x|�i/�P.~G���RD�gPD&(����^vZ�Q��1�JT[	v31���+,�)�4���D�s�Vqm8���:���I4�O$�m&�x�����4�m4��e���n8뮸��Kk[���H�$�ON&M�I$���e$�l'q�i8�I$�I�I�G�4�m��q���a'�$�$��e�I&RI�ׯRI>I$�I'̭��akJ�aK0Zҵ����6��������a+-iy�^i���%疷��-l-k[[�Kκ�8�n<��<�^a疵��V��kakiimkS�K�J��\m��E�+[em-k[k[�R{]MkU���X�H,�yl�E�����!|P'�sއ��tvA:�P'3���*|��p>�����@w�"Oֈ.#��k?���U���OH��F��2O�`��{�ln�Q�ɗ�k%	5���E.x���T�����!Ҏ��xg���kڅ�x�|_.vi,��-!�b,{P����gu��:��|y��ܞ���H[�=���?v��}�{��w���k9�{�������;�k9�{�������}�ֵ��i�u�qǖ��um�k[�[�%�����)��̒�^ :x��N7���@��8�p�(Q�S4���p��3�f~��S2������pj��(��&_4W���,��#�'���i��K�C�K�.���HK���!��H��'?pK
S	iێbp�,�sɚ�����M{�������6{�	x�Hy�4e�3Yj�̰�Ҕ��)O����9
�w�R?����$1�l�%�bڷ�}18{Ωm���ˏ�|델����um�k[�[�%�����+޽N��33&�{N�%-ߓ^�c����{���?��?��O'=E�P�s<�q,���<���d��<=��9�`�� ���)�����'�l�~���y>� �,Ɣ�����QS�i��◇GF����]P�˧�xOV�2�R���Y����j�0��h����0c�����cz<9	kd�Zyku�ێ-l��V�ֵ�ky䴔��Xe��}1w|>�D��K��2�Z��RA�6]��6_��|�ɖ��jhs�B�VБI'P�`%�
;�W'�v�8�.ۃ��&�>c�F��������ԲvS|ʨ#sW��h���iD������nvB�M��������I+[<�2$A!"R�N��i��]X]n��^Yk����'�/'vݦukH��E�K��n��ښ��������E�QXu��0L$K���?� �qsGy���g�?����"i��,o8o(b�}��.-���G'jp�^{�6>�a�r��m�٩���j��Mn&<����T�]�fgI��s�j�/�+m*3�&�������y�k9�+2ε��%<Ӯ�Ɓ��f����=��UF138_��e��[����en��ֵ�k[�%��蘦;���$#V �直1��r4�9��|N�D����i��uǹzt���������Z�d�R'х&2ʝ��κ�ݪUT�Z�pq���˩\eF��ե��X���eU��j���u/��mJ7����K�k_/ߚQ�]��v��mg�K���h��/uOu$�����!��}9���u��w}uLJg�L��Miq�L��1�'M[q�X�&��ff�mGL�/}��b�W���a�%��q�]y��q岷][kZֵ���R�Ya�_�)Cx�������?9��?���g��J�0y嶓O2���"m���M;?|�V'��\���\a�L���Ϧ�zS�҃?E�_��2l�qV気gM��B�������陙�=i�K�������믷���\��m�-98%�%.�|���Gb�/4�Ƣ9�r��Ov&s��F��M3���笠�1�����j;	�F����-��q�yl��V�ֵ�ky䴔��Xe���{�&"c).5��H��q�@�p�(A��z�?��O��z��ѝu]�mauv��, �5{����l��;{��R��M{����hB��Ҹ(���
:���Mm�)����c��Gϣ��/C����z1�^c��P~z'�b4��b�)����;�͖���]Q��N��i����Yo	��8�UX���e����G�Lƒ�����mk[�6�-����Z�Zַ�KiKIe�cM�^-�&����%Pr�T*��
Ne�ݞM�|$<6��0R�*I�8��۵�9��Hw�S7Iq���Ŋ9�U�;:Wn{v�K�L@��	��H�\ya��b1!Qް��Cco���b��/"��5kF�n�!l�)�EqцHKIbI�bh�L�0<0�)m���Iڇ�K*��L�.��Pg�i����L�QO��^�e/�L}ť¢[}�֍4�T���*��ó���Kn�pO�3a��L��|f#f�8��u:k��E�1�[�"��v��➙�����ǜ���ɨӏ2�ؤo{�fsI~O%y{��jw���y	���%�1U��&4T:��oȘm��Sm'��F&'e��a�|��[�8��an��ַV����R�Ya�u\�H��S�+$T�(E쌄y�F{UP�(���ߩ�N^.�A�'�r��� �D���G���?�M٤��>��g��;�6������<��'�Jk��2����2�LL�|��m��8y��h���}�p^�=h���$#/.>Q�+ɴwc3i�q�Ű�J���Jf<���G�3qkN�0}g�S_3�FSQL��r��7�Jb��V���hD򥹜ì�gm�yo8�-l-�V���ֵ��[JZK,2ے�Jfy����Et��a8����2rlnffd��\�4ӌ1����-���c�>�\e�m�mU�p�ZZg-�Ki�L唥�}3����|�M���#���.+�W��/ �����e ��f4�dE4��� �g8�H�4ʢ�.b��1���'�<��J��&��bn�y��ߜT�]��Ym�m*5��g�{�>���^9<MS��b��5Q�u�W�\}��)��O�ǟ8��q��an��ַV����m)i,�˷;��KĔ�����4��p���߶�g�O��r5D��l��NG\ӯρ;��G5��a!,,G�.e�~m�W)R�
���] �����A����4�L�9r�)�ǵ�'U[|%@4s�x~�8(#����/�?����ˊ��V�ܙ��=��b4�)W0�n�f��̰Ѭ&qa1W��&��)���R���E:ك	}�Xq�Ƿ���~���2�R��*�UVkf��q������?ѽ�?�e����t�>8�m�m� �-�_����~�n�m���X�=�s3��""ȑdDDYm�D�DE����"�",�,�"h����E���E�M��"�DMD�m""��D[DD�dB",�����4[DD"�"",��"E���E��h�Y�9����&�km4D[DE�DB!E����DE�MD�"Ț&���4X��4MDD���&�h��&D�dDMm���"Ț,��h�"�DM"$YD[kh�DDDYE��m4H���"�DDV�DE�""4&�km4H�DD�h��[[h��"ȄH�C�3�DM���"""�m""Ȉ���"&����4[D��E���mmD����+l�H�d&�-��"�&��"""-�"""Ȉ�-�""-��""D�h�4Ym�D����b&��E�H�,��"Ȉ�u�β",�h��4[D�f��D�h��DD�dKm"Ȉ��""-�"kmdYDD"ȑ�ȚD�d��,�-��-��$��h�H�$��$�e�H�H�,�"Y"�$�H��K$H��d�D�D�il�%�Y��$�$I"[I��M"D��%�i,�"D�I%��i%��D�I�4H�I"D[I"�m"D�d�%��,�[H��id��i&�$�,�H�[Y���iiY��M"Y&�-�H냫3��BY"D�D�5�%���$�H�D��$�,�"Yf�$�,�I4�4H�H�"[H�"�d�%�%�H��Y"Id��I,�%��D�Id��D�i��H��$�,��Ki�Id�$��3�h��%�[kh��KI��Zk-��$�ZI%��֒[KI-$��kD�$�K%�5��m&�,H�,I��H�K$�%��d��%��Y"D��k5��X��[I��ic����[Ki�D�H�K,�KiibD�ie���M&�H��4��m,Ki�"M,�H�[H�$I��i4����-�h��dZ"ZId��4�$�I$��k$�h��im&�,�-���D���9fq��	m$��KIf��%�K%��
DY5���,�D��%��E�K$K%�-���-&��D��h��--$��e��KI5���i"�$K,�M,�KH�-&�[�4��ii	ie�����3�&e�l��e�m��m��5�f['|���	m-�d:Xs�m��5�ٵ�f��l�[#e����X��ųhFhM��l�f��!��ɲ�d-�	�����&�LІ���d�B1	���,!f!m�Y�L!3M�� �h[8���9��h��D-��i���АPI��$-���-6Y6�i�I�֙��M#Z4�F�<���#$�4��M5��M4�HȚ�M5�D�kMD�FD֚&�Zi4��i5�$�kM&���h�2��k&����M5��k&�i��dMd�M&��F�i��d�D�M�4&���h�&�I�֚&�X��k#$�Md�5���5��4���R�p�I��i������M5�"ki�i4ɢkM[M�k&�kM[M&��M��D�5��5�M5��4��i�Bh�&��Mbi4F[M4�M[M&�k&��e��5��5�I�k&���M#[M[M[FI���i5�i5��4FX��ki�i��4Mbi��w�]5bh���4&�i���i���4M[Mm5��4�X�#"ki�ki�h��i����hMd�4M4��D��[FM4�X�&�i��ki�5�d�[M4�5�����5��2i���k&��&�4M	��&��h�d�ML��i��2[DE�,DDE��[LDB,��Ț"-D,r��#E����4X��4�Ț-�h�,�Y�h��DL[DE�B"-�"�DI�h�,���E�"Ɉ��Ȉ��DYbȚ&�!h�"[k""E�4[F�&���m�"m[iD�D��h�DYm�DZ$Z,�BF�7-��"�"E��dE��$Y	�dKb�mBE�dKm"E�"�#Z%��D�dH��Z--	m��Ј�"�-Ad%�D��"B���"B�,�F�8R�nBE���HZ�H�hDY$H���E�E����"B�DDZ"%��&��""�4M�DZD�""�"-��!dDZ$H�%�25�h�h�ő�5�D�B�E��B$YD�4�Y�����e����h���D�m�-�Ȉ��"",��,DE�dH��[DE�b$MD�[e��YE�"��DZ"-�""Ȉ�m�[D�dM�"�,���D�E�4Z""-�-��H��&�DE���L|�y��ǻ}x�ݭ��͜g���>��k�F6Z0̕6�[�s�e�����{����_o��W�Ϗ������������~�u�?�x���/]���;�����~w���q�������,���������}��>��>�3��>_�?����{����o�������8����~��c��s�c�?�����������G�߻!�6ߛ��o��g�o��&�~Oɏ�����q���o�����}{��߻��<?W�?s����fl/���G���(��n���:o��6Ͽ�&�_�7�;kku��Y���,�s?͞��wf��7?/>}=�/Q�Y�s�+y�����o��t�V�_��~篻��]�p������{��Y��������ٛ5���e�o����1�Y�mM�k[n�;s��8q�^~�9�7_��_÷��3��Ǐ�����}���nB@2��e	3Z���3P��6P�l�Q�.���_�?/Ѧ�g�{ߥ����L~�s��#���C�8"J��6���œ�?��������Xٛg幏\���~����o��������h�/��>��7��|�s�������~Ǒ�����[;o��?������������߻�濧��?��fl>���#_o�ڟ��s��N3�����韏��,}��6͇���cfl?����m�����i��q�C�vx����]}��{����^��,�[}��`7�����n��}���L���m�a�#GY�<����4y�}�Ms9�����~>[9�Ǎ�oٖ�u����m�:L�m����l͇0�o�ª�����>����o?�ٛ����g�,����}���������_��_��~������u��o��~�\�[~�����~���~Z��~������[���7�[�}���ٛ�6�pߛ��?��6��fl=��~O~�������7��g�?����>���ǽ�/����������h��?&�؋v�n���������Y7���&��p|�{w����?s�y���t�nۯ���yy3ag�_~�m��:w��3����c}���n���[��}��߷���������Y�LS�^]�6��Ƨ��_Ϟ����g�1m���������=!������s�O��� ~s��9���o�ͼ�W<��8ߡ�O�w���O��sc��m�/������rE8P��a}