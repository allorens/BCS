BZh91AY&SYh��Z�&߀`q���#� ?���bK9��    |                         }            ���U�P ����� � P$�)$)@���)$����I �J$��R 
��(%B {�R�AB֠��֪
*��	�I 	PQ5��  ��)U (��E PH PD� Q@����(U   ��T -D h�� 4��j��0M ���@�P hbP �P
� �Q@$\i@  �P�b���Rҙ@	R��Y@ Pa��i�dL((�E�@)1X ҀX3B��Di("XQJ��T� 
�URp  3�P�6U�4�PګUP�5��%@����E�w4��
U���PP�U�U.����e]΁J��@)$P�
U) ���  	�:������B��t��: 2�����s�4]�B��3��J�9��h(
Q�^��  q��T
]B� )B���
�p   v{�:��ʜ�
�Nh��*���@P�N��� sS��	��h� �N'sB�E�]Ô��AB�(	 (�%J�P�!�  ��:��)U<�wJB�G�*�UN/sJ
T�T��J�% sF�)[�P(R��l�k j�UM@@
E����  ��
-I�*�4`P�!��
U�aB��j�1B� ZSR�
4�
��hT1���TDU@ P��	R�\   ��@���IUY! ,��P�1S*�"�EU[Bj��I��B�3P��Q�@���EQ"�  �P
p  �%H�,����ԘU��2%��J�Kj��
h��UU��U@�h)U m�j� TP ���  8%B�j�Ab� +X
�M��*��iMIU �-�Q@L���E,
��V����}�   ��֨50T�P	�04ɓ	��T�1%*� �� � 	4=UO�F�%Q�4@  E?%%ID� �   �"�����'�$=C#C@��	��J��jT��    w����}-�튮�7�rի�҆�m�[��̭�^,�6�¬hيr��� 	!%G��
�� "
�UAQ[�I*����ՑY������ghZ!� 
���ڪ�P� TW�2�g���� �Ig���+�Ю0p`�į�^!|B��į�_� �_���� �+�B <H!�ā�@� x�<H>!O'�C��_��#>!|J������W�/�_�!|J���� � x�<J��<JD��!<B��� x�<@�%� �!|J���+�W�/�_>,@%|@B!|J��� x��#��/��	�D����(x�� x��#�G��� |@$|H�x�<H$�$��ā�@�x��.$O!�T�+�P� �� U<B�x��"��@S� �)�O*>%<J ���
	�USĀ� O�%G���"�� '�E��!|J(%E<Hx����UCĠ8�_�$Q8��"	�Ċ'�QO�$<B���P� ��B�@O �J�x�P� 	�T�'�PO��!E<B�x�P�"!�T�
>!�@����*>!Q�*/�|H�x�@�"/�Q|H�T$P<@�x�@�"�A�ď� |@��� x��#�Gď��!|@$��%|B%|B!|@!|H$��_�$q x�1x�<@�$��Cā� ��ď�_�" |@$|B����ď�OG�,�||FSX޳{�����K�b����%�O���7A��3N#E�M-p��+/�v�5eF.rInk�vKk/Ĵq��$�I�]�H;�ě�{�ے�d!�E�Mޓ�l��3k��F�pn��W@wl��î[�@�I׽����〹�%(�j��Pd�㏻�ŷ�\sӣ*���/i���rut`�;(�Y��7p��Ir�G&�'�_.�z��!�
r��&�];V���ާ�5�6gC3�S]ͫ�dTP�sᝓ%���[�Ï��B�Oq-Z��`���E�v����N�[��L���c�a�r#�[�Pv��B{�#��M�E�u�7wU'DE��0����\6��u����0☴q\�dê�n���jw�.�ǋ���a,;���˩�é��-}H'i�6j�@�pP>����rp� ����vtv�Ǎ'�dP��܃8�%덚�wnvZ,�-ٱ� �tt�3:�����9͜�8�f�Ev��(M88����٨�J`�9p�FЎ���
/�V󣓯��.��]��b���p����6v��&\��	kB�^��i5�tE��{�;�ͫ�'���0��rh�W�7]Y6P�I. f�c+[��E�	Y�j�d��ބ���L�X�n�(
#Q䒺�V��B���I�k�I_�ٳ�������lJ@(�E@�l즻��Ǳ�ldX����=��v�F��k�V]k˛&���͚��{����	�O[�*�o�݃r䷸�cc�
�o7�Z��7�샥j-�Մ_�%�.��<�Md���8�O�|::ecK�6-�wB]˫�J@xOw�JyYC36T�ϑ�s��{��Ԧ�s���Vn4�W��y:V\)g\��z�r'��ЍX�l|88ɏl5���mq��)v�[r��7���F������]���wd����U�g�ݧ~٧w�r"���6�v!�y��n&Aw��ӳo}%�X�r��Z��ַ:p����	2�o������3���nt|Ú�yH>�wm�Ж���V�5�7w2��WP��{:=�����������eu�uwtJ#��c����8��98A���R���.�ݦ�W���tΆO��v��*H-����v洕Q.>��'>��|!�l�����8b��q2�;��7���\}xL�H�uM��t��C��h����F��Tg,h敉<�����j�b�H����o._.�Z��,6�!73�l
��%n��=5������.drU����S��l���d��֜�ܘ�'&�� P���4Ζ��3��1���(�ٯ�"�գ�g�Rz�1���ڙC�7"<���kۯ�<��z��ۤ�D@�w�oq�Fi`�1{L�nH�2�#�7��F��Me���i'�h�OU�R�u�Zgv+���i�ҵ�#4�<���� ͧ���A��ΰq���N�r������`����C��w�l��tge��w�9�J�S����
q��5>�����2��4tV�� �#��Hq�V�Q��2"�5Ǌs˽�U�K������o&k�n���^j��C�wSaE��������{&����5� ��dy����\;�4������~���р�N�͛/k�X�ٜ2�:�_bܽ�^&��"�/s��t�i3�M��caL��ika,����]r����������b�NwIw�NM�~#�vVq�%��@��s5����7"#ӫ�0�]�v�/n�Uc���޷�e3fsΠ�n�ͤ�����DՉ隧=�v%�{7]�ѡ=�&��2O3AY�5��7��,����v�(Ҽ��*�a�;E0��3qT�����,�gc5�ud�=��F�;\%���Z�1,��m]L���фRk�7���mx����
'p���J�����b�����E�OoV�=U��E�����!F��0�f��0�|�jyO�▷���=��읋�c髎Ϣ�\�]ByǸ�����\���k�27�{3v\�T;��Svu�;��C��n���WOlFZ{[Zp��Vݫ=*��)�)�䥈�LTڠ�hE����W���d�<)���U�n0�,��y����e<.+&У��΢����Š.�  ��ws�Kh�%��HWŽ�yYyj;�YI
�ذF���E��{oCܲ�ey��*�N��.=��D�=G�y^�E��f�i�.#���U�a֖��;�	���'�� +&����_�Z��|���ʫ�É�vM��F���V�wH��$�>1��vvoa�r�� �J�3��I��ii�n�AӰ��q�h�3Q����!�o#� P�#�����Cm���/���Y�T;0e�K��T��U�*���6����%�Vvr6���٭q`7cu�;%�S����+���|5�������n5Xoww����8@ӽ�;���&�SzqX3M ��Ҵ�A�g ��m9�����!Ů���8`�+S&�x��D��W:��q����N^�xF��zm����/l�9t���"�!(�M��
0��4#C6A���'��T�G^f���8[�w�q"4��.���ļ]ӷ�G�BaC�ud���xK�,PK��!wL⇶kd}20�bҨ;�����B�8�::��	&ܺ��T��h��cJ�u��E�a@7��u3��K���i�#���1��5����jZt��ɵ�@�<oZ釞�#!����-�e�L�'Vh>��{78�:�:��Ȍ�
�f5f;��Rه�y�7��o�f*��7W��B�s�L܌�p�4�����r���yç�;۬I���z��ӌ��E�v�Љ;i���]@f���h�ol)gA��~�h;� �����ܗӗI�̋uYîX��ӈ�]�/Y���q�V���7i8�#�lyY��x�MŃ�&'`9ov�<���nU��{y�
F?����}����5�z�cc��g�&��6��'lY�!㦷f��gVr���Kh�w!��΅�n�`�]�wr[�;�{l�m���_��ut�:TpL]7ws��\�߷xqy��w�'nչ9u<�k7C��xֵ�dח4�PŪ�/|vYŭǞ0�w|d�DX�9�,<�g,�����s���<�94��}�n�'�F.A�|�O���!@���VN�C��`h�Lv��b��{Gخ��9�b��y0{w�씍+S�rv�&���-���B�6[�V5=����_Iӷ���Cf��tZ�ɡ��\�@���Q,L��P��|�'�J�i�׺#��Ν4�_a� 9� w�崺�Dod��uk2�繽s�icwΆ�;�ǓWB��{8�rZЀvkM�����v9ۜ�}�X8Ӂ뷛��#��F��h�³P�'+���`�ZC8Yds�ψ�.��m���ǒ<���+���,�9ͬ
������4��7yA�0�����v6q�Q��BZ�t]�P:sK�GX�x��v�Q$rt��<����c���p;��V.<ش��v��HH��jyľ��a��aUW�E۽;�r�;Wj�����7�̘x�%r-3E����]�a������=&�W@7w9]�`�Y��5��5.$�qB�s����ю3È��Onvı�w9t�<(�A|�l;8[NW�r]��� x�><�`^��H�d�I-:�^
���I�h�B�J���ǟ-@f��)b)������y(�[2s�����AU��SW@����A�ʨ1��LP4�ʞ��s��h���P���;��<�Y	^d��H;:�M-nvl\�'t�v�����w;p�G�����ְZ؟Y8d{�5��ϗ_��ÖM����*��ŝ��ֲ�\FA:���od7���T<5��x�eg5	�dF���uG�f�rB�3�h]%��u+np�t���(����Y�]}^�{p��vf��5_ �RD���!I�n��}Жw
ˮN�ӼZĺo]��r�9.0n����`�Ԟ�������ro���`���1W� %�
�gl�%�{��T��8�:q碛�D���|V��f��F�z��4l;�W�݁\"$	w����k�vb���30�(ۄ��݆j��p����v�8P}�`�la��@q��E��`��Fm�f�.jD��{��r���/2��y�5�8m�z6�t��w,;%{M�8S��q�3S	VB�x��NQ&�\ɤ!��Kxwi�MZ�<��3ȩ�c׽��>��A�{��pzfو����*�Ҹ��Wu���6^U��-���}���g��ˬxl�̭�Qb�c;�;�x8���%݊�95�K�]-��V��x7F�8�ꥪF���Úu�V+`Xՠ�ՇT]4Z®��6����L�]G� ���N��Ӭ�S����+`ܽr�9��r �Yw6���K�] �㚙㘍Wm;�"�*��Z���8SN�)�'e��rhgZ_21�[x4N���xuvhO;�fCg3{Bdسr΅Ep���bU��wT<z��ٸ�["��G�m���jl+�S�@+˖nR����#��J7�A(β �G�rH5�2Nն���YP��HƼ�~�ѯ�0���ܢ�[��f����\SA��iĠ��&@שR�a�̝z��ݺ^�n=�d�<(�pV+л�+u�=ױŻ��sEy��8�v͸1�Y��e���Y`�a���r��r�7+zO`��� 퍞l�=;*wf��	���s5�G�v: ��{2��)سC����2CT��>ѷ��PG,��gX;�[�Acyc��$_����D݅��I�9��VRMM�&m�4��j��l;7�fLxuQ�Y��q���.��.�����ts�d���)�q�[��8�`��1*�}��w�{&�B�|ӧof�a�v��܂ˏ-���o�p��4au?l��{F���t�;�'���Q��}�ع���	�tod�z���D1��b���#��y�$�$� ;'&���p1����x9����#X״�ً'Uûgm谠4������%Y�;��.�}���0C1��biW��@;���6�Z-A���_3�˴�
�#��mA����T�RR�n��p�����ȥڌY��s@�R�% ��a�Q5k�����3f!��X�:ֺ掤��Q�[����d��$�	O�����k�[vD���T�C�.<�t息zc˵�y���(g�H;b`m�I���7�-|�8��n>����E�ݰTf�����ݔ�U���v^fI���f�2d�5w!ß%��:��`k�7P�)e��V
�lag1��
�awU�;J7,�S�S�֥f)�XF����{K4�bz���q��ڜ.����f�Z�h���1�0-�M1�v�3���5����
8��Gj�3踜ї��҇A�qe5��"扷	�8��bЇ�wu%�x`�Q�&�:3�<	uk.9 vK��oh�nR����U#����_-���-��.9��]��q#����,#�;�L�ǜ�^�"�-z��$��ٶ5.th�&.����'�.�j�3���t�1�k睶-�J	�wt�f��F�j�$���~?k���ċ�ʖ��t��������5���u�%���Z�Sljǳ{g�P�3�'g<AE5ꃾ�o�`�gK͓�k���\�>
I#�/n�o*��V�4aY�c7����v[��,cP	E��ZA�9J�.·�����5���{/'���c�M�R\��*@?�	d�kǝv��Y�ԇ��e#����Q/�W{�':��t�)n6޽�������:88��v��I������k�V-x���k�ɝ+X���8D�=1�j�
�s��?�jm�c�{���PF���S�۹�S�,�nR� )� vnm�]�n����_V2�o�lH�Ś�8��;��z�%��;C��50�IH^5r���}{���Ԗ<��q��J/��,3v��!]9�^���݇�!��L�lɛ��{��1�ٖv���JJY&q�R�� 3{S���4䮷'���׷7�x��� HR���.�q�oTn>�i�P[2�wA+��d�1�\�j�͛0U5��9>���X��{��N�	�����v��<��o=L�s;�T���ṧ~��t�fw7Q�k�T�t́FΡ�s�k����) �8(�]���1m�p��ݲ�	U�z��n]n���C�:�'3���0tjμ;dlk�*��{|.� 8r�6��=F��Ă��ޙ�XۯOt�ܢ;Ռ"�^`gct��f�+��5��r��v��C�;���s�%��������#\ �ka(�Z�
(h����l�{R}x�	bR"v^�z�6���[��C	�۫�yx�MSv�KA%8=��uC���*�o�M�@���{�!ڈHҵ:���D�@��0@U�Zȱ0S��^����Ƀ���3'+�p`�4�7]�՗S�\ZCc���e�-���Q�l&����z6]��١eN�q}� �U2�Hہll'{f�GF��ܺ�Gu˥\�p�n�mR��1[C��� �*���B�ӆ5����3_$B�V���t^�,䳙p<�4!9\����nY�)W�f�³��k�2W({&sԆ�ݡu��H��nX����ƻ�8f<fj
R{^�;�5�'{N��� �:}.��{�g��~#��]0��o�p�t¯�_�����ތnۈwKo*j�hU`�CI�K�q6Da��Rr޹���YY��g^9�~��Ч��զ{�D:�Ս�"dˁz��g��<:\���!�	L�z����b�B^�4.[�$k�[U����[=���c����\��y�KVkT�}�������K��^IM��ܞõJ:�UJa�%�B�A��,�±��o���w�l����v�'�,�f��D�Q-�1�^�ca�5��;EEװ{�egN�Y������N
�:����rh_;�9�f�����ȼ~�s<�n2���}�t��.�`=�D�=�D����GܡG�GiǨ����2�K}%=��+�q�sϳ}醳I.���hɊ�N�Ҕu�S6�EV!z�BRU�]at���ɭ�Ϯ�⢘·�w�����OMg�0y��~/�g��W�s������U�
�.5\^��||�R��Bq"���^���\X}�x{�S眃���GN���`�S��;7�� �7�k��P�92�SO'���!�a9�
~]���:B���D��.�f��ND*(��m�8pVKn[��0n���=\�w�-e5P"+n����l�a�=>Fv��p�|aܪ�ݚLZ̲n	�bWY�N��$�r���3��'�΃���NM褝��=���ݓجzݴ,��V�#�^�qq�崤�n���P2o�؜�(w��X��^�����%�4�Xs�� ��$<.��B>��"C��7�@�����Ǉ�o�5�9RcV��)��y�3}^�\��5:���\��	�@'T~�pǸ	�鄯+Í�#��[�����iBFS+2+1f�6�5a�NKy ����1%ܰ�w��ш��I� ýn�݂�o@��٦)5�B�9�ۋx �{Y&��"{ӯ�LG�o�ov�ve�յ�䮓܁{_����{SD�&�4�����:Bނ����Q��ڛ�����{J�TN7yA�bqy��TG�X��뇒���W$�M͝摞"���g 0ӽ�~w�w̼��wå���t�d�r{�x=�U=G����Fz���(^=�����Y��瞋��P��R94�|Гr�ʫ��eH* ��y�$�U.U�XYs���?@74��욆84���f�)�7�[�Ѡw��Ge�띣e����no�lۂ^��-�z�,��|'H�����w
!�r�/�'
��㋓{�� �4AP����w��Y������	-�X�2,R�mh��\���Z��w��u��MIwQü��/L>Z��⼸��J+ԫR�A�WV]Uk�y������s��q�M�q�=eʈ���S�j�}�^$��=Ö���&�w&�y�u�V����Xd�zW�:3	W�b���3��ƛ�����}�{tY�}:��7>�x�0�1^|�5H
g�u�z�p#����5�D�@���֪1A�[�XQ�:����sb�r�:f�w}��"�$ɗF�>}<�?4��)���}��f:���OZ|Mf�>��{�����}��.�뮥����J:6��N�OH��+.�v�؞�;�gk�tdp�yp�ɀ.&6O���d�D�sf��է}�A�ź�z���ɐi���Z,�6~܂v6�^��M
k5Y�wd�[�5������}7Ǿ��3��X�b�Ѵl7z���z�b�Ȇ��W��7t�/�jɝ�Ho��>�����;���wwI�ϙ0��z2�����#�p�9�k&N���W��Ih��$qK}OdZ2�j%��F%�������h<qb	���pO�4W��^��/k]pq��+hg��nt�ݜq%�q@�Q[Ƒv��N����)�ß�����_,<!�S�_�{��dق�+w|Φ��.�^8|��c�z޲.ՍdZ��PH���l*ٙ��N/FV=f�Bv�;Z/��U��o���xH���Ȓ�#^xz��u͠���}����9��8
�X�hn���=821E{sپP����;��^�Q�ߵ�2X�nZ�Ģ\���/aP�����r���z�\�~�K&v�B�g/.��{�
��7�r�F�͑�0�ŤM#��Vn��3�ԓ��0	�5In�ce�E��=�{�_"yY��Ko_O����&=��:{��6Mr2��Y����X���3q2�9XTU�3�����}��9ڤ�˺8#ŕ��E|`����º'ɍ�G��'eC�M<��bC�DK����~��f~��pMn�Oof�Hoa��os	����5���j��:�'�'eX�U>c,B�=P�*���w�]m�w'����xT��o?�����u�L��Zީ��x6��3�V��V�����!E�����KWU(���˭�nu���↵B��;����}���Ƚ�ZGb 5�Dr�^{�=���Q�ٛ����0XmިZ�v�6��`ۚ���}��ND	��ְgY6g^M�Bc!���{m-8Nh�s����\>��o����#svd|C\��]�a{��Sv�MU����F������
w8�Յ�B�I'S&\��J,�nm�&�tY�3l���l�T2���d���m=AW��W�<Z�p�<D��ɺ{�=0��C��3[6�p֧^^���m�3�t��P^x�wq�5��n˨���zgv�U&y�(���.ѯws}=Y��_�1�u�4�v/a�t�Ϝ��ݧ�ͼC%͖xo��H�:x�~�	��q燘�I��t�C� \�^�������I3��\B���|f���e�)�m����ס�Nf��՗�}�X����f!~�hR7���<��Oϝ�w̕�2!ҢĬ����t{�a���G�s\�^=	���xvC�����M��ha��Ϥ
����^wz�	!��i�|�AyNK�:i}�7��`���W��2˚�2���9.�ηw��u�ڊN9���S�f��f
o�1��^�S��A���^����Z]W���� ���fF�2]]P��L��[�IU�X%vO?^G����ߓ���d`e�n�h�JG!�1�PҪ���fsK��n^�f��́�yh�VgC��7g���6hmo��u�t�x�n>�oz�^�w���e��D��q{���>�������(=�S��}|�$7�uH�o�&:-^Dw�)�!���8[񹑚��Gc�Lժ�i^/c��2��Qn5�L߽씶<�,���yҸ����<����gOy��=�]-N�@�gY�~7F�e�ko9�F���k�@���XqGWydw�E{�o�Qs���x?.��Jߖ-S}s�6S�[% �f�������l����[�h��!��V�E꺝��dV)lc��K���V_g�i�st����C�;�˿r��3����96mx0�]��p��ܧ;����UIPW������x]
=�p怕>\���+R��:-?.׸��;���L��{��j�#�6t>�a�h�/%Ƞ��v]~�>�ћ[[թ��� ���h6k����f̞ɚ���w;/�Qبd �X�{��h�=<�I�st�%�����׬�_�Ƈ�~>�=6y>�X��ǘ)[��Q>s���%��h�U��a�n�4B��%Ց��[��.0��+z�M�Zޮ��c\�\����`�6ہV�YU"���΍�cX���Z�k�=�ކ#OF�;��k�g�+nx�m�����o�z��G�{Q��%P�ɢԝ���g�,ov�4�x���PW�4��7�]��Ѽ�j��v.,�q�-��7M�&�L�S����Kȩ��UEۙ�Ǣ�B�Nv��<R�Z��q,K�zO//r���6"�Z�[��G��_C�B�zS1�l4��\��=��^�zU8��*0�'~��`��1aa�K��[-� ��f�V�d�Qv��߼3�q�ꏇi���g;�R�~θ�
Hc�=<�<�Z�7ܙ�F��&��CW5s
S�Uq)cװ���ӌ����LC̔Koy��]<��_��2����u���4f&�hYTZ��x��h7������r�|.paUȫvCwZSn�ڢ��x+.������&��@�&���j"�ڱ���gR�74q�9�ފK�<���$��?<�WT�i�� ��ۉ�һ�=���y��$����:��Swu<�B��\w����K����u�Z�d���B6|�����F�F�(\_9�nop͙3�n>e�IIo02��x��޻w��zC{{�j��(�s�)�zc��,�����{��Jbi@yqi����gT���p���Aw�y�.��-�z~+�-n���1��9g[�Vu���t-4�u�7CO��קa�v�tG���#L+-ь��1=3v��|�;�o.�t�Eᝓ�j�%(e��)Z[�YU�!��%�l"�㞋x�,O^k��j����>_��}�A������ܺ�a��Tn�o�Z��m3FP��T���">t��nI*� U�/�b�4"<��&�ϒg�Z l��D��S4����羶�R��(��5��7���OF�n����yt疼�{Z�s���臞�4z�R�[�q�z�S��NÓNw�y�Y�}����(��p]9�=���M	q��q�r��	��ѧ=��Ը��w{�y����]��X4 ��}�W�n��CVz�%��G*���)�$͡B*ф�c>	p��,T�f�!kTv_	���7!�򢞽��5�����xId� b>�� *YW������ý�w�R�U�n@�`�^�]u2�hI�R:�-�`�P��Z�[!�S0�6Br�����-M^���×'/LkS[ݵ�E�(?9p������Y��7w�̣F����s��n��̇	N�v��a[y�!�f�
�0)�L��Ý=��+6��@#��)#؏wj½�C��8�pz^����1��e:����پ����oL��+شA�4^=����Q�!|jXԻ�`�c��t)�͗F������Õ#>�̬k����3�����Y��'g�&����)A�9��@ׂ[S�SV�El*n*��5�z�=����I��;�e��/����ZXw�|�u����i��?x�,;�"�r~2ݞƹ����ޏ�Z�m̶�m���@/vї��޲G����ь�LKJz�pY�|��x���.�i�>���e�&y�����_��9�\�@�Ç���(Np�fŃݷ����m7�Ϯ&��ݯp�o˷��W�{����=t �<��"�x;$`ƻ�S����>�@����V�(jQ�x|�v�o���v�g4���*�gS���;9FՇ�a�2t� ɛ��%��ˀi Ml�-�.3`y�4��\�Q"ejIjѱP�ȕ�b��N*I2D\T-9d��5��Js�0섛�Ln7�[�}�f{N��GuO���y�7��q�����}���a�(`H�f��x�[8�Q�\�]<7�"9`��I������s����vJ��M�>�i��M�xv��Bt>�A��׳������:��a�kܳ��X�@��n�K�R|���Wfv�W��g��Q76'L����@vJ��gp�㋞�.𙤚�g"�H7T#I����gd��?v�ɼϑ�������f���Yax�Ӧ���")�KTܘ�j�}vM�I�J����y:C�r��љR�6��3�՟{v�s%��c"vx�z��Q��=���G�QE���ޑ���r����%({�׵m�o��*f��=�/�/iHL�b=��-��['�I����K���t;����v�ՠ/tc�@�6�W�pr�ބz9�Og����q����ǉ���+���_<�����Vd����l}}g��M��3�8�MI��k4�����<b�S��oͽt���K�n���vv����]<�A�8�d�9�ӣ̂�Dy�oo���.{�Y9/gA&�V�|���^~sr�Tq﫵�n{��`�ʕ��$!S
!Y�A(��.��ki���a=\��s�s̕�m��pȞ�{Qq6�܁Y6�6�P/@&J=��2��6b��z�ݻv�~tf�b�6�7�ɘ�.��ޫ�2���p����ɼ������g�۔�b^c��Z�UO� l;�n�UE2�*6��j�ו
���e:��W�A4ҧ�wo��j�e9�v ���R-�"���çX�����icc���[�#7d��4�R��
Uѡ���N�G������{���`��Q��ԋ,a�?�O���N�׮�����������w�_-�ئ��٬g6_�B%J�&Y٭͘�Tݫ�9N�$����zl6�r��_g��`e]�g!�$�M���o/"�K��:K�7�\��#��
x�����S�U��{o�f�ǋ�tOg�mD�.K}畮�{N.��q�kW��W��w��㍀�~\�g��$��P[uH⼋������M´�jw���{.�
y'3���GPoWh3��I/��{ۀ��OqS��vb�
I�Ϙ&��i�i�1�� ^'Q(��ƋkL
$�z�ӽ���Ŝ�{�.�.:�<$�p�x+�)}��e݃�����$D����q"����]��S���T;�ﱷ��x�rx�O]ޖ���*l�Í�[o�+�U;�ܭ���b#D^,�І^KV��x�����iʺ��b2�>7�1��qΜ6�_T*�O�kYmyx�N;!�f[�9J�C�U�+Zs&���Ic/V��,e��"��5��5@�
R�E�d3,u�s�h�:[I�<�A��n�LTn&��o0�so&�U��I2e���}���b@8d��Ndp@�y�=�w�8��m�R���0MQ�}My�k���!����a���G��V�:L��(�(����aMf���i��8#)`(�$�&�4���
���# 2�K������yÐ�$B�8����a�'������왐Ao��D^�3�FG�	���֏��G
8QOA��#�h�Mzqr��8]���qʹ�1@�/����Jd��*-���������_�擄�$%�����}�>�/��Z�[����Ζ{����K^xz��;�m�i6>��*��>U�����y{ŷ�����|��"�}d�7����V��"�^FQ��F6�{U�7���w�^�2a��j��/]���XTo%:t؍�T�З�[��8f�����sJ;y�C��v����ΔƟl�Qڛ�d�`皾��a��� e�`�ڟbʆ�����5!�18���J==���o���3�u��է�3e�����#zNB����o��p U|tj��,�SH���NʴS��
��SAR9L����w2��Hk%�%�	d{���v�y`���n���3�8geL^�vjF�5SKkc*��n�m<Փf����S�X|_-η�(��x�V
��K��;Hb���
H�2a Ǽ��A�+���+��I/��v��0�e��>G�z�E�'��VZn+Kl�`ZZFs�jF)���I|�S�	�{��J%����t��1wa%.�w�`���綝�e'`�C6&s��B`w�w��o�k�{�=<�#���XD��5KF��~��ޙ2�&�sjЦ1�F�^kPZB�K��-����b�fj�һ)\;�tGt���C'�����Uy���'F�}��Tﹻ壮%�˵^�q\�vح~�ʭ��8�í��ri 9n�/�}܀�z,]������ha�,0�1��0�h�!2�(��B�0Ba�0�0�0�a�`��QzF��Q;���A��#��O=��tg ��Z�i%��(2�֤nS�X�R���=���5��gv��S���bDh�9]`k��Cv,:;6;e��2w���gp�*��jۯGM��F�o��nw�t]�[gl�ܣ�4��P�nU��^�;��݅{Ӝ٩�a�&;���6ݗ���4��ḽ�L�k�2n��g92g����u��C�6e>�'��y�Fyߢ蟗��h?FA#�I��Qys������&EAh����j�R�qV��v�ܺ����׮��"�Y۲����p9�WZ�� �JbK*��[o�]aC�oww�7������E������L��i�\𛮞1��tg[��v�f�x�)xS;d�������v����/��o�~�D_g�]�����~�wE�����ƅp.�cƮ������C�H�����o!�w�s��[�9�4�zږzas���{�<���f��'�aW�rt���VR�Paj��Bː\�H�����6��D�u�t�0Q��A�{u,����@1�f {�pـq��e��lT]G<xsו����^�j�{ݝ��;0Eѝ�X��N�˞95&Q@7���
�<���$���M4����U�@���~1���=�k�.�<�|�3�_ose�x�}��9��Tn�����TE��� Z�蠃Їa�`0�0�0�2!
!�%`�!B�X�0�0�0�b"N�oY��4FB넎��S�H�|˴�y�}^�;{�C�NA�m���;��k%��T����, �ٴ�/yv�joY���A��(�N��w`�Ռei����mW�9���X�y7ye�h��p��m��9w��YV�sըwl,q7�O{��/yn�Z��®-Ȗ�}�HU�ѝ��8ӕ-*�9g���a�:���7���ㅤ�2��%�q�j�֔��2��F�=��/\e��m���٬v�u�}W�a��g�>��k��>�/��#�>J?g�������u�YV���č��<̗mT�欣�!%�!Ua�L�� O�P��֯W�K���X��l�2!C�6��B$)�8��.v���u���������f���Uo)t]��-Lyװ��_l}�/����r�w����͋���<�`�gg��IS}�3ڇb�7UI�ܞ�:,]��e���;w^��>bn�|�Fe�8AUf��Q��9�{GcbSڐ2�;o�l�PSŌ	���C^>�g���wZ.I�'I)ػz�LfJJHȡ����_�v�xjݢ s�^5��1xŞ;&����[KQQ��%˸�vj�G��<1� žK/5��=y��׆n0��j���qNAj'Ç/}U.��m��܎̋ؐ�t��:�9!�����LNl@oS���P�=�����w�̜�}�&�C�<�|]��#���J�*"	1t������8*$���4H��0�0�0�a���2��(�B�!B�0��0�
Ba	���_h��;��{��2���ƯM��=^N���C��2�Jn�L�͌[Y	Ԫ�-�.n���CQ<�6{/�MW�f`�e��`�+5璉}�S+'g���1��5�����s*�V2 D:�jVf�2b�m���D0�v~��ؖI��yJ�7:q��
��Z��7�;gsx��������S�N�[4/.�{�����qM���x�X�� )��=�Ä���5�ڹ�����<��{d3��'f��srע��tbz'�B�'8]����5����wT��Ei��+�����=98ɷ��kb�v�e��56sJ�w��=�%ğ�ǅ<�=���'�o����p��$ ;��O�^c�g��=ė��㕚���'yv��^��/��B��O>f_w]�"�����#g��Id� �k7���vvLE���Ĕ�(YX�k��QJ���2lmkC);h�n	��FEx?x�/ޏI�^��|�ש��F1g�1���4����Y1D7�4{�r�Nc�(ʸ��eЫo�ڇv����bci
�V�貰<Α@g���xSл궿?*�-^+Zkٺ�Y��%�*w`;}���u�ݚsZ{�ۛ��]W������5z;�{���B�i�c$�w��Q���3j^c�Û��'鐻����H��܊bN͞�}F�ݔ��绣׻��1�qc��-�",��f�me>X'n��Ge�b�^���C&!c��bA��*Tg\�'ؒ0HЁ@!�a�A�b�!��!B�(��!B0�0�0�1����0�ǣCs|�ـw.}�b��b8²��7i�
4�fg��&��m��>�s84���V��r~�}W{�=6s�i\aE
ǯ��qC�2�W��nh[����*���7�I����N.QN#.�9>Zb�X�YJ������y<x�爖���>����1����ϔ�))�4�&I�=��t�k��䅩�|0$/Qn�:���oDY����l!����I{O��Q�^7�����|8���/�i�d�k?kO��y(��d��q���57��YI'� �ͼ���*�Ԛ>�}M��9��Zd��{��U���|eV���\���4n�5���ӕ���{�q!�	�ٖ�w�^��נ�/G�\��z�%�U������}���>#������Y��9��&�R�����o�||���bQS��= Q��{����Z5�/^����ztj���ۭ�;{��.���>,v�{�gs4�"��5nk��]�{}_z�{�D��C���K�|��ʎo�f���C6R+43�6�ۙw���;���� �Z���������RT���������лx*�Y�M���O.-6�¿O��ȃA��כ�K��#=5b�v7�]�Fxo�}&y�/\>�-��yx�rHLŽc�{�y{w�<њ��L�vj�0%����{W�V��j�����]n=a�5[w�E�*!Sp�-��zp(O@ǳǝ�uM��m�s{=�lZ�>S`�c�h��͚�wj/s�_P7���S�#�E'<�ig����6V����J95	T"��S�c��3~��D1�j�{�c���l\rk�����w>x���.½��E��s^���=܀��AV{��<�u����8�?{`d�Z���:y83h!) �-ۋ��0j�pT�mؚٰ����#���6S�2�ܽQC�ޟ?������$%I��6��G	B�Ѧ!}�za�Ƕ�>���rՀ��.9���q �*������
f欧@�t'��m��h�2u)���[�7���n����f���S
X-���gzv>��,æpuo�xqҗxA�[��f�\�����ˮ\�;޵WB�����$Ӝz���#53��CN��Wx�o�<��z���{�(�¢�B��ݎ�����[�����7�B"ˋ��Y*�Gj2�3���Ct n��i�cB�2�TL�ڇp�з���2���h(��v��}�u"0-���t=����c���\�o��n����C{����g���g�.�<^�}1��ueG�^�Q���i��Z�o�g���7�F;ʵ˧������'�^�yC�-wz?aC:�y ��4Ěl?��u��N���d�gS�?fڇ�u��m�N������ѣ�tta�c�k���;�^N�!�`Da�mc�;�e�LdbZem��&���M\�*R�AY�G�,��oE��C���
"��P�KP����{�N
Xf�]M���?��S�ۉ\M�V�Ө\��,��2 �j��!�Pћb ����J���rT�Ù�:w������
Ɵ�E�(��R� .v�V�,��N���%�S|��|T������-��q��'�wo�ޠF t��;� �O�c���"}\3Q�z���:�}=ٷ��o*�C;�@���7O�>́AZ��r%�q�<1zU�{�r�|3��ɑgr�s#��|..l�M7}w1d�	}5�-1�^�dXPn�v�J�d�lX�o�Riī���t���o^��}��VI��;����j����)7�zZ:�1gf6؈Fk���+�J���F]xPC�t�b0���imN���+EQ��E��)3gL��N��sw"g�==�G��db�`D��A/��/
��w@������^$���N�"����-$�"7"��T�Û�͍�zl8!9e6�p~7���� �����}��w��Mň0�u����i�[�B2�;;4.~l�{R��B�N)��QAH��[���	�
n���qJ�11���T���u-�	����OS�,��n6ُvMK�$�}�R��9?�_���<��>|������|=���5��{�t�8�p[�=#�ܳ���5Y��=����}�|��Yٷ6�}�!�������oN>��ˈA^z�)R�\'3J��c�a���
�(�:?6Z'��]��y�Sy.�>�HW��Y���g�6f��|�*����H��y���yU��3����h�m4q*2�-�XU;�5��)��
�����D�_$b]����\�t�����������ǒ�pwi�}�9��5�d:>8���g�$~W�w:���̌�Ȭ17��m�d���&�e_	}��D��m8x|��-K�R�t@�^�q3�wkna{ѧ�^�}˫۲z�2����[�8�p�jx�8�[���|�&m~��p�G yȣalOݳ=fA�n�;�0���\3��<�;�����U�8>��&�,ܳ.p��l|��zKئ�P6�޵��^��˽�g<�3��ھ+�˷;�v�lн5�|���g��证�v��κ{��.j�����:9��# ��;���~\�&�k|����u=�V0m`����d��]	"/b�]-z����M�=٣��g(���MG��I^����&/e�IVb��O%Y�F�ΐ_�c�F�q�⏕��{:ؽ���OQ��Jެ����־1#�Rt�<�0���O��SY�y -���ƃ��!C����`k��0�f����P�{L�,�quX2d����sa�(���F�E˗�1�uͩ�8;{|V�H��X��Q�Z�4@��ۑ{�,�5*'�ےx��EuRǦ�zlN�!ǚ�A޺#���\��L.����4�8W+�c7�=���P�m�iZw=p��z{���a�T�$�W�J�3v�_��s/&�w�§��z�0�с{p�Q��a�5��E��-Xu̟o����Fon��4U[��X������'�'w�H�
�^۰�8��O&8}��� ����;�eѲ�k�=�)(���R��l�	�� ���P��8=�y1s���U��{��0f��$�EꝆhAЪ�wE[��Ɂ)I�@6��ԝ�q�ۻy��b��d�1"͊e�]z���X���]���,w����ֶe%NÞ�T�0������Xa1�����XË����?B��7��{p��ĝ�O��㓞���=&Q!Dy2��{=,3͇�XP��9o���2���c[ؕ�1ݡ�.�9�r>�]l�<���G�0^3�K�b�Gӻk�{�y�[嚈-O:y��L��s�T��N��8*[�P�9ա,�e�5�tVJ�Z�%�\��Rv�!�
ZAV�#�ʍ��ج��r�sf�Y���zm�Ú�;��@ �f3�|���i7̵�TɈ��{nәJ\�r��q�J̧�e��f�J=%��v(a̒��{#F(���)����q%��z�j+8� ��dm��~qn(�:�r��J��;7} Z��֓��2w�\�n���G���B�|��� ʾ'9��m��g�>�6�9��!�9�b�����=U�S����z����y<o@C��L�)����h��~�܅-�')���ujٗSI�8��1��罾w`ޤH����C̶���ߐ�Ku�uy�z�C�`�w��@K��l<R������㠶�����2nL�6?�s��S��w&��.�9z�>'�RԽ<���g�s}�.8}��E�y����q���"M�þM{��N!�L�e���`�[��%�݃/�;�q�����$�<#�	l้���D�$}�ޣ*��T	6��-(nr���j�*��v��Í^��agx�_�"�g��_�����{c�Z��L�@�N4I���"����v��S�T�%�T�Z�=���k��3���R	�C�[�����>o��w��a�>`!Ⱦ���""������4�٦	y5%���a$�,���n�%�	���eN�{՗;���=���>/�s4�k����I��x,=��~^?���=�x~�tw>�ǘ�]�����x,�z�i-0YyVS���九52r	���#&��Eڍ��o�4��3R�ܵV4�s�#�I$$$��������������{F��ힽ���y-y��b��u-��aн��P��0�����Z(��:���E5�j�yR����=�=�u.�@W4�/n���6��L��J+݂	=뻞�f!��F���b���tw�4�m���x�䚌t؟�B����ie�
�UNJ*��?��zh>���u����o	�J��èL�5hov���L�[(����ʧ6���^Ȉ �b����*v��j�ND=��L�m=Q���\�Q�x�ٵ�i����'tN�$$��o�j���ig����WSs�+G�2S+"�S*S*�Q����g�0`��\;ґ�S�kLN�/N��|M�Ҟ��s�;�.��H7t'�մ�p���p���<*�CC�<���M[�(>�� �{Ј���f]]��]�@/\gv��g���O�zk6_N��^;���R�;����c�0�/���gxw�Q��#��wٵ��{�&�on�6����I�0 �]Im�]��:}�3��@�ٹ8x�_��y�@�Օ�y)�u=���7k�@9{7`�1���g���%��:��2x����}�M�,�k<���&i���F�mY�w�ެ��YO�cp�>���NƧ��{�D��'wUw��X��������Go7a��iIr�sm��]=�Z�QN5���"ɰl�n���?�{о�nY�{�����X�/2>�@�@	`8�8�)�	����v��34M2D�~mcъ�m4�)���X��l浊
(��c���>>>�آi��cV��Ӣ+X�[;�t��3�[6�3mAln�51�T}���c��h����ꪛb-AZ�`�֚$�bJcF1�������DD[a�J5���[f����ӵ�Ɲ��Vq��LlX5%m�* �?1Q$}�D��`��6δSQX��cS��ڜ�QNŝ6ƨ��v�PSkMDV��Z6�TDŶ
a�LI%EQ1A�X���52Emm:�A�D[i�(+l4SSV�1lq��i�Q-��)���E4�m�*&4m�LQ4�٪�h���QUlf��u�ִ�Q� ����U0E� �֪։�#��EE6�&ݍ�[f �*"��n���&ǻQu��6zMwe����Ç;���0�~��}�p���e�`vs�+�A��^�O�Lt����uɫ���}��V�=��x�	�^w�����<A	8H�1�n������b����|l��Xi����Q`����f�C���]-��M�ݾ|���"�{��4�p�+�����r9��oo'����<��i�ڗN��Gpgg��6�@r=�G0ѱ�|8�.I�{�;���V�j�բݜ�{.��l
$L>h�vۆm�{6	7�x$�Ù���
��r�����0J�b7'l���[�Vöb��z\LE;q��.6J��y��]#����S\\�[�`\�ᰇ-WΑUU�7��Z��'8^R���S=�_c��t�:�Hf@R qyv�+�ݣ���6t��k5�-���n���[/l��lg%Ղ�+���	�Ġ��w�n���\��\ڒUȂ3���`ݕ�+y�WMr�n��e���_��&{#RǕ���t�h�������Z[����ɛ�V�談��hy8F�+7u������嫘^�tرq]���;� �C��O/3�c;?�rg��:J�k�S���lW�\�[����]HjȺXP�ZɯMc=��﷐��˷f-^��f!��1�Κe�r�ón!-�,`�1�n\���<�)�tֻ|�����q@�t&���+ ����fnr��a�s�YoV�/T��w��E��,�*� At&�7�=�2L��V{�y:@����f���G9�"���0mD��w��f��v�QT�7�L�ҕ�+�š�D�	Z��c��_aο�dѨ9�s&D����w�ɤ7X����yw]�.��<:�v��b��l��ј�:/5��&w��E�0s�u����_Q�Z,��!�;��A��":�S|��]F^ň�&��M��{�{g���䣇I���kc-�n	���[�E�����}�'v�GU�M�����-�5
��@�s�4w3M�UV�^u��k�g��5O���s:�HrF97%�c	&�V�.�z:���]ܡ�>�6�V�<�F��G1V���[�ݹ�2�HvFGҨܑ���^l哆V��#���F�X���3q��g��܋@��:g���y�*��������hS���%�S��������?P'~%==(�9��\��aa�j�O2f��T��Y�1lV4a"7kY��t1��i�)��N>RD7����˥/�\�_K���w\�qb]��5p�@*�q����^�G���͍�=V�*��v���
c2�<���m��ꁝ8�*�Ӱ��c�v��a]�f�X�u�[��l��۝�[oo�I��h�)���PZu� Df�A̷�-�m�n��ɉL�����.Q`ЬB����	:�F^Ȓ7*&��w�Į��g��=LzMq~8$���]��N�p�t�T�*-�^�Y�M_<��Ԅ�g\�p-�A�4��j�\��8��1{4�k���W8Jby��^�z���e6,��k�|HЁ�ȱ�5��;ԗ,��o���q#B�.�����[����j�ov��]y|i.�=� �i6�y{"��Ha�,w&"��Z������~�ϳ�B��X���D����QIgK:eTj��ɶP�l���9��yJ�h���X�,�?d�ǷL9=)��+��`��j���u���VG������~KU#�$?�A��
�P�ڧ��C%tC��b��P������j@� ���O���ݱ����9�ϴ]��![�%�7�w:8����-�$οt7����&���+��͉�݊��Mv��s�[m��2�H�"x��b#l��k��O%�����{!�]��'Nf�LjKp���a��+\�]܄>}�M��|;�m'�/����}ŧ��J��x��8m},r���l�[ޚ������,�bQI��3->+�Yu��z�6��P�p��J��e���z��6����d�OzP�ĥsǱ���n�35�~[P4�U��A����A}��NM�O���X���3���v���Oݘ��'��\���e�ySav�g.S����{;��x���sv<
�x!�85\��̺��9w�A��Y��͇��Uɞ�㕜lV���j�Sݺ��qQ֍<lNsc"���V��|E@���6.���r�"a�D�댡�V��k�t�^uU���q��Z)O� ���c,d!b�t��I���V��R�+2�^Qܛ�O ��;c�K�yS��B8��2t���nI���c,ظ����V�8^�ӭЉﲢUQ\8A�;�H*뿆�lf0��yQ��_!+�}���x"1X9
�D�u_5Д/�*�ݿ$'w8L�>1]��Y&�u��U��4�Xt��z3�ܐ�!|�����};���7E^�H��UW=Xc�7��'Cύ�dpCi��u���e��8�Iv����L̙7]��\Z���Z�����-p��o��@���r��n�	����8Mk:����B+�S�3���]��%v�u���
�s$Y����e.�M���9�\6�`$O�(@�;�����^�O��*,���3\�ď:4C8�On�ge^lH����m��,r�`���U�т�ԙ��(ۼ�%��Ov�}�.�����nN�2(9��'�_��v�W,���{u�� ]=���n�n{���wϷ�6��.U�ջ��%\�	a/�'a���p&�LN��r��#��f�M1W�<�=^zT_�s9y�g"� ���*�-}�g��t�j���i��8��P���iK���jch���S��qtȘ71�n�'X���lR;*,Z��9�۰��V	;�V6٬�!�pD�^�e�d�;\m�2�����叛�ӡ.�f}1"��Gy�7���A����<w���S�7��V_%c�����R�R*\���[�On�@�8�7g�;��Mr����!�Y���{����3�3�d?C
8'�H=��8��u�!�W���5��Ň��q����F��݈oDJ�4���a�$Is�1
���V6����mX}h[���u@2-���D�A���x�<�唯���}{�\�4/N!�(�e��h$q�"��G`�3r�cF��D	����-m�zC<&�u{|����Z���xZ�Xs�VJ��]7�m5���;�R�wo��h;Ymw�����c���,NpȺ�6�;�5��3ur΋�n�}��1=�;��)��p쪡�"Er�4�e�ץ�8vw�dh���M冔���=x�4���*yMdA�����~��R����V~�;��^��t�;�//]�W��d¯eg
��y>�Fy�ރO����ϼ�i������\�������I�~�/ވ�<���v[�n�����?p��u�)ib�y|Ȇ�>�2�.�-��=�ւ �5�L��ƨ>]챱4� u�8X��ABS��I{Z�����m�sG�~s]�z�w��F��A�� ��������t���E�:�>�c�0����Vwv�i���|Z�����,�T�<�ι�jm���iJ���'��Ճl+��zk)��o�-�.�8"b�ݮ=�qo:ke�SYbw�S��0�5\�{k噯���z��M��|�E��.M�-�g{�Ph*�!lH��_%�9;����}��l�a�l�86�ͼ�(Y�R�˟e���v6����D���t$o���a��,�0qk���c�ë���[Vp}N��XЬB����ȅ9�� ��������ժ��dn���Ct��8�I�FGP�S��es��Fn������{����r�鱬����'�g���7pL��l$G'1�q�-��۶�J�����Lp�ңwb둯.�7�Z��p�S�{Xc^Pl�Z3ǂ��{I�>]X��cc$��Y��Ԯ�^��Hꑔ,~�o'z)Yʼ�^b��ood\68p�34��)�K+�ͷl[b�a�4��%87+(�7��-ɗ�*%���tOwh
��J��wX��ݼ�4�9�v�j_gke˒�=V�g/� z�z)�FKXO!p�G�f�s��p�q�b�Q�L���k��j�رyfn���=��L=ܚ6Mt�b���Mz�ƽoaܡd� Q���5�oo$��;+=9�bk�8w�UX��}�	�C��N��V�ۉ�vq���Dq�Ut+��#�k��+U*�iqj�	%�Ɏ�m����-�5��&�E��ۋ��c_B��<��6��;����p�l1@-s_}ݢ>�6Ҹn����^#���*j����7&��a��,r�l6g�t�������=B;T���9����ng}�닓lڱ
��Fp�#>�0U+�j��3�;#:��_�@�n���r�4b``}���<wԭ���{� V�N��wԿ/H�n�M꩖oO�P:�eE�=�e	�B�����MM�vD�6��T���5�\�,L�����w!���2�M��JLnLe�MfS��a6F��Z"\C��b%^��7�8g��'��0�8�"�,O�\�m�nig�v�u���s3]0$-�� �@�S�읻��r�}��v�^����O��K����� ����JQ鳮�m\����6��]4"��4u�p���v-�י\ݎx��b��ɤ�=�9��Q�~�;�9��9��6/��W�r��5��6�(�kp=Uo��i0��|3*5�GH'�wq �F�-��I�S�"#M5\s��2-53�"1��3����t&�o�Y�����5�[�q���#��t�����
\➌�7/H����};�כ�;#��Z���f��i���!笃 �"}��
�3�Ng�-c��n��~��p�f8���8	�yU��&E��>L�o�m��j
˚�Z���q�=o�k��f8pI	Qn��`�IF�;U�������t��鿮a�A��0c���\��p�V�M���9w����w��4H�ì����{�;ʧ�+�B��'����Xl�M�~>��$D֘A�^�h��@�l&��<�p���-���=v�b��Z�IN]Lۗ'Ϟ."?xUk]�{uN���G������w
X���Oy��l`H7qv�����e���W��fL���F֘�jy������l1Ak����)�:��Ɲx��M>��M�Ϯ.����&h1��ܬl<���I�ɘ����:\J-�}�o����Sn��MS"�?6��i$���v��q��KQ�V�c��ⲙG���|���O���t�P'�`ڜ�;�|���z�f
D>�u	���7o�޻��s�=�u��v⃸0���Q�3)nie�0�B�²���@eY�=�[���?&�w7�h�����Poe�|�k!�o�8����A�ugc���ƪ}�"��e���;�\V�(��7b�8���SG^�y�{^䍾2k��*�{Ѽ;ǹ���,6�N��n�&k���`�/�#���>3V~��5T�o��`4���r��<���ݷF6�#n�%�=��֕��|�|�y�Br_TDAF��xXc&~��*�&�[V�Vܵ��?$%	85\��]�诏Z�a�`P�:B�!Vư�j��Mk��샛]rg����l�������q�}�������{�0����]c���fyqq��;�1B"�%,�y�w��ݐ������Av0��I�(��4�V���V`Ľ�K�4 �*���1y{�M�}��o�	�s*M�|�42�Nz�>���}J�0���B�>�Hx���3u76�&��&�i?�`��6#�k-�����(��<�����`g.~D���IFo╵wO�3���wǚ�]&{�ς��-1y9�|�5z�� ��w޻��r1�g5.M���`��a�;@�3�y��%M�|<���(޾^�q����i��8J�32
�105�e�.�!�,ܰ�3��&��Km�Q���n�$ļ��ْC�n��b<rw�=�Y��5z�g��I�H���)^��YM͞o�m��:�Ȏa�5�+4��.�`������{�X;�m�&���zλ��g�%��<��ψ��o��z�e=��f+vN�d��^�A����&e�{C~#��93�_
�
}w=޾xxy�]��5m�gj�W����ۃz��GG�������>SG</�5�]�?����������bKv�!>o��z�e�ͦ�4�g��o��o��E�'��;�&6>�#�=�v,�2k ���3����ج�و״qr
�>���yO-��a����-7�G����o��+W�4!ܽ��<=ɥ�{��#�@	����xN�7t�ͥ�A�\���1��/#%�nǹͦ�CԺ��z��r����^�����#�n?�!S|� Ė�34��K���z��n�V�q�\���1z=�����[���-_{y���g���ߵS�q��!�iB���2xS���e�%D�>��i� ���Pw��m��pw��N�:�^++�E��֢�L��~#���S�۾�(糽������N�2�54�%^h���̺m�[b��n��W�R���X��v�^@3JZw6�KY� �o�WP�z�A�'�j��٫�_E�L�3cڬ"�gQ�ة��,�>ص�Z�{����*=!�!Z/�ӵ��_o_
{�}ʗ�qzOKej�7��� �ߤ<T��u�͟��f�u�-��{��u�kM�_v^����������1�ꣂ����3��$�1	5��Z8��]��s��qI���S���2��&ҙ�����w�����0aEVlŹM��3����of����'���hv����Ӱ�<�i�Bͪ��
n�_�~;y�}%U��x����ڧh(0�����+/��0���{H��qU�?og�`-ךƻ�q �Ә�,u�r]�I��yb���Ïv��X못f.�펚3Diն���n8ԝ�v�qTU��]ۚ?;^�SQ8�\�s�n����D$f��h��-�MU�E�v*���i����1��Nݎ港cpx�ؖq0q�_ �0���˗�r#�ƫ��;j�j��pmE֒���u�g`����X��,=��h�v�N0F+�+N�>>>>�8)���틞�=�mS�kA��5�f3��O�q��ۭ�`��w��n����:&����||~#G�^��=�킊�z0�z&�������F���b��ڍT��Ӹ��F��bnڈշh��C��v�4Y�]zs�=AD����#Nƶ�3�;�����IGv躲m��&6�9����E�<TDh�]m�\�(����=��Z���{آ��٩68��.ظ�탍�8�wm�DQU�q��g��]=5GkO�wz�ck1��V5LGA�	�u��A&�mEv݌PGX(*�v-��#�EtPU!��u�Wl�5�Z��f�J&<Y�
����1�5DQ��u�� ��h���QI0t(b�3�Ŭ5  `|�w�� ��?�E
�B���ݬȶc/�.%�E�XCp�ũSS	�+pL@e��Z�1ukZ�����&l�o�3uK����w��fwg�){�4% ���!>IT7��>�HP����K�j���zk0�Mg������N>���s�+L��;�kO��i5��%��VP+���65^�cOv���V<{V�u^��[�3Q�n&��}�JAљ[���j��m���*���pX�Ў��g:�8_��on���=8��<�L�-�Ò�o����F0J�b�>�"Sdt�h����g;De����\��{L�@�f=[ռ�|wA8�"X,��#�dJ,;��9kk�ÛGv�w��Qk�J%�{)��a~�e5��s�:zkw�\^]���E����n&�tM����8e�Qh�\���'�b%:�R1H�jn�<�"�֎�d�擶EL ]��Mvp|�ɛ��-K6׺�ROC�Wp��ԩ'�1L��Eh�q�w�Go}�o�j:ȇ��_����^s���o1͋jx6���Ƣ����,�n�'�zӔ���J�t�r��.��O�[T�O��s��V�p"]�X)`�74Ñ�'f%�=�d�u���Mp𜅵}彃�BO1��B�3��~��k��ǯ/Eqy�)�ø�:h��$�m�F����Y��}�i��{	�{�f�}��H�4���( p�8ڍʠN��.�Le;�WLn	���yѾ�Ŝ�e!MH��P�]u	Jc�wb< �Y�\�̤� �nyK���3!�깘rb`g����������T+�X5"�� M�Y��Mq$����B2ԨjU����_P�ˈ1p	�C�PbS��S�W�`؃׺��uff�&���vܱu6bS��5����ŷՎ3�蟝��z}'�%ؘ!n�ԣ9U����T4��ȿK�}�2{%���
�BB�*(�n鴽�p�Y��Nj5�u����M�!흴�Q0�͍��wHn~;��Q3�.�	�b�	�(T�R�4AȪ�i�R����7�Ip�u&āP�\MOz|�Y���W۹�bf���ų�a3tr-Vf�A4y����4&]�Ƕ�z�o
��E;�/��Ѝ`���_�0C]y�y���S�&$���Ѹ���G̉�Q��RY(5$g�Ƶ��Ο���=`���0BO>��z`�KDw5+��F;���p�yJ���PB}k;'��H�P�LJ�fLa���hDH����1c�m][�cp#n)	��i�b����b07�=�N�-T)B����YĽC�Y~�s�yGL�A��Yb$T,l!b]�#{8��wW_�F�\�<���D���6`5��h%�Gl7"b� z���!�N����Od�fd�[�'�0��:�q��(w���ڀ莶�%�ݕ5�j"���
�;8/a1#�7�d�����DG�	���Ҕ��y�����66Y��;N�p�vJn���	�v/	��V%RN-��'�`��v�~MZ-ߔgV�v;00F�r����ʻ=.�4����z�&X�LT����W^܊�[;�͗��U<x�h+Ӆ���o$h�B1��`���:�i�P�ht�Z����}[�����]�+T��<^4�/#h���~g�m]؆�|QIβ�euw�1л���k���
��UjW<5�)=X*K�;P�|��!��;!���i����2rVir�_O�����:ҁi�C*(��Y@Y���/����,��Y�zwD���dO��!�ggjr��0�J�(�����Gz�(����,6��lc�ȀO��U��(%�9.�����W�ޑP��N�Y�����@`�Dy�:	���|�mK7�׻h�棩P6˦����4��Dnv��ߵ��[��0Ƕ&87C`t{Ӣ$�����z!0g}����&	��K7�,D)[Jx-�d���#ד��s���zA�a�8�r�9��f�N�Sp=
��kc%w���+�EV��R�Ż��C���do�F�2e����_>��'�Bm����7qh�m�9�v�����W��`��.A�tb
��f\�m���U��Й-e�(��.Dz�o���sՉ��]�{�r���4�z��*�E��Q�Y���X01Q ��f��c͜Y��8( ������;L��m�lg�2��L�<�DZ��vf#���qm�TZ{c����PxdrOId�r1��t����Z���7=�]I����c����w5�~��jV'*Z۸�X�ve@,����󇡽8���Wa���VH��[�� �M�#�b���ڱN2V'j[���D���!2`�@����L,c��ON��~��
&w_iᮞ��������I��wP�^!�S�΄&�rU�3ۍ��3�����ն�2�&�IP�����o	�����,y��i�Bz� ��s�5������;�<�|��t������:N��)��&��)��׵��fˈL=�Ōͮ�˚�Ř[��'W�7!��J��J}}�0��J.��)�yi�ouO'�bdB�
ȧ���P�=z�O��8�k/E�M�������*����r1?5�	�it�~oW��p�{���\��dd�W�}��@r�G�<�cT!ƇT���[���w�*�=���m�����b������ٍb��޺��Ʉ���O��J%O�1�k%�v����H塴�����gs9�+1��)�^��AC����	n���l�vѼ1�Z��xK�%r7}a��o�E:2�����1�����7^��L�QiŹe��r᳨)N"r��ʼO7m� -esk�u�2��Ӳ&��<%�����8u�ѭ���KS$��z�:[�Af8���JՋAo��r|�y,������v D�á<%���
}�!(��c�����P���{�׫�G�S§�ϧ���P=r�hņv2�����wh���z��4Qү���蚛�L��,����Ǥ��H�r��H:"���#��}�.�<'�oS�s�hvb�띃;����{b�8�Dܒ���ș�ݬ`��H=�$"j��_�"�Cuc�o)����b�~���L�!	����lS�T^=����w3E�,	W!�%�8�Y��ME@��f���UkK�-��3�~t����Yqx0��?c�[�?���U�G���G+��-��C����{��^��|��N*
�sf���ɜ-��{G8k�U%��+�1��-^24�ȱ���|�]��ڧ�&�iM'�Fq��ј�oV�^��;ǐP2F�" H<�b���M��3����{��B��: ���I���y_�B�K�����������~7���/�����%�b6��ͳw���*�����E��1#e��q�]h�{�2]
�עD���D���Nﰕ���)�j�����Ã/=���#�C����{Αz�;��7T�j���T�&2��A�n�C�ܝ�%dT[��l8�"�LV=�����&�)�q���k[Mp��>0��!��#� ��y���
8�N�ܤ
n��&����O�p�,�<c
��}���/7ix�vid!�6��Ԑ��;�9*oJ������g<�4�@���mdLgm�K^�סW<���s�L��z�	����n��>Ƣ�����|LZ~K��F|.Qӝ�����f=�x ��i�H=!�ό�Q�B0A����n%��N�f����%�N��p歗��G1��Lw:lw��%ݠ��Hz Ks1���1��Q�0��bt���;qZ��%*���2S���M�Z��*�f�W�-ݛga�8�� �^,����MR��-sm)��dT2���Z��u1�e�gǧն������� �*Xن[OC��bo�ܙ�Z�0,g!孼�:lO��_w�P~����~df�+�HH[EE�'�o�ղ�K�Y�/��C��pw
^�h�gh��e5E����u#Y+�u�w	�.��1�ނjEW������oe�e�T�D�כx�"]����8dSz@���_T�[<~n�'z�)�=r6Lv{�N��z����1��)7��ZEq�W��㽆n�o�P�(�n�gT�	G�x�ޔ�&�V�Ѣ	ɏ�Q��~?�'o�\�w�wx7�����	7IL�V���x?A�l~K�&�^!����STq����a�&ITH��K��G����]v�0�K*[�z�]�[8�5e�E�5��y��["���&P�>f���Ur5qlb��KX֮�Z�s���^�����&J��A#8�z͜e@dgO!�L�؎�p��M}�(�37+�c�ު�E�˕\���U�,s��X���!>����qR��rc��_�i�5��;��X�&�㛝��42�%�T�봏h3�Z�#!0����־	1I��"Q�E�5-���H�����b�gv�d�n+�ģ��)�!B�l�0���r|�òso�!2Oa����R�jށ*F��y���n�=�)�u��5�
�q��8ޯK�Hق�b@�3#z�y2+�-�&�t3�ٜu�c;�ƪ@'�E�"Mb:p����o'F@A�v!?w�T�Az`N[��*��e�[�wj���\%�76^Q�d]s8�KK�@��=;�?;�A^D9�1��6�c�|#mdޤz�n]�0z�e����m&Ves��I�O��dC驘�fL�0��τҩ�t0"u.|��E[�@�I�Ƣ����e��1'\]�TXW�h�vU~WZ�|��>�0��azxƯz���Q/fv��+��s�2-(�y�(�X��:�V莇��9�����V ��o��8��J�t:�Cmm#w�ٻ�.�	�E��
/{!ʕo�? �{ā'�k����4�� ���32ė���r%46TT�v
��2x�=��x�p	���L��{��%�:�`���0u�,�9e�R9��Ȥ�C�q�1�\��^��*	q�R���g{3��V��ʰ���;���((G��!���9نe��Xk�PB�v~��~��� �뷲��kh�Lէ��?t/^/a�ɑ.���x��x�m�_�%�'W��f�lo%8C��\�k����,8�k�t3v:�3>:"�ǜS9}hw@���0���|as�.K��)�v�7Ww����@�3�d<P�HzJ>�e�N�U�6��*DF��-Z�����Fε�Ļ�=�B�s��/��݃�"��$��A�d��|��6��9A�
�ֹ�Y��-(��Dz���[��H��o}>�}i��-mG���`� ��ˑ'BTy���?�nZ�G������v��LT:��,�G66tޱ#���%s�-�]Jl��Be�^Ls�FQ��6����Җл�=;�X�o�jkgk�MM$>C�����#�O5:��խK�$1���Zy��o�.k^e��)LP�����z��xO^��!�X��|���lOh4���$�E*��۰���,�VlB�����^�p�T~93���/r�vc�<���r{[��qo_��얬��<Ǖ��_�b+'��<�Gg;}�n�īS� wv�y5,�WQý/
C�t���2_K���_�����|@u�ۼozn���ϐ�2S�/�:�x�44�8�������/=j��#�ן�v�Ѽ������$��@��{*d��:r�<��酣R���)�yi�n�u9j��c���ulE��x�Y�/7lS$*�O�LhuHLk�r�iC��YU����QQ�ǣ!����������C<|�S��-�4(W��x�`鹜���SE����c��j]�Ta�d�v$xD�]���H���ϓ��p8v��j���u�q�k��Kj��-l�*��9�y���_��²����
{��+�i
�b[[�1�Bh�lTE�u��3�v ��h2�ћW�0m�kr�E�O�*A3�Ǯ3<���,ƌXgc&3�04B/=�.�B�M�/��Kr�߭�d����J�Bf������Nw
Pߟ^�x�dt<1�:���Em�޲�V���ƃ�A�\<����ęH��= L$ �D�4��-�x'�9�kL�3|Ggs��4�������k�b�cޜyZgx��(��dEc7�;��</a�o���jÎ�y22�����"���̚� �qI���i���m,���^�'	���h�2wO�%=$n拨r�^`�'+4ME�5о��ԈF]�E*�AC�;^��K(�Q9e^E�F�7I)���Q(�YR�^Ҍ��%�'�� M��q#�w��u�6�����N��ňM-�(P�R�:3/�r�VA~�D%٪/�X�ٙ�w�X���^��%;����>�pf�'��V�t�w��ŷ�â�o��~�X�-Y���n�TY�XNY�x��н�DkZFX �ҚObQ�a^�1�ޭ����25�W�4�;���*`|u�e�oܴ���a�jBq��r�K(�k���Ʈ{gOMn����0�d�ӝqZAD�f�0�8�ݍ!
��@tD�I��Juz�S�F�[\nK������o�̳IqZ�6��R|=_8����цmَ��v
A�P�}�J�v/;�s@�oڙT͕����w.��M����L-�^�����"�G�"<�:mَ�l�Q{:�˦�u���l�i�mer���8�k��qzryAt��w�)�
�p=N&89��<�^�s�����g�i����������e�s�����2ML�|����A��%�����
mMX�a�%n.�����]R2�5�v7�'-`-2m���}
�Y�����J`Gp#� }�8��/�E�?���턄U�/�S=��y��}&{K�������#�m�n�k���o:K�����^-�1�3�k�K��#�7�e����r�G��5h����:��l����]�ϔ�{4U�FK��9A��z{�뢩9x�y�n�<�]��3�!��b��I�S:c�]�z�W{��~�վ�ՆN��<��f�,h���:�Q�i��PmΒh�yt�E!Z�P�uN^��l���l�9{U��׫�˾�����$wJn�cJ��P�ӱY�&���dٻ��_X;�M���3�8��X���{�o^�qEF9�VTCkc��7NC�|�/w������ܖ�:�هɘ�k[��U���sH����8��Άz�}c*�E�U��ҝ��A�F��:Db	����zs ��f�r^�]����#S+�:A�||º��AM̭8ѥ�WE�oӫ��������-�_��ə��%����Y�/Tf"��h��V�.��G̒����xrĪ�)��,��j��-^�M��Ä����d+̧��'��0���%���>�]���xs�s#��di:��*�c\2��DJ�{0��+e��7b��R��e����6�Hz�čX�@��]JM~���N���I���Z[г
j[hVæ#n�NJ���=��I����#�<Y�������:��b�WUZ)���:��D�l�ّ����2�N�Z32��y*��q^�(��|U�,s��<o�F��O�Y��^�Uqt˽�����E�>�Ow���y��B|�1�qe�;�>bO�w�ʙĩ�����~]�����O7=j���N1k0(zlnD`�o�.����1�׹�v�t'�I*�<+.9ɋ>^���|]�\��${�1v{Z[p�9N�a�W�z6�<��<YG��x(�;��+�ó���<����_`�{�Oxs)w]8���r�za�F&���)�]�G,9����g���v�~���8t��,�ӣ7Gt��n;�ܯ��\j{<���Fޖo>ռ���˜��V�̘;6i�5͜�V�����S�;�k�!�G�y�$�,1��S�c�ץ��wp�o�>�^w>~�,7w�d�-���9qm<��{���^&0h	�6l�26�n��gsg:ﵾ�[���5o^��,�l�@6Ň6�$�$SR�1�7WL2�3m�i�D�uzĥ�����e;IӰ}�}��N��5r���u3:K+k9Y��Ga,�
�ڦ�i5w�Mȍ֬il�lo���Ԝr1BnZ[{�ɗ��b�ޏ��v�Ӵxb�l��L7��9����u��yb��RiTk&��a������z��K^�ļF�P�G�A{Ӝ
�{0�&�wLH��.�a"�����]�6��T]�y��aꇗ9Z�"蘡d��J��ڋ4�흓|'��i�oU���E��j"~��[���^6��rp�/\>9Kͤh!S~` �@W<8�_�\��PL�V�KQU4Sn�Q��� ���Q$�OݰPP�����>>>�f"/�Ml�m��th��tE�PQ^���b�����a�"��������|Z�����")ݞ���)!��k�DU�D��I�GZ����1�������PU1TS1MRk1DIv�����kQD�;b�����b*���M����������`�m$E:4v5Et���H(���D�D^�t�WgZM�QQu��ĔI1L�E��c��U�QET�Gg54�lh�h)=�EE�J��j(�b��b��ɭTLų�,Z��h�$�
�Y&Ѫ�5�Q�݌Qu��Ѣ�*��h��*n��*�(���**����#Zb���f�Y-64Lų����i"vr�DQ�IG�EGZmb
�~hĻ-^�~����xﰈ��ud�������qgY���z=��s��m�ռ�ͺ��b4A���*sX0Z�\���"���*qdko�����v�E���i�jL:��Z�OO�l	1\�~�����1#�r�9Z��vwL�eL�B5��LZa�bz��2}�v��e'�23L����<�� k.=V�;��I�ߴ)���2<�g�!3�`0ZDL,scja�������+u�L-�zfvS�+��-n#�ǜÄxE��x86D��!��"a'W���s��}�K]ʍk�5R�;c@�|8�=�Zf�c9ی[ˑ�i��5���y��["��`0&P�a�-�}�ЮM7�����]��m�[�<;Նr��n�A,��Fq�64c���Φ�rf�*5#���]��g�zN�i�9��uY@�ןSf� �Z��A=yd	b�N3�1���/P䴶�	�EH���H�e�̐�:"y�W�']�j���FB��t[��'V�B��U���At���/%e�!�񍿧*_��:&�P�oB�,���nK��%��tBd��ħJ��,(\���ݍZ�&7��;Ԯ�����M=Ӎ��#adHقW�%؆��f���;O]�ge'�|J��˰'�z�ڎ>�vo�j����!�;cS���"0�8%[���Dlv���/���UFx���K���5�U{�^�Z�����o�A�q$�ͽ"QlZ���!V�:�|�~��>�Ծ~ _Oc.^�/�0`��Feq�L���N�l�'�Y+�<�Qt��/�e�w�xa�ZF4�r�uH ����F�<�7��v�{��8�n@�P��X.�z�rm�u��iZ^F�;5�@;�?;��p����,�*��n�R֤CI{��
W�(��L*�fW<5�I��T�4��0��DóOd=�cvdDˈI�]�K{��w$7��L�L@L��uEs�5�,ߌI�|U�<ʬ+�`��>�̡y�\]���������M�H�}r�3�~e�L��	�{�G6��4-XQ+\u�ǥs�J	{k��93IX����p]��\9k_��x7��`s�g�:���k�X����ږe��F\s?��@ƶ� �Q:��#3nU�C4��泰0����dȗx��`<{D&���1�����3���M6�m<f^�d_&b�*,x.�L�zfa�����7�_<��
��_�ld��CP�'7t�\r}nr�����y+�k|&�����@�P�jZ#��ok����f�h�zO�VQ%�����E㉊�y��Q�����Z�7a ��㐂z	d�9�m�ۦ�x���Ί���j���yu��T�v���	�Rs�:��2��rv:�cC2�\Ӻ�r��8�D���������s����i�6���5�e����9��S[n31%Rd������{!���%?bX}v�
��CK3!+�LԠ�lꏐˋ'&2�� ��`kv�t�C�����)�8G0�a�q>3�WO`UF5u�9R��)^���\�&_��p�����֍ȟ|ݘ��eJSq:
�1d]tX���ǽF�7\/�@���f{\_�ӳ��^�
3��h$e?_�xE���o��:-���!�����YAT�F��c:}�,�Oۂe��A�9r����IP���ǯk��Ox��C��0��w�X؝���Pͪ���L����>4���>ޙI��d�g��i��i0�*�ȍʯJ�
��0V�����1y��H|�ɛ���^��4��G%C��Rt��5�E�{�)�����K��۬�iPh\]f�ݵS��1t�����li��]Rr�5���*���z�9�����q��3{݋�W��̽n���� \K������<���֑#[��SEՍ7Z�������Q��A�\rF^"^9T՝ȗ�^�u��@�z���l�s9�Nk��4گ�%����l���s�������0ݽ�� J�Γ��NB���m�l#����X� ^D;k�ۭ]LEZ�R��_�Z̆�G�Δ��n�[�w�ϥP�6[�g�ժ#<�'\���.rK	�&񁍸��yD�h�Jh�N�r'eCrpb������%OA���&�f��)3z��Kl2ɉ��ʐP��CVܣ�ޢ-;M�qD R���w5Ho[i�����`���	��=�D���f�|=��Rcl����L�q�ș���Z@r�=a��Lg �u�\�Z�S|B�׵At���t^�C�ݐͲ;%��zHz�(1^��)�WX�c���+�9Ջ�+n۰� ��=aָxQe�mFk��&�ݬ`��	H8CQ5��';@ҶJ�ct�:k_�P����=[�?��z�;���+L��	��{]΃��	�&���nw��|������u{7�\�o#^Y�X�ii(Z�;Kg�#w>�8��Ů�;��n|=�pm�����{�������P���	�G(=y�g�M<.�.�Sp�輁�/��؛we��ʹ�Z�����DJl&dԌIu(�0��ǾV�_F>��t��ǌ��M^�9ڶ��,%��Gn�!��6�B	�q�d��R�er�z7ER�`�9؟K�Di嵓k���6
[K]�@��Ȕ��!���iH��])�r�	��"�ג4�������ޱ�����ھ��,��.���C5��*Y����*��v
A�P�F�*Iؼ�*��|nd>^�E�W��.��b+�����HI�hz|w���g��]����O%��[�f����z�.�͵���^�(9��Z��Ǔ�'�d:8#~;���z�7ɢvx�Z���"�����!��c0DR]亼�:W�+�2�k�"��Oqbx��&�`�c!�)z��W[y[��3�y�o�F�>G�|�¼B=Ȋ	�j85�E��'T�9e{<T�1����'�nv���^g.m�CTYts����<���L$��>`"� )֡G8�x�)�Ё��9�u�<��s�������إ���H�R�
x�x�O����`tb`W�
��ܱ�Ƙ�<ѵ�f��^6����l��nL���jE1�&������-2m��Ϡ*�f��ͳ���Խ�'�r�v�:sfw� �����?K�>n�
%4�\�uo�Hϫ�TW5 ��?�-�}V�ާb2Nj�C���v�v�>��A��!���˲}�v��v�pB1,4 k==� �ys�����Mk�ty�=ӢdP.�&��gm�D��;05�$Gu��{:�rnP�p�7W+�Y���SN�r�b�Lq'DYz�o�D��A�4���u��{Aj�:��=�uⷞ�a���򤶙��*W;PJq�j�#.��ԟ9��l�w����5
!��b�#�.��&�M�i�B��՗��X����A�RY(5$g�b�n@�t��EØ��I�DN^�&v	�,�ĺ^�k
�n���.�v��މw{�o*/Os����>�>͞>^r�v�JU��vl:z�&#oV|ed5N�Ͷef���@��۟�OOߣ�����5d�)��aM��h�ĵ���-�Q�Z��}֮n���U��Ɠ�����+qf�em<`����!^D>c�
7#��ȫj��!>����zYX�]�':��m/T��{�j��S�o����հ��g!@�����*by�F��MQ����A�=�1IխT)T���"9�r6_�J�Iї��:=�l�<���n�<&�X�ފ�,���=�.�$vP����R��JU�3:�c}r��¯^�9l營�Z�%RN.�l�	�hUӍ�>5ä*���nc�uH�,���zj�p�K�V���|�(�%Ɓ�8^���O��!��R��Z�]�VH|����9���+P�ν����jo�U(�&m�u��iX��vk��w�~yۢ;n����{|�����_���e
7�v�
�fW<5�I�,HGjJxw��
݋����*�{4��٢v�'{e9u���̛o�7�:��՚�l��.��,)gO2�S�2������z���+)4�of���s�&�2 G�(T>�4�0�9�u����`hZ#"V8��J��ő���xfO�f�#]U�;�2c�[���j`�g�BD	���Ӊ����Գ-�Ú��y��smF����!�V�in�e�Sx���z���w�mKT���^��{��O��PFmۯ<%mN��}�5C�<�!v>��#�EP������k��@ߧ��O�g�q8Y���U���9�ڐ��h�b�N�DFV��[	ލ��*"4�ˌ����I� ƄƐ� L31�{Ԭ ~Tְ{F�(���z��̙2�H�W�D��}����g�k��2�M]�i��Y���E�/�I�oz�7Q|�lvCbzTT�xu�q�&�v�m��q�au�y�,(��6��a2,���Hz�PnF�l�tM�1���u��Z��7��7=��2(lW���m�tfV��Ԩłk�&� f�����Ж~��6k_DK��]�=��%��!�yg��zä�}sE�1��&�:�k�ޔ_O8�D&�^w�Zӧ6]����8��6�*yX��сa)��h5M�C��i��%bv����>����}�w��]��E��\ܖ��T*��vл=;�X�o4������H|�����[a�����O���|�Cq0Yt)��1)���LP�� قե.�9�ٚ20�O�ؽ�P�5v.'t�f�0SL�h$v��L��ĲN��X��X ��(=��v8�d��2��蜭[��v�d�C5Ȉ�`y�uAhi��)Cϯ����"�z����de���2(^��<�E�Z1���/|� �jș[;ڻj��I\��M�'7VsW������[�K���x(t-�f�'�*���S�'JѪ���֮����p��o�y�	��V�Sj�N�KR�3s+ο����s����lC�ۧ��1ŧ@�#���x�+�!bP�b%A?������������6< ��B�li8An��!1;r$��$�ʮ��r-?7^M�i�{��0����������I�MIĸx`>��y�k?��SEՃT+߻9`��tDy�bi��Y�(Y�R�\:�K��R���sh/NdϬ�u�}"|���d�^.!Įɞ3Ydx֮<f�+6� �V��=+�҂^��]8���ql	v�!�Bk�>��Qӆ�4�]�L�7[r��w_��1yj�f:�v)anlʤ��(�}&=�8���f:b�:�(�#�2�o�Wݸ��X,�A�y�<����bD������[�����W��b�%�>1U1��}v[�Xi�:c�2�f��WÄ�H�"T�Xڌ�K4��ci�C�"���a�1BF�O[�f�J�C��-�>P�^Ȗt42坩�r:��w���Q${")0Et^�۞���^�uG7K^�8q�&>�*m=sͼ4�yg��-!	�%�z�}<�9�|�I�{x����o:9�ykY;,؀[(2��6�r��l�|i���"���h��E���~���U��}�D�)(Y}��C��a�hݐz�����m.�L{#�ʊ
�0g+y.f�뜴û�
q-�`��-5>$/���<��''�^�����t�P�A�Bw�d���$۽+]x/x��0���#:D7�(�
�[�ӑ��vd@�1_�~� � " ��bB%����?�����e�Pgg^�>�E�W;^���%6�2��Ji=�Q�a@�f=oV�]�\c�E��g��ץ�8����ò�	^B%���@�>ӳ,C�*��'8���R�er�&�}���\��fĚ�YȜ���L���HP1<f�i��W�A;$���N��1�j�,m'�*�;���wE\���\ż�N���ty�f�t�]���eGe�#����T����ڧ�u,������q��O"��,9��az|�>σ����	�f8Cf�-�`��ң)��^��~}���M����s�z/�'�K�\�GP��H=�C����r9Ān�fN�u�{um�ߩsO:ڹ�N{zm���"�~[#�Kב��'�q���ѽ:��|�@0�R]��ù�e�;�[&�:�C�:Tj�'6jE1�&�������MȊ�,�B����٘��k}à��y<t�iN����Ny�C��;k��.���dRAD�A�@�^A=>���͎��t=��qmi����UB�r3���Ŧ[��2}��h?����0l��cbέ�:���m�}�I����,�K|q]+噵#g�f�Cj�T�k1˛P�X�Y[�ڻ*e��v P'}�_G�����y�ꛐ��gkȮ�\N�ҭU��-�#c�!ۗ���7/��GI�N�Ck#�~[�S��_~�����_�?� �� 1=�<��4�?���pB����ksp�-���#��l4�;L�	�O�ac��{��Q2�u���߂�پ��;�BMs�yf,K�q�DYz�o��%�<��h���g�I����iaʫ;�꺻�V�^׹O�fY�h��$�%�6�F]����<�/CpP�`�$�RJ����:���̎��nyj�B���ۯ6ۆT�X[5%���#8���Z�22'ҚόI;���J]S>��������"�#��V���B}k � ��@�4]Z�Xq���ih��m,�31۫��o��Q��S�"#���E_���1:�Y5�\��2���n��t��)��y�RX�߇/9�29ml����1�-�����N���v�=���N8�q�9�3+�k]v�������J���j�*I��l�	�d[B��ZޠC�`�H8��1��A2��0cT�������F#��þS�Y�Ɇ�	���"��K�qӅٲ�_���l��}�r*_ji�Z��=�A��*�Xv�0ճ��D
s�P/ix�f�����ϣ�� �������T�<
�x@C�h�5�=->:�2��/�;~���f��w�o9�vt�˅����Ӵ����:F��P#3#
3��q��+j7:��V�ݤ8�Tj��]|�FE���o��9��Mf��� �=q}M�Ԇmö��>��"����\Og9��o��Fi�V��'%7d��9J$���t!�Y�c�<��>�YӅa�A�����\Q*��Ke����v�L��s}��Tj��{����c5�c�L�{�(w�"���,�+�m��ش��|<����Z�%9�Z���sW�*�v��Gr9H5j��)�j������h�U�7p�-�1�r�v\��]�|��i.��a��'-Y�Rsb��y�K�bk��Ą�yf"Q��hĈQ:B0-�ܦ?o��/İ(¼�-����j/uҚz�h����\V�P��Jm@8�ɍ���n�S�6��8��3W=����x��@�8�OC�����(2ot�ð=wsҫ��'���^ˑM�.%�LӷTҺ
�M�2�:�����}r)��N(��{A��1��n���z�4w�#���{:vM�(O���_��pӾfB|�)��������g� ��x�9�����x�94"V�WTn6X݄�H[��CO1R�f5����u�c~{z�>�����;`�hA�y�׌��Wȃya���s=�[���E�U��E�.z��]�/���s|xq�-�no�>q\�sǒ�@2���-,�
�V�(�8b�qB
���њΓYT�����/����o�\��L�Թ1��U�7�*6�3�+q��_�j��f\����T;7}g�^���n����#Q*N���c���ѽ���:x�h���7Q��HA*�5�W:J��X��^�>�Y���`�Վ����eO��7�����!Z�����Is������fdܪC�ϟ{���wS7��FA������3�.H��.�7�r�W�ǽ������s��'tP�TfU�]�[.2�`�x��دjhpd��e�j��~2��2��2x��"�̭4feIր󸵽��E�]�C4{�ny"�,{��},�WN<q��/��ȏ���G��m]c:��9]�M>]~����U�B�o�����O���++�~��{��~`-���Oq^�Ͷ]�o"�K�q�O
p���5R����-'XT�ih�j��2�n�.�kB�|3~��p�tGS���v�+����w*�xG�@{&���蟟�,��:d;��P~^��N�8�M)�^R����Sb�8U#����z�I~Ұ���k���s֯%�d��)��Ȉ�Vkud�/�9����5{5�*x��ދZ��D6�(kw4��YE��[ݼ�U���ޣ.�=���<!Ia��Ow12�u:�.\��x�)	���4��͘��zn$И[����NJ���h�bL3������m�)LE@���p(nMD�-:`��f(�h�;:f"(""����"#֢'�������U'�,c&��b�g�T�Eu����5�&�	1���?��
�*�����������H"�4�h���
�(�������������j������L�D�u��)�i6�TVٶ�D�APUQh�h�������QD���Uh���)���b�� �*�#mM�E4�b�+F���4U-HM=V�)��&�)����h��ERTQSDDM4i�]�4A_`��T��(.�h�b&�����u4ŭ3Ql抦"*"��Q��+�v5$SE1TX��t��SBQ]h�
�_mx�cEQ��55U4Ŷb(����*����*"(�{�kEA]���"i��������Z��T���:��Ti��G�������պ�h��F�`Ed��u�3�T7��O�RU9�T�F��Fɺ5jd��<X������7:��S���,�3?��" bbU�RaP({�{9(^nՅm�-<à�^��E'&rD�;I�U�\��\��eP����<K�.ME�9��qwl&��b=yR��u�8��t� q�+�l܊:I��>�tN=�!�ȇ�*I'k����&�����&0;"iH����*H��1�:�soi�K�J��D��Cf:f��*���^_f�u�
{k��O�P��v�@�+��Ŋ}<��ˈ���2Y�X�Q�N�u�{0�^I��U��&�(���z���� ���zH4��F-.nɁ2z��ʖe�{����Qa@���L�v8���T�x��n�lg/>חz�~.��A����Ꝥ���k���04+�0����"�x�����PnF����&�-DD�"�e�+�u�;;�c���39"���I5�7s�<6R�*\&��8;�ǃ9)�E�^bG�SRo{̇G[����~��g�酆Iƈ��/2�-�g.63��<�>Ya�;.V�^2��5_(�#�CC�A����H���46)����V���!�i���pբ�
��S�;c�E�m��7��%+Jy�Rγ�떼�}=�\�xM�b����Vxa��}��s��'Ax�l��d!H��;�]�}�TR6z������<�ŷ��8{�Ƽ��qva������2v1[M��j��Y�g.�|]8�`�??�� �i�D"% �����I�&�m=j-m��'l>bR,�"S���`��z���{gh@Ŵ��H|�Z���)��ӝ���?)W�i �jJca�JtT&	��%@h���}��xOV�ϐ�u�PW0�N]����d��~��z�hv�oL���$�x�44�S�k��W=
�vD���%��N������FP	���3d�&���1��"U�j^��)>0Fa0,��☖J�F�B!���l�8zv;%CZ���^�`�i���E�M��	�ۑ'|v�8�������ώ>��^�͜�e�y��S����t(~nN%�����=�d��#�kumMFb�8,Q#$xT[��_v-���)ʌ9�K�X���8����B5�K�C�Z� �JyָM�����ʭ�E���-l�J�a@q�\������p��n!9��������Z�L�e�:�TK�z��H0����ˌ�Lọ���3�Ǯ3<Ǫ�z�tՠj�mkb��evZ�!p=�y�<����_�ջA�kݲ���Ǥ�$87�����M&��&.�X�hj[-a}:�>�H�p�:|ۅ�bk'af`�V�Afs����+f�\�Vr$IE���ߌ��㻨�����'�8G�d�9Pg���`������
-��W��(Kk#t�PԲ��p�n�	��,�w��U���H�U�k_�G$� cE�R`D�PZ@

{��ƒ�Cz��p.b���A�w��h|.&%M����t��gv���s���R�L�-H�qi1���7`B�r�i�ѣ#�DT:��g�D�C���N ������R٧O�K��=��z%�2�4ÒYA
�%�<�ͧ�y��ֆz#�Z|���Nv�����=M���͞ʫ�^:��L�R�[7`]8P�&�9T�������t	w�D�����є�Ñ��ٖ�oͩ:=���c��'+~����%7��A�iM'�Fq�x�f=[ռ�׫m���=T�]��'�����t���+�&�D��x<��W�sP��/��Y'�R�e�juw�,z�4�WRG_s�W=���~zkw��vl�xLc@#@�^�DJt�����_L`F��qeu�v�d��ԁF�[\nO5 �h�#�4>3¹f��\�`��T8��u1'�8my�9{�]�@l��X�:�.�{�E[E�5 z0�>G�|����Bm�����촚M�4L����z�4�ΊSi�t>���h�ryAj�X���!��a!N�p�`���.[����"2F��$��*� 8���ߞxz���+=�~t_�{��#\�q����a���J�j�t�,�T0�=���T���XP���R��G	�4���hB�Srs�Auj��}�Ց���#񳻗�a�9suz��NI!rii�D"U�P�c{�����9����.>1,K��ɦ��i�k�2����AOZ�I��qxwn|ga�kK����oB[]���w�S���vN���\��H�5�&����'-kL�z�s�
�Z_�\:�1=X�V?w-wf����@A�y�t^��������L8̱���m�YvbXf��.���:�����蟝��Cb`D�*&��]&��=�x%g�gt��Q�Srp������R�{����LW5�-�P/a�G<3�������ڑ���A�ݫx9MU��/���b�z�5M.SEډ�bĹ����9��l�w���h���F��S�)f�W�'(��ٵu�i�v<�2��m�$�P*q�j��i*7Ӂ���`V2d�h1Һ���]���g�HA��[q{����x��f(,�5y,����g��8˴O_77Q���̛Dvj�n�Ӽ'� �v�yaP	�9mAt�Z��	�d	c��\�A�����'0�iz�=�\O�t̘��r��W���x.3&'��S���!s��cԦs�mC;է����3Hz�N�_{:�ǋ��jOz�vho|<�W�ی�L�)��w�=:�A]j�=����神�&�0�D�N�!��K���އ	��1;�3ݳ��޶�;�s�ܖFFk~�1�r>�ׯ��⟳��ߟͷ���߯��?��("QX�Z@JQB%hbf�6����K��IP�bUԷ'���������5ߦv��.��Ǒ��s����ͮ޽ڪ�Zػ��v/��J��U$��6q���-�W�q��i�:A��!ۉ�kW��*�3�s��r�.�4�)��oR���LU�y^�\h����'f�# �r�^�}8���� ����^���6�T���ʎ*���JD6�6Ⱥ��9����뽚�v��*��s����w��fm��Mל?4Xp���7C�TQs`�N�a=�2���I��RX�n�Q�W���Y�nb_�N��P�y<;�G�C�Ϝ>2��Dsu�[��ʊ�V��d�q\T��딵�e&���=mY�ȵ���G=ؕ�dM|�@����v J�������,8X�`�S�\���綊u>ݐ�#�'�҂^��G0����sPw����g��19	>`�	��'���MM�&h媋��@�e�[",�TMKsQ�^�^�90!߁p�h.ֶ�HMT�`Zt����Jrf�:݆m�����D�`r��"��5�m�.�-���ߖ�-A�/���J:�iW���	o{��xϵ������OT��9�p��oG+6)
� �Ɨn/e��o����: ��!)�^�	�_7��ڈ�xo]՛�q\q�dv-�E}��Oe�|�oˢ�6'?�}%q��TW+��s
p������  ?)�X� � D`�����ww�V���܋q��-y�lTc#ú��Ȳ;��'6�����E�pa���p�{�ǜW�PT��:c·�^Y9�I��v��	��5�p��V6;��+uκ.�y��)û�Q%^inZ��k�����������Ʈ�Nh�ln��7qm�P�vټ.��H�t1���B�Ru��Ű�E�T9��L����]*`E9�����T�T��v�Kʢ�V��3Yt)���!2�*������)�9�Qy;;�r�������jzأ�{H0�4!ق�CP�2X��AxNPJ`��	*�o���
�GBh��C!T��#wv�����h�(>p�|�hY�a�,�ze'X^%�u��)�$i0�ZP�֕.��fnu����p�Q�ZBvl�D����o�ZD�9J}}�0�jQu��µ�4E[Iʽ�(�����(r$\���7�;��MB�li����L$&4v�Z������7P�(@5�kŹC�IKƤ��9d��t(~d�4�s�S��kkW��kumMG���;j#퀦c�Le>��=B��o��d������n����C��~������?x����Y�������1����5����	�����Y7Q��x�B��X��e�:l�u����ٔ2օD�Aa�xE�����Rh��d���.a����ӣjLT]�������(T�U��D""JE	 B��_�׿��������~>���K|R�c��K! LE_�J�s����NhH��)@9�'bʔ��e^�s�!|@eM16j�[+
Uk
�ҹ�(%��؞jY��|���H`�guj�*�tգGe� �!�b�0��Hنk�n�\eRcl���ɟN?�m��;FȉS��x��'s��-y�ې�F8t�]�6�Ƕ����!�dvJ/��=$=D�X����V�V%Em�{�/;�|Ь���v����=6
,���t�����0~l���.H�J�Dc>Z�-#�"|�/����_E��b*�dK< ���!�Za�~��9��^�Σj&�2ڦ��.���ǅ���IhhT��K��dͧ�xk��#�Y黙n��wo��*�l�ɼG��
����왶�ES6�;(2�S�$nC�6�'ƛx]]�U
%է흃7{,��ČS$�ȋ�N�k~���o)�A2�-cM'�հ�D���o��B����Gs�6��lN:O����,.b�����ge��!n+�K$�
SM@-<�](o�������G���=�*p}�s�٣x&�w�6��N2_]�{��?ya�����5S�b�pu;�36̋cW�^�I���f�6p+ps�4�ـ���	�6R���M9�W�bv1��a`N�ʴ�ε���Y
��Y���ü������� H�$D�Oy�{��{��v����Q����1�<!c�Q{d Ŷ;䋁�)MfژL��#�d}�N���Y/K��>.�m߱�J|���3��\?�vz2~���J��Ty�f��JY��ڞ����l!A�K�W$O^Dޣɜ.�E'6�sȣAm�z0�����RG��Ȅ��J�{����vUej�ܽ�q�=���4�0���zOȧ�K���:�w�9��1;�������%r��I�D�����'<��ud�wo��U�\�F���Tw=y>;��}��E��uY�ϑ1��J#{3�^B�w�k؇d�huP�u~�S2k��ғ���M�X
�й�;�Z����-��{�0��Y�5��n��=��  �^D?�R�M���"�.S)�S�Z��]8��]cE��&��x�m��~��q���?[�Sè�C�<x�iLZ����w\�~�{jGR��.���kh�j�|�r�)��D�M�3,l�`��2(9���
q1_�->���gC�V3�����Ww�KC�O'pЂbK��,Ť�0�A�.^���l�w�C')	��Z���b����=Cٻ<jĽ@d��=�����`�S���k�0t�<W+�Ap�����C�>H�-cK��o�	�g�XvA�Y;_iSӑ��M@:h;׶��U&�x�p���ndS�^Vo[�k���j֎_2o��\���� �J	J)��"^�f����o3{����9��������LQ|����u]��̳L�CzIv*-�m�e�E����x%#
Z��;c�q�����v��
�t���ۓت��u�جj���A��,��d�ԑ�g�7�5����/G���[i�3�֗t,#� ��|Ǧ ��V�'ֿ��u%L;WU+���Ϝ���>�o:��ƯeEê��fp��r,D�S���S�����sD-;tƼiI:z�b�W�t�+�XZ�R�J���'�T\:��g�$Ao'0�v&�OO�z�\f��v��'n)�s��I��Ju~)P�bU$���tm�W���Fc���#����Pe�N�m����h�p���h�n�b=�J�,�x	���"���A}��f�xaɢ�j�./������($(E���~�� ����T/T4�ꔞlf�X<^4�/#d�u��ĝ��iÄ�����vkg�A��p`����zQI���P�`�&^�+�@��ɔ��;���;fTz3e��݃9kj��P�Jxwf��|yp��,7;��_=�ά�S��~1'\Y�e�WM��uh�>�Y>�3�1���+��j��iV4a1,V����Ň,,����y�iֲ�ê�,��Π�)�`��]��޾4�e��wJE���� ���sqW�R�4{л�׎�F�,�/�3>�o��%�`L��>*��_�cߏ������E�J�0��Ī� �
#H�
��`�g759��uK�t�Ua]k	Ov[��=���i����-^�0���p�K�}=�4��osk�'�ꕮ8.���A/mr��O�P�j���:	b�����38��.�[�jP��W����{WR̷�Sn:�a�Mk�0�9DԷ5�0�j� 2%��fi�;�l��]�������V�&�9>�n�w(��O�K�&Y��񙆐tE���hٿ�D���V��-�Q=>�&�XR+��J��I��^����܈Mo	������I�<pM�S����̺);P�v��T6&���C`38	A��̿zw2���S��&���^4�Wfu%x6�ӆ��=��G�T�}7B�k�7n��uLC�yg��'"�h���Ʈ��U�i܉�U����{w��s֢��-R;^��eK2������su����ӂ`��]�oa%�y�%l��l�A˲��ن��"Z�	� �P��/�`�tL����E��Lq�N}2��������X���`;+�4��<��Bc�bS�*S��IP�Ȼt<@�������_Q��ݫ��f�;�q:��Mc �*(��Q�c���e��+C5�ƙ�u}{Hp����ܓP7^�^�h�t����y@�J����y-Wwb�c�"�U<+~�h@�>���<�m�=�`���X�u5�CqS��@��ý�t��P��˜�2��۝oN������O ��yk��6OT��2~�6~D��~�Uz\��y�Z(�owX�������!���k�@]�}�F�fF}�g��)�6�{8�\+�س�܊���ML��GZ�spV����qS׫t��ں2�I�R�����g�{�5���0E�zv��_,�K#C�w�5/2=��@��UZ�-�;��/^�^��K���${}�����w���������Z{|0#�*�������s�C�cU�}ϩ��$Wl���Q�;9l���v�}��^X���ep���4�5i@�w�����c�7��n9M"+��rZ)坻�}w�o�h��z/6ϭ�]�Ǘ4N����1:D������v�[L�E�|����"��g;a�g�!���G�4�y�^�׼�}�x1w��+59�@i��N��nu��5w3dtVX�<s��3�G�W��0<"���#&=^����f?@���`�ۤQ2��������@p���r	:���e�7�D�{w�2�>�v�_>D�o�l+�V����x��lð���5�Ѕ�@��h-�~k^��7�y�r�W ί���zdlw��<�OdɅ�POU��.�h�6��u+	m�=�r�%	��i��ؽ��Rw�N*���uޮ������KYū&��k�BryJ��T�[^{R����~�}�4<W�X^n�	�}�f�MK4.�+����3�x� ���7:�f��=��j.fP�
��{�˗+^D��bI�]�- B��d��T�g�9r֬��C�0Я<�;�A��V�x�z�nơJ��L٢���/�-�F����TC�!1�bj1�v�ܣ������h�w)\�踹�[�	���[�X��n2Ԭ����\�I?+nuF�CNw��5�}�����h|���1N�sLɼ�a�Yy!Q���.U���{_`ɞ�vO�����U�r&n/*F�U�/[0��ng�ˋ�\��^����ٜ��׉6ok�s�4���1��{D��7G���R��K�9�%��;�\6�0��r{��ܢď�zO)98,�.��5OߞJ��9����G2���}PO�{9e;��6�팚0�E�Ym�R��b�@<uKrx�/��b�򪇻����A&6SV黜�����ɫ´+��{ݣ�{z�#Wn�u�wv(�۾^;�~G���������$+���HF�e����b��^$&B�i@�6ä顙���\L-��.êu9����&5<�n�N�6�D�V��q뻱���om�#q�G�m���b��^��[���W�~g� ����ډ���5ӈ*�4���k(�QA$��������m5DAE�����p�Utu�EEKMU1S֘�1������DE&��S$�NZ(����1�K�݊���Q���LF�5�c������}u��i�T�S�3�Q�GZJJx�R����w/l�f�z�N�|||||}_v��]OVŰcF��:� ����E5U�m���M4�SUEMA���MTX���Ѩ����Ѧ��&����f��w]LPOF.�Y�/�$��Ğ�3=�TEv��;`�����:눨��i���J(�ۨ65m��+�EAU��ݎi��������WN����])��wE�
:Ӫj��%4�=�ű�i��v��z�Tt�5�6�5݈�������tI5E��8�`�6:;jJH��S��N'C����3y��ߗL��MQ�f�e�D6�3���.� �u?�X1x]��V؍f�S�:�gJ���*k[1Y�
���Qj�����X�\�v��y���B!@�D����D/ <<�7��������)#"��=O���-���"#-�	�v4�oL��<^%�u�s�1�ڙ��/���Q�=�����^���`�}h��͓X&�.CZD�)C�<�L(�.,͙R�ힶ�����蛇�.ʇ����g�"�jd�cdp��C�Bc@�P�[��\�cQ<|x��3��:�~~�S�5��T4J���\<�e�{����~��$�T��wuV�5nV�q4�P7Z�2�+���K#��\�J�s���`E@�w�'q��!{l���]ԛ޳'���49y8yN�uM1����ZË�e��A/tꟛUܳm�l��r��\t4!�C�v�I�δ4x�"�;'-#&��n>�E1=*���\q���Ʀy��k�S��_-��7��3z�lgA@x���u��C'���m���/��1�!�GJƚ/r���vl�6u��6�#�F+�;DS��!�O�D��A���/�Q��g����	߬���8oM����^�:�"+��CI}����~��gA�CW��-0����c���qb�eIʏ����9^n(Ǐ���g_�ݑ^���]�N��}��px��1
H��s���D�Zj �U�¥хcb��L�1{���w��=�Z����=�v�h�3�Z���S���̜�����J���t�4��N���#�������H�*D�Ĕ�2��J�*�-
�R�)@B s���WUn�s�{�i��L�]�Xe(r���)>sͼ4�^Y�X�ihV��14����[��6���ʙA����s��͵iJ�����V�&�9A�-��|i���y�aE��8<󖰚���!� �4?sϢ����	X�^��D�sܕXij��{Q�a��,��q��7c�Qݚ�mз�x/B���gD��=� ��U���'8�ǽ.N�7O�Y�>��8�+��9My���E��"7�휼�On�$��f0�?�A�'�Y�>��3,�z���<[�2�_?k�Q%��T�b����#ry��.s��f��JY��ڞ����Tݽ��2s�~�i�N�J"C�����#�UI��Rr��G��-�Ú�������
0+G����=��+�5�œ��\���YRC*g���0�,�n��LZ~I�����`����#m�����2�D���0+�*H�A8�xd䇆�]j1����
=s��M�zL�{o,^�1n�@�4��y��8��C�v{�����y�d�huP���Lh5�w�)9kZd����ɉ�SEEWd������R:R�x�=�p��HXo-���R!���u����@����=t�R�]��W�C�w�*�%�:��Bs��b��7�K��� 8�=_u���E���!���p{�p�{It���q�;�8*o�t�o�J�\%���o��?���JX�B D��@"�Y��?5Vqr��{�ͩf�zwf9���s	A��ö�/]P��^��lb��SXZ��8�ܖy���X�y}����F}[~��q��O�ੇn�D�.&��^��1
I*=*�FSn.�}f��d�S�%����h8Q���nZ�_DȪ�:���
q1_�� �����^�*��!w�1���m������f��,ŧ���!�>���9��{dK��I����Y݈�釸�40BF:�i�L�a+�nǼ�Fe�f�����@��A�v�z!���h
�ˊ�fY1�{�u��}Fi�m�����p�P,}&1���\����V5P�qG!�JҖ�+��)'7cz�i��-m�����R�n�Ϯ��w��@���a��T����U��B}c��._Bjڳ&�q*��=~�g���':��r����3:
σX�.2�'��j�d�9���B��8s�^�Mj({!�B��<�G�Z�R�*�
jrq�uEë|g�H�ހ��5����d��u7���d�=F�u�6���=��N��B�)I�w�gOd[B�Ӎ����ӕ�z��Z��:�6��9��]+ӓ2z-k�^R������)x�fcK�9;A8��3�x2�u�K9�6t�y]�����OL�������yr�G�c3i�H�գ��ަ�,��y�Q�nQ�ie7�-�o$Κ�G���D0r��(�+t���;ħ�&�e�?��� S��)R�- ��A,�����0 um�8�ݍ7���4�A����H8�(=oZ��5�&*��.��K�~g��B�n�N�[��d�@�0����Ƒ�~�A}�=YVb�k酊*	�d]ax��pk�f���>.����>�^t�ʧ����-��
�a�n�����t�¬�熓`�n�s�29m��:�z@-�ʂ;P��K�4	�|yp��%�&5)��uEs� �P��m����t%Z�sx�n�[n)ʋ
Y�̩T��A�sۇ�p��mn��ni�a1&��޽ ɮ�]U��Cr��B�xX�1�\�iI.`�~�!����2�|�@b~��Y�q]Wu��<�T5K8i/˪Y��m��P6tֽ��f�&a����0ཆr���t�{HkެΊ�\�i�m
wA��0��V���,�@�}��ǲN�o�}1�Qe|��4E@f��N�d|�n�+Tj�As.��μ���E���&{f=��� Q5�&�ct;��Te$`SL��5U�6{������0�������63��2p`=�<��Uga)ر�'�z!C?*�O^�&��S����+W<�H�8N`����L執&�5!��3K�]CQ�KQ����qfv��9]�u��J�؈���~���|N�5�I�9�
��\�˯��}�47 �v1f��8�M:&%����������yXs���c����{�����!J�Z(%B$�� ���]ıQN�.�Z��J8s�p��ךE�ۦ���tS<X@��8���/2�Lq��U�OeU�c�ҪZچ�!VÇ;(2��B��G�>��LwbY��Bmg�i܋[�ꭞ寖9[!#]��blNԷ5{�	M���BeK
Or�hY��{i���ft����X*2����0-e�א�-:�t>C�FvW��T��)��1)Օ)�j��C�v��_���ѓ�_��}���X�ٚ���/�=�L�[�6��#6d�8ıbK㺍����U��GOFF�Q����`{����}����|"�]Q��֑*�r�=�Y�]���Vf�*�9O?4Z�K�-�uC*1��;�׀�� ���:nΩ�Ln�2��؈YyG/���ok{��:P�^*�8�Jz��}d
�Ƃ�P�Ʉ8{;�XG�:ml�K1�c��-�g �O-�1<��N0-^Nо*L:��sJ�砲4����ݐDջ>�0�4���e�����'�p*`PaQ��%����i��˒�m\L�{���ߕ�2��m0^���}T��:�$f�N�_�Ԓa7���Fp�u�ש��s��s�����o.�Q�-�E7�H�g�0�J����0Ώ��&��ӑ�c��ow�HB�LR���9I��p�ݨ�/T��DMي���;;��:�e�n�7�����������?_~??u�����)��"A(�A� "
)dB���&��;��������G@t'�z��HɆmǡ��l�)LK(�}�L�q�w�5��J�:P����G��rY��X�<2.��t^��_��2~݀ͺ;%�N[ʼw}WK����z�B�^|p<��~��}�.�1aCC�p��綣5ք56�*�s�����(Z���B0�z�$@"I5�}������hAiidh��r�{���ߍ����f�����ۿN������;$I`{�m(�N��"���ޢ������؜�R'}�Hx�d�-1��.Tz��Sw��l���[�u�r3g��h��׫�ĶЩ��=�W�;=�sΠ�S�y����.=<(	U��دN��,�A�P�������;7����c�<�Q�����g-��5��<A��'���Hyղ����D �Pνr�y8�-_Tg-k�^IM2�e5w�F��W=���S܈���Ivl�0�ƐF�1����}ڳ�{�U�ۥ)��'���j�)��&�}������� �5���mǒ[/�qgzr73�e�i�����pj�Q���MX7J����&�6o��q�>މg���t*��wx}��������,�����>�I�t�ӓ��6�q�{�:#�Uѣ��CVI���u�]����nƍ�-��wI~��"?��@�U�� �Z�
��~��~����e=[:�7Y�`~�'z�$��1I��yh-�Ú�<������a��vL�����bN�=�X����y�Vc9�S"�&�r^��!<�^��#�.�`�Z�Y�+��6�v�+{e(0�a�O�bq��ǟ:�i��Us]�^@P���w��bA�l�l_%Ө���dȂ���\&�yft!���!�9U�B�ՃR)�5�w��I��nJ(́�C&�i�{ ����sݷ�|�. ��ͺ��� ��(K�:O^5_h�i*x���ա-���^�nq���z�	�^��O�nLW5x����}�!ۤt0m��D&-0��]�5GWxC
�¥��e�oD���h~CQ�꼶�pm��a@� ��jhOr�|��/"9���;�5F�^�|��UV������ܬwPny;��Q3Eڼ|e��.hL�rzLVMuJU�3/�='���Gׂ!�Ƹ�EՎ���s��}̳L�[�K���a�c��7VmT����#�e7�g�gmYЬd�EexY�!�)�{W>����^�	rd�7�����DDld}0z���TMى��A�1NJ��M�VU�������B;�/C��f��^Ma��t�ZW��r�zc�3��޾߱�^+}΅Ժl�B|fU������wtճ��	z�}�j�b�T���i�����)ø
���#S�92\م8���� "hT��b�Z�
��͗Ws�	)��A���6q�S:|�\<�
Έ����¦n\17F�b_����󔨬p����R��.�	�,�,k�uk=x�c�VT\9����(>�\ezbyۦj!g5z9)���Gc��_Hl��E:���C�e�|b��Z�R�*�
jrq�uEë|g��_��=N����7��֭s���O�-���a�-�]�'��%:)H�D�IžŰ��жnyёt���)�|�����77isyy
�>�(8�6aU�.��b8=��T�`/1\�$����9H�پ����j�7:��\����N��i�!?WT�׎��T*��}R�͂f�B:�*zҜ��6�^4�\sC��+�92���5�-y�!���:���5�lY�V�aF�n�6��z���Q��]o�\��iIcH�C	O�ݎ��u���p���+���`���kĨ5�J�yX����q�q3��kJ�[0�'��\��$s����2?1f��IwNt2kW�zu�4�\)�mȶ4uP�j%k�f�1�\��^��]Bu����z��h?����GzN#�Rv�����sǨ��ޤgTQ��������o`�E�����w:���~蒍�跏,_��&��Q�o9��t�Π�-��i�_�&/��Z}��(��[�o,���iR1m�j�ыp<L���hn�4���W
��ǜ�^`��>?�>��3�V� �������_�ߟ���Ʀg^f��oH��?VԳ-��E�5�P!tN>�a�r�&����/\�U6�Lv׎*�4z���\�T�w�h�A`��o�2��'W�,� �,8�ba���#]�>�u����oa�eߪ<Э�c V*%ͩ���èZzH7�00l��#���#2,��OMMm�	Y�c���B��|,��!m�C�9�W�Q˼"�B�:v*�
ޑb��zw��,��Q�8�V9�Wb�1Ϛ����<29��B#^i�ظM鋇\��c����MTy�񙻤G>\N��B�9��r����q����W�̡Fң���.b�͋ٶuL�����)��-_gSF��)�	��lǷoQ�nW;R���%6q���P��%vл���|~�6u��w9�?<|�myl�xzv&(p�lJq(>P!#��CH�S�^�BSc�	�i:�.cojZ�>u�m������ܑ2͍��iN(�zpl��$lP.�|�� ���ƀD��锝vnor�pӮ��q�t��,l��x�4���5�����s�����c�`��c@/�c'��ꅲ'6G(Q��N�O��/ۯ>�/v��i��G�)��,O7i��"J�x�NDc������`��*�r���xMT��׳OR��s2�MOD�}3`���ĺ����%*�S1"Ii��&ܩ�SY1��IK߰���Lŭəp�޼��9�HCt�"��؏��@�!@�)J4)�f��m��W\�g#��兣R���cKMCs
�~�-^w��<P͍>����ٶ]2�:�Wt�]r܆��J��./
�{"���]*��qr'��[�s���C�.*�e�ͨ5A�QB#1)Κ�`Z���/��VGs��#�ո�`LS�X���1��Uޚ�� �[�S�Z�f%�t�jd`�0��:��A/t�+�l���xuG�/����3Z����Q� #��;k��vm��Λd�˪Ll2��܌�/��<���Ƀ\;�`ӎ��e�Ľv=�"$1�&��tة�'�\ǥ�@��X�EDje������8�`6��r�(�����8�z|0��!ٺE�<�"!,45��6_�P�&��5D����������/XCP�C�OL76
p@fP�Y�-,Tv�!�.�I�S���OH~1�r���w��8%�������e(r��o&���CA�O���+��\��Z�5�����%ߴ��
�::�,UO��{rlS5ES6��A�S�RG)��Q�R��Օ�F��;��b���ڌ�J��n����}߁�:[�޺��
�Vy�R��aL
6����"�ê�M^dR��lf�n�-63[�w�iN��d�������x�G����N���m��E�	v��u)8�\z���z����sv�n�"�+���M�$�(�h�+�T��kc�ܟr��z����ү�Bb&�c��.�Å��v^�֏�ģ���N��~�H+t�͞��y�q��r��k����	�0v	����a����w�톙<����"1�|yy{ޝ�����ݞ��^n�ᠧ���mj4N����l��Fb�ݧ1b�;�����v�iP���4�ڃ��ѸyD��)��y�oh�w�<��F�y��O�l�PNaq^��~�>���p�N����N~J���x�>¹�9}���lڳ`��x�u���L�9��>�t/�u����\)6�{غ�k��B��������(�<b8#���z(���$	�ܽr�g}�mћ~M푭���:`2]�tY&��'qn��6��*DK)�;�Jz�{5��<���1$Ǥ+4�T��F%�u<Vl1F�lމ��ML�M�8�D���<�m��l�oS��,�J ��<�bc�=�
'��Ί
���o��Z�����U�PJ��s�S3�P�TT]�����>����t�Ɩ���{�t1�
�rPոe9&���+>�r�nN�:��%����w	�>�"Po�<�w�d�=3�d
}���r����b9����OR+l�X��߳�q����+���wc�ȓH˺N���QLV]+U3N�-�3F��GA��J�ܷ��".�*��J�'�cW�y�`o�n�l�ͣ��E���ׇ-��N��s�	Ѽ���d�F7�5n�D��;���Ϸ� P�4g��G���>��Gk��N9qӘ��&N+���r̨��ʙj7�F�i�c��B�!�ݝ�e�,�-[�6Uc:�5��PF�6��.��7�}۴`��z���X3<V�gJN!9U@��b�]²EZ������xћ���$1��֏�N��
���I�7�vDS��o5�^��B=��.єԋ& ��n���:��6E�@�����hj�ɖ�&���^4Sw���u^��\�S��{��g$��/L3/�h��������ޙ���Gs}��u������v��|ͳZ&~"�1r^�44�0e2M�Չ��vJ�ܫ�9R��ډj�v3^w�KZ��F�N�5s�X���n�k��N�<��jӝ��P��.պ@S& �/�ŕ�4��𽚑���xf�H�F��u0�M�!��PS8�e�Q��g�d}�މ���iw�y\U9��:���w?2ȗ4�4����"u��1U�1uh�k7:ն(�N��\U�^ˁ8��Ì��1�Q�!�#M�4ݝ�Mhr���
��Bmm�撵]�b�*��@�{�c^�_���������z1TD_�A[b�()i�J��J�����h�(�����~��>>�D�gTQ�M�Pi�]h֎ڛY�.ä�f����:�11����<|||||���;Վ�i��T��;f�n�i���m�(��]h-b��E֊�GGA������cm����GZ����j:�u��U�HUQu�F����AE�q����>>!Ӷ�s�׮=`�(���ƣES�Ŷ��h�b��:"ib4�uѪv�]t������ш��h�T�lTcջ�[;b����v��n�1 �N���F( kN���*��D]�q6�\EQ2��;��&])�(�h���]&{��6�lS�ɉ�aѠ�@h�4A�;���;�Gl�QƬd�MS��j"*kZ"J(��U�����bclhر��$��  � 1"�����G�)�KW�x��9[-��*a�M̧�H���ܫٓ�NI���+W�*��o}[~�>���~���~�w�S� I��"� `ěؖ���ڜq��bK��M5"$�t�w�Xqm�����p�J�`������%62e�բD����z��L7�F}~��Ή��ɯI���1�D�����:��#Ukb�����i����:�~aϢ�\/N����X�i5؏F��sS:yjw�\Zx.�fa0J5kN3A�ʣS���s��!�)=tD�I�9�N�)ƒT���ry������C�#a!�I�uY���*g`37Jf(]I�-�`d�q�*R~b����٦�ǣן#Ϣ����wjȝ�s�H�ݠ��B�z<-�+�PCuv�5':���jzŧ�.|�M�~���Y�+����m�\�{�4g��\�pƀ`�Za��\�n�v��0�� V@�R�:ngDSnJ���r���g�\�V"���<��{���B�՚�Lhɬk�K�X�3Z�suМ���_�r2���W>�*��8>U�1
¨#���_L�)�I)���4�i
�U�V�����L8'Q�+����Z/�gK�?;0ފ��'���L��'���*$���l���ȱ�m	�K}	6�ep�L�̊��2&�rY�
M`ڔp-�84�����# Ng�����4�?��G��G���vv���/Yo�;�sG��{G=F,8$�嘆�eN�+#
��PjV�	Z�� _!�P��a�rM����\����%�JH��X�S����?�_���2%sL��P���U㲓�YX5l,(r�6�t����F	��~�����]z�M���n�83�TkO�ac������u�w:�P&h�Ŵ�0��z.�D2*�ץ��Xe�
k������H��FBg���F_�.q�{z} fY�h��%ب�A�.�,�\bܿ��0�s���Iv^�ִ�5��:�ȧx��L�#G��ȼ�G��m�ء ��$�k3�EY���..��^�<)����Y�¬ǰ�l��sӼX03���|Ǧ&nA=x`�]��#�x��}Jq?(��*-l ���Ƃ]Z�@�|l��s�\d��b$�ɵ�� �l��8�6d��j1�̇� ��C,{��@Z�R2�����8�/P�=q����I�����g�l�V��>�� ��S��;%75�L�ߜħW�W*�qw8b㚘EWRԲ绝SE����i�F��=�v!��0ӽJ�"���Qw=�����1]l)��=
���}�|칈95Q�\8Q����x�Aθ�F�*�9U)<��l����́{���<�(^N7&����9v=�T��)��+3z�{��7�1�]����	�8�P�淕�s�B�ǖ\~��u���4[ǯ�J�v��RИw;}�<p�;7qt�-��VJb̞��O�%��=�D�7�q,[o߫u�_��LJD�+7�=��F�����Se=��iiy�[�&\K�'b���)��ܻ�����B�l�n1�l3���޻��	K�s�,�I�RX�GjO�û4�|y$¸�w�P�>�/���G�S�֭W��\�9ٹy��/qTXPY�̪Ƿ��$J�s�&�r D������uu�X��<�T4�u�	�����4-XQ+\���\�QzhO�Ȍe�a߬���&�"��5�CgY��3pNZ�HhE�f�w�h�棩P6;�:;�"��po�����OU�ڑ���Q][�g���(!0�<F�zv�=���q�#�꾘B˗4�o+'M���M���.���Ls�����+*o�BГ�~��I��(ǹ��D
wql����3��-F�F�S��[!�#Hz@A�0��U�6�ƀ����B,��̔���_��ʦ����O]U��Q.[��/fG�����B�ךn6�5t�ê�x����w��Pe���n��<t���x�@̣k;���a@8���,�o�Q�Czq�ܰ����\������4@�hdn�D��� �$�/2»�3tHb��ZĚ�q���	~��󽷐RqŌ{���x�����=Ոd� �i�zr�P�kt����H�=k	�T���l��q�L���
����F0K�'2�=9{l�����b��OG$�Li��f�����;�^��(g��G7��p��C�������=Rū��M�8�L�ҡ���3�^"�_�ݡ�>�R5�SJ����z��V����bذ�2`$;'�1uQj0Jca�Ju�X�b	̈�:���W��?8����&p)Fi�}�fbC����t��4�"T8�hv�jjqƍ�3	۹彼�q��{�P	�X�\�,y#I�k�8j�����3c�`��uAf��rUx�%��ȳr�Cȵ]0��J.���<�P�F:��;�SR'"��� ���9�����|J'�pR�eHL�-�l��*���~n*�C�&�p��A�V����Ov6n��|S�L�7l���S�QӴ/��s���R���@p��4��*��}y�7cʄ�f����lz:��ښmW�E���8Î����2w��k&�k���t�k�����0g����d�s���f�8R�1��=N���Tj�rp�ӭ����x��q�©ڀ=r�k�,3������x���ξ��d�`PW̠���u;n����Vp���~����R��x_T�R5<�t�4T����eV*&�:�L9k+Xѻ;e6��la|��Gx*=q���Ӥ�j{^����Ϸ��d�����\���pN�$����Ky�w+&�d�[
��{�B�>��`������o};|�P��)IՀ���"��W�Q�6Ũ��.�4���}�3c��WS��B��j�tTb~$�bwk;Ot�$@"|I�i�[�@؊���gۛ��a�c�7u]ef�{�6�_�;���;ż
/�dEg��@�	e(r��}y6��Y��Ʈ�=]�l��ܣZ�>@3.H���6T�y�ɛmIK6�ыdɯ��tK�q��֣��niE��kw��^>�3���:E;���"����	X����O��
�����ۣ��zX���P��v']	&q��ǯ[ռ�[� �dુ�T<=�N��Z�=䬲�y,��V�(�5��Y'���+�&���|j�Ξi���%D�f��w�0ݦG��9��p�gOT��X�a��8ꯥ'b�j�LRR����[��\:�����uF���7��c<$���վ���%4��p�ƶ�|s���F�[��j���x,@���K��v�����#���Cl�O�ض��Ḋ�7	�=���	���	v��\�`�DY�&�N�`��F�vg0�[͠���b9��N��Qr�sä]�Q��o���iXS�=���7oj�}�����57���E�t>҇m��+�{�x/M:�ݺ2n�����5�3�U0��O�{���*�S�u�������{���1��@DMD��nݩ$���B���rp��HeFO��{�C�yC^������)�N�=�f�6�cꭹ�r�.�AOI��t���!��!�:|���}���0c�uи�5�V������ڒG��6�*k@��i�oV�}
�Y�^��;�L@p��>���>�+��(��,�պbj��4?-F���p/���'�նr+gK�?Xx*aۨ(K����P��ќ�Ή<�T4��Ƚ�b�]������K$@9C�W5x�s��X`�±'pu���cܤ�CN3��F&���-XQؕ�S�5�&��}�������~Kzn��u}Mb8����RB�m�jk�!�4{E�1��ua�[<Cw�w�"���g������Z��}N���\}�<�똰6Tk�o^_����."�� =Ų/b���׻����wm��1�~������Q��W��A�y#8�^͜eY��χ=;�.3���o,G#$r2�C����r��q�J����O�u�n71�����[ۇ��k�"C�	����3[ԍ��S�@�����a�F_gyb����w��M��$mwk�!-�%��5���c^��Q��nH�ʎ�.T��[���3����c��y�*�<5�e��1ySl�/�|���f�V���B[�`�<f��'����n��W�Qͱ���3�T���x�G��Z�08�>��۴���-Q�y��V�8�'KT���W0�AfN7K�:����xۦ;�F�ff����� ��z�K5צ;O�%ۄ�Jnj!2Oa�JtQ�J�#4<�:��q�}�ź�H�GR�P<3�m�N7�HB1���a�e��7�f}�J�,/1N+fm��.���n����"e�(�
� kSߝ�Od��#a�O�:�^�;YS�/�#a���"N^��W�л^V��)��9�i{ �x�ˉsbD�W��)���p��E����f�DR�p�["w���cz�]���9Ԅ�I�P�+��\��T!v]@�ޚ��fd�ȓ
�O��q�M8����n���샭(X�/<���K���⨰��<ʭ]k	�{����n=�7#�.����x������nLW�=6��An�~��dR��V��zW=����*9��u	ֲ�:�>$��f��v7&@~Bd�mO�
\H���,��&���8��^e�Z�4^4�0�r~כ����'���S]�����ȗx�`>��b�l��q��~n��9�-1n�)�2�NB�r&���<�"z�m0��4	�>�HoW�(��H7�e�ws]����z6�;�q�kD�}�5���؁�ʃ�1���=~�U.��$n�Ex�h���3/Lɻ�e-vN<}a���*�6��!�NĖzx��\7�`�V���K��|&����cOj�o��f8�L�4��-�tg/>י��3��6^��>�����dx�{;�ddQ����e͜������	�Hz	@A�0��T:&���fq���FS��eϯ=I�ʪ��&�O:Qi��cĤ��v9����r5曍�M����f���e�����--��$�����{i[�ʖ���d-{;2��(Q��g9�'f�ٳ2����_�m��C�ql>�~`�Z��C��lQ��zv�����)��	�J�'�yR�������я�2�DϷ^���}Ol�AE��@|�0�b�CP�Sm]Jc�n�'jV)�u���e���q�zIJ`��"�]���z��	�[�Hqm:A�]�bG�g�������ZSD�V���ٕ��<K$�<SH�a^}���a=k�@�a��Ⱥ�(��]�3J������A�bi���<��):ahԢ��-5��\��p��=C�:YuS+�𥞒τ��
=Z+б厃Gr���P�Y�����O�~*]*���K����[^4j����+���q������e���h����V��?U}���>ڢMU'��C���6�"ʱns]z�5�M�(5���y��xϻ_��.�v��M�5cq��˘P���t�#Y{#XV�[��rU�8���5Y6-}�VV��Zj�9L#���ƘB5��zK�58�� t��8�0�Gs��T;�nں7��T�:�#l�f��!��Ӈ�PB����u���4ںd�2�*��xq�\��+���_,���M�ė�ݑ�7w->����	�/�b���FV�C����՘x�F+�ph�_�?����S�>ߑ�N=3<�z嘗�������}��F�����v+MU�G;�jm��6s����HfRO�c�C�"���:"��qa���K����c�L�s/_��]�m�����{�҉�ia�0��	�"h1m�G�6~��VT�1-�_zrΔz��eK�ivD�xW�㇥A���K��9ɼ
=q�7����K�}��69�p���SݢS�o6��7�SD��iiL��.th��z��fڇ$�þ��A�����Є��~�iۖ}p2<=�8' ��:��*�)�k����8_�����K��l�|g�*�Sr�w��!�x3��-)���[�tf=z�����q}�%�Ȉ�~KJ���*���1�/^�F�
�v%��n��:	SWz�OG =
x<��������Oj��@�����uoO1n�ɮ>ۜ�hԟ�����p�������ا��I�>�nA�q�q�=��U���P�)�J��wA)R���B��ѽ�'��x?Y���k���W�b��=���n.�!ɟ�~�bY'�R�er�&�a����l��Sۼ	
���Y���m��+���8���'��DJt�ħZ�K	*Ml�qͣϑp�d<��e��oWr��-y!P͍ BR��Ԡ��;��q;ԩ'�1I��yh�XsL�;:ُV��+Wa޻��].�ǟg��[`i��z�M���C�{�
ָ{:�E�mODŧ���K�a���[/����M�g�w�C@<��<�)��
=�"�q#f%�=�d�={ѳ�����ݺ�S�8��gĥ������%VE�'�q�b]�c<
�Pw�	n`]Tt�wb���z�J�4�̓�ʶ��nAJ�k��Jrִɷ�W>����+b�ٶF�pt4q+�۵�ny@� �9u�u��K�u���:�Z�(�é�k-{'�ն$�sQ~��[�S�u+5}��ﴯ�G�h��mi�^����v���NF��t1�Нf9����<i,��ܸ;�gg@h�o;BLL,ss�{��yb����u�|1�
��{|�r�YS�.��6���nڡ���믓����ozʘ�շ�ۧ.R���y
wKɸ�r�\C�ĦԜ��C�)B�w�[����h��r'���o���S�Q5��>��^��Kؾ��3ä��!`����=�IVY\��v�#m�`v�x3Dˇ�������{ӻ=�N����pZ��������gx�z;4�3�R���=����-��I��Ǫ����y۞�-�p�~�>c�t��:��7i���C�ұ��n	e;���2�qҹ���$�yon_P3�Ζ�����]�,{Tρ������9e��{������Q>4Pj7������ž�p�F�R�E�wv�۸���{�9�\]��[�xo�E3;x���!F�᧱�6-�7^:�>'F\\�N<���7޽<���=1�f^����,�\�A��O �7ݞ���9��4��}..�`�K oU�^�����$�@ZWg�����F�.�W���-�e׸���5���zl���9�7w$�O��΃{i��K�3��v�`@��8�Zp��~N`��&�ż���FO��������^�ї8�w��@�O�O2�>�3���ǡ �����y�s���'���Z(-:q�N�-�5gsM֪I��hw����W��;���]P�޸��&7<_g"|��%�7�&�snh�Ew�׶�~�`s����{���{�5���5Ɂ�1�1�ufHI��`sQ���9�v�/K���qh%�����K���a�fy�˕4�S4�qB�*���\,Kw���k��l����9�k���5ƈz�~.;��<�L,���s h�L��z��1���^co�����eD6��P�^��
UM�2b"bщ������zzxmX��߼�R���G�K��Ew&��R��}S7}��ŭ��۫H������ ��x��'��&�7=�5Pƿw����[呩
�nnڪz�M�		��79i��E�Z�j^ӣ^��$�(�����/%j�C6�F ���z�q��	��Ƙ5Lz��I*��}���nmg����#��	����2���gӋg�ag����ώ�І�"�zW.��"����s�>���D|�yf~��̰���������=�s�D
�����^[P��P��f����L����]��x����;�d(!��Ed<�Z̈�[���(UÏN��F����:�G��4{p۲Y�ɴ[��w&C����WJ�:��[����-�kޯ�'�p��K'�9E��S����tl��`ʹp�໧������^�{���ud����x%��NzWW�|K��W5�/ӽ�w[5�����e&�T��Ҷʆ��xũ{w-f���*��^���ܮ�wz�ds���ޒ��д�4,���4�^U�12���+l�s$nn�%$�J3f�F�U���c-��z����F[$/�
� ���İI%�c
�`
k 8~؟���c�AEZ�ɩ��lIER�[Q�QG��vv-m�*��?g�>>>>�f"э�V��lF�4Q3EUQT�$8Ϊ�i�����1�Q[|||~�����CUm`�;cb6&�N��"-�U�cF**�6��}b��(1�����񱠩�(֒v�Em��"��i�j�m8�
�mj����4�j>>>>>>o�1Fō%N�m11��"bŢ�i(�*�gUQẔ1AF�������`���61Z�щ(4:B����lP]�حhqb4h��l�[I���U�h()#�DQIBVͳ%U'F��5�e��������S8�_9�EHEm�ԐRUDDS������P[4��ꨊ��E�SAZ5�Έ�U�"-j�c&�DD5�cZ
5�������~���?����3ѩ���v���[s�π��fR丙J*��P�.յ�Nl�	�ϻ:�){��i��z3�OG��p UD�}��o�}��/��"'� ��i�.���m���	:�:�m�wO�,�ExWd��~�%�?:��uz����Bu,���={�m��	w���t�w������W�k�-��4Q$�a�|�Z�b���:��l��Fq���8ʲ���zw�\fI��>�G�R��û'��\*�
gd�NG�[P]'�:�'!d	o�]Z�_��^���	ڻ�x/YC�{j��g[FV�E��ƻXgX��\��2Ǳ�):��P�
K	mr�9�&�c�7^o��M6�����bj�&�(R�u0���K�	����D&Iؼ'Ev�lNC�N�a����5�
Zq��E�*���zA��q{0C*�d�Xg��fF�*L��8k��v�].��߷�'y�E�M�7@ٓ[/N�o$n@���b�O�0/��,���4k�\I�1�uSf��M�G���f�Y��9�-/#h��=~g�m8N6&\��t���iWGR�]�{u�Ӕ:��+;E�W��\���)=X*K��TD��33�dI�,����}Ƒ����|�!��k�u>[ty�o���z�J��bb���zE^]u�����Z�{^�qw���:j�.@��b�`k���xg�co�j����=0����lݱS�:���2����sA^m�G0�������5�P������k��m�:�	m� S$��QI͚�lĝqv8�,(Z��Sc��XH	���sS��/�ȁ����sovS�u����zn�&,�9e�R9��i�jZ��[����П�>rf���m�Y�7s{)soeXV�[�w���`�G���lsH����R̶�h��u*�tַּ\��b��-Lmn��Z�T��w@���g2�w���x�	�;�X�T�$��t�q�ʀ�JȎ�6�G�h��ْ���ޫs	�c�C��4��cC�[9y�����*��(�ة�I�P�4ZW�g�a�R��]�Q�6�ʙ�Ȳ(wH$=� ҏ]E����MG)��s_I,��/&U��Λ:���ت�Ƕ�{k�D<1��p�9�M�ۦ���uIǩ���5�s��kowT3���=�8��I�1�ߧ*Zڇr��kY�A���'R�����Z��]ݵ+�T�C�yg�#�:k�9�F)�J�j[���D����!2֞���on#Z�� �h��7JYB���cռ55���b�|�I��!���COb�k��`���]И��ކM��RD4D�3b�C,�1�^F��,Uh!��J�ڝ�4VSj�k�sgh͜�N>�vD�V���^��qq�L�0��Z���{]d�[�V�zq�Le���8������+Bb#G})�6��R{�L3����B�����_�T�]���C�g�MZ�ZR�&��~��������Cd܃ކ�'���f��؇1��W^���!�rU�Q:�(S2N��e@�I�؋��r�W��C�.ͷ$�,�o�[���չٯH���*e@-iNJ��yN��<�{�)�������-A�R��R9j��#/�H���)h�G���&5�!1��B�����YS��E�沠��J��ߋ�[�B�νQ�o�܁p����<�����"5�f%:3��c�Ӵ.��Q�X�Ϋy�0��պP�޿g��Qa�H��#�T�@��8u�k�SM�������V�ɹjq��o��9j���
{���9���Y����.݈?	�/�A��>�W�s�U
����b��l¶�s��)TX��O;�������3�G�Y����Lg��C��^�5�DML]��Δ��eO=S��d�[��@��D�_�Ǥ��H�r��:"��{t`�c/�i���2}u5ۺʖ50<<%)W׾�{i���4��ci�C�$@"I5 ��v�ry1Tv�qu��dH�w��y���%�r-��̢�Qۛ�;uj`ҫ�wz�r""�o�6�q�L������r�4�PMf�TX��Qљ�c#�4 �\�P�#k�o)\<y6�9�����r�
��U�N=�=�4��ڃ���1���
^��ȉ��(}�&�kp����e���C�C��ڙ'�z��=�5�۸i�(vI`h%�,!Kغn�Sh����"��M�&D���N"�A�ł�/����?��kV����~=�F�IS6�]L1U+TT�1f�i�ӣ9Hm@��j$���6�i�gH�x���/΋�\zxUҸ`�]��#Ra3]WOyc[u9��9fu�y{��Ƶ��2j��{��
=�Cׂ/K���x(dU�޸���=Rd�g�����	��ֺA�y��Z qyeO�S�2�(�k������l������]4[*��'7�vvEht4�f�'Иt��� E��tD�Iؼ'GT�c^IRkk�z!ĭ�wv׻P�tx���n}�;�(��P�m>�e�h��ʁ�v
|rT8��T��b�+Kȵ��WCp���s\�W���T׼�1C�0g�G���@r!6צ86Ϸ'��g:����w���."�_{p��'q�vYo�gw��/R�@~��-��}k���Ƚ�ɦ"��j�s��r��$��v�+jG���5���A>;��Fi�-�D��@��)��Lz_V��H����_S�S2F\s��Uӹ��LY����q*��!�6c���cݎ`�����o�"z#A�O��u'u�9{^o��ow��|7�'�P���XbR$a��D�VX����b��5T�mm�H�n1�DhqV	���rȼ�����D�C*b""*]���ڰ��k*��5�N~�iʽ�k�zRrִɷ�\���l��n��;�~a�+�UG:��e�9l��Їjt^�:���i�K�Ja��5�����ۓѝ/D�oL=w�q��Q����u����_Z`�53�r��6s�Q�/��C����~df����N�heOWe�j�lk������KD�	������ ��d�wPny;�B(4]�K������7\�^-�}��z�y�[�]b)�l�w� ���i):Ω�[<[��G�j��7q����'z"��wd�� ܌;m����y��CdS��B1�=Ų/8�,Jz'����OeU����
�Ƭ�(88�2nJ�Ra(h33y����(?���s��rnP}jA�T]Z�;Ւ{�iЇ6�
��Lk�6��'ְvN��1ЗV���{l�Q��$ϽJ�
�7��˶n����2B�D댡1<�5�=����
C:Ǒ�):��P�bU�Ѯ�p�q�v����)�z�?le�T�m��J>�0�w0����v�%77;�I�2%����=V|�J��U��A:������o3��7��ڀY����;;Փ��k�z�&n�D	��	����1��ط񻗼���C.�c�zQ�D�5�y�:T�k��@��#����{��e�5j�����U�H��5gv���lD`w1X�T��ΌNM�{�9zyW5��\����7iY�"٬7��c��#D:A��l���]�i�3y���z�_���aLy�o�W6 �d��H����qӅ��-ᄍ�A��p�c;���8@��X��M������Z۝/�7i3�j���&m�u��sO�����\��#�9��9�m���>���W�u��]{*):��(Q��L*�-薃�)=_��Ƽ��0��٣ÍI����k�;|��H�g	��'"��	�=��uf��,ى:��qTXW�0��Uj�|�@ИF`~h���K�v=XNӧ�3f�or��.3�~e,2i&=09�{MV�V��cҹ�(%�Ms�VN��[��X��<�Z�؉���Нj�=�u=��4��0�jY���a��:�z��.������qO>�f�C�KsW�@���g2d	w�\=h���m�^T�$�R�e�Z�i6��i�m8�ɘ�J���0����1���@�r�.���:�4�>�5�i�[��Z;���=0Y7)��I�a>݌A��� �<Xd�3"�E��xc�`3g�����@Ų�3S[1�UymTs��'���[��a�"ʐ�Q3;6�k��_'�7��y�G#��y� h}��`�.�W�)���C����m��4������f]��rbK�V4,vN�{�y��{�j�:��q����7�Xҫ
^��
͈U`����Ӝ�N���R<(ɾsy��v�Q��<6��� ���{��5�Ӧ�ʦ��<T�{r�F�0Ϝ���M���)���{�Hw4^�*��8m�cT��=���*��(�����u�VB��z6:�T�J���eJ��"k�t"��EH�0}�K�j[���M�N���pP��Q]���:��Tl|��c�������8�٦�x���[HN$�P�		���%��N�������ڪ�OWn�h��d�	�6�%:*���b2s����z��;�amA:A�vq���,!�<�\Q\�u�!C��8��g�锝ax�I�s�1��i����p�Q	�s�7�ܗld����r�>�Y�DS�Cji�h~���M���zs��<~sY��V�C�$6c!��
���sܻ���r]�c.
��-����B���*ʞ��r-?5���������ݵw��{���=�.%���@���-�1B1����]_�N0,t���Q��i����#�{��OY�I{�]@���9�K��q��a��`�|�cji�X���5�O5Ӽ��Y�G+=�ʍ�뚽���/]V�AF��2�c�a�4�h��Fi��N9�+.\e�L$�z-o�/v~���P�ԩ����9��@����\b[K�ݵ�\���%��wFF��;DY���"�s�jhژR]g��m}���n-޽Pݽ��|*O:NK�?{iǷ쨄@u�%�v D�	�L�k��nr�(����Q������z)�
U&!?K�1�#��5x��1/A��pͼMr7�b�b�M��P]N����P����!�Gb=^c�A ގ1��3��ƛe?_I3�u7m�-G��ټJ�øvM��<$ �>2�gV3~���n$��a{�Y;f���siWM��nFe����ˎ<�Ks6�wkez���]X໢3|1�l���g���!(w=�'���r�
�X	f����Փ��k��spi�3FҠQƑ�Jniԍ�{�փ1��s��;l)���;�9e\��i2��O"�%4���֫ǳ��y�k�
�0�V]@�\�kak��.V�?P�Ya��~��aM���)W��*��P�s���ZZD؈h��.����p����)O���ٯ	�p*��y$���ED��ћp�m����d�}|3Z+ϑʞ�W���y�V���sT��J��jؽ������g�f��]��t� !">�.��K@���K,��Mf���B�i�J��c�\0�m��3��ogvsx�whY*��2̑�NL�PD�L�\��0.�L��t��r���ƽ�<~�~���Co�<cm9�����W���eT�Ҟ�\�s���p\���=b	�@����S
��}��OE9D�u�˔���5G���K�]+�x�P7��M	��1G��z�vb����9�yx��'����h���~��`��lA=���_uW��CDi��)O(��r#waO#*���W�wT���*���-�Oza�R�Ä��n7�;�V�p�OH쑸i+�ň�[rc����y�ٵeB=�,����DW��-���:'ս"�Gam8�s�D���lV�檏�b�᎚�o�݈���A��>�"�/y��s£Y��4{p�o�z�w�3��%Ή="ͻh���+7�[��V*�ۛ�̞�<��Q8� ���#O5-��T �`0��7��UT���?߅k$��u]?�Q/=�)����|���[�ٔ[�jۿ<��;��v78bL�����B�7�Ղr\3rT�F��q6�/Y���"&swb����]%1�i�E�У�,!;��d$\[jkn!D�������DeT�����pdx��"�7�����Vv�ш�s\�%.���Sj�H��5n����(���&��b�	��>�֜h�Rx���A�RR�m=w� ��b[\g������;����ɐ!d�b�gb4b���PM\`J7�FH�i˚چ�6����Q����q6�'כtyA1�/v1ֻY��h��eg�ֳ��n�#���}���ْw����hH#!�������he�g)��f޺磷\w��&����
:p�¬sɐ���w�nO#������ؾ247��U^�׸q����᥺	#eJ���(��>�����U�B���i�G�R�1�x����,#�@��h��W��W9��h+��:С��\��u����Z�3�y�f'{e�����K�t�*3th��ʖ�n�Q��ENڙפN��EM�m|2quG�o0(����I��{P���͌���5T$��5���������N�wX��cX�&��'i�=�=����:��o�V�r��;"Aݕ2�{���>G;�&�2���g|rR���O�nj����Iw`O ���Jy�Q���_�$=:�xˋ���T���s��<ϺW!r�N�yhs��˼�n�/]7~[�u�����>DϮ�VžZ���M�]n�E�RϮ룣����Z�V��է�RX�3���/��(9�|�>b)������ુ�+�����G����4߾��[��Lj���E�<&����^9���N�bb��ƛ�ȺxIG0c�U8�.J���)
dJ�FED����JVRpa�7�f0��J�y���'��(>1a��f�Owɝ�m�ܻ$N� ��R��]#��t;"@	�l1\�{ӳb��|AZ1Nw�{�Xˉ��f��&���$���E�3���_����W_+U���� �*Ξ������{��rۢ|J��P����5����}�<m5yyd�0�n\�Wy��^����-��߆�5�h͞�N����K��x��UǑm��7z��r�T4��`��n����ś�=oI�,��>�z�D1�t~娔r��컼��Z�Cӟ����{e�wn_x=d9p������K]�X{����6(��s���D�г����9�Q�w�0�1i~KV�yL���l��{n���ͻP���M�>A�m���Y��b!n�����x=���άU��5ENˇ�x�/@��O?7<3��C���O8aҮ�59��6����&�EE���7��R��\�{=j�!�	^,�G���.��Z�{�#v��g.k��Ut���<v��:���H���o��g��L}�\<��a^�}�W�8x�:sm�a&��N,y%fI�х%e%�q���^
��9U�l>^������Oڝ��U�/`PSW�h��b�3�ھ0{g��E�RD�x����E3rb�	4�*H�yP�i6�vci?5�WO��u�f�T��� �Ɓ\��\DT��Q�P�hٝͦ�؝�=ٻaH�~�wB��XA:��>�ή���u5y�#ˋ51������F��V{��J���{J���y�N;�>��o��e����|!*(��8+��x;�ǹ��!Nu�[yT��%�$���1Fw)7�"ftk�&�pR���̛��0������&�=�p���m�ܻ;�6�����<�d΍B��y���@݃�Ff�ƞW�3�A�l�zԧ��s�/$��*�·~���C0Ot/�xN�x����������}zb��;�a�E(°��1�A�A�n��_�Խ&������Ż��[֕�1/P���{\��&[�w�ӻ�K�7��Ϧ�n
vb�*"w!!���
']9��*�)����-۳	�1AV7&��M� ���2 -G_���n|y2t�������ݡ�뚪H��+TL߻���j�"���fvà���֝Jth�F�AT�l[8�������S���Ţ	"*����1;N���j&��6+UA:4�>>>>>>~��6�Z���U\�A��EDD�A����m̆�Tֱ6��8������*66ƪ+lh�[h���N��4�[h�h��b�c[m�D||||||�CE�QX��2��BZ�ƀ�SN��i,lI��IF��M�j�Kl�v�bl⊈uA�K:]hh�Q��ti�[(���)�Ѝ��[`�(�%R��Z��b���4h�BQ�I���ئ�5��Z�:��b�kAME�PcbجF��F���uF6���(-gm��QX�qj��0[!l:��֍S��͈֨��kD��V��ִ�٠4⢚"�@h6�ڊt��~<Ǽ�O���4��z%��~��u�s�Ay�_zF��}#o��{�i�xy���!���Pw���v��"x��y�>��K���[��k��7a[��Ѓ������'-�'���q֞�v��\N�N���\�ü�m�J�����Gtņ:$�uM-~@���&�DI��}�y��R��Pg_�>�݂:_L�da��s;�z���ӵ��iEP�/��o�ٖC��$O�HH�8%_B9����n��X�N��z!���ǫ����ш��ܽ�$h���\P||T�:%�xg8��[t�����'��,��Й�u�!j+o�X �\��N�POO?lU��f��\өe�p,A�?GX���{�[&e�j��Gp������V�*W�]�z�=sNj����$��KSP����n\�a}]qwȎ$�p<���R�~�U����[슱�B���e^�\�+�&�V��H;�m6�oBK��J�מ�x�����b�k	ּї��w�`�in�2�M��pAן�}����b�x�s����A��.��7������W����Nf)�wC��Q��x�~�7U\=�rk��lm����/>jsk��I�]�n�^EH�%�PofMf�
E���F��"ah��SF.�alx[Z�'�Jے-��ud�B�O�J��"���ߋ�=<^�z���sZ�]�^aO���϶yrMO3EPؠ;7���Y�����͸��h���ˌ���#�]T%�	�Y}������t�����Ks([D�2ŖJW>��}y��W��}�$3|�:<��v�6*r*1�2�轼�9qX����ǖ��&��P��l|���� 0�G�r�/bT���[�_��t%rH�Tk��c��ʵ>����:}:<�G�d^�9�fY�#c�/hMv�a�/C�+��|$a ���������l�=��wv�8Gov��&F* �L�͍�Ļ�ve���O��
U�;�Z6�6���]��H�NE<k{(K���`9�k�7�m�s2����s�8��͞��gUx�{�K6Uҝ�s>�g���A&���ّ�-����pWY�{f4�n�����V�UU�yFg�W5�Δgu�J
N��pr2%�95��Y�:�cϚXqҘ؈���umd�
z��=3�j^[����0�J�av�N8�a�/n�n�ԛ@�W�f\���A,���j�Z�vr�$���Ly�m��NԴ��%q�����΂��u�ah�ìgo��w�4�қ�u;-`ж���h*[�o1�;��p˙PB��F�#g7�Z�ފF�����7��כނ<�m-�f��Rh�-T��_�b��-���S��=��R�R���ǻ�PÉ�Θ�;}'0����Of����\���Dv�t�y�	��Q�o�f���w����c�s��Ƕ�̍N p��G>�nS����w�xN�����+�m+�mݖ��������&P�bxyXVð�u�+Q#[f�2��L��{f;{���G�ia>����d��n�ϐ[r7���<�v�rꭺ�>ٹ���5�^GZJh��1�0ݶ���7�[.k��7����y'�`�Th9U���l7LQ�U�`���a�֧���+��g0�D(��dU;#��+�1դ�O
��[[�y��`xD;�낢ě΍M���כt�w�ٰ�z�����饲wUS|�ý����O��Ǉp�Y��u�:��K��Fjrp�Y�Q�I5�-��X�g�KC1������P�
-���G$T���8�1����s��wK8�Mf�]�>���x�����[#��G��ʅ{�7v���p����(lZ�tl%����Q(8p0'gU��I_p��1+��M�Fg6��(�ԅ�a��t��О3xeP#]M{õ�U��#�Ṇs8������p\�2�y�$$Fi֎Yj�-��CX0�(4Y~����R&�����׃���K6@HS䬄�M��V��o��2ۦ���6�Ϊ���ntv�T+���#"�ǒ�� �PR�m!�ȷ	����'�n{����L����
<��=jѨ��9�W]��6���jO��v��9�io
��r���O�g��A>���kZ�;_DTW�7����u��.�^e�Z�9&���ԅۏ;2B����<�����3��gگzo��8}�p���$�sɟ%�`���L�p9�ǟP5-]n=�����=˫�l
6�33�dЭe�%8���xgo]�KC�$�\Ϻz%�7훎���Mc8.pä�7�QJ���zg������,�*֘�����JEӓE��A�porY���'i���v����7�5���I�s�:�$��� ���ޟ}������H��ү���<.kڿ@��圓��$���AL��E�9s�ؕP�����*+��ub�NFu�5n���9�,&�0�/!}�a��O�3���#�9��\���M%WM׹'�ٻ�:h�9�o_���\����}�<6׫��N�����K�@7Pk[���ކw��|}����a[�k�A���"�[A[
6����7�a[V:�&�t�x�\����ᣣ�!�E��F�aUI�>��]]��7t��;�N%����a�W̋vl���"�8q�w=�o|ΧQ���"r�Ԩd�o_�p��e���D����{\T]^�Uأi�z�������i3�GDj���W]~��H|��w����}�%E�6���&����XU�a�.#\2M	�26��x��P�dD9�r:���q]��wy���x�g��o�ĵ�VL�K����u(�������o*����=z�9�z�$�q+��p�b�E�7�b�c|��L���/2矷�rp�fz���j�ׄh���)c��g/ze��;��'!�'S5�%X��˵XM�XӾڹ��gB�#^~��+J��a��D[?T�Ӗv����#.��J�\��.��ۺ�sul���VIt��7QM۵�֑ϐ-��(�;�s���q�R�EU˹#ב�7l3��:�+F��.�56˺�RkC����B6��������V,Ě\���Ӧ�0�'k-mW����痲X8"�9Gk���m
A��)u�H�s}�[3ՓiH��yγs^r��SW�֫�B�$p�",1�x��ھ������F�91�$$gqwaz���9�|<�H\���˝m�_G�-��62 �پ�>Et��.�hWn�O���!3W�5�o�H�&֎�l�Y�}���ê۟n���|��,n�+�sA�	�ݏ�h'/9���po��x��Bl�ō\��9�W	ް�l"�g�|��~��1�z�@m���	;�v|ʧ�/\�������� p�sn�o<J�N������Y1F���ʓ�@���(b^90�S��G��hH��2����.��S{�a7�/�yx]��}�44�����]�)�e޳k�cڷ_+:m�w���	�>|5�c7 ��F�Qo3%
�f��G�K5>޳c��Й�6#���p�F>���Sޅ,��3�F3�wP�>��ݟ�X	��f���bAS;�a��\&�ݯ��M�c��A���U�S�v!����9%^3{�Q��ɮ�wv������X~��N�>'�V! g"�yK�]^Ky�&B�T��D��歈7W��eUޣ��E��Z�E�4�ґl)�l��G����Q�m��Ê�jN���t/Y=�e�,�PT����@�d�搄�=���t���J��j�-�x;�w�M����t
�2�x�*�.���ʐ��[$���Jߦ���r*D"�ۍc�j��G��]ݦ*�W�ү�Wc4y6n/l;�зP�ʩ���R4�����
v۔�"�+*�T`�/;��]��-���M���3� ���&�C��櫃;*��HEk�F�R��S�L,_F?h�l#�v����z�]�=�ޠ��M	�ۛ��-����=Y��m'�ݺ�g������q&=�JA��^�Ggܷ�����6�Bz���ڼF�|�݃�2��BjL��=gp�Su-�kg�������K�<K����O� �HY+��Ո-���ڒw���\�|���+�T���ȮZ������Jq�`�m| l5����lƤ�����ܯ�v��+y%Y�$Ҁ��lm@-s��v�]����X�݌�̓T�	��7*
��c�h��]�Aj�����s��O-�
Gaԟ7��:J�HͶy_v�vt���u�u�@��*Hj$����3�Ǻ�s8���W=�HS��j�c�T+;(�p�C�0�	�&4n�)���tQ�c��1����%�ww}�Y9WLm����	���}�(.����v��ȱ.\��ǖ��u�����d�����0�xAH�V�����u[�WO����y}6xvj���,�p��({��f�v�+��� �PSS�	��Pc]���9�6�Y7� ���4*�S���9��s��忊+��
�qD���"�}����^�W�����$NGwS��=�q��\'����n��w�������͇51��&�����^�\RY&�j�UZ�[���M'P��G�*%�@���Y�M�F�^4�V2*_en����J;U�sM*R����;ǁ4�=
���;�pn�։�'r�={�N+z.���(J�J\��N6��r�d�HYa��� A��b&���s�5Qn6�k�w�$���t$c[+dFd��L���T��e�1t"H��郝��DOҕx��7���/�vx�+^�-G�]{�>�yi���B�@���>9s�bUes�7IQ]�!�$����G��\��̲�#��z�a�N@NòN��ڢ��6d�eV��Tkb
�Ƀ�� Y�w瑅6�y�+�	F����5�{��4$/f��#sTf�>^�i�p�Y��{o·��o!����4<T�������N�y��ם�59|NIjD��NQ��6w��ϻDupc�y)����Pb��&�̍/]k�w�SC��[�Ȫ��X6aVŀ�+\�F��Y,U�I;Oh'��8�����?~��dp�4�3�Ȯ��k^|��=�?t�ΣKP�Bxuk��v!�k.�Am�)�O^:�j0����m�Mõ��A�Z�kF�w)hE�&�jO��z�^��\o��8A����@t۝�39B��:Z'@��m�p�4��J�M�=î��$HI!!�y���z/�󸷉��[���nr���:!0�������f:�L�6�X̚��M�9f���۬�U07_u�I� �=�\Sa��{0��1|{[6�����U+)u5]*�����B�%"�O�Lt�b�F��A;W./s�LĒ��IP��P��>;w"��Ϫ���"8m=5X��<��k{oia-�^#݇���-.��):*t?̮��~�U��9Y���Kw-��ja.�#�N������'��'��Ļ$��G�kTk�<��O����B�= �(6�6�m���&�lls�u_�7ju]���Z�G�P����0Ǎ�^mmr}(|�¨�ɯ������Y�rˣ?msV�H�{�/�S;�_P_O=��͹��}S��w�g��N�;J�S=��C��;����u�~�c�[���jgX�4౉��1C.Q&�X��ڼ7E>*��u��+l��7���-��v$�"��1�7�C.��۸�r��9y�`L�ۻ����Y9*��n�����\m������i\(Ә'
'm0�6�f���3���y�&)�C�> '�q��{��G�+���֯][�opUX8}��]�P-�[c�b^��tz�MA�7r�6V��ͪ�ӠX*��'��]��z�m�{w�WC��켝M�)3uUP�"���&��kfJ��f���\7�8w���@�ia�����X��@� \��)� dO{���pK|?t����*`:4P�g��X16�c�*dw�����Tȋ͉��T��%I{�SbҊ���KF1��'��K�z�_,��Oh��8cc�.��'���r����B��#�x�T�뭖�C��=a��EP�K�owZ��s�	�N�^\�8���8�d�DHJ'z�MXݍ#��~a�Uv�=��7�I��u��N��8ߚ�"���#�� c�n�g
;��xn��������j�^��˅�b�p������{_�Mp�/�|F�����!�k�KV�E[F.����z�[������%�Z���r6d}�<6/ykg�J�<�`j⡏��N�#>���;����^��.<0���)�GX���r�ҩ͞����0�6�s�ؼ�����3J����t?��C���y���<��L�>���*gY����۾aC=��[��TW��*�Ng�[�?	Ēs�yr�D�N�5��׋G��}�%	4��������}W�5�nn(�]��d��N?0O!L[;���
R��Wr�r�_n����Z��j]utU;}����W[���I�<��bw���v��}LE¼��Y�b	Z��xq�����!�G���.�o�o�`�{��h9{��Q�{}���Foq�#oWƧ�QO^}��&I:{ww�������%�d�j�b'qa��nRx�\<q�2ĸ(�5YQfM�<�/���ؚ)��݋w|�r�[��ң��-
����������֑-�{���1:�syhktd�v�>��k��,��w����$;�_�V�����m�?'��)Zs��^��o��_y��-�V�K�r'��YW���Td\7�,ж�LXU�ݦ��93W�z���ɬ,��	��<1�l�W��xM�ʼ�`�x�����鑟i����E��q^�'�;����r���oa#Nm�K�	6�k'rj����^>�	Z =�*�ww�w���Kt���뜷N��稽Z�)���>�:B3�Dޜ��}�gxI�u��;�%�ꔾ���ѩY}G#ބ!˝�P^L�uD���o���"��l[p����C��!���@�C/H��,I	LA%&5��y
3��K��h�V�IA��h4�ն-��bk+1�?'�?g���mgN��i�T������U�j�A3��`��F�m���i㏏����ꪍkh��ţF �*��j�`���lF-gN>˥�:��J2�������h)�0U5N�щ�U�thJ��Y�j�(���F��kM���V���������h�j��N�%����j"lZMQI�(hq�(���ZDE&ֶCA����V"�ŭ(��kl:
&���ѧk(iLF�]m���ƵF��h��F��F�&��Tj��AEQMأK�ӭQ���:uE�F6ɌAT�:"i&h���c�(�
�lm��F"�lAl�)ڱ�$�!EX�1��E�1rF0����1�Q4E�
����b�%Z5S�R�(��h�~$����h�vY��kv��L�r�6a��!2*t_ΪI�.��*�1Hʫ��a��L���Ȫh�̽
/[ȝt����z�@�"��i#)���@j?;*ʴ���?J2�㭰_@`��m�(�3�N��ɛ'{9꺖�RڮK��z�|�o�5����	�w%��MF�_���JZ���v�|���i�ױr\�3<?�ȼ���|�#T��G��y��WH�b����֬#h�{>���Bɉ�c�Ǩ>+���m��(�Y����q�|�^}�#$,���=��==�;D5�Р9˦3="��o��mk�y!��Q��;�|N�>�$;��Ɏ똼sR��-#Z9pU�ni��CE?H�B���]�a�D�C�j�D7I5Y�y�ݚDwXy��R�7܋@��;�s��,tB���*����hf}~��3zƑ6Az�����Y}��M%�i͵"�l��V������{�O�(��d�ތ�;[�-�y4��I��p�����/&��^荸λ�ݽ�&�ٻ6���̄����{�g�}��i'�{g���U��V���N��]�����9��nr
3�����-&�Y1��s
�1J�Tf5HB;��y��up�\1VýB�#)��2��4�{�i���3U��e�ÕbؚÕu׼;�������!\�<#ڵHkg]�q����oDx��q���7v�'FHgy����6(zǘ���j0��#�fu�®�o6v�;~���%U�ہ�N�V�A�c�W�ܡO=ƗV�/�i��ț�r��a��C^x�]�=�A}מ��-v�qk�ٓH��\�V�n�潷��%	���}����f��?�u��Q��:v<��'��S�'�*;b��!tQ�JJ�����`ɧ�w��WV���ш��d��X[.��ٝT:M0r�y%{�{��l(��3Kf3_���k��Zv�	nɡ(e0q~b3���⍎���i+�����.��^�}k1����
\���'!���a�o@~�kd-�;��CM=V��ce�p�]PK�|w_�{�>������%�c�rws�B"]����zp�y'ؒ򄗱�cW�ft^���=�X=�[�	|3�[��3qһ�QF�J�;�J�r
)�E�;:�a����e�2����81�땽�R3�C�;��/v�.�[���¼�sqQ���x���pT��I:��g����G��Gls�-�����(��c=�@���;�4����WV:��Kk�_f%�d<�%"#N���=9\9�U��`�]��H1Mwʇ�j��98R��!0JА��2n���.�Y��_��n���Ϭ;��=T�	�<��~\�P� ������{Sv�m�'.FD#����X��u>��+����h�.o`�%�7����ս<2-���w��fMA�U㹒:i暀@�\�	���RS��`�Ps�>�[��8���<�E%�I��ݩ��}ْeMT�{Y���6�8U9x�p�u��̈́M���I��"�z9��}�S//�R�3��B��c�gb�@�и.er�����6Rh�kx���vq۫�}��݄�����Ҍ���W�
�cs��%GU����~I�y�uk�ѝ򮶷����*:\kC�.�n���{�f���ݽ'�@�^�;ې�0`�����Zz�ǂ<�Z���1~:���ۃ,-}�r�e}��2�<xI�v�W��11��t�h^��1e�P�忲�^4��m����>���Hf} )�ƥy<
�՜x�f^a{m�����۩Ȝ�����qp��%n�W\:��>� ��CvvGjb)Bh92������#����>�o=�����wWЃ��h�����yo�RR�,:��~~��ϣ��ε�L��6�sP�|�^�7sV����J�<+T2A�of�;�q�$�nx��.+7k�N�r�iݝ��-���GxmĆ� �m��n�Cf�+�p��e����$����|�قf�e��y�q�3xsM�O���� �@B����5u��h��"��L{
�u�O���U���O��4�ڞ�`� P�����s�TLN����۵���+�jҳ)u����dө,�EPF^�c��C�3�;��o�8�fJr.D��l+�IiJ�!u�n�%��d�0�`��*�M�I\�����}۱'.c*,fY�w�7��L�s}�g`����8ϙ�|�t;���sr�2��u�w9��T�kj��YrX��N�����Hzh��)�o{�ĎC�|�׽��:}��e���4���G�O?s��U�G��%<ܚiD���uq�ޒ�5saV�Mz��{��]̂@i�k�J���˷i~�''o�U������j&��\F*���F�Ғ�^�b�5�w)�qû9���S6���I�>Q!��<|�,�֓I�6IW)�BI�R�w'TNwE�wM�Zh�hG���	83fמ ѾUS��4��3x".�kM��ۖZ�z���D�Oڌ�����-���Ͼz�":�u4Y���[���{�r�h2��^�8��6�|i��3���TYl�g{���Z���ML ��=]/)��ւ�q�ԑ5*l̋�O����L����b�����"?1�R���/;��g�7�8Sn��ǛYq6�E�δ{t���= 3�`"�6�&p�g#��g���aXg��9�v^�j��*��{��OZ����^��ΰ�D�1��Y�+7�J�kpn���t͇i�d�Ga�;|8玏Ȭ��l~�Zz �'�\)|M�o`Ր�`T��*�\r�5��f�����}���xb�TPGj�{���1��Lŋ� ����.���.h�̀K5��%tL���g�]:��Yڏ�����Ҟ��±'ٮ�;s�zobtY�B �=��$�ا��d��,��/	��㙳ne,�5uW{Q�t������K�[ ��>ا9"^�ts�����Ou���zC�w�\z�3�iI�u�tim�6��26��u�ļ'p�i�ذ�1Ç��e3����F��!e��J8����7��A]��}��ٮ�ꘗ�pڠ��pѫT���5�*����sK�����)۫~���۶`�ϻ.�U���� �"�Њ�b3�s�1�23�(�$���  ��4{;���J�Ϸ�ju#K���dpX��@��rb޲:���޽���^��<{T��.'�����=�|ُE���O�)b���r�í\#�<���/��(r]r)�s�v�	�,T��z��(��*q<o��f�	$Ib
��]]7=^�3\���i)+���v�ݣC4&9
�>{��u\�O S�xvצ]Q�v���Eб3�#WKlfF1���Å-�V�'�o�K���eޤu�ܧO�GQ�]��潀��/8��a��w���ڷ�h�A�op�{{��^���TQ�����X����v����y[�2�[xj���+f��.���W��9@a�0�2�;3�P�sF��^��fi�Ws���v[�Wtr�_p�g�Ճl�3���l��#~��fᕠ�]ű��3���=��eE�_���a�����]c����J��~k*��\v�t�c0��D���ʠ	'�c��!���D�I���y	E��S�m� F���KϽ��C��r�l>����u���E�A�$B>�v�J8���T�hV��l<q���7���C���"R" \�������o ]*�·=��s��`nx=�4&j꽘rF$�8�������{�&���><��I����a�=�A*��OP����+�筣d
{��n��=r7����c�1�s�z'�ۢM;�h��ݩl�b�a���Ǝ�EoQ.F]乳&� �s:%�][:�("�;qj`��n)cLTd7C�$�>x�5grFh�M�B��0��oK�+�^s�ka~=�tw|8�WV$f�{ö�D��垛F�����s}v�yۇAn-���+��cr\��İi)��!��G��=��ֵ8r���O����ӱ�uE�.�p�f�wwJpY�)�5#�}�ȣ�c	�$��[��;1������ �Wի��iz!OJ v2g5��dI֎'yy��EN5fk=Y���3���#"!�ϼ<g��y���;�8�+�*��\o����6��v1Է����j���jՈ@�rǸ�n����WbUB��Qz�<a;�9ݺcs���O��2t�������l�Xڷ�fJ���̚�����/܋�i��k��o�ܢ���W[=Lی�l��X0+�����P��dL�+Ħ��,�����g�*�:���GҺB��M�x0���1�Ʉ.�w��Z�����_t�J�ԍ2���[ϝ��d�c�U�Z eɕ
�gG�dJ���7���5�[���}|;�a}F-}�䂜��J����'�TOK`�O��^���rN���!_}���:=C ��r2�E�<LY���r�hj�"����ݸ�I�Bh�|+:Ɗ��_�¢%.E>��T$m\��3�_jP�~b�Vx'}���JU>������ۤZ78���W����`\�����a���"H,�O��L�=�i�3���na_Zn����/�8X��D�ח��@B�=%�7l�MzϷ1�9Y;s42�4�z�N��qΒl��ɯigE<l3��r	X{�5D�ڠ��o�h윪����0�[`�
�	u���R.i���
��L^(STg����S'��q����*%y�dЃ�!m��ӓ���S�0v�i|�7J�E$
��Ώ����g�>����ϊT!F|����lV-����T��g�p���З[�o��zRV�L⦧Ӑ'�c���]m���w|7앮Z�̍�8"����e�6�_"9߮�N�^fo*�K���{{� ��i5��b��5��^VN��z��#"i����$�$��sCRݟ ��������P��/�>�1jq�M�N�g�����ʦ�^���?'�6;O��K��� O���ʛ�a����u�H����[
4Ȩ�̷3v�u����(ّ������)�N�� -�و���锣j	��ڝ���%`��'��ޗ�������w��|.��YsR��E�.̪Gh��:���Un$���)�܋�|�*cS�xu<��/��������n>A������:z!gGY���RD�ҧ ݍܜ۰DV�t;�Y�d�ݦ[g�=�oh��	0���ܝΫ
�f��o;��q���W�	��1�Z��K+��~��g϶g&,����v#�Q��ű|�{��UZ,����Lt����k��;�#a�Y�l�]K�rL�4���#6p��%<���A�{���(϶)��������Ǚ�ҍɜ�;�^g47p�9tڮ;�t���=�jRh��ח9-�3���im<{E���Uݗ�T�^�qDO�� \�[�4�ߔ�ι�}�]��h�Ͷ���
��滅
�����!ex��HI���v�L�[ۦ1��R�̛�`�4�QB:�豫T�����O7��=m̋Y�a_,��ɞ�0zd���R*���NEO��������S.	�_�{���
�6�ݝ������Z���{�r�Ft�fK ��;�y��]��?6�x��;f�9NH���^ֺ�Vm�u�p�Xhf���w��ro�o��Q���|D�n�j�ea�8o�n�v���{�^���<C&�H�Z��q�S����>���7�v�e���V�_���w�Îi�87e(��V�9�T�V
@�a�|7=����@'���zV�^�Hv��~�7n{�i�
�tL��Y}�o��^���]w^�L���٤S�@C�[w��0��a���@mS��(�;���6����;��M{��CQ�nZ ^��p N��j�ýo�`�PԱ�V� jgq�oCvx��k7�o��ތ3�\g��|���7d�f���`�C���W������~:���:U���7�K�����a�d�ףJ^�d#&�3Ώ>h,�6�#���ټ�K�5��+&��sT^�n�ˑ�z���u��6��G$�������]����e����<�G@*E��Zg���W�!�sU^a�x<:���٭N�:�`��Ga]�ơ��_'�
2�OĂ��!�ų7���V�(��Zfb4���J�Up�L"��g�kzo�k=l�N����~C�-�+��z�{<����2�M��{�p=��ш�l�ؗ���'`5^��]�ѯ(��Т�:��g.���@��5�}������_`t{�{"̇��k�>�}���28��g�
��!���=0Ptc�5�����j�������S"���6�����E��K��'�[��f���B�ܰ`9�9��0��o4��ǾW���A�� ����F�mL�{�n����j�m#�޸�"]��|N����l����q^Ӣ�������Z�՝�y��,h���>��}{f���������?�Aw�?!̍���M�7�Sd��Є�.��7rk+�K[u-�cp��S�P�NA��"m�K�t���rzUE���s}���=�N�[�zv��>[���hY&j+(�m��ru�`GFr;.�ݞ=׵�R��o�*o�n����Q��F���<X�).D��X>�~��F��{����V�b6.阢6tɱ�+2f�e\T�yF��;����ԥ3�g/ ;�ۣɬ��j:�}�#CN���ě���`���;�Z���^'��Y;�3�}�rf����f��-j��M�;�-�z�\�ى����;�S��`�i#y(�Va�,�1��+�cv�-�O*H�>--*���<P���t��0��s����.����2��,��3qN��o���{��pp���,9���	��9�\*�4�Fz�t�G�Wf�0�+;�3����^�`P��ŴF�5�)�#w3n��)<Y���%���Vw�F�l�p��]�@����g��K�j�?������O�_+=�,����"�30������vƊ�*gQSM:��-�QA[�֊c�x�����7�QTUlcM��*
��j ��ڃ[:I�$��]�PQI�.Ռc�������mm�k�L[j��&�gTTV�����h��X���.�a��TQ�c�������1�M3A6�D꒢hH���m��mRkF�c:��������ࠈ�*h�cV�h�ѣMh3*���U��(i'V��TQi4F�6t�}�mh�E��b66���mf���k��5-��Ӷ(�,F��T���4f(����,UDQLZ1S[jk�E��i(�b	���m%[f�mS1�TScbŢ���6փQT�6΃F��v5kQ5N�6�F��E5���l��Ӎ��֊"(�b�T�k��N��0=�}B��^�Rbdd��h7�0fM�,��Z���T�ǳRu2��t�w�b�8q�
-�w�f��|�8�@�Iaƛĳ1<�����	���4�UO��.�i@"� �S=��:z�t���>����OzRW�ݡ1�y����t6c��t���;�YŹ^��Ad��#���Q"�,�&�+	�<��'�TŬ{�5�`5�^�{-5P�@2�S�z��<���gԆ?)����y�=&�щ���^I)�M���vI�Vù�ٝU�h�0r�y#�=Ŭ�{_TMnj�{�_Ϳ�/�0�`���� ����׶tR16X�A~�b)���v�Ԉ㸂$v"{�Ǩl������E�c�'�<U�}�bjn�>�a�sA$FBD��_��h�P��Q!G�l>��g��NV`\��G#���C��='�Ï��2GP�TNZ��pT���W���-m��8,gF��V���e��H�$D{N�3�����Y��8&]�WB4⸶�O]֝	��ۣc�A��,���@�k�vŃ��ߦ���'8��"�L�ϩԍ���R�μΎW'tn��;�b�R��Nv��^�.Й��j�*۠ڵOsTB���L�٥m��F*�N�R���b�PW������S�-�;�����: !^0�𙫪�98����4͘�Z'6�շޤ�9f��}��}��OK8�^�V&.�0��͂VR'��׎���1�OTD�O;Zc��R�c���Fp�� �w�o��I4�����_cN�]�a��X���u�,��:���OM<M3�Ú��o��XL�^bu�{|���|#o�Y$y�%^)&$�=ڟn[�i��Qb�I�M�'o���Đ�b�� �؃�c6�_��%}7���#Ӕ�-�[:Z��nkT��<�^���C�����ao�'��)i��Ӓ�u��};��t�I���'������1�K�VH~��9s�bU6���w�sS�U����q�Ot���v��5��cj���%�7�qF�n��ZI����$��<
	�Wr�[����`�q��7���[h����Hh��N,��|#������ȷuZ6�5�E����>)Z�f��xG���>�u��৐���U�:l=��"QI������>�=����d{-�r�S�&�\bU�NB.A�%�QA�F�p�,������=s_�a �0af��{�����~��A���&��I:��ӫk��R�+��6GStl�l?Z���h�Y6v_p&HNÄ`�� e�T�h2��=���h�gJ$�3�17w�k6�g�@ ؚ�������-�����ۙ�V�e�p�{[IS�tYw�"-X>�v�<:�7���M��ka�;��3]���܄��n�/y#Z;���IxppT�K��tB[E������vfo���0�/v����[�"l=�&�V!Ȗ��â��8;��r	��5)��=�A�����{>ۊ��[gPSJ̄��o-H��3��LD\�*e�����op�F� ����F������B��*��*�u�A۾}g`շ�����UA�5��Z�+��'!�u�غ@�AO��48�fd���������^9vO;H�F^�~��k#��&����Д���ޔ�wm������7�`���{��R�x�ш�����<|�����t�[}���Nc~��ً���"�G��{x��s5�OT_�Ę�yrҫ̋��f�U���v��*�2'���Ǿ��� �_wh���O��y&9���Ckڢ�o�L�7�&��̖�Z{��/�߳�Z�F��d�tV��q�"[;Oe%����+;����ҤU�ɟ,��},[}RA�pX9dvˋN"8��Wi�U�n
�/V���:����?b2�H.}�8%��	Sv��ȡ�@y6#��muv���]^�M��Ly���,������ ��`Ty�ӱ�N�2����Z�&����ĎnP驸Z�^�3�9g4_���8#�!�Z;s�R�ah�7Ӧf매+;n�q�X�S�T��|=Ԭs�N�*	�_OGҷ���E��:�FJǫ�j�;2^S��y�8��y�J��vY��}Cq��vvJ�=_]�2����{�H0{�;ا��g�1�6"-���U��+�^��=o|:�ҿv���3x�	b9�*�Hا;�ܵ���9/+-�j8u팱��x�)U��M=��O���p�z���P�(��Ҩib�7Su���1&/�Ww�i{����Y�]�w�jhg�jS�aj՝��g{�oϟ�����h(��'?<1���n�9wp�ܲ��8Ҙa��3e���_#[>Ґ���H���N.l1��*��,�sYm�<3#�+����;����ة�,��u�:N<���۹~��ݵGI�G�.'άW��p���uϠ���T����S����=��"�.�F�N�)Juр��N���@)����|-*���{9]\�U����%��)|k��M*�����Zl@"�D8����8|�>0�ȹ!pc͞�BDi�C\�4 ��=�Cf:h�c����".����JX-�����W~׬=O V������}���>�g�藼n��i�嫴��zԯ{*��<�x0��߻����L�-y�I@�O��rZ��En�_o�q-�{��>`J�$�	�q�ڮuWJ
��Bک���y���|1�o�س��\y>���f����
���;�a�1ĳ-G�[�miœ%H�wS9q���t�PsPz,���c��a��F�LV�ÌGs�,�t:5�d_c�u3	�;\���v��cz>�}wI�".41d��Y���b�7e�<%���r�M��$m-P,ɺH䬭dN��not�h�E�¶����`�:�*�ɫz��F�L�mx��#Cs��X��C��H���]�=l��pg�ܓ���Һ}(d��ضA�z��H7���{d7� �0����7c�˻y�$D�1�Ogeo���:��L!L>��5�h޲�[jc�#o����f]C�QZ�𔍊�ot�Y���jI��leo�3��~j]��/-� �e�B�Qj�t	���Ó� b�w�d�έ���O�o�CK�9?��0�Z�Ϭ;��^�P�z�͞i�̓wE�L,}�7������ρ�	�-�'�=Q.p���,Ab^�!EX|�����A�%��
;���1
��utruU̡C����͠�j.sr�m�ٍ��6D��#mn�r�����g�ƕܘL4��=ir˞�yz&�H9�#d�>�nIɁ���I+瓞v��sS;U�Ld��7��=�uo K�5j�6���Yn�r]�o�v "md�89Å��=��T�6�<z`w��/_([��}}��ފ@��j�Ŵ+ϓW�8�r�0�|��uiUoq���u"��h;E^QOPyn�\�rp���^]A�k\��:�?4� YL�b9�������;��kd5S�����ӲGH�2�pQ���|��SUt/�Emݫ�iݖ�sy�r|9[�@�~�ǝ��_�vچ�&��d��}&�Oc�wb��gE ��]����X�@fо��+ɩǉ:���:��ٕ�]}\GN��4�Uk�E	[��x��%�>�}3虜Ť\egSS�����ʡ�0�ge�2���Ӫ��J�+�ˤl��C�K8(�?N�Q��Bg���6���/��:�������)�P����%3i��x�����2/�+�d��f�\w��-q>�DJ�K�zv�{D�=�'�ڭԎ�p�h�
���lw/H�l�y�Sq��f����3�t�	␐�x��Q�/�/G:��.����t6z�d<gDEOb&���j9.Yg�a��dH�ɮ���x�;�i��:4�E��x�{q���Ln�d�s�nM6�D�k����[sx�Ɂ2�C>��e�\��9�3�tu�E˻���毗:K�������ɾ*���c5��龥a�G��'F���J�^�l���,m�ݸ��)��`�U���.�hhl�,��8:�N�>e<���uJ���o-^�OH��x=ǰ��ҽ�
38i	`���%Q�8�t7�V�.����fZ[�$��ֲ���v-�|2���``̰�� 율DG�^=����K����7�Sk���n�J������s�wo�馯@�FO���"6���l-Q4�iM�}[�Ax�@a��O�u�l��Q#�T�����wqՆbN;'|�N���4���x��*��&Vv�m�-�S��������Y+ȓ��/�6����]QZ�;��J���#/�`}��D*���fn�E�:
2!*���s���W]^��vA��2�Ӯ���7:Yw�&�	���,��H��^�v�tu��ux$MK��zn�晉�~�5�û����EM�s��8�@��ѝ��������&��q�����R��9h�k�O�.�~'tX�����o�v�%�s��񑗿E�x���gp�ZH�!߃���B��,̟�
��u�b�v�/mz��S�6h
l�M9ޝʉ��}���"�ŷX����̉{u:�ܼw
ʴDȼs��͆��e\z�|;��؅I����#w��� pWW���Í��Q�g��y����̾"B�:	8�` � uk�t�����D'�ʉ��=��&��V������D�ă��݂��V
xj2�dQ��V�{靤w�,Ԯ=]7�lv���sx�	bRj�т��,F�Uj����|�-F}��G5�CU#Bg��r.u$$�	4��M.8cd.���|����f�;��Е�dN�mh&��ĘX�FFϷ�X��;,�*�����#x.�i��s&��z��)�������W�铏�=K3���U ��@�*�t�˹�n�U��.���s5����k1Y�����\�&���\�@7A$X.������˭4"�1A�Z�VE�Zӏ�Hat�
U�Z�����ޤ����E#����P5�|��lm�5�cD����7�:�E�Y�k����t>V^>���|����'++��Je,��e�-!�B��1W�0��H�)�J�	��rN�|j�m�Oj��!��9�a�#��s��E�Z��q��M�bN풖�m�N��r��6xt��2:��jJ(�~��F�v,Xړw�m>=MS99�����8FxRϧ�x���t.��3�~R� )چ�E����7����m�dDDD�2��]!v<x�@h�k�/`0]�Wk�ﳬ�s��W�o�6�a��e��{�L�U����x��#z���t��z�u�N��aK�3�\<�������價����s����A��[�@�u�����ʡ�@uH�`p�7��G�1���~�v�Hb��Z�9�8HW�܏ ��Cq��{��tw҅��MЧ}9��>�~4�ݗ�*a5a>�L��Ǫ����Y��K���67����2i�C0cQ�3qq�G��AK@���E��n`<&B-v�D��/x�h��M����t�:4u6D��p&���x ����w���?��N���0 Ec�(
��x�EQo���x�e'�\.!H�H��V@��P !T BE@��P %Q "C ��Pª�B��{  `! ���  !U`%Ua��  �� "��U_m}b!Ub ��  �$ 	
	"�UX��� � �H�T �!� =���D($�b �� D� � "��"T
`�  ��Pe3"�B	� �UV�  �� !� �� 
	@
	UX��P �� 7p=� @@  � @@ "@B����. @������E�
 ��
�	&O��2�t�z�35]���;"����1k��ͨ��4�uq��垜��Kb��+Q���|�v���h�*+��A�'�����*������f扂CcOy�*u<@�e�C�P�HE�!d��4��� 	��*�*�B��*�0 J��"����� 0 2*����ʪ�ʪ�ª�� �*��  @2����  @ �
�$ , 	  C*�*�*� B��  D*��  2��� R��  P�	@���I��?��/����(
�@
P� ����bc�_��e&�Y�Фv$k5؀
���r8PMB��J�ΖE&@��� 
�����;�4�BK��HHIx�a�Z��Q[��P�
��2o�����c?�����o�?���|��| 
��H�//_+� Egi�@��k�s콾�}��^�rL;ץd, 	!%ڢ[ Q^q�#:��A���^2��k��|�A�
y��L7�  �Tm��8���5�>vmR��X� Ep�fmi� �u�l�Cٝ��?�(+$�k!���?Wk0
 ��d��H�{���*UHJ$�
��EJ��)E�E�R�"�UIDB*)BUQR�T��QPR�JHWm�mV�URJ�*�**�HJ�����m����RQM�D�@�"�� �T�b�QU(��U@�$�{�֢�
ZР*TSL���	��@��R�AR�TT�قP����#bڍ�����J��@�
�ة*��*,�՞�HJ��   {k�j�WhnꝦ�v�Fu�m�;��Z�E�.\4uJ�R��٫�ֆ�Ӻ�[knڮ۹U�E[rӷ!��U��%+�Znv�\�ꮃ:��u[3�R�)H����
"�   s�(dhhhdD�{�n*{5�ldH�ԉy�B������ӏN�H��{�{kz9��u5T����rZc���&r۷k��Wk�;JV�k��[Wu���8-ӧMm�q
�RREi�Ѫ��"��   {�P��ۮ�A.�mV�U����r�wn�7Q�[.�wpn��j*�����wJp-j�ӭ���]%J��1kmջ1[�E�WwwN�]�u��v�@64�P ��   !�z��M�)ۺUU]����ꫛm���v��ݩN��ôV���W[;��m�:��*h��]s��n�8�[
�N�5��M�UEUfP��T��   {*/j(��Y@4��T��Hr諻�R����� �3M�QwZ�P�����MGU����D�TTT�S����+�  Gt5�@�{�P��pP��mmӺL:M�mV�4e݆8��N����ҩE'q�i�Fh4�:��
Qֈ��T��  ���=�Eݰ��&�:���h4���95:(j��5U��t:]�� �wH t�	v�րuӥ�l��A ]e�JH��  ��@��6�i���K����˸ t �-� �q����`  wt�� tܧn  �0t���u�T픩*h*��G�  ��t��� ��n�r �-F t ;��    1ɀ: �a�Р�K�Ӏ@Tɇ@h�)
�B�5J�R)E+�  �x2 ،  �,t  �%����`  ;���t ��� �*� �� j��@�"��1JU#@24Ѧ�S�0���L@����`� �JJT�  �	�R�  4	2��U2  3Q��q���	�DEKX�-7(���8��2̐�s�(�^!��@�� DE{|��}����1���lm���ݍ�cm�퍰cm��6��������o���?���G�S��/�U.��_��۲#E/	0J�Q�t�M��M�*ZUj����J��X�ʰ��#���[v��g 1�����gJa�K�p���D6�ZL5P�G!��Jա���q6DIde�7X3%�Ic�6�j�ۣSE�d�!e�ÁJ
���wi����QLf�W��:���J�BP��q�T5a֒&�#�Δ�{�u87�nە��cB�G�G��1���B�\��{��Ux� E�Z]�����AU�]�K�W	Z�t!�1�'Ljb�a��j�D�1hͰ�/F9	s_��f��C�mK���"N�mӁ"&p���Jλ���"�_ch�B�/~���$�^*7�4|^��7WM[yw��Țz�>q*�����gn�8�^�{�5t��?Zt��Q�ń��ӮD�d���`�Z�w�b�<Kj����)M���{���
��2kj*S������sMYu�-��=:�ڈ�bW��3�ۇ/w7�d����"[�`0ŀmı��#s0P��d9���[1G��U&ӕ��[���[� ��p5�n�䚊`�Z�
�c�/7-97l]�e��n��a��N���,R�̭iÖ�Ӹ��� ��]��)�7r��fS-���b&3[1�Q[dZ�vi�!,��W�m�t�b���q�y\e��kK�}y� ���fn��pU�+p�&k�.#%���a�զ�ۘ�V��yW&�˥�d�f2X�C� �t
�e�Y���ދ7���X��@<
Z.�qڈP��n�6��+ԩ�{�vë �N i�r�ۺ�l�&[�1�uv�+X�E��7*��֫%�:�0z��p%�[B��SFV�@]EF��ۚ5$m^��`)�Yj���ѧhd�*A �n�H)cf��Thcx�;�wrj"-�qԤ,!T���TgCZNfd�V�:�ʊ=�^&k''�ʱ�c���6�b��� ���� �D�wpP�Hq^��U�zUV�t�+%���mn]�Dևn*mF����[XF`�����c"��OYJFu���#P���'%����R� �9u�eS�z��B��w&$�FK2^���(Kכ(K�R��f�땂�X����r��^|�,4��VX7q���Q�r�۽��c��4�%k�,�Y
�sv:pm��+sD<��@������d����Y[Bm�q2�Mb[��5�1m����V�h�+(TkN�~	vYw"�Z��LH�M��������(�٭Iy�^e�Ŕ+F�Yie���i]�m�`LvlG�ve�֚�1��`:�A�R;wWR ���%b�E�YBD�Y�$`�+Ϛf�e٭���]ܧ`m�Iw���g%����V�a;�^Cv�v�����d�Ti�z~���ҥ��m������])V�t6��w�(�tZ��N]�'k<y�^�f�-�ȞS��lV�I���n���M��j(
��5.eB���Akkj�V%"��Z��.���@_E �b�/8�4�"���G0<�ϲ����	�f,�ۼ�2C��V�b8]��;MP�T�ou]1�@���d��'�-��k3/'���H{k����gi�b[�O�ڕ+e�CNc�:�NËj#���Q٦�whޥ2у����ChU���
��T�ګ�B�Xu�<O%U�%ݭ,Pk1�W ZfZ�2�i�J�����az�V�I�h����b�v00+KB<7X�r��Ǌl&�e����#R���ۻYXiޭckr�Q�	`��;M�n�
LRܤ��[��W��mYN,ydi�Ua1�JD��ݻi�wcu;R�g��2��E�gN�ݘ�l)��k�U�)̑�v�W��5���B�j�Š���v�=��4մ�v�˚`F�Zd�4�"�Z���PT:{�:�3M��xY�*���5m_ї&5��3��#_iǥr���
�c@�q^;!g���5i�Ov* ��#�Ywe]��H��f뭓."g
zY�J�e��w���R���x�x�l?�#�2^�w��E�I�@*��l�#�4mid��6ݴh3�KU�F�u�F��ܘ� �&�e5�� �Q������*��@�;.m�&E�B,��;%�SS�0<&[4���V9H)�o]�m��0�	^K@mn��J/4�GZ�Ś�&��1k���@�q:�A5U���Ӧ̂��������fh�7wV���M�i�2���<�l�1�bÌ�3RevGd��ˆ�-TnΫ���)�jm:l�{Vs��)=A�I�l��a���B��\:Pxt��vV��j�1����������Zׂ���n�T	�&X9��%W.JZޠm�Y	��f`岷�rދSl#�����Z�sl�YD���v�C�K�����+rJU6�	Iɀ���'���m�$�m�]ʷm���CR�Y�ӐP�x��`�J�Պ�@�j9"��X)�a��:�֋1�"�5���t��ژ+.A�6�1vl����اl	�XŶ�v�4Kߖ��Lv��y(R54 ��]�٫r?�;�1��m1<��Y4Xƚ�X��ѣ5�͋,d���,BF���e4�"nmӭ�A3mK�/3H�fLvL�"qcW�����`]^w��LR�C'�q��Y����3-4`KR�X���ÚN�QR�^*��UԵJ�� 0�X��fi�[��	��Q�%UY3L#n^�J�a��R
��"�f'��͸+]�,f;%Q��)F�Ǫ��FV�.ÎX�([�MQ�V�N�&�'��,��z�Dv�a4�+t�@K������u�;V*�i	F�Q���5�bb,V��L%��Ei�#���1=U���F�5*��H֮RFe,6)@� V���}Pdu��Ѡj(+3a��m�FԷy-!�U���ͤ���tfla�[`��x�:��i���ֺ5t�3]�;��5	Ź@��l���l8�iZ�U
ۛR@5�����bE�ؖ64��%A3�L�7M�չ�bUp�C37�Y��\�LR4�ì��(�r�R%��-ÄL�p=n�V4�nޚ�/	�j-��B��V.@��۹M��b/uԫ)���EA�]����j�>vN8̻���\f�����.٢�8,Ӆ�����-$i���q��,����d�[�kS9��b��WvtLw�6�EV��K�w>;��x�/�V*�L�]�K���s�^^	�u巑@F�(Z5R�9y�m������J<v=Ʊ�G�x*�*k��XT�W�|5T�W
�3V�1�rӤƽ�P��n���y�v�����A	F�`$���E��m�:nK#i9{&�G)U#��Ѡ兵%���(Sʕ/*���5㸀�]O��v������
���
��՘�K�������f� Y�;[#�na)1s�ᴱ�5�
Wm`S$B��@ 2�bY�O�ר=��5A�NL���+@��tt��d�Gwr̐4(S������Ska`l�����r��=��i�E�XF6�O"F�X�.�X��4� %dn=��(Dk3	�VɡLX5�W0Je��i46�W"Ц)��ѰjiY����(v�0f��P�+V;UmKw[>q��.�k�M�2�m�қ�Y�$�Ki<n�;��e`�7XR�� �=ٱ3����V١n���M��x�jT��ve�4��z���j4�)�ݰK�DC�偐�L�v�@��VCq^�[{SZ�NӰp`h�����mdU�����x�l�� b9W�2��2�6Rp1��Y{K �Y�lx43"�f����4����^�۳.���)�+9 �&�&���f�ȱn�iJ�}v�1\���%zh
v�#�YoH�:��H��m�/r�I�N+Od�F�n�[׍��T�aHvų���9�Auy�n�╏!t�4f-����ȝ�hS����B3^\��ܐ+ �@�f��t.�J׈�o��q:Pj��R�2�;i�P�D7@����lDp-�y�]�ZB�u>�T(���5y{J�!
O�O�HDJ���ͩ���Ҹ��,��kp[�&���g\����ShM8KOCE8C�ByP���j���cd�� �m;�3BN�9���|��킞ͣN`!�+k�A`�Y��5�W�de^M��Ry3V/5�ReûtS�NBF��-=:̛E�s>x�-��aۥ��>�d��EloN���35��ʦJg�5f���� Ҳ����|v�ws�2�j��۶6LʱCY�X�(�1�R5��b���x���4�,ۤ�D0�U��J����+�@^��]�P�1f��B����%�Y�m������*�T���Wj�QMV�)�Tkvhʅ*���A֙��Z���
o#�y�q`@S@V^iN�n6�.�e���@�*k�� �:�f��.`=S�Xl��쪊�<�#*�gP�A鲁�H�4(����(ɯoe���\���a���ôݥ��N�R@k/5	R��К,���Xt(��W���j�ufKmT�b�ĥ�D�����9*`�:,��+omҔ���ř�ś:��C�E��>��(�ڣf3X��ZӸ@6e���c0����t
-�5��:l�0�&��ȫ��2�j�`�.H0�A	V�^��
�o&�LuA�R�,V�Q��D������p@�h"Z�dD��/�Yu����ONkG�b�)��*H�+�/8kx	�[(h�s0��-@]�%���֠��f6�.��g;�����n,����-��d��jCmK��f���˳B���@�R+����Fd��,�oo�ۘ�G#r[O(aW7n�B!���c��BCI�u�M�m�XL�����V���xCeZ�@nA�l5Gh�-)�2mGE�a�t4��[�6��bIaञ
.��i^�y��M��i[��e�wLQHy@�3�����ìO~�ͧ���T�ǅVD�m�h�wJ��.�s6���ku�S��ys�ǵ�qia�!��TcT�^EQ��E^keУ{��������k�(Q+���b��t�*�fiv�IIm`ʃM�WĲ��;6����Ѻy���[�dӣ"����pV,6�-�t�Kb���ݤ���3/cհˤi�����E<,0sSw��ľ��+^��Me�G)�w�`�����q���i;��7J�"�=�U�zU�d�L�-�.�W0L��D7��!��DPз`��CM�
�,�gR�U�7x�fLĒ��.��Z�0��ǳ(Ҵe�ǷO	bP]HCP����,�8�P�`ͅI��5�Q��T��iѻH�p��2��kS�� ��,�Eތ�2��;cȑ6��E��с�Y
�o'��ӛtd�Y�^�JSL�ѻ���f�u,�Se�bQs�o`�v�{�e5��������Z�ۨ#�l�fR�T�u�,��k{���V���\�w� 2�Xb���ی�ء�U�M�ׁ�9�b֡m��U��%�eK"��p�f�łE�F��Y�Qj9��-�ڹK5�G77I�P�m�Ұp��w1�XIe-r�ҵ�x�J�C��Gt4��km��k5-c�V  dݡ5mm�ElMW�N�a�x�@M<�j-ݬfR
�h�>��� @)GS1G����6;gr���YZ�2ƚS�w1m���m��0$�և&� ʋ5݃����P�i*k^;י� �B�f;�[�ܠ�͎f<'v�^V���ZdԠgm}`1��&%���t�c!�,�Z�L��+)dv���Me��
ʙGI\�"�Ei�((-)+�`�ќ&�X��
�]�]�j�}�*&�O���n��f��ӭ9�ڤ�It۩e1��f���(�:�Slk� �4M�R��a��V�2bn�LL$�:���l��U�%���R��X�X�[�$Bb��#Y��4#�*z�28sBW2��J�7��NmA2۹p��\�ejP�(O������Z�mCH�q�7R��H�@=��5��#�-M4F1=ˍ�z���pU�r���-��Vn�Kw
�SbKR����T^�W���B��=c*�����֠n��2Ѽʍ��(h˙�D3$p�j��O.�*��L޽�������:�h�J�J,�h���5l��Z{)*1R�P�ph[�hmcK*�#8uR��AUX�me�fT�ZS�Ԣ��dSq<16[֐ ���꩘�G
��E����R�a,v�ͺ�l;�J���n���Vbh�f����cqV@�t�i"���uj���nK=Y	��"�"!����S�kU�1&mY�#؄B��	�z6Y/�sTx�A���n	w���e=N+&O�U�Rm)��CE���!�z�2`7(��v���"�4������Զ[����b��X��`��qb�����ӌ��@��P�]m�ŷ	��ER�EGg ���J-BVV0x����--��N���������P�^���A��2D.�+Y/,彺��	��,�{��p{�l����R����L�`7��pnU�e�w2�V��)x�$l�i�v�&b��l�lF�$�6⁙Q�M,���0��j�T0�Vi��l�(K��[e�pU끫U�����i��3�,fKG�3]�B��D2�odq�f����֥���Rn��\5&c�F ��n)�[{#�Ka�X�%�.� 9�o&��/E#���j��F�5W�S�)^+[
�v6�CCn�Xfjt���6(n񸔖���cV�.Dh��j{���X˵qa����l���VS��`	me���B�jG���n��QHb��2�3F�k2�c
ʱ�U�QؖCj�V�5��(>8�є^*�Ƌ����� �˙|����m*B�7��l��]�SIغ��O0�1r�Dv�0�5�)���,�x���`�!��ss[}��6��8cL�ܶ��h�nM}Q*��3�X$�Pv��y���#�Z�d�'Jqʏ&�j�2���6�8;(����ް0i܌�` J�{z�N���Sx��0�[ա�:\G�t�S'+�ѐ5J�ɷ�9f��w/�Wek*X��zd�s�%y��D-k:�ȳA��h&�'c޽�A�s�렩]@w_V'������q����9����R��-��7L'�D�!��K�>�9�%���j��^��6G�YF��}l%��	mq��ۦ�a��6o�R֭��g�$I��7�X��7N^"�w-n�{�:�'��[
�'�V�t��ue-W����z�f��a�E��I��s��b���
�S�uM����P���_�N��y���F����1��GŔke�̹��$\�<���1e�c����	�X�҆)|j�ɜUI�{I�3�+%N#T�4d����z
����:��7�$Mݝte��qv���[r�Z��]m��v���F|��cH!���Z��YiR��v+��I5�M��]�B��s'l��~p+ 5x;4@���;�R��H3/*�ݏI�g�k���W��O2�R�L��R�Yљ�5��\��Ț����n���j��.Pb����]f�D+3� ��Y��s�|*��e�4���\���:���e�+`Ե�z�T�( ���g[�f��{Z���l�}��b^�\�aZ�r���:3��Ǻ"k�{*�]z#а���7��tDw
[E��Oz�bW��iC%Ã�{�9p��p)QI;"�2��bv2AZ�įF�ӟ�f4;�t���
ѷ�8]���*30���\�9y*s|o(f}*"Fgr��í�-�Ԭ42���n�p�x�򡛜��.��;x���p���s�3h^h+�>���>3�����T޺D�����ӱ�u��Ѹ���Ϲ)&8����=���E>�Z�V�n���SZ5�=9�b;{V!���0:6���v8>�8�oX��r֒뻱��܆�˚���$���dRq��;9�4`�܎l�S�	�������uL������6�]��j-�������u�ni��Ol�e*|/��^�s��pK�Wi 5�j��r_���n���y��V��Q�z��T��W�|��Z�)N�q��b���۪�E�Z��]ۊ.�(��Hv�-ar��麜p���)��Zi�^o�D���n^[�ݡ���^��t�]1{�\�X�#�����/.H��x������<T�"�=����.kN�`^1 O�u��[L𬡍�}S���=����zB�|��slu�o{{I�	jP\ج��A��ӅЪ�9��"�Bk�S��*ů)��GQ:2��Gir.��C���qRO������<�Cy��p���Ꮹ>v���i��A�9V�ckMt���[Tua�w�FY2`AP�G�,��#�M�c�ؔ.^�s6��osEd�I"FC:ֱ�4W �ge{�R���`,�鉢\n%�<��ĥ�� &2� Jm]�5Lh���É[��]�TT��/F��Z�Ӽrӗ����Ug'ح���/F�y�9un%a�V��ҡw�-�,;�i�ր�+Z�����)4���)�:�;�P��3��௯�aø�9��p�Zܦ�V��R�t����w���W.6z�f��K�@zS�	�Ú�Hz�\�9���>Ɲ+{��E}�.�q;��]f�r�ewX��˦7�+�/G+\�+��u4q�`��2:�F�ǺhU����!���K��O�X�����(!w��07���xt	I^��u��C����
Ǳu����])���,��]cB�O3�SdU�*^4��cu��#��t�v�¨�S����޵��	ou�/�;uQ�q*�|}�(1����M�v[�-.�#�ό@
̎��L��q�U*^Y��Y�f�ڶ�<`��`�y�s`��9��	glp�]n,�sF�RK��b�m��n�iE�ĩ3Z꾻'����R��]�w�.1j��̒_�N��u;X;*5��mSIޝ�95_Z{��c$[�V�q��,����Gy��yژ��%�%Ւ3(]v䝭C![M�xU�{@�w5�s�v�����4��+{2�2U��F�4e�X�T�3�)�"��\�4�>�uȋ]I���v�'�ad�����u�F���x}Wf5�P���	j�v�׳e:�U��:��@é>rX2�\�ܘ��=&p����*r�:�LJWeFX{��}�]����Ў,K1�Ag�WWWg�WS�c u(vf�z�E���c��S�q��ŉ��8��;4T��=um�7Q��:��&�5&�E�"��v��c�R[�+�r���gO �����Zm�f��oGot���2���R�<��9���2u+��]����EKb����.�;%�g��e�T�^?)&{:w��_�5~S<6���%f�Xʛ���-vJ�I�fF��SlAզ���[aWR��9!ɮt�N\��dt@��0�ky�u�N8K�oy�������s�7Z��Z��u�
��\�lJ��O�0�s{��/�WQr����g`��篳��_>�c�Fm\�MN�����C�6*�����v���X���R�!�Cj��e�
�G��hw� v�@�n4O��P���i6�Rޯ(�ˮ�B��$.L���.8�վ�K��%ӗ�Ѵ�g����%�t�\37��8=���eږr
|SfR��&��o"Ĺ�k5��|�`��t��\���o[��c5�&�nqJ������,Dҝ��'�����8I�I���6�S�8������06�9Z�ofA.�Y%�̭�t܎n[c�k��Y4���=]qvT}{hZ�zU":�vc/��ŕ?#;9�μ*6�ոY��՗9��2�� 
'�+��v�֭�%VP޷������,�;����R����~e��zF���MZe��/�٫�Y�ic(t�·�.���ɛ}�)4TŷO	�i�#{]Δ��G��u��$5}��hV��2u\�L��8v!�26ӭ�9-��qu�
���w$ׯxbs/@ �J-��@I��+�N�1De�<hI}W��f=46_p������Q���5k�Kt��kWS�]�u�{�O[��J��N�P�{xF�9c�1۴q��2�1�8nW[�'h6�of�9ݶ��8�u�����,�r:�x� j�N�unAӔo�m�=0�>O2�5��l�W8洮��&�j�SR�r�D��K^4������������ۭ������c7��3�Ke����eC��H���b���[b<���|���	H3_f��5S�[�|.ґ/_�B��խv��B:!U���j�Ef�`����X[��,�]���y(k����	��vŠ�؏p�6nU�{|���2��e�"�ƫ�z�m���j��⦳&��k��>q����R���`�^�:=愽˰��e
��@�v�� �^�u��������h�^z�7~�tN�՗��h��[����	�d�v7;���\|:�?���HI��P���۴eǻA�0݋�k��p�Kɽr�X�PI���YCv����ٜ������x���IJ\a�X�� ��V�薝7��4�fԫ�{�wu��ɏ.T��N��\�E�S�e��d���9\ۘ��Yh�l�φ�"$Qf�����w�����+L����5^.f�j̠�� ��\'�(D��5h�X�����:r,����u�/����ĝl�Y�խ1���*9��*�`�+WM�/&T�P]�`̰�� �ZN'���k9����k��	�l�.������١�Y�N���O�	��t���n�'��V_�{+��H� �i����Y�)���@�I$Vp:sW�O;�C�ȩ�ߜ�Yʗ��.���Oѻy7דn�	���֝c�s0oV�f�L��A�������C����"���{�}�+T��Nb���-ޫwӍ0���
#z铪��΂m�Ckn�wz��5���,��J ��K��V4��A�䊓cOW@U��wQ�6�/0�}e*ܬ�R�e��������#i�yL���F�T�Sr^�F��m�W,�+]�E��r޾��08������N]��ӻ]��iN�9vc�'�gTy��l�c�2�j��`v!a�;ϧ7Վ�
7��� �r3��U��,&�L�M]�\#�u�q+q�̾cv�+ي9�+� ��wn��:;�ݷ�JE/�jzw�e�R�oVg'KJ����&�	=���%q.����R�&[\���X;6�&�m�"pꛢ���ޛ;G�:��V9�А�u|�� ��O���P�ꥇI[w�|��+@�Jve�R#�B�^��eU�2e�ґb55�"%��!H����T�+�-<͠�(��)��9��7A�i�^MN�YE���
��D�frﲭi�F�/7m0S�{���yk ��8��hV[��d�H���dՕ�	U��6u-`��H���PV���lh���sZ}�g7��sv��y L�&�A*�����wLe��.S2 �h��h��z����Le��y�<�M��urm`ř;�-ۈ�r�Yf9n݃ݐ��Q޴k)K�v+��tY*[�K��Z�_u����Tmu71h�ʔ��EmݴGc�)-������Ҿ����C���+h���R'����JL���2ΨT�B=.�\�g�7��k#C���'��E�Pe��c����no]<N����2sZV"Ѻ6� 3�q���`�Eg�ޮ��4L�]9gV+ޮ���[�&��n�[)=B���ݰ��S���Y֯�4�4�\4QS;��w�p��ai�R${�����fs��վ�.��Y�)Q�]Lê���U�Ӝi�.�� fs�F��.����4���n��+�B�2��Ī�dd])�i�5���H᧬qMCx�ØĢ8����̢�yN�m�i
��ڬ��ظ�3ڒ6����+�����d?=�b]|�6���z%qZ^ˢj���ZU\�(�A5��c+����z)�i�u�!���D���BP����];X ��3�\շ:���c�Z�Ɗ�4tj��t��M0u�G|�uo^��MӻQ���ˆ0���:t�U�ɒ���W�P�{'A��]2��B���:ܝM^<���&���i���Ǜ�i����PL���]0���Q�SK<�}N(.b�{��f������O%a��}�b7պ�)F��A73Oa��nb\�hk�c��]��j��v�υ��F)�lb���/y:����YL�eõ�����0�ԟ-��&��$=X ��,Ox����<{�=�S�.��}�$)�%@��� �[�fu����y[��-$�lڱ���"ܔ�:2p�j�h��Y=W�h�^Ԥ�ؓ}���[�V��M���y��JP��U����*-X�_!�� �.FJ�xF
1�Y���v>h���$�;_vK:m.�8�4Ҙ����JNB�MK�_uGc#��:_t�����eL*[�R��հ�W\�h�s�z�Ӯ�5�76�k"�	WhU��]ѧ%|���.H݋1����m��vS�9m	k�2-r��)RiV���v��%ix7팵v�ʜ�Ć���qe���>�I��֊�x�!)|:G� 2��v��=���.;�;73t47A���m� ��C=��ƥw�����]"��̣Ϡc�E��ʸ�G�,���Gf��{PGDk{�/��E.
��S�R'c��v]8�/���t~������H#�VrV�w,�y�mqQV�d�-S����:]9E���$�\�U�#h[ȥ�*Vu�|�}���ف-���%��Ω���2�RO�������6jR��ל�9�%�@��9�\�83$�eB!�7� ���Ԣ&����>�h�y��܀&YSw"��-��%����|MeM�q!���"�p�*��v[z�eMt���|��=sqT���ʙ|u\�l�sE%;I������!lX��|+�$b/�0J��1�wS{bu�!��wNZ�ƮT;�
����dE��;�{���ʋ�u�ǲ����>��>8��ۭԫ{&RF�}6��S��L��Ѽ�C��fԷ���--<���[cb17��fG�v,�
�yĔ���PU��x��9���rfm�5�]�G�m���K�Jt��Z\w�wM��N���jwhϺ��s�V�{S�Ԛ��vD�Z�uҐޥ��Z�.��U�u�s�lp!�_F�Q� em�U���=�����@5r�t�։�Vӫ�7M�ڍN�)���2��M���h.�6���vw"2e��]�V�����u�֓Y#}Ή��58�f�7��\�g&ijQ�
]5�/��|l�����2�6����-�.���־T��r{8�5�%F���ȝL�`�p�.c|8J9�;�w	�w�+���u��:��*[¹n��m��Q'���z�>J��Lp�v��1�G1��;�u�}�4�H�£����3�:�lk��Ћ��:;R��oG)�t���	�8�喞��P� ��z��$�!���tE<�Y�ͭ<����n��˚���Wn�_K]l;���#Z�]�W&����+�a�9�^f�I.h��R�n�uټ�Fr�3���	������sG��5�w��<�	��������"\("���Qେr����k�g^�����ˏG,k�Ƙ,	�i�bD���.��cqb�%���WM��V�!�K�f]�k΃9���	:^��`7�e�%��D\�H���-�+~���J������
��=�" @����`c �c����������?�]5M�쬼c���e�e�N�i@��;`��-��(X���Tˑ�X���n�U��{L���W+R�=��@���˲���2�A���L����c@�5l*+N�&�_q���g-�D��J�qq���]"N�ծF�P]�2�Y�h�8�q+쮮j[�2�u�С�U�%Y�)և�L��3T�K��
��h�4����3.��m)���܌e���i�n��H[}}��;`��ðV"�p�򃐼�R�¯q��΅����E��`�[���zS��1��s�n�8�|�v"f��isM�x�c/���o�\�]iо���v�F�����a"|������(h%�L9;2�/F�
��vA����W&u�Z��M�[���}rA�V2�ᇲ6��qS�S��9��֊��v���7�|��/06*�13j�xu$/�)�`:9��a0v[�M7���.��o�ǔ]ZV��u�<��<x��F��� 7��䫃8a\�txe��X��_�P�:wA���33>l�4�a���Lb�|���'gq��G�s/�/_>��Ø��.b�;���F��z�@!��n�L�s�5�(-ҕ�W�bp�ơwǻ2}[��[��v�
9��U��륢R�qk	Ja�Y]�;'wQ�@��X�J�WS��.��r���x�Z��z��]b�\z�Oj���m���Yݬ���%������u3�"�K+���ƈ�*9k3+��sr�
zQ΋[9����k3v��u��횝+�z�l��>
�9�O�q�"���Η�&�O}��w^˴�����u��u�F���M���'2z��	�@�ʂ���P!����s�1v,�es�S�K����&<:)�nP;c5Jr�E����8��_	dT]�7�of�v�wW�2��������9%R�4*f����-b�[��yH
90��׳����N:*sv�)�A3�	�ro�V��������e2
�r�n!Y�����6�1[ռ+�7��ݤ�� ؅*�r�f;[{+�<�A�u��[�C�Æ���GJ�\��:�@LWl��������F�Gs�Ρ����T��iL��#ʇ+v,6d��oF�!q�*���Aga�>��iSΔ��d�F�1�vv�[�a;f���犈�D��9[�:����vR��.

�n�Ҹ�*�{�X�5CJ�t)���#���2��k���4AJ8E'�\��!!�-����:������6Bvp1/1b�쌬�+J ���e�%�E��h��W�s�s���ݨ{�w�mXv�M�hvr���f��M���L�Y�y�"�c��Weؑ�2�q�\c�U�Q���#-XYӥ���+��-j<�e��JP���P�תup����8S�l\*�jk����Eڷc�)q=P���t��}������6�Hc;ى��u.��5�@p�`֊]6\kh-PHQ�E�س3(NN�"�v��9�|�E�#Z�	�yVu��)��o��!f�؂	EN�z�u�'�3b�m���Z��@�;"��K7��ܽ�Wx���}��쩲^��� {�ƂC��ec���Rw{n!V���[i���5�&���E=j�Z9�?b���amZU�pn�¤�ݎ��	]R�gЈ������l����\-`�e�]r�|���'ʺ��N�!b��U���Үo2ç��%"����1lw�k�q�T�&R�7Q;R��Z�t���:B-�X�;��7Fcx��v�	����
�r�9�.�Kv��x��y��̃�#Ki�
�)[R�vg��뚾�,���W}�ͫ�������xX�F�A�3�8��CY��I������p�_#�C�[/E��`���˄-,���<��C��Mn�W��낝�N_N���U�5L�
Њ��2�t�S0%I4͋�0��M	u]���nۘ����׶��ed�����Gf��o74�y4��/@����^�{2P����m^&��iv��\j� N���H��w���>�=�9�U�ʾo�uVܸ�Nypvc��UKO;Pw��u�C^�f+��K���89��M�G0x�Y�/G+�H�`�/��x�_w<��i�DU%Pt�[O���l�Krt4E��No-݆λ�!��V�E�%�.u����Ne(��JL�W��౾w��R�5v�p����Wc#34ZMӡk,�vJͤ�=�7��@vJo';IWJ�wR+mݶ`�2�B���B��u��E[���ݝ[L�jƭ@���EW�"�i��Hz&�V�^R�W�!�Yu�*!-\!V>#��`��SEN̰h$3�ʞwM[��^�	fuF������V�Dz�G1���	,s�>��^�ݴD@^�od7�:�J�cr�U┅��Ɩ�mm�S0�qtC���F�Q[VvwjQdJ��=VB�!�7�E�g}<�h�ʚ2�R�X�]��p�[W���F�������X�c)J��S�I�t)8�Ċ{� �7�v�]��Ǎ��u+vЧ6ѣ�N���l�fb��p�s�g�J�9x��� �-֎y�\o7$���k�1��1e5r��lE��t��a+�GJ�!����a|6k��8:���>���Sn1���Ɓ�\��.�>'q��%p,��u �V-*�"vB�Eu=��E�$S!�E���W�l4��kJ5���:�����5f��$�r����D�%�)\�ݽz���2��W}C�&i��s�N�v������|d��No7����PM�1�=�Z')�6�ι �
] �ށSx�k�yAVs�z:�,�n�\�����rk/RcNtϮӼ��*n�sP�=Y�ʣJ��c�-�k/F�	�Mp�C,+$��&-�X�Lgh��Ss.�D;t�o�ՁVRVe�J�^#D�Fń�h�oMv��-]p>����:�Q�cn���j��j����m�l��E����o��P(������V{��B�w����邦ģв�K� F�gp���U��9�r��כ��WJ�y�3��҅�Mڮ Q�s��3kU�[���U��a�Ntm̜�T����@v$:�F(l���8�)S.5y�^LweC�9sܰ2*��5��	>u�0���-m��p�tr���a���u�����
R4�B��q۩���p���2��n��ĜAG>J}�����Z���M��������r͔���dj�^ �g]����q�aK��I@X�n��;J<��ٸ6>��b(�f>�u����c>yVq��:�~i�]F�y��e��K��0`�6n�Yl�kkt�F��O�Na�xqK�eJ
�u�IWP㸦��{y�B�mI6,��spuљ�ɖ4p���oD�9��+D�yV�S�-�.��Ic��Ɲ��+r�8i+��r���rhBejj�� ��Q��3vN�{y̳9�������]��R1�A_U�����6�O1V�Sj��t1��n��+oj����Y͕�Ctfݽ����E�[��a��f6W!�˧�Ҭxz��uoN�|\�ݛg+�u����rq�R��T�\�g�Ŧu��%Pos�.Vᥗ�f�AZ*�koK;3rӒ�'��Å�m)��&�5t�1�����dޘMٺ{���ֻt���|&��`����)��T�T��1�}dZ�h���4Һ�(媒����6ڀGI���
�d�M�]d�� T���� ����*o�+e�;tZ+p��G���պ�̝�ƒ�qn����0�KꏌΆ*k��um�)3�
�K�Z�<�aZ2�Ac�Z����=ڍ�
l�K:aM�y{N�J���2��/S����y���]�wI )+q�E�W8��%DK�퍚(��ݶ�����Pb� �K"�#���B�У�v��&F���s�9�e�N�S]Ѣu�����WHC�+G(�d���Wr'�uu�K�]DN5�{�5��1$ٔ�ꕹ���Z�mw`
u��� ���#f,��?�Ŕ�Q �ѕ��W�����b�:ىJ2p����'z����;6Ц����_oJ��8.��>��ERA����NwGz�[y�fi�(;���)�ӱ�G�VW]�����D��,�g(W�X]�R�y[���gH���"�EW;��N����!�|	]c�F.t�9\[-�ZSRNy���hH�
��]퉄uby��6q�C�oX����a�A�Y��ͱq%��LF&��ul<:C,�X=8�۬1�E�P3�C�A�F�� ���pf����@���)����]�s9���n�4��h�w����ྮ	���7M�t��{h��r˽�a�Z���$�c.d�3�nn�(����'F�ؒ�x�{*��<��|��{{�K|�B�1&�f�H����6b�b���n慲��^�7l��R��Nm����:�!:Nf�[����wsT���e��Ni�x�J���{O@iۮ��F<DM\���g-$m�c��;�[4[P&qi�fwQ�y+��m��拥�Hv i���k�*����7��n�k8i�2�b':�$��㫒3��}�e�[[ǭnΥ\�ܝ��rGm1���fr�ɛ/Sm����U��;��(���hbĻ��H�[k{Yf�Di�z���������J��^l1l����ɘ6�_R=�jM�2�LrbU �7�ҵ�Ξ}�v��QvA��������@jp��lj���dX�Vl��S+�xg"�X=t�=&━��Uݦ&:��t�f7
������f�wk1`���R�cUv��[%]$*�n��Nlj�o�0`7�z��e2Z��:T��jf$�>�͢�M�V^��ӺCL
������,�'�c�C�."�л�oA\T�7rEc.f�QWqw�Pu������8r�%.�+r�wCm�o�n �Z�_U侊7�r�[��*ow��lyg���39e�żV�@YU��V�ᓜ#�{�����2���P\ �.v	J��u�}�tS�.��C�;�ۮ�n��uo!E�
M�V�b���iC���uo�+Eu�ݗjn��9v�*=yJ��L�|�
�}a�6=.,���2���m�{L����0wk�(\*�t�v�|p|�b7HM��b��]b�PW=.��U�Ie��z6�f�.�+CQ��6f�1mq��"浬�̣:�
	K��pC!X��[K>j[nۣ-�� �b�&�ɸ�:���^]y���j���g-ܵim�i-�i{+l�N� ���x��Bj��w�&�ZH�Rm�R��p�1�	K8u�c�qJ��E�Kh�J��{u
��[/�l��}j��m��*+���Т��ɩ���&>�F��NC�F6���8���%�	u�diО|07�����%q�2����vq�-��I���-���u��vլ�ju���� a�!E��8���@�b��T�`ė^V,�p�C���+��3�Ԉ$d����x���v��GU��=��Vy�Fp1��,I�sn]v!\�!�f:e��u��J�T����mB��\��I��gu1��r��[�[��{����1�]��J���_ʠko� �t�Q��:H��-�u1��o��;H<M�2�᪐��M�w�B[����s� x�S92���NP'&�w��;�U�"��F��rgn���N��\��h<ٕ��Ԣ#]�<�^��Ʈ�N�fp?�Ns�ѣ{H�զ.����Wg���C��k�t�i���/0i4Nh(�#��'^2�	�d�y̬�c��F�	=%����yv]Kw	�:v:���������t�ޫ�Ҵ�ks�6F��';Ν�;�����uaVe%*��XԍEb��=��+���{��s���R �m�4�{{w��kή:���k&��r�c�E���ۻ�Z�
�պ�tU4�py��:9w|CL���ZE�@�u]h&�q�?�Z�o(�27�*Ţu�ͅ!L�BF+�Wr�Ll]{��u�/��M�K�9[��Փ-O.9[Dkr���}{SsC��� ��rv�HQ	��N��9�0̛�k0�1��4V�f*��EjW:�ǲ�j�,Ĥ���<썛b�:�f#څN�л��P��}AA��V�Ñ��#غº�[t��e3ʱ���+2ulZ���ٽ�]l!�_$��Vj��{	.;�GM���.;��O�ƥ� '��'Y�I\�1�,��.l�mGov�j�W7'�n�C(�5R��fG������j5��Yg�QФ�l�)v*�R�L(�'#���@�}է�J��vH����%lhHSK�;����J�c�bIvp��aG��[\s���p%]r��Y���$Q{t��ܓ�aS#p��+��3L�z�v��B�l�e���hL˺�&����W��Z�)�#;M��Y)
��Y5���'������p<���vWf�����VƸK��s���)8��0i�k;�͹�����8V{.�tU�D��*�ļ��Z�s�޸����]�A��F�X�J�4mG ��tŒ�1u'r�қoQ�fm�*k�0(�mG�U���u��E��2�=6΢��m�Yy`����Ŭ\D�|��dFP�a�)p�P����+��=��\Qce�wO2�R�P|89�K�X�����n̸s yӶGz�T{6&�f�J>n	��{.ˌ��\�*$���,�Z�+�Ȱ��'{����8Q�C^�5��B��n��P�l��\�h�TCR��y��#FwL��+DS��)��V��:7�8}�c`�t6˟Kn���;Y�9�&��Xh�U{&��c�Cq�]�x�F��cF�XZ�&��m���m�r�M���y��ѓK���S��)�y�a�5��<`�x2�[����J�k���i���VHІM�8۔4�v6f�\̒p�e��y�u��K�=��D"C�ཿ%o�(�Ǹf���@�B����s�s7PZ��.w��]m;�YO3��؃%H���:���+�y;��.�_7D�m���f���T���lm[��fo�,·eH����ӷ�l�{]����rH�.x�?k��7��,�'�)xG�Hk2vw�S��_�aȹ�t��=��%�H�	Z��;�ESl� �����#���ͧӚ��g�+R1�TIԷ@���zn�IH:�ϲr���Xkn��t�p&��(��Jc�z�����h��Pg]��1��m����� 3k0�RK(ugR|��ƍu0ik)�:]�"�wm�i�b��8-mrs�y��o�n^u�)�֑g��0.�Z�zQ�d�KŎSN�W���<�J�n	����YՅ=����{�K�&�j��/�c-N&QB��>��i�R��]P���K�s��@���o
��ݵ��R��y���`�ޒ��_����ZFd�� QD�\�����R	�S�#9��݇7h���^s���A��
�1Q�F���}��v�7]��2C{���L�F������]������
��*�:e�p����V���Y��˟r�к�.���&�[�*XܝG-Q�Ԏ�U��Eµ�yy�b�}X���;��&zaA�L\�d��إ(�R��5a�5r6dZV��Gi��竦�X"��WL��̈]p�����*���z�lZu$�s�q�D8TT9��UH"�r%"rsvia�U@G"(]�(�����8wt�C'=Ԉ���B�h\��j�P(�i�z��E�*�.�'Q2��]���9h��ҏ0�XA^���t������9Q�t���Ȋ

ui��#�'2�exb ����9A�r�]Hi���ia[�������$ʇ��պ!in����绞�gK���P����i�ݹj.�,���T�uJ%�A.��B.���(�0��%�0��C��A����օNl:t�R���ңA��hI�U]nExz�I�df(�w9��p���"[n�H�f(h��
�D�4�#T�LC:]+���š�[B�iH�H��n��Er)$�]]0ws� ��wPL�36V���UԓU��E��$�]*D�J
"�**�y'$�$��tu0���s��z�yД�R�� B(�O�&�:�58�l�Wnv��<ew^He��J:��N��&����G�3\�ձ�q���6��$��okU�9�oO-���g5ú�Osh]����߃�ʡ�R
�WZR�h��޹S�ZN hI���G}�OpwuY�꾂�Vl��3��m��Q��~y�VE�}�8ՅW���0�'f��ur��D��rw2�V�9��� �}i\�^��l�Z���֌;��(
�����/}��=U9�❙(���С�:P����k��/���^}���ڵ����3ږC��d9��w\�_w�ܓ|s��Wi[�Fb�6'��d�׳yʱ�o��ٟ�,x	����������]�=�3�s���*�(/z]�;�t�?=�_�_oD���'w�LY���C'�J��D��vcǹ#MsU���t���s�ˎr)�«h�0_�G�܍�Qi'Gx�����B�B�5�Ҳ�OD�ZxQ9�6x���θ�!��[�ܮ�r4��:�*��3P����VT�nc�oF/����v��ʩa��p�Oc7
HJ�vU���B'��L�gyIk_{Ӣ� 7PI�$�q�{�q1X�DE�}e��)�h\ѯ�����nsi��kvyŻE�������a���Bc(k�x��Y�-�����N�ml̚�.�]����;�c�'(��f��.�q�ݧ�*�:��` ���t��N����w�l,w�_��gd�v��g=V�>��\+�Ph�{D�|��B���grݡ.(C`M�SN�H邹ٓ;�ȇ}Nt�vH���~�c�m�{l�p�=>i(�;d�5pz��2�MY��*�SQ���3�e5�vv���\�����Q�<�g����UT�g+hO��m��J2%�u+ۖ�כ��Y�Pˆ�t�v��al�η�����]7e_At�8l�dC�r�SJ=�~��7����M�_yKf,/r��@�yz��/�n*o������d��U�P�¯��6�G��@]����x͸_囐�y�F�_:B���lt���&�*��ˋ�b�|�zwn6u���͜w��O�&�s�cq��7�jP�Y�e�փu�3��/�|�pd|�H��u���di�S2{]Ü�)�b�;,F|�\��p�h�ԩv�/bV3��N�w�V�t{��EV�.�;tp}7�օ�U�y�U�4D�6�mƢ �����[�,���[�R�hr�W�)���KR֦�=Ӎ'x��Ս㒫��\�C��5>�t3G�2v5�a��o27�	��&�د�wY*�f��ϳ�枅-�%�^�Ho�N��'�����ۮ�3����\A�y�뙜�T�v�"p�5�s����փ��^��z*UlX&�[<O�ĺˢ������cn@�O2d;�>7�>,�noA:�F�`3�XG���Kcw����Qr$�'G�KO�#~j�TOǠ��gs�{������Tm���.'�y>]�\u��8����E9EaL��X�J��c^i�.���M�ں�y�vwn��YQs\���\:3���P�Md3"؈��*�b2�5���v�pyU��q<
�ٓ{29�yt'�:��hؗ<|o{m��tv&F��\��s�z����޷7�kރr���HfBn��XZ��2W3�y�A�-��"��t'�7�;ow~�6�P&����s)�j$�b�u�\b���%��l�˹nm�7ǐÚ]n�!�[0����ux����e'��md�(��j��@��؄gW��>�;�5<\�C)���a�#�����׉�9>I0�J�ժR��޾6}����P�} l�����\2v%�f�G$�
�G<�q�OpB �u>��γG^��0J��ඵL�}�0��L���w5נ^���C@ߝ�j&S����h���bU{��ڻD���5NJ7S��3d�J��ë�uı%�¯�"c���u��(6��m_R��pSR�nf"Gf�P#�h���!�{};Zuq�c�&�f&�����ڌ��^�nv{ʶ2C9X����q.f�}<L���	��<�7�ow���7�S�qe�ֲ����x'�
��l��>����T��1���y�M�'}�'�7݊#H>���Y#B��ڰnp?Pok�g�O��+�f<���8���=Z�d.7[iv��bh^*���Hd5�����8C��6^
���{w� ] �$>4�L��ҍJ;B�v�C�we��MΡؚώA���W����6nR\-��س����<�td�����ˁj�ުs+>��1I�#bZ`�#�!^��$h��0���[�]#Bݢ_ks���>�T�͚�Ȭ����E�]PM@�:��a��Y�tV��itՌ����[�s�Ud��h�Ԁ�k��]Q�[9��]�#-���w>�s+�C}g�F�ܬ���j�ߎ�tegӔ�\�u
`#ڃʖ��{v'��]�)7oG:x��\a�g�/NѺSB*���Q�:�t
���d��(�CC��A����Q�� ���
��l�;�؜�Hek ����޽֬�+eh�ur�4�ub̽�v�[]�4�6xS��{[3�{�;���F��agE9��a�1F�S��lG�jtrvV��)���6dg	�����`��,�f�-nc��s��˙:pO	�Հ��;����2��Z>��jY ���F�t��T�����{μ��핦�Ԭ�St��1�>6d�Rx؍J�sG��t�|:���s)�2���m/��K:�^�'x�;ڟ4E���l�2n��N^C�?u�G��Ն���訅J�7��|�a}��%]P�����+ʫ�z���3���#����%l9�}�G,�v�+I.=�f4��PDN�K('q�	���F\��p�����{�e���a�q�r�=Ӻm���ÀY�[�����x�`�x�zl����z���#�d��s�&ޓ
�1���Na��v�g!���M>��Q�
Ќ\6|-}���Fx��LتO/�G&��Wp�Sb��n��̎�5�o'���N،�b�FH�|�!Kb'%�mFd�OsU7	��nV�;�c뉦��L�k[v��s�����tޑ�n��}�����03k���Y�ʲ&uH����A��va|��,p
oM�B�w��y�x��f)lt�ɴ��8��UaT�����<�����OY�Pq:Y��5ՖT+�^�\�}�ݽ\��A�t��x���\�a���v�v����`��"ͻ�&<Ct]�0J��i]�Gu�A��o3H4�����p��{ͬ��cY#�4Ee.��`1I.�VV"��e�[tՁk��p�,��;��R�e�%��Tb�%�*-ѥ18��e[%�M���+=m�і��nF�ȼI�F����ơо�!p�fB?:!ʕz�v3�f�򋫽��܈א،�j���Q��&���'��k���^�Ƕ�RѸ�zu9�����75p��F�I�ڽ���a�	SL+W�Љ�f6�G��>�o�{]�o[���z������׎���;8W<Hw����V�>��\+�h�6:'��ؓ�����BI��N�D<H�L��1��*ui�ئ�D;�s��@������̙�{^�Z��F��qv,y��3�.����Vұ�#Og�T1���|��-�����t֧��ѓ�@x]��;�A�7�T6�$lK��V6嵴�G�j5;�U�_V^�<�14�J�ȹ]�\Wx�q'�l��ꜩ�ҏ{ŝ_/�c���l�x�,y��>���x��n�r�ppQ��W7�*,
	�'9�޻:E$�!��^�c��=%Q��{����d�qj�Q�0��P�<�j��k9� �l�2��FQ�^�2�	P�Z�-��+<o�¢I��ܮ�-�ڳ��`�э5ۋ���fe
Ѵk�SxD�y�v+]`R��:F�smik��;��7�H��������`R{]�A��FkB;�m�QOG��m�߇K�q�7!jO1d|�({\N��g�}eY����tǰ�[�i�������SFN�q_�J^bb	���W��8�]W��r�S{mjŘ;�]n��YZ����>.F�B���ئf��wr!
c����@�R]53�ŝE�z���k���ГW�̅WYg��(�â�x���aE�I�We+�k\�x��>'�Z��{�
�lo��M�'���l�ړ}���9U�	�QE(�mr��7_J3�j�'&p TXg�{�98��wd:oJ���I	KOT�.��D1)�K>�y�vu���T�n����F.�*�2�Иl}�"��FŪ9�6t�';m�n+�Jr�w����[���ݺC!eE�_'�~�p�N�2�&�X�Ƴk���v����	q��6��;�HMJ�����zzz�1)r��?T��p����t����m�g�������l�]��RMx�{0�d&��(�'� �F�y�b�Ou�!K<<9�܅b�s;O!oO\~�U�ٳ�ms��mm�^ї�\-{Z�h��4e ��~�3=Z���*�D�.\/�+�e�g����F��E�_&9�2��Y��jD���L��Y;���C�ӵw���.z��a�����0rJ�Ez��:G8�Z�i�ꝲ�{*�t�2�NwQ%� �7XU�R�v`�1�\N��7pOj�«�ԯQ�~�Ԑ[0��odd&�q�L
�U �\R�$`�ZD�o60%!{ʙ�oSR��p3͊ldO�vfat�%�͓�i�ɦ��!L��=ļ��UǴ���W4Y7j��*�57����+{ԏX��R�@m��W� gYuG~y�0�������}�'��7 �_s��T�]X�o��]�*Ꮃ�����p�����F<�z��Ys�fw���9��.��y-�>��b��[��S�Gs�WNz
�sjl �������]�[V8��:��~�l�
Y�m�0o��U����-U���Tmc%�>�8m]�ҩ���0 8j�74�����M���r�ӑ�.^G���m�4�Qt_�j���gg��ʃ:;�!�UX��{
��؉��95q��p���6n��r*��EJ�Ja_��}^R�G�z��8!zǵ^%�t��bʤÑ���b�ʰ��ђ4� ed��ͧ`{^�Y���1\�G^�(U�����rc����YK#�#-�>�F���U��$�b;��s���,˘����f㚞&�ޫ�ӵ����v��9lGo�$9uȞw$����V�n��4�fw55Q�|9L����ZII����7�1V�V�@��uA�c�8��3������P��dBt�:�̳�74AY�Φ�wq�ԡя�:�Z����0�i�u[]>�Cr�z{�ǆp���@�<WDx�+�&�;��J����᳂�X��D�!_e����E�����Y�� ���"u����K�K�v�X�m#�T:��-�$��E�`�)��<�����ff�ɫ�H����v&�x�	�㸽���}֏�t�S*��n)ؖ������������_KB��1��q�ٓ�I�b6 �\ׂ�"�q�\���r�ݺ$�{u��Y��%^���P�<�\�w{P�/����T�m`c@�@,�]�}� kws\�Gj��� �MT7�G�T	XzU�z���<��<lژ��|�\���Iì���W�I&]�Y�����Y@�/��%�f/e��S5�Z����&e��yȓ�=�a~Y��\�D�Q�<N.��:�l�Zs
�,73��l�A��.�9��[�v��"�⮙��R��Ӏ�P��8,�0�'���h�+�!P;�cd���'s��M�]�Sm�қ:K�Ɩ�7jl�������eub�j�5���	L����u�.m�6mV��T�B��Y�A|��(�2Co�E�ڔ,�*#:�^�Q=NFR�`}볧�f�!�i�W,����}�.ܭ�ǵ�-�yFm��(68�c4�ϐֆ}[���v'l�b�в�ai��&�ϵjp��I�m;~����Z>��=Jd����]��s�;	�L�j��s��/��z�*t����c�}Zh�Ux}�x]8��_0<*��M�,T�����v��Q}�es�C�d�i|�Z�}�=+ӽ�\:0x�W�5�0�/���s����ϼH����|�����$�bf5�����?{v_��ϔgp��Ib���)u�#�P�M.��n��ф�p-�՞���:p���א،��\s�7Xv�V��L���Y2m>t/gz[���\\���e��\ ���cwڼ7���Xa�m��f�*i�*ȂU���*�����9%w\�6>ϗ]����a�gg
����~��L,�u��<��k�U�*����R2%Ď%��̬!��ӧ�=�������Ә��Eᘩ����g׭�-e�X5��g/�s��/�es�p�U���A@`D־�P�B�t��`]0��l[�J �)�`�����!����.\�&���\�oةA7ޛ��b/���%�k�� ,�G�(��
�DX���������4&��Xh�mn��x�*T���9�=����jƮW�k��i�!Әju�ɏkiq=���bY�Md��K��{B�C�Mb�wΖu��:�'m��O����qh-c��2E��Z�%E¹��`��d�����޳ϯ��mǔ/�7�V9��u��n�L�fT��Rr�*��L�����vlz��\s
�d���(��'2�5��K�乷��S�[&<��\u��v����#'�us���wk��2-�K?{G5�Y�;g�����:)�^3ҷ��ŗ���M�k��<|�1�{׍����AF�qm`�ZVp���V�3#��3�P36�34�=@޶u��m�O�;L�X��N�Ϩ[1|�F$*��nH�b����0�K��/)�;(��<�<�c�|�EU�zoh�C,ǲJ��jm�.��.7L<&�c��『�x�u���$\:�Ӣ@;uaV֙b@�T�׺;�b�[�Qf�����&􁪻��G���Y���	��uͺ�v�а'}1��^�-��q(���)�(��̷�i���[f�&\���Z��i�V�WiL�Qy�|&�n�,��B�%K�{9��T�!���V�J�E��g3N���N�Zk	R�:����Z5Փr�,-���d�qk:�LZ�)m���^��dz�_K���m� tu�2�G�_nF,G���"��5���ׇ�������������"�]@�[��E��U�۴c�\'L}\f�Z(�Juv[�g�}���a8�kr]��u ��p�N���]�w\�V�F\b�q�D��.V�d��G{V�"��u��ތ�Y���P�|���69RI�zT���*ʼ������y��0e�������dњ�i�������quI������]dr&��=�:����iﮁ��L�z̵	�;�,J`��3*��<y"Еծ|x)zK̚:��������9�i��a�:r㲓C{���޾y�<1kb�Ӯ�]����؉U�+���d���si�e���l��f����U���]��z��Eg�q�]3���,���*�R�v`L�Q��j�귓l���ࡵ��ۨ��W�kwZ�h-b���	�;2��6;4F�o�
�4�]�X=��ǰ��~�ķ�wS�+S@۝uc�`�k��$w�EX�\�)Ϟo$E� c��
�]��RT��������/�On!fV�;�����k�����ȧ�Yw��o���v����V=̥M���k���#�;�`^���`�ƫ�� LT���y&5��r�c�����S�@��$���JI(�E$�ܫ0��"z�IUm*H���KJB�-�II�����fQT{�!AedQ�"��aem�J��s���Q"U+I	a+��g+EYD�c*�urnzbX��9��F���c,�%a�DDk��B$��s��j��I�%�{Cs��p�F����Nbi��.l��rj��a�J���9M�J�I,�J�+�DG"�(��y��Y�̜��B��Ĥ�;�p�X^��C'+�2�8�k+�tT5�bXRB���"���";�紒��r]OA�N��Г���"#�E�Q���	"�]7)���54@���T545�]p�V�#��SI3"(3
�DJ�Uq��+�XF�Fa���AT)�
�-bd�P�bJ����)T
�,�H��k<¥L��$�C��CE@���B���̭��&���V��ѐ��4���w��w�kN����K*]�feg\n��j��N��b���B���ö���3/����F��K��w8����Ǉ��U<~�ȡ'�97��u�������'&���o#yC������>;_�}`�8��9���b i����>1�!LA�I��0e��:�j���Y=���1>]�9S~/��ސ��ܝ�����]��V�~���=&xI�F��|q죕����d�v�N����<���S�|�;�}q����|���&~���qߌ�k��N�U�Wc�@�����~7Ϟ|'�nv�~����������������������zBI�7�<�~���;�w�x@������&������
�\x��'�=�V�w»n���xx̥9;���bHbH@�$��`
1�����Ti�®?~���7�'�_{��ߐ��÷>��ݷ���q'���v=��zBv��|�rrnw���0����xI���C�?F��s���������;�Q��Y��:w�i7����?[|w+��{���]��M�ͯ�i�S{yǿ�{zO)��}����ӏO�90��wl�����;�~��x����O[��O����;��D��	!��d�EW��\ߛۼk�T���?Q�����?8�Q�]��@�O<G�oo;۴�C��y��9P�����7�'��x�������Ǎ�?��0��}����h�^r���|��	��������˝z+=����*�~��_#�o����yO	��!����9�'�޻��aW}q�����~ǣ�xL���ې�n��;۵������oI��:v����������n�=�G$��df��kM�������羥@� ��Lc�"�Y�DF��NF�n<+�w�V����^�z��~C��!��Ǆ��{w2~w�<&w��=!�7�$�N����o�rs�1�H�F09�����\⪊�}y�}}�_Qg�E�~�O(�"H�>��	.1Ex?�8�Y 2#�@���v�z��V����y�M���o�^�G��}M��y�����]��-��͐$�
�s_��!|љ��WK��c��LA �4�@�����@F8���$�h}1F�"~B�d��U?;_#����$�����*�ӷ����ӷ�������'$��$C #�@������g5Xjhr�nj_�@nG9c��Fx��u���
�@��/A��ƐX�1jg
��;CO!f��Ν��t�<��@��&T��oh86���9A�s2�<:�;�7O��U$��gՌ<CV��7wr-S���W�����q���H�Q"��OZ�Q�<����x��aM��_��~v��~�I��'�ޓ��v���r}O�c�S
�9|8��8?��A2F�� ���<��\��]��{��{g�8��yO����n�� �C�BLG"����"$�"ù Q�F>�� �� ��C"<cÐ�H�a�B����A�Ű^�]�#˗��ҫ�?l�P��(I�!!�}��#r��C�[��N>?~|&����@x�q`z;g�"���{�������~t�NӾ~��<~�����Ϊ���s;��F��Ӿ������M������bw&����]�<�}}PzO9��&�P(
(~O��ׄ��1$�~���;rr��N��۹Ã�bȀL3�v�b�@6��R������n��޳��왟�����ޓ�~v��~�ǔ���ܝ�{��Ǆ��?8�>�'xw��x�m������s�j���/�?;I�����i�R�z6d
1�3H���tY
��ey��?y�֧w� ��0��>ohA�0��}�����\}C������pI��~v���<;ӵ������ohN��~���bM���xO�����O�@xɍ�$�&�DE��h�¨����y�Le�O"L0�6��C"H�^�������=��'&!��ߞ7�~w�9�����&����z;���o�rs�=��ǔi8������E"(���@��F�&6�U��������ւ��و3D�3�>��O�?|$'��<�];ô�=wc��o�s��EcL�������}N��n�_?~������r���o�@�>>�,�� ؙ���|*�]���g��d��-�����dD�1D��������5�	���.�F�&���o
�Nӿ�ߞ��򟝿�w���
o�O�o��}x=&�P��v�SϘ@FO����DQ��S*�?\�_�s��t�1�!$"����ь1��(�A������o����%{O	��S�Z����raO'�����Ǵ9ǯ��>�&_�������'{v��b�E��.��>\��ݝ�9yՇ	�P��\�u��\�y@����/xt��v�[��Qs��V�|��Z7ax��s��D�����y�.��/��U��]�ۭ�9������y��9:��V�m�|�N�v�%/rN�,�A`dᶰ�&h���\�!F�ie��c�6��������|xD���(N7�����N�^��~���H�y��pxp�˴����='�J�ϸ97���=��]�1;���'���0���<�ۼ���޻�o
�Dah����c%���3i=�_��$���S1 �FUP$��&��M�=��ǔ¿���z����!�0���yO��&�����Ν�Ǔ�<&������X$�]��=t~CǸ��?V^N���o��r}�cAW�T�~S?��|q�9�?�r~��»(����>!�0���}��˾?�s�ۓ��޾�w���p}C�aT���X��7���(G�nW{v���?'��oo;ߗ��{�<�p��F���|�>S$���(�����y���;�b}��?;y��?����ڣ}~��|eߝ�@���xM�����G���˾����s�"1�ib���$�]�f���򜯳=�^㾳D#&�$��%�A&_��<�c�ԝ�ǒ��o�nM�	�y�÷~����������3���yv�>>�����t�?�_{
~O.?8��F�ߓ�r�}��������J�z�y5�����G�'�10'����������q��c�Ą������!޻��o(Rw��\yq�>>S~|8�z�Hra_��G_P��"�������fm�\�=���^�,�Y�U�f*'��'A�4����~߿w�p)�;��xC���?ՏO����;�Nq��u�0���qG���&�<����x���#�Ȳ ��}���&�>��A�f�~�&��@� H�'r�/�� I�;�
H|b$�`{>�dI>�<�=��㷔܄�;��)�\
o�X9����,O��N�m�������ڠ�}|9w�iSx���K�)��o��	SJ�羙���EO�~��5~���$W}"8�"1DuW���� z;�ߓO��w���<PI��=~��y@�����m�ۓxO���k�����
��ǾA����ߧj��Wz�u�y�w���ꟾz����p�]&���o�����_{���@���E� #�=�Ő> ���v��ߝ�K�+�HN?����yL=�z?G���v�	m��B���`lժ�@3,�k�����|$�b㥭�۾|e!ٜ�wR�9	sx�v����(�d@̷X���Ï���I"˯a�T����L��1+D6AR�lE։Ց4,�Gt^�9ܶ�ΔF�!�T�txеE���Brr�̻��׻���u��4��$���Ӽ!Ʌ~X�G�𛐐9/��o���]������GoΝ����o	�!~�����W���~}���o�_c_�ɾ�\s�'8�����㟏����Oןv��ϻs�w�g�� LA ���	�ſ}����s���NL.��Ǻ<|��L/��q��~��w�צ"�b$�a����wϫ�$�"#�>�QE`@}ݚ�[�b�[���n�U�8�όD�>QB�1�!V�ϻ�)�ޝ�<`��r�v�,ro�;�![�F'}O���?&��S����|q�?��C�y��c�!0(�bD�D�}�������?�w�����#��~QgnM����s�k� y���&�����߯w�Ǵ<�Ӵ��ϧ�.Hx�o	�''8����\
o����{M6�a��Z��4�1'kp��Vϸxu���'?��}�������?��߽q�L #7&<@� B=���,��Ͽ?x<��I���������L+�o����SyBM��~��xO��T��$�v��P���������69'?ݵ˯n��`�+�W�� /!n�8��&��$�� �`q`{nYȀI1uU@�� I��@��DI�>�Ȳ �:5x�iH㐒H�R�x�'���ϧ줂��k��~���� f�&"I0��%$�I�����M�ޏ7�۷��_3l0;!s7�o�ǥ�+�0�i�N�L}N� ���T�v�I���]݃\%
���N�\���8�ޛ�~X�}3/��.�(�lK��E�X�\"��!��kq�G��٠�]P��W2�ė�1�;ǅ�1��*�ꅒ=��ܷ�xVw����(�[��l��,�[ȧ1q�#�n)�W��ܰ�������mֺ�eK/��[~}��vu�4��)<���]+���ݑ��ޥx:�����v�:0�;Y�9�o6��9�W}tW
�ц�M�m�Dޣ\*�������\�I���ݶ�of�^�8u0��ڗyrC�4��[3/V�J2j6G�� ���9{��^|�2�G�`0�Zxq�%�aˊ���	:�=Ӵ����w��8YvD)؅��.jk~䱐X����2�����'�z��+=�|��\z��'$ɐ\�)��/�[ʬ��]�J�S��pOe�,���h֍OBj�E��fw;j��a��j��'8�F��ɝ�9���(<�ӧ���,���͊��s+z�7˛�K{�;��O pϦ����Z��Ktg;մ�nF��@j�;g"g�r�t�ɪz�{�iU���	_$,6ZO�|N��4\��PڠP�������7�*.�9��9���_i�7p�ˆ�t�������N�%̹Sp6Z@�X[1Oj���G���2/ח����f�����'���ѫs�������=�cP������b��%Q�HO3��J��0�\䫋���֦��\/�nBԞb�3_:iMq�@z�^��u?�k^�!�����v�K��2<]B��@m�ą��^u\�Ϡ�gaRD�ӕ�){M��#t��1���s	��C��T�-�V�
�-7�)���W�Vno]n����r.�S��CK)�ұ���Ve�jYIG]��=hK�̼�N�㠧�n�J�K��ܩgX�L��*f�7��G)̵N����d���ϐ���w�Om9o3�i���@߄�i�������7c�_XHW��@u�
=뱵��^9g�e!��.)�>�>ѻA3��,F5W=�c���uSd 7zB�p����o�T�h������R��L闞�.�{�ϼ���7��T���b�i���Y=���b�؆.����}κ���,��D�r��0�������޸~�d�l�jYcp+UG�W��J�Y�['Z�%XS�j���˵u�M���Y�ۑ�2�Иl�ǟv�(�3���+Ǜ��ܳ�b�>z�<(�����<� ���<>����w��s	�)��:i��t����W�q��F���RɐV�L�5	]���L��*s�-�Ӡ�i[W��zv�՛Bs����.���NPj���(3I�Ĭ��~fcON��&�-@1��I��2�r�w]��t�B�W]��V�JǺA>�:���2�֢KBb%��W�/U�W'���9�Se�И�.��
v���a����n��((���0��y�z ȭKdt���)�SA�D�Չ��vB���ՓE�3��;M��^�.UJ�{@BU�O3���䲍����;H<A���i+c��gh59�[�LD��"�gr4���������]�hS;�N��Oer�<'<'��x1&Bm^�F�����6��"*��&Rw��"g��9���l�M��2#�6�N�˜���%^��sNfI��o�;���=�����L�w׊�4���q��[ޤz�ћ�	'��Cu�d3�7
St���O8�fmOT�F�@&�Ϟ���/hx�\��ld�sT3���� �^`[�%���{j4%玲���|�ѫT��JB�;��۞ā�:��S����V��q4#/d���F0U\��S��<^ߝ@p���ЫL�`�s�E�V(ʉ�(�.�Sh�oGN�Ny����]}3�>��ԉ��9�!	�������z��[%�f�<��w.��<���υ�`!����9U>�_�w�}�T��z�����EE�q
�¹��W�BqT�o����l�T��ϲe���"�\�\W���L�׷&m �8���g(C#$1Di�q�*q3pjWQ���t�l`w��(t���}�J�m۱H��>a��>�쾈a�����Wm}C���T��N�7jC�vC�X}�҆���V�I�XM䊻�]s��YW0�ML#�#jꑥ������ז$�^Y���!ݦ�<�R�2�c���U-NJ��޲T��t:gn�*�kv9f��ȶ&d'��MW0SR�#� �	{�C�/�����S�]�E0%`�͡菣��y^>QwHϡ��s���W\>��JV�r�P��N�����2頜䭓�I��э�SSTb�8��}p��~.����s+�}�؞ϕ���X[Q�I�Y&V���0h�]�/_?VVQ0�Xo��H6�Ȭ���#�rx&&cLcx'rZ*��M�k$�x���k����H�9��sL�#؟ˍ�;I�b7�3�C~�f�ww.n��C�}W�/����E٫F_�y�L4.�7=Bj�f�p�sڅ9l�z
8�N��"�$j�0 �<V%�����qځ.]	���ʃ27��!@J�Ҫ3)�j^2�K�s�V��-�-J���˯�A&�~�Nd��o왤�ľ����嵿gMl&r�o/�鋨uZ\�^����d)�s��:ڼ����ü|�h�pA�~W��@��Y���Õkf���ŷ�y@�:B�l48����ܸY<�7�]̻Uc��Os'>!�V��0g���Q7n死��j*թ.U|�+-���@#x�c4�ϱUC��N���ȣ�׼+Bk;�|�r���WP�nhN��.��J����s3$�Mh��z�c�d�`�^��`í�B�oj��a����w���u�n�ѝa�;�N��w�\��ݡ�_�mԥ���S]%z�9���9����qLA�[&�Ӳ�o��ѕ*�J}ڙ�$S�pwﾏ���wYP���P$�6��]V9G��->&����~��}+®!�r���P]$�����+�N��~4����ϸ�`�	B���q;0�d��ɛ�{�M˭G{F j��Q�{�/>�7*�;�9��{�~lv�m5�����;SfHt2xԪ�tKfvK8
]z*���]���f��Øx��G���V�7��.�n4��EĜ$o��\��w+r�ܜπ��ʑ��lmD),�̅�;|7��^�F���:T�E���`PB�@lU����oJҶK�+of\K녟Ge��X��a��_%��.������E��f�*i�ݭ�`��=�����m**WG�'�ZL���7�>��|Ƽw�\@l��+�$8���.�'<|/���ӷ&�(|�Z�W:&��N�r�!�G2gy�cS�Pyդ��k>�3�[ӳ�c��֓��YT�v:�Jǻ�,V򉆁kI-���f��^���[{��fYͫi��f�t��޾>��M!g����XOWP�Ar6�$r^WRsSSbY�M������%���Ϋ�=�.�v/3]�-m���Γ�I䙕#�U���;3B��w ��$���H��N{4X��P��ހ��u-���60�Lk�yC]�V9�����͌]��ruD�f�X�X�Δ��| �V:��{����_�k>Spʛ�J��)�2Ļs3�P� _s|�z���;ı �3b34��[D��.d�9w�]��-���L���͚�x��(dBn�Kߥ�d�D �*;Bx����3��-�u���7tt}q��ގ�Õ��Iݑ!��з���N��^��\�����T��r�����nGm�#��w���뀌�z����s�U���YV��d�H��F�-��RDs����nn��1�6F}�	
�^c@�V��]�&:���Or�kL`���i��B��4s�zbo��݁���(;^\��B��Xe竍�ߧ�_s�K�[P���Y{S��������7�(G}a �r*����d�[30Q���Jk4�^G88�,bʈhd�+ a�G�nGz��N��}CL�y7+�.s(�j:8QI��oJ��0� ��˵u��sB-s��K� �2�щ�ao�}�3!������:Uŀ�)�E����&�L�heV�r۹��;�Fhc����W���PjON&��IfcZ�i-uړ�����L��-m��p�\��c�`4�k�u�o������N���:A���׹�i)�Pd��K�J�˝l- �H��f愉̧����۷i+�����+��k:��8�˼Ǜ)T�h*7�\��zo��L���ӭ`�o�:c��&Q[:j&��]2%n2C�=VБ�{��(3��G-�s+6S;5RpUdp��j��*g����N
�4��#�2��d`�%�Uh�7b�V�J냺*"n�C7��f�=ˉ\+�p����Kk�h��PDF�����5��������J��[��J��ffog���t�-��U�gf�eT�|X2�����¢�tE�w�n����Ԡ��q,P�L����b�am�ݠ�옳���"	)�`9V�6�3i�{��%� EYÔ�ik��X�T���h:M��ͤ��IqR����x����`�yS[Ţ�s�Wģ���֦�!��U-�^R��NYV��۷#�Hp���Y�bj�����SH��&w�H��驙����pc	�+6�������Hܙs%��4�#�7pK}y�|�0��x�CX��s->�L�ԥ�)�:�_r����q�բc~��)2�{޷Ϣ΍p+0w#ʬ�Ҩ���z��=U�O�-�H��K�Ɠ1�mK��&��uD/�<)��ܗY�S��m��w()E�(�L���Yu�Lj���r�E}�P��ntA�f��B�5bŭe,���N^�06�F�eӥj:-Ȏ�#����ޕ��5n^5hp5��Z����G�u5m�9�{���N�Li�nm���:mlqWV��W�r���⬤#���o5F� �u����l��oPػ4c'�oA2��-��E;Hڱ�=�(�3m;�{b�>=`�]aK���n����kSE8�P߳�U���bJ��K V���ţ�h��/8G��7��	�eJٶ���S4V#���t�C�͎�.��	l�5�3|b�@��"͓y h,j0�F�ܲ��W��Mu��:�����h�P�6��|F� ���/�R� �ݲ���I���jv�&�.�Ң U�N�Ew^���J��o�6�[|vLu���}C+IQv�k%�_i�V�&�ꔾ��
k�w���[{��r&Rզ_	:�؜��իỴcr��f�E�0��E�`��@xѸ�޷/9.�Z����ۗ������$����R���/f_WQ�z��׆��j�Т�3lRyG9sZB�2���m���3F�u_P�ou^Q�XrA"�c�+��xMFVD���-���� �9|�ٳ��1Ԙ�^̃��w!���M<�ET��\Һ�h���',w҂4��(Y쫩ڷő�{B>����Mh�n�z�k�u�[t���C	�g\}y�X�{�E�n�V>���8���l���7m�.�n������Jdm��ba<����V,�\;[;U�1J���� ���ٷ&��sgm�tmh)���r��/7*�=��r+a""(�'s$%s��W��9r�Z�4�*#&[�Pй�䉥fTh��d�if��<!�R$�+�u�C�!z�C��\��Βp��� ��NG�I�0�喋�t�ݒ�^heE.��눕�Q��<��QQW"�!��B-���*�H�Sb�2�U.�(����+L�I��'%=�w@�*BIR��=�wS�+n�v�T��3ȣ��֌�E�YDP��$�L�n��{��1�����9�<�G=<�wEԳ4E�"]��I���U��'5��qĲr�O�=��<���.z�t�N��Q��,��6"�mX���5t�nI�ЉS�u���+-ګ��n��)B���8�����\�d�����r�I�bWY�9R&���2V��e\(5-Qv����!����[�+������\
=��8>�SP�|�E�CvV� ������y�7�=�0[꺜��GV���\� E�湓R���興�Z�֧��NL���3�B;�B(�gW$��Rɒ�zd�̆ռ����[��uʍ������t���әr�h��.:W�:t�r���R�U�D�af�1��_*:��s���K�<�('pd�Yl�N�x�k��ۇv��s)�F�KBA����;�J��=�˸�mHhW0��Lq���S���[0����F|�Ιb���R�C��:�1�$�Ӽ@2'PS�dt�I��xȎ�(㰘�0�@u��X�`{��J:��fv_g��/�cI�R�ll���MZgq��x��/!ћ�	'��t�Kwu��go����rwwXP���Z������Pt4{UA[��/p�����=���4.g7[;��\���2���s4/�g��2y-A�9�*'��Vܲ;rB�jjw^��*^Xϊ�yy=�zM�n�jY{2��9-Vp�V'�Iک�2<�7B�Ø�V����Oo��c���e"�Fd�V=����������k�E��(^��P�����r���LE��K�QU`"v�r�[6!(#�l	�4��b�q��CAl��/60��}Lx�h�]�^�7%L�Gط��Ј��٧��N�L�{�Vj:z��+T�5-�H�C������^X���)��n�w����sVP�/��\�U���Q������*Ξ��o%u�<t�ڮ�߇TEFr������;"Y�ʘX\2�wz����)�ӕv
7�S7�n�_i>Fŗ�{U���t��Qa�wI��=3u�#�/Y�ۉv��+F�\���N��l��]�����jWC)�i��U���	�HZ����_Y|��j�b�zh�w�e��XD\-��ʆ��_��QZ�O�7��ć�g�A�ث�l���Ҙ�W���C���d�O��&�l.��'�_Q���j*f�B1���
uޅ�o2)���P[����'�ˏu�\{���uP�@�S2���]f.G5�k����ܵ��9!�^C�u��g5K�BR㘎��h(LƸ��N�C�B�aΔ#M����ǥ���J��&@�ұ!��s�&���q��;I�b6 ��f.��y<Y�{Z�H��UT`k�v�M���L�c9��h�ۡ�<���:c(k��SENK�4�Mr���'�1_�u��9�����-+J���+T�����3�ȑ��g�q�|�y_}�(�����k8H��轔���\�sJ�h���gS�R���f������/P�1��ަ^�V���}{������[r��8L�l�^�w6A;��,gY��d��vb�1K%p�o!H���۶oM/�$�e��U_}U���~[�]���u��J�b%ә/bo�NB"Ʀ����ޡR��OMc�3��:�M��M��d�)��Oqζ�,F�K:�x�]�/�f��F�%�
��b+lMU������q�-�w]��c�r�3늻]f�a���zA��x��^Nݽ�8�:79�Lz��a#/z�S�wh�#��;֍C� �S��B�C�}8ֽ���"w�N'*}��}�y��@a��j
��BՎ�[?\�ȃ֦o�ֶ�;���$Z�s�J� �;c3/��k���r#�#����<�م��P�� ��5`�}<q�x*z�����c�_]�f��[XeC�����D�����d^\k%����Xry� �Y����E�Y�p�(�[��s踓��@���ꜩ�n�*���*3{o���T>RXZ�����/u�6!C��[Xu�?X W���~I�qo˟T��I_D�&`���n����w!r�ˍ�\rX��.����4|god6�݊��Q��͠x�{.�+V�������q��T�׃�8S�{D�x����u���T�6WG�u�c�[�֝i#��_#�d}�G{ �*�Tj���M��Y��2�Ո ��zs���R����[_�8�Q��{�t��{E������m�d�j��XA�#$!\,�\L���7�[Qa�Vr���0gd�v��ؘ���Rē�/{�.J���Tt�C�Z	;����A�F�L�9�N�P�N��ӂT�f\�f3~������wNb[��\��Z�K��4�o��6*���7���E�sRy�oWZ�3ݻ`�4|��M!`�Ҡ��L�<y1,Aߤ|���%,b�kWmZ�Uӎ�j�9Ez�|�5�C��ui]�=\I�`�d��*ll������Z/˙�׾��v||�F��a���iS����*n1Q`P�M��p��V�<' Ң���=t�j�w������
t4A���ξ��<��i�F�Ww��^��`�q���+�'}��f2�����Ш}ZhB*�X�k�l=��x�zV& �+՟5�J!�ޏ��N�����W/M�=����a��}��^a�֬(�|昊���`��4�X̙���\�5������sG1xg�/�dՍ��aA��s�r�_f[��+&�&�{]+��a�z�����}LR�M�<�%i�:�j�X�[�⣤�=�Z��l
`�p�2�n���׊�*�K�AJ�O@�S�}1�Gv�8L�J�N��V�B|���ȝǚ^Ҏ��3h��(f��  ��U����[~
h�;f���}��;*��mqj��g��g��~��3�H��]lW=��i*���S�Y��,	��J��E�y�|��1��ҾP�Ld�������y|)�;��Vx[�����g_eۺ�8�hE�w��܌�9���`��UJ]�b0���U�?c�E!��ȃ���|+����n��3��3Q���]Q���i����n=ų!K8t�^oh<�S|��4�j��
Y ��CI���/a�;�E�e�!ݘ�L3Ӳύ��懣:O�:U�.F�KP��H`���z��춈N�)���u���ގ�_�u3qF"��3*鑩�O�� �t�3��S�$��O��r�Ǎ���+�;��ڥ!�!wP��.��
v��2a��=�����u��,_{o�\��qⰕ[�o�P���������z��j����(e�o�\>�f�X�}�4cР�^�K�Z�3ѓNfMC@�29���r8ɫL�!d�ᐋ�/!ћ��h����6;/jz/�uaR�7s:r����(���a�wgh@X5^���d� �ub��]�@���ۙ_/��fj�	��76���{/	n�.�x=����a�|����Ǭ:�[>�v���H,�k*�-�
_v�᪶/fV].yjr.�ѐ���G�������t����1}�3�H���JZ54����ԅ�{Q��j�ިS�������M�%�T��iLi�ʪ:Y;3���2��1�S%yr9�-Wl0��y]�3t�G�Z�wݳ�B�+&��c�-��7����<^��u�뼩�U�4*�(1�;�#�n�>7W�ol��t��M-R�vt��Jcd�lf�[��X��'41����۝7�s$����U���^y�S7�RR8CpK/���}� ��r��,0:&�9&��f��7Y��=�T3��ڳ��Wx>�l�K����Iy�6:=��Y,�pr�Z�yqV��f�����g��rszPO|5�l�5A[�Ŗ+�{]�0V�Gc�8���&&,���^ޢH��,_�,�;�.�u֞ҫPǾ�j��$d����eٷC�41�8�^���y�Z����?��d�)n�W8�s��erw��(l���Z����S�l*��:��f�T��:�m6�{.�]b��r�)�����%oF�u,Gdk���#Y�=���W,���\���o½��l���OjkbZi`Xߵ�Z{�޷���>�����f޲S��Y�R�a�'��G,SN��:�޻*�#�Z5ʗw@	\���,�0eh-�M��O���n
�!b����ӮKI3+R��x[o`�읔\��.���;��IJn}_UWպ�>�=�qω93��L�rFX�i�ʳ���Ƞ�UON�c��;}�LM��}���C
���T���p'�
��7Pj1K�����gNh��܇��\�U����t��y���MYU.��P>��)5e76��1#bV���t8�+�����:ʑ�ѮK�^�w�Y=,�r�B�N�T	r�MR�e������oٔ���>�H�WsY:�����E�=�1M��r�s��&_PDi@vȩ\2ۊ�#y���G���GCYP�#{!L_'��~m^X��&T�ΆbV�ND�M`t\�օ�VN5k�!�U���h��D$;�:{E�.��a��vj6���=̔D�Oq]�ʜ[N��qG3��;��=p����+-��A�D6#�&4ڿ�*�z# �XF������"��r� ����w��M@au���f�yP�c�SV��4Cp����ka�ӿ]Ի{d�fܫ�k��������MPV���5¬]�*�!^��Ӊٔ_0<>�O%���^����q^6T{[^�y������3�ζ�L��;N4�w"R�&��mqc\���7��;�{�xY~T�;���W���.ʗ��o�wL<4Yx�����'|�[��>�>Ȣ�����wz������ ^l���j����U}_6�u�e�G|T�!�y���ƫ��B���q��\3���.q����|�����U�f�OG+��Ɔ��@�\�{n`�|����ÿgѝ�F�p���^���=~y��1�U��������HAr��@��ذ���܅�S�8�p�V̂o�I�h�Aq��!��� �S9��p��hC�b\��䱐X����^f�O|���sY�U���*�vVW-�Id���7�[Qp�9z:��h@l�0eR��U@���,;f����[b=<c�!������Au#1B<j��f7�(0�sp���{���eK��}�/:���d����\�C@���ߠ�$&'z��������v�c�k��SJ:N�b�C9=5�����M!g��� ��	���H.U6�}�����H�ޔ��^�s��Ѥ%�n�A�,�K>sl��섮M��<� �(p�*���+{e���-�9��ޛ�����Ş_*���8nZc �DaO���W8�`P)��>�|�ܯ�A�32^*�u�)�X�E���>��5���R{��4���d�.�������`zmuFU��}`��q&�FD5l��Ɇ�tU/�k[���F���B�����VsK�kQ%��q�s.��m[���\�K����ȺȽP�M��DDXkU������jW*ө�\)�����m��Է���������w��Q���{Dt�U]mђ�X�x]����Pxh��d7��B��@f���V8W��l�Լ�{�X]7���ec�شd���{�v��5��uno��2��9����^�P�H��:���8��ss��zF�����k�s�S�'\�2*wC�����3�l���:Z��cj/8�Xt�:s�ǧ�˺��=#	K�[�d2M�޹.����ɱ��H�Xp^O�Ύ��Uj����*�e pH5	�ǙcTCCS�Y 0�����C���ϝ��;6m�h��Q-��2�wxc���������Fg����NL����Y�nF2�Ь
�}{��^�[�ݝP5�~^�Z�T�A���a��*¸<oc�n��:*ayP�u��$�O�fm��t;s��p��{��$i�5rKiK$ޙ>2]����u-RV1�����Q\�gk���T�g�hF����.��?C4*I��jIs=n)��u��9cr6�ܙ�S�Yt���Ł��bwStt�+��֤1T Z������Ǣ�pq�ͭL�pV��p���I�`{;�,�	A��N�O�K��F�oP��8��S�2<����!V�|흭3�N�WJ���N-���� MO�b)����H���b�3jg"�wg���X0�}~T�7�?�#ˎ�+v��xu�z�"g���7vEz���l�X��� J#5T<�QC_Sk�t���z����tȝ������nꁳ����B�)^�T�A6�l����T�VsJC^�R��F��f�7=9�ג�o}���^����&z���|��R�F����B\�2hZgq����R=��wC���osKo:��fg2��ސ3��(d��J�4����P+��E�R����M�gcoz1s9P'ڳ>&��6�\�>�&Us�Ω����mZ��j��1P��-����Wu�CYNa�zs蝼�8Uۘ���.����w�1��*Y�o��w݋6A���N5r���#p�"��𺍘��Ԙ޳nTH���!;���5���s�C��O��]>��(Ʈ��}��p�pl��۾.�	��Y�{
������v�b����l�S�v����𭆬:��6n}Ip��K�iy��c�}%��H�$����j�;5�;啕il/1H��SL��=��^*7Dm+f]�L���Ӥ�NnVd��9����f���q�_.�R��̬k��8��@��#h��-8^!UV�N0����;f�����Ah�vfe6��7�om)e)r�z�ھ�c�k�Uռ�6Р��XtwI�F;�s�Ҿ�{&pu
�_;+��
�A,�����mp��)4Fd��[Qpx���v���v|cMt=��,^���M�z��>��kV̟e�������5w�l[y��)hs��r�L���U)'���H�!G�)@�asm�g%�G��/�e�R�P�N�k�W�GY���$�b_!Km�>������0ݦ'8]s�e#X�䝇ܗ�e�>��ʝ�>�w�	�V�=7����1>3�:��y�]�$ۧ3^LN�ɤֽ�	��W��
��o����X[��ud[6D�GV��Uv2 �R�ϰ�:��|,����λ�bㆅcC�߆:��q��j��#��MTڬ�h��\�U�3N=�<q��aлA�ԋq�V�"� �C��nZ����3���B��Ӷ�d��G�cu�b�|�R7�ka֮�S���w�G�	;E���6�S<��r6^	$.ʆ�o�\<:��!���v�F6�Qێ��M��`���܍Mgc�c��՝o5d�+�?G ��,t�B$+��r�r
�-���λwKj'��vo#������N�L<�O#�a���c"�L�î��z���g�����˩�8�囙����R:r����}P��Hu.F;������n�m��̥���1waZ7��J���������{��P-DB!�-��8�0��4w�X�MU��������{�Fzi�M�9+p����xr�����b�~��Msi��ҁ�����j9�X�64
��'B��p�ځ��@HL��Ha�q����f�B��l$K�Q}�p�2��E��WB����pZ���j��H�S�f��̾�y��p��]o+Wpݩrc�����`}|�#��-��VΈ^+�
��P� 3�����$�4���Πs@:�!ua�D.5��,�ZSm��B.Vc6Q�|�&9X���mc�-����4$�(�ըm!�u0İq����db�lr�m=�Z@���<�&yYx$�B��3��y�|�\6,'JPX��R�]�^��+M�W�R����U�/�&��8�j�X!��{4��N�ӊ]�Mw)Ċ�\��dE�]ͶkZ�C-()�ѷc)\�+�����:֧8�t]����,�h��)�t�"Y���p�la�Y5�*r�����P��h�/I�+V�{=d'���s��i��c���6���UԆ�Y�'���\���ǁ(/���`�ő�+�L���@s�n�0F|7�t4ӵH>'Wu=��o<Ͷj��oe�J�� 4̏y�|�=����2�dJ$`������1�&{E�s:T.�����W���	\���O=��8������r�*�	i9��-3�܇��*�^�������h`��ss5Ϋ�����fQVe��]P����sS٨�D����]k�����Uj�D�J��IWW5�np�w�����U��=/=�ZJ"��Iw]�<89�Yey��^���K���J�'3�=MݺT\�D�H�@��u��e�T4��Y$tR4�<�Q��Wsr�������UQ��Ҍ��9�{���3R,��ĭb�{���r����\�w2�*��3T�*��S�waI���z燐�\BU*�)P���՛F{��B�Q�Y¬�*A
��2�*�6&T�j�I��NG41HЪS4�S6���YF���Uh+K���K������.����KI!BSTXGH����]X��w`V`M����Y5f�������V#����`I6v�ɇE�4��QNʔO!����˫=�����α��K���j�������}:(��
G���؁dGv+�"�FH�s
a�a�H�
�|������G˴��9M��ħ�������Bt�:�̳�Sz�ۙk"�$d�|�N�7��ue��"p��ԍ43{�Ӊ�q�w0�o:y��9��N����P�=��Y�(H����4�gWu�;%敹�8���U�-̊c,>XJނı��N��طٟw������No;�[;�Nh�'��I̚�ZL�r8��i��>ձO����;��9w��$a�il��Λ>y��r��>F�O��针�Ў��.��J����S�q��;�'�� �bM�`�lj��%��^PX51m����%���U0��dJ�٣{n�d9qX5-�zx�ʭk�ޣV'���N9g�.�k��B�N�T	r�M@�.VX35<~��V�w���*��������Φg!<�`v�G���SۮK�O��j,�����
��c�A�k��r�L�r��*���P�7���{�o����@����a�����^�
�g{9%�)	:��vY
}�y�w¯s}���++M1ՏI��n��(�Vө\G_r{�\�:�<v��$���u����Es<�vՠ�i�ĩ���dv\��u��m%��wX��c��1,����O��u�X�z���&��ڟ� &j������W�g���Aa�vk`�����z��?N�0j.�]�؞��
P��-�[Gy<'uU^h�W��Q�
Ш��`��:Q�\��@#x�c"4�ϳ�UD5LaE�#�Y<�ZG�]A('�E���p�d����uF�y|-X�m�->&�)p���#�su�L`�.��S������ֻ�N������>�^���W��������*��Fct̙rg�UN��/�z|%y�x��f�`U��0 �_d�D�ǵ�Ka�R�6��R��+=Z�:��߆�A����[��m��ve�lV_���vqZ"��X��_{]�%d�}H��^<j���A���x���j��Xc�]���\r��CI�P(ٲ�j�Ү�_�0S�%���d����� �B�@r�F_v����_��Oi2��|���ݟ���3p�����UB'��ɓ����
H}�.�����Yy��U��;��޳��e��Ɓbtr��?m���d���MP��M�U���l��Q���Y@��΃�:�B,��ԧ��N���W0E*��Rzm���2;i�坘6E�Y��#��]l��>���vӮ;���ʒ��@ݣ�.���������4�$�����]
O�X�mXF�i����Ԡ��@�N��i�NgLx�Z�;I��%�S���=�Ay�@�#Q�� 6�׈U�\Z��X�w�λ�&������.9b6	�C_;gл��,6ZT��	���p 13[w�-Y/�S�V��T&D�ӥp6���n��he��t�}�A��? 0A� =��f��r^gOV_+Ɗ���Fitu|���p��8��M"2
}�6�*L}���c�SLm�g^W6𻺬d���q�ZJF�kf���1�:kl���O0u��h��ww"Ӣ�#�i�!n|��B�҉�{Ő~��b����Y��B��^A^�W�F��;�d�O�]��d��{W9.q�gcQw(Bf�~�������ќ8�ϽV��0��č������zu�ua����W�f_hg�6�Y�}���^ᖐt�}��rə�6l�T���V���x����]�qYQ�b����P�f����VT6:�WQj�`���ٰ"��\��|c�����C��Ϫ���<��CBt8��a�eQa���*�R�ɖA��!Xh�N�E��8퍫���O��շX�6��K�B*6)B�o�)V�K���)�]����{N4�9�Sr�V�{���ȏV��̭�f����a���G��7��рl�^�D�˨]���U��{�2��c0}^��V�?5���" @�k��o=7�T��X�F����M/�����]WT��te
y��uqGe�����a+csщ�v!�S'�/��Z�������d�3�;U�n�Z���1���{���o.���{�O��K6x�^״pS|���O$��K&��K����0֗W8�]��s�4dFi���d�ס�H��i�����f�ͨl�����X���o+|��wrٌ�w3q"W����ڙȠ�ԹC��뽲�{*�mW�z�SH�{hć���e_[�ӂ&gDTJ����g
D>�E�o낝�7��f<�X�?P~�'�?E��j��L7CP�^C ���������!0�xȎ������R�rZs�=�ͣ��-Eȣ�-�Իǫ�Ӛs2h��!L��M��*�57�I�M.����Y���W:Ū��)�3t"�On�9�D��X|�Zx��?e��i��V6c�{>�c+'_T��c��U�dq��3p�]Ѹk�s5��2�s���*�|N�j�W`T�.�3�Y��.��خY�y���/�+�;3['\�W�hW�[�p-��N�8"�b��[X��Y�e���8�
ڕ�7o�XY\��p�=K�X�S௙/r��寀��M�x�ڱS�kI��n��ъ���,ۂ�@��ﾯ���;�S1:������ѐ���;����Ӟ���]�c��������m!^Z�����۴����W�GO1�����2,F�l���F�s�MPz���]E`xx'�յ}�,�~�����N��]��Gm���x��R���]Ya��M���W]u�k��Q�{�z�C�3{E+S�F�:��9������5��2��PФݘX��,�ղ"��()��b��
�#ʀ!��AK7@��Ȕ��$s*�UVq�6��2g��J�V��ɦ�1�����P��d'M���̳"Ȏ�v��3?&$$fl���W�y�)Fo]�. ���!�ϟH+����LY�U�r���N�zU�I��l�k<K��;���j�Uv�)�+�X���ʴ��[v'�����\7��q�^+�s��=�s��mgYt����Ȱ©�=4%q2\�"� �v��E>v&�x�½q^��$�g�6�����}ɻ:H��h��M5-"��Ў��=H�	j����S�q��N��&�WKـeֽ�������P��o[T��p9�V��JB����4��ƚ���l�-P�.P�џ�B��a9���Uc�˫�7~kv�gI�'[��ERcM9^��]�L�ʢ��{'"܊���ɣ+� 7�ᧇ�ﾏ���ֹ�3��n���c	���x�������%���
��f%olܛUv� ��d�:D��KZ�pk�eG=�,�s���!m'pz�K�BkVvj�*x�D(HΩ~��@oBy���Jò�6�Za�3���#�f2u�w���w���}A���ֽ鼿9�����z���U-����L�u�+��'���ڼ���L�L9��+o'��`��xu\�fO3�U(=��L�F���w�:�!��������ad��]̻T�.�<!Wռ�]YB���.��9��+���P9�)���Z5��w����d�����
�@�/.�TH�|��gu����^�:�lh,p�R�S���m�C)3��'{��k�F)���2�O�:��C�ߝ� u;�'~7�E��n�)����T)��d)��:5�E(��DY8�x1;Hpxom�Y�&�����c���x;��V��ۮ�`@4;Uռ��rp�V$u���{��Q<+]�Y<��]l|��$B9*����ϝٗ<.�)��6>��9��[nh��I��Jg��]d� ��`��*O�Tl�$����T����k�5D�*��\������"��yoR@�8��&���J��|�R���;=�cR溤@$3�Y�Wq �|;o��r)H���+S�����,Z�',<r�n����_}�}�}xuOCǓ�5NM�r�\�%>U
]EeH�U�0B�fB߈v�o���/s�y���L�4����V�{]�o&���t�X��!���xL�Gl��T����G.55rX��&�I[���«�]�����2�\(Ӕ-�l%M;YZ�hD�d�;;�n1Kj,<��G�/>e��z��ח�S�
vr���ym����bKѱ�!;^��u���M�Ď���*���i���8K"^s�O�n1��tY��-VVN�
g{.�ڭ�Z�1��O��P>�,s����\g��Yٗ��M�ob�v��A�R:���n���XJ���葊�H�Y�z�	M�;�W�2�[�u��V|sz��8�f:b�v��uM#��;<��ͧ��T��v[����8֞��rFO���E��yf:����[��j���Ƃ{�jA�KZ�mt`���es�J�u]�n���Y᪄�t.��]�kt�צ���ZIwс�W[I7 ��g\�ڥ�Ԙ�׼���u�3�'G�+��v/#Vj=���e��y�*�����邞��|;i凧]B�^�P,=�fO�Ӎ��4��f��ι�1M��;k��f�/2tt��S��'�G�}�}���W��g"��<�W�m�(>+���q�mU�ϵN��}�[��=ȁR�y4�/}��y�j>����xҪ|���k>j����1��0Nl�Sӥc,��]:��i�VV�D�rruEDaFnrS��Og�"r�lc��~�'YM��n���k�2�K�J͡��9,sӜhnl��R�'��U����%���'���C0���	���{6����2��W]�R�mr5��X�ga�M�}O��{r��2rBa=��T��4���.zZ�z���j�{��{&z�޸����aW:���'K��q5K��f_.N���D�ᤗA��o��	=�/Z;�8޼fv�%sr��og��6闛�O������I����	-S��d_��rV3�	�M�s�Z�Ѿ��Ҏ�Ӆ�k��XC���_%_J�.����8�3�4�^sq20��*74	���N��eX}6$�ee�se6��O>YF�;5ot�[�����bp�kp �4�F���2-�yŊ;��:���Z���/�IףJ�B��պ�Q�Ь{;(G2�+�	�Ne>��=X9ڝi��\�p�`�i<�I����ﾫ�o��k�Fi�a{��;��W�f��=�S{Ӧ6R�}��ss����]��{wx���=eؗ,γ�
ޣ�!<uq��U[&;k��o����vZ���ٖ������9Ԍ�90��/�ôG�����\O���g�?=��$�k�W	�mm�<\�����!�iiƢ���,��3�__m�©�\��ϟ`�On�3�:g7Jm9�± Z���q��wX�z)l���k����S�D��>�h���~o�;���|0�s6ʉ������>���+�,���8B�Ms�eNg��^�ֱs����w��m�;���#�ӭ���Ta��:�7&�=�����-�;O�\o�2�[[��C�}a�;�#���+�%�n�6���v�Cs���&�ǳ��ŢM���<ͭܶik@z���2�DY����v�߳{sк|��&Ҝ��"�}�A���*�@���L��:���^Tg-�?]�X��,=|!J�T,��n���ۗC:�q��@�ya��G���1v'.ѿ5������hn������菾�Y\����ޑ���5G]�h��A����F�]i��/����Q�7�����9g9�`��W'���w/�e�q�	I�pνp��\ ��uN�o��η7��Y�|�=;e8o��mb��٩l�������D�弋�v�U�Zc5����:B��P~&���K����݄8�j(7o&�v�q���w��+��y�K�ke���	��t�B����Z ���+�BP]�-�p�W���Z�l��x�dKȯ� ���@�ҍ��6����_l�gry|��msA�j�$��D��\'Ba�����9���s�Z��Wi�G�uf�����j��k�W�n9�6�UT/5ak�b���`�NM}8��w�Sݿ���s�9��cw�)+P��\�]#�3��]����8�w��2��ڴ��M]b��;��=A���2�c(�^��^��N��Wf�9������KR�)��.�|�P`�BY��r�`��#�N�����3�i�*}Һ�r�,��9����QC�{n��̦�a�j�ҮU�p�mR��X�nf�|/l#\ea���M�Fj������L=�5�!��{�Ū�D<�N溂u�B X�y;���Q����We�_`��a��k�n���)��dS��D�t�Bn�M��o$�W�����Q���vsc����p`��}w�26f���;6�	2is��*u)�W7.vI;Fּ��y��H�G��	4Kp�!��=����,�![8@�D9����	�^]�NnVV�Pm�6�CW���+����F��T�4��X�o��S-Np=~B��Z�����V�{0ɂl��Z�����O/-�;,�����Q�m�r�#�󔲎h�d�v$#.eM:���0%���3-�Op�W����#:V���
�=Va2˶��ij����V�N���Ow �ݒ�{t�#�]Bf���z��N�Z��ۤ�a�������*�#��(��f	iXM��2�3i�sxGG�#K�353|��o���S"���*r��A�pC�;2����!�G�_X��OR�t�Î��*o�[��4�yK<&*�3����d�ML�ˠ�y8�f�c�Ѯ|�+�uϬW�oqpF<���p�Vs�tn���ĦSi�̫hˡFnsWϚ�+�T}V��]�P�� 35�A_M��P�[�mU���9��ŗ%�7ja�W�*�@.�]K�@uĐ����
�㮨���)�rXs6�ǖr�9ĥT�'�33t��)����8�9i��B���o	��m%a�:e�1�f��h��
f�o���U��hu�>���x!�X�ww�&L璠};��o��xz�&��hNVG:2 w�D�\w�ʃw����������5]�Š����U�D�O�:�a���;�d���wv�]ʸ��/�Xu�m��E���ӷ`�-j��]%Ջu�[��ORhp�]�j��j�ۭ]��.՗k)^����W����8����w�aGul��n>$Y�
�YucqV�o�Q�@�q@��䆦G�w=)3x�`976Jr���:������yיNK���ټ1��\��Ʒ�]G��Z�2ޛ�W_㿣�4r�â��2�>�(�f<T����:͢�`-.�<� S��T�����J�#�/(�(���ʙ�C`}�ȹ5YA�ׄT�,���~6kL�@Q$\�]�p�͆��fc�s\NWdJ&�T���6To�{U_vn.9�q)pӳ�8ޟ�������a���#�\�r�L�ҋ��5�/�1�m��6-'.,B���̧1�:��I�v�+]ǃ�>��cՅ�e{q��f˦�s]wg*l��T�i�r��u��+���/$7�i��5�41\`�[Ë�2.�nc���W���W;Y�Ͽ�y�{����jU]hF�B�G+�΢d�!GU)*������4�e�u9Z�\���Z���)�"�&TY�E\I�*�R�5$0Ⱥ	[PV�KJ�L���Hy�Ri�E*Ab�:uX���I�9�&Y�XdV(�V���UU2��)D�0Y��D%$���Q2R̪)4R����f5B��\̌B�:�EՂsCZJ��"Y,�8���O0ֹU�U*T�Vi�2BE3e�JXiQE*TtY��jdb�4"�WN�I��VQB��SP�f],+��D�t�Q.�Rʪ)5�Tj�B�wK�U\���u2
%6��"+	����H���2�(��Z��h�I����V�,���9)���QT���!YQ�ERYG���^�����v�(i,�v�(VpSR�Fl���Q:���7/�Й���q4r�1��Ds�9˷���˓յO�"">�Cp�.�Q�3@;�'��)�<A�}io�;�iv�Y��ys�ȼܼ�I5Fw�u�b�q����:�N�v���ۈ*weY��]*v���x/��֥V�f_:u�4a����2�zϷ�}�'��Qd+z=��fM/�MGպ揫�-���也�a����-6j0�]�8��w]��y�Ĳ���T�1���s�s���T�䰞<t�b��Dk��m���uc�n��7�����u��q7&���
K+�$���v�0�^�X]�\b��}�P�ז7F���퐘Gw�bm�"�����{��77[��|��&w
֎����a.��U�h@j��QuyK�7���^Y*L�X��k�8K%�>������O)��O�N �8���;�ó]E�3��u��aV���Rٗ�/���*��"�%��ɕ0��+9N+_e��Z���n�	ùSX���T/�.[��r����P/��v���M�g&���`���ZqRuč�p	]R��c���b��6���t�M�-�3X�������+u�p/6!$�}L�n-:>C�>�ɷꕿ  ����x�ꭡ�+���H�\G���֑up�2�,UQ�[����Kr��P���5��Sꃷ0�znw�9�1<tr�;22���UtP5�3T0�ݬ�Ir-��t$�S���%⿨���k�s�Ųw��k���1�9C�É;9����О��<q���7;��sB1����~��~VT�F����<�����[��}�p�j��b���7��%�_s���\�����/!U>a>e|��gg&�؍Ud�$�봵P/���9WӁ
�zܵՆt��c�]�2�����Q&.�3�����V�������nV�Y�>�wW�Z��'�+�܅�7
�
�yroި������{\��X���%c��=5��a�7�5��5njֿ�s�P�M��;O��}P{�3Ҿ��=��]�w�۫�;�OYq(R��#�,;�}��f�G��0M����϶�.w�f��Ѓ�[)�b��9�hժφ{�+`�\f�ўG�$I�Z��wF@
����Vu��d�T� Jt�|V���1��
�j̕ɊV�Y̻�ĳ`[��U��}_b��h�S��|�\wW�&�>�nF�]i���>��\ɘ��tﭮ�Kt��r�k+����I���q�x��¤���bu����=m�[ƮV�������Z�C��A��9��g�>�ɼ.�˔�ӷ���2*m�hS'>?%Q.e.����C��;��幩�Hk�%�]���'�3-c���7��v�B���W��f��h�i	���^�NmՓ��Y�Y%�l�_K�.�¤dk8���!<���<�=�4��y�hwS���\�ٺ���m��+"�ؚ=n�?&�->�8�@n��@�q��VG�˯��Ȅ�խp��p:��~�u�0��{�����3��M���{�����w���ǟL�.p辱�-.�ׯj��i�&J��*9�.����.߰�m^r�j>���ǳ<��Ķ��a�]
j^!}Õ�F]b�8�����lRʱt��Q,���T�hGc��V%h4���ÐY.���]�XC�>�|�ǳ�u|�uݙː]w��>�I�kFԜ3OӘ�`E�vC�ҹ�R�c�b�3�-ţ�׶*��9�OO���#�k�m+h��}�m�ͣ�2ϧv�<�����ۉ��9:��d��i�v�K���Zc[��rR�W&{�ί�.s6Ȟ!�Q��;���i/��n9ꖕ9�n����[�I�g�>Xj3�mũf��㹴�N`��O.�wszz��P4ͨk"y��������e���`"'�Rl�F�o��d꬙�8Ԇo��_]�f͜�A�ȍp��]&�j�*��є�a�Ճ�]���p�e�%�q�I-�����\��p�DP��:��v����c}�^i�C��;#c�S���&�.�9
٭��ݱ}o�+����k�'����z���t�B����Ȁ�OJk�M��jc���Y9��'�Ȁ��=y�u���}C���\���:�,g��N���w5�/,�F�-h7o��{��v��[.�X�-Ljk=��Q�e*&����XkNνDκ�3l�G�����9�v�lӖ�-��}�2*AD"ɒ�7G%�N[8>�E�P�y���vuI|测��[���kz؉�<�{tLc>#��V�Ӹ���qY�֎�mp]���kz��}���0M��ﾈ���R�m�[�蕕5*�gk�N���ui'/"[�y��7�ҩ��sg����~��쪰��ß۹�_V}���=m���¨��W|FNo^��W8Y�f:ܜ���M4k��Ѷv�[Ky�'9�Z{���!G��3/$øJD�Gz$e���U�=���{w�r�Ή���Sy�ߪ����ޘ#X��:�1o�u>�0#����}im�����>Hn,s�+~���^N�ߠ�"��_;�q;�ϻ:��ҧ3vzi8ULx<����.�';R��Շ�^zϧ\W�Qc!Yns�m�B�ݟ,��s�ȍ�er=�+YYT-���pT�W�$b'���%��e�h�J\��U���&��>3�`,��#!o�.�P�ʉ_]:�P%J�C[[L�0Nݽ�ԻGU@:��r���1Rr
���V=��v��W��K8���6�f���#-<TL��T�F�]Zz%����x~�2�MJ�URk��;g{l�m'��9d�r�JT���l,���B���{��}�Y�К���E�k�����{S��&"���wR|+pEu��aM���Ѫ�]�:4��w�V�l���}��d]Z\�^=���}�˳�P�k��]�-+�nI����D�������z�!-��N��F��f��;�V�y�i��n%q7(�MݨQ�D�tNsKXO;�È�noCOu7�9�m(w�Sݗ�ΰ�r;��ݧy+%V�w�jT�uu"����q���Y-�y/��y���)�?�gOj�����ď(�Ȁ�՛G� ��=iAUξ�.�����JV���sn$���~T����S�zm\e�Ց�+~��2KBީ�I�n� �&�!΄������/��a\P�v	N]�n��Mi������ϒvr8uqT�On����s*�G�Z��)b�VFZ��-H#��ν����L�.pZ�ls��Hc�:>�X]BG����3��;��c�[;��V�/S�6-cW�L�醞t5�T�f)ݽ�JDm��L�'�Q���Q_��2�'�SL7OsE����nj�J��=�G�usH��Ki�ҹX�r��b��9kɻ�E���;�zD�,���i� ��ΰr�SW��^.�Vv�K�k�8����W��0���B�8}DG�m�%<�X�Sd������Ê�z��|�>�w����n�=�߮O5��O|�Hd���m�����^J��{��=]�49�wA�I̜��Ҏ�["����l<L�y�d�MUS!��G|�;���R��U]媺{�����wY����c��l��k��'�S=A@B�9/_l^�[�Vx���	��K`j�V�&�9�[��\Bi�Dj�nJue��3�M��i�Ud�`�\�IV�}W'��\�������2��s�Y�g��%[�k���4nz3�a���w�5���l�V��k��񏪕vjg����</x���� l7 �A7��b{�g�oN��N� *��$0��[��N4�^��ob�����'�|5f��6��ܖOP	��7zʵ�����.��i���\�K�dk9%oQ��H��o<��~0��l�vuُ$�6�;����� rV�٢!u�ν���Z@�Wvr"��DJh��<;k��I�.�#�-vۭz��ս
d-#!���'������>ݱa)0ޕm��Mw�}��A���ïT��1�d�*"���}����O|���;Lx�ב\��a�ui'"�m�<�Y�;EO'�n���e��z_U_v5�7��W8��}Y���^,����
�P5�m��7�������.{J��9�b�\��4��w��ڷ�U2�î�V������r�vh.7���a�2ARʳ:����n&�����:����8�`�9ӓ]�d�y��T���з���{�ߪz��@yձY[MIFf���|6�2�Y�����-���#��p�V<p\���<g�>�3��wZ�Km��4��P�5�1:��E��i�+=�g`�R̝_fG]�u>S��=�N�눐���J���QΑ������v_MrQ�;ݙsr�-Xq��.�8�2�R�����]�f͜a������|6Y6�6�7���Z���U�7.��2��G]$�e�p��XI�U.���yya	��\�v2��lP��sfQ����D�#"�ۚ鹤u�K�.�����ǚJ���,�2�U���pk"�Q_d{O�������I�F�Հ�[&:Vb�:����h=l��K� �o�U�qv3+�+ ��'���k�2����Pܣ�c�G��Y/RE��7P���go�%q7&���P%'=)"������{�wV�Aj��ʞ�\J�{a8޼nv����?_#��L*�םؐ��Sk��8��L�����Ľ����⫈����`�˭^��cN˶�E^��1���+���|g�
-dD�e���J�q�*CyF�;=�U�ᛅ�D��e�ʀyVR;G�|�wٺ�����k�i��M`���/���u��y�v�����ÚEl���G�[j�Fi7���x����N0���y����N.��7Owis��r��9Kb�m�f��`u���̜�yç�*� ��V/~�&�q�wU�c���u�[u���R(�wN?�j���UO�
pZ�Mi�<A�}ih����Jf�1�3�[۹��	Nv��\�*����j���e�h[�»2M���m�R�t�4D�V�ע����`�B�F����k
j�u��R����γ.�l��(֛����������n_��=�,v��*쐞�S�ɽf����"����Y�NI�:c�%uq�Y�^8���4ۢ��8m03�)[Q�����V5�_)�u����XS8yVΩ��D��++n&�3�N������+=��.�"�s��|�X1u��Z�o����?��wA�\=���컩j+������<�I&��5�q5x�w�n�u
��u}j\�al��EY��s[�ͭ�sU�C[��3����_�9�S=A@�e_]$���T޶6��d�C�:���+۫�&�9�]�����-+�nM������2��l���)m��hA��.�g�v�\��Z������ä��!�찅�)��Ӛ/t�:�qW��"aj鸎	-�8��N|K"%�>�O�q��(Z/�ui�9����uVPٛg�k�����_l!�q��idKf^�d\�,�or�-�k�Fi�����-�Stp�󦶞���}C����X1y��n&��y�t�.^D��%dT)iLk9 ��v�'������7d<=+o��SN��,o	J�:��YZnR蝀��qN�nu�r����՘+�q �E|����'h]�K�G�ẀR�k��L�Щ��+1�S(�I׌
���Ws2�}|��c�/8�2��\^��Ȟ�%�7�ɪ��x�s�H��Q���s:��A��)�YٌA�O�|_5s8��(���+Q����/v�rn��dV���ڽ�7�F�lLGV��;]9���A����༩JK­0:��E���,�/����O�fU3q���6���Ҵ��=4#&`�c��uǱ'|jMC'R�Mvג�`(��cx+��Ծ�t�������g#8�Ġ��)���d�[����2�����}��}u;/��Qb�!HY����ܳ�:�Ko�q��ٯ�YJ���\/�EV��JMͮ�'��+kwn\�ݤr�!X��/f3 ��Ț[Ш㫪b�f
���忦�A-��ݭ:mZ;�+���� oU�e�D�jʉJwl��^oZ�ao���Qu��v;�pǦ�-3�u	n��j��K�����'J���C'�iUIZ2�����@X����ҥk+F�*]��m�;*E�`��֛LР
��'�SQ�ᩗn��-u�.wo�2s��Y��eR��K���{�f*�J��>�:��nM0�
�P�m���6KFuwcʴi��3�4�¾C��6��w)5]�r�f�hl�/"6�^eA��z�%�(.��X�x�Cf���i���k3�X������f'�βԺ�S�6�n�X��4�)��F%	q�U����,]���OTޗ�
3榪
^��&�� (�Y�� ��y�{]�kgd|F�_#l%�I�&Tʘ�c���Ê�*u�JV�m���h���s{����$k�@�l!�G��5����D�C�y�j宸:O:Q=9�m	ԃ���� ��}��F]��j͵�HY?��5(�'r��U5��G͘��v�íV�4���4�������z���ॅ��f�^gR!G�'�0r',<�}�1�p2�e�#�Dꛚ�E��4���[٩gojXG��Pދ n͕��1�r�٨|/6&;�>Ѫ�uBKB��e�"E�'�_V��|����<��(H25F!�\\tY����ݫ�ѫ���ʝ�˲�C�;j遴�$�f$k���ُ�65�L�eAW2�:SXo�RŝtU���0�����@v�v��i!��a�]zFP:��<qb?���{ڮ��T�+pԾ�r�I�6um��!��fԳ`�k�g7�#Z�2ĝ����WrPG��IZm�DR�f�Y%L|���+�[X8�Ȩ>W�gJ��*�sx�o� �.`�e�Z���]��l8�@[���鰛���\����z�X&u2�y�R����_"����v���|XNõ��R��ݔ�v��AN�.|��s��UypK/�d/f��=b���n�Jz�A���*H]�g,
U�m&U����,���g+�4M�iZ����Y�U�XRE�.*��H��(2,��Nhh&pT�̩CiE�V�^��EId�)Ah��R����huT�2���Vrʂ��DXj$kC	)�2�TCUJ��Eh\�]̶r�*#8�::�MEKD2E4��IU�w�2NV�lӤ�9GL��!v�:!�5LI4�.QZ!P�B),B#DP��Q�����:]R�ie� ��eVȊe\*�Q"��vkJQ++3�E���4��`��ژ&�#�dII$�i	$�֙bQuReJqP��]2.UU5&�%Ē�E|���A:�!YI܇y��U�_�����Ȯ�U��[���#J5ۇZ;�Vm��Z�\]n|���Ϙ����2�d�Ȇ�G~���"��ת7[9kt�ͫ�E�ME�i�g���M�=9�R���۽����f�U�����x�'g>\�սP9<�v,�9*L�(Y�r�JW�N]v^��QV��%]=�������}�x�g8-3C^�!� j�9���d�39p�s��{��K�X|���Q�en2�U>cS-sӁUݮ:��*�
��O)��[�v9��梷Aw�ʡ}Jol�X|�r������q��R���ؚ$�w��6�K�*G��uq֡��Nm��͵����dc��-�|�3�cg�������Oe������`���0��Y�Lځǝ#�p�M��="���v�z�
��$K�k��Y�n×����ώ`J�V�o��X�\.�����2�����GU[F���M܇�3���ƂNa��pI�x�(��FN�f���^�u��m���J&$m1K4�8�:��&R��ޥr�A�x��F��ş���l��iڵAu<kn�N�)��OF�n��q�a�|�b�-���Ѡ��T�x`�ٙ��}Wʙ��(�'���C:p�GM��\Ș����/��@K�s޾��6k�s�@�r���D��|[�q��S"��6H���NI��D�X��e]%�v_���B�	G��s)t����t����u^F���k]F��%�"�K�oe���ob��2^��c��fg7����2w|Uݙ�=EJ�\u�	\>3�Qup�2�^3�]��,��rJ�>ʮ�}6[�V�
�d�����O� �֋�m��I9ێp�7���J�Y��&ugڋ�*���r��#����VF��Uk�'uB�
�7��fv��oQzs��ت��]�k����_ZSs�mM���ִ������ײ�jw��Kgi�u
�:ƥ��9�6�Z�3�V�nM��V����vwqj,���J����`�<�V}ϡ��m��1�[�v��*����4Ak6�n��7�}͠g{����X�y
��.�rg��/(��=d�i߻��T���M(�X�Xt�m�}w�&+��Z��(i�|筱��+0���Z�ಒ��b��R�q����]ֺ�T��Y�Ǚ�p��},���I�}V;��:���b2�<C����w
�o6��r5:�%m�K�	.Z��r����DD��u����]�}ӔgGm��6��No�s�;O�Y��Xj3�m3�Q�dQ��l�<��W;s��q�J��%����(oSo����u��b�ۋ!V"�wD�9`7fz�Q%u]v	�G��܍p��m��浝U5��Y�ac��<|7��xg7 ��x���q�I-�e�n�T%��6�j-Yf�.1yZɆ�#�p���fv�%'"��P%'7�%l�L��I̬�\�嗽�%99[��*��?J�{S����n!P����5�s�SUط���{�;T�5��8��N|K%�5��f�s�0�S�ϪB��)&�9B%^濥H�eꖟό��E��l�ϥ╒��f�#�_oSI��;Um��r����\e�ՐJw�pٺ�)9xWب��&���ܼ1��NBt' ���B�w�j4�y����/c�ϔ����*�_yE��~�.���k���V��s4�cYY��4��yAiz�	�'V�5qtk����z�]A>�)B�Q�K�e�� ���xF�}�V�]�]4�����w��PؕM�8Y��������d��zfv���)������lӐ b�"{����ٝ�'U����״�Upێy����K��N.���Ov��\�7EHO_p�w���_#t1�9	;9\�^��жyk��\�҉�	�l�|�m��;Տe�p����O��?*��8�S6:�74���wp�Z��t�4�qQ���9:o����&�N�A���/!U�֮)�vDvt��;sv��ej��8���y�������QXQc"��>v�m��X� Nlv�Ƶ>_�X��B�Vd6����E@�:���X����=��t�y����h6
��.]�щ�s����C��k��ε3�\I[A��Pa+S~ͮ\r�o�6**+����'+���cUo���~�sv�Os�m_Y�*ssK�����\rO��5ٮ\F=yj��Ggc�;�q����2�=�:�}�^i[��_!zx���C�j���+Z;�8޼nv��IT]���+��Ln���=8��LJ3��S�We���P�H<�O�r{Iu�	"i��f� �c�8Zc��2]�=Q�VN;�9jx�Kv,d���H�fp�@dXg1(��Y�/�*�8w,X��J.-�g����m0P�h߼;#�)��{��]}
�_�W�bMV��;�jJo���~C��d�m,���S����z�q<)-:uSnLJ���GM�/���E�����z�i^��,�ɸuKp���r���v��u���!�[PSt\�ͣՐJj�LU{[5����7bK$��ٗ�Kq�"VE*@W�OTHN���O=-|&f|�ϖ��gXfVd��ǽ}�Φ���T>�ě�FcY��2��J�l��x��-��̞��Wk�f���x�'es�OB{w�c�g����N���/����o֓f���ټ��m�©�\൬��Ǽ�����'���*9�-9ݿ�_M�:S���7:�U�o�%��N�`s�u�' �r��wE���b^e��j����({y���xlԭ�@�Mz	s���}-��JC/�u�N�t��^E�����=�����#�V-'35�l�8�6@�]N+-����m��Iowrl���WWC�b�KZ���OM4���q���i؛��[	2�A��Sj���iwJ��=��I�N���Ϋ����z��1�X(
�7�4����P7��n5��V��X�}�Eݴ�q��v8��}:��E�׉�v{�����jg�
Zӑ�)_*/����ז��UP�������l�;O��������Ͳ��']d��C���]:F�.V�����g8kr#XyA���e[�/��c�>�5�$�32�?���I.�4�	=Ϡ�h�ʗ�� ��e�&-�8�ڤ�蛕G�k�J]7����L�ym���6�&�8�Z����j�+��*� ʸ���}`H�X��cZ����7����O�zz�&�;��KݛM�[�)	F撺$�V�ژ�)��ޜߧ�z���ﶱ�i|�4�{�P�����Ǭ�Hr��*z+R��-�6��t�^�z��f��yQR��G�	]h�m�����pێy+#svjz�u@>��t�.�ub^�Q��'%�̤�����x�'t�¨��ya�h�P=:�p�JU��7�$�u]�9;Ҷ�8=�/+�����|���Y.�� �՚<��u܊�N�r�ͅK�+�����ܮu�G7�����9��S�ݬ�.��^��{�զy;ɛQ���{f)���g���ʵo���4b\�N���#[GM����rj"qu��������������8�Q�R(��2j���r�gz$e�.��}޷��*�Z�7�]�=�.�m���U�b���h>��4z<|ֿfyIZ�����f�he�s�a�O�+�V7o' �>�9�.q4T�k��(�nS���{�5>ЕOZKbvua�n��)�OJ�%_k�C7�*ۉ���s���E��i򣺯���dw#I3ڢ���J�V��`��S�YL63���=l7�	�c{�U����K8U��b�����z�'R
��]T�6q��f�v���/Cw�Ş����]m��/��ɯ��5@�U��Kae��^�਻��Lf������[�C]��_���M�4vcc��E�=�%�q7��Myηjr�����V�\Ʌl�N7��·M2]��ӻU��2�t��ު�\�qWK�p8A♰������t#{��5\>Q�`d#D���1�;E��J^�ׯX�8
ǵ�ow*�v�k弳l�;�GAs�
[���$�y 5Y����èH�kZ�H�}�]c���9�X��n�X&B���o�c��G�q�Ĝ��P�Q/vns����36�1T�훭<����/�W�|5q�_j�>3��E��[2�^)E�������q�U[��c�\��� .uqh�d�4��tf��5<г`�y/:y�㓘u�S�=)Rv&���]��.��/h�������=D� ]��-������
�q�>���=U[�;,\���޷Óa�W캬΢u��E-�5oA^���ë��ͽ���y�jv�1��h~�E�Q��T���릶��������T�
pZ�lu�������ilT�>�g.Ν/�X3|o�]�Ҋ�]��չԾ����s���v �]Gf��[Ĭ���Jwl,��U�V�M(g"uEFXϕ��t�H��ΰ�.	]�3Q{}݇1T�m���g��s�c�OWt��n�&9��Oj��
���fս�9a���kA�.���㰕2O@�S��@jE,�Q�p��I朱�hP���D��,�̅���rx��[�<��^����j� ��Q,Ȓ�g��̤{[�h��4�i��7f;+�-����d��4��X9uO�C�6]���1�}��:��}kB��+�����p��d�..}Dm��k�!�g!�}���`�S=���U�ӭ���$��Yjƣ&�5�g"y�ϵ�{��8�>��*N3Ҡ����܁�e=�IN�]�N �rZ�÷n��}���u�+��蛒��GW4���:���_`p��t��.�y�j�6t�k�s��ns,Mub����[�g�-�k�7�k0I����@����w���8�m%/9��cC`������})ot�q���:aL��G�� ���^�C������箎�`§�"龾�_�^��ظvĄ�zG�s�H�*.��]�,V&oByV��g_�I�.�Lt�ˉ[����]oAo<��k�9����4���}X��^2ں�Ĝ�M�<�\�IS�+D�D��;�8�>�e���8���)��F��[�OܯN�k��2��yilmk�J�/��m���+�X<z��f�ګ�!�B�K���Wv��� �;�RZu���r����F@�[��8�}Pu+H&uԬ�P����gs{�o2Ԙ��n�"�L˥,�&m��WTy�+&��(-��X�h�o ��Rp�X������S�c}����it�������"�K�<�ѵ����w��
�r8-c�"/DtL_&��vs��݄�yn��j�������|�q�*���}=K��r	i�]�O&&�|KX��ggW��e�T��Y�c7�����}a2�C�O_U�&_E�kQW��}�k�G;���,���^�YR8�Y2�!�1�G\�7]e��0y��q:��[�x��g�������{��s��ƍ���S��Z�$%q�J���.v�877���6�|�>υ�Hslt�ݭ޷|��Sդ�L"��2���9�\+WWɾ��nk��M=ѝǊ�\�U���\M˨*d��@�$��$�a�7��	=��Ca��cR����Zv���O�o^3;q
����G�eE�]7[�q��SR*-�{��̼7e�ny�a��x:Z�����)7�����z�����1{����b9��r`Vg�j�j�Y�ܝ}$�άw+v�i�"u�}K,�Yn�\zڻ�,��6WeZk"]v��$��y֜�zZÖ�g�H<y�� s�n�}%�#��gd���u��}�iD[�U��򭒫H�|{#k��)Q\S(��[k�w���p����f��U�d7۰V��B��#�6w�(gu�5N�9|�̾�z�FQ�:�3~��h��׽�>��/,7�ibX�i����d6A�]"{[�:�s[�h�aͣ%���ʢ�� �=[�0Ra[��*���u<Q���_hf����KB<1��z����.[�wP�x噖���X�����!���FRyC�P��zVz���/p�s_F#�1�U�Ν�;*`)ԕc�ko�C�O-�C-G�_,�m�e<�$)�V��h R�yZkf'�|�e�P��I�[��VƎ�Y�U�t%b�q���)1�^�᱋:S��Tt+*�=Fv��Y���g�"B���`�
���:�f���ϱ���p��]�?g-�]k�Z����%)K`Vf��d��gt=n������kg/wziU�i�����9�M��Z��`j�%��lmcc���K���+�6���5K�#4(���m�Y���� Q��6��fF�f e��'��3&r�X���é�򬂲��ja�7k�MX��\8��.8�X��l貍�S�+���+b����U(sa����>�/��q��d�x���d�Gr��sv/����	�Ɍ��B[k]r�7�A��d��m��R�\���\�D�������J�'��r��~*��j�0�
�s��!T��[���vhXޡ5M���´@j�j����R�.�|P�����9Ǣ|�չƺ�����8�jMB�bЈ=7�2�WR��4`�6�]��A����t�:8�NK-�}��1���]*�rdL�WEt���]Q�8��W��f�c]f_!x�S���A�`����_N�6�jo���;��s(^VK�8�W39H�a�l��xd�����9	7^蓫�՛�;���m�qR�*'�Wm���5�2�ٴn�k;�K��\{����b�w��M�իid��5k�a]R�'8-��׌�v��;+�=��"���wP}%l�+�_i�YA�Y���"�tt�RR�t�Wth�n��h�t����t̚�[Ļ�3ҝ~��Z�=���h����@w(m�����A��WcSn�-��+u�w4]	�w��+@v�Q��n�>�!�%&iK�8l��V%Ǣ�X�h'/M߅��H�6�2ʟ)Z�3�;�2ħ	�U�ܨ��Fa=J�c۷�]��%q��iP���B8�F�D\Mr��ud�oN\݂,P|^��H������Jʁ;�srf���7�4+��o�rf�����6R�[�K\�5({��۠f��K���U��>1"�+;B��ȈBH�J�ZW,�$]ӂBMPI9J�R�醂Wfe]�,����*"��.�4�EUN��3Y��%Fed�*'��*��I�0�ATGe�Ydf�4.�֖aZ�#b�9g��j��*Ԣ3���P�H��4�Y�V,:BMR4��% �T�Vt2(�L�je�X!&J�%UT���#Q)R���Åˊ�K��S���d"KH*�KZ��$���8��PU�ď2*siy	ܮ\�Wq�p�Us+��w
�Ҁ�T%��ɹ�$ʨ��%��Ą��V�ft�+w`��В#**�V�Ե.�Up�RL�_>z��Ǟ=z~|��� �Ge�J�������*��D�x�}:��	��9���3{8�����JS�-�WՕ��Û-�0�Sk��c���<SID����O&�1�!(�M$ⷧ:��J�xCJ��lΥN#o�v�����_�I�.�N%dTvu�2mR��⼤ޓ�Z���Y_�Wl�d��r�7I' �n9��,��t����VrK��0�ؓ���c���?-�<4�=��{�ى�g��&�;<j��]B����on�	��rjqu��\��K�2+�x�th�
�Ԏ.p���p�ٻ�r,�;���<U�� �t]<u$����N����/!U=�+�ϑ�����{���W�ƶ?���:����wbm�N�曓�N��,�nTC�GD��;<���a7�JY>��ݝ791}�>�$'t�n"iC9�Χ%�;O�܊�ѣ#��}ֹ��v,��6\�V:ʞ��a�9��˸��<�*����!�]v�X���(��3�0-Mlb������f��r8�M��7�l�9�8M�r��]r�#�����atKWPN���8�c���5��$K��#Ob�þ���e�E7��%v�m�O��Xk�or��;����X5���J`N]��F�Q��d��V�:Ꟁ�ޔ����O�l��^�31�a���f������u�a,�7���Y�N��N�(�YR�d�<#A�x��Ծ�pA#~���tw޹���\-?c3��+���~gB����R#����{}yG��x���j�6NDJ�{S��ns� �V��uͮQ&1W'�L-*��5t�pin���e4����{�i�׏eu�M�їUm��z�ꭡ�7ù��Y���/������Kf_N��+��yݪ���3o�����oP9s	�M��N@�}C9�U+�C{Kq4�K�̧�/%��\��̅�2�d���wk}k�X�t��[�# �h���Z�˵gͫ���_ɸ�
�c�	���5����<�������U��m���Y�Iq}}��>)��\�ս��^������ۥ Ũ����d�������ޚ�o[�A]�fZ�� <s��:(/C�an��R&�n�u2V�m�G6�X��Y���vb1�a*"��c����Ƿ8��&�W$}c�Wh��ܶ2���Ph_PYj�:5��nhzGf�ďmr�&�s�ʝEk&7*C�1���t�H�E�xil��N���S�s+�lu�k�x�F��fi'��wYZ�-t��{;��+n"h����/!U�a�#�����;�����Kg/1��Q������臷�������M���v�5��^�5��.Q�br������}��6����`�t2���S��y�H��$�l6���N)x��׍��e�����z�u
qN�Ne��g$���ਥY�Lځ�y�ȉ��5�{�>tV��񊓐T�e�,Y�\��[Z�J�+vK�{t�Ֆ�wW���vF��}9�ws�v�Z�A�I��nn�{�m@0$�/�Iuk0횿�6t�k��RQ��ѻm�ԺPα���������L���鸎��8�.d��wb��m#�6�q�{�o���q˺o���0�VA�*����E���)7�zu��o�%�M��-��V����V=�&�`Zd��Ҁz.��>4ͶXܹ�h��(%4;8���g���,���^ĞϬ�d\�gv>Yf��:���nb������.��+Wb�]��w���|qp�w�n��S��!�in�8�u�J��%�-�Kf^}/�&�.rg����`'�3�Eس���ɟv�����4���[*z�.�6e�D��\j�S��u�0�h�=oh�h���J�[}Y�/��^��QĜ��k�;Om5ae�g3�J�(	���+�XA��z������x�'g!s�W�@�sxc[�i�|�|���5ن{�k����nwU�=�K�z7���yS"'�ld�|�ִU�r���\>ۿ�`˥֖��K��:��V�|���\�p`�k^*ޘ�����7̳X��������x]��EC��&8��u������I����Fz8u����!���8���,���7�0K}\��M��A�Q�vT�唛�i�B��V{;��d^���WO7�f����$����e0�;Y��P��m��oU�׃tD�≷7-+D��]��A�`ec|�W�v?5������gij����̭�����7P�+�t��<8�{[��ՌƱdj�f�|��Ǵ����{}\��t2��N�4&e�+��u䭃��Q���v�r���VڢƤ�V���1��[s ���r&_r�'nH�t{�qfg�(��O �+W|���򥜻$4����>3�ߓVj/��P�SS��zOόF�$��|+-+�C�ۮ��t����K_��u�3�
�������q�y��El�XxW�s6�599��O!)�~�X�l'���wΐS+ �D���p����P���^Z:��T�ı���q�)��󚇙)�nد�/hм�[��}&v�ݾguϯ�($+���)�|g�,�&̸v���c�u&t�J�s���;Umj��BW�N�@|�����_ȹw�����p@Y�,���V��fY�����N��=�؇4���5�x���n�7$��ܬ�uYOK�Vێ�k/�������4<N��~���w�\U���)v�?M��M���g!s�G>}���55�j����y�Q[-MI��&spo+4^�ܓ	m��\�m���d��d޳Ҩ3���]�ӂ���hՋRzzi�^9:ݦ)�iV(�P�\�R���P�F��1����*�V|�v���KS�Xv�N�qm���m�(��+���+2���txY
�i��c\+�3Ш����;�:��T�
�WP�^�˃��k�/|���8��I�k~������):���,��T[�w��}�{9b*���:�w|ߥ0�9v�--�h��8<�M(g'TQ���-�C��r	� X�#�O���s�`H�X	޸�CV��i:��	g���}����q[���]kB��n�s(�5Ac�%��e�@���`
gd��o��\u�5����}Q���N��]Y��[����ֺ�4�񹣲5������*B�=o�FY���}��n�8��W$���\-1��´�nMA��;���v�<��r���}��X����f��y8Ͷ�Ζ������"$�ǎ��yVJ߻����pg2޳̙M%/9�{��fh���LА�9����USo�DW�J��DOH�_U���x���o��{�}`�}�ی	{ҵ��p���zN����^�P}H�Y��;'1X_R9��|B�0p��^���
���e*��r�g��t&���Lm=�dsk&��^=�O*���Vmuv�ӧ>E�12ue/'><��� {��#9]�ɩ��S���X�n��Y=���ܜ2���
���]�<"W:4��D��!���ѯ)�#W�Հ�1�Co�X=��9%f�L�@��'��bA��YD]]:䤸SC����x�7WS�&�}+/��1�6tѝ��#&�kΗ�ڌ��J63������o�W��\W8up�v�˽X3I��\�I���V��5�	|�[��V>[7���{b;m��S��
pZ�ltVH����x<��Y]�Xq�m��.wlq��whZ��lՈ�x�g�r�yR�;�c��½�G23�]����Y�GGb�٭En��0>˘�w�m��8�Ɗ���S�����O�b��ۧ��s�{*ߚ]��,���+��7;��4����q��|��ⷶ���&�.�K���z�帜�W�Z���<���L�Of���(\v>u��L���{��� <���o��>� x�K&ze�q�*�E�,�u�S>줾�x��&nR��QB�ӕ��q�j�T[[�>`�;�C^�p��y�r&�Z������X��EA�����0y��\h�ax婹��>������W=:�]�
�V���-�s��-�L�FfPy���p��V�W��nMB��8I,\pIdB�v��XI�X�A��̸�iU�g�/��l약Ӑy�gFR�n&����1>W��쁐j���5�g�"}o��7QB�Go���\��Ϳ��hw��#I�W��#'���- ��!.��O��C���������.�)�=�Kz|������g�=��d?{:g>�g�\:��	��'��¸�l{x]��l���+w=v;�o�-0e �x��9	����~� <7������L�έ�T��0kO�q�T�w�Oz��Դr��b��V�B�#q["�䭑�z���̱��
�^�>�P��]�����]٤��.�n�P�ƈ'��Z"����F��{�rr �͗:߳!��]�t���5j�'��]�9�^�{ӓ���Rg�.�ʆs�b���l���|����G���ZkF��{�˖ w�C����\փ�y/1!/�^'5ߋ�7n�*���B=��{uw��].25��vl��nacI�-	h�$���R���u>g�A���P��r�s��7��(�u̪�,Wy��IP�6kv�����J�6�˻�)�k�v�{�>H/�<��gYW6�A�gNYxqc�zL�`��U7���zǲ}��zw�w�����ly��u�OV��T�p�z,z�������NB��KTf�^y��I�F���7���a���ra7����H�͗Cõ���'��Ey��F���{�T�Pt#z�s�[U镑<��2�����S�:���;�"���Gzm�Ù���L�˿V`�nB���#�n��:;�2!�^K��zD�S�����Z�赦����Y)���{Cг�*ȋ]�^� 7��C���A˵~�[���ܘ����7e�[��M�η5v��=Ls��r>�����r��X�%�!H`�/�
t�[ّ^z$��gG�_�E=]yw�v֏7^`��e����v��H�Ui ~���ù�Vg�.�=4E����fo���5pPϹ�dVW�������wޱ:c�lUê�Ũ��LǙ9�7P6:5�QZV�����>���FG
(9���(2�8�'�lF�i�1���C��;��*g.{nz���uv�wy�*�ú�.�\:�6qY`�|�V	8��Lc���`3������mG��t����G��i�^�N�X9���5s�"/�3����.=��O���:�<�g��9X5M�K��1D�9�NN��.Kp��&�=V� ��d3{���wamB���ٸ������m'���E^a���Y�};�S�{ٟ�(~�|��I���U����5����R	�-�X�J��e�*~�pS����M�z��j�2}�썙��ʑj�������ƃg;�4�FWeԯ)R�H�~&m��>I^X�޹�x���#�&2�[@��~'�c�a�\��v>_Bc�ʗ�j���W���x��ٹW��l3�������ݹ9���u9X�S�ؾۨ����1{�j��
�������sj��F��qd{]���jtXL��o�А��{�F��
�e��9O�4�H�^��[>��t�".��N@�l���o�^[��v����`�~�'t%��w��I>��j�V���׆\�aB�
�S3�FzI�X9\MCο�Jk����{�������/��y�w�v\���Y�@��?K�/�M���X�8�e��O�&���/���޻>�:�F�B��������b�I��3h�A�3�NT�~/��M��eD}�hW9L囯g-J.k��>��;z��{�>�����ߤ��(�H�������U߇�.P%wv�e%�?���+qOҪѥ-����UG0R�˽���3MF��&���K����zFjv�����Y�D�C�*���f�hN�ty�S�1;T�$Ek�'z�je���l��0�����h
�l�$���J��<�.qM"��,��f��"\�	Gx�Ҽ0�*}�ebb�1S���q�r؆[�╀k�T�y��Ԗ>[y��*Wi�R#�itsXvo�9#�R�������ouV����z�{���c�|y���n�b��fG�cν�JY+_#N�z�`憬�z�ne�G%zXj�(N���v������n�dt0n��(9J܁�2\����VQ;ϲ�S�.�����g�]��o���g*Z�C��ԡ�?C]u	*�z�&��Č����^Jb��w]����9�v0�gGk%�s;������p;{]Ӂ=Y��'Dhnا���V��[2��������/��ڒS��c)RW�8ynˋO;	uh�ntJάwI�Or����	-E�����L�S)F�AT�q�
RT6i�ï���@8�.
���I�q��Uf�8����C�(�Ԁ�F��l<��}W@.+5�
�kjm�Eݍ�#A�H�Eӳ.�dGW%
K��&�eu�|�i��=K����{��]��	�\�E���e��y���Be-s)R8�e��uqݹq�pv���Ճ��
�|[u%��ו�)Ѯ�UhǨ�[��e�_[�Ώ��3���j��m�%_ٔ�3�n���U���Y�j1.�j�z�ĩ�u�kwt��N�HD�2m���V��W6`�xi�+S��W�D�6%>�n�L��qD��	����wK΅ɝ�x�,6bz��m$z�(����<�yo���rJB���"��W*�����3���O���R=iwX�	'B�YoK'��l��͗�Q�f�ޱ�t�r��.�'���-���Խ��S�>j��p
���/�T���K�/o�n�&�r[t�p����WG����gW��f�}�]$��$�:�6�����=��}�ۂ����ث��:[�<N.飋�Y�nmg(���[K��v��������Qvl����Z��x�%�����媕��}�|����[g/[�j]��oF<�,��t�s���1^�,�K~��W�sX�EVk2��4�`�7''��i�Y��/��Q��C{I��H�L�e�]Js�b�f�H��`ة��NgKVp���N�4����%�L�h��#��	لw�;za莄�{�����{R҃2Hf���1�/1�
�깡@{���)Yƞ�����#�/�]���cgZ8z��-�ѝ�>T�]��b�ѽ5ԧp�ꙇ ˈ;�!gif=G�价&t��Wq#,��GN|�u��&��ۅIu�<��z��FY��#eRo<�ӻ��N=B#�1�"@�JQep�ɧ$�����se�eU�d�2��Nt�
�ls��`�E0�g(N˅�MPJ��:�UTbPZ�͗�'��(��H����*�UEP"�ulI���(�Wdp���r��*8�q�8�T(�E���,����R�"
*9�����%TA��Ws<�QQr��(Vh$G.Y�E�AUs�r�T�!9T(��\����p�Nʈ.�J�V�����dUp��*�W��ERL"��
�v\�������A*�Iu�r�L��7P�8U�(͓�9J,�!$�A�K��fr��q"+D�{�Tz� ���#$�N�U�Lê"HH(�ػ��gI���E�ֲ��gP/�k�y��{a�����dyf[u2��u�voH�����oa�;�p��I�4h�WN���C����v]9�u��\U�����>��T�w��X�����6=W��}���G��S��=8Vܙ�{u��:��j��{�'��C������B����^ǲ^wf��-jU{�B�=2}.���6hI�a�
�9�>�*v)��Ӟ�������f�o�)ot����E{�(1hCw4@��^�cSCǢ�w�	��ze{�+�}';˥^���g��W�=��ǒ���&�����%���&7�)�l��9���^R��yf�����x�./����&��=�O��3�؉w�?��}����]���A?_Y=bf{�^;t���|d�B���Xߙ�F�����2�}��.���g���d�ڡq�$��]�����sܔj*׶O�]l�ᳶ�ܯ����r���#Y�_�d{�/^X�>��r���X�m�qZ;��(�<�މ��t=�б� �s�=�����c~O�+���z��r�Mz�eb��76��e��>v�mX�Y��>�3�iҋ��~�g���#������r��87v�EV϶:�lS��U�é�W�7��X�4T�F�z,�����ǯ0��Vµ˹�@g@��nu*�Q'XȨ�TT�C�׻;��������K���<�{R5�1.�^Ѣ�!��H�B�ww�F�|!��T�
�`7x������*�z��sO�����f��u707dC��<nmW�]z|���Wc Y^>�Gh{&g�x�jw�Kޡ��|2��:����kht��O���.��\d����4n��=�����
Dx�hv�ϊ��=��#�֮4�,���m��t 5Cڬ�v���ܵ)�U�=蚨Wwj�3��Ҭ�]�#����O��l?W��G�����D؆�d\���^W��#�.5�C�W���TW���?��}?������A^�I�>�[���K\��S�;�ʔ�5u�U^zȽ�9C�Йj�S��K�S���[�9q�_���}M�:}��8:�Mˏ_�����-a�7W�a� ��#}q:-ڸY��&'��|>�7d5K��|��@E1���˱qB+�~F��w���@E㝏������2@Ϸޱ=���.e9�Inp/���iᾤ/�i�)��]^r���]���}���B~�������=��c���r=Y�V�3 $�d�hK*]��i�eI�G��}K��tX�)W�2#�M�M_�?@c�=^��˽�~O�!��ߘQ���B���Nof�ʜ�7���s�o'��ur�MX(����tCu�(�M#����y�uJ��I�S؅z��������o[���[�p�bCa޼�/@R�W�r���6H1C�]cdl��XYʼc��%{�-rX(*s��E��+�q���tޓ��^P�%�M��.ss�ȴ��P׮=��,����
��z$���!�U	�b�LR�"�㸪��6��th�zk� ���q[��nN���]�{ٹp��>�aVv�����L��{zrp�n��� �r�����_pV:}��8��$�yg�}�W���c{'�M�Ca�\�-��=��]�.Ub�8��ʣ���k�b���4���uN��Fwā��7^`����ww����N<��#�:O�p3�f�<�~���%�ak�8xʮ��}'�_���^�h�q7��#�T|��ߡ��%�����^<j��2�;����凕_��;q5N}�]z�N@�s�[�NeG;���H�����ŐMƯ	#ʦ�����*��#��׆FX+ӷ�!�A˿X�8�X{'ג�8z�"s���O3�M7���;���/޷Ͱ>n;���mt[��G��T?�R�&���ݸ����Æi��&��m�5ⷽx�E�{���{÷�s,�C�9��eQ`!�0�&�|�u��r���F�В���ڴ�Ǯ�_T���4�oz&0���q&�Px�,��۹V�tp�N���ʍ���,�y����d���p#J��3{�7ةp#:��f�h8�����I��r�[�l=8�}�ka���#)�%��z�'F�-�5R��;V{J���Ep�E�y����>tv;�2���+��ܼ�Bf|�K��'K��{��ٛ�=���|�z!�^�񼒆��Ȭ�{o�!�N�Q��	��[p�1�L��W���3��p�Ez"����fF^a�9��FK��lF�i�1>��d��S5��]�c�z��u�� a���M��ʮr;^���Ǌ�'>Mg����Ǉf%l�9;��9B��X���q�.�Ej��!{~���.)����r�5{	[�g�O�m�ڎ����+�޺���ۿ\�%~�>�L�lK�`?~��x�t
��t�{^a��.�7���B�����j�r�����9؏y�X�޹�y��=�K������]#e���e@�w�O����V��������{��P��˄�?f Ϫg�iǎ�Q��ܜ�C�U��!+��6��v/(�U�)P������d�4�3N,�l;����k���dQ�Y���x���u�o�����:��:�>�������yu�:r�������,�J�v����{,��O�Ǭ<���|t�����
zE�΂:�ގ=+Y�g��(b~�[3�k���q���w�H���,�N���`I��'e1�s"�����ev:��J��Ũ'�8'Awۄ��+��q���c=��0������T�w�z_D�gֶ�W�pq��	Y��MK���;��{��n�b�>n&�k����#=$���q/:��I�+�9�K��Vw{�n�J8���9������Z�F���ޝ�ᑁ�傡迅��=�`۩��p:ӽ���X���[U�S��NF�^�ez|\{1O���<��OfS qAx\
W����4d����&���{���}�ϫ���v�����o�ߤ�e�Y# W� J}�xO���s�e<ҷ�3��p��ν=r���깾-��>��doz����̋a�'[TN�I~���o+e��o�"���6)LԪ^�E6�9g�}��7�W��zu>�48������6/ ~s��>˾�x����*~
�g�w��r`��.�dJlМ5Kλ��+�)S��<s��Ѷ+���'��N켯9|��F���Dz�qV�-	���U/Y�l4=��-���q(M�����.�����*|R�zt{ր�xd��[2��W�W��D��Đ'~�o�3}�7�]ow�I�R}
kς�n��.j�a?zԏl��3=툗{2�
ߕ0�
����D�cZ���ח���'��:\�l�m�jS�G�H�Ͱ���޾���7�#�0�غ�D�A���u��C%Wyt�����5��
�õ�9/��Ht�.&*�R���o��o�^�_��4]c�Y����L�HK]X�kc�Һ��Z��V��l�,�'v��]9�F����ߒ����=��̱��x
��>�{�8G��P�%:��r7K�\��(z(uz�/%�ʠ�l�g�zox�#��{�1�g�~���sD�@��:*%_�����U�C���
�v��'����^�ҭ��Gs�ٛ>���#��}m���]v�<�{���z�פ�߫|�[1�a��j���̟QUߝ�a�׈0-�H��s3�����OuQ�̫��>�i��������x=�;�$N�n�P`n�z.��Ƚ��>C��0=뺍�鬭ʒyx�o�zM�����P�C}��l/;R�Q�khv}LOdU=o{ӆs=U������M���Y��
É�
�Kϸz�'K�Ǿ��{�o�d��Sq���Mm{�j=>����ǻڙ�*�� ���)F��q�sN��\�����\�{��W���{�Cm	�=UY��Ԝ���qM�:U�(t�G�������M���o���p9[�g�ΟG��ު:'��by�R���NzP�iy�bD�.�\
s1)z�t�6�a���d{=�nv��[0��RdR�
����ܵbؕTov
WD<Fj�?�,z� )<Z�E�]v/�]��R:ȶ�룶T�S��h��al�����'i2���v�5��y�¶����;�J�[�����s�m���ު���p�����)�q���ƺ�i���.�x.�>��r7֤p�n��NPb�	��P�v@�T�q�=oN�٬g=eVNzB%�^S��2�(~�$��N�]�� u�!3-ՏP����_f���}�������+�=�\2Spq?cc~�#��u��gL�ެ��� ��a}������!o�bNx��o	@H�Joв����!O�<T���z�?W���o��˽�H/W���}�nvp���;U{����x:�U�J���Q���h�ԭ��z��=�b2~�AF=ޟ�o�z��^i��3/�$�UƱ��� ��C9^��gO[�p�m�.�%�=�U�����ǟ��g�Fz�K�W^�ޯL�ϼ��' �n�\�
�v���z�A��x��w]\E7Y��rQ6Nϵf�~�������͚#��qn�N�S�F�����}YмZ��ꛮ�םӊ5�y��t�6	��z��W���}U��p��~�ˊ��Λ������h���U�����y+g��*�U�\8]:�MƯ,�mQ�`d<�0u��%��H�[}�L�T���(��ry��%u��}I�?d��bͣ�|���w����`�7l�գ�/$�@�,$*GR��0�KO�X�����D�}��<j�5�@�V�aN2��(�:�����H���+�������V��}�۔���Js��M����`�O9L.޿�iX�&����[����5���1���s)D��Hϓ����~\T�G��(��}]�'"�3�`_���
���`���S���D9×~��w,8>��������xMV+�k�k�#��@��E��".>Gn�ϰ9�b��HT�~9v�տ-ۊgWx�7��4����\]���)���O8��޹�r�ψ�9A, �T8�Wt�}h����{�:��7��}�r+)��^��w�e���V'�ۗ�# HLϕ{�Z2.ۛ�\��;r��3ܷ�3���#�y|��6�n=�^�$%��\�O��`��U�KeB6߃oN�]{QW�W�C�PW�ME{�ddO��t|�1�jP~��8��9�8z�g�"�����>p?Z=�_��2^����V7�䎖R��X��X��6��� ���{#�9r������l-D�l���W��j��OH��[@��mOm}KԹ���V��nZ��D�ҭOE����j�<%�&��Л�����y}�6f�~̩��o�i�G��t��0�����m�W����~Ul������'�ǅ�(ؠD�f�}���4�X���`�;k����Vw�d�쭹K9��BV51�$�x�ul˂İGv�:���bh�4��{���ިW��
�a(�EÚv5������:��D��oJXO2��t��S�	�q%w�w�B���p�{������]���2�!�=2G�%���mԋU�N�!T�'f�Y{�}w��l��8=�ދ���L�!�U20�nC�Oوo���}j��n(��nN!��#O-���}w�Ҟ�o9W��=�5�잮�[Nw�[ �i�i�q�B��
tXL��v�T^���K+��ޮx����kU9��WKȺ�8-_�;~F��o�G��c��e����7�s�Y��1���$�XD�}�\3�<v@�{�9�ھ���lO[���n�M�h?T���.y�Ӳ=x*M�#���]Ҟ�^ћ�;u�"00<�T=�p���ǯ6}�x=/������g7�%z$�ɇ����9��^���~�-�f)����2�UOvS P^�����ze���|�f�^C�,�v2S���^d=�=~�w�|=��yV��N�YfVH�J2SA\Hޟb��j�U{d���L�J��7T�^��.�=~��-߸x�����w�X9�Y�Ȇ�b�g�ݴ�.�iU� �FHB���^�^���U/
�)��a�����)��{ا�=����6J-w(4̹\����P�t�b�ϏGp�3د�ܴe鬑r[�,��9݇�9h27�a��0Î�l�gW)�j�stw]�Wȵ(�.�0�r����ա����J�9w�}�y%6�9
f����语حT�4��RXaw7��&����ϣ�lC���e+�"[4$���T���gإN�{=5E{rN�x�q�C6�g���'��$�{ p�������-��*)z͌9MZw���5X��j���GD�Ȇ��������l�W�}XM���]3�˰T��al��8N��W�$�W^g���jǖR`��Y���9�����Z���zfw�]�ͻ�"�/�k�te?H������m����p�V��\��r�ƥL�/ݑ�y�X��K�P~�L���̕ �ν�g�߷�]MƮW�ʡ�u�FNJ���K�Nv3����l�/7!�7��#Y�_���
�/ޮ�|P���\2ǜ��{c�{Eh�<��v�������׸t�B�d���?M�,~u'_�/�-�yy�om��3{��S��W�G:�nm{n�dp`w`�^��!�׷�2��K�z��K�VM��__��)��왟F�9��W��)C���W=���3q�۩�T���E�+����w1���(�^4G��`��L�Ʀ��.���?e�3Z��JYFN��rE�|��~*�~�?��ǀuu�Ժΐ�i
}t�Cq��D���dӛXV����2�݉V��U��E��3��O�{]�ʵ|϶���]n� �*Ⱥ�)��x���\�2�p&ʰ�㩝#=����C���@�}s�8�u��}0_uu���<up�[zkE�A�Y7�"ucv�o��}�WKsЎ�fԣ3���v$g�;+��*ft:�X�s�u�<Uƛ�}�k�oe�ͥZa�V�qe�#8t��:�3)���:��-�[KLo��:d6$̩$V��I�0v�M&uݦ��:O����U�����ؓ�;]ȑy� �U�
�{f�P�A��WZ����7������N�jeH�aԲQ��P{E+nics��C+��
�ll+Q�&�i�c>�6��wy�4jG/kI'�Ud �ޠ�\��tR�m���{d�SN�$�b��܈7vs.�f��N(M*ɲ��o�aR�]ɼ���ȩ����ܢ�<M�j7Qq�?:�����;��o� �����5���z1���!9���\�R���7k�����ؾ���q��]'S����j�^�Pv��έ��� ��7q�'����Y�WVg1s	�qYH��Swק6��:��i�}l���4�������u�Yr��,���v�co+d��coqU��%���׹ɯ��u,�Kw��
�����-ܗ\h i^��U��oj{Ԧ�Ja-����4�o�Z@3Ԫ*ɣ:�W�xw��O�{9�p��]���ɀ�ZM>:���:�C�MVY��h]GN��ss7��`�>U8��ĕ�j܄#�ջ�Tt��ٝgw5����c����u�V�UA�Wgj{Ye
����P{��D�sj��$�����<ꎅ���ox�]E/����V6iR{@��5k��Q���ݶd	�]��������1���ظp�#�����qw�4 
�nj�Oa'�!dL��	��Q�um��o�z�5���e+Z��1��avM^>�*�溺u�V�O��Am��3�u񰭮�l:Ծ��ZL !p�Ui�ZW�n7�k]D9q%R;��#J�y}�U�Z��u1����JX��T��}���wa�,�(�����O��"��g-���31tΚ;r����[��\���=� +�RP4�6��$�(pQ'%a^.�L 7 1*��W��X���^3z��GJ�j5c�yS�s���N����G%�\:�X���3�l�4��F��]���� �7�٭'��PS��#,s�4ae�r�M��9ئ���A�l��D6q.%�ܢފ�����������E��*��K������ż�d������su�_sJ���X䁧B�����5(�h(s���|�:�w�ήp����3��̌A�tse;�33��u�wK�]�7��(<"#�vP��u��*cP�!���z.��yN#�|+�t�,?�8�Vk;�Ffd�2E�`�7���L�=�sU$�}�qs��_�Qr�����VUTJ!��2�9R-�e��2N�P�҂(�w`8AF�dTD.u��(P�AAp�"���)X��$U�	PW��Ty����(r��e�b�y�B�ʇ;J�s-M\��JԊ�^Hr��4��(��s�y��PQr���Jdp�Z�ZQy��H�N�'D��8EA]Ԃ� B.�B*"�P�Gq�.PQ]�s�l��R�#R�h\���:��*"�+�%�ڊvh$¢.UͅVʩ[�����ez�r/	5i�W�QTAG���AG!R�D*�H�Q�G ��E��K���$�\,��G*�]�&D99�r�����/$��������z��"��y��Q�����AL#��P;M��슬��a���z`�N�GAu3�8�GSL�I*L��B��$�"�Ƅ�)����K)��&m]��<O��:���[ה/��X�Ƃg�-��S�n8y��D�>ܴő�iuʸ��*�1���'o�c��{k�c̱��D���k�����Bt�<z=��^�q��9U�:��r�r�+�e�@ �T�������u4����2=~��������?l���/�]'�����ͬ�+��з±`�`H=��H���l}�u�^3��>�~���#J�H�2�=�G��y2v�T9>�r�������r���I:O0SL�Tۭg.+ɫw]{�LNŤ�5>}ו훐u^ϛ����x�Z������92A��R8���$W�T���樂����jo�����(g��d^E{�T�����̐3���Og��պ������M�\��/���T�{�w�F:r=(������2���~����i�����Ι��g��{���Z��S�X����^ o�bX�MڛŖ�2{�)�x���	���~� <4z��{���Ido<+<W�U�3�V�m�X��<�{7��\�ێ�����	��n�@hv��j��|�=u�ء�T�O������
��چ`{m5�����-}�ܔ���԰%��t���wS1�9\���zg�����&u�M���@Yܡdc��[{��F�5g�K���}Q�!���5���;��&�s�S;}}5�87a�m�`�i��k�.��;WcM��H����cN�A�n�s�MZ:�Z�ݻC��7I��&�s���:|�̹}�t���4s��ޜ��>۩� �D3�]�_��p����9�e����n/����I�ח�)���}s�k��k����[�S��S�F����n�{��=�A*�eA���{��_������k�{zu�ߏ����y�Ǟ\Wgnt��մ7�fڎ��>H��jF�*���*�����eV���'�y�y�/ ��\�~w�w.I�_�[�K�գ���O�y9�-��-)����~�uS�Y�=#"����.F�oֳ�%�{Z�E�`��;A*��ʭ00<�9͑D9×~��qܰ�O�%��Ug�pYg|6��I5r�$I�tg}���>�+�Gn�ϰ0��B^����RǱ;�Ob�]//ߩ�R>yۓa�{:v;�^����s,��9��ed�- R!��zsX����V�d����G��Ya�9�^���"�)��^��ީ��o���wn\M�����M��I��i����L�Uz(9��yّ�E6���6"ߖEg��bC~����<!���ٞ\u��;���`�Smf�-���ͥyaV㭬���.�ru�	'HQw����z�S�7�9N$J�=ƟS/p�vm3�]���B�.�c#��%@Zv ���єa;��N;��+E��+���25���Z��*���I��D���>�����?�UH��etS�!�27�)�9�b��*ԭ���lF�����X�sT<���t�]�1��j�@�UxT�Ψ5Y��n	�ʮU�^��O�#�`�����>��7�]�{dς^��V�Ϯ6%Ө� B󉣢.��X�ܦ�^��vjߺ��3|�/�x��*}�,˜m߀�xzg��%�l��?fT��Lq*Y=��d��Kn/Ț��a�Px��,�x���/�~��;���2�!�=2G�%���mԋ�W�G#*j.��n�$�QW�:�������a��_L�=����b��}j�����ݹ8�!Wo�G+�f��w��aY쪣�Td1ckҲ'������Yl�G��Y�u~��~���[����-�]�j��Wz#������Vx~6��?�Ńѫg/��9q�3}�[����`�c��n�����8����9g�?U�q7�F�*�t �����_��O���Q~`~����E�[Ş�h>�&wv���D{��6=����$���ӷ\.XDT=��FT��ܛ^`�Rj�C�ƷpZ�ڻ��v���p�lS'�.��7���잭�<��HO�?_�Zu�*҃����֎Y��
x�$�䫑5�q`�g���ݮv���<&��[�	�S��}N\��|��\�ri�覔�R?�P��9 IT0\.,�7�X����['ٓc���s]/z�{o���S�;�f�Gn��0^"��/ܴ��*��Hڅ��V2S�c>�^d=#���z��ݽ�yV��N�Y�a�7��V��,aq�X� ���<N]�^��{�^�{=y7���	�|z��.��P�ƪZ3kE_j^�qV��з³��#��@�j�9���K°�l9�g,�o�֦�+��=8�_�y����'�ٺ��c�][qﾰ���\�\�ʀa��Q�]Ƅ�^u��Y���.��{ޑg�y������׳Ӱ=�=%����z�ht�+�C�Be�� @^�c�϶�xS�8`ۧ;��}*k̅ޏ����L�~x�~��=���`?z�g��@z�ĉHy�F��jE�^���=^�w|$N�X�:��G�3��.j�aD?zԏG��3�R�fo�v�W>��u�%�^�:|*���n���ۯ1�%L�����ݏk��(c��d�}X��4O�$��*��0v�\C�AU�6���Vˠ�l�M�S����{߳��'z�,�f��ݍO?f؊l�|J�p�U«Xuը�W������D"�G-�=��
*�rtb�2-�Eb~��+�.Y�'^ATU�k�T��U.ѹǙ��#����*ʛp�;�,Ee�X��{Y:��8>���-\�G}��#��Ė�Ǯ�5Nswf��1���f�=��/`���;P�D�������>;�x@>����xϩ%=s��&���g�+����h�dԯeV��ݐ*�w}{~"���
��o�Ԟ~Tg{�G%ff}�Y��w�>�ּǝ�'���N����P�]C�w�_��=��x�h:[��~����C�bz��ަ��;�C�Q���;R�ٝ#(u��;���w�k�d����OD�Q���,'� k��}^0|z=��[�Yݞ�ș�t���QҮ�S�.���0� �W��MQ�n��Pm�ӥޫ��=~���pj)A��uw��V�t{�����>�yȲ�
B��p)�ԏ ��+��TÇ��n�ZezQ����9�v��/=s��c����\�_�ǹD
�y9A> .�S��K�S�j�t��F���g�z3���sU����79K�Ν�{��.���Ϸ֤p�n���.��+�C��i|,�b�ez��+��(�0=�:������C>Y=�e�x���� do�b{=v�Ղ��4cb}+8���rݨ��L���P�X�gs{x4�kk!N��/��k��rp{�An�Լ�k'*�EӺx��&�J�����r���Z��X�b���r�t2��#������	
�u�[MT��=k���˯3��F��mf��w�'uvo? %�ď�]�Ey�\2!�7�6'��������{�����c}�����X�A�PϠ]$2�5O֦�e��!�8�Sps��z�C�y�-"�z�rn-��W9�Nq��ܼ� 3үfX�US���^�W�>=��{�V�ƽb}�<�ߍ�d1���<�k�b=	/`���W�O��a�@/�`�v����h�����ߣ�߈��0�}6=����{���N��fʖ�wr��*���^���G���eT��^F�g�k�B��)*�{�S|1a8s���זצ����y�AY�2z��)�x�C>��9�Dg��y9v�w�R�7'��7Y5�;������9Hx5q콿!4����{z]U{�T���yם�V��ΐ"��*��fZ�>�j�+W��!HѾ���c��Uh�x'C������ݯ��W��R����ؽ�Oi\�h�����ж���p슧;s3�ة��='�;3Ļ9��J�h��ϩ���q� <��z;-0wز	�w�F����Y�;r(�8r����m��YG�=�M����W<@�� �w�g4M�SsiS�u14*#;�[��9��-�K&��,�mڱ�c�ۭp����8ns�����s���=�gb�R��)5�id���S�M�Qmr뱮j���k�U��Q��x+y�[J�8�9�|6�ZO������n=~�~�x�S�"Ȏ�v�� �P�.+r2�#����&0�z<ʢi���^�{�U�.a���g�ފ��w�e���|=YFVNPB�`��x�d�êU�o���i[�؟@�\<�1���ȯ�x�VE7���>tv;�2��*��v�g�e�g����P;��Z&g��AL�Kw�E65s�+~Y��bBX��?T�9�\�]Ò���>9��T���ʫ��%r�E�QԌ�uiW�{��8�A�%�O�؅�>�
7¯]�i�}��ޏ]�d{����
�uA�ȁu�%yUάv�1^�y�z|w����=\���F�xJ$ۗ>�{����k���bm۸�T�75P��GD\S7�=��PS�ݯ�)B��J��_��y<�ȏyf\���y�O��'�/#fn�*B�*Y#�mg�L�|�p�p&r����|:Ǽ:���_�=;󼱐��2�>~�L�헷��}�R	�+�'�/'`�s��VaA�I���ul��}�;+�y*���܇����}s>�[�m�!�?��{M�F��r?�Ԥ� x��r�Y��[�^~ޘ}/�|��Ş��^SmU�Y�ssw�e�s��g:��}V���y�¦:y��G9X���e�����Z_�J���u�Z&6���e��vqWGP���*uB�8jU��Y�u]��&{*��:�,m9Y���/o��-��4�24������"zyL� ߻��P����7K?W�>�*���ȗ���b��ճ�����龻v��~�w�A\Iؙ�1��d�!]��G{,���绫8A�m�2����EW��_��O�����u,�^���*��d�}&�;�/
����zFǲ߁ߞZ�F��7v�F�@�z���\��Q�o<w<\���A�,�e�X�g�bO�&���N�����O���'�n�zm�2��\���Gc*��w����^�$�
���9W��4�.�O��=ީ��o��yW�ק�(G%��tl�v�|��J��OD��td @S9��p��7^��U��g�&�y���>v|��cޟ=ֻu(�Ӟ�;�oX����U��?:O0\���M�:�Y������ё�i��3��,�+9ݵ�/=s����:�x����W!�nW*a�/��ݲ�����$�bιܬ~�e�N3=�9S���������~�@�����늶(1p��p��ΉFp��'?e1����W�=��Ҏ{4o{9�m�-�{��k�:fº��v�AHx��K)HX�z�������l�+�N�,�\�N��wyV�0���N]l�;z��2�"o۷��[z�E۸��3��_e�z�.�����Y�����:b�n`^�?x�ղ;�y]���\��g��;޴�'ղ���_L����R��_`��#������,���U��(	�s�c>Y^��'!�d{�\�����?zԏG��3�Q.�g��{�u���K�(�U��W�x2BP����o>ܵ�llBT�/�q�]�k�P�\��Tt�̪�o^z���g���̜c�T.C
�C����t��;�M�dyp���JWo��>�t-<$=���c>�S�8��� �h�G�W�GWK��&�p�=������������͟N�ߖ�>�>����h��{,w�7��k�exk�Y��X-{�૿x�.w�dxZ�#��s�3}�g�a���t?Z�~us�	�3�ʩ�T����yp=�(��N��_��x/\<�۾Ax~��L��k�S�){�7�q�֯;R�Q���.����N��Y��q����S.v��ê�c̱�K����t�(5���|NC��#o���w��
������W\���V�	9u�%�󠖏kK��8�i�C>���G��*��U\�1���wx<\�Ɠ�{���X��6��ԫ+T��t����3�D��J������9���&���JC����g���7�&�9��.���������3�)�Ց�0q��n1��J�C3;�E��҂=��h`.fpЉv��9�:�7��<W�����K�z�ǹ
�/��C1Аn9��A����v銦�C^���B����<b��w~3~�'��.=n{�R�(���"�!��( ���)�Ao�S��J<�fJλ���Ŏm�S��5�k.)c�i������+�^`��tw�7֤p�n����O��l�z����Ǽ�徎�@�_��<ǵ1pPϙ�ȱ�,R�o���2@��z�����J �S�'F�Ww{{��U�
�LΪ��yّ�SC��\1�7>O��؁��=���}#�K�o���H��{?&���IX�N)��"}�Qk��D*^��9��h<�?�SprY�"�c�o=���p�巀`�U�G�&yպ���A�V*�{>�W�qN���}��z��lF����1y��Y�V��BK2�&�b����'��6�5��� �ӵ�״E�5���櫻^ﶗkGM��5~�]�K�߳.q��]�C�zf��l��A��H�^\�C;'O[O����������c�Dyw�g����N�w��O��u�����\��_KiwY�뫑�$�y��:ҋ��ڽ+�`�5��Y�`�J�E��^��]���-�H�k��y=R�9k�,b������V��sh������.F���d4TNgN�d=�	�6�v&���S1\�A��&)-�v[��%-Wx�ŋNw�;tt���Xꎾ�:Bji��d����k�qcZ�;Lc[}��	��O�(��T�+�&Y{yO�Ӱ�_yz��qG��{��f4�U�f��5δXR���փҬ�����[������� ����Ա]���H�\nR�uy��b�M^��-5&�F�gm4U3u�H,e��.�~a�m�[��Ru�hj�H��N�$�lvA�{O�[��+iA3�ˊ�P
ݖ0�H���=*��͹�|ԉ뱘����*v�\_ݓe�ɒ��L*�>ַt����馂�d�Fj)���tSs��E����4��rj�8u��5��l�z�ZMq�b�e�G�M���m�8 �������|�w͡	n�'m�uw��md�[��bJ�;���Yg
o�Y�uu���h7��s�Q�I�=�[��V�Ȳ�{^�ZDyC�4��J���=�	s9|��L����I�C!\;S�eGK��Q��ҙ:��K�Tu��=]��Β嶖�kL�u�D-Ȗl�v�S�44�u��fh�zfB���E��)]*��aVTZ�1�����s���6��7���w�v��C�uj�	�J��Py���xX�p�ڝJNto%�� �L�\̓z��f.���_gp֪�ؔnbf̘���R��gh9���r�sF^;�(Ŋ���rioWd�J;��t+8�5�n��Vq��5�3����7w�t�(+'QoCcE�����\�5��ΘyJ� st(�9�tԞRg�e�ES�D�v��n�}{Q�Y��X����hx/$�x���k<�5ca;^���R�C(ީ��DwWJ�\�vS�xF터��ocJ�m��Qb�@;O]�-;X�>G%�ɜ1�m�V��L���Wj��ç�����ne���-���v�8��T\�'37�'�B.�j��Fed�֝�1۰d�v��oB��"�w���渒��ٴ-�vⴐ�ķԺ�A�e][^���8+�@�r�V��b	Ϋ1���3���g1�ga�S����ʡ�|9ۙVٹ��lm�m�����OS;r�o������c:��5$�4^�Xk�]i�S�ٷW{�ǰ��d�����e.v�=��LZ^��:��`of�ǲ"���njpLY��@hÛ�fuF�a3.u��Ү���̷qc��!yB���vxJX��[tq��;B]ϻ��ݖ�v�mJ!�Q��\� ����t��������t
�%�B�1\^gj�;n������zH����aPj�V�;�N��W3�ds�<ػ�X�*�T	a�*.&躕gJ �&^QQ����9Ы����%I�"�ηZ�I""��7%�.�ZEd�QI�u8y���^��abȯ3ّ¢�/Ν�:���Ù�A�r����.'ZY!A�'Q�ADV��EEB*9I'�\G2T���R��5I,R�1"(�\u"�-���7EФ�"V�\̊&U�%6���LZ��΄U�]�t��ZDS�g�����K��99��:QEPz�t�.sV�%e�벣�2=kI.�T���*�\��dgNI�Sn뇙T)arQhii��D��L��d����Td����I%�KK�E*ʤ�u6]ĮG�QT��Q�T�9M�q�*�dQr�/$�'v%`TDNB��T��T�52i�XWM��󬈨�JR��!�EB �a��%߫g��E�ƭ�Yn�W�vֺ\6���t9�wgk3N�PX�.�Yӝ8�ڈV�]��D^�u����:c���9W����@�5��"��5~��Y��ww����^WQ[8�������K�bV=��2�z); -�K�۲&��N������ݯ&g�H���]�����>2�;c=�-F��B�%՟֖	ߑÑ/uA-��	E��ܰ��k����n#�yt���:��y#�.���l{-�x�	�z�iʮY��Ȣ�˿X�`��NF�U��ϣf��B��M䮟W�N8�9��}�{-O���"��B�|*�W�w��{wr�Jsz�G���n�l-ۊ�<{�P���c����\�9���lEeY#�]~��O&ۏ/���[|�Y%~������ٻ��Q~�Ȭ���5z�Ύ��e���bz����=�ٽF{��ST��������3+�'�9-ߤ��f�Jo�"�+�Ć�[����������-���}��{���Hb�@��	Ȧ��2��LQCV�dT�{�T:*�C;G�Ň�n�"<��@�w�����
� j�]CylH��W*��{���0��ذ_����i.���P���DޏΜ6�Y,�;��S�	��1��L|�W�0�T
]�\9z�C��ĕ^%�Z���>��ul��|8B�k�C�3�o�e]gp�w����Z��I�X�eK�.�Gfo	I^��őK��=�(%�.*��Y7�EZF�%�~s��#�N|��K��{���V�Ϯ6&�v�*�T�0/l�����%Iv�y�<(�UyX��L��V��N��}�wr��������ļ����ʑj���<�ў�D��weV��R��^��ہλGvR`���!��_�=;�;���2�!�=2G�^�K�_�^�G���*��Ԯ��#�\�$�ᒺ�}ì2<B���z��Oوo���}j���=V��w˽���-u�
�R��ܜ���ZC���rT�t����|�� �!�8Ӌ#�齨��ʙ������>�xďf��G/Za�]�r�{���+B]�^����歜����A���ҽo3��{]�*����F�;�����G{,����I�7�E�o��D ���P��k�9�LTL�9��V��:�]�@�s,�W�N��§a��zFǲ��u�$k�3iۮU��
�]0���S)�*0�~���)�,��y�2z�[ؓ�ɇ����9�{�{�~�-�b�Iج�.�z���R��r~��e S
WώU���4�.���_�l}ީ��lw�=�W���3��ɭu��W�N�D���M
%,�Cկ���[y�:�h�w!��c3r��g�d�A�A�{RعXX�[�,[���O��̋�x�[��n����l�.
�ms)�'S��oV�t�6d�3���m-���,N:��pY|z�zܸ�UXF<go�dJΝ$�g�����Ֆ����^��ǕC0r���=˯�g�&�#F9}�����<W�t�c�ީ@�F��Ί�D�)�	?<����\��ީ�\}�u�)��Cƅ�V\Ƕ+�����u��f�K��N�}�hw��<F����lCȉ�Z�2��=bj(6hL��_�Nx�>CQ��M��\�t��̙�S/:�����27��3�늸b�L����&r�moaT��-|z����E\�s|pOKO���޴�}[,~���{=�X���d}���h�~��D��bX�R6�+�	d?>b��ͬ��~����}~�����Q�7�}Qa�-V�bk����+�P�t@3b��(d�����nZ�66>J�_�#��̰r���i�^���KN�cx&�y�˹��{j���X�rr}[/.����s�{��O2�߃+�[�U���т��BK1�g�~��{��~��g�+|G�Q����n�å��)�|�}��]w��r/�@�Cw�y�6};�w屬��z�y^M������������b����i�Ῠ�s�f��� 3�X��06.d�m������|n����u�-�NQ��i*�K)��L�v��k�og�<�v��x����F��>�g���)+�L���]��&�a;o��Q妮����i.��M4�5�4A1*Km�m�@�����{�;�~��@�_H���37�垝����?Q�N<�$��v�ﲪsM��+��έ����<��r#�{��q�۾.���O[��M{*S�^�]F���FM��H��a��8�{��"�����h{"2�{>����F�d�e�9N'�l^�������Q��S�)m�ύ�ho�9k�o�r={Jb���� �Y�~����߮�;�u���Xk=��~˥��^�G93Z�E�d��,	���{G��+��\d� 뢼�	[G��H���h{���Ƽu�SSU�#�:�o>o��3���s��z像�#�`VxCȜ�����
�9���)L��ҧF�=�K�o���N�|��u��\W��g���}M�:v�����#}jG�n��NPa*�ҵ�y��Jk�$����xT9��@l=P��C�ȼ�+�Z�`=� {��2@��z��!k�?��늫��H�����kЪ�ձ3-ՇBj�� �h{S��7�66�H��;�����BV��C]�3|�z5{:g=Y�L .� А�Jm]4:y!O�<T��n�w���3��߱+"��:!jV�l��mFckMIk��V��	P�{w�Vq��d�vp���2��-ld��i*��֪�gv�V<L�lvή��o)y�e��J=��{K5kJ���|
V�5�oL"�|�s�.f{�FW#��Ӵܾ�� W,�۳��μ�}�<�/�V�lK���V�T�k�P�
�C��F�E��U�ԅ�[�v��(���G�Jl�؄��C��z$�Fq�`�/�4C=5���;�j+�+����� _=�,����7�8^f˖�wr�z��c�zf�G������H�5�����m?_��n5kѫ�4Ї�_��b��]�Y�2z��&�����Ϻ�k����iߊ���Q�l��µT�C�D����Ƚ�!���7�i�dA�Y��ww�ꮇ��A]�P���9����w4Uh������V�܃^�ð=���j����oé��j���ٷl�k�{ظ�(����]�w�~y	j�"�{j�r�p숪s�5FVE׬t���ϕrW5��٩��-g�c���炙=#<��zF�-�x�	�w�F����Y���H��>^�U~̌|n75�D��}�<�ܠ���Z�����q�������z�O�E����!� ���s8�����ҳ���º��ݗj�,ʊe�ܘ{��t�z+���g�ψ��2�p�xNa&=�IT�"
�C�gNw�`WCȫ�:����cI�钷(��9�ڌ'�W1c�}
I�֖(NԢ�I�6��4tydϘmk�S�#^���{�pm�Clwcme��"��o@��n���ٕ��E^o�N��Į�yn����e�����asd��Ϳ
< �D
�P��l4�dW�_�r+>������8�\�!A�EГO��]7�~Sw���������a?�܀��3_Kw���z��6-�dV}^�$0VV��>�]�Fן����Xlx��}���?�T�/�PW^�5Mّ�O��sPӹ9@��3m��vi�x�`{(#m�����=]�c��g޻�I���l*��6Q��sD�����]ᾪ��t�*ix��B���NBk=.g�V<@�k�O�6%Ө��S ��鎦�c�)e�Z^������c,s�iK��O�s�yf\�6��{~�W�O�>���/�u#��{=o/�b��;5ǽڊ�*�@w�EO1���F�GvW�7�����>�y�X�޹�x���#�-��w�뺫>�W�U�R�*� �>�># ul��v����C��dd��z����R������Gi�u�}Zr����nN!�܃^����+'���E��{[ �q��^�z�(��F����>�I,������������Y�G?^�s����~8�%�VF#`�?��#�w8V� ��!�畃xt9{�zF�8^�D,��]��,>a��v��Wݓ�7%;�P�ۚ/9t�SG��=�Qֻs-�ap��u����G�>y��5p���;�U�"�r�9m�R���+��)BM
����d�7jf��cӮ�{}#��X[גN�oH��UpR��B��ދ.�-H�n�S�����3LW	�S,�ҙ�jx�*w�x�����x���������v�,�'��{:�s�6t�U{ ��
���+��e�n�[R}�0����u��W{)�>�ي}%Ǣ��7>c+��YD��O,��`�8	hz+��r���4��^d3>�hQީ��F��/��端+�u�4�彳��Y?e�q�7Z]�i:���ډ�&A��<�9v�zz�׆G�דw��l�c_�|z���.1y��H�Gz����YȾ]�YMS��<L�._�lj������yQ~緻��'99^�����~�;)���>���dz�q`0�fR�P��.*����B7=���>����N��u�����b�;�<s�=�='�~�@��{ p�_�*�6v��w�����xW�8���9���TQv�a����2�I�O��z�ߧղ��~��˄��=�j�/�(�U��j�T��-����x߬b�h�K!�d1p[W�
�jG������[P"�����/e��n����6�pF�d��+B�hM��/r�Z쓋Y"��u��Mg=Wi {j]��
ޕNU�i�+�� x�}wQ�EL2���bgv��Է�j�b�>�Ϋwo1y�������Ž�����ǋ�=������s���)�/�����0]/m���/�R�F����=^�}�+�����v�X�T����̟lK���#�H��^<������k���=��k����>����\�׫G�盐��bϢ�aǺ��ȇ����Z0� ��چ����`��8��ut�?5[z��ʿj>���~�n}�{3gөߖ��>�^��W5˵^�~9�;�	y!S�%��蕀k(����>���^�#���㙛���N��a��^|�$��v��Q:�y���Um���}���^�^4���Q�����|2��g��Φ��*R��o�㙡�`f� ��3������k��~���t��ݕ�=�OD�P����~9N'�l^��=~ϧp\k���۾�=��C�a���&��Y�ޚ�6� �R�\�xr��Q�w4蕱��i��> �s�����������6��~�<��\BE!��H6)�ԏ �٘c�y�Ͻ�������Nn���ݺ!_����zL��}�=ީc�����/D�- �?-%oG�'z�����������0��o�)���b���FҰt:�G �<���i�<����;���2ŀ|2�×�`�o�0�Q�@�.�S[���7���)��H�f�c�V�SeU���["�M].m�<CQ#��2��2"��J�lϢG��NGUy�����d{=�nr)�gJ�ט/��7֤p�v��
<v�捕�[Ư��|Dĥp*�����j�����(d3�y�{�T������q䝾�Y�������xN���ު
���:�9Mّ�E4=�\2Spq?c`ߊ�o�f�r/63��r{d�f{p=v�G��gL�G�<*�P	�ؒ��3n[@��)�;�� {1ǆ{n�V��j���Y��W���o��˽�~O� ���tR��;�yo��w��?(�>�]f���
hx�~�dg�z��=�b2~�C>���'�.�lװP� ƈe&�E	�����vRS+��z#�R�Ξ�W�Z�6�w��]��!��]����q��zrO��G�L���ܞa�qk0����j�w&���Y^#˾���g"f�S���>��9�Duk�2��.��.���yم]ה��u:ǀޑ����p������p�i�diŞ�U^�U��a�fdW�m�пF�^�yq]��w��,���dy��d�nw�߇S�1�ļ<�U���u�+�����/��;%j/��a9�����Ic�1-�@�sݔ5Rx�e^2}����-���u*k�_>z:K�.|rm)aɱuɤ�D�Z�ˆvp�Yoq�Ӛ�Y[;�WVc�f�`ۅ�-��R���w8~����u��$���Ul��89 F.�c�W��@�>�������WsQӻ�*��3/"{����H����A;�B/N�p�,�Nw%s9b���e�)M����s�Yv�+u>D�^K�����q����_�ǲ���
�"�ۤ7��� g����x�FN�| �@�(H�)ӗ~�[v�Cǹ0����{�^���\�9���J>�˳��.[�x�n�Ү�Sމ�[��C��W[���W����EdE7���>tZ����&�N�>���/��H���=`i:I?:�f����2��ߙ���ſ,���Hz��c�q볾7��= ��2:=�}���lSC
���NE7fFA��*'�f��#ەD��~����OR���Kζ����2��;#�~7�5Y�ȓbU糲l���wg�y=y~I�ʽ��z�O�<V	9	�������լ�Ȟ�n�rj>�͇~W��;�Z��z3\���Ռ��h���\:��h��U&�u�p���D�����6����`����`����6����1��S`���;`����6��1�m����m��cl����cm�cl�[`���cl����cm�m�o�1�m����1��6������6��m�o�����)��������9,�������_���0�^�=�R�X��U$�T�*(����J��HBR*�
��� �"� �	U��D��" �n�j��*B�B�%5�UBR%�!TR�)�(�R�@����TP��TU@qh��*K�R����H�"�Ғ4���QI�A�)(��*�P
�B�E%I���"���A����6�Q�a���R��jmj�D Si��)f,+P�[kj� ��m45"iUR	 P���yI  ���֐њ` 3�QFR�R�Q�1ҁJ�q�� P(n�qJ)@��˸����T�%+��(T�-5�(���@��)�KMR�̳��@t�M4;��T�;��hle$j�n�d���R���4lD�	$J�TN�  �*��Szt8��t4�ڧv�IՇs��;9�iݣ�[�;uN�UU��uWZ�N�U�H��"RRT7�  ���5�kkX�:%WfV[��J����mU��p�5[m��k��UT�â��ɻ�R��ml;�U֭��0��j����*J�%P�� �{�҃����\�U*��tu�mv��[kHvR�T�p�5bڭY�T6j�6f��Y02TQ��M��U�MP )J���Q�=j�mP�����ֲj���X�U���lR�j��mf�b��UEF��ѥ��S�T�kZ�%JJ�"J�l碔P����m����j��)��%BD�B
�3j����BY)e�UR*��Z��b���U�,m��U�5UIJT�YURKǪ�����������Z��Y�A-Q6ZZ�Jڂ�6�`�j�MCj�F���Z4�mZ�E6�&��6�)J��hTJ�D�� �P�5���m�@���-VP
@�a&�h 6����Ɋ6�k�	 	  (  ��eIJP�# �4`h� �E=�	)J��hC@ р&�� 
�� OB`�@�z�����M�S�=H5O��JQ���`�# db`C Jy*��J�    0��  M(�1J�� h�0C� �&��?������4u�������{Υ�)gw��}�����e~)	5�g�a<�	�~�%�F"uD���������$@L�J�����W��
�����OV_�Ŧ?\�qG֣��"�QR8BRYCy���YB�Z�4�HlJ�:E�*H"Iԍ<=��;�ËF�u&e>���^�_N�1��{ޯ{^���}���m��m���m��m���pe��e$ ed�,��Q$��A���)"��I��Hb��b�b�((I2� e� �I��I��(ZD��b�!z�!���$�H��1DRD��I1R 2�!���RC,	$�A`Db�F)b�*D�	&)!&Y L�!2���		�H�$�)!"�d$�`Ha �D�!1D#	P�� ��BL!$�d�IP�L���1H�#��I*N8����Y�m����m����m����m��lm��m��l�m��m�6�m��mgm��m���m�/���%��Y�cn��V�(�k%�e�T����[_:N}-W.�RUm�<��Z�}v�J�������Z2&͂Y�w�@];�	e_��8��h�{�q��]�Y��͠��C�-��"�M���a���30���-�J,�61���8p-{shl��m� ޝʊT/J̧)7L)-
��d�,h�{2�H�0�f9)ǘ��.���5桶�i;S1�F�T�5�$�.&(�7r�7s���=6�L��f�sg�X��{��	�z��RT�ab8]�ģ_d���ul�)H�Xw�u6����T/鐣L���R�ޅ ����6ɚ�;����
�ȳ�,�����:����J�����_;R�V�4�:�鹄@j���p�� y�-
K���/,;� ����LT���:v�,���j�_S&�l���u#�7�r��7T���l���I*���zkl��ToT1��jj�j��nQi�)[v��[W�f��ԢR�Y,�d�c0�lm��n=D݅�)E�߹̤*�����P^Z��U�S%��wZ�Z�y��p,�re���7h�(�`Xdcm�j���:"��K�O��(�;Q
�2�_p�ϊ�3]UDj�UU���u�rٰ�%�x ��y�AOi1[��ؑ���[���F��t[B���p:��f�;w0�Q�i������k%^�v�o>Y�!ȭ�+,�n��v%ҹc�E�x�ٗ	�e�l�Ma��v�&��B�*��dl��23,�)n�*�{�^���:F:�-?�<Yz+,e:X`ir�1��{���_Z�R8�E�k��9��CtR���*a���b�iH��A��s[ӛ�:�nV0#N�a܇h��K67d�6c��	B�,�Q(P�:��m��u�/j2�t茗sQ��a��a,���tH¬�,��Slb��6˄�/M�Ն�v+oma��.؁%�V�N�l�*�	Ie'2؋3][�P`k���Yu${��]+n'�lեj�$��V��m�b���f�F��m=����@�l8-G&T���2 �7����
V�b�'�f��w	4 ����8/-�5�4�.�!�:͇,9+1y��j����)�@KXq LV���ra��F�ݵi]�ۖֆUf5/�AƮ�ۺ��q����"�I�jT��z��̭�����-�q�hx��g)@5ɳ,6�hF���&P�~�yI-�9-Լ�&5u�J5XJ4���3C�יQ`�2��J6U����鮝;��CV��@�bm�hae�Sua���hX�'�Ud���eh�X�lڶ�t*nmen������Mю���B�{A1���Ynm滋u�4�F�mf��������M7�48���C�7
ií@v�<ώepS/vQ���o詹���-���b`��A�e�P�0���ś+Y4��gMD��敄���&�7Cw�aж�f�	Z���CeCz�)8�J�]\ݼT]��L�:l,�촴�&�C�am�3kv��O/F�eK���n@�8r[�Mݪ�%��-�yW;�];�cq�lK�'C.l!]��\4�*$�4o@X"R�t!��3ኁ���G����Z��w&�cvS5l��ㆆ�S
����"(㽺j��6���\��*�U�m�Ff�[�S��ec�&0j�Mku��;Z���w���ԝhT1*;����wKOŖr���`Tʢ���$P�Z����ckiI�V�Na�� ��k5�p���Է�dtE!T�A]emh,�mۓ.[z�dZ�c{�:����߈�[�"9vl�����fX��7E ��*�C����RxTKռ2���X՗*�Ed�W@��o��W����)^R�����1l%Eg0�Y�f̍f�v��r��
s^B��&�����-5"���T�b����T�@�7CNDh�Pe��M���H�#��x�KA�u�`WH��#�ԡN��`Z9�.j�Gle��^�T��ײ��%L�t�n]8�ڷ�g�C�-C�U#v��W1m]�yO6�ޞie�����H�x�[)��y�Lݷ��$S`
#td���\Os%��:�Y���%n���Y��p���"�
F����''If�/�)d6��/-�E�Ý��(`�3BYxb�E��!ݼ"�j�T�إ�v���H&3"u�m�gv^�,�C6Q4�^��baxcK*�5�eE�64���[�U����*��i�b��j�[�V��n��6&**��bt��Q�MK�����Z��-E�,2��)�v���^�M��E�!�v	��V���ǲ��ǵ)KؚMf:PR�H�Q�ղ�������
̇fFkoS��b!꣋��LT�N�.�'�n��(O�/j	��oI�wQ��q ZY`�pİ�T��\y[���E$)��++m�g0 Z��v��h�p�u�Y9�@�r3N�)5B�bDT��LM[��b=��Z���$�kwl�Ӷ�P�%eZvM�!$��ale5�
:�0"�DeU^�{�3�*�/p&[�Խ*km�`2��aś�-Zp��Ah;��j�8݂�����d���fkP�ͱ]�ҕ��\:�@�*f���h��t���+w	�Stf�ح!#̻�*<�y��{�$n�K��ȕ�2��Y��[�f�=2��{���D^v�5��Tkr��faV$��R�Mp�{6bO�����F�໲�5�&!���lf��VR1��j73[g�xPH(>�*�Zŋ'rX����E]5P��U����u��%Ƀ^�de����=��� �f(����R�;�m�����֘�)�;���PsBnK�	�[,��Z�Lp�S;����=űW�ڬWP�Z��Ie����J�܋7!�fS�H9����� �F0sBb:�r�e���f��z+mS�Z����Yn��&ޗ�$+u��-ݼE`P]��*�֧Ƞ��zH�4 ѳj�*f�0�ص�"�!Gv�ˤŀ�Ԃ��Gm	[��� �;�YwPdۏk4Ķ"�V�YZf��;��ؕ*�1��sab��P[l�1&��w/nd�]��5P��i�
����,X�7��·�sn*p�J�3UP7��,Zi�E�`R��K6%a ���D�[RY��6�dו2�v��=r�B��t�j)wz�f�*1�5y���5�������ucݽD��Ҽd�$��
j�D�3M�faK�v!Gg�;�Y4�Ę�KEc��V#V*�ej/]V�s*[��ӎ8rT�	W�qY2�V�s.�Q����ɴ��;VuQ܋"9㻫o2�
9�M���g咖QWu˻��D��
K���s��3i�{����!X*0��ra���11�YOPoZp:'Y��!���[��RiY��3Q�^i����A}��-�VXl��
���qҤo6�1�ӑ�ݬ$̆5Rb+Mj�g^����Rݖ����6aNզL�,IQ���åPu�|�l4-��n���j�MF��.���]�,�ν��Q�f�i��֪/l;�l���xq=l0�X�ɚunl��ڛ�aU�I7{h�d�!��.��fZ�V�tL�}�Y����ḛ���H*�. �6��f
7���K!\B���Kq̺rE��T�5a6�tMݸ)��s(���2����Q�xp ���e�t�k^]hi�H��.c���c(%[L�2��FM�Z7 �&�)�A�s�(��\Xv�`I8X(�b
�L�a݋,d�{1���f	�:Q�Rvƍ��y���sN3�X�#)	ʳ��N����v��8��cm�f�\ׁ���b���e"dB��e=k"'���t����E�Y�����.�&��L)5ֵ��r �"�kk6�J0�3R���Ӳ&bțǷ �Ձfj$Ù���v�����VobʏI"
4�/#h�+Z����{�n�n^+�c%�mMowdl��/)�;D��X������NYD�p�ۏSf���S7`����/�mA��l�)����OkB[�J�ۡ��G(�喢f�ӖfQ;&*{x�� �+qM��0$0K��734<��JAG7-�w*\�N�F-`��R�Bw�{FTK*�sD��f�d�V,�S#]�m�u�B�7f���H�Ż"͸�M���rMbUc-�X2��X����b��afˎ�����a�����"a��8� [�V�#�Fwh��r�ё����	�e���Ddy	Z.b.
S3-뼣�YQ^�f�dA�r����� �a���5�F�T����B)JB#""�v�[˄j�.�9yim�R�V��Z\7x.[gt�Μtb���̪��w��$�_,�U`��vt��vęV`�ǿEYP�]9�mf�V��+�a�n/j
��2��`��v5�J�](4�t��&�����j�i�u��f�9hL��a�yj�̰�����"�XR�V�C{+Kr�&@s~�@d!�c���#1�Ktm"
U�bPZ�R����ջ�n�6l�v)�N(�e"��Hi�i�K�e!d�7Gv��f���V��i�Qd`S6�.�z�{��M��2�����(�j&nh���.Қ��L�DƳ(Y"�6��W�ۅL�5�նv�;��˘B���+�D{[6�KwF	�4�b+�۳8IZ��Y��6Fس�����F�-F3��4�ʦ*U���,�`ō˟dI�L.G��Z5���;-K]�r�F*����S�bʅ3�Q���*'%�l�x��Y`��� j�x�fH�'�]�gh�X�(ڔх�>�Vj8sY�b<�r�&,�L�UBH��Gj-Z+�7��Դ�%<�$ti�ɕ�
E����k����[E]�h��M�r�(U��I��R�	�u0�ŗ�Ea2�0K����,2j5t�u���b���*`��ga�7��ED�fL��
�¥c�DL��"����0-��g^�'�ܙ@`H���Q�,��E�;�H��y�fT�m�ٶj�hV��P�h+1�H�v�����]4�`BP���{����#/���z.��մ�0ö/�X�,�����KE)�*��D���2�����Q�ېU��%+;��%�fؽʎ�^�2٘�Kr�lv49)GE-���($��e�ؑ5��]5����[�o�o+E]H��&�i��6B�ՙ/e��1�0^��=t�i<q[Sh�h�j�a<��d�vj�5̺��n��7F̳��0�YjCj��,���n��B�҈�h9Z��R�urXXaKv3,ٗ��ju�shѭ��o�20�ԳE,�(DM�.YW��ˏk1���6wq8qV�t���a�L,����(_�o��R��1�CvR"���-�w��52�e(%�,�Z�F9Xv?�*�1|��-eÌW���ҧ�"��B����eIE*K��$�7ڬ����KZ4�E�wm��姘�.[�q�o����q��k?���g��ڻy�q,�(�y�F���p��[U-%�ؿ���h&`����Ͱ�8 ���4plT�V��k��2�SU�vv$k�N��+\���:A��;6���l�L�UO],Rw2mBׯ�]�ՋIBﳰ���3�d;7�fZ[��{27L�O��Y�\mt��x6�H���
��&�X[�v��c��7m98��Ⳉ��K'f�]����8�\ܻ|����*fV;*�-�9�GmHL��17�vp�����4�l�{�c��%��ts�bt6�T�gH�%b��F�F
w'^��z�7	�n�����o<�e��1����a�5�Od��!���j��ZUn�YV\���2�%�l���7Ǚ�e�H>�5ޗpҸ�\t��'wN��Si��q�kK3N�V쾾�cnd=��ɅB�K[w}�خYG�����5U�֛)Y=�/���s6��Yy�u"���W�#�yw�'̱�%
��Mޱ���6�3���3�ٍ�N���a�Y7;��fM�����ɏ�M��uvI�ku���Q��a�u�+�uӻ1�q q��>K	�q[�3�p�"��7rM��q�F9�nsES�G'VW_�֦���q8s8�H�{
Ɲu�t�&��c��f<��3)�
Nq�%��{����V��@��*s�a�rɼ���f`�L�����j���v�.�"�Y�,�����/����؆L��ƺ���+��s�j��k��8�E��c���b��>f��V�_>��N�f���r��	��풆�!��NU��yy�L�	�=����_.�N&�ό�S�������,`��pwŭ�����׎�e�����V]�ǻ�[�[�8귤ɗ!�C}Ϭ��ϧ�����l��_E@T��a��ǕԗK��[w��j��<$�.n��t-���i�l�3Vm
�:42��F*�WXj��L����w\͝-)z��֏do�>��]��j�+.�澙'y�Q��A�^w��B{�!\o�l9��ԓ�}#��_d+#���-뭅�"w��։:d�Ò�N&Ew\ܣ����eDU�^��X�'e\hH�T�ġ%g]�-ծ�)��v�|�X��y��pT�/zm˺�x�.����;���V��y���r��3O�v���Q4½�s3u>W��w�D�'fwbI�_q9�,��5gsJb�->�;������/�\,�ҹ�>=n�g/LЍ#+Q��u[Nk���x\vA�.Uᠱ��f���}��Y�S�q��"p�7��ȺZ���D,_G��$�]�J�LřɁq�2P�d汓��],�z7�&".��omڰ\Z��K%�TIT� !G�mn������]���м�;
C6�dD$M�������J��np7V�����n�����VU�*�R�Y��HfGS�̮�:�
鍁wU��Fܢ���*�Ǆ�6�
5��9����#��r��+X:�lm�i89���ǞR{�ҳb���ɗ4��$8i����_ʍ^&��u5K�9.�e"�]aj�h�w��5�nwN��u�7��dY��wD2��)Т2�Ej$U	��s!G\��B2�$J+A����� �c�H��>�����yТQy�*%*4����yh[�§��#�צu�\Uج�y�&�w���7fJ��8#�=�
�Z�L�pַR��۴�뾥ғ�.q<�����n�nT�v��Yf`U�w+�gMV��tM��:Q�x��_.�hߔ*���,|(�MM���{�3��F��x�p(-Io]�
�)��]��������vZUlE徐��ۯ���3D�('6ݔ�>��n�
�*�,e���;��ǢȚka���ΑGX2�Nfvfm�wZop�agW(1�L �IR��õ����ƶ���d�i�p�:Q�Ij�ə�T�y��X�"�k�8j�>��]@H����$!�ϨQ��v�Յ^��3^N�٣����{$��5I�k�t����9!�҅���M4n��0�ͧZ��*K�����E�aУӌ�f�s3&@��c5�8r-�j��ڳ����U��>����e�Uv�ɓ�;��r+t�>K�l�am���B�[��b1�PZ,�UmZԱ�`���b�����Sw�;8�`�[�A�]oE��X���a���i�Z���̴�n1�!��Cf��ٽ�k�q�#��Yչc/�_k?q{*"�ǔ�.��Ӱ1|��G�s���s*��!sf�+t��Y��r��=���/l;v�J��r����=�j��0tw��5�h���q��[*E�GB	t<�F޴�o[��S�Ff�S4�B
:���Y�����%V���J�7�hm@�Ļ���F�Ɣ��ӳ���zz��$���F�Nޭ�z�E�X�d\�h��k�1&���0��h_w�jRǸ�CZM����캖
�-f���J��.g
��d෬���6x�W̊�pfVUY�o����Pcz���7�	�O@���=�҇��Z)r@��_th�����dJ��ޢ�d��L��GP�rm��Ź\@���t+)��Ru���Ӄ\	k��f��9 ��2R��X���4�d���6�7g�	K�:z�u�bf��wP�83!�s3eM�]i�{��q[em.M�4/6����-�Q�'�6;D�E�<�4���Zj�6�G^f��&!�k1n�1�m��q_SB�UF��-�V���=�^��;@��Jٍ�]ɪm̕�vIj�E^�>�A�}�5I�DI�(U^#f��V��VY*w(뺴��]ЋK�zy3�G���8�������]G o���4Q�N��l|4.��;���h*��m��Tq�D+1}RL�C���Ț���'*�˼�w�w�Ď��V�d;��/K�U�s#��ε���e832֩]�0��zJ�"=p�?G���;��5t�	���w$d�ճ���=�j̋ q��Y���H���YϜV�����3���2��	T��Vݔ��݉E�%�Z�n� ^*���1˹|']�:��%�g�3��3ʹOD�M{�s��kj��$�C����G-a�U���3%_7M�!��gu�'��|�8˗���;]b�$�O-����<��.'0�eJ:�Ҳ�sW�%���w����y0C.�b�lXN��۝4�5�ǹ�R�&��燵�eByR�<�u��ql�M�Y�4��X�[jX�Z�0�7�
����o�aO�Ȱ0P֭J20���ZBvY�s�i�r��
O&:�Ai�u��ؼ�]Ǜ��(a��œjG�K��ax�����c2��y���v걱w2=����񯔡�GT��gU��I�j�N<�F��OZ��ǰ�Cõ2��\���;l�R0�n�����������xc$��Xhc�ՑK,N�ͥΦ�{و�{�k��*��6���a�c̲9��)v��BnT��-�-�q��v
VVj=zrbK�w��g��%�S7f��g�5�G��好l[c�]�۠���J>�]�����1�m[!�%�W|�&����p�l:5�ۜ�co�_=[C4\ޢ@�ݬ8�oGK�ġ��[.:[V����G�æ��x���g2����y�=�A҈��t�B.�����:���*�a��>��%աi�����������#G��u��h뙹��C��n��\�E)�\�����fa�#NܖVhZE�Q���l��/�4�{lf!Zw6?�dy$�����Y�|��J�uw�'a�w�[�jr�e�Q�a\z��� -�+�֦�mm+�Z������r��3�F�;+$��b�U�:��R��R�]�H]c�Z�"rh�6f��JK��ݭ#���p�����1�j:w�1�Q%$坋�gq�y����^�f�1/F�4�c;��u�':��ݔ���r��ڴ�
A�/�L�sk�E֫�V��v���$+n@���Vd��f�X��j��4�3 �i�:�j�' ���bf�Z����#����i���1�1�涍ږ]wv�Fv�D��*,S����e�o[�w;�v`{n�501|P�%W��n�ˇpÂ�Qs��
���9��K9���n����f��������o۹�б�,��m1G3�bn�ť5��N��ٮ��z���X�Ae����1��y�+���!�������]੬�7d*�7c+��� ������:^���K�r��:۹])�2�G|�Ø���\Y���USa�FI��G,YK��ֹ��i��[ҍ`�lK�v3R�����G�sK�HU��Щ�Z
6�iޕpcD_;�N��8��i��Ҷ�j�۹oJ]}�����X�=��	��*������i×��'��/��#�[.�
�}�ۇm��eȴ�L�v%\1�tb!��:�A��;CM�^vA/�U��=}�4Q�B�%�z��(���.��ӅmNj�8�4�R��C�~��:~��,0����Di\��������,c��/10�;V0V�I6a�L�,p��6�C�#��d�+[����<�r���T��ؘ��C��le1�]�]؞�8���n�1����+/5�"�r�q�&�t��W9���:m[=�!��sj��q�6�����ơ�a�YH�=���m-��7�3*�]�$��N�un)�yV�����(�/x��xg]����l�՝�"]�r�Vص�(75��V�dU�S÷���l��"�]M{R_A]��(�����P=K0����UvE_v:��	G�����'����x��T��37�>�f.��*{g�l���t���pq�)�#ӡ�3�X 놵����+�(�RZU}��3��TJf�3/�vH5%�B]�7q�����8����6�O�1�nn@��;�$mOb�ŀޒ�-;�CBے��;�%^1����3{�N��$,��ty�WӢX;o*����k��K~���|���ᕯKSj��c��D�{��y)����Y�m�+Ut�7��=V�Ӣ��ICH�Hָ�����qۗ`�[�s2}E8A���F�X�R����S,��ǊtUb���g�z�h����Ƌ��&��rR����p=���K��������Lʜ�&J.[��u�on�oq���<���u��s��I1��Pִ扛�M��Yh�3��87�;j�8�/uqafm�B�IR����E������X	��B��k���N�8X�e�r��|WCEJ�Ѩ������{e\���]�ɭö9+A��nɢ�9�F	�0�}ݯVE�ÓW���X�ݔ���:P��rs�iL�;�bg`=>�oc9;M��z����ዔ#�H�f�G��ÍN��ݕʉ<1��+��e�� nIpsS����5�*�3���zv�W�<��;�kk��p�χɋ|H�H���궙��\�H �۟?,��I'b6�޲�<ѭe$HI#���*~��v��WG��%g��Y�����X�%LÜ9$�U�ڴ�mǙrٟ>���ոʹ��B0��HVʝ-uD�6�G{Nfuh�8�yS+�_-�I�voα�kk3�c�m��V02���[���}��Z�K'��[ͧ��V�X�HxOpƵ�WG5>�bv�=��)�E×]WJ�M��̓D�MQ���ˁ��.�],`B�-��]z��陴��x�V��	�p�y9�>�_�MR��Hw;\��d�H��j��C�W>Y�Js}�o����U�%t?m��졵6�6�_qT��S\�[�j���ܢ����e�BIM�0�_n^�ҙ���^^�e�Ye;Σ{݋�r��,�k�B��=%	��)X�6��pݺ\_gJ�R�t �3+�&�cA�Yܾ�̻�Q�Vre��1�p�й��ݷ�w�5��<��w$�����:k;(q�^<�YF.��Q�2��#̱���M��{�c��%U�<
=9{�:(����e��O��������<�'Gµ��$ êW=)v��Z��uV�j�S�zh)�|av���R��W)$�$�)%uUI$�$���I$�I%��OO=�&B��&\�TF+3�`���oQ��Y��DR��s�>�H�o��u�w%��X�-��ݝy���TE�O��.7]n�r����f�&#�U��M�n��Tv¸VoI��[��"؎�SX�z��J�i9nrη�ӏ[��:�i�����WXz1.��d=\�O4����o�tY�]�:�og،8����oWe�L���t�S��Y�����>��n�8+iA׷�J2<��$޳�o�EW���&�՜��ի����vv�ք=�[d���&�{�Y;Y�oT��#�@��5�U��q�����뢛O[SqI�H��@x=�^��"\���5�ݲk�3���ԟ\����wb�c#�U������n�S��r�'M�<eA�R��]���|���Z���`��w��q5�v�Eޤ��y�܃��l�W�*���-���jU��z�.� �m��t�}:���ld�.�2-���U��L�U�h˗��$�z&v"��vst�{.г�P�Cc�.��jL�8tծDfZɘ~��U�Ʈ��1�k3/M$�	$�I$��k2�I$�(I$�I$�#��֕�Λ�u<W.�h�n�$��W 7si��u��bS�-;BM�V���fv�Z)�fЭXE�Y(���6z�T���x�J�-�ł�`�f��i�]�m��Īr�y��]>�P �h��p�r�z{�V���8H����q�W6a��9m���w��B��e�wD�8��)G�`k�$���Ql'ܳ3t*����*��t���iȫ���V�v:V��c��p�����B�rG2i痹vrp��7~%A���5m���wkz�w�mu��*���,;�X$���P�7�;6�S��7�����t/�m�o6.|�K;�&����PA)�XwC28Wv�vL�+�#e�ilc�ٜ�b�Qfw��ޮ����ȵl7+br{r�t�}b]&ᚁ͟u��d�3�r���iYf!\͞�p�q��wW:�<o�����!��ڤ�y�������N�8C6�un���-n���"k�Vv�t�����j�)Qk�����!T��+��P6v�Zr���o�����I$���V�I]��I$�J]�ϻ��f��wA�tw��b$�� -�t�1���vM]�.�L�STx�ط'9ܦ�N.����:<eWE��']W�����Gr�9%�F[T:W!۴m��83��\��ڵ��c�W\�;�n1X�.S���ۜ�����e�yjcV�}˟vJ&�j���&��o.ĸ�/��Je��(B.�͔y(%��na%���]�)J7�)��6�g�r��"��dM$\ʂi{�\�LH��ϗbZ���u�m:<�I��ܩ�S��Cr�j��:4�����'�X�
�LA���kl�C[ɣ��s_*�>%m�c�Z����q���N#8V�w���Fi����հ�!�N>%p�M�.�5�dd�1�k��.��{\67�6U��޾΢��<I���wIi/zq�#/���������ԯ��"�-Z��i�����lqR��eA�ݓu\ے��mmI;6@Q��B�	�n��[��q (nZۧ��t�ҳ�]X3�
n`���db�T Or�����ifb:�I.I$�\�I%wwv�I$��IbJRI-\��1��[ỹfbUv:�������y�wc�x�"a�i=+��m���1�Z��Ű7X���bL�¨1�(��Sa��i��J����&�;�֘,���,���F�*�|.��]k��8�	2���k�QL�eiu��(��/g��Զ�)�ZJ3�f��X�U�7_�god�u�3�5tM�]nq�s�^[Ҹ���oit����H�N	Kh�|k�)R��n�̆n��%��1��`���Sy�|�g^�1�|G5�8}{]-s�]9����l�ʳ3�ǅ��/�r!|v@�t�uэ���q!�3qnҗHp��n�.<�@�?��j.�K�U#�G]ɛ�^v�л��U1:.Cl5i`i��غ�=X9w5�2��̬O+B�C����BA�$ ��)���Y����=Q��ngJI�����u�ệK�T�{�pukvV����W)� ��O��#��9���u��3���"�;ْ����,�)�������hAo��U��6{-���N�
:��hn�ݱ�����7���R��f����djʹ-u���T�����=�
�邮C\�{պ��[.����9Lj��"l���Ws����o�Y�w�l�1�>��)�W��N�
�EF�vf.�C#]�C`r�
�5��˖�y�푯V*bk3�"��R��A�ŵ�x�n��k��ǲ�wv\�_k�Rd+�E�mרlއs6v�6*w%����)Q�7�+	��.L��#I�åU�U���*H���W>`���Z7V0�v9�w����>,�Gt�c�lF+ښVT�+@AB�+2��k��N�#�{����f�>�Ĩ�p�LEnoP��)���j�N�/����I�'S�ʓ�4�pnR���D����a2�1j�B0�L�ZR�8�:$��QЅ��r��S�D^AEQ{��ÚO��j�\�в�M]n��TBKguS��\�Ƀ��x)�,>WU��!z�R�4���[i8@�jŜ�7-�Ved�!&�r�\k�(���VO�������������{g&}��ssi��Ѵ�ua�Ƅ�\�L���(�����Su�C5c��q�KO�d��N��f]�99�5��ŷE����
�1y��>�j,�w(b�9j�1q)�C�y�4J8q��r��f�*�2�&�h�k��@���\�\�@��;oQ�M��G�����e]�x�䎺�K��}VI�:�(��9Q�xwUrҥ:�9��Ϻ.\���C��>�d̺��;z��XM�t�&E�+Q=��Ś�$�US�W�KM��[�{���]�dY�+��XZ(��Y���s]�4]j�!0��Z7�9텴�q��2��v7�B_M-��q���˺�DI��Tw_���5.�ҋ5���,;�_F�u�Λ(����F������V��N�Ò��AHN�eIi�49B�r��Mە��)�rڃS��p����$2��t 8�j]ݩXeu��G����f	,�\f�u�)��q�w�#��J�A�z�lk'�y��mc�.����Y�o�Rm$�K�j���}k\Sf.�λ[��=u8��VH:��z��i��9J��F�b���_bw!�,�ɑ���3Vǖ�s{*	��W)�Pv�W�sruM�c�P��u��Z��C��o�k�/���xc9��T@]I�-d(����.4T�v��5�b�.���U۽9�&cjs6n��1}�O3A��Y1QݝW��2��{�DF�V��.[x�X)
ۚ�tn�P�w[!�,����K�{,.��tvfw�ݱ�fqzksN�	�Sε>}l�d�P+�؇4��c.��L�pru�e�j��'�]/��T�eS��c<b����oL\���J�-+yFb�6�a8�v���l�z���Sx+)t��l�Ε��W]�pC���:�.�uo,b����O6���Qw��p��Wc��S8l������%ے�7��*�����Z27B�v�+ѷ�9��]���Y���Z0K��B�r��I�5I��b�X/nd�7y��w8�ہ�C!���ii-�zŖ�+!���l;ۼ��[Ϥ��da���#��nR�w��M����q�V
�zm���Q�8�=��G"&|��L=��t �X���n�Q7tb�=������nYF��@���W]l�x!h���M�;Wq�4Ό'��8`��ٚ4P��]��|���a^�C
XZ��V���"���]��Y�C6��Sn�uw*��A��t�N�DκDQu9AQ�)��Wj�� ���g�J��5�aS�x�]�@xNͭ�Eͫ��sֹS
u�ͨw
[���*�b�:��y�&��R+.���R�o]�5d9E�*B;!�;�p[�(k����]a�7�G���{��]u���<w#�h��m�s3��J��Se�yj��yB�vq���g
S�f��}�a$��cc ��vV��fж�Ŏ�=�E�D�E�Rme��uS�QW	��*�&p���!V��r���X���.wQA}V�z/�Ru��ӌ�50���Ѽ��Q�O���uT"�jwE�����?��6q�+L6'xy���K��V*	�B�[�a˾�u�ާ�Ҥ�'���T��5���R��K��f�s�]3����f阖���=M�ٯQg^�U՝fwJ:9[W�J�=�3%�J��8��9�U�V��3�t�E]�n�*�]+e�ai²�Z!�z��;U�H�]�V�0�HK{�D�TX��8���Gٔ4Z��N����U�E�ugmv�L�n�=X�q�����_=}w6H	��n��9oxn�\ɷGe�G�c;B�Mts���6)�TaC���e3T�Úx(�ٔ��h����Q����Mk���_7�z|j�3{�UWA4�yw�vN�;EU����M���q\�O9ټŃ�������[��Aju����!��O.�%�i����:YT�5C�_t�u���;�2�2��ݻWE+Ҷ���(pgF૶���]rn��r��Z�78^�ۇ��S*�12�����[�J����ZwNꬽ��2*=�2�m�<쌮���*n詉S�]���;�aѮY���e�7Ư���Ӿ�k]vu��p�1�Y�±r����C汷m�,����Y1�݁]��M6�sm���,m�깋[��vT$�V�l*Z�XY㙊�=�{��F.,�9d�K繲QMv��Jf���3�w9�T�)I*�����w?�3q�\~�����g1��p�����?|�1cH��I҈�?���`��8
���rfgc�#Y��щ�]C6�7in�\3;�a��ʎd��o�rU����f���i�me�*R�=�{�5�9mcs_c���R48��''U�!�X�1�v*�dm\�(6�r��|q�&�Y�w��n�\��G��?���me6m{珼Pŝ6��f�;㽶v�AkjV�Д	�9�]x%�v���oj�}����&B{-9���q�)z��ܰ��5ʭ+g��n	��o#eYU�Q͹�p͠A�.���˼���'��B��.�ZVf꩝;E\d^\�:�h�������Z���4�]]�Zu��r�U[5"�5:ӤB�A|+��c����]�ݢ�<w�'7u�/�pJኬ�Z��ׁ�$�6�]�{\\���e<M��a��ʱ֣IK2�[o���Zl����	L�Owujz��}6�k �A<����ޔ�Xn�p�y�*�X�e�E�*����o���6 nއ��U�
��hM�����K�3���81J�)}[�wY}��㶕̍�� �3D�kZJS�%�n\�﵁��>c���LF�UPh���bz�	⢂��1Z��o�}�ib�D��=p�K�]����Q'��\(��\�}�{�C��~j��T���$�t'+�<��79'���.�������̨"�����]�$�I(�8��0�Vc�}֡�(��p�T�,`�*�V�V[qKQZ�z4��E�-�QQTT��ؑ^U2]A���#ȔB����G1��
�*�Z���V8B�b�EDTJ�U�ˆ�)�YEKm�d�PV�Qb�b*.,X�����,�p��)VnQ���S7
"��0*��"��hR��AQ"���j(�S��^Y��r��QRe�Ba�߾��_��g�"
�r�ne?Ս�]+_I�0_l�m7���<q�O<��k�����ۉ�c�T�0��{r� ����Ŷ��e���������Є���P��B��n,�P�!&0�ݷ�6_{�@��k3��J�분˰��:sf�{���k���;եeJ;<~��f��_,R��0Q��ЖB'ÅF��v���{�q({�kF��G���bޝ,=Sp��)a���&3=�r�{x���:�mZ�����){&VXؖ��{CnR2���*;7����y��o�%�N�ܜU�=�ތ�[�]d�Ƙ2���7���Ra��H�	y"K�I��{
K�0�������Zћ��6�'���J�bsA)�d�ͮ��$�ذ��"q�W������ϐ��}_A���mV���@�9�wP����`�ܔ3[v��f��Tn��?1�Qݴz�x]]TU��/*�f�IR5��ӐY/����5W$y�n�F���Š�{G,�5��F��{�{����<���F�B������(Bfst�z�s�u1s^آ�Υ��w(]=�r|h�|N�TԊhȾ�#U=�%�ٞ�y�\�K���;��uo�Q��g`�=�#�-ɱ�%vȘ}Z\)|Ck�~�z���.����/싳c~�ݮ9�nM��K�r��s�s�Bʭ&�k�O��ü�|�`B�[��b�+�����üt��"�E�v��Ɍ���
�|x�ؖ�}\W���ɞ�LC���ޭ�!+���	�.��I�x-s��в���5x1�K�.��.�(v׾��mx=]Y��*�9�J��g*W�n���3��4��1r�u��/��fI>��Q����k,y��kn{f����Q=f��XU��7�.���D�Jc���'X)S{��]o۪�ԯ׉����\�@�\of�J]�ݺ��@�t6nHw�����{����c�Ut���gus}�p{ǹ��U���<�Аx�3fd���t���S���=��7*�4MR��}���Y�n�-�p��K������g�̳�K��m
Ώk�����	��W,��\�/3vm���1/�-ƴ8ZfoU���֧�}���d�3��y|1z��6dO�jx�N:0Di���ֲ���>w�w՗�stq�X�Y�X<�X=o;�T�\�{΅��3Vk61�琧d�!eF�mټ��5ch��Ql�hB<�����>�_R�_��w�򎽧����8$�#]�̔�9�f���N�y���kn���Xk�� t��Ǚ��>C�ԿXTro�S(j�:P9�m��sbg3F4,��:�j���r��qzH����|��"�����ɝK����W:�ޝ]F�.I����*���u�b��v%#K�h&�Ј�Awb�Z�*iV$���v����k��Wׇ����.��L��V|qƈ��
�+����)�:7A��]��S.�w�g>�*n�>�N��2v�Q�ņ���C��	Z�[D����4�C�E�������35k��]�W�p�*���Rق��t�"��5��,�9-��Mw_��SH^p1z�5�H��]��_-�+&1�{&k*��:�����>�Rv2��M]ZΫ\����b�=�V�s��mϳbnV5͇�1��٤����TK�|h,y��J�+�\7�]q7E�^�흀E^-�(CSya��fs�_~Uu���D@"sm���#�X����r��N�7yC��MC���-U����	LnU�#a�:tܣӍ�Z.wKm�\�fg	+;;���L�2,�v{(6Au�Q���9+j�u>�a|���o�1QT; ���%is���yrg���	�qj������RQ�:��cjP�Fu�k^狎�
�U�;�ش4���v��Q���{-���'V��Q*־mM��.'��فH���8櫤f̓���/]���Y�V��!%��+�pp>�"qRs]�Jl9ROMR�S˒�=y0q]���r˦��o�:^�f���kZj���:���B.<qu5՗<���$�+L"�o:I�����[��X��7��A_M�x]�ot���E]Ekg%��˸I�lzm�T�]�Z�=�	����{��MH�绫�a��զ�����>cE�q�&��zp[\B�nv����k+:ѹS�2��4��3���8F2�O����KqY��)��{���X�N�����.FT��*B�EaS��>W/tJ�N��f��ԯ�,u�!�G�t�F'[/�<��J��Ά�d�U'K쮘�6ֱ;Hn+�{�}HF��ۈ��z�;L�X�ߕ����=��V7G2o?�Ww�/�f��o�.�u��V��̞����R;���������I`�;�&���{}�n�7Oܓ0Y��Aч��'����kd s8Я_3c^����(��F�wv��O=�
~���o��g��O3"��չ�o��w%�on�C�T����q}H+�v�1�h�z��Y��[���T���cO�˒D�.y�X�'�eD�Yt�s��GE]{}��\�]Ags���7��=�%]Pe�;k�*�H�P��#a�EK�ڛ�n�қ�����ܜrٜ��-)�mp��D4,���QeutZ�P��5�wK:)�� �n�*駱	�{
��+�sr���\�;kv�n��	x�fn��suwq��SK�]�c|H����d
|�Iܳ#��X�:��`�8��$��#����-��;[�V^.�If1��P�:Z�&��ƛ7���m�������l�WWE<��O��u�
�1^��ЕN���������]I.\%:)qx1,Q;�eN�S
�z�d�z�n��:UU�7(���:P�4���W52�s؛~g���s��=��̭s�v�j��iPk�p.mf�2hW������h��q�'�����9T���%��ly�5��k�:��	���(.R��V��1!XrC�>��@nm�z�.�C�1/�,�q:�Lق,Ss]�ݮk��L��e����蚭bjL��qCv�IVU�,ju1��r5����?A�f��ߺ�*�~���0��p��s!QNfa��j4]F�H=���W��iU��9��X�qL����˴t�֍&=�\��{���Ǜ�Ip�Ө.�!��q��hJ��vk��1.1@7WV��eL�N�_r�t��Uɚ~�U��j�����uf��yn�<*��nm>�ܙ=��6v�������Ժ� �}j+��r�_l�Ӿ׾��[
uG��j=��p�%��zJ}�,$�9������NET+±��ǂ/mvçS���N([m�QBT���w�"t��}~w�9�a��3���]��H̓�Л�s���zF3���Z��g;��9�.�r+������N��P���c��f���*��G�3�c�D�V�P�+6��䧚�r�ۯ��4m4��}�=���wL��	}ݤ���¯ԥ��3oqi{��^(5�b�����Ą��׌�Њ��-������p@��RQ�%٧4�����db���v'���@�o��W��!�y�%ws�c��D�6���9[�mX3�����k�+y����ի"�;����t|3(5���˙�K�����ɷ�	�h�c��!��թ���;-���F�<�y�H�*i��Og*� �Ӽ�k&\r��<O�/f���{�U(u�W�L�W�r���`������=�ι.)��;��/bN�nU���k�i�����k��
�׊�����l��awk��6zO4J�t��N��f"�����7t�y�)
��.VU����[3/�B�[�*O�7���3��(�c�wQK�U��=�,�LQ���^]n5Jjy;�3g�z�:ܢ�*dt�#h��!H+�����TG�5��#b؆�Kʸ��B/ع���唨,���wb0Y1<��T5n^N�7^62��y,���F�U�r��]���F�:M���X��ۤ�s�ra��-u��=�p�������&jl<s±���-Fk2U����9Q�Q�AZJ�n)��]�,�KH�+`�p���Dl�yS�/�i����9����t�DG1ԤoY3<:�B�5�3ܲ��h��n���MVsO]U�/�č_G���M4��&{���u�P�̻ǽ�fC��>��M�NGQ�@n@=4ә�7�+j�V^s�w�1��Tې��l�X�����:��o�t(Y��VM[sqt�U4�/����+��:��Þ�����ͳoh���KN�oO9�M����s��P�h,�7�l!��ִ�~��C�^�3��c������;����@����N���<�5�!)���7*��`�OD�W���n\�����4yj�g�S�`h��7����=�h>`.>��99�>����5_�,,ߥ��T8dȃ�-���6�\:���X�rܫ�gm?��aJ�wܡLv�Y�t��WG�
�6�^��C>�Չ[�=�!95����q^�Z2�K��dbYN�N�ʷݛ���au[�Am�Ù@�S���J�%a�HKW�Wj{j���9�sIݽ(�����i&���H�iZ;�9�k�bU��7�M�����f�K�Zw�we �g_:�_7����B>��J���ցM�@WV�q8r^%�j�^s�@<+)s�7:�'�-���UΤ1D�:�-K��U�n�xC�H�+jt��֨:�J&���EW?��K����/{�+�8+���y�}G`�Nטe���&Qf�Ė1v<̮Ӯ�V7����A��-G�����隶�X��I����E)S��OR�a���wg$�V�z���;7]\]���#,�Ʉh��f�\b�t>&��Ԓ�v=��[q0���i[vgu��!��v���|{;�h��dG:����:�adj��5�r���V�Fo�K���P;��Ҿjnb����J�oIsj��:w�n�Gݬmo��b�s3j�^�TO�����X����hpp+��FC�,��V�$�Í�Q̗cb.��n�k�S}*�v4�rBj�8����k�3�����DK<J�&k:�R�t���m.	>�|����q�rT���s�v$�[�C���9Yk�λ�!%[7A<��m�F5״:�X��7��B��m<{VF�ZG�uI�c3����2�%���؝�ܵ��W.��)ڣ�U��vx�gE҄.ɽ!��֐����n�3����i�^Z��f^��DqX�W��Z�o&��Ϸ�P��mI�͔��ɦ-�໴EH���\���x8��mk�G���q;I;N���wdWY��U�#���t�Wʵm0*X'-�ea�Y����8˧���z�.���}2VuQP�����`�䯌)H��7�o=Mμ��h;�(���(��{!�^Y�}�C~������UGv0�^��Һ���<��"���M3�;=T�ک7��v�I�+��"��fH��T��lk���
D��Y4)�+�˶�s�a�]z��E�*Rp����=��'m��������"/�/��{�=6�RTI$m�0��*Q�+#h����ַ�g�i,fU-�Q1Ja��TŔ�EE�m�QP^��h�2TQ+)[*:��h�R�U]Z����S�1DX���]%���+2-�{����$*�EE��`5Ԑ�]`�Z�������c��Z��k�D�UX�*��p��.D�3�n]������	Lٻ3SFr��ƪ��r6r�9�UE��UW2U$��EЭ:��yX�v�2-2ڗQWB�B�r<�=TW�aa��j��Y��ɭaqE�v�8,ݚeEJ�nU���q4J���5����\UQ$�&��;��2L$P�K&Ҙ�nL�F��*���DmnZ�EͶTZ�XdU��C�����R�Й]JyA�Ds�lӓ�^T����51��2�d���6�jb�zc���]ޯ�m���x�Fsk���{�V�+����8@���x5sUS�t )J�m�Ҷl���}#>_^�s���$��"Gkk�+k.���YǾ�G�l֯����=���k��ℬ����D��<�\u=;��;" ��!��D�zE}��[B�w�D��m=�t�T��n�1��u�x��������?w���YS����ˆT�.���yې��2��LT�>tQ��W�^��+�?H���C�����+.x}_T��=�T���S��u����p��i?s1z��}���d�S�e^_���j����"2�r��uJ���z�|��$i��2�e'�O���:�λ�2�|�V�� }���O�긌~+�6��=ݿD��
E�����=�)�5�ų���BV�{�,�:���Y��\ש֖by���_�2o'CQ���Je$�vz3'�t]F�z�H�e��YC_b��*�[��9�Z���gM��9��Uso	�m��W��*�'��� D����>����1��r�Y�p��B��i�;f[�օ΢�Z;?j��ػ��~L��-��#�Ĺ��'�x�թK;�c)�۹�We_&q��|��}��փ|h�ھ؂ysyO194����*����Wr�u}�x��yK3y����.�Y���B]Q�g���2�{�+�زk�k���,�K��k"��?)<�
���e��/+럩�6��\UVtR�v�F�.#t�.ڮQ���?�;���M2_�]sn+�v�S���Q����.����&/�)���/��M̳�؊��ާU�ȸ�^�pq|���8w��r�@@�<�˪�f���I����*]N=(�\O�ͫ�ozy<V.SW6�T��S��]�p��6�5�?T�<w���=F��Rz�$���V"ם�Zow
�Y��LF3ς���7yĞ��*>h�>��/�I�DD��W�y��>�>f�J��PI�:�:�WW����OYk!¥�s��TOXn*z���40$^O�'F�F����r}k&l�F��������-���TLzFI��>V���c�i�}&~ݼ���5�ݎF��5՗�-s9Oգ�Y�4�}��U���'��٧2~����JZ����)�gc��V}�}z�4�����*k�νs�t���}Y7���
���O�8��������P��	���������ΎRD}�2��8�_w�E��Sz_Ս�h��01-�3�7��q��5�EHP�#�K=���ؾ���)�6��w}��F]�Su�l��* ��A}^�s:~\m�_U�����5�T ��*�?�v�}���a%곏}.��*��!���GXM��lv�g��o"l�����2<xpX�hV��e��Q��ώ��u��Nu��B�Z;lA�ћ��̫�m.h��&���L↳é-��{+��7��]�I�����P�S��Ut����tSȞZy;��W��+��:�(N�=�I$b? w����>�pz�$�+u�u_<e`�N���'8�9�"}O�v��k7QJv.�ݑH����Xq��uc�)=���;�����gLƸ���6���_g�`�z���KQqp���|�ѳh1|�KRN��=�~�F���qH�;tv++M��wj���=,S_B�3���S�}�3�=� ��H�w�8�_'�'̆Т�����7�U����>Fx}q�x�PY%Lk�d���:��T<;��4ɞy��o6J�s_H���|��>3�	�ph�i;��+�:Hw�>Bm'��&Y:��Y&����PX>�2u+=`k���'Rm�{`dƳ�$�`y>�RM��2�p|�'���S���=�I�DxY������!<OY����&���_RM!�2vΰ3�i�N%B}�q���I���OY5���8�:\c��տ}�mϪ$r1[��0��I�8ϝ�]��W��6q2����r�yz]#�#[�("����6���(�V���(�+֣:��o�ʏ<�t��OZ�@�O�;;;mmls@]��N��U��y\�����m�'���l[8�4����>B`͆>Ad���'\���'�6����$���d�I�������w����OY=d��N�X$4�9�&����Y&3Bx�`fٴ��'hq$����'Y<���N��f�'�:��/�&~U��]�i�>���T@��3g��w�6�|�Y6�q�c8����P�!��!��'S��O�$�h3�|D�GX+������YlzO�dOS���w���$���I3��I8�l�2On1	�C%��+ ���@g�DX�}�""~�B�[]������=�����'�X!6��(wVCha��u��3>� z��ke �ٻ�i0}�Bz��l��,3}׋�a�٭x@��iL{��<�ϖ&Y&�P�&Й5C��d�h��.>ƟRL2c��0�s�$�z��x<�ʾ����������HL�
ɤ-$�O��$�'S�1Bm��C��t�yhq$���`��3���:���=%BP޼�OxI��3��b@�͒��<ݑd�+%@�&�|�!'���$�2yd:�`�8ɴ�1Hm����۹�?�7{�����a����3�>�cx	�4���Y'X{�1%d�>��VM�d�)'>�3�	�OS3Vk M@&ϼ"{bVu}0S1���� 0����I̼���w���M �{�CH̀q&�d�RNO�VM�3d�'̝�<3@�����~�q���>v�a�Uq��Θ�6AB��E��3ppO�a�j�i�K�����o��F�[xD�A��l�d�|'�^�U��O�5��b� ��6�rw��v�@*�i�����폢�=U��Oݾ�<g����;� �2�)�哬�^ل�AN {9�B��OPY�X�sa$�M���+$��E���}�H]�W����ٽ���${�G� y2f���u���$�Xk�u�+���N �=�1���a�R=d{C��	F������{k6>W����e�,'�[2L�'��8�`���a�,�!�I�8���$��)�N0��0�'�X_}�_sY�N�3���ޞ m����4����+�I�v�L�Mv��C�d�|�a:�F�L2q3�x��2n�`AC~���3뵟|�t]�(��Dx}�@�㬟2kv���f{�$4�MI>O{a>z�R���i�����M��>�{ �?f���[Y?}Y���8쁔0�3�!�>��d����p|��O�R{��I��N fyI��͐�`f��$�T��<�{9ӭ���^{�g����OPXՐ�8É�y�	��C;�����0q���&��q$��Ɋ�'\�8$���XN3�#�}G������:��ݫ��Us��4̡�Iٛ�>d�!�6ì�J�=����߶I�}�d��	�y�&�Ry�&��OYx�=��ӌ��w�uޛ����gwI0ɴ�)���|�!����d�V�m�Y8ú�d�ݝ���s z��ke�q�=�2�<^RC��~��d}� {�*�����ZC�|����0�Y'���2�6�b�L�2��q���fǼ�ꁤ{ȏNuoRro�z�몳��ͺ��}D�̱�m���S5��5�e�]�X����ZH!Ť����K�]VΏ.��/��;��vJ3:@����_A��v��y�3�.�����j7R���q[��557l�ԓ���N��O9`�OSx�T'�u
��)3l&�:�d�2m5�P��@3-2u�!�hm!�au�6^���ؽκ�]�q�G��}?����O,���,'��&�d!�yĕ	�8�d�V���m<7��S?d�(�{�����_|�jY�}�4G��L�_�tŁē��hO�9�',&�� e�;�I8�~�T��%@�VL��m�6�/���o./���s����M&X{i�4���c�:�>v���Ma�	�;�	4��w���o4@��VT�����#��Z{���o0��a����L�9N�l&�<��I�2n�]!<@q�8�5��d�I��0�q&H�� >��O���_w�]�.xw�RtްJ��bYO�3�M��f~�8�Bd򇎒N!�C�'�^$��n�
P�X8ɶ
C��}�L���s�s������aP�'w[ąa�&~�XC��.h��,�|@�1B|L��d1�!6�=�<L�3�� `�WVԩx�>1�j]�'�Q �k!������'g{��N�|���s+Y3u�;�_(}�<t�X|�z�����������/�{�k=�<�����<I���(i�wN���X�I�VC��I:�������f{�4�8��"�m=;B|遛H>��H���!s��Y2ǆ}P}�d>@��g�g����L�O���N2���Y=}I���&&�N0<I�	'^��sfk��oF�e
��J�V*�2����z��F���Tf6�ɠ��5Q���fu9����8�*"&,ŧ/p��}Q:�Q5�����Y�!&�1R����zʲ���bGpv)T�vkl�,=�jҼ�o﷿��<ǘ�%`~�8�zʙ�X
Iq��:������N����$�q0�5�1:��l&��:ɷ��xY�<~�׹7�5�'�������{ĄǴ5�I����`
c����ϸ2u	�>I�N%O=��a�F| g�zd3�}���G;��W~����[���I�l��d��qɌ����J���yI0�l�.'�u0È)&m'YXa�N�|��d6��u��o�s&�F��!n��rŔ}�q� χ����t����b�|�Xi+'X���I�V�X��e�|�b��>��"�R�_�ouw}�e�� A��guBq	��I�M� ��	�U�x���"�i��gC�hVM��ͤ6�:�b�>a�w��W�����z��c��Ci������,����N2u���`}������'�� z�Tɽ����t� �c T&=�Ь�||��*!������)��`	#�}�#�,���>P���'��6��hE�a�b��	�{��P���$�u&�e� $�9�	��d���x����ޮ�%ABw�E&�Ry��6��{�	�N33�k$�<Bi�֬�I��$5��N!6��y�6�2zɎo�V��zs>y���wV�&�'w�dgT�&'�䕓�VL���d�36iyC�&�fn�]2�Y�I�@>#�ӝ]?e_��5=�%k�u��tx�m��vsx	�>d�b�͒�I>dY>́�M�z��/��K�h�>���~�x��}��w+���p�?	�ӝ�M�:�3����N���,�]m��UT���B'���9�JӨ�9"~P�_o=�zoHY��R��$G2�����v�5���u4l��5�f�<�5���=;���]���[�����5��d�+ q�ot�'�,��!P�'��s�!Rzɓ�`��8�z�Vύ�E��YRfy�H8L� yxgd-0�>tq�j��t������;��z�d<�dn�Ad�15��q��RI�T;�B���1$�&�d�Y'5>�'�����g�n�����W��$����$0�g�N������&�y�I�:�S�,G���N�By9�ORu'̨k�L��q����v�䫸�{6��(J���}�i��}`v�q�m�=�>Bc4�2�4ɤ:����8�{gY4�Y����2 �����{v���G�V�j��3Toǐ<d�'w�6��&��q8�m����I��ɪC�&3a�O�Y:ɤ8��{B|�hdݝL�M3��Ϙ���/�$�]�G��=��}�}���pHx�y�'X7I��LLО'X�m )�8��1��q��&�u�����=���k��"=g��p�|�<��pt�w��I�&�d�I�8�$��i�	�d<L2u>1`!�p �z=��bS��5_d|�KOR�;�'m'Sɪ@�}N>��a��:�ge�q� �z�7q�OR-Pr��2m;���=��c�{���c�d�C��0��̜J�ɪ���5d6ɶ'_Y�}�@������'�v$�c��Ԇ��5y~�{�O���,����l!�O��N$�2�i�I�f(u�hL����6 ٱ�y6��0��+�K����%�z��j^Z~�1*�j4�إ�s�q�ˣ�{��:1�uG���7*��(��n?�rQ"�kU�X74hn�$ ���N�=tz)�f��.��-F����(R�(�v�r��%�{���|H���,�>a��XpH8����)3\�Ǔ�E�'���(���4����۵+�H����|V�����H`�P��хtUM��������;��B�+�A�Q�<n��Oe�6��g_N��{)��N_H{������R�D��z|V�~�S��֧yfݩ���
έ�����t��;c����A�/Ӵ����q3R:���`^�)���Ѿ��4�O!����U�U%_Hښ�`g��D%-�9Y��}�no|p�����P<��Ǧ�VF��|�s\i��;<ݤި��w:���]��]���|m�P}�V8����S ��·ِ����߿M�����_z�=ҫ��i�;g�+�������~�bMe�c%-���nj�!��$aY۱S����:˹�K!hȖ��ܖu�����>[�s%����VX�d�^7eub�����B�DӠ����E��d �C�����ʓ��w��Hqr{\M��C]�j�\���z�o�x�w1��Ù�,��+T�IE�wW��s6����]p����֨;܆��J�B�>W#�.�Yx�{p<���k��&̗�}����2*�r�T:C�n��C���M}�QtТ,9�"�/.\cF��m�ހQI�@�(]�̆u!yRo(?�Z�5p�C�\����}������v	?��z�L[��^ۘ�$��+z?�=-��fWsÀH�f�gVl��'E����h�i�k����q�����Z�����VF�SNT�zT����Y��h���=�{ԡO�x5!��
��{��=�϶��v�VV�v�D�(��ƙ"c�i���K�jS��+�x�U���'N�p��a��/����v2�,���&�$8Vk`nfvc� ýjšK��36gq��.kn�	�՘��t2���,�i���aX���?pÂ��s����oe<B�T7o.T��7���9�7���,�OaZ9�ޟ����2q{)�~Y�P�%����������g���N��]��Е�m�0F[��ԗYќ�5�(e�{%�'Nw}%�)��k�B�y��qVm�����d�t':�9s���o�+���uiH�oK+��Ga��P�H��a��\��c�:f�V�+��s$/H��P�j켇 'h춧*qgFn͹�;��;�:�3�|�9/ >[*P�;u�J����OvnR��U�q�2��ܸ
.�
�~[V�YL�G��R��UD�R}��%w�EÚ�J�)�v���CnC3��P^�,�oP3-@R��^��s�<��)e������ܡ�D�^̜����I<؄`��[�li��Α%�ݱ�b��.��]u�w��(+	=�w�󾴌9��k�C��5�ϑ��{���:䱞�Uc$��Z!���`��t�k7��N�w�xp'M��er����H�u;����A��R��ގ��Y��Ψr�b9�g����i1T��p�*�k����c/w���.rG��m͐�� r @��3��u{�0OAݧ�<u	�s2�>-U��c�o:�����Dן����ڔEi`�U����5j*��b(uՍ9�V��0ֱ0���kLY�YV�UevM6�J��QA�ep��mJT�ۥ2a��Ͻϐ[�6	s��IN\�$*��:���\���Iy{R��{���OQC�����AU^\3R-�G��!d�X����AZbඪ��k�kJ#���|b3*f�mvv���f�fj�3̌�R��j�3*����Ĥ�ɢѱ
(�]���TRLhL��"<�r:��y*b�B�8��ETb��(�V�
(��Ub"���Qu
��*�hU�rerH��Q�#Ur��\ҙ�/� �jq�y$�n�[CR/*���vs����[Z�s	F��)��)J֤sӗ9-L�Q�"�I�~o�3���Y��j����d#������X&�rv^�X�c�,b�P�l4��*�H�7�W��꬀	������_o��~��
}��Ʊ��g|��}!�_��D:澭�^&)=�k���vگ}��gu�^)�O%�]I�d=w�=Os<vv6b5C��s2/��ݓ�)�n�]�>Z��뜁�S���G���;B��w��M)�甆��&��Nja��dt��P�yȁ�[9���<a��Nsk�e*~��.���[T9GI�<���T��[5�'$�UqLWn����ߕ��������\e���ɮ�ڃ�ݮ�eh�~�it4�خ唨fC���0�����B%��6�x�C����
���r:����>���ޛ�K}����lc=��aM��!8�P}��Wv�׶����Mm�kÏ�!��J�Ne�9��wy�ū��U�$�Qr1ڤ�}K��¥�|���ӎ����w�U2Mv��C6��_�D钻DS+�k��2�#ׁ���s� �}�|H� �����>��������o��d3lz��k��W(���,�OV��p��V��G$e>�42�l��5�LdW^5ȩ��w����^���姗����QR�jm�6>��u����M�WcB�-q5����2��3�&dμ�E����/Q�Z7����V���9r���[i����{T��5�dS��5!��8��f�s�Hw$���\��b;���mT�c*���>��	�lV�ɝ.qf;���Ey���������sG�n�?ll�{���Ͱ�f0�e���q0ߵæd��>��Xsb���rq5ͮ���7]�[��s��k���dm�\�2v�`����d����x'�a�
u��9�.���Lh���U����EF��ˁ&1��ㆴ�s(�zF�ok#���+P�'7��w|zF]���f�s��7�/Sț�+��4�sK��B�q�����?$Y�I ��]��y�.�G�|��7�g�*��
��yO�1C��"���i�����Dh�P�hG:ee\.�Pmox&���nu�򵲨���]$��sx�-�'�Z�p����Q��a�Y���q�R�UH�X���D흣�焙��Yn(��w5�&0�;#ג�w�����mx=sN��𨢅t{���]L9��ۭ��HkOFԻ�4�I�*'&y`iU�f�_��U�*��zi,zm^�,I��ân+[��8d{v��gM�]���m�m�]$G=�{N�d]�>̞����'Y�{'E;N�{J�N���i��v��ݭ��'����
�*.k��x|�	ϐS�j��y�ɿV��@L����6�ŐK�����N�_�:���u;oN���ܛ�\dS�\��gX|�����6ej@핢oP�{
;X3�,�xgv[,���|7���n3V���kW� >>����#�'�������뻣��d'�S�o��y��L{l*�'�θ���#7��8���k�q�yE�{�>�_g�f/9��p�y�eP�K�6�%QbT[��S�}O����y;ٵ�|/���e�LU��oc���B�ǡvo�_������j�έQ�N��]�_w$_�\�����y�{�9)V�i^sf�-�璋�U]k��!�Y�GS����|�*�uo<YY��{��mUz�TI��<J��� v�w8�U\_�\
�<�N�SSc�Z��}<�Tf�f�3ۏ;�""��*��
����XԱD*��,��w;W�������tLӗu���b�*�w������#��#�-n3��[�x;�w����v�o$Gi��"Nr\�������@Iu�ɕ�*�$e���H��r�۽C�&k�땎�NbfHA��Yɼ��s�ub������.�������߿o�w_g��q��\�^#�A�A���lT��Pŗ��.gSK[�un��븷{f���r����s��8n���C�d�?f-�����>\Ḯ���>R��[��m�)K���R��D޾��� t��0&���Ub��v��dޗ���
��f�HޕCS�[Q�Ó��hQ��֖��z�J��+���g�����\���$��������s�����f��}Д����SNwv#�#�TǗR�j�GH�;BȾN��8�A�.i�o��c�{ދ�Am����N:ב	���~R$'r0�k�TC�VN��p�e�j,>K6��^�9ٙ47W�g+�ru����]��:������'�bs�2�Y-
<fV��dK��4�!{X�1�z��4VtȢ�T�PЇoc�}�U�ꙗ����:"�_nz�er+�;��w�=�{��� ��(Iks��W��=�vkVQ��ؼ]_%Q
/�'����5�F�<�������z�#���t�vߤ��RX��a�iѰKВ��$���r7 䭨_��*[���^��p�5�l&�z5�F��sz)��o��i�q?����W�6����k�}YR�=+��-K����n�-ֈ���6��M�.��NUώ���=]�׊��Yɬ�~��ŉ���fz��y�*���NM/`C��`��So�R�uR9Dܺ�\M{9#Ac̷���kR-��c���r}[ �7B-m�	�ƚq��a�Bá��U$��{���:�8��Y��8�^�9�5%?�w,ey���d�Y�׶�Ǿ�����G����f�1нF���r«b��NX⾣|�92J���T��{��X�e�;mJ�\�1�Q�3b�b2�1����9=�~> <	��z)_w���U�1ض�;������0��rz�iy��{�>DmWkO�����:xavMЈY��$̷�ʦ�-��6�e����(^ĩr��J��F�&��O����L�y^xn?�2�rԏv�
�mr�H�<R�Rm�\G9�ծ���u��;�-��˓����1�I0i��n�'"��ȶ����)�)��]x�#s{�Ճ�Z�W�	�%�������2�Vo5k.�W2�Wb������*0���F�e�g[����&�}<Jw�ô�IS
�YR4:���۵o�T^�\�#-�G���
��WÐ4�B�O�ʦҝ�+p=��Q�Uj��]rWv��VLN@�nG��:k��ªN�aѵu��Y�p��W[�ͤo��R(��uu�5��n��Bv��Ƥ�����絙�w�S�;1�&[��u�
���6�c�Iν�Ӗ�������
R�$Ǟk�﷽�����R��Ž��T.Զ6�)[��긬̊�����a��-�)�X��kEX�-�W46���eT����}{XX��,,�
�}vz|�Vh^�ƳC��.�D��>��7�MW�'�3��w�c���+���s5�-����X��vG~���J�0#}7�6��Ҙפ����U�٭~�g�?)�y\v�a �F�\:���(�vgTB�]�����,�J��ٵ|.-��ag���,���J�_?Z�{&�=0��(2�C����5�%7y�����"1��dk�V�'XV	��aU˥ϵN'-���T���]$hd�a		g��!�b�Z��\KL�ry1�9Z�U]���G9�;\�T�c2��ʪ�i�+�I��gA�)ˍ�޷tC~O�)�y��E�jc6sI���t�ι�Z��(Tl\��H�8��[�o�VV��{��w�'�����"� �!5��s}���z�c��發��E:R��o*�6Z5�gb���w��M]��"��+��u�'�[tLS{�F,�oI�ȃ�t�W�PM`���X�%���$4�3�y�԰����
n�(����k��F=z���ׂ89�6{oL�e�yy/
������f&T8��oJ�ʹ�&��>\l�A�͜�������EU��v{VLMۙ��W���gVc�2FU���X�Y��3ӳ��O&i�P���P΍S���yw���gf�� �N�,z��b��X5�v��b�3z�oNsw����.M�2����������6�X�N�Tgu��/��I�4���efK�X\ek�z{j<��Ȍ϶��`ú�)�`�Z���{]/5z��bmI2yu�h��j	`�Ox\��YIݞ���:GEl��nD�=S�a>*L����D�7�V��V����<<H��#����z���ص߂�1�h�"j�/�Z��/�z�U�G:��MU�rbN�|R�;���W�8�������R�#��/
����t[Ԡ�}m��p	�p\!;��n�>���s�/��7�
eIK'[j��r\t�]�s�b��v�º~�}�Ɔ�ʑwv���ϺB�aG:Fim���B8�GL�����s�"s����s�j��{t/�Gx��Ȉݑ�K��;><�ЕW���PP����������[F���+�V�v�ٴ�{a�=�Se�}�Mq��"�%��z?_�?m�Hu26�,V����yvj�s�|�T�L���OϨ5�ih��9�Q��^h��ma�""�S�j4�Y)�AŵUT�Q��6��Vo4�e`�Eo(�P��D'$����²��'�3Q����+l⬳�5�t��{k��9���>R��ս�]C�V6���Y4�[ø��N�ťخ[,\���=��H��Lh�(�l�C~� 9}�|���UYt��ː��k�+[����m���p7�R��*ţʭfp�t�7І4��d ��s�Ʈu��R>T�pjMe�[�u�W���h�Uo�2�#�x��>��K�f9*��.|r��u�{�isU��T��fA�E��uظ�k�gĒr]*wlѳ��T�o��䵛Z�KtꢼR�!=$��  ��+����uPZ)%�n-�Ռ���-�a�h�!w��8��J���S?/]�g�Ni��{�0g+���֣������#P;[�����uEL�`=|z�:�au�=�Z�|���'Qy�\]83kם1�Ӕw8��]of�+{�����7�y<k��9ł������nc0�gl^͹@�T�M�:2-+����ǕO+b��M���jYXX����X8��W�d��!�]8}D̀�5&wp�Ӻ�s�Pch�9���uT���{�ai���r��ITuպo�����.��V�Kt/1Ӊ�W��En��"1�	X#4�m=������֛q�J�ˮ�	N�LG�Y{�
�]}�X�$�]���Q}f�t����1`���V�&R�)Q���적�&�"�������z5���!�m�T��#*h��&�7��4���A��`ܷ�MH�,H6�V�R��)D���u�Gq_ݹi;�zC*k�Y�o�Y����q'OG��U��u�%�Ėb<��oP�{�7�V ���Q,87�Ȣ[�E�]��vч�=K�s��6Ul�et����6`{�8��ҫ9�;ҁU�e� J��WP}t�$trˣk����9�+�^��hVWI��wQ����d{ԷN�ww+�:�D��'dz�AiƯ��[�-"�$�Ҧ��e
<��v����{a��;yB
q9����C@09uD�t''t(L���3:��Q�=:v����2�n���b���n�H`����u�7:��Ct,j��sg-�s7:6�%o����N�!��h�Ux����X�R���aZ2F�3�]P��dV"�*)\`�1���h�V��0�

�ة�U��ʊ��9DL���\�B脶�
�/j�n���ϼ�"�����&$������Ihy�iM����O&��|?��"|���m�DT�L<�DU��g�dl�k�k��,�K��{ޛ�S3#TȤR�q�m��{9�B��<�ɌCS�DT���R.k�g��"綍 �$�f��{\����\�C��X����aA��ȋ�2�"��$:a�vìk�cNb�v�9$kh3Y�dX�ixj�DbQ̈-CTh�]�QE�Å2�m�B�	\T�(��۬%�kcT=
0�B�v�R�&ȣ���ʖ�+Qh�e���m�S;�̪#ʫ���ʓ=<B25=H//Dd�G�����u���V�����ث]Kw����qq��Rt�|쫍��w��6��Q�fq������U�]��}D�x}��x
���Ցc3���{&����
fz���^o�X{�����پ��}l��s�y[C�F���`���b�c�9z��ȷH���嘷�����˔YV\�F�f-m�]���v��
\�Q52tC����3�9�.�!�Թ�����ja�����=�G��
�(|��.�t��u�6�{�P�羾�j�*�u���0h�����_@�0�Ƚ;�e�<^q0zO���[ժ-Â���z�+�L%&�agv�WFߞ�~�/@9jG�V�|�
j����L]�e��S�gf��8 ��p^ܙ�Ы�/sݾ�)R��2c�!}cJ�gdx9��J_Wm���2��Bۻٛ�[�%��:�N��[:cE�{�8������&fv��<�w�q�Q%�5�<ۖY����ufڷ��%N�gXъ��|�Y:��e�7�≫��/uH]�b��fEm���o����"�����;��罺O�����y��~j��L�8�Bq/��4����;��S����6)qV+�m*�آxt腟K�xU���q�n����gA���N�����*�#�J����NtּO�J���n����ʞ�H_��1z��l|�ь�kr�K�}燥�[���b��ܪ�R���6��n�Ky�'qsy~�����¹���(p�Q<�~-q�5�/u]�&y��}���|�&atM�x�,�[/��r�mOnBu�77Z����eT��ni�� ���̺�Ө�}�}��o^�f��]��B9�L��:�;9]9�g7Qs1g5����V�/O��L{6W�ݞhש�[;��n����gQ�&zŝJ�ވf�a�Yc۔�͚��n�JwȠ�4^dA3�7/�X�ݣt%k���sE��;;rv0Н�aO"��:�с3Æm���P��1өi,�Ŀ���d�H��!�<���o���ߝ:���\%���6������{5 ����;�)dX��vP#D u��.;�>�η9���8�8�˼M7Q��]���"=�� �\��'Qն(��Z��k���OJ]��-�(�������k7'�wrU�&i�狩UqLV\��=��7�΋��������T>��κ9�y���5��E�_1&��Xq�� ��s��
[=�E.��Y�9%��&�C�A5y7��`ǽA�4��Gu�y��T:���S�Q�Ӛ�`j=�\,�-Zm����_,47*�d�^1�MC�ڔ�A��[�������>�ܼ��"��tY�=-��=|~���l�fE�v�NT�p��Ğcx��ho}33��}��C�o-`��\x���|DV�+�r�t�Ko�;W���w�Iy{����kt�(��`7؛��^������g�o�o~��䄊�x��<*^v�}1�tx~�iV�3�fzE\��aI_*�����"�:��~����urxP�hP��C9�X����b�Q�u���R����A�3�:Zi�ŃzFsw�����־0�\�rmn�n�Vk7h���S��r^�(��{�E�&�}sz��w`2A���1���=�GU��
��2���MıZ��2�_(�Js���{�No��'�Z�8xz��Tu�c�{�RS,>���3%����4���������n݌ձ���ܣ����	��5����e7j�Y��<>�}pMb{���O�<�"���.+����G5D�<n�'��{�o��	���7&QB�PWD��w{���rһIh�ބ�����jMѳ,V)\Q��;�$z�PXAO��G��˕��>82KN�.�W�#�/�Wq�|��F\�ǐ�[�w뿾߾o�w���,!�@��*�6�}F�
޿ʄt��d�s
��x\PU\��U�O;���2��G�SY!K�J����5'�y>����z��w�߀xJ������G����z�pߤ�lA��寝�����/��=�����i�4r@�r:�H��y��Y��mU>�����U�Ln%~�B�,�{o���ω�R�:g�%�z/�sw�)6M�9�5���8c�5�VrD����'��~>�	K�%�����])W����E7�&�婽SS�պ��&R�<ML����=��\���ѫ��iN����^������k�5z^=ҞcR�0'pȬn����] W��ގ�g��G�x��U�wU�9�ټ�7c�V��Y�׻b�RD?O+����Û%^���T�t%�w{�S=]S^���wv�SH�|4�ǝ̣�Im���ķ�O�/��S��SI��l����7�?� E����(O =:�y�EB�'�z2z��i�_D�ޅ���m�Lj��7+�c�G4�	{Nz��=����eZ��^ʓ
[Roc�^+��������&��m_,��`����Y�nH�es�(`f#V�R��X[bxg;a2�v�kŕqLGA��5Ֆ'�R���㤧<�]��	r�o>�U��de�)���*��崩J�cF�IFkV��	3{����DT�$LU��d�W�ø��J�[��PY�n<g�G~B�DMN�L�..���c1!^i�˛s ���SɃ�4ѯ�X�
*�>���w)�p�/ELe&�Ysf����Oo�˫�Sι��<�z���hlG�h��&�H�;\��sf��E𽽡w���qZ)p����wi����@��z�����n�~9���ަ�d:�9��]�?�!^���]� ���y�c�+����ӯ|��|�~{������d P }�颔�r�~���+n{YA�q*�j�ng�\l�W���9�\���m�c��jn�'��w=*R0&�e;��Y��d؋=�o^��n�}��D�`%c������E�(��*����^n��k��}hlųƯ�j��G*lέ��z#�ZX��X{z}Bz�r�A���.8����kz���57gm}^�Ѕ��6ZD�$�Xo�n��(��(���,fE������bzx��դq�[H�I<G���a��}�s4W���ԁ�#9h�Y\���y������:kU�f��&z	&�ڶ�V.���s��j��/զF��ƵH��D�$oHF�r�mh��t�λ,rş5��Ż�<q��ļF��2$��?������UL��I��j��<�[�h�q�qf�5�� ��\;��e�CS���=�0L��)�����s�B�)��\�/�o���%Z��_��m���v��ؖy��H��㢻A�)F{3�cT`��	ӻ]�����Y!"�d�����w�wO�a�$��G:�����3Gf�hQ<�ˍ��B���Ss��G��?\�������ۈ��E`?1s�|\R���J�f�CF&é��kTL艁�	mJ$��h��pdJ!�����^~#"_/ٚ�G.����D8��X��P�%~`��+��kkj�
�����6�խ�[j�z�jg�
b�H�QƦ���]6�7Ge���[��_����^H_-<l߁�VGCM�y�*�Y܊�+�����X�a�<l�V��Tp���S}�=�ia�����/�툌���Iȅ��u'�g24��TL0��R)�Tzg�j�!��-�^�{z[G6�����L�w���巍�>	� �Z~'04�u	<p�}.#(k;�Δ�6�e³o%��a�����r�L:H<��#H����%�j�ǐ;�Z�VE-�eUԻ�d����TLa�R�Ĥ��ױ�,V��86N9��4p��@��Y|�'����Mt@V���r�n�>���Ar�thnj�/8ڮ�>]��� ?$$RI$�go[�;ښ��;ZhgJ/6Y[(����;~rN�&8���z�W(Sqb�ΛHR��D�/�3o#<'?��e*�R=..f*�A�����;`����-*a|�6!~�BR�5��ZtϽϩI�wl�5�6�s�xb���$�?;�;䏒����7��	_4L,9���:~WdD���z�=g�啖j��x��1�$��/Z��W�xѳ��)t<�����Y�b�$��蜀����k�_$G��b`^�W���F,�=�*r�wzzI�����O0�0L���_b�H�ed�6��5v�1����M����҇��c�E+��I"$g;d+�r�8VܳB�*�ر&y�qxɶaؿ(8�+�L��#�\���ù���o0ۮ_^J�J��;[9�|:	gݑq~��ՓN/�����=�9?rw�Ѩ�BPȸ�+��yF��!*��4�*��N>*���̢��D�`ɳ�Uu�Z����V�'��p�٧{��tƴi�_Kl��-�'he��U��Ek�˵���~;������~BHH�@Y�������yX`~��v0(݊�f�Z^3�@#�R`Te�|p�>����W]���k�H�l�~jB�T��}p-���j��HZJ$�۬^�m,r����7ѧ�'�jYf�]6�7Z��'���O6{�֙�4��)���آ"�p�D�k��d�f�{Lݪ�7�BC��zc�9��M��[]�3Աx%�5$��m���¡��ԥ-ثr�(�A!#ت����a��`[2Θ=��2�� ���uD���t��8�ʺY�4Ѻo���^�s��(�R/�3 �q�l�v�E�"�爲L�����mLM>OT�E���T&T�݌B���9�-����^4�O�4�r󸶯.��9_�FI�⍂�+"�9]P��d�z�_5���?^u��L\�4ڹ�p�{(и9��22��&�|lPZx�ꃌ�- ]� t�d��UĹ[�����4u�;��D��9P�#t�y�i��['[�x�oZ��_;x��!,^��"�P���ֆ�2g-���=��@�h٢�&L!(�Ss^�gU���_a�|X���YK+5��+�e�V�U� dP$oP�a��.K���Hrm�F��6k+����� �/����,�*X��÷�
�1v�4�|�p�@(}aL��]�-�e�I�X{t�ཱ�t�Z�yr�}��0�2�0�tFD/M*�#g*�o.}E@�l쨄�dj��3�E�}9Y]��m�su��.���}�)�=e��Z/���ԶУ����=�Ư/:��,�b�����)m�D�.�0�H�׵�ZwE7w�������}�.�^���b85�\ap�m��c.N���]�ؠ�9�I\���no�vfl���	�h��
�{V�ֺT����m�W��ڛOw�vM���K�E6=ۤN��?��c}^�5�h�t��guA���X�i�E�L�v�w���°�0;�Fj�8x�[��"0����h��٧���6�]����� ��Ou={��r�ƍ��3j�>y$��tC1��PH�r|���?��3~Bn:�H��e����K:�5ڨ�����q�O��z�Nr-A-T�xH���mX.P�)e�/N=Sw(�]��ڻ�����a��X����|]f�L`7	y,`����rs:.�.��u%����(�i �Rn%k��K\����'���:��	�����+/5�8{��v�7Y)s�o���w��9���yжh�p�r]Us��cx�b#d�}�"�Q�e[�|Gv:��&:���Ȁt��#�)r��j��V�<f��-nb�N�.�ڵ��S�͔qӑ�Z3�\�"��޾=�tcirͳ�d�)h�� B&C��ٱyw�
c�Cu!֖ɗf��g_jB�`ÄrO����5�(㪾���9>yV$xw�C�2u�Z�-�I��d~�YD����s�U�T;Ʃ�ڹ�4�ÛU��(.Du�]�w���ެ�Irj��u���t�q�n)E���F��J}v�w�ִx^�#����k�+7$����%/��N���;h�����7e^��0sء�p�Q'|�`�ҁ��{￠CB'���(����P��ma"*ԕ�5��bT��\ݦ���42�;�g��>nb����vCf�6�8R�1#��&)��Kdˣ9��R�f�ذ���}��6�ԣQ����z�F��l��*/:'�h�j�t"k�p�au�{���J��-&y)8��#�z&��0�mm%m\�Ckg������U��՞6�n�ԒP��圬[(O
g�.�3*/��2�L���w,'e��W�P�if�jA+��Ԫ,�9-H��AN�0+ҕ��y�������TZ�P<�V%ˡѶ��Wa�!���E������&�x�HFe�Ά���죢t�ڇaŞ�hMS�zUе�"]]U�S0�l�[&�fzh`c-�L�9wgm�+U:���Z.O���T}�tΰaeJ��S�}����eC�@匛]ʷW5���j�����B�jr�������}��w�U|�H<�_}�|9ϻ�_�/ξˡB>�W�a$Ǽü���K��郆Jt�=Un[xwj��A�I"���d隥_���
�$�bDgH`�ĝŗ&0wޛ��خ���=j��#�S��Y����W�f�4��Ҏ��r?��NzI�s���e�r��ʬh�|�_��UyW�=�|{1�j�T���4;[�/`]ƅr���]�hM9�k�Z���һ�Ug�����=�`"�d���Uo���k���"���k���B2g��ĕ����'�,v��9�<\G���46\S�g���ΐ�*^��"���ͨ����`[��>۹�5{�ad}�H�:|kn+�1[���b޵B�j��$YiD�b��i���]����%�D�xώ1��'�c���Z�|��I:_�y~���'0Ή�Q�A�&~�^��JW���O^u�g{-a�6ȐCT;$*43zz������K��q��m�Т�t���	�;=R��L��Ú����|R-���ڈ�X�on5��=T����{y�������@P�P�( C�w������W�v@��<V�#����H���.�H�k���D%�5ΕTqE�N�X�#h�F��)S*����u�Y:I'`g��b��vf��0�b�5��{L��"���ޏ#�ʸ�R�V%�͟W>;U{Ŭ�p0���T϶"A�?�����?8�=T���0ػ�M�mJ��r].g���ip|�.;K�y���i�a�G��G��Fnvx����v>�f�c�
J���v�G�h^���5�b)H@a��A<��S�v(S�a�P���	ħę�h��pdJ!���й�^~?z��LT\����܆������J�x��a{}>������N/ ����lNc��ع���8�p��L�ؓ©��Ƌ����̞;hY�f���Q�Mn_c�D��>�>/�T���k��B�G�T.�s�h,T�lp�c7��I��s}����g��ܛӘ���ꚱ�)%�]�w��n�1ڡ����ބ�����Q5ӶN@�s4�����A�3���t��Ń����x�U)��R��<�!��~�߈��	�"�d���7������8t���D��8t؏�L|�e)��7�&s'J�ɠ��)��m�����ї3{���H���4��Q�<�%5w����京��O���?8�7>����5{�S�-��vD�Qza�(gT�8U3�lr{�OND1jx��_)F��:3��T9���H.�#��ے�;y�������&�=_=�e����O���o7��#��2)Y�eŞ
;�7��95J��B��8��h.���^5���޹6)H�
dmE���9��w-)�@ޥ��=˘_'�������V�5�F�(��D�����g/����Ib�ѡ�1�43Z<�|�z�~;0K$�8�.�U�+��N����FP�ⶆ_��h����@���B��6�����񢯯�/{��5�$���S�s�]���c���]h����#��h���Q���{�qU�U�������YF;�b�[ͥ�2fa.�0T`��72*�ػ�����v.Xm7���Gv.�0nh ����89�#G%̬Xٝ�>3���yto������B~d XXH,$ {�>���;���'�9�:�������>%�ϷK�]ʚ�
## s���/%](8���U���'a��g��v�pc�L�BDO�'l�p�F�pt��C�X�Y�Sx{h�h�&FM�[�uH�(Cb�K��b���GU��s���+�x�Y[�j��/���m0��ޙi�X����8���v����w:���&t�w������a���r̵ix�_#�R�L�҈���y]���S�w#O72y�w�>��^H�����j�0o�B�g������L`";f�Δ\l��2��t,�sg:8��n����#�͏+�>�ɫ���q�^1�@�0�$�Y�MZ��;�<y-;hHyj����x;���j4de��k$M�h�;�$9$E��W���TwVW��9��u?���S��gy4cځ޴tB���5��͛	�E�=n��UT�˂�y.�=�K�dC�2���2tݓcyK����0�^���M�ۻ�XL�id��n��_�tU���	ԏW^$�S�i����5٭��\�[�a���hka��18-Nc}���ޫ���{��7��HI�$"�E	$<��߯>��+�`Ӂ�{3 ϲ:!�l�p!��W<E�ޞV2��C�7����X���7�����%w�&�*�@%��>��1�:��/i��/����/R��aw�vPL[��KOW��	I�$�h���=��-j0?} �+ŧ)U�XH'ۦQ�q��t��Q�"��Vr�G�̠x�7 �\r����Zڳ&		����9ӏ, \�C��. ��$Q�lѺ��R�_�_�HϠ�LH��^ơyw�n+K7�n.�X46����]��5K�5�'�u_?��ㆲ��\�tLk�s��k�3j�IۄI,��c��.\���Uj ��v����O,��3�`o@j4�W:]y�k���>yI�Z���I^T����L��z[���<#zW�Kxv~���������Q��DL�QN����T��＆����"b*����]s7-�B=�=!e��[�,�J�?Q��W��+G7D�gd�ohY�C��,F7x`�:� �U����.�����Mk�/Ҽ[�n�U�ڧ���x~#��� 
@X�<ַ����7���nm�\}�b���>g��5��=jǖ���a����˿�;����kG �fr�֗nIʆI��=�0���|���b{��+�(�%!dy!e�{��i����=�[�*�4f����#�#�/�~�B7�J����x,ᤉ�ZS���i���y�	�\�Li/^="�c*:lz�u
���Mkh�t�,�ވ;ا��m�P������,z���D���!)fz�i�RЬ�3'/,�U�z�s�0I,�r�B�M,z|+'s��|C�c���\\�g�S<�]�os�|��-Y�:�jQ��&F�q�J���O�òq��˩n���F���aT3�v�Lo�<O����0���#�-�C9����.�]*��0F�}��z������%�
�ǄR�崍ŧg�D�}L�퓚�*&:��B�]~����	�Ay|����T:�rB��z�M����S�����u꾆���\_d|�;��+�:܈��֩W29Щ��RÑf����u�+!�������
,�����s��]�.�+��@���Dχ���=��u8&ST����1s�b�;�;�Q�#�!�<R(D8žw�B������)�k,��}]�Nv���J]�
jY+*���'�\�p�{�N"��3��eG�:��2�{�v�ѹ�5/����|VGCM���qǗ��=�]��齊�Y�^�2ΗԝE�j6p�s������L��+��m��,���oݜ�ɢ�b{V	�T��� q_5QO���?>��ߐ��i�G�D$@#��)��W�b`�p�jQ��,�>�����b$�[�֮�5�p���Δ^C-@�3�p��+a(�T8נB+����wO%*
"ߢFD�P�s�s���El#����nQ����Q��b��8��9��D�R�p
_	� �c�i�VNp��ϭp����,�.�h���V+\C�n�Ѷ]���ZCmB�����:����=SU����i�x�K�eF੄6���f�d���A���־�6��,�b'�ҽS	�he��Zs��I)�_~ ��E ,�(I���s���_�/>��/|ה���T��<,lB�n���X|r��w�f��Gձ2�3�!�ڈ�|��~=A��S��	�tZ[���w��eY���0:|y�w��wW�!�H;��\}0	<j�U��U��n��J�U������f���n�؍s��"8��%��
�H��3�O2;���V��_�|Dt���'�KX��43����&:���z��i޵��z�S�hJZt�.:<�*��}YC)OY��=lWa�����0���wsӭ���m;0D,Z��Xkʾ�܅�òp�lH�5�'%ƭ�M�_5�<�8���A_�eo��1w�� �G��%��P���"��*	��h�T�O\�
u2EP���9�̎�e�d�P�}{tF�oϞM�\'`U�/��E�uFk��=�m�>��p.|��Q~0R������az4jn���n��궗�ƥ%�o'�VU?-�_w/ll�l���$�᛫����V]D��Z�((y��r�X�*eφ+O2e.b�.�3���?>w���C���o��:>�����_�!�0 Y���[�����U��8ƾS���G��G�R�5��Y�������MW�ɳ�l����y�(?cg#Li�
���Y�sŚ�{L��;�BC̛O#{o��J�}��Q�Z�\{�$=6���{�O�E�Y������&�� ���M�uC-z�hB����o7�c7:٥۷�T�[C���o��L�儬������م9��I�jH�l�w"Qur�b�o�f��y�gS̮!��ԸѾ��w�:�0�G1�F�2�uGYR�i(��WOU4����^����W��e*������ٝl�T$?�d�����|����f�bM2������^�2���s���]��	�_O%Z�z!It�݋{�‟m�?\M�7��B*c+ϋ�$����r�����f�sJݚ��OA�J�5�[G�Y"f;xc�+�*�����<����*E�X��n8��:n*__	�NձE.�U̵��$M�4����y�-�|�U֡�N8��}�1g��^Y]�{-�<r�2���MM	k��r��b�m��C�������G�'� '�	W���ߢdX�����D\ W,���#��ÑW�E��O��3@�d])�O9[��̇���:':�Ey,��X�e��V�G�ʭE��7Y/xh�忳w�y2l���q�nN��8V��E���H���j[���Ҏ�vn$�߉�#��ZǤ\o��+���;5�+:||w���]��9$~}Qjlr�������vY�(31x%Ė��	X�->S���s%����X8�fb���`��~��9�G�5ٞH��
�%��0��1f1��hr��^�V��l�t��ƴ!)#�$7J�A�f�-��zp�AQϭ��z��5�7�]
�w�=����0V�gAi�,$N��\���NK�����������=x`�?V��4&oP��mO����1J)}��t}u���M�A����ϲ�q����p+�O�\�L�ӭ7a]y����#���C�����;1�#N=��;� ��R�L*H�Vt�eF��ժ�����؇睪mJ�c�X�1ro,YWb���9���}��a�U�F��kz�55�e�޺�QGv����Eȥw]p�a/���
�:֢c율!{W�:��t��غ���f;�'n�;Oyex�2��Z4�Y����f�Ҵ���y������F+�6��;!���H��fLhv���:����yI�I���,Pyj���Z�9��(����A�
9��OJ'u�)�+<4<�w�B��;�ͤ�gl��vտ�*��4���|��&��
���j��S̠���1C��̀� g {2�;��2�U�]Q��1�M��vs��S����8��:n=eM���p�3�v��*1F�vMւ�5�m7�J�7l�
ܫY�\&��
lycq�^�E���Tkr��������8Y8��0�Ӻ�ó#�R��5N�f�l�v��x:�9���i���_j���Q�F��9�g�lF�;Ry����Tfp�L�оj�2RF�O>8:u�ر�6�r��2��XV4�V���ko��3�RR��=r�	���'EY�C�7*iv{+�z븷v���P�}<��+�)��mXbȪX����!��3��2�Y5��Y��k�xk���)֊���.<�sB�up=����MN�����3�v�qD��r�M��!ݧ&��mk��*���Fn�`T]�6����#��Wj�3����C�M�@yK��Ū��/y�������`���gW]a/�,b��Nvp�]b�Ӻ	��W/�wM�-����uG �P�ܒT���9�cD��qm��t�Z{c���.���@�;{���{���u��Rn����/^J�d�=�|ﯸ�K�
c�d눰 �=�N�G���p$�6,��ٲ��-�����$(��a���i��u�0Ĺ�\�R�B�:�G�m>�3��\6��b�]�x��4��[xi��V�r�����t�J �(_�W��غ�o����껬�i�mv�K]K�%C ՋM��f���ⷆ��Uc��Ius�/���$�3'b�*t�@$^�.v�:!�ѓ��b�r{���@�]�㳑EEo%W������9b��U]G�U ���l�p�=.+l�X�u�$�%�9�Sh����xPjB���׽�>��g)*N]谔9fz���F�3[;$+�&ɞ�5X�]�{�>Z��	sȦ592�(�T��15)9y�xL�Vp*�2-aR�
6%j\kZ֍j�n1GE2��ʣ�V'=����J�Fф���h�k�^�����4�#e�6�����V��L�ن�RrJ��&�G��q�Y5�skd�2fE)��i��x���EƤ�"r�R��S �ʨjɓ$sJ�$�� Q(��$+<�B��t�;C����^0�fI^����	qP��h�%6�&sP��Q�Dp�P��EZ�-�*� �ds%�E
+C]�	4�綗��^A�:Z�j��3Ϝ�4W�n�o�k#�<}a�$jh�x�9gD�N�o�oE���ʩۍ_k������x�^o�䀲
 Wk��>Y�?�A �#m�fGU�3Z�^؉DN�k�ʸ���ܳ4��ؽ֖���u�С[�rI}�Qm�f���:x�R6�V�9�8������3sW��8/�P{�2�DE�ͣ�/=!��rg���}��e��o7�V+�5T3-�p,(�,	NUT�ʂ��0K��Ҍl���^Mw{��*�]�e�s;�E䆠�jY%�k���P;D21��o!��kRu�r3.t�*?�*�ȣ��ر�W��g����D�ޭ�[�-��{D7CL����Cd�4>��	�1\�l�t���y�_�]#�w���VE>դ0.�#��qD��L\b\�K�?nѬ���zǹ�9ȼ��	�oe�9kՌ2ό:���Ŏʞ�W���I���ebծj���hRN�ş��S���3����"l�>4�Oz���m֛�՝|
y�����toi���I�e4,D�@��9�륾�C���cnMGv�*����+
�e�;�T�X�L�y�΋[v�͝)ቛM��zc���]�Ϫ~B)���c;����;�]��~��7�ϜYP���)�P���`H(�y��_����k��|�H��j�N
�*��}
#qK.�Yt�"uei�g	[�eH4�+>3Ɲ��x;͠��U!�"�S�� �~>�~#~������t�=�� im.��w��l^���(i �;AcB�?R&�x�!����p������O׏*h��k@��^P%��S��/��BR(�7}2�[z�9�8h5.�L��� -Q���K��%�)�z�	��V{�n�E��Q]���A�cBSd)Vƒ^�����H=������2ﱻ��.��l����*DldK��a�
}� �o��������hw%9⡆�����<j��b���@J�h5�elZSU�{Gj��<�p���H�C}��Д�զr������a�������^��%�(�'L���%��/�É:���(��o|��o����t��VI}��,hk�
�nFe�AaX���j�պ�uȚ���ѭ:|z�ə���+:�-��r@��X澻����������)d	M���W;Y��9����gFr(��j8�+2P6h��˭�*��oTL�Wu8���p=�;Y,��%m��DY����s���) �U	�o�v���v��H�s$U�H�Z�2��Ad��"ۏ@<E��z���Y3Ⱥs�A}F/����B{#����ӷ�ʨ|P,އ���p���;��e^|)U������g���_,���Q�76r�x��^�^ooG��gs�҅��l�i�!x/��ۅ�9T�_����+�%�{���e������E���Ǧ4�FL( ��D@|&d��3�cȺ�=�(y��Jsˑ��.�o��+z��Z{�>�]!7Oc�ܨ���Ԟ�#�����+k��FjЂ��Լ`X�����z��ͧB��m�OH��XD>I���V���~��N����+e�/7��E�x(�M�K�(��\F�16�{q�n�7o3��\t�r�:��`c7z���г{aӶphه�;[?����,�*��g��Sv��L�o+�����vV�]�o�{h�����?�����H�
 ��L{�����W���c�y������/�������{T�S_��H@�΃]�U��ҖB$�Sb��8䃱K��#j�^^"��$�q�kdSd�x�'M�A���t��0@ي���"�uP���I?y�����`�Rmc��X�m�7PtӺ�U�>�Hg�^����'�U������nVrz�e���%C�J����FŅrϴL�x;+Iϯ��,�6�|���T���w��0��&}�,��xcBV]˃�n"8��V�c:W��S�ua���1�Xb��h�.`Mܳ��p�N�����-~�M������˩H�/�{?n2lW��-c���z"�z}o�~��}��K"�T�E��-��j�^�g8�EZ��x��{�Y���>�ǐ��*s%�>����n���G9A�b]d���9�h�/�>kO�̖|If��R�K��*4�����C�P�`1�YK�bj���w`	��K�����8v���A�,9ګh��+�;˜;�z�H�rs�7nj���.B-�O�*�SV35s��/k�W��|��������@�s�����o�Z��f�|��b�P8am$�Bv>;[g�OA�=ƟW�k�#�����sm#�CiJZ}+���7�J����a3e��8	9���	�s�����*>5���_��q��tp�������D��mLM�n��ũ4F�E���}�\Y�O�#�C'�'y���37N���+zҵs��J�݇���Y/$�� 3��du^�45H�0�ހ��/q���WZ�R�}9J�pڱ(�0/y�J7�%���,X��LRæ��'�DF�K���B_���a���ڠ�,;~0z�K|��|����Q��e�z���^�1�,զ�d�k9�,;��:H:��<`нJ?1z��^l�W�ٽOџ}�!���I�@��܉�&I֦�Օc�"�Z��&����|9*�1�y�6h�,��?��!.ұn0��L`S��$�띭�����l��d�\�����
�xZ]�TYe������'wN����Gv�Ho)�fD���R�7��,�OQ�c�$�1tj!��V%pő;j���p��ս����������o���I'�$X`E�x�X����ׂ�ٹ�E�TC.�:dU�S6:$�p)F͙��qgr���]�K%qs�u�8l��`�^���q�(�C`q7jED�A�������yJ�|fu�5����(m�gl�Ю�����2{]���[κ�����8&oOb=凄�*'�)�J�z�^��{]=w��Q�>�{#iL� ����v'�T}��\:�$�E������Yu��詂gXɘmك�t�u���s*�8�S��);�T[�qT���Yc�6	:F1B3.���:w:Qy�L��G9K���4�]���N9�Z�����˓��A#`@��hx+>��?���^<�Gv���9}���MV3���lJ��:�o5�"8�"=�GP��'�VP�N���X�PQ#�x��.��ɜa�ѝ���,���*��gX7�݋����v&����K<s3���yNJ�w��,�]"9�X�Y�1̢�JてGL�f�U�N�]��w��bW>�\�vL_aZ�T�1+�M�
�d��p��#2��+N�]��w~���ܵ}󯪸�`�"θ�0,b������֒B��>T2�u�����z�,f�||)Y��R'�4M��V镰Tz�A�'w��s��<�N�=�^�����	�$�Q�Z���z_�9���_s����!�ɸ�j��������<�*���.��!�����cv����ش���a�Ce���5�z�������m*O�Y����ݐ�!��%��Z}j�e\񡈞k��T}�.���X1n(u����GNj6�{["^�⫗�!��lmq�Z������h(7N��:ɲ:��zT�@��n/a^N���!�Խ�W�UZ�Vت��%��&Dg��>V�!���Ӎ^=>T>��ҖY�t�l76s���"!Ds���gpל���ō��>�4��a���*��d"����zkq�#���]�F�Umt�A0�d�K�i�����ڴ쫮�ILcxEb�ٯ�O^7k5���;�9�&d ��fuu0x�z���)�\�$ڏ���y�+��^�:a��a�"����j��ǃ|�g/��x��y�����P�=Sƣ%yD���Wͱ�_7�S�>��b������ݜ�8��>�/���!X؂���=�>�l�V�ԕo��WW���M�?|~!e]��G5�#f`���⻋Q��0�u�R�qaȰ�|f�zX7���w�:���B��A'Ko_to����{� �!
ݗ�=r�W�es#)g�o<�Z���ٝo+��F�J�B�v�G��#?%�XkO�$�_��_4r$f*�ő���C{k�G����TlŞ����u��kM�:�����  r��)f�4�s�y��i�u�LL(�n��uL�Y0]t�(ɬ�A�gg^��a���'("+P�|Ĉ�gP`�R�DXLdR�f��\;�f����H�W@�����g�GN�6;&�X��pvHd�^K)�l�܄��B�ı�����!�s:.��6��B�O[U��.[/����`�4[z22�3D�s.�W��[�1�_�-��N@�@�ss�̡&��ĉ�=��gK楫��7�M���[V��=�˕:���.}�T@�_�H����}�=�:��dfB6mM㾮���Ňr�{�<=KΒ46K�����S<nd���ult2�uH��՗M�ob�t��dQ�7�dME���I�ؑ[�\G����8�i�����%�iݟ
y=jǖ���#�b]�r;3ʾkO�z�7���+�:�oWZ���Tt�^@�=,��$^@�0D3M�
},�0�;�����e�ޕ5�3�s�k� z�;�W��M�
��34!m3e�N����K��YQQ�cΕW=P�5�/ψ�A5��B��"E�hά��վ��l/����1�*a�y�Р��-�����'I���p�>u�����QǺ�"��2L��I�4����x�����;K��O�}YQn
�Y�q�M�xӡ�jح��g�A�΢��k�K�K�5`W��WȆO����sf���c��c��;�N�&�!r�d�;^�|����Dl���N����r���f�iPF�;�-�g�W�˲S�ݹ���,ܭ%N�ݲ�<������y��q፼���\�Mu=3�N�U�d��o.,��s�v����I���l:�t;���s㈜���WQ���S��ǝ��K��sfP)D`�Jp��eAG�u�����u+ȋ���R|\�E<�	�Ș=�ğrF`W4.�C�0GcԸ���6!J��l;dH뛸$Qy����j�����V^f��D�r��X'ޙ6���ֻ��P��y���c~853�
b�(�+�V�q��~��'4��\��ͷn��8]�q�	�*eN0�&]�zL��y��lO-��_O�-,�G�,TYf�v�bm�CU޴�^�S��X�I����B��=��q�z���OY��ئ�j�g{�S�{<W4�8�8��f܍Cby��9��8��,��p����ۺ����9�!n'����4��?c���e�N��7�'�0����uަ.Kk18�(�t��+t��6��Jh�w���d����ЍORQg6�m��dB=�u�^�h��`+�w-�jsa���[�j�� �
�j��FVP���
]��L=x�Y�V2yc�gv���R<#ő���o=$��*���"g*�S�m��X��Ŧ����7�.���L��j���0ɑ�T�G�b-�:� Xg�}����ݝwU��O�b
;�m��������+nNvO$H~�z��=��/[j���(�9mwek&��M[�`�]��-gb�'�Q)[�і��O�r�$&��Tۭd��i�`��2SZ/�jѠ�;�����շ��ow���!H������+lާ�-�+v�Lܗs����k-E�N��ˁC��:�S9gp
v�vQ����x�N��ɶpP�VMD�n�Y�'d����$a}6�ݡnrW���9�o�6CӮ��Ȼ��-h��c�S��is��lޮ�g�:Ov0B���)�kB����s�L��N��Y{$�a��Zs���wx	����2]]�d��VU��%@��3�9uX�ը��"�9�w1�����]���U����Z�K'��ܽy�+&.��r�j�b�Ԑ���p0l$�h���Ԏ6C�O�:Plg�ZG���l�k�[�C��m��Ko^<{��$�[+��֔�5��
n�P�N�*P�y��R�n��끜�pƬ���Kk�����7���@k��ca�쇲:�f�*4�n.��.�/U�Q̵:�c5����9|�&@Sm��$��˾�����&)�j��l�{ϛ������\a>��VK-K�̣�P�c:t��.��3��/ps�H�����`�Ŭ�j� ���3�s��T��d�Zc���M�)R�٧.�^��wj�{��z��H%��;ӫ�Ɏ?�{}�f���i}6���	j�5m�o�Vs�m8�b�BDk�9���
�˖���t�ڻ��b�n���u@�].�D�T��Lp-:v:}�m�M�I�58�D���R�P��,��+�1Ι��v���u��W�A$���I+��ݣ��:ѹ7(��"��Eٺc)�|�t�/���u��oV��\���S���D�԰Vu������noq9pP�k�/9���͊��z�ِIٖ�׬�Sz���gY�JT%k%UB�
��UKUDKi*ѣ%b�k�ߚtX4KPR�P�m��J֥�F[A]Y���[n5�kZ�b�d+*V�am��Ul�QQ��ֵ�i4�Z0V� ��"�`�ԬT��5�U�J�ڠ6��Uu�k�ZTYYd�Z��i�db�9�Y��^�iz�zI�z����iG��Dn�:�T"�G�Z�iBx�PZ���E)*%�iPKTX�X�����Z�E���QEV�Z�X-�-+��"���t�Ԣ���WB-�ŕ+R����V#�ł�Z��Uk��Q�ԩR��T
�.�|�յ��{�w&.�k����V/mV������_5����z�h�[�kt��tq>#��q�I�I�w5���d��"��`$���D����M�"��2$V�/�U�
����7s����$�*29�8 �v(���bP�8D-�L%P�uY��=s�C�6�Mҟ�T6�����yD8'Or���cn{	����1���m6Hx����ϱi���L��?*�z��y��($��y̏��>��K2�w�μ9�`�&�B�7�m}��gۯ��(Q��
/u���Z�������>��T�X�g�r6�"|�i�s���+`ڟgd&B�h�Z���$���,��]M�IS�y|�?�,l�Q��f�"�e����VhՔ^s$q�CQ�u���)x�W\��ƪ��6b����*�|��"{i�rj��S��h3�}�a���=�\�K}W��GThR���[<�(�^F�r�`�}�"DƥС���Y��F���lT��Cw��G���Q�勩��{܁�8W������.�'��f`(��䱪S�.�Ja c���i.	`�B$��W�lu�(����s��S^s�X���9j�a�#Xǘ�ȗ�����v��CW,�FD2z(I�J��>e��(M�l'a����Cȃa�O�h�f�z��*Vf^�u�Bφ�e��#�#=8����ō��}`9��iO�,�ۜ�W��y�?�غG�4�L���#�s%W�$q%	x��:�'�)(��R;������.����,��B��GT���'���6�􍑓��
�x,�|�d�Y����k������e�����cc(،�=䎟y�_vo�S��n��l�$. yw�������L�Q��E4!� _ֵ.&��>���]����'\�ҳ'��2p�$���"�H�U$�MӪ4��
�ʷ7H��|����
�m^��ޞ�������/�s#)e����A�n�����f�қ��xmBC��HB�)>v$�����"}j}!�#�k���%��qк��`f+�^15oy1#�����ξ�<�f�v�szkPJ\��ant硜��E�L�yճTq��c�i�k�[�\�9���=x�t����U���l�V��p,櫠�+3\{� ���uW�Cw�uY]�Izy��x)D8�n��u2�,�.�I
��c��ʲrg�r�����I7G����Bܒ���<Գ���E+�i^<fW�+Ӕ�f~��EIچ�K�V}`�v�z4dat���0����dd�:�n�-��_�w�ԍ2��\�c!�\@��gE��B��iZ�A�3"x�>m+��8<lmǯ~&�܂_�{)��t�3��<<�;�{��o� Gak+Z軓e�{H�ʑG���"��ȄI�ĉ�4;&�/�S�9K�Wv��lO�>���~ZF@ޑ��;��O<4��蛪���BڇKo��S|I��4�<}��_lų��!)a��0���U%����}��Ҵ�|�$�79!Tj��x<D�|��e
�@ܔ)`�(z��AR0f�f7��Kz�<U0�6�;�31�d�5u�4�#8#vcAr]Z�T�1�|����h���+�c�]������r�o<���dXq�p����F4��m�l�%�ߪ��{�'&����7c�ep���r����nvu�4o��Z�����O��i G��`����1��0邹��짫=t����D�G��a!+�Ǧ{���N�I�Y̟ ���~=�E�;��K�NZ!�r0�j]�8)��K�ّ=��."�}�G+L�<�)E�\�j�M��C(����z�#m�6(wA�U����SI=�G�^zC�^V��a���^o��=�GE����s_�'Y�`����lv�Iq��_=����u�Ru�"&#`k�f��2(����Lw"{J�H�7/=��'��ֳ}grǆ�T�W�Z^B_��؇�TQFn&�x9�W�e.�)/���t��I�J��=�˃�h��*�N��~#fxU��*\v�w��T��ꉐl���7�r�ٵH�H���)_�~c��'�T��]J綦V�PY��/�y��և��X��������(��t�3�V)�=��L�eG'hU�:����n�c�<=Cm��7_o#rذ�S��[G�hv�L��&:�eoMM���s!>W4�<��U鷽$�}��E��#L��؎P�(,T�tm�2Qۀv�~�&;%�oYV��9�3�pD�D�<W(�������q�jFPT�%\�쇢5�Y����TÎ�1^��k�8󟾈���)�~�����sb��P���J�i,=<A�X���H�uL7��-C-��]#
=:Fqf��+����"�J�!U53��	qIi�A��bW���~��#u�ֲq��sF�������rN�U!��^F�|H#Zփ^yJü�ןq���-����2�y×�>��ƚ
��Y�S ���Q �c'�㲲ksT�4��Cr�HJH�-w����4���k5�^k��:��W���U�z\}�F����>��5���Q�Lڡ��uF=�
��xj�	��c�9b���S�ǭ�h����b��^�<q��g)�D�*��N�3��N�B�zV��a!9� <��&�X�qS��`x��4'p����ͱ�%f��XկRfZZ�i�\r�k8)�M�w��PHvuf�1���c��sD���JZs��Ԅ�]�7ݻ��D=���HB��NR�����>>?l���'(pؖ�wv�quQ`�_[��t�G�j4�A���)@1ibN�|i��v�ѽ������L؁w;@�p�F�pt�ۖD�%Z�ö#{�w{p�
Ӭ�n�]�L�!�'*620�	�o����>��z��Yb�|�[��8r�|��{Vk?}���ۖ���U�2E�ܤ�[���\��[,�'�pE���J��:���/#�q>�f�$�9�)ƔZs&߹�{ꗻ/ggX�)��=;���p?l���/L�q H�F8�y����"�2��5�u�I���G;���mnK��߲����b�_�C���g��P�-P^�Y����2���f^߾2l�ْ�P��.X�.Ђ�-Ù�]��#�'��c�Z���t{24��\s����#zb��"�$�u#��Z{� 69��"�����O��9��y�ں�{�����U#]�Z�#�:Y˹2�h�	_dC&i7S�9y�y�f�h��QN�V�;;1��*�vv�yj��K���V����D���Ӻ�|^^ji��#^�M�R�}O�n�Q��L�ڇE��I��r̙���ˉX>��a����Դ�ms�I.6v?��@�t�XH�r�S�a�GtcDlDѹ"x��qи�8���4tt2��t1;R��N��Y��T���Q�D��#�A���C>2������F�
i���]��N�Ȝ���S457ê0u���J5�=}Q��� �^��wU��k	'����OC��,�Dp�޺�k��D#�5��]��N��kV�(�BZIv�cj�Iq1n��bG�Ws��UR��D������Cm�F�d�˜I{�{
��_��TI�fƾ.yM�}\� �Y~�`;\Y֙���GE�x}��Y���U�f�/D���8i!��e��,��G�b߲q7ĘEyp�[ý��%����}�:�|x ��5�Z��!�����v_F�:�k�s{��z�G�~��'���m_5H9�w,uY�K#]�G8w`�e��:���c�5ׁa����w;�U���9�j���%��_Ov#�F����b*�q������n�r�Ÿ����f�ϳbS�㋟�o�\F@ޑ��0f4v}N�0�*�\%j�y��Ml��Ok�S*ώ�6[=�����HYa(�H�7��B�I:��Rm�Ou�z�F|�Z�k�W����u���J�ՙ%^��.�-:|�4	;�����~|oˈ�-�r��4&�ЇvЙ��nȳ�I��_H�2/D�?T�	ʛ��~�|��TH�_�j��ZI��&yJ2�*�v�2��<�	8F�� 3~��GW�i�;7Miҧ/���bf,���i�W~�LٵbY�+3��v ��>�]ũfy:���۲�cD����wc��g~飢ۡ���!�w1� ��~{w�j�yRD�2�,Ѹ1�A�>Oˍ�rN��h�`�+?o�݇�C�͒����|����{cL�@�]�F�����z�*6�FE�����^ٜ�av�G��Q��e��,�6��:�jn��pv������6*�1A�[��&k.��w����Ɛ�J����տS]�̫��"(��nE?1s�"���4|]sE=`�Lw"{J�J��2�pp�z�v�mR;��j��m@�����D8�R(x�V�e��Ås�2�Ӷwq�N�F��F��˃�h����w��ߦ	8�G����X��mwM���ȸ���h���O�o}r�ٴ�c��/]{#@R�w׮s�.���s׀��B�s"�9B�X�������,��.#�8F�ۻYša��ݽ��L+��|�x|I����4+S��N7!z��"e�R:栮�M��'W{�����g�V��9�,FB�p1Cqe#��V:%=��\���� r�ޝ�fy�dO���5X�@��q��p�aH�ӊI�ģ����;��J2���b{a�daߛ�8x���W�Of%�����9QR�y��\ڒ'a��6�ےt�U"y�?���v.�L	��:��2TG�ιݵ���w�䉮<>=B��u��QQ9���ԭZu^]Y2.ˏ{��m���O�4$+��ʽ�I�ڄ�J1w2�˘�O�6��s�^��2s��ld3���T3����&i���A<��p��ϯ;��P�ʛ��p
���1�������^3�э�q!)kH�ַˋ��3�s�}�1���Z�K����%w��s�<KiG͝�zv
`�q�E�x�С|���5���1ݭ^��{Yk����$��N\}t$�t��M�جs*9'f�x학9�&f5�fgWCF����'6G��%��e(݇WT��]e"��)��$��h�r�����#\���/rF�(Y�5C�3�q�)a�rt�F�I�U��=�ny������j�N\;��1"'9[�VG�/tF���Ltm�Z��7=�����I��s2��:�r����L@�m��U;�yR^�gVO$���+4S^�����%ࣳկ��ᘬ�#V�����s��J��l/Ť���u�j+�޳�Q��Hi��E)S���}��l"�:��9�O�0>
�+���Ȉ����&?�>��'��j��G�:TPg���V�kwJ�f��|�gVj`�q�\,��nu�����A�3:�l���$DG��Q�e
��d|��a��؍Ι]��he"��1Q�q7�w�l]�E��3��&y�JW�;��fCN��,n\V2�KFc
�ۜ��Ku��As���n�v��fdn���]�ˇ�ȳ�VcR6v��Ǭ_D�%P�*l��t�P�i����)�?a�����}n�V�h��,vMjV��a��'P���岫q�L�C����5��B�aw��DYA �P��C�Ώ%b�I��Yd])�o�F��v����f�A�nu�ʵ&Q���.j̑jDfAL.����l�f�	�:�DZ��O^`�u� H\���T�>�b�\�5�`7�X0��If�p9�$KM��7y�t"D��}��k�'on�:�S�쮫�u���.��RԺ�Ү�\�ѭݝ�K���-6r�N4t�v�89�tk9���u�ۦ���j9ݖ@$=�Ǌ�K@���9�Y+L뙗��b�a�RZ|G	`�ZR,2ݱ\-I��uW�6UMS��W>mi����'���L�p~t�]=��{�ݽfž-�e��,��\^�b<�f�]-m�m87��8EFY��E���gh�w���d�5h��v�9�=���kG#��p���������d�T��۷���VBo�^���mK|���ib�d�\Q$vC^5�Oq��}�-��&�i�g� �vr���l�i��1�r�=��Ʀ�1�f́�w��*�g|]�όz�6��؅K�љB򳮍D
�][0p����F�����r��P����%��Be�:��I�rWb����p3�}*Χ(��ԛ5w'���~����h�о��?m��A�렘w]�n��9��SK��3w��n�+? ]^�iJ�ܺՎ���[ї�8��*�q,�-U�ˬg�h���om��\l�Y�T��Y%�P�u��]�ض��r]r�H�y��n5��x2j�m������S�S��l!V	�[B<i��v7Y�������b{���,���W	RQ��tv��{7�oT��R2�����O$6��Sn����r����u{ݒ�E�yO�0}�x��Q1aR(,%E�X�mYQE�o9浥ҭ��(ʒ��,��9VQ�yFeQ���G��(Q
�kZ֍Z���T�#%j���Jł%e�D�F*SZּѨ�Kh��+l���%\���t������7[Qk5�k��AA*R6���� �V+kJ(����lyi#�*I$���
��*�eJ��ȖԩF)X��T�Z�J�EU���,Z��EK"V��U�&z&b��	hydPZĥR�1-*Rж��,�Q����j��J��T�ȭ�
��Yb�PY+�V*��+$m��$�%�&ꔞ*n�(�}�.@)���T����Y�ݍZ[�8έ���fl<�mF���I���:2;�9rWz�O��K5���z�)��r�43񫌨*���7�g��H��`��:z8s�Ƕ�ҳ���kݲ�X�OG'�m�:;���4�П"�0�ƣ@5s3B�r��o.����q�>�l�䴉�V�8x8����~�5���V\׈
L���6�%x�ԥ-�^��y�/��_d�OD(A����Q��K�)��F� �N�Qw2:��t#o,}X/�8�~q]��n�[�g�6@a�=�!r�W��������|}>��Q�p�7�gc�	�D��Ou��wK���z�G�0A�R5�����^=J��̉Gu�8��w��Ե3st��Q���r�T'�I9�)8�j�WM[Y�9�6"`]S�]k.�Ρ���U3a�0حc�.�q��Z,#)AQ��G+}xO�O��7�vm?|��> =�3j�6�Í�A��e�q��IZ���ߔ�Ҏ�i�]�צ�ۼYI�B��Wq����k#I�Gp�E�Ui�9���o�C���(97i�7b��Z;gm��D��ga2���%E\�d�=�&T|��?�$�N�F��a�Z}&A�~B��I1�O��8��ր�C���`��d����pO)Z��1*�❿;I�a�И��H�E5����c�T��r�(xR>:}u��Ły��qdS�L�â���Pn��[����z������ػXl߲���e��{���2q����v�o�U��Nv5�g8�;Q��x�z�x���3i񗥆U�\r"�bFo:��C�2�Kj�8`4p�0��&3d�C��x����9<fcGiYgN�r�`%��]���p߅d&r�N�-2�{ ulu=������K���u7��^b���QX[4U�K*��T.Z�4)#
+����h}��qV�T��Y/���	��GP�+��q������*��r��S5"y���ͩ�̠�/!s��F����F͂�E�r�,�y�c>6*e�]��d�;(��Uj�Ђ������5f{q�)��K�g�W2qUp�Ց�9[k;6R�i��v�Юs�]q�8�+��#�k-�o�zFζ�2�K�*#//�;h�\P��:�m�J;*�;�NJ!�mܛ�'L�OM5\ǋ�Y/|�'�;��'ŉ�����:-��,�	,Λ�*q�C��k�y�'Bt�]A�΢��rP7�kTkR����s=����^�`qr��}	�O�:�����I��*lXv%��".ы�Z�����G�s�K��"h	�!=Z͠�^<n�I��$E��ˑ��Z|�%�q
aeDC(q�\�����q��H�@�1܉��m�Hm����Q�l��֍�LdJ!����������/�Ɗ���ս�{ۜ�����4v���DE�c��ٸ&+�'�,tȚڤlUc�ց�!s��֦z͊�Y���N"��i�#�8l��2`����"}�\	W76�W<�9e��V�Hb�"���]�(QK�`�)�_^��3�E0oZفr�q.|��Z���GG�gִ���?!/���G��{+՞G&���뻐|���l�gn�֤5rv�6���U�������~;+��fE�kYYv`m�i3.��NN�vy��݇9�ϩ�vV�u�p�V��h�����B�=oR+YU����h԰��`0�QP�P�`�Cp-Cqe<���	��Ѵv�̈́�.CQ�T�q3�A阑��RM�q�R˱�����jWK���N�B�q��ʦqy�T4�e��/�#ſ���?�6�����>��,�6m=�D��5�_E�%�$�R9�88a�H#J�OO53w��?;Q��ˋ���E(މ:)O���mŎ�L@<�B��g2��%ҕ�x���&8��=�!)F��kyq�ϩ2�3{����Gj�ֻܽ�=�K�=~=M�� O\d�g��DU�6���[����W��֖2<�
����X�����o��Y�>���_����EN�C#�oVc����!�Y��<rl�0u��PkqzP��T�Ƽ��y��j�N�m�o�'|�ҽksG"��3Q�:c>��t��Zms\��/.���/&�s곴�&}]�����z��+	R��h�S]��g3����i��\ �&���78A�j�Zx\��x؜췂��P�e�vsu���Cj���5p��n���t���}n�j͜®��YC��4Z������D= �F�R�{��&۬���#���wӕD�ĉ�T�-)��0�d���|8f��=�ݚ���=x�[c���~̺:��X�ν�����.a��:Q���p�^;�/���"����p�4>�N,l"�'Tre�ɇ�M��U��*�+��흺�lx�㢕��	^�t�͎.MA��ݍݬժj8Ȱ���Cݎ��G����ڵW�Eȡ�_σ-<�'z�=�}���L�-^8������ϫ��4�=0+h�<��ʲzff���S�u����CM"7�L�㴥,�+�8��3T��0%���a��w��[U{٣��Pt0cNjGǳ�]!��� \�����*�:����U������aL�-bTZ�� ���+��JzE��t|X9����՟xU�*4�/u�ۢv�㬤��%
������]��#�!z�)�d�XǼ7;zf)�`ν\L�*��{��a��s�����J(Ч1w��/���9�VK��k�Z[:�n�N��[��ީ)U鳩Q��`k���$sV_�==?%�+,_��������z��j2˔tߊ�6lL~7C�������Mq�$��W��z.�u�zRW�n9��Ɲ;`�W��cP�x:��Фh�J5�=}�%+Q:y��Y4����J�P""ӑ>ͪ@�	H�-�rx�]S0�`������v��ҫ�H��=[,��4�h�1�y1B'U�>7����/�ó��]e����8}�ծ�c^bU1��?;h3���턬�Ĝ9U�
��D�ݎ��N⦯?ta����vTd2��o�ϰ���8%��fۤ�{^�>#$���x�S�̣z�h�K)!���,��M܎�9N@�������[v�KM�[�qa����YΆY�X���;�p٨r^�y[g�Uր�������;��N�pX~�#���{�ʩ�����g�u�f��0{K���uE]h�+���i��~	\��]XЉ<� ěB_�:/�͙���~��-��8��O��M8�,�|8l�Ȏp����2�,��YRwSҦ�QV�՛��f��(�����Oz�d���jҳ�����Qr�g�Z{��s_�2���׋mï��H��#��逝�j�:�~�؍5���=<��E�H�c�U�={(@Q́�Kd����:��Y'�:bN��:K|��i�ּ������~�l��U�or�5�g�ٝ�C�{"�z�@���y1�)�i\�J�`p}2��M�'�)h�.p��K�L�,Ή馫��t,�7�Y��v�x܅�Nu�v��I�Gz��R:��O��AnU�ʖh�,ҳ"@�0�FeC��F2u��4� �1�+�#�Pn$\2��p4t�?(�a��=�v%��Ɋ��W�=�\�[�'����=���<X�#�L��#AS,DfN�;�K�u5��q���uĖ��֣�5�E)q�k��,eL��ܭyo���c�>kJ'´�$��Χ�j���O�����h�ix�G��w��RK���ڹ6b35�mcd�Hd�W�=����Xt5,N����^l�0�m�`�/��dJr3��;�N�>���'���±�l���t޳ՓOH��9<�%�6Y�i���q������2pé�`�}A/"j�����Ô&*� KMuO}��J;.�^x{�7��D�(fP�G�%�p[��d�v�_��/���g�`��5"���Y�l|.0�L�s�4�285���
!b�[cP�y}yZ����a����@>��L^�S��G��;kOML^����_xF+'�Z(��w�M�(�F�ٺ��Ħ�S�~�US�f��|��}u�����4z�ztI΁�e.W.>�M"e����c=Rp8`�~CWg���V��c�DKl�='aY{����NϯC�*�3�iY|	qDqy��o*��>ָ����]����ӎ�s�N@���6!@9'K��T0�."�~By�ir{N��Y��Ց�9��y�N͌�ӟ��A��B�Pu4
�.̻�Wi�;T�^	xު��h��XC=oR�0ص����ԙ|��MOh�k;�/�(Z8��n�J�f�|��Őu�;\��TAw��|ǎW�'g����T|2�Wݮq���D2����s�;���p�U|�J+���%���6x���8'N�	way�[�v��h�h�P??K�r�'�ѓDu�﶑��+��3�j{ݽ�h��M|D�3�HAz^%���ߍ�aF���0]2wT�[����&�E�0�*h��6�ꐎ�UD3��2$p��]��	8�v��>�B�>�o�_n��[���$�YD[\n�ث���(�A�
�Kɂ&�븞���]����殤�,Mmq����}?4�"u}`���j��ݹdITBS$��������F�P��k��Ց�(m�q�\tF=�<��qx7������T|5�}����^=.c�Lv{��Ehs$]nRF��'�Ӵ�.s�۴�	�Ĵ����?0�����]q�!���{)Ɣ\����=Q��7{TT֝y�����t���
�3A#,иʂ�"��HN��J�+���j�7�0����5�
>��7���r|�����cH�FLH-Z�z��O0���ee���N�H���]�7�ђ���u�H��Eon���Y��|w��zS��]Ĳ��O��(=�|t�8��@Ƶ�I恘�J��Zݥ*����Ògo>sB8m(oW�=<s}�szkք��q�(�ق�*��}g�;����򤸺I,;��~Ҡx�()n�+�8�!���`>Ww�,Q79c':fj�f�4�H����Z}>���66�����Xe�y8e���"�w#Cu{���\��qi�0��:�}_\�j�˙Fw�u�o���nb�ѻ�7���0�k�-�p5���]Q�<
�غ�7�{ȯyyj5��y����6Z�4%K8�IgA�H��1�@�rA����s/���쮯g�:M<yxR8����^"��8����cP�y�A�4Y
���-�U�M�F2�6CQ�V�/
�	'�����<h�k������� ˹����-dt��D�||a�4=.K�yW��I+�'{��Ǹz�C%�j쳂qRx�w��f��V�CX���%SS�㦆ۆ�*�Q0���/��G>�Dgp��V��'�ғ���
՞�d����0e��7�F�o�=��{�!w��u2qMf�gh�Kq^��N�v�[W�Z�]Jg�GYԩ.�F��v�d�U��w��5��nm�7�U�ř}SO1��b��L:�T� �^@v�
Ӳ.��w˘��o_x��m;��i��Lhv���Ȣ�E���g��;��1�7��p|�U��KM�.��u屌<ޫ������-n;	����7�)�ɘ7f(�;�e���Eȋ�@n.{%鰉����:���Ȫf].&����Q� �����z����Do ��
�h*ZHwF���^�Y��8)���zY8D�:^��h��̬���k��ml�쒷��]�8�SW�0Z6������CQ&qu�A�)o�߳�J�=��:�]�77�H��Q�͆�H�ڥqe��b7��`�ٶ���nji_
������P}݂�n_a±;z�,������X�ۗ5q��&���5����&���>��Jw�c�{hX�2a�0�G�'��]n_�q��L�F�M�·��J��l�k>�\���[��C�'�	��:�04�J@�n�`Č$�e5�s�!FW��}Nn#��7�ɝ��P��y���N�Y���n^@��#����W�u�������I���������+���B�RL��kB�sP�.�Q�+4�"ol3f^��Ocń�|�Q={}]Ӣ��ܷ������K�r��u]m-z�,NކY�Vs��p��D�ݑ���6]�%u�����*���#����pb�2!��Xx�ziu8
��6W,'R|�H��Ow�z���$�M�k5L�b��CC���p��7]s�=��W���;_t�F��{�e�e��_���ٛ�:4H�y4��������R�U\����WW�~d6�.7��!b����m�<�+`�B��7mP��6Ĩ��}��E	��]����2�������;.�nP�Y���SVtni�5ގ*����MŜ�ۼhU�j�ٍ��3Ji�mUI�rC|��������0���zG��8p�vu�j��_dv��)G��p�s�|�\��nx�ʰ�3���e`zGuX�n�gM�Ƨ=���
�3.|���Ax�%T
ʢ�X�%ab��Ͽ{�AMFҌAZYQ�J�"��V���cZך�ƵL�LBjt(
3�,��ڥ[Aֵ�jвi-kQ�{�j^b�I9s/+�ih�X�]kZ׊:"�j5�DRa�TanY�
Z���4J�j��Q�lFX�EW��W%������$��yAfZ$Gk�dH���J1B�(����Kh%�XX��(-�KJ�F����F�¢4Ub���I���g��WI
�r����aE��$�-������%j�R�Ⱥ�s��\�BBT5I���d�-lp϶q]�)���T��	їf��)��=5μԠS]�,k�bq2NSq1����ڑ��ݭK �ŒMk9�����Y^QhC��&4{>�:� K4�m�p�wlZкc��}����~��"��oi�֭6Y����*xO=���"��Ʀ)���R��}�.0�Z�j�񞾞"�Gf�i񗥇�U�6y9���/�����K°0�1�ˆ\T�TN�W�t�?}�S(��j�*0L��w�>\R��l#$�Q��5��2����^,�u��}��H��}&vT�[����HB�X�/�=A�8��*�j ױHYQ]olle��n����:������*І4��D�-G8W���R��K�q�"�Rn4_�]_'�꛹,WOe.�����3 ��p6������E�������I(rjs#��{id��=Y����{%�CǾ�Y,�D��#0+��w3ގ]�/²n*\�e'|��8���Wt��<�fF��9�WXz�rfͥ?P7R�lV��*q��ך��S�6�R�x��ţLBV���H哐�0�R�W1҂�wjnuo,�S�1r�D�zO��9����X1!���ˌ�����e�ڜ���+���i���F�>#N1\`qTt�,�#h�R-ě	Hys�y�3����{�pk>�i'�h�.zC��e�Z��!D�V.7�8�h�m{eL~��s����!���N�_eDB48G��ȹ���R�F���h�m�]k���ny<͌�&qzI��Χ�j���G�U����!�c��.l��gW��Λ1���y��3e�F�PFNHg�܌2�:g���D6���m�#Ӥ�Z�b�ȵX6w;�}1��W�g�a�9Y��\���N��ב�{|tc����8��S���E{]P��r��K;���Wp��wey_��xNW-_��-8��1���#_x<>$�Zz}�����0.g�������2��콫�⚑E����nk�!W��J����#z���c��=5ν�)���甩�����������;�1��I�ᕯ�C2�ѳ��V��8|rf�v�����<�8��N�3fk�K�s�{���c�,eY�-zo�/�>�D�Zyj�_�����ټL��4�T�������Y��mBh�﫻�;Z��g%|�m�M��t�]!�G>Y^��}pW)J��C���0+/��6����X]��o}m����6�c%�5�ο7���:�r��m�Gm�:��D�p]�����^���ţ%����F�R+���A+��<����}9�{�ȯB㎺g+��fr�ַ>��(��T�sK>C=n ���kK�����ԙ����eM�n�[F��lzuD�J�ǒ�ܦ	�4X�ڟ4*5��U5�������c��jk��cZIұ,����ꙟ\aE��^���I���.�3�!�Ó"}�_����z��`kqzT�G.73��VC��ʼ����k���	1��n-��w4r<f�Htϭ֜���s�ٽWׅ-/�2x�ܮ*��~,;��~+�n>+���ܳ&���I��v�JwFjl�(�F(8�+�ʄ# nI���K�_�%���+`���>��hw����6D�5�ۛZ�')�l�����w������j�.r\�n�p��M�ʌ�=R5�39����ޚ݄�	������od��wLMwi��j���ޞ�{�{���ΆeVg.�&�����D��)ʏ��&8`���Z�ױ�I�]�Ɇ��eɽ��ةplo������U��YVf�h�6�[�<�a��Wvcz�R7-�]�m��gOn��scƻ���0XC��2n�ӹs=�7�[,_=*,�Z�YޗB�}6s�x���v�h䖷�h�&��r�m�4+֭����'�)������x��5<i��7�tg�����/�N�_3k1�1WL�1�z�.;�����6w��	��V�/x�������r�0�Ua=xg�"��֟W6{H[�x<�{yRvunK��5!����[c,�L��P���(Z�C��c��>>���)�`\���IL.{�՗�k�(�[s�MP��*�A�:���|�f�Ai輗��]FX��ƶ�jy�fT�ĳ�J,�j!\�j�P�a$,ִ��v��9[o��w	�F�m�=�U�����(�=3׽�VS�͗���Z�m�:���zk�ڝԕ�Awp��\��y�M'��Tæ��!������Y�V��u����]�|'4N��WQ�ۯ3����8�;I�K۲�����{�v3G�uT�U�"�y>��|5r�H��8k#��(����N�����f� l%0�Cs�j�V�Z����vC�Mg�a�z��\~U�+�I����[�ȥQ�vM��:���6�񮷯�;��%Pc�����[nJ�i�G^k����ny7į}:i$Ou�´ѧLv��k��b������ǈ��i����������p�7C��/�e$m�ߗ�^T��H'��<��Xjә��m�Ҁ�-p������Z||w���]���ظ��a��B\�T��ow�Sͨ�f���a��xK��g'�l�k�~��cˈ�ޑ�N�퐜/Uw�n���;��;0����Mt2Oے�f/c�%d�����r�2'J_���J�
W^�)]ށ�2f�%�%�Y(���E�T	JS�p�N�N�WY�Feup{�[앦-8���ŬJ����zW}��_Bv먺\�u�|�#�ֵ����:r��[B�TH�&�`S�(���0���&�)iK�f�n�N$��Hg�p+�����0��|�:	o.Ea��.4���{����m������\�g�	������D�"3�p/仗��7��z{ ��z�;6t�Z��-!�o�y�ܸgs�}2i��<_B�{�1���E�4�d1��5���{E�Ģ7�#��Wt��6�K7� efy-�bI�ǹ�^���]L
�x��4�-;ʟ1��}��+���"3�	]y���Ȅ'���f��DH�0Q-i�2>,l�͠�#�Ǎ�$���q������v�7U��AJp�UPumė�z��\�����C�,wt_$���fr}R�H���h�ĚjQ�:�)�Ck�����*�O[�9�.&_�7�^�D>�)>4S�^��jŸ��"�UH���rN�Ȇ�[�=��f���s<.aL�Ƶ3�S��4r��.�~9�Y�f��R�s$:�wsl���4Ջaj��̂�"<Z"�v^P���]dc��,�u��ȭ5d<�����f���c�>��7�R�˝.��'�Űh��Ll����٥��h����NN3��s�y���ݣ����w�Q=V~�w\+$##]P��P�(,T�tq�#i�B���{{�������Υ����
�S��s[�'��9M]��BJ�����������W�s��VԊ��Ps��Bp7���xOOv�y����=7`����c<������H���GX����RKJ��kk��=������6p�}��W��mJ�`𧝻R�@��Y�.y�Iv-J�Ib�GE�D1�Y{����D��͉Go�I�*�X�}�ٳ-v�����,t���ay�"w�o��1;6�������T��{ѝ�G'�$XU0tGA(�
D"$M,t������kM���]�񮗎�^����:�i�	�66mD�h�S��Ǩ7㴁=FM�㶘c	7�;%M�nr���PkS_>�ccIz^%��OҤ�h��t�~B��R����Z�����г-O��gy�����=.���k�����i6o�O�}�n��R�J�/���9����HT���]�b�7:(ޝѱԮ�8ah�\��n���d��S�|�w��¼'�=q�q�'a}hֱ�9"8�%�Gmz^꺫��뒙�'�W�Ma&6qD[Z��w4pɂ����0���u��skQ���J���5L^/�=<|i��	{����v����j��t�a��ܚ��|�rXv��0�ztlkHU�wwV����T�;:0$[��Z�J��n2!�ǆ��5��5�Ras��Zs���r6��ܧ���N�����&����S�u����R��t�C4}��d���~՛n�����y�s~>ܘH6���ݵ��;�U>�>��|h6g�WS�!�2fg�Rl�ɇ��s������:p��t�Y���Y��V�S���z{8-s������*y�P��<Qq6�::2x���3~S<jА�®<r��H�S�7��k$ND6J!.>���iVG�Ҕ�T�hr�����8h&/?_]ԗ3��*�DǓ^�}B���0��d5���U���u^����s|W���O�6r<�A�Μ��=�s��L��:��$�wq5�!�g;W�rή��[�,9�V��Vj"#s��Y$�� l���kGD+OySZ}\���5s�[��=��o/��sBg%tI~p:�(kh��K���Pa����Ҟ�D����]�I���2͛������;�0�z�/�/$�Y�)����^���GC��}N�:!.4�ޠ�"Y�w���͉s��蟍$�ޘ�O�������{��֣O�r��0
FӾ1��,c|o���B��.}��jpL]���Z9�#�YDe�	�_TبA���}\�K�B��w5��K��E�(֣�s{'z�H���Rq�����H���Lz\��!\�V7�V(Y�@ԮK��ۋ�l#q���WT���z��<���8�o�N�f�ǽI��u�nt�fsj��Y	On �ju�c���j�*ר_��/��T�X,�����'03b���.�������fA��ٻ�>�(n�=�yؕ�u�Է�z���Ֆ.��۰�hdz�w��3�F��w��4�:ݱ�oe�f�p�\JS��W�N��1�;�Kٖ�:r�C�֮���ܣyK:��5<eΦ��u�s@��@w9��oN���3z�9W{�-�^�d0#z"��Zù��Y����z�x�j�7�����V#w[v��Q%���Qv"�bD�H`�\(�����4���=�Ǘ�����n4_�s��tFa�S�.i�{z�ktL�K$���+%�=�9j��x��;陛ڮ��W�
��,��X`��=~��*��WD�!dQˇ�[ǻ�������7�AZ�w��&t���I�/[OЏ��o=^i�u���a���2�=oK��/}�i㶠�M�h����oD��/=��w�PJ��D�Y3��W��cs��x�t�F)���w��s�f��P6t������W�U����F��±q��5,:;�F5���J酸-��Q]Ȭ�f���w%N��_,RyQ1��Z��v���|����Y�#�m�oZ�jY�bR����-*hǌ���n����^Ix�,�7�XMe�F������3�f��3�]��F��tL�4����a���џ5����H[`e`F�Q����{��|U�u��n�3�	��-����=�e��o�p��Ѭ5�6.�n؈����s���p6`�	��0Pztϔ��R���76	;'N`�`��/����60�:tV|�kw6,mop���\�_�#ْ�p��N�Z�
�hn�(��u:�;���Ǫ�oI��\�bT��1JaYt,�\�b�|'k��^Vv@��v��a`<�[��$�s0���٢���N1�L�|ik�o�M��Hv�teJ�F:�E$o�|���	�ܲ�r��VM=���ϸT�!���$�z)u�w.}��{�jP�q��շRX{:��Z;l��Q����Wn@R﷔x��>��0��1}�3�v�W�{��w7U�ޔ���{_RX�ʻ�-�<2��dp�v�JY�)�0��;}�᧧-��q��U�R��ި�Փ�d⪰�QZS�I�!���i׻�E�����#�k�a@��e���ev�d�zYO����3���;�s�©ߏ�Y�!���1D�
z�!6�fQoyb�8�r`[���L;��1KΝ��w��\�eQ��0�Hż�X���f��Ht�%L�S�db�ϰ�د.n�V���V�w�]���"�
vh�N���B���|^J�9MfB���0p.�Jk���^S�����7�EU��M
[�9v�v���UJƽR�n���Ah:���1⒦w�a���2�n�eH��]��s@nu�t�c�__r8�b�31�3�N�����oV��Y�3��A�#�!�y�z;Rů���t/���Si
\�zTސ��2�*���S��p�1��w���kc�n�t�}�ǝ�mr�7�3o�\�ׁP���!�V�
WWS��F��	}��Z�gLŗQ�.��4x�{2����l�FJ�Wg�$��ݬ���f�5ݛ�I
���V��pڣ�S��Q�wᘳ3�:��ٽ0�V�+"�Q�6��C�\6�Hycә�b��	_e���e���ʖ�X�+������v��36��j�<�w�ټ�M��cۺ︊�+o��#�I$�H�R	"~'���H�h�'5�<��vJ������}H��ɨ�ʮix��l����T{0&J��.��5�t��Q�0�,1��a����[R�ֵ�ji���"�T��zA�<���QfaX,P��k^hѦa)�6����g��$�ƣ�ʲ,YP���E-��,�b��-�b�����"�m�<�+]T�Ih�"kn��e���hG��u("8��3�
�DXѰ1t1+r�&�*�R��5	!�����2!$��&B�Ꞅ��fF��qݜBT/fE�2mr&M�啓2.�z����v���B��qZ�:�9�xa��Vog\�ٕg� �m](y}�)�f�.�˝�:�+�nj������K�؞�c��6�������7�X_+T�oKx��̹�_
�B�]0��H��o!�,z��G���)���f�TiU�$�m�H02Ҡ�=6��X�ێέ��k0��oJUq�&{z.9�p��-�����Y�o�fV>����e�Z�5���Nn�6�:&�<hPŮ&��)��͋+z���j�ؽϻ�>
T�.j��Ô#
bg'�$�k�'T�7/��5;9��a>ܥs�<MH�6�G�S�cH��V�<J�\]y���)ݪ�;���<�\F���ʋy���p�+tȽ�=\�l	�˒��*�ʊ]�p�M��d�Ϡᣁ����h����5K�b��=��z�Df���.BE��u�y�G�^�^e���aB3��x����� �j� ����-cz�q6l�2.�K$ni�ԯ���73��: �2V��-�"c�J�W3P6����F�q݄�o���v${��A܄�g�������@�{6�y��ቊ9�K:R�}�$k(oq�q�|�A�+�k���'��o�}�s=u��nb��U==l�����\V�2�\�.W���#��9�<��~����]X.yeC����s��:�}D��*��U��d
���8����x:>�D���m)Vm0�kM[I�DEK�*o(k�d�5y\;������ix�Է&���9	k=ԏni���j�\�!��ԃWU��#�][����������ʶvT�W�e=Ka�eeu[��dn����b�l�X��fNV:�{vV:��zrr�����rĞ���[7|_�}���
��aR+���,VK���C�CΝd�Bx�V�G7�U���C���8��B�l�Br�����Q��$�ѹ@�,�2�B�)n��闼uoGv)�#�0n��żw P�{y�΋[v���7�6m����殇�:��j8'`׌qO:��_{�y��[���R_O���D�׷*�Usb,9Y�����y)�N�7ٷ<�&嫩�˫�e9(��(�g=,D�f���>y�q
��W%�X|�%SCy������j�O,�㮰!#6����:][os�R'�����R���I[(�u��z����ko�L;�Z�����Tۄ�P��)�ڪ`�"<1�$���n�v-w5d>Y�LG�]y�an��ɰsa<`Y�in�<����'���ͦ}Z���ѱ�c{�\�.�A�g���������sY�I�`X�P�D���&q�ySk����cQ�$��v��4��>�q��皍M�9	����oEKm���ʭ�d6��]�q����v���.�
'�t�r��'jkg3��Ck*�)q�T��:�\�z�����]�hTr�R��M��q���k�ur��x���=����d
��
ō�|�.Q�Xe�6z�e��J�+C�����7.�����\����-Q2���y���1r�]�j�����	��Cɽ�Sx�7n�-�U���3׾��sU=�͙�!�W�'2F�53{��3�o�&n:5��~.��;�ĊG�>o)��&����E]����w6aނ�4/yHNoS|'���ׯ3q8��G,=�����B"��'Z-3z��{���U���k%K�}Il^k�chnW���`O?�_4o�M䞭���ꮻ+S5]�q[��p6$�}<��ޥ�Ri)x-r�j�\Um�J�5cߌ�[�u!S����Rzv��i�t�����;�������ޥ�>���')��հ��S���m��]�7��VW�e	5a�c��u$B�����I��U� �����v�ն���uM}@��}�Z�!*�l�l��20oD ]2�R��M'���c=�Ɉ�a|(�B*�\���1�d�4g2j.�Vs����u��6���~�=X�
������Y���雳B�!<����6�2ܹ���2��+v�d��9
<������[�Y�6
s�T�D��x-s�TT�W�`��$nA5x�u��b]4h\]�ւ�U�T�w"��UnD���nI��N��j��%wE�炽�V��U3�k�`w���{y�s��K_����l�V�,c�a��8�\�j�oU�]TqΛeV�Nr>\P�t�}���Wdd͙��ٰ�y�<oc�|��}\"ڳ�0M��N����10��7���ػ�,Z�r��Ю%H�r{L�b�a�d��f^�+O�/Bp��<���a�%�ځb�f��r]�-�~���p�7l�
E��*g7X��� ����z��|�=y���6��-��3U�۰NgW�z&��;�/IyZg�!�/�㫵��k�v�5������`pQ52{�Q������WҹT�N8\�{9��l�~^+d��F�n�����҃Ƨ4��jb؝
|+��5���x���B�*�,����uǱ}rx���qӵ�o���9׼������O��LRI`ְ���ztI\�@�5���uj6��rvu��*��t�ٝ��C�2��u@�"���(�ܨ�;N3C��N(K��u��:B�6��,؎\V�*�^E�ؑ�L���[�Ķ�E����]X.yev�qݻ_	��r��J�O����Ƨ��2�<�v{J���m*�^W�B[����y�V979 ˎΘwSn��q�OemI|����<|�CԈD,o6�����KH��ݔ� W-�7�����{�(����j��i��_5x�����f�5�s��R����XH-cQ�37�z�
����/�^GH��1���s��[&X].t�ŋ���q����y�h�a8�jo��T�H+���޺5������7�]�g�-���zUU�>?�3����kN�٥�s�̯d~���.vk�ū�Tg>�^�,���j�OJ���H}�bU�Ig�q�����rY5a73���Ҍ�~d|N7�9fo�P��y�)����<�U�w�����ʝ���W3�X��q1W�Ƚ{ݛ�}�\K��j������NO��h�.����=o^v��xP=V�2�]=�U�����'o՞��/(�25ݒ݄Z�*yÒ{�L�;�QʔX[��oy��"��X��0�-��ӌ����e��cב^�N�]�]�T	E<��W�c<���vV@��g����8�j*q}{��s�*��8�G2��vΩp�L��X�mh5rt��3~�f���ղ���O�5+$�N�������s���Ar��vj������X���m��U\��۠^H��ﺡ&����=�!������<mEr�=��,`@�*i���B;5,�)Ґ�J��YW�yf�.QðFJ��	\�,��������ǟo)o"#�������=>+\Ԑ&+t,����Æ����ƱE�Xw�`��D+k�E]�虧,��3W�D�z���,M���'gX��{F��8=5N��zb�	���T�'
����n����_��o��qj�͹�X�F��k��Ԫ��� ���FU9��3�Y�mfd�y=H_����f�Ui��1{X��%[�YѮj���,OrC;J��]�'
�?l�����/�(:�'Zi�ՃzMŃ�3�P�Q����Z��>ޱ7kyp���ICQ�����Y��=�Ud��CNoU8{
�K\���qr�XS�u��LW�)�k	��u@\I��]�Ò����϶�R�v�U�><�}�7�>���5�8���&�Z��<���|��0��\��_f6޹�bwv���y��4u�y�,�t:��J�Bǧ���;O{*yə\z�1�����J��鐧=�F�d��-7w��H�Zi.�C`t���k�d%[��94p3zB��Or�ձ���[S#���6V��Ѽ�����+�������Z"�:�_}Yhs�5����iR�z�1�!_^,-틱�^V�|�o{}�B3N�������t�'o\�W��{�>BV�pt��w�S�6郒�.+$�J�B�:Ɍ�<���Q���\�Ϊ�+��2*�
�g���u=&W��}[`Lj�@����gs1Q�D�'K�X�����'��D�f4�C8�'�e����\Z.:��S�j��v�%b��n����h�s;�fW+%tC�%��/����i��o3-\�W<�\mNzR�v��o*�_�N�JJb�HFp7�cX�ߚ8�M��۫�.n��e'����y#aۻ>�j���ؽ�e}��2�������A½Q%�ʕg��ώ9́7)�C�1B1���E�泗5�*w�3Oe��Ҧ���Y��Z!�L*��k����ݻސ����w�?�s�P�����z�E�X��ٵ�lN�<���\�̤'y/i[R{nJs>���C��u&�F�`��֮�|�����f8=l�f�sf�/u�� l�w`K�{��x�>�L�9����2�"�O,��nČ��v9;�|��
ꢷ뵟|ڞ��鿌;$�p���gή���kee��Y���fsk�ױ��y�.��ª'���AT\@J H@Z�Y���BI�b,�`��F�����L��z]����].�fg0du�?�������G����3l��X-b�Zŉ��h�$X��$&u"F0ZIAk$�d�	j�""���;`�c�<�+�
 ���(("��(1APPPDC�
("�DA���AAAPb@DADA�"
s��&L$��􉤅�@���C�&u(���y��RjK���4���BBI$��H%�U"�̭(����W=e���=7W��h[��i27�.�,�L��:���_%�fHg������ԡ�}K��KX~�^UK���ФL�!�k�k�B�$ '�F��߾r�'`��_y%�l��	!$�ة4C��	O�!UD�w���xzè����Њ�d7�?i����O�����T��9�	$�;}���tI�$|/U�nr=*�T����#���bI;��)%�i�e{�cX�*����G��me�Պ��&LIkf�H(˝��s��J4��ǆqL�J�����H��9�7J�Y�2Qɤ��L�&B�HI$3���E�`���	I&�C"-�Z]c#z͵"�-s'��)S�{47�ѓ�� ��Gi$f�Z�J$Z��XH��QE�3���:I����tq&ǭ�#(Z��{~]�MFi�~
�󄌷C�G�e$�w��'�s4dy?����k�Ga��f�jRZ$ &N�,*j�:R���ݨ�#��[�`��N	�=�a��.{uH���<y<N��Un�:S7���;�����K���4z�O��6:]���/Mx��P���:����=���!�S#au)��Û�ȭ��R֑UϕD�(��P���	�"�T��
��KJ�#�q�Y��%�fI5���mM"䋳�܍� �$f�Ê���**M���,�J>M��L�PI-%D�i2Ov��q:]FĚ4ھ�T�*3]e-k%#�a�Sd�c=����=̳��0��	��2d���}a��9��Yi�_>k;�=/&�N�����%{��?�J7q��R;9K;����Ο����|��'$�;�#�t&9#�C��',+�wR�������9�����Q&1x��>پn�la��%�	��93�t�L�R�Ҋ��o�b��!-�!��Sd��>��5:���<}��sN�K�#�z�ڍ3*TQ�/�w�u*J�K���ׂ�
c��w��7ԩR4M���2\�?۪�??��v�I�]��D��;N��T䎤e�X�7��.�0p���Ȩj��B�W���qe��[�I���uZ6rf���$a�T�wTV�W��p���P�H�D�>��.=}HݶďB����������BI2y=x�M#��v��32�Ve��k-�_�tz��M$s�T��Ţ9E��ϙ�$��4��.�p�!�g�
