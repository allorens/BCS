BZh91AY&SY��F�_�pyc����߰����ae�}�}    |D�    �   �S��`  w�@      @ ���h �   k�c�P (@  �   
 1� �`�� �   �`�2�w�vs�U֗3�u��e�ݝ��=�v�Uu�-{�>�N�]|���/0�[��(0N�V�tt��u^A���JP��pk���A킻f����v��(_b��( >��� ��6�������m��A�f��p��@ݫ݀���8j�/w$ ���M�9�kɤw�;�����o� 2�B�h4����4:5n�svM��	�aћs���� v�[H=��<   >����u���<�n�e�s�p:��tuܰ�w���ݱ����w��L���x�wx��wluNh�m�9���Wv�`:����8�-�Ͱ<�  @ ��zx(��;��9�G��Ug�`�k]���æ�ݶ�k���l��;�u�
��T;�x[�ħ`8s6n��nl]wS�6���gn�ͮsvl;�^  =����e͖�-b���d�N�hgs]X�l]�]�V`��wv��x����UJ�����nM��i�n�Õwlݧoo@� ���)���6��      /a�  @    4 j � �                   T���JT�h&��� �i�ɣ Ja!$�H!� � �b	M���U(����d`1��I�J��i�4�4   � �U"&К&#I��&ML�S�fL����L5J���`##4# #d��'�'��7�p���Z�f�_�g�+a�$QP��0�"����@@?�S�����
eQE*���?��m������������?_�ח���u���Z�DH���[�T�P�g�U��~Or�* n(��Dl�Yѩ$��n	.�DQ����R���?��������N��*�3�s�L��U?d�C�����.^�w��*=�bs��)ȹ��V#�E�>I\��հ����bbt�ҹ�9�D�	�Yԫէ�&��v�Ѵ���O&���l�7�4Mq��g��Iʒp��6$l�=Bzb>,�!�;�M�6sf�C��ɯ"f�$��!�l�X�*'t�D�#���Hɾ	:Yh��<SҺYdN"WZ�&�;�!��z�Nk�DGmW��n��(��`�D��H��楉cw*�<��ҝ'�pM�I�r�l�f����D�$DrId�b'WM�u����uȔ]�&DG���t���R"u=��]�V&��H����]6U�H�R'<��΢#��Å�D�r�.��(sS]�����:�".�a��ei��H���pK{)�W0J9w+T7(D}8"c0�XpoҴ�epٷQ��"`ܫ0��Mf���6ܤN����Xpw�Zt�R&��\��D�:5��2��nR&�JD�2�l��	�N�ӑ#0�5�rI%tGr	�eWY=�U�j�rVd�D�0��='K�T^�=���J���U��ӒXԳr%�K��Drx��el��t�� �T6�})(�U�k}�!*C5�K�JE��1�+�ds%sf��LI��'$��ZzD�vNN2u�W�1�<<�S��4�G*W�rI㌃��d�9"5&;"o"a�j��Ux��A�ԋ���J�q*�Xy�t����9 �Sޓ�Ee9=�J�����/B\6j7	��!���~Qڎ�n=�o�[���{٣�o����ZWX�ܓ�����;��z��D�x�kv��A���O���*���eVI�\�#ɜ��r99��.M�ƥ=�rRΜ�+�;ٺ�U$;���oea�u]Ȟf3���S̓v��D�Ι�vj5���z�n��_Ę7�\c�MM'F�t7���6r�7El)t����E�OO���;�T���O,����8v��d��8N��LH)�'��+eN�"v�y3	xzS�n���p��>'�|Y~����A%�/	�N�ԏI��3]0�I��I��q�{�]������D������Rof�oroe7 ����y���P�ITa%���<�<��$����u;L��βw�<ɝ3l��$�]�z,6Hɨ�OFM#��HvK�&����rC���3��Y�z�ɶ��ԛ{H����:�I䔙�%��$��H���lN�bt��C��A=���d-���䎑&�$Y�״��o�{	��6'�	��p�ģ��;��9%8O�:���ID'6�4��2�'��%$Ęt��͒:M��:�[�%�d�R'�"l{	�!1&8�4��D��8���<I�Yⶑ�Å�;i"x�z�DDxAׄH욂z$M��&�0NbL:S	�;䗰؜��H��'L�l�Fa8l��D�u"%):l�lL��c�Jm��D�����'p�Ј� ���I�'��`�)<$N	��	�"wi�tl�u���O")!�t���8�{�2�^���Y�_R$O$M���8oeؗ��Ɖ�:Bk4{BZ'm"bN�؛y"t�$þ:xJO�G�H����b9ډ�p�:�
���Ώ�z�vMa�ږ;��'s2�d2�z�<�D�|��w�z50����h9�ԣ5ӄ��D너܇�\7����r&��E�|C5�t����xY�j�8YZ���j�6��>;�пY�w����%U�JJ��ᅓfj�"#�TG<V`��Ĥ�p�6z�Q���#�TF����r�k�?O��jp�>>�����Ș{����':���\�;֧���k�:��pk�pG���Z��HܔC$������rr<��먘d�:;�L��4�7����bp�5�H#�Q:[!��%z�X���PFUDF�Qd6''�i�D������0�c�V']�N�q�TD�$:m��#���"t�C�3u/�wꈗ�	�Բ擢,��r��o*'J�SH�L86I�";$DRL8V�#��D�0��L��ɤ�u(Fr�#���{jQM$2D�����#2�'m��� �Ã��DGݨ��8C{�D{���n�0� ��N�ri:m�N�����DK�R�:��"A�x��L=s�ǳBW�H��l��rpy7ܑ&eD�Z����Ȟ;�Hx�M�5����Q� �Qt �j�Q�!L���2i8l��;B9(����!�C�I�n�8#Δ�|E�K/�x���P��N�ת#�<RCq���ӧ8ԲdB�������ܽ�HlA��,vf�=��d�����ji&��5aL��A8����QtÒa�:_F�58#IM%y'm��w�:���'N9S�<{[,�IF����q���8Q���7.ʍZf�����wq��s�7�ޣw-좻�+���UD[+�
�p�Y%�A���{e>�^�0�0��8%�'�����l{�{�{�~�?I��O��7N�uc�YO����y+�+ѩû��Y�i+����ek��pl�خ�\W3���͎���J�#&<*���\��8]�.5<s����㹧�ޖ���ߪf����${����}Z5}�Y:�Y�K�b�u��9�c��Yܐ�NI��[�c��*"fڙSӕ����}�����f���S�+Rd%N�u���0�'��Hp���q�^�M�F�/�}j�:��U3%ԝ�J�ID箧�sݨ�j\w}gӌ�L��7��������F�.�*=I��`�U�U�S������_yi�u����n.%>�jr����}$�M䓄�D���΢p����<�F�D��������7�ʡ��"ܭ'�RĶ�"u�H�r�l�����Ny��g�DG�+��5�e:����D}����5)m�D먈���}��O�"oە�-�L�JN��V����R'|��XpoҴ�epٷQ��"cr���P:f��K6ܤN����Xpw�ZA�D�nU�oe"Z�N�m�V��"m��N�+��u0�f��ND�2�Mt�rIE2Dn%rRx�T:�ʪ;U�Y����a�,��ʣz��'G�T���y�����ӒXԳr#R��#���'�ʜ�o^$8H �O��:Y\(�j�Z�D����JN���.�x�"'�%a̛�ę;F�7��>�G":��85�^�xLy+��窓c�N�n]S�9$ù ���H�N���~j��U�C�Y�(]LURa���2�� �5�#�u=��v>�fOT/�ק)��t�:f5zn9����T����{���o�[���gkf�y��B&H��%���	���U�Y�ڮ��FN�l��y5�.�����2K���y3s܎G'=9%�7S�<�����7�lޥ��q=�����)9�뺟�����|1T0����G��&`�P��+������|����wg����`<P�1R�t�C��[�y˜�h��(Y̆��54����XB6d�g�fS���!��1�n���8CL��o�K���T7SD
B�)F�e/wh�e�n�|�͙# !�i��2�3RM\B
p�	!�5�u#BJBaC����)
2H\s癧"�.p<��14�:i�i���i�Q�!>2}���8�
tX�����FS� 2��$�x�R��!rh�b4�!{����381��K���mQ�V',�Je4�!	���5�f��HQ����hR��L�{���< @S��R>isHЃ<Q����G1�F_R��Q������pt�҈ӛ�nA��2�c��(1�њD��!�'w=͝� �h�+Kv
p�H#�2k��4DA
�9ya�(�R�v�݋��h�"n������c���A�
3 �-gN^���'�3�2�eÈ_KM p��n���%��ѽ�Y���!Q��1�>�DR��/��EA�8T��\�C4��(iB�V�����;��M8"������˃�t�3G�#W!�HeJ2�#G�C��Ґ�)�?��Ҝ(��(���Fq�=�ىB2�tB4C�|�VS��D�&O�w�b� C4���44BN���P��E(21vŴb!��d��-\F��D�X6��0�Ϯw����DR�q񛦐e �"
t�V�˳/qr��1��nn�̈�gp�z�'Tѐdb�[��A�fD�ZRӅ4���<���3DQ�)B�,�te4�M4C4�������Μ �sY���Ap�!sf^w����������z7��v��k�ws����a#^]��؟�?#v�`��'�}N ^<���t|_o:R��[-t|x�*F��8����}�άpr��{���8���+��_�-ؘ���Sf��k�.kz�G�p�D����8��Z��!<�&�rL�pJ*>#������BZZƯ��vq8��x�|*C�\6=bl�Qe�������uf��D7������JGmYwMt��i4�D~���!UQ_Cj�F���wM�|�Zeb�8��y�ѷ�{N�d�AVo9!��{r�jTW�`ۈDh�ΔK��Y�̜�y�Gu�dL�+c7t�k�G�7����GWh~��Y��;�	��9��Nßi��w�{�|��w��H�F?����Mb���ZG�w9f����I�7M�M/�>�6�Y8Gg7���K/8_�V��G8�oCd��������<�A�ϭۥ"?�ҋ՛��M�.$A�7���r�kb�M7y��%���L[����p)f����C�'6��M]���A��Xoti[��P=��'�b�'v�I�}�Do�Ev���9�;J���(=:ཧ2�`�h�,߸_���Z+q.h)�u7�4�n�%�tҖ�[sP�wy�_E
Z����_=��>D{q��SM��ߙ^�}"Ӫ���>GWO�Կ!�w�):�S�F�z��ڄ�lY�
|Q��Hu���~��TcCK}F�Zl�\՞�e��El��=4�>5 ҭ�Jm��N�?w�|pl��}4�z�Zi+�p��>y�����B���3���r���n#��
td��9�{"�+��1vL��\z�ny9�p�����Ҫ��H���׳yӦ�o,����N�i�b'��;Nd��63�;$�k��<�g8.��!�A�ty�"�-&�%C��h��K�it'QN�"q�� �Z���ʉ1����;)�xA�!��]�/�闆�MI�o�&�K��c;ޜ-�?��DǠ�NL�͋��b���N!���Z4ߑ�t��}E�Ӿ���rj/���n(�'�wHv��e�d���lc$�]жȾ%Y��L�&r&��	�6?A���(�$wԇߙ)���ye�ǭ5���N��B��g�p]g�,�A��:N�N��7w:�VmY�6>#N�&�|�{��<�!���'s{j9�^c-�7��A��ZC|�#O���Q��5�",B���5!��Q,/4>PG.��u��x3�;��;0�(��+8Μ�_x�Kf����w����(2��^��穢H���-/y����/�9�;ބ�n�N��q��H�+�d�$F��^����p[ё#�!I�Lt+f���Z1�u�q�pì0�Dԃ\��|i5�\�7�;��>G�63\8-���M�骚U��3b9�A�y̗,�ǒ3���G�L�Yʊ�t��O��繛�͢�n��A��{'G�o�K��W�����:��I�o�w]�->�5g�snw�!���y��nm*Kx��Rn�8>2O���ډ�U���7k����U:A���C�=㊎Oے��3�iR7�>�g�œ�>�}���X��v�mE�S�{�|�m��N��[<�����K^.�!Y5���S�Mh�黧�_�zw�ΣS�GX���y�՞��6οۍ_��)+=����t~c��q�N���Q��1Z���vB���,�3f�e�I�;�Gg}���Zӝ�y����D���&/��B���Z:��>gq�BsG�Ixk��|#����Ť�V�#oI8N����:��9�~��)��9�1u̘���E��f�'! }�_�Vu-u6O#����]�h�Ҷ?-�o}��z��YJ����q�z��{Mzw�F͸�^j���C��5Х�Lo�۱gMËKيo�>�rb�f�Io�md{��VI���5ѸP���Q��g��W�zV�����⥱29���S��N���\8�6�I��Қ����{�F�%�r#\�=�':��nK�cH��͇#��:?|z�SI�_xг���hoMtn�9��[k�vˊM�],魑鿴�p{�s�S��}��zM�,e�/��Og{��I���<�	1Mgy�cγH[�>�È;[��������\/ԑ=�C�+�!u�*WHᮕ�]5�[�?B>e���8�s��7�H��ҹ�1�9s�m��Kq!�#�o�+ħ���ǋ�t�f�W��ܺq�g�#D���rt���9sY>co<��z����4�Α2�������K��=��in����~���|1�%ʹ�f�f;������q,�Y�����՝�"%����q��>�b������]T��*����m|8 �tu��wȽ���1��!��6�����EQ�Q>��
H7��!�VBؐ�OB����M
A��9�?M�΢w��$�����>�r/����׋��'���~����uH����~�����C���i�q�����_���Çf��-���8٨6��ÞxA�D>���W�y�m$$��^��;;�x�l��h|�n�%�w�����w�ݕ�J�Sc��W3[��D��$q?q�:&�ū"gd�}�|i�K��K<��Q�#�q�m����Ԯow�9���5�f�u�{Z�{$\B=���9�EC{��q����zu��gi纗��c�:c� =Z�d�K3=�mj�?vf�n���=��J5���k��ts4\ B6�A���~\�C˟sg';x_������[�uz}4��?��/���'S���,KS�����g{򆳽���_Q���r		"	�Y٭5�u�_.�k]OeI�ƞ��Q�n��k�sYj1�$EUD�d��:꩹�_2Y��h��jo��D�	 ؗӜ��Smb��A-�B�g.ʃĢ �.�۾K}\�U�ßz�}��8Os�۪U"���^s~���y��;�?Q=�Nڙ�����y]�:j���7��6g,�M��e�U#TQck�fX�$������ք
ȗ�6�lbڛ��p�������]�K�h��1�.�#�5�z��7-Cq�5z�a��k�&��n	di}���چo�{�$�E>窊�g�׎q�����I{�����W����m��;9����D��w��庹��!��nv&ݘ��,�3�O5qf�����ln�YP�(����:��7��·��-��Fc���a�j,�/d��"Z��+�O��ۼ���U���j���콳�8��9���om~z��o��"��I�>������9WީM�9�6��;�w�:�����7�ӵ�*��O{�Y_o=�3Q���Y�*"��=*Ē�	y�6��ݙ���,�\�>���s�i+�K��'��]���x?<�z��@��g���Uwm�"=}�����BK?h�N'ӧ�MU����:�3�,����b���7jRQ��������ˎ(!��)��#l{�曫D�Pj��۷VI��cr��M�WG-�*%-U��J��,�ę%j(��q�EFWT���UZ�I�c��-mYV;+-�Q�r�Y��v%�8�m}�Qp�B"QrUe��^.cDPm��T%�b�)H�dv�i �4�X�j��Qn=�m��ɩa�%��@�QWF�!^��y�6*۲�F�o`���eUK:��6�k\V6��ѶX�R}n�$�mRU&2����29��:8�ZWD^=J=�^VUr�+Ri�-�T�qQZVZ�PR�E�����8!9۹7��m�1l�ȁHX��;^�ۛP� �o)g��ӻ�tU��Q��`ڎ���(�6�k{-�a$�o4rJ�R&�ho&X��ｽK�ƾ�*w�wuI�Ku�����M�N�����s��]�Z�F���$%�eN�h��y�ɾH�d�!��RI4����T�8�.��jDV8�l�}����7�����;�D8h�q�[��o�U�|�R9iU�s=v������l8�֛�����b�Е���9�m�MMt-u�ly)rجm��lv�Y#|W{8q-�q*�UjYU�)j���Z����k�L�ǐ�8+F+-TJثhx���v� �YGmqKTE��(���]7�
&!�U�ΣE���I�8Q�̎42�l���*�"�HZ;Qj�IX$�bi(�B�"eL��ERPuU
�I�;�z�	���'$�CDS��ԍ���m��(!�9�*vb�4��뵢�NV�Z�X�~�W�	�T9UR/�^o�|�rZU$�^�E��!�(�g��W�{�HJ�Mpr���ӊ��8)]���\�������/yDKn44���p[&��'�+"��Tk���8���?����rU�!�Gg%?/�gS����ճ�T8�1_#wa�W��s��Ŵ�թ4��!PIՋ�҆�Y/)5X$�(��Im�4ǍD˞�ŭ=IW�q�"���Z�I!VG�$��j�R�8w������kG�ѱJGg/���ů�{����4�zJڶ�Y�����;q���sܽOڪj[*��Kjk���&>:�����lщvUP�2�VQb$iʓo-q$���Uc���$RϺ�4l���kb9�lt��!|�?s��.����n�U���Y�f��.r5�����wv71V�j��%m4wԉdF�,Nq��s�W=����t�>7jin��WB)=/�NmNتmX7)�du���&�#�Hz�N����7���v��_q�V4��*�����mq��S�����X&Wb��|����n�u�W�rk�D�s�QwwtQ�*�S�iE��Ó\BD��&VF�Ʈ2'�Īom��ۢ��ZL�,�$Hi"�-p�ϻ��ݚ�{
�P��~��(�^�������ס=�� @���Ə�(�F�� ������t���?5}��@��J\R��'��O��k���|���UګǪ��[Ux��U괪��UU�*��*��v��U��U\X��]����UW��Wj��]��V*���U\X������U�ڪ�Wj���V�U�+UJ����UU�UUTUUTU]�/[��@ 4UV����mL��ڷ�T-���y�Q��6Z�
���iikA�H��6�T�j+׳��WUU�*��iU^��Uz�mU���b��"�������W���ګ�iU_+J��UY�U\�U^*ګj�v��Uڪ�b��"����U\b���;UmU���R��U^����Wj��iU_+J��֋�&���q�Tm�aV�o�Yj"���M�,�Y66�5h�*��65��j�n��H
�\J��"c��;������U�U|������1UU�*��v��U�n�^+J��U|���U�U⭪�Uz�*��UUq���Zz�ת�Ux�j��[Uڪ�ZUWȪ�����W���>���Ux�j��]���v�ګ��{��aD�1T�,H [l��Z��%�X֋lm�5%�r�.JѮ��Ѳ���}_w���[UmU⴪���U|�UWUU�*�mU^��V�^,Uڮ'UUq���ZUW��U�W�Ҫ�X������U\b�J�i�mU�W����V�U�*��iW{������U\b���UU�Ҫ�sA&��V��Vc�[�]#F35q�yu͵h��xj����q���qq���U����t�V,�Q6]( TPD¢�$U��׏m�����qm���mqqɪ-�8��j�Z.5�|��~��o��[j�J��_��={����!�(���W���?�5���i����q��d�����1' ��"'O�"a�<tN�P�A6 �"C�lCf�Kb'N���`�p�0���`�'�ق���D�D��DD�<t�QblDN��'Y�	bpN,K!�D��D��,�B�B"pDL(E%�tK0�0�blJ �$A0B��f�J��f<x���&$��D���L��aBB �<x�ȺJ}�W������+��)F"1� �
"C���F��hB�Q����2EH"$d�%R��CSѐ2����E�!�~E6�LT��9��EJ1R"C�ǐA�Jб�Ұx����!"�$�)W��)D�CHPPd)H�8Ȳ vc�v��:���:XKJ2���A�F8"���h��
�����l��4B�1�����T�܉�(B��H�X1�ED2X��n�kD���G1����AccD�eDd���T1̔@�2�B2<�1�B���QSFE�l�yUB�X�YHTX�J��"��61R6hɚ!��Fj;�*^�(Bd(�\aFe)�:�f܏F4;�
�1��#�ۣ���W	�.f�F6J(A"K���0W-Ҏ���4������3iV��1#I�EH��V&(!ܓ��8�Z:�IG���D���Gq��iҌ�D,Fi�b7g$�UEUH�������E��868F�N�$��*یm�5nT��4X�N�Z�#d��2%�ǊQ�v' ��u�"��u�Tp�k)m}���r�P�4����x����'
u�'f���bK��	=��T�(�UVB��HD����V4�mYH*Ģ��Ur��ۺ��Q�i��tN�o��i��\���D\�A��ؤpo�J��uY%�jUEJ�",�CiPiR�)rK��N9H��lN�ړv�'�ջG	
���W95��s�~|����Un���F��*��"���Un��� �ib��b*���V��ߍh4ib��b*���V��߀�Qj,�����[K[ͼ�μӯ0�κ�6�{|��m"1�4�"�&�R�lC
A�(ȅJA���-&<�Z,�J\v}4W4ܧ4�(1�`�h2��cb�$ �o!D�:$Б�X!4��-F���H��bb���Od&�k�*J,kTTjŵ�D"H��G

E1�Q%%�*q�s��*�Jn��P�c�f��3DL��Il�	�&�1,H�ȢQ�D����0��ʁ���
��X�����ݏ�W)���
@щ�+�fݸ?/����N����T��W�tgבd�]����ɢ���UM�bB&{ި������C��)���`��&!)��c���j�]tt����[��G�o^m��!�$[n�iI�&���d�M�uu��~"|tDL��	���g씔�dq�}ԒI�|Ou��e�ٓN�ӫ($,�����OGF�y��J�Q�̚�m������!�!v
����L��D�豁���+����*�F��o�%�X����?BQ"�fnŬ"F�)������r��\����ܦ��Y�hi�8x����˃�Z0(�a�� Y��N�]�`l�|l�������a�8B�b��/�D-�n̂1�n�C-I$�2�>���\����@l/I>v��,6�h m�>�a��t��5��d��a�.��'͉�G"7 djBbZ���2��QA�B�p�?Y�fB�O͠n	��͙�'#y���D�P21��a�cnM�G�1������,Q��ƛ�\:�0�˹�ʩw�j8��ΈIJ�h0��
�<RC�<||pDL��	���f�x�Ww��o�y+o�$�C3X��7:3�:e���y�li���h��6|���D3ieZ����F@�$�Cj��(1Q6ɗ.x��� �?~\$0�Ũd�r��-�WCtYޫ��Z���#���f����J����"�"����T
g�sHΜ�i�3��^s83Q]��h�˜2��E4���O�N���Y�Q�0�:l�M�GDe\�Ƈƌ�P�8&TFRC�8�Ŭ��*Z���c�r��B�3S)�G ��2Hp��
>��A��#�)Z��ᮌx��!,�ȂD�ҹ�8"eY�uw]�crI�V�cN��$J�C��(=IU��^s9�G��%]bƈ�vzzj9ƆE���I"B���&�B:!�o4X�&��I�B�!%	�\z��C���L]h0��E|�Óm���I�{R�fT��U&�<����fJ���#E�I2��v�������Yc%_��k?��"�A�c�>9F�j�I��4�p� e��+wX�h���g�ʭ�h*}�#)��5!����G�7s���[����M���SֶY8lM�g�>:"&	�t:|x���!��C�gےݔK�x��IVtN�I$��p��vs���Ô3+�^��@�ꃐ�_g�R)2��Ѳj���$T��O�z���U^���@��Ct�C!A�.h�,��LBV�˓(��%J����NYL�<a�~�����p�C���A]*M'#�u)�#���$����e�rWa���	��|D��0x9K�!�͘l�b`��:ӄ<y�.�Hx�g9t��JI:�.�t�����eM�a��i��~�6<��Jd�Zp�h䒥�N֏�
�]2ɧ]D��|�x��c�s!\����+���yw��@Q`��HXt�oTH�x�F��8D��˪v�T�}1�єd�%fH�Ƥ��*6��ɸ8t,�Ev�^ƶh>v��e���JK��h�Y�6|Y��:ӄ��^ϐ�+-��DL�(�bUrI$���a�����rv��o�Ǎ:іjÄM��Tx��K�Ho�q�J1;U�VPTCERY�8w��ߺ~�^9�f�U�A!�8FB`d�/�gq��d6d�R��)l8�}clx<u 68�>h��i�m�f|nN|;hs�#���T*R�2i�FU�����Z��Q�,�gL<��y�^u��<��l�e���J~��B@b(�X���.q��,��"\�4E���;x{���r�Y�!1�U���D5���
�eH(&2�'�&{9�na����3���M;uĘ݃��Hku[TFЕ�"��Q$�I$���EI��qf��Z#QI 8VM�ucm1��)���I1aq�ƈVMS��馹&æ0�p\�ao2т�lF�e���X!'�Lf�#Cn��f5�K���c!��7:f�xI$nh0Ft�$ YNm5�ɷ%Ut24h~�NC<���?ć^<x�"�%T�b��ŗ�b%�,�ƪ��Öǐ�><�rd����8g�F���:"&	�t<&C�M��gH�%]_�4��՛wn��c��$!jK5��I$�%�Rj�!��d��<;h6Q$p̚v��w5E4U;L�F�F@:tpND��&���a��$�)ڕ�����ګ�`h��ά�^M��CFi����h�+�$�T�"��U�E�+
�|�D=	/宾���7�Y2|c/t�ÃnJ�ogĦIUA��7����&��W��Wkd,���xО&�h�ɷ��$��K3�6�e�KK^'ͥ����Ķ"ZZ[,Z�-���N�Zy��wmo�[]G�{\^\e����<��/h��<O�
&�x�#�L(��V��~F�L�KGï1i^F^ao0��G��ah�Zy�ٶ��|�N-�8KKO2ŭ�m�E�����c	Ű�E��LZi--&ش�[�Z-8�O�g�D�+��h�'�Dp'��r�z�������K%�����'��������y��I���xvOd�ș<Ŀ�ܕ��x�D�<9rww$�&�'�w���F�FR�Re�J��Zq*-��t�&	I�7�:D��T��|W�l�kĶ6�-:�Ih�Z[�-�I�ò!rxa�T<hS̛�T�d]I.J��q��0����Ź?~��J��ݢ���>�����g,8��^NFx�ݗ����R��9����z��������we	]��<�nr.�=w��$�!�Z{JϤ�����c�"���#���ݎ�HK�/��{���c������=T�������p�#�s�]�C�^���d�l���~�{���>�Ù�ɏVpW;�w��9���x/������{�*��w���M k2ffw3���UE]�{~Ѡ32�33>�>>���Uw���5�3+33>��|}��}��|��������Q�Yu�Zukm�u�^m�Z�yi�e��'r�kL����A+���r��f�XuS���.���duP�M�����D4El��}݇&��r�ڛ8D���7���BHM�a��0 ����ZO}]�3�VUg�ǹ�i���!A#�����n��8�8Z7���m[q�䴓.��'Lg��afs��l!g��48�c�A� xa�4@�\)�[v�":Z3��O�GD�i\�;8=KI	�p�B:YiQ�4p�cU�2(\H�}� �A�1��z����`�ڏQ�*	��>m�A�*��`�����XX`"��ʕ`�ð��!���y����u�\u��-��\�����S�9�K�pF��$�c���QQPHQ��D�_t>*��B�� P�r[aІ6��HJ]�U�S�S�� ��b��<��>�J<���4H1Q1D��R�
293tH�!	*5�01��t2�����,Ԅ��a����(,�<b�h���3�ĒX�l�e�I�$�[i<p��7Q�-�vA4��ѥ�CLK�s|�pac����|1% ^�6����jU�WC�����:z2��i8�=����G�<d퉂��N�O���$Z�b@8A6����!cCg`i F�%0S���"lM�f�DD�0O�D�<M_wBTw��{��8S�ň����4�pA��y2;8�t�h�sv&-@ʮL^؆�]�¾<[�E��Q� �)KI�xL����T6!�q��]Q"���X(���>�o�'�b�i�ڪT,�wMiD�B��#�QI�mRĞ&����R$�K&�ʹi����S`�E<oX���$�P�f� -ȗ�*,Т%�(���p����oL��m�h�x@x�1V�����ʹ�S�
���bq��%��|��@�D���(�=!b���)�
�L'Ĕၖ�$�hb��@�Q�En+t��=D�A�=H��=�`��%RPA!C:1�鴢U��r[ z�a���Z8I"R��}��O����X@����(!O�(J�LYA�����j
4�p�.n0�1��g��. ``Q�/�l\0�SOF�<��9���g��)��|U���y�^u�<��a�\F�#���Y�5z4�8"���DԄ(hp;���Y���W�T��|�*���D�E2b��m�t�����xa���ba�a����p�m4nF�x�("0R�t�LL�}Jm�KD%HR�RH.̅�2�/A@h�(P��"'�(p��	�R%z�A�H2��	�I��Qt��e��YeM]���l�� �x?X�|��!	H��J쁐�j��6R==�UT��]��h������Z-�P�(����r��C���шC�*�6�E, $"X��d������ϙ~eoϖ���<�<x>(���pt�{���a�:5��w�TTT J����	N�a�Ľ�W�>b|Y#4ե��%���&b`b��Ð�t�3���j*1_���d��=��Q01H��P���b��J�A�%����B)�����g۔Yu���m���&$�
:AR̠���-J�E�G�(�$ޙp�,���D�;��P�:�:b���M��tm�
u��	�+����6K�u�ބ>9I�#D\��]�!r�wE��C�ČGbA�1� �$�� �G%uR�<`j���鋦aӲ��#��䁁�C�|B�7������HRS�����<C�ˬ������m�u�q�κ�!C������;zt\:#�����ֳ3)���"JB��J9�;��[�x����J�*SP��Y�V�#*�/�Ja����E��;!)Ax6���@d@�� ���Htd8A�	"8�啋�%��dh��F�FG����n!��!h̜D��xyL��ϧL�CNh�L���uR��)��ы
>|�<0�@vh�8�$��+L����я&'l���Zpqtř�b��D�sz���M���l����7"A�9�(���S�V��� �a��8���FCd����tz�L�5[0�'�Uj�����*�ح�4��m�R������H/FGe���y���yמy�C���|p���.�hF���J%D���"X1�D$�T��,򨔂ĲkB1�vK	�ҋFC�HӆB2TN��2�;.1��7�Gʈ�9y���$�i�"I�YcR�Sb��&iX� �VZHEmD��q���������@ѳta{��!��l�2Ǵf��1�ɩ��0�a��!�)�c(32��봒X��ҧ�_kl�J����-��؇,h6@���R��P�w��OF�*�y	<@�w��Ta��bu��c:�����bA!l��l<����D�/��i���� ��X({�"+H�{ͨp�on;/
a�u�<�a=���;b�z!}$��k�V��;h��a	T����!�}g�Cw���L��(�q$�TD
$W�Al��F
�<++S@�%9I$.�^4IB�!�D�\���A�"%e���TKa�ӌ�!vSD(����b�+#>t=x�(l,���0��'��舘"'�	><'�+|:IjL�ph��.��B�Prͧ�"����$���,���B�`Ã�^��Nd=�%�$E�;��Y����[pӺ5AD��;��u�����>���F޹��[1!'��Ө������O�O9�H�XV�W�W��3ixd�ն<r06`B��!P�F6H~+���*PR��Wd���MT�L���p�š��J�;lr������l�IR�͌4Az{�ĘN(2@���!��et��(u �8�Ϛr6��!�ş0N���0DOa�F9�!�!~:��_*r��eU���;�n��������4�;&J�68o��>͆xl�m����d��ԉ28`{��Ca�z�A�;laC�/���m-�(�`����Dy&	AUIe+�X����U�=��rف� �(h|h�C�1M+���Y��x�5�=&F�!"�����:f�&b�!�Ha��!0>h8�l7A��8Ak?>�t��r������WZV��!�C�ω{V�h2�t��9G��U�~<b�0�UAVÕ�@�`HAU��ǰm��?+D�v��|�-�[e��?â"`��<$0�{NI'����hZ�:5�K�{'+y��2�%�A�.!�ٍy�("g9���������	_�YYZ}W�$�Cf�ԧʹi_�V�ix2��)�Cx���G�bh�ӓ�Cж�[mD�e�X�2;YlI�"Є��� v�SV_2��D��wQ�h<A��	�F(�3����H;���a��Lz68S#�!�a���
\�$�%�v�`��C�����Sdr6�¥p=X�h�A������\"��ܱ���-�	
C�wׄ�d!	*��#�F���l�s����|L��b��t��mْ�D�LU�(�U�Kb��?0�O��%�ext#�g������t��1iť���lZmlZ[ؒ��io1V����ɴ�ZDh��%Ԓ�",�H��a��Z0�E��m0im2��)�+����Ɋ��G�q��QkbҼ�y����ai�[�-��O�o�~Ke�mD�4��O�i�Vͥ�ť����n
O�I�RK<0��m���8+E���ɵ�V��lq�%��Zm8��G��u"ش�+f��Ӌan��%���kb�+b��b����ir|�][-��o6��X|�M�7$�0�-��cO�셓Ēx�Ļ�w="\s�8]˺2��i�B�)iĉiV�o�u�N1�^f�I�����--��[�[��$��Z-��������%�.��9�OA�.�ZDm%~#)ygfd�1fX���Q ��4��!�Ȏ�Cf����,4GkDf�4�a�xA�C"b���3��!�RzLу)F�i�T�F��sB<�x�B �A�ڠ@��ТLF� e�C��yYDR��B�c�Rb�(��2`NB�dE���N�k/6�p�����4IOHw�}�Q���}gy�H��ke��&Z&j۴Az���>^Bj�!H�)�����5�YnT3����Z�nJ�-|5�*�dM�����m$��*U�Iם�!S��)�6]�/>Mb�&'��7�Š�'��%! ��A]��r�CF�<ψ\��-h��f�!���	߇\K�p:�yl�1�i	�s���4���T�,Z2�Zx��u�{h�)����p�Ә��a�x��)�$��p�6�����O�ˠ���q��Ψ;)�7"�g�h��D_��^@i�cY��$" 	��ٟN,�8p��"�s�8��78�ԻN��[��<�(�����+�(�cb�*���|��r�GM�}.h\�)�ҏ'�?��䎩=�|�������'ް���r/#U����OW��u����i�y�z����ή����^w��y�Ê��[�51_/�������v9i|��7�Vs������ۙ����r
F|ｿ]�S�}��{��q%�o�޼k�����;�$�{�Zm'Ѫ�y�7�Q}��t�
���q�-�
;-r����EA�+*�V���	;]����zT��v���1e����jʝ*ed��$Z�o]s�T{�Ԣ��cv�B��B�L|md9-�,�X-Qq�Į������"��+*�Y+S�W�����o8�\����v�m;�(�Pu�7�+��˗�Evkm2�s�t��Ņv4J��z�;��&A�M����!k�j�H��}�+h��ϧ4�U�Q���N֤�E�L����Ȼ������N;��n��]��H��#��Mm�|�?�~yg�}��}��®���k3+33>��������w���FfVff}��*�}����}��������f}�V*���}wy�s|)Ӯ����.��km�u�qǑ�QŸ��6��Ͱh�*h��H�RfP�E��?j!��`���m�1�zV�.'Z��tQCaH�bv�!�h�H\)���.!'�%A�I����b5R���uD�R9$����ΩK�D�*I4:�X��D��GԠ�LUUG*D�t�BY�t�1�6�h�Nd:C ��m8�R�e)�ʲR�����#���!M�r@� �E<4I,8�ޢ�����;K����0x��p�6����F
TԬ����H�diV���`��wV�,��m���Ɛ�A�<�c囫VU�����|�u��Q�.�.�mlk#AgB�lM�?7Ee!�l9
�	Q�pr:�����$@۷�
�E�.<�@Ea��M?�#�8+k��!	)[m�mU%S)aQZ���F�	Q�Z�V�q��;0y��W��@��1E�%�q���13]|�����Q�[.<�Oâ"`��<$0�><|>�>-�s�'7�N�1�c :��k���'��	�=U�5����o�d0{��
��]˹���S��i�)AD�8I_2Xgm��e%���HB�XN��c��<>�6�����)����˥����h?�� %:080M8Hl,uCaa��h���0U�FB���#E�2ۂS���Ɲ�40m�#!�y��*h)��G0wA��o�i��'J�V��:�0�6��VbLV�X4G���7_�!��	6��@�b	,İ�P�C9��MXe���!���x��6��:��8�����jۘvph�*,�멈UTABY�I�k�>�c�@8VP��ˇT���)2z|B0!*��DC��Fp���6�p�jxS�3֡+Ų:%Ue��D�Ü��`��7��07�u���"q��n�yƩ�e9���9�k�a����T�"����Y@Tjd��yǭ�[�#�j�l�$\C%�$*Sa�:�@)�t8���k���m���`��@��#a��������� 0s���^�<2v����K�9�0ѡ�a��T��|F_"�el�o�~mo<��<�#���q�����)��`�&�_c�1��WB�μ)�Q�J�������,�����	���li�}Ԓ̟G�Hy?.���Q�ac�\�x���Y��KRm�8��c����|IfLRh#A��1Ǌ>t@�D��<eZ9�6�j)���b���銥��H4�]�XAm�p0��4�x6�|8�L�S�0��!�0�p�E6�Ǫ��G
$�n�	��m�v��Im5cD2�(4@��V;���0h����)�4݅.�p�|�Jhc�-�(v678i`�0�l����oͭ�y�q���׉Ё��d����a���1�1ҔC*+�Xѐ�HH�H�Sc�P4�i��T�"y�it�f���q��B���rX!�N5��`�H3����b����m�	HԝQ^�Qv�iH91��:�%C�%D�S��m�]U,ic�5����H�Lc�HY�47���c"$DB �V!��ţ��ȳq��!���3%˺��x��x�����Y�WOeR��c���� �§�����7v-����2E @(a��i���^!	��ZG�TCZ�2t�r��0�UylKDљ$$��a9�0F8c���}��# `u���b`i�!��m�X `ܥ�IO�9vi���F��n��j�����ؖ)�@�x<0��Y�鰏�Ѕ�����`|@��m!	H�RBږ�L!vIf=��bй�\��&�<��Է0Go_�äAA�d1�� �1�I�'���G���i1x(�F�p���N�4|"`��<$0�><I����z�I\{�Z��c�B���J�J����m~ �X����:v��Bp�@e��\:�Z0s����&�����"Z=<s7D%U]T.�/H����P����6�hrFE�����h�+%4thj��Hp���H�X�����
BJ�(�4<t�q�������A����9u]Dd6&X�Z헠�4b��l�1�������8�-R:�B��䀛H�<l��a�oV������<�P&��!A韽�ᡠ����h��`5���z�Jn�e�e�u��uo����yמ|t�������`ǖ+�a���
�y�̵�ԟF1�c 4��Qp��ѨOF���5Hl��ОK ��r0�����F���@�A01cy�G�������|��[w,��2B[0�������-�4gd=�.�H�.�"����,4�';9w��Y�	C�����8ǧd��|�>PAV��nj���i�os��0,��#���%\��0���L� ڄ6ڤ1Y��Vk��8<cOƙ:A�2@�#n���el�����u���>���t{c�C���W!��.�5e�ڪ�*�N2���:˯ϖ���x�<xHa�<n��n���IEL�ѱMV�%���_'�SM4�M�	I��c��$�)�
r��%�9)�P�����5�i��$s��B,E�9��)h�0U���T�"�І�PbNa�cQ=c�"v�5��bڱ<���R�`�0t��:�<$ uH�#22�F��ϳJt���� 80�U�������h'�@��|�7o�V�Ч+�Hi��7$�%-�&bhp4��6�td�(zj�A�0@��v����t��!aE\�xvI��y1`|@ӥ�BwM�t1.Z�a�&�y���6��<�2��Ӭ����ͭo:��8�����n��!�&Q�b�.2��c.<n��C�����L�)AE�װ$c4�E�dEC4���h�F��M��6lF��؄���e�u=�9�*�(V!���Ediĉc�T���ېiؠ�I ��3��c�H4l���72Ao?XAp�-
�h�F��7N̨Z���,�(!%1���_q
��q�M�j�^qa��_1�H�ю�� h`Y;
vŶ4oa����;xI$v6 QO��A������S���%j�J�WX$���Ԡ��I�-�?1��Id���F���G(|�� ���zڪ1��י���:�=� I@�}F�˗
�0��.`t�o�6�Rкe2=`h��'�6y��!q�MŰ���I����2$�
4����0r��>g��6D��8vP���r��駃e=���J�U�yim?4��??6����Oavl"Hr�W&�B�8[��&J��.Ѷ��kv)�\ \�+/5��F1�c 0�.�+|���t˰�2hz>h��V���������D��S�h����4⧣����ѦT_V O5�	%z��Ca���7c�KN` p~v�r22�~�Ja��U��d_��*Ɲ:h7�p@���H[��tA���Q�G�AB��8��lv�����1E)a�*�׻�y�06�k��ԦK����&�ƞE��?J(邮���8�I�0�	M��*�T�q��-L�}�ipAڄC~j���Ӑ�����$�f�)�$��	_!�il4�J��-�ɤ�����[l|��%�2ش�۬Z[X���%�[�L��KF�ť�g�:O�D�$kg�d4K'�X��;	wwK����˹���M"�b���|�%�V��E�i��?%y��^a�-?$[����E��Ǒh��ylZym<�S���f"��S+bӭ�iiii��ZD���Z-�[�M��E�ŧ��-�I6�*�r[n��d��&ɲx髑�t��+Ɗ��O�in��O$K|��b��+b��[6��E��lm�[����i�؟	�x��'�d<X׋dH����w$�%�K���\s�,ZU�ela4�L���l1V�M���χ�p�|Og��ƅ<><�[+N&�ť��x��io1W�0����w����;	w�'����2���s��8�I1^y�������7���wr\��#1<׽3�������8u)�=�f�o�����g^�w$�{ͫM|���[��Ny��s��yo��5n�{~�>���_���Z�h�)#��}~iq�j��C��j>Y�k\���~|���&v�3�}?"�[�3+�O��
�緟c��U�U|�}��o{�����f}�U�U|���]�sFff�3>��Ҫ�X�ܻ�������}�iU_,W�]��֌0�afa��[k[μ��8�:�8�Q�L0 �I��c�ID+���@��c���W��=+��ܯK�ߌ�_)!��Y5u0��5br��(x�ݙd�:�2�l]�M��B�1���ah|�YB���Ɵ��Ac�c(�x���Gc�Q�q1�����L(��Bؙ2�X��[lX!c�@�A,#���2�0�&�#�Li��Jf(��m�[ SD���-�F�i~h~�# # �|4�G��axF��٢2S���գÿQ�U��+� �$\�4ㆪ��J��r�Ep��>iƜiվ[�k[μ��8�:�8��5��X�9.[v��Lʕ*T�P(��-�w��|l�2�A˚g�������i��E�%x�!0i�����R�^�CgaL41�Z����h�B�$N*:� ��Q����B���,f,�#��i���$��X;|�Ṁ0C�D-��D�K|Y�Kuw��;�abB'F8�F��l!����`�pǎ=``�.>{ƌ��O;m�B0<o�'��p=�O��HX���v�����Z1����T��cR��s�f]/X$!�Ԇ<�8��b}�P���1���2!�F�}G&%顃!Ў�>`d�����y�|�ti��i���c��C{��Y����4���O�??6����<�#���k�q2ɣHD	1��A��J\��p`�Q�C�\\\�|Z:uv�!�,����	<��揆��!q��.#tz��8"����(�D��mf�����R|�Ѧi�Kp�
!0Q�"��RE�H�)S�9�X�N�H)U�AWM�V�r���)+�ċ&���2�c��ce�e�%�?Y���EEEhHB�Yޓ9rb�ak�`�V�,Dj��M�:���(m���;���y�Lb쁈&2@���; t�MQ�68~`p�d9􄘅E��Kh!Ճ�� @�r1�����t;z4C�'�E�T�l�"�.F;��A벆k����P��|ل `��|Ӓ0�e�4�����6��9��n�T�po���gR���B�8C�<i��^Xƌ��p0��j�$4��'�ZX�X��1�丢^8��d�)�u�J�_�x�n,���P�t�C"�1b5�Í=� [�'HI*����<O�m�����C����m��m��ŭn���8�:�8�nhd�m�TTV���Gk��LA��m�)!�0���LU���Vz�Wx��G�C��'S�(�B �
�%1ZW~J$
p��`z���0||sx�M8�����\���
h�:ԨQ>e�M����"�������u��?3�<hx�CO��cc�uKDL@�4ϖgqF�"m�C��b�sJs`B�0�'�Č�r�P� ��	PL�B03��a��c����J��%"">�M+,�;u��aӁ���f�p�g�:u���Z���<�#���|�Y"&�qÃ.�se�8Ȉf:W'������А3�<�WR�������=PQ�`�4�1!�:h�e������1���*�Ӡ����w� A��6�I�mXW��x�Z�����J�!?h�"?%�ED�:�!#���v!A��%��@{�y>�����|l!x�|4'\�~NJ����uA����c�`d��tݭI[A��5��Ad���r��u�rI&�CH�Ũ��8f4C���#!C�����������">�|�c�Z;&���N�|��%&�>|�Ͳ�-�?6��Z�[�8���㙯a׵5(}ւ�&�ޢ���$T+ǥT�X���؛!��i�փn��ɜi��;��#��BB�r�
h���Kq[`�Q%���&&n��^e\�f�i_?5&��y�%�$d!�<,`h��%�a�7���h�c�hJ!_1��P:�h������X�2B�]|6>2YL$%@�a>`p�H�I�6�����h`�ybQar��������UAc��Z��#C��BO��%�+Uڪʘ#-#Ͳ�/��o��-kuo<�#���4��N6�E��a!s�܂)�s�t�m�b��x�d�-�f�T+�W��[Q�Ǩ�y�#^n!���B�ֆB�[�����u�vV�8�I649��$e���[D��=�R5	�3[%$VOόm������f�,&8�epd�,���K�t��J1�ck0�9����a���h6B�!��&*���M�e<���(�̴=`]}%�C����p�vh�4�
h�3���x4&HF9qe�XW}�g!���0D�Ip�a�t0!����C��!A��l8ο00@5vCp��UL����M�4C/IǸ#����&[��7&b�ӟ�RR"	YR%
P�Hحc*�X�uGb�b� ���]K@�$�0�T|�̲X��/�R�\��u�;���U+&�&��>:�l?-�|�����Z�[�8��x�����7����@K����$������k��TTV���q�pR�q$�V!a����T#D�����W-�dE�� M+��(ڟ<�!��p�`xo�n$<�2���B�������堄0�Cc��4��zB�-�U6�I'��l��O����B�����b��|LyT$&"d"#Ƀ!�Q�ZD�� Ą	Rj�*��]V}��>��d�D�'�I����c�#�iC༛�2�p�u��jfR���IN��a�BE
^�Ȓ,H��U���0���Y|��yn-kun�8p���p�j��	$��~�EEEhH|W�ʣ
ºcY����OT~I���Ёd3L70���;�ˀ�T9t6�� �~F�A�`��JÀa���Nìp0|��������$�a� ¦�K��.'�Pc��"�H�$�� [!I1�GɈ���"9�3���S �E�6;V��-C��BCP.1o���c�&�B��y>h60p��d�@�0Q�	TA��a������Q�H����:�$ƒ6�#BL��rn8L��968m�����e�x���̟��G��8��ռ�qy��O&�J��PF�I"5Uv@ԙQ�q��Zf�:�\�,߹�**+BC�
J��z�cbݷ� �ς|T���CL<6i���j8M�����k�h��� �e5�eT��%-�Eke�,���pv;w������p2��d8l,>2�Scx,v	:}��WE���m4�,� 9/1�o�t6M6!�"��PA��܅���4&�a�ن��C.
@��}�,���kI�	*류G��%TN�&GZr�6�XD~r�����D�r��a�
k���		"`�M�����Ҧ0���b$��i
~�VSi2�%<�<�O�W�h���ɧ�H�u�-"��[7��f���b׉�[-�-��[��KN���h��Z�%���&7%����)dY"]7x]Ļ��'q.�ܻ:��M1r|�j�h���m��Zq-+�b��+���m-�0�[O%��iձ�ZylW�żż�α��,��:��b�m�ikbө����[[���������~a��?'Q�䭭��ܖ�Ka��Zm>Ki�ìq-�-4�[���:�-:O����<Oۑ�����I�-+�b�c��-���#M���8O�����Yg�!?I�H=��%���\M�{I{\�w+��D�lU�Qh�[-o���=N���k��[--��[��KKq��ilyl-x��a�&7%��4�K"Ȳ-$�id]I:�FQ�"LKW{#8d�FZM`�FL �[H"�h�l��D	:�P{���"D"�!@��G��S�؅raCiVA�D!
���cɜl(1�Xi�3M&R�� ����@���H0C�)?�8M=%�Re���B�(�GE �"2;��K)�����T�Z��[2�7o��ķ'�u��\ńڱd'�E�ŗ#-p��8s-~���!�2�\>o�{��=�0}\v��.w9%���)h��t��r�����!!�xo:!�����E]����H�F2L���B;�S9�C�CK�18CދsI�*�aGA\AG�!Q��RN��5��*B����z���$}�����iFɕZˈ�ύ����ܝ�h�Ӝe!���=������pA�J,������	��{�#sK�d�lWn����)�(��ܞӚ^E&pC)kBh��L��:!�Z�h/93y�{Ê>��Ż�Q�h�t8y�ɽ�S��:BD+}��T�F�����h�D�8A<� �~�����$v��lg5����^qO�}=w�����\�$�r��}�������C||����a����Y��_���/y��g3"�#3���w�>��b$��B*�B�W鱦��l�rIa+�J��u�T�����U���pD�V�t��I�$�-u�i$F�%����ZXڴC�4�M8��q&X��$�udY+��a!�u��[e����R&�ՈQ�"&�U�%E����aX�h��dRR�D�^������AT�[,Q"��g9�]k�q9$��f*�M=�"�"�*�B���I�ܫZ}۶i#�BEnbr)޺���N���D[$ډGlc^�7[�&;l�Pڢ{o%9W
��G������qZUW��˻��32�3︫�U��o����̼���*�Uz�-�˿�333��}j�U^�^���j�N�u�u�Yu�[Z�Z���y�8��u��D4�EʉE�V�@��$RA��*62�&9 ꣙VR"�Lt��B*tB�1'�D��l���%��ʚCTY`�X��
J��$8�eK]-VWk�-RQ��*EcvȊ��#�;J�Y!�b**+BB�	�\��J1�)r5Iq�B"�� +�r���t��I��y�?�sUN>�W[��D������R�^�g-G�%�(�t��2�3���4j��J���}X�5_�>����B[��<jH�?�M�5�.�U���lt��0���d��N�W�r���U��Dl�a�;��0����X��p�����HC���d�̚�4�� ��a)r;nޘ�}�!�΅����;|���>�����I
��C��2Ï4�+m������O�O!�e>f�ɷ�g0�������s�l���ZEEEhHt����ߩu{N����C�4��G�8C�M�J��:Kr��˯����h�l�R	_��BG�\%W�!�N�~���N���4Hɶ���pٶx��81��R��hE!1��$���іEr84�D�nw�)�����2}�Q�YCaz�e�RL�;�|�!�ǃ�֞�ď_<~밄6 _Xd�upi2�7��~t0ql���q�[y�帵���C�Dp��'��J�l���e	�A�ƨRs��'�����	
c���;�d�4z��g#����	�%u�p`q�(p�2��7�*���+�ꊟ��^��kfJ�E���z:c��N�
!y��2��*$ZL��CH����[D�2"ĜN��M�bI����x6�Hd0B�����Uj+��^�V���3 H}_��=���0Cד͑���ƴ��!@�4�g�sr��l�ԄI�B:�o>h2��R���v���0a�,?6ӌ�ۭ���ַ���8q�m=�"|cɌ�ji�^I��**+BC�a(>:C�*��W��I'կ����h���Y$�?8���a�G��Nl�:�^!��P�����d*��c���&]��z?8�g���IO����{���a�n�UC]p�%e�Cd43��9��)�A�^`'ɀ�S��y=e]\��Ŝt���68}�*��?k#1���
,t���)-���i������Z���=wu*-���	,�v�ZV��ݷ:�d4�4��i��Ϳ-ŭo-�p�� u|h<x���Η�Pb)D,�Ɍ���ۃ�L�#"i�*)+��Ѷ�� �*Dy���Z�V�R���E�E�A���
CG �"1�u2�2�l��(��:p����W\���e�"��K�6�mQ&U�+,-U�*��.�fa����7s�QQQZ�6j0��F����b�Db>���n\t5a�lu���4Ta1E5T�p~`�BEp���2����aDN�[U�G��ܩ�ճ��RD�yK�?������r�>ú=&�h-��ܱ4����uKr=z�C+O�$��ç!���x�4Y�X`�A[��L���aJ���\#5F�d����n���I����&��!(��K���*lUz$�Y��b�h�YF�q�����ߟ�Z���y�8���kaI�^>EEEhHL�J�x�a��h�Y��'prPT��wE�!$g�����kD2��B�}��5��W���YA�~�0��yc��K��I��ӆ�C���F[��
z^�v�Pdd\��s8E)��Bj�Xh�\q��d�WYZ��F���8�Y,㧮�"����dzmރC��uW.�ã�cA�1#,M�	$�}��`�cX���WE���{_.+�Cn"�y�����[�[�><x<x�N�h����|���;vd���"���$��VVQ�|I\HM���]�t��pt8��px������9EK)���\4<�c�oÀ�=v�ч��'�!d8}P��i	���Q�,��FʋB�������9-)O,�I�����!���ѶL�:���9l6��$<�$�0�<trPQ{[��,�&]��NG.�����Ѳm�.���i�Kh�4־�~Vr`ۈ��4�N��~Kqk[�?:t:tGN���#o^`��m(���6���Аh�ʺ�\"H~0�+���]k���F0�F�̖g� �s���D
qتou2�[)D��Y�i6�v�RTؤCnI��biєh���,Y�|���C��Q�S�I:u%���P��cA�z<��J��Y�:�y4<R�IU���C��^l*�k�)պpx2o���H�z�󺽡rk��*up6lzҙ|>2!��$dv9�W��+յh�_#�>iƜ~m��������F��̷�S	&q���	��e$�\BEIP�jJE$ev$�%���+	Z����|�ш��HQ+�"�tTP�c�!�f�)�ݹ`�c�5d �l�!�B^l̃�%���B��mY�$d� �{kp���,��R']���4�k�Z**+BCEl��jl���t�u���3�����@x��������2��<<pC�Sѷ�O�p�$�C�.ko�$2>`rXHk�FC/ñ��[k�8tzB�]C����e�	BBBcŢ0��[EφJ��ǦB�g�9
��4ûJ8s/h�6<���m$~!Ot�N����4!�M����s���_�d�M��%�4�x;a4:�X4==#$$��̩W�|Q"$07R�_�*"��dm h�x���T�|���N��O<�ۏ�-kyky�Gn�C���&����V�ȈT�1I�*�'x����1+/�Y��H���	��+eee?p"dv��Ī�.���#�ؐ� Vj�44L��O��B��ex��պ�t�!`�IذXV��,����/f!��m��r9�����N�����}�&�B�d"DH2�*��������J(�j�PB�!�d�M��v؇��p��YX�a�+���J������%)�ѱ���	����D<��:*N�)�e��C4d��2Y��??6~ � ���'��"A,DC�&����e �ADJ+$KbX�N��xO	�`�	f	�X�&	�&	���,A�	blN�D�H"lD���A:,�pD�6%�f��P�� �""xD�H'N�m�強.N���|��|�y���)$A�Q� �
�<��y���V뎺뎭n2� ��"'DL�"aӇᲄAC�	G��7���"���=��_׸����5>G5s}��{}����趡�~Y��Q��Ψ���7|�us���n�V�ïw�칒�}���a��yf�|�ۻd�������l��w���Y����N	|�����~�����4�<�9W���>�s۴|�8]���=W��S��������/z^�[b�:Y|J��D�+ݶ���ώ�&ƾ�\�k�	T��_u���Aw�w���6J��ɯw��}��|��W�Uڪ�Z[����ffg3>��v��V��뿷����Ͼ�V�^+Kw�������g�Z�j�v����z0�Q��i֝um�������#�6���BC��**+BBJ�p���Ěn��Xf����ta���8�ý�r�a��یB�q4���d4�490o��N��?����Y�x��G"5*W�J�-��M��9~��a�&�Kj4duaAi����0�i�P��v���%�`�G�;b��Y���`���h4ݥ㑁����$��i�F����0�:��|��yo�8��ַ���:tGFp���(�)�&>$����"���$:h�E?|Q_�$�b�z�N�'k�<mTV�����������0C':}�U��ă�(���D�� �ҕ[b�B�ē���9�=Ј��3N����t�,��C2d㗂B:v2iɆb�{Ca��ǃ����#��	9[!�N��#�ֆ�	�l`�E����l4�P�Ӹ�C�4<n���<�`�(��&<��q�ŭo-o8���z�t�,C��SG��F��'#9�
1��#e���i��!T|��#�V�T�Dve�*8ޚ��\`0�,ѡ:ؔ� �fn)�I���I�'RGD�HA�]c���MHZ[�k����	2r�"(�hN\���\��Sǖ4����%�u��"$��q�?��A��a��9`Q�g]�����>hx󡑰�u�޻�I4<M��_��]բ��X��5�����~��A�0~:�n߱���W.7�Vb�:�C<�Q+Ao~<q�������y�*�pp4=t�xI:�ԭJ�b�8���j�T�6��mB?B�M�J1��U&�:�DI�5� �N!{�~��3s�8@�р��:��eˀ��y����ڲ�8�ξi�Z�q�Ŭ��ǎ�8p�٪f�v=⊊�П���[<}�*��9���C����t�t��n�'����;�hԢ�IWd���&���rM!�,!�4:��a�}J���#����TÅ��A�l1<#��J�D �5e��E�Z��]���c�B�s$cZY�U��'kOU�yl+.���Nl���fZ��y�J�M�k����c�$�+K���%UH�F��jk�V��G�m�_?4���g㇏:x�Ӈ����2ڲ��eV@fI�
	 'r�QQZ���x�e||C�ʅ`}\#N���Z`�f	&�� (-s305�|6���$!s�-u��ð�Ƹ2���np5�	�Ə��*�$ KU�c1IcX�Hw3��Em�PÏ�����|��M��$���c$�Ð�ϝUB�����w�q�	Ag��BB�ϝ4p٦6�(��A�t���'�*�����*�"��<�B��B���ƃD	=�NЁ�D4Q��_6��-�ߜZ����8�0l�!_@$sh���	�J�3g�����κ���LÌ���x��7g� ���	"(�&!�12F�G��c�[�������gx�4[�A�I<�������^�I&�><�C��zU�����@�f�dv�
6?:o�Q*W��z����� ��:,2g�*���l���؏��f��t8`��5UD��FG�C�f�ބ�����C����K!Ҍ�,����6������#�6�0ì��!��e(Rdvr�t�i�47�n�����F5nB<�YБ���D\I�&��T*!�J�.n�r�ňX�m��k���Z\YZ���{mEyZ���*P�YkbʩJD�%�S,I�R�
6�pQ��~�b���#���Yt��SpdH�"pD�bEQ�i�B��K%UI��`���Jrl�����f���ka��"~�(�������౰�u�����B�m�i�\�ǵ$'�=l Y���	*��P�U���B���J�������B��V��6#l]V��c*5��r�� �vu����0b��b9hL���<�.Q�ݶ��*����cm~3��S%_>�}Ye&HЁ�d,����<VW����*��C�p����?-��Z�Z�q��`���,������ Չ�5�,�Vh�=�Ȩ��	t�m�2�U���&�8M�R�}���0����W0�>>h�1�qX�Ԯ�G�rh��� 0����\@�'�:d��tu�0�z<y�d(ن�D7��_�&L�sWy���=Tp��5�ϞcY�V�0M)�+��k�6�F I���á�y�G�u���7�ڣ2H�$���:�*���z�8r?p�꺖}�H���9�&���qS���Y�]�E�am��m<��?8�ַ���q�q��q�4��xo�g�'j�K��vo";���:����J)�lx���=��md8#u'k��OV�7P�+��j<u'1q\}L��W_K�%��N0_��q��b�!S���h�Z|��!��(��eTZ�u7�"F�3D$ĹP���Bq����8�[I��I��@�X�9z(a�<2͉��饰�q�Æ�F1Ș$���Y���<ds>�r��LW1��b��q[���q�δ�����Z�Z�q��o˟g	'X�%k�&5&"����F��f"�7)��SUW��h���	෌l~�J�!E���R�9}��|>�̅����prٸX���8~�#��H_́I	@�)��*\."2�K�����P���N���AO4��3옢�U2�IG���[���۽<~041���*��)�L\C��`�|����,$�ѦL�$�Ft�`i>�Z����t§`|��z�c����p�!l�؛?A��~Y�l����@�$�D艂pDL�N(A�A(��X��J8"tO	�xL<'��`�0J�	��D�A�'��"Ab%���H%�pD�6%�f�ؔA�"%���<"a���D��gDL�:'᳇�-�+el-���,���Q��$(D�'�'��N:tD�[����ֶ���y�^m�u}'ᲄAA�6B��<��RR�"!.�Dk~��AX�	F������BJ,5�SDAR��?i��O�u�PpH!�Q�)F2b)J2qaJ���8n�C;�\�@��
����.<��2�8YTaQm("2ӌb4e4e�1���Dqd;a���3I�&K��܈�y�|8�t;x�Ĩ�-F�
%{��L��C�l�CQ�h���9xƓ#1�%5�7A�m q�C��<4�+x<EEbx�48��y�N=�*V�";���h�BT���E�!�c.!�4tl���G�
B�'�nz�f���b���uX��\�9��Rr�t�$<D$�
}υ{��C��R�碈ݑQ#��M`�6���/>]!�"�I����+$�`N-ro��'ѐ�;͍�m��}�NDU�h�]�z���T7t�l��xt],�-ߡ�B(赇&2h�l�'�9�ydZ�`�e�ri0��u��O�ml�����3���Ɔi�M�i=��Ta���Ư��7�3����g+�����ػ�w���I�(���q�8��|��j��9�\�AF����x�č�=N�
D��W*�ESI�-�rB	�ҋ>�*֢��koS늒��ө֍#�ys5���-�Zۭژ��q�M$��������I#��Z�;�������R(�ۨ�v)�pj��☜�RE�(E-�X�U��,ڵ^rM8qBy8�r*�)%,-]��^�UF�x�TwwV�6֜�H���ϻ��K������eLz�D�CU|��֧X�ɶr�5QF�c$MǤ#�뻻��s\��_������O�V�^*���������mU�W��n����333���UmU�ۻ�������}��W��������FC
0�/�i�V��qk[�[�8�8�m�����F �(�!r2�"B���FAY[XQ�*�;fRے�\�`��"�,*B�tehlPB��UHB!0����V�D!VX$��P���m��]��*�m:��+�-L�
�2���T�Pđ[m
B��'R�Jڣ�*����**+BehM���i���ED(��D�KĭjU(Q����xp�=�e��f�d�~llwa`��T��O���f\�Bw�N���$���a4�Q�Ϗ�N�{9.��Vx�=8tP��@��t�m�=���'c����Q��,zs�Bzs��7P���*�X���H��t9��q<t?#�MF�4|a�a�*!F$�1��TBJ�ƞ���t0�ꡧ����!_]�r�ܧ	%�aan2����y���-o-g��ќ�ݫ�Tݶ�E�n7�,�y���� J�B�����a�ha����HA��C�v9��>_c~���3!1����̘�x�ç���E;x��e�"fT
�����|��B�6�J�ѶR��m[:eߘ[Y�3��X�K(U
" �,m��m��1�K��$+�]�~+ݫ3B{�aN�!xrH?�Ø�Y�1	f����U��H���4��Dd6c�zI�a���$
+f+�ɩO��:��|�N���-խ���qa�k1��<і5�*RD�B�Y��QQQZ+�,.����V	�����Əs��^�_>��d���&XW]�����������鷡�#�癉8�Wǁ����P䘠�+k(�Zlh�Rn*K)RJ��V��En�B;����{!��@�����������A隕	P�$O:�@��t���Wa����$�N&\�u�l�۲�4-�������Y+n�u<i5�x��u�Xa�[��崷�~qn�o-o6�8&�K�P��ga��G\EEEhL7Xv��U�;�-�el���|;h(��t��BI�zM5
	D��%�bF�m\#Qai.%�#!*Q�x���F�:���頁�ĄH���r���{����6������a��:s�vq5��33�4���}ʾ����6�~W�x_�"%$�ծ.��J�
�Cg����882�&�>��IC!�^����dQ�txe?��^�ZGXq�\m��8���Z�Z�m��oȌ2�� "��1����p�+�,� �Q	�F2�֒݊SX�-���^,F�t��pѪE�viDqd�8h��I!�]P�Gi4�$�HR���#�Hk�L�f&�V��5�;����14:��僙IX�Q�:J�N��b'^�#���[6ok�F6��З��h^e��%�컲B�j727��\n!"��E���a����$��;#!�p�B�	�o!�G�Ywa��<:]�Q�:�`kc�ٳĒPg��	$$�,2a�l6x��̍��<�A���aF�|z���:cn��h��>e��̏	�ԕtK�x�m���&x9�93���#�y�cC"��Y���.wo�P�8��ϰd����k��T���U�a`hw,�:'*��/�(��0xˍ����mn�o-o6����;�Ij�-p��e@j�أ�񍢢�'O��U*��ޫG���h��$�v5�������i���T}��p=�BQ^�vZ�8m�pH<agJ���U��4�C#�!;|#�T��|���RYi!���1�7	Md�<`l:\pnO�F�GA�������#C���˱2Ib�Ň��x�4\K�М�YII	'��X6>�lc>VKW�U��z�p�Ѧq�[i�kq�������ێ!�6Y��x�N钯-��g��������]�����B�`�(X�2�(4X�t�l%�(�QM�a=зN�&G�҃�፦�C���6d�ׅ����q�4Қ!e-��5�����{�kI��U]Vj7$d	$���4�8��
e��O��9	4��!Dblf��j�õ��_O��l�|I�"2E���\�[�|�(�ٱݗ!	>%U�x��q�R�����>ua�m����[��o-o8������~斶62���D�%E6=���EEhF�J��p�u�sCWV�{�bU�~�a]�9TW�i�<�����V1"��<r	�L�&��ի�Ϡz�]<���+�%S?A�(���e]�߃/B���b���r���ҨBIѮ������.�h��Ed-�0x�9�
��ʻ�Re��4:7�HHF�/�&���?���|A�B~-t�W�x_sA|2J�K����i�$$���l�6��e��qո��]Z�Z�q�Dtgi�x��bG*Pe)�)�f�!K�EQ�*,���,�FZ'�K(�ALAiY�i�2'��(�����!���T�	�r	ZV+�&Q�Vd����x�]�SH�;J�rA*�i�Q�Q�Dܳ*MEN�db����W��y��˙_Ȩ��	�B���V�El-D2e�V+A)e`�X�R\�fA%�B�,�<?s���H��~X䁪�L+�����0��e՗}q��$�P>�>��&��t<s�!�ō?��ؑ!v\�lz���3��a�A�����ۭ��r���Cf����_C�A��p�"|a�A��@���W+�}^�!���|0H1��nG�B���	!�Ӳ���I	�#LI�������QR�<���|z�I�Ğzl�X|�/2��yŭ�����u�:3�^���F�c�\��X��E!u��V��F����X�{�**+B5R���W��h�kA��R�d|��
��!��dק�6[�%J�.�sA�����c��� ���	�!��N�^H�<���fȲ]u79R�u�*V�X%-W��Y?�
 x�T��i
ZTԻ��L� Dd*x�'�n�?QNW�~I0r�T�8�W7��놩��}'7�&��;�*�۫�TL��ʲ��i_y[������[.?%�Q�"A,DDL�"A�pDODOtN�8l�A,AD��dM���X��`�a�`�&	�	��"a�<p��X��O�6 ��	��"xD�f	�8%�bY��D���""9"x��P��&	��&2tN	��w&�(J<��]ZE�Yo#�2`����lN%�8t���B���[�n-o-�y��|��Xx��Ǐ<yk��9�8�&�O�i����m�����w��]����W�|����{�x}��W=ק7��=�#�ߨ��t�F�G�ڷu��Οn�i})���t��w���^o��[�}����fNC����{Y|���}�<�&�[ǃ�����e볯�M��w�^�w�9�p_[n����e]��X���E������r���[y<���swuTd��9̛�ļ.�}�]���I�*�!���hӺ璕P�{=[��v���I�%�w��Y�J{fydY��[��i�:Ό�����������Na��r�ۭ����/~��mWm���fffg���W�������L����}�*�mU�����������U^*ګww}!�a��0��Z�qkyky�\Gm���`����?]o�[��O�ʂ��4C4Ң�S�|3���I2_j��!��x��f�0s�''djVQ�s��),�Leldpn |p:tS��}�O��`�n%Ԡ�^$�e��oi�OS!Yrg��$�W���I'����<�7=�oXP^̒I$�I$t?�Ѧ�L���������?���~[�-o-o8�����{�����Z�cX�2�3�=�"���Xaɭ6��	#�\�\&�3,v�a�����*�J���ؔwuf�2�VE�O�Ñx�k�!,�Sn��X�lB"���B�T�D��ع�sCg��cL��I����=��U�^�\����p��gҪ�D<�I������fL;�^i���7$I����,(��)���o�,h8����x��{�b�4:gfF�z8��G�vN��-�����\Z�Z�p���s ɟXQ�R(��)�(h�$��@�R�c��ǹ4�w��hiT����l��)IG�I��c�
1A��E��i1��X�Tܓ���h�.63��6Rn��7����dCN	��K���ڕq���e%DH�q:�-��d*�L�cc��淄�J.]�������F��E[�)"lD��-�G�$Yab��7�gN����)����4��Q�{}�a��	<8`z:����頁��$!*T�
�0ll��a3#�}�!�TU�:�:�s�[G��t�D~vm]W�D��NT�?h���ՃJ�h�p�Ú�wo0�B��B�P,�rY
�c�&B�X�J��풪���*��*Aҹ�r�WY땳�fK]Iȵ�0�8�1�>e�V�����[�yky�]Gܖ�]c���9�=���z�t�󗼼9�O��Ƣ��Xt02��h6v�X~��TB2lr'xG�G�tטC�ń!GͶ���73�˗a�:p�:I�-	a���	D(��z�Fۄ�\�r�>r?$��ٲYd(����J[r�TX�<
Q$~�rA�S��ۀ���|"@�D����>��4~��:�0�7�DA��VH����I��#,nN��/�:�����[�[�:���6�n�.�%���QQZ0��yFڔ�t�J�^NJ��r��!F<�2lڸp�x�J��H|��é��0��^��azx�"?>��RA˒*�r�����Ę�,%�X��<�������9S���&%�M9\������?���|t6��C0���]��v;�L��w^(�(�����b2�e�w���-�Yc�[.2������[�[�:�䳤҉*�4������x��>�\8})7�Օ���U�ߏ��(ᢄ�c�M��)!F��Ur�T84��J�64�6��4�?��`�7V��Y���u����鰘��j�������>z99pe��N$j�K\�$�)]�v�H��jǌ���nV�i'��zWkj��#U�귒�G�e�^[�qkum���t���iQ�h+��"�DtD-4L)!HR.\� �8��6�B#g�ej�F�k*fA�A2�)k%˔I"$�ؠ�7MX86nW��LB(��|k�&ԍq	�Ubv��b���G[i6�bNV��9
8ڥ(�5nȾ�clm��4)�9p}A*b�<F�e����3lZ�5#�XA������H0��]�����^o���fe1�SYcM��^�m�cN��q~�$AŻz<�5�|�=��vr��Qɱ�^ �֏[�>$�v09l�!�߲�0�pס܈"-s��Ǆ��45B�+�1��D�+G
�d&��}�� ��V��F�U�M��UXLLC譙e1�:ˬ��^q�n�����㮣�nL�kV�F���p󈨨�SUZ:rR�����t��$�C�6P���Z��G�ǅ&�5��+^��eDٱK,U���eUX�r��]��2���p��hp��(�!i��4�|��+[J��l;Xx�lO��e��H�nu�"� DH,���L�x��H�	���x�����jiz�	���R�)����M��˵�8�n�������2�μ���[kyky�^��#�Y��l��Ɠl��
�%�^�+�����QQZ6+
��x���c���k�F�8<�>+�C�HX|I>�唬�W��#��}���`�)�UYe���E�T5�IUR��1"!KJ:P��b��}��t���h|���%I	Q*��oU+gY8�O�޾�⊦�H4�B������,F)ۮ�SX�>	gߊ�䯩�bC�"�e&븋�j>=E���|����/4���-n�n<��㧏��,Pҟ�r���+��"A��!�*���X��$�i(S�h�o��**+D0�W
�h-��a��s>�C����Aw�<���@N����$�j9*��$nUk�K�b�������$�5IP�S_%C�z�I�
��8C��/G��ǡ��=Ol8�=8�Y�0b�.���膃�^;v�}����5����u���C��5�q썔UH��J�Ҵ�W4�`�����_>i��>��0N� �D��""t���6AAA�F͈�&�N�:'��0�a��;��`��0�8P��"X��BxD�'�b"tD���g�bpKĳeH"P�$DDL:P�$�D:"&	�8%�'6lJ��2|O�Ye�Yl""�Fy��<�B'�Ǐ:tD�:P�$�y�yխk[���o�ae� �'�X&��Q
͓Ez��E����܎!0�(���3M� ��\:?�jШx8�D2��#!8�sG�"���H+K����Dg�������f��G��BC�Ith���(�(v�P||�qs)w���5A�
�AAX����ԟ�$�i��]����7���ϛ��	9:(,e	9�Vƴ�q�2�>�}��:�ˎ�C�ܚl�]��ɝ��8��87Y�m:W�HX^6q�7QH1��P�b=Fq�`��� �oirS\s� �٤�p�����׹��A�RlTQ
$YQri�NsV�m_"�D}!��26X"��c�2�H��q�й���lD�|��p��:���̬��7(�!}D���8�F�^7/�2��l�f��"6(�اe&��-�+�օMi"�*Ə3Q��i��S��3�<ʹ����Q�B/!%�+ ���g!��z3�%�YI�Q!	�o�' �ʲ��d4A4�!�������R��c�t��Ng=��E�ؓ�k���V�%z�w��S���i�,����?��,ļ��KϢ��}SG�u����L�V�sx-b5)�#�G��&�k,Q�$sv����ݮ$)b��GuY�ى��kI�V5����5�7rŖ?J���O��lm��v˕֣m�I�K�WV���ԥ�MQ�
�+H�U=JCv��H�-����+�T���T��D�uƿK��Lzϐ�i=A�-țvi(��{4Vƈ�w�d�$��[<�m�Ɛ�8�� �vV��,rI��6��`�H��6ԁ�������W5Uw{�{u�^����}������*��v������333>Ϣ��Wj��ݿ����g�U^��V��ߵ�����}U�Un���A���l�κ��Z�Z�yky�]G[e�s
�TD1��M�*<�c����*��F��FcKF[D$�\ �2$�U�Db��$L+˒�$��(�B��Llc�H֊BX�VK���GP7!P��f��q�ԤUG�<krE�*��!4��1D��.�%�=�����hulؘK�le������vJBZ�%�,K!b*$�"pj��V�����_6��� C�Ҕ;:��|�`>a�wF�	���e��i����GN��	W|�[�d���d��Hu�N�F:f��A�6�%����>��|�l�����\�pӆ����D--���Q��5����b���<�2��p�>�@�0�2?J�J�O�#��~e柟�[��ukq��um�+��LM{]e��wrIs�!�3w�+�M		a?������|����	�T�ATT�����x����Ԓ@�#����u�!���P��J�bE{���]�s���1�J���[�B��VW!"�H`>��'���+e5e���Lک%%�:@���0�_x��:D����/���O΄��0PSӧ��G�C(X�x�L`g�٢E�����agK8b�[�-n�m���㮣����{�u5�m��.RJj�n��			9c9�2zL�*Jm�S���1#��C����]*�QR�U�x@�8Z1&�1��ep�������n�!�\T�XbArN�xuM��qLKיU�wV��*<*�.��(��x�Ւ�euw%IX~����rp9�᠎$&���$&�1��L�v5s���6�-$�eJ�~$8�
�I/,3��[T.�S���u&���t��|�.����[�-n�m���㧏����{s��\�s��4L�/�			�1�AR��g��~x~ч8�a��ͅ�G����̅<���,�e���d��M����`���� ��f����/�v���:-��v���N�,*B����;��8_��L�dx<	ݑ�ӧ�ITVƹ�A��5*�C|D]��>!'+�տ�X�	.�E�]]�,�v�C���<ѧ��Ã�c��x$|PI��t�~i��m�^y��V��Z�q��<p�K�[9DA�� �d�v
F3`�@lc���B�Bő��Y��M��-b�Qs!R�td͌��QX��n����S�eTD#l�n4�Єw-!T���i=q�uX6�&F��H�^�+M�V��j�P��n(뉩[S[���Ǳ���U����$$%�4ѱ�-�P�҃$Sn���+�7TnTA܅x�G1Yct)l4<~��9�&�o�'�X��g9�~1VY��BHeXS*a�����&��<;CK�I��XY�5%l�F��
v�ߡ�����$*���tf��`h�8>��:l�L5�	���Nb ��y��5�B5�dؔ[��b�46A�ʠ���m*�$�R���6W+gՕ��,,>+U�j��0�D�c	6�P���m��qo<������[�:�:��~��{�(ƞ�Hw��А��S_%H��9�VK5N����u$D�US�p�/�n���WV�FN�C[Z�]�����%bU�|?x2�GQL�vΞyÑ�4~1��_�CCK�G$&46(@����I�D��J�Bd�x#�oH	~�x7.f�t��
��I�f�r�Zu>&(�i�Y_*�ȷ.d��FV�����������J�z�t�#m2���qo�8��V��Z�q�Q��{��=�|_�l�f;D^~�ùJ$$g��4�)rbGN��c�Ãi����A���Ѱ�d��*T��:�!!%r��A~���g:�1��u��E
1�q�R�&-���]��G���WЁ'�վɣ�C�̙zp��'�a��
W������P�h�T,����	
Ҷ}�D�S�&�J�|����pх'��%J�c��3���p�gu��-���V��-o8��h3�Ε��J����j!�S�BD���L���N�><Y���$�-k񹠳��?����r�A�4,CW[�Qԕ�i!��Be$�LA��� ?�A�pmɤL8�1�h�ۣ�\�#<�~}����v�aC<��:�5�/�y���$d���>3���e5%@ټ�>$�F�����a��Vp�f�^�J�֑���/�-���Z�Z�<��㮣���#a�
qb�4c��e1�R�+�mKI\��ƕ�Q�l%bK,���ʙ������!����5�E��L�&;�ǈ��MQ�HH��W.V�*� �lKm�����;�q5���V�hj�;F����i�b�JeF�29 � �E����U��"X�L����%���f���!�a��E$-���a�+[�x��QN�r��D� |�O�,����WU�۟<�m��a5Q���*y	��ka������x`�8d�D�.Yl0@�ڿ�����t�h��>3��ޝ=^��T�i&Y���"�1�R��9���.�j�]W�)��x����~+pR���1,������/:'$h·��c!�]i�_�ykuk|��󎺎��0r�`��a�f�&�K-nܲ��O��"#^�9X�K&P��	9�W��_�����|4�:�m�Q����Hh%����|�c��C.���!��Cc�d�נ\\���TB��	"�񈂄��/�:]Y�����A��&Dլ@�/5�ѕsJ�t�����F+�s�ʀv&.�=�c��I�c�΂í���Ew񺕜�Zi`��i��å���� ����B�B"pD��`��x����� �"CK!�l�blD���<y�Æ	�`�&	�C��Ǆ�D��DD�8x��Q�6"'D�<lNpKͲl����8""'�� �Dy"#�(L ��tK0�,��a�^a�$x���G�[���2eh��G�y�q�y�^l�D�8"xD�����h��ae�Yg�W�E������{�M�ky�#��K��V�y;���?/���+��;'��T����N��gk��U�\�4�r��s5���4����y��p�k�uMw�}s���*�[������C˟?�o�u���Λ��;���c����k�r��P���G��Uf)5�z�{�'�Sy����ߧ��~:]�������8zow�G�u\97A��{޼k���{��Ë�G��Z��_H�vNk>$���z�F�߰�م��Og�w^�/���W�&s��SP��ߘ��ky�4�wuB����z��N���Nמ�J�c��y�=�o���kՋ�ӕ�"V�s����V�M�|Z��3�W��}����ޭ�/���7�^ۿs{�\�Y���g\ٜ%^X�vߧzɭ{���B���<||;���������iNΜ�'���R��T�nl�Gs}Þ����us�I+-��n�w�u���O�������yݓx�M.\�>����/�+�_rK�Ty*�J��o�w�g=ε쐅|�c�>Ϣ����[��~3333>Ϣ����[��~3333>Ϣ����[��~3333>�U|������0�l�fuն��խ����u�u�]�HHH4��h�UU�r=�k���p6*Q	��A�7v\�(���a�:3���L�t�tB<S?�c�
,.m�jy���IQ��weY_�<V��f�������þ*��i-���y%OՆZ����T�;�.��k%�'�����2:��Bx}�e��&j�����W��摧q�Zu�m�-n�o-��㮣�2�#d<-��begY$���*�i���|I�[�<'��Qa�.C.R��G�������(��-ƥ@�EdTE��qKs�8g�O�fd���c��:�FJ����'C.`�}��{G���$!/�߈�F�%��[( p����s8ʱB�����ۊI	�
��+��l� OL�T���=��G��<`�|2�y͗���_N�գ�y\���$���H�L���<��Z�����[�:�:��G᣹D*2�(B�Cl�0��� �d�������[����A9�ސYX"��:X"e8!�1t��è����C�(�HbW"�(X�B.&"��(82呖���[\�"�6I�H� ������I�h�8�BAS�$�H7D$���Z�������9��"�T�+�5X�ǯ��W��t>;(���n6�o��:Φ�9K�	�;^;��IL$�iC�A�^��2�Ucc%J2 l��x����x�I�3��)����I8�������x�m��n��݇�V�FT������w�lr	u,����J�	��#��EN1�C���S/�������Um��?&E�B��L?F�!�:S��6�������󎺎����?;�hBzL� ��̋�\��$�:�,���<<���O*�F�ݖ%`�x�"}�-�@��	�!���$l,:cL��&�Cgq�2�a���ɫ�f�>�VÇ��>�ڂ.��DR�b5v`Ŗċ�j�2�HIG�	������&��B���"B2ĭ���5��<WF��GP�� l9�%C�/d,�0�-�̭��[kZ�Z�����<#�I��8�rT��PŲ�Ό	#��
!�w'S�ޞ:�u�S������ȩ�z��Dd�+�-X����'����1d��L���iH!ZB��s2E�b�Z�;]++�ڦO0�V>-�o)3�d��:�+���^�9H&����\-�l2�+��5�c<.�l^�܇�z��w��a���UV�'�!�8[̺ӎ���n�o-��㮣��Umר���3�̐׫��,svI$�C��aM�����406?44�P�����c�����k!$6��.�=#���x<z�*U�:i��ka��� i�а��3�h��
v呷E�pt�M��h(a��^ݔ�T+}�Ǉ�K�4QDa*Bx��-�g�jH�	C���Y�̖|`��ͭ庵���ܝqm�O7�	EV"�2�!�!���4>n��rE�:,s*%L��GX�!��*53tՋ��)Ym&i��
(�&�W��!)h�ȦQ�q� ��e�86R\���sRq�ѷd���i$$�I��*��Z�*9)j#pR�ڮ��**Q+���I$t���X�B\Py�P�Bt�B&B¶2��u;!]�Tc��2bB$��O��O���t?����z%@87$c�秃�m���C�F�g���+.53A8�{����Cě+��F2OÙI$�hq�^$�'�����Y@d�3OC�·I��[nǅlە�Yӊ��v��N=+,�Q������
�F���bu)�b�����dM�?-3LA��2p����I<��%V��t���Vˍ?������<���][�#��ֵ����+[xH��=�i�{�wT�Hp~�6�����1������U�Yun���Ö�}�C��ԣ���9���d�����!$z�lz�],�Bc��0u�Ѳ'��	%�7��q����8|n�$q���2��b`�I�+0�w(<��<�=%c�g�d��%1�>z(���D*���ьQ��t�>,�-���mo8����un��6ˆ~�`���� ?C��$�����:
���ğ!��O	!��p9~5���0��:�����6��X4|I����p�6!гj�N+	$Ǆ���6���K��=���2IF��ka��G�D%V�e]��*�b͓A�F\��JNQ���Y[��v�հ�I����t�H1��O%UZ�W��_�a�[����Z�mo=�<��ëu�q�i�Lɍ���wc�Y-�1	RS$��VoRI$9f(d
�\�����r̈́*5`�"p9WW������XA*7�"�YD�\e�(B����ʚ26E�t�d��ؙ����0�'5I!�4��%�<�rۣ�ѲJ�:��!��p���#'ɞ9�C��A�24Y��5�� lp;5����J�c!�gG���0�9��_��~�a!���4�ն���˾����S��\b������0%�4ѺP LEP$QUl����!�J`�e���!HA�U�-nR�$��&YI&L�*�e�eiJe���ٖR�))T�)L���L�,R�̦R��IKd�R��)�RRf�)%2����$�e)��$�2��-JS-)j,�e6U2̦S-L�^��fS*�f�2�Z�2�R�*�RJI,��ɲ�>�V��d�YI2�e$�d�I�̔��%)&Il��Ie2Re��RRd�$�-�YI)d�J�K&JYdɒ�̔�,�K)�ɖ�\�䲚J�-JSK2Ʈ��,�J��d�2dԙ)*[2Y,��2Y,��lɩ4�%Idɓd��e�͹2RY,��%�-�5&JK%�&�ɖ�%��&�ɓRd�ْ���dɓdʦ��I�Rd�I�-�L�5&KId�dʺ��5&JK%�&�ɒ�e��d�dԙ2jK-��K%�ɓ%��e�&MI��d�dɩlɩ2ZK%�&�RR٤�dɓRd�dԶdԙ2�L�5%��&MI�%�&�ɩlɒ�d�d�d�Ylɩ6L�L��&MJ���u�,�K&K)��[2Id�Rd�d��d��Y4��%&[,��R�Il�l�$�4��̔�dҖM%�Ke�%$�L��U2d�$�d�RRɔ��YjY4�JL�M)e���4�J��i)4�L�Ri,�JM)�l�J���e)E2Re��)IH�JL�Rd��RiK-�K&��T�M)e�Ie2RJdʥ$�L���KfJIL�Jʸ�r�+-�����+5������R����e\��mee�Y�++Jʲ�k++J�iY�VU*����ҳjVkJͩYVVZ��T 0BuF��!	I��Uҵ�W+6�f���+5ee��������Yk*�Z��VZ�ʥe�������m+5�f�)�0
��!��"P1`�0�)HT
�B��f��µ�jVZ�f�Vj�e�+6�Yk+*���YU�rV��++ee�+6Ԭ�+-iY�efՕ�b n�,A��RHY�ee�+-YYj�ͬ� �*D.
R��$%�el�ڥe��ڕ�iY�+-iW%k��Ym��Ԭ����Yk+6��U+6��V��k56�R�T�J����T�ʕJ���YVVʛl�m*j�Ml��ʛYR�T�R�mMS�ܓ%)J�R��KjT�ʕl�meM��*�RՕ6���k,�e�l��,��5l���*��[,���m���,������YU,�K+Rʲ�T��jY[K5if�ͬ�ԳZ�m�eYel���f�Y�K-e���e�,�fԲ���e�l�ZYT��YZY��U�U,��ҩeYe��m,��-K-�����ʲ�j�kK-����if���Ym�j�Z�i[,��me����fԲ���YZY�-��e��jY�,�,������!p9m͖e�e���e�Ye�e�-�Y�jY�YfY��,�)m,��2͖e�e�e�f�i�T��)e,�,�,�,��YYfY�fY�jY�R�-��Ye�e�e�Ye�e���,�f��e�Ye,�5,�i�jY�YfY�jY�Ye���,�Գ,��,��K,��f��fYe�Ye�f�����-�Ye�Ye�f��fY�fV�,�5,�2�K6Ye�[K,�2�K2�)�ԦSJҔ��S)�L�SR�K+L��)MJe2���YL�)L�))��,�V��R�2���R�R��J�S)Je,�e,�)YJ��S*�R�2�R�e)[�\��i)�ҖR�,����VR��L�JJe2��%L�R�%K+JS)JiK+,�����YM�,�������ʖS)e2�S)����R����R�R���R��M��L�)��lS*R�JT�SWۙJTҖSJ�Se,�4��,��4��ʲ���eJRS*eiJ��L�JJ�ZiRʖSR�))�f���R�iR���S*R��S*R���e2�))�2���J�l�Rʷ]r�e�RB	PD!�������*Y[,��Ye2���ʖVYL�,�ee�,���JYYee��ʖVT��RRʥ��+e�ҥ��kt�ιZ�R��*YYJ���+,�)YJ���VR����)e,���)SKi���JU%2�Sx��R��RZRL�R�e��j��F�j����~a�Oë/�Jh)N������1u���V��-hK^J�پ%��~���Q�~���_Ȟ��ަ�?����t��>��q��_�L"����C���Ύσ�8��D�Du��oBP�P����O�l�����O�s^<(�4P�3�������kI�����������`0"���%?����?������������T��?� Z�u\�9[�o{[߷�����žM��ZZ�JD��W����A!���������?&�D���P 8�_������!?�(���� ����)���#�g���<�����?ʝ���,JJO�'�1
i�����p��|�dfa���XLG,�BB@?�S�����II��� ��b���`��XZ�("�T� 
)��ED? T.�Ȣ D������A������܊"�Q�`)���?��X_�E�����?!��� R� � ��� �5 �E�@#QX��1�
�(�DU@�@Tg����E���ů	�������H���D?�n����o h ������O'��'�E��������_�`�AP��F��m��h��h��T����������������_i�������d�O�O����� �|��������
���O���������P ?X��+�_�~�������:u���`@?�~ݩ@�c��B a��T@��?�)�i���S��2����X�?�����?��cc��,��+��AGNQ�Ё"G߀0��2,�K�E�K���6��C�֊�����R?�?�`�� P:����7�����R9O�%	�;�(O���"�)���N��~��a���\GJ�����d_�b��M���?�N-C��������������O�?�r��Ce�Ґ��'�]���0?�B~�������@�"-���������������P ?3�����H �k����m���ŋ�1bƢ�EEE��QQQch�bѭF�F64lh�1�1��ţcb�QF#1�X�F#c�F,Q�1��E��cDF"#DE�#DF#Db1E(�Db�Q��F4Q�1DF#F(�Q���#F1�#�"1�#F#F1DQ���Q�1Db���#F�F(�1�1Db���#F(�h��"4Dh�1�1Db��E���#F(�Q�1Db���1b1Db��F(�Z4F1F6#F4QDc(Ƣ"ъ"ъ4X�QDTE�#F4Xƈ�,b��(ъ#h�(،QF#F#��QF�(Ѣ��(�DTEDj"-ѣF��1EDTEDTb�1ETQ�F�4hƊ1�F�1�F�*(Ѣ�,hѢ�4bƊ(�4Q�Q�c�1�(��Q��(�****(�lcE���6(�cEEEc(�QEQE��Ŋ(�F*(�(��b�61�(Ŋ(؊4Q�QDXآ��EXѱ�QF�m(��EE��h�EE�6�TTTQQ��(��hأEF6"�1�F1(���c1ElcQ��cc�E��F�h�EF6(��(�cQF1�Q��4c�cF"�E�1F"4E���1E�1�1b"�E�1b1�#b(�b#b(�X��F"#"�DQ��F"�E�1b(�h�(�Q��F"�"�F(��F��Q��1b1�#��Db�E�1(�Q�ƈ�Q��b�Q�E��c���1cF�E��Q��1c#4Q�DlF#DcF#�1�F#�1#F�1�h�F�h�#���،cDh�����cDb���h�"�m6#cFƍ"�h�"1���Db4b+#F�����b6#Dh�(�X���#"1E"1�#(�E�#(����#DF"#DF����"4Db#DF"#DF"4Db��"4Dh�����#DF���#DF"4E��b#DF��"4Dh��#DF��F"�DF��"4DX��F"4Dh��"4Dh�(��"�E��1�E�4F�4F�#�F�TEE"*(�F�h�QQ4b4F�h�؍�؍�Dh��4F�#Q(�Dh�E���؍��Ѣ4h��4F�h���(Ѣ4h�#Q�lQ�E�4hѣF��4h�4hэ,F�4h�c4hээ4b4h���b1�4h�Q�DTF4b��c�h�4cF#��1��#(�E��#�b1�cDF�h�h���4F�QF�#F�Q�X�#1F1�ъ4b4cEhшƌF�1�c�FƊ(ш�#Ec(��cDF(�Q���#E�Q���X��1DF���#Db1Db���#b1Db��F(�Q�1Db���#F(�F(�1�1DQ���#F(�Q��#F(�Q�(�b���"�F4F(�Q�1E�b�Ɗ4QŊ(�DZ4Q�X�cEDTEDX��(�F*1F��b�Qb�ъ#E�F"��b1�c4X�4QDTEDTEF�h�F(ň����"�Qb1F�hѣF��cE�(ƍ(Ɗ4X�F�ƍ1�QE�Q�E�1�c�1E���F��EEz��_־V��_b�H� ~H� g��?P�8i?P�8���E>��Bu�����򁴑c��(����� �*H]ݑB�?���A��C	 ���?���?H`>2p%?�e3�06d-��ܙP 4?�?R����Ne��G�01�ԥ�p~v?�������=z��w��A*��͙��`���������������1�m� �T��?�������PZ~�0�����O�֦��?po�������~�?̒0�Ԡ��"��C����"�(H�s� 