BZh91AY&SYK���'߀`q���"� ����b!�    `                                      ,  x����     ��      �                      ��UJ
������$�)�@� Q�
�
�J���U(BR@�P�R�� �UT%@R�Xt  �(HR�P"I��| [*�qj�ް�P���%�Xtu�@�������jWTU9��ʀ�a��   �T�RI
o���hٸ��=*�(O��R*���¶��{����Хi��é_W�ҕ}�{��� 4��
*� �����:�@D7`��@  â�JR�z���JH� ��x -g� �`9��^�{ ϸ�O l<����vt}�� s�� �z� qp   h}�E@R���=>@v� ^��K� ����t{�/�r 9}� �9�@� �� z����������� 
 
X�JJ��^�$�����UD��*�� ��`{�����Ϙ�` y�ׇ�A� -����:t� yz{� {�J������i�q@   ��H $.��d �J��C��B� @\8J���y �`rv �@�  U �J����RDEH(��T �Q*� f���`r @N�S 	@�7`�� e�(�����x   [�H��`�� g� a�����  ��Q���wX�݇��{� ��T (9򂤕*�%"@H%	�UAB��x � `=݀9V@,�$� 6à���5F� :��p� ݁���P
Ϩ�@v ��� $9 n`: F@9�%�� ��� �r >�    PS�JT�0 d0� O�Ĕ�T ��@���ʩCS�S��d24 4�*Q�%Dd4��F&���&M"(eJ�d` # b0T�i"i��O)�F����D�'�������m�i|~ ��z���=�A�5��q��H�(�6�]~`�(�ʈ�*y�(����(��h	�O���S�����<Q�誂����J�|


����}�ٕхD�0��
�dFdA�U���e?C ��eQ2nʎYUL�"�e2Ƞ��(af,*a� � ��S,�XL�
�d2�dL�dL0&XC,��P�"e�2�n�e�2�dL�����e�2ά���
�:e�Cv�:a3�(t�0�L���e�2ȝ0&XC,!��*e�2ʙeL�X,��Y�l���2�0�0�i���W,�� � e�2a��2e�0��2��� e��(e��,.XC,)�e�2�ar�erû	� �(e��+�#�W,.X\�:�p��G,.X\��axar��2��VC,�Y\��d�Y]X\��dr�hɖ,�XC,��+� �2�Y,��2��a2��D� ��C�C,�U�"e2�(e�A�*��DC, �YE�,�YA���dP2Ƞe� �
!�,�0 e�@�*��AVC,
Y��eE2��e�CvA��a2� e�@ٔ@�!�,��Y@��2(`2£���x��Y�4��b(i��Ę�]����-7	�m��ݓfr����������ä��(��0A\�+�� ��1���WEZ�;�+ڻZ�s3LQye�I��]�]����$�Sw([3�or�Xjͳa���UWLY�,���٦3�N���xi�%Χ�n�{��g+�6�����Q����&�L�^�+��7nkvT$�Z�cY��(V�~���քL�s�λ�0�6���'�{�gҀ��Ý:oUS&��64�B+�Ի���Uʆ��������:�k�]��O�ڻ:$�F楬�N.s�בD���!e�M<U�F4e:�^��U��Ǡ��r�����~��N[��[a�.�g�F�)�TOw�u����� ����ɧ�s��M�,�=Bc�DYu��D-]3DLR�����~�ɅR^�7e��8�LOE�h/i\2�y4zݷ�Y9и])�)3�*G[���"rqoE��,o��e]
��D'�m�`t���ygcx��d��v)��-���"^���1p�����sgaBN{�b{b��Rce���OXK��z�0�3�`H����A�9
��Zg*��A(�;�-���=�Ϝ����b�ҏ�,sTM=�h��͓�ë;�-����]دovzqE۵��ɳbJ}z1�ܺ�iDAe���Nݧ��L��丳������V��ө��s7Y:�YgQ9c�����3�c�n��v�.�ӗ7ot��@N1ۓ:�V��H��'�Γ�I>K/>��'�h�E��5���(�;���O4�c��]WEȫh3�h�6cIe�>�k�f��Q�H��X^����Ơ	�l��Inw]˗ۣ@rU�-�>�b���������5Ͻ+�7b-;C@�i�����u�1)���ys�ֆ��cɵI�W�v����S/al��(r����r�C�M���t=�j�[ɵD��Z������]����ۡs�͡:�� ���j��!�A\8�p�$/X��
=�G�k��۩��f\ٛ�v�Gj@�6�rr�6>Mn��I��ŗ�����5�l.Ie�\:ӔE����Sf�;�»2��VνO��{$���}8���Z�	Ϗݽ�tZ��t�orikj��7��]�8��A��1��Ք(�3lxa�7�9�p҆t�hƔ3	}y���e��u��i���&��V�N<��1�9p:����Uқ�F	l�y��^���3����q��hW������:m�0M�t�+Ӌ�m�,��&l��xpd��t�����۴���	�j�:r�:�ʠ���{.�Ղo Jj=�MĒѻ�G6�(�\�-����,�if�7��RE�k}��F��;�!��I�R�i�"�STC
A\+�fP��Ӣ^�v������{<�^�sF��zE�1eq»�{��1psR"�7��H���w�S��dQ��A�oê����t��f��]�wAkHD�m2tquC`,�7�d���/���p��d�Hw 4���J�釺�{����#�;l�}��uL��	�龧�r�ci�����5�<8���Wgai�o<0�� �ou"�vr��S��6C����ٽ�6��f#�v�����mf}�Y���*�����Z\tv��9�=(�L']]�Gmy>�1��br2�wN�gU^Fկ���Am�i��h��9Cb\Ԯc��Iwuf�g�S2ٹ۝u�릝�4�3D�(7y��S&]а��kPӵ�ݺOlٝf*뱛P�W�md�sg�79�m! ��:2-ý:v��iޯu�'|P�N�g#sSJ1�c��<�z@`&�l��Q�a�l}����M�㇛G���v����J]���$o(��8Ӌ9+���m!�M�uke�Ν�4�]#Jo�,}:�������7��ǟMm�y��Η7i0 �H��Ck�k�+����3S��ɘ�`� ��bS�˚tI{D��Id[�(fDjY��4K�5nr��gCΖq'PanM�vcn��s{j-��&>'9��X�7�F����Hc�@���&�/
 *�b�o�6[�,8D;�ƞ'"��# �2(��d��CD,�A\0_���u"�]��S�J
Ǉ\<z�<�p����.��>|��VE�����l(�d�j�"�v{�Kf�{��-fN�>#�Ϯ["���݄dW]�tq��,t�>�[��L�;��oC(a�J��cb�/�H�Q�L�Wk���A��G�������_n���3���+�V�������=�݅��  2�rW����5�[P.���Z�jhj=,�C+N�����&���rSQwL������1�|���f V�֌&�v=���h�b���f��m��N1b�Q��1�@�b����caȺ�q��K�1�sq��8"nFo'Y�,9x�D���F1�K����]�U7;n�/����%�V�8OuYor\5=�Z�d���G7��lˆo<W@�D
�wg$������� ���-+���`��y��m��NN$����6�֮l' 9&�����=�v�W��}[��6���;�D�a-��z�a#��^�)u�{dɹ��n�6�ZM]ë�W�;�!ڕ�:*3������{wy ��_ud���n�-\y�0T����b��r�tA&���u]Ç~צ���N��wVnnՐ`� 廌`��˴IJZ|64�������"��u���3y�X\h��rM�;E*��35�n�E5(��=�p�{NkQ���^�^��龫uE�=Zyv4�9;��:`�[C��6�m�)/'t���9�5� %�5���(���v@����M�;~J���VUg{`�C7m�^��ͥ8���m��8_gK��.�F$��%����{D���{cK6���vwi���@l�:���-�r��X܍G�G�rq�w]�z��	�Ӛ��z3���5w`�gG
\���w1�Z��wOy.D�0�s�;�z ��\-�1��Y�6
SN�����V�Τ��b�EZ^.#5�زA�tre��7�pOm��u
>M��|�ۜpሖ�hݓ�5bpagCXf�ƺ�v���BJ�S.���w;ur(`���;�pB�D.�}�*閄'n����y,�^���d(f�3q�J$:�W�4������T��B����fҺ�;�l�SeLu���43{�\'�����ɫySɂ1W�Pܵü��t��c(%T["�Zd��Lt��hÏ/.�)f@�49t��՚�zM&}A*<d���!��5����
U�V<5i�ec���[�Ծ���+�z,��jxe�˷� !x��bU���� ݹ�(˭���ŔI�wwi�q��D����r������+c��ذ���y� /�a���{�`9�	A���K�A��N�D��B�hk�U�hie�n�rn.ǐGN���˝,룣�M��tx+.^�A��L��3�ծ�v;j���te�v�
xF��^���[!�Gۦ�W`n��S���س�H�_ƌvnD:k/[�Fގ���qr\8v^���d9�Ņ�t�x\^�ΑnF�>9��)�[X&#�f�0�;:�D��8�7$Q3�i�6R�Q��1:���(����D�H]��m��2�r7q�
5Eκ�E �u;�or�_!�>��
�Lߐ�
��'i�����L
u���_n3��kZ�aw���+˺5A�<�)��:Mg��m�ڍy+qA�s�]3Hj�"���@�zNl���ͣ��no��p���v���Lʉ2`׈�{�c�]z�K8(�:��l��N���+��-P+�dA���T�t����� n&���F)��;vG�Ov�u�gs�fM1�4�9���%qB�w/P8���5�X����+b�6��ý���uPn�BІ^�v&�,��6^�s0��[sl�ޘj����� [r��8[^r�-C='6�~���g�q�5N�\\s�E�)PW�t-Ș�V<�;��wU\�O)�Q<��P�@S���]����FZ��ʷJ݉(Ut�|!pP��^������@�ϰ.{�C�2l��^v�o��3~=�����v�C`�����Z1��kf���Ҽ�|FIϘ�Yx�Q�Ɛհ�h���9v���g8sF�j��9�vq���s�w%����2l
���+`Fs]��j}�«sk�2�+�Aٻe�N<-���3:29�K�����Yn�FR��c�m���Y�}�*1D�c{�]�B�
QrdK�N���܁D�����sy��6F���d�X+�$��s����å�؜Ӷd+�o'����5^�ե�sw�uv�����'yq�kM�%�%���B��ũ%��.M��ܶ=�b{'�����:l�3��Z�>فv]�7_,��
|Θd��35�{.��������EmiY�8d�3�8������w2�C;�]���c�=�\{(&Kf����p�ظ;NhĎ�e��u[oFZ�V���f�&�.h��"�F�ܽ��+�Eқ��˃jYTy��`�n�Њ�Ӯ5Z[9��s���ǧh���gL���K7w{N�vd�s{�ރ ���$��غi���ӓA��۳�K��Q�z��E���g]{D啶@1��w�`z�<i��wc2��Շ�=#L��3RT�Lj���3g5�./z�t����F��������K ��N��Ϋ`�V�����[Z��gE�0Ϋ�qۻ�ns!1Z:��Ӎ���M]ځ|9J��]h]���Õ�Ě\��9-`#/qA��%	� ��{�o7�X��9E�5H����w��w^��)�v��bp�d�,Z�A��� {t(���X��8�N��st|�_^�F:3T��B~B�tr۱9�m�i�U�N�l-�v,��6���9� l�r��3vz��nm$���/y�̑��n܇"<���{A��D��:vQ����.A�f-R���){�gs@ǈ�Ӯb�靫{s���V��a:r��\v�E�C3�AyS�rg}H;�oZê��K!d�;x�8V�n�&D�c��t.�Ns��9����;��H�-3���sX�@#�$�wX��%���F�6Q��I�WN�N�IH�:	��̻�V��k8'2Я*W�r7UP���-f��pd寮oYX����Jµ�q�b�C�� {���d�@�8E�#bs�T6ػH��tp	���w��v.����;Y�1�T)�'�Z�[�����5��L�%r���8��Q,\@GmN2��`�.r_<v������%�u���x�.s�E��0�r����EZ$p�4�sgV�GP�lP����Z�Fit���Fi1dqr������tɼo#����gop�{:'w�nMqn�����b��E��J�G.��v����橜�d2�Pn�S�}�US��I�uX-�H�Nr13�	I�Ʌ�կv�mu�Y�%�7�j���ځz��N�`���GWNvS�wc��mE�9�� 5����c��p�;��E\#.��.�����.����ܱ�v�~7�: ��|�^��:��bԒ��'�ʭ�[{V�n�Y��7��fϞ�v�{�{D�h�桎���	ڄN���e�<�::�q���Eƈyw"��:0�q�4oN|4�÷b��-�<e�*���t4y*��y�;�ѥ3w��ͤ�V�!A����ZWr�ˣZ���{݀w�sx�u�0�'rZ��Ntŏ)|�i�ւ�5��>��|���<έ�zճ���`��
<'e:�`p�s��,} L�zܛ4=��@�n�xR�^����Bl�Kr��� [�jjY�&��b��� 2���-�a���[6�&���(����:�_A��Κ�b�M��|wEJE��[[cGNfo>��'s�
Ǭ^���&PZ�4�	���그iĨ"��ֽRcuN�H':�tq���3�镔�U��fp�ǳ������M���O���w�g�k��ׁ́����c�d�p@�w�ZuGŎ	�E�o�w�$O\��]�F��{n���VWv ��М�ջqj��h��r4�x�a�G]:��s��Y;si�˺�<����ނvQ��Ur���,�ۛ�e=�Dz2�9v�F)��a�=�T¢ggt��/2VVOS��,'�&A���H��e9�|�뚰aUҜ"m���U0kc�ٸz��h�](9Ҵ�z80;�4(��r\I�;-{^�pɉ���3���������0r��s(������ɒۀ��z[�D�#��C�z���<�L�:l�ղ��e��jC�`q�6�۵���	�Ƃ�< '~�㷤Ca�H�^<6��joyh$m�ⶾ}�3\�Vx�Ǟ�x��ż
�o1v�]�7b��6�&�"¼2�#�����;�po���=�ȔC)�I���^�Q�|Γ0(w�{n	����7w&�=��ޅѩ��R�r#�e�H�O�J�{_��7�3��A(�wn�h�Ih(�⥾m��Vj���K�ǯ�lI'|w}3wg��]�v�4cx�k�y�q���l��}��մہ�S:J/^�e�m���0��Y&��<�����`��q��`ػ4\��d2�%i(~*�W����,����v��5s�N���O�,M�yc�I�|g�����ѝ'sMH��J���N*�W� ���C�N�~�°��h��7{���7�&������`?��9w��0��*�"	�
�!
@@�T)B�UZ@ZD)hPh�(AB�P�h)�� &$JZP� �T
P�@(H�b�(D�Z
�
T�
EĢУ�Q�T�(&!)TĠR�bPJJP�U�)@X��P� $�@(TJ��B��P
P�F��� �
D�T)�F�Ц%1�DB�\H$D(E1 b�R��R�A�D� 
E��U���Q���E���(��EĊ4 ��X�@�E�L�_O+:��"�$�R[�����>2��{�^��<�G��0�b[�f�˥��͸���^3��ե8��W�.�z��U
��R�9J�p�Zv9��z*�:��~T�����N�^��=N��+;�0Q۬rƱ�'q��{�@˼��)"N��@_������~}��/-�?���������=�w�C�[m|���h�㮼�s�P�M����ڎ�_OE�׽���nM/����a�Mh�۫-ͺ���N����U(ŏ�Eİ>�V��H�;,]^I�\^�9ޓ�,�w��HÆ��鍝���8��{��k|�
'��^���	}/�0�e����U��*���f�v;�>O�t��'S���fr�Fd~��|>\*~�ٽ�(ϲy�G��Vv��t9����샽�	�4��΂Itg��M1�ǌ����_�C��Ƕ��YR{t�
sڴ"�o/��z��z�<�3|��^n�ў�[7���Kw	Q�㖑t�E�o//)|����NX.�}O����z-6���a�Ƚ�#�uܵ�zA
@V�/�g�*+�o�TiJF<�=��'�2���{�o�����<�цor�����Y/f��{ڰn�=��/�	�{!w�o/}Ӯ8G��5��6kjo��.�?W����B��7�n���ߕC/�Z�[M��gnx�˽��<d&��.�gt�	Agp��m�ظ�맃�o��g=w�<�]Za��d'\�Z9^�6�	ڠ�d)kȇ;K����q����ra�xz��ɓNP�Y��ؼ�^�wr���K]�t�0��}{�4���|�E���P�ϐ�qo�0������}�f2/a9Řq�p^ ۓ7�ɱv������[{���{s�7�2i|��׺�+ۧ�pa�d]�t�����L��=�����s���E��|�v��^+&�۞K����i-�κ)�}��т[����r/l{��&��/���.]Z�ޒ�=���	ǻ���4���:�rI��)�.��.;v��|����B��p�{�G�OM�ǝ�ηO��w�V=�����i�N����d+8=YW,��N��b�8%s�zM�u:g��U�^�ܽ��v�����BAH���Jl���)۪Y\Ә��n�=������7s�Zo{�O����=攣���:��9�Q�����sv�_��[�)팦��w�����J���z'Nq�Q�r)��͞4�~�%G��'��=y�^)�U�x�!��{������m�Q��焋��ݖ=�������/=��(�vv0�N����;��F��1b�]w�i�}q�r�z�d>��4��x�Wa�=�~��bh2��tNY[�����و�{��b�����&Y��w���<a���~��A�d�X���ʗ�&�����o�=�֩�/����u���)������j���b�����3ݕ�P٧n�R���ó����;V�!���3����2Qd����_W����y��{�K�ԃu�匕�S�%<�������>�6�<uj�Ol]ݔ�q{!�g���"��w�����Mg��O��,��1kk��o�:�{����޴o�Wy�{b���;<ם�5�8>�ڗ.U�f����w������G{X�<�xz��I��~�JY r����Ǽӝc�����F}��G���^�VN���|oz��/޼�&1�庂�����8�9�C>�ơ�{I�FN�=!1f�j�|�f�-���)�`F�<w�s�w�3��h�^_>Ə�I�����út��wV�Yz�v�c�C�$���s�6�|4���a嚼V�a!�r��b�B/�jkK}�T�<W�;w{W����B�'\뾕�N�;��M�����X�O��_=��H�Tl�p�zj5%.�O��a���{<��0C7-��pR��:�'�{@|��ȁ?#;=�W�A��;�2�^�C�O@]wp�9�c������ő�=�o�=��e���5�`���lug�����i�8���p��օ����(�Oz>0^)�yӢ���s�:�M������l;�ۭ�f�_������{�.٣�C������� [�љY������g����w�Q����������3ۤǋI�}W�I+��l���ި+oYA�ı�K 8�%�k@����g���[�o%����Pna[>yv���7�G=�m����F7�z4�h�׻'w�ʡ��\3J��wa����㞜3�X��Z�اK\������|ډ�F��3�6Y|u[׈��鯏�i�܍&��|7�����p�Y��q4��fOi�j<�G�:Y�gjYI���v����H�-h?�C�a�)����h��eW�e����k�.�83�o����M����V�z�����u��d⇱��ܫ�}���yo@s	�;w*�5s� ��858���*�P�L��߆P�駳�gNg��_��݈���R�|�Eݷ�f��_w����~���ϟ��{����l��5o����
���9�����,n���8x��\�f���I�����;'S�A'��5�<����rZ}9�J'������8zo�G���\�����v�)�{�L���d=�>}ػ_{K�uס���V�����޻�N��۝�L�F3*0#������������K@�I�,�u����reܜ���7ް�V2>�ҿ8���N���~3�%��vn�#`I�kD�����=xn���e�f�kh��q@��#V�B��P�*	� 8a���;������<�3�|zx�;�7=@K���`�rm���q��7�����w�
r?4��=��G����o�����dʶ�;Q�<�<���cT2���c��Pw�5�p�����ި潄�ې�[���b���߽4"�Mo�U���q��{_pE�=����~�p��X�ۥu�o`B������ܫ7 �Ʒ�О=��7��nx�|�ae2l�sqc�t樽{f���=��LɷڄP�0ߑ�w��>�8	V,���v��h~�+w���n��h�������Yѳ�Jl~�\�!�8y�-+����vx	|X���ɲ�������\'��y�v���H�L�z�M�f���1z����ޝ�-�ū�=����Q�;��wBJ�!�g��;=�v����Kipۇ5��7J�V���~dp�F��zx�o��˕�8a�zd���ov�gc������qo_��N��sE\Loj5w_;�d�#�=�o<�t`>��J�*&;˸�L�OF��D{��F}����fJϰ���z�]�aqU�;�ƺZ� �^�i��3[�{ޔr#x�=�	3+��g�/�����5��[�.Z����C��{��$��Ȼ)аxE�iK��NL�o%�%��/�g�8E�w�j9��y�xw�����y�yW���c�6�|s��υ�18fG�OwO{G����I�c �X=�>���5�ZY�85��sq�~�����Y�����dh{j>3���`��o�{{ ��.��OxxK<x�}�{���v�z�ӵI��7wR=���j�jy}�S���N������g��e�9�.,�e�F>�8$޵�z�͜�9��j�\�y�piz����{�\>>�+�׬���]���G��KZ�{S���o�Ƨny�x��;���q�qν�<m"��n�ۧ���nȇ w��O���c�����ͅgz(����=��7�}�+�;�XP�~e�Y�ő�r�uz�����3�����ݦMg��N�����|z�/,]9�^`w΀:3O�
����h����!��f�ӽ�[-�
���U�g�`��wF�>�wD<;�<s\�n�:��F�&��޻������|;b���Fz�}�wk'�E�:�_oy�z�d��p����Ç��[>2�FＲS�bΙ4����Y�p�}&vՒe�W�<3�9�"�ݛ������{p�}���g=� Ś��|3M�*ش�K�0�f�y'�y��)y����
;G�׻N�w<�v��[[�tL�f������ԧ{q�������fo�zI0-ې��K׷�,zd^k���e;{w�w!�����xj��Jo%�7���`�{W{���n�����N0W����׵̄<��{d��/�D_e���z���n��j�����|N�H��JJkC��¾�j����0#c���h���/�WY�5�}ٺ�/�=�n����I�틏�o(����`W��:P���T���u�(1�պ���U�@��=�������ԯ�q���=����`�o<�lN;}�,�db
Ĥ�ï�	͔�s{�)�>�L?�����=}�ڋ��C���ã4�bKf������ᩥ��/Pыç�<J4sZן�>=y��U�n �y�V��[��|��=�]����ު��ޠ}�ݦ`��=�r�=�ދl4���?.�嚞����8�.y�{�i��AT���Q�yp���6����S��`�U��A�~xk�v-7���>���J��~�T;�z�����<�Jg��rt("�<��'���&�s��t��K�u��>����f�ç�b��Q�����y{P�����55ZW8j��TyN��VDAņ���<בFy#����ۍ`�on���L��������v����r����N�t���!�{5e݅-ږI��O��,GT�?U=���-��������w�b�d}�t�%ynRN���P�=t�gy�g�Y�o��_U�����t�4�j����V�M�D�y/��ˣ˾�p���ٳ�W�(��<<�OW:�k�w��m�U�hQU��C��<T�%{7#
3/���أ�\8�
;v'�4�)�MKMZ���{��sxY[.�p����.���
�ok��s�������>u�un���ʲ���`٣K
N�3�~��v��w�2��^�2<<}1E�Ǌ�v8�Md��̶ �2����C��{���|C��]����;�>��2@��*��@a-�O{yv(!���WU�w}w��9:�;�O=c����z���L[p.�"�]�G��Υ��=is/-,j��<Go�͜;�^�,��n�'�֯y���}�	�{���q�~��Oy�<�}���-��m�W�G�J�]e��HI�鏋�����fu���a���S5���{��e�7sL��f�����)K*��A��G>7Ӳ0Z+�ӆ�|�ѳ�ܷ�
�}s��9�2���+��H�o?{��_����w}�k^�%���d�/0��z��]�=��]'[��&����˝<lkft�����8�]���yn��Σ+٩;�>�)��V�(�����?X2�;ΰb��؏b@����HR����'2,�} >���*�(c�+�������t|.p��{�}�W�%��y���mI�a���9uQ!6�2.-����.g��J�g?cHy��a�:�7�K��6S�+�k��O���^QO�$���W�{S����^���t���yE�(�P@$�n�����I�]I*������[pY����}Bf��YH/��ݗ�_p�� ��Ek,�Vjs�x��O4��Q���>(N�<zr���s�<y1s�*�/�f	��K��y�I8V<�8y��� {v���>���Ӂ�7�P�o��'w�y���@	����ۯ}��Ĵ�H�ļĊjIE��p��g��k�,�M��I�ܻ�}^ x�G��� ��ۣbddy}��Rg@��Y�0�8���9N�o�I�<4�,��[�h��1��hǽx(�'�w��wOI����w�K�_��P�)�0�Ck.���U�߯���^�C��s�9ş	
�V��կ��yQy١��=/&'�����z#��`,Y��{�JwܷM�a�<��u����v�1�{+�v��H��o�����v��"�?]t9�M�=�{��|8�{��sǳ�|����v�_��*淗�Q�Gy������ Bg�51[=�BP�)��ȼ ]�hƮ{x�؆m��)�2�U�Qe觽���!� ��w4�o`=���]%���I}(���gc~����p'c�we�o��oex��w���\@_j<����r��������� ��|O�Lz.A�����Q�rݯ�>���0|YBi�ݞLW�W��.�=�L�|��o>��
�=��cuI��pJ��q��h/��F<��zƲ�����W���؋0���7���{�������C�=�LC�VlKˌ8b���"p2���6�t�)�}�Ov�K���~�n�3Q�Ȏ�zv��}��&���vmƞ��n�lo�M���=�M�'����Ev���m>xl���O�����G�!�=}$�8xR�� g��t��%Û]�bzC��u{�X�j;��&� ��9�G� "����N�!kBy'�N�=��Tɞ��%�!��������煭�<�Mv{�p�'�˶Tw�fi��sE:W븬�XL��(�Oq�Q�����o��To^����{zҧ��_��C��b�|�(�.if��>��^^>�p}7�/z���/�vP��C=�?U^���$���r�r��vxG���-�z��Cru����zeǩ�э��g����w=�܎��d��Zo��_[����S����}��k��Q�ϽT����osb��q=<�Ϫk�5�<"��eۛ�:���s,���S�z�l��K�yg-��������ӭ\U+;�n�3z����l�I��u4lݞ�/'f�0qɸ�9�^Y4ӽn�hI�/=�xv�!,VvY��s<=����2�xq���wo/{��V��y�r8w�a	<4��g|Fw_L޻����}��y����G@�1��C�g^3�����a�����L�7������}�Mݳ:��������{��/�|sK��s�V������̻�z��4$*,D���ڭ�@��	�vz,��U�76��o�ŁK4,ɇqc�oΘ�m-6�-�/W��>�Wփ���{}�߳��~(�������}����}�wggY�g�^Nߏ߾��*��n\1ѹ���BRk���u|�-幔U�E��-�חG���y����zO���]WY�2m9MY.��lM-ԏ	,h�#�U�{xݬ�"��n�mY��nb��J��WCs����-�3�u�y�V�.�ݻr37kX��B4�Ѳ����F��Ig\�|�#	L�١�-qr�\n�Nݵ&��4M��q�Qs�4F��e��EZ9m���3�{n�P��N���m��os�p9r�Y2�Fm�<���v啊���J�gA�Tk��K��vx�
��	ɻ���az��J�\rx����un���3�-� ��\듛`8�s7\nW���M�Gn����Ĳ�e��"�	�Yfs6�Ƭ��h8�h�m�`車�On��#Lq�5�c�NѲIw<[��τ�"�Cye��p�ۡאC�aU^q��KN�N,�3��O&�M�m49��mN���ol�� v�6��+��[�BW
v��Imm���9��<����v�p�f�ˋ��N��Rb�����i�{�
w#Wk[�g���b����V$6��s�,�-/U��i�����L�õ�u@m�Թ���kV5���6�S[��p���s h�nCО� trR��&���A� ;h�=tZ�`�4% V��o:6����u�#ɬV��]��nN�<]�+-�W<rѶa�HXj�L]e�k�;rR��p���U�a�a��[��ΰ�;@���9(y�e�t`(�7d�ҵ"0�]�.�{H�%�K����]b���nX�2�j���f��v�K�F��D=N����J���u�@,˦ͷ'F�.҂�kڽW��An�SM�䳍A�Gm�屦,4c.�0�eصv���'-���edk�3.al���Tks�����z�N㴵Yٺ�^��k���d8{�6��1�'f�C����L�<���-jʲVa���0�k���P#
:�F:�[��5 �E��m\k{r!�!�!�M\l���خ�v=n��J��م.�CU�ŕ1B�Y�)���U�f�r<u�s�7:�������y�.�n�{*=�q��x/,�4���i��v[ku��5�ہ�];]�c���,f��6R�,a3c5v�bᗈ�L�Kّ0Kb	�݌�[ɝ����Tm�\z��笅Fgi
S��lA�e�:sV"���(Z��э�uք�Y3�d��:�F�ؒyzֳ�c	ـ��\�T��+��s<�7馬��ɘ�"ͳ�����ac<'R��Wg��Q`�&q)]�0Ǐi�]Z��ؠ:z�:���k<���\V�N��Ba/f�3�e�3Z6�e6�A���K�8�1c�2�f�36M�`��[u3���1�JǊȤ�c`a�0pq4���
�Ŏ���2e�r4j8��@�7b�NI�G<�x��h��kk���D	iF�a����0b悱�8�H�8�j��6��+�:��n�6�n0m��v��=I��noOce] 0��V&sJ`k!l\����u��F]]�ZF��&$��7;k����+�oee��\��F��]�!u&��zra�o ��j2H�Kx6�u�ΰ77x�5��.���A�^�;t��K���Ss���g�烥�g0�^{D��/k������K�M��g��Ny]�����6h�\EKz�Ȼv[Un<�$m�Fbv�{]��x��"�R{V�C�O,\���3ϧumn���K�1)3-�K�n��O9�ø;=��nE�[��k����-m�Rݎ9V�3h݂[A�@"�(��蹮����2=ӳ���k,�hQ}��i8���q�\k�ӑ��[h�㫯GZֻE��蛎nM�%��n9���z��\s�u8�ölyȜ<�u���Gn�vy���0c��9Hќ.�<WY�l�`�x�힕�v�ex;oG]�5ts������%pm�t�9Li�2]e�7���.�|�km�3[L����6c�K8�1���H]
�l�M�m��I�Ŧ(8��O�n�&�Q�]x,=�xF験�
ҙ##ձ&� ۓlRD���1u�4l-���й��7\h�p7sk�5N������ޞ6�β[��2`8���u۝�Ք�K��Q.8��:��t=4c��&R1��N�rc�V�c[;�\Y�r�%�8{1�6��G;�l�O(�k	-4�t�� ;T��X���p��ՇGU���:zn��ܑ�F9*�uy�m�΍�F��؂
���O)K�N����\�p�\��ͻ�Q�^n��&&m���e�J��6�Q���zd����V1���n\i�Ŵ�6�:&�&�,�,�Ź�7=��g6�>�r��!�fˡeU���Wh$3�K��ٞ�����4X-ZCF�w��Y)��6�'mv��ݖ��ͻoBV{wnD�r���i�ٞ��k�`ˢ:�닇e��xn�����S���f��ׁ��]K6�r1=�ҡ���<�;nR��=r�k�*��j+S,��T�J����s6�읁�U��U�bݦqgTG1K]���p�/v�3WY}��m�Yc`��;�s�g��RK#4�j'eՎ"��n��K���VF���d �fa�t����t�����<�ܮ��\���rEٲ�sEHn/*���5����OGY�5yf�Y^�֢�X|J���
:�����R�jBU�]/vPB�/ ʜ�9�K����2��\�e���
;�KMe61�[�;�[e��C��^p�Yo-����r9���1��9y]G5�����^2h�mkV�v�3v��Cד��:�à��g��9����N�s��\�X^�ZX��E[�ݶn��ҧZܽ��ŕ�]��L�|I�@����Y��w4�e�Yq��a+n�P,���u���=bCiyΜ�yy@��c��$��<�F��Pv;k��yq��bI�u��,ڣVQ���t�C3R8�.�$Gf��p��"�<�v�[y�X�:����Ҏ���\喽���I��]C�+��j\����s���Sef�
���l�	�ܽ��nYk��g���VxcO.�vx��*ng�7e��bhl����\�,.��k=�]����.�I��$��;f%6�jYnݎ�nw��-t��k6�]"�nεI�CǶ�>�=�y����eb@
ƽ�u :ܛ�ц�R��!"�*����[^��H�y�d�{3Z��@��ժ�����yG�,�n3ʜ�r:Y��:�HK���%��E͉��;�M"��s�oU��o6v�S=t�&���k�g��Z�n��':ɹ�],fu %C&Y��̜改�X5�:�т�5�1��:`痗�w!ڴ��L����S'7b�.�{^�m�ݽv�pz�Y�hm������y�b���r��0�ÓiʖSa\l��{Q7n_#����NƘ�86n�e,�[R f@5b���%��C7MR5+d]6��B��gp�Wn�6g��q��,�X�ջr�V��.S2�g\cMc�����$\��*�׉�`��;et'M�D��nͻ^�6\�=��������Nb2�U����e7��K�A��#e��nHM,�����JJi�X�����К��9ś8ׂ�5jq�ٸn��.1���E�V�zݶN�xC0�s\���(����vݝ�o-�<��۱�������s!�'U�IY�@,�h��-M4ԣ͹v��<б���.��qԸ�5�%��zm��-�sI�ؒ���'%���^���=<(�k^�b�Ͷ�(�Yb1��6:�Q�6�#oV�A��/�LO=�W[��˹�d�kA���'& �)�mN(�+b��C-���JK+
*�H&��g��sTAVbTr�kgi-V�cu�j����%q����ɝL���p-�mѮry��Ņ��M�D��B�g:m,�����u�uu!�]P�ْ����[����r5ɮ����u��똝��"ݴ��$t�t�����
�@ó�d�˪�B\�K�E5��˴8z�`��B^-%����E\�8����E�Ҳ�p��M�Yn�w6d1��B���<7(�kNs��F�W�hL&gaxVgMXu�-���T֦ѼێF�;��^�[='�uۅA7j�!5���X��b�T x�=g�&�k�1J0�q���%�l�v��M�v��6�Hv�v��^�����C=c�j�G��mF��73{N�볓��lU�k	G"9���q0ݵЮ�Nq�<mj�{Ji�X��=vCZ1mO m6y�G\p�Ϟ;�Q�kh�]�8:�Ry3�C��q���{9�e� �к��鮌Kj��`�e�MB�d�y�Pr�mY��vu�ʃ�ٞTؑ���5�-ԫD�,rru%�ٹn�E�7V�Dn��R�R��zǕ-�%�c]pe��z����6�puk[0C;i�3uۀzc��nx��o!��s%�8��G/F�\�
�<.��r�λ:{�\r/���mLt���
�5����ѷ�n�s��\�)�ے�`kM�͇1��Zmb]qp��/���km��l�k�YC� d��!ـ�����٭��aL��X�nq�cc��:�^u��K��� #�����l.��;�R�MΌ�aL!3f�h2��"�^t�9k�G]6uVsd�����f�&������͓�5�n��Ϧ��M�u�å�����{tڷg�:�톲�k���7]��f� ڲ��\u��z䮜�noTt�Ʊ�ն����,=ql�P�˱�n�g�f���r�Vw0����i�Z]v�`u���]�tt���D���S�ut�$㪕�%+ֳ]f��J3�M�,
Z�VoGi�甗���R�K<�8�Xm0F0�c��fZ86,w��Mn(6�q���o׷�㏕��>]Դ�
�{e�f���QC��c\�Q��˃Y�+"�S�IR�X*�QJԕ+XW�Mڦ!R

EP�Ŷ��,1�AR��1 (j�"B!���#X�-��X���b�+*�R��5�(��n`W�Ȉ-E�l+*J�U�c�"6�R�� 5�҂��,(��U-�++
�Z�EE�V�Ɔ1`�(�(�U�B�(�
���ۨTX���&�m
��,8���TX9C2�@�Ь��ȰbDH�!b��ɶ�)/��(�@�c8�C��T��VAH��Y"1A�((�Z�*3�SiAJ�P�U���TD*V+�ǌ��j��"��* �Qr��Aa��c�G�KŶK�I�>�?=)V_m4��՜33cf,q�KX�� ۮ�ֹ܈��<��9��pF`�vk �'������ހ���g�Rv�9�[*鈎R\C��M�;#<bo3Ĳ��.�{v�½�셫��K]�ݣ��6�X�r8�W]W`�u�{ulK/S۷��a61֝�Zv���ژȰsf��⣗�f�=sJn[�r�A�I�DXK��va�6cG���K�!�cF.��Se*��»W��f��嚱�[��[�59u$�jOٟm����zƙ�t��3��h�Cf�]���X��S��*��>1�C��tMQ��q=�^�q���VPt�vj�7B���|ԎAݵͣ7��C�-�8�]<;^�\s�������:w]cw5&�]sk����ⱷg[����q�wW'jz�Q��݌����Ĥ� aoK�G�ڬ��y`]Q�j�q�0\�0�v���B��$m��L�A�3י�X�b581C��W[���tݸ1��ٔ]¢8�.�!F�y�D�Q�t��V�5�t����M��n^��S.�KsIl"h�2���h���,н�e9���hƎ.�N)CRR#kb)��ӛ����Ōj]:�3���i�bꥺw��k�"粉������Ja����<�� �aF.[�F�ٞ�W�Z�۵��L�<b�Ƹ�]��$�5��S�Q��#n�4�V7��&ܵ�9'�7Yl.:�����v�r1�����&s#>�d�0R�[����u�e�KZ�VF-b@�Q���%��Jf�
7J�Zl#]40iE��C���\qokن-�J�盵�N:�x�{v�<�u-#� QIm�������m�%0�eΤ46�e�՜�y��kK���g�g�g|]ڽ((����,W[ �X��Y���
X�K5X�mx�����Z��-��##��]���z��5�kb�[��؂�76���`������N��Y�-�B�瘥X����9q����*(<av^^����Ֆ4�̴�h����h,�K��R��F��*V4	iFѥ����� +��C=��9Ca�������BQ�	Z��@l�/Xơ͈�N�Z�����U�Um�+XB�@ak{�q��<
�ݑ^W�#e"�P-Kii%��z%�"uJ���l�����ϒ�a6	P�	�zI �E�I�Ӝzܤ�5s��W��	 ��Ȃ72h�L3wvf3'L\@r����:�2i��I3��#��րI�t����b����D�Pl�b��N�)�@-� F�`9�$��,���=��NldIˍx�$��ԓ2.Ar�z|��i�c��Y�˸c�v��	${c6��DUnd�Jl���3>�I�H�Jb�@��
� A���q%[y�@N��A �6��	�;� y�;�#ZM�E¡υn	nk-�m�[�4;R����/�l��ʒ�'gvH"��������'Aר�A��q��@��{����Rp4����1H���K�!�f���g���G�7�hׅ�F�e�4"籭]{���������'g伥���}�<r�i��)�xi�)�H�Pju�ˌk��ׁo��sK�OqxW�һ�� ����|N��'�d>5M���v35pV��:��Ґyh���>o�����דn���1�o�VO���x��Y �(=��S�N�)�Ai�5���h� d�%�7��$m���L���� ܧ��KRL[�K�p�|�>:Ց"Rjma��C��hԁ>�̏G�m\��s������_�WXBr�kL��7%�9.X�e�9l״��� ���Q��g��A���sF��O{�ƭA �m�Ąkvik�ӕ�4�)��k�ϲ�Yq"@Y�!h_��03���YnoKE4	+ A ��q ���2�߳s+���g�D�N��Nv�x�� g�l��G��HU<	�'�A���T;o�dh�<�q�ۥ⸸���z> b^�q��o�>�;���=�ލ*�a\�P��ۅ߃�n��B��[�K��ZvL�2N��2��:_(�i[R�͵�$	+ob ����� UX��e�m�	�q��o�n]3h�ќ����8�||�8nN�y��c� s.��I[[� ���|�{}~����C
��J�{]�az[��uZùx��G\�F����/]����A�#Ar�o�* @$�D�#V���}h�:CNU>ȷ��I&��=G���2�&N�2&|Q����{m�T���ku�N�}a jo
i�NœI�"B�����y� �.��` O��b���ȋ�𥻢�x��cZ	�a���4���8�����2zɠ��l�uc�@$��� сչ�5�k�����*�V�����y���1�7��WT�w|7ץ�g��{#�M���D������U��x�������透 �R��ު��t�J5t�t��,�k��IS��<SC�dC���'�o1 �uS�%f��ہ-�8�nI��].�x�Z����vc�y�GZx������N,�@�g% �\�Vq�N�?��N�N�Dz=GXA[���*Q ��D�y�*4��߿P&�qfnh[�H��6He��35��^���im3�%n���?J7^z�_����/�ΜCV�>Q��_ZH�� �v��5�fk<dѸր@>%N���b�4�	"Ļ!6�M6�wx�1u	!]�'�,��vs[;.^J���'C�iւU�m�ԍ��pŐhb�� �
ʸ�I�&2�ݪ�FG��F���2��#ĒUm�{��!�d�djD���yq��-�^�޾�xFp{��+�ߓ�?E����#:��U�X�Q�����Dsw����!x��X1<T�T�}A8d̐A��a�3�eG������Q��ܙ�͜M�p��z.
��GN]��LC^{gnx��ٰ&���K�>����?:�^C0s�c����s;#(��Es�\���\�!l.ʦޞM��O�盎�'<G��8�)�㣱� �n��:'X2c��C]A�,��\v9������6�ts1*���g��z�p�q�=;b� �a�6ܧW�kVkc+���F;e1Nq��9��8en���?___�Nd��,�p�KG�2�n �Bͷ�sD���M��(�R���H�p e�N�L�gE3�v"=ƌn�m���ʽ�zf���s�:�5ۈ$�n �Q��a���5W� ^�H��%˹Q��"�;�Az�c�� �)��M �D��$Vm�G�m�A�A�0I���,�^�>�k��.�'&u� �{q ��|e/8pa�����TM��	�)�� �!�� �����H鸈�%u�n���ʽ@!e�B�^:u��r�tqZ��3>�&���n��,�p�òʳmm�N�q�v臜]ti�b��>zC�&Su��׫�O�8v� 1k�G�VEN�>�w���O�>+sb�ʰ�;0A��e2t�� ��٩�S���k�E�EĲ��w���i�������?vm�\&��H�xx>��h��x���	�׎{;79a}�K;���X&C�;ܢ:{wH'Īۈ�1k�A>:%&z��D\%����u�wI���8�g $�h��;yy](*��[��O����{�4��H�,�r�r�|"6 cL�c"wS����!��	 �ȶ�I���m�w+X� ��}ax��4,E "o�[Z�<u��@��؀A�5�V/�����_[�N��:�wBH$f����9qr��3ל��ˇvذa��佼n������>� �!��,4�p�I�Sp���v��yO�.�Y���A���}�)�2�:E��C4N���O���ˍ�fܗ�A��� ��7�SK��0�k����̫Ɋv;:fU^4["�O䞷@o$���q��닪�у�V4����|��p]�&E��к$5'k���L���gu����W7��7�}��B���V9�Oj��k�o-����[Z�	%n�$	B33�,�gE���	/[+�>F�7�2�d�l9$Wn �I�ݢ��Q[Yo��u���e�4K����Ҫ�d��q�`C�3"�l4��[��;p �A6�ѭh���/E�)��sr�n�:�N���1\J��+D�Bk��.�Fs�hZ�iwo;fD�e�|�T�;xǉ� �K���ϖ��l��k��A��	�ѥ.�$�,䉐n6S�7a����c���&� =�x�1��y57j�k�2�=q��#q�I��r䁿�Bw��W�`jJ�kf���e��$l��pr�(; Y�!��2��:[!���10cX/01��� �}��H��6�7�m���^jiI��c;�h�ut���<^s�� |ﻙ������՝&7�u�|�}��{��Vחv�s�����N���ǉcQ�p]�p�g���H&�V@ys8��:�U~���3�גM��V�4n"��z_ϝ���Ȑ��RF�0�\�S��k��F-�ۦf�Ͱm���mT`b�����w]����d���F6[ǉN�0�gZ�"+:{KZO����CE���32&
:��$��E���,�A mZ�	�0��tv�i0��[�FヂT�$Q3� N��� A$�*�	�hM�6ֽ �N5�@>$n�b�@�\r��M�c:�Lj�ݙ��(V@1�qĂr��@'��k��R	� ��Ǣ�І߆j�s�|���W�i�R�ٹ�D����f��:��@ΰ����?u����AĿA�/����L�(n��[k�lz�i�����i}���7)�Y�L:e	[݇z2��5oc�8RRX�$�H8N�ݤU1���]N\�rru3����˖�Gkq��6��5��H#DZ���ۣ[	��&�A��t^���Ù�q=bό��t��JœXHY�����.���j��ݮ�U��;vy�k�@�K�&* �6�m��ͬ��F;
Z�]��cDԙ����r83�3��ݍ.�v�EEػ%�p]!���#T&[6T�;H7V�q4ۜ����)�`�u̹np��*�HզCb�,5a�p>�}�52b�[�}�|���[b	$ck��#q��"K��G��1� HMV���.�؄��C�����|=�t��%�����o��y_���`���n�D��p�����1j�J	 �|���c���t���h$�*��������,�Ȣěڝ��Ol5d,�"�F�I����P5�����L���zB6}n�r�tCy�:�DM5k�3�;������B<O����$-�
l*�E�RYߍ�wqX5�Ha�,�J�\FF-f�3]7nl�hǷ6][v���~��D��G[�Ì� 1$�]��O��-�f�5��f������c[Ed;]6�O��܁ ;�-�p� ��?�[k�A�l�`̈�E���<;�Ӣ�a�f�_igU<��ػ�-10��&+ꬨjOߺs�^�rw0�Qk)awg0�dy��wb��,4o~C0 *�x� E��x��"�)��t�ʐO�k(�%؄��C��U�U<	KmǠh ��Ru/���j�H8�n �%�b�J2��vfb`�O�'���,�XE��J�C��Ml@$�֜R�����ٗd�DG��!��� �W�\dA�$v�dF�aE���� AUw�ӊ�(MG�ߗ��F��y��B��L�ڄw\�����n��t��3x)wS]��׵��!R^�K󯯙�IWW�ӊnBg�kq-F���{�>e��.�쓲�:�bh���v��ͦ��k��Dy!�ϊhڱ�ZZ.Nx��^8�,ᝊA��5K�ڂ.3�3��������8|3����ޏw��������H�3���,�x�3�?n����s�;�����VV�]�L�˳&��/Oc�=����r���aO��;�p�D��nr7�a+<���|��oh�mS==��>�ݯφ{@cz)�l���Z���\=���9�I>:(�D���V�h%#M}{�����>��p��_$��ӽ�;M���ӞG{9研�!�e+�!�^q�㝴�sy����M�0㽝L�ݙ����oc�q��ݞ���j��;ݯ=��e~.��=���5{�g�_�����qHJ6�wR=tS���0z�͙�GÚUSG�ɖD�<d����wx�<�><��в>�W���t����=�:%�{ܽ���rީȁ٥�;7Ȥ�{ц�=�^���f�w<1A�M���U<�c�q�G_3���t�>�Q0m��)�K�qIs�G�ǻ�p9�]�n�����+�Y�2m/GN�Ƕn�V�n�����.
B)E���ܙ�;�iz}��o���kI���Rִ����zh�޿,�'�.���;7�Sp��\yw�o���{���b`��\�2��1vwv{�.�&x@��;�Z��T����Twr��i�{�?X	��q2��v_+�o��8����d�ny�л�c7������L��xnM�ް��׭��r��J8�P���z�ol⼴p����$TA�r��~x��\�V{��{�g����w��L�vb�vwX�#q�Sv-ۋ=��F�^�۸�=�l��!����\���-��̝��l�C$K��w���"<ޑ�G��M@����ch1_�-�Ũ8��j2�P�֢AA����m8�P�x�b�"*�LC3-�尭���J�ƚ:��F�
����K�Î�37%Me2��1S(�p��Lb�lJ�Ʀ9�m��e��(��*�)�u7��#<#
�xs	�A���X�ڠ�'��x����<_<���Scif�Щħ(qĊW�1����Z���6�~�^N+I;�1����x��<�sp�b",��c��E0�TDԩ
e�J~W��;�pJ�[�����q\r\�2�%I�`�SJ�3Vf=��`����@Wj�Y�t��L��ħ{K��;l�.�i̤���`�����Y�u�g�����Y@.gp�c8��e�Tmr�q(�7�rNv��/)�Ӯ=楉0�T�i������9i112���^Ձǋrx�%�Y�s!�]�s����2��fc�C6�{����٥���D�K<$[{�)�k:�?	�)2��VR�?!a�<�ubH�;�2+1U#mf�{ys�q㷸S,�q��R������c����ry>�Ǆ=��Y
Z|�����Ʋ�{����J�y�_�jfE3�C��DP ���|�e���~���P�%O}��!�;+V����I�;T��H{�Ｌ'�m���|���ac1���S�ߺS�~�^e�ݭ5���ڐ�5�y��c�}�!!�O�Ќ������5+���9�2�3�
�)���u:0+ �����8LI:2T*O7�{�âJ�>���������x���h9̓(�mg�5붱Gst']]�iT���[c��[�q���{����R庸�N��0������0�%��� ���}����,
%HY���e�% f4�h�j���ԣ�������i��D�lC����	������~�Jܹ� �P ���} �ĥ	����x���}G�w��V��~��c �
C��}�d� D ��>���m\dcn!Wc�(�#�y�?er�Gr��߉�a���:�!Kd,����r� �
ߙ���w{���^��9�����e��O�o�xLC�
�d�X�����aԕ�>y��晸[s4�ä��aS�}��a}_�}����8��
�bb��s�������T�<�w�C�R5���|���9�3�~�9q<����r��Mc����X	e�C��	������Ŀ���0��/{2b�S7s1�f)���<dS�xȺ1q�]�>�'��M�Ϝ&'FJO�������csU���rC�� ;�u�R���e�i����]����㓬��}�)���PvF	�Nz� ؃��@�W<m�88�^O{ɻ���n���,�N�K�f�v��{��s�j�N�5�M��R��ŋ>�����	M�̼=ć���;�!�Yl�-!�}��{�Y.���� ���1v�P;� �±��y���"���`��<�zé+����̷D���Ǥ���§w݇Xu9c�;���t��f<^�>�7��>x�|	R���Hv5!F��ߞ��8�}�H�]���݁��1��>�=�4|��J:d��ą���Ad?%M���!�:�Y�3��e�}�>����|�}&$�
����fy������VTߞ{��!�>$,�ݓ����e4G�x����1��c;�^=��!��B�C����d�
�`T�|��u:���e����е��(چ������Ȁ�Κy>�`V}�~�6�iw�Ru�O����%��
����N�X�o~��ϻ�s��`~�,���R�HX5��i���Hvv�-HV����@�'��|���O5ˬ4�)D-Ӎ/��j4�ؼy
D'i�.f�9b��^ͮ&��ӎ���'���͈�[�4 7���s���U.���>���g��i�,�m�)WQ00eI0Y���E�K�ʙR&���c%ƌY��W:q���Y��=r��%�k�Y��N�\7o)��B�[�m��!1�e1a��U�Su
�Q�7k��1�5]͍�S�vlP�T�W��S�MF���j+���)�:�n<�����4=Wv݂�8�b��[y�]k�)��(t���k�v��B
�L��p��X���t����S�{c�Z;v�=Ҏ2A�Zٲ�������h\�u!ϼ�8�� VQ�Y*o�l�'P���XY��ޓtT���s�l����ޣ뿾�$xO�2�(%M��D�B����[��;v�ft*C�a�����GYl��m�Z��4�_�TTA6G�(��@�1s�{�M�vC���N��t���}�@]�n� ���}��|4�|����[�nnS1�:��K�y�8�,��+؇�w�9:3XJ��T�o��˻����R��(�B�}��t�{d�
��s��&'c��߳���.�z�����0���N�<��q#�����
2T��}�dAa��Z���;�bR����{b^�68Ӟ��A�>���p�$�Gm֦nZ��r��	�5����묅���� t\d#@�w#j�{xYsz<:R��:��fC��;�<�:A�IP��
��y�yXu%`��<�|���BY���-'
\��h��q���lMŲ�k[��~��3`���'落�w�����)I�Zg����C��"llt�<$�<"���m�]�ϡ����~i��A![��|��bu�R���r�V�樷>t`}O�U���H }����M�֋�l�\*�U\�!U/Q���ƔD�C�p���RD��|�fA������"+���㣶e�|(�)����ŷ����w.�=E|_\`�v�6�}^�هx4Iq&I����	����t1��{߼�����>G�-�պr����I�^9�#�m��T�Z�=�~r���
ZC�<�yY萩X?~3����o3�����Y�"eO�wϼ&2td�Q��D���{�à����?��1';; �H��>��������f�-��x�o���OD*Ă�����N{g��/�<罩�!cY
�|�q��n�v\�~C}�K���|.j	�сR�|����>~ֲ�d�����v:%7�{s�'p����k�s���C����~�|�}IXS~o�����*J0��3�~眬�B���D�z�p�$�y7���w^,�M�����iak{ZFWU�T�&Ѹ:�u�n����z�kg���O�⩪���w@�����c!�B�H{ϻ���B� �7���S�
�~뵧>�f'�￸LdAa>����䕅������3�4s�RtaS��{��ì��T��5gL��r�(�E�tz�����*B���yڐ�k$Y
���t�I^�%��hf�K�Ě�����I�DV�6IL8$��<$� �:�*+ ���P�%M���ȝ�'Y��@��n����鸨�3Eޙ�(���g���\�b����oN�lRV\��)���h,ʅ�C�0J>x�;���(py�]BmR����j������yt���ql����<m���wB�����S9�!��B͙c~E&gMH�
�z�΃}X?~��y-����o��bB�!R��>���!��0+*eO}�J�
����߽D>� "=בЏ���>y����r�mݩ���O�>�*|��C����
�������1��Ǿcg+n0Q�DxfS�"<$G��d,��߼��Y�y���T��	;Y��C����˲K�V���\�t)���ͭ�R�0�[�As]
o�?�{�|�m��d�?b��Hs���VAg�R�z�]�w���8�����n8���"=ju��hm~�;�f�0ȔRI?_H��(Uh9e�2�vUT<k̀�K�5z{m�o6���I$OY�$�I�ۚ4IX�=�5�^z���Y��`�L�'�U��I�`�M�c�2'&t���]Kw�)Ѽ�I��"e[�q&BJ}��`�Y0L��Y�]��51�S}����	���3y,��L��w\I>��	g��z$G����1����F��u�j�,X�{ۛ����@��!m���%���:����t��}����s���=��78��Vw����zSd�t�In�H� -����@�Ȼ�����O��H%Q�g<��|QS'-��,��!$���2A$�;�L�b�G�h���h`Ί	�8r]�����:^<���x�h]<�F���5#;�,Y{��?X1�����Sѐސ�y$��x�$�Itw@�c}�z!3�o�ud��C3xn_D�g�@0�Q0o)iMY�'җ�y$L���Fv�u�_��J�2$�) ���@�Ypt�{"�z�h�������)ҙ��b^e"W��́@I��;	YrG`��I$2/�I3��lwH�IW��3��)�|�u�[7ӽ/{�%�b^&<�K$�o�I$�m�����]6u&�i��.�
ER	n S%��c�d$�J��s���é7v���S䗒Kcc��)"ݝ}+�9Vm�{T��Yu���B:#�s�#�g���<��-��;ǒִ�P��ba>^��x�G� ��g����;��_`�A5���ã���~��z��̥�V�#��S&�u��n�W=��"S��]Ռ6q���D�^���mW88yL+cǷ]nQ�.mn����ƹ��m[��l�x�j�y�b�$�G\��un�J���\�z�
���{qہ�7$�ɣ�(��s14�s��lkz�G5wGX�+t&��4n&�e�.�t����a5bzA��ٹ�`9m�!ֹ��b	��6ua��-��q���X�룰֨���\�:^�sA�f�,��ˣe۽����-,S�����y�d2I$�9�ϥ$�M��&R�F�3��̽��Z��Hw�'��C`��NX�tΐ`�U��Ή��ke�ȉ�#���1�Iy%�q�@�$�H۝"	%���u�m<j'�*�a���RH	�cL�RIy&�ȓ$���B��"w5��$�I�#>Iy7gH���*�j8�r��ŝ*��Ze4Ss$.�S��J�̉I%�o�D��Kc[�O��z��i� ��}ؓ"U��	��f�
�@5�fb��&�n�e{s�T5_vE�I&��3!W�N��'ҊK�[�HH[Ż'S�+���D����ՙ��նĖ9�[�iG�Ş.��Ŧ��m�`b���={#im��g����Q� "RM[� �	v�t)	D*\VTt��n�4ML��RH&��Ob.AE�Y�.�l�L�@ ��3����c����D��|}�Z4zz榥O}-���kD�ڣp�c�Bˇ�������ɕ0���ns��e݉��3Rm��T�L�_�������ݬfBp�I�wG��	!�/Ҥ$����\҄w�|�����A5��I� ᪈��J�K�vKdHd�I+��&�f��;��M�fQI-�~�!.�"n���`[�B���;��|�{�>^)��M��M��*RA$���<A��Lï�
H�4�)mv��΁r:UT�5�e�).�|2$��17[�q/�%Z�jd�I
֞�$�g�L�H�Fq���ȇ2|�z�"���k�9v� �茧m�v3�փ�@�+�?~����ˬ`���/�V�CJ�Dx�b]$�A$6_���IEș��-����.��S(�$�ZzX���ݼ�a	��3�	Ob�����I[�"��O-\�)$��&R;-ڤJ$�
U���-�x�j���R]h�&	L�wi��'�}�j[�H�I"<�޴+�mӋ�jf4�y!:�q
��C�aV&2Y���8�����i��.��H��i�4#�k�K[��3ӝ�B3,�&�$�Kآ�@yI��~�2�A3b���dΐp�Ti��n���u�fe4�bC�I$:�L��<��m�?�]J����,L�y���΁o)iMo���L�$�?>J��Qi$�:���'ƺ���H��H�Iy[�q��5ƍ��4Ԯe�9ٹ� �9E$T`]���U�s1�c��vfÎu�=���۠�bsK�?.��t�\� ���Φf]{�9�TIy%�ф	&wv�^u��.�[iN�ߌ�W���+IՇ	Z���.���S%�����uDt���{���Ht�I$���e �E[�q�J+�Fj;S4�ڒ|��	�����B�N�R�)�Ƿ�
RI+|r��&��8RI$���L���V�dJ�n�HY���ćx�b�����ӵ�ӓt�̫�-�	H$�J�#ϒ@ އ#����������b���q���uucU�.{}4�u������.��V�BG|i�\���>�+�zXU3���ox��%�>R�)\Zԋ:fL]
��]P�H
PIy/�fD���t�+�x�	-��S!?��d򨽑�I{UoK�K_#�9�[FL��&j���9M���t�n�+��H(p��e�p�Ř�n�Á.��k����csم���+w�S�K��bn7"���Ij��y	�ZX����(w�R%I+~�o�85d���*��L˒iX<9N���S^-����Hc�Ȓg�i��r'!j��|�%�l���Y��ػgb��(��!$����"PHߟ*�Y�6�I�;��u$����ekگ�^�B��!0`�?�g�TS�+;}l�C�&{	��U�&RV�v^RI#����c���Dc	%�"})x.�)�æbC�L��tȄ�IS�j�Mo�,VY8Z����T���	$B�^��[K_w���nI��}�,��Fr~�g������}>�G�d�W��6��SΔ�~�߶��_Y����%^�ǽ�t>S	w=}+��S���yx��pK"�����q<^������zY�ru�zW�8�o�+s��:̙��1��B-���۝7�t�g'��Q���랶�Nwܩ�􇦷�x�.�y�s�j�{��
g���F��g.ۡl�t��L���>˱?Qލ?Z�X����I���7���s�a���u��v�A���%��$��B(�k=�7/h2	�����]AD|)bB|/f���8}G+o�ݕ���Z�l��k�B[��7�N��*s9x�9y�͒F��6j�L�v��Pu��/{���{|��ټ"G�'�F곗Q���{A O7�q�zj�OU|h]����R�Ɠ��݃q�+E����g��Bz��������}W��͢=�}E��l�]���b���>z�[�R_yl��w�h١n�y#|%����כ�=��1L�-�*�ׄzf�՛�|�d;����p��C�j�O�:��3�f�ks,�Nj�M�u�s�|����=��u7��]�L=�� �:=�?�8����4�E�h܊/;�W�ɵK�J������aP�.E��`���V��{�¼�ӷ}�E�������HU��C�t��{���n���k�M)�{����+�͒�"�s��s߽�^���)���+��1=�x!��Y��Q�ׇc�D`���r�G,��^�: �{^����w����c�s`�=��'��ON/���^z�}�����<��(��$X���Z�.X���l-���Xq��]�����}���J�9jiF�?!��.R����q�5�b5#s73q����n��`&����LH���L�J�,�Lu:�ؐ�f=�<�,��v��y����nn�nҺ��P�9�«�� �VT�+hbV��.8�X,SPRQ�Ef`2�+I\c�0������+��bhʨ���x��CQf:_Ƈbkh�k�:�� ��No�rt�'��,	�x�
۝��$D�J��!�U���CPK�ɛC�CSSԩ��W;�=�Er׎���7s���:d�_�kKc8��2U�/U��KP��ͭ�N{k5�ҥ�[�R��@Ԭ�Q�x.g$��@d,a F2xRRc�ly��EJ`%�8��S�0Ķ�iPPm�e�b0�IC<W𚼫Ď�`���*�^�� +ў�R��Z��"���sl�ˣǏr_Vp$���	)�Ɍ��X�����Wg'ց*� ū ��3�W�����O<���W�)ܱU񕜵A�X6�a�c�U�'�}��ĉ�k5�hCL1��۩��m��r���9��"��/X�qbk�gk[2ssc�k�sҺ��oホ�nn7R��ǮL�>��t��U���Q�j�j�6Epq�:�\��@
�Zj�[R-Ɔ.-J-�U��bn�����B,i�;-l`6��n�@k����H�d�tr����W.,O�"����^�Y&�5��*{Kֽq�'��/F��k/Eϭv�nl��i��Gm���p�;z��M5�����v��u�w^L>�|.żA[n�$x���bM`n��/�:�k�j�4��v֡��n탊�Wj�-�T1֎4""V*��`�bAe�FU�M6%�b��0�9K�lU��(��ݒ�&� �:����V�6T���C�grl*gYv���uv�V$�[�Q���7��Gs�3�n�X�+D�X�}�]�9Y���]&ń&Gs�oq�k#i�4κR�ѥ���M�m�K�BR����Ӗ8nN��<'$ ��i�m3��eS5�ˍGJ�����4�A�z�n" Kg6}�6����s�S��/��d�E
�4��t75H�e��7-�l��3b�	I���f� �fWghe⃛lL�^.���[vƁ:U�պ1<4�����z`���Yw(����pn��E��Oj��	�G8��K�[��0��ٲ�N�,���m/�T��o\�S��<��t�m��q���0��:{v�U���y��t�qgh�����K)s� cb��-oG+���u�n�F֗�om�F�Q����ť�#����uӰ;��j�Ҝ9嫇cn|jz�}����o\]ڹG���w��a��Zŷr��-yS؈�7N��jѯ��$=��bg����/����ۙ�3�kl����ǁV����<WI�n���$�mO9t���uV:�t����:l=�� �F#��tF�p�j,�.��[���IN���"{6BX'�iO<�q�a����dxx{�5v�G���q�h�:��'Wla70��B����/�A��¡nZ��!m�G[����=�I�q0��מo<nK+772�]03W�m4�����*̋aJ6[3q�L1��F��R���#���α�r�/u�Nս0�xws�19fbض�`���<�k��z3��n�LGp�,�X�ϋ�3�8��X���48X���QM����n�&.���83��k.���[j���%������>?��L�����N��~I$���9�$J�?F���@��$�(S���vFT����&��^|����Jw^v?���5ti�D��6��L����a$K�gK�I#�Ϧ}(�M����gjݩ�&|тR���6	N��]����ڦ�]/$O>��2��YP�w�j�4]�H�{)�e��%^]`�k�]ػ;�iiJ:�" ���IE.������%+��X�٤6��=��)w4ܴ�%zxU�X"��,�*��E���J��'��D.��Y��j�i	$����2�	 �gL�����Ⲵc��|}}m�B��!z�������o��n{��ݢ�7��Ny6BZ��d����-��t{[�]NGI"i�`H�I.Ι!,��Tv�ZE\�rp�Ӳ�䗐	x+|�cbU�ԈӚC�x���<`�����ϑ^ի�� ;� s�{�k����綉���ߎ�F�2�Q�mR{����|�%������0q�B��]O���	��Tʟ���1;"@I$��lȟJ(>��,���Z�H���2r�;�-)�z|'ҐI%דey"E��f�y����x��:�� �Ov��w�B8	N��]���]�&n�>iK������î��M�l�	fI%y�	��CwK6+�';�"�4v�^��M��&Vb����N����y�[q>2���3m'��xb>���3U���>ԉ&R@-��(���!�������4����6��#��+�]@��oRY@����nndZٲԗfY��>�_Iiy����8M3���A*͘�+�/%л!���Zz��/���]��:nD)%}�"����	�k��4��y]�>t�J5��1��,F7F��M���ɑ2���d��ݒ��@'�dб4�d؃W2���`��.��UI?męA%��O� �J��<�s-�rN���W�Kwf	dlm����p~�v˓\���f��ѳ�?g���j�m�8>���iћ�TѶ�(bOQ��pM��� kM��$�H.�����>��e�%�4�vC��Rұ�dehw��4��"y��L���B�e�$�K�2A��\��u6���8��H^�W�ȱ%�����f}�H$���	�J�;u�^��$�8��^BD��"e{i^�!�g�g߷��˭�9*�jUws���L��q���n��-���qto�^��s85�v�߷�Q��>2���2�Y�"($��dL���y33�����{A_vȟJ+�/Z���%�tU���Ö.�(�L��D�X����,����2JIb��y	 ��#�(%[�KSj|�=���l���3+��3L�"�;�a$�K�L�$�m�u=;󽋠�H$��]��@$��F���U;$�ْ!ܚ�s��r�%�����	A���J<��Iz����L�[� ���n/��1�{��_b37��ݏ=U����Zδ��:{S�#�q��{�X������y�\f�U:�6Տ9R��ao%��Q���0�P��^�o{����?|�'��j;�A,y��9)���bA�~۶��1Rb�eBHrΙ�E2^@$ި�2�&��ʖ��r4�m���t]Â�}gnv,���hI���c�r���!�]3�7Rml������t\��;����H��|3)$���U��Sp�!U�t����VuG���ܻ��vwI��%��(%:0��Nk�&�$B�cL�K�$��dA2f����k٭rs4�!�K�,]�U�QF�Igd���$��,X���-��Az�|�H$�mF�>�RK���d�se$�̭�K��%��v�7bl�) w��"R�f�K۽R$�	q��z=0�M{�/Uц�WN�8t�8�*�.���$�$�卑"��{�=������F���$�ɑ"QI.Y=/)MY����Lt�Ò�K�]L�/��8��yg��(���)_^Ƕ|�����ǔH����L��.�d�V��6~���cMK<B�B���1��P�D�at��#�hͦQ5ٰ�B�M4�eq,0B����5R�IR�6�i����Sc��:����ѳ+�F'/&-ky��ur]���J�G�)ϷY�������n#�<����w+&��n�֩m��T��<��]]Mrd=���p-6��iR��Gݢ���)J��k[u&e`�<)��;f�/�<�fm�Ejf���ZŻ6;s`�]���kJ�jvֶ�ֺ	�=��O��9�AC|dF�2A*ܘ�� 	!�'��)�lU�)�ƀ�:4̢�Iv�ȃ7�Mh9A:.wcUAqər�i�9��c�C������	I$�66D�y�������^I��&��qS�tJ>M��)�8gtK��M��lT�T���V_:$BA$��׾�""�e^��K2:D�$�/k>t<����:.�Ȑ�K�.�,�7Jm��6���O�P"BI%I�e��Il?b�7t����ՒPWY�$J�lđ!�����4�	����y�ܕ-����YHezu;Փ�L�l$�gԟv^|�H�7b�J�4�vY�쎽�vf��;����H��pvRˉ��`H������f�:����70>>��:f�p�$��-���$���"	 ��~�2�FOr��N`�̉�PIZ{�y�J�u����wp�
9�h��Q$x��כ��OU�SA��i3bɰ��E����ʴ]Pdy޾E�	��� ͥ�bvt��伾WďYح|͵�;MK8�c��P�B�k�}C�����?��=���n��w�m*=�(&@HP�L������%tn���ڷA��8AݍU.933	 �7ؤJA$�D,�v3�L
�A$׆'�����(�7b�)	��
��ft�;�M��쨖ܑ!�˾�5oZK�I����`^J9�HI$���Fܐ�ݦ�Nc6|��â����r\�w��*i�i[�̐K�6$�D���x��ɵ�t��7r�D"I��Z}(�y�`O��i�9�{ai�E1.�L�	bX;�5Ǣ���8��q�,V�q�fhf�P�4ö�=z�"��������+%̅>f�(]z�= $�	!��"e/q8�%�c��˓)$�}�2�mM���d��f�]S�  x���1�w_s�z�H�W|�) �_�D/$Mu�8�J�����wPtm�r� ���m��>��^J��%���A" �� c��P6!�^y����U����{p���{��3��=ܠf�~�6��:�%��m ܢFw޸\^1�h/�;��k%�ȆQ���������ϟR^I� >I.��D�R����N���U9�R��΢�M��.Ze �I���	$������"�hY1V_��Nռ�%!W��Af.S;�M,J���(�J��D���۔'�D��9�$��L�	 �7dH�RKS�K�y�k�Q�'���� �!����筳��ݥ�W��i+(�5�e���_;��7�,g%�~]����YW� � K��C�I�wU�^y�W��/�̄�9�.��q��_ I%���Ι� 2�}]p��O�ƥ  ��!O���=g[�i	�V�lF�Iȷ�;�HgR�f,��b僱�'g�0%$O̉�$�J�2l;�_�I Wl��I{TgK�"wPtl9Y� ����ĝ|e�.���"�Ϝ��^�I2R&���HI����ܧZ�
v�0�s�L�u����(�zx���C���{�Y��<VF�m �=�no�a��eo��(K�>;��l?�[0�Y���׎:�}w�����;<*J�������
7�O�!7���N���@����L�L��-�0O��d�z}�J�Y{�&BK�o��>ʐA$��_�KZ���b��Ho8w`��f,�tS�{b��]d��\�7;\�sz��r�_?��3��I�?7$�ye$�W8� H$��G&�r�8���UsR$J.�O7B���{��$�AܗA��]�3�D�����k�]����I$��oҥ"R��� J$��̞qn:w.;.�H��M#BE$����iS?6̲@$���>$����cN��E���O��[�l)$	+��3)�WlŜ8L�v5T�u�R�k������$�Y��Ȕ<�d�d+��Gz�K�{$�s\"vrӔ�9�A,{5�g��������3�X��bi������ )I$���&B@%�}"G�x�;��-R<K�:qSUظ����Աma�;���xh�����&y�^zZ���v���',���ϻ�7g��0QW�@!=I'O=>��.	l���d��̹m2m�I{��љ	6�Ѽ���+�De/X��F��`m�of�8�1�vzz|����l[׎ղ���x�cHRڴva�v+]s�B�{O��w�mf^��=�lK`��[6�[��/C�n�frˢq��v\��O�.ד��{uًWa�O[t[];L�[<m%=7=�T�۰[E�띷n�3�"�S���k�tc;��iݻ(�T����\�L�ʎ��Mb�\j��۝���`K�3���-�i�d�H%Qo� $�HOgH�	te\>mD���ڬ�~�) ����ц})fk�M,]����,����A��K�8%˽�47B �H$��q�d$�Fw��))Un���[���D�a�4K"��N�3Ъ�S1fR �Sױ&RD�	��y����v�*$�W9gҫɃ$wl����`H��I.�"� Jn���*�M�3:���	/$�oFe���^I�қ�~��Օ��Y��@$��,̥�ܥ��]ˆg,K��fg����2�����En
E-�X׼��I	��3) �IN_H�d$�7a�T����:�ǓD���vL�M�����s��<���@ۄ�`:zYx��$�����Q\��� ���ۑ&e����>�
A-�n�M�4���0S0OGQI%9}"D�2�m����geU^]�2�����N�Agn�fx�DT��B{��~��^���;֌��<���_��E+��y��-�p��Z���*�i�������:\y�g=� �hG�$��ν��D�;�H��I%���JI)6��a)?b�몏"o��3Cr���K<6�:�D�����F|�J� C���r��4N+���y ���2�	n�tHbS�Ⴐ�%;�L�3ػS1GBU�X[fj�s�K��I�W�U��*|� �r�ʁ&�VƗٟ*d�绑G[�Ђ%S��A��I�fC@H���S -yBsT�:�v�$��$L���̇�R��I\�q�)��2�x9�~��/䧮�y�ɠ5��F��{qx�T���<n�vx:�Qf�:u������R�,!����]S� �H��l���	s��I��49�@��jQ�R �@%w��)�b�Ps�gp�
B��2�K6h6�]�y�2JI
�}�!$�I\�q�Ey*Z�]�Hϻ���hᒐ�޷3\8!��z���5J3䉹��"Q��&o%��=��l��������������ۣQ;'��'�؝��}r����c�_n�A��<IHx�=�����у}���^va]< 89r����'�MG��������x{�ڼ�ܘ�,9�VGW�s{�@r=�����g5�}�L�z#�;5gw��1�ׂ�a�!�C�h[��V�w!��V���/3��w�{�'�p�H�X�_xB_�jo�;:���֓�݇<�h�H֧yM���=�
�Sv�W�_P�{��Mw��F�/�����מ<�[G����ޘ$)"�w�����qtz]�QE�s����Ҝ�����5��x��E�c9`w��/���w&�����x�v��4i[��꯺����nM �|�%s+u���ޘ�՞���S�k���f�m}�u;FS(B5��3y�i`%�4��`g�>��yjui������&�{��|Mz�H�f�pu��cF>�^�#���
r�YW��;�1���o��U�>�~��}w["�N;��t�x�wX,N$�ݜ�����g���~���Zi��Ƥ�W�_b� ����yo��֜;��3��w���&�ԍ^��7^��Oh���F�4��ޤ�OG���˼�xJ��qT+�_kՖw�A�Y�����t\凜�}L��S�}2����y��vk��|BԖ��D{��[�ĳ�X�μ]�v�瞆vP�n$шSu�~����kq�����׷S�p]���ilk��f�x�{�-�'��^���x�案_1;����_pN�]�L�����h}|�X9 #�'x���[�{���������/)�ߟ2���	��G}Y�'��������:��Aeke%@:*~)Qg�jII�b�E1�[q�VV�����1�*T�b�1��N3n\I�ƒS�'Z��|TH`:���Ci-e���%�Q t���� m�t	�*wD�YUH�F,R������9^�`r'� ):���0����k*��)PiB��F)kb+YKLL`�����-�QH��J�iFV,Z����%�
��Ԫ�(�Lk�;�,��l1&!�̬�X�+"�v��� �Y+�5���TP^8�*:�u'''�I:AL2�,��2��p��,�B�UdSP��+ee+F���	ܓ��V@��K��2�6�Ĭ
�u�D�[NId�s#
���:Qಲ����((�+Sp����r����FF%P+#Z@�
�+���Y��!Z��ʊTZ�VJ�T�h��h�u��:�.,� H���ĔV1�m�w����E��y����I^C}
BI$Ϫ>3){3��K���wgrY����Ì��3a�
���Kw�Y$�ܧ��H)��.08�i3B҂K;��)!Z7' �պ�8��ﻱm��bp���<j�]$�ɓ�RM:�*BI$l�G��"J�� My�!�!�'��f���G�����P=��B1����bn.F�n����L�',·�����v@�n��M�>d�I,�|3�I$	GvșI�jq�9��6�(�d$���2�;v�ٝ;�gpħ(��e$|o�]��n�Ǩ��k���2$�W��L�W�)��D�E%Ο��#�ЩC⠀KӚ䰰����*X�6��)$K��H2JI�<�w�8�ky"R�~�2�	$�l����n;����쪩vKL�6�+T.G��N�3-4�R	$��3�I$#��舴���D�zp�''.�RJ�ޑL��f�����K���R�K��ӎ{6E�����l>��c���U��;\m�7����DT�(=���|��	H}��]���ݝ�g���tT��J��F��	k�E�H6�ʙ��H�}"}(����T�%� �7K��[��b��	'N��Eܺz��K�;Wn�v]I���I��i71�-�dhK��������tX�?
��qA�����V�I��� �ϯҤ%���Q3�]4�Exc3(��dS@�����wd	f�L��$��]{n�E��oB�kS�l�A%��L��7��"_���u�����)�UlΙ���"Y�D�w@�s�tf<J32A(�*�!:x��~�=�^H��@�����L�R^�aa��>vw�R��Ζ泥���k�I*�Ȑe$�J��$�O�D�&k�bd�܃) ����`�"���	g�v[�M�/2��K�2��H
uV��X<�- ��ڑ3�Hmfę�I"���@�G�o=�s^�ǡ�7L}7bc��k�����$�ۭ{�vk�b��8����u����yF�mvڣ��,�e��Xϸ�"|�x�V�JE�h

�H	HE��{��-�.۪Tz�	zw�^���>}�q�v+��`�1�n�ٖ�UE�w7����{<\zU8�6�|�<�y��ц���ԋ4��`��0������uY����bs��<i'"�wmuX�m�:����Z�۶�kCH�ltvڙ�S����Ԭ0�تZ���v�d��$�:�7Z�g�Ee����,y6�)e����Qõ��v��v}f�{�얛7e�]嫖@u�|�GW�D�֎�ı��Mv[���L�3;;;�;�O� ˈ��WY�%$��}�2��m��7g�"�I�ؐ��F�"��g�g�U�1�>���U]4lA�&*�l��FA"j�^��I���e��\�V���ĻS�*�)c8�����w`�f�Ͻ)$�N���Rw$p%{{f�J��)���X&�^@%�}I�$��g4�)챍��ݝ��,�@o]�Kn:2��ȡmאN�c^$B>Iy']��!$ �s������d;V4FIx�!%:Ø�|����%{��d$NG>J�b�)Z�˷/ρ�򻻙2�31�;-"_̙$�G��=_�oPv�RrX7�p��x��%���h�:�e��BcKA!��f�n���~�����,����wyn̼ϒA"mE�A>��LJ�~0Nͨ��g����I,h�i����ٙݓ�:d^�$��2�%Cσ�����0
h,&1;4��d�����&����fo\��Σ�&������k)���"
���[
d�"%�:%��l'V�'��i��AȒ��K�܍���!(@R#B�@"R
� ��G���jI 	!�GkL��A=��RX��;�����]N�I�2
d��3�I�D�f��}%��
2ߥI �-G{ss���	 ��u�Ҋ	 ��yL����
�v!���e3�<����U�4�1���	3���;3i<�w->yfC�J�5�	 ��׃��7�Z����߉%��B������[�\���
�J��d4�$ON�Ą��A�~�l���30����I�kw)��N�s��S'��a<+�2ɍY��P3�vdm+�AD��j�jB�{G1=2��l����Q�eu�/�uh�\�(;�%����-BD�5�Iy%��Hۑ*S�s&���'�j�RK�f�L�]����&�g��U_�l�̤�Wݓ.�gL&���h8D��Q�d$�C�:$�I%����Nn��Sg5	J�����˻��Kʔ���T��U8��I/$��y�z�q��
"a��E>���t^W�hQ�=�O����ov�'yI����w�_ocί�dν�L����'"B�U�d���> {���$�H(�!y��3�-�����Ǥ��_N7Х+�D�gNᜲL�&���y���	����Y�[ �,�}�)%$�y�Q3�����~$�͈�آ���U�dJ�XJF�v$���
nm��d�'�N4��-=b*m�ٺ�3)�u�T��H���2�:���g<�B���ʳ�'��gx�����R�����w�����a�q���xL\���sp�8gL�\��� �%]=|��Kg"Y �$5�y�R1T:m���WR(%S�Ф$��aa.PgtKK]��)%r�1c*$g*��"u���@R�@%����$�B_+���H�*V6�N�L����K��0-���]��R�S3>tJ	+k�h��I!���q[㻰�<B����K� ��y�J���.�����v%�JL��=}<��p�=���$sUq0��7�!���2�	�|>��>Ѡ��
�i2e�в�z����A��x��R}¸�}�}� ����ѓ��@�Q���a�R�1ަ��亪/�W �0��������J�J�J"R*��� ��|���O�/!/�mQ)�Ӹ`�S<����y�J^	 ��O���Zo�i<�NV��t���I ��q�ҊI�Q�eGF�
ѻm7c��b��D�vYiKQ��](qon�/f����30�V�e�CϿ�^�Ojv�*z7���Iw4�>I$�eG�$���ws���V�.�)�������c֩���vEӱL�K��$IUwO���Ůq���g� �Iv�Z�$K˲�DNY��ˊ�J]����/M�]H����ii5�T���$�?@�d$�{I���0�o�$�9͖�J($�gdɒ�dd�^,�dh
<_"!w���X$KcF)��H��{$L��\n�ꚵ�r��fI'i�i�� +p;S�3�wpS�'~ؓ&|�����+is��p�$��^��	��̑>�RHr��rH��K��r���N�����zi����j���L���%��43p�᫒��Ȟ薂��=ܻ���{W@�V�i.��M�׭:�ל�Z`q�/��R�ZP)i
 b@R�h �Ӥ����v�.ZV�:��c����U��������nwm6d0���a�,�-��r��ON�^,f���;r��j�u�g�t���}�a*m��f�� �nY�3jY���aLV9���ۮ���
ع68��5���m�.��r<����X㮰׬��#�a�ݘ�OmWO^.b�Qn9y�3�<lr��.ɲ &ݺIs&v�K<l©c��GBs�ͷIɵ&�`��;Z˔52�Y�t��)�-�?������3FL�3�5Ŵ�H��or$�I$�]������ء:wX!�wL)�l�(+��d�%#i;�ꓝ���%䗴�f�Z�um�	![�"e$+��K�K�.A����/M"R�I�����Nƪ���\O��Iq�Ȑ! ��K)ٶY�A;�s-��u#��e��Ƶ��$6������3�%��[���z�@�_��o%]y%"p��<���Ak\�3�vmݍ��á$f܉������NvF������S���'�i�1�2��>a.��"��(Z��rI:��������a ٶL��p�їʆl�zt݂v^pV:M���ۚi�4����Hӳ3B�S�8gg%0/�������	Q��H$��֌�L�L��K8��{fD�K֫:^R�TJ`���&yK��Ze/$G�����[t �H�
��'�<�2�T6����<����~�=�6�==�T^c�-��ic�wQ��4��k��㝵�玱��<J��()J�B�*�����Y�یc
HZ��^RI%�F|�%��`k��1�[�T��g�R4�rRv!&��b��"	I�e �;9]��	�3�ɪ�L���에��G��4�]qI5]�9`�L�S��5�+V�m��,���>��H$�6�4�I%��] �B��a�t�@Y��y	,�7%��)��gtKSSz�I��k"L�1��ݮ�$�'ʗ��IMq�"Q^I�}"O��6	�/��{<vΆזԚ�8�-�	I�C[�;{k���|�u�;t�m5n��_}�}���ş�~���UH$����2��(��/�L���宵�kZ��yI$��~ƙK3���vfd�`�Q<�fR]�m�lfܵ���ر	�H3VsL��Iu�H�g�l��6`����z�K�l�)�wtJ��U*i�i���)*��%$G�Lu��e�����TG�\�d�	�t錨���j��篮�<���w���;|rx/�����	��,6�u�������奤B���X�
)P( ,�
?y��{�������7���1�u��&W,�R�rS� �D�='"�LY��͛�7��de�|%'�1,7�$L��I]].�.vt<'%�vkw�Im�<�C.-&���,��Jc�'��	$���H����
�Rj`^Wo3�R(,��(�����乞f��ϗ���w�/�}�f��c��	�.�]��qX��Q���mp[�95Ҁ�����IVw!��-��ޝx2�J�rJH$��;��f��}��������%��(��T��$JC�kHG83��aI�Lv&dBIv��7k+��_b^D��J�6M�yӦ�]T��	5�o�L��ʻ�X�Ա-�%a�@���`������9�D��Kȳ��"imoUyߤ$JX��$	Q�j��yI
�D�E��(:g�Tj�y�y],Xs<3��y�wt��"A�I �(��&RKY�[�@H�1���R�[Ї��"m��(kkI�H�j1�)��0|�tm춼�<6�{�g����O�{�l��e��w�k�Wh���~��uビ=g��@S�#@�J�� P� ��e��~���g����&`�L�/��0�@$�=�H�=��z�z�#T��z��W�I!�Q�/>I �	s��ʽ�ڶƿ]�h.�õ܋CtI�m�h��ִ�t\VM����0�[��&���)����yݏ<�GtH2���W�R�	�H-�יI�=Ƕ��`+ʆ��Փ#���KTg_�	�$���{@d��3�%�[�Y��"R�IPx�s�����ۚ��?��I$�Od�2HC6��ДW�n�W�Нݽς3�}��#��P�4��p����$�;{�d'	9�,�R����38#@Io��S�K�	$�Kg9�R�^h�i�����`���%�3.qM>;q�'�	q����^Y;�2A$�t�v��⑛�{L��VKO�^���d�E��(:g��'��:	d���K�E��"[a�I�剐�	\�<�QI �28ȕ~���W����=^>�g�����=�W��褣d;*Ș���	{�y��m���ٮ���x=�؇��[�?W�Y�A�O6�5��W��+��N�W��s�x�-v�H��o_�p�\O�I�{ms����cpd�����(�����o��n���Ѳw�a�ۋ��w�[��8=6a�wec�:���i�}6�ɝٯpxlMf�[-�r��}�w;�B]w�&/?����Ra���&4 5���>nt]Xp�|��{ܖ̥t"{��}k�q4�/#��>/��} �wz�ە�u#��{@��ӽ�Q���c�y��^,�{���pNYu�s�c82����N\%��'ry�e#�ǖMas7h�r����iG��Tq>��wy�D��ǋs�����yg`C^v�A�j��KN^=:�h����݇��=���<P{��w��kW<g����s��!v9��jѕ{(S�w�<�f�ʎ��:t�4:���tk�l=���K�	��P+E�~;<c��g[�u�aţ{ŭ��{��V$A��yz7���|׏��R�����[`λ�<׻�f�9�Fy�]��Ny���|��=�'d^G%�z���|��zv67��OS��`;�o=�l��ʬ�8gpW�����'�ݛ�>������Œ_c53�,p��{\O�>��*����b㫳��l@�׻&�"���p+�^����;z���L�M�-^DQ�s��ƻa��@��,���f����MC.�Dz���C�x#�Л�O/\�E����bG�=nzw��"Y�C���T��X����N����k�OOa�Sy�D�H��X�$�XS�R��	�x�+��r�P`�d1D�TYm[cG-�Pb��ml
2$�x*���&"a-���Y<�c�Rr�t�1JN�s�+��r�s	I�TT��,�F&�k�+&����������Ke�'$�
��rp@�G[c.Z��4f��V�+Q� ��f
��մ�D�5 I rES�'"NN�����
�H�	"B�Ċ�t��"�1�AE5�)���$����*b�YsK��%h��R�h,Y(�u+#�$(�1; N�Rc�(��D�pqG�I��U#=I�P���pVD���X�5dĘ�PP�T��J�Ub ��de�� "p�@ Ѱ++.�Ep[���R DN �Z�)),P��8"H�B!$��tZP�@����n�W�������BT;T,"Jt@�gη�k�1�+��(�Q%m-QV}��h�s��ܽC8f��\r�s�*j4�� �f9��f��]Z���޹��k���+Q�r�ꎮ�ˬ4 %&�tn���wlƺ�$�V�aΖ.郁�-.������<d8��,f��7ZEV�U�Rf�j����.%�"x�����YrS9aFm���YfK���eɨL��%Ƽ<�����]-���K�$��S�,�e��gM+<W��ދO-ڎ8���".�v f�uhkm���b��[=��7���F��%��`ԯ:"�ur�RR��啦M��n�J�WX�.̆1[J\%���"I:��g��*\ŲX3�mV+�n��:�������4�Mw�G:���f����Fu���)䃱�[-9GD����P��X�P�n7Cˎ)<u[��`NXS�V�����Y�q)X�6EY��.�ֶf{cy����q��(�͑(J1�v��A�<��#�9�\�9�F8Ϯ�n,7y�'�y��68��.��=��=m�|7a�;����OWꌛM��wn^�Lc\�l�2�ܥ�Z�G)Ef��v.�7W��%�3#P�Zu�W!��Nv�Y�����[nnن��q�� ��0���4�&�7Uy�ek��s/2�"���h�aanW�a�E�*�j�]��2��1�ɖ����8�6��n$*�4h�F��:��J��;��K�}�WB��mka���6��f���`(-��)W�d����&ǭ�ݖ�s�0��5�Ea6ީLrl�]u�u�îV�:�3�SH����X	��i��`�㯜�]��aSh7f�=m�Vd���fV��S`��Z��W@C[`��7��ܔ�ݪ{I��γM���-�l��%v7a\n�rS�D�5���M�Nyv8F,cu:�����I8�Wx\ۅw]B�Yhd����,b7,vئ�:j,*��SDf0׌Gע�.v�+�뮮v]\n<��t�X�Ɏhy���j�k��9�Z���|N���p4�)��J��x^a��h@�� ��,� ��U����i�\����1J�,�]k�(�Q�1!sh�K��0pd�P�m�j�����1�N�+��n�Hou����W�cr�<3���8�of�99�v;p�c�}�zL��e�حt7V-��UГ\�i5��.��I�+gn{S<�3��u"n{YKm�b�-[!�qT���[g��i�\�ۚJ�[R��lݹ����c����]v�e<�(×�c�f��2���spp���fܖNz�p�)rj��z�q� �P?'��H_�����@MJ6e�	ro^D�I!ϑ�I9��g^L�����$�':��RWI5.��7���RQ�*I��|�,V3�<]e�Q�ֈH���d$�<��fQA-#^-A���YԞ��$��,T2w!��--!&�ן	I�F�O��^dv�^����.��˾�����Y�o>�PI-���e �l����� ��R�[3Zb�ӊ��Du��$Im�y���=�bRI!����o"�P�e�����g{��K�N�"��엙R��*�=�-�$ʩ��1�L����IytfȂg�m��iJ�^SO?��;�}P��۬�	E��<�����Z�Puq���A��K�]	�P.�y�}���ft���k=�H���J�vO�^K�OCHJ�M�[��1
����ւe$���2�6�$)$��b�$�)�GL�D��V�o�����)��݈iCPq���X�\�y�8q�n5���a%��]p�A�F
U�;�&c���������H���:׋�9���O�����"�Aa�r�9�>v�h[g��yӽ�l��~�%��D�%���[�Z�n6JU무�i�3:�f7v�GdO��$I�cNCI�Mj�o(u�Cf���As�H�J)$:�zZR�Jm�����i	۳[;'o��3�i<�$MDtO��%]��2��խM��DMj�]$_l�R8l�t�N�]�U��fC�^K�V4�U^!oo��j�D�w\�&BK9�%�%���փ\�����u.P�N�����9v�9���E�1��5K�f%t+k��f�d-g������1}~	n����H��;�$�Z�z�!&��RNd0�w���5�o\�&R�S�Ғ�r�fE��('g�T���ς[;��g]�U����xƤ�H֭����H�׍ J�$s�5Rnx�k���Y�Li���e���0�u�H��I"=}�XV>�9�m|4/ݕx�V�^%�j]z����gptY)0��)��b���g���K�q��t\�d�ŵ3�n*��Un<eUc]4߬m�g<�xCĊR(R	@D�YH
�9���KV��;�s��7խ2��l�5&vd���j�(�~�Pe�=�Q0�jډ�I%�ժ'�$����sNO+�V��I!t�2Ҕ�S̼̝�g`��J}|�BD��D�ȱ�]�~�k�`$$Iͧ� J($�>t��9��x�Sq�V�p����.���]����,��3n�ճq��]A�4��;[6G�����r�;�`Ļ��ṫD��q���$�Hk�H�J��n�|k���2[�Z|����WOҧҷ7����wt��Y<	�U�E�(%�U�, ��uӏ�|�c�/$��k��L�b��$J$�CUfK�p��活�]̋���N�"OS<+�D�GD�%y-��Tݰ����o6��Hܶ�J($�܎�2���"��p���&��m��94��*�s�&�]M8�J�$�%}="e$^��(�o�l ��V��㙗r���B��B�W�c'����pO%/x,kO���\��f��y������y�6�_z�]���w����B�i�J�fQ�(�"��R��1gm7�]��4����;9!��
�J~��@2�D�SdK#8^8�yn�Ml�R��D��c�/O��+v��HJ.��Y�/|���wzifV�i7�K#��]oro;d�;��z���m�ed1tA5}���2r�3�,i�l?b�)$��ݯ� �Iy%�Oҥ!�|9i�ւ�lc�sϔ����P���Y��'җ�^�vfwN�AvTN��2�z䦑�q�m�����%$���dL�N�7B�$���i�>"��շZ�){w�a��.��yy	l\ęA%�i���I�k�6�'5��:�"W��l�&BHn���I�y��d]�$Rt�*�sĪ'��Puw�$Y�q&RH$�u>ʟ$�1�ډlk�7��]�� ϭ�	�1wdX��&�M��*QH���S�V٘�N÷[i �����2^I�~�b�I$���L����"��_J�q,�z�����OF���L��o;0�����[G��H�|�������mkŲ�-�3���0�y���[����7t�s�� ,P���@B4%JP�@P,"�,�Q���Bݼ嵼K�n��71��7qe��>��/=q�!�j{Z�4v���<��:0�\ïm�u�yƓL��n]P���S�J�V�̴,FR���f�n�i�=8�S�ك��6Ѓl*:䖋��t�ْJhl���b릶f֊&IɎ/j;v��6jX�Ol� �^1��ۖ ���u=�<���c:G���;*��g-tka�{8��v#9���Pv��Q#��c��D����>i�d/��Ҿ��;����f0��(�ؐe$@;����K�Ϝ���W4�B펑2�I�~�!%����d��g`X���,��S)%�#s�z�]����C��%O�^I(��S(���6����C�鮖��5���l�d�gI��*�����ϙ IG5�D���sC��N��K\(I�\ת$ޫ��gI���.�����L<��D"����D�j�$�U��H$�J)��ϒI%�!�s�7S=�Cy���藹Dϫ0M��;�H���Q�g�bRI%y�
�l���D\I*�j�) �Q���J)$�G-Q+�j��M�g\�Nċt�1.�L�'�f������FX��������M."�-�A�vdMa>�t�ŉLm+]�82^H���S�D���f|��SfA�I�^�趸D�K�7c��Rز��&p�Θ31�%��)"=a:0k�؝]2�F��/'7�Q���::�5B�O]s�|?�~rv�G<?e��o�o��.7E9���M5K�ue����i<�]u{��{��B�(%"�R$!o�<���w��$��G�d��� ��D䨨���*�&�[SY�r�����gdg�xy��<��5�ʖ�e��:�a��� �ޜ�H�w� �{5�;3;��v#�ve��t�f�����]^�H5n�`F��I�u�[q���cc�2d�{�00t����'��4��`�����W3ج������;]�� ѷ� �ìn�����갰K�Νݙ�r��;�|��P�-��V�a��m �9��Q��k�ϓװk�Պ]?u�dI$��@ �m���C-8i~s�WD@�	����Ր	Ν��)�S)�zd������/E9܌���$�M|ޏk��ω�CI�m���Ύ���YEӹvgL������;�"E�D�I>��H�'{i�Q�qnL��ϸ^����s�{A�M��kِ��s1TĽN`�۱{cr��ypl�'f��)��E��c{nٶ���<4�4�J4L�x���L����o��~|��|J��KZdC�NYj�k�Ҙ.��!��8��^H=5�'��c���$�v:u�zN&�k=���	�u�6U�vL�L��=2$ O�FND��)ێ�;*�I6װ	����~���$����m�l{�}��>O/�:��Ku��.	P�<GM9������Խ�/��������۾��a�$���Ȉ	���I ��ӳ �nu:xvf�p��L�H���;7���ӻ �r� �T�2$�{���a�qq���M���O��rgĒ#w���A^\���f�St��c=����H�wfd�LL�6�̀I�%ղ$��b+�rmˬ���G=�H�O��N̟tYW%Ӗv.���b��K�܅��!Z��7�	��OLߒ �N���d�/4�|�ӕL�?��������P���M����+�a-k�Fv.�� ��M�R��;I����hur5V�݅82)�EЁ3YNck��W�R�H�(�B<~'o/�I�ۦ�ȇt�8F��I4[r�~��A>N�3$���Ӱ$��������)�_͝�Y{R��C<�^ں��P'��Z��]I`�t���k��s���un�; ]�wd�̒H�'&Ky"F�g(0��gZg.�ߢ� �����>��M��ٓ��
y������I���gC�ӝ9uI$����$�f�P% a;�4c��/�Č�%�:L�Q)�ϣZ��$�l���_-P=f��g���P$�뜙�	��g$c�4�%�ٙ"S1S>Oӳ3n�p��|��`I~��'���}�}-��nUE���zO�8��Y�;�w�fAw����{�'��Y�Pf`� ?��\ϻ� �_�H>���y� �k��4�m�Ì;�D�؟N��\����L��r�1j`T'��@�*詸˖���Ω�^�o���js�cߑ�x��o�Xۼ���b��Ҕ�P�E�{��ft��L0�.��m=���bAO]�胏[U@N3�n6�u�np�a��%�kU$m%�^y�l$m&䭈�v��'n�S�w
n��֗��# ��lئ䕆�\�����n��;-=kt,v�2��mYF��ks˥I�zݐ����k�W�;ֆI{BL,4�l��h�e���5��#5Jj�M*������z1���I��[�;@=Y�u�]A��V�[@�eb�\��v u5���|��dC�D��"}����%�P:��`����$ۥ�d k��D�H��`��.��t��; ]��F�a�m-�У�N�e\^� �H���$�s����%hd�&����~���M��ذt�
i�v�&C��zG�ȧ{�➎����'�x�Ϸ�>&�E	fNS;�]���3�r1ldV��e81k�|VG<|	'��{2	�%��g�{�b z��^#MDz.��"Yݘ�E&
Klt_����b��D�슳�dS�Q�zx� �K�d�$ޝ���G^��;k�f�;>N�Y-n�]#w+CY�n�u�8P�"ͺ�i�Q#�Ͼ��߲���wp��x���|y�r���Ӳy,�0+K�x�Q� �M=�L�'jm�1�'E�Azdq�3$x��#�����P�˚߉�9%������S�b!�!���g/w�K��"��6{Ҙ����.����b����-����/)�%�ূ@.w۽|V�0g^s���U��q� ��r7���H��7�'gv)�� UnTL� FeO����_�;���tA�$S���$GeG�y��%�2`���95�����!+�X,���H䇈!GuH�ݲ��N�6��� {߳��t%���ܣ�o�����l<��~��v�t��Ƹ�Vd�"��fw�G3�x�NC'x_a�B�)�G�;6���s������rp�ss��g6����5�.X���H�.�2E&�>���EF�����5���Ӷ����]�7NL��|r.v}$m�T%��w.�Y�̂��IU�;��c�j��{n�q���덝� �H�}�|���ֆs1w�}5Sn�.;��}�N{�;��wκgc]e�x{fr;��=��g����z=�O�hݥ����6�e�#;&Hk������Nt'���:z��;�j�Ϋ�����<w���x���5o�G� k�^'�J+|�dZ3�Tz1�4f���&K8,�#y�|��o�{*Ʊ����:޿������i>��|�{��k<c9_�!����{���g��;$ӻ ����]��i�-Jc����|on�6c��IJњ2��<K�[����۵F�~���Xlj�/���/t>`}vo.�=z� z{����o�O�y,._94GIZ���}�������}c>�=����ycݤN����=\\��f�g�v��t������*y�b[q���=����֎�����=��6��/u�}�!��=s����G���v��xxf�ۇ}݌��@� �5���L~�&�grr�w��|���֟}��s����*�pf�Am�P�B��Eg";s�j���!wt��f�x�/zJ1��6E@�>"�y�z�z�{���>>��G�����{=�oN]vw.�=��������|T���7�]�����a��{!Ǔ�7���A�5�c�ٱ�Ri����{n�����L+�J5��ۃ���y��ꏌ��,W����>����S������S}(������C�(����8w(y�^Z8{q����W��K���ߴ�ە���h'f[_W�d�z�`�m^J�t}����z�w�v�@ȇ���=�l�*��
{~C����Ҥw��Z� ����Gk�3���7��ۃ��)���,h�����2`��\�j�G�`�U�"HX
Ċ�D\M�:��3@�FҴV%�T(���-'J���%�ĵ��0�l�f�Z(\�CQ���8��m��Ym"�R��lVE��'E�I�ml4�:'�rw5"2'f["V�#$y�*��R%: -��V!��,E�YdN��
�8��kIXW������+ȣ±�1$"�E�$��� $ �yE"rI�u: � �葅�c�k�8�@䘚��E��a���� ����8)9��9!X���"��P�eF=¨�� JF��^!B`�2*��1��ADE���YeA�بŁj�[(G�K�R(�Ie{�8b��[-y���/FB�FD��`9:$�$C�=	�	�0H@NTN��0(��(�1���X� �3�O���������.:zd;�}0m�֢��0N�aq�Oxwͨ�����tulO��#��L�Ds����~ݗʗ��H/�"o3�r�0.�4	�S[A�A���U�k�[6F�8� �s{�$����A#[/�Ku���P�ju8���nБ���x�q/U�ݵ9�>�(��ϭ�ms��0jd��&L��w�K�ȓ�Mk�� �G6_L����0������ sۈ=S��!��D��g�A�o6u=�$�R���v$3�`_�"	_s�A ���[����}�����r��;�f3 �׀I׹O�{a1(&[B�O��A'���L�N8f,�v.R>�7�=L�T��߉�zx ��J^�"Ao{�{�cYJ�IS�Ή^�Է��}����ʂ4�7�7�����7�	�l��k�o���a�F���>Su��^sB�:^��z�L>+.���������v� 6�k�N�3�%�D��L�$��2!�q32�=�5�-S. �-�� �Gtc�>@�m���~W���r�/2r�kz(6�m4v���Z�U��n;8tK6�{[B��wx�d<|D��Ă	;ё�-Xcv�\Q��q贶�gċ�拢��ݝӱd^� y�#�A�����i�2�vt[�"޻f|I'z2�򫞒�q#)_Ih�g�t�'��B`S��� �O\lA����Z�|�9@�+oE�H��ɐH���EHr�\;�3�_�^�"�9�wn�푓��$�����$	��l�9�S5g*�9�2dO���\3˻�)@�ODA�|xg]Kku��k��$� �N��} _�����z���T@W�4EvI�#�f��=8����4l�Ѹ4�=���&ouBQ,#Z t���f�e����kXfN�.��{���<�^_�/Z�X�4!�ե�譼v�a|wK�YKa����������nx�ǵ�,��ke�#��UoE��LC[�E!+va��U�����d;1����cL�^�=w:ֵ7/d�. mנk�F�(#2�Tnl!�9+�ы�q帣I��6fl��i\��%�� �e��e�65��{#�����uHFj���f�Uu���6�صv�X���5�LE��,���, Ҫ����r��;���r��g)�9r]�����3 �I��� �H�� ��1y]L���C����I>�z �Foz�����@�\Kǈ�r��%�kn�"��d��vǠ�b�v+��6���_�x�p�)3�9wtR/;n��e�^&efz<�{��;<F�l7�x��6I�w,�$�L����f�$m|eޢ�/�{��-]���t�x'+�~~�gP�T�û�1��5�͹� ��_z�N�L�TA �l��I���A71���lS����]�p��4��y/+��/U7$����B�g�[tboz~}���-��X�'�m�x�%ec�$�q�zD�TZp#�f[:= ��u�훥��p���%�L��̉>�x"+\-s���NCbU�q��W#CL\к��r�x/ptl������o�� ��n�дc��]K�1�a]-b�P���֙N���#����,}�$�}� �O�W��� �����F�9Y��F{/�M���wb]���xp%e�"4.!�3GLx���!Wd	��F?GLߒ�D�,�����y5�"�C�Nۊɡ��LGcư��x��#"s�|O�7і�;X���O���G�{�x�+�� ���Q� �H5��"��ڟq�O5>��q��d|	=�QK%zİ(�v!�!{�j�V2�&���Sn�HzSƭkpOS�E�~�����c�}�û�1���1���m̉�%�Ow[�8��<��|B<ٻ2H�W]�gD�wr�Bh5l�VNs�)wY����lω� �e?��������fs31���ót]���ڙ�yQ��5��~����Lm�"�
�A-Q�sT[�<���������o@�B�h/C�}�W��ħ��R��	5t�\�f�� ���nߦA$v}0 ��{��(8fvEڄ�g�`�n"�O��y����� �ٳ�]�v��qD1污��d/��p
KPջ�����l�5ڛf���(_j�5�2	����I�l��eCHa�����NcQL�ł����ڞ4�Z�x�w�v�25ٽ/lr*��w��H�8 ��������$Vt��I#����6lttl6��늇�>��x��i&��g���du��,5hy�p��|�f(I>�Ɉ��/e��ɧ�/2e��*;G	���ؐ���HL�ݘ�GB�P>�,D�O����$���	=���b�iH��fr���[35� �ڢL��@ �L6r�H'��}<G��<�;�gE\<��uh�u	Z$l�t�U�T� �c'g���|=y�X���g�wS}�y�h�&r�jVد� �Ϸc�F�z�8fN��ώ∆ �@3�@��SB�Z$_e�{��@&��l_K��\k:<Yp�$�[���p�t�-ʛ���2��7�*�uz���A�Jg%���O�{���$L-��l_D���v�pռ�f�|{#�%���+�I/�$*��g�Hzm�q,�/B��"��� I=�}2	<�;��*Z�)Ƥ�Q%�;;3��;q{���mo�3G<�*���0��<H�9��"D�y���'p�$&KgL�
69�3���͐��>��ْI=�N�[8 ��d@���38ww.��g#fI �א圑�Fa�z�8@$3;�I#�;�I�Έ�{��ٍ��=hI�O�<���2��pC�x��%�����/~��K�2n����9�e��a�e��Bd��V��f��-�n7t�P??-%��:O)�P�/��5�5`�s�J�m"��p�-	i�#f��yԛTu�B��F"�Gd�5fX��g��yN��{[�M��;p����z���n��γE�����:�fٶ|WbM��u��v�ԄK�sSc���1�^	��P�1�v��7�ppi�Zkk�913G���@u�{A0��^-���,��6�1�E���4*M�s��5�mv����9��Eu�#N���3GeF���c5�.f.�>{�w�(jJ�;}�9��cę��$	��D@4!�9����)�~1�I��vL�kכ�ߊg%���O>\�����m�+���$I�����A�� ��x�0���>4�T�]�-�ߡ�|��z����E��w�<�uY�i�`	̌�I'5�O8ĕ�	��N��$|��lk2V8�\�9��{ss&��Z�A��5��rtm&�NI>��t̂gK�w`̙�"���؍�3]^�l���ʻסa�v�H �����4��[ӷ!�������i&<�K;��
E�Zwn3>w.��ҙb�.H!2t�g}��w.���v�o�;ĕ]�W��nq ��B�71�s2	�$����j�D�]'i�o�	�>�C�2���y����������q�s�7ܻ�eX������������
���e\�dⅸ1��{&ʺ����ht�����d��I��I~��@$�X�{"�t�h��|S9.��h>����H��
�RϷՂ�ot@ �?_D�H�s�h���N�U{|�Ytk�s�YQ����	�� x�	��wO9�c�۪ �6�bK�勆NY�ρw�x�$���&�}����	�� GtṽN"�5[���z�?_��ذ�4{uu�
�m�i����e��݄1tu�f�$�����~�ڥ.�,�'�v:^	���I͎؟�ֵ��$f��|� 6^@�F�R�;�vp�	����$Nh$�#�|Vr��I!v��"{g�$�nj?7��Gn^?P�;����v,]'i�lC�$gc�$A���m���B��zೳW.��l���Ǟ���vt����v(7*�d;���{�ٰr��i����+���p�`9u�{��.���򽿾�$�k�	$o��L�αA��vwr�G�[ާ��Q&`[O�C�qTwD�|	;ϭ�٣o�L�+��я��Igd*$.���H+�˭�=)��gS>$u��	��3fI$�>����}�{�):7%t+i(�7�+ڗx�av��N�!Mu��Ш�:t:�ZH�%˄��<-�A'��bA>�w�bú�J���KW(s�tH3���1d��"����p�-_Kd��uw���$�~���$N��G��߬�w�qΤ�ި�\ɓ�vNaT2�:d�/�<O�+�î3fW-/�呝� �@'y� ���S_�%ِr��U�3�pe�)��j�� �{��<O���^�8��Z{B۪�f��Oj���O_��*y����/����o~�`j�&eV�>�n���с��_�׸s��8[��.��'�'nL��G�<>@�������I�gw)4�+�@"�g�c�S����/u's<tD���$����(�s�r��v�\!�s7����V_�b�V6&�)䈖ك,X�5P��V튵nv�E��b�����	��YAwyEmL�I�}� �2�PVB�w�X܍��oY�}Y2I&��"vE��\�H2c:�1�Q��Nǧ^�nb4��D��:+�A<�ڠǏkR�3��3|z��,��;$R$2}�̪�����n�m��v��W[�$��؀A#Y�T�6��'�8.�z��6�R�m��,��d��	�Y���}�ݒ����nG���=���[b!9f,�'h7SƱ�n��G=��v{�K�Lzi�}�j.��}m���.G/,��#��/n]|�?���ٶ���P�����`>E�ef�6]��z	po,���q�/m�n/!�&|b�y�&��W7^��g\7 9YS̬[���x]ߗ���Ι
�]�6�eW��� J�����9���;`~�<Ҷ��������N"�OɅ�~;����޲������7ʼ�O�ǽ鯠r���y(��C^�ƒF{��\!�+��=��FI��Ҝe�>Ꟗ���f{/K���y��|,� �|�=��n�/{���I�` �ڄ��Zu��|:�5�?��+=�.h��1F�����#vN�`m���g>�~�fyw�#�e�%��%�q�וo�h�	�d����5uѵ��l��3�h@f{��Ǡ�vB���`��j7|�v/�]�J"y�_�>e�^K���.�~���g�\6)�
�m{�����s��\�0l��	zP䫛x���q�0[����O�e��]��(���G�Zq��Y���&��9�Z��Sxc"v���+�j�"ôp����'�g�7�/}�:�;��N�tYC�/]l�5��������滱*������w���눠 �C�4����"ww9��=����Hgz�#�ɝ���2b�P�Z��ܾ�S��]�3_�n�E|�Z��K�=�Wa�^�ǰO{5���w;s[�ZB�<s��;Ľȍ����3zs!����e��U��X��rg�y���񜃛D�C�=�� ���،U���w��lz���	�0���]���+毠��ſ���tzw�{B��|�� Iʦ�)4�`�	 ��ޢ,Gu��I� yX	�����Db�,�q̨��
UE�,�q1
�J��
(�耯D`�0�����> 8R�� (1Nc-rּeb80��*�R��PD��q�Ö
X
��ʘ����f�6����*�'0V "����:�b�3J.�&:0�z$���H	"�q ��!j�j��r�ıQAX�$H�䀝1)��Q@	� �1��*tb�8�=crD�`�A�Lj��!Z��P�T�(�m�  �$A�V Z���J.Z��e���*"ָԂ*r ���*؉b��1mh6��Z����e��X����-�V2���IZ뎠��������1��;z '�z;cg����@ܧ���3�j���ןV��8����b���=���U�vFɳ���D��c��	@3�^}j�:k�qD0䣜D�3�!��W&_mN�::xbn�RW!�3���8�N1!eYn���mym,V�X[	]Xju���J��K�`�wnvEx���oa:�=��+�<tZ�z�aB��	�k�������78��ml�\������w�X������S����m
���䔂Ĺ��>J҈uG;.9�:w>�z�lO������[��<۫i']�:[t&JpogM���js$��D���ٕ��p7\�2�GM��v��rR2��`%���.wWk.i�ڶ�t�-굌�9gS�����vS&�3�d1�&4��ȴB`3͋/dE��on؞,U�t:��jJNTn.Nܘn62=1�H�� Cqt\E�E�v��	���*��^e���1r�v�r 8rmX��0�Y�=��a�z�_2��N����ѧl�rf$̭p9�@�:ɇbW�E��d7���l��������-�^y�᧥�m]Vs&�y���ˣ6�f	�x��c� ��s��� W��\7t������lc���l��Zz�J��O�bl�kA��p�y�".u�Tnqմ�K���n9��.���-4�3^c��nhٱ��*�H�&
X)�67�M��l���s%q��=77U����1ƧBvڋ�/�o���7R�˯�W�<�͋c[Y@l�������H챨�l,^`�7gm�Q�5�4F<7e�<wi煵����R�ۛG���&��7������c���űWa�-�E���sd7m�r�cq+kf�k�٭�D�qz��QT^��[������PйKel�e4`����w,�lJm�1֯
��܀F��pE�OXƮ��{"�\i����=Gn {%�cN�ܱ���:��!�G��������7!i�t�M���x�R�n^i�T�f[�h�/a0z�e�����gh�K���- ȍD�Cm����#{d.�ñ�t'Wf�]LL���X�ο���������g��s�%�x|rv�lOi"|�y䝣ե���k�֑3��������Rmr<�^K����9�1 j4e/&�A�tķD�QvY�Wk��ٶd��"�7;�J�'Lܙv���#tٽn#��9��x�������(eX��KoϿg�Uv��ao�P�w����}�������� I��U�����i��qy.v�PO��I�D�!�2J�T��gă�z����9����
�O��%��C�h-��z�/.�*�$iI%˂�&2��,���'�|��'�
�ڎ��'��v�Q�Ion�ɓ�y)��)�gd�B�v��1t�K��`	*d1$6�2D�vś��+0A>hi� dΛfd�3��8����I�Ȉ���OS����Tx�D�fȐF��CH꺦�������������[#��T�I��{,OIՈ0�m�����&eq��{��S�8��	�q�S3�A�A �o>� Ov�n�x����J<AQ�3�o��E;��݋&�����c��}���m����h=P�k���E<���l�v��gx�IWB�2l����i�U�'}i^��2��ؚ"����צ��b�M��ҥy�WXd�o����.C	�7��L��G7�'��pv5Δ/i�Ԉp���bT
�i�$�n�I�{��sx�6�bA"�/fA ��lz���$d��,��O�͖&�mL)kOlƃC<��� �M65�ѽ�Jg����}H��I0^e�qj$��Z5����O5�ǖ�K0�ڛۙ2	[wG�F���a�hCpd�K�LC��q��kہ)-Ӏ �ǉ;i���n㎹�J����'�={>�]��5M>�����I'Z��B�CZߌ��={�>&j*��=3�3 ���6�A��ca�E���#���qܫ��i�9��ƶdLi>$9�b	�׶� ݓ�MgQ��}qW�$�7�P`���Θ2i�5��>5��@>���i�n��*!h�~�a�^	��W��b�Epw�.�qz1꼅��z���lN= O����h��!���^PǨI�R
"Iw'����H$�?� ��o�p�9���wt��Ī���97г"&I%��< �ON��$�6;fy�N�3ދb�bz�=�%��.dƂ}j6G\^ĝ�=}�6��p��KmTA$��ُ��>1�;������ߐ�n�mMc�F�!���[`\:���%e�RlNGv%f�&�n�M���_>[>R5�UV~}b.7� ��Y�Nl_L���i�ɺ5dUVɻ�|Mξ��ٚ�̓;&g�qϛ3 �q�ݒy�Sȫ�A$�ǳ�O�9gL�a慻�(�J<��f�>v_��f,9	�d�h��&�/�A$M���n朅[[D�}0=��2	��C��.���H-�s�ꭉ�ָD�Gtv̒O��s�jl�u�/8��\_'V�i.1��)w�w堓�k��~�����'��3�I(Q�k|۩�U!wz��"H���?xx|�1�@懣��G҈vt���(�-��I>9q�ʡ��I���A9Q�"|H7���07�v:\l���H�����n`��J�Bv����g�yc���Kء3�=���|�
d��h�����$�|��?vTL�[�2��M���^�7�A>˾J�$b�ȤD
�vz�<rpT�A��va�( I���H$�t��m�4(�����K(�#�r�2fvL��½T3'jd|s�\@*�^te�5p����� 㯛�>$�ޘf�},l;&I3���U��xi�m妜���$���$�����I;8�k��9ӄ�wޙ&�x�����&i��2< �n.��r��b������ zq��>�ѵ��ëj��ƚ/b\H���ϸvw~��}q��y4]�������5Pcl0�'Ke;�pm�Uj&��n�/3w�W��`��,燼C
m($Ò[Z�A��2<���h����W�4��<WR�kMś�҂�[�֏[�2h�Ëv�U�[�j;vy�$hF��Ks�uy�3�z8�6sfv�i2<O;�Pz��ZO1,[u����c�F��U�
K�Z��s�X^i	e���^B`%�T�Ͷ�m��M��Yx�&Zdceƍ÷�v�������S".��wƐCg%L�㞶�Xq�i�f��4�c�����1zɻ�����{��=��Y�LK~~SL��I �e<:q�ǈ���rÅH�"A>=�Oj=a��"�Jd�gţ�	�Z5�f�i�Ȋ�> �uDg� ��~1�J٫fm5e�ut�y|�`(�ŝ�H����@$�k��*�6CWf��_��m@�|	8�c��foS&ft�������6^kc���ꚽTTǟн�Ac���	�x��jޘ��=��o^�T��{��Ɯ�b�9	�g��CD|I���|��L:�O�'�~���{0	'���_"fa[T�D���N��>p��א�9�����D,��n�q�#N�{7}�~���A��NS7{Y�� �G7G��><���n��4�'0O2B�>����8&���dS�!DwL� ��\�}���Y�;��Jm}|�%=k���0]�uϻ~�$|��^��R�R�d�w�m��cp��ܯ��?Gd�K��՞��W^���K0��h�,T�{��i��_�J-�0H$|��H�<:���y�Gc��^E��b�mn�A><��	��/����q\\ѯ]`F�KX�c�}ޙ$�VԊD��bY!��E5Ç���$�͍|�j.:dHc��g{��Pz�z��K6�$-��L�2t�ɉ�T3:�d��=;�T� E�Āf��� ��]�>'ĝ�،����n_A&�����^�8�b:���iὮ�������yyE���y��gv_��o��ft�q̆�D=gD�H;ӯ"��JY�[�jzE��/[� ��,K;D��L�$�\<{p�[M�xܹ������ɒI=ӱ ��q���D����E��x����S���f%�TGt�<� �TG��{�z,��I1��n{i���EEǟ2�\Ɍ����x��ۛ4:m����x_��-H;��R�6U�q�7_�-w�.����������W�d�m��>$�u�o����CbōQgֺ�ASҞ��������1 M����>:��f��Cck��M4F`����� �����]ӢY2~��$�k��g:�l\wChѹ�� ��D��D�s��x�+Ƨ�2ێ��On�m����i �YWh�H�l%��,��&�:;��i�Ɋr�ɉ��^�̂A'nr=H�΁ �΢��D�ΘK��-�$��ο�ą����k�333��^=q��E�v}QQ�I>7��$��'dW��a�91b��w��Lr_' c�k ݾ'/k1���Kz�D�Rc�t5o���� �>s�$��0�#C��z�|{:`��c�nQA���D�J���=Ǯ�Hܵ�o�-�� �N>��F�a_O�a���F�ES��.V����nZ�d0��4�m~�(\����2x�݉��-�i]d#�2zxd^�� 1��9�D�B@"�a��y����DW>�*b�0v,CH-�q�|~{܉ �3�*�=qS�i�1�$���yի��7����2�y;E����8w3\%<,�W;)����!�9$.�s;];�9tK� p|������D	�=oL�>�7jU�Ȕ���'�?D@"���w� �;T/�0d˸E��T;^fD�.��j�P���^��Hn}0H8���L���<��M��C�2fd��4O�\4@@�zހ�d����v�\/�}2��cē�[� �};,IgD8gA3H���Fn⧜���H2��O���2	#�k*��+�f���قES��JE���D�ʈޙ$k����f�$ukɂI��ٓ^G�s��熾��N��w���1�檖g,2w.�{|�wsBԲON
ׇ7@A��wў�<Ƅ�}5�;���x[GOzL+ �В"����f�(�1.	 ��l�q0��qk�-��G�SP9���cV;m������L%�=����]�;L[Iѵ�U�z�Xl=k�_-ܧ;t�7(	�=���m�5gA	�95�L�/f�X$�&�Nȁg��8��ֹ��g�np�ݲ�m��;��h]��0y��[Xf���XF�[�͂2�B�j[b�-�6{�;%�<�\{^nun�v�ڱ�y�IdNZ�0�+�b��"9̿=���֔� Š}�-�L��@�A=�Q�PF[Y"WMT �{�}Yv�ػ"��.��8a�`A;��XV]43\�K�5�NC�L�A �uG��c�gg�L�3߰T�)�gN��,�Ϸ:fd�A윈$7v�b�lIg�`���$��Y���~I���b�>���%E>8~�X0�F�I �r�by"}�����NEE0&Zw�A>#�Q%�"���}���Q��ⱪ�b硔H����I>=ё �F�d;��A�#Q�f��$��dX���p��"f�-���S�r��b�65��bb����Jv(�,R-����$?��5���:9�\�3F�lӏ�]�s>$v�^u���f`Γ0b�e?6� ��Z�27y���O��f�l�l��h�e�4�HGAl��T���C�SB����ɘ`�B�o��@��a�SJ�;�� �_\W�$����@������d�`�4��H�m�ۤ��.�/�_c�A��S\x"���Q�;�:�$���ts�W�gH��Yӧp�49�fvw����]t�m"�!�M۾;ϝf��c���;F�&�j< ��D��~)��:��@�<��&fN1$���t�$7_:d�s��L(���}8�5p$r�Cjqtn�w#��H��Ϟ9�ܵ�m�t��l]����{aMƛ0w�����'ƶ[`yI�|蒶c7/YiM�x<θ�/%��'whB��Rr�E�Ui�� �sq$��O�5�,��Io+َ0	���J�
T^��j���C�~�s���Ӌ$S30w	�"� ���D��\���E���ٙ��zyz{{uw��~ߑ��5��Y��o��뎧�eq�F�>��A��ظ����WNo[>Vj���i�z��7��X�8�@�`QJl�Ky�b1@���܉�j�W}��^�=�D���V�x�E>�}��.3�s�H��PԴb��|���|���\=}����6W�o3����K-o����s�w&�u+ 7P�ni�d�X ����$Q��BwpB��8�$5F���:���'�W��,r�+�(?���VҮ\��D�㾝R����넢�O?k��>���&���Kϯ�����@K�,�`�G�"w��]��#_-�� N�1n���!o>��zS�,�����eZ�����<�؋;=
��1��Jo�Ex�z��u�K��VI��G�����+܋�}.�{:��o���o��n�H�6{<:x��Q��{Ϭs��;�/Oy`¦\q��4��)�o���5�\����@%!ӎ]᫽�y8��0R�0�3��R]��p������º��{;S�{�����X�3��)���`�|dڋ&��"j�k�;OP㟯��㳖8�bm�)��=㮟T�?(��p�0k�����(�.-�{��&v����p����a���4��{�x/���,X�|��Е{��[�mY��Λ�ޘ�|�,&|=��Ӈ���Pn/�z�{#���pٜj���|l>�oX�C�kδ������3Y���6U��������H�Л�_{O-�l%�)��SbV
�i��&���}e���8��@o4=o��<�ĚM�CA�Ő�/DIB� ����TkDH�����mk"ZS�Fc%BՋ-Q"0�8�Q�
Z�^ ! b��@�"�9"��*\�\�F��
*�Z��TF�(��(�V(J%"1X9�`�b#Z[�0b(�8��*�dW	UT��4j�#��3)X��Qq�*����UD`���@�9�*#��Zё���+� �m�c�X"� �Ä����� D B:1DX��!'�jÁ�`E`�	�J�J�KTcG-�U`�U�#���(�bUA��(�j(�eb��F�*(�TD��JH���� qX��U�B!�g =�Â��H��D@�%XD� ,�x��w�Ve51-*e�FzF ���?������w>}2	�*�'v	�N	L��Gg7E7i��t�l�	&m�'��z㧵�d��Ix�-��'�װ#���1���;;�X(�k��c�U�;YqM˄��I>��2I ���6��g3��τ�4�.S0G�m�Ջ8�]3�8�X�+�&*scl�Tغ6�'4i,�♈vw��cǉNE�H$�[�E���虁 �H���*Gl�X�%ܹ4��+�"�=�]MϤ���Q� V�8ÎE�!�Ko
��^$V@8�'�E�)�Y3� �Aˎ����w,����\h�N���>&rwfI��GDO8�d��LQi�Vt�6�v�s��)�6xX�n�I �Fǣo����/��ť�LZ�@�h�r	��S���}�g�`���6��՜�w�Ǵ��}�L���h�u�.�"�T��}wy�}c� =��y�2~�t��:	8%�~��O�֮�5\)�%��q�$�;c"<v۩G���8���{!�I�l&XC���R���u���6���ԡ���s�������Y�F�L�����:f|I���$�}��J��nj6+7��� �H5�� ��K5���v�t�l5R����:�=wSO����s� ���P
�N*��4�g��$r/�΋;2r��:�kT1#����u92�sp�:7@=k��� ���(��W<t0�q�b1�h'�/rL.咤�WE���VQ�g�$�MDOH�L��NBc�=� �ܬ��ӻ�u���6brVӈ�#y�@;[]}����G��4��yԱ�Tp���!�r�4	�����0��k�3*Ǟ!����l�q)s�px��^�R���'|��r�e�# ���JH��G�0�Y�5�!,�i�,�cT��,�n4��� $78�	�L���ݗ�:���Ns����eI�Q�q�ս8�N.#)�ړXv5l�<\�=�6p�W�֣�U��b�ņn��i9N���%�-o.���x{v�
�>Q�㪉�݃c���*�6�KZ��6�V!5G�[c��R�F�h��vr�,�]�]9���z�)�^S����\R�9i]�R"8&U�i4�tb_�?������]w���Ϛ@9j��r��gƚL�'���{[!A;/�,)��3�,J��؏ ��u��v�z	$�ƸP	$umt� �OQ|�9B %�6ӻк� �_�N�b�>=	�<�|f��$Ij���peT��@$�ָP	9[]	�Ӳ����̜��"O>B�ݍ)Te�&Ɖ]D@b	r뢼h��p�fr�)���W�_�O�;�!N�$C��)�ϓ�$�H����M(gcoqe1q�fs�r��&@$�X희�4ë�1 ,nt]��`�����d����Ofn;&�!@uf�[k��bi�&��߿B&gvA7��l@`|sr�$|Oud@񈴏P����F��9䈭����չL��E8b���/��{r���k�`��-&�J�.ٍ-�ʇ��03ֽ����Hg�~���
e	����(7�͘�@��9�B�T&�ߞ�wR�_	};�$��u����x�eI̾�O�OG���Ι�%L�lL��E�/�;a�Fk�<Z�ud��\^d�;�K�A�(35�pY�3L�Ҟ�9J���1�>$���n`�=/��2	�g��х�W�6	���H������gb΁v����G��|kDh�Z����^x�s=dω$�vDH�n�*9��{W�+v7�������(�$���&+Z&��}�cg���]�����ibF�pX�m=z���^}�C��oy�;fI��w@�	����7���c�+/����$�Q��'b�&S3;��Zd�]ĳV�;<2{+6����>�Q��+���*!yd�=TsKZ�����Ckm�'t�N��|]�	 ��p���/��t��K�Gtn��Z���˽�����(��P�+������qK>���x�B�D7�x�ӽ����]��7�.�I�Fu�\�O���P	����ӧg%�S#�bdȳN)�n� �n@�H=��G� �����F��sC�[��
���
t��'L�ÒA���h�r�f�H���$%n�A.w�M�`9˗eG'$X�I$A.�����N!�֎&;xݺ�z�egl�O9�8���c�|�}��X�v.�'n�x�̼xl�����:[[^�H�ץ��< }�z@ܐq�tS)��� �ݰCkb�dQy��O��� ��$ݵ�53�g]�΍�,�:)�%�J�҄x��dO�$�9������򁛧� X��A>��Ք��pX_� |�Jy��s�KyT��I�;Q�2H#f�ǚ��U.�����Zw�75U��ࡕIY����6���&m����w��y���]0��W��$%Z��)4�jd�0�k{*�-������<zz<�nwIӒȨ�܉�� ����5j�j�\�լ	�q� u� �A뮈���U��C�'�9���r�=\���Ӭ#�Q�ۓ�u'�sŜvR�0^r��u���pS&f���ӭ ��݉�'Z� �7L��Up��h ��ӱ ��'e2ػ���ܱ��.�͊�]er��1�$�ݜ� ��] G�T4�c�N9��PHʐm1!P:)�ϛbzD�|k'�A]�+c8���u$�/#�dIێ�>π�i�N��D��]�6�~�b� �N�H$Gll@�z5VJ�����n	��H�ne۲g.�������mP�J�o8���o�*n$O��ˈ'o��01�j�s�S- �2ɓ�^��7l���iɆ{k`a�5��׊��\2�wl|���,�{�i�8��ks�Z%B	��|��k�NL�Aww�D<B�Z�&��[u)^���	I1x��MaG�K�ƙf�2\Ɣ�9���v��=�eud�l;!��]0�)��p6ݔy�x�s�+]���#Ů�=U�lKL1����i�d��s���.�]�-���e�w�W���kv�禆�6�y��'k%�����ۚx����{vc]�lG)l� �]G[���d"Mv�6י*�B�)s(h܅�:|c(ɳ�n^mX(�f�֕σ���R�����%��'NK"���fdO��0K2�;��`��|qp�L5��ʙ ���|���6]�Ν�L���ǥ��ȃZ&�كS�Uj"�,I�0 ���F�@������|z8��8N���A�{��k9�Tk�l��\A�������y.̈��y0	��xߘ��P*���N;G7(у��Ċ�i�A�y0����'eZ�i=�n;H���#zpM0d�]�%�AY�&=p�y�v�������&�2+� ����#lBur�i��6Y��ywr�X1vN�.�+�+Q��e����e�°��{���\y'������فp��$p|��$eܼ	'�S�3�>�� 6�`��$��H����%�S#��fA �>wӜۏ%��rC���^����i����ʡ9�V�R�;�N������C�lȫ�x/{��f^�,����o�<=���;Gn�τA9{ �K������U��ws��EK�o:`�fQ�9/o �|f��$�O�5A�{^��{@�� �}յ�>'��d;2wA;H�ϑ��ל�DV�%�-���n���$k�6kq=\��\2��m�w{	����^d�="AӰ"��q|��}Pn<È�$��d�$��ǖܬ���>��������c�0h�n�+ѻv�Eђ,��E�O:�.�t��t��g��~�	��� m�W\�I�k"@$�Ot�G�xh������m�� �G\���I�K$8~|�㞉��^����=��$�w�#�	�qWk^}������΋�%�G� s�Lω$�ȂH SJ����";j"m<�tX�^pC�cN_����N*)�&�[-�>yg�����/m	�_x��F�L^g����(��S0� *�:$�|w�`Ef��.�N��,̢OMÚ2"]�pL�$���6D�H&�: ���_NV;E`��T�!if�;���Im�x$X���i9���^�{��I�� F���8]ľͪ^�jy� ��NĖA�fgt�<0�ч<��������e��tY�M`���_����{���]�#�H��ׇ�D���l憬��������g��K1gN�Zg�ds��1�;#[�>e��E	͜x'�{�s�$�#U��϶���b�˲�t�j��|� ��������<���Kl��-���A>�u��~���gd"K-r]9d���x��V.^ �Ac���9;/�>=��#���y��^CsGS>��رh#��
�~�����ݻ}�.�a�v }oo��X/�-�}Il�4�� Թ!܂&����T������"��S�o'.�fS ����@�����Q��t���SkP$)��$��H;����~µ��*����g�ܴ�{t�v�-�9�F�A�eZո��ᮣ��;���`�8vd�v�[�u߼H9��	�9�2k$n%j
wZ�M�=P v�c��A��`K���1"A�g��yGz]F�|�	�=��A><�<��Z�Xn�cǳ�	&S1wL��ZAi��A���ȒA �t�G7�ڊ�� �1������A9���˲bC���*������N��H�\��oa��$z��7�7��wZ�Uӗ�`�&����PD�M��r�Jgٛ3�H"�*"��!��nQWvz1����w��E}w��l��::^Y�w}��w�������핷mF�	��6�=�i|<�;���yyl��=�������C���h�W���?t���W�y������d�WB"�ù����D�z>�sJ�x)G��2{y��<�ӑc!Na������/�.�^����؆��ޞh���3�c������a-�PlO�4�t��d��]�Gt\"�zH�G7��k�xc��5��<o�G&�&��St���o�fq>���Mö���v��6t�$�G��+|�;_=�@7����\l�ϩ^�#ܻ����y�~z�6!����<�6c�^=@ll��wm:��<���y��`%�4�B�����!F^^znpT�x�<�kF�Rj{��l+�2��I��y{���B����_�u>�Â]�n����s��Y�=W��g�l{�g�@��N��L������y�P�{ˑ(g��}���wެ������XM��"���ݰ`���qSީ_o� �g�Nhe�Xi���]��m����N�AMζ@�����Y�v����{�rc6y�I�{gzo�Ow�g{(�,�9*����ғ�u}�I��w�@���',�:f�_g���vV��G's�y��Ǥ���wx����𽚙:cro-�S/�[�wg#�daV�2(����3�ξ�Z;��k<�Kz=��Q�����{r�{��:��B���O��ǵ�d
�㨯=�އϷ�wީny�M�azn/H�r"�w}wʈk��ŵe�- ��B�KaF���؆NH��X�� �I*qm
s`��-(��q�K�%�������X����A`�EJ ��ί<�'JЖN��6�b��L���j�QbKG�J��Ps�6���ֵ�h��T(*�ZZQQD���J�
!EA�L�K���R��+� �x ke�0�H��a�)iB�m�3�[kF(G��¡ $�i@�����dR!��+Ig9B� ���[��R0UcZ�mD*XմX1���p�9d�D��:'"1XJRRBD��^�9D�("Q*R�R҈�/s�*�) "H�PX�(�U[s3���K$��1��F�JԩZ��+� B��D� �Eg)��
;k���"1X����D�"'Y?}BG���M��f�2sU\���\)C�ɪ�3�I4ٹs�nI��γn�͛k���n9�g�yx=�@�	v��zw��[�:����{9�7h����B���nq �)�isF+Y^��rk��"U��	K�k��u����x^��%B%�)[��YD֏i�Ve�M	l;EW0�������l��7hp˺{8�+�3��"<�ix���Ӆ�6�g5�s][s����lo6�e��P]n5�(���g�2�X�)HDId�b>K�hх��nU�`M��O�j����q��:fj���r�s�)�c���Zy�U����G��ԛ-�'�EUM�5�i{Z�˨z8O&f����p�-������#ܚ,�AlӰ�.�&���l��!���4^��!fC^�c��^v�}�.u�Yqh�{o<<�����v4�f!#�Tם��p�T�q��0��Y����`�gv
37+��u�޽��1��P\ˁ���Hk*����aI����MT+)uՌa,o2���uՁ+�m0��q�&�E�[c\��J�7D��2A�Kj�V�L�mp�8�M���:���i�fwYPlm0V�e��3`B��&A8kT��&�;yw�W1��ۥ�E��.�/O��ͳ��<(�z�J/=iaJ�fj�l����]5l%��3�nT�6"�WU�.�]��Û��n8p�VC=���[Y�6)D�.:2�X���f�j���7S�j�A��eu�;g��=ת!4%�+�f۬�)p\Ӷ^n)h�)����W��n KXv�mU�ؽVV�X�*FŅ�UÚ�q�]s�S�<Τzr�[-�Ϸ;���	e���q��cR:�[3h��d�l����mN+^��f�FƷgM<Z�eܺ�\�j���pbg���y�$S�uex'<b;���k�^�3ۭ�w\���T��2:�m�%캷��&�nGΫ�u������"L�XR��B��B=��I�qʀm�n�[����l/�.�`���[q�Fzܻ�t��q�\�Yѝ�Ä:��z��3�3�H��LX�`d��)��LL�1�*^s�i���1�ӹ8�tah�5Y���eA�c���u�&��x�k�&)%���M���
'Z�$�%WY�5���Y��.|�:�wOnyC%�'�"�Ih;K��&�V>u�F �.�VE�\ݵ�����C</V��j���^Й�Y��V]'t����9vDw$�e�����{��$�/��(�:��XuSk����$��tI�~�D�p����J縂	{�nqZl�TݡA<��2H'��� �7�u	�Eq�O���ޠ�x��xM12H/��Cy �u��U6��Ck�>&�w�@$�{��$Z`��`KL���V�G��s&xH�����0$���I/r��7fV��t��L�]ȑ�fm˖dC���#v.�!��h�oK��Cm���T��	"�e�����@���>|?>�l�I�F�R�SR�1�ܩtk-�emtT��4M����8b;4M�,���$�᯽S�=�1 ��o�<gej=���q�|H$ޘ�[���NBwrJfS'�� "��vԺ���=��l.��Fns*��ꥋc�	��cE�Vၳa�Pݛj��e��&��k�Nd�vN�1���K�:��c$����Au��D쇝�"�y><�f1`,��fN�'j�~Vv&b	&�[�#�NM����A��,Gn�Fx�w)��$M>�pI;L��c��ꨨ�q�H�{��$�w}0I>Λ�V�Ay�Mjl����9�0�i���A�-��Cqz�r$�W<$@h9h�L_D H=��D�Ή�1IM�l�7S:D%�ؿ���R'�\��Sr	a&�{:�7�0�!�լ�7Q�~~|3]��tX9"�ܘ�H9��`sf�$��^G؇��@��@�A������@d�`�Jdsf��$�3���f�}�+e�ǉ�=�}2w��b�n��ˇ���9~t�g,S2���ƈ�H�{A ��D0��A�;���g鶂�ٸ�Hݻ`6i(���8�����\��<������~E�Ȃu��QYV°��j%�������}��$�j^�>��r���)æN�&h3�ᴶ�l�ГR����\x"	�����+
[�mgx�QoF"��ޠ������2H'Ƴ�={��.�-�!�_��Gl�ȟw:b6�iu��u竧���[�ئ`�')��s�u��:=Z�fv��ؚC��GyoϞ��>7F,`Kw����I˝ȒI'ݝ0/}7Ҏa�����x"	��2	�T�1!�`䉓9�����s��k3����L�v��A ��VyiZ3��}�;�nxϘ��فd�H�Ι�Ay1Ĉ���VN4��H}ō�d���L�I��ُE���� �d��	8�e�ozOB��]��ˏO�gK�$��~�/{w�5f	�G`��t.2Zf��d�e-{:#���_�׏��+���'Z����nC��o��Jl��ŧ�Rc59ǶǉO�ށ{�%�2�A�~K�N�՚
O��v�濙7�ړ3D�ؾ� �����z�ǁ�~�)�f�=��ܨ8uvL�T��hݘ�	U������t\;�X�Sg �b�U�Ho`E���y�c&I �V����:�.9��Dk抪��$>��+��۟`4�?� ���d7G�������@Ǟ�� ��Uy'č�~0Iu&���e���t�]b��2 �E��&A��>�Av;Y�*�D�X���牶��I7�1B����gL��c���3"�W6l�n˽��J��I2n1�{^�yߺ��N�j~Acj�z��S��L]�fS'K]G�	��{���TWZ��M�m�����h|��׾�>�N�=���uB�!Mu6���y��=,q��\d�y�'ǯ<�6nkr|�,$u5���|�O��Yg���x�P�)>��f��yA�08Nm-XSږ�B��WK#j�+F��Z��S�q��lܚ��E�9�Wg�.�֥�͋v8�n:BBwbӺ�\q��[׮tIt�v]��f�՘�֌��A���h�W[b�l�:��:^���Q��xm{C�H[u�6vE�s�ñ� ݽb���vA��vo*렣+4ʏ�h�4�,t�R�q�Vmat���W�9�hсr�]y�v����f�N�jػ�ۀM��]MՕ�Vfi�KVB�y�N��:L��k� �;�N�oFD	�]��i��/� e\k@'��ޟ'	�A�ϵ�:d�%�p�֌�g�I��O�#y�A$��qe��������'�"X�%���}ȐA:WZ�0e�����ўAQ��y{�2d���i����$@�=s
s��@_�.b��I�~�	z5i-9s�����q�1MȻ',ȨA5�ϧƺ1��6m:�ٵ|�p��v@'��}3�|Hz6=��!�����^�����G(����\%�@�f��e&�Q�.��B49%�bڮ�狺1vI�s{�ÑQ� �5�}H'Ǻ1�^�מ���#��;O�5��np�
p��ˤ�"An�� y�gI�C��&���G'CG��O]՞/��lnψ �}��l�yH��E�[Y�#@�tu@H�F5�,Rx4�4nO�9�q��A ���������z��kl�d�I!;�%i�鎙>덁��ٟ%��Nk1��;zd�|w�_�FT1p�E�-Q~ժ�+�,5�Ă}~Kā�=C�F5o�P�ϴy��Ļ�L�=v)5�AّrD�;Q��O�k6�#�v"|�S� �ddč\���㓱�]����k]L,����e�i1a����]��[�W`��A��mz~~}>u[�]n����G���G�������m�^�3���[2G��^t�o�Ւ]��;2cZ�ɏ97�n�ҽR�����$�O�ތ��˟ϴ���h�ڱ"�l�sf0S�gN]'isۿ�x���н�ǹ�����7oI�n+#�LC���'�6�6n�*ϯ*�Zed;�eڣ��v�o�+j��h�4�{{:q�_\0�xL EͻȆ�EU�|H9�/�2x�c޽�CQ&pĠ��C�cV���5�����7�R���#y李�2�.��.�>+�`A�IVΒE&�
�X�l9$�^�H,�����O�A>�ь 1��d�|�qG]��ЋZr�-��5����n��;
�V����b5'hg�7���.�k�&��H:d�� �OsD�p����m��0�E����8��/O�Dx���1�I�3�;3��[�̂A��J�Cm���6��ygSA$�4�^���H%�;�ۼ�:U�����Lf@<Z2<�e��$�C\al�;�'b�;٫:�	9}�EF�AN3�:I�I�{9:�rÛh��# >$�qw�$����q�������o�w s��/Oc����*�)�;bp�-�,�)U���nl�t3b2�#�t�`���T^��1'.^�p�Y���b����4kvA-D����������Θn*��9�s��ĥQM ����$�v�c��-]�[h+Yq߀�`���C���ָ��.u�V�<���DtMkI��`Q����= ��-�~@������;�>$�O��b<[6��D-S�^y�V��U;�$vX4�W��'$L��t�n�y�6��kmɽ�y,+��Nd�m���n�}ź����G/p�f4���1�I�;�3��>�ͩ�;2b� �7`�h�h�la �_N��$_LA�L݉L�8L�|x����Ԡ�^����y� �ۓ#U�7(<Ѥ��,�ێc7:�7C'b�\&v.�ԃGb2��v��5��c H욹	9{1 �u_S
�z���(�y�.U?C�g��+���Q�Oۚ�-�����`΄NU�U�T����$ʳ�"}ܻ���wIʯv1� �>۹!h�`�ZYX"��`q]f��4FYt��q���s[3�+������G]=����;�#��n��D��{Z�zm�[�n��e��4���8�=6���u�VѢ��7n�xe��h���4bV.Lk��M4�̫☷a�l��.���d���HݱK����!M�#4�b-mv��	�c*�s��X;[�	68�;]�[�x����۞ݹT�v�,�[Ê�Ʊ5�_�_>q~ [�k�}����%�v"$������>�m�=9=3�|I��x�#	L���L	hD6uD |#|#�z��m���I"�& <���Qcn��=St{�ƴ�(;NH�ў�H8n��K��	aڶ(\�K9�ްO��ɏ;����L��61vL�4Ц��n�s<3Tx��@B�]�I~��P"2ո��mi4������Ħ��M3yW�]��0��OH�r}��س)����� ����-h���flg��m]���cp��m��ܐ��aC�e�]
�L�Y���K}����V��Y�|?o� �̘�'�{{2��2�'b�'��0�����33�S":#�H9ik�~�������ݾS��=�'6 j\��}x�|e�q���؉lb�u�5��&B�]㷲j���ʻݫ���Cz$S�q}�2~��x�yA�&��=?3���o@}���mgn�,|���ne �~H��O�g<���ȓ�[O'���]�w�@)l�G� ����>=r�$RN�3�"���K����I���5���ob@$������h�fv��~.v�����Y�.��:2�û|	�&!�A���6�H�m$�܉�%�A��u�C]�ub���wH�V����`��4�.ʡ]�n��t�mv�':.���n�.݊L��`p��ė������Y��]P���"��4 I/��3�E�Β]ٙ�3�D��p x̮�,�1ݓ���>$���oFԒI�ɀ ���gn2^�!�͏2���� X2���ٟ�H={1Ĝ}�,���ztxyg�.^ݝ]]]]z�4�ڤ];���ϭ��� ��ǼH��z/
!P��B��g�3��oeAf��1[���yo[����|�Vj�D$��mM�#3e{bY�t�u��2�����B���WN����	(�#���_��v���h	���k���})g~��1�i�CǗ�02^m'S6��৯��E�+}�;�hl]�uyTG�����u�۾G���O:W	Β܉��H�Kr(%۔Y�L�q�?no�ڐ� y��p�?�ͫ�]��&�������|(����+��F�6����x�ー<H˼�)C������0��r��|G^����L���s�g���=WY=E�J�1ܴV�|�����j�j���>��F�e�n������[7
��Z�G������Wr����5o	<L|�������kWB�]��%o�ݞ�F��R�k狸4fXʜ��W=P�j{��g���>�H���J��|H���|<�w�����t´`Q�0�S�NuE�ў�g�-��|¼���c���2a���h���H/�%���ǉ���|�~�s��g����{��a���%�������v�>�?ol|PҴf�i}��4�hi<{�Т�~�*x���7od�m��5}t��$ O�R���v�8�b�!�qa�F��郼���;8;��(�/q���gvo��Ӟ�o����b�ˏ��<�l�(�6��q����}�*��ֹ���t!���b+AT|A�����Uij���R�(]��F(�,Y��2�UETT��%XA^D	Ő �U
��������T�%9�
��$zĉ	 I��#�@ #�P	9c�zpH*W���8�p���qm�RWYSP�[T�"B���Q�jD��ڲQ�V�!Z�k�"Z�P*"ԡZ���iQT����T��YVc�N	+g���"++P�`��Q	T o.+fQH+�jDJ%�Q�� �i[J�X��Ub�]�`�R�����W-c�U��+SP�D��$�DQJ����������ƨ"��(��QEP`""DPD�`�(;j�e%T�䕎5F�F
�dU*T���H�*��xzK57|H]�2I� �z�&���oȤኙ�q��;3�9�	7���E�LAvy�-T���##�|��fA ]�4ԂE2d�����r���G�^@x��M[�X�{�K��Ȑ	;�1#�W4�k'��q��b�1�f�	��.L�vt9�;%b��7t����z5�7�n�]}{�{�Lu��2�w+ι�I&�f �$	Օ� �y�'I�l��5r$�]���΍J�w�g%E��!�tGU��fݽ�l�O�;�1��9g[z���_'��-��h��Pݠ]�g����(��G�ϒ(�\����M
)7M]I��q�]��	��Pb�2fg:,�@��}��-vj*�}	>'Ҷq�x�������.���w1�;��IKELU]����۾� ���<;��Np���8r5b�V1��ݺ}���x�.�_.�eU��j�d�4�ZgA�=�	7��vdy�O�I��Ly��I��ȟg�̱0'�xO�wD�}�_�<	8ݝѕ]vᦁ�`��e�/��WW�.�Cl1�d4�y�z���s�cg�T��v("��+�'Q(2ffw_/\��Op�I���	ɹT�q��M�DF�|a��43ad����h���a<�8����Y�27�	$�����$�c�I*3w�;�ӓ+r��<��w�`�@/9H��I>3��o�OK�=s�����s�A w��u�S8)غ-B��x�B�Z�s�x�����w�I2��2I'z0|[.yT>�S2�	��O�ya�����p����I5Ѱ!�1vM@#�������$���uo{�p�0�t�t��4�+�&�.-(F¡I�u�.?�}3Ћ'��`k��Xw�E�Y���Z�to�� ���'��(��f�гW�}�C�`�N-KN� �cYa��	�敢��F��j{N�5Ξ��]#�v.ֵ���6n��\�
��2�,M��M<��|4<�p#ӱ�d�7��m�kt��Ɯ�s��v�8b��.gxG��T֝�Ч��:(;p����˺\�h�֍c�k�8��9��vm��$����$��=c�n����m���i�:ڻ.�y�b��X�r�p�x��MPb!;�㖭�d^c��j���!��Bg�o F]�&CB!ٓ�d��s�(�r�H$wFD͚�e.��4ݧ�!绦A>��q���L����lSF�/|��.]��_^�z�/}�5�D���7�c}Ͱű���3�bAf��;0t�>�ȐI��q Ո������Φ�	{�ɓ>H��=v�YX.��#3�:$�����]%��N\�ğ���H=�OCDF*���q H���ц4��L���h�q^P+z�(�y졷�ԸLt�ngvd�M�l@$����a��d��Y0���mZ��Z�!���:�3� �������n��Q��gx���hffw(8L{��� �N\l /%�Oo[�3�kYm�1�3:vd���"v�̙���;2�Az"	�O��^٦5$M�M��8m<1�};K�V_��>�(I{��]L��3���!�/���ˆ�Y/֜G��%fI3J��Qp�/#z��È�Ëo�a�,�s�� $���<	�b�Y�z�p��&ڂ	�2d����pAn�]
�v�����(/���	�]m�%�bAf�:A�y��˚����ݬ��U�@�|��m �C��KG-3J��'�.� ��4�fb�:HkQ�Ѱ��nD�V	~�T��U]�A��m�~��\([�d|����.�ƺ�V.�B�1��XFYa���d5,�K�����l	-t=~{���ɦ�t�}/އ�L��9$�?ntɭl��A�(.�� G,��e�Tř�ܠ�L��t�$��v�}Z���U����D��f�v>����d�A���&,l1̃)�
;��	 �^�	��#�l�K��t�����Uf4�l����cfa�dߍ�4���z�3�H6b�MEЦ5҆����,���Ji���Y�����^rq�9��*�)V��!���|H��'�E�$���=3#������/��H�h�rO��fA ���KM�)��|0�2	��ؐY��w:����3�I�&Wr"�t[�Uz�<H%�w�A ����d�9$���&�hr�-q[�s�ے�n�t���F�;q��UAab뗇S��'��GUcj%�31I�$8Yv��y��㽓��"��B�.�h�$�^��=�y����p�8,�(g���هW�{+�#5s�A �.ٽ� �H;�/� �o7z�֖P�Ƙaw�ʂ���;��B:�f|H"�fQ�u�w��\���#n{fH 7��<A�Oe����v`�P,s����v����P�Q �F�v��������u�	�נM��O�0�ox0 @�{�nh��*;j���L���<S���gQ��'a�z�RU�Յ���a��`��N�<7�i��wZ�fg���4�,�`D�·�O�j��N˃�x�=�$��Lρ$M^� ���X5D6�<���s���fRF��=n�G��Gs�➸�m^��r]�㣶%��b���р��;�!�~᭽s O��L>$���Z=<��U�U�c�A{-h�p��á2x��AS��|�w�s-���O��>팈 �W����fB�s�}l6��d]�i5��Nsߜ�Od}�{�{���[F@�I����z�[���X' S�~�:3��F���<q�b'Vd4	�l�L�-��}��W����w��S�3���T	�N�vOlI|�l�6ᢩ��;�o �u]�G��龐m����ש�xܳ��n�1�'C��u���{��Y�AT�7�G��O;��б��ë|���*�=��^��hO+}��'������F��S:�]n&��دa	Y���˚�mܼۍՙ�Z����5ڙc�\��9.�4&�[gX͹�pGe�ff���Fn��NͻKA��]����T`���o!sGL��6�\ۭ��m��Ɂ���P�խ�H5�\�����R�Ai�����Mv�,n��V���OO�r�Q�;'R���p�Γgn6��!�j[��6Wv�[��T�-�%��զE����]ha���ͬ>t����%K-��$#�TtAi���	Λ�k��=�FM	�aH�/۱�/$9^�A� �w;�!�x�lۙ�����q]��׍xɮ	�>��AJc6�_kel<���-hrY��p�L�����%]Q�=>.��㕪8����*�	 龙�Z�2.��tK�{����:��&V�����@;�>�~ɐI>=ј_�ۄ����$y�E4*�H�L�]�0NK??E�E�����͔d�j�&㷢A ��6cv��.}B�K��n-m�s�(%����آ�7Í�`�����,2N���v�I�Z��$T�ź`9��{� �Otc�e�y�4�]��i���͑�F�Hdȳ�Rf:6 ��_mN�u�a�5=W9�T��/�n��M�N��%hz��1�����6@kxW =x�s$C������3������MS��8�0���$����$����|\mb��v]����@:��Pg2;��r$��L$��&���N]���y�A>��ِO��ɏA��'��p�L��w��ҳ�`+^��ލ�|H�y�$�:Z�n{����cc�$�a���t\3�]�Iָ�A�>2s��ˡ�3r�ln�3z@�~��5gCG�n;SZ�y}��nI2gp��� j�j0�62�J݂�.+T$�ֳ��;����p�L�]�0N��y㣤I>5��Ă�a�:A��[��qr'����FVⰋ*d:��Ux�ި�M2+c��FvE�w� ��D	���i�A}�"T���=�e��yf�RI���9e�2LlA'Ǎ�C�H>�d�R�4g8i���	dv���[������A񦭉x���hQe��Y�J�m�L��^P�/J���SYK�;�����>���x��:;�'�ē���rC ���ܘϜ6���5�7y0	#\4I}0�2�t<��60$��������0d��	��{� �����~d24_VW�	��Ù1��1^����a��~|��� r�)q4���Y�G9k�[��]g[����+V#.��@����k5�����E�:%ۇ{��؇$�����5Ӷ���%�����!+zXG��H�L�]�0d�̼tt�$֕[��ʗ���[�O�Z���A05�r����/n��^/o�@۳h�JPd�"���9�>=�A�T�C�s񼽠I4�᠟:;:d�g�w&8�1A����ꞛ�M��2�����#� �v2�D�A��@�\u9z��-�w�*N
�f�͝��S���I����}��f
`��S=��k��U*�;��S��N���c�)�;�[���.���J �rP��	U���w$2236.@�A�r45�Jk��
��|9v�A �ѻ� �I	W2`qV<�3�����0ƺ�	=��5E�v�<^��Yr��e����\��*T������0p�3�Bq�/��݁$�Gt�Ǹ�~Fc��h"b�@6��]�AظgD��.�����2��v�� �V�I$N��z����)���s�d���^S_�y��Zd�;�80*�3$�Mt�A'�0���xoZ��S����A��ؐA�v ��4�d�A�()������Ei=��A���A&�q��H�����tu�3XJ�ʙ���0��P`���ce���#ν0�e#W�=�Sd�I���8��_������'��ߤ��ꊂ��� Qk�����G��PD\}z���o;�cdp�����������"�,�� ��0���
��(!"�ʈ$0 ȉ� �Pa@!�@�l:�j0�� C(��m&�H%l$)3$ ��HRfB@)-� RV���D!�@�PB 4e��������C  0 0
��0�� C�2�� C��YQp(��+����ʋ"��*,2��*,2"�
,0��*,0��,2���+(�ʋ����0�̨��*,0
�,2
�*,2��
,2"�
,0��ʋ������ʋ��«���"���8���d@UhP *���_�����8����~������C������t|��W��~_J�
+�������*���W,
����~����Oy$������((�������:��c!�������q:�{���>
ǣ�UA �
@� �%&A�"E%$�@�B	DI 	%E��FTXIQde��VIAa�RTXBTYBTYTXTXQ` E�EO�$TX��0X����S� QiJ�(@������y�_��5�=�>x�����<�ѧ�<�7��?�0���7c�}���|�����>��z� �+梂��(z0�!� 

��{���"��O�0��l:ƁB�����	����4	 HI$???��
���	@o�oר~�C�5��<��������TWP�~�TW���j��ǲ`��p�f�=�א2��q�*
+�nS��a�����p�{N��@ ���������+����׍���C�?��d�Me�WLZ-f�A@��̟\�~�                                      v  p  � @  @  � �    � (h  @  6�   ( ��                                               Cx���f�.mو�&�Bb e` f�Y�AL�Q(�a�u����KN �i�"
b�C@@ �@q׼���!�� �U��Ms5Qng�\��΂� �P�LC:���5D@U�� ��� O{��Q@�          �J���94�ƍ4=�t�eUs�.cW ��x =
)�S�`4�^6��W-J�2��y5�Z�� ���ڔ��(UM͢ {�� �s�AWf�h�L� S;u���y���px��]�@�N� s��J �j�r�0� uBM 5��HE@        ���{��a�A\کR�P�� w�U9�\�:Z�M;��;\ :K;�l���   i��  4�5K�c���Lp 1������/0�1r�p 7v�������@�g@]b�wT)  ��           oyjF�wKjV��\Ǝv��70ӭn �:���vҍ�]����5��R�8 4.ܚ��2�hB��h[4   B�5퍚�`�` Z��q;�R����ШFA�� �v�nw'Z����.ƜMP�f�(�( �   <         yҞ�������0b���5��㠭�� ��J��L۝�T�nn�i�1sh:��ڪu�6D�L�sX   x  t�3J��+� �@���0�\�I:���ڂ���ց��T���U:�\�� 5=��J@  S�&�����  5&FF@ �ʩFjRP# #T��i2�R ` M(	=R����i&a%@Lڶ2�IS(i. ���� �$��Ng��!$ I4I����$��!$ I?Ԅ��$a! ���?Q�����s]�5��v��M�ڣ���F�v�s��bY��が� US��=�%�,�yP���F-������5���uz��i�b8�Y��A���1^ �l�r\�����Uhklܙ�t��h3DX:w5��V	�o4΀��:�z�!ͅg9�hK�v��j�YX v	�ߜQI��x��f��D#ԭ6�.6f��;.͵�ch�O�W������q��3��vױVaKf�p����#�\%������чr����v�;,�Q���l����e�ٻ��� �N5��R�s��9�B=��	���F!ib�o���͗��C�;�+�n=*rD��0.FN)NoD ��xL���id�v�0�pc{���|�=@9w =��d[���C��PpY��C�rs�5��gwR�[��<�鷝�0u��:.�A���ۑ�P�	���P��-���ܷ�i��?N��w��f*����L��H�U�7����k[AKv �����b!C��5hDoq�Vw',ღN��(�x����cYVh��ONatMd���D�<cy�T����e�.�@w��v��w۵(����$�/�L�UUp���q2��n���$����\�-Sַ�[W�7�i֮5�y&Xǽ��q���)��j\y���h�%�����֘�gn�o�6��3zn�8��n6��3��i�59���8V��yJ�
�)g<ݜ4{�-�öd�iǮ-��e=\��Q�E���]��"��ugkSi�ܱ�SOa�Jw�h���ڟiH�:)�A�g-�����u$�<�r�ܠ��б&U�D8c���t䡹�QV�ל���rC�-��\Kg���w"�ť;�]���h��!'�xb��t�kȨ,Ӓn���ɵd��nnm�&�jGVvӏ�d<�E��1L�b9 a�z����o�qv9��:�}(\���^��g@�G@�������-c�;%1C�I&��~اq���x�]���l7�5i��d;�Y�x0�[˂��i[���a|��ػ�U 
Ҏ�syPn�[��A�ݣ鳨�3����4#�xǷ�ü�H�wg	E5]��u5;ݳ���jg�7^U{�������mKۨ�܀9߮��o+yd����~�SͶ��x���i��h�}��97J�����+�*�_k�'�r�S�V���*��Ӓ���=�N7��ڷt�5���x��V	�y�����I���F����h�g>(�ٲݿ�=�����;�z����h��6W��d�.�+OWv%5���Fj3�+WZ��2quG.��V����5a��g>M24:t�t�� 1��+q���s1�<L��?�NI�Y��*P��E���ʯi�A
g�@��}�f��jD�
��W:v��jl��D�ˡb=����U@o1���:ր��˯Aq ��u�t�3w��z3�Q��v5���;����;{��uOr��c\5m�� ��M㋳�z�Nr��i��$gk ܐ�Mx�X�D�,�c�6kbv^:�E��@`{�pv2L�.�����N�{�� wLo{�.r��P��5;NS�`��vP��I�;��)w.��p�m����t%0t��֝ �� ��h�^tt�ɫ�=�9Ńp�L�'��w5o�����c(�"��j�-��<!����8�+����B�Np�+�7�`��_-���\,�-ٱ���d��h|+�]�&��X����c8 �^n�1�뽪��!K��ʮ���q�X��=���@�#jo�s�c�R�"��)��z��s��NN�f��6�y���Ur��$'6cS�n�u�\$u�0[�o[���������
*�|pp�4���{_amgi
<�Ǥh�7���nRui�wJ+7�owdi�nk<,fv�\8�2�۹�V���U�^td\�e��p�G9b�ѷ�.Ik�F���pF�`a�"1ix����Q�����k��x������q�ǍŲ7vk�p�DD�Ừ������U��/�U�xL8������(6���������mELhɪf��.���bq�bC�9QF��{/rC��p���1%9���'�heu4"h�4�)�ra�����"��4��^㮗����ݤTp�4NUh&�'�q���q����
���'-o�^#�����;�e�u������)�"i��E.���m��!�4��t����YR��8YP��y�� �1�Σpn��7��2���EB�ӹ����ߎ"��z���]b}�Q$=�e�m,1>��״kOBYu"�7s�����%��'#�m��7��;��svm��U#e��At���x��Dc9%�1>�ݱ�ۀ���[�!�ǈ'���*f�gN�
;��]"q�F��;����r귄�����Y���6���é]u2���f�^��o-�C�^ se�o�]}�N`P#�N�)����#2ŔwK9x\�<$������0w,�����9x�Kj�=Z�߬�x���Tf˼Ƽ���'��C��a� ���h�E<]s%�*��N<܌ΝnZ�@F����/{U��!�RvW���Z4PλDN��D��$�Y4ױ�5�`A�OK�(���k�;9/\|-�-���!�")�tΛ���'ei��)zux_"�t�S�mc�Ơ����2s��C�l�J�m�m��<+;�ur��+6-�Q�P�F�0�׷�gsѬe�x�l��+�I�7G��:=�����k��yx����0����S�&4�b���N�p��9�5��^A�Zk�nZT`������׺Cݲ��)��^U�	� Cfoc��m�F:�F[=�x,�/�I�J���o#�����P����2�|���MxLrq+�[ܕ���K1�z�Z�4��T&b�k�l�z�Cw;ú%*�	��No�Ӄ�M���Dл.��qYY7uT��p����e�:�؞*���q��M�,m�)4��@/��mnKj�b�ѩ�~���i�Wd�3��-�%�f��_�u^�n��I�)�)�k�7�&�h�F+FL.k��n!����7�51�!t��a'
�@���e�ۉ�bK^pc{E%a�T�!��J�}�K����;������AǛ?+-�NM���qa-/�<q�J�v(tm,NI���w���9����#q�3��z�	���]O�̹]�PղN��I=��ɰ����G�'��Y�������NLƑ孁CY���*vt�,`�z�;3p��W�@�G ��ѝ�(�G���L0��:5wy͹k�\�m���@�S
����+�d�4������a��V���~�=������0���D'���˫�'Le�\�� �TWo��:�_w�����(�.o�ٽ�M"�����^��;�n20rq��F�9��C�N�5+[���1p.''W�W�fMô�Mɫx���Q�r3Nn����&�xg<����v�@�\S#��.�e�9�D��	�N VX�Ν y��]�൝t��]���[x�;N���Wl׳g���s%.�bs�ŉ�ڷy���$�l�v��ۯ-t���C���إ�q�^�W4��5wV�����X[ߓ�B\Q3�޻�ʠ��#��쨤Z+��k��١a����]��\��J�=��x�+t4�����eƔ���"Aé�=�5����v�ݺ��n�{I{M���1#�:�:4^U%y�CI�5g7y�t���G��)q罣F,r¦+6B1�������fn-3*3*/��~�}��ډC�����%��5b/5�����6Q)�mg1�q�|�y���S�����Ávv��PY���4��6*%.�t���G7ێ���{`��r	?�p,�����x��ϊP18F+��Yw��eaВW��z���ۣr�׵/τº�N1,�4����ئ.9	�G.��$կw:L�ׁ�\�w
�V���z�����rN�f�����k90�m��^[�jf�v�0;p��A�-8�ΗŸ�|�T ��M0�r�ད��C�AZ0^����;�`���7>iЬ����fk�¸E��Y��E��{�~;�V����{����N� �(⛅&��b�N��g�Z����u���Wo>ђ�z��J��4�������_S�gL��6v6�L��w��>o��i�;-U��8��}r�Í�"�
Ʋ�ke|OAdo�hsn�Æ�l\Z3M�q��/ y�R��yC�:������fw�u"��;�ˬ��S�XS�ћ؁ћk`�פ��c�:*�Y����ͬ62���"=ܜ&n��������à��.��M}����7ck`'�f-ⴾ�f�[�;_jY�	�Cl0�DH��F'_�ـ�T"	qlt��{�з9Ar�;ɕ&��bs@����廲L���Ӷ����o�rmܼi�F@��3\�ݗ�k��8v���)����$�F��vޯ����c�������F,6eh�XZ޻׳����.�{��45&']�?0�����'=g_i��~eթ#����^K�p��7T�t�V[]���O_�,�c��Ӄb��v7a����������ɢw�t��ޘ�i�w6gcP���Ŏ�u�H�YJ� C.;�h�r�Y�3����kM=����yլM��)�rd��zPZ�7�ز��z��q��)mw,1a3rf�vi3m0(�7Yre1��&R�q��h=ٚ��`Y��F<���5�M�2�Ҭm+BW'�c˵D*u���A5��SYT���I�2v4��hٵ�8,���G���n3,jj���4c{���,��4��lœ��N�S�6۝*�:��!*6H���[2(��6ѵv��[��ԱYɍ�&KyThA�U^�t앍Q�f۳5�U*dKzb����G�ڮ9YO�W���v�}6A�]	�p�0�a�=xn����b��v1��~	2�&`��/x^,�Z�ok�P�Ԟ�Y ���0F��Y�j�����OOl�`�{;:N8�������O�e��t�nt{$t�?���t�[��hݴ�݃C��"�80�u^|�B�-R5"Ƶt�!�o�G�6S�J��͋z���5��a���ČB�蚮��i�$Gb�Wm�>�\z�&q)P�gt���[3�4Ɋ�[x�V�n�o�K��"�׍K�����N�� }�R-+�c��OM<��WrM���NU=�,��D�=۴����L6=iN@�9���+ä˚��h�y��41��m�*�p��b���]��/I��83���=u�� /7tAgbOs��s+��c����6���3�Gk�N�}Ý��O�o#;s�/���㉮��� :�ю+��vmq��(pVv�&Vn�t]#^	+�p��ǠP+�����U�$��hdn�%�ۮȺ�8T�+A�p�xޝX��&�%��@�_�!_i���.G�Z��yۂ��G���q��,`�xxps��2H��.�`�KE�ŵ�nnɽ�n���Gn�$��w[��ۃckD�v��$\2wn[a�q#�=�Z�O��*!�w0"D��D���#:�-�髻��@���;���ˇS�4��wP��k� �
��ON���N�(���ur(��` � �wp~��wh�׺ 0���ۭls9��0�Ug틔�PcF0]� ��.&a�6N�3"��P��p:���l�k�aR,[ٸ7�8�s����� M�7�VgC��E�ұ+��ǒ���٭N�N�gY^��X8�u�;�z��:o,J��U�0q0���8���@����f�y�%�N��1��<<�5�:O'N�s���}1�4�5�a�9�Kz�ͼ@�v���<�Հ�M�gm吢d�9�3:�A�#%�sl. 4d��.{n���y�Y��Gr����t���ꐳ�QǕ���ù&\��x+��Z�v�d���sKx�C	�=���_]�r{�.]9��5`�0��V�[p�r;�����������N�ˏ]�8�ڭ���	�D��ZB��]����p}�h�;�E������x�9�47�ͭ�˕?�\���
�ܤ�jb�g)�8f�=�J��?u)�w�F�r�����c�u���y�{5���y�/x��RHRH�!�<�Z�Q2jˠQ�Ms�V,��~؄�yv�����z�]M�����(�P � ��w&i�#׎�;FpW��M{�)V�ݑ~si�e�E�I���ٓ�z;{�RD.��^��8G@���m�� �F6/Gbv"x�A��U��wT{ݷ!h�R�2w:w`�$�0���U�(Qւa=�����B159-Û��-�yѨ�A�0��Zjc&x�]Oת�"dJ�~����B�;�5e ��pUGj¥��u��$m#Tٔ�8Y��4��9vZ^Vm�|��m��y1�  A�;M�p,7/%�h����L�{yp�tf�;W!�WC+��r��V޽�<W^
a�OI��;�Xf��N�۹'c3.�e�xy�{�	 �+$�
�V��Y �Y	"��$��a$*IP��d!IXHT� BE�	 ,BI��H)$�d�"���E@Y"� $$I��"�$�J�������*@d ,�) $%d XHJ��$P�RIRY	XBd�I(I	P��@ � � �a �BJ�VB
�	@�RB� � d@$I$ � �HH@YH(,�( � ��	!+ (B ��d�$��I"����@�@�P �$�B�$"�$�I�"��T��R ,��P$Y$ �d������H@$$?�B�x��������a���{�:��Bx����]�o��RfV�LN��������c�A�m��,����1���������:W�yт�|���yN^Sa���'{w����m�U��\=N�u��q�M;ǈ�0Q���_~S�w�K0�چ�G�-K�]M����8;x�� ����A�?x�5�5ڹ�bA+�;���,�YE� �Q��F�i�Qo����<b����g[ש�_Q�x�'��3��ƍݮ3�;���W�SE�>\��H�1'�6h��g�m]�z�7���c-�n�A�,�wC=�{ui���5��]��/�����^^>+9k��X�p[�z�ձ�`}���4ܸ��|2W��Oo�zz���5�`�O��8(��w#�����8��?���S\7OS��i�@�>�C��5�
F�~l�dΑټ^��C]}h�e9���޲>y�}�&5|�
w�Hh���s5��\�_e�dF�E[>� ze�]VN�f�!_��jU��^����o/�[��o���)J�u�~��k����8��Xz��)���ƇR�<�S��gw�'�)�)i��N�&<ע֨�}6�I�>�p�Ul�y���k�۝3�E}�'�}�I�b���@�A�`��9xK�pq��V�K�{5�M(g��G��~��8y>�qh���祴ޭ������j�v=�;�2���L���^ڵ�a��~��S63k���o�FP�7q��]>�||nx&�!��_:�md}ǽ�D��x�9k��V ��X�H���g/��t�_���	����\�3���%M~�~{0W�q�{���[�g9�f���W�{��ÏҏS���1� �ժ�������=���w��a$�yK�F	�J}{���y*8�.���8��x<=�&xu�Ϸ�"�Χ�{5�w���u)�_{f�Bx0��_;�W5n_
�(��uBom<�,�dH*=����5���N���w�7<�|v9N��`�wda�e���]�߶��藺��5��F��z������==�7�3Pz�;����!<�hś�%�C�{;�o�B���g��wr���&�`{�3�'�/g��_Jϟ۝�Ţ����n��K���'�=T��Z��nz��v�t���o�P���WD=<�����rι�<;O�mi[sިI��c���c(��{��1̞���=ˮ��3��g������u�,~
�?ݞ���+�a�>^GT����;���ٽ���.S^�U�"e	��ý��N�e�c�qb.����Vh9|�J��tP��f���Ӌ_�dwg����e�����od�w�P=v��fዉ����G�r�z5p���K��W�AO��{o��>��4ВV����uPA���1W'�1�]S�#����a�L��oM-v�Pb���2��#��VEh��I�j9�X�P��]�{�փn��%ˏ�ܧۏl��v1��e�<Z��[����o���?`�p�,z��;�o&T���ڞ5{�o�N����z���+d����2��7s����z��KB�'�޹e���3yzE�2;�m�;�?twݑ�g�f�q�;{����m�'z�w�垼T���|��� ȗr,���p�|�}�����P������ge6�,���0B�{q���d�����d�i�m�<23���B�����a!Y�l)o.����'�Z�(gf�5E�H�=�=�����vg%�G�(�N�f��S�C��p�n�O�=���cjf�����h�/w�J�/iZra��"}���]G/\](�g^9jgN�+��~
q���H�'���D�tSU���Dg�weK<�y���}�Q��5n����/>1d\�^��c������e��x�(�8˝��|d^���7��bz���5��o���8����.����<���(X�r@�_M<=���)���hv�:n�G~����vE�h�7�z�}-�+�o��xz{{�r�h� �}�lk	��h��)a�Õ�D�s��{�p�T~�ڲ�s:S����ٱ�xz���O�.'�X�.�ذw�k�V�O<�=��ʽ�vs�,�o�p'ǌm�qd���9N;�=��
5�A9�2��
���'A��w=}�ߏ�x�d���4=��!0MT>��Z�S'ά�`��@�{gk�y܏��V��+�[t�{7�u��TL~�)ow�{n_i[;ޕ>
B�E~Fy"%X��0;��݇u9���n]���{�`�Y�!��-+��nϚ�՗P�˿VU�<��g�B-�3��I�B��V����V_ab�*o�WV��o�p��L����������Ҭ�M��'�g0p1�&_\�U852k�����[�:��.�u�no�8F�f�+�9�m5���:���Ar��T�&�+�g����nU�Ě78������]�U���[ޙ�1{V�^<F���f��?��oBOEsV�`�X�x���|q�Ψ㞻�F]����swD>�V�i��W���ȸ�U�]��{r���WI��<���|/q]�<F�G����k'b�`���w��_���|� Uur��2�ڣ����Q�ó�ͼY�lqK.�F��b�D��pegҜ��z� ��W����;s��{���cA��d�n1����ȫ	����܇�Y���˖a:�{K��_=����o���:d�����������	�gNL���o��w�F�] �n.���[��Z���r��~򣏛�������o�/�Z1=+H�~���㞰�aQ?;������Ȅ�v�v�����ΚQ8jb��q�xy���5p��������=E��~�T�N��5�m8}v�Cx�oT�w.��@d���'yEC�F���Dq�n��L���C�7�"��v�Ǐ
/_F]Y�M'��-�U��V3���=��wu{��@,�]wӻW�νCw#x�>K���inG^P���'��s��zxOg��,R�|7���� ^��uz�w�g��=�΢{��'�l�t��\�'�,����,P�6�Fq*��D�_f�n\)׼<����Q���`��"{=��>�ۅ����vf���xa���5铣��ι�u�N�[��M�x�QS��ɷ�ȴ
����~>ל�۞^�[�����-�haG�S�0����V�hS|y���$op-���M�{Y��n/VY~R'L:����X��V�c�.�wn���_����~
Ž�/i�c�#�����#�Í ׆�݇�W�Ը���o�94����Zc�����Bn��}3{}��Z�vѝ��s�U�r�A�)K۝��L���)֞��S����6'v���� �f8��?P��DF����:Ld��U��Ί�ׯo����Ę.;��]�T�xUWv����<.i��>��A�Is��;=�=_91������v�yg)����ӂ��f��R��O���~Y�.�m9y_3}媦���=Uꋪ��f]�5�d��z���[%�v#�{h[W�v��Y��)��c�E�P�&���L��.B���e�N�8_Y�yG��=���䳻��ռX"L�:������K�{������-a(,c���g�IT�N�n�|ZfG�3�xk�����ԉT{�ۃ�8��\�ʇ������O�c�<'�������t;Ůз=�}4�{m>���=�ⶁ�yS�#��>���)��T�vnn>5�.m٨i�7p{Axuw_6������Ni������K=)/��ޖ�1{=�1�N�u��w����n�g8��n�-E�h�@hW�������LI���(��9�et�Q��x-�ӻ�˻�@��_Z�h�Wuۉ�ڈ�إ��+~ǪW���[!;t���\��0��q�z���;رlFv:0�q寱���<t��F��]x�b;�x�{����;�5uOS׽���P��<��f��ͣ1��N˩[������=��,��=F�)�b���,<{��n�U'�7������НMso����:�1�r��&���j�C}25������?^iO\Kz�횔�ֹZ���)^>�(�Y�Zwr��{�I߂��G���U�N���:�n�Wtf�$Vvܙo<��ׇvPG	�L�^�Of�9�y㪃9�=^bx�o�`�_=�f�!;���G<!������d��>�^�qi[ם�}���1��#|Q}v���6��bk����qx�r#��p�d��^j�<��b�S����C��Öc��.)��mD&s�h�kM����<���<�Mt���s3+���!B/�V5D�G�<uι�͌v{�/{f�5�n�0z�<�U�;�A�n�ҝ�m��O���SV��+��W���^�.x���O�*^ٝڈc��y�m��Gy� .|A+7(^^� )�O�r_�i7�<'�u'�Ӷr�DorL�o��g����WJ�p9��@VFʽ�d6�s ��=f��0_I7)�
����)=�jۃs�U�����%v��	�[�r�r��`���lgQ��F�0j�xt����������wqLCq{=�z�~�"�{|��?v9�T:)hѮM���z�ˣw�9��SS��[�Z˝3&"6�df��.R���ͨ�7}Ɂ�w�So��ƽR=i�ո�����{��)o�S�|r�JЩ{g?`{���G��{B�\S"�������?7۹�L.�~$_뇅�6G���^�����	�w�cˆ�p�f��[����re=��1j��c��D���V�6����X�
�w�����hճLcV�诼O��\�lۙk�~�=�]!�����|-���ݝ�%����Wx��_�sj}�FL�{|�����<vO$N�V�1��KT�E���{>r�9=��{ç.\d_�������_/b����Q<�⽻Břn�Ud_�BY�x���9�ݼ��]� {�F��~���&�y��e�d���x��j۫�1,]&/LWN��ih�c�.O��϶*��Rg��[p�jL�wJ"��x7�QUMZd�w{ �"���]��q��a>8l��"���o��Ӷ��[�_zwX��t��]����i¤ԋUp>�c:�e So~�H��ٿ���`����sc�^,Tl���KG�VF=�=1&�<��]C.{�Z�r�n+k��F���ރ���M�u���V����W��N���{g�]�,o�_1�n��&��X=��59�{=����ܽ��K���O��J��]���n�5��R/����u���d�£�{"~Qwb��?G|�<�n�M�a�7m���ѕ��ܾ�Vsך�x�h�N���=,]s��{��j]w��yoK��8
'��ٶ�>D�9L�G�v{=�w���bɛ��N��}걓��>�{�t�x>��o7�^y��t^~K$��ϱv�k�UA�҄��7f(���5�Azχ��3Vs� ��t��@)�_{D���=�M�����{�P{7�֔�m+_��c��٠8�K���<&��l���f�Ϋ�9d�ѵ����#P�ј��=�d^�&��O��P5jb�Ѕ,O'5߇QY�6�ƣ���o|�]]f�����Ctc>�Ǳ��P� x�/�r,�[<�3���	�]��k˝p'O�:}<7Fl��7}�{�\1A酂�h`��+J��{3��Ʃ�y��h]"f�r7����9壗酸�n{��Xf��]���-˷��ll���ճ�s��K0��R2���=z�m�cS!N[��d��g"��ncc��;8m�� �d���c�Ōs����q�ź/�G��$�o���(�aH��&}��]�*���`��X4�zsۦU����y�sm^X��i�.��$�-��t5�ϋ��h�h�ݵ�0�L;�T<���c�{�������y�g��+�%���v��\���o��ou}�w|t]s�;��ׯW�]�ރ�`�Q�k�M�&V����x��
=��5����}�<7E~��r��.��(hx`c�l��:��>oQ��xۀw=�oV6A�@�{D{�w�ۭR���$�xZ�|}��vBq�ӳc�G�=���@g��q�H�$�뽾�5�z������s�۲��1)�=�����}膗�	�'�Ƽ�R'w�:��E�<�]�C����D�*F
{�����Qu{��L~�n��Ǘ����U,������.�_b�0��F�Y��[�^:����y:��%��u[a�%����)s�'����_�u���w���|İ�^�P�=v)߷� �ő2�Wc�U���3}��s�+�X���9�M	�k;� W�}wFV�qy�䠋���;ͺu�\�t��FS7�ޛ��\"+�s�5q2���g��s����� =y�"��)>=�Z��;`��:�q���~~�ɝ�����U��� n��.�ph�{;"���|K���g��]�VU):�J��@��H]CmgتB怜)u��iCO���������VB����b��<z{/:x��w�W\����u�S���ណ����ض�����qc��k����^���{/%=���;�t w�r�Q�ð��|7h��N���m]Κ�v��xN�O��oc�,��G7�V�6V}yn��c��{����m����d>��p�+�{R���>�+�X.�f�OW=|vI5��n!�]}w�gX}?Yu:��e��K���8��X{F���,�<g�G�	纹��G�������)��9�t�4�=܇�{�F�����0��ݶh퓞Uqg�a�)c�|��7�a{����r��L	Ї��w'�L�6L��?'��@w7�ַ���G�Zc�1���=��pŷ���/���e����}�c�f���$����?����"�#\��k�ԍ�q.��b�U��s�d����nl��M��m���ļ\L������cGh^.8�N��U���'eM��	v���Bth�[���{rG�`�$�k��l՝��Mkͨ����h�i:�Ѯnz�7�ϖ�n,��u����&�t�w�.�lC�i�vOO2����|���!;v :�0���g��ܸS���v]v3�kk:�m����{.�ϵ��ۮ�է�/A�����gm�9��b8�^��v؋!٫�=�z6�!�qΌ�.���:�`F�#���h��e%#��-�E�J�</a�"��S�����ua��Ղ;x:F��kӘ9s�<!ٽ�(L�d���,��Kq�-۷t��l�Wwi��p��`\O&�a�۴gֶ㖎�O���//M�mrPnnv���Wm�n���m�<�N�vn8{`�Λ�8ϛ�>�>��>ѭ��`�uy,���vۀ{k$�	\�^��vw�]�WZ5ۍím�y���q�N�y�6+�۔���^|�]���`�������T<]����V�۪�v�v��cqvȏW�]��wa�;����]�*u��͹r��)�본�mnۡ-`�V.��O8Й9���\��U��.|Q�Ym��t���rm۔,��ۓA���X�U��BۭΫ�eݢ�g;"�c��mc�۞ۗ͸�Ÿsۆ:-vf�3۱�q���q�nz��l=km�6���y��#n��X�Y�f����Ǡ��*�f�e�W(q��^���rqзcy0���Gv���������Xc=4k�c\r�wQ�Mp퀋Ic�J��0{�ε���h8<���Ԕ�f۶����nWm�6�=k��t��	gۗ�ѝv����4`�C�1Z��Jw\�n�n�{5]KV=s���BZ��N���i��f�� �m��Cnz�+�%��r�f�jj�fۚ57g�;���v͔�O#�]:�)F���˹7��f��&�<�z4��H���ǣ;�)���m������#�Ԅ���5��;:ړ\C�q�fS���kFӲ�:�%�7"v�uۙ�'d�#�{�kOn��v�[��Hb�7	��ۭ�;�z�6zzzZ���Swl�����:1
�s�z�"��q�^�d�<q�6 ���<b�E��m�έۻ:��z��:��"vp�<&Zf��Q>�܈$y��ݹ�;����.R�Yx�.z��.7"v7���:n���ɶ|�W�u�6mc�q��Cu����n^L#��=�:�p��$�8�e�9޵�r��Q��n�m��˓/=B��fܜu��8�B�b;kv���n���F�u�ռ1v 9=)�Or��c���������I�m������W�mnF�ŇE��s9.y79��]�Yqک�7\�s��sё�<e�n��Ǫ9��z�b�6ڑ��]>l�9xUA�L�A����lu�6��ɶ���g���ݶ�S��g������v���������^5h�'+� �ْ�`�9��cvB7X����w=��'��9�<ŷ�{�k^�y��ٛu���qcT�QtdZ���Gu���q��\Vx��[h���l�ݩv�nBON��ܝ��,獍;vy��N��Ŷ��Ӱ]�3���ظ�=�8��]��Қ��Tqm��;��<t�k���C�C�fv�������]����K�Hc:��ytka�f��x2쯩x�z��gg񣺽[��ٖؖ��v�in�Tx9�� 4iw�z�i���{`v��Z��@�x�[�seqv�w��=���Dp=�͞���NW��;b-��^��m��r��Lqv���:�vg�m��w�WV�!�)����5'V�w[tbv��c�1Ѯä�P����<�؂c��(�e�T�,ns�C�V����6�g)���N#�;n&V^yÍ۟m���v�[m�\���㓵��y�i����:����n�%�rDݺ#��c�xQP���.zn� �c�uw�3�`�+�W;��u*;�N��R;;h����eݍ���jsկb�-`�G8.t.�s�]���q��s�{;s��p��\lv���ݱԆ9�T�n�5���9D���evI�ݗ��(�ၣ���6��#۵sҍ5����r���ȝm�GEUmeư���mm�J�=Ov�s�7Kݎd����il]����ㅜ��̃s(��嬧k �m�r��ua�p���z�ci1�M;�c���۳��s�����;cF��ll���x�}l�נ�[�ݑ�[�Og��{���ng���eE�N�nZ�w��K��y���;X��v�ʙ)�x3�]�ʹ�u���	=�N3����BU�l�q�@�Ƥ�4;tݷO)�u���n;q�9�c��3׮�&���n�F�1��T�G:�<�f�]�90��j6�mu�!61n�;=��5]��уp��e����ss݄E�Jw �r[{g�:��nL�c��۵v��:�TN{�#�u\�뛣[>m��&ܜ;��^��]bv�XUڻ<h�����Pb���-=!m�X��;pxݔ�Y�i�R�T�	�����{k�Y�q+��^g����իY����`l:�Ӈ�K��ɝ��ힶ�ǇEj�3���c��1��s��nM�Y������V	�9��(!��1��c���n�S�/=��Qz��cr�O���C�zr��o�`�#�1�7��\��v���` s��v��������U�n�����tݦ:��l���la:�6�8�|Cg��ӻ����ơa�	ts�M��7��8Y� %sѵ�1�xݔ�ִv�К:�2��^�뵽�GP��\pst��)ˠ�+��n=�h%N����vΤ��[�;��n��-�]�睱�e�;��]v��<�j`+�qgznב�uhb�l��v��>�Z����zw��/s��y;/=��^��n2�75�۳����c<���f �۝����7[cWZx�/��M���b#�\&wE;�uOm�ѷcvb��/<��Jqj(��^y�պ���y6w�6�q�A��r�O���m\ь�{[�v�z�ŝ��v磶\�a7@y-��N��kE���mٺ�oWO��ճ�P�I�sϴ>�b���gc<�.����m��`N��x���ۢ�z�8����1Ldf�M��1r�+Ņ�ʖ:딳a7^��i�WHDv��e�!��Ys��uu��v�f2�r����a6#8���'Cۻ�Mن7h7\�OZ���ڶֹ�s���]]����d�D�[b�gכ�n��������'v��ptc2�M�8���W�s�I�\썶�Z�t���ݻg�'���ìuױ�]]\p�>L8���`L�_[*�����c�֞;�ɐ=gw6�'-��ە�q%d���γ��s�66a�{7Yژ	�fű��G8��b�.�z�"2ylh����]v�� ���Oj�gWk�1��z����i���f�n�۞�PnN��^�����	Âc�Y�q�؞÷eW/c���c�t�kҢ�����q�Y;)׶�^wC���[a�ׄ��̞�U��l�Z����z3�^�8·4O`��Pݮۣ��ls=��h�;.�m��؛� ��^8[�8�e%,sn<j,nǢL����y����Ӂ��ӛ��.q���k��O��¼&����+�H{w���Ǘs�Nx�Wn'�ͺ�-u��.��Zm��g9ӧpg�_�ٶ�n�d5ҷ��m��*3V���oe�����6z��
���@]���6\n.�9�
�t	s��3��1Ӷ�&=��z����x��U\��z�x��n9�EŞJJWqW>G�\]��m����}���Z�ܕ�z�&p���:'d���=9H�1�GS=�����Қ9v�l�S��nm��<�Eig���g��^���ֶ�9�����[��)�x+���Ӄ��Wf�#�u��x-LnpnU^u؞h�x��d6���σ���m�������v�n��V��+k�B8w�7{;vF�9"+f��+��՞o�c5̙��^�0��-���N�9b�;Zӑ�wZ�c��Iu�wQ]���v�<��z�ζ\ý�d|��,kIv�n�6۫'g9w��<X��}F����;u�{X�gX 8�6����	ǋ��:ǮW�XU�FN8=6(�����gFK��x�>v�׎<�WY�խN��&I+����}e�rqn;s�뎳ݱ]��:��kɒx�}u؂��h��n�ۇ�%@�����/�njNץ���,xy�m�Uӣ���f�L\�%��(��R��쨺�S�5�b;2�6Vy�ح�=<պe��@pj�mY��C��G���N8݌F��s�O)^��c@�����z��Ge����b"�Zw��盔1�8n*w/n���=���v�E���M�l�ݎݠM�Íβ�=�b�ՙ�ܝ[l���n��z�]"�h��	���:kq(<�paM��s;G&v�n�]�:��<�&�9�l#ˡm`jn��n�V�Tv�v8��r�/n�n�m��0mV�ړk*Uã������=�X����Z3]i�u6���Z�׮f2/Y�o<=W�8�nhθ���D��&�ڮ6Ee�t�/-�{mۮ���˶�v�5�j��CqE���b{K��m����]ۯj��v���n{6�]�pp���<u�t��n_8e0cѲq�:��v�e#���.���m��񣓙��ݜ��s�a�����9v��8z�GR<t��k��sǋ\�D=����FV�U�2��9��"�ϰq����Q��`��su�GR��jNh�20����Q����̈́u��Э�6��7
�]�����v�Z]v�RaK�h���.
:�ێ�T�?-��p����+��kF)�QP�B"+iY"��`*�j�
+ �PX�a�B�H��+E��&X�FҤU�E×J )b����*E�	*VVE�a*Ep�+$02-eE�Qd�#im����1�,�sa���ES
�	��� "�,��#
����U�Y(�EYYX�Y
���"�$��%E�A�02iZ��1l���(�������IZ����Pq@�Ub%lQ+
�n1*9�D����VH��,(�jE�Y�bƴ������*��\\b��,Ţ*��LR����**%Dp�0��(���q�L"֠a��aR�UQTT
���Qr�����D8��\8pa(�,*W	R�a�J,+��ee�b��D�kEū"��ѕ:���=�:��nl��V��=n4�$ng%ohc�n�ܘ�+ζ�u�'U!v�׀�ur��W;tc��D9�@��vr���b�&6��}avH��`4ym'6�9N���W;�e]����v:;��H�Ѐ�sh�v}�ՙۖ�S�a����mA�7%�������\ر�s�3;��u�Q��4S�-��UM�q�Ǝ�����ΰ����M�^���&ۭ��;�ult�(�T��ӆ�eqC�M�Fޱ�FNyzk.��қ��u̼�[u��سݶ��X�:�Is�`����lki�����]��zr>{uy6v�;��m�e�O@MT����Jn����
�Ǭ�q�xx`Ȍs��u�HKdݭ�3�i�5�ݰ�OK��Ʈup`9��v��N��Kmu�O]�lG\nQr0�7/4%�`�ur�n�m�n�;v����M�\���ݜ��E�8��=��/�����/[�����l�7a �ʃ��u�I,�i�Ho=��5%���1�������v���1�b�s��Y�T87�����9�s��9����;7�99��V�X��ts<{]k��Z�֞�W��W3�d�-\qr��ob��D��q�nj�:d��Q����y���x� ����v*���燶��u�D��t��G ���]��[��Eo�tWh{)�o$a�'1ۡ3���u��s���"d��#�7����x;;��]�;6C�S��nUw��v.��v��ڞ�q�z� �tKʹz��Q��x�m�br�i��F�\���/��mn���n��|�ό���\�����K�h��d�v��m�VG��m�J��81��Cl����:��Y튎���fSu<�̏ln��<�z�3�^�v��ٖxvq���Gn�������ݻW�u�m�;��݅�d(�`��RF�6���>3�<�.y��v��oD�Vt�]5����=vM��v�v�a�2�˰s�g��s�]��pq����;l����gc;v���l��G.�gq�;���xq�M�rcv�eȜ��g��kK���p�p7 ��ѥyw�c)�v�/s��;�U��i[�nJ�)LTÁ�h.�p�N]�a�;��L�e� m��]�TCo	����L���(��q�{x66|;>G���{9�s��ʛ��������q��/�I,z2_{�?���x��v�o��/��ʹ:㐓334`EGA��#�y�S� ��U�u}o;Ȃ|K|�D�A�� ����.{r̞����@���b`M@54f�B�Z� ��/"�$��h�ǋ	���'�^\�=�L�P�&b(P����ް^isMoJ�]��$i���|	�ټ�$�k���b�(�yO^b�N�$rz�=�AU(��l��0�Gі�m��4n\)���b��U�v�Y-r���gz)@_QD�P�I�su��X%�ݮ�tݸ���1^�#��r��P�����{LԈ4b6-u�A �˒+\Нȋ.%�'��Є�� H$��+�6�a�X+4[�������I��}�ٰzz�b�v=[�C�"�c�s��O����=��}�4����w��x�ZDF�*g�݊Օ�9i������	=!vdN�[ �H�8��%Z�$1K�g֮�x���}.xQRL�@ET�,Ӆ�`�v�4���9��v�*���OMX �6}���%�L�i�JIW5��Q55�	.���>-7h�����u�B�{BWF�u�듌*Pfb�Q2b�
�=��y^�v���[KgL����|�s��$�OR�>'�ʹ�X�2��n_�Ca�N��X1��a=��yXv�����͆ۥ7������7�?����MG0c��Y �]ֈ�m�+:n&�+ڿa� ������@1߃��I�8M@Z�}ͨ���ᐞ{ӥh��ı�A|�A��ė3��G2�#D�SfL��&R)k��I9ͻ�K�?�q�J��ѽ����z�;_���Sp�E��=j������_��JS��y-(y�ЦAe�L�z��>Y��ئ:��ell���ɛ�~$�r@�{�v�H�*�	����j�A�]���n;X�rf��j���|���b�QYq>?���������KB8�`�I-I��j��~���a,��ۖ�A�۵�H��d��U�A[93M�f�E��������x�;j�^ö;h�g7\��8�\wMMEWh�q1"�
b�
�<Wb���ݢI'���vuf��[Ix�O�������\a���jg���k����I���	V� �$����>$x�x�_�V�4��u��~�����&�E���^$����䨲K��NDV^�	|�Kē��!	�:�UV"41)?	>��t}��3�~z�Y� y�kĒ�6B���5cQv�L�Gu뿞{w����N�n�U@r�{�x9����W<�F�u��^K_7c�}�VԨ~Ε{&�_}������V_���z@?o�xh)�S�Ђ$�ܣ�|v�UB�Gt\eu���e�A�b�_��4�r�����������������/n7�\q������6Cb�ܗkgnpqx�p��\��~��ߣ�!cm?>����@�H��M�J�� ,հk��3�|��!�̛��0(H�&(P�������֫1�Rv�;�I��M�O��i��QۊGf�n�
�t��tB����F*b��,�)�y�Ȃ|kx���#�+"�`�K;�b�*�;D�pWꊙ��"h�[��\����(��߈>��h K�m��q��IFq]l�LUP�4*H�H���#�H9�h�"f4��K�Λ�B���%�nL�a�5�Q�s��b_o�)�T��9T:a�B�����,q9���=R�#y,ه���i��{�NTU�f�m��xU�qn;� XC%��5�&U]J�a;[[ٚ���6趦��v��gɻ=5��K�}�2;��$�N7��mMv�ko�:�Ƴ���s<�1kt�lmoOj�6�j��t��rC�٫g[�������Tv�<�z��Ͷ��x� /]�W�p��yܱ��s�L��I�:�,v'h���-�pč�0i�`��t󲅻���c�xҙ�n��mӅ�gt�v;3�W��kL��[V� ��::������?O�Ӧf�"�LԂY�����4'Ā����Y̗ۗ��Q�\�
��>H��m�(0&$�},�`��ɝm����WY���A>$j[��}��H`�Lb	��K�F]جсP�$W�(P��Z��sv����à��v}�'�	�h.�1cE��f��R�fv��=��#�n��$�m��,��Э붞&Y��D�Đ'�
�QS350LM��cK���-d�dM&�iJ�N��A[m�|�Yu�r���U~��7��(cX���b�	X�~I)��B��5���h�9K<j�K�������u�b�:gYO�I5�h���l���9S绕7U���<H'y�Az��.bh�Q�5 �2Zٰz��1��]���� �6�O�g�xh��K�}���kl4L�wf����Eĕ��3���y�p�3��۷��\�C����(Mz|���K��"A ��]yu7�M��-dK��x��sg��2jb(�4RM�Dud߈y<������}��%�|H,��E��H�
+�hP��ou2C#iMEvX"������M�H����2r��Ǯ}&O�|e�M�9�H�=s`�I���m�F��[��	$-e��$ZM�a��ő�ٕ}nN��ηR�A��3 ���n�{���f�N}s<3��/��Z�Y��}���L,0O���$ ��D��K��8,'���������~�m[D�I��}g�������+��}7� �9�
K�D��7*q�]��1��`$
�j)�XxSk��.��d�d��~�~��xc?�r'�۞R�6�~G�,>�^����]#rX7:<fVݘ�]u��h<�>�w|C�F�:v���h%�}�yB�IsK���(%�����}f,�S�~g� �I������<�U��l�!;�g��$T��Сg����v�0��яG	�$w[�����C��k�eP\uM�$��yD�L�(��vm${{i�˸wܼ�o����q�qOc������}�ݦ�TMD��Dc��>H�	�>m#���FY��{�;K�}���'ܸ+�EL̊�4b/�;ix�pf����r���HT�R �	�����/�x�=���P�iE�XJO�'wm�q�v�Y�&�N�I
�5"A-�ix�C�E��3"�UT�6m���s:��A{�/An�א[P�=$�/�}�g7o�^���T�M�wi��E]�t���T�]S�Y�#T�V7o�����혋o	׃ۜ��:c����(�͐Lu̇�yV�9�(�q2?4���~� �P�Az'^��	[I��#��HO�t���߯�~��n�;�֛���]V�����n5�=�q�h�֮S��g�W�{m�	??{���tݷDСήMA �6�Au-E��>9
��`���m�'��-$�4q��R�{��}��h���O�2 A!�m"I�5��Z;ܢfр���Z�;��fIU(&�/�_?��Q̴�_E]^��|/�>������H�1�|Qx�2���K�Q����y��t��Y��'����yE��H	_5Th>�؏���l+ϻ��K��l��ے�x�
xM�C��8	�|���������{������d�v�N�čx��#|t�#�Ƕ�X2쉪F*�����P���)D�����ÇgZL�{_b����X��ڜ���P=��Z|P��xӵlO*�yΧ��g>����y���u�K��zͻ`�,�;D���\g��	p�Gb7���`�D�����gl�ɎU��\���X�(q�t��ہ��a�\.��u�	����{ *�B���l�[R���t˺�{�k�.��z�M'�3�q��l\�|Gp�M<rn��뛗w<�M!����L�%�Wg�n۔@#��s6��y[&��v��aɭs\�]4�@���Z�Q�<��*�c�s�}�����6=%�o����� z�U�>$����;ӼmodEg��r@���I��C$����V���><��J=�Wj�7��I;R�z�V�;����3ݵ�����w:�	��MTL �&�O���#�H.M�{�!C��H.���J��\�+�T�̚�"��Nڑ
��k������$�F+�H�[�շZ��ԥ.�����7N�Ǐ�h5��_��j�|ݠiɡgL��yH$b��/�з�/����&hњ5X�c�5˩��su���<V��JQ�;mI�mDnQ.�ϰ/��S6����� �=7����-�ix�V u�Q;�:����$W��T���8�; �o����`Ç��V���}�%������y�.�� �٭V��`~O���>���~ǝ��f���1��X�̂KW�a����&3�˪�6o5����`��EMLMA��<��I/�v�H$�5�{��n���'U�$'�7h�B75 �����+�v����7�	)�b��Fo6� �9�#���s�\�ذo�O�}>ɸ�D�Z*��m 	 ��Ջ�t-u��$_V�%�m/O��j� p�=����?�x��ڈk�Wl�no/c��S=�w��50��֫t��۪4?���2OY���;�ƈ$���I���:��8hzkSA��a�0L]P��&j�D���%OE�u�u��D����D�.��&[6C;G�r���`��ΓMM	HSOR ��Y�W�>'�C�r�!\nUH�_g�eh��oe{�7=�������m�zm�u��1��_t˅��z��z�Iw&��*��y��}��}��M��^=[S	��C�9��`(眹Kf�Z7{��u�z�
���M�)^b�[������Þ�*��?�-qȸyb�^���]��3�� �Ȁ�T�F5U�<��xd9g]|���Ea{s���ˆ9=����<`^ZQ��K�S�ʙ)uWtF,��^��=yq� {l��Y�2=��JN-�>
��@/}{�͖#�{)̟7��_����f秐�^�̐=}ß�j{��s4�M�a��P�N˚vQϒ�����j��yZ�os%��!p�:�e^0�'g���k���C�#��v�M��{5'٫��g2�M��{������ݹ� ]����;�R��CoabQ����5�C���i�g�^	-�&�"�u.��\to�:���r�Y����<�V	�'M�³��h���9�}]h��uW�Z�Y�NKU��:'e�pt�)�������a�)\'w�r��4}�1	����w�a�=��7P鷪|v{��='�]:0�Z[�g�ůo�Ȓ�U�y�}"
7�����=���^_�m-�r�bK��Nk�43����!Y�h���KNƔ���ȏi���zy�;�O(������>[P~(�]���²I����#�vqu�&]��1�W��.��r�ݡ��񄶤�j�?^\b�e��1��Q'7�q`��C^�ׄ\ަs���L���w�ܘ�dPP�Qg��q�\Z,X%�Q�*QDEkT�0�jn,ia�P�I��0��RTQ��(Uň��VڹH��m!���CT��(��Y1i2̦sh&�\���0�,0�#i�\�P��f�� �Řń�AaP�V�^Ǽ�G����x��g{�E����h��v;�+�;�����xg�p ����I��L& �e!��,�eC1��4�A1E�
E�8�Qł����%�.0[L "�VJ�E��
a�C
�0�TXT-��"�0�a�B�b�U+�U��D��%L!KL�.(�(�ap��03
�1J�+*�qi�T�
�����`�0�fS#�2�9�,�*L�(b�\%�h����P¥I��S
���ݎǓ���<[%�f��XTW4���ͰP(�;����|��Ax���_��()"��f���VەU�����
L���x����v��$��6�b{3ϔttօ�{�������o~�m��[�b�!Z|��[H�6;�瘑 �=n�(�oz�+,�L��v�۳�@����s��u�m�qx��T��׋�.w-O�P���^�HL�(%Q�����">���t@ �\�=f��Ը�3&/WL����Ğ.��;&�Ԋ���L�V��5Z�C�*m��N�$�Ѷ��$�\�G��!]v�o���R"[6��<&ո
�}?L��)����'�a\��,Ϋ���;�J��$�O���aT��9��ϰAmآ=Ky"I���v`��ӏs'��_?��n��>�V�����Q󋟫�w���||�u�����f��jvn��O��)�|X�&k�폢:z���X����^34LD���@"Im�
�X'^�&"j��*�j@�q�X��(��wr7��Q0@�&���Z���ۮ�bx���1ͬ[�ܛ��=����ߟ�D���-��*]�I�[H���R�bfz*S�R��.^U&"�LH�6x��d�҂��*�I�U.iH{��q�����~�}P�=�¦�m����N�]�su�D��$�R�:��^ ��kH�^�i@}B.�A�SR �j/u�����M�N��O��v�^G�*��Q+���z��� Ep&0�3�`Q4��M��I&X�������I���^�4�!�yb�(��O�:��wg�sasB�4L��]��f���5�����->6�s=���v��������R1�����m�Cg�p��}v��w$��wU�a'�=d(�^���nՠ�:ݻq)���{���6n��˷��f��n�{]Ŷ�.Wpݘi.uo������F��äL��s��������W���i�Ֆ��4ݿ�;1��nvv9s�۵�>@݇�]îՎ�;;X���v�6����ٵˀ�ø�m�ػM��<�X�6'�M�]2xN�����N�-����7�>�@�wLڿ������$W�&���z�~@�����K�y7�-WH�Zn���ѽ��^$=�i�Ln� 16¶f;��0`��To}�"	'ٺ�@�If^H�v����{ķ�+�T�5$ȩ6x�'��z�lA�������@�C�myqY`I����i��O�R	{��\�\�����K�|H$f�a�|H�M���"�`X:!�z��_<#sY!<e���=Jv��kP�nSsX9pn#�y��=S����u��Ns����/�1��EѺ�1l⌬����;S'W;�ܯ&���{cK� %m� �c8�8�{����@/.�NRm {Q�9���f�����*�p��f�ș@?Ħ+s�~����o���Wr(�Zݢ��*H�{N��p���Q��d��1%V�.&��TZ��nT\!4([��.��q�f��@�Pw�4Fj�O� �.��$���/vʾ�YR�Rܭ���'<� 16¶���n�9���ӫg}nKsz�H9;8E���׉�P�
jI�Rm��m��ݡep�Ix�.	)kK�ۭ�`�uE{3���t���v6Zl$��N���0�n׎��B7��X$N*�`�W�k0g����
d�}�:'��XJ	8CtN�Xw�\�����͖�\@nѵ�<I���ֱ��8.��5U":�z� ���$�hEa�|��9�����"�j�$N�p�Q%�x0�'�O���e���W2�A �F�z�$��[A�d�c������޾�Ծ�O�X2��M"�wr���s�H�.�޽H��}�$���]&���-���g_�{�qoF�$~�|��Ba�nIow�nݚ���à���`7`ڟ�·8�A�+�Kē����;:(ȂD��h�7p&c$��o�񗷖>��iA �s�7:yeHݯd,֑֠�0�I$T��=m�;9e��J5")��M�-Kă���'Ă�X�����/�pϑ�8�7�,K����/0���cT�c�ns�nl��)�,��������������}�� �����A>n�����ȴ��$���|D�>�>��YY*!߽��8�%a~�z]��W9���T��;����AI{����^��?u��﹣�8�P(�����g8%`X�k�o<���@��_^1n8�J��:��q��Z�幦F�\��M{��G�ed�������0�IP�J�_����ﷃ��1��0�0�+
��{߽�Gr!Y(2�VW��y�7{�<bܷ2��mvaq+���`=Q���q�b�q>@0G�z ��ߴo�����`V���������>�g�_�(Z�ʾ��+쫈�Oxtgݴ���X�CxN�;�lv�����O��S�7��ӥ�{�,���*���cw����>���@�@���C�+?g��w)����n70�
����$�T�
�|߿h�g;����'P>J�I�~�ݜH,F�(���<���H[,7����Ă���2#������?�"����k#��= ��׷5����7=]�������?������qs��78�
�����O VX�Yc%g�w��*AaM��=�q �}]��v��)�Q���a�@�<%#+��<�
����v��s�8qq��g8%a�{�0+R�?L_Lw���ށ���ߥ!m!Z
����T؁R��'w�wP�AgJ����1�s�i�C߳�h�IXSS0�*2&�ET̈^|�����>0��R��wGĂ�D�{|�;��W�ׇs�k�Ԃ���]{��nb�m!m�w���8�^L�����i��+���r$��w�8�9����Ok6���0��������P*T*J�����a�aXX¤�{��{Gs�G�{2m�������Rm0�Nt���7.p��L۳���{�0(5!m����|)�������L���
�����7*T
ʟo���q ����߿{G�JÝ��D�֟Vt�>o�����2�;��_^+�Leܦ��3���TY���%ǣ=���&	����7����'����;|��'�����É�o@,M��O\�{n��o��V�n;FI�9�qٍn��.-����厵�����N5��셻���q�I��v�Kjz���;��1�1�l�����'�p�};a��)�w��2d�v��u��������d�||s��r��'quCon�������SÎ�Cg[y� ������/m%��"qj4l�)����M��]��mt�ѭ�����x�[�vwշþu�r�Μ�1��9����c�SS�n�XFϾ��a%�T�Þ����3����@@{��0�0�>�}�O���*�\����j�H)��w�u�`V�~�ta;W��8�
�I�{}���@�����=������2���|Ʉ($����~��Ă�RpO}��h�N!Y�>��D�C������/�k��~��� 	���_ɜ8��8ѴD�9���A���!K@��߽�i�!Z���ι����\aǷ��*|�R*{��ڇ�J��P�{�߽��q%a~��v;ɑ4j**dJ�������*�e'%߆�
Aa�?�����%��������%`X�k���u���p�+������<
B���w��
��G���Õ�4s�N	5�{�H)�H�'Z���ޒ�[�.��U��Ĉ,>>��Ì80�(¤�w�����8�d����g��`�@�����7ߝ��8;\�Ԟ���$��ڞ�k��9���siB�T�>\�q�償����{�s�-�9������G�
Ԃ������!RX���]�
��9�{�c�{�� ����u�~*���h�VǾ���%S�q���q�s�`#�$z<G�}���VS�n�_��!�yFQ�u��KQ�v��7�7����'7;M=��1�w
c��yq��"�Wvgl	̴r:�9[��������<�2VT�S����@���Z��_o�{�R�/�����as�7�����X�~�u0�7.+s����'��~���ed���g�70�R
w��{^�ֹw���u��aF%���{�I�*Ad���շ�"$�#Ӄ�&1B�b���C��;��1�����y���H(���F�)
с^���T؁R�>�K>��0�+)grg�ϳ`.���3̕����V���y���q�c8Í°�
�����q�X!RQ
�;����q������m�pvq	P5�o�6�ȕ�cXk�����R@���K�����WBb;��]M>ۮ�s��
Z�q��i:-�j�6մ�g/X�Dʜ��E|�}���rF������w��\���N�2T����@�lIP�J��\��0�
�}�yn����g�m���Ѵ����������a��6r��L�˜��ф�_�_Xp�0G�3x�M�>ţ\� {]�����-�*Al�_k��R
A|.��~�}�ނ� �/v��s`cZ��8��+�w�q�Ʌ1ssKw0�¹���A��
J!Xo\���J2�X���[�Lv�\_��I���K#�w�F.��;��Y�ϕ/s���d���N�H��;W)"���9��Er��(�f3�hR��&]T�F6���+��F����o�i
�z罨m�`V��ݷS�1r���p*��~Ѵ��u���G����gJ��\���F�0��
����}�ۇq�aXT�=����$λ�^�Z�Y�ଙed��s��Rl>���nL�8�\����{��`pjB��{�ag����ϝ���1�͟'���
�SbeM���jg+(�P����a�
�̉�"�'RN+���ٹ��y�c���nIۢ:�ױ=o8��dxI@��*��M��H/�a� �_��2��%B�޿w��3��P(����� �DJ�siѮ��8>����nb�m!m���{P���[�uG�;�p��0c;����\�����@��1��Ξ�K��󏷞h�d�IP�+�s��8Ì+
F����6�����h�������ߵ��4�:��'�@�<gg)���3L��q��m+�����x��R�{��ѾJBҐ�w�no��`�{�h��}�N(�YSz��jg#%e*�{�h�IX\{��L�S74�p�0�{��A�o���7p�AI��aϻ��8�2XʁD���{�@���F�,k�{=�a�y���k�����m�;�u/茱����ڮn1�SGt"��{���G�哾Zt���,���\�4��uO
H�B���7� �<	��{P�A}�[��؎3mnq�����6�+(�YY+�~�tm�
��fe��9�}zH�'�gsZ����aP?}�}�i9��� ������@$ظ����2���\I���SQq�=���𝓞q�vqe�v��SF�H�Tk�:�I�Ρ���55Rj>@�=y`r<`Q�
Z�{�h�
B�HV�
�{z��T� T�9���s� � ����P�8�R
C�߽��!�%a�_�a��q��9��k�B��0��ϵ�
M�*M���݆�c��g(ʁbT��q�T��_{}֠l���Nf�׳�{��o���C����9�[��	�ۋ�Πm:���i�H,��^�}֍�T*J�IXc�kǹ��~�>��>a�
*J��~��8���d�ed�����Rm*�1Ô��g�\�8�P7��>ߴ��m;�~�����hk{�򐴤*Ai����@�P+(��=�C����w����|�2To^Ȓ��;���L)���[�q�W?���aQ��� @��>w����-�栩�o���R�o�}�@���Z�_��5���l�-,7�{ڇ0*�2k���i��%kǋ��_��,-g���c2�W��Y��y����Of��:�bQ�[����W�e���{���w�3�w:�nyɍ�%�ݳ�R�x�OM�ˏ��=~����f�+
咷T[ ��~*�y�J�b��n��m����X�B^�0�����*��߷|��M�O�Wďd>���H	[�n���%�-�jS��_V�f�ezf>���=�Ƿ[��^=4�p/��$7��
�MC�׹V{]��L�]ܣ�����4���F�O��@�y<�oǧov<�>�^7ݑ���J;y�)��y����|��<?v��&�d��3a�n9
f���qMe�6����z�������y�`�� �K^,��H.{{ݳ6�s��K;}�T@Q� u����Of�2J�������4,���̇�,.��O��:�t��!���9����6��O��.���?�
��J��?d�x�����$���8&���q�%58텱a���f��������B�-sVA�p�9{F�8w݃����g�eKNJ�%��%�9<���=��^�V.��\+&�]��m����7����./݃�'��郓��9��d���>=���x�~�m<������[�"��w:��^ڽ�}�#6���L�꽁�z��x{pY氊��f��'���u�y��J����z�wJ��-�}ΎK�ޞ�=��;���mh���sjݏ�g��]���D�y�;{��>��PXu&0���`aRa�����P2�QR
)��qC)2� ���DXT�
�C
��pȢʩ ��a�db��i���6	��m��8#ܝ[	ܖP��E&[�B�,F���̓s��6�V.FQ��fb��e	�DP\9pb�%*�(�[e�Ô�Y����AAk.rRT�aX�F,+X6�Qb77\Z9n3Ha�,*W	+8\P��J�CD��
��Q�&QdÆE�	��)1��"�4�W�R)1
�X�EJ��&srJ̡�a�X�T����8���K����-k+����a�&\1�T�`��YPF
�
�+%fY���b��J��[���)jʒ��AeC,���۷w������{nVv����\��]g�.������1��m�����cq�ҳ��q�qjܤ�n;rYAk=�q�M�Yx��4�on�I� ��ۇ��{�[6�*����wVv}M�u�;��;�t�v�{�����{7f�v�Hu��q� tk=p�zx�zP`��`7�ˡ��y���6�{y�d3gu�9:����'OGn�����"Q8�.Е��vue֍����6(����6sیbM�V�=%�ד6�N�-ǭ�,<���)�;/�s��H�]��#ٟ<tq�Ӏ��$(�+�Sz���6\y��q�\W�ֻq�{M�az6M�]�����Fngnݓ�d��'j�ګ���ɵn9��t!�I���CY�!��l2��m���x86�9n�f�ݎ����#m�UnX����z螞q�6�\e�tv��^x-:�!��p�Q��IK��x�,0uX�ݞ{g�ؚ{G�u�=�V%�]SՕui�n��l��C��v�]vϷ%�۰۶����G6�4��W�p3�K�ݠy��痨���ѹ������c=x.7Y\e�;�˷6�$�9AD���:�b��&���.�6��������Nwl���:�{5��o!۫e��t���ci��q]h��K#b�ڶ���.KփO�g���n����$�@C��;����[m���[1���{]'m�[,�=���s���wj#��t7��u��M�5���q�$Ž��8:�fK�6�ύwHa�K�^|��M�qy�h�n7<�WPt�:r#��Бz#�`�H@�B�}��wa�S�}��s��y�i��/�ݳ7y_F;�9 9�|�snGuy��n92yك[y��7>s��qۊv�2[O�&D�yR�X%�tyN�.�%�^[^!5�6�H0盝��h�GX�ݵ�ܼ�M�;nf9�n:1j��;$�=��mi�p�H>6Ї^��v�� ͓�y�<q��7']�UpFKk�'�4��{��j�X��:��9�:q����3�ז�&2;&5�V9��Z�5v14e��Ez�6۸Az�,c��˸-q�죤��DP�mt7X�m��\�wYn�qع8v��v��<�W
�݌m���k�����M��0��w\s�Ō��������ػ<�lbn�ݸs�ud\�n���pwnyֹ�;�wb�R9m���ӷbM�d��X���1��1R�㊝�1�-����NS�U�I5�8rD��&� �O�� �7���@��%ed��w�Ѹ�P�J�O�,{�����A�G#�-��	#�O{���$�����2���kRlJ�+lK�b��Q��1a �,�큇��x|�:��k>X9�+�}a`�JB��[�w�� ��+*o�����<	� }� ��k-È|��j$�)�����s��q���H/���h:¤�
��Xo��چ�82�� �x�����FU]	��� �|�`V����P6ZA����|�}�q���V��)sn-Ì��Mo���"�oƺ�ȯ�'�}�#���밁��(�������8Ã
*K���q&nL�^w8��^��1Y+���%��V,��T�	��M%a����x�R�=�w�7�������V����|��߀$ @E@������8�2VQ��P���q	+{��w�0~����:m�.U�\a���<�Zxu/W�=�m�d���܎v�X{g��z}��qssK}�<¹���A��	,B����w��q�d��J@���#���y���M�|��>|�;����R�!X}��چ�0+��s��_�3mnq�6$����8�)��ƺ����ۛWvb�UغYF���� v3�d"u��v�����ɬ�-/o@�>�ϐ�����fON��{�>��v���������I���s�̘B���?s����VaP?���m �r2�9���V������ε'�I eٞ�dԙ�3Tb� �|k
B��߽�h�
BҐ�`U��qή��@�9+}��P�82VVJ��{�}�C�+
}�<#I�L$�S�� ��o?ng|��/����:���IP�;�~�Gq �Q*����@���cX�ߵ�����^�a|/*~=� G�f.�H/&>Ѝw�����w�Ě߻�N�d���ﵞ��d�k����]7��Aag����q�T���~��}��8�d�������{�6&�~_��۞̉?}�QU5PR��ծ-�΀�(�7F�nGgF�ze8N����������q.p��7�@�J�y���jB����F�)JB��{Z��B� AvwUV�[S��φ��z�����(��~�q$�)��~>�\���m�8Ì+�}��60�J�I߻���6�a�{=ޏ�8�FT
����m�T�����k=��������{xu������w�q����ܺ�b/f3mnq�6��繣��
�++%}�Y�H(X��g�,��ڗ�q��բr6c��6�:y�^��Avl��e�器�y��^��.�`�V�t��~$s�\f3����=����c���		����0�V�ID�����GpB�Q���W���d�B �=��Dȡ3B"h0�0�>��6��[�����4xD@���	 �*Al?{]���
�YDǛ��a���,/�.w�Y��D{��>�yA�?;��1�b�ƈi'��2H!���G����ϟ}_z��@߾�vq �85 ��������|1��~�v�Ө���1�A�B��ᬥ)n��Rq$�����ֻ��^{qq���N��6��Z��7�F���.mŸq�@�xI����q8�YY+(�^��rm�hQ%B�+9�wۇr0�;���?w8�=��ϡRv&=���Ă��������s&�h�>��3���b�7e@ؕ�����Ç�A�<�N' � R���B�HV�ok����H,��s��8�2VQ����75Ἶ�]~��h�Aa�3�����G53]Ì8+�}���m%B���a�s��pg,e@�T��y��{m������+�X���sa�A���ß��jx0+��\��q�ks�@��'��sG���z��翀�������f��IP�+����Ì8+>G��>��c�F�<�7�_�bw��h|���{�^���G��{V�l��˱�jz�o�{@��C�.��x��_.���T֗N���=����$ ��FVJ2����I��������ܗ����p�����Aǌ
ԅ-{��a`��H��mtQ_����N����e7*Ae��}�q�J�3�@�@}���0�A�ٲ�Etu^Ti��scC-G]��+�չ��*u�m/nC^C��z���Zƾ���}%)�U���c��۝����I*%B����r3��e@�P/���l�"V�~k��_��l�Xk���j�R�-����ڇ
�c�ӧ�nmŸq���q&���G�ed�r��?S���8����(y%B��/��na��aXT�?}���Ă�����~�cwi����{�@���x1�8p�f���w~�6�R�{߽�|)e![���9�8^���s|�S��+*w��ڇ8�P=��{F�~��TB��D_���T|����MZ�������L!R����8�2VT���~��@�V��_��}���~3��;
B����ǃ�=�wXp�J�g�8�
�I���4q �r2W����c&������k����+
{\��Ì80�( }������ A�\;���Y ��4`E�b��aO��e��;F��v3fU�^�ج��^u��n���mՈ_{�qD{��=����=�I�$bᏴ���m<x˻�Oa��������o���n���!��i皲X�;Bc����A�͎���n{m��{a�p��;*=�D�Ջխ�x�z���.����`�^�����ƫO�v8�"O�kнK�p�2�`䭝���N���ݎ{g�l �t۬M�t���f��t�n�7l7
�q�p��q���Ј��ħquی�.!�۳�ӝ�oZэ�L�q˝���26���<������ݶ���\˟d9���콮�|v��X���r�n7[�]�l�`�_������q���� 	X~�=�0,jB��߿}��!iHT�����@�m�
�j�z�?|28���~��z�b{����8������m�.s��1����R�}��$�&~�������~0��k�8�2VT
%@����m�+�`V���wP6j�m�����a�����g�`m! ��-͸n.3�N$���h�q��T����u(m%Bĕ��9���z�y��*J'���h�N!Y(��Y_����6�@����1�7�q���m+}�=��<�;O����Z���=������H-�=��Sb@ >�C�߯��s�q���S�� �g|�4m�+���?�%\g���Ă���h>a��!RQ
���w����g����y�x� �w߶q �8��_�o�����B�Þ�}�q �����w~���p���Vu��v���nֱ����n[]�/d�b��]A����~���#�5Q*~�@ջ�@� ����i ��%ay���xa��#>�wt��Y�F���0��VJʐW�o��i�
���8�sn��K���V�?wA�����b�w9�UZ"n2����MAP���Vqn���+(������w�U��.��}���rq���_Ʊ��j�I ��3߷����H-�
����n�h*eN{���8�2VX�P��λ�ӛ���{_h�IXS�~y����q���L�p�6*����la����X}���8�2VT
��~��{7���y�|~@�%`Q�
5{�����!ia�w��8�bDM��
	�I��Y/������=�x��n3�c�:��J�2U��~ѶM�RT*J}���8Ì+
��x��X�=�?p{�Y�w��Y�}�FVKW��u&�hsqw��L8�.3vT�X}����Z����{��o��������9�cZ��~���{p4�Sh�?s������2R���� a����˷�s�9������ڭwWnخ� "9|=�<�iJ�G�����Ź�������ů��v�{�w��`{�h7m%��=���6�P9o��@D ��=�\8�F���uf� �����ǃ�{�1�����mnq���7�i�)��A����{����߽��r�����IR����0�
°�,O~���Ĝ��2�s��u���w����?�� 쳰�����B��!���>�{������w���7�BФ+G����X߾��^l2^%�j������,���4�w���嫎5p��0x���r�J
������Sڎ������HN����/w��Y�� ��eM~��jgJ��
!������8$�,=��6�8�s��ɜ���Xm�_k�h=�����v�޷�CI'�a����9�J2�����q �8��}��{��wI��!ia��}�C�os�֜>�r�7�'��=�N VQ���W��ލ�i �}{��}��3:~��=�c��0�
°�,O��{Gr!Y,eg���z>�~�"�淡>����G�ܝ���Y煓�!b��sx�:�OLq���>mx�&�MK{�Ċ�� ̃#����p��R�?w����-�+X���/D @A��`.���>�J���3�{���J�2T*��{G�J��w��ss8�m��Cl80�/������� A����؏��89����o,�8�R
�}�l��
Ԃ��������ciW��V�q�ޡ� �O�拌�Kq����p*m'�s����ed���__�ލ�i
$�T��׳�wG>��ߡ���(¤�����q �r��e~���I�� @�=�����4*hB@� �/�퀹Y�0�n}����@;3�6�yHV�
��}��SbJD��7����%}���_D)������v��_w��k�2��g�AdB�{���=���������}��fуȽGs۔0�M_��2��XrӍW�<� ��I�=*�~��8����'�m��3���s��� ��=ރ�$�
���چ�;�|򙾷[�@�T���vq�R
A~�oz������Xw��<`We�|�~ӯ�懦V�\_o+���V����J)����^u�u�"����jx�.p\7�������$pd���^��ލ�M!bJ�X@߳~^G�>�9�N*����#�O}����9��ed������M��#��2f��Q*&��I8D|�����>�<%>��w�X���Mepmr����^0+c���e6 T��~���0����|o�����QL��{G�|$�)�w����\\g6�n��W������V�;�G#8���� A s����?<�靪W5��A`~�,k���P75H4�(���g�_�!|�3�-L��
�*_ȩ����sG��~�7�\�Ӿ�hd������5(m%B�+
s�{�Ì80�( {���m'5�:���5w�a�ᕒ�������i��߱�q��\`�pݜ@����s�t0,jB������m ��پe��yuOk�4��
���^���*T
ʞ�{�C���YFJ�����mD������y��ɯ�Do�'�=5��E(CM�D~n"�?>�N��+��So�*����uN�^�{f�7�����u�o.n�>uKʣ!�������_���TkM����i���ɝ1خ;2���y�Hz�}��(��n潍�ڝLl���xV�L��n�t�V�X�{l�6���<�Z���:�����ͭې���6�pۑ�n�%�8�}�S�������&��������-����Hb]vů.{qonOu���[<�kg��4�p��㝇��m�;�:�J�۰�tnܓ���I���=�pN⋱�řt83�N���ų�H���lt�b�˛������隹�s\����¿]{����B��V������d�ʐP)�{��Ă�̯��~:���X���ځ�T�JB���jx����kgO�s�Ḹ��q8��罣� ���~��ʷ9�6����2iT(���>�nH,80�(���{Gr!Y++'.}���?3њ����Y @r�S5TDT�9�*Ұ�?s�������_ B�}$A���b:���d~�t�� ��߻�ڇ8�P�K;�~���}�>G{�j*��I�������0���r=�)?#�������Gq��T
���߽��x�0#��������ˡ}S�iHVϾ�����^�����ѹ�mn1�6����4q9++%e ��+y/�4�O�&ǰ�|4f{��8Ã
*K�}�h�NVJʐW��oRm6��~w�o���<�O�1sV��v����;{a�b!3�7OT�6�WRXk�������)�e�M������a����G�
5!m���ѾR ��W��oP4�@��ξ>����� ��Ok���pd���
!��~��!ĕ�>��qs��9��r���a�aI��/�YD#���twj���f݈S�/k�uv��0߯��@�e�5��g�*;�����<Jw6���]=��'��s	\uc�D�j�}�E��鶁�GRI$�?0�����q���
s����8�Ĭ
��ﹽ@�� �xE���jENf��j��x�1Z�:x�ˌ7�'s|��N ��U��oP4�ĕ
$�5�w�����:��ߡ�� �o�~�������VU��7�6�@���o�q��s�E ��/���ԃo)����%�
Z���Ѵ�������B "����������ۮ�����_��;*C\�����g�����$1U5&������;m�!h5u�}��b�Wb��cԈ�ۙ��zh'	K����'cM&C 2ke�ļ\-aS�Hd�Vr�f�)�??y^��i�O��^$�+�Y��{h���X���_�G�L����X�!q Jim�A��jt.�9�$ֺ[c��'�]X'ľǩ||ʑ�+�$H���EEMTT�Pl�X�����"	U�*��|�wweܻ0���Ԑ�7���b��۷���|�	,7�'ᚼ������}�]�j�v�)^����������7<;���f���o����}y�{C{*�X��{�|<�s�t���;E���v\+|��^���s�� ��[5yr�7z���"�Uز����n`���.r��Co�'ӓ�[ނ�k�주�g7C𗵃��;�� ｎ�����|hJ��zdޙ �s�)�t�
��ʉ:�=�9����+)�{��h�l��doo#�������6�Ձ����w���K����״��s�n]�Ȝ��X��.��ݏ�J��F ��9	j����p���J�X�j�e��Y�;6y!ד��eOd�.���x�=J�řX��2 n�n粲uLk�0����ױw��p�_t{V�Qzh��jg�sI�+���(W���'��fˮ�����5q�V#��zx�fƊ��̚�Nz���^�I���s��o-��?n3�X����6G}t�-�.����UI�%���^˓C�{cǆ��*�n��La�z����S[xG]������=�v�[�ǋ���Piˏ� w����'N��݄����W��`�Q��;۠��=�x���o��t�W&��������p�\(�5_#%�R�wb^i�T�%��ö��-͋D�C&ҍ>�}�x�m�6����fgg��X��O
����,�`���5$��c�����}x.����-��o�!x~B-�vmK�[�ڢ�fqJ�;���Aqhfن�L1`a��)s����-Y�.�`I��Y�P�i3�[Y�mUW�S6Ȉ\�Ʉ�eţ!�UB����m��Qh,��(e�)R���J�J�QeV�m*��R��-��b��b0���ip�4�,1i�Qf�aqq�\Z�a��Y*a�h�Uh��f\��TÅ-�X�iRVTX(�+j+�6�dQ�b�3�c#X6�h����KV�P��iQ\ن8�IF4���*��D`�*T0�L!Tk�`���-�W��C&(eT��L��*#UZ�eIUh�+m�X�AV�T�,p�bʙ�&�R�H�V[mi2�E�)R�3mR\Xa�Tg{	��N���� ��1�R�a��c�T[h�7�8��0�&��
�Z�ڕ�Z�[V�mFT�+%AV��X�����	���C9��X���1�+*�m�E�,+3�de��$�9����
E߷�X>?v}��b%��S&f&�շzH�N�-#r���mY ���/o��Z������7��� ʷ���ki������cur��m�^+3�3�M��8��$�cH�}ͤ�7��ʚ?~~v�����Qr[6e�k \�2��sf9�q�C
i��l��~�o�[nM�w����Y �س�>$�_six��Dd�P�Gm+�ImcH;U	�����)���$�6�v��;\ �;�$��m I톶(`��IV�����{d�1$UQ�:�-� y��x�A���ѩ�{U]ٜ�XH1gZ$}��$ub.	��������](:S�^$�^jGĒ/w��H����څ��&$�I��'��-�,�'�inl`UJ��.*UR�yZ3���u�W�T\�����<������cq�?gy޹�}K����9u��
z(��$L1F "X�2f"i/w�� Hg%b���Y-��D[��D��Y��{�ꃧ���
-��&��0Ȯ�	u^Ĵ�mȽ����7��z�ƻF�\��{�ٙ	��4H*���m� ��ڮ����y·LC�X�y�"A�|��;�hς-��%�0g����{�]�gޝ=0a6����;U݂���nB��o9ʄ��$M	�0bd��x��$�F���
��Em����${��z��X�\B@�K��*A���j\�f@$��h�N��Y �>�kVѺ�d���w[���DQU3ST��.�U`��c��wWZ	��K�Ƃ$�wv,N5�#�J��7���3ޒ���´�/)�sm�i�$�s}/��tAj��QF���a�E��,��e��[���R�1�OHu����s��x������)5��j;I�˜�GnL;��΋P��6�K����p򼝶�͕�L���W��y�X�Ӂ�ɺa4�j�'�c����؛�^ncf��\y^;�m���'W��l>�vNk��쫱�ù��#�͓�m���]n�0��/m������kl��b�#���w,v���փ�F����85�nD9���ۈ�q�
7Y��!I��7l��V��Y��ez�����.�=���Ɍ�{�۾��wJ;M_ޤ�$	'�g]س�I����Ȱ�V��� �ww�>�0j��$�P�l�Ƽ��*RA�)Y��-�|H'�:�|H�Ԉ�1��^2]�2j}Rb�����|O�y�� ��+uij�w����wb�C��mD,ۤA
jb�A$uo]����:0j��$�7y~�O���@���մ�;�_
"�2ҿTw���B��S6��]�#�IǼ��;v����hGm�#^g$A�筤f2�u޽�0�
��H#eͺ�i�6c7�*t#�)�[q;d���۟��g4��s��-��x�Y���w3�$�O���.�Ķ�9LM�g�-}��D-��j=��G)RHM^���h�W�O:�v@x��h0)͗�l�^�Fu�d�;[�ȯI�ۓ_[��(5@�Wzr�˥#�R�XMV�9�#�[�x����� ��_g�f|�� ?���7Vm�C���x,ȪB�B��Ӹ�@��ݠI ΚM��&kn甭�	��O��i3��ԚCl��R`��h�o�_�J��ϫ�Gvw$H��w.���=т�>M�Kč۠rjD��52b&��'Đ���q4+���r*I����|K��'Ă;���^s��ͽ���q��f����.ݞ�g<�\rq�͆*�YT��g�yzy��&Xi�������K��J�='�h�s���I'Ǻ��]�qnA�����	�� N�A��5S5B �9�XX��V������GĒ�H	#������Ф���u��@�JR"���n�6��P�n��!D���Y�c�Z��3Z:�i�u�|{~�q���G�9���yn�*���ٽ�..�y�(����8�{�����ӣ���{�� HLcsǅ��lؤw]ݐ^�*�I�j��7�������"R���`3=�׉�wVH%�cB �\>4��-&�!���S �ULED�DC��������j�!n��'�}��$��wv	!�cC)�Ř����?�lɺM;��^�yƃ�c�ll8d��jm��-v���Pn���[�~���l���8���4���w`�@��i��Z��(������ز�ș�Bj�e �ؑ2)TU����I�;����!�cH���N�E#���{>�t\�Fjb*�LA�C��d�1���Y��Bs�T'y�	 �{Wb���1��ǳ@��G	d��_n���+`��U ���lX>%�g$H$s�kM�,��q��Ѽ�`xbC�ϭ���{�lY�!l�t�B�%���T���\]u�췳���F�4�vr�x_����o=�8b�x�礐$�w��ji�׶�1F(@3QM��q�@#���<���>��@v�� �9�h"G<摊Ȼ�?��g���ߴ(\����/�غ���n8������;�6�H��t���u������k'S�/���v,���g$A�sBs.��%�r�k\��U��1����F�L�T�T��1a�4�;e;8�t�ȕw��f�	���8�_��_���I�3&��D�@�]��1�;@�|q��C�͙7�N�� A�Y�x��9��d �g��-�����yϲ�P� �g/"	�$=�iA��]s:�l�Ϥ�W���ʁ.f&A�114����@��Wv̻�4�q��n�� ���$�;�X����5Q8H�h��fB�m���g%qU:^���]�=��T��?=�a+a���TN�oO��v���0���/}���HH@��^ˋ�9���521��B�(qU���nq�83����=)��H-���6 �O��`V�uk�4�1��|��|�X����9�kH�L�����/Zu��ݙ��]�/G5��-�� �{sc���5����C�⎑�7ێ�S��G�ugu����lr^�G �j��.Vƞ�s���W��G� ܼچ�T��ػs��@(�f�͇Wrp%;]S��7��2��E����)�uP�c��Rq�6I�����	� �TMA5w� ����D�{�U��)G,Uƃw����z�]VpmDP�JhZ�a�����|>��e�|<8eUUMk�I�#֑;�]��a<�;�Q{n��μ9[-4
@�}m��I ��Y ��!p]Sr�a k�i�|Gu+�����55fR�v�vL"����(�o�x�A>-ҫ'ǳ1����� ����N�A�ȩRb�h�6C��d�V�5�Y��Lu�$Rw�	 ��W`�^f4�Ĉ�?L�}���M���)����M�ZX�=�n$��<;&��A\ƹ�n�5���w���W��,�:�Myx��V,�Ay��x�)T������g�f ?_���=����D��wS�@5�s������!}Y{V@����L��N�aI������y��������;��J�toX餬���v��< �����|��U��~�ϒ'�u�Q�3â�u}���g��""*� �J@�U�d��gZ� �1��8�Z$�WB�w����2�њ��"5޴�:��R��ս�,�Iw���G5�ogu�d���˻ l�fMME�:8�v/F��z_@#n��	w٩�M����2rbڞ9����Q2Um�.n3�f�mS�x�ֲ��b�:���rKZ�s~�C�dT��0b�	/�N�`Y����$|�m �註�[zU�b��}� Lb(��4"bd���HSO$�t�F�*ݲH'oq�I>m�K��0}_�wg�u��h &! �l`����$���$��h���#���W�
)N�'�n�!ϑvء�3=����/ֈk"�Ei���!:#k�O)ӊW`�cf+uNY���=�m:��y��O� }�=H�t���(�ET��H��Cq�gf��k�C=V�@���ր$F����q%LR�FR}&_���6IX�=�o�` `��X�Ȭ������q+sD���O�޼������e��[�h" ��Tj���q�c��;g��q�כ^l��щݪ�:��5l���~�	f LɊ�Fe����'�5��I$o^P�g;̋���k}h�dӉ5BjH��B��-mX+y�v�m5�� H�o�'���.����t�_c��Z��(�uD�ĉPi*��/	v��~��Pщ�VaW���]���!�|��};s7�l�2�c`6�wF����.�Z��Gjʲ|Ofc^V��Nk5�}O���e��1]U�?X�ʅ���,r�u�@���w��=����U���˾�0{IM��?W�b9��S*U���� ��v�q�]���x}��:��!�9Ƣ��������,Y ��3�f�V���	ʼ�I>!��$=�i�Y��Y���i6T�S���q��c\GKaz���vm����^M�XO�
kS��-�Ze�Ix��}�2�ו`OncH���V���z�I	=��Y%�&G	1&f��_-D���P���ܥ�ء�� �ګ$���/ℾ���9!���|zh-�40�1��{�7���o�#���$	�w��#6��>/V;(�sF�ə$Ы�W|ө�Ŷ�IR}~��|Jk^$ټ�vovqN3�E�V/j0ѓBhĚ�`��� ����e�030D�\���$IU�	�b�KĞ��h�ZȪ鎱��k��PBt0ͫ�i���l�>*�k�^QA���<	{�8�=�e3}Ԍzp��B<��\�X��!�p�7`&���<�@�D\O/g:�z������Rm�H���þ¸�z;&��������1���v皚���f��Q�H����p� %�|e�ȉ,CL��� �pj�$����O�����7#�K ��0p?�ȣ�É~�����-�;^��H$����2dh���Y9�)����n@�� ��1��G���V=��
|�^�7�4h�����ts���h�����a��{\./w�L,�_y_`O�=y��;�C����,'9y��3}����a���[x2}��/��5�|���W:�#�vG��5��B�ؖ_��*���x��B��,0nX��{�m�7�R��������%E�曗��K̀n���)��B�:qh^��yxf���<���ދ�3ڒz�����fһE]�^԰Z���z���ʏJ�K�g���%�`�#Һ�Z������h��5�����ǎx)=������l��Qx������o�;�ֺ}��Ѿr��o1�^�d� �٩F�+�/CS�.�,��4_�;�e��k�1ߴпz�j;t>Ve������G�Iz{Ӈ�Y�:5�S[O�a:q�8��ז��Par�G�$�������*��9�R!؇��x"����ީ��=�t�:�~<�����w]z�wSyQ~ߊ��n4����7����5�%~|�^�S�]���=��9ۓ!^��\G��c��
 )�ֱ[dV��a����0�Jb��E��ҵ����J�^]���Kn%��*>���iP*1
�"��m���P���(�V�p������0-Kh,
�ʥ1H���������p�fQ8;��ڞ�Cø9;�ÌB�\�嶆p[0���-�.ReQEq��m�#K�Ua�ŔI�V9�j������Ì�Z�E*AE�-b%ŅC�El��&�9��L���B�R����J�"��0-i��L��Q�&\+�
��e�a�aŢf�$U�-eKZ6PF��(�fVb�ƴ�,�+1�m��\U��԰p�P+p���1���<���H�r݀�x��*����1�i*
��b�*TH��(��h �[ �kl��-�bZUKj�v �[�[=�g�=�m��TciUij-���.:��`ˌ�7c����v���!��J%7>[����n�hh���9kkn�A;��oZWby�n �rg�ʚ�v͎���ne,�vw.^�{I�$�vtq��N�7uκ���Ih{n���GoW��N����8�g�6ҁ�#��A�j�X݃��7nk[i���]���OU��v�ei�}v���n9��n|g��k��wz];n�� C���@�����qk^��]9v��n�[5ӻq@Z�B�q�㬄���0v��mu<E���ٌ��V����r�\�c�g��y_��7�=b�˜��Z��>��u��B���l��Q���ٶvݵp�;q���K��U��y��p!�'[0I�F��n۰Sر�0۷�.��R��s����j�s�\�]�0v��c�JS��mÞݒm���ITu�]���rQ=W)����'gn3sˮ��g��;:��wb���_l�3��{��-۴��L=�)�,Ꮌm�凮�
ݍ<�Y��/L%�n�9��pe.lʛr�)��ri5;���0�ACx�]lRn��z��ݗL��cy��0�,�=�r�`�G�������O�=�O%p������Wiۻm�jW��ݎ�\F�N��S4���I��J붷�;���׋6z^.�y6q��[�UA��ؼ���hM����'8��P�`�K˶�'=b���y��ԋp������|"�ז��xA�K�f(�`���c]d�5�����,w�:��
FqyݺS��l��2�E=A��ιȏ����m�^B�5MսrX3m
���crj�.��>�.�vu�!{��3S����ل�pN1�q`<mk��*/�Ws	N�3��C��㴡ݞ{q`�n�ۇae���q�Ld#���#��PWB=`��0�>�����۫�k[���l�Ÿ�sO`����<����������w���;|�:�e���ό���q�����N:z���i��{;�9�3�b�v#=V�MgZ��{���#���ݣGD�z�LGs��)c1Wc���\yι�����۝��.��mm�kŻ\k��X�p�Nԥ���U��x��e��G���9cYcZ��>��<gGh.�=��vX�rw%���rX0Sv�6�����ٹ�sН0V+n+�w�m��C�m�F9;rog��ݺ�z�l�iC�<�]�<f=�H�Wh���<Q�մ=[fy6;-���U���]q�'�a�ہ�&�=�������[Kgm������ ��W� �o4�U�]�MD��uf7ۿ�'O��_���i��%�|�^�*[lũ$�֊�庐$��h"&�;�`�2�5�
.N�L�bLM
�����8���A�YՕsXE�J��iT�'ć�����;4f�	3hQ�-d����ogĕIj@�F�m"	�֚�4�7�@'���R:f��3M
��Wm�	#�ڱZ�t��b��I"�� ��c旉�=�q�ٲ�����9�쨇�,H6�Y�3�,��&J�Qw(���k�س���(�ݥ������U�F��rZ��������*�v��e���D��ݠH�C5���e�K��+γ�voX�>�<���	����{w��?�T_���m�]�|~����_��֜InTh�|��;W�����T���+��BM�o��b��{���ǯ�޳�R��xp]ݓڱN񖊪�����)M��x�.���$�7"E\�G5��|�"N��u�yx��b��EZ �]�o.���[�ėiu�A>%õ7��Xѩ��UF��r��9x��H�P6j�ȓ1F��2Z�|F�Ƽ�x{����ĉ ��ڿP$�,i(����rv�ٽ���m$������Z�;�u�ָ�QO]=��En�!�����c??>�?M@n�&M
�Wz�'Ğ5��Gă���3���e ���v�$��WG�Na�j�fhI�Rl��i�y���v]��u��	�lO��4�C�@Wm�Fm������uD�H��(�Qѷ�pA{y�)�0gEӺ��*W+��7d^�{��0���ݯ=�����D(99>'�wDD�y��\�Xm�:5�wn���MI}������y�|H:k��^!���;�6D��LE
�Bm�]r&4����M����$�y�ky�i ��S�F�GZ�G$���b"%��%Ƀ�{�&��l��{���n��'�;�ax���A�P�(�5fav��,f�E����`SX��jx-�H��`a��vv��%"q�C���sM�iK[��1=���z"{©�ۻ�����-���@8�H��#���` 8�q��*܍� �����H��r ��Y�!L�O���}��O$��jM�c���$�����s"���L�껮�'���d��9�	�Ω�5�Y,,jL}9����o��Ox��������	>�h�C^�n�Pt��`:�v����_�2�W�Lv�ק��ǻ�,Gf���5���Hp�"����2^gh�8:\�Fê4x�{W"uG������;�	��6D��LT��Bm�׈"$��z7�T��wy9D�%j�A#��K�'�^īޒ3��D�Yγ�ׄN�>\v���%5�2gt�&�{@���	Ɓ}}�,�	I��M_���� kv���jl����t��7n�H'���� �X�0|�D�N7�hѿv�f��s��[��۰A��ց'�P8:%&�Ƴ�ٿt�X9�|��/"�Zw�#�=��{�R�N�u#"^��O��kA�']�9��$�M@�lt�ns�lUtMF�Wfe�A$���l��d�F_���s����"s�gV��,�52�l�`�_���q�麡n�H5��i0�9"A �����q��=�ޕ�)�UA�O�M�A�#i��#���Y���!~�k�5��{ƚ��L7K���x����M�ws�1�c����BF�י�rܳ.K�hݭˎWq'd��;nB�_5����;nŮ�vu�7n�/��T���f9��V�
���������螗�\�Ƿg�ۚڅX�+�n1n,=fM��i�Gf��;<J;��Ck��y��M=<����eL+�ō�Ż�mG�.�[fWn 1�N���y8��Ϲ�ڣv+��V �D$m�;Z�Ě5e�lY��O8�������67��,F��-�A�q�6㰭o����A����Ͼ�l� ��`�@����芽��2c�V�$�=�b�co蕨&j(���pWz�ֲ�-��5v� I ��ܛ�$�yvH�SU@F!��of�`�a�R'�4h߮׵�X�	�=�ճk�X�ix� �W@`/�w ���IaKğ�޾�}�N `���#���|v�sn��צ��v�nh���)�`ѿt��/�z��&0��bga�L�Ud�}�Ջ%�kH����˃Bo�z_��jÓ���v���������|݅���W;�+�ꙡU5�e�3Q^1F*$T���r쐵���OgkH�-�Or͂+�݃�}������Ń55"jM	�{/I=���M	C��}���w�[�j���/>��hC٭�W���@�Q3�%���պ�����購z��~�B
����.jo��+�I/�#��
#���g[�$ �~����O�A7�Y}��=�3QET�X���`��[`׈�aV����yv�����h��m��Yڊ�ffUR�0�y��B�Weu� &���  �F{Z�P��wT͗sݓgvv��Sm��oԨ��fJP�[�p��Y��M��od��tW筰� gkH($���u%�͢��vܗ���MKmn}c$ůoY��nݮۙ�K���1��R @M ���B)��,h�7�5��f@@|7�m0 �y�@�W��̭��u��y�ﵿ���ڂ��((�S�U��m�{�=���9>�mn�
	� �֬�C��J	/����'}}�^�@.���UR��U�4-��q�.��l���Pwe��F�2�rR"��8�n9[97|��u����c���RC��A�ѷ�x�[��D#��8�J��3t'��k^z#��ߵ���!~�y�eF�蚈L2[ot������^����� d�޶��g���� vs}v�ѓW����{��a���QS32J�RƐ.y�6|��λ�)EU�9�g��C��m��g�d3������6��g���6��q]���$ِ�����>U4�p!����sl<���?n�]�)n��`���6A���Gdu^Lzˆ`�����g��׷�HM1�,hd�|��BF�y�3��f7�~L� ��� Y�Ϳ��z�k��.�hk<�7��~��٢��RPEJ�Hv�I����Ͷ��/�n��f�����<�d	���@z�@MUJ����N���z˿s���D*�˷��_6� =��L�~bne�L��MG�ْ�zyO=�e��*~���֛��5U�����	l��-Cy&���ǔ��
}Ֆ���}&�9˷6~�����"o� _�?{蛀�**
��m���` ,��w
g�ySҧ��}�|��z� g�[LS���3.����d�
��3q�;v��vWzI�r��m�l��L�\n+���QQ�&I��ۨډ��$�R��|s9������ (�v�`����nf��́ ����*�ԩ
P���6*�����qiX��ucUW�ؐ����ݭ� ����Z�Og�G{oL(����L��߷E�I�Nz�m�@�T��������3ϛ �{��Y�55H�f(*U���۔{iN[2��Wf[��� >���q .{���2�������m�������51U��������m���bq6��z��Ͱ���� �!s�[f{3i���[��Z�S^�l.�r+�op�h�
��p�p�]��O�s֬�n/f;�ays}�����:�(�##$t���&���=rj~����}�竴y5��֞=n�Ɗv ����1�PA��6d��.�O����n�����F�����2=y������4f5拞�p���{=Wn��v�<U�6��';>4pk�M!m��<27ݗ�q<��7Z3�\�9ɷ�Ǚ��kHө��d�)�|xۗW=�����8;�9�\�"m�{y�e�O`� ��M�^��{]fcc�4D��lvyF��ٹ�)=S�0/V�������emѦ�?�?q�B��[a�D	G=�]�I��X�SV�yWW[�� �[���z���a0�E0�Bo��'��$��~�c�������;h¿w��0�Q?v�*�گj@|�kީ��I@�s�p�!^�ͳ��ە��b��� >}�� �!_���`�皉	x�	62�����y�ۏ�}t���ݻw�>��;i �n�]ܨ߇���ȑ���?B~��M&	i&XȐ���v��ͻ������o���Y�m �B�o�L�ۜ�A�'/��~�/�O'qH �@� z�����v�g8�ݹ4����n �w �۳������{l̦�ԚLOPI"��H����i0˕����s�.|	��i� �y��������f��(�v���m0AZ�f/�z}��D|PՇ ��:��X1���ᴹ�wS�|Ũc������"�G`���ǆ�5k� !��>��<:ڼ�jED�}l�����w�b"�ڮ"!�������EWE��˿&)L8�TTD�@�����l@nu�� :�N��5��w�/�~�;�`.����,��T�
%TTB(p�o��s�[}z���z�b���o�M� �9� 79�EWzz��Mw{/b�^�m�k�j$&�R��UQ-���I�I�Nz��A��{'%D[[�B+���h����|dnsvN�O�Z��]�������K���k����o,)6lఽ�"�m�^����mT/l�>�[%�LK�7�.��� �=�� #s��*u*U������Ͳ 3^����`!����1��ۙ��ޜ^ �7J���~ ��[ �279���)�&D½�mEÆ:ow Q�{<f���_������ �Ow�3H����|��/�_/gD���������2�k�1��.XV�o��̟o(V���w�3��l�q����o+�pu�f�e�@8q�C�^��
�پ޾S^# 7v�8�}��;��P��Rv��*�9���j����������Dy�9D�F�I�-���3�P�{���G;h����&	ͻ�[�uHub�$/*��V��$�z�q�;�K�����W���7�{x}x{�|gf�rQ�����ƻ~]��^�h�÷2/Hm6�w�z�����џp�qYv�P�>��nq�D�O]���P�N�����{�u�-g;���3�j�y��}r.�;l�W�UWۃ|P~���m��j���~�[�ٸ�_�yo>�>��s��Y5"�+���>��H'<���lٵ��nM�;���1��xDÓ���������9�z��\0j��M�~3�#�	t�_4�ʟ����������ߪ�M���zC[0<������,�r�xy�9�����g���L�T��{1j�n�]^�+.ҵ�wt�i_�k��N=	����%͞s=s�z���o�F_�f���j�a	�aɽ�؝ѯL-܇�ћ6^�aj�lsw���ޓh��@�Y3h'/c�1Z#B_	�b"�=����	c����Q;=9�66���b%��k���v�gM����o.n_ܾ�ن�T1^�V4>�B͗L�{�oc��/�`{Q�'�E�����'�;ު�����ڂU*o�V�L��/��һE������Z��2ڢ�ե���m�imU�1"5���iR*��*,QQmmdU�(�J�eE��L5���[m"0���J%j�b"��mk,�UR�J�aD���0�U����-��Ԫ#Rձ�������b�QQb��(�J����V��!klB��.0aC�iJ,mn0bb�V��*���1`�EV�Zb�-L`�j����UA6�Q[�TX��\5TEA�UE�
�.-E��1��e��Q-��Z*V���*)Ym�hV��k
F"�(�G�,X�
X֭�-�V�+X��aT����JR��h0���V��F���5Z1�����E�(�()R�E�U�����
�*�UQ���Z�-�����EQEV*�-h(1�)iX�*�*\4�V�@�vu�;�븆����a�S#U�f�T��'�iVkY��5 |ﭰ@ ���:` �}��͢_vDtD	��I	59Ka_�M~%�}�f�@�7��ޅz:nN�Z�{��y���@#cw��dD��;��̻6;;�|������a���mW<84⵫���]�#�֟����|�]��s������&���`��0A����`�E����.�y�Ӻ���3 ��o�݇Vy�"h&�K��HI+碻�w�}�{�Q���":;޺h >=󸈍��W���Br%}�=�'��Xx�L&��hث�P��6 �ʧ�$�m�v���� ���6�>�s�6̡��'��_�kt{������r��|b@�޻+� ��i�IZ�a+�rם��g��{��^��N�l��{�{{V�Y�g-�5l͜I��ʸRrmMT� ��m�sNZWv"!oA_�ľ�n�31�>-dDj��%5�0]�Zl�����ټ�&�x�.�k}�M>v�� �;Ͳ�s�1�_>_7�~�����Y�Z�m�NS��-��nkz�]��S�`wiN�n:Ύ�g�����u�eLMT|UM����6� 3|�` {�fz#j��`���v�����DD��᭷��R���MQ-�]nvb�����P�W��� ���󸆀���f �j;��S�q;�f�ۘ"j&"f��TE��W��q���� �}oed��^� ���" [���π[\.�C/)���^�O�>�~/l��P �����v�y�@|B��=�1@�R���������3T+�&�n�����` {��p�ކ(���_�]�0���1  ����m�_�x ���&㳐޵��l[�Զe�(�3^�h����A���V�~@�AF_f�gf��wDC`�i���:?��wn�~��Խ��s�Uq��ơ��l=��p�c������r��g���<=���V�.���糭�&d�7�3��"�n$i���#۶����,�5�;Rb�O\�W�����3��4F�j��:�j�7nC Q�:���=�2s��:X�<[�$��Z��:��j�j�=���R�t�^���۱�8w�{ni�\�7'�tFБ�]���cT�qm�0������T25�&�lg]�G[��]m��[�gpnq~����;�OY�c*dB�~��7��x����v�2(�w;Yi�u�� ����/�*RD���>*��v�i�����(�I�[~�M� |������6�d��v�4��^�L>���U**aL��f�� -��l�G�w�~���>��񼸍w����!{s[���Y��<)��4$�q�_����Ӟ�\tDyc�<�`|=��l ���|��ن{~������z�e�E�fh�T:k�mkm0�"<֛ן`͡=�DCO�ݙ����2�N�3!ϧ����t�� e�00 %��>y�]ͣni��:�3���2�:��i����:��~����R"����w��q��o�� �vî��T�a[��)�ݙ�|/n��<)5UJ�T��
��ٸ�n1|��]��^���ûB;��]3*��N�%�w5��[�5t�/�y�g�>=ĺgص�6�������@e�>r�]�MG�_]����}����|�� _�y����]���x���@lߡmL��)*��lU�[L�c�i��D[tMﱲ:�=�H ��o�@ ��L;�QT���S2ٴ��7vl�/7{�}` ^�v�  Q�ޛ	 ���wp�*@��1�_�'5Γ�'>ްKxZx�4$�q���	�ݏɅY
n�=������d�wcx�@��,��]D�(�����c���E��b���f�3�u�.�:�9������U5Dғk��ͶD���b������#֢gg�t^�xH^��� @
�5�z��U5J��R퓽���+���sK{���Qy�퀀���3#ѻ{��n�5/޶�)�F�T�%5$S"��&π��y��&,���N'c&��P��<^_ݣ�1��IB���}/k�Ob����r���j�a�"��t��M�k�5(ܦ:���>�qw8q`O�`��ߺ�v� }�{z�����絹���}���u[F/��Z�m�q�>�uzO:��a:
}��b ��٘ ��"_6va'@��� ���b���MLʹk��ϰ>�[��q��m�P��M{� ^�>�π ^��f,B������W�UFj(�BhЙ�X{j-v��g�����w��C����'g��[)�h=U�������"��ҩ���]�m�|��� �ۺ�tN��o�{..9���L��n���n2(��UEPU)��������܊��t�Z����؀�|�F ���6�k=Z\F�g<��]���\{�Dڪ��ET�d�n�,"ݾ��"�f��Z���8���`a';�O������K� �2�����ϻ����W���@ ?o}>�  �;w���\�X�Ʈ|���q���&�����M���0�v����s��q��3d�V{�%�X���.#�5���j���ߡ {����ğ'�/� ���ra������,y��������P��_ �ۍ� -�kl�.�۸��z&^f��;����pz㵦᳴����_ۇ5ۈu�C��#z������O���������fW����;3 �o�m�@$�6���u9�)��{f�"=u��pߢj*M	�Ro}+s�Ј�����)����}�� �;ݮ�u涙�+]��������$����a'��9^�� �n�� \oz�Jz��NNw�[d�ך�L����SU4
J��h���{i��a��Te� �u��| ��;h�ϳ]�̨��"з{[���W��TJ&&��0[����>��x�;�-g"�#� ����C@|-��� {w�2 �����(�rK^.�����y����B�g�y �v׹�/_(�Q;���t�n�x��p?���qu؃��,�����{����ſ(�e�"�<i�
|�z�x1�`�m���F�N�=�vઞ)f�ˇ-���{nq�sַPk�b�y��=�#������*@�so%˷I����t[k]�#01�m�|��I`{<𔹞y�%��l|��V-���:�6�ic��'e�b�l����!�x^����<I6�*ۃ������"�q�bg��{��8�M�X�7f�m��QJ7U�(�`݌�0;�v�X�W1�g��>��O���T��UU�����"/5������Ȋ���5��N�$��x�
#�ـ�m�4���}{���ȳZێt'���eWg��z�n�n�w�O���V\�Y�	��L &YiM*�o�U�۸��gwc� o&TJ=w���]V�$Yy�i�|�~��;�>���[ģ��#����H�漑1���f�ov�%=O?�	8q{��h����x2�n�=��ŀ����0w~����7��D׼�	{��3����[Y`�郶���o�HQ�Ǝ"�x���;8�l�Wu������wP��͵ݫn�
.o��؈�D��D�����v�{{%��@x��	�=9�m�S��2 >����z�=H�Tȉ*��vkX |�K.׍�fJ���d�蜾��1����J���'>0���2�tP"U��3�֖�k��ri_qn���-7���"D��<j�����'�� @w~�������d B�|�i]+��0K��������D��u>�b�"#cw�� >w>���k��booff ��vf���H &Y<O0��޹��{ �7;q��=��m �B��9%lm���yޘ��U~����X�PUDUER�tж��@ Wٯ���/�2f�w>�*"��fdF|�H[�悂L�jJ.�^���жvwQT(������� ��r'"� <��؎SvI��l1�؊�Ki���z�0�o�[S~�U��8Ā��[`_g���S�^͘˘��Dr����3���;��T�#U��PS�q��VE���p�
=<�� {��m ¾�6�	�3&�io����{��0�+f&!UH�*�b��m��|	�kI���W���ϝ9��9P7�k�|���9+��i��O��f����y�oD��q��;-�����:��po"	��ޝ���ڙ�����$�k�w�@�����O�y�4�/�DD�MD�D��O��x�m�O�VyϨ Oo�� C��l�^����g�MxaT�,M޶�.�� ��SR�U0��ͻ�wv<�����!x�u<v� ��<��L��33�m�K�붎��)�U��t6��aD��Ӝu�v�/f���=s��n� ���Ϲr�
T���L��
s��	 	�m�C۽����}h�\呂Ó�颱遖q��<i��J���` ���ϊ\�/S C���n�fb =>h��1y+�9��}�8Dj��*�LMAL�W���7���g�#^m�6wq[Y/n�� >�O��d=��� �uӱ$*(Q55�.y�am:3t}����H?cl�>�wffD.���ʷڈȚ�S��ݻ~��1�~ ���ߟ�Lvl2in��Y��#�e�ʱ�p�8+�;��b������w6�Ev����%���{[I���Q�!U33QE��?����"{}m2˝�y�E�F�s����|;|�6h��m��I�5�K �����Ɇ��u���iJc[v�h�ןIۖ��</����~�5Z�Щ<��i(�7�A$��ڭ �3�G���n&n��" ��ff$���2�%<o���$$�d���g��ym�@��ٙ� ,�󸆂�<o���f��G{G�4����<-�.}�p��Yۖ�dA��o�U.�W� owff$ �n6�*mS1SH��E1�]���qq��{�F�W����(��v�@!u�4E�Oz�E�e��vlc*� K�A�L�'·��d@-�I��z�̉�u@*�~�� 27��DD.����#؜��%�%������x�O�l�K��]�x&W�%�G,�+��P􃡛B>q`OT�w��݆��x�ͤ��7P�����}q���������֯���wP�Y�Zz=S�w�h�xr�3�u�{�lh�n�����ؽ���w=Vˁn7��'��%1��w=��W ��E1�Of�y� �o���xSc�~ǋ�}�'ws�}_wnn{�+)~��*Hڛ�H���뛣��5�	�o{�. �o�#��&��𣀆���Eb���w'��z�F�����Jw&wy r�<6f��A��/'0װ�O}�k�,]��ͣ̀g����/5�چzX�<�;Ln��|���K��������0d��L䳳֧�������_bҳT���aɸ��D{õ�;9�}u��{�ܾ����O�t����U�ɖO%#�Z<��%�]����G[��@i�輯M�%�Nn:�'za l}�˭z�wΡg�	��(��R��4e�M�Ӵi���sDo��m���`��^���a�;�w<o:P` �w���x~e���B@=�c�;w�vm������h���j0�{ �ut����Dj
f�FB،�<���s�s_{�ZC'���כ���1�<f��$��d�Ǘ=)�CJ��h9眯=�[�r��|�R5I��8�(~S�K���^t��n�	(�)cՔd��}쐏,�o����{�0Ipw�c%������w�A�� ���������ctV����X�U�
()P��ڍJ.,�8�EA��"�ѶX��XU��J�YU��U-�
թ[U+F�V�2���Yib(�H���+F�X�+X��Z��	b�*��EE��!l�[K��ZTEb6�iJ��Ԫ1EEX�Z��E*[V��TF�"֍��H��"��)�U�j�U��TjQTdEV"��V �m
�C��#DXڵ"�V�b��b��[c[DQh)Am*1,��Q��"ֵ����UE���ؠ��-�F��*�FJ�mU�a*"�a�-"���[(��TT��bDDPm��J��10�+%��"B�1e\Ym�ҭTb�*�jիF���H�KB֊VĭEF�[kª�(*���*�^���k�W�����w�ln����7�!�;���X��="�z�p^w��m�SAt�=�C�	�v瀍�z����[�g��8U�0u��9���T�¡v�v;ͦ���J����6��;��:��n�J���o�㴌�5������'���llw%b5��u�;�*��*4�"�5��֩�ȑn�G�ٟCή��.��Ò�р|�tvy[^��;l'j�Ai��ڽ�=��m��>3�u�Ms���G���p/1�m���/��y���t��rpC3+x�!�����cZzP٣s��,x�7Y�]����&z����k38����7B�g���;�OK��ݽ��:�#�y�+nN֭v�wt;s�'ӫ��[���c�k�X����-NQ��t]�;d�
��:gc��GS�m�f����s���ɯnqٱ���m��vx�,]�{=��7 �8�����A��m�z���N��\v��p��\�vzK�x�Hk���E��6��ݽ�P���r󳹥*�箪����Y����K�OZ��n���n�ǹj��N췊;�l�Kq�x���:��9D�n�	�t��X��;GU�۫���&C�����a;ud;�����|�^|r�y�;F�a�1\䧮��91�!^�燣!�;-�7;k�L�p�tjz'�s�'hO&��nϕ��;��u�>����A����@�m�V�c������ j�|��g�]D�xyR0�����f����u:y(�>N���v�ۜYzQ�"�a���<v���m�n�h��qI;b�] kl=qk����ŉ����l�m����n��[�t6:V��E�9��#��^����Pc�x�l��A��\m`�mvzcmu��/mOHfMg�w+>nk�ل��i�	�,���M�нJ��;v�)�{�.����n}f��v��:���Ib�cH�{upS��A�]ۥ��r[��y];q8�4�^��q�kg�]WMc�E������1�����;��a�O;ۯ1���nÝ��q=ru��=��'N�c�"�ix�.�����nlb���Y����v1��c��8�;b�v�Hh�Tu�]��]�:�l�����h�3A��譎������0G8[(�8ݻ���s�ɖy^�]��8d�U\� �4�=�\m����r��m�{n7k���m�c�Nt�3TM��i0��q۶cdQf��ݵu��G>�j�=���3A,S���?�� I�p�Ia���5����##u۰A%o��AH���L޼̈$�mZ����bU�QBhT�^���j �B��N'Y�8k˶�a���D.��l��7�w��Î���N]��\F'����Q���$����M�Fs���l�����pD��4�I9��OЛ�75����<	�6�_��s[�J}��@�Y�BI�~v� �����_��9�=���ܵ�����	%QLhg�v� 7���������q����}gy�` 'KU��#���f��8j؈j�s�|w�ڮU�� ���N��U���rه�#gc��9�x���J��*� (aO�-1�a���VB�z� @}��Ȅ��z͑*��9ڗ��&=յeuޠL�	�)TP���w��DϾ�C����ˇ��J��'�u]Yʵl��͈�Ь�E�7r�Y�ԛ�s����iV;f���ut^��g�~y������Yy��� ���o�>�~�ݙ�p�?`�^g�ξ�	��̘�A�Q4�a�T�Zl� ν� ��`�z�}��w��>�S���@���8���d�bd�%����(��=ѷ=���un?�b@m�7� ;�f7&�w����tD@5jH��eS��&���W���߉λ���m�"5E�n��m�f`!g^ތ��軁*���pn�$��L�`�ܛ�[]��na��{�`��p�u���������h$
TLʢ�����q��n1 g^�a4>��3���m�}���A]�Q�&��EE�&�I�f�8�b�j�Y�{[�	o_vf �|��N�Y7�BqU�
;;B����R���)TQq���!g^��0� ��Tro:�㼒��*�e�R��k>��V�����߽گ��^D0<�=+��NY���˓nڱI��	��pR2M��e{�O��x�Ϳ� ��7� �om�w��jh��"�d�D[O}[~�.�}f${�׉` �#:�Z�A$>��%Z�h��K��$�{����Q1�4@T�?����"�m�n�����r��Wc�~o ,��� ]��q]�5��ef�!T��F}��*���]լa'u�.g}��y࠻j�~K"�_!��&���&�o�{����$ Y�븈`}���Ao&=�V�w�����$�λ�]�Й,�2���<�>^z"�{���" >��� B���pb�YZ���w��q�F�`��,I����h��8Jͼi����]_�� �����"g_;�h.���u�"j�*�3J�Fͬ�gD�#�_ s�o�"޼VJ��׍�[�[��Dup8(��*_j��WG����#�o��e;�/9-B�U׾����a�]��ؾ�ʶc�A����a.�ɑs���� ^�����'1J&h&fJTC`����l@ �ټ�a�Z�LF�Ok�
��n��	v� {s����Ͻ�w�w�ʏ1��`(2���$���;K>��X�
Ի3*��L�S�[u���~~���ݠ� *v�n��L �x�b�۝٘����fϼV��hY���d .���`��sd��
U1J�����f` ���Y�&}��]�� uw��	o�ﻻ� b[��eH<�nBn�ha� �D̪)���i� �>�^�<�fUf�� ��Ͳ <�y����E
��B��)���gb):����f4����0�ߵN��N�t�����ݳ�=�����LҨ��e�?` }{m3�l猕�^�0>���l���π޾m�����I�G=�UǨ��&�\�A,���\��ȫ�eՉ�q�e^�����Sok|�{�u�,j�p�&aJ�8أvo���tN�L� B��*�W�i;Tg<�/X�|�:^��X�۫�ݹ�ܯ7O�f�;K��+��4�3�����6{xn-�3�	�m�,[��m�'O��{u��N�[ �KS���RXK�\[��"��κsΰ����n=��[�]�r��#�nM[<q�v���@�'�׮�s�nr�>�c[eۃ]��s��'�3�I6���덛O�V��\�ɫ����w9�4��<���%U7��y~�B%Q!%*#?���7 �{� ����owʕ�O"5�Z]�I]ɼ�WRd� �2hDT�^��[i�{s��u�*뻼s�o @!N{�d'���nC�[k������\�
�()R�4��Ew�ً�)�u����{�C�^�ٞ��罙�
s�m��Z�����2��4	�X�~�|�\���=�� I�;` =��͇U��w� 鷛���C^��A�1�:oۢ��@�ޑ���1�d�n7ّ�s����V�Q�7T�3��A��ܚ�$�4�g��G&�][�v�f���e��'��9I��[�A<O��a�}���'{� �{[��@j8�ۆ���gf` !Nn����W4�SQ3$���`��b�Y\������q8�uXTX�r���^q����y׼��ښ�������4��ʀ���ya�`N��g64N�G�t��z7����Wۋ��L �su�C�)�m�
���ggo�\$禴1p���ƽ��I8E}��q l�'z�ۿg� !Ov��> Wێ�/nh�4���R��]������V�=����u�����������Dg>��q7N��O�� ^y����+��)QS*�c�}�m��o�sq�̿lO����+�6�c�"4�a&Z3���u��������UK��a��v�um���P�;;[6�y�Gm��8�혨��JU
h����� �5ݰ �9�f`8˘�Ɍ{70���́ �����ncS%LW�4THٵ���y3y=��[�pz����  ��~u���o @���PI�Nb9w��/}&D�$�I�2 v��?�A�{�0 _V��m�-���6p�y=邥ס��S��}�)mwwf��U�W�Fk؛��7���ا+v��k5�Uk��a�Na�t�]w�˷�� �w��� ξ����p���	j1�_m�M~ܨs���;> 3�y� >׵��p�o�(�I?���N~����)�I4M*v��{�� .�m�Sz���s+րf>t� }�}ّ�߶�L�[�?1x��s2�@M"�J�P�'�4�k�Nֻn����[��힜&
#v�$\�����~ͻeD�k� ���N��޽�  �������:�&ʒ�����	��w�fDm�.�L�В&�נ;�K�  ��^G�3���!��%��n!� ��ci�$q����py�+�k3DҘ"�������� >��m0��y�2�uSk��^�_ Y׽�� ��ퟡ�ˡc���I�#g�X�¿��B�͞��V{, (�n;��Na������oS�P�*�m�7g�'�bΠf�t��,{ͣV����;�6@�,���O?y�Vy(�����b��b�Ȍ�]��Lc��ވ�[�b[��EED)�K�]:�� A�͹��z���^�H9}��� |.���d�fkta+ko�y���W���,�Q��P���{;�ɸ�\cI����sή;=*�%���e%~�^�Sƛh�Ys~��ݹ� �{���"���h;�b������{sUkK�	� ov��k�&�8
���0���Ȁ���.��,+�٭�߀7����s��iIa)w�ϸ���t�öZM`V~a��35���lU٭�ȃ�Ǔ�ȀH.M��&��޾�����ݾw�G<^؉���6�6Z)�����קЌ���b�|
�޻��^V����{3*�$Y�����z�;��J�U"�I����^s�Ȁ��x��>�&5�h��H,�e�@ kΧ�v���}��Z=>KV=�����6�x,��.r%{��~g��y���$I�6�����[�{o�Uʶ��`zǾ���W���>��ۧ>Y����ę ����:��희g�0�hp���s�^v�ޡ�z���Z�Îݰ����p��n���טrI��� �n�Y�Bޞ�ź��i����7\������c�+c��w9ru�v6�Nz�⎞���ӄ��|����wh�=���+�:4�c�rs��Y��a�I�J�Z q��C�Uwex�vph�M�'L����M��9'� �5bl��4�I��M��ɼ�������s�Msʶ�óر-���g��*R
�W�,��p�A�6�� @{w�3U����+��ֺ�
���@��כM��>��f�jj$�(�m"����9;S���B9��/fm�h�{31 ���&O����}�?\M�@+ lcOL'��� }��x�{a�s덈��շ�"�6� ^����=q��z� ��"hm�5�]�V�΅;mW �U�@ >�����w|��s�@|}��0���FR��!6�2~?9���&=7�m(�|����g�չnچ������wq�*5��xz'����3���u��\����6ݔר�X�dh��>�gTԊ�J�����*�4��&j�7�
��p��3w��� @�w.� �{w::�oK&;;iTDͼ�'��QB� �����p�tW�zN�nnW��+��3��lZ�/xfnЅ�Zk�����u�__���ݙY�J�U{gMS|�OB���C����_���$�/{{30B�z�́��.4X��uL�(�����&b�*)Z�x�3���^�dDD���ǍQU�e���j 7w����!u��`��.�P�QJ�i�nV^����]t��׶�o;�`A{�� �����ܱ�ۿ^��NXX�����0����� gO9��k[�cw���I�u�݀ .��q}~��A���Օ�W)�{�������N����2�]<f�ms�Ϯ�Wm�'��@>\���o���>��&d5B{�=[�f` >@����`� '��p¼RS���*O��ݚށ�B�^��	��y�bǅ2%&�0
��E�X�omf��V��÷y���on�}�M�D@�D��vF�_=��-V��s���*��*R
�P�oo�0�ͦȀ1$ȿF'��$��uS���we	b��ܖ�-��0��;�s��U4�7�����x���4���Z^�����v��/�����M��V�n�*��%��	G������{ۉ^,Edmf=��a�*=�9�o�WWz�Sz�u������xz��������}`�����eɁs�B��{<������}�\�/���sE��oBJ^é_o���$M{�A��<==�!�.�u:�o{��w���Jl�ky�ŵ�O�����28�&��W��(8�����O����j�����֮;�(�<��ì�ݽ�����{GY�b]�Q��}+��X�/dXt\=��=���9�\������<�}:���K�et����)9��dÛm������<�Ӽ�OQZѠ��F�����W�����}g�K���)��j�c�擓�˯n3�B��\WnI3��M��z7��pq�I��
�����{P���޾����{*�g���f�����-�S�w��_]:�w�c׆r�7�e�Bջ�9�
�	�z^��g�a��Ti�Ǽ5����ԣc��L�۪0:8d�yN����z��x�ŋ�����x?^'�8�OqǕ���{���m.-�f֒�o*�z��el��Y[Q����ݞ�cr$^�O0�^��C�4co�OE����I��/=|��ޤ8�:��ؒS۞b`��Ʌu���{���m[��OG榬�����|��ֹ�>�+y� r��Uf���F��|���Ԋ_n]]�o��3�'>0��{��f�ߜ�9�˞"*((1Ebq���-��(Ԩ�[J��UX��m+V5(�+Q��
�B�mH�(���
�R�b0amD�[aD[j#m�+X���*�
�@�+ER��ic5TŔC�UA�[���e��D��Ԡ���Q�V�-*�����%�����-��"+EKeQQ��J�؃m�6�[h�b�*Q�6�TE�U�***��H����T�D�p�Ym�J��(*�����U�J�ҫeAdTDdEk*[DjJ� ���V���J�P�K-*.�e��Db[U�Z�EDYm��k,U�iF*� �,`�����m�J֫b[Q�-J�ba(���X�ŋ����k%J�-����UTDKF�QF�ŭ
5b�Db((�����U��R¨5��h�%J
ŏ���Z� ���l���6�@y���D6	4ӛ0����X��?�S��d�k@��m� �{���>{o{1�N�L������ޛ*�"TDҨ�dE���ɑ��<�O��UO�T Fg7l"����� ;o{������N1�G7�&�	�h�P���Kg��v��s�ݑ� �5'�k���}{~�
 *�DL����6� �m\4 ����#U#��λ���ϛl��y�8���X�@�@-���W������2?���zq��˸` >}�n �|�2 ��9�D����t�MD4JO
��E�I�O�}� 2�Ȟ��wkd~mߐ |���l ��}٘��ϕDP
�T�B7]���+�1 �@ �^�x� B�>�Y�(-��<*X�G�<[�^�N��z���ۜ�&{�H������s���[i6��_=�v���8 �}%o��ˍ�Z����/6zҔUq&�sG��� =���۲�y���Ǵ	�v��f��dF|�o��C&{�bb����� ��������ƮoVKf��V1��H#�C��i���a�������"TDҨ�g��4ȁm�<��>վ�`,�O{���(��3�2�A�w^�dFz��F�B�
�Q#�޼�0Aiߛ3�&p9��z�7��7�vf| 	�|�́��	.�љ��s�x/`a$��~}��������w;2Ź}1�{z<�-׽� s��I����{10
d4JOor�3��4������gs��6�]���)����ʲt�x�7�����u���*& T��s���`��r�gl,�j���l	 �wf�`D�u�@nSidY��uo��/�{x��n�k7x���A���NCAɣ��:����=5칳~Y��(k;��8&��ryvu�8y`җ]��<p��e�V�=Vy;9�s�2��6�ln{{Y���ݍ�F_vn���=ng��g�ۡ�s�l�Z��FI���G`ƘL��nݭ�sv/F.�<�3�5W3���]�'v�R�t�.ny�i�V�s��ݷf��y�_j轮9ǂ��h�63�l�3�Q�\��X5�؜��v�6�<Ը����6�v��8���U���Lv��� s�M�g-�gL�]��v����,
2#
ǁ;;�ًg$�N0���>$ջw������{�����֥߻�$���M��7Yc�$�'�u�1��7�����_u{y� �k��A�q� ��uyQws��=ٝ��G�1
 ��DL��.��i� �g,h��At�x��]ۚ ][��@ �g�C��P����4�j�F�w�s�,���;�� �=�� k��$��q.j� /���	��f&L�i���MߗO�N4��dX�Ԝ�4�5V����DBC���s���˕3�2��r�">���웵S��72�h��.��Nӻvb��uVG��=,k������ޝ�7\K���~~�&vq�>�k�̈���˶2�}��:��{����٤�Kg
%2^��ﬃ�%!}��%rX�/m_�j;bQ��p�W7��DH��w�.��C�:�hG��v ���vs'���m�a3*"��f�Q�
�a�r~�_|� {��D0k��ĀA*�W��Qŧ�~���Ǯ��LIM}4Ɛ^��Do��ϰ����1�.�S����D�e6�"罙���4 0�8FL9��}큡��$/{��wgfb��u��������p	8}�����e,O	M�7���� �^{��e�
�Q{��؍���� =���$ ��͌��T�}�߹��ǀ$��)��m��Uo�Ϝ�>{g�@]�]n4�7<����T߿����0,��LdF�:�� gvs�������}��㵺q�@wk����*�LD�TL�Ъ�[L%Fj��y<ݣ��wk�,�>�Ă ��i�5*�����gϳ��[ٴ�MQ�IQ2颻�q�B�ݶ��	���B׫�~�a�u=O)P��G6����y�6}�@�ayڇk+��
�۞տ����ZI�/ �g�՝��_�*d��]�,S�A������G�A���"0_�[L=�2�hDĀM|K�ʪN3ݱ*�rPV�<� ���l :�����|N^�z7�>��vdF-�AҡB*hQ#/�� ��{M3�D��K�����fDb!W�[_2�:���c�ܟ������|MXm�<s���qDO���Q\d6,�)�	 r���}�����dn٧o��^gf` V��d@�]om�	��=�.�>��ٙ�	 ��{[L;�y1D$�,��hHK��!g-Z��{�}���Q]��������Uz�j.e�2�_[�K\�U%P)��J��B���|ȁ[�l��`VfN�Ƴd���A
��� oi����-��L1���(���f��;N&Y��~��W�m&�u���� >ͽ����ҿ��q|��l�u�m���x�S��u5{���c�8P���_/\����ٳ_�"w�)-J�<i���:Lo}q.XF�?��L]��(��< ���m0Y�qT)&	��c�5�SdA�o�y�2�t��8�����{V� u�fD.�#��Nʾ����7c!�^�]]f�"l���u[�`��Z^��B��H*����P�4(�cy��m0����  K:��0":�VT����}� �u����Qx��LҒh�-�y���
n�7h*���F5��[`� �~�A�{٘�	zw�U��f7�
���z���,0K�Z0�ǵq�:��a|��E�}��s�]�%�ބDe�U�� ��{3\�U%�B0�F�����!�U�a$��U�A,���π U����ޗyWI���܅�g�|w<����������A"��,��n8π@��m�?w��V�TRe<��o��q*���f�ܨ|�h�K����]vWt�Hep��B���ɟ�z{w����[}�&���-{����`-F���3]���>���d��ܚR�󁴹%�S��Xarym�4�m�v����4:9�����w��9�֜m5�vϩ�Ce��Y��ukr�p�v�#�:����y�\��[���&���[����=^�h����3�4Ak˦�n��{rn���S�l��Iٞ��k��gF�]n^m[hc�E�	���A�;t��7��.\xwB���Ecd�ٕ�Fޒ�ۇ�ۅ:�S��v��[��/h�����t��kM�s~7���LT)��U� ;�y��(��v�9z�E�(=8<ܧ��vf��*3R���Ŝ���k^wW�s*��o��D /s����]�k�	#t��c����st�DG�h�$�"�`H~�ﻸ�N��n��6�:=����o�c��{٘$����?g�lL��X2Г	}�غp�:}<P7~�� @}��l9��$��ݳQ����s w����`�a��3�����?=uq]�<�a�U��b@ufnf �B�֬� C\�(����":�N��θ��F��a�*�ی�.1�N�x�n������4��[L��q�ߘ�`��J/���v, )�m�D�]�a�s<�/Vz�����3 )�si�^��UIe5�C3	�J��N���z�)�Qt��T#�΢��r��b֟]�&�r�u7�P��C9���p)����eƷYK�=��Ȋ�mi�$��&�m7���`A��qs�V� I/��p�X�L�����n�h>X04(�b�gc�2 z� �x���̷Λ�� !O��q��`y��Q�fhTI�%/G^=�uڕ7����~��w�[}�က�5��ՙ��ցX��>�;z��Cwq�&�QQ1U0�+5ט|��,7W����U_�4'~E�7q#��V�@�K9�fD#}��}�U���"�3�5&^�y���vg���0q�po]����k{v�v�mK}��� �0)��n�'�@?��}\ϘA�k�̈i"��ٵ�P�(B�� @|m{)��
vr�JB"K-���"��&7�OW�{��� |_z�4�%���3�>~���L�ݦu�G~���}ǳ@m%������ o�s� >A1����gn*�R��d�Uu��EP��O��ǲ��r���B��{��i8B�9ޣn|'l'��ǭȘnM5�*��5쩔;�v�3v�� ��7�5�7� �t�eB��jTQPث;��q��s#k�J� �~��F��n#���˾�ˈ�a���{�ra?�p�-�Xl7������ǝ.bp;}��u\4�7_sq���A[qԷ1G���3�i�rE��3�B�51V�V̀�L�\o)�R�XG��������r�h(����s즓 f���D���G\U92��G�s.���K���1 �w؃l6p�1�!��=7�B�O���߶�� 3o{3/Wki2�D5ּ�O��ߢ��9�Y���ԗ<W{ݎ1 �/Wm�D0�������s�lh �u�fDD`�]��{p�QR
j
�TX��r���u�7����y�X |���l"�m4Iw��r/jf>%����F�Ϩ��ǚFm�[,x�Μ=�Ytz��tŻT�g{����뷆n�n/Dm�VD��x�&Z��J��30=q'�vT ���QQlU��p�@<�l�WN��(�)́��vf �]]�� ��M��B��(ɜ��J:*bD!ln��ΰ�Ӯq� b
y��v��s��מ\�[����`E���~>���;	8Ny�۠>�p���P�{���2���s"1 s��M�(����a=��d"A�7N\�|�7z�]�� )��a ^פ�uE�*-�9��j�x�J���&�Q1c;�p�>�0 5��vT�*sރ����ku�@�9�ϼ��OO480Z�F(_��������˜��"�;& �^m�` 3��2�=�?7&��B��m0�1�QT�UUJ���)���mfB��$�]�����̚�s��"	���Q�����K�z/�&�vՅ{��i\��i�rC�eI������.0�Ń\��sA�^��ăcsr����;���{��$f�#�|��z냎)�r��'/�9d�2�=kM����{��o{�=�~[�a����k���U;���?z���7=�	i�c��rg�w�C��{�f�%o�P�y��-�;���|~x�[�ǺV��H�����Fp�2o^�D�`雹�.;6\B�4��Nb��Lz�'V���w����/�ɶO�t���_��5|�����i�����{���`�3�Ɋ{��:T|`��V���{=\w{���]HU;��7ٓe�ΖJ��wҵ^��dn�n�9ik�[M͇�|&���ǚ�3�ۢ_b|�{@V���x5�{��a;�s<N�G����ط؈�8��w����E%���[l݃�d�1�O��پ�<\��&%��%玘�j��w��V3Wu��E��Y$�p�o�L�فt՞8=��\�es-��n	���=\V'a��˦h�#�����=��p�x`y�y�E���{z�'qu�RVN]�,>�����'��CL��_�w�8� �^�5��F�M��*�0P�}<E��/A���8�d*�嘏I�U���8��i��o��� �ӍI�ٹ�}�(~���Ӷ�]pӶ��Nf�}/�}��\5���{{���s|}s;��w��O`r�6���]ˆ��b�����@;=�\<=�5��C{����s��������{�A{o�,��/K3]���$q�]s��ae���ٽ�<,�b��C��Lfh=������*0UŢ%h����1k*�
�TV#��[F��Uj��%�DQ�Q[`��*[UDjR�bAdR+1UDQR�V��,��+*


�Z1Ub-m�6�[X#Q�R5�mT��6��Pm��Vڬ[h�
(╊�a��Z�k��e�Q��"���na,b1a���U���,U�Ь���TR�UTqeE`���\XЪ"�XV�؂�[b1V҅��H�dR4���R����T�����b,F�iYmV+i*F�����`a(�* ���E%���UX�aF��(���F�V1kA�mQaZ0D�)XT+ij�Z�b�"*�T�f-�* ���T�KeH�*"V�ҍ�
*��QEX#S	�"�0�b�`�h
�����UPUU"�@b(�(���{��w�>~rg
T;Tm��G=�r�9�Fës�/U\��q/c�k�cv�pF���ݩ[�"���m��rkj<�Gukg��Z�6�ӣ ��v�����xΐ��;l�9�S6��x�\6:z���<��5a�um�Mpd��l�5]��y'uke�h4�ܫ��6��q�v-��[����\�]Ju���+Wm����۱�kl��v=�t����1h�=8$��;Z^�������.�q�s�h�K،d��x����fzύ�'�G9��U��L�����Z.7.��z K�nb\�n���ye�V���R��*��Ǌи���Џ� <c����w8���r{����ڶ1v��ug���/��skY3�æ"�b�8(�k��+�3s+)(vMu�x�N�lh;5�s��g�.N�w<v�a��ݡ��qF8 Һ�=��Ӝ�6ۭ��xC���SV�.竴S�KcI�W��M��M��
'�{��m^Y;�����nv[n@���9+���<\v\�p�ֽ�f����G�����7fs�X�Sn�Kt�W=n9���Y�ڮ���ɝ׺��Ggy�<��y8{f�rFO.�oe�-��ԛ���r�J�z�������q�v�#c�ۛ��]ñ�f�v��,;'6��=�nۣ�z��:��u�v۳6��˧6�Z���9�a�n"U�kly:7l���<P�˻���ଶ���`�{to#t����b�T1՝qw#�t)�y�<��v{>�z�n��N�&�����ў^ :�\^����m��#�J�i�:��u!ú�vS���=K[��ٍ�V��8s����h+d�Oe<n�T�Y�݋sn7n�{ua�4y��֟'��Ԓ�ѩ��1�n�V8wB�1��I��#�ݎ�y�z �$�\E\�5m�u;�k���jn��H[G[��Ɨ�&��݇vų��Ov��[���m�N$�%Ű�����u��=��ϓ8�2[�@�As����)�ή�pv�0x��y6�VFy:e�:�Tj<9{n�vw��D��t���\j���p�zw�6۶�^��r\n\�+�;q���dW�ؚ�X���v�ۛ��9��gv�A����8��C9���Dח;�ԗ0��j۟7CrQ#�+��
����n��@ݎ���ő��ݮ��
.5�)½vm�=�|��od@��Œ��õ�q���EL�(���Mﯓ >	y�p�@$�_vf�4︛q|�},{�d ��=����+��l���w�0>����v��^�˸Ј���^�������k-ڻ�甅V{�&���a�$�{g��	�u�7n�꼸��TI���z� �%��"#�]����*��DMQ%A��3�n$���t\A;O�& |��� >}��o���_�7���W��O�Z̖���h���c�H ^�;&Z�)=�О >��[��7׼�$�����z(�-����L��6]�E����`aM�&]����[�ф��÷/0d1Z�pVDn06���ܣ���yj���*���T���r�����  �g7m�ۺ�}誼����Y������8/,�l�L���Y2OzG����6�+;zk��"�O3r��sB�x���*~��~���h6!z]��U�N�X`���[�q]�0�Gf���ufȃcOm�+�,̕��|@{�ݙ�/g;2 ��u�ޘ��3v�	<��*C��l	0���f@ ]���s���y[�]S<"	��o0�s�4��y�;!DM*���������ۑ�W�? y�y���3y�h*���#�����/���S�q"�x���(B����Ұ@ ���(���tOf]o٘�� �n���""���ԋ8v�9r�Z�����k��a�,T���g���G�=�-���Xu�Q�y̧g�����w�L"�Ԏx�����u�>U�y�
�ՇJ�S����0���Y�5j���T���dE�K�r������=7����  �n���W��D4��(�v�U�����5:�����6�	� �����@{�� �pk�� (:ny7;����s�V�h�}�w�<u�&�z����)��P��y����=*H�x�K��o��NըZE�d	j�+V���'	8`��0!'�{�b'����ʖq�i�!~�ޓ�˄��@�ڰ� �;�X�}�zn(�f\{j�����a��G�4)
"iUL6��t ���,%�#������he먈����mI n��N�V�o��ٹ��~��L��O|�%��u��+�񓵍�]W�5G/;�A��\����~�UJ�UQS1�#��V"*�u�> 7y�q���Y4�������"U������P*S*jG-y��� L;�Ur�����Q��^c� �fDR�ᕒWa��η}p�
Q�DUT͍ {�������� ����kSG.�`x�_����$o>��<�FFԡT�M�P���Εoy��zgs��F�]�X�@{u�f  {��+.��կD����N�ʖ��d���f��O���\��unuz2\fNP���1:&�Y�3.�e����B���'��.���$}ڦ�?y\�R�6m2$�_����$=��!qo���[�ƀ�|� �����s �n��[������v�a���&4���򟛍����N��ڞWm��:)��?#�b*Ъ��z#��^RLz!�&�,�@3��4��9��ɢ�ת� H�>���<�*��D���b�z6� 1�~�W���ٵq��O���I��$�n��b�$�~} �ojae�1Q��r�מ����n���ݲ���\0>@}ݯ�"3��ڰYZ5jJ �U4Uȋ�:��^q���Hy�n0;���@���b+ם�5��ܧ����'^���nD8|�m��ca�~��I�KǴع�w#�Ƿ����{ٙ� #�*$�.��DE."ɫ��QYR �ﳴo|���s����{2h6�j�K����n.����j��]>�x�A����3��ݓK�ETR"aR	7.����*X���[�[��1�o�ͨE�۰����k�.c�A�u*�[�q�pq�Z�C�]�q�����u�;��O�z7��6�vG��n�x��y����N�j�]�����nz�]�n�4\;pt�ma��2���W�l��!/N��s�F簗"$&�H�M��#����������Nx6W#63x[���>�m;�:|��	�͹�v��n�qڣ�M�������m>�Q�OTQD�S���~@ q����ᇛ��P��z��=�� >���ٿG�4)
$�UP�[�0�ZF澄'���7� C�n����8� �z����o{B���?����n&[x��+!�s�x��AW�M&�Ϫ�"������،Oy��0
��7�y��)�IL��7%�֭�%���t��DD��0@ >�޷;y�j�oéA_m�<��%J��*�dE��y0�A9�4���(���]A'�J�O:��Dv�sy�;�1��-W�l��q���Z���v��Լ�z{]7����;n�Ƴ��A$�b�&4�U	UTjh����j�!�=�6�v�vf
I���w񱽭�"������O�**��&b�w�������'��#���d��7��`��[��������׼)/�X8��*|s׬�w���̏���G�qy��J���霔�Y??ۿf����4������#q�^Í����}��1D��jA�ܦ������L����Nq���ik�a����@}���ML�"QU1R��tm��o��*p� _v�`�#}��;	 ��L[���)�;ګ�	%��Ʉ����Ɔ0�Sϯ���t�V��zFIC�bo	�]֊��"!ww�3���_��ח�uY[�o��/HlyD�{�Ւ�:1�9�gWp�l5�����Cl�O{���D6�eS�3~�Ϙ �����#L���ը�^�{o�@ w�z@>��)���@6�0ğ�'�1	�$Z��;.�߽�A1���`�$�ƭpIZ�0��*���$�^�*Be�S)�wK�ND�r�.	$�_VS�=9/����������Ӹ:{�y �gI���>�Ow6�OTM�'{��gPfm>W��#i{}p�ٚ��E��� ��vf ��6�.{�zSDIS�jG��E��M���B�r '/1���"�n� "�:��Rpʪ��G���o\Y�RU"QU0T9b�w�g9���Ԩ�a'��u����Y(D��ɖJ����w3&��D0�ܺ�T�ap�<�7 pV�X��	�PԲY'i��w|�/��`$Q|k�}�Ē|	���D0c�p�W߳}�^ŮK�a$�I�g?0�ı�S*n�՝��r�vT���T��e�+Ri n�M �+Sa�,�+�;��O�g��	��l4�0��X��/_��""'Y���y��l��}w�> ��� @"��6O�3�UL�Q5%/Es�ʻ0�3��P�_�4�v��& �~� ��vdUy�z�����ߝ�L�.��Ǭ��v�>ջ��5�W�w��^�f�_CϏt:�n��<�f{�#�I���j��4�#iJzF?pF��۳ٿx�h�J�4\G��y0@{}�>������~��k���� ��S�����u���}_�>;��'�y�a�� �"��=wY�۰n6ֱ,��a|n$�t��mu7����~����T��z��mX ���M� ����Ii����h_>�L�	!�|�/=��,�W�J�\��=٘ lTN�G�DN_�h�˻� �.��q�]�����6������tu�M;��o�>�Қ�����U$�,��{^L>og<�@������ꢲ�� ]充A&�3D%{8�����54`�4��ڽ�?��u@�� >;�� vp��R3Ͽxߓ�tJ �Y����6�2�m$`^��@ ^[�j?=
� }�� ����� ������1cے���EOm	�װ�s�Q+�Ԝ��.k���=�$��v_\��	��C�$-����a䶸����pxn�M�G������^��w����X����+�g�*N��:�G<]S�J���>7�Flu����{-�AF�ӹ�ւz�uf�d.��<�0��C�Hh�#�|g��p�8��ۤwv��e��q��Jk�ϝ�Q]�������rjָ��UL����j��۝i�/�l����N{v��t�'�N��D�Am�ۉ^�q�[��&�<���WL��N�7U�f��S=-m�&�B�{,��t�6���ԭ�cc�K��y�f�-%i �T��܂��������$�}�r��-X�w�o���5�߾'�鰀�����\EϾ*�%2�7������L{3�2p��E�z ă}���g�ޗmI (�{��T��F�/�����hb�ay�
`��>�������� }��˺���ʗ�@ �o�2#Gw�ېYZW�*�LH5&�)A7z�D������x�S����w���y�O�2"&o����'Ĝ�	��-2�0D=Wl���4ͫ��������� ��m� �:��ʇ�{��.�����q�u�����M�,n�)�]D���Z�!��I"��P>�Q�P$��*��倀aur ��Q�ڽ'�!=�w����|ǻ�ې�p�)O�S*!5!7}�D%���\ZsN����x0:�E͉=�����b���{�d]�����.�� �9WJ�<x����sԀ��cw�{ݘ��o`| �����[Φ�TZ�5��j��u�|M����0V�\??.��$�L��� ��̽&n$�/��{��ޜnH�>-�Si ����IR&��L���ۺ�{���V��J�w9mI|�V���w�����"�NWe����~F������2��0�{�B ��<�w��u��֭������:�A@.���������&�eK�����������A��d��\7I��y�k�8��8/o�e���x�`���SJ`�k�i(&D��fz!��a���_� �S|�$����	9�w�`�ē3-����R���T����� �ηA�ݹ�� ���}����K��#`*H�	�D�VI�{{^}��	�������V\P�'X,�������%r�{�V�wl�;w˽�nyu�B�K>��fE9/N�A���LYY���1���	U,���f�:�F4o[�0���^�o��/n@�N��g��w�`��aB�=7��8�l���;��K^Nv�CwVe��Ez^��YA>Aw�Dk�˯Ͳlb�?QE�6z�����)�w���\�]]�s�QsP~ܰC����LZ�{�d��	{�l-��v��;]�te��I���&wc���=0����c�i��g������f�����*����r�>�T��Q����3�����Xd�:�B�猶g��p�(2������:���i�A�ߣ�S������O�ρ��'u<GU�Ü�8�~��]��:�G�6*J�郏�rB���˸�5f��=s���}� �/-��gwt^��xҲ�i^�z��I��]��a�� ���ހ�w ��}���a����;iȻ/,ػ�}��� �ӫ���w�k{N��MǨ��6��\�������u�y�ѯ9(�b>���։����/�0�y�9�պ�w�yz��E۾���=����zr�!6縏v��ۏ��,�.u��=Y췚���࢞��t��	X���mv�}��	������b�B�_�����l
�����ɂ�ѾnC���&�zѓ�;�V�Ҁ�{T�p5T}*6y��u���n���Q�ɋ��
�I}�+�G~��;�@����5�L;9�ś����Mo,Ӽ����v��g.�Т*�b�aU�HV�b��b,b�++F(�"�F�m��*,�L	 �qB���@���E`*�T�R�Pc"*%q��P�a!KJȠ�P��TQQU���D++�Ȱ�m�m��m �E�YZ�`)�Ub�X�H��1EF ����%L8a�X1fPQb��C�W�!R���+Bڑ-%L5!���6����Պ��AQ�b��V��+$�%`QX�e���n0L"����jE�U���U��l+Db����X��[��PA����"��R�a��
EX���)�W�-�)X�PU��aQ`a�ie�!�4**�c�*A`�fYmX(b�EBVE_I�!���s�$V�S���v�nf �T���Q5��]3�^2�y��=;���6@��������[n\;��9Ҹa&�f��Q6���dIT�R�tͬ��X����؏��kw�@%�yn���s3�0�e?t��e�����p`@bO$�c���*;4�u{E��&�6z�չ5n�����"j���j����� ���`  ��{�Y���E�V^Sa ����pT#���S��Hf��'�D��ݣ��o��J��lv��`�e�D#�H��똗�7���+�9_К|f\L��a$���fq��m* =.'��WϢsr�D�ݹ� ~;���/	҅?IQ�����UTJ�b^s^� ��ǘ |��9�h����Ș�gr�W�L�{�}u���:{�V�M�q�`�7B���䍑uQ�ݢD�ԍ.��q� w�ˇ��U}+�]Ӽ����/��T.[���NzK��Iώ<; �L��t��/�@{��c�ވ7ס~y��DC��n��
���M�S�z^�wn��ѝ��ɼ���A�.:M������۠�b��8Lax�'�j�	/1��%�Ͼ�8�����A�Y�n�ѝ���~��Ā�5�T�SQT��%TTK[�SL>����.�ì�����@}�:ܰ�
��l �7u�E|�g�ϧ�I����Hi��m0F�gz����"+s��|�22/�TI�|��� 7m� @�O��4l$��_���_=����[�Ĉ�<��@� T�m�@�g7���j�/�~�/��I�e���
N�E��+�w�B��};�u�kQo�� �m�@|�ӈ���{;3Dh}�����Z qT��/���5w.MW\�`�h���]u�Q�-�����w�-y�e� ��ͣ��<ە�n7�ϴ�5�^�����5��a�.9x2۝�W�Hxtt��nqCG��l�v��%7b�������^���<F/fͺGļ�ٞ�nw�'��T�i6��7��z���n.��0���pq�-w٥�d��m���ּ�f�6�v���vM�\ȭ�n�7��tS�v�y��A`j{�e�:�:}�:�g:�=�ݺ�q��p�����5�x=k��z�X�۟F�n7���c�%��m��R�6LF��cA�fwO;����vy_��؏��jI
����^7`���`�����+�����ޅ���7dD�����٥|�RU1E)t�GV{��^�6]"�q��� �m�;�<�I��8]WbK���X.�)���RJ��*%� �ͫ� f�s�"DLNOA8�> ߺ�A�����:^I�$T�ETUMA&/�{�Q���r�c�Ȉ���٘��w�R�*���E���lv��=�J��&f\Ovc� њ�6���u�dt�T@���Y$�x�	'qƣ� �w��_��6����,-���׮y���:�۝��v��F�d[��玻�6o�����t��T���?|��� �w�9�������z�=�>R��<�鰁 �w;3@p,E�>�5Rf"�*B�Ĕ)����n�&�,���H8B��;]�4l���/���m�{6��͚0�l-��;n��L�ȹ2}�y,���:��Gg��������@{w;2#�;i2 "��}Q�O�s����G�I��R+�(�7Zug�1`B��m� 2s\�_uz�5��|@oo�3n}$�����$�)�AC	�~w���;�W��l@�en����vkv���|>[sތ��w�7��y�) �l��XD��! �C���ݜ��ȯ)���=��� >@٭�A�$���}_w�H���~�K�D�q�^�R=������@Jus�s�m����EͰ����R7⾪����E���İ @�5�`
��h##���:���*�{�0 >�6�ՋÚ��)*��o��ܦ�W�G����{{�� i��0��|�f	.�|���J�}�oYDgZ�S4Q U'QѴ��X ��� 7}4\W8];=�S��z)�r�G��zX>��D�Ah�9F���鈴�y &�{�gv�p��Y�'6�/|�s0�����b��@ z3[+ ��V�K�J���W�%L�5�^\cN��w�Ĉ�Q��B��is�-  ����͆Xߣ.�~:�cW�e/�� �2�{�������;���Z�㶗�/#2�&�jD�}��s3����A�=�J$�C8�d��cѭ���垷B���u盶9�sܓhx@�X����߹��m�ma��Vo} ����\ܠ�K�uV����%��ڑ"8�@F�+�U2��+�O���]���A�s�\'��}� I!�Ƃ=7��Ɓv����C*fhP�0(M
���I{��ȼ�Skz��K�{�|L�֐$�x��(-y)�(�*�q�S�5g�9W
��N�Ƃ �3�@���������7x���q��95C��y� �6��NZ��9����%��:��n_h�6e�ʞ۞���G�L1HwҐ�:j��x2jմtW��5$T���nV��$uC��zz��pc����YaF�Ƒ>#�;�7�P3�!s��x7Ln�pm�we=�wY�g��$4���=�p֙�Vf�S$������g��A\~����綉�yCQ`�x�.&q4z�X�w�q��l�X�o�q�y���W���=*�f�|O�#>H�O�� �m(wk��g/��=�zj�fmz��H����D�0
un(�J�$���$	�)�^�2�&����P��ԝ3�
ng=|F��h�I>�\�X$J^�}��-j��??o�eWܹ�6�$�R,�+��O��:#�vP.�����_�<SR,�\����fŚ��e�Y�N�y�"�`��nR��w��G�����φv��T8aϽ���p�o�P�����o�^���og��5��שy�;cgճ�I��۳��A�E�S��wa盶���ta��b�\;���O/b��}	��J��z��ۭӹq�Y��N���E���嶰i����vTsM�#�k�1C��t=e�!*��l���cě���o6�F̸x��W�����t��u=��U��q��N�f[�������8����M��s�N�
�[�mZz:�t�F�nt�-݉�6�N7[L����v�\U-�ܴ�2{<wܨ�MJ�U ����6�B�C�"�!R��-�X��؅�jᤱ!� �D��3%g���<x)���`;#*���7��I �MM�J��"KŪ�̮��U�^�J#F��jEDML	6d�����Ё2��ȧN���ۼ��]�8SR,�I���thفצ�&eO;ˣ
(՝,����rI�-�	�Y�	���۪��\���I(˻����d��$L��4*��Љy�E��Ӭ�5�l����'��h�#��=�I��JD#�	�x,?�L��řl��#�^Gv3ձs-\s��멿?�C}�մD�F��Һ �����6���\���V\x0�ޓ~+��^$���`9M��l\^MY���9�D�KG���.�&��G�!n�EL���f$
�����S�]�s%��w�٬ǋ���rc���h�E���0����x���A�B�Oi�[QQr����W�"}TI�2f�I�Z��۴ �Wqo T�J$��$ͻ^v YL �MCp!��L9L���Ų;���Fo6� �/=��O�ic�-�� ���-a�H���ԼH$�qMH�Da=7W}�H�RD�i�خ�Kb��3s�/{n��c�x�T���D:=�,i��Us�u�hہN�>�t�����S7��u}���h Oo7kē�v;�;��Fe�ִ�=�ݢzt�X���""f�#�y]J�t�DMI��մI�;ʹ�$����~1o$m��KM]<�	�WEa���H�B"ǚ��$�t��Q'����],8qQ��©e��Ff^)jpm�&*��iCY׹�)�q��}1.�J W~S`�sϝ�܏����Go�˭1݌O�six�@:y+�څ�b��Td�E<��v�L��̀B�{k��ã�H�@\��g��jop�[z� �S�$�D������&�h��(�|v�
f!�����2k���v��x��%[Ɛ0�V���|N�RI��XzB^,��cu�n�-j��\�2����9-ʑE=��䰌xP-��������w�[Ɨ����w�3��iH�=7�����I<,"CǍ�}`�
�gk:�l�����O��� �x�� ��K���/���UA:���lZfעO�-�$A ��ۚ��{�QNN����;c�A�x� ���D�35(ER��s�a�R�y��f;RH>w�� �m�&��J�"\:�o�ϵ��؂���d�÷�AG|��~�����F�|P��7�sH�\�����(���f����=���X��j�N�^�Y�W93�6�B�[$�}`I��؈��Td�@�݈"	9ͻ
6iZ3�r�qΨ	{��>%�I���/��o��&�|X-��l��[=ktɍ\f�p�ֵ%�iE+��6�������bLTL��E�[	߄�G^g$	|۴
�BMonX2�r�]��@�t�QR�1�X�I���d���<�0}�9��F�cH�K��@�l%��p�q8|��4Ma33B(�A�B��m�$A ���I�0�s��7"�_r���$�e�i|Okm鋙���""�� zb�檽T�Y�L����H���^$qx���eģWwb�$vrԼr�K���&jP��_u�"���:���As�&p��wd�B{܂$��?z$��!$ I?�@�$��!$ I?�$�	'�@�$���$��	!I��$�	'� IO���$��!$ I?�BH@�~!$ I)	!I���$�RB���IO�!$ I?�BH@��	!I��$�	' IO����)���}� ����9,����������0Vρ`         P ��P)D�BU@ � w�H��U*�A
���RT�Ȋ�w�ݩ�v�;�v;�\�ws����I�zy����iLz��*����F��ݺ�k�<�6��ӻ.�� � <J�U!g�۫��g]؞s:���%h{�7����*��   V����� 5vţ=՝T�pς��U{@)��@�@��: ��
��A�}
Հ �s��EU��EJ �@V���]�	� �=���p ��b�)E@xz�)��R�Q� �7L�V���8û���;�<��Gw[���    Sb��OPh14��2i���"��`�UJ�`       ��*�
RP`M4h�b@i��%*��
0�&�d����2�S� ���	�!� �b`M�$M &M1$�Fj220��Rp��+�c��%�+-/6���X
��,w" �p?(4#tUG�������!qev~�����?�����A�B@ZUA��@.��A����{t�~��]]|tE҇LY�WktcwIQ=�ݠ.||A"?o�ܿK��4��������m�[�wy�����&�۷.�&�eL�L����\tsO)/��t�<�:[+5	��Z�+����T@��F<P>%5�	Ȩʱ����q6�Lݯ����{4�����7�:ܽ&3���sm0Kd��0�ZwSX�w3��7��܊�ΰ�-]�`��@�K�q6z�s	��r׈4T�0l��1���r��[����*f�S�C�7mԺγYb���7qv��a'aP�4�hb=��{`��3 B3Äŏt��l:qnD����^TY��cS�]��!JI�ɑ.�5eiٍΰf��\b�����wt��wC�8�[���<LnI�<�� v�I!f������O��`�b�gCn��g0W�X�q�4J�֚�^]ܴ���)P��6:����
ћ���rN֕�j�Tn�t�{�(\I�c�5�/��W�8tO	5�צ]��G���KR�-ˤ�ӧ��MHcq�x��5Gscwbim#���j�,�萍L�Ŗ,�ix��x�en���=���Ks���/a铟�X�ib�ʬ��gQ��t���v �7���;�V\s��^	Y�O^�jFYZ�; ���Ѡ�8�{�4���"{N��8;�@��*l�XTL��h�IV��d��=�w^�I�EV�����Su����:cҮ�reO�t��G2/yn��Sc�`d��C6R�~���-�W�IwN�ǁ�8n�=Gp`qT�8��Ƙ�#�P��%�[2 �Žk<���=V^or �����"x]6sƩ�O��Eek�)M Oc114�s�j��O�,KJܳ.�#C�E�qeN�>���r�>5h������pɽ��wL6"8v�9
UI��5Å"'L�5��U�>�t.��=ы�X���a�`��@�p$IO(fa&Ŕ�ec���b��f;R�m��ci�{-�*�o�=-��N�9������2��wh��7�$b��I�9��$�d �q��}���:b��Q�7=�t\ݳ�Έ�M��(7��
�&�۳{c{j�ݝFn wa�)�t����;'<�����#�tɰ�}O!\|�4^���ķ�x٦��׍C�>�x]��ohL�5�8�H��4��{۷��'v�ۇ:X��"�Y�&�-��7�<���_k���/6��f^�����pv:��շ$�*�;�����P8N�]�ocB�����v�w� ��%$�~�߀6���c�iի4�}�kP-�6n���̎t��wv>�Y睋k��������v���\��X5+���wt-[l#s{��C�øxEw6W�^�IV�Ƒ�U8r(5+t5\�$�h�$
���nT)݅��b���8u��@t����5�������aʑͪ���7n��{˔�h� Γ�#�@)�����3{E
��-Y�8\�WJ��VE������	�0Zٝ�^3;�O�D�����I]2@Y�s��5f��n)���?	�r]wy�v�/L�:���n<�ׂ�E��[ک�g���r��y��d4n ;:�e'�kz��S��׬�-���hW��V�}K������b���k��E|�7��u㫻� ��G^誏tu���u�m���x��U����"� !��
�q���gU����M!�݀���Y{�]a�/U�"�V�م�K�tA,\�Fy#|�R)K�!�q<f��W1�:� �Ue�Õ;B�n��-�ƫ%#n�G�����_^�aSJ,�������Z&��g,J�s��';Sx�-�,Sl�k�A��+@�$��M:���컬��V�p;tJR����PFM5dԚ��x��-wZ�p���C���k����G�dB���}��u�;��Y�0��+�>��X7b���nu� ��Q���KKz��ŊL�v��.\#�#f膮�e�g�<ӵb��-͓�]���cZP�*�Y��G%�i8���x7��NE�z�d-�ß��i}1|Zek�,ɖY�f½;��(��s\� Rj�H2�G匋�n 
q��"��P@
�"*2 +  H��T��� ,��TJ�� 2 ��"��P*
�� H��A 
��"*�� � �T@� �(@B�����7vm;��vM����[k�D+ZCVV�$QQ��ȁʚ�4��)�GCzv�[����X�u����{���.>�ݛ)�G\�Vr'=:g��A��Nh�ì�����K���:r���5Ǿ�:���|5n���ٛ�7gq�N\B�y���̀��v���2CmS�ɹ�J�Ȩ����_�����;�/Z�u`�}	�A�o�g��O� �qz%�v����Y���׀��}�ݛ����0�T������>� ��{�;�F��uy<���P��ǅ(q=͗r��F�?��*���(ȚK������Wl
�C�vj�а,<�v��xX�DZ_��O!��{0��j�g�64bc��X[���*S��R�"`Z!aŜt��hG��@��W��y�9��\�}w��C����yxޏY�������`F,����dO�{����I�U����Iv�5��n���0�ž�:��3gq���b����E�z����wU-��3��n���F�i;n����'r\�^ן��ñt-�%gh^�+t�,zl��i��&l['M+wN�u��#�g2M���[��#'(�&فZP�7j��8٪��9z	2����l���]�nW|�kb�]���7�^���[�~fv���Gn���%睔��c#.wt�D'dҸ�X��Ւ#6^�%�%�&f/6�U�AoA����=RkyA�<�"�xXh���^����6p`.����9}����β��k*�M���$��n���}ef�v"�2�LE)�P
�gt/P4Խќ)��`>9�w��O4�?d�7��p��/3;��
���/n�:^�W��j�-�|(6�3�S�����n�>��O��B��-��G>�L�O��7��n�����k[͢��[�';���>H��X~����<{���T؀�$�d��ݥY���KxVڦ�Ui�+;���]�t���"��n�w���m
����Nʼ�?KI�2�3��]as�c˷V�S7�"ꁓ�vK�R����)���ea@����UN����2��X�&n3��R����б�q38!�zeU<ֵ]x��z1��I�9�N����6_jy�	�οz@���&���=�2�g��]�{O���=�wy[�n���a�B��,�N�^�>�Z��f�ɺ��Ƶ��������Bݪ�q����jč�zoB�1DAZ]]D�^H�ȧ�S;��_6��7}�����gym�wd�U6$��˫��m8�w���~��-��������f��
����t����6��&k�;���Ks6ч�P���� ��e^��}��4E��Vh��]ۗ��V��);~�-�Z���,��.n̫4`fn�s�w�N�^ۜw;`˶s�Y��xo����T��}}�� ��yӪ�f"ow�;7��Z:yd�]%P�c�C��Qw��wx��+I��#��p���Β�D�|��|��fy��]����ފ��蟻�U��&��ѻ@��+r4�f"N�/b�ٝ
6m��y�}n[� 3TK����ܼF��U�#��V?v�V��`gk7��
P	�{��<�h��c�F����&L��{F��^[�����U�p�ZΨ��)q��|x�����{Ϟ�����Cc/p��=����;�-���x� ����א΍��̻��}�uk�����_W����՞�5o{ai���]Ώ)�U�����A&��8f��v������m����D�`�Af̋�24��T-�s�^F���nl��/zUާ�b���y�I�2�B��KcX�Q((:�^5�'q���Y��k�i4ɻJ����Fi��Y</V��mX��/;�Ǣ��:x�5.c�"��{��z��%]q/�7N�����E��r9��F N]H�=�	۽$�}��o���{:���5V���/��O~Eq޻,� ׭�<��K>�{Y�48q��ŗ;�^ )}�.����L�f�%J�ֹ/s����P����C&�p����o��|��/�.7�9o�4v��Olp���n���x�V�;������;�1��ԀE>j�칃�9�/Gf�H�
]2n��AM�-x�A��,�(|���e�GAo�H�Gp����ǦY7X��z����P�$��D�������w������_����J�JEf��h��ؑt�Q4ն�4��f�TUζ͈���Ha�����AbZ��ҮpU��9�K��f\��,ZL���`av[�hjJ2��Fj1��[[�A-�h�F�$��!*9�me�Űn�X1[f�0,��7WQ��^;C���Q6��;C�f�lʎ0��+���ֳIcae%jf��r�X��K�-�9�mKl�h�8ΰR���!�\��X4\�ٖ���]��ٰ�\֑e�VUͭ�.�P� L�Y����h�����.Y\�j�9�u�
Fhc(��"��,!P܌�,ԥ�l8��9�cV�(h��&6�� �,��88�ʊ�,�FKa�H�.���-6B�c4��,3M��.�(����mk\��u��(n,��NX����L8��%ٛ�+y^rr��D[�]�
\�gR5�,tu��k!e�n&Y0��$.��-�rk�V�QZ�B쮹]��L��*$7+x��8׭�eLX$�����*��1�]�ɥ�ofR��m��u���V�-��������ѼS<MUfi��b�@5\��D,2��6&��s	�����WB��7Z\]��m°�[�@�lek�c5Mp��+kF�f��0�	Yc����C@h�B6։\�M��0�sUu���q8`��;Pn�Z�Xl�-r�pӭbd�r��v�\a��"�$��4�)G��b#�-�Ns�!��Q��f����vSJ���vԫZ6�
i9���sPCK�7
hٗJ�j3K��SgR�E�	L@�r�s:�.�Ĳ�J��v�:��i�p�.H��{B��/j{idd� \J��2�k���.1qI����sK-֙Jb�P� �Gemѵ���u�
�DRVhp�zǋM*����hj���,6�.b\X�]�����%��ld���k3.�M�TB�Jk�Q�� 5ck�QHX�^�n�a�����d�V�dTq�������ni��\�ɔ���[m&���L$4*��TcuP,�P��k��h�p�F��Jcg�ᔠ�%s��=�4Ŷ�C#�Ƴn�h5���V�d��s0��&v�0ؐW�T�u�A�4�X.��m������`��:b�m4�5nŎ�j�jE�-#Ú��2S0�͖�.&X������-�Uб���8�`�Me���ʹ�x�*t�5��l.0��\�5���V4�k�VZWZV\�6�V�����*Gs3����X�kB��)i�r:�/Z�ܱ&4�`˻rܛh�l�Cn5ں�����)/ۍ,�����,Q��+y���j����(J�aU UUUUT]��YU�
�TD�-Z��QB1�c���K��2�p/3f����m��,Z�:���X̍�k�̭�Иf�2�\03�tw8&1���	�1uɴ��#s.1�
�5��ʬ�lYb�б��T�#)�Q��XFƆ6`jSћ�֥�6��\�41k��Z�"fh3���w�,���f����H��#lm�����LbF�Jƣ�
r,V�@,�T�Z��d�dQԪ�VҮ%E���7weh(+��Uj�Ւ�e%ܱV��#.T�1���d"#D�"�J�ڒdƖ�"|T��~��{��`�#١b6l�M
��Y��-�B��˹	J�!Mf*��D���]��	Y��\JMSl����p��e�n���b�g]e7�1�&F�ŋ���9k�d��af��Y�0
���ev�ZV`�`̣�3�)��$��r�X3��Z���m�K-��\��s��5G	�S#��ͳ)`���5MBQ��4t�n���l�5�a̬���*�&ć2�+\��)F	F��B��L�p��R��r��&�AU@Z�����\�bie�e��j���ҭ�9j��xq	ӥ�ҙ�[�^eZ�z�ޠ�)x"F<*�m��[c#[
ȷ�X��VTB�h�#�"Q)g�c�g��o��zz#�l�)�$m����^k�o�w�Z��G/ג��ҎQ� �dsݡ������?}g�L^�x纘 #@�hş|�7�Eן}37���R�j�5HwȮ�Y�*��B������緻5��L
�PD�F�n&6�Q�!5��[T��1M�7�|��U�v5�SP<�?h'��Ӭ�yř*��#�|b���)��|L��mE쀛Og/N�)�s�ٳ7�o͟:ZW�q.�t��k��ʸ�$��u�)h>u߾�/��me�p����`e pl��c4og�]wÆrV�w���o����byد�%�:x�0gmú
�E�<�Dc��c�&63@6}R����3��<�9��_�Լ���\`���a!��!��o�"��q���ߗ��}�SHNûa�Ӵ�d��3-ҋ�;25�6�=�߽�i���^h��8�r. ,�#7�����0cф
t31��;⎿�_��ǡ�2Oz1ض��<����sYy�<Ut���y��"�rA�����].f5��6+�[���SC#� :F���A�;�8����m����&grTz�_k�i^!�	���y��{z���Z���H�'��|ə�ƶ���`���+m\|�'��+$j��ü�����&��T:h����9Ѭt�-�G����0��2,��̦�� ^a	
�a]i���4i���%m����ò��T�]E�u����y�im�t����#�׵//O��q۱��9*<���Ӛ�f��At�<��&�:k���D)7Z�t �� �ߦ�#(毓���DԪ�B a�ǔd�zV��|v-,��Rl�/^���o���t�j�t֚�{���u8�����z���~�����@�##<g���!�/��z��ҎQ�G�Ucf ��s��u�Ș`FnW�yE���q�����	��lP���P!0L,�G0a��=�|���g�k:�^�ƭu"wޚ�t�&�[Zw �<�(��ؒ�(���]���Bd,nll�t����Ga����GA�2yiF&NK��?U����X[�3��9��Τ�Ϡn�=�F�x�o�P(0��h(����}�_o:��S﹭q�/$y�߯6b��(��#�Q���Mm3z��Nn�q"hj9 �}�)9wܰ��f����E�7{�Z;а<�}MkȂ�D���ណ�淒�Ρm}�5��j}�����Pn*m�����΃�8��E�ݝ���><n�Ե��x��c�=�γ/���$Q����ZS%{ޙ��v�񊮚�}��5{���o}����fP߯�|�����VB�L��J�"�-�<��b��H�����alZKQN�^�n��]mc�v@ ���wj������Tk���f�b��lb��.��/��5��OK�b�)�ksٮ;M�&�;i�\�1#���f[�N1��<�2����SHy���рsR�|,�r�צf'Z�z�2gG�b1nhu���]�@ "7RKAf����M�Y1>�>�I��'��)��_l���e-�6�?]�n�Ҋ53�y8/�3�7���h�X�EoͿs�֝I\H��y35�Ӧ��N!7=�یh(ϊx�A�h���Q��ͻ���JҌw�)�a���m�)�^n���]1׵�Wt�*���3{�{w{k�^�Wo,ݲ{{�K���KK_�l{�<7g����n.{�;�UX�+�+���4(������Awt�͔�U�Tn�;|��"(���ٞQh�Y�!@�bNn����U����z�f[��9���m���H��<r�=�sAlٝ�8�D)�źM�����$,��'��;34�ь�U��ַ�MH�r�-^��Q���ǳ�X�ٕb��T/���l�ڦ��f��\���^[�N��	*���g(��l�mN:��ji����w������$�_�ƿ	�D`2Txڢ6����R�F�ڻ�	*1���c�"2 �h[+H�Z'�h�)x�	͋VF*FP�iV�0$H�E���"FBI ��$H4�*�ձH��##$cMəudeFA^�� �au-��"C���1����[�2X\UD�$��T���m�Ɏ�eG�TQ��Ji�ܑ��j����
ǩ,�	 �^D���+�||c����?�!V}p��^�?\y��S���
����te�}�tf�贈��fʬ$P�{����8��b�S@�L�2��6N�mGRV�}��r�z��s�"�Z}���:�N����yg_CZΤj=kI�\���B��W����v2� ��[9�{;�ۦ���w>J�[L��f�K�h2IE�!
!'��	t{�`�1mG���{��^on�����V��6��LW���c��Q�Q��=��H�#~�i75�3���@� �fi�ϢW2��֠�I�xލ&;Ci���xk�nr<��]�[�o�X�U``�=�t�9�
,q��h��8���"��b颴ka��*���m����ѣ��`�h�1���4#[�̷UqQM�eH�����Bx���"WӒ2=���-���9WrA*=Oܪ��<����D��Ϲ��'Z�د����D�zƶ�Lk=8ֲV����5׊�'�k�0�rvnvw�ԋ>%ż�	-���\������� �$G�v�7Ψ�1P��u�Z�v��\\e���ٌ�t��06@�Ɵ��ڌ��ޯ�8mEv�׾^h����+���<I�n�͚O����<b�1����x��ċ�Nw�}z����e���^{����{7>٪I����>�{R��� �ky�[M&�a��O9p
hT��,m�5J�,kRԏ�;���M�GՆܐ]5���Яz���ltƺ�0�o���Jv��5�޴ic�bA
�������OS֣�Ot�ޥ;�~ߵy��ek�/�F����3������!i�~��w���3�����F��f_�>9����oC�V���:�]l���6<��o3y�tf�B��G m���ɝ�ي˫r:І1��y���o�^ugu��q�m]��7��뷆�o-4�cVO�]^b��.��75g�C�ӟB�1��k>����=�v��P�4w��Dhu�|�11����=�!��"�U��[��㧅�Z���A#r�o��ፅtS�V�� @��j�H�p[e�G��kF5%s4�ʄc�qWK�Z6�C�Տ.*,�(iX:�`P(0�иj(���^x/��^t�}*b�$��>�7�͘׾��3w���/Һ���3���u�7��۴��Nِcno� �}
R�n?���2�ͤ��z`�^JM��y���3�J i�@�b4!cfAA?�M8��fw7���5���*?C&Ѳ�S�A���y�1�g~��{X
����'_n�CV��fbz�C�k���=����tƼ���QrD��=��֥�ﷇͱ�$��|�oU�h��nSs����G�E����u�pYF�+��p��u���d�{B��]�
 �����v�����Q4�٭8J\��w����}�O�>>kGW���h���+e�.���~���F/۳��5iIw�-]Co��17�/S;��7i��%��o>
���ݎ��.ʱW\k�y����d�p`T���wOJMi���{\m�5;*?3�	��>��]$Ns[�����'_�/�}��Zi8�"��!��gL�E��V�����":�^�B�~χn��Ҝf|1w5����E����4`�a�p	m�)�a�����@��&v�����Dԍ���k�l�
������{u�s���8���^�;�j�Ci���F
�!��f�k�ƛ��{���@��ɒ#�T��z�-l�0��!SN�گ�����μQ����Rr���X�7�^��ʽ:V���Ⱥ�G XPw��C�}���o>�|Y�ӳ��4O"��˼���x�t~�EG�u����6�F��.`~��?x�u�|�}���c�.��F�v�ל����Y�-��%�����A0{��#9Yٱg>����p��o;���S�H�+�����jgo�V�h^����&W�v̏'�!��c�p�R�%�&�r�߶Bp;��E?��yr���E�Q�^,�-��%H[� ���*mmaM�ٮ%-���%�IlcThJ�CU[0-�-�Mv��2J��lbd��a�, 0�H����D�5%Ŭ�Fءl�[��҈�*^�Yl!Ju���	e�Z����#m�����[����=�Z!,����^����&��pKHC�e!�-���KA	`x;`�,�����;�3kPcjL1��7KT&6r0�#0�R�J��,1R�\�Y��;n�&�jD�A���ո�&{7R��[6��讅cH���h̪�j *�<]Mq�v�Z*[����{]�֬c���	0�1�ƺ��X��,�$�F�8�, �^@v� �n�f��.U�X�n]6a�WA�[���P�·�s`�%bR�\��)�VėEɍ�X���6"�]�aL�0JP�MlK.�uB�X���a�ík����&f�U�٣�t��h��ܮ��1^a��mZ�x��&�����]��vʖ7��5��iNyHk�jf8Ֆ[uy�m��+*�t
�Q��~�_֔Vc@����`&v������U�WJ��P�����^���,U~c�
c����y�7����d��;Ut�Wi���߷y����f���w ���B�Z^0ǔ	�B옏:�6�8��n��.<���)��W����vX�@t4��������<�����=��s�S���/���.�o��݄������T�hW��� }G� ��6���/�Z�Z���z%�ھ��77���#`0��Q+�ZMB�w�s�m��E܏�9;�4]�-�奋����}����>]y�:5-�]��o3fH���*�H'��|���=3F5��^W^67�����;!�%7a��{w?{��V�~$�9����N~��Z�rF�/�~lӦ����޾v�᭭��tԫ�������ˍh�M�X�2={׾����C�6S�LQ ��<��`ą#j��${=��+����-��;�tLi��7�xc�٘cĂi��}�1��B��b�#���l�F�����~$u����C־Msͅ�k{r���C����[Y��`�Π�orn�q0 C&=(����j���{�{.��&���z���N$�i�Z����l�ۤ�ύO�>���P�#�O�y��5��{��J�>��lƢ \	�C#� X}]ŽIA� �鎝ݡ.3��Iw�����=�qR4$K�SvfȚ��Y������[Nܰ�%ͨ�n&n[���j���ґn�F0�63(l[VYXD҆�����Lz���d�*<h�{�75���屑^�0��4�U�e�Yǭc]w�{�M�Ԋ�'��κyN�d& ީ8r��F�M˄}'_MY�hKj�����%�129�ݗ.\��>�|bO"rO�i�܏�q��q?���;�����qs�5���y���{��?$�P��w�B�j�sq�H������;``dǶ�͒������.<�eȪ#��ۛ�I;��֌>H+ă��3�^�O.
�vW �{��E/�X����ɣR���dƩ�.�y�(C�bx�!�{\y�۞��O���*�Ft� �&53��C;]r�;��D�L���� ~�2<x�
��M���g���0#H0#3���ڒ��81�[:��G����VPc\"� ���M�� ff��9�"& �� ��֛P&jYa�^q��Nkn5$D�x�F�!v�����T��V�n��*r9������}���05\DU,�,���4�D��^��|������������?��Υ��&��w�u�pYH�ҍ�G��O|�O,-<�b�!���n{4bk�ݼUz�\S�o��/�����$�^�.�X��G$k���3e���u5ӐwY�4n�ze�sqN�u3�ޣ��魵��;���6T�{�<�ۯ��(��o4�$����X�5�+5��d���`��Ei��Ҝ6ݺ¤"a��m���������3e1*<���a�,��͎���b���/^w�{��nj�A�R社~����J9�(�����2C�`9=�!��r&<;Z�8�}p�����^���DG@0#H��֝��|��l�أ��u�&�ue��T�z "l7	�Kh��N{x�p5<��U5%<=��&���oS3]N?�}�̈����piU���E���Jx~xx��u���)Ȝ�LϿd����1�_�_w�^��М�S���r�l�zx$C��oH���R�5���כ1"P���%
|�����ecGZ#D��(R��imU��(S�	d��>�v�Ú}K��I��T2��s��<|�~cF��J,��@�D�m��B�@�B����4vJ�J�J�?o97y�"P��(Z�x�mIB�)B�č�%
P��"P�(�ﯼ��p>�B�)�߾���@�"P��U�4�� xDxG� ^_F�u�iS���9$��0�ݢ*�O�G���oLv���K4�n]�ME�=�=�����/��x#e��x�Y��\�΍�y5E�����<x�E�@��;����p�v��B����y����&����x�灃�(�tI�˟2M��'Mmnf@*�}��"�4q-���{bw��5�T��C�jFc!-v����2�cBӚ,ۯ���8�Y��� ��=�%�m%\��OX�%R���P%�ƴ�o]L|�>K��/R�4:[)ր�x�	o[}e𦭚��V�2���g��u�����Eb���o[��i�I���,nj�P� ��!�R�m�,���^��D$ay��)�䄭��$�P�7�^S��ҩB2�R�rԍFJ�
(l�  ?d(R�+���҅��j%
m Y�}�ٍܼ������i(R��ԉB�)B���
Zj&�P��auX����4[Dh޿����J�J��F��B�k[����
�����B�@�Cd(�IB�)���3���K��n7�/=��~�����J�U��-�'��R�+<���&�҅(Z�j&%ZZ����Ѵ�h�(R�]��9��D�J�I�҅-4}%
P�
絁��G#D����n�4m�'�(R����J�@՜����Z1��J!!�J�hܔ)B��߷34�:�;� ��J�X�hD��-����"P�HG�8���.�y�9�kI��ٜm���=��s���UU5֫�5�<�9���y�����)Gd(���B�&��:� D��-D˔)B�(H�-��S�ym�Y���0��r]�����6�)�?!iB�-����j%
�cA�o���K@�B�-%��'߿g�4&Ҵ��)Bָe�bu!���-Wt-��I�(Z�'eZq ~��ɚ6�|ƍIB�)B��D�q��h"n���}{�B�-%
P�
R%G���Ti(S�o_hNM�)B��5�(P6�(ZbQ$:�����
�h�(^�7��ə�6��B�Z��j�i!��*҅��P�
P�q#UƣU�Tj'�@}/f3�˾�>U�F���l�s;���ɽ'�?�QTr�7�0X%����YMJv�Ֆ�Yb�M��n�e���l�&"c%�p [��Ivf�M�un3���b��p[�$�L@�i��^s�{�y�ġh��bP�@4�(R�(S��)1�[V��B�)B����'�{�nf��P��"P�_�?ei��P�_5���(R�6��p�J�7r����Ͽgך1"P���%
|��(Z3]��s9BѦ���H�[Q��D�M%ZZ���fh�P�d��w�_�o�B�("P�h#�pJ���(Z����ʭ!Ĩ���B�gu���Ѥ�N��-*!���(Z����@�D	�ZP�ġN D��Q9%
P�?�=����mb8�(�����2�hH��#Q��F�&�"%D�h�)B���Z5[j5Q��)īK@���m�ىB��(R��G�{�-�9�]�l5��U:f�}<}�|��}��@�i"P�
P��"P�G"P�
���Mƈ�5Ͽ}s7G�4���J���V�)B��5��Ѵ�J�L@�(Z6������h@�*Mwٳ�pI�dD����VV5V5�8�ihϾ��J�!���HP�y"P��L������Pq(S�(R���(R�%G5�O��"dl˹�Yyv��w��z�4~h���b(Z>Kj҅(P6���4{߳IB� p�P�G�(S5��fh�|�: D�k��̪Si��J�h��[E�D�!�m-(Z�j5[=ˬH�?s{�y����(�@4�([j�O���f�3���f�;=?;W$��S�Y�h�g\~x{� �=��?g�q���3Nڍ�=�Nf�r�$Fw�SJ�ȨDY`	��RѹE��5ff%
a�<�>F�e�Y7!z�j�{�陇]��!ֱMȢ��~���-�@
.o�ez�,��c�и���6Di>�Q���j�l�"db-�8���=dfVeX����<<h�����'ٽ��\b�z߶uk���w3��:��������� �����ːkO��ɚ1��}���?0N5���}5�u��T��y�Kjd�׽������):�Groۊ^qT�䦅�
���^��$��f��lFC��6���,�����7���&�z�ȫ3sm�f,��V�n�K��9��-�d+4�a%��h4�;Pz�a��yJ�f[��4�͈��6L�m���A��1�.+duʌ�b�Z��|n�%ǦH"d�s�4c��߹>�Fײ�����2b���z���Ǎ�Jnr2<�fi�_�� \mP�Le�R��1�Q	�$Ӝ��8�q�S�-�Dk��"D�qfΣ7&��.X���~�PP{o�Ȣ�k��}��������_$9�}���uNB-?I�f��я'-KIH�r��L����0�\K��cƣ�+�}�g�}~G�[I�ق���u7��8����H֤}����kڝM�T����w����u�1b�"a#1�)-�Vr#���P/`A��+>��m��������ռAx�*�Ɩ�������Q�L��!o�Y�Y�)��ı"�:U�6E��}۫� ���\Ab��7�5;�zN&�8��  �D�,��e42Dp�\���Y끷 �]϶2��݉Qк�lIXЛ�Q=M\��,��xx{|c�Ws�4�L&j>0�^��ή��oo��&��ٺ$"�*�33���ם�"��N'&#���^��va8��I��;!\�����}�L�Sz�WmJv�>�K�8�޳���ES��ܟCi�[�I��71dNEǮ��w�8:���@�z����:!<�S�3RVd��0Z��-x����[Ń�߽��E\䢃U����yA�{W�^��Ť/7�	�Ħ!�4��I�}Z���"o��� @Y���A�ףs����5�7+����T����vt������e��T�r�[�3)P�)M�'��:)�JB��'-�Ν7./-$nǮ��Y�gڐ��F�>�p�����㝺��b��rE$ʺ�R��'U~�� Kn��iDQ��-6�JTY�Ky!q)J
XY)C�,��-�2�A���Ai�ƥ�EDI.�@ZnR�5�,���ZD �FI1Dz^�4��yMy��oP��*��"�(����uij[,Բ�l,(��kz��ʊ-�F������TLj+y���ej7\Wa�Ҋ��ѿG�e[�,�ͥ/:kVV�M2�8滈6Y3˴Z���ƚ�:U%���Ym�Z[c�,!�Ř��FL����� ^769���1��f���1� �J-і,!��G��QQ��&�8�L68�-��Ɨlƌ�t`��\��R4� �ʆq cUY���B��+�s��릈X���r�\Te�cp�Y�.W��̶a�H�U��F,��/6ȴ���*+�k���[�ή�������3��&֥�6����UU��T�)Qp��VVX��-��8�cPR�$�b5�˻c��;��o`(YQ#ct,5��D�M[�SW�"�VmpM���ҥ�lh�Q��$�Q�㣑�@���΃�bk5�*YK����=��([}{2<�n'/Hŋ!I��)-�,��������~�Уx>|N���9F��ҟ4A����뫑��Zv��	n�m�Z�a<��y����PH��������Y�g�#LL�{?Ȑ�VQ4p�F�E���{���U���fI���[[�Ot|����٬���)�ʤ����]k���	�C�b9AD6��Aa�aA-�oiN_8�]��q�����R�M�|=�_�T��������͢.AȈ�jNS1kJ�j�>���#k�}�Wɫ��c��	��6�N�V3��)�s1�a\z������L4�)&ل�N�{S[�P&�� �k�
z���	=S�8lCg �{s���K��s����M����*,N�\�Ω!QFV��<=��*�5��S�/�zn�`RwP����a�a��P�ϯ��'��웺
���MN�����b���)�h�n��2�sރo�bt��U[z�TCܪ�ɹ\g03-]p:q� w߃�v�'�+�94x�ω�w��:u�|O?U�ctķK$�0jf��9�7k��ѭ�KTf��6�X�a�Z��p�݉��8m�CS��@F `�
�"�v�'����d��ŧ1d[���ݱ/z�[Zτ����k��ߗ�iU.A�����Z�6��Q"���Ǻ���7	4�2�i�QM�v�}0����׻^Z}ֻ�՘F�8��89G�Q1捯���b�lr�[�S���ֲ+Y^�.�oҚə�3�NT���9ٲ�얍YRf�c�HJ��i��33�}�~vU}�sk*p���rSr);n�A�2�r�N]���*���
TC4�	_1�y��s_�w_
�[������V�38UHuRk(c�;½��2�wf9R�(PXA��H�q	4�{8�����]E���;�׆ ��C�;�r��d.8>�O��)��s&����rt]�	�3{S*\d�t`˜4� R���(_l�c���j���'��[
P�e0�0Y��Wݩ�����cN���:�)�ڛ��TFnc�8��^zz+H�7}5�74�2	bc��'AY�>'�����/(���80��ٺWXR��m|=�w#KDAH%�,B��fYb�l�l��;2���}<n�:eV�)n�P�-uڴ��Z&����h쬱��+�4a��b�C���G�8�>�ݗ�Q���yҚ�5yfY��˩�tS��
�&H�z8��k�i����:)^�fnn4����y�f;h���N��f萂�_}�Gw����g��ec���swI��G����rBw"�'t�}��o�QW�zl\��MVg�w�
����h�o�6ox�t��r�4���}7 ��}��O��@�i�,��}��|����Y���'+�勳�6�9�ު$�_q�����ur�%�9u�����w'O�z�� ��ף��@��3�5{���t��-5�y���o�s.�������zwb��~w�뛗ѱ��>���|o����R��x���yK=��o�������'$��o&��ܣ{�+�S�}�L�)���Ԙ=�N�媰�rw��1���}$�潣�p��#�mz G���Z�wv %_M�q�1k�&.�ټ �XG�j$j&3L춷AP�����#�9�xy+�ZȤcC�B�LcI+��ǲT��e���mx&K0
"eeت�#J�*f\̸�1DQ�)��d��.,��w.�J��#��ld�RE�q �V�j�]��--UV���QDT���$*�I�FX��~{�v�ۊvZ����}��đzd勿�7E;.Sg��ϵ���t��u����#vJj�k�}ȇ��P�"��'�7қ�|p- NpN�+��\��
zw%]�]rS���a�$d	����ƹ��["v2&��N-ltO,Թ$W�S����]\�T�L��7�|�w߽}�%����پ���r�:�V��<�q����2@"�n��4��1�f_�2���L��^��n�s^ޮ�)��w���H��NR㛂�F��變#o�#�ZS����/ҧ�� �J�i�e�Vٹ�ԵK�VC6���g�����i^ҕ�v�8�m��Ba�6�Ə�U���:�Q�&
I�JI���|���j��K���Z��Dr����R2�q�>�Cìރl����I'�<��ꈽ�ʳ�� �cr��eJ�hDKPbAA�Xh&�4�4�'����j3�;Ԛ��G����������;�̩��s� ��ӈ;���5C4����"���M����j���B���JnV5tjQ.�	D1)�
T"�oo'ˎ�]w�s3[)��l�	�Z��f+�MU������oC���W ����S��k!��&f�	՟���1��N��JB�^��3	��}�Q��m�Ʊ�3}�g���l��MDL��n�{�f���z��Բjyjg.��'0�gtmiPv��!���>��Q}I�7��6�e��{�S�/؉�m'������^|���"k'�z�8��;��X�BL$	�� �a��B�������C��*��3ff�S�Ne�
Fa����%���n�^p�c�>���&,���n*��E� ��䦫 k��z�Eu���;�!a��M��q�Bc�nj���ѣ�
I�3�"��6&�-�cA�Cl;��B�j����җ%Z���a�6�d5�`�#���IDP�V�0���A��}���lnbqh�N�2�a����'*�Zn�)�]�U���9�&�VȎ��@�\���V*&fZ���@d��-�ق�껹5�mV�1�O���N��p&�;9��B*�E�7��Y�����vw����C㯊��y���j릹�e�����Y���}��.+l�Gk�������������[�����9�ړ��H�ʬx͐���]Cd�o4�H�K�_M��$���`��cl���V�!��c��>��Z��+�wp5�8ۜW�/����FfMf�s0�̍��]ۑ���. [a&�)���L����\\���ŝ�_����K�>柡E���ro���n����/jS^�rD�]О�T.qBӘ���^�u�k(�..�)����u�"�-͐s0h]N,�H��B�X1П�������w�]b�����-�rr�U��:\Ԝ�Z�bi`�F���Ԛ��ϧ���q�J�1t��$��V�S����r�F�p�g��t������ޯ{��.�K�{WL3�nH6�;�x?݄Z���}� g=a�^kF{�{@�k9Q��
	�%qTR�"�XSc\�� r��i^����;���S�ȱ�U��ָ�>m_	����Ƕg^����F�L
C�o�g(�sE�����9��܌Y;1�!�E,
� �1�^��u�9*��n>�P�a��T��� F�§1�2�B�E�s"���}� �P>b����)�ri�)h��,Ir�""����WCM�QK���*�22�(�[��"��-��]�TKq����R �˻���JEUB5�Y!�&5�QT�20���*5i"0�H�����e3���m�,]��Ё�+����X�ԳP�Z����1�3u"�m1jJ�PɁs6y��H�I��h�[�Q��~Kk�b�V�f0ɮh*���͢�\�q�B�=p9XP�a&�eMJX�ŧ[���zҺ�pJ]�XX��1q�!41�4`i���t���d�Jehַ7MA�,�%JklKe!lr�+eiyZ@�.^4Ͱ[�Z���cL�-]�7�).���J�)F�ه�i�V2����l��%(2��rڜ��ibE�qaj����f[�T[��k��ͫ���29)x;b�T��7F�t��1��ؿ?B{��[s�[,4,�i���\A\5�&	V�,�6��j�@��Llhf�Ё��.���R��I��8f0��e�S*�5�T5�{����=*�� L�L��\e��
uWBd��Sc1Wt�L�t,=V�k1	�ғ�7����6MQY�I��h��ɺ��nо޷�ԅ0�
�Z�a���x�/��V���.m�"j/]7ԪI��;	�t.�+��»��y��ZbW7���j�ۨ'�牜ا~��˓�(�ȕ�~�_��mX�ǃ+�H�	7�%�Ӝ����2+*�V^.|�]'d��*�������G#<��[=׸��Ꭲ"p�uel��S�"w_���2j>��]ŘF]B����r�N���~dL^���&Z��#	�&	�>��I��g�\�vE�]�I��5��T��9
��}z���`�p�[7^�v[�}JN�C�a�H�Bɴ" �c3��[������E�Ѝ�=��w�t�����Γp.�P���Ca���B
�S���3��:�s���̔ǌ���2 s��(����;��.=vm��N��=�ꢽ./}�9M�������_:�������)G!59B&d�q���ᢪ����Z�AkZ�*+c4X�ba`0k���R���ܣ�:[�\Fܖ�e�J��Df0�� 
`\
�i`��5	�����ͮ�2/@�;|�3�����Y|0�Z��������+ܻ+�i59|q��6�4*G=�)��-������w�av�7d�Y�,���!����ڦ�occkt�Ξ�Τk;�P�i��sø�og�o��:�_燧~iq9f{�z����m�W(N��'1f�)�fۧ�Қ�������U�;�,ӄ�AhCP�0S0Rm�v�O_8d�UO��5�T�}������r2�2[��ܭ�yov��ǔ�@���!0��ؘ��}y��r��]#��L#�fWW���7l���e�Y�%���+�u��޽�O�O~�� �h�鴝�$���Gm��m�8j�+�.�Mq�3*��;"V��(�I��9��U>�e�U��2�n�}��2nq�gv��P����'�e_۫U��1��E=~{��;>��_z�3
��MOD�5,�,"�"���7gJ~�>�\[�,B�r��T麅!�]s���-�(u�f�cx���
��,ނ*e[x �c`�a-B�9R�2�q[�v%����TXgm0ch��6�Vm#��f�G4V�;�b�j]re!�L��t����d\t]�q|�$�Ud%��9H��N��'+o%5��0�V�Ò5��N�)���d�Q+��zh=1q���.���h�"@��0"���va�ޘ�ôE�����:��vO�vм/��e¹�����[��7��_������ɚ���Nb���ݸvn����$��>���痷H�ɴ��w[��a�󘵤m��f	��)��j��lr�ܞ?e*"�7�[�Sؙ�$TF݋��8� �޽�<����V�f}�*$ƭ�#4^o��S���.���}���n���^�(��37�iT�A�k�j�"P{��w/M����bZ�uU��+u1�j~C@�'�d���8�{���}���":S�ڶ���C!]b�����ا�ė�>��8������U|]^w�-��7��T��gcC���2�}���f���\g[~;�Sthw@">�[�ޝ{�׏x�\�2f� 
�^�EK�w`�a�V��M��2H��BP�D�\�IH�F�X����t��[e"���S$"Ƒ�DE.F�.�,jMŨ�M�ZX5m�\���K�PZR��"�EF\l")JL.�2�+p�E��~>���_v� fHZO��gҚ��b�.9�^��l�>���<fņm��Lk��۩9|ǅlTIt�ywZ��G2��w<�\���k�y�L�\��}��N��I>�k|D��	�������э�u  /ﻞ�U��.�f��ө��!&e5���i�}���\�3L�鴞9�@� L���>���C��Y� M���V�^�"p�lv�2��k���t�n�]^{6>��G��%�7E~@���w���r~rNNO���:�aB�ʖb lko-��%b+�6�1����^hT��eZL��J�e�a3��2#�[D�ZSW6�6V�Q�c������Y��x�լ7d]��2։�m�o���H�>�I�Q��D�!v@��9[�GsP�@QTV�<��^f�n|��f��!EUU<�	DC�~%*N��5���\�`]��k��E�Om:����a��:���jxE}�ScmD�Q���,�ǳ���8�'sNix��֭���g�K�.�t'$���2��I)jAa`��5	��o�m=u
��y�8��צ6�rF�\Ă����캽�1Bc9��۝:����s���>�[|e��ܬm�;Gl��fL�]����郑��O��b�*E�4���S�D��$33]����6%�$)==f\�[[^�>��̯9��kjp��*<z�&��Rr�o<qv�t����o׻}yzqԈ�0j��i_g"*�wq��e�O{b	aZ����0�o��R}�0*�RF��_d��TLyK�� λ�<���f��y���ؗ큷��1�c#[Oо����j�,FK��x}��߆�Dp�����Ko�o��w��AI!,`G5����ۉXF�,��0`��H�h\�K��D�����U�+
ge�@��3��uι{�����[>�������o�R|�lȬ��s/��+
���e<9�EQ�"��˗���(�zs�~�q�q�u�fL��qXoV��1�� ���y�;t�Z�N�vVwo;�Ц�KI�\�x�ܬm�ĭ�';FO�۔a�#�ω\�9�����^�|��������&�}u�{�@;���;<A���AAj�sQp�l��c�"��n�|����Ǫ���n��٦�f��6���A���Y0�:�C���_�e5=��%T��g���r�ϣ�Q�y��U�n���"t%6R	A-�F	Os��\�=��sun-�NWy!�dݕ�O���4��ì��V��Y]|i��G�a�������/ea����5��:�����3��.��Kk���D&��hÆ�(�[}^�N������S�[U�1�P����K�?{w=Gv��(�Q���7Ψ�|i���B�>�j��))�U]؊�g���P�=�����mn#�P�ns3+ph������n�YK5�zx��/GF��.��g/Q�3t�$��U0`:���lx����Y��iE林uϼ������K�#��s��η±�[rm�>��Z�w�ZSa^-z��<�X��w�9�j���4yZ���_ݻ7\��Ӹ�h�����]E`h�ltԑ��>�y�^��h�h!{]���h]�wOp�c������ �*i"*�H�(�pc"�[RK���6�ccQ�4D�#p#i-� �*Z-���*�U�j�R��]Jj�@DcZUG���ҍ"ܔ���H��T�A�TDq��bK��D�EPm��crqd�u����O��F�Ѻ���Q����cF4�t�+m�6�Y�X��5JM���l��T4��BhMuX��5��[q�kbd%�q,Jip�����f�h�`���IJ�����Bg��L�q�	�E��!LiB˩�1����Pܥ�`X�Y��KZ�0f��]�4��4
�u�L�Y��t�[sb�ţ61,`�3Gl�57i�y(U­�NY-V�Cm��f� �������)c���h�kej�B��4`	u��5��ֳ:�uiZ�$f[F4.�X�f"�U]���5t�1�b.��B���y8�Z�]+�&�Ie��.rBqa�uLX4r�Ĥ�%����ǆ7hn(\�6�pœU+K	ajںW��Q���*�Ƅ݊&�6�3 ��i�
0[���ީ"`V�5�Vs������N�93јFE��)��Q�.��$\�+y�8��s���`8��C���QbU89��ݶ�/���	X�$�(��&�Ok��}�1�	Ǐ5҇��~U���ߨ�_R�y�~*G����r��T-���/�ц�	�F��Gr۸��Ϯ�����L���=I弙�2'^��>�����D� �!�
a��L���ɡ\�&Dϛ[�e�qh��`�u#���͟�/@����ʪڎ� �cj�Hyie^���u9ʙ����vN]]E�A�OH�# fU[��!B[�
*	O�����粱�<v�R#O�B�ʼ����>�lK�<�Z���\�#ؾp���\,5]Up��]��^AAJ�v�k��4�M
��[Fσ�����CI��e�HL�e�;4��Ѫ�]��ι:f��kn�"jv���X�]i�ڮ6�ݑvV��nsm��oNh{w��$��ƫQ�بi��g��v�TbR���z�K	����C�|&Y����4�u�X�M���g��e�D�mf�]+�!,":���\Զv�Qj�c+��aF�� ��M.w�ϖ;��|��~'���������eˀr�/�s�# 5�mf��j��ǧ*��f�5".�&r*��u�F��� fH��S=�.�{'ƩmA �:�={�~#��Ͻ��@E���m9�#B�+s(��Pf:�2k�`�z�^�6鼅k+1�[�p��}�����2�WȽ�q�A�~�W��ł��~(�79n8�W"{��L�{���F)�v�ߞ��_�Ν'̧��`d��8ӑ�}�w tݐ�.��m�N�H�3V�덇�{"��	��'�(]tzn�9�;��=T6�te�+9�rt��۵@r8��:�\J&AM0�(�]�ɮ�>�k�T�Q[\i��&���%��F^7M;�3���~�"��aN��n�i�38wg79a}����pxgU�Ĳ��eM��yR����	ݢY���k��HS2鑸Q���������w�����zzgӢ�o7r�=�%����Ȫ��O�(��V2]O�gR�䯊stC�������gb�*�����q��(WfM�UK�-fVw�cpކ���Y��e�-R��[L�w����ZK3׶Y`�M�f��Dc\�!���n��V9��JV&q*͡6fj!7 �%=��O�Y��;�s�f�ٷC�W�ۤM��̵&����'X�n�}�ҝ�m�U�z]��*s�`^���ٸG"�l�H��a��4�__p��5i�pA%�ݭ�^�����E��n��N)l�����I��*��4��ۼ�8�� ��U$Q�\�����`�K5a��lKӖ�%��d����ޞ:���"�&5�߽w�>���1Z@�T�t��n��ӭ0��ӝY��U)�X|H޾��xD끵��������x�UΠ{J�9V-^^�.mʷ��Gw]���wh��N1�9i��\~�SwzӠ5��O�v�����6����0&g�pg�>�J���19�2��0nC��"�@���6d���n������s�r̸���xQn�gu��j;� �os���z�@a^^]ʫȓZ�[��B�$�y��\lƼs�)�B���}*a[9�z����6�t��블/E+�s6uE�"*�#qn�r���4"&H�I�@hED�ZD��\��L��հT$%*�j ���IiAAH��rZ��hTlH�(��lm�D�T�5$��Xd���K����5~�}�o���z�V��̺���Me{.�ٻOg�-%J��\���|�z�{۽8S���it�iۿ-bn�3�->�r�y����5�Tk��e��l�[��
%eμ�E��N��p��NU_Yt�8���rET�Y.ΊF"1��`���wۚ�;#Y�����J���뜵�No�7�_:��1���W�T��%ͽg-=��~���Qg���qn��*�Hݡ�C~��~�/��}���O���yJ,e��sXl�0�0@�.j�.�h�kfF���.J[4�ص���K���n�mV8�܃W8��٦\fX�[�]���}��}�ޯ5�6�5TWɬ�Y]�6:7N�{�e�����'�3���"�� ��'��?���My���)&���ej-&RM��!�	2�&����q�d�e�';��;�7�6M3�]Z]��u<^��m�8���8���l����2"�B�5K���X3O*���.�����i�n����30g���*
'�*?�0�����h�ާه�=[%��r*1�Ve��f�];.6w�r�3/�����r�:���ꯕpyW'.�D�xZ����ZWxp�4���B���7���Z��%�u~y�~�����Ӷ'0���m�=~����]u <>��WK�M�r8�i�9wp"*1�݌�R�^��8{}<DG@�p�\���W̗�nrU�Z�ۻU2[�oy��x���fҜh�V����ψ��8��2�(��F$�;�u����#	qQ�G�wM4�$�������z��'�����.��V��Y".�뫒�;��4$F@06J��p�����F�8E���oHN#H0.�gt�r�"�n��6�ƻ"��ܫR��-��6�A���k,-[���jK�a�˴ĸ
�ƺe�!N�Hd�5�e��dV�.�c��B4\����RJ&	�S��iS����8�Ѭ��0�/�LR e��f�Sp6\@�D(O�;mB����h�M�7>~��{+���v^aթwOa�z�v�ty�$6{\��on�+����hX��8�:�\i[h$�i7BN
m4����ڲ:"2=���t	��z=�U;��`�F�vzpJ���K��/�-�1�p�+��
�DA��3,>=ʛ��}����9�#c�=�%���q��7@�3@�b?�����*6 zD�B����2j2N�N	�t1h�]2�{ߞg�o�7^_>��P����؛X|nƝj���@�! �*��NhD������S��f1!�l�d���`bR!�J&j�R�ǸFI�o>��:�W\Tw۵Wg�f/%MiɩK6���9���I��ic��ت�L�vh���y���u���p@x��b I�O���)���φT~�Տ�
�\�z}�̴:�/��$��=α:67O����2���gx���Ss���1�Lt���/g���a�e�H���0��Lzc�N��dk0|�`��m0�Fw}�[ʁ�z����Եt��{R��5�g3mGL� ����ӯw���#��u�i)ƽ��^f�g�[jrT=�׵���e|gk��Y�g�h���'��{ ��$�-*I$�O�E����E�x�:�@D67��a�*���k:ۡE�=7����끤?M�X�e��"!#.P� B   � �X�1lC/Jv��n�8�Z�A�N�C��&��S��[����&��m��[�V�e�-�c�ckӥ�?�Р��F�5l�@ψR̋�fNyf�=H�"rk�z�ߟ���c� �!��
 �~Aʌ�Kc���%�����?5�0zz�Q��̓��w=��	GO�(��0<��g��2Aِ���l	�Kbƌ~�Q�	�MI�++Ak�«��B9p�;�x�;�I���{0�n���0YBj�k�}V�<����	픂�p��y$SVCE��ug�og�Fa�d����ýCk���Lw'.C����|�P}=���D�_Q����Y7����?���?�z4�!�[N�e��z&�t�������|!�jε�)�Uwtv���zI2N+�k���=����]^'������#4�����ےi�����k�w��ܪ�!�,�"��{ߨi/��EJ^6�Mv7C3 �M�C�>���`0o�F�ٱ8PO��wO�E
"����9���߬�͉1j�
Hx��2u���(��%Rj��"�X(>��"�g1�xj�9�@D%��>Lo{w����6�װ�����r߼x��;z�m��,N'J���{6H�I�!�pK|y6������Pc����'�U�o��4I����1��Ǫz���>���ZoM�ln�i��28�G�����-�Mv�����c�D|>�I=�ߤ��n�a��w[� P����WPg�ʒ۫��B��ߩ��o48�F}�M���y&B��H �!��_1�I��<��|��D:��N	}�~z9d�4���u��[#	����>%ٳj;8���]��BBe~� 