BZh91AY&SYm8�b�_�`q���#� ?���bQ���      P ��B�G�D-������JF��6�(�I��l[m�4Ѷ 2kB�����*�KMi��
1*�@,�UE5`�6��VjҋZUYe�cY���jV�-f�֖�a�Vl�!�6j�R$ՙRX�f��CDնhZ-����C<��6�m+ml�ڌU�@Y(����b��%�[fF��+fT��+L����-[5��Z٥m�bZ��m�-���-Sj�[��Y��6��D�-��8  � �G�9PږZ�:�6����AA���qI�kma�i��UJ�j�L�s��Wv�ti�p�ԶiF�iHfeeZѵ�^   9���� �.��@-����4 �k���Рq�v�$�M�c�:Р��w��wcp:�Q���p*U�V�P�v��k6Ջj��`ll"�   ����HGn�� zR��{ީ )K�f���������]2��ޞ�]�=Ǫ)JW9�*���I��С@{N��(( =릐Vƶ[)[mmiI6�
�  ����UW�x :�{�}�������� h#{g�t�({�}�ϕ�h&|���4����>�)IU��|�J��^�k�z�(
SǩGf�M���Y-�ȂQ<  g�JU		�S��� �S��
(N���
R��y����)T5y��)q���]4�w���5J�������� �Ҟ�c�BH[2i�X��W�  ^=(T�O^��mJ�8��ΔJS��{΀�wO{��W�m�4Z��� � ����.Ǧ�t�i�׮�YA;���%@��mR�-�5LM*��afUo   nVw�(�r�� �#����4P�v�Su҆����5MPi� j�s�Awjࠠ-�[�Qs�� �SU�1K[-�kٶ�E�   g^ (/�v�Gi� :�� Q��U۶p V'\�
��4C:��j�	�
 ��P[�i�����m[d��  �� �h�K4 4��� ��n �K�@k��
ݗ��.���g+�� Q:�V��E�5%X�ŭ6�1P*$�  o���5�t˗��1���-]� ]���n�������� �6�4 ��Πϑ  ��  �*R�0�0 &#M0i�S�R�U �    d ��d))*���&�4bi��F�hT�U)F       �(�	�j=D�G��ԍ4�b����M$�z�IT4ɑ����˳�<z믭�흷m[v��oӏ��rۉ��ǖ�p��r�%%a܎��:�!�C�~���|>���R�$(T�Q)W�ъE*��V>������~�������DW�T�U��i�����"�}���t�n!)V����-���F�'��t`t`z � Q4`h��!�CFM�$4d�D��CD�� x$4@ѓD4d�FM4H���$ѓF�4dс�&�4I�FN�2h��`h��F�$4@с�h�$4`h��	�D$4Hh��ѐѐ�!�	���	�!�CFCFCD�����0D��(��F�$4@Fh��!�CF���!4Hh�!�FCD&��=1h���$4d�D h�с�KFM4`x$4d�F�$с�D4A4Hh�с�I�!�Dh���F�4@ѐс�&�3$4`h���CF�4Hh�����0�M0�!��MM:$�$4`i�!�!�FCFCFC�!�CJR�$4d4`h��	�D��ѐ�	�CFCD������(��M222$���F"��&�&�MM��$��4Hh��!�!�Fta�!�C��04@�!�D��2h��04`h�ѐ�	�&�F�M$4d4d4d4I膌�04Hh�ѐѐ�!�KD�$4I4`h�h��MM0�0�������C��D&	FHh�$��HHh��ђ@ђђђHh�FI!�$I4d��2@�24`Hh���F&�$���0 p@4@��CFBCF��! h�ф��	!�&��D�4@�@ �	$ѐ$ф$ђBh��	!�	��D�&!&�HMHM �$�4d��!'FHF&� �!h�$4HрCD�&�4Bt@��HF@&		h��ђHh��ф	�	� h���CCFBFBCD$�FCD�$ h�!��ђHQ$�ѕ8�*�Y
��S�)F�$��! �$	� &�M	I4Ih�	�$HD MB Hh�	4d�4ah�FB�4a h� h�dh��!D� x h��FFM	�D82h��&��2hɢ� h�F�4I4`hɢ�4I�&�04d4`h��D&�$4@�FM=,@ѓD4`hɣ&��04d��� h�����4BhɣD��!�D��0� �4`h���@��M4Hh��!�CD������� h�h�h��!�D����a=���!�y�~�z�~up7P�K��d�SM]DfZ�tUP��dT�0-�ͳ4��^PN�^�ڻ�m���N:�֎hԶ\q�[&=ѩd6U9v ���v-�*đ�S9+a��Ү#��o���i,sˋ6���ql/�	�9W���U���{�RT"A+�5���YS���RT�fM���pX5���������i�n�lJ�V�6f]Fjޟ\�NeBq�,�5�p]˰LZ�F�\�KiL�Hi�c���CM�Ӌ[<�R��<#4=["�lhMl1F�:R��83C�N����P�F�܅�U�)f-{���N�A�+�++��E�B��FJ�ݓE��f^Vd������K�(=��mH^aX�F:d��F��0�^�N<W����@�B�س����e�ݛOhY���kn��]J�4c�.Tf[r��A�4^�.9Qm����Wv�f�e�v��%�}O���0kLf�7DȈʗ�PUq挂�%휼��2��e�q���)��*
��$�7���H$eDZ��j�9r��ݍ�����}o3-і�VhanP�e��8��ڵa�-T��t�s�{�]0�t�f~s�0ɪ�1�VlA�a;���q�)�W.�j�JV�0㊕�(�탐�3���� 	*'����N���ˆ�Ŀ6����.e���e�j2�ՖplL�t̓�m��o2�I�U��fE��w;��Q	�X ʖ9��/sA���bE�tK�$i�C�pS�q�(��[�"�$؍Z@�Ysf����������Y�K9o�XX�i?�3�j�X���bī�k.�/{ a���v ��0�f@�jw�7�5����Θ��9�3d{0��rm��X5�A`�r9��r����,�L^�
�[u&�NE�yEg�A�P��V�)e0�f�o +�NÓrJ��KG1LY�޽����l��%Ou`hF �{V�I欘]<~�E�՜Mo��{�gVkY��̬�M���љYT-�X*ૹ��bOm�S+c��C�AHh�b�'5[ޥ��p�	>���5����l^��]A���Y���D֠�,��]��L�ȍ�n�XpJR�D�=��c����l��ZӘ5�NCAэ`v��'KZ��zJ��6�3@ޔv��A�)�(�zA��u0d��v�î����jh��L����R�E��.,G.�n�3,��<��Ɍ{u��+C2�m�mI��,��h��
�8ݕ�*��j�cY�Z&�F���n�ƴY���fQl��t��JT����FK:F����{m"ڷ��Y��.^�Q�ƀe�����b/e��6�C6P�p[B������I�h��n�*�{p�0]J� �iǻRG��+qo�F�R!Y3v�7��kѺV�5`:�X��r<5�^�5�1�漹�F�N�^��0fޡC�F�r1n�Ud��rLwwGT�r��ʛ`��&n���v'u���$�shn�[~x 2l�M]]Kuhǁм�h�E�)����c@Yi;��ar*�eS�Ì�1�<�F��
���ò�����V��!NMX�NP3S�M�.�e�JJ���MW�Q�F\UhͶC�V"wktC��n'V������&�� :��R��u7a7jT�0�(�гU��+�G��]Lxڗj��.^���1{�(\�#C�Y���-�3&���M���o�J�k��%*z� r�զ�*F*�C��P�mm��Y�s`���n��Ʉ����\7p�rKf�κa�V�l�͜ZI�sif[�z#�[b��6ބ+<ra]^t�{���{c�ɤ+=87�p�A����a˻
�"�$���뙖��~F�'�a�
���˦.P�������X�������,Yc��J֎
��glyM�@0��ە���ԉV�Ǭ�z��7�s�v�8�������T��J�$�����,-����f���Q�Ng�R��ӥ�Z�6�!\��)�ՠ�o�B��4r�2H��ƣ��]���n܎���,�2��<"��*���Jm#D��k�,�:��E�k#�W!��cr�D�Ur�7W2kr� ) Rgk[Sn�Ob̀���pa�7�V^�]��Y,��p���`H(@�0X��$uf�-V�t�ۛ�jk�Bߦ�*#)��̛krj0��V�7�5$�u�Bl����e�v�U�ef���W[�Z�Z�aaP�5���"�aT��1J2�I���,��B�4�-�F��z&i�(��f���h8�<��Ӽ�`��Έ1����.��bœAmDC�i��o2�q+U����Z��_,�<�T��F���v�N��2m%��C*Pj'35,��mہ��Xι�S�[��Y�H,���3bS8l��U"��ww��A慯Y�۱��h'�q������6H����֢�Q-��<0:�Ɖ�QV#�-�L.l���%T�dWo��RQ���M�ia�P��,I��)���6��pi��W�*��m^+�(d�[�����Y�[HkP���1#B��œvl��	h=�6��r�^�N��CT\fy ���H�h02>��-�g�\���Њ* Sm�x�Br;�x2�R*�ԭ�U����:Ӊ�.-��v��[�!�&`����Cr��<��i�r�.7.�mL�r���8w5Q̣ ִnP�� ���T�^�x�0H��7��������ݗ5T�����]f��KM��q�t�v!e��Ni��5�݆ebe�sST�7-A��<��bnl` ��ݎ �ۆ��&���c�;ܪ�j �_�����T��%2�m�:�Y(⬘X�L���Y6��]L^�f]�.N���4m�_�ʘp1�l�Y	e��Sriѩ�ܴ��#���k��x,,�����K�V��~�ō�e�ȿG�ei���@�:�0)�Q�y��-��B�̽�p퇮�,��j��x�f�0��4�� "��-���<���lTsc-���qZ��0�ƅ����Y]3r���7rXf�{F���f�U�P�S%�e��H�&X��b�W�9�$R,�{�u���w$�,�˚�9���/�Bʗ
n�5a��j��H�];�a�'G0�[�4Q�0T��Zۚ� �k1���Iͻ�c����ڼgk�汫��C+�T)�2�%�,�X�U�Z�ISo���Rml;��j-�u\�6����3�mX&��
��0Uj�yc2e�u{N���Ȟ��/7h],4f����Km��˵ՙO;�W���C*���1�H�$�����P4�l]��6���n��V)	X�'�6=R��!��U0N�X�?�I��n�z~Y��>�J�&o��eGx�ql�����՛��j����1Hvx���Ʃ�m�D'�JY��*��MLkxŃ�Һ%u�򆶠9��\d*21�;Ry��,^��P�D5oj(�U�A�a�v��1� ��ɬ��Q���c�Ea�.� b�Av�����<�˫�n�7&��G���a���Ԯ�	�����չ��k�
J������0Qzk�z�RS�:Ͷ|�)��sU�YŶ'Ɔ��n]$6�¢fB�]�'ln&MF��V5����8�F��N���Ē�uh�y��[�]�w�VW�m`VN�5]]-�e�9�����7
�ӣxX��um��˫Md�֯3w�b�l�����*F6a�*�S��v�C�!����ZT��Ulx�$�u����m�ǚ�w�< ,�od5��*����{�f�`�:�-܇n.�Ų'v��(un[����m
�4I�&1[���:���q9 �ti�1;���6�Z���ۻ"�*��Ǒ�˭�X��ɺ�*�ۻ�X6�d��{�^^Jң��N�6��[Y� vj����2Uh(6{�
��ڲ�#*�w/5� ǲ����ܸ�˂I�t�"�m�6��P�QkW�5a�h2�-��rjJ�Ɛ��;PRT�ܽ�8����f�Y�D8��^Z��w�u��đ�/%��8�f�m�����3�F��fؑ�+n���8jL�CE��n��P�p*�m)�D��0�I�͸�ͯbe�(�/c�)��ڹl;mTs0A/�X���ƞ4��zUMɶf�^֑��ٺ�ݨ��Y�o}d#{2����a�`��q�xw �ͭ,]kʙ��Y�E�lՈ�Z�!5K���eR��|�b�4�ں�Ƈk�Xo���UX[��Y`��+̦%:�R�B��٦-3^�(��Z65���y�ob�=�DV
5nf����U�umc�#)�&Jٮ���aZBDUk�H t7����L�v}��%������wefr/��л�����Z��-��
(Â=ȷsu��c�S���%]
+T�U��r�dW~ku�B�B"��w~�BM�&����[-�R��Y��w�ӫkٙpk`��Rg��epMXC��ϳY$������7h.�^bܽ�
V��5ebn�7����z�CF䳌53EkJ������Ѵ�׎�+*Θ���Z�Y���}�s�k̩v�!�a5�ἄ�-�KDU�JY�D�cwH8�"R��co>j�/w-mG���ٚ��4�+pTB�ވ0[U3l�J�n��]��u��s		\�HM��K=X��\��$����纓�|GR9ySdb=�u	���ۗz������±Gw�Ja��k��H�b�:4ۛ{cw�ו(�	[0&�4�\nV%
Z��U��y�3D�u};�l�y��ߕ`w��M⻗�(��X�&�JK�)`l�ŃK[8p���7���^����x|�D�$�܅i���N�K�\ȬZ�5�Âv\D3j�d����f1ePnkB�-[i't�����#�"�T�6��5�I}ه3��Gk�y�^�:݂��A˷!�z7v�<���駨2�,o6S]b��ZOy�Q.R�.P��X5�Jn3��,��ݼ�n-�n��u)���ދ�����3N�u��:x_�����˼�iH\ƀ���܉ ]`���仲�T+f�@!H���m9������áQ�S�\+a�7oVt��vmXyF�emmcK��K	�xwsq��Z�e��՚˚7 ^e�ȍ&��DN	M��(A��-ʎAx��"xnkزH阃��0���/oH��CԱ�K���f]���!p�Јr	mMڬ{M߯n���]�u����Fv����gLT�j�%�˺��F�)�&��h���SRS��R7)�]�u�m*�"t�.���Id�=�����fMgpC�h+]6EU�!��t(U��+N�n<ܽ#���۱�K+)қ���,�(���2Ee;�qjJ��$؂���A<�1=Y׷EP�]G��0�Y�܆��Ņ+��FN�H�ʭ݈^w6Cn�g��;!���x�7��Q� �4B��*I�%���u9�����3�&�X���݌LFY�o*�,d������JCn��w�ںȦ�If^���d�ɫ8�fmM<�U���-.gO&�S�4�}T�[�{��#�-ÃcP�S��Z65�@#X�؆��(!����{�V`KQ#k�7�L�ɬ$�IPʛ�6�eڥR]�$U� Y�1�8Y �G1��;|��@�ǂ�Zv����6�i�goA�W1J�M����V�b6�mu���|���4	��i,X���:$`�g^��GPؼ�Usp��v��&4�v.�HS��Q�+t`Zd���̢�,@Ʉ�-QUL��ݰf�}u˝\G��	TMb�Y���E�5����	=y#Y�㫹a��i�r���RIv����"n̑6XB�,!ʵ2ɕx�g-`��h�`'�87p����Y�󄱢�+j�d%2̵/q�Z��d��6�R��[h�Q)�Q���ا�����yv�mj72�!L���,�+iͤnňN�l����ړ
)h�q�Ō�KȄ����s(PdᱹM�%�;��%}�E���
�a4u����ٰ��9D�r�+p�d�&������Â�t^�O5b���R�)Y��6r���	�Ml�س���9+r"�g4*w�׸�����6�Q-&��ܷ@�f��5X�6YCf�nP�:+&��`�+7mޒc�[oE���[��d�v.H6�a�� �2�)����Sr���.�I0�%"���v-��TN�w"vRٴ�m@�h;@`.�D/2U�^\�=�F�F::���'^�����:N����b��5���Y</ڬ<&K)�Kf���M��+nh��U��LtE��.�R ��9͖uTt�^̱+*^J
g�5J扖�U�� 32��e�9����G(�՜&�xpbƦ�G!�x7EZl�a-z�lm���Ɛ�jO�[�ˮ$�/����L�x�4]���Y�+]ՒV�ػ7I3�x�c�g����Jz͚���h�.��,�д�6�{Z7i��Y,&sb�Tw[D��{7��0ЄiL��I�"�f�t�;�R�,��f���ʎٌS�˅S"�9�Oj,+���W��ِd�rr#dp��&=í�;�n��u�P�.�m��/�u�7�pKI��6�a@D�^�vU���ٸ���r"Ѡ��rg5f�����5X�d߸3�U��%���1a�7e���J�*LIK�37h*x�{!�Zr�jf�q=�Z�W.:��ݗu��̒�ŢG��;�W3�{ �j�l\[�0
����l�l�"5�+���f���VlZµ���c��E�>�S2ҩ
�#Ǘ�Z��l�`�N��{~y3�ɋsC���4���J��絷%�������������o�>_?� �?��G�m�������^N�QN�uz�#���9(�Z�	p�hB�uY՝5��,Wz�v�t�q.}�4E�MLuk��w��30?�6jGhϏ���8jY+uEp�U�����6�u*f��۫����G�x#�L1&�,��Jɘ;mU�����(�AL%��0��E��B�ٛ���匝�w����z��Yi�z�Z��<�wȶ��D_qp��)�-V�NU��G�Ov<�RVW��[�y��6V��k��|�p*f��J�[�w\�8�w>gxe���v�	�"�`{�v���f<ZKW!8�1��x�CpG�Pj6�	�����$�ks��o���Q�x��I)*S��.*N\5��]��[:�e��2^���:A�T�٤�"�V0��ԇo9㳏
y����*�r�6I�L�e�H8���eo=��0�{��q��k��[��LЪ�nf�%A�G$4��HՌ�ķ��-k��v��B����;+^����$soq�Ğs�㚾5�8YVK�T���k.H°�5L9qp�G�k���ݒ�q^M����2�����v��p0I�T��kr��+O�=u�1>-
��Ӹӽ��o�-V��_eu�EUZo��!aָ�:"�����6b�R�I�3�:�&�{�XAS�V�@U�-G1bʭ}6+��\�;7eK��������k�m95�YŦV��!hb�%��]+V��x���D+�i�����(l��7GsC�]��]��.��یZhg�+]�������yR�n�>x����Zڋ���LW�4l4��6�K]�3�����gJ��Hssb4�hwdyM�;
�r��ЪM��O�ݥ�u�|7ofv
F��z���l闊�sZ�냑ɘR�L��SE�6p��V���Q�,7g9�V�5pY�DK�_��:��Cw�CX!���N���]�oD�}����'ЯQ�+�%%O1~`���f���M�6[4v��,�
{8(t�[�*uֱ�-nʌ����h#��n���;pJ��6���&���)�%/k�^%ut�z�Lg��C�mJ�p.�Wc�Z�D���ºa������w#+���jLg�#�1��٨�DQ5��a��te�{Y�3���X�3[bkε:�@��63�:;*�M��0p��Q��B�r򙙖�j�`LS(��p�m�kA�gHV�Nv�P�eCXnVs��^,I�s��ِ9��V��;�{�o��+�2�;H�p���MuB�y*c<���ykiR��:�%��:*`�G,pS6�a���FX��>��u��i f���`}�pD�U��C2�՜v�](���)G��Q�|7��r]֥����+�]���Y�Z�3�M9#IL��{�<�7ky-S+fFUF�e� �f�Ay��ۭǒ����]`F�U�Rk�S�sk/F��9���E�����9I��J
)s\"�jC�G�*�}t��)��|;,���w�[s
y����i�V"���[F #��><֒�U�pn&��IUJW���ı�x�3�K��-�n�o^V�o�`\�զHnv[$�g��M���Y-3��b�/�s6��MlZ�P�����Ykxj�Z�3,�2�zz�^BS���g���mQ��آ9c��f����..7�۾HW-��>��0[��slfU(�''fIQ���_iq�r���5V��[i=}���Ws�|F��
R�k�S���Pr��E�f�=ԙ4ʊ����(󻚦v*��{�tA�u����+���p�_���v�u���yo�{�S� ��:�wN	:�[�2��m�M�jh�=��\��m�u1В]�ɞ�b�Ooԙ�&�詭�ƞ��Z[R38���<hŘ0��%.'`ڶ]�#&�4�Vq�5����e��`�y��)�1���xܹ�5�0z��!m�t\q�F���wiZ`g��4+.�#��b��Ie�C3\�,UX�^n�{M�u�h\�P�L
���x�g�f��3���\(�Z(T�^VRt5M��)$+V�c��/b�lj*�o�̝�V���3naP�W�.2�R���tZ���+�_�c7]	(H��5Y��a'q
�VZι7U�Y�"�eAQ�B+�|�]u�vܠ�������q��+�����VC�st�<E��/t�h�!�X#��q�u���[Һ���d��	����X����cuHo��t��ML'z\<�o@��=}����X��Vܺ0ڋMfroL�x��M��;g-ӓ�;:��Gh��&��cװĵ�3�,�*�`17\o)�fn9uC՛i�A-�2��*X�PA����l��,���;L��)��i*l��3P��R��3���U��	��j�cq> �v��f��!�}��Y�o3�J�LΧ�yE��[ns�1��,>1��ɺ��Z��#f��t7�T73jQe�U^�J���m�5��r�Q<*!�-)�륢�1�Q�\#��������r�G(�>��Z�5�Ǒvr��e���Q�3���x5���r(��\�ȻXp�o���2�8�{��s�V��{1�� �k�t�JV#�[�;��Ȅj�!�r���8F.�l�7R��{�s�c�oo.Ӗs6:d9��x ��&=Mz�Y�qu�S��L.7Uș�XT��e��1`��j{�
`�P۝h�5��O.s��LF^?G�@������S�g���:��J�T���Q���5���eʝXڠ�tʇg)�Pp5�w@��j�ff[y8;�]� �2�v��V�].PΚf��ݩ��U[�(K�It �S�X�/g+��17�^��v���d���ו�J�EX�i���3o
g.a�l���g!U�2YT�޵o�P�(hW�����r���y}����脼3.��j\���A�qjD\35mq�z5d\�{
]��rд���a:�[�g;�̊�m�7`�/q�Z�mۧV7&A�3gi�uT�I�-'�r�Y�r5�BK��sN8�7#s_L<-�d0��7g�F�]�n#G4+$e��:�:�M�:����ȅ��9�U�u:Oi�v�c���"�<)#�����oV��'����]�p����J���v�"j0�$���O��ɶJ���P��5ަ��:
�9�O_tJ���di�]�{�*�zՓÇ04�ѐ��}4�[��U�2����j�mp�/+��1T�µ��M-��C�U˪��d�����B��8�2oC/yc����X�[{�b�B��l^�-#��5l��Ss�I�[8+3(��{׌�u��b3c��!�4�-fY8����a=ۖ�N�1,�t@�`�J�������K�ݟ=u�Cu���Ժ�P�+��$ۄſ[�
�r��{�����QJ�|�4F���x���C��*j�U珆A�lo�����iPK,<�w�A1�j�@�G���`�棏�u��e���᭧w��w�ҩs<��)k��g�4����s'�<���f&g��ړ�gn�b4�f�ɯg!��%K�ެj�f��6�FN'��g���[�:
˙�B�1>Z+���2l�F[���vJ�4T"��A��R:��)�4�U��M�e˫��Z�Y���ֆ��O��z��4����2ńS'd�Ç,�v�h��P�dz���w�讦^���B}�o�u�)�X�!.����m�3�L��W�^�kV4��xa�t\�r$ڽ��Ut��,�t�Ė�0cw��^�$���t��7qVْ������4��y��yG7��Pwg�y��Y|�W�u���e5gg9�4��qK}Իesp�5+OF�&P����J� �5۷(�\���A�Ѳ�9F�gN�ʧu5E)�/V^2H���3*���W�j<��p��g$YE؛Qu�Ә32��n��x�Vʹ{s $�6\��q�+n��ɝ}�,�ųt6�i]�<s#���
nj�k��J���������qX$���$N/��7V�KF�9s-�wr��܅ͮ����r��Rr��[�.\q�{�.��B�wmY��i�y*̲�4ouY2"c� ������RnT��F!�#UN^�c��̩s��{�s�j��'r�3K/n^c3*Ts�4��z5\��Ж�b��)+�Y���]1�\"���LB�
���ۏ�J�Dͻ�o��]��1��̧�<J�7��FaE�b�{	���6]ғ+i�<�� ލ+��;�.��J�-�5NW\�sP������k/!v��7�8�gWd8E�����.������a�.rY���%�:�*(�L�3�m�5�q_]�dllm	R
͕���x�wjmK\����WXf�讠9)µ�!84�zNfI�����R�@�H�J09����H=�'m��2m��n��V
�����u��.���c�d��
�a6�G����7*�L�P�2
�ќ�y&#U��I��i
F��r<#D�}p�����+�.s�I��l������6F!�8��&4�=�����\�Y�ԺZgL�v2:Q傺ܾ2--�c/�+g���Z�.}�:�-��=
D�s��A�b�=���&3�u1�s4P�I}����K��B��OeY�Ι�X(�	}j�N��e�2����
r��ɸ�ۑܾP�4�ɦ�-W�i�$eiڎ�]��#/���n��X��!ӏo���+~�{���Z6�:����N�l<X��t�^�n��rn�5�ś�7z(��g�vy�����6!�Z�!AVdBL���3�B�g��o"��wi.{�OG�gQ<ۦ��E�om�����Ƕ|V(���VU)�k	��eFɌǣU�(�m��CJeod�B���]8�H�O4{��v�r�ES7D�$ \�]w�5��t�>��u�mG'Xe5��#.K�݌a�����}c`��mn�cg=�)�qۑZ�y󗶵=n.���H�M��[%.Uɻ�]}V�L1�Q4s���Vb|�ӭ&gP�	sh����L��i����^�����4��d[,E�������t�J931@�B�cbuY���"u�rմ�X�T-��-�k�Cz.W�RŅ��#C+W�(,�uu��]O�"q@����8��k+��e(v��;�7Ӯ~=�J÷��7Nww�Z$ݛt͉�V�B똈��3n��cl�γW�d8
�e)}
��N"��{�I��D5�mKU�ba��]�mMy�%b�����MӺP�K�lf�g]\��W�r�\�U�m�I�I,f����,�|�[����އ}b��\&g0���x8�N�Ų7�M�x^�mS<4J�c��L�ݶM��/s�N��dh�yS9e��/9px�cRި�DvWcy�Dkr`�Z�,�g�`t�V�*�H�Y;�-�q81F2��(,t��eނw79�R�����׵G>-dB]*s���ޖ�|.����lt
��6�QL���*m�Cr1)
�q��K�p�q(N>�V�N!�`������zv�h��)����ț���h�ʹ����UϔwyeYnon�CڥM�rɥ�p1��pC�\�G�VYp#V��{�bt�G���ٚ~�/^Jyb:USNv`�N���ً������x]�ݜQf��*n_)F�l�.�`��I`�7��F�k�ʫY���sʳ����u�X-��N�p��7�V����,R���p�JY �<ue�Z�.;ӣ��۱v��s��{��k�/%8.,��89�� V��k O� ){��*���B�Bq{r�%�8�]�ɽ��֊R.�v���$��d�Qw-�;"���{ͭ/7�h�G+��u6-�֩�+|��`�uk8��7tdBLe3P��RJ-���,�ٛ9�~�R��MIY���v�T����W�^Kϛ�$��6|il�m_���Cg3����A����֧�x�v���yW'*�a^� n2�����;2�e��˘�5fv`1V�pt��\6��s,R;���̪��96�7r%*Pm��F�����OD뭸x�� �
��In���]��oT��[	rh�}OE��V�*�b���]H2�����+�a�dA0p�[D�ܥn|��Π�^��Ʌ��m�_a���Rv)�e�:3��}�m����Ή˂Ų�}��9�;:Y��%
p�R��VޙNG�9q�t�ݼ�Y�;oFB�[���v�����G�S�$=�u�t��m��YД�vq�T�׸j��'�@V[���K�b���Ql���-!#Yt2k�Z�F�̫5��G���fBfG����0��k(w�nJ0uC7g)p]��U<��i�;b��o���蛸�n�9��)��G������}��)L�׹��h5�.f>J`x���x�g9G�t�A���7;2�(u��\���;_F$���̙�Ū�56�WL��������+fe�;,�3��Ƕ�
�����w�Q��gp���1M�ˀ	@�ƇPC�����g��C���>!�'����rf҉5Ϙf�Y��������'ϗFyl�����'sۍ�Xw�S�V6��p<��9��yùG��l"��3Vٚ�&��qޚﻈ�C�^#�g�to����z.�����p始:H!�
7�i�@!�ێ�1x`��,����֠=�Ǐ���{�����|�
��d�i��<�d;�Lz+�U����ݽ�Ve���5�
B`�$j���4	4P�$�q8��d=��SB@�I/ElquW$��D�����͛'$:�f��I�g���,�5��P��q�n۷v���^l��!X#�z����������Q�ں��� M�Uo,<z��e����/�������jk;�'��'M�����<�#o�pp�<�nͷ�i�B�+���֐�7�|9��_/'��^���?�������V��ѿ�[ޤ�wx6r+��o8j[`T���EpN��v'�Ч���Ι�Kv��%H��'2��p14�����r,��rr*�鷵�S��=�4%r֝Ս���޹f1�;/�37Me�����ܣ�/���j�4��3�����y���)@~Q����7���JGU%�̷R��ݔd�-n��eP7�xW���^b�L�sv0B}�S������ك/��J�-h*�W9S�}M��v1B��3���U��;c$q���-q[h�?f�B�cn�k*Ȼr��`��HÖ�&�XPՐP�H��POE�\�lw#Ej���TE��-K;Gl6���Ճ�m�=G_Wki��D����kU�)_muu�k֣���FL��rAU���8�Gn2�P,K��1L��G�����+N�`��.�I֞��]TC;aZ���wQλΩ&�huz&4Q[=�:q��T���T��|�p�m��Y����t�_u4r���s�GF���F&j�t�e��a�{��c��/�{��7ld�%	�CR=���r�oT��fC�U�E�{��g�p�ߎ��s��ǗsvsE8�t��5`�鬃��g.<��@�fk�����u��:�U��V��mu�������\�67qgK��ef�$�(���<���K�J��o�p�[�%ת��-�\�k�}�ћyP���I�5ޭ� ��b �A@� � � "  � �AA� � � �w�'|3��sM%p��Km�B[ѣwlǱ>�v3I��8��5�ע#�2Έ��v1��N�v�J�_d2�U�����w\��)aor��>�8����V�lķIJEF���癝ЭE�ܨLf��gp��R�9r������&����a��:���N��9g,�s�s�v�eCD��ܭ۽���e'N�|�b�`:�6����	����7ۮ��ukL\���i��Qg�UXC�]u��ڡa��v����'ax�I]N��2��m���qwvv��<�J	�K�V��<��.��f��&ܼ1��W��;iύu��15&���|��6o˖�ǎQO�Z�M����uh�ՙy�rӇmE]5��V�G��w���l� �����
J(z�U��`�1�$>7I�[���y��^�����;6^�%���>�����^#�k�si¥t�®���[��X��7x_	v�)�[]m�����]WCHv��s�GL�҈i��/5챱���&�-WOSf�n�nnd���n�yq�t{s��ۏ+lrԲeh�,�A�ӆ�ZF~ѡc�Z�9u�W\�AH��j��4�b��*!)�K��������/'5.su�Ju'Uܚs~uQ���VUKI𺏲S�K+��B��B�{394�z**·�hp�����Ax1A! � � ��@AA � ��
AA ���m�mJNnH�-�z���s�W,5�-�����K���S�ˎ0��y�����Z8o\������#X\ݚ�
'�����c�tu�TS��Ɩ[��}��ePM��Vr��Q�B�N}�CTf�|�R�15�����&��*?h�VonͥPL�v-	y�$�L�D�_j�(m�#��i]u35F6w��Sf_(����WTє�����Kf��<��8Uh�dQT|O0apZr^��Y����աA^k7M�8ol1-�Rc�����n|_%XR�v�Yt4Z�:{�NZ�HGJ5���:��Ba۾��n'�S�,d�n=���N��fzd�5��i�0e�̼gr��=�8��p|�fcqX���"�&�ouo,Mҭ�e��8����ұ���(���J�S�+{��-hÊ���!>�1�m��
�	\ň捗uu/� �A�����,�ZF�8L�QI��_%�`��^J1"�L�uSje�f���Cr�n��2�g$`�n�O  �}��G� �{�R�Y�������n`4�}���Y|�Ϻ�,�_:ī��7�D��C��z0���}ֲ<If�X]yo4��I�6á�))�Q�s��w��ɾ6�;J�U��x�`go,-��"�n�rx�hr�G�ɀ��̈́��A��.���m���D8Xѣ�@� �A� �A! � � � � � � � � YˮѪ�C|,;�:G9Svx<�⥑[g���&֒���J�-b\�#{.`C�%j�5��\��9���q��}H�"�����K�E��y�ܽ�H�D��c�҅،uT�,4{^�J�H
k
;ҹY�b��m�����of�J��0�3�RuS�4�i��_#34�Ж��bb8��]l[�y@ui������DMy�;��z�gEvR4%�j>+72�ۙ~�sqG���tI�$2���.t�����r�b�l�mYc6�U�a��#z�.�^h�V�dT�����s$��CI��H��藀�2�J�Cnf#r��{�&���|�u+�x���H�d]���Q ���x,�!�V���ɳ��č�
�e�?Q:�0���/;��&��{ZԪ^�O�6A�k�,Y83Jf����]X�1pR�.�ҞD�'�WՑ*�L�%T���N�wE����$s���7��
-$L$�����>����c��q��ۻ�nbh-x�Ҧ�D9ҕ�$;H(
��5�%>(6����K�5���`'v-ipR���>U.�� ,�=��_t�vO
Ùmb��̣u�@����5b�u8���c1uLZ&��@(�Ѻ��AVl)Mˢ̮�M��Rl�gz�uv���!��)"a�J���s��˗�у;�=�#t��[����mc,X���A� �0AA� BX� � � � �,AA �AA�`N+�fSz�,���Wf�2�dŜ#���L�� Ρ�ͅ|�^-��!��/SѦ��a�k�`�l16V��U��A��m�b:hM�������
��uy��UA0�a���
��X�핌Js�����[<z�d9�MŢ�W������,l�Kr�n�ifg�V�!�\�Q�J�?Z�k'�$�W�kT/r��=�S�5���!D�<�UN�-�T��x�a��LI��2;x��OO3�f+,l��	J2�m�C}CM\��!m��o47HWlӸp�J���Y�X9ͼ�ܣ1Y'��fj�n��We�Oa��<H1cv��l�	neV��QdLq'Zmh�U�m&�����tֶ�!����z7gr����e�< Kc��sJ�ܚ����.����S/-���-G`�;'S���s�í�����%�����Yg6FJ���w0��Y�4�I�r�z_Iå�F��8�o��U��m��
P���xpa���һCF3.�>w	ZK��2�'������`���\���OJ��s6�n��
ds�U��.`�!wuv�쒻�J-Y�n�h�Xz�%��J�j��P&��P�q���w�v�!���qEwZy)��>7�ݵ�j�����"L�ܑX�]j)�V��b��w`�(���!;06$��V��4�ƺ���O�׏5�{Y���JÁ Ɔ�AA� �A � � b�A �4AA� �B�/a��Ve<�w�ntʲΗ�sZ�5|�|[J��MLZ���6�#�K�/X-��,1����v�fD�;��F0v���a�Ռ�WSUU�͎�0�va�m_1�nI"�����M���4h{�^��C�\����$7�ӗ�@Q�`e}�u��7-�uvT��+�+kWv-��F*VA��)���IJ`TEZH�<)��_n�3X�Y���ُ�K7����گ������T�(`�|�Ձ�eU���V=����ʔc�n�r�a\ԖT�-����es=�`�LuΨ����v�&��˗���N�jg�<H�4*[�2��)=�iִ��FlOpod[� ��ח�+��aY��di�t�tt��p�����ۦ����)ۉbٚȢ2'/�����Ὢ�b�{��t�ᬪɂio}���	fĲK�u�����{V\�y^��9sGNQG�u����7����z5��cT����[�ps��Z ����Y۴�T��(�̊F��r w�P�{.Й����)�f_�()9n8a�?q{r�(c��[�1�j�����i���Y�L9��V]��8&+�iq�jUrA(�����S���7dou���uشM%�c�=2����qڵ;kr�]�y���:�[�eX[S�Q��:g�X��,�(!0� ��AA� �A �0AAb� �8A � �A����9��B��3b}V9\��S�HeR�T޸�L����sO�q�nt�3@�EǠ���Eژ�sZ�rH�Y��Y��`Md�4l�#�WgY.)��,e$�X�����5�'4�ɣʻms�u�V�t�����QuDu��T&|膻���-�Y����b���z)-D�j�U��BL=����ąk1ӎmN*�t��\�vkeure����]� Yl�y�h��t�j��/���A��]&h����K-@��n�R�7�-:Wk�u�턡�8ѕ���Y6��SEUO��Q�L�Sc�2.��L���Ce��n8�h��x��6��<��-���r����.���b1m�!ID]+�fh$Cw�vVIsp�M��@��uۓ�@ʴ�5
]��a�������D����QKc�Gdw)��}Χ4J�ٔ{���:b��l�H�;3,7�7`�+���qt��5;5>�hpl�rݠ�m�m�gQճ��>�B��ej[�rBiA�/���u�!��c䆼\��SA���VͬCI�4ɢf�����i*�!�P=�4�ɒ�+K�[��0��#���mu쨮��*�0���k����&x�����Gmqx/I���& o^k�
А��I�Խ�x�+�>:[M�ea͚sJE�j��b�6�`��dA�u��xg�E�к��8@�AB � � �A �0AX�b � �� � ��+.���ż��N��NRd��+�֚;�r8��Z��G8���=�@o4)���t��V�Q0�u���M]s����\140a}rM�Ur�Q<���mM���CSi��?7 ̣y���=��]�����s5�κ7�)e�n� ��Vh��LR�障�d�%�Li�����ͻ��I ����±).�C.�N���g���/��D�º)�Kq_JQ6f�z\a��}���^����^�ۓB�;y�2���A�t��f�6�X�Eu���~ySes(.l�BzMeS�о�c/�mαX����tnX�0�B�8�`��k��,Ywӽa��zu��QT���I�]f��͈�O-�I+�<��Ɋ���<Z����Y�`�Dڇ��� �q�![/ol���c�C��o��
?y�yNwH���w��ؘˈ�C�aɚ<�3*`��{�Y��IpW]{�܆>Â��MWZ�^��M�R�*-w0��փ\�z�kQr�2Mٸ,[OBK�]���G����Q*B,�d��E�MN����:�w���{��-b���3�U���q���+"����{Iƚ���%}�5��J��ni,�c:�ت8t9���eL�s��df�D|eY5�����R��V�
uqe�p�9����ߩ�\��%)�l2�o�E����C΋A�WG��,(O:(�'MM�7���#':�S���MJ��B�h�(Vmv#P���+�i�*�롷E��!b! � � �AA �A,X� � � ��(AA@�7>���u�N��E�B١�X���oS�a�X8�TX��部޿̴�^���\��ۤ�/�A��䄂�@��mn�Գ�/�Vmgb�H�!+�yt���D�Q	G�^}�r\.�1O�$����':*6ߗL������V��/�dh�d���ÜZ𕘳U
[[1b/.mb��E�!��ȵf'ǰ��Dw��P[��
�@��Q��-����S�B&��i���	K"֞�++��惤Su�p�o�vϒ��oC=m��gZ���kw
���i�FJ@��y}����i�]��Y�e:�Y��J��͝�Z��m���]�|�n5UC@@w:�^l��.}|��e�!lR��W۫��Nj�5�l�Ժս�(�ޗ�>�=c�lff}��c�X��5���r��]�d�^ݪ�ij���[å0�J���I�bV�2�y`E�wp5����st22?�"#s���a��0Sl�Uv0�lӺO���W,���>��8���d{��-�M֩ ��p,�wn���t��n�6:�j���o1ω��쫌�G-���"f�w�
��9
�L�����{Z��8.���h��v7k�}x�N�z�Q�<|�\[�]f���8�k�¥�F�%v�#똬gv��f����n&aݘqn��3�M���n�؝\:��`W3���L&$�ف>Z+]\�wR�	]��Uغ%G�BE�ј�Y6*��l�hVv��1SH�~ET��&nh-A�b��dX�r�����x�b�D�x�ukz�쩵o*+�2t�0V�f���u��.��n�ٌ\v����A�1U;Wß+�enݫfWT�gRq6}	 �I��p�.ٝ5����Td|�TZ��-ZMC㯯ĹT^v��U6�bpJ�ѯ���^�0P�ņ���ʆn�*LZso�q��eE����U�:�Y��Em����:�(�vby�L�4h�8^�zA������9����"���uYMc=��)̪9�U�^%�M٢�m$J�Z��b�˴��Ka��hm������s,Ṃ�=��Y�v	B�@�(�f�Y3�D_�Я�NT�m�=a,�rD)v�ӏ�tjY
V�l�o&5�}�[�*�tK�)h��QĖFi^���5�A0`1k�P�|G �~&G���an��Y�f�;����3r��fk)��>����y��	uV���.J$�S^���anm�4�w٘�v���R^d�p����:|9P�'fr�x��e�Q�*�D(bƯk]hV�f�r��I<���+6=�����ƶ�䶸7����0Kآv�]�챏��0LJ�����X�ώ:D^Ki2Ȓ
�[k,f7Z�2�-� ����r$�6E+Q[�Ҷ�L@��k�ܞzS|�}�g0����G����^����g��|~����8u�����n�^�g����c�;};��(Ѓm�y��vY�'����D;&䤪N2�24������z��W�#�5oG	}}5r�d��I2��歶�:N� ��kr�1��d�K�������cl�0��o�L��2�V^"��OO�8P�����:����b�M �1;��oE��(tu��:iQF��<�M�*<��1�֣ھ�I��++:l�n���B��O)frν��T6v�y�A��W��:���]{{.�r�l��vC\Uc�s������Z}���n*��S��UE�����F�h���Z�w\�K����\T���b��M�M�M�W��OMXN�u!��TW֭�o(`ެ�/*�e'z6F����d�[t `�g�+��Q3�V4KhP-D�W+J��F�;hA"N�y��]	��������wD�A��m*�lV�5w9�eL����Ll��Y�]oQ�ǝ�l�I��"�kVZI#ݘjŚm#�뀧m;�y��]��&�Įϴ��7���a]�L��������iX�Ӱ�B�lչ�sۧ��>����!��\5�v�p������sf\�䙵3��r��G71p۹��Yf�۪��E��Iv��N fY9�VgU�4t�n;�7X��5@��eΩ�vj��^*-+x�e�×�+Ĺ�ǘ7��s+x�j�9�y0�g-ż�j)H�(��;*�����KiZ�*��#q�#{��8�Q��G�-��B4��*:~����;I�)6J���DԊ$�)
I�4����2�)�??Ĳ6,�!�I��DY<hM"���[@��h0��&�R$��܈2 e��A�5��ʐ/��JE��8.HbiJ^f�c�L91ƹʪ��.9�����̮as���	�����/2�L�2(��Qc�jU��+9��Q����F"քQV��N|:t�1;R����B�{�([QDr��0b�[�aS1�-X�33���æ��:�F2�+j`J�x�ۈcQ�Q�Pg�ab6�DPQC��*z���4ӧF�Qxw���1��m��J3ĬzY�1�)�b*"�
J*��Vұb�S�ONΨ�*�j��Uz8��s�Y�,Q�r�Q�\�b�ѩK}o����+�"a�����^!�~y�1h��h��}�Q^���~���-[h�b�j*"ᝍ�Y"�P�������8\�^a�f5��Nc�PTn8�4�Dm(�r���9��3[F�%S����p��k�'�s���qL���çO��ӳ�}ʘZ�[��b��f-�嫈�NfY�~�q<�r��2�eA�V�җ���TZ��\�-���fPę���F����Zt���zt���AADR�[1� �T�D�P*5�� ��R/��Um-�B���9q2�W32��
R�^�\[F ��a�+m[ciPm�QE
�K
"���\<r9����TZxն�ڱR�#�S�F�[DPZ!Kj�{�
س���)��r�R�_UQ�n�
��p�x�9�õԝ:Cwd�f���w>�vv��(�a����z���rԝ�!�R`�w�`�n�z���Or�.�IV��
/�N��]�e<��ޝ��F�ئQ�\�X�}��?+��A�.��k��t ��6H�:�g`��1eM��.1{���az�~���c]�-���9�`���}��ׅz¥��@�v��庞�80�p�G��_�}o�����C7K31�'6^ݳ�Gl��f��^3�=~��oQ6O�dA���g��~���J�S�a��g)��3d��s�>��n��b����D��+x�k �^�U�������n7�;M��7�������� �8d��zG��D��������7 �a<�<�<'x�w��پ)�y� �ו-���%;��5����<����z/'�M��9�n^���w��>�a�E���#�f爋�8D����nO�E���4jNq{��I��g�����Z�Q=[�w��ғ���{�%7�B���������$�2��Kޠtmm�-+]9=JM;�����xE���g��֍��$6��^j���!��V��t�D�_Z�K��V���+x�ƭ�s]9oL�W��R��;t�A����^eq����I����Dv�³�-j��D5���Ŕ��f��Wr�ɉ9�y�� ���=��Ģ���k��c���^�G~�6_�^9��;��,�;��W�>����L�i��!�o�7�{���}b_{��H�/�K~�k��p��z	|�D6�8^u���]��}��w�#����Ž���g�(���;����H~�Uz����W��j_����-����hl���� {�4"`�W�ݤ�m�F���I�'S	��������K��Ox�޽�l��y����l��k& �+I�7�=f>�O	>5׳�O@�
���K敛�ǻx^ِ/(_�|χ��h��W5��E�!�:�����������n~����l�����]e`��t�����#��]{�s�4خ�M�olW�؋�^�N&�¾��I�;�	y����ӄ��y�öI7�'��o�n��
kƢ����0ks�]}����0������FM���l�85�|IL\�EGڦ�:5T��.�Ua�[�X�]$�27^��q�����Bg��Cf��חr�ۛ��WL�����l�w�i����<����f��m�=�7����{��vfL�r�f3�W��p!���z��kdG�=�Mx��c�H�>�{c�}���p�C�)ös1�U]L�z4W�<:S��%fg���ǿs���:z�|��<��Koo�0����Lx����t7�R�?���2�z�/�{���"�E����W��'��j��~�ߖ�K���@�r�!z`����]�UK���why��K��[�;���x�凑�v)���G�=,m�ˈ�C�gh��3K<���_��x�1�=R[�01�hB�H����=�M_���Ut���y�~3|���s����zܸ�\��!��T\�
�\�'N���6��@�z����*z4f�	�"Os��5b�8� gH5����9���9,���.������Y���y��goc�L���|5�c����l�Z���wV=���u ����[������r�tR�b�W�Z�7��Q�j���z������4�v
ϟ���w���E=��@���%�WN�+F�`3m��%�|������뵻S9.���у("e��Z�i�ǵ�)�PAok�V�&�,�y��F>�\����ven�z����Um���N�B~�_�����"�0��>���{�dPP��*���}������?��OY2\��ѳNh�W�<-�x�|�z�+:[Oۧ��A��2�A�i����ĝ�<f��Ƕ��2UJ����Ƕ�Ӽ}��0z���f�n�'��#^L����Bq����n������G�8����4m�ì�y������(k��ݓ�=y(���%����2�����_)*��W�����`o>~y�y2h��,gv_r��:�}-#�>�z�zL~U~5��}Wb�}�1�~�Dm13m�O'&ˍ�<	�-O���yn���o�73�y�]����T��q�ٻ�U�Ի�-��K��D�����K�E������.};���,>�z�ϼ����=��6�~��z��r݈�k=A]W�c��n���בּMąѹ5Uc
�P����O�q�RW���ޟ��(�B�'��הe�Α�%*�#,��F��y'+�p��S�/N��}�B0vb���\�Y�c}��s�rO��#�8�V`�6����s�P�Ig�J�6�lE�&u���J�E�[�lptX�Q+]؞�A.}0jh��H7��P��~����q��c�_my�(xsx/�~��{���ֱP_�
R�k��-�=����=��.Fg�;��4@X��x_�a]����Y�|8��B�3��=�D���shz�	�{��H/Vy�>7��ޭ��
�t����s���u֌�"�g�^{7@F���A�7&�OcH�����K�b(�4�j7��;�:h8x��ͤ�&����k��V�������ߣK�yѼ��F��ޞ���ڀ6��H��´�k�z�<�I=�E�dSh��y=æ���˹̷���u��[�p�GLwNn��k4���ƗM}�r?w��m;��*h�l��t9��6{2yWTG��uj��|=�|\=4��O��]ҽ����&z{�90yB�M��^֏o�.4k����<��*���q�u��wA)��MC�rK� �u��}u��V\���������꼰���T���v��!�Gt|Yon��win�bGKK������`��������	F�Go�Q��90�M���3�����lvf�Sy�.�Ά-ˎDVS���CS����f�螓�/��/�#��=��ѕ=Q�<pye��~���:C�_-<7���]�]�}Tq��p$E+�{��p���7�ɹӧ(��;�O��k1��9�����B]���-�g%?z	�Fg/uW��<rY��/���Zm�
�����**�bRzqƴw`�X����wo���^��d��	L���~��%��#c�b������dvu�؜s�/tn�?���+>��\����tClp���K�T�����ٲ������4o7�����p���w'�l�<͞�� lS̛��40�<�iu=}�,����'`��l�WX�����O������ן)m�Z�%yu��^>2G{�f�f��?p����3dײb�����rf��q��/�[����Y�˙��O:`�l�;�^�K]��m'F�Ķ�c��2�u)�����S����lE�^p�m���3��M��s^s3��G�V)DfX�s�4�.ms��u���TF�nE��oyCh���λ�/�[�΁.���9��v���Y��mm�ʏ��/o��^P@��@�Ŵ�y�p��U��sL���by��n%��>����g�޸1��0<{s�H}m�t�8���7��#�8��<�ǫ�Oߋ��P��d(M�����-�7|ڲ	�l�1��
��+KF��7�'��_�~�}2��\`��[���������+�5d{/����;�t�/�`�ߨ>�]Y��Y*���ޕ�����o��C��d�+d[_s�oOC���g,�ӷ�r\�����1���x'tC�\˵�ȷ��Y�Ƿ����V�^9�U>�No/��a��ma}��y�au��*���W�n�y������&
�ݢG�-��Ƽ���"�A�z�7������ ���,�޶V~�����@�$��M~f��p�G��"C�{"j�dki<}ϕ�n��@r�������3آ2�w����+�ȹ�2�2nj����yl(�1"y�)^ɶr��uT�E�(c��w@�k{�\/�i��S�������'�ˣz���ِ�� ����.ջx�(���nJ�[N͕��b��k���=������9�`�K�����{�P׍W5�έ�c/î���g�o���혬/��޹��9uȊ���3%�W��u�;������xK��k�nT��y�{=�޴��"�ߘ�m�]}�D��#���I��{[>Lvhu����a9�H)�:�7�N���RA�K'������������۾2��h0�G����d���mp�{�����X����ū��V��G9��=]��9�U��
B�|켞��k|,W��s����ts�48�.`q�1�[���sTʡ�=��m���~~~b�0=84Ef�n�'��Ǝ��y�r*Z{���"���a���x� ���y�|}ϡ�sֽ2��ܔ��_������D�������P�c�t�P�c,>p7�gN|�f7~�+k��~��	���lm��B���D{iڙ�n��9A�|F��)佼P)|׼3Փ�c����i�X	�fԲ��tO)L;	����7q�[9D��ТN�y��f�ֵ����Z��3OuZ���Z�\�yX���[;_���H��L���� �Q!{��x�z�T���/6VO�3m�WQ1\{�iƏ���k����~���W|�^�Y��_��[4랞�Gw��'����Wk5��n�7��H^����a��(	�N������ڏˇ�!7�_���0Ps���[2��Y�'I����걻d$��p�>Y�ޚ<^v�=��1�Ի��Z�a�]�׶��G7�z�WDxz�C�Q[���{�0c��(oN&:l��������îȉ\1y�y�m�a�=�ZwS�*�6� -(� �r�M���s�ă��ðY�tS���]vO_��\'�ɏ��Wy<V9?}���k�8:)�CU��l�c�ζ���9�L���QDLܚ���&���h�=�>O�o̓�/ª�{���z���!����f͓�������M�������^[���q������Utf �փq�������jQ�F.�~����:��ĥ7�����N^�ּ�G�6W��Uw��۲�L!�3�;��Y�^�E*�>F>�OQ�2���v7��K�&�-8��f�f��̾�t�$B�'*�$�����o6�A��c�����X��=��ת��ӻ�>��M���7tܖ���cO���s�0k�ݷ�֎Ù�ٝ�)��/
����x���
z���$E�;���w�b=��o�	i�Ul�J��/��p�̞ߟ��ή?��x%��|���>���%s�k�^�~����uؤz���/cb��f����p�����Rh�0�ES�x���o�����}�.x��U���4wht���;I/��:{c�*�ؽ���WAp�h�d{�f�E��������NW��y9ϑ"��a&�/,�H3���5�ާc�-ѝϽ]�tr�%x�+����}t�t��_`��v'M,0īC��+� ���ȁҳ���9f�4�:G���	/������}h�t�� }��fX�\!���R�[��l;�^�e���Y����_k9i쾐�7CF�Y����\���� �9F�J�y9�g�e�r�dͼnm�srC��S�,��}��hƞҡ� �vз��W5�
dC)�*��wI`�Z$\woI���cKB�O�h�g=�*,�/�`�N�8u�>�G�]  K��m��I>&S{MZK`���K������zmCm��/��5'Jܘ�)���٬�-�n
r���<EjK�{��FEw$���^֬X���s:Dy�Vvܫ�@��1�57/
Tg_DN���`a4�S]�&0��M��8��Pʶ

�\���`y�3v�F�Tw�
a�iYk;t.s�}�ݜʲ0oS��I<�-sÝ�/RB$-C��%j
��
�%��3��/)#\V����Q�\D�v���Z�nE�2�賎�@q���4�&��:�oD.�Cf���ûG���뭐+�uw�n��]c^-f�����6.wU�*�خL*�J|�����qbӬ�x+rPKn��F��JMT�n��<tJ���Ewnkv�c�q(�B�1��]s��e�6��)ng���ӭE�)�c�Ko����)�Ӳ���Ԡ�G�K8�DHG��	a��>#~w�O4AU�t9qzz�1)�>Օ�궉��J�9p9y�Lա�l�/�VC���Vwz+���|�'�>�O���7�dh܇9�����˼60L5��m 5��]�!5��w
�B'QFٱ�&��db�لD�����:ޔ�����[��ׄ|�tӿ-pM�4Xu���o3�ge���<#��n��}&>�u��.�Z�5�{��Wg'��4��y)%y'��b������>E��\p�2�B��y�}�{�FJ=~�^6�i�)�K0Z�Y1�[�p��DGK�gMrbx�7aw��z�繓f^�� �ܾA̽c�`F�;1�����nrj�ev��|���s{M+D]ͪ�ù,A��8ℳ#A�F7��t:�Y��%]���r��7�[�}n+4:�&n�N�ԫ�T�DnL6�d&��ꎅvh��0e3%@�I�P�eu���Y��Z�*k��nڝ�ش��&"�Y-a(�u�N���"r���l3e�ܬ�C�V0b�W8c\z�kM�.����̷bC	̒�ʗ啎�d̓�Q٨!d�̝@�y.V�kN�&-�c�N�ٵ�!P-i�S��U������<èa��Mr�������LƟ^�3j_n� ���fr�[��R�	�6_.C$�`�{�em�\��u��N��h�c�:��]�ɲ�`��G�kt�j<��&�h/��:��߉�xKfv�lZ3��%�y
���[CT�uN(5�����h�	\��3q������E⡆�3C�fOY���2n)R@�³!�"��-�p�\�Y���NO9/{'5<3K[��Ռ�޷���y�e���[���,��\+�m�˙��(�q�
��cL>�1�-�5Em�m�&<:t�9�Ǯ&%���G1ÙCA9J`���Ԭc�,�����8��{�g�f1j{Nӧ�D:1QJ�U=���NR�����fX�U2��f	�.9B�a0AѪ��V
!N4���}=���X�ڱyi��µ-h�0Q6��DExYQJ�0�E�gs�"0E8t�ON��+@D`*U}@�* �*#֢�R�r�����(�S�8zt����Q\j�D�Qz�k*�hW�����KYER�`#�e�em�\R�t����֠*��b���*�|�r�������PT\�VZQ;IVa�����;km�Z8��TEg��Y�
5�H�U�����K*1S���:�'��Q�Q-�q�
���V

�j�deeU�T�Ub�����Lh��"���A^R�#���U���*
/�xC�2�}+�T����"�����ǩ
lZ��l�r��vn��øf���*���y1�W�TԪ]v�7*� ��&xAހ�d�ٸ��:����k!/^�C׉�=^v�8�_�stרk�,K�_�t<�OUP;KQx���ž#a4��|��o��7hkNnu3���%�?d��R��y�t޾Kyc�8�z?q �^߯w�������)S=��hj �i�;o6&��y�^�rR͋��ƅ�� �_3v�?������%�W��{:l�c�h] K���p9/"0X��U\�V�ϰ��a��u4��M�f�&�{������M}�:���:a�V�7���U�I�>c'�s�@�հW�$.6�o��Tg6�7Ȳ�a\bYID�>�i7��;�0ݩ�'��y��(���U���,�/�m����!e�@"�=����;�fS�c�
b������j��z�Ԏ�d��_^!���`g��;P��P�,b�E�6D!�zzY��}%�H��6�[g�E'+=�"�-�a�^=_ۻ�q�ֹ�.Wn����W��B�G�:m�1��F��S��uL5�M��8�O	4��X�sѝwM��V���@��(��!��VG�|��kÐ���Umt�u�g*���E��n�3�Z�^��S�q
Μ9Ҝ�ڱ�˂��nN��-�5nY��G���\���<#�UP٬b�L��oJVdz�̗�nǹ����'���h��2w3w�͚�/vc�f˾qީ�����돁oX�\Wd���pxf�	��(g]���w�� Z��s��N��t;a0M^��q��"�D�����*��@$|�y�&���Kw��܋W��Xך�b�nc����r�W���R�Dx�pP�8-����JhVD7��nw?�V`��*��n�ù�k,rz<';�k�]X�\���Nd�iDgۥ��5�V,m�52�ܞ�>v`['׽B6���Q��QÒ��RQ\�~,����q���scȝ��8f"/�-9o;,�"`㫘-�����Bhq�.�	�o�Lt8mGs����S�-�N��}O���ClP>!�4nG3æ	�u�P�Nldha�����s��0�$�]�nu*�eL<V�p�E�heMa��� ��>L_�bu[$��`I�xi�����>��x��{\���k�*����Km������9�T��(�3�f�P��t��N�,��|���a�#�����۵L�j9#:���j�!>�����{DH�W+������eEÚ�X�|���N��}�2�<�}�:B�qP�J���Z��0�?B���B�B��^,-�\[Ot\:�r���[��V]�q���,����+�M~�<z���&�ϣ�<��ۆ��í�EG�nK[/���Ǧ�
��[y�TmM�>����6��vD�v�5zN,:�uI��s��׊c�Y���uŭX�+f�%��|�xc'n�f��×��y��R�n�4A%6� �ՙ+z�6�zǨ�`�k����3r#�������	�{1���J�5��E8��[�Ķ�x�Z2��&zu�2ޚ1���7�A�{��`�_U�'��?^�F�J�-�	�J$g�c�a��
z���Q�OZ�i]@�t�z�-�'���#���Agk�&`���c}���C6�d4".� �.��ڄu�a�n`�ax�K��a�\��~g���8{h8Z�*`���O)�K ���h�awt�r����n>0z�[
�Z���$E���4�R�W'��~6H�]��?:�W���&j��Z�=I���n��kYxh/��P�̝qv8�,(Z��3*}�4'�}�P�=�3Ƹ`�6�q�ݐ��T�ngb�&�d����������̙�c��a(%�Ts`e�#����A3*����4�;�0p��g&y�bs�a�e�ۜ���m���Fpι�c5]��bS����~9Sk!����������3����a��:��b�NհK��ӗ�����wz]��ӫ0�q�I*�k����y�+����!և�Q�t�Y�\\c"⌇a�Fϝ�Ϋ:�>;e���0�Q��1͘��?�f�![u�QA�^�$u�W�I���C�^�k�3��KФv2��&���\�s���2>�|&��:�S(4�\�5�8ָ&��Ow1Y�9�{��̗�!�j'+go���6s�b7�!��a�ɪ��I^<�v����?�@A�^�:؅�J����A'�2>��]�W�wͫ>�ʅ��M˜������,������!�S�loRVPB�;^ \m:j�L\:��L�J�����yx��[o;9ݜ�������(�J�M����1຾�R�߰&|l ʅ��J�L(뇭����eqۻ���!~Wۤ;
����)�=�9�F�
�sm^��"�c%{U�nf�!6n�m�1,�'��Ƽ5��Hc���-f����ʭ3)Y��>y���W��>��s�#
���BcɔWk��J�d#�k���j�U�9�Z��	�[�i-���������M��*9کE��̓�gT�s�bYX��))L9��!J�?�o��<����g(��>ܷv����MX[��'�QiN�z�<�L4�r��SZéۨ�S�b<��;�x�_G%�m�l4�t�-��D&b�(Al��̰�B��͏(qU�*���~n�PZͮ��ԜK�B�;�v�����%�{���P~��P`����BdF��	�N�zK8b�0����Uz���߅*��J�欉eCr���e��\�np�Ve�Q��XUr�:�Q��t�UN���i��`Y��#nO	�r�"{�R���ib�5��ᕛw�_nIgb�|Y�8��r�+�-ܴR�콼���1��v[*�oV:p�z3D��O߀�z�{'���3�M�x��a��A�w�y�`:��k�\X�W��D�n���MY���W~�2����y���׀ܪ�d.��~@)����4u|cD��/����J���ͽU/3�7/7G��,{�/���}�	�y�(�s ���(!vW�Ug<��۰�T��dJ�m^첏�o�ܡ�2��O�c^�ŨH�b� m����:%�Xh�w�hf$�T&��m�j��g��� ��)}��w@H���A����{��`�u#?yh��kt������]Y��]6M���8F���Кa�j�/��ӛ�L�]����YA
�%�;��N���eg�7�+3y����ֿ}�ZfP��������p�6�J������L�v56�H��s���`�~�+�^Z���w��#D#I�[E�E���9L��j+שͦ�nlUu�ksr�m8n��4�����ܮ�`({�bኸc�]�>j|<�Ɂ�. �H:�ᚘ�i���7goR�x�@��-@��qxd����+�xZlw8��-L�����Ѧ�6<2�Z�5+�L�;�v���G6��I���ӎ���6u��&ˠ�9W;Mkim:v�CB޵����P]H�$�yOD�m��*zV��.���#��ޔ���諸�#D%���Ĺ�t���|�fn\ta\�5چnB�>�����5O���[�Z�,6}���/�0���'�G�9��1��&��Gd�P|��L*MVa�\�-�uG��/!B`Q��	�����|�K���������n(���Ck�sa�WQS���V_���}����u|�	���Á�y%6ؘ��>ܞol�TCQt���_M\���U^;t�Mܶ�qaL��y�M0����#���>��r9ƣ�?i~�+������~��<F�lغ'�5�����t��;A�>�Fs��`|5��.#��y��}���r��[y`y�#vxF{�+��[]钟��#&�n��`���m�wf��ǘ3����ۅvDed4��Uy5�V_U���61�e�vO�ㆅ�d��c��	�����q�]A~��
��9���~޻�P�"���c��eL�h�[&�C���'D?>�)��w��N]�A"e��/������9����ݎ�\�2ǖx�	����k��=�r`S%[�_ӝ�����D�1b0@s�u�_zo��3�h
Ы�ڥ��l'�@3�ߚ�X�I�=�˖7c�/,Г��6�n����J�{_�4�k�$5rҗ�k6�*VNRO:�+�~7���|�#��.�%V��u������o�x�%�OE{���q���E�,�Uy�gp&�H�G,��WN.]-�M[��"{gqA���M3U6gdA�6�y��z1����0矷��,g;-�"f��2�[���8�!���kmjO��o��;�g�F0�=ŷ�{�U�������w�/^:�t�Ʃe�1�Wdx���Hj�Ft3׆l�&���x��'�JX#�;�W��/u����]���2�'���Ym��O��;'�P$~~�ߝt�g˴���52�}=���ޑ����f�zoM��hx��1��=Q�:ɲ�_��Z�^S����0W�RXS-��n�*���#"_Q��Ԣ^�1�1!���Eä��:�Pnos�d��D�6��i����υ�0���SO+c�xt���>�4�ڨ�g����E� �؆L,WC7�/z]��ԩ2�Ų�x�ct�F�{��\!����"���Ɓ~�/��-�$�B1�r�L9� �X��2����2ܩ\�N	�E�	���t��;�����`ަ�@\�=�|~oIC��pǪ���%\?,��b�wQ`*�y+�����o�IcC�ӷ��C��%�Ç��|r.��3s���q�)o�4-��Ru~5t,���V�TXZ���jT�j����y����DLVm7�˱�m3T�zĒ���ﳞsXy�+��$�̍..�X��(����e��-��йpWBt�>��۝Zh�&��ƻw-oW�#i��
<��4����{�f]�doR�:�յ..�wk`'��w7Î���D�RŽc� ^?V`��0���O����@�,�`kd�pеnd뎶=>Z����%G0ɺM�1��'#4vs��<�^ú��@@�ft:H���hL3ye�,9�i*�`'�u(�	�e�FK4��ܾ�YoZ�;z�x�KsV�̨l>���0XCypƇ�&��4O�|~�d�o����ӵ��/��:�]#ݏ�1��-�!Eyg�Q'���x�4`��5>XBn����,��n������Wa�B�1�z����yހx9�T$PG���d^)�X"@�BA�;|W�{xJ����@U.YJ�E����Z��dcH����vd��� �����քu<7C��C%�p�]�6,����S۴Fx0Pнb9���vŚ�r��o�6��C���~�s�	Uk(RJN8|�Gv����a;�������f�Ռ�S<	���g`���F7���R������e-|���!F�z<�<�T:��Z:KH��������[Jq%��HOex�f��<�x;��%��.��ý��b�x�ua)L:pS��9�[7S�c�Hp-�����!?#.��Js,�;B�}��0��0e��.�D��z2��O^�U$�1�:0����O=��S�4j�37Rܫ�x�F�+!�R<t��Ze\����]qW������Kf<�yˉ�*�s���t:�M�#�/QqA�NfT��Tѡ�M���'P���M����k? A�����N�r�9����_x.�^��N��2.�7E1IJ`���UD'>���	>�S^���]w�Ց�gXS	d�h�H�@�(y��0�P)�u��)�-��:��y�ק��ȡ�$A������W_
��!:.Y��B��L�{F��Z&�F�{���PX��#��3<^;��2���9d�����P$0�w���B5��=)�OIo!����&eE�P�-��t-Gs�qvj�t�	�<6F����m͗�j_~�c�?r�� �|��P#��A��4�;������ޖEw������li�]1Æ�'�b�_�OcԠ�����<!t��@xN����e�q����כ5Tu�F>c�8܄��VGS�>�zc�OT��*�%�y�7��"�
�^�{c��7ri���mF���K�t�Hf��I��s�-��1_��h��%�>��]��>~� Khsќ�3�N�hz�;��L7M��V?��wWw͜a�z	^$@#�K�l��凞𱥼�]3Y��}؍�\-��xo:������V~�3-O!����L��b�~+h Ô���zW�c^e0���in�����[�j�%�>Η�>���<����;k;8/WSJ�}�{*?�m+�VQ��O����g��w�*c�s���/Ks����aɲYo�#�q֩��9�&/;L��;���qY�;Y��?���P��@��gQ^����e_� ��j��i�,�(X��Թ��#�i�&=�^Ǳ�K-�h���ӷ���2r�5 0�577����5��z��^��!��Ŵ���G���0	#�����`d��h�3�jg^@.Bu��L����ϭ=�\k��з�x��U�;�
�xaz��-/��ÊI� i׮u��r�d��o����x-`�-��q��%��>��������l�O"���E�{\h��U�5]�k� �CZ�G��6C��A�@C�Σ��)�|1��]"��Z��6z�dy�UYȼ�"�d<��l�Cy�%�po*�`�pzL������`�j��/��9��v�eك39��$LҖ�@oFk��#ϲ-� B��M��sۓ�E��Se��s.{1���u��_ss���5���<	=�.*���DO����C�=���^�jk��M7h��؋������r�/uw��_�apW�a���U���i+�������������-j�	�����2Ms�����܄i�k��I��c�o66�_��"��wf�ԃW�4��  ;� ��P2	��E�=�s�+���<��)cV��LJ�ud�`����*���S׆DpVgʹ=���ƫ��-��(e��:yQA�g"�W�})�k�C9�u	�ƻ,�v���ח�e�ǈ�WO�jT�JunF���C�(��l/��|Gd{�e5���IM��$�"��=g݌��D�֝�qb�72k@�ِ���.ʮ��5sPʕ��wNα���q@ʹ<��L��A�Gx0�L�b���/
�ko(s���X�c�;�7R�u�³�Cp���e�_������zKsR���8`��h⾡G%u��oZ�n�d�������q-#[|+��z��w5��-�+ƅژ���}��Bm�DTUM�B�N�+�!���R�[='r�g;pp[�B����Id��seYw�T5�L"�b��I�v]�n���P�c{�$<�//,ؾ�R}M}'n��b>6}ݨr�,R�X��:1�>Kۙ�vG�8r�$��]���v�3��q�چ�ʝrZ�*��O�}X�h�������W���n\��CJ�o;�k���/26��[e�	Y#�ÝrힻY*$���f��ZVmu�^W�J�B�Է���i���y�i��Z�E�|� ,�0�ݮw����U��T��b�\K�շ:��/2�՚DU�������&Zʭ�l�jJ�F�3�k�^��q�J��Kq����9T�,D����C/D���Ĥ.�Vk�J�Q�.�]� S�WP�Փ��Tol=��!ޘs��k
�G��O*��c�T��=�wf7n�Íɖ�*�cU_�7���������{)=p��y�Wx^����:p�w��#�7Qd2+�T��I��>6$�"�"�=���-�룸�9�+U\�7�����N���y=u�hS�µ0,idҁ��Ư��s	u�좳gr�&0�;�L�W��nސ�#��͋$p��{�.I#���[$�*X����3ot�p��gH"�����n�v1���;A��pk-)15Y���.�)�=I��&��R����� �ls��&���K����t�BZ�m�;j;Y���DȢ;�k�t��J��q�&��]v!.y��ۢVnda&u��B�pm�~�e�;kX�{�pU����7�1�+��z]�6;lHx��(X �fu�w�}��s>��+6��,+_@P��L!h�h���yń_e�rj�X�s�5*��H�������)��
r�}��M�;j�x����J��L�d\3;\�v���E��o3{��wY�����4��ي�+T��=��i�Nm��kŚo�ح;��i�GR�ѥ�܋FޜU�ixTD���u�dՏ������e>�6U�$͆�t��y���n��^h�鍔���}S��7vm��\W��'��ʩõ��΂�)����ғn����~4q�R�GA�
d	��E�bz���eNy����]�����6��*��X�Kyl-�1����O�OK/-H�zi����Tb>X�.�+��XbTPX�(�VD`��-�B�ON���,ekR_iTE-�EX���Pm(�Cg��b:a��vu"��j)[��m%J�"̵�f0�T*AH(�{eQc�b�+�M4���QX7e1�h(��b�e�UĭkYSX���*�Y��*�bp�M:t�F3�8�%��H��-I��b�X�����X��8�x�|Jt馞�:6�Q�!屹p��+'��b���UkAH�*�q*u�H��)Ӧ�zt�V�P����0`"�*,������D�O�U<J�YE��1Zxxi�N��UB�88�~RUg��*�S�l+�$Q@X�B.!U1
�Td1%D`�XUb"���Q�(�U��A�$��������}���[��|=:r���s���\�o;j��j�fp���֢�%t�n�Ĵ���X���Yz'\��d��m�1���*�J3wVBO�8q�V7nV����6jhǴ4�ܕ�?��P�@P�A �A�A��a�������v%�fh	��!��u�K���Ρf��f��1���ޭ�5� �PH�B�n�;��kI�f����>�A�x,)�xp��9`��6M�Yԓ�~df�W��c�&g��k5;�6E�/�e�i���X��CVS)����<�g��B��2[�k���R���v~�?3��'];����n��h���C"��������D�� ��o�k��Q������Rf_Uu�]�ݐ9��^>ݧk��Ơ��c���~kO@�Ǔ}"��h0��`����9���@xg覗�U��"#%x�&��'}rnd�p���-� �ٶX����ޜ������F��1�+��1ۜ�a���B`��
��M�S/4�7�����w����	eIuc9~���z�7�P�ki�F9gM��#|�fV>��2�:&��r�o&�}���A���4�`VhR�TX
k�	�����{y��}����d���i܏��*���?���%;�헧#}S�w,����Δ^�}sW�z싮��2u�!���}��ht�z�s�SB*��w$}B�������ɲ]�}��,ɥo*�7M'�f�'�^�����bk�p��u:u���5�����]��X}&�`�F�����.F��[�K�1˔���!Y+L�c�o;y�f��L*gT�؟�gm�)�j��ڦ$K��î�n�f�v�J�>�YTG[֜ŕE�>n�?�"""��(���~��Ԋ�[�y��-Ö�0kO�����C�[ǘO� �F4�B|`T�)ձ腚f=�ʻ��2��C;�CzlԔ�LS"��9�iyGf��ߙ��8{hA±���J�6=;\U�T����i�B^K�{��Q;)����a�B��O�T�<�]����vC�[ΣrS���3�|,���=��̂��z��u�dQcV�`�k�����:�|�����K��ܾ�GȮϏ�Ҹ}�/��X_����,�p�[$^���̜q��=+]'%�;
���цqj��Ō�P��5�j��������>�jq����0̲ok�kVrT{��<�c>��mSd���3N�	`�-��!~]�`���D��������^�$3-t1Pcq���WBv�Ხ��5����oL+�D��L3v=�fN��<�yg�Q/��u��+8��>���~�2��K�����,U��0�^E��oHD=� ��Ca�ʇP���:ᚅ�ZL�2�<���n╷ 8FRv�?K�=5�Ƒ��Hyj�Az+4PB���M�Ӧ��m4��WO�Z���?]b�l��g州��R��˼"�c9�ұ��d.T�MR���WP[T�}��-7�4�!�����Y�2��%�|�Xg�hL2��	���C7����3lV%��c��}Fj[.�_��m�	�뮜�2��Ço#�y7��υ
(Dd���0�{{���ߗ�>h������?�yv�Jxt}��-�\���`�	A��e
Up1�D+�G>�5�=7o��/�fmF���LxBll��q%�m�2W�R���F'�=�V��X����8�k-���\5]�Z�L�J�/����k�JX��s��.ODOyk�-�����/:�hsǥ?Xe0L�+D�e�k��Jz��y-������u���J�P�n�����a�`.�4 �_hW�3%:��,��eoduc	*���qOw0^����p�N8�k�-�V�gb�&mQ��З!��Ƒ*�ey��QtÑ�k���/صRą�3���`���16^���]��E�5����L�=�������]B�Z~k*lg��P������Z���|<��%��!c��_�l6�����_�:�	�c��t�2��k���)��C.��^�������]�!�������ں��GdAieT�l4\�i�m����\�Wa/��ȰC��״���yO;WRͽ)�w@ ���/�+h����/;�os������ܙ�ͣ�WwnFD��5J�����#f](_����]�\U�ne,�1J�+o=�!39�D�I��pA�&w8��`�b�]9��� Y޺5��ӕ@��`RG�᭫��%,�jN���Y���1u��5[z��O䟆DH#�B# �"'���r�PB�������1ә�ĆQ��dϧ���,Ƽb�;�g�U"E��ˮ*�E^�:w �8UN�!�.�X���3 ''���a��<�{K�=�C��������!�ӛ�@�?�^��l�D=0�a�8�D���/x�wH=y,�{y��^�c���<7��N[�"��R�O�F��Ȋq��g��[��V~��z�ݡ�~���L��<A�U5�[&)���.�ܢ&�Б�{7���<��N���~hd����s뚟O=^�2�Ҧf�5JѦk7���:o��r�3��������3f���^<��w��ڲ��Q���]Ƣy��6�fX��m鳧�#%kpc��ϒHO6�5.�.�+�Q��{i�����(t�m�)wMؑw�9�i���%�l<�{dY*����xĲ/~IM2�J4�`l��|m�t� %�6�3M�h3�T�u�����cC4��.͐���@�:N?;�t��1�ߗH�44�٥q�K��bCx�==�e�ȸ}��Ř����>��}/���uE��Rr�T%��r˧�l��Ө��*t�`�](�QӺY�wSb&h��nڬ��9�T��Eo�eD�:gU'qj���X�eOx4(���w*�hǽ���[\���IY�װ�z�9qG�\���b�y3�E&ʥl�rV�����r�>�i+]�f!�vGUb�e��S���N����9����#$D�"$���$�ߜ�������:�1��$H��S
�����מ�Ϲ/8��B=�)����7��gT�B�fxr�7P�km>>�-���_:X�%�qy�%�����^���/����gk�ݤ���F�d��-/5S�Us]�^(Z�����DwD�$:~�Kf~��|9�@F��D��s�曮�_[u�M�e	�)��<����e��u�v0�/�~�d�̨�*���b"�'f��&eo����N�/�p��F�����]K�>�b�i��X�Lϵ�y����{�/y=\<Gƭ$Z�G��nF3�t�x �i��^���B6��I86��0�H�بq������3�����0Z��������O��E��c��^����7hS��4',�蚆5Y�k6�q3�e�)];+2�ZE�=(��ǯsͼ�ȗxA�� ��ŧV&-��������Ul]�<"c^����Hev����)�A�L�M����x9�)�0(F0��I֒��k�f��/\�eR��!Us���m�a �2Pnk�Y$5r3�.6m�b��NT��=��졵�����{z����{�4�2I �CFp
�f������-(eQ�*��z͉�ݐe;�f6�l�O�t#��#׆�o^ߵʱ~�6*[�m���yB�k��byg���ι�}�K��ʷV���s�%˾r�~=A��T���C~{����0�"@FH�"0��O�{����>~��1	���"1�L܅�9mCT�Z���	�Z�,�.�g����>T�Q�b'��oO�k5~��	b��R'��T�&�uϯЃ-{b���ZkZ�~����#,,������L��C7&N�������~��?��r#����_����.�L����^�~c�qy����=+��E%QN.�Od[B�:q�A�gd��beC�e�g'WE��\�yC�2ڥ\ĳ��!�"���2�_;5��7 BF4�r��qL�5��ћ�3�A��!C�Q�,kr��j��I��3l���s-/|r'_���(��������v������z�?$h1�S�E��
'e0�e{��ܤ�~*K[.�S���εǺf)�)�g7	cTs��Х��,\��_<j+�X4�Z�HSk�+g�Z��3b�k%��J�Q�1y�9�I�}d-���8!Ð����͵&X&6M�fÙ8��Xa�Ko&厱<]���O�YN�?w�z�q�,	zy���B,xs���;3���,1�tV�Dմ��3��ܩ8uKŹSuP�E�Ec��,)p�ڏx�R����|��!��s����w\���`u���b=#�-��V�� ч2v�	(��bm���/�{{EeN�Α�"T0N�w82P�U����+�8Ԝ�����*F � �"0dI������(�`�t:��^��q�i�j[���\�r`C��0<xJa>x��"������c5[Ŧg/9�%ۖ�׈�'�{̞�]������1eyM��y"���Z�ѭko9m�^/�5-Y
+9ۻD�xC�Oy�x.|�(��I�˞)�4�.���g#uN��1m���� ��{Ǧ�nF5�[Gd^�VHB�5��m��ۢ����}�䒇���c�ZӍ[]���'UxF����g�j[`=bR\_���e�8OvM����f��z�e.�:�U�zY~�/_w*��:)���i�9��c+کng��qǥ�f�,ç4ξ�Z�29�Z4�<���=;��U�e+(�����~Y�F>�n�o�PZ-@�[s��>s6:C!ŪKW�)�g�는�5zT.�KNc׵�վ;�alo��ow�*�V*��sl2����[ϳ/�{z!'\Ĳ.����	L��ᮢ��Y�<P�y�|�VF�E��lw��z]�nƑ*�(���QtÓ	�]F�CrMCq��X����IpC�QA7�u��fN���kVk�Q4��wzn�j~�HW�⵾�ö|�q&���O,*;r�Y}�5w7��x�F�%���n,��׏-�R�v��5+B(�;{0��)�\�:�.M��V���r�v,�j-��dd�]�y�~o=���ϖ� �� $��$�D��0�F�￾�]
�b��i*/G2p���=Q��A�hQ�v�8�Ut=1vs���`��I1Q����mōKzL9j.%���W���:niD ]]DӚ�XYw&ȡcQ}�Ts����S\^t�L3m��r���St�se�9��8x��=�zG@�������Ͼ�ޖ-���dT��M�Η�a���5�8�,~	A/t�+��~����&��)�>�.m�kJq�$��7sE�M�l����ofۮ9Rc|�M���>�zc���1�b�:��wjy�D�C!����{%�S�rd�n�@N^�yw�3ʻŎ� ��I�ūv���5M�IT[�
؀�v�=9�����W�ﯺ��ل8���\���� w��Yj�B2���z��펭�:)~��7M}��~��/fߋ���v��79�f�R;��� ��m{��*��
^Ô8>�ٴ��-3?j�;�0|>��/X���k�Q������؆Q���^1K/=�!�l�!�Z�`��9A�fͧ��V���,��.���ιR3��o/�͌���D>=���{#���b���P��/Ӈ=���z����-j�#��7ۡ%ۓ�𢟈�U���W��C�4-�ާM	�ݶq�w�G&&�oP��KGcĭ;R�w����n�_A��F=}D�6�»0u^9
��K-Q�a+�Uz�#$�� A �#�3 ��=�Z�[�ݼ�є��5O��\rÏ�Q^�܄���(2j��4��*b����=�9��d͕�����ts�V��k8�t0d!{�K2�28��@�H�C%W5tB	�1,��Ji��Q��b#��zy�iX́����"%[<:�& 瀙�����}�\>�{�~��'�)ͮ�Lo�N]�nE�{z˧PɨV��ѹ:����4D�lk��6�H9.�H��x#��$�\��s^-�+�\�A^>J�)�aǀ�<����>��/��|��Ƌ�m=Tڝ^�>����_(l�-���E��A<�^���:��i�����6@E�F4�t��Ӯ�[sU?V�C��M��>+g�WY4���5�w�Qx�jF����r�����<�G�E~�k���T+�y�7g{x82]v�]^�\О�M��4��ޒ���6�cԧ��S#W��ݐ~�	����Ok�k�Ҁ�����@���0����P����"�\�a��uo�C+׸$�Xw&l�u	�\����z5���P�e9�u�W����~m/R�$^��ғ�Y�6�IY%��`6}og՟�nEV�;?8o�1�܃�7%�L+�\�U�7D�:9X�[�B�����w��ǖd�L?d���Cb;N�P�[sx�TZ�����M��
$r����6�4��]�������n����� g�v�Wwk��߮g�?��"$�D�"B�$�������߿o�{|��ߟ�y��b������GD?�,ss c%Cv�k���r"�j4kՆk/�s�	^]4]�#,Ť����f�*�-?k+� ��o�~|���e6�m�m͠�눽
����S輽�=c�Iv����!�[�Z~h���%�pJ��p̪��v)�sn�<l~�c�uW>��±�6(� ū�d����>lS-�d�gOeZ���_St-/��NV�xg�/���z)y#���p{6TU�j��_��	�8�Z�W��T��gI�F��DSe=�Ҹ�8a�̘�v�ɮk�Ѓ-{��i#/U�L�WRΛ�;h���L0[ߌ��t�C���y[���{r]�H������2�#j��ލ|�X�J"uՔ�Z�*�qw8�z�K�*���xM�2A�z͞厡�;��_�-�Su�7�����v&L�ˁx	�~�I�.4�Y}w�xg���E���rѹ69ZX�N`��6�Kʘc�9X޷2�n��O6L�"�<^2��7IV]���q���=�.�ֆ�2�<�]�ށ{�\h\�P��S�x���9ju��@�]`��uO'3���0픋23&
s��2�vMGa��\�M�}�qeB6)i]_���5�b*���ټ���=2��y6;��J�!�y��A�i87��E����>
��.P�t\��cɛS�*VxU���u��y�s��usPnlSs1�Z4��s�U�(Z�O	������W6֪�����*U-�A鱾:�@$.h�r�uux�͋;M�RJ��%���ܦ��FW-粒��S��yWU~�+g�(���2=jkɻuL.���;�I�ވo:om�Z�ۛb^3`̎�7���u;�iw�I�Պ�Ό�A{Zq*ņ�����@�3(���n�䲓��΅ֈ�N�n���ȬA�¯.�h1*緛v�,"�k���cCD����N��{΄�Pyk������L�:��;5��DȪf	�)M��}���::*�lAX��Qł�]c�q�ܔ�:�8�Rs$x��oVm�on��n�2d[]����E�Y����yG*s� �M:�&����K��Zѧ:�wGXǠA�7	4��^=��ZN6+r�<�������� �rͲ�]]R/�:<X�ͱ��ɛ��T��E5�潛jފ��Z��l�I����m�;��QШfG��{�Ҩ-��[�g���ۡ'�Z��2��	��N���]橎e���Z�:��r���oY�R��C8���7wz�my+s2��H�uGIѡw����F�]�X(�5a���Y[ ��q�ް��{���3:,f��n^1�,�|��A�;�7���&^�H�"ܛ��b\hs7�֝�ɰ�ifr��e��1bQ����u�u�t�jh��]B�g+��G:�Y��JpKV���9�����uZ�mj�;��,�dr�r3�`��OL���u�3��%��e;�d��9b��թ�D�s�ɛ�
��g&���N܊x��N�U�o����6����U����}ь��]�P�mݝq빼�ˑ*�T���t�:8�
����6�_p�:X��8-��Tt<HV��OWT����,�j�خ��on��{1�0��ݓ4�� ����C�'�o`��-�Ґ)p�d�R����I�8�`��܍gո�g`E��ܱ���^֌���Z*^��Z��7% u&j�Z�͡��Cf�\8�e�'Z-�yU
��_%z�#ӳ����7�I�k�g�s�Z��xO�Lk�׃U�%M݇,m����,,��� �r��y:�&�ŷ���R�ы�{�7\���z�
RnGA�'d�nNOgU0)w������V�@�S�Լ�X��j,XM�gv�DdV�"Aʖ�f������J�y��@R	q��A����������$T��[W��m�.�m�%d���{�����$�$�)+f��:i�yw��R�1klK%-mʼ�ڑ��띻"���N�����Pא��� U _���"��PF<-�Z�5��eIkb�d:��N�M=:O�ORs-�6�ǌ1����+�V�0|嘬\N3"�a(�����ӡ����2*��!�TEu��u8��+{h�`�Q�$�*�0ᧆ����!N+dm(��Ƣ�XU����*"��dr�{�s-�FJ��f8t����;�1�ޤV�B��ٙ@�b�YRQ�*�|e���)��Nxi��=��R(��eE�P(��,A�G��.yx�kUE"�[Y�1Ƣ)�M<4�t���V��Ě�̳R\j���bES��k�5�hZ�B�pӳ���,�Eaݳ9R�IU)l�_��>f��DX�%yK*UE��aᦞt��O劲����	Q�ml�Qm9�R��s���*�*�R�QYU��.+�Ŗ%b�eh�������*(��-J�^u��TJ��ѻ�q^�{.�������7�c��A��S���U;���Ls=��s�ec�w���q#
IIB�v�����! �"�$�D�M���������K��}���5�C�n/@K�~�2$��L*��熳P��%�[N���̧�&V4�5�j�:�&�����b�b )��u�x_Y���gu�5�Uh�c'ʵ0yY���d�4Ϙ��X�5kۇ�k��>�y���
[&�еa̜qр��8��y5M�%�!�ņ��瞙zS� ��M59�K�|
�����1���0̳X@���ĩ� =M���0�YG���L���3N�U-�G�Yz/b��!���`?Lި��+��K ��[Ol�f%����4�&S��	�nס�}0���5�-���N�Sq/Z�i;���\�U�?|7�0�!S�QY����D��R������@G��zdjʦN֙��f;ݨ�U�׆�q���DFc����Ƈġ�Ǆ������c���� �;��w��!��D�h��am﮶���s���+�h?|�;2J�8�ϝ���I���s�T��3w#��ԫW�"ux���*�ȗ�:k�5�L|����s�(�J8(`��H��c�5=ۻ֎�C�8���@�v�<���/�A�*�&�>���ma������8�rl#��++�ě��~������tinu���mrV�.8��*����
Oc�l��7Wj�F�l5�VA|;6�͑�2½�S���#�zFnP��|'�d�#A�� ���3��0`=�0���F�vI0���o���m�2*�
Or�(]��נ1��@��v�[&_	嵃[�����yҨ��p��5�E�j�B|���S�*SC&�EP���Y�~׬xOB��*�$�t����ɐ�U֞��B�	z!���^Gc@BE�H�):��d]ctS����8���Ն��)	���\�^ډ�����1�F.�'ZnvQ��}�l�`TŗHs�1�צ��B�N�l�W�SrO��_��oG�
���n�0wa�'N҇eOC�Nٜ�קj�m���ik��U����2�.�k�|�I�X[�?�/���=<���:�P��0�ݾ-�96�]��-U({��s$R���@�^�<v@qF�c�=�ér�L�ڷg�z&��e,h�'i5�~���o��a(%��D@��eW��1}0P�!/���pɸ���{|����k���Pe�����K��e
�m)���*9�OK��LXgc�Z9�t,���ۛ��h3p����jj�V"?-����}�׫��y_���ey�g�|3�'�Uqλ�dwo�N���y�Z�Y��
��-ީع:�aͺ;x��\�μ�fOۂ�6���߰^�>�I�-�>!+9��͝�2��u�h蹋�Z�"��CC��c��{1=��w.�H��繙J�;�{��0���hB+�'��UW�� ���2��D��K�"I$FE ���k��7?~���>x�&FpЋC}�b��bjL,��	_JL������"a��~�ﶎBJQ���;�ݗ�gYw����Ԏ��iƽ��O��~0Ϭ�ƚ��ʿG�z�ݧ�hn��	_v�_gKnu�iAt���CQ�E��z�<���5QLP�	����?<yK�t�H�a���Dd�t	�idl۞7(1�S�W�9A�ٳi���P"��0��9�#8Uz�vM���8�bY�2�u���L�\6��=˃Rn§&�bS��t�
$N��Ǫ�r�ݰkUV�!��w��5&�eD	A�l.�gt�8�
t_ɦW(����6*�Dz�V=�(~�ej��'1��>D�` �ai�X�i^F��'Eш��vk���{��mZ7|*�Մε2�vO5y�.���Δ5���)��aj��E�U)��V`Zw�m������n<6��r6�(�.VsȥAmsj�����}�4[A���Hʒ�f��]�g3����/1��^��Iu�S	��jp��1i��O ������?`b'<�
5�{ҏ�9��z�G����Z�/gU��:��b��Rv���x�'O9s�����¡0V��nن�Wɺh�;�b�O"\�Y�����	S��L:�;�U4�S�ٍab�n�3��C�E�{kZ�����[2�T�.�(�k36���]9p�Ç.pۆٿn[���)tb�2b2T�%1�&1I�U<<<&s�J��+<�K���>�D���]���/jG2���w='�t��v/��\��l{T�]oZ1L�ݘ��"u�	�)��Սw��I��b2m��J}U22f��v������wuMX�~h���XZ@�*�@4u}��఍Ӧ�+��ux1�k,��c��c�֍n����,���w7Y/?A�t}x���X���:
�_T�({��t��f�.��Q��2�wL���m�8¸87A7�E��֢�������`PY��9�01���[���D�m;f�n����A��oBh���e���'�DY~h���"]�����؟����Y/�L��T�sn�׳���[ҋ�%8~���0Zù�"���`�����k����Ң�)\"�5���W>4��J�H8��bԖIQ�gћ6��aN� �K\���Մ�Zώ���'� ��C�=0���Lc�6PB}k;'�j��α�5v�Mm��Ɯ����2��
�{�EM{-�|1rÞC+��r(o�O�n?�_�)�O�k��	��.�^�^�m<��ǄJ�C�y��S�1����8`���.�5[ϯ��!�z��tR]��{F
�Pc��H���e]wz;q���ˀ��t[��=8,�
����&$��u���i����f�gd�4�!o�|���p�?�!'�"@"2$�D�I �HD@�"�PlY��|+X2�}�A4+T�a,���N���=*���|���A7�v4x
T��X)��*3Grv�Z-���M���Jsi*�J��^GN0�ض�Fq��ҠS�����Q�����Ǿ��yC��Y�l�����T�a{-S�\h��/N�x"Xn������_�0B�6k/�o���{S ���!�Y�n�'��-�L�#���nK�ӱ<���Yc������I!�~t�����ݐb_D���{�Уgi0�X�9�Y�I��RX���j$���D�\G=T�a��A�5� ��/���yW覯��B͹��.�TX>6���-�8sI뵮r�/!km!{^L'��O�C��CC�`�C�w�[��LhN	�^�U>A�	���D�X3Tҝ�9�����F�Y%�&�'^��%���*9���:���C�8a�#��D��j�������,��}M������3�@��	�i�@�~�ǰ�3N�nm=��{���z�bZ&��IЖ�gwcu
�'��u����l��¸ĕ�"zցޑ��Ϲ
+���|-}^���2���3՞��̩�)��S�X��{�4��!��>IfJTFA�P>v����U�]��ZL)���p������P�S>��<^u�ft�H����ȶ�׬����ڽ�ǩ�UkL�H������ۚ��(Y�xW{�dCR�a  �!" I�	74�s�߽�Z��	�,G'�)���GvY�[�<��C�Pi�.���:�tJj*v��m�;�<�i~ӟ�Zg�k���U~��2}���~�P�P~�+�a]5M�&�
�/!
׆��-�.5��_r�^�`?|B�,�_+��nr���P�л�al�uM-��~��s�c�+W"R��u��ޛa"�*��3�BcN	��!�s��Dcɞ�WM�Y4ϻ������ux�KbD&�0-�'ݔ/���-�QYE�<�����q�f
����OHG~�^�����|���Є�0,�No�J`T"�]�2s[m�=��m�O�NT�SG���ރ
enH|��By�f��FI�f��N��d]g����H�aJ��S?I*�����������x���Ks'�rg���cH�B����EL9L"�wR�qש�C�GZ�����jZUC1���6�54���>hy��}08�R����a��KwU\�s/��1��l:9���x�,k�t�~j	Ļ���(8�w�75;OTs���W�~�yl|1a
f^�^g�V����z
c{�������72pi>ѽ���b�-�u s�o0桷3x�ښ8m�,�M�w��`ͩ	yg��QՓ���}/t�,�#L��d#2�n�vOv\�ʏ.�C2����;��l�k6{�$x���K���V2���2��c(X�V2It��˧>��z�k���3�b��
�vJ�a�Z���k-P�zղ!�����d�	�>a��,���T��L�9z7-`[�a��^��kb��q�Y�P��<��o�Գmt[�:J���D�L�B��n�� ���:"�ȇb�vm�����؎T��������GG	앣�ܪX���o���[�����x�,(!�"u�˲}���"�Q~����� �i�-)�=��ա鹖؇e>�x�X��p{P(E2�/���c��!��mc ��Cuݭ��	ƙ�w���/��C�4olG�����]C+�Y����"�'�z��<c��GQ��7�*	��ܖC!��L�^�è���#&<�ٿ�~�-3��V~>�U�eN��U�)��h�+��l)f>��A���5��(�Y=�e5jq�j(���6�����N�Y�0�媡s��W�p8B[CV���I�mV0J��H�"Sm�7�zњ�{��a@��|�$9����IE ;����l1,"3�2�q ��������'�1,��Ji����C�p��3�(����'iY�%PÒoe�B��L����q-t��Ԝ#a�,�ѿ]J��7h��ZD[dY�4�@��3.�V~���`X_F�V��Y�i<�:Z�׹n	���s���]T��m�>�tmR����$p�>W�r۟� O���FA$�!V1%�����1U7����q��Z7
����|j׶~y�� ��Q%ٲ��`�v4�/���'E�ᶰ�mܽb�0Tww�!��k��2)�iXv6�'X�~C�Q����'���;"!?�Z��u��j�5cot��0F!�J��1��h��k�Ú�����}��#������:=1?��3��Tm_�z��`5���Q{:f˦�}�&-?,�y�.OB�_�M��r�{`c�o_;�䩲&z�v��d=�D<1O^�3M�ګ�E߰�/�VP��{*	zK ���|ER������,�x��Y�p.)y������_�@�u���M���k�oJO�c�o2��`�V���*����}�<��\/>��`h���p\D	�'��;S��.�� nu`lX�`h6F���}�L����[|u�ȝ��糏�Gè4z~߄@�`��W>,�ӞU�d���U���S�{;�P���P7�n���d�y���ߘ�+	ɔ4.(����?�{>��&{��[E^`��dCΒ�_;��]�����˚����)t�����e)��߹��ī���K�%�bOFU�狫�^��y��ũ͵ןE3R�0m��"nԡS/t�K�Ai͑���4�,»-3J�ճ�#���v9׈�:�fh�&J�����@�8q�m8��@ʼμ�u�A`��)i�����{�s=s~|�y���w���D��$�	��BH#$�FC����B�&C�M�iZ�DƔ!`���s{����CzO;R\+Y�$�G\΁q�]D�J��}\�E��Ϡ_���8l	��!�.��>]����k|�(�&ū�d��
3��E�w�(hڤ�Zc��lS�ʟ����Y�����I�1�	��M�ȫj����vE�~�N�}�	Y�4�w���u�,��}ϱa��)�_U�J1rÞC*9��dۓ�E췭4ɑS̰��#:c����3�#q�%\�LdJ*�E�2ڋl�.W�q��"z�"�	����c��'tuW-}�sx��^ޒ��Ad��&f��	*�U��5�(�cB���zB�f�zY�4��ک|K:4;����&����m�sѯ&E�&){�E'��@�t�}��æS��,�J�!��ާ���g �b�[L:���!�v��}RS͂f����6r&Epkc��\����n��6s5=��uמ�&�z�c�%�n������4(ߎ�aU�2��Y�I���m�E�f��q�s��I�42$DJ<*����vqz��u^�4,���*�g%���Pl^{z�vh�boe
�z!�t�&P^	h���t9�.��:Am�868eP�;`�������A#�����ɉyg�Y�n׮�}�K5s	�Qf�R����*c�9b��$^���X�wV�N�J�S�\��qoFb��l ��?��$ D�� H#�$D!@ � �I��|���|�Z����St�X�}l��1��Q��c_��Ӌ�J��"��;��k���m��YA�N87�=+^�PK�X�>"���C���s/��P����!���ez����ŏkW�d�����i��@6˪��h�4�{�KsP=˖��|�J\�Y�+7�ѡY��x0��A�6�na�����n�4�&
a��÷k�R�C����m1�Hc�лʯ��j�R�X�Zr�O�N���{��"�/�kzA!�%BF�f;JV�n)���w&�����B��=���6��\3X�	A����ؗ���P܌i��Y[l��L`��Ak�O�n��u�&p$Ȑϣ#-�t=C��Ͼ���I��ofU�ߦ�(;t�s�'��m��1����J-L�\}#�κ���)YTu��EMF������z�8�����s5�y��N!\�z1��mT�5y�	M����+�I�h�|L�=��"����&♅
��7�o�[�^s ��߹ė�q�`� �|�O5t!)��_��u��0����[9���X���ke%�i8�3�1��f��=k/Z�4C{�aF�2ÜԶ��g#��&i�<�R�]2��U�E��z�bx���Қ���(U�y&�b�>��T]ٝr�� ��v��3O%�w��6������{S~����M5S�F�s�As��YY���%�	i��3�UoA��j*`��]]d�o_Q�� F�mj�z�HIH�CeE�S5�wR	�FY�",?]\�(L��޴��0�gef�ntK8�(/��?L �27M���K���W&c{h�w�d��R��ά"��+.����
ݺ⽩�Jn&zO=S'�%��	������.�e������!Ӯ�Q\��%�EVfJ΂�	�*�%�c��e�}|+ {sB%Ef����!�0t��,��o����p.���yϬ��Usqe+3s����縬�gJj��ܩԓ��>�#�.;t����i��2�j��]i�x>����OW�`�X	,Ϲ����d��e��EW٨�E�n	��USB��+�&^�<���S�����NΙs���p���=v�a%n�X���_�QlA�V�k+.��,�]+�b��Y �=�^N`Rqvv|k^��e�<��o{y�w�|�K�n�\�����S�>�{&r��$u<�;���3P�s%��o�����M2�N]�SΏ�}�7��34�Jt�����r�ξ	t/TRإƻIVl�tT0��)D�7����>�ۡ΍2_[0��0��or�b��0�zh7i.5g|�z���t�J�n��N��n��^,�L�V]�x�4_lc^dƔ��Yͪ�f�W��qvt\���p�s��j���\N�����J���s�Kʴ�=݊f臢�w%��N�Wٓ!A�z]�8&NNEM��dΧ2V�'wF��9�N:4�W[	A	6�sïz��`�Q���,�� ���b��Oۛ���uY��������{4F亲���q$y��X���lwI��I:���#Ե�J��g4�uɢUP���� ��(����e�n�D�nl�<:�G���}����N4�f�^��uܠ��A­����l�F{e+A�M8ӽ��/������Ayt!�����x+5�t�>m����
p\{yhfl�`i�pt�5�i��wO��K2#�m�����s��vW=�z
-���f�����i��e5��1X�i�{�8�iؗW�*�,�SiD�&�p�)�6�yp�N�����Ν�l�l��<�l�-IGs��YX�ngl6d<)��B�kSf����c��W�:�;e̚11�)�_W��G��@F��b}w��!&5�WS��q�i.�6d:���sk�`W�j4�م�P���6�۵��RǳM��d��BKLK����g��r�Y�v=�$'K����f�klt��[���uKQ�J�i��o�$����fT=�wM��V�t[T�t�r�QY"�(Z���]�;��������n�	�	�%q��,B"�0(�z3�S7�=^Q`���22+Z*��DH�N0�G�����X�Rk*��4���:b�U���i
�р�TdYE�J�ZP��	�U�a��0�H��^	ӇN��"�E_/�	J��Lh�W��g-�ѼJ0�O���姴
ã+mZ2)Y�O�N�R�B���ŅZ_�1�`����p���8�%���hɂ�����9�+xۙ�<C�QJ�rX,[�Lp�k*(� YYl��9څO	��)��\b�`"��)
�b�B�V
	m��,�N�xp�ӳ�5��1�
�5�1aD�9y�TaRW2��Ę����V���,aæ���-�Lf0̢�h���j
�g�DE̳�X��q ��*L�

��'Ҙt��鏎Z!FQYQ��")�֒�j�U-�)L�*Rҵ���ţ
尬�Q��ZЬ�!R�keQ#��!�
$E���2ғ��v��q���M��8Ǒ�3j&/n�G��/.��E���(��ζaG����M���٩�k��R��![�[��WU�K	2sTw� H4{|�9_	9	t��3�ն�->{��]��;>w��s/�B�BDHHDHH"`H�"x���P��ȇf�x�G�=OM���C�h.�|��By��|g��	9�xc�StS=��X�C�iT_z��5*H�-w�R��S�c�'�;�'9Tr�v4�T/���E�]0ij�K]�5&몣���F�zY��S*��P�@Լi u0�>2p��?�4>=���(���N6�ݘ�fl����Ƣ*чV⮇������Ƃ�0����]���a����������7z�T�0'��;���x�1��!�e�	Q��Q��lW�G�X�X�� ������*�i�ꜩӼB��|��݌�jb�Y�Ň=+^�PK�<���+�f�ͰsZ��1v�N����
���~�n~i���7:m��T��eO�L�q��y�C����FD��y�s�R�N�5�(�?k�<<�cC���MY�q��0͕������PҞ�2���{m췡��!����AA	���b���z����xQZ�/x�wHn.�9�a�*���&q�ta^D@"}ǩώ�_�[����?g�?����>���mW������36H-Wl��
�����Cr��c��}STڌ�ځ:�Vf��s���Nw����Ͼ�8g
�]�Y���먺T�+pL�'�u�I�P=��;�+3��|��`%�z�;u� 3���[�'��\�ӻ�ܝ(�2&1SK��T$@B߯|��|���������>(m����f��K@��#&�۟���'��6Q����s������N?&'y�R�^�����'�{m�rTͶ�ڭN0-@r��͛OC��02��b��)��QTFXBa��`r\���R�A=kV6��;��ټ�MBњObWN0Zoq�͸�C����O�W.��V��߁q��%��@$<��P�U�^�q\bYO�,h'ǟ�W��~Et�=馒�V~����<o>��iݛ*a0R;p13���cǂ������g_5Qr](��K�N�����#�y�ϑp�<��`�ƩU,�SYl8�6����]��3,/(`T��q �4�ሥ�+9�R���9�ǣ�|���B=����g�q
͓x���$�p�^�T�HdJc/`��������H�]4�O@~��9�v`�<P�mFȰah0�Ƒ�8vvZ�����,v���(�U���Tw=��:hdmI�a�a��������ݵ�;�Ct���̠AF�N��="�hz;���oJO�x��y�b�	Ӵ�g�2�Y��g`[��ce=���c�.���Sx�%j7�h�9�����2��2q��n�2@~!�ͨf�P	�s�s�w�Ke�JVupcO�3󛚍��<�C�d�6����c�/)y��$��;~o3��>���y~a��� ~ F@ �`DID	/��s�%M�6��%�`/}��e�͒62�n/���Y�m|���̖�q��T�2�6E]��ɛm��S����K���&�k��0Bb���^��d��t��ȵI�@ӓw���D8�����4$@�Nk5g�����Lh|Q�7���wy�(���fxGm2�{S �[�_Fv*C��v�-��Q��q'DY~h���J����T���������x��	n��&0��1"�-�z�}���[�����d�&a�[�Zy��p}|PF�d���j�:��S��(�i��ȼ�G�w&�V�A��A�rY$7i�n�rt8=]���v|%���������:m޼$`�>�	;�c����&�8D�5�1����o�h�fՙ�Dԫ�a�-�ăz�`Lv>5eEÚ�΂�pXs�e��F�i���&�<���3��VK_h�Bl��n��쨤�i�)�
�AaMAnNH1b��Z*VF�ǤBoGA�}�N.7W�1��oeQ����z�+�-�]�'��^r��H�TS�~��&���f_M����F}ƆY�ĕ�w�ܥT�8����̗2CFJ��
�eX/�TLU�+s��NKҤOc٨`W�t��Ua�-+]����f���ük��Q���|���A��F�3WS49Aaw ��L���
(�9�zy�������3� �FB# ��� �#	��}���B5�������26���ޗi�i2�^b��J}K�qӘ:��F�.(�*�f��}��݉����0px`�!?T�#�{ K.�pS�T�z)����9�����f��&[]�=�V�a]r�P	q��l�� �ڣ^�P�|���'A�L*����e�TD�y;B�ll�)��f<��L�ܷ��H	��vh���8}j�&�	��	y�U�hY���vf�f%�^ KmU�\Rʋ
�hr�e�XG�ŧ� �j��!i�t�%�-ץ'�#/;��.�v�ܨZn�n;���{�S%I?��sѬ%u	֯s�K��z��4���:�����?o��g6:�7b���Z���e�X��a�r�ƥ��8��8<ߩɄí-t뷾���v0M �ؼ�HO�:��,�+�ٗ⢓����A30��T�o�L��f���W�L��p��":�*�}��hy��5>XE=0���Hb��y��A!�܎Mŉ|�x�Ÿm�1	�{��T{9i�W�`��`���=�$�%���rq�x*wMKRa�)��fw_D�t{t-G7I-[�GJzZ���1s�e����1�m&aA�,'32���[S�i�@�E.��nv���qY�2gAo'�r�	��i��\SR��-iV;��ưܑNaN�kEwRКfh�c����7�R@�� �	 D FH"D�AAH�?g����>w�����k�%��$=7�pG9Dd�;�My�\m:nj��������Gw+�<�$y�t��Μ�ݑ'�X�R�Ę�ve^��ʥ����
��e[)�P������o6LɈ�l9�3�Cj�BE<�m���g��Z�����;!2�dJ~���`��z��s�k�]D̥|1e`�60��� $vW�i�S�]Jc`����	�L�J�hx��`���Cb�Ъ����(8h5i2(���L���V�z}�2K�^��&nM)��/��*R��"��j�3��_!A]��N<��������A�`��}E��/��KCEV�9�KOnDN�V��vG������<�Kƿ$�h���Y��ӑ�^�	�*sH����P�]���/y�I@�P�֕t=Y�O�eAc^]&�0�{;�����k4�׀�����FZ����|��cZO�cX&ф��qTa�Z��3~�D1.��nON��`Ǚ����V����E�3��`ݯ�b[;I���gO���{��̧�s���;_1Bw�e^~���	�:�^~?�Z�_n��Qf���C���\��R�������W{�u5�s�_8�����;Է��4��?��C�&����vx�OQ�*�_^ض�l#�m�4�q�(�Z�S�N��ֹA3c��ʏ`/.e{�'�wߜ���.��I�A�H��# 	�"I�������y��_�Ǡ �,k	�������h��2�Y��*M�a�u>߉�N<�b�fk����NT�o\=�ƾ�f�NvTg!@x������D~[3 ' ��yu���ʿ��c��fcj�����+�tE�j��g��(L'����l��{�H������7��sd�w>��e��oQaK�I�8�;�O�Q��xg���-M^C`��z9X��N\-ޫ���ۗYK��B���߷hkH�Φi��L��hч�gM�-�Y�o����q������;�����c#)�Lz��cH\�3m����������f��U������Q����i�j૞u�����8�.��W���Jm�r�5Z3I�b���h��9��k9l��ʿB�ט����"�k~>�kC�dD�C�+�`�������5d�I��@�P��l$5�-��ot�(FSz����\��?�X�������?��n8na�k�jL�d��������Cbi{ �Jsa)�#)��z;$H싇\��85>�k�t�V���t�%�]FP˲����b����VS���p�nM'1X�o��f
_~���G(߇��~�,;�3�¾���;ѽ�[3��\�Ip\B��h���$��*�v�hr�Ԇ�wȫk\�=�X���s��ϝ�����n|���O��Dd�22D`#`"@D�4�>�����>�y�P���w��K��Ω'����)RU�9�P��FO�GF0���5AU]�1=��H�!y<�-p��ܑ8_�V���1�K��bq<,�yӜ�mx���*�AR�~�Y�� #�+��#���#L��g8{G��W�����1�����r��Y;:�y���}���$>M"��Dh�=`���q�N
��jE7?t�V�N�kѲ���m�
c�Y�����q��tZ��uDх�D�����o(>_yP�'6��T/b�(|�������Ԯ��f"���TG��i��^/A� z,�����7M��/��ӳcNΪX�d��V�I��i�V)�6���P��LW6��ڼhZ��|�T&��m�/�q+�#ZD(,���X&7�����B�ėg�i����q��Yz/l���ʳv��m|�'x�C��p`D��yg�����́�>�^_V���yڼ��Q醓uV>JOxyDL��M�Ϫ�q�c�<j��f|
��<}�1�7?6�હ�Vd�HY�����y5�3%r��ߢ����ߘ�j�~[1xv�.��w��R�L,X!�@�7��	�D�w��y�}�:����ݾ����D���P˕�k�v^M�sF�+**�iV�b*�%񡛽$W��α����ѝyj��V��H���[������? A��F## #"
 ��5:���B�Ho�a��y4�]�Ҝ�&,y����5v��\�Q�֌�e��Z�Vi÷�E�%��>��\C�V3ю�똨s[������`�N���%h�}PNF[mk˲�ث��Q��df	zsk�tȬ4)Z���>�xsQf��/���n���O}�*��^����i�D�JnnwL��xO�$�*�%8�ض�h��v����ASZ�ۚ=|0Pem�l��Hq0�2ۇn���H�)��%|�)=��<���{�>c)6��yu����/o���xpZq�|�Q����!�=�}P���8�E�rR��v�����~"Z����v��A u4 t|�+���*|z{5�r��
2�����c[�\l�xd��L�E��#.�3���ǟ8q�~!|v��y2��Y�m�(�M�-�<"��A^�+\Z*K mt��J���yY� �H&5
�Xv����%A'P��[� �� �*�����.q�zV�NK�*9�����W=����0���R-���䕕����=���FR8!\T(�fM��4m��I�t��X��GE<�������Q��H*Ļ8mb�����{����Xa�x��7(��wU��Ԑ�nbۂ�]gq��9kݽ�8V��#��Et���B�L����W��B��Q � �A" ���⬤ax�ɋ�p��5n���:O�?�veu�Xќ�D��%C9�S,X�@��Z�:���d4]���/�
�`��|�|�~�/4Oִf6l��E��������k���g�{"3a ��SqL����|��C�y���T[#{�� ^E�K^��Vڝ��\��!��GCPDcH�xcY��q�Yq".�Or�����]�=�^7aF:����m�Pׯ�Y������4�m:j鋇ֆz�4�	:N$�6��ޱ�_��s:��]Z�t&�OWd��ƽ*B��A�Z�P*M�|�&��Ϸ�h�_�IA~�W6�O�,��/��8��0����R�a`BW���D��ё)�J�@�Ǩ��:�$�=m��\=�5�ze�q-s	�U�o�*�:��0ħ6
��7V��eV�rE�®h�B:s����=�����y�ʘ	<�ƀD��锝:Q[�Z`�ںX��gs4���t8�2)Ja��|ᮢ���0�r"�R�3"�3�֐�Ȍ���]	�3ѝ�u8Do�Y�xk��+�ϳp�n��P����R]YG.�Б2�Vk�2��׀��������u�GWCm��~ܒK��N�MFr���5�u�-y��	$�ț�mu6�e�+e����t+����K��qQ�]}n��"����"$X��{�ܱ���B��Eޱ侰�5(��x�N)oX���-A�6�zh@�5���	�5�V�Wg����Տ���!}�(��"�O���z����ʂ�t~d���d0�p�im]�Y�d���!�+b�a�����i0-ZVP�������1@��Adi/N�d6�yA��e�r�_�#1��/`�]X���S�)�z;��o(X�2�^��T���"���r��z����tkS�!���X�_aڝ4óe��/��XʇPc�=�Knk�^�o\�i�s�~Zwc'L�k��9���(֜��&��`�k~o�O��N��	vG�i��K�)���!Ϥ��XFW}4Y����IL#�
,���&�7&5�&�wu�F+e?r��p�0����� �u# ��k���)����Hp�>9�"n��5�֩��=��Kս���2�87��4VPA0�oP�w�KL�r�osci׷o�e|4=0�:D���~��G>z�1�.J���!� ���r����`{��nX�-;df��ѕ�x@�=k^���(����h͆o}���O�6�0jm)��R��$i�ӽ�k�K���ꖨ�9!ۨѸ�A����r���{�����1Ѱ��o�k����v�B����@^6� ˫��p�
�`Dw`��woG�����N��5���
����7%��s3`��
���y2�d�\h��R��DV6�`�p�R��g�{�|yo�ve�:]9��V^�d8��X�H��d���p\�n6t���	��2����f�k�쑸ޛܬ�jª]i��j��37��2�CyV��ցdKбOn�:U�o�+�xv�ea��d_-�k�Xx2���[���L�kB�]�Q��/m�
�\��0��9�Yk-c*�"�7�	�kd@��@�.��13n�V�t�\��n� :�R6t^Pޱ{:WM:��R���֥=`C�;�ކ���z���.�Qm>���V�k�Z��:0M ��S6�[]#��@i�q��WgձK�C8V�/f,�{�4wgZR�M�l��r�̈́e�C�.��]��8�5+�P�q���t���S�14^�
�6L��E���[�׉�fEO��Oh5�e'���(�F
K�{[5ؘ��֗�s�V yӖ�a�X���s��n��#3 ��4�.�#9c�j	� n���="�с0���m+���w�`+��E���Jdԩ�k8��ّ�ݮ�����e�ܡ8"LwMi�u|̛��-Oۖu�ǝ��t���aw}��`����-�����tQY�o��uO*�.��PJC�E�9�l���]#ܳ���gڨ�"���b��0�gia61�+������7t�x�r˸�x��Y�p�b�o�o�ʹ���tJ���V��O���i;�	�t��N�b<r>'��Um�l����pF��&�kHGM�Ժye�5�0J�3C�����e�����a��u��E���fh���������Ȉ4�����n�u�K��$i%x�m\Ū�8�ꗝ�;�u���,�n%�ޫVi,T�0Mqb�}nu�x��.o,�A�c�]3�L�x�s�*���p�N30�$���p��X"��u�����x�p���m3� NC7�m\�����e*mQ�n>YM��d/�Al2v;u��&�'v^Wc�2��k4���a�!��H+f<���YQ��C�Gw��4ڙ� ��X�}��X�ת����.�? ��:-THXs1��bd
��"mf&�خ#C;'9-�#n�d���]]�MB��Ö�}�IS�6#Z:ݝ�&���W��f����Y�@Om������ۧ��X<����e�� ��]��b��t{����t�e���̙X�s$TjfPnVE�ŗ���J��{0�e3���N�r�Ł�M�.�u^�V]�Bڠz=�;u�V^�W=��k��(��#�u��M��'Q����x����ɏ�*�،�S,��A��D�E
�%q��Jʖ��!U1`��bt�����ګ"��6�Qj
TV�
V,{LH���J��e@R(���FA=8zzt�R,`�i�m�`(��6��dP�k���0R(,Z�P1��ѕƉ1�Z(��'N:t�1�01Ʋ�%g�}���/9rJ�[U@-��b�".+0j,Ym������ӌ��P�#p5�E�[+
-�!�p�����nU����	m@X*%B�M8ziӪEMg��UQ��f1CH�RT*,+S��Q[eq.4�1�"�e�*�	���ӧaִH����8b�$�gNqmb²�H�*b�a��R�8xt��B�z� 9g�"�de�`�"5��0Ĝa�
�ʅ�s��Ƣ�X(,�ç�N��U�KDB�ƾ�8c�FFe�ܳ�;l��c�d�4���S,�E���Q�r��B�V8��9j,��`�����2��!v��geS��1��V��R��R*kC�Gqm��[E�V�J��M�T�lƖeVv�Ƴ�Wr���l�a�?��?
�Dd��cdF ���-s�E��>B���S?~t�w�aŴX~/鋏L�L�o*D׫Q��T�ɦ�*sM��uۆl��YO{�l7U��Z�O�B�(|>��a���`j�
�J�fYPFWA�v�E�*�#�g^�\ �Kj{)�ut�
��[Z���IP�C�?��'(G�f��CI)~���'+w�s"�!{�O9w,�(�b)9��Su$i5�������� ��#���Ȇ���f�O5>��m&gn�r����*z�$�Bb��E*�U�9��az��y���b��l�k��+"��{��yЂʦ47�r'��0�-�$��b��M����5N�e�ak���,�h�x������Z$i��F�\T<6���Kwb�&̮x�2(x����w�{����YN�˸�n���y�;(�g�1���?v�����>궰(g�Ѥ�!0��N��m�������� �CcH�"��<����xmls�Yh�&�;��J�ݍx�_�>,1�k,{����ZA}���A�� ք
�����K���~��g���^����xɪ�fZ�\��� B��U�n�%5�nnoruK�-�9���;�v���c���.z4��Qև4>OR�W/�����-飯������᪫���(�
4�1�6��B]<��<�y�dP�W�z�xP���"���߾}�����Z֫��b�=b���b�Rt`��;h��b�n[A{�<y�ts�x�+ii���o��2��)���یq���ב���{�Iv�e����88������{�NnX�Lމ���A֩��cE�0;Q��ڳ�/^l��������v���"�y��ɼvO�֓�]�����v5W�O�+�����ؗ�U\��"�A"�m)��t�Ñ��3�	�V�a���	29�i�e|���ڃ�1�}�]�"�	.�n@�VV�mx�1��l�T��y���tJ	�8���K���q>�7.u�6a"��8�.�P�5K��S���:ū&7��0�N>�2%2�F�%3�2��k�;��qTsߧ�8*cuA�ϵoe�;yt#���u�+����)̀���B��]�6q��hL,��P��:H�Ս�g���ϮP��rO�����ޑ}
S./ &*��"��ۉ[��8��ۭ��z*��O�z��v��z��B����� `��q�{.�M�~)���#|0����_�\aV����j	9u����VGUN?)�ϗ��I��F�@�����5Y�Q�o�}x�$V$ݲ���ɚ7kWh\�ȴ��I�X��G.�d�wo��\G��V�u3�zp�ؖ;*|uRp������&?��$���AF"~�ߚ�߿��{}��yN�x?m&V�x�=4�{��l:}°\4+�/^D?\�%�t��B����K#)ET
UN���Z�0�ٝxe�f�%~��P߽H��i��(CY�6o=�"��s�ٷM��o[��Y/�[@�A���,-ts>�Z�@/m�>�*Ai�K�粖|�PL�q��Wo0N&0z��z@��d��ҵ�y(%�Ts4'�K۹���"��]_Zz|�p�vd �f^�q�"�<óu�es՜�l�k�0'(q�nc��>!��[�9�5g;
�7]{lCu>�	_�<�z�4��q��g�s4Km�J�
bK����l3b}�����m;W)} �l;?W1e|��\�6г�PyO.*-���fWH��&�H��=vz[q��0��r�CH���N�N�=�1'�ߐ����N�����S�/�~{��G�"yU9d8�4���Z�ݲe謐� ��4��i�WL\>�V�er͡z�}N��[��c����k��5bE+��KkP�R��A���x�8��fͰ�\�C��z�C����)�W�����_�u�ݘ�]P����[r,�\ª7n7G��Z ���~��=�0���V@�z�,��A�����ڋL�z�ۛ��Is�e[�"9�h�93"�
�՞fS�� .m'�_[��N�1o7��۾���b�H������ϴ��R���@���`��̞@��l�0����i�@�!7�_*�\����}�ί�$�����x��?��7Y��ձ"�0�� ��|Ce�j�BSqxNǻq��3��U��C:�0��<z�X����r�)��Cdȇ��	<��� �Ƽgr�S����*�;:��d��9ᴺ]�%*�׭qϗ0��È�b�R�MS����^a��1y�`V�r^y��R���<S*[�:�sb��^ w��3
��yɪN��%z+��R҄�-�s�Q�v�8�����'�@�,it�~d���}����*,�OXk���h����~(��<�i�}Bl�9�9m�C�|n�27dB s5��L�3��tf��t9@x��d��
���j�OP���V·��t���v���2zE��#uF���y�/lԳ*�n�P���w��k��w6��+�q���;12��V�2��.�H��S��I���f��A��@��4t!�{�>�|/~�d��9����6�/����}�f�Ɵ.�[n�ǘ�L���-�o2��*�Gn����ۜZF��o�s�7ą��f�Γ�����0��!ѕM��Ǚ�4�S+���Ҭ�FhY��V��u)�2��ʜ�KT�@�C].�$���J�dݫ���w�|�y���� �"�A�0�˯����<�0hy���1�r�t�t�r�>���F/�T�M:$��`��0`t\�������%�ݣ���H�p�K�*��A�s�CHބC�"�=N>L�jMu���Fe�_���ߧ�GÎ���׏�UZ�X݂�K��&P������ǌ8�ش��Pɉh�!���Cը׆^��x��--> ���ӛ��Z��tk#�Y�������0d%�n��* 5��:S��(`�g=]�Ëh�輈#'�^S8�,��`�"Sl�S�d��U��Z�ԛE���MJ���<�.�;#{�b�Ui�U�W��.ŇV"���ΨM~��6ͬ�(-LD[E�؄5��I�$��_����s���vq,��?��M�߬Ш���vK̕E���,����O=tBd��±��mt��!�z�H싇U����5��^_f^���B�z(�3�lm˰R/g���Q��Bb��EhR�����(ا���M'Y��y��4G��D&�v���_�D6ۖI蘴��@���ߎ��ϒ�r��r�~��鹓z��&52�i-��#;h�odÊ���ZC��|�NX_��d_s=������/�y��U���M���A̶ȥӎ�+¹���B�7�l�&�9�u��a3�r��ZQ���z�%�C��S4�{�O��	A��E4�;��~���s̿���~r��.���d?�=(�Iq�V�p���B��牣�Eǝ�.��+J����+���_N�YĆ&���D1��6ܑ���W�:
=~��M����]͵y��kD�N/�8��S�Q/��"^"
H�<yPh����<t�q������f����'c�dQOҘu�z~�c�#���4�,��A�;�@�V��g��o㇪�bO��U
�5�����j2�oP��l��O�L����m �c�-C44	��;��TߨS��S���>�]a���ג�Bǫ��3�r�^CR]S��x��#f��jbU�ȷ>�[�l[9��z�Fh���_�I��/X͟��
���P׵/-ك�i��~�uZ�$2�3:�ƾz�<�����Я!0����]��3vm����!5�5�m����-��.�Z�K$��Q�o\?`���$�y�,/�Q��D_�'��=8e�{VqȈ�@�s�2�O�`� �(�L��uc=x�g�M�T9��!��'�eNUu���U��ZE=�A�Y������r^2�dW��N�Wϐ��Ey.�V���@�����Te����xz��3��;t�$L�m��"�'b~��A���rs]�ͽK�V[T���%{��okX�Usz|�Iz��%���c�ّ�w�a���T/�U_ʥX���!�{��ۛ����.Nq�%2��?��V�t��2?s�� �^���Fpԭ]s���W���Lm�ůi�R������� ��X�"�	�N�7$p�����!2�F"S��%A:��Tt�c.��X�b����v ������6��7�5�x.L%HqC��5O��ۃM�H�wJ��x	�����M�1W���L������y�/����Nd@�ƟC��S �y�%�{��3Ig��N�gL]��6�R0�j�b]`�ǌ�|����ʂ@�` ���b��"x2��.��ٍ�Ϫ��*�|��ޖ{�B|\/	�U�\������PX׵X��:hNֵ@C���C�����zmc;�D�v�bN'�EԼ����U�Ru��%Qa^���f�J��kml��\0n���в���f�֎[�D�����p�9nɁ��/UV�N8�q�Z����%G0]"5�E�s��v� �њg��B�~^0`3h�-~���aٕ�]s��H$2�{����E�˹y{�Rx�C޸R��/S{8̀d3?�y��?�a7���'�,�Ne���/6�����exf����W��y<Uv���x�|6��{��BG1��Ó�vH�MUn�F˰q��[OjJ�pR�e鳑�0'�&�ً���s�^eYۘP� o6�{�J7ôԵʺt�x)�1��sA{ќ��o�:i�y�����m�����b0F30`�`��䛝"T���zfMO���|�9�*>�b��O����Q���
����Ԏ�n�ԙ�w�y^>z�0Y��B{��lk��������3��I�����9�v��,������ݖz9��K��:@<ł�1~�6(vB/@���&|�q�髦.u垵��{��yqrӎ���aa3 �:�*3&��j���[j0:aT3uv��"
w�+�{=ʇ����_�j��<�FQ�g�-�Mp�9�b�d�.���A�	�F�'���[y�[K⯇坺�uc���~��0�\([0��E��'v��pH���CM�j�Bt'��z�v*�e�K�����l�ǵ�<�3��V���}jgO���P���D>Ä�ƀ��kK�	�8��0��͢����3���E�.�c@$�0��p�.����k�ٮ���-v<�=f�N�/���{FiΉŁ�y�r�j"��Ӧ᪥Y�z̫�oP�1��;��f��.�!<�/�W���� �40��s�R�w��qYJz�ŧ�1NX���a��'��m\�Qf��dU�n�y�B4�%g�Ci�'�>�p�F�ɼǛ܋��O�p#*	�0��U��k��qt·k;T)�''C�vY�{	q�Uo�Ω�]¥�#Yj�w�i=��#3IJ��3X�C	�٬q[3;�9�\ԣ�)���|?��}@
b #B""f��'�,���3�s�a�`���!֑��a�Y�(]�*�=R'X͕C��K�E�5霓2�:�8�BȽ8x�����B9�a����ÞN�F��]�:{�k:k�?+���ē���E��Z�ڐ�9�;!�X�߼<�~V:�H����u��=��ʰ�Ϥ���&gxpź���v��>3�P�ʁG��J:�"wml/�l��U�8���?`��42x��W���V9VHs�cCua��4��p�,ߣ�C�fz�ݐ��X���~����o��O���+gy}�������_���n[4%�൓����3� C@���زO��oF�k�y}Bhoh��ܬ��#&<����Ʃ	�ϭ�Y���ޯf��KL�eP�����Zu~��Iz��璖k97>2�ԯ8��o˰��z�C	e�v�׳f��c�:��;�����"���ʖl	���$u;�<+�Uo���v�8f�%�y�ɪ�Jz�]8��ݽ4��Z�_��*��1�fg|p_�����]��y�R����E|w��?z�A��l�x�@�c0��̓�ww�tu��~��H6��W(;�O~<(���t:�]qկ��䭅�˙�\"_�V���E�e�F��1N��6H_[)6���m�.��Y4r��x�o��k����F�"A���;-�w�W���-F �P,�d^�Ji��4*���ơ�l��S��(T��Rvj&�j�;����0Xl�4�'�ҹ�e2O~1�G`	H�T1Mm~�zY�ϔ;^�ԷtF'S���τ ��R�o��g����y k�{m���{�+eJ.�Bb��JJu��f�k&�+�-7h����ˬ�N�Ϣ@��$p"= :[��n���;�b�oM�d�����4GJr��s�]�m\s��iТ��]4�A�֎���	���aᎾ�D�v)Ơ�2v�p/S.�bw�m��������㸂���Q�l�B��&$�"3Wјo�Њ�ݾ�}�3���'wᆖ��_�
qk�����ʢ_�-ݚ;pB>��L���[��}��7g�U�3��;:��0Xwy�k,{�=>�4'[<^h?��B�v3�M�O86�]�&C �h�d��ݹ.������4���ɺi�" v���[m�>X��m���1�ݏ�6x;�1ឃ�v���G�![�8,�n�f��do��L3s�=�N��?�|���
�w�1���fȸÇ�Uy���2���f�Y���칻,���m٧ɋ�K~тVӘ����[K������b���)^�|�)8��e�xm���;��R!�%�3��2��g�e��X��>�q�X%̫64ŝ���pV]%<�NƠ	d�6HƷ�F�94C���R>�͂�p�3)��IZru_(e� pj;[��>YX��T
�ٙEV*o[�:
���z�鎺�3i#��_:!+Y�i�16JD[�@���:'9�Ms�:�rTtf<V5�G]����o�{p��s�d\&G���۹��7�I��hn
�J���� P�����F�Laj��$�'Z�6hm�� �f��{e�?��Uf��v��.�^M�`t���O�"��A��M����4�e]c���j�L}\&�wq^�P	�Vs��=�˴��w3�9Jh~v�T���ER�`�	�������Bl$]δ{C��Ҕ�UԖHξ|�l}z��R��g�a�ݵ����ö���@z��=��8�1rD��@�L=\��d�yg����c{[�
h���{�c��8����ڮ����Wo�М*�b�!2p�+.3���ˎU�'=�]xe�F�'�R#u��|������t��ӗh���^���w=�����UWACn�k1Q�Ov�M�Γ�Ǚ���*�Ι:�6_�t�y+��*#> ��e�&�_
���.�8�hP̏c�此��Z޲����.ם�@��k���=�X�0��9�-�Yˉ� �?��|.��k� y�LA{v2^� 駜Ӧ���@��	V+�!���6���,ͳj���P�-#t��+��v�ゑY5��X��q^k��Z]^�L�GrDd!:��XpWZ����̭�]3,��>T�]H^W�Zݗ�B�
��4AV1��/u����]֑2�_L�[���Z�lܗa	T_l��3\Uy�����c���o�s�<��k�.�2�8H$��Q�l�vF1Z�孭���TZa
�w�ṰՁ��8�а�:���;X1;V�T�����w��-#`�y�^�urR���kVA��Nֵ���n��]ͥ��&�"�u=z�r������/)��8_;��Ȭ��2��S6
M��٫�(�y`CtNL�U'oγ��lu"nZ�a�7�U�Y���Aa3�tN�=JyH����{�n���&N+���N�,�:ыI�O3��z�Ϊ��Ym���Jah�qR����ɋ�]{�]c=�w���fF�]�s�v�|����������E̍��Ev��˲^�]yxj�#���sF�N;�z�I�S����9oo��v�Y�,�#X�뒷�ܥe��w�vonZlY�nIٛ���=���ܗC� �$r�	]�WੇQ�qQFQB ,���I���q�¹�T�8ٙqC-"���z�`W��k)k�*L�1/,��q�&3�m�E1+"S�xt���{�bc-�-��֬XJ���b$�+$���
�/�q-�H����	��ON��=ALT*K|������kS��(�J�T��8�ڙs,-l*E��2	�����Ί
�R��JY֠Va����y�b*�^,V"-�H�T��L:xt��J�*�{B�r�7�ǘ�E�°��P�jJ0L4�N�ڥg;B�-�$�"e�q5�C��	�"��T�XO�L8i駧@�m,�«QKh�P�e\Ce��˹��\���̵d������X�N��:u�.B�@�R*�jV�j	S��r�D%Kl�1�L`�t��ӝ��c10kPBb*9[��B�T
���+1�,�
����KZUm�G�s,��Z¥Z���m��s�������(q9h�����*�b�����L���t�� �7�f,�Y�:��v���8��k�Vr݃:L�+
sϩ��gs���r���Uy��(��y�vP��7c0�6�gJ�S�������ѻ��_Q=������-�N�>g������,�F ������߾���߷�wL�4?�_~U����D�� �-��$�!�9��>����;�M���Q��5�P�L\��D�+�e�81=�_ӑcα:�	������*?yIO�G�\Jmꋋ[j��D��z�,���+�8�J�!��6b�j�W@�t��zw�Xt���)�;�Kc�B�]v�֯��zg$wZ�ڼl�(�����{P%�%Ր+�;d<Û��4�ic����^u�B�x�Z���x~5��ʃ���>	0�R�B�����5 v� [�}Я*3'X^�+��!d:��4G7�\)��7=#��_Jnj�Ƚ��NoV���!s�m�nI��Xb�}4���=^�?������}�.�@���*�)�����+29�M���|�(c�.yAE��A��{���/�!�*a'�c�d	e9Zr^�&����Λ֩12��Bx����P����8�>�(6���@�u0�����ǐ#���<,���21X���;���K�/^�
7�E�
�Y���C٘\�
�ƀԂ�aR��#�����L_c|9ϊ����)��t�uJ�IOkf6�_�~Ivvd�G���$�M%R~�e���z.{{��[����X_5gF���t�_4ft�Wb��KԖ�O�+�S�}˘�Z|��L��:�\�ɐ$��f\���q������+�0b"1�9�>�o������.�X��h�?��P5�O���%QaV�y��*��kO=8}��:�i��#`�	�����t�bP��hg*�͖�N8�=+]'%鈕�UPs6�.�TI�W\�v%�l-d5��B���^מЏ3:�7'vf5�u�P�J��m�uAe���vf��V�:�y�/�$k.���^�9������0��~~�?|��d�:��&���F��w[2����l9L�AtRz�ۏ^&dI�"�Ư�c9~���Fy�Sϡ��-U�#_+�W���u�o����Q!��3`� ���1�{���`v`��3����z�kn+8�aM,ή�=:�j����ƛȎ��������4���Mfb���b�7ېa�M��\ݱG:�����n��.{�!Y���S��N1�����[\7:���G'��?�����[�L\:��g� [XN[�#��F2W�R�Gq�ԛ�܄�v�q\�[gMdK���ٴ2�P�u<r�wFc����-B����a�!��;ګ�4��O���'L���,M���C��a�{���)ܠ�#�::ŲsX����_q������g1h>��ZZ���?�N�ẌW)��p&`�V�i�G	�wx��su�[�oV�mU�J�ۈGP�C.�AK���w<���'P趌�ߟ��E.êu�4N`���v����\�R�-bQT2�g1�����n�8�L�z逓�Rn�ދ������C��#�T�PtBx׉�)���Q{�Ź��&�ŗ2c���ߕ���ɝR�y��ӳǵ�#M�aR�K��q������y�tQt��T��<S*oS��/	�2�	_uBSj���79�-V*�B9�8M���)Y�P���*L=x��eH��t{m�\��Y��v�� ��6n�e�P��2��L?���M�G�e�Ñj5�1��i��k1(˞!��u�0zy���8zB5�KHn�Hp�_�LKj�u��V�+ֶ}RD�9��s"��O$p�q�K�J	{��PD�vB�`�CØc��*h��Ɖ�_}�wd�dc�s�k{||�V܀�47������骷Ϗ�2x�S���J��<^駳[�S����k>Z�o2�n}@v�v�ғ���ӽa�n_����҃��H���V���-�Ox�s߻�|Ȱf�����X~�n�;3�gy���x�;O����t�:�M<�s�����Nr��~��u�[~�WD8j�*u�����؋N}*h���5~}���?�$ACfCLb7��o���O�.�GQF290�v���Qz2*E��o����9��fX���ݬ.^�����U�w=�l;Xo�����Qf�������w��V
�T��ꋅ�#����Yp��n�@���;�X�A�t�����b*����i�F�����/��T��U�3�@����T�a\�����S7d�[��<"a#X,�s������Խ�u�1�p+�_.���t����&�C��~T��d)����vA(����+gN����H�lD��=�Q)�.�a@�f=���|��3��,D��
�K��MM�ke�}��p������'��"���oү�Λ���p?q��6�%�$yܧ~M���Y�D@d<S�ϷB}+��D&I��Nm)�#)��n\o;K1=�/���\xE�C�?��`�a��T�L9��˰3{%�wJ�I����)*��Ox��Lcf�o	a4a��њ������
!��Bm����;z�Is�!��&P��g�z�B�'��f��z�X���Bi���6��i��@~�lO�b�r��˟Q�c��ۉN,'�S�����	CvW<Y��C�*;��|w<g��(�1����ǽOX��o�/#��X?,z�C�uM���N�8'���쭖	�*d��Wk�A(N*{ͽ���X~����cN���������)�|[<{���{ /��u�[N*�͉!��U����>��t�QɼOK7�Xԩi���u�}�IeiXr�{���
���=�(�ƣ�n�ׂ�߬eO�=�]�INk������L�l׷vl�!�B��ݿ��gn�w~z�"b�L鼽�E �K��g�k��ç�Q,kX�HX���E�e4۵�a|ip�C�� h��
�Xe1=|�e�G��N���0���y��Xصw75^lu�;�Eҭ�����Q�C�(���s2[�_}��4(q�/o/PG;�}�)�Ev�����{�8��,K'�E}�4�|g�6���*+����X%C�G��1�g��z�����V��tf~��*���(`��va�ѓP5�c�{�{$月��W��vrO��A�U�+�VI�
�H���X>w7��c��yy�sp��ɅZP�[A�,�vdQR�Z]�#��<>e������_�����pk��/h���hv�V�xL�.��B���}$ƭ�x�b�B�e3L;�Q}�ޠ��y�o`@�j��lJ�#իu�G�B,����kk�Y޽�ǻ8;�stL�	w�qտN��$�1�Fəb��[L��ճ��I���6�=�%��۰imup7�:����΁������M��aMeN��kQ�F3�6��K��#�����^D��1����u�>��#��uu��lX��~�����ol��2��JݕOv�;��>�ȑo�A!� ����_�x��XǮ������vι+�<�K����Z��@���2#�Uo�X��P������(+��{l�V3�o���K���a��"��)�F%�uSL�{�Me��͞�!�ʚ�(���@�UVW<��%^+�
�L�n��Ɋ�/c����ʹ,Ia�k�]���T;W*��b�w~m9�Yj�)DS>;<�l���H��D�0��#�^��Mϴ�� ��G�T���p+�5o[Cĳ��	_�M������7��T;4��r�gy#u�&��ʵ�v:Z�z:[i����铀�c pn������@H���,�<�^&�����FoII��G˻t�Z���p�2?�Yۼ�Z��̊[�$Om�w��Q+tm]>���B'�w���Qt�?~��=�I�S�|�(~����2���`�e�~���7�`ѵu/��a��q�"��*�oi'����J�ά�q�K�7s������:>���ރ�t֮� %��6+�؛�x��[�"�!��WT��?����Ǖ�@�Ƅ�9$ ����f
�i�|qN�DP�^�A��աm����������^1ɦ��m�kz�x��g4�;��>���ှ�5�'��˳#]�P2�Լ��X�wY�9W�
驨7��!R�so�#e���PF���ڵ+��+Q[v�I���b�g��MJ�Y�=B\����7V΁�Y:1���vC�;o^��[[{��S��!�7����X*�˩�gL&��u��k̲�
�=	ͭ��]������S����1�V�h&D�Vy�x\��p{����֙��m�]��,_[��OL`N�FF��O�Ϟ�I�����~c�Zd��O����*5l�s�׎'�EkϷ��&�ѩt�����n*���1��(����GH��*3��f���qH(��O��DK�g����awp�H�] ��Cz�oC��1�a.�ɻ�F�\[>�p���M(D/*ht�
f�u\R��*��j&p��I���8w(��W]�K���i<68���&�X8 �<չݱ��V����W�v珓�������Mܛc8,y�5ci��ƃ,��s���ol���^t��q���Qo� e��Β�7�<����:�my"jjS�`�/#)>����8ӌFES��&|w��j�UA���F�n���l�t;����7�����6�ik�ǖ76�#�Xݤ<�/:f\e����\��[��1��Z��/���~����X�
����%>�40�����+���:�S��b�����l�i�������V�?F<�ry�;dUт7�����ۣ�YV�4^<_<VV�D�*,���������-��pʾ�+.6�o��S�H��6�q��6���Q��Հ���Lp��p� �lT�v������S�x�8�SJ���	��edәY�X�mu]�:oons᱊_�#�d\-�@��(�0T.��W����.�����1	t,��uO������F���*J\d�VT<�oT��Ɲ�"7w2&}D�d�Ƚ��.U��{yr�&P��Tӎ�)���Nc�9A�U��c��Z�e�DV�Mx�}[���ۋ#{ksKxdU�nŋ5�������r�y:%ϵ5Mw�ުk���T��᱓�hd�4,� �g�c��(䨒L�0���Űo�~Vw�ApP'��1$�%|��g�q��vϜ�Ei�'����>�)R8�S�<{m�\�Bڎۃ;i�ǁ�Z��ט�5�uoc�m#���\���`,���B�w7z��-��oLB�.0�9�2k�x7�Z/ l��D�c���PwH��g�k��l0]4��U�C�{�ⶺ�ct��+�A��'�]oԷz*J�S�,+<�N�X������cji�$k%ᢔ8G�G\�
տq4۰������X�iU�yU�#v9tֆ���pa����X��m{8цB��&U"0`�3��$����>���������
��}��	�:�`��n���/*�V�y�{�m���ҫ=�B�e������b�����#���dؾgK��H��B���2�%�*��ǜK7�H�`xO�	��dtr�\��X/QC��3gOo���/����7lv��ۂ�e�����Ҹ��>W�~�}�6`�R�2�X�k�D�u�z���צ1W�4Z�(�����Sm�íj��e�WK�w�Zx�f"/����b=�]�c���H1y ��m+�T�q��z+�� k8�7.m�W��"L�nY�	�#y�p��\+!X�n��k����O\��t�vF����J�3k�oQ^Ȼ�(�W�Ɠ���w�9���k�;�Mr�<�٧g52�p��d;��GrW!^q�fD�n�1����Z����F�a��=\2�����oV��l(70��m��ձ@>�H�J꡶噀|k��Z��h�i�9��3iP����ȷ���!Oc��k5L^��1���y��;��t���*R�2v�U9�f FTB]pM8��Þ+���(i�^�ٯ��R�Ҹ�"��;#Ha�q�s�t��l��ռ ))��@�{����Jz�/"��lO~�݇�'n5���zc�ۺ���m!���]��9�H��9�=�^�\��q�X5��u&��\T��Be57�s�Y,�'8!�Xw����7��nt�� P�z����*D����{�à��i̪w�}z�w��c{��M��:��s�K�M�c�t�:�b��s����.Ƨ��+�ݢ���l�,1e����ܪh!���n#+�W795K2�%�w���hSWE윰���35�/�IL��<
,k$`X�l�A��)):�^�δ������*�Q�8F;{Wejt�ݒ��� M=�p9�wPP��A�y��*s�Fv*m�쁠�r��:���˾�|Z��\��h �+Bl{�<�m��إ�Erw�o�s�b&�J�]�dk���Gx�����@l\l���X4q��k[�%�(��8���iŎط��򎂷��*z�l(�L����	{��Q}y͕*��.]:,vx;�oXj�&E�u��rV-�H��x�G�?�.�\��	����̈́6<�Y4�̢�k2V�nEŃ�vlu��n��_��K�춮_���VH��\zo-��Lɼ��q�$��Īaw��ثq
XJ,�w8�^9��HYwg9\�#;�7V_Qe�YU�+4�G7s����:L�ulUl#wn��z��IT���g�/�T�/	��7�n�Y��Ϫ�i�T�A-܃�=5Y��{UKLEMVh����.�plv���x�h��;{��>K��Kg�Y�jT�P���'[��q��ev��9`������l�N%�nL�sc�x�d��Z�HYo8�f;j�9�쫪���.��1���� 5���Y�ۡ#��� �bS ��Y]Z�1����6��{���I�=�X&$�M��X#�����T���e4�NQ�.�:�1)4���N)n[��lZ��v�Ω{%�'T�,t������vﺘ�/�<TO����LV����ZH�VmƲ�0w�l��"%nF�N!��N)>t]l��NqEu]Lfb�Nb���WMA���J{t�0./;�3t�vn��f�sJ�n����J`��=���cݩ��2�\��5��l��˪fRX�H�#�}�����A�V��7cE����L�[�_\�fAG&Z<�����W��
lsoo>�ܳ�ԧ����>�QF��d����Q��ׇ��Yْo=3�ԙlr׺��we��QT�A�@���n`���7�T2�aġ�����R�¸��"[*@�iű�J�;����Z�{� U���̜�/���{$Q��t&�	�Ҁ�s���a�/QHt9�4ʐ��$Ö���2��̹�6Uj��A��a#���c:��oJǕ�
a�����V٪u��vy��S�R�n���2�\�I�;#Jtfs��@���V`�������N��0.�#�**�*;2�W�=��U^gR�eˆU�Y����R��Z�F��o�����̓����sw%�˧Av�4kt�X��2�A4M @�Q6��c���lb��T\`e�Aq%��%gR��[�0��çC��4E���ri
�Քb��KmJт�ܹ)P�F�LqX)RUaZ���=:w�A�Ҧ2c�Zߦd2ѭ��ѭ-�
�K�3+o�Tʔ�,1�RҶ�S��t�k���.o9�ҵ,m���
�e���˔*w
-W2�\(QQ<�ĩYRг{a�,̫�L8|>��jAb �Q��Z%T�(�*+ZZ�QE���^&e+A--lX�H#\f+\CRTD�:t����z!��J�j�pkY*�Q̫1r�ek����
�����Xq�V�O#d0�������֙����Z�V�¥��1�S��>ZF{x��PʪQe�+-���a�ON�H�r�9U���,B/K`���E�mQ�Tj���5�Y�39%.U,J�+Q`�[b%8xzzvv�6����Em-�SY�ŎV�-�Ej�,+P�)�h�+%Vbf6��iE�c�)����d��.	��P��DUK�1�(�R�̋
$L�����ߣ�o��}a��[۲�eUk[X/S��ٻ.bh�%�ozbJn�ȯ������k&蘤�N&�Wpo��D�����I��hU��Q������0<jXS��o@q�*���i�ݵ��Kl�r��n���tfE;��olv�4l1�G�`<e�>W&}u+k���-���z�-B�j���2g�]��z�`�Zq̃�AzXte�;���dG^��D�Ť"���F���3PD9$h����Z��j*U���s���4���Ty딁Sٗ�����C�r�/�1Mt[{̬�릵�����U�<�+��w*�Lt���QYgHAv6w�ɨ�殷����B�\�{o���SsN�l��OA~�����VZ�=��Y<V9�m���pu��+֌��.�n�P������m����C���׭E]��G��1��A-8�T-�:n�m2�4���`y��OعU>�B�l����H��I!.�-��$���k�W���=o�F'�B�f�S���q��R:}w��<kX��������A{�0֕�kk�5#�b���ld���Nđ^�99 ō�Ng\J�zFV=�y��.���i��4��������̮�gd�hv��u3�`7ŭw�5�'C��¬�,������]�F)-˻�!Iƨ�-�QB�ʑ\ޅ�7rD�"����p�����e�\5>�!�[>�+�ݦU��Eo�}�GS�]������[�ݨ6Ǚ�0��^��ʦ�i�"��?ˆ���}jI�~Z�}�����~=7J�5C�UX}��viy�'vM��`���Pm�k�q��S���nY�o>6����l�e��Ը������"foҲ^�)>���;��<�z�j�^���L��i��)(zyO�*���E���ا���L��(�\���L�_��>A�����1����~8�|��{tɺ����1��K����=��9f���N�`�O��AX;�<+5iF`Ƚ����"@$͵o4f2�ъ{��du|=M�M�k�7؂"<�����*��z7'�uёML��zk�=�Ep˵kVA�x�{+�v)̌�{B���#Z�\�5/��7,���p��΁�A����ܚ�M�su;���'gI�������(���@voL�Zf�Iʊ���k+N�9��Wr�N_F���C��W�6�7�A	F��N��A˗ҡ�(3�������ډ^8�'I��7d͓��6Κ�^|$�W_I�c<owP3vE�VO	���V�F�>�ߔ�qN�t�РZ,#�����fU�UQ]��o*�Z9�B�2t��� ��&�CZ��\K�1M�'��n�˥���`�D�W1�4�˅��k�X.2�F���{3Yo3�vӖb�_o���o�x̪���2�t�t�x=D�0/�!��Zl�z�Y̺x���� FdUӝV��P ;�.D`a�}{��R-+2��|.i��WY���76u��ں�=��0���C��8����k�n����5����V���K���\�>�Yϒ;J~��-��ns��.�Ɓ�����|�}��%�g�W<�)Ex��]c"K��M���u�h��(T�gN!�4qxv�C�<Z�n��-ފ��*��MLN?t��ʹם�<x1�iSyfV�=A����NwXv¼v�I#�|�ʲ�u���gb�����%��,�][�������$:Hs�#Ҳ	�r�e�y�{ÿb�<��0ZѱÎ���pb�?�_E���zWlY�aΜi��.4j;.�hm]����:���eq�3�_Nx�+	��gu�V�"i�{��5`�z^f��p��l2�PK}dhd(�zĨ@9�9"�*e��Vٶ�%�5T�f/�5�-�V���̱���h2�hw9�pΫ�G(Ktm�d!�;���k:n������A�x���G��; _�_8�C�Ӧb^�.��5��M�\GI��Cx�$�.׏9k������o�!--B^&k83{y�JNh�L��ˍ�GP� �*�Ux?�\'6T�\Z1���0S47��^-�TF;��=T�f��2*F��;3�*U%��ɢ�6��K��'!��~|2%�E�O�jÜ��X����jx~S߼�rVﴉ��U[=�MNg@��:hvj�}�Oi����Iw^C��,k�惤��sg���\��l�C��I�U���P��)�]��1�!�@�B���-�R�]�������Љq%����W4-�K����CS
c�a0���~�ۉ°@͓���A���X&�3/�iܻW�e�0����C +��{��)�q��������>�CO#��/���aʁosc�Vf���/��Gl��W����R�t�tl�툫�H�6��u9`+7s`W-'��;�_h�����|��g�v�`��-0ӛ��:NT��렣�!oC.@-/�c��Z���1f�{����\E�Q�2!tu��ؕ�^h�U⻤<�����uMI�,���cg`z^aò������g�pw.���q�W3�ۖL�*g̵�0��!�݌ަ�\���nT��K����Ր��&�e��o��ޥ����n�7�ᣰ<w�|�P��2�^�i~xΘ������u�o��K��z&F��i�^6Ǹ`q���
����s�>����`[ʂ v݋�%2g�u�1�'�i�29�:z���O�1�����B*ѡ��vnp�s��xǘ��=ı�hQ�T��?ukF�^\?!�]Y�p��)�3$H�<"{,@%�V\6_5Dr����Q������w�`w����:<BMw�Y��%YS�:t@�|نߞe�.l�����wr�l��;]D�yll�D�h�u�#�]'\r�s7�����6�ۉm>�mc٦L�V�C����y�}�`Q����u�e�d��%"�1I�_	�quJ���o
�F�*G���%��N��٩	�n�.;r��k1 x�K=ň��)���my+.i��e�
�Aâ��:B�G��d�jBj$j�;p� �#2��J���\�v�ji̊�vY,��le��y�t6�_d�sϝ���V�^��΂�acM#B��K�钪�n�/�xLk�ՓaUo�$%�:���:���;Ғ�1�V�ܗ����w��������y�T�%��g���W�n�%~�H��zʜ0tMY�`8?n>q�"&��	;����m����ښ{[�)v�鶴t/�����v;8����r%��*.��J���F`��w��(?�r�3��h�Z�-C���.��ʫ���4s�x�mQ�i��g�a��8;�Sk�p���n�k�V����Y3���o%��55�(��xe'��0w[oS�ujKݨ���=�H���l.z8x�X"/2�TH�ǣǤA��w*1�K�Q�����J�,c�U\��_�1�cs�����NMF<�衊��K�4���x�s�$�K82vP\�+��z�G��p	����k1]v�3
{)XJ�b����J�Z��p�O���K�;
�&H�Agd��
S��O����9z7w+Cf� w<�u�x*ke�*T��W�:`-L�C�Ζ}������1�}�[��I�K�׷m��8&�f��ώϣT`�
��[�a�}��O9��*�!Zw�(���3ϡ������+����6h~��E�g���埤�w����MN�㸰	0�A����Z���YŎ�� �h�l���	Ͱw�g)���qx��yH��7�i(�Nm)�e�g�owR�v:�o&
�x��mS"��\>o ��B
��2OZ]wQ._d�MWi���웤o����(��B5[�*�]̆��(�Ip��H�;UY���-�2��S�;���đ���l�?��.�{�P?E_��l���s^�;�ۼ����	�-M�m�N�l�^�:Trx)�Z^}|Z4������e?T�n���ǵ�>���t]����;�ُnA��n(p� A���EŚ�]���
�����8=wy�-ް����R�&�ų�����fu'��	��u=]н8�O2��7Y�`f�K/�S���nu3�p�k ��쨐=a]L�2�d������P�d�[%M�������Ǳ�p���5�<�� g7w^�q�{����x�r*(Zh�@9��咧�_��.���D�TT�T�ͫ���LA�=&�d�\����}I)�,���DO��>�\�ju���M<L���b�}�����k�o�[�\`�X��ތ��I�Դ�>ϩS����c���a�`@�7��P0o0(��ѕ���SYD�U3ohmlm,�3۶5^.ި����@Ͱ��� m7��@{�jȭ97�s�57T]�fx�����->޴���AQ�h纃�`���4w�ƄQ�A)P��nKRqO�U����Ï��wF�Ƃy�&U�2"�
#� mU��<3B��qk%b���WMmaI����ܹ��/ނ��o� zq�pc"�mV�@��΢�)C��=ު���̵���vd�"@+�VJ�D�dY�k����Z��`p�ou=g�ȩ��a�A�*S3k3�*��c�H�Y̬�.X��"��DW�>3��;��k��aPK�{U��8�am�`)�{96&v���ʯ�CY�@g%�E�襅O+GT���רt۳V���9R�I�����]��h܎���VDg�
c��<Er<�LK�h|����,��|��TV(���q�~���!d`��XM�&���Kq����T�F�_�MEI�����Gj��4��4΁��N ۤ3o�%��1)���񷋴�i�i���zRJ��4�JnC��|oH�	!x��zo�>����f#�CL�p�Yѻ��H��%� ��>���H��e�E^��ށ�=�Hz9"1���az�,x�.65�[���Ȏ����X�r�S��y~���^d2=b3%�.�B��3݉M�=$������b+�C|�щ���߫�ݏ�B�l�������$�=�]˓ti�<m������YO��v^p�{��F����`_˜Gb�nRc��<;&W�/���K�e�ځ;`$Ml.��6z��}���sN�\j��;]m�.-QA��w�T�qF�tۊ�<�o{;L�6tEx�۝��l���R�%3��d�R[�!J���F��s#�u���X2�:J����j�=�Q���L���^�d���t�����Ko�Ay��ؽ�L�{��ƍ[̛P�N*m���#��ۛ��C�
�=�$�ŃD�P�FL��n(��{Ѽ:�6;Hq%<N�V�c�b�u1�͵��ðWH�ng�R"TȘS�s&�_�Ѧ�it"Th�x�����{���y Qb8��z������3[�}������q�D,��S蚞����S��9b������o#���{��Oa��;�I���c���Y�-(�����������ˡ#�R�V�w�)H������PFc��~a5��Ѿ��s�9���()*�������7�|@���c�;zZ���nf��ɧ�ms�B
%�0�W:�.�i�t	)P��m��2Jdol�*�nh����"��HfF:؈��;҈MlzS���IZ��3]��x1@Hx�Xو��ݐ�O�k���Du�!E��ůvzR~T��l����*'$�����}$g����d�*@A�pY F��Βq>~@�����Ɂ\��J�}L�̹�,gAf�WE��^�J�qc���O�N��=��]!k�1���o'mY2f��}��V��]v��3+��9_������v�*G�7�<��۸��"�	���P�P��]������[�g��W#Ρ�G#׻�Xٛ�;d�49�u:L�32.c�R�-r�36��Õ�fX�;�VY58G*��J�.���E

)x���5�|q�a��ޭ<p�3����js��
�Ȩz�W��)�DVvQ�����B��
 ��䬌��m:�F4���ǥ]�M����^�}�q�e�%Sv��Y���P�gy�j�$�1���&����}�=h)��ޢU����믵d�W`0k-XxW\�)b��no�Ry�.�vt���D)N�s4X;SUF��#�)�6�1��a)ӈӂ=�8{Vl$$Ђ�vk4g<sv�9�vq�8>�9ތ��g�9��c΋��-+d�f��z���Z�̸���b�I˪Y�2;�X�!=��s���)e$;�)�(u�Ga����:AAi�,C�3!ݚ�C�7+����	�	G��MY�vPlq��Ȳ�]���o�7kk�����y��ƒ��W�����%�p{ؤ&M�{6���m����[���;�O)��	�������oR���<�mL�5�%�Cn�R1�C�t�K���sd�Q:��ϗb�֪7f��f|z����o�`��y!�^P��+ٙ���%�0���v�#6 ��(WK�m�A��O4��.�=D��)Or����nf�[�S���ҵ����Z�5,XDi+�-�;S�uw������;�=��m��N9��AnI76��x�`6i�kK&4���͵o6�r�nM9�d���q�ىD��1ꋹ^˜OE�d��58-oL;�,������}� �d����&|%֫�`		���+3�R���!s$����)��Z��=�jR��C�q藍6t�9vJ�*#��ۑ�|s�l�I��N���l桸���;�e�Ql�kE��2�d{!<�V=<o{�p����7�Q�O1<�����������2��(]K�1�H9Kp��X��ؙ�������೙�:��r�6���Q+3ۉ+�jJ��΅j�����v|�Upf�r����LZ�0u�L�AM��m>���ͬ9�	]�W�@�fkAIc��gk�׷©1���p��!Xr.���f��2ID��X�q��+��$�Du�9��#�^�]���,;]fC5cL��{��N>��kT�L3�c�ekT�omG)-1ZJ̝ۧ1�J39<�bˏ���M�^P塂�'P�1�fu%C���6v�<�;NR�*�ޜ�o�j.�c���ȹ�k�!]rA��m��,���;t��sc{�}�hWW���fJs����v�c�y�6�rm޽-S�ծt��W��?����p\><���GʞF��a����<����]CS���f"eFE*����C�Y�_le���s.x�N5�U�#�70�����^�"�)�*)m��U�խAUnf"���8�N.7VcYo0�R����qJa���ӯ���2ذ��Z`��bZ�
Ue�c
e�m��%�����L:t�ӝ���aG����*�e�+-������(g%�,�Q�H�V#�̼��L�����,m0ᦝ��§Yz�����Yƣ��Z�lmK�d1�8�)���-��kTJ�lYD���
֥A0�ӧgb�ƈ�|�m���k��-ZV�Z��\����R_�g,�QT���DÇ��ӝzW6UW�b���k,a�*�3�-+U����J2�����QƸ!mF�Z1יN%e0�����ةZ���\X("єE�kJ�"�b�k*�0�h2�Y
���çN�8yz[)�0p�\m(Z�Q���I���嫗
�%�j72� �9�NxRqbB�s	�mKV����E��l�Um[K���_.U�#ܝE��d`�ĳR�X{y4gA�X����*pڰ���Kƫ�
!5m�$tE����wm�t��avܗܳ3Nɉʲvd�{[�{I�wt�Sȭe0+4���p��3h��4�S��;@���.M[����c?/���+�&"d��@Fb$���a�;��K�~�����	�*fX�����8��T���tq�J����8�goC��������Ͳ,���� ���K�ҭⶀH�R�����#����)�Ά���6�q}ܜn`j����n�t7��{�@;"�/�EfK��������1ÓXM#AP�7@R3_2��ǧ�m9��򦂝կ�Wjgwz��a+�fF�g��#�6�ЋK
���!�`���� W�&Q[chc�v�v
Z��~�gA��
�~IP4�UU^?�VEr�;�wd�zD��{�W��D��"^e)آ!�d���<��HIn�}��E���{���o�4��N^���3��;�גP�e-n�������T;ns�^��,��[{���F�sg��W�)�A;h�۶�)�J)��m��]�EI�Q�V|��د�]����C}w�c\���t��e%���uW�<D�
t�y���wpZ�w�=f	44�eu������rRI׸*<��0f-�Mg[{vd��u�mB�����@e�L�^�f��.�ڞ퇭}�7$=��{U��mՈV�զn��C�
OA%*������o>r輁�H3����d���_o���"�n7����"�Mgs\d,*{�ɢCd�W�r�@��S�Ϲ��i�@7����t9<uJ�\we��]�^sNI��<|u�I�xr��p�f>��B��2�b_z\b���=5�C����Z���4�Z}���F�m)����U&=-�G:�4[eX;�G4T���ɞ�Q��Z�֒�+�Wc�dD������9���α�.DChw�����z���%LGS��:�y.��b���=��g���z˵�1xH/Vv�?�Cq��!�E�m��Rw�=Luf����j��xfw	�v�t�Ckk�Ч���h!ά�@Y��~�}}O��Ft��笾�>��TH~�_�~B����̭t}
��nE�<��g�uA���(���7%5�@;���+^}l�D�sξ
�R�����/xH�|��X%F4��
�6nzk���Qt����l͜�m<6�V��T*�-�ّ�n^��w.�&&f��j���ٷ�6�Qkp������_�h<n"�0�h�nA@�}#Lwu���>��<,ɦ��wdY�<��Ԛݷ.��"]�����lÚ��O�KNz	H���Z�h�,�"��M��+��`>ё H��}�h����娃Gt���\fS�������367���z�ر�a� �y��W��F��ԖP�@��xmd�\�ea�"�E^���u���P�K?�W X�ߢգ^�]̓Y��j�Ț�9�u�8u�f�I��=��4�4��1�2�r#��=�ʋ�ז㮗>�[G�8��#�o��	%!���ju�\*�ȑcZʾx���ԥ����2���m�-{���Z�vG�"�<��l���NpQ���eۨmeS�j�4�s�"��R{��t�G�q��BT#Kƴҝ��sZ�'����g�)�i`]�	�GY��I
8��O�����mД��.h��(��AXت�8ɻ;f���H�H���~�o�f	%��mߙT��&B�r�/m��h�����;�P��I�ť�G� �id����9�/K�Z2�>���v��:�m�
v֍�!�L�ly��fS��\�;a�ȹ���~�������n@ю��P������yܣ�Kه�M3��D�]6N�<�f��H�.%n�7�$m�#6�k��u�#�M�#��a�����v�!"�/���v�'�Q�Hޚ�} h�r7�_�(Ȝ�XJ����3��Z3�b����3�4t�����4M9�:!�2d�д���4D�>�)�or(�����&x�\��+�bS�ɺ	ʉ����\���/>���Њ��tl^[��<$q0EV�!����U7��K3N�U�+E[C���r@B���Pa�<1 �r�o������T��]�>T�M-J�WU&��@�wrl�Y�OC��J�I���+��<�@�x���#��>�dx�j�� ʮ@����W�n�ǺZD�
.�[^�n7M]ط3��{�	�{�,�)*�eP��.���4���l4]���/=�s�+�΄���k��#�Zec,C��x��=�b��3�G�+�;�%X���ipx�X��d�-�oF!�[��X"8"�%gH>�]�˫�4��X� �ɧ��v7kXܻ�/M�Yd�:bt�>�|!�\��v�F4�(���'k���߷�}��3Y0��6X�)Jxe�Rt`�:����t�0��%*�c�S�۰��0��:/g�"i��i�+���:W��G�x���	;F���3b`��72)��m��2i�R^}ː�N�ky¨tV���@ţvy/\�~���]7;8�c#�w��T5��m�ϖ��l��j�B[�ɍ[>��;i���U��!�go���ї��v�!v��l��,n§5�v��A�����|�}"/�7:8��*֗�ot��4��g���;l�.����]qm�ä<d���v��eH~� ��E.�D�ԧ38ԣu;2��D���+�y{��av�u\�}]�h�U�yNWP-VtcK>YzV����~�0=�n#9�0홁�d�پK�2���I{�Zd=L�EVf��z�[Z��jGPm��$uG���͚}����a��U�3�~��C�z�J릘��g3�MNݭn�M 'P19m={��4]ٮ��6��꽖i��p�=t�u煨�՛�5P��?Z��WK�c�ɤλ�%�Rr0���/F�o���Rw��ƫ8mpf�d馩7'ry�03|/���ͩ��c�~f�:h�0ی8����<�{��`z/�O�1	xЧ��$��ġ�=�^��:�|\r"�:H�qW��c����/��������/��ZM9����)��<M�{�@z��D�T/�$u��%rtu�ٴ�]2m���sm.�7uƸf�",*��=�	c6M���A����'m���hc�4�{�댋�v���4/�s4h禡
��xj՗u�+|8�8q��j��Q����6o�_Mэ�n��j�4�;�'>�����?NY�ZWuX=���s��Щ'���Z+Z�I�*n�t�F�2[�����vGy����%���\����j���x���N�;|���݉��|]���]�Q��)���=z4L�
=qӶ^�OEg��s��R;���/NH�m��kFȱ�Ľ���9��]�&$���\���R�}���n�=�Q����U[���r�����%�7.o�|�����*G!����ͫx(��)�{2c�(v=8V�Cv�G�:�Cʟ}�\Qg6���teΨ2O>ᷬ���݂��bM�}"�f��Cp�[���LL�U���/�'�>��}lw#�C��Ҍ�ϙ�0�o�|�F�e��<lDb��]O�u��R��w�wi&��Fݙ��h�U�PLg��6H�o0K,F�e�T��Uc�����1�ի�F�5�9%U[ ����m��a�op]؋��JQP�m������f�4_ez�#�I�=G��P>|�:8���)/���3;�^H�j�1q���t����w��0H�z1����fr.��K3���U>�5����<��3�΋��ޠxo�� ��w�Z�g����z�&گ���ݛ�3�
^�hЊ���p��݄X<
�8Nd�C��z��k�]�M։�ނ�ߴ�=��(U=S6z�dV����{9=W#q�,�b&�ا��q�i ��D���W�":E�E����׉RК'g"s���[�	�~�j��*]W�/�H<�����v���oUɋa�����S0r��B�݋�_��+�[\�8b�n�r�X�om������#|R�Ѻ�HbqL��SA��ip�+�=(���ʹ������̖�tZ'ZX�3xM�����5E,��A�{������T�M�Z����P脍�JFV���C�XL7m��dSl�KC���z��H��
Dcm��ލ�H�:D.hZ�N�j6	��/�MuE����2Ĉ+�A��U|Z=]%Q�\o]�ɵb��#cS�<"jNl��.�@~�B�d�6�����(w�vݹ���ʛ��Nd��v6@a�,mP7�L1�n2��N]���KmU�M�j�����D��
X?��8Ꮼ�]�]���{�E���E�[
Q٦Ki��VP>ݣ�g���A��s���Y���_g2�&O�K�E���u���h0�X�k��#�~�f���9I*o�x�f���,X#�0�C>i��p�Ȼ V"hq�<[�A>��ŷN�U�뱹5��S����f�����`�F��į�â[����1����d�&h.�r�t�VķfX����39�)WX����9H����|�R�:,嚔�-�A��9���,'�Whc�K-���M��ҷ�v��ᒊ��˻�v�o>�&�� �C-U�M͒ӽ=�Ey�V-]�꒞-���͠Jh}�S��w��[W�Ie½߆�ŝ^]H�g �,�%~���������|B���w\�U�����l9�{-��{K�^�K6Mӌǐ�w%�/�B�'�c��p�w�q]��;�H�l����#Ņ+2W[O�)M�9��O_.Q]�u>a���p�w�f�EM�*�b=�!�R���k�z�!m܊�r��3�:e�0�fUn����Ѫn\�#W#
)>�>���+�*T�T=Bo�Ճu��"�[�!��&��P��%lEm/�)"Ύ��e5�66�Lݭ�"��Nq�A��C]9����b� �qk�藙�y�gܕ�N�D��H��V9�J�����?Hk����cV�Q
O2���~����

���cd����\lwP=O�	���� W�CM���O��JV��l�`���5�j����O�}��mt�L���c�ޮif���@����w�7fZ�g7}�,���APHV�[�K"pw�h�����)Z�}a���� u!�z�Nɲ��Ž��k�'n�ב;����˱W+4hL"��=�x�xy�L������O�c(��M=���oE�J)r��\��o��%�c/���1@��/�]��%�31{;�6�䖪��FC����t�'��X�8ÌF}.=�ԛܳX�W@o)��E�([Q�us�M�P�Ý"A��g��q��.�^���G�.��j������m�����U::������H�� �F�c�
���+��3�j�`3���s񼌻����HrǙ��`w�b��,P'��2������?e,�QFV�z��3Q<
�/���校�����ܙ��=��ޮH!Y��Ta�!J���������ml���EfN#7�ks����j�n=c�y��B��j�D�D-��Jm<�	��@f�˳;de_0i��v�4�b��B:�,�B�n� �@�ٕ<�34�6c2�����:��#��;w>�n���@)���*@�n{յ�l����|ڇv�?],������=��L����wt��!��;��v��+Im����^}0tP��d��}y2��^҂Ξs���8��Y�`��1ce�;�R���T묎�R�cĸf�w�Gs���sM��\�_�ּ�XB�)�X;Z��"���M�<@��X�UG��QuF5����RY-�"�H.)�T:�wb�KSuȵL��l�`�x�X�G�Զs ��B��X��r>�w��X���M�Ʋ�]j�}�i���֛�6���CV:,�t��̼�AL����e�+�>4��C��w��.�����u,����ٱ�/D�O:��8(��v�s^��/E�FU:nǅe%=6�j��N�[R'av�o^��7h1����2p���]8[ئ�c��Jΰ^�6n͜N���FH�b��P��^��6td�>�)�h��f
�Y,h{an����<7q e��õ�8޸��9�7�jw\�%5��ERBs����k��xw6�A��]a������)���R��`Ǫ���->�\)��+�|�d5Ιo{��;lXs�gj�}b�t��fQ��[�<#w�ٷ�f�tc��+�d�����!Ba�/^��H�=ʵ1��y]��j�eSy��n�چe��#Ί��9n��Uo�R<�o�T���呼��n>�FW�zާ�O`#I�ݭ%R��\0k�v�掜�X���*�G���J�ĎW[x��x�
�z��T���)�N��ș�Ʃ���k�"�믓�n`��j,�^�Ї�u|.�#��_iU�h:�ܶy�Q<�>e^��ҝۍ�Ng���a��J��\Ͷ�k�B�j���W�1�=�X��,S�>�08��R�Ace��[t�ZK �&�2cdr�Ƅ{u�m��N�N��:Б����ɂ��v�U���Rs`��o�G���:=%��t��pK���%�ʹ����z�t��p�QGn�ԓ;rpm��Tܧ�%��XEn�IԎ�M�u��1ɸ��B �\Bid����Ӝ"�&j���0c�3s���@��w��lZ7$���D��ڷ��J#��&C�ٕ�w2����lˢ0@(b,#9��L�ۮhc�3oo5�0!�Qó2�_:�fc2���G\�汮��o*"o(���{p�f��;��dڮ�Go�r���;',ƳɈ��Ǒ ��G�E��u��xHm�|��)��*�`���(���J���je�6�Y���s+ ٷ�q7t*�͢���qT���6�����ք����31̨�.��e��y��Z`Ψ���K/mY�n����e���fE;Y�����nÌ�|��vÒ{����+���� ��o���v�usN$�
��fE�Ϧ����-.nim�&:ڦ�V����Q�s��X?*�+�K��!�s,�
fU�m���/
��ڪ��)�f�+�L::t�V����Qb�(�W��%g,�0T�����9��:t��ZΫ]�^6*#�#�b��meD@��2�m(���33
%8zzvuQ��z�1�*����Ĭ�E�Z2e�H*�b�^9-��Nr�A�X(�8p�ӧ|B�/YDA�m�D�)s0�a�J��2bzʪ�8�V,�Xa��ӡ��oS2�8��n1�Y�K�%J�����Ӗ-[�d=pV,���<0�ӧN��1�Ʊb���1S-TTFާ���{��d��1\q'^"""��ç�N�{��mZיq�J�UVV��̡�� ��s�*e��RR�,U�R�0�ӧgUl�|��|h�(�Z�CrW�QI�������Z"��b.R�Zآ[X\9JR�Ŋ-AkF��b��Ԩ��X�DRե-5�j*�b�V��e,`��Z���f�����?V{%	H�KtU�9�����絙�g���*R��3�$F�jvH������W�Sm���8�i���1�ux=@�ג*���]:����n!$2j���^Z���QcOPF|/K@5Ďy6uwx�z�����-kն_[߶f��	<�u:6�O���*4�\���s�d*ƫs�$���,�S���|�C��d?R��Ƕzz�e{��J
�܄]d�ܘϙ
��/)���V�CFt0c��\dDb}3�����*�p��F*/�~��iЩ%~�����>�@P�P����z��z~{oo��׵�busq�v&v�	\7�ݎ=�^��`f�m�h��.��GXV-#��n]O��I�}ǋl$F���=A�{��G4�ɳYN��k76��ox�D��b��Θ��p}/Ǟ���x�]Ua�Z:[y�hk�{��^���ljwb��5ƽyށy}2�x�������{/�f$_e�s��̭.����[���4�
�e�x�!5���e(�$|�gymB&o����vr�����D�m�P��o�J�{�\��aء���4
�v��W�Vf�y9t/��;��/�Nc[+�r�5W����	��E�������ſO��
4K���|Ī*�.�v:�3�,�N��9�?5m�޺�W� �����T�KG�A)���љޅ����؆I��c�������Oh4Q��B�c�~��20�A\�����S�-mJ��>)����6�0r^�2 ��X[�T��&w��ם�umXcv9�){emnU=�^�
m����i�d�,�I&<e���[����vs�]A�p��a�)X��-�к��Fd%���Q|��wQ
����8{�
���<:�`�<&}2�_�WITzS�7zC5���[O�R������'E������:��bS��uΚ}ֱ2j@����]��c�v9u���<����	50��X�`��3!���D$5�������Uv!�����uG�(�k�蛥=={ t���/�tY�G���J�1��f�����_�����x��^�2{�,���9��ڔ�/:��"�%��������b�-gmy�D>,��;&�.=c3Ak���]���"te수2�]�l�:�Wd�W�A�5mj�9S�'^�W:Y��Ul:\N!'�".�d��]���']����PT�%�s��7�ue�Jh]#g�M���]'T�F�Xh3�t�		��P����9"Yt��s���\Q�mw�%;���pR��7������~�o�G軇G�48ɐI��VͶ�J�~���dMLޓq5��Z+�ح�.���8�f<��U�^݀�"�<_jAƧ�5@�u�-u"���Gc�hkΈ솴B����LJ�;��B`0�/�+Q�k�6����=��?W<�������$t��r}�L|��c�3���뷳uw���㴥�P�ޥf|�
�i�X��	�CJ����v#�2����@�1X��ĮG��ʅ�*�u�:F`�̝���R!�Y�V�gH�?g!pݙ"=ˇJ�zG:
@��Rݪ�ǯ�޴:j%��2�%�%�@V����؋��;ҒN�R!ވ��J/m���r��ޓ8�2�)��J��p��+�U�mlz���	]�eu�����d��aoj�Ѭz�:ȣ�16p:�W�������	q6����:�q���GU���1�_fL�S�ٹ6�)��Y�0�NY�������yf���[����v���u��qw�)k[����^~��5�Ө8���[S�@�	���ip��k��4���c{7��8�+�%,ݿv�Hb�*PB�?ø&×���u8���,�dSS2�C�zMvs�Z��q/|gˋ��0��a]���L�`ϒ�T.�ԁ;�ĉ��@w������QzY�wl]>6-Ɲ����n�Tȼ�xv�J��n{lZ�~#�	`�R_i���[I95R%67����g&��L�enz��2��2D�0b.2�/�7";�X�-����w��1�ӴұG�4C�~N;�43�G3�a�̈
ⰾh���khR$�'����
�=��Ky�&K~f�#�F����y�ٶj9����n޿�,Y�� ����w�<H0{^��3QOöZ��4�j==�oF�G��w�v�W=Cq��4��b2%�ה��D6?�Ξ.v��U����EC�[yGZ���n��yK�زI2u�4�PR�����k�v�d]{%2�S��r���~zá�okK��|�U���9����@;/i�M�dѦ隷ɯ�(x��S�Y*�h����3�7sd�lP���X�v9;��y4ԣ�C[�������u�k��>�CI�J�d�Z!�ь��}��k�~�"�4ݔ%���L=��+&��5��	f�{����T���6E^�r�a!��74�}AS��2���y�'{m�:��Fv��������y)좔�ԍ�u܁�ߦ�[��Ty��ET�BA�-��g�
U�7s�,���4ds�9�%Q�$U7WT��<"A�R��.��WwsS�,�=ph��t^�4{�JW�uƽ�$�P;��3��t���� �������|hHP��S(txu�O��ǫIPL�D'՜��T�-|M�]75mӻ�����a�V�t7�!m
����dEk��K�R�ZPq/����{�/��nP�0�ƻm��#6.�:�-�`�`y���;�������gNg$�}����LNH�`��0#,l��E�ާ��*�k�x(��;-f%��d�	��{�yɺlX:9uk�F�V{{(���w+C8)���ƿ(s;5_A�N#B��m.D�;��J���^�:R�P�lM�(�Y��9Qe7�k'�v#ͼD�N�4��/�\C�o����/����7�����y#��;��N}�N���������sB��͔p��gδ�fD����UŲ��_��f�X!�9K��r�<<�t���c{�K��P��X��[D鎞�x�z�s"n2_�kr�wk���0��ǂ�)�輾����!""3#Z�v�wk�����Bۄ���E�h�_��ѡs#.�O��:�*�;vcb#�wa~uBkM�~��`�c�-/c(%�ꧢ,�n�ʛ�[��nE�a:;['������,��v1�*%��gA]�1p� ��D�-�6�g+PC{h�09hq��Y�Iſ�~鎟�����h}SZx�o��Y!�b���hG�l-�T�H�u�T�s�h�V₆����l��]q��Em��@����)�l���׶�Em��^2T1"�eb�b�̪˼�-r}{�ޟ��[�n�eqhE$���ʕz�r1yY���N��ըj�ʑz.�f*A2Ɲt���V���#a
vH3r�dMw�:]a���\�2��6�6YW�ٖ����#�z1����B�������`dJ�v�h3��h���Ľ����w��EL�3���j����� =����Nl�������2_�i����'��ﴛ�n`������e�:��m=�(#��U�&�j��߷��s�U�������i* ��y��k���]�ڷ��r)A3zz�&�T^t��P��+]��n�ZЇ�m��3g �����Xe���?n���N)��ZEu�ޥ^}9>ӫ(��W+�t��{��D��j�H�%�]��Й	pn�p���q�H��H�\��W4�U���!�x�V�mC������h`Alp���WT��\z����5"dp-����܇�9����W����q��	*�����]�!��+|;M_Mm���5�h�"z@g"$a惢����|��,�zJ�FZw�[j�4��2g�\�O�5�u����A	)�:�GE<l3��0��aE���6C�%f��K�]�Ӌ6�Rە�\KwA#{����ެ���P�1�υ~����_��7���x(i�8�#Dͬ��o\t��8,���,v��
�nU����}�'Cv���gHon�I*r�>;��.�y1o�mʧ�V\Җ��+6W[�0��J�U��N�7��M�������4������U��+�iIZ;*[C����v�vk�'�w�ވ�A{kf��p6�.�tDj�&�t�t�\��󵹍-�����͑�ӁZd�P}���馠 u�Dc�+�b#ռN[���Z��m��;3��_v{��x�@��<Wy��@k�[NC����[�v�\���_31C0q�4��>���|��kkv�K��:���ް���[���Uaqa�[�E���$�,�y�uX(�\_�#0u�=�Z��S]Jʩ�l��|,*�Rzt���T#��VW_�g<��6�t/8p���A�g�zc���Y�^�P�oLF)��۳��bH����K=e4I�j	&�/�� ]'���#dj/��c;� � g���[���O��E�koc�,��d�S�W��[�=�a��!];�v`���gg@�1�lF&L�g{:�X��^|�/�����J�u�VOE��u�z��vj�諊��モ��l@f�c1a��Y���t;(eٗ��ݎU7��Sn�����=�Ȭ�kH24�R�ﾙ����>����Z��}ᆼ$,�wӗ�{4	�~��{������=�n}�E��q��X���F��?[��UF��g�����sE�C�H8{^ �7Ս���kn�hۺ�.}�''a���*�����D�%�X�%�M�!#wÚ"-Kͬ�Pf��5�bC!�"/�F�OO^�.t����ɶ����!�"���ҜӜ'*!�el��a�

���T+pMx]FN����m�3��l���MM�kg��{m�����X��hG\�Z����;3�vAt�F9��eIJ��N�Ϋu5�=!�LT��@�R�ko3��y��,������s9$��)3��O�?$���oj���ڹJpP�A�=�:��J}�4.���G��%�N�=e����656k��y\�go*�i3�-~���븟7�>xò[�s.��K�!N��s7����o7vZ۱������/�X
V��\]T�o������J�:u*�1!Z�&��;�<�FpM��α�e�*X1=�4�p�w�� <�?e`��!l�66�϶��i*(K�mvy(�7?�:����e�<��T��s�������`���������snN�C���[(ԤiƏg��k�́�	����F-�<R��*�\�޷��!��prڬz�����U+k��a����!��EK�U�zJQ;y�j*�Ni���p:�$M:�dd�Pq��oo��^GU��ih�M�C���P�r����s�)�������;Fy�/g��}J|����'_Ċ�f��o
�%�`��;p�[�t_Y.ota��s�xx�-�.n�D��_lf�e7G��y����R�#QxM[�8�@e��2&�4�;�;ݝm�1�����[�
�:�>��F�1�F��g�r/��>�.wL�1�{�Y��t;���5��װ۝ָ��M���f�m��}�������7�u��O��E}���~������V�4�Fx�p�(�dEDQD@	   C�$�@HF��FR�F"��R��޵�`h�02Jnd�@����B �   �$   @ �D  �2 �� @ @ )#  H)   @  � $�D��� 30!�D� �       I   !�
AD�IP�  �AA  �@�("D� H� AE  AAAB ")� ��$DI b� �@ EH �D�$ PPQ�� 30E`�"� D�Dd (��FH "���E@F(��D@�Q� ����(Ȋ(��� �QE�"$�������DQ��(���Zb"" ��`� ��$��	 ��$��~Xݟ�JEt�ERc��_V�N/�_��ë�������o���}�wv���\Z�-4>ߘ�����m�7~{��U��{��O}H�\�|��_��y��&��.��'�?��u_"�w{9:Y���l�����>'ѭ���=�w���/&I
V1)Xʫ0̒�B ,� � , j��1���v	I* D�I  �  A�   	   � 0   �X@ʲ���(�  d  �0" 0�$�� 2 H�`d�"ʬ�PH�$ I# �D�� dd���#$` $a#�d�0`	 F,�0a"�$��D7k챚�>~G�����S0�BY�<'5���̸�xۣz�=���?4��yޚ[�}n��5ڷ_{�������nt�*E*�?W;ʽ�.��v%���J�u�a�\6w<�)V^��kJ)W�K��i~��[\4���>�{�l�.�skr�mR)W6<����~�}U"�pma���U÷��9ux�^�Ƽ��U��}�����"�p{1�5"�{V��խ�u^�f��.�?w��r�e���߾�R����8�L�kU�i~��u����ܼ*E*�[4��[���L������h����d�Mg���=f�A@��̟\� m�z����E  ���(*�JU%I*ETTD�) *�P*��T���TJU")U"�T��%�JRA���QJ��J@5�D�k@�QPI
$H���E�HJ�U$�B�E@�5H%*" ��Th4F��()	veU*���J��BI	H�EUJQ�HJ�T(DU*��(��(T)BRU$*!v�Ju����  ��i�m��M���4�j��
Sm����� j�"�B����T�����f�5�K-��m�Fl�43Jm�l)�d*��((�%(R���  �AF�4(P�C8w
(P�h�
t�(
���X�Fә��U���ѕf�I
�Z�e�Z�*��U)�c*�Y� �Zf���d�*TT��Q�RP��  ���fL��٠S,�����L�*�fUeil��`��*���j��3m��ցV�V&&j�hR��J����ERIU!U   �@)��PՁ�5�f�e�j�M*��ح�eT �`M"�1� Sf���V�V!T�1TPS`*"R�R@�*�    ���`3+�i��6� ՚klX�E ث �Qi�*�a�m���H�cV�d�"%	$I!%
�Qp   &p&�50h$k2e@�jm	���#M��5�EIj�Kl5FCT�ITQS*E�*RH�)*�7   �w��j`h-��h�����J  5��(����1�  �Y� �e
*R�R
�% Q;�    � 1`��� V  �F�5a� ІV ��L� �K `�II)J*�!�ԔUN   �`  6�    �  -  �` F�`  6*�  -)����0  e�$�J�%J�)E
U�  c� �0 `MU`  `�h VeXP(
C,  R�` 3  Pm*� ��  x)���* @S�0��� �7�<��M  S�A)J�  ���P�&   �Q	�R@ �@��Y`�"l��ش$Ǝs��� ��B�+�d}�;���v){着���ﾅ����I6�BC���~��BO�@BH�@�HHo���~T�s���w�Gr�̡D�a��؛@dD;�ըe��ڵ&�h�@5%Ջ��CY0�#rC�~6��@�j
�w��N��V[P���"��e���(�@gp[D1 �t�J;���,�&�ʁEkSӐJ�^3�UŖ��i���z���vj?�Ь�ZeL�pA@:zf��j�ME����L�>��n%x%*����6�a6rfTB��y�K.Uˉ�V��ޅ$�1Vᤄ[.��OW�*H�jR����2�j�̒�e�֕"J��m*����R-DR*җ,n]�ƕ���\�ȗ����B�أMGq�f\���\�Kn�v���b�-N��6T��hP��Ve�����Y�0 ��W5�1�r��.8��`{!�RiEl�3�m�����&��Y��bS�DFѥYr��v���WN���
mb-��S�SFݧ�����u���w P��]+��R���<ِ�����V���2�f9r�y���+�5����r��6��BX��f�KҖ�ܣ1Z�P@�x.�M͸�,��yIPo@Ȭ���=P�f���h�t�Z�9��Զ:ŷc�M]�n<Xm7���F�W�ګ�l�J���]j��ڬ�t��9,+)0�i��X���:6��@������fYT�]�����S����Ƕ��t�kwl0�0e^nĉ���a���,b�34c.� M�4�ݠ�{�)�&KLxP��Nf�r캽���%^,�'�0l$*ԋ��"�M�v/S�Rݫ�^,X��/jm��OH�@T�`�zIt����̸���N��Z���p屹@QjP���4��ndZՓ,�ą
xM���(�im��&VQ�;��sD�-m5�%�p������ެnS(a
��!�� �В�^���xe��`�+$����ȍ<�I�*���3�{
�GJ������ m\y�$RT1`)�"���,9�w�+v摃]���yv�1��e���
�f4]����W��ˣV�m���U܌�7Q3�# 8�VM�3&�E�r����ݠ����k0�G#��B��S[���40 R[Q�ݩES�,�i��Ͳ6v��^R����,�������S.��`͹A�z7v�� `T߬�T��5`#��a&���,!MMt%��b��R�hlU�����ӕr+�V

L����v�A�U!b�S���Ie��L�m*ͼ/0-����V�.�æ�<e8L�r��*(�ѥ+{{ߤr� �K�%R{6�1�Xi�y%,6���//r�Ĥ�Wb�1;��nJ���+
$���i\86V�Ϟ��2Ȼ8���cV�Nd����S3�eJ��,	�CjX�Ĕ�ݻk#������ے����`;���[3�i �*��:�j��j�vTb�t�y� ��\�m�`̺�J�MA{pK��ۄ�lS�H�BC1`SeљxF�M�Hm	 z4�
];Kgζ^�)=b ����6.�L8-M����!zܘM�IB�X�e3fճ���fJM��军��Nl�Mm�ƍZ(��NT�Y�oݵu�(�V�ej�ֽ�׉����Z�YQB�n
{��&f1R�ܿ���u]��D�V]�
v�+�]�Ս�'5��owv�J�5B�|��R���w�ffJ�
� a���������U���6 \��.[�������2�Y[F��K2T�e��Pj��敯�B�7���r��#R:����j�����\�[�XĖ�p,8ҺiX7@��>h�fJcHŭ}&Ib�ڙ��Zt�t��̅��S�*��˷��ܴ�[�l�M20t�M�q$�%ۉ�[N�b�GD&������/3r銑���*U��*%�+6����+d/uw[J���[��je�"�$A��\V���/͊ީaP�>�յ������<�2ȸ�Kua���5��p��m��VM��G,�����^�F�ٳ�{�!�	�j��u�c�Ȋn�j��S&]IjmI�(ljD Y�mD��I�Vn��L�ZƙR�I��T!�Om^Ɗ+�p�:�pK���1����X�m;4�2�v�5��٥6��g1��Dѩ9��M۔���!���*����oR5�mGI[���*�	����v��l]\�K�Kwl�a��"�7*Q�����D2�Y�C�\xi�l�yu�d�!��yD��6���B�н4�]Kd�n��R�k��v�ֺ�QyIYn� 4V�4P��j���omձ��L�7��2�Ч�^,9B�Y5f�����2�%�ȇ�w�4̀ɂ�
�.�s]XJ:Z"�[p}�>�B�=��$7��Ɏ%�,��waŕ�!w-V��Fht��ۡ6����6��ӫ�+ ��r� �k �"��y��;f@�r��mѱ��n�"�z� �-O�x�\k6j1d��%�V��e�v�3>y���f��E	���I�ԗ��F�h%�0n��i?��w>������
2�NZܲ��)T�4K���E֩��4�U�˪�iu-��-�wvT���ӣ*[�2m
C��4�+5�YP�ɕ��c����Ĕ���_ŨR۲/֛ۨmkf��ƅ��h�lx��a�-�t~�b�����ZC[�!V�_�u+*^��U��6+Rc�O�N�DBp����x��XM6��%%�[�Ĝc
�g]�z���c��)3fd��e�W�z���2�i�t	N���M��Z�(�.��ܵ:�J������6�4s4%�mKF��r퉮�Z�:��S�)h�"�t�t��D�V�ضf��o4���p6�U�5�#���`Ӵ%@�	�j�ę�$�U��o�i`��H�A\i��-�
8Nk1V'i���9J��jwE�D�2#g6��M9j� �n)n����[U4Zgp[PTt&�5��f����pX����[�0���d���2�]����T��oF�ͺn��u/1�1�N�ZՔ�Лa:�<�o$ƞ]�Ʈ��n�
,$iXL<S,�"�էP�cw4rY%�;���dGa6# ��ű���S�J�gVn�P"�]����6Zk�ߵ۔7p+PHU�t�d۬��n�"��l��ܻH彆�8)Q��I���֐pfe����MV�QMp�`�M���B�9�km*�%�{*�Kf�bk`�`�ڗ�9I�h&ʧ�Mb0/N�m�Y��8Ջ�d"�d,!�j*˄�K1���;���D��Z�*�*� ���(A�j��2;f�-�ӷ�����Q����$�^d��;zf�2�En�me꣙���Wk8i����tc7Z�k����*R&��PW��@e�l�f�tK��r��wx�^�1���r�]c��n�N��6��-6��z!a[(���˛m\��&\��n�Z�z�)�����Kv2�S
#O�1���n(w`�َfc�/1�Sh��Q�ڭY[Kn���t�jХ�R���n��rV
�5Ԇު�64�Й�tm����+_��� �|eR[r��ѳke�[��dMSY��q��@��b�m��4,^)1�j��&�l:@l�2�a�PL2��෇#0])�����ʏx�������m��`3%X�ǒFD�!W�AV6ܽǦ����S���V�b�x�n�[�"�#��[������Ť���T�kl3�-jG������.6U�S��K92���8��h�֦ӑP�����{d�W�u
0ؚu������C��{QID���A�oe���N]Ŋ�2L��8uk����6mGh�[�����O�kJ��vk4��ֳ޻)��3e��\���N=��Ywḙ���������f�8��5d�K2۹ea��c�քX�j��T��Gu����R���55�VV�����%ز����J�PR	�R���SZdi�r��A�^hu���k�{Gn@��)T���lL�i�u.�h1��o]�JhVt�C��]��q�j�Љ4�.���J[��Ƅ�eˀ[{e��jeA��V@,�hb��fXb\��(J�If ��[�Z�%,�,�q�ݺ��L�˘�obw�g7����9�J���fD���zH��ѼN�t�块iwl�F.�<9�����C1���b՛�n��4J�m 6��DUi�^jF��l�2/	�I�܈ڛl"��"A*���V�����Une$�ʱ5fi�˭l}!.��Y�TB���Y��̤��N̨��˫�0@˵[t��$��
0U�s n�Y�t�_�y�7/�*�v�{�z[9B��o(,�]�Z����W�S�Z���U��J'�%����lm^�C! �t�t�e�+K.���C�6c�V��8��S��aV/�����@���(V�s
�7m-Kqf�H���f�7�Ze�ط3n�� �i�vּU��]*,�RdʼNJ�&�{����&�-��mI���U�p�oo5jn�Z!)��NɆ	�n-d��
�d�Ѣ��*8օ�S���q�X��ic�3 y�aYtҹ��!��u��fk����m�Œ���㨔OI��y��Պc��Ў-�6�d7DQT��v�����FU��2[w�M��ˡS��Gy��4.�9�р��q݀�eR�[J��l������1������!-bi6�����淮��-n�hֱ.��1���fHOu�ޑ��U���7��WV�f�E�>WM���^P��l��I*b�˗����O�,��!��x��cxi�M�-R��pꕪ�-�]=�7�hG+��RA�<�Cb����!����yQ�Haa��
B0٫7C������$d֜rf=���D�h�t"u")�(��	�~�n�xS�³,�{��oi��Ne�-��r����N�K�y��D��e Z�u2���3+q"�Ғ�C�sJ9.*�%M�/�ki�mF���?�d���nn��{iW�n)�%����،��AdU�z1���ja���Y��^#�/n2�˥�H�!,�v5�Y�e:b�1^�˨ke�-���5�vm<,5�[��j�����$՝��@à�x�u7p66�m;��U1�Jok	Dm-�@��LZҌ�#LS�$�[,���	���G^�5Il����t��F��76�%)/�EC���ϳ��q�zP�d	r��y[u�*[pJoŔ�[�Vd
�9�*\����McWnm˥�C%��5���Y�rͳ�m��FӀ9U�����7X��r�����m�`�h�C)�Ƶ��J�XF�J�
 �{h��d���=����X��n�ELr�48�ojGwL���J�@�v�l!kd�/5�%�p4\�X�鿣n軙p���^"S�5���BL��n���˧A�)!�	�qfV��E�>��C/b�S���Ȟ�$jKŸw4���It�5o歺�C)��H�O��.�mlIS�>o곊���$b`-Z�!I37/^������х��9rd���X!Xۼp�9h@XIdX�bu�6�e�f�)���d�v4�r�%V�����2�SY�d�*K�)����,����y1�jU��6�])x�-��Z� ��1i����N�1,H�u�wu���ƫ.�P@˻��Ñ�p2)�$K��u��Z�梯*ʳG$	�1�,en�Vfh����n�	(\��Cbe�Z!G&����Cgƙ"��-B.�=�T�$i,e���+N�7�4�T�X��+mWiGBU�V����Mje��Ī^�.�[w�D�A��7�
v5R��Hݨ��n�G|6��l����"�c;l�Y)��L�����w�]�o7-al�����mT%+k*�[�o72�F��F�`F���.�1�=B�> ;D��sN��9OA�!F�t�O,*m��m����_d�%[��Z8��i�(G����$�I�]��F����b�fU�ChKۏ�4���kt|�V�y��$Vw�F�%cy����Z���0��Rhm̦V�34�PM1nP��-�ay�ՙ��Z=dܘl7&�������i����l�"e��=U�P��sC���Hz��.�ҽ��ڵ@^�#tc����Fqɗ��;�m^�K6S�M�`�v��rP6�^��Zi+Dˌ��h!�*�w����H�KZ�51[��]��D�i#`R��q��9E;�쇩-��Ʋ�(�f�iY�O�w1PW`B���Z���2�(�j��Rܠ�Ў ��Zb�Q����W��X�4e�]5���Mw��x�t>T�&Q�pS�
P�RE��Ժ[�AJ�쏛$�D���ښ�Q�M�d�.�b�ABэk6���W13gV�<�b5x�j�@L7�'%��lIp�Z1^)(R�4/F�GG	ŋo3�6D�;a/�U�t�=��S������Ǡr���HNR����,�̕�C��&J0��OQغ�S6���3��P44��+.
)�Lu2��34��!X��ʷ2:בS�!���=T\B�G,ݓ�&�s(��)�Lژ�6jyn�P{V��eLSY{X����l)��W�5�)�$n��DCM��oʖ]JF��)\��ѵ+YL^��հ��h�R�:�P�1	T���&�^����b����C�,����w����>P	lVVց�w�04鄓�l�φ\�k(mcՊ�T	���5�]ca]��Q��JR��i�@m�y�$�)�4�n���OƁ���icF��0<�J��̈́�V�5Hvol��y+̢�o�͡�3#���� ݶ�,U�$�O@�����ʗ>�G����r֊ˍ�)�f���j�ƖU���lKCC0J)P#3\�sv-m�>���8ʮ��C���U���}X #n骰OHw{���T��9�.�V�[�kn�F�Ω��Z� ����DFT!�j��H�p��N��+��9u��������̸��S6��_u��ov�))�f�͍��T6.rד}�������ү�T�Β瓠��@wh�喴�v鬮���n�j���Ya������oyB�q]r�S9�)�N�a�(t���j׆�?�nA�8�������n�5+��͗[����R4�k��J󕭹�0�x�� 좣[\s���� �.��D(�������/@{����vc��԰�M0�[�1�<S��ٷw�hP���w!X�e�|�����CZ����k[/#��h5����P-L<_N��:�]88gW	%RV��cq�yk7�Z���`'��l�c ��"���k�	i���-�����w-�����/N\I-]�m��Ku,�N9���&嬗Yo7��5�!om��%�­�;S����ۤou�=U�x � �����u�D�o]��[�3CM�k�}\z��.�]!t_0	�@hsY��=����NVwR(��;e�����/�
�a�<OUb��A���f��Wǌ�:jVJ��wk���G�;^mhs��m�2>�e_��)�KV#.�^̟q`�wn�	���y-]���*Y)V��WA�qh���_*(oa;gb�^rt��4���oP,�k����d
u�ƅ��Zl����sox.5��S2�7�-�M�?�OR�z�E��>zΈ]�e�.�٤E�f�'ӻB�8l�W��rW��ެ�2Vr9� {iw)�2�j��lH�-N���ѳ@xu[N^���]Qv!�!f|���wxxB�q2�Hȳ�bH�S���I��J簾خ�s/��	x�_RY;:��f�%�{B]%����-d�\�w*�s.r�d��w��#�Z<:�qk.�V�,���SHB>���'U�|��Cv�;H�v�h}��k;}e��o�)��ޠz3����5�tկXw��� A������n)�}\	���ox��nT]�.`�=Z(h���~�k�|3bں9X"׉�܋�+�Y%vf8���1��jm+��M������n����v��P	C���t�cb�fM� ޖ�GI�V	�&:(Ӄ��T�@3�K�n��si�WSx�����u���tY�xi��I5�6��෯��+.�K����!��r�J���#I!|R��������`�4OG]��3]v���pj��y8�7yݪ`�8G���].��E��Y��-�ϲ���o5$C��6[M���,<���m��9�ϧ�0,�Q,��Y�.��Fh���[o;8�.�2���u�R�VF/w �5�w���d�w�[/����tg��,QU���Z9ݪ�I)u�����p�T+Tԓ�9��h�ʜ��KY/Rt���v)�8���DsD�fҍ�hy�:l��T��inT�j��`�]�`9ق�̼�i��bӧC����L[�ߵ(Qѫ�@~i�p�5�������S���yn.�U}�e=U����f�)��K�GՆ�����哃.�X���e�g�h�Q ]�.�`X�M�.e�S���cջ3��7��,��dحp6�ӆ=9r\7	;yj͊�T3;�D*��4��\[ܭ��7�u��v4�\G@٤�5�E�����K@X����Z��=J�'�'�V�oj�_�������\��B�i�ih�����Wd�q��(Ri���7�3u��i���5 ub`X��sͷ�/F>GP�Y���Q2 �w�ra!�h�fK2;�(+��hTw�"�4��b���B��o4��w�.�j��+6h�}:�KM�5Mi�iͱ��IC��rTE^V����Q�l^5E�+��'��h�6pU���C���3�b��lђ�Ǽ9K�$�ߚv��{}���q��u��wIcD�6����#{j�Np���nꕖM�ya��`�{ok�c&u�:,�����B63n.��Y��s��,��c-M��`�W��-�/�%ݝp9����;!��j�\3/+��3�JK���6Փa:���;�@6�VG��m%:���}G/X<WImu���F^#c%�ym�ܫ�y���M�u�aK�O�y�8�ъ���K
����|W5�5���OSv^s6p����{�����s�����A�t��f����;��t��\Wi���x��`��.�4�9V�����]k���6�;(��|�@2t��ڀ��0b,�5u�qY�j�Ҭ�{�k4��:���޽ֺ��-c6�v������E�ٸ��@�?%�1h���u�&�d'U����V �qV���Zΰ)#����'YWDC��Ht7��ww=/�ôo��!��Q�:k���Yu�z�]8;*��s��9\���ۮ�+܄�(]�=�*N�	����`���l`��U�}��BT��qv��3�deɫg'�b�g�
ݷ�7�����D��@�DoJ6�sy8g!����KҲ��:�T2��CE��7xu\�mʖȬ�2��񾀌���"6y���r��t.v�8��;�_h�7si��c0���'�E��%wpJ�%�X�>�2��-Hf<���ׂ��Ԫ�[��c��!��������S��7(����.�@,8������q𭮅��ƨH�OF�j��JA�ׇ+0��n�S��#��K=h��=�E��DLo�Ö/��H���/C*��s����ƟQ�&�Kyۍz����dFd��9�κ��R޷g����rWn�F��u�m`}��=�`搰`Ͷ-�qgW.7������M9b��X�AE�)6d���ֹ�C�h4�]�,��vQ�����J0�m��oWrݬ��t�36�����u��'��D��O���b�\�-�$�wϮ�)X�ppC/rV��L�4�+p�8AW�P�<伭�鸶��r���v�ut:c�vi��i�� ƕ��|�����}��X�+������βx�l��w+$ ��}n��T���ot���p��H��4��7��5v�.w�#5�������G��� L��
���C,����\����o�wV]��R�b>��N�Z����o�qzan9���4ĦR�F�;qv�V#\�LoԢ��	+]1�k�i;����+�vv^'�w�H����9_$��u0�C}�j��=7:S���; �#dg��ԙu;��#W
]���Ŕ�B�K���󁱐j��i�|7`컴�L�F<�D�w�'\�Z4��hAH��'0h4��-��f�U�k;{�\�ym_�I�Ը���Ɩ�9�'N���9��0���eΛ{��m�V�j(��m�U�9i˸M̮��2ڟ7�槎k�y\�npo�Wʞ ��*��%V�=�I+S؎ۊ�*�F^q����*���y�YO%I���o�h��/B��F�`V��U�ܴ�Φ7Q嗔�1��sr���u�=\�h�L�Q� l��@���;͡��](�� ���3���T����[�,w�аr#cF��C��n�M���`�]}�w\���:�r���q ndw>�Ky��J��l�}��a�k����պYh��5+MƴU���U�y�LLwX!gKIŖ��SP��qw�결�����*�-�r�h��[�p䔢��N�AJy�X׶�^w[i�3����_K���ԵW�oWnA	�B��s?nQ�wڅ�����j�S��̭��1q9��@Fe��&��FVr�խ��X)��loK핏i�lд����E��B�wu�������[qe'�0Se��2�@e[�6�olIQ����@O8q���yf_Zq.[t��'V"N}���|
2�w9wzU�:�M	5|�DB�d�c��Mb"g��L2�ob2����]�2=&�WmD�m	`�.�VT�t��}H�mrdf*��w'��m_oـ�-T��tSr��ϒ:m捨4��[zؑЗM�Y�>�Y���93�i�y�Jn���=@��L,�:�EYt;�0iWdB��tCiqw��ﶍ�h� PX˷��eӽ���oY#�]�ے��8�kW3�Z��^��v�T���BE�6��Z����ȅh��M �t`�R�uF�:�=Gs)�je��*�6x���k~G2�h%fh�&�cV/Wv;�W�HX��]N����Pb�\&-�u�j�y�Q��G'R��{L��s�"�y���i0���{�ר���+�uú8t��N��e���<���K�Z���y�u]9u���h+XP:�u����ɱ�=�l�J�������9�^P��k��I���ӭ�GHe(&�*�c�j�5L��+��AѨ�
S�4��q�O�>{��G�a뭤�4�7}y�R�[��(ݴ2�[�x)�=Z� ڒ��I[S���w
\���:�XU�n��R�5Y�Ȭ��V®�}'mwz:�sG}���륻h��V%7;S[�wP�Ç������S��IJ#���*�\*��OKݣ���s�0���p�j�|D�Xw09��X�&aM�\�V�MB���7=�0��U���=/t�A%3H�+y�bҺ6�9�G��Ι�k�E>�ެ�_ʸ�V����e�&���y��5���ɻ�V�����C�.	���e�f���2�_];K^EZ���b)G�0�Eî;���z2�K4���<�;jN%gH�X�&vP��hx4�iw9�Ӽ(��V��V�kD���F�ͨ
MҐ��\�ނ�޳�����Tt4a�b����젰Q�سO.���d ��������%�֘ y�[ug=:��!i�b���]�Vʹ������L��q	o^���]qc�odT��e�f��S{�֮�Z<AN �;�w�Ƙ�RJ�stzY��ܓ��7D
��9���!�V���}��(�fV
{�� ����<2��on��V��K�׵�g��R��uz�]6��M�a�!
�����&��`^� S�F6��ݸ�ZU������]��
���t�Ҵ�PT���m�]q��k��-��Ӛ6�����[���EB��`�@�nm�]١��mrl`�OK6�JV���"ɫEA��D����	�d��+�2�^�H�_);�'Qѳ�T�;m�/I
��j��̣Jwt衕9O`��rS|�kpl{܌�U�^<u���a��-u-{�(5tﶺ��S��}�^c��c��&�TsG=	�M�c�j,��]ňW(�\\�N��vu�4���n�H��"���;�*,����I�W�q��}.�,2zu�0������|N��.{���m�\y1,gBc3�����]���S"f��d�[y�rs�6q��h���ʝ̔	�
��i��oy*��c�&gb�U�h��[3fK��J���:+Cë���	�m:��%㵳�
H�pG��n�^^_#�
���wE��eo�G/��]��8�����a�8���մW����׸����=��}y5�M�fѢW�ż���6#�h%��K��n���f��vur�0/y��#z&#뽙��G/�.M�.qbw!K9�t��;������Ȋ�o8��#���51�k�Ut����vsUq��p�6��gI����~�+u����TQ5ڽrr��-!�j�U�h�x6�H0��"VE����9
mڜQy����i�H���z�Y���d���[�;{�;�(zI�w��ҞS8�»b���K�ˤ��������n��;���S�|�3bz�1.r�+1v�
b�H�G���3r�[t�ub`RN�${c����|r��֥��#�͝�k�S멦�՗ى=n���TΡWڥ�;�%��<3W�\YK�<�G�,�DVVj��2-���q��9j��/u
�)��9�w���t��2�2��}5`�LZ:]!Y�.C�6����.c7��|FaL�H�VT��q.��"�k3+*�on4�h��MQحRq�}0'o�p*f��%����3�i;����od�:�޴��4q�O�֒7_R�2��'vJ�Dָ{c{OK!`tr��Ր2���VAܩ92J�<��O��[��Z*1��ԔڻެUa*��c�[�.�gj��УÎ'q;1��9����W]J���1�.��U��V�,���өM9:�`���Y
�xJ�W]�'=�&Z��\��S�
�6&�4�?:�9 6�TU�9��8���Ut�N_Zf>�q�Mᕸ�{��V�*[T�;wyHQ�h��bu��b���rr[[iS�EΜ�I�P���.�߮��!t��FEVB��ܡ]�v���a�K�S�E�iG�T<}�7m�ז�ߓ��(:�1�x@dՊ��hU#�Fԭa�@�[}ˇ!֟vG'vV�|��'\�-�z�@�	������h�%���Wt�{�8x<�w��2+�b���Y�́����L�t�q�}v ��!ݖ����]��}�+�e6+���Mn��Ր��%�x�4����r�6����Zr�#��&s%��M5��ј��\���Ԡ����]�� �ChkwQ���v�+��
�_#|�g��V�9qR�m�go�<��Wаj��
�/b6v��^�]���\�;�^T3W;
�]�P��f���p�ͅ��`�Fd|�������W{��%��q9ƃ�P	����.����Q=�� ξ0�����g�������QlR5�v	s6;�;��mbN�ik�a=�բ�S��9u�b��f�'qŻ�qc��#e2E�58�N�d9�w��p��9�e���7��5�����J��7/	6���S8�9�y����v^� ��L\�8�W�<��#Yv�ǧ����ZӜ��%���:���rk���f���%�RI%�l*���(�>���$?d$ ~B@�����ǌ]$�-:�4���<h�IQ��dp�ʔr/��s�[�æ��7st1���\�qH!-�݉Wc����r7ۺ�v�@�M"#N�АCpL�>�Sr��+-���F{5���p;��P�W�֥��nr�zb幫��|+�\;A��Z�]^�3ّ��m�\�9(Jˬ��V���(D@�pv�X���:4ko�K��;�uc�A���8��$��lLl�s�Z\��<i��z�+v �ʻ���d��0�U��֍f�J�L����E4�uD^�Z�fYN�nG���q�e/Ue��7K�%z���jZb�����d��ui�Md)�]�f�ӗ֥
��PI��I[V�¯;Ev�o�L7������pA�v�JI�����u�����V�$ځ���e��
� t�k_c�A��H���EN�&�����+�%;5�Ԩ+ש�x�/����u��ə����"gkɯ�>Sϵ�fEWp��*)օ�l������ך]#���7�ܬ���j{D�Y��иow0�B��R͡\�nR�W��dUܩ�&c��fUv����)�ܟc�uo�ꇺl�v�����h��$H���n?��)v�q .�7)�b�f�i��V��F�y\7��W���-�xK։Xc�n�z�KGs����=yw.)e!��r�BX�Rق1a�ؐ���>�B���`^gV�ԬT��(���;{��Ze9y��\���qHK(���kH�:���.��&���e[��F5ι�'q�
�����J7G���9>�L�ƫo5qh�z*�L�ܧ*�.�=��kr]�n�N�9���3�vu�����Ռ�tzf�4f��LK��xk,t��?��s�e������s��!�����5�kF��'1):s�d�+A�}i��!X�^^��W֮]a�����w�6�j��½A�ŉô�-�gV��씲७��}�Fdh������ZU��&�R�ی`�b���5�kuEI�76ͮn�V2�*o<�t�&^��j��EP�&����BWp�ܬ&�y]�Է��CW��w�wZP�m5����׺)^�ڊ2�nG�e����Xw�4���.r:�[��Z���j�qO3(r�k���>=F���seKB�j�']��7
�5m��L`;��4�%��H)f�@�/�X��4o��r�}���p��b�����5r�a��ZvdY�Z�˦��K�o<�r1G�s'^�m��`������a�W��w3Eضh�Iv�m��QuryR������R�3Pw�vJ�yl"�퓸�ޣ�pL�c���G!�f\��K��Q4��Uӂn��buZv�FZ�E�l��+�V\[H�0�@c��9I�;7�¸#�������VF�^��j�����9T5���r��b�{�OS�a�z��V�Ē=Θ����(� �eV:�A�-ݹ�uAy��ܷ��2uk��X&=��wqe��5�֎*Ro��S�U���Զ����GCzwpF�_)���D#ۦ���t�^�e�)�6�wX���YӔM��|h��Uo5���e��w-��v��]�WTw@|�kf�*b�ݦ����ܫʣu#������-Ky���oe[��׻F[�Iq��.��׮�픠�;��-��L�WGX���ss�^"�-3�in��OwW[<v�ţ�#}��U��s,���\5�M��PC*ذ�F�$�R��72��3r�S]�#�)���Q���7{U�y��o3���6-W��;�Qr�U��*.�Ԏ�tF��*]�C�p�|�+2��`v��mՕw�2���x�j4-r�L�]W�ms��+sW/�<lSK����F��6���ZyY�%5�:�$%�ۧ��9���֞,8hd�k�s1-��һ�u����K���7��v�gl�sD�8�[��sk(�Ϸrn+ϋ���r)�(���#׶!��nNv��KkJnc���r‛v]Nsڧڪ0;{"Q��f�/	�m�΍�wA�I�W`��`��(�J��uui5�r�]���*��+,;23�"k�H�Ɨu��Z5f��a��^a7�ZF��jvG���LF��S�3B]k��&����R�8'gb/��b;�{���� ��V:j�W]A�;ꐩH^v5A�*7a��L\/��tuw\�J��$+���M����8�C̽Qާ6�Vkso~R�ͩ0ۛ)�,��v�Χz-t�fwf��USP[Ǭ t����8��GK��*:C��nJ�f�Dm3]ʤ�})f���w)sr�rιSq��;�u�v�}2|t�a��([� G�k��֮�Ջ�q��c��Yõ��X��x���T�sB�Ts^�BX�\��8�b�X���_��Qx.i�s9j���U��rcU�3�Q�LZY\�cR��D]�鯗W!|hYn9f�`��%M���-��gM�#�hJO&h��_���U�9{��j�c��$� }ZD�c{D�3sj�'x-�y:�&d��Z�D����^H{-�B�l]b�L�œ��	�h�*q���Z�O*��AU�7�� �LY��/S���R��
�t�������w�'QЮ���=�����]��:էw�c�C�h��gا`��g�}`a� ���afq3X�mN�M�n�T(n�rt�N:��;j���_ZM��,N�u��cK��y�S��ZH��&i_cw��Xp������}/[��K���л�02sCo�8*�%"bY���..Ʒ*˄X3��J��\�;��w͋�ڑf���T��̤�g��u1
�ӭ��
����-ly�����E�Y�0�Ѵ�*F�v.��9���сw%����u��b�6pr��$_w�NE�]	�G,��ܼ�e�i�k)V����у�lJp�`_>],���Ci'$k�䬈V�b0�[Wx��w��YPa{�cnodvH���YF4#Y�'wGv�J���Gz:�9 ����-�Lr��W.�#���J�罢��8����J�TO*�\%��I��S���41ݟv�M�3���Ujf�'�j[W�)]���'����'�����9�]L����2�K79Ii�	���ͷ��]Ӯ$ըU)��p,�'X�LU�]�����w�l[ U����]I�k��|�����Ī��m��O(�;�\��F󰾒�=��M�aȸ�ٚ-He��B�j`�#�<�A�`�W�v���y7uk,\��}H�p�{�*q�Q�.�-]�y��Vͫp�ZJF�rg	�����԰�h�R��L����ˡI��:a+e=Y�:�DV�z�����3:<���m@:��%���9��:=q�Z��9t�ڽ�֭�Y�[�q�7�;o�wd��˔K*ұUxi��]��l^�b{�����H�j�-������]XX����:�F�c�;�@A�#�^���#qT�xfFN�B�>�׈E201ޅX;{ 2�H���:�]ͩXa����Z\�qɽ�N��Ύ�ٻ˸�n
T+�H���]��RWm`��͛�Ȟ�G�h��u�c
y�M..�-s�(d����t�Ai�v+�mŵ}���cݚv���	H��궺F����ݙS�Iܾ�r7�yA�w��+��e�̣`K���
l����S�}��]_>[-|���j�����P���X�|���9�KVc.핆ڬ�v[�0ŋ�����@�FK����L_b��l��42M�����]�N��g��m;��:�um�us���Nr�l4���{��M��ѝJ����i�:[�BPR��;%5k5fe�t�3��Ԥ�bw��Ր�����Ѹ�뽜���]��7�n����`�k�XA�yf��Uv�Ʋ���=U��g#0���Km���,��GU�Ʋ�,��	�VgZo�.�)\��5�ҡ���|l�t,�yk�����TfM�A,��j���*ݝ�R�K�+8���;�@�O1l��Q���*�ܽ/�R]����;���g*�U��d��a��}LLfs�v�s�.fکt�}��\�n3pT��>���:�7g��Y�p�ބ����f�,'��\m�ř]F��5xl�=\R��ߎ��V�ԥL#2չW��p����F��V��h���k�NoW.�5�T���&' ty��c�&��\w3�SA��Q��7WV0���[O)���<�qHG���7�橕pk��$�G���f����p�7_=^sK�+V��͖o��f�/^2v�1Rb]. N��A/��c;R�{t�T,k�6j��+�����5�9������!,`}�;Ⱥu?�PV���pki�*[v�b;GkI�W�3Cz�r�qlm��4��5�'Acj�n�v(*v���j̺Xr���m�b�&Ɂ�l�YN7V+L��NX� �Ȩ��|��]�j�2)k�TFz��!\�U|���\W2��)�Z.��d�X�R�0+�f�^o���Z�_
�8�D7p�T�+7H�V���2���FN�7m�r�6�B0�Lfn��+�o1J��XÀ,��)GS�Nݹ����sUi���R��s�<�,�ڼU��EM�Vk��^qhKXK&�F��)i*s|�"�b�E`�S��]�goc�'n��e��+���8 �.8�'�\&��e��ΫY�]�u�jiD�M7�Zx����I»0�|��!�z�0�ӳ"E�9g2�u��uݕ���A.�v�g+sK��Wvwc:��*�[��|\�{����%C�Ho�+�T��y�J��u��ۃ�]��R�7��Wd�m�@��b���{\�ԟ��f�,����, ���*��9���ǜ�_ �rXu�Z�]��ES�R-
�۹Ն�=dvǵ�[4������i�;xY���ѡ�.sG+,�|����"�dwe�R��-��e�K�$�5"O,�lY��T�Z����w˪:t� ��ƥ*9ۂ��k8n�i�V��v+��;�O��7L�@ `��c�0���<3��Ur@����jՓst�&23+!��T��MT�}�.�s���貺'�o��>�2�JV��{�)Lu.*�-Q�V��4�Xuy���6
��"�}|W-9R�}p��\;k�ۨ�x����;���j@S�o���{-髚*��*��0I�9ê�V��#�/y�U��K+;V�%�u�*�1�LôBM��ɃZ��u����	+��C4�ouK̀i*6(+Ý±fp�e#��T�V�ز$�uj=ޡX�f]+S��j��p��Qm=�����9�;��VR/.�cS��b�;��%�p��ϹH���/r�v�dת�3�\�m�w��>�}���Sz�s��/�c����v��.�p�u�*�H����~O�V^˵,,Y/\�������Y�(p<�Na�)u�ѺPٝ]�:*Tw��l�zf�SM jDe��n)�+31���B�#�<#��u���1l!]&%�Ǖw%���:�A�ޣK�9оޒ3`�Wm�#9}ζÔ�hݩ]��w+խs���u/N�4�`���ܹ	k[3[�+k+3nҦ�z-}�4��L;E��6-����h�t�_d�ʮ����P=��3�ܒ��3g��q�	4Q��^P�2ģT�j�l-�d�Jn���y߸��4N�@�
����x�f�2NZ8����ֳ�E�1b���6�.-�gT��pu�+/h��|�y����9������?8�:ܭx�YK����|���{g&�v�b��α�"8�J��==�Gh�%���c��3�v��@����� �#�ʮ��+si�r!�3���N�`j����f[�|3@T��`յ�}*ի-]v`�|�w{8;Z�]mi5S\�u\����֧W��З�����=o2�s^2�J���.��2�!
�V�Wä��i-u�b��/G\
n۾�����ݧɞִ� >v7o�Y�'�ii<�t'{�i�P�;��Xƚ��o�`��1+���[w � Ӑ�|]\�|�*Y�N�q-��e�R����!&;RmY
��v���m_#n�[�l��'qto�r�ˎ������f���J���4+�%�t� �p
�B�|�v���l�m�n F�@]�;�</)lq�]�2�`�2����U�%۽��xyE�g-�g�A��wC���J�Ԯ�(p����o�U)	��)Bu�Nj��[���s�]��� ��{V�f=ܥ��瘐��9�z���=�lDwp�vY]�`�ְF�&�B�c$;��0�u(���"kT;�m�
�o�U�Wwt�eiG�����#��ch�������}�^ ��C�n��d�rU��IW������mֈ�2b�ѰK���!�&��MR�6QZx�E5�=��E��Z罷�<�wB����S��6�ް�۫S�N�>{�8��җ�����ލђ�jÑ���'M���F�ղ�t(u驐H5;*�+�sI,�Z;w��eN:zV�Њ�^�����Tt�H�[�X��X���]7j�������q4k,Jږ,!c4��W�sI���ہ�6�3v�F�]��@���8�\1��嫌����)%�IP�xq=*G�9����ҍ�������S5n��t�wd[I�,�'5�و	A-mDn�r���Nn�����Q���,��ݼ��2�Y�t3�&hmd�I|C��N��-���G;bŗ7�]1�=� ���_-��l�)�-��pG_ju4N�}��b�^jx;��ڡ��
�6�lIQ��/J��)�>��Dgzfue>U1wPݲ���ܩk�����fS5wX�4+e�Oeպj9@ݷB����/]���<ζ�:앝�0rw�����Q�X���t��17[�E!�����o�r�� ��&�}��������;]T�nf�Ԋ7r��ڶ&�8�����5��R�Fv]���Q��z�Z7ٗ�ѾO#4o+^F[Lvft7+�-�K@���s�`7�ᇰ<��ʔB�^�j���K^�y��FQ��NI��W#�ڇ�[wτ����C6�k\d���̝�b�p�d6i�/FX��*�s�7}V��c��}�2�;�j�W��tՆ��ZG9�/E�TpSŒ��}�QV�[�~i{ܮ���H�=��,Ӷ{�݌��i���"@$R����7vpÖ��`gh�;�8�u�=֯���;�q�87wJK��v���;j�n�;�zb�5�f�hY0���s�p���&K�����6��\�Z̃Ge�E�OA�Q�i�����f�gj�������weΩc�rp(%o1V�%�����ljv�SX���L�WB'��,���*u;�:�r�|͢���ʦ	��E���#�.l��@�!n�>��n��WH�l�Az�n7���{5��7�f�����k$�U'i�
gj&J«h��dw]��koR�br"�����k��"�c�c�GT��7v����w5�@F{MǎMk��Wo11]��-]0IY2��O�kV
�k-dG6][.�r��{ҟZ9_�A*M��~����y�q�)Իǻyʕ����f%rfN���m��� �!Q+O�W,Y"������Ӥ��-ԙFr*�)m���I^EV(�.�C��&K��Yңga**5ۜ�Bݨy)T�I3+vET\$�I=Bmg�v�FcJ��/LY%&r��Vz*ɇ!�u�v4%7@ЭM7TR��I\�*Ԥʈ���4(���#P뮢^�Ӓ^IS8Ry��"dR[9�<a)�����'k�]X��T53�Ӭ)��g��1��D&�T*%�r�$�"�Xrl��"Ȉ��fL���p��m��XV��i�r�7��DD�Ü������5&�&���h�h��T,��V���,�j�yZ%V���-H��6�\�4fL�r�e��M���݌��%Eu�QV��<����NĩR�$� ɍ�B�r�֊�F4��4��Zq�r���g��i�]n�#���Q;��.�Ѩ����c��T���Xg�>u:B]����X�k�+S�V���kj��{Re���Q��B����z�ˮ��#R�w��Z]R(Z pFC���/��ޣ �~���?���~�"�?<�Y΃�p�h�������n��L�kNn֕��F�E�On�s6!���b��B��b��Wa8UiK�嚇������֭h�E�ڿ�L����p�N���tf�F,5�!�'l�:A��9n�N@1��� �d�G��2�!�;�%V;�+�cn�t�0clm�8�U�j�88�tTE\�����0��T�/���.�=���6�WyjTwO	�oi������."�%;��� �0x�)r�T���"���-��0�|��F����چ���}���a'��������b��N5�o�k�I���K�����n�θ�b�*cs��X:LL#����=��4���b��Ld����t|6`e�%+X�#�^��q��!��4����:�M���A�
�Ow� ��b�[L~qR�>�A^���F�*�eڱ�b1'�h�oK�;���}kk���z]�2#xQ��л��-�݊�
�N��{��N�g�xD�r��®�}|.��
Y&���}q�,��n�߳kW%�����G�d�y[�v�L��9�,��z�^�E7_-�-�v���#J�8��_K�B�Ph�u�@�}^�5��"��Uה��h`�2@�7X����_ �e�븛�z�'M�F��gm	���ou7�Fr�[]�� ,�ɋ�j���F4<�5	^��4W&�-�'�("D��3��� [x�^�W<��ț���?{�Q�B�v?��g���xmgqus��^E�JeMˤ�2�Q��_v�z�? 0A� ��ꜗ��Gx���ج;k�^�1�U]���wT�k�:/�yX,�d�M��uC.:b�<a�e�y��AS�]�>�w^���v$�N2c�ꫨZ��F3���P�T	ۄ�l�qxg�`�0�����|�R�Tio7;QB\�pJ��cb7e�{401|��B�#�(�s��Yx,u�͓�Ø��QmoD� T_�K�b�����C[��Y�s:��C�2΃q�:|�1���S��u3�vڍ}r˫�곾wwHIV���k����Xi.�:@�}|����$c����J�����ck����t�e+l��k�b�?7�yW�(U.���`����t}�����ڛ�]39*ğm�ܧ`��X�#@��謭Ӷ�O�V�تZӝ�՗j��㺕:�
��A��
j�ckZYu���y}nwd��w�n˧��K�X��:�7��K����s�j��V�-_�+A�����R3�!��lˀ��7�	��:r�!��7�g�{��_l<���:+3|��ѱ�&����ȟj��$J���ZAg��)��3��;}b��6��VC�r1\v�����P'�fĎ��FV��e����K��S}��\k�Hf|X�j��B��b$B
�G9ɥ��r)�湭�JfXD�����q]u�RY�E�*]���
�LC^ʖ�U�+!��m�V�ۑn�F>�()�T̬�
���D��48��WU[V��$DҞ����򅫘:�v`�ߠ��" 4�A�iy�~\qq��UŇ��E7J�j�q�mU�ՖztCg�`7�6�@>PQ����Z=�@㢟��kn��9�}j��Y1��`�a�K�����8C\�%aM"EB�����[���aOs���w��.]bX���tc��Ь���;�d5�&*#�vh�s��
��]�&��x1P�d� �O!�
�^�tm�.[��]kC�����F�������n�MIDe�i f��8X�Ǻ��v2h��8�J�{��h��N@�T�l����ҧ�����u˨��k*�W y��M��վ�L���=W�B0b���yWJ�{�/��z�{άJ\�ˆ�y�|�N���i�MCS:Ñ
N�Q�w�^�d�3,x��
��6>��H\WJ�#���q+%��uLE���f�D�@:���xN��X�u���y����{#B�Y�6���a�u�׸���X�)���ƛX��A�Q�#5�앍u��^�p��CWQ;oۜ.Lu��l����Jv�N�'�4�u���ɲ�V���R�ԭ!����U4�d衼w���m{�i�*CV��l��.�_lM��߬��$�5/�������y]d�\i���SȠq]${q�����`�Gpʫ��E_cQ[K�2�u�1�3e���zC+���4��
�����l�|�4H�0�Swk\l'��qQ�m���:\E����=L]L���A�W�؅�[����C/ ��7a���
�:��ƧyB�,zi޸����V�~���EH�_]�f�������N/"��a��ޤ��t�l��x��]����I��,�u���R<���ӏ���./o3.�y��g{N�C���X��m���͡L}���-9���	k�ku�y�����@�*��L�I��dc��f�W9.�>�p�I<f:i��V�J��f��*��՞U���u�{����n��ۥ��ш��4`iv� /�\
�C�_]�t�IX�0��u�@Vz�И��+�R��0뤀���� �p�BX�+��Նu� ��e�Jvـ+JE9������)ݳ"��EI"8ҽ&�q���q=OSTA�h8�0�_AY\~���[�@��y�_D�Ӹ��/X�����\�{�3���>����ȶ{M'W���ڕ�b��?TsT�y�r��L�V&�`턣J�%m7҄p6�02w������L�b�b3.��{ld6���
�z��[<;:-KYi`��,=|S(���}�����ͨ9ye��"�-�`������M�&�/k�^*��1��8���d�#7���_�9f�nX���5,^oD���k�+q�w�������o���)�zb���eo;�;)`�.��@axx��k���e9x�M�w{�]�ަ������n}z�
�k!�2�#��q܈J�w%Z�(�ʝ+;i�v�s�#/E�ͮ�����?�P���7R�/�0��T���φK��dC��4�s�*��Ms3�&�H���˷E�ߵ:�}Y\�#��WL�b��D�����L��q�;�B�����{�k�E��T��zfn.�ݽu��1�}��m˖k�7�F��]�mګ����eb\�����yu=�h�;�tY�5�)����s����J4)�'D ��Z��#�Pb/�-�+�r�������DT��65#�gvU�+���h���]���,$�R;����k�]P��W�%s�p�J�q�.�G:���[��V�<�w�r���Y|@6LJ:	;S(=��SK��vA�lV��9�wD~�{�p4��hO%OO}�C/�i��y�2m��������m�'�v���EF���T��06����&r"����c��}�F�1��~�P�+�RQ�W[4���&1i;m�J$
@��ZH�[��(E}�������e�븛���t���2�y�*�q�Ք~v`31�@]Bt���]F�Ƈ�&�PF����{x
^tE���i*
���q�uu�<\�vk"�4(xV}P}�o���=�V�������i��-Zf�+{o���ؖg������L�ΐ/ :`�*��Z�%���.����v���(��u�,+T��(�M5�U#��_r�d�&���xPˎ��L��u3k�:ze�rz���_*~u�1���g�����Nՙn�0h�V^��b�YqL@\t���53n���ۻgD�_M�V̝C)���8�tu/���[��t�h�:Uh<��/���ݢ������oWgP1����ݠ;�jo�k���G{:k��e=�5�(A�}���+�k���N����O%@��N��fl�q�;yl$�F��ӶX����.)��⭉�Fδ���A��s����q�~_�p1���%e�6���3��1�1 l���i
���
�?(P�Cp��O�Ď���'"�{'��S�~�D�Y53�l���6��_T��Jd��I1|��zy�A�ܚ�!��gi��s�w�e׹d��Z4��:.R]dU����U{���l�<�ɢՖ�@��	Ӥ�%)����c����;�+:nN���LLA<@�w�榏�t�~�V�8���ؓ+�j�	����] B�М�V|��܌=9�E-� �	�c*�u��W`8D OJV�)s��(�N��\9B�`#�	��������:�uכt��E�|��0�'*�&�$QS��u�qIg	���SF1�&nk��>��2dRrޥa�T�Ƣ%�F���P'�i6O2���V'�H�δu�Z�����3��)#M�m����U�^��tN�j�H���=~�M�z��7Y"o(��GuM#v�_l�j��/���ވ�d`���]�Z�B�@�q����� �6u�}5�5�NQ ���G!V�]D�������짎�.��{+�Ȼ���{u`�z�#�z��'�ƕ
��4�A�iy�'��\�L�&�����ی�+�{���.tCg�`7�nh��b�O֏j�@�:+l7��7�r��9��߯���-�]n��s!�.m��*�+�SH�Q
��Ls;�[HL�T��O/���70Ċ�,1�V��R��Rc�th�s��
��K�$�-�06-oS]o	;�%给%z�b��=:^�V%R��.A������ZN�2�@Ij�mȡ�!�=;ۍ�zchV��t-V���f���r�>ϻ���r��ʩ�Pn����ކ����
z��`�i��;7�J�{#B��&����#1Wm;~�*�UwJ�)���ݬ�h�x���??n��8't�J���5u��|:Lu��lӡ�W����xF�M���Vl�t+ݏ�u��p�٘���WM&Y;���ڿ�ڭ��Q��N%��b�Җ_WЖ�N�y7�q8��SX�j�K�-��y+��dA�1�mޣ(!J�*<�NX��;����EX�ǯ���}ۑ�$򬳏kCtL���b^��P���:�k��l1T/�%��vf�I:gs�:��aI�h���L���;�kunH�P$�������>W&���Ty�U�� l�7�����9�Y2���\ �h-��N����t_�2�T렊�3A����+:B-�P�4���UmM*��5{ܮƣ�*Q�0h�"JOi�4�)U][��&�o'�$��k������'ۇ�Z;DG�㤞eW��])��M��c�ƻ���͑,é��OF\�/R��������Oޡ$�� �!�`�㷶��s擲-mY��������Q.&X�6\���#i�t�ћ�L�#�<Hc���53�7GOtg%7[�̡|j1up�� V��&,BJbrUR28���)���;����اoR]dE�$L�]4/�Se��XAq�7�]l!��e�"�+����%4�1C!di��$6�%��정w@��:G�3�i;���;�C�=G�j�.F�B0
�3�b��ōQ�;Q`O��<Q;@�XC���s�b�Fe�[�m��m�w9R��u�㪪���@b�����a��uT�6�}�m��ﵰ~g:p��x����`MS�0ʛX�kq`\��|��R��Q�pCs��]�f��P�S;�e�M�u�l�:���{�'���C^�iNP�*۫���rau�S���h|���,P���
̍��v�k��#�pi�b�Gt+8&Xg'E�ܮ�z4�K-V�V)��͉����j�]��A�t����ҵ�
��e#n۱+O�+��+B���g�gț&t����^.q��=Z�����g����Oz��&�5X�1�(�#~c���ja�hi]�h�EO{jY�%�n-m`�D���L
�7�c>uN�7�6���q�(��"ȥ�3��I�=HU�ZUhB�ON'fS\��Y�o>em4����ٖ]�m�
�͆r������;o�G��\/���YD��. ���uH	w�j���F_9�f��O@k%�Z��}HG\���)��W]H�Qa'G|]��H״�:��<�����9l�]5�t�[R���it�柘Yq���1�n�$��$�D��2���Ԃ�d��}N9�����ޜ�h.4&�%o�s��㑧�6��\!�g�����u4'�4\���vn..m�:4:�����E7_��c~k]�w��*�3�T��!-13���]X�EK���t�l7�����EA<�r8����Q�xcN�����L��gyz��7�-:6�V9,M���ō�762B�+$�5J���^���篣���j��vqǓ�;�+{2�v-Jkb�P9���'�q�z,L�j�b_���1 �#r�'B,Bo2��<k%�AD�c]:��W!��%�zE��[�6{5-�g��W�m���H���hRfJYVZBu�5�b�v�P��\�L2=�,:��u�aZ#��հ�U:��*�s�ND*>O� ��PM���%%�&>�����R�v��0~���eY��$�_)1�u�us�r#�Z�8�P� �Q�����{ۻ�����.Sl-�ƌ���a�,q^g�I�0��.Ɖ|��Nmb��|�-�έK^%�t��WԅF��Q�G~G������}���*=�r�x�>SO`�)�w��)]<�spv(�A����U��f���S#Yr`e��32>%r㌫&4��v��ګ�j�,;�&�}��\�P뷃QSY���ZR�����jj=3N�IZ�9` ���f�n���t�`��OU�|�s������Z*_.x�	���fF+�h;9i��wo�O���K�IMS�_����8���h6ѹ�����d��W}���fQј�8��u|!×u�c;� $��V>�7N.��,d�i�o�5�iwq�;/l�vA�:�&�B�ٖ�=��tiV�b��Z��f`�k���>�Ѣ't�vն���"��WkG�WM"��n�M��.�]�0�%����/c���͙0�l1Y�3au�JaEx��wnER�1�N�� z���E1��F�f㫽��u��}�uv�U�e�[��=��tE_'�G1�]�	���Ed}�k;4 C�����pڄ��-�{QN��e��l`��	�G��\�
h��j�=5Qq-��^i�p�\��f)1e
ڄTV�w��VY��U�ɹ@)��-���JSGogE�-1���,#B�[\�W`pXN�\\�;�mEg";O�I�~��V#>��G�+'Ƴ�g-�Kz�:^:"�@4w��1�^.�Ji�-���>)�G���}�tf^�)��m3�b*���ٻc�>��e/�9R�ec+��h�wJ�=�����Ʌ�^]Q(&�Μ�NݚM�/��-�G��n���t�7x��hō��Ye��Cc�.1a�MN��3�lO9
e]x��^�n�a�mӫ�ů,5RT}���A#�Ȇs=����:���+����ͪu���A�m����_,�[f<]��.�38Vb��6*>f9���p���3�շ����S\U0�X���6��A�ǩ�����Kqn3Ons��v[(=W�&_P]Bp�u���k�.���xe�.fv.�|��z`C.�鎜���5�u���;�Ե#����3J��F��������쵍��U$��|��%n
1��R{ۈ�9��[�Wr�u�k^A�0�����Ҁڵ:3�<�W;�B�ӣ��GŻ�)���HiQ/�!S�fFeU���dH�Tf\�OID��@�3D�L�4OP�'H�32])"=E��sP<�4L\�H�4�L�K,�RZ	L���-��	(У-�UL��Y���"��E	H�2$�2�0�JJ-0�%6����/L�TP��Z�ʭ�5LT�'#M�a�D����T2��҃(�pȴ�Ҕ�%�ȴR��J�B�&�K�vG�DH�E+�*��V�Ja��Yk��b"&FZD��᪒��Y���G��iiaG�&h�iJ��+����Y��^��.n��z�]ZJ�"�V�W��XZQ���*��Rz���zn�eeU"I��e���릘*Fz�^R�ei������TZ*%���T�Q�j)D��e&�y���B�ҫ�5�O%-O(��4Im��1]P���ѽ|~^{��}��ُq���lWnR�4ȩj�ו�
U�y�gH<h�]��k5�
nA �
Í���ڢ�eĭ%���7���U��Ϲ�_3�H,���3W�B�
�M�-)<���(.�E�μC5F�ZZAq�9�<�eCY�Z��+�O��a ���s}�[% m)���W�1��>�����u���9�xx�;5�}�so����%��MUE&P������He�d���z����AfWPn��ؠ`��'yAm&�.�3F;f�e<�)i5�gS�-6�Y��^�
��)�1����������uNokӫ�D���b=�Q�E��d�ɖq����>�$��d���Wl
I�))��\��S-�I:���2�)'S�l�]a�ePSG´TX+�U��g$�^��6��}�{�׋e��-������m��s���H*���a
`rw��(�B�ܲ[���<�aL)8���Y2�(R3\���Iii-��a �������̘@�Pø��w}�+�ڷ}���|�f�)&_jc�'�j�s1d�>r��Vj}u"�$��7�b|�H,���`�=B��]Ȣ��[=���R,�a�=�Xi�&�����~�h��"$@6A0(���_���Jd�Px�8���-Y�% u7,���6ϙ)1�!�l���l��I�)�&��௨�3̕�{9���ώ�ؓ5D�lRh>��� ��Uޏm�="�y���^�C6J����i�	4���)�Kai�x�$gXb�ߘ|��Ѭф���%������J��!�*e'P�S%p���X
O!I��1'���D]"j佁ѡnV�{3/�ϰ{�b9'��,��,�2�I8�K��1�ʰg�M&P�J�G(0�!l�6��H,�e�G��2�U���Ha'�RK���Z[ėUHCG�G�DLǽ��ҭu�n?]_�}����!�nɅ�IԴ��ظ��Y8�׽��L�q(M{��,�%0�����dٚ-'�m���k�O�feцm2�Y�a<�a��[�]�
�bDH�9�=�O:��� ��i}9���ԋ)�t]��̖�ɞz��T��'�}zH*�d�Q�bÈRA�f��+:�L����M2a�m��5d�m���)��q
|����r��4����#7�(�i�b��,ѺAS+}}�E������ĭ̽X�];H������:a��f���wMD
�Vz�����S��]�V����Ӷ��/��^���}�ȧ��8��zΩ�rJ]��f�c���᫐@Ke.�ҳ$���$���FY������I׉����l�&j�m�fO�ra ��C��,�%]@��锝aiğ%�����<�ai��ڳ�i ��v�.Xq`u��RE��%�#�����*7LNLǲ��&��w��A}L�v�Y�*�����l�v�_ظIoo<�0�R`�;�:�d��:��4��
d�0s�q�u�ף��2�o�v�z������E��Pe
I�)�^薅��C2�a�L)�%]�x�i-
L�I���Ka���Rי4g���8�HJ����S4�L߻s�3ꓬ��k��}�E�z��q#�`�14=��I��N��L�i ���Pi0��!i3T
�N3�	�"�L]u�L�d��4]��T��'�һs)�d����e �k/�q*k�����^o�ǿ���>����._Ze6��ٶ=�2��S�KK���C	-
~L��R�D)�fgh1��ަ3�-��UD�lU��1�;��l�tMU����I�[�v����/.�{�v�D} |�1�H�%�"#)���L�a�-����n��/�̗��0ɖ|�WF�z�ɤ�B�I~�cTB�Z}�0�d��D)�r��a-'^8e%0YL���'��k�Ư�^��o޾��|�x�[���V���>I_W�z�a�C̴4n�����ϐ�ys,�2��9�^q
I�)4_�j��--�|ۆP>JaI�Za�%��+�I��6��cn�eS��0#my%�D!@��#���S,���3�Y����a��ʨy
�I�-���&u�m&��b�S<���1L2�%�3���<�anP�5�Y0����Ί�̤T�o������WyS�rM����>c�}"��H��0�]I|�f��0�Y�2UK�HZAɎ��&U�2S51P�a<��l�j_�
I�)�&w�`�AI�)��}�4���h��bJ���	=:���_GK�ќ����z�Ch��L}BD{�hG���C���0�WA�Kg��Zm�ʯ�	�N0�b͡�- �Cy&�|���5p�h)"�8��r� y)�d��\�&y
c�c�s��f,���E�����Ί�*3����Z[;c3ٙ�z���:�W��k�E��pv����-�A�����^������^��h����r(Y�ۺ5��/f��E�E��n;}��9�M<M�΁�DG`�{��[W7�3�1s�	õֲ������u�>�>�o*��}����г��I���}a�2�Hg�i4�a��3�-'R����֨�3�y���6��)�u��3,�:��j�s
��)'�U}To�/ڒ�ڣ�2�%kC��h��DH�j�c�@u)��c����ZKM��C�)}Ru/����C)�ת&��JI��X�l�e��Fy
���Z����4��<�>�γ�Ɯ޺[����Yֱz���e8a�e-���/�%���Z}�XVE1�{P�A�I�s�L���[�KKۛ!L�jK���:��
�^��;�q@�P�2X�|o�1�"G�h����F�1c������^�����=%$�
t�Ҩ�aX
O�����K��S��l����sx�a�d��uѻ�"�U�xI��[:�WF;@a�N���;y�Ĵ�ϓi�T�|�P����ﵼ:�����v���YF��K=C��>�>�?G��z�L�CJf�)WSl���S��K�Sf�C)L�o�M����I׻�cL)���޸)����g�D��O%��cx�=�����Vk�[ڽ�^�ُ���D1$��Դ��v���a�B�e�+
B�|���'P�]�xɔ�3	l-8��o7yB��J^Ԛ3���M!I���ؓɦm��Y�_���[��o��}�s>��>e3l���2���T�M{ץ`)<Ͷ빸i�S:�U8al�['YL�KaoYM�dQM�N!i���l�:�">�>��V+������v����yk��{�s���U+:�1�HZM�ꎲZ����e����m����L���'�a�Ұ��AnY-/�$�a��URm�a3���J�
�&��� }���!���$�Z���I��[8��|βB���O��`�M$a4c�)8���0��Jx�h_��b�)"�2�ؓHJg��Ϭ3��d��N���*��ʂ��2m�Pz�{=�֯�3�����ǉ�S%&��Q�X,RL�ZN�R�u�+��`RO'����	�Q
g���P�KH>���6�gY�->�,+��=��H8�m53�4�|�hJ�]k��װh�]d�>�0Z	�Z��K��6����u���t�+�[	p���V����H��hm�2��qK����N��]���3� �����8�]�u�5���,k�΀ L��F�:���a��y���L2� ������#�m�s����aķ�Kg�n�P���ꂞKIhR�Q~��q0̲S������̦|򨖓�WjNK�1-X
M����'���
N���N�al�[����0�[z�xn��U�ck���s���N$dQ����q$T��-�g�$��,��������- �1vm��D��椾��KVa���@�Ry�}��d��B���bL� � �=M�ʺ�[���{}�����2Z_�'�w0�2UT�z���H,�%U;A�,R
���I۠�m�K��u>az�g�|�H,Ɏ��M��-��j��J~a���Y��1G�%�o�׊c�eGO�gg�W���6��N�:��KI�_{l�J�RC��$��ɶ�_N���2�I�h�?6�`���*a'���q�(�P��G�J�a�nծÁ�?t�������̜<���1�r�/Uik����
��{$��ҹTk´#��Rw˻�uggE͗���|�\'���
L���3��^B��X�OT�4!�i���dR�㨦c������2Op�c\���ɹ?�}�u 7�aC�w)��M�U�1��4fAܘr�j�;|ܽ5�k��@]���U
����*����\�Ӂ�ޟ��آu�Da�����љ���ℋ���kL��>+��T|����]_*+k|++|����N�� �5�|�*���l���o�O�ݱ����NH��E{O���n��(��<���cڛ	��A��b��<��}�|R�5�8��~
��u)�Wq��f-�[�f�1��{{q�035��տu�S�kVk�r�`�E���{��R����Y�K�h9+��f��̀
B2��r���}�F�=�ն��d���w#���>��1�6a�J�e�P(��tt� ܝ�;ԜOdr@8�kZ��Q�N�����Bi%o�2z\i���u��e���(�����ߤ�f1
乨@Xd�!������}M�Ơ�x`�k]�w��*��?`��-2.����_{��?W����5��@S ��EA<�s>(F'<0w��q�ߋζHU�kZ��_��~�������2�~|hqU�P�uAa4�o��Q�.8�%q���):%}������ٽ�.ޝ�J���?�tɋ���ɨmցr��M�,����ƾ;$OҶ�����M���b����{���&��ZUM&�x0�B��T���S?T@!3G��`Z}J�N��j�5:�<*O#�_��q��O��mT���4y7@s�(L�P�������x�m�������^ �T�Y�����Z���e���Uq��~ri��	�م-��\]�[������J����U���{	�:Lln�L�o:}��.t�����̆�|�g`Zj�v��{J�ѱVe�2��P���e��ǳZ��f�d{[�I��ѫZk�����{ըt7��M�7Ǜ��b�귊�β���I�A)�i+Z�z����6V���^�PIq�m���+�R�5NwO�K���K9�"���������w��y��:c���(a�9�����
L=0�o�δ �si��֖��>x#Q����{'����ېz,���]tt�wA�gU�&e2y`�p��@�ޛ��{})$ n��j�Cd㟵r��s�R���J�V�6|N���Y���((��wB�7�����f#Q�ٕY,�k�r�}�<���<#v��ţ�&"MG8�2<�f�N��{y��JJio�J{�N�}��<�G��{ų��n��b���	�X���9��U��m:\WI���P�*&z�]mӕ9jb���;c�p�Ȃ�Gr���*�L؆nGJ/5<W��:k��%$��;����ҵ�>]�K������eѫz:q�]�i��l�1��m۸y�_�zL%*�n	�Vg�W�}4!;�uu����5��^Ĺ͸�pU��	�%�,9(JS%MG1��J�NܘsB�����y*ʽ;���j1q��'I�l�9Xn��V{U�� �Spt�8K��ܗ�����.���j�yО�7b�h��d��bfc} >Z<2V�<)-���������|���3:nS�	�ՠ�T����D��۸�Y�z��N4 a���j�V9S5��˜��]�k�NΜ�=8��\E�}Gl�]��1O�U}_T�Y������J�
���d�F�4�1����9�i���s�r|H�J�ʸj�Lt�{ݦfae�`��0��c��}�+M����
��4�Ѹnb5�C�T:V��~'5�g<��U�����uе�0}4��E٭8�޻�I����!���b�C&^~�m�KՖ�/��UY��:��!����{G]yϤ>�s�ff@�����۶v�u�	~]���K{��x��Lr��4�l�
vx�`����P�%�1���ˆ�eF���R*�kw9ѣ�i�/���c�zM�!��O\��*":��l�΀�y7�Ôcۛ�^1�҉�'O�Ī���>�SI�N��6���j����1��
6��6J�ytL��Ib6q��Bg������1�WX���U���>}�*'��۠8P��Y���o9ĕƽV`<_¸V뢸F
��4�)��8��4����*1ä"p7���v�Vq��[|��}��U��{c��]�.,P>�+_	M-�)�<+�����(s�>K�jĮi	�{��[ME��e��5Mx��&���VFn���]�e�|�]�"��Yvh�'Z]%"#yK�Σha#��)�h�^���c���D��v�YT�(��;��ћ�VT�|4�$��g9r�|��ݷ��6�ـcꅌ}O�U}_|��ǉ]�=����&�r��処�GE��<IUc��є�P?1A��N�D�:���[�wK��q��T��9��y����z��\����g��u��+ce��*n��F�'V�����2�q��2b�R-ӫFmL�>�Ȳ��[g���椠	(�63����xE�8.5��vD�m��&��Y1cbu���Ak���x�������];�dY%Z��ህH�jb|�W��+å��8���[VY��)7�L�k�,Vӭ�o��ԫu�R�\W��&����4�MQ\bs�ѩ\� �l����OKo�]���Z��N 9`k�",	N�&8�8�:̣�t�v��uLׅ����犻&+��2l����=!���	��7
NXZE����O�,����i�6�jy�?(�����)��6���Z;	Lh��ʅq���@t_�(�+��	Z}i\�5�Z��z_�"�CC��I�z7�?�O�Su�'��:z;�3�O~�vey�3ޭ�牡��1�������vp[Æk `ѿl}���Lh�@�'b�:�#%`�rTU�u:[�
R��g僔ph��k��,;�D�cT�9�e���c,���vs�
�N�2�(�-�S��\4���5�q׍uK��뚏*�n�ՙ�mbx����?�������C{��ݙ
?�ä�TA����䟳�<9yԀ���c!�;�D��/CG���ɩ�ggx��s��Nb�Wih��˯A֡Vo�k��� ���BxyxBC°��5�Y1�~�{<"�}�&w��p���,���bN�*,O��@$�`��t3\]��9m�D�B�W+��S�´�h�����"�N���*������BwR�Xc��:ӉUB�.��0��BF�LvB��`�i}�'l���vgD%c����ݨWS:~��f1�dN$���r|sO�m<�6�9WxT��s}��	��#&��W8�d8Oİ$t�5 �����}M�ƾ-�-�v�؎r4�;�\l��ng^�FT�6������1b��]�@p!i#I�Ә:P���2[W�R�ؑ7Gx�N�V�N"���\N������k��7F����A�`󝢨Ƈ�jJ�&A�]h,�ِ�V��uA8��U����1a�M���q:`���Ǝ����ZM�g*�mA]�}ڥ1@͋��2ŏ��u;D������K�Zbg9
��7��˚ܾ��c��I�HvrIWWU��b,��)^�Z:�J�vv�b��5%k"������q�k�j'�:�R��q��w�e�kzĈ5�WB�G�G�F:�!U�NU����W�ј��*�%7<A� h���5��/T�;��G)�VJ�Ƃ��+"Fw�ϽCf���w�ә��z����Z�����������$�׭��k7���7sݪ�K�qX�8Aͭ��YLU��ӽWP���1���&����RG*�AmP3�\�x�f����g�
��EtW����yy;�o:�^m�����TEcޱ��]�Nk9����+��ַꈫ6b[� ��vU��q�r��Վ
�4�뻇
B1�J���_,���U�3�A����jhw�n?��#BJ�^'2]e�s���d9���\�ٚ�u�i8� LZJȾ�P�,��g�U�/涸g�Y<.}Iu���oZyI�wu�����-����Zn��$n6e�W�,�j9�e�����{%�f�x�^Ҙp;#��yzG��.�&{���&�Na/�.�R���j��?uFH�G����ec�v��h�%���5��}%f�,Q��x�8�(!zxdV�9SHă����������R�~a���2Q[&�u��i�{���X�2QJ�3�
�]ٵ�F������[[PLh�|�@��kA��1q��v=`�:�
B�F���H�u������-=��u�6���38w&��*ʸ�g��n�]�%���V+r./��-X3_}������<��B�Ɂ���N��f��Wk��%J�
� �8ǽ��-��,l�!��+�vGû,��W��-�]�v�XOR֩n=mp�ܚ;|�LO�9��ן]/��CdQk��9��V:�qW3�^=�;�+�.��R�m�
E]n�hU����9ER��OWu��O4�_j�9�pa�b%��ø�n���4b	�c]��QkD�����΁+��	O�Ǝ��bݒ�
&�i��Vm�q<v��&S┫�Y�P�j��*�;���n���3�]�2�ik����<H����D5����QtDY�����ՙ��֘����`u,Ui��T*��U�P�VS�=�)�-��u���/x-�L|8����4��Ek �;>y+��h�.S$�]�6�U�:��
͒;C�.y^<#:��߄F��Gh]-Eiw��i�8��i���b�K';��r��]	��}�p@%�-s��2���ӹ�*�9ŮR2S���4=ttsвe�c7ik�Sv̢��^8����ڂ�7�^oZ;�������F1A�j�떳xR9N�g�I�x���k��j�>W@RR$am\��V 4ż4����+�-��k]�Qf.B:7.�Z,-4m��g�VAf3�M�z�ip��Uˈ��};֮�i�E�3su ���
����Җ����ᵗaMn���P9ی]�N�N3@�KB�x��v洰���9X�T�:{�a�V��]�݀%���+V[��0���Xyp�T�HR��.��Z4�o[�F�9M,P���ׅ3d�B��Mؐ�ѳ�@gd����u6v�$R���IAB&*��$-��t�5��N�i�sW� h�L,�O�Č�o}3zl��*����yk�o�}��P�+�����p�m���vh�]d
k:��o8��A���x�2y�׹�+�����K��d)��*嚰�^b�8q�T�*�Gz�nղPt;�k����_w'V%��Eh��&��Q��o�gi<��)��Km$�7��ݡ�޺�������pvn�� �bի\�x�`e�܋r�1.�n;��������[�]q����Vpq���"[�JJ�M��wB����T�F�Z}�Z��`jD(ᔕ�v�Q��u#v�`�+b��`��P�4�,�N�+
���oo9[��F���s���k�N���=�A|�륫��k�J�.�Ơ��Ė�����˱&�D_��y�gMM���@�NKe3N�x��Ў��Sz�f��c�h^�j��6�g%�;;J���S��o�c��Gm��;)��'�R$�x�>z<޽�}�)QZ�I�a�X�����nD���i^��*��^�a��k�QZ*j�UeZ����P�;n�N��*�2Xm3]�7#3���2�,"�2����="�LнK(�%�!0�Yً��a�YjD���$���e����Y"�hyE竇l��������QG��Ji��Xd��y�aEBU��aZ^y�䉚����iRA��H^�.�Z*jD�Z��h��RL��M�ʂ�s����ĉ�"��fZ�iZ�&E��"����dQa(F�+��&�&T&�Z���UTjJy�a���IRI���4C�$L¢�=5O0�Ip���C-52C�J��2��	r#E�-OT�BL�P��J�,��������LU3q4�*�$k �i"��.��R�镨��f�*�����RVXY��ed�a�e�7F����{L�����N��V����<�P5õKT1���0���ei�k�������]�sp���O��?�U}_U��}G�w���L�n<>�(Bi'��`�E0��T�{������}`��w�737�w{��r��f1��=nc��Pݻ���C�ޓ0��v�Ó�6�����{�H��ѥ��U����� �_�N�q6�`�����$yh q��U��o�����݉^K�9)����y�	��\k�I�G ����9X�u�B�%��.=#'p�3��+o��5� �g�T��d|6S7�������c�0���K�6 �p=K���vJ��Dmv�u,d��|R�����^U���xm�uz����C��CF�V��=�����s�JW���AK�5�UTTr��z0p�Y�ڲ��D���J���3:��h7XC\��=���iݮ:�(<<����&���~��x��T�:�b@Ýu�b��Wu�A�D�+�3�7C��k��o7�S��1��1����ЧVx���dn�#�v[����"�Es�8�yخ�$�b�H�V��C�k�1�׺:Y+�̽֨���_��Y; �KHi�Q�k�+
��W��Hf^�4�2�TP���請/�7��}�k��r�}� àګ�����ͪu�w�����G0�wTTc"t�N���X6d���U��7�Ow�s6̾4�";;����G|��;;���j��R��K�D}��������>�҂����qS-��F��L_5p�T�e��(j=m�����1s���CU���2���q�a��=�X-���yMs�b\`ʧ��;{{�25�R�ʽ[���E{6g�J���xV�+�`�<'�/��A�f�Z|Y���oaHѶe˵�.�u���O�v_�fY���9X��� ��[�S,xW
�Oo�&�uVX���J�oJW�#\L!��:m�=*jx.%G�*�3>0�v��e6�r�t���$߽�#��?M�����;�3c��{�#[����R� ��՜�Qّ3
m�:��p"��>��}I����;��\��"�#^:�{�ѕ���z��*�2�}z��E�$p��|
g�\�b�����m��&��r�`����C�.02;�y��~�d�� ; �r��H#�M���q�XW�\~ڈ���w3Az�ȫ�k����8_�ŲU���*���)�y����i�8<�g��^����c��aXv#׸S�JQd�����ҡ�)���sZZ�ʔŖ�[�7F֑��\��ң"gbx^fNs��'\�#Hk��-D�u;�=ہd-'b�g,��L�=PP��qwfs�Q���!�z��~6���p첖nL�EJ�)���V>��W�UW�����{���?F��rT�y�\�Bu?qD�!a�����]Xz�v�q]7"��Mn���6����Utc��������&:Y=P�J�#^8�#y�"ԊͽW[�L�@����Rmm��k�M���n�A������蔍�Խ���L����Υ�_���h�ϻ~ò�L��&w�{����!O����hJ�5�itZ�� �ks�э��P]�&�����c�T���<9q�H
�k!�uN�*ڡ�[;pW_���H�=�G.Ͷ��z����h	U�
��
f�����*� P��dk�����yz�M�)���8�M�ϩ�٦���q��<h2R�?X���
����ժ�s&�h	OnE��K:���h�xS$Tc���9b4�І���֐̋	8]#�4��D���m�O9#6����|~��J�9qt�柘X���
*c�e�Yd�(�^iWGO96����I�P�1��Q�kU�R�U����_��H}-mrf�Q���	����C���Vv�6�O�ޖoYc1p�n�.��}�hL��{���|g�W�A�Ѯu�+�:a#k4�z��\.�iҬ���U�۲�^r����'L-yڱ�!J����-�ŵ�
�6����>���Nf��HW�U}�P+������]��'�P���ZS���f[����x`���:���kp����pG�k�@,���p�nM�����(��� ��{���놈��"j֥!!qN]��u�kk��c�e��n�I�����2�~u\hqUZE�8MO���1���ʴ'w����^��:>{��a'�pF�M�C>-�&����N��h�ҭ?v�q(���X��k�u�׋�P��."�3���c�#Q�L9)��S�:`�&R�����n.�ۧw�*��w��h�,���%��{zW���mLH�̚7�n���ȺU��B����ur\����$���=5'�1�mm��˭�9V�����r������'b�j�P{��6����u�@��&C��P��hB*�U���罬
5M�_�<�W��羛����k�M�Ss.
�/gַ�Vl��@����P7f�5^����k;k-�r��-��kFp�v�p�FY�o�>s�����ډܲfx��+���گR���ڗt����e�)�Ft��h����}Xs�kA!����4�`����p�p����X�⹘l�fe�ӝ�%��3��f�nbw�*ԀMH��{t�|H�m���Ď�V�����Ҝ:��ٻ�J�\�Y�DqS��&oP���.�Q�_h�&s���/�f�4ա�z�*]��vǢ"#菛�4�eI�ؑ虝d��H��|Ց}N��q�ںnU��ѵz�tω�k5.V�L�����ԕ���FJ�G~�����ˀ�	e��=�����޸}��Sƺ�Ҹ��6�CC�*5��Y+�Ю$���	�
�*e���*�}�~�
P; �a�岫#�x�Ew������Ծ~�G�������W �
��עS���\�Tbv���T��s Y�˴GN�����SX��(Bi'��$�@��ô=�:I؟k{�x�y��j�ӓ���ь�}'\9�t�=�#��Vj�����s�Z���y�?r�Q��P�"���^����5��d���v�M�=�#���*k� `�����8�����Z�`��Y�Ǿ�ƾ��$p�����Vۭ�]`�*�쬳�yk���K��i"p=�/fɀ������)�L^�˭�L�a6�{y�{��F�'���}�{�O�"���J��v�^0�a��3�i��u!��d�.�a���2,
�ԇ3�K�����ns���t۽��-���au����~Y�X�n��VS��]2���z�[����JƠ��@W��EtQsq�+�$P���WF;���ë]�p:�wB�J5{k�Qb#��n�}Үg#��+c1{������*���-��e#G�ت��u+�Dޞ']_c�Ӫ]�0\D�xj�7&S��GJ�����ew�޻�p�L�r��_s���]ԃQk���v|a�����5oKX���g,�����+%���Sp��f��4�,R�ʘu�4)��m��W��}����\V�w{�xӦ��>�-U��3��q�}l@	�,B⺦'����L}�fvlL�q>I4���r�|yX�T�2�io��*�S}ҽ|�������j�㶶{k7!Fƞ���b������
��Y�ٹIp�A/���ض��Ӥ��5?F��P;9�Bj�Tnme=kb�h�i�ʹ�Q��6��wQ�.��(]L�T�W}�h4uH��B#BiO��]�*{��w��Uz=�HM4�m�2��Q��QZ�J������+��n��a�A�(��˱�6w*�s�)ތ�\L!���['=2�ǣ���8�'�����o�[��I�5������<����~��(���~<9�9��c��{�#m����D�����x���j=p��1���/�72��ڥ��9�9�i�)7շCj������VH&]�5O���
f��O�}i��Yϓ��P�z�F�i�z6RdLGQ�w���]�}MY$\�:��f�zo��S%Ѥ���KJ�×��}D}�Ҥ�f�oSX �>����":�h.=�&�&�e��Ɇ;
d��ʹmV���'����ky��e�L�"b:��XJ�
g�\�.��)�f2	�)�����iڥ7������{��d{'��#�������y�кSe�a���},�+f��v�ʴ���Xg���A1h�a��0�;�8�#��U�Ga�G�t�i�k�{���	�ď�*d.���Ӵ9�u�b�g��Q�S%�,rP�u<Q;@�Xl���᪩F��x:�J��U�.�1�Q�Eo=�3��]�Rr������OK'�,�����q�w��&}��|��"�>�w*��-X��N�� :,e#m=�	�m�#NL򲪐�w��;�(F��ܱч�t�?lހ@��;��g��ٕ�(�=����=��|�1he��ɴ;�-1�Q���jٮ�6:ڶ~t��r���Ʋ�סe�C�*J�D������b�j��m�U�g
--�:��C+�.�����>k��ឱO.��&pU��1N�c���s��R,�������T�}q�|k��%��5��f�,A�87Y�*s'p����ڧC��Mwi��G1�b�{I����aNAc��_׹��S�Gi�R�N)�NXm��N��[�������"�bk)�����V�E�*I���l���}�m=��3Ǿ��J��bI�)���G��}����w:�;K�Π5p�E��1�n{~�LG\D���dB���ne�q���e
��%u=+�lh3=_W�c���@,�%w����u��^���?������q�4���S�S�5y���K��XuC���~��v`q�Ƅ��+|s��_�4���kr��Ž�W.B�sYK60?�g�
:���I@H��jiO�]T��������n�1�5�t��u��=g�*%�!
�T�k�� oTA��I��j��P-:}4o�;u
���+�����W��{(js�OD=w��3�B48�"�k���K|���預w*Y��sN)��T��F���6�/�w���(d�EKnp�\K0Y�.=];��u�@�X�%��nl�g%QtW����R5p�C�I��^|0�B������ڱ�T}Y!;��oqėޠE�g��}�ß5�8��]�{���mTH��O2h�ɺ��Mٶ`�1XE��7_�,�c���i
y�(o�ڋ����G]ի<F�.�����]�X�[��)'_'�ЂU�I𲫻^��!�:X;/%KMq'^�+�&I�.�
]���g�V��Ue�6�l�$s��E�([�^�뾢��ԫ7���>���>����[��z�w�ٌ$��3�0���{����Ʌ�z��jN�ᕸ����/��OU��/��r\	ԝ��}eY�hUB*�U��0]=��a��FLы�W��m����߹슕t��
?/gֶ�f�Kq��Ϻ�!]���]?��=���;�޾ Tn*�-gA�t��g����9�~ߑ;�ML��\�7Nuzߧ�=3n�>N��|t�2�� 0��VE�:���?j�mW�kk�q�1�7z]���Q3��K���V\��uH���ѽ�p��&��e���NxF��Sa���p���%�MQ鈓H�D�릗�T���4����>�C���~���FW��7w�o�R����gO�W*�_x�������>��Z�J���r|i�]���ʵv�y/yun����S�X�&�b��~��BCI=�P�=Ċ����kvX�!jMm�픇t�uͭ캃��s���,`���1�>����1��n�C�rY����5�jE�{�o�;OnՓ%�%�uF�ᴂچ��6���ij���jlP�|,WP&|Ȁ�l$�ʹ=h�c/Ҍ�g���b������N:�+��NA��ný����{Y�[����`]��2����|��G��z��P�U��=kD7��]�w�:s�3��}U��Oz�#e'����'�N3ِ}���nㅗt���'\8�{0FW��Bj�S��j��'����{܀ׅP��xt����Q��ܜ�Qs�9r�m�bC�@������ό��D����+��& ?@l���+N�������W.�E3!�F�^n��P'4�v9��t���`?�?9�8n�U��]�IL1"�1��+M�:��Rxsr�tp�j�ҫ|q	����p��kBb�#e�D���:ů��>��j�-r��]�bET�0��H#�u��\&�� �S<��$���b']ԃ_d�v0�t��qJ�����/�7��뮊��4X��c����F��9/��(uTȋ�(��gaoQ��MQ4�n��Σ�%#�A���8�s+i�zMs�!��]D���np�l�?q����5�{�S{Dt<5��}<�yZXq��'���TO��\<�SI�LH�t��;qZɧsYq���N��z�^i�*CVo#f�\.��e%�lO��=���;�U�W>{9ڵa�<��E�.f>K���f�����)�%�f��S��ka�{����e#C�;�V>�B�X墇�][�Eքn�l�� KV6l:��N��;�IN�9�Q'�rEnZ,�ag'��g/u�֩l�7ǭ!����=�]K��f���kCpt���I�k'���Fw36E�� (ᔥ���8��G7ըkm�\�b&��\��ǎ'x�lx���'k�����f�A�ͼ�iu*Tr,ܬka��%�ج���f�
�A��T3����;�]]Ek=2�WP�;���]a�A[-!�+r�裠=g�6�<�/EP�ܮ�Kx6n�>v�s�� �E`)w�v�,W��Lɏw)ꔠ,*��.ӕ�"���=F6��6�Ӱb3�S�5l8�1�0
\��=s-ͭ��2{n�ڜ�l#�����^r��푲� �E��G;����� +���ܕc��_q�>��{�l�#�7'��$����t=�`7������+n��}l�����L|)^���(7�w����`���n�Gk��4�Q����VM�B*�SӚ�R`2�Y`╮��rtJT�H�s��ɦ�DEk:t�ù���
=׷ @��nFդn����J��s]|���̽Ӂj��B2|��M0�>��2'��4"�ؽ_wG9`��*����cy2ս���t���`+��S�r�x�:�r���za`_Y�E(�؂њh�mvU�'(�LЈ��|�y���лy�ڜY3�4Vs�����1�Z[�3l���ŵ����WGZ���׈:u�Z��t
Mf�\��;��'pF9��bB8�V�'���3:���O_k�!�E�gT�p�F��V�	KrL��V�W\��lu\;l�5�\6��z� +�c��k]�4��H�`U���҉mZ@ʹ�,.�N�0]c,�A�����ݽ޴����]Sw�_R�!Ή���-Ïp�_09`�&�[�b#�ڲ���}�ͅ���ݽ<C�Jd�v��&��'a�����n��ծ4`MuLxE]b/1lR�G�/9u��\��y���z�>�oبl��G��T�/H$ub�n�HѶ���K5٢�:W��i�U��M(�C��s9���.䫆�C��Y�%���G[�|^��9R�;sTީǫ��+c�qEI �KW�M�ǯ$N���f�.*��[��N=O0d�K����Ω�������Y��V�]�YC���� -�<�>�n��{p��L���3���Sz�{�v'`ێML.\�ONk&L6�0���{�sr�cg%�7ojK�ퟭ^�b�9����W��>�V[��RTce��ѠV�|�r��G�juc�c:��:β6�6R�:R�V��VY��
���.���,��$�t2s#@�44=CH�"<�7t�=���(a�if�Z�j�Db��U��^�aX�HxXVa�dJ�Eh��j�^$�V�b�RYh���g��*��@�b^!!R��:G��`����n�6(bA(���Sg.��o<�b�I
n���h�Hg��m&�u�]LT\��R$�t�S�,W!
,��		̵2+�S�v0�T;m4ȴ�̗Q-!(�,�,ȱT*DĲ�S-#I�խ����[XM��F�ˮ�n�f�$^_,���m�Ai�I��v�X�kmSj�UQ�e�a��^TJ!��GY�����OMSM0�P�C�v�h��b�C�MK��Y�g���b`�G�iWm�ec�'��Ӯé�*�yBNV�*(��g���O(�l�Z���<H�5%��q�4r��������7I�޻��ıԋ�ᏻ�"�F���7�q5˷u݀h�m`��i^�����F��>���w����\6��?�k��5�3[�F:4�:j1�e�t�$��;�!7��Ԟ��qpt�O��P�n[<�x>$V�P�*Q�� F��30g���B^L�O&�]��j��qthp����.�Kw�\B�c��_<<�낊%�x��7=�n��L��V������
�������}V���O2�_c���23����%�r���[��;���i*�v\D��1#��>��Rj�Ic��C��;NBrs��?8Ւ:Y���U�q]V��L�"z�Ā�)�l��8.5��vJvَ�����77)l���ʞ�Ƹ*9g�bUb��Ζ/7�W$x�$V��B�<�h\R�c/�2�j*�L��}�:�ojӨ����2j�8LZ%\_Cr��^Gh���l��F��_���*�4Ľ�a\kW!�g��\�2^@r�הDX�DON���Xc/�d���N5%dh�{LU�3|­-f�k�V��cUtn2��4����Yv~�3�Jg�-a�j�r�}t}����JU�������Sc<�v]E�T#fQW�!+U��Wr��e�q[!%<di�C��6ɇg�eؗkpeutI�S�$�o�5}PPj�*S����5e�wrb��8�.;�8�+F�-�:IZ�S�;{\ �oi bF���UU�UVL�U�{�j���͍�٭�N�qh��Lh�6!lrw|qs��E]=�%���^����^�&+�!b"�Լ=p�Zϸ��[7�/���1��
��]Zqx��n����gJ����I!�n�~�i��F�Lp���D������ܽ|��]({�G��nK���Nm��j���P5ݦ�U]�p�M[Xg�ƀ�eW�i�Vo�R��^��{.�vbO:������iZt����g��}�S����S��R��?X��35�I;�9����	�+���Pb06H��)��t�qs���[.����3m,��*w��jI$�#fv�";�}�Рj#�����ӣ����������;ݹ)K7I���I9���	�	9ih
�k��.?5����(,���9�2��-'UJ��Zkd�E�jǇ�
��48�3���liA����ҟ��S=M��j���:ad�1�ͅzwC\�|����[���߳�B�%����Pd�,�}9�h��`V�������7x:8R�(g�_�WԷΒ�KX0�Z�n��V��+�1,����l����ti��D��9�.i���N�T���$�]�'sO��#�;���k��ȫJ�:Ig<5��{�V���uD��YRŴ����,�F�9ņoq<�[�����{菣ﾪ��뢭��|�n���掠\{(nBu�K�Q8dK?/���v}a5��&f�8�������>�k�e�P֪�0$��?�t���b�%�8ļy 3���;���Xsd,�!�֖�6Y�"b[��tW��޿�Ԍ��%P��&�y� h�X���ݝ��֒������� �dq�୬qR��7�+��}[j�EB��M�Q�:2�Ф#e��9CoV�j� Z�4�*�U�V�㩛\)���Ω���]oץes�F����s�R�0�}0��=�G�W����6�����dK�C�4�v���
��.��<&��+ȳ��t�Brz�}�$'��/�>�Ξ��F���[\��f%��� �����Js�?���NR��F�q �`����q�1��:9z��M��k�˺�|Y9���Q�8��m\�w J��5Y�[��V	>�sQ S{��~u�N9�WKjtGC[\&���h�j2�bv�wtGQ�|���%�]��r\r�����ˀ��Y5�S/�����();��~I ��7$��ĕ�ºk8������\|<x����xӽ[�c��i"���;|��H�lj�V�8�����lɞ�mx�.�/�@�@`��yKvm�9�]SM��x��z��́��M�w�>[��!��9�����}�|�{E*�n����������xI4�m�t��^�R�����`�����h:�v[�^f߷ wK�eg�����q�G�j�H;PeC¸�B��� "���w�N+�z���3��׮!���rj��|���+�ㄝ�*t�*��W��r瑷=�V�Q�3�m�BR4�?�_i�]��uʰ_t�]t"!��B��տg]cCT\�o:ظT�y�_p�O�&�[��e�>;��&���׍��O��7&nc�wK�c� c�mV�`�/2���9H�.pCe����f'*�DwS�2w��j�z]bD��O�YD�w㢝!�+T�xu1 �������]�:n���}�����ɶJ�62�F(�����}/�k9n`S'e���.ǫq�F��e�$Ķ�]���>���+����~�9�r��Ow5eˌ���UbI��,p��M��g>�dLcSpel>W�V��6��G��s|��)G�̏�W[8��%�7hNٹ���YY׉��g����;tBŝf;!�ti�����X�'�H��/|
?b�}~���Dw��-��m�ZuA����
�j��嫊k�L��g��&w_+h!\�}ٮM̬Ju�e�x{�=���������Yi �:�T�vGs�ܬw�r���Ú���nڮ�6ܨ��S�c�����:���r��p�K��>��+��Ory�z.9�k!�:�&&�3d���ӿ#�}ih�r��k-���o��;S)�׼7v/s�%,Vdl��݈Ξ��x�7"gtT����U��U����R��o���O�y��y��c����s5�5�.ߔ!�GC�X}�X=1�⣅`C`׾���M{�1��p�[m�î}jo��]eN��S!Х{��,J�}�`�đ�\B�����)][��eㅴ�{p��D�Yu��!]�.5�\M��j���]�[돫�:�KMAI��s����j>y�+{p�el�����Ӝ�{�ۙS���/���ݵ��\S��3o�D�V�Z�a[g1���-8�GJ9�"��oLf�{}�M΋�K{��K��Jdd��:���^=�mu�n�3�Ld�)ovV)X:H=��d=�k� d�H�Q�|������Q�Q��婼��R����4��_.�VG�i�vu�����̼����to0En���E�T:��p���UuN�9�;��}}�[T�[��������<��7��D)����>��%k�r�vb�ȭ�j*���4�F�faƗ5a���W�O��4�=_��m�VJ:��Ìw	��n�OK�y5ӭH�O��L4�hTg��O!���R�Or!]��u�%�lu�o2弚�[[�]�ک��8R��}�S|�/�ֵac��y�o�^������lY�m-�输����oy���y5�ō�ry�ʗw�<�)g�w��g�~��p�nNv��������܊ɫK�fE=9=�7*{����=ͨWf����03��sUH������<z\�QjCٝ�49F{�3��D�:ɾ�~��:�@_R�#k�[�����q����t��Ȗ�\�͸Oz����<����q�զ�e��k*T��tF�j�0�1��E6��_9��u�'o��.Mˑ>y+a�EI��T7� ����J�<�v�n]��F�V]aD�ʞk;m�*XWd��D�U2^��y�o���dԘ�؞���O����z�LP��X�"\��+�><�����:�{	����CEm7�w5�����;Y�6r������»��Ri��3���0*�/�u@X��یp�\=o�
 ��E%S�ݭ�Vf��]

V��A�	d쎩�F�{��h�MT�5om�[P�Iu��=�Y�m�7p(%��G�}�* 4�⺓C�ЙBC��;[j���n_ܱ��q���t��()��ޘ0�KB��'�v���ɪ�]�wW��m�m+f�n|�h�x�T�f�
{�юt�b��r�װґ�e<IM{\����Ū�\v�i_��ٶ*{]�|l��c&u�.r_>K�YYA��I[sy�F�q.s�	����c�fط�i\��f.,��yW>U��xLFS;Q �P:�
ܚ��s�g<o��K��۳vH�Q�<����%��W��k�'���<��±��-
���N����U+��ޮ�Z����Q��ֱ�k�b��y���P����7�#]�4����
�>�C�L��x�m[M�:���3��y3]Y$:W��vܞ�80nB]� F�NVs�Ǯgs���0���`��v�A��.�8�mem�.W^L�ꐥ�v0a8hq�����LL��$Yw-45l%���#�w�'/V��]���m5�Ƨ�ӟ���{-mr[�	iKKhr}]7��ދyP�Qⱶ�e�N4G`��O��2�\s|�S�ϳ�.�ƬI\��ӤK��,n\��&�+蒘�¢b�!]-6�ކ�qۑT��3�g^�W����|6�����ֳ���K�Q��4�fu8<��.3{fr�7�pO��{��*�:�΁��� �/�uB�SΝO2Y�V�I���x��_��.o��Ox��Q��08{�$�Eֻ/Z����)ߟ�������,pը�jOQ�v�Ǡγ��ޝ����EMk=on�R��)<��<����+:Tm�:u�z�0�Z�i}H(p5h���_.���������}��^��Q{Ȋ�<��)���vB�����P9;�]ы��4�֮�f����+(�=�:�EӘ'kr��7:��\V
4��Z=�9p�IuK{��/7�Ia�ڧtnjn��Z��
1��Q�7������f�I��]�M�n]�'��rk���nȥ�훕� ���`�j_kaV_.�ˠ��;��A��'������N>s�}�R�Y��[4�S!thN�c�����Ɖ���1B��n����\_4�v���W�R;Q �s�Z澝��*���6on�uHV1�٦y��u	�MDsLTCn1�#p�|����\�u`�7gd�:���y��]봡'SP�M����c]�<������`�@���t��ZY��u�~���5��y��vz������8i��Y�x���S�;��Ө����V.�/y��rD��o����V\KT����<��]h�GEܔ��9�'�/�l_4�"��b{x��ǁ�[KENhq���=�}��H�����6���=�kW�6Cǈ_;[*��Vv	��)��C�؟�sB�R]u�5�"�,���C����<����1]6{u���tj�2���F6��o�!�>�7Ժ�����j�Ц@ՉO�>�zi]l����N����ڔmuq�O�h����q^��2Ƽ��S�^ߒ�d�b���*�h�ή�=�t0�9e��kEEܐ:"Oj�œ�����ga�f�������!�B#�o*c�J�hsV���興��R66�&�/���O#�=�J��o/5���i�5�3��'�h����3y��ѷ�0��Dw.����HLF��{�/W<�ё�d(�Y�^�1�^�[ٯ�X��!}�%Aỏg�J|h���I�eC��{��}SvE�ڻ�RR����t��Aw���`%��j�oo@��3�OE����qZ���W	�
��ʈ�L�!O����d�tP���s��s��Zc��Kk�PL��	�{�����ШN�[�k�Y��-�����w���N�c�6�V���vNo,\Wܵ��w�n1�#p�EڬNw��`Vvw ^�H����`�ʃ���f�����z!cSQ	����ؽ;.��<��˹�����ԡ�:u������-����ڕ�u؉�%���Ѳ���/��v�ʨ�f��c�^���w�O-���C��+S�?%n�4�e
�u�* ��*7���(;�٬7����
�� ^[B�V�o^Wn��ҵ�hNȌc�X1�w�0MH���kw9N���qm�m�5ס�� �QGyr�����2��nMk����y.ӽmK1�i=m���,���7�����j,«���=��6ݴ�r���;V����n�mj��w�m4����!�So��r�ő���fF�'u�U����X<n���J1�+��A��e>5�Rp��=�z[�e��F�:I����z�K��ٴ�j����C�,U���X&��|�\�ŕo@�N��z�E�����V��b��o���V�>44�wuv�qۺ�e��j�:��M�F�
S���$�M��i�܋�z�7p���B�X��^�
�����e�6���⺆d;֣.ӵPX��F݋�{��[�uZ�ڨ���*����S)�(z�\QP�X�%�\C�Ǥ�)������u�J�04�͘�s3I�^��8WH����>�WP����)1�t��\��n��|��\+U�s6V�w�VR�|U�բ�32��s{��wiն�8*���{$�W��^�G��n1��,�չg�V[-��k�b�l�t��4�q�E�0���h⃙0f`�ɘ�mw7�b'�;J��IB�r+�TM�W̌��$��ʛ�.�9P�sBާ���/�:e�nN��Q=[�[�t.m������@X��aTw��mj�B�����U�ی��++E��+�N��7LF�mfttK7£T.T�8�nywWy8o��u.6ٝذ�cVo9]��5ip*���i���Jd5�v�}GJ#��MлT�7�U+,���]8Q�E<�8�¦���1����s��5�6��m� ��)�|c�Y�e	X��Y�V�d��!s�����MAmm�J�k�s�m���#!y�wPE�m⾬&��b-r�-�U<�y+�uad��$Yvͬ�̞rE�Ֆ-�[So8ǥ�<1�C�����6�*�&*���̼�|�Le��z���In�<�����BYzks�8$�ւW�s��QS�s�U��Xd������+�#1�C��4��_F�维�%u��p|e�潼�	o ��ej�r^��д�I[m��[]����={�Z�nu��R���f�I��6��O�jV݃�V6�p����Xt���%���>4�r���%�Ֆm�F%{rjs�pC�Wv	W�R_H+�UX��*���rKK�7�S�e�5���%�3��t_0�軔P���]��9�5x��[�x']2�r�nh��yA�K���ѲR�\Co&���M�t���{�3#�3[�
�3�dߔE�ͫ=��/Hсo/շcG=�����v�T���k�����g�t�;o8ӧ�#]�pm �f���Sr��dћm=iԅ@���@'9t�+��@�;W�b�����\큱h��1�˄��2���o%���B� (� �b��|�eEb%�D��D��J��<��-p���4��s�	RO+ST���d�g��g���iQyQiXjDUH��f^�d|d|��.��"`��),,3е*,�!���VXb+�R�|g2���O)P) ����J�)L4WBȯB���Qr�L�D4�Et<���%*�sʮ��[%��a����#�#P�7��J) �r�KHܐ�5(�R����r�C"�%7%�5(�L��OAv��1TSI
/,*ą(UB��fñ�"�K0��\��f�h��Vʔ�Y�u1#,����^r��GH±@*
�ʡ$�����h�B�$�HY^Q6ک��+���4�eZ!R��A�.�R�\8{3r�������p��J*�k�yG�D�E4� �Q"3T�T��<L�S���ꞣ���Y�QDTDAzICA,�=#Eq#���IW�QEQ�#�9��F�.�3(#�z5r|=��ߣ�¼��7�����6��҃����b��䔻k�Z��jg:7ʆ�SD]�m���a�d�b%����y�τ�?꯾���y{'�׎�WY����k#]{x��V!�Py��4�ӓ��X�n'"52�?9�6;�rV#��ٞ���(���U�몹
�� �̱Aɻ}y�q�x�6q�u����Ruu�q?_$*:Zl��~����2.{ݓ׸F6v���ȵ$�SRU=;S����}��Q�7�M��}�h� ba�*/P�7�;�N/l�����PK��s�ug:W�in��Z1F����US�YW�[��)�Wn����C�� ��Ƿ��F�Ƴ�C*�o��O����������=T�OmR��g9��B�Q�T�!���I���E	��mwe�;�j
O/�x�dk��x.a�J�P]��AsV�t�}y������Ҕ��b�]���>��\3mn7�3�.��1F��n��G�Efbi}tƃ{Gk��⺾��Ri/���!�a�� Θ�0^f�v�`E�|3��͜*`��6��Ȯ�^�:��	��8;�fwX���{�w���F�j��ժ�9�\a�$��wofY�d|G,˘Q��JpSte���%�uwwҹW`<峔 *u�8�a����go\��}K{��m��Jj�ke���菾�m��-�h�Y#l`�����3y��|���7��;pwz��	�Yz��U��u�'����r6��9)��ќ�����t�b��F'&���[�e�4&�q�
ȍvD�!���w1n�y��L2\��=q�K4�gV;�7U)��u��[��e?\��Dé�wiJSENwr���M����n�+���ë�}��c��p������GE��m'����5mDM��Ix39�[N�S/E�|�S�+
|&�����׆�^��8��fW�Suy��=��\l(u����w@!7��֩z�>��S�y�5m��^AW �T���`Q���l�,��;"�Has��z�
�ekۇ[�m�Σ��1Q� s�����>��)&��v���%��eh���6��=��kj;l�Eh%���/J����z3#�h����t?YDZp�<J\U?G�'������&���wX�O�:��N&��@o/|�Pk=����vT�h�����0]']}{�oZK���[�FWS�ŵ��3�u3�k,e���v�"���˷i�JN��������{��
ĝY�����Tbo1�V����4���A[`d7��m�J��$.��o�T8�gv�Pu����O.9���ж�q���m�hm��Mvc���I���͒�\��}__.�O�|[������˱��i�N�Yf!�"|r����_g���>}�*7v9uF.ʎM!�b`���Čpm"�Ƹ*�F��_r{P]��Y�P���ǗS��/�U^�;{#�q�zu�w�|��a�"�Q��t6� �ra�]�$Lfn�R'�T�4�-q��M�M}�4�Cn1�7	���Z��NG�Y	D�����+�s/#5ⴝJ�
{��mDs��vF��qE�����f�ṏ�|������";��M�o7�\9�yJtP9��g�k�M)~���{q,_�Os�w�z�s����kg�fy���[�,�ev1��h��"�ױ:�V��@�[�8�jM_Y�g�_m��P��E���k�Ӿ�E���g�z���v��T�p�u����'��n�
���8�R�{����io"��!�f�R��:�G6z���SA��)Y7w�5e��gs���}��S����>��k������Nя�~�?_5�G	�W�<^�F��[�j��9�|�:��:p���{_C��ߡgt��ѵ�V{1�k�N٭���q�P�g�@�uet��~�,����3o�~��������蚱��WBW�Z�-���6ާ\���T.��H�n''�9�y���%�p7n"Ou}:���*W[��f5��ʧ��^9��N��e��V^$����(t�h��`-�;��uR���8kI�og*�[��R�cL�v�Ǧ-;ŕ	cw���|��V[kk�g�w�[�#y޵5�]��WKܽ{��uC�r�ү�P]��|a�	h���fwee7�Z|����I8�շ���V�`��ʉt�"B�Ѷ�Q� *���x9*��:��=?_i����7��hTBw�t�|�=�PDsQw֣F�s�9�{hbXvA����Wʅ%pR��V�on�%j��V���"�YNY�����^�����)�%w�;��2�e��9��!+/��/^� ɽ����9r�ي�����C+ꒇqR�K2��8Po3�Ȝ��_��"">�'cH�\��~�~��D�ɬ�u�K\�4ø�;F�a�Sdp}�d�rQ�h[�u��x�ќ��?{�7�������=�h�G�Mr�Z�拉��^�U�Ibט�b�LB��D���iM�,����:�3z����<��vn�X�{"�%�';YULε�==�����v'|�����O�����k;tn��KDL�9�zo��l�Ho@��r����h��V��S.+�v�U�k��.��u4N1��۹�w�a�\/~Ëp?B�V�{��w�k=�kމ���2�b�h[:j��o��v�Vxˤ���qt�C�Z��ب�ܦ�-V9��ǧx�Uok�<���K��V����0
�%�D�@��*�����l8s��2�ko�nb����'���A-p�?Ȏ�9#[>�����u�Rw�������Omd+%�9�`J��*�r͢��������R����Qt��K���6>vw{�UGuu����_�
��|����$N���l��G`9uun�r�J�𐬮S���5|����ux�m@H=�.��
_4&�t���}�}��yor�v�Z}�����p���[q�n$%��P`w	jv몳����(dʷ�o��w��?�kjzk�ˎx�d}�3^
ϛ��1�or��b
1qsoy�B��;��>�O�7��5��h�x�ԺQ�"�}���Tќ�ֻ���n��k�⺱q�I���LhL�[�[T� ��;Կl����o��b����X���sܺ�:{:��Tm���p^�ƴe�W� +�P�G7�\l��;���Q��q1\���9� �ŕ�یʷ��<��MF'�����9�����S���w���Q��k��W�s������V+��R�
i5jʯ��?\W���,�"�Vݜ�Y�b���e�<�Y�n�Q�X����Ú����_Fݛup�1��q����+��f*���Ȍ��7);S/G7��Tu�=L�,��#3)�|pTr�y<��:�)!n�ecn��[B�V�naS������9E�I_c�Iu�k����oR:�)L9�쨙����ݹ��k�9�\ݝƄ�:%u'ي��y0���+���
��:*go_6���P�lF�fM-���U_UWU�Շ\����句;�vϢ��������g�M�z��l1�cv^^����T�Y|����k��3���-s�n{��CT�T*XW���Cqx��#*�[�s��-�*���vu������U%��gm��wVm^��y�8�)���.�������UDV��:绪�ñ�%H$�����\]�T�4�����1����ky|(#x�%Lq�;���� �����KN�Ryq�=���=�(�::�p��]���Q��P��;�s|��u�.�O�|[�O�p�%ǫD��\�
=�+�ܛ�~�j{��0����r�]�c2�0����U.q5��Lu�y�
m�.Y�B�;n���jt�=r_ywX��^J���v�q��).j��h+�aJ3��y��3P���L:;I�se�=j!�a�nv֝���ҕT������ӕ��lS�&���oUb��6Eb�n*��*�%�E(v�����i�]���F�f�\cq���I�9���3:���y��y4��씅�5�86��lr������=}�r�hT�juG��D�ɨƞ�_7�<�@n1�#q0��?r�.�D��3 ��7��ڷ6�y����[_o=vک�X�M&�]� ��E��]ڱMZ֣x��`S�he�VrZ������֮?N��������T���#]��=�lĺ]�V�1�������m�Du-����������^�8��y;����8������5�4�z���Ir�����?Z{1��E�U7zդ:׹�p�Sa�-ۈ}�_"B�֖��~�'�n'Vـ�K�ҥĕ��=�ܐ�%�z�[Ψγ�LwH�LR�&�ś6e@괛��nzUD�CW��j�b�or"�}p�\)��]U	;���׶n��tˈ�����}_N�
��z[��e�o�T%�F�\�H��ʝ���u�k������l�_>D$�"��)Iϵ'�p�^�bs�J�d����&�h�p�@��E��v��^��g��y�{#������q���K�٧�zҔ��: .��=~���]u�P�R���݌�R�u�RN��C��%.�4~����1w�-U9�'M�>�a���j�r����U|]��$��u��a��Y�����ޒ���۟>��42:��t��J��jǘ��y�p�5ٮ3��9R�+�PS�oO��Z&�oOڄUs|���7k�U�v?�wTc}���w�q=���t�|�K���Μ{�*���t����1�7�N�K85ы��&���;�;B�7�P]2��An��a-Wɥ���A�^����5�ξԎT%�i7�����`ٷ���N�r�]2�N1�u�ے�&�y�mR�������q�B��Urץ��X�Ϋ�����/�����=<�ݴ��Fb؛�٤�7�H,,��]{��ㅽ]k\9x����UF�7�tR��f*��$�w�߹�|/5�8���s�Z���9��Cj�R�7X�ecs�_�9��7xۮ����U'�fr���ݙ�f��Gؓ��j$�����˶N��L���S�ۢc�;��f�hs&���q�)nD��7�)�)�*N���t謧2�gb��q�:m%����T���φ]��Mm�md�;��v>N�x�A�N�ԦmM��aY\����@�g��8�Y�ZC����}_W˔���o��a����5Ss�&;c
���GKM��z�ᵽ��vl������X�L��\�VQ��!�E\�;����\ip�669��I�R&�3��;�sΐ��d�f���Җv�@����K��W؝,檺v.Â�ͯ�:�XZT����T��{އ�ޒ�M}��x�=���	���U��.b�Г�/���v5���I�j��c�m=���q!g�@�*63t�9/����1���_JZk�)<���]��3^q���E��5��7]iqQ��R_RpWڴ_�����>5�o�ٷ۟C}��x����qd%:��W nkq�ո\Y{��0R�]p[}�BMq�'�Wj�k�m�`\L-:\^]���5^�o쪙ҝ�zd�9�m�oˠ[v�f�fl�\:^k޻}7�./��;a�q*P��v�t:�sR�%�[e��D[/0��'����,��,#�1����\h˃zr�U�Ѵ�5α4zԻ{t+w�V-\��Z��u�iţws������:���;���N�K A���n::yuZ�z�-%f")�t=��4_ʆ0�$E��`���X��ˇGO�X�H���[���s
�V�̨%um��q
k\���s�����wv��'0�EuL�v�ކՀ�p�"���+��vu��Uϙ�}�0�)�*��Z�+�G�m�;PK�A[q#ҥ�9�Qe��6��]�{����!j�4���2]�P6�$L��J��imutӦVq�6�Z���U�:�Z��/m�§ٯ*6��u|�B)��J�ۺt�୶ޮ�s���,�3y�NGS�u�Ƈ#β��J��&�|����:0L�3U�B�Rf�Q}#ε��8���K|��{M�ЈG)��Vz��ܹ���4um�j9���X�5!��c�����v���ʅ�3�^�«�N�tns��c�Jν���V�A}�71�yȬӐ:���p��~���vr�}ob(V+�̏���[��*���w�u�bM٬�t����B��4+����ψ����LEZ3�}C_M<�U��Ľ6�29r���a9����H���JH��mDj}��h�;��Ȥ�P���ô�M�<�0���NZ�]���q���;�_V�ݰ�Y�-5�6vR��ս�챛C&C2��Uc|�J�[JȜ�T������I�:�00��x��%���շٓ�ܹ�%n� 󭚈�t�(�r#6����+w�f�l����uG�Ea� X�R��|�B䘩�b����KW�q��������t��s��s�l�F�͡)o�t�j��K������B. �1T�)���]��̭�n���\;,}�p���-��WWF�@��}i�=zeh�Y�G��Z��Z�2q�t����Y�%�5[Hwe�`-��̲hvK��YJ�Lb荻;M�[tx�&��C%3��{Y>i���eѺ�PΖ#o@-����0��$ws�#"��a�UZ���*YUg5���N����mݽU����ޙ��og[J�������Ǝ�e'A����Z�}0:������m��Q�ǲ���Dvb���\(�L�k.g>�M]n>��L��w��PԹ{��9*�D {U���YyC@�gskS�Fsđk�u��`��#��u�V�,-uӅ�3�w��,{��G�XӢ��O% o��h@1�RF�8E���k-�}B�5�:8m��L�Q	����)��thV��;J�5o���Wt��+8�,e6�$�b�Ce;J�J��jj�Jə;;�h��d:$���f�*
`�k�:k�X|S��l���4@�0u�_S���y�\Y}8���gR��q�	�ů��5+ol��/z�,�5�w�"7�l�b�9�$����w�c�Ol4�,� �h�� �I1u=;Y"���۲�䢦�WS�yAW=�6���u��Ȩ��E��"��Y!TJ.QR�&�)n�^�QJ��rF�h���,�iGm])I	��eg:f�mnPq��/lHd��(bNy�2���"�M��Q�\�f#�KFͬ��D��ђQ���+�Q��e��U�%3Ă�<�򣜺-�X�d^�M��L#r³�%�����Ig:X�Dg��2H�.BRue5�a�hj4��.a�I��Y�Y���<"WO<�"ˈWE�۪����R���	�jn^�(�T��nE��4R����S�hZ��M<\jS�D�ndREE�x�۲*���6.�Xy'=�Ԃ3"�0�/cl�zg�y'�bf1Jdۗ��H4r=h��Q^�/*��l#��R�2��t��JM�fTI�GUF��Z6��nq�0�Qt]ZQ�H��$�@P��mvE�u���h�L�����[��u�a�u��[�*�f`�W���A{N������o&Z�1�b�����P3�����;Z�==����K�O�k�bjq�
��vD��>ƌ�� 4���S�Z�Q�q<�sloV+��J�
y7Z��Dtk�m��C$TV��i��+,�ǫ������/��sV�e}�*�K�����7�?�4d�������T��.3��ܤ��2�_7�L�&���.�C�(����8���\H/����~]�qn	��3��m0���'�������K:����4��kz�.�saT��\�D����F9���Ւ+��C��}gtTBI�p齸U۶�*�:����ur��S�N+��U�Qxs��k{�R�2�[����{��g���:h�Wj�pM���x��X�|�x��X��SJ��o/�p�^8[I���-{�\�TO%o�L��J�m�ʃ�W�R��e-5Rys��ޅ�2+���l�${�����\j��e�O�7Q�y]k�<����NW���O�aY��Hs�[u�m�דpߙr���ُ��;�{6�J�E�'b�[�S6kZ��C��&!���W r������{k3N!�)|wrH����Kr�vΤ�l� �R����Ut�ZW'����weo��AJ�zJ�&/��T_R�����4�G��\�#%�V��kƸ*���ڈX�(�w��%���Z�d�[�sbS	\-쎩I�3�Ӄ���z�3�+�m�.Y�B�g�A�ϦUj\v�ĕ��֕���[^��������w�v���aJ3�����K���%j�Sq/�99�pk���r3�ԋ��i�p�v���������Q5��6�f�r�2��֐�wA\���<�sg<o��MB�
k��k�u;~4�瘘
�o�cgޙ7V��'o,ǵV�߳�,��*Nz֮?N����q��̅&�;V�`��q�Nu,��f�5�������m�GRѷ��(T�޸zz�-Ӕ�3V���jgv�I�5���?ٴ��|.�~_�j+j>�?q巵��ЭY�W^�������L��:���g�ź�im7'^�4�Y��)iU=m
J�L7�0���:c�����k*�H�=���$f+��z=n�����~�]r��>S�e�oT�]�w9�!�gZ6�+ΫEdI�4���Y�5���O;fpޡ��|�>W�WL��R{:���H@	ejW'�G�=�;�۫�^��Dl.�.&/��!�J]lL��)�(C� �̨}��<T��%���z�5q==S���-^�cM�E6���>�������W�n\�[��VQN+@�)Lʤ���bR��-���y�n]���LՇ���XȲ5��()Z�_>W�II�uR��Cs�#闼Ss��<�O5��+�s5�^�e��}�0T�p��v����(&��xf���}�k�Oj4[츆����񜯥�W���z`�EgE�U9V�T\�CR7z��a��O�ඔ:Չ��.Y�D*�mv�+�UA�P�cI}t�	��=��8�Q���&���;�Я�j���K�f�3h�v��u��ur+�J�%m�Fo:�H�|�9�������Nh����R���.�U�YO}y=o*�z���f���S�����'gbo1���v�U�D{�~��q���!��������������V����˲�	$�o�B�:��fnً��c+B��okN��9R��U�Xg/KS:���#A���3�8ӈ���"	�uK�Ӆ��������՟���J�Uo���_4&���)��dLG!�y����^ͺ�q�ܽR�4����
��N!7]k\9���s���F��-tf 0%��왇؊c�zՎ�X�8�n�r����_Z��F�Or�ٽ�֐�+:I^�U��T�E��톔^���+F��b>���;5SϧLI�ݝZ��ݷ&���w�7�<�Ҽ�F1�E\�Φ�Lu�|�����u��b��2�K�?+�N���{���γ��es �TK���_�\*���T�%/^!�g��������5����ѝgj"��<�D>��lw4�#qnԋ��sN*��$VS��Vᬶ��t�Z���T��A�>V�����o��VRq���]E&�\5��c|�n�����5Z��	�3W�*��u�:�R�_�\sƻ>����}����ӹk�c�հ1A�+�1Ԯ�&X��T7��t��I���o���@�δ���+;;X:�*�g��k�lV��Vd�ڎ1%�@իk�H��ag>̭��u�k�\`�%̰�ܻ�Ybr�3��6�)Wk.��0p��m�=n��H���/1�=�}w:EN_�{��E��0\	h�Ϯ�r���_Ao��}��h����E�>;�rS��U�s����;�����Z븮�\v�iuWZ̧lOb�"pd$��w�q��Av�q[��)���y7��܆D�'DQ���R�kӨ���)� ��\O�P��v�u:�
�8�E����aԘ맪D�bme���Y�ᾩ�i���q��F�c]�1�l�-l%J�n[s��[��,�pk�\���y�Պ�'SK)�����]��*��#I��j�b��O9y��ۑ-�yk��{�6������պ�f�)z83g�z-��"A��Q�*��p��e|�{i����;5�n�I��к������}�������ۣK����yp�U`��i�y��nS�ٹ��S�wW6��s�u�k�����#.�Ts��s �W���.��3@�eL��*u�T��k�xf2 B��6����������w.���t�3%�T������t{����(ͼzi�b�^�c�.�/:�9ܔ��^:
��CQQ+5}
�q�}�.�3�GJ���Go���RupV��2]���]�S���о�\��cm��X�6/�M���s'�|��t�7]��{�J��m_vkbn��I[Q��3�Rje�/{�+�}���]��;��5���������\�,�t���QIR�-��8k1���4�;�}q�v���ί��������*������ZBN�#�5�9��L=���V�[x����9P�7B�zJ�b����C����%���;1?E�7��|���WglpS�<u�;۝
���V�W�'"���{��ғ��ZI@w�d3�)�v��4�\B�R�Vp�(l\�c)U�����K؎\��o����!J3�v�;�����ǰ�dU�#/9%�q�ඦ�Wd���֤[}3��0�q�������=�0�mg=�ђ3b���/ծ�U���>�5��5.{�~>�nmW/Wdw!��0�D�I��n�ȬRW��`*��gb���
%����Ɠ���Ä=��
��k�y�4����nh�{l�mfEY� ��f�?i�z�ާwdMKé�����hokt���4m�.LƫOcYD��|�^>�@�������Y��9��~��ʧ��j��{��6��,��$�֮w�S-����3��CS<��zdx�f�9y*q<�s�u�t�}Q1T���Z78�|;��s�]�t�jւ��.D���W?�Qڇ��H�s��"b��=֣@��ug��;��'Xˌ]m4O>�W��?{���sj�!mN�����z��nޗ�v�����u�P�3��>�՝�ݱ?x�+�&�]J��w�������/��� �s���2��F4��6���2X9�}z���uY���,O��Gu���f9�I|u@�K�x��)p�+P���I���D���[����+�PK@܂��ʤ��m��� ���o1�i�_W�����9�b����|��w�[��m��u;�$�6�SW�����r�-�[X�dk���ˤ�?w�ԾF`Q�*ً�޺�"�y��BH1���Ɯ���-*8���,�;�P�I�cM���p
y�\�R����Ԗm�٫O1x!�{���}��P��,_Eλ����r�Z��h��E0��P�-q��[bBsr������<w���5�ɓ5��S)FM�%QN�+��c�V'�p[JýZ�`�3��V'/J�2�M��o�[ϖO��Zٯ�kˎ)b�ɥp���/VM
�KFu"�v��ʯ����_ig�.�k���#7�}����0�'�d*ۜ��R���є2-E����(r��Cl-�Ȟy9��e�d�GZ�\\l���fWc��SK9���k�����]�<�H����OfN�YN5քCۥ��O��<����skR�u�-p�k˨=�-�~ �����L6Q�RV`Nv���ʶ�M�q+�m�[��㜾����]�{�J�� �6����v*��t�^�\�ǿ`�hҝH��>��;3Ϸ�]��p!ʙ��_.6��޶˘$e��\�"nr�$�:𨟯���a��>�K��]����A����tw{˼������G��9�웏����ʸ	��jA�8�"�nA��]F�Ԯ�q�bYe�V�cv�y֡�ՙ�����8tR��:m�b���[�։@=���
���L�(wϨ
Ne��N%�R��<i�9]	��t5�pb��a�:ع�Fl����۬����K��g�Ѥ	3��%�kfX�}Q�}N�
�i]����Ry�����=5<�~P���l�p5_�_"���Λ-N��M�^@�ܞzSn���<�����UV��C����M�A��csV�3}�"K��]{���7����1�ڄ�ۅ6����e�e�y���p3�r\� �.5������KM|Ry�����ͧ�s��Q��р��í�W����(.�^}A�%��>��r�O�o��f�2��mj�:b��8}�O�r�Qp=��H�"��.���Z�Ջ��}����ǯ��i�:�����o>g0T6�(�e �:B�|S�+n�-���W��5��K�L��Ӊs�օ
�L+�˂�|q���o%K/����kLE���U��'��[����bzq���2�}��*��� ?	@x$���tf�hM8a����}�j7��	:��c�5	�;P�Q��E@�-��0����4���5P��݉����TbcĠ8��܎��e�Nh���JB7H0���i�m�����]���^=����hˠ���w�{)�l�v!A��s)7�%t�M�����jWG[bY.�[Џ f�]Z�[ʗ%�S��B� �ǧpp_���r[U������~yX�9�녮�L��e���k���5Q��Rov�/Z�=�������VL�w�ox��yͮիr�^Ʊ�|Q�i6�t�osk�Wf�X̢�`<U79Ry�ޥЭū6*��KI�[��
e62����������rÔ|��v-q�4��V�)�TF��=X[�6{}��~��P�����Mk�{J�@M�^ru���F��ކ��0�+5�����5�&4��)�{mQ�O��Ӯ�0y�Τ�T�2�"��z[½^�~�d����>w��Xj��Ĥ򗗯��X��h?��q%.����%-5�I��h�n^�7����"��Fh{O8�7Mؠ���E@I��	u_R�u��;�	c���E�q�!���5P�f�<g+�t�"}�������G��7��d�܎f�wS�1]u���vX};�/h�&S�Wl�@�9��L<�Z���J��"ÍV(��E��U�5V��D?�Po#�����ת��S�h� �yj�˦�4��D�:�L^n�
�Ӓ��E�]�L��xeCs>h-�XE�sr�`��84��	��V���U�5�Fs�W%�r�PѺ5�^A��(�f�&�)�%����ヒQ�k�楳��1s�il��hnV�jv����Ӧ�ہ[�7
?Wo3�!��EU�wuz�J
Hf�N�(-�C:�V���f��/p�Y5�N�d[��oW�j�ʵ�o	���Ӛd%e�gI��Â�Y���x	���p
���Q�zJ���v���7�u�T���+Q��+s��]�V9�%�@L�]�k*j�����}��;�-�;h+O3d�j�c��g�Ԣ�U����%6��]uz��*���t�ɀU;ڒ(�N�܂���%��.r�g:�@ v���K�^�n�R-5�(�{��\6��s�W�p|`��NĐg�볖.4iΝ6�B�V�yN�"+3Z<u�7�Fz4�7p^p��J��J�����Vh����2N��e]3��-ޛ��#}��}�f��q��N�i�u�.E���.&����d�ɻ�+���N-T3)ph����_��&��Z��yY�Y�-��p�GlV�7x""ao}�ĕov��K��m�t2����ep��9L�"�&M58�ν�Qߵ��v>�v+8E������ն:��@V�RZl�+5��-t�����4Y&>��D��R���:��Ҥ� �l<5��B�6k��XZxY�J!�W��ͬqh�*LB��[V6�����osYeɁ[�sN�b���klښ���k��]�%�cu;p��uGϢ�asb��4�[Sql��u0qٌ	�vuo벆#�{t5�P���'H*��T�E2���y��H)[��^M�ue����ko��閷�IƗ2�]+��j9����3p���V�]k�4�xM:���<ѻ� Y1#,�*;HF�}Q�`r�K1��DAYK
��+�äq�Ǹ��k��
u�k�ĕ�H_>�u���O(id��b�]�>B-�ۗ��i�s~u4g�K��/(��VU��w@B�D)Ѯ�t�`�3_Mɔ8Cru���V��Wa��
�
���<�l�+��|%K��&�b](5yi<�����Cɢ�6��j��I����A��	��;�W'J�jaDff�_n`����geF���6�'Mn�9k���c�y�D��雉Fviɥ)P�uz�	�Ue(QÇ�C�s)M<oywsν���Gx��d�#N:�+)V��Y�oE*S��"bcR6�h�ڎƖ�VV�����^R����Y"�t8���}0�\�D����/1�\Z6�e��slf��
��hdMMt"Z�:�r�s"�� ���'c]�m��P��.(؍���-2�Jhb��WZMdp2�(��g%]P��r@����)�����im�f̓�	�P��lX�8I5�a	I�涇;,����Y���Sڅ�H<��ѧ�r�ã���44�4�h���2=��DQ�\���FI�s*��d�5�q*�"�)[L�$��g�]5A��a�i�G�9�0�L�U��r����Z펄xfUfH5&�:��ȼ�ڤ�Y�c
ܓ�m5��u�K���ܔ�s���S1B�A�1��w4L�L�d�E:�L]K��"���iYUJrE��QQkWclH��eV�ѵ�k���U[VT��)ZeL}�yߝ������v]-N��Q�;/p6Z�|*Jc�m�S ��\�kJk�+Y�NꝍJ1k$�塛;%s�ɗ	�wn^�~��Ջ�l���z�ca�v��5�!Lt������Ż}uq7/sA��sR���#��(�v��;��R�)����/l�@S}�i4���v��]�Q�֤]7�5�0�7̑�ٛݩ��ZKT���y�D�?��;�h��Y�sڧ<�k��Á��[5d�������:%�^Q�5�|k���/>��G��G��9��}Rs��<�4o��cq�N��[��\�×sӎڨ�p�Y��=�]�=~-V�H:ei�ږYR)oo;���y*ܮw�{q��5���|��P��c0?]��ț��P'({����g�$����O�m;�2��sx���ͤH[�nk.*�v���<�;�[��ѣy%��¢b�!Py��DKm[�͖� d:i㧶 ݳ�+�+��{eJ�W|��s��ꄴ�0�*���g�
 `J��1]G}id1����/�zc�Ԇi������=�c�tݩ��+�i��U��W���]+�Qd��K�_�z�M��t�n�^�˱��R�m�>�_,�9�Y��B�ØO ыP9Ќ"o���Zц���;5��������Tӻ�6C���!d����s�3���H{顽wn���/�'TX�'g���|e�7w �^o=��̍Wi-p�=��M��@�*ʤ�Ε&U��K���t�[�c\N��놱}���Zͷ����_Z9d�sW���j�*k����'r�-�[X�f��x����+��-�Z��O���澤�Z!�����i_�ޭ��EC�r�wa>l|�7P����k�}�ϻU{����U��ri\�>�Q���0��ua�Yy��*�s�*S(3���`�s��f�=���t>z��)�z��0�7�<�����A�n1�q0�	�Gh�\��5)��Yo�k���g���3�7u��{���&�]�Mֻ"~�:`Z���oaI���f(r�M�jv;\O59�3��I�-p��A��yU��7�t_Bʋ�1B�+����?w0��aL+�1��Ws}m4.��vNZ�`E=�q�xܺ�]Gj[����l[�цh�}�9f��m'�qFu��ǎ䬬]��F�̞Ҿ�ҳnLv�m̤����C����+<�K�5�]zD�#�R;���x��
�ӽ��	�^�]wQ<�m�_nV>e�-q�dk���+ko�R��\k�Js�q�2�r3M��+_��'춝z/��7�v`�OWx�1<���mR$�J�qʿESs�SxTL_$ɩ�v�S����Lw�o��{�>�7�{[��MXq�-9���b����i'�p�8��������I&����f��UFu���zX|'�a]%l;�{��$�b�oRT�4�*-�Yp�}p�>�7����+@�ȵ��fH"�R:ZiUC����E�%Gy�ᬿ���M=�6����}��Q
o�x9�p%��BK����KM�s��k��i��]�X}]<g'�ye,:����(9_oO�A	h���r�O���7?^(^��^P�Ц�ƣ�b����r�|�]��cJZ6������o96���7��!�i��ve,����GQa�a�s�C3��9l���pZG�����Q��w�<1��i�o���x)��^�ebdW_Z1�%��i ���7�����փ�.�D��H�^��L,��� ^6��� j��9�S�n#����q淟3�+���t�|�S�H]CA���L�&�����y#j�[�w��5_c���|�����q0�	��v���-�nQʳL��j��|���^>�Vw,�9��o�j9�&�q����vE��9{��A�$��1��/Ṕ�ٗ�Mf-��ē��8SQ	�;)����ng��y��"ܸ��:J:�%������[����/�N%�:��M���t�Ҋ�nx��g���	WZ�ޢy����g'4diy�7�������VͿ��负5��{{�+�u�fQWD��9@[ѷ'�zz�c�j��F`�qi'p�Scj���vm�9��em��ڃ��h�n�����ښ�NzUD����XS�6����o��W��u���4*�:r
�M%����^�I]Q���-^�Dc����έ��{A���Nh�c{�Y�p��奥d^��R�b]C]�����;�9ۚ��12�Y����%o��{9 ��Ax{`�HTe�� �n�a�����ѷ��R/�-���e�y��i�����t�B�JgzvU�J�me^s��\�1�]M3�Μ�ھ�%�kFi��%�Qdvֻ��(�"OuN�*���hn��p�C9x�nB2;3��Ҽ�k�5�gV_*�w2�A�>U%.���:�KL��&m-q[�e�d���iu��Ύz�,�r��黁A/�� �!&!.�KTV*�{S�5�ϻ-'���P[�O�8�p񜨗H�"�}�&Z1�gyӅ�Td�қ�sW���E4�!�Ԙ��;_K�i���v�Y�5%_jk�ۏ�ˤ�wÚ���#�5p�������k4��%_m�O�e�S7�ՋԿ}
�r��X��/��n�[5q���7R<=�^u�|��5~������.�{yW���2��q�x�t
�>?������2�v�j����
q�''�߶:G���m+��W���ĨU���8�!����aO�T���u��7�/����s���:(�#��+��}����޻G"z��mK��t��&r�|
4r|i��ǥ�@6���~֯[�w����+8~/iz�].�ڇvfM�C܅���\)-�c�\,���m⼟��/���\ל��Xۋ�!Xd,�#j��'��bܶu�xu�J�!�,���� '>:� ;��bv)����8�̛�����={s�qlb��7�����:}�>��WϝM{�b������]���߯xߎ38n��׺tH�.��땸!>(��O�y�å�u9GE�T��;���ny�x(uO��}S��z�wg��1��Je	�&e��^J�4l"s=ae@��Y5��]�i�}��\J��x��^�fV���z��
ګ��]�b��r�B�VT��K���Pg��^�F� �	��֟zȸ����Q��ֿ;�v�5�ֺz�x>����Y�/沤u��x��AS�ϑ��p=`h��$Y�9�Ⱥ��>�����}KNF�G���\{�s��Ü� �6K�s���,	U�� R��X���v�g���_�Nx~����:�7���9ޑ���gW�\>����f�9ozUH�Rt�7�5^�<:x��)T�^�!7�Z2<�����+����S0�:�E�<x;ӭv�ќ�ֻ|p�`��F@���IJ��
XW�և�y��g[���L�z����5�*V	]���O���q��" 5Qx���z���E���5���H���0~�ڠ�\`�Ȋ�'�OlE����j�� �JZ!44n��,[<������{D[~�\PrV�����Qy[��iн��C',�}�/����=���I�44�����s�6���8γ�s�����h34��=3U�GP�,S��s:�ۥK�=�&ܮ��K�z���&��h���s>�V���zH���z��Q|v�#z�x�Ü��U}���[�N#�~�wZ�p��@����X|�5
m��2�l��_N�7}@O���s*WOl�U��wK��{P�UTzϼM~��������/�x�|6�����Z˷|Ch?z��������E=�*�ݯq�YP���1�>�W��K�׶n8�������K<������&��n�mhwR�踥��{;��\v����^�,�~�ޔ��`���AX/��]_��%�^C���̩�zx�ۃ1�P'tÜ�q������<��W��?}=>��i�ߧ@]wY���r�"�y1�gݫE���|M�*��>�VUi��c�0� o�G�5/����s�=�����ƾ��:�<�нS�z��C6eᯌ�B��R(�.�N�qyd��;�;��,�}��!L�w�׉��~>�eǼVW��vB�c�}$���e 1{4I�3n{�ͺ詗��5@��~�8��zG�¢=����[���sX��2��3U@ߤɛ1頯=B���7�&s��_�9K��T����n�� �7Dd�[��).ͫ��<�9VU��O��
�=�>�ɔ\;{�#�a�X�=����;ԧ�n�� fV�N�:��Z�Y¯(T����ɲ�Y�qw7�IA���)w�B-p���N���|�+��T��]z\�sBq��4z;��cr7��~w�.�TVs��}��1�Y��/��H�'��.H�_Kjr��]7�$\��ў{^er�?d��m��Y��z��a~���>u�!r|i��|f	��q7�+�d)����t��굾L�Z�F����y~y���zǊ������߷�#��LNÙ.iSG�D�u��/��"�p�P���]�v�p�CgЗ��~��G�q����h7�����g���d�)T���I��5�;7�FϷ9*�O�{��r�x�Fc:!5~�?O�>8}9�}�`i�)\�鬍���#o���g�
�3Cb�+Mj�����G��Wtbן�ѿz}���dw(Ĭ7��6t׷9(m'�e����1�巣")ϴ���1���1�߮�[�Pu(�o^<�����ъE��]�U(��?N[�7��>�;��^��qJ_-J�8\s,��9M{+3������_�~���r��Y��g�~갮�E�l�v����C���6j^���Y옷Tr��ͧ��^�4x���_d����֬E,���C5$ʔ+q,��!�P�J�P:���ذ =�nW��/_����1vV6�����\J�-�bu�e�p�Χ\�U�v,Zu&����:۹k�x��:�g�n�+ZZ�Tm^��ϳ�Z��N|�^�|�bu{�8;7&��9�2��N��I�v�׺�{�5B�,���uT���r6e@��^w�SO���y���Ko�>ɝ����n��S!z�v<�Q��z�{Fz͍��GD���=�,z]�^���r=u��j�ެf:kν���Ŕk/{�'}4}e��C(���ϑ�rk������#=�3��{�Nw{}�n/���v��^cW��xť�,��Oi�~4eS�L�n+��%��m�y�z�c�0tm��Y�`n+�Z#�O{��#�~���.nPqD���J�0�L*�Q���Wt?��j=�,��d������g�=�>NG��F��|n#ڪF�{�~��u��j$�&u�X��j��n��u2)W���/�4;���y\MϽi��s�q��z��o�F���f��,���[K�8�1�0:6�<�0/��`�X�GȨ֩ϥ��1��ζ��g��������^��T<^���R뫬��3w�Iw�FԐ�=$d�54.)�x�@S���j�m�j���+>9}8�c�ѓ~쩷����t��H�@I+-�����fL�T3�j۹M:���:m�O��{���4�x$M�a*�Yս�\ް�-��&@Db_n�b�6:૬|�j�Q$�<h�rѾz���8;x��wlS�W)bp�B�;G�%*K�z���i�I�0�������Q��-l�ƪc��܏yUP
�?Nn��<WE�Z��=d�l�lTX�� �B�O@!����*+�պr(���ۇ�:�1�O|+ͨ���L���>Utn��t�^O������� �)�*�����g��V�o�P����"z���Nzp�;�iܬ�^�O�h�C�P�q�b��,!뙽��(���^�=�Z��{R�^�mz�{����wK������W�S^�����;�p{���>�����I�[����.%k���Ƨ��L�T6t)9'F�J�N�`V�G��~��u̬���ue���\a��9+�w�W�F?}��,�qd����ȱ��Zd�˴����^~���;9֡o�n����-���~��xo�����Օ<nωJ���Fz��W����t|&G�6������~;*�%�}�=�)z{o����<��\��<I�_I^4eT9��!��W��<�#E�xhF�/�8:���y�^ӑ����>�}q�)�9���-����$�D�G׳}�#E{tУV�ٻ�e�I@� ?K����xE����3�r�OhYǄ�9Xth&�mM����7Ĕ�FU�E7�okv�Jí��n�O�h�r���[��ڼ�w��t���n==W��m���6�ܸ��-w)��Ү��wX��&�[y��8^���bU�s�u'ɑ�qѺ���
Aփ�Y����
��u,-g+�ۙ�9tٿ���L�S:_b�t���ST��z+�֭�6_V� E@�5XK!Lh�b
o&%$¸ݙ���,k�]s3T�\�[*Ѣ��lBU�W��]�]�N�l�HS�HY���rS7�-9dC�������/�X�h�
,C33f��]v2�&n��U�`5�Ÿ�J��,����X�Cj�9nY/�d�b�.�+���}��QN�ƚ�/R꺏F��:Z���L��3���lD�
݋:�|M-��ʛ�),����mՊ�S�N�,9ͱo�f^�)h�s�cXӈ��-;�F�� I���a>�.�ƪ�V���/.��XvkO�����e�6qn�&�eJ|l�l�ݎ�S��R�L=�d���_MP�("�V5�����teth�w��k-�fꅼ�.����鎧 ���5�{y��ua��E��IV��:��3�-c�e �iH�AI�\���[y�bafN�UnEGs�ڷ��Q]�v���% (�ai�:����^^CE�r�w2�5��;��G��mK�3+(�Ĺ}$�`�9�<����T� �iY��/��F��H�0rľ�Kf��m��>�M;Uu�"���n2z��<�9���j�f֒0��V�XaF��\�qS83�}m�}]8SV����p��̈��������bg�W������{���5�u��{+{8\2��O�<�Gf�]�3�;��x"�ޜ�b�c �|��V�G��/��]rZ���4��2nF772�j#d5.�e�5�N��R���Y���6�մ�u:�ٳ!�ʶ͍��G,9��%x
��@���9��ھ<]c7�nJ�oVWQWW	*�'���$޻�]�$M��A���d�t��]��ȷչ�Ue���0V��-�&������GM*�zWWo&ٮ�.u�7;V�Qe����E_;-s}��6]��}]�
�3��k�E4��j�9��J��ܖ;�(�6�];��٧L�L5��RX�:�p������u+�2�u-b�u�0��:�SZ���u�+�����J�;}���u��^a���A>��dW�����۴e�9C�t媜�pzf�|�#alÒ�:=ݙ�9"3�ԹѺl�;/�����+Vn�v�txli�
����]�uf5P��AK�h��Hu�O�]wEk�����FL@�����-Y}���]�υCC^؍���<�+�D����J�`�\�O��{0D|:��퍳�pKx�x�`��k4��?5ƕZ�lb�ܼ:�7;%�U�Oh��1.���*wK�c-rk��E�qnR�t[�dё�m�9��P�[mC�+<B���q�ư�p�6-rm���D�F�Lm��uN*ed�*�"�)A(�$��턑QDHIV��k�f��F�Id\�De���`W���\�MO*���N����9Z�Q�&\ɕ�]���-�h�q�C�P��Uʱ�u����WE��VeQ9]�e^ٌ8ax���	�)�؜St��$��NxTu��L���du$�駕jQ"qf�-bE!I�T� ��Q]ԪQ$��v��$�Z���**�e�Td!��u�hg=�]����(j6�uMIm�(4$B����ȫe��Q\��d%U�yU�%$
�RMN.�EjT':eKY]m6+��浞�#]ڍ-�b$e>J����aK�P�wn����)��^bz 禯5=�Ӳ����un6�Vԉgi��|f��7�"Wv]�=��*�����3]�;�L阮_����MՉ�n��>�H�|s}!��j�}���g��,�xa�Ѕ��\f>�p�k��[��|�r����C"���ϫޤ&�޴4g���;�w�iW������;N.���8N��6[��3ˌ_��e@��@p�#	^S���5����;c����.�0��{�6��_W����W����n��" 5Bx���z���|}��Cz���Z���,!�Mџ,[>���}c��d�<l2z!�ՠ\O������d4l��1/��n�㵊�X1�8������F����W�7ޤ����}�@u�9�)�3��3/�ʜ׈�f�8�E�T���-
�EK��7�_���G���+��_?z��d@uC.:}�&��*N׎��k��1辅�䃡~���d�86)mxU���q�������}�Q{e�����=iO��xC�bҮ�����܌��<K��_�kC��i�qI���ǯ��G�/W�Fk��ktX�Ej��'�]@ڷ)�{�yՂ��eN�O�ݳ0�BwL;�����u��j� �����ŕ�0����W�I�74����;�F2�1G�K"n�](t�je?ϻ`�Ǌ����5�O¥����@|y�Gp:�	sOD_gpP>2�r�6Y��N�Қ��n�u����yK��ד����֫�v��)Ĭ�@P�ݗ/��gn�v^���`Z{;-N[w���Iz_���+�i�ʑ����3A�s�:d��{b��=j����w�j�I!� �E�;"�:~���TsS�{θ,�>�/T䞻���L�5z�{s�kU���/؛�>\}�l��GL��O���/K��l{.=��+��^��/�`�h� M�o�N�������͇$���@�n5��>�~���#ޟx����<�!�b;w^2�EV_�}�LޮJ�q�>�$Q�0G��R�uץ�74'��G�;��cr7��^u�z�޹����4̅8^6�^z3������C<IUX
D���[S������.[��[�3o'�w�Ӌ��r��~J��q�'Mǽ~��@�>5����u��A+�f|CD���W����TY��y��~���C��=��p�n=��u�&�̗4��$灆��3�Я7�G��w�g��o���u�1���>���>����{�{��_���d��©-H��أ����Ȟu��߈�M�xUԴtn��ƴj6�W�7��O���s`?��$U������q���F��qX}Rgx�lE��w
 ��v}�VmERn���΃���G���9Y��q�.����t�{D����뾹f[*_M��nA�mu��y�NޑVI���Vu[�-�2q֧ {���j�QR@�qNF�����_�)Wd��ب�O3B�+M^�|n9z�z��wF-y���z}����}jm�(iUd𧻓OzY�2O������>�-m�ȧ>�W�Lu�+�d7��Ti�uޡ��9Ρ���������/�� ��+bL>��aw���7���J�4k�0>]�˱}�{�UK=����9�CƯ��U�=8��a]̋϶Y;P�7fDVW��kΨ�^�i���vjh�v�\�����n;m_�:���>�/��'��jY�Ł��0���/߰�;j~�>����k�����R%�f\
��ǈ+Œ�ϙY�K#��ә3�g\��"Mb�DϳW��9�2�σ��GE�����l�\iw�n����׼{>v�;�Yz=5�bf�����kw���cز�����H/>x�qS>F�^Dq�z=^(�G����	�Μ����5�V���n����/���,��b0�̳�x����KS)����^E��!؞�0fϲ��V�I�}��!��ǲB�|�l{�|�)�.K4�U� yL9��`����,g��Y�Ɠ�,v��hZuhs�
������{}4gZ��]�N�Ҿ��R�j��㫶�#����}W.���N�]wea�t/4sK0k��\y*������W��oeK ��i)�(��q������q��xJj�*s�f7Q���0\s��w9{�ٷ=GO��\M�w�8�#�{"7��~�R6��@�[ R�K�?J0X�GF�>��7o���犸��Xh�E?+�>�$G�����þ���mתٛ�̂�>�:�=�u��g���EEog����2��:�l��@Rѿ��C�%��1�}M���{I���q=���a;�v'�1��su.��d{�>=$��Q%54%���
|��\�MW���ύD����6�r�Y�J��ZT֓�����Q5Ϥ��&azY��}^�tZ٫�Tǯ��:@��A�c&q��\qK�|��?|��P�� �)d�!񿏲���ñEx�s>�Ǽ��%�\R9��Ǿ~uto羠[��>�fhe��ېiO�T�Q�c�-�aL�W��'��ǝ�ݧ�\���>��YP���v�>��7�b��,Z>ɜ���MTz�H*o����J��]�c�g�t��������O��q�j���k�c!{�K��z�_�^��O�� F ��������Q�}��ΒǣuNQ�u*�N�j�ny�xgΩ�<��^�q�!ΗN�r@~�E\u�����)M�ر�Ci���	WG�6�;�H`�e�?�\�QS��g���Bku+��p��˒�zK65(͹G���G��;oU�U��e��À3�؄j�S��Q��r���v��2���n5u�)�yqW�U��l�+mR�3��f��{��ߪ��S.��+��̟^��_��Jv�טYi�Q���)ה`>�N��T�+�q@�gj\.�������]!�_�PZ���ş������C���R3�@oI}*�;骼���ܑ�/�ij��_�:�/����<��:ʑ�sĞ5%x�U=�3D��zS�\>����a�G��l��Ʒw#���r7�<^����S��u���-�d�s���pv:r�;�;;�lz��z���w3�Pȵt|n)��7���GzG��!�^�p�=5�>�W��T��ܛ^�qA=y����g�����PnPȵt�r��Bn'޴4dyﭣ�N��w�FCO�$)��r�V�{��~1��>5
���[�"�^S��R¸��C�D����=LJ�b\.���g�^��	Wq6���}^��fK4���	�bbW����ۈ�7tr�ko�>���ʞ]�ӫ��wr�2�H�dNK�� >�\K�3隄d4l��_O���Mp
���6�:�֥_��W��q�n;��m�j�F߽Hg���� :����<��E/~>��lz!X�uj=�7�wm�пo'e1fǮȫi�!ǻi�ѽ�:L����бe�
6�4 S����az>|ṽ2v�#���W���i�#{+q]7|�)��V�B�q��CK�<K����ᇉ�ӲBW]���n 2��}��Y��`����UmM��h��R��/uǳ�y�Ѹ{+�ѷ�P��e�O�d�o@U��諏I8	���z	��ǧF�8������v�U��o�h��D���l��;y��+������l�i���p�qD���F·�>ӢS�'z;��_mޏ���Ⱦ����e����}4��~���K?>ͱ�˳g��@��6j�W:�;��W��K�sU���8=9xs"Q*��fe�J��D:��>n��/b<��G<���̩)�;��xj�C��»>����H52�63����g�I�q� Wэ�"�z��'k����ȏ>�/T䞸��(m�2��㺦�+���N�+�$*�н���9P9�>��4��M���w���<�+�����S�xvQa���v�r�T\�/4�ę�L�t&|:�Z���P.o��4�t��tZr��+>���+���϶;y�ɜ���׹}���7���z��& �R�����.r۫q����;��c}��W��� �
Ř'��'5~�<�mG�٫���i�$�X�)*��9j���o8eޯU߫&�M��])M�1%�&��϶�U��{(�ug�)}+�9�k���k��u<��J)��6~5ݵ��f3Y�xY蘙�23��<�Zj:�ւ��Ū�Mx81��1V]:�+��n����Y���9լt
�(,ǝQ��Q���i^o%���=�ix��<��HN��޿\z(����A�p&u���VvD��3q~�ۣ����%��O���^G��z�q7��H���v���H�> r �n{y�W���8��%l����]{��̫�x�y֍G\C~����>�~�����|�O�<e�K��:ܩ�B��jK|k$q#��Ru/��χK񿵣Q���Q�~�"|r�<O�:�)�C,F���zs���$z�rvA0��V
�}=�B�Ҵ���㗪G��Wtb�y��e�uM������ob���[U쀷�j2+�a�Pd��&\	�����K>�]�Lu��í�3Fj�>s5'����Gz}Cќ�z��ޟ=q�B�;�R}��z�L.�;��w�������K�"�}:�_h�=���d'U�r!��x�zh9���2�f�Nl@8�ݘ}YF[���9��/��7�h�Cq�NDk�x�m���uU�'>���^s��u���rN\t�:�f��{�9ヶ��^�>=,+���u3�J9���F/;�W�%C��+�u�#���=5�����B�~1�@,����8����q���4���#��J�@F����x��l�Z��YK"��pWKu9TՕ�zf�ʎ���#:�����dď
�ST�7��Y˞!u`�H��a�]��]J�#Q�:�>:�[M�pC�9r�ѳ��v���n��ټ��wϳ6�f��?�z5�pJk�~�x���҃�I�;��h��Y3=j�M
���v.��߹^��Ƭ��qgĤ��bI�;\�2�j4���{�x�0H��n�h�|;˩x�T��_C��bᬩf����~ �c"*e#=S�.�^�r�⺺�����^�^�ﴥz27�>gs�u����c�\ܠ�e�ĕQa���P���󣞎��^�o3w�ɞ���px����q-ߴ��9��P�ǵT�����=����9Nn��v2J�v7��s{�׬@� ���F}�Q>��p�s�q��z��둷�z�����~}R|+}53ٞK�O��ā����}KF��C��6a�s����~��:<���D�����k�O_��=��IZ��P�B�GR�:V��b����qֵ�;�wU���!��K�W��|vsļ�:��N�D�\��3�'��K���-l֩c��hvceF��獯H��p����z|���+����� �zl�**_V��^����)���m����v[d�N$rK�ٝ��t6ZZ2��u�yMq��� Ի]p�i��&�K"�V���;n�:j��%z���P�Ֆ#;z���ie=�f�ʵ�V��t�X3��.{�V��juՉ{��$+�5`����2����N&���8 �ףQ[	Z��W��n3���o\{�����{ή��H�?_���f�\w���>%@���lF��͈���Sr+���Y^�~�^�{r��w��{k*D'�_z@�eJ������>ɜ����ۙ�A�2��=������gC��CUO��=�/���Ǳ�׸�|����;�pz�=�<&��j���/|�����ӈ������ꁳ��NQ�qR��;����wez�5�b�e�Z��+����~�?87n�_#w3�N`0���"��d֛���Yi�Y�-u�����9��Զo��ʹ,�3���?]!�_�Pι�4<Os�0���}2��nv��Oz�(�<3��׭5�y�;}�5C��/�E����~�,��e�qeH닞$񯤯����0�"�gy��^�3�o�������y�W��o�x�ȍ�Ǽ�>����7H4��_��/���z}�m.�`�D�=�]Q�S-�_��E����y����H�|s}!�������}���G��>��M�&�<�߾�F�P@�Q��R����j�����Rs�Z3�}mRJܽ�2�W�f�S0ĩmpǋ�6�Q�ʹ�}r�ꩯ+����湝��\Ö�1".���bsVnd���.�ܝ����b+��KfU̓�Ҩ�ۛ�eW2���թb�r�:ݕ�1h��څ�h-�W;�	��[�1+��g�=�N�|tW-)�>����##���g�f��ۥv�8�Y�P@���IJ�ς��R
.�+��]�\.�^[}>�⳯ö=��&����7^�\M�2Y�D@j��<LOҽ]FC��ҳ9(���U�R^��o�vH�q�y�}�D��&��ՠ_���Dۙ��B27��T#q9=�#�FxN�*�^T}W�����~7͚��m_������z� �dX:�)�3�f{K��;��ܽ.2��Wo5��#��O�Z*O�r����{�=�:�)�E���DT0����h�_����e��o$}q����r��i�qOk·e���{p���1�>�W��3�yHr%/���w��P%�6����p�q�*�L5ckC����I���u1�ڬ��MY�}��f ����ز~��v�~��f؆�˳g��@���̟]�Af��N���ŏ�w9/.��
�ծ@����u^�!z��/~�	��i������3*��.&��pMK��.݌m��Q�u�����y�
}/ޒ��TsS��<�нS�z���(mDGC��9u��R��5YF��)�s�Я��|�j�(�a.�˨�v.�K
�|mޜUb�]ս�$hKkw�Xܡ�!Rͺ�Nh�}l�2��JȢE�>�y�6�[��YǙ7�����Kx-Ԏ,��ڍ�i��/)g��e�]m�h>:�/�݋$�B����P)Vd�
sjMg*��@kw�����yU��EԔK�ҭc�A�gl�l_ڏ>��������.�e;����o��\Tyr�pN:�w���S�]k]���2p��*ԫ��us:�����ry`�K"!���M�q�Ѷ�X�[��aҙ�Т\���a��,��h���q�5�Ǭ�i���X(��(�)�q�k���D���o(��r8��쬢q�B�+����Gw���2V�,A�+V-�&d�ʣ^ŝ��{aT"���!�t�� �y�M��5�KD�b��K5v�2�9J��lYMɻ���ah�p�](��w�:U���qW](�lȊ�U=[.#b������(x�<��1�+4����Jw �dG�*�Rʗ�/[Qa;JI�;��N��4T��9�+�c��n�ꡏ��'����ɝ��OV�]����}j�m��r����t�^�U23�'Z���"h�e��[�A� �
���!�,��3y?�ѭ�Nmń(�"�Y8F1a2h	>���Q˸zv�_�gnm.-S��KFmKιx4h�:c�Uu�L�Z�ʷr�Z����fRޒ�{N�L�T�1�z����v-W%^��]��Pf�Ǚ]h�\�T^DcLM��P[zu�,�y�����9丅���p�<�W;�)�ؖ"�$K�ո_ZB�{�jw���\*Vr���[\Mgk��|oU,L���Y�l��p�7�վU��kRɛ>Q�m�G�ݢ^��O1��gVBd�r[��5h��Mޚpͦ`
N�^�]Gf�9��H����&nT.ʝ�v��υU������A����xqAt޻n�=�u��[�a,�i��7+tU}�e���z��fYPLգ���C�V������[�	4��,��M�kB��k�_�	���W�9�Z<�g�����	]��3z�*!F�� +Ē����9ɹ�eX�ztAIV871�V�)aq�/�����0��Wo�sZ�����
�P��A��2�;(i�1�����_#2Qf����ZY�e��ːzW3}`ԡF�u���o0�i��8�,�+���sT퇫��'u֚Wյ�A������w7��D9��;Q�瓕�1��j���� 6�WI�ҏ�u�i����9�2F��gM͘�G\+4I�v��t���l�X��1,������'G��7�ʧB�bwQ������{�o\t�dfGoJ��{�M�����6�������38�t��!�.��)jn�^㥛��WJm�����cډ��j�GT ӫ�zHяB�}o�~:��=�fc�mB���C�\��D�Ÿ4_g;�
̄M�^����z������]K��]���2��Jh�tOh'��B��Gi�fH����*/#6�gZG2�B���ӛI	<�P�86��S5���.(b&���tt�لB����,ل�ͭ�QUtaD{WN�͛WO/#�="f����^^�2�=leT���X��yԈ�yM]��a��(\�-�e�da�j���PF&��$�9I�S�3�����F��Qa�ȼd�P��S$��E(��!�T�$vՌ��WZ�@DW#\��k%��!��DrZT��S.�d!��SD����ɓ	�09P���v�˱���jQ[n6�#�A��\��&(�P��ꘅW�gk�EQ'�a��vQN�m�!p���=�"yy��3�Yɧi�f����'��䭸�Х���\S�]�&HFcP���6�L��F�H��".`��`�5:v�(TO$'�)b&�(���={t�D�L�ڕ;�N�O�_^7J�Wnpξ��+,��%�{#}�k���f,�a�1]�2wo�C���qN������L�����+���_���*|�7W��e�}jߏ���z�SI,�t���I>��xz��$�Lms�\޹���.�7�2�����Ϥ}��X��Rf���oVz7�
k�Ea�n/������b�U!u�^�9mՉ����8;�i�o�G�
�sc%\�Z}�;�;vC;���ǻ>sY�υ�e�$�2��R$TKjs�WP}�S��j�<��ӗ��֞	�޽�y���U�i	�~����.O�}��Á%��ez==3��։��7]�J�ɕ��*���ʢTO����#��\8����m�z퉿��sP��9�^j2pQ���X����`6]�5GZ3���#�8���v���|ϫ<e�����ʙ����y��R^����[�+>���F��~7���M_��C���}9�}TA�1�&v�a�g;���^@{f�#h�zw�3	�U��\�����5j�Ǘ�G����s�Fz�Q�>촰e3G�vϠs�f�#���8�'�L>��1Q-m�ȧ>�W��1� #�1L���kf�M�U2d���+U�v�x�!��Ԅs��������t껮���7aҵvg*�E�����n/���X��(�+��Z�EKP���op�\�r幜�p��W+��]a����)�I���	zAuںH�D^\\�YئW���|��\=�Sp�>z��"�w����=at���[�v�w���2v�w�2�8R�r�8_m��d/Uyޑ�N3�a�NC�U���R2�Y;_���]"*�~��3>��6�j}���7�ZN��5O�n;m_�C��q8�^�w��'�ݹ�������g�+fE��$��G	�>*t)ɝ:Jd�y2�V/;�dC����}GY��KE>�c���;~N�ڏ�d�	��6&X�'�Ϫ}GEԺS�2�W]����e�ǸeyW�d�9֚��Wo-����\wdCw�ƫ���gĥc(�ē�v+�^q�u��y	����&}y�A��=��{v:�5�}��=t��D9�F-��f��'���KS)�,A��a��ݝ�OUߴO~��b��(�D����Q���iN��y�_3ĕPf��3��O=�=�y!.�eMw��Fsǲ�w�龸����r�y�gѾ�������w���~�þ�
�"��G`��� �>��#����=p�Xh�S򸛟z�8}9����4�Ƿ�#o��Q�UE��m�b��2,�!\�i��i��Q�X���S[RG?2�Q��o̷�O��cӅ��I���EXy]|P��ƚ�שb��ޮt��I��ض����UC��ˎ��C}'S�˾��pn�8�u��C��o#gX��� ���΢�Ng�M��g�2�/w%� � (��q�L���r~(fD-֩ϥ��1��ζΥe5�륓�0��ee^+�S�zO�9\O\R��9��*���Q/)��N{�r�z���Wbw�O�(\q�c޻jo�BǊ��ӌ��@�F@�t�&��'��^ߠOa��}^�tZ٬�������zG��٧�nԆ=��E������f� ����T)d�!����hZ�V���-�z��UG�O���ݸ|o���2=�WF��W��8�!����ېj��zVS�Z���v��+Sk�U���z�n��nW#���7��>O�h�Ͻ@z��ۦ+��,^�{ޞ��jE�ܭ��yO�L�l�,���W����"��6���x�wK��W�u5�0���[ƥ.��^��@���_�^��g�?���χ�:���~�U���T�������uaB�x�yh��@�mV��}�c���c.�p�Y;�ü��'�ڗ@y6��K豽�쉫�S�Hy��r߯���{�z���?m!q�*x��)q�xA�^�w�˙����4��`b���5����:�C�JoL��F�����ʶ�i õ�#���\�Km����R�`�'���Ӹ:;������S=3E�B��1�{]K��,��x���y�\b����Û�	SՖg�T.gHm�u�b����˷��Pa�zȽ��z{o���z���-q̹>9 <���G��K����uM=�W�;0�FS7������W���G�܍�Ǽ�>����Yh8� �<o�#ý9�7��_����(}Q>`5Q멖�.+��7�X�7^һ�<_��p[SJ��y̌���)g�;�)��Y �,� r��(�|ܡ�j��Ͻ(J�������U\=Z�wu�U7�G*����'J�������l��%��U@��I�)̀��n�~�2��17�2��g�1��la�u����MǷ����_�%�Y�D�O�]GLs�g����w��+q��1��k$p�O���>�"}�NM���@����d�g~FCG�5�pd�u�.�wk�߈��}^�qE���P�\٨��z������}��P�.�^���x�&j
���3C�gt��8*K��.5K�r�\{�uTT=��h�?z��J�(�_�R�Y3ʹwS����ɓQ�*jO�G��mJӢ��xU���G+ۇ���Xe��޷M��5v	+����N>�u�ӗ�ob㓘��,l�㽵82�إi��KU�O+ܾIk�+���c�}�^�Is�+.����SvC>)9�`V��^�e��-w>:*�Ò�<6_@�_�����(�Vv�r��ft�3x�,k����o����t~�?@���l�q��G�5�kC��86):�{;��O�����,�ܽ�*��<����}�ӛ�v���k2��N`0��;�����K#n�RQ٣������+@
�n�2!�z��z��/~�	,�neH�|Nf�����������^�9CyV�p�J����Z%f��tGD*�?zN��j}�:;�k��9'���:;�}����^�lg��Xj��˙Gk��<�tϠ;���+���_���+"��;��o��a��6�fo{��y�b���q$�̰��3��Tϔ��s�\޹��K����w]�uݬ�5��uU��[��M���#l�2��I�� y2�R]u�sM�	�7�o-[�*�cW"��}]�n�K��Pg��ǻ�xǢ�gY�J�,	�"EA���=�~;S� ��{8n�{��~�ފ��$\��џy�y��'{'��~��������ȁʌÀ�S�l�Lmǣ0ɸ���Z|���O���醊�_���O����#�ӣIQ��Hۏ��lM������~����'�y|�ā��,-	}����}I��Ԓ����v��]ެ��k�_q� V�PL��w-f�6/��K{o�P��v��r鎋t�h\�R�����s�[�Ҥw���TɃzK�th�>�x��ܵ���FEb��x� ��\���Pѿ�Z57�l���x�ޝ������<Lg�;W��#�V�=S��"����'¾����"b'ޤ*��ѹ:_�ƴj6�W�/�ȟsfž�!xW_n+�.'}k ��kąG�Ӧf�*�R�h_��Zj�S�q��#���a�Ӄs�V>�\uz�Ǳy٣�@�/����>�$�Ȳz0����TK[z2��Mw���.��idY�4�O�,�z�wB�{���~�=�q#b;�R}��z�d���a>�<�G/:E��S��;\f�x����p���#��CƮ3�a�N?uX�Y�#/e����׶�^E<�\MZ�;��:����H�Ƨ�N��/����gΪ����x/9�;����np�;c���zƾ�K�|�甗���:v�}�3���Zn	^%��p1y�yC����v>��2�@��G�|�z�����z1�V���n��+��������G�81�1���$�W��p;���d�;p;����֏��{=j�=��b�eO��R�2�W��.*g��9�����S%hܡ��sU�V^�o��y��iT,����n�V�g�ޱ��RE����	��x�}�1�
eb�2Vqy����j�k�m
��8o;J���x]��l�WEh��pW�-W`�KpfP�Q!ώ�mh�� ��&�t��5���_V�9sWI.H����q�cr=���Ͻt��9�F-��f�{L��2����~ב�ȃ`ײ�f���Yi�V�!=M�k�>���A�8��� �������R \�j�J�$[���Ru^jT��x�T;���+-]����뉹n��x�9׾��j�{�~�����Cۗ�'�&�[���K�� SQ'�H�
G�ʬ4e�TJ��z�#��V��#Os��L�%��l*y{ �[璯�;��~3t�>* �&@��n��ॣkT�d�[f��i 'o}�'�G���U��莙�&����׮�d[�,ҩ!���A�hdS���
|��F��c)�l]S�S�ڴ�����A��>��}8�y��F@������3>���5p'��D��Qg�/��x�.uȞ���_�zkzX^�;�����t/:�>����*,��.)d��C�>��Y���c��������^ӑE���P��/u�{�j���V�~������{nA;�׬�9`����^�gg�U�o�||��R��m��ϓ��8����{n���b���۵_�Ⱥ��Y�b�D.K��5�UwW`��Pظo�1m���Ӧ�sO��{����w�h�˰�Y�Rz�T	�����z_d�vއ�-��I�mhΗ'e�2��������j�U�+�ݲ��j���w7���v�!7{�m�Ỻ��R;͓�E�����r��@�0�-�l�wY^t��<r;���������2��u5��?3[���/������{��ٛ:�����>�l�rrN���_���L��v�U��vH��]f�wW>���%�1�j=�Վ����cn�t�ȲwA�y|��d֙�$��=C�g�ν��'@�F7l*��x��^�^�C4����g�܌������!�Z6�����&�-gy�����W���L��O�d^�_�=�~�/U!��e�p�T�3�tug�i1��%X�^|���D�g�z����o��p7���������H�{��yN}�u��o^$3����O�3�����UB����50�*e������t�X��7~��/�_�5ѡh�'U����|,�Fk�]������C�*�2��P7 ��C>�t�gޔ&�zd)��uٿ]W���ƫ�jKk�A.�~GȜ<�����U3(�W��� ��E���%��G�� ��e���>�l>�4� �!����&����>�TN�%�D@j��1�U�?߿T}v����Y0]�f]���j��j�]84��L�'���+u���j�oV2 {ñ�j�	0�ZwR�E�v����-^�F��+�Hv��7Pc�//���}K�A��c��g]��2pY�1g�uL�S��}\!�|0���s�k��w&t��Y��`IU׺�袼^�Ly�k$pOΘgޤO�zp2_�8O��9�L�Ix�v�7�e����^M{��H�O�J��.r3n��l�m�j�E�ҁ�� 7�`x�����V/ʭ��;�՟�?�)i`�f{�ʜ���qR�v���㗺���U^6�W��j�)��������� ���C.>�Y2j�*h��=8=u+N�{>۴��ܯnF�:Urtoѕ�gf�)+H�z��oD�>�ˁ=?^���3gx��P2a�����O�踤����q�^��;+���zC�Ѫ�G���!��w���h�{z,_�2����a=�Ni��3F�X��gӕ�z�����{U��u��}Z�z��/�hw[Hm�ȼS�wr��ǱU�7lѪ*��B��+*:rgN�S>D��LQ��"�z��&}1��G���>�=نf^�y�_�M����n��Q~� 8[��#���>u��T/K���.�7�S;��4xk��&�ٌ�G�_ګ\�_/E�wm�����}5u�����M/ܪ|����4����G�W��;@c>��꥿p����+&�Cv�[q�9��ʓ:`n����YH�䚴q�V��T�gB�k Pͨql�)�|"�Bm���	kٳr�KU[�����1�s(�%��V�7�M��f���vS����+Hۊ�혦���2f(�]���^��)F�d���b�#�|�W�Ͻn���#p��,���A�2��ȱu*��������-{�${�H4�i�Nν��/p�n���#�z���Pg��G�C���|.K5�%W�X$d�2��q�/.M��^��ژ;-މ�[������+|��W����7����D�� j�/jEF�1Ц�ܩ���*� j*�L{��~W}�h\���:4�{}R6�v���n�\z���ǉޚ2�9{��O�4�� W�끸�_f@U�Z5ߩ���w��|rp�ϩG�Ùo;���*� =Ո���,)'�=$�P�/����n5�Q�	����D�Ǉ9��zP+vk�KG�����x�l�4��\�a{B��h_��Zj�S�}@����ʋ=���e9�z�\Bo�h���7ɚ��>�$�"��0��O��DK[z3v��\v+��"}~\�`�q�oRs���7���M���	��ȡ]��|OW�&T>����R����S��U^$�z��z���Y|_$�Å�m��dB�W��}�5��vz��Z̩���3ޥ�}}yA#���<%t�P�24L��\Jܔ���0��qlb�sJ<�e��p�ܢ��y_S���X�8V��V�T�=��v�$.����[���J���nQ%�}�r�����v�fuGN]/�1W�mai����]Z2� ���+9�`�6�Uo!tQ�����T������)�Oٴ��xƱG�d�V(,X*��G:k�-�ԧ]gWRpb��tߒ}j[h{N*Wqu9��ǭ�R���őɎ�E�[Z�m�����]ҳ,r����!A���9�0B�,*=��]*V[�������,XK��s��1��NQZ��P2/E�F��|RF�R�U�g��Cub�m�ް�Jghj��.�úc�4sO�9f��RSj��``�v
��r�'S�������X���mfv�P5	I�7)Ѯ2�rK�IR\�]mʽ�2�u��Y�S��)J�S5�6s�ʙ[�v.-�`������H�mB�W������ͩwM�ˮ8���,*�V��Z#a�G.��ҟd�t9Y/��W}V�_�z=��Q��\J-�%�r<-�	!x�-�Y�O6��9x��Y��tH�AT�F]��Du��`�h��"�3[�1�0ܹ=��ʎ���z�c<uU�e�[+:�a�Y�MT�?�0����fJx%�`�Ǌ�i\C�e��)��Y	�ڟъ}Yz����DS(���u<�ok����OH��b X�P����1�
ͱVK���R榴�9��i5�/t,�p�@�����Ҙ�m��7GU�:��=����3��߄�'���<��)�;�K�)�������83�pq�}7K�D]��F^�6�����v��{�%l�n�a�ai[�m��\�1Й͊���.�Yn����*�>t�^��XE�%{Pͻ��-�������]YS.	::�ɮ}z�L��6J�Q�	�UҲ�ž���sR��zjC����<r�\�\r�Y�⯙�Ȼ6)�Q1'̛�n�մ����K
M_P=�v��r|�f������僰$Ѿ���L���؋Υnfd��Ӑ�K�F�����5�ٯOt�6�k��)K:�-�J��]|�Tڛ9Hbm�N������Z]�d��ҳxjgJ�17C`'�k�rR������K�����+��|oK��Q��K�V�Q�YK�i(JW�7s��Yw4���㝻3f]�s-��2��R_Nu��u�p͙�FN�Cr�J/��o��]&��5�#|�G�۴�����^w1�Z�G�*ɴ��l��-��ėۘ3H�Q<��Z�\ۭ����W�qJ�������
⺯��+�oN�v�Z�:�S��rG"���@��a��q6���z���X2<۠��/�F�p!��ܒj�b�Pi��vl�B�*M��h)	y�r�͕j�͖:�%=���JԊK6�䇯�N|	�,ʌ��v����ʒ���YF���x���Z��J�v���Z�4��a�E5ָ�aK�]=�ܮ�s��ر���H��i^.\��E���ذ-��-̊� ��cʼ�6dZ�B�4���7H�,7*�CCUЄ[jQd��ii��F�X�44ªHҌ�d2�*��ĎfE������[0��0����I�P{T�d#�ď#<H�4�L��d�k:��s�K�;H�y&��i�l*�R�c�4Z��Re�h3�3�U���N��IJ�l�"F63Y2ݭ�'���9�.s���6���h��ss�'!bXW���G9{P��g
�y� �.���G�0��\�k���%���XB�J�񆩺.�L�gT�a閊QYY)HE��1N�t�^���=�l$U��JK[�;E���#����6�6��X�N�����R�3L�%Nj-t����Z�(��^F�Ξ�l��粊�sJMg�Z&dT����b($�$w�黾߱S��q�U�j��Md�;��7w2����iHwwG��C��֤%����=���T [��p4���Az1�����m\���L/�Ee$o�S�'N��w+��Ϊ����x/9߼�y�bt{Ӟ����odf��U[�.�ɿl�t��}�K���ʮ2J�(�̸�������N=@��=�v}O+/�Ϭz��o�p�7|��̙�k�t�̱�O�T�������%��Vl�8����W���~����>>��g������Y��Օ<nωJ̱��b�gȺ��ir��s��׍�Է�<8�:�#=�1�l����Y��a��f��w��?��xؚ觕�@g��^FmyTϑ���HO�-��8�ף7�>gw���A��:�A�,�����zc�z="M���˒��_��z��:�ϼU*�>=�7�[�a��s����|oڪF�����S����_<�*mb���p(��zjKCu��\yU��G���&�޴�Nx�2����+�x����ū�_�]�ۥV̲AgaAQ z�u��/��Z+Z�:2���Q��&���4=����U��Y���O{޸����~2%��RCW����ȧ=㻅 }>3h}����2�R��C�c�V5�4��z�e�.�;&^���#ot�Ή��R�U]4�M�:r�X�np�3r�m�蕝t��	��Mh��zz��L�2�4c�rs���r�����;o�8��v,<T�3[���0� ��7�N%Ss�*W.Ѯ��Gw\�mW�����d����~���n�IPL5�{5'5v�'�xO�iJ��Q�Q^٫�}Lz����p���\/:�>Ϡz|�>f� �����ؒ�KǬx�n��B��׸^D�ޝÿQ����C����~����?_����>��z1�Eoe��x��{�'� �\F�~�[�h�>�)|o��ۇ�����ޠ=E�}�Nl��3N+.��^��<ݺ�ߣ���Pr|����6�S�x�wK��q�̢��nE�C ��>�}}~�c�ܢ���UA�~��ţ6}�����~��l�w�NQ�T��N���>���fGeEw����!���d �_��U��?i���8Qin0xx������=l�3�w�� f�Q��;���Q�/}�����
���~�W�VG���8���Ƭ��qgĥ���'�u�z��ν��n�eL��W*�#�P�y�޲.7����W��Ez��X�mF��魚�5[����"��%�}'�k�*���3��,�uP�q�{NF�G���\{�i� ����߉ԫu������ �p빯z�5�L��Z��5Ì�ы`�U�9c��>��=P5(g��X�6�K�p�XͫȬj��x]١å-��$m/�eu�Srv^�R�����Gq��ˁ�1�2p� p-�=Ցh�����at�&w9�j��~��}|�|��u�^|?s�O�^�O[<e>�bn<�������<*}�V�wq��=W�=5�>�@��8 r�,	
P4��2��񸊖�h���a\�׏q{�'6�ho=O��HҮ=������0��f�A�A�=0}$K���/3°=ܶ<����i*�&�}J}�CB�y���ƨ���&����u����3%��D��\��.I���&�4�N�f�Y1�ޯQ���{��G��r4r~v����=87�z���{"\pW����軙�=7�ϒ�a���I>�tn(�;W�p�o�l�m�ڿQ���ԁ�W��Q�w9F����WW�*�ѵHٿL���#c��բ��~;F�K�q��q��=�wG6�V<�d+*<�vZX�4}���9�{�O�d��a�4rX���+��ׅ\F�>8�^�؎���Q����T�q�|�ь�ފ�ip'y�������Į�d�Q���O���Tq
�ӳ&�۩^W=%{�0��G�|�^Y�#�.#}4���a]���҉ݳ0��X�T�L��=�b����QwuY����'��!�Mꂱ�a�8�O�~�W��%����Q�#�X������UՉy0��9��g<"�皰��]�o���X�)�<�f���έmχ+�ed�}q���%sԆa�[��w��W����Ԫ�w5[ V��c���+����)��_d��ۙR3�6G{ļu@z��3}ܒ��xe�|W��Ui����V�`�17d\*�?zN�^���s��Gg Ӏ�ja���>�^��!���.�咆����z�_��g���TtϠ=��W�ջ��`Ё}u3�Mo���M�~���oq�F��ꚉ:�K����z4�r��@�mg��Sj��$��D�ZzU�rڿ }��>Ӑ�>�Y�wL͢�Y�\_I��A�,\T�B�b�vo��q�/mw�������bo[�ޏS����_���ݐ��=K;�%Q��[���nj��GE��k*}zHm�ө��+� ����k̯)8y}�'O�^��r|r'v �s%EC�n���o�f	<뉲}��h޿+�>��W�����q7���#|ϳ���;�[�2�;�����&O�� 54Hu��|}|CF�Z57�l���W�����v��u^��r���x���<�>�>�(�!|���q��F���kF�V��b�ȩ1&_Q���9{��Y�l�1�nL]�+��U�ރi�;w4�2�HIV{w"Cv-���V�����}�^��1�h�����l v�Zn�X�Gc�����S�ΡJ��c��gV\�{-�2�rt�c��n��� �ֺ��>Jީ����}L���:8OL3���K����7�|��e�1\�鿌�/_�V
��=�B�ҴӓB�ULwdS�>+��i�#������]ы^~�F�ޟ@�dQ�]>�$����d��>�5�-z�A�VV�ƥ�6j��ۢ~w����Ɩ���U:�C�~��p��M�O���ީ�p�����g�i#�U�����	�c��n�E��wW���v�߆D/Uy}�5q��z_�h'a�9���+=����7ސ��������v��O��K�t�/��vڿ�U^�qz���v�5����m�j'Z$3'3?VyD]���,���v�/���wYU��W�G#f\^u���%=^x�W�9��_�O���Y��K#��s:�Êe��3�]O�踩t<���t
�W>^���C�����`���g�ڸ��z���s<hx��X����q~����M�gs�-#�T8��3A��3��C��z<w��/f�kܷ<	2Q�.�)��T:�o:�nA��$���]1>ȶ��>�`_o�|����}?[��)���_������\on����sG>�\�%b���W�(KW�5�]4Z��c�bO�)�Л�[��,�z����:��$՚IB�����=��+{�q3�}����cJ;�^M�k��4;��k�tjh�7��ۜa[)tƵ��X�:0 ���ww��8 �W�YJ��-��Z���t�\Mķ~Ӑ�#�{} =!Le��56�쵞,��2�3Z�Y���d�� SRX��)���&�޴�]��8�a�;66k}�pnγ����g}^�fY ��)D�����|�m��^���M�q�^���m��>ζ��gt�������^��p�K5�!�DLI^SB�=��X��F��\���JU߻���w�W#�U�Ã�+>8}8�x=Q�+޿\M�3�*�0�v&g<a��L]�dNz�r�����FCY5�TǮ#��ʪGD/:�>��_3q�T?e�΃~N⧶ޒo wwy2L���/*�w��Rݸ|o�����]���?W���������{y	��̧|�{�vT���D��p>#M����;E���R���T>���v����̎�©	MGe.��ϴ_��;�,V���z�oc���Pr|��w�Z���[��~���6#x�I�u]./��k��7����Pu{��fl�㓄�~����(�ɻ?���	�{j�����Ծ��޵�����c[��y!v�k��s�?�T����8�Z!��Ŕz�=�Y�|+cV����L+���4^uM�`���uR�}#*��N�P8w�4oS��],�H��\}�z�˷���
��j��Jd�
���][�%{� 7��PꟲD:�G���_#��:nd�٘x+=�>��z��h�����W�E�R�f⧨�4׀���.y�<�z��R�i�~�B�VT�Y�zL����f�@�g�K�NW���_�C�2��z�o8��ޢF�_�=���������_��
g��k�|Q�֕�y�geHwsĞ5���*a�Q�#u��o[�����+}#��-8&�Mٜ�T��6��nDҟ+t�d:�A�	���I�T��_P�ν>i{ʥ=l�J�O�Vׇ����S��'���}�!q���:�k�Mo��� [XJ�7(U�Az�|Fo��j�ݖ�3�(In�`k.>��*���ۊ��0�gb9�y3�][���*==�5��:H�A9�9,%�hp�����}�lv��w{}q:o�_�&�,�U�����*L�E{��^2�'����]FB��oZ�:�2�H�`��d�ޜ���lLQ.x��S�w���M��>�!#g�����2����5گQOޤ��ͻجYxL�et��cp`�����Sfcw�v� DUtڰ��Mؼ5���u��ܬLobej��8U�7��t��qв���+7�!M]=y# H�v�o��fDq\N�)�V�}�[m�	�o'FHmM��W+�VN�s�Tל�U��C�CN]u���z��*z [6�:��қ�� K�ߊ���U�K��7�_�^�<8mCf�ڏ��T���\uz���S�M��@w�:���O�dҘeM�:<lzJÃ��ׅW�0^��j�I�F��;Z=(�5^�{>��]���^�~�p'��(�����8��C&���oүe�p����^���֯�&�Y;�����mޏ����}��{�v���p�*p�D�%=/:��>�]���{�<�t�=>�r5_���~gՠ��yz^�Մ�G��R=�55h��4���W��ѳ�wl�{jc��Zn*e���i�*17dZ�S��Ϧ5�����m����|?m����o��#�Z�$�ܲPۙxh�T+�U#WK��r:g��O�㣟��D�O���	�jZ=h�z;.���:V��~��g+GD��:����KG�S�1q\�9�W	Sh�u(���<��T�ER�sG�*Ԅ{
e�����,��b,+2�E��z��A�,cvvr�F�/<0x�e)�X��<��mҞ�����k��p��G����Pg��ǻ�xǗ�pxo�ё��7���F��k2�����t�5��6��H���P�+3xA�:remv@�� ��J=�Jol70R=v4��*�ܾ݉��� 9Σ� �w�܎���t�����7����S�q��[�:��yW1��k��C��,w�ɥUչܕ;�q 3�OE��>��o8H�oף#�k̭�ʎ�G���7�����Y��U�^:�������ф@ޣ0�Oź�l���h޿+���yb�>G_�F��{��H���N=�rv�����U�Gz�퉸��@M�7\���2�h�Fc9�[g��Q7�A��p[�o�q�v{��v��Z�ߌ���,T*�Ԏ$dK�!W�K�s���D޹�i�tI�+c*{^�N��{�]G���O�|}9�}�`�d�W.zn�/XU���=�A���P��UR&���j��5�����G����4o�z}�b�c��d��E�ц	\�\P�qu#���^�1�^�NV��ݯ��w����wB��������y;�2�&3�L�ۗ�.v�ykD�q��|'tÕ;�b��>Z��p������#���<j��Vt�X��1�ȼ�EY�A���E���-�G��a_���P�������/���~�Ϊ���@���􍻭��K�=�}WQ=o�8;7&������N�93�I^&���_9z{�v5��t��"^,��[�.�UWH`E�6#�U<�F%�ζ�l�GQ"�3-k��N#���rͷa�2cs\����KHe�ᱚe�p��zK쥝a�X����J7�m�x-9��I��jYǲ�Jʎ����%:tyM[��52���P�]�4L���u��]\�3��i3���VG���;�t]���^��ne��<�>�������
6�]��u�d�� �K�Γ,R��]Q����cU���>%+�,e�"*��������6739�'هD������Ȏ3C�>���"���c}���z���9�F/沥���4���]q}�=�o;ܗ��^3�O	%#�]tļ�o,C��V��'���@z���qKī{���˘�=7h���o����F�$��3�*�qFX�w�[��n��>^��=��!ɨv�v��ݝ�[�>�Fk�p�߇�Q/a���I`L�@)����F_�D����d����6�i���䧜�o��u��U�,�Y�PGH��p�C^GL�q�:��[���gЗS}�l�>ζ����o�{��^��p�K5�!��u��S��gz��N�"�{3����������\���W��A������Kχ�2G�~�����}���}Fc��h�Ի�m�'��D�]F�[5q���F�r��楒�r��1@~�����BO�HI?�@!	%�~� BO�@BI�BI?Y !	'�����BO� !$�$ �$�!$��BM BO�@BI��I?9 !	'� !$�d �$��@BI��������)������Y��0(���1"����M))Um�@TPP��Ek_F�vjI-��ET�R�%U1:��!;��D������j���EmI Sm*H���7v�]�l�h��]Z�̪���n�\��U��Q{{�{��/X5�ce,���5kݥ�e������U�����imU��komu����];�#�n��{Ưq�:�3c[��!&i�+5�M�ݭ��+i��6�f�ӻS���mӻcV��Ά����Sjh�]��l�e��n�m���s��M��V��Mi랖�v.�[� w��5���g_/m���Ʈ]{�y��+Zn/]U���ʹ�N�X�O]�^u� hyλu�\3s8uA�]�7]�iM�V�-��o]�si�WL�fV���[�v�k�� ��Y+�]�ͺxm�+==r�yv�^z�u�
(���� ���������� x}{�E z4QE��GE�ѣ�}�@������ (�E7^,�[�w�	��[���M�  ��|�E|�ۻo��g{n�U�3�{��C�z��v�ʭ�������{iCU�^�kʊUL�]=�6�s��l��Y�F6��4K[b�g�  ;���h鮡�s�F{V�sӽSCme޻��ݯZ޺�^���R���w�=C��W��[`�{U��^: Sޥ�vcl�v�٫�z�����l٥���ezwv�l��n��   >�>�}4����wi���h:u֌�)@h��{oY��:3��V�lWo^����γ�.����n�U�{8�5^��NuC�A��{�f�i�jE���H��ҵ��� ���֞�R��k�oo]
it�ܡ���ב�3]�s���luTѡ0��y�n��'�:����ލƯ`�w5�=w�R��3��ǽ�����x��R�-��������؝��� �����)u��h�h����{��[�v:nÞ�S��ݻu'�ҽ5�Z��ڵε�4�wG����Q�e �iՏuo7 6��c�����Rz7X�մ��m�l���r�   ����n��,��+�3�mǡKV��{oP6�����'��@{r��t�n��Q�KM���{v������z��۸��{hk���[ё��k�m�]ۺm�G>   9ϊ /������Kj��t�xX��{uݩ��m\�N��hl�����]�9�]]�˙���m{��^�m���k�m�@]���ܵàu�m�nPK�X�l�n�]�T�fɮ��  ���|������SoT��֎����G�v������x�֕�d�ŻP(�t;nWJ��E�kˀ�:���ѮTͶ����Jts�T��̪J�2�E=�	)EBa2�5OOL�UI@ �JUC@` T����*���� 	4�=UM* 4x������������n�p�o9�]/��<1�=S������~�u�}�^��BH@�s_�!$ I0�		섐�$��	!I�ID�		���}����W�����DP�^Z�Z4���8�܂gڙͽ�$9J���/�#,`8�inb��Yt�*v��l��J �����WN�Ř�=�C4jYڻnR[j�L������h����9M
I�v��'�YH���eĩ�E�h�m�ںٟ
Q��w�N�K�٦�$>�|��<�lȼ�0���*]8 �Yz���Q|(�(;t�Ի�S�Z?�d���çl#q�_�U�n0f¡ˣ�h0���%�Ż�M���`+Z�,�V����]3n�S �&�߈9{��� nX�������.S;��2��[,%�5n�uv^��z��f
W��%!�hmi�i�4�Ŵmmï�6o�!�km�� ��ۥI�p��-<������(н�l�̙d�-�D���d�x�oj)$˛m	�@�ب�
d�f�T*n$�y��3a,8��~ͫ��J�w�-�x�5��Wu�씈b�I[{y��E=lbI��X�29#��i1[�Z0�PQ�z�Z�q�Yc�e�!���M�Ebִ^:wN+/�Ѭ���\����A�bm��-�#un��ř�p4s`\f'�¢�ɺ�e���~ԀD!(����ŉQy4�WJ:���ٓ-Պm�.az�,3Kdj�nr۩�p 7-Cz.eب�!������C�c{C+&�u`�W�Ih���
�@J_e͕��n!�^�M]�мF����?dQ�t���ׯDiٲe@*��1�l�l�Ac[q]3��/s�p+(̙WY�-�lcY�Xh�d֥p��$:v	�^�T���(˂�"�RTTl*�h*W�:b�AR^9&z��[�[�<���i��8s.��*n��f�e�Zq��3	�0��d
��;�S�|�I��ͬv@����)�1=D�<�Ӯ�bZ�֭9v��6Z��!5���ZZ�(Gf��lљ���k"���v��ʳ�Jj�n7MQ�Y��^��BŁwOb�͖���7x̵X��Y��o6T�
lݭ�n�Jj���d1'�IxᎱ`9��Z ̇j@%��
��f0�%X����iJ`&�Ы���P�Z��g� q�Gq��.�z4�3���@N��		k�K݋{��v�u�!�����6���x-�^��TC����M�AKE����7�3I�W����ؖ��⌌Y֝π���rdW���H�Ч��TnlL�{��n���e1�cCH]���Ep��^ն�?�i�k��g�-V��]��#�M�Uwa�nȒ��	�"M�,튀սZ�����Wx�¤�/�IR�J�mG�!��<W$�a:��@������8�AJf�v��e��V�A�ĵA"2��!��P�%�"0��J��&2n��O+	U5��uv.�ŉe3D�înT�L����%���[(�X-�r=�A�-f�/L�����/(ڱV�Ud��ZG@�`9q�YF�
�Z�A��ևe
�U�n]�xPt���{\ٙ���;ԘI�}�D@���K��G�nQXO�ú(]R�U
&�bR�
�wX/>�Xk �kE[i�;����lPє)��dǢ�КH�`��!��܎���F���ѱ���c=���\1y�	�2H�D�N�!GM�bQosU���*��X�j�AJ^*|�&��S4�N��[.5�w>���t�=�n�ުEFe� ��m�!*�^������U(�R\�:�� �&�.ic�JH������z�|�M�1����7�q� #lB2�t���F�7��h3f���+.�B�6�:(��m�l��'���o�l�b��YOt�v���CY��Qˠ5; ��{C%d�iܽ�2R��	��ʊJ9jV�^*ݙ���R�݁�N]/��F�Z-*R8�fIMecM�b�hk�l��"U���ؽu/m��Z�f���̼)�O*�vm0p�Je*�D'�ŗbir�c0���,��f�� 4�69gMYdB�Lm�W���^�kj0��Ն��̚V�W�Y�������2�,�9�o��;�އwѭ
*��;Zk+ma9��;Aeդbd0oBU*�f��K�r�X웢,fk��%�e,f��	��Q���Yv�ٲ�mF���ѕ�س�F6�m;b�Cu�;�+�v�V�tH��Mk��t��]�x�Z6�Wf��C-*�A^��Y�ޒ.�1B�ՠ-�T�A���M�a��3N��rY4���ꭲ�k�Y�Y����QH/�������k���&���JТ&�d(��8���i�Kq�zN�Y��wq$��ݲMy�%(��	5[�x���f�r^����w40�89j_�a�͐�/�c�%}z��۸~�܀O��JI��n嶃�ůf]1���j�,���)˕
�h���,,��%ȥ��ͽ�6Y�x&\��n.1f��ǯ��:ߎ���(�9B#Wp�Iڹ�m[j�Eֱ��\.�WI�Z�7N��e����)B�]D+)�3pI�=������暱�%�7�E��]���:Lvxh$L��ӂ��ǰ�c��qc9�x�k{G]��(�#W�2b-�z�6F�_b}g~Wtg	СQk���[R�(��$�q�Elv��0 ���	g�,z�5)z��sPU��F;�i�_;�kr�Ik�Mn�(	+6b�A��*��]��jE��ǖkYp��T��IFjma��QwZ�mf����ޣ�-�a��H%7��N��1ޝ���5m"T�:sEa�����;jz��]r�z0M#"��!�H9NdÂ�.X-�hn�`P�R��,�"T�fMá�S���&0�v��x��r�]��T��{`P��(�fLzų��w��j�X�c��տ���[u�2�Ђ�lV���t^#��[�`�@�A���jLu���K�"��d�Pv$�0��)n�;�ml(T�NX�W-f�/���q5������t/�ܗ�#�M�����r�����'&k$3cY�T�3���V�c��m�7cf�Ku���4m-�Q��
`�W�m�����3Tkl�yXf"��%A�Ս���d0�T3md�uN��9,�dަ�����R[V0���+��q* 8&e��K���R��y���B���3H���WhT�K���H-	Y6waĄ,G�^X:h���Bi葤fXLV��*�ϭ�/krZmd��(��Kaь�����m3�$�@j�`4��Ye hL�f�L�1��Y2Z�uiU��*J�իm�������Y[A�m�D8���Õn�(�j�]̰���@���kW�^]e ��Z�Da��(�,6��x����b�()����Z���A�-��Z�)�EPfL�L;8!�{G`7rK�,��٨�"��A���5f-t�˘#d�l���V��"�p�Q�sN�Y����l[>����eV��j[WZ7�֎�S	5y����;�k����,�0ᔰ��`wi�n��Q�ٲ1�B�3v��֋f�KE���Qܬ�Zh�ۧ��L�U���#x�ĭ��T�!n�����=�j�:��N���XR�|3Yn��W�yg%��n*,��lU�h�L��	�[.��<j���;�6�3�[C�e�p'����<nw-!p���qY�ał��n�X�Ӽ��2�u�yz�k��1Q���0:�5*� ر��ב���iH�Cz&�6H�����[[�(ԫ3U�,�����,jh��F�6Ҕ�հ�M[�b�u���F}x�b4��a���
a�Q㫔��Ɔ��F�n���J��o0��e���h
�i�5KL���:ɨ"j����Mɒ򡛹���A�q�h,S^�D4��R�CH<�v�f`e�GFP��r:���)e^�p�!��X�rM���ײ:.�8��ك0���c�E�ym���Eֻt]�����M��ydђX�61����F��F�1%�����-rD�U�/$�9�`߷lǂ�nRӹ࠙x�MҼy%!1�ff�@̊�N�u��BͻLj�|���Bj���i�H:���F�fM(��k��M�)r,���8��&$i8n�#C���*�+-cn�w$�-P!�WN�虥"XVs)F�Ye����j��2P�R��a�5=�d��Y��f�`��1�()i���iCU�t�.���~aEB�wv��@ӓm�%��c���.Z�ʦݜY2n[�ܻ 쎴Zy@��S	��̍*�����������7[�F���E,�ij�c�����ZZ�v�n�s6��j��Nd�i[ȡLj֩��kC��.!�B\#�N<^燯�a�v�����N[�/�R+������^�A�;qi�u��A[$*�0[� ��km'�7���j�G���S)!�m�XM�K�qq�eChfG1��u�'�R�с��n�sI�:i�Bei������ċ4�ȵR�i`�>�V�r�5gF�
��*	����1��yvX7Yd�ɕ���߅��M)�|f^V�ܫJ�̧H�Sne�2R�븡��M&����C�lLJ��j<fї�m����&�=�� �1<����D���)V��ҳr���Y���x���8C�>{f�,Vh6����gU5yDf�v�n�;kn�N��we�+Kr=EX7y�������q}�۱���gh<
y��a+.�1B��0�Q�"	�E*̡E_٨��È��v���+QQ)�WH̤Tq�e�����[l�v�[��f�YFf�)P�F��T�Q�x�����Pej�����y2��Sm<�N�[Xw5<�6���hj���Ǘl�V�:S5(��)��n)������ŦU������
�,R��4n5@3{r�8N7K y��)
�X2�@^G>[��f�c��@�Ҵ	�'[���5n�l[�϶�����FƪkV3���(V�jֈ��u�,��b�2Sr��Hi�4ZQ��bwX�wK%���>ҰtKp��N27�y�����nT���8e�{�2��)d[X�;yVT�]Bm�v�۬U�2��0�ݥ�z����4�'��ڽB������;��F��w ѧf����{WB"C�v�wݣ�k9��Ń�Ck>l�����\2�ܵyV�p�x�4�\�*�ܝϨ�[�k ��$WB�@qҨ�0KX���3Tc6�"� dڸM0^l�s]^-i�E[���SƁ�͂����P�Z�=�[��)�;�h{�h��p�p��ztʔ*]��*�S�4�y�]��e`�� ��D�Ȭ�V���j0��V͆��AQZ�4M/r�CXݪ��i���Qł��-;6rH�(�Á+��t5j�)���őt\IE�ň-�Z���Ö4�t����ie� -|䊹4�5b��30e�M(�.Ïzö.͉��q*�J��h������M�y��#�6#$\(�#[AA6�T! ���5�U�Mm�Tu�V�C���U�	�E~H�,>�,z��څLsS�w�B�PnM�ӱ�K��Pj΁S&��NYz\��#���6@�+6[��.$F����ۉ����{�Q��i�!�m|-9�d|S�4�ԅ��ʴ���pX��VЄh��W�ʷb�H��B	�kT�{��O�q�V�ә�J���È����
� �����^�5!�^Q�.���j:Vh�Zz��2�J�M�(��$, Em���ٶA0Îa�o辔���ݕ�*%5���m�.d��X.��NJ0���2�J��z!����C������m'��m6mˊ��dn�cU���.Y�s,<;��^�x�*yA�4�A�@�8�gwN���+C��v
rm��NM�8�42l�`Y�4�N#!|a<��h5aLg4��d�K�-e1��D��"Mk#�&@#�ؘ,�6�x`oL�9{����mXtΐ�RBq@�fᥗN������3j��.S�����8���9A���ڄJ��=r[Փ!�`L��i-f3���I�a�yZn��nlg)@q2&���vw��$�vج��Xn�����Mi�h����b�ܠ�%o-�2/(�M�v%f�4
T��T�1k�p%3]!Mm�4)��)�9󧺨I����+�.O���J�U���+%݅,�tYh���lv�t�*�=˪N��,�ݤ-)���~Pނ��j޹DI�]�ek�M6�k��t��[R��fLGH҂��A�#u�B���]�s`�.9z2�����y��̫b�-��(&���1[Ogs]j�!�Rзe��8�m>������(� �<&�J�;�3n6��]�zK��@0+q��,ee�S�f�!�t����"X�Z�׵/`��J�f'vA2�֓Nf�fkה]�O害2濄��/i}�O-+F�7J�r�J��SȜ��x ���3u�x����b��ě���IZ�I���+2�;B�ON��6ڹsr�BT̸Iz�&l����Yc1�4d��H�=��Sjm��k3JYX���n�k
�T���-V�Q��C��O��)sa�^�7�kp�;�����c"؍J��'jX��$Ƴ
���:x)6�7v�'�V'��7r��V�v1��.�L9�Q�<��Aʘ�nӺy�Ʒ���^�@d�����L1M��@Vh���0�T���V���xA�7lSS+g�j#��d���.Q�*�@_bT�b$d���Z�N��n�:̼X�9�G�����R��tm���0pO���v��N���h��5�Nm�ݚ8�}�E�oӽ\ |m��Ƕkx�}�:��]*M����[Y�Z�V���3��`K�8Nc�Jm(.&Ǽ���U�𣛋y�WW���'9��ܬ����$�DB㨗F�Χ��ni]M��.���v�@1�:|w�5�u�{�1x�-޸�u+�Jɯ���� �?.���tx1��JP4���9}��85'�R���ڔ�3p�s�&�;�
��%L�AJ��m�	�Ϋ9���#ܵ�0�����*p��J�9#0��e���ޞ �ܱz�e�U��W�.��܃Y;��hI�=F ��}��rTb�[�)B3������-Zhpڊ��ر�>+��6��{%�f�|��g�T>�׃������/&��F���F���,�$�y+�π�Fq�d��\;x���l����1�5����`�������Q�{���!R6� �=��i���JBʧ3�8m��Н�U�=��孃���7�I������d+�ya��Z�3�ߤ�j$�wC=��GU��6w7�#v+�y�!c�a�H��{B�_pO-Ԏ(AKE��8�΅����9k��μa�M�w�n��_Y��:bf̔��PZqh'���Y�Z�ޒub.�@7�h*�i�L��ޫ���e��R*���W�q]l�J3�`A]*[{�Ł�(�����"`3��c޼���B1����_�}���ۓ֥��n�duX�КL�U�	�tr�rx�t6�eI���Vuf�{��J����v����b��dw��z\��ɱpS���ǝ��&��Y��������ua�(d/�7jf{�ݔ��!���7�c�,�X"��9#Ǆز�'z��NuB�"��ʹ�,��N����l�]��@���y��4��l�DNv�3�z��Ө3�Ƿz��(bk�@V�t/���)���Lu��"��ͤ��8��惙�}��j��遱��!ݘGJcw����X�M�B���Hv5��BX��+]����6�#�=���2'���<���Xޫ'�������W����,l7Є�RWD�ŸӬnez�w���*T�Y�ux3����lv�
�	��V-�Rmf�c��S�*qc��,)�Oes �(�cX{sF�u^P�٭���0�su���?x�ॅ�=�'�Ԗ�i��`��ƝK]��u�X�����;!2+��,�Մv�vf�\[�p��{����j��T)����m^m:b���Rt'wr��{+�!��ݤ�� q1���P�k�n
y4t:{s��h�l�[�O���"�3X��f����f��rȬ�SW
!:J�Y|�>x���K��m���^;�{�����(B5�lJ�&X�GG�u4^Swl��t5�h���ΏM\���Ww����t%='�^#���x+����8wmz{:б{��+{���+_NM����@�.L�oV�f����!�:Rz3�����d��ws-0�6����=7�k����'VGy�"��{��D�2d_uhd�_L�7�����4���k3��T5��٦����ބ�^$.X;����'�E7=�"ąǊ*�ˢ�N��d�gV�hgi�1'4��,�z������y���� �v�i��� ��w;8�ZS��r�������uei�,��7&�f�����K���J�c���5m:�R�|U� 4Zɸ_�ڃo �u��b�l�7{xI���(�W�����A$������Ft��w1��ql����\����_,"\>W��:4.�1�ұM�X�|YV�_��/1�Zbб^k4ؾZ΍�*N��u)'i�s�Iqo(�pYہ]�oN��P:db�ܽc{Z�h�l�����u�v��v��!�Ky����	���r��;읣��2/n�A<s���K~~Ŕ�C�����\L!��]��z��`�2�m��+���K�㹡�%L�dp��n�T��� p�{�¯`��a������(dr��+:]��'��gOt�V�N�ue�{��f��g�
$[�Ov��ܣ1�Sr��\Ct�Gs~n�:R��ގ�A[���q�[9�C]YY��l��``�g�]#:gu�bK����|����E�85��i� 4��ɉ���I�CL�yn鐝���v+tS!x�p����T�Zc����3Y�î��g4��{ʒ�����4/#�R�D wIoZ�0�4݉�,.���w�u^�p,�lL�E��yw�J1�_qr��ʲ�x��c�h�	:d#��</w-B�^&��A	�:�q�S�gHٽ��s����{Dݜ.s:(Z٨��Zx7�i깚�HB �Nr�>ߘ��.��ˤJ�o]���*kgF)X��a�Y��qKl3�e��~��73e�ʼZ�ڽZ�e�sx�]w���/0Lǹ�9�+��������"9�{z]�-.�Eݼ�aU��R%�&�W+�r�9�q;X1k�ܕ�DP�O����/�c| �����R�@�	��z^׻[��,�Qk���}���,b��;{=��{'��9au>�}\\��2}�����Z�ă�w���e��hp�*�f�w�����b͙�0\5&�|7u�/)W>тT��!�E�>��qh�Q���Ϗ����וY�4����ѓ_�8��c��i	�a���Zw:�Q�k�QK��_CQ���uЕ�mdHg�/<�������ت���y_h��֬Ֆ����.�aQE�n�T̮{��5��WM-^cU>}Y�]��'�K[9�!G�jJ�D�N
3׋.���8,�/�Y��ֱב���J���C[��c�$r|{b+�4%V`k���[�����r�8��S�k1�3�l�/yLF�S>,+����vpY�����]��O���ٮj����8ٝ�+�5��ʛe.r�3�ċn��T��]���f���|xD��|�U�>pun��U�k���X�˶��:[�^,8,�3sukiNY���#��m�{Yј�]̉�?1s���*�9�S8�攋���"���Js���w+\���:j��u 㺓���i��D�t�R�0�B�{�R&m��"��q���=����۱�Ua\�;�+aӌBq���ê�`&Z��6Î��
Ʊ��&v�ӵNI��[e��*۷�.}���u��9���T�!��FZ��}�wq�� j�֫31_�(�+z�Ï'g3�v���T��*��Q��k"�{�g�����㊻Wq�ӻQ��W�n�$R��W����w7��3:�,wuX�z���d���JZKE
ӛ_�P�D�۬��1P���i���]��nIὛ�{v���=��C��b�};kpQ���)�[�����\�qle�J�cV�;�]r;g#`DX�����gO�<�s�lr�0�[�gr�[{Ѣ�K�w�c�wK:�,e�w��_2���-��#�>k=���,�����*󲚅��d��9�k�_��=���/�sxq\X�nf�A�H�i�ȹ]�U��	�wt4�F� �N.W��)Vdv�YJWMj���������J7��EJ���]������t
\[x�eUha�re,�+Y_6��h/��q�a�d����*�/:�������86ԭ��&[���\��l��&��wm.��O��l>�En!���Z�9LU�ao�:�U���'G�3�KV�!3t]=�B���Ӂ޺��͡;eh�t�(Z��܈I[E�/y�UEo����/+���X�I�mk9c:� �G*s7ZkE�z�k��*�q�i�{+d�\��� #W��}�2��xn�\�}�%W��� 96��rh�`���`�^n���N��"��-8=x�HNJ���ǖJy�l忭�N��Noue[x��b�m���vq���s;�}h[��D:e�lL�6��]^e�{P�˭���n�<�=��u �[�"J��w(m�٘L�n���F���i��Z����Y�ڽ�8�կ6j�%��o���E�퍖-X��wY��QQ����si�0�`�Y���T�']�.*�gl':�@3k��]�`�:�����J������=���*��gɊ$nJXD���ƶ^��b�u�6���[a/83@v��Ź;�k�K�ZӶ�ʔN��.��1�=�D���3���m��3s(��eɜq6��j��"g1\\]���J�Qs5���n<:w�	��sw�j�r�p��Tm⧦���_m��I�92PW��5���<�پ��N&�]
��d��E��t�U�QD����x�.�6yc�__ӧY^�v#��r*�α����ً�wYxq�i?��;����ѹ�L m���Yh��ݻ5e������Ոc���>�Yᇻk�!�&��MH#,*�e�.ܖ��m<��;�v��+PM,�nL��n���S!{}�jW&�v���]Y�����/��Yv��;pF��T�� � �ݗ�+tGdt"�і���%]�ݛ�FGXv��F+��Eɬ�Nuu�8
��c<gZ�ɚ`k�U�ou6�2jӽ]gMl��G���wao.�(T������݀��>/��s���(�l˺Q�^neS��[�����ʀ���ﱻ8z�CcF��� e�3#[]N�y|������`������qKym��v��AN��2W����������7���i-zv���m�����}�2`��C".V�"�]�=�� םu�ʲ�,��EΧ�uj�M_5AH��}o�
}gh���Ra��ц\�3�ϯ���apںD����;�}ٞb�b:�{��s�pA�p(�K#��Ţ�!V�����8����jR��My�q�H�L��-����1K^Sa$�n�~�K0�9��TV0.��v�9�ƮwNPm�ڞ�G�k�0�uN�`��(�	v�Q�\
�f����{����k���Q?^7��s��/g+
��C���Z�"�kR�g\0>Ә5r���h)���<���ge��'u��\h�:��u�t�y���] h��u��W���h[�ѠR��3b 9EmMgI�/�
G��+�2��@]��?Vw��֍�]�X#���rB�.B����`�,�=�q�����\�������	p��#i����x�z�i^��uL�u?t��}n��X��j�b��"�gn�E���0Z ����D]�Є��ܥ/�M�.Q*R�C*bc�l��W"��������@r�ս�,��D��jo^v�:ݫ������Y흚WŒ�^,�D	@�y��n|{�Hu��3�Cyˈ���5�-�MG�&w�ڜF��,b�
�8����C���Q��mhvZCYY\��}��I�UKV��#�U���ȳ�,U�:��Mv�$�W���eR:�53kf���uZ�r���������\D�.>��L���y(R)�<{�f�ؼ�v�F[�mʽ��${��v
r�|Y�c��ˮۮ�>a����s2.O��!�F����LTgv#;��u�Ÿ��{}+w��j���<�؍ �R���W(�\:U����e�aF�IHP�W�-��/��S^���-Vf������ƻ�|�S3Z'{S���+��Ns�r�����E��gOs�Y�נ�2T���L��6�c[�ꦚ\K�*�e������;����s^�����=�Ah���rU{޶Qz'�n�r���;��+d-�q����d�)i��}�$�M����q��<���+����Ա�ٛ�P��BM�1�Oz떇�eҖ�������P4�v��3����BR<�@��x�J�)7��/$}�KL�$pc��X�G�R����Zр��nJU�tK9x��G,����kƶ�m�A14�Y�S�Ƶ9+�_���hvT�{,�4=�x���z��	��ץ]l�8>�����h�F&,�wJ!0��Php�G�����c��e$��+9�G�)������n�
�+W>aoQ8!�K��Z�ʩ`��T��;�7�\"Lݺu7����1s�U{P��2�*�[/���a�^�B�@NV��"�?����Wh�,��6֢1H+�H4n�i!u�R���Lt���9�;���+�<��_]wO`�IV�Oi��yp�j���l�;�J�IL�Y�vx�ت�e�ϴ.B3J�]���=|u�.]�{�n��v�ɻI}�a��V�F����r�&f��٥��Ez���jo�ahix�{)���>j��P�ZθՔ������F� ��k]z�����K���+�Z�w(!ti�����%�De��E���^iF����]ts.l�=ܩ��ؕ�tv!Q�x;X"�屜�[��]�p�p<��n�ey;�n,����_	;��Қ»�*����|(�ty�öֈ�mp�o#��!��B7.��*We*�������<}��nFrh;����Ҿ�}��p����k�`�QB�8�R�ޥi*v.��SJ*:Y�U7]5>�"�{�-��q>��{`��+j�޷�fke��t�V�^���w�T��Q�~��������!�6����0�E;
M�-an� E�$c<���sLꛗݴ�5���n����j��c)u$j��G��-�?!}]����-l����l���5C�"SE��c*k�;N�#d�N�O����$����{�)=mL��E�d�]7onsS��ր���v�*ju�XOG\ѝ�4&�I �\��� �I�61���HHIOs~8o��w��T���]v��Յᾚ;��js`X��>�{Ͻ��[|m9�i�h�7�OI������d��9uo��M<|�I���\x�l0}��^,j�M�T�*U�Sl�����c�Aaӛ2Z/m󢃇�ʶ�mj{����^.F�����h[=Z�*ə�=2��7�����O��Gr�j+�>'=�;x"Ѭ�j!,���^I��WgTEĲ˼�{���׽�V<!�'�-JJuYZ!���K��>a�
�bj�d
֗��i�Ґ��!k���!y�%n�٣�9�Eo+n��<�F�d���vݎ*N�}7qS�F���c}��a�Mh�R�j���=p:�$��e�8ՠ�[�[�h���_+�@2��{����QD�u����Rֻ�t�ۮ�( `�L=��˦2�8R��"�����	O%�)7����;�Qga|��e��.�+�q���ljs+/�܆���+���ON�Dzk�ګ�ݗ+�X.��h*��li�M��GA�N�APllߙ�k��)�;L�4x�s[�CB�R��;�_b�y���V��p���m��4i�jP7�Q��頠��#����N��ޅn �ŉ-����	��tôܵ��v$��l�;�s�Y�����n^���X��h3����lG�t7�_��ڎ!����n�o6#�+'ktR�˕�k)�#�f�v��$����e�(�R���
��|R���\0�Wo��ۃ�m��u�_2�ŕ�iE(&4��V2� na��L�]�[� �:�}�'0!�v�+a�f���v�;[^ef�u}�4*�L �sfX8�p������ޣ�U�n������h*Tt��q�ܣ��)�A����|g5n��E�حH���q�"ٱ��^�7F�\��P�JJ����i�h�PR帳���.�{K�Zs �ݺ"vn6Y�eXO0`��nքi��zy.ӡ0�v��4�`���f����c
bY�H!j<A�'8�Y u�Y'K�Q�z{���v��)#��m��9ȵ��!����=���Χ�Ba����1����B��
j|��/,����Y��g'k\7��54T�2p,��N�X��P��}'4Μ_>G
'r�^�Q�DGk%p��Iu�}s/�ɭp�2h3S�O;ϻ)��i�܌*{��t.۽�%Wn�E�Z30* H	��������_,�{���9��9���	���-\� �6����Zu;��Mٹ��ܚblE ��"EE��;zgT5-��7V��}Z�b��u�pk��;�NLSޗ� !ά<�v�����=�Y�r���xjJ�V �
9��gh\�t���8��WH�|�����z�a��ޭ�4���z�^�=�����=���p!�-)6r ��\�����ǃ/�_AM�ᗪK���$=3��I�{7M�w�^�b�����n_�5.mq�aU���;1-zn�`L��nw�@	���f���SQs��95�F�`� `�V��w+DC��e<��կ���[Be�� ��۠���+�h���)#���D�F�7�3���}�k��.�3�Iu������ZI���7��ũQ|�:i�7�Z9Lã+%[2H���{sՕnՑ��{���$f�zp���ۙ�|ΞA����V�B<�kG�w5-�:��YV���s7�=l���8r���cC-}�zi�МR���V��],!k6�2p/t�0>�>��1�M�网uv�6UJ��%�v�6f��b{y�<u�זC���aCа�_Z��倶��٦��K��������<��v�Guж+��7���`e�ݺغu�G<���:��p[a���AaYGX�D�SF�3H�ٳ��v)�x�R��Hs+�~ư+H�;}�ʟ=l�>m�ZM�S���t���@
9(�뛀��0�;�6nJz�V��.��$q�6qV�sC�ܾ�c�S�˺У@_Β�J<��K��әZA%W^�,+=��Zw��)�s-�f�]|��9���l�Ը9�-�i�ώNp�gj���)�Pg 9h�2�����8��gG+�
vUN9N�Ϯ�!˒p�H��L�]��a���ʒ�+̪�a��羓�1���xyl`��gK�v��va�C�̢�h�#A�ЩFi3��g2kj�ڮ]rgQ<���y�K�G{y�s�y�M��ܱ�)ָ6�[�.���ή� �2�Ų]v��l�y���L���.|����c�đ \7'6�O1w�[����tt
����% �GmU)�r�\������ZO��c'��$2C��=���g_cu��N�w,�8Gf�4}�wu��λN���F�θ���L)m����c�0��S����1CV1؃��<7)�M0+p��zR���f�S�.�%XKW2WP�wr�&�J䫩��Պ_b�u>�^�Y�5��_4:�,)jaN����4?�w��t��v�D�
;
����D�nn��8ygvy�mZ����+��ަX�lx�`�9���[�{���9�6*�P�z���{�
SW�&B�l뮗��2ضڠ�HD��̵��p�ڟpU=e�0v�^9ۭO}(T��o)r7�wk���2G �N*�b�v?��7Tg	M�eù����=��+V�:�',�5z�R�$���Ƴ�s|`��G��^|�#f���W�[�`�E�+v)}�T�P�;�wRh�����^�{�s��RW�����ꚫ��0d�sH�%�@���{"R�L}�p4z������u����E�ӇG��\P�-U���V�'}�����s����̵ ڷ�P��3#`oMݬ��I=-�Q�I�8ckt���9�\�:�4��툹�ڮɝ���;/[:iX�	u�8 ��Wnuݓ�D��ldb]�T�E����sT^��HP�l��A϶b��;��|zb��F���=v��v�t���q��x89���dڳ��0�O��7�0}�OzSOM�ӝ#�%KT�rW���W��9��*�)� ���\
�XU�"���=6%m��l��#�H�f��*�t�jY��*V+×�fq$_>�z!!+8�GJ�gZ�k�)���=;�3TZ2a�>�GhXr��Qyf����0$w��ˆs�72���V�j�c��ې&��L�v󋮮��^:b�㔬��ʹa!)u��o��g�y�t[�q��/�=aQ�����0���v�Qt;rU� �D�Ww�	2�U�%�S����eügi����ZXJ���*gY��*J�}ڽ�(����ur��gA
�U4b$ݿ�#@��[�����v�+{vY%[�w�9S���6���>�u��Qִܗ��*�6x�v���wn ��ɐ�Ӑ�]�Σ��W��ļ67B��p�c�8B��t�������y�78
���L�"��Zn]��kl�ek��,Y([�62���n���3-�����2�4�B��$�f��b���*ݸv	hڃ�cX�Ew2X�,*�YY�;r���_�{�"�!�� ܋�:���r�wj�[�����y�K���<Hf��r�A ҫ|���
Ƃ��*,t�\1�`�0���f)��l�P�����ھ\�0vմ?f��'�;��!�կWA�Ժ�g�3����g9(��pe(8l힐V�#mhS��B�����kR[v��k��i���D��\Et�4�fI+V�+z��|���oc�)��$��kl=�pDm �;�!�]rb���_*��$ېj��]2Y���oٷ����y����D	Ւ�AX¯�s�.���4J쬏�ڒQq�
���b�M�����o�8���}u��;p��$�򽆮8� c�Qǻz�;̰�cg�sȮ�UӸ�r�J�]��.�i��jd��/#�e^a��Gt4)��x����像g^mgW�o��+wZT*�M�Go�Z�N��������}�.�f��	�Pe�X�m�	�ŋ4�<��&�&l�>�X�J�s`'\X�S�2�U��l8�w�;6��]%���룓��� �>0�����4o��h�\@X�]ɭk����f�ѱ]�Ø�A���1zs1�`#۩Uw:���3�
�NQ�+f5��cz�lt�/s��o�,�ڎ�r9t��+�&۬�p��ֳ�reop��i�l3րx�,�p�D���n9��"�^U߲��w��=�9��.��V���8�r����tT�A�'u�wy�緣w؛����yu��2נ��4���^�$X���\Su9�����4���u�E��K�Sz6�V��H��!V���ە�v~|+^�u�P�o5eбt�t;t>v��.t�Vg,���W�Y ��G�k�Gr�K�f��ڟ!U�6i67&�[%gp�Z��SC,��j�V�v�K`��I��L^����;կovm���7�z�d���9�;�|QA����o�4��W\��L�?Y�9�|�84�ה���*���c�o��U8�Fr�p��C�]W������#��(�0U���o�ai�n���xB��������sj�K�jx�Un�"�h���ɖ7P�0�	���,3�q��e��j�>�2���`('��Ai]n����`wh؛�t����/`��@kў����Z�l1^�]�/���B0��<�Mkt�au$A�MԂ�A���*�lWL����
C9�:��n��뙬L���	�r6�6G��HvB�v"4���,Z�	�.�5-6����{O����9��Y�u1�3Bn��)�a���W(�n�{g�D������l�ǩ ��^�ƨ�"��p�NhW91b�繐L�ۘP:��J�\9��򦆼�D����OS[鞢������Ǐ=%�jͽ<�J�;�bYkSRB��dV�Ս�F^YS���"*sG
��N��\FnGRQ�Fdf�v��JW�z�l��Vq�
����2ɞ#��д7��O�W�)�g ܻ��Y�>���:�U��D�9#H��i�c���|圳�%�a�u I������	�r����Q��o ���2��aΜ���tލ���h�OO�J�ŕiN+{~�z.��Ed�V�X�����:x��;�򣐳��`����dw�Ĉ&֩0tp,��K�(=������u*��"��Hr�|�����@p��ޜq��_e΃�SR�(0��F���	��Nj��S��"�j�knr#!�:ۏ���&�dǍ!�����U�;/����[�톮�s�tjv��q��hp�3�0H7t)R�Y�*��A-� �>�b��:&�kK��-N��� �w����aO}vo��%Fb�%���W!]}��� -%+NY�`���f&0zz���x���2����<�V�0p�t��JqvFt�����|�T�� Ć�A�63V14؛��}���3(��Fݗ�Ҏa�%��:'$g{e�tofG��nV�#7$����YY\�{C�ޠ7�@��s�����l%�����3�����S�bզ�$}k������|���=3;�ڤ%]�4�6�Eڜ�q��#�F��N��;�r���IZ��q�7y��Nk޲��m݊w�Y�}�<�:��Nd��}����z�/���~�v����h�����x�d������ݐ����*�dJ��H7�o`i��\̤J��aKɪ��M=z/+����+��d���A�X��lW�m	�q޶-���v���W��nK)6��զ�ͳ�{�Z��&9d��ٹKG=V�e�Þ�դw`ɯP�n��i@A�b�R�43Qx��J�䥑��RTq�[����hѝ�:����J��Cպ�#Ӱ�[\_U�C���Zh�@u=�{���%�<�2�g%p��cY�t!m�$(V�={03��=G*��C���M��N��v��`*�Jr���t�BJ4n
�Y�.٢r������q�;�R���v����D�ۺң�S9vp�(k��V�\Ua�H;�X��j[� �����4���κA-���u�<����Ά-#MfL�P����0N�h��J�, �v��>|5�;��"��'Y�P�{h�2�t�ڒ�I�,��yxF>b�LB�8ԧ���&� '��M��m��R���ǑO��(ޛ�شa��������4�g���o�D�'l�z�E5-���rh*�Rn	q)K7x5�Mo_P`�aci��1��#��uoC�{��V9��/nW�8�I�~j���|b
VM�ES��rf&��s�_M�i�m�He�S��5tj����yB*zA� Y%;|�`06�P�Jx0e��/�Q��vɜ۞ML^M��ׇ�4��nNt�J�MY;y�30E�m�`G͔mw �5ݯ�ϥ����kkWo	l��o�Yp���$*��7��f�V��
�0�tfpa�R����Q����a�s��ھ�MI�+K9���6x��|:�%����)�n�zn�뾍YZ�}ם�^<�NM*`����oz�����u���`O��l��n�y��l3%p�喢tb����Ve�
���U�S�"5�LI>�ʏ]:�����^e��b�)nvb�J�S��[vu鹸Ci����P�SD̚����3Ԏ�uh�j�E�� ��T�+Sl�.N�vJֹ�b�ͧ�44-���Gb6=�ԝp0��:�v�XW&]����o�.�Xᙼ��iS!<�!�9�Ou�����	!I�5�}��揻-5�py�t��`�>���;u/5GQsù�gxoF�۔y;�к����o��pձ�<v��o�9��N�uUu�����s�v��h�f�c���wL0��v�F��;�)3�]Tه�n���n��<�c\͘)�/ёE�jl�ʟb��z�$�D�fXD����s�<��R��-$�������O|+���ڮ�����"Hsu^�Vʁ��*_59�Ew:��1-rg82:��h ��K�ڒ�vk�M��<:�.�띀�7��)T6yz��<�,3XV(|����[�#����|�2�5���qu+�ޭ���r��;��1yم �9nm�睮���a:������#�9��݁��LawI4�1~,�	�^Io�f�؞5{��}�N��8���l+��&7�n��:�m�7C, 
��4];�w"��C�R��)���-�l���шl��	��`�\4�Ō��@���}q��S+#�i�290k�c(#;o`��Rk̾:$��T�6��XKӑ�K�&�M��OZ{F:�;����艇�!�s{�i�1���'�%�n;=��(�=�gR��{�nK�S�ٮ��g�nu2�J}��:0P|��țE�)s��w5��_�&�ՏA��>�4�_=*�;�OC-��L�m�N�3.�04�������x�ܒ����W��p��� � E�����#m"�m���X�#Z�2��R�L�J1\��1QA`�����T+"���X�����P�3

J�Ɣ�,(��*Im�*2��P�A`Tq&"Ȍ�����X���������0PRT�@FA�U���+b�*�X���l* �,�eBbJ���bB,�%H�k@��h��h
���m+�`
�Ņ`��%DaPR�2W1�B�P+,*&5 �s!*V!1�%U�L`b�,"��B�Rl��IZ���X�J��c�Y"�B���Y
�(�W-��dX�)1jf,��bc
������Q@F � ����~~���U�����<V�xh����덁]v�8q�)���k��x�pW��h��"�p�L4j��3�.��cX�Yu 9�����q����^R�>e�s�*�n�B��Bf� UZxk�K��5t���ۗ��޺�Q/jϹ3���yp�.��(e���o��	a夅k5�W�{�1S��mF�3ٹ� ��ލU���v��]������T�:২�!�ʢ!ݫ5�k���������5a:.}��&�N,K�X�k����f�+��(�I��8)�K½��U"h�N�q�,!��f�صx��y?�[Ϸ��I�+�dO�[�=�?T��+A��x���#�oj�#��qz`
�/��&7�멏!���凂��h�춪��X}���K���v���3��2F�|�[K��O�>
�s�բ��М��L��YL�Gn���#s�C�K�N-�W��Ԯ,��Xb��0��5�Ԗ>�Xح>n쿦�c�J�"Y�l�w3����g�e�긡ݬ����r���zw���ah��#���)h_���g´K����N��.%�z��^�a�������絚��4j�����hw��k�����/^}w������,��S�u,[��$ ����xl�;5hLׇ�ݫ}P�l�:EV�v��ܓm�m�7�@؋�o[�v����1�=$P��5Ҧݜ.�����2���Y�֘�7�N�%�)K��]��F���Z:|�3�H��/�LP�\�J�iEza0��NPضs���G�[�o2p�WK�L�+��Յ��u"��x�$�z4�k�o��FE<�.��Z���9�������3�>�I�D;�ߍ!�جv;���t��Gx�G����5��
��=p]�w|��M�g`�B	^�{ZC���<o�K�j�t�DK�h--�u2�,B�� @��9��ی�V}G~�t������9|X3�a����=�Kx����(D#�g���^��<W����e
g�*%��>�=�]����i�Cz�����}b���繩��D� k5��u�]�*�.���&�J4����Ji���$��9�.��}.�3�:��2��|Y�v]Qgr�x[�b�ޘ)%�'��"J�������"���DZ�tؙwıL�Pp�n���:�����5y6�>�n���	�g�x�ꤞ�B���w��d��r:]do�WZ6}5xi�yTA���3�ȁ*�Ҳ�(o�V�E��0�K�l8��;J��e�ꩭ�FFS��곚{�ݣQ�__mp�Z]{*�[��dĲ���f�X׎y��YLi��gT�@��d��{��b�93�Ϗ�u�$��r�����6l��o�89�(Ż��R�吻:�7g'z�/C���i�c�|�X&.����Q}/4����g��>h�Ӹ��;��Q��.��Ɯ5�<vӋ�f�����fP��Ǳ�9�7W���j�"�u��4��<z)��z�������Rƫ�,2(_��A^�2S��־���%�K��;yy.���x-K.w�m��s3�GN۫��w��V��z�u ��n*�������)�T�`I��7Ý�?�v�˦hp�Oo�uL�M=Ԝ�r����0��z�cx�� t밺�����jr��N��w��eL��k�֧a_G9�q��6a�xw�c��q��&)�]�=��ɵ3���W��7�J�s{+��	عU4��nY�w��ޝX�p̭]��޿��_m�?\z��Xs�˒eQ����]���lg��]<�X�_t:k�ϯ������ۦ0��N�f|������k3 �M#}�;]��Tт�FI�͛�;���6�V#�8��8k��:M
�6���#]A$�j\m[-��W�6�X�=��,��f�l���\�yO�m�b�͹��S��w��g�o�n��:L��`�Pm�������v����n��˒�ݓ�Κ]:���B�nKf\bz��R�;��<��}ٮ�Ǹ$5�nM�0JvJY��U�}�ʫ����m�M�\�ܛ]=^u�n��L[��[�Γ��]zz��m�WO#�К8��}��}����U3���'ӄt�Jv"�)?e�{ϕtxn���ɭ�Tv��	�_�r�)����;����
�~������:UP���0��>���ꬂsږǟ�9i�O|�(=��l��;{U�¶�SqZ~�/e_�Q�^��(?V�W�_m���L�g�S�����x+;:�|����%O��f?���};n�"� c��AΟR����W��a��}�Y�庖��g�I��rz�Vot�qG�zk�(�T�cn+���W����Y)�-�npu:g�G�O{p9����ࢍ��
�~nHf��^V���"�2��+�	��<�C�j_N������Xr�1�����]ڰ������-�2�La.�:��9B��l�C5Z|�_��o��1Gzkد���*tw1���7(�(r��QnLo�s����j�EՖ���X�:���L�Ͻ��ɰ9�_�q�{��z�u����:W����՟f��_��6���;ï�ٽu��sv�$8X[�|���}�S^�"oeНlX���,��G�\�g���&�w�K��Z����#�υ����R��BΚ����� Z�%1�t��O��;�l��@�o>��%��%ܫ�xh>�x'�+�˗Y���Vzt����̗�/O����:���{��z0T�K�:�t|��ͣJ�d��1En�T�/��h뱺̰$���a��I=�����VT��0��8�g�w2�q��C����0o4^�Z�����p��j�U�sq톸A�9�a��Զvw���뻤�7����~�������j�rގr&��L���$�㱝�����>	��C�Zw�ꩂ2�W��L,Q�?gxQ֌0�ſPS{^�p�Ե�J������H�"{t�I�p�w���:7[��n9���8��Al�QhF��x��`��v<���gZ���h��[㌷��VQy��|,�6��xa�u����C�j �6� �=(7 �
�c��]�2gJ�sܯw<_b�i������	��v��}��qΟ�-��\�ѕퟆm�������3c$�����Ʒ�8�3�!�H
�u�~>N�e�p^���S�p��-Լ��=�&���rn����S8��:���q�����1�{�\�S���W׺�V��6}�#�~��cy�A}�qa�N�^�N�}Lu�^���r�ru���k9U��-po=�� ����}�;6{�N�;���J�M�vb�%�v;���o��`t.v��f����]:=@��k�s�`��ul�G6�#����O���Η����쬑��Se��
����Yˮ�[ۼj=�C�+��Κ�<�	ο���&K�˝v���z�g
�;Gi7]�rA��Je�
wZk�p��v`nk�W����9/Dm�]�
T�p�y�b��7x����[��_u��z��6OT2Ln�#��e^���u6����V�hi9���h�˃�=��C���1��6�#/��Xx����c*�%��*��-�g�a^	M;:Ĳꥼ'�ˀ�7Rd��PP�].	V��G�q�q;��B	є|;	_o4��{Y������nd|r�V���v]�yW3dǏ�ʶ��^�����{<�kQ�}�^j���2co�\^�����}�V��p�tv;;�2�}�R}�r���I';X߻w��������5�=8#������*_��wEJ��r皋�:ky�P�>��=�mA��o���ގ��Ŝ�.[�o�'�����*EF���jFf��N����3g'�t�w�~��9��T�h����F��S��#Z�kE���p9:�Z^�Y����>��M�}K�Ѫ�6ϕ�n� ]�1�����S�7���ѷ���~�kry�M^��k��}�I��4ټ����d����ّ����ea����C�6Ǚ�x�l�t�;���z�sŇ�:�.�F!��NI���){u�*SY�ݙ2, ��v��N�{`��h訕j	\n��@؍9�!�B��J�?(N�[�����ɼ���=�0�&���E�����6{��
�(��'�(����{��K�s1��Sw��G6��-�_�E��q�m�g����߹߼���<�=�q�^�<��������S�&���N��u���T~gΜe��R��nGg/3�^u1�����qv�Qy�p�~��}]<�<�����v�Z�����{�;�Fn&�{<����ɂ\�3��� �|/���;w9<�]��)w\�;%7/'�ى_��O����J�V�%gMӪ�=���ۆ��/v�]z_l��|w {\U|e=Ϥ5�aɷ0J��z�'�������^{�����+�ڗsݟ=v7Y4���S�D��ӿ�a/#��i��{�Ղ������ۋ9To����U�1`8�g7-]�ы��'*�鞹�=���K�>R߯�w����~��x[c"��c�n`N���/y����?��膏4��!�=1<P{��vxy��c�k��z�_hy}�WVƩ䏖�iz��K�j9s�I��A����uF�b����2mJ�,p1��æ;��o8f���M�ȸ���Z/R�BU�n��6~'h�qu�c�2�LwqW��rУXgV-[��%F!&���h��V����v�3��=�s;�n���~g;����7��أ|��p�Ru3ю�=}Q\~�D:�{�l�Hs��`)�����z���=b������1��y�瞤 �'���l��n5)��Arxѫ���'љ�݂d��Z$c3�/CB�-�����ƧNG�O{\��wI�Q<
��;c��Ơ��R��Kb��|ٰ�����J&�.s�y�ni��3͏s��-��z��u�K�Ԯ��ͽ��d�Ivm��	ޗ�9��������ֻC��Y�N���ɷѽM�+�7���+d�k=oe;n�s���t�}�:/s���qju۷s6G����z�G=�Cf������w%ք��Ju&M�UQ֥$�^�%�T�4�㏇t�ϝ\xe=rW���K߸^NG	�,)���J�?��q��Uu=}�L}9v���s���]'���{�)�
������\�dӋ��n��#�]�y��̱��0�m�vm�7Gq'�tX]�b���/�8�����(	�o�Dۘe�S���:}���T�+p���5���՗`z��G~��:�Y�&F"c~p?�{�*�Z/t�@�Qܛ��P���`���;
��5��{%c�*����~D��-���f�X�K�;\�J`�����ir���ʛ�)���)�{��m��o�y����޿K���K�L�SÑ�hk�ٯ~Ү�FH�r��թoS��xb:R��+��س�~g'��^_m	e������]T�}�귷
��6�h�/s籜�{�-�l<�fUk��vE�|*��Ǉzx�+�D���ܴ��C�����k�rl���=�ۛ�ĕi6�=�Q=�~�^��E�_�j/pC�[6�`:���bǌ �:>y~»�Mo{�6n���Y�~-�Lu}|���s���^���qzy�wL��=C �̊s�N>۝����t�v;-{Y잯��R�;.D|�h�#"�m�ݝ����cr��>��+K�d�q��(=��y���춫9�'-۫�9R�̽�n�vXYVwɵ`ûRƼ�X��K�W3�r�d� ���2�[�x��ӷ2s&nPJ|'�w��˂N�3q��p��k�����D�SVSp�5��u�݋|*�<dTQʃ����ȝ��VPu�VX�K��/7!��`�1�O�C{|�b�ӂ�/.��l��
��=r=̚�rM�D��X2�OT3�.l��/s4!O\v`����aW�b]᜻i{r�s"�흽�S�>�l��m��H����\���4���B���R|BsLu=�����,2�tO]����D�Y�l�&��x��ʑl�:�9� �6����W^�c�G͚�Ô������L`�I��0�jC���\v�ӕ����$3F�~��)��G�Rx�Q�`�F��'��[����v�)v ��ƻ�d�,�����5R��p�cv�b�䐡����eA���6���u �+�Gi�Ή�E�Bi�z�C�f_e� ��S,�QuT���O�}��f�}Xl⌜̼wV)�k3��T�cGN�)���P�R<�ǯ2��.fMN�]�ڂ�W�קǶ����5|u��e���X�V�|i$�:���,p��(�x(.�C�t�@���$�ͼ[D�,3G�ީ�MW�㔸��uNד�jǕ��b��/kN�GG5
t4��/�5��k-4w;~Y��;�������F��2�}pr�E�^��р�G�f�u�Y��2�aK�p���Yi.e���z����}F�坲:���0���ʊ��A�$�U�o5̴����^G�ű��]�	�VP������fd�e��yz��(KT�l�)��ȭ^��.��W�b}F:��	Kb����p i�_f��m��Yq�Eo\f��YUOCBOwD��oi�{"|MW��ڹ8Aܫ�( �p��Nۄ�}���<�R��sr�v(t���@��J�E�Δ���Aq"�u�λ���ي�6E�.�8jUJݻy��ʒ�7�|���;|4���96�A%���Y�k
Be���R��#�m�O<�#MK9wP'+P��6Ŕ�����&�
��d��C���e���di���S����)�޳,=�]��(�@�9;�n��O�}FS;
�wۘ�gd�}�d��躣ZԞ:�s U��wc��]n��8f��G���=�2+�L�����#9�j�O���;fN!�b�ϼh����l�7j1��c9���-`i�2xf��iw��㋵�j��v���ɗ��DY̘5@[���]y��5��<=5��59�:�R�����!��a7"Y-��ke(�[07��G���;m�1�vUj�w.{��{W���AU2��6k�R���Y��_@Ĩ��Y
�ĩ$R( �G2����)*�E�"�aU*
�J����m�������RTYKam%ADk-��m"�mAed�,mH����µP�e�

����"�eH�Xe�c+����
����Vc �)PX�U
Ȳ�L��RJŃi-��L`bLHc0B
9ed���$s
$�ԕ����a�5�����Ơ��E$��h��
��I�*"�)YR
�U�F
�Q���Z�m����"�iQ@̢��$�Z �KH)**2��KB�bE\b�@R5�A�*�4h
�<^
������<,,[,7j��o������rQ���J\�KO�F�f��׹���㧅�S��}-R�[�%7��Z��%9���P�ڛ޾z{��غ��:(ro�Oms���ۻ=y���'|���~��y6\�ʟ\�ʑ�N�"#�uz����������K_(�)�}��!�}g���7�8�^>׹镚kU��$���e?!o5���볎��y*��\�*�3m�S�8�F^�Y��b�ݺ}n�zf�s*���[�ܾ#)�{�P����bО��}���xXrm���8lg�ɮ��w8�7�����{]���`܃'#RH��b�p?�}V��l�W��v��Z�7���f�۳��T���}O��F���s�9��c;�S;=��5��>N�N��'�9��ؼ��qu�\���7���T�GQ�%�27
~�fUl�Wf����fb�4������yph������gJ��Z ��j�Ҿ<2�`����jݦf	��i���fvxF3����p�{�;�V�
N�.a�@9_����_$�i��1�{F��ie+��ɺϯ�;E�q	�&�W��ۡ�(���f�-�UG�z^
_>�0��N�dӛ��+�{��ƾ7'����G��ʞ���1ծ�A�������}��b�u�:�{<��K����=��H��f�&����^}��:��`kW���0-W���N�Q�0zGbT���{�{�6n,9@v�v��[1`qf��o�o�)���y�ġ�t<�A�a�o��N�����iu����͌�̀%1^^��W��?8%��WN��ݴ�gz�i��{��\�3+�^����ˎo�N�����^s��q���Y���:��3^c:u�M�}��7_Έ]��u�m�6���.=b_h�zw�-y�ծO�tŚK�~����Jw�.���y��_��۠��)�U�sf�[gM=5vdR��u�J��u%Xn��N��m�s)c4��>�j�K���>�U�����*}��$5�`96X��߷�0;�:#|=S�_Lk�ʰ1�Dч��e�Z5�s�sb>��d�2WvZg6�ޞ92<X�����(i�k\y��,;)����c!b:�j��7:���l�e1U�\��'�y?'���	%�Fju��i�E�;"�ҭ��/7pژ��3���Q�$���C/Ӱv��݄���L[��XC����4�ޮ�?os��ޓ���綑��G;ٺ��oĹ�|�B9���~&����a�7�I��=��#i�cʸ�8���ߟGv�7}���{&�5Ht�����sH��J;=�y�O��W�<�{���w��\��h�y����I��l����Nd��繋�s~�����z�|9^}[�+#�tǏL���oܟh���-s�K����޸ۑӰ�\E��]��9웗�n߻���g��+�����sm�Է�v8����F�:~�u�=�����E�.Lb��N��q�-��\=��ﱹn�L����O{|*ZWS�?Y�lJ���S�q��üyO%���:��f�zd�A+�f�Q[Rr����>���k�k'�����"oΏQӢ�;<�J�M�{�7}�/�~����>�8e�pq�J�er����a-f���g�/3�/y\��ءFQN�ݒ�N�:�-�����ϐGQ�)�kiļ�l&��n噚Zn��� k����J͘Ө�":�_m:���A�X1��SO�ᘋi��E˹6��Q�"�a��׽\�N����tP\��:����ff���S%j><���W�|��p᧍�徻s�(�gI�����5U?]z�D)g��H�peK������jO?)�|�f�L��RV�V�����V�^m��A�s�xٟ�Ԟ�d2���>nk�W���>@�s�'SL� �����C䚲'�`��U~�f�JyK��>�>�_}R��<���6���):��'�0�@�=<�O��d�7�]�i���%N�����N��|���'�?y�o��[�1����ú�yv
d�;�0'P��Gu��I��%J�u�"ɽX'>d���?P�d2j��Ěd�=��:��}��$Ĭ?d޹���O߿{Awӫ�����4���}d~����A��8��V�)=d��c$�7�I_'5�H�w��P�i<}O'�2q�����4��7�<�$��~
������e_�d3��@�L�z¡ӻè,��=ì�A`js���O�P��0�I�'��{�I�MM��W�I�M�OY:�2é'��L���U�wP������_�������A����$���~d���xI�CS�è,'�s�u��P��=I��2����Y>d���䓨=�!댟2q��<%K~���U��t�i��̏�R��'��5<���B~5�>f�8����'�u��/�k	<C�jo�:�d�3�}�Y8�	�;�@�'�Rzk��O��gu묊U�x	�\*�P.چ͆�V�C*(8m,�{?b�b+��{�L��1T�uhF_>2��^x��͞6�ι�I����1�7�Æ�ɂ�X�Z��v*��$l@���fl�͉�-�"�<���_N���Û�r4F/!,��ng������wl'�$�Rc'��,���&�FY�I�V~���[���OM��|�:���'uN~���'����������N�~�������~�=����9�t�'5�'f��q��O��d����OZ��N�YBz��:��8�m�Oƨq�g��u�[�	Rq'S\�q'Xp��<��盼u}��_�{d�a��d��	�߰�'|��w��u$���2J�l��C�VO�qe��?2q5��I�MO�8��m?kxd�V֧��q>�|�w�^���&�S�����?Nw�I:�Ù��6�l��nI=~d����'N'�y�T�H~��̬�1H�>C��OfS'�q>�o���k��^y�|��r��r��>{��d�+�P�������H,�a��o�&$�,_�i��>rl�&�7��c$�h�쒤�|,��~���6��]L;�0~���>m{�=d�vY'�>OƬ>O̓n����}d<��Y8��h{>�@��4y���OY?2y��;I�Oχ{��M2wz�c	��ַ���=�ϳ����t�	߬�
ɴ��6�l�I��O�7l���T>d��!�C�M���s'Y6�js����0���|����>�G����VO�ՁW�ە;=��I8�2v}��Y'�k�a*
7x��|�����M�XXN2|�a֤�f�a����8s�u�|�'d7������?s��d��9����K��u�@��N3�'�Y����|ɮ���Y'�<�*V��
��VJ��d��o���'��<���&��}�H/�4�<�F�c�߻}r����ɹ_�?���;9�0��o���8���¡�� ���rC�|��S'R{�2J�$��
ɷHe���2w�4��~]̉��#��P Ɗx�q�������Ot�$����=�<x��#0���M;T>5�f���辣�5�&_�V+��^[�oð���!�<(1/&��Ɣ�j��ޗs�va���zn��Aה�h����k�-^��7�/F�1��ol�/�~_ee}�����d��&�h���$Ĭ?Ns��	��w&�q!��(q��}��'�?�O�'oVK�$��ԋ'_-9�{��g;�7�=�{��VLI��c8�wVi��L8��d��N!��βLJ��>è,�����8���;�Ԝd�+;�!R|���~a:ɿ���o17�w�g����~�ys�W�O|�,<v��je�'����2u��j��Y4��<5�@��d�ɽ�'�u�7N��LNyN�m+!���zÌ�%a���J��yB�~���o� @~����}>d׾d���h݄��&���:�|Φ���0�OS:��>׹'�i��>~��'�q��N��I���ν��w_�����g?k�?k���Ԭ�w��6���Nv����M�ϿBz�׾a=q�L�J�i�O��,�$�*~ՇXq���I��d��u���t����s�}����=�&�i�m��M!�)�M�a:w�8��M�$�]�2|�����VOP?{I�Y?0��!�?2u5�q��!x��H������e�u�FFw׽�k����ꇩ6������8�Ĭ��p'u?a�i���u�o�&�;�@���{���N�O�<�+'���%d�������N&���履�����������s���k$�3�$���̜J�ѿp��8���A@��ݒu����q���ޙ$��&�;��8�q�y�Vd?wm�ϻ��8>�}�ow��:��~I�*C�c'�ܦ$�!�j~����6��d�V>��:���6{ܐY:��\�߬&2w��M�d�v��i;�<�3�����}��q����O���IY'����%a�!��l*O�X)��'ٔ�i8��Cl��mѿ��s�!�9��q���{;����a��s�l�d��y������ȳ��gfJ��¬`m��I�x����G6�Ϸ�j�����P+�>��FV�)��7�~}�5���u.c�s~��3��|:HX��kG�J[�*�E�,�����QDYF宻D�ÂWN\�����k�}�OT�yw�z����J��|>�O1gF_{�� ��&�i?��Bm�d�w��c$�h�쒠�07g�>AI��6���ML,�i8���m��N3[���N��<�@i C���¡/f���N��^w\��w=�O�'O}ͼd��Ow$�u�ğ�&���f�59�?E�uw̒��3vq
��VO�@�2m4aa8��a�4���~��i���/�7d'��w���>k���t��s&�'��gp�'�'˺q��>9ܓ��O�i�k��i���I8���$�RL>�IY>J�P6ì�?w�o��>��;s�|�w����M�~N�Ö�m��`m%~d�7��d�=C���I:�8v����;��$��9�	�>d��	ԟ��%ea<�=���~�/��s��{���IY3VL��'8�M~��d�x���N�u���l�a���%eC�s'Xu�sǸ~d�
CG;�P�OPY��p�G�~�;������5�b����<��8���$�a++	��N:@�):��Y�~��N2�CO��d�M��>N�x�Ϸ�I1�}gX�LOw�:��_W��촗~��Xn�7|_��*�>���o$�s�1���d��N�>�O_?e��&�Ghi�����u��$�׹��'Xy��XO��a�Y�?>�=G��V��s�3� >�����Y>J��l�'=J���V2~�Y�$�&���_,'�t�OY4�2Ì�ǩ��$�	�T�?2u�~��>*"��"���=W*�}�?#� ^�M!��Aa<f���6��t�=I�O��zw�̛dѽg̓����'�2|������M&�����T�<�u�^%{F�/��{2�|(�!�}�?Pda��O��!ԜA|����I���:�d�3�o�:������d�'��=5���|��%d���'�d�ϡ��H������
�VPO������m���&ֽ�2��f��ڥrbw`�[��?1��f�L��ø����5\}���wЬ��р`u����y:R^�+��rdI6f�=GI��0�e�<{�=��=m�J���'܏dEo������l&`��W��]xɴ�eROYS���L���N �k~�!�N�O>�Bq�Xh��:�a8���N�o�	�9�:��M�$�]�:�=|���o��{��9�����%d���ed��hk,�����k,�	�*~ՇRO���'R�=߹
���J��	�a�~î�'Xxs0�'=�����T�V��\����ճ��w����_�'����q�|�g�J�iŰ�+'�?�5��~I�hˌ��:�è,&�f���N2�9��I�N�Cs��?}����^uّ$�^�ͭ?����a��aԜxɴ��yRO_�;�d1�m��%a�Cv�䬟 ������5�M��k��S�$۬�C�8�~7�`��겧�,�UwU�bRb�2xɧ�w�䂁�?k��N�~d�k���<I�Մ�z�ߵ�ē�rs�IX���q
��!�d�Q�p��>����\�i5���]��LRW�}���C��{d<7��u�o�{������>v��O̜�'�M0�o\�M��4s�~&0�CGd�	�t��䬛3�w�5�/�w���ܯ@�OY6���=a�i��:�Ն�;��3�:�׌=���'�&�M�I���o�d�M2|�I滒a����$�|��J������	������9�z�}𺫺��~�IRm�'�(I�M������3����q?}�Ci+�'P��ԓ�<��4ì��G�?2q��s�'SL�	�|f^�M�ȸ�u���~�P�@�'|��q'�d�*I��ĕ&�Y?e'Y>d����a8��x�Ϭ�d���]�iO����Xh�p�'S�l{��o���x��z=���R���Hv}�AC�OPY��u�5�a��u���IR��nȲo��d����M����&�6���=gY ��=���G2��B��]��=�*���sf�����*��N>[K�@��!�׹	'FX�C�y��v��t6��Ӑ��PЗ�e��;G��Ӡf�vmM�ԉ\㇤O*�9`�}����G;vd��]WX���w���?C��1�@$�}�^ly�=��֙&%a��������0�'Xw ��OR������~9�?2N0�ߙ%|d���"��,�C����<�a�N2���sǔG���?wf\{߀��|���������:}��	�
�7N��LO����M��5��z��>eC��*OY<��I:ɸo̒�2NnȤ��'S3�|���o~s�������vyCL=a4��8É?y`x��8��}�$����è,'�k�a�N%Bh�=I��2��{�=d��_k>I:���x���k\fz?��w{���8�'�O�a<vɤ��0��٩�$����4��(��>C��A|�XI�CS}���$����q*A�s�d��K��.��ڄ���޵߫�{��J����:�����zԟ�8����d���d��f��N!=��C�'Y4�$�2u+<����I�59�'SL��r��|���:������w�i��'ό'}�d�&���]�:��'ϟ��+'�ۤ��?$�*��N�gM��� �N~���'PY4o�%IĜeN�y���e�ذ~O�L�A*z��u��-����}��m:���}�2q'��=5߿Iԓ���$�6�(|���!�C�����S'�u4~��i��3o�������|o����t=d�V<��6�l���������]��a�gXm�'̜�ܒz�ɩ���N0�O�$�6��Z2�|�'�l��'��y������7�>�Ϸ�g��Y'�i;�����:�s��:���}��Y;��dN���|��bM����&�;Ϝ��6ɠG��Q������G̏�϶{��v�����w�}�͡Y4�ö��d�jad�$�i��&���q����������ݰ>`u�'�ͼd���'�]�>v�ğ�;�$�i�W��s��ky��m�?��1���������5�E�W��^܇�Z�N<�cT��}G=�����W��:�ݕ����yp.������<���L�]��/]��5=Tz*#��f�Q����`ܪ�v�j\���p֭��8s��������N����ng+�l>�z�<�W�UU9r������y�CO�G���	��8�d���@�N$�4aI6���Ն�q���:��}�����=v��̝d�	�w6��03���۟o�͙����_7��I�8ɦ}I=O̜�I�;�0�	�w�+'�Y?ei8�l���'�Xu�'�~d6¿2u��9�Y'��:�����߾��Ϲ��i��	�c�d�O�<����'�Y����|�����N!�s̒�a0��aY>J��)8��M����	�O��凭a6���|˭g}��zs=��Ot;�0��a�����Nx=��'|���T1��}��P��S�a��u&�y�T�&O�VM� k,�����ߴW�Ty~�A��¦�̝$��W��~`~g�~xɦOP鿲Ax�L5���I�X~�0�����ri'Rw ��OPY��)=I��~I8���~���W�,(���~���3����8t�&:@�N2q'��|��C�4�ɦI��Y���n}��$Ĭ?s�:��1��'Rq!�w'�8��V�!Rz��?h�y�կ�տ}��9�k;8�|ɭY+��oNY>�q4e�'���,4��CI�u��N0�k܁�4��/������o�O�}DMC���B?|3��^��{�4WR�p���·�8��V7���4k��N�k�2J��q6�i�'�{�8�|Χ�?0�	�j���N��O��>C�'/�}���/ؑ�ݡ�a�����x�<M2O��9�Y8���<a�O_R|w�l�d����'�uI댟�8�e���M2���ԩ���	���	 o��s�Zu�j�Yu���޵��qY<A�r�6�s�u�I<C���s�	�߰�'Y6���]�2|�����VOP?{I�Y?0��d=g�N�����ԩ�g�����^�v�����x��VVs�`��06&�+��Yj��lh��u�nS�@��jȬ/,d�s2��\Z�c�X\�2�<�	���[�d���az��m>>p�t��7�u^�'r��aW;��!+v����`��i��(��x�j���8����&@;ʄы+��W����.[��p��謰��R[���n
c!�H�ƌ|0in�6����y��돻���		+2�y�&�������r�=Rtn4F�D����/+G-�y���XK��f���w�m[M�����{0��G����G+s�륎]���D�=�k�ʓ��L����j*�"ũ,�r�S]i��Q�M���s�Y�ʣAfܣڝ[���Ɣi��k쾄��p���%��Q*���
7���;��F������ӫ
ך1M#o0n3�)��V�xV��[ ���v�����m!w/�n.Ӕ@�|8��dE�7��c���?&�ZD���K:�)���zl��k�Yc���o�G��Z����'ѝO`��7��q��Ɵ�|��3'V�`�K�ťcλqd@h��Cr����x�s��kbn�;OJ��XRqJb�5؋"&�&�V+�ˇ;YC-`��0E���t�R�4Fj|M��B��F,�u�2* �z����eI��͈(a�C�w�k��x�vB/�ai�ĩ����֖̺W��bY�-� �n�A��3�m�����7z�mn�f+�3+�[�i���\�l�mh�wuxsn�lߏ���F+��u��]ld���A�94
�.G5^����E�e�%��Aӯ�d���L7���uy�:=l�����.y�5;Ѯ����|�^������W�p{h�S���{�,����Ƭ��5Jh(�����j��^�M?��;x��$��oS&WNy}�Y��S��X	k�/�8U&(�0�|��uh˘�"R�Fg�U���JIX�Nnw����vAAx�����ܔ#y����[���`g�u���Ç�	�����4��|[Pfܽ<�Bt=׃q��gJ	����}�.�u���J����6��:bo��2M���n�8�^	�m)�z,��LT�����^%c�^URɎ>��zݚL#�%���'-����Ɲ�y/2�~bn��I]�f�};*����r�f��s�a�"|.��̪�$��CN���H4�|g�Ǔ7�:�k�����+t�|���*�;���z�Ʊh���x��э(��A�]վ�z�h�oIW��eݚ�C!J�`�l!�}q���̽Џ��Y�F��R��w�2,)�NPD�芩�W�~�ۛ)��c�ޝ�F����c�s\��@���vi�I�-%�hN��׊�����e��<\M��Kp��ru�Y���;;C2p����	:m=����D����z��������.E�V�V-E+�Y�B�11��c�,HV,�jE�QkYb��E�)�[U��«�V�+*(�m��
�V� RKl�`ڱa
��FT����&0�Y.1�
��[k���&"ʕ��Z�Kh(V(��YE�dD�aZ���Ƣ�Ed�R�U��P�KhV*
[HV
E���Z�Qb�Jъ���TPR��T�q��2�UEU*�[J�a+XT�B���+V�����P��ʆ%*�U ��+%�Qb¢���lQek��T*�E��5r��FAJ�+Em�a��*E�*�	�QOݻ��]^��Ţ�XxN�{{<�M�^d^��b�d������hw�M6q�wF7����rݦoع��<��_W�Q�s�������YuJI��I�
��
���J�{�	ĝC\��Y��7i�M�0���u�>v����d��VJɦ��|���N3��5���ܮ�������9��d<g���f\d�Cl��C����C��J��7���'�G��
P����쓬</0�'XOzY&�R}9�?I���|_�|y����o���y�_<앆��Jɴ�2�8�2m=˟wFw7��Hf��8z	nj��?^*|z�A�sBE��N�|j���펣��is���6�?B�7�\�^{�m[����M�h�~Y�p����a�핟l��-m�;3��Ⴗ��~f�`2MJ� ���w\.I���]��	s�t�˟ZAf�u�>͍89���vǇ���w�����pw�K�˒����t���qv׼ {�#��]��$�s�ɓ��J���{��&ؘ'��js۷�Z�j~!��lgs	�ϰ�uh��>����:�n�[��2���������x/!��B�`~���x���=ه;�~%�#A�
ׄ�Y?xA[���kOn���ٛ�� �/�{�z.��*x?$���%b�� ���ٙ�AN�7ZBq`�Myޝ!����f�usq�Eg���	/fd�aa���ؘ��]�)�x�z�A۲mεU�ѷ��Q�.IsT���駑����_UUC��;�Z��t��:S�a�z=�^_��~}>woη ����z��@֏M�]��˝�u����l��+o�ʎ󷀵2=�|�ٔ�~���~�|+r_8gJ^繌wf��9|��u'j�}ũT�b�>��y��/��ɻ�L\=o'������s�n�n����aL���G}�{�&U������8^ۖKy�w��$��m��y�����T�:�)�`ͫP�T�_k������Aj����3��[�eh೟�q�lE��^��/2�v�	����*�l��'��:�C)��9<��=C&ds"��q�t�]n�P:tW�c������N��#���|5����J_s�`����U7��l	ع�9�:���\c�jk�������<�'z��?5���Ϻ�������}w��"|3&vp��t�|3�W���Kc�i}Qhx#nٺYL����m`0h\�K�|pd=�a����a
��aB��b���nx, οs�|�UĽ��v&f��|�-�I�`Qs���y�j���>̇��]0l�&���Ήq۲w=K���q*{����	{��?A�O��of��g���.C������>צ�Ko/��W���;��N�����@(�����]��f9�j����Y�g��?I%J��9e�������Reږ�����uF��J_7�&�t��(l[��;Z,H��&ؗR�xL��G5�Y��O6�(��z���;"�ލ�%Xr�p<;�A�I��z4L���CĽ��W�[����f�.S�1Of�6�_?N�ӂ3��O}�qϲ�"_B�-sr:��-�3l�B�N`�z�Ϸ�,�k����8$����W��/�Y�7D���P��>i|c�������V���{T��f%�r���ʾ�w�ݞ�Z�}=�7W�@�VE���s���n����c�}\�LZ;��$�8� ��o��7r���`/T���+D���0�%�Z�/!�ya��V-u��h�;��a.g9��W����w*�÷C���)��s���ń��xg�	x���@\3iz��ԕ�ᢥ@�����kr)@�$�VF�B�L��S��`�-�xGFqB!�ڵt�m9O���:d$]�}5�~C��	��玪LG,��ʝ1�=�[��M��:�/S���JS��}��C$��}HO����q��t�1��>�s�[|��:=
��Y5}���w����ۭؔ����OgނP�o{1�״��%Cx6��L���&�䬭[���am��o��.syܻ7�Wf�{Z-T�1�uw�rIޭ��n*h�u1u�#z���o?\z����5�[Y��v���G�˔ܭ��Is�k��λ`�0�����.�ލ��9�Ԣ��M<�vcU�n���RlT��u�&j]���P��s}����qٻg�<o[�Os�x[�nd_s8k�/�D��=C���7�k�l��g�`Ԟq�;�u���Bpv"�W���z��C��1�p�u|j�;�~��k��w��p/g@���֊���T�+68n��}����v���f$O��Cs��|�NGn��~ߜ�*��u;{�|��r^+�B�8r�yN�����<-��nT�c��)Ӧ�����@�a~�6q��ۆ{뼭��y���:�;XGD�.zՆ���͊N�-<��?U�朇� ��0bs�����V�	�*�U8����U��ݿ:��ueu*7ƧY�y��Ʌ���E��;|���_o���\^=1<Z8{L���+sF�e���݋�R��2vf&�J]|t�O];z&�vz��y���zl���g/{���caL�����a!=�c��uy1�X�}޵�p�"�l;�79Է�r��I�d�f�}��]�9�Q�U��W�����z��hp�x�o�:p.?z�"��`K���RU�n"�g���0�l-�ikS��-��=�rn8P��Z��;rI�{ֱ��Ijo����V����{����(��d��^�(�>�y�>M{�7=���f�`���\������^�K��P竒��!7��[QM�x'��Ӭ9�+�2�\��K�a��_.}v_�G��]��u�.� �Qy�U��.5���dr5:|�@�ĥ���T�_p�bf�̳3v����s��Wc!&�r$�El�rA��9��7S��zb�@ܓO>w�v�	��c�Zs��*��E ���`���oZ�{<�|>}�ܨܕ_�x��y�s�_��;��7������r]�V�w�P9�&�ե)
�+��Prf�s�0��z|���T�)�	+�ܞ�oy��@gh7R=�yHTd�`3eX�+����n�M���)�ڭ�4٪0೒ؤ�C��+�_��u��K�)=��9|�}33�}��:y��P	x`Yw�=��,�F;�GKx;]⥨1ްuyr�\9~��C�ҽ��ዊ�}�0�����=8#;���a���<���3S�+�A���G�OU�v�����BgJ^��;� 1>O���7�9;�3]�:�4{�l�/_�ǽG���u��^��ҹ�7q��vQ�ge�9�����U���H�^�y:�1NB_$2v��}-�^=%���Vl��_?5c�
Rʇ���m�;e����y?�f�W�gob�o�
�W:EJR�R��7�cʻ`�%G0�{:����j�NM����QR�o�</MQ���k}��!g$f��\�}s(Hv'x�wzItqbĈ�3R�,+W8�;�9��Q'�g�0����n�>��������=���;�&�k����t밓����coz��W�1w���\�&#����05'E�����vܧj�[�m�7[�T���r��|윬����ֻx���z@���u�(s:.y��OQ��7�>O�
O5�M�g�}�eo8s�fw<���Z��.�x���:x�3ǫ������볦�O8����L�2^�":���}�v�ɲ���}�io�n��[�]8����;1����kk*�i+�v����:�=��A�/FT�bXC��qӁt���g����l��56�f��L�z��N����l���F��J;�U�}�i7��z%�G�����ȍrU�-�p?_A�wN�;�D��N�U����eCM�����7���s8�8Xs�N��޹Ù�J9wvj���������ʺ�����-�ң���vؖ��ĝ�a�((�Ga�F���*��+��Ւ��$,+������"����y�/ASF8T<��:���X�ƶ����7��<t�^�'���@mI9�	I&��{S��~������^���{�������Ň�Ƶ-�4�����~�o�=�o�)�O�?oc�|.ǃ}�z>�pg>�8�S�~��=ꕷ��I{Њ��;��+����9�k~��	�i��\|�Z�X��'R��c�cZ>�U��Ֆ���G�5q�^��9�v�̖o��v�K	�Lp�0J�~6Ux�cجÍ��Z�s�͉�Xu'���mO?E�|;N���_�Z3��B�YӺ.��x!]����ټbWIј��i�XsŇ�������k~�*�)[�_
��_^��)�{=�nj�����ܾ{٬��7̚���k$���F�as�}]c�?`��;��޹뻮:Vbڃ����=�뺜��N�_4B�>w��Ҁ�u�����Ǯԕ���OgtF�>����J��y�K�n�V��	s\<N���n�W{}���}�/�fwq+&��Gwf��[�c��l��꿲���a��a�ա�*n/u	�1fs����L����eG·�N@���n���.�z����"��.UxbW2��w�!���ef��ۛ����ѳʙ�
�t�w��4,j��e�b��������g�����w�?M�8�;K��J�T�r�;��(k:iM]�)va����s�����ǃ�n��F"�9x[�nd�d�[ӑ,�}�7��58�Ij����`���kF�r_�S>p?px�;1ы������h�H�{���c��׹;����I�К`U�0x���{9�{���+��mc��9Ԝ�9,�����U��1�g޿3�ލ>ۜ�
�q�=θ�P���ӂ=��^��q�g��r��t/*<����'���w�nS�{�m�X�m�����ݓw�^����%���p[��lӯ[�����v7fr�ak�����t_s���o#�a��#:���&��d��guI~7aS�4���k�H99}/���{_����|�탈^�����s=�93\|���a
�Ώų�oI�8�h�<Oz���+JO7q5�`�NL3�c�t��2����'5��+i��ӏ��R1�.�(�zZ}3q��`GB��nF���Y�X/p)�jѯ�&<X��|��M"��
�jnʔ�.7���c���̄WP��6e7us�s�������}������gh�����K]��͛L���x���L^&u)����׷���k�ʷ%�����sOm�ns�W��0�T��q2bY~�qu���X&of}#�ֻ~tB�tP.R�'+Iuv/뷳�7�)_��}�s��ns�ϮI�S�C�/�.gH1{�C�$�tf[���D9W��76oW-�͗��mw˹.�"��g�q_U�3pG�u�����Ԧ�!_z��`�f	W|e=�`��<�U� �5�������o�f]��u���z��V)�e�=������;�ɛ�oj��f.^;+�z<�;�s�%�C}U/��c_���f_��;�#���<��V��h�<�UZ������5��ח-�9���n���yə��{u�W=~3��A�;�.v}��/*��:��W��ar�yfD��u�=�ZU��Ohѥz���W��5�z�Ph�o�I�����N�R�:t�� y8us�/���9#�Gy��	��������[H:umqSYem]9��
�D"��!{�t{v؇L\D���W�uF�,�5h�ou��u��n���'�܏��ƙ>z����ut�Yܫ8u[Ȁg5�s��|+dX��+���&%�N!���?/{k�xكW���胕w2���'K>������s������/Y>u���V��o��γn�np1����B��M	 kyh�*�*2>gX�鼩vQO����w�R �H�Z#A�ʷ_n��xD</֖Q<���±�
N�2��X����\��2Օ�ߎ��i���$��4>cp+U�a*���DA�R�ƅ���E9p�	�)��$�sv��)�"��p�����9N��u�����At]!�ɱ�����\�Sv��w�x�N�@+��M�� ���.k�!ŕ{ћ��)ؼ���M6{�3׵=�I�|9i�fA��ݖ�T%�O[�3c�x$)�u�e$E;g����B�`ӫ|e;u�3ѿr���xg�#|�ɕ��Vĸ��u�(n��	Z/&����6��HP�,�ͨ.���d�7��2W���������\L��O){�ˊbl��
↭�ݺ�9�+����6�� [���gg7�����#����z�*����=Tl58̈U��N�r�����F�O��4��j,�9w���V։ѕ�2N|&f��2ͺ3���Ě�]�������tf�e�s{�6x�:W^�S����o]�Ǚ��}��Ao�9�ide�����eކ�¾��f�L�����i���ɫ��7�����o��U�l<��"���q���4�9Z�ɋ�؅I�܀�gU񮿟�����c�چ{ϖ���;�G���n��a��*|sHf�=��dR��4�-|m_?í���VF�'��Wѥfd�`�tAW֌����&iC7 ���fmmsՎ#�
���Ja?t���5������>B�,�@��xܧ\d�����PT#��7��]P�,���]���m�p�w�W]/p\|����l��,��ݮ�/`n���"���k-�����/>�`ʴ'3�^��p�$7�N��]�Tn���G�ɷ��_aR�9L\�e0��+���g-���η�b�X	��n�)��}��㾻$����*�O8D�}�������m�,0�+4�ThW��p.])@��fS؟�n���Lj�E���$��D��S�YM�lwqS����s���r���ھɄs�6���Vb2b�}T��[N�ԅ<{���{���2���U�4�y��hD��Ħ{Z�T�!^S.]+�}���^�	����6F�:A�B��r���y�}������ �*"�"�������µ�ZѢTQk�Z��e@�KJ2���bŘ���b奭��ʋ�
��+b�A�VVڥAb�J#X�)U"�Ԃѕ"��,-���kD
�Z"�KE��,����"*�+%*Z�DQEV�+Z��R���R�H�T��V�keA`��TYYX�YR�J�
KlUX"�-�0J�*��H�ER�Kmkm	UP"��IF�R���Qeh�ŨPF�+#l�"��VAs%`�Y�VA`�j
e*0Rڢ"����KATjV�0���e�jQ�EjR��TXZR)[��lD�R��eRT�-�F�V�(��TTZ�B�DF�*"@EEթ2�P
"�4�+���|
�r����zs�N�v�t� �����[ځ�;dXHD/��f�wf5o��o-����g$��������}_UzGxQs����՝�VuoџN���g�'^��'�}�VM�c:�溝0���H�+�n�i���/I�^s��=&�{�K�2NW����^�zo�&�|M�Ц�G��h�vy��ۖ�^��z�c�}������fܓ[��<hՍ	�ʇ������/�ԕ5��e�{�{yɮm�\�"��5�s�6n���~	:	z]1��<Y%�%��|�������q�x��&����i�A;:��t��;�4a�g�6�Й۽�����x=�s|6	s��~�lv��]G��4Cx-x}}ރ��a��Wڧfq{͉�aL�\[w�I�\r�zz��\\U������QY�>#������Y�w���I�~x��(�E��}Jv�kT��vFk:it�	�\.�8����^P߆�{^�<�3�f�r��~OϬfL�Deƨ�YY@@��>����Sղ�ғl;��Z��w�i�VD��Tku�#�-���[�m���n�����E�ו�p��2�M7�m���{�3"�O`�-K�zi�
������V��s��+2�}ݞ���%��9r��m��>{�$��*M�au��M �JB�X��9	ܵ�"oo�vh��3�β}&F"n��	u,<%hۥޔ{ү	֍]Ro�����y����8�rV��n����t�������`�星�vo���.���]:��nf������?����U��z��x������	R�	�j��+��6���L��>ڹHg/;��F�[���>�~[|��v�y��[��'�Qz}]:3DpTc��Om�9{>n3d~�y��֥y��hq��}5ДN�-a������OZr��/>�K����;}sޱ0��� �F������ٛ;#�	��[<��u%�Q��]͚l��<�^S�-և)�Ύ�g�{hU���[6>�%t�05��s;�xx3
C��VE�5g.�%&�A㻫xj�2���5�sS�8e��z��r��S4�ҵ����n��o]'�����B�1��q�R�Z�>�>�C���۔�����u�eG�̣�gyb�킰S�CTv�؏#�]���n��������}@�������]J��l�����%}ni�5>�f#�C��6f��ͧK�M[ghÿl�\���Q�8�M��>����U�������{��wEڋ��m?��!Ҿϳ�o/w�w�LҬLu���U�}��y�#��s��s��/�+���J�$�5p��!nz�ܽ�nM�����;�K����U�a�+�gH���|��j��G�О�+��x�|7����aˏ���C�o�)��;r�u7�xJ�>]�Kp]dy�9 CRw`�p)�0B%�NW�����f���ɴ��u7>��Q�vn�h���X{������zVlq��k$�ӏкe��f`緳�����_j��G=�Խ���qҧs�{�E����JS���L��_o��S��f���w��%:�����{���ƥ�"=t�le����Nn̝X�e���3�Y�y����4�֎9��q��ñ:S@miw�(ۋ��c����N�u�(w���5��ZOn���LxTڻe�]nշ$�3�}w�ɹ1��ξ�1�D�,��� ;�_�J�Q��g�1�o%�6��l	�=�	;���/�,��{�Y>��x=mk�r�)\����k��ד�u���O9�𷻸����3G<���j�#١�~,��o��h\f1��pߛ�J{�w��;G��<�:����ZU�Z�Æ�p��3w�`�ĸ~�L�3�s�+i�f;̫'�U��N9��;6tx���ZZ�W���1&#��n�ó	��&ysN���N�｢��z|��tE��ͺ^[ �iY�c��&�y��������s�k��d}:�k�9�\���I�K��Z��|�������2r<Cь��Z.r�QGҶ]�~�Z4��*+��R�M��2fG�3��ڐ���/*��Y�YZ��.���ٟw���'���",�E��3wJ�5�kP��ѡ܈�Z���)�v�ma7�zxg���?�%�;>;�Y�!�����8�*�:n��eK�h��w�t�\�t`\?Om~�c���ЭLx�_��l��Vp�j�]��A�F9U3���G�S���^�#:���7�*-�_q���2-�s�W�VT;�<�V�Z���T5�u=J�n��׹�������������a��Ϫs�C5��`'\e�C���A���[��7�PI.����Euk[��*�%����+�4�g>�&�<��.�G�䤸SQ>8]-y�7V���9z��<��#���(&�4l��6��L�01������M�HG��i��<�H{
�v�}����E;i����V�d9�^,��#��6��p�P{cu(�K���B���^qx^m�3�fݘ�s��w��PzV���_�wR��d1���M�.�g���LN����5��i]#��σ����x�z�!9*��J!�z�!&�z�1M��6�OiZss�K��%q��AV�e�ƅ�X8}�ĳrٙP&�s�#LW��:o��Cq$�;��β��pU�Yh�v�,h�qT]O�Q��6r���Qh��u'1���R�(Z�0��i�o�vC�)w�Ƹđ���n�줕�#zk=H�gK~�|Ä�J)ޖL,�P�Υ�C�q������^u� �w^�t��������)Ť겎���B�kNU�!�fƊ�ҵ1X_N��nt�C$#6.����RLF�O��'��Z'~�tY���˽�f*�1��	�Hs}�������D�H�O�0pe�s�;[5�;��s��zh����ogKY�o�}�}_W�ݱo$�� 4L?�Uo�b���r���b��;F�,�V6(q��34+��W�zs�����7��e��f_U�C�����k~hq�nz���86��<O��?
ǁ�,f�K�nPx�m"6�wh�Zo����(S3Jk��4�uO'/NA�^�����{ms�)	w)����1�J��, �� ���kR��t]�������~v��̎RVr��kt���{�V`xeH��衽G>�p�	�H�h�=�iX)tR�]���oV8�n��1�=�^1��,Ϟ�ە��.�p(|0�}���a�}��I�OG��'fg�:�m���5�_��z���%aʄU����(���t�˸Tǧ���K����:�G�Z�d�F�����p�ʲ�-;j�zY6�9c��+�hX��j�1���zq�a�Q8�Y��@^*�~Q{ǅ�3�/U+�Om٬��oK@�\K�5wu���+�J�XgX���a��yb�4��|��G�>w���z�_�T��Fצ����ɉ��δԺ�]c5�����r��/ԇc4%k�y�K�}�zj���+�Aឍ9�W+G3L]�[.^���#�j) 2�ٕ0�e�N|��.+$W3qI�M�<k[�G*���?��5u�I�P��i7����ﾩ�T�!���9��>?�������,��鮬f`LtK����Yq֊׼�zQ�ٱ�\�z��J�fp�s�0�'5�#jP�[<kǴ�-/R��}ۥ{��y	e�M����e =NR���T��%ɮ�qXw.Rߐ�3�c&]3Xo~;�W��g�F�Y.H�K�9����������;��|�V�B`j[9��C<��p���6�T����P�*��_%�kk��U�Ԫ/]܉�Byg�,c��^ھ�Z'�|��7�~��Z�;�i�;����4\��%�L���:L��<�����y��r\���ǉ}�U^�6�}8��=n����i F#���o)���2��^���n�9��w���RV�{�c��9�¤���W�������D��Ӹ��9�%��
���������2�J����w�z�a!�N����ǎ/ß	�Ho�)+�^�Y8��y���]����:���5j��>Zx�nd���pIJ׆,NCo?%�`v����Շ�A���O���͉�yO�:�y!v�sYQ�c}�XE��n�	V�*}T+�E�ן*li�4�҄�^�{UL���E=�o��v��^x\�wh=�[1����/ol�P$����vӫ\!'��91�R��\&Ǟ��y_��|>l�y��3���e$��H�,�\EX�J�D�h�g��`��r����+=ǭQ�pՃ�}����H���?��؈�϶��]/-�T�pL���/wKE+�RiX}(��SF�y��&�P���2Li�T$�Z�
�A:�/"3h_"�o�zCY:��M���OF:ں�^����P/ӭ1w��;���x_�b�t�xd��{C
�Zמ�
��o�i.5��ku�|�d;WY_A�t��e��n�=��Ǎ�Za���֩~�q��ySe�n�U�z�cۋ���XΨq���k��>����s0{�'Jy�;��֝�ǋ�e�������h�U��)֕c�@v���_�t��r�?5-깕v8W�l�K=sh��j�L�cr��/���z��N���`��G~zjD�z\ �T����u�{Xs����kܳ谳2��!kMlԝҡ�.�<o--���y(�*)�ֽ�;Ѓ�Ug���u�	���c5�`��E���O��.!�Ds][RL������8=�d��O�Tc]Q��>|Ӭ���wp0�X~��-wcm�4�YJ�Ԣ,+����)>ƥ�f���5'�ث��d(fuò*�@��q�P3PX+�u����6o�k��w�.\E�nwK�;8�,=�+Dq]{1�~��k����M�u��N���`�îg%��P���F9ࣟ	����S.<�,��D�r�#�>��w�<&J9�7y��t��=am �c��p�en�jf���.P��CQ��}G���y�3���z���+��Y����PL��4���k��ܽ𧗧)a�Z�4�B�G�z��MA2��wop{l�i�2zȦ6Y�%\������UK�-'8�z��}Qakn4%b����{��>�hKZ	����wI!��rI�2�]����5s��en�\���Y�4���gt뷈�����4N�)�1/<���^{Kl�{N8�
����F��yh�aZ��}c{��m�{6`�a�H����LpSԺQ>Ь�f�#�;Fz�r�z�i��5��$-%X�?\�����8���C	��Bg��O0�t#<^R`���%u9��.�ۣ�B�?TB�xL9qps�{6����AC7�^��jFB�C͢������Ot:���f�ǆ����yX���A�q������ǧӒ��XWt_���f畂��0u�X�h�JKV���Ս ��v�ר�KD>����MS�
���W$e�3ޤ$w�o�g������-�.Iv�'�-��&�lM[r�LylK��|�3����[�#�2W�׉���Gp�|3�j�g���}�}�W�x�����6
�FI���� >S]���)��VS~���c�U�����%�o4ӝ.d�]8��e�-�m���
>�ً���"���OČF��/�]B���]v�J�^s��q����`ɦ��+K2�ws�>��k���읐��֋6�2�m@���˝��
�7C�X��evD�
��z�Qp��a�����R���8�����2�n�>ɠ��A�����t���cI.2�#�
�l�hdSW�Q��G�Ggy{�6�c6�"<�ܓ��y+`����֫�:G���Ŕ2��v[�ߝ-�<u�R�y¯}�Ѿ.W@�h��O
��Z�v�#�2��hN��"��8)�v�OX�]�	��5(ez[Q��{xp7F�;o5{Y��7����~�D~\��	bP �:Ԯ�5��
g�*%��qYA���O�&uk��}kP�zƿ}+3O{��b���p�%� �$kK��N.���]�tI1^���S}:i^���|W�����`Fܬ�?.�'��a��eه�#��.���Ӯ�d���& o5�����e��1>�7v��K\��ʁ!Ֆ�]V��$x��=(�iK������ih�i-�+C^��>�s�Q��xgl��=�5�@���7i��Ļr��-��\.����)uj������o(Pm]��׆#J��W�nI;(v(�ʽu����Y)0��D�g�day]�D�i������5���]�E�Z=X��5.,�ʕ��� ��V�Hŭz����4���<^�w�R�̨Ư,�M�f^��7��L�FsḊ�V\��in
����F���k�Ġ|t�
�L��}�|����rIn�ȹ����o$(�ȯ������˨m��J������r�>�/Z%;$��[�-H��6U��6m��PO�������bC+�[��	����'v3�. ��vu0�c�n���oA1�.j��<�un$�ۢ�����s*�gZw��Z)��������&j�ul������%�[)��#t��,Ĵ�:�F]Il�g+X&(F5:�����\	�3)�(!դk4�!�jP���d�[2��]vJ��`�fQ�[���!��v:fuS�Y5~XA��r�=f�ty̱�$����Fv@���5�}N�跩�r^�ܠ��˛�8�F�Ewv)}]t����g]k	��[wnb���2Nt�{P��A�&��GVl�LY�\�:��w�maF
��F�J�j�)����u��B"�т�X^Tt�]�¨f���s�E�`��n��r�h�i綈��l:�x����o[��r��E���`v��y�(K"��<[�����F�3R~�﷡#�-GܾT�k�!)�GL,՝�ۓu�Wa�o<ItV�*Kb�%jqb4�����-����?����o���ZP�_��"���0�NA^�{([|l���WNZQ��$N�<��;y��-p�@_�BN?��]-J9~��^��ZX70*�s=�r���Z�FgZ�3�Uq���[LXKC�֜�m�wN���C�W>�Y����!�a����3P����ywn��q�u��3Pz�2��;�4y���f�A�a��Q	jgl8�[�͕�^�|����0dT]���(ms�i�]\�Y�V�{�բH	]���H��G���O����Z���8+x3�wHY[:�Fb��޸֣ؓJ�����b�LG{����UѐPy���e�}�j̪Ft�ۛ����(3"�1���t�������(Kɷz#,�'9�JX�Ρ�O�XFu�ѷfr�z��vX�u�ێ��;4���zuf�[ӑ��MDoҜ�T��%D�,��*��Q�")��+b���E�Y�ˡ�Ř��EK]�Gͤ��e��v[����j�x.?Y���a�9�_)���Ĺq}���ҝ'�%㬰3)N�
��7V�듸:����Ͽn�y��g�~�,PX()Z���B�YY��)Z"�[%�eYmX*�P�.``���[���ʊcK[)
%E+Q@̡�
�ԭ�j@�E����J��kV�(�*�,R6ֵ��QF,V.&&+�T�F�U`�Ym�6��R�����+2�(E\B�bմ-�-eDT��\@X�Z�+TU+"���`",e�X*
�EDb�!VءGC+B�b!+TE��%aA�+TJ�EP2�d�0�B��iEP���I�T1�Ue�al�����m��1��T.f���e��r�@D���J"�m*+�qR�-�e�kZ��*���+(�խEQR���,+*�J�m��iTX��KjԔk�Z�*�TAFЋD�
�#*kb�KQQ�Z�B���*
Ұ��@m
�
�J""��D�B!�uHvS}j�|z^.�z��A�㸵�Avu.���6�ko9����Y'cQ7�l�sx+<�.�d��0{q�=}U{S�>���[����B��)2��>���~�]����I[��s1��9E��N�������{�]I�ţ�9�b�葆�0�/`�p�����Ӷ���t��(V�,0v�q��5ò��e��ח�ħ:\��x��h۪xEB7R��e,v��l38.�����.mza�q�&�i�D�Oo;
���?C6�j�Ї��L�ږo9x��R/j���5A�H���'y��um�����*:^�h�M���#�=��e`��1���O��a��O������oLͤ��9�CZc/m����^>B�d�p��^>�٦��E�����W6��l�~~�v�2�d�]G�z�Q`w����}�-��2(w��#p��QG}dY�$�M��g�񞈳�,LIh��~`'�� {h��g���fN�05-껺�j��JO�&��JL��sUlJ��N�b��JEh�r�U"G��hO,�zQ32:	R�U�:��6���Wu���w,8���*��8���s�)��qt�&t;�5^�K��ZhY�� L컷xvQ��΍w�!�N=~�(�Fچs�R�y\�n�w�b33�i󣧄bk��⯰.�T���y���
�(���I*v#]b�;�����c�:�-!D�v��l9n�{��df�ݗ�����5?ź(P���F3�+�� >	����0\�K,�y�=�d���d�7�v�eQ��ݠE|Y	<��(s���jo�M�.�V�7�}7�N��עU�"���Y��.y]�f�J�L6&&��$�K+�����TnsD3���_�4Ж����(gpuy�w�t/S�Z�pɐ�ϥ�G�*������3ޜ���т�.J�Jȇhd6����0m\X����cNIJׁ�Ky��r��-�Qu9�;�-T��U�-툓�H�myh�����n1�	���B���פ"���o�n�����noG����T��tʞHO�e/�!�g�Zk�����u��߈�P��ؕ���xd�N�l�j��.�8:Y���և{�h�'���U�~��#GR�`=��4G��̶���/��O�J�J����{�&.�S� ���'�mq�b`��ay�F�,S��<&M�|���'y��C²��M,���v�%�<o��oc��Z���/{N�i7V�Uy�K���d�lc�����"�]�9�<\M)�L�L�!s��JYD̸r���f�OXn��:����K��}G�ˡ9�5rx1j��|��N���ٳS�	��,@���L��,��u ��
״�>�r����y�m����������L���p�u�|������k�:
�{�_GcQ�V�-t��l'�����R#�o�$�&g;��������h�zG2��V��j�IcpVZ�`�"���z��)���\���)�w=Qա�Ie﷧�gl��xE��Q�	�f�l�� t�ρI��l���\�����~2���3���U�8����&d��	���~�ְt���]�ͅƸx��hh������W��y]�����N����L���ld炌��� \z}��9,�90��z<��0z����Aֱ
�!�DF>�ޘ\��f��,)����C�r�Z�
F����䯜<�:^Ӕ�3�.I(c[A2*��|�OSJ�����i��ê��8�~� V�ᙼ��i��x�`�5��49�<�juP� K3��z�S+w�`{�"I:�,r��w��������-h2�#D�B[��K8-%��h�K�s�Sp�L
�����]�ܺoxJ�x�	�h������m�OQ�B�%Q��hN�{�O����i�難ઞ[���Ѡ���s���i�S��o�u�z�n�b:���92�GI/�(�E�-=�_J��ES�g��z�Tw6�ZL�N}�QF������K��;;<�>��u�.��Km.{Y1��W�_K�K�ǡ��Ǖ�� &�O{y�/z���r�W���.��H��2���.�O����C\���ҭ5���{~�W�e]JXs˭q�3�^���5'�P��lp���:NhhJ�+ft��� �m�w�Z�z�?�o���ϯ)�ͻ�^׭@y��/��X�=�ңXcA����8���\�ny�$;�sn���?Ki��X���A�q�������{��K^�蚾3&�vF��2��/u\[�Ou��Z�ł��e��UﳅY`����U���Q@��s}�M�kؔ��%�ý(? ���;�rT:���̪�������r��.�+3:zr1���r=�7�#���`zi���g|��(|�c�>������{�Z/��~�=�i�����Q�:���^��B,V�y����Y��a���Ծhzq��ϧ{̳|�S,mNs$9�`R�#`�[X*���uDu�[e2.)��(�ye��s2��)���7��o��P��A���`wk���#��\\Hf�we��?!��nmhꠊ>�����j�0k�3Z�ϴ�Yb�k�#��k����!~��C�بH�*&fu1`3-�C��Wk��[G%��d*��v�"$<ZR�3y��ˣ����٘ήa�c�،�6���i>���q�Z3�u�:�������|�Fy��OV�/%/��)E��DWm��䈫�L'A���A37)����K����� ި��rMK������u�O��g�NЖ�C��Ik��B��%{J�b�T�3/���J�KP��c_�fi�Sa�#����d�`�$k]KF{�?a�̾R��ݭ���\a����{�uf��ȃ��]�^�Vtb���f|�x�b��0H{۽VX$u�3�x*n87H��}�}������ck���|2��s�8哦˾;�b�D�4=������,Z>�H��R���tS���/'�<c�ziղW{ο	֍�M@^g�K�&8*v���"4��W��y����b7��C7t�j�{l��Ʒ��yu�	�}k�kڳ*mK߈�C�T�A�G��N�P_@�֨�>��j>:�<G��=�֞��v[���<�,�-w�	��O͝r�$!���@�
�)\]KXt5�5�#�\�;��M5��Oz��X���Wo�T;�4:w^D{m��P�D���oj�5ۮ���/�%�?Q�({/��1x䡗,���L���͒n�]��{��PFFn�\��=�s�fs/+xX�/�(���e�C:n�S=E��0f�;0j��#��e;���|��s�#sś�����ʦu+ �__
�ME���+w3!�T��Hz�Cb�޵Ūi��U��&�>�.0��J�|�;��bKG���OixU-vjJ>]q_Wv���̲Ϙ��Y�w��~����������ʺRT4�KRֳ����U��v^;�98О^k~�U�k�/�b:�&�s
�#!�������S�x�>TG	4��-�g�2_`�~[�t�F��e�����wZ2^�Ｑ諼�������oKχ2�z��;��Y%�L���oeǸ��r�{����c�^�eө��t�c��9��}�\�d�r+$âa�i祟xt�˘7������I�i}hP�Y���04L�f�*/�������g�����ط|*�M��<����.J�J�gk!��}gV`���^L�v4�,׹Yc�y�Ƕ�`��]�k}br�<*�I*�H�,�\E]We�����4����i ��>������y3���dD��q?�˰�d�K��@_^���"��V�{���A��c���&e^z�����w�V���8 ��.q�����p�ئ������{��h,J�q=c��T|��V���� B�J�5Խ4��C[�Yt!3����QVx5v�y-}�W@U%�����wą\Wj���i�9.����B�ڻ��L���O�H�ӦW�&�pS$Ƒ�<�zאy·���U-��P�@{7}����5�j��S�{��gJ���a�x����ߣ�E�^�M	�v���[���{6@ݝ��=�^��$:����||!�Z^�iOz��c��S;}T%���R}χ2���np嘘 z��=zz�׵�@�����3��q4�k�kC�6[�C��[�&���`���U�-t�+���rsl�"v= O���:N��L�/��VΧI1;�<��w���W�(�.�`������K����Bq#��Q�,B�Y�K�#�Ġ�p��;���{C�q�r��1]-C��ث����S�ݩ_�7��h"Q�ݛ������zj�ل��cL8���}�8���:y�83�m
���3���y�!9�tH��b��wS���L͝h��Nx(��[ޯH)���(�/����U�[�Y7�,=����T(mJ�D�]���[�_�)��鑕�,��z�W��6~�E��$;w2��ьk�&痞��n���n��@ἳj�!B��qM�F�oWa�Q_�U�ኻ��"�߲Y�����A>�&=������n�nV�X���^,~�x*4��R�*B򝖉뼧��1$��#ο�}�T�jl�ӽ7<����+�] h9K�I���L�ƃ��P鵟:�}�;�u�{�����ɗ��v�^[� �T�,�*b�~?Z��H�I�]��=~�K��/�؏/��8����^X�Ή���v�xJփ�*L%����5���u�^�z�*OT�<���_j_�wS��h���⦉p.�1}Ҩ�m�4%��Xy��o��f�]��=��Fߛ��v曪�Z*L�JE�Ox��-0l8)�](�o��M�����7���Z�����9��}��tɈg��ƥ���W�ِp��$���Oæзw�;�DXoU�*��ϊ�>~�H{����[%�7��л|v�w����3=Jխr^3�M����-b5��-�T�X���8p>";x=�k�5��tWa�e>}�K^��rK�7�e�&w-+�`��ӧR����&*�^�"��2Ub�ִe��Qm�x��6����iO�-��]�o�,=C=%�Օ<�2(ȁ��b8�{>^��yZ�L��'1��Qs5[�X
�*��r�p�p=bg�����Rܲ�N��ݖ�2�x�.L�z��-־�NYD���tŝV�k���K�����Ú���"GR�.#����R}��F�
�<��z1Vwb�x?����n���]��O��+���:��'=�q_�<]gm����k>�,�ws�>u,x�t����;>�Z,���~�v��; ��}>�v�*E�8�Q-iE}����|�_4<�Cۍ+��/�]�x*����YҰ�3�)r6
��ʪ�0]Qu��X�Ȧ����>�7�}�Ƭ_m��k��Y���d+�%ۊ�`wk��H𲸸��f_���uA�Uط���S���a�R3�a�ݎ����7����C�5"#�@�ɥ��˩���314��4�*�wo���w��E�+׾OjLdNugǧ�g��o����A
Գ�\�o���,�sok��[K���;HG�='!��N�E-i�Cz�\�vU�,�$������跩��|{���2��iǕr��·���#`9Y~2��p*>|`��]tN'VS�2���0WB�C��>���~�f,��0RV�B*�s1��}V/���j��>��-`�6��	֍�M@T
�����I����h���,�}���E�@�Y�h��
��	7ݨحuui���:n���V�K�C��6���;̯nI��'�V�u�r�;׆r�mW�Z"�i�2j�枱�2���{Ě�h�x��L̈_�>T�m����[^���W^δ��
�z�g^�m�Jf�a[�������8�=]���������Q����w|�K�r'5м�LpNס�j���Y�w�0������ھoQ�us�V��$9��V�[�^���g�}���T��E5�5�>PmG����ˢ��kb�ٽx
�����l����~�cux�O`�v9��5e���^4/r\�,�ɶ�mt����X�U����f'R�B�g�]�}n�*�)ʓ�)��;7�N��d5e���(|���_
�ME��q_��d>Rީ[�	�ZO<��Ys��ެ��OM�²(��줰>2�\f\�j�T$�z�l����J&����b���d��͠��('�%����IjZ�]V^J���v[��"��*#Ӫ�z�ӹ)t�p_��l�]���+�����MNQ��*#�$��W��4v�y��/7J�|�{��J�Tr�W�m�=�L��ntV}�Ny�~P�/�m�6Usf�*+(T�q�1j)9�#^�.?fw ����*�q�>�|�����ɝhm'lmS�r�S�)^���Uuw�r]������^S��ׇq���¬�=/���Z���#�^�FV��i��aN&T�4ay�n(K'��3�R�g9ݸ�U��o�tS�fi'����2/z���esȬ��-q5FPt���j��0u���.���=�yƶ�2Z���I�ivźx�Z�f��&k�ͣK��[�����b�X�9��@���L�� e�$"<�*"��Z�����g"�����6W|��z>bf�dI�ܯ�)�����r�ѫ?6�!���,>�sW�8�	ƛ��U�[8�G�.ǆ�� �`c
n[��d�s�R���Ȓ�7�ߌ(i�Ē]�)�ә�h������Z����k��Νtf���;#�.���XT��(X�EE�0�1&h,gU�+=�p�\t(�.xW˞Q�nj���3���^�U��s�L��b��|wDG®�ɛ7��GxV0j�Ƅs�K���cX[����)�a.�-BP9��}��	��̆��7��|��k�&���X�3�ސ; !b+���QF3JƆc�n;sMLX�S�iX���$
I�D�v�g+o���T$A� ��g��T+�t1g�.��B,򹈑�V�$ǖ��Un#�u�M��EK.ܽ�(�Gv��:��fo
x�:�Y6����M�T�)����$�7u|�i�3l���`+t,e^�hަ؊i�j��ĵ�X.��o�����Q(�,K���Z�$yfH#Q��*�V��*�z~9H���`�
�ҫ�3�Pv�t����-��zK�Q���g��,�n�7���n�����h�����S�}���A�9��de��ǡ���6�j훷�<�eg0P�7����|��p��!�R�k��:���8����+�e����ܚ����|�9�����C��گw>�0�3Wq�f87s�jYµ�:P�칤U�Y�O	�`B�૖��up��`��:�ٰ�Z��Kl�9�v�]��98��.g�:>$d"m�-8Fn�}��5]� ۍw�	0f<�1y�J��`~N<X}<��%��8n�X����PP[�Ē������h�b�w0����.�V��y҂��a٤�K�'+^
�'oc�E�3�u�7��*�
Kr�9x9���gd�С�#��YCGzg�@�*��,�uyV�h+1Gڶ��Q��B���}]�7�&�;/�ԲE�n��P4WCsV���y�� r�rהʵ���N �.���@��X�����+I=0^'�Js��<�
�R������daq�z�-�f��F����-��=n��xsj&��ߣ�0.f�C5�܎�Yv���j�x�v^2�����-qQ�z���Z�����.엖T1�q�T����52�hw;�eB9��&pF29v���^-M,`f%G�/��Q�Z7!<�U�`����R2}J��X���X
�[B�)P���-dD*(,�����T**�,E��**����W-��*�UQEEXŊ�** ��U��X,D�$q�"��J�cZ̲�\j
�Ȣ���
6°D�(��J�EX���+QjT[lE��TE�*�AH�b��*9nXJ��"�2�ز*���m�YD�V!��b&Z+QT[JEb1F�X���6�m
�C����1��b�Ab�EAAQQ(
��K����dQ�TU"�J%J2�"�@D"�,DdFG
�VW-EU�DY��2�.R���e��m���Oo��
;�k:�W�[�|��6v��������2K�X���W��nfu&h�Vӂ�烹��1�r����n����K�{o��:My"O��C�B��"i�����%�a��aa�y�U볢�C�USzH�w����8�i�K�I�Ծg�2��Y՘�eł^L�����]��'�en�����7��J׃�&�¡�����R/�>�Z)4�k��~>��Ƙ"9�?_�Bd��v׸S��u��9���`��Q!�_N�eO$&��2�Wx���x�HJ��}�K��ٛ�v�߸��q�i���"�>�M4#D�\t����w�y2���wJ�=�J�Ľ�_�kԴ��SU�->�J���{#��'�����׀W�
�����M������7��_�K��U��O��	_;Y�=0e�����7��y��Y�wx���ޔņ4`��k_�^�^J���d�^�V�q`�3���^�n��]�-[�\�8�����Z'��ۣb�/��k�V=�\�9���5"8���O��XF/x�h�s��Vi�9��	���BEڽ�Ics��X��SWK֦S�+��Ig��+���(�m,�Zî�ϟ��)����Ⱦ9���p����g)S<�.y��t���Ak�yk
듳i��I���M�л�=_4{k�Om:��%�J6���S$�a
J�"��.�l�;z���q�ղ����������'៾�v�<؃�3lW�G��M����S�@�~���kܡ���Yk�:Pg����\'O,g���G�gL���U�Y������n�&<�4Á9��lf��=h��u�y9�9�k�����ǬY�%�H�j�˱���|���Ʌ���Q�2��R����	��*�������>��&��\��śA1|�}��0�.��n�aL�4_w#���7�����㜮�=��L��%p��H�9K�I���L��_��{�K����EO�����{�����m��y_��19�SK��RÝ#��r���K�W��T�D�\�����o3~��:}�	yp�.�脥�{������ZHV�\�Ӯ2�:
�t���:��M��^�i�V����ݔ�bV^*�%����v$D>�V9o�M��{���Q��v��K��fD��"�_�"��\Ff��J�{�+9�7󂞥҉��Qtm��K�����H�=�"�U�u��	flL�ْ�/>��3�XԱ�*�ِ�N��ML�o��)�wz�ج�%`��(�B�wP�m�7:�7��\�v���߷p{N���K�8��u'8��Z�O����_n�m��=p�^�&�af\�V�繎���}�uZA
__\�v��]��ǲ��=7�B�(��f�\�޿�}O���=G��+�!�c�d���jߡ^�\\����m�(5�!�-�w����=�|�����Ɨ��Z�|g���p��V���k��O�>����ˋR^�Ev���~�v��Fn_�g�]���ی��d��%w,��ӃV�qgԴ���#�fmwE�.�X�/a�=r�k�հ���]�M�fg��a�}���=%M�c%z�â��N��U���G��h�`��{�@�!��Q�`ϻM2�V�e���RǎMv�v����;��#U�+nUe{ ����wxC<�c;��"��(u�����Ҋ,��a����jW4ĪZ���Ҟl�ǋpo��>�d�\��q�eUq��:뭲�42)��(ŷ���Z�/�������%vZ)�]���\���"xY\\X(&e�we�wa�Ә����T8op�|tҮ���� ���7�1�kּ"�䈛.�<ZZ�S/ �L{�+�9�-ʝѻ����%��߅i���~]��3�s�:|'�g�NЖ�J��kR��`�A������]|���
//ws��K���*�~�\��ft�:�<�]h�'b�|��b�b*�n���r�!~�ϐ�b�lE�����-�4T��?�fP�P��������:kj�E��4��Ӟ��i.׻�#��RΨ�O���j��`ۢ�q=�n�� gQ�}��)�������~t�҇�	Y�{�Sa�#�\�w%���}�C��l��-�<P7�����x�	�U�}x�0���D:�Y~2�����՗��ͻ,^���dA~���m�B�¶��y�����Y�z`��9P��S(T��^<�c����h0v���N��w�a�V�*
������c���g���&���שz{wqƮՓ�{8!hlB
S�Ä��ΜW}N;,���a^ڲ�"B8q��<�̹M��|�����uo�V��$[���{�o,�c��Ä��;�X߰>��Z�=��Ru��b�v�kٽx`����u�{+4���
����w�d]�k����2Dem׸��z�<���]�Lr/m��KXY����p���z�wr��\M9��[~:�zkM��j�g�[jeT:���P�/���&�u󋃹��̹a5GE���9��)����6�xVJ�����=>��>1%�ҟ�	�/ �#����#2�;e�����E����bU���$�����t/l#p���N��x�p�H��p�'"T1�ȩ_]m`�ݸI�>��	l��N�ߣ����ڃT��"d{\vc�v���z�ײGLժ�(�{�c�]p�X&�ĺ��1�
�����ܹ&z[�4q��}��q5,�P��])*@�s��LtEh��������y/ܼ�^:�@/�w��`��e��w�g҆�Á��<TDi��KA��(�N��m�ޙ]�|r]m�q۹��Jۄ{�e�/&�Ef�;�l.���j�}"�?a#��ئ�Uns5���#�ĵ��5�u&t;w5zVܬ�:��N�ڦ=ܹ���W��b��Y����J���'D�0�D�H���E��mX��9��q�Z��T�z��e��fv�[ǶJōfA����x.�4�җ%uL����Ca��m�i�u���w�؏G\��A���v8z�x�)Z��,NS�~�I*�H�%[T�Z�襂��Y�"Ζ����yx�ꤧ�E�e�>r�ܣ䧒}d�X�̡}{O#�7�{��*O>�9�
2�̮<|]���O��M	Ȟ�q%�G yV&w�yv8C8WI���M��J��+PVP�um�.,��)�t��]�Q{�&.�O�4�^��~�ݔ���h��*��w7<��Ū^�6#����w��O�>�i�+���q����Hdr�5r9>��'L���9D*uT�v�l*v6�4%��5_։]�3��r���:m�9u�;���37�>��*�z�m[f�z��ʵJ&~)+[P�&g�i��k�֬du&P|}S��@L�	M���Z&�����bƍ�zb}jL�n��Z՘Ǧb`���ܕ������A���m{�Ԫ\-)zd3p�26�D�iX�wr�}z6͊���6Z�ly�\�9��x�e'����-�t�&-~�p�������oW�.��K���+iՊ^��+uh�bG��՟k}3}[@�b��f��O��N�<]G�=8׹Ce��*�Ms���ޓ�����m
�s�Um+���'%�[�p�|��9}) vg�}zVF�nW\k�i�;r	�HفJ`�\GZDtU*��[Ɩ�fo�a0�Nx(����P�I��{�k��'om�X$���﹄�������D��"m���y�7.ۼZS�Խ�b�y�#�=E箎g�����r] i�\���cYA2/��C��-�U�6'��o�Pn���9i}�7��p���YϦTł_����@��ȍ%�^�S~�=�m7����r�BL6'��X�%��"�`�z�ɐsK��f��#mxG�;���X�z�ҷ���ے�	˓q�.��BN"��ŭ�j������P�w
H�͓�v�N��S[C���ݔVW'��t�Z�4�|-~���N�U�&����{lq�ĵ�a�R����l��	kAɕ��yi!CY�K��9�o���/QO'kd��\����59�{+u�1�Xay�m�O��!���iY��,�(��^�V��R�.��8�~�;s�疊�����i��O�2����U����n9�3ń4?��k^!����f���'��*鐊��H	]=[Yp���>�nc�ّei��y�c*�c� �9��qz`U�z�7�c�6�aǹ�k�~�M̓6;j�P[��'�>}o��B�L���k
�C�7��W⎳�l����G#��rg�~�z#�Xg9vF�ی��%��	�84�+���b�r�[Mu��ϧ�y:�u�Aw�+�*�����f`w3����GOv��P�
�G^f����g�f������jE�'C�Ѐ��*��i����/�w9C�RǎMv�sՎH�O�5���<���G��q{U��
T8��(q�Z��Q`��a����o΁�ӊ�7�
��cP��j"}��A�G/4.�5�wP[$8�˛|)
�e�X�'v޳��=n۟-ےp�\�5��m�;�zD��zz��8]�@�1VR�	Y����GXy��s�p��׽�<�}�er/,W���LÊ,X������g}�'z߶��~��*��^۾-X\�t���E�
��3�#�
�l�,�SVW��SM6�w{w#�g�}��(�0�,Ǧ����v�Zt�qqe̱���Y��@�rY#=�vq��֔54W�z��q�{��~�q�Z�:SR"A.�5 ���ξ�pz��v�OHk��OzCyᮒ,��ԡ��-������]������3�{��`3��!3�����]S~��bS�[ːL���,?;\�7,k𕙧�R֞��jT>�!2A�/��L�򶨝0�$-�ZU�Q��a�i�o��Y���E�qǒ�z�W�g������5]F��CҼ 	�v��vY��H�őخ�;.��5GV���o���l�E[O����/�� o3A�%�9D��˸p?R���@�p�nS��rc��ܢ���MĪ����T���.�>��]���� �:�8K���(g�����=��#,g��|/xg͕6n�u�Hџ^����b��cl:�oz�И�����E���f�u�͟
��`���|q��Z�Up��͊n�q�Y��-��~����R�i��E�G2��@��K�J�n�KA?a��@�"�V�$tqVz\
����T����|�ǒ��2�+�Y&��X<N�yK���^��+��x�v�ȵi�k�4N�DO|����x��pz��ǧ����{#��ln�}i�b=Ӯm��� Ǜ�y���N�[�J^u��\)=l#b���3)����7Ч���wQr���s��������wtՙ��mL�K C��P`�z�Qc��A{&t�uYb�@��_���fuKxo��۪���Y)@�n"�D�>1Uq�rɫ�P��)h���y,n3�K�-G�T�e��'P�Է�Ӎjπ��]>J���8Nq�-LtEh�~�GW.��PzM�O����R�=�����҉�1��P�X^�5wO>TG�N
����1@��3}��(�z�L.
Uǳ뮴�|�\���6Y2�ɹ�Y���<o�j��]�ݹ�J��;�������8	>]�(t�<�^�.���S�le���O�˙I�LS==���s�]c>��$鿦'�D���/�A�ﳍk9n��u;�:��;c��^�jK����n�7���9.zxA<�?	^��_o��_�p�E�����[f��3��/U���{��l��u��O��9�ٔW���m��,���3D>V��^o�K��t��Aʇ�w�\Q[�
������^�	x�̹�gC��ɺ+e	o�؋���9+�y9��s�����^!�3�������2�w����wcNIJ׆,NY<*�I*t�_�T�"�g���Oq��>��o��tlŇ��J�qB�˶+Ӯ�1HN�e}<��։2��̶%�ٹ��BL��������ׂe�Z/Nŝ��V�a5n�h�
d������Op�:�0��s �C��"�Z�`[���j���Nߏ1�ՔPȸQ��<G�z��9k��Δ���7e�;lX�vg=�hpJ!�᎚O�������Y��>Ռ���;K��z���-qFl��ӻ���KÝ�@�m��4�8<\������\0�<�N�=Aa� ȝz�{5��W2�}�zZ���s��zJ�V��M[Z�t:f�?���e.X���8զTb�>ۍ�\�h_��e�`ۦfr�?5-���H�W�K���YE5t�j]ۧ���]{zM��|U�>�+�G��,�ju����hzq�r�f}Yk��˗G2-X��`�Ի��kP�J[t�oe����4�=5��L��Ƙs��c屚֨|"ܫ���J�ZJ���]�n�]�9N�_R�V��,C:���h�|j^�m��PI����z� ���0��Tey���f�)�ib��k��X���\%����N6k�N�w�������;����I\�<'���U33�T�Š��]V�#n�%4/6�#�o���dR�2j��x�H�%LئwL��ʗ��]�\/,.]�І.�]�2;j��V����K���'/7����o�I��fQ���Ѷ��ۑ�9���B�b�VǷ��K�E_a;6�Iއ��ɒ(��{��	L:{O\�˭��c@S�e�즑��P�5�0,��>��e�B �XȨN�)Xzq��j��0���r�i@���՛��9� ��J�����n�D�%�}k�X���0���2fӉؾ�͕��X�ċjk�`ƃ���V+v�jTf�� ��I,�V�~�����p��Dn��B#�"�r��Fw-Ita�E\�9�t�{��D=|&��٭����z{,��A�'6��T��<�7u���$1���LJ�>��<:��[͖ɽR��|Vyr�;��구������5,��ׁm�����q�����nS���m���n�=K�C�\��gB�9Xj���WrV�6�t4�6k[}�r���u�X�t�!�唀W+5-�p�m��V�"��|�WRof��Ym ko��Gf�!f���\,fڔr�w �u��;������;��au�#
���ωR��;�P^Q}��#�f�]b�{����%h�3��Qd��#j��&����u��-�b�b8�=M��!V�H�ʙ����5
z�<�y�.�(�͇�^�����f�1[�;��cX4���޵�v�����NZ�dun�k[������G�uȞ�{��׻�f��U�f,�~l�2��^V��{�Vjԯn�������DBBⱽ�����d����1��Zv�:T"�B۰b�wL8p[���t=Y01K��ù{5�y-��ٷ�uθ�LL���Z���c�zl���sx�v5�ʇw5��-���՗�gT���ap՟��"�C�K�Z6G7���1�Ԝ5Ӡ*v�k(�2�f[2�c21(S}a��^m��̖:�M�r�*�eQ=	=���G��e�U	Y�Hjn!!�^3G�k�ǸI��w��Vm���`�e0��Y]��B1A��:�Vm����A��v�!}�7cc��vm�^�ҹ��Ԁ�*���Ÿ3��`,�6����9��n�N�m��p<�-+����ޞ1
�LQ����U^�ۄeLtT��V�U��wŷvR�@9b��L�GT̃q��B�dt�M�F��)��5f�ۣݝ�U�l�c��E�y�t���c��I���ެ���/������71�/����=c��{8�	�$H��lTb�E��[h*ņ0�TE��1Aci*Ab2,��L�
�E��¹h,F�X�j�Am�1�b�E��$Q�UcQA���)�QA�\��VEUX1U�EX����8���Yk"ŋTQ-�cRL��TU����V�UIZ�HնF-B��\�(c.6*�q�1EDm�Db+V��"ũJ�UX���[f%\�R��b$Fң��b�j�-k�b�
1�kU����@b�EAh"��Z˔��#��2��b*��*$H��F�UTJ�������r��K)h����Z�
�"�e(֪*�)kpb�5��+�Ub�����~���Ѽ�NC�ֶlNgo83x9�����V�S�lŻ�,�tdz�h��X�6�F�ڴp��a��޹��2�?6[7H��v���C\���G5`\����|���Ʌ���
(�[��a=�L��3����z�l*x��P�DӔ�+�6�Y������f��[�VV�ù\]��'��嚽j�d]Aob�<��Hr�$�1��TxRzvy�;b�x���<�՛�sG��}*���}S/NR,��=S��L��%�Xy���y�y/S�]��}3��)��^g��Ǳ�-��pev�y|���>i�˅�T��%�ʄ_�	`td�^mx˽�*e�,�R�F�U7���\%n!�L�dzyA������)�OQ�Bˬh�̬��U9��2��>�@k���_��N4�U���<pSڬޔ�����'���ך�M$�VP�ա�y9�x��;+4x��q{F,���P5u��>
�d"��'��յ�}*Gc�Ɏ��q��Ⴀ����0��-���AεoҊ�2�S7�ws��ͷ��Z�1�>W*�h:׈�N���{1��zV��	���׆�Z�k��[Mr���`Y2��+ Q�0�1˱Ƨ&�}�g3k�=e��7F���;NK�V��\W�K���>,�pl۫�#����ei�W=���7]]������hI�sp"���u����Q�����*.=���0�u�<C�gHBA����aw2�N	��%�uk�p�P�.����Pɲgrђ��Ou��5jW0Iy^����=��nji�xGE�yW�{��VX8}�ĳr٘�f�A����A�����;�WwsF·&�_�8fCW�-�-:�P`�Z%�s��-gե��(x:�<qF)��v�>�M�̧��Y����z3�GGB��R��C����������Y����,zf�Kҥ_����sS0T�МP�M���a\X]K���EUq�uDqے��ec�w��aH���2W���{�Z�������M�"��V;>wk���W
	�4���zQ�d���r�x��G��ݗ�FՅ3|�)}Zb �\�DK�h�Z��n�D�z���:"�OO�V�y\������Wܭ���ޜ%o(0_޿I�_�ϡ�&#]OmTI�:�э����IːP�eD����rܱ�+�KZdPޣ��tLۼ���^�Gؽ�줪�UA�.�=�W�BiA�\�f���tGw���t&-�6e;��h^ژ
��cWz-�t�N��I|���g`�(r<[fJ��[n�F�����k�:�����]f)���o����+x.{�Q��/3��%�1e�n�����7J��#f�sÒw��.�Z&��om��I/ѵhM���g�����׾S�U�0�̶<%u�B+ah��5�;pu�1������iK��+_�SgU���ZE_��8�֌Y:ne�9��/)>�@T
�p�n|��P;�Y���pշ�;7�����sz]%a�*Ö ��n%��Ε�K���g��{iy3���"O��Μ��ႚ�m��ڱ�φn�4y3�L&�=�I󞷥xGy���C�Ns1�j��v)����:}^�zd�δ8_4c>�y��W=v=+�6|s��9�7V&���%�*]a7��'[xw1��tՙ�])CU�du�`��6(2�ٙN�/�H'��x��s�6mzd�^�}��V��4���S*�ԯ �|`��I���c|U��yܜ�7�2�d>ӷ��ȡݿ��xVE����=),����G� L����IR����pݞ�&UW��FVzQ�̝B`j[���%��P<��-k+��~@��zN_��6�I��sNW����Č�ő&9����ÏMN]0�|��$Z~���(���������:��H��*n�o�VZ'�f��k��-�{"���uC��me{�x��n,�]�l�+���ΥtZ�B"����0���J )*��؅�����E��
�6w�_�uvGU�-�,vc��b}��ۮ�5o�}B`���V�.��p;�5zV�#��dˣ�g��>�U��z�F�5�]M��=c"ϋ���@�#A��S(P�c/�3���Qz�󊆑��Y�u3�Ë�^���ѽ�s:��D�`���7w���VWxo�^Wmb�3��R(RK�Ǻ�W:��Ca���1n{����R>�K��*�J��d6^���MFuGsc5��,�����KɁ�˱�>�����<*i%�)��)j~������ړ���:j+3˰=���K��%S�H�Xr���	��L��Y]͘y�of;﨣�.S��S��zr��ۼ�7��hF��2M��f�y�K�2��&���I�M��k�H��N�{>���T��1�f��?P#��ȷg� ���*.pHq�N�u�V׮9]B�g$��^m�g��t2#��';�G���l��t��r�I�I�}�T��m;�-߭�+q�/���>�[��'�o.�7PP��A�E���&S0���s�'|�v^����/@ �x�wXzjd_1q��wg������)�[��iM�g�\��&o@�T[�.K���=�"�����;�5����.��V����6�A���N5}��cd������rk�=��W��k*L���i9�p�-��ǽ��5��-tJǡ�.Xv/O9Nh���_n��+&�'�c���;I����~Kz��v������X��S]u�Y0��_�iő���������{K�HǦ�K��,:��x��hN+5tXY��h��J�?J&�I�;m�Em�"R�CeT��i�oMC7�0�y,i�s��S��˯#�{��>Y�B��V5���dl�����[A�:+�Ċ�/�c�����3=�&�3<��ynS}��7�-�����s���|:?]J�,�.%���0�qvR���Z�yy��H��W�Vt�-��t�]����\*)��[�Y~�4h*�#���t>�����":�4��;�Z��ީ�P������R,�1KB�L��Vh���Y�$l�n�9b?b˲z>��k�\�e�g�ܾKZ��C�d��X�L�Jփ�eB%�&�31��j+wpZ��^�}�?BH�U�*Q�%Ǭz�Pg>��X7]�0J��e[D�w�v�r�
~�t0�/Z�q����1�m�ѝ~�ϯ�!��7Bp4�ǵ��˖� �᭡���t���F�8������ۮl��+�htRɳb֪
�y+��\�<����Bd�v@���,YJ�d��q��'��W�� ��au���A����$V�Y U����h�N8�
UQۜn�ˈ�y���Vk���m9칗�=��n�w�n��Y;aY��h=Feu&q	���>��鐊�ݧW�ٯ�;�.-�~�����X�2�E�ά�<G�&? �;Hf��Ex^W�X{	�����ً��>��6�åi�YI��ǀ^�U�z��Yk
�>+s�ж.��@<k3u��&c�^�oM��q�iq�~3�#p=��6x�7��>�)������i�ȫ}1y�X�(E�\G�}w"��*�����l�w3�t����u2�O�N�y-H��ѐ����� �R��V��R�Bӡ���.��L����,;��o`��j�n�M���o/�W5���6��^�Y<W��mL�qLP��D�=�R��:�k=�+��zg��N��	R���8����y��::����$��4�j�L�,��;zS�o�ɠ��U���~��u=���N��E>�]l�Ζy���c�T��y��v�h\��>�\��w.62��y|�V�>Т'��@|�$0fL#"������p�%�z;�f��=���E�Y�wn}�t�#��nf�bܼ�0��gC�:1o)�-�cJofN�V��]o��P �I��o|V�����k�l�Fթ��~
.��p�E�49V��-��=zr#���W�����b��
�/)�,?[#N�ط��!�g:ç�zfq�d����m5o��S��̠AoԬR�v
�b�C���!������=����S�϶ff��\�l��^#���%�$������iWiϯ���C��҈/���śƵd=���V�4:|z�{�Y�a���˳?F�#�"�˪,��ufb�]�}M]a�>�%N��s�`�Zс�'M�2����΢F�o����z�(;�놎����B%KVpKi��P�S��^��}���Y�{��{�o5��:Q����;��O�P�ʳƯ��Cᛷ�C{,��nE��zW����m�3+�����l������SǴ!,��0O��R��-�^�Y����L�� {#;4:"�=��ٚY�O����v[;5��b�9h���l�6(0^�3���o��zMd�6��i_mh�*y)N�ef\�:3F<��a�4�5��OT�G�]�3��9�e�̵ܽ;"�%�n�K�.�m��;ҋr��E�+3��F�f�&7o`U�5�J��nVG�q,]�'/Y�N�:�u�r�V]���a��N�nL�q��p����ð��s�^V.�W�,�c��c>�C�dW*������[���LV�b��X�3!�T���;�ɂ�J��Y�I`|bKG�Ef���<�36ky��D�b�&�~�[+���d�Rޯ	Ƈ�`3��TԵ����q�2r=�^fH�=�E3����D�8ОX�/�
�(o,8�S�t��1��I�������g|E�Ը	w.�U��v��r樽P��L����d�7�R��q<�o[g}�;�f���v�#A'��b��^ٕ�Ea}x��g�hm�[慡��%��ӯy/=�l��~%��+	0��D��H���B���,庌\=;*yx6��[�˦�x��d�y�O(^�TŹ�d8s�/Âx�5�GIt�
�~ႭdW����X����~�c��Y�h3"�y0?v4䔭xc�')�C�)%_t�_���׎�g�Z	e���ݧu���v������ۀ��z]%e��.�8�G���+yv�+Ӷ��������y�h7��_4N5�&M�j�8h��{=��ѽu����Zf if�հ�ʎIw�g�5��8֯q�K�]G���#���2�wTܭ���ὝV�pL��8[���*[;U[K���?(|5�<JS�0�s�R�t�jQy�p:��'�۴>zIaиN��x*e�\/NC7|�V��B4K�q%`��1/��x�l�}�9�ߨ��g�!PԬh
ԫۑ�-���Sz�ү]�Q����u�+1����sD�.�﫽��ۯ	�ط]5^�~�nx��cu�Y�`���ߪ}V�-���TDDl�L������V�r��~j��i�s:�G��F?��{=���L�T��.O���/j
�,�`��q4�O;��h��Ǽ�G���SK��Mv�Ц:���s+���3l�atGC��	;I����~j[���v�d�7>���b�*v�u�Bj�2}D/();[���X�`��8�ԉ`��E���xQ�N5�Oc��2bח���UN�x|z
�\��hq�:�E������K~zj��f,d���̭P��i�3}��}{�u�@٭kOZ/%�,�+���q�46��T�'Ռ����~���o�3�<����y�{~I�[�qb�3��~�,�D�R�l�0�!Ƿ�0Wy@Q��)'��Hv�9+;!�����H]�/^���H�r1�ݭk���ОkRk{hF��>��fVO^T�F��˘����y&OwPTb��^?g>�c�i��C��qR'���Ƀh�q�4fU��3z.�p�s�S��;�Om�BZ�	[�$]�ډ�8�!�A[�i��=�tp��g�y\8%�Ĺ/U3��~�'s��E~��Ϋ��~zhsA�V���ܽ�<�9�)j���192�)X(=��0�[��neݱEg���x���]໇��P&V��[0��WL�2���-h8&T!��e^̸����2��?H�4��-%�x��ϛ��ja���;+u�1�+/�m^㊯z�m�Z<ϲF�k�gP�bD2�'p��>X�|)Gnq��-'ٽ)Z��]�|R�e(�R<}|6�}���Y�S�cń8h�^!�Dpvo틃�<�c��.)���rlv5,��{-��x��x���p�8Fc�����jT}S<~�Ҋ��-�̥���w��6��s�"��,n=���Jִ���8L~쵈�_>LxiKs���dZ�^3�UoW�V�d����8)��">��9vF�{q�2l�ܷ�ܶv��5M��T^y昗�2��x��
ZE�P�*��gE�3�ĘܶfE��f���Ͼi�[{j��I!�%D��{��bod4lzCז@�o�n�Փ4���>��A�o�3t��$�Yӎ,�2s��GV���f�*7� �̱��Pe�����|�Ck\�V�G:�1{dL�v�V��)t�n�=�븱v�cb�)z���ʌ��Wu2�p�0ی�2T8�����X�'�*ݽ$�(WDfCV9�����6�屔��K����U��ԖoZ�p9�t�W\��Ϝv!��(�3Z8���r>�u�w�e�kܬ�p5�ů/gPn���En�&;�*�N�Y���K�ㆌ�=J���w���su��z��̍�c�z+��Q�Z��k���	�Le�Â��aY��2�N|q0�e�eIq�7`�Y�|�D����@�Y��-�'�������N�l+�ԐQ��=�NVF|v��,�rJy[��W`Ș����N��y�}�~�9M��<N-��J&X���e�j�֣�8<�ϱ���6�s��J�TbI��G�[��=%_eZ�83^z�\HXq��]�/A��6����/
ǌ����]h��VA�3P'.��U��-�T�]�Rַ��ّ�-L� ����PZI�xR�����٠������uYʜS�V�5θcM�y������`�����c/fp�܂�X������)o
v�ul��Q�ΏY���t���5h���=�
 ��Mw�M�iw�^>�';w��N�X��E�����/�ԫ�y$�do5��*zh�jݍy�
�e���.�Z�Ժ�d�6��nl}F����m�2v�	�lt�P�����J����2=������'���xt9�]=�y�l�\�՗�Cͧ-��la��k[ַ*�9���fi�NV9p���wj�k�U�=U�t���=|�#s0�zՉ��T�U�/3y0WN�o�]�@*
'�]P Y��(ǍPչ4.*���d��4�k|��  ʵ�w�V�6��I���a�h�q�z2x��:3�
�:�=�Ȗά�Es����
�r�5EN4�ƶi�_ft�/���U��M�iN<���/�vv@<M�#)�`Yr���m�R��<�km�+���уv�Vcoxpbt��E��wm
ІbAQ�%���|�������y��a�8�x)XN��U�z�v*;�]�B6��iz��*rN]6_V�Y�|����,8�|1�E��@��w���&�W�D �������_d�4��er�W���
is��v J���5�$lFĬK"�-�s{8���5���C\��SsE�+��k�����1�BZ�)�ua#n��é�"��u�7�,aK'2�S�|�?,����2x��z�WTi"ps�y�[�C����\��i�J�0[�;�M:��_`B����w'����ٓtS�|�7kJ��ze���9YNp��sn��7��p��kݟ(�cK(��TGiP���HV娫1m��(�b�TVV,Q,3Q�L���1�1�*�T`��"bQ�b ��ʂ�\lTQQ�1\j���EDKe��b ��QX������b,*�.�UD�Գ�fYTb**����"���"�("#QDn%*�V"��EL�m�""��l��j4J�b�1P���3,�Ȫ��j�-���UQE�QB�Ub,EUR�D�Z1b*(+P�R�D�E�TJ�Qh�
ذ+Tb��U��2��F8���*�UG)DX�DV#-�aEX�DTE�X�+2�\m�QTDb�"���@�ګmPR�R����,Eb*cATUH�X��*�E���h��dK�Ħ5ڨ��,H�*�1-���a�K��+Z�h"�L�eTKs+��f%�(�e*���/�=V�Y�R�][1��]��p�
n7��w�΃�txV{g��{�"G{�P�����p˵��8�u�`5������/?|fu�Yh�9���R�@�9z�*�.���kifU���fK[),�}G�N��/�LΩc�>����;!唋:���қJ�t���5���!��Y����ӽK�-^X��&�r� u/��鹜x��mu.D2-U�;7�T�$rQysz/z�#eu�+g"����1d}t{������X}��c�\�H�2�oON=��r�o2{N�V�jU<"B2<��e��6��3|�?�B�c����f�w{�|2�Ц)�7[���`�.ӦZ	��)�-��X'+}gqw�=���u=�43��������z3��]'� w`J̭K ��vP�z�TJ����07,k𕙧�T�ѵj~M�_��խ�����y.\;�^a,��	#ZZV
3���ҾyW)k�����z����؀�B�-���y��~煊������HjΌ
v�˳�,��t��u��֯'�W���a�G����I�b�ޘ)'"�9���(��>Y:ne�'���tl����J��x��x<��-}��i#�4z�fg`<�?uu��'��5L|�L#0v��S>�����J^d�dJ������vu�����]�ԯ�9���P{J���5m]�4��XR���M�F��J����L�2��JN��u��^�~Zv�;ҩ'�P���qc^KDt�^��0YnJyL��'�k���j�Uh�N�*�P�k���z�ǟ���j�{p�-�[ҰJ�Dʞ�Q���!yS�y&{���cE�^�>�u���1�x��pz�������o�>CJ)U]ǧ�^������󕧳��`ӺU�UtY���YA�\*�:G��|�!g�x�B����>���^����&^���\�;��i�7�i���3藆�z�=�����Q���L�=I��T!�a�̇�Rޯ dP�{&F�a�=�R{U��'�����b���n{w�k�z�0b���H�V4b�:��Է��q��F�ǲ��U�H�5�{s*g�+���ҽS�g�R�/.]��w"G'�=(��v
���S�w����sv,U{`m�,zDx��h$�'qy�Ӵ�|�\��+n�l�e����t�(Vzt�N�M���ݏ�^��g�_ӽt{�P,��j �>}i���^V�:�nx娆�<2�lU��\���vn<\�V����2a�|�,x��P�H��9�j��k�<��4��~�# �C7��(�������w�����x�:��wY�.�yk���]�' ��J���d�=��Y�{1QO�ݏj����\�d�-6=�|��,t�I�#��?Yw���'� �s\�h8��(8�8�k�������gyu���t�5�t/V|�L[�.< �����H��)rH�eV>=��|B���4����R����άϖ�\Y/&%P��)Z��,NX'�Cs)$�.�>�jcK�9ο@��b��tȫ�������<��:I<W�H�6�,=cI�E}�]�]����D��<X����$%Y�]3��Lŝ��V�a5aЍ��m���MT�y��`�I��_�*��5���h�e\���9{�C�aC�������jm��>�{����-���*�b�n�F������а�C��k�����"\/���W���{�5�#������r�_-�ǚ� Zo��[K>�z�u�r�����Ǖf&	�3��zK���lk���8_����k^B�[aşS���	�ұ<�����
�Z�3;��/%{���vZ>�#�P
�ҬgY7�H��i��R�'����C�aq�p����T�%?%:��5thx�q�#tz%F��S¾/y�t��ml�5u��r�
y:�m�#Lȼ�lN�U���𻝰��Z�w��c�5���F�f�zC�����.�Q�vl���*�fd�Y�3�hܔ�};����i.����wؠ��A����V��f�h��p���#l�N���)�WH�zjD�*��r}j�4*e	b�7�O7�l����ţ�{�І�����R��>���L��=5�}�	�uY7�DJ][c\�ハ��x�FW�?�z�y��E�\k�'�~H�j��v;:�4�3�c(.۪oRoXo��K62s�G.V���AL�ytY�,�4�.D0����nP�K��}�߯���Ű�f>�F*V�3uS�
�s�g;���<Ѡ����yj��a^yeZFj�7/vtF��$����BXC��:�}�����_�OT�,�ʘ�K�a����+�=���nwH7=�-�<�Ԧ]໇�z�.�/�ؼ�:�K˅�˶{�	BZ�}�׫ꏩ)�6�v�\{����gM�U��G�
ϟ^@��q������A���[���V]�ee>�ճ7��T]���Q3�Wj1}�U��З»��>[x.��^��^��z���^�Ӂ�r�A�2�𲚘Up����s	޺������H���!�Mγò�4�T�\/�>������\��@�P��&�n%�X�������n�o�=�+�����3��4�W��F3���|�^0�QF���r�4�34u�Uۇ����<�l�{����n��3���!^�1�2m+�s���|�E_"����r)s�Y�t�ض�e�8���!T�b[oN�w):�Ϸ��KAb���E�ά�ӷ��,�F�Ox���Q$mI�eZ��N0�Z���CؗW,��
�6V�>����f4�zV��	����o�.�X�Y�V���D�d{�?{U�.[>��8p>"|�������zUw�����Pτ�3�q.�u�y-ڧx�N�^g���	P��PH���X�j����%���6�US��Р�{����cq	��o��(|�e����j�Gi���"�J��v�e�Y�>�)�M�������3 �,x��oW\ۇ]z�f��\fUm���q	�9{w"�`�+�H��p��f�%>��ɬ�L6��:��N4=��e�^4ͮ���q����!��-�Ϻevӓ�"X�}
��E5{e�>�<;�1��[�V;>wk��~�!ō�Y�zƳO�4�v�D�z$#"\�{�i��������ja�Y{`�B��\ѱ�t�ٗh�ɥ���S/ �L�M(�<���Nc"s�>1�=L_e��y��~��Ju̾X�����P�Z׊�S^�Sސ`��ckp��sPP��G	4=B>�'vK�\E�b�^jʰ�Y�-ѷg���49�ED�{�Z	P���0�3	{*:�;�κ��\���cǹ-��<��z��N<=�/���,`B\�A+��vB��ʉCo�� ܡ� �#�.�}��o�u���o�<c<1<\}7��ˇpK�%���$/��ү�fq��ҞU�6�p���qMþ�����uz	�����|���0��.�8�i,��Rge�ː۾K^̬��4�N��I�T��{��X���f��I[��.�:��9D��wıHj�~�^���u7��,���մΌͼ0��({z]%o��NP`��W�Խ.F���[�t����y��]�g�܀�48Ӳ����<.�c�������	�{p��-��z�#��:V��#�ǧc�l��8��(oV{jY�k���R/�׆__���k������x�Z��#��:{�Z3��7Tf�d�V6��:ҿ)y�Q�
Oi����7�&\;��Y=�g���2���5*Zÿ5Ղk�F�\�;��Mi��j�ʭ�0UC�3⻺mz�$�}7\�� �0��4�S!�n�d>��[��dP�\��V{���챁W6+���:O�0t�ע�|�y"��`V�C��j�Op��U$+�Vj�*���/���s�v�jLm�0��-�9�e��G���|Nzc�K�q��K�M�	�W�Q�(�3f�����w���������r���-g��w�E��e�ڿ
�����M_
���R-��ΌBN���S�Ƈ�g�c��:mUr����W{���Ƚ�m@�K�g���"��.�ϝ܉�	�zQ2�����^'ЋT�^�-�8.:�l�|v�A��c��Dq���h6ئ
U��Ӵ˩S�/T#<�ꞎ�7!�/י��<[G2\=�y�g�"�kW[.Ƞ�P�h%�D�uԙ;w5]7��/2v]Kb!�d�N*��ֆ�_N�ڥ�}���l�	XI���D�:D�#��q{��6
��z�C�wS�Z>m�yN�c����P�|]ՎTŹ����%z�!}�GI�-���b&�s=�3�jP�z��6:���ux�g�9y0?v4����X��
���%��_��[cD�������X�M�4�>�v����˶(��r�������Dc�}٭��:��A����~Myh����	�qp�8=�{} Ož�(�NtU9O,�sdx��X���;ȋ}�M�l�m�*�<�:���N������1�-V1��`������*�lr���L7����w炨�����C���"�v���ϣ�hz��;[��.�����wxNT�n)M���'��"ۆ������}'oe��̲#y��*V�lu:�tb�勚9쎻S�=:��v_^�da�����i	�xׅs3	�DhXi���t��^)).�nx����s��u�~�IF���i�꘠�ܱ��\M����b���r[Hi��O�^b����-s5Y�"�$�c�o��x�h�'�k]q-���s0{�8�W<��_0T���m��4�����q?%�ОZV�j�T���0���31�X���^	j�/=��]p��(vf%];͛w��ҵ�V�}J'\U���H�H�K�_Χ`��o��tW�W��<��{B}8��^���Yk����f�IإCeT��L��禡�zE{�sۮ1k���nO=\O��}a�qI��h�ֵ�t���]�ͅƸK�v"p���A���jW��+�i8�AuDL��f�]�G}3_Η+�;�h��q٢k探�g7�Y(�u{=/<��d�����q":��^uZ�է�
��ֽ��22�x;<��H,E�9��,'�8#8I9[�����E��ٵ�:�f�ڞ�8]j��LB��1� CX����
_o��]�:Uy<u�8��^��������exmc�{{ͤ�W]�~�5n`�n�>p|�[�!�ru�b�ܪnG��9g���:F9h.fU����:oF���l�m�Ձ�oyq�+���]�p;���Z�[�,ݳ�]�Y�6b�nZ��Oz�<�<��T.���P%�W%�pud>���]����K�v�ڑ��fmOs��>�E�ut���f�+��u��|߆�Sp�[�lY������Ob��Gm{�V�[�g��y�]�Z�JB�tW��Kl�G��7v�/�!};�ZΡ=�{�E?W�]/R��6�VD������'��f�7�����:G��&
O����-�gNWh���v�� �v5'�P�f0pE�ά�e/�غ���k�*0�Ig˨/Q���S�V{�^qx:��]Ly�^�ˮ���럏 �� �v�1�/��~�L��i�{�)�/��I���g�h�W������#s�B�~���	�Vf�R��ݳ]����[�>��ӧR��
ZE�dy]F�����}�ĳ��fUt�^~���]%=�:C���Xz�Is��({]���W
[hZt9 �Z%�d��7��Q�a�!���{���_�)Zar�r��K95���N�{��E��q�U��}J�J3�7���k+����SipP>�`/�3�������,�ǭ��:�NR�KzI+�={��/�<���=1��[��o4.Ѱ�WL�����G�]qݣ���bC�At����/ueG���"�{
���Ō_u!Y	:t9_<q�P�ۖ��xN[����� ��8�+iEza0�jr�r�C���<��nT�n�Ui:j���T#pu]���A�$�w 4L>���Ji
뮸��Sˆ�1d}tx����c�����<W�!b����'���� v�b�e��2��v[��������/����W5��__K�=�9��zd���b����T���%���e�L��iK~�F��o˴S��xO�4�fFw����s�y/S>36fq���a��%]jWK��=�Q(_�.C�����o���bqs��II{�K�_S7��p�}/0�p$���QB���	���K���'���k��|��k�?Qՙ��r� ��|�$4�T��Ꮍ�"+�k.�Q���e�~~���k��k��,n�_f�
J�r�nf0q�-h�哦�˸Uc�~�Ӱx>��U�VO�D�4�ؽ���y�x_�Zv�87��V�`9b
_N�s�!��^��R{7�ya��#x%e�gt�0�||�\��Nס�c7o>q񏥓P}��:n87,���C��!�]b7t��`Vυ߽�k���^�ަ�GW�}�3p2����A����v{_%�ށүl������^��V�]5m�I���<6���l[Cn8�=;"cT��Z���Z�ujP�z\�s8����B�g>�ڔ�'��{�<�6���\ė+�ÙM��y����.f�Ӝ\�ύhTE�
�#B�/mY�QJ(�9��#����3c*�닀�uw��W���O7���3$T2k��
��/��8���u�X>KMA����x빗��k�\��Ɋ/\����5 ��ٝ\zC딌�����;#:W�D�y Fo�n��ˀ录 i���7ލV�;�@|M~�O�
aͱ��8��c:wТZ0K�7xՁ7�s,ɭ�$�q�K;.��ѭ�1b��@pP�E�0h�CNR]�gh�y���j��Q��v�T� ��d}�X��ꣂ�2f�"��pY����������pVCE����{B\��aǜd|�9g��P��Q�s��ݮ�Q8�XO��/-��si��D�zy�ù��p�r�6I�Å��uڸP|!�-C�lp��/E\�(���<�xgJ��X�.��Q�Ьsj���x�� //z�D��$��\���ĥE@�ʺ�&�)�P(XK�{���e��),x�j�z4����!�w�R�2�=lV�x�%������L�Y��N]��;���8Qh�����Ω�DR)kAvv�ˌ�V���o.ĭn�/�U?5��B��������"l�S��ZzOy&m\(����]�~����(77��Ư9}e�in��D.|��.��Zɛ'[�(7E-!�m���v꽞^Iae�|s0t��֝Ƥ��(�t��9{b��b ��}��ٕ��g2����[���e�a�Ҿ�ܴj�Ч�]����I1�7�5��,^:��r��-n�:�tE��]r��,Vm���}/�����Ƈ��Ea��=NJ�����n�X+���L��yf1�i)����ț��r9Y�ҷ�g�_ _>Y�-�����+o\-_h�a�}v:	�R���n��A����o�^��	�:ɍ:�溰q7��PN��+o�k-F��;��I�cި�.��K��/��aX�э�7���V���q�	����VӾ������0A������� p��+{t�se�f����I���؍�<)=#�ӻ��[;��5�P���4y���wE�����Xos/����V&����-����;�l	8a(�A���0�</oj�E_n�5b%M8��ܼ� p�au���N�:�x�*�|�8]k���m�C1���{Hj1B�ZJE#SeK;��z��3�ZNY�P^�gt�#W�]�4�z���E[y�sD�\�w-FPm;����l#�����U����d����)뢑_xԑ�Zż�Zs��ԣ�����o7ˀb��EQ�R��*�g���cEX����E��*��(*�F1��R(��0�\�ckDEL��Ĭ�E�ն�1e�-lQ�ƪ�)`Ԩ�"�DB�ڷ�R�iVƙDB��Q"
���U��2E+Tq,�Q\��(&Z��PX�ى�Y�1�hTD\h�[X�+R�҃iQF�b�ы�QUF�Pq1�1�0ʱ(�R(�eUE1(�Ģ�-�U��mE�UUUQjT1Y��5���V�FR��V�aTb�
�%J֢+E�dL�Fc
�	�(�\�E�c5�1X�-�$�EB۔�Q`Q\h*�8¢e�����m���R���UF$q�EA�RV*̹���a�EDr�[T[K�-KlP�����*%EjTEr�a�Dm�ŎZ�m\���AdUQkr���W0�R���[F-d��cr�����9�QJ��(Ԭ�*�����i����]$՜-��t ܗ�j�ظ��ر��u'�%ݳ4f�{)8�=�E3����DY3'� ݴ��[�x5���Z����F�;9[˯�Oe,P�����F+j�㶤W�V`�:����
[�*�8d���bf���G���^:�ݝc�F�U��Y�����Gk��O4�+v�\�����V��|��^�3>�s��B�d�p��zwW���ct՗�[j�b��^sїކU����u�-+���P���j.��+w3!�)�0dP�\��
�x]�!����ގӪq{<�5K`���`��/.Y7�BObE����:�fS��8����U:��<\�,�S�EW�t��d�U|�Ky`��-�Ԫ-��3�DL�c��\O������H�rN%ɽ�{�k�0w�X:x�x��4M-�ئJ���v�Ǿ�1��G̕(E��!�<�����W��B���y�`�DP�j�|"D�%�L��w�֙��x������ζ�0�{�|�ٵ.��9-�G��Yw<�I�� x:���P���b������2b�%�1�QYDo���,��X�xW��xB�`r�-�d�p�r�������V 9҇�����ņ��l��T��.���⫺/��(�&�1��[��u �S1�.���^��8�)�?^�lSI��J6)�^WO�<��~]t�z�7�� 7�q��[�񗛷&s�	W3|h�e�wv-[=�sc�^�]ğ\�u4/«H�VD;Y���]Yˋ;	y0?v4䔭xc�'&��,��*�l���]�a�I�H�}K�E'�\5�b��mV{��i+.(^v���W�n2�Y�yX�/?w��	�#��s.�`�Y'���Yk�E���p_2�.ZpzU'�X�a���4��S<z���*j&@�&4�7�bvR���M���
ڢ򷇩���+hO[�O����q�Se�Q{���'�GH����9�-�MB�I�\/�}���zC̏j�@�d��y]�!e����率�A�'�/d �d���r���V�j�t���n�7Թ��\��%uC`c���k��m}NfJgS;����5��� �gw.n�A�|Z�IX�e.X�j�T��{|a' ۦf;�����D�ޕ,ukHo�T�6�l��T�n�R�������gǖ��u[�p=5"X��hpql�����__��u��p����z��xø+-rJ��4P�wp7�&ZG.T�w��fCj�Ũ�W5�2M��#����b�^�6�<.��m0B嗛�3ˌ֫򝼙鯆l��ዙ�R!�IǼ.��'��I#P�½wo\����2�-����̫���Ge���l�WoA�[����t2pTW��|Q8��	c�е�uՇu�A�߳�:����[��f��=h��O��%�;	�;��Ԣ�G��8�Ԗ�w�C�P���0�ld炎\��W���l�\C��]�t�b�9��޸��_�d't� �;�A���y�kON�O�\g>�\*9��[��e�t�I�nh��b�H�W<�	B�BEJ��w�P鵎���Ꞿ,�W���1�j�3��&
����l��g��C="�l�ZI��,	uk"�?��I�/�}o�����󅳩�2B�I�kr�l�{~9 �	k�ɕ������CY\���ixnU���n�Yí9�e�W�o� ��n�#q�=�մN8)�1}���U�Z/YB�ӊ�P��)���]m�
�˝L]ɤ���%�.x��y"�%&�=KK'l+4Y�Gw�~Y���]i8�;��P7ՑD篆���U�33����C���c�,S�lp��G�鱹��ɧ�
��2�Ѭ��r���<����P�傟AC��igޕ�rAO@��[���X�]��7)���@k���3#��P#gs�EVj�p���Y�n�x���Bb�����y����}喘UC�^���j�yǨ�;r���Q���N� gY����t��6Hpa��ʹ�%ݎ.4%e�<yTb� zN�Xo/��'	�RY1�wC����~����G�m:^V=.>��N�x���89vF�V��q��%�o�K³����Z2V���9��J��ZE�L�m.�{E���O�k�{I3�s���sv�M���y�}�����unJ��b5�beZ��8�@�U�(x`t=oʕ^>�]���ޙ�=�4�1gե�;��RǎMv�u͸u�������\|��8��t��U�x�~�!��u�U�,�D��(��L&jr�K懾�h{gf2��L��e_����| ����6/��/�KK���+�����L7�y=���i��:�\"�`���u���	����;Ly�/#��W�n��������ֈ�c'?i�g��A���K=U��'���s/!�=�S�"h�h��KA���h&e���c�����߸]�@��3�Z��n1Sz����fq���	a	�J����J�.k�}B��Q(l)wf�_�uqp�I���y���?msW~;u1q���s�ʻ%�d�旊�N.�*����k�J2���yh����{AY���Ɉ`OZtթ!���gc=2��u�����ޝ��E��۶����w*<�7�����A�r�-F#�q.�����b�p���"ԍ��3�q�5�g���yz�&�9ʜ���v�z=���{�,�	�Oܬ�1*���՝}�L�0�Ƒ�q�%`�H�U=��~a�A�&_]e�z���/��1f}�0RV�B)˶���nY:wH���ӴO�g�əO�g�KɴH�!�Y���fm�gO�C���+}�����8�bu0eP����,^k�s���ܻ��/)�D�P��K�����<Z|@��e.o�P�(o�'�g��9D�}p�.O[Ҽ#��*�k�L�l�O��)yև�ꆌg�z<9V
��9��X�{�떤�c�Z�<�T6|p��8=6���u����4�x\t��ȼ�
[��s��n�wl{��\~���2��^>g�a��\��:.��u���{�ج� ��<X�ަ�~��l(VJA�ýI���'R�Rޯ"�{�ƽt�K��Z�Vدu[=ޞ(��'��aa�KG����=����GpY���'P��rެ.����w�zx�j��9 y{����.TZ+�b��y�#8�1p��b�fr�OV��|�n�����ٻ��c���8MU���T>�mL	>MV=S�2���G����=gg7�Mװ����i7ܺ�=���O�K�,�ˇ����U�D�sD/1�gu7֮�'��n�!5���v��e��ju��a6���]g�cM�Һ&�W;�K3k=2�݊�z^8�6Dq%��t%�L���t�3�ܹ�W,ު�q����j����W�z	��_{���S�l��ꈡ���˲(0*P�U[;6b|�>Ӊ7��g�Y�e��z^.��:��	�T��r�S��Ed�e�N��)P��Ⱥ,��>��9�ށ
Ռ�B�[�,{����п,r�-�d�p���w���e��e��A��h�KR�P��`���{����ŝ�>���]�9%+^+��^Eó,�^���3�o��T9�/�E�V��z՟E;h�ù�J���ؠvi��L����y���uA�S����F5�L�4e}{OHJ�S��`i���L���-G���֢��ɨ�6���I�#�yW^�m�f�m,��\�\�53�S�IK=�^V7��w(/��O�J�J�Pt=�B'��{	��E*�n�%m�uҵ�/���8�S�x���ɷ��+~/P����,A���8K霡>�J��cO������"���,�Mf����#�e˄��s�x���e���fr(	REPv��f�]�kM����+M-��=����zf���^Л=� {w���{3k��U��kx��;O�����e����S��T��b�m{TxjR9�i܇���g/0ws'�3=�W�D�a.yx?�l���q/P�w3��M+���TL��O��l��O�����!�y^=����v���.X��T���D�������i�M�3=޴r5���ۨ��G���;���%(�,V
\Z6ϥ.z��*�x�+�/x���7���ٰ�}v�t��5�Z��МS�Sxø*3��
�1Z�4Ug�~��� ��0��ƥ�n��sǒxV��0�y,i�s��ߣ5�t�E��]�ͅƸ�.!�+=���Y��=�+����*��u�D��L���0�ld炍E���
g�G��K4M_����
��\�1ֱ�*m4�u �SK�?!����ּ�L�����$���צo]jW���'K�`���\�PƝȫ�A��6��C5֊��9�]j7|���\+�����hY�_SşK�b<��:G��u����z�.���[0��s����m��b	�{�s�y�٪�%����<���f�+��q��~���\&�����:u��k�8��t�C��⼦�90�<�y������jZ�{ka����V&�I�gm��-L���G���O�1���E�`^�SIdS����GL�`ȕ9������J$w�����
|����x�N�Ks:�ɀ�[\���j-�������a׳�}S�h����U�N8)�8%v��DCo	�,}»��>[e�����X�2{�K^�fvk�葼�R��ܑY�e��৩`,���pi�L��|�p��e���S���y�%�{O�鐊5N{i�j�z�����炾�{��e���;!�I���-X=�*|�7Ҋ�xe���Lw�m�(5��C��|��k'1Y�οJр���pEp@{���y�t�<��iZ�c��������������x��]q�Q�x����<��vF��2�����+yd�^��V�q#�W�dyP��^p�,4�����O]Gi�bP˅乘wå��g���W=���to�|,�!,i�Q��xάɒ,v"}LK�8�L����n�r�Υ��>�b:��}qb�}z%�51�t����<��(�b��E��C�.j$�(��L&NP��ԾhxN4=�'{̳e�:Πh��0�UΝ��0�������TGX��Y�g"��6!��b��>�m?o�)�؛g��&���R�����i�-��/ٕ��#��B5�hk7�k=���6)N�sɃ���og���:m8�i^HV]�Ø�m���2�iy��(eD�	q�Ķ��o����nmѐ*�2S72������We��+�x[1ǧS��G�n��n^��+ڗ^��ڇ�D�+��>����;��݇�3�^�6�D8�-�'k��nK�#~�佬��B�|DEv١�H�����;r�P�e�4���l�+�U�^RnN�N��T+޾�佘�$�l�u�O����-��1	r�.��+��5�&zײ�ǲ�t���#��K�K\��~�Vf��.�.>Cz����^a,��HZ�i^���m�[��2ur�]������z���;�o�+"�]�^�՝}.��U7wi�@���\y�[xR0�=�=�[j�=��/ú�Y�z`��P�r�nQkG��]�/J�ާ3/{D`X�蕖����
�|=��.\9{V^���sz]%o��F��<����]]�����O;�f�[ ���N亼#��{n��L�J�������]7ݱ���P_rmg��rfк�âv�D�c�;O "�*�
ߠ(_
v��x�0��U��:ө��{�y<�x`��3�u�{#�y�6��wTPӶX;�f/��^^�<} �P.2�-�l�G%a�<ష���^c��3t�8�ۙ�ΞT�Z�q)��ٞ.x-;�{/�+�n��gA�+����ǣu��v%�+�yIB>F��P��&n7W1�������7�;�nQh]���S��������x��D��>�Ȯ��m�����v���-����5�3��f'R�j��p������^�kN?w�ގ�V���<Y�;>R�`�gR��P�0|z�Q&C����}�-���E��j���%^M��V+}J�"�ʭ7}U\f�M|*{���:1	:�|3���=�z�Tѕ��1Cܰ�t
�y�kK�qyr���ȑϧ���'�����.9�����}>�7�Y(Nu��8��Ϻx�x��5�M-��"��.��v���^ǜ�k]#hl)���T#�ǲ�*��~ڣ�g������bw��:�̏O5<7u�7�\��0�ww5���5h��s��>���U�"Ü��7%LV��l�J�L7��D�uvk~𡶮��N�a�$���$W�hKY�u`�v=��;�C�]�qK^�ɐ��t�zeм���{�z�*x=��D,�t���j,WU<sY����}�ƹ_�i���`5�ql��F���;�M`��I�P��Iw��-�%�Yb�}*����I��L�0FLC���F�;0r�������MZ_��s�U�ˍ��mZ�b
�n��!�2��ԡTx�K�9Cz�1Ĝ�X!|TZ"��;MD8����A��2���9��eJyA��vK�g�d��<H^;�8�H��̙lB:��&����[��1)�F�u6]1Y��*w�QKm�.�u1��9;4�y`�}T��J�7m�i��c����a[r�"X�����(��$o�S�|�nS��Iݷ\�Q�'G��8��.¬໦��%��ê�ުC9_�M�)����_]G�6�uc�X��F&�o�J��çw�^c��:'����˦5�Qs^�F�츳jD_;�>ޣ�΄*��W��N�\�>��q�h��h���V2A�+w��7h�(�������v�/bGI�62��Wt!<e���0��`�I�Ht�˂�o�u�e}a��Wa�k{P�2KtZ����2LⰉ�&Wj�c�5�8U��h�l��O�;Z�2-�`�^ѝ�o� C�Ӯ1C��l��v�~�n���Z�X�ia����sO�2��^�&F�M��=�\{�����u��Gu�ǯ���]h͍@8!d����9)���ٙ�=;��'��,q��4��K��u�{���x>�3N�4�ٳ�_fU�v�;{%�:��뻒��B�9��/:tI=�|9SHtn�	��*��m�����W��'��%w_X�WwD�����,�2``u���)�o{QYop�� �������B�����E]�Le\�RN�B�Vq���7��7��fL!ڜ�԰���
�>�_9�{�}�f���ve�=č]�v&�[|�FZ���Ē	iN��WSq�Hܙ��$u�ݶh^!��f�8��gkAWبyPXUr7K,�@��SJo'�o����;�$�O�	����f_jܛ�ك�����&�rx�>���C��v��Z��;�%���,�w	t��a�:���(��%@�v�Rgcx��j^Gםo^�\'w}.�&��:���^sV������%�5J:�P���%=}h�{�\ʼ��e<��y���[�v��b]����)uX�ڛ���O'����C�f�[�uX�J����K��4X�L-zWd�V-����n��↺�V���ȵ��M)'W�HA0I�s!��V]&��Odz⡆�C��qZ�v��61�缐S�ۚ�^N���=����8���h����̊-ǷG֚4s7�:wB��+'%�Ӓ�
4_7}ǷI%�/g�aPOU�� ��a{�q�p˧w��J��V�V�,Р�=t"+��F��"Z�<J��^ݴ�}��D�.�y�ٷ��kۗ8�}yyWpI������؊]�pE^Y�"ڙ���~+i�CcEs��b��m�����/.X:��H�y7)���7d}�!���hݛV��;GOoS�M�"D�޺�����C�(4TUF��maXc�lAJ2���b��ċ*���X���-�ī��1��*��ee\�c#�W�.68�Lk-���[aR�W.*f6�#l�P´�*(��cm�L�c�GX�Er�����RQQa�eb��*�m���S2PDUPPW(ұb�,T(�f6Y\k
�R��
�F��eB�k��Ve���iEj���E�eJʘ��,���E`�����YV[B�����#2�aR�E��(R�%A[f8�1+%�kr�R�����XEPW+j�DZ�V�B�[F&fLA�S.a���J¬\��Qb��
��X���bfX�Ԣe�EV2"���*9j�Z��(�
�2"e�J�
AE��X�X����©iP�2�̹Z���
�Ll�+�2c+&Ze�(*+jV�m �"e)mkj�E��D@��
(
�
�
��r�6ͻ��v������r��ZDR�PRn��wا�O4Zj�w��wR�l�q�/F'}R�\��.��qM��Ǯ!��j��%<��'uA��i&x�C�^�\.��Ct���
Wí�ﳠ�wǼ��h��0����6�(t�MOZ�D���P�c�j����0���f�,�=֝�Dp��P�:�'ﺙҬk�
6ǈ���-���M����dǝ����y�>����]�{��{.�V�<`k|D�}X&�izz���cO��z�ܨ�g\v4u�S�ݯE4`o�Ӿ�+�"^K�����ِ}{\D�m�|����iA�5��nj��A��\�L�����e��WV,YK�+�U.X�s=��;�p�fMܝY`�H"m��$:n�89Kz�".��X�t�aE4��O}N��L�iċY:m N�7���{~�\�{�l�E�S�O5Q�N4���E��Ֆ�M~�(l{�^w���ɷ�d�z��� ��=5ݖL�Cœ�o�@#5�t�Eʤx�Ƹ�cYCݖ�vf8�7�q$o��c�,|���6a0�9ࣂ�oz�	��u�8����4�.^�%!i���qʜ���:���	�'/��5���}���/:wu���t�@-}�wq����R�����	��t�r���>Y�{��y\B�&�ǯ&��&���WàCy�ڃ&�u���� *��ۃ!d�j�5��n���$�s;≟{ir6
�Ă8��îc��p�en�)�拎�,׼!��"I(���pײo������VE\�:U�3@�=���t�iC<�S��]����Sϼ��WtRβ�b!U����	��h���kI0�E�uk"�0� �0�Z�hp��,~�D���Ӯ����x�)xj>�(Kyi!_f�+��9M�o��7s\S{~�}yۈq�m��)�z*�'���HW���m�54�s~-�7:�y��K�Tș~�弴��0R{r+<���৩t�}��T���������ww�,�dd^�xm����x�j؆����*�{1�|�\�N��n�����th��LS�o�^�^S7�w�ٷ��<׈�����#/�����A���>~A����Y�X�t��-��ǳ돃��'��x�<�����&�W�c����F�Y����{M�27{�}���|'���թ\YKH��u���[�E"���� wQ=At͵�4b�I^it)X��{��'ͭ��[���_�,]����9�V(��\��NH+s+r(��Ur�ɚظ�#�v��K@5��Q�aH	����)ku*lɑCW��x�#�x;L�x�j�J0����.J�KD�[t���þ,=C�Tݧ<�;m�"î���G�+s�B���^��:�i��w���G��^�PV�P�ZY��r��K8&�z�FN�{½h���f�l�#��3'y�9G��k�R��X�(u�j%oiEL&NP�+�N4=��;^*�yr�f��S�f�Θ+Ƹ�R�#eqq$����뮶���E5{e�d}�izc��EO*�kr'9��S��nՍ�1�ݮE�xx�ł�fc�/C��c�oy�s��h�#k��<��/�e��d�kֽ�Aڜ�U {�M-�S,P��9�{�&x�J�ge?<��u�ݤY�W�|����Y��=38�[�%�&��CZ��满�z���urvok�g[K��I�B8��'Xr+3Ox�b��7��ˇr^a,�$��ۦ�{�Zde*��v��EJM�uBr�=����Y���Fܬ�?.�/}!�:3�BSY����=��99Ԑ�z��"+s2���5*���,?�1f邒��B*��`�������R�~���;{Yu{�t�)��J�i������3����GX��#��S֖J���'sK`��'�4Z&��<�v�҇��,���]�d�+���H�k9kF�f��u���:�k�nL�0X/���7�\�޵/������	����v���yL��Æ�r����Lpu����L�4Nn����	�����nI�|���ܖ��_�,��w��vY�|6���<�����C�r�u�nY��~k{���Ǡ�0����$�s����y`��b0�eW�"�/�k����@�g-��������S5�����}������C0���}�:��
�Cn��=.��8��d޼C�u���i{ļs�����&��o�^��u�ӬIAx�"ر�'<�U�~���KKiv�U�y
�=䚋����fC��-�̭7ܥ[�ܞK%�E�ɜ��nF�a�6;iZ�i��\c,�¡&��R-��yы��������1D��׎m>>�ڽ��Cܰ1�i��jZ��E�ԫ��T^�w"En���)�k�v��D~����#����%�I��P���q^��<l<�Qi&��d珧ȭ0�M�QП!~~��V�G+��[��x��}��/v{x�~�t�
jvU��P,��W�9fj�k�\��״+.��B@��{�����-�X [uz�0P�n�:�������K�of3�VQ��>���1R�Pڂ�:ɺ���,�p��W�-U��Q�	ou�L�eeh:�x;eq�5�.��
�=]lF3,���s�
�t���e�{������.~]
ח֡t�yp����c����Y��d�<��d�s%a&v8�d;\���Nd���7�:L��4��С8�mX��8�}�z�1{�*XL�N��$D�3Xƨ����YͬW]��:J�P�+���V#֝����Œ�`~wĄ�V
���.����3��k��9L
�I*�"���h��.�����`K�̾�V����vw����kRC���wlr��^.y!=��I���y�/�i�		K/DC[2p�o��~Ӿ��>�LşwKE>�M4'"XpS$�t���X����h�dA�Hk�#�t���y�����hf�Mm�����t��E�v�<9�kݢ�*���Y�1�ݦZ��vL���Ϋ�Z�O���:��pVq��x��`�Q�����Zљ���.��L��wJc��ܶ���I^S:�E�}��\D�:(�����&��zUU�c�f^JGl�+�ZsM����k�%c���N`=�����x�� .�s�f�G=��&�ZU�m��CO�Ǉ:�ope�[�f�taK���E��~�CJ���9B�p�;�W'E*a`�`��^E��y���e_|L/�p!Qf�@Ja�v�t���m��z�"�Ԇ;������*)f�X���$���n�����ߖi�9=n�O��^	i��:ȣ0���F���s�]E���պ�wx����ʷ	����>\E�N�<�G�=��Oz�����9i�)}ClțB)���P��3��}LnAw��c��5��L��ƘK�oT����^.�g	2��wrN�lm��;:Agp�q$sU*�p�x����لÓ��=r��^�S=��a��4���U��:�:gY�u���śA.�]H>�o�C�֞�=�U��h�����/}�A�a�^�e���A.���Ϥ�r] \K�I���b��w�:m`uP�ut���1:T;T��z�tۻ��5��'�br�LY��l�[ȍ%�^�~�P*�R�N�SZ�{;�ex��}�+4���Tb�)Za��	��0P��$3�f�+댿�uL���5�I9�Kﾣ��u�t{+�f+/�h���OQ�B�TD6��qG�QY�k�c��)JD�.�^���l�#3y�a�H�ᖘ6৩t�}+�jq�!�����6���X3�n�D|�@fgܻ/wu ��^}c��.�糱8H��MA@C�W �v��Z�(�I�6������G2�u:�-	�t�K�Ns8(�{��8t�6�|[�cF��/e�%>%�\�BG'v�j7ؤ���h��[V�`r��[�!�}���ڇZ#��I�{2^D�m��<���W�ٌ��oo0nQ�c$��,�޴|`�ۇ�0���C~�W�����=sC���?Og���Ә;�7x��f9\pX��s8�0'���/}l���P�����~�e�c�h��[V#U4��M��eK���3r�{�#q��P�I3�h�[�gR�L07�[��:�*�I�y������k��� �:jm,�r٘�f��G���۶��fD�i�*��ӗr�5շ'3�d���z�V(p!V�p�4�YZY�����u,x�t���=��\��_bND�ݷ��ܼ!�	��[k�C����<�K~{J(�za0�jr�>u/�����,��t��uk�n�`�Oח|8]+�:���G�gʫ����W[e2.)��e�_�{N���<Yj���uq�m�r�M�"�}��g��r-#���.$3@�v[�\���GX�MnP��ܵ°o�{y�&=�ah�	gGm��"*��pRi��)�HǑS^��v���y�e�V������N�.S�� Н�l/�Y���&��� �PQ�����m4�[���yFI�zϦY�m^��u�;�ʏqv��};�_��R]kG��h�Y9I�໦����|u�0Լ�Οr�K�N�Z�x�g9լ�
���s�[���3��u�L�w�;%�X���@�CZ�k<����K�Q���̔�t�\^.J~v���+3OxSE�9r�ܗ�K?W��=�Q;h��������"
��U�]ˮ�>Z��7�z����s����dA�T�HUu���P��߻#��g.ꎙ�4� Y�v]h������f,��0RW��0y�ɵn�ok��=9�n�A�v��>���s.���K��@�/��a���#����*C���˪�e$���]�+VO}�����!/�[�	c��(g�����g��T���2�{*�/6�מ��������oy��3v�#������j��$�2����yg��MhC�x&����/*͕�3jbG��uU�l�(Y�R+ޫ0?���c�l�<��Y^{M�����PӾ��;�*��'�ܐ�-&��AU�+�j��ȯ��� �6(2�ٙ�;��Y��?���n���^�oͩ{`�����֠zkM�U��UC�X�(_>�I���]���O�z�N���Tw��;�|n�ZW�RF��ww�Ɗ�RG��<��۫Wvv��QU��f���ĭ�|e/��F8��$k;�W_�iξ�kMV�=��YY�F��0�۷��
�Ϋ���j��|��eC�Ź���s{�^M����E���^�s��6�j��L�{&F�Ն��m+O ��mO�Z=)���{K�������z�_��WoGydVɕޫ���~�E�CӕtJ��N�b��DV��?6;�&��Vz����[x3 �X��Q���zQ3�҄�^>�ky`��a�G|��9��H��쏶S�M�w��2�Au��t�yt��G�'Z2�MΊπ��<o�(]��T{]�3:�w�O{t���#'ܵ=�/�3���O�VL�Ch)�T��r�S�)^\O���)-�D�y�|�t��D�H��K�++��\��������X������l7�%��z�簃��|a�Ò�\9��z%�xU2:�����l;��	�P�����T�7l��HA��m��ݍ.%K�br�<*�I.��E�WT�X
Ϣ�<>�x�4�u�=:��O�Z]wݑP���<+�����Y��T�Bx}�e!��+=��ԖuNN}�a�`�w��Ke�W2���v���)��k~t#D�pS&��f�և{�h�#�����|�����C�J�̾j���we>�xtG�3ǳ��ܪ�`p�a'|k�z&�l6֊�͖��S,|�p>�:۱^FX�W/y�t���f�m���&we��[����Y�һ��n<�K�(|=-���)򷯯�}�վ��3�M���.�ua붒p�=�=���h^m����r��=�ǈ���-����ne�uN���ކff����ho��˪���^�=�bU��`�Pȇ@�ǲ�Z�'�����s[��{�u�C�Ӄ���k���%�	y*�2�{\D+l8���k~P��E��������q4�OK��gӵ�ۣb�+6Z蕏C)r�]N`=
DF�U�^����&��zUs�L��>u�r�? Է��	j�({�������gk�v��.{�:G��)پ��_�MH��R%�T"�u7�ܩ���ƞ�z!�R�3��A�W�uh�r+2�IDv-��	��ރ�--MC7e�.P�f|��|�+ܧeQ�K<�x�s�c�ӻ y䍘���Gx$GER�w�[Ɛ�L�w�0�rs�G��Y��9�<F>��C[-�-����T�H=��<q٢i�\��Wo���.�Wzab]�3V��<�k\�
�x&�o	~�`�+�2��c*W�VE\8����a~O޴���>߹�B��d$�	'��B���$�	%!$ I?�	!I�HIO�!$ I?�	!I��B���IO���$�䄐�$�	!IHIOB���$�脐�$�$�	'�!$ I?�	!I���$���$��1AY&SY��M�Q_�rY��=�ݐ����`��|S���_>�   )@��	(�
�
^��U*�T%TT($()@ +�eH�'ֈ�EP�Q*�@��yQ` c�CF[uT�,��ݸ�fj- �n�,�PmD\�n ���veB��j����-���շAN�u�*������3]�u�pIt�l       H��s�B��ʩ��kI#�mD �p
�Λ��Yb5�u�53w.�;�9�r�
��8��'nM�]�v�&�n�wr��QۜܹW]؜�KFE�Gus�Sp2I۹��M.����i6�ð�p�� ����Gn�3f�Z2�A�)IRD�@n'F�)!IEZ-V1����ej]Δ)!`�c���ɥim$�)$$#�m�b�$.MĻf��R�!�I����SU��{�* R	P   S�C)J���a0  ���`��J�`  MM4� T��UJ�Pb@    �"��	J�&�    ` $A�� &��SL�'��4l�A&�%(���i��    �G����S��������Y���QfR�o��@��-j>��������%�����N2$�y#�>EZ�j�H$#$����f��%w����Վ��/�S��Zj��oR����
�	��!D��/�t��"D#ꨇ%	�*H�*$���I$"�Gs͖}˸2x�$ƒ��88w�N�+u/�g;�@2�  X. ��� (P , @ qaP`T)@ P�*
� 7��{������I$8���'I0�4�$q�!l!0$8�Hq I���8�	���Hq��8�	8�`Bq�0�q CL��'�-�,����	L�BIHB9��뮺��e@0T@�PC*   �ะ 
� 2�@2�P ��v祦�_d��������9vܴb棚�KνOCҖ{4覜t��fim%ef��R����+���ҫ^���-͙6�l�l�� *pH����j���toC�w-=������8�2�@�c��wf���f� ;��K��é���i�v���-X-:x^n1Fehv��1M+��N�Ѻ��#R��Uj[+T*c�YM@0�<NnmH��4�=QH�h��/+9g ��¥���;d֖�ۢ�q���Y�h�!c�/[e��Oa��|l�/*I(UU֫29�չ�ia�l��4��*����2ie2�q��줟*cmr<��ؖ�>b�����su=i-1	{�`��X��] Q;�hڭ[Vڻ��V�^\�U^f%
��P�n��3��k ��Pf��hj˫��	�m��Uy��kK��n���d���B��ѳVP�p�4�����V�D�-[mX�d-ki���q�]��"���Ul� �ʳp[$֗�Me`��� �X4�Ws~W����BMԽ/ ��e���{Y�mI[���G����FAO$bJͻ�i�
,t��/,�5n}�w+~t��f�Ft��]�4�/�K�*�g�ݻ��B�J�V�faE�.���2��Fb�w�U,4)肮�c6���M�12�Kor�z骕��Rky���x�7\6�C�h�Z�ʍ;f��t�UI]�������������0��YV��x�;�Ib�v�8KCxwXY��vn�n�P�
��m����v�K��
�7HB�����2օ�(<�v�8�"�
4�݋A��7Q��J�����rTXK1��1B�|)^��*f[4	�\s�kq^������ڣ�V䕫lJ�z]�*AR�쒐���
���ǎL��Y.�:Ķ�pV�Ȕ/o-�7�Vҡ{b
R�a+�QR����Y�ֻ���E��	Nt-���/m��QF��t�x��ѧN�[E��]��F��;\2XI�2F*⊎a&�1VSܧ�]�P���Yop@>���!B�r��Y�h��M��n:g�vUWKG��;�H{oU�;7@�t�ְ��V�e��dV���]��S"
�
r6�VNٽSn�ӱ���ǲ<5�ம���a"O%��
ס�+�䭰0�P��01���S+#��$w�yqn�Cy[�k!Ւ]\�ٺ�ߓw��pޢ.�U����]ʑ�V�$�#֑gU��hjg6��e��\&��7����^"�䖯L,�Ց��M��zhۡ�T��&�^5˴���l�ˣ�
����T1��Xv�����gβV@wj2��V�B��i�֯�'G\4�CI����-��Un��C�vc�T[SD �ݪ�A>�1�1@ko2��\�"�=��� 5ā��eH��ӭ����*ˎ�g��Ɠ	VkJZ�3(�(ʇCۀ�ԫ)N���߯vF�R"�9z�hF�݌fD4�����qndO켲l�5Ɠ��㻖Q�.�٬a�R��P��5���ӝ��Н�$��Ƀy���5er=��,"����]X4R:���bh���j�hU-L4�Q�b�A-��)�CAŘ�ԁ�vw�S�wN�lR?�{
����F��Fk�m��!"ѣX���n��Tכtnɳf��kLe)��Q�mP�C۬j����������p|l�Y`21��X��U���,����D%�!u�@��ʸ�^C/�P��;���Lv��e�l�B�!�Gzn�*�i�rG�&X)bf: fY�W�<�厵����/(X9%i��ҥ� ��tM�vq�kP¤�/k"źZZ�&�nS�ī�f�!ʚȽ�bց�f�k�e�-�$��w`�ܺ(ҡBk�*��Ыh꿱X����V�5a���÷E��R��x���V�4�`��rٮnӬ|萊f���:��G4�Y��X��о϶�ʴQ����5�2[	��n�dҫ��B�7/D���Xl�����2��%֪1�Eި+0�Ca�Q�YY���[Q��{V"XF�YV]�Z�x��nH��h[�O�YE�g���6Z��1���_��3�W�oDWY�[�ٌ
8C��2�`�(V'Ԏ~��I	���N^K�׮xB��B-�SN��Ej�-U�R� d�i��4,�#52e�m�7	
F��,���7�N���[�js�m��M']l�m�KH��d��5�w�%:f�m��N7A�W]��'��(q|��,�U��qE[xL[�Jt�$���A�E&
G��P`��N�����X�o6,�N0��u&.�6���KF�e���Ɲg�ֱ�[a .|����3�����tPK��U�y�]�����uu�z�۔ל�^��T�vQ�ŷ�p^�m}~K-*T?����>��}�(���]�&$���FR%C(��%	0\�V���s�1�M�q�qc���e�7�l��:��lL1�LBKH��/�Ȯ��<};+�A�!�m���Q�p�.͔�.�1e�A�岈y|�`y&M�+Y��X=b�%��lW�J���f�(�w�M�Ώ�,'26��J=� ˼���b��t��*S��sIS��=tU��{��2Y۰0g�Y�MN�xr��%��p�Dd�RwiF��l�al�[�3r���]ø[bK�urrj����D��ĪnoP�j�������ӰUI)��<:5(��l#�#�A}7��{��gI4�׷E��͛�tw�\��� �Gi��`������h�T-�[�šx�J�e2�f�"2<��nĆ���F�.o7��Z�,%����(�b�Y]��ht�����@ºs{$((t f�������r���;p|�⫩���|TtG!;�W�j�9=�c�`�<�WM�@⎎*=ث�V2��z�<��	�G��=���l�`F�El=�4E%�_usu����o)���W��w �軱�R��4�fc�菉F�nۄKAwN�(?֯c	q���<�wvN�,�j�Fr��rS�{��N�M�Z)P�y�~�mM�ɮ�$��8ݾP�V�����ԡ�M�(�-;�=�{���V�Cի�Spi�t��L��5çL۰��Z%o{sP��ՍWV����qxP�u�:g�Er�W�r	��V�[�����|Dg2��YSxộ�p�Lި�Z��LA�� ���f1��;n�l[{GbQ����4G�0�+�ԟ�ɀ��jq��rr�9��\2�b̦.6s�6�bu�w$����(��5�	�	;N�\9Ț�֗-�D��=w)WR1K8����{w�NF�;˒[sM�?-�.԰N��UrO��w��+����'��:WJy����"��u(Q�*f������k'b���j�tv�w\x:v:؆	�(m r�]�ۄsY�ݭMp���Sj�*̜_��3���D��[�4k0�ixՌ�Β,�Wɔ{�D=u�Xˬ����r�\��Kx��nӰ��3> *˖��\�KJ��2^�R�k��x
�]'�K]Κ��^�xf ,viq�f^��F@)��W.s{��[�*d�;din�;37��&��������r�2��mrYoi�y�V�i\w�0��s�U�f�M�9�w`���ޠ+-�	�J�����.�(J{ ����R���s'0��L�V:q���UL���_^m����%p5��Q���|:��9g�'�,�Q�JNC�:JK�Z�7�ސA63��/�E�v��	�B��8�z� �d��ޣ�y��-��e+W^xʗ�:�)���wUM)8�^oD��1�SIe+Kٷ�AS�U�W�
W'mo[���'��(��q�@%)��';�oA�Q��A���7:��릋�C�ʴ��fI��j�f�J�r=�J�Ѭ¯��;]\+����͇���"5�d��c�`�B��aweIw��m�����w2QSo����nW��q�y�Z�3p��:Ň��S|ͱ��W�̥�1�Y�4F%�0DC��w]�nh�.�Y}Vf~}���V�q�0)þjʥz��݊ơ ���or�c�� �z򜹗�l��ӂ�����ge`�$yi�^t%)]�@���۷ւZ/r�2��ftޥ��<�7$�rP�7�B�C:w�5&��)7't�a��7Eܥn�I������[A��=}���W�5�Ԥk���ai��(�:�F���(�����s�
�36��7����ٶ��/�׊Gb��zT�Yowu�0�4�Dv򝟚(���+j�'c.�vîYŦm��4�e������n�Փ:ieF`]t���Eݥ���ɇv�r�uL�1�r���GlmB��&�V��愻"I�����=n�h���L��(�o����8���5��єԡ�]ՙۏ'j��.�n�r�_Nȳ#��g%e��_=�.Dʒn�y��!��vG�C��"m#HN�����fhزv�ܸ�pt���|��k�B����"��Nz���Y�3v��=�\�c�$�Φ�8��ٻ�~~88;�5�R��n��~{�o��A�l�WΕ��Z�$��߻K,�r6kܥ��yD�XȂ!�r)>�f��y���R�+���m���^j��➋��D��FZ�u�tAC��ʄ�r����,��o7�+l�\����Y��o+5&�"%՛�DPa7�k�ەu+�	�-��w�Xj����<@��[W�iR�)�f-}���3�"Z��ݫ[�]��C�,�LT�����S]]/�2���W�6�U��f+5a��;�C�۷x|���ٔ~/.�
|�*���0��b9]X{�vkGfFF�Bde���r<�nIrI$�T�I"�$��%I$2M���I$���sw���0r	ۨ.��q*�:�-nv	� jVp�8������\�F���#&F���ZV�ٔ*���n�&T�� 9�.�RD�e)5�z8�fU�P���Z9�
�&��I��ja��c9=�H�1�3����[�Q�
�3Em_L��L�i�1V*�"E�$�5��wx�%���埯����Ewhn&!��%w%�4갌�A����=��IRI$�)I$�JRUT���JG%�$���UajLh	�X{&6.W�S5�׶�=�5k�\!]<���J����{�ٮc+9��R�4L�!�r��Gr�g<�p�vd�]d�仧n���e��.�,����gRE�F�7ktAY��,9���4�AVu��wj��E�y�|s\�D�<����bPv�//��м�%_(2��`�o����S��!�&I$�J�fd�d�I�$�H�%h�����x1�Ws�:�P�I�w���y��Z4�
0�`p&�U�]ݶ�2��٨���D=�%�W�]�R3�ejܲ��c��;�࣠;*��7f��on�X�WkM��2o_"z��0ł����U����,��ʁ�y՛��ĵ��E�7�JB
����g(��P�a5�y�3��e˾鶮ݺ�]'�I:I �)�d�ʒfd�M�I�l�HD���c�5�{�f���e˷����S6��F��#5±�w�D���
�ub��� kwt5ގ��IupIZYxN�-�w�]u+mK@S0*��{o,�݁3"�.Y=�`!�:&n����1(�'�Qx�Ifp��.c ��V
���ǆ��5yȅXz0u�����͐�0Y�l�����7:��n�k�:4�W:��>�B&!��ms�����nt�H$���t�A%�;sd�t�A$�	$����[,w��P'�rI�p�7u��tA�t��M�gE-�BT�2_q���e+a�K,�h˵�ҹ���뼦*�b{������٬YS�3�:޻����4�Y�~9�h�";p�w��Z!�i�����m>ZƵ��78�j�j�*W�o��b��Z�i�mg;a�+�P��_[��&����W)��&�ƙ��uLw2�uR�h�	&�$��6I$I�L�;rI$�I�I$2M����7�r�wM������8�A	k.GW���J�b�D����ը��nr��L��M����T�/�v�Z̨�Jʭ�����N� �;\�'�k��$���9d']�Q���.^�Nk�Ѽ�?uF���H���L�b5�n�:n��\x���u��Ⱦ�x�^��jڌ�R�,&���*�w�j�}c��|kV��E,�TQ���\�I$r�A$�$��:�I�$�H��4���2�`�o$˖�F���d<�ﲎ`B��	�Mf���;����tvu(�*"�\�h�����+��sW=ll���N���v�΃ރ��S13(�j�yta��Hd�P��E��F˃�x4n|�f���J�9SU�.�Xqb��4{�T�2��O��,n#��[��;7_v�46�̫d�@,�Uiy�%��������r
R�6��aZ0'�{����I$�$�C$�$�ݕ$�I�$�H�������������9��"O
����]���b�֬���A�Y7;zη�]��������\(�%tk�/r�*ЩB��}��`�gN�x�뷋I�Hŕ�]8	�Z�h��r��M�5^Gwٵw�`4ހFR�*��ypE���[;:"i���yX�7�[F�9��v�܊�-�.���M�hm;#�a���n|o/kٝ;�!�$��!ue�[t�]C��gv�N��fr�^l���L�ŭ;h�֫�ꎙe�����n)�����]���j�Y���Z�l�ڦznӂ ̱�)㘃�}��
�o��;:p'*�ֵ��L�{t�SǛt+6�˭�����N�v�2u ��ܣ��Ȝ�%m��oj.���9C0mX�}�*ԣ��-<v� f;xຜ��11|WG�s��9�D�f�V������B�������J��{�uk=3�������  ����M���$����+Rf�_�j�F.�hj2M*G�h�>�F�����G�KiE�J���YU�Zb�[�J��VXb�M: ��*d�M3L �c��,�$�?���%����-�M�EQn�1E�)j(�JI����:4X�F�%<��^3���02�㞹�J󫲆���xLx�CH������o���nm"�G��#K�T���m妯yCe��U��3'<`D��QR��k��aj��_5bYsIP"�����R �z��bu<�X?iI����;��`ڔ���(��Q����`\r�w��Ηה�=�E����rT�g8;��枕�9�9e�ڒ��0����G1�ǡ�����s��s|���`故+ ��UQUG+�&�V�E�t��]�Z��zDQ�m���F��{޴ei����R4�P�n��kТ���Y)4�zֵ�Z���Z����������b:SUP��Im^��i��V"˺حSZִh֥.��j�m��R�1s(J�m�wWMSIiT�|y��'���)�}oo�վ�p�1OM��areW�ނ��VA�̔ m�RmW���k_�R����������X�l�]�<����ܗ�%^�v�e#Y}uα���1���2ʣ0��lsS��,��wem_�y�V�H�����٪���Т~������D����Êt��n�hCo�[�U$Fg�I3Q����3�ڄ�D��x���:�#���Ֆ^�r����'<�i��8�JT���w_Sh+ q�o��ɮ��^����<Ki���/#@�7]���`��T3�e�L��^v�
ܛ�@cu��5�����S�u�g_f#[�FG � �E)�<�� ��y��GnϊkUL�N�{~soN�K���1��;�a%���-�Gw�7y�.c�6���nĆ7G&Ѿe����ܤ2`CU\���w�Y4��:��K��x=�K���z�[�vvZ�����h�f��m7�n��^�1�Z
m�,�wp�(���$��DM�_Z�<�P�s~�{ڴ6�0�M��kTUw/����/M�!����l!UV���g~�u��|�<�4�b�e�˶��:+�����X�HN4�,��:H��#�D	[����}/��j�1~��l+B��\���sr7�gG��7S��Uu�ˤپ٤�w]�ɤj�+VS��qޮ�z��g/{��m�j"�U��S�+.�Og]�u��n�F�#�m�y�5y��z�g�;wTw�C�c��Y�b�&}^v������r�>�>j�ѫ�H*�'���)�N�sSC;|���]f�<}~����޻�I~����k�9º��)-��-�y���M��n�ݫ�^}�N��BB�"�p4(&���c�o���=����io_�ݞn�)p�4�'她8�5�����k2�ea�,U~�a��\@�׹^g��ڣ	��k��i�,���}��hS(m��U���,U�C(�/t����sUb�����
�%����.�U��	IIBO�G��m>w��;��ƽ�;uڋD��T6��Nw�1����}��^K���/4S-���z��k���h���1�_SY�m�̳��5�2n��Ax�U-��'�r�8��CƽW�������f�9�-�Q�63)�7�{;<R��no�FEq�T�UC�u�b� Q��K^��&S��Y�6��R����T�e�m�s��՞�}��n�}�⎄5���~:$5Bv�]{�c��8}6�P�Q�G�������v}ܕe
p�x����>cG�]n���ú�E��O�(�e�QuYG~�1�X*��������ܘ��c�V��#�E0�Я��aV��5NyU�+,�ˉ�0���KG�+���^��Z�u��y�e^=M8@��N�S��5目w��x�v������GP�i��3Xv�����o=����K��!�Cy&�.7Ж�ܬ,4�I# ir楽Fݫ�Vo�CU£62�}�E+�y<}��
��f
L�4�KU^��V"_����Z���sna�y��]��z��[��d��L]Oz��W�������<7M}���@Dl��u�<v�5�s����PV��i��E2�3{u��;Xݛ�=]L&3KF(�p�8����ϛ�;��#��
e�"�TL&+x�u�[�v�i���p`�cUxu�9��uA�y��,�bv��WR??��V�K寬m��u���Ux���ս�L�`c��5a�#;q5���ە��W�]��Ԭ]P�u��@SW7~u��X�Ab�,���:c~9y�{�ϗ�g}�(�u�x�]
���-�W�A\����/�AX4R`G���_p�����gEh��b�ML��8oZ�y�)�;�Q1B�e9N���+O1�c^ֺ��R
<�QBӺ�;�m��������M�ڣM�����Q�_y�ϻ�E��ͷ��ڣ�igY��=��� ��e-�h�Ma��e�M�ϻ�/`˨{�(���Y��2��D�:����m��TW�d���&��Wtr&ʒd@��n����.���1_]3ɗi��co��6�vӡ�6Μ��|2��Uv^?i����\M�0�!��Jt�e3<Ƶ�k]���èe�,�O��h�1����ֽ��e5�2֪e3�u^�D�ݭ{>��V>h��֊�������aǵ{��쇷E�o�'wY|�6�fi��X�2m�z1`�\�u�T�y0��y�xsZ�a�:�MUO2���,�����ܧƾ�3�ߵf�:�J����Z<n�?s�SM	�A�A7-^���զ�i������}���c�j�W>�?b-��7#-��Z��r���7��]u�C��"�me�`s9��U@�ކ��M�H������\�;fҳSN9�O#U��@UhLtsO��|P�U����x�L�k;��32�a�	�˟Q�ȅp�\�*l̎W�PO�0���#A\����������a��m�0�qGY��{��׫����K�/W�q��X�=Mo�絇��a�]n��Mb��K��o��tv��9��u��&�{�o������@=E�?�����{�e�߅�O����v���/��������1K����0��eQ��#7�~g2\��i�=�?n�}ff<������f�h��곈�Ϭ��&�]1Rj��X5�V��*JQ���A2�:�9���g�G"t������Vj\f�T�wp��-�xA���b�W�2����ں�ݾ�{� n:O����Y
r��:���ں�I;�8R�`�Z|z�37��f����ұMŞQ�������:�Z�&=���/l!��8�l(��J�D	�Q���!�؅#թݺCq����J���2�w|�)�:ڬ9�j<�T ���򟴉{�G��}0�.�aY�[n� ��ȓb��W�yf�Y�ֲl�q<_�.����[����59(�Kzh1�wE�]��H�Xtu�W^����᎜��wK�l����U��mEՂ`��L��Ĉ��t:ƞ=��k�����<Q̖�U!I)� �H�vZ����z�-�X�U[*�޳���j�l�--�5E�-�^�����21B�X�!i
��ZѤU
(���eU�jۭkZѪh
�[
le�$ֵ�e4]H��UUWV�Wwuֵ�����i&�PX�W�kZӦ���T���cu��h����V�n�VO�+>�㽒��}�_R1�+���E�Ͼ!����ڏ������I�Pe��5�b������l��L�ɔ3�E%�:Kpr���_�{���r�to޹���4�6�e]}���}���q�u�:�s���[�����
�:�B�j��Y�]����5���b��<�3\M2�W�9f�'ڠ�~�^<�9�c�
B���3R�<�m�Փ���ky�q�IN�^0��)�b������m��A��:W��>�5|�4|®��u���^s���i�]�7Gک���5^U_߶�`��<2r��2��R�[�N�@�n��[ޘM!����)t���%�{^qmEb9=UB���6S�Ӵ�gի���Ç�QR����N�_|{|CS�XS+}�a�)��}�W�+�p�h�*��b���UߍG������Å*�TH�����Ō�/�zΧ�\M�z�cve�^+i�>ԟ���]ec_>5����A�*�?M�/\�Y���L�gl��k)Ǭ�*f��e�+�i��i��y���*|���o�ʳY����:��\����ۭn����v���o}���S�ZJb]w�%>��z�Kh�F"4*��(�O�;��Mm�9���1dM��V�=[�'�6�0z|�ԩ�1�Pg��c�]�}Ͼ�޹Ϟ4���6�M"��+�
��Y��S��~7�h�j:ϱ*�U�i�*|�w���8gS��ZKg���əS9)�U�"=�Ss{_R�s�u}o�\��I��W�__s�jL���Zr�&��4��U��0z�I���z� �e�\�LE&�%�v�{;�v��ު�M=lM�4U~(�J��F��|Ǝ�*ZV��AX,U~9��n��k4���Xk)�������W����Y��%�oN5Y�c	�i �g�\��C��zXRF]�|�&�q��q���W�ts�W�K���r��1~�X>�Gv�j��snP��ɟ�}P�k7��S�U��U}��QSw�,:����h��OFHk�y;���a��)���g�{�c�Nٷ}�����S�eɒ�O�W��}���hP�a�J��[z�)3_Aޝ�՗���2�3o_3N:�O=z�&�Gƽ���B'~�O� ��U@�v�ݔq3�{�ΧYL8&���Q��E}_r���o����g���W��S.{B������@��*W�����7����5/�����*��@Ҳcx*U1��k�I%��9}��_[zλL'�W_&��r�F�S���E�ѧ��b�&)e
�^��ߜ���T~�Ś8T8=A_Q��޹�p����ӶZw�S��l�.�̯������2�3��(�u�J��V*
B�5=�|�߻�3֫ɚ��UA,�������h�?-+镔���V�ʢ�_�u�֓�,E�	2T��q��=���|�:�N�;y�}�����z`I�hϝ5_o����A�jDƱ��7��)�u2��w5��ٻ݇~��O�nN{��t��
1C�GQ����҂S��U����Țo��z��o��캪B��E�V���<O�__y�/��Ѵ��h�(�b��FQ��~Q'��/'��ӵ�Q���.�SL˾Q��s����������c;�g(�����tp�y�����G�S.��&��|�M�X�ӎ���:�u-�6��Pg+՗(��K������i8����)i���}�����>BZ(�xTƐ�7��Y�7U;��e����!NyU��o���w��<ٺ)�V�<g�<Mj�ᗒS���#�*�B��fp��k��鵷����N��y
���`}����$�  �&[���P�DW��Y��ӯ[t��y�;�^0��m۝�����V�~����@}xt5F�B�?W�s����F�ӟv��^>�&��mɇ?AF�����s	���0�~�¬USi|P�~3vw�'���B��O���v۔�>g���xϾ�s�	�a���ӭW7vq���f�~���ۄ�����a�iY���̡�����}�N��CUx}�w��G�����CY�U)�a�����z�W&���ΰ=i��	ZU�,b��b�2g��yn��^��C��tu�#��ꪒG'�������T�x��9�r��^s��{���+9��3��8��NN��|��߷��������^��(x.?X����>'�x����/��
�f��1�Nv%J�Ӽ�G��9�?t�g��eΪ��><���Q��)�N]a���gn�3F�ƻ�O:��'.��ɯ���NXW�7,~�7�~�}_&���s�m��TGi)�����w�q�(�t��k��ӕ)0�f�^�q����&S(��͘�w��h��{�׍kVSB��/�"�z6���ʎ���⮬}H���^��[��L��d�mN�Z�D;WD5>�1r�#&�f��z��|�v����{��r�!�9�f�!��dW��t�S���>#/"Oӵ�L\��ܯ���1�k3{F=���>���}	�"5�T��ξ�����Q�:���CR�R�D}t��c�b�W�1\9�\p�o�'�n�����{��lϪu���Q�վC=�m^9�g׳ϺQx�3�2�LT,��W�+�K*����{�.�	���J~���tc���ڃ���F���,UZ�����0d4�V���n�Q��$n��!��!���4�Twr��-Gr=UR9~vo����u<�~Wl��Q[�m���=g�ow3��z�L<�o��GR�m�����o~z��f�i�����a��ko=z���ߐ�TqTy���L���(/>�+��������T�(O�P�㞽�3ӭ>�}��g��!�h�5 1_x����x���IX��?������2A�MI�s�p���ѹҪe�}�x��gY�L�9�}����c�������Sfŀ ���T!o�k~ü�{���e:�,e������R���T���x��=PU�F���g:S��h�Mb�0T� n�Wd�n��T"��K��T-	�^a���-���niӶ*�����v3�3J���Wt�6̭t�++��t4�0��;���\ݲ�7�4-%��J��h]k]��9N��j#�&u��kD��S�F��G��U�h�v�v⧍�6l��Yx�Ԓ��P�H<�L}�[�|��&�%�z5�g:S9ӌ�kw$vGZ���zf��E���[4��`LǢs�LztB���4D�(��qDo0E|�����%����Q;�7�p,w'�*w���9�3�i��/t3�0~�i#���vdW���'o.�]Y�e*l^���X�BWM2�gt���
	`��{\�\�>KuLђ�u��%Y5D�V�6m^�f�u���N���/w η,�F+�7q;m~��ұ��Z�E�]��3;������j�`VCo2�@�?������b��ߕ�Wԍ[)R�A[�?�ɩZ�[(���Tj��Z֦] �Eue�S)oZ֌����"1j+
ֵ�hEA�,��R1��kZѤ��Jh]2�U�ZѥTEE�,�E�ZֵT��.�-�we-�^��hP4��S�����˱�*- S�#)�i�=޵�~�1����� �CF���N����I�kLV�m��X��s��6s�ؐ���$�Uu/s��=�s��!�Q��m�V�)�m	�(Us;���3F���M%��I�����`�����!�Z�O��N2�
AC�,6
L�������)���i ��~�9�2�L)�RAd�*Z�CUD��� RA`��
��iE �4�82RA@�RM��}�}�b�� ����AB����T�B�C��
AL�S��jH,�2��2iaO����]���(�3�n(���Y��S
g) ��ì�Xi��)�\�)��)��	��b�R
��$����}u�k��e������)�2RAg�3t�AH) �)�Y����-�|����2S'YI8�$E=�޾�q����JH/�8��4�"��)���
AH)6
Aa�
@QH(ZJHUQ �il=��Rg���}����08��Yi�֜n�ZAC�|�é)'P�����R
l@���$����l���R
�w�ާ�u�d��i�
@�S0�i
�,��ɶ�AI�) �k�Y��Ì) �
A@QH)��}������M>X]V'Y����u�o�=SS�����J͑��Y3F�ԡ��ꪑ��I�XR|3,-��Rd�S%2f�E���*�,���:�-����|�al������vB�i�d���O=��kp) �u))L���R��"ņ�Sm$��QH�ì)��RAdٚ��Xm�TAJ`S1�w>����P6�� ��� �4�L�H���H)��O�8�JH(*�����}��w~�m �)6�I��S �A@QK@���SH�Xa�?0) ��%"�Y�JH)=���׹ކ���i �A@QCI) �su- ��
a��P�Jde"�RAH,�%$gF��z�&R
M�H
,JH)��
z��L��P4����Y2�O RAB�LXe�$�!I��'��|E�XRH,-�H,)��H)�B�Y�Ԗ�Rq�P2}E��]\�
`m�-
E ���w�W1���Ɛ8���) �����L����Q ���Xh��i���$��'P)�Ǹ��l60��P(Jx�H���R
Aa��X�ZA@QL RAaۨZAa�u��) �#���y��JH,��B�C�)��i�d���,)�d�������R
Ap����aiv�hJd`N`���;���y9�}�g��V�,Y�����,+�}�׼=[���h32~:���z���/c���&�ͤ��aLXe�0�
I�) �a�i,���Xi�$�$��R9�y�=��oܑ�Rq
al7um$�9`RAC�m �m��|��i6�R
AH) �S) ����o��[ �I2�Lި��� m�Ap�i;��S䂐R
AN%r���-!�Q~���۾٫�[C�2���f\3�q�Hg��p��T>�>�D}=�o5Ǘ��;�{��0ͥ��L=N�Y�v�/D,Qg�\�¨��B�"�NS�u������ԯ��q�0�0����ޟh�>����PV��������^��T�rZ�pc��MAR5���.���Ϝ���:��8�Қ�#wv�rI�G.޶u�-�z�3i�	�_W��������q>p�z�C
�6�=������_��cYܐ�rnڗG��,�vc�������fM����e-}zDJV�p�	�Z�����c�׹3һۭߚ����^}�k����@�����uxv�0�e]��*LX�1u�gGޣu ��j�����|�`���[ܸ�P��R�>�x`�He��%Ya�*H��US�w)ft��*��>$[F��7P��b덽nP��rz:8oLb�W�Y9\k^?�|h�R_�����]�.�������H,�����U�Z^xz�;�u�~p$|�f��ca!�V�;�;zhl.��+[n�e�hS�	��M��о]h�9|yM�i�>eFo��oG��ɨ*��-`��̶��� {�j�fFg9'�Uk�ϹC��왴��Q?���\���R<��9�:��s{��E�(#0�:kx#+ �B���b6��fvt���ƕC�C��z�k�9�C템�˫b�b�B6]�����(�>�}=�lCݢ�
����{Ńb���+����Ŭ
�u��'�7g�vLK���h�$f5H[�����W�����M�rB�d�؜� ��U�w����ꉟ�#
i�SC�d�Y���ӹ��)�l���8����=�&O#�Z����G�"��|�+�d@g��I��Sv�+L_o+rK��ea��ܳvv}vo:������1@��pS�8�ҽ�8������C���Y�F��4�J��k����� �h������61sB�t�����,�4/^	M.bd������w����� ����2�a����q�ft�e���43ss���@X1V9~�����B���
[����:)��R&(�׺L,���>X��P��?g�c�3�a�CJ@7�^F�X��X��PH�߀h�EW��<�Ob)/�93Ss���D~@������W�}�%�A�ՠ��ܤc�-�oX�O�߫����d"�b��=��)���oq��������x���pP�f��O��RN:z�j��x����F��u�s�c�Ϝ����*��7��A,$o�`������\���NH݂N���
*���♮�z/h�z��xz�]ݜ��b�N��N�g=|�K9$��'��r�7{��[��k(�`��a�kx� �=�Y��Zw���e��G��못�wwQ31336�H�?�ڮ�������e'4�}��
~�3����tOY�h�+Ӌ�bSE�r�mc�Тl�,����L�k�{��.xs�/q�����ˠG>Q��P��Z<�j���[Y= ���g�큁�C�}=0{��Et�y%�����}�~�MtN��~��t˝�NѮK㔦�t�(˅��su���v͕f1!�Or�-Y�W��(��G>Y.���>�9A|k�u�E�Y:��aׅY�����Wθd"~����5��j��3�կ��fN��U[-�졖J�Qȭ���1=o9��tu�x2�)�^�1�#�����̱(]�"�J���=���0�V�S�q��Y��k�]݃	�v�Oz�acf� ��B��86��%�hjW�=\o�ӣ��z��!)u	*�� $a���^Ewfn�u�ve�� PǙ1fF�//2Mx�u��G�l*Q͗ߐ�Q&�IƸ8M)1�,�{g��[S���M&�����ռ Qo k)ST���(��1ۻ2"�:���x%�wQ����Qr]�u��owv����X�028A��%&��p��M��iB"��d�H ��װ;��ɜ�Y|zoWl܈-z�l����R,U�[l-���%�CtSW�}�**,U4�cDX��gZ�+A֬��TF,j��j�UT���kZִ���ꊊ��U+Zֵ�j�Q��n�m�ֵ�֨)�SKZֵ��(�"�S-2,D��Zְ�LX"�f�DADT)�DK�y�x�6��_\ۊ�l�a�����|��
!�}���d��7߄b#��ǦP��A�e�%���q=�o�L��{�H�eW�O�C��,�E+��&`�,Vg�jݤvw�Wސ����B�f�׬�U/V�6���Gi���R�
�I�[�sdWv���K�3���w�����U��3<<�R9�w��;���o�]�i��ek�QWn[P�Lu��Q�9}�&�/���C��`�(((
�;�������mp�Z;�m�/Z����xg�Co�C�ӧ���Ͷ4its�H��/d��f�aS6V��7v.�h���1ߡ�_��2�Pz>w�Zy��{̶=�7���ޝ��/YS�?��yH.T�D|v��3�����d���-;9;���@a�CŇ�W����D;�o'q��Y�#���bd��[Q܎O��_�_��EH,�d�@P!��������?Ԋ����5��ӫ��v}�1j�TNE��ⷀ���Y�� ��E��X����h�;��p�Ufne\8gc��ޮ�����uwtin�9^m=̡�l6��Y�!C̒�	rb�o�0A��'��Ӛ�k0aTx{`ݨ`v����8����(����ܕ��Vnj5�:�'۲�Ns�s�\���oY�����XA@@P��H
H�9[��N���߶X����	��)o�Ķ�C����_��icr*2��
~ղj���l�rM���~���<G���p@ʽׇt�V�b�ֶ�
�-���97��v96��= �~����|
��o֊�Y�-O8��u���d�#ׇq�XNa�]�u������0Rf@����GYϓW��{��~B,��,��)`F�U/���z�����}�ĵ�����L�߫/
���d6�ǻ��;L𑡌�������"�e��ָ�]q/(k9n߱�yY�OX'c����U�ȿ�@)~#lA�/=��3�s�۸�upXp`S�<T�6���آ�=���v�m.���o����ډά��ބ�ܮ�����׫�J\]����ʲ۝�s��@?0�(HE���Fb""f#�m4Я���(W��&`R�O�G�?P�6,D�z�e�:EOs��GlA�oܳ_�׫�^���NF�``h�%�NW�25�jd���K�ξ-�SӦw�ڱ��U�[�ɼb��Q�0���U[����3ѷ�W�S���9�{_Q^}�ǝ���kmF]fgR�=����S�4�~�:5���A����������P �d �a �B���_��k��O󿱒�}�;��ެm�����Z.�c�������~,�y�cPΦ�]�-��\j*�>]�j3>�ٹ�1��s@�#��-�Z�_��xcn�F�+e�^�R:<����<hף��;�5�E��:�w�\�Y����x�v������8�j�v�i];b�zq9�v�S�k���]��	��@RA@Xd$��������~�k�x���:�B�=�xN2|3xǱ�������҇��~���G���KH=/x���z��,xq=}Y��1G��*V���e���Twh��#��5����s�a���b���"bz�_ܰ��j<���T�JaJ����Y(�"��xؼ�}��6J�H�}�����$��XE�,��>�����S=����x�� U�%W-پ������\���X}I����(�7A��9�Y����\_ɂj܇6ݮ���;D�Ɠ�]�F�=%�Ғޯh�-AG�]=Y�w�ޗo��`����7�&:�;�d3m�=�V������ς�V�$����¦+M �o���I�n9�po���7��{�Ї�`
H��P${��_���q���1��<��8O���ߧN�X�����t:~�{�<}������`GE`׹��K�){�+A�Н6Y����Ǳ1}�:�^�2{��"w�N�mFM����l���5{���g4{Ӹ]7��D;��}+Kw�-m��vG�DE/i�8ެ}�2�|_��c�S7Mb&��i=�+�*a8�X�vh����e-��Ԯ�F��㔩e�ō��.���G���B�T�Œ���5I��Y��-Ì�
��v��4��)�VC�Z6�h�3)�T7����J�Ɖ�ѡ�$5al�5��1*���Z.�r�q�Sl�b�ԭ�v����֕����´��w]��^'B/�E'�E
����ol���p���J�
�+���a�e
8eD�� ~���6{FΰKp;��W�;�줚��NN�B�!p�hW�D�&q�̒���
�-�l��¹|�3�K��F$�V�r4��M���f��(�OGX��FլҤ�tf'G.��k�����uTUgB���]}����I�d�M֒'GD�v�h�G��Z:/��ɷ��3�p���Ѱ�E����f�kj�sٳJ8�v�O9��eo�n���ͩ�
���1A\4#\�ѥ����K�ֵ��1EAӭkZ�",sU��(�^��f"d��)�U�Z�cQ�&j���U�Zј�(E)*��YM%MU�Z�Т�j(�Y))]U�Z�csET�2��P�5T����h�F��	 }B� �O���w7>��tR�gu\㈎F����X�t��[^��op�X��+g3��*_e�r]\�/�������d�I"�"�
H���o���w���#Ƃ�U?�*;�#�Z�jo���kJ��8O�XM��l�٩^��T�o�O��݊��k�V��V��~J�ڃ�n���)8:&WB��/x�v���Vg�N�_��T�n�<��b�����ߏ��|�#Z�~��1|�U�����5x)b-�6��[V3%j�Ӝ�����%_(9��@�]���� |�E!,�,�P��}�q�_~���5�߫��y�T�5�p^-�-�|�BǋC:��:��X���G��R�Q�b_fiV�Xޣ%�v�$�}q_5YVJn�y焓9˙h`@mY1u����;��F7�{�}��'��=GX��KF�f�\^
�kr���:y*>�W�+�4�ٝw�����G-�HF&�d�2�y2�ҕ;����H� Y��
HL��}�c��oԈ�?�xtvz������6�V6�����L݋�L�>�U��3Ҏ9�m�q��:݊��R�ݛ���h��`>�C�;���oe͈ZLn�ݙ~��V�]�d4��7(J@���e&t�ǌ���yo�7)�ؕѣ/�������wcy��]��]�[�EN��Tc�}�r��Y�{i9��;���t9�u�s��9����I ��A@�߽�}�?�u��pq�2d��&���`@�j�d����y�]]��VO�r�B���ܔG:�&]@��Ҭ��m�ѯ�����הSP��9���I�ط��G�ٛ(s��LXxnFP?*�(	Xb{��o�%�hkk����Ӕ>8鑂�m�M�މ���k��\��w�$��k���x�ʜ�<��NU�ȍX�˔97�\�����@RB(� ��̸o~�35�*g�W�]������ȠO��=�p����VG���3�3z�3�s��d.��A����"k®5����ubf���l�T�5\����Qu+�+�F��G�,�]W�-ݾ�/ï]F�1<BIh�*�cs��5�.s��k=�뭞��:*P�ss�R��p�_�s�Ʈsw�z��i;]��s��+��{�!?2E�(�)d�	=�����:3�qE�����Z�'�r����PA�����ݍ� �84�j#�J5�]M'��S8�����O����q�%����܂�us�����������dĽϨ���Ӳ��FK��?Jtg�g�}��@�)h�53ٙ���r�s�ĸM]X�c%,�Z'?J��i�����ܥ���^S��\����o���H(��� ) ��_g_~~�����%����r�eG���ϊ<�f�6�

����+����%p2LM�;�ԑ�(\�z�e��*��� �
�ǽ�0T�:0�ۓi����7+eey��ߪHy���7�7lm�dv6U�>��uT>��t[�ǝ̼�5��T$D��[��ޅ��x�~���4�����6����A�e�qR}5+�Ŏ�(��wB[�p�s<�x���?�0�(�)�����m�������e��:2^�j�͙�S�7�ķ�CN�
��4e�<��m�H۷� v5�3JU����O����ޱ쫣[s*�>7H�p7]zgrIsb^�M�k�C4�xȮ��ݛ�{?w�N�>�`�k<NV���L����;�`~b�9�#���3һ��/&��:�Gdi���L�db�y}���{�_y�����H�
H��X�@1ܛ�k���3�oߝ_q��De]�7��dп�>����F�k��S㢄���t+�8}�74��wl�̻���\�j�e�vrt��� շ��/3�ߢb\3��[5�F�z��;��D�y��������?��뾸C�l�嗔�e�V^�m����6�	X��W`��j���|M9lk�r B��>���2��?$Ya�@��=����4�^�l�t���wL.\2�z���k!��Z��	�}��1�7&�M6��س<{Z�Ö�(׫ìh����_��[,�l�""�������-vϦ�_�/ԑ�׆��E	�(�B�7�G�5Hځ=l��JtQ��N>y��X�������zw����cSR�H�o��Q���y�.�W�B�r)=#��lh#=��6�!������V��z.���^7']�
�$���68f��-6��5!@�:����Bq��\ٕ9�N;�[{�778��t3��T�	�ԫ�ZU��δ�0a�E ���)��z�)2��ݔi��t��������ص���;�5T-P�Xbf��x^-7��a��p�N��G)U�[��T)
�����L���T�1�*�ХJ3��em�����r�<���2N��c�0Mk���7�'{o����%��R��ð��`�үgS�%�U�� (l%/��qS��o���X3�l�3�-�{zѤD:7��.�ʛl�.N��tĵ�H�[��CN�5J1abquyN������܋x��}ScV�ٰem�2�,V�[:[s�9{��0��ݼ�́`�6�Tv��*�FDn���B1sU*�F����JkW�j��T-F�JTUP���^M�U5H,�44:�kZ4�3E��S)�J�Q�#C�ֵ��C)XS)��#UJ%U�aZ�kZњ��V�IUMR�T�j���Q���W�kF��!M"*(��)M%(�U)h��zֲhR)�))��J*�j�YUAHʪ*�B�UIMU$��j��(g���p��Ve��γT6�ٲ��m�r7>�
���Ad��W������������5�>������0�H�[e麹��#�%{��L8k�I6q�Ow��֦h�5/�\ꆧ���V�z���b��|jb�P�86w{zsb�{,>[|���v�!�����jKӝ���mE�;�D���pweo�6O���>Z�9��p�rՍ���*(hZ�aw �V�WY��Nz��y�sz�w����"��P�@Y'}�{��6���s������s��v���,6��Y�Sͅ�Uv#���3ѕ���H눎�<V�ZzXҴѶ5#ɗ���vy�)�����Y(1~Z���*|����G��<��}|���\tɥ��}��p?=�|�A���o��?u�ulKo��7Z8_{�yI���x�Z}���;4��l��9�i;�g4Е���_���]���߭(�R��w�q뼫x�gX��n���WJ��4N3{eC�8)������5�WLQ�#�Vg�.T���������0h#�"1�Y�}5A9��ǆ�n�;���	����]�vƪy5388�4U�>�����B��􁂧�/e-�]|m���n����b�0#s�������̾��[��E�X,2{U	J\ًa�ʰڑ�F9�?W�����s3��LL/{��(~�g�l���j���t{qG���7_���Bn� #Ub�fU����{�Y���r贰Ú�0?y��$~>w��/�o�����ٴ�>p�-�S��h����U���@|cΩ���S���gՑƤ���N���`����y��n��x�������p�RҀ�*C��(�e�w}�_y��<�;�ߔE�$�y^穐d����:�l���Μ��&(�v\v8������~�#='٣wрmf�nnM{�����x'XE��D�i�`o7���<K=�d�ؾ<߮:|��$j���$�[q^:.���5N��w,�>~�a�2~.��v�k�`�w+�C�ҩVz�H��J��_d1!��KCt�M�t�j;�I�_�_�EaE$R
B{������o>��9[S�Y9��u�3Ei�8Ʒ���S�߅{�7��I��#^�\?nX���� QkBc��έ�ˉ���v��v�wk'	�[�g�ȖP8�ޛ��h��2�w��P��M`����O���������/O,�l2Z��(;c�W=ˊ�|�8w�ӂ{�͕���=w������I̀���@�I�u�O���ֿTWW���ؤ���~�<�~~�S���.���g�7l:��Nģ���@�Ԩs1��Q�,��=Ga@}x�{�/k�Z�ա���7�K����)Z���2M���|�|�뵕ae=5&�Tt��T^�E��kH�7k/'���ߛ9K��sY9��l����Ra	��N��R�>MN���U��,�Y�(C�}���f�xa�]��ѧ(Zndr���_��̮�Id��/��ױ��
p�{�� O�(8���غ����{/+�rcr�Q)�8b�B���t8�N��ҟ�7����\d]{}Q8�@��*x|�:���E;o����b�8ܡ�\h��<�+��.�+~M��ه��w�b���bd�u�#��⪫��~�����,�����}{�����?%�Ll`��Fȋ�_��EB�m��b#@�~�r�)�+=~;��g�,]��hM���5g7�-֪}襁\>�=��&4b��9��Q�F��`r!8_H����y���)�\g����Yf��y~������?�r�kU���6�/�|Gg���Yc0��i�ʛ�KwҰ�(9�(F[S�2UW��~����ߔ�R , ���?���7�s�Ni�y�(������;(;��Mi����U�R%�������:�n�/���L轢�HK��6�d.<�+u�Ɛ*�_ya��^S������5e��=8����Do�:e��ל����)Xݝ)g=y:NTW�L���DA��~�ft��կβ����pM���֘w�d���ɷr��MBX��S|ldܦh+���i�Z[�ɺ$��G�=�a�ow��e��I;�8�]�dR	,�y-�퓚�܁�� �k����sf��ᴝ"6~\�e� Ȼ)�Ua/�0���f���Ѣ�ط��W8j���e�E4�q�����9ԬU��0=ņ,���ȕ��Y"ݞ��y(W���v�p��p�5RP K([
0ѣ(�={����r�S/���E�n�m��:����r΁�ڽ�I[��E��rl����;6��5���ݖ���2$�������i13A����A�8y��� �k�u-&��������p�P�>|cX�N��q���u�M�}2e�R�}�e�0�1�v!�����f�IjEǞV����n�ޕ����k�*o��k�ޕ��&���]���f�i��EH�J�-B��E`�UR���ތ���*ҥ4����L�RR�J�R�Zֵ&U�((���"�j��ֵ��H�T�R�(�b�H�Ƶ�k�cIE4��"U!C*�-���AZֵ�kUUEңt-%6ҷEF�YM�U5Q�kZֳ�5C@�"!T�5AWT�t��V-��4�ֵ�dӪj��V��USRꛠDm��j��lU����h�j:V�,�[�J�ꨶ��]QT-�t,��ƪ�l���u��T]U�Q�����[nz����K-�gV�,�c��,f�6��0h��)�{2�0ҕ;�w�C� �"�(,�IZ���pg����4��T�0��!B��B؞gw%�)����{�R�o��鷪��ĿxӴ�3�����_h$����ߛ ;���ꓗM/�<E_z����վPk��<1W��s�<V
��)�գ{�.���p_�{}{�bJ�*��j�P�S-��Y�\��aZjof"�g]F��V>������v$1�������,X��P=�{}����sX_�:��r'�pw����^;�����cr
���;�>�m�C�k�k��5�+�Q���k��,��`<����p1G�n�}z�p�P�T�����ŗp+.���-�"+1�����7�����w�/U��m/®dt��t��42�>Z4.���v�䒮lKBy�����s�w�s���b���n��=��ׇ ��V������[�KR���tE+n��lu^��u���r`^�g�77���nA��[�>h�MC�n�r��Ysh�בȡ�����3��-pd[cT�x-�[���\{�KכA��ҳ�޸8�SB����篷Vqa�s3+�<�(]�d�6�+]�&�������c�::�R��&O�Sr<q%���3���̶�e�#����Eep���J�w�H�q��c��o0q]�<3h�MƠe��xq��7���n}W&�����X��v^M7WU<]ٸ��=��F��Kt��}�'s�)���aߺm<�@{�;��cxt�aY��S�J�ɞ}��_�n��.L�bN{�� {�QESwc��2���[�(�r�O���j�h+�������y��k炩9�z�c���C��ߜ������k(�/0o�z��h�{ڽ��6!h�����FR��Μ�յ�yw�U�y.^������}_|(���X��2���ٻ�Ddf�H"�S�";�v�͙u���Z������~��ۄpY�oK1��"ˇ4��%��w&�-����d:n;�-:�VXiJ�G�UD�ߓ�z�Btc����o��X����1�q��&q6#�η�h�Mm֮������q���l�n�l�]*]�F���/���3���I��4���](�i21c�V�>����fg���<yOWN�Yx�؁��Kv���f�\f++������ꡫ7�;\X�/n]��ㄬ��S�� ��j�fFv8��Tp	���
��0b�5�'���َ�c�}O,��3�Z�;���/&L\y��	�� u���´�Wa� �~�����fH�vVz�I�@忋�N+��ꂯr.��@���x@Eo�ą[�1LO4~�_}��ۇ�኏oV��HO���� ���r��(����c�8ҭ�0�n�Ε� B�d������US��~��C�z��Ѭ�B�>t��]��s��_?!�^�y������䇅��/"O ��=8�5�=��5\����B�|��A�{�c_D6[�C/*ք���Ź;^�����81x���}%ȗ��o�Qy�����Ȥñf�,��o��v��ww@t�/�9�GY��\���m�i.^��X+d$3'�sg�(�^8�n�)�L`�¥���r�F��׮�����GuOB��,��h`T!yq�wA�r}���H�[:�� ��'��ۼ�k0���)�vr\>i+��� �e�+���.P�5�����M�ٽD㍥�i[>b�}}j8�W���Fߞ ��N�Z��]�1��_P0}}֩��-��r����#�n���x�R}UE�����ʺ�'�'�7���r�a�w�/�)��I�8A��r�[�5y�����#/��W�}>��`.0F9����dVL�9.���\���O*,�G���8o6]m���4Uxl�7�\�\{Z�f��[����nzp���j�������D��A��DC�V�Zub�X�6c��lfg�l�Ef�2�t7�a� �F�V��L"����C��F��܀�=��3�l̷G�f�5[�+�S%��7���%��-���;)v>5t�NZ�S�y��ڵj죄�^@�&�0Q�����|�T�m�Zm]�ٻ*Lt�wV���b*�ow"b�P޼���X].]�Z�]Ҥ��76���8�eIFPz�Ʋ"�%w�6*���k��Y���Ҳ��T�������W���n�j*T���5[� vz����ry\mu�挥��{ޭ���U;me�7r\����8$n���u�J���CԈ����#�q֢!q��%�w_
�3I'F���$B�}�Bf�&�S� `�f!:9rL7(<ț4���)�5f_pY{�����Ԕڐ� ���آ�&�YK]����YE���Sܕ�nU0���u�+Pu(��������ꀣ�
,.�Wwt�%(���AT�F�jkEH���*ƚ��]M�]B�F�I]��}.��MQE  AP4��� � ��݁a���D��$� A$�EP�>&]۰,�4Q]��R���V+*�����kZ֑WM�R�j�ں�*�*6�QmkZ�u���*����ij��.��)�UkZִ��]���2���P��K�Zֱ����)��)��]�m��R�Z]��TUQBSm"6�*���r��b#W����o�ַ��5��c��QY�OUPc.�~�38Nk3F�~�U�Y('Y�����6�g�e�",���n�ٱ�Wq���D�Y����ثp"H�y1��Z�+q�&sW����y�����z&K��4sV���D*0��oe_n�!�a���+��kw���5m��Z/!�ﺶߞ��հ������,�9�R��Wg'U��L2O����|A[��F��!��}̏��Ѓ���}�I��_�y��V�),�kA��W{�V�#-l�	��/��!�g���0�ӱ�S��+�nH�MڜP���/��&5���Z{�u/iڜ�����4'_ρ�9Xs+��3�]�����U-˺��瞨)޽����wW8�6/�6S�c�%����[���j�{y�<�����kN�x�Ϩe&���˿:x�����3��^��������NA��T�[J��VUOfp3d�<��*g��,u3�iQ%��
�\�]���=��9��),��2&��������^��.97�'"����Vs�H��!�ӆ!�̶{�3���E)1��=3����wQ,cV�:�P�6&L�A���m7�z��X�j6lt���uԷŠ���i�Df}�֏��h�5>���yΰnϘ�v��_�ȫ鮍�itX>��:ć{�Ⱦ<,�kos��8���?�Y4g��|��N�	��*�c�$=h��g��賲���M��6Du��/����W7��=#��Q�7���]�(����}���oe
�\M5�j\p�'�N{}pn�O��{u�.ǋ���<Y2:��y�� 0�x{z1~m��<i� Pݛ�zor&��0Q��Xk-��쟨o-����b?`g�uuH�<<fj�@��V��;�в��A�.���v���C��1����8��@�@1�6���X�^6��L�"Ȳ�|+���L��Ddr�/�7B:�|��\܉�+��=~��Oص�Ux��vm�sk�d?{��>W���;@�@G�_�d���H a��;��_�v��T�| �soY������x�=]� �'+�5`����C׎Qo�9Eu��zJ���HE0��Q� s��6�2�m7��F%h���6D�Z�V/5���Νx��R��Mn�U�܏qi�E-d���V�}�o?s �E�8��=��q�`d��7="M{l]��C�V��Ʒg��͖�����]�|��K۰���T��U���ذ��3�U�u5��Q�w�K�i_ywL�OF��5��k��)c�~�/بE�o�����]�_K��Έ�zZ�P=o���Ƚ�X��S�ʙK	�c��q������.�JR/�i���k������Y|��M&�A���YT�4)������}M���>}�/�=��@�Vh졯p��	\�t8?��_�w�^7���w�AL@����F	��^+��97�ͨ�%��B�b�\&6f��~^^�0lz/=Oǁ+�Aţ�m��(�@��Y�*��,(G�°^�hfV���t# yM��Ye����m��ZX��%f�wvvU��g�7c-��t��+�U���g���|��_�\X��b�me����v��zk^�ׄ�_X{�2vz���^��;$#;�Ն3)0y=i	"�z���_37��0]0<���8f^:�S��z
bi���f�u��J����b������t�%X���FH�c�f�ȴ�<��� LS��\��e���΂�W��̐�ߚpRoݫWZ!��3s.��>�3���z���~���,��>�s�AE�q<ܖ��,�3�җn�܎�eǞ��Ey�9�C|R�h>��^�կ^ܛ�E3����-����N�ya�$�^�^��)|o����Z�q�kV�8;�0�]V�p��NPhS5��/j2�#��=�ˋ��ٺ�,Z�}l���Qj��kN��7YW�S.s�փ�:�>���K�g%�"C����]�6��EUྻ��]nSCZ���N�f��²�
�s`� 2rwNyȤ�Z����qU�Q�o,�f�A�I�� ה#�]�r���
�5��_=X�Qm�]����-G�fЂ�t-n2y��v�=B6N�뚬���Vh�YH"�L�|�iD�vo��:nC?a��>�yu�R����^�0eo�_�1̜{M�7VƮ�\��;�(��X�ŢB���g�\���=���(��P�cI���й�+�Z��gNm�V��������I�u�Iz2�T��ŋ'7/�bdmaD*a�:J�0᝽�֖Q�#�e�w�:��Ȯ�F<2���i���h�ˤ��o�h�Y9
ᆳ1E��*X�R�Z��e�M��*���EmK.�c\��c3E�jUH�7v%40����j�ֵ��i�ؔT���H��7t�[Kzֵ�j�Em%�IH�(��ֵ��V�CWh�P�M!D�HM$Q	D�!]���I6hP�H�
�(�F�HU���j���-T,����[�����k�ݶ�UEj�.��[Zֵ��B�1��)�hj����Ⱬ�m�RUU�B��C����~��0��:�iܕ�{kE^l�V�1��ܡ�!���IY�5��V��|ڕܜ�<������;k�z������/�k'�[<��nߍ�e����"
�յ���55`�?i�+��=�rG��sތL���p���ۜ��*���1�g�3�3�����&�b��{c}~������[��g�3�/=zp/qU^�i��_x����v�K|$�^^��>lC=��zv�Н�wb���fd�u7#���|Ÿ��g*����ǉ장��O��̛'�X�s��(�Y��EÆ���ڇUj/5�b�#��D���o���c0z�2ȥ;^�mέ���p̺У^Lr�ZG^�|O��
59F��h�~�7����a�ŪG�ɓ���=������i`�����.��O���h%~G��u�t�W��C���f:6��F�4z�t�f���|�]轖��ү��v��21��=�|��΃?`�����P�������ݶ��I;8{�ϸ��O��N�:�3�w/v���s
H�c����9����N��HFb����u�k?{��\�驞��ц
��Ok���ŃI�Ǧq�,�o0�x
̳�ݽ-L���1�Ӭ�e���"�������r��\Ė+�.-?c�쁛3[�~�-�w����9���קB�"h
ܯ5����,�����G�F2��M�ͳ�Q<�Fx�
��$�ϼ��ݯzKV*�.#u`ͬ�|�������{���E�hܴHKt�p��X��i����wVeq��wV�n���e�؜�ރd�Ո�n.nLf:���D����	���`�vJy��Uon�v�=��r��	���M����s���To��³��N����Q� ��/��Z�lE^m�du�@w�C��y@�7uꅂ���t��W�g5��xY�Gp6l�K5�Y^�@E��XW�h�8<<���xoY���8�F.f�j_[�Eb��*ҙH�f�Id�<��.F�O�G�t��kˡ����;F���Z���20-J�C�Ϧ�yΣ_�.��b�&.~���G��M��z�zn�l��,ZXI��7�����V|��o�y��9�=C�zs�v��=t�R�L��`�����<�V�{;�aR<��}6GfA�4o����(�ysk��^hR��i&O؋r<q8�][M?T�}3�������}��}�~g@�K�[^֮���h�7�7�+
��o�5���?I��5� eЕc��ތ8�=o��R5���[�V��9�N5��h�1O���kǒ�l�4�l���ɭq_L�jw����[o�lQ�5t���{em��3E6��������ug�������#�o,țz�R&����t
�r`����v�Ի�˂5���6iQS��Tf*}9;��N��*2�wN��G���qᝂ28���ԣ+�l=}�z�`=��'
��Ps�Q�M�f�g�V9�(�z�K=fUuq~�{�O?ms��W�c 3���6�ރ�J� �@tBc�w.i�M0<F
���"Ng#��^Gw����$y�K�r?������W���B��JxșN���o�v�ų�����Y�c�]��=�MQ���C�6�c��զ�b���3�u9��u��j�L���XՕ���&�O5�0�x�-a�3�o�e<�MS&<�1��o�Bx=]�ќ���]nBs��k��T�����&i�.���Z�.m�a@�
��Q��H�DwVv�3@�Kv��skw �*.Ƈ!��I�����9�<݂�{��y]e��k���P�#�1h==�RD�������B�C��b��e��w��w�;޽z�۫P�\���G)�ܴ����8�e��ӡU�����b�k��r�Z9v���-1��_7(�^��>-tY��pp�47�_.	*t:��T� ��!5���#��GƦCV%��vh� �6�����y,�F�wXe"(`��yX����n��e��H��@)���WI�J֋]��u=�AV�Ƅ�zĩO6��	�kV-������(Z�O"��&fܟ,"+R!�ЏUݼw.�D�`��e���P���ޡI�Φ�ljAn�wu��FG~(�Ç�Oz�m�\Nʓ��"��<�����å�֬}:���L�7P�ͫ[-�8���55���(F!�{��X$�A�1�'+�uKˉ�s)������	��̷D��C[�6i�<TT��4��3���f+��Zӛj��R<'4n ��pk
s3��0�֮��9'e���&�R�}ε�Y�-e=T��Gn�vdB�V�պ�O�ѳ��o�1_ �UZ��)����<ֳ�m�.��Ij�tT��ֵ��B�5cR�J�kZִ-*5Wv��(�SE4Ƶ�k&GH�U�X�]We�%0kZ֮ ,���
D�$�+�W��	$+��kZѝJ(IESUJ�4��jS`�
��Ah�$ >D� �)QU@iU�kZ3��)���BT��[[m��m��TURP�TAQ[�������g�]Jp(��׮H�*Gݽ����5Ge�Dvv��U4Fϵ�M���t<���+�>�2��ZRޝ�~��S&�����J��FIc��s?>6��yw��,.u�F�Y�:��>g�zx>���������W�3=��"^�ێ/Vk}��go��17q����1�O�Y&�ɪ}N[[FK9::�P۶&J�E���m6N5�
�"b.�9נ���I�޶��$��.V�Ω�������,J�=�x�sGƺ���̓;^[�6�?�]�^�r�Ɔ��틾�*+,É�DK��	yj��v����H�M�񯗴/k�	���;��O4]�<
�<����������������(6&�Y��ѿ`+��ـ�դ�W���O�e�Q̱.ˉ���L��F�7�7;��9��x՝���Xǖc�QJ]")o�[q�g���*��;^��x�՜�/���^�Ï�@ww�o	�X.}樜��0mH�͋�֧��2�BM��_Ev!���P��-��@\z�ڥ��ZI���L���Z�zl��L���R�4��g�:ڃec�p��[&�
v;n�u��5ҹ�l�5����[Y]ME�VҚ�P�sB�v�V���q�8n��
��S��b4&����m���1ݓnf�׆#:#k0�2���ypM���!�9�uv���[���~i�ar�o�͍�v2u��ۊ^�����ú�7��%G���RF��w`�,��Z�%���%	J\}����eYmH���w��	�xq��������~x"F�q9B�����_y��G"G`*"�^��v�bP�]�yg�=�iz}^͌��ԵTI�V\���J�v�V7�T�H��c^Y��U����u+��\�L�&S����Ƚ�`��3q3~1Y���AK�'d�ӫ��5y�>O�.0��S��ݧ�?	~<�2��ӔOB�(�ͨ�q�e�W�]�;<�_f+ⳡ�^�\����]��-VW�t�](|�j�>�-c*$E����.���C�>&��
z[�M��f�����7��|0yo`5��L�$&��s={��������.)UGvAi�a���]�^����u��W[I���-�N����_KYtJ��;x`�|��P�6&��L��dW&�-g3�=~&'}f&��Gxߢp��o�k멕s{����^�;י�V|n&���&���檂6�/y�[;��:D�T!�c�y����+�ǯ�P�j����K��^�p���ۂ�)��p��}4:w^ۈ�#��y&�iƷz���c�����(s�!$��b���{yU���5���4�����b�P�Y"�(J�#i��2��.����<���=��
�n�1�^�6��r���g����V
F��}��s�$y[�z;=���1�x��qosZ�y���{��|h����^ӳ]F������c��a���V���dܩ���C_��������p�KqQ��v�����3�f2nO��V�+��Xټ�򤦷��G[�NA�Ve�|���9/r��c�Lj�l�f��q7��PÙ):C���g��:T��p������`��'���ɘK��+�x�t;ߺ��	�`��>�E����O	�O�8x_'���E�u��A�X��2f���sh��\�X&&��9�;���v���/s]���V������f"���3��+�������gi��p�Z̟���x⑴�f��w���R�(Mҙݠ��a����J�4�G�z��hU�NS���A����G3˒���i�cD�O��%�� �Nl�l��_���GZ�{�YP��.���]S��8i;�),�eErX�.����m	�7���;1�헶+�敾�����'^M�ڜSI�����
iPUS�D���K<��C��E��@�~�*�j���]bQf�K?��?�{2�FJ�oq���-�c�,9��R�TI{� ���-abKXY$���K�ZD���K,-$Z���T��cU��"@d!4,D��"H���eP��J�*0��@b
�@b " 1������ 0�J�@D�@� �@D��@A D 1 1� 1 ��#��%���H�8Ȱ��A3�C��JZ�P�I(�%IV�O�'�!g�jB$ �B)�7D�����s?����?��p���&��U�)fC'�t�s��Y�����~���CJ�aR��p(�a����kf��I@%K����GB�+T$�G�#_���:�u:�j���Y&�v�C�$�(^H�Q!��U!JE�\�'K��lz	��\t��Oɘ�+�c&�#�704���mx~��1�m� R�W�D�F��G�j�����RR�#[�"`h<�%��3q�Lr�P��m����$£����G��Z���>o�	�6Pؽ��j��ˋ��𢳷?ӿ$�RץW��t��X����V��3��mlV��:Z��4)�YI`� B��@@/�P�	1��[!!�]hTH�J�*\��~(�	Va����L�oz��-���le�@�m�a!�� �A$)B��	
*�qp���$���d�eM�����"ץK��햚a�p>��Ni�J�Z�����!g�a�0<�?��k��uF^Ω/6,�����v�aSJ��zD���#�C��ލ�كC���.]9���E�D��v-=]Ső��:�+8I��R҇�:#^��f��37�����ƃ��"D"�|$u
��:t�f�3hh�cAu)��[��Z$X��Ħ�i$"��������LEF��{h���Udp]^İ�`�G�ef�%�J	vH��2fل��p�RoaJ*���̌%�Y�Y%#Lj���HE�I1Xb�����3���R�}u(��������0'�	��3 ^%O�d�	��`����&�0YI!s�Wٳ����6"s�舑�t5��$�k�;��[7���������[��u�t'0�ڟ�a�# ���D�XXW��)���Y'[a���R<��$�x/���O���MI���ԴD�GC�8�e���KT����h�C�֩?�4���D�E�u�2v�4M,i����d~�a���O�t9�pN�pG�y3�#<��**3��x���^R�WT.��ޏ�eVF�F�\��C�լ�U)�4-3fʮn�{�^�>S�Rb�ˉLt�˲nZh���S�'(�FXڛ��|U��T���i�ъR3Q�e7��l���u��t䤺��4T�,�pib�$5�O7e';D%�c}$��D?�RG���"�˞F�	�N���8�M]*�����!�r;!�*L�a��]VL�ee��he���G������M�QO]�$t�����mnI6rL����"�(H	ʀ