BZh91AY&SY�W�ݝ߀`q���b� ����b@/�           7E=���0���ĩVͬ	U
�(�р��*!B�%R�UT( PJE
�*��UJ�QVf�m����T�os�)UUH:����Me@H�ĩ��E!����%[j����kUUP
��IJ��*�D�iJ�Qx j���`0�	$, Z�d	T��1IH��AUTB�S�	R��i�IT��T*�4�(+fF̤�SXF����j� 4 Ǥ� 
;��(�[lh��2���[�7Q�Jӹ�p��21@��\ iXe�@���x $aې�Ј���Є]�T�|�� <�+��<m׭�Ī+��N��@wnU�L�*P�t{���t�R��=���I[�.yTR�%�����l5}�*g�� �SA^�����.���
J5��jP�ET_y(� <�=�h�EQ@�/w�CJR������s�Wn�=��R]��q�R*r�=���<�=*�������PQ*W�<��*�Qs�;ʢ�T=�`���ћj�F�K��R �{���!绥(y��ުh4�=ޔ��*M�{ީJ�;��=P�
^�^��Ӕ�*:���)T����T�D���<*{]�v��ٌ(U*S`���� ���G�>�
�M���)R =�n�j�C#��J�&�%��*�����z�R�G��:�Iީ�;aI*��t�]4$]��uJ��QђH��u��RK�JJ ��|�*����J�EVh,�)U!�7׉B���8t�J�3�u�R�ܣ�R�PVtà*�M��*�Wm.:�� ���T�u�4��2���<y� h�����@� ίox (�� � h�L: ��vӀ #, �GR��F��B�}R��� F��B��1@ �t �`�t�t �+� 5ۜt �` ��� 8�EI
���m�bTQ��R {|  ��� ��� �  wr� :�;�� ����@���  v{���t[��  Ψ�/-R �ج�>�)@ c� �� 6����� j����V��;�@9������ �h�<|  JR�U %  S �JT��(i� �A��d�C����h�L ��4�	�L5<�%J��@     ��Bh�J�0  �  $�JB
�A���  !6�����M�<��hhhi��'��_��?O�q�a��\Ȼ��{��x�6h��rE�>�g��}�9�w�V�ϰ� ���
�" "��S�DPW�?`��,�����~��=T��( ���I$�~�H���H������A� s���w���Ƀ�X:b��LbS
`� �%�m�[ �!lb����m�l[b� �-�)��i�l[`�ضŶ!lBض�K�m�lB�6Ŷ!l�ضŶl[b��6Ŷ-�m�0-�Lb��-�-�[ضŶČb���m�[���m�l[`Ŷ-�m�[m,b� ��m�l[`��Sؔ��Ŧ�m�lb[�L[`�ض��-�m�[�����`Ŷ-�bS`�ضŶ�`� �-���i�l`�-�lalB��Ŷ-�-�[ضŶ1�-0b�ؖŶ%�m�l[`�2�6Ŷ�-�lK`��6�1-�l[b[ؖŶ%�m�l[b�c�����%�m�lb[�6�0-�lK`�ض��-�-�l�Kb��6Ķ�m�lb[6�[�6��-�m�l`�2��m�l`�ؖ���m�1�-0m�l[`��6Ŷ�l[`�ضĶ-�m�l��Ŷ-�m�lK`��6�`F-�-�lK`��6Ķ-�m�[�6Ķ�-�lKb��6Ķ�XĶ4��4Ķ-�m�lKb��6Ŧ�m�l`��6Ķ-���lBؖ��%�m�l`��6��[0m�l[`�ض��%�m�l#ضĶ-�m�lK`��lJ`�ض��-�m�l`�`��m�l[`�ض��-�ر�l؅�m�[ �c؅�m�[��l[`��-�[ �l��c-�[�-�m�[�lJ`�i���-�m��l`Ŷ-�b��`6���-�l`��6�1��-�[H��"�[`�[b�LP`lAm���P-���E� ��F�l�@��� ��@-�)lAm��
6�� �Fآ���`�[b#)l b [[`�[؂�V�"�[b1��Q� �� ��� �*��@��E�,b+lQm�-��
����[blm��b%�E�
6�آ�[`lm�-�E�
6�`lEi�-�E���Fب�[b+lm���m��`+lPblQm�-�E�"��V؊��"1�-�E�*6��*�[b�lQm�-��
F �Q�
6�Vؠ� � ��؀Sm��1�"��F؂�b�lm�-� -��U�m���Q� ��@-�-�Q���`��)�lDm���E�*��V؀ŌTm��1R؊� [`+lQm���U�(�U�(��[[`[[` [ثl[b�ض�b[����-�-�l`�2ض���m�l�6Ŷ�1m�lK`��%�m�l[e�#�6�-�lK`���)�Ŧ�m�[�6Ķ�m�l�`Ŷ�`Ķ��b[ضĶ�-�l`�ض�M�)�L[b��6���-�0-�L`�ض��l6���m�lb[�6�bF%�m�l`�ؖ���m�li��i�lb[�6��%�m�1�-1-�l`�ض���m��#ؖŶ%�m�l`��6�1��m�l`��6��%�cm%�m�lKb�ؖŶ%�m���-1-�O���Ԩ��?1�ϓ��J�+����1?�eY���y�&P[l"�VƎa(�w�sr�r��n�,büZ��X�.�P���t
��ŋc,�X6�����	��	�*���=�ޝ�l�%
p]D���Ūz��FL�h��*�8�-w�lB��r�EZmIF��b�&��)Y�A��4�
��b���mݣ��mӣ#������p7�&�&Gj�UYO//;6f�5��m�\�������Z�ʰ�L\��3V�n�ҀctR��BZT*�E@3Z{x%��Ks���w]g���<
�tL2!��Ri���9r��{�i�$'j�Z��w!0G(9/*�-դs@r6ɲd�㺭MH�RG��+ +j��qեux��M[�h�J��2ݧl�ڕ��f֊��l:6�JU��G	��0����d�%Ơ��L����6m��|�u��#XU�r��Y@Ӣ[Y��R��`e��x6��",Y�Ȑ����G2�l1��,�*�n"�j�%�̔�X��x\���'s%ov�h�j}��;�;D$�5 ���f5]����)�K^�	M��:I*��YX�(azc�'���yR`��݇c�dbEf��kl��nN��+*�w��\�$��̷����h%.�;��-`U�E̙�����74f�[�X�cV�
�7L.��RbA]8��YCX;����.�K�ј��ݶ�Tr�&������rɒ;wIދ43ɤ
�]�W��������$��lZ�^��J�
*;�1-����փ4�P�l��aLuxƈ	!J]I(m�X��6��ʩZ�h�n��1�3���x�˰��]��t��YU��=z"���4I���ͽ���"�F����טsh��X��T`����=j�g�ڣ/]�5Cpm�Z�R����6�ݚ1Q��vw3&d.�L�GCq�B�1��Ɲ�t+�b�v�^P.k��7Ѵ�&�31�wEL��J8 uc^H�4�HҞn����D<�Ɲl�ɀ�=�*����jd�[��-�P��H���%���,�b��օv1���R	zM���W|tWY�1���Z��W�^��[��CJT�L8�*	5G�f�)�� w����A��n�����1�i*p�g\���f9
gڛ�J	�y�yu(����mHVfܨ2�$�i�Ze��Kd�������M��.��,�bܢ�Sb�]D/��;vӮ<��9nʂ��J�;��
(�km�I�����a���`$��m����=�d�;���1\E�G3&$D�a�V�0v`CTW���@��A�A$��Z9��+3�U����C��dwM�WO�4 jI��'�L��t�1,h�ͼm9��L�Fͺt�$>��hE&���"FM��)�He�`��4��uCFDTjã�X9.-E04/�e�ٛ{���v'Q[*yR���d��Qi�w@�-��Pz^��sY�+lỂ&F�h�Yln���l�l�^;�ܫf��8��-�����Չn�Ja[B@�k6���A=aI���qVL7����JEV��7fR�d�in�Z�ue��B���Mi�.��I$ä�Id�x���׭��.���J2��"�J�1��pm;.m4#r��͑m�z��h���7�ˢA]v���Ɂ�R��J�m�c�`F����`�Y�2���C��L���[&���.e�{u&,��+T�t�X҃�2R�:d��:��/Dn�=5�TJ���+
��M��a`f��{)(�,	y��[��QX�0�T�9-��D�1=Y-3����`=�2�0S���ů3.��D��U�d7*n�(f�*�-��z�aZ���l�X6#�����Z.��N��:ځ=p���Bn��im8��@jz;*���u��0�/沨��j�r��f͇D6-�ZZ��T0���F�b7�l�.�U劑H��쒉ʻ����=6�&$�ff��W�a̻���͡��,Z�L�J ��t��V����3D��mͭX�m���݋�-��i6��v�^���$�����u#��5�%��b�s�ѪVKE`m��k)Is/.͖f=M��ej�7"��Q�7��ݬ���� �IMfJ������R���-�Ю�Ť	��Z��3<���m N<�6�)�\�ʴPNm�jUh�2�B����#�M;l�Gse��n�:�
7�[+j��\��%35�bݘh���.�r�q�H��(&�m�%qEUK���o5J���$$FX���ef$)��V,�)��4k �GX��A@�Ġ�\����fŶu(�9�d6�|��S(���.���n5y�q�	�Fo;N3n`�o�8��+���h=@KY���`*�j�o0�BY@Elར]�,u��o�����Xe�������L�3��%�Ƞ��I ��$$��l���MB�0�W�vC���!���1����m��]e%��=��p�{I�`V'0nM�
D#�S�X�oX������I�hhY��h@�ɪ��-�o�r�������lK�ܫ��,f,��F�Խ(S�CC�:ݢD��K�(�U܆&��؞���2�^I(ʸ��i�خ�@�2�晪MY���
n^7�.U�1Z�G08�
�Y���A�m��*��5�����a����j��52��I�^ƪ��Z*Βڼ���4%�.�ƞ�]`�}�-���ڹr՚y�T�JV���z�L0 9��K�̪"M���XV���,C1�،�JΩ��QT�v�L$ɱ��sn��Ԛśe�w��$�E�K)�I�=)cZ�ʽ�T��̩�JieZ�5#2P�)�f�(j�7��U�Y���F�e�e�����V�*fܪ����+�������+dw�j<�ӞR���4ٸuD�7b�Ѹu�hl�6Gfb;�]
��66�RT��۶)��M:A"f]*�xA�p�t�[I��).ck�Z��6J�f"@ʹ�j�<E���R�5,��v��i�Ic����"�V�J�D�Œ��I��9B���r]'yr�^Y�X� ���ӱ�z�Ywו5�4A9��4�
�+/`��	�ٸ������ZV��]�J��e;v�R�(���3��Eu���,l�k$a�/p�%�̒�GO�\ݻ�Y�onushz��{I�5$�ֽ6˻%��5����{W��ǓE�" ��B��i� Z��f�%�s&�X�'(���D����hXˆlB��6A�a�݈�1�&V��P�ҳ�$`��$��q��-�O&�U��c��]cwB��Le<!
ƃ�[�-r�V�
�ఓ���4��2LW*�#n�"靫��k��b�6��c�2���3��Z�c*R���ӫ��>X���J��@���8\�Z-���ٚ�P7f�y���l��حєee]�Wf�CcZ�a$��v�Y�$�q�y������I]�ձ�az	�'f��'R�ӉEZ�8i��A�(ث�����Ӌ]��K����1�S�v�7tmZ3)�*ht���z�A� �1�9�-��)i�+ ˀ�;Y	Ѝ �S���h<���l0�B����Jp`�r���p��#�X�T�dY�A'c.�FPEP2ݝú�T���������A��i[wdU�������r�:�GnLnLڣ��E[�!���%�cnS��KG4���75��U���N�+@,Jh4ɹR�љ�n�!��0�C"� �-%D��a$t�ɖ��VΧ���r��XW���-ևIn�0������n�5�N!5T�,��QI����-��v$I���CX�l�5�h��.'�%`J6�D�u/��N��$�Z��y#�mU�)D˹Mm;uK���S$x�s0�Ǣ�Ѽڻx^��M���-���Z �kSz�F��B񂮉�A{j�G0�sJX�3,[6����YE��U��i%��Di�������Wr!���^��y%%*+�&b�C�F����K�x��+h]��)�V���n�}m�ˬ�G���.Pf��X�0�ޭpV��R:z/N�P���l��l50<�ڙ"�\%��v$V���-��t��0N�w�ˢR�On�Ve�^R�mǹ3wm��: �F��yY�0ąȲU�ne�p\D��^f��UD���
��{1j��@ec�a��R�K�R�k�V^#O,���oƂ�q$���.�+D�Q#@̌�kU��e$���R�RFȽ��-���'���U뵹���](�V5���MnQM�ۨ������j��E��:���Rr��!^$ ��#M=d�5yW$$</qdX�6�J�ʃn�!�8���%u��Zb�26����:'�p7{b�-M*tU���e��9r�w�u�0!$���ԛW X�QX,m��iW2�A��#x^͖-�����.Kڰh-lïA.V������dS�ν>Aҫ[�Hʹ��i���B��E�.��-eն5���ʆQ�Jz7Y�SV+XC �P�#÷I+��V����Y,.nZ"d]�u�4�C^���J�Zb�r*�W��ۆ4-���2A���MM+�Wv��t�;���QY�	����F�Q���꧄�5`ɕ�[�m�%�[w��ٳ���n�����Fŗ5�$�b� V�1�SI@X���F.\;#�wb���M���5ޫsI!�t���AɅ&�͒%Z���t,��F�;ub��/t�˹��j�#�t���I�:̇�����;���6ZǦ���^C�UEz4Hr,,fX��9��7K$�nc��%1�mK�m�5n�lY�˥^<hՠ�1��-PJŵ��R^ފx��-��h���jl)&Ŧ�I;8-��Z����"#��k�F;�2�`���b^�D2�Z�td:�M:�噀l1⥔Ҋ�8����FJ��OXۙD,�s�Z�f�'�;IF[�+5���Nk6KSD%5�Qz�4�l�J�S&�F�ki�FM����
��7 �ͱ�Y5Ś
ҕZ�FYf�.���Y�l�%� 4�,��U�!���J(�#U�4i���h�R,��\�-�-nQ��H�M�x���[��eг!P�W��b̽���¤��x���=����-�Vf��fl�;����uV��&�a��)!%���C7,�ݲ��R]K�	{-��+-8M�=U�3j��o2J����hU�˿a�wYSf�ӡ@��vW�aM���n�*���u�f�O+f+����	�	����a�n�RSi+��i�s��[�6-P1Z��u� � �� h�E����b�b���x�q�)a�2U�\��gK�w�iZ�M9m���4���=S#s.��$Nm4\�z���8.��5�-7��5[��
�u�4f�0;�B�3�}��%�ep�(�w196��0�Q�*�U��<۔��,Ȍci��̺�fe�R�;�r9+S�E���l�>�r�[�[te>���������y�,���e�͛E��F���b�n��n�+)0A�d�E��䈷��pYJ��wXQe���1��I<��+wOY���w��(�V��%Kk��R�J���{{t��GJ�6m�� XCi?7��y�R�]C�t���l�^��z-�+E�ܡr^+w��n���$�i�G��K�$K�H��^�8���V�ڲ�9�ا-5�*���8�´�Kk$�������k�a1/)���z�ax�L*9� �F�u2�V#HF�yGaY~����-e�`��z�q,�F�; �+e吱�љ�jř1P�抰��{��^n� �~�+6�_$�ʵF��մ��N�� i��<�&Y@�s�ˉ���iY�ru�rr����i����Q��\�!md�Q���q���,Du�\O���JDڜOWv�Ws�Ű�,�-%���P���'���d�Y�[*��d��g4�Q0�(��WU�s\�R-.Nшҍ8�I��8�!Lvf�8�1�B���m5��Ճ�O���KU�m+��jZqcN%J�4�-���W$qu��ܷ}�-cI��ch�Jj�Q_$��Y6v��	̓��:��P<oK7���,�E	�x�+�3֡�d��oOqM]���*X��"�N*��Q��4⴪%��z�Eއ����*Y�4�$�7g���q:a7�C('fWp��1):F��M��tSD���s�[D��n��,�2��h����'	�p�6�F�F�RPVO~/&��q��G�:z'Y���Н"�Ҩ:R��7�cĞ�i5�dR�V�wJa�qR9�ߏ�C8J��7�Y�A=�E��
U����Y�Z�N��c%�Ӵ>��@qLΚzG�N�q�!{@%v#j���kU�\��4yg+D�I��9���6L'�n�F��%Nz���gt�^��fNm��F�/��Y�a"GQ1��Dޙ�YqB���B;�o�Q�����m>Y��(�bXNO��d�D�*ɳ:p�'��ge�l�K9�p�"I�L���0�&���eq�qdY�c!	�54�&֤�����v���O(
��(�9d�6t�����ΫvL(��8�I%�I&�&F���L;ţ����ݮ�`ϨkqMOV|�'J�L-��d�a�t�gY6OKd����Q���⤜KTъ�*��8�,�rM����N%���P���)W&���MKbiSU�ZT�T��J�9�9�]i�|���V�T�DڍLW��QsM�ֵ5rRՂb:��kq=J�kQ�N�'��ɠ!��1�	�x�'5Zۺڠf5P�iJ[��x�$�NrѬ':�][ p��of)a�:e���J���C�o4؎;k��j�VJyݒ�Z�s��Q9�Oi�'�Jj�i�j�cT�)\DI$ykO�iL�Y����S���.�}���w��������}�<���}�'�/7<Mř�Xژ)t�<����:k�|��c����/Vʏ5Jb�0�n��n��I&��ҡ6]ڙOA�୫�i�Q���R��a2�{׺s�;��SCr�9�R"����Ylp��KE�{��\^�	�rQ�姧U�%��ݬД�Bר�l*"Wgo��	k���˲)&uh�ս�\�
;ץ-w��ֆ���F��Gy#o�A3���e`�7�E��,�b.�YNcԮ���$�o��ѡ�=u�L��}��{��R�c�����wJۤ�3{8����&��o���)Xή�(fr�+<�H��'g����.��Gv�3ss���b�|���Ŋ=��r$�u��kz�$ }�U4���ΎJ���:\�R��/R��n���s"	�zi͝�{��u�b��(�tL`$V��dsĳ8��z���_X�C/�Q�Q{[3�����&���)}%ul��+qE���ڽ}֐�U@���G�q����Y���Ў;ҕ'�w�(�Y��Qצu���E4�9p����\��8�-������;�<U;�N�Z�8�B���$���Ͱ]�=�kqr����{��(;��]��\K�P��	�Y��`��S$��I�E���i�b)Rv=˧���~<��ø��b&�fc��1ܔY�%��o;�],,m��ۗS���H�C#{B��3I�:3a��$uI��Ս1�oG"�\wӘ��ޛ��v�2o�pq�ƌ�mo@��{OQ6-b����4G'bV/���ӕ���mf,��}���\è�$������-j \��Zp<3QB���/z�Rw�I����j[�3���fE+��KĄ��;	�k�v�7�j�O��g�\�&`wBf�+��M�0�Z\hW�r�)G,�;}c{���x�B�}}�3��ܥ3�|���g�;ݹ�Clk}���z��tu&8;�O��a<5-T����EhS��<g/e�W�|��V��u����ʛN �.	[f��� �\q��\�3�²ĭ�#̷�9�7"�*Ֆ�8�9���ga�2;ߧ������w[��p�s6Z�8(T13�W������8��k����B��������d<����4����c�×��|�\66��$`�o,���l<���ɷ�nѮoe�Tę����dyoqЫ�=/-3p7��:LrJ���n�۰�ڸ��2WRG�}b���A���5�n�f�yv�p�8����Ky�C;{��+���	�_f�k��{gWKp>��Im��R�+��0�ε5K0�]�kq��r�̨'d7�52���y�#�7�w%`��o�G��!zV�f�x�[���M����d��]w�O������nHu��F�"�J�[3$�79���-�N��b\��6�Ab�83��),�.��{Y[8ػ�\[�A�oxZ�}ڔ۶������"�Ј�īe�����|�1M]y7��z%u��aQ����$�9K���p��W=����,�����w[�G�a�^����R�FR�%!�,T�������.�|FΖ���Xb<.�l:����!l,�fG��C,�9�y\�����
CnI�;awg��|J,����o�ܗ8����m�k�AN��Ѕ�V���Պ���}��E�%!Ǟ�Bk�� �^�ȝ�@�bM|y-�U=�]ǩ�e;�I�<7V�s*��b౳��怮E�u�:�/n�G��^�:�y�"�o�(ǯ^�u��+�[L�cu�}��C���w.����"���DG��V�N��Moq�p�[|EQ��rfwE�-�����:䃆n'��!iq���9�Y+gU�=q�R����#Y��έӭ�����i\=)�#��7f��Q씯{��sRu�-B��A�WJ�1p>��Ɓ'\�����	�\���j��WE�2h��	Vܐ95�SkV+�w���$g�z��Shև]:�)���冦9\%��/0�\�Xf��ɫU!�guӁ<�l�i�]]@n�ֆ2�[l�Be�l��j�P�|#�$�݉Q0���^�R�j��=��3����[G)��h݋��ȫ������u{�;�t�ۇ;�Y��k�QW3�e+6��vZ�.	��=���ʧ�Rׅ���4g9�(TVFm��y����nLw�FA@ѳ1�`w�m9��wY�_dVEk��;���z��D�m���Y��Q��m��I�n��N�;s]�xoYǲ��-�tG���vgV���T�K-3���ې�JWm෬F���}��.�L�!OH�!
.�F����MgW|��v
Mm���=4�)V�ۗ�ҁr�7�(gX���T	��!��i����!�wV>	�{���t�2��1��Le��`���zi�����*V���\���+�t��w���e�Ī�ٻA�݋�h�%�L�����9�R�M�#��HUէ�5�f��Ӌq���5"=K��v�R���գ���y
\Gv�^���Vs�]���{�PhN&�h���W1v�<v��вE���Ἐ�Mޖ���`˻���Qrl��E�&Վ�wv�c�!Х����L=�F$j�p�<3���lL�.���U��tov��W�|9���Ȥn�w4e]��_��.��&؄��sA��J�r�m���U�:U�ĎJ�B��Y�*�q��R��Γ��^�G1i���������W	��K�2����L�y��U:sԨ����ӵ3u�pY�r��-kU��j根��0j峼q�[�v�&ҬJg��@�!nm�>�6%]���1S�v
6/"p��^Qu�$K9��n�oo(D�fu���{V���ڌ�>���}T;.�4�FTz7:w�cs����n��*һS3������JZڑ��o:C���B�ef��u����}<(�]x�HH#b��暹3V<�V��t����1^��.�lgl�N�o!U�K�0/���k8�y�sv�a���G�p$�ehb����\L�8g9:��jV��`Ƕս�MrI�98]źv������gd�C��jŃrl����~	�X�ǋgK��v`w3ze���!�0���8�^��=M�m{�+-�r��
��S[S]�T��w%51�C�_7��.��n�/oFX�s*�e��zDa騕����i�X��f�F�Q\P1��HoN)��vW;���5�z�{�.o *���W;��+�������K���թ�놭�Ӓ������v�Pv��=�o�i)��tU�T��_��ʛ�B�.ýw�����u ��/a��u9"��ؔь.�kMr�ZD��2�&�Rfa!W_7�gf��H�_Y���BsgX�]�:J/�o�kwE�\�`�ʼ�=��y�8r��rɉE\�P(QY�]���e.=
P<�sQ�;;�D&U��4�H`����|���՗�cj�ERvK��(B�܄�טvڙ�p��|6��{Yuj%��z��P몃�fLޡͫ������|�J]�Ǹ��\"*3yV�T�_/qM��)!}r���5�=�n���N�Cd��%d
��c:v�Rb;���U���x{{�녷ϒ�5��z^w	Ÿ�'#ܻ�*�D�X:kk���2p���R�h�U�������m9��m��h�\��5P��m�3oE;!�:�<1�-	��6tY���\�ӓ���7q�/39�cй�u[8q�ce��o�|��n�5�x[o�����V�w���VV����qGU	@-�R^��H:1�&Og^�tyAY��nA[{���2�3qs����6FP�][�7	|K5YW��\�Y��t���K�k��b�b�Y)�Bg%н���zv#�M���]�Sz]wU���t���]hjb�sny�VyXd�JV�-)6�ft7���m��a�cڶ�΀�XI���k4K����j���St��+'S,j�cn��ת�^�ח,��ݥ�9-U���������:������e!|�
����+Mڛ�`���H�W(�]Jk&������������G+��J^���7�ԛR�_���*�I%q-�^\s��#\9��/������JO���҃���^���s�Yګ�6�Ԭ���ۿc�Hs��օr�\��{ͼ���:��!�uIe��������T�nelT���q��v��έ�]��(=��gK�6�"�0�V�\�^N�WjF-�0�o�v�6�+7Pl�_gK��j���1b����3�4Sx�)(�n�������꽔A}�9a�m��޽�t���J7��Yw
Ԅ�/i,�������P�6�iX\(V)�D��9.�Ȫ�t�#�t��s@����aE�{&u���/�+K��sU]Ҡw��sc�%���C�*M�)
�MqJ���Z"*��ڸ�ٺՓ���t��t��WJ���+��������/���p�A��.���Զ�E���\$oyv���ܭW�(��ג��W�Z�3j�<��;��i�hkVI�H-=��RKk*E���Ӑ�+zcw�u�hWg&�)��	�$�]ه�,�/T����0�����=�]X/t>;����]x�)n28&yn�h�KD�Kc���32ڱ32�:N��*�Yw���zP��9��Ez(��e�k�:#�o����N͕^&k:�c���AA�l�J�N�C-mr�)���m�ƌ�w2�KdNX���e��J_K�i�]*]v��
d�j���܍20e�7��
�J�R#o%�2���.��G5N�m�lͺ|���0y��X�4��w
�;* }%��F>�p���Ԗ��ͽ�VR]l`�G��z�rL���!�]��[Y:��Z��]��5N��8óA�/W,C/�m���1i�{7���-���}�kgs\����5��Rs�S��W`�e�W7���+5��\�ӧV�&8�ݚ��v����b�a��kj��Jƥ:����J�sJCc��r��+���7m�aޞ��B�zotpn�ñ.��f�j͆�7Z٢�-���Kn��Q���Zdt�7�;A�Oӝ��i�@�+:�'����Y����1v�u^U�9;�Xj�u+{�,f��ث��m���������;;�����M��]n	���sK:��ݻ��ڷ�)5oy�u�#��0L��[=}E���\��eQ�_ؖ���l�w/&=�&V]��W\U)�z5`��d]���K�L�*�*JR�E��:�vc��R���iw�`y���ky�ݼ�����Rit�0��w
]PN�i�E���Χa�bK�Sr���"�0��]��jX{�λ骦e>�]	j]s��c�bM����ojIn�8�N>�rv<�,�L_oh����N����z9w�&�������̙u(!�]�f�S6��3#Gq�9��\�8�i�N���#�~a�^^�]�YB��v4K�ԝ�UqU���_P�\]/#��s6 u�'&�����W)�S�3ja�`���Vt�W����%}}׍�DЮ���8��m�8;��k�"�V+��2�و�*�}�5l�(H:!η&��f���ۮ�w���&lbC�ź����|�Qނ���{�xz����,��j.��u;���Iۙ���ҵm��:�S��1��/Ը�BYp]�%i�+�1oma�Km7�[M�gS��NV��L橣���w��t9�k;���I7���GiJ�;-��f.��I7[@��5&�6�9`S{B]"q��&�M)�{�kOD��^_��4h��o��������K���X%ֻd�"<�ʑ�Ky<����H�t'�<��]���]�oIJ�6L�gz���>�;	dv�;�
侩��Dܾ��%��Wu�{�ְ����g�9���m��s�k���<��gr$����J�����

�۬�s�2��y��I�ȥ����<��Wt+��U�ɐ̫�=�� �������Y���n���y*�G�VD9��*�����u;�� ����� �{wa��yR#��.��S^�2y~K�ג�2 r��9�큳�Cw<ޝ�st��>y)G��y$ 7�E�4G^W�W=�����)�_)��y9��y�*�:h�z�&�~�"����5h��Zv*\@�����T�g#q
���TO`M�����"�j�<�y�T�	����컯9B���L��v(��W��ݤAP�}�����p�_q���?����Ϸ��7�j����&&Z,�I�ʨ!kl�ћ��n�L r+���K+�]X�]=�iߘ��X��Ir���9Z�iѺ��)�r���8ݜi��:�����W��C��aL�=�c{�M}����Z���kܱL�ײ��"����Ӷ�#(ʐG̨�eS����z-���]Է�K��j M�s�g��T�<wSz�b�s#P��x{0���T���ޢsnWP��rt�B��h�q(+���(m���7z�NM'�)�=j�FL�Tk��eT}h��s)�C���_�-n�V�Ȟ�݊���5um��,<�^�wʷv�eA�o_>{��`;u(�ϰ�����"ә]%�\�z�.h��p+�Y���w:Tnn�HP�Y�Ư�K%�k*}x�:n�-#� ;X!I)�S1Y足z�N�;�<2�Eέ�tZ�I�@��fi3�������W���S�*�&�y17�	k�v�([{��oߺv19Qu�{Ԩt�����;.������)��K��E���˫闁���z�#�@�Z�$\z�
�P�|ܼc���ͪ�� ���v㡶9�p��𻚍p�u�U=P�b�fm�׭Dm�/����y�ImG�����3&v�2�$�Z:^Mx+��<�6��_�����;z�:q�qӎ8��qƜq��>88�\q�z�q�q�z�q�q�q�q�q��i�q���:q�q�8㍸�8�q��q�qێ8��qƜqǎ8�X�c�8�q�q�z��8�8�8�8�:z�۷n;q�q�qǎ8�N8�8�ノ8�8�88�8�>8�N8�8㏎8ӎ8�8��:����$���I���W���3�v�۱,�"�CC�
5���5���e!X��)Y��f]��:����bnJ�-
�Z�!�m�1�y��[��ڻ�l����f>�-�&����eU��`�LVS|+�48ڰ��w�e��J�)@���m���:��W�J�ܠr�*�r�$��F1�\A��B��f�D	Ni��Pe[���ȡ�;(K�+��օwyp����s��yu*�q��XV
�R�rBM���f���yp���Nk=��+�m�N��DYwY�C[���[�2-9؆�pd������9�"EŽ�*,��,S���y�T�����a���rpQ�R�����u8e`����v���b4��!���&硕�w�sR9Af[�AB�fS<�b�'u��49;�x/d��j�.-	WmQ��5C��7*�^�D�(MC,#pi���XF�_t�]����9�$dVQN:y�^3j�U�C�޷����d�B���b��R�m�"��w�8�E����h>��i�mз�"uIY���t^j��2�т��tM��c�IN��z�H[�Z��E�y_b���/i*��t"�Yj��hQo:0j�4��3�>�Jc��[ٿ��t�����\z�q�q�q�q�v�8��q�q�x�q�q�z�pq�q���q�q��8�8�8ノ8�8�88�8�8ノ8�8�\c�8㎜q�v�q�Ɯq�q�v�8��q�N8�;q�m�q�:t��o�8�8�q��q�t�8�q��q�qノ4�8�>8�q�q���q�q��g����<sJ�L>���A�sRh��mp��)u�Zȝ��f��kE铲�7R��<H7Y"ٓ:�
R4�;������+Y��-V�05-6��ൺ��;�����xT�P*}�>�u�1E�ѳ�ӳx5��qVM����-�8|t��쓌�v���[�WB�\�N�U�ڣ9!%���NW@����m��r7]��td{�nW+�!��u�{��f�21V
w���4f��&�%�!�۩�V�=�Xw5���wU���a.�w}���f�I�,`s�2�2V�0YA��f�yL�-���À���VY��N���#aɆCX\�W{���۳�V�8ˠ�+�}ޤ^G{$��Y6���h�@��ȧ���N���H�3wX]��>J7�]\m_sL��(�2�W{�hV�T���}}����x�6���0d���::��ڭ�d�����z��d�3���5:�/�8d�Gj���۹49�ubZy^d�����9E`�7�7E���w��R|�b���̬��9@�h�6�A=<�9�S���۹�.��f�鵃r��TaX�rT';�eU<�X�mA9��d�c[�vX��F��8>M�#�[6��jnU��e}'{�;)��v��Ǯ>8��c�8�8��q�q���q�q�8ێ8�;q�t�8��q�8�8��q�n8㍸�8��q�8�8���q�q�x�4�8�>88�8�q��qƚi�q�q�z�q�q�q�q�q�8�ۧN��8�8�8ノ8�8��4�8�<q�q�q�n8㎜q�t�8�q�8�x���۽��m;��ڲk��m��;t��j�G3���}�.eڋF�V�1���k9�y%��᳷W��C,X��TO��[O0��PCe�S�Sժb��F���/{���2�T��k�^h��3���J4�j�]�%`݋�.X<qA��
�z��㈇̓]J�X�ܨ�<_$kI�q���5̃��o�/��2��R��']��f��X��:�rL��E�xQQvW�%#˖�l$ Z���Kʻ���H���}�Fή���3��^�=��w��u�9�I}Z��2� m+V�ѣC�x�ڵx=�I��b���CtV�UN���{��`�ˮ�sBv*\^�������LSx�]�L��]yt%�v[�����`Ѫ�ڌ�&�����U!ǯ��1��(���xvkvD���ʌf��C��\�I�wwJ��vP�w]�S�i�)�����K�=:���)_e���T��IϨ�%m,�f"@���]kT��w�w�y��l��h9t�n6�h-�^���u�!YJ�������5y)*O��+k^�%�Zܺ�c��(���6�n��K-CF��g��4`�Rj�ެK'{��u���ƨ�����*��K:�o��Li��{����P�Z�8��q�F-���®�y��c	|�jG�7]>͈;�P�9��/ �
tf��[�!��c�]G[���e5d�
4���*�m�*�:WR�)��[�6�{�nMB�0�M��v�m�r��J�s.�Zlɴ�Ai4�*�f,������]�Ɏw��B�db�mN�k&�R��])��r����z��F�#S�wpȎt"�7X�͛=�]��\� �A���/8���b7%ͼ���3��J�/;�K������)qoZnԻI:��T'E���й���`ۀ���hV@Ƅ�T9mJ.۶���Ej<�����*�8f���԰󡣯P$x%+9/<M��+7N�;u��K@y�j��j�͂Єu�<�|!�Z��+��$�yݗ0�V�Lx�^��!y�ao��������h[���1���5w�hق���I}Ւ�d��w�fO.ŁM�1ֶr�*a�|�u��w�%e��}��l�ر+�*]����N�\e[���e]��u��F������X��v�V�B��D�P�Oz�&;6��Jn��{�G��B0�]޻��p�<C������iC��*db����d:+�K�~����"���`�]����d@{2����G���֧
���h�om�K! ��%�Ͳj���jא���x�;&1h�}���hfw�⤙�yz��p���VU;x�̡O2:��;��ڊ�î�WN�=[�6򨫃�G+��1�)-��++�u�5�+���b�Û��V����/���#�4}������nM����.rsa�ю�Jʹ�vw�]��u����kX\�\�*Zf�V	D���-�p�{²�Tq�^�%6�z��W:�][�nH�N�r��+�^���H_*b��'������u��n�l(�v]:1bS�yAY���uR�W$�M�X��.���zj�����=��󺊧\kuɜ�!�2F�jS�Ɏ_�lƚ��8����f�u�}�JZ5����#U��VMLO�n9K�۱F��dX"�;(Ll��,�ZH[�\���ǱZίyÓ���sr�gf�/�r<�=q	�^���V��.b�aR�'�޸��b�8�������$����q��Z���<1b��|j�6��c�Ŏf�d��~.Ȃ ӭ���
����!��yH�C:�����}�ž�Od�s��4鼲�߽�w�(ή.���'^NM���mp�'N���	��l��у[�xe�gܙ�ht�D���t4&�A/zL�餙0��˭fkLҦz����2�Ӝ� Z�bm�xc�8�rm�\<=�\���t�ixv��Fڊg,tx;kx�	@��Օ�J�t��A��ڸ7 �^|u8ܨff��_Ӷ���S+��-�Ok���A��격@�����m�J�7f���c_�k7ݖ�'E�en@�g�{l�����5W=�i]+�I,��j�轚��K��+�������.��6��அ��Է�ǁJ��������ڥ[J-�`X�EUVCKE޴nM΍D��M�1"�khfS�}�f�V�{�(��T�ʄEԣ�Sd^�p�}z��FS�6q�������B��N�������NDo�ou�ȎոY !�],���(�$�վ�ڲ��[�SׅAx�S�\]��	Yyx��PUWt���ד���(K�$]O&��&�oY�pH6��[�����uj�֧y����OR,�&��ۣ�η��������J�o[��6�;Z/`ᷕ�΃W��7M��?fNX��q�|������2��%��dMҾf�3 E�\Z8-ħ�}�V���7�������ϩ��k6��K�L�۝�/E��oM����%x�VBH�TjA:��++۷a.��t���(mޛ���}x��XIH���N�9֥�zc _>��71|r����,Ȟ�쫥�`��u�YId�'O�_$$ �t��D}�WfGG�_K7;�FC;g����J�oS�]��oz �U6ծ����ix͆���o;:&�犽�)�׫�TV�r} "����g%��p�㏦�7�ȼSZ�X�c�u��\�h���-+�'
s��uy���ҳ���z{�h�����G7DΗ^�D=�Ӟ��9R�yP4�Ѫp���lh����Y�����#7fu��O2U�$%�5z�M���1^��_@�V���>�zZ��:L�SQ���Hp�{2�P�wx����dJ�$0N�EhV�*J���Va�Һ��Ks����;�����q�S�P���gn�C{�1�<�n	�{N^�ݢh-����5X2oi��7	p���� �^��&��j�6{f�n_�Nuq	1n�FgUZ`Cm��k�ʠ�_��"�Њ��rL{�٫m���(Gn�5�U���F9q�,�7�2E��ut�T.�4o�%��.�抺�L���]օ�-���eYS%������U,�fu�:(x-��(�kg=���["��$�������r�%�E����]�{նj��H;Kb9٪�/�d��C�SM&�䫎���:kLv6�l��m���t���KѼ�x�����K��x�֨��Ys�d������Y�HL7;n���g��.���^]��5-H.��|��)emT��r�]�[u�U쇕v:�Am�C8y1ܭ�N)ҭV(�� �3c়��c'��bG #v�T�9V����j���mK5��u�~�}hj��dQ�Zv�E|��)��S&��{
��z�Y�͌��A�:	��"�\^ΙO{9e<F�]=�U }�*�n���Sk�e�`��,:f�]�)eU�6�̱Ӹf��T�ѷ�y�i2%!��w�P��ly�ڸ��\�R�6����|Zѭ͂P�H���,�������������֍�Ϩad�:�����A���`�`ʖ:�܈f�]Xe�4�Kc�H�d4�r��9۶$�mq���ڌ�L��:&C�VBp�����#��/��c��������I�=�f���"��(�퓳gl�ǁ�]�q����r�Ź�Wo:��&��7�u{��J'��`��=�9��6sNU�1YG�Ы�Ůl�C�H���؁�[{/��̤hP��qkYWy��0ə��y�f��ʤ&#7[`�ŕ7B�'�͹˞r��gZ��er����-+n�u��rT�3�u�ׅ���hx	��[��ۀP���t�/��v�u�kX�vm�S"�b��$:lwhu�=Gbt3K�b=�cW&�b��C��p5c����d$�=�0�ee��yj�j���Y���<i\�Rؑ�|C֖&��:t];��p��,�:��֮��4��o׽�Z
����U*�E���O�3]aݶV4S�Qkʮ��x�e��S|t��6��i����~���C���Z6��Iz ���;���34��_��g9�<-�`���%z�\��ĳ�P�m�YU�)��ĵ�xQ�j^���v��Ӭ�MЛw�*�w�^�բ�ت�{�`�EP�G*�!-��*P���r[)79˱��+�SW�iAd��9y+��Y{;Y�<���ә�穅�Vod��h�iJ�ww�k�p�_pܬ�撓i�]@�Qj������]�e�L��t>s��6L�Fs ��������
f���o��C�
\��4B%�H|~���'�P2�]�J��D����#9Q	��r���m,�\�o?�� U�l���>�����������Q5RHEO��A����_@�L���Z�@O�D�	��j$�J�n�LLH0�-��a��`�Yn(�e Q,�Q��!���-�m�$�$�`��Fde5q$�(!#��C>BA�^a�M:f�`���((��B����A��i�Pm2�p��"c8�17q�Y�!�9l��h��K�d���$�!�E}!�I�(B �C$��I�AF�s�I����~��T�,$�%�)�R
�FRJ(���I��L��1�I��O�#�+��UN���N#[ӮW:xjᖻ�
�/�͡���SY/��Seǯz;�g]�e"�;0rblyQ[c�rNc��S-w86Fخ�0ʢ��%���w
��}��[��'S��]�]B"�"��wX�X戴�k%д��WJw�9J�w�/ ؎���:`�4�Nd�K+��\�[E�s�P.bl�vnq�r�u�i��=�g_aw��I�b�Ah�뱼�p��[�h^�ɗY]�9Hwm�_NZ�ì�s69���\��_]��')�sڙ��U�˻�Z��|��KfK�y�`��b�mڄ�[��Q��-<0���-y�[�{�&��7ZL�h������.���i�/q�q��/�녭U���[5����'z91�QF�x���j��xm/��K:�ֆ�u};ꍃv�b�aӂ���8�lQ�sk ���zj�V��+2X�ݭs�S�%�g���jC�ZumY�w���8A�)ax�Q����	ʌ�6�n�a�t����;{��M� ����e��)a� ��Y��N��|��}��8��:�ܞ��x<�zG�N�/�6m��=N/�2�S�3F�v��z�M6�3`���I `o�BQ!��јB������IB"Dd."�h�D!D��P*(2���M$�!@����2A!��A5"1�j@�.�B2HM�Im��B����ȇ�����h��M�C2�H8~)8J �1ƀA�
e�#	�R"�*�5F�E(% E&�qF�!&�1M4�L��"SoĵH�2���P"�
0��$cnG]0�PTY�((�a�L���@�b !2b�Ƅ���6�D$�F"�I��dB�
HII��MFj���m4�mH���
	#�����dQ4h�$h@�0DY�~aA@A!"9F#�!��!A$%|�$�E�$&�$��1�L���@�>��	�"	�!	aB�,1�RRH�S�A#!p@�6@�� ��26�B!�"���t؄R���F~(8$�0
�Xm|B"DBSEF� �\p��R6bH
� di)��hR
%0&J/��DR��@��0�S�|�)5
�.w�oo9��w�z��z�k���k�nq�!�]J�����I^���K����c��=}q�z���N;i۷no5�����z�"��w#����6HJ4) ��R1��vǎ=q�qǯ^�q�Nݻq��$��$�!]���</�.IF�(�H���:vǎ=q�qǯ^�7���������Ib�Bl��q�.�I�L�c5nm���)�wk���/.���!�y��^��s����ǃ��qO9rm���w�tV�8����+�[w:�.����<�Z$�r㻍�$69m��rMݻF���Z�wL�r�v�G4�w6���[\���\�\��n]t�v���wwn�[��	Ws�9�wq���w$�H%�s������8v��]<�t^U#��Ը��,�^��^��ꩴ(�D�,�R����@C(�
,�ۮs�1.�?<�o�=�޼�d9\��������^:������G;��۲;9ݷH�&���*f�{���K&��lB��z\�@�Lm b* M>�{��A�@�I
�a�>�B@�eH��9������A�4����:o[oiE9�$Ap��w>��M��V�9��r5z���������<�g5�Kԍ7Ǧd�E.$��0�J�!��Ԃ(�l�i�f4��&$_#���8�P�T�k���!�	("rD.���N6"�F�I��)��I�
e�	H8�1��a@_�������h�QQ���d���5�����l���/�ْ�4�$o�$W��'�p����]��ʥ�c.}�E�T����>'K����E�6׈*�q%j�I�j榜ѭ��@�e�3����Id4*�d]ϫE_��4d���sa*����Ie@F�j�X�{�L��C����9�4� S�nD%ZD��Gs�;�Ov�O��v�v��eg��w�_)"����2�N�`��W�U�Sd˿�2�4N]��'^�IJJ�eJ��&̷�	#�q�c���$Y��=����7��֯a�۟�2���Z_g�� 6��+�Ff��H��4��p��h���e#$�bU��<��e^�2]�{q�i��ݝ��H�&�-�j#A�B3 8Tf#�(�F�+h�@�Sff�,0��5��5hؒ 7,0㋨�ddG�kb�4����0_L�:83�Nb\�+��o�z>�_v���}>1��V=����5kV���
���GV� O��k�H}��r�����u�TN�D+�`�b䢳���Tx<�h��c��8�
u��Ɯ:�9I:n�т�����>>>o7�� �`ǊWu�`o`,��`�.�W[<��17%%��CԺ���n���������q_L�*��ERH4�4Ϸ���m<#]ٜ��!y�}��%�6'2�^�d�Y��RX�cd'�)F�E��Uϝ�LO�54��2`L{9����'��_��RU�^n�F�y��1�o��R�VBJV�4�R���*��5�����H*e���\`=D�g��p���u*���7#g�_}iO������@�Y� �,���]�K�y���>{0׸v�^F�k3��vM�V�ON��Jȗ��A�P������h�\�߲[(�f�ژH�two���%�*���t�Ao8U�ؑB�+hJ)��[bJ�\W�yD�$9��)h.��6ʔ�۵]�e���{����8ѹ�+�{X�Bٽ;8�I���7[�[�n�]�v�r������u|l����hIY[廳ל���!���@x!���g�S�ed�2��SS��p$�iقX����,l)�r_rݪr|8F�y�/9:�x7�ukx{<||||@;e��ܲ��4�7A��G~�ל �{p��T�[-����ݍ��4v����|îf�A������Dld��[(ϒ��wZNT��-���iQU8�c��:��-�Z��R�϶4�(�C
�-ʆ��9�L2���Լ���ꬭ�q�d1�fǜf2⌧��۰��x�;�ԍ�U�UTC�(K�4�fTdʯ<��g����vd��{t�娎�X �y���٥�$�|m�����j�Y	��V�VM�L��֝H�f��*L�Ü�.
u���⁯��%
¯;��V�wڌ�I>	�����ªu�	�$���`\@!d������yi��y>o���A`�c���Ww=���k3��YL�b��.枂�+��l=�Xr}�yH��lk����7�[	��U�t)�8�=b�n�����A]���(�zЧѺN��b]�{�Vz�ޙ��\���#�ZB(�v�)���xp7��V�6����ߎ�)�+��o4���bHq�\��9p;�f�>�o"��p�w����� vƩӆ��PH�W=^J��ۡ)�``�}��?%�6-��7���m�Հ�����y�FM�ʵ~�Ƌ˱�/Bi� o/��Ym�I�f��P3�H[�N� ׉��l%I�,e�����>��I/�.r猪��a��� VǠfJ�#��*ו)ioX93��j���f�IZ��>۔�On��Ko�F�:��ˀ5`�(��c�F��ԣ`�}(8sGi�n��;`�%W�#/�{�"��=B�U�]/��Bݮ���^/hZ���eiu�e�x�����f2͸�IPC��n1�S��}C&�5�~s���ݮ�`+é[�L�&�B%T������d�����ΟK-�D�i
wI��혼�ô7���i��T[���#Ny!@S����N��H��l^1���1 �S�N�z6sal4^�!e�q�QWg�X���Y�iM�c�K`��9k&F639�$��6r�Nς�����Y�������yh�4X��S��ٸ6gA@�]<yj`[6��bk�wtW3�!���Ղ�������+���@>>�&�mL���.�����㻣���.�	���.'�k�1�Em���\5�l��
�N#-�on���l�C���Х�Va�%�i�h(Л�]6c����e�SD����YI����{�d��3h�r�t/i��"�y}�^@�!E��)��S���C䫯��7]����?M�)U!����^O�a��$F�e=�#9�����Y�ιk�0�5}�9��9��c����7��]�����*���ý�.��B��;�
��ay�U>M!Z�T��j���B�5�@��,�b�<��E�Ym�o6�_��n2�"��5UmE��Xم�i�Q�4��Q�%�4���̄JaD�к����2�h� n�Ļ��cMŠ�)�kz�TO�f��d�F�Z�0�V3M���ܗ�w�(�FQCahY�M`����Ԉ�e|��_϶<�Rg��r�-�M���Y_������l���i��tgm�RRє�3�rQ��:e|�?p����c��Lߋ�*׼σ>�<(��B����r�jz��gb쀬�~�&��\5��������g+�ҝ]7#�/t2�\�U�պ>>'D'gӨ#-<���V�����
6Sj�+gt-�u���P5�N����&p�b@W�%-�{��f+��YY
����E=����F��W�����7R҉�R^����Z��c�2�ɴ��E!����!��9a����.h�NB���o��
j�X�C&�gv��Ilڍ��8(`�A[ees"���f^�z����5)em������/��^�Y��&A|	C��9Nb���=$Yd�ݠ� 6����_���N��wzR�i��2�q���찘4���Ok=��[�8��������5.v���2�M�J��J0#����@З������JEi
BT���e��e�k6&�f�QSki��M
p(_�kzWf��HU=����DzX�F_�^��͹u�f�)��td��n4��7�N�+~ß}ִC�ܹ�7�E����]|�2���K�~> �����G-;�k�ȫ��}�y�E��{&�¥��N�`�S�ojɝ�˾ν׬�]]���)�z�ozxU �p����-i���{���ȩ�R(2
��"���Zom��["�"��>���C:��jB5����Jzly�Y�Jd#w~���*�<
e.N�5�J�ջ�c١����$���UA���u���~�KF�ц�;��ĳ�j=Kwa%��"��䄷df|�3���3X�%�Ƣv�j�ffF!c_��eȄ2)���T9�2���rZu�=��F�t��S~U���;��a�c끖2�϶�Ċ):��m���fj��FuC���1���ml�(��r��s5t�<��xI����hN���������g��cG�3
#M�Փu��Xa�P�f�봒�T���wn�_.'��Z�{o(;g������Eř�����8�#WvbZ����s����9�i$�|���2�9���Zʓ�_o��wWS����Ѯ1;��:%�eħK.�krռ��-�9����|�����]���;��;[1��pv�3u��7����e񾛸�s�l�HA�i����g93P޵=֗w�x����VA4%�"�u[B��&�����^�~5�&��CWl5��/���с����A+�}W1��{�א7N�I�f�oig4Y�Ks$lS���|�Q)�U#B* L�$׌�k��+`�*Z7�DH�Dz���2��^x�����z:!��iۇ7�x۴�)B��ׅ���T��Aۊ�s��3N�j��ENT�īa�rEp͍�(,��*܅U���jS�]�jޭ>u68��	����gw^�
]���]p/��5����I$*�ɂ�#*[mZ��x^��f&)����N1B�9�k��H� RZ�T�����C�%Wf�T�bl���{�^�9[0F�(���:��؛��4���6A������;[>a�S�fǨ��9v5R�!���Q��y����b���T�R���{rчh��̴���S��d�[��3����a'Ϻ��~��- ,4|H;b-ȳF�B�-��r��}��#���U����BûF��Dś������_=wo��'��R��!U���b9�/���n�w�]��2��k|ʜ�,һ�����Y4�!T��%�iGF�H���[3]tT�ZPr$VRE�}��vq�|�!��[�7&��Qeyr�$�eZ�'W�n�x�%\��}-7>Ib43����!Z�z�� =�z�1�l�hvvl^a�@��-I.w	մ&�N�;Y#i�k7(H�>���b�Ԙ���l�R�K�Q��Kh�7��<�"��T��5P�&�>�l(�wf��9��L���k���)�8��;�c�S�&�_Fܙ�S&Z��^�J������z���4R9~��M�MI&���܊JsYv|$�$i�6&��/�)��B���Z�?�ԧ�6K�F顏�ʚ[^M�IJwƮ������,L��Z�_N7�>Nƨ�\��Kh6�����������,^\T�ӌ���T��ے�e�^�1��oRX.�B�:��R�IǩO:�mE���"��Qk�#*#^oL<a�+6��[�y�^�?$�Vbܛu|�j1J,|�d�PS�.�s;D�qDo�E<9Gɺʀd],�,;�B�*�v���1x���U�����%5\	ײ啙܌���c��]�����_��ַ7�w
)��C�W�#g6ƬW����t��f���=WmnH�[Ӆ
���^��0N���`�u�}��/�'�B&v��*��S䒐�Z*]^3�L���' ^�����f��p����%~�N): -7I�0�.T���vuӹW�d)�%�ꭅ;i��ro36�{M#����!+φ0���i���Y�EHͼ�b��=E݆�tf72ќ��Q#�nϕ�+b+)V��	&u���2�g	������دJ���t�6�D�K$ �*�%4�5�A��6<g���u�l~��;A��d��l��ݶ��HQo�T\�^(ՙ`ha�����h���k�3wr��q��T5�:Z7	�tI2)�ݟ�����{�}�eZ^�{�c=�qdv�5툸�ӌ�ز�@hoU�¬��o]gL���c�ݕ���e�����l���}�������w!.oNܵf��Xv������]C�d�Q���v,;�z_�MSX��/�c�8G���n3G H�f_M;�@xX�
]�o��ػ��}B
��2�̭�l ��Ɇ��Y<5jP�4'I�-����M�X⭰j��WX�ywk��\��������،�1@��X��\�<��pJ�v�ǎ��62��-�~͸Y
627j����2�ܫ9ڳmw�}kUi�Z{9u�Km�}@w<+7B�`�3�P�z�=���Պ��@�+�n٧b��bB��4���:t�oQ\��C��4�Gdo��9i�[|�R��-urNk��2p.��S�s���m��"�&P��Zu-�h��A�2iR!w�jG6��vUͳl:�77K�9S��J3J���M�Dkse�x�"M���y����[ڣ{oܩ}:��<�wBiqg�u�U�ە����G-i����B���.� �&颠.�#V�k��L�#��xV� 49`qL��r�;����wg\�Mz����%�U�Ʉ!�4�;U�β4-����._E6�4���ۍr|.�5��u�5��-�ڢT7�uQ�d�a}6�Z�C��-"E�X�%c�,@�0�xrC��H($h]��N�sh+��8����W�~���G�r��@K����у�t��h�I-cg8��l�6uY������TB���]�Vf���M�c]����zS��*�Gu��[���a��1��ؚ��wvE�A^c٩
�9�0.��˹O���x��D�㔑�-[́��y$le���9�d0-�ze[�W�fI�&9.]'7�}t���ϸB/��絶΢DN�*���6�X�b\2�<d�z^]��Y�.�6Œ]��["�0E1�o$��ϻ&��u��gf�n�&p§_5���������+��]�:#�&-2��Q�W�3�����1��)x�ls�V��K]f�9XY̹Fwhh�c��J.4=�I96CT2�GLt]�]��;/Ӯh##��}5�H��C�]e�k�K"oa��Z���&Iaؖ�B���n�S�!6�d��踞9�Ե	�0��kr©b�����*n�P���)�WQ����U�Z��O=;�55BZ�v����lؽ]��#W]M�����z��C��d�������	= lȊp��Ǣ����\���fV���Z���':��p�m�&��	dM�[����*��pS3������|cK�,dS��b������E��;S�O��1���~8�__X��>�w�%D�����JcDf0Ϯ�S��I		����o}}}q��||}}}x��O>�y$�$��!I",�+�[��d�2*a�t	�E <��:}}}}v���\qǯ__���o���|߻�������P�&#��7˷'���/V���9vd`���(ɈJ��,�h�S"(�%�p#*5��ޝ����F��LEz���� �*4fI�"g�tE�����~9���Ҿw0��>��>.����+�n�˝޻Ʈ����Iby��A
"��{vzk��͈К� �j�krK���:1��Lh�]\���(��1�Ÿ_:��tB��MzWρ��$y7��:르g&^o�:lm��٫�S;�d�`�� 7nb�.p[۔mJ��O{�U~��k�Ƽ||��	�*��� <��`�oſ ���Ȗ|�������I覀̧�*��upZ�/�����
���:�9�`�o�X!P_Y����B*��^���WF����?��W�Iw�ȴ�D�@%��M�{«g���v��h��K5��5n��=��z��]�@9�����A��)�3/�s	�zܷ��\8x{�=�Ѕ��ן���c����N�<�ä�dz[�9�ڹ��S�nk�O�:e�3}���t E�hmn����P+�"���_Z�@>��O���I��(E��^�#ö%"�=�/���0�e]I/(��K�wD �V�Ys�]�M��<k[� 0颼��V������}B��nM��s�7ۭؕ���,���,�W�`�2�Λ���D���LWr�`-�A�4��\?W�_u��ւ�af3�����c=�xt:��X�XI5���ߘ�Ȯ��E�jJ/ɞV�[���U�����y�x z��S]Ue�=��b>�\yE�,n��5���'�ߔ_��!4��[����ct�����Q��b�����w������f��J��@h�p����Y�<7�Q,���Q�/����tέi�h[6�n��XnSN��X?���y�cO��t&>Uj�6hA��QX�Р���;jR��� N�WNGϴT*�cwf�-�W����m$�J�v��Ǌ��ͧ�dc�3s���>f�����M41�N�1%Z����LC�����4�Ⲉ~�6ԏ������G����E�f�����w =���T$���s�~����B�!�Lp�WA�2��v�L����21d(Ã'����zl�+�mO�r��?V���@_�s��7��[hy����D�x7.��[Qo��{ffE�p a���7c���J���86�<Z��xH�H�G#�����~�/P��е�I����-�=��{�x�n�J�n�ɢ����:���D3�d�����C�����ʱ�� *�����0�á_�oH��%ϕ��/�]�]�����;r�0Qr;����������w���.��Bt�Κ)����b4t	��Y�upK��R��y~�y�j������j�]�x�AN#ˣ� �����5{��f�eyi�P����;�H���M�k29�K(���W6d���K��݆y5����C��Wr�5��q"�*[���7H��Ʌ��k�����"�~	Y��q/�V���������ИSW��������U��+�;v~��2��B�6��_�Ӷ	�����c��+^q+z�rB��3R^om#/i$z,��3
��hƷ��r��`%�7������na�T{��e�P;�Y�t.F7��R9���8�r�t�]Ɏ~=�ۺS5uy��Ve��ݕUwo��<�D��-��k���ʖT��+�tj����p�e��[%єl�خ�����
�Ϧ{��f��Q��U�˯����M�9�{s O?X�T:�g��Ȟ0�өX��Z��触�*=Ҹl�z=!����������m`F��s&�w	���·)��p{�� ^^�k��C��88�yf�v���U�U�G�;�Z1t�>_Bi��sB` �->��4d�gmu�u��n��YZ�<)L&��wE7s�1��>�->�sQ ��@Q~
�6`��|~�ώ���kt<V:�:P�����R5�<zS
�O�����7��v�S+�N:�xw��-��f�?0ޱYGp��P�]�_��[ӯ�^y�z�@�$�iu �U��7�>�5�+��K�k�0j�K�I��?Wk`K���l���0}a��ό��ͩ��Ⓙ��`��� ���V|}��>�	��3�2Ը�'�3�.ny�H|�4Է���h�e�9Jk�ݕ�`�9�װTxN���k���Y|��{�Ju�`��Cq�pjÁ��O�Nb�FM�g֋\[Ԙlsklgv<�҃z�8xbp74jD�w��O�8%�;CX������
0�ύ�p���ĸ�u�f+]v:���|YY����`�܍gho�{���r^VK*L)b.ޱ��Ί8+6V㻲[
]��־�϶��St��׍^˘��+��l���o����9;L������rHGj��U9f=hi�ڹ��K��7�y�a� &��"/ ��}� �{#S��)���V��>��2�0J��x;��IB��w��n��g5�����yQ�w�$�Z~ꖽr�/��A�e)�O��[��f.	ך�7��78��{��;����R&����
�|ۚ� �>�����f���eK.�$t35�p��u�0����0�w��WT+�gIa`�遠�������D�]�����[�{��:|����]Zv��P=�5�dw��Z��[զh���}�!��{ӓ���Ɵd)�1b��j'%Ů�ս,��m:o_��P��7{eu�ɼz���=)��(8�[�#���	������d��y�s��4� Mm���g���pS3X�<�!����]{ޞ#V������;#�!���ڝ�Q���v�쒼i�`�g������ 8��~�1LP�6��v�HH'�TK�:������Cu�v�w���{��&� �7�Nb�j�z�\ ��/K�Ӟ��d�M�b�8�[.�y�.�9�����×�;�!��&�@�Ο��m�>L.��R�P�>Jޯ��$*��/��y�y�>Dt��|o&���B����[�#��=�u�:�MK��N(5-�omȟ߮�H�W�~�fǮ���n����w��?RJ[_Uj<��c����p�ø�X΀��EL��{�:�ڐȲ��
5��k2s�y?F1��b���5��]��p�l
�ï�z|F��A{�j8s� ���>=#7}=��+���\�MwWs�w�9okl��T�e{b�l�
�!�-�D��m��k�T��,�J���e�5%��Fy����g�zu��(-#����'���u@�;A)��$/�x�Xy��h.o�g��e5-q��˪44l�w��iu�G�6��~[�z���#/u��h�!���G&�RކA���ŧL��j�;[��iw��q��e9[Hy��O�30��h��1�[ia' �p�%.�_8��5^D-j�o{�:t� ��� ?���Շ�|�*�[c �U�Е�N�����j��;.��<���
�8���xokv�i��>k�i���X
����T�SGou
a��&�W�F0�{�}�Fxo-���l�e�c�:�"��'a6��;c辞�Gv�A����T���`����JL!�D@h�*X��ɪ� ��Ô�^���z�����������1��ξ�36��"�w�T�{�-���@���-��� �ݞ�/�W�1Y�kEyQ߱��"��?_<�nkBc���Cj�F�V��-O�j��ݿ|��H���+wJ nBG�X�8��v
���m��1Z���8��vQ6z,�s��w�=�������������6����m�r�|,H[k���<�5����]�|����G�-�ό`�c�RI$�~w�׽�����l8�p� P�
&���s$��)��t�Ssz���[9��Ñp�����Yv�&wz_J�ޯw�d�KL_�^���i��a���c������3��2�
�΢���LM��A~������l�ͱ��2?�M�����:͞3  �F@�y���H܂�.R�_8
{��q��1��-�O�_����r֐��o\>���8X���#L��'��r�0�W������Q���{w���x
b^8!2oCQOuP�ă@4��DW�������S�KyP���孴��Y���>nOk��=�b��;<�`j�Ws���w��Ф`�I�D,�-#�g%b�K���;�׫kkH��fL�n�]Y��/Aj|)Q�,6�Ʒk���IS:�_mǤ��#a�Q.Y߽�lM.���a�����1�?x�|�Y�ٟ|`{�iO�Ul/˚<��9�&�k��p�זj˽sy��w��CԙT�����4��������c��f�
'}4��.ɯ-�u1{OC��9���[��&|@�Xu���erO�I���8-i���n��4p��������˓k;��H����ݷ�ȅ3[�� �Q���{;q��v(Kx��q^�Ǝ�f�b�ֱw-ڼ�h4��F(t�_$�����n��t���gն�֒�T��'r���s��3�L[R��n������j�ҳs��3�y��j�滣�R}4��h�c*)2�/�C�����r�g7��v�x�L6�kҞ�������k�2ܾ\���.N�p�G��'�3��D	�X�j������%`��ջ>��8�<��6�N{��-Zk���&v�Lz<+�`�M@w\�n���m�������c�X>�gs�x�>����U,����������^���Kts[U� �L��=�va]��q|%�� Mv��(a.��[B�kOC�oB]���1��5����t [ޒ��5�A���7[�;�u���=%��ˋ`9��=���n�5w���Z�'TUQ���]+�x����d~�}%� �~if�� �;�~�S��}G���D�uu��m�����p�:m���m��ׇ��οy
P>���a����]S��yR�Wp�Z�K.��6"�~j��W�س�k��ަ�F4���~b5�s�Ct���L��{��Ʉ��$�ڦ~� Sr~��4��W_�kQ �iQ`x!e� 4j�o^�!�e��iw� l4ǜ<;;�1�OO�����%��/et=��ɽC��e��i��H?s�
;��Sy����eV�'�y��:����5���]�ԘW���龻���cK�p�8��X��Z�{�o�W�^+����Jkčkd�ȴv�nl��et�S-�kW�J���<���yl��Ǔ�l����#�M8;^�"����̋���( u�2�3�u�瓣8��7�k.�Gu�|����4ݛ���u�Z�5����K>,���L7�-�������`�������b@)�$g����Jo&Ã��A�f��/ފ�o���O�k��~d4Q)����-(<�Zaٳ�䷂m��4���k�m���n���g���"�|Nw#� (+����Hh���k��*>��WOl�:Z���A`L�:��`;^mٮ��o�*���y/�b����p9 !���J<��Vc���μ���#ϩ�C�>0�^�^Shx�D��}����xt����fNy���T�I��@���F������ �k�p;���HG5��m6F��42.�uxN@I�^(pٔ��;|`i�c���Ï��{~��2�Z2Ώ���lhK����� ����~q~���{��xI���]"��!�YtjTk��[���F4)���<��oL>�b�o��{�e�!��/�xcA�V@��'�4����܉LgZcN*;qűAR�����Tyk��o��޶��{m������l{�lt^xb6�ەV\���V6����Z����>�a��'}B�:���+�W~x��@񯳭�c�+0b
"�k�=��:7�σ;��`e������?	�c����>���ɐ&V�׺��G_r����o&[����4����H]x6���N1�(>���ؑ� V7�ɴq�w�N�ugA�o��fk�=ӇvM5���o���z�s�~eo�y�@>�cBi�*�4*��AO<���ʟ9�> �&�K;D=zX��gڢ58|�%���=���=��)k�B�����C�|\
%���y1��!v�Ni���-�-�C�dޟfǇM�'�&m8����c>�)��Ȳ�c���k���p*���dns���ǝ����:[jvB`Lo�{D�t?��k�S�=7.�*eC�����]���5x��7�8��a֐!��~�->���^5�~��җ�}n��\�qz�|�"��qT�F;�M���������˞�П��.�H/ں ����=����K>A�&�=4Ȏl�˝�����.����D3�ɴ��h~��w��:�y36[�Wf@�9W4�\���.����� �x)��R=:�A,�����K퇆5���t/u/:Ù~}�Ω��R��=s��w��M:�.s���k�y<�Y���e�J��H�[�R�=�yw��MqϼS7������h`2�w�}]X�%��ίd�6@9V��|7`��MO��k��ja�8�QGj7�-�=���[�������薬yW�*�Кݔ�9T�3��fz����j��'Z������ۑ�y�CY�=MGLʻ�j��a�Z��\�U(SZlӽ��D8�,tϓ��8����)_ekr	�c����{Hھ�l�������wG�:��$��vuVL�pls1����N�x�xo�y���i*+"hh���**+"2
潩ߞ�{�� ��=h~&0/ʸ��f(Q���f��4���W1�/4��Go*��1� ��6Q2��$���Jm�`�,���n ,�A�`����]��#��t[�n�I0����;u�t��L=��"K]�5��p7��q�#�^��O���H��U�ȵ�z��lX+s:=}���`��?�u�4dA	���K$�wM7Go��+�q��?<�S۾�״p�vV�]�����x.2�1�N&����{�d�Ⱦ��x�p�M��y���䅷�F���/*���<��g�[S����� S�:�S��z[�Bn׫�@g\s.��|)��'z�WB7��7����cp�!�:�;�|ǌ(W�����~��6��k���^/��/7m���Ǯ���Qv+�,zO��ֲ|^F���0�_�l��!�����5�o���87��Uݒ�櫎5��e@���@M��feBPK�o�#�|�����{������Ҵr�qQ�u;��$��6�7�\Kl�Mw�es�W��z���{��6wTܣ��BW�v* �|}�\��?v|Rb��y�卜ReP��`�n�Y#\Y-j�����M��G-okz�ov�T�:�8o��#x0�{�k���D��]�b��H��n�#��_9$���3�Na��Fg	�n^�:�3j�H�ۼ�]���wW8V.jA�*�������c��T�[3}�!�ᦎ1��7]�2��hu�k�(��*_��)�.�d�Z̽�r�u�&7����w��m�жlk�t�)��S��qa�7�=�n�#��{4���J0iҁ�EQ��U�'��r�+����i�rp�Y���@a��9����]���ї���6Jrn��"�Yk*�Y,U�>���F�Gh�F�������1�����f�Y�r�,�n9��m��S&1�ga�kݻ��+u��^��#�/M����+�a�w;fuJ����9K$���,�Ӳ���Ƿ�;!}1�-v�
ȕ=ۤ�K��%c����ОZo@-�$���pޣ%�Kf�X�wq�u]d*!�Nn��F��X������Y*DݸK�[Γ�y}�ۮ؊�Is0D�.�;�-�\f�ևf�T(K�V��b�k�n��Q<e_^V�;oV�^t��sy�q�f�å�Wm�����L�g����W$�f��l�JKX4{���]%����ne�y�Г��ۂ����r��̭&z����h�̈F�P�K�D��
��OGE)a�e�~D�P��SDl%D�N�N ����5�	8\L���Ӳ)���aHq�Z�H�#�M0K$�1��_ȢӶ�J8�N��7l���ps��^=/��W���+46>�g�sAB��=ޫ�N��R�V��Ot��l��[d7�:��6^�Y�A��VW�fX݌��a˷BBq_S��Wt4����V�}
o�PGj�aC2e	%���;.����/�k_��;��3P�x�����U	�+h�[+,�r����.�5�&�#t��N��z��]�ىJd\�VΞJ�fe�E���7Z��f5�:�ڍ���iP��Z�qm�ԝӲn	����I��VՎPV;4:U��՞������T�Ӥ��Rt�:�&�����y"����HT¸wo�Ka�ٜ"̻�ڸ����P�)	s7�3t��_�����2�Yu07X�6�*��lI����X�"�ۻj�G�b�cT9�M=��ɆeRj��P���c�%6>�X�����Q� է;������[j�ܸ8�9V���B������=Sid5;k��(��C���e������k�K�RE�Yi��P1���U�:ξ#�^�n_Pgr���ǰS�|:�.f껝�ǈ�׶����vݓ2��7��jz{��rw����*���9;���Ƣ��Զ=��ke������*.��m�t������x?x���|� �K(R&���"��A�HC�I촒$�����뷏Zq����ׯ___^<m��ׇy܋164BF����̦4��(�`�=}}v�����___\z����׏o[���7���lb��wE��[�+��N똫��K�q�<��W6�'��~��������}}}}}q��}}x�㧎�l�A���u	Q�bScK�.���ZJ4�@���#ԑ��d��T&�1b4�DY����m��w4��\�/	$c%~.�?z��M&"�X�Ҕ������]'��E`�3��F$�lFwV�����z�k�^+�u��U�d"�K}7^=���RE��Bf.��,cj5���wv�4Q�Lb�|r������}�{�_]y�]�z�"��H$)�1��-�ѥQ�$�##���AH�E$�?�%�B�JŐ?��J��m���o����Η�m_��9�e�Bp:�`�i�b����mخ`�e��N�14� ��!�	)�~i�������'��ċo�bm2~@��/� �r($\o��q%�1��L��I��"�L�D#	P�SsVUl�S(ݗSUe֚+W5�U~@�AA	�� ��ED�[�y�|��>E��.�ݽ�ث޾�C����
��;�Tj��Dqo�PuN$gO�Sp-?�;k�=.�$���Xn�Zi����>oK�C�`�v���T������ �>75Cߓ��<3o���Cz��SL+�Z�J�-���:0˭��[�� ���^���@2��^(���ɿ���O�C 8��G���1)��b�e���i=��g�i#g�� ��W�%�_�����j�!��2>���^��ά��ዝ&���t�ؤ{�Ti��==����n9�͠�i��F�C�y��Cg��A����g���O��,����.�O.���â�\ ��z� �ɫ��C���	�>�Q^Z@�pcx��@=�ٹ�%x���4�â�Í�5�kj�OK K*IV�J8����R��Ԏ�/7�y��,���
<*`s��`>.�;��1p���8~�`�ɽ^���=I�7Fhm��Ӹc]]Uo,w���oL��X
g�!7�tt�.�1������_#���9��촊�+Sg��g<i��B���+�f�N�[A�O������B~���F�eĈM��is�}������&e�Hsvf'}s��ղV<.�Θ�iS�2V�]3�*�[��2e]�4�t�yN�J�BS�����ј/���T�u�UݵM������t������U��oY���nl�ԯ���
�{���'Љ����h)����� `<<<��ҧ�OZ�~��α�s���^�+�޽#��կ*|����ș�>
1��;�Ͳ"�p]L�Oo`�\J�aL�F��w_�����I��ݥ�j��{�І���� ��>jnekόz�t�n��$#υ����A���
�rQyj�s��0	*���xw��#S�E��(�[�7�.`��uC�2O��L�r
qIt�|d�OT���ǯ��Vה�����藾�W�L��hy�0�[�Y�\^
��)�=�������H�Vh��X�8<Xr��j׶����X���W�$����/��L��n���f��c���o�s���렜A��@���L�Gy�m#�<#X2YkZ'�W���8�k��}������La�w�sܨv:��DS*�l����0�8(C�w�C6�ݗc��(�[7��U����d$!v��`�$��wў���K��`��=x�[����l�,Cպ�Äi�Q�xGX�N$E�1e�n՗V����=ڃ���>4��Nz����L�#7���G/ ��9f�Y�5�2��0�T�s�1ֶ������ߎ��G$S>-6�	3̙K����0�|�s5��
��d�6d���sJ\Y�m�6��m��1�����&D5���i꾓��E4�8�L�L��m7}�{�i��)��iX(,��|�����T$$HC$kK+�XA���fU����SF�m^��PYu�eԕ���(gC��/�� yK����{)�[�|Y���ϳ���<��o�J�]_����%/�_�p����������APuU�YF�(�9C�8���@1��6�n�zk�bkn1�w��9Z@;]YS�9�H���ǭ{+�R��!e}���#|���� �˪���e˸n�;`l�F}�yր�%�o��#(a�os�7`�5��<z�Ɇ�̘��qkBqS�/>f}�׽Z��l; �lNK�&)/w��`
k��
t��b��ݦ��4H��E�F
Ψ��m�.c����;�X��pt۳6�dOQ��pqA��T_9eΘ��*9�k�M>�{�|F�ڭ���.%����64����vt��L&�1j{�]��R����oڟ4��tQ�:�nK�M���ڨw�:�ۛ��H����^�ڎ�dKq�~mw �SE)��}��Ua�a��Ol�߽ Ο�r��>�����;#�`0d��S�6�2q{P��L�sn����P����}=׽�`��B�mY�J���oXw1)CZꫪ�vF���rP�����l�o� ��j��|���K�������L�xC��슢��<�'/"c�v+M��uk��D��M�v��<�;�>�W���"�CH+M �QQP���{Ҿkߞ|�^�׾^�kd��/϶��z�\�-!� �v/��(h���5+�_�)r�}C�K�i�*,�	���@f�C4��&}�DS4؞-��a��V2�1���F}��{�gO]�dߟ�|���l��s�h�2�,ܥq���E�{Ctr�{g�5���k�8�]	�Y���æ�zދǵ�l���P�;<ê%�fυ��b�z.�w�Ob���Ԅ�v~�@j���ʫL3��?����_-X)S=��8�Q̟Lvjz����)�c��lP\����s�Uy㉑n�[XnO�q��-�:GO.��1�In��9��g�mh�R;��Jl�RCsP��O]̻լ9+��@U��@Z'��_w<p����Dq��iN�,�j���ِ:��#�q@�d���[���C�q�S?<�o-y�#%
����\���5�����){dB���5��E��O��~�l{��S%�L�myΜ�����-=C����P-�;�L9�Q�>n�%Ɯ���N�ˑ}Vtd��iU��.�Ҩ�-u^�M����;O�$�/��8�3F�	Zk4.`�Ǚ�)�zP=UĞ�A��*��K �V�U�7X�y���u뮮���VRlwE;�ڏI��I���Nl��M���\��V�m����Ux?�V�J�$hi@��� �{�����[;�}����!$�7���ǥVŝ��ȥKFM��Q2�\7NId��J`���y���G�G���rj�k���L�٘����n#�'�t����7_����h�Fi�.p�!���tj��/Y��=�J^>����N�[�
����Z����;��C�))��#؇,��R���íqD��}�K)^{s�pg�k|$����F���vL�qC��箪�� Wr7�i�A�D���i�z�$����G<C��GA�^h�wUEÒ�����x��{	�R���O�#�{�C�x���b��o ˢY���|�9�:��X�8y#�3��׆n{�R2�;���S@;�ޢHOg��p���YdM>�����&S�������:��8��,F:}Ւͩ�{#�5���1�_��k��֏Lޚ$�ȃp;�X�|��A�!����P����W҂~S���sK\{e��{�*��R��.���(vά7��}��	CX�����-6t{�w6m歚u�8�O��QM�98�{2�=��^�R�)�g璽Hd���`��m�M�@U��*����Lt���έ5�WU�ʤ�*b�^�\�]��EjY��f�6&�N��M��0ʔ�9>�o�Wv��k��^�z$���q;+�٪��t��6.t��\�b����fܽ�fa�4i�rhw�� ^�y���Ҡ��(�^����'Ϟ������c�
��v��k��گa���IN3��p�;��vpEN3Wf�����`����pXsP���:���[���A��,���]%��92�oj��A{[X8a��X��n����ϩퟃ�{�@���{`E�>�mf��IҖ���*8�e��$��ʂ�����v-��N6y�	���p}���,�5�[�eNu�K�;ÀޕE�Cy�wYyʽ���.;�I]�D�1���^��煦����7BlF�C�xP�L�@1��r���ҜM�s�09�����f���D���g�:��~dE�pH�ɛygs&%ڐ��r�Կ1�Z�$��	�^�o��j��.�ʸ�����^mv��}V+��E���d��r��C�Siz���
ÒS������P�a�f�0�uf���q��v��kӽ��8z���>`�ye1�(��E.qܡk�aZ�v��)'�L1�ۯ��P�̼�Ks�g�`���O��O��z`ag�h�\�,_T�U�ݺ�fzA$�;��5�$��wf�����uu��J�N�n[ٶ����{�-'s_�/����M��<����:�����jT�Ӎ�ipT6��f�9�۔�����я���o"C��ͮ��P�u��{��=�{���҉P@#CH�M"�����ݹ�����1������8���PfJ��W��gF1����Ed��8�,��q{JRx`��牝^�lV7�sG��1\�T;-z*�)� `[:yחx�s�g{w޾����Y��]^j����ӳ��H�v�3 ��|:���,M����*m�C��9��{�I�OP~���+[�̥V]^�;�F���ʤ!Z�y�����|u]�j�lVh+�I�KN�mp��t��� ���ϣ�3S>ji��CZ��0>�~x��>��&�8�eoR�Ҿ���PS ׄO��-�_q�O���Y~'��=Y��7u�軬b�v��r-N��rlU2�s�W=�-�^F/���i흸'��G�Z� %�����v�;a�����ض�l!%�LO?X��st.�[쬄qY^S�V��%�c�=�������{2�#l��^>{��+�xWמ�I�1�e�c�Su{�us
s\5�G<�`x���Du���^]���S}#�4�`u:NA-�����1�e�g���l	�UT�dYy�wl�D�/V7s��V]�E ʹ�)�;}\xNa��Hs{׷$�>�m��҂b�)�JC��!ܼZ��B'b>&�ˤq1+V��C&L�����Ч"�t]m]v���
�h�R,HFtb篮.4t̅��y��W:w��j��Q��h i�����F��Ȣ/s���߹���|�|��	Y`tu�p.�_�1��-}�+�����I��T_9b"�^�CΫ��F�{:�8Z����h`>���Xp�xU�m>�W��<�vo��Ճ܄�k��,±��;�p)r��d�#u����I�G���6��^��Ü%Q��,^�L*����xk-��Æ��ι�z�]p#ʪk͗��6@�����n���G;]]^]mu�'OMއf��� 2�6z�Г��}���K֨-�oW,��������@f�D�4fe&����������2s��G�%�M�����ߧ��Y��3�tE1j�<i�s�����li5�GSv�;�!��pr�H������&��A��۵�I��@�Gr82��e�G�ҷā��_RQ�����2Ƌz`k��G���K����u��;kUj�K^OT^�0�V��k�E�Hgyt�L�)�L5��1{�N5�̺�k�r����;5x�I��v�B�jn��l.Y1�͚���ǩ�𤘰��a{��'#�|��x�tj��N�*�f�3��ES���3ik0�,�Z�k��b�����s-��P��vd{*`��:�n���p���-�<8��Ç9c7�{�T5Gys�,��r��8���k9�yYpL�&���ו����P��i ��i��*(2(�H�"ù��wS�<8��L�I8���3�љ�m�d`7�o��p��[
�g������y����C��U{ݜ#���Ui�P�O1ߥ��缦v�1='V�!�� ��H�Ɓ�^'=�4�s��w�xx�W睻�zɽ���������ߌ'�-��u�pJ��R>^=�՟9O�:�Sw+���X���Y٪�5�[1kt�� �I{��>�����}���k���gR�S'U��1��ٙf~L��\�Wy_E&�r�O@>G�^�W�2ͷ0Cl�O�����N�n�m�^e�-ʂt׻[�G7K�z�<�t���?qcg��{��� Ꟈ������u�Xt�34�
a�Y������_���Y���]���(������s�_��x����W/���e���V��{aݵ��\Èl흢�~&{�v=>�^�G�T���n�S�w$�\Ki�a��B�p��ʃF/uT�It�#��L6�Ʋ��3�3��9^ �w/�:!��/p���vЇl�`��� �W����%�=ѕjEϯg�����0�����gX垚l�je\���s^�ϥ�Z�֥n���s[˕�^!�nῸR�&j���=b�Ǩ�3�+�q6녮=�𡓆��Ke�ܝ�w|m��b2��S�ɸ&�9_��<��y��{���ߗ�}�?a���hiE���U=�y>���|���UI�����i?j��t*	(������y����s0����Ԏ��U5O�S��elp)�_��;���A�^�׶s#c���_�)�}�N�� ��/�O	W�m/�hc�؞xtz�D^��E��=���G��yh�-/�hr��0uω�=�Ebq�ۺ�X90hzd^)��hq��`�MC��x7r��qM�Z��[�#�s�;q�L�fp�4�!��V����l{j�ڜ���@f��U܁,��*�y��jj���	[����u�j5�0OGP��琍=PyY��#C+{;	��P���Sq�������j����:��"f��]�mAY�ßJ蝟/�ޜ��G�)h��~ a�`\�Լ�s�A{<��d��\�u��ay>�g.ig�C�:3�y�>��4�h���^�?7��|����}��ԙc	������JA}�/^w�xa9�����Ŵ�A���nnJ��w�;��������f�H	=�����1��#����.s� ������L��_����Y_�����,�07����2��S�Wmc�aW ��b�!����#VU����^u����j�ά\qZ��F�>çh񮔍8;�@J���b콕g6����o���-�/5U�Ւ%���-�t�%���M���������ݭ6f��2$W>��%�K�����M�(�<˾⸝�j]p�F�Lv�i�]���-���VP�b}Bj�f��N��׷N���L�0�85��[�C-�~* �l�􊥛����{]L%�B$�HJ8�Y�ah��d��{ٻ��M�����l��]jGo���(���5��9]}5��{��K�(�'��m�&���%WX��X�A�4�˒�˫�ճ�B�x��n���Qz�WT����T=�}�����a[�~�r^���^���ҧ��)uc�b�c�$�۶z�6�}Uǫ��yI��*f1u�(s� �u1��4�R�BgwU��W�-���o	ǎ�e]\�E)$�Kt<
�٤�i�W�S�W��xȮj�u�6�#�U�Y�X�mE�5MQ'p�bv�����-7/k&sa�ö�5�cf���٧G*ٻ�d���M^�|mr��`p���[x�8r�^'+/3�#���5�a���wh�r`딺n2�ɴ����!�k�r��"fVaw�L<)!�����8ՂH>7;�]�аC�)�L��R���6�\*�	�]Wv�s��xN�1��Ϟ�+$��.dk���᳏�C�y����!'[�]�l����Eٸ�Uw����f�X/��%�x,h��Z`��E�E�<��B��.q�x4 ��.��Ho.�H�.t�ͬK�9�9>{Y7���8-m�7o��oV��]a��v\v���}�m���U��DZ]3��Әis:)�tP��Zc����+c�}�s]��֣��*,̢�)���t��
ӧxYU;8.���y�q�f�������}-=��Q�枋���p(BtY�i<�B��E��|��ѪYͶ�#F���5�"G���M{�z��[�n5=�24]<�����������˽�u�(M�H�qh��MԲ���7�q��me�ߒ�ʳ��tlsr�_J�	d{x�����Z�$`0�Z��������	่���"8Z�t����ݔ-�zh�mk��E�7��w�Jv�XY�y�,� 8�ܜ�x����Q�����z��Ә��� do��"�N�d���j�1-�e��l�.��N��{�U"yka���{�6`����B���Ơ˥W�k7(��
��)޸P�y�6�!;�q��]��d�3F�9�����^� �9tlcozr#DPh�o:�	��m�*)�HH^<}x����o�8���8����Ǐ<w�2�I$�%��ﹱ&�W#Fƀd����뷏�6�8��8����Ǐ;u�$I	.A<���5�=:1��`�A����㷎8�q��q�O��<x�ٲ,7IU@UT�P��	+���)5EIF�&�J�I)�4HBW����ж�e��W������Zοv��X�,_�ڏnk�QF��E��k��P�Ih����\�ع\�捹|W��_��Q=��Ebą�w���Q�;�Ih(�+��6�E�҈�4Q_�V�B{�6�F"���
H*���0n�畋 �O�#�d76�ΘWI���˽#j����v#��w���ӟ��}.v�����
1�r�Ĺ1S�����Q��}B��4
SCJ44�!�{�{�'���-6����X��{�Qx�Ͻ���w%��Q��.�ʇ*e̽k��֯���ؑ��[V�C_�.�F�O5?|���%H2rM�@�K�P�2s����\�fs��=�oh�qa�*I���a?ha�{�AN}�eoPwz��tu,p��B����\�o��\w���ڬ��о%��=00��ld�f�ݚ��ۇe���a��6���*i�ֽ�v��ZB��z��`x� �>w�`�"xjI3Z���!�k/���v7}�nOl�v+z�
&%=x�v:��Z"�P0-�>�;��:ݭ��K��}����ߞ4P3�@��xC�=F/���t��fY$�"�ʗ�n��P��H(.��N"�;;�6�M2������L� M�A�C�!>v��QU�6h�[�&Mxc�mT�!t�VMCδ{M�����b�l��Y��֩�|5B��'H��Bw+���ꂋ��g�A{�z�I�:�q>J*^7�6pJ�*�*=+\=����/P�<���	���t|��q"�V}�;��W���yA{�����Ȅ�M:����Pi�L��q,���C���]$,�m>�*;9�;�U]�l��V%�t�����O9�D�B�#�aa��m�T���۩.�埠���T��>ƱH������Ҝ^������S"���� ��ҍ0 �"(���x
]:T��v�� �D��� �����'�}�P���Ui�)YE�i#�}��8��/���Q&��U��7�:Q�ޥ����ix���X&PT�{���k�?=J�����t��=�~��>|�k�	��+`"��1L�t�&�2b�o�;���>����ŭsy���o�k�/(`�/~�'H��}=�6}��'���<���Sq��/��&c첶�s���}jw�����<��~i�۶dJ�s����/p�LI�]WyI�U>Q���͏�T9c�q-��<a��cH�#ZD<'��פ���{c5���G�5��a�;���z��~����i�V�=_r`ΐ�&0�zp���$i��qu�6�KK��ڣ��:qkR�2%�`�a�����{���UR2�Ű�p���s
ٍ��m����˻1��W��C�<�͞��^7�R�F>�%�ҌH�����bv�	����׃N ��k	��Q��򨏖Z���+�V�?�����}>� ����mt�i�M�ha�WUVAA#Ru�r�MnW;X��U�;ή�X=�U��q���4^yfY3�!���k�X=a�ts��ߨ��=��A�Y�E�=�I����B�Uңs��X�&�\������E�o�<<:�
��ЁM  W|߷�Sz��?JZKɔ��lwS')iB�2�s�H��Y�:r���n�=_�����)/�^x��P�z_S8}���yXC���N�%ڹ������W)�-��/BXł�������p{Č�4��ʹ�^��./'���$���V�1%N������"{�EvjB^;}t5U&`�ň-- !� =����{kr;-C쓋�߹�b4(Y��;��&�-��2b�u���&�Q��i&�Al����1�T��D;;����g>a<61����B�B�&�ю̅�<���8�o�f>�zǄ�;.����ȶ�m�thL�;`./�D���������r�;�=�t�u�u
���d�Ľv�#�:�y>~��+8��:��}B�o��)��(e1�S�y~�d���%?-��z�=-ot���M��s��[>����y�/�	Ŷ�l��!��Xv\�5�k��e&����]����lc��x��Dsw{}�E��-�N|�<��cϐ�m�0CXΕ��l�7�y�RD߸Zu�[�F���xtݜZF�3M� ��4�K�Ư��"�~_�?h�)�R����ݨ��"��۰�V�Kζ&Bf��j낌qpwA�n���F��*�[v��/g�������YO��/�떾D�糶�1��+_D��EP�u��{Hݦƞ��H"�xҾP�]�U�Ё���Jhi�UJ!�xz'�Q'�:{Fz�}�xnO@I�n���V羣�P�<|׼�_�|�!Ғ����c|v^��V�7�x.ϡ���k�z`Kn��j�g���'���} *� �걦TS+���9�ă$=A�A�;�s�xmk�y��k��[��"��6��}CaԽX���#x�/���	$
��E���|'1l^?�C��'����_1V_���û�Ҥ���Ҿ�tQPJ,py�~?Yւn���+7�Fm.'o^J�������k�K�ԡ�|����r�Όw>��0\&Qk���7s;��s=��Fߡ�>���#(nֳ3ZO����מ��R�9jw�D��k�hÞ��
�P�X9���A�[��W-��B�O�_
��5��@m��nty��\Ut��z:=.���&0cu[Wj��l#@^�������a�1k��5n	��Z��J���9�ϯvㅜ�u��|8�Շ5y��~X|e�8^7����~^���ȳ����yU���钣B�P�h��w}{�*s��ZȼC�����T�-��V��ٌGW,�S"ѢpIp_n�ց���2B���)J8^`sc�
���JT�7�����}�J7����E�d���7r���y��iF�����|���=���^��D�<<s ��W�bz���MKjp��Nڔ����y����-��󽂹�q�ӛcN�rb�[q��J~�vtzOy��%�9���l��+>>���r��S��F�ߺC�i�����c��؞@�5��u�� �S��]�D�`�g0g�O��V�]
��}]�[t>7H��e&���: �����n�x�3>�ń����A�����,|�%��-$��>Ցt��&��s
����P��]ϋ�e۩�0��M<����j���a��;��(�va�?1wڟ%矪T� ����Q���ڴ���e|͔K�3�[g��\�|��ZAT��9�����\!�:�v��$��xz�5������tr[Z������h�r�{���\ ��X��B7:�5Y��B��%}�Ǧ0��GtHv�h�v)�ۨ����A��~�w§ӹ���؜�B@���&:�6'�/
�C6���B��Ws���^�,�@O\K7'�c�e�h�a1\�QP�;�~J��hu�+��w�n|eI�)[.�i?3��<��rAY�0�wY���P�e�؁�u�D3Z��n�a�!d�QJ�(��}�ޠ���.I\*�3��(�#�^����0N���A��h˗27l|�;sD}�X劢w�z��������4+M�CG������Av�;ط���^a�=�T�m�`,��鞳$�9@A�P��S�PS�Q��V�6�j��kߦ�[l{��8����琏yTUj�}{��Q�I嬾�qj�.f�=���E���������Vhlv�P�H�>�
�μ0}5"�^���M���r��Kq�A�ye�T��p����0���3�z����q�Rmf�\�:�԰a��U6g>pu	Mh��ss{�:Es����5�cx��Ui��?��g��Lq����><�m�o���D���j)�>p��^9��q� �#ƀ��]�K�\VW���E.�u�?-���4�mxt!���VP�x���ρcٽ3ܘGo�E7[�b���z��$�N�ʩ���j��?\�=k�Bq���[a�m��GH�I���Y�O�5�sX��� ���m��C�Gqt�H&������Ǖ����?-�8�'u�}�,�2��7;��2�;�����2^eC���%����C��`��3��>���z�[^>�_,�<�05�v%J��}�UK�$��&ӁQ)��y�����l���-�]h��RZma�cJp���;�X-���9�Q��+f+�.��J7��281����|���u�Bĺ�J��9�.h�"�u[�[}q��o;[���J~���������{�6���}"�]繲eq���x�!�5�'N�T�^���W����4l����7�{h]�ԥ�5�k��	z�h&�|&Ƕ5��9��g���V_gB��_xL-ʄȖ퍒�	S����)=��+^�Y[�-
�R�P��JO�㍍����ӣ8p���0�Κaٷr*�Su g�m'��(ԣѯi������6��5���������xS�tHa}���>|���U����1�$���������sK�=SiC�g{�J�=�u�j���Q4���XXa��))�t��B�s���g��,�������s�ت�8�u�9s��E�~�L���Yff�j��O����)�0����O����N�]ε]w�M5�Y����4�"C^�'(F��Ô�#�6���b~��Ec�y�'�x�斛:!M�/y��9��b���O<Ǡ��^�i���{�~�7Wd�Թm��7�C��2)��;}�0�Uuf%y�>�)�QIxi����v����>,��>�B9�ў�^����80����S�R�I~'34�w�:^����<� �p���u���w/&��}�3��^��y��+յMC���L�D8����T� �WZ��brŘya�X�#U��g5�<-')rh���l���E0�2�OoЁ���일uS����P�89���d���:gIy�U�-��Ν&Pv�*0�Q(M3Sz�Pŀߘs�y�?�)��)������PJ����
�����4����w�+��jߦ9�
�H�>~�d�4ݲ���YN"�R�-���]~vk��k��������a��5����٣p�g*/�T��j�� ;�W����v�w�p���a��F'����ض+�c��� ��X��Ve���Ǩ6��(֑��^���<��g���a~&��!�%"s�N\u]�[��`s�k	�xm/RW���:޺r9�ZM�����s�G��w�#X�xk���y����v�H`���1�,���&�@3~�-�n{�Wa��W�>�ۨ��[�}˿{��<�7�� �� �"������}�-�����,6�ư���ʓ"#;2uC�^�2X�����h�2
��t��uTG����L��\&9�:�6+V_p����W�4�w��ui��!C(w�A�(�a�nQ���zC���	����L���>g/"�:� LO=ť(f�{����a��B'�tV����W�Y>�.�>��j.Uwy;{��Y[=��KQu���D� 7�[�b��_s��Q�ʎ\� D��\���&T����0�❛Z)�z���x�9]{# �2�<kP�zu�G}��=�N��%7���n����ϥ��44���Щ�pz�飏��o�b}Y!�:;_�ee}�>�r;�pi��,�W>�o
�ѷv�Br�q�����P'���+� +#�7Ю;�W�a��r�Wr�Ԓ���5�9�y��Y��WKgx�eu@5RO�cX`_	�T�b�(�a�u궟oG65Y���j��A�}�|ڡ}�	��<�Y�8�����6p�6"S�H����m�6���>!F���PZ!���C~]�@�]bz�
j��Ɇ���Fʿ���0[^����ݝ1m�w{���x���a1��=7k�=����B�>K"}�v_�f��lcgQ�W�Ḷ��IaƆ���c�6�m7@��d���^Es�% �w���ݦDR߸�����t�����EzmL�BS�n�FKnL}E7h��Q�0y�盛N<q���OU�17��s|��po6�@�e/%� biQ�"Ϗ���dڅ�h�s
9���s���I���!���y��|�y��~�9���<54��X�!�B��}�긧���lܛ�/�J^WRIr�K���>b]�9,��'1���za�<��eu%��Hֈ�F�F5ذ��؄�&������|�6TօoIV�)�}�z���^dd�-�sR:0�`ɠ�<���u�J�),gtѻ��ک�.K��NU놳��y��e����ߝ�O��4����?��͸�;��,>\g����XJVt����(|~�V�G���~�����r!�h���v��m\bO8���N^�t$����ₛ�j/lK��#���,a�^YnB8����(^�vf~�~��sRXkN�ua9�װ
�;A*|��> lP��&c|��U_}�~:���p~�����ór}��^��a��TO=��u��@��E2\����E�T�w���euB���8��$_U��Nϻc!!}V��c��c�c�������+��J�u<;�ٟbt��@���)�W�gP�~��+��Q�FRΨk1�?;wW:ͫ��EK]g�ܕ�"���d^9����p���H�>�
}M�����g�����l�ǃ�Z2-�׹����r�P�R���l����EC����Ϟ�,t,�����"=U�������z�����V�&`ك�s�z�q\��B��1P�V����V>��\7�~;�rLi"�n�[kߠWfϐh�5��AlLO?Z��<�����.�l�o����뮇���Tº{��4�3����1 ����ɷ�<����Y�C��X��\���j����{�d���Q(+�3=����[�:%^�$+E+��T��V�a�n1+��>ʰC�m��5&p��β�6T�IN�S�mvA6�����^�l;�I} ���4�:у7]������3QU���L[K���� ���,z�8�9�7Kc�us0���x�eJSE�h�6���a����B�%��a��ˬAĦ���n��C:Q�?�r�jV��`�mtF^�VM���c���ovN�Y0�^����2�:��WEY�<}n�Q	���f2P]2��x5����}Z�iq��zw^n_KcIB��Ŕ2�kʄ����zupThx�+s�_�q��fnvm��hg��W}g�#.P�8�i٥G������X0�p�*=y���B-�f5�2�-�6J�:��%y�W]ZXe�k�Wz�_J��#JA�i��;A7]Љ��85Z�����(#�S�V�
�_#o!�^�8w�WF�tW{��m�1�`2�\U�sB����/�F��l]�����Z.�2���I��G��t�X��B�gm���6��..A�ΰ:�Yo�\����'r��F��x�s ����vt̺�d�L3WV^�`j������&U"P@�X����n�h��0����91Bk��TM
H�B!G�$�RT�]W����ܑ[�et3*�ɇ��s/)�V<�c6/�h'Y{9����d��½1!�;���ܺk��C�C�_2f�īJU�����usE�9��A��5֖x`�A�4���0*���Di��>@����A�Ims�3.�oQ�6��"�;4��W�l��yu}]u�3�uc/n�jN��b�Y�e�X�J�݂����3n������b�^���(+�f^2ݵ��i�5��_mc�ڠ��;���zB��R��m>m�A]�+�����s�L]����f�hwA��&�;T2*��4[���(Q׵��i&�*N�ʶ�CP$�#���j�;�9�o�)�S�V�2n�w49_S�bK4�H�u�S��P��I�8ȁRn��g�@��!�2�=[�m��o��sq�U�U��n�4�mo��Z�G%_�������k���[Ps��L�� վc^fn5S.��e�U��������xəUt��r�H_\3�����.惲ㅜ�b�c�Q����*�ƛ�2H�y��!�ب7�����f�Nͧ5s���A]��T�0�Z&uκV���]H5=k���9x񸃭��u�6�a!��Ju��ad�'q�N����'%�%jkp�~"�w&��n�i�6
h,Q�5s��{�{�{x���N8�_�q��׏<v�7+I���s.c�o��ch����W(��z����ݼ|q�N8�_\q��_^?7��z���]C�nQ�b���j��w���+߾�*(����� H�HHȧ>�>6���8��z��6��Ǐ7���K����%cL�Wƹ��mȈ�Rl���Kh��j�d�}6�[�\��o����bM�Š,���lcF�m����\"�[Ź^���x�X�E6��\�%D����	7ۄE��](���X�nj�F�`�^�\�+F���F�5O�^x�8U5�Dm�������Q`�\��b��[��F�cO:ܢ#a*1X��s`�H��!�� ,�#}l0j�E�Fa��&J�Xdڑ$���)Bچ��H�@���NBb� ��F�R������1���ȯ�t���a���ݻ����;eߘsl ���\���!�����u�(��$�Al:T	P���i�@��r6ȊH�>i�T��]U+p���!�~dY���	��a6�Q(�0B1��(��( �@�@�.M\@
��2J$FZd��uf������M44��򧓕�|��v�� ��8���u�0���Db>�X�z�� B���|ǎ}q��|�zOoHg>:�C�w��0��/$SǶ���3��8>�ㆺ���,[!ϛ�0��� ��Ǐ�k�P�\���)V9601��zhN��P�F�r�\b���@ה,t����!�o�ß��"9�8�4�Gh����V9�7N\r�Z�R�/���Z��*eC��q,��!�8?64��5��l��s��<P|����S�-�"��.�/^�n��	~�����o�/�����Iz�d��ҭ)�w���.~�1-�BdK) ��aD���;�'�~�
f�Ű޵�ş�6,tm�j�tS�� :�m�r������9_k���>�z	An�fou��7��qn�;=�1�{��G3�0���c��� �uTG�-n�����Ŝ��C�Z�.��Lp4�����D�]x�z���H�><��z�LhZC����O���)�/z�C`�Ѝf.}1Z�8�v�zI�v���i����魬p���/E�05��.lF��8R쇙��k:F�Q�2����՟ (�M�*Ne�'اip�e�*G�^�JvtӶ3��������ȮͶ6@^��#�d��[�BsV��9�ݩ|�y�9h=%[���r���ŝt�^��HO*]H^��N޵{�}�r��>��)��ha@��3�r����6:ߺ|�u�"�ݿW0�%r�������UR�33�>������g���=������R����{hw�W����Lh\���͛�{g��S.����їU��9�) |X��\�"��#��%q�������z��^TO?r�o
�n���)�Yz�@�*���V��D���.������=_d���hȂ,��f%�t��D�d?5H��Tv��9��Ъ�_1a�VWT�& ����#���
]�b�fU��+�N����y1/��=5���E6P��涸9"Aȸ~���[TwH�r��jL���[5�b����ѩƩ�\�Ds.�t�d�bz|�>���à?����lf��b�w"rX�k�A�z�G=sy�f��p(�o_AX����Fi���~vz��i\[AW^�a����k�����)��pȓq��R9���sϏށ*�ܢ�9��u���	��G��>`���S"u���-���Z��L�8��'��ރ�y�ޫ�W��NNuξԴy>����I��Fk�ꮌ��3W4��"���U�y���|�RW�-Z;ﹺ{���%��V��c�9���)v�Etb�-�X;��5m嚫�e��ofIRS�ŝV������7�y��q�Ǻ�O=ѯ 7{�7>C�؈(z�5"|�ł.���bK���=L.�i�MI+rEQ��_���?H>o�-��R:��$����x�G�ط���X_�v�{����D�����]�RK�`O3L(���(- ''��	&S�Ҏ ��0��7:�mNv�,n2�p߬ڠK�}*��޲F�SW��,���g2}����ھ��b����=)�uXj��z���z�96�E:��=��R�)���j�r�XFjx�g��;[�����fq���~��N �!����V�ߠ`����*�}$2n������el��GC��k_����q���t���� X~�>��Ƕ��	[z)�zcv�Y��u��N/�Z�ܔ	bQ�gР㉸韗k��<�Ku���g��:��0�O{�يn�I�7������B��֘[_���>��L�-L�8Go��:T��~�+T����8�^����P�ύ^���1 O?w)�es������.п�]�{�l������B2���f�Ú����9dƳu̼�L)k^}ts/N��ȌPxR�<�*��n���#Po��':�dx�!��k�y�)a۹�N�W`�reF��ƭ^��������jF'j/;bGz��\݈�E���rT�z�W����^!����q�ŏ2��̚�ñ~��!������X��A�~��&�{��A�,�:����q�b��1�;�� `��v�ۈk��n˩-#r���P7'�`s]��2%�{$vgt�[DX,�f�Þ�ej���M7Ć0����3U����D� r����Ģ�חE�G1�����n`jyc�n�*��3�����Ü9�m��2�6<w���\�;׭.�҇Wvq����z�g�����`:lu�!���^O�J�
gX8H�!��s"�*!�O6u��=�%�,�[CbJqI��BOm}PX-�����LDy��N���F�Wt�s҈7�(��h�����1j��l'3Z��8�E�	�e� �>xY��1oO�=�9qx1�h/f�&�r�o���(-n���Q1)�v:�����`��sR�����i"�)c�P-�<�<��7�2y��VES�g�ʄ�V�d�(��W��u}9o=�l�@��b'�`to��g��N���=�V~AZ�����Ֆ<6��X�-�J^a�~�ۺ~k�����k�H� �s�T��o{2Ŕ��1�U��j��*^�!�|���x���=����RBφ�0k�\6V�����z�Ż�VzE�d���h�A�����9��l�_1ۻ)W*�ɭw�L)����y ����!����(x�}R��a��ʓ���V;J����Q��'n��y��;�i�����d�a�=Y_��1��~���yk���>�XZEw���wr���f�A<�L-u#�;Zw��j#�-�T�j����nP�)Z��6q���2׆{��CX����8A�j�ԧ�n�^�ݹnO�7��]�dsuèW<r�^�ȷ�xm��2(�p�-6.-��t[kk�D*7�j��Ǳ�#LO?.�ār����4�hgdz"��fNg`5DO�ͮ��e�T�Q@b�UԆ�&�S�'g�-L��)��&�K6:6L��+i]�����m����9�.(=�eN�Pbк�����8n.�=�x�-{�\�v�gZZ�zS��uO2����s�{z����@�4�����C��F9���*]k�ѫ�|ޜJ/x)��A�&\���9e�X��r�ϭM!g�����P�a�k��z�3���?N�nb�*f6"��4���~>��
���}֩�j�U�M�z�dҞ��n@@oE�]�TKp��3v��,����9�$�}�M"w�C>���P��=��
��7y[A98����5��y:�Ϯ�י�A[�C?e>����F�V}��or�y��rŞͻW]f(�/�}�C���A�լ�ӦN��ِѳȭͨ�pS����ڎ�=ajS=[S3�s�E�+~g�J޳&�g
'�m������O��}˸�aP5��|��<ö�4�͖�F)��O��/϶�N�Cr�����s�P٨f6�&�!���d8:�c���7��Ϋ��\�	\���6��X�;M��s��r&l�3G��ĳ�\7�����h$p���i��~u�ȱ������婢�X��وH��-2X;vu�ޠ����j�z�R�n��p�8@��!p[a�ancآq���Ծ�Ymv�c�z�>{�T"�O��O�9T�(s�R�x蝹KL�ee�����W���v���&�����0����בOM{�Yt�t��-�h͋��q���}���Up�th��@�Q�݂�cX���ǦLX����H#<��}��3/E��Y�Y����Xq���C�ޭ��lxu��"�c��~�=J�cz5���5��PJ�TZ��Do&:�;���W�X���.겺��W�Ǔ�B?���h#N[�?�4c&8�:���Lu�<'�;�Suwus[_��5엇�1���DwO��.з���*�f��=�ag��&kG�)�k#�NNN�{]�ޚG�r��x��6�T�=�s2ܗn�w���x�~X��	�,��n4�1:\��]�o�'k�V:��N���o���l���;�W�b���xXPk������ii���@���~zk>s��'~�^C�gҫ�MW=Ϯ��r�����X���L��Ž:�X<^6�W�+������,���bt?�{�A}��[n9n��T_9���V�:A�3L0�ы:��z%s���~|_��A]7��F���u�-���(�v�ϕ��]Г��V�<5R�1~�C�[[�=ć�I�҈}�ބ?j�5㽯�����rr����y7P:7�\��R�er\o�î}
�FV�H<Dw����}�q�\�{���ͬT/������!��^ZƮ5� ��x���x��{=Z��y`Ƅ;0��6y�|DsSH����.�9T���Z퓧9�Ѹ��W86��0���J�O��M!=q;�-4Bgf�8E`V�szhox��q^��+`6�e $o�1)�v,��Qz׶s��{���Gt��7t!0�I}�T�4 ����ZDLjz�kN���thEn�O]���h�%:!�.2�3ٻ}�wg��^�-=��V��ΐD�1S��O�[�e�/���*��}�4�}qg��Xg����?�m�SX��+i�}ٷ!�O;������睂P�0q��[�Ȅz�0��X�A׹b�����K;����c}�,�D��^�ܳ,%�{��<��R�<!�k(��u�����_^�n��]]s�X�n�\��<�a��lI
�I;���ӱ�^;<�(��j���������jݺ!��4.m�^�<�̙K�o�,=�-�� ^���IN3ꃎ$\�C���/�)���*�:����i��9�������a�����up�����<�cx�UΡ]bz�
j�ܜj5>��x�	�u���=M�o:��7N�c�]1������mf��Y�9���ܤr�L�qo�L6ޚ9���u�!�3R�0Mǹ7���q|��/X|��+��hH&��^m������۠���r>Vt�iÄ=��fT����xpQ�0���װ<�kζi�s*o��]uye�$�������c��(w�Pz{Ҽ��ji[G9�ṎZ�&�W7�gI��5�+�0s���I咨I�wBe��9�2<RB��d/O�<ϵ�:��b�%�]���u�=�w�Y])��},]�|"�V:bXA��Xy\a�	3��Pf�hu�P�mB�z[{��"����Jq���,�[!��|�ے��� Gf��]"?b�!{��9Y+�uQI�]u�j����V�{�
��t���h+L��@�P��̮�ͼ�m1�8Q�+�LfF0�ai�6�N�G��M��̨:�`Ӽ�M��9!����ٲ�aTd(��
�,�*�oT59�]�S�=γ�W��xx��{���xH(#��s5e�)����S��;�48_X"�j%��d��\:rt58�j��7��O�NY�<O�ãY�b{�fۨL`��l'3Z��H�Jq�:�	��rmO\�H��l�m~�V{ꀕ}$r4?�M��]�#'�R�x;��oR`K�z�.Ĺ'a<�9�����x-}�-�_O�O�0p�B�$_�����ϲ$��t_v�{�I�c��b�r$���!��z���Ɛ):L�c�:��\$<~򨀫T�v���8�Ԗo5�/�����ߥ�l$��_�	���.�-|g:�LL��� ��:�!�!r:�e�w��-V<0}�T�h��1�f��,�
�R���P�L"\u�G��M�X}�V&f��w9X4pv�0?���Bs��F4�d��6��h�����b��oɤj1��nن;'Jn��x$9C�pN���i.&|�S(ί ه�:�b����'��Gg���Ɏ�L�V����n�3�v0�2	���-4W�
V�Y��Ս��2�S����'J�(��&"z2�pٖ��/�Z���wJ`���{��z��L$e	��8����@kz��\`ve�2�?/��ʶ�.�����\�86zd���Ff�S	���+'������chٜ�k)ir�`p�<��V�� B=�ap:�/9C���s[�Ԙ{�_f�ފJ�C@���#�r�k����������6�`�)�)����<�a粰���u�Ǣ���S��<�)��;MJ:jw���9�NDs�|�6��h�	l,9u
U8°�:���Tg9k]ʽ�=*\��q- >��x��r�������=�(�Je�rig��1�9a���P�K�K�cƷT�����=;��>-��h��F�����~��28�h-��Þ�>���,	����	=��\��0�S(�T���<~��Df A�����[ԉ��D����ydvo�b}���긜�f=����FN��޹~�i)fl�I�3�
Ltu{�֒��c\9�Q,��&����y�:��Y��{Z�Q�-s2��u�g�g���'̶�W��O��d��v�O�/�p���8x��kR~���5�@���C~m�}��!�^����1|�S@M��Q5�u�2�Rٟ���0�������T[.�Z�sp_F��������V60�G��E��ʤ!^�%�Z�ǵPT<1�M���e�DMqθCN�W�Z�}��m$(�ʳ��z�%Iw{�Yt��o�-��=����3��(�5��5{��́RA��93�|B��[zv���C�k|�����ժ����]��M�b�U+p�'q/�G+�Ӻ��4~Ta��hc��Z��C"�P�	u���1�Ve��Y��u�)գ���wuX}�<�RWJ��w.�+���V}��ml�O�e�U�{GQA�}q�^�s,]0��S�4�7}����W-6���1sщ=��tYy5>�J�)+J0�p��$�P�gS�EL�T,rL�}��y�n$ÎF����]���:�������cд�]Mq�i�w-���)&�}Q�."��018����[A�{z��H�p���3voL��{��ڙ��ͭ�搇:�:��Aڃ����4�U�<Ǹwg/',^n��5,z�ʘd��»Ρ�:X�gJ�E�6MPd��G�X�-�f��L��cqir�61�ݫ���e��vWB$a�4zImnw' �jt���Z2��>�k����O��̓ڜD��.9�mÊ�����]��^��c5J��r��Lv>I]�o7M<bh�Vs�Bſ-��48���أ|�.��3;�m���Xu*�/��u1]�ǘ��x:�_n2��Ƚ��/����l��ai��U#2%��s~�.w[�nF����w�t�%�$���z8XeN��d�i��]L+}�m�Ul[>%�
j#3ʊ6EP�T�G)���T4�!ո��'�4�H��]T"Z���sz�|Q�a������>'xus��٘Ab꾒��ϙ�u�
�\Ђ�׹!��.2���3��У!7�M�2�P9o$f��d{'��yԶ��t�_.Q�v9,��0uo9u�b�`���[��M;��i��
b	��J),T�l�e��u�Fʕظ�e�G3��ӆ���hqݷ���.�I�U�Ӆt�¥;{b�e�O�/�3C-������3��B�����Y��3�oAw}���[ݚ�T��Asj-�asQ6Wkns��}�:��v;GI�<�+�n����Ȑ_�?��g졘���K��@6[/�c��*�Hi��'ў��^V�Go���

�<t=�&��J��Ɛ��׵��Z�BcpQq	�݈�+LT\�O9�p*�o.��8��s�6ew���hi�iұ2�\V��A@*#�&o���j�8�v%�zf��Po_F����������Zw�
�9N�z����R�&�\�^Nͭ���2�.	m5�(�ؘyX��������q0�u8�۾�r�s���T|���F��4��F�W������AcWw�]7(T�RMQ��x9��U�&�m������8d��z"y�K*Ѭ�r�\�I��sI�y��8œ��ʛ|u,|�]PڙX����&�)������+
hNw\1�	d�Gx`u�g�睕���$���#��j*"�sm�~����0$���t�ǭ�||}}qێ8���4��Ǐ:@�dT�E� �lZ*+���nh�22#"�!����ݼq�v�=z��>���ǎ�^�Sp*H�%�/λ�۔sslc�7-�c"�o���o������q�8�ׯ�8��׏<u�������ەF,b�] �ԅ�P]ݱ�λ��lEGwm���#^ZWIK�^���s�o��r���E;���.+����6����b1��D������l[�ίsw.�G0��_�̢��+�1]۫�s�F��~����n�$D*�D�5TH�W!뫚/�:�S��%ݫ����c^.L�wh�s�ݷ^uzW�3�s\��׏&�7�#����Vֶ\�5����dL�{Xf�u©ʙzx֬��J{���n�I;�'x�P��ũ���ѷ!9���~^���W{���W���}K
����8��a�9�NO�z1�*�ϟy	�Fx72�\����V�Д��,~)��^b�Ui�B�+�1r�!�.����܍cl&���R*�L��u��u�܂C����U�ޔ|����y�y_VO;y�������RWlՆ�m���I�O���9�{��~\�)��������d��/�c� (̩���n��Y�-D�I5�{;#ֽ�f����u�2�dW?���X���q=�ǝJ�4<D\��jx���;��Dz5���}f�E{�����1�qzE��7H-�Z�I��u��9W���jTë" ���8"%�y�@2ňxnׯI�m�������H��t��p^�(�19����1�É|=�(��+(�;�r7��kǽ ���۱�Z�e��xA�����/�m�C�w�.;�OsՅs�UR3^��/>�w����i�a���oR���ڴTSW&��NӺv�j�X*�Yk�F}T�t�9m�1�R;��/ʇ�����
z���Q
�-^ޔ5�����<[z��1�NL�3���ˈV!
��ۑ�JK������X�[�Z�ž���,����ԝ�n��:���r8&�*�³'�V�i��7s����w�5��
����
�߻㴍R���^_�H�<5��1X�1��s4M �%E�9d��,C�gg�F����B�K&��=����F9�:��C�q͋�Ccгj�bS׊�b�P�=��U^[>�ȶ�<�����F�Yt٪����{�%��f�~08�>�/m��y�5M/�)=w@��I��n�O���,�yۓ����f����x;'��[�L>�忥(}K�C�y�o.<@��[ѓ���{�}h+��R'�|��}ch�L@~U��cXv��Cݽ0��F�4�f���[$��n���׭�О� K*	�t罐4a��K��B�;B'�"qƌ�_L�Z���8+;���'~����Æ\8���W�ߧJ�g������Cܷg�S[�e�=.��ʛ}79�v#���u�USK����bi���{��cn]�~�2�)�p�ڶ*�	ܦ����u��L��~U{�S?1XP�� ��^S��e������@נ&��SȮsZ���7��;������xUk�]�D2�(��6 �>��F`ܩ<�`�V�O�!�|aW/ 9�i�A3s�wz֮��fwtU����w$��k���7|w-ph��8����"��j�z�;�6pgKzÚa5��V�=��IzZ&����}�e���	g.��P��b*��]�_sJ8*<n�p�߫�¼<+��٣�%������l6�}6X� >WX�W�e�X0Ǚ�eK���ّ��tt�?X��6���RW�\K�׃�h���^��1�R$��{3��3��qǲ�V�a�}=�-V��O�k�2�5��HO�Ƹ�	�y˚���{r����{=_Z�꒡�ٙ�뮛���D����
�g��c��v<��F15�V��A�;�4�{ýȃ�G�8)�m�k��&Y�����RFx����'���,$-�֠^ب��Nb9��>�{�:ġc�/t�6I�eD�ӹ�@ߓ��{*}!��J�n���4�2����g��Y�4l�c��sߚ,h~!����d�ёh�u�WH�O�9~+��ni�(��)3��Oˠn������^%��+�gP5<����v}�d�.�����]n�1\��� ��J!�b�	�u���Q3����C~���P���y!D�F��s�/7���<x�}�e�V���{��P�k�#�n�����C=X��
�!�0��w7�+{�g�V�%�lԊl��n��C*`M�U�k���8�E�P�fs�oY�^f�������f�9��y��X#:'��w:�Ω��.�emq�WoL����\�C���r"��7D��n^1[�$��O-�����us��Y[�rD�j��cw�����䷙C�0�Rbݴ����<�oyּ�PBR�Tс��M�Bm7E�h��>g��ѓ�CK5�y���<�<��
�c���Z&r(�!�/�K�ʭ3F�7�S���7}>�O}A���b��>�4��s�ޭc������s}Ga��#���\w����P
��C�dܮ1���p|i��]�[^�+i�3g��Axk�s��%�=��)�������0+����|@ߧ�;F�F�̆�[R�4����[5N �tjy������<��ئ�� �
:�v�n��8tff�ƨsk�����ޚ�eXdO\v�ӊL�O\��v`ҙt,y�/x����{F����>�y��)��<����G�x/�;�,Pu0��U��o��0�	z�Ҷ"z��_a�gGP��w�~h�L��o��r���l�ݱ�X`'���t$�OS�e����b���a�x .fcu#��ȶ�S�+�[$��Q���[S��1��[�T�c�f�uJ��{���}���}�G����ӊ��J�PX�`��%sĎ���K`$xs� ��b�cZ��W��IOr:2��+���N�f� Qj��gM�d�b�Gg
�0��߮��>�f�a��φ04v�\�GW>t8�.���n��e�K�6�\8�Vԥ�WpD����,&V1|��έ�(F�;{GL�Kܽ��\lS5{���<�`��w҇���n�U;��^=-:Z���1�ōv�p!߃��'�yǺ���0�mU�ޗ�]Y!���k݄��S@S{	ӂ/�;�� [����ս��%v�ڨpv�O��w�?1/6�ٓ�thF�&9T�5Awy���Z�}��,��Ѽ>���넉��J�:�X﫶&=�������,����	�f�\�_��)tj�O*t�\G���<��gq����)'��,�aw�Z����{{��	��罡^��A�������z�����O����"���V���@���A�#ߏq{�9�B�^+�U﹇v���μ����AqXbX������������)J�pu�<�g�|�4(�(�J��:�����e^��	�8��	�=��O����]�\��n r.���D�י�z�9�Y�zIFm%�C������<����)���{�A�^�s�Q�u����,RQ���+.�*��̳_n��^~P���c��&�rp\�+���nO�*/�������jۀ~��Ͳ�m�9����.������"{���/]�w���
�	� �gT���3{+�u�(U�� =�6<�d� Ŏ�f�'����x)�Gc����w$���U�5��S��U�Rl�i�73r9J���W��xxW�e��6����]��a��{a���yt��->⩮W2BA�q�T�w4cn��o5vFV�k�4� 9����a�r�j������Å^�6��{��$����i��V�%�{1_����{�=�+7�=���z�ϵPeq�C�J� K�����j�����YB��d�>箉Y�^'[�����z_}��W��R<��A^�����kq:���tYN(v43�eoޗn|��������l�m� S@ݤ���ބ|hyX,��8oF͹r�}�����e�c'��-=1�=��Q�I;�F��X�{L;��܋X%��G'���/�J�M��-���q{�p���W���Ϝu���9��_g�hW(Nq��,�ݞ���`jk$�]^|xñ<<�6�i�� 'Ps�d�ݐ9;�?��b�٣j3jkduC�.AU�ĸ�82j�(5w)"�m��g·/N�@��^�=��)�!�&]�$��N�1�6ц[U�pcn(�F��ע��C�9�ˇG���To��"1i̽��.�Ye�suX�+[|��j❽���F�,fзp�n@efb�k5��n���r������+��t��*U'�|x�wx48��o�(�c�^�g�񺲅�����hރ�_W��{�>5�|'սdaIX`�a5��˟�of(2��7��C�jCMb�0��/�9�x���g&��a�J}����W��>8-ac�>�cx�{]�B���&Է'��<�[T�E��n�Sɟ�����i��[�#������%��"y��H�)�=�x�w\����^���;�v_�������L��]�p[O����s \&����9�]aONfl�kB� �sv��Чس^�0J�22��0tu���}�~{ ��ͬ�gQ*/�w��R����~��� �5A��Z������<��_�u�71ޜ����A��n�CӬ#��j��l1��N��J�����L���pq������Ʌ�!.k�/{������_�����'$��Ja����S޺������
ܭ��uA������ŗ��Å��L�Ƶ�"��D�p�3��t$��:��[Q��:)%}�:5��ӣ#S:���:�; 0��f�Κ�>'���"��M�� ��k^ʇ�N�D[\J6/%S^X\�(<p��kU�Pg\��'p�����`r�Z'ڨ�S=�����cj&�ױ<�kַ�3��9fNk+Q��Po�I�w-���^o��o͌�/#x��H[Α�w>�rJ��"�����=��mS{МQ��R�����iN
K�7�G�yW��b�n]����ۥ[��ː��n<��wp�y���=�=ݝ
��Yv���;"��P6Ql��=#!��߂q�C�yy��bn1��J]πf�z��r ����Z&�F����4� {����`�	�gqoìO}Au֏m'�$����)����/|����M?*�m��InU����UÚ���k��í�5A&9�8��À���&7ٕr���R)�b�׮C"]�,p�l�ݲQ%�M�M3a���zO,�Sp��Zc}K�����G5ߑ�n�Ρ\�Y	�;Ut������c+���j6Q��3�F��;����y�[f�N�����	��L�}��N��zz!�����wk����JҀ��Տ?'�{�sg��^�.�<wU�tTm�T�5����xj��}��%�=�n����� ��u�9N�68�c�\o�a͛�I1K��6��)�`U9��b��=@O'�mtg���6�����@�4��n���Ħ+�����Bn��[��%P���N)2�����k�ЙP� (r�8�ep~.�Y��`�� q˧��2�&B��pH�=�]����p]K��.�u8��As��-E�x�G��Z���9��p�"ū�v��}�.�r�[c&ģvË&�V-�K�[@k%��fu�|:���S{�L�]Ԩ߫��<�a�Z-����zg�ϼ*�h����}#ZD<'����8֭�SB�%ԥ�_v�E�o��O��ۣ���T`�WR��L�︩&�a���=���_�����d���\|�F�/�s��w�Y��8��_i��̪ e�b�l��Hptj���<^+>H�SW���26�nn��V�e�Oϧ�я�Ai�ۃL���϶:�@�uvx�U���ɴ���Ý�r�͵���Ax���Oy�J}�ʜ�wlgw�pr�
#9ܻ=R���U��zl"\tI�Ǳ/�Ud/e�͎q��zP�7�"�`�����2k�4���,���ၢYDXׅ�ς^��dzjL���L$r�!Z������Q]=�f���7��u����3��
`X�,����K}�?/�����=����(Y��-�EV�M+m�s���ugû�AVl�Xh���)&�,��W���zz=>p����^0�o���1�4���W���P����ޭa��m��9���4F.�f������>�!CɭO�2�vٮѬ3oN��C�[�!�a]�=�n����
vV,��k��m7F�d�M�X��quW�U�v�a���mgi�n�i;:Ӧd�K��o�9hk���Sۘ����nZ�j� �1�:'��^p�~����@U�n�\g���[��< �@F%��׽(���O,�g}ׅ5+��g�b�{"�Ԗɛ�c7��[*0�VG	rrT����q���^�JAm>^s�aM�c�X��Y1���ٻ�^@tcΆ�o`I1��~*��*R�5�l丈��P�]�k�z��/'�@~dF��u���@���^b�w�m���}K)����wQ��%���4�Gk�^}�����Kr2sV���2���D�u~w����C�����`?gO���5��e
nOjU�:J������g�b��.�{�iW*��l�C6Z]��~w��oa`1���{�E���D� i�ۣ͐}�-�٨�V�E���he3"�Wz��u��n�m+2��F<�|����f:�ш��J-�A���g9��z�����3c�4|���گν��v㢣�aOD�lD:Ӊ�n����8���L��7�&S̔��u[�s��`���4R���Z^S�/"7�]^֥��VQW8�b���QzU�'��0uuս��[̘��  	5^3s���E̝�V�o�E�ň�ͽ���W�_^��!<,i��խAaNWs�U�f⊆�=��pʙ,ǀ��u3�j�t�M�Aꏒc�hT��==�Z����}s�	Z����PဒX͇�_<�v�yhjj�3g]�O�wI��7�TV��Zi��RS��v�hY|��c@7{�����Ѷ���a��f�mv�o^�	M{CFgjOqsL�4�6���dZ�h����^Kaoy��9�W:[�問iJ{�,��E@���ܫqs�r�{�����i�%��Ŵ������QD�s�mE��vL�ޮ[][��{�;��т�[�t�{b�p@�N�6�:b���&�d�Ϻ�d�pC,[>�P��J�o��g��37E�X����{�*m���3qU�3nV�M��.᜴5yC^�]�IP[�u�b��ܞ�@�Rb�U�S+��nH�6���+��I��Nq�\�_nLN�
��պ�J�r!x^�o�sl�ov��`}����R�َ�d�D�WA��2�CЪIݛ��}M�Ձ�*���!J:;�yẪ"�Ȥ	 �V4ԯ*�i��?(��Cx���>����M��$W��J�z�[J��4 (e+�*����4yj��dq,�e8 ڡ�i�Q-M�����-z�)�F��6C������יi�sht�x]���hHw:Vc�h�+�9n�V��C�7O6m!G�Ğ��GK�F�N����gQ�S�����7��*��=ĵ�G��nY
���]�zҷ]��^�јw���i���R��S�g��iޜs��s�ǳ4� x���:f�`�J���r�F��khuiN�5�V������[��ũ�6c��鮾mt���2%!O�Nwtq�r+�{+�e�����g���^�+��2�m��wVu�9�Y*Y]:��n�8j����ͫ����t��r�z�qf��7��x`M�G��&m��e�V�+�5k��6��u�]�Ʀ�x����Ik�Qq�&r뛻�dhY��t��^\;%u�l�"�mhZ��V�ge������hj�C0��
5SOt�1�g��ש��_;��S,͔��N�*���Z�㸜�Î%�j�FT���E������NZV[��D�,�n���Ǡԛ��(��-yɹ.6yU�y�����N�ӝN���=Lb䮯K�ua�/j!
�.��\�1⃟V���u��Seo,���6�ŗ��w��E9�n[R�3&]�-]�7�����>'���tH@��H��:x��;x���x�^�~��ݻ}uq� ���[��wc�ʫ�͹��5_^��i���qǎ8������۷o��o���R� �.,�n,�Q=}|v��o�q�|q�ׯ���nݾ�z�� �X�ђ���m���9�͂��ъ"ܯƼG��R�5A����B;�Z}{�s���g^�~����\-���]��*Wv���Q�O�m�μ�z^�o��P�*&�H6ĽPTm�;�zr�lZ*7�o<��E�N|^��:[���Ƣ�k�v��6����m��La��$�1��$�����"D�NZ��J8�iB���$	!O��"m��sr�f^�k���qXڏ��]�����޾��m�ٸ:�j�gV�Fմ6��r�:��Na��D圧�=i�%�*%�
(��E4�_Z�RB:tId(UB�MH��!H	`���0P@��J0�rE"�Aq"b)Drq4(��eэ��*��Ȃ)BĐ@�H�_H�MO�H�������p�q�t�6^+�se
s&��UENpW�Mӊ�����SS��9W2:0�{	h �Q�o��@t~�{x��TU�cffY{iE:׌���ꅔ]	9{��X�Wg�[�����p���Fg*Y=�k����^��k�E�@��$.�!-��W];�}J���އw��S�9cVn9Æklwz׆m�{�@�@�P�%�����:���U�^�a�+��,�Ld�@w�(xz�k2�������}
��zԪ�{=V�Q��qN�mtk�+6ٷ�i�g:�X]
:�;���u<t��Ou��s+�f�"[gifT�70�5ӹo��"�u>�ղCQ�~�_M�	��Z��c[�y=���V2tL��������r2(�5��|D��l�[�1��ݝ������X+�l��v��ɐ���0S|C{�B}��l�`�iljF宓kaR�����L�����3������;������.�[bOU>U��\�Jx��^<���m]�`����c����|��y\��>SF��^�N�r�{�c�¨q�r�k����3#G�w3�\���ΐ�x;��pj !�E������{��bV޾��d��U��|<�a���q���ӫ�t��񨄝�Q=������ݐ��|U6c��å��D�>R��<Â�fA��>����=*�#���O!�`6g]E{L}�> G���{g8	��H�r���T�p~p�9�p�ä@�*�IR7+�����+u�D2Z�Det��Fj[��w*��8 ���x�.e
��f�6���͔�6����r�)W�>���#5c�-�p�9n���K��"ȱo����h)lK�/��|��H�R�X*u�̋,�
l�L�$cf71�4o�r��������ծ�Ճ���}>M���l�mq*��{26��qkL;<	2]���Ft=�����ez�|��0	b�l�uk��D�нu��4�H�d3�V59����aB&����D� ����_�3��\���%����j=n���l���"���S.��v��g]���S��Ph�+�y��ͪ��k�ꅩ���`U�M�ٚ�����JΪ�kQ�2M
P��X�O0qQ�\w���!���/����.}��$��A�b5�L����˓ú�;z+3
�u���~�T��SCA�%.
���v�xgr4��[�g���">˶9D9E���{��jϩ*����漝N�e�hAo@۞H\{eHI.��l���p5�Ⴄ�)麛o3$�bҎ,�__G���{��=ǧ��óvA�5�LiP�����w���)4���v��徟M�F��UrW�䧊~(��Q�F}�m�� �h~>Ђ���B�24";�'ē���5r��Nm���L�U[T��}&nvQ�3Ks��O�1�L�Xv�|������w��ߟ�զ\[5�E��j'L�Tf#�C7�Ƴ<�ׂ�J����3�n/B|��n�'�;Γ��5k����������m,�y����A����UDf���fw�� ]@���"��[� L�,��q��Eޠ�5��^M�6<�YĪ��j��sط���S!m�O��ǩ�\�v��B��[y�m�b�#,��m�w�j�{ݑ��-986��w���xIy�s =֩^�t��| ����:�
�ePOCިw�������aA��#�yJ���g^szq�ޓb����������H��7�{�?�{>8��\�[���4`���O7
�MI�����s�;z�zp�����X����q�X��c%��B�T��r�MS���)�A�F���,��5R���syp<��k�[�e���{��O�?&��ouג��L���6�(�v�N�Դm^�=]
R7�R9�.i���M�m��[�ve��g.�$��C����nF��H�t�垪s$_[�[8�)sP�Lq�'%N��N[�ǧ4o��\��=A.���3@[J�U]X�>�s��p��u?��" ��~ 4x���7�	���w9~*�^S���Y`�	O;UWyZ�s;��h�}����ݧQ=��OIwgm�j����Z߶��4a��6y�x��l�;>%��n���~�/��D8g�}�Pzl��BD�ު�H{RQ4W���=�.X��>��>H�0`��o�L���=�
���ޔ�ҶL�ܬ
����y�X똊2�xD���Qf�p��c)�f <ϼ(��=҉��#y�k	CC��4̋K��G���}2��S���^�݈��b��Tw�)���)Mh��<�����Z�������U�׳<��8�DL�
k�����N|����^p1Q�kP�	��s9^��>�P���v�<*��l����^5�n���C'��["��0[c{h��	T�������M�^�f�U��2���"�B�q\D��"=�w�<�e"��=X�I|}�P�1l����<9�pn��w/`��JA�[�2sy>��#7�3 �?r��0J��� -a/��f<��""Y���Y᧡�Ks�ڮb����tR�H j- �_�Y��aD�=�*ڊ�E�������+;�ˇWZ��~��mq�*�zߧ�Hffg���2�;��u1�U+)槨���Xk=ֽc�R�$����D��YF��7��ռ�n�\r�[��P�ZZ�5�j�c6�4u%�Ξ1�i�a
D���q��7sW�����u4�os�u�b*|DWLy��7���3̔�A��晇���j�Y;G<�:�遏-�K�n���o�}7סp�v�hj 3���g���.��Y���1u\P|Ͻ��Q��e�ݭ��
�`�;;N�>����g>�.��u���>�Ⱅ��2�<�e�1�Δ���U�� ]�~�
����o�M�l^U8]>���W�6.��P�E��-b����;w> -�+k2�R{2wW�wwoGor>T�ו6[䁺�d:�c_�CYz�Oڐ�I(�fl.����˨��I�CUqV�~�Ɵ�hr�-�c�b���{0�v��:,H��{�.���!N�꣈�)�л<J)��3�l0Ƿf+�x��I;iag�S�J��b��«վK����unʰ7����坤��g+H��3��������`��gL�
G{4Mv�B~��7��7F΄e��j��(�9�!���~�5G��ޝ���:g2��C��n�х�{^���x�)
�Y��4�h@\1��0��K`��T�'k�ws;�E8�)�Z����V�L �;E�ܩ�L,uV�MYu�����8Eq���.��u�]��rn��j�w�ȾC�5�:0��b7��$�ͻͤ����Y��"�+��-H�)+J+m]��	�Y�v�uE��Emn�K�7�Bv�?��JɎZ]�6ް/���ζ��ʕr@̾9�)���z�c6�y:4۹,'���y�����{Ώ{��Kq�iё~0V��n��O�]�|bEj�2D���/->Z���=��sGse9�C���a�({�49���@Ui	T�}�U��u{m&���F�A�n��gdK�,%�Q���PY�7Z��G^�h���-��:��`�onw��4!-�ۺ�u4�,�6�ɹҏ�c�?�x�v̩�����MZ�ͬ[F�1��ܚ绩���qL���X����c"�ĤK�MgoGj�0��D�y͙�]?H��{�?�:w6�P����Cl��R!�Eo��.�f�E_�R׳66�A��g3 7��6UM3g$�9����7�ɝ[6c��[3��{䗿9���g�o�}5j�`]С	�����Mm����N뜝��W밗(q�r⺤�TGfQL�ѷ$��oL�����4�s��":�;72��;Z$�M9r�}�Mʀ�_a�.օ��p��
��]��7sK�-f���A�c>կ.�v�����@-3Jzg�uP��]}��,�
z�O˾��&���{�7*h�T�t�5�ՙ��l�R	��ce����o7���IKҬ J��q��*��pfn@�푾d
0�8�a�����WRN;Qk��������5y#F��m�0��Ajؘu��xLx9����|���0��)��-ƅ�Es\Vr�.gi�n��2h7.�����W1]/w��]����v���Y�v�{F�R<��P5��&GBw&&��f��x�>��_�! :a�wTR�S�����e�{���s�Vg��S���|�_Yzm{q)�Tvx�>�П�*��	0dU<�C�1vfq4uok��X;6���2�P�Zٵ�-�6@j
�X�~�{��1Ai��W̮u�G������+�$i��ve\��@���ŏO=q;�R��Ƿ���ޮ�03:���3�i.��B{�Gmܝ��K�X���\[L��@X�S�՚"��q�PK��˻��r��~���R���[e���IPuQJʤ�&`���<AM���U7�G+�����=J�O���7��j���chli�WN:Ÿ^T7}�K{�My(1�5�c�\�{h�vw8�s972U�{�'��:nA%*y��ʉ�O~�������:����/��TVsK6�d�hR����U�]d�=��P�m��7"�j�����c��F͞y�����K0k��ffu#�ϗg����7u��(V�9[��;Ki4�Z���B��xJ���6�u�B��Qb��Olֈv�p�rߕ��'����V���I��X�kᜆ�~���\��bo�f�z���gb�wA�ϸ��W�x�d��{wݗ������|�8\��ǈ`���BS���1���Ev��U�-Y�1l���0�ŷV4n��p;��L��S��Kof���� l�Ǻ���y��M�=^r�Pk@W��|�=bN;2���n���)YL�~��^,W5��N��b��fH~�lЙƎvsG�r�'�=N�Q�ʀ��[
ӡ�\W�I��p�-�>s9������IK��y�sW��Ou�^pϊ�� ]&��|^�`���@*)�D��d�7G3���x��満<�^^�yۘ��������}����3�6�����M�`m�[;�A��`��ry�|慥���;K]6�e��4��D�z=�ĉ'	\����Y�g+x�˸"���Oyإ�~�������lﾙ�+=����g�޸{�z���^;��WM�o[�0�i�j{��/_�ղtPE`(P���UW\V�Z��Yc_��:.awr�F�'%��Ո�����j�Le�X���:��&c��=x�B�+�Bff�Bģ��q�f��Q�P#3�۾٧��~cá\�q����C����IG����W@���&yysy-�1��Ԡ�����~�s H��r.X!���lV&��yy�0Q���);�����;����R�/8,��U���5�J�)�������	}���ס*����⣗w���/��d��m�԰��=�v��+)�tp�� ?�M(���T��=ڸ�K����N-�FC��m3��<����"�O�7�z�%�������S�iInw�FWd��7��������?�uzԁ��cR;�#ɪ��R�\w��۫�}Ԟ���c2>}�s�_O���/n����]�#��,-�{.�6Y��%Xu�ႹM�޾Dm�t�ܩ�6V�>ZQ��ʛӵu��۵LAu��*��S�l��8�Kx=��V)�Ց%����Y)�x��Y|D���tݕZ�ܽ6;o<���2�dQa��S���o4���&�KCVb�|4_+��S�����X�sl�nQ�o��G�k!y�#n!;�kl�I2�N��!f�������Nrin��o�+�vVfUTZέOFV�;R�y�ũ�5�N[�9T�n^YWĭ����v�f�1�fQ��3��v�.�΁����iiWO'N�%7D���]l6�^�T��i�Sl]��Y=�]��{l���ފ���:���(يE��a���#*�u*��(K���Ў#���^�@��/)Iy������/�����8o3�C9��\v.'�4k��� 9͠�����V:��m���:��"]\��#���P��k����-�W���c��;�U�m�2,_'�)��W��	ޑ���B3�n��M�r)]}b�;�F��CN�<o����z3B�AzU�xN�Y����;o�Vl[|:��N�u!y�
>v7����Mo��0N�z	�ugV�l2.O&ѹ�IԈo���^*��+���)�x�D�g0m1�s�^t�yI<h�V}�
$��C�i�%-5r�s�1Ӭ��](���68;�>��5�9�ĦW^=���/����s�|��m�-0�K�`J�+�M���mk���t��lwv���uN���c8��'����B���cr�yY��6t��e�k:��= ��1��Gt48;kC���t[n,�Ĭo�M[ǫ:ˏj��h�ڤ+d�hؾ�|���Ӿ��Z �yH�}ض�AA�n�oi�7��M��&6z��sU��v��|!�O��%a��k,�/�ym��7�wC[�fl뮖�]�+��<�����p&����f(m;���÷�=��ˁɛve[
���lQ�[Y�cw�ڊڳ}�Ȯ��sGt�U�����Z������x���Rlˮb,�+o�X��v�z8�&�{�)v�Ṫ��.ZKr���ʳ�Q�#wd�vR]�y�G�%M�s�,����U��h+l]�r�gy*0G�z�%�ѹc��b_x��德7��c��\x�2�Û��}�ݡWWL�e1{N�N��,eu��U٠�s�m\�MM�����>�'.�����/�QJ����G�\�%�ke�R�Z,U�S�m�w�������|c�X�aCd��k����k���t���w8��aƹ��U����C"t�H�A
�Q���nQsr�7.W/���t��o}}q�z�����۷o��1�j/�\�71���]I*���RJ�D�=}x���q�q���z�>�v����ʁ���_������nZ�	P�Q�۷o�v��q�z�����۷o���!$'���T	R�K%��|י�'q��ۙ/~yx[���¸��/��o�o�q�9F��$�+�]I�Z�xג�Nm�9��wv�n��ђ4^7B� ��c&��"��tW�F�%M��9�ݒ�9��J���7<x��݉��fKI��wvh�%U$�D�$5�2y�0�ey»܇o>���e��ͮ����%�Ł�`�y8w&mYFG���]��w}�7�[����o7�mY����9���gs㰦k�[ 1��Z,3�tܒ�z+_���7�0��U,ø�Ucx�E��c$� �)�����q��vbZszNgd�<�[j��h��� %8#M��L���$$��T�]�8+��T���~�!�I��>B'{���±+�qwM��J���VxMys+��h���D�4K�	i���GQ;Z�<M�]���+T{��8u5�������;+8��)��[M"�gX{�T!z���v+�^�����Ɯ�z��(Q���)a��=>_H��Z}/~B�X�P�(��T��0n꣆�a-n����w*���Y#�n�SMB�k�;&��ӕ�k2�-��~>��+/��o��r!�9�פ�;�ǻ�]�T�w#i�&}OA��ƭ�&f]Rұjő�*�m	޼��1�ݰ�'�͙t��3�}��2Әd;ﭝ�w��)�3Gi� �������|�Q�����n��I�Z7�!�(����A9֊��':dU���΢a6�h֮�����{}.N���w1�%vѝ�����Lk�rgo����y���+[F؊�c���=�%���]V������i��������XԊ#^�5w��y����ٳ
k�kbt�o�]��b���̧���\o�	�����m�6�N��7�u��S�v��W6w(L�B�Žw���$�E$�R�5�Kn6v�4Î���-\[yU�V�xtS�lb�+��{�5��
f������A�f<�Lͫ9��&��c�mR�K���n�Y�g������^EN�t#]�Pc���'�<J�=�|;��@�z:%�mO�+��^���Y2���ܟ�D�r!�mya�7GkP`;���/�`�PK*�;�Žm���L�'*�{�ȣ�O"aa7P���BBz�_o!��a��E������SYXJ��f����k���	Q��
��ysc%�� ��j>�z`����urb/+�ɪ�lv��xbd�V*�-�]��M/�7,��3���V�f��뿳g� s��ıkI-V� ��C'��̡�sU%���V����#���M�ͱMolŧy�鼆�p��M=���\͆��=���x������Ryu���^�}�9�\��	���[���r��1w��`���X�&�֘�X4CSM��z���b�wV�m7� �n�j�`�0r|~nu�;�S�ia���
}xkכ�:�q��]
BF���^����wʻ�7� �q.�[���0�@?O���Y���b4���]�=B9D�Y��n�F̒��7���s�wq��a\��YB�DW{�G�9�{|��-���u���/�O�����#0�7 �:]b����ސ,�&{�5�*�Xw�����-�e1���x�����î]� ث�&j�5��z�[��9PI8�wo���f(��_kd��%�5�n`���k���I�3�|�n�/B����v�Ċ=�;��8�F]��幵����9�XT�n���*=��}Fb�t썍5^&=�B;uE*�R��m��1��U4pz�M�|��汝��"6�����ι�����t���ѱ�Q-9�j�}�R8C��sHvk˗�mY[�*U�!����iΡ�!5��Ǉi���>x��/���gi˫�,ը�]��!�67�vSk-*��C(��}�J؂�����2�ضY��Ҵ3�L��w����y�޸�{�R��]�#<���O�C�*����}ն_i%������6%o�܋v{�߹α�b0`ұ��]�g@������dY�̩�\�x�g�3%1R	m��B��h���2�y��14G4�U�2f�2����Բ|��Z��u��=�F��e�xź�,(�E��خ��؄p;3=�W����S��ݴ/H��+��,�t��6�Fu���2%wavC��l��:5L�5��(z���y��Σ��Y�E&Ԫ	-f=]X����(+�E���gB�\؞��`usM�}��2�m��z���ܔ��T��z��w~�V�S�xA.~��1U� Wdny�f�Փ�.����x�ܸ�S\��o�s H���}toG5]�x>�ug��_j(�챮��ߗu���ܒ�>ٖ�{̱�e(l�,�[/Ø��I���,��*�'C�����Bm���u�N\A4ޟ��L���oE�W�̮{{��8�����U�k���t��{˫wT���C_�)��uN�x�g�3�U������h��:�ep/D���i#�~����R���X��T<3�G�H3���Q�%j�(g.��w���j�Mp���N즥��U:#�pFDq�Q�6�Q�`�Uܻ����\��6gxWp�{��2�SP�`q�iȎ�t�Y�UD߸��䗺vʛG2�J�;.�Mֶw��?�9	-�����7}RøϠ�O�OI��fmA�Y-�����p��$�|�|+�k/ƌymn�׾`4t4�h`���w�tM����`����(�����$��O�Q�Blz�yt4\��&籁�B�qN'�&U���+3Мw��8�����U�p�K�4,�
�	�X�g�*�P�.�����H]̰HuO봒�,�O�>�B�}ggw}��G����"�?H`��~���j��F�k�I��F0��+d:�C�as�����Jlw�n�lOa�#Hw@{�T!�0&^���G;2�L���T�&�*�,���x��ī2� �o����G���	Ki��G/�ڼ�,WOK��|�`�����k(at��)B�GFKW��Vd��b�|wI��#���q�Z5w�Vqmj�C���`��g>��q�v)�s#Af�����ޘ���+T��p_x�24�k�칧[ޛ��}�)�u4l��5y��QK4mW�x�Ύ1�#������B�pW�n�m)sn�uO��z��3��y�ImT�{}7�=����c��ܣ������7D�)��vl��榛R������MD��:qG%�[Џ���H�\�9���Y�>�`��]<;�	�Թ����	�)(�ݓ�g��Xc=8�n��ɭX �Y3Ug5mVG��>'M�P�q�:9^��>���*��:��1�ǳ�Y��uxh�x7,��9Z]�1�Ru���a�fH�"����
Y�!��BlW]�צ��x���7��ݘWƂ�{�c��0iaڣ!���=���g\�.�)fw�p��r�	\k��T���������%��qv�/z��l���/3]t�쑯>��%IGj<d	�n<��r����xF�mZ�R��r�)vH�N�l��[�I�*�՗ն)|��
˦q��G{{S��5h)�& ��(�5�H��1;�mY;���as�{C���_�+ZV^��7J׌4EwWm��9�fY�x�,wQx�;��������]�t>�R}]i�)S�q�9�Wq-�*�\x���Q8%��`W��Y>�dV��.ft���N��6fKW!��2�o�7
��h3�z�$ �A���z�^�u�g�~�Ԅ�X%�o�f�nei�2Ԋ.�׺�m�F��
P���Mʱی��\V,ڛ�Тt�n�)t�T��E�Uҝ�s9,��b<�8j�N7q��M�G\���r��ᨀ��xL�N/������MѲ��
�m��y�����<�Ȼ�q��\:��ƺF�Q�fVU�����ۢ5�q�6�>lP�r#�p�jњ�_F;)WwH���㙑9�U�V�3	u����gÝT�y{��0��<�Q�����(�vv��5�(����r���w����꣮��y�B1;��0%{OW�!ݰZ#�7�ӣ{*ʷ���t� �,�(�[Ĭ�3��u��F!��ui'l��i�\�d���G8��b�M�ٍ#F��zI�Bf2���wfw���L�#�m����\��s���� i��#ޕ��Tj`�fݺX]c2C)�0�G�x�.4������e�#�����q[�&�%�PއU�HSw����y�يsY
I<�`e�SJz���-l��hQ�W)���[��9
lGtB.��X���퍢����$(㾣�n)���5U\>��(�W7�~
Ҙ�OѶ64��5۪�U{�!>���ǎ<�xg���@r��Dm�)����jD�e���ӻuX�v,��{�����C+�h�48Ý���G�@��ڮ���G �L*c�\�';�s-�V�2@�o{��Ǧ``-����9]�9=���0�ϛ�픥��r��k.K<ۂe�s�:�oLಇ��;c��Q��ʷ�ֳ��{�/8L��+UҤgݺ�\�{0����Ww��u�{ ����/@!Ou/	��U�P�/)T��zC��C�炖p/Y�A Zf�;�@�P��E��Ub��dS��u�.��X֘p��_I�;3n��d�������|�R�CL��=�4]Լڙ�Ӆ8&���V�T6�1X% ���aE���ɸ:��� �yd�cT{;�lz����y�ݝr��ڣ.����X��\�L��}JT_y�W�����˨�Ә��M���_���<Ϟ
��(�Ǻ�M�}
��z�ٗ�ӛ%�oو�w���*�[�b^�4�8,��X�z(���}��n�⢎3n��.Gl'�Թrr�<�]#rߤ�G�/d{�������F�b��k��Af��fA�7.�c'�Ζ��[>j��l�܎+�r6V>0�͋i����qۏ:t*'ܞtZx�;��<ci!���]�\��L@���q<8��0)w���:r�Rv���2��MA����kv�N����e�C�f���i�D.�
|K�bx󒞻�e��s��[7#�T�U�-��xf�x�`�g�s���u�.���Â=��ǽPg�{�N���
K�g�Q[;`��0r)�!F��x���.n{P}�8 �9���)�槼�:q,T@��>?|#���|7�p豦J�V�<�=Ƀm-���2P�	51�5{��}��r��h�=򂒭�Y��PDd���E��S�AT���l�����s<�-�W	&���ަ��v�y���K��Mze[��:�sV�Q��X�Wֶ�o7���Td�J-&����{*�N'9* �R
c�Yz�j�.�7���vU��1�N�+>���!�o�*ϸލ����R9(�
M�1��)���i��B�A5D0w��!��������H�`W�T�}v�^k�/��p-�^�<��c�<z
�?��ח�4�O�}6����Ws��x�%��D�d���j��<y*�O�8�o�ޱ������&.Su�W{Ÿ���z����^�|���%O��ji�*�������z06euM݈ ���������x�����vfl�[�d��仺�p2�}��!Dkx8�A�:'o�]*-��`����[Q�&�鱊y+au{���K�&��]\�WN���U�`e�������Я�E%����D4��������:��;hEHِ�EH���vLolم5˽�L��K�u�S٩K�y�1d�1K����eպ��E��ՌǷ�P�n\���n�}�+^��-�|�Ꮝ�&�N�_U��v+�9s���fTW�ך�͆�1Y��2wT��
�%��3���]�!E�ǻ�T�3qe�zb��_�sy�_K��4!�/z�P��u������יl�X���E�3��w�'wn�0nu��o7al�c�ꠅ�eiɫ]�-էK��2�R�s�HgP�|͆��([�Ū���hN48S�-,�u���wCkQɯ'�Sq��jĩ1��U`��l�ɵ7��/^�;���tit��j��hm�%_;w�J�P�<����j�+Lv�NPR�u��6l�R���뱊��zyC9����ܴ`W�ctP�b�&+��C���겊�*׍��1�uV�r�2ސ����ة�\��?.�.�^<��>��2/��`'����m&�y]������fsXgoj�åڊ����\�ޑ��5��/��报E��x�짹�9ݡ��u��P��Æ��Γ��_\*��u�y:��n;����opev1��a6��˧
T�M���rn�t����v_1�N�s�{�fF�b����ڏ?X�A�7��Z������y5Z��'|�������Y;Մ��G}kP*՛��0�.���gT���h9Wm�:�a�.f�������M��j�NkK6$���V�ʜ�V�c;�%l�ap����5��l��ƺK�E7D{���6*��"��$��$�>tk��#��!%���8!��E,�ű>F85էܺ^��C�p����.�2���V��$����o)��9�zv�X4�1�>��BX,w�QM��N����낶����6�N�=%<F�;�#�9����@kYw�\��,�7�w��ہ"�4����gv�,Y�=*��>�0 ��:�t\��\np��E��ܣo8�#v������{*��
㛸:�nSN��f
�Q��B�r�n����s"*��]R§�Ccw6˗�Ɖۦۥ+�ɧ�4C�@�0Z|s�_;��u�^-����o��}4KJ��Fx�=.�-��7����r��O�:��	]�.�N!e̻�;5�թ�̼�a�<�D�$Fv-��&%δ��yr��W\�P�Y��L��e�.��1WI���/q����%��v��Ǉ�6�u��.��Ԇ�ʖ�]$�k#C6������,�1̼��������[�e����R������x�rK��^V%��;��5 !���&�׍U�V�Zi7�u�\��W#k�.�R�c����k=}+zHF��� ��.]ݶ�3�ĵu�*Tf�W��V��V��|��=�8;���Q��㪶]D ���?:� 	��2�9Ϯ����6�ޗ>܊��˂�{���;��������ׯ�8��^�~���nݾ��������zt��(���FI	UT�	'���U�v����8�8��ׯ��nݾ���F#r>���DNuT�.)rHHz������8�8��ׯ��nݾ��$7
$$�$'�&�4������1��;˜���y܈C�B��\���\^��蓥�\7x��S�IzV�x���J`̌;�"�Q\��]s���ǳ�Lb��j(�6f�M��������@2�yvI���HX��n��뫅뫉�@�u�x��z]����v�9�S�9RD! ܻ�P�|I�H�!�����[���l \@��'$��	��#�!�D[
fFmC���p `l�����Ă�nϩ������nĎ^�����pp�pl7}�pi���H7�@s_cw����5�!�5 %d�B$"?$
DF E���H.`��Q�#q���0�İ�f2"�""�&�!�q�c��i8�NO�	��Lh6 �S%��3d��P�!J8X�ȏП��%H�����R3fYϼ�<<<<(:t����t�,#����}О��r���� qғ�k���^2E4�7�k<[��)Ɍ���R,t�L��ϬF�f�i�p�UUs����P�����ܦ��'��d�ʇ[9����*����	��p�]y��
��df�gˍ�7�TW���fn��g}(�D��^R��4%�H�`w�͗F;_���>��Ti��<�;؜���(�!�A4u��\C�ϰV��rhJ�mL�Ms����gKn!�֯"]�M�6�̓A�V+''�=����bB0�֨F{;�fQ���ٳ×l�����r(�	i�!�X`��^�s����(�ϊ�z�Q���uW6�k�V�\$r�"�}����h�>�}��,C�Yn�,�J��9n����<b�x����[��+�yw���������Me���X�l^5TwYR*�y��"�ʯF��� �Q�ö�K�&'�L;�b��U6i��7�α����ʹ�Y
���c�� �N;�7(Y��+e��ot��T	X�!�۷�+��Fb8/nkuk ����&�0�g7�]nu��+=�|�f�3�J�̟�1�7�d���OH�޺|x{�5�{+���[�r4�;ޮ���O;fЎ�����ޣPt�!��\�d��~����η�S^�i(���q"X>ķ=$5YR��!�3�mV��+�������
a�1�#�sz4Nv�w+k:����0w<۞�I]������W�a��ƟYϲs&k���21�q�^�c�颫��ݰ/��@;= �X�^�R&K[���ǧ�:(:V+���}ݵ3���5��=�!�������G3��=�,�]3�>���a��|����ף<���0z�]=�`�`��a�J�-�u�j2)��L��Å�}q�Sӱ�h��{�˽4tX��͜0�4�{zdǎ�N�m��7�p�sxЈ�T!y�f�䭇�̜܎3�}���@���re���L�2�e}���ȯV�#�p�I\ӷƑe���ɵÅ�y�Ɏ(���(c�Y.�s����k-��X�ma[úlf����D^�"��*�����+ut�i�,�2�V�p�wL��]Fڻ�<O�zgD���5��	�[�L��k����¼</�n:����/�wwuh��gwv�Ԑ6 ���a.���z��7׵��箯�*��>�>�'���<��#�|�B@)4.��1n�Ѐ�
��̫8����at=���VNxY�@{[�zB�0wc�^!k�Y�H�S8*���oc�>��;�0tC�MЈ����S��8��t>�Qn�_r
�a���76j6ܟ�梟�bg���
�{���m��z��Pw�)j��Ko$�<N��8%���=�Ț��q��kj;5�oIo`K&9e㺗G�PPU3�'���8D�mRt��pi��Ñ����Vz<�&���q�ڗu�z}ܐ�����f�;�҆^�째�wp����TG���[5��9Sڣ�ˇi}+���F�k��j(��u	�	#�� �GO�\����^^�w'�[N�>*�@��R814�-޹}]�۰��'Nq�FI.ڽ�Zz����
׸f���@W��0<سѝ��wAS��s�K��8b���y\t^�w	\g��~9�Ϛ�(����,�=\eH����y����T�R��������a��d0�dy���W�O��U�b�����뇲�q�Y�I��Ǻ+�[��l�
Y�o�ˊ����=<�]����t3�=�56�Y�+Mu�W�ڛ}fX�`��gi�ڧ������y�gr�m,p��(�q�S�㱒N�8���R�Nv��ۉwyR�Ö	d���֨@�M���*@)�O�ppJ�Z�"u����f�XHE��Nz�K�E���R��r��6Fe�{0��CSv3�U��Ͱ�]��̠pTys|��:6}�=�|��^�7��U�W����4�a�� �[�ii���:;I ��_7��<{ay�%b�t��lLB�������f��kdZw:�׺\����R�sY�OC�8��ر��1[�cy�>�W{aO���gOTr���2\��V_��p�;:[!���	��ս�\斫�n
�4M�Ux/EN<�o�fd�ň��{7��<\~w|2��ŵ]�s�J��e���t���xӌ�������7�N��N8�I�������S�=�_�<<||||��/�U+�:I��>��U>��ܞ�ҝ�F:>Җӄ��*L����9$�c���]*_�_��;�R���tn*��k��g�S6��Y�� �\�!N��9�<�����3�;���"v�V��Kfgp}���N�k?3\�vϠ��z%�{�6k��c��8���0�nM��ӛ�	�!���p�GeF�͚��⒫۩������� Q��ӕ��vf$3�g&�y*;�ܔ���yI[m�<e�ly�h�UN�t<�a���N�\g�;��\�|+�<��d+�!Q_s
����S���m�7���}���yT�R"lb5�{��zLEg�/��畟�t�2T
��<�+���ֆ�� ��=�٭}d�;^HƲ��͉��ɫ��9��N��@�x݄>�~�#�.s��2n��9n�3'���Z�_����T"�讐h3�v�@C<L�8�w�5��>#��l/�Kc���L&�6`曳����[�q�sݕ Ͳ�ɖ�^@�n>�u\�qt��wT��ի��svtvc[α�����M��Ѝ �F�i`���Tۑ�}�ASWv�v��ڿ��q9���N|���̬��2�ζ�mtE~���xlB,�j
��n���	S�O���<��0�!�{�F�UCvʪ���X�p���H�]>J����*�Hا20	g�c�Z�}ַv�٘MtB$�f^h�j:6��{�V��)_+��i�m�t����r�K���4̀��w�ש�ug�2dvb���:�����X�����KL8��6+���AU�Р����#�vtU��hY�H�\���:6r˧�Lj�(&gc�w[����$'��~�� R˚֎�����Y{c��t:�WWR���ߍ��ꀮ�����r^`��f���V�9����w�Uw&E&�R��_�C���2��ql��Nvi�0�����AyHǉF��⦊�=m� _k_����&��3c�i^K�ão`F��Y��lA����꡹�Wt���}�NWs�cm�Yi>�j��A�����X��%{�����5%\{��r1�u��WKi��*�C��o�D�.zG���dD�~ #�(,ޞ����u�b��3�]B�����"��Υ�	��,ٺL�oOV�Ǎ����n&gp�\���lc��=�su_n�|<�7_A���hߌy�śȧ|��YcMP��5۪'�zg2���]�)M|Ƀg5����r����_�Vl�fwJ�U�6��#T�l\ٝr�v'��jM��ܡd�z�w*�
t��!�}�m̇'�ǖ���F��iSz-UY̗�ӴV��@�{g��2��X�_���P��|p{�;�!���ɓ��{����x��˰fR��@�%1ԅ��Ez��l3u�~z��f3xBT?b�?y��e�������#Ql����x�pv��U�������}B�y�����ݤ�qb��֍`�!Ou!�D.G'v*�Mb��t� 0n�9�,�h�;����ˮ{Ӂr��Kʥ�wb4r��@�x�Gz:�f֬mF���fy?������=|��2���V�d�έ^�� �%H�R�)=T�H3OM�uQohS�2�3��ݧ�#`Z�k�NW[�ӥ���hR���VғnԡU1�*��:%&�"���t4L�1'����u�,���7o���o�.�T�����E�}�:Y��ГF��o$�e=��¦֝���}���T<(}9?����V	7����|�t�*��w-�Neu;�=tL�M%Oeq�7�s�R�C&�����F������%!��ٛ�h�>Ω/Rs�R��O=ù����?`��ܮ�]�b�ͽ�}�z��5��eQ���[�K۳�`��[��dG(o�ks�W�i�m�Yp���|��#ro	���}��(6��_{MC�:#�ջ����0�%cYF��ijK���Au�@vR�l8?�s�5��j��;�V�6J,����=Թf��U!����kdр6<�4��||�f�"0N	W͋��0U��wNd�$[j���'u)���n��P��fŏ;f��|	`@�k��mP�zi��ޫ9*�*AW�.�;�~""7Z�f13���s �fP�XCr<���X2�f�������]	�"�m�vk�[�������ǟ����߸Z&1J��MlA��Ӥ���k6�)�sޥ�	�A9<��y;W��ف�����Н����c�Z��G{�)]���+ŤS��9�-nZ�]W�x��=���ޯ0��y��l��jS�T<]=�s�w65U�UU]���h�g,�I���'K�c�,tIh}�nC �x[y=w\MI��؍���%�]��+i���L�����n��^_g�� �C�<���]�P��������V��R
kOU��*�o|�3mNLz�k�@�Lʋ��e��ҜW��Ȼ�>��5����jS�y�w�K�e��J��x׸���ERs(h[�a�����u��c��W����9�I�`��N4eUv�f�3MB_%�:EN����؞;���p`�S��m�8�99ZN�=�yW�-����7V(�:���͗��٦]э�S�&��qfw9'���1��è��M��p#�#��~�ҡjn�z��g�"(�c�܎�Yԑ �"�(�u�g�M��������DK�nol)��΋�vz�ܪ��,�[����m�jYG.q%EHc^�ӭ:G�N�P���a�q�X�k���s���|��{:c@��n�Y�R)��ϲ������K�w��p���,�8�V�Ni�B�]����*o%3V�=W�	��h�*��(�y˙��V����1��3�|�z�>����L�@��I��i�rU=*"�L^�}�u[q����>�`��遜f\QT�r��L{OvΜm�N�%�O��n��gЙ��>ڑR���5ج�u�c5d��E�rl���>��7���r`��k��<�fd�D����_vm��4<��n���Z
�'�q��|�^h��Y7���8;�
1�����3���w��ie�g+ך�޶��a<��^/q*��9��j�b1�8�Rxv������J5�j�~1�jV���d!�;�{�kH��v'���rRe �wAЌǞ=C�(-���im[��:�#ä
� �+mƶ�u�YV���Gq�ˉ}�Ԋ�5 J=�uv�i�:�f�4�E=vcN��F��r5����s�o�[@S�uS��� ��K�[?>�g]�r�������
����0�f�Q���laʱbQ�L���5Ϻ����]aZ.���n��\��0��1i�b͜��p��W�^-�n�n��X�[:�a���/����kۄ���dֱMIwq�H��N��被n�fɕ�U�[[��.l�|탒��kuVSlC�V�����na��v֜ʣ�&��9����g�|f)��칖<˯��:��"'fgvX�?�S%�zP����.��bպ�sx�D�}{Ɋ1�n��7��ڰt֮&�6	��H�ʓ<��s�̮�MN+��Ȫ�2>ܹ�u:ՃNYlAnBmܡܫ��/���9���Ei�t�&�*�ބP�M[ aR�Ws��}�l�K���ȭ�J���q��|c����P�f��b�u�΃̲���K��M��Ƃ`��gX�h�*mJ���:��{���$T��`���}o�,���J���V��/P�Jz2�:
�a�/�N�A���3�f���C�J�le-fy �o6��(��U��X1]q;�;��1d���ʷM���7&�I�-֮#DS�Um�ӧ0���6
���6][|Ȯ�a(^��\��k��d��7�'&>��P�[����I
�(�Y�j�Ӯb����=�!�M$�AI�D��d��!7XÞ�	�p\����tԨ]x�����u?X0� H�[�H}� �b��iSK��?I��7�g�b�(k�����:��&i��(1K�t���W�$�u�ox�۸�VF�����y���G��5����-��|�3��ΐ`��(Ty����{����,�s�>��� "^>K4���L�XY.�(ޜfYQd�O�[.S9h��#'ol��E�w���>|R�}�v���Ï01ʓ���Ǫ�%���
y��,�U�}Tiq�GǑ�&Q�2����
d�;�a�*4�T�#|�\㳓�W�{��]Zt�sZL=��h8�Iul;]����uu���v�+��.�:J���TB�f�딊Ȟ,Ym�7Ų1��m�ԑEf�b�6�;s����{��^a	A
��	X��[�/�s#�v!���2;ھ�1{�V#:<�a�����|C�	�l�xnc��Ί�.�s�_W��J����9_Q�{-�^Kqhg��X3rV�P�;�I���U�dmήg9:���ܹՍн7��ZǍrWS,�#C喱V��[&���K����ӵGA�۴��8#�F�����|�zU�n�Aۍ�t�Ŗ����}�.��6b�9�I+&ڵ8����DT�̎�s���_V?$�w�]��I�;��q������=d]痀�* H<aH��sN��o<�4.�J�*Tc$#UD�|z����׮8�=z�����ݻv��P�*I1ˡc�r���;�9t����&+��ל��~�{�{��8��qǯ^�}}c�nݾ�]q��dd��WwLe(w#(���FByۯ��������͎8�8��ׯ��v�۷�O$B�v�t`Ċl�h�"�	��wA!)�q


]�bB��s�%%�\��%��t�M���ܐĖ1�La˦4��K	~[��!"����ˀ'��~j�� HI��.�"1)��Y)�y��f�]�F���dz�э�:�do���8��DG9��,QI"��v�W�-�9���,��@J��gQR�#nP|�iS���=��M��?'%}���£<�U���<��8_�����kh�K%5:�{�7�!L�Sr��6��25��0Uy.����0n��"S�
ۻ7�;�Xk�����9�K�AolzE�_��\Sr��*|�����"n�m����.-h���%f{���p�eSۖJ�*���l_h�vzjݍ	�r蹪�g�)����(oH��\�3�7�꣜bE+�߻������;?n�F6�*&�S��<]�bm�͆a���ΘS��5D�3����ʃN�������d%]5Y��3�d�x/\Gd��#��9�{9�W7���X@��?v�<MPS�{n��Vb��|��,s����*�>�X�Ț�v�K�{,���=E2�	Z�!���XZ�ϝphs�l᝟�<j��w"tk���ȗ[�섁k͂@7O�r�/3E�|�{���
�ec�.فhx�#OJ�3_v��J={������ʱm6�K؅A���&iHL�;��/F_'{O��м�6��Td��c�ji4J�����Ƈ8��]X�V�ejL!S!���3j�۾Q���.7شrؤrVl�j9��ѽ��k��յ��}nz��o7���:6�hJU�ק�!��Rj�O5T�ih5�
7��ٖ��e��w2�բ*�d�u>Y�a=a�>{�U��Wu�C zoF�Z��D��w[/2��Ntj��T�֔n�V&�SC�r���i����P;6���M���Ѵ�@vuu��=�U�5o
�p����R����YGn�u�u�(�y���˗U�e�M7��==nV8���rl�x��Wq�i;�'��v.3�ܐ�8��u�RՕ���W1�5�MX�#8t�{!z7C�1�ށD�����Yt[F�fMZ�e�Hc��+W/yZ�SH�?_�瑒ÚR�*��6`��q��Uw����.���>�:Y�-m�.���w]�N���LDf�}XqUiG����3��c<����B�����6���FO�:ԑ�eu;�V��v�v�T[�ՔsZ�D��G�H�qݪ�-��m���<�2
����|H��	^�{�B��\P~�u���"&���] }�i}\m�a�Oc�q;\����wW�6���ӜJ'��EqcJ�a���������[C�/���#���j_�0�w���u;q����E�! ��_�c{}@�Ɨ%J��+�S���=-BΦ���7���	��U5���G��������v,S��T)5�5!�&נ�E2���;�
�|�L�m�����ki7Y4�$mM(Bn@������J �U�E�[��0���'i;N�D�l�NA�p��x�I�`�ח3e�x/
�@{�N��"��Mj#�R;o/<m�(m�����#�xoj�^_H1O l5��Z����x�x%_s~���wBf���)t�R����L`l�����g_y�j�o��mL4m
��Z�U��H���"�{�_w��%mϯ}�¨T�C��b�J�0#������ɠ+��t����K��ƹY0����8�wf��Lf���w���Js�'��v�U�dM��۠�j]�+U�m���ʋ��&J��,Mj���}�Zơ�*��
��n�e̾ �%ҋbj�;�zx�I�ng�\����x�WM�2hRKӁ;��p���ϩ]��DK�g-Z�"�ڍK�s�\^NI�C���y��of�@��,����N�U����~�o8OL����X�ᓽMGfn�m�td��*Q�\����vI�,���p���=sZ2"]u�ݫ��γ�s7���B�|���i�޿Ws�;��!�n��eˤO�����2�[$�^w�}��PI�)ryKu_(n�¼O;uW��9�LL��`�sc�����F��z{}[4j�'����zHS*�2�����ڢ��/R�ȤWg�p�4�p��\�X�dk�f�S�U��L���S�`^�����׼*�VT�#5�#��~�>x�������U��$��W�Y{E'�E������h�N�~�gd�ut]Uo�E�߻eg�Y_H����)
bVK`��q����p�E���y0��̣�E�%cu��4��?��w{drCQ��#rn
�iV���Pi��ي���[�赥c�k�弋�n�j��%*�{Sn^ 񣶀��xP���m��3Yu��+�:��b��~y1���@�󗪔�lKF�_��I�A���I�ϘrM[ݘs��������7���ʪ�����S�����	��}(�2<�Ks��e��2a
@�@r��;!�f����/�^�����L�o����@z��>�7���t�i������^B2�֓}^')�����:�
`:1��~�����1Jy'lv�7�k�˺�����z0�>*�=V�8s몘�����B�}��>��r}z� �z:&���j@�v�wH]�M�cn��g����	�-1wsU�)��vwE��`M�M�ݎ�z�C�-�ٟ5��V�)���6̒�L�O2;b����q��=EO��}��Q����@�1c��iZ�������gH# Gl
1�}6�bE�U�6��)l�~ȭ��<�D<������v<vq�׻���bLW�{hlQ�]c���U@�ڪ�c��h���_�L��
�<e�z����q�Ft���h�
:���V^��0�sý���S��P7=��h^��͜��M����:b�h/�jW'.���{��b-�`Lz���"v5�:��uޔ4p�]���Ӎv��E$�5[�[�@�n�T6���3�z0P����� �a�>��Nӥmz��~1='um$M(Ԙma ��0>o!�ﱲL;��*&�g)`���ffO}۠�ʢ��h���Le�sB�ޭ�������y���H=�n�mz;���N򓰧Kj�RN��uݗa�"���t�-La�P��|ΓD��`�q�M0��|+_^5�ƍw۫�u6"�O��ۏ�اS��GDp� d_*h����u���ڞT�O�pg�KF�U�+�H�yH�=���,�G�tϞ��.���pq]o|rs��w%8�/�V�֐d�J�ۊ�u��p����Z�ձzE�8�X��:n�5�HjU)��}����S�����g�?�-v�&V�#���&8�WA������w:�Ǻ��kp�7�{�f<�S_��*���ޱ���z=[�+��n�Q�o%�q��4��f��nQ}�vM�أ���<��"��t3����K�,�I>�R�<���n��Ewe���oK�!��/��뭺�5�:��ݣ�ڄS�\�\����c���i}�܆��/k�@�2b��"�V����~��>> ��ت�2��|�rZ�߷&���T������b\ݡ�UC7%T��ʜ�"@�-�5K�<=p.�\
9tQ;�w�|�;� W�ūyQ�;rl�<V��ɐ����(�pb�߫as[��D��e�k0��9qƶ<{��Gt�и�g��=π���a�A���mҚ��{2u�{1�x�@�z��ϔWv��^ǌ���p��mfd��71O/���eڒ6�t�v��v{�Ͱw�hM?��C�`�6�;�G\5�^O^�oG<���fHpz�WY�v����ej�N�$�͵0TU4����N��)��}��2�i��m8�t)���5B˻n��Y�\�h���ҳ���1���ɟ�X��6.튨��q��8u#M�(�3e�]�|�=]��{{i$�D���Y�o�<8\�~���i�W6�zηn"0�k=ä
Z���Ќ��:��ԃ��4���g7 �p!�X��ʚ�ӱXU��u{g҇��L�P�_,G0H�X�p|��r�MuaMO�r9�HM��}׳1��RS���4�o��M�z2�X/F����&,�N�c���ھ�\¶+�^��%_���� ��|��O)Re`�D�@C�Oz�guV�	ԐG}ua�f+��;���-�!���/a(�i���[��y�
����ܮ����A	��/K�"�M���yx�Y��e
��4��4+�"����:�,c�N�uܴ-��2�:��6m:t��__&gg��>�cL���,���*c��O8���0S��j��;�'�h*R+��7&i�F���>���}�v[��6�9ý�c5g-],-���i�]Lg�wnω̋v	�������ƣ���f�L,U���,n�%@�b�t�o_q�����3�ڱB{�xɥ�4ޱ�r���7'���� �1>���%���w;:-34.�؁��S=����-�~�@~K�`Ԉ����U����ТJ����ZB��P���G'z��r�`���p�#H����7KTnVB���s�hEV��횼�\�7SL��8f̺�(p�4j�	�&h;�h���D/���,3�o��;9�|%;�m�����"Uˬ������"�H\Lؒ�z;�Iu%w{�~<�ӽw����u\t��ތٳ�QP�'s�yJvq[�onܤ�=5��kx?�����{��r�H=C�gs�	p���[4P}�,���X u��`7�M�?������M�����	1{FA����L`�<����<ʜ��8�Ѐ*l[��J%��c�!ހpWN߭��4��v�f�V͖O2^��'/�;�^h�[
�/�����Y�Pɢ6'{m�iӌ��B�pD8�g}���z��܎���r����Wj��)�*�-d�Ma�nޡOqg6�R2�c����L�R���M�V6�q�a<�$�x�0Z��#I���EDϡh�QB%����C��^]꼒��m'ѽXJ��2r�u[�X��?=U�ǽ�Z�Of2���1���8R�l]����wsU�fl0l��=���5�{��-�Sy\�RW����+lȲ���>Z��d��HKz|���'9F�����a�m��d��qZF���5"�Ww/&Uܶ;:������n�OQV����9�&��M�yW��J�V-�w6Z�f�تV��s�s\�bcҴy�%�=�j�̓���U��������������2(��G�á�m�g�\�O��yd�QǓ�7�9R�8`@�S5�N��5�Gv�6z�x:���c��3�7:d�l]*�Bv���i��l#��,X�'������P�<��j�>O�Av`׵��.럴��q]9w�s[��M��	$)n�!W@
�a���� w�oK��k�5����Μ���5��V��J�Mړ��-�7��D�v�����IA]f=�B帮w�uȔco�im�Q������a{�����U8�G�M���u�ct�u�`�P3[�<��Z�w>+���p,{�w	 ҃���P~��s�>�iC�[}���9�T2&��3�Oh!�Z=��#g�Q��d�V��B&���w����d��V.)J���<ԩ��	�O튪��}������G� k�Q��o���T�t+�Ȩ��n;9Z�����Ub"�,f��ɕjjmSU��ͭ�,��R�R�fY�MM�L��[Km�1��5+ic*�Զ�Sm�%�i��UMJ��ֳSmKj�M�1e����ŕ�ŕi��Գ2�55i�Z���ԫMM�jV���5*�k-SS�k�*�Rښ��ԫMM�56����R�6��5-��V��i�mMJ��զ��55��V�Y�MJ�Զ��ZjV���55i�V�����M�զ�ښ�i��MJ�ԫMMjjkSSV����͵55i��MM�5-��V����mMMZjV��U���5-SSZ����kMJ�ԵMMjjm9��)�B!b�AB4�MKTԫMMZjk^`4��00Q��B�5WZ�j�jkj��V�Z��RԫU-KZ�jZ�H� A��E(B+U-MZ�jmj��������Z��RԵ���ր��B�@ �Q ���Rԭ���֪Z�کj[UKR��Z�Z��HP(��B(�AT�6�R��j��Z�h� B" A vZ��-�jU���KRږ��55��V���ԫ]շ[SSZ���ԫK�K���Zjki�f�50%ݨ�	�$�* �*�%����ic6���!J�"E�@jU�L�em,ek,e�1�ճ2���m��������w��A$ 0ED@�O��W����<��>�j?��?��������������a��ؕO�����۟��?p( ���~a�����Q}H��*�w��>���O��	�a�J�
 *�g�G��^�k�y���~���D�����Q'�sB�*�"� E(�55���5��5R�-5�VͪVҵ4�Sm��5DB*0P��D"�B�RY�Ml�K5�m���jU5�֦�U��Z�mKM�-�)kR[V���j���PA$T � խ�Z�Zf�i�jKj+i��*�[R�iMjT��5��զʴ�jeZl�MMjj��ʴ��AHE`��$H�D�EX"n��J����֟�*��(����)  $���@���߯�~��>~_�4�?wШ �A��?�ٯ�>ߙ�]�m!����a����?K� *�~�?j~t��N�W�( ��!��8~a��-E��?� �*�
~������A�((?�+�������E g����}�����E ~�����<�?�3�}���y�=C��?���B��?��W�E @�h�|Ca"~�����Pu?�A����^����;Љ���( ������J@��@~� X����3��"���t���w�j�-����.}m����ޟ�1AY&SY<��H^Y�pP��3'� bD>|���)""�h���	"$�![E	JUUQUEETEQ(T!@�����D��@"�*$U��DU	eY>�]��Ze
-D,���Vٵ�[f�[Y�m�4�ګj��Qf�*$(a�UP�kt��B��ki	�l�(TڍVƓK}u�m�mfCI��f*�RJ͈��
�63M����+,���0�m�lҪ�M��6fZ�$�d5�6�խ�5@F�i�Mm+ŭe��i���Uf��+�   ��ۦ�S����@i��][p;iH�6��UV� m(w�]{��� �G[�UJ�T���V����1�j�j�w\�;�d�+6��i�m�[����j���  np�(P��J��Һho�O�>��Ht4�SF��S�<����ض(kt�>r6
�ۣc��mZM�9���ʣY�k�������tn�v�4�\����MP�N�7,n�һ�jd�MmR�E��k)Ymx   ��=R�7n�Wwv�h�*�wR�쁶��N��n�Gk�iT)�EVi�ٓ�V��TҖ��9T�Ԑ�-�i�� ]���:���6����U4Ve�wm�XP���  �ZF���6�3�r��]��X��`Q�Zf���c��FU]��F���]ͱ�:)�꺺�m�u��k����r�m$[��V�B53&|  u��J�ۇ]*�wt�
4����=�Nⳮ��պ[�:Ѣ��N��+7p��N���GZ�vv�k���G6�3Z��U�-�,+[d��  M��րs��t־���ƨt��:����Q�Uwv:���n:��{hz.n��wwkv�`Pk������/=���2�;5.�JiP7�  ]�K�.�H(P����ʢ*R��y�ʕE���U�J�U�K۞�IP�..�챮w�y�AB#8���R�]絷����Sl���SVd[k2V��|  o|��C���B(=�s���!�z��UR/oyM�*���HDS˺R��w�=�P�3����JEQ��s�)Ii�z����,ͅ��e����1_   ϟ)RUH���x�	^�=��wJ٪A/x���R��{oyOCE"�z��T@�����
��	yḤ�=�x^�T���y���5e[6٭���Q�mg�   �w�^ڤAOq\��W�yǔ!���nT���� Q-��y�T	Eg���)*
;�� $�.�7J�҆�=�s��"J|���R�L@��)�IJR�  S�!)J�  ���*(  Oɤ�U*�� z�"&ʪ@F����?�������	�����SUj�L�_&�`���^z~�����1?�菾����﮶�w��ֵ����Um���mk[o��mk[o���ֶ�Z��������K��{���?Ȱ�c���}t�rT�؅�KpQ�r��:~1��ajp�7k/!ʱ[lZ�y�Tu���N�����Xra;B��B�2��;3S:�c����Țؕ]��j j�S�4�cr�e*���OK�E����&�Ӧ�4~��+lBlҬ����E�������y+��{�֏ٯ(@)�Y�%<�gk�1�Y^�
ɷ�kU�v�5�)`�9���qcX"U�����O�P���Z�Q���ѐ5hԃ��{��f ��@ɪ䠍l�PÑB��f)���(QxM��ne����1`�RYu���F����ɼ%^�Q���NA�Vh��*X��yW�0��#�&��8�[�2e7� ݳ�� n��yN`��J1x¡ywnM������EP�me&#J&^�m(�m[.���u�i`����Ũ:V��&V�o�B���0n$u�D�-�Ebߎ�m©n[�$��X*�lkM(7+o�X�2�}�9	��0�rz:�[�e�-
ɺ�Hr�T�nΧ�����Yl�j��b�����{6�--�6���V��7��˷q��5�+����)�r-2£%Σ�+Q��'kp|�tsi��A�J�꧰��V�6�ZYBK��AJ��V�#Ҩ\��ݩ�뚷��ݒ�j��@a���3%���&�p��7v��YN����t�j�a1n��s`5(B�#��eԠoj[L�����H�i|���"��lܖ�����MB&��Jn�$�&f%��N0���݌��4�A�j���"�5,wx�S7Y��$Tg5�٘\��kq�W�L$�X&��]]��9�������Ib���UXt������Kn�7��)�Y�X2n+7Spn}����I�g�x��T�zTB�+��.nEi�[x��vE���P3fn�o`��HQ:�	XM�rS��3[��*]��F�!�*�4`��ۍ����6�3�	`AM�36�W���ř�L�Yy�J@�`Ճ,8~�-�^�[�,�.��ʹx�L�Ԇ�$�Jԫ���S
n̻
�i�V5�Эs 1���j�3 8)Jt�-���܃V*����E�v�-Ee&�!�+j�*=���ZH��B���N͂��f�hZ�r` UY�,��f�Xӊ0���R��&���2�^-OoT��W�s� �6����f6f��t��"�ĵ���h3{lE5�
iQ&�]iLGa:y*�h�Z�{���'� .���*5&-���/5E�hm�7ejr�$77��lݒ��e�U���w�6�kt���r�ؽ�J"B;�)rIH�XiӼ�t�c�y�k]cd6�L�>Mku���Z-gl���.�%�h��d�nP�M9���Z-�����e�����zc)˫��3�{N���ܤF���Jʕc@R���U����r�(�j�X�c*���� ��MXͰh�R���׎�֩� J8-�)�b4R��*aa�B;da���E���Xx��*���D�q^�k�G�h5��Z�_dƨɕ��M� ìDs�I��)���vHݼͣ��ʽp����j,���k%��QC���8M
�Or�	�����]�(��ܫE��*論��4�#J�N����f��SH��<��T�D��k{E�@ńG��+�*?�e*B���)�,УF����Q�Y��9�+eK����d�����#u�:�*ƭ�\�ە��+q�Q�x�F�٬2\��F@ں��Zon�VՠY��x��\�
ە���Ή�W��*yPޙ.}�; �Ux�hR��R��u6*w��sF2�0*0��C,�Ӭ
y�j���V�ה	Z�o���>=�"w+��crU�',�2���H%6P� w����Ul�R���V�$���آe^hQR�W����K�2��F�DȒJR������bқ�
���-[��û�D+�R�M�nf �O`�B܌�I馦�XTH�l�L��Ȑ�fԭ*��
��5����wn�4$kX�� *W��@����Q�&S�0K���n!w6 kf���yr�J��	��F��d*O6��bQrܕ�>�
��{3TݸN�AV��@�4��ab�S���)�h��Z��h�`ܽ�l5A��vj��L�GF��b���G1��^�Ղ��mnc��4�4�_���*���v_X���XVT���!�Z�P�6:u�q�ʻt0
%�j8�&n��$�e�5��-���8i=�۸�.Q�R�l�j�R`f�߶PF�m��*�C�O�!���Yī\f[�mR�洅��e�H�5���Lv�JAY�Rv��̹Dѩ�~�%n�3�I�uɤ�{�!�4�O2�^ۗa.Y����Y�3m�]3pr4��g@� m2��V��[��cU�5!�Q�v��2�j���X��m/�+��IQZ"@h(n�F�b0�*�NP)�����%Z�5�4�R�d-�Y�NX���9�:`ڙ��Ȗ�]h�`�t�DJ@7��d�i��f�F�ė.���oc�����6.�U�r�L��(�`�Ӱ�W��kq��"&[wY-��Q3[T$�{�!	���3���i��(�hۻ̈́lH^|FS��(�*˃J-b�V��2��Q[�.陹!�X qh!"��R{��r�3Si;)%�#Y�����D1��l�jj�Ѓ.Yi�.޹������Ŭ]^���N�!o�G���*���qkڷu�Um�ݷj���b��)�e
	��w�):�� ��@u��k2\����b�5u �p��J�`���g��.�޵��Y�0�4��&�RWfΒ �5��k�t6X¾ƕX��<�K���h�2Qu%XܔNJ��&З+
���!P�[�Y�`ƛ��ۺ ������)�����wkY)Z�)n=�F�d��OX���ջ�F�b���>�͝n��Ʌ6��ݓ6�/G�+c U�ޓ�Q��,]��dR�h�[0E�
��n����Vv�ax���n�S�����wO1� Y��x�v��h��� ":���V�y�.��x2^�qI���
�e�R_�ݏ�,knL5���(���A���1�6�	(���eߜ�/5U���>t�w�Q:>y�ɯ-îKLj9\����Q�V�t(Lh��Ǎ]�6-��������91�{Bk�����
nP2��k(��-�m���hҚ���xr���H=U�];e
6@.(F"�`Q��+0����n�#��XPa�fِ�4˖T�����60zT��9�� �'�1ǌT/w
yF��t�.��[�Xt��b@�D��۱g�,��<XR��B�����7c&Y��/���ЉQ��q+�p�ѯa:6B�4^��O^HEڬZ�k*wIm�y��m�YN���2��c�#d�i���q��g��䧐m�pJj<A,D%6���<�+s4K�H�O4R6��KZ��C��lT�'Q�.ݪK�M,����l��F%�7&�����V��D��^�d'J�ͰJ6N�2��m�dѱr��D�r臮D����!���dA��Xj�:ف�Gx��֑���RE底{(ݚ�5�{�� ����0���t�����V�
��;�@�Zm���iN���*��'E=-R�4���ı�h���f�RL
��5��h�,&��1u��oQ�Z�*�����$O2#+u��5��uu�U��t�,��� �1��1<�7V�e�]�{��X�5T����yl(+��"�+Xr�۰�ҵR��+�{zrFUc�/�IJ��F��dT�a~�~#[K��Z��5�jү��s��D�ZuSwx�j]9��n�4#d��r��2Br����
���5#V #Jr��V��sle� ÷&��36Q����ʒDZ��t�rH��g2ą�rե���]6橥Tu>�B��H��N'c\b��,�X��t��v���b�̍ ��6;[���rGD��dD�P#d�u�9�曒ޗ�J�Ljkͦq�����l�;e7X�n,W���6�[�
2ݹ�9o�/n���Vm�0�KUx�R��a��� ��u�+nƳ�<v�a�${�N�́Z³
n��Q��%���QݡYX&��/\:����m
��f!A�xCD�L���]�d:�/��@�m��5��'�F�5���N�d/H@�z>!�#v	��bY�d�2�y%bl��n�Q�:4�3^1�m���7���(Ѱ�;��]j��)�#��X�Mz���X��r��� �Y��В<�zLݭsEh0<1����͖6c�q�f�\PЬ*�m�&`��`�ݫz�V�Y1����$kC�+%Z:Εb� mɹR�]�!^%�u�%�{B�7�M[�m०���%��N�����7.�`H��T�B�ۤ�J�(KŪ[�/[��VҶ�ժ�#t�Z�Y�起7t-B>�j��f���D�Z� �*�!n�oL�L��nM�U��]n�7-DD��DM;���0<YZ+c��فa�$bę�^G��VȖ��Yjø��4Ef��d���SY��+���b�n�QM�r��������̩�0��b�9���K���b�2�6�e5r���J\
���|�	wh�R6���Å�΢E�C� Ĳ�Cl^:,�lR��p-ߛ�2��&�OkE�+p�N�.n / ���E��Q�'eݱ	w��E^֕�.:ãu�v�0n"�U�7��d��A���(���̎b�	:T�Y��%<��c\#C ��b����9cZD��TU�
�)n���̼(�͖��]`�BZ�v�W��`ʘ�"P���Fٽl:ۛ)�vX�ؘ��}�單�(-{u#�%�Rj�5xv�h�E���Z�ʀ��h��ý�	!��*0:���{h:�c"�Z��P��	X�ĊY���7r�R���5�R��L�����SE+gqL?vW6�=�I�I�&�@�d�b�F���e����fڈ^�ج153*%��3"fӹLb��iIv��M�+�7���v�Ǭ�[F N��u�T7,�8��:�P^n���^%��`��;S�ȷc�7�f��pi��^3���`n�T�
��T͠�T�1��!��$�V������n��"�֦�ފ���Ƴ�Y�ע�R��I�C��;�1S
�4#Mm��\�[�
��D��1�+*�;��^C�ii˳�)�e�C��A��sf�ܭfS���!�Eշ��r�|lM�ۂ^����)�Z�#I�u�$ml��e�s2YJ5���nL�l"�*yTj� �v]���g��'���#�.
�oq!"�q�Z�HL���Rf��[������$f���FCA�����k#��`���au��+n��Ҧ��1�ˠΕ1�y0��]c��C���[p�i�iŮ&,�-��\�������BQ�n����ن�-ӵq1�81짎�� f�&o�*��fit
�7v��=y�Brk�t�+v�������i[�՛ݝ�fVIH����H���*qbYY��Ss�L�f�Ս耪yW�B�`��YZ\h\��5�Eʱ�[�0��d�(j���^�Y�Ɏ��mliU͚V���Wx��(٠�U���y!�FS�B��[6��tc���J5�ar �H۔��J�tT �lՒ��\Z�y�ޓ��f�wNA��R,6Z���#�Kq��[�R��VJ�~X)*ɣ,36O
�.1 �hJk��=���r4L����46�w�&fV� �������>U�j�9���
�U�M����Ņ�wA�X�hE
9������U��tw7G��; dm�����kJ��OV��N][S,ZY��`RS`�'�`����rT���]-�JWL*�	l��C��n�rӫ�eS�IشV�VU�^ Pp��@���,<u!ͱ*����f��C�`gt)BS���餒*o$ԩC��M���T��SmM�C3s�ᘋ��H@�D���V� ��o(����Q崙ѕfL�&i��g�.4��t5@�hےLyl(L��f�[�)�nm�95Qۑ�&��-�sw$�Ӣ�l�h���EGc(h;R�Z��E7~�Q̬0a_)�p��v�;6v������v��S��X���ע�Cp]�2z���pV8����\�L�A�Y���L�[n �����)��mȶ�^8UeC���ݗ��v\.����Q��VL)��/pP����ڕn�:���[/�ҡ3dH�0
����G3u]�0�ƘEn���/v��J��3l��k�J�%3
L��ޗ`icj=��B�Yb�h*e�[e�L�T�Add4m��-�z� ��s���(Y���`�%ЩA��i����Q7�Vn�F���#n:�Xɚ��N�Ŭ�������5n�=08���+)�������eֲM (�©$r�������.Cj�eYC�h�]K�����p�[0�f.�7 2Vb�O	������b03U޹��'�8��N�2��[�R����!n�0�*����P�m���n�ͣOsJ�"�u�=�*�;�AZi;V��4�\ �n���v�2��ϰe�F�i��r�l�� ܴ��6�S�X���Ǯ�u�f���V>�q���ލh�"Q,Ў��t%���G`�b�X��N�����š����b�LnjÌ�}0�2���h�&ا{�6��b��-f8-'��[����+b��/F���+k,�;pM�N$��j��~D�B;���Ȼ�Q���|�i�l��;f�B\�Krv̓�7�A�K�S05u���������
��2�LŽ��Pc�Pљ��L�̹�j}�ԕf'�^j���s�Py\vg\�]���0��G.����ѭ�(S4��W^۳8�����V��-�围��,��YG�8Qq��+5�y9e��K�lI���۬���w�m��t^�ù��w5w@����y뀔X�WS��c���v��w+3��L|�M|��X�b�r�p�₎��r0��6�Y�볔1��\��vZ�ʢg�AB\1�ۻw8���uRnT�:��c=�ɴ9),�\�J2ej�:���X(�;,R��_Fn�HBSh:r���r���IWB[��FaS�*�s���|M��>##;�Zw���5֘�C-ͷ�{2��m掤���M�4��-Ln�Z��_Doq�P�eC�J��3��MN�ml�z�N�S�|5e6�A 7��r��6�9�CL���7��]��AOu�`��n�vKw��ؙ�.��%N�R��k�0��xR�=}g;0��I*晔mI�ơ�7�LOy��t�8��r���F�P�ϩ�.Y�v�$�hN�M�)�Ak6�wp-}���1�����A_hQ"�ȱ]��m�ۻt��s����
�v��H�� �i�t�u�V@Y�r�=���M�N�TL*ıv��'d�Wa'�>�a܇ԁ�մ�%pGcwP�穇�9�zh_gX�x_T�(�Yyұ����z!�Yʃ����ab�$-�\�$����y�ge�u�֍�ռ�/ ��(�oT<[�#)��ʐ��̡��5!����a�+��z5<�>E%:�*2EbF�C]xK�Ks�f��.}��]r�H��?�q��)��}+&�t��S6I�o7�EY5���f��i&Zb;�V�N�Y�]��N�틔"@l7&�۩�ٱ�z*v�F�׈3�ʛ3m ׹΃�䂋�<5��*��IWٳoL<�WYH�3�G��r�ˆ5@�n�r+Tn
�s�PT[�0e��k��W}�$}Iegǀ�Y�څN�ڤ5�{�����7 5�C��Y�l:f����8֋�p�>O�c�����tS�$f�J�R�tv���b�����0�]����¹ڦU\c�qɺ��Ԍ��+�:|n���G��[�U&t�c�#z�m��ԃ��f<�#�iD�H�vI�&��*޼Y�%�k:�oa��wmֹo���W!�;x���.�i�j-�7 �}���:S�AY�
+��s�졝Ss��g@����4Z�]����ҝ��;��x[:b[�̼g�	�;R�m�agƝBR�6jj�I�I͵��SAmf�`Z��M����|��N*��Ll��ᴝFwp]J�w{�ANR0�t�GS+��J��C�^�ݽ�a�K�oj�g+
+	y��&�bn/TdG�g>�������-
�kv�v���f3��g\�p_b�x��	B ��S;����5c�j��4����[6���Ey`�"�GQ��oq��}f�۳mb	X��i�RD���6G�m'`�]��U:�K���xP�s3�d�0�:�]Ah�w;�wc��,�Oz�	`�(f�͊]�$���b��#�:
���! 2�H��L�E��Okn�)���<�A�X�.��-�+H�jqܖ��dvJ�\�sY��(�#v��2��9�'{i��j������rPH1֕�t���t�T�CQਊ|/�U瓗<�N�Ӧ�X�q�yΝe]kCС�z�8�o�nd��E����U@��L��k���� �&^�a�h�b)v��+��5���
�{A��6'	Ε� c!7�]2�3�GjP����fn�j̓����c�7��������e��m��1�a�1���$�7,[������dU���κ�۾;2�v��WyIj���'H�ɀ4Osʑt�h�H�q�6���QGBT��V3s��R[���J�ɗ3�W��o(a� 5��\��4��ƾB�YY���۾h.�`��v��5�+��Q��F�[[���֓�Tn��b,s�\��vFi�����ۏe:����[�L�7�K����870��O�e�&�fV���@����gV�*�,r���n:�}�>��V��E���E��Y�����aur�J��M�(�(��}F�bΜ*N��d���3hɵ��(�c�fa���:����A�0Ѿ۬U�VJT���#��-������+��B�6k��=jZ�b�jF�_,E�2��KG��sd#wR��{��};��S��i-�cnZ'���ytτ�2����wܡATC�S݊[�.nK�w��sPu��ȕ��(��������d��M�ܿV�)W�d����=�Z��&ԙw�����e9D�:�����lu��v[2ò0�p���-b�S�O����ƺ�c<ҿ�#Z�K�
�!J!`^�r���������T��wP/i.�oK�hAû7����u�ښU�S�|@kVoGPf���#F�o1H�:�w����Ѭ��(u�C�]c�����§f�ۦw$�h Q����9����%�:���͌h��� ��F>�޷�xK���$c��m-���Z�6%Q����`1�>�;���-��j��[�ű}�4	5�'U�nu�3�D]���D\Y5"d�9����c����Eק��e`��^�{��t%��S��ж
ݍ�y�U�9s�y�nJ*�3�V=�����{_9��rH&���Y+6�v]lOs`�x=Q�-j�gn2�=ν� �H����	���r�j�"`��BM�%��4����lf�ֶ)W�|!䥾e\�ǻ�N�s�Zڌl��:sR��Y4�֍tur�c�+8_!��t�ۡI����D�d�i���e96���]��*b]�`BH�FK.��t�B(܃�Q
�,�L�V��WT��deK#M8�5��hiάr�{97�oo=W7�̓��h_�{P>!����!H���Lit�a��Y��*���#�6��aķ6��k��m��ѽܩ2�S�\��d�p�gXw8��`oC�
�$Tp*څ�0�dT=]����8u�Ԗ��ҀzMdДi*
U���{]w-�������d�ョK7J� [��7R�A]>}�^�C��y�%�b�s��'{�WD�uk�9Z�4���;ki��)Rn��������#�bo�l�
�� ��ŬG��R�G�J1��Z�K�ٮ�e��}W2�LP
�P8 �0�.���ǅ��X�utl�'y��V�@�WL���eM�Ǐ��6�c���E��x�i�l��s��.�,����B�T���X����o$��+�3��m�9�w���7�YShQ�X
�h��7���5���.e���%At��@&��L���tM�#B���V8�6̼��KMd�Ғn�����_E�o�={i`ڷ��z4gk{��g�y�e���9�>�� 5Ǖӄ�]S���O����u�c�3^���Rq�I�Wm󣱷%�mN�J�/�� �EpnE�ݮ�7{,�5��E����t������*��̮�reehˣǉ�}32�w$�����'υ��)�<�1��Ǧ���Tv��<K�;��0�����=Kf��n��k�sL�F�h.Y�V�@����unR�>u��I�d�֪0��u3�3Olp��Vv��A$����wc�}�뵏4��'�U�y>#0�vJsx3r>;�����)ffJ]ٲ���_aa��:�W.E"���2��Z�y�]��v(ݳ��r57$�W��*'(Q�V��WKD��� �H��r�ښ+7h��6`8��p6 �)��&�Kmo6b��ו��R���n�V⾘�X���؉ĻC�h�W�1�PM�����t�	H��n���Ʃ��Y���A�N�So��q�QU��V.�{9��i#� ��,e�_Z��Dit���ܸv��X,��;���u��o'9W�vaKW���iͮ��^nq��ء�>���b��Ż� ����+{@�5����in������5�\p��Z�b������7��e��ǋ��*�qw6��5G��K�So]��#�m�vFz���Mm�ٝ�["�ޜ�^��N�_�2݌m75���Q�w���O�
1'KXp�j�S:A�N�v��v--�[Nw�*�d^����Ս7C�_d��a��;�d��wk��*R���S|5oJ��#㷿Kp	3k�W]��2W7�P�`���Lw��si����G�-��Ã��w/�ㇱ0�9R(�|l�	���J�Es� ���c,���mE�p�:��p`u�Ov��8�z�V�]�է�V�kobG�_bb�S���6����]��Z��%��Y�$֩�f:a��7�tj�g1�m�L��[��K��|��\<�|_l���)jR+�@՗3�;�n �V:["�oV��A�;�۫|�a�)ft�O=�c@�����V^��Ȁ�q�ыaỳ�]�p�o*�5,��e\�:e�.����ie�6XB��4�S%����(�u(y�6�ػh����m���7wv��WL헻�@�H�j+2�GW� SFѬ$��>��+(���Y�n�2�.J��m]�Eq� ��V�Kt�m�4�엘�vK&�h�L��3C-ˑ�wn�O�1�k���Y�z[�O�V��r���0�hN�jtܓB�U�O�����1d�>U$;,��n]���҂ej1SԊ�:宀ֆ<E���E���ו��@�^Y�n,Uj����"k��U�k�̨vN�F��6��Iۙ��Kth�Y�,]�(���iJ�0��k6�Q�;Gn�M>��}z"��N�9t�J���4ew]*�]#P���_Q��Ne��S�rƮH1k�j�pv�U�˔�LR����S�����:���F���58��V9�k��f�+ =�ۚ�g-���ݒ1=� qݕ3�;u2���S���O8�u^�#�R�
д��m\�w�d?o@t��!�v��Bv�����1S=��׹�˔@}bM��ˤ���1u�q���
.���k+��{���mn�d.A��Xc�&�ޭ-nڠxɇj*=��F2�Z�7N�5�������0X'eڅE�9�S(-�tx5(p�T�ף�����@''&w�ofT{�K"�Lf�H�ʺ(N��4_Tf�h�LQ�Պ*5���k���v��.]�NZ���R�.Ku�QL Վ����<��X�)�t�]ý/��+�y�Fq�࡛{�w���$�$圝Q\�!�9L��I5O�].�=9����z��Q�y�R�(U�i^Z�8��ۢ����b�5k�+���O5Υ��uܻ0��\�ݸF������o8��\�Թ��eV$.���,��4�m��C�n8���7����R�r�mj�;��u28���h�V�Z�����C0^�ӯ�j�N�: �E���t��O4B�!h�3�X,a��5�^�at�������%���"�jۛ�ė����`��h�#+wx���e�i��������!�+����p�Sa��9˳�[����|8�k��Ӧup	��e��=�c��l�ŕ|`c��{����{���y�s\ۡ�N_QR*�zl7�{o�7s;�\�9\�[��˘[}��͆��!�ƚ�	T�|�^�u0v��4��먅�DH�6�Jڞ^���8^򽔐�75��8`0�����ɋ����$@8e�ڐ+�x��u�c��R���ր]�b� YtU*�i�Mr�X�;ja|�k�	��B*��1+Ŋ�ԱB]C���Q�.�z[��ӫzjFԖls��j!fQW"�]S-�%lO��L���V�X�9�C�h�[2h7�*c�q巣h�?,Ҁ��4�'ٮ�� d˧��������&��՝���F83W���4˴%�S[�X\�M�Ji�\�:^�q$����W
�a��-;ʼ�D����(�)�������>��scb�;Y�X��:���j�0m�u@�ԏ7�?F�eX@a0�vu� �;9�k�/�6�v�jnU��3fó�]ۜ!�q�:�񮭔��rC�r�M�Z��)'Ձ� �#ܩ���������z�}Ӯ�)론9%��*��	�<fm(S	m �+�ޞ�[x��'��(��%A�:�Pr#��!���5��S�ZJ@���`5�7تYupZ��K�zi���f:1u��٘���{JWv���J՚��{G`����,cc/kK�9��%)�S($�IB��Y*E\��yV���;X��\��9��9F�\�ߐ������4�����J�t�:;WRG@�����EKNK��ξәԈ�j�m��]�
�:.gtHDYC7:�������oI㭲����HJO]mB[Φt�P.����<���x"{ջ΀/�U_+�.F(t��#�%^
�j�X�����*�1�ޛp۔�5����P�d��B;��*���U�96!�	*��;E��{7�	�Ռ����p߭@�I�ܑ80��q}�(�|�*G҆��e5�:��˶ځЫ#�׊�q0��ϛ���u��\	��w�Su3uk�a�=���C���1�'C�R����c-�܅e�@��'�O��ۨX���:����f��l�k�{��!��A	D��tQ��t����_IӰ�Rc0Us��N����x{%�-r����G����G�YZمVT�ڄY�l+r�E��L���ot7*�� M�.t2�&Z�b�7��i�=ev��!wz���ʝw�;��Zs�GV�)]1vk0
�1��)�]�dqto.|��r�R�m�kճ8mY����$$�9-��T��7�h��HL���l�a_h�AwYi����֤}ֆ���1��PO�K3�5|�����;n!y:���eY�6���)B�	d����L�J�z\�oTNf���U�UUT}����#���>��#�/I�R4&}��/F��n s)	*�i�l�f��T�ISF�vΘ0H2���$�6�)茁�1ǝ*��Z���-`�Ľu}x�t&t��U��"�8:����&P�������v�ȩ�,���)��Q|œ0��O%2^[p�p�X�f5����/ �G\Û� ���Do��²��;��y��D�X�܈���M�w]����,�y����&Q�K�-�R�đЎ���W�Y�V�|�j��f��i�&4�����/���8ls�p�˥M�Gs���@�:���Y�}�QO����N�R�,�Yg��4si�;�
�qVt�1��Geج�5��'�>���OuvU���[�ķr�f_S�)m�CLT�A#wK����xR�U]%]�\I�Y��.��Z�El�#��2���©v˦6�Oyc�B��9t8�c������ܸ-�������D��k�����/�R'�SSI^��o���*N\�wI��9�*f^ܭ>���'2�CV�.��M0�k�w�Whڻ���d	�XS`��>��zK��vH��<xR�9m7�̔j]�d��e��۹5���y�o���d�ύH{�m�P�Х�(m��\�e�h�^�B��߹��^bR����d�yA3�v��L��|L�N����FŸr�͢��4�8���Ml�eQ^
Ra��VNx�|0�wY�M-��q"6R����/w�MW1�)ɉfu
\d��*��=���e+y.���DT�m��f�XXѝ���aAd��1����5Ջ�V�e�:j\M��0��S��F]@�H|��d�3�]�rт�S���t�oT�-���Kn�b�g]EZWaJ�ݺ�,2r��`�z�_NQ�m��\�Sؙ#(�{X�rН�|�}u.���-� ��gtqTֈh�7��a[1�;�7d�30�,�����^�`��i����G�^�i�� 6�jI�t��7s/�l*E˕:"?���|�<��_�J:wUM�Y�sh�hP�&Hl�emP��1�:s�(����9@����TC�i�a�������
]�J�*�M�ʹP�Chq�/f4��w����jf�f��R���H󀭬�_�}���z�^>uw��;Yӆk}�*e�f�j��4a�SS5dZ�e��r��� q��HpR�8!�J����q��W�`�V؂��"�j-J�\��h�st�H�(����w�lƔ}�ѭ*����<�xkNOnɹ;V4S����K`U�U��H7*m��k�{+(���������Y�8�xM��5\�4nh�[�t]
)��-�������ܡ���S\�L�56�r�$vW*�]G���@<J�վ[.SX�ղ��Ms��ݧB�R��Dk��ԍY���pЋ*�t�Ka��@dҧn�9W8q�T	�{Z�K1�����c*3 a��h�i��K˱}bY�Ơڔ�c�|���SY{K�ik�"w7	���wP�)�I�BM�i��՘	'�h��t0t���o륎G��Y0��J� +�5��V �Aإ����U�f��� �7s��滍�1�@��q�1��Xn�� ��}���9K���<9ݧ�&sD3,7[X$�`��O��{�E,��
��c����\k�99tB4U�LܛdϺb=�Iب�j�8;3mt�1�� �rEm�������Dt��ήۊ���i��-��L�4�\�=�}�]eů�,[6�8�vi���20��S�A6��V���}i͸�S]o�B4�o]�+N��� 鸯vuG܀�]�Z�3]$Q�z Kkd�mt�����L�A�l�" �VJ2�������]ٛb�k�2I&˕�m�G+ �O�Pג���c]y,R���x�$.�-�&��X�ΫT�nD�Ѽ����:i��`Vm�0�:f���٫��
BRL'<Ҵ>0Q9A��s+j\y���1aK�[%7,��]o$���o|Z��t'B��ә��Y�4�r̺�.�����,N��b&ev�v�7><V���(�eۖV"�����Zoy�P��
��K����^�Z��hrJM�
�9�w�Xr�Z�h���P�*n��Z�S�C���w{kj"t)����UHH�B���k�1eE����f����&q��9.c�⛰��̗H5�/�a\�)h���q���빲}��2��X���7kH��7��	J
YZe\�ڵ7�c����N�m]K�ǈXX��)�,=��D�4Uw�.|�X�|�=�U��<yԗj�s��)��D 9r�/裼��W�����xK'O��][�ZήR ���PpLC
S�%�)��@r���d�H�0֘E�����:��n�u�V�PH�Un�Gv-˛N��]3�,���|��A܉ςc�g5F�Q���a��ɱ�C���f�s�L�bV�4F��p�k�����n!O��� �0E��=����$��-�����3o:��hʻ!	ӔN�=����V��#.�l�y��Cv�N�9v�v���z��t���^�R��7�k�ƑY�3J���{�[��:XT{pI�C`���%ۆu���&;�+�7���O���v%��iS�k��P���A9�/����OV�+&Jw�K\��� +J���r�@�ӮP��Au���κ�l�ɂ�r=wC&���w�JRcObCsu�Vް�!��Nw�f�����أ�,�J�c�N\�2�\)�5����VgĦJ�&�JNm��Y6��D�4a�YyV� �VV�b��eʹQ� �LQ赠N�F�=�sx�{{SO���٬��i�ۼ�>j�{�{�m;�����T���u�������k[���MO9��eڽ$8w���+���$�\)��O6�ܧ����l�.�q�FP0�� wQ����F[.R��*Đ�a��3N�ܣb��+a{�
s9��:��9�ܣ,�����W�2�j���w8�T�T���zJޚX-B�R�ݦ�ɂWr��5#�GeN��F�����C�F�F�̰)w2F��	��6�k�`͗��V)]�nb� ��oP��Ru��j���dCv+�^;M%̥��{�Θk��z*ƵG��%�|�
e 3�	ˑ���:l]��f	�CVphΊ�\ջ�`����.Z���E��� �Z��^��A�̜���]ϸ�kj�\n�We���OH������0lL/��W,���Z�Cn���c�Wu%hU�ޜ�u�I�4iw�N�Vw���%�HR�F!�c7��ʔ�W�%�v�9]�ț�4Tz�9{)�J�<4)Z[ǊȀ�'�Y}��t7,
K�u��-����S�e�lm+̕�;N�[�M�%�
B�kZ�)��.C��j�$�U�wv��bj�Y�L[��i]�*T׮��0i�8�%��{��x�E5Kͤdi(�;��y�l�I}�'����
����r�D�[�Ӯ��Z��_M�����s�g_\cV4�!W����wZm�φLnpb���t����
�t��.d��|�4z
�Xk��Ý]cUm�:�̺����¤7s������;��ֽ2o,�v��iT}!�^�f9�7j�5+��]�U	�����Zδve���G�6�7\���L�c�k�|�#�"��緵n��Lv���G.4{3p^��'Dyg���I�D�^[.@�3V�,}\
�W%4	6����U��p䈊���,��P#�'VW(�`��⮕�5)q]��6�XAq#>V9�{7[��P���4�F����%�V�̮YwdJ���Z��º��{oU��u��g�����S`����^��{$��Iv��w�T�T� ]cLB��}[�QY��5�8[R	2�mE�j�
�K��%0o*M�Q2F����N%H���Fk(�c�Y�(�\vڹg���r���Ylv��שA���w�:�Z����]upIר�Ա���죍��t�3K{���TI�]&��me�"UG��r��1Fh�ۺp^�ݦ�1�VntY�q��*09���_`����Vo��zn#�(q<O?�:÷��ܭ�0I"�=M�\2�.�f!��8s��ه0�|q����UЬ%d�š�d׀�/�u0�9؅�
h\Rr��Q�T��J}H�L���jq�Yq)wG�4�.[ŻQїB�+�m���Y3y�fM�R�;N��8(;��㢙�����t�z������[�aYoT�G].s�l *�=����n�V��O턅uM蓖�jN,ZB�I8y4�2����Xw	AKޒ�*�`]��Fv�*+]�������[�c{)T��y,Cn���Δ���r��+��[V�ܼ�P�ʺL�R��q%qv&���g+��SEN�Vu��ω�Y��P<ׄO������ӓ;+%�����e;Ov�CY��Udor_>Ę��U����>�&bm�i�yCrnL:�ܣ�(p(Ǫ����f+T�tdw�Y�f��<0�
�\q�׻1\��K�T���Yq�xI�P&�㪛�[Ma���������j?5ii�&�>H�[��օ:|2�&�ټ�����l-FJRa�T�����.�hff�Į�[bS�jM��y݅Ʊ�5�n��J��>�oYI�����e�r�d�!�44��xl+��+��U���H�`�}B�s��ٵ�fWe<�nH��R���L^R鯲��u�:��[Lc�m�<�\�9�ad�η���	�֋uozYx�(w\�E��չ9�@`�J�չn�SYӰt�|�_*&��W\��� M� �M��o\�VM!h�נ�{����2}"��v�l�e�Z�J¡Ai��>ѥ�m��}�8�+ݍ���������.�_dѧh!��� κf15M; 9�Վ鹒���wBe��y���p��(EY�VR��:�I�c8@���W|@i:F��K;q�h�nɷZ��]y���E�/�W���-KC�DS�+�W|�V�R�y1��R��;'8됂��e�����I�������Vά��F�����R�fj ý���T�+q�.�2�힖�drR��2W]ky���u�{��uu�EȞ*��������N�D:����U=:�U��ӛQc�Z�6�2���e
f�X��Vom��duӨ��¼Y�f6�tX�"R䀨��R}���+=��:�{ۤ�OHu� <�O��m̕)2z�쇜.�^Ct�(�r[[�R�iMG
�*�u�բ��l�XT��M4�$}L�rŽm�zW�@ob,���I��ay0�ï'o-���w�F�&�� f͜�S3p	�
�kwuJ�^�K�/��-�>�\oEm��kmF�,ռ�{�݊U�N�*:u�����r�6cS�Twt�$=SY��$""�X	�a5��ڹ�m�N��\)�d����m`��f����9>�^%,�9��
��F��TpQ��%�1����,J�\U}�rEZ�8���+B�1;.,�3��5ۃPw�`�W2�2��n�0!�aK�-6�� -�ʇ�Y�Q����X�f�5��Gi��=�d���s��b�sA)��r^
Ю�k;8�	�*3iKu��C�03�E3�Wiե�Ҳ����O0ii���P��|zTtfB�w��q��Cd���wvMUfy�;MO�4,�h�s*����<iJGH���M�*oi���]�^�M�Tq�z����oIݚ}��Wjx��ws]8<���)��v��0i�yw�-9w��:��H��\h�,�˹�ҧ���?����gx����l��ɚ���],v�m��p��b���w�K��ΧF��]K��(��v�0A7f#��4[�.��ql���)�]�!^v�8w�J7n;��cc���]4S��^rÙ�S�7����7�&���t
������f�Wnaz�Ա[rjk�����v�T�s�9�&�Rh9��Z�ݢ�a5;&4��6�v�}�/u]n`E^¦��Tپ-�� �N�z�S8���gGOF��G��k+�
v �̎�q��C{$�AaMX�&���O�2��쎠��]qA��[]��x�gD�N��Ep+�f,S���c�_CR�F���z$M���M��f�؆f�	��2����%�cU��P����B��
����(�a��$�1���*���R�X�.��]���1p�5v1���\e�k��/;N���G�e,�p�J�l:gQ�T�=ð���+(���@�pSd����4���]������QʌB��K�%X*�A�RP��Zzw�:4�dý�f��5n��5L>}Pu"�5dbO\cm%�.�z����yI��,��0�Gf�\�2��eH�.8��[�R����g+]b=���y�D��!������vV�8��YYrAD���6�*4��@&Kw�z�"o�=�	wt�4�J*=R:Ap]�՜쫻|9�V�܀�\1�������{P�%�#!�"�H�h�=��}t.Dî��4Z�N���7�_PĨm�9��0	{��w�zK�ܹg�痏`�B�e7|7�lX�����J�u�z]ۻ�#�{�Dm$p�i��'�;:�#���r�Z�2�H��c��P��e���D��OpӪ���1��`�ء9�������o����K�� ���Lȸt�i��h�Fa�`��8�qXs��'�D�#�!qk`�6b�x9� 	��X^�ꥀ��S
6�Q�s��\�mէ&_jdp���y�1*p�lԉE��G���4l�ҌD�9f�N���f�Q=�ר8�����l	Ž����B�����i�(��-#z�&r0��AM��-\������*:<�a��8f�[j�û2�#��6<�'(��D}�}G�}?}�s^+���z���8�g���T�I�tfӤ�Hz;�x(�Ff�ָ�z��)�F@%�c�P��t~p=�����n��� ܈@��K��t#H��2�{-͟M�1��Z�]9��7����ްPY�jË��p�
Y�Y��u�����es�q�ƛ�mC`�G n���*��/�Jz �(����0�0fO����\����\q��U8V��]��-�Δ9�U͢2���}�P53���
��]�%]�.�t��j�I;��(ΩDC��^>��q"�K��m�.1RS%��Ȳ���
�h��ʇ�+{����s��f#�]�}"������4dӏ���yU*Np���J�+\7F��Y���n޹W�m�#z�WajĹ�KJ�ncٍ۹��Z�
G���fm9�G[�V�qjq$��8��̡m�u��y�,ܖY���!4��t]�v��A�n�ʈ���^pf���J/�D�:�K�b0��.P�������S�-�m�{#��qTj����n��V:=3b���T|���R����h�o]X��8Q@V�3�����;, +�ZKU�#�%���:\o�^e�y"�x��3�YU��¯6�!B�q��>��ږ�f���V�Ą��owf�<�K32��G[�|�֎l��R���QV�������߯�)�����P�������.�"�(���!��G2"�v0#\��A΁����wn;���wss��R4�T�+� ����mѓ!�$���t��MG9�(�B�$"!�������2���u�S-��E��D���&	��S!���M�˦�%wtr�Th�hĚ�d�FlFL�# 	w]�C0I��΂b�9��r�]�Г�d����s��# �3�(s���vawuw]&��Hw\D6����
s��nC24�:SI�D�a�0�%��H� ̤��6Xe��E���s�%.�1���\����u�D�H�2r�(3wp���u&/[~�߾������%�����D1�j�K��n�hތ���������^�a�(��㣫��%�Gq(�O,�U#��|��������EoY�n���j�v��15�]'�kd�c���{swV�Q���ۍ\���M�� dX��U�`��/�:�z���6���tU���N�@�g&{��s٤ky�MBu�Ww�ߙ�0Z����o����Ƽ+�6�롋��^x2驤�V��w��������i]����0��-q\.�b�>�j$Ks
7��$�Q�:FN�r+��[	`M»['⍓o'����)����'\γ,�k��4��ـ3F�8T/'9Mɾ�X�v�C�Ŋ���qNxXX��u4�}�5�n~�=mp��Q`����i��o��a��G��f?���'Es0..�@{�_���0�{��yLG4�{w"��k�5�Z�d#�([�O��ƶ�v\�'�IH����&�B��bԱץP�N�ƧJ��fn�.;�*���s1r�1���.R��}G�'�Z{�Li�Gá�~Eq�d��c��UVb��i�ӑ�2����m\0��_���$�x�W�!8��<;���:�����]�4ɏ����I첒�nvn�Ӽ����Fg�xZ�E*�������㮬�9��g;h���P�T d�2*t�Y샭��wL�lWU�R�c']�E�&��3��(����_F;�{�=��:0p� �G���1�$2����y����Z���J`����H�9xg�[�b���mA�cVī=S9���2�8P5��S�<�`�]�z��'_�[����]�鸊4���a�,����
�h������2	�X�[]� !ɪ@;�Fc��&͆&���
������ٰ�\S�����@~��$iFy�7L�;�~�}�R\���.�5ϣ��wJ�0�8Blh"8X�`ڪ�S �\j��m1R_��a���e���W��r�&~}΢Er�ɢ��5��@��~�'�Xu�(�4X��Oa��uX��A�|�MM��p�,�*�8s�k����N�=?9)�q���o9@�?��Ʌ��Rzoм����]iS�Z�Y�\kY���h!���#:ECɄ'[��:�m����gV�]D���z�V�S�t���]t�wB8<�늇��S�9�9�J���Nխý�5ޝ3�w&��v�vP5�*��TY�j���<a 3����fuY����1�r(D0o/�YV=�[�eo#P��-6���H�|�fg�ienM��jF��:E�sS���� �7���u�Kx����mE/����T��ٍ8{�6����5N�$U��9�])}(8����ٮG���rV��(]�V��M�`�b� ��|:��t�j����
ک��OE�S�x�y(�i�83�*���8h75��}K"�i����a�:�@o�$FD*�����cv۸B���<2/$�%�3�I/�0�����Mk� ��f8u}��d���Br�Y�5m���B%��� �A�:l8;+�}u8žs�!i��f鋪���ɡ
��鏱Ö-|X�Cj��Z��7p:.�J7��TI��{�m�L�Zx�]4�O��L����Qx`��ы�!�s�Ge�b�ʜ�����k��n������w�QU��F��HQ?`�~��2:��e�qв6f뺗
�\�\�/N`����,MBuR�� V�FGA�SǞS����������s�_��V��=��9A�t#��\\AyX��Fۺ��PΩ+��	�xEIZX�[����y"^v��O�f�$h*��`®]m����f�+�� �yߋ^m��"u�vr����@���E���!�3`H�v���<*LWܓ��As�¨���:@�r蠌হ�u���h�#  �$�J��<���;>}���,r��b.uK�V���M���
�9�lh�+35rC�V�ύ(B}��v��6)�qG�N�w�e��Q��C�',��D���֕
U��	K�
���	���3����>=�{���<�"��-��z�zk*��R.V�d����/��E��j� n����0v�A���KM��h)����n�(��{o�p`bݨ.���+��x�*�7w[�Ґ{l�V���hEBq�"Oo��|o�P�%�ߨ��#<s�Z����ʇ=1�*�*�o�b��S��f��쨐�z�:i�ЄP�X��3�,�P��-}�be�^��F���]���@τ���3�Z�e|�1��oh��X��l��j2��Sn�+)ȭ�R��ޒ���{�֘������4"�<��#�0�Ή�b,Gt�Zz9�a[l�hO|
��t�1O��x��bc�i�@:ȹ�#�g�)��23�+�[�.�w*�i�=7��Q7���}4��4���H�&G�-^�e���|UƱ��7�d��W�_�xD
Ǆ$�~��>0���n*e�G \���[<��84 ��#XD#�鷽Hv:�����h˨��x�<*�$8��<L
fb#.�v��`�h6�C��u��/5��Q=��l{O��mvRR��n�T�rd~M�O>݇���Y��=ٮ���3�-��-S��*;5�����sҮ�\gL66�Q9Ջj	K����5����ʵ)����ڝ&�f��L�֌�;Ed��XW�"��]�����H��q�+;��d��T3bD/�AQ l%0-c^^u�gT��ê��<8*�>���}-�f0����s!㘛اv̋�UQF�A;��j�_v]Rw�Z�v���&��^�(u}ӣ���(-�,���m��_9�qYJ��Z6���^�RQ��;��H��@Q�"Ꙛi<P>ޢ��?T&�y�r�֞�LWj;kv:�~ 8j���n���%�=uFr�P�]X�
Y�˃$���`�/q�Mm-�|��
�,�!�s�ix���.0���*��Ơ��wպo�+K�zc�v7v��e�ǩ�r�4"�z�K�s��
 F�2/#]����b=z����Q�'��f?���2IG���K�}y1�b���Y�݉pY�D��P(�$��l$3�m�Q����8����R3ʎ�p����>䔿�9�V��R�v��ƛ�8N�[�=W5���"��w��+!���xm�x�'�_.:�yTk=���ư���Y�V�g0��\}'$����Am<B=po�ޑ늼��*��v�h/P����uP:V*s����>X�L����cu��v���tY9��
�X��G�����$]�;Y�X��o`mGGR��+���V���1^t�#�1��N��v�=W���֥7��w��ǫޒߎ}g	�tW�:+�Q�\]8��^� )V [������g�
��+P���^��PR����a�t߱{�����&���=_�@����c��}�~Z.��5�m�ƪ���?hn��l��-W��G��tX�!���Ih�U2�C�>ոN�J7v�H"��E�1(�F%oO2x\i��m\0��_@��(�H ����j1�ȥ{<���
옒cx�t�-J`�z�#��i��q�*!��!�@۩dD�#���U��M��F��3�H1�	��k�� "{h�q)u�p��	�q6��N��/&v���u�����S�5�g���ƾ�"N� 4*205��©��۠ ����^W3�#4�)�V����cF%��=+�OJA�t�����3������K�!�סL)ڔ�l�.�� �;0���u��&�pC �N킦m��4�_#5�4}��ߒ��S�费�]�X��t+�t�H:��x�n{��|<�\�`.���(���C��������'�*�k��k����7�N���5������n�$��Ad��D���W�)l��Y��$���خ�z�F��Ƨ^-/r���(�w8x��~GK�6R�T���8�z�'W�\��Iݏ�a�P�!򙁳*چm�5�ZgJ���~��x*�V���ˆ���	����r�N��� uC�z��s���x�uD�S�]ޡu�Q3=kƘᬬ:8o�g����*L!;m�V�֪��Q3��)<��IX2f���N����f{S�U�8xkˮ�ڝ���2��'�Sn`�7��<���Y?8�y��d&@k�_ż��Y�&�����9��)�U&	�5˴P��� � �߽�V�<���J��"��=�͊�C�����^�O�����&�L�7����CBf35��+c��f�'��c��GỮ��ꛒA%cy����Xk�:��A������r�Y�5m��3�Br�K7�t�{��fgw
��z�!\�9m»���ȋ2�E�T�9VdB��鏯:c0��m\>�*��',�뢋����s�0�I�}Eh=���@�\;�S&hb�T����[#�vl+C�J[�z9,[��vb�ϧ���>�CP��"�h##�)������N�R]pS�ߖ�U�9�7��Uꂵ�������v:Ǘ���l��ү#�&��p!y5�2����v��w,TРN�V�>�,z�t�ɀm���aRf}�j��]�	��]���rr��ܡ����UBdۼ7�2q�C����e�(NM1�����K����`o�j�1�3u<�� ��2:�x��qi��1\S���-Ui���3�\���AyX�n�m��4P�P��+��� ��xGL_Ϋ[+%���m�Ԛ����h0�#�[G ����sh����+�^}�ZH��=NmLJmY�sÊ{�[
�M91�E@���F�v���1�:,�.b1�U� I��ɷnb��^�iuX�(VuO�(Õ�/�r�՘C&;]���J�s)� |id�[���J}-�|:����QU����ٯk���*�� huײ���B����V"�H|��m�͏������΃�!��Ɋ�U�+=ȓ��C��qg��HV����7�5�6d���a���������.�Fw�
��M����+���<�H4b��'��ΔK��f��xZ��4��	Up���gڊ�r�φx:�%�9�x�����8s~�c]��_-zu�C���x�{�?|�����;��i�鯇��뙁���V�؍����1k�Ʊ	Y��/=섶
癨�*!RB� �d�|O�E�^,]C������y&����a��o���p�[w�"��瘴���pؾ��9���.]c��k���{1��ԡ�U�__7WD�cA�i`e�ל���9�C�i��rwAnU�6F�;�`�
�E�&)�/!^&=�Ze��y�#!ܶ{"�p|u�Lj�1=��k�'0�7z���qUZh
�G��7Ԅ����J@�_d���Z��a�{;q')�w�ԗb4��qN��7��J0i'A����Q!ʦ��C�-�F���l׽��:���nB1����n�������ե�6 D�G����H����ڌ.z*�Җ��kd�����\������ڇ��d��T3��J��va�r��Tk��ߔ�����<"�B�=��<�n�1�ޗ�!9�P��N\S�fAS%���fP�E\��oN8��<�S��h�L[�2�C��*��0��� R%�_B��'�qp�����y��+��rD5b@��C�!i������!��P��%��WD��1R�.L�Tw`�¾��8����q�[��=f��Ŋ����\ H��)�"�y�&����r�6���6xI�K�f�_��Ρ�P>|F����!itj�p�u}z��Su�f�)b+4
@�9���f���fK��-:�R'���������Z�.�_n��:���ѓ�\��O'pV���Y���[�o�9'�O?�䤸`Y�v��r��)�pVC|^��4��*t���w�7���;줦��>�	�ut�T�=]��K�.���0<��
�<���1�]�| �
��:�/�A�'F�Y�I̑n*^����j/o/�ޘzb�k��rU1]��1@��zY&�3uA3ّ��<3_Y^�o��'�q�<>T|`�ʥ=���$�����Tk�e-���1  ��U�6��ՎZ�Y��2g�� �����sXe����W���i�uQ��Q������8�gl�~*����~�B���G,�+o�?X�'Dp�<r)H�i�"~~�o�����ĥ=�x���Y�S~�d5^�e/s�$�GC�ng�C����1�}�ku��H��I�n!�@Ta���l��T��*��k�m����:��
��u���6o;x����967��f���9�e��?!��j�S8��8%���������;y�YW('A�����eR��aJ`�z�#��F���q�)��!��`K��[7��'vMΖ�����+�uw�<�)vy�b�Ru�t%�p��y�>����x֔�ziW��s$��-zh�F[�}ϛ/r�1\�f���i��YKM��b����W���.�U���Q����L�[R���L	0�y׵�e�_α�m%m��U)�6;���7�<�ʌ���!�75�(��I����/�i�x�ہ�x�ގ��ӂ��Gb�F���Yf�Ԯ�Y��"#T�18�T�r䇹@M
�Yӳ��uŜ�#�*�Z�m��}w3��:a�S)6A{.�v�ʢ���4�-���'[��"uJXN��Kn�r�n�ީ�{d��'l����@NY�)S��W�q�GF������йr���A�s��]E��_q:�����1�Y0gSu-�|GG�Ct2��=:�}�Ml�v��M;��h��d��������y8
��yqզ
�|��D�M�K"��4]�*Xq#1i���u�A�P��u_Y�f���=��mLu��n��"qߕZvŎ7���=�,V���!�_=ꛀDS��@^ն1�d��1kw�Sx.Su�h�V���W%���vW�����̗�l����jI�,v,Jws�5%�h.ͫ�6SB��x6��e��,��
zsl8Q�\�@u��9`�܊��&���|qq�)�@s]���p9YJ�a�Q��us
��M�E!�v;�.��$���M@5юr`9�H���%$3黳o���I���u�bN�Q��t��0�CV�D�Z{N���B�#�2X�σA�\gv�	n=�ofhE>��:���!|�l�l��u*R
X5a�e����$�����e�����^5PQ� �2��O�#�V�%�	����}�^��PY�
s�vC����~y1�:�G�LJ>��,Q'��hӊC(H�옔��U�r��C��f�q�jS��y��j���lC����	_�6�,��ӝib�4sh�+Y���\$Ta� ÐZ\�p�Ś�����4�7�B��N�gVNT7y�H�ջY��	�vp텺�MuAI�;��b�F���~mBr��7�^㵵��1�)d��=�P�(���ADV���sb���յU9�Y]Tm#+nEm��x�>�F�y���Hge��0�E�wKF�/*
��y��@=�:8�r��3@�8�U�aR�b�eH_<��%����ٶ���s�0b`M"v_ul��T#�O1IY'P�4��c��J(=��!��5�c�WV��cH�{��)�)�����B���T5�VD����u��t Nat�����+U>"�ggn��It+[�/��w�՘��<̕�bcd�4eִ`N&��kfl�Nu�p�c�˸���yG0������#t�Y�c����!N�(\pl�%L ݉N�:�E��}$�(��Z��e@���d`�hsX�.�4-G���6�3�򹠂��:�3w������VE[�-��餙��ƨ�T (��332aH�I�;�(2��0��$F�2�
����!#�ԌX�E�Fhۓ�u%�B��D�!�H�wn"��"�r����Lё��!�d��CDʂ�H���#MBDL�!���؆.Wf)��X�F�%"b�a�A��AJB3`�wpLH1��&d	
77K%!���b��r��Q(��E#)��J$R&��L�`�$�$�L�؉�	�&I�$�LRPh����w\H�(YrL���$b�	$�"� 
>�>5�mv���jhY�r��[��2��P۸s�J�2цXSk�X�:OV�CNv�:��W��9.�H�����R��ڕl�:������u��_���^��{o��h/{���zEx��Ž���cs}|W��Ү\����^u��m�W.W-��m�z�?ӫ���_����~�r�������[|~7����T����zc��^	_���}�^>v����/>��~���ͻ�~}��~��գ{_����z��r��®r�?������v������/�{_�{^-����������}X�J/a���c�=�P��J}�H����������������>��鿛w�����{U�����;���U�~��7��|���޵��7�~ok�o�oKO�;xۆ�?������CQ�|_��_W��DeG�y6ASW�Y�,�F�������k���j�+��7����Z�{Z{�ϟޫ�ޕ�^��z�����m�|��}^���_;�����\���^a�r�ޯ�{W������^�=��A��)�Y'o�|k�P�p���cf�[s{m;������o��-��^����������	BW?`���G7�W�_��x�~}�z���zW����6���77��~_�|��^�6�/�����A�yBO�V�e�;�x�� �w΢�W�O޿�w^��mʿ˥����m������?[}^
�4D}� ��ɺQ>1���9�}�#�>�|���o}�s��￾W�W�-���㻦�=My(�zt�,G�4��G�}��_���W���|�ޛ��^/��������{���_��i���^�>���+��_7�n���������۽����mE�+����׭�<��\�
����E8�m^~�&���R¾��ү�:�6ᷟ�y�����5�����",G�L}�sc�"$}"!��O���}W�x��_����o~��W��U�{�uy������=qW��p��j
	�3����l�\X��ꯋ��}��ս�;W-���1_W�}��5��� ��}�~�P�Gۚ����z���o�����������w��}v�M�����yצ�/kF�o��_U����"G�/r/��lw�����>�"�_��Wv���}���ռU˛z��ﾷ����x����ߞւ�ۿ�~o>y_U���������7��������m��6���ʿW������ܷ�B ��3�������h��QB�뷬��-VG�|���9�� ïb�+(�d�i�2WN�.ó�mM(>�dTY�M���N��mN�n�7K�:p��5>Gv����Y�4�u���T�Q�D�-��;�&��S��YZk"ڢ�<�@V�� �}^���{k��ׯ]���zZ?/}|m�n.o�������|�^֝ڽ�?�z�_Z�}[�����|�龯�x�/����~-�o��1���j��urǥ�}�D}�[߭���y�2kc�[��}sno��׶��]��W�z�u�o���}uM�����A_eLUT��}/O��xUW����ž-�ߗδW�o���������F��{SZW��&����Zzߍ~/��w�+�^-�\��o?��+�����ү�湯Wy�����_/��ץ�>5s^�w�zW����[w�c��|DDP���W�1�X��>����?}������{Sv��s��F<�>-��x��}���u�o�x����kF�����W��7��ߝ�TE/���-?ݱ�z�{U˕�y��zo�;o~W���-��{����v���@�j�s�l���t��]e�>m�7���v��/��7�_~}����?Ϳ�����կKx�~�{Ͼk���Z����}���>�J�>u�sn�۟=wj5��/:���Ӻ�����&>��>�7/q��I���z��5��uw�ţ/mx�|����h��}������~�������>�����>���{o��1�nX���B�{�s�W�}G�"�ν/M�y�s��^�z^-����ۘ�� �vY�{�����j��)ų>�MsW�z��/��-߽�ݫ�����^����x�o����zߍ���Ư���=-��[�wޫ�}o��x���}�^�~�k���|����o{]�ו�d� ���d�=�������""E��|W������nU�����m���6�Q��:~���>�?}">��#���Rms|[�z���{oKţ���/�}_�x�W��������__��okO��6�AזTo�L�"��w�*��X��[�\�|�v�����5����zZ7�����[�^-=�_=_����m����z_[~�ok��U�s���������1G��}��z�}}��k�?|��}��
�d[S^��a����7.���������}��KF��=��<����Ӻ��|�_���zk�������-��k��^_�W�E����ֿ�_��ן:�c��5���گ����{��~��oJ!�#�Oί�'>R�Wq�XB�q=IT��x�|���:�~�F�A���\���tmGN�)m-7�^93lO$ӨR�I��L��y']]f���9C����� ���5�:�ٓ��M�R��R�L�Y���E��I}y�����ph\�ɰ�T�{��J�'F'���G� GͽQ ��bh�G������oO�����5zom�o�Oν5�����Kx�^+��ww��k�꿛��y��_��h���߭��^>�",� �DA����X�f�yޘK�-Q˨Ï�鏨DH�}�)��A@��^/���*����ҹn>v����+Ҿ-޻�}���/��m�{�}��^�ޛ���Ͽ<���w���x{��^-���+߆,D+1�����[�^�VU¬��]��]?�`�(|�H�#�d}��p�D��D��_������W���m���׭��W.�������|�彯kA�����{��}W��5�|�����}��j"0E���$}��^z��;F��f�:�0y_��DDP��<Lp� }}���]�������s��_�޻���^��X����O�d}�KD@ DE}����+N����;���׋��߯7����3�z~�#�"D} �p�Q�d`��m�f��}r�|�|BF�2~�x�r�����������k��y�����.~W����﹨�����so�?�ߚ�����r�����|���nm��=z�Y�CA }p�1���H���ߵ���V���W�*C�Ɂ-�ku.B>�ُ���_��z��+�_W�E���+�������{k��\����b��[�^z������_7�{��^���o��}�/J���{߽z[ҹ_�w�~_�}����>���|����E����V�w��!���m���~�^�.��/��Qo��x��_<���u�o�ۼ�_�k���m��o���x��~w��؋����W�O��~��7�żU��ח��[�&~�g{0C*r-~*�Ϣ"�H��D}�}����o�x���W����������ڮ\�6�<~_�_ͽ����߷�~W�~E��g����m�y�~|�Mͻ�o���x����wW�wo˖���Z���ga؟K�G�F"D}��W���_�x���ߞ��_�F�����G�"GܝG�G;�m{=r2�Z+ zбY�D<���5+�_�Z�q� s�����b��:}-�f �/}	�h���r�)ݳ#EBQf�^Z�r�N��V�G
�4��{��>�h��7��M�G��j��e��2����y>���<mSc'������;�t��oV(�'��˛I�|oZ}Vn�g��{Ԛ*p�$� IѷPdy�5_q.���9RY�sv�4h�p�� ��9�Дa����t|�9;A�����LZ%9�W}*c7��͝��{��Ӿi�7�$D�@���/�f�N�A���D'y}���SZh��׹J���'�%/������אu����R=�t�zᆺ�KȦ(E* �r��gcb\�M݇����E�*�����˂�	��*��;6��0��\���Ѱ�
�&����m�+��w�>�ޠ�
 F�uC5ȹ��,�9�p�1Ol{KOouqs>�|Z�;�`u���γ���Z⹜}T�vmD�Nb�����V����<�Ho��p�PT�[Y��s���ۄ*���':��4�]\��
�֢��Θ բ�^�ʀݺ*��8����n/0@2�%�"����@�㭽��V�^=a����k+���C�<��W�Q<��h�ƩH�i� �7�uK���͕=Q� �*I�l<�#��\4k[_tF5�C��'�D��=?\�|~�9O4X��ت^�� �huAo��s'd*��-���g{ގ�{�y�¬s �o�o˺eX��uh�uD�/����ö.IO�Y[{M]�&����  �:��+<����;±�e��ZC�ûN�ݛWL��mnC9�Z0�	t�r����}�pM�f �
��l�ĵLj����[F.(�$�D΁�Aȸii\ܖ��/�E:�EIa"�g~����C/��Q��6��8%��5mS-N�����Ε�A X�b�]�EW�J�����E������.z�0(~ވg*w��S�9wV��<gj�&��� r�3�H5 
���'��<�1t���Ŀ.F�X�m���x��B�����m�ĉi��鸣L�I�i��H$�@T|e���]sʏhWpBS�^�t�K^T�nK=h2�����&��Z�^y�QAWqtH�'�3��;�S�A55z�a��sYК4'�9�P�9T95�n���``�`���Ug��T�ί�ȋ9�P�s��\����v�f��4���9��)�Y��{���K� ����n�>���Ӥsn7'�����8,Oҧ��r�`��4�;u6O]�W^���s�����d�oح�kE��!�����Dc�T{B�
�t_�L�Y_�Gs=/�{ �A�t���P[����f(/�nr�g'����o4�q<h(U3�XG�Y�t��MB�R��פ/��λd(���);����X5ƋJm�;!�x�{2;�탢�Ҍ��˥k�w���3@��Q�5J��ĭ�Sዌ��&�[��xp������^�i�tc�0N�;��p�m�jI;C'jo�W��`8������P	;�V�����l�s���4 �ǵ�W{V�J��	��#�E���@��X�0SX�J-V�:�g���{���%u׃���*O,�{ma�:�,5v�����Crx�V�fp��d�o��
���0��/��\��ULC�ٍۏ��C��þ���-vֹT��jj�W���/pOPJ����q����9ᎃ��%�F�9l��j��S�OK�����u����{y��`�g��c��9��@��U/���&�+�.���:c0���Z���6�^_s	
���`S���n)$��΁�C"�aOn�rc���!}�����6Ϡ�����
1Q��G��p�v�ʔn }���
�����B���_����h�߶��W7�F��~�w���qΞ`o�{0FQtP����  ��>�JU�lO�SOc3�p�nqe��1�������#��h�yX��F˚B�;�=�}�z:t5]zwS2T��r��SS.R��ڦ?�a�w �F�~�Ԇ��� �D���ZՖV����5��j�w3ɖ^ �zѻ��z%���3-���ٙ�U'6C։\7�Z�H�x����0%��n���V2[@�h����X3+������Zն+���f�̡{�/�|3A�_r�h�s�.m�:�):�h+&d���j�=Zw�^���D�V=��xR�P �A�i�=����>��|eP񪞺��8֟��r����OPͣ^�����8��D����њ��ҋ�[�۞z�wsj���(iί!.>bdu8�3@ɖ���B3��qs9�=v�v���|������^�=n���%&�`a�.[{�Z��Sa�r�p��f��AN���Њ�q�"Ola�P���zb�ܸ[�F�m�)�Y&�������IVw��!���T��=��:C/�FA�@{�Exj�A��
̯w��{�����T�X�0<@�c��j��@τ�����1����/h͙C��>rm���rxxXE������g�[8/��+�0S_�r��Q��*M�W���DhꙷIc���l���͈���P�6�Њ�R�ɠ��J���<�H�NkA�U�)�f�;��g���U�P�w��B�M,�8�+���qQ�$8sZ�=��ϱ{b�e����*�^�t�]���^�tm�K`秨�7���l��MYAue�ٛ���^���8y��������o37̗S'����sW35&���N�ܘ�Lʱ��@��U��jZ����sZ�Nĝ��ݺ=4Ť���ﾈ;��p���������2��L>����L��p80q'����q��!P��Ԯ�Wn$�s��%S�GYb���=����c����Hv:���ٹ2Eԏ���C���G��wxr}��_Q�[4�TI(m��)�d�?#l�Z7�~2�ѫg�/-lk���^�~�S�!�U$�9�tzb����C�n�1�A7��Ȅ�4T<u����lo/X�N�ə��6=~�0� Tt �١(��
�G�b9;A ڢ���A�������ws������+�N�O��ܑX@pD��.��i?�%]�d �!	�d����������n���1��@(N����:7�#�j��X��+��W#Z[��n�IlsF���u塑�UьE�99`iy���	j�����a�
{o�����z�Ý�ҳC0yXc��u��iZ�E�@�N�e�k���h�PU�L��V�R�__�r�}��{é���� ����gi��kտmoL=1k\W3����϶�F���5��Lം�r�0X���=����020�s�tVq�+kI��R��v��1jn�,M@G��ԱL��ɽ]�����M�ݭ�Q|���zbOVkq�BÎR|���f��9q���W��4� J��+�vg4�%uyyz�%b������sh~�����%�56�J�3'��LeA�1'��g�Qa9uX�=�Pwѷ��[�d�)�9;Ú�t�d��zӵ�.4��~�7n��+8���xn���C� ]���mE�6P�]��8N�޸�F�����q�k��k]t�E�%h?+t0֡�:.7~�Ɇ�q��c�QT��z��̠��rsZ򘎹u�F�{�������B�������^�{�`+�2#���l5{���Pp�p5�(uƗ@`Bs�'pً�j���V��ʶ�]�b������o*�_ ި�$p��Ñ���Fk��9�e�ϴ����ڸb�L�.�f[Ϻ�6��v.|N�ea �N�!�%1�S1��+U�Ҕ�q�]�v#��=�{�SVD�LU��|K�*l�iN��7)x� t�
 ���'��塃9��W�k���JA隘�z��]�n��n���qF����,�ȈW�@�$@_Ǖh򿂩����d��b�=]��.e�� pi5lay\�g��M6�@��cȫ�Ȑ�Gq��F�)֠`�����E�5�;�̇^p��d��[�+�R>���5��ǌ��8e�M��G��}���0��A<��}$[:3@$���̧�fj޸�+J��u�[9)t����Y�D��A��2�	��܂�Sm����U�v"�ց��iB�/�v��`����������սP�m�ܚ�@����5�T95	��^C5��!!;��*�u1!q� qe���P�i�ª�����RS9Gb4�5����%�#�L�<��9�u�WO�*[��
u;|��u�C�K7;t���vh��>g�RӨ{�q�O�������Je���5�;�9�%5h��5G^��N!�@�f�Sn�F��<)���n��f�l��G	;e�䂎`�`X�w����Omc>�Yz]W��.��/�H�n]z��Գ��>�9)���3f����^��
�=���^��dA���ԝ��̆����3;��J� �@��|�T���
a�Q� q��lgʪ��p��ҞN�淪A�����a���ۏN>u�*o����pȈ�6������; �1��B�r��"Z�W����Ӻ���"t醀��A.�iw*��a��ª �K.�e#Κ���d��&�5�7)5y;S�t\':"Y����0P��s�t��E�11R����9b�D�d
7�'.�t���Ɠ�MD�c��؉=C�75�L�����31p�IwU��/9ث�Zt��P��]����3J��#+\w��O�&%f��0VAd6:��:�0��J���{��#��Нa�gR��n��L��pk/rt���@OĐ��o%1oX��|{/wR�fI|k1J���rg8&��^v5��*WZ2%�;Cƺ.�l�}�r�in�2�Az&m*�S(!�+�'�JΈ��¯u�X�7̕�Q`49�$�-6��U�Ԁ��x�E�f@,��y�εۯ�t)޻��3A��sS�ٻGy�Mn�Æly[��E�Gj�!�q؝��F����m1e(���Z��}�N���K�b�����r���L����\ׇ�H���缸Comb��	ڂ�n�E8������1 C
QR=�3)�P+����s�Nv2���n��0HJv���J��R��̦�b�$뽙�S/v�m�q/F�l2��T�Z�Z� ^nN=V���h� � ��2�A��`eu_!�\/v�lNh�ް�H��,ƥ)	���ɤVGEjv�m�p�Y����K�M�ܤ�P9��\����i(|8�j�Pt*Yg�W��b��h�r4 �׃h�8-b��rl��O©R|wM��\�e�ͮ]D[��4���/�`�>غS<�6)��<�X�ջJ�*�"�� Mc��q��_CN%u6��{�1%ܖUͤK��Yf�l�5�W4�ysHw�,C��GW_XrU���C�O�����o��KS�HK�-;-����S��ЋF��]ү�QM����f������-s�m��8�����A;�,�����X��/���Px�u ��eKy�y/M������Aǀ�dַ5�]ߦ�wN����f���f��R}�S��m������HM�K�8s�B��9�u��a[�9fFw-E�����nb.���t&v��{[�v�Bl�w*�Mvs�Fɮwo�kqV��V8��]��+��N˦�F�"A�䝚z�q�Y�-��cX�v﬌Ԥ�����5i���"��S2�c�t���
���<ޚ�V��	�`;"IS��v��Keb6D��
�9�s���Z;Q��.�����]�������|�f���O�Uk2���Iҟ5+���]e� �W���}����Ù�&�KH��`֓�24pJŢ]�L���Ɛf�7%?��׫I�8i�uR�Ӣ�ș�b��Wj,v^f,/[&���v�H�wvf$�:v�5I���AqZ1foe*y/��I��9֞9V<�zn��YO*%Lׯ��팂�^�P�ƋS�ܽ�d���pST�{��lĢN���#��r�s�>��>�mR��:	̧��f&z�S+����am��Q����3)��Z�'Xt��	�{o�{j���o��֘�v���k�o�ߟ�׿��~|�����$FB����!�˓�EEQ7ə��p� P�d�QHc���,Q$&%�r���(�$�+���`�f�$w\�3AM��D�I�Lll�4�Ja0�h��w"a,��	� ��d�C2R��))�1w\M���;�%"��Đ�';9\��$Fw]�»��10ɛ#%),�l�h��`�w)9є"`�D �&2�ݻHDL6R���.\(L�f��Q�Cdwve�¦wt��$�"�75��M�Q
DA�v�Q�e��D��R� $�t�1!l�)�$k��9Zm���ҋ�v����>|�g7���{�+�6+')]*�ϻ�ך���h��:u�w�"�)Ic��Q��������\۩4��0���� ��b6� ��P8�_$�C&g�<��4P'��bw��`��쩌�5���9�Ø�p��۸x;*Q�G)�1�'�P\�E:��|����(T�H��ˊ)Tp
��Ɲ�n��]&�:�s" L@�A�-��2j9�Ⲽ���Bܺ�����_�{�낝$r�������ۧV ��L	Vyx�h!�R���N-�G�2����V�3|hf�
�u�C1�E͢VX �8le=Us9=9#V���}wxX��t��R"u�v/*�A�C��aL�����1�:,�Ւ�>�Gֆ��UG\F&E�G*@��c�0�+��Y�Jk���]Ѩ1v����f:����]�æX� �\', ��g���ʁP�\��s�N����r��
�/"M(��Ύj�g
U��X��C4���sB+�q�n��� ڷ~�r�&���S��`6k6	:��u�Z+F�ϵk�
�G>��b��T��~�f��쨑��D1�k����ܢ���i�j|�q>�:�;�2׷��Sւv�;V��<�`#�
��X���i��J
���xy�4o�}aE7��^j!���<~���M��N�7Vg
ڇ�G2P�[ZM�x��k1��^��H�[���1�D�d(�;e�QZ�+���UW�W�˺S������5�����
�_��J�5ȁ�Y�m:�#��u�t��Ft�W8\-{ܴ�Ȼ4ǫ�xYj����J��n!�Z S_�r���x��尸ڂjO�򳠧H�dDۄ�x���h\n�U��tT���b�C׊��*�sjx�c��-|'^\i�6!���g����YUǬ��~\W�s��^�t��h�������*��C̵x2#TL1���}��;�鸔�U@�x������hz����3��w�;�����2M�Ϡ\�"��a�C1��t�oz������4ԕ�@���x�ڊ�}<���9�*� ����	�ʆx�}rmҺJ�u]xN9��Z�;���AWB����t�M�;�dH�l'P+�c�����u��Kvٌ�����'1�7bU'1�.1,�k1��UvD�v���%�����f��\5Dt��TG'h �^�lr�ﰺ}ˎ�W�����'���bۺw�i��$�(��F34�x���P#���."v�%�±�/�����T2e��Fxr�V5X���(i���q�z-�j
`;�R0A��1���=\8�j���@h�@8��mI�'*$hS�є4���J��6�L:����>�����<Bg,�]��LS���0�[�q�EW�}U��Tʓw�<z��?�~M��,y��&�>�Z�A�j�ǵ͗u���A��ds��et3�!�n�Z���E�,-"�q��P�Vϋ���6j5��
bt�^���Qf@ЬW�RKΫv]��͎ V*���SQ����6[~�����i�4N@���W�ϯ��e�%�'��^��iɇ�-k��q�S�1���m�I;NoV���EV>��5���b���6M�b�'��26�|5�4��W��j��|�|��pͬ�ӚE.u�ai�8/�� ̳0����E\�E�60�.'*w�L���u3x�R�A�7M����5�����s��mR*,�+l��$��X�$sSՙ�i�%�"��� `���nka�1K�5���1��m�L9g��,��ܾ���#��dA}��#W��BC���]i��Aͧpً�Z�7m𿒜�3��_{P���F�	[����7�˺�kґ#��#�ģ5��ӑ�C8.0��+�K]u���l|]-��^o���ۭ�����M��r8+Z���d�.�Y��ǒ�=��ϡ��v�>f��Ѕbu1;�GY�� ��w�o��*�?-Y��˔��Vj��E�נj:��꺎�uH�����sv������+�x�~�����Vxރ^L�����pJ�G�}|Mlvrl]mN�����	e"AD�
�.��"k�w�q���A���z�#�4l����zQUf3�p_��*�!�ܩe@�:| ��}5��v9�B�0�i��W&���';\�6y|�+�cS��y븝2%��,�EF���*��c-�u��EB�_[����*�GS�� b��V����ŋ'a�Z�w�dHB���4�Sf��i� 䨚�X�p೵!�;f@����5
�T9)��[aC N����O�b#�vDE�vZ/i8��(���Q�~��gDÝ⾒s�tQ�F�t<��@N����*w3b�u۾����|�����(��O�ªQv�O<��4�;u$�l���EP\/"���v��3n�N�m�*@��vU�m�U�:5�8�,��L���{�{�஧X��(�����һ6�u�u�:Xo�5�Tl���k�סR滯]D�՝yWZ��1X(?�]G��S�ȃ�����\��n����o��[h�sD�(V:y�0�&#��q�xU�a1�H�K㕝/`�r���Cށ�m7��O���;so x��o����+�teQ͢�IY0��i-�^�+��'a�o.2�x�m[Sy�S��3r�ڜ;|���G)��S�� l��]BҎcvԹ��}�U}�}U�w�p���u�����}lgʪ��ja��k��
ڞY��ǆ����a���[��_r���E��q[U�DC㱅��%&7�s#!U1ptc3b�Ci�ef�>�q�Ⱥ!�6�vNt��<�1_A>�%���Kܪ����Xc��BYtm9l����+w+;�E��	:�!���1��(D�q]$��D!_L��m�tY11SG���9��4E*�x��z�-��]b�A`3��j��Z����1�$�t�`��UIp�L1y�mӨ���-�ױ-�EUa��*P���,rۈsn����R�}�L��	H"^IN��w8CjŨ���Ͳ�g!}k.*�+�]>;�'@o��#�0)䗖� ǻ9�/m��\�ۤU��nL.y�Yaq�[�_�:H��\������6�F�:���ڐ��{��E3��р�Ǿ�YN���Ù�%ic2|jh0�#�[G>.c�xo�׼O^l�T��~O"��]I������ͺA��:ꆻ�x �"4�x�쎅��XKх1C�Fse�Bj$Q�,t
6D�nP'c�pY�t�6n�ƞ��ܗX:��w���P=�X�|9�Y�\Cx+�͘%��s�pWJJ���4�F���;ݤj8U�e�G)�@*S�%)�1ʏlP�Q�����9Ҧ^��/�Έ�V��ayQG1G^���oq?����>��VͧK�1��Q��s�¨��N��w���I��:�:S]`0���5t�]3ካ��5mpu)X�UT,3I� ;�g��*|�\��f�]���|dv�M������eoWEx)?G��n�����cŏ"ŵ�4#�\ȇē� �|^����ح��s���S��	�en��,XL��� ���:�2���m�^��s�ջ�V��~ÁD�)�ަFB��j���X�w���t�Eo�g��N���K<Մ�'N2�]i��0ŵ�t�,^�6~DܜJC�Ҁ��}�xв�'P ���ߧ�=[M�C=����b����p�&|o��,���B=��A��QSU�h/x�S�r qJE��w-��u��D��1_OM�Ŋ�j�ӊ+���v��V���d`/�28u�����Q0�_���N�zo�Y\@8
5�'��G=�vCzo(�g==�]��
>@�֑�%�J�d3��M�ޤ;>u��:��9wqv2�x���'=X�w\ɹEų'W��ZO��������`bx��T6R�b8S�|/7-.��p�����M)㣼��{��ONe��r�"�[gn.�.�����w67\Ȫ=}��a>�!w�/�"�s�����P���I�h���N���?}��G����vݧ:h�;'�p>�4j(��E��q2�a�S.9�������uk�=�oS�����,G@Q f�J�T@1����B�=��2�6a�z^��b��L�t3��RF�c2�W���K/�.�@Č;U(�\�U��Ÿ��(A�U�G��\������4GJ5�5e����M6����(��;\�]D��/�fi��uZ� ���]���'	�@H�J�pp9��M��9`k������B��G�%�ڡ�Q�w�0���o���!R�Q�"wV[	)�1|X!���4����\a�?5P�[R�1�r}�7i��������,Y���<��R�M.�۾o�}� ���6��(���07����su�Z�MJ��S:087(u�������G��o�x����k�)�g�w��� ����m>wS����EDcN�ٷ�I��E�b*q��8M�@M��@�q�����.�	�Ce`���W3��Ky��*���� ��íRe@xz��Lm;���M�3rI�hSk��	c���'O �è�f*��C��a����I�L�.>C3n�(�3�h}���h.<�B
7)	�.n}�[��(ɣ��O+0�R�s�F���SVQ1�N>����Dp;ӪlDDDD|.lb��f��kw����'�2!�F���ۧ���ֺ����to�K��E���{ՕH.�@���`@��\���򘉷쁆��~�^�"�na�KW�I��=�Z�k��Z/�3��I�Ƅtf�&X�
@� ��;��\D�Ln|�o�2emM���Ś���w{4���B�L�$Ɩ�^�S*�C�4|:���+#�����^��O�l��m����ױ�)ʇ.�BoN��j����?�.�JbI�g~V��(1���)�lT<kGmk��4��r��NF���~�N��v7�D����� =�Oh+�<���s�57��cĞ�<�������N�����t�Q�~�N`�P���4���R�(���;�p��v�EK��ۀ��ՠ�3
0���Z���U��0���6n��r�8d��k�<[_���c9]�C�I��^D3X"�!�'T�JO0��}{=u-n�����U��]_#��wM{��zf��ox���Ht=�Yq	��p%Q�n�>ܱ�_R��:�L���U$0(��Nr����`�%��l�b��>�FY.zY������l�����]�{�PS���St;Y��b;C)��fw�0�x���|������
�F�Z��s���8�ȞN��_�'ʼ��կ�s!G��菾����g����;��?P��-2�>�Uyn�;ΏyKO�{�u�];����XK��3���˩u������{p=���&�"U��������
x:�%�K'u��9����C�J�db�@H������N�u�>jI;~�s)0��R|���N݇�st�	�� �G���U�~��n�S�<̈8m���N��f5ú˳���e�^	��9&l)��M�TN�Վc�jg�"��By�����N�ޝ�I�����猢HX�7rig2T>��Q�����-�R�u�k��F�,��ޖ�ӛ[7M��Wc�*���R_T�]_d���>�A��W��#*�W���eF�㈖����:�Y.��/�U'���a\����W@��$9�2�C:�:v�Q�/-�m=�+9\©p
~;��rR�]R�8;�@h��?���)<�b�i��黁�R�����
�f����x���m����k<�}���W��洨&
h��N�_���F��^W�sa�{�23�Zӱ,�N���_t'na��x�$Mύ����ە-7�^��%��LV����n��w*����uT�<M�*��3MOh�"gF�N>�����㦳�w�䥐���<���y5�K�·ې�f��r�%�5�zϥď&kk�X
<��3޷y�^4�[]7l�vn��)�a޵��
��s&aի��0^5TƖ��WN\��h�#�MJח�}=�r桾��b��f.�n��70'�w	J��L��!u^+��;��;줞&v�'��8Ǽ�������Xn1�W�Ts�9�>W���w�r��/Ce��sk}�Y>�x���X��&�]�7�.3欞���k��p��Q�Ս�:�t�q9�oVLeջ��]p�Ú�-�;p��G8�O��gT�Y��bX��Ѹݍ{����So*{���gO����yFoE�}�7Q�߮�'Bc��T���3y��ۦfq�eA�Qf#���u�����u�������TF�B���;A�?w�ϗ�[��I���ѫXԯs�%��US�'�����N]3#��h�٤J����Omꗓ�'bjNs��Y�3��}���]��䡵�\�x�(�W���0i]�k�:(n�a��תa{S�DJm��`5w�f��)�g��
�n�������d�mL	m��X]��j��V���VZݷS!� ���>���ٸ���ĜdU�'�;ev=y�}N��k�Q�[Y�"���+�FG@�U����1L����&Dp���5V�x^�a�x>�a�3�!l�19/!4��E�օ87�M�N�B�B�����q�$�Or��t��6�lx�F_w�y�]4-U���*�R�<b1��_�k�T+��uۭ����;W��}	}׽lve<4��^3A�/6��4W����c���K̷�3�#�F�V���k��5U:+����lvh�Ol���ib�lV:�5��=kv��	�ӣwհd;�[0�Xt
ň�+s(���7Vnf�a��i�1�7ma��<�Q�g3�e�H�XGYd�.�7^I6���:���\��	ee�+��RSD���W9��]� �P���©,��&�pNY��9(ݔd}Xr���݆��qYLHGt�q�f����M�p��B�}��u�3Z'"�t��pj@Z�V8T<����R��[��s1�o-s�릌�[�v]t_��؞h�������e�4��H�
�Ԏ7ۧ�c�U�ĥ�Ev��b��B����i0/�"�.;Ƶ���ԙ$��j�ۦyw9rݽu��sm�b����kz��|��v�I��kD�f��{�_cڶfȏJҮ霮���Z�wqH�WW&�QqX�{L��iʔ8FP9#;�fl��&V��3��[��Z�����5���mr/���oD�od�����;�A(�,.���l���cO/a�ͬZtQ�wx'�E>��b����]v�p�lb��&{z�N���)�f���A]x7�uɤ8�Qt1eNZ*J]xi!�Ӹ4o_Q�aꖱXn��r,�L�(.'d�c�pi|��b�o&JJڼƑ��=R���I�v'^Lظ����f�q�x�Yր����K"���&ˍV����7oVaj@크*�.�FgVM[(�U;ߑ�jH��l��=Ǣ:�ְi�3�*��\7�@5��Q�h��^���*Sol��{}�!9�VI�j�Fu>�a��E�]�o"��f0U���E!����s�7��$�A�ʚ*<�7��0b��"��H�w�17W�eV��þ+ B���N�i�������)Ո=��<khf�N#5�2!�I�j�(YXu�B�5��a�T�����s��sNmq�"���q������$E�ٛc5�c�[��c�>�2mպ��&az���;F��2�j�X��K�`u��w�*�Α;�xR@���A:׹ɻ����垱`lt���Ҧz�_D����NU[_ T
@
(dē$HP�1&#�42H�)#0f$���I	,�2�2Q"#$�M@e	�S1#$ ���F��D9ĊIbCF2�6LFb�2��&`Ȧ$@�9\���]�"$20�%#P!���%�� 5$�!�����!�Ѣ���%2ws%$Ґ��"*"Ț�h�1A�ˢ �c2e2�����5	�d(���a����IR�4�I"J.�,�J�	d��Q�ܻƒ�%0B� �������bGF=�g� �%�f��� _c�/�c)�LT���|���.T\���ȡ|�gީ���1tu�DG���l�s���;���\]f/L��]'{�s5c9Q��Tz�|�o�X(�lS�m�z�M�eD��'9���jWZ���r���`ά�y�ݞ�wW:\�QuH��n��p�w�<�m�i�W���.���ʼO���V�!�P��RS����ʚ�y���8[O9k6��Z�TQ��a'�x��wd�o�ك�b�?�I��),!.��vF����#z�,^X�=������E���RcL�~Ϧ�v=w�m-�E�c6�'f��v�Փp�s\'�*3���f�L�Q�.�`s�+]�]|Y�kp�0s�qeW9�i�|:�ᷔ�>��q��5Bo�|�ү���e!�G(۪3/�NwIs���@n1�W	�����C��]3��c)1��5�.�O+��<��x�S<�;+���>��O���o'\��3&B$�z�="Ij�نX�od7�g���
8�|7L�eV�	N��t���oL�E�����r�yW��$������Y�@��M�'JU��c�:Ƥ@����;�=e>C]�j�{ȆN��+t������節����xW�]�6��{0�sj�f��q\9���"��^	p����ٮ5EtnK^s)�	[�%��U�	O:�Y�����'mƜ�\�t~Y6��~�\���mw�-׶�EC�nNUE��qTꈌ�ی��\2�5&�-p�V���y��>��cڞp�^�^cf��,#���I��bVBJ۝Ë�
^�����X��\B�o�w��� �!��1p\/��q*Tc����yss���ۭb�kg����x��=u7y3ڔI��[�D��q��¢o�Nm6�姼��������;�ڝ�'�.xߎ��\Ie�W*k�M�놳������T�U3K��	�m���fm}8���H��\���W�c�{����˝ֻ5k�q�_<��}p��-;Q07�Nہ��*uU(86kWx�^�M�d�u�t��Z�R�4e�k~:��h�e.�u���>���:`'�އh*}j�m��[�v�8:��#$��|U�
�0+�Ε[�MP1�R�U�Y����.�כ���&�b!���6�h���֎{�Ol��菾����h�\��Gg�=�)w_����C�r�]"�/W�O�4t��Hܻ9k�b�s�{��W�d]z<�-
��҇Z��<�۸�6�L�7S)6�+D���0��5+s.w�V�˜�o��m�pBʑ��kO`�;�7�=�7ְ{��:�'?��T}�M{�:����s{�fo]J7N`�);z�g��%��us�V�*?o?Z���hv��z:����Ñ���b�oing�L���὇5	�;\�+\dK�'�Rځ��^eD�z�me��6�ҋ�ƃ���i!P�=Y���z�Wދ�:��-󅺪�X�JK��>�:�];�ר��^�������*��|��r��=�N�r�4n���s.�{um�j�JK��79_D�Q�v>v�y�/�y�q�8T��Y�Ƀ�������7v��K�v��*p�}���#
����m��n����/I����d@�<�+�՝mP�i�W�t��Q�]��l+u�_8��<Dx�����\Y>��W��2�>�my�n�0��a��י�k$23}b�4����aN�;i|2cBf˹9Wf�/�A�?K��ᵓxD -�uv�m������Py��<�/A+�/k�ƶz��uAWU�I}Q*Td�����d�f�ɛ���\)�Ɛ�[i���mŝ=-{�|/���=R=�/tC�N�T��N�N�Uf�2��(o.1�ڈm=���Wp�\�������F(�{��Y�������=����:��e^�R�۩�6�u>���>���g{+�Y��*�8��-2��y!.�
�n'���t�<�7y$N�r�u5��u����!8����al�n*���@W�C�y�gX���ś���[*�ߥ�4vC�=�#H��R����V�˚����7;s�z��|��TO|9��w�WJ����%��Nѭ�MN��{X��N�p#�Ws�*R$K��u<�D��q?'��}�>�An^,[f�]�[ca8Y\fZ���W�J�c�<��v��C�*���Lʡ��7���f��6�*7�t�s#��}�ht����:��R*ҫ��7n���c:ۨuyj8<�ލo|w
l�ϕ]�*-B@���+����Kjٓ9��m����q�h�`�Z��/Vܖ) ����=�c�mX�˵)�j޵2��d����}�9]���^�̩Y�z�.if�Z��[�v���h��t�4뷮~"R�T,���ز�����f�闗��;���;��r�j)�toyE��Ͷ�Ϫ;@�������b��5{�����N��m뻹L������=i�6߽�'沗�[�y����l)�򵎔�s�%a�*$����x��B�V��Ö�"��.�S��k'�*�u|e�c�^\��T!���ߺW�� �{�0�M�������{)�M\�DW�W	r��j9g4,)�h_)rmTK��wn��Byx�떞�AY���A��5�M��g��B�\�9k���D���ʚ�1'��X�m<�J����w[3�}
�}�9���J��wRatd쾙��a�At����ꛧ�5s�=9R���_r��(Ϧ�	�^~��?[X��<	�eL�pJv(��0U����k*C-w+�*&�1C�&G[�cX�ٱY�ɭ%����[t��zL�-Qv×�2�s���M�yp!դ ^S��|�^�cMQPq�!�0�
ٲ�)���۝S3h� \�gI %k�����荒+vNkp3��:�g,��x�T�eVG|���f�V�6��YΉ��ٶYJ�Vk�;-�6��7��hSo :e�M��� u�nV���:Y���/T�d�bS�w_%�j|�n1�p���mξ{4UpVqne��|K��z�rqjJܚ��kOѺ�$�U��q� ���=�4��;��i�^�����n�/J;"���N�j|�|��z�k�-_�5!C�p�1s1�79P��Z�v�-mI����q}7�ӓ5�=G�:<������k}�˝�s���d>1P����~�Tz\�XQ_��y/�̥����b��镂�>z��Ƕ��N6�N����j����3�fCޫ�Y�~�|8�qХ���w^j�kg��x�2W+�|�]�pZ�N�Q9=Q�����E�.nq�}K��kV��_{0��2��՚���t����q���������s�g�[2�F)�4�=7�x�>�����q�k)ǝ3��Ӈ�LS�"��s^�T9����>D�7�_=뤻./��p�( :MזH�K>��{���:{��\#�}}�D��vNt���V ���]DI|Tr�/�(������G�X�Fk�5R�#���:���\��v��=�/�¹S_bo2�[<&�������c�U4�ji�6�ep�'~��wz$��gm�}*��R�'�o
��^Yik]��6�qʈN���]B��ؠ�dt�t���%��_
p����rsj���1�b�	wB������p�E2Z�ϷԋC���mk���9����F�����١W&��޷�`��yӑ�B'7\�ѩ�Tl�uy�0�MJ��Oo��\�M�w���O'÷r5+��z8r�\�Q���{�<���6Nkw�rt]�߫�{��:��eN�_J?g�Q����V����Gl��zRe5.+�V���!��t6�%߫�4�8sI�;Q�r��C�'�Rځ��藘������
��0�WX���كYD*$�{��[s;�ǽ�Z���b:�J-��Z	L��hCc{q�w�z�Oj��%�ݼܖT�����GB����j�sn(�i�����.�z�;a�]Zu�:.ù/~��5g�
%j���[�}��f��P�,�3^[��W�ҺָsP��g9��'�e�7��:����Ƨ<:�}���CgӼTY�I�o{���x�c�ȫ��ߡ���2�B�҅X�jB�]��3j&�*R_b���ڙ����O;�X�"kj�՜�Ž�f���仆�n��z�}k/��)uD:��OV�)��̃�Z	���;wq�ݯ�w�m�ƶz��pU���>����~����L�V��9��C�CHs�M�/�t)Τ�K�������yW�{��mN\Rfpcz�z^z���[�ҽw��p��Ol��eoˀH�	קۖ���� ��/#����V�j ����[c���7-�QG�,��	��)�o���nt�݌���Rym�����t*}��㇌��g1Rwԉ>����̮V}�?��֚T�O��g�u\҇Z�Y��7be�I:Ƚ����K���{|ÚM`��&��c8��tj���Pt�Ԝ�ټd�i�T��3��4�nJ�1jIv����(C�����on�g3cf.���\< �ce捑�F«�Y�}��֞$Z�W�B�U���;��ܽ��Vf�=��b�!;�����*�ȏb�RQ��^(��<�3��O���P�9ʗ
e�}�.����o�*�+,*�sY���fGS�p]�Üw.9&��v��'��q�fkr�e����oV��_�9����O4�M,p�7�4�\sVOv�WeD��G۝Nyug��z�TrA��3��>g:�Z��E�G[8��2�na��c���d=��M-N6�ؾ��f:�yR�fs���}2�f��*�Σ]�>�l��:�?zӟK��2��~����j<ꋣ�V��U��T�c�m���6w���v���{���[��������nr�C�:P.�8��yF���c�:������>y���f���t�ݾUs�'���-��2�q7�{�(����;o��S�L�r��Y �A��U�y�a��㵂�<!/���&�	���qw�ת�hLzPƎ.�e[����:}������M�PU7���MШj����ӊ�����an���ܰfؚ���\;���9C�F�ƞ3������K�N3�a�i:|,����++z��D}cUgm�l+��v�K���~�݁�tsn1����+9F{Y�ui'�6�t�\���M7�);��rR�/�¹SX��p�,p���boE���:*��c�S�s���;�h�_r��w
�4���+(����i�����n���7\k�W��8ͯ�3�K���캏�܄l%Y���+�6�GM3K��<�gE·�6�;ש�lۗL�)����4�ev%�>�=����� �ݼ6�A�L>O��o���
��@t�|�\��B��X��[)3���ֵVz�6Q�B���Sx�K��&�;��8U�t�2�E�R�8����Nq`���cf�+rj%�O&n��ԑ�2x'Sޭ�ϲ�sB��x�����9���Vԙ�����W<��F,����s�/{x��KPyХ�!�.�;MNS�uQ�H��3yy�eFs}1�L���ci�,��B����@��A]�Z�X��#�/y����޵E�XA.af�-�ro��j>5͝u���Cֺ�{)⌾�o3�j87t��j��>U�gd*w!SO�'�~�/}�DA��%.�̮��IN�e=J:�A�.c|�8����]B4V�r�<��T�,i���p-N�;f���>ݝS9@�љ�ih�Ecc#5p�P[�(�J-2evr�g-��x���s䣝����{3!�/-7�ؤ�h�=6.���[7�6R��ih}xa�il��Շ�D��Z�r�Y�;+H��L}s�K��L3����{���tYQC����Ս�g��ό枽�k����Z�3B�����N
j�����R0aK740%W�M��Y�먂*����q���.�5v��m!+:�-�s�E�)�/�]j�c�1̏�W��B8�����C�j��Sb�J�@�`�GX��!�;/��]�ZVk����Rw��7V���9%��0�Ds%"�F���q��kX��+i��󾏹��]*�-,��`ۥ�֩�Qa��ո�ު��n%�v>W��Nmr�]p���b�w�}�8���aH��kL`N�Wk6�ې���)����4��w� ���(V3��L�9�)�2�ڱ|�f8�������<y��o�]:�	���6�һ jۺ��Ǽ:�+�&p�yQ�,�6�e!�ep{�;�]�.,V,.�����đ���{i��<��/K=�*.�I*v�c���n%.2J�ݣ�(k�ֻbV�˱��î�g8�T�
�,�4yp��(1Z�-d�b���{L�%g+G�N�$r��u��S�Y��s8�t۬��2�神)�RU��R����#rS��+�Jp������`ײ��coFƺ��i)avo���^�A�ԮRNn=&U������V#��so�
�X����̹e([�"o�ﺞ]GVv��C��0�8ȫh��K��X�A;�핰m]0yt��TWYX�,R��s�rS[�s���Η�-7Ct�4VcKs��q�,jD7Mu�]�v�a������)S��a���oi�}wY���U����1��o;m�K6
&��E�Պ���z���+) �R�.K�T�_wk[�v9��Q��@5Ĳ��4���;��)�j���$�4z�k�Q]ؓ8
���il��n�>�.��b������k�鎴X������V`�Y�2���(C��� ��\N�[������a�<<.�-��GQ�+͝t/��Nrm�t�w�d�J�!0���%v��(�r�ѲvZkIf��i�w׎|:'7��v�=�a��.���F���]�|�%�WWa�M�@2a�޳�����xضL��V㔦#-ʁ��"���St[z��k�Vn*=��u�u�C���*�!6�x�C��ڙ��+���eA##�i�'m����dL�e\����J��P�ThQ]s�w�Lh�ňIN]r�Ѭ�]������&aA�I,�#I��(�$у#E1�� ��2��wn#wnE�\.�"�3��IIːC ��1B�d�1��P�(Fba(�hȒ�i&$Bs��(&Gv�����F�1%@��0h�Г&��$ALMA���4wu+"�J A2wn��c�
:Q�����$�i�!ID���t�0��r��]�f�b�$9�ȁ!�˩D��c0ɔf"3T(����k$�C��Q�$a��)�f@}@}\�k��l�9�ǵ�d	VfC��;��嚖l̓��Q���D}��cЯAk=Ѓ�#���Էgm�6yIS���#��V�6-W]��m�����n1��'y7o���f*�{
�u�����u�\�W$��{�q�+�'��\��}���r�ѻe�u'���֐���{����/Ub9׫��ظdt�qj^�ϛ�����c[=t!�rܽ�-c�A�S��\�D�}X�J�ޝ���{wzGA]�RQ��yٕ=�#�I�5��1w����TƏ���_V�';Z�S07���E妭N+��U��ڮ�9;��	e���fB_%EJ�p��V�� �=�1ն��yx�mCi���m�P�0v�T���\Df'�޸ϱwP�e³�m��)���Z�q�P�T'M���}�N�ĝY��q��-S�x�t?�n��cm��)wXV�q=�P񜯥�)��6�-H�;��Kl�����gϵN��f�\�W�w���`m�b�..`n�&��R��	����џ�q-N��]7z����A�h�"*��w���F��RT:#��x`DMz��k�r��pv�����҉Vr���#��8��Q��<kj��Y� 
s�J�Ѷ�-��z0޽�G����<��뮻���d�Dl��4��j%nd'�_iU˜��;��0(��sO&�F`L<�J��6清ѳek���>ř����D,&�n�zK=-��k��k����R�U�~+W��:�:=�MŢX�Bq%�L)q�V�5*��c�4������m*��fP�x�!ݺ-�v��9[	8�4�1���&2���K�Z��<�;m��G;ɻ��wHj�#hrY¥S��.�o�fx6��:� ��z�ŏ�]��'��\���s�V�v�OS�g�S��MݯU{�7�Fm��*��3�]G�=)�qp��آ.{WA��x�+�F�D�^�)��[��C1���*�����.���r����+����ٍ��nu.ϥ��������U�@:�菉���&�X�m�荮��:��H��LۆTM��6��X�Nu|��w�p}��={�h��כ�����Y���r�evV��|rV�k���g[��5��-�P
�`�[w��Sj��MX�ߟ�{n�i>��-M%n����.ےR��{�k����<8�I���L�N�����S���>��;z��$�n�,�o<�D5���,��򙺿}_UA�w�8��p�]�{������yx�ki�|Vr��nK�U@��xm�m���Z�6�Ju{���?��5��m<��6e�IA�
m�Vn^�o���I��͘;�8��J�$�ێ����
�nBq�}:���b�����<Qq�/=/b>t��0cL�b�����&�5�nWI�X��VN��]�p�s��*9��鐈Y!w�p9��Jח��8�)�w�e'�M;�7�ä|ҩ���^N���#�|�X ]��s+�����h������靎I���W�TLDs�5���U�p���"�onL)��uv�%<��y=���j8sI��h����dke��������#^��ZȮ<���u�F�<�-��xӞ8��ˍ��[,�n5��M��U�����U6�|�++U�L���٬���X�T�9�[�K�bm�{M^^���Ƴ����<���ܨ��t��p�m]�8�%�%�b�(v��A�7�c�+�1FY2N�jݥ%
�%��e�"]�:������s�tή5h�ꆲU������qrU/m�/�-���Ж�dU�>q��Ls]<�
������^�c��;7K���~Ò�Pr���L���L���^�}�������77�f;O{k�G����D�;�Ë�����v�=�Ʋz��u|U�T9kN�{Ѫ�C��s�*VK�*&�ss�����R�w�\I�K�~6��קU� �7���=��-�u}��}}��o�O0h2i��3���f�ږ\�V�s�˨����\IJ�K䨩����oqX���{Iy$�~�J����{�A��tGh��zGH���0�YAj�HtᏧ��GeTmu����k���3�.�����!}�F�J$o>�Ŏ���=�ch*փ*�ˆ��-�a޽�OtT<g)y�������ÎmRʹСoϼ�����. �-��#�B��4�7��h6�6�j˛�粮as����tGŇ�X����֮\ᨏ6h1��5L��[�3���)vQ�oG�\��G��PƷ�]>�}�]�-�z�sz![	wZ�̌�s���kו4��E.ܩ1�Zm�g�ֳ��`�ܖJ�{����7�;�Η����"������`��� v����5��w�9MhL7�+�;"r�
|kU?^IF���Zub-u)�O&n�[�J��bbX�Aؙ6���\�D�]N��kz���s�׵U��;"����,��4Z��W�����fP��m�9x���s���uQ�L]P3K�+��:)��:�W���᭾s5�S���]9�[\S��ә��mn�I0gC4wh�p��/TFt�޻��V���k�ݯo����z7MZ����ٷj����z�M�T�_c�ظTGK�
^�����*�C�E�)�Y�=̜��;��f��ʞ����qӅD���n%�w�sÝ�:�&��d#3N!=o����O��g v��+��{�JXk#�B&Q�V�.�!���<�k�Z{p�9�7�K��ʎ���旺t��yT����mT����˰��a�uemJ7�A�K�b��X*�/�d�ʲw^i�lc��8�D����$u.�q���e�/��Y�~�[�N!ϰ�����풙�vq�[�).;B鼫�1]!r���<6��P����E�M��0�Ʃ�6O��������UVj��5����p��OmN7cl�\����2�b]�l���F+k���͗m���dҔ���]��3k�r���nP���f�b_m"�w�5S*�1��5�cm���u�V�S�ʉt�R��
�kP2��|Y'[�vDi�~��\�[1١W&�:�����2�:�Y 
c^�8���z������%�t�u|#O�>��M-�޺��������r��`�A![--�r�����w�Y	����q��Z�7���؝dɕ��m�>�0۪�q�9�L��S\�P��vF����ۚ�}P6�
�������;����2�nn�,�U4�Ú��y��q�~�L�όOz����'�'��)�6ܼ[z�~˫W���k�4���s���k�2�a�ԯ����Lj���]�X���+U�L����,�y|e��x�o��y7a��8q�K ���/u<�%���@�V�B3w#l���r�q��P�[��|(�x��á䦘�Z����Q���=�Nt�����Ka̰��ں.����{݈9�n�d�ϴ�:����3��*�_P,�b�NƽV�J�W����}�~�Y���y�v��:�\����^��>�������MnK�$����m�W���oJ^�ojs�Qݰ\>)U�zb꛾�{<�w�oq<�.UF�p����K����:�������2�����L�����'�6^�T[�A�AM�uF��a�M�R��ί�Y.x�/�[q�b�����	!|�ɴKKU�Z��p�\c����Vr��Ua�}�;B;m��U����<?�A���k$�;�]�=��8ko-�y�v��djz�\�_f�w;3�i�v_}�N���-��o���K���o5�/I�~LJsGw�Js��ʕL���u�RcHJ&��al�n�)��^�y�!x{e��%�w;�P�~Y�y���p�g �
���i�jV��r�v]P��٭P�4&u#����_���A1p�;sP�\�q����؜q��uv����u��Cl�Őb�����6�A��`��[[�@�|˫pmNl���<��뉆�K�S=\3�<O[�~,kW���n�N��W3�f��M�&�d-��7��Y�5�:�̥qTm���sw�g��S'n�щOoIuO$�P�p�2���v弱yu�v�cT+�|N&�����RV�\��X�~�x��MD,p�7��!�N�$3g�94z�m��o�Z�W�Q���y�Ɵf���s�z�-M�T�!+�ٲ���n�xu�;I��|H��3M���`�����uvŔ�X���AP�ZĶ58Ξ7Q�O5�����y0=�_MO���Ngv���5�3���;U%�t�(E�L��Yn1�N��3b�ș|���ܔ����^��O_<�ޭKGx����>����g��u<�Ʋz���&�d>�
�p�N�Q9=_D�>��ՅD�˛��v�\�z��F�8�m���u�%�S�*g_Հ)/� u_�v9}�6�p��i�\�G�Ҡ�v8�8��m��؃�`>U%GH���-E�z����lj�j�kUQJF�t�L���y�*�_]4Ǣ�р�n�.�JԨ��ԋo�a�uN��9�u{@j����i(k�
�SFr�kz�5;�Vͮ�(wa/z�Ou�������c��'r_ii�P��'>���nq�j+��'�g]���aB�7^r�s���K�J ��J��b��������2䬆�쥾�lb��=�[Z�\f�<g��;.�ܤƘ	FnVط�s`���p�'�D���Lo8�Z축�w�S�ٲ�
d��ՠu�us���fw{ڔ����H��S�V���wmʛ�x���bw���y@/<+Mo��M��'�gqIs�ք�7�vr:���v������sZk�z8+��{�������b�uⴕJ��l��x�J�q��R����f�\d5L���m��̩X�%�r������k#v�zPB���\�^(9���C�_k��WP�U/2�pԹ��L�f2qf��e%���YW�����=�;��usI���Ûβy���&��������.b��➢���t��|�;�/�>��_c���#��(ˡfmy���]o�IVĆ�:��d��ɇs����9ڗ��ta�)�,k�����*o]��Œ�m8�w�Hi|���۶<��땩�sS��%����**�(��rz�]Aʒu�F�9��mq�T��᳁�Oq��u�����Zc�f���"���}GֆNt�p�;qGb��넥��o;���85�����ۅ��f��{���[�z��Wҡ�F8�¢w�3�1�U�:��J�֒;wq��R�p֪�ƶz�����uT��*9V���ޡ�z����u��C�p�/����Z{q
s�od��_���zv}fE^}w��`����n��i��T�N��p�c���{jq��+bpU�å\ŏoA4�^I�'�xWeI\�ZɨR�\sֻ>��8��'O���<�4�����>^�¾�����6��R+}�	���8T�5SB�ۂ2-������p�OW|Ԉ�J* j�6�f�\�P�[�F<K��Ǩ��>�l�I~���_W�q#�>Lw��{��z����*�`��{�rv�kDGeKi�w��Ȕ�S~O�"s�ћ��^�^����=[ۗ�["ٞ�0�E�D��q��y�/b|��w��0_8��r@zoZ�w^���1�xM����B���@�,��.`F��SY���U7iL6�J�8�Duܼ"dNL�®=q�:+���w�'ז��t6K��'�L��d&�6y�o���{F+{��(�)m��c����{�ʚ���7u��󚴳%s����e���)2���-��s^�0�����$Ý��2��K��.R	�]r��h�����J���7f��v,c�l�A��J[WLi���'�x�^U�"��r޷�;�%L�7P�HB��=���l
���W�\�Je�M���qO&�:Щ���7��#fH>l&��dV۽��Za���m����Ç�Q4��b�K�n�c��f�aBu�V��x���s!g\֏KC�(�.e�Q�:*��V�$O{,��:�d��h�}�WY�����3N��<����}u74F���kS�V����8
��7�$��B��M�n��>nƞ�qfa�q��Xz����>ܴv.�f�B�p
Wm�0&v���7!��a�[�t���qw7���7N��
�_(�PL-=�q�f�A顛���.:
�sŹ�nj�$AK�7��/�u�y˕3}VM��Q��rb�����U׮��K�[ظ:�P찞k��R�hw$�k���]�Kk�h��H�l�&Ȣ:��h����<3���Z�7�<�7���\@��:����g�c�1W�$�V8nty����]����r�7��zm��5i2]mE}�K�O!������M̮rK��Z/:^�P[W���Gm��w��Æ��(��-;R�1��ԃC�˳E���T�ʛZ�CR�ղ�ⳡ%��=�B9��W�ܲ�뭚�Z�'�]8�Ŏ����KrÙ֙S���
�Z�r�
�i�І��w��R��on����N5��]վ��Uq=��8�ri�Pa� i�zN�]wH�s�e��쇃�4���te����pf����
:����ɔ�P.-���On��t����*�ŏ���M���O ��V�֧S(�u�O�58{46��471䠒%�P�� ��k�:�	cal��ϳ6�w΀��˶kKpU-��F:s5���m�̶)'���#����8��l�%!l����Y���1pC�]$�d)��݆�Yn���V����!y-�u�sG-���Zs�$BwK÷�����=���gD^ƳugK�0s�s�샓���Y��ܣ�Ve,蒼�����yji�=p�x9��xV�`\%6͚�0"��r��<J�앙i*�d�{�=�h�0�ֺ.�/���oS�r�5�����t�1Ӻ@u������B�R�����K�]����ڛ�%��X�U��W���D+z-���JJ[cx��}"�t�Wp;���}�J���f�9�W�fv
X�aڵqd�E��I3~C� ��>b��&(�&�C�t�	�)"B�0h�c#4��3wsM�4�B�ʹ��c3,�5�v)79�,E	�����Q )L�$1;����ѳ1!@L��s��2$�-&�(BHƻ���$l(�����	!2��E�Buܝ�Ҡ��cN��d�f�f�ZQ"	4"�1b
I�ɚ6.�ɤ�1g��i�u�@�9�+���lH�w�Dn�s��L���J@&��:�(%`�Hb�����B�rC���i�
�;r��)L�PH��k�"%��3)	������:b�]��u#)�X���l� ��
�T��
��E�j`�88;*-�l��U���M��Ws��P�����>YEL�5}��7��]S\�I��adLk�������ѵ"z�hQS�Od���M.�N�MbɎڷ}Φ�8sPہ��9�Y��@n�즶�Z��ɽ���^��>�}y��Ȩ��:��cO�f�k��x�yJv�nw�srwcz�z���IW�fq -�/�3�6��V�Nb��_L������d�u��m�GN�_J�<7�OVOj�������ўz�E��ALa2Y���2፝�G18n�n5c��8sz\��lՌ�G�#������D����L���ʉ���
[}�K���tc[=uc�*�Q�Վ�h�a��A(ʤq��v��=�\O��76�}q��7�	��q\|-�������3w�
�@�r^�L�;W)\in��p�_��ki�|Vr�[!���p%��ky�Nq&�� ك�~�}%*�=��ٓ��8k��ltE94���=�r�{�D9�z�{yG�*��,`��j�*��7�����]�F�c�2���`o���SIHu'\�`��d��{�2���O	:�+�!iǤ8�_s��b,<A�}D֜�9�෮�jVP��,\J��y\:b��"I	8�9��B�ʜ6Ӯ��m���26Q0Dr���䄻�+y �E7�	��P�kZq�K��NK�_r�1��TO��І�vLd���i�2�֙�e4���Z�0Sl�DK�h��]�69��=[��=sN�rn���9�/���\�7��f�V�Bt�磈]JNk�|/�G5v�1�S�W.u��bs��T%�5���tk�J�(�]�N��n=��Q�����k�0V�\����>�x�S=9��kq�{ja�.p�%<�w^��1��	�g����/'O�����=����79��&��lK�C:6_�֝����o���w����N�|z\_M��V� 
*gE�I�U��8S+.98�q�Yۈn�9���|����{}���b�\��A��5Ӽ�Y$�%�޸�Qp�뿓�H�~i{6���a���} �Vv�O=8�[%ߨ�ʐ�yZ�4�7RQ��:��(���R��o��wt�v�Ss:�z"t�v]�Q�9�mA����<"�˪<���ǩ\h7W����]�	@�1�V5YW�Nۍ�,���;�],T쥐i∳l�3j��9��'��^D~=[�����s����?���"]эd��f#��l�j��QB�u�˞.o�/�
������}r��vG
�k�gw������Fml�t�\��ʁ���5+��=ΰ����n ��{�d�\�K���j�������QgK�fN����D�H��Ե{�X��8���;e�um������m|��C�n�eR�������T��l�j�n�8	T��E7��
]��,k�5�m|�t�:-}�D�p�O���e�F����Θ[��iXw�q=�O��]3P�J"�yg��g'��☋0;��.��Ъ94��@v�Co ap���s��U�]�s;5����l=sr�'�Ғ\�7��ڌ����/h�����U�Y<=t����W���s��|f�j{Kʭ�d��K���5�:�>u�a
�VAd���sDLZ1V����FZ�����1
G�)dSr��U�eK�>�MF��euu�\�{ �=�<1m�c�d$��C��㏇=b�u7���6��}N�L�I1�s��)|�!Ld�Y��b���F�k*�w҆�Km��k�
n��S+E>������ʈ��zu���C�3�;�]#U��w.�d}Mp�⃛�S�Q�H���+k5\��æ�M�O�x2�t�YV����k�w��s��l'y7>3�"���ъuoF'�K/|���U�9w�mN|�����T�����fܹ��YE�n�{�a�=��;*�m���T]/\(�K��Ę�t���Lf�������|����W�m�����z�%C�q|�R��jj%_��x��t����r��f���������+�j��/�%G)�1�b�,��܇�#�Q3m���M�����)Ψ[�*�����^���q�0�]R8�m��8��p��c������eR� 	[U4�-Z�i�ըp3D���Os�V�j���Z�qy��Rt�[�/7]�z�P⧩�Tz�0�(�k��w-��V�`�K����m��p��s�:Ə
Y^��*�����\|�ҥ��~z�lf���Yl��͖��~~����ݸ�=�|����ܸm��b|����]I�I��Q�'��{���n�uw�nR���q�Ը��'|��7���5d����K�·ۉ�wB���O��5����u�x��|�i	D�Z����Ъ94�v���bT��W��N�80W7�Nm�|�J����	��J�ˈ	��#;"�>n�č�[.|�6ÿ�ȘN��6清Ѳ���N��r�v[\��A+�qK��Y�c��}'�sޭw�Y�b㝹�|���&�!\�C̆�
o)��˔�j1d��V����,p�9�������v�ceJ���k���c�\��􊏧��t5J'����p�Ú���e݋߱�E����q�����8[���ԝ�_�|z\S�TY�2�:|3lE�y�j�����3o\6tc�Ȼ���e�_����f/���N�Xz�j�c��G�k�����q72�?��<��Vt��g7���63UQ� ��ہLl\납n�6&�v��ܒ��t1ި8��^�=g�w���S�������E��z�z��
��h]��I��ۣ����L�tLw�Q@m�OT	]f�|�f'%�Й4nۭ���Dr���X�KǴ�`�/���t˛�}�M>mtV�/�%���Ȉ)tc�gF���dD�ݸoUF5�ך$�oon�>S�w�9q��A�I�T.��ՅE��&�\K綧:�Y.-e�H8�w�UU�-w1G8f�`u���\��4�wἿ����ʚ9x`x�bN��$�s4���<�n�N��D���=�U=��j��P�56�k��,޳.�df4��}���+W܆�@K�}'��u���]`r9�G��1oO�^�ʕx��p�Q�p��8)`��9���赵�;��p��d�����-�a޵�`��g*]3EHU�}��it3�}�ݎ_=��RJe�;�.��+ysW�o�b�L\s�.˗��<$�~�yvǂrY�YM�&�by<�xG'5�xzP��=Qջ��J�%y�����:U5���Gsћ�j{Db����IT��g���;��wFN���64�n����
��A��W�6 ��l�1ڎ�c�9��]3z�n�춸Vj��E��r��q�$Z.�f���	��ܚ
/��;x�i�u!�;`XJs�cb���5��Ǡ�<(���K��<�3��R�� �:�^�{�I���!aL���hֺ����]�+���v+���OcΆ4���5H�'x�;Cr��C�b[
]�Gn��=H�z,o�%���,�A:��g?M��60ո�����>�6��-�ީ��t�������|U������|��W��m��P��]�X���j^�N}"���^�o�A&�l�;c�-V䞣:�p3�M�TD�>�pc�p���i�{��{ı�j6��_T*�\�2seL����uT��P��_`Q\��p��FT��K���T�#=o���5��\*�9P=#�jWL�X|�(�U
^=��]��
��Ϯ%���9_�l�\O�~|�JU_.t��-�
Z�UVj��4�j��c����9��m�_/�I�0;�[��/[6f���{�q99���|��冾)v_,k�\f��ʉt��1��okԼ����ͽ��/;��l஦g'�$ƱwE���ѧ;�׷pXI�Ɠ.��v��d<TFF�=��v|�e�/^�|�Rkw���Nݧ˞������ܷ��xBt�8?y㙃�lhl�&����X@��k�F�n��X3+�}5��}2�P�.zM���]�Ұ�^�'�*!�9Q.��>gek�Y�/��;��
�K��
f�fJƬ.��4*�ҿ�|�hwv��h����u�gWy�\���y\O�K��"s��M�uJn'�O/�;�rw�9Yx���5��WádZp�r�4��=)ޞj�����ʓYG�Ԋ�n��$��"n�w:�X���c�kT8j�Q/�ۨ��ܞ�S.軽t�+�r���YL��_�6�_r��[�r�A͆�+�p�>~�)���n�E�g�Sޮ��{�ԑ�qN�Q>u�}���վ���w�7���"^_p^�\�A3�39Ҿ��^�Pb&ޫ��X.9>w�_u��	�t��C/���~L�o��j������V����<��8er�z���Y{z��fLJ���=mm6����&�9�/s�Uaf����r犇��8��@���:0'��p���<�n���/H��ɼ�{\4;ηFHo��C)�w����a��=N���R�ƚ�I���5{웲3>W�B�<��n㙦��n+t�)����Z�;iQ���e�GI|�[�O'DM*������ jۮ���=�9�J:�[:�ʆ�����T�ܧ��.ƶz���
��$���}��K�5�u����#%�#�Q��o�Nm6�姶�:��J����;�E������_Kq��.$ۨ�i_��Mbo.5�Yx�m6�����p��r�u'���}�t����3D�mTI�v�d����~���ϼ�J�5���]u�S�\��U����I�0��o326ۚ)w\@V�UR��x�Gj�����f�'�*U3P��K�i�%V���{4'�O��'�=��T�.����'�W�d�wӔ�J���.��i	���+s g�d�6淣�4&\4¨�\�7��L>!9c!M���T�����{qr����.r^����vf�퓜�$��n5�Y�~�nl��zE��Q[�N�N����_�^U.Q�r���59m��f�(I���%�ѕk�`ufI���V�
+R�Z%F���{w{�qgH4T�'0秃t���@�vfiO�Զ�GA��Nk\I-<��*�F�dY�Sy̬��vj�ͺo!j�� �7x��D��u����j�%��;Уvvּ�B�L�t���R��vT
��VaX��VU�ޗ��Þx鈪�Pw6˺1ۓ���N��y�$���ݨ�^OMD#�M��<�]u1���*&ŷk@�t���=�Ax�#LNz-�Ts�o��`8s�2�T�>��h�'M�]�����Q1O��F��f҇0�ʍ��[�rk�Sy�����NmO�N�&��	��R���髰�,���<�ɫ:ŵ5�f}��3���3W�<����|N�/1y
�3oՃ��dnӡ��>K�-���\���(���t��sM��:��*�ǎ��x�y8/g�5��׊}��׋�d�_�#FU1$�v�|ǗA���޼�q-���d֢���^�u[�3+|seK�.��D�Lo�Z�j8�'��c L�:�F{�)�ϻ�Q+�ݦ�b����7 oU�Ć�����>�23�޻��q�/�����L�Kf��=��4%Ϧ2[�Z9�����R�p�r�.O��7�E�vԏK��z9�'����������!C�����Z�;4[�I��!Z��k�m�x6�տ�	gZ�ד�,�Y<Q�Nfim1�%�{rfNm�9�їʞ]K�1������w)ܟi�-�7R��ʔ1���0Y@��^e���#L�t	���1f'�ӆh�;�cH��]�+�1��6��f�)�:�c7�ܬU�ܳ����[�B�ٙ�&jc�rˁY��P�.>�կ+(��lW{�[�	7�q�����ڕ�a�ROxQ3g7�*�_�T���_gaZ��zqmcءd!�UH)��uƮ���t���ڇW]A-2ve��*�V��f�e䝣�쇎,�ܺ����������3s\��Ӵ����ڏ�S�K��:7�u��v�ǋ�-}�Y�e?�J
���#$�PC{�.������$��M��|y�j��̊������k9ײ(�=z�ջ�\b�,#GlGo*�A�whc�๷W8=�[Z��؛�/���X�;1��;v�6�Iݻ�6=�|��z�����F��-O�aJ�b̫x�5� �JoQ�O�xu!L�t*�Y�k�Md�I�`��DQBrp�ši -�s8�
9ܻ�� X�͢i���mB	�-�����]w������7u�s"6WF͹;�>TH��ʊ0e��-��T�n��&<�e��6#�J���u�ҔWGZ�.l�l$c��@´���6x+]Y������조��e(�"e�WPK*MC������wi�fH4��)M�3�NV�n���^���~u˛v"T���3ci��+�\���Ȳ̭|Ng5������7y��.Z��%�w2���岦|f�;h���L�$kPۨ�7x�FMh2��\�'O{�Sj���S\&%�s�e��'9Mŏ��I�]������J7G�0u8r+g���ܲ^�&��c�3Aブ۷g.���Ȁ$�Z���5+w2�RX;zJj���gn��W�>��i'w�Q�0��WY�*a��&�"����c.�=����'�ƉµM������y���&Ȅ�e���F8�J���5k�kU�(
���V^ͬ=a�}(]]��&1>�)��$TO;F&hE��e��rU�8�ha����@w\cl�R�Z*�J�{N�l+o����\�r(�#4ŚM�#V5b���3m_�"�M+U����2�Fx䉱�
���O��Z.�,���r�9��V*�{�̳\2(h��㖏;3s��@�t�:����fd�d�@8�m�?�h?w�-�^R{�|�kL�����Bq3*V�Af(f;��c`���y�n�S,�mZ��R�����!L�MEPN���Lж�5�e�/�ިz/��w��Bt�(8�Z�cW��������Z.(ou������Iz%8��Z�"�@�r��]$��z1�	ިDR�4+���ep�:�va];D-	�V#ح*k:Y��:o%��
|�zS+�8�NM,��N�R
�#���� 
l�^���H�N�˻��FK���D�f��`b8a!<of�: L��^ A��\�:L%����b���he�s����2���H̑#��7��7u���w��C;�Ww$���B2X�rSDɆw\���:9r2G��c<�L���.���r��iBS��;��r��c�����#���+�����w;��$Ar�]8��;y�(��x�n��یGwwG2Y��b]�n��
.�r3��\�!�k�:3x���'ts2��&�Ν�<��!$���v�]wuΓ�"��<w\㱹����s0��Mݹs�͸�O�P$�
�F:�&1��2�h��{@�4u�@���K{^𽾗^�x�+~7�=�V ���f�j� �iM�pd�ٛ��.t���r���*6�`~�u�c���˛�[j':�w�"�%�mT��>h=��4}��f�����{�B��>gpQ��v��8qoh��3�'����W����3wS:�O��\�$�EÙ"���]���\l��ʈc��wB�M׉����M�O�I���Q�p�b�q v�P/ib/L����P��]�ϗ�;�w��)|�1�Ϗ�D��$�+c�!���n�/�342���9��[�6���w^��qE��5�e��m�Y���0�{�U������q�"��h\�S�Aҏ���6:},z{��U����b��ۤ�̒�f������F�]f=��k>�i19�~���S9��77S?����s�e�j�{���lמ
�R|�d�}r����z8l��@����s���㬳o�K�W:�cI�!M��ei�-x�{(N���Mi�@���`N�V�6^���/zq��3�/f�F��j{=�����ɤ�6��3��wh�?ra�z�d�j����.��N��5ؖA�*R�+�ѫ��XW�P��E���ÛY�b�Mruל����D>E��Y�`����0X�軝��0gq���v�η�;%?�)d��f��a܉�}A���St6�p��puR���T
� ޗ��Մܕ�W�3,_77a)^^�{73M�T[іӦ�O]!?>�
�$�C�ʨwF|��E�L�l�	�[ֺ����K�����yH�ߢ�C{>�>Lg��֎��I���A'TL�ꎨ�3�0%��N�!�1]��/(��\UE�S���g��>�#�W�\>�Mo��t��n�<��ޏBqWϲw�:k���]�Jn}�h���޷]��1ȳ��Q7_'U�;��K&����G�z�~Ż7*n �0�|\��^����X������2���]��v߼�@�3=��~�{��J��mJ�5�@z���N򐾒����ioYt'�ldA���Ȭ��&�+g�qWx�v��-ز\s�`Tr�z}�&���$��$a�=��H�W1��E��H��^�>�u۰Nq�|�m��� ��+�L���0��E�K��R_�Q� 5o����;��dm%p�J"��wQލ�G��%�h~���Ƈ�Q�������V*�.����������O$�+�«���k�Ѻ��c�h����!u�4+�8����E�?�`�o>�0�_�NC!��u4�R�1��ٵ܊��]-�Tۼ�x�<�sZ{�t��ts�� 6��ĩr}��$����X��j�s��0��}ۈZ���=[�8�I��/��R�3O�����ff����.hi�`T
,����[����Ϳ��xu!�R�踧:N�l�꽻��G*�dgcC\��V[Q6U�2fk�=i]��ӛ�����6\7$��3�Mه>��N��L1Y�ˬ9�9O����~3�6���6���]d���E�]!~���{��{|uT9ɝ;_�W�� L-j��8�5�u�mŕ�����X3�n9�Ѿו����ީ�</"g�(�(��4��#��!�1q��vߣ����sR�yRf]L6v_�7}�����u�P�RIU2¨<y�r`X�yFs��{��*��f=Y!���,��O�btx�}�[;�O�{�^����+���H+>n�~90��j��<¿0= �
Z�IN�O��(r�tǆ�8k���r���x:|�;��D�t槮����rM�>�>�$�<��H�.[7�L���;��\�ƻ��;�hY�C]B8�,a�Gg�O���j7�-K5�y��%��J����z�j��t�GED�;�=v,*M�n{eF��q�`�k��T���]�7�S�`�<H�%��_��a�Sp��)���4��:�-T��ҪM�@Gge�H�}��쮗��)EF�BP�J�ֹk]�q�mm2���¡�	���q�B�Ԯj��l��+�H�6\I�DƲ���+뗻�����̤V��@˥i�(��Κ;�;Dutۧ��#�9 o3�rXdtn�-�����v���V��k]UIaI-OH~�*�wB[�r����m׮M���io
�\&��n�����������S$_/&�}�$5Э�%��1s{ܹ��{��+�v=s�(R�vUE˲�/��ڒ1���\����(��!9>��&]��%�2�5Eх��b�����5�,m.����]R��j[,b���۝��o�k��>���d��<�%\��\@���M]�G���.]z�{�Ԟb�.z'u�ӻ����r��)�5CO��(eF�_���$�>�鯍ڎ�^OL��p��_����_��	>��
�h8�S3�Nl��.1����Ts�oϖ�	tn͎�L�v�lo��M©��x��|\�<\2�e�y�k {�Mc>�~Q"����e�>�L0���
��Qo����k�M�_�r��d%=��(�P3�^��ܝs;B~�����q���KL�o�z�n2�y,��D�~��c�C�_�-�_'#���(=�=P�oL/G4��j�g����@��uum��Fu���!�8�#�V�t}�,���@�Ɖ3��	(�fU�|(�;x��Y�Z
:� 8/p-����+U.}`�����kЧZخ��]�����954jtҨV�IGT�i[f��uc���K^޺��V��	�~Zi=ʦ}Q%���b�e#2|疇����n%�}Aτ�p��ړ�#|�u�����F��>�Q%��c�)��Q�������IP���p��Q�;�]�m�Ly=��#:m�@v�z�]Cu^�Ӓ]ÐsQ'����l���w�}SU�=�U~�W>쁺��N�p���vO��<���y�������|��]}���^���b�}'��zQ�^���s�@xso����'�3��uu	�3"�y#�F�'�z�.�2���^�qy��`�9B�t�7��u�v��2����q��#ƣ`b�I�����ʱ��]�Օ^p�R���!��M��W���j�X�.VC�j�
���exO6�L��C���1��_?���ДF���Zd���R�خϾ�y�Uj:���c�p��ۥu��&X��� �^��P�C�u|�zfv�����uBj��=e��.:A��g�7�L9��c�Q{�����U�����s��!��ze[�A�<X�6:z�z��� ��"'Fj�¼N�˜h�/:s����t4oN���S�1��j�Nm����t� 4Ѳ�C�.�8��Q��\a���o�S�;��5���Q��z�����2�_��E�!rL]�����V�[�zb�S08]�⛯��{�t��yp��6j�iQWYQލR���o8ZϢ�LNz?~��M2���$��-�ʊ�_a�]��
0�~��:'�������d0�w��'XϾ�)���Yf*��rc{c��y��gw�̵߬��s��x�w�ޞfp�S�<�#i�0��Z�/d�u^~��v3�U�I�R��d��
���F��H��p�� �<4g��z�� 5qi6���	�:�b�Ү�u/7Һ��ޯZ^R���,��Q���j ʨwF|��3�{&\x9�^���䨞C͖�{��E���}�|��G+���=QӠ��&p	Ts�����N�8�cɛ�������c�T�~�qd׍\kw��2�>di��j;�2�O��~�{}꺇^Vڵo9�*����?LmL��ϭ��7-�1=��v;�4���\NϪ��<�8E[q7����=wu<���}<}� k�2H/�
=+�j�n�1量�/�Le�Y��߽��=5Q����kJ�V8��u�X�K5���	+�"������a����1p���k�~�[��٨X{��s����
�x��H�˖u��;/h\�j�so 5����]�sh^�N�o�&���E�d��V <n�B�T�7:�6[�J�*���z��fq�Ӌ��X����WY��|�I�4wr�{��v�H�/k^>��&�G��Κ&�5O	��s��kj����
��MMDi�{M0��ѨG�ڨ����/Ҧn����SY}�\��\k��֣Qͭ�,�9X�`�r^jb�d���94d�S��Y�H������'�R:7���un�R;g�(�m�:dz�!7X=.s�s�n2���r��S�AN�?ENi�qOi
���ˇ�%�a��Z=��jG���Br��QM��giu˸�@��O��J���V_�ck=l���_U�xp�jy��r1�|�S+=�v�x�j�����w�{Vl��/����ݲI��3P��r}ǩ΃�L5��c!U;�L}mK=�n_�`�Z�MW�oKfF2���5o�x���k�*����(���G�/N�-*5����1k�3^�:uX>d?�5�G�9&1��v�n�Z6�-C���={	� uW:_���öo�#�oV�u���P���Y���¨Ҩ
���^2�a���~���>�<�"��$�_L��'^1�<X�ގ��a�/���3혨]#�j̳���P���h�#��v|�=�֣o�i�f�:ɘ����c��[���j�����OIC���]�����D����"�
��f�ᕕ��h�&�A^ٱ���ّi�3��*��Eh&�s��Sb|n�Q(��Ls
�tlt�:2o���D�eV����y��Y.�}�N2&E�ؾ���E� , qp��o@�������A����.¾S�EBS���҇*���,z1�\/����}G���������Ǣ��N�ax{j|mI�� $H��l�T����!�r�V=�>;0�xd���Je��W�GU�m�5�l�u:�ᖥ��"uc�Oź�J���g�qO@�7�j���g��� \�s����,g/����;jE���p�改������g�ܠ!��ZC&3��Ȼ�E���X�i�\j.aC�������~�����2��RxV�=�PHo^Ept�1s���␭N�I�83�f��w	��n^�Ͼs>d�@�`s���/&��f;�V��Os�mVi�Y��{�\��)��P��l������ƤuwmR1Q�Ί5�\~��{�i�o����{��XD˞��c��'��kk��4�Xڅ�xĽwB�{���@���@c}�ao������+M�P+�Y���s����5vdu�y�X_U׫�C�s��6V;!z��������v�r��7(ek��=�O� ��7j:�y=4�Y,�,~��rᅝ�Y���sg@�ek����uW�W����	b�L4WSQ�Nɸ�妹ЭG�Cʲ
Uef�i�%ì��*���2���R԰[���[����D�c�gm�d!w(3�Y��KO	�g�Zfg;��Aټ�Y�V�.�B���0�����������Iu��,c=�bs�o=b���h߾}�b���Qvǹ�/� �y�����iy��'}g`m�P�9J�@�&��u1w��̯t�S�z�ٺ�ݵ�bw�*+���<���:�:B�F��g,�5|/���Z�ru���~���u�`Z�30�w�8��;V��=>��k��u�A��x�\Tϑ�rW�C�C�}�0��4��jq�NNBsT�#KC|�r���}t���t���0��:�R��7U>	�<�<��^�=)O�w:�4�Ƿ�6�2Q���s������-K6�$�c�\*�Q�̒���7�F�J&-8�}�u*8�\D��ﻤ>��E�aw�#��0�2}'�:@Ҿ��L�ю�so��2��(�N{(�F|w��yB=�0��3�n9ȳ��ԋ�MW�搖j:�ަל�BsW瓋2���~z�_|/K��Ky`�O:�1�/�O��7d��O�:�d<�`������A�E�>�I�$�W�P�ӌ߁c}��v�&42��e�\Oi���%�׷���\���E�+\׹}�9P*I�d~���5�n�9s�5�������fSU�AΊ{�..�:KӇ)dV��ag��u��w
�ø&:]����A�������	qP&;��И�*��5����}���L��Sm�^�C5~�W�q��W3��Dz_�1K��s���>������b�������gR�c=b�����l���u�8��8J��4t^�9Jdߍ��ڹ���n��gj��Nr�e;Ѫti����j�����\遅��2��躀�����;������.��y�[����{r�c:6��*���oʔu��V�v4G�O	�n��օ��|�t��ceY;U����IŚ��S��?VV���ZN��K��뇊�;1��p��[I��}��W���i��U�w����.׼��o�$&OO���_)�6+����E� ��j[ށ�:�}�9L�/�cA�NxQ��|��e�,������6��#�x����{ �,lVMi�� yl�6�@�U��`K�����agr
w.5���sct����=�G,�)Y�xh�T:���_B���CO+���(OE�~��{N(��oyw9Wɇ�N�1���A��PJ�Q�-T�ȣ>G�-Obg �O��a/j�U�G��PW�U
���ݵ��|��Dr����d�OWJ�Q3�(�=���z�,��ia��
�u�&��yD�8)P�ws�8�q+_#+7C-���o�z�wT���wx�7��]���T��R�f'xbX���}%���4k�c�)ͨ)V�H�:�c�z��&��(�PN��f�2C$hM�!6�<�n΀����P��HFKk��[y4�;���4���u��1)K��2�����V��:���Vu�������l��E��g����;x չ7��L#���:�ޜ�5Q�Յ�%�8ʩ�c��.��L���Z��,Z�{��IY ��r��tY�'RZud	��f��%���xHM��4"��
K���p&h���>�nP9L����0�M��!�v�GJl���_0�H`	���A)� �e�ۙO�U�b�hd&��l�1�.�G�M���HK��33��lQ֑jF��&�%ҒP�%�w���[B��iVq���{#Zo�I|�U�%�(̬����c��
#���]��]��Ջv���K�vq��T��z���+��(c먚�"d�<�K����2F0:��n��<�W��Рȭ�LrY�M�bC������|�lD��b����G�MަED�<�ÝXw1:���5�����F�l��l�Uہ6����`����;�ok4It�n�9]�Y,v���=M��f��;��Y�
4�Y�|�/T���y87y�3s$9vQ�_\�V����/�.�g>YJE�>�=�D�5`!ܻYS-3�3�k���g0vY���+�[ �>�!А�T;���7����j���I����(i��5���|��gm�ˆ��*��SV�s�	��L�Hv�ߖ�L� ս=�L.��zMh���9	Q�E���]t�	K2���R9}�mv�P�z jX��6򲬺�BxV��k�t��'j	����t��%ұ�`�¥��2����������@c*(��1V����<g���ږ
|#�BTj����D��n�5ܕ9��e��ۥ]ʴ5*��{Y(�C����~iCg�Ч.�a(��U��|r�׽&J�4���)��J�@R̺���PZ�xwM�K�k���Z��ڠ�]ڎ^H+��pQ3��-ΝI�}[3�|̾SC�$l���b�wN�n��3LǸ���kR��s�Sɉ[��\��1b������Hȩ��:;�\�|۝t�v��m�!8����|��S�}�8���dᄙX�F�t��/�&�r���T���u�4v�c5�|��NڵA�'���ݞT{�:�,h�zu�«Ԫ�
h��:t$ږ��{U�
Z;����+5|O��#w8=jÖY/@}����4SA=�.�ЦkQ�e^�]�\3Q���^���#`�V�T��R�����#��G՚̓Y��v��V�}ݔ�R s���7��0�$n��wH�(�x�b���]q$��w.�����o3s��L�\ܤ�:�s4wn;��.Η.w�׋��"����np�;\��˛�y���#s.]��.㺻���q�s)wt˷t�]��)�r�u�]��wur܍�wA\.�\�ۚ�����%�ˑ���t�sn;��]��u���Ӝ��������Ȝ�;8])��wn�˝1�As.Y;�]ۡӣ�p�rB�wuݢ����].C"�;�;�]ݻ�%��N'.��\���wL���s���G\���wˎ� ��%��9n�A;�L�bE���]�F�q�;�\�
&]۶;����렋�qt�7M̅��I����
&�#�D�� H?C��<�������t���V�:��f2dV��u��wPkY������{ݜ٭���u�kS�5��4���b��sySU�ި��/�ROd��t�ǓLַ^¾�H�|}�q�w��ϙqf��䗅��<>ӗ�u�6T06ٛE���b��~��n�M�-�2�[Gc�#O_���wꝝ�K�瘗�e�d'8f�x�8�Q�P@N��?��J��X��o���O�팃����s���=B�;Ft.�g��g��£����Mx�Њ��	��R*$�>pa��[�C�b��� �f$��8�8��i=&�j����
�$��i�{M0��h��6����ׅLg�ܭ��҃���l����h�6��e0�|9X�S�i����/f�94:�ʌ(S����+^-�ҷ	�h����~�������J-�����cC�(����K�ꑢ���4����qj���d�\���.�¨��*"��Q��uZcݎF�w=r�n�ڟ#W>�k{��mu��GCdqf7�a�)vlO'��\�k꺯��c���q����і�y8��Ԍc�+7�M�߮����I7tf�vc�y<4�l�\ ^x�o����ǔ�*^6�;3��J�������?���vd�^�e���c�[i���W�]�ww��k-�Iy>��c����TG��zy��y a��:�Pr��<���WKܠ���a�ؔ4詑���ʕ�t��2a�u�q�Z]S0�n�I�R*�r�h��`���F9A����b����6���A�~"�c���#�+��Jp9u1��=���ӵQ� {���"�j�#ܓ�[����^V���,G}+Ic��9ꅲmr��7��.���J6�9��9q��*��N{�\C���dS��w��|먡�����N��[�㗮��+�s�����u3�1(���2�՞P=���3�r{Tu��W������_�\�f=���/�^.*��� �<+�:�W�KޟGzP�|��p�E�8�"�s�����x3B]|�lt��|;jY�Q%ўD���l�T���ǚ([���W��������Q���O��г��D��MG8jY�"���d	�܀u��:˅F~ÃϦ2^v�^��	����uK�{�`�]����z�~��K )d�3��CWd(���c�kF������S��i?��q[x:�7�w|\�f�.Ճ_Cn�
iy�Q�)<+�R{f�����b3�x��]n�����x*S�ؿ̭�
;{SGb9��Yd�%�Õ��9�d��gB�1��^�7��&�u*����Z��Q����̧\��w4�"�t|���Ef�.�Lcz�v]R>��J�,ti#ݶ�s�jk�<�L���1���v��%8�Y�;F�2��:���r6�������Rm�P}�q�p:���)n���l�2�����c��G���W�i�/�oz�;m]ыM�������|����q�b5z;kq}F�L8|�w��[ShNx���k�٭,f��b^����$�;�1Q���9t-�-K���W��
�}�-@Q��d��0��N�W�t�Qz}��ƍ����xr�(q}{���`)�}�vv4^r�M�7(ek��y�$���v��!y=*]Զꦥ]���ڞ�%���+F��x���Ƴ�i19�y���ѷ�`ټ��㝖�	�)��z+�1;��^x)��Vj�'ME�v��?I�d���:��y�l���֧�{�����{zup9�� ������Be��:6��)��Q��(��^0���:�\fx�Gm3�\���|��ץ�p�e.9g	J��@�/��7�2�f����� ��i�)ę���4w�=���>T���	�z��Ϯ�>���u��|eSS)���O>ytx���|c��� ��t3�c�}��<�{}@>���iR��y����Q%���'ʡ�Q��˨ج��Y��� r��Kmȷ�0�k[�	L����l;�z�@$*z�.��W���[H�f��%�l�1B����i_�!�쬕d�vA}�{�L2��͢��o���3� \�Y�4�7�'n+V���86��0+o�v�kB�Y��)�f��܌���AQ;���k��s��������]�{NIv� ��I�.���aC}��v���h�K�,�Q�_��ۊ�n�!��ZS�=��H�&���4�����k:���n�ʆ�}2��p��+>񨅽\}/��c�_��.n�m��i���G��p������V�̝>��!� v��Nq��,o����Ɔ[�,��=�f��������w7:=�Kbc %j���k�mL�Չ�ϫ�n�[5��-�!��+ֽ7w��Jv�\�8����u��-�uG��	@�k�4kL����P���v|�3k�}4,5�S��	y}�Pp�y�뇢7�R5m �}Θ_��(z���	�əW �|l��pw���0I:s%��J�M��/�=e_��ٮ�O��h�G�.����h\�=��ܯp@�4C�Z)+���(^���82�^L]|��6jβ�����}�;1��Y���bs߿^	Rܑ��坻��������i��~��շT��գ��:6�������B��Gj[ށ�ճ$}��gc�.D�����]W�!yϮ�J�x"��P��=���ڂ�uw];e�aB:�ƿf)�Y7��m,����"t������f���/h.m��f����	�v��ȝ9Ӯ��H
Ǌ�0i���$� [�3�4P�u��`�p��z�
�����t��#Y�|�,ź�Xq�x����{*�,]d֛� y\m0%k�+��Tn��]�/(1sx�8ig9[^������ۤr"����xA��ii�] v��\��"`/&�*��{x��D�p�ǳV��XyНhc�A�mP�<I��AS�^o_�oLE����]R����ٽ�a^�U��Ro�n���|�&3��Gh������Iܭ��~��Y8���㶟 �^(�B��1_)լ��+����w�{�8��(�e��5Ǆ�Kۋ��p�r&��p@��3�H��h�Ē���ۭ[�0rv��#�̃q�P\��	N�f�+ӳމ�Ez�t+�����0d
=+�kc�o���O��+&��B�Ɛ�w5V�c�	��Q6j�Q5�O�"T$zd_�^�<.��3��蝯2kv����,�7�S���_�9��jj��k�Ы�I55d��_0��Mz�T2�)k��c6.��)8�Q�U����5ͭ�Lo�9X
>�T�����}�%��q,47�~�:J��7�{�/*���VT�g2*���8ݣ��[w,ͫ���c����&C��)(N�|�.��9�&˿u�[�Chר3�خ�QzhՕ�L��x��X�@�reʻ�-R��6-:�.֬�`�5����u9��4U���V(̐�"
��D����qXRy�#qe�Q��$v#�y��Cm�Ò_cC�8�=�Vk}���{� �XR��nP��amJӢ}��]���Q{^��}��Ǿ�p�.�@��𗅜��v����Q]��{�4��A*4ǹ��}�D���<�����)��<m���S��0t%��ǲ\G9ZVz�B��yM��N�1�'tÿ�+�n��;{L��}��i9�����-p�V�aL�`/y=s�r�ݛ�Ǫ�E�]!m͓w�a��َ���G_��=B��~>��w�̓�`	�ݢ+SZ��$�=���Z7ѯ+E}o�#��+'�T{)o>���ذ�p-�Q���ʤn�����������.�:����=�o�u[��]�Uz�u�H:�I^�ѵ&P���1p��鯬�;_Y�{z���9�g}�}P��0�
#����s��^�So�_��,�}�A�p���N��R������tǃ�5��́QA�>�B�R�����_7�j2�V�?@�Sǆ�X:@)+��l�L���h�Y��	?�+�+��ᠻ�WNo�7;�Z���;���G׷b�:yAÖ��"q�TU.�.!/�`�0�V�7,����;5e�v!D�6L?e]�}t�[�e�[)=rl�ؾB��Cw1����6�:�ٺn��)mLʼ;6T���f���L���=۪J���Og#�\nP}՗;1�������cB�;����?ڟ��:�3~-�zW����0�N��z7e��EƢ�<�U=��=���9�d�;jE�'U�k�R�� nh��`�p��;�Q�KU"��N�����a�[xuo:�>.}��eڰk��Xf�]32xM�V��V{��������6cຼ*�*_��[¡�j�F���Y��%�+P�s��}�,}۶�VS�$t��/&H�*�s��Q	��Us�U�R;�RF3{�E��b��[(F�5���ʨ�d~�ꌊ��Y}����a�	�Q�uc˥�U<-.������>�&X�՗n��c�X�ƃ�����ʍ~�f�Z����V.a���0�+պd=>���FA�����ר�ЃίV}��a�cA�^j�NO��C*5����Q&�>MA�Q�#��Ǽ7qo��F��-dٯ��**�)�F�����cY{2½���Q��ѿ>X���S{]'RyQ�=��)�. ��u�Y�^���,�	����g�rl���f{:����3��i�Y���M퉥Ѻ�kg׿�s�J�c��+���o�n�Y�`�ZH�;~��Yu{���V��`uf[5�`��6-%�q���]O�/)й�6gR�U���C:���Y�V��
�0��]� �T���:��g�kK-�� 8�s�������~�a���Ug���GD�<��4�Dw�z׌ru��晆T�Њ�+q��H�=
������e->���ݯ���g
S-d2�6hyhu lh�����
����z�'�,�tm>;�և��W�+�]&}G@�a�PgW	't�%,o:�J�F��R�G����c�P������ې�z���PjmK,"K�1�&�GJ���m5/`�����"�σg�o��T��gѮC��E�a���u�0�2}'���9mǟ�Ϸ*U�y����m�ຠP�~7FY|k�0�%�H�O��7�E��v�E˕�Z�&zG��j��xө����\���g��#���9΅�{
�Ń�5�c�/�O��\��9܏z�̯��{#�����q�;�d\�QI����(�0���܅|���K�?K�Ñ��]�ъ6��.ϰ��*.���P�9Jh�$5�&�LG>�Q����_�,{�Jh��0�m���%���uHTord�|�-�uG�Q�*�k�ѽ2K�Pr�/��]�]_����vVv!�B-��wKw��(��՚�囔��S�2Fm�ͪ�4����Zs�et���	���t�
�JI#2���ɲ4��t��u��ٽ<����V.���z�LǝQ+r�N�(�R�(�ݾto&Ј:��l�-�c�\�(��-�z��3R�etgBP���U�CӼ����]����L/�q�<�y@���3��7	>��6�^��]f�i ������M�^�ǃ����9z��z��������C*#Z3Q8ݚf��gkg',ltc ��=,m��
Ⲑ۩zN�Ҽk諬��F�N�z7�-g��br�1�M��F���(�zp�����#�I�Ή�QgC���:.��'t�6�ݐ�}
�{��c/��Q����ό��.��m�ӻq���W��t���'3��������ɭ7N@��[}��{�JV�GOn��>s�&�3��-o���E�uA�QԚZO{Ru�[��7�E���#�K����Ф^�������z����]�r�(�ѥ�^��L�����yCH_/EH6���ƾ��Qe��4�����|��}ն��9%�/BB���~욯t=�	:�f��x��/�$��;Ft���v}�G����ǵ\>]g<�n������b�ju����>6���Fx	�)@��s2��ۜ�ݡ�<�>>.؃�b�+����C��n廘:��*����"�:�b�#��Y�/(�'�7#j�r�,�ӵE>�T���$�z�޺�<[��e{|�nU�]�yI錨���d��sz�<�ڲh��aѢl��!���[ݎ��u��4ovY(�htN��q��*=����=�3S�~��~ۉۊw~0��3��8 'Q@���4�c�o����gf��S �W�1�8O��:.q�g���\sY�ӷQ6e��n:���D@j���`�T�����ީ~o:ܣjը̮\T\*m�sj������s���͵`TC^~�Q�&��L��@o�m�����
wwޣo��z�/�vͫ��>�3��M�ւ��`~�:�*�����L"���p{�1_7�+��K94�+
��6�E���1�GwrH�\�%�����yK�Q�/�b�v�y#�],Q��`���7(+>�S�lW˭0�笨��Tv�Ku��E��'�u�w��:��c�S1��&���Cm:l\s�J�0��6�9>ӂY�s
w�xwq�L�E�!O;D��t��ᕾp�oP�>���Y�uu�4^�L�@��_U��^t������[<6����:݇֌9 {s�uX>����3!�N�c�b�߮��6���A�~*ꆻ�+рغ�o;ǅy2�uWzY�}E�9Qk@�����SZ��rLc�oӃ7^V���ީ�<-}�i�g�ީ$N����q\�
u"��mZӳ2��E�9���%��k���	�/��U�z�	�e��e-�k2��v��5����u��]Q�b@��hV���o�Wm�5���B�`3�;����^\�
�y�]�ڼ��M!�W­
��e��n>��^�޽�:.Lw2(Njѭ59�����t�ܭ��A�s�z�w�}��+quН��]��c�r�;MkX�Ҧ<Tt��Ƕv�#
=ڜ��X)Q�[L�z;R�F�{�VѠK��)/�N���R�,�1c�����O{SYɴ"����h��uܛչI�Y�h���VL����;OEa&w>�9�I���BLM��a86���XԸ�7YҕCDq�o�2)Py�=�{�T�h�I>v�t��I����� @�2�Y8Y҃�T���9��R΍'GfVt!<5}�4��{�(��֜�U{I��9�)�֪�L���&�VN�Oq�� J�s-�իgr�׵e�S�}�9Z�I�eؾnn�Dٛ{��"T�C׆wK_rvBv�m;�.m5Kz��ލoQ,�C\v��$��	�0q�Kt9��
�҂�+Ъe]gGR�ݳ�b��>�霪w=���3��%[�k՗E[����f���s�WchG�:AuSB�wI���s#�faj���VW^�i}P��m�'9�s��ru`#C�����;r���kX��G]��iTˠ��75,q����*�6�������;*l�V�#4�=��z:��\�u1�.�c_ 	��jn]���j�c�� ���`�ɻ|Z�/FƱf�\�|�Ӳ����\9��3�6�Hf�X+_5���޺���̊��guv`�
�2N�ŷs��2�!��И�lM.�TX�˭��]H�Zh�sۂp�Z���q����I����`��+��o]�F�T|^�ɚ�T�ؖi:WoKýV�Jۦ�x! �N<�Ƌ#[!n�>��`7KGsh)�s��x�7{➠�2��2��Q��Q�@�\���]��A�:NV)pVm,��`Vm
k�E�C��N��ӱl�t��ۭ�:��Ч
/$��Y\xɝ)�*xR�l�sg*k*��
�\
��I��cz�����M�øa��sݦz��R�I����n�p&�_l�Mحẑc%Z�-ܙf&\F󄭩!9�H��[�.�Jl��?K�w��s ����6������2,�(;���賂 v�ƸB[�����s�;!���,r�bx�f�j�t���qM]��P}K���w��j0h溇6�g	����찗r���0[�\AI�yI�a�5�ˣ��6��}+[��9�4�i %�e�T�TX]f5Y[�# �}�%�h�/���J�t��w�u�Ա�!h@i>�Kfs�7Gk�v*fC���>�IT����iV��N��4z���u	{�];a�+/��1*�!O$� ��]���p4>�D�4��4��Ҹ�]p���Yݵ�n�W$�	E��JN\�吹EF�s��s��h9���]bw;�W7Nwi;��;.���%���˩���W7:���ɕ��%ݻ1�� \���hGwι�(���Çw\��.��;�s���19u�]wn��L�������I�s����5%˻��뻹С�n�h˗w\��wA]t�6�.�����ӗ:��ι�:��5�q���]�k�� q�Ewq��;�ȧw���Q.��әnW\��!�����������7H�ۮ��8vr�P\�w;�]s��)%���\�]��N�5��9N�iݹHƝ�9˛��r$�.D�wh���u']�Is��昬PDR�e˓ "FI&`ɻ�bB]�9�Q;�MΈw(W�	6�}BWl��R��F��"�enWl�l	]I�w����R1�9\�2eq���ebʜQ3�\�\�=+y���=ޡ�����@���ph�GG�.��
��x�C���e?\wg�c�!+˗�ۆ�$�|�s�z��N��5D	���ى�7�>�,�E�P{z����gsm�)���2���R�#����3�{3�$Fx	�|��V����O�҇*�~b���>&��H�f��;s�)�C�s���a�e��l�K�<�}-�%��5��f�w�קR�:��{��㷍9Oi	�o��dڟ�D��t	-�14{�ϯ-����Q98���L���*�{��<{��ˎkNڑt�W	��iK� �M\L��~|�W�mg5��-ݢ���0�\&��*��l���f�V6�����Fu�T�v�a��yƛ��OG�N�d�B���F�<ʍ�
:���G9zK>�����;n�E����j�$�mO9�ul���QD��D��h\W�i��zj7�R������yW��o����f=X�.���Ôzэ
 (�~Mژ{_	�S�ubx��<-�c�!U���)�0*��K�+@vw(�ͫ��rwc2��1���mmeqwS�j�,�ɐV�n�$�C�έu����]N�j�ʻ�ޝza��`WS&���6-]E�Gz��<aoo�0��3VVw�QV�u���pnu����6-Β
���ݞ�ń���'	jB`�����]m���`���VqǦ��;B�;(Mَ�����7
0{�+7�3w�!�o�\�O�
�^��K��;��5C�'����HU�Q&������$o�*�rϓ.�fo�z�s^W��Gl�69�����ԗY;��3�Rag��W?+F����*�n:}��Jh<�_�762�y+4;����=������d}ɬg���1�j^�k��e߶���.����Z�=�9�(�3�d�6-t��a��k��k��S���ft^b�����ӎ�Fg���1o�-;G����� �
e�]#���V�f����\D����ø�d�ۣ��;�Mh}�9�F�Ux���*�Ǒ�*��R=xt��U�WK�dwv��/
���0��+׃5Ŀ�s}@>�z���Pk��R���$�3&�t�~�
qPf:��ut.���Rx�����Sq;���k��s�����t�S�'�{կ
���x�z(ܬ=j��5��# �]P(z|̂���u
�{�t�4��؎r,㶤z
�������žk]��r��� �Dچ�t��kި��']�%�L{�71*��NV2ͩӎ>���Ҳ���|/X��z�D�Ň��/[�!��Z�B�AӾ1�-�>�7N�=N.jŖ:$�u02�#wƌu�_rW�
]2��ڔ)�6imj����)ek��W9�߫�2'��A���:~��@��҅p/�ޞ�RF=���S͍Q��l�����f�c=�O���v��2.]QeI!�� t�
�N{�s�|F.����\�]�^��<��A��Qe�h��j.��P�9Jh�l��dEFv&�#�sY��ذd#�2�Nײ��#C�)�D1����7^'�=>}��`�w���5d���R�W�d�eu8 Ͻ���+q�g�Ũ�*�����H�u�*�L/�eS�uC����j^_�U8z��+�ͷ��E���x��z���YW��Gf�����~t�N{�!��<dIQ,�Y<g�7�-�KC3�~�ӣj͇P���S�M��������j��ǣy��nEї���=J��4xo�O~�X��7�׎~����?�����T�g�7W<���G��\f�/I�F��>���9����p�V3��9����U�],>��	�A�����4�@{��:�=�Q~�~��P�o��-��}�>s��k�0�ѱo���Q�;�fza����F)��d��]��gfn$���g<L�9�����t�9����%��e��˓�"��ӡ�Fo,_H�$���w��Ej��qS�2�.�� ~�i�]�"���h��u:a�����K}7���^�t<.76�b;&K�u�G�J������r�!�j� {ykr�!�0����/m���Ae�$�.}��*��+[�6���8�Ԍ�5�f�gFՖ�W�F��n���},_O��v�Iڄa��S��5�}2m���`y(�S=�
Z�=Fx���g��3�}����߇D��O/��*֦N�*�-fs�z t��\ �<��h71$���x�E\�hh��Ī8i���32�ދ:6���E��v�&����C�� l�� ⼦��dVx��t/s\�x49����G5�O�����~���SR�\$zde�Y���ؽ���ܻ�]��彄xZo���kIp�%�>���]3-M��I�;^�G���iٻ�O���o���8ͫ��r"�J���7:�S [��|�=�8�J�Kˎ=>q䃝Sɲ��
v�_)l�6;�����wE2�My���)�{ꂠFo���j/��}�B�jl)S�n|�:pT���0�.zʏ�k���T#3���W�Ĵx��u��t�7]���R�����U'�Ԃ:*�Wk2/ۗ�4��^||�輦b��m�z�l¤n����\dy���]�i&�n���f�̩��"}vn!*%���h7�'VR�JMٽ�={:�����u%c�U�� G&�v�_c���Q�pgW�g�{��	�^�ޑ�7��UD�}ckC���f�#�n�t9����2TI��^�b��CC�]��}��f�����B�Q��|}d�j��O�c�����o1#���ǗŤJ�>�kΡ	��2!U;�}����d;;o�s����7`ãz�쭿�t=V5����i/�o�ʴ������6Z�G��c;f�Z7ѯ+E��9A+��/�'�.(��:A���ng� ��y4������FkZϹLw��Q�Y�Oz�h��%VZ������?uu2�Ex>��򘸧#��r�u@^͢�Gx=�V����K&��|�����������L� ��1��b��T��UO��y4�0�M:>ۀ���w.c���}��D[C�T{��݅ֈq�2���P<�>F*'��ԃ�}o�8n�w�yT�m�=�4P�mՍe���r�v�M��t��e�
4���1p;*/3�N���4�\�NJX�f�,�1�W�����ѿ�zr���5ڑt�W	�3.n����߱j��3~��!VՙV��j=[S`ɕ2�Ȇ+��U����!�'=�e]wY·u�`��F��+��^��vk���+�ǝ��n=����ܥu�Ns�Į�m���e7&vv��*Չ,�f\\SL3��Qi�}�P�� ߇1�5rJ�Ò�;4����bځ)\&;
����q���_�.ՃPۨ�/�t*���ǳ׻s������RtW��'�n	��U+O��~=xT4�xo���,�1^V,�Q����׾����ܫ�W���Ѩْ;j*
'�V���{�U����LǪ��%OB�'��7[�%����m�Q�\~�У�@�Rѿ���'(˫�K���3�ײ�������Pq/1ׇ�I�h54ܰ2�]B�_c�P5�2v�L>���ugY���
B=�Z2�w8���#v^{�\,+�z�����h2��P���7(e}��E=�N�9�I_�&�߬w�Ev[�:_�1FW�ɂ���eE]���g�y9�^>�
վ�Џ�@��kqU׳G.̴��m@�u���_�K�Y��z��w�J� z#�X˙�� �����&G��#�����k�ڞ�;�1r2x+���tK#�z4���9Vn|�@ο��#��G�^�Fg�����a��|NeA�Q �R���9�;t�����^Ą��q9�/��(a�u9Y�n�U���uF��+'�C_4b*�,K�]�B��
BoQ�xUƬ�\�0����h�-U��%��7n��[�c��p�q��H\��B	e����M4+�ԩ�Q�g*T
��v�� "�ض+$m�z+ךN(hO�=P�ٽLO��l�N��38�t?=�G�=Fa�=HTha/T]  W�f���^�2,5�ڐ°�PȾ��o�mGe|�px}ִw�jYakz-	��q�Y����BW�p�b���3JgF�������M�}�C��[@v�z�黦�O=�r���d�^<.\ɧ@��$��gt�ì�7=�[�:��\u�F�^���\:��=5���#%�i�r��8!Q2Hn�T�<&�Z{}<~��]�FLqq�\�ݷk�Փp�^��a>^���׮�d\��͢T$�W�h\E9��c�\t�Yx����QU��N�c�}�e�C��M����B�R�5�$v��~<��E��j�]�ɓ�J/:����Mq����\��n�O������;���@�I�q�Izq]jwg����.c;Fʴ���X�<ϕyC�x��dwr�z����L/��P�8�M��cdP9&��t���:'�H��B�j��"�V{�{k���uZ}� ѯ��żf�l�V�����#��ou:��l� �:�C��>�q�f�>��(�-~W�wm����\Ҭ�k�)�i��ɮ����-�E�`u�Ni�9�u�e3:kK��TN��9[�?�1�gr��:��a�*�^��k��Ξ�"qE��w
�2��7�:��2��~W	w��AɎ�8����K�t�^=�Q����������z�T�u�p�d?ap�Z'=�T?�YL�~�&��&P.tT��t\R�����y��zb`�z}>��������m@��XϾ�)���Yf*߮�����n�a�	�:'�l��/����Re��rv�<�`e��F��P:9&�74.�;�{䰿����������,iqt�Gr�}���VU#qN@�j����[�p��{-h�gϮ�~{T��N����E̵�wȒ���.�U�������Cz�����ӪȄ-��C{>O�-H7�>�5~g��M������~�(UD�?���dL��O��JүZ~;�C<+4W�o��oϯ�bW:9r��b3�N���]�9���@��,� '_�&���$�㰭V
��ë�JZ��ևl��^C��_���}��ꑅ�����t�-�(���U8�2;}r�^MTnNv�E�N:��kG�y�|�a4��M���A_B�Բ���	�}�ymՅ�9n.v�U�7)2"X*�d�]�DP��P%΍;G4��Ԝ�ն�w~>i��=kA�m	&1Iۉ揷P�]%�@t�i9���̤v��+��j;��Ζ����eZ��'X1�9���d��%��3�Qmr\�)r��:��,��ħ���������+�ꅽ�0��0ϧ�}�|8�m��k�Ы�Rh��������z��}/�'d�,�f`�&�B<<�����
���7:�T1o�ZCĽbb(t=�a>m��U�>�\�b��M��A}.�P���j�YQ�GV�\kzu���R�w��	�E���V/�jc���#��9��G{	^�
��W��b:!Q>͕{�:g�Wh��&�}�z�jG���� �B�;*�J]����X�]�t�H��J̸��a�W�P���]��Dv4�r���u|߮���d��`�1�Z��%�q����j�狄����'��ǣR�w��fGYv�xW��t�����F}��\�r��W�8�t�70�L��>E�9V�?{^�is����c;f۵�}����:�4+_g�׸�{���C�U��äefP�Xy���<|�Dv�0�U�Tb�o��"�i��󮢆}d"�aA<EL�L\S��a����==�E���oA���i�1�rp�,����(x8���/M`�j.Gj���{I�2�\�fw2�h�6��N�u6DU=R�f��Z�%N�d)�՛�g*��w�WA|�N(Bp֟�����z+��(A:�q _r;;���A�ֵÓ׵<�{������t[9�?&�ޙ�7�l�>�� �1� �,\T�B���6��g>�2q؝�"�Qt+���/��.܎7��C�A�b:.�t�i�N��� �1�*��gPt��R�<E��|���a
��ucѮ_�F��=~�Bt�W�=�!B"(m��S+���.�U�� {��n(��Q��B���h��'�/�j/;jE�K���x�J��ϲN4���z}�x�4�A#L�j�s�Z�	�¶�GTo:�>.}���X=�Y�{
|6����J���~��3]32|7�R) ���5R��n@/�o	�К���T�liU^�:�#�T��t�3�%�O��)����h�̑�P1P<q�/�s�|u�n�9��ǐvwId,�I{�芈n\~�Т9�D�ɣZa���9F�]X4�_�V�O[�P���F��2~����|���qZMCr���5�+5����d�
��D6|ߑ5َ6|�G5E��w=�X�*Q�ƞ�v4^r�M�Cr�k�6������VPM�F��g�YeK���R
�$�Ehk����4i;V)\ϰU�?yk�{�dc�[u�ZV�Su�ѯ���2��[���C��KO��]�U��MѾ	�R��J�*ccx���=⍸0�/.���7�ҁ��ա�����:��{H�D�}ϏʟG��f�;kl���/�8�%̹Nt���`W� ���+�8��������槧�yep�N�t�`��#�{�i��(񗘙�����O�|d����W)4V�H��6
v`�,�ڒ3�년��!j�*�A�����J�fk��vK
޵;���$��m,�*f�s!��[YB�F�$kvP���;�t_Q�"z5�od7���䔤@Ԥ���֦�U��P�s2T�{Iճ��x��;�����W`l�Jِ.K8����=�U݅ld��Kuқ�H�VΛy�j�rn!�*|6r皹�}��8�?�+9ڰ��O1+'��X��5�.�X�d�r��85�z
o�RD�8`������eԼ�I��6:�:���ĵ�h"��kc��u�MO�w{�9vWFH��.�U�h�)ϸU�O��'�B)�w�p�,�u�Gr�����˾a���̐	ȣ.0��\lA{C�{�p�e�:4��S�����g�y9�5�Y�hiu݅Ws��ò]Ӄz6N"����<��MS�ig=�%��p�Ow�̤N?��Q��eŪv�f�.c]�{��S��oe7����x&R]q�3zN�ȓ�K�:�g^�F/�M���m�0�n[՜��ś�-�	��}�lͧ��J�숨��Fl�\� }�u14�`j;b�ɽ�*���i����2a�V���-�4j�.K$�͡�і8�ڠS��&��+��w�ڸ\�=DvA�+�
�=�sU��d�Ӭ,F%��i֚�����i�s�4����]���g*:ep���;	�\8�\�p��e(ݳ�5���o+	��}�q}��6���6VBZ<䱵Ml����w����.����KXtP��ytT۹�B/j[�`�a�{±��Zݶaa�
uz�fQ��r�f�i�%���u���u�M
�����`�v>�xh�	DS=M�W.��um�Ę�iI7]*����y�n��f�(��=Wv���c�k�1��7+#�5nhe/��-̠M3sP�1��A��t��Z*�:�{�����Ӵz��a��zƧ6���C���"�\��F5�N�Rۊ����s2���E®����I��g���An�<�st<	���c�G�U�c�|��=wj��wU����رY,��y��(Ծ	��n�P�u3pT��N���<�-��6$g��y�!�bp���C|`0 t�����!�����%����5�o�2�m��V5}r�$XM�4���(�meɐ���;['.��y88�0�v���ǹ}������u۹ڑ�p�e�v�w]"�swa4���Cfnn�n����C���@J��t(;��i�vv��ۂ���lBI��tF�N똂��p��9��-3��S�:�`� B7E8㻈�Ѳ�D]�v�0���&B��`D.��`r�0��Ph4)��$Nnb�)�ԐP�.v]܃#롙�dWuq ���Q$HRs��"19q#�ts@��m˻�n\iA�	1�;�َvL��%ݮQ#ݹ��˝�A&"X���PD�BR.����tƸtRfBRH�s�#��%4T)AL�I�����;����bW.�F�B�$N�H�w
L�]��1 b.�wWH78
�$P�����\��  �F����ʍ!y�5\�A���Z��k[����۔�Ef^Hp�{ �|2������5���nKG�k9n�g�)	>�P0{���ҋ�_�;��~x��ʮI~��ޖ5�|�&V) x�
�告E���a����f^ߕ�~��@�c���rg���Eap;=��T�d\����eFk�5uo0��3*�{�E����>��g�e%V�.�k�:-��h�DX�^'���U����m����ۄ�Q���y�ÑG���� �����{Z�<�������Twy���<$����Vv��n��r��Mhy�h�����]$���瓚�
�w[�)��(I���*g���7{RW���_A�}�[Q�Q���ִw�e��K�bmD�s.��;	�%�1�֡�#/M)��Q�q��l���!����;�+��r�Ρ��]
�fv�ܗ� �<�0#�#�g���Y��nд�<W�+���{�B���吱�����;�~둲�_���p��]D�!��Px�V���W�w� ��a;�5��ٛ'E��0�����G9�%��}�^��r�7��	�^�S����|v�.�_���ׅ]�PQ��t��Dǎ�H��df�u)cv�	��5�]ʕpS1=��5Q*�_1�lי�P)���hxh�4?:���˷̥��8el��q�G�Sڽ �@�o���L����6���ٴ�l֡Y�bc��C�k���H��K�6����-�}g�MCj.��P��R�5�̑�B~|�R��9#�~���J�䋏�۹Vxv�"#cw!Q�ɒ��r�ZP��M�ֳ�����'����;Ŝ��l\I||��(�*/�wr�k�SW:`a~�2��>i2A��uB�/^�K&%�Κ����a�KUٯ��-���T^ת;ۮ�Oc�=\�E�;�	���y�*g0�n����d��: �G%�cgC�N�ةzN��~
�8��Y���~��,�ye��ll1���8oak>����ߩ�M3,��I;;s?��:�S��	gI�o�ŰeD�5C͛J��ۨ��.�A�o:�q�g3~�[f*-��Y�s��z �?(zX�u�Tǉ��
Z�(�rϩ΃׵�Lm��E}���rO�s�v!�-����}ZQ<�D\���h�o�n�ཧ������@{Qi�5Y���ʷ���'Z0c�\�y��t�Z����O�vZ�l��IzAɇ�F^�G�o��6���푥�j��V��I_���}F�X;��WWO�i.��e�y(�LRM�-C�*���\t��cIӷ.�~:��0�p��t�k%愱�I���D��$�7ǻQ�<�Le�����"�쩹3!�kx"zA
����>ew^�����Nz�98*d��켤/7��%���b=ںb�5Z/�:	:�g �Tu)�ى�;Ǩ��_:vk�϶)\j�w��9[�٣�c�T\s��+�}P���hK-� ���0�k���\EL��ܻh�,��7y�7˽*��+��=����9r��D�CuL���)f���8�d���Ï�|6Vs���a����k�����P�mZ��~��n=���3�u��5>6ȁ��!��+ܪ�-W�����[@TA+Ŭ�0�oYf����/�pχ��m����(�11��WM3]�}�\�.g%��&��0�s��=��s9��
����h�6��W��	፟�w������n�k|��n�_5_�$}��/s���F���xʎ��Gl]��G�N�w�9q�~�Q|��:|�4(��x9��?��閾>=�.|��e���67�Qo�!s���S�8��b����y�o#�t��4,���u@����Z��]�aeƈ++�N=�ݍ��i��WU�6z�7�ƃSP�k��Cu��7��$��{*ĳ �2��ś�}�3]�yqA/��W���Br�]j����Z����w�ɒ����9����r�PiU/sI�fP���Q[F���<y�}ż�r�L�]�.���lsL꒠ �`TXԻ�;'U��`:�5n�Dø���k	�C�\n��y$g��yZ�+����x���.�Ѽ���d9�ط��s��"'�{+A#��9�=+پ$�����ڌ����!�;��>״ǣ�Ik#�X��ߛ��k!|=�w��Y�sE;�_�,'z&}�⍗3f����*�.��^��g�bR|]�{�[���-���n�3��{�[���גQW2�T	��|�%�����Wc��ؘ���Xwx{%��Q�ȸ�-��'�=�t��Q�z�gղA�X��2��J���v��B��.�<�}�J���Ǉ��4���q�P�`�1�;jY�Q%��):�~}��C��f���}2�yh�K~��>g���{�h�<�P�ᖧ��7�@Nm��������nS6٘�q |mL�Y���Ov�G���ӗ�xj�"�y�v�B�y��l��;:+��~��S��9 i��@���Ug�a�[�p�_��<o����};�w+��yKuW1����r6��[5n��������zP�|���~�Q��Gv.�ʺ+E&m̃��앐e��ZǦ�=n]ujҦ)�$K������r��\n���&�g 	ñ]!xD�f7���d��$t���Ō�z�e�/5d�V�f�}Bs�Z���pbpiJژoHҶ�NB��ǫ�������Q�9 ��u5��U�T���i�}���zK,��{CV�j�C�e�{2GmDT��(T.��E�YU,��<"����BH�uEk���F+{�C.����Т������ڈ�1���������M��}ђ�%�?�NYU�΋[�V���T�u���nX�ơY����d�<vKbW�+ܺ/n�;����������\,(�W��k��c��ʯ5C�'������>KE��������"�͢N@��6n�:^N�#�M���լ\25$��y�5�୛��\�o����n���=b��Z7�|�6n��1��Wм��u�f�@��4�gk)B���e{`K�/4��Ō��Q���k�s�S���8s�,y@���
|���t��9�â\�D�h��vj= k[p}J�01׭��Qw�7Y�*-�R��>'v���gUCf���x��'��ly-se��4�}r��E��}��~a\?&��!5��kQ��~{t�}eS�3�'���㗜9n-�A��O��)z�jB
���_D�7趘{���螵����PL���0�?j�����ͮ��8:2��!�`ME	����2�9�.��u[7�U�ޮJ'�W��BekZ]\]MfmM���t��9O_6;ܒĽT��։���]ȅJSag2���~�s�'d��+�N�`�]���;��N��>+=���{	sE�6I�f2��B3�d�7�w��Q��l�1�}9趀�;^\���g/P�a��+�zNIw@	�D�BU�z[7FQ~8���\Kv�׸�2�z���p�P�q�;�x��۩P��=Жs��<�@�n`X<�(V��t	�\�'G��*w���x5�:�c�_��f읇n�n�^��\�gaA�@^��Z��}W�A�;���T��m�[yD=�p���g��}��ͺ��My�*�R�52Gnׂ�g�W{;y�������K����Ws��͢8Wv�C��%�<��:��(�O�}�=��$����og�␗��d��G)B��V�"ٵQj:����ښ���W���>r�H�n�������e@�7X�^@6<����Z��#�Z6;��/k��]V��C"�fvjno�S͉QHgx���}wC{�.f��� Q�9,+����Ez�mԽ'M��x�d��n�e�ʴ8x�%�Z�tk��]�;N3�<I���)�M3,�?9'gng�T6t;�*s��-p�
�zK�v��k��v�]8P�
)u'SHQ���k�ʒ�jkp��s[�/v�h�l=8l�����k�t[1�x����8����z�Ƀ��(\�gB�[�bV�ЗO��^�=E�Tu�fL��+�� �^I�F�&��YL�RudN���E\�I5�r���AL��=��g��3�c����x�78Ng�����3Rm�!k#Uhw�vi�zU��Y<զ�-\}����v�5�ct�y�!q�{t�Џ?pO|q��0��(�rOy�f/���s:qt���� j������N����h���h�j���sZ3kfݏD?w]�r�(�D���3�:�F^�G�o%��<�Q푥��9�s�ϪN�E���p�-�WZ/�ʶ�ȹ@���.�C��Jb�ԙϞM3F��@ګI������=�1����=��܎9M�C�t�e�O����3�O�J���{زv��57�u�/n@�S�n��g�>]LX��u�o�8�TO���a�g��Q�@�Pg p����y��Z��}8S� o�*�F۬W�ݵ�u5���k0�mD���']Q5�T�9���*n..�g�ϧ7���	� X�{@W�����L>�[�C����_�2��Kn|][|)�ヱ�u��ʯ8NJvk�(���g���i�w�1̯��TuF��F�����-MN�,5����k|Fc>n�]�i)K�6���K��#��;�ٷ�b= �3��Ip��~��l����!�ݖ������V��K�Ѻ�I����/�ҍ�ϧZ�] z�Mi�q�|z��m�n\�=�r:��M�
��Pfs	��$T��9S��4������ܗ�����=�G&���L*�/M�_izw�f�h���ն�z�K/Q7/IF�m�1�+�F���N��60���Ӷl{��XF}��,lԱ6�c7T�r9��mo�'Q|����t��4,���v<c��󙘷=�N�N��)ܚͳ�x{*�8{5<�{�ƃSP�k���M��������I7d��[�Iފ�q[����9�2���,�>����WY\=�uX>���ϱ�r}�X�����?���P�K���s�fZ�ma9��1�"�c���#Y;�k������x��9�Z����O�:=	m�	��*�����l\o���':N�&���qF����G�=5g�j�<�˧����*nߨ�d�π���y�8iGq�&�;��o�u2�J*��c(L�w�L�LO�7�8��Udy,0Xu���~��%CH���(
#ٴx�}�[;�Ojq�iϻ��׎Z�
�g��,�X�j,���N��褴��ϧѾ�;����p�ﭡ�)��y�<�Ltg�x�q�Oi�r��O��.�M�8��{y�����BZY0�P�D9z�)�W�t���í|��
��ei����W3v�&ug��QfEC:��t�:uB�TǙ��5K\�yWN5Ї\{M]ԡ ��1n�\Du8���UնwS�ƭ���0�V�rlԲfWF�"yw:%����I~;S(/;w��D��ы�>g��8޻Z&�s�P뵗�}-G�ج׻^�'�e�;�f: ^��g��a龿z�[X�Ay^G�!���75>}�c��_�ҕ_=+ӳ�G���`��J\��@	�Id�P#��U�a��\<��l�T#�<�h�q�'�k���?�����E�C�L�䔞$��|H05�
�_Ȁ|��#Oq�,�ר�J�C�w:�C/Ie�ZN�Հ��e
�GI#�*
zq��zO���Xޛ��ÎɯM��D.TC�m]ы�߬��������=�@�R��a�ڞ��zzh��3�7w��<�����t�*�X���1ﻺ�
�����s�?}ơx�8�1G����v�y�W�/�x�2y���E�jn{6?3�ʩ�e5�|��Z}��eW��Ӓᷰ�F��t��ź�eا�Ԋ��D�@�v�w1����d�ݝeE]ep�jI�οz=sMo@^UJ.�t��{ý3�[�y���ѷ�A��Azg�sc�y,25����."5�4k��)��z��	m.3.���ܬ��QBkqj��1��0 ���͠�b]%��;����w�au�0;�`�I�C� �Yz��k;��c�⤎�\3;3a��1�����3�WqI[۬f!�o��Σ+��
m��;Ix��8�$������|�CR�p�&��sJ3=�l�[�Z�ܛ7�L���GR�#a��˂�����i)+$1.},	�K �*������Qvڼ1�o���(��3�Ʋ���do��&B���C���ǫ&���!���A�E��}��~a_�ɳ�Mhy�kQ��~{t���kޥ��;A���D��1�k�=^S)�rwRW|��g�m0�������R��[�֞�ۯX^ڟ�I@�@��C�Xȉ�cx�L��{v�8�}6�V֬����Ϭ{^Q��`]���r�a�O��r Nk�<�J�ǋgh�/�=����&<���;�B��[>X}�;����ë�둷^�e��ӂ|m����6� s\�YJ���~���9f�gQx�|��n��X��f��Q7P�W���K:���9��y��uXU��+"��n����:����*��d;��l1�-�|�}��6�2�j�)L(���>"�Z��>�A���	gm:7Ev�\lß�z�B�'R+��q/��*���յ�m��յ�m��U��m��kZ�v��km�mk[o�j�ֶ��յ�m�⭭km��[Z����[Z���z�����ڶ����[Z�۵mk[oʭ�km�][Z���5mk[o���ֶ��j�ֶ��kZ��Vֵ���kZ��b��L��>ئ	v|� � ���fO� č7��>kQM���k
I�ZeQ6*ٱ��M�Z�i����[|�'mT�ښ�4IZڛKmѨ�˻N�Y��&�V��)f$�`�`Zֲm��͛.)ҟs�im[EUk6�+z�鱲T��K�v�'f�]uѢK��[a��V5-���M(m�VR�m��[Um�ɭ�ڍ�v仇t-��+�����ٕ*�2��j�Z%��]��WVm�6���Ʊ�f�[Z�]�Z�5;R�m�Ye���6U117wG,E�ZnƤ#v*�ʤ���L5Q룩��˝ƃ�  ��uu��rϪz�]���궠Ηhӳ���ӓڵ�ݼW����C�uk{r�;qT��WwAWZ�T�u�n�֪��M��쩝wVJ�3m����   m>��N�n(�%�7�Ը��'�=�f�z(��(��-�q�EQEQg�qEQEQE�n(��(����qТ�(��(�zp袊(��ܩ��(��7Ng�i�c�wm5����ۻwf��Κy�  ���J����ǔ�r�*��tp��=�a�5�ӝ=�N۽��۸���;�QRC[F��v���Ǽ���]���mL���շv궶�h� F�   ����gZ��z��p��W�g��ʼ��cx�w��iA]�c�z]��k٥�Xnݘ����OC]��Ps�������{���lvd��^z��խ���v���F�m���3+Y�L���  ����N�nq�랫v;w:��Ӷ׳���Chm��@�wf�*�f�kv�;�5�u�K���==z�7���z���v�ݻ�ޏ\�E��u�޽�Sѯ79��f�^��&��J֔��=s�|  {�Tձ�ns���l�)�:�����T��^={����{k�g+7����{i�罁5�Tft�;u�w���{�R�Ӯ�V��v��Qu�czhzm����9��㺵�Ve�6�3V�  \���S귥�3[M�zt/v�v�������������]w{w��{O]<���^{�;Y�M�W���W{I׷����5���]��=rۻ�٥ok�w��ۚ:�[SU[Z�j�+U�YD�  F��:��ۧ^�,�ک�v��S�zt�Z��e����;�κ���C�Ol�u��{�j���w�{�y�^��w;n]�w���]m���ع�ӻ:uv��y�M���V�=w�ηZ�f+W�  ���t�����\s�5MuݼgS�	m��:��ym�u��y��٧UM�Ӛ�n�^����ާ��{���5�ɨkc�nWvu��⽻e=$������U����{%f%5�mM��K�e��F�   ��i��{�zk��򻗆�o]�u����z^����9�[�tk�ݫW{Hw�����i��m�f�M���clz�;8m�S���f����]f�> ��T�(0� )�)JJ  CB)�IUOP� )� �*   ��MUS@22 I��zb�jQ�z�e?��?9�����?(�&/��XjA�c�:Xp�=���<��z������$��!$ I0�		�BH@�Є��$��B�$�BCc��y����?�y�����ޚ��eQ|u�[Y2�aʆZ"��F�^����L��T�hn���+[3{
�c�t�PU��F�l_��t㵸�0���m8؁�H�[GA�n�)n��[-=y�������	up�G쐺(;�o`*�2[�w6i_J��O0�[��8��b���}c"�$f��_ff7�,��iY�(D56����,�b`�m&��lb������y���	
�^7�Gb�$�AA�@���f�^����\������ŵ�<��#�/DD[ ���a!�i�%��dÜ�h��Q ��cN}v(�@c�YDЏ&�e=�[ha���+G�K$��x5�3�-�]K�VP�����s4L���ȶl��E��;ǀ�Q���k
*���62��Y��Ә�L�A�V��b�:��Ŏ�ɏV�=ĩ<n+uZ�<�{���1Ĭe�׮٨"�M���f'HHAw�F]�wJ���t�y �dQ�T���,�EU��U�(��Y�/B6�cm�c����gLÛ�J�n�i�&D����J���r\��P����ģ6:�S�������f]m�gfR�	G~7vjS����EnR��5��^���L�V=�[0���n�3��r�*��]3�혣���4.�`��,��WL��X��rMT��E6�Pwx]�c���~Õm�n<��7L7S#���f
;uu�J&Z�l����ur'ܺ�h6�mn�*�c`��ٲ��a�P���hr�|�]��k�Q$-�1�"��!��KZ�X�Ƶ���A�������XN�eE[�-̎�a�m\X1`i�q2�#�%�kP��Ko~O3R���3u#ԻI^��[H��Ղ���S������oI�aّ���[$���z"���I�m
(��m:%bp�1���
����nC�Q�̄�T��r�^23(P�CE��n�Z̒����{�k��O,�	H��Zg�G�-S]�/3j*�P�3�h�%���B+Z��2К���e��ڊ&qn��\�n1pѲ�*��<'Q�uޥ{K1��PY��]�l�v���j���n�F��akEĴY���DԞ�(]ld!D��b�,:�l�df�����f�m�f��(�p�.S�r��X�E�.�����L͡q[z<�"�!Mݖ3Ŷ�k�F����R�3&^���\�X�֠��B=6�.+�^�VL�ҭ³�@,a��+Ǯ�7V��"�޽c$�O6���U��[Z�o�4wH�h^QE��X[0�&��=K�oK�AFcuԉc#��u���K�B%]��QS��\eD+sj��(	�ĵ��l0�а����\�#:�X�ѹ�� c�e���tY�Vj7��'�9`:S��Q&G�c��,�eKۢ�&7� �4*f���\,F΍�(|?��V/��%[vr��,С�Vali�-�˰�#��1k��Z�m�v����Y��8�Y�� �4�$��3jYg^-)×��@3�\��)JI-�ܺd��\����8�$���E.�n��m�`F�u�̼�i�7��Y�R��Fc�q��5r��V���>˨]��T4��'�T�Ӗ
	et8����	
ݓ++SZ�P��ި��΅�*9�oMܺU5��$��6V�k^�V
b+G�k[�y�	v^u�f�U���HTLи���9�E����ݷ��+2$�h䢕n��i�ஜ��R���,�HJd`n��P��>�b��턇[Ǆ���q�O/(L�MX�Q��6�9z&B�%J�Җt�tc�:����KW,w6Pl`�]a�Wy[6���m<*V�A��/lʺ3Y؉�U�͵��S�l@�+/w �a�g&�WǗڳ�?��:�l��ZYxH�6�3g���$�Y��K��Kl2oqel8�
��p�&-���
y�"�`ve`�,�:;�]��E�X3�?+��PU��F�H-��u�x����b�
ש�v�ޭR�bŀSq#[R� �I�o$�m��l�5VV(�V Le&�s@ǫ-���H0�	°huT/�C&��i�OB�{���f��C1H����PHp���4AT�{򢤱���;�RgqZCj2\��8����^	�
��Ƚ'���0�t�Ɇ��ʫ/�ѥn��
��j�;�`�A���y�jN(R�ZY��5�Ř��ʂ5tvl��N�pC+u�@�EC� �@m���0��P�fQf:3b�h�\�w���!"Yn���T��1Y��0��EY�56i�񘘉P��t&i,�݌-^�$�v���ȦPVu3�-��L&5�� Ud�b&d�� ��h�����TjHm�PFܻ�%���A65]e��O��6 �1�o�G�87nX��K0��1A���Q.�IZr��`L�гI�7VH�*�jM��!���a�Jř�9v̦֘Ȣ`g.�S1,��C�!���SEnYXa-�y�u"��b�Yj�C�`f��ml��d7b`���Pؤ�Ɠ�Yr��I،y��knr:���.^�iE�Z��5��]5��n��I��SckI
*��C�"�H�u[�]��-[0�1ʙ�f�lkB�!A>V�8��`l�[rҚ�'�^B��p(Z��;Gh���\������1>ݔ�P��q���j��q�J�M�I&�vZ�Q8$iJ�FhZ���0����S��e��̒E�֐n�
)�e	��<֭���'�!��!N�R�o3q�*�0)>\��o��p]��[�5��Q�7���y�uq)�ki2.�N�m]G5���8�¥��t���9���A�:Y`I�g)�ii{�c�Vu���Ʉ�u��v� B���x(l��#hL%�2��ئ�)�� [��ۼ-	�괷mݕ��MҼS;�"�)�LF�4�eiR&�˷�\)e�d�^\؃��솤��7f;zՆF逺B��3��S��r����ٟj7����2P?m9f��X'e�.�l �Fe��:��g�[Q�w['Ưt0��۷���`���0��:�%�W���ѩB�6E�-�ըG���S����ݟ��J��))-�s&����-�5���t�Q9��V�Y8@d[�ELRC��kX74kU�����Y,�1ŷZ� 5*Y2�Å�nXJU�u�{��"�ySC)e[8�ȥ$�JF��]���e����&[6��1�|�sVD�%A��SWH�Ք!�$��T��컠R2��J��f��1����UcXc��n\��n�F��#ZT״�:Q�^ؿ��7���4E{�it\�p�n�f��*U��R�3�f��ytS� y�����da���R�ԉ�HS��v��+H���Vli�[�Ӛ�|��2���P���l�"`Vh3Dw��W-G �����ha'Y.���L�+C��)V�G�І�`���I�`-Ӏ̓.��Lb�gP�Yj��֑��]KXkV����R����ֿ�[Wl��W��8��ݵ.��f��TLni�k6c�&�J��5k״�"�e,3U��a[3v��*�-U�4ۘ�5mG%]-��h:��aS�W�\���5���ie:�y���v��.�e�1:Zvʲ�Z�����B�ݻC�P���'2�PI�aL�7B�C��YN�B���:,m�ժPFn��\3-D�`t��>����!W���c^a$츲�=�P�N�9�aX�Ju(�[3]���2 l�v�r�㤐Z)�[��V�5��	�$a˽�vdZ\yE�Y-��֪-JݓG�L����˰�}�oe�en���VV�,dl��C�"�;,�X����f���Ҭ�F�4�ߚ-�&µ�Y(c��*j�j����I`��Q1�Tiec��`&X\�E�65z���u��J9�b'�/@T;������&X�ijR�L��[2ܛiB���T<���`n:4�ˡ�4<[��W�C%U���-CX�n�X��C Ԡ��Օ����!�X�X�ܲ�����PAn�9��Ԕ#âj��*�E�h�z��a��m�4B����h�DiTݐ���[�q쬏Xq���!B��'��|8� ��!'R�j�T��G��Z�,R�U�BF)ц݈E�4r�#3n�h�u��c���h�!��_�g�q�M�7�)f$�`v��@��Z:Ec��\�t�-��
�;EMةե(���z��� �����ʰ�o4Zٯ�tȚ�m�,
��N	�0�i�� ������>��!�m�w4Q:�ڂ���
F�Mo�gJ(���B�P�˯��ńZ&����7�UV��t,7C��d���.��f�Xn�����a:�X5�#qn�$���[�5v�*�ܰ�U#�kVеc"YT�����#��
;}��`Hr�^�T-��3���
�p���N�W��Cl�v��J2�h�KR�H��Í�L�(K)Wx6�]�r�65�`���S�J�m9��.c�nY�m#͏뱓l�{�u)2�;��@�X��i�A!��Î�(�E˴ږ���k��[C$7��kM��k]d[ZA[w(��b�0"��(�33PuI��7��R̲�mǪGэe۫��>�GC���B=�Q�ZXyd٦hD��&���v�/�ӛ$	��[�x������Y#���D�A-�U)�3��Gf�k�-ݪ�0�����x�K�����m7E�!0f��aq	�f ���/�&�F����`�khJ�"���[�j�#б��KA���J�R�h"㣥E{z
wx���UY���#��qn5�� tAs[z���9,m�$��F���֦�s*1r��M�d�#̚򥃐���G���b^�����up��wIM�r�i(�0�ϳ/-	t��aTv����ֽn�)�@�	}:���� ���c��͛0*'7l� #XJmm�q,�X[m��Qѿ ��97��w�3mni�o
��AA�Ӣ�]Џo1[�0/%6�bb45��^��n�x.�)cf��2�	VqӍV�aЋ%�l7�轅<0�Zl1$/	V�%F�]��mR�p�i*�xLݻ��3YT\���قT�u��I��R�޽Ŋ�h���-6
8р�ٸ���`���b��1�E�J֡#�V)��#C	��S;��LV4���6��Dd:�)��X�(]3PY�zF8���^X��<oea�E�H^�٘ݬ�����ɠJ��+M�*ؓ�r+t�F`66�H�e�V#x��4���@�\���Mm��K�X�,B��]R�a���������R6!"��f�R"0�m�Tk4`D���9+�Z�7�b���Q,)�,��˹�a1��Y��*p6U�u>�1*m;�DG8v��U!���KT信P�) B�l�H}k��3WwB���ʇjGCOl
�F��B��0�z4���*�����2�%�Jq�.��a�Y�fYX���"���i�,bܳS���.!�q��.�!�n��ʺƶ�"d�Eڛ�e1XҊ/-#���d+�Y(h��"*IZ�2CFi��,��Ԃ�ޠyY�`g4Z�J�{5jf�L�.QÎ�e4�4��(=Z���gF��4Z�2U�6���η��1��^��v/r*�JV��cwK�
olT���Y��)9#ͫ���X�)�Kn��'��n�X�#��ꓵH�Y�q��U1���X��cV�Zʽװ��,�u�)K2��Лx΄.���9�5��Q�n�'2QaF���m�±���ϵ�	�ѭv��B�.�^� X.�t�X�b3[�H�,1�k~�u>DZ�Ƒ��+�/!�2�8EHو�9p,�P+�
!���	��,��H'^^�A���T~[*�5�`�;�Ad�JJ���(n;
ҕ��KAW��u`�j�i��֨6�)a�T�ՕVޜ�B2FT�0�<����1�� �,�.�Ր��2���u�SPޛ(V�M����h)F5�m`��t�Y�(;U�B���.E^Pɩ]f��[em!g��]c�6�����:^�Q^+U��&���:���ή���`bӬӰ,�0]m�f��g-�v�n�
0���m�vP a�TŃ^���AXǸ+vFs� ��R܂�M�z J�v]���Q�ܩ��Y򺺴٨��vm�b�p�ͳy���B��LY��[t����I������Ue��l�=����bP=F��e배҂T�fBƩ�o6E5S�*`�E������#ֆ�@CS,Kt��4\�<�P�!Z��4C�X���7S۠�i����i��N#1�4J�0c6���L�s�;L͋�5^hj�12̙�RbV�V9a1h�=��Eз"W�\���^�Bm̫(UÊ#�zB3j��oi��Ư;�=�uO��u�>� z(���iP7GwUY�Q)�G(�w����P�CZ�u[m�˦W���Ѝ�gm�x*����R�";3搻�F����4DBGJ� �އyX+^.+/�V������ ˼F��7V���d���Rot��E�5�@~������L��ˤ���!T��e��x�:�l�e2	{�S���s�Ԥ�^
�l�ɉI�x(ͭ���@�o[phQ-�F�whux����Ee3B
�yJS.@�֒yHޓ���v �MV�+�1Kz�e������Sʶ1Vېغ���ܧ�������q���=���JΨF5�*��47H�!潁�!=ʭ*���J�Tz�DZ:u����O6����3�5��8l(�й�ܽNug3f�`\K=��{ Ov]<L]���s��R|]f�Or�}� �s)���5n�ʶ�)�����qv9H���ڣf\/C��f�/�L��*vAQ���&/��x���2���1;T�mf�y�uԖH�2Y�Kh㡢�w`�6�2!����*ӉG�+�S��k����+��c
����H>����!���waT��%�-�Ɖ�>��0L��@��m؁+�jY�AJ�N�7�֬�BT�d��0�T��R���a��P.WaTN'���v�d���=[$�7'�:J��L+����#�q��l�7�%��g4a|�/�R��tN��s�F`#q�cA��-e-�KY�K��\W
��Ǧw%���/w>0��;��d�QdclROX��(w�Z�
d�f��*v�mL,�edy���2�5CnA���o)��N'��z�ڡ�Z�t@����7��ՙ�U�n��ЖVͦ#&P�b��v���m,�cpl�T.毡�!��v�V����7a�'�/[=�y� u&��c�H60�[q�LqL]M-ŝkkkEN�5����u�sc��)�o3kwd1��au1�6n�f:�du.{:��x|�l�˺)��Jv 4#/2�ܸ)DG�R+H��k�!� �)�czާ������j�;N��}z��C�A��*<�j����7/2����+K��d[nx��؄v���H(Д�%��pQm�k/Wp�����*�����~�פ>7s��;X!���ܽ����1Q��,j�@<�=uΐ�R�NL\�5��#��m���}Lm�od��J�|ZG%�Z5=��s3�X:�)I�]F��n_g2�}�1}{[��m+3�]�0+E>Ӂ&-����CƏ�_V+Dt>,�C"��2�T	m-�Y��XT
��xR���^r����A�����" ��'�k�s\i��=�񹷸��\Ӂ����m>��^Y��A�h㬵�)Ȑ6��uh��S�Q��&�,e�Y+{�_j���RY�2,�
/H����Q훉�@;�
�k&�v��|(��h�K}�K�cŽveZ �Vʊ�*j�􀬧�T;
�܍�nC�%]J;y����1����i�ڪP��w݂����4�I�%��oj�����m[��ۅH�kr�od���{��8'4�q�j�+x�k�j�3N��%�Zb���j���_u�Au��N^�OI3�'�I����I �SGZ�l���P�q�+r<ʞ0����*Pq&���ژ�,moQ��ّI�.����û���e5���
�p'� ��us�ip�^��$���+>�Ap��o_)pٶ�Kt�C�3f���γR�u��(od;6�S��3�B�TO��3����]O�L0�<@	8�u�I����KBZr�d�[56�L`֫�:^��絍`t�3�j8u,����r��U���*�y�Q��y�+�ݪa|UL�Z$�O5=؋p�kw��իvN�3�h �κ9i�YI^0�	Հ"��asX.���S���qsЛZ��5N���<�&3s b��މrP�V��Vq�n^�aJ[�czfꆍ����\�V�,�QSz�k�Q�>�g+��tG������A����>Gw	�m;��P����ܲ��;�9�G7k�ݧ�/����n��{����x1=NsQd�V(��t+E^�iީK&�)κ�b��{oR,\��z�c��:���w�V�#��@�G��l�gʄQ��*��ps���"��ky�h�[���[I�R"�n�FOS0�$\��vekA�;\fsV���$�IJV��X t�CԹ�X���^�Ju++�h �D1j�|,M������{]y��x���0� ���n��4�U��.^K۩ݳ�q�p�� ѝ�S������
���m\!Q��7H�laT�ܩ\X�m����참ud���%(�W2�E��+;V�`�s���[|OU�������"��"4�@V�!C�1�W�ƛzV���A2\եi�Ϻ���o%�A�GfVB7�ؗp�Ҟq�q�踻-��4ɍ���]u�(�{��5.s���/�c��˳1�_`f��èg,A�-optq+�Фm�����h�]�Q� �/��0�T]NL��n$�4.���N�O���>2<y��J�(4Vn�J�\X춪J��k^t�XL9�Lkwc�C9Q�ɤ�hP�jol��9SUn��~�`��MV�<$�ܩ9A\z�=7�
,噗�����u�ݠm���	0�ef�&8Q���ܛ]�@��VӺ�8�QWq��F����2�2�nK�9չ[���aW��;�l�5:-�8N��I�t�X�45k.|^ȸ��
:���L��G�ga;i�d�j?�	�4���_!�,����]6�C��Av��qA�)4��E;��:����r�ʗ�`�+&R�qZ�R_�w'��=�FH,���+M�|z���OkSr�t�C�o.jb�+}wZ���w6���Ͻ��d�^��>R�42C���HiW�P������K�oɕ�"��S��41�VQ���������X2L6��g����ޙܣV�;+}���T%Xp��t�ܣ��tm̾xm�v_#�@�&v���63���$'��̲�G��E���W@ݍӻ�<��zN]B*j���T�W0�t�0p2����j�iբ�wz�J�hG�rf���2�U��v�������N���+�5�5�e�3��uՑ��6�|/�\���cv$�"�������Y⬛�G�!���m�{&t�
��XN������+OT;iۉ������O�HףL�/��;����=�?5��sզ���u�mߊ�=�&z`4$cN�%��_ѣ�q�"��}��>DgS&2�.VeXc��q�*���/��!�{e�v��!&:&c�Z�p/;�hLw
��r�5���ۤ��}z�1�;�:-Í�b�J]�m�p ����Ă�9I�i�S0�à\GM	ԜU��Y���⩏4��Ge8�>d��ӕs�粨y�lL�u�cC�K��<V�ѐ�v�Cr7��yծ��t��ұ���=dt��oj 7sq��Ȋ�0���6T����V�-8���0Y��I��낔f���ݏ���諝[c��s�s��(wr}smAB�l�V���&�7�-�IβV��fk;t+��6R�����zZ�x��5�̎'o:��3H/����"�3X9�6�_6����5N-؏�D��Ш\j�Ҽ=k���<�zu`�u���S3l��B$��}�	���ja����򓱅�_c�6Љp�\t���x�*�c��qk�{d�-H@!�J�ĺw m.�V�5��g�8�Cow!<�N�����:�+4�s��1�\�KZM���C5�9v9��k�r}�S�aﶳ��n�v*"	��\���vM�%uu)0r}�O$�Ʊ
�Ɣ�'qN>��b��nf�����2i6����/���G����=��+���$˗Ӭ�U�iK;;�{��n�jڛ.��d��P2�Ie������/�[[F��o����n�c�V�U^��C�C�ԁ�����J�Pۢ#M<[YϹ+-� ��\��~�to�i1M��P,�O�`��
� 7�b蝗��72^L֓n��e���m�1.ؕ�$�Ui��h_\���櫈__j�P@����#:̚)^��v�'҉D�j2a��sZ�0�^Cłށ޻��X˸�3���e����"�,���U���ܥR����O7앺,�d&��F�Tgru�726��n⮨&����4�`᱊��9�
eG�tZxs�L��r�]N�xp�V1<ӵ��G~{�:��]���.�>)VV���ϣ�OVV(�E����Q=j��WAJ��K��%C3U�vDq�8�\9)|�S�*N�A�k�ʂBw�i���JP��<��t���l�]��18m2-oj�ס���v���(ҩ�Go��Lٻ�^5]�x�P]j���ɲp����˭ڙ�μZ �T���O2�ȥf��yb���d��^����A��W��R`�l9S�P:װQ��3~7�Smدh7/�v�k��D�9U�R�t�$Nv�g���D�oZ������5�q������U�.t���sK
<]�������)@-2�N���B���8�(8���Y	J��鱁�����@ǌ�K�����A�y���D8��h�¯��7�Y��r��m�5.�n��eM�60Kոʶg�4�_G�+w��6�r�f�tk�
w���W��L�'�����pX��1�Rӈ�����a��X��G�(V@M�' ��A�(��:�7���&��q��V �2Lzw.�V��{K�H`��b������f3�%=b���8!׆,����+3�f���d
�EE�@����mW!��Ћt��r�dŕ�R�b�Ճ�����2��ɪ;�j1c�q�O7YiV&E��[�&��P��(�����О-EL�+��am�ײ%Bw��0��V�%b�f��H��$��wsqր� 4���5�*��T��jL�z>�����,�z�����bU> Ij���B3�ʕ�"�Kh���ܮ��\(�v]LA�%�+cj���
ڲڔ�:������Zc��t���m q�Z5!��o�|�ʵ�d�I�םKt�-�%sN��DpS�ۡɽX����ǻE@�ұ�<f�2�fҎ8��k�jfu���ų4١��>Et�P0�����:BE�s����-�_f����74��f�,,����N�/6�@�ȼ�ms����p��U�Y&lmKĩiΤ��ç1����u�bvv�pI�V���\�[b��,�i��WK���^Vv �Is�o�F�J�@ɔm�|K*�ۏ����:*VK�"sO�U�b��m�}��mxj'�3�W[�ӗ��*2�-�3F��C"9]щ]*�mwao�LV
�.P|yQ��֑!��\T83PÌ;e佫f��+�:��Kx*�82��2el�b�QQ@��+j)�#a�3e�\�l�`�Y�fఴ�o0�"mwV�3�ض� WTVx��+����=Ӝ\�v����yd�Ӳ�ɕ��)\�m7؅��B�e�����]���TѪ���םA��6��2&EvZ�H��8�QˍBLds�Bj��{V�}} =�o%e囖x��IG��&�,��n��9�U��#2�y*�p�c/�����I��UX��N�q'�]�1_|�^E�q�:F�����̼:�mǢ�X d�Ð����C����lcc�m���B��m����h�}8��"dX�י��8��#���ƞ��)]vEr��Z����\ut�@��
�/�j�����l�bsxCI.��ݰz�VJ��e�%uS�ޢYqٷԍ1[��+)ٌEw�ư9�뀕0YL���7rc2.o�����-	j8���}�d��ct���8;uG�t��0��MU���J����sb`�����)��n���.�/��U��If�R�;e]�'E���%��5V-έ.��r���� 6��{/�v��4��x򗪠���7v�������,#����_<O�Q�J��ΤL˘$��Y�f�s���.Pg��Us��U�3�Ǘ��Lmr��.���EG�����,�Yuڮ�����+2�i9�ĮIHU��!�FT��A�p^��_Z�����h��m��u��GG!�ɇ'u��1ɺ�����'ƐY�b�i+�D;D���◲i�S)��X��8mT��o>cEJ�]��^}/UM���.��փ�AW��0��	M�(�L-��-�3nau�i���c���oN��J������^f�(R$v��@�xw�I�pt�wQ��nֺ�	�ŪR�9H��԰%u�(��)��䠔��+��FV��6��#���f�
��m��w��w�E��Ѷ��e]���Q��۝��n�M�#2�AT�Ӓ�[�y!���ՁS�jm>�U%Ӷ�l�T��[<ӻ��˭��7i/omH��S�$�ܴ�j-�dS�GDڌ�,�׷Md�Ւ�X��ٛ���x;d����r1��]�:s��W1J��ks�8��ҺI�8� ;^�W\���H�j�#{zv��3�N�[��&�ͺ!��%n�tY���[T�5L,�ŐfU��`1FHU�]KY�ag]��.qخ&��;�B��f��uc�%�bRڵG8��r��E��y¸P��D��=�̈́ܫ�O��L�X�yG(t�".����{b�UsiNɚ��>ܭ��T2����D[�LJ���@�!��}�����t�׀�hȩ^��TVVZ.�%^��1����l� �Z��-�r�p�YZ�hI�<�����h�q�5� ���Q6���5�4�X�]��z]5,wB3w(D����}뜬ɻ��սG{����vsa9LHᩳ�:T��F��m:�]m:���&�8Z�{�E��� o��<��N�z#ofԬ{]AY华<�n�f<��<�9L���G�,�+n�(�Y0�aoI�W���(��].�J�6=���!N}:voF��F������p���3iJA<鄺]���id��]:Q��L*���:�BgZ4]{���c[��y(q�s/m�Vo��ǒ:�t���|�9�II(���T���H�f�w0�H���3z}:�^g_(����G�,+:Z.T�<�X�s��ﾯ���������z#��K��2\e�	���w	;;D1Rf���5[�5����*m��ʻ2�<˱��8������)�U�}��K�-�C3t�%�W��s��e�os@�2]]u7s!r����T�=D�$�h��d��u�v�f7�j�X�tXb�^��^V�WN�%[{&[��Õ�96����]�v�b���{1u�Xܾ����ʖ
��Tj`u�U���]8d����eض��hc��39�U}�J���b�$�[z0�H:>$���h�%n��V�B���4ou-� ���,o{<-���"pٛ����c�`�(��"��{T=�c;��Pc����;�R��*G.`��բ��	
�܌���A��|ʠ�nq��Ra�+&;�{8:����j�;X�U�a�;��Rq7���-[�71F;����d����u�p���4AH�N�s���q���F6_]�F�k�n�R��]�B��%��1�:�)��mJu���Zti�H/w5�b6��t+%,�i����Ël�73,e7A�é���P�Fm#m����R�n��b΍I/n�6<bVw[fn�Qi�"N��n��)#�^���R^�ݒۺB�$u��}ojbM�s�&�k;Y�2�.��s�T�tIh�{i�z��[��m�ҷ���p���ۗ����I^�dN��o^S�I�2VP�/d	ܧ��B��M�VBHz+S[p�z���}���v��Js5��	cP�(Z�Y�;�2B�U��M�8(���c� ��d2�9Q����hD�2��L�ZT�(��c^����c�i�@Ӈ�(ÝGy��1-,��5�q3�+}h咰�۳r��1h�����(E��v�oq46�b�4�R�%V��Ą ��|�7��3����A0��D@���u�{[Lh 4�����_uCen�w�t.��z�����Rt/�G[|K�&�瀅F˲p�w5��E�U��oL�� Hs����^I�L���v��h7F�Հ��b
��X� �0gbtG%Yϸ�9�
�X8R� �	��'Tێ���z���Q"�&�U�S6s��N����n։�D�D���e�+�N��Gb�]+"��X�=j�12;6�b�Z��A��PU���b�2S|����o��9\��6闦���	g�1Ru��F�I��V�ň{6��*Z�%�X��)��P�G��%�Ǘ�Ch^�y��3M�:���K�SMݫ��l�P����t���#G3F���
��Qº��.���!܄�Aa"�<$CT�%�XڿA�(�V���]�f�'H�2s��.��3����oz�\�*e�X^f�:$���0�Zj1C��\��g�ΩS��eMT�@šG\����� d�0�x9��W�~�
x�P��	V�%јanj��Wі	뵫u�Ő�B��门)�j�Z�-lW��-}�,�M&��'3km�������g�,���eb��%��+��ܠ�1�ŗn9л��#D�gPT�n��)�Ǳ�Ub^]��tH��њ�W[b�f�V��4� V������I��w�[N�gWG�.�JR��:Ѝ����[Ŵ�V_Mf��͗��0��[�e�i�.�pZ��8��MJ��D��՚WGwA:	�u+c|*�f<�n�yKV��8%���]k)՘��
9���h�Ƒv�,�*i/{l��j68���N�Iy�r,)m[��wB�1����+$5p@�����LX�6+���<�{E�h�;N��u���fq�%�,�:W<#'�+�_�/T<]q���U0iгEa�Jo	�c4��*����A�_lJ��'�6i��pU����I�a�grW�.�ۉ-�����iq&�coa�*�Cb���iU��jMb��,�D�+�� W]�-�D��n��m�_I�k:�U���X�(��h�د�spC�n���J�[VÖ����w�۷d<`ݲxv�a`r�"�9T�W�`ǱQԠ��̑V1{�ɩ�u+��c쨨�a<*�G
�w^ژ(#�<�Yup�F����>���Ua	l$q�Ѣ�Iv�/�u��b��n�oq���TI�1��6/lF��@��7O
x4g0�\�	��Zc�@��/h%��R���-r���+XD�;��f9୳t��j����iYw�6��,K��j��n���n���L��cR�o��ENa�����tWm�8�"����l��.u�zg�+���(�=�~W٢
C Pnj��g-/6�����La�,�*��;p)�i��k��JPj曕y[WU`K��Fw�	��ճ�-"��|a̼h���eIy���y�: u��̭�����Ҕ�c/�*V��6���0%��#olYqY��������p��`��{K��o\��uԀvU��}/�,Lt	��.�u6����i����B�1f�\uz�t�2ek��>h[D-��E4�e�InJVa�$	6{��w�{��Nuҕ�mI��5 WF f�M���[3̛�L�8xV>ԑXb�4,44>���ڹ��;�O*���޻�gl0J�D5���'��X�6�ʽ�b��PGD���նC�6q�\p�4�;�-��.K�j�	%�	��FT}�'˛�F�t�ʽb���/-WL�ٚ�,��A���2��%�(Q�5�]eǻl��,���짵,T����6ƶ�'�N�*�{"iF��j�t��˨���Hʾ=��K���͓����u�/D�r�����ڇknG�\͚����;w��m��|+��I�j�9m�뽳¨7+AO�t$ӽPcG�Ue Բna�;Jp���29HTv���q����6";[]o5:cA�0yj��c	6͹#
����^֊3I\����;T��<0³.O��˖�f	�%;Ŷ�\u�L(ܫJ�V���nX�� 1-
^}r��++s�g��y�rk_h���)qu�2���yB����h�+��U�;�i�P.��<t���F���ȻF��̡�>ƷQ&�D�H`��0m��E����h�Yݮ�K�i!�����X\wX�r��]�-.5��d�9賑����ǲ�\�mIgP����_R��N��u�����md���9lֱ,��wG.�5��ssB!P�=,7�f�����X�
�4�u��������}wCx��2e��j������Z�y5�4�8j�3]%���"Z&w
�ur�K%�����$ĳ{t�Rb�ܺ�;%���$�e�gn�Rq�2�Yhvѥ��ݾ��{+iL�Y0Bk�&���L�ץ�en+ǧ�N�dJg]��%��aSYwG��2�íw�����7�H���������u�N�Իݵ��=ld2���2'G.����+]���CC``-����e���Wa���@B���}O��$= ����9�ܶ�Vr���./wۣu���v���\�敁"V@���.�	����2�o��Mۀ敇�ˢӮ��"�M(��l�%��q�1��A����ǥ"���L����]�-	R�R�Y�Nn�5�uML'����cZ�#:�h�`d0:����wҏ�y��p���(�%����Vz�i(���0���*��j�^�E��.Z�*���if(n�o�Lѡ)s�n������%[�]�c�i�v,���[-i��WJR>w#�^V��D��lT�1l�u�A����gZѮSܸ�8�w9me��[O����o/(I��Ժ`�N����w"6�
��{��vv*KX��Ӽ�M��lQu�wJ�r�V�v.v�U�o!]DN�4)��^����i�/u�Fr�e�w����2��+m$^��7qS{I��O�x�V^�!u�h!��|`ݹ�H��I7��]���-M�����#�_DOX���kUh�F.Q\�.�I)NW�'ud��z�ͣ�ۭ�0�RAYI��&E)2��	���7vU�H�zt���h[\$�&�][AI��z֧q��s�8�+��`T��(D��ݲ�����ݶ�3����hͪ����7/�2�ٚa�T*U�ÕN���N�xkh�s���§r]�㥊�L�c$�38L��L}'p,�"h݀��uo^Sײ�2�\weM�x[\�t��A.���ͦ� U����w�a.�3�,4r���S֦���j�U�ȼޒ�uӱ7{�*�1�WkKiӊ�du	��L����I��#�/��f6ƥ��򴨗z8�0��®"�k�P��{����X^l��5Q&)�B�L�4���tGl�L�fv���7a�p�����"��D��o�� �G�qXf��1|]���ac]���+(��qn��[�k5�
5�M;e@�	P5�Vi��z��n��12�eJ2Y�^��R�=�C�uv�B�-�����vr�@�����8L�P���rT��(r�un�V�+ov�=�b�q�NB*c��b]*a���_eu�EQ�R��P�<��4[%䇩d9x�#9�Rf�ʻ������) ���Y�n�dށ�
��#cD�8,MF�ή��l� ;W.PwXqv���p����q�Y�h�u��w F[:��730@��1M�8N�X���|�g�6OW�ֈ��]-җj�����9P�g�;r��G��d�
�uA{�(�q�a�ݔ0'�0v��G)ސ���;�{)�1�H���we1����K`;t�2t��ls=V�ZQ�����a;#�J��QQ�a�f-3E-�λ�F�W`Ԥb�0H���s�$Y$gr�:1�{[ طR����x�F��=�i�/~~U��,)��]��7h�\S��"v)�Ύ�����{��_YB�$�֓&�����6�%�S�o��6����,0����3.�]���[�5�P�oO?����H5��n��ML����O�g�Pni{�f͆S����e���Gh�B��X�.P��W=VE7�˭���d��F%f��^��%
F���ێ�;h��2qzb�����s�kmE̋ɇo���6,.�-۶D���2Iv�fj8f�5�nB��l�fҢ,f6 S�h�w<�X�@�l��f�c �l�m�b��f�v�^��0�!��qɱG�&Ph�=�Q	]�H2Ρ[]�}vn�ew]*����VNNR�RW[��7��3��	X���n�!��t��E�I�,�7z Wr�
5�P�H��^�@��x�Y�P��EѰ-�a� �ւqս}ٸ������a����Pw�թ�)&@k�5��G��
DH��U*�=;w���qK7>��u�;�颯K#C)�3-��\(7��	��yi�n��̺ �:��:��c{t��r��"��r���Z�� Mٸ�4�L��� M���YMErm��,��IP� 	9����)k���a�^�lފ�K��o��� ���]Z�2�n��͖����XokJ��sp
"��F��f��",�řDZ"��:wVt
�V3��nQ�ĵ�X�`�0fA-��T�a`��(�'|�}�XN��u*K\3��t�F�=q���e�i�/*t������Xӂ���8F��d6������T�F���f��ؕ��nN;��`�B��l�)��c�.���ٴ��t2S	�	�N�i+�����jRCw뵖�P��µ8�eu��
��U�Z��W��
�1¯�<��,�hI� ��"eb{�*�x�w��ΪpKB+�R륉h\�VK�.�HbG6� �0��x����c,�G�]n��d��n���r�fu�\��[|�mf���c�8��D�N�&�9�I��	�H�p�qm�oq���t�49���|����U��Iv�Z�L�9xmj16#m;�Y(q���m���aYe�h�u����R���Uu,�p�_e�uζ_GHj��[�ؠ��m�:!�u��ry4V�MG�{�(&y�t
�~[���e��}�k���{лM	�u��f��Qu�^Y̫�%��uB�sx;�
:�tG�"�	�Όuh���i��\�w)�'Q7�P��;�W^6�$h��<��̝o�5e�P%L
���q�����{C,=��<M֓�
gw��o���l����)�NÕy�3�A�N�覫�0�}�a�΍��e>��l��.Ӆ"��9or�֐�g)}�p-Qf��K��:1��+n�sA�}�t�)���7�%8��T3��yN�����tb��K�Yb<8:� �|Ū�)&�����zkU�.`�3���	�Tt���bҹ��n���tjN��ˡ�L���n�� W
��I�e�p� ��qZ���G�Y�;�U������0�]}�[ֳ7���`d��ƶNL[]���13�(�F�y��W'�!�`g'^�p�ծ� C	��##�z�|�(�sQbGh8���@��I�ٚ\��A���evE��YjC�R��cm��o��' �:�ت,sE�s��������ll�ѐ,�	����j�m��GT�-_b�G";;n�e<�Ci���^f�\�����9�mÛ*#�lL�ѕ�o+>(����G\ֹgZ���̡oY꼻��
���)��)�j��7�X#}�Y[V������*Wto�����1�Cn�Q4Wڔ���zgP��[�di�V�'L���Gphͺ���FX��L*�����t9��[z-ʩ-YG/���To����z=�x��DX�����xu�+N�h@����8�[����6�u��(�� ���Z{C�F��;lb9��3�se�4,|� �z���'fq�>�T�i!km&�*N��DuY��zR�n_T�����\7z�q�B�D���
���{�$�E�z7��R	��*wFȽ{j^�c�)0M�=�_Ä����ޮ8ľݳX��հ*�r�W�qzM��W]B���K; Ɏj�/Hu�������Y��b���{ݷ�+���t�	l�>q�w��z_Q��츸�ty|�*���p�S�ؼ4<�$��a�t�G|-yQ�d����q�x�1s"���X%��� �o:����7���9\-��+�!n��;�ڧs��6�Z��b�M�z-Lü~�[��opw��Ւ����j:s8*.#l��ܗ�
N��C�n��ye�}�b(�IQ�6c���cpD%77�]XBd[=��A=���{Ch;�3�&��̜��o�MY�b�<��u\Զw�f��&�&�>�'Nf���6��o��=����w˽D:UX�t�*k��ξ˿�2����X�WFe)6�o9]jQ�om�9w�R�VڼI�˹(ͭ��/��07QT`CEK5R.�N�Y�^�"��c�,�2:e�=����6� �A��-sY㠼7�ؕ+`Wi��_t_Z+yHB ���<�(���Ec�r�\�QXcW*Ԭ���h(�"�U��̌+`ŨԷ-S-�E��
D*TUR,�h�328�ȫL�r���cA��1�R�ŎYr��m����b1eE-H�R6ň��j�Q��Ym�-�lK���&1E�`��--*6�X�V��)Te�1"�V"�R6�r�®2cLm��(b���Z�
�DFT�Re,���,Q���D�!���S)k1��fYf51)��3��ȰP\d�f2b
Q@�Ƥ�J��DR6�U[D���.*�Dc�Z��*TDj-���Ĕb�cTV�jPEC-���ALJ�iKJE�d�P�U)R��B�U�*JZ
����Af[2�1��d���EU+U+�)���:�6`�(t1���e��+���4�H���[�Q}�m�#8��\K#���D&E�)jU48Iywlj���7N��� �RpN����A�S���=�P�
ϔ���L�ooP�ێ�y��ݨC\{xv>y�Vu��U�*���R��t ����N�B�k�5�S���D�1x6i��e�j�Њ�N'"�{Nn�/m!�"b{��wԇYwE뚕�X���DO��������'�i���e��������E��ذ����2"S����~̗Q�ȟv�-E�̸��[d>o���wx���W�LR�Ѵ�A�:�����>��l	�:�Х��b�\�K2�����+u<����i���ڶ��|+��<�R>[a��9����J{WUE�}VR�k���\�h�� ��y'�30e������Der��>���įD�!ప��G�Ν<�žr���U�LS�:�_&;u�.��}�	��4��~ ���W4Ñ�fn���m��_CP+�$]e������~�T�~8����j���f��6%D�I-��Fzǧ`ռ����,e��]����Z3^s���\صSM�0���@$�3���o�u��=�����AgJ���*Yy%)�1%5:\޶�v���״(�^=uK����syP��� �5��p�ۨ��B�y�⯫nf��Ͷ���{\�5dK���_�;�y`��v�N&�Ap����o���q��z��������tO#�W�E�3�W���^�r�8y�^�5��Vy5O������:&אf����n�%;J���)���t9��+Bs�k��:|^�5�沚�?V3�o]$���s�ϫs(jy�Vu@N��9J�䱬q8��=3y�:.C.5�{�&8L�5��Y\2c5n����V6�5q�'���or�[�z.+!������y�q�*��&�UG|꧂ݮ0]r�v���|�m����:�S���=�뮱��A-�����V�&.�����FG�9];�E���\�MBp�s�^N��sÎ�ѷ%u����/qW*3ئ
Mi�Ϸ��z��ՇX�(o-c0G�$c�V'y����$�^W��K8�����2�*.��ot	��.o)��W2���]���^�9X딚'\��:����Wx��YA8�V��\*0)��r���-8�2V{��w�綋���c����x�S�׵��V�R	�����MOQ�Y]CZsӾ+W��֧KZo;w<��W��C9��n��C��3�Ĕ3է.u���9+~��Q��}��/�@F%s�$c),���
���ը�����o�V�o>�A��޽[;����g֑=�3�.#��y��nS}���˨��LR����Wx����V_������Mt�9|�ЋYp�vm��J��p�VA:�r����sI+�����L[o1B�Rz�Ћ��+·�y9/}�D�Ƶ�
���V�\��T+@V��T_	��yx�LR�%=��ڏ=��R;&\*�Ͷ�[�ChÌa��a�sҨ���f{V��|�C���զgT�Z��B��O��Gn��*���s�����V���gg��8�w\9/�|�=zyS!wP��2z�TU:��i��Vsmʻ�^4��*y6������>�X�	�T�!�ۀC9s��y���˵H��6y 4+�w]ܜ>�=[�,�Ըm�E��|�$�osC�z�:��5��v���\{w^���l@���(r�r��U��T'�'����lŰ�ٽ~�"�M�|!�v�E��K���m�a��m��ç����6D�P���[o����z�]��M����Kxs���U��To��Ȥ�ל�;G}X���`��`��ޝ��3XX��GS�}�v[���:QI��Q�2S�c$�Y*�\�p�i�X���.��W5N��d�׃}��UN�Ӫ�N��t3�������J^����g�Z��OP�j��P�Ԟ�ԏ�k�WѮFt�ٺ�1_��B���C6�qϮ,�NJ�>�;�E<���|ڭ=j�h�}��ִ+����Y������ޝ�X&)�ޑ�L��:�<+����M���wΜ]~�l��ڍSMm�o�=M�ܬ��5�%ñY%�H��W��S���b%�hbO���Zǩf�S}�+
�i��쎝5G�s]�p��
��\èPe�:������A;+�j���3(��Y�^*k����j�vud�MG�oJ�/�$$�[����7��Ɵ�� d�;s��M8ӮE���E�]��-�N�l�C+j�wr{�5or���W��z���r�q�
��\�>�/��=4ӂ����ͽ����-��Z.���k���3B;ϫ���2�Ɔ����fp�b|�k�������-~�[��Nelr��b{�k˺�U�[t/N
�Z���Y�t�	����UC�1<�D�[�9�C�Qh�h�4o/�}͹�ۃ/.p]�^O�nyۭ��}U	�7�c#��0V��`��>���zRMO\Y;��2�k��S���gBsY*�R񚄡<#�q��$ ��ӄK��k�����'�pz��>�)�u�=Xkg���:C�]մ^�I#�DD�� E�[�B/f����~�������r1����g{�?"߸��Ed?f�O��w�q��0W^��Yj�1��GnN�%x�����=3͠�5Q�7��Y��h~��N�TzNAX}��\�t�ۆf+,��ś���c]o��:]��2����W���RҠut��Sub��-�F�Z(1K9�*�`�u��{)���J��r�6�);�z�t7#ٜ;u\z�;��o`k�!�bP�&���y[V��NTY�a�uf�a%9Fa�W��/��>w=�ڧ�x��A������V��?����tJK�7���Y��l4��uE�{�1#U���k��qb�TJ*,Ѡc�ݾ���{ƭ��\��\U�qY\�:Ue�&��}�O7u�ns�L��yR��M���N2��<��pbu�����F$��];�/�S&R��d���ِk����<J�`��G]�*A��U�{G��A��[�ѦN���u�9O�u������Q�t4nW��U�uTK���.����Ǔk�T�!4���wj�'t�C/'LR��R� ��D��wzLIʥh�t�5W��]M�u�ܧZ���
io����UO��=�'�L>�`wlן9]�=K�CnpB�\xk���go��j5un��ܲ�>�颌���<�ClÈ�� �s��+s(jy�⳪uvҭ��իG,䘳����^An9y��"и�\7�`��<4��[nv�/�3��Sy|������2��v^���Į�]C���f����#����L[��o$D�;wժ��6���I[I첔0>璚���5����io:�u���rD�gM�>��Sk�"�w�9���[-
O���>��3�c�;_%�Vi�\�bry�n#djUg?�Ѕ����d#�]I�+�x�A���$��ϯ�ʄ�58��^D#���:}�.=����t{ZY;4���!&r7��˼DK�c�QI���-:������⺬��N�7��{��d���ޱ1��N�'�����_������.#�W���.�ZlT�dZ����9��������[��x��*Ej'8$��G��j/Xߢ(f��C���8J_^5�ʣ��A��� ,^M�����U��5�oYy�uY���֢��0�jz1��|�q<��3/�� ��6�r��J̯$&�˨/������W�����AϮ�U4��[N��v�YoGf��
���=+{w��fD�ަ9�Ђ��:��؅�)~����	�U��h}�S�>��.�? ��Zw����XP���;)�y;�� �+��GS�4�9;WH�΃d9[So2�0Ҝ�6h� �C�!(Z�#2�w>{��>�]@��zw:�n #�Kgki�o�����Ej|�^(SI�_'�^t>�ԝ���C��^�ړ�c���z��@Ss��
�1k�^(S�[ƽ)�Zan����4Y~���D.8+�v�-�h�5�hy�ۑ��y��qف�ۤ��ޓ����~�Tݗ���r0���+���~��e�[�%�/D�L-",���Y��m\;t�B�OO1�-��[6�jR��罜�jf�J�un��g��n�.=�sp��'چ��Z�m>R꼓M�0D�g�sk����;�aJ�N;"�{Nn�C؝9΁�*��ή�w�_���]c��W�����:P�+���0�u5����)Ό��T�a���ԇU���!����Ճ֟BQ�(�ݕZ��4�9�7��������l��Qb�
?����?$:�>�]�� y��=ZXN-��Sb��@�Z���EB�+�QYƤ�h����Y��^+��Q����z����k�S��M��˾Kj��<���Ρjr�p�tY�&���m.�jom�\�d�N	ֳ2Y���qf�z�@r#љL�S��{е}<V��X���N������%<���q!;�r�T>��&�m^דu�Z
�{��X���]����~ߴ�^�z�+3��sRo�ǒv=�د^62yqSj55��~�c�jP䷋�J$�x����>�rd	Ѷ��N��HV$��_4�{"g���{ۗ�õ�J��(�T'������j�qԘ�_$-B؎O���hᴒ����7�=9�AަT~���F�D���U.x.���}0u��2C
O�#�S�w�.b����n��k�Nx���.���xW�^w�;�9K�u�����y'������D�-�7�~�*���=�~�]��Z)s�	<삱ד囐�����Rw^ቇ�w���[���~Q�O��=.��o�Z2}��d�A:���)x��fވ�)K|$B��T��"��VNG���8=�^�nA��A�z�='V�3F*9�A;o2��X�JmLI u_]�G	��;I�3��V��q$��p]s4�x�b�í�+�l�]����`M�&h9̩��톙fwK�{D'[�Sx6��9���]˒��K���Lfj/u[��R���NGm����[������XH\}G;_T^-�'K�+�c���پ��I��y��4Fe�}��Ŭت�w��)���w^5ذ�ʄVt(�C�*�Q�_$=�wi���]\��{e�~�� _���U'kE�8��tj9���[�^�Z���,Y��ݠ{m�K�ǎ������B��g�����L\p�(�4��Y��O5[z.��maoseEDeZ���oе�n�+��Oi����Xg2⩓u�o7������)g�O���t���n++�7���q���F��z����=�9܋}��[zk.K���R��j*�1X�E�Gt�U��_u9&��~��5[�=���Q��xܠ5�:���H6��:�K+r�]7'6L�ڮk-��ۄۨ�캁�p2��Y�{������}�zoE�lK�kԭԊ���dV;�f��S����k�Ё����x>ʹu��j���=Y�JXEhy���7�vB:���L�w)�xD��K-��'V���{V�#a��޵���	I�nG�T�2r� Y;Z���>�L�!�U�ݳ<|h��3N��m�*����A��LX��� ��(��A���DD�]:��3V�0(X<;jΌ��[�BV�2����
�l� �i`�;��f*�@�����ʕ\|ͭ�4������
���4`�{ �n�ʈ��ͷE+�Z�7(���xb�{�������*멧S^�^9�`���H+��NbV�`ףj.L�ʆ;���S�� ŋm��5b}�ܐ�OWb:���Lw=���@x���� 7y`4���;l��Yf��$&Vd���;�[Y8�Ք�M�M\Fl̫�3xts���k��ٵɖgc���S����r�<��F���T�Z�i���p�-!��b�룼����9a>Z�]���l��I0����'n���ց��k�U�Տ�+��Jm���3�]Jh���,h�q�P_��vSͪ{����a��/�q�N�x�t�y �k�V12ʹ�_Uˍ����8�,�Ayt;jҩ&e.˃�.{Rʴ�4�A�.���=%C�舯�U�uJ1����66��X)�2�
F�ۚ�1�%W��R|�{���t]���`5}�oOV�Y+nle���)����M�_�0�BN�b���}�l/sV�6*{vRt:�sy �����T4���4U�K��5�E�5a�AP/������V�v���5c+p��3�$ղ��5͌�Q�d����=|'^
,�e�3W��$b�*m3l�ǳ�#���4.�]�pe�
|��Vc��W��Wf�k�Զ6-=]��-g1�a�2z��u�-絭uՠuh��eCA�n��}۫/��GtI�Y��.�.�W\;ܸ�W.#2�ER�+qM��V;��D�L^��.d�S��NT�d�)�zc3�ø��jVf��5Ѕ"��6�1i��]Y�LX(�q8_�}ݳJ7��&Uï����0K �$8�z�䂃���[4��g����N�v2�s�:�l�$�\�;p�(�j��ݵ3��װҧl♲�@t9ch5y�4�f�C�YYM�n�8�eVI(�<��X�^T��:���M��Z/v���d�]dnpy]b�v���u��X+ 7��>�k:;a&���Kٻ\����%>�=�2�{"�kt��J�)k6�e��U��6���b��]�$�t&c�8��^^�lV��f����r���|v�·[��e�g��]L�A�ƇT�J׎c�]_�.���s&���9���jɝ��������>oO%�tg%d0H^�Ð��k�X���I���Vj���V(*ʍl��F����E
�eF�Z���Ҙ�cYRb ���TT��m�b ��ň��T�b�@D�JUnP�mQPS�-������,�
cQ�J��U`T�[)Zĥ��KƊ�11�8�(���b�DX��*(��A�1�X8�B����[\�1Lkkb����(��Ъ�-Z
"�,�mP�Z�Qb+�ZZ�ک*��U-,VFRVUETUk(�-J�"��%A)UYm*TZ�P�������ֱ+)Z�(,�cX�mj-��čV�dA-%�k[e�1U�[iA��+Uh���X�*�iF�E(�"1�
"�`Tc(��1R�J��J2���R"TFJ�`��DX�m��Q@�E��T*��
�.�뻾�U���2���}�u�[���4Ybo��u����i�1�t���ǻFH���]iNk��M�J�u�WW�FD��	���Q�{>��j#��o�f��<��lw�k+Ԣ�'������,f�OV<V�ן�S6.5)�edBj�a�{FGL�I��M�5�Uc]*�x�u���u���+'�Ӧ���э��}ڈ����i{�Ȭ��������s+Q;jx�BgPN���[�/;�ϲ��.�m��7	;#���oMJ����+�Lf��f�<�Y*��t�i��K���v҃p�?c��W�q�,ᑞ�'K�+�ګgp�=/�[W7��2�����#[k����*�N��B8C�tu���^( �ܱ�����z�!?Q=�L�5A��jp�s���sÎ�Q@̳E֬�^�w��͵r��q�.����b��P���5�݃�ܰ�U9].EíQ�%�f��8������Ҭ-^V�58�Z�胓�x�fW�s������Ems�"V���̒���7(X`]`��D5����Ֆ������i��/�g�f�9�x� ��+�s��lK-ڥr���L�4Hs��쇷m��U�n�Q]��R��m��p��%r�qj�r��_m�� ٌI�%e��&���cː������ʭ9+k��i�S��S𨎏b������$H����	�nf��f�k��Լv��]�S�{�;�RjC����.��}��}��o��fRBn�n]x� �K�U��*a�i�������+����/�������M�ܬ*��f��tɥ˛��p�|�=
i���1B�OZ���f��=�������KS���(THP��"\��}k�^(SKx���{`���]�s�q%'�:�����y`���-�o�)��^M}�[����4�iP�N���k�3%��\���x]�A�Z��Bs�|�og�,ӝ�d�sZ۩䃗�Q�4��<��k�^>��5��YB��]�y�� �K�ۅNg\����P�捵�5�mXr��YR����)^|a
��Q��([��ĿS���X!�ۦ��"� �'�X���s4�<Ru�8�;਋\�愓a<�p>U�j�vB�N>(Bv�%�:�NE8:���d�e;�KޚN`���d��6�3&6�B�zwQ�ݽ@�v8�|�Sm�*)�����
̓�=�&�����ߩ��4���*{^st��D�bs/�][�6��#ù�{�y��*��U����漝(�N
�)��e(;Y���։K�vb��S]gB��V�����k��{wR�8�h�;�Z.��ZZ�o��x>��M)��j�2W�ϭ��V��Tv<f�7<����=/݊6��6��v{ɿ��x%jU����=�6�b&��>��G��z���{a�r��oi����>��[��yF}�\��b���ַ:�u�F{GPq��ˌ��c1�O&����]�����y�����;ݧ��]��i�[��P96�w����UrAF$��w���-��gh�WBܕ��<��YNs�ða�#��2=�p�0�	�^�q'YX�m'8�>?s$N0�|î�'Xy���{�
�jb��ٿ5;[s�P�p���ѽ$DF�i���w�q��=���I�:��-��Y>Aa�:��8�r�$�'�����maěe`h�C��d�>zw��&L���Y�"
��z�t-�w�\���h�.����n!c�Y����YתQM�l��sd�J�~���]��ETn�v�:E�7����e=&�V��^���������:8Y�ni�w+���D�0��1���'��__E�^�2�.r��z�~�껪�����~a1���Rm�	���a8�2z���ē�z��$�d=-:�d�-!�>d�Q�m��hm<d�{}����/�V⯮��u�~�1�vz>*CL�2q����P��p��=�|��l�a�js�	�����^N!�߽�LABy�q
ɴZ|��GƐ_!�_�vgEUVg�)ҫ�{����;�k$�y=��'ud=���'i�́�P���oi'��쓩�'�=O����g�9��$��^I�@ٌS�����u��W׫���#�=Rw(I�N'��O��k$�h����!᯲q�>v�Fs i�ߣ̝d�����I����~9�������cŽ	W!�� ����z�LJ�y�ԕ&�Y<�N2|ɷ���	����4�l=C�+�CZ�'LN��}�?$�I���2q��5<v�[��x;�ڽ��-ӽ�����Yٯ�&���Ӿ~���u�/���>�IY7���e'>d�����i�����N0�~����'�z~�q�`�=\3�ۣUs��O���ئ~��=���Xzɴ��AC��Ag����d��xz�:��s5��d����d����&�z�5�	�S���O`�1(����W�yE����#���wzͲLeC���PY&'9N�q����&�i�C}�
O�<���XLd�}גc�I������[ lG�h���/����}��t̨�ފ�X4�2xÉ;�I�'P_u�$�C����LOk�m*ӝɤ�I�*�܁�O�=���i& k����a<�	�g��|e����<:4���R�����I����'��mq	�~f2u�RoVO��/��	?!�>�O&��>ì�J���ri'>��]�@��!�l��PNM��YVc���������q��0Q�hTku�����l�3��Hs,>�z���,ٽ�^NS�\"�-�;���폒��u�K4
�K��
(� ΖY��{���3qq��N���.=�tG)�Jܼ���4U(Z�6a׉O�����/O��^0�`S��q��=�E'�l���,�$�Vz�Rq	�n��,��4�Y:��^�M���̜OY&����{�p�z�4��[��]����P��d��'}� i��=氓L��a>q'�4��Bi<d�{2�2M2���8��2y�Y8���&�q'YSp�0<�{��w�+4,��������Wv+�����a�N�a?{�Y:��l�v���i���LyCl��0���d?'��OL�2O��{<��I��!�{�z H[ͯ�3�����'�-�x�Ԟ2�a��Ad��;N�I:�|̝I�L'�9i4���s�'XN����I�:��-�Y>a�=��x��&${���T�y}��Wط�'��o#�'�I�ܡ�O��<�Iԝd�~�2Ad�y�_�LI��ru&�0����I��Oӻא�I��9�|�u!�O�{�D�\cV�������nk������C�'�)�'�La��I�S(u�o�AC��d�>5̐Y8��y�;I1��9�R|�&�z��N1c޿�עG��=�%������}�_8����y�b
�����,<-�$�(�m'SS���'�>d�������'i���������'�#޺�c�1�`�P��!�T�xv����|���O��O�~�Y&��ߵ�1	�u
ɴ���q'�6�p��d�z�mI8��|�N�K�`u&���==S��� M5�|v�,K�ۿ~��=I�u�l�������2};��d�C�w^I�XM�XVM�dє$��~SN2|���������B<F�zԏ�_�3b�ڞ�������/O��4�auOXm�l�1�i? s�
�����d��?x	Ԝ�䘕$�}x²|�@�,�d���1~������t)���Q62��/7��l�cQ�ܱ��;���D�Z5�3�(��s��Z�n�H�g���36��粍)/"4d�����kVˤ��޺��d�S�Dx>��܉���H�p\!�{��߸x*��q<w݇�j�z�p���Y�{ܝ��~�#�`?���J�'�?j��bV�8ì�g,ěAHvs��i��AI����'�'R~�k�1+	���,�1�x�E�]y���͸�ޑ�`�h�"<�6·�z�$�����'�z~�u�bVo�8��1�,�N �>�;�P�&���o�AI���<a1����A?�_�o7�I�7����ޑb=�GY� xe�XI��~(N2yM'Y=I���3�N��ky��+w�:��1?r�d�VC����h�=(��"�ˎ5��M��= D�'��גLd���+���vE'�L%��䟞�����a<��O:��?�|���AטI�a���P_G�D|^JS;?:��}��bM�N�]}��VC��?0��N�vw��M�zo�߲Ld����8�x��Ȥ��'���$�T��Xq���i�$�
�����������[���C�9�_��"x���3ē�7�:�Ĭ���p�'Y>~I�,̚I����O�=���N���!�|��{�q�i*y�Rxc��)�~�1�d(���ob�nw�|DG|����8�̝J�u��N���Ì����u�o�|�u�6����:��&���ׄ�`{9C�Y<I������{�׫>������L�SI9S�N0��gO�6��a��d�V��&�u��Y��'ue���8ü�:��L'������O��I��>yͯzG��z���&g[�|w!�G#��O�ٔ��<d�{2��|��:��m��Ì�J���l:����H,�C�y��Y'X~��:�oO�~r{G�^RꄮS���Vb�G�{��G}�c���Rm���6�̝OL�0�I���g�&�rÌ�J���2m����5̐Y8���g��L�q�E�_f#�6�/1�"��|R�HIhS��j��W�kI��^��kiuP�A�N��R5*�R#��@��R�!��^.�¨'B�(^杘:v� ֻ��(��j�\ݛ)�膯�<����{��SF�����4�F-h	J��P@�Ր����f�D��=舀^ci�u��{��>t�|�'Y�'�����I�{Ͻ�LABy�:�I��h|���I��O'�6�N2��M��b��#�0Dl/.����w���t�]��>`xó�g$����'S���x���O��'�漆0�C�y�b
Svq
ɴ���>d�Q�m'Se�B'����MK˞���3�.!�{�I߲m���z���L0�.޲~a����u=d�'�����C�O{��I8�;�$�&�ޤ��J��"�p���O����S�u��7�%\|I�O�٫[$�<���WL���ɶ|��z�����p�4�����'�,�w�	�>d�;��a:��9ʏH��N����O��ޥ��J��VJ��O�6���XO�>O'��I6���I_���a��>垰�$��a�'R��ACi4�ˇ��{����:� �u.���,��[��8i�i'~�xLea7�"ɷ�
��I��><�`u<?P��I�=?X�����?k8�c*M���:�x���ŏy��#��}��eJ>������ ��&���}�2s���$�N_�&{d�ټ�d��̰�i?:OǖC���=z���i��1��?i�z=� ���DEZ���d�˗b�~���i�O�Rݞ��&�����̞k����c'�漒��:�9H������u����'��Rq��=����|=G������U/����Wg|�T��8ϒx����~C���Aa>g�>�Ԝed=�ܚI�O���s��>d����l�=���8�x���)?:`yl8�i�O���.�}��w�������m��'��c'�,��~C�8��5�~C�=�s����~��:��������N�|��G��4��Oy�y��㫪<����C-�׾_ۡW����/�g�яn�:{wyԩV(~9�Zi<�b�w2�}�����*ژ-�A�j�,ayV���ǝU�3���sd(P/��$�TΫܞ���5�:�)���;���:�	�e9�3�XR��V�g�fͺ���(q�`�C�X�\������3�9��}�����&��e��eOXm�M{�:���Hq��S���a����I�}�:��XNk�u���~c����D!�Y�긥�q����J7����N0;��O�d�����CI�&��e�a6�O=��
I��:��O�I�N%OMs!8ì=9�v�:���ì�Մ����Nӗ���ݝ��i�Ui��Cޱ�������D!�_��ؓ�m�Ҳm����!�x���ˌ��:���Aa6�{aĝe`~a��d�T����'f��������ʼݶ�勯��#G����fc�y<a?w�I��Oӻ�8�q��y&0�C�l>J��-!�>I�ze�I�La��I�FXq&�X��	_\��͵��y�M�D!�h��!�}�
����=�����wyXN'̞���O�ϼ�1���:�d�-!�>d�zad�a�}���d�F��{u%w7�����}}d����^`m���t���@���=��6��L�>I�O�=M�;��OY=�޼&0�Cӿ{䘂���8�d�@��c>w?V��|�MT}#�=�'L,��3��5�m<��|��YK�2q&����d0:���x�I>@���'S�O�z����M�Ԝ�� =�|":�o'j�)���
��~�P���J���<��>d�{���'����q4{a�J����8�ԟ;a��d0���N�z����8ŏ{�@��R����W��7k��CI:k���8���גbT�oT�ed�e'Y>d����'��5��=�ԕ�!���8�bu�����{��6E����U����NgD�����w_d<d�=;�	�>d�{����59��LJ�|�%d߶���'̝|q	��_�z���i%~���+kh�}�wn�uV�S���H��g[�`Ų,��<��~u�=�9\k\.nRa]a=��G�И�uM�jN9����:t��ǐ�(��z��2{b��&��Z���enfE��^Y..	�fR3��P}�]�]��|��_^�� �@��-×��$�/�y��>y�?g���1+��m'XOپ��'X��AC��Ag����d��xz�:���k�1��;�o$Y7���2���I��~���걨�]׽�n��8�G��h�}�}��'P�k��$�T<7�Ad���:�����I�*����2y������Ow�y&:d����I���������`�͚�/��V��"#{�H��l�g��6�����I�'_Mo	4�P����$����&ҡ9�?$�M2����4��'�w^m$��멫�^��}3]��s�9]4�_��=�jȤ���l:�|�g�x��M�L�:����!�']yI=C�}�:�2M3z�Y6�	�,��l��&y����3��1�#�j�bk�?D1�p����y�����m����dR~v��{�u�i+=C�8����2q����Hu��/��m'�~d�z�4����G[����nW�p}�ە�H��!����ì�d�Ԛ��L�$��5��`}��'�$�&���I�'Sܳ��L��Ad�����Ad��&�q'YS�u�
�����Kb~V�u�=B=C���L$���ә�Y6�����N���&�{�ui>s^i��6�Ɍ=CS,����S'�u=�Y'����@f��tN�g>��,�XD1�p�=�$�'�8ʞ��H,�a���]��a�gRq��l��@�M?2~��I��{�I�:�Դ>ed������x��s;���:��ϻ�כE{�"��"I��>d�V��M��'5C�d���{�:��bM�Τ���ې6�O̝��2M��w�$ĝH?k�wz��|��no�k�����;>B�~Aa�`z��:�̦0�I��ya��m�u�o���6��hs\���<=�|�$�OC�aԟ;I����$�x��[޳���5(�t�[���T�4Y��B�k�r�t#S`�`�.�o?�W�m�#=�g,d�r�d��:�G7+$AԒ�xf�d�sY�vυ��w셖�$K9��"R+l���}]W�K/�LvX<�=鄹le�[:�aTIul�Jҟ��諭��-.���f����d�3�5�|& �<;fЬ�A`�q'�:�$�I�߶ON3ٔ>d�������I�hh�a tz-�(1�yfb��Q�������zO��ɦ=�~�N'�����u{��& �<7g��J��P8��g�XN2u<��mI8�=��&�2��G�=��5}�mٛ�s'r�[��a4~�̞$����������uY=�����N!�;�$Ĭ'����iY<2�ğ2o�c	�O�G�����h|m%x�o7�F�T�C�6�kT�I4�fw�:�8v��ğ�;�d����Hu�=;��a:��ܓ����VO��哏�����2Υ�e�cJ�7��t�Gޏ&M3���i'���W䞰���I�Xkt��M�=��N �=9܂��4��v�R~I�w��ԓ�9d���{�G�MH����`�7ںn�ޏ��{�)�Y>d�O��@�>��]$�C���u��=���$Ĭ<�� �L|��N��
C��P�'�>�"=�=�`���>�Fb�$��s�k�h�1��_k�1�I���"����Xu����'�(N2&���$��4�:���u��
�����$��?s�_A�yFsw�G�aK]�rf$�=W�)����V��K�'ƨo
�C�i1է{ޫ�k��#��IO(��<L��H��{��ckȡ����V�f����5��e��ֺUr�s6�T9u�ɡ^���R�ۄ�k�z]E��AX��F��i�QO1l
���^��1���X�N�D^��1)J��$��À����V�+��֘���[����`�SCo��jI���xf�O�?KPW�i��[4_L8X$�F��xV>��,�t���o�J�ܵ���U�L 
�s&��T�}���.��|�4��я2F��tD�Zܚ�r��� ����*7G.w�ƕ��sK|LH��:�m�';��NF.{M2]�[�b�hQ���%�}3n���� �w�ef���?�fScU=��/c��.�LYg��I�ژ�N�m�0�.��*��d/���B`\跩��;��v53�ylt�9
;���`w3��<o����kJ&�/4.��TH���{��An\�r���y,A��k�=�~0�_�B�W!�뵣X�rW`.������3�ݨ��.ָ��X`Z�}�_:�VW=�{�N/��ô���iz�G���V������tl�K5Ѐ cW\��9@���fM;}���5�;a��u#�I�p〵*"i��ɮ<�3n��h#DՙNm�äoh���˙u�G�n[B	�`ש�U��c��X�Q���ǭ!x�e��o(���:(W�:�֌�ر��9�IK ��ԗ|�F1j�U�Ef��@��Y�4�p�J��px���f���`��Z�Ѐx�Y�Ҕ,J�:���L:�Ց��}4���c������;�jP�l���:v�
}�]�D䬼{5Ʀ'h��[A�<p�ۖ$��)����Ι�V �غ�(�Qdwt{-�ܛi�`��Y6Q���&���ݼ�����Jֆ���,|,�Y��7n�	VU�E��Z�%��*
������D��7za� ���"z3�d:w#Vj�)�6�f�eb|)��*��\K1�%
��A�� գ��/JZ�s&AN��;s�K��9�Q5w���Q��d�jPz�U�Yꕊ���\��<��X�����]�-�s�4�s�rʄ���c���z)�:�uhWC������aY��������%	�@/A�؞�v�*Lmč�V�所v07teZ�烐7[��ga�[r�9y��)�)�R���EV;�Yrf�"��k�v��$]C�ϲ�i�T�c����xr�ơ�Fo�ͅ���:�O���͑��LV.�p��(=l�5�7]����6����ZHW�E�&���eK�;H��ɰ�W�E�2���a=���b��峕E(��� �"��\p��iWu�uݖ�L�+�B�'u����`:c�+C����o�y"�N:ֺ]]��:iڍ�a��n͚&�	m�i���k=\��؋y�˺�@E�	�f����+�!������Ϳ����Iԕnޤ�A�ųtoX�F�Gqm7�����Hbh�59�O֝HoZ���B���9������]�E�)��U�+�c�x�  < m��Qb*�h"�*�
���*��U"�����Q��V���Y�KZ�,P��ʬP�JŪ*�(�[aPm��TZ�dm�����kU���RQeh��PXU����%J�ATU��YRڱH�m��,
�Ym+*�XUB�[e�-�Udh�(�*�Jŕ�m���m�*�QQ
�B����H��Y[EZ�d�m�VEiem+QU�m�Z�j�DV,���!X6ԢQ�E�*�"5%A�F
�j���R��(�B��ZJ�U*AE��ʂV֥�h�b²��-* �*�Vb%�H��XV�PmЬF)Y-��UKjԋPZԕUZZX��X��-�VV��I*��*TQej���(ZU++m�kEJ�J�FԵ��Q�P�~$AD/�ЭU;�|/6Ȓ�g���݂��Ӯ��it��+h9.�7b�ls��Z���U����/�%�^�B�;��UU}_}�o�7!�hU+�dU���Tt�W��&���oҳ*k5-{����ɳW����]�)�� �ͩ|������M����ʧ�*S�k�e��4Ň�vz��U.:b�	�k/)���/�)��]��MiD�^p��;����������ښ��Ǣ;���xʃ�WR��礑�����<�ͅ�l��1��{��U�d��tX�~�o�Y���d%*~#��g[E��܍z[W.�yYk$ÎC�[�c�lTئ8P��姍�[wj���A��³9N����}T;����a2�XJG��y"����!���L�VOs�u��+�{
���{��r�a�Û{�QF������R
Ƚ2��K���uE����7���[=L�/��d��&m�D��c+ԁ�~�,�mJ�g�Bx]�O����.osQ��P�V��=��<�<ՋC.6���a�VŹ�6p�B��o`��sM�������˺�8Թݭ,Goh�P`����[R��(��p�VKh���۪�����g����l��e��͝Q-�x�Xs���]r�v~������8�.O�ت�����/�'t�6.�ȉWR�d�z#�EP�]��z{� ���\�⼝��7�5��݀���L!�sv0�OԖm�{eC�<u��j�6��vk�����o4�oҊ1W�O�M>|�����VK��j2idju��m�tRͨ��U���_�m�_%:�V�7j_�`�nk�E�c�+�GJ���/co���Gd�چ�c9˵���:��ݸw����/��(1:�U�C|���9��SN_.��m���:5��D�S}�+
�ò�J�uԨ�L_$.�lt�}��r+d�����WB͸��E�hؘU�����9�L�,iK9�V���x��.�Q���m=��t=�[����N��2��3O���rO��ryӵ���dk�^��Խ���No�	ソ��GY���!p���R���3�TS�=Ri��SPZ̓�|2�ta�8:=Y����ƅk�r�n#m��Q��5�io͗4�ڮ�ạ��&���Лf�5X%�7�.m�$df�j�������J͗�1Ҵ��*C ��/9H�[�&���v���D{�'��T���D��u�W5�(rY�V:��f�[V�W
�feN���)r��{Kc��{�am0�Ԭ��H2�߷����8ݺ�v��dGn�v)Pm78Z���Y>ȳ����,I@nx���>juI;�Oe�q9��ӛ�tZ�����ݦG�����H��^��Δ6\Go>���'J*��^�)�;�G��G\�׃*gUD5����~q��X}Tut�'!L[2�sҶx�w�q��5�jv��d��
��	>qۇ��g��.�Y��9����k~��z^��\��'�*a���ٱ	����4g�X��z��?*��+P��c�ii�N�kCa�(>���{=�ɳ�t7j}�oе�i��Gۿg+o�}[2V��ޣ�C�����MF����	��x���y�p��Fޚ˃�����u�q�T��eݼՍC/C��O,b��W$4��;7�A&	�F��v:/i�K�;@���XT;�|����P�lBA�Z��,�ڷ� ሠx�EX�i���ҕ��e79��uo5RT/�Q�\�]_l�乻��E:��������c�*yxg83��Fc�r���p�{��o���\&�ʢu�ލ�wH"�n���6_h�m��y�h5}Gf�m�v\h�f������\��T+L�ꈞ�E�E�Yy���x�8ץ�Ϣȕ��^�w�:i&�ż�F߃&j�y�=���\~�*d(J�����5���>p��3v��p��00}�@!=Qx�T2B�w�!��.S�P$����������ک�:�q��l#ݕ�nf�Yv@���xd%S�+XǽA�����ҭ�V���W�<"y�V���02k6���+M<��s�1��^x�jW���RoY�x��1�m���Nb�޼ݼ׭^L�r��]f׭���F�6�9QP�vEy8Ʉ9&�B��Ou�ݤ:����K�˞sU���T^2'�A�rj�z��)C�]�q�b��, z�n��w��Z.._'B���Ty\��]�k�]��7�Y���h4�� ��X_+���"�'�@v�[���9�_1k�lʱ�.+�+Y�Hm�H�&t���<�̤�'�)B���f��S�tW{�ܓ�/���W�WԴ���=��[���v�� ��.ʡ�*���{T�Ձ�etT�}盨h�9�\F�;�R=�$6G�QB����C�SA8���N8<_	��=Ld�e-��/{Ťg�~��C6�q��4��]��n��v�U�t>\�+�t���Ыm��f��'�Q�����㻙��+�&]�4���Py�/�g��*y6u1�z����E�$zI��U��[k��z�ʢ���'S�
��B���k���Y!�A�6�ѓ��8�Zw�a#���gh<���������o���
b)=p��su�u7�궺�I�A� 3��'�rw�u;5=�;G�W����&����:�Ӟ�jP+��q�����0����[F9�����t�!�^��p��^�w]���4b"#G�[�z��#Q�m\���X[�1�h���ߟ�ԩ`��e�"�,u��-3����"�^b�KZ
i�e�c�|�|(ԯc�/]x�Ys+�x֚'6 �J�u'E��n��{�꽞52�UY~Ѫ��aCK��w�*C(2e�:K���*����E��PU��_�#�Ԩ<�z6���j��ҍ�ޏG�ﯚN^���K�J�D�\���v�jݺ��7
�yee�8��^�ќa��o�����}.'v�y�9��aV�2�a�[���&�!{�`��K�\%\�.1�0�y:]�;�U<1K��=�r��)�(�O'F�NH��SȂ�֚�Mm{;}�<�k`�t��;�U'���?uj�vCA�촵.�2z^�(n��0�Ӵp۸�����"UԺX���f��d�5���gJ�}����i�jv�s���zZ�oaE��>�|Q5�jڵܺ�Tn���~�sմY��~��z^��W�<V��X���5p?HNe�<��]:I�)?�z����SY.*/�ʵZ�m�hT[ow")f�dSy�T������?x�3��&3k�ݡ�~ג��_b�<�Jz"	���o�C'�����CY�k�dr[�棈:�\&�N�|�ĝ�%���T���w��B���]u`� weI����[I��Vp���)u�e��y�+�k�nL	��x�$:�"��\���:�s�r�{�n<B�Ʒ�!n�f_��,�+�6�����L%�;y-UY�c̎�K� �VlQH�=��)Y��X�	T��nJ��������O7�џ4g`��D/�3��]���[�vJ�u�J��L919���Y��tj��&�=�ل�;�E�zk�Av]@�����9�+�6ĕ<��o��[���W/C�T���s�J�;�~���=���Eͦ���Η���[�P��\�+�I�k�o��{�������P���X\j�ڔ,�Cl��L�Pc��pS�ה9,��|�qۭ��"M�!����y���o8����S|���r���mes���h��wQ���9��)T��o4��&���l\:{NnBxG1��1��ލ�6�]U���I�.3-+VZq9��j^#�N��Ek��ֻ�U�#aӫyܖ]�F�|���do';��EBp�+�d�;�~G����LP}Y,`���s|�+����Jj���2U{5�ڠ�&��Ţ�9��0/���?�O��W7����<7��g�<��[|pܐ��)'�:j	a�7;n>Y�ߪ�W咲M���0�Aҙ*}�	�Cu�9O7NSrX�ܔ0�j8C��ϵV]�Ӳ}�Ji�E�w�1��X�#��Y�׫3���X2CouO�_}�W��r-���ZpV}�s�����t�ʍ��]��|)<Z8U������y7\5m���A�Zj5�4�P����=�'�{u�y��b�mɯ�]�/�KH�'��^��6'b�>���Σ��
��1|zl�}ǂ{�{�&�S������&�{�ߟ!���І�핅w;��ŝ���$������73��ƚ.^�}��������w��;%-�5�c��O�~
�)�D�c/���|�k.�͸M�.�ɡg+1�
&�k��u�Q��QL�E���b����
b)=5�+|;6���V�~��HߜR=&Z!{�{m۩�Y=<V@\�.��gX���Si�j{��q��V�3�d?,\�Yq{hS�Z�m��r�tU�U�{G@ړ���\Kj�����ol�r& ��	�p\��,����lgEr���(�S>��)4n��:lu^zP��,U=/-�
�n�i��@񹇋w/krGڶEW1��٠iXV�:0�(Ay|Wt��u�Rm,h�gg��l��fp7����|��)պrHB���Z|)Nbn�J�����W�UUq����zV��{q�y�:���mZ�L�,����z右���bDY�^��O���!ƺ�GO���pU�~V_��Ȥ��9�u��A�%�����X�-��n�鋬U��^"'y�~TRq��Ǜ��$��:�'GI� E�Ol�K�-�n�Ԟn_���g*�*Q[4>[}hݻw7ku�tle�f�_w-4O2W�P�6��Zkw�CX��1�(���t{���ʋP)�k�Z��K�=S=Љ��{	��`R���%!*Ek�X�X�Y>5����jX����Su��C�Sӆ��]Fq���-u�}���&��L59v��5Fs]�d�� zw��!t~F{�Jqߪ��P/�tC���Gz��n�&��c�����ZcI}84OU�\I�\���$k8�U��%��܍�zx��@��U�Ȅ]-9�6{NE�\9���Ѵ�Y�9C�C� �"��U��\�])�/إ�n1�Q
_\<�2�*�<bM�% �e�O:7B��b��d�%Wj��y�.�}.^N�.+se���)�Ӻqu�,U��j�~�y䱶����ax� ���x��]oBE^��/T�哮<Վ����J�Ne�3bZ�C6ʎVc�em���,��B�S��Y������ޤ���'j��?��C����5B�F�M1���mJ&�Ku�E�ڶv�\�Ir��;]����A�N���|%oKY22A��pJ�H�Y]T%��Q'c:w��ҀC�:�����x��Rm}}=l�Q�{ɉCne��k����(8T1�J%�h�~���wV�ٌ;;g�|V��:���W"✱7�6����b���`T'%s24Ud���N���Ӟ\XC��Hoc1q�G�ӷ��g4�K�Ga�EB��P��X�s\������S8��s����1��MO��5�9+)��S��G`T�H'�)�%�Km��`���7~�q�i�f����G���U����C
���0��ē��MV�<�>vgE*��ؗ��uT!�S�T;��B㵾�A����.0�����E��k(c��d��Q%�_3Bâ�'a<�E٠���#zjh�1e3��a*��S)v{ț�Ȟ��C�x-�W��ܪ��bv�[6�|��:�\3�0;�f���F�ab�f�"�i9zDO�NC*�#ÄX&>����U��wU��ok�� �0(��ȸ��ȶ=�Ρ L<��A+,��2�.��Z���qQ&a]{}��$�(ˢɮ�?��nv�E,ǀp��[a�Gu��N���ZA�7U��HG�d���H�r�ݏI�9�ΓA��^�-��,`��t͞�2���s�j�
��=w"g��z{��*����ݩk �@4s�V��:9�5��Nui��v����.�<� ����<�`�N��4�6�U){todKpp�C�C�s(�G��5�\�]}���4�P�ѭ��i�$*��a͹�k��e)�m��֠^�0�C�ֵ>�y��I-+ՙ���r�@�*1zvn�yzn��g
b>�m��`�gt��WJWù[K�Ѓ���p۶�Y�ڵ�%���POP���Z�7���W��!��`�����S8�ن�L��/�:Ȧ���*�h��Y��K�3웱z��[nuF�X;�@���E�rC����muu�2m�M��гo[�gN2���Dp�#��S�^`N��qmmay!��$�ut��%t6��,\���Û���;ztf\t�&��Ѧf�دQ�#����X^��^��o+�n���v����$�Xv�6��%�.�ՏlFFm��L�n�������w�L89h�mϙá�wʗM*�7e�VA�w��u+�#(r����ר7LXM���5&�w���L��7��`��ob��9j�Yn�CnY̛o������y˧Y�/53Z�7�6w�9����5���j^�!��;(�sU�2�,[�3nC�9K����f� �\��ũ���Q_D��kr�a�͊�&�Z'Q��)p=��#��e;�-��B�.�4l�i�W�F�vӭ���<����������#]&�֕�U�]���� g�l���� a��-���RИ�Y����k�R��5�����o�uu�9�ja��?���M�@�Y\F�' IT&�ZM�M��SQA�c�yj����sj���}���������(Gcj�k����׼�##�����#����I=�F�ӷ´\9�ȫ`$���[s�:N�:q���pB�D�����sv�>�j#y��⊜=`W��e���:�cc��	Ց֝U+�d]
C�m;�	��2��bw*I��0e��޽�t��頠B��[����JիlM"v���yf�p�A׮��\]#�O%�@I�ue��J��&K������H>C�v������X�nmi;h3-�����]6 ���n�+�K�c�9J�Ԭá��jn�+���]�������d e8Doz�V`!ծ��������F��,N"�ӫ6�7k�պ��gB+FD8�L�$rŉO�8t�/i��	]y�n��3�teW���s�ep��PEZ�jJ�������#R�Fұkmb5R��E�������cF��
�P�҈�ZV��DF�Z[J�Rm�Z�-H��Z��؈�+*Ԩ%��Q-��`��1���[R�+mIF��T"�Khյ�UQ�c����Z"҅ER��)m��iU"�	XV��Z�Z�PU�R��`�
"(�TVV*J�h�QH5���[DJ��6���2V���h���"�!RVDEb�ѭR1Z�UQIPZ1H��J��R0m�
0PYJ�amYc"µR�E�PQ�XV,�J�B���QEX�D�P�,PP����T*TQ��+*Զ��V�RX��X,P-���QQ�XR�����UQiR[KJJ�X�������E���+J�YFjV@m��EYJ�k*R,--eP�%J$��(�-�+B�KaTeFʤE�eA2(��(�,��*DH�KPm!X�jT�޳ߴf���O�"V��6Լ��`��I��dv�Z +5i[t#��+9�L��g�ƣ!7���a�aǡ�*>�����ji���6/vf��޽�A���p5��m.�� ��P0xV��r� ���F+,�M�ԥ�Z�wRi��D3�mK{4�á��`wΨF�B�h�����Tb�����$�C�izs��6�Tp���bu]��g��k�%cn�w
���A,��XWe��ت���ZNד�nP�^�OoH_E���v|�iՀ5��/11�B��Wc#��ӽysN�lԦ��1L�L�Q���������z�i�t���=�YBP����wf�Д)�v���3w_��8t�o�m�4��t���a���#���6�_����\mF�4W�f55��iI�;�כ��"�L��Cea��!K�G��hU�Y;$ZZ���*���i:�m֔o������(:�T��Y��S��@cC���"n�w)�:TA��P�+w�G��8>���yBE^ײ%���>����亅�F<�j@����<�V��ʓa���G��wt�}2�j�`C���?����[�T\�X�_I�^��^�5Z�<-�������o�o7&
�Ï*A3���C*d<3�N�xN�ͽ�D�����\�]
�K;�ע=��tC�"���0�5�چ�jNR�������;}D�fï��B�c���T.4hE�Jq�g`:&#�������]7�r]�R������<���sJJC~��Vpc,V�j鍸u�"}�OQ^���\w4JE�V�\�Z��w�*��(H�i���N&��0�l:�兑\+Y�G�y���Ľ�<����n�,*�#�Y�Oם)��^�wjd#��	�*!����NT�hz������l۽�"�����,:���v���I\�bu:���GI��#�Sް���owO�<�k1������Nj���ya�������aꓬ�C�]wt_�j�׷Q�K�w�n��=N�o�=짊����.b�^Tƻ�x/�3��}KE��7����/�4_���@צ+o�u+~���9fgs���x�R���H넩 �ŻǪL��\����Luêvtd"��x�1����5��㳍X����w�4��QXFb��]�ɽ���7&6z�e��!3J����i��7��n��ܬ��o9�Eb7�o��[��&����c�WPŀ2,�H�!����A��B�v,=�p�;�F+����5�lI��A[/�aA��x{�VW<v�T�}%�+;͑���at��]O���`�c�B�!�T��1m�^�۞*�z�:�S��0�������J,ΰ!ȍ�����Dcz�)����Q��q���4�6�R�˷�Co
����"<�j���4m����蝚rg���T�L�H�S�DZ}�7��W��͏v��m>izys����v���O@�{K�3�]J��eY�(Ww�m��Z��A������	K�����,����z9�R�m����P���	{WXa����R�Qu�'εxSj��;��Z��T�/G���g����a�s»�p ��2G) 	�Cz���f�8fWu��6s����v�	�{��CR�$]h�q�U���Y�ȅ�ŋ�Yų��1�O�]@�	P8�o�����
K�9�W<vtC�J�Q�����Qȴ��YĖ'r�h �q�W�{T+�A^I.5I	g�z�Y��\���3}M*.<}`�W������[B��s�vf]��h�Gܻ-���^�A�7*�C��A�\�4�ހ,W�������$��^�D��4>�2r��V��s�(��R���SZbQ�9E��\�9e]h���]�x�J�樈t{	� C�;ۉ	hۊ���5����1>���k��]��	�h�;]ֵ;5�!�5��cct�����T�Zyg1a �OKS��V�3�D�/0ۙg���-{]3�޾���n�2�v:��D=�od�'n��\Ŵ�"2y�.�����!vA��׽�b�it�{��Twc�}_}_}�W7��m�����Qq~˨�o������&����醄�
4;sm���v4�aWY|��ü�,|ѻ��,�ӡ��S�xtB����F���hL�i�Ct���òӢB��
�Ws���X��B`��2p;1j�_���{�Y���mh鯜��.���a��G�T-�5ʗN�=W3Z2��d�(V�P�c=���
�üH�_JD�b�O-�O�2��x�91[ݶ��c���W�}+ُ�_�0�"4�$�k������Xy&� ]��酗�C1Z�JEt�\nThb�K�C	�ǝ�}ɔx��i(G�"y>lO�ewT�.f_.�Ԥ;�*����� ��|�EӘ�)��=���yu������
�����qtk+5󝮯LpC��q=O��XWU�W"✱7�wg�a�L�S�	s�}ӂ�,���	j�K�y |G}P����J>9�>}82�S9�!�1A�ti^��oWV�)���G,�eSk��j{�7��c�����>t�XF�vG>~������2������C������&�'��|:wfF���S�۽y��]�Z������1����d[� ��I -�B�9X�= �D��)]�N�2̑DoU���أ��6C�F�j�$�ǚ�8�+oU�pL��٨��pr��}��6���O��F��2���)N�8�D�p:N.Z<��ܵ0�hi��R�fh��dd��-�juI'�1��&��ڍ�ǎ���hy�4:-��uRTF^�'M�Ѐ{�SI�U�9�'sj$�=����P�J�o��Z���ڴ:�fc��񙯙w�^T�x=�9鹒�������E<�nUD�'j�3a7�v�w�#|���E6�Y^����_��u��}V�0�\�{2�Ò\�tEGs��Z���<K0Q\g"��#63&f�y��F�V��{3�᪖G��]d|&�eZ��*�;��lVN�����6�0,�5l<!w=�a�CSY��kئ;>�`���U#Kg/����S%{n�ww��g��ߧ���1;��k�(�{} wϏ�Wn6;"�Սm!K�ELx��N�e�H�}�����C��fhQq�uC�|X�.���Zz��ڽOrC��u��@{�40T���-+}#����ظ�xi6,ڠP��ũuȾם�ւ/1pzO��s�<�a4�ݣ����i�}(����2��-��(��٤��/rmj�����ɝRZε*>���K�W	ݝr�]|-�D��9b�V�C��k���}��{V�N�e��1�FJ�K�^�*�8q6s�xMO��Z&8�黺Q��^҅�{���4���{k*%G虝~��
�e�>L�;�R�K�E�,r6�L!h�n�UӖ$�G5ͽ7��Y�mL�e�Ç#��(:�UA\L�Y�<�5��֯��p�uo����0��m�ـ�{�ƽ$��U���#�;n�4\�@�*x+��z����yR���U����qys�ɞ30�mߚ��+�x�=���h D�X׵D��|�����#�yVN�ݛ�5W�_����gN�鍸�Y`!�̝��=WU�F���֞�X�˺P��~�%�j�F�L�B��)8���uwg�窑"R���5:��u��ܙ;����۝|��G�<	��hfl�멨N�@L�r9:E3tX��*�ixc����c᳔9�@T
���q�u&��$��Τ��&%9���9�t��)��B��}��]h�^v]ȿ��w���/�ʥ\
��x^�|F������/��������ӻ�!΍� �.{~nw������׷:hZ��k��p�/�h��^&:���i��k\�>,f�sf{z���2
Wkʟf� ��h��Kw�(�6*��|��{n�`���=���{0K�жʨ}<�Z���R���{�6�,���Sv!�ڶ�y����kX�B���v����}��bX�C��8�b�����3���C���z�Z��yY�g�}҅��"񭤁�LV��CN�z8:��9fge ��U{jn�yi��h΀�B��*x=�gF"��x�1��X7Nz���"�:����� h�P����Mm
͂�y9��,�,ܡ	�.��.{4PͥH{D����Uw�f�f���մ�&Γ�x���
���	��`����L;�]-/�C 6���u�jC<w�����ô<.�g=*h2.d%-1Vv1H
�}�_�k�z�5�w��E��z��6<�T=`.�8�K���Jj�8}ms<'�ˬ����6A��E��I(�h	~�W�D���Z�0�����]�E� ,%�]a�'��R�r�BC�Y4/�k7u�3�Vn��:3�u���/��U�vT7c�	<k�By�Kxoee��[c9C�.��g��d-8��~�[��*cV���
���jU��t��Yų��ѷ
�dM�׺ҧ{���%RX�6�B��;5�0�뒭�$T`��QȸN���mt?WI��\��4�N@�=u�(�������w����~��z���`V�+[e�����|i[)k�2i��TW=�A���*N�Y��Nb�q�8	��' �,c��� �S��S�e�W9upg2�E!�
.�ϫ�>{���NUڊR��S�{���yu���s�Q����ʒS$u��:)4�k��c���ľH�����y��I948V�P�������8�2ٲ0׾Yw!�%�Yؗ<3s�HE	@�������ԗROu�>|�ɐ!"'�
xNd���v��;>�sK�3fX����wa�	=���q���֚�p��	��8;+I�tc�t��`�Nj��D��7��h��yg'�h���z���\w��1��宑8�P��4p�s��{�r*�T٨Z���$�^�@���M�B�e��âVUG#��7�2��������a����w7[��+�2%�b���i/,*���Q�#c�ĚO���Up�r���3[h� ��OS<������z6��LW
P�c>>Z��@��L�q�[&�����7P#�'խ���+������b�zX��ez�;����c�4���p0п?%;�ܚ�{�w���	��ˬV�41~R��|
͔�Ԅ̂��z�D�l��ܝ걣*e7zж����hY1����v�_��>nL�dxF-̠Z�\�˸Q�]��R�6�c��u�W�����b�^�Q'��%�b�A�V��Ғ b諎oێ�H`޻q��G��Uݙ'Q��d���o6�]b���'���{�5��M�M�u�Wޕ\Nqa�F�����K1�z���-u�����9Q�ÓŽ���BC�,u�Q.������
-�O����wq�o����.�1��7K�C̤6�`?k�ɯL��m��BǨ!���|}���ӾS�⃎{�m�X+�k�^c7HR)�!�s�c�7�0$"v%�WT�W�`G���Q{ӑ+)��V�l�H
�*w��,�쉧FpO�h6:�C��ye4�o��P~p�X\ew����Rm�5I�|
K7���zN�pr�a�"�q+H��s"F��y�=���;WH0�m53Ӄc���4�.r7��:"�]D��LЅ'�4�V�|����b�L�0���v(�lste�cIf=	���<.=s�0�4��ΰ����Tbv�[6�q��@����tsJ����]-8"�8�\:�f��,7��\����*6���&��u'�re�镭r�U�P����r/�q�.�dq���#��b|D���"}Y+_Ӫ��VM��;�J���^��Y�;N
�ȐG�򋉮�H��F�sGa��vW"�NZ�bB�7��;���CB��.N.e�eB�x������:�e=�F�(��ECl���7�0��+vv��f��c��2�܊у�id�����堛��=�z]u�i���kͱ_�����bc�
��<}W�$!TU6j/���~͔ɞ����y��ܻPR�9�U
�ꡜ�;8���z/�LۃM��^�m!K�ELxO����ܷ�9�]������ �ʩ�c���R����OrC�lL�=rd�&K2��n��:sbTH��b�Љ��<�8�:|X�)u���f��A�xi�X��TĪo���ˣx���$��J�P���~�!����Z,r7��B�
����T�閈4��vxp�.VՄ9������T��Y��S�&a�E����ڧP�u:���!~��ט�.a�T:4G���B/%������z��{k������T��&K��L�ފg�1��y)Y� è{P�	�ĩ�j�~2��\q��/��_�o$���� ��{���o����Fy�+H�WLm��X\��rx��M��{%� ��K���s�JX���t�)�CQ�c�uON'Cb��1�j��fb-}U�' ��>IQ�w1�J�.�A��G�(\;ї�j����F��w���pVPǢN��������2��ѓ�؛"ef��O���Պ'��p�]��U�@ۧ�Ln��@�vRSoy�yn�����kZ�Ťni�L��軹+J>f��\W�ɾ��e	7�[�4q^&a��/y�;sU&lA}Jp�n�������]�M�"lJ���R���c����p�8�=��:2_;�ondC#N<���:���V�sc��t��۷�����Ы�I�oy�cلJ �v��`��>z��+���Cὂ<�V6E:�Q�M	�Ҵq��
����n@Y1�0j�vY� ,���;�=-�%��lC�m'��	v�b��6�띭��LM��M�P�dA�MA����V�s+VĪ\����g[�S.Z��X��V���z�]��^+l�"���v�[Jl�2��{���60팈\�˱�(�>�X�,΍�ih+������_K��m���Q�r�] ˼7��;u^�ܵ Te��0��i�a�r���4��
>�6��@��h�螶Ƣ+x�qpG Q��󳋇�f�:�8�n]
wן<'�\Zu�qbR��2v��5�WЍG$+����W��-VT��ST�ˋtZ��y�9��j!��Im����i�W[D�S{R��+qK<�.�Z�7��#�!��&h��>��"��t��%��L��MGS�t ���K\�]9�d�;͓m�7�9�M��ɳ|6+D�5(i�M�����LM|Fі6%y��|e�h4��]���hDL�D��5��:@���Ut��]C������ռ�8�PT�ٓ���SK����,�J=W�u�z�3M;u�k�������W�FV���eo�NJ� Mvq��- ����[�u�d,�B[�u8�]�U�-��ӷ�7�:��m��D�y��A�N��O+X8�݈��X��ku��hWŗ�{�A.���h��h�4����8w-�E+����X`H�a��Gk���EeԬ��Vz$��K��P9��JT�r�
u-�!���.�8.�uj�����N�Ev��wC8GM������������kf�y�m$=�7��c�tD,��Eb*��L+@��5��-��3�f3�>���ϛ'���=�o<�(�0l�5��5��֋�O��|;����(Ĝ��9;�Eo*"v�;�8!{8�(Z
�i��djwPqBN�y��3%ε���鵳�8�α{�a��O�f0�gL�h�gn��IF�sO6=гz�n�t���%���!8�X��:�φ�U�^٣nힰ�;Ժ��O�>a�ˮ	��,Ey/wpBs�(KW����9Z���s	�]L%}:m��G/C�!��ZC%s���-qR���.�m�;�����	�BH�%F��
ȤX
B�E"�m�-�����*�U%[dEE�(,YJ�k؊����PX�"�Qb�Vڕ,@P�h�-j�(V���Qb�J5+%B�#Y-m���PQT,j�J�l
�,QX�ZȌ�+*V6�JȨ�U��J��J��*T��
2�*E%��
VVTR��D��
��YD��Ƞ�VKmV)���ȫ"��l��dR-������QZR���[HVV�YU����aP�V�E*Q���D�`��+-���T��VA���KJ��B�5+��"�+&%@m�X,`�T
�h��1��E�1P�,r�A�-V,EEPXc&��PU(�`�ʕYr�Um���-eeh��[h#��YT()Z2�qV V �Q��ZY�3QkT���XɉR9HfU�"�%~�ȫ*�RkS��&��n��t�A5�݊d
4��6�A��j0ǸAv�#(��$ !�Af��'��7D�̎@J������&��j��tX���N�U7�,vV�=����3]ēQ�X�N�@�'!��t�Zv���9�4mnM��Y�n͏b���)�6��9{x���{yԓQ�TMBu
�,��Q��s�Oj��Y3=S���~D�5a8]�H��T���0���vP�٤E��)K���r��.�2p	{�����w���z�'^Tᡪi���4��-���(Sq�����V�+C�nX���kVE�=��8���z�8g��n*��1Mܺ�.l�<xuډ`;x��R�*h��[�F2�*x.�Tp(�XZn1�b7"�`�9up��5gq�dj-�������0Ejs~>J��D��tÁc�g�(Bf�S�c#��Ӂ���zݱ�T��+���s8m���<���}I-�
���ã��<��+�P{bIE&���Oef�'2]j��ظ�O����A(��n:>������K�H_*�2���!�;��F^5���d�D���yL[�=�-a�H�0������q&x+�TP�r�������G]%K��CE�o��n9��\st�B��׈�� �Ҧf
�ᐬn�C�]oQ e�Np����00��;���suhv�USD��]���N�{�Y&.;�yC̈���'�&�\Y�Z�U��K�U��1��Њuk��U}T�o�_�r����09�dЄ}���3ʹ�^�hl���*�.�^|Cݕ��L��gT��rE�}Y�称ߊTƠ��>W"�XkW�)��h
�) �WKF�[&�y�U}�����c�.V꿂�\580%�^�n]��ylX�Y�Lf�+-����׵㶒<25�7�y�!�����Za�%[�J��܍��f	
杹wx����G���&?7t�'ߊ�%��#l�_�E'T�X�Yɡ����0��ݐ�tY)���,Ί��6@���r!<����Ԓ��D�ᛕHE	Pr|_s��9��L����\7=d���&��?g %�zܥ���׺�CԼ�^[~)����2R�.�?4zå������t��p$W�VE�ei7΀��{q"�����"�j�SBk�h卤ҭ��$�W�{T8�ض�����V�����D��Cw��*9� 0^��<�X�K۷��]�u��5?%�	s��̪p/�QYU����Ƅ�%[t�q���rōx}��j�t7�n����Si
-�ݭ��XX� �އ� �5y~�ŌkW���a�?<F�����t6^p��c��n��5!p�G���U��B��y=:�Aʖ]l:�-2��e�R1JYv�]*wj5����SvbJ>������II��qV���cIu�f�\�5j��-��;���-��7��#��-���I���B�@�����b�}U}r�H�I�,��v�@�)�7إ�x����;&��Iǯ`/@˯k��=W��u�}�qݺ�c��c|Dk���*�pѕțxZ���3�e%�΅��ncC�����Jޜ�[R��C��bU�ˮi�>�^��6D�<�s�nhdg�
�CT~KFs����'�}=�?*�3��ۈh�v��f{-�31.w���.��d?a
�8*=&z]v=)�x�b�o�ȿS�b2���Y8��ꝧ���>G<������9۔hw��U�|g���b�cԆ�:
>>Od�j��6��E+�zzH�Z�����Y�Y
�=��P����s�To�]U��5����ՙ<��l��՘����$��cj���a���r�S���p�T���J:/U1��zP��R	�qbi��*ڪB����4�	�XF�a��UB�)�*�D���z����r��\�YL̽Xf8�ou�r�y3�u�}�5����|�z"ea����T�獋�K���K'e�q͏�0$D	c�f�b�KF�Sb��:<Ò�n����}�`X��%�u�t���;��δAZ��7ײ�>�D{�N��Sg��u�{&��`�>��H�̝�������ԻI� f�f��M�r	v�f=F��AR�N�9�,eӫgt���uM�(����@�l!���w|�"��O��i�<1ae��mm|
�3^|���7��Ō���傝V��N�N%A��`�������n$�s������؄�ۏQb�ٳ�ǦG��LO�����~����3��뻁�.�Z�ֳ�L��v�`�6�t�9�Ӂ�mt���x�L
��q3�iS��;/*'7�7���Rf藷Huçv7���ԭ�v������W�$��*c�X�u���me��~������� �U>,"�,<��:���)�H` P��w0�US�*g���WTa��$�`���LpA��yqPr/���������J�����S�ī\&�h��=b�"PoЯ����poH�/�����N�*Xy����s��z�l���q��L�)QA�E���f:�T<�r;�F�D��e�����V�q��/r�B"�3z���3�4ϊ<B��
��O�P6\n�L�����rr�ߞ�Ԭ�+���RK����Y�
=�3PIդ���[�e[��m�g������[�'ٯs��l���2Mv}�� �&��W�}&eD��%9f�?>�!S۹�^��bbPu�G���)�\+$��O\�M0}=Z��S�F<w|/R�a�u�O�׌�}��ܜ0��V��=#.{*��8�7������X:�)vpg�B��R�9��9��Ч�=��+*���fu�(�&y��n������8]o:�B��q�P�^N&�Ź�5�U+���>Ȼ��ml+���l����!�`v������L�� ��G5��l̎G�=+`�s�I�5�6��߈�:%y[V}j�T<6�p�x��6��?��P�P�]6���zE;��V�����q�'�ƣ^]Ȱ��/��*�/�ϩW�z��|D$�ß��ˎ��69m�Ɏ��5��`���b�a�y�i���l�V'�Y�Y�nD�?U��)��݅/y�۠���\��L;�b����Y�j7Ny����dpƹ��-M�;T<����m��g&0D�ʀ�#qQ�\�����XZq�b1E:��r��4]��V�T�67a� >%Nz�F���p9�k2��X;%�a�s%�s��o Q��rPbFT���C\$���",��-��tT=���Z���z�K�H�N��vn7H]��X�BJ��c�kUe��h&�v�Б�'�u����:���z������}k�;O�$����z%�	u=J�=U�C�|b�]���LoK�� 6X�N�h�ב�Ӯ֖54e��28;	F{�?I-���X����b��x7��S���i�N+{��E��7�x6t;�PY�x��x�D	E:��&Z$V)���a}խ��|�)x�R����n�Ԍf���ž�Ӎi�W���K'��^�	|kGnu�݌�O�1��5�{�|R����N���t���GR|�E�T_\��}w0"�� ZXax�n���>s����R���vv
tƭ.�y>U"[��M�p�S�)��O#ە�1�u׺�R���@C�11��o�t��Lj��X�g�>f��b�x����6ob�
�!����HL�'=2�t���Ƈ�E�u�x��c�U,�fA�BƖ�k��FG"�c��u�L3s$���e/-�\5�b�?�����h�ʎ�g���}s�kU�I1���܁�9j˸hd�,(ez\��Ȫ�J��g�����^A�>��gS�,���N�
2�N.�$\L+ڙյi\Vp�(��Z�X{�%l�a)w2WhC���p�:����@N�σ���,߂��g.���]u �e��@ޞ���{9��*ˆqr���v��Y	h��d	B�^"���T��Q��T�[�<�u}����$�'=]4���}�� �>v�7МJ Ts�2�ʺy�򼺄Y�í?-܈�D�:����O�eE����b��r^�GA��EF&����y���{q!,QCt8��;I�&.��{7 �t�(fv:�B�f�ôT\e�c78:+�]"o��,h��A1C#[0q����ꎹz��"Uy�%%�	s���o�%����Q�����)�HJln�w.�.aaVru�=�k�DAZ�@yv\;&+5�
�����+*x,م����4���Kޞ.эQV�Y�e{�*>�����L�)ٕH�>��Aqu���$U�B� ┚gf{�r��2}��C/�#-l�>���7oԳ%�<$a�#^���Ǣ�xpb��w}�X���I�c��k���r�ֆy�8�ԅnh�x�1fQB��Zo�ZʊB�"/�z+��_��Q�P{��*�+�t�7�`����r8>����T�.��j��'+�2փw��pu��aTK��8�V�Coz!��U�=�C�T��[J���,�ipWj��t�
�e�W����R�|���Mp�3㧮�a��#}�L.�Cqo'k��[�7���IN��� c�;un̷}��c�"�@X���H�:�3J��X[������YΤBae������B+��{�ؤ��Я��;��5�7�y[�T(x��pPy����d����38�?������1B��]�u�P�ʘ	�8�.x')�Z�9SZM�q4�K|�����vzM˗�H,�T��a�����;;��H`����=M��8��b�en���N�rwv:��Tpg�ʲ�_�� Rq+H1�fD0�N���=�^�A�/��\P���F�7���Ǣ^,%^t�s�X�g�Rq+I� `td0-uh���˵��6j��z�6bϙ�n���Ìӫ�Q��w(����@�f�]>��!z���ǃx&44APw���>x��GY`z�{��4�;��OVӖ�Cp�<��as�❺��+^���ױ	ۏQr�T����Y	�q����̛�y�dE�㗮�O+6N�MmQ{k�P���r-�b�Y���j���B(��Y�Wr�%$�P���T�m��P�9O2v�ʝ���P��7/vU�avDS܍8���;F0(�U���@���z�G���Oi\"<��)�u�F&>�9ƭ֛��.Q�yI(Z!M �}k�?-=h_J��&v2!����(��+���Q݆ڣ�?�I5t�u�4��঺�]���� �)۷��Z���xX��`�.G�q�u�MoU�zs�+ӈ�T�}U�Bz/I�G6ğ����:XF���_s�KOS�;TSܐ���f�}W���T�ו69�|r�����Ġ�dϬ�(�+
�"��~R�|��oC�g�6vL��̇U=��U��RO@�̒x=��Q2��	���HF���oT�3s�[�9��27���}����J!:�3sW����-
y�Ǒ5�����3�H85�F�{�dM�:�S�a�%C�"y�����O@�*x+��E�%�cFJ��}�)��8�`qr�
؉u��A|���w��Za�����U�ۏUQ�c�ў� y;�-yg�W����U���B.���ZEºcm��u�tu��WM���[�ߤO}���TW ԋ�uBE@f��B��T6uCF��0�̼=�M��cX'���VtW7f�̜1{`�0���R4-S<3�!�r�J�V��IW���{��N�|i G{&�=��?qRW�W�۴�1�	�+jϴ�L`�ܪk���h��gSJ�ͩ��g����?W��.���)d(�#��q���e�̣�+p����J���.��,%l��0ې�)��6'7��8��Ą�k`�|8�\�V��]dp�FN�Λț���w�W
	��4)��Q}c Fk�c2����N��L7��>��=����.�2c�FeB�MN#��9u�T�	���zB>��@�NK����)��7���!�t���������e��P��X�w�R�Ch{�\��Ph�_�����*/t�#��7�4>������#�֬��ǵ���z9���8:�[�%�����e��z�&��Etˁ���ʞ}�JΌ�XZo�#r)��-����#�nz��Gs���]�pe�X�ĸa/��T�ꮠ���f�Lו;�3��t���[.�dL���UǤ��q}l{K���]&�\L�I<�)���x$�ˬ��7�Ɣ���Ã���B� ~󼖘����Af�O�ObL�WN�"ZH��X��7��I �:�A�零e�Kǧ���͏>�j��]Hq�� ���h{����?vJ��\� ��3�F�T�,9������B��,N�e�m���"�N�
����2�w�|�MT^�O��zJ��xBr� ����r%�Vk�WF�?yћw�p哹�����ְEjV;�Hs�GÓ�ޥ����h⼉r�-a���DT�|0���"�
�D��<��%E&�n�ѷ�#c���k�9�nɼewf����M��\�R��U�#�5�0��\��>��rDdM��2\3&j�ۜ���6a���:W�����{�m������bI��8����Ȉ�{LҴz�wy��=+r����T��]�\���{`S�ҷ��n	��v�(f>����L�GR�wQ�9Av%��6��9wL��g��F\�ܼ�8u��3Q�Vө|�s@���i�rT���O���!9~
�x�z|<�V�гm��:ĴxG���ۍaΙ5��B9C����>�O2�:RQ��k�액U�7���㲕wW��}kz�폹�7�E�}Ԧ���%�T8��<V����ӸrF�xn�A�ub���L7�fQ�W}q��ѰjP�I�0������[�ǳ>}!�´���A�}��7K�������F�u-���5���y�
=g����p��
�=ɹ�>՘6�ͷr���~B��St(��vn��M�J���U��c�LWF���۶5^���t�z���2s��S�x��86�t�g��v�3<f�E��˧�`��iص��v�%^�8�E�B��6����dS6,��oVܫ�#:�C}٦;��i����5v>n���˾�|�. �Y�v��c�2v�ShT�8�u������Z^8�������豐aX����RDA��lh`�vD��`�[��@��Q.��v���E�u+%�N�h����sfk\
ŧVQ\�s����fΑVWS�	�U��5цN!	��y5��yɤz��Ϋ��Rq,Nv����' woQZ�INL�9a��\��Y���w�����,�F2-=`�0@�),:�Km�XGG��i<]�J��uI5�5p`J*���S�B�"f������bgn4(�;b�x xΫ:����[��������H�i�ZN��{$ȟw\��P���-�����u��kP1�x��v �K��%�v�2v��#���'�h �U�eF;���#�7��p�,�$��H�٘�	e�]�k��,���K��q�+O9���i^�;Dѥ�Fg_Q��Q�;�sj�Z@V��k�$s	���2QǙ\�^�\J]}��{�9������dY=����/Wuhfsjv�5c-;���x�a5v{a��t�)��"���S�S�w)*sӛ&Ծ����:�FsZ��[��FD�n��9F��ĎB:��!#{�B�_T%��b�o��%tZ��v�ËmfY��'窸���̽o��4��q�u�Uzr;��A���(2������]��J�/;���ޫV_�%X,�v��P�qy��9b�T):�{`,�)r� 
 x�$@���`�m��,��X�U��e��b���*b)DU�ZJŊ�Q(�����ѥP���*T*���*� �(T�V(,Ī��Z�G32c+l�����bb���)2aFV�Ķ�J�ڱB�VVQX"��UQ"�PX
�%-�E�Q��ĩ�%Q�PR�����
,�W2�q���LB1B�X�U��DV�J�J�PYR��Q*��P"��+V6��J��Uk(�Ab��K���aYQIR�\j�0&%Vȹh*�#%JȮU�(�b��Qd�Ѝ�IZ��H�KIE�
ʅb�
DG,Y��ȲV �
,Q\@|����W�ËD��ڌ/J��]�����Ü�PB2݂���!�"�Qۍ��-	��`E9�Z+�H��Q�sv޿��z,�ݽ�<�Cl���H|#F�9�a_N�؃ʘե֍��-�G.Ao�ye)Ʋ����û�C��E!~�p�'ܤ�$�'�^T�u�-8�W�-���\�r��C]{���Vi�Q��l�9�>6�"�f$M�f/-�\5�,s��
7�r����nΠ����2K�t9�S�# T'#'�p�!�%��Թ�Qݗ[�[2�Γ���'jb_��証U �T�)��	�@� ey<��~;�W��K��N�=��G5�����EbZ vi��Y�z��]n�PA�&���vV��@��w�h�KY4���]-6*��H�5���jي���/�Q�1l�@N��Q=�����Z�ou�qI�uڹj�Ec�{Q�zȘ�|����^�,WTJ��V�IO���-�5{�z�]��\ksg����l/�-v��
��)��k�d�czhŲ7�:f�ɭ�'�m����u�O��� �ab;���=�����;2��}���.�{�빜."�\��\*G�+�|Fd���K�d1a��$��Ы1� ��O�v\q��;>�VB�����PW�:r�ޑ�f���آ��E�Y�k��M��S�F�=��P�ǯ F>�[���B�Bs�f����5Iڅ����;��]W����ִܳ}`R�G��D�c�"�K뇉>����~���W����c|Dy�f0���8�t��N���J�~�%�^�,=�v�1��R���|%oNC[RÚ0c)���x\ѻM^>�|�4n@~&�:$F�T꣮%W^�(=�vo�Ⱥs��1(oUb^��c|Rmf$��!��8=�4CRQ
(��
�zL*�u�oǥ"��W��+�9���Z5�[S��hۊ�(�7 ZOX���n�ٶ���f�%Q,r7��T({��lwV���m���})I�&xV��y.�P�w.ͺȨV�����MK�
�*���L ��
���K�M%3[�H�j;�s��XS;�q�Z���r��g�YM![��T��:�\5�p�������m���+�?l�,Fi��U!YVX�
i��������>�d:�T�F7}i�h�]���w���#�y�o����~�`�/:R5�١a�P)8���3oQ��v�+S�N�^Y�lر�H�[9�G��X�u'���k/<�	��N���Ө�K��ٔ��M�",�P[f�)�坵���	9Ҭr��o�DZ���=�S�܍�	ݗwț�Hd��ZӾi��*�(��/��Nlp��c�F��y�..'��r�GLХ5����_u��{��R^��Q��9X&<u�a��h���)��:�\�)��;�#Ԝν�J�V=+��P>x����^�0�6v��z�D1]e�ɍ\������k]jd�B�T�q�Q�X��u�\��k��U�0߹v��2�l�HpJH����uLYgE���}=�t���Kǻ�E�_=��dZo��j��0(E���7�lR	>~��V�j����H5.�f�:��.#��;nX]/.0��u�m�{=��f�wv�5Zc4��Wy���������.9
]F�V^�L.�+�sEZS�y�[{�ٗ޳g��Rֽ�4�!pBb��f,�(߱XT"��j]r=�JÕW7��͵]���{y�[_��,����r��n�l�M�@�r�+�<��i;;��o�_ {/�+pw�	��[�5on���� ���Lz��G��<w�kّ�ݐ����]1�GR޸��uܧl�
�C�"=��=J��A��1Y����婽���D���*
T��Ī��S�F<�o;+֬�:�h C��g�&�d���P�Qn:2��Bĭ�8�����CXZ�7\��+K2�����F*�oCiښ���L��G��G+=�G�l���o,����5B~H=�y���*X+����Bs����i��(!x�3�ֱN v�B���0��Dʄ�Ynl�g��E��5����U`�
]���_��p�,�VT����y�C��6�zOB©�C�Y�P�N��:(of9�[���P�u���u׌��90�:6�nH4]r��t4V��G�y�L��W2Wx��͜=t~��-��i���f�V��!�n��^f�jr��� *8l7>k���,u��|,�4zJ{h�S��`FV�m?mJ���������]�`bX��d�^^Xu.��hw�ZsJ'��M�~�7��d`u��	���I�-#����n5�Κ�4�y�^E�o�.��5[z/0`"p��S7�AE��ŉ6�d�y�7����5SϕK����d�j�s��v���/�Eΰ���)�]B�c.+�u�_U+:1����A��
�i���Xǚ���|z��I6Y�f�y3�]�&X�m���
E�E��&T��~Ϋ����wI|��bM�z߄�S���=ڋ7)+�Ih�����`
�<��ع�3h;�,I��C��כ�����2�I�F��{W,�ں1��\�0I���Mx�ٽ�JK�����_KX�MIw(n7�ŻaCz�Ίp�]���%�%p�H�`��;^�\��Vj�[�zލ�*\V��p+����+%��pи��
�rZ�KiRVsdؒ���$�=��P�9���S�,������
�&x+�T��9fp0�=��D�)��.渺�ǧ���͏{UZ�C��(�����a�~�M����֟p�)i�OJ�~.P��b���:"��/\¢��Gl>����ޓs�<��Uc]"�2Z.�&��,o�z^)���隆��{a��{��ϰi��8�1r����2�@ B�ba3W�aU�n��ʘձ֍
���m���#/Zq��n�$.]���U�5�������Y�~"5@����qk�C�uȦ���$��֗M�'61�ڨ�c��X,u����\y[ig�sFb^�ts~͵|�:�zT}��T�Mޙ%�qa�pR��.dYI���z3=f���mP��rh8|{�������WTb�e��(A��ԁ��Ja�Bq(Q�@��yWq�nt�.��Ҿ�p��̹�ӞK\�}j��E���3��u8+VE�ei7�tTx	ahe]Ӱ"����R���pnp��D����%^�@(yf}s����x�r��Oa���y�*�nsNN��TZ��`��	b󀌴��.�q�Rʩ�j�R����/�.\ȡ�FvĴ6��$v���v����P��������3���zIZ��W���x�3�f6"���ôT^]F3a8:*�D��\�q�)	�wxU;�7���0�(Q���f�}�w7�U��u1z��8+�ַ[ž~��2Ԉ�1�s��S'n���m�ct��Ѩ�:4F����;�S�ڐ'�d`����e�R����H"�'��t��d"�i�3�Ӗ�p�[z.�"���^�]p&�z�)����Ww9@~˞�E�ɿc�"�����e����V��3nߖ]���F�si�k�r�����ڎ�"�_�e�r�]��w�|��ڻ&���L�}��2��k��ge���fi���b��8+]+x�~n�.zK�Ԡ�#]��E�W"��o*E���Z�,�<;�g]H���� �(��Pw��;��x*n{YH"	�~�DÐ���nE����:�5��q]v��]�Y�����d�v&X�L#+��߅/���n�i�ऊ���,N�ܓ�8s�朇���E�sq0�'�0*�5�<_���:���݉��Z5g��mJW��������1q13X��*�����\��X�X��C�a�����R��2Zn)[~~R�c�>_}�I�6Zi	��)�6ݕP�N��D9e�tYyΏ%:�z��[s��x��gn룁T�aq�jq͌��Gv/#ң���J�^��{~a�NJ�ag��cr���w,EC���~G*I��Bx���fvP��%�ĵ�Ƀ�8�a�<6 Fi�s!�e��
i.�Z@a��:��c���0�>y'�d�h��b��-��x�^�Ղ+c5\I�ݶ��tT
�q+ILn��cX�	ʅ���z�H�v��M��#3�fk�K�*�9f��3y�A7+k0��.���[^����;j�M�4�v��y�"��"��,vl�\�Q{T�����p*&�g>Y��0���n�I��EF��D�s��9�ph�kΈJ�Ǩ�j��yX���>����� �iH�m�д�/�K�ߟ�.����;��Z�د�E����x��	����[H����A�Z���Hqnh8�-�~��A�*wcs�Ρi��7O�w���Or4S�4A��z��NҞ)-�.m!J1��\����\mB�S��)u�Xw�w�.9�I^jYU�7lm���
�3�]�L�*v3g�F�1XW�|X������K��h�ݬ�~���(j���i�v��P��o_��Zy��Oj��W��&�6+WĤD�E���z�V��^�6�+��>��#�� �������E����]���K�m:��,r`��Ǡ�i�E@1�f�=�L�CK��A����{�,kA�	rWk�m��᰿�o�����U��Q��<g-�X���*��/b�&�׵��/#�\Zy��P��\�E�E�<��G[۹D"B��(s&mUS,���q�fۯ��ff�œ�0��,��uܧl�@aQ�}$B{U03�%�����/H�k�,�G&,��w�e(E��r֨�����N��p�|;)Y��a��0"z6�[&����[��}�������k���Z�ᳫ�삫XR���P�"��j�"���V�8t��C��@��rx�+OU�B�^��[����p�q�q�XS�_#�.H�:y�zv��,]���<.�ad1¶��Hpܫ�+���q?��;<��n�lM1���t�l��#�i�)��������-�=�/�ܸ�=��>3�d��]*�ei���$�Q1.!:���GI��!����7{���CDϸ�inK�5��ֵ��2�!�N�c�2/f0*��`MB�`�O)h<�i�z�&�^�顔-�m)��o2��'r�9���r�e�)�_l\*S�9G
h���|r�l�ˠ���nR|,E�ky.ڔ��Ak�|6�,u*�+��8֔w�3�`؈�6�]��8��Tw�%o���J�r��R5(��͛r�=�T盀o[�Y�b19�������d����u�qbF��Y�c0�M�u�P[�ggއ9�gK�6���V���^u��p����_���������><}���,0__���f�ܣ�;b-���n����_�8Ս'd�X�U�a�Q�V��+~#ܮ��2x���{�/{�ް�eS��3i��+/�E��X|I:=���T�x ��ݾ��t���kz5�ZB��8�o���i�>������Af��{�MA��P=���&%�l�{�R�6��]����0��b���{�A��mi�Wц+Ĳz�[Iv��|��YPT=�EX��Z����>\*_ ;jvM_�>Y�����2:��O�����$��3�j�?x��-����'Uԥ�o��	����O�H�n���w�yȳ�|�k���k԰�ܽ�"6�i�D��;)=ʅ�Ǯ=šOW�����Ƨ�G=ĝ�X�����Bs+P�[K/�e�}X+��X�,	�D��
ኧ��qi���8H��HP&�Q�8��m��
'v���2��;kD�$�G�6��hJI�.�c�����D�+1Eq�ܢ��v~�b�Ӯ6�p �)'%�v�՚�*^�};A5.�wf�٪��<a7#I=�9G�7HH��b\i�q#2���#y+YGx�e��"��2�[e�q�Wꡇ��h�P��|w�SJ��3�	t7�:�ɷ�b�my	��Đ��_8��Tؿf��k�+���N@��P��4�]��v��-AXpD�
��T2�2��y(�/<�
_S.ΉT �._���XQ
a�D'��rRyW�.��u���67*.�o�p��Y�7�����b���G�|l��M�dW3�H�,�3���7{�Tz6���Cվ����/'�߭9�S�Z=Q��T��rr.��_gs�;]u*������(����X�滶�t��,^̸tB�����F�ͦz�fѸ�.#k��reV�1�v-mp�/N���:��d1r�g 7�>���J��^r�Jw�\C����
�T�w�W	+��."ۮ�KoE���V�9E�6�y��oc�cƜ�ͅ2���"��M�1�/���O����i$L��k��/��8�E����Cr]I��qT�p�Z�MF)a�k�[���/���l�z1	�&tb�G%��\M��ŗA$��P��:%n�h����̲ę�=UI��ɔX9V1\9�W#c�t�&:��ڼ�q�/bq�5�U����`�5���]1u��J�ݢ�J�I��YX���˂�
����จ��VK�f;�g`�V�v�(�Di�ѝa�ő �kӔ��ShD6�a���z��q�7%�12M��T߶�5x{DTt�2��p��>���l*���wK4-�:O`�d�SmO�ZGw,%r2���� n��[y�����ب�#���,�I$�4��`���dܜU�\]�'C��R\���,և2�l�~vop�V�6-`�Zy�����p�a��V�_)�d��%�f�n�/yR9ғ�AЭ�vY��W���k��m�+��"����Ӡtf-�����y#����;��$=�;eo�O����1��Q����̔q�˰���N�2��`��d�%Ћ�9��8`w2���3�Ji*쎺b0]��o70��)�o�v�ul�"�SY[��ɇ�S"��c}w�cB��jH�{.�V�7���7YC,�"$ץoJ�­�}�GF�L�(����C��G�?W��m�9[�n#Z���G���u��P�e�P��j�-=����;�:[n�Сo�����*��Ae^�M�Fe���˵K�y�<�=�;5��Ԯ�ݼ�&�*&����('����6��J�}wri�e�5��$�� �t� �+f�v �<���wzGu�\V�P�����۩����"#�I�0��!�0�d��p�D/�gz��]�g(�2mI���������^ӧ�뒺k� �ú�dwX�q����ߜ�k�Y�����b�����X\�3[�s�����R��o����X�-�v�;�)lL[���dju�Wz���������{E�R���Z�l#ˎzR�ـ,f\�G�����촶Zõ�8z�\�z+�b���gt�Ɂ�tN{{Q��X�-�[݃)q�@�R]F�����@r��k~�4��"�x3z�4˔��2Zh��g�}���x>�n�&���f��\��h��@�m�C�͇�\�G*�-��&t�JI�����-R����K�6�;a[j��t�Q���Q5�{�2��#��e�1]����*�4�_-7�FL��u�
�C��9��b�&�G([Ud�^Z�7���ȭ�D+cN�jA���e���'dQ�FJ�`
5vw��`Ι#;h@;:�����G��}1@��/r����6(��1�t{�P���ٔ��\�|�Z\����Cy�S��]�ت��L7q��y�B�8�|�w-�&���n� s�c�����S+���t�9M��z�(�i8�,�!�j�ir3v�Y;�Z� �\² �
n��1fxh���:j��aN����,�N���
v���ͼr��� g�f`�9���w+���{�_��R)�JZR~j��mAAq����B�TY"�R�TH�X�*���&5A%J�%EW���r��"��ƫQ�i�A�V �X��J",r�X��c�3*«&5Uq�QQUA�e��D˙VD@c,mj�Ʋ*�����8�E�k*,R҆&e�2T�LE
��H��+m�@�.P������RW�*��UQDE1*)ib����(Y�
chr�X�+F�#mbe���XVQ��mQH����2�V��j�RV�3+��*,B���UeJ+(��2�ikB��P+V�
mjԩch�.��w��nκz۬��
�$R����2��Y�6�˂�m��� ��}i(�#�200[YҠ:���.ْ�:�7��ymf!�R7��	� p� �G�N�:����Py��*"�+�'��ta�Ox�Hu�;���G5��;��t\0zZ�k�s^F�^0�D>��C�T�pzR+N��W$JðS����I�!��W"�S���:ͧ����S�����9�W	�o�\<�G�K��5�n>Z��~|��9�5u��(ζ��:ȨI�L��Mz\�TkG��4�<�v�>���5�q�q,4��"%e0�:�7<Xtvùb*�T;�r��dK؝������[���/��k�0�f�R�����n�O��8��_�m��R�o���s���'X�b�l���_���q��xg׋]櫉5�m��D�4:3Wn�y'V,Ѣ^��(���j�mZq��k�Ve��]���i���Q��]��yo��=3͡a���|hË��'Mod�o����<ͭ�W��U����xt.u�|Z���3bV�7^��մ��]�q�GIb��B잓\b/E_�揖ߨ'e��P�K7���^��\�3�w�3B�@c.��m���$��0��/sd�B'bBö)��z_m�wF��s��u�ҷ�>��<-���|(��E�3��ԕlkԵ��N���y�1.�)�뫕��U�B���\��\ü�stJx��t�y:"���uB6�m4_���Ɍ�9�ئ;?z=�6�PsN~4�'k9���ޢ"��jy�!��)��n�w
��܎uL^7O�i�;\�l�ܫF���O��[�MK�R,o p-p��p �uӁq҂7�52����� W
����f�%;�?�Uq��������.CP�6�3�Y8FD����'"�"�*�n^��(�t�RM���[X��ǵ9`�6�_����\l(�"�����-�4�k��A.�9�KI���f��3���f���p���>��}����n�*HQ@����A��d�}|��ܘ�������Au�^�
d�x쵓0��\L����,0��>�!TC۹���F��^�Z��5Q�����D��[�a3�֤է�O;8:;��U�y���.�2nXNܤ�C̤6����%RwJ�LJ^�d�Q}'MF�oaU���gC(V�6�F��\�uu��v�X5�k,!�d�P��5ڥ6=���h_5��Ψv����S�n_�F\b�a��t��t��y��^����N�Vm�$���K���NӁ��ۧb˺dX�x��v�E�������%� q�z&`���]&�Y>7�m9���t���61�<;�H�T"YZ��	�#�v-[�ٓ��n�|�Vk9�:6�i[�go�������0�"��u�h?nuůk��<�5�/�iI������'bI~ܖ"k�ڀ��tBt�f�~S�8_"��C���T���o��R7,�׋%rR$p�z�pK�)������1��疥�Nf*�v͕��|@�+��;W�N�6�mp���<9k�Mu�o�cT�d���H����Ls�Y`��Wˇx��y�f=�o�>V4D_�h��U�c�}���Z����dw��u�d/r��-�K���^k�%�QI�vj�puo|r���Ӿ��"�e@��\Te�q�J΅�@��0�Y���.���"x��HF˛���O�EVu-k�o��|q-O.D��vxbq�}7�C�_�JD6��W����3W��ۉYx&�&pR$�}N��0���K�k����f��� ~�P7�3���"�i��P�0ٱ�~t|]Q:NًS�r�{&s~q�[����˞�{��pTfT#��U��pX|�.	��k�Q������
`M[ML�]1b�Z�_�7������D��<�MLٖ�h��o�?/m��f�|
{qՠ�<4f�E�#$Y�+vi�@ei��K��4��o V�[�7���5��R���I�/Hw%I�P]�%�ыYr��)#1>}�w(�s��x&�7�j]�����$�%ICb\�!�"�H
�+D��,�{aQ �y�e����;umcn���GgULc�t �`�.�����K�~)����'��OyUv,Q8LrR�m��̱{�i�e!v�<hv�jy�K#�e|��@\,z��[��yS�ō���4e��s���JNp���f/�.��<�,9��5�$��GIip�E�����;o'u��x���h�j�G�ƘCuND�w<T`�>f���:�WV�Y9�1X|�H��t�|��os�V9�Q���Gf��oT�Q�9�a92'#'�p�<�Ԓ�a�N�#�e�'�ۛ����b�}t߅/�v|)�"�7z4� T'��s//�N<�q����<=\��h�,��h��L轘�p\��y�������"
6���c)wb�r盧b�K��D�3׶�^�)�B�?��w��9�N�7\'�q�Gr��`�Ζ��n�͙L�B_���g��d�0�Ӝ(�nm�W�g5���MzܱQ{T�>����tP����[.L}�<�W<n�Ē��F �,��b�/|������	*{ɯ�J=3�L��cs��)�����q0K��d*u�����i�{gJ��-���}�;���%���x��)� V��FÕ;�Cۈ�V��$�Q"&���t��Be�ۦ;������8a�'΢�������c��Y����ǔv �rWy:�����W	+
�a��r-���KoE���Vx,F�d��̳���\��nOP��J�ҙ"��[&��P���@��
	Z��xW�!lu�z|���Y�}���)�	�#d�zLƫ�p8U�D�,<�v�[���ր��͹��shT�����=�Ϭs��P�	0�bDO*��K��T3�Ƿz��&0��n_&�ś�ff�8���n��L�a��j��%�t���hz�{b�A�@�-ڞ�2F�u{��Xx�t!Qo�ȸ���ec���p��B�����NJ&�2�#q0P��ɜ�37y7�w�����?=;c�r�]iъ�]��Y
������Ne���Tԉ���<F�2l*q�d�
b���P5��%\��uLha���f�W���> �]���x̓��޶@���.!�.*��5��M�`�|6UO��K��9���gׂ!O ���y�_�_kQ���6���7��s��r���*��ۍ*F$�fYe�n\�!�i�5�o�cj������Cv%�(�a�^f5n��P�yV�H�)��#V�����fZqqpƘ�(��9Sz4�6�� 3b����s�	c�k�wn�����e�hg�=5���Zǭ�a�I���4Uٝ��e%$���ص�F�8��]�Ͻ�t}��0צ���<6�e��]����/g�Փ�d�Մ�q/�ED�'j�a7��E��0;�"���f�z�P�͖%1L`Y佥�=���.נ{��/��mI��f��@�� ��ڽ^/��E�F�V�y��T��l���W#ޓ�YvY��e���"�'CdmM���m�����m�q�s�X�82�{v��w*��Z�Ջ����B�*�#>�Q3�fk�%cn�v�ݍ��P�����$63W7`_<Y�zzw��/��BF��x5g�cܪ.c�D']8҂7�:�|X�,]"�n_�X�;���5Fk��h��>�+��k���Z�kLB(?&З�:��N���o�	{\�Ղ@�cp�j]r8�O�oϭ/���zTF�+��a�4��=�X-�x�%޷(�Y������D#]�R8!�\>��_LT'mS��||g*��i�h �7����Y���E�]����GMZ���<��Ts��]�]G(M���9	y�Xú��7�oG�lr�-;�W��C�9gt��*���J�T�մ��f��-㔒�>������=y}B�Rճ��oh#ۈ�2���R�0������s����*p���瓐a�ꃲ�w�l�Aѯ>�!S�쫾/G�I��S�݊:�U����E�%�\��OY܉�A��l`�<��%��Bݵu�Ԡ��Ayk�L�����( C���� �j�/�[䘾'N�:��x���K��:�NAn�#&Mޞ�R�x�m׎�'�Ob$9�B��T�C�P���%�FΨh�M�N��N�&V���b�S�1���8�M�a��uwa�S�����u��S�EߏmM�2]^٫�6&��k����NWMG9b%:�|��v.<�������B�/���b��]_S��T�D%���aS����p��S�iJ��ʶ��W�	�#
���!���;��	Y]6gVC=w�,�K�����W�<}i�D^�`u��`MF*`N�`<�i��h���S���5��mN��e4x5Xa��yQ�r��G��۬>5�mٮ~�7�?5�pk���v��s�p�9�j�Ӎi�,�${jf����W��Fr�Yu����e�̘w��Y\є���u��Ө��������=0y�������-ޔ	O3����^�h>�8kl�R��h�rMnAF��xr��|����r�U1�`gk������s>A��t�n�o*vɢu�A�u|D�\������O�qǠK1L�7lG�f�&F��fff ��j��W���n]XwVw�CL��� �h��cI�q15�
 �XÛ�W<׬�r��4\��ƽ����i��7�ݱ�J��k���pJ;3<_n3o�$K�������Fd���ъC4�h�Zr!�7�@l�w�5�=�Vܱ;y�����r��[K*��I�
�]T��D��0�� *On%�p��b8{�mtև���nMs���Y�hŇ�Y.�Q�ڕE�+��뢸]����;ӊ���\�9B�/8^��,�Z������]:�"�bc��IC}=/��[֏����7u,5c���ԋT�c��i{�������{����$�7� ��ck��M�z�6_N#D��v����x��&��=Z4,b��r��(w�dW�"�5��Dj�;�b���RP��f?D���N�OS�&j�/a���{ꡇ��o��Ec�q��)�BxeŖώ�W<��[@��?v�Y���
�e���d��,0��P.�# Rr0�yw���3*Q�"�L�5�wCիGUջ����u����K��\�A5O��[/Q�}��fRY.�$��SPpۧs�&�h�3��+��[�*{�0J��Y5ĺm�
ӒZ[;k��̴�,��J���=�:����|T��kg�������SYk���K|�~t<F��G��R�]���u/������@uޡ�va���=Zc�p�]ͻE�:eNMD��(f�S+׳����y�a��^_v�W�L��
//#e�yg&S"�;d��`R���HO��d�5��C1�ճ�0���*,�P�=�],�:�iX=�(+ڋ� ���U��l?��A���+�B�H�&x�v�c�s`�m◙�[U�W@|P�U��S��	�J��㾵�òӢ�
@{����҆�l��wG�/7 Ư�y :š:�����Up�ȺZq�l����g�m�Xg9�p)���t�j��7\Ǿ��A1�]���׉�/إ�n1�Q
_\<�FZٌ��+5	g̴���+��;�k���FS��1���4Dk�4����W��U�X{��t�0 6-�Zb�&�{W1�km��xl/�w���&Q���wR���k}�O�kh̗��s[,U�}&I�+.	��XK<7'���W1�X��ߟe��p�� �(�0c��K*e��Jz%��Mz�\�Pu����'������)��i��g]��
��
8����9z�8dړ0)Q��¡��$6qm�!�:���@̊��y�V�Tt>�͵x��Q�ҕ��MxB��S��cFPfG\uru}���I2<&<�a_�{�v\��"���Y�OM ��`o�����9�P�qP'{Mw6���׻D}11�a}�^=(-��S�mO|sNy�1B�ܻ7�[\k�ȫ���V�}���M��2��r�������O��j/zsҲ�Y�1�Xtv��w�\Iz$�v;����*J2����&*ġ���1ՓzP�04�^*��,t#(�.��jM&#���r�9�q5�3�����{���(c7H�9�|<\��*�|ܾ���~#[J��鞑H���co�tJ���?j�̝�֨�6����_��;gG�T���oP׵����o�s�C���gTP��D�N�(!���k�!�A�t�;P
�7r{Gd�6����S��/5���ip67�H�'
�p��q�_���]�H�յ"v��|�'r�K��ɹ���,��W�H^�f��Qu��s����.1��8����8Ϸ�'��)��8�m�_���f"��Q{4:il��Aڧv59�E*�b��L�
�m;f�;\��)B�R{i̥�㗴8����N#bRZ�ڱ���<��w��W ��Z <��,�ԑ4�Ѻ}0��Ֆ��Ĭu�L�;�t�4$���)+��jMZ#�Y���Md<��4]Y��Ȏ�嫇�J���3r��x�A,�Dw7LA10҉�6���;����0�;�ɷ�.��>�n��Z�!{�E�"V�,tSz12hJ��}�0Э��S+��[nR�[]aG��R�*��f.�O���z,B��mQ3�G]�o��M����nݐe��Sv�t)u
Vk�m` �9hwt�f�� �9x(:����|7�XxE�]�d�R����;*L�H{�νٲ�ۻ).D��f��}L[�2�Q*u1�C����9\�&��]�M���զR[�Owvb��6E뺝��g@'�5.�Ӓኦ<O(U����}�1�kyj}-a�M��w
.\J�nZNa��q�+���ɮX��4��_4��X�u�v�r��Wm<��K<�]N��S<*lCUCa�+¨���۳���gx؂T�yjs��BP��m��=�ݯ�f��}&�7#���]����&p�!P�Ӫ�T,*z'��l���ܗ4_�ZR#T{h(�t2^-v��0-�3�5�u�;������;�*��U��(�e;0����n�{w�|H��[&�`�J�pL��Y�q^]��r�Sxu�����!)]��K>�솅y�v�U����}��k@�,�r�Qc�yn�̇��w����ĕ�Y�ԗkF�-�D�mW8+sɒ��˨�lv"��X�
Wۉ@�����޻����bU�k6�E.R
��ʤD��{ܙ5�e;�FK1�7�W&xi��V�b�g5n��F�\����c�:�Z��ڰ�T]���s�N��{W�������Y�eh/d�e=����-S�ڍ��Ѭ�)ep{(X�V�U���${����si۝s��㏧T��lF�I̫�V(o^G�`���4���yh�t�nd�Ŕ��p��Vެk�i��9�f��Q�[k�W�o@��hp��J�l�v����"�囕ĕ�l��2�
���+p�Ԥ��kY��P���0�p7s%�,k�� �G�Hz�gSb�2�Å���Re�*���9N�ay���j����Oc�Γ'°t�Szv#���׹O�#
p˺��V�˺I�BwZ{��n��v�
y�ib��ܻnjՓ�Z�JGJ��v�p�u.�4�s�0�4�r��fRt�6��\�]��3��V���7]BZ�y�ӣ��o|rM�$�h���сu�ԑ�9���gAdW({^��'m�Vu��q!���F])�kNæ���c1���tpN위i����8�%p�_=GsLp���xJ"��}z�Z �ubn�Tu�yS����l�4�5�4�}m��;�n�T�Dz��rםW++@lM,�m�{f�ڏ+9È!`�KcG���:8�ȶ�(&*b6��l����ҍc�UAJ�ҋ+A%��T��5�Ķ-(�0���Z(��p�B����+��d\j�Z�e31�J�(�!r�fH9f\�j�֋UQVS-J��fJ�6�
�W3��mX��0l�1%���Z�h����Ymr��cTk[���Eŵ�eJ�m��E�kh��-m�*
���s�51s��
��b,Y22�Jµ�jQq�SF��L�5�&d��J�2�kE��U�%�[mJʬ1�&0(�R
cU-���U\X�����n8��1�Sj�kR)Um3-E�r�rY[h�[nflR�E��Z���j5R���Ta[V��l��z6�̇$ "z�(�ʛʦ��U+yǇ��v������tf�JH�ḭٕ���+�w-ar�ͳ��v@e�C�U*3�5N�f�FI��� �+�8�@�<^ڄ\4�f7@�qC{��G��;&^߾��k��T��9c�Sܑ	Co�;Eܙ�K�R<M��T}\�����)8s���m���Ŏ�H_����t�
"^b�zO�,s$�P�,C�{L���k�q �f�z��>���0\�3�~��#o����3�����
6�דb�;�o��ޓ���|}H��S���l1PT�Ʉ!J͸��򝳰TkϤ�S�D���3��E��6�`XD�N�s�����(S�uD����6!���u�0ȋq���J���u����dU�m@�&���p���\j��_l��Y���m�d��,^���(B�vY����i�;�6�e����O9<I���u�_�~���p�-*%�{�>3&k7U�Iɱ7fх��--����a�sU#fH�F٩(k��1��IwUd��{.��{�~^wy�a�By�	̨	��!y:EC7E�S�!�HC%+ܼ|ϴ�Q֨��Y���#�<�ޱ�b�*�G�%�mII�y�0W<�!Ө�.�ʱ�*��si6����=�$�ʓ�d�W|£@��d�thh]�~|�0��\��Ǯ�\+���7��[\H3O l.�_T��V�=�R��#j3���ے��.7��(o9�z8����'Y_�˹ns+�3�;z�T��4q���>���/R�&��Y퓬�C=\I'�b�����_^R�w��!.E���A��\M��tе4�s�*<L�B.KE<)h7��];Յ���f�l�g��P�/ԛ�o{��jy������\/<�s�]Ix_/	��J�됕�ͣ�)�U+:2a
��LFe*ú�{�CbdUf��]a�:���_LJEӕ�)S��Q�Ա�J�Cc���=ˌ�]\~�e�&�[�\��^=V�.r��*scHOL�E�q�X��ô]-8�J�8:&e<��0���=�����@p���஝B��h�Q�aa�R���"ǯӅ;�[kރB'�&�#�����V7��h$N��Kqu����^%�9B.�P
���	.��u38�q��l$p4����U�\>����� ,%���6U�҅r�Z���Ĺl�y6���|�Co���q�'"��by@��"����Ձ�����W�o���{���}m$T�e�5��e����]�y��s����jj*�a��gb5����+rv��wP�EB[�;a}���E;&꣢�N����dw�M���]�MD����C�Oޥ���p�lCp��H|!���W��7^�sχ2�S�/&"=Cz�k�.�h�'1xo�˳���رn�+�Hd�T߈�,"T����/o}�W�.�LH�r��8-S����dU.����Y���T��iZ�j1]�����7ji:){�c��c]E�b�d���T�\' F@�'8i�s�[K:��V�d�~�$�n
�R֌�p��.A�]K�u��K�{�p��owf��)�眕a�`��+�e\_=��J�R�ܪc��Mp���2�\���K{��VI�˭L��!�5~TV��tLc���~kJ�i6{>Nx�ī�����n�ԡ�Y���X��L>ʌ�a�:+�]"e_�����X����H���U~$���H�k\���h��I�*��W^��UB����s�2�����K'G@x��Q�m��i�⽴���E�@^��8Ur��Zx�S��%z�Ot�*��i�n�sU���;�!*B�ĕK�/g���$����jα�O&�E|���F�_�7�,.��\J>^���b79����M�=N���lN��@i�	V��d��n�ֲb��z\f���,��b��6�M*=d�j:���L�=��ǆ�e�m��9�.=��7k-�����F3��<�p&+�3�['\�
_\<�e��`�ݍi���_��w�O	���OԴ}��\jU
�1DrEU�|�P����0� Ȝ#�mFp��ܮ��^+�(Yͮτ���C[P��p��zx�Ή�R�u�k�S���i?c��o��\�XU�DRs����6��\���Ey9(��(p�0c���NV�m*ϳ{����;04�����;�Co�ȿS��ͧq�m=4�����L�mN�����w�^uCt��K���J13^8����Y�;Zo�ѡ<kjV����'4�/ν�e��W�0_%A�%�m�O���a�w˶5�bC=��G��^��2�'p��w9�z���#���z6������U��2�=X���L��
��V�n�_q���yd�hvh}��\x���8�Z,h6�U#�|�|<\��/�'do3��c���'���/ٗ�пE@N
Ţs'ORg�y�hu�f4F�<�p8}ʽ�Y-}8`!&��p@���O�����l_ �	}�ÐYV��f<��U��#Hd�f��)R_%���%���c0�fj��}*w�{1�:�)U��w��܁Α�ɜc�A�%�F��޺ӵn�YK�lt!�[�j���Qy�;�]9"ሞ��A��b�]@�*&�v�\3a<��H�lE�}"θ:rkwZ���U��{��[VJ��X�>�="��B����Nu%�7��ES�Ӣg���Ϝ���8\�/Q�|Q��׆LO��:"��X�:�ki�c���Jp���X���ƻ{��}�����%��5M�#�nl�onPv�ݍU�Mf��u�^��SGEc����@�bm�n6dUz���(/0H�"�ux�p�Y�tؗU��x\�咐f_UpB�K��i�Zz��ک�H��������1���j��4��^�T���f��N���� ��/��C��O��Q/1~='�x�9�����Z�~�C�}#)��U�2���B�K�h�Ⱦ��획�Bwr���;�n9s�����IF�	���z�PD�Q��S�'"�)odL�|�,�*0%���i�L���.��e_��@*�c�ؘ�\�����ʖ؉U���l}u�E�!o��//1�L����O;��M^�ת��׹�,��A�q�Ԡ宨z�Y>����ʏ8ΰ)*���E�e�1Q�k��kA�ᤷ@�e-˻깻�*��V���2eЫ{ss��"M�ĭ��c�غ��D�l�������ˢ�=�E��M�^�`�:�mp-I��Ŷp�|��N���왲�B�b��}orsV*�RR�6U��Zm\��n���{!��B�ïP����o���P�qrh��J����W�sl���i�7Cb��P��F̑FQؒ��E���M���-{�<
�����<��%���'���#�{��49].6�Hr���\�ж�Z�St����h�*⥇Qw���"���&�8����x�?J��Ω�w1('<��������ݡ�Y6vr>_9p?+^�E�&��z��'Y.��Đkҁ.�v���]/{�6����<w�(h��Ǜv<j<��I�}iw��f�g��v�xHf4�4d���7�0]K�.p�1m$�+}�?(~��[�L�3���U�R�@�k����7�BS��C�C�ۦ9̺87Ȱ�[t�fR��!>�lL���K5u���P��{��2�}2U�m�;
6nLl
��5<#���v�+
�:�1���h䁬gu̞;d�)[�����L��FЛ���H��qX���İ^��ۺ9F�J=�-��+ޤ+����ͷ�o�K)�z��5�*�
ΰ�c3���7���jw��/�(��!%�����z2���/�ur��њ�sN��^-�(��I97������@Mt��	إ���L4�<�J�{��T;����I�T���P�w�Nvhuɞ
��+-6#��x�Q�To����|�%z��h�ӔE�=�����A"t�^���.�R���O�]w|f�ʸ׽��@���#��/,�f�f��=�L��v�|D��S�뭣������|�K���Ú����Z=P�+�qM��Y+��dq�ۊ��<�%�㲂qӜ�%�>H���+7�ۻP�Ƹޮ�pZ�5o��-9��pܻ;y-��)�,���'��6�4�)�|�571Z!Ip�1p�t�c��>�x��cÛt�C"��|ndS�.���[S�j�§|��,�A^I/T��<"j&X�40uE�;6.3d�\Xa_��P.�# rp�]"`�d~�=�c�z��?{��	�z˥�%%.A�e�@��M�6{+�K����*&�px ��nʸ�{S�B�Xj\���T�
��z��f"+�q&�tX�V�S�֛w���)��z��w4��x7$�-�y���M�Iv�ڞ#�_�4���[ʍٽ�&t�:�ZI ���s��B���`�u���WbkM�w����X��vT5z��@Bv:���YТ�(i�V�⥊��ӧ��;�./��L_v�ݢN"�z��(z�w�#s�l3}�;b��޺/����޳N�̰}�.wot͢��<"g���'c�%����+\�"���ޟ�������+[��~�]�מpp�ڧ��3f�w�2��E�N��]���sVC��~�Z�S=�W����q�U}B��Gq��Me8}cg=�܇r��za�yJ���p���2`��-Ϣ��a�T�{Ư�Mƺb)K�$��T��56�;����+�p*�W�3[��5�*��Q�U~�7�09�Ļ���&���NnCi�V��%�ThbԾ�3��ǃ��=��<t(\�P�RDx���i�Uo����w�ba�g�
�T���邇Ӆ'��u�l�DE�5�N��!��ȵ�39���o�M*��D%��XZ�/jش�}=l����ơ�����U�۝FW��-�uOWF٢�K	���W	�#]���������o����hc�욹Un�0'-�ֺ�b���V�\���P�r���
��_T�Z��3(R�p赆���Ix׺iy�(M_*:�<��̹��.�n��䡖��Ksuw\�ݽ��ùne	õ p7��Ԣ-�K��w,R�H�7x�w�u>ZDo�����B�!����d�N�%�K2�'�S԰�;��?e=ώN6=��,�쫷�ۓ�-���r� ��o$M^�����G���5լ �f�sW�5T@�x2s{���&)�g�VsX��?j'���}�С�m�jj��~��=bj���ZP����/"�=�q&���4,:*y8��㜁�٠ũ�f��vI��c5��:�4Z��y��Kmys�Ah�)�]�5+k)'j�6�΀��הE3b,3.�딾<Ð�~�w{L"��82�&j��6F��p/T芎�厸��#��C��n^��>�L�~�5J}�/�cA?��8Q���u1?Vp{�O�<���[M�����U�#��r�mp�`ydZzc�Q�~P/j�F����ٽ�Aũ��ڔ]�y}�y\�SY�pP�B�G�����c�EW�>ki
�y�G�ux/���y��{]$���tip�2�����,Zj���t���=�M	CI�/bLú�K �R�պ�^-;�۲��\5҃S]6�� ���5�JhY��+:�M7Q��.���;�Y}"��i'��S�ȇCi`A�<{��]6,���M6d�{��|lg>��4+vSbu�8�di�/�nmԗd�~=��Δ|�����ĝT�ת�3[,߳�|X�.��C�>���.^b�I�r��9K����YP�o˾�2������U8�Uq��_>�����<=Ol�n�bK���ܧ���8mL�e�+���n$��֪�ve>�&?�u�5�[7�b� ��Įi��7KΒ"^UL
��N�x=������PyR��N�[[2�T���34u�\2���x��v��A�-I�1m���\�������i�b�O7k���-��`Pˣca�+M¹coβ�B��LG9<�k7v�͝g+���P@=p����!�r��kU�9f�ꖜ��hl\9�6�]�ْ!�;�=F�^��y�(�/@�~:�3Hvx��I5�X��'T�_���bӠ41RXth�Ĺ�浲���޸x[ywB����Yb�=u�g Ŝ����ҡ��u �Bɽ��$��Q�ͥ=u��i���+�0���q�IJ�V���O�V���.=x�E`�T��������͟ݚ�D�mӵ�t�A�Un^t+�8�V�	9�b��W*֏���R�)�AVR���TꝌ#�AH>��ܒ�祿�ۃd6�6���!�~	�W E<8wG�g*m���]�VX�%��J���Z�y�'|��I����7{� a�#\ur�e=�<m|o�6�Qr\�������eA�;48����iZ���c�d˞V�B̘�m6�V⥈,z�!��[x����z4f7y��=��\���ΩGUB�N;!���<o�τ��["V�a���������R���@p^�ͳ[�)D��|���Ab��n�2]��8-�Y�͂7�F7\:��Fa�n���ν�nh;�re��虠��<�њ�e���n=���*����v+�K�N��i8����cV�ۼ����]�*e�=Svu����쎵̻e:]��LŸo����n2�䞐�U�TR�a=,ުd��{�[
�T�Yтȡ0֍	d�z����YO�U��3yg1��'0���:��օ�>9@'�m��ڛ�]�i*��5FJP"6��yVn�PP�]�|č{��.YA���60�٧�X�R��6�l�6�u
iu.����V3>];�;�jG^�;ә���i�,�2n!HJ*��w��-ī_��.�P��8��5ͅ6���SFȋd�74-�)�wag�T09�Ȅ�7�rF&�	�U!_Os�A�����&�D~F��2�y�c4�>�R-��7m�i#j�w��
��N�tұ5V�EY���%`�\���g<^�{��N-7�b:��5��6�.i4Ă��ŕ�ms��=�p�2�⣽�]�,SeI�v�/K5��hW��Bܭ��{JT���)�s: ���o�R��8NH]S[s�����ap�E��7:��nkan6��2�Q�\�M��E�����>ko(KZ�%�oT��Wù�*�>l����*ȏtpӆ�6��f�����'&��c��ֳ5�Uf�:��m^P.��$�Y���4����V��Y��ڊ*{ְ�V;�j ���*:�7ya�zқB��d�k]�����S-�Zit����l�������\���:�1nV;8b:��6`�,c9�Ʃ+�����f%upA0=�k�.�X����|Z�&(�U2mqۘ�-@u���w�J�r�pM�d�����B|Vڮ�'�U�̱OuGN��Yp�<��Uؘ�a�չ3����2�A��&¨����2��#��ڄ�Ӱ��h�b�Lo�����T�+啕�������k�(������u��b��V撆�G'�1'Q�nm)�0��R'>�^��21�G��;��tټ��`4��B���.�y�绮���fn�-�b�G4��1���k0��yͻ}��D�2�f���m� ����<ڼ|z�WJC��R�2�L���EVe�J�խf%ETpŬV��*YAm����E����ٍʈ��J6�Zն�̳C.J�Ek+�!kJ%bԬZ��ѭKV-��h.ee��,�J%m��©ch��Q1�J�[B�[)���ƣV6-m��UkK�a����J�U�*�s0�bъ�iB����f
�-j���*ڲ�ܥZT��ɕEm��(�YJ���.[m5�q����E�ĴQ�QA��ņ89m���	F�T��������Z[�0��r�b!KR��b��Km�nZ"e+m�AL*[Z+#�X�D�ڱ�b�VD�Q6�iX�m���*)[m�mJ��ZUT������m�V�,B�����2����׺����˩/
��t���w[$���ҋiqrr#���@����S�in$��׺��0â�nC��q��+��X��N"q\��*�{���y��Q�C|���A'�_mw�jf�3��t\6��{
����K�{_E����m$S87^u��i���b���Q�����y{������m΀�B���C��gF"��1�J�n��tm��n�ƹ�{�w^^-��0��QQ14�3�<#��UHo�]-9��5��_Ȉ��)�Y������{^�u��:�gE"GN@��`
��	q��o�"�i|
�b��XSZ�.���8�,=��*J%����Xi���uU�D��0�߱H
�>�YRF�t���=�H��mȝ����=�-a�H�0�A e 2�]"�l�����;��Q�/c����V�ލjt�^b�%�W�3��L��v�������-�P��ݗ�W��#$ш�Rk�_�_�Q�ܫ5�+�ߔ��)��I O�KN����u/H̉�bwƍ���;�:zn*cV�u�E�9��~n]��ylX�Y�L^������Y��8�훩�%hƸ�����J�NsB��v�Y]#MVK�<��.���v����/L��=%�_0��V3��Z[�������˫��9��'YJ���t��p���Wh`�yO9H�]��i˝����2��M��~��]L5�6bب�:rkpZ�=+��U/���N��#l��˺��j���\�fUb���48)���c\^8���,׸�¸��	UTv�c���ßFP�/��Yw!�%�򂰖tf%.�f_$
�j2Uݠ����Z�b�3��	+��J W9+��\sɛ0�J�R�ܪcz,�#f�j�ro������������U�q�����&��>�{q"�֍��q�@�ϥ���:(���${�+�ꡋ�2_LZ;8:)k�M���,`�Q�t���S���T��	�[�ۉ�wz�f���8�<2c~�,஧�UB�Tf�
eV�1�v����[�S�ĺTY���L����#��V�&"�["����+�S�t���rt��ԫoג̆ڞ5٬��i�-�c��.���.x�-���Ƨ�~�LA�D��3��b��f+�z/�9��}��c�C���������c���1�߁Ӣ���5��
�h�c|di����q+	㒓_��,������u�5e�l��n�&��֮�s�����s�p��hsw�=\�R5�ʉװBmV��y^��ns��B��R�Ѿ�t�m�l��}�4��TY�)g*�"�U���$97x����*Ҵ{��/f��]u�mԝF�/Х�������kjǜ�G�|.L#�#Ǟ��n��EZ���y}�Uq9Ň���b��"���7	�Cm�\���EG���n��eS��W%V�5�ݪ���(k��`3�n�qZw�t1o�H�S����;��i�4�z'1�G��}2��ـ�\���r���
#z��6�Vz-�x�v>�(�7~��)�Jo��#�R��n
�p�����MD��&X�0ʝ'Z��ᬇi���rp��?!b���R���o��v(WӲ�B�������1�:����yҩ5*7[���IܑL�:ÚF���,1�m����t�B��>q�ۿYbՉ�Y�]�D�N�3��hb��ͺrzN%i�r׋�A�S&�>#�f�.)�,n�k|�k��ݗEW}x�F����
��QQ4���i��`h�yDV���"�m���:��1�dZ��f�HegW��ip;�l�({�<��<N����9�i��z�����s�ݖ�<��L�ޢ��,�E��45:;���+ٵq��<�<�"݊�u��!���^�Y�´�nC�Uh؟ξ��L�%�W��ChQ�׏�ل
ME�vDb�Gn��N�FU���Y�l�,�K3��8n��=W��	���5NyX���9�����#{u��N�#Of]զ��7s;Ӫ^ͺ��3en��b�Y�5�,K��*�~��bchJ�^��Z@����{:��aZ&���l�~����c;��{��lwn6dUz�5��F �1_8��5�y�9s�`%��Ova�XA�K�����U�at��Շff-�9x�lY�q��5y8&Y*D9�hD��x�u����R����S�.̰K�i�}�y�rZ��]�|��r����~�P#��W��|��Z,r7��x{-5�3/1��;u���7F�޻�B$(��2B�͎�%[?���Z��¹>ͺE��X�[{��u��N�q��O���m�j�h4���0�z���p�4*Xyu�{~���M���4�ފg�/���U�yCڃ&9	�jOaةp��mv�+Q|N��7|J�H�w��Ûހ��������)���;�p�=d
[�t�a��Q�����=D���r,A��Uγ9�咬i`ꝩy�3;,�ֺQ��Ӧ�}���ҽ��z�X���e�O]��H:e����>k6@����K���c3UEH+o��wʞ�q�z!p�jv��V����qd5�2��l]����N���2�I��d��f� Y*�B���P�Rt��4�(s=g��\k��laD
�/��O�����%�s�1��r\Z����.���$��,B�T�\'#���t��hh>L<o�nݨS�Xp=��%_ *T8d7��&Ku�<`��h���N�@�0�|�(s�Է9:����'4�-���~	���Q*}ys9��Y���XoEz�ě�RcmE֦N.��*�ZG9k^u��{��W�*�f�������g��>��OS��Z����u�`Z�.(�m$'��ߔ5�����/�j�m!2�7�5���R;t�*�,n�����]�#qQ�\�U;:2!5�m�V]>v3�{^�[z\(#s��C;�:{ےh��J�_�Q����\�hG#]J��K��e�ܷl{b[�2����%*.j�t�%�A �0�d��5��8$b���K�h�ZT�̽}w���e]i�47�j81��Q������DV�J~`s�/q"��C8���ŵO��;�#��<��ޝ��kP^�0*��e�,w��fU� �g^!j��sn�q�}�zn�eB0��H�v�푡�ɻݓf��*M"ud�O�Uq����t�T��X�]ns�B�giC�$�$u��ƃ:݈y.HCJ�7sDJ�f�N.9�s����bމ[Ӑ֚�eц(�����Ӈ�O�x�^J��R[f�Ll������WR!w=G��~�����ȟE��3GK��|D���A	�Fʻ`�dn�no�9�:Z���,,�Z=Kz�?;t�۹�\�T=���$1\YX���t��qo�&�5H�^������',bP]h�i��Ӑ�z���|l���\ia���xH�Aq�>�p�)�@�'�s:!I��lT*��^�=�*�BPT`�n]��+�;i����(�E��:�_�f����/Ţ��.�5��	W�׏<;R���Q	�#��h��Ԙ��W�g���^���*��Yt��c����R��0<K�q���3���+��*�LR Rq(Q�@�O*��#�8c��T����W1��*�9�ޒ.�ٖ7���)��:wR�"�V�vV�|���{q"�֍�h��qj�h^�&� g��IzM|��-�7���[��~ÔTgLc=���Z�x�������v.�dk���85衬���l�N�+�{-�#C��>~�,�V���%~bDw+5�X�ΫLV�ٌ�n��h�#ǯ����#�S���к啂m�f�)s]<޷�JJ�9��ۮ ������
��sF����-��v� {��׫3���1�隱�/Wk�f&��Z�D�3�����o�,`�3�s����c���X�]����M��V!ʴ8�:/Ϧ8����a�/,�<���D���mh�Z�z�p������K>I����
���{�F��b��JF��\��]AUt�@��-���R�T]�fl�t�u��m�g��k9�����6�ُ�XP���#�4������u!�s<b�˝3�e%�l�F�1���G.��1�-d��L�!���z�S��7w1��kS��ؑ�Q�;H��r�܍v�T���9��P���Q�y���s�r�^���ҍ�0l!^0c���R밎)�F)o4<��E[��J�z�:[�Q�8�q�X��9S�v�S0RQ ����B&*=_!�������秬s�Y��^9N/	q:+��95�kUđ[~���X��C�����插\���@[�:N����� *�9���}sJI�~,:.ùb*�T+���!Bq~J����3q�^>�7hs��e�0KA�����)��]bŁ�n8�Wf�$M'ٳ-�ڍ�	��N��g��b����_Ĉ[�[�m���Zy\�"<bL�z��9�e���Q�u�e�bk�k�DK�q��s�sb:f@�w��r�����Aڨ�\�17Y�ru{[�Zr\<^J�=MM˝T=�����ё	�֑pXcjUb���R��c�D7�!#�]�7*���$�K8r���f�EP�����TG5�u8��s�3`�4�2lýٶ�
��cz���Zѷ{�ET����NEE��3��h�f��&�TTMy'n�a7���b9CN[��2�����{X�!�jİ<ͭ���׀U����`״��f+��YX��00�фz���7W�a�}��Yױ	�ư��UX=6��,���Ƚ���E�ʞ�N9ҿ;�Y|���S'D'�I��U�ny\oN	�Ǩ�*�ئ��¬��7���@A��94V�v�zUr�7D?m�n���s�=���=�L��cL�^�-pQq,�>w{����yv��Uר�x��n6�J��c:]FM���n�]��$h���К��ɧ�]4�[��v�����EU�k)R��|K���}} b�|XE����O�n�̛�*9�"��I^);g"�V!��~^��Dvzep5��È�{֟\��n= m�u��f9�N텵 *�-leN>�8C^�;�͌�ي�]n���_<�{��z����4�9�{��V	Ķs[qQP��ڨ2�̋E]�L
ݐ�.�Ɍ�䀾Ը�s��z60�+z�����oI CY3.�p�-z!k9��0^f�L�<����l�k��囂���3�2��21�iИ�p�˻��\��-Ǭ%�ߧ5�~��y����.�4vݰa�P ����ʢ��3�,V�{��`]hK�@
~u<�N�㘽P;���om�yw7��Hu���A�.%A�j��a��lu0k�1�_r{wj5���^�«B.���P�5~YL]�:�!�jۘ�����}���gy�Z�:�l�!(U�:ky�T�0���--����1���Z�۾���ö�w�޾"�W2G��>�d���uIx�$��R�+���r8�=0�N���y3�.n�N�08�tx3s$��H���Rd��oō��4K���&�h	��$mK��X�虥C���d7#MByw"��p��p�}Y���(g�f��󐖉ұ�l���9m��&�(�ᒀ�nYX7��_o�Xv�����T1�R;��4�/x����=��N�q�h8ڛc��4TykG,���ox;���*j��[�e���O˾���&J앁�ŬmS��t�#sy-l���M���<�t���c%��
^���_�+;���s�N{S�IE�ᦇ-s].�Πo��2[�Z�S�J�X�ꁣ�l��>c�|�ŋ�A���cj��M��om-Uh��|�s���WA��݄�J�~ڍ1�N��TTe��.�E�K��?
�|�f���oCI#4���,}�	9z�K<d��a/��T�z��A���B9�Whqr���c���+b�f�i�.r�zښ2����j,��,�eN@��`
�� o�`��asԓVǥ��:H�M��:'y-0h6tm�*��z	�{�MA���
��C�S!���sU�N찳#["�V�nI���O1c��lx;ڨx�C���Pf�h8}t����.��F�����^r��0��Z��x�kk����xxr'�WL�e��lG�@_�M^�����r|�{�b׿
s�f�}�^)�v=��z�o�ȸv�a�����N{F@�:g*'���Z�:H��a3�|&��;:cV�Z4Zj�4�;�gm�1@����'�G�D����t����d�9,GI�m�0����<�R��,������D����Ѡ��z�mF;�Eq�yM*�1*�!�~;J�k��2����W�����$
�!�����KE��bKΫ,Z4�qK��a���5�Y�,��X*X L[���l;�_X���G2���]��zl��J4�a���WZ�hM���hz��x iR�MH@Kk�V���m	F��lѤ5�d�5|�k/^�.*�!��{����k~�Vѝ+jp��]ז-��X�ҴV��r�*]�rN$��"�IW.�
7tL��p�իE-�gF�b��VpoU�[���R�h�wӤ��O@�n�DV�<��'X%jỡ�wa��7+�תѩ��&큯/�[rA�4�f�3	@AEf�ڱ���)3�12����F)�c�~���1x%E��w)\"o�;�[\�)E,d���q��)�1�޷R7��!�sTo�.k^w'K�UfQJ����'����o����{�҉�m
8�5�Gq��a��h�4�n��lH�6�}�Or#6���΂��Zu��/��d�Q�+.p�g�f�٥�J�?^��w����Ecѡ�ڈ�d�qKd��f<M6$�i3%��g����ڥ%Tr(}�h�����-I�qϡ�u��vF8fI���:��D�sc!*$]��r�b�ĵ;�]��x~��S{���#j�mm	]H`pAH����b&��[�f'/Ga��:��z��2q� �W���S��D�Hu
��<�B�Z�k�<�J^" wu-�X�ĘݾV�u!ƇJ�����2��V��J��S�����b�,>����>�cx�v(�]W0�R�$���.���.�Oy!Ċ�rV� c��o�4�lid�wNM$�${a�.rf���q�H����v]��{ʄ/�֫��4i��r�a���[�U���[\��b@��Z&�Q������'v�#�sB����0��K4�>dT���̑��BC��mJHa͙T��-�wY���n��;���gad˷"m#.�DDml
��OZ	XF�d��յ��"4�*����໩��y��s��Y�J�o)�ձG���)�x �O���ye/A���!�x ��ZOh��(�3��t$��6ȩ§��u��ҵpΜ�m�9{��YТx�0{8w^��YÖ��K����1��DGՙe\I�k \�� ��h,�4��������2��5��\Ơ_U�/�j�n��0;/F�[���H�Z,f�<�d�����2J�Â����X�+f�Q�o���aw����3o�\�"�v�YsM!w�mԥ��TMX*�&@�)�IzOza�q�и�#�{h3�t�tT�dr�З%c�
�3w�t*^G�Nǝ4Is�a���G�E�񅉼�����Ǔ���u���C�enQ[��x(v�m:�wNJ�A�'�\�լU��ӧ�}�,l�]N�ˊ����V���^ε�'a��[�~�o��}L�B�E+b�B��VҌV1[j*֌Q�����Xa�k[IUQJ%�e"��Kj�mB�[miE-�ER�L�ʢ�RѶ��QV\j�(�����q��� �ʶ�B�+iE��F2ڌF0��PRհ�e1q�ʔQ�l��X�a��m��űml�Ѳ�*#S3�-�+Rڊ(���Z��Y1��e�UQJ�JִF.[iaZ#���eTT�[e�(�������je��b��m
����2fZ����jen(̸&G-V��ei�cr���؍��UUPAETD�V*%J"%��q�cQY�Jض�TJ��H�2��h.%F��a�̆`�Z��P�`��R�KmJ�kmZ�#r�(��aq���n+(Ѳ�
���kh�*[F��E)S-C�[��aZʢ+��6�UF�kJV�+�F�а��h��YP����1+�bZLa�!�-1DE�R-F�&%KZ���
5amU��R��dT�5��{~���z���eƩc��WI.N�e�!0��|a';W8E�x�)��V,�#�	�*�����b��\y3���o�@�OrԧT�8g�2��6@���N^�u�W���D�N��Z�юU7л<	��o�jٷ�];\��Y҆�}�R�LWC��@�N% +��@��yW!��^5R����eg��;e��\%I71E���b��9EY�:t�7ؚ�!�XN���j$g�ѷ���l���w�܃����39:�7�ڡ���ђ�Y�ppj�H�Ǵ�Ō�qUKKoy{��}P���$���-0H��4�b������vUE�z��p�Q0�Gg9I�]�v0�����Q�e���@�ע�%8�l2�,���u9?-`���;�����f���yO?bfni��ώ�l��n�vE-��cDV�9E�<��[ ;�˚����cm�S����/۴�2���2��d>t�Nن;n�����8ƽA�7�yc��jsݜ����� �	�Ӥױ��;ד���ֆ>��<���1���}
���K2����.����v�]Oq�j+��\D��j1Ks��*��i�����[?z".X�Z�){n�%=	���çP�H��3++x0����e�f�|[7,�Z=9�@�+{��8@q�.���-e4:���NP΢	*��/=���]4Ζ&S�H��^��`j|�E^��w#N�x�]-��ds�p<9SUJ��o\��6�E)]����x�r4W�4��	��LV~��P��]��﫥B2�e�QΙ���L9�b�̼��!{�ؤ���6_Jl�5�h�3��^!�P��C{_8���]�L�+���'�)93��}��bz-�W{)ק�"��Ȏ%�-/���k	�{�uy�@g�fuw�bX�(�Pk]����Y������\'�$�{��MD�����N�d_Tk�f�һ�Qh� i��!8*�aM#�<�Mi���dC�S�Tj��4��sm`VkM�i^Ur����p\ǢU�"��ґ�~�ch:*Bq+H�t�FC��o���S����Û�����\,=οmQ,�s�v�TFk��{TLN���b�l�Oqץ�*N��n��f�e+�8�x�����׋��b�w���9P��-��^qS�B�<V(�l`g�b;��S�8�����u1?�<)�����E�sU�Zy�f��)�E�t��-��]G�sa{���
����,J�6)�¬��/m��-�Ybi��lᱹ��#�c�ي�-�!�f=��.
_n��c��!�uu��$�I�Z�HU�8f��\ܭ����7#9��d=��1�CV��I��m�JIa�[�浆�'�ޖ����7LVb���=��yo(ͽrJ-i�yUov�+�	C`8�<Ƚ�Aڧv59��xgut�~�zd��q:š��7�����)j���W\���/���gK���S��{��`M�ê�0�^\��e|о���i�ؤzu�J߀����!.&$j,��ȣ~�`1^E�b�{b�����5�Eq�����n^�,`2��GNJK�������.�~��q^�8^�N槲�;-�Dk<��n�עͨ{ďa�����v&et���L�Y��;�9���KM�fCJt���R��,�z��;j�9���^p���W��E�II���5��d�;�v�*3�q���n\�j �S���j�^C�Vl<��ms�đ���]m[�r�-o�S�T�bw�Z�� �zbB�Ϲ�M�����ȆP�4�X�u��>̉���������E٠HZU:��5�Ki�[9æ/;�=��W�`����8���m���;��F�Գ��%ۿ0�r�𬅣�<�g�����U�RU�"kܥ�W�(V8��{8` �:�	����F�v"h-��S�l�2Y[��4\[W�%ˍ�Қ��Ȟ�;OUl�L�K���g��h|9���=h��l�þ��K_]k�Tǝ��Ȼ�^�f�K���&���zÔ�d�B	ә���2��F��ATP�+՚���c>�[D�H��C�Cr����I��a�77���������;��v)��*
�R�y��;���,'���J�^\L }9.��a�/i�Fi�1h�0�X���]�L	Ԭ�Tkθ��{gM�4�s�Vĸ~\v__�u�SEE�#��7�4>�۬
�XEB֬�ǵ�!9���VD��Ƣ�D8J�F<�Js6�g���˧j1���!�YU��#9xPˮ�]����܊U�t��m��"���t�K�(o[5�bc�2Z%�R�������b���}'���x	X�[�M�{��5�d��~��=���]ȳr���b��]O0�W����7�S7��)"�x��M>�׊�[ض�V���C�a�+��%��zh+�I��N�Ur�"5k��֛�6��F��Bj'K�l��m�C�C�1p�Jޜ�Zj�F�'��OiWg�j]��ɓ���Sl��I�>3��E��GR|�2i{s#V�L1�!B�Ҿ�۠��Ҕ��[4Y�W��e��A��y(ĊӧOZd�r2�]�G
X9Y;q���\�pۘOzƞ�Fp��{�,e�7X�яJv���E=|)r�"c7;&�dlt�u����y���rJ걝	X3^+�����T(km��7h�'����ע]˕��t�ݎw���\�v�a��������tu�k^��)�z�;-pw~�\��F�U&9���
��鲝1�x+W+��I�㌽�ɑ1�����#�[�t��
�X�,O5�����l�بVx��A�IV��h�ˍ�w�vj�D�o����tWՂ��<��|'4bK�!�~;J�V�kT2E$���u�w���M��a�(	��/��]��B;RK

�R���R�Q�S1�������z�fNEoF�H5��V�))8� �rRgz�,�p�J�/�-����(�{�����|,9OUf��s�nҁ#Tei7΀��{q!\�\��3Î�穎�ZpUF=��j	af�M[1W�P���*3�1���E-t��{Hqʡ�  yY��mL��՚���g���ȃ��^ 8g�����	VpWS�UE�~���Vcv�kr0Ȟ;�5�={6�&�^uC"�c�dzz!s�zd1r�_������E� ,|=n��F��I�*�ܳ���KJ3�L�s3HoeN�.��찉�@t�cXqڄHb�osFt�ܭ��bй��x�8ϼ������u@�ѽ��d�wv����7�ձ����:�.r�=U;<:�umL�3�݇��w/eG%茎�8��쩮Q)Z9�j�>����N���ӑm��݌`�fR6ϥ.z��&�齭�#�{�������ț�LEB��!kf1��hC��Y��,d
8"��M�qsN[ҫd�nʵ{�<MF)a��v�N�������Jޜ�Rù�1Wʊ���x��Ǯq%ѣr�6!�"9�Ur���R��t
-����9|%\st�DLi75}����7:G�i����(8T1�Q�1�밎)�GU�W �+`7����剾Y�荧�p���4��멁I�DP,r&�\&�w9��B�@���෋mW��]��E�+E8�h朇����s�o��T;}�0)sG�S��0�ʶ	��}�1S0�|!Wp�)��&sf�:��%Ύ�损5��\G�'v�HP�_���{�d.e7������%M�ZO(Y��U!YVX��SH�N��6�U]z��yB�OE�n��F�u{�S���ݨ�Ԏi����c𗈊r��9�٠���ZE�6�5&��qC�\|�Э樤`T�]�M����dlZ�+O,��J��8_c���Q���Ӛ�҉�<�׶"<.�ά/,:gβ��p뉩b�&�uΌ�\Oi�p�}��hj�0WHQC!iYqS����bV�B̎�D��V�Z0�pr��~�`aʇ��7�V�ڷ�Ei^�����Ow�����=m�=��)4�\�q+N���ٰ��D+���B`���t�U��<�;E��S�: 8nWC�)��;��k]jd�ĸ�V��nu�'���]�BVv5���f����k���}@N�o�}��s�t��=g)]a�����},W)ͅ����
��k��j��	tA��e���b@�>L�v����4�Bۤ§v59���=��y��~�4�cy�4���f��N���0j�8(�T�=��pdh3{P��T챞�u-7OOS�;j9�k�#�$�k��|6�{�he��QWf8Apb�5MY�Q�V���.a8�d� 1��.Wl���u{�~N�������5���Vۇ�DL�@js+�)�r�k�|^��[���Knu��!��Ⱦ��}���;�f�\������ߦet���L�Y����6k��/���=n��V��@p��������=��tHZ�r�]@F7*m���pgH�>ʶ�m�9&��qQ1�x�t���[���ClR쾡P����E��ٔ�m������nmY��v�#v�_+X�B벏6@�v��P�:��U��pd�jˀЇ��6�v���9QД���P4�lfƸ���c1%�WЯ�	<୧�\:j����{�C�{�'��Q���=hܵKu*F�2���9�pU�y[�³�'Wpҭ�V���HUH��GZ�u(w���8 1�9����l������߇#�PU�3}���x[�L)HVU�{Pp�n��%uM��6�/���b�L�)�Gjn��ة�~���P�d�'u����ֻ��.-�n�Ԟr�q&�"E�ю{����d�����a8X+���z2��o�k"��.|�C]�zM����y�ݼ�r���,�����W�����ϱޚ�X2j:/&�ؤ�Cns��*��j~��YvKx9;Ԙ�է���Rؽ/~�������������S-cJWU�7&^E��=�i���QW�Eer��u�ɡV�ݽ��3sݗK_;�|�q��Q���^mQx&���Q^�LW��ߞM��T^(h�-F!�g/~�,��fj�������_j[�" =�o��ʳDl�yY�E�u��+IY1�r]2BQ:(����c��y�Y8e%��x�Mȍӝ$��m�P��� �8K��Z���a�y�́څ^s��RFY���ڤ@h�F��nQ�q��nS}�]�t�^/��*�=g��#�\���i��f�p+g�4�j��͸M�eo�ʃҨ�e���b���W���w,��V^8t���"�[гo��Rt];V��kg�p�=L�A���@�'X���T��0����z��.b�EوL)]r�ط	>��ҽ��
�+^M}�nFsڵ��y�WW�{O�+jf�5�����ؒ���[!z��Y�n�&hS����x��������]+������z3�Q%j�;6���(O\���������'��Ox��'S�I����RN[=�	�ظt���:�l��4L�j%l�g0��,z������栛K��PJ^N;"�7�n��8C����*�dV��H��Ɂ֟|�����*e���~�t�8V7�d�tгO#�q��E`��F�!��#v�*(�r�ڷ�eց*�.���s��|�C!�@��T�K`��{7 �k8�dW{r��&1b�7�f��Վ�u�@�
��nI�By��m�8�]�j:s����������{���n xۗy�����>��&x�������:�QO�����j*P��;E��}{Y��Au=�IZ��E��(��{�$:�C��EE�j���#~6�7��_�)>ay1֓p�V̭9+x�V�� 졗��9�˭_Z�:��Sm���,ڄ���x�E�U�b���Q%\�y����[�O\k��&�=����jk-����m�̥zk.K��O����<(Fv�I�uSqв��E��$��[�)e�Է��M��J«ÇfeL-o�];���y����J��1^��{ƅ�z{�A��_���p�+�r�+C���9¼�f�$n�����i��P��i�O��:X,���,����y`k��-�m
s5����nO�VmL����u�X3�8�t�y�
T�
�V�������o�HIO�BH@��BH@�脐�$�$�	'�!$ I?��@�$�܄��$�$$�	'���$��BH@��	!I�IN��$����$��$�����$�$$�	'�!$ I?�	!I�@�$�؄��$�	!I���e5��\0ڵ�!�?���}���������


UQR {�����!o;�HUE*%J�QT��R*��CE�0
�-�C f� �	��za� ��wnt���lk(��T%X  �;���@e���el��J���
暦�R��
ژ �s3mU	kU�l��bk*�R��(ɑJ�
)�5
����Z�����(pP\k6�ѵ����I�+�ۋY�32ё����(2"�g,�l5E�Tkf�h��Py@P	 E<d2��OҘL�@`	�4  E<0R���	���i�C hsFLL LFi�#ɀFO��U4hM1M2d`	�i��A�4���0�ș242d��	OI4�T�G��i4��h  h=@re�S�����iM�l�4"�!��AY- @NEAAf�� DY��|c�G��C��,D�@X%���@M!X�n�Al�վ��V�2��6�@(*�7��T�����c�����;��"��������͚���sL��ɞ�﷚���Цڔ_�RX4c�ݛh�h����Pn����nЬ��6�����V���i<�[����<�@(e;ņӡ��B7Suh���7����*[n�;���,d����ONTēʖ�(S��i��XߦU��q�I���Qe���y���*6���k2�4��Yq��*�%�f�=L�,�Y�9[X��n��En���0e���4��;�[��Zúy�:�@b-����ja�,����2�#q:6f�����v�� ��Z����y.��ׄ�)$����#���F�_d��H�!�k!A���J�\E*�ʤ&���<RY��Gh��xy�ճ,�b��f�F0J�x V]�ֆ;3jU��NY�t,�j�l4��7Q���0?��Q�Z�r�5�沝�qe�q]Z���{j�5��.,�y��ݵ���A�3e�2�"�֦��E��X���kZ$��W��Ve�e)xP��}��'{���+�٤ݜ/1Q�G6����5p!WW��YL�6�+�����vRX+u��C�:tE
R���6���[I,�a���µKYu�B(��-w���\��Иu��R�f+KC�l����tȘ/
*��'�B��U5-��C���i2���7-V�n��t)��r�	��OJkfa"�B�V�O)
Ml�y��t�(2;��<8n��,���U�=�{���m7R���f/��y�&���x�&�ۮ��� �+,V36�@ےen��4 �$ʕ��.�o��VՉPٸ�Sɻ3u0V�B�	laJ�0��R
��]�������5�
V�X}�rJd!/wwn��Ȭ& o!�TJ�r,5�f�;���]% ���U;�3]j�1"}[D4�X��Y��ر�
�ƭC2��V�C)��p:5�%�f!�]��XrS�t�x^�4�����o��;c)_Z�Lqx02b�6s6�̺�����pT+$wC[�@� 6�ݱ��c��)�a$`5Ώ-&�wx���wj��h*h6�)���QzV���9�����PI�Yxy2/+Z�t�ح&�.�M0^b���3)��!��ր�TU�v���~:�-E�5f��ܱ�:ŋ6������F�qaP�2�6ê�(�ٻ�3^:�@�qO��.Gdٻ"��M�w�%Me��Nh�k���y��?��#\�#��<��KOn��º{Β��Z��ea�RqK���m�8�Ѧ���ڱ�H�[Dp���O[9�MhF���N�H��r��Hw���zE�Ȃ9e��4<��e��	t��u�4b��Sb�ʺҳc�����*�b�i���i ޅm%h��x�S?<eJ�5�[@V�����j�65�dU����I	�h�	6�K6�&(���U�w�-�CrSf�0Q��W(Ų�v�o�ie���Bf�)��D+d6l��L�W��`	2�Ic�vX�5*��Ɋ̬5�<��N���Ve ��Y�
�\�;7�n��lFj׌
�-UM,�#���r��3K

8U%V��:7a:?d��t�e�q�4�x�5�*+�R��v�A�ko��:*��r��Ա���iw��Oe��@bǛBb�#�$����ݷ�s��O����D��q6%'🣿 �C�LT~��FA���?M��Eэ�P�أܧP:` ��dt&��F ��*Xqcw033 ���T���̻���:�u�p������Gv#|[��K&��h�Υh>�&�n�Ju��ѬȖZ%�wE(M�H͍_D鏲]eo*�R�Їp��XE�f��<�Y��t�۔�%s�9��JL\1\�2,��ʉ:��mu�]��S����7����9J�g[�����<��Ζ�L��mw=7Y)6��U���A�[]j�;���i��;e�lY�y� R6]ed�^̜3"���m��`W:��������h"3�d�=V�����Q�]���B[ev��w�l�]�j��*j�1��_9G��7a����}7{r���lP�K�}���"�R@k܃��V]t�lZ]�]����;�4�t¶����5F��َ�R�m��J�!J��H��$��9fd�T������Z1��7	�Ƽ8�����J��
1Պ�e��t�z�%X���6L���X����w�#�坛-����V����^�*eM����^���˳�[#4�<�#���$X�7.�*���&t�*�Ӌ8�B,A&_FY�����	�EQ �p��nvi�v#'5*�9�ە��0=����w���S�+�tE"���m�e-n�5N��i�p@�]�
��v��j�:C��L�ܔ\;�%�d4�ֹ�儮=��g5�uѶ/;.r���W
�j4/B �9m��H]���_Lwd'MX��6��u�]V+^>��#�0�ɭ�dr���ɩ�n��1�8�!e�k����Pj}KLͱf\����ﵨ�sa���-����'P��c�2��f������n���$Oo���1��N8������#hu��Y���^�n�W`�wa^ˍSW1�#ۙWju�kH�W�V���Ls-��//!��B�tʌ�ɱZ�G�)�&�sa>�ŝ�n��ǘk��hH�i;]Q�i��%A�w�-͸��v�%I�4�h�غ&k�"1�Y�����E�<�����e����_��=Q˿�p���β�f�#�����w��!�u�����Ox��V�K!�aS[���!jN��mw��-�(��gnl	N��t	B-L��*ET{����:7�j	QŘkz��{%���+5ڶąЊ]�v1�s��l��HmnJ��:���(�I8ܓ����blr�w���8�|��9N��x�I$�I$�I$�I$��$�k�Ӑ���<q9�w#ۖ鴤���V{-�����v�����
IN6��k�RR9}Z�'z�����~�C�Wb�/8]ǣ�(R-���Յ�r<FgT6��w���ʅ=E)k��UԬ}�qf�b�)�i'}�8��y��nƝ��3G)[�Z��
@P�u�6̛�뺘��jH��u1VCr�_�˄�ں�;�Y|�L7Wl�h,��UحM���H!Hٴrv�?��8�3Vc��YH���ԟnjO�:5�u�=�Xظ��������΂�c;�ld��Cq��FZ*��n�K�+�2�/,�ݦ�uеS.9�7�zs�7̫�(;b��ې+��f�Tvr*-�݋�>�w�>�e����,� A��t��.�(r-� ��  ���=5ۅ+9�DR�ZE'�l�j����}7K:�LEFje�A�w4Ij��ֈN�w�Q�B���I�\�e���4�_�d����uG��U�rI�p�wz]f6��3��.���e!���)owAL�9�AV94��n����q�Y��5��7C-Qbˍ��Kr���B�]�zfuu���&��'&�U�.ӗ�-_�,��m�*́�vt���=Âclָ�Y%򱇳W�ѺN��"r���CxX����b���W��-d��h��YV��m�gz��ą����<�p��԰1L�v���;�-���fԎ�7sR��K'F��./�Ϧ�5A��������%�7C����X\���{��=s�L 2����z)���?��7�[X�n����Xs7yaF�Mi���$M�r����ʇE��~&�.�B����Lc�t:X×z�؝�f]E;Gi�5
sR��%kx��.�u�>�J�Jΰ��V�=��މXF����ȝ�pӼ�w\Z������u��^�BԼ�j����e��&����J�N�-N�������a��D=���ލ�r�q����F/�KB"������6e5��"��pM�uk0���D�z�Wc�8Z���U-c?mi�i ,���c�75��#��V�h�RqW�qq���[���	�1(3qƍ,C��v�X�i�[����Ysu}Wo�7�Sf"�1%˞�V�b��L��r#��|��*�8�3	�)4��<ǁUC
]o��
7�_�6���gQ��8&r;����L�bV�*��Ɯ��6F*�_:��ͣ���#����<�٪U��e73�'�-g]3�CB����'��`�6��Hۙ�n��T��WI��Zb�
Z�&\`��[KM��V�و,WLC���ݚ)t��G���`}����~rb�u7�� �F^��qm�i:�b-�zk���uL��ڙ&��
��|�q�[�������ox�HY�XGF	*a�&��ܲ9 �)e�̜��0N���범���	i��P�i��h+�!w	yt��͜��7B��wZ�wQ�ڝ�$$uf��v�е�[co�ʬ���34HV�ַ��1��<K$]�޳�p�`��H�A���0H�c��1��1[su�k�����kι�e2f�7}e��(���1�T0�7;q�����u"��:�}����q�i__TTuj��ʄ]:#pj���2ŗ���ai��vf�����hv�Y��{�Q��2q�H�R��l�� .�n09!W�q��K�8�o	��4.#�Fڍ7�06��Ž����Rс��z��]�bu�^�x�f�膼8�9�s�:��Y��p�#�������*P睎n�[,:$rǓӫG`���8����� K˕zc�@s��k;o��b�oW-�'�Pݡ؈Ϭi�vR�4*.��s��w.�d�Y�S�L�*��]n*O�uN|:�Y�S�-5�hL��6��Z�=�Y��G|���ٺ�3&��pmgv $�kb2����
a0�RzB�OK����ӟ0Me��K���=[������F�8q|����8Όxm	325��q�'�}����j��(8���+�J)=� �]���S�a�%1W.����{z��f	�v�;Zn[G��$4������'=��Wm�SM�T�ݗ@���0+e@�-��66�S�];RXk�<�W V��R��ϗ��dǬ7Z
6tUxt�7�	B�Wq:�/M�_7Z���6�����S����6�ͮC��>5=ݮ�{�y����Ǭ���#H�F�/Q#5#%
��q�b�KH��X˻�b!r\�]�.�mAU���IP�#X�fJm�V
H@.��,��cv�B�(�]�I!lmdI.�K�F1Yp�kI�n_n�?�_�8�u���$q�܍b{�|�M��dq$#Zbw�}������:�#Z��U���;gO<z��x���Z�}����vu-��־H���죉���!��f�
����O���([_�Ŋ႗o۾���:Ʊ�hc��S����Ҽ����M�O��x��/&�þ�z���N5�Y���o��6r���&�֏�W�����	�<iVe]6A�MN��e���SYJt��ʍ_O��M_&6d�F�gɷ�w�f:N'�%jJ�7MzZF٨[mwp��Z��s9��oz�^�rZ)���ަ�/u�f��q8�pZ��-+^����Qܖ���{��6�z�����ׂ}~k\���:�C���{>k���J��_]vu�9���u5�W�^u���Yӝ�X>��H��HQ&��e��L�֟���}����]&�Ba� n���v�EB�,&�����u�Wyt������{ׄ�0N�=h�E��{7��<c:O��>L�*��'{���vch��="�11_5��o��k�c��y�k,�{q"�Wu����k�Cw1vx���������V�"cE���h�3��y6�;��N'�_8��޿���4��m���i���N�9��!��:ni�Ϛ��Aq7�Y�[��|Ő^u?"��T��[u�rR@N�|_����^ﻧ0�:�Dv��}���}t�����u�_p��hB�8)q�c� �w���m�4��k^�s���QۏS�BV�p��i����Ľ��6����#��G���0kI���淋+��m�Z��O'6Cɿw��w�����+ihyϡ[>�\��;f+B��CL� �6�'�~��wtm8��!��(
r��4�^�Զa3�}Q��RR̎���,��p�J��:�����n�k�O^���'R?p��b:?!�׭f���!���yf���\�tq�;C�Z_ү��̚^�+p�@V���>B�
W�2�U�ߧ�9�#Zz�t�mY��a��j|��]x�+HG[f�}7�g��v��~~|�����5u��M����۳7M�w]�X�����0��;v�k1���9�>7�m�hu&g�hU!X�-�
�C9�� ���{*�����]PoP����ܯ>b���i�q����j����ɷ���Q��kI�_8��n���i��~��M���rW���gv-[Ǩ�1Ƶ�~�Sn�>����bu����]c��\�o���:�t�p���2��^����YS��i�E1*!m�
�P8lU�(
ѣS9���~�e�v`�P��|1=e����+�n���u�x<��Sv�n\К�;e����|)���Ǉ�*m��Z(����%cDN}+��~H�����2��J����ݝ�����f�~h�TC�mm"w�^{�sru�_&���Km����g_����M&<C�&�%����Ӯ�7Lc�IưO&nQ���5��s��R�;�Y2Գpڹ��ǝ��moP�6�Z�T�Y��ߜ�fl��v��=i]�WB�O+7�y��S�%��^�E�����G�9��v�F�W�.��vcV�)�2Mk�֓�by����������|���Ǐ����6�C_M�}�[E���������;�>�������q�֭	%�;�;�~�l�C�Dj�դB�>K�}�{[���<M�CIQĽ��'a�ʎ<~� ��i-���������Hu�{|��7d*ߍ�فĴ���0k2smT����4m���m<�\�b����qR9�.���yi
�=��{����M�r]���-��m��5��r�}g3Lv��i��O�u��,�W�&�ќˣ���H�<�)����56�4rq-���q.t{p��N\6��О�qN���w��ԫk�M:k���3O��c��?'�k�s�^L~u���6����S�cV��ﵛ7߬��h�n����ܝ��R�'�8b�м�)Z90�%p�ؑ�$J�%p>l(t�Tl�mu��o�f��+�>���w�!
�4��R7�<*��߽���ָ��S��nC�o�������u��q���7���%i�������{�&�4g�i��|���K�:�\M�q�ZkrQ������7�h�*
�(Y�<l/��VM7��!Bh�>���(a�Ưy�S�z>)ϧP��ʾK~L���W$������?��o��^���?�]F�c���� ���W�jNѻ�$��r[F	�&���1�����&� m�U�v���o�Ƚ�*��C��ê�]՝j�Z�[Y��auhİlܝ�G�i���B�Rf��+�P��C���>.��cZ�L�hE[W���5E�I� �%]ks���)��O5�h�N���ͅ�D��^��.��W�g����%]��S7�u�a��1��Z��S������`��kW5��A�:�w%��v�8"u� ��j6ն��y�T��,ƫ�:9-�('��畱J�L�zW��B�t�d��ܥRbݻ�0�qvN[���m���@�?�f�n��^�
f�M�[#+����� \����$��]ݒ�$�I$ ��RK�K�nմ"n�D��WXZ��*.�Y%)%�b��TnH�6BF\%��UwĴ��$��U�d�Zr*ܻD"+%([V�-D�#m�#mF��F�TPI&�Q��1Ԕ�n�����S�@Sk"�G�&�x~��ۮM:k��4�Qĭ�z�����CLb)��Bӎ��Ǝ?��ĽN�k���Z�׍i��#ﵔ-�oN']�M����v�vZq8�$��'�?;�:���`-i�h���o鶕��ט�SH[V��Zc=�r�4q��F�"�h[��W��Sy���%y8�L��K~_G�<x�]�tM&>N"�F��^�x ;������DL����e���W���'�;���C�J.n��;��]]�\t�kXC��C����|�5��%|d+�v�R���1C~��b]�{1�5y���6�R=q���y����g�X��P�U�A@Sk�w+�\N��y7�m���z��ogIG���6�1-C>��1*Љ�É�5�~�y�8���i��~�����q�4��X���B�,�{,Ƶ{Ӳ�8F!.���_Ñy��[-^����Իq�NW�oM��wJ��u��j�Y����,?j<0p��
��oe<].��ާ���g'�f�e�n�.o��4b|�x��&��ebu�����q:�~��c[�^�����h����Q�mm"u�__}��w����^�B���3�]y�fw=�6�7���C5��7z#Gͽ�&��,�7yu�w�~�n�#�M���9~M}6�I�����g�wםڳ)ԯ���[�/c��A91�a��E_A���R&�z.��_zkl
����b[@f$��ɜ���Ry3_#k��C� ^��]vo)���y׼��y��x�~K�A�}�ue����۵eY�!:�;�X�z}i���@vt�.e����漽��BĐ�K�Vϑb-�{$n�F�|���u��ZD1�(on��R5�6��{�=L7Ѿh���m�� �y������KH%J����q)w7XGӦWN�6iX�y�>�ع�6*�����^����cxz8Ko)Ƌ����W��F<��+�λ�|TČ#n�M�ϕ��Fأ�6��;*�N�6�#��f���>+�-	�*�ٝ��u�^#��
U�[��zo	��=��e�<�����y,X@��tH���r��&�����}�6}��� ������;��+�9�ݵ����Žn�`:�]`��0�&g��\(��˄ޅӆ�WF�3�u����.��j���g ���=��1v vm�v�kM���С䫚UQӆaWU��9ݬp\���Jp,��T�~Cȴj7��jj8�&Zʯ���_�e�`Dߴ�ꪅ�c�>¬R�;�	^�[^F�E\6���6��G�:�����4����������,;5A��u����5GP8��}v�w�6�0��/V,`���Y3��Go��=��K�E�*���co9�u%�$�΍������������}܇*7�h���~�s�]���Y.p�eޚ�R7-֡��M��v �m�HOvSA�-�5fm��Ź�����e=�'Z\�W#�j��i69��u�&z�f�Ս{c��%�u���.�Ħ6��%G�($d�T������g��T8*��e�n���1�Z��\t�O���s�0�K7����{�q�!�1�5m��0�2q��J�{{���3����s����Z(�U�ƃ�Q���6еTcU[@�%F}���ƨ���h�nQU�j��P�F!V�GZ�45Tw�8��h*���EV��X�[U*�Ѵ:�Q�J��ٍ��O��/?[}�%�)l���=]C��=�C
^H�MR�6y��_@;�4J��77�p.yY��Z��
	��������W`{+n��:Ґ�,���k�W]]-���ߧ�n�n�{��֍�r<*�-�jA��f����ti�p��O�0s��k�FY=by't���w&.��P�R?������!b��kI�}�;i����_���P
f��Iֳ�����[ц5u��T����(�\��*�q���#��+KT\�wc��˱m��\5:�fp:r�l��e	�n oi+�#]�ю�x�WWn$�W֤8��,I��d���'���p�JZ���`v��O�w�_��W�AD��"D�p�	r47�����D��JG�L#Q2�#*���-�ĉ	K�h�-�M�2�j%Jm�:��Db�EU�R팂]ݑVB1!�bD�#7pj%F�M]��R,��u.���D��6ő� �y(P?�~��(�{�D�x�JO�������T|�Q�rP�E���)TD��1��F� ��rMWݼ�U�Ī/��檋��� cE�E�~Z�J��(�_{�Uhhƪ���>J��ʠ�!mm��ڭ�T-W5���m5T-u
<�Q{˪��
��W�!�����U4U|�ւ���TTj��5Zj���TOJ6��V����٪�h��A�h���ƨ�%QԪ>h�%s�}����;Tm
�Q��A[B��J(��AmPK���¼�|��J�GZ��}�(-
:�Eij�-�������ڪ9�j���[T_�AƎ5E��T]�~�Qƨ��Q*�i�T���B��ԯ�*�	X�����p`+ȷz4��טE�4F���#���������\������
+mP~R���(�A���R5T~P�Pf�Ɗ.B�ۯ��o �Z�1mcEWZ�j�S��A�UD����}�t�:�m����U[U����Zh0J��U�L�e����]�"k�]�O�/K�+B�)�^�ׯR��4Ԯ���C�F ��2���7�6��z7�7`�^�p'�A,j*[�W�;�^Smx�����sK�����s�1H�L�}�}T���)�Y�v�L�TNw�c4L�c:���w����W;�4��,}3{`�m��z���^@����x;�j�q0Oi�f��W�R�ݷ{ݺQ�`q��R�c��+9�m8'fz���G�;:K�u��>�s��CeHӊ�#jO��}�v��߾�7���9c`�����D��v��!=�v�K
��Z�b��D�5`Lz�{8��W\i�2NPiP@Uͼ��m���}�>�D�y�n,u����x�Jy����n���Z� ��/,ν���y���%q7/#	N���������?�+��{���&^q���V�2��z�nx�|��=V��w�Dج�L�'²:���y��v&OZ6О���q�)�"͆�뫻����ݛKp��A SHw�WfCu<�uG}�:&bv��ep�ƶ�K%���GjR;I����L������~����rDzͼ�H��StY�Ev¢Kcy��Jewn��3����*��Uᰄ���BXZ�ϫx�ݴ-�V��r/dc�'�4���
��:@��2%^(�u�7���qW�n�k�l�JH&v4\3{wqj�"<� _f�_��Q�n���#�C��-�N>��tn��ܷ-�δ�*kˉ(y��kU�K�����	���'�3sݏ�wc�4R���w��+ӷ/�@�Q�,�����7��H�9��U�~Wu��u1�5Z�q�͞*~���@�YƉH��p�����&^���/E���N��T/"�*JFi�Զ|��>ߤ�o 3u>��s���E� �%����=l�ʯ$6�ޕ�/f� ��M��iަ��7n�I����w�� �U�Q�e�.H������D�=��P*�[�ٮ�K��lיoCI��;r�=o�k<���$�c�ˁ�cþ�pC�\�}�+�ʗ�� ��x]3.�V���fTE��6Sh�)E�SJt*ԗ�j�NuX����(��7�]$�yerȷ�g(�x�Na�])"��۟����%�	��?����R���;[WCG*�
�-p�8 ,��u罓�t��P9ׂ�q�P��t�bai��^�qb�@�mnZ�Nx��l��x6��� Eb�k U���B��m~��N��,dV�T�%*���7�<ӱw.��B��3�c����_�J�^��7��a)�X�v��CKJ��MtÆ�й6�mk�7K���J��brn���障ފʉ�t7Օ�.�s����X8�"󸭸0�t-#m&f�t�E�˂H��5ػb�uj���b�E���N���b[���z�s��a����F�Y��n�����s&��}b�!�	���'y����my"�B�Ğ�l�F�:.���]t��\������S��`Llw�2���]���<u�:�����AgZ���R��:���
�(�����L��w�Q�������Zj�"��ѥ�VH�0nK�Z��f��a@��1n�#5�Z�H�3W. �Z�5��ĉRH˄��-�.\�l�d�B�$q�EY"��#�B�RZ*i�Ŕ��ܫ��v,T��1#��l��wc.�	0��|A�����WN�5,���zҋ�_UUPI'A{��r����+��a=�ڇ���V���Ľ����z�&����t�}��ѽh�i[�^�߻ �Iszl�LK�m�c�ȸ���r�9�Y��R�'�*h���S[5��jE��	Ɍ�������|�]~.s1�Y�A=��S���/ݑ��N={�{4��Ү��S��i^9rŢ��:k���an2,�Q:_<ɾ̯_��oq!EM��N�ީ�t�H�ﶁpNf��U�w	qH�w�(d��ҙ�����^�޾睜�82n0�1�2ޣW~Xy�?_z�d3l���kxȴ^��9+s}<�d��1��&m��:}������u|�.9�8.�6r�n[���Gk�쩩�<��W^�?��V�Y�+�����Ĝ�����ȏ#p��S��c4�ֲ6r���c}�w�׹��򣦗����>9�P[,�8>�Z���>��U�tF����]ڍ2"C�8��*�P�n�-�Z�Y�U��;|��YSF��b��`�|rBW�]tVn�9ԓ�"�
6fi�[�is����#�$�|��^�;� W���^�#f_UL�}յ�"�B]�U�5�z�1�s����;�,V�Su���%4Yӣ�M�'��E!�+u�}̍��2���U�ax�EF/i���5�����ɤ��U���E�뛘]�<�q�"E��ꯨ����~����������.XWtH��{�F*,�x��X����p������,�+��;o��Wbi/E��9k���>&fW�^Up����T|:�^=d�h���ׄl˝n�Q�DS�'?U}�Ug?޿ߎ��S��/��ڇ��T�G�Oݴ��v�ߕߺ�7�4E��Y�w�K\D�=˕ѻ��q�	�X�Ҿ��d]f��C[jIA>��Ie��~s�;Fn���(m]AK��z�
Ԋ)
��Č�ʏ��W��Y	~��3�&�p�g���e�G�i�6��@��v�%���ޅI�w>JgC��h%�1��U����VA�� ��T--��uiu{q�Ո��z] ��e�PN�}��z�R�3&��)�yl�|�q�%?}��|�7�_��p�3Z}�c��f���&?��;�g˯|O+�t�uU�n���M�hUuy}�+�&��^�{x�A@��n�AJ�6��ϮaC"}�c���*��w�^N]d@;�|�H�+��{�)!y��E"�Kf?�TDu� ߤ��]�%�0mۜsk�^	�`�]��k��~�nsײ[\1e��9�,MwLT��f��X�vh�b��l�et��Z3ָ^��׽�^��`��A�ex�N�ԩ3��L֗8�u�.���T����d��JT-Y��o�hӭk� ���b�=��X���;j`'qXxh�4F'�{gi�b��gMb&P�	��	N�RR�cs�4�6�{oV��t�|�`G�JJPG��:��Q�+"O����ެN���qOQ�r�M�y�v~e��0e���"�q��iQ�UŨdC<?n�o\���U��E���E_df-��!��m����&�֊���gU�|԰�/zZ,6�[3'I������$1Q�t�3�{��37�vr�d�o
h������JfV�f�u�w\(ub.U�R� ���Pt�p�.u���ؚN�N�i�*)UH)$��-����VѤ�Im��#):�QDu I�5r�Vڌn�,H�H��(F����*�P�Zf�0Uicw��c-�yv,j*ZE���Dd�jEKb�H2�SN4Au9�R�HFIU#J�o�o�o��u�x��8�����U�u�����W��XG��&x�ju��Ө��o�X���[ZEp�u��z���n3d�\�� ��~���L��;f%QW"N$Ff�sʏ 6J��C�u�����]�hqS��B����X%��])��6ӗ����4.�]���k1�-������~��SI��u j"{�΋�:z����CU�m�d��x�`P�E�W���S{.�r��M�v���Q��L-i���'bI�cV�[�5��H�L��U}O]~��|@���v^�&�xo�����=�e�:ګ��\�abx����>9Цo�f����ap���uT�<�����=��(��a�^���m]�9G��ި�����X��\��ޫF>P�N���QO;(����,��R����FZ��S�?l�N�b��9m�@Os!�ܢ�&�[��~��^�6��;inͯLg�5����X;�	N���t�Vk���Y��gQKv3�^i�,��r��Æ?+�~z�	���BV#�I8!җGꯨb����c��>�,�� �L��l鰾i�u��k�_��C������s���>�N�Q��Xl�.�>���x�ҷ.�ؤ���\�$x�ri�\���@���^���U��w-T���I���5�`��CMȃ�1����>�@��#���}��>س�s	Uһ�R6=���`���%�ݝD���*�w��qf6pC���lܼ7�h#p�x�����䘣r���9��4�#���9��}���"��G�bo 4�Gd-�
�C8''��!��UҼ��	�ʺ@�?�+ɉs�c��&�%�ڙ�4OcR�Ξoa�6��o�x<�q�}�xT�6V�x���k�1Q6a��&�,Ku���ʼ5kuȉUW��U�_��>;��B���ы��j;���j+�9�@.�tΜ���\+=*lWF�>���l{�Z��Kng��\)
�E�cy"�B����z{��As�� ��DUK�q9%#|z����Q�cӠ;��r�F+�%A��y>n�=���ޔ���ܑ_����_]��xǗ�r2� Z��3��a�Nhzv���.��t�����(��*�5�0�̲��s��CW���ƕ��3г�5�oǞS�9��{���k���+j���t��K�O�lk�A��V��k\yɌv�j�˾����r0w[93>�h�����];�E۸���څ95u�59�������U��1�+�ܳQ㡾���u�Pj�j]������R����Q��V���5�
�o랺�q2]�?8ş�J�WD�#8I��U��^�oQ��ϳB��|���LƤ�MM���w1��)�؈����KF�����6��ʺ]������,�������
��;Ƥ�2.a�tq�9c���W�O �e-CiQ�����3����kXԃ�
�e��h�������K��Z`"��a����vd���d#�S���S��mG��w����M�����1b��g�dL�_���m��`��m�ŋ2..�NRm�q�����Y�%��5Uζ�Q�>��o���qJBc�H��t�0��wc�R+ݬ��.�	�"��AJ񫼂�j�R���[���7���s����.DpwqQX��--��nZ��U�����H�(���p�@�))GHi�d��W�%*�B4-#X��Z�QV���d�4��"Y4�X�ww��UuWu���~���
�H�����s��������_&?G	~��>=��Dئ���E�k4-��>r�k�XC�pg��Ac��*ў�K
�*�s��ո��q�}%/U�!���-��W�g���8-"���gՒ(iB��&�E$l�[�����9�������.#�|.׽�>��"/-�v�`�t�X}�L��[�=��`Ϭ�y�w�>]��N�aa������?lժ�\�u�dWv���Û��R��{:�G+��hpv�ܳ�:�A�pN~���S��պ����?5��N~�21ݬZ�op�GĎU��m*����]-M�.hU�" ��u�Ũ�ءM��)fs�u[֋�l�Q]Qg��M^u��MܱsY�y�+�U�hS�BIv�0�[��#�f5��PE��~�ʰ�����k�wЏ�tiKۺ,Ӵ�J�Z�
3}=�o<��:�7pC�$��W�k䴮ٕ����}�d�o���^�`hg6�nmYNL���{K�Ph�iYٚ;�i�L�\���W����g�uo�\x3vow���x��T���&`L��Oo��yGq,�6�3K�(:�y�t�Ne4�;��cp�->Gwḙ�s^$���eV]ٯU�x��{�7f��\:��0(�ݷr�U������Y��j�)p�ﬄo��]]3ZF����eB������6�1�#T#緉iηk�th�0�/+�3mh��`�w���5��c2�)��JY�oR:�m���>k�wU}{x��z��#��9������'jZ��-����a)�������{����(I��4��U�ķ�S��O���x�eԖ�;�T�[T�iBx�Y�o��ub�}�u4�J�*�Ս,����|X�n?+�Ӷ"�q��C�o��8ۖT�d�wwcKWB����ڽ�<����{u;5�_�n��f���;���}���O������w}����ymy�k�zS���;���e5�G��Z���xߗ`�k5�E�ݫ©:����z�����%�Tg\%ڽ⻗_j�_""#�����z��WN�Y��HyR�C@w�z&eL&����t�=��.���u3$��u��Cr�ۧ��@Є�׫W�ݑM�^]�f�zu�����X!��}�7��`�S=y����s�()$�@ې��ӟ������곡�~�Goq���+��1e�D꺏���#�*�{�/Q똜�k	eb��0�Ee�/�tc�����|}F�7V�Y�u��7eFv�-3�Df[����Z��Z��b�{#$\w�H+��b<���}9�m�x���ï���XrH�RR�U� v���ջX�5.��eH!{�6�%�Oou�ޥ��<]򚌼]�,A�Vt�b"u��{Xw��
f��*&���k�۸�V=un�j�@ˍ쳪�o)�Z�mqV������4��Y��n)	j,��Ԝ�f�}-��҃�� {��]�Z���\aeն�m�K{u�\����X�9�sx�D�����ܓ^���R�-J!s��&�u���C.�a�lq��ҫ�T]�Y�p�֫x�$�s2�
�3�[�i��CR�辊఩Ժ�����NBB\Yl�UiF�5p�����U2-�e�չu֮��RIJ#KhEj�Hڑ�Z���4��m�-��5"�U��X�c���0WC�F1j,�*�v����������*�r��(M���%G�($a�T����X�n�2�[�(߼�7-�=W���6z����Lͽ����7N�8i@����ə��ğ�9�-{g��ɨ�P�wU�LL�kuѴ��������<omLr�k�_�/KV]f�{u�D�P�r�j)�QS�W�W�'��������qfcK�WE�Y�z�Vg��̷�ஞν��PAis�5��1r�����t��;/,heF��Y��;�F֌|�^s���GkÎxjٮN_7��a�$N�����E�1�tvM��9�:����8�}��}T��|G�%���޽�c��U[�,��O{\ͻZ}h���f�r�z����I�gڑls=�_]"��ڄL����&�Q�K�	��|Yv�]��7�	`|��$�x�thH�������"q��g{�y�/�5(������������v��Ƕ�{��7W�69�,�b%�Z�XT�l�D�����B�mX8��cɕ�	GVb�Zդznd�v�*��QŻ�p���w*1m�4f>��3iH[�ԅ@ӟ�������Z7 Γ�og�Ͻ�UR����}9���='x��3\���n�� fԸ';��Z�.nsXU�al����0�N>'�u79<\��� ����2�^��^����kjV�BRT�n\�md��Ÿ�}�_?]�h�V~�ܬ�e�}^Aj\*�H��ǫ�$�v/�sY�+C�^&�MF{f_Z�K�D��ak��.�T"��-������@]šw��^m[�&�5��a}��I@�93p��GeT����麆W�����:?�2�t=[nY�;��-?8���K[,�}y�O3�K����Di�Zb[%�9P��������,zcEt�s���-G��"��y��������f��<ۘ}.CR���z��ki�]��5�殰���4�+����_,]���o�Hx5�8W�.�̂�?)���k����ǡ�v��Ruo�{�����&S�x��f����K��,�Y��VerC~�yߺ��>�|Y	�$1V��ns���J\���v��u���TYA0q5�w^*�!N]���t���,�^X���>�Q3��\,����ФlV�m���#�:�\R�����zΊ�fG}�Ը���3|��y�tш;L� )�5I#�s4r<��}Z)�vV��?�<$�\�ƿ+����Bu	W��An��}�"/ۉ�w��6={�+��N��}����Oz�&2����3k����o7X�����K��`�ŪwfQ�u|}�(\s-�K�����+7�E�"�h���]k;V�m_`��v��(���+�gLܠ��35�w���E�A����[ܩm0����ڴ�uC�ւ�^!��V��^�R�ßIO�7�J��=R�[�A�s��ܮG4ѧ�\S15�|t���[y�r�Q��`Ֆ����iQ3m���V�q�n��0[��v��e%b
�WQ���8��`�%�ݏ��-⛕��ф�+r�P�Δ��2īήhF��^�a���LE�Հ������j��SKq�J͖����o��\���kV�Z��fBظe�-#�7c�!/XZ��"v�VA"Jd��Ս��m�RIPZ��m�դEnJT[��b��R+rTH҃��+iL��L���M-ȶ������`����l��55���2Ei$��"��E�H�$Dn^��$����ƁIR�@f�Lr���k�k;��|��ÎW?���zJ�A��5_,{M�v�XCꭍ�}y,���.�7�Il$��2�VL�l��hP�IzC�����>F��5�Q���>�r�b������b�{�[��ِ��/i��M]�k��y5�/�1&�ou8�w�(���=�}�zlj���ZDG;�ܩgQ�˭H��!V��Ϊ���/��-�!��>�.q�J����V�E�T�x��:6���zCƵc{�f4�ֱ�˦�q��j�J���()����"���/'�v ���Ŝ��8�맴;��c�:��Fk%��z{��o����]0> y�Vvc&��>��2����14Ft���{�P��Z<2�N!��+k8Ӽz�t�ʺs�K��HoN*��ߎm��:�]@X��R��"XiE"��!��It�t��P���H���ިK��z��Zr�Mhz�/�!�]{�T�q/8� �P�կ��yȨ	����t<=�ii�L��YG�0�k=�����\�~N�{��3��f��V�Aq��k�I&pna��-�p�k�Q��~��#/��=�:�s�sE��!�>˘&�ӭ�C�gK*U>s�̸��sƁ�\oX��X������a�-t�닋t�ŝ^�Ibش�r���'!t_:�Ѱ]������ۛS�;���g��Hjm���۔��,��.MQ�ޑ��O==�W��+�ZK6��ȇ��s�S�����a�nx�^�vG�6ըNч���v�XY�\6\�[�=,.�^�i��)�U+�U�k�����!.y5�0�]���ڤ�C��G3�;z;W.�Z�yP�U!��{�o�虳�5�����$M�g��,�nK�:��9����gx�e	ۖ{[�4�=]�n�f�)4L���g���.x�펢��֡�~/����~\X_v�[6�q�n���B�繭�%�$��Q�9����g��w	�ڏ$�ޫ�V=_��u�#���)����wL/�J��=H�~�ԙ��v���ےbd�|��Y�s�V�1H|��ul�6���!�&�l
��Ξ�6�1EX؍#��:���kUy��Eq��
ai���Č�ʎ��b�0����ݙL{R�P۫�@�W�(����q2�d�;�B';�o�C�� �'3�-W�N�mc�<��Ϟ���yV�[V�ø���_,y�z���$����G��*�S����e����;l��[ʟ�3��F�7s8M;Z�o�Ac5��g�\��P<�<���ǃ�FT�(�,w�X�x���wt��޻�vdtF("��@�Gո�ݵ��U�r���i���R�f���3�G�NU����~�c#�KM�:�_*�x�
�7�t���g��]<N����u]^�XKWÐyO�І]]���{i�J��0g]қ��*Z<��e���v��3J�˔�k����ɜӔm�w��޲��Æp��c	���^S�ˬJ���A
��� UfV>�G��(X`�\p�v0��0V>6�S�{ً6�rc3��Y��9����eBP���&o�,RM�����b�+�g�8$�}l171s`	��6���.�"��J+��e���k�A�U�$Ε���;������ݽd���

`c ��/v
�^SG���٦�Ț��&�YQ�Ғ�س�Rђ�qB1�i�Aj솵zf��%
-TKJ[IpF����5�4�[e�D#�4֐�`7�[YAH�\���֥U����F�`ЌIwur�Im�d�O�z睻SGE�l-K���ˈ�S��7�Up�Ƈ�E�vI����V�:�>��7]2�����
��ܮ��ը�ć��>�'�.n,�e�fd�{.1a�Gd�[��,#����ҽv�ťU�"�s�L1�h�n�b��\��B���]�Y�b�؎)9s����v\`<�o
_tS	�5�������Y��ލ�ì�h��Y��:���y1x�_	����ʽ�m�G��3Җ�Ǯ��p��R��/ףг��H)��!�:u���Y��Li�b�C�ԔK��)�6[�Qѝ��w�s�)H�\)B�l~Y����]=i�)�&X�e�5��%���h��M��40>Ɍ��7��Bb��Yu|�,uZ⮩^�}�Wb0tni=���/�����W;��ƣV�r�T��w���׸ݩ._��+G˜)\pm��+%��C�^�C�]��f�.&�ǽu}����-�wVy�V�^dV޼�u�Xy�`vqEmU����`l�MK��Os���ͻ�S����rO%�܂yF����L�Cpt�Gi$�+�ƚ>�Cngv����r�Z�<��s����5v������ɉ����9�d��s�R#焨(��|��0*3]_g�8�A��3.��bЩsm��H�*ד.lݛ<D����Q{���u6sO$2\3ZH�7>�����|��z���2�{��YW��q�w�ɷ%��$ Z{�5���+o�4^|V{����pՅ��E��@sˬ�o��K���^SYcY�wYP3e=��zy�,�Ե�uZ�~օk��az܈����l�����}G�s/M��#{�d��,-V�v\��Y|Z�f�;��fC�`hE�ͨ�Sos�)P�Z0&9��][ �e=Z0�cD����&�Wsz�Y-؀}�v������$��ወޏ��k+3�)��GM�gBِ�$:"�h�<e��=ǀ�����չ�-Ӗ'���R��-w�6�f�w��vcp�@f��+P�J������_m�,%� �$U���1�k��B� ��u�-��M-N79Q}�lv�et��l�n�kr�#�5�I�7�+��z�2�&~+}Dpa����GG�Wh�Y��1c0���ܻwk�)�7�2�ڽ�<�i����b��'��Y=}z��C!��o�'���k;Nu�=��x�u�q�\�U��q��kˡ9��"�N����X��5��w�#4�W�1��j
\fu��#����F�������Ǻ,�dc�g4�^E���f�1N�}���n��cl�L����}ˆ�����J_+�%����C<E�>��hyeɧ���Q��A*�9gFk�$l�En�ሓ�;����Y\�bw��Oi't1$e���@��3s/�9�Q�@X��YMX�Q��&������ ���*w5�P-!I�x-��S�Ӱ��N�w8�I ��삻�.Wv�e���u��+��`gxEl� �&�\�9�OvK�.`�����)KỺ@��L�gM�n�������V�n�E�DB�q��%�^4n����qn[����U���b� ���� ��2]n;��e�c�G1�n捱5�m&,�l˴�a%�����b�x�(�ڡ2c̼�C �2^c��:���ke�96�gX5��mY6;i�]�힧b�ժJ�,m-���ݶX�%�X�"'��!�¤j��tX�%���QU����j�K�U�.JD��ۄ�\���\��MhТ�[w]ڌJ�0bE���{`5�x7��\���4d�D��w����Z�M�:%�����Jb�۬�6`n�lo�����gι�W;s�!���d�(JX^ܔX�5�o9c*��������V���ȡDE���]ϡ3Н����w0����;y�~�ơ���1��aC��X�{�;�&E�������x��Q���ဒ����>�΀�K�T��v�j��� ���,��WZ�=�S��C�ZdQ����1�3��`�Gk���,
�1�tz�7I��M�E�R�����N2@aܞ�2��Ò�[��b�4���9ͮ�Qצ�����<n�M��h���mM�9Lc	o�]���[�]�<��إ��VT9َ�N��?w<z�Wn�|��mݎ�IxU�XJv�wK�	�+wn젋'�^#�4I-�4��ܭɽ瀽���K�����s{,|����1�J��{���M�� ����3��td�k��1��U��g�T�`OEY2OH��䕖�su��3X�SY����tK����K�t#�Z�m����d��&kW8�{�ȸ:��7(���p*�m�f8�� �<CzU��EZ��a��t�)�ō?�/F?+OR½�����6Y�)�3=��ߏT�!��x�绍�uy�фT�/<e�˷uoҙ)�CQ(�
��{�h4��xW��u�r�'&0nf�Y������p��JR�b)Iܮ�g�Y��Ʀ�B�����|'��Z3'oz&�i�ӡ��仳ʇ���Y�sJ�2+u��w�R)�y�_�uy]q��s��Y���Uy����R�u��\0+���J)��BČʎ�6k��B'�d�5w֯p�m��h8r»_jC�h�׸Vn��ʡ^�0#�kJ�+7���MM;���ќ�#-�I�سZ8����_��������TFa��5�P^{�3�.	j���w���R�(Zx���cXJ#�RXӎ"�]�5�����n����a��1m&�y��07����O�'���k����մNC>�{�����U�K��~?8X��=J�xm���<t �����I!�ͮ�5�WS�nJ#iԷ�o|�÷v!�&�>��ry�q��Z���U������׾�מ}"��6�T1��v�Gn��{{�sO��@
p�@�cRG{�*i�l�ێ��B����9�p��,��p��\KK|�>���5�|�GGeʯX��h�*
���khC3}�q8��{����h��v���u�n�祻C��LKC�4l�#5�C�'q���&'snf�B�i�CG��Hև��̯���~����K���m�>y�����B&�#mF�k>��;�׾nW�~9(�,ԡm6����{�K��6���I�R�A�N�w[y1�N3gv�-Ν�Z8��
Y�@U�@|b"[�Γ���[�A�<5��4ן��ߍ}��+OȾM�m<��KLugt�4`�CHUp�WƇ�,X�[�nXh]��ߚ�18�kw[��������G��cZH��>�~M�C��U��]q{��x���Gɷn%�o�	ֶ��(Cg�.5vjuF�HGm���i������?�~��߳��O��TQ[�J (*���~�(*����R�PW�����NX@�%G�ʅ��ݢ�a}���!���h��P U@��%P�p�����+@�He|��h�@AziH�b��Dw�\kᇡpMA;��2�bV��D͈@R��s�};ƹ�~zo߅�	N���+��\�@_�sy���s�	 �M������@A~	��BIfr�|b�:rH9�B�г �f����ϩ��l�9�$m� -� uK�a�� aQ��D0������h�-V.^�VN ?�L%.iذi�=:��[��0�V%��@|	V/��ӖzSl���@�P6�'@�'��h�]�g�q����p?�¿?ֆ8� ���$�o.�A<^�f�uA�3q�ӂ��ϝ�o+���H����!X1�!�� ��7I�KԘ��_�� �"���Fzě�@H,�.��c�x-�z�pn.q^�wy{�I� ]	�0wNш�)���]2;�� E�FA�@_W��q_4�Iu�
^u�Ɓ��I�*'afy�"����i��?W�:W��*���i��U��O��� �O)3#R+����ke�:���vZP�.�xL?2� ��&�8� �M� �Ӵ�S�ixhd���=8j�ay�=y�Z�G��S�$��a���ه+��N�N�JOٯ��|K�p)�B�GP�:s��z�wZL����~����s���jցdE��t��P�	��\�� qv�p��� �s��q�-�cu᤮4��l@i��\�V�i�,��	t���E�N��iW*�^��AdIP�<	
����}�L� �gn��M��ں̇A	���a��\+a�;	U�+9r��k
���<Ri �)~���rE8P�<�