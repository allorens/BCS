BZh91AY&SY^jd���߀@q���#� ����b@��         `@
�
�  (
�  ���   d �*��U)@(	 
��H(P�
4� ��֦���͕l�ق(PP٪�A��[46�6
-�
eE �hH�Z�m��iJ5��M-�h�SUTU��>�=��hV�g �Jt�[YTp�N�m�m��-
)�m��Cb�� 
��%T�QM ��CE* ����� 4S��T  zR� ����%k(JK)�>�A�4�A�5e%R԰U:0�� ֥m	�:�$�Q��c[Ut5L����4[M0 ��ϥP =��)�h�{ٯ{U�gv�+vP��`�̯p;��z�Yv�m���8���R\�QpSA@A�Һ����xݽSw��н�{ǥ��Fت���P�(]��  9��4��t��=�	m�����(݈u�=
�#N�*��A��:R��y��i n��{*��o;ЯKn�k�t ��M( ��4ʃ6��Vo�E( �{����F�w{����������oxJ ��.���Ɔ�s�ݽ^�i�W7O[�*W�t0{ �J���� 6�g�tvQ�ܪ��(���M�K|}R� x�}]kJngp ����m�z
wvn��SwZ� ��Mt��h+�	�΁k�h�n��PuNe�r� v�8�6�ܥ�eF�h�����2[��H ��� ݭ�t�hn�7S�sA����s� n�;��.��tV�I���̳�K�t`SK;6�@��������d(V��u�i���eU-��)�{�@��P[��SF��6h-��\+5TLt�vU@�ݳ�5B�.8 �r���@Ϊ�T���u��r�h1
UP(/��@{Ϛ}h�LU:�v7 ʍ[��-�U��CT�Ӏ�@��[p�ۦ�*�UmiTT�S�(��A� 
4�Z�4-������O|���� \:���l�u���ƇB��UU�uWYB�v�%T�igP(vi�n����l��Y�{�R ޾4)m�s�tQn�m�EwSv�Z��ns}��)�EYO\:�[�� �nU� P��ݠ����  ��
'C
  ��R�@M4��0F�T�1%QSC@d	�0`��2
TU` `�O5IP���i�a�� h$�JB
�� M42  ��$�0Bbi��@#j����?�������r������?�m��������ӝ�_<�|�ϜC��2�ߥ W���
� EO�� ��O�`� ���t	������gg��� `�I$��z( *�`xS�@��?��~_G�`�X����u���.0u��Mb�X:���u���]`� ��b�X:����]b�X����]b�k����u��b� �.�5�`�X���.�5��b�F&�bkX:�5��`�X:��.�0`� ��b� ������b�X����X��`� ��b��5���bF�b�X:�5��Xk0b�X�5�kX:��\b�X:���u��]`�X��Mb�X:���u��]bk�L`�X:��.�u��]bc`�X:��&�u��b�X�����]`�X:��.�5�k��.�`�X�u�kX�0u�kX��5��X���k0u��]`���`�5�1u��X�u��X:�k��`���k�!�X�`�5�k#X����b�5�k`k �.�b��.�u�k3X��M`��5��]b�X��0`�5�k��d`kX:���5��M`�X��q��`��# b��b kX �@� �T5�!�cX�X
�]`�� b k]`�Au���CX �X �X(�]` kX��]`��Ebk CX���
�Q5�!�Uu��CX��X�@��@5���5����Pu���Tb�k GX*� �*��5�&�1P5���Pb�kCX����&�P�(� ��@5���` k]`��Eu���CX"F��WX�� � �5��u��u�`��E� ��WX
�]`+�Uu���E��� � �15���U�(��WX"�WX �WX*� X0� 0 5���� ��(��
�5�k�� ��5���P`kX�� ��0@5��@Mb�kX��@�
�5�.�H� �*�5���`kCX ��P�k"�P� :�5��CX��5����X�b�X���u�k �.�`�5��u�c �.�`���k����b�5��X:�5��c`��.�`�5��]`�#X��u��]b� �.�u���b�X����]b�X�����u��X�u��`�#X��5�kX��5��]a�H���]`�X��b� �\L`��.�u�kX��5���.0u��]b� ��u�bkXF&�5��X�u�kX���\X��"=������W��"��w,������c�o]n�)J�/6�Jh��A�B��]C-,M6reka�LȈ:-��E*�ӴY{GJ�d��iH1�p˻�n447B�L#WT)e�KR*�ͽ�»���ZC5[I��"B�#AI
����[�{��Ek��-Ry+2�Z�wUVl(���)��`��sD0���u`&�H�,�xSP�Rm�Jp�
2�J.�@�.M̖�a��D�V��F�6j��J1c�nL�ڌ-٦�Rf&�E<8������.��)crPh^
�1Cc[0�q�e���ʱMȆ<�j�jM���J�#+�caڼ�ǭݪ��Ƿ���nM��̻�e��ڱ�l���#=���*�w��M�f�36��oLA�m��FD�U��7j��Ǖ�	�5��S���T�sMQ8�L�.e�s]�č�ZlQe�Y�N���}f�y����ZY��e��Ti�X�o��3�
T���N��'B���.��
Qd�]@��w*o�S�pSp�T
�x1�a�`�� ڳGn��S��1��@�mx�xb]�W����iXZ�Iz���SĨ���g7.�()���=�ohE{=�VY˪ݧX��,�#�E��Ÿ'I��`gev}�/=�/-4:G�n̍��Y8��ɻ�k>;��Gv�!�������Û�T2���9�5u��#6�+�����9��������AA�܃e�������JISY���W�L9�����f�6�L�-��p1t":�L�U�!P9e���Yq��5E]ٻoZ'rۭ�Ɋ�G�T.nf-,���71])yE������.�崖C�EA�Z�Y��Mfೕ8a)-�1����D�������ˠv輸0�rDc(� �&(),���gw1�A�[��8�j�ܣ��-^ʦ�&a̧K1U�r������W�Z�f�h��r�XEm5PI�.��Zw1-p�.���2D\V��peH2���Xީ����/Hc�˭qU�XZ59j9��y��L�SeX��J�s׫���F�tc�)�n�ia7kj��(*k6Vѽ)3q���o�R�m7rȕ�a�dŢ������;Z�]�{{����V���B$������3�%3�tFVP�I6tR����海�V���:�n�nޜ,��V�ٹ����UT�n#vG�m�[��q��E�Q�XY���m�ܔ�fm�tkN	���,׳٫N�-�ۉeSܓo�u���.dk)�p�E7��؉�u��N�#t��Y�fV��[enR�/v��[�O�p f(�e�Q	ͻ��k,�5�WVJyo�i#5Y���5�U�{)���n����m̈��Ӷ*ق�'L��N�&���j��V	ED����"٨&�i����W��T���,#��6�C�p�܈܇� V�J��Me���hMY5��S2�J�{*�4�lL�����{q䂯$Ğ�s�3B�/U�RɧI� kU���vXH���B§�ڠ&*Ȩ�0�j��nR���GU���o+j�ELq��;�Ɓ�S4�b+]�X���b����2`�y�Z2��B��5��&)�Al`6�����T滉nԍփV�j�b�V�t(d&9��ӊBKm�#R��V�!Zq��C���ca^�Vr2�����a3Nޣw�݌PKL��m�P�A�;o%ɬ�M�������)����\5�xT�w�I�&`�&�i$�U�]��1����R"�{�`���엙k^��u4��w�xՂ�ֲt1���� �z(��V?+o�wbi�-jT�Z���\VEǳ!!f̆�i;+%j��m��Kf^Y*,M=�o*�Kّ�"�����
.��G @�7�T�uٵGm�bb,���m0�����@�
�n��=H�
���o4ۉJ�y�V_��Aj�h)W-[��y4Qɺ�R�Yv�OT3͖�Ǒf݊"U&��Fv��֓X�ƆF�ޘ#�v���,l6�*R�e<,m;�N�ʠ��kfV�ͺ{G���SX�yS�uv��0��互nm���W�w3`�t�᱆\u~vd�HGc*�{��`����B�n���Tn�ۛ~'t������6�׮�2���Bedh]�f���U�f�zvƧ/,K���әf�2��(&V3[x�����jg�ak�doI8��5�!H�ʥXl��^j˭�-#6�fc�7cq��]�	m�Hm�Pa�[��Q�V���7X��6ƫ�p�
���׺�KcTF�8��K�.�AQ[6jfX+�.�S��s)�^�t�U��,�Yꦽs�$A�
��P�-��]S0Ld(�I�j˒��f���uB����q��7A��*�e���7*��sq,W����ǲ�UFs5�*�*���ٛf������4	�'L�j�f��l��Y��I��5VYʄE#�/j���r�l��j�q�ٻj^�"�;l�r��w2�o*��������GD2�Ɖ�j���\1�qF"~���ɂt�w�r$����E1��7uM%T [!-�j<۳X�PnZf�mP��{HZ�D͛j�R�ө�-Y���\Q�ɫ2Z0&w��SU�勗m�K1�˓LH�V��P�7l��2�	u��˩�X��#E�6[Ǳe�J�ռ=��R�gm:�)v�C�4J67w�UÏ^J���9Z!�K&Kw��,��[��dEz�[�\��|5�]e�AC=;#Y��E�e�[{��t��t��n
��)�$)5�
ݛ�vB
�l��1��i˼��kZ��q�*�ޚ�
`Ѫa�U7L�Y�1�N7HY����cB�/4�U��F��w�z,�y!�m-�F��!Tlfԫ�u*9���^�m��U^�l�2.��
�f*�3�cݻx�1�X�M7��kj^�m���ڳ2¦���36���@!أB<Q��Ie�M�Q��n���T,͹Rh[��f��3��{�f���Ѭ�X�[�W���b��Z�H5�`�0e�{�՛���.�;�tp��v�.�h&qSx�KsV�Q���j�<��n֘��f�&�PX����U�u��N��\��Ȉͺ<Q���Mke3w�S���%)�v�Rz4�b�k^U���-��K�]=YO%��/��Ť)����Lѵpe{f�M�z���ԝC/mB�j��q�]���V0�i��Ȧ↥ӳ���-8�ӱ��oSu�eYda�:"�1͒�Kе檔�K31����@���Qsb�&d¶R���YxN4nQ�V�l�x�'�3�ØMT�j���n�Żz�J�#V����=����Y���3-7E�q���*=�)�`�tdۙo&����w�7N��%�nax^��f�՘\p���V�`�ڭ����kH�kS�qm<�f�b���(�rE㒭��\V���fY'f(A�	FE�w��Yd�J�wEj�&�x�/J,/n��v�#xQ��E��j�4y��)];�ے�H�+1�,��x�2�6�R���NJH�-ؚיYZ�ҫ^�d��̚�KFA[I@�	�OT��ڽ^cn��n
9k!��i^���$�x��%4�6�pc��;b��"�8��܃O�&`���-GZfh2e;ص呋.�(�ͭ��5 �oa�[[2#%J<C�����פJ�كr�F(��\Z˫n �qj�ZO-[�ej��N�����G]��a!�kAB�:)ݵ4�MK��츶��<݂��g.���͈lx�dTU����a)Ja"8# �Z0i��maSwkU��¨�x�=y)͖R��QW@�w�~&��8m�n�Y-:�a��$��B/!n�nfU�P6�:2��J��Fk2�*E>C,)��	�ɼ�X��
s.��d������x�6F�Y��M���R�$����-"�z!ˉS��7xj�&�ͬ�*�wi��
ʡ-���*�/Z�T1��H^f8Y�\���1Q
��a]�R96��#4�.�VU�{~[��鱸��^��%(��06�C�(�ol��ss4\	�(���*1��]�CbVLUe)U�f�ҳ37vY�lm
2�&�б[�P�UV��7�(�~$�V��U��ɛ2TKux]<4�Wp9L\oe-&�A�n���܆SV�d,ǡ´鵇S�Y@Ь*ؔ71��Z�T��f�0*�a�Y7܂�!.�^�v�ޤ�dI]�M�N��Sj���Ӝ�-�S�������M���WX֛��ަkN�d��ݡb)7!'�ӑtr��-&�ӻv���3h�5x8�w�����g]�nY�5Gkt�$�:�j�K%�I���D�M$�.i�bV�,�bbʛ�֍.���81�a�H�S
/.Űl�]��D���*:�!�@᱄���)�(�[�Rjd剂��w�LA�{r^:y�nSw���7"��mR@��U5GU��7��v�U���J���u�&0�^�8M+1�*�����^j�溵�EVl޲�M�Z,���+%4��m�S-�w;�D�P���w{��`�6���g؞U�oba
.��,��u�Rm4볈�m[#w��s	xZ�y���K�&����Jv����a
� &E���r(�b�VCc)h�c^0��!h�6˄R��t�U��������ن��t�9�&ZGp9�����L������4M�&VT�� FV�-�sQcw׹�c��(;��.��Օr��hɰ��O&<U*�V��0�C���ά[D��u��n�Q���(r�q�4���.�%�s1�)O)���-�:]�Bv�<u�NֲmO:9���ʺ���n0�;[�'5�ת�-�"�Ь��Lѳ6MY�^/�P^�F��x2��jM��ӪaU�T����e�l����F�#�]�F�o��PTʻ{��IsU�֩Z��4�H;�]��7�ljVL7��J����0<N��8�V�e��%����U<	7	��1���;���z)�SuB�v���˼Z1I���X�n���z�i�U�"�c��#L�&�9=��.�:�Kv�Ů��M��o-oct4��Ê�E齋ƱF�L�����K�]aN�U7H�^a~ݡ.����,�n�!(2��L��ᄂPa�j���]ۭ���D5��3	Z+4JC2L����XI���V���Ņ�33ڕ�A��R��H��mAwaa�뙑TJ
�+h$*J2��Þ,d,C4O^4�R�,*��U�E
��n܋!�0�diZ4�SV02�j��dmdZ�H�QF�n�DE��l�:t�*�/�@�"9 7�)^9�1�f����nP��r���S�SL�Ns!b�Sq�.XԈ�O��booF��m�E�;��E�Oۨ�z���-��!�Kt%�p�.���ىi֞l�H�+r�M�Ad�?C3UȈV�L�+)�XhT�����Ƿ�b�{���s#�xӶ�ٌl�Ǘ�أ�&D�e�bʱ����DB[�{�-W���B�ݰɫ�xYyHTR�.͜rC�7j[��f�'tX��c,r�k%z̕�ԓ30�otX�R嬊4�t�c�Uǁ�ʎ�J��-�=�(P�Oel�WVb
��]��B�SD��Js&j��.^E��:�`#r�V�Xr[!j�ۣ�5+�y��K��ts�,*Û��aɃ��;����*���O.�n��Ѹ��{�3i�TA��v��i��S�Rd�ۇ,o"0������4����05tj*�WN�#XSw�	��`��.j�UQ��TTR�Cf����Ԍ�"�̌m�nXS�Xn�����Z�ۨ�N�a��j�E�t�$V]�Z�Q���)�#U'݁b͸�k�E�J�i@e�tRu��S]�"�g%U���۬#o[z��b�#��V����dګCpd&�����2�MD��+�lm�p^ݳ���XV^�T��2�����щX��NԼ�{D+ÃV6f%��U
ٰ��#Z�5W!�hM�L5$sx֚����l����V�s-�f�&s�4av��r�mt������e�wJ^l��e])���R��gNnc9����֜�CjhR��B��㹙3q]�ʛZe���Rm������꼗m���#�2�X�M;�6�$XX��#t�g��zZ�y0f,�Y��!�I	�Jô�ݹO`pe�
�ƙ���v��;���7�Ii��_�ṕj���c~����'Cn�t�cM�q�IF�[qG�{��ʓjjM�N��5y&!@�Z`�&]���ORT��(�3����]�D�l���ђ�E�\T��|�K�t�;��I�YIZ����7��,Yًvq.3&Lk�ż��cZ�.�1&�ũ+H�Db �i��-HdԱ$�Z�$A ��(i�Z��R+��R,�QP8�īQk��60SW=O{�H��\�.��h5�6�J��U=	8T@�]"���+kWH$yV�l�KM*J�m��I4��V����*�L[6�h+���Ϊ,J�<�U�"�M�J��Ҽ"�*��\��I�N���2VE�$���pfu�޹r5��*{�E�./���Ws�D�W���F\�Or�\��j��I_$�U�RդZ)b��z�6
Ė��J��j#IEڟ>:�V�E��(	嘊]�I�f#�5h6��@�V�D�mjQ'��}*����E�-�Ė�H�@����r�#]j%��"�kuTY��f��A�Pe�/
H2�����]*�" ���jMm�Ԥ�ֻ;r�T��$�#dsv��A�N-�E@�����;�Qb@�I$���+SV��H�.̭��8��։+��Z�V☓S��mP6�%t�]ԙoV侪Ex�$�֜E>桧8C!���@���|�/Z��}I5��ŗW���krI��S)^+��[T�1Mr��p$�|	�2�����I4�,ijT�]y�$�wK-m(i$A�=L
�@�X�I�������%����[i�Ԓ��]J4��H�m�G8U{��h���WjZ�M(�4�R�I;�{�5��k7ݓC\Հ��R��X�L�{���ۖT^T�2O�L���V/��� �ޕ��?0�������8MMm/c%w�i�i�����j���-�1�e�Y�f�L�Էz�#a���쩈�^�.�b倜}Əu i���c�嚹��3�'��n�;��3B���x�Uٝ�1"锲|�"����&�ٻ˛MbvU]7a�sMҐ��X��q�5[��0�$�HX���&��g��W}����Jn�%rIQn�(�[?D�f.dk���-:��+�`�l�Pg:��QTj�[�'�d�y�+��u,�ʹ&�v��*��HQ�YkPI1�s:��l�3�[�TԲ��bE셰`_�˴I&��̶.�U�x-�Ĕ���m9��7�S(HL=��fa��(u3V	�"�)�����v�B�9U�h׺8RZI��fɕ�V+��0���U`�+&ܦ�6n�S��.�l�iO�W����ܕ�᭐E���ƫ;�2��^r�3Nf�А92����Z�Su�A�7�����=�.C�
|�%r-��A\LZ�g��s�6TM���^#����k6s���,^������W���J�{�Y�G
��r�'Yn���C�zR�q'QC}�y(���5��;�^M�ԥ�a�ʵ����,�Ъ���Y����ۻ2�n�F��%QP$��8m]C�j���5�)��jj�a�B���悷���R
�5M�%e����r���v��i��M��-��o�ʸ[�f���%B���w��xs�{���)ެt�G���ma����s��h����boU�5���nSz�U�6$B�E⑳�+s��Qt��KJ��� ��}֭Z��3s/v"�/YY�˴�����\�P[�ɶ��t*���AWv�����n_i�۰왋/,�b�N���w�Xص&�}(���կ�ee�t�Nnj��9l�=B��ګV��n2ՙ�O~�o5jyo�m��N���,��܀�dbql��.��"����waR&�MUY���_S\t�WT/á�O&ff�9ҡ��Sί^�2	�v��+T4�MY�tXk曹�0^Y�܍Gv,Z&��໛+,=gN��ݩ���j^V[�2Xqt�0�<F�5/�MS6��U����V^��Y�"g ��V��m�ܫ���#qi��!#H�-�����5�IR��rF�k�ܾ��l���fz�����\��ӕ���HI�k�f������d�&64e[�3�`�j�j�7���프�<d:t�:�N(�	9�3B�4ث��y��5r��G%�kmLarSYHgn��),�bB�N:}W����3k%Y��������ocZ������떆������3.���ӤZd_g)ֆ̀ڹ�v�%�hr^��#V��g&C�-�M�!V�M�����77{�õC��pK��\���̬O�=��O3�mR�\"�[�n��r��c*�+��9hVl׉��ӛ`�+ �������O�x���k�WG�V��I�&�f5�Ҵ�,��`��m�C[��jIe�!6.���X���֫q��+�V�ЧrX��)�ܯ#V���9b�z�9^c��O�� �Av�*�=}\ָgP��c�s�����5Ԭj�ƍj����.Y��l�q3E]օ���Ě���oV�E`�7R7��+�+Ѽǁ��b�w�_a	=��t��=�او�ģ��T�U;��j��̪�,�p�Y���Kun��*�|������CA��W�'mS&t܊wa-*��%�ŧ��B�㑆�����p�Y�ǂ�v�T�e撋ɜ
�91�cW[�!��Ț�V��շ0q9X�K��M��uhe��X�뜈Ie�9"�S��VT���;B۾�+��K�Op���N���Y�tT���A���TJ��N,ɗ.i������vޑ�o&�i�A�*1�=��6ҡ%c��껝;�2�v�B�i�@��c���U�ϤL��*2#^]:뮾��BwL��)Yh��u= Ú�����U�7F�r2�1�u��;Kn�ާ�Fa���p;�_`�V[tR;I���ڛ��V��� ��i�_y;m7��(w�J֫:��r^;7f��<��S�o���=j"�̙tl�c�U/�o�U�cx�u�bx��q�]�}��R��D�Vኖ����k\��!�5FV�Sq��]?��������;-8:��j��O9�ɢ%�ջ۷�,���暢�$�R�J��.��w���"�m��ԛ�d�F�1��>�!e8�fS:*�.��ل3��N��'eA�2��ӫu��Ė�cf�����+Ғ2/g1�4�,a��
4!H�/E�H)�X�6qă͕W{��(^bW�.�1T�{Bj��o�+�Rdn!r:	'�U�D���Ь՜��y5�e(u"�0�۷�N�U�����������d��BSW+���X3�X��]Żک*������wTOfM�";��}nq9�;�Ŭ��)X0eA�6K�*�Oj��|�谅��M+���۷S�qi*�h�a!h�d�A���d�I��؎j����B��TV��Ӓ#PaX�sхJ��fVp�Hn���U�ӫ�.�87ys�zn.�N2�f�J��U�I�����z!������X�Q+ �}Hٻ4aB=�,T��l�H�Yc�G����Uz+�s1Eΐ���$��X;m-��Nr.�])��:��F���l�3�0�X�׆ �M>�O�`�v������}E���X���7�,]��r-;�kz)�RL�<n�Ϊ��J���e�*����]�ڔ�;�{uG��Zb�4�[�¹������Y�8tw���Oa�D�e-kebp؇O46eN�Ɍs��W@������7l0�Z�_b�YN��}Ԣ��ȗ�";�#���'on	�kh&��v�I1�Tf��]�����m�6�7*U�БZ�	5L�iP��"�ѳ0���n�.d�����N�^��8�]��,}�*g0��v"�w%lt�`ӷ�W^vcN��2s��r��'j��z/a�B�ܜo{oǳӫ�u�:�sn����0uv��ʭ�˲�n��N��@�=��Uki���r���v��������f7yx��jcv��%'D�߮9�2���nl�mb�;�ۮ�c��gz�Dλ��Q���}1Í��{lI�%��:�E<s��)*�(:�ydU�%g�����g=�̍�e[y�f���N��fu-ٗ�b\�����=|M$�4��Ĳ#�̇3����R�gUP{��Ը%��ޘ^�Sv��,v���ko��Ӂ��q��X��4F��%N�gt���Oo-�jj,���Z5d��']���)�1Mb���l�T�l���3o�5pw`�6��Z͜
�bQ9gmS6�ȋ?%��g~�f�/H�c�5Qi�\I�>O��	1�tK��2��Ov䌨���lMJ�7ara���3e#�	�9��ض�j�J�F����R�f���PV���&<Ӳ�n�j��6Ɯ:�5�n���,�%\b�&�6�.�b��8�l��[�K�%C'"�����ӹ�Z�s���;��r\{��Ҧws��*ūۺ낲�o'z���"S�C�뼈m��i;'(�^�+�!*�r�y�.'s��{a�S�
�P��{z��ֵ!�������|�+�(�=�cx�&�T�WAB�v�q��&��l����Ĺ[�7:]s�|�n��:oU=�am���.��:]��f�����#���e���"I=���k6���M2*ve�#|�']2{xNUy��R��cG�xք0ދ��������]FoCy�w/u�L��M�V)V^U7�p��m`�V%e��\t�OrA��ʛ�8Ru�u��%L���U�ЋIQ��\�L*���Ι�)*N5`�w:U��+5�r�ƺ�Ӽ�{$��]v ��-���
��K�y%�;!|�J����E��y����5��q�T�E�))���,��FN�M��2�)��b���e�|U8;,N��Qq���k1qՅ��_Dt�8q���N�\D})�T	i��;9�Ψ*�ZWWn�8���$�]�N�-t��ˬ^��i��:�Jz����oIs{yse�h]��o�AA�:es���ɚ�N���1ԝ�0�RXr�Ǩ����;�쥥bʬj�^��%tȻ��K�˳,Wr���v�}-TC���5��u��}��iփo�F8a��ABŦj�
gU�,����I�ݍ��V{��eQ��M�Z��S%c�o�q'�����ɐV��&��2�q�,H^5�.�;����݉l��]ʞ�7"�u����~��@�ʝ0�d�^���V�:��WE�2��*3��i�4�T��'4�ӼF��х!�b����yڸ�-�tBZ��!SV��S왒����M�R�1k�.o���z�2�<��g��ީ��ʨ�t�6�-���3\#3���jE�m̜CZrDI:��5']�я���Z���oKRڬFq��x��fh��әn�)#UV3p��F�a��қ�voA��#�륚�f՚3!Y{3��R���gI�4�in�*�k�Zٌ���6PP�传�Њw�\"�6�N�cGS��9�5ӛ���K�}�]N�E�g3.Q��0�i<�����Z�^�﷪�2�FҐ�8˰ƻӱ���x���-�J�頬�6�.1("�Ĺ4��X�u���u²�{].��Z,��3;.Ц$MXƉE][S�������Y��w.����/4��D�s���*wm��5ka_U����=�Vq#I�O,☒}���
X!�ra˛����R�:�K2�������m�6��5�.C����;�}��X.��=|��YgҠt�i�ܻ�XKy\*�,	әe���6��Vp�Y�!�z���G#�����ݪ\�4d�ۦO+hNu"����j�Ҕےu���S9'Z��k��������$
q��Wg��.��	�޹}T� ���;T3�mXf��ڮ4n�5��|�۫c1��r넍���Z֎u�����>��9�3���[*�����n��z�!�Z()8�\�o^M��R�t-����WJ6����('��KR��h�6��`�$�E���"�������"X�Q3��X��n�.A��z�;�/Q���Q{� 7"[�Y���q���/���V�lS��Y��[&�b�S�[���U��(͕�.�ޅ��&��(�O�N�.ܬ�"DP:n�=LZ�;X�ݮ�2nx��i�{����&e������r���0�T�h��
�[ہ:���s���#�X������!�H��D׵��CYa��6�Ķ�����w�q|����\4�q޵ʕu�5�Iu𶲗 Ւ�"�t쭲���Kj-B�vA��QGv2��N��Jr+Qy�V!�!»b�y���i[i��'	��z��]��2,����u�bY�N�$���}����+7vhx���j��M䝊É���p��1�D<�X�SC-���.�7A��Zn�K��Tsi=���X��J=�WUD�7�Fؑ	�蹓�VKm��Y4j�l�ڤoq�6�l[�y������v,�l9e-�N(�)�,��e��ۡd�4�n�)<;)m�R�G�b�a���f��w[�P��*hܘ�A���0���6�*`׭�r龬��Y*�q�R�r�Q�q�ޱ\:�gS�y�b����m�����q�&�\�	��]�u�t��hފ�t�l\��3U�g;�W-�̢oj\�Ǧl�;;�e�H�o��{x$u�Z(%7pZh���̄i*#2�l��#�0�+ɶ�L�؁B͹ۉ�ƴ���E����q�v�WD��j���I����XJ�9��ѥC�&�=���9�*� \}¨c���i.4�PΤ��j3j�l慦p�"���ղw�h��N�f�����(5��K�q����0^,�/ZMd:pu3�!����9UVqǦ����Zս:��k�M�o�,�����B��*�c���r����&�ڃ7�Yr�/-�N�-�wk3��n��3v�5�<8����t� u�7U�-��Q�Q2/q-�.ɣ��'-�;:�T9��~��E��%�s�Tr+���bM���t
:�Ub�5cwtT��ݳ���]o!1�U{po7G��%ՄT^� �[D��n���mL�wy�Y\�)�uE�w���g7{�ø�\�׫��a�o7�X�Tڬ6m�x���ʓ���b�T�*�wf�E�;�Zrj�J�����{�KN5��ӷ�5�׼����WuY���ݛ�e�r͒�4"[L�[m��{�jwM�ި�w���%�:��j��}�Ǘ̻|���;��1|�qE�&ÈC�(w�u7�y�[�us's�'�����ω��ǽܡ:vc��<<�h�In ��&���6�pb u�5p ++(T�1xѦ�"r 
�V����� �F���&ϼ�$ H�� f7�,�1y�Э^������#�ܰ��(��I
�l���[ND{߈��ٶ����L�$������j�_K_�v�x�zW/j��p|��vu����������T猜��s�	���$�/x��J��<�qxxV*7kʛ��aW�����Þ�T:�L�r�"(����߿�P����/���S��`|UAs������=����O��OԿ�q�T�c���\$@K	�9
Vp�Y��s�MP��6��#��u�wX]�jֆaե���-];�R�r ���hj��!kD�+0m��T��79o�]+�G3^P�����y+�MT��*8w$�ӊ��]aY#*�Xr�WM�Z�֮�sg@�Y0^jT�Ğ��;���*U������s&��G|�]݋���a�����r�D�䶚�0�[��-{[fǔ�s&�]1�_�&���+$��I�����5uz)Ӓ�h���s���y�o��jި�߶f<ۥ�m�=�}�o��]%N"��0�U�]W��[���v�V�L�7��y��}a���W��qgB�- ���/�^��uf�[��v�'*ki`zJ��NQn��2h]��4T{�N#��f��;W(�8�V�uV�[�:�wX}���2d쎛4݋Уj��(���HN���f�=���7{;�~�TJ�ht�v�-�sZ���:6n�Ǖ�k#@v$�]���X̘��'�7�Y�8���x�ʺ���/�x�'y0��*^�t�΄Vbͷ |��
-�����[Wc�F呕�:Ҝ��6��-��u�U��۩P����f����u=�A9Eni�Y�ͬ�na��M�Ԫ7���T��Rod��.Qȩ�7#V�D�/���yz{{|zkZ�Zֵ�-kZ�ֵ�k�Zּ5�k�kZֽ5�k�kZֽ5�k�kZֽ=5�k�kZֵ�kZֵ�MkZֵ�||z|k]kZֵ�Mk]kZּ5�k^Zֵ�ykZ׆��k�Zֵ�k�kZ׆��c�Zֵ�|hֵ�kZ�Ʊ�k}��o������YW�%���MB��@����C�IS7����_kn�Dj��#��ڽ�Z�	tP.�4c̏HUG-W��;ۙ!]���ƅ͛8$���^ֺ�\�g�����uF�c�]^\�h���7vʆ����%䍵���x^��ۇtp��"��-u�+.kzSӷ����9�P�${�6J&d���za��UV/�f�F�[Ff�:���r�Pb�/^V]�dɫ�����*�!��]�iV���}T�Ks.��Le`;�f;,10T��?8&���5�9��w���������]a�k�M�^;.�쳎����D�+M����]��Y�j�GKw|q=�2(dd7��=�+"��tSY)\�����6&���W��n�����a Ћ�t�e��b��Oّ��{�y�݌◶� @E�K��8&ȥm�[���S��2���[l��L��S!D4���Q*�\�;2��u1�t٩WP�9WӶ�qw]:�<�7n���:���F�i�����ݻ5W[oL���`���;,u7��ڱ0�X/N&�!�q��S��'dP�o]�A��Twz�e�:��ogcܲ0G0<�+W$Nؼ���D������S�%F���T^q<��7�/]�w�z����ǧ�Ƶ�hֵ�kZִkZֵ�{k\kZֵ�Mk]kZֵ�{k\kZֵ�k^ֵֵ�k^��5�kZ־5�Zֵ�kZѭkZֵ��cZֵ�k_Ƶ�kZ־5�kZֵ�mk�kZּ��k�Zֵֺ�k�Z�ֵ�k�ZƵ�xkZל��e�}��d�1@�<��#�F!�[��$\�%�nJ9�a9�"b�@V
�n�E�8EtN$ �2j�QnѠw;�(��}oiֵOk��MI�݉��κ�4�+5qO=�oz�\��K)�h�o�V�q��l�+g6��dE��9`��h�2a��WER�ꭩu˺W���q&B�2@�.ZH3�2���Q�u-L�����	���i&�-��U�4�q]�^�[�Wl;y����9�^�UQ�-��Vc�\��-R1����eT]��TB�3�j�gmUn]dx�avfuj��oU[�	���r���1k9B�*v&`��c�ʓ)[�nɖXFƘ�+^5����
�Q���SO~��wmBp���Q��V�(q�VG^��eK{��xv�+lA4�ە:�lb���qN[Rͪ�J�f��&��f�xIT���n��hőPrh<���z�7wlIIU�r��,�)C6�ff��cl�ݒ�έ����g)݋�9-x�ͱR��|�ɹ[����vcb,T�˃���h��Vtī(�%'�u�N���o�J��(=������,�1-G%0Tζ�j";;#":�
|	�s���kTqV��yݻGr��]LŨ�j��1���B�l��QPw"�+2�E��|u���{||xk�omkZ�ֵƵ�kZ�ֵƵ�kX׶�kZ�Ƶ�hֵ�kZִkZֵ�k�Xֵ�k^�ֵֺ���kZ�ֵ�u�kZצ��u�kZצ��kZֵ��k\kZֵ�mk\kZֵ�mֵ�kZ��5�kZֽ��5�kZ�ֵ�kZ׆��z3�x�^��/gfT�[�գD�6�b5םm���/�-�i�\�����(˻vʽ�T���3
�0ff��4�oZ=.���*}�9����+U�'J���GJ��w	Jv��a#��v��n�#��U�P��<���3��{ǨЙ�[����W�N��P���ۍѬ�dX��435o	��r��,�].�:��*f@�V�.}�&U����نE�]L�N,��6;#Oe�={�/�*Wn�N�^��.�	�V��i9Ĉ��$���R�V�{�w,�t�{�v�&�q��bP՛D��̈�)ilv!ۗ3P�&��V�-[�x1(�)��Z�A,��c��K�4F�v�l�/[�V��ik�F��۹������E�����@��Uu��#"�8�n?����l�u�(�mmK9��ĭjٷ��/����Z0ouU�E�4�t���XYMV�}T��OZ����SH���Ƣ�h���%v[��>�g�ܚ�R��IgH�yM����c�k��"�kf�T�H�9��8ofS�-����d��y �&G^�̘�J���.�S�V��[|:ޤ9�s��%:�ke:9x����t4e�C�'ݡteh4��gUU�Q�;'i�m@63F�a�UGK�t��n�����C�'ُ:�od57eD���:ߨ����V��gbQ6�W,+�bڑZ�Ѻ]ٕ-ESga]��C@��2^�^�)R�-�	J�̝>�P������k��K^Ԯ��-�g\}�*2���u���)�ͥp]�Dá%�T�1p�������@o�F��Ɩ!�/wwE.�:���.�k�K�bw�G����i�U�}��S�Y|�}��u@�oH�m��3��\6�#��U�"9I�򇷺R���:u��Ow+E"enlɨ�Q����w�ȅ�Z���I��YCN�$[W��~����L�3��!��Tѝ��w5Ba7�Ǵ��E`�Vꆂ�KV�=�n* N��$"N�h5��NF@d� �]�5�c.
��B�7.F�ı YF��1�rl养��R��ǋ/(n���ʨ,W�.�f����S'���Pe'�-�ue�ڭ��]̻���t����t&�uGd�[J�yc���n���ۼ�;��N��xlF}T��$z���W�R�hj��dVdf����E�<�t���M{��6�����c��w��nd�������yN�=uhM<�t�yk%��㺴,g.o�*C�i[��������y��Qԟ[��ӗ]%B*'4��Tu�T�����Ubn����1lu%J6[��9:�w�8<�*=zkMU<��h��(�C���=B�w+�P9��[<�jZN��ݎ��Cԫ	c6r<���h�%�z$gmR԰mv\�^y���i�"��hG���ﻲ�֣�o�A�kp�O*�b�zR�1�0B���ʐt&k��2u��mѲ��D(ц���@xK��-�*{�c�3~�gS�9[�ݥ��:���'�!OE�����Aͱ�fí�R�y�s}�R�v�_V���EBUM��i5�Y������s{7�n�Lٜ�V�,���b+! \͐����ǔ�!���*۵��&8��m=����K�D��}����ʹ{�����xQ� w��^n��x���+�kz��
u�as=|(��]�[d�������,Ջ��ʻ��N����/�oA��۔$����g,�3���Jk|xX�*�=�v��\r�{
��Wp�UUD%&��P����bf�EQr�B0��uFhXw����1"^��J�˨<%T�7�c�Y�TЬ�nh���KV�|�� �gv��F�R�a��3��#aQ�v�`xE��Jj�.]>��+�2���4.�(e2Gr���cU��=�,���
oB5�c,��Q�x��������N�魝SbsRovf>����u]]U��qx�"��E(h`��썗�^^�G�ӝ�:G��?c��.���S�I[�T��zc!�u�a��w7F@���a;c��l���x�Y�C7� b����gk�t_��8�X�rڧim��ZQpK�b��[Z���0�d����c[sw��Y�GYƝ�s�e*IP�j�1a��l�-�{S(�l���*�.L�ʄ�����J�H���FȽ���4�A���rA����yU�F���C�*�Ы5�
��ؽ���c��:5�Y��: 	|��8������'`�÷"�[�vc�Q]��r&%����r���Y�z��7���yS��}�Wf'q�G8���rG�u܏����*�t��ov�,>4�X¢�D��)r��^ u%�v���S��-��+�.��T�v���lw�U��X�cn��s�)`�t��
��u�5VLR�zFV�� ؉���t���U�ݛU���{-Y�o��\gkqju����N6��vf:�`�N5Ihx�7a���F�Bm�%л^�a�����������iNUz��t�LN�b���i�u�P�'pj@궯T�AaR6FΧ۲���\�^>j�m��4]��d�
]����d�Y����d&�a�8�! ���:�8ɳYgVfH�c���s���X����f�H����P�
Z!��uuSx���O�V��7@�B�ͤ�Ŷ��0n��Si�3�V ���S;nШ<h���N�e?=K��a�)�u��6�/x*���f'�ӝ՜y�:����鶳ku.�sJW�4���L؆�^�oyn���(fI���Q��v;�����b�=W`��u0�����*e���;��ꋲ����ɦX�p[XtB����v�:S���mgl��X�h���ܕ:�[�r���6ōlK��6͔S��^�x��24:;W�k7b(�h(Jv�zq�u������!M�ngu��S��^�Iz�n=��ͽ������a���"dJ���fm	�Ww�p�*YwzrgokʼV�4h�x�Oh�Q���[wxޞ��_s���p�z���s8��v��=:��5�(�\���?45�Qٛ��/�N˾�kVЦ!�L��܊����y���k`j�'s����9�����>��FVm����I@�w[QDН��َ�`:s<f�����t9�P�d�4��5^�����ThdR*�\yުႠ�Ξ��).;�W�,�]\z���2Y���-ЮXs��C��u�"L�h�������$���ua�XL�6���É��k�pô�L0#mg���Eg�N���˰���w�o5��:�k���	Xh=4��3tqiC>��	m����Tja
V��UسN��Z
�S�]��Q�x��s$�Ȇ���� ��v��\bt7[
ĴJ���I�bƙ����[���s��V����ؒC�z��Zo�YV��7%�xʘ�&zI޺n;Q����<=+��K�X��4p�s�.�UP��嶹³j�AX���^���M^q��36���s�����IfQ�t�������bt0m��5Y�Yԭ��.��cQ5���My���`�0�]c��T��J�����dU��j�GEٜ�E9���Ζw�lC���1q�w��Y�ފ���z�WVh��:47��ƅ'uՐ�VQ��v���64Qx�Ğ��1,�ۢslk��+����ku[7�8v��>�[{-ʃ`Sr��w+2eћ%�k6�fG��Y�-=�xtȶD�!�UB�s�{0�\��'�9�rS�Ưz�VIfւ7���X�#�'ٌރ�I��i�N,�b�)��0�ȟ�҃���)s3O;p�&dS�� �b9v�Ƨlޱ7l\�%Ҕ�-�� �*�!E���\�e\�R*��`�PZx�ˋ\:z�vꐲ��sY���"��!����v�ݝ�%���Q�I{&�_<`�����#^Z;͑6¾����z*U����/V��!]�E��փ�I����#��5�m�'w�ޥ�F�b]ֺ�P�]�7��2�{5V�W�U}TU�R�W�����V���<b<K ���V�ˣ"�(\$tv�윳)N��r�ugR�{�LVqw69����E��A���R���z�o^�`��B1e&��NM�����YغĖ�n�$ɱB�J�Ց]��z�ǧ0َmaZ#\  ������u��(-�w͑���i���"��]ChUѕ��sx!�q�I0�$boWl�c���'<�]����B�@Px���ѫ���%,�b�=[�tB���B�Nj�fYzy �N����%��5�J�;�*��l�U��.�V��L�	g���º$d�bu�G�QQ]iX�������v,��뉮#x������k��ԭ^��:���Ҽ���3tjoSUL�Qw��Z��l��ghX�0i���k/R��7���2h�e:V�1.V�M^�`�(��������i�Up�D�F4(�H�+�s0:���uV���.{R۬B;��/E�#%�m�}����hw�L�7�7/u,�Xv�C�ޜ��LE�٨��`�"rZ2��VnD�����Ţ��K��̝ئ�+q<�7N�ЛOk|�m�Z�+�DH5;\�8b�U{p3��^
9f@�w!�}B�Eڶ�sh΍�X�<���W4'�;�����5>���Fb��ň�n�O�Xl���O�  U�����?�����/���'����$���e� ���.0�i��D��
Lj0�6ۉ�Y�J ��?"�$�Q&������e�DP����Q�A�HnD�0�P����I$�@�8�Q��%��C�-Bbj�A"�=J�H���^Lȉ2�(#E"Q�X0�c��2:����0������Ȓ&�`��ɤ؈�
$�C�Y� �>e%�C�F��j�*�l������]���X��7����noe+-�k�v�KG8-7o���ȉ�׬ӗ�³lsޝsp�gn)N�k[u�{yp�:g]�L���;XRƲ�t�6s��	��,�5 ��_j��V*�b�S\��ճ7mӝ:��R�S���<xm��B���et�=�lm+];j�K�I����sb�� 샊�"t^�v��b�f�5�� B� �+Yu}0�1�O"�ƶi�d�h�j���t�p2�ҏWWX�t�U��R��,��X��qlRY.������IR��HjEM��%��z	��+�u�w����_�"U�sH"��X�7���YT��K���k0B�mf�nj�87mD�KX��|ؙ׹c%TD�J��Ў[���*��ے!gh�x"$^�P���d䵸�+:�o]��ł���5W��'�T��KB1qVFIg8U�X���i�/�wH��t�-D�9Z����q���FjL7*�M�l�ZC�sr�ظ)9J��IC��������ܓ[�*��%I;�׬��v+ژ�U��k|����֌����xҪs[�cK"���Q]�Y:j馡��]���γ�\�ܳf����T��j-���x�����Cn6��wo:���f6�M�4�l�a�\�A�B�E��"D�% �*7�X�ȋJ�N/B�L?(���!Q@�-DZ(�*��R$X���B8���#�!$��D��	�����I�W�,2� ��BBb�B�������
" ����N&�d��G!1�5Q� �Q���R�1_�PH�@�m4Xi��qzHP$6�!�,F���F%&�E�:f�����*�8�I!��`��
�c��$A5!�2Ϡ ����b�
�Zۑ'-D�Q	�2��$�bQƒ^�-�l��RBC�"C� �$��DAnFN&�i$D"$B�z��I�)��i�dbBb�C��)�
~nA"!��8�bI �Xz�b�J�>+�]�w�ܨ�ޞy�e3Q�
�Q�K\�cb�nޞ����ֵ�kZ��Ƶ��$,P��y+ǒ�t��$M���,QHj"Eֵ�k_ֵ�kZ�5�A%���X4JHm(���W+�s&�(�2,cZֽ���kZֵ����[��&�ZMAfDY7�v�K��J
��м�_�b�F1�уd������@щݹ��D���$�p�݋��.�4�u�s�.�n.�\u]F��� ���ƹ�suR[���6�w\�w*�srmD����[��v��ERQӺ�X�C��s��wE\����+�����r��d�ڥ�����t嫝˷}�槎�t��Ns��{����f��r��]�#o������&�]��rݎ�J:||�/ZF�嗷λ�]���y��<�ݣ�vW�ݥ���w��7��Q�o%�+�<Wr0�}�x���O*A�ty�0Y�2gw��Q$F��=���>���Έ%8Y��j4"��*%a&&T5Hҋ�(�c|���bۑ�׺��f�v�M�8��۩�yj��y���dn�m�^�{b�L�Ś�ԖcL�n���S��(�B�B$�&&"�4J*Dj4�^L��MR*�(!��$&Fى	�$�Ćmȁ-cLկ���< �{��{)!U��̧׮�I�ƪ&l�Pޑ��󕙲�xl��Wwa�U��m]����Pr����|W1��}3��i��: ����}�W=�h�y5�Ls�P��Itٕ���ۮ�Z#��|^�ő=~��ٵ�W�O��ޅڶȷ�&�3{��	��11CJy}����}b����D��tֻ�ٍ�d���ݣ��)F��$B�'�]0�a�_f�����M*�b�+q��ggh�}��Mۿ���6�W\��4%{@���yG*��b�kU�g��`�ݎ]*�THF}�P9L�P�W�r�7I�#J�E�
��I�Z�07ί9.��ߒ���pv��h4�vFjum@�~��jg
������C�uR�#�_GMT�žEb�ֽ|�n	'�;�@�� Z��Ɉ���3��r���
Ѩ���қJ�6:&ʔ�+N�Q>�ګ�fQ�i�\�m�Ő矿q��'������\�1W��ؖ���Ԗ�5�$Y���<��4�So\DE��M32���2����働m��F4��ħ��N�-�9���oa#��oMa��?L[��� ��zj6��e=�߆vg�b�As�4u��F��;�����1��z�p.�����ys"��~?��;�]Mv<���::*����ޥ��L]�U+���.vPmM20�JَPᮬ�B�.2�V��NU��W�p�@�Sakv�w��z	��u\�6�E3��4�}S��}�b$mp��b�d�����йu{�>qs�v�O]m��Bh�%-��<���U;�ȱ�����;	ݚ�1e��ʝ÷2J\:��J6�1�H��D7�������GbV����]6˙mK\�_eq��a�yڞ>�S�+4=#G\��h�P}��+���>9��v{{'����q`U��ʢ���1�o_��i��Kp����,��)+}����7���#�s=b6�1�#�n�bz��S�l*�ob��)Q��xo.�ݓ��j9ݖ;F򣢉�T�¹��V��]��ı�J�Uz�����:���:#�I!l����v�T�Uʿ�7O�ݕ�,>���*)v�d���0K�Ũn�Ί������9\̾R����>y�)1X�`�N���F'��B�a���u;Ͼ
���ֵM_.b9�])s����sG��!}�S���Ё?7s�Dvʒp�����W�9� ��:IfD�2;x��:O�p��R�A�u[�&	VOq��B
�i<���j���w�@4~����w_O�q�e^���=���4�f�I��s�.ܫ���ڑ��ro����BN��!,��7f: ���+�Q����$!����	��7b	��7�%�!nT�B��Iu��y�U�y� �G\��۰�t�����VK���:�Y�]�g:��	�77�pVm�s'�T�lZ��c;Lj3)󺚡{���܋�';�*6��0�L�%�e�r�{�o���Yc�X}13��Z�y(p��4��4vFQ���c�D7T!nҥF:��@]�t��x�I24���&2	�o;(�-��J���H���ؕ �53�*�Nl���4�#f��X��5Y�3�Nѹ�Q�f%�1$��ɐ,��U&�k�y�8Qt�e�����f�<Uˡd3�SPm�Hs[��2@`�{b��ۼ;�B���/��;c5��y�
6�@��))��#����ډ�k#&�K��Y��MW�D�ѽ��[�܃�]U�]���Qɗ�A�PD5���+�=>Uޝ� �?��Zv[3ěc����MS���9�l�Ք�Sg8��ԷF�'�xuYB��z(f.�~9���wvw�J�TF���ݹ��j\9�p�F4�=B�D�}g��}������9ϔsq���_+W
��4�����?8V��3�s�\r�)�:��tbr5���ژ��ۉ2�r�=�����	3ٛ�6���n��T�F'����Uq!�Y��*��a+//f� r���suV�I��R�>[�o:��b	�w��.K�6��F����3`>{��q�w�d7gb��ͦ��ߦ�!8����G$r��\k
+*��Yu��V��H�Gqn�R`¸����I:`Fkō���Ɏ:�=��߽o�Z��0�g�Ixfe��r`��+s/jS���p�PP߱�
�m]St�En�o^dX;YI<��Z�}��!}̤��>>>>#˥��{fQ�'r1����Ę�&R���'vڪ����,3�FǊ���=#�����}@��۠W��պ/�o�����{��o1U!��O�b���Q<Q�{rw7���m\seb�+^sp�V��o7{��;�qVJ��X>cf@ഷ�u�N��ܮ�5Y�v�r����v���zC��o�G1@aΰ����'C��T�Qu���!=�50$�7�'g�R������y�}��4�*嚋��Z�ᘓ'��d�y�	��N�ήޣ[F���v�}؝r�q����2U�\1͈����G���;`����=یY�Xo>s\��&i�{u&_^��}mbΓ�NO�$(��S��f�Y��<}�٣�d��W��!�hл���n��f�w\,W��!�>�G9�����z;���8��3=(�)�1�pm��;��W/��M��E6��)A+a�Bv�F�p:~/�V�"3<��\Rꅸ��	�TD<4������D"
X/�1��B��y��Ug� j!@g��"� nb��ǿ�Z����a�º���7쳵\ƫ��1�,$�qs���r�i�A�dl���������
�m�p���]cE�֪��壻�.���R�C���52��O��OPU�O��ZX~/ b�:�人�_v���Fԋ�ǧ����E�Y����t oܷ*��������`<��:bv����q٫<����xf�@�"���=�j�g����'{�z��=v��xwd�r�֠vp?F00r1o\��a��6�7V��,�{J�{D��Ɇm�d[V!���pvF��k���4%Ĉ�t!����a�����_x��+��(22�3r������0.z�^���g��qm�wٸ�$N��H[������?aΰd�t��H>�<�S����cv}�E�2��whi�p4��j%�,����3�D��}��9��GUя0��P�9ϻ�p���xiF#%n��F��4�]z����W��1�V�B�RI���5*����̺[�*��kOتQxhD�U��~��q2"��$;Q{t�*��)�8_w[��O:�,<��jpa޸�鞚S���Z�=E-'8�pfn��_C��>>>��¤�˽�me�{�yۺ��������C�F�=�ZCT:躜9�}p>�#y���ˏ�� f��o
��#[���FF�:uО�H�z0>ێ�|�f������s�;<���P��V�.�����;�<o\E�ՙ3�3t�6���Vv��p���K�}�)߳��vV������uua�3��>`�p�b�8��b襭
n>���9�jT���f#�[�'L�L���(5h@�	�6*�V�g�9�γ�H�eѳ��t��O*��ٵ@~�Ő*�68�DH��Oh�5$��x����9�Cs����f�j���6�բ.A��L'BA�P;PB�	\��/���|^�oc� j����:%���k=F���tHȝ�b�� ���k	��{���J9�؎��;o��;���ऻe��t���]�0|����!d���Y���^���0��s�ݮ�3V��Όv�ܩ�4�8/��]�Z����~g��(U����Z�.�\�C�ޭf��)����.{G+�r��V��/9zFӕ��yi�w&Y�7���pW�1�����ʭ}��TlĈu�nT�oeou�2"�-�m�A6��hn$�!�����
_B�^u=Dk��I��������]�!v}M��Y�(o>�tB�̤eoSq��Os�ؒW�����Tu�A���T��i���|v�U�	:�p�`�}�1o�˵ʳ�ۨ�y��&��-�T���(�+o���/F���wc5��yҍB;������kuĪs�ӝ �q��1�.�m�v�5��`a�42��v'�QԌji����$�)�vn7������9������1_ ���I��\�=ܐ�xcɩ7�<��槻����SA�OuKVP�*)+��ς��׎+��YMۻqw��Ջ��:��qÜƎ��$+���,[��rl��Hߕ��"O �KҗGuXZ�aBÉ�WU��:U�.�Xx�ʙ�9����:ov�ՄK�}O$��X����1�
�n	/n	���oc9�*,�}t�7X~�w�=���I$E�> ��|A>'���*�!��.�4�/�:�$��Rr��@�n'��U5��&h��j�DK�pV5k.1f��\7�����y������ڷz������7�ڕ�Η�����np<�[��|�3$�����4 r�P9�aWQVq�7�ީ�|wf7��r����r��A�Ol�Å��Tn��>������F.�	ܯO5Ӯ34���C�5.���u�@冹󄦭�~�M�.������uH���X��rPՔ���4��a�LZ}���Y�t��8��BSh#�YC��n6�:�X��D��9F�����{zL텕��ܕ�TF�]�7��Ɯ`x��Uy��[�<W7�5-��s��+��h��X��D7ܚ,<�徍�v������6�>ɡ��׷�
�%w��{%GP�0ܐ���-��'���{�{���/8K7�+iNty������v_`�f,�W.�#�+6���.۽�u����'+�t8ߍ��{�l�Ok]�W�4IJ��0�P�Ė�
+6.��Q[�d����v��P_	w����X!��᧦�X�Wׇ�+8�m�:n,7ll��
m�{id���� �Z	b���	n�)��U����D�mۺ��]e��U�;\ �� ��<7^�s\(�PL�r�	��Wׂc��9�͹��h���=}��W���$��y�7<��!Fw8��f�,y�u2ձ�EL<a���S�.����V�wwyz5����	�v9ї�Z�0f��lXYǲg������q_�M���l���}��=,0Lx�-�����\U���`�<�|>�.ӊ8�,�=�q��<�}Q,��-Pq!5�]-�=Z�龗��u]�)�jx�:�%�Ĭv��g:�d����r�?Y��U��GG��ʙ}^����C7:�����y��R�����Ԯ�����~�)~�3�E��ћ Dx�W�Z�Y\}@��qN��!0�cn���q��o��|Շ<�A��G8��~��x^�p�����=ч�� ��2����^�@�vIppL���GH�}�ޟ�}��	#��m��$U漑S+��m?��l]7S�ayI�*í�U�MǦ��I[Hnk[X���٤h�*��̧��R��u�մZ�wB��y%�*��$��lPU靠�fĪ���uk$�7�f���a(�O�Woj�mFPw,�uD�O%���2�Kx���ε�ڷpV-i�E+�t6��KtS� Aw�ά5(�����o��siv��U�"�����uQ6\��Q<�f�a���K���(5Q�*mg7�Goo����0�`�`̮��#^�WS8UުL���]TU��Թ�۩��F�򱑌�B�Kquԉb[U�!۷ȦA�N�2Pڳ��c5g9��!7_F��Sg\UV��*W�V���s��]�]��V����ꑡ��kO/W6MY�`�7|3I"Y�ݰ#Q��2�Dﬢ�bT���n��ѓ�^Il��gNV!Z��E�`���n�n9�H�S0��C����-ڷ�M���<�Ռ]"�÷��ǁ��ӝ�ޏc��������^&͎�C�s.�H�Oqe0�J�W����w5A���UU't�̊^��vS�B�Hvi�)1]�1-5�V:�w,dJ#k�����5U���r�*S4�kD�+�\�s\�hmb�w��즱;`P����5N#t�lf���1z�<�;V��T�����3k�UU�U�Q�to�eˤ��B=��R��x���T�|�iR����E̫y�,&M�hU�Z��
��bݮ�\�K E�y���
���L����zi��B`�����8���ds<!b0rh̾�;V����Uf���;�i�������s��6�JE���6K)b�:�C�ڔ��e���-a��a�KfopOՎF��T"�g̷�ɧ���K��h�7t�c���CS/0(�jk��-ujs��eQ(͓.�����jB7����h����"-J����v�"�aLIV;�W��5#��.-Vt�B-9"�u6�E;5���)��J�0&1����X��|`����4r����F��B������.���`�-�F�w�lQ���5�(Sa��[�m���{Y�vL�%��bsig
��wS���mu��H�l�F��`�ֻ<�s�Ǚ��6k��D�q��Ϫ�N�:��r����$�Ãw��ssu��B؛WM(#�bnN�;-ޑ3[Y[���:]�v��������"p�kE�Ye�쉘o���Y��Ѧ��̝�ge����g�;���eu�w�ctgl.�ndF��ᠵRC��ڷ_nE�����ѹ�#�n�}㻈u+�̸ʙ�J�Wg��3B���ƷnY1��ê�[mk���n�Iݛ/�-:�� T����L�Jjo3���s	����{�.�J
���6��u35w{���wSI�)!�w�ؤH�^5ҾM͋�$h��E�o����׷�������Ƶ��_d���%$�" /rݙ��W4a"f���w��߻��������������FH@cHI(��* /]vB�rs�!	$�#��������Z־>>o���m�o���$ɰ븈A�r�5ꦼoƮ�'�v���1����QHh��dr�I�$Z"��b���,^y��
�D�D6�f�.iXX	E�W�ޗf����1�v#"R���Ef���� hb��\(QdLcJ`�}72R�Ϫ��ϥs�b��HH	!" "�(e(�HE6F/��#����w�Й����G�̪'���'Ε�[7q�l�1Bi�U1���J"�r�i�����^wCb�w߽���������j��ϻO{���b	�V�Hc����mci�� ��$@#�My��/���0�y K=��ǃ!�n��m�Q�!�G�:@���*�}�ٔ0׳/P�� �<VP�!cΤ�����v�!e`v�\ )�����!�x�#¢Yp$���a����@�01�/�yrͶ���*f�0� O�M�MJ�\˩�i�FT(��<��2�:��6'Ƙ�D��H���,:.��9E�J.G��%5�;e��Dd��������szO8�I����ߧL�
��2=-��м�o;	�c��/�d����0 	����f�h�8�� ���n,7��bY'HĲ�d��Gc�W��<��y�Av�e�\an�<:Ԯ�o�u
xo!�x��6�u���*�'�-�����*�F�[X���tl����{%e4��SU��aQ� �ql(�0������F�|`
NVy�-���F;�$�"걐�;��-�9���&�{��g����Ry���W�������^�;�����[Ŧ8pn����	m�#������{�| ��a��4��AP�ڮs.�~��w��5��'�0v�n�di�3����eF��M��uo��vl�T��k������)�������ף�i��R�6���#Y���a}V��z��n�L�K�'r�jGu�93w[�(Y�n�l�3��Ԏ��z��ƷyL��d��׶8��}�˾g��'��{`8���*5=��:L.�5�!�á�F�˿P�C�?Tb�f�ߛ���*5�f�@xFDSn�oֳ���^�sϗ���Q�0+���-�� �e�M�y�W���ߗ�H��	�Ӻ���omyc�$�8�y��b�h�i9�-Ϳl��?|>@�{e�u�>7�8z��m��f��'��\�M��,������OI.�U��:!���<�g�@���c�4ؿc�(Y��}��3��S�t.�$5�0@w�S�u�������4���zN�Z}^�"L~ ��|S_�_`��g(�.}�^����.l!��Z"	�J��Ҽ l�f���|�)pZ��E8�dS��C= 3{�da��r=[�L�u��p�I{f>s�'���/\�����Y(2F1�{ȶ\2���$ŏ�d����TD��8��]���H�i�����s6-*�ϭ~;  ^ӈe�ucLQ�9�M�^ʋ�4�ftxX�Ys�<��ǚ��^�F�ɤ\���P�l���0'X��	�UI��oKSo=C�d��9�~�R,��^����w2����eG�ى�7�n�/��F�6���f��3|;���ZDYi�w� �Ôe��_�6^�YSw:,��&c���p�b-���җV*�XSt�LReC��"�*[�p����A�4�@?x} G�>��(�8犉Vb;2��̵UT0��GE���!�E�he®���H0Lh,��"�c�����0_Inj�~�ɼ���%9HȤD�M���7�Ю��4��^!]��|���ȶoz��"��i�,v�;�_[�Y�C��T�c	�+�si�H5���i��?:C���C�u�/� ��א���n���4>00�C����o��z]��<�7n���Ee��uŗ����r�t�Aj�/>ޮ�[
#Ll+�dP��u{e�_@f�Z�����4.���t<'�o�DB��s
��'�	c�	=pIcH�CxJxw'�_�=0,7ed"*S�`�hK�3^q^Xm��z�	.�NH�C�y@o����kO���� .�p���HR G}��fL����҅�*���q\5�lg�	�l�Z�&����X���L�U�uo����RoE��k��G�s@w�p�{3?�PZ`>4&�Y>�;�����=�Z�8ô���s�DѽݽU4ix��`��^�W�?A�}�
��� �����D����f�yE�6.��C2�j#tv�,��pP̵�W�a��[ծ-���˼)fE7�C�y���¢���O�g^��iә�s��]��rb�Ņ%�G\-Qx���Em�nnv7'�(q���W��b�e�V޾�xx]A�*��al�%�����U]�з��<�/QHSך��ۥIӓ�j�Y�Sʋ���x�;]ǟr���u�>c�}�o<�qo��{�I�<�{��^q>���za���tM�1��f�\F�\h�7�i�U�]ܦj���xv\�R�����c>��/-^��Vׄ��y����t=C��|�J޶��"�1�h�/ Kwo
%��p!����mJ<��еt)?�%\�N�������y#svt����8��k~:)�|@�0G�4/�?}�*6�oLߴ�	��B��k�34hз��Zѕ�\υ���ƚx`.���<w�2�5�8�p6�Ss�+cŵ�H��˲����L�mX
b����wu('���7���f�;dbFǙ'�2c���/��Cr���Ɯ�����l�/�
�ٚ���%�t����K<�0b�ަU�u���
LB`���C&��a�+(�и��Pm^]"UY���Ȣ�3�M��S%���3�8�H9���M����'k䷔Gm/ G8��u6"[��`+�-P��yI�Wa�:_�r-?5��4J��L!�q�v��du<��:���?� ��� �:�9�Uzi<P�-��=�h]��ˁ@Z�����ޣ�����c*�%Co�V{b	Lf�-���]V����B�xV�����N�7Y]�g�@ݻǔ��&A��9��4���<����a��"�^���дm:Y�O���a���p;�����l�[a=���J�y��F��E^jJ�Y�Ӽ�������H)�+���~��>�ٚ�BD! k,:<���sآK'�y�L�{x��m�
R�4�쎝��9� <��Qｹa9 K.�a��o��EoB���������G��<�rG/�n��l���*�9���A�+{F=�� �K��4O>�@t�`p�� �����x){���~��!�:��}:>��/gHf���嗁�/@ ^�C�;��b`��>�?��p�cm�n�K�7�^�0�^\/EO��R@�;)�b#��%#
��:�\'Åoj�C��Ta�TƬ:�W����Ss\�igCD&Zx(֘{nOB^� ��!�
���)�u�Ð�w�����dO@��)�w��]E������ {��̵
�������<�����6ݴ�IS6a�bb���.��R�R�W��B?w�Z�}���g�=�@� 3â�n=jq�T'+��Ŗ�e��ͼܽ-��{���ok���+�Ŷ<�j�d�|*)8$�¼z3���/m��'���>��������D=<��b�M��m8��:��m�AƓ��3L�J�]�v>5gF0����$�6E�,n���F��7 �O3.��I;�h\��Ĺ�����Zs'5"0��Vf�YYtF�*��`/S��v��&��S�ٕ�Pg%2��]
���,��j��<�&�Ŏ�YR�9�z�z\"oF����r�H'��U�FV�2VH^�7���~��0L �ُ�`�SjG�M�f���N��ͅ��L�$�,ƹ�p��������Jr����X1z|5�UK6à�.9��Iw�F�|`
NVsȥ@-�Ø	��o�(\M�S���f��e�{�>��z6!)�� !�E�iס|�۱���LZ~K���[4g!�J��&��׏{x��n�~M�Ft��&OO��^06ճGy���[��f4���s��s������z�Kx���pd(�v�|`&
���}Ws�`��ۀ�"��m�-|�׀�ڣ��w�2��^.�qO�CܪE��H�A�t��ހ1Yu�i�ȉ�е6?r������ <���� Q��H�vp�p�ݴ<��Zhtk�Vߘ�$�A��U�G!����9C2���81gC�c���2{�yr��@13L	�ox�4��
r����/ȶ��K���v�άE��	�q'ҵ�LkU������ 7�44^�0�Z*
4F[mM>��ޙ��W����o?|�r���K�B h��=	:�1m����#љ}Bw�"+ZT#�br�`fZA"3Đj��*��#�͈��ЪN^�%9�eF]MN�6t�&����]��o�Q2+�y?[��0³���̭���2Y˟$��h�槪�n�T�Yk���ﯵ󬣙���L&�;1z	JXol�V�q���m�Z߼@>>> �G�uԾ|ж·.��q�J`��T�d��*\��K���h߼,9h85i�T�C�ߢ4aBޔ}f���,t	�E��,����O�*���˝�"��?w2�n2܌.(vAZ��J$gX���Q�;�-�>��S�h� `��9�l)�1�n�J����޶�
273L�!>1;�j�������lZ�0 �̟��?OVT����y�Q���x�� ��S��M"�ϡ��bަ��b2%�T�uE���5���뜯w�xyz����=(�������H�	8>��"�sk�&M���1)ͤhZ��욡u��lXj�����1A�a=>ɶ�c�[���p�8�!�e5 kpi���*�&�1t��ixZ�Cx	���)�5��f|8?E�ӽոFE��}���}�-x3�>x���]$��͗Zx��'���4�b�g�tҴ��4�O?w�<���Pp����w��wbՔ���u�fN�.!x���ȕC��
��y����I�rĮUx���� �>88�Ѕ�G�B��4x:���874��noc)yN`���x����*�
��2��ҍa'�xЊ�_}�aC����egٌ����U�X�
u��D�֕�󆈩��Ǝio�o2�o#QIs{���]�66�,QP�lɒ�=�Js-J�[9����Lf��-+��Mͻ����ͭ�Fҭ�I�\�m5#su�0��%o�
���y��}�:k`��,�x��|3[e0r����q��ԊT�.+�J׿%�c�o��naI��BYO����짇���ٳ��X�!�k��s���C�,��	�m�5᥍�k�L��s�?eMd'[w��l�<3H݃>�!���p,��'���C����k�ѓ��f0�&9� ���U� ��T�׿M�����Ot/m�xvG��,�E}�!�$>a�=�y�D(G�MUf��>����W���=��9�;�Nbv"<��D{���/�22�A�������r:�xy��?��z��zǰi��O/�vB/Ed�(k�7n���jzv��[��"���<٠L\���ѵ�6�;4[L�'�!׹�H�ɬ{��=Bn���JBǰvcj�-��Tuþa�0��5<e�R�O���x}�6��}�M+~�������4(>V@���ʖ��Se��	���~S�C�zZIh�W����ԥ�~k�u��ᦞ=o(���Z��6���E�n�q��I���5ZK/Ƅ<�_��0,�A_x=����+�6�xԠ���VTc��u��������y��r�����F�V���no$��<R���bƑpg'G��������4�xhVI�[C�e�
X� "�@7k].Ǔ�V�7C͉3���Z+/����+r6�����ý��K����.6�{�.��'6�:�u���^c���c�F���צ�/ K�
�^�oL�齎bY��)�JS�|��q�'�q|��T/�F��>�.Ӵ��5��K�.C+P_Iu�$�'��J.��)���6�� >�ų��G���{*�Y��,�d3�؄�S6��U}I�Oa�:^��-?2NX��L?2}i��=�#���;���r܆�o���Z}#Z}�zc���k��J�`]�e��#YL�nsQ���4���^���gs�5?ʒ�AW�� #�������`��),p'��:�tN�rw���gLu�
{�T�=T�e{b�>ϲ��С�D��wRL8�Jb޵=l�33,�,���3s�H��~�/�cюu��&��6�n��y�1K�[��kO�@�����65k�79A��6�/�~��HlPk9� Ь�r=1@�LݳJSe֐}p�s�����0b�h{�wV�S侲U�A�Gmc	�N���H���:P��4��.�gl�+Nz|�ǘ~@\K<"|�[�vL��M<�ݯFe�ނ��r�&!�l;�Քn�j����lÔ�t�U����;�r+z;g�ocݨz�ÇX�q�u�Tu*��0��B��`�Ζ�Ʊo" �JNJ���4�����(�p��u��Y�#�A��ݷU�Iun�CV�q]JP�m�/$���i�������2
���|�W��^ ����O@�xi�<�ň�Zd�"@y�Nnc��'���W*T���]E��A��[q�mb�'��;��Ԕ���Pz͜OX�Τ�N�,8��,:/".=2[gHZf�uwN6��c���^�0m؍kCzO��Q)����f��Љ?��G��F��Ah%7oOg�/�/�n@S�Z�c�q^&%��#4�ĥB�Gc�W=���{�DI,�-�'�/i��Y��^ �p�����`�^�B�>�Bd���s�JE2IJjgۀ�ڪ��L�ݱ�S�]ɗ��m_����?>��S����+���>���&�)?9��Q̱X��N�.��&�/ A`��ڹ�>G�=�l  ���Bm�Lpm�^�`�w#�K�֘]��E��}������ڀe!2��7G�D�apGօ|>{�ʢc�E�>U
�B5��܃���u�F��zh�A1��� �z	����޵��O��!��y�-���/Q�n_�9����&����ٞ&V��]<^o�eys����&�y	����	�ǽ�Ǳ������3l��U����
eZ�T5nS͗��F�����sܰ���:��^q�#�J�9C
k7�ÂŸ��3���t�K}Ɩ3o�Q]{@�j�.�rd��wswo�7��;�V���⑓��7r��T�2Rs�إW^:���Y� uUfnm̾��L��1�ͩ%i�b�]le�-�jޱx�C���Ux�N٤צ
iл/,[:�*Ne�nū�LaG�!D��:�[�ob���m�	�z_��e��B��{���6)�&'1Z�!�e����..�W��y��h#���.LKv�RuJ�޴Uj��f��|�W�T�)c`!��ɣ7�8�&V\��nzL��2֢�p)6 �l;"�h�7SIMkw��R+3�I���3��ȋ�`�,u�Mf6�"�,X�x������$Jn�v��Kx����Օ���KW�<ED��>B��3�J9��Y7wE�M��f�S*Ό8Ҡ�|ځm	��e�:�E�˙MֳX�C����઺<�d�v�6D7�A�GR�5���[E��#��J7��G����j�@��T2L�ݳ59wG�ƐP�Ϳe���� ����$e��ZgO��#k
*����BU���Q�3��CsJkr�A�V���
�ɇ�Gu�`�D*�+��1���aQ�cv�j�)�Nc
�S�[d8�X��)���p�#)���%u�+��A�ʕdձ��v6o��Y+Z2w	���h����Unc��R�P��ŕ�a���}y��(��&�0dn�#��K�t7�,_��մ�LԼF�xBiGB��e\
�[��uIY�Xթ�������IѦ���ifX-^�f�hl�Kʩ��NżD�٬�E��Z�-��8�Zy��`��u��iɂ�������v����ĺ�\r��쥬TU�ܽ����ͅU'F�sp˪��l%~W��*i���PMF�������M�6�!	�-�������VUNn���������of&�VZǓ�mW�wa���KW�G��YO3s*h���气�p�cd��o��:�v�ܧ���+`�4����Q!�Õ��`,V=���J���̙E0��i��n�+���Y���'�%wg6�GҴ�5ۻf��uQ�5ɭ<�t�d��=%�j�+4f���-2���Y	a{g'E�̛)��it�1��loy�kʸ��v����$+)��if��T�Ո%Uá�܉���ڥ�w�o���j�L��H3��bY.�)#��gmܕ�U���]N���n�n¸-�m��*��lvV��uN�դN��{����(��8CI�6�.l���5r��n���J�7���Vm��Y6`��]i����:ָI�V/"��a-4�3tӗ�d����2�\NM���S��W�~:���d�B!���O��bMI�J#$��c$H�������ֵ�kZ���6�IH��! #I������͌�$�!	"HG\kZֵ�}kZֵ�}},$$���a&fI�_�`wq,iC�9#	72:ֵ��k�Zֵ�k���.dd$a2�I$��r%�{�ߗK����j a���wtLh)$E%wta$ �q�#w]�Q��	F�+s�I����ú�BwrL�D�ޭ�y�F���S�3��I))<��)��d�JD���fc$f1 ��q&�0|r$�0R�����G����	@a=u���;�<vFe�&� J#�(0�^w&RL/}\�&��ICһ1D��˚葓�[��{��������d�Zl2�$���p��J6�A��l��3%oP��P�o%Bp����l�iœP*A���ګ�O#,�@��!C����ΊiS
������3tR�	�B�D��(4���q�� ���L�J�6�!�
$�A��f2�!�l7
H����E$2�i����A���	�8(G 뿗>|��֣k#���9�IīW����j��@8W�e���N�\~j>7Wdr��ZC��?8�;�����xtc~�/c��,R�&��ss�^ �`p�b&���%�>M�;����Xu�ƹ�7`dq��C���L��x�O̓ؿDggA�;hN8<B�0�]�A��^��`h�37s���]�xȝ=�rG��?_�L�|���A��x[�dL�Mi��ϛq#;pxT�(��K��w�ho�=Y�=��d-HA��������-?�6p~A�����E��E��NF.��s��8���ײ��E�.q@vBZ��A�#!��m��q>�rf�uU��ݠ�J���Y�C'c_�͏�ƸD/K�܃I�ϧ��,�0ŌY������c����*�/����_(�3��$͘^����h� h��ϯI�M�-z}���tȋF�+
���b���9\�]i���cE2Qp��:[�)@L$�"�p�+e6�>�b]��s�-�m[T�O����T�/��1Ry��w;4�F�[A���P�@������|��,y�/���W�u��IT۵S.�ZW*=�����+?l#P�NYSn�b��9x#f�9��-q�y.#י��KB�.�:Ci��U�>K "=ʸU�Y����}�I^��B��rV�^��VB�Xl�k'%J����%q����YG����R��}���}
�pD�T1�D#�V�HK�q̒���@L@W����DЯ?E�ӽ��	�d@�4�t�}�&A�'ZL�a6�����o_��
mTz��r���b�C�&Y��=�g�p�5��E	2q;��}�'ŰF���[�r�J*��8����U�
�v���dzO=1����PXׂ�P�Bxw���zp�1[N�\���~��c��@�rs�^���Լ㪓#�#���J�­t�)��a���G4�'���;ngL:�=���y`�y�~����Y�I�8��8Ϻ��y(:��4�e>O5��"�m�+��E��F��s>�p�3?��������様&�n%C�.�<��שׁEaNE
x�Ș���G]�$��{ .��`�V�&=��D��~ �[��0̟�a��%V�^�ff��E�V�Rn�[���0I�tE��tg/<��@����;�6��Q�2�i{{`��K.��L�7"��:A�r��!����B,d*1'n%g�k��}��Ĭ셋V�ྱ/`T��a
��빳@^A��3v9/���+��5�Ӧ�Ŏ�^���~�Md�Y�Q?$6v�����`�M����[J����ժ�ڼ�҄��r�צ�|.�D�Q7��po)�e'��ٝ�a���J]j5��Y��y�3	��>٦�a���<���]uϝ�;�Ʌ�o���Ӄ��ӂ�8�#�8�Q36�y�w����x��i���V��ߔ)�����v���!v��B�}�HX��j�PQ��'��\ d���'؝;o{2D��0/_�{r��X�  [@��3�~z풌�a{�%6x�Xby]S"�߷ ^�|vD��'��a�F�?CQ^q&��e��]Nz���pnM-b#u��~k���:�>,yz%ߴ)�j�U}�����B~��<�ԝs�u�ɰ<7A\��{��u�M�^�钝c�G@���0�0-�(�5�Ҕ���\4��#�q]F���Z#+q��WBϐ���3σ|�d�:�#�(�aa�]s<�妟��v9f��yw:������s�PJ?`�$�q��[o�B�}I�H�3��^��$�ܧx�u3-ۈj��P��se��?�y���~�p�]Q�XsWjT.�F��͘jB��=��}�<�뫹��B���;�o�c�?�&7�l@�����A}��9lU2%�Ya��;ө���V����װT�Oa\
�Fk�[���H`�c��<C�y�0�#��r[.�5�9L`�~�e��7��u̎`��K���	���G�(㙲�aM�s�v�ܔ�e�wW�2Z�j�m�
�2���r#n����F��Z�B��uu���+���hd�g1\js,nwlJ3�ii�q0w&.�2]%�����H���<���8���"|޺��������2����H�υ����q��v�y�3�H���:�f�*�S3դr:���r�����#rI~,���b�8��p����y"M�ݳ[��{����,���T�C��������c%�v�l��0v�r_A3�hq�vd-��ht;h�[�����k� b*hdK<x�斔2L=�N���k�MϘH	Z�X�����lmCWQ:���A��Z��
��&�-?4S�^<�#�ZHP +w��b ��M�e�݂�}��|�{*��l��̗Ah6�5$r��l�|jg�=�RV�B�~jל�k�A�p��VGf޳�a���z;�Ie�Ī��j%=���v�-�m홭��я6�>���kF>�౅!}�	��6�� �P�2N��de%�q���L��i͂"ro�����@^�"G<(��T&���E�\포��<�AB�g��&���bo&��	�u{�{�ehA
ȸu����a)fۃ)}`�׳��Gwzթv.��;�l�y�Tfp4�o=pZڔ�]�SY}7�R��cE�ڋqM�mNO,��q�(�*%��Y[�J�+�L�Q��>�TG�	 ,P�k)n�B�n4�����J�O�8�1����+���]3{lݾ�%c;���+�j1��1"���8�(�  dE��7˝m�/�bS*������j{;z�-�tM�8@��]V�5х�ϑ灱l!�D�ژ��"פJz�.�,e��m�+u����le��q6�����!iy^=4�}��CE��kH�#���yK�Ǣ|�D\ftY�Һn�!�_�6y�fBeIGs�O��!�=��C$-'�e#����ox�#1���2�9�qP��Mv;���]<^UG��݋wc>� �־�O-n��
�zo~��o+�"�ȇlu�6�e�����6��Yc߉��W�δ��<?�z�(�x=��u�n��	�P�`ω�@t�}P�p�ĽK�z��FN���	8ō.j}*��ȫY���)�K�&F��cC�Qx>a�7������n�:��r|ZoU�UB�87�g��ը󢠟��O�
��*���l'��F<���N�-i���ZnbV��Hi�f^l���Iv��O�z��� �5��^m���f|ǥ	��T=ɺܵ[��gs���au;�Un kX
��Q�A�QY(5y#!��m�8�t��N�S�4N����c���7�jҎN�t�<76R�N��h��������"�mnҷS�p��[U�`�#��T%ΈZ�V5�2_Cx��р�a��';H���K�$r�	�ׂ���}�k#��o]�]�p��n��}�,��s����{O����@q��3��_���|���tg?3�v�\�����:~O��;�P%�����z0q«f�n6��r�3y��c)L?%���cIv�L8o%�\/Ck��pe�`�L�Z4)n��Q-i������[�!���VW�K�E��O��2.3t��\��[�&%�s�#�.�#�ث�ٻ�%�W��I�>E��^�ƙ��o@�����8v!�R��?R�Lqlʙ�rX�Of�8�t6�$��1���n�P�:����,T0��vl��K�Ɂ�c�$�R���<+��/ݵ��y�僱U��p��ړ�d�2.���|`�(6��ʒS	Q�3_�)�O�
����m�3�`�u���Ժe>�OV������|����?��,��m��4�=����'f����A!!����u�y.�X��Վ��T�ֺy��*�͕�7�;e�Sm���[~Tl�?+I� �>�҅����5ތYV`J������s»)95��m��gI��J��H\��9�ߧ�0~�g#g�(F(��~t>d.�@��l���9c]����dEnݵ;��1R�*~��Vꬖ�)�ʪ#��#��k�E8��;����^�4��]-$�|{�DLO���ꙸ;���e�-�V�+��r��!�i�SͲ�ӐN�S�^��Vl3(Ї���}��8�l޲�:8���Q��qDq� 1�����|6���~N<p��Ĳ4�����'(�������b��k�3p.RL����7pM�e�e�����r�?,�n�a��),4\�k�}�3>�-�xtg/>�x�����e�ȷ�Xց��iu�6���]�,�V�Ɗސ��* ��5����D�������J`�e�y����w���|ă�/��B;{������-|�%r�dy���R�2f���_��^E���(�[����z������_�A]��O��ۡf��>�`� �9���U�?{��.���)j�҅ T�p�8�kP���~��g��ma9k�8�yOl�NT��X(�<H���l�ծ�!sZJAcV� )=�9B���{i����y�^�|�Kc�'<zw9�ȹ�lX���/`eyӗ��$�Y�Nl%%�j�U3]���׿s�:y��x[*�J��M����Z�EN�Yop㋫P�/�z{�Ru�cȽ��eA%I�?E󆺈OGz5�\�GU''iej-��֪����
}}%�}�]0��J.�s� ʖ������Y�V��t&����o2)a�YU�ݕ��Z]m�d�*r�Os�2����a�8�(uGs6)6�䵋��R�[z��l����H[�e<����gJY�޻r
�!�����&���f�Ǽ��"�8�(㊊/|�ͼ��xK$b�zo��mxw�A;0��!6��M�� ��'q=�zc�\bS�qId4��zqp:k9f�)����j��MA8��p�~h�@`鱦7�'��<T&i�hXptǢC�֦~˭�̅����eЮ*���>ǣ�Ʊ ���9/��p�,G02�/3�s�B��̻L*��X5k>�ixBP��L(�V��(%����U#+�,���6D���7���]j�j���Grlze�vb�EtS*�CG7�zu|���=��TC��v��
i"��4������3^a�az�d�#M��d�^�/����ؠ����8�zܾv��O��}ճ���i��,7�}.&%Nc�c%�$6p�`�#z	z�^����\ԕ�3���޴�ط���Վ���X�[�_�L�S��̾�
s�ۛU86�je��g�R[C�Cퟒ��[��X0j�<0|>a��9ʩ����oBf���73Y���U(eٝL���!�7~p��Gh={zq>53����Ëhz�VV;�X*���7;��Ц!9rS@��5�ۘU&��k�ޛ���� t����j�]P���/�?>vaJzz���BN}��[���r�|�Z��1�7Q3j���C�4�=x)�(wc�л�<�����e﮺;�y��}~�Dq q�QF��3�=��χ>I�㮺zPtv��rj�,b���0M���q;nٟ����D��Bn���MD��mD��3��3�O�3�i��}�fYD㌎elep�[�U���/օR���)��E�kP}��&%�{	�V%*��̘����v�j���'S���E�N��.)<'X*�l��+|b��eo~P�M;�	H�C��quۏf��/��ZѮ�\��H����~����҆k�H��
@�y�H�I<@��6��d���H/���B/��,ikȭ���q��<�����d1������v�|�a�3v��-9�h����\Cd'n��2�����2��!iy^=4�G_�Duz����\��z���𪭙&�9:�u�9Ɔa�޻j�欟PL���w*�b�?�z+(�0>��n�	��h�5��:�zK�Kv/L�NhL	m}�Ҭ���	���z�}�ZT-{%�P����T��4���Ӭ_�7LD�3��Ck���|��S�G6����?O0�g�wmy.���-����.&;���ﲗ������>��5��ʢ)����'~zi��&��u34E�
�S��@r�˜u��̲�Z)�bN��K���1Bؚ���7`�K�3}7R�uCi�f�MגyҘq"	�Ѻn܊󨡗�⣽q�m����n�U����V�H��e]��J
���7X���-]oS]�s��:�%�x��8�� c� �=w�}|�����y���	Qb�.[4�q<��"��q^����	��g��SC+t�a^z�h��unp>����V���s�"]�`�#�4�&wuw�G��^��ܝ�r���=�}^[ҋ�Pna؂�֞�<������4�Gzf9�C����vCM�Z�>E2/~��ϫ&)�Z��v9Y&���^H�i��e]�����\�ұM��أ|���@���=���\�2�}�}ka��P%�T�P�Z�4S��]��u�e��
�*P��d���\��^Kϖ�5���0��?F�Z�L.��խ��\b�A�o������RaMH��)z��{g�� (2.�v�qn+e6��sT�k��aMVot�n��T�:�Nl�A:��V��0�ȶ�]8ޏH{h]�I��P� Փu��a�3)ߚ(�޿rM���q�#L�L�p���$�	B���ѹ5A4(xuz�k�~z}��ژ��i�][�c5�N��ʞ.K�"���I�����1�M� �X��=��2u_vWں�<$�F24e�A���g�T��Y�U�f^[�5q�N�(oZNZ["�ލǈ�n`�ϕ��[U�TJR��V���|�-�I��n1��W�M�m�m���t�`��plwlU�-W��51�F�u��Z*�\�M�\UF�^�zK�A��:f���L���($p��R�op��wj��e�țv�f-l첄nm�K��{8�[U�ח=7{��Q�o7],{y�غٲ�V�����h)QV���_8|���zʘ���	�x����c�B�e�b����.�R�Un��T�!�#+����Q��9�&Pf�t��J�=5����`��L���8�:6�UH��:�R�Z�w�4�����{�ükkv�kR�:Z�PY}�3�Z�!e��	t�&�̺��%ˎ\�]��k;d���J���3�m���hIX7z��.����5����wx�+�2u�hL��b��O⦷^h��-�W6d]��W�;�D�YX��R.��cR�J���v��闅�7N㥼�d���M�yP/�]��*Vhh(v=#�&S5Z:�A��w�dv)������	���΢n��M��.J��V��O,^��݊���2V&�2�l�N�l�٧e�h�U��ʡj����3����H�B.�Dǲ�m���\�ZV)�us��y+R�E�8�d�%�7H`�դ�\A��i�b�WU�t��u���fY�nも��,1�^e��]^Q�~�����U��=�SYG�3(�1y{N��7J3j�,ܛȼ\e�O3K�ז9t�luG1�z9gb=CyH��+�x鄤E5-Q��$�|��"l��xP�#M�QP��o`��{#N�93Nt�͓�q�U��*��os2]Y�r#�{Z�U��L�OK�T����_J�
꫽|r*6Ȩ�5�yy�ʦ1��o۲3Ql�ҘV��ݠD��{:��Ӷ�f��������Xb����E��U��J�ʱ��z��2��ƻ�s�]�<�:%fޖ�b�Kj�W���F��f�Q�I�؅&��$�8F�knӤ�n�hT�8�ֈ�"�D*��@'L�Ò�yN��z{��řx�qE�>��vӭ$�0vg/Ԭ�5Y�Gr�s���B��a�Ks̍h�ŌSz��'z��h,Lnvi3p1A7��fE�j��"%k7&1�쇨Δ"X��&u3m���[�4.�\+Pp�u����ad)���Th����%�*��֧n�_RY6�q���F�֖i��{i��e���n[G^ՃsW4t���I҈�X�\6'Ql�r�����ޢ��t�9�6m��Jmr����U�Q�Vf�K!�53&wJ�A]��l�������v�Z]T�U�	 �|D=��d��ut�Rb�1��ۚ�W\���dȘ���Z����ֵ�k_���w���H�׿~^E��%&;�<u�u���$Bff;�H�)��n�5�kZ�ֵ�kZ���!	$! B��̢@�
f
H���l�B1��k_־��kZ����J}w~u�Q�g>/O�/��u����|닺�Q�,�ۤɘ��4�˟�)J����"K���Θ�)��(��q�5lI	��QK���4�<�(]ې2G��$� �IA ���μJ2)3"����X�6C�\��=�ܢ�:$CH�r�2E0����90���azn�C F�g��/�r�|H �"D�	WC��k��9�����)8Z�x���7*��ڷz�h�����cݚ5w@} �lܦb��.����x}�G_�q s��{����ZB�+"�y�2v������M�hd�Fvܦ��-�P��PX��Q^q)��X��!���ي��`���n�[yᠺ�5�C�v��I`}k��Os���>�ۅ^GLYq������5d_�H�V�������Xk܅����su�2���ښ��\`���qm<<9Z]9��Wᯌ�>V�G��x�1AO���!ݙ��p*����m�5���^�C�N����g3��o3ΈL7})š7A���C��dr�C ��FcC�>�i�¼�Jt]���3"N��<���Cy�ў���鸩�]Z�sl�}ٸ�� " 
f+� z��;��������78�C�Y=0���A����U&����.���.6�%�b�B2�X���v1����}�y+��c=}c�����~�0o���/�dv��O߳�~"@�p�q-��.�h�ۡm:����5�BM)�|��sQ����T�p�3gH���5�L�8��aAi�9�'�I{ipa�ɍ���㳌���8�vz8��bр�����j#ʇoT�j��o�
��u��S��/���]Z?P~9�Q��*ޠRm��T��sB+k"V�{n��ڼ�o^쳋�7Dedk0�鱉�v��~z�Ω^��e��G��(c� �8�" ��Òj�XvW�O6o@-���
Os�{�;��3��43~D��t
,]�x�7Gt����A�+��|�Ej�j}� �1;�L	���v#g1�k�:y��;G3�,{[�yz�.�;0#S�~�	>_@Bo�z}�2���K"��)�$�0���^�櫓�3]��F���\���u�p��s�xnk�*�.�wEL-�]ctS&��]u���ں�i��x����2�&D)������!6��M�}"M�N�Ga�����DIR���`m����p�_�R�eK���|C=�,����J���O������v�ԙ�^_c����M�)]Ɣ�x,z~���;�|��q�bU���t��|������q�|��J�ߵ7"���F �0�1����'�{ˉ�HY�@l[ݟHq�{"#�ف�.�q���쪚:[���@̭�Ԣ��Ѫ��n�Oo��W��]���@�ׅ��F���զQ���fX6�t^��Ի'�ܐ�Q�t��_\a�A���t�=�`�x�gD[�D��1��Z�N`k��a*���RկQ�z�F���i�u�T�^ɔ���Y�mᕔ��9�n�����Ł\1c��4䭋 �̘ٓ"���Q��x��CP�T�yeV�Wt�����;�gG=�3�vB	����Eq�P�ˆO�o��7��|�/W���Y��t�{iJ��ôY>������L	��{�*iN[ؗ�J��MY�0�����".`J�a�\x�95���켏��?���7.��=�4�q�0�xi���ݯ\�ꕽ6DF����]�Bp�a����r��i��O\�M�4�Y�?42���9�r�����>5T�[wk�]mŴ�L�W��J�`�ϩ��7'�S:��)�,8�ΉI�a�E�)��s�gX]��"�^����5!)��L�ŭ<'�Q��8�����x.�q��+7�,Ʌ�=����8��%�.b'�y�T�B�]*�w�ApK�K�:\gm�RT*��4��o2W��+��b�ze�{gO"���A� �_{�	��m�$Y���	�{s���.�$�i�iF�2�B(�5��Gd��d\9���Q���4�\Եy�^�H~����|�bTVk>I+: 6a-�d�5�_<�T�sj9�/o���lO�t �И�ڶ<��6��Q;�<��[���&|7��H��%蘴����i���m1�t	w[G��F�4���WU��X3�%�;NJ�}�v�+X���~7H�:�B8zS��cw�Gd�h�JOc�[�'mr�QKV��$�n\@V�pi�Æ�X'�5Q���1�1nU����"�W�lmH��¼Ê*f�<s6��sî��N����ӊ�8(� ��
�E�X�S��%�=xOD��ΡU��<�Vd&P���M�೻����T���3�4�\�- ��ob�<�ȇ,�	�:��ȍ���I�����¹񩁚{'%��N��u٭���	v�Ƚòt^����VdR���^n�e�`��Pp��'��fN:;��.��*��?�/ֽ2�E������^g`y�;4[�Et
��%�J:�6���ރ�ѓ��$VB,D�Ms�rŨ$7ڙOC������\c���}�Qc��]+��6H�A������]�4ŧ��;�:"��t[9��%�!�h��*��`���v7ǚ�33:�win/�v}FF�ޔ]��HA�r�v��֞���y6�f/��Q".6�m�U�5Q�ѨI�����8ʟg#�o-B�� �,��KK�5��`�o[)���x�Z%�L��GPv~u���a��P��za^���#c.��?'��v}(�J�,�DH�^��[�NW=�ȟ:&E�_e�ͩ���%Ĉx琞�4��ק���c�}q±��iGЊ���b��.�R]�Q�ڑ8�R��l���3I�4S�*
��TA�oڪC�m�=+�a�-D���؄��)�+ ��l��&�dZ7z���٠�IҌґ�e{��r{�^Y��ӫH{�Y��ۻ�^����D
�8�8�c�
60�d���v�E��(�5��TXS�[�b��S�<!�A�u鄝����ў�:��Q�u%�^p{�� ���9�Nm#AP�)8���a#r-�tc{=!�'I�,a��L�NX�����j0k΃W�l��t�L�1����%>�$M
}�Lj��;I�=��yt�嫫���iwWT���_j` ^�;ޗmܩ��\�Y�u��+K��=5�(RW%�;��p����w��,_'�XC�$~�X*8�y�
ն�!��֧�oݿA$ڞ{*��֐��4j��0��q�>;
�9m�D��B^K����GH�..�J�úWmvجK)�P5�|n�����T�~���H+� ��C�e���p3*�^E� ��v���QN�R��r^��Q�$.�֡�n�=���0F�3�����e��⭺�k��7f�!��;G/��ՓƇ[�Ǿ�k��i�;$>�:�=[@�:DC�������썊��3���ȼ�C6n,4���0A3"N��<��{�3�N��H���xU�'qNؾ��M�x���tf��V[;6/.��Y֩���t�m�7����S���T�tI����#y\!�G��r����\��Zb'���+�R����J"淉�Z��r6v�Z�w��U�Ě��F��n��YZ�c�������Lq�q�A7�>u���;���ϰS���y���!�ϼ���}�(A����|�p��wQfd���,!*]���E��#���e�^��:��ժv5�Q�{����z�\k�~�V�(7��W�&[�\e�j1p�6��T'H��>�	n�Cv��yX��MGB�;ך�:P�t9A�5j�*�S� �ٳ�㦿P�E<�A�������w��˪���5Ҽ8�2����K	��[,d&UhФ��࿶�/���8��0@���/�c~�X�}ma�K�ַpJ���#�O5y�	M\�S���LD"�]����^����ʈa�f,�N�mQP8ԡc�O�����ƺ/�ƽ>�I�1,��]ʂJ�
�w��ڇ�iW���G2�˅�˘OC]y�H��L>ː�>��Sy�{9˾�:(�a~F�CY��:�3�l��v���b��̋�r�6�>z-�!��!�Bm�0+�b�]�d9����K#8ǥ�n=H��=�C�4�L?5�Zl��?w��
����}���M$p�yR���!275]������3V�qfAyyAh��Y/3]5�����x��.�J������er���Sv/F$�$�MMI�S�X��I�a�SR2a�iD,M�A��Ø��j͜�N1V��m�w��N<���tO�y~�qq����rg/�H�8�i�nd�����-�2���(�YYF	���^펠�;���� �R����O�sQ{w��F�v :���=jD��<�t��~C�&�q,UL�e1�I�oZ��^��V?�d�����i<���3��Y�n��mp������0�]4�vl��ye�Ѫ�ϡ�������_}�N,sۀ"�w�>V����k����Tg��^D>��˘��F��0q�J蟪��f���\���F���ݾ���=�ț�,C�{� �{��DJ�/b_*	`�ma�1��C�0\����脤{�o~���]�|�Z���k�{)���0��t�=z^���f}P�"ՍQŶ����^C�KEe+�z�?y�b1=x���Hǖx��--$(o.zc�*2u *���#�֯�1�/#n-������x^�w�ČSlPH��f�'��>q?-��6��Zf)UDw]1�]�R"��D;� ��yq�Ízn���MXL�Ū�Jr�[=��5�38Ġ�yn\��>�U�;6����K������=^f֧� ��bY���,���n��e_�D�`���S��h��!��e�c���.n���,jL���^YaO�+0�R]U�1$J�Ê��'lq:K���w��k��]JL�Yk.:���ns�/�]�&/�5Z{��w�uw����K���ӳ�B�T�C_� 3��f�iGe!e����l��Sۼ	
z<�����O�dp�}+���	�}Oq踃UKw�V������S�����#�.s�� ��z��,�Cd�s�!^th]2^u�����|�0	���π��X�J��a�G���y�l[����'�5���(ݳ2�W[-��+���O"�>MCj9����2�̴���L ���4uz1�Y�֙TZl��I����C�.$C�"�&�4۲@�=p��2(zJ;��C��ù�ߜ��<�<I�Qm�=/�&�@�	$�t���Ug���8�����ғ�]^J��z�l�wПo-n�p��yI��o��"t�`�����?�ߟ��Y�+��m7F�ǙM�9�1
V�+�����^x~���Խ�h��+B������.��g�.xc0��q&w1p�S�0i�a�8�D�1�?[��WD�ƔU�:�1J~�b���� ��/��O	D����'�_k�����%��$�1b\��9���-����� �Z�X�ɮX��ؚ�]�n,ӾDWK�'ݮ%��M�qiF�aF�#QP��e��V��V7�m���k�z��!�Ͻ?WG{��ƥ�µ�~J�Z���C{�ƈ4��cfg*wN�t3WbO�JGMjE��ؔ뼣<�u������N	�8&8��x���:�����ψ�{�x��Mi��gٖ�FoI.�T�Q�=���yǌ�f�`睖 ����0�]�3!�@��� ��=�Ǧr����q��C��J����LA3�⩹U}n��\gO#���s��BO^��za^��z���i��U��B�=��֨�"uμ.�t$�!�\L�_d�]�F�_�s���.��Er������r�N�B�Wv繋����vN������]�-y��&ڋN�X��
j&����y��<!�A�t&v�,/��b���{�9�
�y��\���9�Nm.����I�(`ghc3��!����L7l�jk[i�
��Yn9�jS �/L��}�&� \&)7H��#�~��;ݼ0���6s��޼����i^>�N\�B�m�2��v�ʞNK�,���Ɛ�y�k�x	���X�لxr�Ӱfw�^��'�f��� �cȇ��:�t�6dI���U�Z��=5��I�3���t�����^��ꦬ;RC���(����6>;ɗ�}��a�}#z-�^�G�c���VJ�M�\��9sS��7w$c�{(�媺+b�w/*\�9���$q+Ӷ��˦�"�0�^�F��^E]{���yP]'��co>$���&�E�6��2wU�ZW�N��B�v6�V�ɋ����4���>����p1���nw�o��-��û����������k�=����}m������2��??4���֚���b�By �y8�zV�NK�)}`v��Ǎus+į~��}�:3j���!���d���z�\�����q�������hs
/�����؂F]���[r�Q�i�G �Dc�Չ�d�s"�K/�����2$w�&�qghI�v�^��U�C9t)�� � �������QY���v��+����z�4�O}��eSb�Owb�^`x>�?b���� �;�#�ޜ�͜�&�X�\���}��n��n������ɍ���20�U�"�5�q�髦.Z��s:8�sE�K��j�S���LC��5�M��Bݠ�|��k(*JN8|��`�0
��5�gB-�X�-��+����Ȟ�T*wx.B��C_*��K�Zɀ��-��u��Ű!8�J�x�7=7���w�f�8�f���KZ�ʟ �6�u�>�%��bS�JK��b6s S�c�,Xͯ����o/���B�s�͕d�M7�c8�S��7v/�잰[��'���˺��j'B�T�KN��&�UUeVm�\�>wY��bCg=���V�{+#EKDN����킶��V!9�ՙ��VOuZ{��N���t�eZkV���d�KyJ��3��v�hBR��}y/+���^$���lvUm��I�Eo\�Z��ډ�8Y�n��2��'Wu��	R�.�:�3�������+�VE���\�%�"n�p����;%�/),���:��֧#J���$�ݘ�v�\��TC������u+j�2��a�}}�N�msǖUt�.>���
�ۡ�4�V�t��>ݰY{�^�qOa٦*�霦��BEWv�\�YT�f�Z���%�P��V��`9|[�wT�x6��sL�U�y�ۜ]}V�_,"����<��o!�w��qQ�	��]fR�j�C�m���U������J�7A�U ^��1�^�gwl�微�x���B�F���پ؄;��({]���J�-'K��W=�l�$������i	P��:�Q�v;�v�3�Vf+*�e��o�z�z�;��y���=˓�2��f��Z]��un��N��d��x�z��ϋ�����gq����8XSW��"M���y=����벮����	U�(�ocC�>�|{(����F�J�i-����/T9lsC.��Se�׷�Fаo��m��o�5&q�a��u�Xw:xr��7��Ĭ�b�j:�-��R�K�-�&Ҍ0{�oR��geY�^���>o��ܨ�]�+�;ܛH��\�����u���1%�s/�/gr�.��Ĳ�U�*��v1EN�
J&���Αp`�6b�ĲIJ�0�P�����-e��yS���*���,xa�{��I=P,�Q�U�QԊ�[��	*�Zz�y�̜�]Yg�CH<�ss�SW^�E�>u�omJ���uQ�2%�No2u
Nm�ͭ�E�6�lI;�7fU�J�m�#���f�[��$�Ȣp��vūvxYW��,A#K����вC�ARȉ���<	��
�C�L���/t3�iN�Mb����'�l���l�V�V�{y������J�B��u�7��O9	�|��]U⎬F]p[W���{
ښ�Yp�HN���_�37C�6�L�u��,�Wݛ �+�p�G�T��9e⬇3u��5R[x�%f�T2%fҺm�qRE��I�f7�i��=8�M�"Sӻme�P��e�W.�aF'�xLI�ɽ�p��v�r+5�CV�t�z��q���8�[6��"�=x^t�&�v+�e1����M���q�D-�@�y�颲wQ�;4ʷ��qj�͋�54O���nk�#����ޅ\D��}7��7��8T(�'0��w���lal���v�)��l+V\�D�wv��nƐ	�o�ɘf0#�u�O}WD�/�%(I71�F!�Y)��{�}����ֿMkZֵ������$���*6�3dБ�6�F�d$X��Z׶��}}kZֵ�~~�(-Z�z�u����qD��E�dD�#�-k^�ֵ��kZ���@�4���B"b��ȍ����q��D�VB#b��$h���t�4�ȣEݮ��&	�ܹ^9�	&�{��RQ�(���꾜 ��0���!�B`fh�#Fz��+�D���wb�y݀��cb)+�r��BRF�Ʊ���-ɕ�iR�Wuzokڽw;�Q%|]��-r�F1�1�Ȩƈ�-�Tb�s�M.����^��z�bJ9<��F�I0[ �K2�� Ԁ�TR�R����ټ��B��y�i՛2���7�ʈ��>[Hf'�˻��Ve��Ѫ53��J�Rq.{K{0��+�"a-6�L�$�e"NH���A��� D�X,�D�L��p�$4RjzG�)(�	��_��^^>>@^���79قg��ڇ�i: �����Ucn8q�ˊ�P��d}��n$�D��{��~=�,�l�0��A3(��r�+��?7%$G]:��s�Y{�q}�����>�1Xjq	�/Sގ�/�)���y�E�y��H�i��k؍�,���/ޚ�U妇�r��k�w�
�pt�~h�B��s�;����d'x�8� 8@�/@����䠱]���Ĵ�����A�)�Q��z��jtIa�}WLO<��wf�#oJc�&���.�Te�Z�e�w=,��Z]�:�:�����~��ġn�!�8��&�V��vv%��g�f�iA/>�{
�����l[��]�Tžh�? ��K�K�C�t�!ٲ�k��Tj����,�����$᥸ow.ǀ�*�>.��L��=v��0��#�O���ӟ�z#��7 '&��a�zY�s�r�xe��=;Fv[sn��fd3�d8e�����M`Їhg�0��^E�/�^�ұ�A�S,Z�I�uy��0��Ly*nq��,v�Ԍ��^��5ؙV>}而[�I�v3JvlZ%=X˝[�{���fj��j6�/<rK�r�aY�vӫҺMlMR=Ί���Ѧ�uj�i:+7���Y��� �m� 5)��[���Y3�]r֛�ұ��"�J�mGXF���&��bv4�L�AM\N:�mҪx�����.�eO��?����#
8�|)E=��W��2��W��04VPC�qO슿(֜xlhg�����n4I�v�n�])�ZM���/?E��>�m���58*��Xn��z���>g�={zq>53�2�e����f����͚�`�B�װ?�4Xs�1q��t����b���'��3�3pӬ�~U�V5V�˥4���ב2��ւ�r,D����B�
nUkP��\Q1,��O�%�""X�л[u^��V�m@JT(�[�g��<�ۼH09qv&ޟ^��7ҹ�FmR�
�Z�z:[ySv/��d���Ϸ�"�����`cH�r�0�a���b�$�>�;׮���35y��%�Om*I���_<�T�sj���y��	��y@W���x{0j�!���/}p�r9�zZ��O�)�3����a>��8�"�H;������'�ᢞ������?j|���P���4,�L��(��E���ᐆ��t��ڶ{�z�n͎�P��O�;�ށ��9�7���D	m���k]<��s��*�%�Jq[��گl9J��W��爫15¦��:��H9jˊ�0�r�J�6ҝ�;¹���l�Gź;��2�ܗ|���2��s��Ê�-A�lD��t�(0�N3�N�Щ7�fª�hVO\N[��-E�B��W�q1�y�z����z�������
�v�8H3ഇ�o(?/�*�NK߻'��C��������و����/�qKt8��Q���P�����C��p`�D&->����%�>z4�G^!�v귄i��'��D��H�p����_���CJ*{C�8>B&u�G~�ݜ6}ǣ���'��̿]Ax�
l4U7��&$�x�f- �.�A�^�=��V.d�]�՞qvKj�gcȊ��3�2.5��0S�=5������zIv�T��2��Ԟ�����%8������e�P�>gm�%���'��zdmʹ�P�>n�!�%q���a�����rل�����#�o�qJ=���<�Ӽ_����o,��]U��P��<ڎP�ŭ@���{)��9�#�P%�Ռ���`1]�}���<�ϻ��&籐�Ɣ#65�xf�"]y�Pe�a5�W�F�(U�,)��������Y�>�����^ӗ�06K�P��3*j�:����B+e6���%ؼ')t��%�R�l�	܋hUӍ�s�W�+F@��ݱ�X��]­��3uNQ��MʛI
p�1�aG��/�uVP�L6/f\+��N\cX�ed�i�i�͕\��7F�����XG�Rj6(�X]����=�p��pn�F��U�Kq8M����B1hў^��������%�-F�M`�SsQq���ʟ[�g�W�xP&U[,�	���5���P��x��i�f�����:sSr�x`��F��Ba� ����]i�i�=�1>3Ⱥ^m��iw���R*��؂i��j��Օâ!����/N�ý4�c��sԼ��dOvJa;� ybJZx��׌q���s���E>?}�}�i7�CY����BsQ]5���9<�����A��YY��6���T�U�y�Sj�c�[ksK��A�p�;E'���MțC�ަ�F�ս��6����e'z?=%G�o�<E�Z��}.cv/��D�����.�,
fn���Oi�����r�PA&�U�h�|��ժ.;�K�w,:x��|�3�Y���frM<��6p�&��pL3Ry̆l��TXX&$��1��Lȝ��I����xmp���
���l����^!@�N�h��)�z*�L��1�D��0^P�S���=�V}3r��j��d�Fcּ[�p�a�2�.$E�>Q-X�ٻ� �X��&O����o	90�z�,����*=��K��7��Z�9*��zɿ����ߐ���;q�m#���Ё�&�n/߄�A2��]P��2�q���{�U��d%uZb4����B��]�0sO���:�j�Z���^u��`�m���>�������� �c��e�������Tu�n�R��k^�� }q���#ғؕr��ךn2�5t��μ�ň�t�L]�h7����\���͜>��n�����*
=уf81�Z�
���p��l*X��>� cA+���,�zr.h^���h���D�[#bv����[,��L�ѡI����f=��y��2�h��T�����`�@s�k�	���4�7�o�Ic�	�%%�^{�*����w��n��U��1�0f����"�DI�t�E�RE8$,��Ȃ\��Ks8�4�j"�M�'��;��mCb(�0���+�w0^��x�B`�p\��C��Kw9�O��ZٚHqo�n<0C�Je~׉�6�F;�=Æ�cf��C
{���C�O.�%�RV�g��h|-_k-(^_O;�)������?7 �L?2�;4����y�c=����o�0�v�#Kv
�2&P��.�`�֑�ʅ�(
2��P��PB�����i�Т'.D	> ����݇m:k`Nku�WÂ�7 ����T�@�9��;z<�����N��UR3G�OE�{gIt�¡�0��:Ob�K�%9���6�X��k�c���I����XF����0>.�ԫH��i H'�A�Κr��T/.V'޻���E:�7�r���*�X.7bh���ieoe�7�ޮꁋ��{jb�7.^�Z@��{��Dz=.���N���
����:�;�k��vl��]ʣU��K�1�Ȋ���"�^��J3wY�k7�^�;��9���N�!���	vO���n}���i���C�o5cyx���Hi�G�h�nn�����Cs��xQe�_!�)K��T��u�R�؃r�a~��B/�H�g�z��_��^��v�V�e���;�wt��4+��3n��Kꦲ�^���ϴf_P��X� ��9Awo6ޟN'��V��yg0��jZ;�=�Ҧ;[�Z�<��	��->�Ǡ������*f�Y�Jm)�	�[a��q<�k����;e�T�575w�;�d���}��B]����E(�צ���P%5�'}>��%D�ܳ�sl�;Rԣ<Z����ZgL��fa���Ɂ�.����^����Z�<���&�;Z�v�[�'���Pǟ�ı�dJ
;�����$\O�æ
��"5��1�MX�B�	��ן#X�ۘS��K.	*S綱=R'�.WG�Δ3u�X�"PW�DЕp�J����gF�3*K�Q,����cw~=ES�qp��x��eJ����[Z�����[���*�6Di��i�/����P�'׆��c�Z��.Ov�\�2ˆ�#����}�aE��<��č�е>�~#����O¸��m0���K�0�¾e�(p�J��b~�J�U�9�ϻ}Z_��N���a�|o��������&�t8t��5�]�r9���	�O�O�4�)^=4��e�,�%�f�G�y��{A�Xh.Z�:�D<2ׯOD�כqP�����L��~�xnʛ�ĩ�owF�r�p�üS�;C /1�v-��ߚ��Z��=E���y���6�"�m�b�'
�y�Z��~���۷�{2�S� �f|s�f�z`�}ЅF��z��#Y:���[��ڴ�n��|:�x��z�~�O㴽~���+B��y���Ƚ�h�e��VJ���|����)��=���0$87����nZ��^���,�:�.���R9xj	���@{�	�̐��;p�%ྒྷů��d_![ӎv'���>�_(�U�/%�g0B�׈q�q����E�'Y����f�P�(�Q]�5y#0�q9mBF�3�u>�|�PѮ�͹���y��s�c�|4=�+�ޟ�b[�.Y�_̗�1h�E=V�	�zk3�>j�׸ۺxv�4.��U�F
�1я�JT䕑��7Ո��u���t�e'��S�k&��7�u�Js��٧��j�o*b��a��ǯ��o�k*�mt�J!q�ab�����/n�Č��y��od����t���^)Hi��=���
!���G�E	����#���[��d�&�����y��k�!�/V�K$�m�A��.b������᢯�]M93���-�'ţ�j��y�����A� �ф�ё+�Qh�S����4}�(Bom��`S�]Ti����ݔ�)���� �������p�%9��R�������Jj~d��,s�۝�[���=��N/�� �}Q���^�ҩ2�0?���Bӥ�aMB�>~'��qqm�'z�}2vj�'��t����/�C*�.�;*I{�2.�p\1��<�w'���ó�̅V��QGny�������p��rsԹn��4�_RaR�����������ym�Ί�Ƽ�T0�'�q܌�2�_�-\;M���"����~�;���J֧�|y���<�]�U�]<�X�����sܩ&1
�ð��TԤd�Z��30���s,�J����=��^��G0�� kP��\?P�u�oL�g��Wf�#?���z�h�O�U�aɝ[�Y�յj'�n��^f:�W%�А��I�����tn����d��99�,J�¯v��pZ�qz��M�\�M;�����Ф�������˝#�0e���z�E��	�/3��x��������r���L���b�o'U\����`�
�o�m��KHH��~����[�vcsRX&�Ԩu��{�0'(��z��E_)�555[�э��-�=Z�3�M�W�� ~��{�,���m�RX`&�b��c�TƀܕA&s���;ւ�"۹�)��s˺Ɔ½�z�d)R���ᘉ>3w,�����ϗ���-�u] T.��>m����`dg@���.2.xi��Kf��O���%�^���4>T̆u�lQyj��^��r3��\m�j鋇�yg�f��` ��(5�vR�p|�A�N�uүa�)��=Bچ�!k��2�j�����Fy����s!��s�����B�ഭ3Z�V*H�^S�S�,'w���&BehȔ��ј��I�����^�Q�@��UR�<�� [HN%�}	�%W�m�[`}"K�w���6��<�^��C�=EPFɉ�؆ld1GN����3:zkw��t_!ť� ��Yq�W��и��}�-n�v1:��:E1)Ja�~��绘OZ���D �-�j��*ΐ��Φ�
s�@��*��530���꡸v/�K��j����Fl���A�4���w�d����t!����v1�Cx�Y�ȶGf1������lL]c:�c$�O�=nR���H�e��	����ƭ=l��fl���)��7��rw�g'Q����7����y���s��!<���Ȯt���]s<�妇P1�噃k�u趘�.�^&�L^�5�X������l������%R�p}�(��K�����PX�]4f9�8����@h�{�po'I���&闳8x>�}w뚙��E��t��sv�T.�T��j+��l%C9�#A����T�.�9W3J�<�zPk�������An�i����C��ݮ"�w�k�PK�=��ۺ��)�!�:�OVݑkߝ��{` ����w���' �\��,���}OeU9/s�,Vn��.�:����z�G=v�p�@h� �E�5��K�|܀͙�փ���ڵ�K��}:6=G�bF���~���e���� ��0:.YzS���fPg_��E5}+�}����`�#z	p	�=H߫�ы�S{dG��p�?��~{�jT��YV1n��0QP��V���#-�^i�q�`J�o�Iw/b��h��01�|]%���z�X�2n	#�!ŗW-�x�-�%,��0�Jm�d��eEW�3&�{ה%{l�F<��*鷹:�1�Zk^I���Uni�v0�S.�	l���ڸ2��jm�l�j�NN�Y��ˢj4�za��kZ*�٭��Ԭƞ+4�t�6K��a%q�vf���{��z�Ψ���'�:^�g�M̡D��d�T�x3~׬��J����Șj��3m�Z�U����z����\����*m���t���Af�W�sĲ�"�+��3�EĪ��ҝ�I���̧Yu��2�m��J�J�b�RWU�6�kcQ��[�(�F$�4(�2,FZ�͆�FA��D��Ҋ���3�VZ�j��L��H�8���b��N�ձ,�rӤ#Њ�X�}v���cw!�2�'dN+����α\��k��#r�Դ��|V>7H��syη����;	x��ns�e��F���3/�U'�C�
U��V�jP�R�f�Dm5q$T�@�Q�0�nXo)b%�ٕx���5R�^1e���tL���-b爽�.Vn�gy�+m�˃��P#�Ρ71]�;�Ն�9�b��a����>Qi�"�o#h�D�Xu`ԨP�
觛j�f���oD;V�9�q�q�*)¦nS
�T��
r[�������B�h�|��W� �jE|��s�N�2�"���T����n�u�o���7�B֓��v��]*�`Y��p;,$���b̸eE��
5A��c��)����1���>]���P�q�
R���k�C���g�9h�M�Ç%��ˋ	n���[�J)l�H?�yŲ�D��e�P�U��+K:�K���؍�Y�j�D���9�虫�{񯑍�IEq�ME	ہ�D�F&M���C��8�ደ�
ER�V�8Ry���hʥ^f�lv��jgv�u�ћY�=��X�q.xen.�ץǤed�3�\�u��̛�93�|������*��n�S��3L`�C�|I�;�f�M.�FFUê"�)�AIΣ��ڍ�7۝��`���w�3�b�7F�{ju�d�.��E�[����޼�O+r����4�՛��j�3xi��c<J� �7��&V�Oq�j��}�3��@a�u�A���Ǣ�F=tӬ����	�,k�:�E��ɦ).�jW7'l7n�*�]O�n;�����,&��G-���饑uU*3l�w:mJlif�7zbo6�n�J�qnue[��3䪨75�x21	��욎�����.�YE>�#���;�*I51v�Z�X�.��۸|�
�<e�j�t��n�չ)��^S�C�»ᆲ��J��䡩����f�@��mw�^#���[&ܠ�M3��9Cov�7�8�'biÛ8E��N!&�0~8V�;QJ���&�t��1P�2y���Ǹ�\OM�6ܠ��]n��umD���ͅ�nr�����&�%�nwNi(���m����-�w�yoo��q����X�`��[l�����[��M�SȎfAӈ� G� �O��#F��]�X*6�7�����|}kZ�ֵ�k_ZzHBBf�%�k�#cTY67��<5�k�Z־��kZ��{�X��W�����~��j@�9��!$	:ק����kZ�ֵ�}}`�����D���/׊�����^64�)7��
5�e���5E�+#�U�u�Ff�
�5ʙ�Q�(�4i�*5�]|�Ƃ1!Q��o�﫺C�L"/l�2j>�����6��lr�6�k�"K�!�W+��-��[Ƣ�A��h���h�1zk��m�π]1t3T�kj�ޔ��l�m�9`��/Ŝ*��WvR�*�ǼE�d���/�^m;ͫS��f�.0�����鉴s69�u����\Y��h(�[G�O�'�DǦ|��Bn��D��a,�S�X<'�1�Ř������U�0˸f�OE�+�?�^�De̎�X�j���_����]Uoso�*%�{�u)H�Q��cW��=5��.0'���a0KA<!�W-UO��q���������?1)��%c�IQkk|v�׸{Ώ@.-�����JaZ���]:�m���ݱ3(rS��^�w�F�|[И�h�%\Ø
'�v�#�,�3��:6Ԧ��ˮ4�?�r!6àۗ~�)��K��y�fE蘴����i��6s����]�}xeR��=s�U_C�]����|9	��U9õ��
�;%s�Y��C�fc{���n�l��WO�-H1ɤ�Y��6�_�@���߮An}R*�{"���q�(T�L�Mnʞ^~��p��wt�ϣƪFVŻ�c0i>��y�z�zz!�[+_M��A���E���Nd���tk{'��@��O嶽�h��Y�����w~�I�פ�[u�����ꗛ�g9NfJͥv�o
����6��+v�z�xY�S
u�˓�b���\��~��A��8?rN��auWD�O�l�w����BSݽ��ڽw���5�Ç���n2�y.�Zs��Q-��Hez}�������1�g�oYy
����	��P�픜��aii*�'�r�^ø�v|����Tr�B<�[��;!��3��V&d�v�k�n�g���vb��`����j+`���wWA4��fP����<2���dD�z��+j�b�cv}��"����@�2�1��}{h��J�G-�P����^m�V�f|�B-� �뛿:/��y��'qA.2�W����=�.sQ��������߄���^��w����������&�*
��z+��N)ʦ�'�T���|n� ���K���c���s~�΂�sb$�i��i�����槽C�ߢ!�՗^��M1p��}�q�tʗH��Qijg �N5��zkgŅ=-`�.��Ğ�7�����
�N�m�[Z�a1.����F��R��}�`�l���`�v�u�j-Ρ����􆶢�8�`�2ˎb}|d�)� �b��E'Y���"�Q1��/un��v���Ix����?�]q���?Jޤ��w�B�����O�����e�&�z��ds�R�r��ܱ
���v����f��6�K-����W����p#;x�з!T�J�F �n��ҥ��"n:�Cq;{WB�3��#wxҵ�B!������:���,�<�{0��UQ-�~������K����b/pjݪpv��w
a��Ǥi���Cm �	~1�q�����]7H�"{\�0Qٕ�o :��Zo���,)�S�W�O���Ə�vw��27���b����cc��ڹ�FȎ[��w��ړ�8��9!nBN+��aGa �
�]k���֟�N�Cch�%8�w%�5I�]5�GV��C�j�'��Q��<\W��c���ʎa+�u�sۿA��5�`��k��w����4O0E��?zC���wfcw�`�oR��Ǧ������7aəڔ�6F�U�'��
�I��l�? ���9�r�\d���{��BqQaDė��潭�W �]T���S�<���@CǄ[u�l��s˼ȇ��i�"���f%E����k�4�.ȟ U��>����Ϊ0rgJ���c�? ��Fv��7�.�߲�O{�b��0�{&=��i�����p��\:ѯ5�ӦΘ�}hg�X�a��htsh7���3x�sE�K�ݹר�X��0��z��U�㇡�8�}sr�<�y��=�JNǅӽcᗩyR�m�8陈�n˨:��u]�-�����N#N�3��k'Ho-����;շA����#�mf(}�x콨{:��s�g��3w�g�B�ü�Jn�\E:E�2���}G��}�gI�����E��9����-������  �I��	��T)<#r&=J�dg�<�k�]^=���|�8�^P��y2ҜK\��L�O��<�&��W�If�DħBm�Gm�ba��2���.a��#Bߢ��������-�"��qk�B;�J�@�f�{���벲[z��^�:��$�53?E󆺈O�\@.-�0Z��,U�vfr"�l��3�^���(+1n�^s��M�\��f\���0��Z]�i�L=���)[��fD�[y�0*j^���O�����'��K����҂ƗI���[���������ꋰ��ᗹ�� Bm0�Ϋ�^��Z�Q�w�Q��-F����;����V��33i����N���>o1�또	�,�vy�� -t��̝{~�!�G_isJ�����X�9x���c�=�[Ek����� ��}��\r���B1�e��|�����>�ȁߤ�^��	��zs�X��&?��lO���\Ø��Yf!�V�>9��S�����	���Z�Қ7gn[�{j��
�Hvκ�]�T���}�
��2#�^��Q�yn�t*���z��
���9Wfΰ��ݵ�/m�����Sye�TwF#�g*Z��v⎬LP��~|�fwg�/7�����?i�����JM���/�?�g����{�Xvz�9��p�Lƃ T�}�\#�t���Y5�=�R��[Z��r˫v�a���;O���H�QNCj~���EKǎ��ا�����3[�*�4�Oq�ᩏ��T'�b�ݽBPͮ �]�Q� b��^ŧS=rɲZzd,v���OӼ���2�Y�L�SST��.@��<tF�E��JY�Y��Sr�4+���^�q��*�)�:z9�skz|gbz��
!�A$��`�FK�"��f=";�&�Q�ޖ4�L�I+w���f�]D,�sv�ڈb�^7�S�cz��[U�>�fp��z^��"X\� yYzʠ�b��51�U��l�:��4�q�d�#��|�*���Xkܬ���& ��z|���c;���XM�aU[����!�q+�C�X��1)̈́�S*	G�jyg����.s�v�c%�@�C�U�PlMs&��F�8��	F�ۧ�~~��W40wR�];�){��R�$sxN����}ճ7�^�6�Q<~ݜCPck�G���$�1�����ٸ"�K���"�'�C)��R7�ڼ�%z���4�8�tj'o1�8��b�R�SwB��JXRX�yS-띭j.ZQ�Y�Z���w��ޛ}��^���Q>�-�z�j�dհ��]��V������B��ú�����A�Z6J��sc�Wh�v6gT�7�MƼ9�G�����ߟ�3t��]��WtK��y��Z`]��cS��z5N[���`�ߜ���\%�4�{�/���Ja�77C�Tjz/��ɤ O4+�c|~�m|{�H&����ٗ��u�MC�,��#��Jv��)8���QR�}5R2�-ݚ=���ma �<b��]Q����k���:�m���B2�#�����^K������A˅"P��Q�lܕQ讣�z��6=�~�9��`���#g�Rq��=4Q5�%�ܵ�?��o�%5V�#/�c��M�2�H���H�z�A�����ka�'M{cH��#�����1���z�
�ׂ{�<;�ע<;�N&��3�䕏��b�v��~t(T��jٯJ�*[+����zTo��O���Q��>�a[����?K̘b�S*�1�jj�s_*�T Ũ��RFCM��.qL��uz��>�a�|���*��A�G'ۂJ��Ks۩ȹ�[�K�X;4��ʒ�x�c� d�C�Ɔgg( ���N�S�SɫhUi�w%��ܷki��jO���f��v�WNꅚ�U�bwC
bP"��ޝ�N���:�e�}=�X�������}�	����*��=ܪݪ����R�f��W�X�N��[�'-��twsNmغ5P�.�<�I ��|||}�Oaʵ9&bt.7�n%5�»�K�.�������4�KV~2.�y�e�K�T�SR�R�<s'�em�t��>�&.��N�~2��>�
-�
e���N���+e6�{#\Jcf"S��F��
Jqu�P��'*b�*���te���l�z ���)BN+��C����ם�H��;�ԭ2ָ	���^�h>Ф�m��k��sքc�G�7=v{�5����������?�布>��0}�8�!`٫��Q��9�ֲ{�S$� n�Z|�����S������mA^a�m�M���f3,0������c��]l�	^��,r��rRX��,S$#蘘��A��յ����D�E�7��_�ֽ�Ĵ�*F�����RXk���B��pྲྀ�4�D4 E�#��/7kQ�Q�ʡ��x0z`���?K�e�bE*g�����iA/mbTs	]S��|�a���i��BYK���"O�Q�.�#�ġ���#�/�veu^p�3R�m��������{�S�L������Ѭ�/b�|�{��c��~a?X���]q����NMϫ�Cx3�9U�j�z����2,��S{8P����P0٬|$���(:�݊e�[tmN�(�f__+�©$_��͋Uh���koeZ�M����UC�!fwJ��Xò���M������<a�T^Z)�%8��#A��QT�ݸ״��
ߏe�+Gq%�I��}��s׎L���ǜS9|�<��h|/"[ɭ���E����3M��� �Uu!�xv&`��l�>������xw_�!�
ye�J�:��&àL�\v-�wx��9;U�ϵ�ޔ�R�����b5�����z��\��d4k�9n���s���ϲ�^�E��ó/�U�CC�q1`\�=ˈ�t-�jR{�A��t�㇬��q5�5oV�ο#+�,�~�f�1 Ϟ��C�ה��ɪr���)��2*�hRtc�2��dn[w�4��u(#���oV��)흣����k�	�>!��kc�ZbXL3>�:]M&�-�xD>�3*/�cc9&|)F�c׷=О�� ��!�ðN��.{�1"�?�j�.���_"�Լ�&t��ȹ��RJ��/e�]D[��`[�`����򚊴��Mmp��Pm; �nN�	��L,#R���*��C��;�0m{��<d��~��fDu�s+6�߫��H,.:�e6�I�}I�H�3�������ƗI���[���E�;���Vs��dcȌ)��2[��uqMΈeƫξ����`��*C��P�69K�����4�y�3Zs9G[�����ͱOgf����qV�:���)+q�2�z��R&�"n��{�e�Q4N�q��s���x7�����l��˜���p؄����-�0�kH��Iu`	�ÚGbT��F^�F��J�s��9����M��=S"����~e�X�<�S�b�����v��r���h0���(4��e���%��+��`e�l[���#�/�ݛ]3�6S�<�C�v"͵���7�]��A�T��Q�ǲc�O\��xt)1'hd�``����~Q�������� �����eUD�
��d�"#��:��ǟ���ï�{htx�Xh���7����nh�tm�쩫����qp�Pn|7 Q�v��V`L�wN�C��ɉ/����0����.hƃkP�nx��VNt��r�t8@��h1��闋<�սݯFe��W���4VPB�2]�c-�gbܕ�a�|Uޅ%�yǆv}�X$�Ӹ"�C�Z�A�Q���P���;��4�^�1�����2���^�f�,�p����f��c�9��BËk�E��О���xUע�gO�,^� �Z������.k^FHb֞�Fq���^=[ռ�Z�;!�BÄY�#�[�x��H���G??��g\ή�
�؅�����p�t��N[�v�L0К�b��-��3ff���nXڱ3l5]s�٥J�Ct�ês�G�mZ�&��'b���w,�n+���L�K���w���͋%��B2�!�c/ƣ��0͢m��������۷іQ$��z�A.xt��I� �hX%b��񹩮E;�D��9��&U��D���5���HB}}+���2Oa�Jr�	e�%I��P��;�b����'�Qk��@��mj��Ϝ;�_y_����I��Sւ{��q#�� ��0�,�_��RJy�1�c�3UDZ���6�\�9��]>G�E�A?�:�jc�l���T;g���zŧ�q���Fe+}�eqd.yW�(��w@� o����r��U�c�.۸���RbwzO,m�s��X���	�=$މ���0�x����`=�7�ˏ4�S�h9��n����{q��:z�]ᔜP���)�5����pms��cJ@��i��So��KK�ݶ�l�ɱ�]K�S���>֑��?\wl��������L� ��ltK��9�k6H�2�ٯ�.��K�}�������Ǧ�&@� �[���dI����b��e�O�L98wo� �,�|��?~�&��m9��3/�(m_ ����x��訌��Mk��*	u�T>�E��jՅn���n���iy�9�Q�0��ԂA
��dV3^I��su����u�r�afZ��e��Ė�^�d�n�P��3S%�j���!��X[uY�����)���	�9�!�ϕp��%�M��Z���34Dqm�)rne�e�2��~Uk�%��]����7��1d��&�a��n18����w8�m�na�\<���܂�t�j��zu`��,��]�yF�ݗ"%(N�0�7���dՂvn���T�
[��vX�b����z�[�sf>�����z\�5=���z�xL��ܷqXvT��K֏{��'-�{�m<�[T�o1�]�1�S���9�.�0b���*t��32�M�{Lʎp��t�U�Q=2�+ ��©2b�iz��E�3�4of��vx��:�"�V�9�h��΄�;˭�f�h�$K��b���t�ҡua ��e��o+us扨8�N-\�s���oC�&��	�=¡��̻����J�-EeDU,�6���&	.n�g$Y�tViN�	�j�w3����B�7���v�����E.�9shm;0M�O�	�sl���Wd��X�m��{�WK���\�/����[}�S�գT���'8v���-4(w;}7,2�N�5���w(�
-i�,V6t3�a.��MY�G�7Zyp2V��v�6Z{7B^��ot��M�ʓ�q'(閵��h�T�f�ǰ��kb��sp`�����ۦzP�׸t,Y6����1E�$�u5�딑��ݒ#�HH��;~��9�3Jʨ���t���+L�3��fT,=Ŋ�j΍x�D��u��2Š�Ē��S�&E��lU�Rҍ��w]�/,5KbRiT��-���͇��6�E1�퉁��Zc"�çS�����r��VR�+,:�t���4����0v	��|�3!�å�-��/�ڂ�A�-�M˔�oI4�fڛ<�!��=�csu<��^�webv�\��u_=\s��vX3(�qt�rl軞��2^��V̝U�T�k��z�s�1��t4�MX٫�oY5n�[|:�+�}��w:)��*Vx�0ż���"L���2�^G����qH�X�,i�,騰[�ij�O�K���zh�Q.�$⦂
p��ۆV7�͑�5�{��¥���Q�"ߵZ�C��}V0�!Z���x�u�`ʒ�7;%Vd�uO�n3+�w�gX��Ҭ��x�rV�n�	v{:�����Ug/5A�f-��m������H�5l+\n�K���B��z��j�uw�"���>�ˋ�����Z�3&[K�� �nd�
;��
7�g�ݼܖ�A[Zj��W�b�]��B61$ڽ&5w@��ق��&��Y�]�N�vwq[�f�oA���#�E�D��=����j+��[Ũ�p�$d2/qv� F�=��5�kZ��kZ��T�BE9� �1 ���l$:��־>5�k_Zֵ����� ��")� �9�$�0r2 d}}k�Zֵ�k_Zֵ�����H�IX�X�IV5�bƢ�cܪ5^��X���x��T7��U�6��_2ץW�DmF��l[%Q�
���g���滢���+Ũ����c�ݶ'��sj(�5�5_m�b�*5x��%�b*+|\�,�llmܽ�w�X=�P̏RL�	3��g�E@� �������	�E	a�������dQS5.�������l�32, �:T�Zz��k�yB�-'��s�]v�9[�;g�W>B�_�mP�@RjF��N5	�aaE"$�H!AA��M�D2Q!4!0/6a��)-0@���f(��D�M��H8KL��x������������t �}z��Vf���������2�OXlwߒ����T5Y]��C`��D�OP�֜���3/�F-�k��=��%��M٨�d��BU�b�o�>���;�lE�x��<!�c�����dz����}�z�&eH�K�-����dū�d�N�H�i��e]��C�=C��`E�Iܓz�[nX��u�����D�ܲ�!����j��Z��R�}3�2��X�F:@{��s[�lI�q���:�ƣ���i����!��6�����ь���_�pe�d�eBѡJzK
m=���e�'׋O�/�;+_3{d�:N��v�h~a�P�]UJO½�8@�����	�{1�ߒ4�a�2Q��n�5ګ�Z��'r"��tNc�$>}�e����2�����}I���&�F�r9p����MR*L?��w0�f��I]Ȑ>�G_������@]66EG�_S2�.��
a���[,����K)꓏d�2.���-/t��׏;� �c�pe��:Z4��^���R��9_>�a�&�ˤ¨vI疠r�����ʡ���L@�nC�ˇ;�O��T>��6l��(U���I�]�'x�וYx�UK�F�+)T­�O��r&�d�"�7m�vN��o.�޽��ݜ���y���2
^�����m<Yn�.�Q�ǣ��__kUū��Ͽ�[��T_p�r0�c�or�;��*�t��h�6- #�}G��}��&���t4j� [薔��H��㱞l��`f�ۏ_��:v[���C&e�o��8q����=5�fEøQ-�01��3�I�8��=+]'%鈕�^�;���WR�~��	9_i�ԭ-�=�ǀ���y���4���3����C��Mc������j����F��|dk/�e���z��^�`<�C���Q��5�'��t[@c�1�$��Z�5�]�^�3"|O�N4P��^}��t%�46v����2���<k2�ϸ�G�3��@�5�6U���j} ���B�gvr%�<^-�lmZ`ˎ:"�������_m4�O�i�S�#!'�z����Ƒy�Y�B%Y�e�׶������S���Nv�/}}�8
�	G�ϲk^��G�i����	˚�*H�F��x�v�P�Ǽٲn#�u�K?�7�s�J-�8*��,mEʕX��2��Q�#A�ܲ ��ۺ�ub��6�d�j��Z��윗��O�������
@׆U��mb����V3�.�X�V��1���6s77c���O�y�7��g4�p1�S��aG6_9Kv��P��V;t��>�u�܇��ǁ�u�m�8_:����_\Ap��M�P�����y��oNo���iM�(w���L��J�R�v�����L��n��<���Y3����<sAǮ�����્����1xEl�$��K�ܟZ�$vQ�x$-���3E��R�����+�F��V�"��T���}���A�"����^��]��$�eWI�A�7��ǯ�Mrh���]ԗ�_��+����L���5^�=�8� R���J�|GK���A= _q�����Wԝ�ϕ�ƾ=xK��u��w�m���½_�D�)�~_oXo��w�A��Dֈx�PҸ�kf'�ݫ�Y�jh�� ꫟e'��9���"���T����W��q�8�-҄���$��;��[�v�r�B1��i�q�M5��3��(f�xp77�.�2n��iH��������ݶ$ �����o������1å3U��%����}
�z/|����_Ox��A�iց�(�w�݊}�s�n�&�!9��c�dc�1&��Y�f�j�o�i���Ӣ��e���`q=p�[?/�~�Cџ����kI�3*Kv���8H�<6�^+��Z3[ӫ#�9��$e&����"U�ƍj�Q2���W�fN��c���[8g	�珏����vZ�?��mo�)��y�":2J���ò��f�M V!���{�/,�=�m�=�.��k�BK��9�������A�N�*&" cGQƼ�K,�>�l  1��+y��ݑky�M�z�jY�	�7}��|C;�A�
P�#֨�d��s"� ��o�6�>��e����Xo���Fq�Ґ	\!��r5[�d��Ry��D5��]Iœ�n�ps��%,�3�OKjF��� J^�����̞��v]Lͣb;�)�x�6�<y��p����Cu�
{
{�ݗ��;�H�	8�\u���1O�O5]��
x�{=�U��f�2�<l	c�6)�	�їܧ@���3<���?g/J]���j�[�B6~��/�	�T�c�f `z%�L����1'��H�IE%ݾ��Ѩw�cd!�������{����|���:�gUEG:�\���um�Ƃ5)�.b��ol��a��ʻl�2\�5s����B��A�����Td���׉�bKDn���%�{*7W�'�3�y�m8r�ɵ�[��f��zOeb"�o{Ee�n�5(X\[B��&'�x���������OL���N���	9Bjn������EH6ԩ�E_N8�)��W�?�_�כ�߾���ۦl҃U�6�>_�9�W1�[����~Ag}#����y���x���Z�Xw�
4J�p�h�*
��x�N}/��X^k	PzITw�hu���b\B��3w���f}���Fb�����V��2���d>��fThA)P��f���a/��Nc�x�I��w�Ԉ>��tW1P���wX�/X/�ҧ��#c�Nr�j|�O��yQ2�o	��ǅq"k�+���:m��C` <2��h���4^.�?X��}��r�R.�׋�;=�8�"�Ȉ���V�GKX<�r�g��37L��<���f�ڕFXcs���U��C���������e\��en3E�ڭ�S}:k(h��}T�Eǖ��IJ@��\���2��L4M�-G���$��xi��+�	
�Bqdz|���N���;�m�Fީ�c�����yIf��e�W�Ƭ���I%�PGO��R�,^9ֶ7B��L$o�sS��CW��D{����\��ng|�+i���M*b�uM�G۬��H0V�&�v�Е����Ў^�/p=]wSB�4lQ��^o0?���>IޕL�mm��'�S�S�o��́"�WpBW�¸���e�0����7a�H;�}��E_��Ԩ$L���Z��Fw���:]>�4c\ʲ��or��7�ޛ�p�!Y��m�4zW�mJB��z;@�d��\������G�������zK�lt��U]��ܢ��g:J�Ψjw�q�zS�%�/�,��>^�%��Y�=צs�˕Z�QJ�_�����b�tɆo!cx=%�ZG_�X�%��F��͙R��t���M(+�,�Un/��s�y�m����i\v����Ɩ`�G�)�c���+Ի5�͡������#�"r�\��ދ�^���`p�`Ŧ0����Ƴ̈h�������:��*�3ŎI.;�~3��!��Cx�7~>����b7��[c�DZx���gͳ��h��4�x�`S슍�u߸�z�~��q&�:���z���-��S"�f؜�(�`������mJ�Tps4�Y��y�Q-$jP�.&4�'��(k��C��tw;5)�Mv�C9����V8��b�R����:{l�t�z\�,UW�]��;��3���dZ;��bhW�(3��j��OJ�k�8gy�ž��D��̼����,'�Y;8�{k<GX	f6�����1�`�u0�L����a��*'��]�Ċ���J��nVk̽b�fTe�ٓ�r��v�%����3���ϓL[��)�{̪K���1'^�?v��v����M9����nɹ󒬈�)��j)���]����7A��x��%b3§����;�L�òR��M�5�M�����"+���% ]��&I%S���ө��_ZF���y��3X�J�~k�N���α���}��.�>F��^�V� D\	�tc}�o�h!��f��o�ȋ;ҵrD�緄Պ�-�v�uSs���sfT��p�`��Y OzKm���m����h�.Wl^����|x|�vD���ʇ�t =���>��*��b���@�����e�Bؚ�XE�KUm��Ȩ��	"v�2A	��Չ��.'JS���-�l� �vY�qO`{A �}�ؚ151�w9�'94�K˫�LC˼�YF��.���Z��� ��9�6��~k-frPS���i��+�"=�������o+s;�S�K�-�MM*鋯e'��1��������ƺ�������l������߬��u�DD=���Ġ�i��Y��Kt�ѧY�DlZ�;��m�Y�|�xS5�_�݀�E͈9us5�Z�%jyw֢8��=��W��վ�0Ѻ;��b�r�� �Ӓ*����F��m��N��I(�*1d7B�ߊT"�Mǻ�Q@o$�D��6��W�Vs۷��%����S��?���D Bx�R���ަ�p�B)�^�9��7^��)�AuQ�`������W,��,���0dgϙ"/�P��z+A�kŻ�2jϮTn�r�@���'�@	�f\K��*�V�"������q\J5��C��k#�e*H��X��]v}D��ϜnV���n��wk�19��9K��]-��{A*���Nr>9���e��;qr�]�	�����sr�-�!jWeDeS��P�Zc����T�-E�|Ι�O`�����i��lfj�����GUK����ѴWi7��m5k,v���m$��K�X�3u���W�)9m�%���{���עifм�V�]%/�����������ī0�B~K�Y�Vګ�ǎISQQ�f�dc�Ϯx�����?����������{�9��[��SF{Lʮ�;˒G��l��AVy�[1^�-�{i<�#:�og��tpe׷�;��4a�S��-����C�C���&��wj+[����N]�enB�IE �t���Av�ˍ�T y���p�.�2��1SfCd����0�H��T;��P��b�Ѩ�����_iX��x`ڴלa��ć
�pQ}��*_t�7j���9xܪ��½d)��Z���G!����f}tO���`�{��@�im7hkă�����ze�u�>W��1��^{��q�h.�3���*����3��ɣQdf��z�Y���� �$r�:$��:��F�xJ�E\_����zr��'�Z[��܎�� ���[j�-��a`�y
<���];m�T�����f����LV�sWs�;��'���s*e�މ�Qf���M���ݕ$x�6�*��g����Doc�G���Y��DAT�q8����a��aٕZٙ�X�t�-�y�KF�RW�zf^Ve��Y+�~�������������̬��x�۫�WӗV-q��	TA:�e)�n����
j211�,�ު�Ƅ��oT���".�jJϯ�uz�O����
k-��< �.�b�}�L���Ѽ����w�4s�������2"֍�<K``��1Y|�]�@ѫe\j�{��}�M����ק~��`T�	W�x<|c��3򔛦���� )��q�KI��ϳ>����n��9׶hc��%�*�;��3"S(������ꌖ��K_Q��a�nH�n�!"e��Z��e�o�"�i�<��q��i��t�؃�����^u�>�k�h��j]��|zzC�W8����ViΧ~��S�=0�
Q�Z�Wa�y�E"J��T5N6�]��IF5�ދ���O��w-n�z-�>�t�z:��˕-�	V�mvtp�Rh}6m�	��[}��)0C0�aǦ;ٕ/�@�:�=�	�������X�˨�{��V0_!V\����Z�����4n���d��%%��Oj��[�,�R�2�~B�x�����^���r�������xR��I�J�E�e�0\jT�SF�qY+Ctv��#�9�su�K�8�oE��U���gW��"[uE8�sil�esusE�r�,�q`�/ʧ�q�ݝ�v��n���*=|��.���n�VoXrK��,���U/jl��cz������z���:��J�c)[Ȓ�cfCףa���혣�����<{RjԶ�K��9�Ql�p���vV�a�s��df�g�����},c�����1�b�yv�&a�6��*�p^�GjgFl(�n$�[�oj��#f沕.}����L�5�ی(0�p;ɴp��/��»$*�<ģo5�nԭD��w_Z��wTI;Y�7����i�Ϭ�܉�Y���m��4,�;�ׁ�X�P�Yf��8��ɑ����ѵ-�-�Sɝ��ܙ�8��,9�/��ؕ�f�VJ��Y����o�8ΆY�9���!4J�;��5����0-���(�%b�SK��u��C;;^3vMZ���ѷ����5�S�z�J��\�,V̿K���83�}˛�#��;&m�������oe�÷3:)�T��2�,�2��U�9�r!#�eCm"��0�5+�o�����y�kFWW�С�*�������tl,�Yr$t�--�$�Tӫlr�(^��%�F��L8&R4~1[�ٖF��[��.�c���0�4���dm�ÔJ��ڬ��/ �%5�"έ-�@%]Mw7���9/��GI�YC�i�h���y��*�yݭ�=\��W�7�;�Wx�T��>`N�U��!�[�!���8��nm3K�Qqz�)t2ԉrg!kÚ,a)	�P�A�e8�d彺9}�S���ENU��'�x��n�6R�7�ҭ���7ob�)��!��#3S�TZ��I�:L`,�A].__lkN��su���n����P6��X�.,�S�ʷ�s�Fnªsw��{Z��2��1����i<�U�0�DT�ͩ�]$��25[�՚ZՐ�vl�b�v�8ߔ�.�p�gD�`=s5p��-�����f�S����z����IT��u�B�\�!������VRK7]^�O+;����(�%�s���p��jԮ�3�4���Ꜯ�P������o��9��%��{��a։"MGa:R���{�
ͼͼlb)�*�!���+�)�ź�K��r�^tE]%�<��m���m̓�;n��CT��U�{}�K���U�q��R.�F�bT�v��\Q�B�!�wk�9a��B�<�6K�+�3A�˽1J��xҭ��
���Ie��vfN9�~vD	$�0� pr-*-���%Y��kZ��ֵ�k�Z־����
�F{��ౣEW����!�##$�}}}|k_ֵ�}kZ���=�H�l"	"$��9��F>������kZֵ��k��{DA	 �S�-ch�|k��[Q�+ڷ����*��5�bب֊�5/K��ڒe�y�W�W*���-��j�6�p����F�r�6صs�o*4V���V׶�Uⱽ*�ǵr��_M	>��0P���x��M�Tp�W�_�L��i���g&u�}sw�u�7�6UpNqD���u�j�W,��}��Я/7����N.u��Z�ͬ��t�zW@[:e���G4�1G����7�cRFF|���+����w�S���5�.��n�8l1�����y�/�z3�̆���"v���юh�Ș�ŎH%��k�x��/2��}�Π���O��Ҩ�][�cٖ�3[ǧ�I<IxE@ȩ�1FLWE�I'�*u�#H�>'�L���z�>������� W�;�7�L�\�ۗ�j�H%ц��\��z�J��MC?>U@Ċ�5
�Uϼ��9��w&H�k��j}sO�DS��d<GHV��N�K'-o[���.����nޑ�A(m\!�v�B��Ux������p�s����A��Y����p��㝵�}�h�d�%�S���2��čy/~V>�qL9pzt��,�S�kK��q��&��I�(la[$�Wdvux�7��	����ӽ̗J��N���df:�&�.�vü���]��F�en�!s�y\&Lk��T�	���I���6Zm��� |c�������YٻT�֛�}+w �:�S뤩�(����D��	��&��C�MCQnQsT�&X������>��oZ,p�<9.�:��H���H�2�^�!gj����}�;b{_m�~��̈,�J	��,��]C&rn��-痒;�㖟��D�Uu�vTULNd��)�����(?xlr�Gtm�2��m�}�ޕԥ8Opo��|���>���8Cg�,7�;��u��Ns3D.��G��"�/��9�0�R�xP��C�-_Fg�j��D��o�)6�� ow�� W7�K�d���3�;�r�v!P.��J}4�}�1))M�C5�~c#7=1�� ��'���Z]ɍ$��@�;D��r!�M�;\�T�[Q���v�H��:�ЋJ}����ϛ�� ��j�M&��NY�l��N��z���RǗ7����j�~ITQ�S���s�j��^l-6X�=�ch��ټ�y,"|Qn��ڞ�{�2YJU�1S������ޏ^���+++�ll��mÇ�J�v`��Y�&��A�*m�M�TN�}��U�y�׻5&MLj62:��op�2��S�%xS�V�uQIC��H� �u�t�6S���4(�C��o�nC˩/e ~���}@��k/��wfs�qM��ڒ&�U0*�aK�5�4��cѴ;��V�jا�M�=��(��uW:xl��Bg�ֱ��v����B�⁐)A�%�{�_��&揢^�δ���8���=�T㹘E�D%���{[��I&䌧@/)�.�@�fQB.Lk���m=��N���>�!���9+/x_.�ڑ���9.&��/eMD@i2�u�a��u��6��u<q�J��Nj��h�?�ꗇ�p�B,7m'�>^x:�g���U�*B���b�U�<�(����5���FC�b�{)�Ȇ[X�ck���>͐�:dxyG�nޏr���|\��g�{~9f�Z����%�t�ǀ]���Z���<L��Erc�:�����󁓓�"��oUw%"��ISʯ(㊬����L ������7�RX�Lx.3�F�J�g���eq�3����Du�
�?)��"Nsl[��#��L(}�Ƴ=7��x�Pp`MY�;eq���Hv��V���7�V��.�]d�ꓑ�ߖΠ�øF���w��
iV��gB�=���in���W���޲b.�l騂�J�u�hB:��KYU,�*70��x����9]/.�w��=!���/8]��d
7o<�[Nɡe��)&<#*��UG9ڳ:.ϸ�7�V�~��`v�x������տ}������x�]�3���eQ�����Eo����Ė�tQ�u1������F�|���DDIí2n&��x�m>��{^9m��`@�`�^�m�����E܃��\�QW3�q���O��	T��#�
��)�ֵ3��!�o����Y~z7���֊Ѝ �S�k���jJ���o�^{�a���~d]�[$��eY�����Ź�bg��	���ϒ������Xu�q%�������;»�y�$t��ϩ��a��L�<(���F<�ذ[6���\�ʎ�'�h��9�U�7m��2E�Ig��$(�At�LNd�³�,V_^�q���s�G|�I�^k���s9���F��U�3:ث�nra��eU�����K4m���m��q�ɥi�P�K�|K��{_%�ۛꇡӑf���W1hc�p���S�޳F*�7sV�����,��&${�K�0WIM{��-]j�����mD��ux��!z"/�x�����7}�g8���PA�Pky�i�����#R�<<�U�v���ѽ��md�Q��k����������I~֭F{/ǧ�RU��J��UNr=�����]L�����r q���P�)�X��T;�˨���Q"&��흟2��W����͔���G��.��<��*�]"+݊�M*�>������Z�)���ƎF��W=кvz���G��y�}��Z����ۇ:�}�KF��������wi���4>���87�A�PcMZ�ٸ;�hnp:�8�x��p2����$�O�g����F!�h+y�Δf�G��iW�U�Ă'vJo�/�gS������:`�Ŭ.��6��O��\Ƒi��:�=�"�-�$���>v���9]���Q��i��H1Oa��q	X{�.�c+}z��N��1�n�R*<ϳ5d�^�w�g�Qn�[��AVd�
acڱ%�t6�u<r3*����t;�v�c�bnM�(|`�@�z]�FaWvrڒMl����^��}�[J]��h�$:S�e�{y��4�q���؅���Rj�F�jvt1�=�>>>>�����7��}��7�~z��\әe�!N("s򤩑E�WhU�Ձ�#.xi-VA�f��IP�eP�nN��K���Y�eGr�W]sO�Aa:��1!-l�6�>=�XII�IU>���eL�1�59a|rk4���u�	Er+x�t��0,!�'y'��]��1`u��f�w�����huS��!n����]����q�c�&��?���C�~m����U����k�d�݇�vm�n��17՞W������e�bK�[b���ڕß�5!˒���#0���������O��KA�3	������-}���..����Q�y�;�mt�mƐ������fk��<Wp����LA��WqY�J|Mժp:f�z����K�-�UW�&��F�	Ԅq�S�VKj��׷��<rv���C���R���q���s�gf�s��D�"B�C0�칷Fb���p��CN6�h(inX��7Z�,�Y����u�.��Ro�.���s�=��X�Ui��Y{v�Ի�&j�6�.1�f���ͻ���k(F�����շ׆Vg52�ms�'}������N���X����[+Y�4��Y��ҥ���Z�׋VBSaaw���Qp�{`:�0���GGt/i'��ǘc[r�}�L0�����N�bAQ��xV@}�%ۧ��w-�I*���)_\�;:�Y�kFokpR�SE:�j:����R""��l�VFmR�*�e�[���J4
�$r-���s#%��:BgݧUuʕqm\��Zt��{fdBǊ�3��W�s���M���ћjn�@�g�m�{˺��e5�'7�6H�U#0���B�\ j��M�U�s&�}P�#0�;����jW�xk�[4�hvD�v��@b����GVK�J£)A�|ˮ�~q+.*�V�ˉ4��ճ��N�}��^��=|�CrF����禚ʍ.v��a��p�ռg�7 �R6�`H9ҁ���Nj��nZ��{�1���2�:�9=�\4�|���r��g�	�	|k���-�4���*��1���g�x=0�xR~�fr]��y�A���0�1��K��h��"�R�)�2��OM˛9�B��E�W�5;�>聆T;�;*�)�Yn:vbM�j�+V�d��v���UV�
�N��n�&u-U�!�j�]�w8#zm���86Ͼ���� o�n��<���;��οo˶9W''ʙlC� xyMGzV����$1�n�����2"��jv���F]˱�g�[Z�jg���<�u�8�fh�ِ�k¨�������|ߪ���K�Ј���v�I�:�W�П0��B7�	�mхa�J{W��y��oz`y�t*#J�&���w��)��,4W�=ڶ�,�7���<�啱���F�la��|�q���,����L�@���C0�h�q�T�Kj/����|-�n��_q�1��'I!�A+��
F_λ!��|�환�u3)Աڛ<���U�Dn�<�$�۞x�{l���E�+�	��V��g[�7�5Q�"�v�Œ{�ǘ���$$D
��F��������?L����P�K]A�kF"�7��e����)�ٞ�>I�_+&����ɘHuҕj��A��N��_N�p����D,ґY2gu�,}l�Ǹٲ�Z������P٪���������f�eV���W�Q*7ّ�N8/�]�y]���N�#��u��\�Rf���χ{��������$��/���u�p.%�q1
�9f�)qkd�8!dd`��U}�T��~��#��s��Q�>�귉�@�ǔ��Y�\]=ܹ�Ph���<�Ƨ������M3Iǌ��ܷ]��-�W\�bu��y��Z'G���'x���m�"��Ғ�@B�2紝$w���♌��Kz��Y��_�3yk��nyE�֍K��ҹ����i����ѵS�/����m�]0�ck_Ⱦ��� �h%ݽэ�d��f���.��3����U���ƽ�`�^��;�+�%ٟU�,���x�E�Q�x�����î$�>�k�t�;�Vtơ:��u�|�lȊ������W�v���փ�T��C�!z�����Y֣a�N'�'m�z�:��r;�;M�A�_���?t��1n��r�\���mQ�f��3��74ܛ���ŭ���<�T��J�kVE��l\TC;j
̧-5&`j�4��2���v�0�1�5���^mM9���#L�uT����XՆX�-I��LMi��WJ�eC
o2j��k1 ~������r�W�sһ#;��^���p2�4	�H7���4�t���6]�Y�U��Q����i<�9�7ٖ�������~ڋȨ��Tm�a�n�8h���@���M`��Y����Ge����|IAU֬�U�;۵��%X$�B�q#dǐ�������k��E�h�ۦ�.��5V��t����R�.���Q.t�p�8��s���-��?fe^=���j�ܑ�h�tk�^T��2�7�~��2z�a���h�ѫ�\���(�B6�ϛ[�<��$�BUA��e��cE�Iߪ,�>铱��`WJɅ�S�"���JJ�ˉO^[&I%va���r&���i;G2�]9�����[\��wIT���҇���Pa��F���`��Uڧx.]mk	��S���jپ�5ɐ;oc$M�����fM�?�d�z��T�`���Ϊ'n��#sBj�.���9tXu��[P��]�!�o��U
[�U�5n>��-Y9d����1�g�Y\R�K�zL����BZ�ݫ&�eԥ-a����^���얳��:ɖbō�*�QZA�)lhq�]����]��7Z��+�ģ�k(�Y��t�GM�P�+�e�QꬨP=:�b�1����bܫ��q��0�/h��t��nɈ,Wu=�l-)+*�o�����0�I�.7Ti�'4�����J\8G��2�h9��ۗ�Q�{6�M�w��-�dVc��V,��o���IuQ��r�8x�ə�]K<�R�mK:�f�_�۽���2�ꐅ�:��4�����	ܭ�n�Kł�*s'%Z2Qܠ����ҭ���:�uo)���{h�⊵E��Mڮ'^��N��2����{_ͩ����O]�@�*������]�AB�s�Ԑji;�׻�9,}�Ash�"���[H�R��M����K���Wp� $u���@��R�;Y
���%��r�ayN30^�5!�O+0��J\��24�w�����ՒT��Gc��N�,�0+�u���e�ƌ!ެ�� �*�X��t���ń"�9FL	��D-��'�3EN��*�E�$�����5R�Gmu�ں4����;t,9v{2��U��pC&G!�^̛�F�F
����A[�Tכq2��e̑�E]�.��K[#�*њ�`t�q?�uXl7y��V������N� �0J�r�)~�X������aH��q���sf�Q���R��0	�����.�^[�&Ѵ&��g"�a1,�܄ʩY�3IK�J��2�L��Gm�ĉ�r�77�s9t�4˽(�c^��*�v�ƥ��%�d$jKvL;2嫈ӻ�;B�zn�-��ԥy����c$R�1J!�t��GJ�,�ΣnC��\G�����2>v�#�^�i8�TT�3�Bﰪ�ۗ�G^�|$�],���帤�����`�w����>�OAF�7�T��̓8!�dYۤ�\�튙�Qj˩[��X/;uчc����r��m]ofZy0C��[U�%�vv�ֺ��ԝ-�ӫ<��-)���*�R�/2]����_M���Y�b�0�{�^��4��p��r0r^j��-�wyY/���9x݂�X��t�ɘI��ٵ�n�پ�/J3��lգӓ[2V�u]�n����οNWc8���u<�3��xL̾�lb`�9Bs1��]��{�����۫�fnP���[o6!�)f�+��VIA��u蘧4j�%}�-�6�$����$��}{,1�q8��W	����n@ݓ�&�W�*���}ڝ䮠ey�m��n�K[*\������酆��~�5f��ו��U/[t�-Z�m�l��d��^��ہ�\�(�"JT�P�~y"=�(��d@dCE�d�$���^�^��ֵ�k_�Z���=�HH� ,�� <��!����#�����_ֵ�k�Z����'0]��ֺm�ݢŮmw��S~�׷׷�Ƶ�kZ�ֵ��{!�M�y7�sok�okomE^#X׵�E�lk��-�sb<[�^wj��6����*ܶ9��}yj�j����[�4�^�j��^�ͮ�Ksnlo�#�� �s�NI�vl2	#��Ŋ5�׶��U�ͷ�׍^�zk�Z/��O]ͷ�Ȋ��Zyvܫ��v��M��f���Hɹ16!�5�����oJ�z��^�8[�
K����I��H ��R.�a&$ ��@�"D��aH���!��"7
�3;n��޽�d�F�S;�!�KF�ͺ�I�;�*VBȢ��۝6�M��V�"1�V��Tu�k"��%S&��MЁd�5#��B�1�"rB�-F��YQ�
,���m�� !��aQ0�%AMB�8ZNH�M��P��O�{�|@>>�#_Dq5<�qê�Y�a���Q ��n=�ݻ�����u�B��]@��Ͻ�g��%�j��%��^�Q��z�T����:A�}���Cz�u*��}KZu��76˽f���1f �aX;�ԉ�૦.�R{�ݣ�x��f��фh�a�X��eH}Y!���OAڷw�SNc�4��G3��I���<!Ń��7�"��-���>$�c�<��;y�<Z��ڮ�䰉�A��=��f�ZS�
:�&7�]i��8������h�R��;�8����x�{�������,ω���>�3��F� �ňO"Ւ�o�pk�,�:!y��NM���F���S�NdA�S�~[�5ևH��֜�St�6[7��R����خ�ޚ�f�`�w3��EM���|P��Pd9.6Հ{u��+2bޗ�����\I/c���D���;(E��J����R����Z��\2�����)�sn�L��<�S�D��ha���A��K�Zt��w�M�%��$܋b���ݬX���Z�"�S��/e�b����}G�>/,ޭ��6��:��+�#�($6Ɖ�k�M���{}U,e�ꮹ���M[<�9���*����я�s<f��V-�o^7iU)*���N�H�t��zsWe00�:a���Qvݕ7���Ym�x��&I����j�fa��am�l;^"-�E+�؛�,�����]���I�R(N%��=������7����l�kf���Wp�/#��6 ߧkp�Z��%(�%�!v<f�eC�G�E@�z*qar�9��P*�;�!�r/�B�7_zs����b���U9dѻ�f��:�n�Z���q���#lQ�bR�C^5q�]�n����۽�J��c�1�r�v�ln���?��C�#Bȣr=��.&bET9Ѕ^/6ͷ�{=��OA�3����q�;:�:U&��:h�VL��q��q��:eZU�����]]o�s�K��̥�I�UQ��Z�X7���M}x8�'�`�T q[o���V#��K��+�����Y0��j��!	��y�h�k��Rh��Uۅb�R�O��>>>>�|Tn�v��bf"b"duiI��is��Ē�tQ�c���tٜF��mkYk�q����Z�{ fZy�FADA�x嶨t[���L�v�w{����}�=ɮ
�s9wI���	��s��7��*��K�w�1[���c��V�s�d��Q�+ӨN�#�-��=-��i-:��,�R�=R�� ��0�ʑQo��R2�Թ���ޤ��x�|��8��}��ك�6��G��=A�J����2|c�٧_�W�-��>/�R��9�T�h�u�z$\�)���n
�]t����B �1��(�H��PH�m���s�kvd�4y}0 4������@�a*��,-�zUz�e�y���CjR��:+c�.b�����'NfD��	d�ȟ.�J�5ȁ]���n�z�*[G[��������o|O�S���ӣ"6
Xf�B�s��F㲎��SJ���h^�x%f��ۃ���Y\���#F�<r�k!.�]2�Wv)|;xs��n�&iC��5���LW:�C��O
r��n��޾I�:�Q�� |||@��{|b�$���c�6�ey��$>��r�|[�dH�R~ɧ8�y�Jx��߻����֪w3`OÁU�"y�>n��!Uc��$��&��B/ù3�w7��g�y���,��0O�G
v��վ�[����x�1��U�{S�q�� �Z�-v�`c��	�uXozg�-Ea����s��y�Z�@J.�\e�k��	���=I�bJ���a�j(��vq�]��K�TH��Yj~�}b/�Ѱ3-�f��D�޺2�T�$���^�^_�L�������^��ގ�#!'�5u�3=-���N:�N�wk��"�U���ƭTH!3+�K��M@��7��V���yϼ�i�;v�,giJķݍC6��J.���>�>��[���֕ȇ���7��|���Ÿ��j��6�.�7>�oᗓ��M����X�5Cj
��U����tstɃ� ^ckNowgk��]�b���-y˰�p��T�.�+�&E��Q� ��Tu�[�jF�]��{Q��Y��E*Ҵ��vvt�;kU�Q��W$�H'dF�#S���F��Q����H�>  ��'�	�������|��G^MF�z\��9-9���v��[��M��)��}J�YNg=#���]-���I�%S���fe.1#����OyǙ����ą�Id�AQ\D
�⨙���#Al�ڛ=1��[�ҳK�RA܌���tQ�`�:�����<r�-��J������E�uf��yR��z̷6�jp�v�}���Ùn�S�o�Cz͒G>��'z�}�GRD��?J3����.�63���\˙y����gd�\+}���TJ14��A;���g�4����|" OU��!��3@ �ȈFb ����-(�f9S�����-���%ca�X[��E	z`8�e�t�}Y-��O�W�̩%�ݭ�z�4�i�[�f&v������	�"}q�.ߨ��Z;A���5<.��//&�2����ۉ*��'��>;9���f��*���0Nʋo�S(��v��W:�i�v�J�fC���!�8�#b�4�x��AؾP�fM�|څR�$Fe�Y�Xgd*9(I��>큇���k!І0�/�9�$���&VU��U4Jtګ�Z�nᬽ��*�w�e��c�3V5��\z�������������\�;�C�0�h��G^��d2W@~It9�O�Ni��Z��qV��۸�����C�h����FK8��1=��W=	pq�#Gu��`�CEw:}��p5���"��Kí f�\�L���v�4׳[��]}l*�z��QaZ3Sq���P=J�����=ź��]:�Z7z����sNdP �Ѕs�,T�,6W��b�=�7��cs;,�pD�/8ˊw��0�-�12f{j�U����d'5"R/xG��|�M�R��ۜ�q�B�uQ'��
�I%T�:��ʺ ��%�3I�癎���$�|3v�ïT��� ->��>���,bN�l8�Fyq�:ُm�V�5��W���iiLi~$]K�p8���>�&�+��Yϒ;eOq��,��7_�gOdWM���
������d��"�J�[o]��m&��b����]�wp��gI̦ ;�D3'm!;�� �+͕�t��H�ٔN�8oy��9b4f��m^�N�������G���d��8��s.���d5WH�ugm��zc�G�Z�`�^u��yU�r���7��ropR�V�Υ\� ��|@�r�f����oC�e>�`� 0����"#���loUnG����T}����.��]��J��'	^�I�p7��#y�F#+�ʟ>i�u���Lײ�cp�Y���7��j� N�m���x�m��p؀��U�{��(9nOc褁}_�w7�̓�+{/�b>�oz�xQ�������|K�?py�t���s����L�=���u�tP�(Ϻ���n�xW}i�U�\,�zSϞk�{3�/��3∃���[i���{n����	Tε�]�R{Ƈ7�y׳���wzOu�/(�U3���Cwu�ɞCU����x�\XJ z�/}�S^�Ib>5�z�GGT9 ���3yA9����D��,���ǣ�J&6�dV����B.J��Bn3R�$=ϓ�A�.yN�ٓ�Oi� z�k&���A�Y$K�pa]@"�Uvb��-�l��x)bU!\^�e�=@Mk^GN	J���3lf;{'��y^�b9�7�\��_���UB�=5]�P�W����u��Ige(v
̪�ӎ+F����/��YJ�6�
(ؑ�b��x�|@>#�u�N����^Y���8pb�Kg�rTS3�q��)�W��h��8�ŕ��ܲ�g����QZD
ށ�m�"�B�$L�������`ˊ7M�����ٛ�2��e����أ
kw��vD�з�mI�>�LxF��4ٸ���m5�/'�Ӓ������R�7�r3�����3
�?R�Co�H���:t���T4��l��-�����
ڷ[�j�h(�g�@� �S�H��u�J~�����K�Uq'c�?p*���@�4��nJ��_c������o/
�S��Zu^��J�t�|��}���`��5VB���q6�_y�k/9�$c���שw=#޹�f ��/�gՆ���X�1vj�l V�^
��c��4
˂��b��:	�>$�	����bM�3sleo��]]��v�'���5��2�}��'b�)�M��"4ؽ�6u��2�m��w�)!l�QXͫ�F5�%����y51�o�q��I��/��5+�wf�҉�@H�x�@F6�"]n
u��X�L��keN��ͺ�V��Wjγ�^Z��ov�<�ԍ�Leq�N7/Wu,�s�*����> ==�w`e����q�&�����5)�5���\B5�VEb�%J�����N|��Ss�5ď���)5=Y�H�:/�ml�B�M�v��s����?E��[��U07^	@{�]�6����:��a��ۺ800kk�"���%�d������ӝ�B`�`a�D�Gku�d�Y�{�㸅T��zMA���w"����fX�H��:���{g�<�J�1��"6���Ύ�y*��Tv��'�l��q;Wّ�~�U^>���X�V���)+c���8�6��#v��x�����]9����x8Em	ࢹ@�-u���;v�*6�m�	F�\�9R*��HY�=����S����d�5n�ӎ�����Tr;2_�H�N�F8�MJ��*(�Ua���0��K���9w�@3��+�s�/����qW/��}b5�;���z�ρ;��hl-�wƝ~���z�d;��n��j���ͦ�tU*eN���өZ��Қ���Ӻ)�'W+M�&,f]�򅼵JV=p�'V�]���R�~sB�rΜu��	�e�����i��US�l�*��7,��,���cwPE9�,(�x7������{�y�A��0�
2F+��[o�=����C��K�c*_g/+������t���/�8�d@ˏWJ���[q^��f�H=ZVF�Ռ�l�
����&!}�"���- ��=P*!�&�g7*�W��rN���9Xx��:������]'���"�{��u�kh��7+�B2H04�G`��/�C �������ڬv��-�쨥;[�w\�3wĽ�	�Z+)N�9�tO[�*g2��A�}."Vū�{Lm���Pdm�{JG�q)^*H�Nm��:i�z��9:̀��,+��给6��Sz�W�P3I��;� ���͞c1�q�d�fd��~�E�S����T��a�� �	���m,כ�w]�۽���^��'��M[?�Nf��љ��7��!��Jx}31O�א�r����ٱ��N�hu&�*O�;���I�]k]�f�p��֤մ�C�D��ݪyZ[O!DV1%��i¦��oqcl�/�L��n(��7
l:���H���[2�G�FP;�h�ٓ�邆��A���
A�	'D6����Q�:RG]:��
�b��	ҥ��Vh��w(��h4e�Ξ�/#�%�K/k�o��j���
�2��`�;N�&�@�s�
V;��f.���q���Y.��9�BVF�9[�-��;���{`�N�V<�v�	ސ����vP���K�n_ir��+F�c�yiU�dO)�UvԵ)�{+�
&k�h�3���+ݚn��^��A��ƪ]�����ޮף�U�}z�M���a��Y�ǔ�|G�z�"���uF!y�Q!i�YQժ�u�ۣn+EK�}��^���*�W9u͹�a66J�uj��h�I�WUx�.F�M�z)*���9��3U�s2s�G�y�Q:��A,��O-�ǠXv���� �4����Ɗ�J,x�����&�_���ŵ),�M`�$V�S�{ �0b��8,�cr�uj�mY�J;zS�n�M�ڔtռ��n�n��;N�[�KF�-;�����-Tb�����������F�v�% V�p�6��*�uorJ��a����GJ]x�_ms�Pm�U�>ɸ(kG:_U�6��O1�U��GC���3ga�U*�4q�Ǹ� o��Ww X8
���^�#��^gjh��Dk��1�]�,H��OL�x`�@��ӈ�؋l	Qq���:%y:�vt��k7�I���uu��-ѻ�P��k��d��r�LzƦx-¯��{�Cg���]̼M�n��{9�MtFe�}�����=�V�JǊ�l=ݼ�k	$��1���[e��`�z���m�
�J��[��rdأ�uRIX�9"N�Ð�+�[q!ݩ�%k8	�k3f�r�/,��δ�9�*��w=��0���(�%N�*��ɺ	Z�:y*���C�d�sTb���r޼�nJ�����m�e��2�P���C����bˋ;�0;�-N�4W_��G-����3��S$��kY]{J����K�۸Yci�9�.��+�NddPvnYI����r#�åV�]U᷹�.	/��D�3N��֗�Q���<�20t�^3;Z�Nmd��ݜ6.Vn]�m�$�r�Y2a�0W7����#�_em��:���eU\8k rP���ejo'
�X�>�G�S��ti���f�P���LZ7I+�QAR�BEh)�nA6�͢�����VM�t��^B`N�����(j`�h�{��Z8���b���@�#��7��2*�ko�m��{��nw�6j���ڌ�pH��P�Y�Y-��+%_00��-�^��m�&ޗ(I30r$��2#��-yz|{|kZֵ�~5���$0�N�`�	x��E����Ǧ僖�c_^�_�ֵ�kZ�־������˥�[ҫקX����� H�����/��mkZֵ�}k__G�q �#�Ǹ<�[���x��]*6�-s����Rܨ�J/����z��{k��r�w[sEo���x���zt�b*��\�y֯���RU5}��M��Q_Z��y�wYKBmDTW��^4k�Ҽo(ƹk�b(ץ�^6�y���wTm�Ij�\b1Y5&�L�,`4PX���x�F��J�2h�X�7�̕	�A$�H�	�#ď/�^�����v�P����dE6���-��V6��n)�RV4��U+�3{q3�7�ON�� �dj�_��� �����v�u�4f�4C3���1ƉT�$�����S�0�t��]f�%p�j�~���Xt��EYM�R���5^'�gCa�Z~�ܫ�Wv����1��^� ��1O�2��_r��k������Nʮ�f�' �kHm1�[m��5��#S��8ݵ6��qJ�zn��:��X��#L?'󀋳�5����<dDb�]ją	�|���p���/Ų+��RA��ݰd����g�#6<ހ�1��f��1��.h'+�u۬M�b-��U���|����ǝK>��2#ӈv�c�qx�j;�1Vl���.X7!��O�l��u�F{���_:�����w���r-��p��r��ؐ�l�s���wwEr�G�j��ե��70}�D`9Ɖ]/6����3/�w�(�=�Vi�Sʽ�aN�5�1}=�rf.|��`�f�AbȣF0��WJ��x5Z�X3D��ۉY�˜`�,���)d`�Ō4�r8�m���Uխ_EL51:�Ցfh�񟈝�z�B��A��!f̺i^��,�{s�FJ��U`���g�������E����l�j�s#Cz�D(�ݣB3וSwh��>�y�S��Ȼ���;�`��Y]:���z��s|�%V��Ե�Ԧq�5�|��*��9��YٚY��C�~�E*��Ɠ��p���,A���yStS����m�\q�d�z�^m ���=&�Tz�=�O���tY/4y7]Mn�k��]�TDq�\s�b$�/�EK�4�K��,_�B����/-�z{cm/h�Үa� V��	���Ғ&/.o�\f�n�f�WXӛ]��3�T}�;]Q�Cq��#d��O~�G����Qk�s�b��w�P�Gr�/\��z{|�]�����7O�uZ1{���Nx[��?@}:ص�e8om �]�.���P�C� 3R��Uw��
j�1�6��.R�]7G�Z�+x�k�E�½�6���g�`���l��|�nx��������	6�;[�
��^�{�7;v^Ǵ7oI3)�.Ҭ���8���n���e�މ����{&�yW��r" $I@c��z��+�Ũ�U��P^�6vn�u+yk��
Z��\á���]x�h��6��W����VJN��)�fh/�x���}��cn�iM^ ���'�Z5�pb8��ZGff���AU=�?K~��x�sy�竧�[������"[��/����7���0Sb{�ޥ�ǹ��E�v�i��by�sb�bZ�Ӯ�p�e��-y��Tύ}-�h�+	P
BAa�d�w�zfgy���Nsa� �h�γ��}�{�o�+#<�5~��~ӕd0H<��÷�y��P5��9���!6e�)�w��vW���b�	��e9v^v��q�'O+���yz�j�I�Q�����;bsK�=�| �k/瞁�'�*4���o-M�9��˰�ި��[}�kE�By��}1^RS���Uwk֌��nN�쇧�o�x��x=5c0��`��k�p�n|aY����nAO��N&Ҋ��>�Q�2ю��/�s���@W@����G������C���ĥ�qnF�k�����ہ<z�h�u�k�!9�-�����p����Vc�U��UN%�ͼ���@Ԅ���gf���fj��e�׊$��S�g��nE������՗J	T�5��wy1q�w�i�q��:0:'�<��> =�ލ_��#s:7�ĕA��\���<pR�ಹ+�)���N��,R��c�����=��2��;g��C�jtಊ�q�Q��Y�I;K�LAA��L���u��v�#�%�l�{��<�֨⪎M��u�C���\���Ǩ�Ƚ&��bio��}ؕ��>����U1��38�ݡm4���ث,#�[�ޖhqhD&�=��i���ʦ���S8�F˫���{\�� u'���C���ˏWJmY���D�IgF�7^��^-����t9e;/J4������	9
�$�v�5�~8��p��z�����ж�Fgw@���Ġ15*���(4/���B�I�r�����$}�<�A�J}�O�o����
9|3cl�ǳ�����-��r��yեB*�q��7�sQ%/eyƎ&(j�[���\�����w��ڋ��	(�~�����"�p�\:iםx�N�_c�O;Oc�-��9�y��N�((�A�-�>�nm�����OD����W�e��ϰ��0�Bű� �xv�SS��uD]<��JY.,��^sp�)�1���L��ߖ�uϷg�����j�5
:v�JY�:A6�G�j^ĺL���E{3m���}p��T�a������=����	���HvP��Y����H�w�G�v����mP=�w�9a�U�V���������UJ>yC�J���-��rA)F�Q�AI�j�j�R[@)��"���.�-P��e�X�{Yٛ��7#��*J�IU?\{��Nǌ����KR�8؅Ow]6�BJR�h�JC�۾�Fyup�lǥc�7=���b�B���Iˮ��8-G���lN�e��RL�)��H|��-�z��7�8�d%Z����`��[":�;[�I�>3�J�3X�:)���Va��o��Gv�Uj]s�����`z<��cyK��}��I�tD�VF���n��{���� �����t$w�V���ݬK��f눵T벨�b�����ۓM��b��g��lV�r���iڽ��4�����ˮGc݁�I�2�^^�ާ]7�TY��+/*���ɪ��?�Iv�ӗt9T�%6m=��[+j5ձ�D���''g�s�,wcqj�g��������|�]�tZ���W�Hh��>o:����
�_B�{�13R����#Hl�k+T����-�ݲhA�'���`*��Q�8t�Z֕%띁�8����V���o��� ����Î�oż�Ė<�e(ʘή���m>�e���/�={���~&>tN�����aF���Cs���g�\j�(ź�,(�(�.Ѩ��{�Zg�s�Y<!��m����@��s��@&�OYFF�u=0�`����Ne�0V�k)x�o����̞qϡ��7,���t�:�*RF�O\z�\��΂�8(�,ɯpkl֡O����,���`�׉Fh��<�@=�=4�&���|�	׷kw��=U�����!d
A�;�kͥ%~OR+�ϸ�fz7j`���{w���9�������������a��T��+�B=[^��J���mҗ=4EDx�1E4k��S�.yU�����U^~jSg$yS1�VV9�qл	�5�?uڽ�܄=�6�.�	@��/Y���[�Kj0N��	�-����4j�7�)5$�Z�<n��c��L�ڴ�h�uA�>7�.Cxz����%}���||�6�&:�n������Q�������v�D�ܘ�K���_��ԍަ`rà�`������ێC��-WmK����?^n��)[1�zw�A�8jB�[�]0���y���l��!��t��n����R4�q�aL*��=�F:���&��G7/�Hf2�Ū��*����vA���ϖ�xS��+��vg���$Z��j��ؗ�b�D%�Y�/�d:��'�����h!��QK�����P\9���=G�m�{��]�zn�/NP'����sY�/�"�7C���U�Xm�hd`E�+�@J.�͒7���j^i�M]�w-�lƋ�4�߰V���O�#E���%]<�:7FѺ:�dZ�XZ)�K��'�a�e��sd�Ez�� s���t#F{�s26�Y�E�r*��M|��k��h�O��{k�^����g۱q��s>É*g%em
�7c��l�7F��
t�V�+q���q�n�]LJ�#�j���gcY�Zh�ؿUu�����QN�#��-FFn�h"久y�CBK}+/mގ�ne
�o��G�Ct����Ӹ5)#�/{�����k��n7�5>��^U@��f	�O��i�ԋ��A��2A�Mp����M��jlv�u!ZR"���v4�Z2�Ѝ��>E��'f_f��6r�$��z��YynL+"�Ѥyħz�0�c��L���3^�B�m���17�y�����"+x���mū�]�սͽu؃+�t�$�?_�V5��P�����7�cMI�	�\�ln���%g�U�[szR��ʏoy�l5��*ש�2�Qt͕X����xOw;�p��Y��6k�@�;��Z���.OH�kc" s�wNP�So|�gu��婅kO�Lڷ�^ȽDQ(Ħ��uX��x�ż�}9U�#�S��/�Y��joC�ȅ�	��
o����������f��f2S��2Gm?���5�~�l�+ۋ�����ʉ�y�N3D�}o)�z��
"���\6��Y�\^�t�u��(�,�Y��Kn"�Q��%ń*k��U�I'��I>$� @ �FFtUUv�gM�qU	�F���*�~ͽ��DS�bp��}7`z���m<�V۰�d�J���V�W��G	���7�xc�٥�Z�=O��Jr�;5������`�r+˧ϸf�!�۾��"�������:�d7v�z�dSc�$�H�n����ׯ�z��"�̷CKq!N�������a�q�GO4v
2�?H"�L!1o����Tk�ղyy7[����$��ob�E�VR��*F	8[^w4��ngf��̰��v�&=S�]��y�<�P'D�Ƒ���n����.z�[*�����qA\�E�[2(+&jlԂ��3l�2�Ӓ|���Ű{����o�s�9���~AU�=YvU(@w����ɯ7H�9q�R�)I�;>���H�gL��2i�'7))�� �~g�g�P��m(�c>^�8�ү�f�7�'����
�Z��~��D����c-y�����/y��JW����:'	��;�xq����ˈG7Qw�(�[�ȪFA\&J��ɓNԪ��R�T,Zn�lI�ں�������+ե�u�N�:-[B���.B�k�OQ�7F�O���5�B]��39�n��d�w�W�Ù��;�U4�r�YX�"p<k.�3i�:%��=��:2�����6���)�e'��>*���ל���cs%m���'�FSjcw6�{�t:n���" �>�S;kc�>�@�}㹱oy��&�3��̒*Ocߤ�>ױ�B��s..���q�mۨ��/q�ngs@���t�wLP���ϲ����n F��(ҳf�54�4m���m�q}r{�!�/��֫�b��/��e��[������tmVq�̥p6�ڧ�`���	��;G"C�N�KB�Ɔ��M%�D)��sF���-�{�}}*��";q�O/�������A�ǡY��;��r�>���py��]˻}/�ݻ*�U{;�7�jSăj_�r���|��B�����m�f�v5\����Ti�.���\�`��ǲy��n�{��<���}��~_˕�9��
 �h*����������(���������+�{�sz��nd��KULY��,�SR��KZY2��1�[5-i�fՕ�f֖3m���f��5-i���,���ښ���ڦ�U���56��V����Z�����MKjjkRԭMM�5-���j�J��֦��56�Զ���-J��֦�Zj[SSZ���ԭMJ�ԫMMT�*�Rښ����MMZjkSRښ����MKT�6��Z���ԵMJ�Զ���56٩Z����6��m��Zj[SSV���R�jj�J٩t�v���6�R�jV�MY�����R����KY�VZ��R�jV�MY��56�Sk55f�m�=oC1��1�jj�MY�[5-f�Y�"�� �C� � �SR֪jU����SSZ �A�T �1P!5j��ڪj[UMJ�SDT �@�`��� �@��P�D ���SR֪jm�SR�T���MKj��V�jmj��j���T���MJ�SSV�jmj���T�@"! 7tCU ��m���56�ԵKmMKjjmSRژ��wZ榵5-i�Z��������jm��m�K*�T7u]�U"�@2[Lc+Yc6��3[Lc+Yc-��f�wm���X�m�L�Y�j�-L��,�lɓ+jd�VنF���s��p0�~��UV@UcPEc�|�����������E��������/���>������i�������ҕ�~�@ U�g�?x~�����  *���0�@b'�O�������h� ��o���G�=j@3�w���?c�A�y�������L$�q������B"�MimM�֦�ijZ��֥J�ږ��+SfڛMjSZ����Z���Kj-��j-R[j-j5��EIB@P�H� ��Z��mQmFڢڋTkRU�j�֥��M�i�JV����V�j�*���6�jk5i��M��KMj[5��-Sm5i��`	`� � H�D"b!`)Ο�!0?��Z~	�PE BA@dD	�?������	���� �?Q��}( 
�Ձ��|�#�����x'��!������>'�~� _����������* 
�a W���|?p}�y@T^>���P U�?�L���Y��C����p}����� p  *��C�C�}�}� ��'�3 ��w���������"����( 
�~A������ ����8?.��$O�}9��O�	���?��<�y�D���  *�H{{?$���{������ľ��E�#��磕g�a�-��������1AY&SY˭���Y�pP��3'� b:[|�E(J�( �BUH�(/�RJ ���P���*!J(" RHB��@�!P��" �URB��)�iB*��T�R��BR�QH*�UR�T��TJ>��"�U��@�H(""H"U"UBB�l%��IP�EDHT�E*R���$��UIm�T
�J�U U%"$T�R
�URE*��J��D%E �f$A)�*+� b}e���f�A2�۫j�nm�kl��k�8m��s��X*v���7]۫�&�j�]j�#[mT��������;u]*���wX�U�+5��ہ˚*��5J�(ITI�  	��(P�E��97�oB�
6�C���Q���Ƅ�(\x���v������i�SZبwr���.�kc�mJT��ӭ�J�'f��Mtv�#�����iSP%��T
�TW�  !�=Y�uNݴ9u�a�t]�r��ݕ���m��F���I�F[v�ݝ�v��Ͷ6[n�T��55�m��:T��T֬	V�[Ma��Z[vk���R�
�$�  nSV4��!CG�GjV��(u�֞�l���h��\;�b��l�[Z{:;`�+!�Te�YV�ь�T��T �*R
� jʐj�_v�-�Cm
�M5V��ڪ�C�*��	T��5JZ�m�i�m�j��[QT�-4��UI%P
��JD@� ΦP��vU*�U���+i�ӓZEM6�EU��2��Q�h�M�f#U��U�޷U�h��j�V�J��T��%D( �'� ���B�T�MV�
�( �F ݩ�� PQ�
 0�jtu� �)��� �VtCAp�(
O�TJ�T����  >����@���@.u\ : ���4 �t &u\�T죻@�[���Q� a�R����TQ� #p@צ�V �9wt�@;�( '5�� ;�` �6C  i���{{A��g@P�E��: �Ilb�)JU$E
G� �z  �`: t ��S:Pn� �n��� �{��t �;� �@� t�%�:  ���̕*��h�B)�IIR&�4h?UT2� "��	JT   E?j �T ` '����@ jyz��Ww��畞�=/�*`�.5�%��*]9����ş%԰�2����諭�������{mZ��涶�kk��mZ����mZ���6ڵ�����kkϿ����^�����������3f�ti�.�Uq�B�hͫ��.���NFv���(�$�>*�z�H�%��=50����7zE�^�4�S6ֆeY�Q�9u��EX[:�N1Su��Ê�����A����J��V�F�wi!�Ѓm�:��B����,�V^��*:ԫ�s��АT*<
KN5�"�b�;��>[>�"���w]ŒP�d�-���];����@Fm:�Cldۄ'���v!�LR�wjZ����A���uڐ�Q�V��C�2�j2-n]�	�#�Sqe�(YVғf͗��҂C��B��r������Tt�-y�Q��z��;�B�)�����N��yok"�c��!2񛹮 ��v7(�9���/݂���l�;o!�z~!x�X
��R4^i��A$h�ۅ:���4±��m"t1*z�����Ң��[��$8����@h�n�n�n���W�|��ڒ�CB�&�*i��bu�DN5i]%aM!�z��j}��^x1�YX��@�)��A�f6� n�&����*Z�P�x(=��6�-VF�0H�m�r�Ȫ�m���a3n������cK{Z�D
�͘�)`�E�nԼU��̺J��4O��������n	C1-����0C`)��F
t�ՇJ��כ�)���a�i�� {n^�e��@@�׺����B�)��]��L�y����G�䥁Zk/�7SAӷs����5�A��V��mmG�X@]ҭh�ת=d57oj�^n �:��w�-k%�j�����:�gi�YR,��(�.��4�#f�E�cVr�ڳ��̎�AL��x�4=l��{T�����+n�5���-������)�jjv�8Jx�Ok���L��d-V)[�N��#��fZ���%ٔ�]6�w �!�me�R�t㕢�`�i���Hm��0K��mc���Y42���^휕ȱ�Sn惊'@,�P�Rf�Jha�Vf���i��,����I��p=m��V%˳.iZ֙*�Ř7�*\Mc�@��D�ҝӘ�̎��H,�ܡw�Jf&���f��җ�=���p���]],r��=m�k�.۫��L;��7�;��*�唫i[t*z��ճp�fԬ�j+71OD'˭�#n���{��U��&u7Gv��+]d�	B�5��z�ٛVjnVb!째�тs�^��Q�9���3t��yJh͇dd �e7��U^&��B�Mj�\�@��Sz�����ƭ�[lӭ0�NA&�t��'rd�<� ]��dɱ4�T��0���
���uEQ[i:��j9q�c5�M�K2�FJ93b.KT�ق��2��{j^���c#B;�9Q;W��[�A����I��,��~�v�/�.Lr�W�'zص+"�V�@}uf�����t��~еݐ���V�5c&���
���%@�Mu��<Y����dX�Z��)L��j�j@�RJ[m6ZQ�fǧin�zf�{	:F7E�Tv�iJP����l�"`Yz-���
»M5M�����+F�n���#�l��yB��0��գb`I@�ej��@&f���EWŷ����,�v����@�a]��TB���+7���^$�PnR����iiF���X6�+!�����������7��I�0`�͋(L6邐vR3M�_`�adnEa��hIz����%�����v�yx-[QVŷ)�5��GvVi��wP���2�F��1�b��3�9��y��i
@�bl�����t�Ѣ�m�	d�@c8��ûbc��:��4Ium�e��.��n��Yn���S�vlQPl{wb2��j��J�/dS�̉�)��+�V���UfQ���E��V`�Qn�%=�(B�wECN�C�W��;����zJ�l]����%�l�m��MխZ�l̀U���ۈ�)�+{fb��+N�r[IV��5=���wK�[���ƺ���썑n��]<J�
@9��jP�\�mةy�5�H�,�)�	T�Md��t����l���h�N=Z������s5��ѵ�'>!��a�
މ�'N�9.͝�CTe.ͷJ�	RI������5O���ǣn;�-=�ŏ5���*�Ѡ�r�f8��&+��Ҭ2�oN�97k�h]ʽ�B�,Tu0�~Z�*4�Z���B�TUw&�$�G,��U@L(CH�	���8�7��/�0��W�e�����hDh�k��}!���|T�b��R��tS�����f&���C�� vVE�#{�!C-=����M��kM��)mX��Z�e�V�6,�A���ҷ	)���E��6�� a���r�n�#�]�J5*�5�� �e*q�w��wm���n.��uU�����v�!�[FV)8녤rfEI\��Ycap���ܔ�YX���������"RYQd��{O�Қ��V�kf�.�\�N��-W��A�sI$\�t�ߢ�0��F�@#i7���"�5���5�̽�.�R-�*���UyӪR��m�	��0���,ܫv�7�ONe�m�A�E�4��el���B�;��d2�VإQ	�v���Y�u�[j�`e�H��TB��GY���~��9Dŵ�Cx"�)Ge�4bXII�HK��(��qY0E.�1
oo\Ś ����{r����rRVd{{[� �3u�A%X�&�fޣޣ[xP"	�w�iT;�آ�H�%C��olm9�2�d4��)EB�Zk#6%m�-�6Ŭ(�D�t�\H��@��؇	��Dm��N�)��\�q�\Q|yjr�T�,XM+�cZΨF���a܂��V��%*5 6k�E�M���g#W>4��*�V��n.�C!�>�gr�2�2na�dE���$�:�����U�/���<��n�Pv��d�G�%�d�6��6�a��D�A�s\�	p�F��0����# �*^�,tY�����,�$�ӧA]�;�����b�l� (�<ݨ���M��e���W{)�2�ӘlV��ic�%f3!��P�N������3WJ����7N�j��ق����M�U(�V�.0~9kX�jHM7$�c�.�Xwy2Ɗ#��$��ssj]ਲ��V[n�nڠ
e��:�5A����
v�e��-KQ�30��]�B�ʅԛ�oo, *'`���zR"�X�,'[�mR"�����m�,ؖ̥
Ӕ.b9Gu'�$�����l8uV�b���U���ԅ�X,�F-���͵�|1JӪ��*���2Q�,๋&+��u�4�<ʊIa�LyB��U)�0�e+�E�hW.��L�u��˦�3R+9㖔ܽ6��Tlh�t¥E�-�"�emn:� F�����ޚUƀ�M��`�j���n*/*S�)n��2�XwN��b�|N7tDs+i�V�f�8�n��j��eӺ���5��v)��0wY�r�ȵ�ãB�Z�����kt5�nbf�(1u%b�V:���#sl�L�%R�e+��6�Հ��˼�O%j����%Q���[�%�j��Y�*4r���f��B�V؂��h�oj�l<��:�d�7�K���b�D�Ff�2�7+"�A��9��77\�S��L�e�c7Q�dn!O�%+/(Sm��63`����7&���J��4dMŔ��jy�3<B�h�|-cIf�3!Z�il[��u�F�v���E�<R֑�ZxP�Y����R�e����RQ�B��X(ӛ���mx�A��7O���(Wv.�,�V�#�,A,���V���7���'E���yV*EW�a�n"Q"��
���P��)�K��օN{� ����k�\���b��I��w���R�F���+~$�����ɧG[��֜���±�^^�g%�����0'��6QA�,���A�1�h�ӱv�I�,�E�PM�J�$�tq�jY��le�pvޫr������Q��Z�k���]����/&І'Lpp	��pkF���mne�51�Xq��*^�u����#�ț�Ty�^�l�wj���X�ڬ�
��ӌ[S>kf�\W���n�kM>���|��"Oqe�l%�`W4V�mF�nh*�e�^��%���	�WXȃ
��e#ND͠��SF\
!7�^=$RD��.�lP�H���2��.�W[�׮�i`�a�N��Sq����IE�x�@�?]k3^��p�l��T�ɺ��Xf�E&�J�N��[6�[GiR"!o\�a�C�@�Rm�H��F��3kd��&]��	*����p؋@T����Hĵ�e�&O�@"��M�X��S�����Й(�t��6�m*�0��[�Y7���hf�W�B�*J���sbv��	�Er��R4ְ��{�X�O/��f�1UBU�1�y7X5�V���q^CJ����%&�" �ܭI�������k%=����%�-M�v�w���!H)-��K�W��1��P47C!+�w�-&jwr��) ���-��u4h)$衆�'E*ae�C)YZDN������OLj(�&�%�YM�45�0�!TbM
�NL[��C�#2�YlMh��b;�H��.u���~4`�r����u�����\{�-�u���E	�*�i�^����(�3T|�"�*�ի�HS.��CH0�Z�T�K�Uy�\D�lj7LFiy��RU�bb��eTn�<#r����k���dR�]�b�E1,���j��F�Uc��s� ���kN�i �X3���& LvskjÌ�Y�W4(���'��z
�M�[.��5)<
4n����YMbE���*ޕ��[ʳd��QD
�I��Xnܡ��j�m)M�%�1����6��ao�&�'�Y)4��wke�T]�nSR��sn�։V��V�&m��g�t��E��F�5FX�х9�@�_��� �U�2Hۃj��U���&HѺ{j�Sf`��#H��tt�*��a֝����ܻ-�8&QBȤ4}V�d֭"���r@�%��n��*T̕��߅�aյ���a
� �[62�<�нN��vc6��e��BJr�����L��N�*���/Km�O]#ZN���U�"�i[�)@�E��ŊX*j���z��S��`���uj����e�Pԛ��bժ���S��+:��n�����)��S���iJ0Z�n�-$"�
: 	�sj��7�,�̆�Mՠ#��5�^S�k] nU�����m�*�t��T34�m���[�k.eDTXA�
�ʱ����%J�`�QD�m�";�筫֛��.$Å�3S��ј�*�ˢ���U �4漎U��Ru%���V����L7&�6�ٳ�KU��a�G^�Ql����MbǺ�}��P�6��8�[�g�Cx��4�VVC��q�NF��ECB-cŌ�����b5\��m]���"*<������H]9B��p[A���eg�Tv����"+d�fĝ����ɗ*��3DZ׉�r�����e�p��HP��`�Yktf����Ml�������w��YkPs^�E��%"�����L��[Hn]a7�/]n,m�t,"ޭt�c�	wI?��Z�V�>
�d�ݖ��������̸�Q�b��VM��M"6nVF@e�65�1��H@�X���%RVU�o2ɼA�5r�۫'cmސ�n`bkM^i{NИ��h�N�`��(�3	؜�z\���.�ǲւ wum�%L�c8��XY�	D-� ������s�Q+h1�)�]�W �E�)�њ��6=�5c�b����u�ǬȐ�֫�i�J�F�<�;w1C)g���8n`�:�t(�)fY���3;T�Թh��Ekd	����tP�wk̷�
�+[v�([�s6ɩ�����7[�y��5�t,�'sj&��E&�v�Q�m���rK�+E۷N�ׁXxL�.�ͦ���$��(�r���We��ҵM�İ�-�`X�rd�iǹd�B���^�i���L�n�����/(�e�[�E�36�藣V]ݕ�+3LU��� [-�`%�b8il�SnVՄ�*�[{'�v3V�
T*EHQ�4�[Y�^&,�tP/&IJ^%J���J/uJ�L-U�<&0��P���%f��E�2M��i� Cb���<�z�B�nj_	��6�ED�Z����M6^$�[���)D�b���c1��SS֮��WVkm70��+)�Zlk���M|�z�:�e�;GZa]��%�z :M@�@0㬳(�#���n��ym}��	�-E���$�w�Md���;��дDڄRlhQq8XMSv�=$M�˒�{Z�4��K��oy��)}6Ӭ�Z�n�sPu�m*EZjY����L�Q����,]Z�1ʌ��q�ʡl����W�F�,3��6p�s(Z°6��(m`��2�{������[�V��kU^4+
�Ma�A�z5�/�Y���Eܖ�L:����XnR���j�X�ILӆ��Y�Kʴn���)�JL�E2ok2�	ei㫶����hm��b�9k6n�ˀ�-�Q�i�[M]���(K���jm��S;�y�����i��z:�&��В (�7w��I}j=�yZH�',���"o&YsZZ�����a�X)Vm:�XG-�m1�������i�%6]m�xR�����le��*�Y��IDk�F��ڈ�16tl�dcC��XZ����<�.�+�*]KYUb��X2�T ��)'������Ve&�f
u����&��b�T� R�Y��6�t��)\V�?�}�.�U�L;}���D7l�	ٜ�;��7�+����s�b�gH�`;��M��g!hoWR�'uc��ݎbո+1�,7��O��5qw�1��W^�S���.�fY��:yGZY9�nŤ[�kT�M�i;�Z=��\v��u|��`�+Q���v��������)�~3�R�J�!�q�!�4�Z;���ݗ�e�O��ws�i��EB9
i�O+w��o1G��709:�:f�V�qF�=�xw��[MN!�Ŭ�7q�l�huօ�Ms�R�*�q��;�tM�u��H�%p��J��e�{\����4Ң�C�ftS=ky����J�6��v��n�8sc֐Z�D�)�b�A�Ad9�g�M������]�˦�y��X�T9��,�ȧ/eMU�Ŷ3����;ԅ9Ъ��$�>�{�vg`�uw��j��]p�ܩ[M֚���b35�ޮ1�d}Wە���.��$Ѿ�ݻ��)h�gX�P(u�pV�e�-�j�>��r�yZr��LJm\��/C���5��_h�A.�e��s36��m&C��:uC�Ę-���v��U�>_uܻ����a��\������ܱ̣5&z��!�>�k&�l���'#���63���'q9��']��.��od�joNuԹ�}j�v�yg9��������G��O�A������L#��NF����/��C�-W��	P�Z�s%��1��*�V�6Z��C׺;F�
뺁Q̺�f4ô�HՌ�k)\[x����ݝ��\�˰֣RD� x0��w���C�H�i]���q.��8���r�/@-�A���d��U
�v����8h��A=V�t.�eZ��aZ�A5����Hަ��a�k�f@����uZ�
ڹY���mc����pDp�ok��!�]<87���jZ������^�#9�N �p2n<)����Oc��C9y�ͣ2�Z=AM��������p���[�W�5��P��i�D����v:�hmne �L�G�I��*�9�%&W�@�����ٸ��1�錾���p��2��YXk��gf�Y�n�5�=�/jbjĊ�����Ӏr5>;�c�E������b��OF躒�o4.<5����S3ksG�+suwP���ކ��KZ#v����ܰ	v���o��2`�I�L����U�vz3ٛe�B��ZdJ��N���YkBi`�]�-�1�J���-.��[6��*�3h�ݾ��r�b�h�,��~Q&���׶�n������+5��Qaě��I��NģW�d�	w�1���W��x�������y�]j���gZN�w�$4۴�b��fU�R��|ʹy�6r��	e��_-{ڑ������ީO�׶���o�� 	��P:3,%��k���Ө
j��]�(.�1�p���y�R����j^)�tH��w;���<t�5�Z뮭c��#(�"�w��'V�ޣ�k�.��1����`*�'��A�ḁ���'�ք�F�Q_&�[mflm_@*P�c2�nz5Y'YK�h�R&n#�V�zw��V*ʜ�b�������Mu;�9�ãjQ�G�.�.�y�L��
X����˹@�״Xlrp�f���p���Ș>�6�ݨ�.y��{n+i�ױGn��9ӾV�s.\Wk�ᶟu���+��0	�Vv5��t'nX*��?�K�Vu�.���r�E��5������n�i��]�������
ǒ�u�(��kKZ�\�:�$��c����p:�Y�P`��sd	����uZG0>��ղ��O0�����7��&�Ghmp%%3�	"���:�	��pCC�nwusp.��s�!��x3���`=� w��3�"}���9J��Z5|�g�����%�4kA�:/5+����u3��:�кݾ�xXX9��cy6�͢�^��YBV.�SFn<kR��'�]����5�[Z�W�Y�*���N5������xo���nCQ�����'e�ջt5F��+��od-<j��Z7���g}�+��]@��*�.���RÚOs�ui�\�7�٪E���L3.�.7��o$�%�xYCI�F#�fܤ5;E�3�������C��r��i�aU�ik���6�,.�W��r=�&�+����vu�־�4�{�nCXsݩ���l�[��W��n�U��w�}b�V�JLXW7�r��� -�$*֩��7�U��(&+����Z�r�=5�%a[}\o]6T�h��p҈�7k;��/*b�p(cțn��\2���X\�Kb��_�)@5� �Ѝ�\��
��Ń��K� ��[�E���yW�f*4�ܸ3�e�`G+�y��1j�AN�!��s��֙ѵݏ�!l��������VTc�m��u��i�>:zRQ*5��
n��b�]$��LK-�	Ǽ��g���υ0+����  ��;U�05x_
H��}gv�4;԰����+�Rm.U��qj�U�Sr�t���m�W!�ʵ��G5�5�љ�R�;;�a�cDĄ��([���_a�:k�d�S����GI��7����:`
ĚK�?/.T����� 8�h�J�.��'WA���L�鮷����Y�+AB�un�pK�:��d}Lh�EL����p��w[I�U�4nX{;z�B�4���r���6�+4���X��͕3bn`��3!�,v��f��Е�d�[R�>��X {�+�*�w��B��T5��y�3vz��ʛL�n<][ghu����6�B|�}�owE�o���]JY`�!��w�S����d�pK!���[��cSF��=�Qj ��ƎG])�275��k ��mh��,p��)�F��nW%b��`��Z2��`6���Z�׻��������Nj4U�R[8����!	'.�����m8x�[����,N�ӗ/H�t��<��Vh��7JK���[w��x���[�k[��ޞ��=��<[���9�J�\���%Wt[���-x�,�	%nW ���K1�ӟj�7(S�Ǻ��1)�Y\��eTt0�4��^�i��L�\+����+���������B*nl�v��4IF�<j�T;%�z6�VD�D�wT�Lt�Q�b��2vաv���Vh'f��{�RNs���t X�S�I+�6���b�'N���nv{OW=��
М(j��y�2�]���e���wJ��b4��@\�uϫ0�ܛ^�	_^zz��47�:�}���L��X��7��d�S5��&vd`,��퍬�-R=������]K4�!*-`��5�g%�*�0=R�����M���WGZ�o��޳�\ӎ��ςm�w��&����UN;�T�9y�Klh�C8�>A�r�Tݯg�3՛�S�˂Uֳ�뮷j�vBu��6��� �;p���|��W���mD��\�.̺T������5dT�r�����eT�v�mr����.V
��7�yǩ+U�:6�9vit� ��l0�rG����\	n'��8�R�6
Õ����1����F��Pu��\�Cz�lB���@h�9�l�N�Z��5j�+�[�j����e�t�.QNDC�B0=ߣᷛK��� �l��9se̥��S�dO����Y��(e*C�%���Z*�].��"�\ޭ��f��UFo�λ�K&�X�L`mb�Q=3�����o_m�(����Q�+�l3e�Bn���N��)�b&���������JJ�U�X�=�(��Vic�;��;�*U�ĈPvI(��S�Ƶ�[�k��q��+P="��/����݊�I���/T]��;��,ᢦ�Oo��Łڧ!��d�x'`qe=������Z�%\����h7����.X]p�r�9�=	��ab��������K�c{�:�m@ �٥�W�����+pm��[�	J��0�n�!�v����Υ�l�9�4f��RV�	�0���)���3�+1�`�+����rM9f8gD��Lw�u.��Z�i_�]�w1C��i��,jIw
z�J�F����Z�2���{:��gu�[c����Z����mF��sor�N�:V�ZS�n�e[}�*.f꽬U�TT5�f	[��>X/+o8Q�t��T	RS�}w�U����U�$�2�"�#��iw���{wV��R��Y�O�k��*��`�SW���X�3\֕\;A����,�M�{S3b�Y��
�5n�g�q�NC)rkƣl������:���'@n� �k��v�̰��p�0��/�m�*�c�Yp���j�9e.{���i�S�n�����1�pu<��i�z���ru�,��5�,�>��S2�]���Ta�.��q���M������Ig}��0a��O5bu�S뾁��6I���S�;���"C�x� �����WZf��#���zTč�}�۬Cv�Q�Ha8�s�I���S��WZx��Oέ��C�ޞFq��������&�T��a��-����ʹ�����+�V;�V��E�pu�~2��D�s�3�ue%�6�.r�8ξ����]��B���/��mB=�(P�ٺ|9��5��z��
೥m���*S;8�v�k�m�[%�w6J���Tx�13+��u��DM�<k@e�fۗ:qO�����6�O�JfbĔ�7f�':����U�<�S"�PZ���]|Y��Z���6Qb��NƳ�M�5*�n�����q�����
Œ�V)��k���@^�X5�N��觪!���U)���m�at�5�í�X�طOL��f���.T���{�B:�<���/CM���5�v���
�:��mI���"뵗��Wv�um��c(r�y_�)�^aA��C�Z�%*�|���&�Yr�ߡ��o�\��.�G �I��������\a͒�B�tlR��<�T'1��=@��mGKWR=c\V�n�)mn�jҺ4��2���d�Df*�����y�Awq&�˹N�s�缟m������:����ʉ�����n؈�
�#���4/��a0l��ٽ7O�t�����u:np��7LM�{A�;K]_�_NDJ� �7�6�ZJ9�nZи�wn|����t��	�7-�~����Vf't�m���$�%j�M�\���p��7+�7��0%�L���IR��.<�>��5D����`��Ux�a��gjB��. \����I�&]�bI����swi�(�ԩ�a�m0��F[�@d�{J���}�{��u
y�!���k
Ǵ�e�dv�������G�ȹ��jPI��M<�{���f;�&�o)��`f7 �X�u\oj���u)x�o�D�P"Ļ�`Omu>�R�{���wq�+{!P��{K��1��E��>�Xe��ܗ��r��S2�r�c�� �pM�諦��4�qan�
�"�����ۮ�AQ-�p�V]�>`2Z��� ا$���Yr�kZyE�`!q9hsy5R �pt������q�̌�:�/>�7i��l8�3��.��YQl���u��ŕ��I�KOV�)�j.=0[H���ec�f�˪����\r���[[t�쭀���k�B����Ȗ�����	�N���Zς�+V-�+�s�P�H���m;��GUvR��;�YE�9#ќFt��v�NQm�s+�-��Tۆe��9ۼ��8�˘��%-��oC}NT�kJ��:���b��*�Bm�C5j���^g��tQ7m��ޒWU�1i���Ty����KU�"�gv���#O��{�g@�(թ�`�Y�sn�٩���]Ԫ�,�tM�L�v����u'�ff�P �Y�)����u-�(`����t̮ub���w|�__,,)z��-u�+%�2���v�(.�/�l�ݲ	=*P�9ZF�����\��� 1�f�i�g4o<�q����Nг_kK�җ;	�»+U&��	���L,����A�Ț�фyp�غDgV�][�����yw\��΁�BN��u��͝n�{b�������W9�c��Nm��:�{����ˀ^<�u�;'FeD��v��<M���3�Tr�����A[0^�r�G��el��3�W����Z�#��Dμ])��,]�j����.u
�WY�,����t����=y�G!�X��˻��v��VN��m�BH��xU&��8f�H���RZ�9���JvH(ο�=KU�;���E�>c4�d�pv�e���vd�I��+�MP[�,��]εH���F��Z0�`K��R�۴�f9�-TFCb�'�CG]���j^@�(vs[����S�e����׎��t�&��0��Wo7�Wne7�Y���o{m�S0��t)\�����a�n�x(���7\���|���[�:�K3�EA���y�0{�Z�"�_3��0An�a(�ܴU�WD�<5���F��GX!���g)zd��ʬzϯs&zH��c�=�p�:m�o0.�<Nc®�k�_՚
W-��Ͷ�M���.+�.�p3#�Ա\cC-��)��O�*ګ��K��Շ]�+�]V�B��m㬜ij*8���V��w!�[�r��e�,]'F�Ӱ_��Zʕ��-� �����;p��jZ��΢���گ���}tS��שl�N�Z��M'2DF*�j����k2,ⳁ����C:�]�p I	�F'��J�	�:M�H�|wf4��4�\��w����j�b�汲qnW;#$=lJV��g7��R$��u�%oJ��r�n"�����K��$#����a�A��C���M4������wq��Wž��|�a�P�ʖ�A�Oe�4�}w��l>Ǌ���,��;�\�w`-��X���F���gu��|�\���̨_
�%l���N����]�zd�,�8��m�#����ն�[_?�m�Z�~�s���y�׮w��w�=�M�f�dh�`�{B�U�VB	��'=2k���޴YM�:�+ʙ�l��K�x�֫���H@KہͥȌ��$��cki����e�؍up&��H{����ȻB�r=���VX�h�
t��p�Ǭ�q�fX[��9���$��`����S^��n}���
�O����_a��\�u����7F�y�R�{�I��V`�Z&�:���t�����,5����^�cph��Sp7(��؀�YX7��,�-dզ@�7au�Z6��7X��E��c�k�G���n,O5�45�;:LvrF���.��m��&�{���*�Ǚ��Ҩ	�4T5��G����vWV�:��3����H"��敤��dw�ˢ�����ͽ��g�l�v�4Vڹ|�n��Z~֍1J��u�L�5��s�#�(�0�s�]��9|#yS0Sa�޹��i۠�����qy�]��n7���(�
�mH���.�#��	�/w�^c4P����f��W\7%��Q]=�h!�����_�P�,'ΓR@�m�U���W�Ŭ:�m9#)U��B�T]��_R�j=���uo\ո�%ϳ�_W_j�2i/�]wC;s��+����|����ϻ�KP�H���E7}؅r��+�O��r�[J����՝Sf�Q���Ґ���۸gF)�|$�־Oq�#o�.�����:ƘRg6����0��S�������G-pׂ���Y����6��2�3��;��R铣r�]5��XB1��V�`�a�	է!7-�Ou���\����Kś���r��ۋ���ێ_cV�v�yҒ��.4�;�\ܵ�d��6+E��guQkt(5m�};���J��b�n��U��Ǫ��˦����X����o�#/7�䶠��;x;]�8�6�nmX�tݛ�&��pU�o�9�o��Y��_Y������D5˩�qt36� �,UԸ�I[5�ȴ+v��8e��Q5�V�F��Ӭ@��J'�G.��5��v���%��6���lt�X1�*�l!��1#�<�:�5t�ػ�>46��t;,�m�(ԃ����ڶ���niOt�+:�sh*N<|
���)�<�գ�T��kp�w��*[ާZ�g�8%[sUӹ�4���/Y*۶��#.�y�U�_�v�\,�qp,����]��*�P��&z��;3U"���&��e��DM7��Mws�5���۷�܀�#�����d��`��׃MŽZhuY�ч��$ux�A�8@R�-�5�2��B"�(�ǚ8[i���c���w]�9/ ��w]�[�Ee�i
j�h�����v^0��w9,��y�5� �D�҆S�9`tȯ$�0�.bEP'0���vm�Q�8�I�A����董6]s�B|�\��t�wt	���wN��	t�!5�QJ��y[�;�;���rw]��eNEa
مތ����Vv��.[M�=�:�%��%˫�7m1���0V)1:Co�����}v$��4jY�9Ѡg#yp�:��L���Q�!��Cp7}CWˁV	�t!�Ӊ�KvV9�y/�ùFu�<��^�$�;T�j����[���{r*f��׽E���b4���G*� ��|�;X��xOd��ɧ�Bs�����uj�.�*��o%�&m;�	 �VO5�k:�u�Rm�;y}��*WsNuţqaR����zF����J�꬧�6X�}L�%���].<0N���ŧNDk�=�� �BC�w�l��:hcA<ѳ��r*���Q�E��n��n�Ԕ���f�go@�+-C���y��Wս�b�	�v]ʘ��wBY�\Rٿo4��W��}k�N�v�*�>g�	|���۝V`�Ѿ����]�xY���u�Ϟ�m�@�V,�E+�z�w��!�5��i\��N<'����d֠w�s׎v�����Y��mk���֕�,�OVn�]
FN�N���YnȓWAՐU�G��\1�êӳѠ��2@��RRH�r�7�{[G��m���/X�48���֞��KjmDQ���R߳:Cm�@뼃����ʖ��`���
n�^H�b�ûR)��c���l�+c�J�v�:���I{`gIr�Gu-O�B��4�΋0�X=;N������z�q<3�woS�a֜Z�܃���u�
X�AN��X�`��������({v��u�b��e\���bt�r�լ���gXd�C�wY��K�i
ڳ���݈����n��_s�N
�^ +Vڼ�v7���ݾO�z�h̠�=\n����=v*u�_N��r���^m�F������Z�}ί�ι�S�3�я
��y:���Oo")��S������Q����[]"�k��-w��7��ݢ�\�x����vk���$���?�m�A�ԇ[�6��J��ch��.Ld�m
7:��:��rBT{ҵb�S��隲��o���Łf[�Q�bZ���ʵ.֓��ښ�1v�N]�D�e>(���3LfF]6��������ףIy4����Q���{D巐9�.�F�w��Jmo���{y���Ͱ.T�h*(��n4�W!�op��4+���ݜ�Z�a4n�[��A.n�f<�ϱ���YLD��m'j�iX��c1�pZ����vb{���q�
� cb��m#VT4�v��#X��Uq�I�r��#逫����u�ء]�:��R�g��b�g;�}0�W��pgu>5b��.Ji%��������f��X1����m}�q)��K6t�U�5�^��?9]t+)�ew*��9q�F�_+e"M2�x`�/(��ѝ�-��<�U�]1xw7\�3S�]�L��@�ZY��;��{��zq�8GZږgp��s��M̛Ԍ5�����\4�m���_.�ċA��&־Gq (��o+xPB"�Q�R��rZ�Y �-�K5���}׹{"V6sJ7�{嗶�KL�¶�����4:g��K��{{�I�x���9`#xhZq>�"*n��+1��Kw�݃���[J2���om-���b�&#K�NէQC���\�����n�U� �4G^+���(�#F=3DU�U<������{��Z+;ݍ�\�h�n�mm�z��}O�5,���ÊT�q���sX Ҁ|J�Jҭ���:�w���J�ɇ�R�m���k����Q�d��j�q��6NJ( �Ê�E�	��p.�w!�i��k���F7�0��7���c�\����!:a�X���L�rִ�;%�9�i�mL�W4�Yt��ӈ���T�b���YV�,]�b<�c\��L�F�^aB��M�򮻘K�b3ٴv�����"�w[�:<4�Q����={A��u2��x��qS�Ww��jy�.�YO8p�]r�+mP_�=&m�N�ч53��Ά.�s��X�	�"��`/E[S6�$(�%�Ǻ���ԑ��[�1r2�顼��'K�Ux���i���A+�ʙ�s�̈́�u����l׵�ުG��H�V�=WS1��+�&�u���
�ֵ��󯛩���7x���I������ -���, ��2%�"�n�q�������+{Se� �r�݆R�[��&�z�7g�[c3t��*���h��M��Cjw�7j�C]�[�0�n�����i�b�`���9�M"�tq��Ej=m#�X�\u����j�T�Z6Q���8i�C��"t�
���y�qu�.�L'�!Q����Uܐª�Ck�)��A���R�.�!_q�o��鿪o��Me�7��0���'--���9�y%mmoZC�M��Yk������6�ݩl��U�V�@�;Qj��Hط��s:�n3�J�g:��J�A0����ԙ@�Swt��EshQ's�f�u=�r����t�������n s?iW|����x�غSW��1�����Y�+3�����f^0�����s��d��j�Q,('y\gݹDAL�[x��Y�04u�2��q�v�+,pKq[
Ǹ�wok�vx���f�h���7���t�ӵ�s�l(���i֛�����X7Fc���BKD��۵�᡿lXV#���a�B�o6m+=6���;r�"eCH���H�l��L޺�1<���u�5$(���˘#�Gr��A��d�NN�rH�Vw`,Ʀ0�$bm4���ͼ���T�K��I�G�l�n�]e.,<X��.R�p��:��#H�W[[�1���,3���d�,�W�z�ʕ�R�{���6(��N��C���8�Rᨑ����	<5f�"5	���xR_[��\z�m�2ō�s�w,�7Z��}�DC���"ݚ�v�a�t��ȭmv�O4>�R`�<!o���S��|V�NX�ͪ���]�ۀB��d2�Ҧ�vmUO�͚�`:�8��]	�#�H�Y�Ҝ,.��0��x����Mt��ٖ�.���+ͧO..$��@A8l����=ʔ�l��7����x��Lu%��=���A2��6��[�}���˵Y�('Ksi�.��ᨺ�����e䣃����	x��ho}�]�8��S���Z̵,�M����/ұuJ��3a�=6k�<�u77_�.�v�cn8��Gk�e��GHj�����t�s疲Cvp�D$�OYE�b�Լ�v�G+�ن�u���8n�b9/gc�D}���ʱ\i����gN��N�Åsb�s.kj,�M]�t6�skĆ��ɵ[ͼ� F}7M�����<b��6�G<�-s�B�QN=p�{�p�[҉7�Nn�e�؍]fh6n�M�2[#/�{��*^jiz4�hh�Ij��]��U��&�[}F�B�{�����jPS��Vt߬s�:�nP��M:�{�].�8�*X>�ZYy��^38dbõ���{�t৷Y(K�J0�t&��������:��z����/:�{�r�v��!]���*�YP��2���޹��^L����:�l����R�GHe����N���Wt#��&
�$�E^#�!M���
��%��w7�1��.q��v��Y��!�\���=]q�x�fm]��fRf���(f��p��{,T�;W;��-��qF ��-�o����<�m�;��(e�Yx���t1�n�fJCE�%f;M�{xM� ��W���^��벓�Lcĺ�����]�ϦPV�S����S��[�N�k�7{�4H��,%B�u�z��[$�M�\`)<��q`!l�٨?�ZzL�h���)>�];�4�^�T˦٥��r�saPL���0�f�;���^�c"����ON9&�&|#<�j+�V�����������s�W0��t�pk��u=�m��"��Ϥ��R�s��y"�Ay�:�M�1rY)Y�"{��	[�I����>��j�,�����/�:��	5v�L�*�����ts���%�I�j^*r7��vͪ����w1��AD2��d����P\�,�Gb.��n��ԔÚ1p�x��i��iq�:�t]�)���B��� ��e�,F�7�f����8e��=ӊ�u�t����w�#�k���U�NhnH1�U�����k�\e*��>cu�Y�w�QIV�xf��n�p<PB���FU�\�LF#��6�h�Wa"%�읲Z�.�
D��ml�"�U+E6�<$ZޜIosUr᧧VL����]�Ҳ�T)"H��k���W(�Ҹ�t;��c��	���$�|q�-�s|8b�B���%��;��V��˥�2���U*�7��R���sI�S�1���K��΄�{+�^:���;Fto��Σ|�Xz�v�X��VG��[��]7 úQR�BM[��a2���xò	�g7[�����t ӟv��n����<��6�Q��s�iyjr�&��(���.���<�yӷ���QW��:s�3w�����^�]�Q������2��Ӳ�����. /",���	:�|E�]�g��j����A	���4�;�j��wn��+:Nwף���k���p��"�Y��-uJ�ڲ���bR�����ǅ�5��6,dA�e�>+h�`a�إ8�/w2�v��+���>��J���ԇ��l�|]��r��"U���5`v�F�q����>�l]�'mK9������O}�Li����v�����=�d���~�f`�n�1N􈯀��#������B�.vЬ�'s�Ji���cg�d��ˬ�S�s��fIR!��;Z��EӾ;$�J�칕u��b,�V�a��&��뫒��2�N��r��>a+�V�T����;i��a�6�*�����;P[I:�1�w1�Qj�3L��`��s��7R ^o-}{B���N���̽o�u�v��	����q���ɚ��0�wG�X�ו�iy{7�u�B�����7:4cwX�8E�5��I�L��mo&�B�uq���{7I[]�	;��
y6�̨�]1(�i��M�z�����(b�Gm��*q%5��놄⺚��DuX(ӹ���t�����|guu4���GJL�E=�s�M�(��e]<�A��ȫ��Տ����D$����{G֧'�-+W2���#��6A�f�f�o�m�mW4p�yo9��/�����1N;�0�1�.�b!�][�uIQ�Ֆ@���ʣ��o9O�=��2#w�&\O.[d��o.��g%�Z�M��W)�H2� ��^fuot���e�&��ufV\����RpÊ��.]Ě9|��i���42�����ͩ�gټ5 �h��u�����}ٵr�,A��&��_��U�b�L��2?�ƚ*�M[��%B�T'�ܓz>&qS[��}��U}_W�|����}�Z�W]<�x7Ƿo(	"�;{2Z!L�`/#u.�1�q,���.z�#�`,���й B�5���l��:+�ھe�t�vʣ����t(e�ʙF.4��J���N����M�V}]r;pd�,u-�mÁ۴��Z��N�.ucz��qN;���N"V�͜��.��vɾ��W������9����J��43�t���}9���K�h*]��R�ˢ:�����6����c������b�+�"m���h)YQ�V�y6�^��iT�y�����]GX:"�e�ܻ�sWf�*(]1�!�q,Uf��\���������[���A�g+�/�8M��r ���V����13Df辵�P�"�[�ڰ�s_Q�a��o';�����D������X�ur�ػ�� mH��B�YBk	�yR�{=�5;p��љ1�952�m��\�%��t�������|7z`�m:8�{�6����t��H䱀c_唗7��%�hЯMl��nt�E˭ץ��6���)$��XT��\�ܧ[�]ua�[BR�-[9��)��;b���cR�.�,`xд����6L�^T�}�3JL��NE���Kt��,�5}��X͉�p5|���o�"�
�)t�ڞ�z�ެ���n�N�F��ѧ�����m�}ي�׭3�:�x��]T��&s��뮅���s��n,�����Fl�"�b�6"!
��c�qqţh�&�#PV�bƷ�F�Q�c F�F�Ns�J����!DlS����1H�Ě��!24h��1��Hq��n5�9��K%DXM%%hQhض�pQ��\k��[��cI@qq��-.sk�'9�cQA�4\\��q���5
")(�m*�d�1������Nsp�*1$`��h��F���
&�dI$�Y(a&��(�����ܔ��\��qF�2D�d������}��Z5�Ѻ�O��I������i�N9>�Y:���x��Ϭ�4J�;	��"Q)�M�z�e���.�3m.D*�����_����<��Ah���TQ�u�r5:`�g�ܼ9�?$�H\�#���7�]x�사uZ)v>�B>������Z���)^#�뷌�=/8��Z�)�N���=����0<̫,xVJ�y���m'�k´/�^>���{	������n��
�>�}ͮ������^b�T��]�����Mp�D}��H�p�j�a�cQKlɖ�2���3���3�>��={�?�Ӹ�\�9�Մ�k�F.#���$�����\V��VoW�:c����x� 1���;�z�֟�z!�&9W���5�-�`��E���0�}�j(�}��*��N
���ZW;sፏ
�/��{�'�W��W�j�.�����ֿn��h%�z{�ۚ 	�`�4eW�&���T��t�v�!z�Um%�t��f?eƣ-S啡\Z�?��$�K _k��4�����7Vc�jwwΰ��5��.=�kO��e������\'��X�aq��@���ՠ�z�y�`�r))�G%]͡.vof�����.al=�����,����WYX�����"�G,{*���Iw��B�"�U�qW����صL,��po#�'3Kv(�p�=ز�d�5LBa��S\�NW�I��T��nv>�0��,Lvv.{�T�j� ��jZ�xgu3�c�芊�T������p�bWvzw��z����n�WS'���@�v�b��c.V&�}X�����ƀ�75�;�Xr�|��ac��v;��p*�����0x:�)]�5M]�
�8�C��$&
U�n(��0��=� �T����i\�pC�TAoIoIV���^��3�=�S<�h��2^�>-���q�%����z�ϸm#;k�R�w&ގcT{5��N$��@��ݰmM���C�ί�b���ef���<#�^S���j�b��Ϟ�"�-βd�6�~e�����4��Uы��z��?jz��JNc�<O���[/}K+�k��U�9��V��8�H�CTp͝����U>鞐�Z���᭾�Lؔl�~���&���T��宆��0�Qx�6}��0=������u�}�c��|?�ʨkq��\���(�o��HR��뗎V���G���N��齽��5M���}Gm/�0#+���߶��Xh���AW m��"�:��M�S/Պc�х-��;�>����\��h̵;��?�ޜ���N�S�8��S��Yϣ���>�V���Ȼ#�p\�9�!��!�u�\��
��w:ƪ��+�+y�b���s�p��"1�ڍ܅���te��L�w�wr!��ǐ�9����I#ǲ	_B7�Cj�q�5.)����t~��׻����3��������j���Fרot�[�5� #u�=Xo\π�Rҫ!��a\�3%{�p�r�tmMD�_�]PKO�^�S5(,��]�id�4YZ}�.�Eu��n`2�n!9L�;w�+N,�<g�QA�g�f�OuQA1���om�*Ǫ���mv�]u�g���Y����`3���c�Mc?\�,��f��f�rڗaSx�$�3�@�$Yن*"ftkV���<.�hǱ�����h>*�e��C%6}YM����a{��mq���EVPG�����t~��~�O�:ѧ�;]��bb�bw>����>D���;��@[�ǂu�Z j����<�}vv�]�ڱ!e'��r���jo�63�l�^IŽ��)���OwM�s�c@5[�ۤ���149�R��2VJ|�U�''�wT�QV\0c+�ܖ�h�7㞸:�H���x��.���2Ȕ�k��yd�.ȫo/���Vҙ�����Ra���L�y?���W�h��[r�H|z�ϙ��Dkj�w��'�\c��W��p�v�#g4V%��^$1XT�WT�βmW:B�1<Cw��e`�>%���`.��뢟�NӸ��j�ֺ7R�����!A&�C"U�YO�
���+K��j/�u�8E9��Bg%��[�!�z�[&�$�����i��V'˗��F�u�'�7����?9`Q����D��c*n���c��cԱԅtU�c��b@��3I� ��+��qb�S���Y�v����ٵ��E����K�T�>&�0zA��Ş�>�J�^���[0���ﴊg.�i�f�������<߂����{��)�Q#c.��=-��*"Ƀ<:&R��{��������{T�c�����U������k��~��;5\� �ٝj��W�p�/O�gc���Æ�����J\���u��q�&\��cw�����b7b�'e�q�R�?f�Ͳ��!�ቩ��?*x]��b��LE�)��:�׌Ǵ�pm������y�߸V�u|E]���QZ�Jin�M�
�T��ï��K�]h��4û}�i��)��ܜ6|��\Tr�P�5X��~]�l4�8b�"�����b���>��&.������d{��hd�ޓ�O�(�O� 7��P�T��dLv�V'6��<>G�y>���E_S��0`�\/6�L�$�/ �}׃�� ]�"���!�5�wRݝ�ϼ����6j!e,EP�Uz�L �C��i�6�²%j����3�����R���X1u�@P��-T��H�߲#�o�D�*���ԃ�%�rӛ[���cp��#_�H�SH��L�"~�#���w*���]�%
�ד���z�vτF����/B�m���T1����J�?I�x�4EoV��G��]��{�u���Ʀ��Ԧ�����?*Km�=󖬳�&<�W����?7n�s<�E}����G���������䆟Ԏ"��4�����	^:��}͒�,4K܏nN-~�0����5���K�7��X���b:�_���2����v�ah�Z�(�]m9�}k��i��I�݅�ZY�����pJ�]>%gSp�[�P���2>G�d�Z:.Ƀl�)��y�����#�-���'���*�U��4�r��ƃ��Pˆ������φص�5����>k)�s�w��1N�z�<�U���!N��Z���'ʸk�;��NP7,�#�綂��h�ɜ����k?5��n}z�
�5�c���E�)u�w!����]�1��XM�H��g2�ܷ�ﲀ��+x�M���S��������s�?@s)�{�$5'Քn�["�2��uh���NҮNw��Qo\u��n�v+�^����3l,Oz�ܢ�ewK0=\�L �9�REw�R��6f���*�wO��u���g�*��EZ�]ٗq�Y��ee�otW�����D���$v�D���Q�p�v��mH���;�{�ݾ���6Ot+�8+�Q�Z[��ɐ�`� Lo�ksA��Z2�ݟ^΍����8���ÆZ�O�{�1�Qi'KG������7B���w������j{�	�s�$';���)]K����C�u����V�?��$�K T=��4��nM������ɸ���L<0pAe��>� ���?1��?m��e��	F� ��xWu%�|�e�N��|�0}�<���L�7
�}(���%��9�aV|����p��#��ļF�Z=�8���{�x1�0�e=���N��=����ac=�u�M�w�A����Z�43}�;α���}ZEktc�����!
I�C�]"~�!�S�w��1;�^ο+2}W|�ӥ+�Kp��N�q�KA�\^Gܲ�GW'9u�.��u�0���U�����>�t�.�~n�p���P!�;?I�v����P�:����f���G��Z_ُo�MTh�&N�n��`-Lr�(�=�%��?<�Xϟ,�ٷhՐ�Mv��(�W�*$|�����,۝��#�w
4��*�gow)�E���}(V�YV�4�X<�e�;��.=X5悇'Ǜݠ���FS�YLtC��+��9Mk��+6�V��7�s�U;��}S:�v�)B�d�Q]�e�mb��;0h�ν��+�m=�\/F�v�{�ɯ�ˀrỡ�QÄ*�G���?��X��)v�{�������uF�͇�?+&��֏aA�3���]1~s�;�c�%b����W�a�䬞�=�C>�i
��5^�\,u{8 ���^�����V�}=����/5��UɈ��z��H�_��.�a9����=��X#�NЮ��Qt"���; \�0͕�_��u�z�V�W]�z*o��~����N�'�����~o��j��d��j����Uz�O��Q��`�:˥��
Q��̞�\_��:.j$�'���ʕ
�+d�}�C[:��d�p����e�[S+���6�+��9L�C�`B��]��p;0X��+��>/7��|��5<��p�J����|�4&�X폮#:C��g��B������e\k�TӯS���"5��ػ�,��&Y���m�ի�K�YM�c��+5����v��^�*��B�A��m\/�/�{>*�����[������d�9����ߩ��܇fwjj����$���g]��T6�f1���j����y��B��l��[���8�ض�����;J��k狺�-�q����f��m�jp�����tD��5>������1d���9��(�f�����L�н�[�"��Ļ����b�K���B}
d����������yP������lՐKG�J�F�v�ie�l��W����.� ��pՎ�l	x��3q�ns�m+.�]�U�:<�0γc4ʈKm�lƦ�s�W�E%�\
~�v�;�q�飠����{���em�*^_���!U핆�]Hw�1ZӳF���w�R���Bw���z��5�J�Ȼ�����`�4�{]X���\���6O�juR6`)���;5Z�}���By�3;V|o�]��󀔅z:�l}��Vc<+�3'�n��+skz|O8�t��C{s��_�6Պw��.!Sg2��[1w���I�Ec���R��C~j{�+{<Lݗ�����!��T�磻}�����>�(;#��*պ�~���j����ꎈ��<=1��ۅ�SZ�Y�q�W��]f��0P�g���S~E�x� �w���^�E>�%��\G�m^��T�w�|}a��x{�I������5���6���@V79�aƫo�����/�y˾�/�O�>�L��U������:�>~�Ab�z��Ǹ�=�uʒ6��*�'�fʭ�w��W��S;ƙ��qӡ�!��f���(,O+��'qf�ͪ+����<�\��7�\*�e����pF��5�8��zh=��p|�:b.����hi�f~��V�%��l਑^����"*���|V��[�Skº|��î�{��״*�a4�=����N.����d�p�EF-�J4Հm��0��ht��|X�g�l�حmLe/bu���\f�F2�����6�e�w�M�V��jN�!LD�a#�|,կ$��-��z�b6��>�ZFxH8
��'{.�o�^8/�>/>���î� <��R�w���������fpX���uMV+��vُD얏�����u�v̋�L�w۱sHBR]�9�%7�L6A֦��)�=���P��y�VY��z}����x,��G�Q�=��Zt�U�yU�����ȡ�i]���\�C�5�d���hQ�6UݝP��'����̊�=ʪj^G'���G�����O���ܮ���,�(��|K��m��Sm�T�<4!I�����#Ɔ�2|�e�����
��;��9��Q�n4��5��A�Ӊ�������lҫeQ��f�~�����J��A�a��=BL�����o	��P�v��mո��%��h�'��̨:�Z��[���o-gmڥ���.�n�n+��4M�W���J����{�b<mc�c�kw���ɹЪ��Xn���0*���Ϭׅc�y�s�k8���+B�=��}'T��X.�+��M�����L�7�ٽ˯�0�c"5��g�c�bw�Q�a����Ly,7T8��h���˺Iw�a�j��2�Ωr�7+�L
�5�`�������Cua/k�F�\kXV��&2}���;i2��X��B��N'f}L�x1c�[}4u�p��m�f�Pl�!n3�5>Ϯ�{^f�ܘҾ��c�}	dOdF�=�c���Sʎ�:[=�KǦ�>-�nk<�}Qo]q�l�G�����v������!��n�Y62�]f���ql�ګĎ_�y��L\»�;��\�Lg��Yz.Ϥ�#�����fx2߃�{u��V߳I�~Ud|�EƔ(Mn+zu��<~c���!ng̿�	F�;*���I�kr�5n� )�03�EL������ń�;H�#�z����:�]fԬ�􋧝�.>^�}p�t ���WP� :8�ڝ��~x*)[!l���0�G�B�
���Iſy���惮Y��k]�P௕v�yF�3 ��m��xf��-)]�K�E����%�]�r���:ݹVsx���l^��q����u�h;��:(2d�76mw5�;삷5I�����ם91��-=��������{r[ӛxu���]+AU���b�f�+�EG2�v�<]toB�o0����h]R�G��W�N7N�+�\Σ�c�_�� �T���\��&�ƻ����jU��_e�����{VG9Gy� Y��X5^3Ů��K����2���K%��F�ZYל�U��J#{Em.�HQ�"�ȱQ��cn�*h�+'^��V��u�XA��\��g��9����\p	H�:Xek"���Ɇ��|�\��r^즹sF��,��{v�`-s��v)Dܰ��c���+���ɴ��Z<�c���up�|��q�s7{�B��j��_dt9wȽ�1.%���-�>��,&+2�p��VfTS��t�x�]M��^1^~�*�H�����K��{�-ˆPV�@��7���!gh.u�#�ܓ��e��,T����N��Ԗ�-�;.�-���;���P�Y�A�o:�������{�u%-\�H�Ӷ�VKM�K�^�m>]��_M�e�ti�����y�b�������;8�
 �j�ɶ��ݮq�3��ҏr��z<�=B��ᑻƨ����k��/��{�퉁hmM�mݙ�Q.�Z, W ����^we*�do
�>J���S4q�B��j�ff�g_/-B�i�΀�ͱ���F�X��,S�2cT��S���/���<D�I];���%*�ye�+a1)`�ٻ�V��S/�X�n,w���Ͱ8��	e�U��=+r>߶U�v�S�7��,�=<l��C�[�#�ućd�f�AS�#5�.5�B�v!���|6���z�u ks��v^.�h�Q��o}�Gٶk^>z%�]���=�M��+BRZ/��F��������!M�� ��ǐ�W��2���S�f��V��<�&�I�|�&�vr������*��Ñ�����t3��93&�=ՇC����X"��7�]r��l�WR�`� �lX��3,����ӕՁh}J[��MU��i�m��MX9u0�G����!]�������q\úNE��a@��ӇT��X���w1wj������\)��!�-b��I0Ć�7ug����0���'�\5����]J�-]<|Pꊧ
�}�3��ڎ��Q�]��f�)]
��]���P�u�����]\F�"£Qn��ڟ+��g�a5��q�Z,��WWZ�����q_\'�9y�w;nN]�7�
�;�m�F�s��flN3����=�f�A�{��,�茳�c��ږ�Թ�E��a�צ�H��M�--��8��j�C�����6�)�G9S��]ά;|�1'�q�	�/V��Cf�G%�;}�r�რ��rIw��|'�}��_=_��w��\�ߴb2�S�K��F2"$Lȸ�$RIe &A2Kss\s���(�!�	I,���!�H�if�9�F52��),�-��H..Tb��Q�P�L�#&%���9�Q�D�0��"�I&EŹ&���R
�8�&a�����qS
*#d�%EF�� ELE&�" � 0��$��F�d�1Hb�$��3 )���*S 2� �L!�F���I*&1�S4JTFd̃(�f$�($�R@�B ���}�߿������l�+U���;ȝ�崰0���[H��Ho��ĤŊl���x�
��i	}(��t��P�B�o����ﯽ}z�����v����g��鮖���5�+��t�{�+�scq��+��.�qq���}r��6�����}���ny�{��v����oﾺ7M����������1��Dn4ݚ�%��u�����]ys�[�+�ͺ]z���^��ns��ߝW����n׾��\یU�pU�����\��w�-q���W�z^-�t���+����������^��p�����z�{�炷x|��x򷾉��y^}��.�t���:�zo���7�\�KF�>���E�+��������-q�W�����o�Zz�7M����wu��]�F��W����Q���T��d�Pˢ��h���H�B"�O/�j��t����;���k��>�^��\j�����x��N�t��m�������9n֊�o���n���q�����n~�m�.׻�{mگ˓_����{#�óۻ|�q�u���P��>��+���m���}[�x����o�[��_/�}�����~k�}��w���ţ�κ؊��WM�ۯ���n����LG�DX�>�D{���t��я���\���4�ˉؕ� A|l�q1�"�}9}k��]��ۊ�.K�o�M�j����Я^�����<m��~��ߛs����[x���������ی[�{�"����p��q�P.��c5R�:��r��G�}񆾢/MX�T�}����_yn���]/��\�t��G������^�v���ۥz�+��6�\������h�6��<�騷���tG�yE���M�]oe�焟�*�+�������}|v���ޮ��n*���y޾5�j7��η�������忷�Wm�]7J������hߕ��=n�x۵���r�����-����[�t�|[�*@�� ����������}��է#"��Ρ��#�#�G�?D��+Ź��}]��[��j�.K�}�|oM���yֻ�ͻn�ߗ��:[���|��~[��z�m�zZ7��뗈��X��"|��~!�k��[=��_Wj��^��ߜ��o�|��v�.6�_~��zo�sn��=s���mϼ�]y�|WKO��7�r���}������6�龶����t�o��w�6�o���f����y���� N�ޝ���כ&�SuβXIL�۾&��_��',��u�x��l���e�64�q��(S�ܦ����l�%n��W	��Q·�K���T�֘1ε�N�F$v�_L4���R��_K��hJ�[��fq[o��P8]��ے[�s���i����׾�ݣ|���� ��X�|�W�^6�یoy�M^8�ߓ��u�6�\����ƺ_���~�o��]/��=�oKE7���n=5�]5z��]��pW�!^|�
�����Y�w�_�6;�4ז�k����U,o���z���oύo]�֯�|}[��請m���w��W���~[������E~m���~����"4Fi㗳d��e܏H��=԰����qh����+��+��~���t��O��t���\k��]^>��h�w�Ż~j�^��ڻWչ��6�������6�K��z뽼n7�n7���mߜ��t�]=����:���;��1��tD���n��^W���9k���Ξ���{o��x�����^��-��(�����w\�i�͍���>���W�����ͺ�Ϳ��v�o������V��kB�Z�\�zlUB�*��B�;�s�� >�ۍs�7������k��]�;.����Kq\{^y�Z�����ݷ����|ۧ�گ_yt�m�sn0j5x⸾��v�͹�,W�񮗋{w����]��}��xU��� �X�$GG��"=-�����������u�[���,x�6������^���:��y�^6��o��~u�_ܵź^�ܻ]����Z�����n�!_xpc�G����"���~��J-߼9z����,}}�dG�!���7?�����v�+��^���u��Ѿ+��oM�n5}�����-⸽����o���y�Z���q�/<��{xۥ�,���I����a|U$�(��U�%�`��ߝ~�W�t�?s�^\��zom���~uw6��n�pj|�ޛ����[v������|�w�\o�z�۵����_��{k����r�*"��u������R��(~�}��y��	/=�r>��n�qqy��ݷ��n�s^��t�o�7>�ݫ������ۍ����^6�tޗ?��-�{��W��ߔF����F>�>��}�'#��8�m��R�>o(�4/�}�|&���o�58���Z��+�v۝r�_yn��鮗ֽ\���hߗ֝r���E����ݽ��]5�z����ǋ�_>r���>��ƭ��}�����Vw\��oWWJS�C�,�ŖX���s�)m�����8��)�s�KΎ:WA�;y]�EI��z��pѭ�]hg�Km�V(���W�$}�������n�&�7��9��b�!��U���;o��
{[n>�{z4���n�wV��_>�w�KY�në�n����/꫺��?�{�K��:�ʽ��W�n/�����j�6�����k��5�_9]-��t��z��^�k�⾷K���|^�������ޛ��m�n����{W?��=}<�a�e�լ�O5����}�˯��������ƿ�}w޸�|mү|��^-��j��;��zW�s�|_�s_��mŽy�W��6���}]-9ͽ7G�G�}�DFɎ�>�>c�x
�>�γU����g���0}Z>�H}T�xk�鮚���ʺ^W��������m����ޛ�źU����[x�7��m�1��#� B/z~��h��=0|5��t�ؾ�љ�3�u�ԝ}P��#�����]�P�Q���G�����@� ���w��z]r���^6����ڹ��m�so���]��U����[������}U�/�x���}o��A���#DD@�n�N�{=�]��*_�F�B��|(_7&g_y�>�P�&�/�����U�q����.���ۥ���n����w��]�6���-���U�zm���_����kF�n=_�u���^5�y���#�#�H�c�r4g��<�x������;���~n�r�⽯7]�W�]-�9�_��6�_=s]q\[㾹�Oܷ�u�뫷�ޕ}\o{�.��x�ۦ���W�p�ͽ~����q_���aޯ��`��>����;�tq���]�.�s�.�ؾ���|G�>�و�@�;/�s��[����~�ֿ���-q�?�uֽ��M�t��~�龵�鮔qh6"��/�t���v��7��H����b��p�����Oxe
���+T��y��t}G� �{�_}l��"$G��+��xۡ���y�Ү���:{��������{�Ϋ��5����v�۵��j��ۜ��_�k��t�[s�����|} e��z�>�>���8r������+�����߮�q���~��V��-��u��������_�uv7�q��������,}^y�ޕv����y�z����J����{mιƣ���DH�>�D�����D�<^�Ŷg7�G�ۍ���_ώ֍ż�Εx�׍pz�*-�.���έ��Z�~W���;���]-.s{W��m����Uv5��5��:�^��������W���n�DP�����5�:�@�!Ƕ���'R�v�wwN?L����g����6y�����i��(�����r�u��6�|���<�`����r�',�f�7^<u;�Er���[���:�Z�r����~K���f<ǰ�"��o�]��ۆbr�`]K�-����u����5�t�ۦ�ۊ��?��79]-�q_��s�_�����zm�m�.��7��9n��9�>u��}d�lG�"
1��<#�<>�t�1�J19BC|�}�S�7�/�.�~_���j�tG*�";�Z)Q8<����I�>���.�߇ٚ����>�|�OZ3׭��Z���@�Rv�lr���:���x%#^=�\*D��}Z$�j&�U�n�c9���W&����ܰ0�}�1��Y��P��l�9y]��g��&7=���Q͞�u�o)^�;^?rwz}���ǌ1Q�uC�d�f�1R��r���U��6!��֗ury���+����h�n]}Q�S\kqXϱ�1;��0�ŃeX̫��0��-�Y�˗��ѓK�jBՇ�3�漸��z�
��^�=��������Cua ey����1f���ŷ���eZh	U�U
�����|<�o��"�w���R���;�r{ ���F�(���a����a�޷�g�c��'����mV���l���eC`;��U�a��M��oTψ�RJk>~�!:"�>k/��5�K)��!�����7X��gF��k�gbw0������T`''NM��P���6��k�����	��n�CW�=����7�M'�F�
�ʅ3ʺ�V�Vm0�u�n�u%S.�R�&>8nKڗϬ�z~!�x�OQ��j�/N��rq�9]k��fͶ�>����)ƍ_��̡�ᮘ��Wi�&b�Z�3Ы��
��v�����wE�Oj����<�d}?��q�E	�t��!�x�Ǜڄ6�p2|%��zR*�Jv����'@�8�1$��Z�OV����N�"��Bګ��l�6d�'���� \�5
��S � L�{5���:�����P^��������3�Kc��Ov&H�������P�+���� 8#�z�xv:��G�� ��p�>��=�ޫ�l��c��Q��.%��&��A�4�tm�o������U� kݏn�8��6q}aߘ���Pɨmւ��1�ы���Snf(�NO��z/D���䏢��,��}���Ng�?T�o��2�dɶ���3Q�DX4��Ǻ�/�.J�w���Ow%lW�9g�X��L,5�m��juB����n\Xg�;n4��0y�W~�%�s�x偃��5Pj�%V9�k�l6g�K:=�����������ӗ��m��,`��~�N«~��4�/��Y����X���-+�h-0�19zIYfǹٯ+�3%H)�``�����t���Q��if�.9ݡP�ph}�:�D9so�n��Z��f��J}�r��B`���*.y2vô��D���}Ջn�7�=�v�r�K��-W��rgU�{�>��#k��_̱R*�[�}u�ܚ/\��7�Z��w�z�N��[�u�~��y�ľXN`5����Qj�#�'�k����P�ͦ,���IL�7Z T���u�0-L1���EƼ�g�c K@qcڃ0�7��'7��/as�{����  ��u���u�<1�cwW�����di�

eJ��q�Q��p�gh�%���.�S�~@R�j��ʐ7
`2�S)�u?X�>0�0[��{i���E��3�X�Q�爃�������v�L��v��B�L}p�:cއ0<7�uz�T~�~ֈ���M�f��j����ӄ�e`;MO��puI-뮾�Nk�ǀP���%�2��8m�ۜ/v��u�N�b(��YP�>_5���I�z=�Ñϝ�e��p��\�|�/tqe8��Q��i����W�@[�����W$yh 
���`�X��&vz�Q�M9\A�U^Wxmy������.pCD;�!�q�.� �ICd��=v=O���,�j���N왙�Q�ѵK��e��#Wc�"���<�]����|[���0{+��gE�	�h/��9f�����N��N����w]��n��P��%�2S�,��1�p�3oE�����&��uC�V�g�̦Ns��c�o�5����n�Z��|�O������1��.|�^���Sul����Gy�f\E��Dy�Fd�c��KUx!�3y:�源�5&+ZvE�1b�[�rY{[�z{�����)���;����i��ubR��.j���{�!�z���5��)[�Իw�`��ր������/W��-Wl��|���3½�2�`ʝ�a�n��[~3�Z�V�8�:B9�bB�KnhS^�"��v����̨W^�2wii7�Պ};�V����ҙ̭����0�Ω��걟7�jX"��ӹVw �y�e�<X�_D��=og�'�UW=�����,/�/x��~�z�w��0%X��:%;{�
�:g��lr��(͉���.�V����X)�&_�����N3J�� �[���sG��W���tn�ߊ���b�.C��i�m�Δ�>�X�[8��V]wʳ���>�<�~����M5���M�@j��iTV��^Ҹ�]�_68w�Ւ���x�ST�\�V���r�����oU���v�3b�Q�n�L�{�Y����:��ட0J�u���d���Bx���+�̍^v8й����^�kq���v��!�cr*��r�fV-y��i'3����b+lR�hN�����ﾞ֦<�w�5������F����o�ހ�-Ŵ̊F��`��؁�N��R��	q��^r{gFXx}P���<�g}��p�xo�Ho�u��7%\) jM ���]jr�\�|�$>��Q��⵷
;g�ai�96��܄~�i�ʬ]Qu�x�=�n'X�<]�Y�'��@��������f=�엇М�
~u�܉[?;��_^���lm}�&V���M��Jݑ�&�Ҙc� ����?*�'h �TY�u�xQ�j��y07�˱Vh���C�S�+Ⱥ�H��Ai4���[=����|=+;�z�^m�}*ױ_o�K��Z~w�K�r���",叽�rv�i�m��v�f|�xZI]���յļl/V^5��B_��&���"����Fhe�0&6Q;_����ܭ�e/y�O�P�;=|]��
Ǚ�^*�Q�u
�;�>��'��#��P����%!�
Ь���4��w��7=�,����ڭ�0-��1�~��*s�k�O۾���=;m�y�3�S��u�2�x^���3D�WXɽ�e�N�菳�M4���=���,JM����@w)ie��%�V���L���'M��{ח�������܋Ľv���<�}�4';w9�����6hY�PY,�*t����{����}_WX�l��-(��5�Q�ܱ�S��+����Sz�Z�*���뿧���k�	�,A�t�ʾ�u�t��:����N�!p�l���{O�ُ��X��M^K�x}��y���7yU����;��bO=�i����3T3�xT���6����y�Qa[��zc��3N��q��ܖ?�� N�nk��W��у<���}��gI:H�=Ek��/_�9��vl:�R#4��(�}�T��@�L��`���L��T�)�hժ��\Q�I������v�q=�rwGw�6��˂*K��(P�X�����>��ʆ���|ˋ�2ݨ����^Tފu[-�ԼO��Q�1�At��F��ε_J(1a�:�8��֣��<���2��ʞ�5Fg3fF�րⵄ��J0�ru�נ"wΰPR��٦��n`5��wU� sO�x�t���|w�J~B:�$'�)V�d�v&ߝ��k�'٧�S��/ԗ�zױ��ԹZ���J_���F�L��LŸ��=e��\�}n���ːxﻠ��{�����������c�$��X�U��[�gr��Y�K�
���/W��җ����}u
�f��
���r���^�zƍ���76ۺ~�łc�<��4����N�^�Y/�nNה2�.�j�=�";�y��x�qi�ْ�a�߫�#���ϐv%����w�2�b�f��%0��mւ���F,	���s1Ub��=�j،���#<�}��z��3�o6V�I���=�)�'~M��`a�P	�ֆ�'��X�=h>ٽ���^��1��~�]�aʵ]����\��x��>�'����V�=t5z�U憾�3l�M`��/��y���~>����d���B�	KˌJE�g��3=�������_���a���ٳ^��1/�)V��V��{��+�X&o_���7��&+���z�T���K�Zɍ���|:(������Sc�]��E��g�+��#�e��/V�3�GY/�PP��g��L�T�{>o+D\k��k�^�?p@+G��C��ɓε�[1?K9O<���H��f�(1��Ye�|ƨ���e�wTy��:=u�z��+Ҋ��g��z��5�tGT�����\S�4Tzf��yR��ex�r�^�j��B�TW��A�����J&u��شQ�QA���+�:�]6����0��鏮Ly��֜Ɋ(	>���������O�f⸮�4�KJ�#���=P���,���w(��ܝ	�5w���i<n�W<�镉��vVmt�l������q��K�J��`n�4��7����}v{�J�}k�S@'��.��w��M�áA�������|'����Y�E���G)*�gw'ύ���gL�X�x+T��& ��o�s���ӃV/#g9���';�F�3��,�f���D]�1G����k_hpM�d�ȷ��M�U+V�Ӫ�A�xś:,�Q]CM\/����ng�����[3�9!�9xV�RԬ�m�喙��+eÿ.(
�vHj�ڳ�fm�wع%v�ۙ�Cm�M�8���:��I�՜�_G,�e�UzfnLZ�j��w���.�>R��#α�՚+qd��f�u�'T�K��;n�.e�-iss �Ն���C]�������Q���/(e���T5}\�3���_e��M�Ǝ�X�.�Zk�>3��+*ul}uD\����Mۢvi_;�2�(�d�8���F=];ol�\�b#�ʹ{��;���@bv�֬*�n����y�ӜȩdN�Z�\�y��Ю�ذ,�Ɗ�">��4L\��ȵ�ʆ�+i�<�u)}���k:ӁN���]8���gm٫@�bR�],��`�{u�/��8R�f�N\9;l�Q��Ư�c�٢�P�����|���;vz�:�cFk T�&�>KSr���<@PXt7����Ѷ�c�b�����x�Z�q	n���w�K\��ɪ��0������Ch�I#���_4������`�t1m�x(���˭�8h4/�mu�6����^E�D�-A��p�/mG����y%�{p�J�֖3;�RǠ��1�j�Ԯ���T̩��}-���N���Z��>8�.�j���ٜ���n���SKg7g�q�P�4c��qIk ���/,�	�Z*�^um���r�Y�3c�㝊h��Ij�EU"&�TS2���ѝn���	;y����y�Wnè��ĩ
�w��ЬL)��'��d����l�s� �:�� $�����p3|��ݰvt+�o��<"�
���r��:���P4�TV^� ��>���)�{��VyVG���$
�y���k4��[T�:%�^>WY-�K"�EO��F7}
��ܡ��*(
I��͙�E��εK�
��d���<�$=-�72�i*̀p��Q���B*�^֣8/ahWc�5/^�9�mU+c/�Ҫ�i���wke���.���k�4\-��+	�ԇ]�Nk�9-p{ͭ���٠'���F
�G�����]�cʻ�������!o7���+!�c*�݂�lTE��]<��r^���<�:z�����W.�Ge�_�����>y\ӛw��6z��C��T��k6�e[W8�W��uW���3J&&JXPQ�����"�(H�	1 H"#L�2Q%(Pl�4�(�l�
a� �l�`��a
,& (�� ɤHKa2I ,)CJ��
()JI�"��Pa��HQRBd�c�e e$Q�``��D��&#d��"1	L��%�E#FA"L���Ș$�ɘҐfe1�ƙ%i2���L*d�D#�e!0�Q��&��f� ��E��H�����ċ�	w����u����V����P�w���l��P(vF�j��\^F���o�����#�orWIv�7�횺�a�]���}�Ճ�Z����-���i��U{5���"���LQiK#���ک��gl�҄;H��)[�eeC۴Q�ѭЃ��%����r��h>5۸q�2���T���$���{F�]���~~g��U�]���ú{qW�q���=8���+�`2�u�N�����V�jHBu��O�ur��G|�Ӫ���ᷙf�F�G=��)���Kwt����Lh�βŸW���\����6���}sî��u����%��k����8r�9�ly��M]���JG�8�F�{��i��Ԩ�\��1��r��i�^�f�1*����Ԙ֝c�u)�;�T�%<�|�o�Yut��͐l^GlL���YQ�r��՟2�5��&�o�H������c�57�}��tI�����}a״[@�^']U�(,���H��^u�jw|���C���}�2_=^��Ѝ�X�3W�r[22��_ȕ�+�m�\c����_Mb��H�����.��߾K;���>�V/��r1��T���o�\wz��#�هiF;���ݙg���^��d�
��nu$*Z:*;���md��=�(�"���8'ڞD�t@,���+��l����y�姻1��cB�Wd��1���Ys��N]Z.|d����h.��6��q�}�Ӥ����Y��u�޿����KO�`Ν��d��TE����m�f���g׌�&8�W�O����ew{2S�o��Y]�o�r���l��/_q1��-9(
YZ>����X8�.*��r[�4�zm-��[�u��e�E�;�]A[��F
��S�b��j=��Δvv`�k=�Q-�z��Kf
�Ցo�~z=�U^��u����OݥQZ�O���1��=��ۼ�m���S7�;<�7~A�-�t,t���z�/|��i�d0�0˰m������q����u_�TQ�zW��>�����ݎp���~;�ͤ5ϫ�&�R �){Բ[Z��z��#�4�d�߬�>�k���7�pe�Zq�#7��r=t��Pڙ��0�|���Yt�%��DLe9���@:Έ�����N��'�aw���y�����x���
"v��,�<��$����@�T�y4.)L1��6���$�%R[�Yy7���磶LଢD�l/v>e��Ϡ�>Ԉ���<��{'x�z����拳�joƌWw~�Ouɼ駫�ۚ0��{��3�O���}���4��d�7�ٯ���{�@�,�Y����c.:{Y��ު}{r��U��f>H��qp�	��sD�^�@o d�j�Cyi��������^�yAaS*X��ZOu]r+�W�U_W�ɯMYڼ��̏х��6�I~�偏�DX�1�漎ʠP��Gmӥ���r�^��s.��\����}��c��W�}s���#?Q����J��m�s�;c�d|�����=\��v��)�4���#.��-���Z�7��y��� �U��}��O�6u	�B�J��{���<qxl��v�v�G��0)��1�~��*W?S��^)T���N7����5�j���v���M�R(�8�mXꞖ�C�Gҧ��������^�����Sx��+�,�;����^/�6 �͹=S�p�LK6'@k����\N���FP��{�Ⱦ��2���ݸ�ؿ}���Z�����ٌ�����4֒�n~�N� ��^,���Σgls��,�&R��U��� ��U��g���+�Z0g�����3�� �pw
�\��:kQ~�w�G�Qu�|�4��Yg�lG-�Y��?+L��u	�Q-S�Yz-)���B�//�~�;�xv�Oy.�[>i��H���ޟ}�C><!%�b��6$�eF�o�wE�j��C�c�Z�f���z�Ế=�:�+��z�#VsH���xجR�ow'��	[¬�`����U�5Y3�Ex6���%����έE�k��2�\>�^VP�cf�p	 ��5�J�ta��E���$M|s�_U}�UT����~�o�՘���D�' CV�C�ʱ��ڵ_M)A���v�JV��s{sM�_%ժ�A\�Y�g;rnϔ��}�%��+�U@� ���
U[~x�ᛍ��s���������Ap��{� ��K��/�V�C���=�I��_�)�������/e���Է��_$ա�9Z�x1���n��~~�(ÿQ�Geߑ@�g�e���佾�#Q��g�7�&-�Pɯ��Z�u������s0��� ���!X�m쀬�*~���U�R���͕��S5�'�SR�2m7@k�5�WH��-��F�7�y)�Ǘ(b���"�|;�oH�B8Q�S�N
+�� ����e�+�:u��^�V
[�����(T"��X�^��<kj�p�(1��2���ʼ�	�~��Nζ�����Oez�5^�vl��8�=��M��B��nW�߯�XTϷ4Z���}��+�� ��2��\�7��}�h>~��;��&2���'��{چk�8Z���aƺ�(�t�������� �ce�=�Nw��Yb�����q���l��G�bhN!���y\�= �d8���]�Ƭ����K��N/�[1j۱|m�✟,���^(�H�R�yN
[͕;�F��ؒ����yn����A�{^��Ա�ȡ�%�9p&c|���Ҫ��jHc�f�o+D]O=��qh�_p@+W���ymw+�Ez�^έ����*:�T��1��ifרl 7\�,�w�=1�7Q����3vF��j�7�i{�5tӘ4)`�������iW��ρ�r���gyw�B��+����G���������QⰐp�P���H�yoZc����\���]��w< Ղ?�`#��j���#���R:IU�Q�j�wm@b����n�j��+�Iy{��0ǭ�%{���~C�'�h6_����]�����Ue܀��OD��0�������޽��3[��R��ONbti�0�!	Jd���H h�{�6v,	�n�s�{�c����)������a�Y�"�"�������n�,�m�r��^��L�&���3m"���5w�n<�	�LM9�r�l��01���G�f4C\������k�[�Z�u/eI��:�=��%rTBԈ�L]R�^W���Wx�rC��R? ����.Qxc��ҙ��G������I�O3�R,���G�Ơj�[�T
v��N��[�&�o �э�4����W!N�y+5�n�Ӂ���=7{)j���]z�b�IO�v(��Hs�70w��K���L�f)����P`�s���s{zI���}_U}U���	��=z��?�R��J�ut��l��.G`K�`�k�Ճ�б�߲>��=�^O���Y^y;_x8�wr`)����3�����
g���tw����$����ɗ��#}�8V�'�	�v�%wy�S��3A�}8��h\Ȍ��l=-[�u�K-���ٿ-�욥	ҥ��ǄxW�-�3/m@!᯵��b}���w��>�ȏJB:�9��LW���x�e�V=>v�=����UK��\h��Lq8_wL��e�q���R=L_�w�T�ԢF��O�ߕG���ü��H{#
!eh����X6ٍ�܏SJ�=u�6����~k�fw���,Ln�+���^(U�C��i�l����2c�Ŏڹ�g� ;�V�z���(v�>�ۘ¤d��pq�4F���U�:��O�ɝ�m�r��@+=�Pcc���ΐ{.�~;+աxc�\ F3��3}��YkRkv�tdƺ2��L���YT~��b���d�<�y���e���rU�/��P�V;�n�3yA��l�u谶�<�����cr�������a���>�*$0�`ܮ]�Y��# y{�q�fEo"йtď"A���+͍>M0x�]�ui���n�Px�N����N��-M)ъn]�����&#{ͦ]p[}٥h���}�W՞��s�	� =rF���bgo蹠����5��p�w
����]��/��@���˫y��֎{z�?a�N{�`"�Qt�������o�`n]6a�y�=�hza�ɘ�d1v,���%�X���x�Q� wؘ���^(�;����Q�@^W����F�=U��� E�q�EAv�&ї'I!,�N�K�pyL�V(����vg�m�w��!����.!g��i.`y��"��鏫�R���2�;ꄵ���f�RV�3��ȸ��-�Ez�mFk�['�ly5W&���nXZG��#��Z��{3��&������zvt�;>���oƷ��tsИ�j���&�ڗ9,�rI�;�q��nN���[W\z0�JxՊШţeP��5�b��&�O'�������y���{�˦�F+�%��[k1��ה��pv�(���jM��WƷ�۝�iM뽦�ʽm+���+�=,��_��y��Nk�Χ����5�e�fW��>�<S��k{=b��y�3��<2�FI�(�vN��̺v�i�>&���.,W�r;��ΗvEm*�����0�Hh�(�h��^��З2d�s(��f�I]��:�cU�k�F�Ź[Q�OU���-�R����vv�f`���>����E���/�}�G�G�M��k37���ݠE�N���=��@jy�O��D 9���wS�V�J~��oC*gOM�I�s���� 5c)�"�ŀ7T�sN�ҧ��{������@����y�rnml��ud�3u�}&7P5���axk�M�0C֝�fRǵV^��7���5�-������=�4Զk��$�K Cv��T��X�m(M,v��!�����6�F�� �Oß�j�{u�ɚv�������1�A���Y�K|gNf�u�տ�t�>�*���G�8WE#
��?y9�!�ʅ�2�� a�jt8V���9��.Z�.�r0ǭ�_�[:=���6��NJ~��`#:D������e\g�A�Jԗi���U��a?:�Ě�<�+Y�0x����_��n��i9�����UO�9���[<�$ɣ�'�j���߹��G�C&���h/�``��b�n���?g��'lE�g|�K�.ώ/����z}G#6V���}I�AJdɴ����YVpxPG����ej��/a�0!oH��Jr�i6�_p��u.7��F�4�h�<1���,w���7�b��V�-|�ִ�{����:�F�r��#�Ć#:�[�D�t$�.�^#Ο.�C��{Aj��1s ƭ�f��Û�o���*�~t^�gEJ�k���������]t��xٰ?�@ؘՊQ���K���|��Ö���벷�"5�v�gp� {J�ŋ~��?����a��ь�#e�i�5P��%V9�k�l?��xRc�,���΅�f#}��{�-���宀�Qna���ײ���eO�B*��hv���"��Ύkس���6����u\.p�]=s��`��:�K�]֬'0�_6.NG̀�Nz�1r_.��}�*X�x�� Lo���U�L1������4���d���%|\�Yc�u�'��m�TW:���3U�/�k�l '��Z�.��5Azc1�{rlH�������)*fk�t]KGM?��KO���U)�C���e|/�9P��:~'Z.�_��!�ҥ[�M�T��K��
>+Ir���@�\Z�Jm=S�順m�&=�Hޅ�ć��`t��`3����ϴ��Y�+�t���.zP�a�Gҕ��-���]:u8��_��X�ы���2؉-�����T>��j�9�]��CW�Ł#(a>��K۔��{*&����"��n��4�u����a=򙞥<sǅR�v�Nz�@_{&[;�L{z��9�MEv��6ͳ�p0�1s�yU�j������F�I�'u���k|リ'ȫ:g�����������8�ۿ/.h�V����������ҴO�z�����q�0��&��S&R�,��W/T�6��$�s/�lj'�gT��Y�Z�I8!���^�w#�=��)�~���\���	� �͐���$,�C�g*���KXV۹=���ƈc,F�%��^�N�W���Y6��^�(O%D*Ԉ��*�B�l5w��fw4==5���v-L��9;&�U�Y1И�jM�mʓ�&~{�X�9�Y��4fL��Z^i���=�|O<��.Wr.`)������[@��;�B�vʠ��˯�1�q��5X����H^������e��ǫ҅���,r�ą>��742#х����3Ö�y���^`�>��:�v����ҽ��x�=j�����m�z�RuLN{����+���[O��qM]�^p*��#pv�=-���,��8,�����*����y�I�<�m<_hSʌ������z�5W�(S����ֶ�����>�!���@,�O��~Ë�5e$d�av�c�Co/M+��X�^_��i�E`X1 ފ�r��3�P�n���8CܻW5e4�����������{ Σ��oX�u����L��s��+~Y+�\�5-r
��I;�E�F�+p��= ���&�`]
J��z,%��n1���r�_;.����,����$v��\ʇ2���\�w]LT�h�
�+z�ݣ�n�!��N���������Kλ��N�z,oh�Z��R�Cu{hm��[����e�s*!,��(�W'�	I��ٻ�!�-/��3�{�)ڒ��j�����Ub�ۂC�ZCZ�¦�Yy�fR&���5���a��,N+�3_Rz��SG-�
�BB4�z���aǪ��d^.Q���kހ����Jwp�[T2��d�ƙu����]���!�ҹ�9Fu��0a�B��t.���D�X�l$mb�M]�%Sl��.
�ն������^�r?Z|�q�Vnmh:�E�Eft�F�W0гy��UE�l�՗y���ڏ .Z1�wu�p�[,C�a�%vq��S1Ғ�q@���,! �)qM�9�۸)���p�s1r�}F-�]�-�R�r��f�g����P��1�BW7}�β!���ݚ8%/�w$Q�s��cU�6����1�ko�~�ȁ��a[�';z�]����sAӶ��+A�ǗBS=XD��C�'�U��*��R�@���X��8S�U>�"��̳L�hmbS��6mf�;H���@�FoR�A�cʸ����6
k��.�sb�`�u�"��չ2,�Z�N
;��F�Zx�͸%36��40jُ�]�aǔ��r!i���t9�� ����߹��L��2�ږe�6,([�Ś�]�h��P��"�ە�|_A	4n=@�3�
�̆�9�2$�t�+��4�#���=Wssul�KFXǕ�7yws����`�ᚮ��]�}�Lz[�4��;~�s�*����p��9�Y[�a>"{��pB�E�G�;w�Ҳq��S��_.���B�TT~7&�|�O]o(�tFw��N��`P��n��R�����M���we���V���֕�wE_]�YܰB;�ˑ1f5�v��K�%oS�Y���u��e �I]�M	�u):�c�R��+��&�O��i"��f�s8-�U��d��)��f���+�i7��ܴ��:����5(9��f�|q\Ը��әCb�U�S=]}a�M ��g^�>��`��Vi��'X7*'\��$S1Sz�,޹̷I���la�f:�f>���k�*W�I�wݼ��Z�;Ζ��.�g݆L�s�[@�j�3��Ӕ����[�H�8k%�傞�V�#��A|�uǼ��Ua�_G:<��H����E�u�vi[����{at��� UK;�H;�C��)���8Y[�m6�\jV�o9�_b�[�jv�ߪ����
64h(��(̙!�E�,�M�B D)F�QbJĒ�I!!"�b2�e6J(e�
"(�h��QAi������j3-�a�Rb��*���(ؚQFIѢ��&*,F���J �1�AQ��#F��&i2cl�43L	��	�E���#&���E�,I� B6,D�4QIBHDș�QF("6�0����0�A��ĖK%&�cZ��g؆�ޓn��(J\�D�b�B��F2�QU���Ǥ�[�;�[x;sU_R1��&��219"�n��)���Uə�}_}_}T��\����C������+ޙ��y`Z`�+u�\#��"=���EN�RKt��C��ד�7�;�)�b<�S*\�x�Ǵ�j�Ӱ����QZ�=u�5Y��=�I�/f���.�@�Q�TQ�Շ�Ƌq�H=�S����РX(�:I�u�x�-��'v�D\�ξhQ���3�<6�O�<>��Y���C��es��یΩ�I�E[Y����8Q�Բ��"4	@��P��;"c�y��zW�+�W�i�� +~�����﯑ɓǃ\����Ǭ��Ft�C��t���:����f%���nD�:��Y��Y��S��r���B}�.����;�LO�*�7o�x��u�M����_����_��;a�9j� E�q�En�P.N}2BWt�������u��V���;5z�L�pĿz�;Z�����nt���9(7LR�f���u{��+nW��������Ú���~�����p��_ZL��c�F}�^��)�&�=�zS]�or*�K���"��E���P-��'y&{�q�v�8�r��,��e����֋4���1�>��xH|����J�V�ɬ��,Ǽ�����WF�a�Lp�W
H�)^��.��m󜂼ޫ"�
�������r�����}_}_}_>�`L�����?��m��"�9{
���<jw�ޯ>�[�ϗM�Sz�v*L�~���e���Ok�wΗ������x������cᇪt�:]gϳ]E��5K�v��4�ih�ʴ�p��r���|��0e��l�r�]���#�^���W��!��5x�G���C�U�v��7��ۤ�����R+�X�碄��=����y��{�LۅP��g�����}�=�q����uzm��K�UI���^=�?Vz6}ϵ{�E��ͳ�U��	tu�7�U%����e?6lR����M=���]���0�O�����}MŞ5��`zq� ��no���~~�r�lG=�"k�+a�ye��5������,��,��`n�*�8�6�L����H��P�GQ������1Ƕ�~����7�|�P�{*&0��P��^��������V��K��_i�pni��˴�ծz��rٶ�5��TvRɛ��/u5p�<��� s�������T�sh�ז�ԙd�ßv��Z��'
��w]#��`�}l�j�jKC[˩�Ƨ^)}����x�#�R~�����^�7=�_%�Y��zeB��#����Ϫ!�)�Bߖ�C��l��}���pʞҸo�[�qጪI�pϱ�|x6�0�f����O��,<�ٗ�hn�S٨����1:Y�Ԗ�P�����øF�dޡ5�lk̐��L�2S(=�ے��K�M{VTf���9&y����\��"�թA*o�f�{����}�z#�wzӻ�q�^_�R�S*F��syU�T��F�����}OG���6~��{ʢ%��+�O�.ʸk״v)Im��w�=S��y���}���v���e�gҒ蘨��g�X���S~�E��Z��%��a�����e������V�.��nG�z3ڍ��t�q��VBz�^��=d����U�)'��2Ó�N��{�������V��ʰ��{�uzR�z����]۟4A�����+%T�F���Y��6��w�ΛOc#� �0wK_}�z�F��MF(	6��wpt�>n&Y����/v��{�SG
���M��S�'uԜu7���;�qo���g��W6S��t[2޺�ڛ�w]a�-v�V�w`�	�k����W�_}�Z��+��ź����<��#�r�>���:�43���¤^y�)쇙�^f�����շ��W�	��qZ�� ���ҽsl)Z�b���=�.j��Nkٺb�Ov��ͧ��ڬe������54�Ѧ�*�m�mA�i�_e��/t��4���5�8�t#��=7�]I[�^��j^�C�׭ʑ�n��y[O%��y�y8�W���C�S��{"���]�ζ#�:��b(K�OI���F�{=%q}�~J����Sqػ��O�v}�9L��C�����f��DJƌ��t{��	��Afח/v��u��)���a\L7L�ȳ�-�ʘ+=�Y�f��$�wn���I����>f�R_�&�����LCb�ci�VTsg��AʱؿRgΔ]V����/ٙ��STiy��c�F}_="u��|���47��X:��x�v�9cj��Q�u2���/C㍇lkӦ�彔�7f0zӮݾ��/����jKq�b\| �k�'5�i��X�l:!�wX`�|�sxJˮ��;��8LKq�9��𘃎�ŉa�|;�l��
1�������=����ꪮ.�^�ONpL���-��Z��w��~�f���?x:�Y'�X���s��W��e�U��қ��k<�mRS���5AK��5��q�,�yrr�5ߧu��\���~���閗n[���S�)O�ޯR�N*S�xR]C���H���~six�f�ZZ8�_�n[�^�k��>���͟+���̍6U���Z��&��{��/s�~�r_i���s�/��;��4������qz����^�{eP���Ɵ��j����O}8��g�Q�#{���׳w5�1b�
�J}�gu6��=�Z��O,�j��*��e�L{H������n<���ܨ��D���*4�<������ڽ���( �[D�K����ڦ ��CKn"�5+'!J�\%�o��	���ù��i�D���g�*��ALoٳ�`%5ⰳ}��5P����b�bo1�L[|���o�]]z�)9�s(k��XS4��ydyAh0J��j1�aզ�m໠�م_NJ�j�V���u��m�YS�+j쬥�>[ec�Q�Nn�I�4�:��B��C�Śi�ɯ���7�h��2�[�k�꯾��M�2K����G���C{��~g���e ��0�y%c���N��J����.驺wl�I�2�;�?1_6��>E��!m;����O���p�s�˳�/d{���Y��KPʍZ�BoC���
�)S:mL�x
q?\�����b�/R�Zu���_����ZLm�;F}��P!�P�`X��Q��-�?,������^s�/fmy\F�[q��qBw4�5�����ɷ���C=�,��T'k�]�����^����I�����r�s�m{d�̧Jy{<�y�����K~����U��~�V��y��~�Ҙԧ5+�D����;3�~�=�?))x�\l�8���/���6�Ǳ_g���^ь_R�.��zz�݇���Hg�^�i��k�z�և5s{Tҍy�peNNTD�{V�SmueI���^=�?g�~���sZ�V6���!�٫�+��:�2>�k��<ƪ9j3�9�}ٹǝm�ӗ�%-�y2�[�]��S�l.��M��EM@�W��NHp�:�vt[S/��!��P�X�w��@��^`�F�_6W�5�|A8T��NI�Q��">�5��z��f.nW}X�;�:�KډQ���Z�ll<z�ORYS}M#�LC�R%��o���qg�l�r����S/R�3�,o��f��C��򜏒��z;���?v/x�#��!�n�i/��SsB*����4��f�y�UL�[nƷ���P��ԝ7�٪�}�S9mx��Ri�+��Чg{��6�:C����\��^��\/���%�� ͭ�MN��rܓ�/U���=�^n�©&���o��n�>��L�{�sD*����V�}!8�+�5�q+=���f�%��6�;���S~BƄ�D��^m��J�Y�ټ2��p�ß�s�f��=��.�Oh�\^�i�:����V}�����k�V}�f����=��r�D�w�w}�+�
�$�{�<�8�N����uۍ�F��F�p2�ϫ��c��y\�z�P�u`��s&�Ə�ۛ��%����{�4@ë'`'�̼�h6�=䰪�^R�&(��ol7/e)�o��5�:0�	���W[!yzݺ��C��V�[��ȭӍF7݆T���:��Ηͽv�/jM�i��+Y�r5:�GSjm�H�������~����6W�;1�Fz�$^/8R����X���e՟@��l�{���l�'�uJ��w m�<�j��Y=>�vg��j�����]��-by��Tu/w�7�2/�ߟ�+k�k�}Ko��G���r�����v��҉K*�Iy�v٪N+%�Û��:�(�9V������^ƺ���.:��+�J2oiҽX���|��$�rm9a�A��!���7�Ž>�c�s���_�*�^�y�>^�{�zV˹��*��r���Uvݬ����Yf����n���.<�o�~x����-�������� ��I\���%/:��7�$��Z��)O��A����|ܷ�,��+��v�N��fP��w�s��m}%z�z�9��<߫��7�Ѯ�'�}�P)J��G�u�������c�n٢@K��,��b��-+���ܪ�
�`'YW"�xL�1�⤞Ӗ�U�F(�;�!�z�{S�7S�+�y��_WV6�թ+���;wkݷ�H��5Yu�f<n>����˗>�$�bh��;Oq��Y���OES�ꘗv�D�`N�h��d�S9]�r���꯫��]C<|��6�=�}R��B����#5앎��-yh]g�Sj%����>�ݛ�Bu�ߗ���z�if4���ʘ+ԭ��՜��]%�e��k8���Oh�kL;eǚl\N�9g�;"��ɝ��;w���ϕ���y�����^p�����qo��y���;�U�ę��|V�}|Y^�D�<��YQ��+I��,p��8ً�e�'^A�9��!��2����>�+yV}6�/n-�9Zߒ�ֶu��sާ��p���/�ԮRZ�A��k������io��ϭ.�8��~��Jue#��d%�:*�MU�_�n�Q����~~q�~��WX�g��(���������ۣi��ӿN��3y��a��B��ly�j�=>�K���ܚ8�X}�E������H�r�{��nz�:��k=Z�ʋ~�����+�I�����4�!G�-�{z��逹[ګ�Gϧf��u��e\{��R[b�J��h_�!V�v_�'��5�z�՗�|���NιXMM���U�N�"�;3h3�r�cZVs����h���?��<�G���1�ޘg=��k�Gw�
��}n��c���@9�'v�F��)J�7oV����Zx�٠�H��i��W{V�Q�Lf��[*����7]IJ��/U�%F�byoCY<�mfuF%K�m<2�O���c~�����ﳺ�Q��+�۔�y��O�m��Ke��ߩ��l�qgZqw�R�\�������>s>�}՗<����3P��l�MѮ?bd�g�VOR�{��~k��x������*�sWַF��}���,Ͷ���I4�/C����6�]�����z��4ԩ��/n�Y���)):�}�kP��V�P��ḷ���t�X�����T���)����e���}-�kڳu��j�E����q�;~��COy�#u����X|]�r�^{~>܉nr�m%�i�\g{dڙ��'��ٙRx_��q���[��-��7i�j�N�B�R�ۥ�-�/}��(���tb�.���7�t��Z�Z���m̮��u�Mq[,i�iN�Q�yj�ؾ��2��]k��C�'w}B�(����q����`���\�G���[����:�p�<���JT��bm)os�'ڍKH�,�0ƞ(���θ�*[��&/�S��b��q��ϯ!g=�hXt�o�j�K����˄���32��]�T�
T��u"�:�@�;(NX>[q�͒)���}۬�4�]-�2��\/��k������D}�_N6���6��W"d�ư�iԱ�[>5o4���N�Д�h��J�EWa��*�'���`��I�4#v^�M��ڋwK:�:;�Ac�շo���f�.4�5`�L�w��R�r
J9]��7�1���`�Pg���ek��.����3�8;>�����I��M����\S@ٜ��yv-ŭݼ�!��6���f�3��Vq���:�a�a`z���ѱ���p�e��At��S��hkRU��,�$�E�̃/�(�@U�)�hM�W��eL���ʏ;%�Z �D�oE�&�gV�Of�B��p�|T�؁pmf�������Z���ׁ&�t�>��t�����QJ��nipٺ���p}sl���(�d]�y�T�.�>�5�E�-�3�-�Z��:�ww+`ں��@v�����Y,caf���}��X��j��0S��5���t��]�ɍ�M!��o{+/J�g'S�P�&�wX�`��U]>vۖ+2��V�⾺����!�\E�vS+$�h���Qs8t�҆�Uv���n�Ƌ♫�c�l����u�Z��#�کrcQ�5a��ΡEi�˙�q��z"Q_.B���{A�ڟa܎vc��cT�ÝX��(����r�G{>����31@
�����\Kl�hn�e�-�Z�
T�RN NP,>ȳ����8c��gH��勂��W\�Tҗ�4�_K
�ЬR���wY}MN�r��r�`���n�ű�
�E`�u���}����Љ�-�t��-t��z���w�R/5_
͌X���k��������n��V ��K�b�r�=|�]\]x�\�M3+��*hQ�%q:o:�L
�=O:'�-Wl��v��H�O~��ѹ��E����+���u�Ū�'�w˝�7:��WZ:��Μ��|��n�*f���WV�r�sT�*�.˵�
۷��S�gx�����8X�Drj�G�6����`����e��+{���5�[l�{β����Wc�CχU>��fՠ.Q��dP�]۠ �f=$�o���v㭚��6ݧS��8����Ҕ��=��+�oj�2ɴ�����i�wu��:�W��"$\*5b���b��4�2'6���}s:�*��0�#�n�M��D¾�Y **�������b/��6�bף7��ܭNc�w���|hӀ��hW1o.��^7F^
��s�X�b^C4Ԯ�0�2�w�ۆgF��mN�ѷ�K2�bB�M�4�Dj1�bب�lR�����*6Mh���Y�(���hֈ��(Ѣ1��IQ�4c`4Q�&ō�!%A�2�i5I��k4Z65�!��"Vj(�""���I�h�hѣHm�����ѱ�1����#h(,U"ѣb��b��F�M���Y$�h�5�d*��(
����٪�����Ї���ָsV_��Q�v��x��8a�̭ß��(��]�@��}�xd�UD�9c ��.�٫�ﾪ;/і/��F9��t?y����x2��}�/֖�L��p�½/{��G�7�]�D��g�u#��vy��{�ܪ{d4����r��q-�~�f��OW�y����dξ��-t��k՟E��OOQ�<�wzCS�/r�V�z�Ʀ���K-���C)�)���P�-�h�խϝ��"^���+��ZE:OjE�{��$����w0v��*�/k�Q����بx�z^��n���r�M���W��ױNp�J�w-�ߧ�N�37���������[�SRѬ��!�\<+���S���R��7D�i{�Y��f��x�7ujA�3��������~k�b�q��>�鸠��݈+��ہ�m|���چ7S���1�Y(�݄|�=��~f��)�GL�}BSU�i�x�n�{��Xb�+��e�I4��c~<)��O�;W6(C'(z0�B��-㋺���Iw3mޔ&���\u/��-4�\˘1�Wwyu��]�W�}S;��+j﮺��	S:�A�(\
�W�%c�Φ�|Ej�l�c@��-
;��T�$�Ȇk�Si�w}1L�Ki�h�6���C�r��n~����k�Ӱ�)*�:܅h7�������h�%���;=�JR�c/|�&��]Ӄ��Ok��vy]/m�{ٚ�����-R��ڧ����N���_ɸ�#藢�e�Pw%o�r���wn�w���Q��~���5���E8F�p2�\���8�ȵ�����G��z)PK�N�rm/8�<��U��){p���>���{��('�9��O03F852P�{��<[�'�u������{���k��[�x�z�y���X驝L��'�h���ZZ<r��Ërz��V�7�^�AS�/�/�Ty��j�B�9������[��]��V���V��=�k:�(����CQ���u��5��/����D7���N�Xݢ�~�qTI{R�k�}[k~Ǐm«��r��@�b��k��{r���^�ץ�h?��i�u�����UbJ���p�H���۷�H�]ٔe�|)���};[>|���S�LPyy
|��X�:�4[Ҏ��٘V�!{#� Ea�t���l���h�{�#�F)X�G���YY��X]$\�vͼt:��{��v-�����R���F�]�`	w��J]ޔ�7뇁�6�\)��eR����<��:?o�FI����ۃ�Ƹ����#��k/�T|����`5;�<�d6��l�mf���_��)��%[q+6^NB�%q�S�I�d=Uo7sْ�dќχ�����Q�)߳d�!,��/n�1Z���5�+#;ί��.�~��8�"o�Ox*��L�ȅ;!o��f�V?\ijn^��J^��z�]�[Ǘ�\Fy�l���
U�����v��Q��ה�Vr�h�~�
Q���-��K���bE��sZa��ˏ;�Cb���ʈe�2�n_�)(ݏB��ß#��5.{Ny�����
v>m�;F}OG������+��}�Y�x������Z��G��%�Y���7�i��m�p��3��e{(�.r�͍hk����d'��zR\��mVr��Ome����'�Þ+H�cF�7��@O<\pU٩z���Xjr5����ܼ��Ct�N�=+��T�������;�T�R'��ڶT%h������������6zc��SrC0l��E�䖻�v��ڜ�wn�1��]��]�wN�tmC��n���wV�;�Mrھ�fʋ�pf����������ڡ�eU�ΔV�o�w�V�8y�U6�QY�uD��z���5���퐿9��V>6H�����e;���S��D�\��e�7&��{ͯ5��cv�*��G��=����n"�$׾ǋ~·�=+lyDﱧ�v�����ϓY:�eW�8�v9�{��]���m���b�U�)_��x��x^�{"����Cm�uX�*fN	ﭡ��w-��~���*��JRr!byoCY�1�~�ǲ���k����/
)�{�j���N���t�ܩN�,���۫�Zfak�h�ku?f5���~g�.��AN��&	}�����6V,�6U{|�����ږ����'�*!��T�f�
~ߖ��|fz'/��ᮯ��ܹ��ٽªi[/C�ld6��l�"��G��6�̈�8�7[�[��W�<u`2��Ѫ��v;�!7q�/j�������<�M�	G\�m��;��(�� z���Tq4�u�\u�����Y�P��(��m�l ���\]W�(�xC�v �n&�oY����k�U���r�_Y�&Z�Jr�Ȧ�yC�{P=��h��j"Vzk؝B�=_j�k�އa��F�����'�&uH�3<�U��T
�p�5���,S��O?�hߏw�e�����ho��ԫ�%M���~�t�ݪ��o�D�9{7�뚺+�X�,>�~GY��[���r�z�:��mzZ��r�E��۞Hr��T�k�]�����Rw�i�v=��q����\�{H:���J�M�9�|��`.�뤺��ݛ�oG;>��#�����r��������r��ߏSحS���{���e�G�d�ͫ^���^�'���݇���I<��=�wuoo7Ƣ��N�G"4���c�7�N�����5sPV=U�p�׮)�Z����o��/sɒ�?�L���pzmgT����^�vVj<��U�9�ǣgz��^^�g���b��,��e��oٞ��>�)�t2����&j�
]�q�Qg]N�� :���@�#X�\�/��Յ.*u�msy����6�s;�C2��Qus��O���+�YVz�<���ek#�wuvdk��p�n�`��@a,�]���h-�|�4ksWs*N��S�g%޳���{ع�᤾嚳�{����/;~���S��e�K@Rr�~��	F#��Ǔ��0�[�m�I��JiJ~�|��S�)�P.�{����p"v�J���2��Jټ�c�{!�7���y1�Q��u�E>�G{^^ٝ�q����]"� �;d)�KlŅ_o��~	`���d���I|ϱ�G�災w죦�5��g3���<C`��{!Z�<|�uF��{������x�,{�4>"2sE1��Ш�Cv�}
��Ҷ���X��/m�W���$��#2�ڷ�.k�ŗ�yѨ֘5��v��a��G=�״��Ȳ��/sl��8�Q&p�&�y�*�N���6�eF��C��'فk4�d�M@~�躖�yn�웤�r-�k�?)�Z{�y��v{�}���w�qA+��]�!4�A�V!B���{�g��Jma�߳�֩�ֶz�y[����53jK]�&��R�r�N��{�ݣr�|9E��x
��)VTr
S�����*�M=-�k�t�P�g��/d��5��³Y�x����35�m�D�2T�|i���B6�.��gb���[�%����Bґ��s�iT-:8�cu}���.�\Wl�=Q���V��5�ʰ�߲z�.���잮����ns�K,�ַ@�j�O}]��J^+�V���V߳ض���j�T���'��6�ϡ�V���I��^�[x��d��=��:G��P[rt�=�j�<���sq�@�c�
�X������)�]�y�q�=&�gz���d�E5����D��p�v��ov���i�7:[#�Zhl�����f��Z��	B�eD�u'u�W8�?_�����?i�F� ���H������,����`��O���Vf�ɨR�n��!C�&��Mt�R��n�����'�r�~�_
�w;7ބ�|�o���*L���叨M�u[Qw�����ʗL�"��[P(Uf�S�vz��ۧ�E��>�1O)[�y����j�z���pܲ�;U�v��������q,b����<U�k�	����KW#�;Y ə����̨�bNr���7��j�au�/z*R��i9�h\7��Uɜ{����b��J���7.�kj��uuq���+Z�(e���4`�b{�]ݿI�וyl�nm�\��Dw Q����.Ȫ\D��׵�ċ����kL;��v��k���9v+WS��>�]��z5�or�s���N�=噯�a5F��)mǞ�#>	ŭ
\��g�[�6���D�nQ�}h��߳��o����w����a�ծ�x ��I^���u�}M�{����g�~��p�nr��Ok[;� g��l�srOA��=�~���>+����7�O?o�T|{�H&�<���Q
����I~kh�[^��������o��?9�R�X��*�r�9,n���׳��ל,�y�.rT(���EA׭�:M\D��o۱�v�*��VS%j��C��)�S�Y���8p�y�@�����i��i���~+�tm�e�a���W�j1F�O����]DI{Q*5y�cv�5j<��)M�;zfV�5���nc��j�g�����>z�$�C՟RZ9��LO7e�#Pu���f(&C"3��e��2�����w�Z9��U02�����Y��\Y̺zt�[f�5	:{ڬZW�5w�p_9�»j����y|�K��_�7x��KU�q�΅od�ɋ���������Y�ܘ�ᥦT�yѭ�y�"͘ե.T�>�)^{\�?�Kdv�Ӳ��\�^�ܦ��Qfg����s���LW�q��Z���o�Ƕ���K���AO��l��GuN�&<F�&N׬��&�q�'�s�V�;��I������?3�L�!o�q����4���S��gm/UZ雓�F�=��*�i[/C����6��v�ǂ�?rr߫�=Q��|I�̌�T0=�Eeϣؚ�/>լ�ɽ�q�*4�Gg���X����֕x�׳xM��p�k7;�����ǽ�+�@���ayl9^��qK�S����Z��s*�=����D�/c�.*��IuN"qy�{o������5��+�n|�Y�D?\�҉��y I�?^�i�ğV�Yq�'Y광y�c�9g/��ʦ������N�B�g^�]}�����K�-ҝX���P���/N�퐿9��V'�A����?dﯦ��6cb%\Q.���Ƴ'���"�+��/<�{`b<�>�Q꿬.�0��u.U����s'��a����'tְ�J��s�u������`$��p���2b�J�����n��&����yɳ��ΚP��Ϣ&^�`�֯{�������L[Y޹���.��P���]������<��M��NI���>�����6�T<pڗ;R��8��n�npE�V4�/�rn�*��C�I^�͞���y˹���q%�J�U�-]�[G}���	]���/�Uȏ�އ=�f����Y�e���}~�.K���:�N�.l3ل��su�[��oێ���ޯ?����+!h
`�?V>�k3�����w����û]#����B��p�5��{k��>���⃳U�kT/��^ٛ���s�ۃ�BQ?Od��ȼ�k��?p^�Uw����Z=�؊����ރr1な�+e�0�{"	`��݅�{�RM&/�]m�>��ߠ�<��6��*�ǆ�\/������L��j��:��o�j��q��;��F��{Pp퇨�Kv}�m@ۘ���{y�ޙm66\T5ra8��
���-���M�4I��MM:�`�aJᏏ
�t�n��:F�L��.�҆R��6\=�]2��5>��Zrԍ5�b�W�1��E�8JU�4R�3�-S��e�6�
����n*$x�Y���+(!Gt�%�s����ẻ�#�.}�^��mH�̧�ս[�d���o�?U�P:�A��n]s�p_tW;��q=A���o7t�E��.��0U�vӣ���]����X�O�T��vPW�J�8�Ѻ�	Gn�6�v�Ҍ=ք|0P�tn�_]�J��׎&�Jv��Ӯ�����fe�9&\�CΙ�8ͺ�w�n���*=wF��c�E��+�8շT����h��c���L�o��_J��X*'�I�I�[�Zy���0��y��Yz�T�rce�7��GP5�S<��ڊ��C�|��.�;{��k=2���]+�l��[�M\&�B�խsH��2�v&;�ࣳd]F$�׈\�w$|E����c\��eWhx�ѽNq M��%���/�fͣ�p�i���[�U�ܾ�y-����t^�՘5�$�N!��\�:x���t����㙇ֶ�U�5��4&a㭺��g	E�@��oiV��àdX�Tu�/��2#jP֎c��}�<�z]��q�i��/�ٵB!2muK�D���ƴ�~�{-^�¬c�9A�.Ll�ճfM�R�*
/��o��U�N����z�lJu�7���5l�J��m�N����qnueA�Bz;WD��
�I�D�Tݾ̘[�.��D�8ٽ�ǰ���v����S��{������o렰T.�S�lv�[�Ծ�u&�*�:`�}��^Jf�d�5�Á�l^�U3}1v#@u�euv{$�E6vζ���7�joZ�B���.1�\N�5�خ�j�Ƈu�T��0��l�����VRRpO,͵���j��-dŪ�A���|����63�9��Ϋ�T��S9a[ݖ�}�cd�]KRR�U���I���ʇ{zŴ!F�ms��0�����辙����Y����g�"�{)�K�X0[U�"��̠�|sR�bڜ��W��b�d��E�қ�y�c�ST�:�}!7B�!|������MҴ'X�L����'A��ݼ�E����-���m���nia�Ä�Cr����ʲ��=j�w�ZWGI˷��n� �)e,wn��/��7�k�Z�֮ܺ���X��j���j�y��p��H�����|�F��Ӭͩǡ�J�� P���zE��{��&Mі�@ф��w�H*V�؈�jqQ�.�ڱ�v�9���K@/��Sr�^���TL��݇�W_Uˮ���Nd &p��+twL�j��i�T��n�w��3�[�fT�L�O���.cor�|��v���bN���0��M��[��-�ugwv��b���w���
T I�m��V�-�Ƃ"�cQPF4b,TI�I�Q�lm��6*��X5�M�ƌF��[����F��Q����5��(��$��TkF4b�X��-d�cZ4[A���%�d�5bclZ"�TlP�h�h�IlQ���T[���c�cX���Փ��D�b1�jű�gg]������+��$쒈x�/��y�slKw�$���G�2�S�:��Iع����q���[��r�R�U�2�s�0ξ�>��S�_�ˤ��CI���4.�q��]�^c�}��-�`�����zn�N?M{�+6��9;�#_6�eF��="q���-ތn��	o+޺s��_��{9-���i>{Mi���>���o�[�~��`��o��OW�_r6�^���`��=�Q6��W��ڝ}��vT���ž�R������ީ]��޽�I�i¢�����Xqmd�͵����s�P��oV�}�wz������3�m/������mg��I��)���OX���[��V�l9OK�y����N�U�4qʰ�z�i�>�e�W���U��N��r���<����Zi�z��{i5��]�s7o�����g�/XopI�f=w
�hy��7k��}��ޢJ�����Fr!�z�	����W'���_I�j��)�з��ax�ٞN�W�Ӎmwk6h��x!�]������J4����|��";�*�\;�۵�
�f�d�����2���;v�\�	�S�+������S�^���q��sV�^�g���R�rw��sD;�q�V�h(ŀ�k���¶�7�Y�װO)�������_ueU��`����y��$���Z�'֎�y��!�ާԞ�����f��9��]�����s=H�=XO�n���ay=�Շ�k����}�K�k�D)����@�{9��OIZ�ږ���uyiVf���Q�+䵫�^�a��q-�4�9��g%Y�����)�y��Nʉ�鯽��bE�'�kZa�.<�!D�Y��֧�="�Qyޭ>��X�����z�M_�Vk����)�m�<�d�m�͉��y�2ۯM���'و�h��+9y����j�]�ٿs�v��3�{��E��V���ZUDc0-�Z]���j����)��Ά���E�j��yM���Y�6�c�9g/���w[>�\=�?�U�0��C�Z����(��ꇼ9Y��ueR>�|;�+�ˢ���CO�o��c<�-�q�}<�/�^�e����y��ώ1�&�ξ�#p*��G�!�9Mj��þ��:��FV����g}�{��hb�{v�ؖדv�$�^)��]H�<�65���C_7Ο:�
�L�VB�W����pP��s������No1���b��a���#%ˮo��}��|<�~�-�׭�:M_���U�9��� �R����Cu��տ3�1 �Q;;R�mKہ��Ɵ���J^�e�.��(]ӵO����W'��7'g@�+dU���*5W�R�cu�K�w-��[��L�z��}■S^S��K@���Q	{�/U�TF,�dQ���yA+S�E#Y��Y��ڱ�oj���]���:r^_���8tb�*�uy1�~0��|w�7���~�~�7���T���Pc�տf��%"4)�'��,���Á���nM��p�l�z��?3�L�"�=!#�x˟h�	Ǌ�V�i����?_�l��T�Jᗡ�������se�uy�&��CvzjK�,��`0V9��g���'P�V�f���t|�w:U�^ue�|���fR�Z
�ڀ^�ۘ���R��ڽ���n����ZZ�xg\T����	Q΁�Ր��wG/Fv���pt]��fVCe�QjC�m����H,��Vgc���]n����k&_|Eo�Dh]��@�ܢjP4�>�W�mdj�\��2n-r��;��^gE{�k�vG��n�3jn��;�%�Uw�OƸb{E��ڝy����mۥ��o���]��Zn{b�RZ���ػ���ޫ{^�-��5��o9V�v��m�,����%}��E˔Ǫ"��g�ݥ/mc�wr�y�[�7�.�%^Æ�*ю�2�k^�p6�-��+[T��OA��f����{d~Qj�l���Tӈ2{��8�MZW�7':Q[���ԫo�:;��q}~h�'^�zϽ쟑��~���Y��F��鸂�6�zt�{��6��nb`��nv��M�㛼�k�՞��s�^�%�c�X}���s�vׇV4J�Wn���l<^��zZ~�>څ��WZ�������;�:[�&߼�^���j�J�������<��O/�>n2��Z/��iU~O���S�3��c���UW���uql��J~�����c�m?i�|�?#�g_3�0a��1�__.�ģ�Nb�c@u���HA��6RЕ�/mXC���t.�}nT�fl�-1��4����0�\�SEuj\J��S�:�o;��B��_I��|�D5��}:0M��V�s @��ǯ��}R�Cnv�u<�بT�VqG�ppaZ��%�Աt�p�����[��}C�=0�<��6����>�w����7��Q��P��=*̌eV�F������Qc�&����^�<H��8�:V7�' �4�c�e�5�;!m} Of�%g�p1?f���w�#z�/W�*��͔ކ�?0����튅L�[�sc�B�hd�>������8ry��<=�饤�MG��C�Q��� R�7m��-z��^~�Ӟ�9<�~K�i�];�7�N���o�G�btc��U����Y��O��/is�֗o��nr�?'ͬ�u]������\�F����c����k{��H>�ֳ�=6��}�����{~kg��;<�#݈5B��w���ٲ/G���{~���ioÍyr�-��k����w=�E'�G˼q���(׳��{�C<���X��(q�mg�
�!P����U?!p�s���J��[, �L�eX�[ԁ4.b��f�-�QŶu�w�s�73wN�p�u�}��ۤ���EbdwJ()�a7�.W]�R����#�L�Γ��o��6���F��(���e�;[E��g�a()�	I:����j�Ln�l9OTD�̸��Uk'n*ě�⶯�u�H}ֻ^I�`Kk:�6#�^ǒ�5�m=���Яq5��Q�;�ˉp-��u6�!�;�3.$������ǚz�7뇁�Ci�J�3
�>��2�:�}�1�]|�'>z�$�Q'u�W(�m��)J��՚�>�h��^�%v�]j�y��=�l��0�U�R���v?���Y�V*#����{XX�5�괺5]Ef�Z��ٛW?����w�s� ���-�g�J�����\��_�V�mKJ�J��6�T�f���Ѽ�hO.�8��{�e8�������q�^Zq-iC/C�l-�[�Pe�}aC��^�/m�fB�;il���T���������H����kL6[�GО���n�A�x�i���ؗ�
��7�ܕ��N�"/�+��暓���ܪ	��J��ߺ����Q�y��.�zEngj�i��nd�1ׅ5������O'-�l��Nv2l�"��.s����"�t++q�h7�:�[g�� F�]9�'u୍�pZ��$k��KA���G�מ�3��$��άv�5�k3��K훼�gD��2�7M��ʷ^�d*���;�Η��˯���6��傳C�{'#�uw-�^NR��L����B��7 [ځ�*��~��xz'I�9�h@/s�>��5�J�}��ykq��圸��W��ϭp����yT��r��8n@���ìd|_{��;[�r��?���<�/{d??9��V3\�*�&����{�(���D�C/(���^��o��:���I�����lzŇp�-[��Vm��}Ƣ��T���P9�yk�T-���<�c}�?C��*���KU�+w�[�o2	;�V��l�z�ځ�t�����|��=�tӤI�'R�e�T]���x��q�=�g��8�����w2��W�ۃ�_�P��l#v�V���K]ص�X�5��)�V[�7Eb�T�ϷF�y���v�����g+v۩N�Sɥ+|�����O����IX��~�7�z�x������Wv���+n��jnVK� ��e��������C�lZ09�K�`#�x��1Jr;h���H���Zx�SҚ��d���m4��ul�ەz'�ڹς9��q��l!uܴ�pn�=�u�J{�1
���yj�[�F['9�#B����]*��-�pL^�l��3�X�xl?3�oŐn�{�l�)��D�n�T�vH�BY5��~�f�
�I�l����z� �2��ϮzɎ+�%U���8eih`%c��Y��'QP�j�l5�@E?�ܻ�8�gP9����f�[>���~��>�mgyfҜ��ҧ�7O׎�V�8�tjްi��7�z=�l�,���Ӿ�^�4����U��s|���E��)���8�p�E�+����x������O��陡?N��W�ý�������g�ե/V8�^r�\y�T7~>��5��q�Mj�����Y���'�X}�/���Q?z޻�������!O��0G�_fE���Ȗ�>�+J�M_��3G�LF�h���qToYڿ��%G��K/�����d�Zn-��,9��ɵ�^�k�9E��	.�'�������(����������9��,��+�#)���*��)zb����2bce�|����v�����zQ��hD-����/\�7br��(lU,v�rd��J���Y�
�z����v���)��wx饦���c�u�Wnܷh2.e��)aO�*�lvb���x��z$���{�n��5�sG���Ni�ޭ���w{w�7W�ޖ�65�k�	������S����鞺�0��
��qz����o镭R�^o�5�xWͧ������/�t�~f�x�A���� ^��������;8w��?tT�Jy@gf�
w���S�V<����޷����7���
��ʷ=0�8���gI\}���N�&�[�ڶϪ��!�2��"��W¼~��I��Sp���8�I�1�\�dM�u[N<|��y�Q�EAw���U�v����)v]��Z�z��yuZ�+q~c��Z�CoC���������{|%�_\<#�Kl�_��(�'�\D��׵�f�����CI�I��h�&���r�;��c�>x��+Uy�;�ILϜao�ҟ���Y�6�9.ӄ[p=��^O�\1w7�,��&Z��4V#97J4_$/%]q��#��7�k���2��e��!�-����{��۴�iթC�]�v��f����odhw:�[����GOJ�J�뾼;�}�)t�x�.�WG�Cə�u:��L���met8dL�ύ$S���]ʲ�y�N�m>c�.�_����Y�~��y���|�=V�����t]z�ݻ�Ci�?8�^}W�tS�Vf?s�_��k�=��w�Oi�|�{Z����Z���SOs|_r��~N>/�h����(#���_�n[���\/*f�^�#��璕�>�4;'��yz*����J�ⱞV��9��/����G�ح�N�c�5:^½��^�k�k������=R�2�U�v�n�$B���R^zs�ͯ}cP��uz+��A`j�������ܡ�IC���j��w���{ƙ����5|wP;�n�^ޕ�&��x��~�>w��KJM1W��~ب�5��'�_�,�Z��~U}%*�N�WY�vw�[�d�������g/*W<�{a�D/i�7M���ڧ�9�_4�~k��?���6z��^��cގ%ꉭ�o|�_�[c�eO�
w��0�K���V{��]�����N��LN[�(�S�\˴gm��B�v���1ѫ�]@h�4�s8��#�Zݏ��X.k{�:�Y�{/o�����"u�OFd<X�C
�����%jg��;b<[�,NO���L���c�Ѩ�_!�\2]���8�g��˛}�'V�Tmn�4�磚*۹1y]}]o��|�딈�j����Q��ÆP/�Z�����Z�XP7��
��^��,��o{���4����]#���6N��+]���@�V:�,f��D[�F]�듹
��f�*���'�u��)��^w�����t��6u�"�f�d��ԍ�a{TA��ʹSU{WY(s{L��w줛wX��#�ŭ�Z�� <��[����.�+4��]�!��	T���9J�J����]����|�J��wǡ��½/�T��
�E���v�aK�&5J���u�9#�#�K�~���jM�����R΂m[�3��Q}{�����c���[3�� ws�s��v��g=[z"R���a���ө�6����D�[�N5��/f�Ȗ�rK��k2��`%��>����i�=��9���x_Wn�e��R�VtʂˣAj1��)>���1�W��љ�l43�T�K��h�(��Zʓl��`Yu�h��e<y��<��Ť�bf&q�:L�v�ռ�l���VCXM��ѷ���H[���Tl��W���q����O�ת 
؂8﬚[�/kn�b��tǽ|�>���)�HQT5��c�:W�a�Ǖ�R3|F����[��eI�z�Y
�Ֆ�6 �6�֫��ݜ?�ԕM��]y7��ᛘ�j)��侱���zu��l;U����v��ˬ�8�if�t���m�r��n
�N��ʯ�J%wͫ5����Z�xݫ⡫^�
�G�e��y[�W�oCק
��t#S��Z��=�;��X��|��)�c���hZa�8���6�]ə��w՝�:��-�"r�%R:�a��q��72w)���Sܩ�gL��j��M1�S�+�N�L���[�z;��S-���u��.cw��i�ޥ��|ݍ��]��,G5���Rr�^hu�j�Q\W[��-����=�8���Vev�L�ؗ-��vZ�A�F�x�����C�0�4���K(p�AV��o�9띍w_@^�e�M�1��Xѳ"Sx3����՝���C����	|8�uʸm# b�|�_lu�wo4,�¦��~�f9�EO��I�deA�������%LM�w�Bu��ʺ\Ħ{�u�a� �r�<�:D1�[l7m7�w��G�gHw����V滀%;>;+R�DƇR�b��\7�i�{�(�C�Y2 ���mu��+4ջ�)��Y���r�ӬFYLY���Ⱦ�7�w�94H���g��l�5����DZ���5�m����6��\�wK���.�3pu���V�+Yy�.+y�V2	;S���d�o�^t�J�;;����	�ﾷ��U�ŦTb��ڀɶ-���Ʊh�5�@Q�cc&"6$i"�Qh�6ŴX�
*4[����$�lh�Ѡ6�F��%��"�F�5cX��
)(�Ʊb�5��Rj4�Dl%��jMQ��Z"�Xѐ�5F��h��I�J���Z5ѬccQ��]}����=�������v%$��GF��q��NxH�����9���.��s\"'0�r{�V;��u��a�)�k�/��Wr������bߔ���5�}��>ȗL�7�S/���ý;/-z��g�y����Ɣ���,z�e�v�VķL�a��Xv�����v"���>df:��s�Q+}5�N��H��=��0�.<ðu�_cFoE�ޒ�Ҽo�	W��Y��_�����#U��Ess����hU�=vΙʑx�mjN���.�{�?�1oޖ��O\Ϭ�ڴ{k<��/2�7*6��OQ�I��n#;7�<��s�������g-���UF1�-�{�#��8f�~����A��T�d\�9�o��u��VT��n1ߜ��ݞ�o!p��m�+�Ié�f<�eZ�>8|��j���vT��O������q�{���l��Z��V�w�2�Tf�s���}�&7�EA׭�:^㞍��ovΟ��~@�x�}Q��i���>��s���K���-{g�/�m���z�{��v���du�E��(B[��NR���;wE�*>���W����ݲ��bi?(q__����� ��n���Vc�J~�r��������%d��݊{sUҢo��ElB)�rZd�}������� �_Z�.�<)���E�AL],-ݾz����_F�<{��^����P�]�y˹��\D=ȕ�<�(�"��o[�썛Z\�;8k�U�|�ކ���j��V���w0�����[EI�`�5n޺Yn�Z����Gq�k��\y��~՗�7�λ��}��{<p|n8�彻���[��uҥ�P�o�Ʒю=��Ϫ%��A�+]��f��/d�]����<k�(�	㿂�׍����|�=�_C�>[�'���F�s��py�s��y5+�-���*�i_̽�rMy1wq ��`���M�/Eh�ȳ1�-�?�e�uO�3n����R�u����~�����2������*`������3^��|���B��3���O�K��WR���_�'��g��˴�.�\��=��q�|���y��d���@o12=���
a�4rX��t�u
}>۞�\M��X1Hw�S��S�͉�+�̮Ӫ�P�������+�ߺz��|��7x��*c~�hye꺈�?���}D������4��
��iK��]J���w+yN � c���v����m,[�����C��I�\�.��;�Kg5�7Uev����w�u��[R0D���Щ��-�s�n�l\'�ܓ���::m=��D�sx��t����<u/	��#�Hv�U�6!����=��^~O�[u�~� ��MR��ٻ��zg}T�|�y��f����oLT{	js�������r��uנ�WoK8/����M�c2n����7Ǿ[��u��U��]��D1��{.�l��9%�;��+M��7���g�\�[#�2�<�_t�Իm��u�U%d��3�
⺩#uW���Dٗԧ)&*s�r�|=�%Ը�dw���q���b�9��C�jI*�XU����N}�;�ȴ� �)j�:�:)�ޛ��/�i��o��<^>����;Y�G^��L��RAP�`�>�ф����nr��ӂK�2�yt��Պ�{��G������w;��9��Y鄶tedɼ�t]R����J=t��΁0
D���ٺ���Jء��^y<ν�T.�	\Ϡ9����x�\��Е���,��c`In�WPa�K;n*�5�8��9�}\�P1����U~��/�g{:1`KWz}ULVC�.iSD�3[�����Oe������ᬸ��M�Cw�&t5g%�4�K8�����be~�M�ԉ
(u�D���}�����v�=ۘo�5��#�ՐP�U�w��4�]�O�A�5�|t��jk:��v���b���t�Y��t���4W�7�K�#V�cWj�=[\���M��J�OB��4{�sOq��X�w^ zo��9�X�U%��;$LD��+��0=l�Y�����=�P�a��p�
�mWIQ�<���ӜO{�k�wM�#�ID�S^C ���˞��4e�^��@��Д_�{ea���#�����6�z���������G�z�s���K��&��s���TD���,��lfSz��1�O��\y�3wO u�`��}��1_�4�l�^w;�8U^�h���C{����]��u�ʼ�X��c�47Uȩ� %��,q�q��5�ڰ�^��dJ��U˫���\"�����*=��xN�/���<)
��ؖ�:�#�MM�r��R�}�\7����9����s�>k�!��Ƶn���p�깏8��*1�]7��G�g��\
��~�4���uՌ��˄�
�O��T�גp��2ǽvNu�Pkht�nh��o��`ީ�(]9��O �@�K�q�r:��~��q�ﻯY��9��=��}��`{��츨K�xT�v��P��G�g����2��c�����3��O��u!��)����~9 ���Ě.�]�L���i�#4P�RVi�Q�S]��~��]�Kmf���Nʺ�
��k��wHo�o}��fV����isQ��J��ѡ������6[��ŽGe�U�G6�t֚���h��oc�FR3���z�ofnLx�4���G�>�)�*e#2x'��+��z;D�9��t귀�>�<�Z�'��+ݹz�}Ք����u�Iuf6�U��f�e���.)�ߠ�ʢ|��f�ҍ�kL�f��;��;M�v*���wü6}%�C�sQ'@�����WڮB���sf|�����t����ZG��qZrH÷��#/����s �JҪd�C'$g�<3�w�[���.{A�u�����6�?}��1�=�|����q;u�|d\9��L�i+��=#�/	ƶ�����9�9�g��ƮF�j�1���g������춮��R(rmV7�?3���I�2G(;F=/k���k��#[�.+�����z��xWS>����������]@�+���!鸃ި����}E�ʿe��z�/���Q�}�8ܵ�r�oU�r��{ ��}|�W
����k�6>E.�X����-��=���� �P���T�ىV�����л���ޠ:�Ǻ����O�]���Op2p?c)\�q=��H�f�Ӎj��t�s7ۉ�N�U�iL�Z��V�n�j�v
��j�ؒ�Z��]��n[��䵎�G��x�{hڃK�/���c�ե� Hg�D}D�u�]��ed���;�Q�lՇ�q��W\���9-���؟ҵ����!V���R��7�d�n7-\w�%�v��.���Ϊ�;�߯p��o���3����3cL��OW�;RW3���ut@S�}'E9�r�p�^��t���y�Q�V��ר�[��r%���m�z��8N`1��).+�Xo�r+L
X�
�����|_7�L���z99��2-���G�z�S���
�@wX��J�=2�E9��T8/tg֯G�q�۶9o��q��S��s�}H7��C��^Z���^�D�jKF���tg��.eB��W��3[�z2��#���y˳��'��}�p�O����β�~�l�K��(UD΁09T;�N������;�����L~��g��N�M����'���:G��p��5�{�g�Y���uƫ/���bܭ��v��>�3�����t�Ek�h`�{����U�g\N_��l�:}}Ss�wk�|G��S_{�=u�l�pvW)�@,mDyu���Θ��3�R�k�u10/��fG��z��mJ.'OEm�����ơ�� h��������&�-�.!�v��#5��~D�8U�R���:�;�4;W�f��Ď%�0pH&��J'�R�f1XyV�݃�Q.C'>�����f��|��v	F��'���I�V��'���Zz��%�-��aإ'��=�g_o���:*��vچ%mI6�sTW�{��:�S��l�{&hO�%����ދJ_��g��;cN���vג���s����\%{dʾSu��掌���rn!�R�:���f�Gw���7�(Y��l��{X+;O��2<{���W9{Zn������N����'�RoO2d��|�P�R|F)��H���s��Zu��u4�\6�U��S�ล�³'��گ.}U�c讓G�x��r��lϗ�fC���x�}���u}6c���K��]8N_���˿=�7\���Cz}�5�u�UU1�S���))�uՕr�W�x.��۶��ct�T{	hs��*`��+��]z	�"��W��������7�<��f܀�d�^(�����]e�}��S���B� 7){ߗ"ߘD_^��� ڕ�wUp�S�ݔ������~��{��xdK�]��?���R�ޚ�W��yD�{�6�A��W_$�q�Ȏ����\�7}�|��EZ�J��]�\�;��<}�����3�1qNB�s\_��p7�x�/�qޥP��y��4�w�x��ʌ�C5����8�O9up{���MX`�g�F:�pr\�W�̉��ݶ�����[��"��f�2�:��
�����uQO�X�:�C;7d�̃zY��Gu%�lMku�iV������c{%Y���6�%_IڷJ��/��FD�c ���`�����B������Պ�{��G�ގ�3�v���㶎x��wP����6ξ����O���ĝ���l�T�������}x=�s��T�\r|q�U[����
9���p�B���ʞ6Ȁ�1�/��GeqN�
�����e47~y�u�a���N�9�c�e4w;�F�q��#/�튿���$�^x]ψe�zh鬡CV<#$��߬�]�)q�=�q�v�[gǧ4�=���w^q=^�7d������f��pW�.~�~R���R���q_=B�[U�Wt�'�����f�t�����N^�cԪ�=t]�����:�Y�hdWJ�W�*zut���U&;�o�ɿ�O@��5�(��3�NJ%� v\��b��Vc��^S��W�Lm��ǡ>��~}A��OS�+�{�F[�WX����T�[,�C�lNa�WVa�����6��{��a���?�w��yU�K�y��l�k���ul�;��_?e��Dl�9@�r6s*÷���l��g�{�4�0���󼫬X�<�gS��d<�f��'��Ճr3�6ݳ��z�po.֠fr�^� sġЋy���l��tx��.�H�{�����*s�3*����)^L���Lzb�
őf�-S�V�+V�_>�}���KgnA2��������ed�i�9�Nk����6a��ٝ����}�U�wѝ��wz�Nz�8p�g���ߌ��J�%�H������o)c��g�����9.G�WY�������p��f��9���IÖ*�.b3�)���|�6u{�����|����9M����w��\x�����jOߵ�P�W��h
�ѣ���?xQ�����PgK�����;�Ih�\l��C��;`�����3�wSⷡ�Y,/<fn��m��7�7�+8��.{u��eP1���*���H�UO�n�0�{��Mm��[���R��&աc��̒t>�;O�u����K6�$���l	�ʡ�l�T����9tT��t}o��y?UOEtG��������ݴGi��Hˎ��Ϥ�@	���$7P=|��Y<��R<��);^>�#Y�w�qW�iAs�V���0����ˎ��i�9�4��Bca],�j�On��kp�Hq���Vmh~��[f<{6��'�'c��'n+��Ȩ�����D�����|��e��B΁ 8��,�/����j�m�������#�������/s=�2���SwS��(�\�/�>�xs��u�M}ݷW2LMa��G�l�QׄZ�t�[��*nҵǛ����pr�=\�����pu�e���S�z��<9iYq��N�ۼ齜�h���Ny(��;r�@���k�yf���o�;����(�zDhU����F'�+�?S���l��*��"�#�(-����̡���T�^�r8_ϕ܁���p�=qlI՞8�{P�h��e��7w\
�u�d��a,z����.ʃ�\O�r݆�D�q����EfS���eb��x;�W&�����_����ˎC.AG�X��g'��uf�eu���x\ֲ���6{M�^\w��}z��7���롷�����Q���Ԧo��[����p��]aw�J�ˊ��p�d�7�j�g����z3��N���������3��xr<��ضY��W����7�b�L;���f������Q�����t��=��wU���W��o��A���K�L�����g	�:�'�,]zkӐ9X�`TB�hW.��eA���s�ra��_:U}t_�.9f���7�ɍ)��ݑۨF;9�v)�Xʡ��C�"�3�~S�w���[3����5��c������^Z���D�k�-2��Fy^�P��3�uF�-�U߹�T�љU���w��d�yﳮ)�Es��Yh?@��-ϨK[��d8����q�"��W��!�g6�_k����^S���.�-���C��������p�
��������u��.ǂ ��#����$�cZ#Q��6��b�gK���g��Y��o�C�42k���b�l�]��¹�Ux��V��'�kM���n�9�+�׉�̧�Awe�C��ӽ<���Ly��*l
�j���;;V�4$�wkv��N\��/����%�y��lR2�\�fB�]hɈ"�U��i���қ�K�?z0J��Q=vG]�݂�Y3�S�<߳(����q���U��#t#��/nA�&VMZ�'t�#.v٨h�Y3P�ݜ�j|�tu��ķf2��4��2� �����)�߂����]<�9|Dܺ�\'0��
�J�9
w�b�)g�K�κ�TM0�x�<��EǩV,[CV�	-	��[a����}v 
��V�_gaig�:����Ɂ���]R+��-�W�Z�s���V�该�Y�rŝp��0���JY���j�+�S�����N�,&�d���W<�E�{����F
O�4�b�7���ޒxH=�9^5�*yw���[}��u��Trc�G:�͏zA��r��ev񐽲4��)&���#Z��в֮d51�i����K��*c��L�6�7鮞�7��[Ne�<�V;�����J���j<��S�Xz�������m�ZŤ�J�s~��ٗL�NV�ŵ����ձ�XI��03�R��c!x��2��4����5N�
�oe�Jpxm�c-�"M�+�FH�;�;L�w}�����Ctn���nr�_Ko�r�E�N9Fnj�اܛ�Nl��g<�)jgU]�Os.ƴ�
���+%򗪝���{E^:�ki�F�/zoa9��+�9�S�B�.��Ӗm �m�}[2���`A@#��Q9�����|kS���<1T����t�����d���'�e���X[J7��\�p�ģ�G�&�KD�R�
���(}Ϝ��=%ʝ/gWe������̽|1v��1Q��k.�VS��ki+[�w�w�_S�ī ��G!���3���i�,ImonP\�����mS|���z�g1X�[�R)>�9Q*�^d�,ˎ��eN�/Jռ�)�umg5�5v<	�q��O���c����O9�g]��u#w�V���;-��0�)�a�:Te.�N+��׶�v��[C�5��֯�="�<a_�H�s��_u���-X.V��f\/�+h�z1>��_
-�u�yشvt��l��M�݉+WG�4�E]������I,�>�ïigm�Y
0=��KV��ɒ���M̭o�D����+��kN�ïnv������5bᖒ5�n	%�m&$�J����x4W ����T�t*T��U�V��.��3o��N�����)Q9[@��=��I!�זj2��ʔ��Z⨱kEE��Z*��F�Ѫƭ�m5b�cj�F�cZŴmF-�U�_Ubո�W�֋WS��Elm��ƱE�qmƲE��Zƶ�j�V"��ɮKQ�ڍ\mɬm�����Q��ű�\k�*�m��q�X�ο�������;ɡ�b��}1�Ԥ�L�iJ9�+��Ws/���+n�d��i_m�S��4�V�Y��l�+=ꭻ����B��L����O�74'^��>�'��ﳤq��W}�YǣM�d��Q^�����<Ult�p�2��t�PQu/��u��!Ӵ0z޶�oH®#��'2gd�Ip./�罱;K�cz�F�5W�@s �@����5��.�:y��6���6,yY泠˽�uY=��'�;w3%�D@j���v�����-����cWᦶ,C!D���oX��D�88������z&����#$�o�D���2�Wl�Vw{��x&�k3o8W����~=���F_ɫ�7�ԁ�Gë��f�Gw���7�(y*|/WmR���J��=}����w�w�;�(�b�ӫ���ϝܛ�9\L���7��P��G���r�z���7�V����W[5��u�2�����t�U�S�j��~����>��7v��롎p^����Iz�l�u�G���T����Oa�S�'.=��nUXca�������oM�Y����<�����5��}�nދS���]����{��b��Ls�.�~�r�	(���*�
��Lh�b*�Q��}��aΙ��A����DJ�E��TSB���:t:��ܨ�1G٭Rg��!�����&���N
�������9KzR}�6��!C��c�FKKW�����:�ݓL9�5��=�m�ܯK0pZ��EW�$�J��Y5��z�=�;�W.�	om!y�ˡ�����~��f=��?EDY0w�h�7J�K�����37�� *ڢ:%u.#���r���Ayv��s���s�P�]�A��U�J��=����<����Qp9����gH��ǫ#�p��Er���s��~��GZ=�չ~lD;��+��Vv��62�el��9���5��OW}�x�>}=�{�q��5�k��ۇ�`���F)ύa轒
�:���qR���N]��Z����oGS��<v}鍧Qj�[ڰ�_��"p����S5�W�UŲ����:�z[72��C��
�ׂU�=�9�/r����������U��6���7*x�"u���?��qU�a�|=���6Y3ӽc�j�R��讏W?!�=���|��i7��#:����2\� jr	Cs��������wme���rþ���Q��MC�o���Ӛ{���n;����q��2K�KSu�F���:o���­g�W���
�\pg���oP���t��Ȟ>�ӞSq�7��PTu{��asK2ܡ��X��{Je"�k��NX�&]byք+W>	k�Y��'w�>�Z8�a<�8�7F?��'���X�>\����3��T�{sZ*�y��Y�^S띁_�n����YX�>����R�6��Rl�v�1\&E���@<Ek��&�����2F퍫�C+�a��OM����]ɋ��̗ǠgF.p�}Qa�sto�ZT#�/����hB�j�;b�;n����2)�a���coU�.�ߤB�Z!�QNJ����[��g��l�Ԍ��4Y�T�<���'��c;���!����cB]�2�=�.�vϡཻ�+kVJ��Bڦ���3�4:�{�i{f��{�l�{Kb��*=���"�4S�&����g�����q�j��K��'�.����\'s��;�}'�!N�."e��qLt������/uOHΥT���Q�9.G�\�;�gx�j�s+;��/.�F�:}�:3�暾���/{T��h�ڟbb3���C�&X�*N�#���%��@ϒ�\x����\n�Sܯ��Q�a����g�m�}���[t����R����t�u3��!��f�/v���z9\�����sHAR�S�v���Nm_z�ue0׏V#�UqQeUA��hʦ.�R7U<�[�>�μզ�%Cqa�e�R�Y�ǰ��I;���.}(5}R����l	<��Q�ɯ5��\Cz��S	�e#JXTP�ߴ�6�v�����$/xn��Rդt��;�ZW2���W�sB�o{�GM��ad������}ZA����G�h����Y�XlIY�V��lwjV�#�%�wq+{.����xXCF����fkh������Ҏ�a��8�8�T�d<w�^���ˉS��<��9�v���T����Ϥ�r NjN�9��}�}�g��t�U�89L��h-6���[�iϸ�)�;{����������,�����axvzs��W�Lp�Έ�a9@�\P��zifև�u�ف���_�3�OwTNX^K�0
љ2s�2��2;fN��T��7�@+�Жw��
��ې�|�ʏ}�mj~���ݬ�BȬ�n}�d�@ʏ@���M�3�j�\@�����-d�)c������h��W�Cn�s3�MJ���K��<w���*;�K(m��1��=P�c��w�����`�z�����z�]���=�\�� :�����2�SĪ�鿎O��
z
��<��ç�>�U�w���G8��n�i�ܼ�~�o���=����xNou�ۈ�G&n�x\�2J���o�}U.����Џ��Ru=���\or������]�[���\'}�^�W�i���^�w߯ý�8{N����
�d�r}'���b�g�z8z]>�:��Vö�F��ҵg�
������W�cc��������~�/j��P��h�7���z��b�1l�38���T�/����&�����ט�����sV�k6��[�祈jr�\߃������)/_v��8;�� �i��;J���hKLpޭ�خOs����锖{���B��b�Z}�9�ø<�f|TS�9X�`,t���*�a�����%st�荺L��C0���Hg<�F�����?va�L�,���򝽮};��[�5y�'�!��<�]�Y�c����8o����PJ�Q���L8��M]��7~���O\��z���n3��?|7��}�'��Fu��>�u�}��~��b���'�}櫬c��)�����Q�3�1u=K���n�M��}��<^�8��b�{�����LNN�JW��wU��1}�Q�� k�3�HR�����
���;u��Ӵ0{�����oH½���ne��5�'mw�]��h'�B��2H-�(�SP����ç�1���	�y
�\O��k����]-&�y��믮&�fK5���	D�][F����0��/-x�^�ժ�.��HC�3;���O888����{�蛇3�5�-;$LK�� ���o�"c}[u=���<��XUve��i��'��z;��=����C5�+��_�t�g�������["r*����x�D���f`e��o�c�JwVW�z�Y|vN'�;����f⻫�֌p��R�o�
���\7N�]��wV'&$����//��Ѹ�Pʘ���]k���n�NMMv5�x�T�й��ds���ֹ�H�K����v���{�tq�cWm�>uRm��d�wu��j�\r��v�T���~��/���k�3r(���;������W���j��~�>�F=�+��{���>��*�vx�.����8f��d���W2�;��a٪�c�����W�^���AV޹yuNy��P��5�N�g;���b����V����'�����Ls�.Z�y ���Oo���u�y[��rZӵ�z;����갑���H^w��g�����G�C��V�a�P��Us'�p����\�F�+"���qu\3��ztj]�����h�\��2�_��'�:=sz�Oz<�][�r�y�{�z���Qp99.����I��՝���+����u�P���RO��o���!�$�}2��<6�yL]t���-F���������+���;r�f���q7{�e�����Zk��ԐU|g@�ȱ�H]T�s�~ub�������c=��1F��O,.s�� �6^KnSy��7�eC��@�a�'dn���?p�}�]V�|���3���r�=�2jk�X��(�3��a���r��n!6e~�^��:Վw�@��)�A�F�`��d�
ӤfU���b܉ғur�@����y�%��z�|�.��7��S4�b�n6D�s�cn儲��&��y�/pᣨ��1�f�s+7�aW�HN����}S��:3 7 Y�\Uk�n62>��Yטf�ߕtm��qV뗐����C�Ѥ�{��ˎ��*�s%�" jj	}N����+�������01}�	�����;���#����������q�I,�O����:�=�Q��+��]��GK�b�*^����p�
�������D����{��%��å^�u�c��,��h�W9�d�P���\�Ұ��*zoWT��|����}fO{@���Bgs�ί���w�1��t|@�W='b�=��1R�^	��ES�f͙��1A�� n�De���/Uy+�]#�1Ps7��;.�V�C)ч�mS�d�{��Z=d��{/b*�^�t�u��O}�1���c���}��q�ɡՓ��V/���g�6x��Ñ��P�.rS����w%�������#�g��q8n3e�{�����U�O�W��ު�;���ެ��S���ܓ�)\����)����1�����T&+��[����#g'�Tyr��I���
�s+>�˄�Vq}�2��m�/��C��^᫓�_P�Ԓ��+\�t�[�l�hv��r�%�<}�0�,�랮���x�``��cV\ŐZǊP��Շ�2wr�Er���:�k�]�8��)+�Jؓ� F��p;��0�b]S�ſ��de��DT�{��u��W��'��-���U��e�e�)��\�9׶l���p�\x�O��S6�»vT���:�Hǯ�����q�UcK���e��ߣ����"��Z����g��ϳz�oh΍�L�}]Hr��]b1p���E��3�A�L\EL�n�x&˼�8#j벲�M^s;�=n�wh�g;d���lv�|�)��nD�l�a֏l:}I{a��7��x����$��=i���:w�}�O9�v���Hˎ�nK�r NjEwl������o{f�U���U@�s�Q��g�0���.����v��u���V�9�Q]�z\g�٬#n�[_v�E�x���A���@zufև�u�cǳo�Ι�n���z�Ξ~}7&'{����;�X���N�� ^��:V�<:�׾%�,��t�!%l1�K�	(�{VQ��u����|vq��.Gu���3=%CX'l�K��2�ה��c�-�q���,�����ŗ�#Gnu܋�n����3���_w\
S�2alz��Ǻ5�o�S�cP����c�fސfy���bt����S(4�R�d��Ww#�Cz�L��sy�1��U�p�dOR�		V��Wq9� �AJ��>�4�h�D���N�"�����S{o���v4j۶,nX|ٖ�Ќ�\�ЮÉ�1��>:�E�$y���̸�7���y�<����|�`��G!� Ҟ%W��ӵF����lo{*�մ���wi����ܼ�m�V����~���qΎL�Qx�Ԛ:FH.������|x��ہ��\W��]Oa8n#2W��W�=�6>]�[��gUp�,}к�5�]��Z�_�g�9�3���㓗3�(Á�O��S����L
��r�p�D�}��+�S���W>�~��;S��z�	{z���\��s���	��)�x�~h�K�+)��oG����9��w��ט9�O��]!�}ݔ�sʤTY�)Y�~5gj�uR.��95 SQo����V
s�k������Wt��S�]hp�D��-�۠�(��DIh�h�l�M2�m]�4+��{龌�o�B�����~��]��d�yﳮ)�W:�}H46}%�'S^�}b��j��I],Jc}S/�/Ꞥ�74'a���ޑ���t�;}�����=wK<�9�O*x{�>Ǡ ���@����Ծ7�h��N���u=>�����.۠�2���}��l�ZR�\��*��k��6Kㇴ�s {z����J!�&=�-(&n��tu��t��P�=�P�.�v�6]�����s����u�����̓r_ui._w{��;`p8�|r�6/����-[
n=�7o�1[��[M(6wJ��ߥ�壮����ʀ�2L���S^��Yף����jyi��G��k��8������q���믮&ْ�Y@�%um���ٹi���~��(�뷲.���ݻ��MR=H������GwVq=��M����d����*�͇n�@5��w���w�tz(�9W�;��LTbj�J��zW 7��5�+����9��B��%�Qy���[o�GM�*|*uV
����F)zn5v�w�;�>eq2Twu����;�qy.�A�$M۝�4GFM��"����JÂ��p��̧��^\?B}v�z1�WI&5��O7˳6=n�1]p�e����8f��������Ox�(�8N_���ʫk���#��mUu�^�Y�њ�k�Ft��g^�R��\���X÷�ݍ��Q��EL�񱫨/������Qa]�����_���OW^�]]�-t��+{i��e��9�s�g�yT3�3�˭ag�s�v��<�ہ���.WR�=��r��N�P�m��u�U%W��=]��������v�e^��ЧK��ݝ/n��Q���U�At����	ʲ�tȫgɮ���gsCbX�oo�3�r]H�����'ȋ�5�l45�yA::wuJ�2�D�֨Z�w����n�mR�y��3���cR��cĨy�E���}���wI�1���P����������
����-��w����>��P)f�BbQ�Sf0>ާqv��Y �#FW4;k&-l�W�������NG���c����8:Ѫ�hؽ%�S�\ج����-9�6&�wM������A��Wc<{Rc��އ5�w]�vV��A���)X݌�R4���9���[w��zr���2�����:�ř��=�����ÜZ����iif�*��� *�Jϗ
S��Zkb:�Hf�vL[�#�?3RJj���ڮкQ'\�W�k���!(��nL���l|{)���w��٫���b��0fR�V0\���ݟpY��6������YP�@%fU�8��5|�lNj ��:⃉�$���z�(m�

��WaZ��V�=�T�.�Wy��\�Tjr�F�謾фgm9!�����<���.�dX,�8�n�б��&���J��y��WN��Tn� sU���gj�� Gx��ic��*��}��쨧L�W2eɽh�΃Cl%1+��,�OpK�_,9oڌX��\�/c�1듶�w�r�+��V�^P�z4���i����C�;�L�)Y��R��l34B���8z�����:�,�8cF�1p�bl޷"�ƛ��2��QP�՘�#y|��	����E�ջ��f��킵h� 7ݔ�[��WJU����:��J�#Bz�Yu�6�QM��:#��X�2��7�8���j
Mc���8���j�@��KJ�k�.��*�5K.R�TnV)��@D:�<D�b���Cr�hX�֞R�c���h��)[�r�������;�K��u_g[��{M�lA��	�9��Ŋ)�@��%�mV��u�i�d�X!E��K��؇L�I�=�6W[gl�9��o,I��T�[׷/.��tRD�����"�^�����ґ����mm�s�ui��sb
W�w���&��W��y�䵅9>ڼv����Z�"`�Z�p��p��\t;s�����r^�A�vMZ5\�9�k7�hXM]L��٨9O30Aj��h<v�u�+�d^��QGϋ92��Wb�S��ʔyxT�\ڄ���u������{-�xa�eۛ�vl�Ј�v,�2�ȑб	�%Z�Xߞ��s^P�	\���{�Q�r$U�mm��}��Z@�M��'me�^_/w^�|��w^��k�s���J�Tģ����&�$���`�����n��"�n��'#5���&��u�ǭ<h�-$��mN*���} ��f9���� �Y�����բ���>�>�������UEmk��Ʈ+q��n-��\�ƶ�k��W��&�5Wh�ŷ9͋9͢���TUF�Ÿ���qn��n9�Uq���5�9���\-Ƣ�9͠�\qW����mŸ�d����\j�b��[qs5�Tm����DZ�[��EqRmō\\Z�mn1S�5���n6ۊ�lU G�UD|EQ�.Ȳ[5��]�Yu�o��}�AA^����k'NC\n�]��)�qr���$������r�ͱ۵����w��5��uN_ۇ�����j�����rz����I����P�R��1���;T�qg�G��F��r1sޢ�}{$�J�gG\T�)��r��������v����OqSZ����D_��=��Һ�z7: �{�Ұ�*-IT� r,{�H\UO'>��V*���Щ�+;ãM��h��^�~1��7$����v��5�c�}R���$��:�)+��ٿ�e׺\[�X��)��oz��P��s��̬ޡ�_ݔ�����@�T�D��1�$�@]l)K+I�1�,_����{P[����?�֟��y|^W#���Ѥ��H���v�\9��R��9\�����GL�͜���X��qR�ǽ�1�if��m��}zsOq�=���ux�����N�)S�4����_u��+$i#��!W/N�i���z�F�ͫ�7�<���ӜONYَ��X$��N_�Y�~�?f��"WE�Z�!����D��4.�V��Sӫ�G'�2�OlV�Ȟ�R�ү7��d���Q�1�q�ȯ�Q��˓�.a����k/��5�fS�`���W����>p�`�x(]З9Z�ϻ���H���v+�Į�F�g�f��[w��X��ݵB�1V�W3�s�;�i"�x��.��5W�Ft���qr1�tF��%y.��f�|J��Ԅ+{o29�"�PQ=��t��QrӭB�);��"�_<E�]��O����ܿ���f� ���Ea������Tx���a�uf���:�|/{�Mﶵ�E�k<��ݾ.7/�ǡ��G����ʱճݓC~�����r�Fr�\�K��ʿk�욧��$n�a8n1Oq��W���I�.��ѽU�wѝ��}ެ��)o*�TM�j"��[��艟x�����9�Q�>����qމsK��]X���J���J��+�������[=�7�h��#�'�~�%��_���G�[GF:��u�<
�C�2yz.1��V��'ʣ3���1��gĥqX�@3��'�ϩ�e\a��)�D�y������M�{w)� G{�1��:�^.���<}eU�F�2������5�f�u�)�9�6۹�~�~?�/k�#�~���_����美�#������YH?|7��Kq�t��i��8g�%���*2f�ʦ\.�2��,>;�\K�]�G9<�}�Dv��U#/��F���h�i��]w�iE�W���\��t	�7P(l�+�sA�W�qN]$Y>�{��0��u���������2���E3�^w���Mw������{���c��J��Sޗ*�]��L��S=r�+h�7�C�e����'N��aU��v
��.�r��Z���y�t2�½p֩��f^�t8��ҧ*Q��nެ|2�啎0���r�m��W��=���Hnaa���9�7Z�/��/M|�kC��x�l�⚊V��E����m���	�Y���U7v̋�2YRHk�� �SB����Tym�|;M�^�GK��E��7�����>�ӜK����u���3=&�L�Չ�1Q/k���Zɪ�S
ukx���֯m�z���3�:�p���E��\O{���������}
��ۀd=7��mn���ֿh�-�����h��ҙ��z�/��|���CΠwW��C3C.9��SĪ�ܗ��yz�m��<\�t�������}�/N�]Cߛ�}z��7��;���.������w	Mei��;ך�ф�[,��y��{*^��%q��W�D������i�Au�7��(��kF�xO�eg��t����C?�N\�� d�r}'}J����{���(p�YP=7�����Nem�+U�����w��O��s.��	�X��Ma�r%��D?nmo��UM��u�E�J���s���(f��B��#B�KL��;Pݾ8h���ŇX-�g�u]"�Gj�r�uĈB��mX3�۠kN2;u��Mr��Vu��9(���=���A��kc�c��n�$v�)�;��"��*�m��_d��m�P@�u�����V,��4���̼tu_sף�I��jQޛյx<�3U�E9�d��gP��K�k;��?WZ7��п�=��r�4�;�0p���R/�Q���Ο�gj6⌤n����:��oWx�����\>S﫝p�:�A���zx��9��9a4b�$�FN�J���bUqS-�_�=I�?:�W]��oH���:G����Ov"i����b��w�f����,�8 'FtE`�r�I|]9�JUb��8�!؛�Ss�Q��:��s�����a�,�B��2O��@W)�b+�w�!ɬݟe]�r������C��6�k��%Gg\N��������|���@�4I][G��i���fc���y���~ҽ��!o�����D��t��o�� ���z&����B2KFV͕�����1f��^�^�#�[�FB���ۅ���Q����GwR���ކk�Twz��u=�.r.c8+�묑mb�����3=�i�^υlT��q����q�|���y��d�GwP��:zr��)߬�)�����~��gu�\��O����V���¯2��Uꇩ��0K��Qҏ�O<ݱ��Qp:71���������=��nS6��G7cڛ�Iʶqt���X��L���,�J�̹O�h���T�h��*�3�n�mn�WV֞� R^<�ғ"�y�$��\[bv���}E��X$�M�#��uv&ڼ"�I,Nގd#���q�'\�vI�ܕ ��롗��7��%W��\��{�8N\Fe!ٹ�T�Fz����ʧ~"���Ӛ�� �F�5��ޡ�>Κ�;���b��s�G�i��P'0ץ;����k �L���&~{]�q]���Hל��D���|��z^B갸*�����n�~�v+�J?�����ܪ����Y���sN7�j���J�\ �XՐWJ��ᜧ;��K��Yζ�{[�܅��<,��T����I�?R]e�uR�F������c�)'K�Vw���q�ԫ�gC5Y<�ap�&�-�&;�gԼ͙��j��\��ߖ�b�S�S���}�k����㶏���H����t*
ҿ?YΌ��[�=^F���L�-IW�t	�b�U!uS�Ͼ��V)J��N�H��P�}uRѬ��ݎ�3��G��w;��9����m�Iut	�R$T���ճQ�����]LWM�x�D������߅�]׃��k�Y�C
��Bp�WTr����������1���������,��*�N���ұ�El:k���q>�M���#/�트�`�	���ʧ�9���b�җg$u[����]Yb]��q���dց⨫��Be���H��"�Hv� Oi������L�h\�J,Naیr��'�[�e�FX\�xd��v�	ݪV�%�Q�55�X�wc��N-{�y\�����he�������%���ۜ��,R���4�]Li�A��Vh�v�[g����Gz|�u� ��W��hɵ�#g���=�$试Ijo�Dľ�*�����/���
������Ȟ>B2y���~p��^ۛ�o��^���$[��5�!�
�w�	�ib�����#��g��&]M[�Q�h��yI����ɸ}={��dW*> R�rv�\��=f=-e��S��I��]<�7�
w����j�v�ۗxO��/>��o����.�V�C*A��%W��lNa��Z�.�j+�����N�_xl�9�=s�o�6�hܫ��W#��q��V:�}�vՋ���g���l-3ϰ����\��\���=���GO�#�{	�q�_�ܵ|=.���|��oF�W	�go�]w�V\{��љ|ѷ)���v'�G?}�Ò��e�X=����Q��p+˝�z\���uc(���4:+}�3�?~���;�'���\�~W�h����ȗ��	h�T��pJ~C�+9,c�bj2|�9S�ۭ��5s]l�=�I���q����b��{t�����b�,lT�#,�WeǸ��*�,�Ϳ��Y��7��'b��튗��"��tc���C�A��V�0�ø�oe--K���^�-vehֳj��8,���
�*3��*��D���1"вZ�����ѭH���n3����DrUk6E�n�z%��v��w��8W*��d�0�|�͜�u٥���/�:��:X���z+�^�����<}eU�D,U;��ӎ{�+���^MV���UN��_]7��v�������;
�YH?@�T�2�/,�RC�1y��iz�w�F�育�.�������ˉ�N����s�����=�d{{��u�dzL��8U�}��u�����U�)蓠Cs����Td=;�ۊ�N�>�3�V�}#
�wJ��J=x��+EY�F��Z5B���4����7Z����|�K6�7=M�Wzƍ^q^���Q>�Ө���;9�����]�qd�P�Hj�r��9�9��cר��7��h9W~����y{�}��ÇTx�>d�Q�����ID��	�1Q/k����$�s��kpu�h�͚���׭܎�T��s�'��x�*<Gp�A�~Gh�<pZw]��o�ט:wڽ���{O��9W����]�����ɸ��@:��O0d{"9�&�7g�W�U+��B1����������������f�ӹWP����� u��;��m�? s8a[����0Ԍ�Rh�xe&T<���,ѸqwT�OB��VPGsJ�~j�)F<�
b{o\�ohj9nughR���IR=���ܱ�'�ua����A�!�����T1{V�s�dީ���5:';��ڶkl3�JUqo'r����y�����8���x��҆,V�GPQ�v��.6���=�L/)®:��/�����-�bw��^῿~�q�,�ߒ�cF�����9���%�_��7B�Z9��k7�Ї}9M�OW���VެFw��O��s/�3�y2�5���Ը9��wXѪ���N�z$�o�u�=LΤ�Mw�y�&W��p�>��)�{t������0�N�+�<]uEVb�ʺ�M�g�",���/k\�ao�P�����S�և�������0���*���}��NZ��`q�%#Pgj6��7E�L�:��oWx��O����g����.b}�.p1O;"�%^C����xda�/��IU:r�~��nbOJg_�X����O�ޑ����V+/ժ�AWW����X��������&���\T��p�W
�[���'h��A��޶��:���'/��~�ʀ�� t���\��/p�|������Kwq���*x+��u����;c�ӛ|7>}KI���߫��&ْ�|���	G��>���fc+i�.�O�;�{��l��@�IM�z�~����{:+z�V�V���h�Oul�o����:jY[
���f?��������3d����򚹞c��)�WW0d��B��;/f�R.w)�Iӯ2�l�,d������$]�J��n�M?�����0�}徐�|�=H��@����t���z&�s=3��4=�&�zv&��37#�u5�����&T�pϋh�{V�I���@��up{�3^��s���{d{�=�Utl�L�|�Z6T�T��u/�Q�R��j��5U���q2Dw���ɭ�t�Ή���T2�!*E28��+��¯��zoU��}EFCb*�~�9�ݷJ��z����QNMǺz���Tp͛�O����Ů�hYjc���R�>=�EW��ϳ�sު�C�W/Cޑ�.3�����ν/��s��xf\�T'�a�]EV�w���R�V+�Gm�e�ʹ �j�=^�uv��#zhn�y<w��g��9������,��I޳�>h�];_�*#�\J���
XՐWJ��=��:7�m��D?
�l��8�ؙ���Jqrt���U?7����eN@v�>f}�2�8�퉞��κ��B����[EZ�J��|&t;��yL\S����渿F��;�����a`9^�̊ q7��n�Q����*�>y��^�J���nL�r�Bİ�XN;�����v02 ?`���77�gQ]\A�F�5���u%4Jf�p��҂{h��tƝ�/->���v�I؊�m������f요�/$��6%>Ɲ�U���*6w��� LN����������L�$�g@�y.*U!2y9λ��<���������x'���oGS�'�w*��k8�z���e]D� $Hx��5S���e�`�U�c�Ǫg�;���([�׃�O3�z��(O���}qވ�,	��f�q��;*|UbW��qOF@㪀���Lv��Y�qW󦼀~�G�Ѥ߻����b�cv����詋|������%���c�1̎������*������=�"e`>�l	$�znt+�s����;^�7
d��?�� k�(W�^�����	����}&{j*���z�h���Oj&�D�D���]��$\;��Jd��M�񠾮���1S�&p�.HQ��O�߫���/zF�۝w&>�%C��ކj2+�T|@�r��Q���񊖲�nǢ�R!Fˬ��QwI٦�=��n5����O��y�2���:��|yL��x�0���e���������}[K��=��6�h������}��q��[=�F�;��{{8�x���e�FU8(���vm9'���n_��!�b5��B��j����Ir���]�zlh���q���@�۫]�66eX���r=�&�B�R�2���R:CEҲ�˛�k_N�Q��f�DK���eޔ�W�������2�r�B�W$U[��"�AI�ږ9N���֙�����4̧���+���t�W8C�ů����p����LZ�u�*9k�[�dW�ݴ�{��N��p��R�Wu�^�U�r��4��4�s+Բ��t�h6�֖f�����ͽ�v�)�������5:Qђ�����s���}���\������X�G*mJ�J�)��0�ݹ�l_d���D뫄-�V�:<��]�+�Z�Ծ4e��̫���Rc��iq�Rv���u!���Naژ3�,�*�N����n�+6㍺�YcU���w+�@Ҷ�u��I4hM�wh;ƒˆ�
I;)
P+�Y�Un�R�r=WCh�g7���_�&X�Z�Ez�ʀ��'lt��.�̤��������#�<˽S�A���'{M|mD"Ӌ"��Ӌ�']����x��y]��
�&�[�r�V1q��HPZMι��js��f]���ۊWR��41�yC2�f}%a�(&.��/5uh jv���ee���ʫ�b�$�������&q �;#�הon�g[�P�pWrݩ��p`˺P��G�v��
6�,)����%�\a��6C�B�ot�j����>ː��gA�J���[1b��/y-�o�����nm0MU�#8`n�}t�
�|�D:$a�VE�[��^�^u��; ��szY�g9��U�U7o�3Fuk�/������4��st\h����	�ml=���3xT��z��LT�[y]Ԫ��n4]h��1Y�5����eISy�t�]�s,
� :�k��2�F�o�}%���sj��=
��嗧�9u=B�Z�sw����z�h}�s1��`�x�gw[��hM�/��jCm�냚@jy�,w�D�T�S�xSr�_&p��G��n�Qx�;F��r3����1X��kp�a�}�0��F�'�2Y�AգE_n,��48i����]�H/[�%#���]B7*	�'���H�e�gn��Վ�"&��-d��mT�np���8��r�'����wy3��ri�D��Xo�͵�D9�b�M�7����sd멸��I�ƜF�[U�ؼ�����^�N}�3�Mtl�7	��'�9j�v4�ϴT�b׽\��W���H����f:�z�hTs�`�+�^�hq�W���w�[�&�D�c�-�k�x�1 ���3Ӵ�U^Wt���s�r8��	w�KmYi�/���������b
k)'��q�Ν[�q���ݶ+���x�S�Q0�M@�r��e�x�9y�kԪ6+�}C��8���ͫ��f��G)*�C;o{y�ltw0.�f��^��_J뿥]�c��rm����\\UpE�lj���Œ�qn8�⢢��k\�-F�Qq�E�j�9����*���j��Tl`ѫ����4X5����-��ѣj�cl9͸��m��q�9-���5%	X���˔n&q�s���1Ÿ��+����qh��qW%QW��!cm�[�Z-��&
�����'8�ō+9�s��q���[��W9���$�m��6����j���s�V$Q��6�*�Am����W.sWmIE��T�[˱<c�/�-�8��o�� ����0�\�̼[Ww��m�c8ڛy�k�*����2�a<�vy�������z1{�ww��������¸�W#qG��7��ܥ\���|��o��y�]D�&����Uъ��8����zr��k�,��Q���Q:����p+˕�z%�. ��g:����ٌ~������
�k.���o���T��<��."e�P�Ю��ว#��,�����o������}�:/��,��|\��߻�Y��9��>�>%+2Ǡ,z*g���kй����������)�k���@R���z����.����<}Q%T�F{ly���}ՙ��S[���S>�2X]�n�0�{�����l�ػ����e �7�,�[�J�+���mn��6� �9�L������n;�>�ry����#��b������f��Ï��^��T��1�6}'�� �ԝCu�Kez��p���Ӵ�������]k�Ow�)UnB�'�3�}��vF\;��V�Af��W� t����~�Y���섢��g0�^[�=�%S|��|s�9���&㻮'.��̖iT����6~r����q�4��Q�P�fg\f�(���������j��wWn�T�)��Bʂ��1�u�BY	�����|޺��˿YHU��\pL̉��i-NAx��o��Ϯ�CzfI�ZL̘h��,�%8�,��o�u�|� �̭Snf�y\����.�T���\��j�1Ǖ#��+�Tzw_\M����S$5bv�qێ`���N~ɵ�پs���EvM_ث�\kw#��>Wr-s�'���3���Q�=p)]9;Ct\׫CMVwM-�N�<D��sv}��E���T<8��á�p�W�|�`��u���ž��P��!{O�^���dZ�'�ޗLz.�h:�a�l�;�ub�|���6�ځz�B�^^�����ݺ|������|}<�����$�'�#2Wܵp�]�	�;ݰwc�j�ڪW��Rޘ��QZϾΪ�;��g�����3���99s?��8�O��S��>�1��//��{�L��r���GK�ށ�]x���	{z���e֟3��Y�~���,z鵁F2�f�:��r}��vќ <�J�c��\��=�L�|�n�GvR���Y�)4�D��ww���5�^tn3uq[U����9\��:�X�wMgz����C��"^Zܺ1˂�0�}^+�����t��	|eTu��n����uL?���x�8θ|��9랪�.������ۤ�cv�
S��{R����w,�2�P�s��{�� n!n�֖;�	uK��@�C��r={ܮ�[�Փ$��9�-/	�n7[�X��c糁�a�<y)��S�|0�M�l��u'<�����v�Jl��PN�;x���������p3�����򫘰;r�%TL�9T;��[��ҙ��V)�������U������=�9v�+�����>�Âtg@�
P5 �sK�8�S�O����g<����w����{����U����wl��Ie@VA�:d
�-��u�Pn���\{.���Mt�T<��ç�0�:so��>���ݝq8n"���X%��D�tnr3�<��Ӿ��ͺ�\����+�g��/-�k|�}�ԉ�����wu`=��J�L{#+���׹'V��]mv��w}#�ذ?dz	�����%���f�.W�n;��=�\ �u�9v�,��{|X�`���Q�3
g���¢^�
��|r�"��ێ�>wrCO!�Q=�2�n��u�v{2{劀�����r��W�l9R(��:|:J���U�S�pyL�خ����i_���o�G�!o]����7��o��e�l�i�U|=0������8�&�u?M����&�#�	�{)���.�0���({�7�W��~�R���{1x*����e��V�=�b+;e]� {���R��c-���T�:�v�|(g����Zl��]��ԫ�e��1ZV>�5Ց}�}�]0C�^ռ��[;;�mC�]�B}	|�t��^]-�NV#�PI(��殬�4/���z#��D�b�h[W:�W!�X����aV�����T��8���^r��]x�WoO��������^w��e�b�5�y�z�Ks��rz�;�`T��E[0��U��q*�e0ƨ��w�S,y��vR�*27bJy�����3U�tntdR��=%|>Cl�z#If��{I���p1�	9\z�����J���Ӱ�(��u}�Ί�q����.3�m=���az·qS<�.)�No�����x	�ݞ�˹n�9�좊����+�u���^F��4ϭIW�t	�b�U!��K��F�@� ��Jf���e���zhMF�8z7�����s���9��ަe��-�|I��֩�L�R<oVi�uߝ��GD/L���~~�B������̭�;ޝ����;�@�T��]S݂*�lټ�]< {�f6�[���V�&����:k�x��Gs�գI��u�����#3�S\�i}I.����.��R;S�f�(n�o���=9���f��;-���^����َ��u�f�̒�|�KSd���
�KӃ=�_�Lc�� �*����k��l���7�M��,@�[�xrw"ї�UB�#$�`�2��(6����y�Z����{u�,�Ek�#/x�VË��&)f	Ş�6��v̈́� ��k\���$��n��`X5*�Kd��D��h����^�PJMaH�9�i݌̀m+��'�%2x���ކk�W���$[��5�!����gx�Ȯ���u�!^����^i/g���秳:�u�Wrb��2_���f�"��G�
�\�;a�	�O���;�2d�vO�Vk���	��k�+�ޫ�z�:�������Ea��2�<Jջ�4�#����'o�_�^t@��:�f�����3�tÆ�}���ʱճﻦ�`G�=7�y>��C��gFΓ��"3&;k���QxN�/�����u]�����x�Q:�m��-�}ƗxO�w}�}��ֽ�˓�^-uEDa0o�Eg@���q�w�׳�J�+/9z���:��~����Uߌ�_�Or_�'�g�hKGF�3�|���M��b�ݖ���*f�S@_@�\
�k�q�s����q��XƯm�a�%��?*�>��2�ܩ��7�[���r��NG���u (X:��Gu>+�ԇ/X�_s۞4%w��]��=���%{��tf3�������T���Ha������<�v��;����҃���e9z�R�"=���Nn���&s�6��2�r\Wv�������::ZҶ�����U��3��L)�z��:*P����wph����X$�Į��J��g��9Ѽr�V���W3մ1�5 �	�&�T�TR�zr)�V[��a��}:�w��ä�Pf6�J��(�fIAq��Q.;�<��8㶈�>�큹����.�}j��Z�ob�aƛ�����N�!��C����zUvTR�[��z銓�;9�7�~�ڎ3��aW}de�ճV�Af�AUL����_��~��z{b�/|�s�U�~�*�teu�1�=�|���n;��r���d�qT�Չd�h9��wS+��3��M{b����t���=��W��<��g�8��b�dw{�&ٞ�Jd���:73�D�j�FVw�^w��Kt���Wd��:�5����+���<��ކn0
��s��Mõx�)��_Vez�����&���o㾨���f��~�xs{�â:�7:�uw_��4��HQ�'���^C'��U�W,���dZ�
�]q�&��}�l�;�u���O�{���|h�B�F=�7�Q�ˤ'_T��'�4�g�F�������z�e�K�p�љ+��H{-Ȩ�𹛭>�[#�/^ӅӓKL{�������N�?~����3��㓗3�*���ʦ����]{#�G�/FS�{�C�wS���VR_t��I�n�#u�'h�&xTA�Rnl���I���kMc�"_m���OG�aNѴb޲�_m㉑���x�Y�ԡw���(����;̈́�Ϭ,�\
>�6w�:�EF����n;JT%�'�������/C�O��W���a/o^�O�g`^���1���g��U>;��&ɻ��VttV�#,��FWK�E�+�z�Re{�u�t�zP_g=�G*�nm��]����ѓ��cy{-�{���J����T8/|1���ަ9�+����&�S�F:�=�yZ���v�۠�r�(�Ih����#qE�L�:���w���O�e�Q^ʊ���FH�޿8���Vm!���A�Ϥ�P$���$r�w�L�1u=I�C��;g�+{)rX�&��Yɞ��^��8��W}�Yǽg�Y���J���7�s�%�$/dY��a'^���=��B��Z=�{��ȍ�WgTO�:�ه���()f�/X�.�+�o�vɲ�����%�S��CV:��GW;c�9��q�-&㳮'UuEc2Y�p���}����[�"g'�NXq���\ ?w�@�0WS�!i�A���}!�������É�����']�#&��	N���荙�fI�l�2�����Ց�p��kf�-5}&���@�>ʟD�U^@�=��ȅ�(T��ܝR��m�ׅj�W4[�<$Sl�+c���Yچݱ�s�Y��N���>��~�Gʐ�{��]�3u����3T�c�.N���u�Z�@o:���z^i�m5�N����sT�Ź�5�]���Z	l���Ծ�.]�ڢ��]���.�0׀��l�7�1Jg������%����]�v�s�&}U���ڌUSz����̖ɓo����5C.9Q�*�r�Qcpt�uԬ8%�𥆮�F��T�vrｋUc�{��˅��cD��w��{"9Q�6n>�Ī�醣'��K[�Xb6|=�*Vt��(�}љ\�����^�=����3�Ղ�q[�;�Y:���N����=�'r��K񎸯V鸮�.1_ /9W.��B����23������}�K�P׼=�9��3�YeW�oQ�7K4TE��w�X�`
XՑq+�q�W�+��m����~�\�Y���2�~�n����>%��_�;0���#�'�+���Y$\G`�=�W��޹�vb��g+��	���q���b�m=jI*�e�P&t;��SNBsi�?OX��xA��d�k��W��w��F�㶏���:��v�6������Z�
�3�@�X*�8�{���Bq�u�I�^t/������К����,y�m;}�㵙��}RͲ�.k����KtS��QA]�J��>��+6Fvn�Z��eqN�L�^ΩQ����jހX[:E����D%��b����[��#��E��-&ì�xwY�i�*�S�ܚ��z�t֋�������׹t��d��
��VJ��y�t^�ѕ��;Gs��3��t�,@���詞���([�׃�s��VoP®#���7��;�z��D0��{�Dmҕ���z<D�3~-�J�<)gm�[���~�G�Ѥ�G=�6�`��{f��Ҭ��UZ+I.yR ��`���0���0��H��x,��͜u�J�ߢV�:��G|x�Vk���z��m̒�*��� �ԅ_�R���i���$��U����q�귎�GB�ξ�>�D��ǧ8��3^���ċw=%CY�V*\��V�b轓�o�]�\Wf���0湐�����7����Lz3�T|@�W.Nع���������g&�c7�܆����c�^��(��{����'�R<���� ��.�V�C*As�]vLq�kr;ڟ�D�!^���^?ok`���p�嚌��^u\��P�7���t����F�'��Ǳ��/��^iɩuu�?�"�i,]�t�G��/	�x���W��.�����}�3u�ib��>�s\��ж���}���q�Qn^��*Ρ���銈�`��[�)��<��:Ջ2Z��R��O,��M?z���bb.X6h�K��b����s n���w�AtU�n��b� ��ձ��SE|Ҿ��#*rW��VSp#7mN�k"����Z�xd�d�u���ZvQj��i"�+P3w��/P�/{Q����94����U��r۵����MC��
+Yߕ0b�hQ��ߞS���'ON�f�)aT�,���'k��t��W+����aFsۮ
�@w���{�38�zq~_�rֹ<���3�n)���4�w T,Lw���^���9z�F/��<x��+&�X������J�3	��֋��Fd��ۺ?|7��=�y��;u��f�.�T����]�>�N�O�w�7�<m�Iuc`LUA`������N����;���W1/��b���+nmHˏ����@���p� ��I�&u�t�W������L_UbsQ9VdnnF�-j�zg���<uGg\��f� ���iU2L@n�P/��ufrw{s_z���Ț���=���B��{�ٷ̎>�;���]w�E��K*Id	c����h��/���U~G�ޚV�����ۑ�ھ{���>�Nq/�q�����g����+�3��9Tr�[�J��m��M\b�x�HcS�㿟�������ǿ�{���խm��Vֶ�Kkm�W�-��km�]��km�mZ���m�k[o��jֶ���խm���V�����V���嶭km�m��km��mZ�����km�mZ��ݶխm��m�Z����km��mZ���vڵ����jֶ��խm��ڵ����PVI��W1�P�*���@���y�d���eg���|2��%�� (��T��cE�I�
�ي��Y��T����j
l�J�!k&�n��jյ�U�V�m�ղ�M4���-l��Za&�i��Y�3KdƳX�3Ke��kYAN��Z��=��ƵeV�֪�L�ɶf�K%�SD��a���d�,�Z���5L�-f�mYZM�k��VZ�[S� '�Py�Pn���lt�鄅l5t4��F�\(R�8�u��d���n���ѐ< �ރ�[v�݂vn��7n^  
Q�X�J �v�� ��┠ (6R�5 ��f��Gdu�)�֪s6�� -�4��@��tt��p�:wq��9s5�k�������l
����w-j�k�[��w� ��q:�ں���:�뺵;�u�V�wZ6�gU�����j�������v����V��Z�;SK��Z�Zխ��5�ee� ��u�)�TN�WU�wU�]����n���uZ���;uݮ���;�Ӯ���u.����n]�w*i�8�]�;�ݖ5*3MkCQ� [ޫ���u���ttZ�p[k�s��5l����쀤�]UweműҮU\[��w-��pۢ
�m���Z���d�h^ u�\�U��vt�g:���7mMj����j�6ݶ��un����R���jۻ�ֺwn���ws��;��������Y���� w^�n��M��뫴��f��v���5�n����w]��v�r̭3v�v��mkn鵪u��m��N�((ۑT�'-]�M���� �V�ڠ�s�ӭ��-�J�WYɤ�v�uPιCU�N�3�f�t�[&�O ��H�wP�w �� ����&�- ���rn�pPծݶ�      ���JEP ɠ  �@ S�R��  �     "����*Hd��h`�4�4�h�bO�J��!��0#@dшc�i���4z��     �BdL&CA��j<Q�4z�6��d�V4%��>����!�H��4�LZ�B�� U���I�䨊�}g�a�eQU�UPMm���ő�TTqKo7?��/�o�?���̓�?�BD���M�API0�����EPO���H�	H��'0�O���>���������?�ڨ*	��/�uƴ�`��A�� ��������f��8�00Ć���?�����x0�߮ZxR��ͣKB��KfK���i��OP7,5[�-4���q�wR������l7N����[m��X���^�kQݿ��Z��-��K#�3�N��F�|�4�
iR�[��S+F�Ē�nD�hXZ���gki��( �:.ht�s(r���ҝu��k�aR�b	��lf)�a�+!�w����zl�p����W	��T5A&Y���jF��,�W1M�� v�soӸ @�����	��i�Wy+l��-���[��u��Y�P�����[L*	�fCt�5�'�*�T���nm@���Nn
�#��h�@)	2j�:)]�C�c��Z��aʱW�1wu��!-�uxqbI�X�lm�X�P���'E���F���r�(&Ԭ| z��b�ݬ��P��(*t)n�	��̌<ݛvmT�fG6�MP����9`:�
sZW�¡�kfVZ�5{��mbx�h���X��Ɋ��A`�,�/H�;���k�JJ�B�5��f`�lm<s*��(kw"�YLTT�̺���B��Q���Eʼ�ݺ9�)e`���X�z�׎l��49S^0␅-��܋DZӗ+Iw��^���/5Ob�>y�4LDw&�qK��c����j�¬�n�݈�|U�Sb;nٙwI�i+ciu�*���h'M��ΊY�u���AJ�b��TubY��p(�"��\+N�
���c��
�%��u�e���=��M2/F�C2#O0"c�uJ��]�f6n+4+4��:�P�"U�XNe���\���F���å�Z���3���7 7�й5�$|G�C�g2�	�A-*b��/�<�,���M2�9��DjU��Uv�8(���f�b�fUЕ6F�i1���hV�) �k�;�Z�����Q��!(l왶��,=��kF-��E�x��U6�f�Ahڳb�I�Mӱ��'��[��sQ6��Ecu65����z*:(S8�q�#�^S���m���r���D�f+�F�H�C]���#R���ӆ����BI��ʩ[��o\50V\���Y�R�h]ռ�gP��:.��O�b�u�W�i�sn�M[K���&�P����R�9&��[�Ha�[�a��ؠSqJ�c1�-��%Y@i2��y��MЖ�4�ȅ�ʗ)Z-��WM;n�8����=� �t��[r�.��JZ��n1,K�j��VBE���lF��tl8)��j�Zi��cZ�2��]�P�.�ݘ��)�]i7F ����xa�>��X��P�zl�LۨqF�UwX�	�Iz����tm�8�&������l*�x�7q��#K��;�e$UkAn�БkpÆ��[fm㻩L��V�����ں����E꥝�7��+h��,:B���Ԉ'Br���[�)�抴7K��i�+R�暶�;cq��M^���X���-�y�+l�=���%�X_43*�N��.���f�(�Pf�������^�n��up�Eآ�PL8Hm�y��.GcpI�k
{3��ӕ1�׸tm0�jf�B�� �u�.呤�R4ؐFŪaK*�L�i;���M�9p �EaH5�Ym@�$�,5��cr�B��u�u(��k(70jk�;�dd�.��K ̬nhnŗ%�)�9�fR\vo�!ZL^�����fCO/!��*�i��!�Vܺ�A�XL�K�YLv�F!��l|V�G�Y�wL�sm�m�sT��0���2���4Խ�&����쿃=�U֋�*�sV��p	�Y��k��`W��*|i�v�&��2��EX�S�{��-��ua-2��S;��[��;,�qQ��H�"Ѯ�$�dꥃi�Iܡ���`��)�(m�HiIj��D�m��5j2n�	��wNf�`�tv��f�$��Y�u�NJ��pQ-�[	�9�wwBQW�
Z�ܘʒ�K)�a/3Zh�˧GS�e���H
�`�]���WgY�E%��I�4��uef�\��h�Ȳa���Z������l�3�@<ȣd:�&R��hi�\��6��(�+��"��T`�oX5��[���u��	�2�XXB��R̃lԋqJ�K�	��A��P���8�<��Lc
��O"��&�9�mФ�C-�����P��ǙB�����%ǵ�nSl�˰��2Qt�h�����m�+�Y#�5i����XX�Vt��ؔ��$U�mh8��-W�،��/n@���A3Eȹ)ͣ�*�׈**ܩ���^V����*}a�֡�l��v-q\
J��7�ǈd����
��섶6�3ww#af��*^;�X�b�����`�"�{��Q��(��ht�EE����f[�-vUʺ�e���k��x$�۽d-;�zv�
A�\�T�� fVT���f�&�Ƃ���Ȥl��>u�.�7��
ER�+];ƠȦeZNRzά�M�t�F���
�ޑ�v�mh����n�m��ڔd'�fG�ݬ��wX��j�&��]"P��7iI������-��*�nV1uf�D���sr���[tH��Va���Jm���ki��f��Ҁ�iU�!4\�:4��ֱ��[֬HS�s1j̆�sq�EV���b*mҋGv����{��T�[%��E�nL[���'.z����&��lk�-�rfӷAj�����y�w�
2)���i�P�K);"�Qڂ��Y��MT��9F�R�Č݌��2������
������Z�2�ᬤQk�"�n�u��z�1Hn�9D�(�P��U���y��,4鉙�[D&֍�beB~r*X�5��+�>�5l�5�D�;�a`)����ݟ�P�V�u`l���q����L���V*Q�KB��-�خ�,�8q������ﻑ<�$h�����XmT���mKu�"�5��MJ��Mҙ�)k�)��M.�맘^�Gel����7
����U;r���nV6��)^^@����Fe�8ee�D[{@�ғ���7cS�mTwy�6�#lK#�j����w���.f`��F�I�!��t�X�q�J9T�^�ɻ����s]H�e��uyӺ���Ft�(QF�|����\�)���g"���7vl�c�����w0݁-,�R�`�H����liRޱ�˩��!*�޺���(Q�i�y[��Al�Ww6�66BS�j:7\��h�Y������Z��C�=������8�H��vq�&����7@w��*Y��ٱ�7&QF�?�*�I���-x�����64˹�n�f7a٥d8�ֳ�P���hu*Y�Y�὎M2DHz��s$���K���	��֘�&j�eAB[�O(�K3Uu6َ�Җ8���)&Xʈj�Y�e��$��Cw�/�iu���F�Gv�\�R�;:�]�֣j�lƭE˘�A���,Xe(*3fx�V�A�#^I��/�׃�
}�
&�e;�Oh��K�r�h�[Z��[orR�a�q�� ��C��䌺�;yu+1'��V����f-�xi��X�M�UM�Vƪ�����c�!F�AǗ2��b��e��ֻ�"���t�!�ڂ�e�v1=�l=K��jj�
�t�Y��Xa�(�/u���Wm�F�1M�p�4��oF�Rd�m�̏�fb#+g��f�ٺn>إN$����7�g�Ӛ@�CVGo]��!�
ڽġ-�e�[�Ɲz��� ���>��t	��+���{��U����O6��|H��PC��6���)��^��`��9y�S�ѵ�IEU����y��V���3���6�<��:��R���!�sh]�-�$�p���k }be����� ��W�Rwc!*�Jk�,�YP^��ШM#-��u�\�Va�a�w����!�E_�j%�uilZ^�1�jY6����1����p\X6������N(˛��h� �s6�nj<yzD��44������ʀ�~Ѣ�Y$�B�_e4�5a�gm^4v�i�Qh��Ұem��+:Kc`��<a��퇯�`�n�RBvVk��M!)i-��mo.YN&0*�o��ƞդD��P��Z�n�Ƶ��֓&Z���ZD���[t�"+U�p� �J6�r�`�K�X�ˊ�i�m*�5�z�=8��ɰȶ��+q)P�X1�ᴴa�S1,W�[0[���Ad�J6�R��Z;-��f��oZ*�ӽ�%[X*���	)�D�e�jB��Be8�U� �@U*�6NH �(�X��d�SS��I T��[؞E���] ֛�
�b��+Zy�+'V�l-�;H�3��i� 2T�`4��F�����]��f�����ߡ��	P�
�ZkFS����qK-ʰ��w�h#2����zjNR7%�䫽��t�� ����ے΀@y�'M�cMSyV۔`�a9��y��1�W�����i d�p�2��FA�YChW�2��o�P)�0d �5��)��ɬϖ?�Î��̴Ȥ{�oe���*}�a�Ӛ�:f���S$�,cilt��
J�wj���v�e�(b4�nC����fP	��`6.���Ú���T��0��M�n�']���[��\ǭ����-����̫=���WYKT|PE�[%k[�����e�3�VX��q�a���~���n�]iÔ�t��}G��|<�9�O����;��mh���9�z�P
ud)9 <$��+y��2SR��-�u�}�� o-.������Y��xw�R�Ct��9���!f�H3d�[��+�z���jo���5ܩ�/B�U桵������Վ����qRd���ANZ�՗�7n冰�������=g��b5�sCY�!<l�P��絲������}���u�>���쩜�b���{�"��W|���!�ܠ�S<�v�w�� �s"�{>��
���^��h�s-�oe�ZW)��QY#��o^�-��򭾨���k�۠Gxn�cK�`˫�H��B�� p>x2���'W�@������[C��E��yqT�+��\��B�%����dC�����b��V큱����jک��V�j��P���4���t	K��y��W;/Uڌ�hi�w�ĕt�((>��l�:v��*f[�mq��d��HP���ύ'ԾN�nY[�E�OpnI���hS�u��97cu}m�2��
�l�ɦ�M�q�.�_P�]2��:���!i�Ήi�����`�y]|v��`(�oC��v��j�C삅�f^r�ko4�/�����,�Ö���]�;��vn�u~�����n"���[Vk�K��cg{GI-s�}z좦��;�����+���j�5�.�XkK��p+�Î��	ǲ�]�H��[)��(�a�Wl":f��-7�b;��NKҋU�5�Uc� 	y�(,��.�s�ǜi]�&�<�� G��0'C��'��_;�v|��h� ��v%�9:�>��8���Q���ȧ�VQS�f�1\�e9ZL�m֖V�gF�F�
p\�r�nX��;226f�`k�A��x��:,���R�K��4eɌ4�t�h�ļ�$�5�:7ZV�����S�ڰQ<А'��D��+aV�b��,[*��wn���chmmH#g�34S�vm�&���J<*�Ю��N���R�]|�0b���v�j���I)vw��f���:Zm��ӗ�����h�� �>�瀍T���
�ءMV�$��󓫭�VQ
��L-��Ц8S���n�W+�*��0:Y1G�#��n��k�6�o"��i�n��v�V����YK�%u=\��H1�,՜��n `���֡��ޔ�(�_�%�j9��b8$�T6��D\K/gn��u�#m�O���gf�%��rh�vhl.�����3E��^��0$�yq�\�\�����{OU �ҹr���
�HV=�+��g����Z����˫4ك������J0�G���ә]�
mT�=�j�C��\��xn�5�;�T+T�B�vgA�N��m
��u0%�l��.��q[�U�Ȯ�*�̸w5�5nr�T��{b;H�.�$��ɉ�3p��E��j��=�=���d4^��x]̭ ����Rr��Ģ}��Dl�	(Q2�4�\�֧Q��6 l���N0��������<a��t�m�uej�i�<B�Oo���-�`G3/�����QL[t6^�BT��ĩ����7:E�9X",�3�M$ّl����0噵ڊ��=)�Ǣ�����-��l��&,�vc,Z�Ӆ59}GNm 
Ve��:�e,�Q�1�91e�w�=�{B�!���uz�J*��;`�f�.�ܝט��`;���6�f�WR���M��:�"P˃I���3.P����ȁ�
���{f�k�`\��*��9�ٚ�:<^����v�;�鎤��Vs��tN
!w��}vV<�W��.��:�E�b;n QTt�p]�5:�U�iv>S[�SIr��T�b5�Q�js�2�f-R��8k��\��x�X� ����X�ӷ��Y��H�
��hL����e�T�ʝ�ݬ���:�d�9SG�V�I_o+26���
Eiԥt'�dCJ�k��x�0�$c*��Z�����d]Մ����MVZ�kj5u.BLf����@u�e�NK���"�tc��fm�-u@�#]��uՈ�V��%���i���lc�E+$ʇtF�3X�{��Vn�K�*��q��r��K�h���s�E]�����eYB U�k�r�m1�u�-�g��jK7.�����ݮ6�4*Bi�ǱY�;j���:͋NV��s�'=��s.o˰��u�p�	�noKə��څdu؈�:C�p
��%ʧX Zx��+K�
���0��]*s�9&gen0�FP�Ԧ+��[R��/��M�O��Vr{��[^h������7���p���2���ѡ��*r��zR�ȳ��wעC�6%)�y=jJ���]uKop=��N(�s���kQ�S�.���{��\�Vo%�0�������������)���}]��D��i��Ȕ���B��:Yo0r�a�zN��mX��3TŪ�//H��s3X��m*��҄�w�0Y���/��\�gn�7�����T�[�B�F�y��nt��r�e���׼�V��Sv�m["�p�
��G�v�v����S�:7���1]W7J!����T&l���~$h��ҹ�Yݴ�m���c��������(�R��#�@v��I�l��(�����v]�F��h�R��Gϙ���nA���?��6��AW���C>�+A��G�!,����9v%��P�0U�-O�lKJbU���n�&)|�j "�CN*3�e.�xo��8*2�����BE�}R�o]i���ʁ-/_5��RL���욊�32)H��L"�#nOq�
-�q˓������b��؀��0�}y���=��RD!�J���L���Ϯ��u�Ǩ]B���5�.�%>����p��'Y��[��b'pH7Uu����gU��f�[�ƭ��)��ޱN0�!a����Ef1E��n�Y{��:��-L�Bc�Nb9l��Ȟ�5|���R���SGk8��r�c[u���A�p�B�v&��yob.�n��6X͒�P��@5G���w�^���ю��41Vvp�U|w��k��������vGk����4z��f[;�10���K�4Jޛ�n�E�����w���
�DMׯ7(#�Qdu^�I�9o�2]�����8]�9x�����;��w5�tWʆʙ���.��7Q2�f�s�YG���] ���reK*<�D������+"{�@:�$�oyoE�']`���yr$Ђ���;��jA��V�ۤYs���܉�Tu3���jz0�ǔ�0a�ٖ�n����K(qAv���d[F4�� V�V���n�J|���1eԜ�V��óU�ƸoI��r�&8�K��Gy��{�j]:�XB���)�ؕ��rJ���Ю�k���Nz"kQá�"��ÌSx�X=���C��֑���SH4�[�]�>�O;�Ç���}�+��
lU�?g���1S:s�͵Xx���:M!Vo����=��=�aև B��yS�H��>�:��7z-ݧ9T^m+��q\� mV�o��c��D�a#@�A�r�=Z��:qh�<�
9���/�7n�Z58kLY���9�7��C�e�D��VI�������au�Ҡ��ϡ�u�Oz�y���i^��M���H����j�J��ˮ�����e�4�T�M�y�+�%�Z�~����ʅ���>�Y��J�7�8�)s�7
���ҰI*[@ʛu��٫��շ���J�
�W�n�b50B���A'�{�L���F�Tܻp�޽C�H��B�eSrvu:�SEFIUu`^�ƳpQtx��e�u$�]�b�1mi�h�W��kz�A`��V���u�{�']�j!GE��a)�y۫J-]����1��+��w��*��u�m��^;�
CT��ƧT{���%7��<B��\�9��yo�c��eG�ޱ;H��A�y��Wf�W^�+�1�W��-͌br�j��	��a�̰����6Ş��[�0�,a�gm�z��4���q؆R���Ǡ����Ӭ��+͸��xR5�Zzy8�&��֪Ҿ�w&����SH<��G�z��Y&`��͇(+�.�(6�V0�3r�N��7���WB�K�m!���R��RD$P=�ow��'��蕵�u(r�!iY��̌Y��z���d��=.Z����.��
j=�D�<����Z��,[d�v��)�;\����т6�.�y(�$DVIO��ݕ{�	p��.�H�� ��	K�--N�Ol���N�y.	:���YMqG8���9�LV�5��ީݵ#�����"�-�^��l��V	�1g:���{��a����e���J�Ŝ�]�_3�a�x�Sx]m��g��Z2��rKŊ>iu�j�.&�=[�3�f��-��-
V�(T.dplԕ{���@���I|M��X��\u˽#����r���3q�ED\��>[\�E������SnEԝғ����� w{�iq���>9\�M���i�"�#�K	|���))E#���#;6mʎ�BnC���	$�I$�I$�I$�)$�H��R�e얤���$����P��lU�7�%�h��I�w遣n�����t�֩.���c�J���Q��qu�+�m�)�H�s��P�_R�Vv62�y�A�@%w�`��-�}a������coC�:d��"�Fp�7��m�Тǒ��FZ�r����a�3#OZw]��*9�=�J�.����'���t���\������B�}��Ԭ��·qe�<[��.8\��O�>g��>W�<�_���o��ڪ"���� T><w�Q�D�?�M�P�F?����v������l�Q1¦f�3��Z���0u�jK*�:�r�WX9O��;f`�����2����z���I����9��jR�^��9�����Ds�2�c��ӏ5�]'v���{[��L=Cm���Ĭ��@�v
� �mܙ�u�����:��>�S�5�BS��\���{dc]ڤ��fb�ȧb˸X�=�g��q�KZ���/lt;�K%�qV�ղ���Τ���K��@ܼ�R�{�`�ב��L�s�
��7/\��1�g:�s�bI*�u�]fu�WWu� �v]Z�)̏���67�>F��N���i�lu�57��1r�}> ��0諝�r��l'�;F�5'Z9�;��(�2���!�(��p_)=\�Rwx���'�]��b M`o��%�{�w�S<y�b�!��=D�p�l#yͪ�Рh4Fm37&��^��e���ь+���q�xn�n���mЕ�v�� A��j�##W��2��"ᤗ(\q���h������uJ��!\��<,[�%`���z�W;���&�=�z{�ݏ�B*R��P�	I.�`��6�N\g7�r�����H��9��h���Δ�;�9fe��j]pP��� �ǝ�?�$ wE�LT�Ԇ5B+��Q���7�maV����K;��tp��`�&3��mт�F��%�u�\�/_c
mu\��2#݂�\�Z�4�ʂ��=��8iɗ��Z��i��-�M�&��Ӟ��ӀI�m�t�����]7q" �G��*�6�م5@W*�y���^�c:�r[�^m��V�1
pTŶ�C"
ŷ�Dl��y�49��k�9Au:��׸���[�<��pԌ?��;:�?���V ਗ਼��k�Ƕ��B��]���V��ʰ���Q�-��F��o#S�������5�>�}�y��m�����c�(]+d�X�����weq���H���v��Thc+(�3�wp��@8>t���q: ]� h��J�j�{I�� �Q�Iʅ�f��S = ��솰f�����i �b��%���k��e�);:[:�gs	�����úҷ�R�S�1]w�sB��:1P�,J6�p%���^��D<L�\ڬˡu�jrV�cmv��������[I����Q�m]�|��\]����]�$L��.n������,@1ԉ��Noi���i"�c8؋TI����������q��+�5{�.�E��>!�"X�&�Aʀݐ�=r�=�Y\�K&)��ҷ�q�����c]){z���)���
�(`m�砉�L�c	��tj�*�ݼg��V0հ>m���9����]��-�<���z(凥�-���8r$Ov]i"EZL���qkk ޗ�V�5�0dC(�]􈮗�B`�fsL���L����h��-"��`ִ����޹E7�A7V^����엚��Zj�\��I��Rc9bY���:�a�i���k�k��:2�����g�g ʮw��9^14<�\*�?az��ݽM#��˻��-`ۢ�0# ��u�3�u����dx8^�]�>I�P1gO*Pl5"F���Z��n����8]s7s�$\C$G��a\�+�0ui�&*3��j��kyt0U��q-�Ḽ웈�s���g�X�}VP����9J�d^����p�͸�J<t��t�G�L�OO�-$��.� ��TJ�uX��4�kTJ7A��ne�K��ѝ����*Ԩl��C"9W�[\��b���E� �:�wV�F:ɀ��C��y2'R����r�f���PB�[�S�m`��`N��\|�����^�Ų��ܷGQUe����CB��->�9.2��q-�w���[�m�����]��m�+�4R������nu��^n�Aq����q4���[{
��+n�z�!Nkഎ�ŦM�PY�
c�$$G�-�un�g^vR!\�a�&�c%N��p�W,���j�!�+�m��8e�v��Vf�(T�C�H��K](-����F�Äa�9�7�U��B��Տ�m��e���K�!�s0h�s��g}b�)��7C{��kWſe��ݡ����3�AQ�6�*�%mk�\�kW-#3:��ys�!�vֵ 8��0c6*+��Q�e�H�^�s��1"WK�2]DU�S��G�N̽�J�EM���#U#�elU��_f�Ǫ���)$t��6�<N�1�O��u����$�8��`�%-˛�(�O�XwJ�V����3+LC�?�Q�'�F��n��Խ�)(�^�3iY�͝!����|i2�z�u,;�,!3�Ҧu�tP�n���(B��#��}6��L�蚙l�42��Z��1Y�h߮��dt]�{���}����$��*��b:L�k(��l�����7�'��i�nV��\�0�r;��p.�w�j��#E��r6���<��!��y�ێ� ����LHr�D��0;��ы
��68f�e1�9�J�P���J�=�o�K�[jU�۩�]읲8�J�[��]'92����=&C�,��Lz3�6�_�WW54z�S$�"�r�:��}�Z+!������7j��tT��� �=I+G���Ԃř����-�(fp7u���nr���������	A���7뼝7�rF�^;�1+ չ ���: y�^J���!�o�*�$WIy��tJZe%ӹZ2�f;ٴ4�=�ķ)����:=._2]�7ٍ:�Q��7.���R��XPu��Ne�}�:��&l=)q��2p<¤��[��(�-Tv��%O�����������t'�e�	�9����g� A}N+�+��V����%'_V�ɿ"�ڳ5@8�v�ʕ����hEM�Ճ���|]�/H��q����\�R�ut�����l��2oM��)�#����:m�aVn Z�m)�4��+r��b��6c���7��ɡ���e��f٤d�/֕[jҔ�dy)�+�ݭ��Υ����5.3�(f���&�E�rK�U�Cz��K�*�t^h�R� L�b�e�j������qa2�V�v<5�a52�c���>K%�wnގ�-�j�'��[��3�{@�n���Vt.mP�k�d�`Ϭ�X3uTH(�2��
� �{k^bs�m��aU���
��9+�۫�xa3s9�$��mB)=-��:�ZM]o(�D8�ӭ�| ���˂�&�bA���0Ԅ�y�)����i|�D��kEՌU �]�[A^d�9�����\nb3�ާ-�O�bw�}���t���İ�wV�b�S��/f
�&k�,�U�mJ�ƅ��E�{3J6��2Zt�s5j�`5�.���++t�Iy�c�F�=:#�l8��ye��#Fl�5����Cc[R]nˑj�;X���8&���\{0��v`��j���ma3������;��n3]��1�/V�e�v�F�X�b9�m��2�.�ZR3A�ٴ�=|yc!h�׻@=T�
��[�-�/� ������t�m��Z�nҤ	�{��Vi��+^�
��ݞ�;�+�vYi��\��u�YB�q3 ��k(�#Y��$�/6̔2`M3A�,�Xy����a��V�(�Z��klD)�_<��]�	��_v�mV�CXW�xD�,`�t�PW+��ɪ�����O��l�g"������P��%i��2�����!�	̽QJ3q�n�l�5Medhh���DIv���YJ$�!�]r-NHi�=�u�wqK,���w^=M0�Q9d�J�=��f.�����]�� �t����i��)
0�����9I�c���y]FgV�9�=�+;��+Aۼ��#����.����b4ҵ��w}K^K�XJ`IX�ru��Y�bL�����"n�)#8�6�GyTq�Xv�"SI�Bvy�uj�0�m�a��V5x�,h�&}{��ۤi���f�m�m�R���[�j��6��ׄX3+d���,�Z��/{���q������C��$(O>]��%��
�� ��h\V��|ȹ{X������׺s�E���w��V�ʂ0�J���A+[}�5F���� B��wTY�,L��[��VA����*z�@�t��yҋuѫ���O|Dk6�K'`n�ڹ��Y)�
��n��5i�K�IJ'd�5�Ұ��B LTB^dq�іZ��L�Ӵ��v���9�EJ1��i(�ʆM�Y��x�Cf�܉w���1r�43�ܶv���%�*�i|��'6�'J�R�C۹/��+s�3P��9%�Z{���HY��'wJub��C/
����z%��fPk�v����h�W�,!\��w��-��.��i3��.�]N�[�Yt��Jr�*_t%����Qs�|��}���x)�
F,��Q](䡘�x]��\Ǳ-�Un��p`���-j���w���[�mrTk��H+yօ��T��s�@�:���PK{��%�]C!f�a���5�p����b�U���հv8xu:�r:��|&v��q��F>���2�箚��ͭꚋ��S�>9�q2���R�R���4;��I�[XU�����}�j�V�61Qlb�Egk+���BHV	Y��G9=�r�&���f�c2]>��{�r�f�*_V
G�[	����Yyo.�E�{���{�޽��(��̝ԷR�5P�ZV��ٻ��W<����*	R5��z��"K�sHs�=48JF���6�ͽ�pq΍y��`9[F#k+��S9miŠ4�T��j�H�V�,<[k8��,����g^b��u��lQn�W�Ζ�G#�U��U�^�b^��U�9��:=�>�Ŵ�3n�U��]L�C��I�]�FZ��^��Q�Ӡ�k���US�f�fkq�w9�=����=W!{�oS����HA	����y�`�rB6�v�om 1f;��K�Fv�bL'��m�R�ξl�L�TNh�J+���iK�0��uxp����8��E�k�%m2��S5@�����Znq��L��Ǽ��#l(-\�8�C.�c�z�]9���mG�v�ث/�:R��ѩ	ƺ�oY��=jyǡD^�s,�u�eD� n���n�k�O�4��R��C���Lf w�1I�7��*s!-> ��PL}�͗�n0�3�f�Rt�44^�\\�IRVlҚ!R.�#J�r[�\iВ\�9��}����>�xg�j�Ř323 ����r0� ��-��h6���'$�eZĬ*&�+'�5���"��h�̪�b��1��3���*f�d������.3)�PVFfQ0NYNKZ��& *3� �6�؍��!�șH��2�!��*06�<b��1��XYRqk
L���',�
k-k"-`�S�T%�)TنYe@DCT�Q��hjc3}�SV����*��PIaUPD�5C����	�F�!TT4��b�b���Ŷ���U�k"&�x'[�~�q��m���[l����t�s<�7��N����t�r�W'-	q]NRɺ`�C��_Q.<)(�����z�s�d]P����C᜻�a�O�*�;����ة�%�[����=-��PW4z�HMF�Q�N-��f�9`W��N[lװ�_[���ζ��:4��U��5VBkd�]/���&��2��r::�ry��v��`Ad�iy��2�]��A�̥��Unocn��;mI=ǐ%L�8�PY�d����"���d���P6k�p)k���y��"
W兦gR'_�3�(�U�H�u�*"��ףz������;)tS���) ]GK\.LT9��Y��W��c����;���tz���n� )���1S��8�͞���زN�׾J�,J�K4U���U�x�`�mSN�T�ؙ
�!U&���[r��o;��eھ���l˱��ŭGY=4�ʵedN�f�E�����s.�JW/p�T�����H���wT����Öμt'U�׭��k��m��Ү7h�rc�-��B�:��G{�W��5�9�z����j:�Ugo�!��W5U{��H&�-���$����M-����� $���s����9�e���EWc��l^ξ��g� H��.(��9�s�]�ԣц��*�wW4^-�?Q��v�!+���������ۍ���ت0�P͜���Ք9�]����ve�H+�c�[oǦk�p$� A�Vj
mf���{�O:��/_��1p���2���M��p�_=�{�0�Ŷ
�֔�Q�>��6u�en��ꌭ��sX��{��bsr�,C� �Z�S�k��֓5%�5i���Us���sQ��RP\����4�c;��M�=������1�(�`�Q�����٢�K���8W��b::^�@�L�_b,$�}ݥf��{���:K��1����&u)��$�J��^� �w��1�������j2*�����M��#�F����b"Q��ꨐ�ט����!v �q`��}p�{!n?��h�u]����rP��Ꜿ��I�h�ţqy���p/c\���W]�y�$>c4����FN^�Uۇ0��
a태��	�e�F��P�Qz��i�vΒ޲t��Q|�6�u��2n�U'��`���%j���w���~Rl�$YN�����Qϳ*��1"ud�EA��:�T����%{`h-k˪�7�=<���l�w�UX���ho����3^*?L�Ǎ�XV�ZS���W1��>T�}Q���`���	��n(pZ�f�ʫ���^#�4��0�j�S{ˉ{!�*�m�t�@��T�vr���Ύ:�k�A���U�f��>��J1����d��K*yC�Z�>]g%�.�EE��=Adw�@һW6�=���ks�M��q���!o��cb\K��Ȥ��g�����x<��Yp���0V>WzO�*����zma-hs�Z4��:R8WA�SEp�{,�ks'�[�!{O:�[ܮx?_���_\E�1��^� |�n���-�K\6��_1[��C�9嘱�+��7i��s�@+,��l,��+��2�:/��Y��;U7�"w��%�V���)�|������uX�i�i7��:p(� /$��6#`k��i�1��=*;\���Q��
��,Qv+�����u�:��4ߴP�����g ��Qv(�š�,n���%��W<���H滫h�n��K�ؼ�/�B2Lͪv��U��,r�i\�u(����SE�d5s5Ѱ��٬��!S[%,I�3�����k=GC8�_���e+2L�k�'��#EN�����Ё<ʸ6ruzJ͡�Rx�іP��~�x���T�qw��K��e��2�m��b�a��I��iA����lAw4�`W\�sv�Z�>G7#S��-�s�ef��L�_,�Q�Gn.}jȊ̒��^Wrp�}�������G�U���E/�W��� ��!���2$cI�[�o]Ɗ���<�X��3�Rw$��ת�AO�x�u^�i�,�JÛ��ү�r�S h�Àŋ���l׭�8�F���y�&��'z��H���g������/U���gB,�pX�/��4��P����I"e����~ޡ���������.�ȩ��o ZP���[id�rg�E4��nם�PoF�V�H��,�ujNs֬K�۫��^>���-��7���N`��^}t�Y�VFuNA��G�r:_{d؎e*}b���/[�cqC��+�";0;
a��{��ݩY��n����sK��*f�w|HH*mh7���=�b�IW�[�w ���o��o���m�wF�Eh���]�_Vh�p��)�����׵�"mC`�D������8zg���/�J��j-̈�b��4��8rtm��.�h�f;ɺ�b�:��RR�C8c7H���n3�$��1X�z:�Z��,Y/js^F-��Aj������ʧ��u������%ID������d������.�n�$[oSM�0^'���1�yp�R����e-��a�8,��b5���Cg��+��+���Ք��^�$L�}�	ز��8V\���0�"o}1T����u�/��x�IPxw�^���FY#pVGB�멓��w�ai���Mfw��b��'#㹊1��Dhv�\0�Z<JP�J�nf�%7��/���Z���p��$F5e��L�E�z(0��<�"h�)��t\!w-���h$���'��S�gىh���T*؞z�<B�x�S7�y2�/�� R�D�@�$��r�z�m��YT����K�x'�K�[\�GM40r,A����u�nj�`י7�s#{;3J�6VZ-ר8���4��~. |)�R��NG|�t�w��:j@��7�ż�oo�N�,��|���pc*;�\��tl
jq�*�͈�/H�������e�ҕ����h�Z�y4�qC�{&rsFP�!�s�:�,HvY��H/��$���k��=��7RL�~S9I��r����sM�����$���
x�ӌÏe��U֭���7h"�Ds�(ޡ!,X4�6��@vX�=�����rE����{�xp��!pX ���(�խ���XH�c��y|�T^�@XKr��]aEE�g2�ڜ
q���mY��C#Szx���sܰ�ݍO�K'����.{"�M��4�2/�wȆ�0C�%�䬘��:-UJ�&�TNu�x��Bϳ�ڬ�g��|��}�k���;Y���|��ǩď�Ը�1�i;<"��KB8`C�-F�8�ڷ"�7�R���E]��d�v�e�E�waO�B9�W}z���NSo�&�G*T�����Qtb���CL�W�uu F/s5.��]]ֺ��rm�]r��ݝͨ܂���rr:�Wh��K�����o}'D���'b�MngZ[ͤR�:��G9��]`�c!T5V�K�Ք��R���tգr��]�v��k+r�}��T	���d'C+0d�:J�ص�/\2�H0�������j9�Ft�\�����fU�<P�y�Xm�M>u{o#��f;y\"���E����U��\��RoTj��^�7�dq�Wz�	g|3���-��$�w��	&�q�ןK����8��&K=[�Z�� CI�A��3}��a�&z�-2*8o4�Z�:�	���!پ�ZSk	uF���W��O�����O�������v�v���-B��v�
�q ����:���	�sZ5vT��"D�z��.r�n�w�+2�0>��!����;���e�[�ꈚ��/�Y6HT�Sݕ�lxz���S	=��>��\�;�f��ce�
�ǥj���NSg[H���5Wdo:�>�"ZX���M;��1���)1G�W��g��K�S�31 ��w=���v�k�qtN�fι�N��}��ѵ��n,����a������}ڌ�7�7��Q���v�L���$���B�gc��`�ي��B�@)�����Un�Ftu*�lQ =��9�7&���b��mgi@S�OOq���F�Pu�;��s���n���r�jV�r���MRV�橰��.]�kU��|�<������|�G.q:�k&dz��b|�.ܶ���F���dW-N.�T�T��+[�{]�+A����fc+�^&c�fu�{�o�26M���}��^7(�r�O��ʹ,]���d�F�J�h����f��n*��B�je��D�D�ݰ���ҁN����`+4f;t��ՙ� =�C��b{α)��^�OT4�U�}HS��7��g��֬V��F�vn����uv��Ω$�i�j�)���_R��X�շqǖy�޾�2�\��1��Օ��^�Gc)#W)ӑ���g��2Flh��z�gSyr�,.�vmm��R7�47����VE#ȾՎ�C4�k�]�ިX�ڑD��N��Ƕ����I���1�s5�d�D,����|�s{LR\�gwm!�J�&3it��0��S&�엲D�qU(T�:������;{)��Z��ѯ���%y��\��7w#<��y��s��Yx�0NZ�ب$����AtZ����^��Yܯ��ܗ��j�3�e�v]�.��R� ck�M
%ؓ4�s{bh��I�5�V"��r�h��דv�#��.���m�LskS�}�I^L��{�Ni���*NlG�Ĝ]��9�_3�x$�2�"�Q�T�c�ٍ-%)1Y�UM5�W��TCE:̈"��	���,�b
��}eE���YSS5F�Q����}&PAo�A��0fc1T;�����`jj�̵�I�eV�mdQED��Q��ʊ"&�֍Q��RALEF��ӵA�dQ��b��DTLA�:���h�����f����m�ժ �-k"7��(��30��"���|��d�NNm�"b!#,"L̬�"�3|QTEUZ���2ʜ���(�Ă�)�"�
���V3\���򧸟�/��yQ2�i}(=9�g��"-�'2Ե��-S㊶��0�}e��͝z�yQ������i���JYtj���G�S.�S���~���?�r������*���SB:S����p��Oо�G����/�o��a;ݚқ@���'��rg*�;����(�$3q��K�fUa���u.7���Q�-Ⱦ��ӮI7϶�,��
����#:y*��˵U���+l �,��~1�6��64M��m�P�V�.֮A��IH���Fj�S51�
�Ae^����%-� �����}V��˸�gS�AF.��CZ���p'�a��kᏺ��=1�����uC;T�aEN^`��9:}+Ks��3fv�d@����U���[N�<�"�:�s纳���Ò�.�?X����=�Z�7Ԭt���3��B���z<K�;�K�c�Y�7	�=�)(�X�[mP~S
k϶�U]�ǜe{3=UM� ���egl��� B�-�9�:y\G&�o\|�t0_jzY�Ue4���W��r/��I렣[+�"�I���N[Q�Rɍ_ZLfX���9�#k�F�����40�,(ެ�\�k�� ���+c�<L'3��KO;I�j�����)���eߍ�s�U��f��Cݎx	\�c��D���z�*x�� ߙXguc��1��!Ũ��zϘ�d�l/����m�j�5���?����hp���	��*�DeZe��5�1mm� �\~�GL�
�M��w:�&&���O��̓�Knh�����X���2�;��ή]�[��y�B/n�[���L��㓘�wq���I��G {�]啾��<|M�Rrs{��q�$��Vq&b2eˊ���^��XfZ͢adɍ�3|S���%�ھ������׷�+��1������$�6]�";��b��3�6�0��*�WgkL���x�3���!xvU�͸�N���ڼ�-�f߉g=���2
[�Zm�s����!1Y���ɧ�]#�ѱ���,Vi�[�m�xAל�<��$��:N���o/��1Yˀ�	nC�"��OrF�5��N���Mm��{ѩ�6"��)�E_4�u@rY��B��'��%��Y���^�͛��7n�� .���W4%fζYY�n�����Ҧܵ��@R귔ɻ�2��jn|:ĕx���@�4�:�%E�O5�w�*ѐ�ڇ�]�E�Q���Ʀ��h����
Y�W9����:d��}���>����7^����ϓR�S�p:��z���pC�4m�2=˾���=�<ǒ�rY�d<��)Ĕ/R�泛���^yǞ���I��������������Ԝ�y#�oqd�G�=Gn؏�;{������@�~��=�oz���=ZB���xw���Fw:6���_#g|Ne�S���w���bH��`}�۬^�h\��!߫o<�}�۟y�κ��z���S޳�r�%��#ܽZ����یl�6��r�S�1�W�69�<�� {���㮼�}�����}�CyN����_]u����m!B��;�%�Cl��^���ԉ�m��z������ ��<��s�����}���7��2S���S��� <�^��i_$߽�� y�֖�����ܽK�o��M`mom���z�[y�{Ǩdm)�y̮NA�q�7ùO$6��B��J���4mu��\���s�-/R3LD9�l�����6���}�C�z>U��ۜCx�x]��a�W#��D����� ߼ �_9�]B�D@������T����^�l���c�zf=�����'�<m����)��\����{���1ԅ�u���/p�!��@]��w߾���w�;�����#��!2��X�8�Rܹ�G	�� �%;yoz��l�_Qh�Rx�$*e�pt�!6^L?�r�	�x;�|5� s6�W0�7���e]뮻��՞�
{���H��b<]�m�!�{;�����R�˱�/{)��wRd��n0�^�v�l��-�>̻�����A�xϼG���'�2�ߞl/2���d���w�d6s�x����L�:%;�s��
4o�S��*�Qu��pn>�1��َ�>[��{�R�/���/��Ż��l/2�@�ئ��by�������c�Ό�����(c��������'#Ӽ�M���/ro�=��̏2ýԽ>b�+�����	�`s9���J��s��߾q�q�}�x)���R��=K��b��ܞǷ2�S�<\���+���'1���d|��3��N|�}�n���:���P�$(�P�2\���<��N�;��}��O%�N�è_%ۼ���y�%�N�y������:��sy�\��>��������d�m�/2p�x���N�P`{/���Ծ��'���y��/��C�m��۫6�oz��=��{�]�i|�8�޼Й����4�C�=���5�'VB�;o��>��R�õ�	�����ώl��/������1�=�똇�ݰR���������;�$)w:�;��{��b>K�m�'�H2�c�=>�gö$|�N��O7�N>��y��L�8�ù`6�ԧ���)�K��y(q��B���w&K̆�b�/�����/S�g�Xf�j��ߎ�t;p��HQ���<O�8?g�ã4����{������U\U~[��B'�7���I��9n7zR��*�M��j�eVG}Z��`�~����H�9�=�T.�x�ޱJ�Sx���_ew��P'RPw)��� w��^���}.FB�/6�s�޽����^m�~��G��K�zk���v���N0%5�{+��k�D���N�7;Ġ�]`�=��~i��v����y��y�ƽ\����������������A�r{!��S����\��+S�b=TFO�O�&}�^�7ɀ����<��~q���n��弮��-���wJ��È�G�z��N��v��:����}����|�޹�{�ק���`m'R�/���s�;+���Ɨ!|���w���#��9�:�ѶNЇ�����=��{�|k�x�n��8�C�7�!u�FJ{�!�\C��!Ľ���^ 8��P��\`�Hh�{��26�6�;ws�Y��|������ޱz�����|�`��hC��^��}���n!�� =��c�{�^d<���u)��C���ۮ��}��={����6��l�!���Od)��{���W�;:ù|���C�w���z���^_�����Jc���P/!�T�O��>��{�(Q�/0w<m�{���R�`�'��&�b�K�{���I�y/p��{�"c��.���s?��˾�z2c��ԥ���`��Ԇ�a��d�͒u/1���y/�o�)ܽɶ�{�=u�\{�k���[��[y�Yz�����mg��֊�����b޽���J�
[�P���v�l��UxZ� z[R���T�٭*^m�+*v#��#�B�Ur}�����d�s\��#��7��|�k�uW0�y�����^cc�����}�!9���d83��op;����z�����:����;w�o[�ӏDt�>�_I������!�vǘ�3���܁�Zҙ��{� `�ԄJ�q��'s�9��_}Tz9Z�!�,q>�ɘ�}P>ý������%�<���� 5.�z�y��dR�����3�s��0�١�`�~�q�)��c�=��1^�m�<��Ng�]�`�S~l<��Cc�gi�����Z������m�rh�Xf���u�G�Ò�/�����m�#����B���C�0;q���ls�{+���5�%��N�`=��xs������o<�y�λ����ʹ99#�qix���5��0�m퀝Ʒ����7x�<����.NA�p%x����:۫5���6�\m�>u���H�)I���΍�z���rW�C�-/V�k��#slS�M;`mylbǰ;o�Hk���ýq���]�/p���ԧp�y�w!I����u�~l�z�6�{�:���CNbw+��}�Gz�:c���}�v�-b������S���d���\��)�1�%�2M��|��|�R�K����w���@����\��5���|��MH�F�x�8��N�!w��9�7�s�p�9)�x���q�`@w����󾇛P���;}�&���Y�H��6T�|����V��1/�O0sz�J5ͮ���o2�3��s��-�΋	GѰ�Y];+���S:9�l�?å�[�p6	�wY���s`��G�|tُ�G�}����_'#n0O$u��;�op �S�d�N��]�y�^d{���_'�=΢"Ǻd*�w7ʭ= �&q�=���l�=��9��1�@�G����s�짐�w!GF��2y'1��D��>���xG�+�t�Vp���D��^��_��/r����Sg�N� x�n�N'i� 9��?C�]��B����z�����Ns��۽w�[��<{��zys+ܜ�r�#����s/��� y��!)9��8��d+�^��<6�N�m��=NHu�پ{�Y�{ל�߽z�2�s=Jy�G�'1�<\��u+ܻ��/�{h�(iN$���9���W�:��\�\�mdf��y��s��W��X��̧0u/��o�pv�2=˨/!y;�y�%�����2np��z:}�k�2�5�Q�{�}�E{�o<A��s�'r��)A��ԝs�y#������/1�q�؏�;�pfo�o�g�k�:뎹���z�@��-!C���/��	���J�o�̾�s>@{�Ru�C�c��u��m�k���n6=5��Y老�}�>ߢ�X~�2�����[��iw�]��u�뭬|�\���]�&�8�\I����l5Gm�kL�8+1�ͫ�K$��^�\2N�k�Ԏ�Աx,���� Q���o�!�����QKr�N��9Z�����h�t�r�%J{X�Ļ�ɼ�x���UW�{m�w�4k�CE5H\� e��Y!y��Tm�8�Dtc6�T4����Â��.�ObFc��E�f+�5ʝ�8Uyr*D���׌�jc'8΂u��= Fb�y�����(�<�7��8Dz��������-X���Xٵ�{[n�,�7|y�6�=�5�΁���j	ݘ���$��v��`�I�c6��u3��u�Tj��{Ĭ�p��5Q���r��՛�=t�8�K5&�%������n�xӫ;���¢���%�.H��{��\2��%~����SH7���6#cXۛk���;��7&�Y�^�:���!��=|��!�}e����4�Jfn��y{J�]���i��\�k���N�K"�+���p���*f6�]�o�磌�;�6Ț��t\�<��p��w��&)�������)�;�~��Kқ�*ě�}��O)�'
у����̻n�N0�c<
9��}/���<���[�'��:��"O����9EG �"v�b���X�N���|�Ĉ'�4M��*�w�-�L���w��Ae��u�f��"a7=����	7�����K7q矰�E��֎�[�}�$U�������Mk"M��<��2�k��F��:��/;eY͍{�{t8,e
���M� ��P��(:Z{����X����>��́���#E��M�聉O�f���q�kO�;օ�*ҬAo_^�N�9��&�΃.s�%)N.�wnT�˩
��M��)�*h��8�j%3����2E�/n�Ԣ�Y��ǻ�%7y�̶��f<��EQ�A�wf��867{�I��\w@�ĸ�Iu�Jb�E�#�oۘ9a���n
=3�fK�,A��7��f�ӝ]B�{|<���y��{�U#�о�:�t�w}�0�(�.��ߤ�L��c~�^mH9��k�·h�X5mǋog!5�0q���,�j�
��_yZE�K���i�
�ge����DÑ[��ju���m��X�>%��+=[�]g�ձ��6♄D[���]��!�3�~����G��E-��u:d��m�t�%�+��}o�
LSh\�n���3)\�Րh�CN+�8&[}ׅ����{Y7R�-�w�gu������lJDJ,b������Zaf;e�خ����FA���ͳ��L�47���8�=�2�ɟ	v8�dޗ�v�D�W���?� 5u�_�����5l�#����h�"v�V�(4�O��ma�i�Z�yQ��{iL��[�<^T�Kw�CyJ�;��#
	�t�Z�����:��a-�h�˅�]Rη�n5��g��3�:��m��\�Qfn�|z�����Ʒ0�6��
���DU󫷐�B�]�gkx�L=�J`K�y����p�{s[͚,	��!�&5''Ǜ��Zz��=ӂ}F�D��X�'	�b��=�>eކ��ls-O��o��nW>� �}L�W3���}�e�a�
<��#�LY��ݚU���)j�Z�HV�/�ذMX��>�)�٥���BI��8p��8pи[N��Fwm���T��XW�G��B�ٓq"��;���ڏu�)c�F(d㨬T�g	{�Պԭ�E�;�����gD�?��o\̘Gk<�M?MX
`�S�E2шtٴ�1�>�����HZ�>��m6V&�jkD��~�?h��a4�,�Xe�2����2j�.�ȡ�h� ������'l1�¢��#	����(�s�02�p�ɠ��q���&j���
����V4�E�w��U�DS$�U%QV�)���Ū�*��
���1�"(������eU�dӵ�3T�DD��# ��0�(� �1��3#l¨���fjMXEVNTTE���(��d��&*�d����jsFURM�b���*�h���"R�XcjM�[������U�8wv������y(4�p��x�\^�%�`NG�9�+]%jM�'�X�Uu����G�%x����j�w�Dwο�
����/�c���	f)��ظz�/�p��<�cY���V�[R�_��8��Q��U�1W�g�Bo�(��M��z��%3�6����H]	(��:�܈�A���%�����Ix���ؒ�'��w,ba��q���C賌9��}_!e�o���(Onw0�Q�܁z��k�G������j��P%5�'\c�u����.<�ςv�9�������[1�ў���b6�N�qϮj�%Y[n���w��R����tnJ�t�^��y ~��BB���Dxyؙ�Z�0�Q�ws�Õf t1g��2VE�ٹ8ghmP�j���ݧ�h���=�a��kڼha[.�9�/�1d�tP��FmUꂍ�&�uDΒ�Mr_�{���ii�8A0�����l@��݋v�cW],,y�%�QM8b\m8�
�X���&�l(h��ã{�[�{wءuv�f,{q�lv-�N)�c���oq��&JXV���<]5W�����u'��ȍ5t��+4��me�Y�@�)&f�/� ���I����9_���5�Z%QG !��/����mߧ��Qj*�	UY�j�YX'1�-\jz6�*k"zy�%����ocm���|�}�ٰ��\��rM{tE[5֢��w	Q�Wd��|��7����!j���[��{:�p[P`�>���W;��|�k��K+��Їv�+do%4d���l݈N�Qա�ܸߣ >)�=�zNF���vQy��[1���,��!��J��Yn�_�UW�W�/)�+�w�s�+��%����5�Xw�R��$8Y5�Ԇ�A��&�w��U�8�;�&��)�U�N��+2���n�ؾ|]�y͉R�,�W��6Ň�$�WDٸ�3�$;�ꌽ���K\)xx$�)��'$V�V���(�Ր������H�~w��>iɝ(��>���-�9�˸[�/sv/��غ�|dr�v��}p�@Ʉ��4m���̀����ۇ-s�̡)*��e��3}"��q}:-ͤ1F=5 ��YN׭��|ޞ�S!�V.W����\���1\�i�0��p��׺��ۣ�VT��c/�	ݑ�n��٭��hU=��S�*�G8���'# /m���4���
&��6L�mwC�]*>��u�ZB��V&�k+W�G��E���[y��9=`�^?�6�.�R��ڛ����ļ[�)�Y〾�B5�H�N`V�J�֦�Qѝ�-ը��&��x��G�6��\O�gy�y�Ȇ��WK�e=؎J�#�T9;���4Z��7n!�f�9��\'pC1ɤc&�5��)�ڳ֘R )�OT*��9�bzIt��L�᮶�6��6�Ai��9����@��y����9\.9q8�9���]�G��i�w��i%	e���ǣ#k!5�5B	a�$��]�f�4;��b2eF��N)��f��y�:��9]A�z���>�uh�iZ��=b�[��o�zK}�)\"�'�/��m��(F��+�𙴳����R�.E╅T��=�z9����ٜ�j(s�a�|�wmK�����������RiF����Ð m�ͣ�h�˼Q�e�/�\��h��%$�Y�^�����#yMk8(�RDKɅvX	T�C6�D!{���׼"���;-�ݚ�Uߴ����6����y���[1S�=��kb�Y�'`��A�C�=�,������!��5�r"���7���n6
�kA�ʝ[�3{p�%��?:'"Xyj��z���p�'X$��v;d��@ag.�R�ؔ����KOjae�%���V��=B���.8�Cbf��R�h ʠ䡻�u{�+$�q�w��qR�(3�������3��~]��"$$�%q]�L�u�XsnGᄙ��E�]��a�gg�rJ-A�ec�Z�e�Q9����j_$��Ch<5k��Z���n��e��Ϫ���yb�&|+�Α�'{U�#�U$n`�雧g2Jo�<�-w�K���3dt^Ď�L��GNx7���H�Q�@��Kb��W�ϼ�z*&������s��L~9�� jS�ryv�溌33]B*��n��j5�7
,�'��Evm
�%�笂�m���}�^�κqZÏ�4"l͞����e�{�2;n�05�! ��^A�U�k2t���g{~O��O�J��w�򸙸)n-(�8���q�54��O���zj�\=w��f��mFge�mK�;�q���u�p�ms�0�\�ڪ�û)�g2,Q���2e=��<�< }��k��I�s;ME�Z���y�j�uv4oW<鑽�4��<��)�b�	��ꫵ���&�S��3(֒NM�_z"#��u=H$�����0�5�/���q�!j,��x�-���p:/S��Md��$�� ����$�c��';I��(F�J�zc�K��k�b��n�Z�NN�S�6/v�+�_mL닀i!r�/=ݞ�����c����F�͝A[�˽�Т�n4�
�
p{x�v��s��
K�3V�-.K*Bt��dL�[g�5͹���7����$�⬎�JS]j28�\��/�s�8-!xy��+�FC/d��9�'Sۊ�.Lg~��I�Ԛ4��qS��NE^��ޜ�����炖�A�֒���(MHtR�o''Q��۶��6���%3��ߵ�6J{�b��sf��d���d�8��On'�ŕ5�2����&�{�:w�Uqk��JUV4��G�Gu�m�d�}]ZD�v�W����Y�?yt\j��v`DZ��W�vv�fܴ������ȇ�	�Ǻ
S�2����H�zL]zӑ�A�OF��sO�!�Z�:���:δ� �b��Z���EFr�q��0^BOp��1����D��И։{c+K�ζt�DsЈ�' ���.���H���j�_�#��ߛ��iծ���A��@�>�"��n��>s��&�o�6p�d�m����uƎ�P�h�.�<�!�3������$�=�zx��R��D�
�I�m���{i�E�r����].�+�W]j�O9>�ޗ�ӂ��R>��]O@����c��dz"���[�p���MN��˕�KR��)u)n)SB3�J+nt+��[g����zu��7�C�x%rF ��L%���Q���AT���k��K%ڝ�:�+jQr�F��7����?��͒	(��5�1��Fײ5�T ��N�c��V5b|��/}\�?mcG��g&��� �(>��o)mK���k}N�7V��iR�3r,ղ�t�C��Z�	@�£z����ћr1�)��yWS]<��K[�(4�Ġ�/�WD������^�<��$i�uw�M�Ks�M��;:��WC��;��R��3��7�A�o����OeT�͸�؆�Щ�f6�ypj1�_iU�_�)Θ��0��u'b�U����~�pN�tyQ���{��.%�!�Z�QܱM�0�8�
Xc9K����䮅z���������+B�69v��w&��mV�fu)Ѕn]"�k����G�o0��'�>Gn���*�Hyj�e��̩ר�<��R�8)ߴ�b�R�<�ĥ3�:]ҠEd耒C�2�7�_����)�.狄�3�3���꯾���-��w�z-+��dЩ�q��⇸7A%]���\|�Mv��`�ρ�k �)2��6�Il\���VRw�U���;���ջ����%�zE'xNǔ�� gY�5;��f(�8�m5��\�C��. U���y��]Zj���힬�U@���f�� ^�vm/1��^��9T�pp�8��Z�j(¨EZÛX~�ԥR��GRw^���|�1��Y]W|,��3ɞ6ӛo�F]émn���A*�^�}+��G<�l�Yӊ����J�s�aCתg���X���G�1��(��x�Fs���&�ݥk1>��P�JG;��<f˘l!�8[�L�w�y�nc�`00�1��,���*i��Vj��^8�H�u�O�`	�m��,�ܭ�UQ��!������������^�V4"�R�i�ٍVa���T�X�E8e�`a�����)��b��,���o^h�m�����^��]9�ֲ�Y	��[�vv`�縰a<4TkV�y���f-߅��LN�秲��G*p�(O�@+�u]s�U*�*�sϱ��"�Vm�$����)%+��S[�>�$
�s��;O ������Hi���j^�E���,��+WQng7��2�STT0Ҧ�n�Ӕ�)]��y����) .�,����z�<���U�Y�(K�a{i��w>��y]� R�;�I�Н6�YN�|&���]���oQ�]�Vՙ�A`e\&��C4Y���(聹�a������X����!V$�X��I���ֆ�!ݻ.�}As�Wo>&7��n̮�;�i��6 ��)�t�G7f�NE��SՉ�}{qiV{�4�C��L&�Vк��w������M��On5{�|�t�i�lU�T�-ʔxd�f���!�(���wIB����̥��J�	�̈7̛к�k�^Sp�+d�t��n]��5�3�;ۤ�8�mJ-��;\0=:�W�
�m��BFX�F�S��&�o���:�U�U�e��AmW.��Ń5%��=Ӥ1�:�Ի!���Z�2-�f��t$�x�jt���	���mZf�OLUHJ�
�ӹk�ʹYɩב���A,7��i݃�ޝ�eѕ��UF�+f
�b�Ff%�5W*Fs�v@S�Lu70Y�-�'��y��� 9p���&��Iޙn�,D�վ�1̧�p��dF���{d�Y1�%iJj�^���k{��q����O�b&&}33UEITU�dDѐd�>�eMd�k5�&��f���{�ӶAR��eM�kXL��2������`��*� �aAME�Z��)��"���"�`dنKV�6�j�YYe�`DM9PPR��d9!TRS�1DQYJ-DِQ5IQTR%m#�-ALA@��SITQ��F�(

F��0
��$�3
��(��������
���߽���tlzo�:�c/�	�!�֩t@\����
�&���`JWUB�xG�ޏD{�4��ț�њ�r��+��8�C�g<Ux�ܠ*/=��Z)�T�3�%+�q�^������+�L���\�yb\3x���Dl���c�w����6��[(N�M�E���z��Bo;d�CU��LOtm�g�i�qÓx��X��'lm�O��bZ���V�^L0��|_^'���Md�� �*t�>m]�<�0�;u�Fl����>��f���Ûtf�A�Êc��Iېo΄��x�ׯx��ʥ�;66�fyNBs6�W�bઅ�jx�^���ۧ汛�5�UF�����k����O�'׳�"u�=�X�WO,�d׽���XY�Q�0�u�ңR���SÀK"���x*��hdS�⢔k���¾��T���zZ���֟D컛1��~UW�UT�9���PA�Eh ��σ~؎����u6���n5�`Д���YYWLҘ��1�LU�3Pq����PU�&�T{`�6�2QB6)���[�.�b]o����S��]<WaU)���.�j��@�R���'�wW����I�h3Z<4+���OU��$��{8'�﹢�_  Ty|��pC�e�0���v)kA�%��}Ԁ�j���f�쮪����^<�
�`u�v�s�KT�L\��4S���\��˃9�F �yjRbG�Keց,恵�}oRD"�A��pn�'�ژ݅}*rX��+���� ���{D\��B��)}Nf��k��lG;][ږ�ϰA��h�_I�f���m&�^
�p�]�`߭["��{�9YbA[�j���R�VÛ9ѧ�1vJ�X���>�ie��%��ږ4ڬ<�[�t`�;�����&Gh��b�ŹB�XV��46�n��$��������ԋ}s�'�U�&�b��{p2���7vL��؃��#'.�#0SX-��x״�p�
��n�*�H��!-S��jVi:�ĕ�3wu���<��B��U�1ַ�`D���~z�2��l��k�C�r���b}pxb��s�塺?p;ȅ��!P�3J�7�>;V�r&���?|Τ:��ˆz��x��.��=��s5�H�k�jKv||�O{�KX�U�]/��1\>ţQJsή^��-<�Y]�=Lq(�)��# ��.*�h3L/Ǆ�j������1b1Z�<�(�� jܪ����Z���K�0���^��B�E�˵A�R'e��7�S-�y*��
ah�^[|)S5�l�;V]o�﷯�}���*�U��Q�HM�n��j�Ʀ��R�e�2z�A"���g3�O.����W	rQ��&�oS�b�K9�`���x^�F�yv�x�[�*	�VbL{yj�o;p\R�4��aq�E�[���J[64s��_}_UU���z�%�4����8Q؀���T�BnGmԬ��m�1#�'���WV���u�y��y*b'4��k��l�(�����z]
 OW���值T~��	yh�x`��V�������V�>��������'ѓSw[U��U��*x�V��5���z�a\�y9�c�$��;p':��Xž�&�s�5񊷮��I���hc�k��=��a�f�
���t��R�X���˗R��:��8+׬BꟅ)��\�s���%P�[�&�4��4���6e���Ow�Sҥ��V��pA�=y��}�ʱ�"��u��v/���M���#��<h�i����Y5l��o*"u��A'�K	�8����jff�;rv���j��k�BE\�r{i�7�p�="R+�����N��c^����m㥴K�ea;ns�s��Mh:%�	�7�����r��c��v�^N�n�o���E�:49�y��u��TU5�}�{ސ�i�N�G�Bb�s�Z��������xpuf��᜚t'�����&�b�P��m�ϹW�K�Z3O��^
�>�m��������z)P"�<4<h�7� T�5��k/���hqG��{i����X9��O*+<��8t��Ld� �CżB:gbT�Sꊋ�u�-�2�w�@�\p��5]��s|�w�A�c�#|j�����-
�`�du�^�쥒X����jw��$�3����UK1��_;�`�gֈV��zm�j1��/�t�o��ƺ]{�+��VyP®���X�!�oVv�m.�p/g�[�%Td��"r�n����Hc���D֊��{`�`�Ҟ�߮fW���]pd61N�V�#��q��W.�"�z筤}�8my_n�m;���庭1�x.��^��Ia����sؽ�X�CV?SJ��zJ�`��	��'��fu�|6��[qq���a�� ��Q]a�y��W�W�V�ڎ�3;Bz��l�dÓ���&��[�0��T�*��Y��{:f�� x.���$lJ�W������v���@St�I $���m\X�����d@(h���g�Pm�.ޥ�hv�����;ǐ�/�������3Q���+)���^��{Mn�+�P?.�X4p�PA�����ISAܮ�zNN�j�@#��e�@�|P�jJ:�"�+�����:{�p�k�Y�Ժ�F���W����x�+�0���l�ky7љR_���Lt��|j���qT4��x�09������t�vfKn�-2��/��*�Q���,1٪�o.,��{�1L?Ge���Nm�v3avWT���/�x�T*с�7��D�U���[q6up��z�-�EP���c���'}ȷ���-stz�=���cn>:ѡˮ|��g:v��NY��\1)M˼=d�Cs�Pa�,/������d�T��q�]L��2g$s��
�G��VUG<�4e��;�1��NC�
�x�����(��]���HP2�V�>Ofr�;)��\�S5*�3q^�\.�}��S4��v�۞87�碆I 1 �h�q�:��əz����cGp,xu��5z<HCo��{��妽Q*�Ʉ�u��G#[tfd�pg#h�ld<��.N�v4&�`dU��S
̭\8 ��l�$�Չƭ�l��=	��re$��X�*sٮ�
�6 �K�`D���~z�1�s8��<�f��[�����S����;��;]M�u>L�oT�W"��}�*#�5����@�{�p�Zk��:̿���jD-�8�"�ٺE��F�L�Ʉ=�O���X �F�\�����w�T.ʝ[���)Pb"��[���0�<��N���*!�:.gNy��eI}6Ϊy��C*)X�+rj�΂��ڬKR�x���(`����Q[�oi���XE����z#�X�$�3�>Y`,�F��H�A�C4�|8IA(][W>Պ�X�&�y�0'�FQ��r�J�RՃ��\*�g��� �{��ؒ� ۋ�5�$ĉf�U��cN�mB�Jah�^_���A�Ϭrz���^l�d8|4P��C��J���
?K��u���N�uő���=;w�]���ph#���^ձ�2��áІ�Z#��H�s�{�wvԸ@�g�x*�w^*m��W�� �s�<;�>��M����/O;�y~B��+"a��r��[4�K��(y��۠����c�
�>�;���"��xS�P�&�a���@w܉Rn����]>7�
�־��а:�Do% ud�[��6+{2�"��%R_��J�*��L�:
V�v�RB_��\�o=�"�����0�cSry��!�sʛ]�7u}݁��(뷵}�=��2z	t�0��q����2�z�$�6���%S��:S�6 Ѷf�ޱ�f6y�`�p����Q�/xd��nN�إNk�8�8VBW�ȓuUO &��1>S\�\��}�U��]�'WK��1N�+���ea7��G�S �ӄ{����4`�諙���+^"%�Fmm`PK2y^���79q�R��  �xBx{�j��֌pxH��W=9M�3�>��k�&ﲣ.���Y2�c��')<���׋Ã�40ܿx�~���\Q�qPdD�Ũ�,Q���,����o}�^�QWx�<��	�y�Q1xU�"(��� � T�5�]�߲wJʗk��ו\7�ߕ �r������@pUӚ��>�wwq�����Y�S�l�R�[,R�*,]��g�o¸��%Ҵ�n߾E©2ϕz��p�჆�����+�nO>c��y��ؼl��Z�.�(�i�՗Vhp<5�p��@�腻�W3���t =,r��D؍�ڼ�������75��]G���GJ�琾7+��rm�����������;��������mPS>�p&Pѐ�ܩ[��E�,<��e8��Wc*,pႡ��Q�+�rT&U�K�>��8��A5�W��&^ؔ(ɐ]����r�n=���Gf�rVTJ�-��Q��\J���]s�[�n�b
�<�����␷�{�ׄ��s��z�������EMt��Y��c ��r�����S�V;cR(�n
�� BD���!	�~�=��n��\����'6�"��9
�<�y�����yA��^`q�g�B"I�d�z=T=��KyԺk|jC@V��杺T�/��<)���o>�<�!8�����Z�����6�v#��])���S��-�l���WV����YD�~(s�PrQ�|B��r$��o;�R4-�2�6�K&�W��qQu6�L��`qd��Ŭ����`�)���*fؽ:{�Y��5�R��ͦ��ӈ�+����]��=L�g�����-��wVi��C���RTA_��>�إ9��f����F�k�.�/�vfn
k�G�F�e�l
�̩�M��=���UŻ�}|�k���7��޺7I�:�QB��C�mÐV���h˻P��)�ܝp*�v��M�7����e]s!b��{.+K*@��m��=�t���%�������X��U|���}W��a��]�2|��Z#��[�|���9�ۘ+yҬ�gI`SV�ط���E���j�v޽G�kDm�t��J����ed��-N:�t*�erx�ݦ9Q���;Lt��X�iu�0H�X܍F���y{�u��I:Лӗ�}Xph�(n��R�}u%���`i^L����p5˾��T��+s8�%�gn�|"���itm�4t�M�;1�6iGg���R�*����Z/�N����n�9NWu7���$��c���J��Ƕ�{K�+:�\���޹M��v�i�:�#r��y0QQn.pU㬙�^ҙ���4�N��aRJZ@�5��Nťa*�z�̗٣e��q7rl�jVZܻ��3h�p.�vw#P-�-��Q��|�̴�.����Ԣfr�q!Is8����̽Q.�,�r���w�����(N0�y[����[V������� 㫍><<dn���K[;�)5�^�4u4���ǔ��/��ef�Ŏ���(2�f3B��qa�zK�]t���78���gv̭�ob#�u
�����N#�8�y� a�ƶ^��GA��B&í�*N���@�gv6��v��3cI�㺖�ʿ�8;�*���A��طl�^u��X��)̢uI���̠8��[Q#��'!�9��a#cnWv��7�a��b�Ǹ�$pQ�@_er�;r�OC���g��.L�մq�6"r3٨�n�2�U-JA�h���hj��J��L����%i��J"+�r�b��
����)i��


�����7�di�� �
�P�EMfb4�KQ%P�E�4U�k#LP�ETm�V�ȥ�����(j�&�����"�6�B��K�U!�T4�ِQBѪ�̡̱2�",���
$v�Z�����`���,��2&3
6�IF�ʃ0�)�
)s# �(*���$�P�+�'n?��u�D)c�~а� _ou1�FR�k��v�o�Mfػ����'bʹ����DN_.)5*��	��i٨Ժ��L��^���]5P毦Uc˩�� �3�%����nE0����i@��t��~5p�r�@c*���㉐�v�̳S�̎:�>z�о<���p(�h�(:e��1�;[��A]�������t�җ&!���F�J����T*у^eG�=�7�IjvtVOuFK�n\�5�1�{�\#
�T�s��9C!wT�ɶ[�E"xxU���SI<��
�僧!��@���T�挗�8�0Ӫ�UBcb�t�g�kxfG*[LR�ݹ�ȃNJ>׻���-���UV��d�. ���!0�ؽ�·2C�yl��+\��~ �פe�{)��� .��v`���j�N�9��t�����]&%��vn�G�?es����-����<���5����s��8�=�>`���l��^�}X��皭�4�"�,����#�T�{�����Op�씻Zh��k)͗x:kdi�jP�wkF��W}�y՝`~DD{9�m����+rsl��ut*qL蘗Ά���|h���Y�<|WD��+�;A�k=2�H��-Л�)�������Q�x	����Q�L*��U�������<*V�P�;�7,S���0�^��-��q���xX��N�1A���5��!�ˊ�S;�F�_/�wk�]��r�g���"xALgU��08��u�-�=�ݝ\ �=Z|:%S*[$Ҭ���Ճ�.a3�|+�CA�X�zw���|�X�h}G�B/w��d�]���h�8��WP>��{�M�{x*b��xP8�"���P@��� �l[��x��#�t�s��g:d7k�,��u
Z��t<(�l@*�p����p l�g�^Ľ8�=t4\�H�Xߐw�2�b���U�J�á͞�D���]������W"���e�W���
e��c�T�$+a_wZ�w�0���V��iQmd6id�Vf�}*5�^s�{(#�n��i1��fi��v5�ߪ��-���{E���.���XP��<5�K�FVAW��M����8�*�U�s�z,UXA��Ty@��S� ��8���Ii�|.;![}q��dV*���(�񊷮��F���x-n�n��V��%��n��H*��g!�R��{A^R�6(���h���1r��+\)K�*qӓ1�D�-�=,���ڹ��M�J�S�0%H&�ym�&�Y�|<�����*�P|��JI�Ț��wS|K���0�B��WD�8�:N���2��Q�f{7���ǙBo�{z� ��%%���̫6n^��PYGl]�ޏ�]*�G�qh�<*��N�Z�hZIy%�6�xp[�J�Yq6��6��j���;50�L�,���\.��T��f�Gp�¬/X�����T!�ۧg�'���6�n�-���e��V��톻{�2�m^��:�ѭr��[�㹝�]�}՘��QV�U�"=EQ��XYOOYLԖէ��!.O:t.f᾿�6e ���"(�Z@�4D�
��ܲ���\�ou1qz���C������m�P���*�9��s*cPA�fi��}8C�c�� 8-����hԦX�q�SP�M=b��Og�Lxp�|*[;���G]�eU�tK���P���l�ι�c�����P"ڲ桺{A���w��g��~#�Y�h���W�N���~��y��R�1c�'�Π�H\;G�S�s��;sw�����/�V�M0A�ʬ:������7	ۻ|(uf7���N��:򙚝շKc�NO;��f`܈�V��4R}s�%���أ&eR�u�5�N�F�5��F`Խs�v������j����~$_�N���`��[��U|��A�0��p�W�����6;ی��f�;i6��|]��>;��9R�oU�So�D(��9f�HH�Fu�#�{a���GJ�.�R� �s(+ɭ���侏g^h���J��e0�! 7���W;��dm���׫uy6�[?���;Ss�^��韷�]3�t����+)�8S˄V�>���LD�c0z�W���xX��-��[._U��O�}nN~�\��{gue��M�ay���7���p%�8T�:�W�n�~[7��ih0|E��ѫj�fb��B��<_ƀ�IZE(كU���ԑS1s
D�S�����j ud��ol�$��H���#����T�l� A�_;5�)�Xd�=�s�wU���,j�G|g�z��ϫzVӡ�\w�����N�����|+l����MA�QU���TƶFB��
�J��mT�<����obk��P1W��X�/� ì��
o�=�P_Y䄼�wκ�t�w��k�50S��j��G�k����*^�m�aˈk-��s8o&�4��bT��D#�(�|��S���G���f��)UX��^�e�����p�'D',U��ǀM.�]����{WZ29{��{ބ��z��^�&�0�&���k:;�u���֫~��������|=LK,H)<�w�:͋�BQˁyffo���/��-�$0N�zb�z����  �����ZIt��6y5�Zʻ�����u�{BT��U|z�굿�+&|��wU��i{`cy�Q�m�m+2�[��e9n��W��WS�i���9��ЌU.c'\���Ǘ�,����J���,�JR����A$L�kn,����j`�
��.�Y�(4?)���]8�K��	�Ų_��E�+��தNR�1uHh�i�f�'�ۿV�%�����%K�@�0z%R4I����L:=�%�g����O6�/�ӟf�G���dݶ��%ӽ(D�n,�)S����^�Z7	�UЙoG�Zi]�>��i����2���v��o�������2�^ .*���}�OC-�\�"
��k���i������k���Nw�et��rK|RJa��=7u�f��B�T��@!���H=�n�v)��q�^�ovR׾'��Y)��Af��P��k���*ݧQ�.{����=^�G?�� Vx�<n�`��;��;@aO���pM䧉�|Ǿ��������j�p4l��G��%RUF�I9��Z�M�Va�o����R��G�ª�E���Ay@�z�){��ԥ+*�Xi���,_LPz���q���־��а1D�U��+��Z����ZE{��ǇeE��j[�E���4�8*^�W�|�F�ҕ�qv���Ҧ]x1L*IW�z�7^<=K���~^ƦVBW�Ȝ��Kq�rz֦�Άv�z�>�s��hx�7D�>Ú|�|-����r��5�(%{��9��L��5t�g6�?�欹�m	׋؂Y��4+ 2�m�$�u21
5���=���QU�*��N�w�x9�)�۱��	R�j��]�����qO{�Sg��T�$B��#�0т���tk<ՓX�#C*�m��m�w�qב~<#�*�u�  �xBx{j�ʚр�oO=���;��U|�eFEј�+V��aW�n��h����j��$��CJ�Ux`"�ժ.u�����]���쭇��t<ot�jU��������|�|R���� ����]��&�����h��י�M�O��w�@N4s��U
��=��rf{�Xf��!Hd ?�l�4T��L1Y�T�D������o�opO�=��c���©Y�<����J��ű��)���=ꕵ͵5�ס~3���j��D|�j�S6�@v/���m�q��B��/�G�D����8`�wކ����f�A�Q��t��5�+�e�E����Ȼ{'
N�9U���%I��_E~�m�L��W�ua�%v%b�,ߣY"��W��G �æ-!8c2����AW��M��,��{m��{"f.c�/Nާ3�'��P@�*�����p��ٺ��� Ý3�P������� Z3��Sc�V�#��C�Z�^�Z
m,Fa�+z4A�Q���j����xK6$���TMb�=�I=��!AU�W7�� '�р6W$6Ҭ�;��dN�-�����ú�P\�:�M��UӕFf$J�;2�R����+&���6ƺ��8~ju֣��T�fa�W�=���u����YT%�8�F��`A#��e��ꅊ�8�o��Z{k�s��p�>E�+��a���0�>$K�@;���S�W�s�|���'yJ�)�c��g�!R;���D8�hq��Bx{xP]�x�~����P!�躩h�=@SA�%V��񭸉'�g� ��W����6���4����� �=h�ܶ���ˡu�R>�n��'�o���0������b��$6�ٸ=R����ǳ�ik�\�+��L�q�?��ʑ3:*U[+v4����s&eW�jԹ2�t�� ����[ S��na�55ʜ�0��j쮪����v��T���8E���Ғ��xP�v�G_��-�� cr��3��mC#��F���Sxz��Vz���A�����R:���p��X8g#�t�kK/vz ���i��O%��X�;�	w�P���nтp���.%C�K|[ٻ��8/ܴ|����,��{!ڛ�6�d�SG��Qݱ����NI��N�au��i��ԫE�	bŃ���j .�li��g���p��gc�
����kW�p� ,���*�c��V��'��}cA�|�K���r�2���d����1�kU�K4v��ڂ�����v<��O+����n}~<1M˖���c��Ӆsê	U8쟲��Q��L�f������Dmj7N�W˳�
+:;V��`���]u�&�WG�p�ܼH�b�Qe��x�p2H��8��=��(u�RaG��n�!���qΖM*�oVT~��xD��Y�:���v\]L����=\�P�3-$��u�/�Xp�LT�+0�u9�W՚b5�we]���lN0t[a.U�bm#�kş�kv˕�G���A*nPbvGf'�_#�O;)W>R���x��h��[��3��tm��{��}-oѩݻ����P�VTB���&�擩��,TB�ӛ�؎� ^��i����7��
:ço:0��ēJ�P�w\.��)�,�K��C\]g�\П-�.ø�B+�0��o�`��j�y\vf��O.��]^�����3��"m)�C92�X� ���I�Qٯ�zRve��D>�,���z�#} �6�[D9���Nq�����i��e���+P�Lk� S��un^L���1�5~8�|uב���b��ݮM蠬%���u�hQ���][a���ntv˦���Ӣ3-ܜ�=n�J̰ӕX�q���%��u�핔w�<�o�����>\�d���u
$��.C����dK3����7�L�����ڤB�緊R��'�*����A��AD��K���Σ�WGM	�,b�-��nHiJ�:��[��vλ�Nfږȧ���~��ʯs�aS����u�7�K[Sy�*4�,\�6��N�h(���3*��frN�I�u��L[�*:aֻs���|�6iw����+��pi��&�ߞK����OE"�*�Z�#����trO��5ȯ�zܽ(�]�,>���i�ll���߽�1��}Yx�Ay`:��I�AI�����ʉ��;�ƾ��S��pC��M@=����.̢���q,}�:��=��T�
�}����.kN#��0\Rl�k!BE��A�����n:��������C,��2�

�S�q��A�dfц��G+&#!���l��2ɦ�
�"��b))���������3��3(�-fjŌ�̥�&!�#,�	��Ͱv��*��l��2�$��(��%Ȧ$�+$��2s0(&iZF"H�ʵ&T��Ak(r)��,��$
�����]kiS%�dc�d9o!F�(p�hr�ԙ
Rda(d�Ӑ�9:�]B�Hju����V���L�_��!��`���7k]빜�=ð��(T<ŀ��;�mʮ�J�Ο߽
��m��S�;u7B�J��U���|¦���ǽ�Z��|
���5�$�GAwS&����ኯ��}f���5;�ì�6��]�\:��p�e�����3a]H��+��mfKWF٭��P!���ܩdKv���� W��0*�Ѻ��MmgiE��Ip��)R�C�����ͳ�=~DZ�3���ഁ���z�=h�\���u���0���1�t�edD���P��y V}.:C�F�os{Y^����_�yp�P릩����j#�?3.!�o��� FNP �:�8@��a�q*u�m�Z<M(y����J{�[���1,��zׇ�ٺ$����EEE�_�X<��������ħ��2�ձ0>��N{<Z�7B���["���57��%�k$���Q6�����FV�ݦ#�����\jp�k@|��B���a��	�z��w��%*i!z��{��Hu��4�4�ȣ���/
	S�J��]`�hoޏI�y̧�n`*S?FؘF��+��:�
��k����X#�S�����u�gLb����	n�d�4%���Pe��&1eU�ƃ[9��b�j],�O���}/�~^\ja��N�����{,����i��7&�wS� �Z8Bhx� L>��|j�::#,wg�I=�0�6i��kڑb!a��b��Kݗt��_MY
x��%�z:h���O:���T ��LK����^Ҽ�[�=�PC�8=$U�5<q#EJ;=h
�Iʤ`������'{77�^��(<>p�ʼ+�@P�[G�=Pq�\3�
�������{��	g���o���4O�
�@�
��.������킬h�
��k��8����g��h	���/��|�K�Y�G�^ɘpW�Z�\�ǭZ�+F�yMWZš2��{��+�X���GG҆hZtGÀ��"i�%o��#!	���·�
N�6���p"E�����M�w��X@C��B��=��l���)�[��YL�[��u��g������u�=�������#�Rg���g�:�\mm���i)+�*�6�5	���VD�n;+����SI�3��:4^�.n� VFܽ��=��{�I�7s�P&Q[jB��k�N�3q,-� rm��q[q7P�*�a��37�Z<�T9ʬ?j�8�k����wE���s"������f��K�r����
[�AV���"iCڼ&���"�^����4Cˇ���@~��{�$ҫ�;9����fV]lG+���pd�v��Un�ݛp@Q�k�h��6[��s�^��uΠ�*�P��M��F'@��������eK��:n�$7ؠ�/㫆8�ʔ�v����@S� ?k^o�xl�,
"�Z�g��}]�S{8Z��p_��y�{���>��k�_�nVSqk�K��W�pJߣ��u$���Y���O�V��i(���l_��g�P�<���ÿr��nx���u�_^��i��cB	9��ҥ9��$�y-f��FL8F릲�˻���8^%���P�a-�H�l�ʿ8�7���:��m�� ��Z�f���u�!♡�W�����%�`W<�sg�W㯕x!��r��P�A�D�Zj��C%��=����oVi%�k���>��J����6�/����eJ�/;�,0�d�����[/1p*�xW��8�*�{][�f��.����ry��*�8xSG��<͏xV�b��v�mx��s`#�cJ���޺*�s��l��%�]w��9O)]�NG+3�ژ��5[�UL6gvrF���e�tBxS���xp��L˸Rћ]؛�Im8Jܭv�۞9� 9V��d��<%��cGp.�|��,�Pu�ƺ^]\�;��[
�p�^�A@[��Y����Q�ux���(T���V]-T�����oO>m^����&0�������4��C9e�lNYF��_z/�����F������M.��i5��	b�Ń��]	M!�hEṙa\�2���S�x`WI�n�f�F����G��'N��L�8{�����tp����*�m쁙�r���ȡ0�g%�EG��*2����f^�s��ܹb�ߐ�ʝ�}�ޓ��U�D*�њU�=
��~���xV
�}���^�w���~j�U�����ND
������8�A~8����׹��ҧ�j���|��'��>�[ȍ��,��k5�:�NR�m�F�78����A5�a��2�U�A�jU�[$ҭ��]R�K�"�*kb���HȘSy]>R�]M_��g�(�P���'Q��un3ֳr{����a�X+��^-���C_�2d����x���H��qXH�,��4�t��9^������x!�����E,@�j�����.��x�T�J�Y@���է����k�:������v'q����p6~U^���w���j�0����/�������?L���+�f0&�/� �kg���s�#��0��84K�� ��b��D�O[�9���Q���TdI�g�˗;;1�}�VGT(�j*���}wz��sR�"Y����@t��ƞї:�Z'f!��7di�ߺ�����yՑ�|�����ukE*�U�ثî)B�����
���d�ʓ���8ڦO
�q �(pW7�;��[� �RV��cݼ(�=�3Z��`�8W�IV��	~<=�إNF�r�8Pɮ|����{�$��/W���Sȍt0kG3�㬀E=��:�T�RcL��!�7>"�n�5��툅�Dт�ފ�V��������]�����S��<���t�r�Yw^�� b�<��A�z�*�yd�QʃU	�%F>'�)PoL'��9�sV�ѻU�L���Q�bj��)6�]�����`�6�5I3�%m�;�v�.<���ԛ��@g�SL`����i�ʷ�#Qui�rܻ�*� 8E]�w���I]�]����Nƽ(ׄ�Em1h�ʸo� �؍��'{���U([$^�iT��>����� �8e<��֊�<�M���'!�i��M�'gBo�:��2r�����6�������@�����&�3���Y��:�3F�Ү{���S�[����l�v�G_ƪ�_U�C�W��ͭꓻ"D�/���;���'Oi3�]�T��#�p��u��2c�:O]P�0{������EX){�S�C�N�vd{��ŵ#����W�bૺ���6_Q��j
���U�Aj�o�5\���m9yG^@R��� �p�\3���1�yo�Yi<���:�<0ob�p�f5)ǖ�%��Ig/�K�� �[��"�:�������<��8��/��A�A��
`�@��Q��[ ��o,��Ѭ��j�z���sd�*���L|�❡ux��w�`��+zք�2Jx
�e��G�(x̪ΙFM�h���ʮ���M�r�����ʊ�~�hv��
����)0�0Q��-\ ��8�L
�u�4R�3��K�S=J̍�B�?5:�Q���_j�*���3#��s����[>t�V����x|3<�x�+��N\䉹��2���0�+�B�0&NΊB�&F���n�j_���r��7ft`��	�}ϋy��&뱐g��E@�'Fz�#��C�3C�-!��z�J1@�R�M&��D��'*�uj�BL	5Jxi�x����w{��5験���U�q�Nn��l������"���}���c(]����.[SZ�Ͱ��-�ډzG)���Oz�\�o�
j�!c�l;9�7V������F���_=�~��kw�Y�������`P�z��H;���#�	�=��`>;��%եsc�����l�ojU{eO�t�#��dF��u:��˃8kd<���B(䉿MC)��a�@���l��%���7K2���vT�4��S�+����ڽ�&���e�D'²�*���O��N�MN|��p»��[N�/|�Ϸ��R1SVg�N/SG*�ts�y'�gY�=��L�{�9Yc��+)�S��ٱd,W2�.kw������w�ȪM���j���5���� :C��1-��m&��T�F�T��]$Ժ�߫�\�emQ�m�E'��p�2����~�b�*'4j��=f����������;�.��7i�<�(����Yȅ��T+�^��x�|O��T�<��Y&�7�q-l)S�I�\\����Jr *��@�WO��g-R�/�[]��ڱt�yxӨL�bl��I�(J�f��~�ݳ�>��	C/���gd���D-���+r�EpSD�Lf�z1��U�E�|�9�T���k6ɥ��R����O�e�Rr�c~����G�*���:�@���^�\0���N>�;=�@?bi24�>��P�P-0*��K�l�[CYʓ���+���:���q��Ip�˳�2��E@���x(@�w��}}�6�M��H�k6�g��q/
B�g�ٱ:�ʼ��K�"o��d�o��+ռ���VO�����O_ZP���~7C����=�������A�~Ձ�4Gi�a5<phM*�0V�`��w����V%M����|;�Pxx1!�O���L������>�Q��w8�,K��2����v��`}J\��u�V"�Y�qTO[�^�L�����L/�-o���Wi���z*~=58�3�1o�uX�A)�����2v\�L�Y/��)8�zxM�x�S����U��9�n5�h��b�nnl�j*�H�Ey���cQV�$���Ybc����L�3UݩuP}c�{��98+<('To�F�G�Õ�)N۹�-i=Pu�P�Kb��c�+��ູ@t�B�;X�^�7 ��Ǎ�����]�ܧ|�9t��a3w{4U�f�`�T�S�`�Uۥ��cQ�e��w46�$^碥�?o���o�l�k�S�XCC7�<�X��fj�%�_u*ef�ȫ�_P��	n+K��u75�x�(���q��˕��<���ζ�+SZ{2������C�5���)oT�I2�t�N�tV^*5�Kd�lTɋ �L�T��v�o|�&�:�AN�t�e���W�`P%�	������Qh�$���ñXb��*dS2��M��W�Ň�d��Ƹ����Ek�f.S����ݼ�8%X`�f�SM�U�Hf� ս�#�,<�uF��Vu��!7�[�'Jw�Z\a��Lw
۷&SﷁyWSE�����r�r��j9X���D��!�].z��œM�3z��c��D�NKl�� j�7���k&#M�[�v�M��\��q�jƬ��At&�1: �f���z��Dfˏ�����j�:�d4k���4�c��S]бsU@0f���r�w_
'�×,Wɫv�<�&g3�t����	�9�%]E ���q5�������Ae(�v&+s0� ݼY�6�Z\Y10_m����t�g9�n\X1C�{�.�@(���CF���$�.�>�E	`WM�O%ն1V����<�9����$m<�����rtN�mBF�7}yP�K�f'v�d>�jd�a��;�����6��ՅH(+Tz=2&M΢l��X��g���c�-�}���t��um8�nۜ,�E��9*7N�h탯-��	E�&ޕm�#��y�3U�ro��+z7B7Z��+<�5��NK����_*���ۓab흳."�Gu�`�����JĜ�}�غ۝RL�����!U�@UTdRP4�%.]�:�De�B�D��؋���d���4��	FK�f�$CB&�ZƓ"��*&�k$��"K�TC���&fdNө��h������m��j ��C&�Pa��&FC�@jr��.FFf	�o�D)��aa�P4��k4�j�j�,��ME9�E)@Y�bS�P�ff���j�kmbDjU�}��}DVJv�]�cV�]M��VdVq,cz�h\_
COE�jXw�m��\��̻��P�'�N��z*��+�P�\J���M׏G/��rG	�
�$��{���S�:�p3�����F�<=B�p�֟-�d�>½�0*�`���a�s�^*����u+b!a� �z�����GV�Ή�s�F�V�:h�zyׯ�B� 6	�/Kb�;��O:0/yP�0px_ԍZ�?���"
�;=h
��(��OJaB|,z�7�xp�40��Na�t��Y�R�[L��`��P9" ׶�Yh�O�U��\,|��ey��*t��U�����tP��Dcj��x@�*�1�*\H`˾��~2�� �r��2?f�WJ=�P��]9�HR���|h��NU��ѭ��gw"�{K��)���p;;�d��Ul�ʽV�����xÃ�_�Z��R���F=��ɠ�E��L]˦���/_���n���Ҧp��uL�5l)�C���e���X8�V�⢬V��V�pe�pi���rm�{k�x�]C�qA�^T�b����к�k�������,2��2n�j��+J��h�>A��`���oE)T.���j�5؞�hL጖L�\FV�tyP����ãq����e��M��G��B3������7k��Q5��8ӡ��Åˮ���/{����2�s���5�T�OP����EL���y��v
�	'����!\C��u<v���_*��� � ,hѠT��Z�o;3x��T����9t�t��P(��� o�r`����id���S�ƸS��g��p���Z�oƵ`��;��@VP��5�x����種
��xV"�f<ĖG�j�v����LT&��Zͭ�hX�[�>$K��T�X4//ik�7b)�]q�Z[re(Y��Κ�J�Ԇk��O��2��p���f\l�\����]� #	��0>81ہ�����V�>S{c��*��'{݋���A�J:�ƀB
��=i
���dC�v�H��
�����
�
 wpF*]0���.m,�L*h�`k,Yzy�}��jz��*��f�|`i�N���g�  �;u��)�=�Q������(�u)��ښR�C�d(خ���G�s�5�QxF����: #1�:������0��t_�2Ԭ�+����YV��MOb�H�B��\U�H@lTN�V�%ITdm�po��j�D@q�����U9��pg)�D�^%�ɣ�i�̌^^��x{Ǉ����MXa���xo�ҋ%<]��ͻ���5��sq'�7�`�x{MujU�Ʉ�B�����A��v �(�*u�\;�s2MA��2[i���t	
LK�+�J�pŽ
��ISؑ��&���v�zުl��\fjz�m/1lK[�:��zU{�(Cd�p=�eh���1N�4�+lR9�����}�ν�
<%%}1r2n�8�z~����ͷ�S&fGW�N�e�Ț4'��������2��N5��b��Y�_zt�!{��P��B�n��4ϓ��R�/E����`��j]��	Y=az�hc����D}�L�J�*zK�}B�·�=�&�J������qsh,R������j`ϔ�sq�s�6�����R��KF�q���i��=�Z��]H�T�/$^��:�|B�~��i�f���Æ`J����*�U-�i=ܯz�ixا�W�v��d�Ҟ�^� ��Y���j:��-ǩ�ިp��j�;B"����)�ʂxݚ�AŠ�ƺ�w���s��!,V�(��H^0��'󮿔��>҇]5O��n�70s�zwu1\��Z6��p�t!l��+�ꉬ�z`O�zT��D�lS�O-���P]7�^x�=�{؍��r�VV͘uw:u�Zr���(��Z��X���=̲8�.���S��A�[�D�\��0^��'Y�"������2.��_}�V��k���P~jUvxa+�<:gG��S'ާp&��Mm!#��{���$���zo����EU�k����R�\�N�F�ɍ��6�7}Ҧ���V/���W��`��[1oEN�Ǧ�B�?$�s�ٝ!�[%��g�s}9銙U�b��S;���F�J�*̭w;Yxn��&��g�xב�5��ЩV�p���k^��K��*T��zx"��K5�B�^��j5J�"5�<<����iQ�\��2�6"��J�_V��L��Ԋ�ڑ
�"0h�P����Q��37�E֊�k�ָ�#�ʥ#�x G�ʚ[�&ffv��o�j)R�[;T��j�"��+�a�F�����h�*|v?�Ǥ������T��5?7��VhB�*�ѯ	@��9����j@�❍���\"�I��we��FT�9��~�q��*o�v 9�ä��\�w��Ҋ�!�cK8fq�J�:.�[�ɼQS���*f�����7��ޜ8_��Xр�hc7H��iW��d�����3�.�D�����nCf� �^T���Qji�5���r��.(��;�:�(\TT���q�WNh:��1j(@���V�eշ�ngd�g}[��,ղ�*�T�jq�K}�p\�U�5��n���I젩{�qX�`��xռ]��x���\�%3p��K,X��T�p5x��s��}^?¬�p0F��/��H[ˁ1pŕ��E�Cjv�a�"-4�@��oK<�#\(��� ��j���#0�7~��gJc�.�p��Τ
��X����R�p ��t�Ի�5��4������^�!ᘸV�N���JLʥ,F\bv����x�+Z@��p��9�o����4�ʩ�+��,�5P0hU�;�;cɚ~z�����|z���a-��{�T��)?s����x�\j=�p֩����qK�4�9��z�dud�T�N�Q��]3���j�d�D�TAa[�g��If�g��z"-	�_N}�^E�)�����Ypft�86��ǘ/+J�чމ�R@@�4pu�h�>`q�6.���)�뮭��ɄО��3¸��詚�J�����uJpS�ߴM)�N\ր�]9����9�<��k
B����n�4�Vx̪0�Q5�+(���xr�GP8�`�`�5lQ��C"�Ոy�d����
�9���x��ʼG��h�z��*+�ŷ�Zeg��}���[�ˈ����hG�K �����j�͗$�.��������YA�ǯ�Z
�¼��h�����r�b�>�ꌃ�Rk�)���C-�:�ʘU��-�ȩS�Ð��N7�:��Q��rڐl
��ũ��R"c],���ۜ�}�|+7���Au�=�,TT	˳[y>0N��w�_�1z�֪�L	�x�f�r[ksg,qC`鍴,����#��+���.���u��a/��z=�l�������W�C;���B�LޖI��sb���e�lXD�SY�.+٥Vy�y��}w����=�h��Q0q��E����#��<=�v6�c���>�ܩD��8M��W;���ROo�� ��j��� {Uh�vNCcc&��|�LħYtvMjh�ā�Q;����Hhk�G��S�R�r��~ � �x����pKW=���
��4���G��t{j�xU�0Op�.��SD�Mʒk��y�URT�I��M����1�}[��#�oy����&z��J���Y�� �y�Nw�%ӽ��h�K\/sc�x]���h�:�ex��#�w��w�>h��J*è��Ǭ��+S�v粣�^\٫�׏uA*U�LѺ�|���K[7�<��)N�}�ZmQ9ޫ��C�~u�w�K��*���%S;]�RT�)� a�t��U�'-���gU�VU�]%��d�f�WL�j�S�5�
�%*�~�z=�7��lf�T|������<>��ϑ}k����:҃O�^]'ow@'���:�h�](�:�˦�R�j�p��1�d�a��[��wwJh�=^@Q��H=�n�⿉������`#��/lS�{��Q�Z+��Q�	��E����s�f5�I�M�V��<ҴݚP�R�;Q�9*���	U��B�b������5X
%�h�z����4}ʍ-\:�hs��edy����V�s�Z�,n��ӧ/��q�F�>/ThL3P�����sq����qH�	F�����D�[�o�*q �����F��x1�w�ǎ�b�R��K��w�p�8`�Lp�	%P���ݙ칻�z�H	�����m\<�[�8r઩4�����n���;��3�$��>��տ
�ϔY{`շ}��2��8SMVt�H�����b��R�m�|bK�=uq|x���]9T��J�ZN�uұ�B ��ڃ���5�G��X��V_W�TU��Ns����M�g�0Z`_|B�v���{��{���^�U·֥X�t����R9ǂ:��z��B/�s%l��gzU���V<O�3@z|֌pxZ5j�r����wFa(���=�,$L�CYs0Ъ�*�����hB�*�ѯ�(�w��V֫��{�Ա=Qp֣��
���/�w��ׂ�r�8~7����U������+� �hmyR:�M#Z�j8��p*���QG����2{z3ga�'>�~pPoZ�!��(hL�_y�Քsٙ��鶪Bѫ+��J�˿^@��Z�b�g��3ۈ/%���&G�E�+�0p�X�yS��t'o�Ϊ.Ҝ��`D�sJᝳu���e[�2���^��B�֊ߣ��ù��]�9׺�Ȼ���)�}�9�Һ:z��1n��Iuw���)zW�XH��4����$7E|�JXeG�[ӹ�%����,H��-.�����
���#I#��F���Z�r�o+�c���B����V&b�C�����&�e3�q��l�hD6�Vh']�9�ì|�+<�+�k�k�����>W�f��䝂��&h�{JH�m<���R�S]�C �=���0(o5��Z3D2#�@���Cc*㧆u�|��yI[��8��Hp_[t"��ε�Qko
d}����f�LגXVc��Cjr��s�eG�{^7X�9R�1S7��ݣ�Z�î����h-�+r����zX�nw�չjQ7f��e�����L^��v�M������zmrJ����%����V�<U�	!Oyu)L���moB)ڈ��R�N|AuûV�q��z�zzR}{��)Z�(9hX��	���`��M��˗��X+��mu��*��;s�E�h�{���9��J�a��v^�>�s"�P��v����f��#������T�Дo�t9��4��nbLκϝ��B�����+72VQ�ɍv��u�Jb.��(u>�*CK�����%���N⺑*�7#-B�R�ƀ�HVs�֔iQ�+��p�J�P��N�A��8ёsV���P�/^��`�J�)�Q�e��[�wWi7�\:��;C�8��d�̝e���K�'Qׂ�v���UY�$��,rݬ��=����Y��s��r������uՕ�ze���.��	W���i�3u��|��æ���v��(2�;^�0�/q�	�iΛѧ$=�S2+����G�M���T�9u���I��:�e���o�Q�MM
����2��_a�ڲ�.~�k$b7L��pRmLY#���םi�Ò��cZ��TV!�[�30U��M�H5�yf�_p:�k2����h��E8�s���I�d��H8�]�I��wŶmϝ�m/A���kV���ki5��0�
+*M�E���X��32�0�ɳ$��	
hhJJB�:�Z�"�&�����iʆ��Y��CFH�d�!J�A����ęN@d�ӑZ-��FYkX�*ֱk#RĚ�ZZ��QHm	�RD	�V���"�\���(rV��L�L��5+NђPU
f`��u&A�ـ�X4ف������P�(;H��Je��A����������DR��|n�w����ɣ�{��r�E[�[�;�JS��F	�r����;�˰c����>�O"�3?G�l�s�3�+/��A�Jyp���%V��cbD,)�ܥ"xTd�bܝ�.���M�	���R�p����{Ro�A�9Ԩ\t�1IT�]{9ؘ'�	 �!���_l��4���=�)���B��lHw��t��yʩ_*�]��d��Y�k�����Yc��ć��u�c�ʦ��S�`��V9�œ�7���d`�X�8�h�k�<���Z�ޯm��)��� 4̧�P	�*�L8h׳�^'���<~�Ǥ����$�����I��c�؜���]#�Sn���5�O�����&ﺊ��q�����f��J:�"AW=FC˹����w'	�%��5F�9���{Ʒ���>U��#��Ds�P��r-���{��<�Z��y+�&>�2kv�db�u�!��w���]i�U�n��	���G����Qt�V�G��d!O�n$��W^]1�IjSe$	��{;�`;��s>���};ނ��	5_�n�L�'�"d�+2���*o�X�	dX���ȁ_;�U�im�Y��TO
��SFk�;���zKK(K�\�3OeuU���ÆP�����i���=ᾫ�#(O�76�gn�%NJh#�Ѣ����K�������YWBד�t�q�s����4�0+�Rھ� M�N�@v@�
���.t���p��|����7��<��C��<>z��� bj�����M`�x�OczpVˌ�d�SF:��a��c�����r�Q*��!o��+���t�,{�(*>Z%�Z�� U��Fђ����F��Y
Ծ�V	O�e=,`��;���F��F���q��W/���&��I�xת萾gľc�@�B�N��Vyy�yh��=p�3�u<�č�mˎ�bճe�'�}�Y��b��ӭy��ŵ��Ӭܣ�XЫ/�SiL�9%�R��x����R��c&�w��6� ��G�8fl�,�_E���ޟr��)Е�~�ky�H�Z$tiW�ЪKA�ݷ}�y�Z|O��xV��+N�.��<�K�)���y.��� �|L���g�b�Y�F��r��G�ګ�mw�>h�}��S�/<{�t��hlR'����f�#�Ä�*_i�,:n�v��S! gn[�U$eS�.�L ���W��|�**�p��V:��{�M����L���v�j�;U.q���vk�S�zX=
$SK���V�Gi�F耣.:A�m�t��������SˁH��\�m�=�Ň��O��[��.,:[$t�����W2����`I�r�fFut��m���%V4a88s8����
��Q6����\��Lz�\�Eb�<txX��
�K��1��}v��c+��h��]\���^u>���n�5��L�4�������n��T��/WGxFHTn;�[�He�����'H��d����.��9$��BٔOI;�@yc�
��l�h]r���>��EmĽք>/AL�ۘ3���慃����p��p�`�W�h�a��+�ߜ�^�^r� �z�b<)P�\�*�K.���4%O����Y���ԉz�ʘ�B!+���Hkr�n�֝�W�G2��xU���?C+�����g��Q��bDf�?т$��SQ9=.*(Ls�=m��κ�=�⧕Q�sm�>�"xs�`���:D�V� /�G?���h�kC��.��e?��mΨ�Y���ux+ռ��Yഖ���|81B̾U�UP縝}�@�2�e5]0bT�e嬄9 k(;$l>����Z�r��F��Ϟ��z��}Yz) ]G�V7ƈ���Z�h�����^%�=���|.M�%���9y,@�Sǀ��x���Q帴�"14Px�U��t�^�+�`Kǐ��������[n]��d�3M��������lhgW�o%Ų��G�U��5�L�W|��Db�NH`b��@��zT�˞�齳�a�CK<��豚vlR�U��~/�'�S;m��s��K���{�)q*�><���*��Ae���wW��Ą.�O;[��p����pKw��p�S�����86� ��$+M{�rT��{m��>��@�fn/�Z+hL��R�Vl�!���Q�T��s��Fw�X~��q��=���>��V�W��qy�ln��L̸��" ��t�s��~���V�N�P���JL�^��g��XL£8�.R3]0��m�Wymk�&K�Gd�v%�wv��i���.hȜ�P���N]��j�ۊc{i`�*0��_s�3��\��^W�" �8 ��4tG�(:υ08��xJ�#�slY~��R�����y6e�C�}zѝ)�ߛچ�$�k6���'^�5�h�]�iu�2΢^�s�/���j�(4�]�g]t�Ө����U}��j.��r_
y���r3�Â�j�(�Q ��Æ�l����x|'���>��z�	�R�	3jw�NVE�R�!W��t�O��i�V�9�u�\��,�ꜾX`�uA(���b�.e����2^�#q����lF�8y��!⩚>�Q.�x���^��kDp�Bf[�{ޞ��u *
�a�,
���i�Iچ���Px@��S,�����w�����fB�_;�\���Z�l�׋AX�Vd�y�Mz�n��}=��pӔo����T*с�Y(�6w_s���.eF@��.eF�����Vޗ]|���k<�_
M.�{��=t�z$g(��7\��u^�^�*�����X%���zn�����|?M*e�]O.��3j^�s�Ãzt���.ǸNL^f*M�V��4*v��]<VՇ��H�N��S��8�jm6���`�=���=�,'TQ���K�a�k�O�R��ZQܬ�z6Dݨ^�)�(� ��/1��m&�^������郵���)��J�Ô��4Z(���@K�Z=5Z����b	�vC�<.a�M�9�N!�;6�NU �ZIb�����i��p[�'C���³�������|L
�*4;Q�J��)��B�,�T%:�Z>S5�|=�e��F�#�J1p�c~����@7U"=�Tʜ��-5�V�f[T��o>�gӑ �o�܊~���u(*�����Y�+��x�j*�j\Ծ7	�E����
��9��1��Ȍqp�OƢ,�28���� T�rV���N�=^�u���4�(�'����V<>���A_j��0yq�B��R'dD�p�e��#����t�,���S|)3P/��������{;Cy6���Cw�GF��P���ڏ�_dD:��c��z��� 5	ݦ��:��gh�N��ǈ���}X^�J]ٖ̂��b\f��@�r�nnIPPGƽQ� ��K����q]�����9C�{���Zр����8Q؀Q�;N&Z#��#�bx{�)2��^iݭ�׶�T�SuF%i��e�6�|0^X�%��Q�]
 O{)�P�lmQ�q���h�u�����[���OZo�I����t*� �f*��xS��&r6�ųp\#a���XNM����~!澿�а|1V�\+@=<%���6�k�<�4��,�j߃��HAK��gB�>�\5%X~��}�\�&�zxa"Q�8�^�J�xF���j�ܩwf�Y�yiB��GIsҥ�PB�ƇU ЄCץd����>Y��d�;H��.=����#�,@(`��U���@V\Q9T�s�e3u�t�j*{�����Y(��i̧���	���kF��6�֑ʐ�yK���6s��E�s�|��ڌE��[Z]���z0��-��:������>f&��.e�2wH����� ||$K��vU���f�C�3�I�2��w��5TzeL�ձ?j�����s��E9߷�V���lS܌� U��務��Z�$Gğ?v��C�ϽPR�!�82M���ٮ���u�s@��ݳ���jMA�T.l쇳U�3�$����y������;J��:FJ]Sn�#�t/o�o����c��c|���I��m;�&v4vX�i�%��k���� ����2�oM]��{�6��<���"�U8!�n����!=�ι1MU�W�<K�nV; �-lm�b�{��9	`��^2�ܦm^�Υ'sZ��1��oo->��h=�B41���ڒ���O�MiQT��N��o���T���mE��v��yZ�N5y���G���m-�Z��e�䠀�U��U�ȫ$�F�����Ҧ�zD�Զ�2.� Q\�tu:bCgsI�}a��3�)=�,	O7L��e��]h�_L�B☸h��5�r�4�G�p�ZWm�3|�n$TLs`�yr�e�y��x�-�\V5�{v]@3^��2*[�y�xS"t�([Q\5���`V�WÀșB���.���o!� �
���g8���V���sx�vu�
���q-�K-���/F{ad&�I�QMR����X�_���������Ǯ�۳3�'	�b�[=7is%�N[98D�g�z-iS|�������G}q%7\��=�T�����`SB���؃B�Z���A�����c�nw`[Oz��ÿ���Dm�]C��V2ƅ1@zd\�6�C��Źs��(��9��h�j/,-�א�Y����5b<{�m۴���@o4.��rJݿ�a�D��6�E9�Wu`}Ångw*��C�	B��`k��x7M��~.?���.>r�CsԲ�]���R��xJt����v��Ь�����:3�x���D�F�]����Vk��*̗���ՐΥy}L@�ڛ,P�:�]O�O���)����7���/!�ղ%���[�و����(�#��"�{a�l�έ�J�XV�!θ�L.��ըbͮ���܃qĹN����aUpU�Y(�S$�qջ������:�;�j��Jo�	�5%��8M���=n&�9��d����9�g&[� ���+�n��z!.�#���3E�r�#6BDC��_7ۇ��[9Is�0�2���<)l�6P(9����T{��kKW;�]d�8����v�|)�WJ1�R���뺷���o��������5']8�����_�I���c�.gc����w��,s�<{����u���w�v�����G�����.k���cd���iK'��Wu�;���rK1�+2�̈f�[��J�uNq��y��E��͵q�*t����.o)���P�+��������q��<Ƶv��I�/2�<��'���M��ܫn�)�l�B#��m��0P��s)� R����V-}�)r�c�|.B�T)Ԝ��{d���s�v���&�@��,�&>����\��V3�2�ǚ�B��}� ���9�EՎ�K��z�=2�-MI$*�u�T�akө���mq���Vfm>�	�����]���ӕ��Q��sg�nM�]h��_S(IJ�S�����X������_,�R[5�'q�#�Ihˈ��q��)'\�٭�b���wk�;8�~�P��ݶ�!�eH�Y���T�!B�T��ǸsX	�jZ�ʵ��E�֌�,&�Y����N�`eT�Pe���r�3X;�V�fHR9dJe�Hd��ԙ�!�C�Pjw�#R�	�aj֍Z�E&��-E���-e4�.M jL!6��K�D�8N�151&A��f`֤�V�P�PkkQ����&�RQ�M��j�� �C��()��3|M�Xd���XXe�V�R�F�$)*�Uf�5kQ�M5m���i�bѰ��T³��L��F� �ΐ"lN���i۬���Ƿ����c��7A
Jc7W�j�s�t��(��o��Pm/���7^|�����r]�U��9B�&�O-�]J}���N˶��:c^�N�n ��m��p��� %�r��dwM^v�R�F��[{��q%��<+���x��8;ee��8.��u�����L�cB�{�������JÈ5��gza�"��c�-��[q�ě�!�R ~+Gq(���]���J杓R��(4�.���y)��2v�#J�q&4c{ؠ����yTIG#�@�;�B9�v��y�V�wIEO/�b�k�(7'���>���m�P\oR�(�ى}����Ѯ�u3�����&��cub�d��%
��w>�a���Y�J�+w'�,�	1��͵{2=/QN��5�MBq�u%��]��y�����9�U\6�gv{� p׫0b����~�՗ŭ�MN�f�7N�A��F��Q���ܺ���Û�F��1�4�@q����xl[��}��sXmt�B9Τ`�57�����qn)�|0�7GN��kc�S�J�<����QUج��%���z�)�[�"BXpMr��*ŉ��Muu-��c��W#�bf�W[ٌ6�����W�&��x"��ݱT�:�wXL�=��~��傞�:''�[f9_ȝ��(pu.�/4��&-�}�l NǟjHH�6��#L�q�t�S�9B�[�[��5�m~��ђ�`�՞� U���l	 ���ؠy(��:2���&ⱄod���rM1�9�~�Զ�|Z� ^#s��[�{�{��q�����F0��ī�֖�9��S��<��SQiĝ�	P�U{����9���U[�<f��=��6Yɭ�r�@�7�;����DPJ���C�AS}P����bܜ���;=F')F��p(���ے���u'�⋫���-΋�vv�7o��⬎�i��R�"�� �eY����X|nN�&M�Q�~'!�uD�����$؁����f��h��+�o���@��m��W�@]��.�	�&���������#�쳨��2�r�t��H�3�p��Њf�.��~�E|�0mۄSX���I�����=��MK��2,�E6�n�X�ʬ���D�ӗ�j�L�fvt�Hb����ŵ.�5vN�䖼�LѲ"�%��5��tf'lL�Z��m�#:4�p��Υ��<�WB޾}7 ۥ,� ���]����Rl殚��{m;��$��қݬaEg.�d>/��/��UE1}��!���v�s#]7� ~ם�B�"�+FA�5(>A����_��
m����>U\�I��#�0*Oy�^�}tEZ9h0pC�s����kX���o�=�#�d�0I����=�I�}T��'c��OSE��� v�#	�U|R�}����f�y7����D2rY����lED��R����U�w��)�+)A�U��mm����vLI�����{��1T���IP���(�&�U�,���d�X�\�U�#��y߯-q1ֶ35�h$j������c�����4xUǟxL�U�>��A+�j�>����V�3NC܆�FЂA�s�L�nX����=F���3�#X�$��P��A>�pc;���`@��y�j-��˿b�:�sh��\��3�.�*77����dGnt	�H_M�Nf$[���(Y4�u�7�u������s�qV�?����Έ�5�>�;D�[��O�D�\Q����7�w��%����)�V����v�ߪU�j_CK<���w��./Gm�9�L�Z=�Ѩ4�Nlu@p*ʆ-�5Β������|�u�Ҏ�ofg��T,%W@�f#puֱSnV�m�9�m�N��Z3�����7��/��vۮ��Y'U_vPњSp�a�6��)���3�̭[�7&�j3�9�i��b�r�1�ܸq���fю�sӣ}���9��Լ���U�n�sh�Ŝ�!�]�|�w�_9�J��
���3���cXI�n���U�Pڡ����z�Ȥ��vtiǕ���c^e�y��Se|���Vxe��)��:���u�F���x���{~�7�z6�s�n�뭺���Q�ye��.P���$@�����w���ң^rǖ,���t�����F��`�=���M�3��&� ���>�q�sg	�6�{{Z���&�::�5��� ��pO���^�ש�N�{<�Ǩ<��:Q%��4�rD悹�.Q��|ㅇJ�f��uX��h,<�-� Ŧŭ)1R�΃�*��j���i�shL>��a�3x஽�����B����6^��}̰�Y(n�{m�Q��ۉ0�E����,�9Z!�G'��^�<"$��e�Ha�ݻ��jMeGk/H-j�ZJ9��(�}��>a�[�:�BBy�M�{	W��ͣ�7�ޔ��x�wlaw�^�:�e��䞒�"Z��sZ�&8Z��q��Sun�-��}�M�R&�8��>T�����]�)�'�¼�s�Rg��dZ'dz������C�B�my�P�|��hx��޽�2�цVE,���):����F�x,�ZOR������.�&�2�V��΍����9SUڼ��L\ �Ɂ����'c���rh���Ŝ���$�����7dg@����K�x7�+j	px�
Ly��[mi��$ާ�&ׯ�2uݕop���p�4���FU��y��闑Q?Z�ݗC����6�rǃ]�n��j�_t�=G������["����9�e�}a>)E��J�����D�zjB�G9w�q-"�P��]h%���.�΁{"UԱvƐ�FN9�g�Q�c��Os���)'���l-i��n��m_8�C|pq�;<�}�������[k�pB��]A��f��߃�������Zb���ž��u80(���b}O0��Y��Iv���n�)��6su/"1VGn�-��B��'M�iR��Ԫ��͋�}�i��1�*	�O!�B��c� cmI�<\{WF��B�K�O�?*�x�}�7�~GO&yޚ\g`dƖ6�ȩ��j����.����ϳN�w��-�OJ-�S�դ�Iz'�_�|�u�,%��"�\0���nfW�4�-���5nw[��\��T�� �9ukK,�C�'�'������Y��L�imզ�M������bT{9����Ҁ������_�hs
�C�^g�N*U�E��-嘅+2#]#�{��S�j������]�!_�u��r�yc�Ѝ���\kj�<�-;s�CwuN��]�*ݽ�j�>Һ�eYK{u��n?�X�E�r�yCu�J�>x_��NN��C��G�]����(Jl@
�E>����������{����sY���:�5U���:��B��:Z{Y/^����mTWS�r\�ޅ/����	t�ñX8%ɣ4���ʺri��w���d�G3�/�'%~+FSa	�3|n��/����-���t��'�R�G^ͅ�]w� :q
��eS�]��%e�O�m���3�(�[ǧ���� P-�ۀ�g��oK����y	��]v�M���{{�*SO�ߴ���1�`/va� �&p8X=|��*�1�E��i�;��Ya���k ��|6yl��=r]Q�f����}C���D��' 	Fn�����p��K��B�
�2�|0b�.�ݩ'+�\�*�#j�S�+N<�"�Pn�Dh�Í����[A*����J`�ڷ��%x�J��&�|mNAnҙݝ��2�,�m��`��5q�]��]�Ţs�4��ը���;{�R�Y4R6�����)�Z����w)����Y����u�]����(��|6�K>!�R��82�c�"��2�*	��XX�Wu�wZ�*�賘�Ŋ�C''����p�˴o�����M`tp��Sw�o.��'+��:+��]g�\<���5�OE[#�+y���9]��e=H���l
[��z��i�ƭ�u��nBJ�}��AQԶ�vB����0[����-
݌��':Y�;LN�5�����y���,vVn�n��Pdt���z`�D���w���?Ih*X��u�풻���z�+����Q�N,�,1g*��24��S���~�K��c��U�y��׆��1��i��hT�v�cZ:�%{W֪n,�n݀���Qؕp�UŴ$gl�� '	��k����[;����[A�X�kѢ��r�]Yn�S���e,�/
l�Fn�S�[sz�V7��������J^�s�Fc�VeM6c�sKF�b�̺�z���	E��u�}:�����J�x��, $㵴�X���Q��z�6g��-^K楌4��|�<b��Ck��8\Hi5%�p�O�#O]lɀ��H�9�t�ZMZ����㙚��ivcuXbkS���s�|fqH���i����	�� 7>5�Kw�i��5k-+a$��J�K5���!S���a�o	ρp�Z������O*H�z6�LݻpbK�G���W�8O�1�;��xe$�oDQ�9N���j��;��U��9��D����	�s�ӗ7�R��6�3O=c�|��+�-j�� M��ۑ� �oW����9�/�hC6�_$o��#f�4��)�p�ҍ)U�.�b��=�NoWG7��z��0|.�
 V�VY&�f�5����Z��o0�h"�U���a�k�h�G��E6m�)�R�*̵�f4��ؙk6�kX�Z��h��Z��Z�2���M������9;M���56�NٛHV񒚂�mf�hJ

��0�(ԘTj2MfPh�Ժ�9���UB[cXM#Pj���35�,����]dkVj�SZ��j�YZ�ֱ�05�
�u;�m���� ���X�d�d��:*��&"[Y�fXeE�fdNf��(��5�ִ�PD=gM�W�:2/hGGA�D-�"��U&cב� ���.win(�;�1�ܾ��_�`S��o]�5ہZ��k�	�E3�Ƚ�:f�p�p��V�#�U網C�"i_$RB{�3s�\�W��X����gw:cRel*�5�	؋����*�sQ�9��	4m��Vc6�]F��X�"��>�{���)%��[ް^��'R�߷��_N�0Ap��ow���d�����l�Π�P��g��Wf�>Oݵ��!7�
-v`9'�HThD�ȫ$����.�=��5/\]g
�h��j(��ۧV�m����:{ �z���ۑ�o2���|��ɭ̃[�E��9(�fAN��J�?M���A�	�����"����FR�1h�׳����o@0I,܊�/�g��� ��`�!I�ѹ7����~��:�+�b�{�^񤑃���'�Ȥ��T*j9N���l��$u�NK
���0Z%�5S�����mɾi��%�ӣ�`5�e���A�&f�����ɧ�-O̾�iy��ɪI_�$鹚�F��Ӳ0�[P�]e�>�6�=:޺��x�>dn��%)�W!�t�^Eٷ���(F�3�+�N����5�[pnl����w�Lu��Q;P�d���A=�����2z*̗l��jm6j6ⳳ�O%=ʈ͖�a}��xyԄ?*��yR�'s��Y�J���;&;���=W��+�Nc\�gb0�wO�7�i�|B4��AfS��h��r���95������iQ n�v*�yM7�VwR�D�#7��կ�@l����ȳ���*|jo�%�*l�B�Π�އQ�4����C�5���{R�������h�ڒ���~ƺㆷV��	ȍT�Xם��(���K�Y�&{�"PU��{�H}��K��uc��܁̱��%���=!WJ�e=�������-c���-G�D���6�N��UJV��@!�wxKZ��G�N��&��&/��v�Ym������s��<�"�	q���l2�+�$��c�}x��,��{��t�U*�+��)�>�4j�Z�&�ӽ_:��W���{��~�w�٦p��):��(�MԿ�<�\��R��O;�UjZ�}Vx��ub�����M:F�ĔI�/Nb�'l�J�-��F����sGB.�� �c�q�v֟.c׶���݌uft[x�;��1�ſ4�!W�Y�'*�����ۜ�Ft�s�QR
\���GFl�t������~v[0�7Fu}y����L0�vJ�Tu6�41{4ԫA�W�pK0�K�c���;M���0U�T����cy�x]�[�e�Y[�W]�D�v7�mz��%�7��)>��=��i�0ܐ�^�7�!�����T��.hy�PT�M�w[Y����t.0��ĥ�ˮ%����3�R|�U��q���y�c�S�휆�f��/o��}�|��Yˡ��$x.�^����F��ɳ"DT��=�-[�{XW����V��Hْ�w��z�sP��]�`�>ܦ���Q��t���0��<�yņ_srJ��[��*�ݶ�����]��g����Xn����Kc%��auC�X9�!ފ5�U܌�e�˗}����h�9C����.��nb�I��z�����t�\Tp���l�Ƴ�{w{{�:�Z�*4�sT��u�jg�/hs�������y���zɨ�2o�
�U��6 f�7���H�3�J��ߨ��ҍmCSaj0�K>�T�������Q���V�'n͵\"����r7Pw�S#�Jy���l����E�d=C#S���̽��50T�e�]�COki�vwiz�5-:�d�*��ޭ#�<K1���Q'����mH��I��{�_C2�
A�{�US=#]��Wҹv%�ɴ���b����yG�$wq�ӥ�����_-�I\�e�`�/aE^ܘ�rp֔tc6��㹥�\!��,5� �u ':U<�So�0��+1 ^�Y��Q^��25כӐ��>I�Օ�&.�2^D˂:��6�܍&���J�>H@��sn�f�dM2��uH��������Px!�F�s[�Cy8�n �S�tt��'�4\��69�<\���Q�`w������[6�]:��N?hs��4�ςxŃ�ݿTi#AR/�ߤ��3���Y�A{���53.č%s+�4׮:͸�Yzu�{�}����X6��\�|�4�U��u�����d~�s��&X
�yN	d�Os�>8����-2�}���4�.�W�+�j8��[���3�GB����Qv�dֲ]��]����d��+�ESՏh�$���������^��Vg-A{k*rfjƓq�2n]Zz�J5h�$'��;"+2Kgb��d#�J��(��\���М�m���1��԰��t�=Tc����ԁM��yN�]�髌=h%�	SgWI2�D�-��s�[5�c1^�wÒ����y'`Y7��-�0}S��WeƝF��=��〾�����#ݍ4�OMGt ���9����uZث  �X��z����M���g-
�{q�]\�� ����cy^��\gn${J��s޽,<Πn��m��I�,!ґ]�Y�F��������@�FY���	��r�4r�_{�ۗ���4�Qȧ,�n��^<�{*ܸK;9����;�K5� �}�F��x�m'���~�ALRv)||߻*M�'��SQ���nE��{ ����C	d��=��	>I�`�車]�v"���g�5�'_
�]L��ru�u����5��u���N]��i%�rh�7=]9�Wyl!�);� �	��ݫ��ޜ�k?����ږ��
�^��N
�Z�~9��89ݜn0�S�z%�b�����X�K��o�\#�a���PX��z�jb�+�:xT�,G#@�芓Cc�d�z$��S�� �,.�{���>Y�nYz�Q��xԽ�o�4썴�.�v�$gfo5*�kdM2G���^�{-?�V~�oN�3����'J��[W͎92�����W:nd����f�%mY�M��P)sR8%�1�2��S9��8)pŊ�Zp�a��7���� �)���dE�[Rl���^T>(�iv�:0��\J]1˧�Ҥ�z3M�
�S� }�&�/�y:�-�t\ų3�ӲXE7=W�_�6��m{h�./rHC}��˸�W��ㅔ�5:��o=P���{��׹9� -\�[{��7�({��+��ޜkF��ME���h9�Ӂ�E�G	��n�N��N/+�Ox����	��H�zH@�k焙�>Y�����vk�2�aW�efF�2���!�]��͚�we���QI�boK��c��P�u�=�1�� 9�q�����nY���^�C��ж�U�<�ң��\��o0e���a�(9�������>��EYt�W���$C��ߔ�Cr��ũL����c��V��W�a:L�B0�ێ�U�r����-�g�*��i�	ERIƴ���{L98)�]nD�����Dnk�`�/[;Тj��Lw�bؔ��Y���(��P�_��ƅ�9~�V�۷0Kv��RQ�F_��Z��C_D7�w�OC�����Ko�pB����+�,t��	1�=�J�LB�|p �3M�鎨���НC0���#�'W�[�� j�� ����doλ�u����ϰ��?��T}xe�U�,UA5a��%PT��b`�*
�zbVH��L6�q��9�6Ck��a�6?�ÿ���$(��*(�(���*(",����;k~M;���LK���&|0N��`|ۇ/�(n�.{����kAPŎ�70=�/�N��q�h���!�v��#G��}{i���[	����8`s�iצ�����y��h�{�n�˰s�*	���~���5����?���A�P��TT��}t	I���O���c��`}a��?��?�O빇��4�4�i�w�w�>!���}߽T�?���?�����"���rĔЩ���6!9t�����v'�0��)���d��p��_C���Y�����A����E����sAPH��nc���ͳc���6��T�?u�үamT!�㎌��a�h4�G��a>g |}���*�����\>������6��?q����j&���c�|����~*o��O�n�����A�܁����j�������T�q`��@���x��'��!���86?� �熇�1LA?��g��#���~������.���|��?0����Ó�?PT��K���?P���|7��p�4Dp��>ބ�s�� ��A֪
��`�p$v��@�65�}�g�����tn�
|M�?A8>:EA8 ��RA�i�}X,�t?�UA1%���y�Xp������׀IƲ�p�.D|�M+�?�tC�'o o��Ӡ������ �'����a����S�S�A-���_�+��~@�����������	�C�D��>C�@�����l���h�g���>���O��G_�}Jm�_O�t��*
�}�������� k���`�������_�T��&���N���������'��>�O�������|� 胐	�G���ؘ�@���?�@o�����v| �9?%< ����+���i֓���>f�����*	�������N~��-�>�7$���a �>?0~^�}�a�ß���tn&��w�=�PEA?����� ���N�S�G�~�����A���?��<�����x�n�ߝ~�!�5����1	��������Gߛ�����)����