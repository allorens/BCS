BZh91AY&SY a�N׆_�`qg���c� ����bDw�  �u�[a���B�PZԛa*�*!*EZY6U$�mcU�٦ږڔ�U*��R��"��Z�Z��mX�f�D�2̑@�b���#l&��#F���֫a��Ԇ�&A���T4�2M��I��*Ŭ��D-��Z+32�l�c#M��h��ٓl�����'����V���t�[m�ءsn�V�5�l�m��Dڠ�j�kVͦ���m-�l���f3i��kDeE�ڙC6��3�ڶM�b[Y�Mke]���Vڭ�M�\=B(9��k*UY>Eثl��hth4��5���wb�g�l�C�]��7Z���� ]����:��Un�WR�-ݬ�l�-E*l���F���) �
�>�}ttw)�ڀti& ��� ��c�4P�ج��\� ��־�i�G��{�� ���� (�uRkYV���4L����L��@ ��|��z�p B�X�݀ w:{�:� 3{^�A@;���WAя^�֝��{�v 7���=��x ��/m��Yf�)�!�$�>�  >�P �y�xiA�hyӽ���4���B�睯x�҃t��J�7�@��^�ק��Խ� =� @�� ��t�J�tL���6�U��l֏��  ���  ��à :��4P�Ǽ�$���zh g�� ���t�]Խ�  <�Ǽ  ��q\{4=ޅ��e[V�����c5���� z�@�����@���@^�L;�@g�t@l��콕�fV  ��׼ n�
y�n�:3q� X�;+al5��!��ml��=�(  ��� � N�n�p 
�v�Ҁ m :� E�˝S������]�m� �7  :��0�2�[VV+fյ�}(  ���q� ��՜4 9�\P
�m� nN ["�@j��w]�

rs�v ;���E�mj��m���I�� ����T]�\ ��qE 8θ ��  ;�� 4�` �b�[��� n8�h�]4���mP�cj+Jj��@��+�� �}�@�ͷ��e� � (7t� 43�n�Puˊ e�� v�sF�  %�TS��JUC	�L&	��L�&S�R���m�44 h �JU( @    �JUS� �     ��R�"M�S�<H�4 =C@i�@�$MI&A���2bz��z���3Q���S�_�������]�����u��p�"��1�Mw'�}\��tvo�y�{�*
����UQ\DQAS�QUE~��E��G��y�?�?�~�������>ʟH���ݕUo�

�������%O�"
"���������"c �2	�
c*�2�0�2��c�0�0� �2!�cȆ0���c �2�0 �0����c �0�0!��c
�ʆ2��(c
ʆ2��c
� ȳ0�0��c ��2�� c ��0���0� �0!�"c*�&2!0��&2���"��&2��
̨����(#� #��)���()���c �"	�!��	�����	����	� )������� �¨̪���������������������2�
	��������)�(��(c��0���L�c*�
���2�(c�2	�)��0	�"c ��&2��!?��S'�o�� ���J?Ŵ�(?�ҿ���ZX��!N�R���PX��� ��%���@�xέ��M`�M�tݷYPh�D��K)VS��ނ�B�me�<��X�0�Tp\���uX���J�-j��-�QI��~	:f��X/`�n6pʟd3N@.j�o	QZ�RE��1�s�f<£���O��m-/,�ze՜0k���d��Vջ�IiV�3r,e�W65
� ���.�빠d4	�j�*��m�4,M��*݅��hcI �E�	��.g���d��u� �)��˳�����W|q��~ǥ't꺇�3&։�%X{JЈ-���Y*=[4q�eަ�nY"�L�7�rՑ3#�%���sփ�t	)�22��gA�6�5/$�pJ�)��^l�Ƿ�r91��*�:Gs1L:U��r�������W�.�Y�r`��Fò��f��*��n��ө��U/0�F�j!��[��(���P �n˰�ta��f޻#���0]��x���T1ɿ3�[�b{�`�^�N<;u������
[+E̚d90�,m�4�I�%�@Qkn­{6����@���� 46J��ذ�[!�b��"�rhf�m�i��32eX��-�ZpU�ᩄ5���R�Q����`ZP�S�+�eޚ�0��s�q�"��e}����YMT��c�(4;En��q�Kt�T^�K���"r��I������Ƅs1d�D؆g�L`�$�d���)�b�]��e�(eh���]L���4dmX�G^]� V�զi	�b�X+&8��򱜔qIB��	z��l�<���X݉n��ˠ�Q�n�]Cp(�
�Pm�.Z���	*��pl؅iQCm�l��B)�U����N�S�[>�]��R��ȃ��I�:�oM�4�d7�Ba���av%L�>z�����x�����SL*GC��Jb��j�'�:	�i�[є����דu��V�C ��`ɢ�^2���������%$�^�����6JYi��������n��Pڎ#6��Lh�&�X����ؖMs7� ��,��[nT:��3 �����=�2�AtV7�U^��,Q�H�3���-;1Y�#m6��]�p�7'�n�.A���G�|4U�w&	�b5�i%a�4��[��FE��73c
�v�%�A�T�X1fX�1�ӇO� ��C�:,s/��,��mqG��9�APlGL��F��.Asv:��[���򀭴������6���Q�4j|-��*���Uٵ� 8�3!��t��)6��`A4�F
ݤ���2h����Mjq2Qѕ�hn�ث�.@��V�mK��HԢ��hDʔ�ژ�0.�����kN�ސޕa4�][�t4*)�j���Q��C;M@�S|�*kkEe�"
�`��%`[5�6�M����1�Yz�*Qa��ᔱm01nn�4^�c��Xѩo*�i'sw4�ĝ]z��h@���ݸl��hą�@�� 	] ����]	;�b�;����pP�(���
u��D)L]�4�[W�Y�с�D�\F0J���xF��b�H��JYL��R��j����C1�WVؚ"�͝�i����L+�Z(%|3�P�zR���7J�*T��Q�R4���[�U�r�c+rC�ib;����MnC�y{4��T��	��HJ�e�t�N'��О�K�4��UbU໶�<��d"��ApZ}SEH� ZƯ2�d�g��D�ڎ%��Pfn-�ۦ�m;�K���{xR0���JK�2�|q�4�<��Bi���+�Q�E�wQ�*kf�a���lQ5�Eէ��*%n�)5�5݀�Mi��5���0�O2�^ fi��VY��k����@�L�Wy�P��{E�����xj`!�cH��(��L�������qì�]�r�KЩ����D�Ź��sm�˙K1)y6����Z[,�P�m3�����`iS٧�E���X"n���c��1ȶC�b`��۽�F�#tͅl�b�.��ŧn�`��q�I��/%/��L�@4��h�Vm#�儳E��-�i�&�;Z.�	\ ��Y�d	1T�rƘij�7e�.��������,�ot��5�ƛ��iR�G�QVeņ�B��	z���X(}�.��a�L(w&�[��Pxi��@^f�ڙJVϥ��ՙV��"�kw�̼�]	���7�oX�S)�E9���{�F4��u&��Q��Y&���A6�b6���و���ԁbYv�n�G`D$�<��2��ʍQ3E84i��JRP$@��y,ӕ��6�^��>���E%xh:+���\)���{�Glu[� p
Wr�~����:16�ts�E�	�X�x�0�V틲00o4�o:����b�F�7���6�z+Xm1����tՙ`�X��[�n�̀j�A&��W.���;��N��Rz���Q9Wm0K����|�����\4����c+��ol�)R��5��/��ab4�U�ɬ\�o��Ve���9[�I�{$�ln���V�8��l��"���;s��]�������fv "mkݘf�.
������7	Џ����OtH�a��sr�ڗ�J9����I�WWX&,F^�+s2�[��h�L��ֶ���WF���&�ב��ar�6	���_I��tn�TE�V.����R��dH��`ڑ��1�����3j���D78n��M�+\�	��J72��
�ݣ��[�^���̡ѩnM��L�t�)v7R�Ck���6a��õ��Oj�3�o"2;{-ly&S��:�N:��#���oVGub��CI�VP�!1c4!�v���Kn�(H���BEL���+N���GKn�=2-��"�ܑS�-��4���jĳ.X)�̈́E#0M�e��E��5��n�gF�I�m�2��	sj�yV4��1�š��[�pjy���CN�V�
�+(�Z�Gp&a��D�,���M)U���<uM����r��)�z%$MsuUwŒ�<H�k��A��)��ݰ�0f�x%N�ɕ5�%ں����Ϊ��[�����.��)��Ǳ���E��V<:(F#��42P�]�V��*1wA��5��i�f��J�2�*1oh}`=<�*Gg)OCVI6*U���Ǥ��%r���`�-�*e�(C.�+ʺHT�I�E�l��ڵ����f��x��V<Z�P1Y��b�4PL�R��V�	ΰl�
��h;�,K���}T3�;��v�d.-J3IB��� �`��Or��
�m�^r���`�ɠ+NQ��{�X�t�A&E�o�}�6����,Ň���].�ʌ���-�_cח(�f4��(� L��K^�u*i�ǫtn�l�%�ɩ� �cpm�t1�V��(�+%=x�7�����9@#yY��S�Nj��Ux7F[0�+q^+�"��6v��K+�����e1�P�κ�5C��a�w��Z��|n=�7*d�f�¦#�ZJ�0K�����@�$��Պ�Gj#���F������U��D�0]C���F���K�N�p]5bV"7�ٻɕ�����A�̆��,a���f�{.Й�_Po��KF`Z£��kW3[ٷA���5�C!}�[�)#�x�Ӫ=p�u"e�i�'� $���J���+��1�T.0�EQ;չY%iZ�`N��Jڗ*ن��NJב�A��
��=,����r�phӟ\cb�TSk0/���N�2�Ͱ@��n��P�J�k���<Zu�&#�I����3Cl�5f���z��{�ɩs2=^��f�4��hx^!t����/C��:@�Ҳ!%� �)�YC$�kUaڬ�e!�Xr�U֍�flnb�93+`y�J��8p������`ɹ���E�
���B�z�#z�K0Vmc��6*1��ˡ��RW6m�+*`��M���K��"6��H���k�[�)"�otfQ4��Ȫ܍���z��e�7seK�O�2�Ac �#�1̰��ef�Q[��t)`�E� Z�Kr�Gr��{Y����U�/��m��x2,mLQF�Rk~9���'mk�u�����l+ש|F�΅�c����0f��l��dK(V�wL���2d�*��hkq8���vs6�VH�^�/5���v1f$!Ʈ�1�����2PE���E�_, f��JëD-��Xn���gvm6��֪��A5�3�Y7�k�v�+ݳH���k�^�ӹ@ t+���7bx�bȒ�Օ %i���W4\y3죸�N���b���H��R�{sUu�K9qڈ�n2]^�[�bȑ^����)�����j�X�2�Xf,f����D���)����B���b�!a�,����5&Xӹ��y2Ơ*G������wM����젹q�k�x�Z�=�cJ��QL�KY�N���]BZ�+5��9���ѩ��i|)�C�N #��#j-V⫁YZ�Æ�+�)x7lY�Ac5ef�(�:[P,w��r�.������rЙ`��n���[x��3X[���0dlLK*���H���dH��k�ژ[���-���k%�_f7d���/��[thT;�u���nh������I.��#���ZrU�
0T,�x�ָ"K�ƶ[�oF�>���U�"��q���!�o@�/u)x)��%�a�r\w*-�8��Qܗ*�cF�+���¸�jo�_V���IZ�5����䌪r�E`}#�M�sQUʄF��������*1'�S�	^���fzҒѨr�l�����T�2
4�[v�0ҍ�!w��l��{��Cb��`T�o�@Ӄn����"n&�2M�V�LE yy����m�%J׬���/tڳ�Ξy�TK�4m��VE�V��y�F՘����ݵSq�q�����{Vov��C@�{C[�f�G���c�JQ��{���b7�ݜ+*�P�fS��s��d;�m^e�F�U�+*1b��2�����A�ĭ��/Z�Ư�j�em:"
y���� �'IX���IVF��ulI���)�F���Rڠt��h���c���`*Q��sV#����o-�m���!b-���/�p�[�}���I�Յ���idRj<�j�� �)�&�>�0���<�s�S�:�ic�"݅4R���:Cch`(�"2�C2�u+F��+q�v��̈���$Y��d�]e1w������n�D
M (h�F���J�Z]Y�r��� ҙ��
#��j8�����J����Zu��FR���]�^�٦׮��tZ�(ˢA�6��]7��jJOsQ�مH%A@� \���5�M�s^��i))�w*$����Q7B���f�M�ZT�@��Y���׬T�I�
�je�̹�bU'[ύޑx��tj|e�F��>�th���;[�(S8�h<�&��M3��r�Rz���f7��i��c�ŃwDʐl��{�Fћ1�wF�j�.X/YtM3��ЈWp]��klJj�
|��iw������WeB��P}h�Dl��Ĵiɵ@��:��e�=�6���:壝�����Թ,,�%��aY���d�MS&VbAZ��N���4�R+Y�^#�ͱ(�v.b���v���p	N�E`�H�2�J�`L���sLV0�he�ה�x��3nb���r����lX�ª�F�U&f5csU��Ɇf5�藡`$�k?d
��P�V6�+ZOre^B���5���"�� �k6�LJ�J���7q�05�i1[1�¨�ەyL�̣[Sʷh4��0�I��a�UL�ZW]:����]z��1v�͵���m�v]a�ݽ/lm��0K��ۊLC���a�-I�����s*S5{���U�qlǮd�����TJ���]�{h[1ȫ!T��1�[�JD������4Qx�=!V]��ɔ�\��$���15�K���^ie�y�E�z�tki�Ro[F|6�4ؑ��T�����{e�Y75�D��@J��G&DqD���8�����	�En�YX72�f'����B�i�e@f9��.9�wd`2-	X�YȳJ���h�:��u��&䣄h�rÉZ"m�LRM��T�}{�V�V:�������CR&�ep�MY��=�`[į�M����hǸ��b�F�YMV�Tu��`���lE�6�n0��I�}��W,�{��5�x7de����_PL�֮T)�ޮ�*�W��5kU�5�GXX����6�b�wf��N�Y[Ytw4��rm�æ;�N�	m�xw����;luc�	4U4�ٯ������-��N6u�j3I!�n̼�Su
�"`����4nMw�4-ї��-V������`5gd�������X�TN���3N���&�]�$ǓtEn|�;�S���.k4����^QT
7�e�OH�]�lp��91�;vt8�w�l`�0�e�*$mlǲ��+6L�x��V�KN:0�4�����ք���t��w�Y��Ցx���4b6�yk:���Fk��Z�0��f�Z9�h�1�d�0��9.����I��p�<ŅRhll�)�T2�%�l��q�Nښ�`c̥%6��Y�c�\�+ح��KZ9ӹf^ł��d�fX��NAu�-Pa�)R�����ol�.fLJ&��1�M���*����>cI݂��쐑� )�C�[��2hY��	�l�3������G����7ܸ�w�:AZua������R��(wU[]��=�n%iv�(-�a5�%"�CvG��[:cv�$�<�gOvv\����#�ƞ�,���%���ӱ��� N��JmZ���h��#zc.����B��9�6�a�Q|B^9���L_����U���?��������J��y������%�ɷ"ž��K0-m
��s;���D�Q�B��GH��9Z�(��ݐ�� �2���0C����L�vD�R����� �:�J:�ڏ{�i�~,�<r+�Tٮq�B^R	�ӑ].�F�œ�,�#��Ɵ6��a���X��U��P�@,T�,�xc�T8�,ȮE�t��NuEMk�
�.ara��6@��S��{PenAQP�t�*�^M����N٫5s4H!;�du�q�$�q	�c��^,�ޕ�N�o.�[ �(a� wW"&�%�)�jr���uV�=6�XgJ��ؑ�n��4m��o�4d�[�����l`FfN�`�{�ݞ��A�iHO]iE�O�%���X�E�ok�s�,e��m��¢�[`�牜DO��qF�s�",S�8��):Oi��x���X/�����5y\��-��c��*J̊`r[$�˳$�7kl.��:c]E��6.,ԃ��4`NCT�DZ�Vʜ�V�w&p�"J�(nk�����yfՊ�ٕ,0�;��i}�|�.X%�Ԧv��AslR���n��ۛ�	�����6�+E����.(��p�u�LT����p_<��8P�WBzu�q��a������˻ptӋx��� &˯����`L;�K�+��u�1+����K��m�q��b>��E	��tm���݌@꘨g^WN-G:���V3.Υca���Į�2�*,97Y7WN䄃P]Z[����C>��p��3L4a.�<n�#ʐ��e9�~&�횢��u��C2J7�x���Rb���r��%c�nT۠�B��js����pj6��Z���l��@L�'KT4�m4`����M�h2�s4"7�++�sꅝ�@�Ѕ�S��Kvwk�-������\�N�V���ܗ��Aٹ�\I�bs_���Z���
�c���$��dX����WT�]5ar:�����y��)fԅiuiA0���M��n����g!��G��C�劷���7v\��s�\�3&�^�]�ue��Y"݆�v�;�E\6�6A���qLR#�j��Hu�ˆ�b�n��b�2��\�.���Κ���yγ�_��fc좝��o1��3�O8��c*\�f�M]�^B;�/,�T��+4�'t�*6Y�̌�58sѿe�{{k/V���(1A����ەd:���P�0c�ˀ�1g��o��ꬫ�4��*��bY�}#�GqWQk�&'���}��[��33uv�q�˺R&�!K+%��(un��@��J�Z��,j@��Z:,�.�wʡ���8��^cP�B,�7���n;ǧ����X8�+��Xk��|<�	Yʯ�f����Ч�9���hV�0h[�] ����K��d��3��?�簙;��_�Fq�����ޝ���;Cg8�燔�O�����Z��K���˼W�:�ǋF�aBr;���e\
�;�؅�|���'PUݶԡY;���v�
��q�N�'�,}7]lG
������i��QIs5WM�׺M�u�hJu��2�Å��ᣚ�V��u=�)����������j _UԎ�um�ŉ���z��g�;�����5"�ͮ�xC��ڳR��Ϳ��K(���NWZbV��Ρ�C]�7+���:��+��ɔ7z�u>�z!w�T`8t����g�-�����po>�0gi�o�xa�z������B�qR���PȟIRL�.��5%2i���r�Y�t�6�ټ�
�гuBE�5�[7X��4Ȓо}�lآ�k]7Gb��.��u��񩏗v��(VQϞ�uG�;c3w�ʩ,p�K�T���<}��ᝁ�w:��ź$}̅�i�t�Sr�+�D�>WyE�@��yA�v��{�U	��KQ� ��j�6�
^�}v���_aT����,{�B&1���I%��x:ܭ\7��e���v�#�mB�9v��4���W���l���c7}���
@,��p��A9=�C��)Q���C.Jyi�	��bS8'c������X�gq�<��@ܢ�h���u�C�W,{���-G��-dۀЬ�W�B8Ҽy�j�5���b�y���� �^=�O'h��ێK��!�3-hbS��EBv���)��[�*1�VV�.����]Z���CsF��v�iYr�=���E�������0�]�f�`���-Te�R�)�n�٢���H���ʹ`�r����פ&h�Y6jt��}�􄺮���r��C�꺟t�ak#�X��ܖW�U|p�и�Zm>��;R��M�/ɤy�V�}�m/Fϊ�V�C\r�=(W�%k����i�k�G-R��[j�Fu�Y��iL��Jo�]�Cv ������%(�X���j��r��u
q(�ܰr���ս`�0)p���E�@��ɳ����Z�,�}�6e<��r5|Fl�O��i1tX4�j�^�N�e�MoS7���n�fD7�w.½�����nT�(�+wo0ʝ���aeI�9X��@�<G��R�
E�.^��f3(�<���9�ٕv�Q��y���l�ٓ���R�P��M�o%�qݶ��M\�X�n3������v&�]z�*����V�Jr��k�2q���s�M���=:z9�=�ZT0G�+����݉���t"Nm�}JS�i�s��f���$檴��ݚ���U��z*��U�폫5V4z0����K�H����l��˰R��1��v��Y�
�!�
�� �-�`�����|s9��w�u�jpej֕;��.�Z���Ϯ,_�3�i	q�޾�r��6�b)�4)f6��R􉱜�iu��K�{�n�G�h�ҷH�+ik���ܦ1gU��A�R1{g�Z CB�\���J��|�'�����d�obn�p���;%� �!����7�bOgv�m;Z8X�+�_'�b$Z&�T��eg����gX�\;�U8��
W�1�������\��K����7".��c(n��y�[]g��������[�����w��B�~�3�L���[�-]�^`J<ْ��ӛ�45T��"��4%���+x�s�����n��̞�NhK��u�.��bS��$c�T�s<�T����]R��=�;�˃Hڭ0ou�wSt�kId�hcHwB��frky%:�256�Ze��en�U٥�N<+�\ڐ��4�i�1m*�U�Mf�`����z�i���K�MH�T;4%���/�q�#i�g+����#������%:����Vs�&d2�u���̔#��M�Z�[ʈ���F�-�(-�
������K9�٠t7�����p�Z�C�l�͵�h�M-���	�J��d�/e88�R��P�R�.�Yû�7��\����h{2���O�y��f5�'G�H���+ovh��<�X�[B[|^������Ѥ��9�;�Z��@��S`�L�مopb�T��^We&e�{98�S�Y�\^�=W�iK��3��c�!N����^�+W.P����J#e��3
y8��kP�,=)����W��ns�&m���D7��9ݢc��Gt�w]ټ�#�7gJ�Q�`�"p,��'���p�P׺�ss�i�-�0��E/��8ȷ�㯙/2h�ܑ����bǶ�����Q+�9x��b�Nc�o�WV��s��C(ض��Y�7w���(��rV�a�D�����}nLV[��Y���K��Ww2c���MR�B�q�ƛDT1�׫N�@mf�7]v��RiT���0F�:`S>�z��&��rLc�1E�6��9LW5�;-�;l7Q_e{�I&;��M�</�u�3H��#U�>�چmY֐48��V���Z�xM-\^p���s�-���6i�ѦaU�;��
W^/��حǙ���ø�m��h�{N[��8D��X9^�
��ց���4ة]�e��\7����X�o��o�����kL�3�<��+4���i�e������ÇL҈3�B��q2�zR978�6l�w�:�nɛO��oc4!�c�v��؁��|�%���[;z,a��خ���$�1'V�K'S�H�5��p;�.hl���<O�� r�{�Фr���&�F;�҃M���=P3��]���8!��Ul�ͼ⸎�����r�pr�%�w�]�3h��4Z�F��b�D͜�Ɠ}�&�$�@H�.v��,| ���T
����\�����m�bv�<v\Iz�Ԃ��8�oF].�zb�[���hP���S�[�����̼�*TmPѰٶ�:���]���y�m����wJ��g�Hz�KLULD�UY�Wtx�P`�7a6��/��+���V�lݧ�Hn��Os0I��xu�Ī�T�Z3�.�`Nn���j�t_@��,�7l7�d���8�e-m��;�QT>�����Ɔ��t�ܜyA��,�f���V�ǜ��q<�m�fޚ�4TF�_�I��I�R}Sr��H�\�[,e�I����\�5����]�=�j�sV��z��b�s7z�x!��p�à���-�֖RѲ�u&9�r�-j��mE��k7��+*R�R����4o-ͤF �CGv5�{A[�}J��d��}��;l4^TU����`��b�Á�7�ö�N|�x��w5$���Ӹf��A8M��WKr�Lc�t�+��-�'Wc�ʝ5$�q�}B�����= �>MlR����u�2up۟gK{�E���2'1<��P �̬γ}�������3�z ���a.�=`��-�@���ͮ�4/M�����3��y�Ma�U��\,�3'�ݵ��S	a��/�ՠm����ن,�&� ����ݤ�6�t�(b�b
=�m)u}`����H��.�2�,6��I���l ���,hIل.Z�E�S�EV�6+�3��:��*��sP�N��U��HYn,���4�	w���H�i��.�>ޤ��akG�8��n2�9S��lВ��k��tA�d���j0Jvs4H�i��c��;�[4���	S93Vo8�wڊ�3�Xɺ�a��W�/1i$��&���*��lr%)����NCP�1�]�Gn0
��޺��Df���U�V=�-Z�X��f��f�MQ�+S���f=��\L�)����M2Id�WTa����]7qG��f���v�Ù]Y�Ԓ��a���t* ��5VU���X�����D��Y7~�6i>�k��}bpcP�`L�hƯQ�t�]�WM�̝�̴�PA��$4x�i���t]X��\�d��B�MŚSޙ�/z�Bu�d�Z+�]hS˔#��&IG]�@@�RU*���i#^�fٺÃ2��D�h��O;i}}*�t&��ʥ��oY�R7�}��gJ��,�#t�
�÷nouaL�K�1R��z�Κ��k1U��Yp�l��+w́��ԌR0qT���G�{���c�|�b�,�h}����%AԶWK����U��3�7�<3p�%�LT𔫞��%�n���$wF2#�9f��8n���RͶ��৙v�PS�b�+$�xvt�Q1Ȍ�$�WoRt��I*Z<o��&n(�X��w�༺0�W)���]E&�<xvW!Z7uݾ���+Kpn�d�VMl�xfN����U�IZ=��QK�BTk�)��F��HNF�f>9���Jbm��@T����dM�ӗ������ފ��ktT�rk���G�2�8`Vf�F_oWb�l�S2�kv���.�6mؐؕ�d[�a背E�-L�qw|�|�<�W�>鯶���ܵd���v��Q�T��dN}��9�V�P���m��˦��J7T|\�H�iNU��W�C�����;`��8%���Ξ���Twz�,�Bg_T�o�g;�&�ǌdr!���GI&�R%W��Bw��Z��k{cbb�p4����j,˭{pȯ����u��j�t^�495WuKb���괴o�3i̖49��2���̘�t3�S�K;[ ��Fȱ�u�PڥZu\�nfa�;k	�NFʇ{`ه��*`t�>��u%��E��ry���:��s^fp�Ҁ/dd�$47������� 瘇j`l6�Gwd�X7͉J��k�8�,���Wv��U2}KrlF��o)��a���o�zZ�#)$��>U��c��(k�0�T�_ww���f晧2N8�hQ��2��:��;0%˗v�����2Q�GLirZ8��W��];v��./V��f�{C��.��ّS��g*z"��g�C�Oa�V��I"�X.�cYnf���tYs��X��cR����E�{]!5�&K;G���eOq�F�m�6/1��f-Bwg]_�TvJ�8�墠Uǩ�\X�9�d';Cn۵5�4���)�#�dʝ�>[�L��M8�l%0����iI��30l�jv��|�nu�X^���|������q1y�9�Z�=I!�a�C�Lf�v�z���0n��p�+%#Ҁ\�l��t�������7���t��G�0�ײ��Pɔii��8\�j�g��0ۭ�:C���l��
s�'*��4Dd����+���1�����*�.0����-�{t}ݡ��R�c��K�[��KWn�J���F9ntIn&z^�Vr���6J�y�oWf�[�A�n��a��^bܳ�y��oN%����yK���i�ݭ�Q�^gs��+��1w����؂	�F�޴L��o���ިf�s��pU���I��&a�k\w�.[*Du�qnL�N�����8�t�C��+N�X����(A_/��c��2��lU1BXN��"��y�_K
"�SO<}w��g�y2<��� �*�#X�}�������7��G5�fuw��Z�����8�,���� ��������* ]����G��?�����������������������?��O�_�ǟϙA�EH�6��n)��*fD�
y��V�D��{IQ�l�V���F��
�V��}�����x��{pƉ�^���Hp[:v�׹0A�v���F��G�AÙ*T���S_Km�٣���ShRڌA4��L�V]jޢE�X��c� b�`�!Y/`�&!��Si*U@��ktM/OvK�Ď�\�i��t�ԍ؃g�r �!�B=��U,L՚�7rkK��fa���ς[;��Y��O(g%��?J���8`Ut�>�	9�,�;���06�v톅��^�f+xx��4.�7�:]�qsH�
:�.�/V�eg-��܈���8���Y�Y�t(m�T�]2t"��X:�<��Q��6�%���|�[�u�v��m5�HVV���s���;�]v�vm�J}Q�<R�E��|ik."�HfQ+��.�+\�#�������Z�Ug��2I���f��r�X6�X�N��M�!T�1��6ގ�F�)Wp%�.�y�ݷ�bB���2�����K�Rfc6Ң�e�5�H�]����b��k.�����m�݈�ƣ�u��$G�H�l�;�cL̄��i�d�WҬ�)�Хvb�4w��c
�]���y�P��Hr��ɶ��l��o 8���΂*i��ŝX郟gLԅ�S��+��Z�Y�j���=}�=�1�p"!�9����������㷷n�۷nݻv��۶v�۷n�v����۷q�۷nݼ;v�۷�nݸ�۷nݻ{v��Wf���u�9q�|K
i��d���J�8p����eh�*��93A�#A5�2)�^SUv�aӿld�owep�1o�E�[t�:f:�ۋ�;s�pSůf�#���E���ڽ����]�Pm��oi��[�o�;�ճ%[Z�]�u8M*�U�т�>�ܵ�1_iu����=�sj�`� )G`S�K�CPy}d"������c�8�Ǒ�\��2"�k;LK���;�-+�kj����8���xɇ#���e溁N �s���pŎ��v�;�r}�cH�#W1�"�	����zb;�=	kt�ȦE�n�[��ٹ��L��3a�f�Eֳ.����l�o"�2,H����f�F�s��V��v�6�5�"����k�ݼ�:nwmP���/��b���}e�0:��\�����6���}ʻ����b�h�8�F5�� &�Z����v��,�6:�M����볔�YԪon.�%[�f�eǪmj�(�*!><��G�}��'������� N]v��̍�#�7���Y�-WUD.sk"r�5��Q��Sf'aL��Tm�:��V-�{�2�+}��pP�ISJ��=Q��sb�V�dT�k���jH,�s+�W'�h]S�թA��������d0���G�^Z��vc�A�:����;m8�굊����.����՛�`�c�_s^��f.]pӛ�h<L�N�n-�/�qx�����>߷��nݺv�۷nݽ;v�ӷnݻv��۷oݻv�ӧN�nݻv�۷o�������}>�O������7{5:��:��y����a�/-�j,#�={5���)��p޺��ɮ�"4��a밠�K��ъ�eab��n����ׄ,�#%�z�ٲ��E8zcr�Q�2�����L�@�7�F8�ƺOSu��$�G{�S5��jЕ7F�9�Oƭ��Q�`���V���z�����U�\�d��	:�:vf��M��{3t�$g�*��"|S��;����&�sl�1e>?l�ܡ�U v=Л_f�뾷�`F�W^�X�&q_p���5؂H�_	<5��5u�v��R^p(�]>������-�j���E�;�%�ʭ5ð�y0J蕋 E���!�D�]s���>��`�u��o7K�̇>wN���rwN�j7(J엦9���|�n��]j�u�qI�Jێi�a��נ2��C�t��̖P���,��c�Cn�8��;��Z��(V�Ȳ�9�uHH1]�mV���(f�1���Umb��.��4�������%�wg6�<�i]����tc��bT_]< �j����GL5�L�p!��li|�ĝ�/�U*<q��̇�Mc�:�]�(-Rn˘��8���2��<۽��>R���`����1k#�\�7�����1|5�P+��ɹ5_7.h',�Q�f�{����}�f�b(\����YB+�Yl陽�K�$1�s�d��������t�36�T3x���^�Ƀ��B�1�X���l�I�pPw-�)���m�+;V���<F��������-�B����.v�7��S�<!5�&T�xB�7���h�ⲱ�lGy�Rh��R\�Vn��>�� �E�oJս�D�[��̓V F��Ȼ�o[�'=�˻��������k$:v�c�[����;���_fµ.Q����kXZ�]&&���"|Ee_c�q�L"�Э�P�z����
;������} ��N�]3���΂����9�k���b�`ut�n����<��6�#AU:��(�d��P�$ᩂ�VVDѬηXܜM���7`��2�mm�u��Yh���oyAWQf�9G��hZ��oa"N����<Q�l�qs�v3r��ʭ�8C�����%�
34�Psӯ���,��j�`�>ː8��{Ύ7���F;ѹ{�L� +�tJVt�N`�e̋r�kj��w+Y����F��,JLҽ���P�K�V�agr��R��q(+p�u#;����VB�j��p���*�ٜ
�gȥ]��eJ7��uI�V,�rGbZ�Z�U�h��^�g��,=߷T�u���h'ӝ�yc��Rz�\�,;���=�=�EG�vw��ť��Y�w�9�Aáe���M�{�l]Y;O/��TL�Z�햹qҳ�l���M��FP�n�p��M;�����6�8��k�7���Ff�Z���6#��F�(we������;�!ì�m�ג�UY.�%�ztL��k���{GW]�.�o������}CLJS��:��]� �[��uf駡������u�nwn|�u�ggA���Qo[2L57:���A�:ʆ��Yt���1X/i���ܔ�R���hV.]��l(������u�e�q�|>�按�1J�{l�T�r�����%(j��&�˷ԘEN�Mb�F��[�+I��e8H�鈊Y�;�]��h@U�{XvM����|�/(]q!�C��mq��A2
�y��Z�Xx̤�v�AFj�7�9�hUڢ�Q�2d\)H;�RW>�Ӂ7�c�ds�/e_G:;A�2�������5݄d�j��&4!����ݣ���@T��Iq3GsB�↜֎h]��E����PZ�L�/lgJ�뤇�V&���`����UB���g�,�ZWH��-<^J��m����s��u��8���O��b�9n��.B��}|{ �R9���`�r��48�eq���[��d[�G[�Vf��s*�w$�:^��ޕ����:ʝ����΂��Ɗ6�z�����K��Q�wxpf�ż+����D(�SwS;67@��dgG��l��ݑ:Ԩ��<q�®�P�n��&�s�^U�Y���3}�v���q�ᛘ��j�N��ն{��N���fZ����PL���O�����u�sn�u�¹I��>+H��+���5�/�Λ�e�Gr�e��^e�(��T�&���Od,v-Y�+���-�!R6���*�ӕ��:.�1\�mxU`1��V㐳�>j��ő	�C"Kw�����Wr}28�Yz��56e��@�o-�\�2�<��԰YtN��Im�v .)D![��T��]-��RWwM	VB�rӺ��˵F�J>�moV>�H��ZL)�N�<"w]Y���o����޵�P���;�sQI^��7*.��5o��i�Y��82�!m��@�n�)F�6��oz�v�om�a�r0�I����`����������{{2�f�V0��QB���6sakp �����YbQh�JtҲ�Q ��i��Q�h���5�����SY&t���%�Q+�GL�s�b�']n��f�|t���Y�'UJ�7x�Dڹ:F��4���c+�T!U,���'�V;���|*o<5�a<(q�9�9
Ζ*e�a7L�LSetAY,��[.�=�,g>eQ��y�T5A�����E��&��WՃ	��:ޝ�7\�ؒ�p/�G:C:_K� k� ���%N�h��n*U(��#Y����r�\F��Œ�+�fq����[X*�隊g��빑��-f�jSX�]���<v!+�������޸5V��}.m�_Q6,U�Whq5pD�V�?n&�F&+R`C�Ä�Y\1���޼����q)(m�R�@� �s��*�} ��8๼$ݷ����З��z�i5;x�P�n�eq��cx-�9j�S����;�nJ��2����7����ZPڻ�y��S�e,2f�q`��U)Ç33{0�&�^V���١����v&����i��BΥ��a�n8oE���c��*EK]
Ha���3ϫ�=�F���(���ĨZ�jt`��=��Q�F�[͋'³m弄�ʃ��8(M�����s55g3u;>�]�����պٻhs�h�ij��䠓,m��_,�4^rYׅ�c�e���.YZ���>�R��V �:���1��0+�r�̯���)�-��/����[��:^=3�킷.�("���]6%�:�^��8�d���n؂q�U�ӱ\�v=ܚO�5�Z
pIKl���9q�ZMy��)v�)� У���X��!������7lr���:�m�X/{*ۛ`����cS�喔��O��0e`����28+:Ĭ�i���T����(q�횝aŌ.ؚQ�hI��5��.�)Bn^4�)�����Ԃ�R�л6�YM��K;��[�>|q_ĚPMƞ�mU�ݐJ����yJ^����Gͩ��f��(}ñ�o�!�؆�q+2��O*K�Ŏ��*6+��ېɗ)su�K����lQ����j�{wbG�4Ԓ����g
�5@�D�Z�Q�.��,a������H=���tq�B�5�2��K��A
śVJ�*"^��A�f��\`�sA�iޭ���
H%�������2rN�(��U��ޓ[���LD���A:r�{_V8a��d�$�+D��9���6����,�,f�Es�YCT��sS�;X��n�s):��j=G+���+�Ҭf;8���ݭ5��b7 eSt6a����pG�tX����[�������_GC.w�{.+|^�Mw$7�ڔ�ț8n��e�=����`ԋ�Oj����Xc\�%9�z�ǣ,�7�maX��Λn�d ��������o�%xК���X����8r;���v���X�� N�`�r;H-ܰh��0��zDؓ�9ע��f�h�۲g5���KՆ�Rl�M�$�.��m(,�40V�ٹ)���}W`i�Ճ�`��S�G-�ך"�C:!��zh����m'HR��vݺ&aZ�gi|0$�9��<��7o��:�.[�W|;XT4K��6M�*}����"df�;C���ȉY�T�z�3d}�y��J��!l-��J�T{5|�c��J����.`�[�|>�4�3�O^�o�h��uE-���p�+dAb�k�c7�݄�;''���oS�t��4�h_P�om�d�L��2���y-����ۨ�մ�;܅�mBڷv�'%,����S�*�c(��9Ա������-=�ϝqF�F����jV�u�2�e*�@�����u�&��Y�9� �� ��՚9��(�<j�h���\�l�ͦ�+���y-�u�.I�o$�ˁ�	Gݡ�G������[s��E��\ �A���.:&��z�Y]�16T�uQ�ﻊ�8Bѓ�hak���Z{+{z.В�	�*�<��+&o&��c��P��ώ��gg-s���Fw��m@$oo.��Cr��7d@K��vPJ�t���#6#յj�O(Ŀ�ŭ-�������_*�/��H��@��i�v���m���PR;x���@̇��%R}nA�h�\�VJu3�^��}ӣ����t�ҙEYt���̩1Gkv��`HN��u���rVf+�1���f]
�+8˄P�"���cjf�YL�SpI���"pή껎�rR7*�Q��]n&�� 0V8p�/�
��]���~AX�����R�`���`�Jj��o&쫘�$�%A��ة����)+(e����=
�2-��v�o�I�8�]��V�1��3��W�9$%T�9n�,0��N�K��fn�l���P�Vҕg0�}����A
J!B����/gb�**�z (s$S������(��N�p���l�s��t�s����nAqԵ�3�������J�M��G���*���w�䦊��Q�{�o{D������*�WpɆ���Kwt�"����ws�훷�rqըTo6�s�i���:���97�3�������CRq@�
g���Fc(g��ųRiN�ecϊm�V�B�j��Q͌p�:���5�[�\�ܳ���f�%�0IH��g�Y���JvܧYC ��˦�XФ�� d���X�!�ll2��A�Qk=�����'y0�o��ή}��+�5���H�>ҝV��TWk&,jK�c�K�<������ji'�䕱,�S .@z��rao����n�y��5��i��ɜ�V���Hw�FМWQ�Kq5`��-�,U9Z�]WX醺���
��6P�%q�J��Y�5�+c><3�U�t���ì vY �'^v�-��۬�,.����v=[X�`�)�t�kF	�\���zk.�����ۑ�3*���+�Od��w+��S��z���~A�d��Fj�;���;�;����5���?ATW�d�����?����w��?����~-�~�����;ޟ[ޤ#�H'L���a Bm� ��]���Z��*��!��,�q��\�8;�;C��E��Ne�/�R�>y-�kޢ�m;�� {9$��(�R��z�Y���kb�������drĹ�K�w�����*�����y�T������rZ��;,�	RP�EeE�XCFk��J���r܎�9��`����}���7�z��udT7��]rl�֓�}�����C� ƇAu�`�2`��c7b�Ǜ�[,N���4Ge�ae�ca��"�X�G!*Y@��D��6k,�s�sEGu0g8w�q�ʥ���:��f5��@�P�]� .i0��H��8���:�V��Vz�G�(5Y��=۰s� Y��U�x}�t��8ǩzlPW	�Ὦ�h�2A]�^ê�	q�(f��ɺ�m�x7�b.�
�x
��W�*Z,)Vzc;dK�gLwM���MvV��xn+B6R�r(I�c+J]��'m�l�#u�r7��g+��a��DHuJXuM=�����uʥξ�V�e`=�k���̂��/�+�p5�z���T�M�3*,'o1vt髴��Ż�͒�����E=#]G��6�qn�r�+��w]�x�l�7]��.`��W>/i6�mVӵY�RAB:x�4=�v�6�nv1Җ� ��ιΆo(z�{r�o.�T������GI�!��<��ᷢD�yo;�*�NH�GbN>��.�ԑ�|2��@�`�ˠ�Qe�Q`6�StBT]�K����=	�H�����k��v�l#�����G��Lڞ&I��<���xus���m�j:�yR��Չ%��F��f8�������q5k8;&NsH�*c�3M&CFINf:��6��kNZ"q������"�����1"@�5!LLFf:�Z$ֱ�D�RjPxyDE6�ɮX������K��^U\I�D����=&C**�s�m��r�'����<�Qmp/(�jˮU�E�l"/#+ĝ��tO4���UV���ĊJ
i�b�	^�Ʉ�B�wH(��d�Q*3<*�͞^6��g
%I���R.�N�2�V�u��i�3"&b�FQ)̷s\kV�h�3*p��R<����J�/J��p���vz,a^m��=ҹ��E��+��'NĨ��Uc�I�jĉ
j"�J�E����'�Y2�93�b�E�p��E�yyt��*���4d2�Ȝ���I*��Q��0��5+UwZ�s")/�L�+íXi�l�54�#��IR4.C�;V��Ւ�r�.���t���x`y�ud�[�*`���e��I;��k�*��e]��["om��U_+6*��;�rs�#��b}��W]6�٥��י��<��
2XAw��½]G ����|���{}ͻ��P�Y��������xG��8OZ�6��ψ���UB<��+�(�
���8:_�^���'�l���^�ޫ�D+�P�4;�%��"����XMGm�d��%3_//)6�<��L��6 ����>y΂���Vf�^YO��Y�e{������]e-�`j�������rCi�7~��Fa���0����3*>���Z��a��Q6�
�H>�P��/e�w�rFWd%�y\hz�X|4�a(�����7��y���ʕnzaK3�n��"��.`r�}`W�֠���r�-��n�#�q�܍�b�Z�'/%������ϲ�=�ݏ�JD.�����U׹��d�=nԝr�9����I����*n�Ӈ^��~=K���
=U꾂��6]mS��-[R�V�fn*Z��癩@�T���Y�UQ0֌���B�[�L����G^w����W��Z�Sq7S���7��@����M�'sPv��sг��T���Ģ��mt*��H+���1�xP����zϏ5/�V�`��u9������?xB�`�>g&{�gxL�Z�~����I�\/(�;("��T!A��y����j�5��ޙ�f���.����1xy�K��=��zCV7���F�ԕh�F6��W����p�Y�ɢ���6��`�Ϗ�V�M�}7څ��R����a^�\hκ��{G_c��o���An}�c�����+�sw���9��^�����Lq4�*�,}��eL���kPWy���yU�gs���v3A�QF�w������̞�녠^D�h*#l��v����w:�A��r�� �_����я�y��쥈n@�|D^�VjO�(�6ʡ�����q�R�`�oB�F(u��6�G������c��C�r0خx�Y�zNغ!�� ��rmYs]]. �ݽ4/�����8���w�Y�쎂�UY @J�l�W�q�`�K�Q��7z�;�4�L��?#3A�3/���:6�pYN4��vR�J�r\0SE�Y]Ө��Q��+�2��^�nS}&8�ԤނË�6�X��Y��L� ^��V�Lw/zS�<?n����ޥ�3s=D��eU���(E`�;�]���Ǽ��D^��o�9�o���k��eM�1�Uf�����aK���-���3&|d�ߔ��Y�'¦5�U��k��$H�Y����Qf�}K�A�|��^��5���nH�m���)�wb��َ����)����n,�Sb��U�"��K��N��`Ďέ^�u\�g���#���TY��s�o�
a�Aՙ���	4��ط������_����؋�r�N/���D6c�1m�n�'^n�]�yZd���	��v�?h��g�v�T�9���u��3�e�[x׹�~�;=ק�b�R��T߹�Mn`���k��<�cm�SOOAv�G�}Y�^������.y�V����^�ھ������H���D$tL9K�O
�y+B�4���
�im �Q��qǶb�	�J,<m(^��n����Ȇ;$7���L�P�σu
�{�xo9�r�M+o������V4����}�Y�u��vۦ�o��UO\�_���¥t��˚y���}ry�(���d��Y_}��؊����tU�^��
P�:���A!n6�Fң^]�c�'�X*�#�w��A�o4=��O<�賢���Vkc�}ں�rK�K8�c/m��wFzr�P���w�Z�J���8iĶc�jR��I�}<������\޾m��l�_Y�^0k*W����:�7��XT{��J�"�ND��B�Z�ݦ�ˀ�u�N��t�P� ����ٝ�z{*�]Ƴ���q�v/�w��Ug"mJ��P7�u�9�1��zS���b��7:zvg��%	��g�$qw"זP�\����f�ޣ~X9rWԅ��-�J^�y{>(�ϩ_X]���:=<�3}I�}7ϓ}��^�sΤ��'�}j�Ƽ���w�9W�%�>�o�E��w�v�7u���}y��)\Cr �QOfN(��� #�Nv	��O�ss׃���kʧX��ȫ5q���H5�����۫�l���Zn�qǻ��&�bkvY"f��y2�\��H�s�L;PI��.�(���@УÃ�F���m��QTrP�e�5�'P�HTB�������+^�W��lw� Qs��V�l�9�,����{S�����T��|�UX�N�'�ʜk�}-gz6��u.��ͩ�e�{s�ܶ��QZ�x/An3b!��zf|�|8K�5;�`y�>�}�g �w��da.�WTZ1��(-AX	j"�z��d�q�����ٚ�1�cʉ�U�Dgf�*�}����佀�-�9�H�_���f+�/�>R�*�ʞ^W�~��h�a]��yOZ����=��}3��}�.9a�X��=�*�h�%D ���xc�;Wz9s�4�W�!g�?{ңU��`ޮ�ZY��^�������U��b5�n��$�ʻ-_�����W���nw{T+W�K���ܭ�
m	K��>�H�f�Mq^Q����!�Q�+^�m�6��]z�������q����m���٦��0\�8�b*�7��0L���&�Ʊ�)�k�{3P��W:6-��]����D�+�.gsT���,E�<�<PNbB�f]�\Uhw�QǼSQZ*�*ֵ�,Dggח[],�Ӯ�/�֚���#�p��2G�9�c%ӹ��{GzVN����0y���@�K玠��jE��a�Y�wdOݐ^������3�I؄���|ܻ�oݯ&�Ҝ��y�Q�(�<��'"=�H�|��~X:�,��r� �r��#"#�"��Y��DztR�r}��8ԏ*��ob��0��9w���zjjK�ݷ�C��Y�Z$�S���bQcޢ��-T��$q��ַ��W�)�=}=�;�>r�`r�D2c�R�wG�!�A�l�.���Kx�z��d�r�Xǈ4=�SI����_vT��V�@׫��KC>l{�:Խ���^k�~���۰�{�s��w�D�o��f�<ZX��p�+N��(q_��J�p����}S�g]u�kO$7��ݱz*�9��k�Mv���7b;=٥#�|6F��[|0+�S���An|9!���_^f���j�ưW�ք�cg���M^��G��ܸ�C�m�8�=P���Ei�H+�#\��@~Ϯ_[��b�i�V���y����&�-9�	�w!R� �h����]p��kj�Sn����6�B����3�� ��ι;�����|�����d��4e��? ��R��)!~ސ~00O�f�O��+��<y����)���ٟ>���B��>�Ͱ;!P���ʈ�)�W�q~<T���Jχ��@��˓�ߦ�]#��Og_ѹ*�>�FE�еZW��.sU�\�ێ�yg���U����C���y3ɼN��7��N�{-�3Su`O�	�yϳ�:z���v��~�2b��x��R�7�z���Qw�JWC�t#�����<�{��v/qT��.g���c<y�=ʟ�b>�a�[��5Ӱ�}G�?�߁s-���3%I������m����n9�&U�i�{�m����(._P8��x]��=*�w�vi�ou/c]�b�l>���,��;����t~��C�;�U�F*PyZ�q�T�z��Ut�H�#k
��	Q\1x�:#��0�]!�x/�k�v8�a53#Y�����նY��Q��gq�6�=����r���Nu�B+�`W���v�UO��V|�+h�dM�s#���"�ۓ���o�2�C.��L|L/c6b��-���YSZ����yZ�=b��r�k���%~�`ߺm��7�\˗r��#7�C`- ���qU����������� A��s��|�sg�`8��'�����W{�I��*��dG���m���+w��[\y��d�.q��]^ע.��7�/tM��W�����b�HjW�p�?��^�0*�{vf�z���q�;��W�*6WlY��xf���E�*of�/�~�A�&@���:z�[ƒ:��Vn�f�\�̓V�x�{����z9����у�>�.�;O\rK>3IbG++3��v�Q\B������;�"ǃ#,h
���Eg���%�QY�M����#�#ѝW���&k�>�t�xWi���o�7pOi��G�m�y�2ʻ9u���IATn�]�`tt�E�>�N�>W�Խξ��A�`b*6J��a�wf?f�]�,��t&(Ⱥ�PJ�y>"�c;i�*��y�؄�4��\^kV�כ���3*K�����ܚ��2u���T����a^��>�Y�"���/ȣ����UNBo��m�\q�G|�2������Ѻ��������~��l�K�=&z"}@��>��	��v���������_B�f�Gm�={�%fqF���e�WҲByCW� O��z���^Vgzzw�7(H���_��%/v��NJ'�쏣��
F}s1xR�3U�R~B�����}j�����O��(�J�}i�T���?s��߄gW�����B�b'��[	,�@i�c�����lY�Gw�\�
[W�ٶ����z���:Q�i[ޜ؟��������V^d��O]����C���[�3�]��{��꽋�S���W���]e�{�(OAXKP�H���3���[��:9��=]O�����Gog��]�V��佀�kv�$z�>�f2,:7�{�}|A�IF3^�=^��j���|�}^���)X�mb�� g{���ߥ]� K��#k[��¹;�\V�� ;�Pʐ�.�Ous���R6p���rHd�sO"�݃WV��	�!����{��Y�9�ڮQl�K�cYD�jM�>Y�%���h�U�7��B)���G9I�vuG1��*�H��vi��D쯕!��RB�o|E�|���p�+@%�6�RYw(����]�������U�*jR$�����7J�������#{�D]Y�v���[���Q\#���̕~F��Y�w}�u�7%\B?x-��;�fF�1@��>�R������X=f�"(a�Ñ��;&Nsu͞η/�m�*׭�g�`���k��l�zªEH�M����6���;I�P�H3��#Wo�gL���z^�r���~�o�e���Qg^�zBr�k���ᎁ���CƄO�^��o�������6�̯%5��e�g��v�3��1�·�k����tDX!z��]���3ޕpڢ+��f�yy�6��O�{���oZ&M,}|Ģ���mt���y�K_C�������7Ơ��<!a:[�9v"1��]Q('�O /���}�u�t����^��h6�ͥZ���7K��k�X��ph�|�,��0�6���r��Xn�\{�CY����]�c��a���v.�%�-��d�
Q9��0���}t:���7k91�S�6]꼻Ŗ��vi����q���p�9#A���L�*h7���b̍�� 
t�S6�ft�j0�N�*Iպ�=f�v�!G��b
���hlۇ:<v�8�Yy37jV�t��9yp��c�S��R��Sw�r?u�e70.V�Ʈ���^��c���	�G����� x�0݂�G`]�M��u��T��i-\�&�Y���pT��[Jѧӂ�hEy,Uܻ�+)5nniF)V�lpX�5��`2~\x�7U�<t��i=kwY���0uPN�'�VJ���x�m:`H6��(ق�p[�����vu�I���n����q�ޘ3��7�yb)��FTˮ�H��Q;�]Rր�`Q�#��չ3���k�ݮ嶝��5��{Fy���)ҡ���:fZ3�;����2��f��ݶ�]�^���Ela..#0d*����J��q���!A%�~�/r�����Ut�ꩠ�1��.�ir������jQ�fְ�Ӡ�	��/G����6��֙@��u"C��5yo�SM��V�R]iZ雍5H�9k�f-S�	g�G+��̏*��yX����x!������E}��
Q������!"�w�o�¸D���x6Y�o�D��!��_ACt�am���m����t��W"Ê,�ݎ�J�`�Q@�E�b���X�o
5�l4��ŗ�`��F��|��*ϊpt��#p�!����s��S��]*�>lVi�ʏ��\�$v�JEq���Y+TZ\5�\�u�V�ޤv�4Jn!��fU���6����f��.L�����D�+ޛa'�U�\��ʙZ���]�uև��t���r:\ͥ[�u ����ŋ�r��o2<C0�q�H��ܚ�_Nx���\w����'gn�T;^�0E!���f�COR��spUѕ�v�L��X�y=�n�"�I�jΝ��YB\�}r
.꫆
����t���S/�v52��!�M���g(>�ǋ:͹�wV��vKv�������V��\�4�>P�bѫ����Gt	�E/���C��T5�m�}��x�y_VD��J/�,��3���:3�eM{���Yv��)��U6�E��L�X�h�J#��wf����:�Z���+��K.9)PFo	�o8�v=u(�[���Mk�SV�+�L�W*V��w搗�{��^�:j����5�1<�����n��n��:oM���ͳRk�,$��	2�h@˘�K��C�/��kDjҵ~^�e�A��=�҂[�/��_��γ�`̆��N���rbI��4u�o���z����m��r[��z�D��9��8��P8�wQް�w���޲+{����]aM�ΠGU��z칍�%��Wnw.<�Ni�9���o���O^�����eeb,�k��jQDW==ٜ�Z�t��%[]��r�Z���Ǘ���ۇzZ��� yW��o�j8^��V�"�IJ��Egp�D�a�1Ƿ��������,��.�Z�d�T�`Q���ʙDxD�����ɴ�ġ�5H�L�	!EuOH���2\����C	W%I<\�b%VIUU\��36�(����猝=W-I��S��kU��њ�VU
�Rki2�LHy]ы��Rg��T2䪙k�ꑑ��GD���r��AI�W�Y�$*$'���GO3.BE^Mv���Ò�yZ����ĉ=:�!�P���6�n�CqT�"���>C���E�J��%���Kl��Ģ��Z�UK��c�/rjT�Nk��]�g��ZJ�
�B�S���d�(:�nU^z�Yۻ*�N`��	��pA��k�_u=ܘ£��Z(��ס*���:eC��-42H�^O�T�����o���_W���B�@u<�ħ�T_�;V~z�TG�'��'.���������f��I���ga�S����N�n���;�dEg�޵`o�Ϛ�R&����07�������T� �o�qY7C½��+��V�//�3ު��g����>�_�(�;&�9�{��D�c4�pU����<?}��y�*`�,�({���#��7�՟_-ǝ�����zv�X*�A.����(_��f��ي�3�>�g6iNl�f�t=c�
��a�8}�4E���y��/a�.��	MCrCj�������G�р�c���6J�וc���O�4kߡ�Z]������+ '���ќ�V�S4�>�p�klI�1�}[R���<5È01>g���s�)Dd:�q[�.����V�E�ǍϾUX�0hZ!��S˰�{D�)�҉1�5��/X�F��1=�vYpxߣ��w0�.����%�6�Y��<��\�/�V�w ��	��VV$�
�b��JGT�3>=y|^�
��@��Vpx~�	��s�"�5�k����%�s�Z�s#=�q#�Iط&om�M1ٶ�gg5>U�]*ح�@��i⽆�^�jp�ir��-eO�'�c�roD���d�,7�5����2@6�<��D���oh���P�� �^�4:��)�H�S�9}��I���>�7ݾ�zz���2��R�S�#�
�f(mz&:��&f!�F�2�e�� ���T������mc��;i��r�\����@e����t*
t0@\ `�L�������1�v��ޚG�C���NP��'�T��==3�}����/��`&�	t(���M��s{j�]Eg����x�E@��FeO��X(�7!h�� 4��n�F9#���"KXzq�&h_�X���@��K+"b�:0��~��_X�oGew���U�®aE�FdG�qH9o��o/i��=�A�=7�^F����$TWݴb�]'.�lvJ u};�� 
��eLo�.��+��ͳb���#D3��/᳷8>
�M 'Օ�IW�9tD2�xJN_�twMgG{�;c&!�6�V���"C��Bg���}�2��D��}�������*��M͎��f}�/Bl�{�j�/�BWE1.`R��`*�sѿ.��>L�p*1�Ƿ��Nԭ��0�n�I��[����A޽����!r�Xuja��0~�R3�I�!�J�rך��^b���+b��[T:����Elm
���~I@u�57��r�2�Z0����U��Y�CGw.W\����r6:E����-��[��zp�抳�nb��Q�n��7)�DFu\:��K�O�l���;ˡ��R$^�����;���z�d	�5v\� �P�`��,G�1�H�u^_����z�#������U����Xj��)���S4��z�����o�15)�G��w٨z��`i��xo���$F��ċ�!�T��J�����)��73��#��^yD�yq�b��K|��Q�S�>٨��Q1^�� 9a>R*O&':Q&�s�_M�ϓTE���3���N_��1c�Ŏ]Vg�LI��;�Mԡ��r���Ƃ��'t��>9F�O?��G��l��[mM�v�c�ۡ���Ub+(�S�(��Լ�7�^8�r�,t^K�V9Z��5h�k�n�S� �_0�V�03'pOF�?t��Ө�x\`օ���b�̽��i�1��(�
�9`�a�\:~�L#o�~	�S���%#:,��$�vlC�ߝH���d��}��B|�`������Pg�xf�g�sѾ5�R5EJY�����#j�F<���gDJT*g !P���8�P���;�����q���6!��0��s��8n+���]Se���-p���CbT�鹚cʛ�Y���ࣱ`��ո�/���h�^�A:���Q������=�Ҍڥ{�b�S��J�_"|-X��O �z�%�Z�r��:^��!Y�0p�]�Ž<�W]�2,70!��:fƲq��Nwe� ��;{����4d��p��O����N�}l��qU�*#���4����1Ѻ��l<����,B"G��v�SB�.�1R��ܖ�O���׏��+\�C�zOu'?DTgz�s��XcK>�]��`��xk"s��6��������$.�Ǆ�;�j}y^�z/�q�%�~�PC��`ţ��ȝ9~�µS�:������]R�5�48R�G�K��г1�����1�K��U�Z����$��w�;v����O�ӛ7��LS[�B}�.�y}�!ΌpX��a�{3hϰ�?o��7q��a�Pc��n���㡖��=H�0��������Ǉ�t�/?쪋�r���F�yԚ�,{�c�-�^����8����$�;�Ns�:*¨�_�N3^�W	Y����T£/.�I��3az�ˁ��/Ĩ?O������BhiF�}~�w�%�;�w�q�@V�p��p�w�b��db�r@�Z����(��U&3�"�K�w׵t���Av��&ቷ�
�(@��?1e㗫/�y/X�	<W9��&U�<�tT�������{�]E�_��K:G�����M��JU٣'��ޓ9;	(ڗ���#�vݼTz��C[i�Eg�64ۙY1��5��i�:%f��uH#j+�H�L�LR�*�wt��Q^4��H']�̝�r��� ����/���}��'	1�=s�����"F!F��������1F��o:|Y��|��t��e��J���d�ܼ�u;.�ô�
?A,�.x�g�@��O���{ro]j}R�>�H���g?B*�YW��s��g˶�Z"aZ�B�7��7���V^ڰ���q�m�ֽՒL9�O��B��ڏ��_ZTH;��ϭp����Vj�k�%@����N�w�UU]���v���h!��ճ;��{��|�
���}Q��bs��]x�Y��S�h�����kFdw��x�D�{�������
Qq|(��v��o�Q69}(ّ���| ߰1�5j�J+�pA؉��x�㩃�������괰U]/����C�ό�ܻ�g̷����y�W6r�p9�v҅Qׯ#���>�9~���=��A��5�F�h�)�z��=o:z/�>)���G�j]��݌�����cX���x�G혨h��W#�q�7㣊'��B�C6�����bl����z����P�:�A�X�%M �5Ͼm^C��c�ڣ���gb\���:�Cθ�,�y�븂�͚9�oZaT����`{����҇f�{��59iI�og�6���	�����l6�/��5T&�l������X����T-�VL���CRO��$��o��(W)9�G����l�|���P�M�U�Z�����I�0 H�����(�s�EӀ��,zm��+��4�ʪܦh\2X�bNQ�}[R�=��>�Skx����Q X����k�0s. 8��
���611�`m:rfQw����Z�=84v>�O��6 V����J�vYpxߣ��U�����u�K��'L�H�9�S}��Bsu��ayE��#y?s�΅�O{�ł=\kC�����^��X�F���?�z��(�"��#~vK.?��Q"x�5���;!5_���&���,Q����NP��
�X�垍������[7�c/Ѱ2V�$j����רw�˱��VV=�|���#�zo%��r����D�pU��:Q����a��Oh����;�dAkf��UG#�����$5�+aE��y�tɞ���Qϼ��~��l�P}�l*<nJ���T�[�bA|&ED��D�*qb���WP�m8$���E��U��c
��Ñ�������'V9�~��F`z��@~���WMˣ[����=�YCT�o��a�G��XCX+e\u�u �]z��`W���ϸk��/�v�Y�����FA;�ʘ��:��L���]��Ztu�Ak�Μ\�\�$��D���m�M�Y��J[����в��$g+�i�D��+�5�6�AF���]�6�o��}�>������M4�;�!R�����8f�ig�c&hx*lW�F͍������ګra��.�z������2$g���8�߭����'=װ�#"\���B����p�:�F&!�/WGo#
�N�O�Ł����F4Þ��Ô5иI�؞
�ϣ>}����b��!y�"��sל�9r����#�E���}��ez�|b�d��)���ځp�+c��ȕ(��Q^&f�X4bj�(��+��t��}޹�,[���ps�*�r��uq0)�v=�7����fg��2G������lS�~���躖Ď�BژB�U�`�x�دF���cS�H�71�:=�͌S��h�z� ���@���+��E���, �>�p�#~����*�;��ר���-��`l5/�M�b�`]xg &Q�> �X���>!a�����Z]��o5��l������`^�f�>ն�ބ�]����E�M�"}�֖o�,�K����<vHw22���RZ�`տJ��7J���!b����/�;�@�1�&'!��36^ʃ�)+M�}�ʡu�����t�QE'Ƿ6ƥXc�V���^+�ʚ7?WOT�0=��l,.�{�t���7��xK;Lz�7S+2nF��䵕yU��̮���r�B���j�Wb9w���ս�vX�yK0]oK��6&�o��
�������(sߞ祴��@��'�l@�/�AQ��.��Q�^�.�H:!}:t��m�JGg-R _�C���zXՃ���p���v:�	W�F �r�}s�� �y7�o���3Pӏ/f����;���/
��_�Sr�h����h��=�	�	��W�U�&����8d�A���)�nTJc�ou.Q�}���V�3�`�}䍯��F_�q��_h@�^4���6*mϠw�K#��K=r�s�Z��ޝs�Exr���N�Ѫ��9�j�jH�߇��szF���uQ#o6���~�C�!�I[����NƎ�&pwRbj0R���o�ϛY�l�˃S�/Y�;8�l^�xi�'�D����%t����5s�[uvN��!���bߛ�dO��eV,��%׋ഏ����ʗ��Q�Q�F��c�B���}��\��8����3�ӫ��lc�:��z�`W��������=1���u�iؘANƇ"Пd]����|��,� �U�����7sVx#�թ���ؠ8���w���N�M���fa�;H�W�s�R����^�6���^�D$�>W����mU]*�Bg�+L=�,ˊ�n~:/{ƾ��G?8��[�/' )��K,�Ϭd�{�cu��BdDVq҂��Jxn=hi�l�p9z�]�]m��S�w�%�yA%Тv_;���҄�m_m�nwќ͛���:>��T� �H�_DDD|#���Z�A�Ha��g�U�r���j_��Y>Mc��I�20N�Ӟ����D{w>ۇ��3>;L�'(����1�P��j�3`/V9p4�������>9Ps�G%FL��Z���b�]�l�2���0<6��&3�J|r�w�b�3����rcS�6�L`\p;��D�����0�g��Ū��t K��"z�/�u�j^��'����tc�
ȱ�.`uf�,��l�z�
���g�<A������r���� �fhǙ�ڌ�i���v���ev9�a$;����Xn����t�{��r� �>���s��g�g֬�GM/�K�9�X5w�.�i�2�'�r���O����8�ٌ]�	N�JDG	��S0b*�����1���K�R����4�RtB��	ϊ���*���nx��"aY��`���Get�{���$5�N�n�Mt�KI,��=��t؜	�,CR\g�xz~�C��wK�������5<��'��T�z�X��ns�5��D��=�Y5�^Z�����#���3�<�W���w��0vlT���`��~ћ��C%f,4�����^
�Kc+t"���;�gExUO�	Dj�o�nvs{y9��'e���� �=*Tv��H��u,�-�S���sZح�h|n��#D����q�Ʈ�w�:�:�~���f"��f��=����y���׼k�:��eqvPu�����ïW��:X�]S��3ު�e�#ފ�~�3U9��7��]�#s��:��y{���=9�O>62f�6(������߭�@n��7�>�7�Y�u�|K�j���!ƷV��V�� �o��lҝ��SG�xU�~|6$7b�5�Oi$\�C����
��e�#����Cj���c��Tv}�K�;2���i/r~B՝���Gwop�=�J@��"�@8�XB��h�	5n[�3NR��i�q�E�[���꒦����?V��*����{��uˮ`;�n>�m�rB��)�A��OpI��=�k&}�D s��0���@��}=@��A�+�B\v��dA��~�S�N�,/S�sF��g/Nzȉ���¨��F}�M��9��Y��HО @�@Wы(RC3�z�<z'�2�^�?����sH�X�c�jp�&qϦA���b�z&1��L詇%<5��*�M�1����N���],{%>�>��Ѽ����h���c�Cۨ���fb:������Ϡ�꯫���w�� ��
�.�(r�o���1v�����T��B|�=4��n~��L���ǈ�i�WT�7��y(]_bzuUwU�14�8�{:�2��[��\2��S�&2Q��ǯ]U� %i�آ��W2l�3�D7P:�+ J����;JN�U�/���b�P�z2Pp3�C��.W'&�ݖ�)vU<"��1������9��jl㛍l��lU�5:�X?`�ClA*މ�c����)�bI�>�@r�Fl���ua�>��z�3�.��}z��Q}۫Z8nRo^�/��xY�u^#j�8�0*ޗjk���k�E��V��ZxX�y
�92�ƛ�9Wl�-����[mQ�S,[M���M�y.�F����&�?uieN5�9��&�]1r�M��unP/�5ғ��i���P���{�m5���F����88��&�k���mn;�t݆��Iv�0m������=)��"䦽��0�8��!�X�tm-�{Z�v�K�:���N��]wDj�̢���tY�;��5��c9�6�
Z�_<9B��*ƚ�&���]>!pm��{��:��[GX�X�Ź�N̺��y��u�
����7��!c�B���d�)��}��9�4(ek,ob�;3z�_V?���}���l�/wdb�AFL�E���[U0�i��j��k�3��Z;>�١�S�������T+s#�����g!�gRm�|�q�Jm�q�P�F�'�28/����]���U��'--I��da��Po�7&�"�.#�mcN\�-�T+;Q������h Ȭ;���V�ڕ���镰߆V{��'mjN�Cو<I:ަ��N�*��/+o���1f��c�9!D�G'�����C��f:ABv��4a;�
��NKPۃEaZn�»,�y|���"�Nq�	���kX͍Z�愨�T���w��U6TNF�4�`�e��tYJ��Mz�SE�ķ��� ��±B���T�^��|Vm�y�G���c~1;Z�]�V���)FB�+���)aGa�U�׼��V�`�-\�����w2l�;��*��S�BW[V�l��z��
�{�J;�P���ٝy��lrVA7:�Ζ����D�V�����k{f�,ՠV���Ƌ��R��FyrX\��V�Pb�$-�r4)��
x�e�B��cwc':��g����� �U��Ն���n�M����ne-�"�⬼�t�;R�%�BmZb�n�YZ4�}��R�����]�+��lԌ����+:4��Ա��l�>'4]�uZs.
:���&C��S{)Z�G:ۑ�<8�NA,�y���%.
��1���N�s�ˣ�r7@�k����,�X���2͋�8$!���pv��&Ҿ�R>4���9"�̹pV��HX���9�)�͠��F�.�b)��`蓒�/�a�5�h�����y���q4�Φ�˛�����'sۊH��QP۠(P9d������~��hhJ��NQW�����r������60J�q�����U�QNE���+�$�/#��6�XхkZ+VX�VD������(���Ҧ.M�2Z읕)#��2�5���"��!^lN�l��^EDx5����&v���̉��z��.J�ԅ��{$��	հ�L��*���=��90錙*ɪ{�@������g(9$Q�3hQ��*�3$�s�(L�&�%���Q�\"ri��m��$5"E7�6�ޯ@��<�
d_j�=��ކ�m�N�g!��7"�״�}��p�z�d2ol�竉�#�=��}�9;R>K�b=�޵�p�o]*g3��yD^]JvT��o\�93�'zۼ�L�;�]A�qd�V�5j8�f�F�.��o�6=a�r��v� cY��v!6u�+Dp���96&3}�$�����k�0]�{&�`��x=��	�S(�F�?:���0���Vh�3��=J�"�Z��(�i�j���y���u�T�F���|���V1�.��B���(���-VQ�'�0Cs�+�ᮙbI��'z�~Q���e�R�F;*{<V
9��[�5y�N,.��v�k+/�[�=r�vT���7� t0=:&GD��"�Lx)Q�t�+E�����8$���^)��=�֝̽Ƭ��t2�Ͻ�b�4fE��N f�i�X�� Lp�1�WM��7���axzG\���{��Uؿz~���N����Lm9�n�F Һ���s�5;4�����
����>�Cs2#$c�غ�{]�B~�[��5���ߡ��I���q��[�U=�����銬������^�Q�����]�_uy�)���i�������ќi�=��s�k�p���z'�F{+jR�����x✉[Y3��z~~��SNc~�}2�L�	4�?N�����V-�b������=o�X&#�z��?���/6�B�t}AӸ�Ⱥnc>�\�}n`�N�UV���<f��/FQ~�WIۦ�y�Hݮ��V�,�ߣ갅z.��"��y���U�g��d����q���P<=u�=tz�fn��"��k����'r[Q/�^�{w����V�Xn�'���f`۸��^ӗez�T��/.X%pʒ��N������n���t�7N�킾�9�3v��Q���nVZ��+^�O���%�1�S����B�T�4�KAB��ϝ{���b�����}�:���3c�	��m�1ɨPa��o�(9&� ���a�;��'���?�6e���<�b��Zs�����M<�X��f{�f�N���N�x�sۡ�O�p��]�h�D^��r�<�^V�Y���j�jl��BϚ���ET�z����"��1�}��Q�1��z��
�9Xe���U��������f�+�}��	��?1u���ݵ�9���D�r D�	0�@�
$)p�X1Ǖ�p��G?�})�S��7���c����eZ��c��P��F8��)��@���D�u�B|�`���ǭ@0|���<��z�*nP���q\66G��a���`k.g���S�%Z�s$)�\	��^����էs����Y��X|�@ϛ�S�W0}%UT/	�]��<6����IV��	�#�2�̀!��ڿxy�ڌG3��Wm�k�����\�"$�C��u�V�3Y5èD/8\vW�^�Nǽͪ�F	c<'vC�zڝ����ou38;��5�L9oh1����P�{����z�|Į�n}�M��v�D�v!zr'�~5dxh�WW��W�:N�"�{�,jՄd(�ING��MAu�u!�w�K���2�"R�%H���%rXI��b�ԬȨ�����N̽��0��>L�T�"y�l�+ػ��K�* �W�B����>�>� �qN
�%�W;Rz�&�W@�T����:/+ч@�eǣ.��к����-}Rޫ�����>�@�k��?�^
umDvV�
��K�R>X�>"s�����1�K��/���3��;�����V\��R�{b��A��g�A٫���dme�`}�AIfvHw�V�	�AQJ���r�z8�ҕ�n�v�x7Ez�Ӄ��4�6}3b��6'G2u�7&��S�^�w(���=�!b7�uRR���j_�e�~�5�I�20N�Ҝ����k������2��}�7�0"2g #,��/!B�j�3`��ˁ����s~ �d<�ʃ�Q�Q�ȧ��=�׾�g��=����E��H��TGE�`���k��9��3��S�L�B�O�X�l��z=���_���q;��%A��t.��/���K�3�O�a]�+�fvAW�~iTN�>3����~��Td�="G1F����"_Iϯ�#����Bps��\��׊̫���̻])�S�+��.#����"@ КQSb�:\?"L��%����`P�\݊~t)M���i����[��Ȱ
��#1�q��p�s]N�'��R����(v�JS���^�Հ���DӅ���U9V�U�1a`�C����Qvˌ�ή�v+UДT�kӺ�0�_>w��s���}��7�����E��&EB%�I�yyU��s�����-ۄ�����R3��Ү�`�m�,U�&�B"A
��ITn����5����A
�_�6��U.N�b#�i���?R���}�V|�M|tT�w�O���y��$�^���Y�4�T�����V!/�vz���bq8�ŋh�F�b�>J<���r*<<��n�$�?1�YS�=WD�����Y����ؙ^}4J����^����̭�Hž�ּ1'������9f�K��|ge��
��pc��/��l�~q����o��_�_�H<�w{�A����3hC�V�Q��mv�����>���3B�w�F�h���~���\�{93B���2k����.b�g�R��
�!�n�·��5���ɥ>>��D�p%U���/ ��/�PDK~�`�0I�����l��VmF:����gb\מ�Uޫw�������hu�Y��g�t`,#���/M�8$չn|����͌���q�x{�.�8�H�z��?��Գ?mQ�Dw�e�>�`;�nd_�q�s઱�c\�G%��gޠ���llF-���j�B�^�7S�%�e���;��]�VK���3���S1c��b��3f+ﲠ�@��ٲ�9�{��r���;0����kv�MƦ�/J̫
En�.�&Ž �����x�f����l����;��S�I�A9��{�|�߄�rD�w~�@q�r�)'�������l1_T�N	�"�~�8�����&&g��5���'��H]�3�Z��6�j(��
���?O�-�Ȋ1`T�dX�fa�A��W��Y�^[���И�1��ڛןX�W'��)�>��L�^��_1��L�5�h��\	<3�tq�*:o�9Z��B�K=�m�1��?Yw??�ߣ`d���� l���E{w���jzA!����7S
Y� �A��y�ע]�*�~��;~�Xc��?;l�d}syϯ���L[P"G��K�F���)�/�\���ycr�j�����{T�}V��:�{O��{M�z��q�&�
�������aZ/�t7�ę>^8.�O�B1�9}����w��v3�3s
-*3"��Z��٥��\�$TW�6�}8/)�{j�e��y◲>] �
��o�U�J ���숤i)��C��u��of���4<���������"��srx�Q��{e�Ϳ�ں���S����lF���y�;����������46��x���t�)-U������^��r�ۢYs.��$�ާV���;$K`�,��0nQ��R"�/H�M6�:r�eP7�0���r^�fo{ϻ�q��<�,>�Q��g&�l��xl����Ǣ�s�B�0��ѝo�7yߟe �`FdTC�o��߼q�0O�����^rj{� ��	��՞�i�=�a�k�p���z'���>{�E%#"2���ǋ�y�J`u��pT6Ɗ�#�Vf3�W��>�S3�i�~� ��/G����&���HC�ln�!���l���-�Ƴ��`+�K��}�y�r�_���sX>�0I��k
�;��Y>��JG���X5��NF�u��ȧ��>�a
�]KbE��Bi��#��~�0uh��y8>કt�1���9������61�eXK�;�B��g�5�=B�a����~>Xv����%��Q�y�~C}X�P�^�=ɋ>�ns@.���4%b�+�<�w�epV�T�ר�WR���ǟ���N�js啎V����G�8�/[3q��ڛН�X�e@��b ��Vx2.jWU�q�<��7.D�o�㶨8.p�a��=�Vʵ�5'j�l½ǝyw��5Y'j2�VV�'�F���3�Ӽ���a��-�廇G���c�+̻}1����Y�Fc��,�����D�þ�db:,�)�2����D��1t'�UuL>>�����T!V=�%�W3���ݣ���:I��]����	�d+�U���I+[�l1m�)w+HW+um=�w{Zg,g� �;_V��E�5���-��T7���j�R�L�vMAi��bC�v7Uk��i�:u$"�S������c��Hr�J��!��ru��  ���_G���~�I�N=����� ��IS1[�e��db�S�%_��̐�Np����J�'��jQ^������es����?b��U��\���]�Z�[	}�+����M��*�D�����oޗ˵_-��� C�3Ҡ:{~�^'"{լMg+		�9;Fb7Qap����f��Z��}���u�>�E��DP��)�+޾S������gu6&��0�������7�ޏJ�+�l���u���b0�ϋ�j���({�!^I���{.=�.��],C�ރUX&0
�H�L�<S# ��T:�Y���ѱ�_�U�R�@�г1��p`�J3�Tf���k*�����y��zkX1΋gҮ��t��,��������R���ڟYy6{/����L�Ls�`jVb������@q��x7k׾��٧<6}3@X��.������ϯ���(�by��aNk���vܿ5pԿ}�|����#��9��E>S�,�>��j�Q�P���,Bż����Վ\/-�~3Y |p�	oI����0�~�GRצ~y��z��B)�,�=��ㅕ�:@�f�2:1�Sw�mV]��;>�O���1=C��R�n�ͩb�H��#w�Zp�4��G��-V}�Y�G4��:m!ٿ ��jS���i��;�k����wϜ�~o�U>�Q&AA=�c���s���n?L����'"�
�=N��`]���̋ /<7:���5��l*Z��'w]ƫU.
�|�)п��?�р���o���qT=[����`-s����0��d�fgWR;Pl��冫���x	�����Q�$��\_T�}'/�#�GR�2#.�fc��ej�;f����垀���NI��c����@g I�� D�	��;O:w�Vž��I_Y��p�z���Y�O-�G'�U�~�]���q����w�;�����{_�3�H,K�µM��s�5�&I�";M%$)���1#��>�²{f$f�疞^���|�?��g���"iV�������
�vz���8�yǎ��������(�gt�@͕P��+�����mJΫ���S����R�;�Y����'���� ���5�Eջ���H���_߻z���Pߦ)�:�6�+��j��:qb�^�[yY���)Go���緆��{�:�* ����r#���]l�Z�����7�f&��¿x��F}Ѳ����S�A]��*��1G���݈V(��T���:	k��!�#���k�i�lE������k��{HV��ԃn*t+'3����]��$�y[8�,=�פ��Į9���E�Hh7�j)w�!	w�o[�מ���~o���>�fA R)�my�����և�8�5�՟X�� [�o�[�5��:�~�ئ���9�Jv=2�P�������<��.Շ��^��D����>�ey�2Ñ�9y4�Wڷ�Gg�����b'M��b�&���'%�O�hX��Vf#�"�@x}�H�	5n[�*�r��p�9���p���{�?P݋��z.�0ʖg�#b黈��D<]s��̋q�s�+�
�ӧ�F�*������^3��j��=?O}9�1_B��$xߣ��g�f#�1o���h�z�L=t�R�rZ̈́�9��}�\
�6$�>���*P26���%�»&�*�a�n��Z����;�pƾ����]��S��3��D��o�I��ThX��׿<4�%;�S�w�u1��>Y��Yc!JW��m�1�j������yw�[3՝ã�rW�NP����z���O@��ة�%� r��`�p��$U��:Q���Z�1�n�����`������?.&�b�(���_T���`��ycr�W���ѝ�������ѣr�,!<�A)�ns����9@;�o�=�U���u���rY\KEV^���5q��;���|d���FS��꽪���}�s�����X�����ٯ�G�Y�F����l��C�%��z��ڽ�E�����>��?�EI�T:��{��w�q�w���g�� �*8)�2(�������(��~�]C��8��-��|�/}�zG{=�W�����B���)�\*��\'��7�KX�� LXdz�e]c���I[�T.�c=\�$�^�S���@{��"���0�l1WQ{=�>3{4��d�}�]���/i�����;�w���h�������;�:0y�bB���BM_�s�{=Cb\�eTF��k:7�<5��� �\����
fo��䃂]zoaq��j�aι�9蛎��
�S�*{ʶv��ڕ�"23��V�{"���w��z��i�~����/�;3-8���)��}��!��c��b���VǺO���V��P��|M���n":�i�Eɕ�p�]_���;y+��,��:�R���n�9~���V�<�X��tL7�BA�w�)?`�q�)��$Q>�u���!����ŀ�,��4&b����X�F�N	�l���0��Q*��a�o�z�a�Q8�,0�>�p�jy1g�m�iw�Կ|����1a�l:L�)'���_�Jo^��M���-LIW���U�m=��S�,�n����t��$���Gs+wF�����g4���a;��*錭�����z"�{@�B-��$T�))��Qp5����Un<e0�H�gRy���J��e#h`��Ϟ�l�$v�T��5W�Շr��틫c� ��k��t���K{/�0�Q���Ç
}4;T�;=��w*t+3_r�YO�Kf�s#��H�����/p�ێ���R�3�7�*U�,��1r����HS\�;���j�!�����YT:�h��2�Txc���Zs�?�I����Ӫ&u����F�ok�(Hۘw�jۨLh^�43~���\�%F���U�J�)�8٭X{�!Pe+��j�B�*|���#\���p㹝D�͋�Ҙ�XK�/�䡿m�8�RV�h��x�%e_T�eFC�}�}�Β5�B�V�Gm��%�\@�N-t~2�]b]Do;M=�p�ʶ;�
���
���ji�쫛�}�՚W2���$t��HFU+�N]Z��/*��[�񭂺�t�F�_l\75#�������]y���u!�r�@�e���ɻv4cb��|E�s�������x�Z9pn8]�����J�x��CZ�&�3�7�n.!K �uQi\7F^Y\�k�IVQ.���@V��	�a#�\�X�N�Yjr���[�\�X��S�cy��rf���|)a�ټ�OlI���ƛD�P��9q�K�#�tB�]��ю���x��z<�KYSdբ�d��Qq)1��+�\ך�:�.t�(d��G�%�2�v]���ڔ����Z�ЗW)�-��Z�>_ ��T6��"����9O�P���Z��ǜ�"p���5�wו:�ui��R��>�{f��y��s5�8�"��N&����*�ma�ۮ������g116s�Wg[�e]=� .�	jR�����7ർ�� ��=��.�V\Ôp�uˬ$d��{�fU�%���Ʒ�� �:)��� ��@��7Hꛫs��.ܞ[��X��Xt�o%���A����Ș�A�,���-�"�s��,���#� �e1��ݻ�4���Ɨ;p�%^�-����Tѓ/;.S[CJ�-Q�aȌPe�M� �eE�p���=�`�J�X���RD���ל�
�Q�k�����L��L�{��e���%M�wF�H�	�a���xfnǴs�9M�)5�u��d����^�6��]��$���Z��ke�#&��o�1|{s!��MN�B�E�$�@��3gv�6AV'ک�E��;��h�;�ma��x�M�ʨ4��m���2�a%=k
��j�q8�=�Vxͨ�%��:������C�9��:T�Q�����[8������ˏ\蘫�Ϸ�܀�W^f��`�ܐ`�3��ِ�Q��Cv�n�~�¼�&���N��@����z%C�+�yќ�^��gѲ��G�%l��r̔j�͗<�Y\鞞����-Uј2O�/�ȥ���v�xux����hɽ�xɚO]�(��OqZ�Ɗ5���.3Xk��==<==/WR"y��`�Oo�"���rל�+`Û�)A3�'j��x��{#�Bc�a�\�k��ϥMʼ�����
z#����h��VϜ�y*�t�׏^��u���&ԩ���<'����u���.�zܾ�:޼>ۏx�I�l��׼z��p���[W*��$	]J����'�A�.�h�y�\�����ɕG7z&�y�Mޤ��0�5KY$��כT��-6l�T����;�ݕ~#̒|;�<U�>)E	jz-'���oc*�b�OE�%U���"r�k1����C�*�0��1����Tٲņ�+��s9ك;�z�t}�f%#���W
���_UrJ԰��,�
�v�5 \|?��b5�L�+�+g�9q�#t�pcb��T�r�U�igt���[Z��$�qŮU3t��j���Cj����}�V���מz
?L*3 �����wŹ`��F��B>_B����V����G�8����j�jm:0Xk��z�{�":���s��fb����&���PPT���/@Y��	V�F��@@k6aZ��CS�b���w�V�G�A��yɛ�7�a�<�/y�<��g����Ŗv���o��N)�U���Evs�-�*v7�n�����V�D��Q��+��0��'�W[��g���ʠa�x�f�Ӡ���g�e��F��Q�%{�b�k�	��x��cʕw�K��c��N?��a�Z	����P
�3s�UUG�\+a�ܾ���;U���c��<OQ ���{�`Tۯ��+��	w\@?{ըMgÕ�����b,4n��
�u����S��i�q��3P_�B"~��.�B�ȿ�޶�o+};�L�wSbj0/S[�[�T`�C�������7v�?����q��mI�YC܍�x�E�z0��G�q�e�~����)�㺫s:��r���dF�}����o�/n��`�ȚS�E���O\�3ن��I�C��l�8�O�#�KYqJS�E[�<�����iE�>�g�!�1R�T��E��,�"��XbqaL֯�6��꧱Z<MjC*�V��y�֩���L�*���	�^�._�.Q�Ef�����ei��y��7�|YI�6o�5��<�~q�E�"�ʊ�~��J]9��Q��t��{R��淃��9�{�%d�}�͚��'bb�u�nE�>~�^���c-`�@�7���P��� ��Ϙ�~Vb�5n^�j��x7kר�-�tqD�p��3� �b��ͩ�g��S�'����Aҳ�ݷ/�M\5/�k!�ɬp2Ma�Yێa­��������z���U��uK.�P�9���Ѕ�v�V9�Վ\/-�~ �d>̍7�㋚��Q�:��nzȎ��9U���)��rÄ�lZ�,s#3���{���͈��/�T��>�S��3j��"�M.�=p+��8�)u-+c�?���Qk3�#U�D��rutY���1��o�k�e^�x	�~��Td�="G(�W ��"_Iǋ��ϲ%�1���l�J�b`_a�����@�;�N����tn`=ˈ���[M�!�D�nݼo��Q���\g�����5JT?�T����d#IㅿC�������g#�[��&����c�|�VϬ�@�Bh`��u6��v��I�����D*�В�AҦ�����~�;vf��OuB����}�fi�P~x������n�7rF�kV�2�"7�ں��z���x�]
%
�#�\}����S7�m�F�*�rAӉt��-�*K` �k�6�_d���B�h*��itȬ�*�}U��98^[�(Q5�O�E	�Q:����Ͽ<�ӭ�Ɖ���2?h������B�����t }W��k�z[_%�u����9���򈽧�׷+��\����ώTX3�g��G���U�^:�~`����U�a8U}D�o\��<�<g�w��"�Q��O��ժ�7��������`9X(�ņ8�O�Q/��lu����_�Wu\������]�0�Dr�b:�k�����w���0�(mWg��=��ܧ+�e��|�|��n��7�9�
��Ϭqb�x�b!��9vk`pF�Ӄg6iM�<���>s��_���\싰X��0I�����nw���=8��o�X댭
ho��V�s|�gcc ����E֪���׈����S��ќ�V��+��7�L�8���o���ְc�����>���@��QM�Gge��U9�S��u^�+��n��{�.;��.�_G��_�C��-��61`}���T���� 0���
q��dA�~w^���`�{*M�f<���b�~��u�K��l%<�P'�o U�lI��
�:1����{�[����T����Z�!�v=ܛ�C�J|X<���j�c�okoF�H$]��R�&{�6��,����ԧ��?'d������i��m&�9�z:��g0��O����4�C;�fS�_eI|:�#7�H������eVd@���y���}��vq�����N��א|U�b�36��c�T�tL�L�aU���L
���f�uG����*�$Cŉ���2��e��
R����mɍ�y�[7��O.�=�0י�}f���iJf�ꘌcjO	P+�%���c��Õ{><�k�.�����to����w�ĝ��g2���L�����j١HS��_�Q���}K��m���6N���<u�w���5�76���=.3�:&E f�xI���t��]?J�}c��b�Ȓ
 ׳���>�$�|�ϛ�S�W0��*�Ȱ
�&+&�ˎ�'�k~���x�ӄQ�>�5%��D�3B���*��=��{Dw�ZS���i]F�F91Y4�_�&H�y%��}i��`��3D�'ka��y����F�lH!�����	�؞�`l?Z�0qƸ�Б�(�CbL���<=#�T���y��}Y��,9��Ss]�B�Ff{g3���pc�ilK����J�p�xj�~���Ep�v��o-��0~�?��`�~0���~7SV[BHx/ܴ�X���M�D ��7�#k�hvR��&���R��+�T�]U����n5���mAko��h�F,	T֮ڰ�"$ӛy@L�}��E�9v#�XU�NGrn�۔����M$����} ��#0�/κٞ�w��㮈����ż�<�#;~�9[R��DՊQ�Q*[�����q�O�vtR��z	�N����.�q��U[����<��l�d|}[�z>���D�bF����3��߭�����A�?�ȌkW0M�p�HpWER�+�F�N	�l��Q�5�I����|Vo
!��V��p�Sɋ>�nsK����)�c���<�u,⇴������õ���tb��艹�D��0�>9X�j�`ţ���fn3V�Sz�`��_�sU���'�PD����&�Qψ*�}R�
��ώVz��5h�t��x�\�bS*�b��bUZ�ҩ�ѐ<�n<�p-��rg�.�3ȋ�yu�#<�q�潾r�c��Z<�]x{;nR����g���c=!�zZt��h�IH�΋1�tL�$lƽ<��tg~�ήvg����ӋZ瞐���W'�Lb޾�a���h�o=:U1~�
˃�S�N��aX��*�}V�ڱ,k�NZ�wx�@��)�50�S�A�/b��9�cS��ӟ'wQ>���ؕ&���s�}�'ވ�D��3�ea|b�VV���6��]����mJ�ȝu�/�[�������{��z��Km7�a&�JD���*�dǳk1��0w������&c�	��ܕ6��@8m�rd�O�,��C6�4��sÔ��-�_����VeP\�������w��pq���F��]M����o��7�Z��}��Bq:E���w���Nך���M� �2��@o4U�W
?�?
>Y���3D������a�����G��w���'ޡ{�X�u�>��`�m]39~�P�/�TdO�&r�JX������;���8�j����
���B?{-�2'�X��ڈ�K�R�0e#�u�S�6���L/�d��R3����w���
0*B�x���c��}�t#}ӟzsf��N��|­���ޠ\D��b�~7��X�¤"~Ϩ������%�p�)�rӥu��_��:��)�֍�ϰ��̗�y��W��O��9� *�<P�,!`iY����r�����d^�O-�rL`~��m�׸q��f�ļW�Dz�g>9HB�!b�j�3`��ˁ��.��	�lz<�Z������BS�&"zXu+b�:��]N|rÅ�w�b�,s#;���o[wU&�'_t�w}�ܶkT�Н(Lҩ0C�r&��� WƄ	q�`Q�s��Kȋp�Nٯ~���ٔJ��wmj!��o3Z<k5#��B��Pe	Z���h�1=R�e�OQ�H��k9f�/�tT̘H���c=�j���7Jol�ږ���$��%�\ɝ���S>̳�v����tY��B�RW5"!s����������@&ׯ?>�q��׾s�ǰ@Z�q���7[x�pk�e^�x	��g��z
�t$S` �@5�ʧ��-D�s���n}s��yo��8�r���4�{��)ۛra��G�rpL)��wiw�1m�9�:~�~��Xf�L)qb�S��󽇴�8Z!ч.���w��p�W���x$}�@�[�w��+DL[(Dxt�����o��t_T�9����jHR'�$����ب��da?���+�H}��
��/�u\�1*�"�[�S����ߒ�
���O�_]��w�W=&�}���� �Q���?:Ԣ=10U~����C���N|,��u>��
U��}~���5X�z�dE`^�c~��5j�M���3{5�q5��\XaӃe�#1Ycn�}{;nu�K��$��ղ׮������f'~]lC�w�
06��}ծxzsf��s4��3��j����2Hca�N���_��E��	�M�︱n=�[� ����~�����/m4�ﰸ����J+��M)`35�!P��U�^˛�' >�`�<Q�i�#Up��ͫ�{ڻ�ǲ�T�����O���42fK�=�L̼�a�N�B`%��O��	eU�vS��n��ġ�ɝC��P>Z��G9ͫ�r�q�[�)^��&K[@��E`-��t5û2�yvYU:	JF��E��j�%bY�mlWQ��M>�����Txם�>{���k˾�����9ί�v%������:�1Ϣ��g�Am�4��6}�Y��	���=��OyP�L�8��;f0O�j^_H��#b[����!����2�S�oFvET��/ê�zZ�m_�Z��)��O��0��>�����+���P�v6�WvT�B3.�m�Q��'���c��W0WS�s�:�%�6�j(��V�&�{���7"7ծb����ńK�b�C�`�\3:z������jo>�c�T�	�'~�Q"`��5"�O��g��~3<h�x:�؁/�b��0�в�Bϩ,�n��<խ��1�Я�)v����{�?���N���ޭ��w�T�$�B
�����ʃ=�X5���!OC���ܫ��Qއ݋|���������>3�'�UI3/���b�(�S��9}R�U�:�Mwd�{{��q�w��Bb���'g����K�
tL�3Q5LP�t��]?JT^�ZX�XH��u�`����=\,}�%M��x�ª���0��3p�N�ϸ�+�]2W�4��g^2�+��3=�-7�`���pw&��C2��<hݝ����ԟ=c�)�����]
�^����5��o���=�劼�O�ܵ�Nn�T�B��۫t�Ǣ�`�Z�OhF���u1��5j=�9��wR]�v�1�������￟P��}���O�eo���~�~t�}����+�P���Eg+?(�����4���z5� f�i>�k-O��^z�g��P����]�S�;�כa߻�:0ySbF�bc~�#j�¶��z�kxZ� �����Cb\���B��	N}�]Ӱ_Xm_Vz3�4Þ��Øl�/c��u�t���:<�\��8���=s�/�m�a��*�؏�3���S346��s�S�\���qu�#�2"'����+Û��C�P203���r�����M�R�����R��qc5�B��tu��<(�S?�ڃ�Cr�i�`&�kט���]{��lSύ�>�a
�eZ"���<Ȋ͵Ԗw,�͉�bwDX��b������h8OL�}�SO�X焕��Mlw�w�F�|<V�:�#���Qb�,���ʅ��O&�����a�~�	�c�����zg�lE�כOw�)��{r�TOM�"v+�$>�(A3���V��[�b��75m�6:��p���[J���ȟn��Z�T3}3��O�؁.}b�(*p�2�,�[��]#~"cA�=o�N�M���%C��ѕ�t@n9���!g}��4-R�j|�N��2l���/}e �6~&2eu��ս$��S�v�J�u���47Ԃ��W��k*��`
̙P��ëj`�ʠkoc�!Is����\�r��}����>�}G�|�ה�l��*��@�Ԏ�I�h�ttg�l�ZhP�*�8F��r�q�Ǟ:۟.��w��A��Q�R���)��-�R1�c�Ϫ�*��)�][�g���M�o;}hp~��/�a���1�M�[�zt���aYpc��qN��j�ѕ8ߜw�ss�=b����v��$%�V��/��U��)n ߗ�@³��1�\���Wu�V��K�v�=���P1=,d��%��_���T;�o�W�/�ڡ%}�o�����*���G���.����k��C״��V��j�jH��B؝R'v��/+};u38u6&�Wh�=vl0��ek�.��/��!�,�6z�ǁF��`�Q�ѩC��J���JL��K�9��m�m��uD�a�vN��������Cx���7�6�*V}Ց4�8�_�҇ۘ��i�͉)�'��N-L0<mCZ/���b�{J��淃�:�m{��e�C`�|���7����=wj��Y��-�9A���;1�p���/S��i����K EsHy~�יm!����iF���m!(���Y&nck��Z;��YY/֕>w�����r�SS�A:F
�2���B�5%Y��.��l�s��U��Aܾ��c��*�,5z3D;��[��^��n�]	�n�C5�f�[^.0#�F�We���#Ţ;����t ����^�̅䛲�K!v�us����%��j̲��m�
b��r*lCmWo:��6.�u��M��7��ɘ�m�Zi̙�V��V�:�JgR؍muې��'���֞=@����V�w�P-��X ����%���ʬHg.��*���$Yx���!J�_mY:h�(��k�/���old�\�Z&�X��C����ǝ�		 y�|e��ua��m*�n�:A�a�y�/�`�:l'�b.s� n�'/�w����	��OtEM�P����ڗ�d$��%_���n*���ڱT���wSe�VϱX��,��YwwX�Z�Մ�ww�@�#*iwy����,ˋo�m�E˼=Y�]�=F�liȎx�#�Ty72��kXհ���Zs^)�f�T ��>y�.����t��Ĵ��xA"�)Rqe� _=u,3I�5�Ռ��E;r��{8бϦ�
UEv:]7�v
2�iB�7�����u��u��/y�c ���#7x�28X���o	-�B欖�S����JLH#ЧP�т��XB��T��Ub�U�H�ÊUu^&s�TыK��x����@M�ޝ�W��>.W
N��v!��(1H'y�{~Y+v����a��9���rY�w3w���հA(���_H-�AU���}.������X]��(���LuD/3�c�C��C:���W��'u�w��6�5l��W%8r�G[��t���oM�u�d��j��pį���/�t���r��j�fQ-�6�dUy#.U_9�}�e��f��!Љ-�×����������,鷙	��>���R�Ʋ��#����>�D� �yqծ����W��W8�l����v�A�fz���[��6�0�y��*ɼ�fK;Ge	D<yr��H�umdܼ��K4��K$���ʧNw�f#a�Ie����^�㙼b6I�*��RdrN� �-��),�-�O�,ü�Z~���,�"�x(V�P�!���/Ꮽ��Ū�}4l��eM�K��j�t#��fc��j��r���Cx��3W9,�����7�xN��T�ǝk���ӀF���QhVdҊ 7کJ���2���w8���5�:w�R�y��;��,��ѣ�ruv4���:�Z���먮�殒Ύ�oݧjE��W_`*|��������pצl�G�Cy�*;�����:�f�46�A���q&ٲ2.K�E��5N���h�a���Kn�z
C�v�u�5�*!/>]�{�)v/Z�u�Tr?��K ���׷���#�̙[Vi����b��zhe�iMm���B�4�0���
������ӧ��ǧ����0�(��5�g],�1��(�ey�i�k� �"M�v�w�|����HFZI"�)�DfW�I��J��b.BF�J�Q��儉AZ����N����y=�z������V^e) �I���jy"bX��(���G��������g� ����iZ'�����ՈY��}OeW�*��I
����yrĴ�<5rj��))"{�{8\��d1��3�BԺÜ�DP�3)JE
�DDMJK٦�Ԫ���G�P�N�DP�-3*B5���-�ce��I���I��X��a��E�B�a��Ct�ѱ�I����e��7I}q5~��X׽����s��Oi�o-�p�k�]c/�@i�������+����
}����k.�WWI_5ck�;x���9l���!���R�������s��s���<c<�|�8��l��X��7R��`����E,+>F��eM\5/�k!�9==�#$�L�L���O ?��t��t磣����X�p�r�.�-�Վf��c��<퓽6<c�M>���j72_zu�����A*�}��>��BD�S�=(�pM�p�w���YY|*���<�E�R3#���ϵV�1�:P��mT���\�]"{`WƠK���+��	���11-Q��>>�Q��+>v��Q�k�n��+��Wn�2_�i�S�&��+�(�K�PW���%�n��@�@�S�-^C;gl=���0m��)N\�ts��o���*��o|�ߤt/UE��Apu����&��fo�Rb�z�;��5��'��tr}����@��vav�fb Xjq�y�i� zu�s�բ&���� �M��Q�)��K���":ƛjN�
��'�_�M)��7Yw���\��>�/��9��(Ӣ����%@��	�b�ީ�}^�o�%������ou�2�j[4��N(1m���ڳ�Ԣ=>~�hK}_�~?��x2%��2R���K}_��8_Q|�����߶�ur����f���w�κ�0�̀!W�6[��;��˕*�wBջ7��IZMuY*��.�Iko0F:�l��lnN�3k]���f)(�S�Vi*��١�Z�5�Aّ�z�����rI�� |?�W�|#�����3�q�MvK�������1��q�֠,�?`c>j�H���>3{5�h�	��}�c2g2��c�kP��K'����}9�z�ь���u�5ߠ(~��tj����?���o����;S%�'���1�/����������g��-Ǵ�b`���5��`�*1�w��=�{�ǧ/�S�>�`�����sa�8���j �C*��^�0��ӊ�D�ܳz��G�Ŋ6d��x�ĩ���5��_9�1. �,!cM�/7�q=3�s7�{jm>4�*ˣ'eLєٱ��5����X�A��|}4DlJu�tD6��*8�X�o�J����`'����c�cs઱�`дC�0g�W�����z��[�W��ы:�S����a�x;���Xw��:<��Z�879�u�K�	O@���V���E-Q��~���#/�t�HJ�]�g��upvM�\��a�кڛ�C�T���>��J��2�������{�)���3.&�����tT��2�,���RY���mɍ�Zٿ��<�Ӯ:��sHŠ)�D՘����~�.����gO�߲��&�։6�R�i���/���ne���;*���Rru)Z�=����+��cc��u����K��Z"{�00����ӂ�|�1�U����2��8�%�O���>��G����>���f'm�z���z� �����+��K`RT�1�ԛ�3�=!`���� �-F`��~��f�/	p�+���,�����a�
{D�gL�D�bi
p��OG�ྩsێg�4�Ń6-Փ����(겤 �\�N,>��`rG�� �D�11<$���:Q"�=x+.�����c����,_Xp���&|�l-�'����Bݧ�\?u���P�DM��)��zh<~׻��D��!�<6�.����Y�G�K�����"�+ϒ����#>m�E���sG;���E���i������T�;Ziz�]J����������:lHϗ��p���E�U���h���{�tB�Ob_���y���3`ɚxKs��/;{��g�a�A�G�t�J�/gFs�"�q���t.s�8���3�[R��Ñ���#��7Vf3�w�ᥒS�3O��z���#��b]1�ߒ�r�Ջn���]���[~�~�������nx�E�R�����^���"j��0ƛ�b߭A��N�
�ܽM`נ<���]W�ձO�G�{��u�e�c�M��ѵ��x\V^��:h�_+�ƭ���z�h]�9I��l�7]�ѠM�^҉�� *�,�V�P%�:_T����q]{x���v
��Z&^�솚Y�Wm(''��«��3{�UIuы�D(<�W��VU�8.ĭ���Xcʽ�ܦ����dP}�޻�{�}���=���za�g�7�XҮb�ǎ��p���+�F�N�Uò��Gf���bN�zjO�EK
N�S�T.|5<�>�ns�w�Կ)�b}f8�:U2��5 �>�(1^�2�@3bD�PbC�B	�s|�R�`Šyc������}�]�.f��`_������ܖvm����k��g�d�DJ<SϨ�	�x����՞����3.�g�7g�V�ﭞ���⁀k6a]���pOA��=x!=��=$)p��+(L�A�tܡ�\&<N[��} �i�S�g!�t����)H��W�ͱ���;�ݧ���P�	�=���>=j�������3��Ypc45N|�DJ*3�U����U��&����4e	���
���t}~���Q�/b����1�\���Wu6�o
�ῼ�D��������p�����-x೟����~��T J�	��a!9���a�z諗܇��>�1�;z�;�r9�W�P�Dx)a��4��/߄���.n��%U6���o}�F������[�#���6^�`ސ����3�a�y��������a{��3�T'�s��{e��'����8���˭0�/W���r����%F^y�͎[�48��v���W̜���]1J��M[���>-�C�<k���n�~�O���y�Z��{�9˹���Q���s��Xa�GmvK���?>.��>�5(~�)�ϳ�������N��>���������aJ��],C_�`�ݮ�'�����(���}��g����yU�v����PjE�9�AU�Pz`���]�5��m�`�F�L�2��Sl(��.�c�2����Q�ʇ�-	�����|��Ib�-�M[��(c׽�U����s��ͻ�>�~�`6����@H�P���
s�E��JQSW�/��I���~0e��d��>X�A�2<'v�OGG�*���T�38r���y�V9�8V����;�Gƺw_U�q�"��פ�l�[�M\,/vT<
�J���R'"�u�"�9a}��v��y��R�!�z�ȶ�����Z�ƧJmT��"�M�'���@�}�b�]曯t�����c�r���Q�K�n��\���W��/�0�)�@�	�L������j6�!�8ف��}"K��}y�Y�Cw�_,f|�����Ǉ���ڥq����,q"�����Y�@ְx2B�{���=�m���~-$�w7���{�ee�v�V���un�xg���I��f��u	.��o�<O�}r�I�hTe���"���cny�b�4@�-���ySn�����uuߜ�]w�������Um]�9����� G��7����1��}3�����j��a����U�~��8e���x�Fϙ�')�̦����vZ"a)�
��jo��t_T�=�";3=�eF�_��}1���\UvH_{D��A{U�Z�Y
	�Fjg��p�)V�T辯t�ڇD��ή[��O���'���Ʃ�9�qA�h�E�����YRpUı**1�R�LwG����!����=��b��Ζlt��}J)����EST���́G:c�&{=���U����&	�!�S���J��[��F|�y˩�k�w�
17�������q؍�R�xo�|0w�3��zi1��F��H�W��>�Wև��@oo�>�,[�LC�5��2�Teq��x;z'~�����w�<��;���(��H���W�͆����a	�y�i�!�{���o�Ӻȑ���p�71��#W	�X�wꣳ��;��vf���z�Z��`���>�KO����+�7Oأ�=�J�Zم4��,*�r��ld<	�q��v�d���ᯧ�
�6.���|��b��a^�����
<+mp7�gN�'d�T+&"��/t�ܢD3��/')�a�<��5�����Z���MAҞ��[�C����%�$��:��Z{����v��Q�;zt�{�
���}�E ǫ<M�بm���b�I�>��}��|}��i۵k�:��(�����k�2,8�S6�0�d�?=�%o���_���/� �u��d{^{ݞ�9�(/���bxߣ�������7%�9���Js��Y��UB�9Rʽ�;~G4>�e����p��+�m�U�0���u��3���}B�jo]�R~N���#�;����6'!ʨ#�d���^V[�B����P20� �2�e����z7�7=r`�D:f7��k��������c:��]�-w��<wB��C>���f���0�-����ea�����^��=������Ӡo���b��?X8*`ݘ"8A�ϵp�b��U���T�+�Y�aNJg�
Xcr�^@z�����q�)�2LM�k�9�G�3�����S0�]=N�Ak�8$ϗ���� U�(���2-p�S���Z{�6����E�G��-c�,`���Ŋ�f^�f��iQ7�{ڲ 
�V�����cJ��>�9�m9��ַT� �o�s��`Pz��r��_~��DC/��Y������<�#��pq����f��2I��
5k����,
����xgkr�FF{һ�(�(:,\�**�`�8���w&�51��nX��S�<�y�؏Z�����_����Ǳ�ܪ�9N�*I�G7.�E�ۢ�l�6�Yۤ=�S_1����
J�ٺq�3���;�]k����e	�P�����>|��mgg���b���T�s�U���6���xSs�=Ӑ^v����G*1����z<��.�2�?���	3{ʎϣ�9R�6�D��4�{�uf`����F_����$lD���[INJ�!�J�r�ϖ{�y�}#a��B�ʟ�蚱J>�w��!3ҫg�۽=w��q�>��E�S�`L}Np�8nuU[�����'#w����b�ONU��kdE��A��}��:�D�G]��B,iW1`�x��M	�3c�U����]kQ�/���I���1ɨ��0��6�'>9o�aΎt.7>��bϲۜ.��\d:��O�*�I�"sq��������}2bL܉ؤ$>�� ����)^ص����*�
?i��x�;u�w|�M�gm9�N�,��ʁ9����N��
�v}\e�N�2�;A�sr��=��yrKG�zF0��Y�
�ߠ5;�z0�� E���'��f�����������5\c�Xp�>x5�} �i�Jt��S��>�])�2�*��~�Y0��ß�k"[�G6EԜ%���P�:S�r�<�DX����3�۝
mM�g(s�]�gms�$�g�qð'9��.�gNk[��&s�)̷�6��U$��8����eRu0ʢ[��й}Վ�+��U\�S�e���k�U���#�� OY`Q���|߼u��|��־��u��BS���0x���o��zw�b����1�hj�"�z�n�}���Pg��6��3CèM1J}5]�v�s��M�/Z��U��*��{s,Y��8��i�#gvE���`�f�nf�T.�
�s�]��h����M.ZMw�p���UIy��0pK�A(�G�
�xj�j�?x*`1Z�X�zۚ��NE�b���b��׷�>��q-_S�D�?K[�"o�{]���Լ5�5�Jh��n�*� F8ݘ�d��w�B:����(��~ˏF ʰ�uu1����ƶ��*V���s�Ǫ[]��޻�2HuEы�����3}	�22�c�1n=�a��o9�l��7�'��5j5�)u�7�����1��1��ƹ��]�g�E�|��Ib�-SV�J���0Ȯ��w�����=�_�/�\�GD-�tqD���9��߁WDx9��A�JϬ#vܽ�U�Ƹ4����j{��]q��$J�f;��d<	�p3�5�F	ݺs���
�=2�3&��`T�A�p���*)�3kh���-���:kNg���P���R�6S�l5]&�vn����Y�6
��蜛�2a�ٳ�o6�N.�s��*�HIM��3)��w[�m��l���%T�/�9�y�9B���ޮ�6�&�����6�oN�g���G���>��>y��d*�^��qM���%�Կ5���ʃ�*9*"t�ȦDz/�p)��tɥ�+/<��ֈ�Q�\&<}���db�r~�Z�Ƅ�B�mT�p*D��O\
����i����.��gya�F��n8� �㔮���]�w�+��Dʽ�/�0� �dM����3��򺩹����$<�6�:���]/ ���{��Q����@,���2Þ.��������s�6l?�Au�q�޺������8~���Yy���eޟ}�7��;p�:9>��ERӺED�vN�nw����Y���qh��*X7����ex����1�N�e�\Q1"c�*;n@���L��МQ@������('EL+���bT
'�E��z��5�7�#rK��h�f�i����{�X!_����>�bq8�ņ�A׎՟����&�>	�o��H.:n�nOyy�1�u&�-��ux�/��"+�@X��R'�޽s�����-o�ވ���s�d��Kȗ�������J߯/�3ު�����.�!��~��^�2 ��n\Z�{+�6hl���Q��P:^�{ԆRc��չ�_+LoM@�t#�:�m����p}{@�B��'AXMڭUm��۳W!���h��l�*�V]!��r�a�x���8��a��O��{u�bJA<U3`d��,�M��.DP^M�:��4V v`��\��ϋ�
@�C�Q���õj�tcT36Uwu_u�_39�Ň&i#	]��u�Ӣ��˅Rl|q�|n�6AʀBV�S|4�3���N�B�+�ꓹq��u!lc��<���7�Q���"��^n<��g[<r�_lޕ`.F����\m,�7�n��t�#��}*TH��Ж��t;B��35#Ĥ���`l��2��66�e��u�����ꕛ��Nq	�fm^�30�%�Z]�}qbؔA�vh<���S����,'xg7ga�[�Y����UԠӮ>be�4d���g%o|�!P�����5�p���5�U�{2������.08�f5A¶��ću˕Û�vķ2�s�S,q�BM"��A���T��Ƕ��{j��U��L"*�}�<���ȁ˩Q����`�_J��dPÙg�"z��0^��c
#�Y�/�->�l.��/�hF���K����;v�!j�����\��G$�Q��+����c��@���s@y�V�][�O�p�U���p��)u�[�w�1Ś���J]r����tX�z%
D��.\�S�B�����KJ:mqW���.P��y��f�u�<�B�V8�fR�s���ma�ԔGz3+�O����$��Vʮ&��X\��V�2���qsި,v�\��u3w��݌�b�M���$�����I�p�Z�"��"�r�cn��V&����C�S�`X5���{
V����{��K���d��F���Z�p�R(�dꤎ� p��:�#-0�m1�7C�fζ<��F������G&la��\V�q>K��^u���5�(�ȅ��!�i=�;opU펱K�$V��t#A��:�5OZ�S\h;w7�<8�=T�I^��%	j�o�)��L"W��Y`6!yג�ə�q�{a��R�(�'o3�p�^�����t��LD:�/��#y�d���X5��t`�nwR�j
\�Or�����}�����]�w;)7-������7Y˪�s�#�L��I�ΐ]$`�K+�zX&�L������V�S�"�h�U�0=�>�p��T�+����X��]*����椼b
����q�UҴ��yq���sk���89U���ř7��/_r+�^���"�*�F�Z)��Lo��uВ��,�P��M��gƷh�î�N�5��=}�n9a���ۻ�`��tZ/9饨��ǎ�ZL�0�x^�Y�+�4����q��KY9��*�y��MӦ$i�R"�|������(雳�y��fI�}�W�,��y�P��|�WQI������9�*l�,�"2h�!Dx��~hhٍ.µA�l&L���ֳ3�3�u�̭f�zt����Չ�kZ���֊̈���{fa�>M���BԈ�,��y�{!
�.�|oc�("�,�[Ȉ)���bk��Q���r�����vP�%q�)$��\�'�9��$�垓9��1H��ƶ��J�P���%ʚ!��L��-��DDrB��5�Q�NdM\B��r�z]\��
���f+Rf�)��'T"�yW0��\�j�A(���\���٨g����^�<�u�|ϨQ(�_R<��凥M���Er�5�ey��^�̋µ �r��s&Ѽܹ<��3��(������B&v�^�L��ԞԨ�*�H��[B�ܽ��e�(�����T�#C��ͮ�3�£�r)C ��7#$��r�QDBoDf���)!1WM�c�ʎ�D�E���)@�]��2�_[�8s���T�*�
8
��U�]՘E���T����A��� ��>�  �{Ǒlc��%��6i᱓4<$lP�%͏_��"����.,[�iV�8�s{u]��f�0��V��K�,W�����9�Npl�f�a���
��.l6'>>�g¼�A���EZv��n��欲�?>���[W��<X��]g�6��US�*�_��)?H�oVNNh�}�(�!�G�є���r��klh��b=9R�k�Dlmx8�~�ު��>��ƎT#}t���
��̋��U�S��lb��`��yN	�}=���|u�7ں<����_C���w�bܯ���_���9�u�K�sa)�9��h�r�u�:U����zz��������@v *1u(SP����/n����k�Ъ`{sMǦ�d�N�s~��{5���d̃`����L:A�I���%�f_,�w�}�na�@���W~�^Vw�0�f�����yw��}��В��c��70g�<�Qt�Ea�w[���uX\���*�~� �gh�)�x�����G?�
h�#�P�<;����I� ����<��>��Q\�"uզM.U�r�N�꾵�����X?�Ϯr�G\�(#����������.��]lz��/ܗp�v��.�a�4Irp����\�r�Յ�k�k5�n��Zѹ�6�օ2:	:�o����8������?L3(�ϟ=�+|�9�.����^oEO�W��D3y��n�F}���p��򚉱��D򸍮�h�w�=��	Dƌ���]?J��o�pI����xU��
��UwƨgȊ��4+n�J�y�Sw��X�^.���sb�k���m8���9z,ߣ�W�&��{VDVr��0'~�"��>��V>��<�w�m:�6}��d��p86g��^������+�>����M������q~ݔ�(]�#a�~�#>)_�p{�a�lK�3�hT=�-Ͼ�����7m����ʍ
v���f ���(t��/ᮅ�ϓ9�
�ϣ��Y�
�Q���c���!9�%��=J������L0<mC��FrM1�Tۖ�lZWf�}�����r���>Z�O�|�S̼�5ݫOQ�N�8T���z�>�;�4�S4吚��~y��ݮ��~�w�
��H�9[hc�{��+__G��F�R��c����i��"ƕsN<p��p����)�Ų�[��zg�t����^���M@�<�躔�����T.�s��[s��,ļ���O������ݒ�nۉ��Nq�ݻ���
�Z�\�8�΁'E9�Ѣ$�FpjZ*�!��d&60�M�bns�����7v�e�z�f����:�rV�s�$8�rn;�o*3���v;�L��f�#8���^ds�����g����p��51&Fc��O�4_�F,v׆p	�f��;@}:*P�g��+G�=���{�W��x�eE+�S0=��M��f�N�&��53s�Uz|$NGX�.�T/iLǅ�foٕ���)�Q��)�{��t�Г�>�l»w��=���=��P�Z4So�;�?�X2�x��oz�0C��P�prՇ����D�} �m��N����IH�fv a�
|&R����s��v��@�,O��$A�󾹅�b�c<����f�ӥT��
˃�+�»�)�,�ʦ�=,oK��vl\�	��퓿_�a�zM���(
�S[���ӌ��W[�k�
��k�&e�#��:���ɟ~�*n��x�E�8*-�����NpA���U�u��MOe�2D����BX�A���7Qk�l35�P�DF�"�b�H��޶��<�q��£]��	���f�Ӊ�#9�I����a�7�cK>���pjr���dO��w;E��|��{��� C��>����z3�_��ь��t�?{-�2'8ߠmMԬ�a�\fǯc�g��3�}��|Э"H�B'J�`���e8Jպ6ݼ�*��Q��љ����,��MlM
̫��W}|o��HVY�Q�T�}[p6N�4�\s��9�ԟv���l�D[����]	Dvf�V��������1���^y��
̀�鿞����lߞ�Ϯ�(qc��E�]s�Cj�.5R7�q��8�J�ʁLK>��ȷ�e_��5��ws�q �;��e�=9�Qy;�VÁLO�Hl��>tc��-�Ц��^���9	.�v��A�wa�������ã�'���߁[�Ǉ�t��g�N������_�X�>�.���>Q5Jpk!�Mc_H�U�D{*��=a�G�U(ɹBv��!�m�j��1���3az�K�]�R��k!�|r��ʖJ���BD�S�=͘&J�z���4���e�{-��23���\���B�mT����4����gW;�	��y�� ���r=)
Ps���/B����I��tL��z$;�X�hٯ��T���w�P���|(�w��"WI�}y�Y�@���0m����S�) �\�څڳXf=��1���	~�؁�B�
*lT�K���S���f��{�� d�M��*VEv>�,7_��0�*!r�0�*B�48SS1]>Sﯪ\��2K�\=�G�P"��yU�(>~��e��9?af+�pc^K��KFi�|h�-v#�gp��`f��mLRV���uw};}���5<�x
���3�b��@�%�Lۓ(��F�'VU�xv�
�`q���&9�ή=t��:_�j�������ǳL�>�v�}���}@|7=�&?�����"�~�nh�_Z���}��>����t��L��
[G<k+�b�`�Y�7�|�Gv��b����B������M�ςqA���yO���ʓ��q'���R��\_� �����*v��[���r�� gv,������'�`j�H�޽r�:T�m�zW���& �����`���������Y����+r�ь�����x5ߠ(�1��n���k�t����%�9�Nl�ϕ����$lh��@����7�y�߯�>��8�߮|d�q��������|#ѫ�̛Ϻ��͜�ɣ,�LԸ�{�\����bs�z��Jj����G�1��9t�Hϒ���~m^C��c�ߪ�ϗӪr�� ��ki^yGW�S8�� 7wڱ��%�UQyoE��rjܷ*f�����5�66�ٌ�VԼ����z�e����u��G���q	]1�\�w��s"���*�r���ş��Ph��v{���"N�Ӛ^��sWӯ�`x1?g�����ȃ�xߣ��N�,l��%�9-6� Hf 8QȎ��0[?�,`N<�v'�;DW~����S�t^c���m%v]�#&'�NW����@b��(e�x��~�4��L>1�=�6��J��껔x؄���׷�T�˷��>FLp����C�F�Eh�3����ax`�|������w�e��D3���>{������W��I���F.��0�����xct.���^���>
��Z��Y�u��ʖSs�>�ML�^��A��n�=�]C�F�Y��,d,��7��F�B�����͕�j��^~��<x]g�?Yw??�~���U��B��Q��!R��c���ЅxZ�{��{���H�;�c��բ]�>�]ӥ�;mT�<v���";��6��>���p��Sd��O�4���W_���Ό��ũ�W���^G����Xg<�c�=.0: H^�'3a�|f	�!}��&(h��6|��aW�x9�G���3a�s�g�v��c��C��޵��8�L��6���t�FϿ�d�O���g�w����{Ɗ3jfV����8�ӂr�X��¿�]u:�T9��hx4��!�[����_������������oG�~��|UU�_Hd�
�P���5� �Y��aQ�}XN��XX�ߎ���٩�3~N�������=��-Vz
��
�b1Hp��ؕ��Ͻ��+6�D��|�x�#{����W�߳uY����5fo�7.�,S�[j��W`,�:�˃������r�\~m�~�i���Y�fJD�:}z�Nݾۼ}�
Ȇ���W�u�Gnp�eI2�`�F����y$\��:�Z�=i�@�ë��YB4�]%Ҽ���46q'�u'���������b5�۵�_�Da��`>R3��ujc_A��F`��{�Uc�����^b�������ږ;�<�[�/d�7�1�pn�����,xR��&��O�\�0��Ԡ"�J���-5c�*F	����۬�ݣ/�~W���S�]lS�~����)}Pċt�<�M�!�\łq�ঃ��c�OJ[.��c(��d��c�,>K�7�b=�P8l��EԠ䛠��ʅ��O&&I�C2��w/��WҸ�?����>
h(�j,v׆rdę��N�$>���5�k\����7g���*���Qʕpy�#֠[��ٛ�V�Sz��X�e@��꺘��=0#��\Q��3Xp-i��Lq�(t^N�ڒ�{�T�#v`=f�+я:��р�Ț�(Ri���%�^���{�Ʒ�v�V(*pr̓��p��A��W��%;-�R03��<g6dĺ��z���N
�@���P,_�Px�߬�����G��ɼa��N�UL_�}�c,��۽Q��k�Q�#s����Z�s$)�\	�퓷�n^�q�֢>��7K��d��ԍ�5��zԥ}��X-�F�	�5eSݑdp)�v��?.6�n��=oQʵ�e�������ݑ��Q�b�(��a��US��u��L���h��{�7@��v�9K�2�B��c���wJSz_r�;���s�l�3~u�����}�Y�7��u�m[���r� 3sӅ]�X\+a���ɛ*+�f)ϠOel4����1�}���\b<��U/	��		ϓ��[F�-p����f�`�
E[�G�C�u�sj�_�(��y��+\�>��u�LMF�a�{A�ig�ck�.0�mK3q>[=n�����vQ�C�xN��V������\z	t���b ����FD�o��P��O&Z��T���)����E(�XN/�]3��7��~܃�-�hN��sSҼ��!���t�#|�� {׾�y��a�PBl��W�a���������l�>_>tc��-¨�O��bU�P�	o�	Chd��f�[6�8���w�Y��e���D��~me��x�e����fG�s�5�W�����PԱ�p�6�GM����9���VDz�T|�3%�c��z7�\�����o9�P^[�B�׊d�mˀ]�2�M�o�T
��V�)�����?x�>��|�/~��Ut:�N�,]���̋+��i��*�ʄ��OB�R'�	ވE�ś���虰��1�Ǝj+��j��'}K-���g=Tj*5�޹c�C,�*\�-r�/����K�C�����-g�"!*oW��\[�73��N<����+�����`���zj��;��2H���9&�cҸ���N���ǌ�1��8����(M�?[%ǢX�����-]l��b	<W8/\�&V[��� ���Хge�C���~��4<hH��
����}&��9ѵ�o=f�M{&gފ(�Y�}��w����]��;r�ô@L*A��\Sb�:\X�T�zp�_��~��$�]{�(��g?9s�O����8Uٟ���V��V�D �O	j|*o��{њyUWB�U���k$��d:�Lv؈V�JN�
��'>*(`*��\+!F0���J��X�m�{�mow�!Y��;���%x%������8�Pb�9Qjxl�`uVT�l>SY]�^Vb�Y<�bLT>�X��.pY����8X��Ȋ>���1��U"Oj6]<y��O٩~������ߗ�3J�X*�R����z������9޻�c-�G.�!�3���}� ﶋP�;��`z��}��[� u��>T�9B��C�����#N9`:�}Y�s�s�f��Y�f�o�QG83ٴ!ƷV�7��5��g6iN|�]3vxM@~�͆�ʨ�U}��{�ne�*s�^%�LŃO`.[H_R��sm�ƈ6X=-�DPbƼ�۴k���QQIAևQG_�0E�;yG�X=��PA�2C�V���5U�koc��|4�op�;UIR��X�t��vX�H��5�5x���u�gN�w!�P�"P�AIb�� ��nHm^C��c�ߪ�ϣ��sy;3B¡�=!�V�$�n;��(�s��p?E�,[3�jܷ>UV�����xkll��1��ڗ.-��*�ϱ{�����2b6q>��<]s��ndq�m�
��D�`9�:���&��v���秩��z~�?�V����	q��dA�<oъ|�L���.��~��K4"2������DNn�W-yE����	?N�]ы(SP����/o��Lu�^V�i�����G��6:��:&qϦA�W3�D���W��$���%{�0�t&�Dk6&���W���W��^Y��	Zrc|խ��w� ��#�ճ1}P"~BL
ISϳ&�f��:O_Y��y,{*�|�k�N0���t�gh�Xb��?{ウ�P"{7��*�gW{k��A!���aԸ󜾩3���Q��܄���qa�sj89#��Ѹj�N�����_%��'�W�n�ѭ������#���Lߗ��U�®aA @z4כ��_��c����)���?`�%;����GI3���ϻ3(�+*�6�[�E�Q�g��D�Rp�9h�Ѹ��76vv_=��8��8Pt�˼v�E
��F�XT��ii]/b�;��ZC�`ٰl�x�5�r�^IG+"v�Y�i�l�\����k�LP=����3)Ebh_iV�P���`�7�e�6Jh�]���ҹ#,�C�^ǃ7:�\tQ�euF!c7v����C���-���gX��q]\1,@���K�2P�w�M��܊*����2���9jn��Ea[���h9f�Z:[d@Tyb��hubZ6�S�Wb����ؔqʈd:�\��v�%���Z���i�<ƫ�(a�]f���y'�/��Y9p�w-	v�1ϕ8��[G`=nï����KO+\��з����=��]�"�2w-ǂ�,�Q�;d�ά�;����q����p6:�SMS�E�:��׽���gՒ� Y����;H��}S�õ����O�a���E��Z��f�6uk��܁0*�GY�e
ע������.��H+R��B���Q��l*yO����ۅ��x�.�8����+S_V�399gn^����������0z���)Mmd��:�[&�<Ǚ��y��i�X�{����vk*Gׇ��|�x�o�Kޮ���N_�b3��cv�b`�g5+]k9\�i�B�lzjLx�U�
�W�X�9���M��(�w�LL$�s���a���	ו�rXkf�O@��[��.-mZ�n,�y����nr/"�ҳ�xY���!���v�.�g�n41��j�n�6�N�MSӎ�V[���D�郘y6��f���lYJ��*i4Y]�	*��+z�<�X�3�d����My
��xq!֨v\w�m�}s1�KU��Ѳ�oo���!���'��,T�7Y��A��9+��w���Ɏ�-��z��,n�t�Ǩ�|��☛��&e0xJ�����wu�����K�<.�@�:�[>Ɇ�l)�St١�ޣ���>˸�tΗx��ɂ��ܿ�(�����`L[���CY$�ׁ;-d2���_kC"]:�q@����1�RY]C��F�L���MZm�q/f����]��{iam�1c�Up����e�7���3�Yw؎�I��tn��
�Cb��1%����K쀮�5B��ܠ~yr�cت�iveX�u��;�dՊ����g#�0I4�\�ݭ�BT�����	�Ƨk��@��L�JyD��
V�U�nPD��C]�6��2���r�ijȰes}��S{s"Go��]5u�ME���qf��q,�J�1|���x�X{�����7&×2�M��Uܖ������Y[�(N�[��lԅ��Yj��e����[�*���3�鰚���ԝq�.u����{T/����A��n�gs�7�9(���ԍٳtM]�����1<�U=�4�V��5��;P��p�"��z˞QE��A�t����zzy���.�Ǔ7f�e�#1�(y�o&EAW��yb**��DjJ�Y�̢)��OOOOA�WFX-]E�E�B�-5�vVV�hU]Sԍ<���?>�u=�Qfd�zb)a:Q_90��<15�(��=�۪bRnUK�W1,K�r�{nEEB��#�I\yɪHDA��عPMB��,��T��x^�YQ]"� ���J�+ڴ4�#�R�2h�i��bra6܉����^�mM#����!�UWV�;&лם������\0��>���sŢ�q0�
����"�x��#Fe�>vnfhNk�f�#2.�9�򨊌�R���<.�P��U����J_=f�Ny�hJA^yL���"�$�Ùs,m��V�^B�G�3֪$�G:�Y�`zHE0"�[�J�Cuʥ\�ØS�-	��j�T�n��ec�U��}}|�o\���va�MB��RN ]'�0P���1��3!�X��4sܻ+��J�%4�(ë��E[·�Օ���T����6�q.�!a�N�����<�ߜ+�v}��?��G@g8�׃	��H��\6�e]7/E��;e_{VDTܱ]����ݻ�ӹ��X�uy+��3�s�B��u�ѮLVM/u����]�^,���[�vYb22��sV��p�a��L���8-�،M_�pu�?HȐ��L�Шz���[��l���ou�G��aQ�g=�����֋��Fq��j�a�}���L������T��>���w��f�{w�^�D�碭H�u}1�s���fzM1�Tۖ�,�瘠dc�E�wb��sbni��sq^�}S�����Q��Ҹ�Ⱥnc�Sp>� ˆ�Un^����GL��N�1�;�<��%����"�h~�����1W�|<-EԶ$uJ���B/J�� �x��aK�3Qk'�p�=��G�E2�+�F�N	�l����SW��Prp���p�'��yZ���:��}�]C��gkgy�J_�@���f,vo�LQ��D�)��ԑ�q�}�Cr7U�8�Y�����5{�ϗ�����m���;P�5�P/�53@T�nD�ooWi�� �(�ِL��?Iӏ��;}[rc���~����xiy�j\5�e+y략�Qp�G�ckF�&遾�,,�c*У�s_�S՜3^˴W1i2�P�ۆ)�L�婫��yE�i��r�W�U����mh������\�������6`�NA�1ݿ��]�䶈W�U�Ӌ+�{c}*�Hԝ����y�-N���3�&+_��k��˟jP��!�����)��l<̓yX�e��3O�~N����IH��x��ˁ7[BhQ�w�C���?N��w� !?DXC�Ĉ�'���� �yHq`�f��������zz�W���n)����\t` ��8�DJT*g>!P���8��v�߅��ʆ��%q
~F$���DU(�b�Q.;/���.�3��>� ����r�46%M�����T.�
�s�
��4�]e������=�Ls�Z�d@��X��A)�E�7QaxV��_�2*�����E�_���-5�h��1Km���o�c{������4ÚO���ϣg�.<n��t��P*��ʽ�̍��G��@})`��Q��+�<S8m?eǡA�H]LC�����FD�u�N8�왲F�W�\i������T�5�5��F=?�}t/�S���7��.gƘ�?xC���$���9$)��fzX�m1ޖ/`�ߺ}�Q�'bb�U�aȴ
G��E�xVE�%SA2����q�X2U�11^�ö��:MP8OZ�r�U��SxQJR��]����5xn>)��&��e.j��I���E҃�����6�u�.�+��Y9]ڏ]��.p�����o":���B�t��f�$�KWf�MQoo��*���1�n8�]�h"����
1�}�Ľ-�5sP,�f3��K߂v�8ϝ��t
��:{�Npl�f��!�n��>!7��
ٻʃ��P�k�O}!�;M��Wi��SWKnN�P�`�Xdd��9����Qv}'�*�,�����x�`^K������Ŭ�V?}U��k�ByiK��y��>T�TD�s�V��v���.�C��j#�X����`]��yc��y��8��	҄�*��@d(313w%�=
vd�P���BO���@�)
�9�x�������'��>�Dʾ���Q���ub_���t��^�W/�44�;"h�"��X�k�%�����Y�i��}#���g��7\�/s�9���ntc���q;@���B��<p4���Vi��z^n=��fj=&��j��s�~���~*��IUF���V��V�!P�)����yװ���{��s=�V�ʗ/��Gv�JHS�!<TP>ϊ��p��HNk�/	ض���O߮�}��U���@cD�dX�w�v���ׂX!X�g�;��'�����O����T'Ѧ���l�,������D��A�9�qg(�uf\)@ރE�w�-t�,�V�jKb/����$Ϯ��Kj��`!&�}2
&�zvpM���}-y�,�
G��eO�j��z���Ur�gQ�+�	+ݒo�Tiq�v.�Gk�r�?��T��*��_�O~�j�h�qaS�;�5��D��#��"+�@X��?�މ��l��Z ���?2��OȊ�j���
kB�j
qq` ���}r���3ýw��m�G'�z*��VT.������Do�l$��<�?X��LYB��C���ŋ�F�΀��7p��=�'��Ub	?����hj؇��x�٭��sd��٥;���:�
�ڷ|����l��rm�BX*��j �C/�!��ͫ�z,q�Tv}�s`d��&T�3s�f�<������nb�P	�PC���5n[�Un[4.Mc��v�W��ӥ���L5{ዑ�=��8����#c)���D5�0V�GvrUV9O�lbv
C��zc���g7�A�W ����}=p+`Pa
��
q�tDu�Y�S��`��Nʚ,Dȁ{�t=��s�����j,f�x@��+�W@V :Qb��"���Ӟ��l4+�EǷ�S����ϝ�7�]��S�џ�8��<\�P5��PW�	&n��L��߭��_�u�)V�X	�I��Q�Z�S�|���X����g�`�����]�=�5>�N�I��o�L���&+v�7�m���5�=���pӗ�e�ΩmN)�̔��-�b�k;�~b*���^fl����ΙWY�H��8Q�>�u�����9�	U~ҍи�Ig�w��&7�Zٽ�<����l�G_TB
nY��n!��v��[����԰*c���*�|y`��~�]ӅH7�q�`�����
�'�
5E����Ԓ��M��)�EԨ��_T���X(��nB�!��~N,>ϛ�Q���WB�wll{�ə�	t6zޝ#�blJ&+�R��~�]C�ߺ�g�/)�'�<k6,���^%C�y�����}�"0w�}q���a7�ulm����Y�Gl�a�S;1YW�:�����Qٴ���!�Ug�\�٥��d�B؟@߄�l57{n=�����fq��9��'�_˙U�<�1#��q��[�&��9��6%͙ɚ��h�H;����ί0B�,t��W�_AH�͌i�=��s�k�p������ledV��tՋ��<4�t�-H,�<�C|*�#�"���W��},�}&����t���Zb�����;Ӧ2m�'�7xGzq�1쭩y��+��t�#pE�s�#�>�2M8nT�9t��v�}bw��'F�e"0�zolK�7��[pS�;XJ�>6�u�����h�~�֪�JPVZ��'^:q���Gx�[o1���ҭp���ȅ<T.�F,2s���y5e�h���7�5�-��F��T�kh�@��.� �����B��������]���&FO� 0<z��m�>�W���lH���y��n!�*�9P�7x.7���M�(]��ՙ�1��Pރ61�&V���>٨��(0�z/��9a:ux�8�hxf���ї��j�ca0yd�ҽ����fSS@���b�b��1$���bC電��}���^�T_i��V��r�"/e�V9Z��1o�8����j�jl�j5�PL�FT�OVeO�������� ��3�X�
�9Xe�Y��R����5�0�F<��pOD�~���_�Su{�ow���/dK"xA���Q`PT�e�8�˷��6�u:Jv35
^��(�S���c���B̆9x[�&_���$1�b�O���0� =��&�*G���]��BVe\Wg�kw1���&���:"U��\�|B�<%�ɪ�^��卿G���ӱ�1Un����jc�Ao�(��D����2�͠��Jǧܪ��{�(��B��5�Ӧ��ȌU�F3�J#���	�R�_��@��V�5ʂB[��?�7QaxV��W�P�DG��yw�ȵ���,�R�hKT/�Y��OJх��m�[�HQ���:��
�ژnᬙ$��՛~�{3����Vk1E���
r�qu�R&�dݷ�t����p��,)�����˂3Qx{�H띬T8��ѽk�{���t<y2�~{6➿tK�����{���^�6����wS3��ؚ�^������K>���K��u�����}�BO~����`���*��!^��}eǣvN��!���b����xر��Vf#���R����.��dk���Tz/��=t,�3]׮��)ǫ9�%:_��}�
�����81J��3��晆YA����W�_�?�%��We��*�6驉!���غ�j<b�p���BB�5�����ݨ1�x7~����Ozi�}�� X��6Kb}���n������W�W*�,`R�<(1z�}vܿ5pԿ}��8&���ݺs�� WRg���AG��rԿ~��	�W���v$#�}�3tڕ��2��^��0c*
Z_/m9�S�|;|LI�#&t?�:��b�t.]���̋!y��U�LhN�'�o�z�������@�Ԙc���Bz�
�����'��v^)z��F%�7~I�%\�
�2��w}o�TN�>3��78�CL❑4=7�a�0���̬���tmFC�vO���E��͡��D�l{y�C�Ñ��m��ti�N���V��F�f.)W�*�fΣjbӽK �o	����ܫ�U��r�P]����ђ��yy�0k����nmz'�~��)��/1v��r8�u���/�����6�.lU��9���}}��z��������]:�%;snLsܸ��k`I����z�Q_z�x�Di�E��)	玿n��w,r��;�Y�o ���_�
�1���*�
�T"R%{3H�W�q4����wC��S},΋U,�Q��cM�'aWք��*���E�d0�ea�k1�=y՜��$�<�2�N@���,Țu�k�}-��B�_�z甤$���h�G�#�k6 ���CQK���U�;����E��=J&6�5��^ �06��W�g�x�_Zb-��t��=?Q�����R&��L�٨��n&�Q��:�h��=>M|�:�K/!���T��O�^���������Bw�15��f��e���L�*]˫�%b���2`�u�Џ�*BP�p;U�X)q� �bf�x�C�~�����͚S��0�{b�}�e��gu]��6t��@�b��B_��W�(Ϥ�FWΆ��=x���;>���ֹ�%�ڵ�y�֝���"%���CT�V\���>�`>�g>�V��-�����b?~7��c�ׁnl�+v~X����Iμ���fϒ�U�nn��E(���<�H��{�|,�n��J F�By�
�;Y)uX�ׂ ���Wsc��,v)���-��Q�����y�Ժ=f�ȳc����n�4Bz���(�͝�u��I�}u��j� ����VÓ�m<�/M6��:��V�;�q���U{�E��{����oBP��i�Ioq�=��XcrP}$v��miq��㇕ʨ�F}�Rw̛l�o\��c�u�F���B0�-�K5u�}���q��Wry�������c|��M��*`a�z�~'�0�,�
o�zz8�꼪<i�J^���}���ϭ:��X�?@���~VA�>ؼ���Y���D<�t����y��I����
';@�F���]~;V�E��y���3�pE;��A����}zT���-��ާ�E8��յ5o������#o(��7��`�F�@�bG�T&���.o�5i���6�=�Iq����]��W}u��������V=Q,*��i���yG}���:b"�G��Qֶ6�[�W(�oR��/�������7���x������O�1�����`��EH�ὤ����!.<-k��ޤ����c���; ������,�!O�F�kWO�$���M�t�b�*t��u{� �	}-o5{]ݑ��7�b�#v�r�̏vܝ�R���&ܹ]�v�.�u�n�N����>�))K�TG^_:�y�]]�Ey�m�	���=y/��t��k*=>�cvsk<����<5W�^�3W�ϧ��|���;Xg�#�wQ���O�E��y]/�ǗR���8/h�"��^ky������k�~��WO��tދ�Y��|�w��͉����8v�������������y<73���e++3�>�|`w��]�8{f�ln�)��/��n�n^HwQ6v�<�UF�L!�׻~Ki���B{�ܕ|=,1�A�̟W��������_GX+�����n��),ߙ�����G}�~���˞����u�Oc�c�t5j�
��io1y��X�`	�h�]��aw��FW�Tw�e���I�M��@}e�ݗ�+܏�R>���^k%V}o����NDLM!:\'�=:)����k�k���x�[r߷���� �9���o����Vd��P[�۵������1p%h�����l�Ζ�4��҆��T�kL�b�o��I�P.�V��:nԟc�5ݚ]�bi}I�L`�5%5��z�\/��GPF䚯��^�9�o,������(;����;�D��U�Jn$ч��;�oe�0XG:e��[S7(����[i�Ӹ�EJ��ݧ�D�)E��O
*V:���͝�/S�.�u�*$y��c���"�}DzY6Ԡk/(�P���[������*�3��*u��.n���)�ְ84�w�ى�4��V[�yH��)�rf>�ْ�Ne���d�>V�ѣ�Fw)i�D�݀�L+���M�cQ���g�WJG6���\�fnN��ਨZ�ڛ�].Х��ٝ黸n�dħ�E��5/ua߯M���y���3�a_v�t��l�\��HPBH���}�V��E�S��,� ��%���c԰�Ri�l2�USWVf�����q��@�V
w�c�r��=*��$� I�*�^�4�S=��͡j��ϯ�k��9��r���}����HHu�����]�2����ms���*P�J*��*��P�SM��k
���^�[,n�v2y��v���3�OEz�Nu|D{ע������V�j�1F�u����XR��ٽ��k�Ԅ�ˊ�����w��\ڻ�y�5��}V���evH�IJ�\&��thJ7Zm�uZk�gm�)�i�h�g�����XBW���̄_H���c;\��Ӫ�ء]�5��u�n^���Xzppӛ�~��@ݘ{8�s�	������˱��X�A��#�6�[�d*��'ڭVʰBG��K�ծ����a.���4u����^�̮i�́�鰕�����tY1^��`��\��c:�3j[�8��V�z��I��r���z3�"�/x�D\��.��+L����Dh�}.�<-�ef!-㹍���Z�Q�}D�R�7�k�P"#/2Wr�����g4����9�Q�Xz0���f�rԈ�M�`��S�9�.�^��-�m��^Wnh��'^
�"���A�m��9��4@q�/�>�ˬ�VP]�s"�n��QbpD����iV�c\�K��7y�v�G/u�`>�L,2���b�LN���4E�8��+YB�]XiL�6J��v�;S����[U�vkS��'�͒w=�k77���s�`Hc��Ა\%��ђJ�R�>�H�;J
7XwxD[Wu�������Fgl�sP�I���V)�W�
]r�SƓ��Ս��M��vr�h�.�|%<���§�cu ���ǜ+�ד��t��c�$��7��c��u�镳1�DW<�Nu./)�{DWZy#��q}o);��/2�Ͱ�>��N7��e���q���<��$W����Ye�9W���&���Dp����(�V��EfA�DU	�I�h��!)�5h1��������S����dWD�<<5�K��c�7'��%�zV�\y��|��<-JkZ�e�U�e�S���������Y�%g�T�y4����D��٩�QV�T<�z�����ym����Y�
d��|5�D���됟P��ޱ�2��c��{�
�FJǷ�sG�g��8Ox��S��D ��!G��:6���ș�^���P���!2��2��H��G���.	9�$�_{eTW��B�Is�D\�
"�>��YY�z�Խ���g��=����Z�V��D�ǽ��1��n�>�I%EȲ9�yԢ��"EUSDKP�B�TEl8f'�3��th�TN]D3�s���v��+�D��(�:�;$*�;e��ѺTy$�̪��=T��
�T�,��'mg����^5��0ccp�EJ"M�.�1w
�(��J�vۄ�	�����ͧ�r�^w�� 2f�Qƻ��+�LL�X�	۬ם#�(��C4�C�U�8S���Q��1�De^mN4:P��65j�䪧d�������V��B?{��q�kՐ��H��FB[��~z�w(��giB9^�b���x��|A
/���ң/����:�w��{$�Y���V�U!�J����-�}P�^���\�Nyei�"/�������I��'ÒB�m�h��Ľ>Ud��l�AF��?���!�X���5yg���6'����B�.�����fԞ�^����u p��[Y+�0	�Мn�߅^������>��:����»�"2�����^�]���H���٧�;���J����3��Q��+���ݸ�W�WG8v%�<�r=v���}co%^lKh�C�[]�g@�'k�,�E!�5%p�hĵ�$[�i�	������6&�~6�����-�|r�P�@�!�
�N�6�Q-5j�(��p�nK�Q��3_��9g��£����� U���^�V-e"��3���̙��u���(�	�C޴��ح�.z���A��@��Fgk���'j�����;��K6$�,��f<�{8f�<��s�3h(�9�%��Y��̎�c5T�#�v��>��������%�m�//�޼�v�OAx��6��/_g��v^�wz���zz��ÏW�2~aP�_Yiv����_U���Ξ8M������T����HN��!��.�h]B����������z�y.�+��s*ew��.��Ԃ>*�Z�Z�A�*�T$>7]|�k^WzE=w���]��љ<��׉ى���}l�òǯ��&��I�U�Y�f��h�Ѿ�8m7��:P��d��]{�����VWXJ�"TeOIu�V����r|WA ��4�g�����w)� Tv���k�&���%�����=��y]G�<CΦ����}È�j��[bӆ��1����ٷ��2ua��t�-,r��æ5l�o(�i�B])��7P�z�.{W�������/m��Y*��t��q�KEY�g��Ћ����b�w;������2Qa�Y�o,�oWZ{yX2$�9�<�3�Lwv��7c�қ�2M4]�}8��RE]�GN�٬�h؜'X�^D������`�����Y��e����y)���v_G�q��G�Z�>��N6*'�:ۋ҅ݚ
+��m������@�$���[=��m侨�kCQ1��mYحݎ}�1�ݡ\Q��>,?�8լW�����y+6m�^����x��<�S}�,���c�~�,[­������$w���������5��{�gy�ovW��!�l��у�/�H�u6�JD.x�=J�M�g��˙��5ݷ{�?�nJ���Cr[u�����8�6ہ�:`UH9[w9܄�����k�s�>,�����D����7�mk�|-]����WE��o䱗��>f;�]n�`����Wq�:A���ٯ)��E���+�^�ϵ��#W��L��M���G��qP�^�l�zww7�l�X���U5�+8�-�-�k&�˴���_d����r{��D#>@X��C5!�;�JL�.~ϊ'9x�r7^�¥,L7���̙�pR���3�9�P��n^��m�5\�j�J�0*��av��5j����>��*��c�3]�D�`��@�ڛ�`����w�F{�:�����Nu�&���BjhL1��[��լ���ri��Yh&Ƈ�ȂO����Aİ�J�,����������~�1oo�M�d�Ƽ������^�������f8�h�4�eyu�\������c_�|���=�6�������2�-Y*��D���ᦾ�m�n���zO�d���x�����I�|��}`k�x��c�4)̛�FLM�r����c��F������������zŁ��G��k�s�>5F��`�����qOT;�zwm�����WV���?��N�Ϣ���Y{��=�Uw�1}��o�q?s�%�#^��y����*�z���-ɍvae�ǔ�@�'�ׇ�<ϙ�Z��y� PF��4Kc{`���dI۱y���g�{B�������S	�x���>�g�.���!�lgu�さ��\Dp�g�O�� �>QEYk~3����L��I�b7%_�<���^���c�pd��5����sF�;��6!"��b�%��KsX���"mr�G��j�SR��`�3�'�[�38�ᡉ������@ub�9m6�]��M�N4zt;���Ʌ$b3���2���b�!�TG�t��C#����}[��r�
��@ާk��w�s�V�f��gܺ�1�[�V�<C�&w�iQֻ�H$���r�vn�U�}����j�cT�'�},��f�+9W<�_A���Q�W�9P���4V}��^��G�K-�3J���}��rR٪�Kם�J#ג�Ӏ���w�1��>S��|yc�%�w�^b�����L�<x���q>�l[I��`�_�pP�����?\�C7���[&�a��ex���Q9�ƺ�-X�T��x5��\�:��U����W�f=����z9�p�ӥ��ZT��O��岬uD�m�9��&Í��t#Ǩ�uxnКZ�Wo�߉���M�9$-�ņ��y>//��Z=S���b�Q��O[�ê��Bw[Ϫ�p��f��kXVZ�����J*��iC9v�nӇ���5�l�CT47��꽳;9��|3�Jti�f*���Fx�;�� ��C���[Ý�\/��'<5�.�4([zL�|��ٵ{�5
|F�VKS�
'l�+vs8�R��D�]�����|�	�i�[c�S����� �e>��t\�8��Y�C��$rM�Ȅ�k���$�ne�BzVʝ ��s�ewwz7��Kq,=�+d�����lM���n��s���1ق7Ķ��g�gqvo��U�ؖ��և��mz�tʾ���۹+ډ4l��l_����Xm}�V��x�<�'�lw�]���t˹��+��Ƿ�<�u�%���`��Y6�Ц�{j�E<��лL����q���3�1'���3A��4M��z)�'�u�˶�mz3{�P�v6�=���b9�CM�Ϝ�����tp}����w�f�Sr��o�3������#���J��ܞ����T�j�.?I����Iw�E���J�r���G���uǻ�R���yy#V1wϭwXZ���c�?��P`�5T����_L�S���tۮ���{�䥯e�&�V[�,{��`�A(�;�gQ�{��.7�A��y;V�w�,�9�s�.���+�/}�W� ͷat�����Q�#�"�K�ᣙؒ�Y�t�酩Ul�Ƽ���RZ�Z��CҶR�z��5��XrJ��=xn��ٞ�D<�m![K��7/Z��\�[Ѥ�rIp�&�Y��G�NJ�x���Y\��y0�#���L��U����1�7aUP�e��Y�A�����4�`�C�yGag��!��Th\U�p��Og}7�&H�h_��g���T&����7�q�@o�;�[c,D�J��#I۝�z3�Ȱ�����c�%�cTƭ��9�\#}�k��$�Oܝ4�N)�^f6���xߘ���z��Ւ�����n�o\�ӷ�����̕�ן*����|¼Z�&���m���B�F���[l���x�i<cE�+ �W_���j�+�x;�o%tȳ���g#��x���h*��5�E�������s	��[xڷ��������Y+|}9��S�6$P��t�؊i�>�����րf�Y*{֥B�v�JP�����̓��nJ�ʂ����>���N�{�6�kb^�I�.�O�PSe-���2Q�ޞ�q�6}�A@^�Xi�y5AG^~Җ�8���(j��nB���q�	Z
���W�	�]՘���V���׃��kh�a������;u{�:2�ur$V�}�1N0R�O]��e�'Z��I��.��YٛS���,۵}�e)zD�ճs4p�)8�-��RN��ƣ{fd/�R����f����=�<�u��W�0k�_3[W�
/�����&�.t��W>7�m`w�t�_�F��O�bd��<@���7~��e�zr���]N��H�_@��ƾ���$}�Ǉ>���ɾ�d�R~,{���J�а��{�G���Ծ�]���z�sVl_yc�Bd.zWu��K$C��8"~�����1w%g�>���%�w�����*z��G�w�~��Hj��)Rn+��z�/?��o��:�q\O��^��͉ս�fim��F��fc����Fh#|/�	�ؒ��kMd�L`aU2<���n��赝�|7���=���R�/����,	�:�3�}�;�0;���79���gWj0H��ᮾ�ְ
��z;��ɰ��d7�Zgb����Y�?k�Y��yhy��~s��vQ*��Uz��/���][�x����P��o����'�E��S��?Ϯ�J�X~/�\�=�eO)(���;T�|�"5�ʽ�VGVwrRӴ��dфb���sIY����j���6h��VӔ�dN�N��ݾ�e4`�I��y�\�!��NY�4Dt9m��;���4Cb��oS�+g�8ί|�vvl���m}����3��ey�Xy�X3�s�ihI����k��o��K͍�� ������}�f�^�����J��/�&��
i�	�x��+g�q�X<�߇�^�8��5���a������0j��+��c{�$a��m�L�ϣrWwo)�v730�����o
�6:�7���N(�y�Z��c��|��WY�W�;|A���t����%�lݵ���-�/3X���̪�u����뱏8+�%g���%�y����V��e�}(�0�_>�py�}�-��r����eV��ps����Jh@�[S\�gǖ7�-��{7����_gx�(�D��i[8�����c�	k؎؏>��=��P+W�\�������6�f�>����� ���y]^]�K¥1K������s8�m6	�Q*�a�����w%��\H���!A&=gY����s��K���j�U��J�(����u	�����W��!�!g��uƳ[�T+V���hp�%ZwU��۫b[Dj�ݻ9��Z3����L��Ԏ7ҏY�}�m��}�R�^}�:��+
�,J��|0�岰�O{��>^+�g���
��}�u	��+��o��{ڄ�HwͶ,4d�vÎ~ڋ��}�z�w��L�2"`g/VϬyǁ�5xN�x*�p����͉ZJ�O� �ElҋKsG�O�`�`���	�����e~�hH�:���0��xV�?��,�J�G�E�g3��Pv�l�_��w�������)l� ��@��Q�xT�+����h� ��96�Z��Ο�B>��ד�� �t�DIq!��Wg���_X�"�1�����Xo�3M`H���$'�>���}�ي����
1٤��k�G���!
�_��oT�Oc�S��}��w9��}�����Q�*��(!�$�p�
ע����u$��i��뙇9!^A5F�$���CQ�a!�h2Xc�$5�6�!�[�n/�{�r?Zϼ�g<)]�~�\��U�ll��7{��]o����n�b�9��S�[NJ�����K�@T�@���Ԝ�2�tom
�v-LV�:V�Q�s��P��S�2�3� �vq�)T�~�%�>�!b�Z7z�_����HW%�#����(�8�Q^f2�tu��t1�����:�d����� 'i�nzk&�2��/`9.Gs���
�E"��s{��J�m���F�ta��P�U���b��q2�ٺ	n�Vܫ$3-!�NM}�ʹ	��Wm�����%	�(sZr_iW������g���2�9y������%���C��M6l��y���}�f�����Cqm�-ʲ�C��)��t�dB<;ckUZ���Z���R�p�3d��tv^]J�&9�U�p�-���y4�}����\}�҈�y��B5f��=�)�iuab|�e̳��+�f����ۥ��9&�v� iW`�Y�C�\�yٕ8oʝF:��>q���+.�����Ѳ�5[���ԤX�!�b�q�͖��W ��0����:d��t����l��v٧�0���K�ޛ����9E�Q�-��c��U�wi,aE��}gv�Hlc7������ہ����s�j|O=��U>��f�gv�Q43g8(pm�V4��b%�7N�5B�=ٛ������31��Lt�����w����a�k-G)�Ѐ��#�f��ܺ�i�\;اX��ͩ.Ť�Z`����f�_jC�%��/�i���Aޭ���[-���{���b�3���v�ᕅv��g�)��PV&�
���nH)�܊�뛥��3�v;�K���3��m��o`4�r�BuH-��&���B_%}�L#�r(�� k����1j�z"�a�|��kw+]�05Ȟ�w�m+۝u0����γǩ�>s�˚�1�n˩l�S�[�oq�v�9���WSE�³�([�^��2����<Ah�R8t���uШx^8չ���:���A�B�P����3���-)'Vm"®EӚ�Z�YN0�.t������OG;[��o�*Pt�J������n�V�yt6jR	��YR�T�7��v>%�l:[���C�N���gE�෼J	�Վ����ɽ�^6+F�d��LnW�r���Σ�m�x��n��9��\X놚Q�����9t;Zcy��Ԫ6����)MJ�c�<ܜ����Ϊbj���*�D��:,-@�C%U2/6�>W�N5	�z�!YX5Y�̒�c�؝(7����dj�|��y�ne���s#J��/��](����	��Rݼo��ԗCu�qܮi���R�\ᔘ�3��[/5����ź�*�U개B�d��|�o`�낖�!��l1�C���j��yדe��: 1,�Ʈ�rb���h8�p�@w�l��es�I��̸�����A�k5NZ��N79Z�96���3����Z�?G���D,����I: ̹[6��.I��-��a^E3�0�.�E�#0�u�ԓ�ʝ>=?g�����UD�PD��kUB���)�L!2
�����<�OS�D���,h��35kE�A:zzzzzz��:��(���XaUDF����@��B�W�A�NBQJ+nw4	�.Bv�g�^S]�*�F���;J��q3+�r�!��(�maQt�C=����c�'/�U��!�
��0��-t�(��f�O*�Nu/*KТ�3<��EU$�xU�T��^�]�B�-"�S�Ȋ�λ�Dg�xn��`��Y�-QyW2�j-T�S�u�i��Y�2�AEU;VJ�����
��TTRzy�ș	�QxS4�:TTyN^��m$ʹ��Q$3��̊�:!0��9���*h`Ra�d�Тݛ�M캗�H�X���Js��2�+Eݩ�rL�%�V�yB�/��Ϊ'YE�u�l���\f9�gY��Vowg'��S��l�'B:��t "�������f�a����wKg ��7T�d;��0Lt��r��r�V�$O��P��5��ƈ����_��'��ʓ�\�������>�$qꢠ<��&0a��x�x���ݖ�䖛�ف6��g����J���TMo�k�l��������U��G+6��&� M,��]�c�������6<�}W��� ��JѝS�)ٱ��;\����� �g�{�8�эЪ�1�}��xI��K�q?xtK	W�{Uס��yG^��F�|T�՜���=��yݑ�{m��8#�(��D�\+��{���w��*�y�'-��7�]#��OgXK�����;�ud������i���x.r�J�T�8kr"�3�R�\�S�=�e��,4������~����0����;v��LȻ���]�~��?#�����䵴��v;��3TO�������vɒC�<5WW��O�U������v1�+��G}���]z��lo��>AmQ�G�����g#�p3���Mw���c_��nt��jF� �]B�)�4 ����n%1�_��u0˨�#��*��R�%�K�o'f�B��ӧ��J�+b�`���6E�L��NQ"�����I��ֆ
g�"�y���9��_[��Ck g=?gДv�G'�;�;�^�^.{.�b@���Ԅ�i��Q�6#�^�S]3�������BP��{�y<i�fNQܗr�(!���+�C��Ə��b9^ӌhuQ��-���e�G�s8������a�ϥ�mD#1�u��u�x�n�7�Q��}��b1�۾�/~sկ����w����UMe��U\�S����jp'f�YG�iW`��-�L�ϥD�X�>��}�W:}s��d�q	����K��w��Y){0qn���k ���.�UU�_Ǉ=?��.��܁;���q��?>�+})3������R����\����:��=��h��a��O��]�������Ꝧ�^F=�}�G���0���t�����ː�����ƨӼ��>Q/�P�@I٪���g��O����t�شq�U\\2eG��)2lv��Ya[���c��C�&6��7W�
��*��#]�.l���;9]��Y�v���果k�쒦)���V����?&�F���1�l^�l�⫫]rG;�N�ӽےhx��B��M�TE�8�+��+�ы�c}1a�KbSF.��{��������/��\�	Y�:;���O����,�OϿC��v{��]̆F<6���#��Н	�򚽽��_�M���;oX�ȫ�g�*�V{Ւ�J��D>�(k�f� ��'�mn�~�槧7ſ ��ⶮ�b�����`Yߚ���Y�׷��F���R��DX~k �3r�4�dیH���<;\U���|��`]����Y4�K�Cv)��;�\�3;x�Ҕ�G�q��[�oN¢�6߇{e��ޡa��(w��+گ׽��(��@�C��Z����i�b:��fJ��i]��¥����т>�J���7��ϵ8���s�V����w��{�.}�C7�[�\���Bȁr�^�4�{l����usU��_v�&�n�n��ޗzy��gJ�,P���(Z���K����쾝��83����s�(uJ�ؠ�לvr������.=��A7 ����u�U�O^e��oxZ��\�\�zl�H�&�7�I2�'�W\�9R�j�(v��k�;OgS��;mD�@Wq�l����*V0������w�+�j>�z���_.[AH��zgwˁW�����-�Z��9{�$!�&lW�:;~�i��I���Pd�|}d�v��n�m+gWO���Ui�ʩ<�o�}K��Q�x�e�&�C7��8����<��D*_�]��0f|!�v(^��H0�c���+�������\U�eA�U||,��4ȟ^]��	Y�hւ��y�D�2���ib�g�$�C��7��ؖ��Ԙ;����O�1۬z��f�����\Ha��N7x_o���Y�;���ƫQ')�;�ׯ��8{���vk&���a��k>��Q�~�g=g6�ԵN �<����l�xh��ۜ�����tD����PZ�U���ɬ���s�o5�n�x.�ʹZlp�PQ����bc^F�0I���Y]��(|��-�`��&i!>S� �&7���mI�w�Bl��;&+/d͙Vr���S8�$��T���+�����O-+���R�|xة���b[P-�Y����q��g�kn-�ѹM���� �0���ݧLG�#����RC��|��a��Z�-��:�>1~v��z�_Vzs��T�l^d*�	�RxF��Y6��4�ֆ+�k���\Wx����Lwm[bNu���eKO��|��8�u��-��-��d{3����̟n86l���'OC�P2CH��z���jiӁys�����Q��tY;H�\�&��ʓ5s_.��N@}_Io]][�u����u�P��Y�����Uc���w_�^�[OD�Wv��]�E�5���b@�p-y�V�
6�IŃ�}�4��ܫ���s�vk�3�u��޽}+kT~��`]BA�u����}�D�o�\�%~�U�ؚw�f.��7H�0�����*��O�8��U=����}�zZ9�Ѝ���V��U�4�fmoҶ网Z�u;<1X8"@�@�����z����8琉��Ǿ7[J�bWu��]\J��X�%�&{�/%��r�%�+qn�'&�'���#����7T��b����v���ޘUAJ*�w.y��|�0�F�i/�ͦ�K.�,z/�	�w'G5c��ֵ3�sS3�
NI*�;��bkw���=�}��e1iæzh�c���~�b(0��[k(Q�v�`��	fA��vJ1�qx�n��x�Z���Js���%X���57}lL��k3_��gy�4{�[_a�z��l��.�-o�O`��T���\���V�`��是�B�t<P�{��ss��8��S�1�+���G�[ �+§Y\/�	���!��o �e}���}�;��~�3b�eSt�ђ|(>����#յ�5��f���U�ؠ��(e����_2��+��; Ld��WsV�AM��Bi�'(�v9PCpKb���D��n�o�z��\t5�a��7�YX:l�K��|�=��e�4��*��;�+�k{,�­z�65Q��Gkn��e�s�S��.��N��=�5�O�f�X^^q2� ��=R�}TO��Ε\u�X�ڬL��K�}�K��S��={v�}�~�W�PX�����f�2��swD7݆�v�w��렧���1�!������^�f�u��j���_݆c�CB�.ƪ^�o0Õn!n�6C*��s��ά����#,Y7��j��V����c�=��uG(D��'+�'�G���}���Ԣ����6�B[~��>�W]2d��_�2{�Y1�oz������c�Ƥ6��g�;�;碕�������Dg�}��]��_J\�~�M��8؃����f��������D��3�	0��*��ġ��	���y��8!�5��b|���&O�VT�֯N��w��]�^m�`�ڴ�8ǒ\-i�U�v��R2�h���zU#�D�lxn��	��jZ;�{P�G��A�/��o�D�]߹ǫ�B�5��>��]����We^n`���p"�B��ö��Z&T�5�����D۴۾Ř�M���7��e��WVߋ~��#�O\��
�F{Ĉ����.�	E�w&�~[*%��%f�`y��w�-�P�k�{'���q�!!�ωJ�Zme�纽��y7��0�:CK'*��MRoރ��u�mt����^��pl"��D��}��3���dNؓj��u�x�rfP�[��x�,f�l�_|P������N�9����x�l9/y"�m��Ra�o���s�}�c\�sf7Vɺ�iwo�Z�+:�=w�4�`�鑸��%��H��20�����Z��ϓT�QY�v��Ւ����E��w�H�c�u�µN �lBWt�P2�{�i�1O�9k��lU�87�.���FX]������-�@�T��N+��v�ߺ[NG��u���/��(����o���״I�k��g>[��hlBv�d/d}��4x�����`�+\eۨ}�"�O>8#��U�'[����>�J�t��w�����/>�J�}�����P�B|���uW�_C��Z�����1�q`��s��(�z-�l�*�i�8(c/Y���*�����r��*L-���דiC7�5�`�]-Y����-��YnbNg�iJ@�0�&����{z�xz��X
�
��L���cے�bX�5ऱ�ÿqLֈ?/���7��E�|ւA���S|��A��P
�M��\#�����/n�2�&$���8]����k�����˰ɮb�VO�WqF>�v|=W����Up�����$�R�ܷv�c�g>�8�-%��EӾ�N=,W5}�,�ÎG�����[���F�d�;IWf>��
��5;�6�
�rN@b���!�`ߦ��P��E�0����U��w]��������}���Z�k�fcl2�����:�F�i��v�f5���m����s}(��=V��K}�s��V��X�k�����oO�No���v���,�<P4��s�W���q6�*\��ٹW(�)���q���O��=�����xI`��|��a�$[ϝ��<�Z�}l_ٓ՗V}{È���Cr^D�A�\�=b)�B��*�&�z�j||}�I�=$mojļ�N��V:B	i���C���ljݮ���Wzf��{��.�'��8��Շ����6!GP��>a��~���O�'�{͋��v/l=�5�#z���(=W�<�$��JU+��M}��	�}�=���g�����R8�>[D��1y�]��ק>[~=�ݪ7�.�l�ٔg�lS�]5�X�,2�2
M[�V ���qR�pub&�^K�h��?Gz�2mN&Ve,l՝�!c�G��������fyX@��%�	5�ҵ�k�utb�V�]7^������>ͭ��#��dGn��%=��bwXR1Va�48/H����1H�8�;Ӥ�	o����]|�&ׇ&�iee�WCR�բ�t�S�����fn�9�}
~A��G����z�x��)�>Y��ߗ����p��rM��z�E޽����xA��S��w�u����ǎ9ܖ�`�ޘ%yR����нa*7�\5_�OLK��j�����wztu��{˶.ow�S�>��%��H4��g���;Y&�Q!��0�������0f�3�5w��{}>�|���16<JX�����{��>�{�+U�+DzD�;�ߥH{�Oј�V���}ɱgXV��&�=�Ǭ)����&�����J���\O��
��^�=���z{�qa�>-�x��&�+Q�Y{]啵���1��Q1�&$K,X��)���_X�a:T���tՐ�,�D�y��/#k>Vn�����fāAHP�-?w��>�umL'��(�N��nf^Z��3�TJ��-mjV�vM�Yg��zK}m�
F'&��̕�0�W#'5[u��qi���hnr]۾�ޥ��H���CY��5��T�*8*�n��2Cκ�̭�l{�B��7df.�p×����P[�瘌ܞ��u$����]ۦ��R�������h�E�w(y(���M�cD]�;vK�ft�}���]Sڤk(�U�`���V�5�gҔ͓�A�*������{t�3�}ٓ��o���!5�G�7(��8M�߯��֖�Z���D��Um�����5�r���AG���&��*C�����P��+m^˶w����E�f�v��+A�rdU���L�B�}��Kr$�l�zhe՞0e[tx�\�W���������I�m$I�5���_"��!}��eݗyHr�+'e�w���ښ�Γ]��:��L8s�*چ�\w%S.i����񹗤rz�P�U�
3e;�Ӎ�r��Tk��VP������j��rO%c��������@_:��ΧCK�����H�nL��(�ut�,l�;i俬u���ۮS�Rqj"��<��������_+.bĊ'��kM�b#5�Ң�tn���lm�B��ӵu{w6c���y��D���sd��s5�X���S��.�<���7٬k��Z��:sY��%�n��r�wW��G���j��hU��i��v^����s�'NV�c2�6A;S��Qshn	�m%�������:&r�D�ru�]cr'˴= B������}��!��E��u2^�[�`\ur�/*�cj�ly(�q���8��O59Q��[б�e����V"��}J˝��V�S�����n�S+��-�H/ʑx5|v�Ww]fUZ��	�,�غu�ZӺ��^g�N��\]�g�q_]�ji�d��V���wn����{Z:.��Q�I�SOa�Yu��l\tէ�-�M��B�=f�27P��789��X+slvGM(`�;���	(<�����
�LXث���[z����%fG�>��Kn6�&��Y��B����m��taއr���'j���b�rn3/r���`�oJ�ߠ����L}�s%�Sr��e�<�U];�����v�i���r��S�[�	���U�U\и+-�Z�:e�f���1�5��� n�V�ICL�����=�.�n��L���Z�7Y�2-Ų�gkY��׈��Gm
w��k����D�Ngh2�{�^^��K*�]�pE�u�2[:2\Jt]QA��j4�Gr��_	D&�=��^x�笫��u��7"�Vv�p����m@��N�&+Rt�F����f>Q*eG׫Mo��v��B�T�$��]�ʛ��.t/�
��@�.�W�evJ�����b]�E�d��u;��y�w�a����愝��ݐ8�L�	�>�j���Na9oD�%�u8��J�Nr`c�����W�UUSQfNZ'VN��U���&�"�ʢ:-ݢ��yE\y{}zzz��.�	���U5$���F�Ty�BA5Шh�*����8z(��xǧ�����K�i-a����)�:���+���'�I�B.I��9ؕT���QUEy�DTV��{�d�v��{3��Y.嫑����Fx^�vN��N��US���T��y�zEa� Ƞ��Ր�I�ʊi�ԋ�vC<L�+S3�tʊ/j9��u<d3�AffzHE,ڎ�^R(�Ԡ�AD����rʊ��aE�]�=m��=<$ݒ�#ʢ�2<�EJ���$(<+�U��O/<����2H#�K�6��p\��&�&�bj��J
"�5f�E⪇0#�򼬖�yz�Y^��d$!Y��=!�i2��'*"��Z[2�D��Ź^9�h��Q��[43�PFfo�+�,�L����@�)�����T�w\fv6����nf�r5cuT�U�:�n�-n������E�*p��_�	�������<	��'ܽ� PChKu�����'+޼���M�c=??A4��e��������{>���:2\?`ج���y�Pqa�oM;�����^2�w}�����E���ۏR�_�<�)7L@��J��d�Q��v��cj��Ʌ2��s:5���{A�:������U|G�@&��WUs�����ޑ��}~��o/{�H���Y���V-����	����y[=�mW�g�����ӷ��1|�hM,�M}����C���>3R|��vo���.��k��rz"��q^H��u��?7%��`��F�G:T�ݾ�����w��1D���e�,��*"��e��������F��NF��n�Q=�A΅�*>�+�Z���j��!a�zs�!e�D�{�I�����"��4��݀a��G���x�vk�Uե-�[�:soe�]����ԅs��������p�n8�҃���8�)e%B��@u��ݢ5aX}aV'��ب0�ty��U���0�!��`G��%��#�M���?_{��_Ǝ�1�7Z��y����8�����8~�Y>�b#V'�����w�W����Y���`og2��/9���u��C5���Jw#�*"��v �-v�6z-��uI}@tİ�D�TFy{r$�p�~�$�E�%�A�|
j֛Y�y�v���Ȑ�6W��٩�%�e�~>yG�<$�9�;WX͵�)��L�+2w���nE+OF���M{�#��@�[�Hޢ��_wSKL��'�㿵�Ѥ���9�U�osT.��)i��"?= &w�zU����7��(�Q�M���ꃦ1u��1��������? ��I��ڰ��io�	@���glUVO.fb������(��_|@���@��By�λN,A(�s��F����ܒN��R/5��>��ks��	��Kռ�ˇ_W�~p�~�3Wd��O��s3��-c��\���5dA���K4)Ж~�s�k�[��~<Wu��s���E��Ź��OF���S
1�{m��q�֋N9�u�p]%]�S}]�;��^H�B�-�nE�0�h�t���������d hd�F��ߧt���"�Z��!���|��N=������4��5�q7k�׾��$8z0А�N�o�����3{��m�y�^�PEX������B�%���*'S����5�9^�������U��z�~�5f�1(:L���I�R����0���şW��i ׽�nL�F:��Ό���~�q>ΰ�\���^�Rt�
K��o~���S���jo���ݙ�=Y<�	��ԸM�J��,"\X�c3s��'������8�8�Y:sy���W[`�m���ڹ�ouXl�/}���WTa�ur�c�@��z��F,��w��MEzk�����oӮCǮϯ�sY3��`�fe� ��V�G��tC���<�*�l`ӈX>f��t�E�őK΋��_a���z,����ߪ��{��+���x=b)���b�ҝ����2�	��B6�̺�-�`��[�Г��֯:�e��d��љt�� &c�۫�4-�D�=c�a���d`��wK}pkf0�N���k���g=��C�2hR�i�FPw4Jݗ�"�dyeo]	�y��s>�ԩ/y�@��{�,�g��K�������V�T��(�r�����;^�{Nz`y���ުQ�T��a-��cO~�j߻�t�У�!���lv׶�y��G�Y����f���%�޷�kQ@-}W�4�|g��\���Zݨ�D]�G���yV?6D�X(u{�S��Y��3䚫��6Wu�zp-��>��ח��:_��=S�������o���]|���q`��g�4��[_D��P�Ϻ�^����>DA�E-�T羀�@�k�=�x��)�����"�����S�	�N�%F+��ݦv�hGw�b�A��{U��?_�����<�+Q����\s���>����Q�:a�s��i��*�S�~2}�?v��娥oރO���ش��g���;�$��bU�xW�ߍ5Y��'R�_!,�e=�-���1;��K�)��c�Ւ���
���i���~���3ۧ�v /��Ģ�V3�V<8�����+��܈��(��
�6��dVh�5�4����2t`��Z�'�a�Q�TH�;aly��38�Z��K]�ޕ�#������̂���ͮ��3�`�
��ZM1�G{Q3��,���΃�3;�
��s�^�M�:´��MzW뫛;��>�;�\�0=����z>š�7>���a�:�փ�ĺf�yx֨2��}���G7�y.�C(`���m��:�h\��y\o뽁sj;�UsVxsa���6��5�7�K��}AK�0KO�z")މ��$W��L�������I#�$��Y;���CF\�*��{���i�|��P^���liq@�m��YY��cϛ:p|�=�xaA����!mo�������u�o�4��ݭ�.�i�P�ԉ
�'wjɜ��r�.����S��Ў�(#r��lέ�K�:���-�P]EN_H��G��LG�f�3=;c��q�YW�|�mb3��h�=7� ����iA\Wgy#�U�ӧ�=��hC�Hq����C�0��9��2 ^};�Ҭ�/B�/�n���=����ԅ]L��м�g|=��7�7'X��d�w�&���Iȍk��r�&��*6�0vVC�2 Z��k#��LFk�M�����%�d��ރ�τ����C�8�.��RN�st�1�˨g�{������D��`��G��f�ǧy�إ�z7z��G7ٔ+�����>9�����J��vtF��s�O�����f�?�`a?D�9Z��$զ�Qc�����s�1�X;����=B�$T�^Of��w/{P�IM|j}�Sr�p��Hq^���]9%����1P�֦�o}��<�	�n��o��\�B�o�!�_�c�3ִs�����X�̴�^sUG�.T>�Q����f�A1�˽�� �k��6z,#�����v��JI^uu�tb�������N!|7�y^F��M_ޜ����u혪�0��=�����R�9�����Շ��}��	��E}ں�iD�Bi�TVd�6�z"v�y	�\DYw]�4�S��N/yа�BRԃ��´wSK@2�z یw/sK�н�dT���)����Ts8�p�Cח}ɻ؉һeI�)N���^�����y�_���J����1��,K����ڈ�wY�X���8��6���e��d_o;�2��çeI�U����T���C0�<0]��9ř���: h��;}ǈ�`v���#�<=<�Kf��@ޕo>��ۦ���!�N��l�����n���yzSc���$t����n�k�e��MR��&U�>�7~�~c͚����6�˱�}���O>#���`�s�n�j�K�U�v��j�}8J/5���w�דh�x8�ն���W�������^��>Vؖ�Ϟ�D��m&lp��"oNl���>���*�a;��~������am�i+ �mg���
�{�k� 샗m.�́��x�Q��?h�DG�9��Չ�i�C|=���9���BF�xN���l����}rhnE���69���0�j�v��o��H;�=��jwc}9��^>�^�=�B��R>B�lXh�/��nM��$0���N73>��c}����^=��m��䍎���ZՕ�"\w��vk'�,��s�jC��39[W��#u�T�ۄo�N��2�mu{��vސ~2�)����疓�+v����%P�m�3��F�Y����T��Ƃ�^0�3��]�6��һ���t���5\�hG��t�e�F���e��*]��}�kj9���{$��4�%u�}W^��\[��	f�gѾ����WV�h�K��y�bOL,B�˦9oz�Ň�ɷ�k���\���<�2�S�/&��4�����v3b@c����`M���,3b��MH�s,N]����۞P��i��sٷ���O���C��R�Ń��g��(������e��x�Vg�PSE`]j�)���ܗc�BR��=���t#�AxR^��p`�;LW��)���O`ڰ�����������=�ޢt��<r�K���?Zφ����c�.zJ�RZ�]�x�Nz������`�ގ��������y�^��+�g�z�I	�[ե����v���{}�f��}*��r�8�m�sݻv$�Y�&� M,�����������?Z1�C=C���*�} 0e��Һ�o��R� H�bT����oE�x��5M��^؛\���L���HB�����_S�;W1�*�Lx՘�?u:�è��n"ӗK
nK��szJ�ognT�J^Y{�4��U�2F�67��Yp�beD��ܥ�jZ3[�Q)]ٲa�&>W0\��rGSj޴��{ߵO�1碁�\b~�bBP��u�~���譈������������o�C6����Jh��.�?t���jgNy{ޱbZ���<N����]Γ��tuku�ذ�:�������z�������gZ��$���݆��Ǡ��q	��JX��������HЎ���G o��ۉ��L9��ѣ�ޯ_����%����F_���0�NmpK��#�k!��R�wTX������;����� ���=����|����Cʍ��y�;��o%^a�G�(�`�hY�n�z���r}�|g��҄��x��o���6�=������S7~��d������6�a��ͣ�	<xO2NP3��<��P�E�����>>iY�9�(j�B��Hu��W�Em�a��mXK��|���+2 Mu�?��%����^���h��Tn�`�5%���U�7�kln�OFB��(���|R�8H�u�v�vskZ9mV��Yԏ\o��E�9�ثyԛ�oUL�x�|��zV�p̛��əo'�<�"�R���llQ�ܧ����1�����Yb7di�x\Wkn�e��u#��}9��"�8�҄}��N�*a�C����ܢ�;�]?i>73��hV�7Y�D���Ʀwq����h0$��=�3�Y]U���*��JP �3s�d�to����ȼg�`��<���${�C܇YA��߯U!YʌX�p�;���)2=�
'0R%u�6 ��wٍV�]�}�G^�^��B_>�)C� �u�4rm�N[t������hB�ә��^�T>텂��s��&��>S�=�&��d�un�K��~��& �&�v\b�A�T>I��k[�r��jc�Cz}��Z�*�5�В}~����}���{}"k�U1�Bw[���{ǘV�o�b����]]߼��%�X\'�{k�%O���	̾_�����?��� ��򂨮�U@���?��
�����F��g����TAEbaA	�`	��&f�G��@�dTt�.10���Ī�Ԣ����0��ʪ�  C(��b3L ª�  C(��
�0��0(�0 0������a�UVUX` ea� !�U�@ �EVUXeUs0��  !�U�UVEX` eUa�U�UVXeUx�@� XeUa�U�V UX`Ua�a�s��Uִ:@@�@�7Q���0��?�(
��2 �p<O�/����������x}G��������?��g��������ɏˊ���W�?��~g�����ww�~��������Q_��H����?��2'����S���~�?�U������?��7u�������?g`�Ï�����{�� 
�
ʈ��	 J��
�B��� J)*�2�� �2 �
�K �H U1�A8���,��_��O�*�
� O�|���@���~��������w������?w�(*��~X�'�����ٮ��	������G�z����Ex>އ�O�볏�7����
���y��O��"�}���DU�~��&��y�w���G)��<?@p����a������_����Q^C��b��~?�}~���C�~����ϴ?P~�?@<w���*
��~�d~_̈*�����]!�^?_w��������~��������I��Р�+�wA�g�L@�C�>w��{_�G�}'�W�ADE8��`h>�\��"���~�_�~��=O�����)�׀�:�%��8(���1#�|@  ��@ � @    �      Ҁ 
 
    �    f��(�p��d�>�Wkf�t�V*�+�UVL�e�-��Zv��m��ҝ[Mm�4�ū�.صfi�kU�&�M��QN��dڱ�[=�G0Ѧ{h��v�[M����Vڛ;��[I�)֊kf�km56��&ŭB�Xʙ�6��m�f�T��f�M�e6ִm
��R�4���V�Z�fFt�P�Y6π  ����[MM6���Pֻ�:�ݎ��F�I�;v��Nۦ���vi�S{t����I�v̮�Z5�c�u����J�����PSO7��Y�jڌ�z���;���T�Y1���l��   gqȾ�"�J�CFC�'8��QDIJ�&t��D�2I	"$D�y�\=<D�L����������%J�7Om��]��V�#�^�;={����Ξ2Z�m��y]6zkl�^��kۭ������[3+l!M�����4z�j��   ��J�Xi��l-�V�����v�ҳ�n�o��z�n��˶��\�Z����u�7f��wuӞ�n�D��m]��w%.����{�{������ҷ��Ȯ�f�,ՠ׶K��j�R�wj�   �}Ү���U[�-_{W�m^��yz��5������s�[�CX����U�t��Zkj�v�[m͝c�Z�6���xsŵ�#0v��:��7=h�޽eie	-����l[3J�Io�   6;��Ϸ Z���n+��NZ�n�k�Vw3�fX�zp.�U�S�{���޴�U����U.{i��QM�ֵ�q��ia�o�  >�M�{o��Ӡ��5� ���iT���w���[�j�O���z�G�m��h��p���]�1�ס��*�چ�w{�n�v�Wm[k5�V�AZ֌�  ���.܀�κ]4�}���2Ѣ�늫�6��M[5�x��* �:7Y�چ�ýz�[w��64  ����A�1�Ճ�Ԗ���[��[[e�   �� 7��  �׏�F�N lo[ozN���ip�7����A�sA�M�z� ��v�t����շn.�F�Zmm2U�T�n�  s� V(Ə���0t �+� ��b�t{���= (�C J���SN��(�� ��{��+Ii�,�fm�e���-�   w���:k����@ G�  �w�7� �^��J�h`�:�/xt ��=����< � /y�+O] 3�S�)J�y@���i�RR�  S�b5)J�  ��4ԥ)�d��� �*   e*
�� '�����D�c����t���}�]"��1�K#j]R�J�U�,�_��x{�q�����m�o�1��6?��cm��6����m��dcm�������?������r �����d�Xc�4%����K�	�b�@At���a4�:�7��3`�(Fh�/c҆�J���QZUi@����B�<��Ǩ�4Z���#�ΧNY��Mԁ7��S�ޯ��T{��X� 3��Z]&�\|C�%��G^7�#���͖��x�h�Tv��N���ݤ�t*��N'w�s�@3�pq���1��o6R5-X2N�����&,���{��T�㙻F�v⁧�9ga<�	�����9닉/Ē81��Jtq�:*U�\
�LIe�)��v�0�@+�t2��y-[0���ni퍖ʊ�cZw_.����p�Ց�:l�2wp��N��Q-�����L"�ƾv�+\P|���Y2�j�H\�ts��.���;M��>̿M/un��e:��wz�O#�J��7/i:�8)k㉶.�r}~KA �v�Lx\��(�17N�5�urt�����9�b8�W�\E9ʄR�N�K���j��h��w�b�uK�^�HE&m Xk���闸����n��{���n�ݩ��n<= �)��3$Ω ��<;��@�o-�6�l�ݛ��abLIQ�p'�Mvȵ`Қ���6�v^���m�­h�#B��`��7�X.5�jh�$���_��4=��zf�#IЮZ��Y'Y�[��d�p,+3�.<dŝ�9hYv�g�{9�|Vj��dS��7�B�,����J촍;�IN��a�Sv+���V���vn�aDqg��Ms��a� �ɘK��3�^�w��i.s��懈*�7��ǚ[f=O�pS8� ��o&������ǳ���C���Xk�
�.���S��+xUm�f%��H �&���Rܔ���˝�tkN2���-WwOr#�����bN`lΫ᧷G�uh�n3n��&m�	wR�ަv9�7N�T)��뢵���	A��)����r���5�5;'�pr���3�r�S��6:��G��voæ@qZ��I�
�[�ܲwn#	�*���"��������=DnJ�U;�\�D�/�����n��������2r�A�!�&���tG���;��;�V�;7L�,m��sh�x嘻6�9"��w��n��C��������pb��#� :^�yʹsɜ��r����E�-O ���t�؅��t��89PJ����Nh�fjä�Z��ܬ�����N���ߠ������G8�"a��V�*D��	Y�6��O@�tz�]��EZ�S\_	N�)(��D$(
��z���S0KBk<Qf�h�7	����j�Ѝ}u��q�:ʫ����A�)TF�J�^%2�����t��é��K)2�x7���M7v�>����Ĳ���N�h].�r�ܽ�\t#6�F���5�mt,c�*�`�(t�/Fm�(�N�W){���/�;{��G"�:[�r3��id��W�q�_Ct(nt��S`/y$1�k�^:��W���3m��umֹe{���4�xjv�2��9uvN�U�՚͙�Z�v6��H:�apMב����:'�qh���a	J�=(�,]���-�t��!��k;���B^݉�vi�_h8��(�ݚfG����_7]���X-�-t6fE���F�·if����Λ�!3np�q�^��/��4�.�1E"Je��xk-	W\n�N�J�����/xg.�ٽ�tep��RNt�`Q�� �ɕ>':��J,F�õ!��%Æk�i��/���h9��s/zW�R����p�����N�Jܙݲ�n��̑Ŕ�sÈ;q��������I6�+�կ;�����4��G��;�cC�L�]e[�|�LJ�^s�r4�O{;�4��r5�%n�j��Q,�H�Q�[���G=cO%��ӭ�x�UC����W=�Z{�Ԍ|��	��z��;�j'�����W�()�(lQ3��n�7<]���7,1��)�)��"�N(I0̰�of�+���r�q��&�{u�/"Fk3U���Έgئ���ba�9�g'�2�M#Uݚ���0훶��| y/��������<�[�fܻ�-��8F��o#dɠA�hK�����*��b��H.�iu˭�rl�N��\{u#Qy��#T����{��'��dأ�d�)�x	�L�4��{6�1 ڗ���o.I;j�w-���-��3�8ї��299	�ezw��oE���,^:4��o���E�8��`d���V類����Id
7��6-D�G ���&��=�ݸ�N����������p��f�ۓu���T�,߇p��y˅��7�9H�Yj���c������#8��ɭ>��[�e��>��Z�NCcqRZJ�|��z��-�{���Yۣ�_9wZ܁W�0q���:r��M��hC{'l׶[�l�U���2���$�(�
L�2�y�L�M&�.�,�RĎ��ѹҮ�k}���	����[i#d�Ր��
@֠/�9�����pqIw^1Doĺ�9Iu�:�Q't�p�4�/Q�wA��x�v�I����=��;�7@:77/0�VA�-��Z��9��ˇ���Λ�ԗlOw{&+��\�o�i�"]��5!;%$.:$4����z9���s���t�h��Oo�XD{�q�.��-q�˷��分^�٦��{�F"�`����ǋ�'R�����]#������Oh�wy�����S���Cm��y�`xcֳ���W����lCN��MC�[���ވUk��;y�q[�팸r!���8{�d%��Ͳ ����N"��3Wgr⨸�-�k:^k-QnR#K�jwXf�v������8�1>G6����G93�Te���P�f��kF{ܥ���F\����8�n��<nk�X���.�y!8/7���~�=��bLݼ_3�� K�\�Q�5�(@��tb��;���5m�Wm��F�B���94��JE��v��)� <�D�?q���_ ��������c��9�u�ܯ*C&��n�5����^�;���:p���	�3D����1j���]��>/R�_��S����l�,�s��¿�Q�_���9�9��Ph��K��B���O���}�E�n�UW�7�r3p-�e`���G��r ��Btw�J��同�Y�R8J;�uZ;/�pa^m�w&��E;�7�V�m����dx�\`��\`c:������)�F�IL���?\/��s�N��Hk�lZ�c� ��1��GR�L p�a�נ��pdڙ��k�{˖�'����g0�ĵ�F<�_33��r= 'J�3M����C�9���<[t��Q�+EM���܈Ȇ����XãySs�+�� ԙ�@�%l��Aֳx�:�e�?Hf��:Sjsx��w:ӹ���u-[��9,*���DB1ݠd�ɇ3�(� ���vkn���u����4�&��;z� K��nS	���tַ/;k��˝��!�̯k8�Ob�)ڧ\�˚n+Fʶ�Q���߮�8��;�]�E�L#��Kv����Ὁ���ټzv-䳄�f,��-a0H𴚊�4\xގ6r��.-�[!v�9H�n�/�ʉ�d8����_���5�M�E+E�h��/�-�k0�|V�S���"��۝�O7 �v����a4߭Q��>�7VZ�,ެ���mɌ�RZ`�Hk��Y3B����էt����n�^���EN�nm�>�#u��QN�v�<��2��N޷%:��H�3G`�v���52���9G�^�iv����Ƶ�"��0�2.��k�э��{��:pv�TL���<z�c���և�wan����-��2L��';����	YZ�f���t�T{[#fQ��3�Õ���=���TN58��,�;���6��,�I�~�)�4o3[����J��Ƃ�01��^�1�'A-CEB��HēG$R�ns7%-a$s����\nh�<�{R�<���8^�8���C���ڥŊ�wո���!�� m-�w[�a��b�;Fp���b:Ogol/�ӛT����t��$dH&ua��&����
s���wF
��&N<�s:D*�fpˡ��BgR�kI�m&)AF+��+1�u��z	�L�Qo��;��\�,����R9$�#JP�O����@�������ak������yӻ�X-�mX��m0�Q6�zsj��j۩w\.olcQ�B5�4GK��N.9���S^���44�a�D���{4b�w�7��; ���0��,ݚ�T���d���ɶ�76��`��Y��.	s^	2���mVu�������CS9TY3�����l�[|7�q%�d��D��2I�����B���#�,�#���I�q2�����Y�/f�|a��Pn��"��3Z�e�֢Z�!׻���ߺ[��:9�l�)�,ӻ�aw.�In,�7x<+��]��:^��e/6"�u����׍F��w��p�awz��@,@��������oF��@Ë�F�ľ�wHIW/ZG]f3!�^��'��\$u壸=�:�/����Gu�Nv $T��]�t���w+�됆p���ݔ��ΓH��
=oV�A�XWC������YԜ;�5�8��� ���R�oF�6F�nu*��n;F���S+1n�k��u�ru�J�E�Q�nW��Ƭ����i�	u��p�s�Z&���V���)�"�9��Fi��pXH7V��ڏJu��b�O��C|4K.�
tǏNɕ�ٜ�ʍ�����N��{�j#�Sd�f��(񢩜�'��6_i��Fs3�\z�^��"��&ٗɻʋ��ʓ�tj��{_�b��]ώ��&6���6f��(��V��X��#\�s׈Bd�m�r��W+� �Ϊ�V�q{��ֵ��N�W�}�9�B@ҥ��< ,�-i���X�p���.};��k{Hڗl�
Z��D:��"���=p��,aV��2<��ګ���^"=��Oצ���qM����t��^��3�и"�uء�!ǌ�3K5��[��MO��T8���Rݘ�)�Ը(v󎭘i�I��Ï��S��'6�$3��A�
��6r�"��3V1�i���p�Kx�7][Ù�e54\�؍�C:��⭊	�=�w&�	��|�q�)^ H-�Kj�-�`�J�Kef��{��)�m[�H��A�]5�f\�C���!bj�����lw���*��"� ���W_5_<��#T��n����Oz�0�1.�k�*��[y�-�]�Y�Fl�9w]v���N8qƀ۰����J���p�0�<J`E�u$�\u��T�h%��4$ ��t����cWvM�׍I�n� d.��vL��V�,�:�N����RNN*񮹽��[+[�"���؞r	��bgoK�xH�XhA�zoge	ܑ]zk���:��tc���E�:�Mh>Z�
[ë,�p�*4^	��o�$�i�E8k�,�s�h��2�Ii�Wgl�.�y7e�>�4�5ǥ\Ѧ1�U�P4MqBIjV]R�9_,כoUT��FD�j-��3�dM8WV��[u�A3%��f��l!����q������w��q΋"djEJ0�uҤ)������^����%��y37�zl��*��;;7&��+hU_�v਌�6��ۤ��{B�Iq9�p7����wL�F.Y�q�X�@�Ʈn�y�� }�8�Fk�{!!�����d���
h>�3�L{�"p^�hҧ;�`1�X�jУ&\���X�W�Rׂ�Ӷ��vt��ɜ��"�ۮ!r�vcpr�{&�wc_�i;��m�PM,}^�
$kս���ӛ���tޤv���*����uA؆��;;w�����"Tܪ���U��e>Ѫ���X0�"g#�c(��(���Q��+P�� �>$���N��y�[�͓*���JF�o^���<'m}�%v�9�l�!qD�ce�N޹��J�`�6���n��k�x�Ťs��L+� A�0P���&i��K$;/1�gp޺j���e�.�&�Ͳ�8�Nca�jW��HkŤe�X�Th�p����:�_��SM�v�c.q
|'k�X]!J�3����/��G��V��
�{�Wœ��lSh���@����:z�[&�Z���|��u������z;���} �Z�{�����I�ళ�k��i���<��3�(t����V����r���a8��/�A�ץ���Ӑw
k���.��<�D���mx�%��2��������}3ݜ7/ujcgX�]`�d��y]�S"N;swɢ�o:t̮wa�хB\�*m�E}͙�E��-Gg]Ot�ʄ�
Ób����ͪO���ѐ"�ոr�s�On���j >G%n�����W^ݓޢI��ת���yP�w�,6.^��qƢ�ce�$���%�hL�vTy��rwVU;�N�G��"d���wl�i�ū�m�ĸ�_uǷ�$*��=��9q���$t��������ז^37H���w���nn��6�-V̈h��Hy�.��P�^z���xv��r9�|���u^��㢩f<zu�����Ԝw#��.o;z[=�d�s���[$��3�R���ʹdѹB��Of9Kp񵳝�Z)�z̦�û�D���^�b�N��֯1��+�(g\���CT��"BTc��'��&2��ˤ^@w�X�m�!�0�ZO�U��tSt;$]�߯���'*Z����^P�Z�u�S,����:����@g�c<0�r�2p6��K�\�Jojg	M5��Mr����ƞ-D
D���̵�J�*r���ӛ�P*<N��(r���Ψ��(l��uLKyP��r�H��͖�8L���]n��ge	��P@�뾆9ھBI� �E3k1��o-��.&!����N�+#ףl��0N]j�غ7�sbt�����.N�C�Q�k{RG�Eh�����4��R��ns7:�a�}�tI-�L����Y��ʘ1N4�d���Anԧ�������ƾzs�U��_���^��6�}�����<�[{/�{s�qH��O<�=�GnJ�������,�yA7�s����e^��ŀ
�'Tf���$x*�Wj��?����st"ؚg\�A����puڵ�T��c�]i���D�b[�th˙MT*R= ������1��.�P�é�f�8�ړ�^��v��y��y�/t@���:l{ebɣ^��؉�&��_:�8�2�'`�4!1Q:f`��xg
�UA�WGlv��*1�*TS k�{����[��oSȲW`��K��b�x5�H_��y�=zM9�PT�k�TAٜa���b8Mdk.�EJ4�VZxnuq꘹�#�&�ؖ��y��.g;5�v��'d��8�;����fвh�G��z�d.�#�������Y�v:eƝ_>an��l�2�*^���h�h��^�\4��=L�%��2 �|�uv��2�	 �w�Ȱ3w�\�.�5�X����ѩ�`ν�M�ȃ�i�^\�wq3�L����Z9y��Z����[*,Xتȫ�b�"����s��y��������N���z�4dC��s� �s��9���v	<(^���l�x	Wj�#q��>6nh�nQ{,<�����~t�S�$W��$�M	�Ih��Gy��?:¨f>6�,
��!ͺ�3H�c+#���eǼ��˚"�x/+��jn�v�j��X�252���u�#NCOKX�F�^B�K����]�eiYLfGp�fx:w`9�����=�p�B��Ww�YJ���ɧ�i\��[�oT��.�s�[6P�(�F�5���nz�Vw�xN�~x"`a��np�d�7��ۣ�ƨ�:�Qc7s�<�"�Y�~y'Y�qȨ�Z�L;�&��ʏ:�i�����zH\��'�Z�Ee�g5Q��Y ̋a�w��b80d�w].ǔ�t�w�����?9\���m���3e�m���&�Gu�&Ku�y������2঻��/�U�뼝w�Y�=���&xV�����y��gN~���V�����۬w����U@��9O:�GI�f͗L=��{��!��p9�P�Pc8���Z:�ŵ+�@��[��y���z�#
�/r��ts\)��|��VS���4�� ��{&, �=����E]��|!��i�}�I0e�AŞ�G�o�K�ݬ��B�����<�}r'=�.G8�#*P%��>ԃA�Li�^n������D�6�.W^����d��owl�J�h�Ԕ�QR�sp���&.�{�d"�v�]�Խ�o�bH	ۂ�Ĭ��ϥ�Z|)�t컬�L��AYȺ�qb�"6T��I6%}1nӇzܺ����B���cⲭZ�n@��|-P��gN�D�C�������#{K��WrpE���rO��Je��(���8��4һ'�A�g�S�,���K<e�������;�D���x���'����r�K�|���K/|&@�������\�����z�����[����2ֵ(b�/r������na���s�5�܇��S�qv�[Ֆ�F0�!�De��p�'��T%b���)%���� Q�`�r���Gh˛�3�ͫ&4��WU�rA�}�&�s�x�s�{�󖍗�I�?d�d�\:�:31�u�_ME�o�jeS��1,n�h����#�Z}�˚��B��a+F�C�ywy�7��g=�7*F�����]�3�H�;���&�)N�'�/��] `��=�� �HK�r=�K���z�O��!{�Nt��l{&�Д��
�.�YIl[Eڏ�3ջ�P),�N�;��r�[�)�z��S��\�a��:�av��ˊ����d���C�MX��i^Æ�ݛjl*�8�6�R9�����ҔN�׎�9��a+6aZ��To9�e����]х��c����Y���d8�Ƽ��gz���W;%`	��-��c��|����;�S�k~oXS��Ua[���T�6&���3���_ly���iE�q�˽�y�,Մ,5���$Яx�=�f��b�J�Ӕ��ؠ�PT�| �f�\K�F�5�M*�*9���3e�'q%on,Wơ�U`r����Zs�u�6Q�:�G	 �6r���#QE�1N�o=Y`l]�,@�ٙ��xr�툉J��N���$��>��<�|�x��]��p������%�����E���h�{F���q�잚��a�V�+)�/��2��k:���\���zU�� ��֞jr't��Jx��}pl6�8\Y.��h�,��q˻E�8��J�͓w*M˂ -jꊜ�j����+qZ�F������3�ѕvl�3Ʋ.�:��ȮK+����׷�����7�B���xrאf������;H��=78��q��C��0C���n�ܭw"Z��V<��M��:�hN6����T�*�4StS���9c���9ΐ�a��3G��u��D�f���O�#L�VF���裮�0��x��\[�#q��������N�;8����.����B��\�kcռ����R:na���4֗L'.��)��)*�۹L+o�ا`���L�ئC�r�&�LP�\dv�7eҔ)�Q9ϱN�����+�;':�"Nڷs%���5�ub[`�C��H/9a�6܄��|�bv�#.w��<[��-�J���~�k�+#{=x����؛���\��n����s��E�0�Î�훥�X��˃���G��R��׷\o���7'.(G({��iX�����Iсr@�I�ǟJyӮ׸7�H������)�xP�<n����\�OϽ����S�'�'���yO-�~�LY�VV��:B�٠o�Ć�y�yP��Qͺ��Ok��7p�=���[����b�x��gh��Y\w�GDq�r�#$Wkl��ͭ��d��YN�n���o0�5F'�>��n}�Y�2���9Sl�3���.�$�w���;�N��ǧk���\���+N�'6�H-ɩ]�9J��Uc�DCz/-!�5�^�Z2�U��T�F5�N���=�b}��m!>��<�[����q �uCi\PH��̏����o��Ł�=M���m��Ϲ4/��ˍ�ս�
{�{�S�(ene�4��$����:+adȾ�&^�bMu�yu�"��hΨ��Y����D"��{r�I�dG�V��=5���5&�S��/g�� ?xP4�V(�vbq�t�L���n��z���q��3�P�d��m;���Z��C�������-��񽻂SJ��e:�*-���S��M���g��2!�f��j%�x��J�6��]o[���QmK���p��x��k}K,H.��KS�F��70`\�u	�I��4:��%iOh�Y�sR�N[��¯���γ1ټs@i|l
%�*ck�j�'sX�S8�H�F ��=F��ugF�#64�e�����}7<�A䉕Ն��)E�YU.a���?urU��<1U>{@InNǪ��2��G�����^����o��S�{! ��c��I�f�r�9�v�l�;I��#rT�ld4p˖�m�����V���:͸�nPJ�i�����++�}��=�bX1rT@�DSvW��i��R�Y:�u. J�*6Lؕ��[��-`!�8�t�PY������#����+?of��Q�N� ��Om�:!��R�1h��+�����U%�����gV.!�����\��D>���ݶ��:Wi�v"-�UEt���;��HLknE$���M#�a5u���t^�>� �ޑ����`/n��k�p���c['0���$PO��ь#���:/��=�%�����M976��N��5x�s"�V*o+��&�w��sn\�]o4mB;%cA(�v!R�O<3 (.y3�v��Z����^a�f=��}{ا�������⾬`�!�����ӯ�I�|X����Z8iZ栺��,Z�����o�]��h��!�WC��`�J,�ۨ:�{3r0��G��x=3�y{��GTI�xZ�;Vm'���T^�<��\�Y�B@���9�.n�z��\�ėN*�f�v##vgV�,i���B}8�z��ʘ٭��bB�֎�%c%h
��!I��5��-���-0��ӷ�i�Z����j�����H�
���+>�֨��r�������峻ԑ����w3L9�۽���Ӥj�1�b�|����o�=��q�ё�
]6ޛ��-�F��65��Z� ᩗw/a��9� ID/)���+�jl���ސt���q�.�;���=�<ӽ��-^�%�ZВ�%0�WE�gwg��s��#ۧ)2����#�
��B�[�ϝ�I��Ӓ/&{�L�Vٿ08[��ЙiVB�@���2U��M�����A&`�!�n����[|��B�7�čT�N�޿������{�:�k\�}�!��.�~��h���󷎻�1���mՅkU}�U��go��i�=T���J{4(��ԎYp�`]�i
�a�;3��u��N��9d�=��`n!�b�(�z�\]a$��%�xr;4��Oƈ<vվЙ����`�u��&?�@�n�XU�^�vp�r�⠷eFer��=�QmY��sef��q@a��v�iƠ�Y��$:E�˷|�t�!.���Y�Q�$3�9XP!�+*�&�g�)c@�1N��*�X�[��M8Z�:p�%>�M��
O ��]����Wv��_OL�Ն�Y��Â�S��t�Ee9Vzެ�D��	�Nk8��ʹV
���e�cA�S��7�+� �9�|>�1-w���ݏ��9�m���f�i�[@�=ɸ� fE_=���S�q��C����d���v�F؛���:�woN�m6�t�.>�8��ŝ���;��.�e;X���g]��ĭt�ɲ]	A���󋖙�6Y�������aGMvJ�,�H��D���6�b1�S���*��Rf�.)�lk*�ӌ�A�Tx���뷞�.��ڊD�H�ZJ�c�Iu8t�w��<���&�;��q���:���ms�t�GP�S�_>i�5|��&s��'d�ũ>�(�g,}18S@Ӏ��ٖ2������/r��Hn�{����t��!�<}�v�bX�Ĵ����yr,?$V�Q��׽8U䵺/1pp� ���e NP�E�U�L2��s����ͽ�ӎ|� [��E�}�F���:3�z�'�+��!��O�+.��;->�Ӝ�?]%�4U�ޒ���b��'Ay9��O_;��"���՝kLUw\܃+fc�ڒ�9��	�+��;����΋̼�Ҵ��o��[QSځ^U���[�^k���WYź(r�h��y���ַ"6Z���+=�������xS����p0[��%K1��Wy�s%#�5��+(���eP�A��q
��ni\�bw��9Jy���x��{��ޓ�S`�}�N�V:y^�D���w��V�z� i���#���W�wK�q��G@Xк�`_�A�r�!*AI�s-���&'���2�]��n/���dG5Ӝ�H�z�������U\@�>�,^$��w{(�ѣ�e�%E�9�oH�n�ՠ��^���xw$��=K/r�]�o�)�����y���{[�M��;��8z�Hm&�o-J^�2��AJ*�ڻ}fbYGg]��[Tky�$^ҫ�h�]P�X\�mTwX�̣̎I+ao�i��I��d�h�b��_'��>�yV�J5�X4�O�:��l�WH���0�vP;t�Pr���i䔙}�����Oz/%��)`�\�7b�K�@j�=��.���꼳��K=w�EJ�A�DA��9�Z����!(!	�w��Q��@P��T"#CU�>�Q���Q4��%8��Y�J�'��첶6o;��ўQĸ�_��_���;5��kH�\+��2�-՘zG+���yE#P6Hz/;(u
9�Mŉ�+�u�s�l�\�2��XČ�$�p�t$e��5V��p����"r������c�ga��m�A� ��L^��w�fD�B�]�۾�2]RO8ޝ.�]9iބ��`.M�Ί'�i�՜Mnf)h8� ��vv��Hܺ��)7�;Y�NC�"_Ri�$��P�6�م)���J�˽�RM3NN$h��J��!�ڌ��G+9)ج�8��t�L*��]O(:��b�{%��r��i�ʻ�z��4:F2{�g��5�y<�y�B�g�R쑗�X���1cv���x���y�������f�ʑW�2�a��pQ�6D,��2�K����ù��rq�-�3�����]�8�ˈw_oEv:1�U�:"��M�݇���\�'w�[�J74ve]��J�}i��.MW����ۛ
��Ğ�4Ӫ��~ĭ���=��%6TVf�F�������x~���<=�};C�O~��T��h�q�$���땽:����9���1Ⲭ�&#+ih�r�܀;X;��.� h��ՔgZ��b��.��8��
�u�"*���m������Z�s�+m������k����ۏs������Z��ugl5ڱ,�-j�ѳ"�tZ���k��^��³�x{	�oFN�`]�e�f�1^�o�H���fQ���3pX�����!н���݊��g%O��Ga�Y�c����TA�^%����盔#�r(/�4������7���g]����x�	�F��$���
=M4�����n�`˕���o���|�^C"m���y��³�k%�j:���|T[��J��8sGYad����q����\c�E���:�n��İ�f�zk��rg����: �}KrU��9C��B����v�v8a-f��nm��TU;A0�IV����1�b�j�R��lmf�OJ�����ʩ�"��ޤ8�s^���1]��H���^��S���U�Te�X |2���q�bt���Dv<1�|}76�x;��{���&���m�gVpC_G5K|��E��r
7�$I�N��86����Qk�͇�n���++(3s��^3y!�p��=帻�w����KX
�^�:��ذ��{؇�߳k��,�X���9�s�Q���mj��o� s���;S
�9O+y�%"Q��lS�⽲'a�ү	&�6�(��c��� 9isĖ�2�'v��U�yxϟ�Ih��w���{��}�6k9�T&�m�����S�;:l�bQ�.�ZjfKŃ�0��"��5&���Ec�9=��+M�#�2�fK�V���edˬ��MÑt�Nw4n\=�}��;�nr�qE�\SP8�OrD4����Yʈ'�v����$��)�N�g��7�x�������y)խ�~k�-�}��y�y��r�F�|�L�+�J��p--�׷5z��W�M��Ȥ���N��|���7"��8oVr���V	]����F.�^w�߽�>)̒�yg��� v��碟ڜ�(c��w]����t1�B`ɞ��p�Uv6�!�{��Q��Xq��}�:�lZ�Eap�j���S��z�m�ӆ�H&����s�{6�$�<ˤo�`�qL�^K��\ϴ.��A�=C��S���"�{%n)Y�2�*"�7�v�����M���mi���K.^:V;q鄖֍����<�-(�mY>�H,*{wCV��&b���l��kaD���V	{o��I�l�0/�bZ��w�� 4am�=���o�!]~�E�Z��v���6q�Cgذ&W`2"��8�V���q2�o�T(�*�0�'�ews�f���!�X�m֊3Rw'E�+e7rm�[��&k��A!_�O=��/m8�[;rE�;���4JX]q��l{����Ը�F;�uW^G|��V�Z��jƆ�1Eׯu�{�a+�Ma�V<��O��M�P;��X`�`ɗq�� <w
�|`�����KN�v14i.;%Ǎ��h�5_{{�4��W�&s}i���(��o2�Z�����́kӝ���;�9$��M
z�O�n����N/��Ѭ�Ѻ�S9�@����Ond1ۭ�oZ��5��m�k`Qh����}2�,�8e.�*��2�����C{|u
�l�Ә�{�����i,��֥`�m��\�9�tbEC�s��*�}F;��.�m���g���{N,/��U�ye�2�`��O\ ����$G_k�)�'��+��a��1[�a;z�ۙFH�Lg5�; �/����1�t���X�Gr�L�R��j�6z� )�rf U�A�k��P�2�D�X3�O�e-q�&�1\�L��ڴ����Ȅ)©��~�Tvi�EC5e	`v����R�s9�{��ї��.��T�!�&1+(�3 �О@��f�i�w�a�I�Xm�7
�p]�y��)FCk�ņ�$E-��,���{��+v=�T�����;"l<c�V�ǚr�;1�4BS�v��#�Tz����+��5�;�'q\�l����ZOv|c�36؅�9cu��qW��T� s�Ӟ<��U��Y���Z�c��A��:��ݝڮ��y��-�N6n���ޑ�?K9l:N�@I-ɴ�'3�%g'_U�������@��raN��Wzw������Ә���{0��L_^DӒ�e?��guǇ��&V��nĬ�6���dvq�/lj7���4��X̐4\M=-,�p��Ռ��r�gɷc��:d8�(���R�Ӆ����
�� A|>Ű�;�ma����`�ΣP��V�O���"\����r�/@��S7�>���i���W.���ŬoJ2��s�M�\��%gEƩ<��W��fUէ�u�Ȱ�E����<jTSZI��7�Ct4�N��ěm�L��
��>��m �#���s�=]���轍s�GG`��b���6˻0i�1���WE(���ùi�s���c:`��A�����w�{��l��i�"����U�
�c������Ly$Boqs��x	ǸS9�j5�1*��2���	�%���.�-3xy�\��b)�U��Q�X/v�0�U�g�`�l虙ӤaQ�­]5.� )�(L�;I�		t�2�Z��Q���m�R���KT���/1Kʻ���-ku�X��F��4aVe�D�ݸr�<qo��k l*�ث�m��=��2�a���S�*�L�%�fլ�UK���\M{�H�����ѭ�}0뮡1���'#���Ws�g#�Ɍ��;�A�S����%P���F�M���}�fS�s����w3d.6v�܄ezA�	^��a��n,�9Ɓ���#���G�\1�9���	;�t�r���OUth'����#��u��	�	 ��}���^v8)�9$�{�J��lFU���Z����=I�V��3�UӬ�X�Ru(��	��B�|T>/i�I/�\Xa�Reノ�|2��9+��༶������n]����=O%�3�=�����Þk^����w]�Jˆʑ�<wb����Yخ捤M�.�H��
�Q������k��%�2k�ZH=.�QnĚR��ݧ-��Iƭ�
��H���"���%o��[�x� &���h`S�]F����F�����v@l����l�	o��Y�5oI���8�}��Z�ڙ�Z�5yZ��+����O=���dP�����}��'+<�)�`�`�`�A��f���.��vh9�.�B�]gK��V�F�/�<R�t��͚�!Cך�5�[
{k ��W�/yƴ6��U���0�ado��LW�Z�2���G���.P^��'�sc
O > �_x�8�H깩>T��@��|��еn�6�����\3��W+�l��EV�ܘr��p�J+(D��i��Tt�uۭ;ZY8Sj3����.��q�P2��v]0f�nlh�Ƹ'��`a&���mT����V�u#u��n����,X�6.��:/" F-�K�������+sX��N��\@t����y��;�K��] 8��=�y�eb���Cq2�s;�_;P����Ӽ��X<�R���}�}<P8v�7�ejz� ���*�J�c=��H�ϥ=�!��fɗOu{��x}U�' u�C9&:��ܮ�uv�N�:�ˣ8,���A|�ݠ��� J�x��=a.j"�
vub4����(#��}�,���fsˮ����f_Oy5�Q�F��;�0h��R�M��M�y�N1����nEW�u��hU�rz��{�AX��Gzh]#R�k+�dfT��W�O��<&���^b�4��-��)@�3,+=6t\����:�&3Vz�l���/�t[���G�c|p�Xr��Tҩ\��[�N����!�X�6�܃gk�N`�����I���7[|.E|�*EKDfЫjvR���^���Qf�:��Q����k�k�壈�A�fr�.�Q�1`=ҞM)K�[�F�LdUb��n��<�en!�Żû%�%3��ڻ,��|e�|6����#T4��j���K<g8D�[Ov�,y�m�M<N+w�U�(��h�0;�G��t�S���1U���!A����b����֓�wiǻ{�A3���97�(Sj�v�L�sD�r|��X��}��C�u);fuh��1�{2��Zr���J�W����d�7^�;��|6_C;��wO0ו{76|��D�ۅ8���&{�L�x���!�քE�bdp�NY��oJ�m-ZH�����s�TRj�u�w{Ѥ�k��c^F�٬r�<jXx*rq]e>��B�6�3�hܖ��|��=�+�\ �t�߻��R
���p���AM5��f	�&s�!$wm�V�wv��c�zeݶv_���!�&�ZPf��x!�-��RJ����&pT���j¢v�5�����%dO�`מ�s��<�Q=w�=��_��}���aG{N �61,�Ӌ"�J�u��=u{O�0���R7%��6�`n��b��Kpan��b���l\�ȝu��t/q�vQ����V6'1�M+�ҼO�q�(����v������Sr���|
KK��מ�!��2ɂ�U���3�@���ц�ܶ�p�E��m:׽�\��f�����-��Pb�v��p�n���Cŷ鏢^\����<��E��;�3���n���U`��pkx0h�Q�A�m^h�JpU	;��)uh ��`v�i���ޗ���� �բ��^�l��s���G�g���ڵk1�񃡕��\V���6����(7i�N�� �c�Ԇ��U��Wtڄ�����ՆQ���	ݩAʷ���x�;U�n8=3h�ʗ�X�.�þe���%�1_�� �(�,�p�c�=y�4�H�i��L�>�ʆX6d����X�1��̗�N�x䆮��M=�SR�eS=�:�JM��'aƵ {C6.���/@O�j�,n*���Hs�[�����p+[
o{8�GF<a"ڋ]:<�cɒ��d��`����0I�/��q�CWڵ�[�P|z�U��J�&�ib�	d%S��Vu�z���H�ў�ԒWy	't�]I˒�ֱ�;.+�F���T���%����\�e[)Ҭ}0XV�(����T'2�����݋��w)����"�s̽i�д��+p;\]m���G�]�A��5X�]��9T5�u:]󴰛ɍ����}9n��8�s �}�qo\IE�� ���:�qhZ���o��iH]VY�~'WQo��g�n݁�#`l�+�a �[N{,/�5��=۞�|�3�Ye-�Ooys��X�@
��zc��1�сa8��H��RI*�X_z=ȏ����&OT��<�~��e2Q����}��S�
�n��E�#���J�I{RC7(�k��ܱn�djp����`f3�7	�=;��;x�*�]#�z{�}���1��-Ns�v8�Ŵk,��E�I3�-��y����*no����~���-Z�&zmÙь��[����17�5p*r�p�J~���fh 
�}�J
��Y(b�	t�L�G�O���7�C�}�Bb*,���̅��3�K�b�wvX�
���4�.�Og�W���xF�}k?_Cϻd��:q���`���N�m�P����$�X��ڜ#.��������Q�f\꺽W�t6�C�Sl�t���s��N��5�]�u�X׽�ۮ��ֺ,^U�,����1�@ʼ7c0x��Po�B�5�]~�?��Π��⮑�|=jG��h���x�צ�x�,�"w3!	�V�Ӂ�L��FfL ���`�򔽫���ӫ[ָ4a�^Z;#�PV�i�pՅʓ�d�[��[��x�.�8蛙3�Ξ�%D����n1�w�z��\v"4�����-�!F�w���=�ju�=J
Vi:L�m*�ʍ7�.u�L�I"�584%Pm�����w;-M��&	3u��S,��(CW-��@�e8:�iW\����#2��`����`d��	Z��l��JښJok_,���Ŵ������W��-�T`�j�"x鵸~+5v�߈�!�[n�@�J�ƅ+V��3�S�LE�e�<։X�7yȅdٝ/�5��Q��9r�����a�3{C�RΘ&]��QJ�q��C��W�t+NO�B��p��t4L��!Q�[PuM7ݰ���b���A���N+�a�l��t1�,N+�noR}�(�]�U�gg3u���b<tU��i��Cq��'�G�d�� �(��M2φ�7"�y1+!�%>.�P�𦦆JsF����V4�ܛYֆ1Ӆ�h1���sؚ۲%�����L�}�}A����p���Dnr�0ˇdH��-_'4T˓�g&�Ѩ��_����6qU���8o����[VnQ�MS]#L]�Lrɥ�꒙��H�QˎmY-�&�贎�{�P[Ub��#�&�d���7xʭ7n�[�z��Yґ�[���4w�p��d��v6~k��\�����o � �}��i�]�$+G�{rwb���B/w�\�V�N�ԯp〗6�AD�+���9��c�!#����O�b��,d'���~ u��5�a�zaؒ�P�z@��i\>�;#��E����l�������c]�sB6��b2�s돂/��-mAZ7@������<�ݷ�B�6s�K͇ 9�=��e�	7�;"�"^�h@{
L��W���71\�Sf�t�]��	�SN��f���k��qkիe��q��=�
�Y/2Ăf!W��� {����{ۇ���mƨ��cm���!NvVW(������qjE=&��+�ɮ�-��L��:[�_6鹂'A�M�Ŗ�G��InԾ�U(��54�Kw8�3xפ\�M��zĥгw�c�L�]q'885aڒ�4�%�ɵdMf`���ñɞ�I������j�f��&cwn���X�\�0��-a��w���[�b(�v��i9��Ù�����w���m�K���­������]Ω1X����N��}E����jɂ��K���в���8q�+�qZ4C����_40��M���z��e�,P����:s��h�3Ε⟮'؞�W.��C��\:nGwoC�=�I��ڋǞ0���C|��N���gz���i;�_u'kl�:�i������� �U↶�*A��Om����{��c�J�A/�$=�:���f�����I�P�[(i���Ut�pjy����M�A<7�m�"7�ZC8.�@D_�h�a#�����8�l����K�6.�$�}��=_fÝ�h8'�t�(�M��b1�h�6�>�������L�Tx�
�α�vz�z=�l��J�v<���`�Ղ�R����KuP��e!��$(S���r�=++n���M���ד���s��1���5�^�@����c�#՝�g�ܬ^�B�������Pu2+E�<�
Qu$��*�w<���Q!ʻ�NHb�J!�����*YX�y�Q2a���e���M:dUar���*
��	Va�U�h��%�s�S��՞�2��Ua�����tV9�Ot9�T櫑;\�#*Ðf*4s')9����i,��P�.�:�Ep�H�E�e!{��4�AL ��%ii%��㇂�AZ�X!e�ygL�C�k�E\�s�'0���V�-B�urwin;��B�Y��h���R	��a��74�b��Ԭ�U�/3���j&�A�+t�ڨTeVRH���*CN�+*Q3��QD���Hr"ԋ�u�!*��`H^�]�q�����2���2N�=Ђ��u23"4i:��I����
H�D#����H��W��a��[�$�Y%��W�5;�73h��͊�����;��s7Pe ��Κu8fU��t�;l<��ʊ�=�m"���6��F	�:0�i`��{�L�o���F~Sį��j�yM1���HEf����Nzr��:} �P�Y|�����4!Q�>�OP?-#�����zPW^W7J�S�� ,z�鍃��N���K�t�9�i��Ӻ����4�6�9 ���NW���`ǒ�ǻS=]ټ�U��??M���0�|5�ָ׷�0�^�.*�{P��G�jB�4�G^�D�����3v��?8�������C�P�_Φ�]蓙�q	�n��@��*��zϊ��3�Z01	�O*��T���0&"Ӵ̌V��-�6w!]}�n΄����;{ZO{co�6C�G������:!W�,T���P	gv>�-���yLB�_lZX{Chi%�{#sQ�l�K䕤s�'��c��XYFs&�l{|�����ff���������;�c�Зg#��H<ZRWoI`�څ��^�]2���K.ܤ�J~8Ω�I��u�]�����}�[G�Ի��o�IX�'�KI~8�9¯��1P��*x|P���c����
�;\W�g�*C�g�+�o��N���mݭ9
v���f���Y��*�e0E5{���XZw&�� �Yz�*��2U��g_G
��Q��F�5���ۘ�5�2+�fb��W,�սׄ�g$��u�R4�Rn�:�ޯ���=v��r4��Ke9�!T
���n��^83�W79V�~�6�1�o���:�����}�>��oN��']��7pt�g���[xe�W��s�`I��� ��c!d!��k�����V�An�?1A�M����;llU,�G����т�u@?y��A[>���)�J�b�Z5�Ó��l���6i��{�5@��m0��!`)�&x�>V.xhy���O۔���FNV=�n�5]��W�����)d�&��n	ή�����X̭"�x�؇���Ve�FX�5Ϣ܌��5j�з���kU�RO§����9U?c}������UYʎ��r6|r���=�[��R�&��ȴ���ǧ����>Ύ�{�pTu�?_eY���@�n���G:6��8������6+Uk� %�}H��h�:��u������꫎���C�)R��O}�'Ŝ�>� �T2��.��x<�d6���h�%���3[,w$)r�ʚ����o�:4�"�I����S��2YG :
����.-c��ho�eQ����'Ⱥ1�a`�;���prO�sx��&T�῏t�2�\�w��"M����m��-�q�̖%�;I��Á]�fv��e펻0�$dM��r��ۋ�M�2�3����>�vc�m�B-K�Hoi��|ω�~ו^�����.��4�������N�%�J��~y0���cG^Σ��qG����o�Xz)�
#�Tf&�,Gۨ��M���
�&��Bo��0xm9l��ۿ��V� �ϩIj�&���bB��[:��*�t�;��}Jb��N��\9B�D;P��}�m���B8a�ȱ���F�[ʔ,$�<�Wt��a#j�t�p�q*X�#:��
�f���0�L+�����gX�3��'�m`�2֨>���%��bҒG2�"��V'�r������x��UVԛ@ʜa���kUB�Z`n�	D�9� �Hc�R�����D��k�;�dח��m����><�����=A�X�TTQ[�Nxs��[�����L�����F���;R�3A3����r��X/��<Lo>�E3!\�%ƹ&�ƶ�@�)�I��1]�/N�)�v*'���	�w8�/N�2s¤�G4�Ѷ�#Z�6]�'�'��P��òe2�b��2u	�ؕM�][�F��\㫰p�����k�H߫:͠�s3Of�j�W��%�t�	c4\D���c[x����Z!7��Cv7�4�Vl��٫V#�X��ʘ��F���2�OJ%�*Z���w�N�#4��C�ty2�>^��P{�������W!i;��L�X��j���`���E"����� �p��׉/@|�Ťu�d�)��c:#����ʺ�^c��7F��J���,xA:a��*Nr�+�1=���,�&���4�g�����[��C���x�<���gLS�M���|U! ����و��T7�%�8��6.�U�S�9���H�W~����VY��N��O�ͨt�F3��R�P~�QU�t��`�hNn���*�I`%����yqT:c�eyF!w;�@�%R��>*Yޥ4a��t�w(S�0S�E��xFN���.�,�.�����~�_��|+�aIͣzY��v�}3C�p�	@����|�F���FG80}�UP�_qn�>��:kg��7e1�����W�t��8w�C>�~e�)ڮ�qE���
T��M P�����Y��U	1O��zqt����`�K1{�֒α�@�7Vȭ�7�asǸN��%�(��)F;:��4���;T#��eU�D��-u��
Ӌ��{)�X����{e]�z_U�W|��м�<��JΥ.�\f���YY51&q.�6`��a0�%_ci�R�D���Z2�!)�R�N������<>���y%�R��2�n�ĸ�ѼB0�aL��۲1���ke��X��a�ǌ���e���c���ӆ�87�c���)�f �)[F�0��Drf��\���e�p[���Y�؏��~��ͳHͩk�)a�|~�����e�"�+���&!R� ���(p��w��qv�����-���!Y֢%�!����}���3��T�y�r��T�(d�Kj��q/��������d=7�EJz����Z�I�[Jy_{�N�~����/����\ޭ�$	T�4�B�� ��1�X�ѕ:��m���r����7U�e+�6��{��-��|Vs'�>���Z�n�!�q2��x����f�mC����8�4��窎��Qm�f��_�f�2��V��Y�`�`�� �R��:��\n6�y��g�{K��$�>X6�T�����u�~4��u:�buc�:��c��'7c�jD�3ܷ7T�j8&,�Fr��j��� ��ŧi��;�_Ω�����.l\�#����rX����Ӵ�A�%P9{���~�;$Rk9|S�4t�$*�Fu�,utx��-�	¥<ۣ��l��˭$��:���-���\:��Q"��$فW�-Pgg�R(�(	�V�Fn�\fl�l���_q
�`lNA�����]
]���z�ڑ+�+�g�Y�j ��.�}a�C�����L��F��ìj����V��/�Pٞ��IZ�5�ѕ_W�SJ��AF����X��a��ܕ�Em���qt�#T��Gr�ѱ��;9�*Rt���zK�쁳���ۈN�̷O'�W��.D�	.�5+|r9�e����[�/�iW�uw~��悤�o��N�[[fP:�֦qM�Ơ�x`�z�#�9�Y4�����65��#f�'v00M�R�s������=DIKjq<#�:[W��{(n']��u�#Dҷ���\�7W�{
O�8�¨����:�7�1��)�]�����S��ܹc-��	Q��z�(���x�$@f; �4vH�[N���G���֌�5jr�o=�p����.�L��ѥm�ě2t�:޴���/0
;�ϰM.�9]�ۓ�ߚNh��T/y)F����o��Ď��̚7�:�\��!%#Վ<��:';��>S���Mt"c9Eܘܺ,&yX}M�VOm�gr[�	�{r����w�B��졭j5�i�e5F\��=-�Γ��\�ģW��3^�n�u����M�ljR$���uoq^�m��cP)��r��oi�q����|�(
6����Qf=�g$>��]i�дꫨ[�N�|~rv��8�e��8g�]��{�+�ݫ�Y����n|�n10��0�௫�i1q�(;���t�Ӫ��pTo��Ʃ�f�>�M!'�::�z�S�'�'1���9��T= !���u�n:�.�u�뙋̵�#�A�ĕ��ڝ�[?[��W��ݳ0��j�=�	)���!�&-4�F �]�ux8o��]�����<������h�uEg`����_[L��t�t�4[��y �Is���*�k�M%)����aY|cu�p�5&�ũ$���n$H��ｸu�8���!�0�UaꟗF�L`2��'-��C��v�|U<0�ߑ��?uNŧQ�����H4F�s�%�XkTZv�����MT=��?!������gS�hu�J�,�J���&\�E��$o�t�p�Qb�;�����}�	����9��[bS׵-b���Kv-)(�-���sս���B��j�؜Typx��qI��ƥuLKmL2�c9T۳t��3V��u�<f�7�Ʉ��Z�a��
u`�R��Vk�A�:ث��tC�Mq�qGZ��|��6�{׏�3C�Μ�_���!�:�_�Q1ؓ52݃(��;ֵ�;λ����9�>���%\8��0WΩ	�2T� #W��	5X4�F<�^|���V�EU��y�ܬ��[\�f�6QyX�n��͈(�W�R��`<"��X�*xs��-�tq�G1��H<�\f��)�ag�s�K��b��k�m� i�31�\�k��,��*����a
,����BoZ�{��O�ᆆv�(Y�����%��M,�5yÌY��.���kp��:���!!�@�>u�֦����U��_�;��L�r�'����ܑ5V�.+sא�uv�P����k��c�Awk˕J�����G@5��:�!��*�8�^\9����b���o�J��,_L2#�PT�� +� 8��T��"�b�\���:�R 9���*�Á2w\�s���Aˏe���],1A�8Ueޚ��J�K�5��Zj�A\N�"�u *�e�-�OE�*�Z]y
v{�k2[�j�Ib�oS�:<��y���u[g�A�A)͙`+�P�Tr��ԶuA�1�p�8QaXc׼M{V3S�f���۹�:&�܊�!����y�A�%�藗E���d]�
<G�\~��pC�����Fչz��K��V`��]a1ǅ�w
|6��̺`9��I�*�e�*)�e^^S{ҙW������9��-tK���%df��w�qӊO��~�d@�,D��dN��h%]|������� V�^�5�]Ot�bƅ�!-��@�l/w&�F�1�T�l=ْ6���6hv4��Y�g"��C�ukT$
N��I�����\Y&hϨ_��{�; ��(M��|���t�a��4FZ�*�{��ސ�n9a�Wd#z߶�P�F2Oc�����E��P���c;6殭�8ԁZ��wt�!�9�W1�-W��"����k`���dK��{�ʱX[X��26����0!�j1up�N�1�ޔ�f,F���9n������9���r ���#w����w�&KJhu9�3���_��u��Ֆp��J�k��Πl�+wh�ӳ��-�[�^R��͕�+w��T�!��Ϛ�K08��㴂�*X-�Ē�5@$���	TL@X��v��z��r�k
F���I=�1�Y��{=���3��[�j��w�健�-���/���>ZE��G�t#�8z	���si�Z��G��xoq"����m�rׇ��T�rL�z��Ґ��|r�d�4N��[W<D���#��C�%� �H'�j��˶%fnPYN:�Y�����I:�0�؜��zw�qۗ<=����NsF:��.`�}o�Ӕ���R��p�=�w��1���؅q���ϗ:Ҝ��>�1-m7RG�����9��n`�=Y�M�g�wVl'�\���{����^B_On������6
6� �]�tχ{����ꭽ���na{�Vq+�YL]v����#}ۊ���o��+���Ž`���T�4�f�(�`�a�B�EvU钤;0&-;L��V���g+T�U��2�"���~����Q�ys8}e��,%dm��i޲w7غd�}K�"uP��&+\�ݴy���+%5��+�\ܜ��2��Z���r+��s[!aej*{	=�C�%���L�.������׭e�lźTƚ����(t�>����{6ۤvFH�9zAĦ+��E�4&�r�Ǚ�/O�m[�,�EX6� 1�q���c�y�+Ȼ�S���h�x������P[<0_=v��F�������6�][M�@H����&/s9jP��'��E��ZF-��wb���-��ý�7!:�$G�|���ţHa�!��k Q�sH���.�)���{A�l�W;Q�z�#5�6`��ê�<F٢�U�B��7����q��]h�#<�ڑ�e��\��[�s�C>�˽B���炙i.�Ct����Q���j�^Đ|���=���w�p�WݰҴ=��Ű����@fR���p�]�]m`UyKzV��k��6�W���<Z���IJ.��n�<���(�h;7)�wj�mܽ�JA0K<���r��ò�t��x�5��FJ�\���'(j9�2]/�������I�oDjf�1�cB�Z1���d�_A���}�	s�K�e;3w��=�A=\l�A0l�nْh����d�N���
\�vƨf�##�rWG��S�ө��}oW���iٻ �me���!޸�s�P�P��d���5����{�/x�z7�h��p��)J}Laq��v��Z�1m[��Bv�9]X�
'�v��V�&�[��3 y��s-�a����m��GRV �����Z1j�ͺc6�xY�KV�]l��0n��]��b�ዙJ���f�V)�,vC���x��vݱ?y�&����K���u*kO۹ƕ�hm�"�٨d���7}��E��b �-Y"z&�αɄ:&���}˘=��K���7� �u9��������,aϲ�A��p��aOZ��k}*G�H����`U��}g	�t´lu}[������>�zb�vr/n�ŃDOe�r���V\����>w�
�]޾����y����k�*�,�w���2-?
e롽퀿�Ո�l��DK�ry;���Dk�Z���ޡ�6�2����[�~�u���8��wN{�{J�(����1ʆ]�7�UbX7׶eAd��"{���������m�ׇ�OHƽY�X�f$E���1�3Kj��܊���f��TKC&��[����e=�/S4���w5��%�Љ[��x:U�|�3�)�q��8�6U�z�*_&�;*l3L�����>0��,^@y�oq��fV�$V��8Z�w�3���o�^�Z;R���]�_�=�vx<��Z�Pr��t��-r:��{�r��aR��}8y�e�҉wR��Wo�l!d�閉���u}�^�k��,�4I���ɒw�Wns�T�Ș�8��$�(`N7�u�K��l���t��[��v޼4��s�$o����s�}��ԩ���i6�K�u����7�|3}z<b:���ʻ5Z�$��&�mM�w�\�LA�nQ�E6B��7�s���w�34Lv�6�&����?�T",�y��W�,�J���n�׸�+]v�fi�g	�/r�	�=H���c�q�6]Ԫ�x�,�$#����U����pd�-̀�Ww[��Ƹeo+�=���nSG{���J�+1C��"@�߃6��_=����;�b,�<��#��&�Z�
�O��j�,�#�� �+wh�h�����JJ�R2B��D��	2���UK��9.���t9^�B�D�eZ:9���#R�	<�Y�&;�wi��9%Q!!)K"��BL�2+"!ݚz���u]�<#�p��t0�M�t�0�
���QF��뗜�s֨!g���Qd�"V.륫�y+���Q�(��r�4/7*̥D�5��P�0��B�q1.�W�Z��0�K�V���H�����S�N�沅2�ԕ�sW#]2�Z�Z�3���z��E%��zVfe��h��J)DUU�3�"u�1C"�w!���5T�JiR�.�0��9�s�F�Vb,��$IB�wr�n��,�wb䉻�98�EVs�=�D�]i���P�uqSWG
n�\\�;(���TT�w@��;�j����(��k�z-2�E#e�t	H��>AR$��Y!�]j�{�kK�B�|P�<�_a;pc2�y�7�*T?:1{$	f����� �E�'S.U�}>�3�EPn�(-m�>{|���0��}Ns�L*����P���p�Q��_�j<>ݹ90��?[x�����\o
����_�0$��q��gT�}�@B"F���q��>� +^���U���*����xC��ۓ�7���M�	����}��Ǘ{v�z?A��OI���Xz7眻�%�7߰s�t{v�щ�=�	#�=$2=��g�GF$�Cs�>� ��> �v׹�!�W�iR\��^g��x@f�'��3�|;��yw�k��3����k������zBI�P�����z��x@����۝��S�s��xW��0� YR�;Z�f�3��m����O��ǵ�	!��_��� i�>��}��
���~��<������w�ߐ��˷??~�'��>?����o�ސ��:_6ܜ�����0����xO=>����گ�?��v�sjo>|��N�oO�6���۹\��������H
�������,�gK�$x�>��Q��G�?k~� �>"������1;�i��_�o)�lﾭ��z����� Fջ�3s��p�!;^��G�<&q�ǭG�w��<�G�o���'��~C��ۓ�{�?#�@G��VD�V��>���~���8E&|�����Ѿ���]����p)�p߫.��@��F�>��}��P��?jE�	"���13�!�F3��
�녟��ra�ǟ<yL��۷!뻃�N��u�������o�N��'���|�ߐ�����o�{��}E�c�V�����ku��8�,�g�o����.�oi�;ݏ����[�zO(xMz��w�9܇���q�0����O����®��	���wA�c~C������8�H�;���G�f\���W�`�X��4���=q�/�o�ɹ��x��뷴��>~�y@�����=;ý�N=>��V�����97�sɿ!^����Yg�Ѓ�"H�'�}���I�$|�V!��r6~ś7�NY��>� �}O�9��݃���o�i�����~[���}��ߏ���0�~v�Ǯ���L>�۽o�yW|v����xON�w���������9Rv�|B!}�O�?ko<4�ݸf��8�s��yoN�R��s�O׾�z�b�{F�v�,���i����v}/Y)�6uZ��2����P�e��NUۮ�}��0gs�x���`C-mk�Hֈ��r�����خ5�r��+MB[���rV�hë�W���YP�G�|>LL�{��xS�q��!�Y�>�������}��<;�����O�9?&�N}o���~O�9>���\~C�aC۽u�ˏhs���w�$���ۑ=�9����L���6 ;ۭx>�������q�n�e���<��xv��M�ڧ*=�#�z@�`>D@������?
}M�7�}L(|v��>Ƿm������R�Qֺb����G�}��@dx>(<�&�BC��7~��rs�8�x@���ǋ���M���z�������|/�� �����?}ϴ�Ȁ!.�vߝ;Ӵ�g�ݿ�����7��� �{/n��8~����O�iG�Y�>��bw&�y��.��S���='��C�y(?'�O?\��__���ݹ9Z�4��o��.~�<	��yH��G��DxC��n�6�/�q' �����Q{�I��y�?QF�{�ϰ�g|đ� #��d:��xAB��	��bw�}�ǋn~���:v��^r�b���aBO�`����Āg�F�G�z��ջ�ˏ���/.9��;��Nh��'�DG�s<!�0����7�돨s���ݼA&_��ۿ���?�˿���_w�oI��:O�;�bM���<'�n{�o�s'��2 �şg���}�G��|u^r�M߶s�)�!�
>���pG��!�0�,X?�>>d
ǰ!����>��;����M�	7�$�@w��P���|�x@���?�Q�=����a��!H7���>?'Eq���f��^���@�<+C�o�����{��:w�i�/]��W����5{̏q��G�g} L!���#�>��|$�dx#~c���Q�fH������Ei�������V~�Q���/�6�?#�<G���2@s���~��W����Vﱽ!ɇϏ���U��ӻ���🝿�w����"=�p����Dx=�hw}�R��>�G�����G�n
C~����M+���g�>��$��d|=��Q�L/�|�������o�����NL.��{/{C��S��y�>@g�����@"<O�i���#�>�nc�}�#���)5O�mO�f���QlX)�r�w���C��ܺ�z���R�����h�>�]��b�:�Cz-"���u� mȘ��r����t�:��ѝ�cU�rd�x�{v��r��B{� 1I=�]���O�8x� ��[�W[������}������r����~�w�i�o>w�9�����yO<8�ǣ�M�99�k�F'|C�=���S����������>��/�I��#�@U�~�;.�����lb�xT!� 2>ݨ��Q q�XQ�����z�w�I����=��J^�ۏI����oi�8v�N����<&������o�������A1��>.�FOx�Qy^�
>��	��|8�|��ȿ<`$�Ă@��q���$����O�����ܝ������w�����=&O����{C�<�?�ӷ+���'� ��!�z�>����>0 �%�ʪ�Ξ���i>$ �$�G��~�'��q��G�o���xC���ÿ;To����˿;J���ɾ������;�`	>����#O������'�FC��� i��_J4%�q�p~[j�G�߾{yw���=��]��I��}O��?$�N<�w�{v�ߐ�E�����ݾ��'o�}���~�]��@��{��<�\.������'����$��|Ǡ�|G�2�eg��G�ua�^��+�l!�����|��>!��H�~�!��.��s�G��$$������!������ԝ���.<��H����n��O/zc�� "<+��{�G�}�|�ݣ����LLSO��eg׵�;� ��|�������A~���^U�����q���N���z|8�|Nv����99�?]�	�]�S������ǟ~�]����{:X�<	��{�n��]M���#�D���˝�Q��I#�����M��G�nW8��< I'�o�_c۷�܄�;��)�\
o�F|�rw�ǝ;U���xOa���ڐ`��|}�I��n������]�s�x7s>�#�h}'���jG�>�8�2/���=�Q������ 2 _ �ߓO��w���<PI��z�����;ӿ!�-�ۓxO�cü;]Nǵx!{K�ay_о�Tj��~Q5S7��c�$	>g�Dy��L|�ߏ}�}O��>���/���|C _k�C�aDw�� |@��G����0��q��� #�=���$x����	"O��d/��<:Y%����H��ٔ&�&b��:��h�/ge7��;�>�u���Ƕ ڟ�^���gO�e����F�Z��xD��X/Z}Lځ-�&P��-�&���k�Y�c��y��j�'4"���#0�+t�t�n@3����U#�6F�S���v�p�"e���H?}]V]e�7�ÿo(xL+�S�r�x��}v����~y���oΝ����7�ߐ�[_�v�p)�;��}�7�/��/���.9�S�~��.���s�~����T�£k|�O�/|�} ��@�9��{C�a�o'�o��n}���<&|�c�>F�C��x�=�_�xC�O�����y�}'՚�� �z�}�G�}�G� "~��AI��Q��i��vze/�����,�����_�;�[{~�מS�;T}C��˹�T=|�ɾ��h.�1;�{q��q�7�yL.��Ǆ�����͎S��6| ��b��<�Dx���7pi���堫��]�7�>����������nM�/���;_i���xM�	'oo~���=��ޝ�<��O8\.����~NNq�8�W��{NIhY�C�i(|}$ a�ֳ���y%\|x\�����~�G�"8}#���o�< ��}9o�@�<��ߐGO���~�'�G�H�61�
BL+��O�zO)��&������<;�o��@�����x:���7�/����j}T*��qn��73�=���}ğ H��1E�� +Cژ���,�3�!�{���g�G(�I��� �>#�^߾��'�~#���v='����o^����������1��)�E�#zj|:�I���{����/{I>!��������rl��C$�EC`q>�!��X��q��^􌿣��<	���_D@�ϗ.��+������9���v<��}�i��Z��x��d`�w�\ �#�C#���F"���n�1��b�We^���P���i����	�Ŕ���<�8�&Z�'��ߒ��{��sBB�|�>�nz�Ga���.�>���A�v.F��X���4�y��G��ч�Ө�.a��/RV���dߵnW�k-��s�\��K�}�	�����3�H+�m\O�j/[��b<-&�׃X����U�u�r���j�2���GZ62U�89%�aP��ϸx��r��9���'��ܪ�\n]��@L>a�a/f)ׂPg�����q������G�N�:K�R���n��qT�ƈggEt��'�c��b�IR�`bҒ��ڼ�>K�e��me��A=��t}��!�N`3P4&�+|s��_��V�� %��<Z�{Yli��D<[��z	��,%���;+�zu���_��Vd��z�#��F����>ĕȢ���ہ��w]���1��ƔTDI�<��#�;�N�h�m\C��2�ꖄ�|�Iɭ{)w�6B� �^`jS�݂� ��!H�cX�+r�B4d�\l(����i����O�PD���zz���2
��+h���Hɔ�V0�!4%��
�k�}cwL�j�R\&�y� h��0�����Q?H'y@��K��!��Υ�Z��"c8��t�7���ک���M��]�{�mS@T�!�#y`�J�s���uЇ'����mώ���^\,�wh�|�~rjܠv�u�QZ��8rdR�ͽ1����	��� (�:��ش�����3'��gGe
�ۂ���h�C�=q��/Jǀ9��<�oZ3�)ɍ�u="k�Π�b�K������3L�p�F�4�r5��;$>�����&�C)��rU�4uL�f�<�p�_����8���Q��W���%Z�g$��V��$�gO����QQ%�����W�V0�w����g���0s��Vq*�	��UHklv��P�v�δ ��C�ԭ��R�^��=A�s��<Xom!�Jߘ��fg�w!1��.���vR[�g��c�aڨ3����� ���#�ܔ�~������2]�n��Z��̌�k������b�&:Z���/�����n6e`�ɨjS/���¸]�]�@��6�1�$+L:���颲o[����ep�T��s�L-s����s���9l��ۿ���i��7�4��Ǿ�]�%��*�G��bX�2ZF���d�(�kV� ��<}>���,v;�[�`}7�+�罢�^���^�`�c$��X+3�21���WP]�7�$X��@uv5U�����J��ll��a��`����R����6-�N��;F߱�Ux��C� �JH�g��N�w�)�V�>b�:�&��SQ� ��}E*�P�j�w�l=F�7\s���z�O�Ʊ�9:H�lCd;�����؃0�I\lԨ��ҭ;ԇs[���j�/|m�{Un=�	H���]c���1B'S(�kZ�y���@hy���ReȞ�k�[Cd�1�Ny/U>ƽ���R'�f�Ê�����l\\,���h�r=�#(�U��������$n��Cw9r1�5�����0�{�󫫺4���b�v>�g~���R7���K�d�F�iL�!v�1]��7���6��2�ɱ5�\��Dj�CE��7�HwxT��i٣q�F��S����<��9(�M�ْj�\a�pf�N4�c����/MlK�j��F��5ꩉ:�7b�/�%�޽|JQ�O�t�*=K�!�eݯ@|��1��_�9��C��������L~�n�;}�e>2U��7��u)r�A-�k7����ݽxk��
)\��i�F���i�9����L��e9��Q��]�f�(1�J��㤧�>4i��o�N*�휩�d�4�lE��|���N
�����X~tb�䃯�
p�|{�8��s(e	����YѐiPjt�Zj��R�`�;��d����u��]v'�.�sNm�Ҥ�Q�0���l]|�B$� ꐏ`sC��_ �9B$n�a�Cwe��okT6l��R�`N�ܨz��n�����yd\�ds�7���	���֬�(��yO���O<�aט��,us�yN;Z�"�Y]�	�ʼx���(���:1���P�9flɨe<�x�èv��\��,ɀ���n(��L`��}K!b�e�޻P�4+��o(*gE	����0/�e��x��ϼ�<j9[�u��`���j������ sq[?Y���4g�/�T�vA�|XYY|F_�0)��*8u���E�xr#��co ��>�6�Wʠ'��騒�q*z��"ƷK^�v��!��U��)5q$��z�c���d���k���[(�K.'��h�����4�p��ݏ+5i�������c	�)�X��A��mH����@6�y-��F+2L�SB��m��Y��φN��tu��]�՛��~�DKix��oY�[���;��X��[��x>����p[�^R��j�W��A�ꐇW�-�ޱm���lY��N�T��u�%C,j}`'0�éU��vԮ��"�\!ƞ�`p���ylS�4�Y�ɗ;�6��=3tE�ܰ4��CC��OT��0��YW5������N
�J/8r�8�x��*s)^���2�c����fr�T�TiY3��&܁��	��L��t��7ޫ���D��3���7�����^B�?{_�~ݠ�즹u6�8�J��!�%�]���ʽDɜ3ϋ5b��%��^��ՅI���̔�%�gH��MH���Z�XƱ�lה��.�#��r����Y��g��՝��Zi�������Ωx��W�=�m�+)9NwU�	h�z�Gk��{
I����G����ﾯ@�+��I���6�����L;��-����z�0�S�b�GI)D��e�����mi[nz��(�3��U�deKʺ�	d�+C9߭1^�ʥ<��_/5�L�U��=��GÇ���z�!4+\�q����$����ɝR��e��#��+���<T70|��H�Y)��r�r}x�:�<��j��_��Ek�G�)I��v�7/[�������j�GON�ˈ�pً�J�܉��� �1<P$��j]�r���2u�Ꙅ%��	����r|sG޴|����3z|��̔kS==+6\d�X�#9e#��*�g"�����]�v9�����=�WzŽ)L	sW�[�����0�(9�]D-$i<�‧�bs�}-���d%��]��}|�>*y33�T����+R���u1����A�� ��F������b��������s��-�C>-�'�("w��hÄ!�W�Tm�t+�#&�U�1�k�;.�ƽv�b�P���6���qlu���9r�-�Gb��7^��Nǆ��\�M=����lc�B�J@_���e�ם$����nler��M�K��f�*�l�y-zn�埱��\�m���>�V����zBQ�VԠiD��q���������m�k�x�z5_�kFc5*�&�u���f�̝4K��kN=�R���+V)[5������E���ν��6��y�����U"�d�&�n@��8�I������4��=�s�U���u�\�oh�1����^����~����O%:�O�M[�����:Tw-�\j���b��V�t��v��;$�Ga�F#6-!7���١���t� �GfJ�G��܊��=U<~�?S*͞�8��Du}E}�`2����<8�����^�T-ui�J�L��g!:�c���	,�(��Y/ 	�8_�}��U�=�+���AF,��Ӯ�k��$hb�]L�!ܗ/NS��"|2]�n��]i�F�rg���KT(.6��?7�����Ҙ���̰�0�ߚ��퇗�y���R�Vp��W�I ]}^[i������=71H��)���ϴ�`��g�9l��v����JZ'�B���*�})V,�K�Bl�$�`�V�u�9�E�S�L}�k�Hg��4�G�-�ŏ�l��OiItɏL�+xm)�7���6_4�i�
����2�^ɳ��ryOM�F����[XP��ݭ���qa��)�A4���8'/��һ��R�e���@]�a��:*Y��5����(�M��껁"��u2��# \vKb�>�q*��Yǘ�Ti�E���9��\���[��>��r�O�|p��t�MtВ��]�<ǱLB���5�R��/����\|^��2��ݫFi�S&�pF��1Pͻ0b�)Ru!OJ����n�ub����/��Píc��Ѥ����v���WC�]��+U�e ��<����gv�uy�]���T�Y�oT�
�?ly�$��%aܳ�B�Zެ��o��Wm�гG�e�w���+��[��t��0�@cZL3l��w�w>_nh�p$đ��ˠo� �X�
<m�+6�-q�(gf.�m
/v�	8��ֲ�X{�ӗTR���F2���}3�tP786�.�ub%#n*f��m�ȷR�V/�<��2�g㋷f�ԏv;�W�U*����|k�J��"m�壧g�S�"���V�덃J���s���\�,�Z4��o�3�+A�4��w۔*]��2�D��c�͢t*��7)�>
�BF�ܹu��ʟs�(_��ohr�	_X�͋lB �ޢ�W���Sws�6� A�����ڛ�b̔#<袵�Av�D§!�9)	�we]N�V�(�+D��/S��,v�9�n�g!�)��Ϯ��������74�5v*u�إ@s�*}�G���~y���+���c�����e�g9C7U4;t:��
��a)f�'!dafj'�P�ʏ	��T"��}>�.<'����qw,�]�8Yv��$N�N^�.�⳺�8�9M���h^�אҋ#1,�:��nu�wzͻ�&�68����̳�����+����TNfKuj����}�a�����̛B�샢^ag�}C�.���17�$�#oV��l�}�d�Zz�s��~ӡqޒ�Ȯ�7�eA��s��[�Ρwԝ1m��Uv��H�w��`L��0^9��ޭC!�%h�0�@��%��շ!ԩ�oEkh�Le�j�'�.���A���?gȫe�k ⺙P�bQ���^I-\��3��Sܼm��*y&};i�"3u��Þ��TS���?yM���z�r����=�6)�D��K��Y�����+�WY��Ύ����q�ʺ����[��0�k^uY�V���B*�R�Cq�e�Ƴ\ON<T�h����^��|���@�"�_P��K#��V�]�E< .�vI�*NF]>��*A���3m,�eY�nCV5m���vd����J���y�*7J(l��=(�r������5|Ѭ�y�i�3j���_{/������ޭ޿��������=hQJ$�f4��)"4�Os�F�j%�vb��f.��
P�*�,�"���H��t��#�V���r,؁Ib�TY�3f�kWv�����Jȳ$9�� �EY�f��H�6�"���&j�R˪��wv{B(���Q!�D�"�ť�K��"�V���(�������xT�����TP�Q�BJ��dI��H�S�M�\Itr��
���)Q3	*�
ZDs:���4SL���A�0Q"����eJ��B�J*�B���C�	��h�,���ZPcS	C%�K(�iBٙt,���+@4��5B���F:���G0�U-K22Ҵ�+��%fJRX���Z�(K�x�e�Ԍ�J�)��%(�]E�H�y7-WD�����k����"�0�,��TU�Z(������0�V�QY�YJg(�D�6%@j���3�i�>?�w��\st�o=��lX"��Y"���6k�u\Kox��X�����tc�[�S*�a&�E�������C� ���W�_ty�j.�7vD��3Q��V]3��Y��,�͙��U����XY:U��j͛���K���f�s"�U��©F���2֨>�1��nť �����������{ךsP=�U�ܷq�˺|u9Ѥ�s e8�.���"N���悛��qD�@7\�3�O�����J�>Lmtc~ߜt���6C��vw�_�lA�S$�=n��t
��M̌�|�҅���0��ߞ�aZUo'����>�j{)�1p\�%�#X)�Jŷjg;���}���@�`&��F1Řue� ^=�7��,-�~�ޕ �}�h+eE������ݦ#���ҁ�R���WJ� Q��c�MyY�q{3�*�ǫ1�[-�O͎���/B����SXO7��)a��������7�^\�V�Χ֗Cf�D��X�v�u=�ck'�9�#���(,A8/�u)���)Wp5�����X3e*zwYSWW�����[7���@!�N~h��u.?e��"���������)����;�W���sK^�t�.7Zq��^�2�7��_u�f��(d�sxs"x������+��`7���$���}���r�m!.f�n��l������ �9a���iHA��Ơ�]I����+k�\�ɽ�������ｘc�{�CV���/Q--S<�G�D�j��*�e��
��К?2��ر�kr���*�qy�Ԡ�{y�T���[�E�l�4����[|Nޚ�#�L�T;��uH�N�eE��21ms��]=Oz
��lp�]y����:P��Ib*uPEf�V}���hН�U��r0(��7I��]���9��ʇ�@�	׷�	�i����t=*O���be��OI��AѸ���p����x����	��b���Q%T�|aX���ᇖ�=�����Q�����n(�?QJ��!���@-7�>�nv#� �K#��=��Y�B���#	O�-V=�ƹ��X�B*4���M�Ԛ���e��p\���#j۲2�sH����]�g.��v��3��q�C,�"�:�W�e2�`Cx�.����c �ґϋ��/ ��S�S*U�-p��v��kku����[Y���N��y,;/��Q��B��k:Aے�W;�|�9��G�3^�L�X~y��� ����T��Aȼ�=^����V�d�=<�����md�2���'\���\�ȕ/P'�g]��������(:+9}b�H��+(�Y�雼�4���޻�odKT-��3�<d���c��5�B4Ŗ�w���S��{��syI�����Ͷ�h��
	�k?ʯ���6 �L����f��9p���W�>&�?A;�",�U�)�����d�셞���^v{jI����B+[�a�5E@�@B�����$��^/��,�����.��QJ'9̧��L�lh�&�RA�{[zF�-Ne��v1�}45��d�5e-��c4���=�ݲ(�<���K�a9ZjFLv%��y<F�L��_���'�h1M_�OkT����f�t=�dAP�$* is�
�,�GNnu *7�c>uNሾVt�*�����5�i"QO�uc���~~gmTv�����K�<���J���yh�(ͭ9X��Y���{��3��3$�Q�B��l��sB�.�O�XJ��\[P�K�P�D�Zk:�p_����d�����w,Gb�}��߱��|N@߅l5S�ou�����v�u|�U0��A�_bWp���� h�^;��[�LnM֎����<�;�馡Ajږ��y��0;j:㮩�bQ��6dK�\���rИ�[5Jj���x�Iᱯ�B��G�tc�EZF�U�nv�B�w5\Uq��裒ѧd���i�Z��{fE��J7V��l/ 5������5 ��E�jor��0AJ�9�m��f�6jc��f?}X:ws�{G�� �U���}=�}Ҟ�qW�������������D�I��S������A��PǙ��)�V���|h�x`���0��E�r���W#8k�OU�w�>>��1�lx�Z�'2�E���y���S�+�*�T-,Nض]�Z]S;��L�Hh1�<>�W�w!���z9��~P��:Y5���{i��Q�O�ۂ0W6� ܢa@b�*wE�#��8���}���Af�M�;q��}�NX�WEù�z���Q��Ja���p/!�`�%U)3Q҉�;���F��Xy-1��wڣ`Y�\���W*L4r��J�q���pڨ�K'�4m�@s�{v3�Ǉ���)�ؖ�Љ.1�\�+>�������
�ځ{55�y()�{��`"��c�/ܰ�5�E��j�����XvS�d���%�*�<8*+�i1q�(;١������@KO�Yp��;�P�t��~�V(ǳ�)�+�	���ChD@�R�e)�<�o��U��}m���T�i�8��u����p�N�Ew�(�������z����x\�ن森M@!���u8����Z*2x,)���~�=��o���H�y���\���t�V�Q��r�6�uf�l}َ�����fn�(SX��e��_A,���-�쾫��76����WF>�{�R�x�U��O�F�����|�I����"�J�-D�'�;���{e��~��9�FB�bm�A�K�\9§����R�Y�Q�
���������J�ȭp��aY|cv�{N�6w� u�4�3�o�C���}:�A���x����t0�YH]oG�Dit��0Xo�岾��Ni��5Yw}L�z+g�]����1\f��rA�	� �m���-j�� ����̳~)�绶�/1����{Z��w�v��痠ax�%����
��ٕ́ _8�D�+ġ���ơ^�E�bAӂ���SF5�g9�p8j*�ZW��yBM@i��f��cgކ��a�aW�c}Q=-�p��ߓ���0MG�#K�5��	'PiLN�Di����S%zNU���9�`����}�>��ܜ�T8!���`7�&�@f��d����>+��[I{d��c��U Cg�\uJ�tt�oO\����8C\�%�_M�&v�fk3m�P�I��q�x�j�c8c��,�3�-	�{joz��<0������9��f%}�`Rp�7�O�js_`]^�膬����M�ó��=�F��*i�s"R	!��PR9��X,TfV���&a���Q#g�f�����'�t�#����@�:�GX�.��Ny3�Hů*%�*��w%�m���� 3O�G�O'��h���T��Eh����>U �1_J�8�鼃�f8�x֫Ȼ�0SCyU�w�%�t`)�nX	a�魘eRԺ��7$����RÝ��mt�K�J~�����"�����Ω�Z�3Z��,,A���Q��,s:="_g`�sv/�D���U�*sYf��)s�Ɗ=z��z<ѾwPr��^��Lp�{S$�N|_j�6i��1^P5C��f2tm�G�E��B��Y9��j��{.��ǎ��J����}�	��X�>��	b�ſdq*��շ��ځ�f���=`�f����L6ܙ}�OP�
HԊ�(�T��u�zf<S��4�����h�W<���/Y��+�~zL� ��LE�r��u���1P�*Q�5wK(}<,<�i׾ɭ�h+V5�������r�CϑN�>����}֥ó��� ũ-��-�]��b���M.ӽLg��YY��t^��
T��!��ra��F8U_(Og-7�}�F�dn+Ô:����K��k�اV@���CnlOe+w���p�y۳�/�t��|L1D�;$"=��+��*%qb}�T{7:�b���c�ݡP����:0��^��I�sЃ5BOK�����[�]�{)q�E>c�#qm%����9"�������Đ�#��Q`���`)�_i�ʼUcx�&�9o�b<���̑p'�Q��p{x'9���U�Nج��(�4#�!�"�{���S(|�iX��vJvٌ&��kp�O6�Kł�����
(B͘6��3"���s��6�mgc�>��n��ǥv/S9�iƩ�-���t�fA��Y�+�"5-�r�퍀�cԬ$3��A.O]��du���
����λJ8����!�>����d�X�}`Jpu+�S;j|��;�P��1�|\��B.M�q+�Cgv������ϛUtn2�r����b���zY<�P���Ր�D�ܻB;�ੱ�^�ڳ�H9��~]������å9l}��.����NM�Z����G+NQ��R��C�J���7�j���3L_��s+6�H�q�kȹx��:ac�AF���EK�}|��n�z���\�F� ]v��+"����#���v�]{縼W���+{���j�@	�,�ť�8�ֲx�'t��U,I.�N`��:.j���o)�#����ó���s!]��%�P��-�5��]l��-�ɱ+}����m*vr�"��2�Ib�P�;nL��3�j�t�HJ]�%�E�:B&��k;gA\2��G��h�R棧V����,�M�۫�J~��������F�N�N�=�/�S��^'�|�سl�g4/��z�πWR�9��-a��SD�4{2�!5�中T��*�}al�P��s��Tq>}x�Q�2��Z��GP�db�3/v�w;p���z2����Q�J�qt���4C/�f�c:&�Gֶ*p�%f���lOn�ƔR&��%�����oP㑬Pr��B�o�G9�9~cUCg������)�����W
Q��5�X6
5�A��X8�-=�魈�O��g��Xj��9�����p�gLry�͏I�k$S��cH��0֬���F�D���}s�f7����bN�zRG��I_�졸�wx���qY�a�����:�;q��sH��]��X��޽w`�� ��H���u(���g��8Ar �n�j�4�'�Je�6r�딏V}	_�V�j6Ҩrju��%�0t0	UJL��O3�
,��:��'aU-榬��#9@Z��\Q���Y�m`�s������Mm�ɍu.6Me8�^���F�OQF�ﲷ��u�8�nq5;�WD�KjQ袍���m�'kh�!�X���� �fqq��4���c�����\�ʲ.`���4Ȏ�sI�6;���^ü�*=�ի5Bk�I-�7�UÉ�����M�U}^��o$n�ټ�,�BRZ��fW~>�p��c�j��یv��G'���>�rS�n�6k^q�*y�ك��z�4��E���H�	�e���;u*1�͋&7J=��K���:%���C��s�S�n
�|~�4ʳ}嘃����T���Z��Cg"'a�so���ݔ�tj
%| �Sr2Σ8�s1̳T��o�	�fG��WrIV����v�v��z<
������3R�Vft0��K��L׶X�JG�����la2]�n��uƎ5ui]<#뵝�	�D�]G\u��3�!���ȖY<�e��e�߰���%룙8�bѢ�G9j�rI
K�@-�ۆ���	�N~]]0n�ea9}cOkg:�����'��~DV��]2c��wW�k�'��u͜�Q�FƣȄ�pK�,��<hs����Lf;I����^�`�,b�BzK+3�21��:�{z�-o	�־^�G Թ�Y�|h�K�CE�4��¥k�0BX��ò�K���e�x�|�Z‫薧�b�=��r�8#����W�<B�.�>j�[���=F�`�&�ĩsи�K}������6�q�9[��jPX�(�į.������al��i	����혭���)��*b���<]��"�iKCO��F�����9����ь�VO�s+2��Tb}q7����������	���S�(Cb6C�d7��_(�c��)�n4��`O�Ʊq��9:H�8!��^V��T�3�X潽_>��ˡ����rx* �����F�����W.�E3!���.h�6{95�J�V	��s2#P6�M���Ȣ�,ѝYh^-��^������dJ,#'��γP�0�u�4S1�T^�FI����.�T���s����<sp`"4F���z�IH@�̪�C���Z,2�`�l}?b��� ��eFj�!��/X��5�����Q}�:lύE>9���A�O��j<9]��")jU$s؇Q�)���]ﯬ��!��R�[t�b3�3�]L/�T��u�G�L߿e�;��S�+�`�}F�4�To��`᫸B�D��:9�� t7*��=y�	�Yjk,VBg���I�����E;}00�ՙ-����i>Cm�jt�Q���1n��;V�r����4��Gٟ[٨�*�vi}l�+b�[O2���Xέ�8��k��|�˦D�ק�4ni�8�h�N�R�6F�v^A'.�⭛����w�
w�a��b÷L�0���8��ʳ+p��\mw=�X�Әl�H<�lT�]����3��#Fb;�D�Q|kG'	�#+������>�����k�u��~f�C���6���؛�<�ޱG�V�͖�;Qy��-��I���3� 1g������S8վu;(9�2,���U���/v���w�;6���F�Uk�\C�tVkL��8�bA���&�X�]�NU�#���S�uۙ�ɕ�nkU�z�l�xd;$/�sf)d�[�n�g����W3s7P����&�r���\�ͷ|��$L2o�Y��y��	�q�*�|�+�H.���-A���3':D��?@z�DK�&�wЉ����B�F�h)wv�ܥX���IV��$��腎F�U������úX��%��a�l�^���z�F���&�)��:���s���V따u�t.��P,F*��F�D���\�ň�*�4�H�c���V�v�����=�7A��g����L��Œ���Q�Z�b�
lF%ê��̡���^Fy��b0����u��Η�.���{'g`���s	���X:YQ�º�[���@Ӭr�UEۑ��64V,79��s���&U�:�Ÿi�}Y�gD�u)�6>�d�0G]�J��(�G�j��TO�	��y�섖��j*�9����NxYrc�닉�ÓT��VJyXf�2��G(n�Ϧ���R�V�و��F.�s�z6er��$�ޱ�R
rƻ��tON�M�U-�"����ȌuǨ�+����a�v�'J��#��O�o?"�]����B��!��!]�#����1�h��6���z�lI�/m,O�E�z�����N�FK8��}��<6k�ۧz흫�k1��}p��eH��-�ts[�Ǜ�v��ʓ�Z5/�ٖ�l5�-��s�/�j��v�ق�M�D�
�������Yu.�0�nY�K<e7��G�b͒�̑���Xᖲ��uk�n�~&	�����a�n
����޿�����وP�ۮ�������m�9�,^^Zj ���=�ϑ[��g��st03f��6�v�/S��(3X�&O0��Y�6a��Ӛ�]�Zf���⎦�4���-ɗD���K�7N�޲�N�U�z�˷�<YH�<��H|1y{����lh�wYV��ue��=
���!y��9���{Y*���w�瀘����pY3��]���X����wJ���LW
A�n	ľ8p�$WF3�i6��%��\y����KiWd9}�8@&t^�5VC6�H���Qмγ���],R�mq��#궈J�O��L�Ź���*j/HE���D��P��!W9s=�ʔIL�R-�ȕ(��w�+��"���F�wH�""���*(��P�%N�$E`�9y��/ZJ�)ad�g3-B��JR��K$.�UU)(�EU�!�GE��-IUP�΁�EF��VWRC��RHX�Q��3Z2��]�sLMd�T�eI�s4���jF*X�3��e�J�D��2�2ULй�����+� ��(�9L�+)�$�3:���A�TDdRXd.�+I�օcL���%�#$�2��,���ʒ�Y[�XJ��aEs������#D��Pr�IP��[TBZG"죝#J��H���Es�a��q	2H���+EE04H�"障%B�C	@��Nm��R*")�H8S�@����X�w�B�9Lb��QϖC��#�:YS	�9�)�0(wt�����1�����"�cGR��~��""J'�=隣`����YAF!w>جB)*�4��	�N�. T�"�uPEP]ؐ��G����|�Hڱ�8�|��L�vT�Z��b�ި �V���ylo�+��t��{K�X���̭�>�-]�\�	�cMW2v�oO�ԇ�K{��3[�Rfy-5��gd����|E{N{���w�O�)v\s��m�:i�}Dm�	�#���߹Wr��� H]�� a�1!"�1U��)��S,w�1�'��pX���Yz��������ӣ���q��E#8��E��ǌz��ZE7�nF����	�P{%�[��v�W���I�,����ߝS2)L���Oʆ�s顝j���XgT��]����4C�}��q�8���ڲ�$'R�/¶6��R���J՞f��أ�o���q��\�}���֭�2{!� ��亁���W�zI�a#
'j K�R]a��HJ�v�x�7�Ϊ2����G�sƀ�ؘR2ܰ4�[V!��@�2�oz�UC:aS�JF%g.�6U��9[{�RT�ԅʼA�e>:��G;t����X���,䨠�[,��S�d�k�W=J��{$̲���;��yI[*�CI�k�^SK0�Ú������Zv<x�e�(����T�q��qS&�������z��wle�`��|�&޻�b-�.�`f�f�A���?m߶b����.͞��v3��J�s֜�_���P�u.З��}#�k���O�o�fW����|P�p/\q��7��=<�Z^�+m�)]K� �y�4������%~d�pR�A/��i�W�j��L�B�N���X�Ȏ��G�~g4*���#*_��-�eh�S< ���~J��^�]�l�&-�L�Ȋy}k���>lB��sB���zX��(ta�6"������ob��]�j#6�K��tal�P�Ss��r�+�Е�U��qalnI���{&�q#x�����г�j�[�#p��Z�ae����1��v��n��v�t�v�vc������zK �@�Ɉ�e)��|4&�+|s�r|Z��1lRQё%��Myw����W���hE\`�� 08�2��G�UZ�E7_��Z���ka�qi��Ӣ��wr{U��md��W!�m�kT`D�@]���H�����t�]4�<�d��JFI;[|7T��Le+Js	ыH�j|����������b]u���,Nv����A���6�Wv����m�m��H�e��ɮ���կ�E�l��	t�/����� 6^�Ͳk4��*ub���xx�Uλ;���n�!�"[W��{(js�OcwH\�@jS��N�V��0�_A��'9��Ao	����]�[�Bݚ���-�&,1aPۭۨ��ݔr�|&̸�d�>\=A����@�H~b�֍F�%P��ɺ�^|�0�`�Ņk�4�:W#�[٧n�|1�@|�c�[qF$c9\,Ŷ�z�����gc����>�K���>W؁M�%�I�칓�����X�->�Z�^ǋm�ái�W�	�2�<T��S����;ۯ���ҫ������>�	�e���u��W�u㘀�v����mj��T^-J��Bq�C�T�!s��9F��ieY��gۀ7�3�U�*>�k����)��u�o���qxY:;x� +����|�S���BFs�v���OL321�Wf�$NE��(�ٕ���K�����Th����D ��܇�ɸs�-�O�]ѦqX6�
y<�X��S;<���&KJ��wu��3�!��2�'�%�����{M�Pb�r�vƆ���Ӧ�ݷ7����[)c1�鮳Mr�S�䌗[O;���սu��ՇV�udC#���7��3�T�v@.u�����\�+b��j�z�\5j��q��Y޽�F����.KSn�w���O6��R���۫��3�5E�������F�����)
߲�6�3<�@�=>-����b@��)�oW���`�x��S��N�]����	�/�S+��DN���$�W���>�9ۺi4�V{���闊,�|>�P��,v�M\>�6������Y=%��9�@,M�ѵ��i�iQ�;A��[��6�����MF�eJ�����-��,/��[�{�n��[��`ć�@������0+{$9�F]1خ��q)�Q�T��
?v�֛����s+��� ����Z���P'�⻧���#��l����1՛AK�Mՙ���B��؂�%q�S�n	�^<"��WiU[��P`Wo�3�r��$wy�&�4Jp�-옑�D�`?�ڙ������r(�C�5�:�ЛǶ�*�]^�r�%��k9�e�=��4 f�J�܀��l	v�Q01jY߮ +���#��F{ ��^{,�J��4��6�]�����Z,3_7,j8��z��d�}�ssr�,����V�����h���3�͞�r��5�F ⊡<(L�$w8����m�.Cz� b����ug|��s�m=��\��d���2*�*�KsyI��o�swؖ�o6��iM�11ʳ8���x+%��;^K�Ν��c�x�L;��z��DF�(W+�����+%��9�1��f�%�KE뺑��7�ќ[X�5}��XL�َ鬶�E�3�g�ݾ� ��L�'_4n9�A����|NR�
k{��|Ǣ;f�X6c	vG��U�zs�����MT53��K�ofe��E�����),����7��C�9�f�^��߲=q*�z�k�[|N�n8�:����7`���IPء��|X8�=��.�lV!��P�; '�`��2/pz��r��l�+ �My͙z�ꇪ��.��HE�-��u��}s�R�F�����cۺ	�ё��lZ�S�lgm���Ӛ>[)]�\�	�C/ ��;�鸚�O�곚S�jL�� o�g�/��5���%C�|G��PR��>�!�یt�c�#t��Y*c�4��һ�]>��� �jJB�b+L$V)��{�M\M̱�C0�a8�_�#�l�
c�5�V$K:��摔H"/��<\�D�_
�)�>C)���G�Ϳ�b˘ފ~Y4v�5�� �u7��؎���6�;]B��x�w���;̲�-����eif����-ЩnÕ�W�R�P��7i�����$TQӨ�5f��@�u��[q�Čo.��ާ�W��B�8��pF�M=>s��&n�����x��+�Φ�3n�Ǡ���ϋ�����z#�05������_���#X���̤]m��9N��ܯ|v��Ϯ���\��	ԶG(�cc`8ǩ\x�3����a(\�..h�+u:0�A�1/U0��j�1@}S�DsT�x�/��[��j�C�u�E����*;<<mn'�B���HԺSݾ�M��7
nXZɡTb�c9C.t�襸>�<`{j�����wڐ5�#-F0(�ɱq����\�J_+���D���쉉/z5����i̿p�1��Ņ/NI������b�f=�i�PʱQ3��ˮ'9�X�zI��6��P�����J�D��T�g��qUYg�82q�N��c�Ck7�J��|y �-yc�wF:�G����wNr��kH&f�cKv-'���1݇_"��Y[X�K��@!a��i�fC���֫���\G���Mf0n���}N��Ru]T��צ��8D��0�����������y)����1
��\��j�b��S�gΙ���*�K6��N�5�hn��dȨ+iS�s�}�7���4��OT*�����>���fCc�;��J�Rg���M��,��K��Sn�]�ݽQ�SU(uI��^ծ��)J���(�%��r���x	���������Лw���C�e�������~?V��`5{r�ȮDqt�ƈa]���U!WWjX���\>�Jy5�.�'7\�d��`��(	���_]R0�R���	�J���]Q:�Ǽ9-��� ��c�Z��d(ղRV,�$�6q�'6����V�/	ƍ�~�\���vh�!3��I��4��qx��Z�z���T���@]"s#ˡi0k��!%`��*��[���Y�=tC��2[W��{(n��J��*X��5�	;�r�T7���n`ҳL��3ޜ�����g)�YTj��\��T��-�&.5�n�x�%��J�b�S�f����kSS�1�?Z5�RA{.�}�)�J�b��Q��C�_&�y� h���bJ؋))�'3�)�� :��,�~�Bf�?0��H�3�f=�>��H���Ⱦ�6L̬Y�G�8���4y�m۝�1�JI��j�T���'c����yB�j�]�2M�T0.`mS��Vgr�m��c!��������_iXe�����!S�^S�Ey�j ���C	-��*�1���[7Н�VV����KsVu��.�:We;�l����A���Z�6�di�0
������7�r�Xy�m���F�Eu�t㫳Z��k��l���vR����B��G��"�v�"� �^��F�7Pj�����������]��C�n�;i�<l�졹����<nD�1�P�YԪ��c�Q�|��ɵ�Eu��fRB�_*Qأs�~��R4�e{�{���޵@�,~�o����TOemĖ¼.&-4ͪM���-�k�o(S�y�C����x^�T��;9_V��]�;մ�k��hk��+�o{ݫ���>dWVu�i	��=��I˛�P#���ʽ���<�A��oF�Tl�E�_K$�R�n�������M��ѽr��r�i6��ݛ"����ȁ��M�uK�c���\�Q�i���ˌp�4�5B�O0:~+�ڀ����\%n-.�΢�g���Rޚ)<��x�?���ן�VnWPy��y�m=�K�Dd�������z����ž������A��ɑZ$��T
{����B�T��*�`H�~B?w\Ok�Q�P�[�2^Σ|h@ݪ ��X�ݖ �ꣻ«rĔ���嗊���F�.��ȕ�Hif��ю��B�f+���@���㜡r�4�G,�;qu�\�F��J��]1�^�fvr$ެy�l<�V3g(2��M�:�,�RaAZ�;�Y|��V�M�矪������sz�*���P�D.��h�)��u.���>7n��#��A1*��.�:f�p����R���6b�P:�sSk��*��_;T��}B�&�w8��U'�5�Pۍj�]<��;pN�5TJ'.�0�cǱV1sS�d٥n�;��O5Q��{�zyfU5dLb{^�i�������#���%_J̯��z�#��}�X����Þ��c]�q��4�b�[���z^G>Z��[�ؾu1ћ}q�eGju�\�/���"�N��[Ğ�mmhO��������������ώO��ӽ�U��&���A$G��xpߖ���I���>#��̢�`��u��T���΅v�)��7�kF>9���l\:omWn��b�2��EW��D��v�f�����7��fV򉬹s�5�R�a�j�6��?"
�h����8ȿdQ�%x��=�n��Ϸ՝�E�s��-\d,	#ۅC�U���q*����i���y�g��/���+r�Z��?6j��%J\�`
��dZ��f�����6oi���-X����0j�-J�����(#��>ޜM_�磌�xq-l3�'�:���뮰�R�qż�zˌp��Ol���V��C����5[��\�i%b��%�4Ryq���-���\\����oQ�ֵp���1Awϲ
�&/JK�wҟ��wttnzA|�+;�hu���O>S�wS�=w�9Fa���,�Z*#Jk2��n�*s��x�t�w��aޥ�a��5�'��@/v�s��w��n��8���G>㕮%Q��r桭	�hE�x*�`�z�w�=ĵ�7�=C�-������7��}�_7�5�0�q��
�9#��I�ne�=
�u56-��A\����N%�q���S�pڧ\5ǻ�_b��
�]X�d���^W��"��� �[��e�K�8��F��ܫ������y��:)'�7�0����12�'ci\�W�9���b6�#V��_V<)���Y"�����m��cW˫��y{sN�j7���ќ�<((K�՜��]�"�g3WTo�f��3Yj�c��4��\�n���-c6��kHw1�(f�b9�l�؈�� D���c^��Ϝʷ8���u<�q;)����A�dı�G��tWs�Y���M2!���\��Wb�4�<�L�\q_0<�{���8Ӿ��*Aܱygq۔[q�z�[��C�n:/,$?{=Z������7�%�F�U��}����Oy�
�`�ŉr�n�_fێޢ��ޚ�ӈ5e0�67Mu�����v��![[��Nl�)��kE�Kt�XN
��홯n���,Bޜ�9ɓH�ww�-�u�ju#}i��|d��Yn�ZU�$o1w�����H:�(M$C{Եb�Ծ�7}Rw���� ԲŚ��nZ'6L�J������Y��
�tQ� �5�n5j8�搷�b�Kg)�w5C�3v�R�-"���fVV%��ɭ]`N�c�}o�&�pQ}K91x��²g723V+���w(�籛Sz�F�>KN�.f�Ɋ�L�h^|��d3����/�8/k���6�ε*�+��k|q�C��	.���'+���/
�۲)�A�Q�m^��`��Y=��w��/������sn�������l��<6.yoU�%��<S�ڦ�n�-j�T]��o*j u�ѝ��ЖOxA�<��fz�|��J��#\�(���G.ӎ����&x�S���
nG?E����u����[_TZ��Lz}FJ����W�	�Z�Y�Tdѳ/L>���y]'���L�'��k�sZ]."���:�Mw�����=�=��nMJ+�8��P�Nm�W�������#|r������;%ɑS��-�[P��Z����s �u Ï:�:�h4�\x��\R�hv��������r6D����g]n��Oz�����\S��V�����ӡ�zT9|�)V����q�Mk��w]u��<���C�����ˉ�U���!4Vj�~��О�r�nq�E��MYS�����[ն��zg���=&!�S��| w%0�6eܸ5
�u�/5������W
ܵ�%ν�ۼ?6��j�ڷ����[C�xqSp�Bln� wڭ�^toD�%guESzT�9�6�Y巸F��{h�V9!�z��g>�̔T�4w�:<� �:W���H�mF�5ǉ<PH��Qob���E +1�/z>�ޥ���<�urA����c�.?jK�%�P�V�Vv^�9�8��.fӃl�p.���5��
���:}d��Yjٙ�@�	���U���3�ޜ	H-!ɦ�{�M�;^uY�:�Z�]�Ҧs���mG7��&F�*EmC�a�6������~�Q tU���\5��Z��{'<�_wP���2�WD��f0�vŘ1�J�R��N��\�Vk�V�^�L
�=�HpD@�sܩ��_� �/0�f��U��4ʻ�Lj�������}���T|P�Θg.��*�FDlL*��#E��X�T�F��s�Q ��d�X�2K�(�Dʨ�4R9UQ�t�Q]�Z�QGT��vVt�Z$UQ��P��+,J���S��+0�S:Q#�0�Q�IF�U�2"(�B4M@5���Q2�!#�˅�D#EP��*LQAVg(��
�Q�T΄]k�g*����eZ��$֡$�%)��"�f�]�(�T}E�ug���N9�I��C�����9�$9t��S����ZW4��$�\�4�Z�Dz���E�Dh�u( �0*"�:Uz-[�➥ʤ�=�����D��h�"�(=��Α����t�#9HA\����QQ�E���Ȕ��躑T�H�8Tf-P�A��Ts3�Tg���Ar��WW9@U^s�#��yRTV`uwk�s�$��	�ۺ���	9����=w9Q�����q��t�Aҧ=�ͺ�|��Wr���������E�Q�y�`i��ՋH�oK�Y,e��D�fj�L"���ќ9e[Z��mE�`/��}��U�P��b���B�;�O3uT��G���2���m�=�m�Y���*1�gN;櫴.�a��L�Ü[��n�ۛ6��r�]Ÿ�V��!�UZo�]k���$�J��*{��H�n��r���x|O�ޯz��I��
����SS���tl<M�v��|��+�LmÊF�N�ŝ�B�Tq�06`� �j\��
�ĩ_�[�z�՝��sN;9�J׭P4�*��;�(w07
�-���A��/�m{-�_��Ǝ��;��o��?#�վ[pi*:{��T��I@�7չܣR:�N�5�o���]��6���S��PS�wL%et�Uym����r#� �\,׉���Aޭ�OtU�2��3�!==Dml�T�";�'s���8+�vW,�b�|�s��a��̖�=���<{=h�[[x�;Nـ��;�. ����U�Lw]���e�Hʴ-���U)�f/.u��n���q����c��t&
��X��v�\�t^�2_H�B㻻x�K�ܔ�6ﺊ���E���6Qǻ)��E�����}G�^�/C��gѧJ�8�e뚎��7ܞ�s~K��Co�+���m�[��6V$���I�܉�,�C`']nI�y[�kS�1X��6s�bH̉=�	��S.;�M�֮s]�<�O���v�{2�qk�b�ɻ����a�r��dֿ���Z��E�6���+7_F ��E�WLN�+v���t�܏蓫�w���ܬ�2��k�k5���.g����}��ZCŞ9+�&|���پ����e���
�Οk}z�����p��6Zu��|����
���}���*�X�Q	��\LZi�)����k'��uJؖ���zf�{�Gc�զio���ѥ��q�ՎO"j爽�_sޚ�k\B.�W�(���v�?g�X=�X�\#�Y��;�����@�Ӄs�_��,e��[���om�@l�P`>G� /�����^��@Na��O%'䴟:y.���5�����&W<��7R�k��.r=9,JV�����C�.�.�=��R�A�*�]An��mQ ^Y�(㛳���c[�H�Ȏ���G����3˃vz���A�Zܳo&�Ͼ��������1�{s���;R��S{k������Έ4�@�������D�,�C����뉇��f��W���oM�\}�羧�|�L�/M�����]F�9H�������9�<�B�����o�vV�Q�dHn��V'D�M`]�Y9f-�Ă��J��+�#�u����示�E��X'V�������9���u�ǵy&ڻ�x~{]n{RT5B�ě\ƥs�S����Bo�����媷�Z�{=�Z>�^��D[����5��i�ܶ����昚mƻ�Y�tD�!�֌ʪ���(;yJ&��`/|�s=[�O��O5�a�{�zyf8��u眆�+z��-3Ыu3����%fTO-}�w=ܛ{���p�<m^6r���ɾ�iW=i�p{����E������+E�&�r�ڙz˃y������+�rq� ƞ�1��o1�.��?T�9�4����������6.�����N�@<k�X�P<�0
�ok]@�8ڽ�દ%BﻧQ�DL�_{�6�	������gZ���A��wU�l�dQ�6s&D�D�يgm�ɝ�U��� �=��sĨ]�G:Q��{��}�fTs=��1�~�LJ����@7��l$l��԰mS�e����{vr��̨*�'����o��u�z5�X�S��P���u�1_G$ؿ�7�{3~W��r��Y�1|���%k��ә���94�J��P��+�a�j�6����Env��B0�R%���Ŷ�H/���V������+b8��CV�-M<wy��d���w%f�ơm�2a08/�-�Ib��"[�w��\���)��֋�	��\�X�N���JT(t�Ϧ
��S֮H�jg'�����B����u'~�����?��=�N3j-�����=�p`%�t����y��M^9zҮH���p[J�;Գ��|�P���JU��^ͺ܄���{�(�ez�:�ǅ.pu��Tr桾h&*2#1�k���xL�A�&�j�v�;}XG�,�'�n,��"��9�
�+M�«҉��^�1�	�w]x�tGK�N���sשF�U��'F5����x���t%��8gI|��`F3E�7AG��,���E�vᗁ� �*�/�s�q�lt���Z�#�z\<�R�b�������tU��2�v�m{�9�5����y=h�����a��q���vɚ��m���1��9n�W괍Ô"�5����[����MB�
^��Ɗ�Y�zp����I�T�vC]���Wd�ʜZ�7��k+�O�)�ܬ���q������O=s;�I+���^���؂?S��S��V/pq_gՑ���jOz�gSVWu+��PS[���Gje���*Y< +�^�Ha�p_�ӛ������Oҳ-�je61֮ns676m�ʎC3v��Cs���y�C�2XOj%�i
��Zi��Rl9o9Wn���q%��JΊ�UX�\��M#��n���uW�N��'T%z](��|�7��4�cV�����c_U�c/y.�6��0��KG8��R�u�[���$,��Q�I�z���+5d�5��}n�ۃ[�(t� 6~��|�jRyJ�X��j���C�Y�p�Xh0����8�Cݟ��*7wF�\�uʗ��׃������B�t��Z��_N�L���`����c�Wt	�J!����H��&�{Q^�;����t�Ͷ�ճ�j��w.2���i��h�����D�l�e�������w�I���^q�4�R���E�|�?��٧��|%
��6:ޕ.�'HnM�k�r�U��[�P[��vF�ͫle9J�1�w�
�љ��ݶ�c�墣K琳�=��t*�ƞ����Ye�;�T;n�z*o�4tS��p�[5K��Z��҆�'��r(�=V���7H�P�C�W�{�-����-�m/@���g�f����^��Kl]Vo\cg;ָ^H=A�Ԙ�6�[���B.������x�j����yx{�}�n9uJ�by��T�'��ka�ϧ�"&�ݰ��+dd�Pݪ�N7�k�Uj�uֵÚ������~�f��Aȵ�|"��̒��c~�ocj�K�ߖV;�r��k�k5�ܣ΍�v�:/����·��Cַ���م���V���&2�;�2����9�륕�g"�yK��[��	�$���	�<��1'\�2.��\/�,P�C�s�1l��q�a�l��/=�����7�;�И�yL ��nx�(Bڳs�
L���ջGO��p�7�CP��(�q+�@֐����$�]��������U����9?Rh#%�hE�_��gUIL+��m4���66�,��n�XX�o�R.Ӈ˻�k(��H<�*���u5�ꆯ�-��M}35���y�u5#h8�|�!�}r�v�u�Ȥ��V�s4xt��d��}��[�6�Ɛ���x�M��I���=QH���С�%���ޝ�c:�J�UG�JTj57���k1���c�MP���鍝O`�7˹ҋ\�wMƖ��*�[�PRy|��{�z|�8k���s��LM��:�[�C�σ�	h���Y�oV'�7����nZ�S��r��j��X3sS�aPY����D)��JC��B�}oV.9��0��f�F܁��±���,���6���<�I��t���]BR����zg6/�u*�SwJ�`	n4Q�����\wi���9��p���n%R'�܀s�@�R&60����h.*�:v��F�T��hub���W�n;��76:�+y޿P6��% �]z��>��k��v��i�d�e��P|�jS,�{����߰F��'l��J�ڄ�r��mEF���P"Dů�bJ�e���f�K�L�To� ���݂���=���Oj52�Ꚏi���k�V~�DO!�)�*	��;h㞞�̮+�U귭:�oj�V�[�N��X�M6�mDu��k�����ʹ�-C�;��{�3D�ʞZ�;��M��r�ָs�	Ĝ�I`�T����ȱ\�6V������e��+F\v��<��1QU0�Ybo�*���]=��W?���՝�is�]Ǳef"�V�}���J#�F]`�+����v.�)�:Ŷ����ts>�3*�o��i�6���h8����y+]�cc�l_Λ�=����/l�E ��l�@�9=���s�U=5��.����OY&�\�{�61��&����U4j8�(�e�I����s��R�qż�����Ik�Nb�s䷴f'�T
�o���I^*��{Ay�٩�7_�4�����Ge8T��j �]�����$K�D�s�C���-{�o(/#qg���F�>�+S���3\��b�{J7G�ըs%X���}�G��KS��,��X��C�̾���i���*��7\	^Ů5V?��ض �(���E;=�U���#���i	t�=o:��z;a���*;�|�0�JJ�1V�K]��,�q�Y�9�3Ғ#�L�p����ڋleD9Fa�����)hc0>覒�o1mX�1��N��].^�6�	�@w�`y��62��3��%(�}�o8%�ƮK��~�B�>�-�.���o��;�4�7�ä3q*����t��͆��u56-�J����SWO�w�_kE�}S\��7��:��w�^�}�pP�Ho������-���{W�kS�m��H��R50�Sa�4�/=7��+3���3�)x���y��������p輹L�o'��-y�
N@������u�������&�M��l^ʘ�i��@5[z����vs�_w0^sV�s�I�.����{m>k5���/&9ٺ�C2��1��X=x��~Ƃ��<�?f�v��������W[u�{�n�96��zȁ%e��M��&�V*�W�~*)��v�x��47���>�ѩ~��_V z��ϬW����gT�H�8v\2b�N�<F��B��u\<�]U�V<�h�I�55`�^��ٸ�g�GDҲ	�N"��֪Rn�'�ef�do�{���ۋ��I��\�v��vʆ�8ش�6�6.!�{j�vS��j�Y���V�*�E;9U��s�:�6�I�	`s�m�7�"yn���S�⦔H幗�ʍ�<�
m��U8�~Y��d�ȝATbT��;jd�(�2�NBZ�T7q�h痍���I��ޡC�9YBP�8�I�3���Ov��_�'��y�D`��%�4��\5��m}�h��Gw|�J��Č�x�R��zU!�E��5c�w���e�sƻ>���ʈr�@��� �:Oo)�V����l�k�Dd��%��4��>z���ni�Qw�<��zə�\vF���c~T�#�'�A��f�is�X�i����|�a������t�Zz'�ͳ�x��"�P)T@�J�5K�{�Q�f�pkI`��R�QUy�/u������-e��{qU��o��y��g������r^�����ך��n��$֙&�v���t[Z�J�g�ݬ���X<�!����5�,�t"��|���;\ƍeK�k��>�iI�9�v��ͤ0"�8 z�t�hX�odV��ٚ	�z�#S�\i�{P�P+i(s.vIۄ��N���Ӷ�Ö��z��#ux������6^D�2�;�HI�W���3�c[����ˡy	��^�^�Y��5
f��q�秗B�ϗ^�`p��H��V`AAhNӓ=�W�6'�NH¹�X���U�*T��n�屡i�&g�#���V�{oEr��{�����L�$�rg+zJ�]�bF��8sK�����@�8p|k�٪�Ń�ûz�G���ҩ�Ubo�Q$(��i�����G�̹�˷��U%�^L�u:�\�
o��rZ�'���$J�i�Wu�jJ��A�-�,cG/�]�_'�^����rR�68��..�\�8>�ΤV#�A�;k�L��h�bm-����I�A�mN�����c�4Y2q��f��m�X2����!h�!�� ��=�J�!"7�;.��@�z��C�3I	�|��~�Z�&��՗�'sz3fJ}�b�Qȱ���(��X {���B��b�<��٦�5.�t7^�Wz%��R+�(cT%#�{���'��ix*>2�ۨ�nݷ�O=$�fV��}sg'9�C����ڝi�/g#�9U�9h4<���,�3^v�O����WbX����B��`8UG�3(�Z^�-�e:=���{�����v�ܚޫ����.X�]{	7�V�KR^*=�Kg��CVl��y�xUh�,�l�X����j�6Fc�6��S�L����w�,m�7Y'3Uen\�mª+=ڔՏ;kkA]7`��5�Cs�{��Q�8��h�<�v�Ca���ܭڌƭx�}����܇�=x���W��7uqHY�k�#M�g�!�$V�oa�%�^*C+�)�)��[�9;�1���nJ�/hg�sSH�o�{�,�lHΨ��c��W12���56��j� ��]*(*(@�<VS��1֙X�i!�|�1�D444{ˈ�{/\z�ޫTn�uN�t�8��4�kF����}d�9�FM��{
�<;ZjHFL	��_KHlV�Ӑ��2��MN�L��N� ��w�!�|��v���ZW,5��`�%|_U�:8��-#{[�Q:����x���k���]u�Ӛ�L*,���U$�q��8Dz����)!��hy�<�/}�6����_�-��C�ކce�u%ɓ�̡��j�ނ�a˷�'L
����C_\I3%�qݔ�������+n����4>(WaH񝼀-�'(����.�	�B�h.W_0=[;i�����z�wH��͝2�!Fa`��Y��U�}�7����x�NU���B���,x������o|(y3�e�*�[Zo� �P`�h�]��U
�"��s��) ���J-�6E!��է9j�N+�!�,�r\+���Ԭ�:�L�Qsr�G<p�C�
��9FkN�
.J3J*Q*UUrԪ�-Y2�2$Z!�Uw=�J%TM@�@�ʓ��v��L��aT ���TVaF�Yj4�e˔�D[+T"�I˅Ҩ��WZ9BEJ�"�R��U���G��:lՕDQj��+��HIEs���tP�)I��#�O%ԮQEU
�C�Je�R*�i�WD2@�Y�s�Ӳ��p�:p�̄�wAqZa�-L�u�w\+�G�l�3QE��z��m	
�TE	���"����a�9�t
�ʢ슩B�D�4M�*ʎA�ΙDp��肻��v�(�Feu%d�B�QQT�J" ����PMP*"+XYU�L�9PB�#�c���Ei5�t�++��"���W9�R�5��l
��IΒ����d�B����6��
uO��ّ�x�W��}��v�~Sl��%���k��鹴����7�N�#��赹�v��
7�<����յż��L{�VN�Mr�j�ҭ']k\9��o���V�r��P�7ٽ���6�$�%fT�ѻ���+��_\-q�f�Ys�`p�V%Q�y	��5q�3(���{�V����Le�w
s��y�:�s�܇���.�^�9�]z�-ٺ�c2�*�>G�wbJa_�\Z��ڜ�{�ys-TڬO�F�xpߖ���I�+(�;%���a=�����+���=��k���)�+��l��{��}����9(�<�\�Ýۀ��Wr��r�)򉬹9�1�5J��+灬��6���{f�b;l�Rml';d���?a��?x<���z���Y"o�%��޸k1�΄��4�<��W�O�3K"Wq�MB��%���)+�A�􄝸�vF���D�3�`�����9x�dQ`	�Zv)|U�h,�+����Cqr�Z�&��O��WV�l�����϶ Q�^9�6B����:fl�(�^�T3F�o�Ąk���R}wV�h|n<,�#�o6��u��s�C�iu����M��R���Q�'\�Q��. ��ͽ�ѐ��6���w�"�oл��t�=�ۮ�h&��9�su��Swۘ[c)�(}�R&E{HG����z��4�i���1�N+�>[�ýo>0TBo!�9�!u@��h?�l6򢶦�mv�ӽ��58����^��Z�o�9M�h;a�#p��U��JRu�+���/'m�`3�Tۈ����y�je���MsLKn1򳮈D]m�l>ބo\쳷���o�PW0_6���W۳N�����0�ޫ�L�E=�ʹ���P���D�
-�Ωy��_dw=���|���-������ݞ\��)����s��\F!��u��Tf�X��.;S����)I$TLO>ҽ*��L�5�E����#|�LyW�f"�Y���طuܠ�/zۜ1��b�O��źŶ��vr���4"#d*��B�O�b~�����v��y-U,�[Zd[):4����6��+�!Ќ����p�R5�H{1�K��M�Mi)�c�s4mq7'r}�Vr:(��U۳���,r�3p�ʜ,
䴦!Ocܛ����JSϻ{�3,�sJ8KP������U�#���瓾���T%x\,��I�q�ۅ]���:���{��j�����e��D�mK��p�ƗJ�0�*��M��|�x�mA\�p'�*�g�gbP�ӳ���-��{S����
�R���硬1\. ��җPvm�㭓���I�,��5�B�s��0*�I\b��[�2N���lt^�YQٯ��ݧ����ڷ�)JU�������cBJE�w�&�V�ԫ}Y��j@�S�wQ��u�������9��w&Ef�j��X���A�9ݐ��n�)�p�P�Ʀ�S�P��$du-��R��s�k�Қ���r &�1��\�5�0�q�f@6jqtjN��9r
��
AN6��5t�f��N�����t����\�����3	1�	I�l�+j��]ß�_�D���*KEG�W;k�U��gZ����d��޾"l�p:����=�f������PK|��Q���ԪefӽJ�ҎR�9�+\�3D|�܂���.����Yhd�ڌ��L�vC[�&�ӵ�.����Σ��o�B�2�]E[]�}�	Qg�*�� <Մ�8v�]�wv5�����F�N�#��kj e�K̨�Z����K��)&+��A�Q?d��Iio��;�1Z���s:��F ��g�1�7���I.�L���ST��e�7
e���yi���k�/�b��x�%Z>��s��T��ˉ;�o9F[O��lgεu�Z�R�!c[S:�3��b��G���es*�쭸���)>g��
R�s��L������1͑��z�6���(����U�5o�ͪ�*B���1r0�^��d�zCW��-=s|��W���o{h�DRG;�}�.k���zۼï׬3�ts�Y)_"��>����{w���0q��M�� {6/�%�uT�O;y����J�TKtk�I�놶��jۈ��om�S�Ͻ���a��q\܇����j4�W��ܷƠ������6�Oq��=��,��u��p�䪜����|��P=p˹*��������Z���p�O�
VA�=�߮.�ų}���� �{���Ө>@帓�̓1cg���,��vyc�"]r������Ǝ�����G�P�uэ^Ӑ�yJm���������0y�t�Ɣ!>ϛ�,�E}����-�O�6�:����}f�x�Mp��fW�M��'qZ�5~�����Y���u`;{p}=#�,��䳍%���s�7�H���b�i�T|��(�ek���:�������I�Ci �	��bz�O4����\/�ȡ�R`f�`�9,-]�cE��vs��;�������Rqm&��6�js��|��5��L[=x�3K��3V�����Y����na��N�k�*�Q�qY�UF�ؓ,�O���
>��k�~R����ۏ��J{~YX�#���Z�ȍt6{a��UZ��GZ��!�샑�-�:e� ^��^�Yo�%�1����ƥЋ��r�ɖ��w��{���5��4"��C��n$��p�f��Jڡ�����k�R�?Y����٦VGn��\����GC^�Gyq�e�.�.f������7ouU��Rȧr�p�j�����t�N��N�z���K��k�X��[�=�)Lw��m(���YKr{�a�N�<��/���{�Cs{��
�R{�8�n��_�0"�,L<����ÉR��:��j��O��d��ҾIӼu;��rJ�E���^�>k;o�v��ھ��?�0��Yn�ȇ	�?D9M�e�*�5)@U�Ҹ�ا����y���"5cD>�hՖ���T��bj(pz�s�jzU��E):��P��c�����[�-[���NVuv5.$[���*@�f�JK��-�	;��pY�Z�����+'s0�u-V"��|q�P]�삏�-y���щ�?�9��7צ�K{D8ڤ_9Q��%���e�K��X����9z�:��2��yw:��q�r��Jýo��o"�3(��R����V����m��F��������|r��9�M�p醅BT���.����7r^.�����=��Bカ��eċ͸��vC�9�&�q��W�RB�Q�7��/9�����e��i�p��֔Ja��OnmN��T� �\íPS�o[��2���Kt�.��ux�T��G��\�bT�x�u	��dC�Va��ݩZV� �L㔈��ދ���ݟ��Y훚�������m���\oZ]x�9�����^�u*�t2�_��."M�7w��C��\� �N#2��Zo��*ףne+"q?[C3�^eD����nU�HӦ�U)��� ��=�7�IC�O���fV�~r�.���b�+ɶ�&�oqi���Ƣ����lf�g��R|��:^�����s��{��dH9�3"�FCkYyWx�N��
�M>R�������r�[�/ �z�8li������j�}�逭ķ[C]�cy&��}�f��-=�6ף�'���9�}��:���]FԹ��	\it�6���6�ifs�'���+�l
��ta��ڟ���`l�NA�Q�=.����R�q[��F�� ��[g;{����i�A��;��A��Tm$���W����Ba���v)Y�{�=k�5��վ�[���>���&p�"�n����yC/�T%ۙ]Ӝ������;}��'�ؽ��(}�s��8�hr���@��=8k�����z����Du�]-|Cy�X��G�}��ˤ�����o�H�buvY�s����إ*���\�֠*Z�;zv�{2,NK�&�]���Λr��3,�y���r��;B������Km̬���M�U���q���{�Fѡ=!�^���b��2U��}{ݓs���*m>H諃\� `���\�&��\Ն�8t�����K�Y��6���j�
��cdunJ�5K�w�Z�u��^��3����G��W�g2׾���n���Z��ߍ�ǫ9�iJ,y��|���Aum�u{�n#�T��)m����;�E�fv�FP}U��X��'�$*��ok^涷*������k�=x��B�/eLV�`�t7S:���ne9o)[���ݣ6#u�ܤ������g���z��t�Z�j�z���EY��w��7��o�b-^Iz�J�k��3#cj��1p=��L�z�26Vf��;�9P�̨*�>U=��T5aq?Zi�)�����#��1ω��)g����iї�",��?fʐ��� �Qd��f3j��4gV�䟂� �*�*�w"�>� ����g����L-�om�M�W}YJ܏B�{-yw��<��E3ʖ������m��SK���c��X�]�K8����3]��T�i>�5�pU�]p�z�sPc�����<��z��O�[.�P~�j����*j!Zܜ� ,[��q�<������9O8��@b������{u~gH�����WQ�ΝR�Ԟ޸kn1�ڋ|��%Q{l��q/xZ{�G�� ��,U���7���k��m�8���������y3�6�3}��a�nفk;h,���l��:՗Nbeg1ʝ���C��z�*8Z(��:�	糲������/�Ǝ#R��9ch\f;Τ�3�#a�������=�
T4�o�5�7����@�5�k7z{�;f/EoRӏ�9��Ì}dJ�L�!� �P:���Â0ZT�ar��I�ܦ��F���U59���k�WS��#��k�hl��5M�jQ����OfT��W��T�ԝu��Ûhf��nms�̌WMc %{X��{0�U�l8�B{u�6�7>���+��tl$����;�M��^�G��-�Y�I*�zT�X���~�׺�W�v�����v������VR���u�w1��\-�8$��b3g�J��񥓮����!sY��X��e���~ʵ�M�k�y�<�m���nV>e����8�uif7Q�(�^	r�%��5s΍_��0s��6������+*����kZ=M�	G=�ŏ��G�~~Ԋ��r��i���s:���w�bអZ����t�(wb�6�f����{g+�A�A�*��:��n�j+J/"q�/w�Y����)V�}�7��sٚ�/l�}H�l�.���48\�:U=5���9]��OY&�\:Ol֚ɚd�M͠y��ԢQ�H?A.W�=,�$M��F�)�#K��ƫ�Q�:��4�:�����ј��U���k+�)+�TD������N�Ѱ�7����Vicwd|f%�S�fHl����)-y��x�yj���K�3�\�Q�E��޿��ې�訋lc(�!O|�<Pv� 4��F;�3�Ye�:��J�l���(�{"�j����N��BԾ[�|ufսBb1n^܃<v��+�s��5p,Y
��[b�Z؍S)��Jlnj��(><��<߫;O?4V00�S�x��kX��- >o.���Xc�c˙�U)�P e*:N��wi�Gb�e33�g}(��k/4�=��0-�ъT��{���Wnm��P�������p�ø�5^_�JDG��]�Z�� ���kz��<�~��RNMκU�w�TCU^�Y*;wb��Vb\���д.�M��:H{2�e�0�f��_p �P�����<5&��!��\�c��uP��ML�O��w\��>�H=��4���3cwM^h�)��b�
�meK/���@B9�2�E�we��%��A�����b��I)�D��_8;Ml��d^�@�*p�[$#�L���!���z�ж�B!]d����Ue��+y���8��a���ju-/����@ٗ*3v�IhDF���}������Ug���88dz7��FˌwY���}���{|��fN���3�(��JNc�s�^�����j�z�Y5b��@�]�ɦ�ZBAqX*TV�{��]�B $v���c!�		;7)�y��YMؓ�q��>��'wm�K1�V��|{�������L���9���w��8���o۸�m����U��ch4s���ٷ!�H ڗ�Rd��/{��U3Rକ�}ސ�w.Z��&Äs�b$��/]$�ՠ�v]�x�Q74}���mpv���Sq�4����.���亳gbP�НS�z�Y�(ps2��X�[�ţ�M�Z@g���ͻR�a%*���N��yk3��b��WB��`�ZV�F«��Wl��gd�;�udE�<�fө�t1:�]Գ�_F�tԙ�Ʉt�ytS9Y��\8nSR�NލCInm<!J�������3�g�����l7pY��]|;'tz�K%?���.�ؔ��4���>ײ�T*b�3�bq�},��<��A�¯
��T��}E��+`�t�B�))b��Y����{[�$z��*��j��}z"T-��νq^[���h���S�T7
ZC�7���Mt��cU��+�PY0�z�O��@�st7m�t\�p[ݶx+X�H�i"I��H��];�p�U�,)4�͖��P��B=�?K��w���H �<Y:Ӿ�f�i����5{l���e"V7�t�j�]{n{��=��\9I�Ȯwή%t�ʞ)u�Ɉ^b���t����N�O.e�ꏲ���Y;Q�>̄C-9�>]7kC�Y��q����*�Ցt-��_n�&z���Q�͑9x/vA��;u�
�#�7��Y�un\�i�3�Ϋ�PʏErE�Ӌ0�O%��*}�t�ӫ��(dPJ�9�,�V�m��)��-����ڐr.�%g-�����;�J"���:g*���U]��,�]��(%HOqȧ&Q�Ur�Dʎr5*I�p��"(���C$��%Y&BjDRZ�DE��b�!TW*2�Άu�TJdY�]���t�hD��r�p��ʓ+��ED\�=ې�G�9r�.�����U[�/-i�G ����)��+��9�T�T�u �L��ؚ��!�iDF�<����9�̈�
���I�tOS2�Zehyݦ�Q�z \�8��Dj��Ĉ�\륞{�Äp�,$Q*���r�M��z�*s�"@�ʊ���n�tM����"+�$N�wJ*���"�UW)$y�|ψix���0�f'X9���
J�3�g�e��'K0�b�(�j�n��Үs����Ked���/�B	u���pʳ�v!��T��N>7[��1���Ұ�[�0Ro"��(\�W�uy�|U���S1ws�Uߨ�d��fln���SZ�;a�7�L3۶��A��/b뵵6-�J�
�SQ6�j��[���7�5�15�n5ۑ��ƫv��9Ż\�%�C�Ф[�e|'6��i_n�;�Op�ɴG�ߚ��8�p�n��4���%��E�Z���3:��W��_do=�g3i� #z�Tʼد��E�l%�^�~�[�T�A��}E���7���Y��G�9]D�uɮ���rKry�^"��Ƚ�ד�F�#�̨.�	������׏
5������3t��:�\aq6�v�6.bۄ�wV�9V�
��ra���4pe�\ꭱ*�.alTrM���z��%bp&Ȭr^��j���W�,q��W����ڗ5����^�|�5�<���:��kx㮊��)zm��3QF�
�CΝ��ӫlI�vIӧ�e
*�T�3Z�3Xk�̎,��.m���˔Gv�j���ua:u�3��+��I�h��-rx�v̔��B;qo�S��#lRZbd�nܚi��ocL��W{�"�	5&��}�{?v��`l���[S���)Jx1�'�����s&�Gԕ�q�T[=<�����yT��τ���E���̎�U���8%��qe;��m�c��o�52C�����T%6Km�/��nNsF�`l��W���|x��q���N3j��8�Io'%�N.z6��(��.��BE{T����'�ѴhOHj�RY�
�M����녒s����B��H�BS�����_u.{��}��Tr�|�}��rs9�厔Vw5�U�MÖo���}n~+\�����kE�%�ʧ�I����U�f���t����E�`�ǥ��U>u�q�;��T�Eg2'���d���q�F���U4��c�:�c� Z�}B�]Y��
qK��f{Ҡ�n�d��'���Nuc�:��tuQ���N�z��)��g��u��ה{�8��=H z�&%|�܆\�\��o�K�;X�f��ɗ}%�5oj������ӵ�qj�=z�w����^"?"t�w'��n��2ݿ�T�h�`Y+AD�Ӕ�X�P.�Sxf��9���74�\������I�g��)��<~��^O_(�C�2�����`�(�6�^��2�T,�j�)u@�nk40*{:ve61֮<;L��YS�-T����ҭ��gL[���fV*���5хŦ� :|��4-�C�����~[<�T֑��Eh��~z!�
m-��R�Ǩ���s������-K���剽�v�gϳ�|���UF�l��
�S�NLz��Nf[�Yr�u�j��o/硬�ިt��Ʒ�P�@n㴃�����c��M�LL1��:��ϩPu��F��I��k���E��#Cd`��s���r����^6�
q�S� .F�Ғ�U��!��v�^�͆1�W�'�n���S�Â�Ɋ?w���Rѣ��{����x�Jå{(=!�^FǹI��'�T�����9�]	d=��\� -K�r/nh�]d��;�h�&�vrg* ����V��D�7 eY�E�;@�!y�,��Y���8����3��h���r ��m7n&�� �3��l�v�ᕒlBC]
�fC�ד:v�J�d�;5������N�*�F�Hy�+]Z6֢6�-=�kk3�����8���|�v�|�Ȩv��,���ث5�5�ՙ�k3�Lz1ݜ��/@��5�����q?B�L��l��"�8�-��S�^x�����-�o��jx�S_,�&�q����-�q\M	�8t����k�6T<�8���z�T�Iε��C%���j����R�jo��r
~��b�y�<�n�kr��G9|�y��x��啁f�İL]�S�k~��A�d��鹇���V��q�c]�t��s���wԳ�^q�RU��^ ��١{���:ωc��h�z�v��4d8�i3*M��X��滯�Z��̿3B$��XqIy��-龖�d�u�5J�-V�}�7����m�L^�ɛ��&8Rt��֢�����FԹ��pbt�Kb��k-6���{I���ͩ�.P�"�SPz;��[o�W�w^6K~-�^��ũ�䊻�%��
ѳ��p�YDȎ�Z��mo���v�tւ�R♣V������օ0��C���yN]_c��u!������׫�ڊD�wH�ޡ{�#��U���3�YЪ;���9.�ѳ&Vnv%];9, �*���w�SR��+���4��uo�DI|�+��Zp�V٤�P���0T�s5������{D��}��S��Srp�7O���Խ\����6��U?��Ar+��:�(�}�;���-Ia�P_�۫�}����T9F~D)��)��.W�U1���k���L~�����\O�9��n��M�S�g�B���Ꝺ��t�.�';���v�rj#��y7��l;��4�>�!F�7�+%���	��/\������]|�T�G4����U�+'h��s[�a,���nZ�~�,�9���ݚ~�\�b�t�JYkBs836.���9ǇwpK�"�9~ʵ4�|s͟�����5O���Hӑ�y�ao{.'$g>�����$
�6k�2��#��w����w��m�t�u�H���3fR�Y�s*��9��[�lf���՜S"97st��m],Տw����4��3���r��[V�´U��U�pE���j�!���e ��m�l�+75�m�2��jK\��O.f��٧����)d5����ܻ��RD�X��#�FZ'�Nr
j��C��+�z�|�5s�������1wZ���(U�}��3�����*CW�'
�M>R�mf�k��w�����r�>�G��U�;����J��8V�7%̓����э���E��G�:{�f|Q���s�
j��mb�!�l��-��<��U^ꐰ�n�-r���:ny��?"
ʦ�{��g�'��9��9�3��@f,��id�kd�����Z��^8[_&�٭�C��0Wϒ�5�
�FΩ��M�yx-��iP��~R�s��F8{_[��P���}\��}������i^�}�����t�Ơ���g|�f�[c+�(�H����6��z�#¯�`��V��`[���ক�w�`y�L�co�
}��WJ\,&���!u@��h0y��R�7ت=��� �Z�������wu�v9�[��	��!�k���D��I���&��WR0�\�y�hKhr�St�����Y��;D��}��T�W9&�������n�G���3uӣ\2w���ȻcY@'��Fb�e���}=����G�c;�>��}��T�Z�oJ!oN���:�4''9�����g��T�2��V�Kz�^ͣ��4��-��y����� ԋ:��]��'����\6�E�n|zN�Hd�9i��)W��Vm>嵫%�5ء�6�]��_J,g~3��7�&zrU����c��O���M8��if������x�����lD��r��>��kE�na�f�Vy���N�);S/n|�F�Y|gKz
����dj���IvQ�B��S���虺ˁ<��r��ϾS)��Ujޮ���4>E�v�6س�ULm��#[���UW:�gW�%q�%VƢ!5��Q�W����`ڣ��Ͻ��{uE�Hl��}ca��^z��&�����T�,䯴\,h�;�x���W��{f�r�*�0y��;*)�RuFԑs��u����%��)奼�������ۃ[���GCa�8@#S�Õ�n�����Wgq1�s	%�N�\�0��k"�z��e�K;���&-��D�TM��'�]�Sb�7��*P����'���4*c�q�)�˕�襇~�D�R5�2�WB��ۢA���H�QƖͰ�G�\]���6��B�kh\�+n߃���n�i�*��:���n8Y��n�јh���EVGV�ڞ?o�Z9�֔�)�����e�ƺ�m�f�g�
�p{�֫I���e-�AO}�?Z/O5�oV'ۆ��˦kv��^�8���r�m�e���~Y��?-r������E[�yOO2�gK�Ӝ�J 7��hT6�*�(��$w��pj�{A������s�P�n)��h�B\桷���\*�R���4MHٽf���:Ȼ�KȫJ�^����Mm\w-���6�VsЛ�j��dS9��$�J���R���Ue-�����eN-uf��Ui';�\9�92*x4�P����
������?.yϜ!}~�S���g�?Vt�ջ<kY~ӹP�L��tF�� �����S�%ֹ�R߳�Lz��B�f�`7=s����h	��n� +�Nk7�
�/p���o�����/!���daTt���u�ٱ�׈�J"8��/�għr�/1��ԫ�O�#���=� d�Ll�x�]�ا��U�x垛��\4�j��E��.����+���8�yd�.@)GJb�+�.�g�`��I5�K��F<���w���9�\;�xvzrN\)`���e�>U~��^w!�핰7wx��y�I�K#
����~���x��Q�w�~�&.B�������?O:.��+�ܮX�:C�+�g�]O��:��)tσ����7�t�}�~�O�W�Tn�o�IkV�,�{ǥRZ�
^�>�ܐX,{�>�U�3�As�k�X|=>{���{��n�����r]��c�f*eK7gĞ�.�1q�T�Ӗ�����ċ�~���P�#��V�̮��V.�uey��q�Ǹ�ߪ���B>$�3���o�[/5���/�6���23�y���(ͿD���>Ok̭�P��ڪF۪a���s_" �,L�w����9֌ڵ�}�6��u��ʢT�֑7ⴧ��޲6�4���diAϩӚVK�{2�u��,ئG�:�o��X�gQ��c~��_W�G�a)���d.��hܞ�\c�~�jw��}�1�DL�|�V�q�
X����M_����}9�|���=7Y�۱9õ���lI?���^eҔj�;`�����e������C�>zKE��`��(*�tݛJa[!��qy����Bp�P:޲.��4%8I����P����{TX���n]4��"����̥:�<�*������F=ѿ�r�,��ߤ��!��Q�r��}ʘ�~��+�����I�e�����Y�g-�Q��.�����a����4�b?K��b�T[�M{�����#J}@e+Bv�h���u{����WF��W��~ ��,��*A����8��P���n����МǗ'���8�s�����'/��m��d/Uy���R��eA�]H������,��M�6�6�wff������H�\N�]/���q�u5�>���+��B������6����f�K�1m`�q��"�J�k��g��g�B:��\�ӄ�c���ϝ?_��N3���(�)�q)��_�B�O�jy���3��'0/�<P���W�>4�<�^��xɿ_�����'/����%#�e�]xw�8h��sB�<�ey�3��Ur'�
�� �q�؇���¸�3���k�|����y���xyez��윮��F��$�/Ƣ���eQ��Í�W����)��Wm�y�>��'�g�7��C�ț�
�K����_|��u�����
�H:ᵪ��-S:@r�#z	^v�h'r<��γq��H��N���sn%x
��it�@�K��Q�����M���(Z
��y�зu�1��J��+�r*���v�����J�m]<^��DC�ƌ"�+D��ؔ���p���;�y���3on�5w0��Y��z�Fҧ�4��m��RZ�xm����y�㵏ۗ��"�����d9�p
N����5�fe=ỵ�|��Zq�[��V������G�ͺ}৥��u'��G�lQv�:�y�dA�o�D(�/ɒ^�1�+E�CDl=Bl:d�xX�옰�2�*����]�.�������D8x�6��ż�[���R�*�tn*c��]�i���Q~^�r�J0��X�oi��X��T�%�8%���.���t���b8�FQ/F��P^�My�(�0*;�jT�	O���[�FXj�Sv���0�4k�A��i4s*���4�\��H9��%��e,���	zc�;NL�3B)'$���cAlׯ���f ��NšxO.1:���R����~�^�E���/g��<֤�����%���;��K1����9'wa2���I�'�"�.�lQ9�����_v�s&\���e�k/��
ۓ+%l>��Ǉ|}���T�5�@沟}�������$��VP�;"e��y��݃uM?V8��N��H��t���)]�o�C��7:�;JF۲k�	nwh4m��U�V��;�x�]G�j3����,b�Ҍ���o�];q麷b4�R��w7r�*+�J0yH�8���mQ�ۉ=�ՠaY���x�%�s�3�$Ǯ���~oo��T�[C��sզ���C���~Mb��t6��5Zpz +x/Zb�Δ�W}#s0� bJM�Q{ܹ۱ہ�x�χ^{ʖxT�,�A��zP��%M��@�e�a���h�g��W6���r��=͹�r�خ��y��VgPK4t0�D'3�1��#���ɼ�%�k-�3-�gq�+��/1_i҉�7�ۧ����z����<�<q�	֫��7{�66��쵓oY�(���-¶a�,,�=����
6��ǲ��k�*m�D#g}�,I�G��w�ݻ����X\��Z��f�&�<4&���~�#����_c�@#E@�6q�Q+'L/�U�1��C���B�J�&f���'b���ɜo��n7��7���-�*toqɴe��09�����Pn�yV���u�r�	+nM�7=�s>TQ�׭�P��&'{��Fzf����W�~ma���`z�y/���hlw���y���[�\ǚ۳�J٦��y@
0{�U��4b��cm'o�41�;�k�mCO,���Ԯ����n�hQ�6.1q~e�ٟ5��ˌg5F���ޫ�N�NE#6ct��	��>:V�%�"	E�]rN�I�Jg�^���9�1��풡���Z5IP+��=l�P]̥%�3�D���
*L�ɔ9P����!Q��V)�9w!�i�"L�B�<�hF���.R�^N����;�%�p�Xk'0#t(��p�����ud���D,fj�/wnWJ��K=��ѹ'��uӅ���]�Ds��H�s+�E<�3�0�qШ�j��e��U���������&�Y��Ĩ.P�di^븂WU���<�ۥ���r4i���@�Uz�dJ.�9N{��s����
�:�i��z�\]�C2sqf�Pj���J�T胳g42RRCuʹ�I�D���:��{�&��'O)΄Ru
4��T�%=�(�=���9�De�p��E�d����@^-�KNu�ŏTa�Y�v�IS�i�r���kbK�<��
P�fg��f����,�I�J�4:ɛ)v;�V� ��+&�n������u�?F����W��:w�9���"7�<z����e������d�96�#���#�s��}�6�P��o�3�25�r2�(J�}�H�A�z���{=ꃑh�X���������G�d�P���G�DĖ�H��]y�߃�
�Z�8g�/�����lἹ�Aɬ��'t=x��`�}�WM��Q,�߅L7����TU���?o����Tۅ��3�Ƿ6R�Οh��=8s������,��2��l�vy���z�ѥ@�?e�R��>k*J;д�F���WFםxdW��s`l?]�5�O
3/����ո��,{(�ݬw�&ݣ(�;g���7��q���wtm�F���@w�݊�>ɓ_)�(�[>oy��3�O��#�C<�W+N����m�R��Gm����v�d>�W����e��VQ����h��}7�o������B(�P�a\@���9�i:�{;��_m��u^쌏?R�s��<�?8��V$��kk��:�1Q�S��'3L��	�,\Ue^�*|�j� ���_�s�3��J"2�6��ȉ���X���;���{��_>З����Y���n��F���.�-l�����t�z���k
U�C�p�ĕA =�`�#lcU��K~�ən��q8�^�uf�Z�k��I��Ф�\���S�W��jo&��ovRW �
2"�;��Ю��dG�V;�a�~��<9� �<5��w��T���i}/$�vo�g��w�h� zֲC���/��ׇ��;Uó�³�$��r��7%�=P�I̞��T�{.א��eҠk>��w>��7����e��y�W���G��TB��:.-�'���T�g�3Å�L�=��h�@��R������E��ά<�����O�������:�h5��,st*���4ז	��cj<���rAtg�O��X��W�J�-�	������G���Hgg,f*�%�]����^�~�3hÊ%��<��,	�R�Ⱦ�m�F���Ͻ|$_�߯Fh��ѷj�d��x�{:��z����4�T+�rQ�� y���o�W��f��&}�S{Z�ٞ�3)F��=��wZ^W�����q7�Qq�3�J���	��"ez�%+����&��5<��]ޜ7�
����#Q��������9�L�{נ_ޜ�I<)��ƦEdx�kzn�˭��ޭ�)���|���j�F�ޟ"|s�>��@qD��f��$w�tM�:�)� �e�����/:�7R7NY�m�{8X�蝪Gn�.��9��<[��^O���� �ݔ��H���u�Ir�UÒ�S��)��z�)��4�v��9ja��.���.�� �M����E���6[ll�]�Ԋ}�'�faW�̓��߫>6��*9����+�1i�Y��}}c��n��1�4,wx\��o�+�j<�FI����dǺ��1S�X.+{����Q���~��1B���ޛ�Y�v�,UN���*�B�~�f=k���;�Cr>��"5��(fO��ǌ'f�һѱ5�5��WzǾj�#��C�g��t�{&�|��#/e��!x�̨w�Ue���wmO?Z��E�fv��F��Y������9�����P��!z�6�+EGzrNZ��%ٹ��<^z�޸��F���{~�.ꑒu��g�*1�߆I�K��w���Jo�a�pwP�����M�ٸށ���#�:o�(e@��W�N�\u:s�3�z|'O���}��\wy��^���X������<n,��z�����z��:޿U����B�h�1��3�M���k#�թPsk�06�v�T��=+�Y	�-}��FLR�NE��.鼱=�a{�!�Oa�����n��lg1�S��M�*�Rx�I���(|�����^UOz�@�L�z7yzV[����h4/Z�(����Ȯ���Sv<��=�5��tb�m�{���Oy%G+�u�H�ѓt���OQy���;ܴ��t`u2r*b�VJ��L6����t-���J�
grA��GdD��,-�]`#�bIB�Nz}]��O�{/O������<����Tðl�� t���o�G]<��5�Z��Z���^/}1����\I��"<oǴ��G^{�F�zi����,�N�s�sm�nVY�N�}�gǤ��[���e�߃�F����O�ٌ��:�;�N�6��̿i��B��Ep��]xdi&ԉ0��u?I�J{�z�={�r6�W��T|j'�tt\7��!Η�%�[�_��d
��� ��3�����F�'���R����xg���hVϩ�2o{�z�T���Je���;��u ��Y=@��G�QR��NV�����1���>�P��S�9�!z8{�v���Uѿ���u`}��N)i��/�Q���
�ا���]t}t�d��~J����!�6ݷ����q��R��eA�]H�6M�J��G���,�F31y~�Q��v3���ؿ�K�t��~7��<�ϴ�/��x��]���?Vi����u�z7G_�>fp�o��(z�9��*�,�ȩU�n#�*#�G�:~���g���B��F��5��r�ks�F��޴z/%�=�n���*Y.hw�&Y|��x�}����\J{���ZR'�d �̈���4t�G�f��'�����t�ޫ�l�Ոb/=�8>��e�I�/���F��ǹ�*KaU�����eY�L�2K��)�m�ۚ�37W��s�u�����C�#%w)�ev-/>q�K�<�O���;v����~����Ք�3�?���Lw�+�1�1P�a���J%�`Lm(�y���)3���>x�N��4�a}�=�b�����d=>g�xy�W����K��UI�B��=P���`�I�����t�/�#�|���~�;�y�>�i�t����|m�ׇd�pV���I�6�̾�q�zn�*�[�u��<�z��ȱ�F���q^�A�iߴ�����H���ۈsl�m�i}��twh����VCv�5`��AΠπ�X5�R(j��~��zЋ^�Z��F�
\q�����r����x�g��z�� }-j���}����>���T����և��lneB�����.mq��[֧�<��/z���z�X%�����N�}r��hu�| Nq=~�2q�j��w�1�O���}�D� zp2n=��:���K'���o�=1%�z��~`�whū��x܌��΄�zx�yu�f��C}>��B����}�X:��t�tT���f?��&���c` ڏ��1j���W_B,��ɏ��lt��~j�f��3o�L�l\5P���`��S��i�,�9m� �G	c(v'd�=A��0:E�+US�󇡊�����e�Ěq��}/_C��=սv]d���M���ȨWyDk5A������ZǒA��������{�����to�{�{!�د��&K�w��]�����ʺ�]���0�p/8:���V����zu��.�O�h�>�W�����ݮׇk���ӝ��%r|��8mK�1�2p+����N���<�n���^�vFumཙԢ�Y����J.}�_���U�`�^��7����&7�Р��֩F��e��NVF�\�ߑ��^N�Vv�uk��=U��s���V{�c��l��\�A�v;(���۾7�F;���_Y�7�׫�{��B5�
�7쑎���s�P��/*��+�gNIۋ�O�A.�L%�77��d�b���}wF�K�����C�������߽��ϕFw��T.���Ǡjn�Q�C�T<�(�W�Pt&a�mU:���E�h5}^�>>ß?O�VG��{��󿪢Q��՝�<�Ϗ��8}�A�2��|�t��"��f⛫q����#��6�.��`�[ؼ�h}�q�_�����fهp.J5��FX�)zd_L�����ח�����{�&�uՈ�3R���N
���ڶ܎��	�:(X�J� ތ�Щa�aR��8�M]�
u�Įi���N/{lհM���Rl��9�L�j3y:[����� z�AQ�Q���Q�w�uԥx/��b�'��rR�'n�0�	�*�s7�����}]ѱ7�o�ɭ��O���aJ�:6ɖ�G�~Ҿ"WtbS������p�j�f9����ԓ�>�GϹ�Y�����y��~�N{�Fwު��*n#�	��!u׍gGY�3�˳���Ǚ��T�+a�j*5�Q�����Ox��S�Հw��f�s$�5�=^���٫=R1-�m(^Z|T�3�HUºh�ĥ����j:�W�>��'��}>�s`n�GO��I�X"���K��ə��M��D��f�ڟi��z_��Q�y]ы^^�F��4xX��Kx��7�,r�M-<�X4�d��!yQF}����oSΪ�����e���\��%{�\zT=S��ެ+^T��,��c�K�Cd�.ԁ�����ג���Ȼ��n�!�B��C!:�"��>Y��IV��p`o�ԁo��(o��0Ќ˭�;b�b�<G�7�U��4���'�o����+�s3�s)��y�D/]F��h��NI˅,;z��L�T�7ٯ3�̬�m��aWU��S)��|v\
��~{œ;�3���Kg���$�$>�����zB��{�����c�[��Xsgl~��"�h��p���Wq
�z��yһ����\�Mm�[QqXul�G:]�4-��q^H]�L��;�R�)alv��W鯐��c�wn�h΁��s9�㣉� ��;�uv��S�I���ˤ�v6Od����2	�:�ً�t<�#f|��xN������n_�ۜ�	�E�}�$�cվ����sB�,{��(z��G]W��s�����a�i�x����D��Q�h�1_�{���J���]G��3Zb��*xݔT�	>T���uJ�9k*����Ϯ{�/��v���{ooVk��;������qɹ�B����,�&4�����������:Jg���疛�7w��{�&����^�3����*#nSq@�Lm��{>	�"mo_os͇c�:@�q�#��Q����=s�ZG �s�qߟ�Gg�DgG����f]�Ϸ�z.�F�,�[��}���l�?ArD�:�oL�|7C�F����O�ٌ���l�����v�C�S>6h�����½��"���	�(�#~�O���V���Q��F�rV�œ?����X5����z�|Qm�����;u"�.K �7��yH@�>� E<�/#Oþ�������-Y&�y���"ǣ�]и��x��=�����`���K'�|j��h{�X����!�����ʱ�dLb�v�3s��	����Q�T���j��wt��7Tg�#�1��T��o�f�w��c[.�-*l�����y�`X�U��I�t���.�i��O�7L�2�΁ V2�a�3��䭾��y=���+�$�E���9IKܑT�~(3��4�~�~�>���]{����_��k&�}��d����܏��c&����4����*�E�&��t�)���=�u���_z@�t��T�Ԍ��d��}����U���+z�po�k-��S�'NB�~7�j��L�O���^/;�pw�J�u|*/O�;�ި�{
kϹ������daʉ�=_ӡ�UVYѕ*�x��Q��#�!���m�kSY�X���<�D{l�������ӼY;��\�(Ozk�EK�<�O��kz�c8zf+sd���*��o����@}1��+�1�1P�a��:R%r_aCea�����z��EyGq����^�Y׫R��^�T!�K���>g�xyϩX�Y��埈�A��)���p���<07|B�\u[ދ�;���~��ѭ��ϡW��O���\>7μ;>��
� bƪ�|�o��ܽr�z�$ò�v�Ȱ�����4��W��zs�3��<�6o'�R�(w���g�c��Ӑ(>�*2�����i�����>��Bo���^�R�Z(������������"�ٙ�2b�x.��"V�z�H��]����e��:��f�OB�IZ���:�����l� lz֡���9q�u�(-���IН	����NY����oo-qȓ{C�y��'�Ӝ��!�b��;s�g�٩)]�c �nQ��k���M�w{����X���wo�L�;��|���|}DL��H��g��::�5z��/�ݏ]��y��v��V�����{�c��p�냪~��8��P���
}��W��n�xO���r�Fw��|�%���ܩ=�~�0�ԉ�|=87���D����˖1��5�}�$�NX���+�¾;^�w��5�W��9�>c���>�
uD(�߼��0�l
��߳�4�_�K�р�Y�O�W*���S��H��{��F���@w���}�{�L()�F�{ҋ��'2}
`x���F������N���෥�w�	?Uq���^��ԥ
r%ߣ��k+]����WF��p��}cz d�R}�~����=�U���v�pNf�y���<����󂲜��o�T���&7�.����M*�=�DyF׶EH�}u!�+���	k�3�u^�?W2�ޫ�>���s�g ��M2�GN�����/k=�}2��i� ��됝���管�^S�y�p�7'h�|'�z#�u䌮<-by*J�rV�˨x�U��=	}���ݞZ�F�aU�{�V�3J
���,�һLgM���1 ��:�[�aq��h����j7<N��p�{tN�x��9O�M��C�A����˞�-��{���Kܓ/Z��@Мy���{��L�)B���H��s�p2o=pr�����!;H۵]��0�������$k%�����\�2���;9��R���i�N#6�� 6�������`�f�f����,A,U��q̌�8��͐�(�|78��3�B��w������ �������FF/3�ہ4۽��ۧx�̵e�
�y:��5 ؽȝ���Z�ޡLa�Fq��������j
-gq3. 5;�_���oLV��Q���8��e�v^7jVn��-�_)"��b���%��(�Q���F�U����SQa�����{%0o���n����y�m�V�r�u�P�{9]���Ș�-R�K�p6oc�EV��+ز;f	�Ep��¿�F��7���+x��GD�ϓ=�]mm([��{W�x��-�$	n���p�^S8a�tFE|r}q��!ؾn;���v���-MR�i�+,24vF���*#Y1����&k�m}{ 9� �ӝ�[K5#W�*��zO:�	��}����j�|�wח�ke��̵B�23Nl�}�7���s�d��D��L�Ou��Ո�>]Tl����ୡ�b&��� ��\�oWq����6
����͐�,r���nEx�����ќ������-CM�/���F�{�z�����;vm'�N�O;j�����E�Ɇ�a��$��߶���y:�חJ���Q���ӻ�n�:�;��G/��?towW	��]�G��^� �C?XV6F���,;F��^��m�GfDR����N-���0A�\#$�V�X�4tV�r���ݔ�G��4P���9�<d�n����nn��X����� �F�DW�
{M�3��X��vu�������)x������UI��m���w�m�-b���r���5��1���P�;N%O��]��9e�Z�6*�:5{׻l�7�A��l͖���;�k8o��蹶�R�w�7��\��g��~��/�/L��}�|�>�B*Z���X��5�hf8dlL�#$U3J�-[uwRnXe�n���vG��sp] 1*p�)l�W�	u�]a��#:�I�0r�ō�w��2�1f�Ҳ��Rf����L�f�m��H-�ׂ�Ll�Ú�[|���G��l�/ok�I�Q��%��z�x���ᡫ�X,�$y�^;��1r)�o2��_%�R�T��o`�豲%1�؛t���1�)�^���h�^��zX����Lθ�Yk5���5^9����J�¥�@$̊�j��=|���^Gۧ�l&��$���<�+&jdE,�q���ݽ�1S"��&�E��/D�	wTNP��39s��=�3���Z��G0�L(�l�rri�Ry�%wwq�Đ�]����'��NBh��i%T[���D�^�W�d��8��fw'+��fTn��K���м��;��1Mj���p�:JN�{wJ���9��$�U贯w<9�^(�Yx纅��zG0�etw[���2���묉�nw�'%�n�h�����Ȋ�q	���,\���R��
�J�DwwRt�Z*����v�B�)��
sp�H�Uh�.aq=�̚��BtB+�=B��.N�Tl�Z�2�9��zD��'���R�q%iVdQG9�z;�S��J�u�#��TKͨ・sú.���ՕQ32���H-AieU(�."��vwH�x�0�5Þ��
N����^qyS[��C�sH*��r0%v֌2ܨ�v�2�l{�t�kj���)Se�*?���]z���].�ΟT;���q�/�ݾˇ��ʣ;�\;�}�ʙ�l��ݿk�ܝ�rIu2Ǡ���Lus�;�Xy���}�|}�?O�T���?z����Vϓ]����(m�G�~�T`O��:�Uxҹ,�n�M�?_�a�]}B|em��ߟTW�/|���q�ȃ7��\�iU`O���q�-��wP|5����Č���y�|�ҍׂA�����=�2��0�xN*a?��f�ʾ2���rTWH���
�Ϋ�.�n�HLj>�}�q7>��2��=��\8�������SNd�����W�������w�n�SY�^ ��e��Ƣ��Q�����Ӝ}��Z�z��M��}]&}�綥Ÿ���S�&����7�$L�ԅZ�h���~7�F��5~�q�O�>9Ӿ'��Q�mҬ����Y&���i0<湶`r�c�����+�|�߄WF���u�d?}�+�0���3r�2�{ަ�P���]KҚZy,�X_J��x���<�֨�.G��q9)���&�y��KYr���;X6�b|�GB��]v_9z�-܎�n�r��/wZ,kv�uz�]k��ۊ��0�{.�le���'��*�;��e\ Ƕ���Z������-^^�ܕ����+�e"p�ɨ����S�6����W�]�����<ڻ�o}A�߽>�`�Z�,�E�{0�U��3;p-<'$�S� ��io��.;oo����>��m�h�S�80}P�O��W G~Y����}�}�+�&�c�R�g���8jW�>�/���~���v���/]Aۍ��Qޜ���hK���j��fV�q�9�cBP�Bf�TKKC��Tzc���x���\�=����}�aċ>��6�w�������~Rt���d�g]z��N�����+���6�?��:���3��G�4��JG���u��U�VKv��_f��b��Н�<���ۛ���.eG�|8r��I���_�o���{�g޺C݆o�R�F��$���_T�TʯI�Y�į�����lrDo�׫�,G�������� ��~�=�&^�-j�5rKa1����1��w��������]/���⢽����W��o���<�����0��W���:�LM��}�77��x�$p�n��/��.)�\MϽi�>��\u�F�k�~"����~g�q%���[��Ի��'Vs�O�|B���Z�ݦ_/?[��/x�g/��k}11N�v�P�b���?\М��z�� ���UѶ����bh�M�����q�����>�jƤ�Dl�g�����E���K��%�-�
O�\�����{s�[������Q��⏤���끸�/ō�u��HvD�[f����c�����T<����vO�������E9���A���Q���4-[����z�|�F�b;G��7b��{�3�C ֨�9N���
:z05�Y �7��!_W��Ed��w�ӧ�ks8�Eۏ%�7�C�r~UT�������q�_���K'���eGe�PcмX4��7���B.M�єu�}�q�7��~�=� �ޯ���X���T���^��(�ʍ���
B<�a�s�]*�7[>������7�yp���8���N����ˡ��Z�ߟ�[�5L���\�'3~S����i������]4O��~7�j���k�|5��x���e�x�\yTj[�Kk}�����3g������χ��l�wUYgFG�*����Q�����~{{W{l��zn}������^���Vq��=�:nd����|�Kj��r�)C}��j��7��`we.2<���z��<�P�<�xVvT�,�+�0���I��pX���E2�?&�N>���my�i�5�6w��y6/�Թb����`����]�B��y��r���9�3u��*���Χ�Ƥ5�[���n�d1b��钴[ȗ����\�+y�F�k^�H���������b�*��*���!���qr�o�9Y���?��t{"8��G�D(�����=���>�<5NW
]�#n.Y'����.��5��8E������G���Z����L��F�w#���s�'��}�����z�xvM�n;�4�s�&��5d��`�����qt���wG��ޫm;��H�|w�x��!�c<-S&Ǯ�v���z5��.��Y�P@�,	
W��l����>���	��z��3�GޕW���Ƀ�oD�/No<�S�������z��w�P���|}DL��H��^s��^I����>�
|�w�����>ζ;~~��o=냦�=^���d���<L��>^p���7uxjs7��s�7ހ�9\o�H�B~v�������d�{ޭ��뉧>%P29=bbNt�yޣ;�]K�2=�[F�떏W*�x�6��n�Hg���� :�*!�93��*�$��EA�8��u��UOSS�'�3:��8�tTܶv��)|n9�n=��p�W��{ޠ;�o�Q���^���{�Br=YM��1k�*���mY�������*9�\<��]�}X]��F�T̈́.�:�-���wBp��Z�1�k8S[�2�s\	LYz����V��u�s74�3���ƍĆ*��W;�4���4Lq�-��k"p�ޅ6��iuEEm��v��jMܮve]�d2n�2m�����h�W��Nw�o��D?U�nNixg�d�0�Z6�;���t\Ru��t��[ѝuNd3��{�%��SBǡ�K##_�x���=4�6g�q�� ݊��^n��Z��TH����'�]����S@����q���U��g_�x�顺z#�xV{*F\B�N�0�1�K>�����Q�V����z;�^۶r�S%����~~������u�r� ���rr�L��#U�m�Y�j�(��������G[��q��y��� �}>'�<����=��ϕF�Ad�VȘ�qb�Q�Nn<J�{�NI�>��K!���oNLG�Ĉ΅˳��z|��G��f/q�tK�>��^�/V�C�e�!_\.ό�G��4��`@��t��r-eo�����ӿ-q��h�{<�����ޅ^��Χ�q�όߌ8�Q�|ITe� ��}2۞�rPf��{�媷��.D�ע�q	>~��^elw�i�l�8\��J.<�� '�S�pяz�2��u�#���L����G#�ʢT��ϋ��<�:4��}������;�f���Dg	�4���×��k#�q.�L�Q����x0�72����3i�=�*t�:���=N5#�j��ƶ]��ֻ���~�E1�<onK��s"�B^�ʒ�w��}�:��w�B
���){��� (��œ�Um�9�,��{�\�iR�뙒;9*U�<��RD�Kt���-�G#zѨۄ�m�>���>��m�נvІ�����x��k���$�>�R�nI�P�R�Ѫ��o����W�7��>D��;��k�$�ˡR*t�kx��/ë �MzfB���f��.{ƅ�:\o9S���#�|RB���<d�����^�1�K��~�@�gΰ��M(���dLvH/�Av�Q����_{�t�u9��gnzǓR�w��І/z�SG�>��X(k��se���L>��a;Gbl�:M{��߭��R��Ka+��q�{�B�W��ޡ�K7׀�dШ�eHˍ�N��{|��;�#��c�_y���C����9�|O�/���~���u��y��L�r�n���˅	��}�ךW�rw�����C��˽9�+ģg%����~>uK���u���Y���3d-�iME�*�1K�n��5j�5�;#&>������<���W}^m�L�\x��a��>�8����Q��:�b���MO�A�2��,\u�z��:���>�J@��vNݏ'e�js@��;|��ncjՁS�e=���|3�m>ZV��=	7Տ�;��c�FH���|0��'�iFwV�uyV&�������P�e��R⼮�n%]N-��]GM=��w�er��\s���ES�u��h����ﬡ�^�閿u���b�z�Ln?W�V}�=����*Q��,�����2��շ3�/,�ܜ��{쭟E��=u�!�>����	�;���\?[�7<�.J4�$����+-�F����uǢ�{⮼�]y�����{�q7-ߴ��9�� ��yQp�y��E]���q{V��y��@Ϣ$�L��7�[/#]X�r������ZDxߊҟ�i�{��ßO"E��]�I��~!����3Q�Q�PB*��D�u��/ŌA�#�J���1������t�{�٭oZ�h���%{�;�^2+�2Z�&��D�^SB�V�x��s����؍�ޫ�Tھ��CR����O�2����N2]�
OC&=����߫��!}��)�~w=_zf����L���zw����w�w#���wB�y׉�@���;��R{_%�
g�g�Az[&f��u��ONev��۔�WuG������]{�����8�!�X��T��W�2״��Wt��{	�|��vpuӭ�q[/����/�m]B���9���N��Ǣ�������������a.�)56t���H��S����T׏���[�3w��J�*k,�7�wD�3`���h8T'���,��-�{�d1!��� �.C[���B�za4�;� �"G^��#�Cf&S^鞽q�����8ǥ�,#��	�)�i�s�/��'fq��f�9,+:��_��h�9��{iTyC��q��T�]�Y�O�XIsĨO�����7�a�����'��a��f���_���LZ&� �S�����xv�=^W�s�]k=��V;�:��Tg��M����	�,Jٮ*���C�:b����_h� ���Y�o�C���/�]{ǝJ��O
�ʝ4>\fY�����o�c���/�O�|:rf�ty��bF�z����N�exy�Ez����a�nT3jQ���H����<"~���$�����v��T_}j�o[�����+�'��o�=�9�u�ٚw��C�J��Y����/����OT�~U�[>
5��z�KN��}ޑ���u��U�p$��ڻ���ڮa�e���(҂�`HR�f��-�25�w�}^�!5\��M�N�:����ȴ�[��p����~G�FY�\��S0��f���"�k�21�������+O3W��p���r@�
���hp>��u���]��g�pt�z�Q,��@n��1�Dw9nx��;~��[�n�H4qԪW�+YQ	��Y��,���g*�TG<Ehy�"&pP�UuC`m�)5��h�;W#vCq@�a��5��{s�^�sN��5-f���'�y�ԥ���A���nӒ����u�s���Q��4-�v%f}��z��6�G��:��s������3��R'�=87�z��g�&�ωMe��6��L�>^l�Q�;O��&w�Q�r���\?��f�nW�/ޔ����� �T?B���Yt����;���%�<y�:�׃�u��z�BR��?mǱ��{+���9<�}B�zY�ݾ:X	{�v+��&5�Z��S�ΏH���Ϣ�'�4/#����.U��7����s����y���#m�z�Ϸ�@����ixgƖO�L5ckC��i�q�q=��Y����u�Z�Z���.j��C���Нydf�R�}�f�Q�~�t����	��uhv}U����A��h��I�j��}��=��� ��+��U��g_�x�^�ǰ�\ȴ���u섪�{�s^v�v��h��Tu�{n��EL���5�}���#>w/ޓ�ǳ�/:Ad,��k�E�9��_�֭���.@c	B��vҪ��[*�@Q�Y;Jgq�Beh��{����z�y.�>�~[lVt��_�������3��G]W�b��f�z�<���8�r{?~�x�:�ǫ|y#4���Q�T&�j�&�Qc��`�����H�{���
�ԏ���x��`�F=갯�/����O�(�鶖�W6CIv#'�(*O���c����jp�9ΖW=&��˶L㕳�P$Ǝ�Q�|,IK������'�x���.ø�S�X�d�+�g��w�k���e�$��� y2:�]x嬢�xg�����{=g�Z�9��]hpϹǩ��HgS��^0�\�iUA����FK8读�TW{A�IB]�mϛ�����"���z2���ߣ�CO\G���7�C�%�D@�ǕX>}�k�/s[͏P�뉾��>݆j9~U�}�d��y�ti+=�#o�U16��ZM's�^o_r>�s����rANx�2��Ø�W�Ѩ�O���>���>��z��2�~���J$/��m�2KF���f���?D�ԅ\+���e������W�=7g:�*&�rc�İ���]�Qq�����6�\�Ǔc~�v(ǟ<�A�"�7�r��+��0�C���$�n����zE��]wF-7�4}����c��d��Y=a�����������wY�X�HR��V������wz�o�t-�:��=��=j�P�s �d�@ɇϣ�o'���ܞ�S�c=���ԥ�kR�����^Gz��-�X:{�4+��#7�����F4�{�)�/M�dD����{�_0*/�蝾�@S!����������G�_3q���g5VS�<�t��?c*��;-sVl��*n��=���~o�[9&j�`�h��Fu[���Q-m9������'�km#x�F�-�D����I�d���ԊƁ��t휱�C���:乯��ܾ�m[�x����y����,��Ջ�#Hw�xpG�Փ���\@�[����v����5�p���yfۦ��=\֊#MX��� �2��p���w�� 0HF��;���A���%��WK�c�%�,طܸ��[�0��	2w{�-Sy����ǥS-Qn�m�'e�˝�b��S�+F��n��N5��r��E����F�C�� �;w�E	���Ǧ��Ѓ�hTP�>�=��OMכ���7�����r�� ��Wf,3\�#q-7���Z�H��i�7�Y(:�l�l<���S-��w�	�/H�����m��5�]֪�)	-�;ՓA,�K�U�48���\T��X\��xݔ�6�2�hɴ����\!�ujCB��JW��|��l���=�	���G2���N&v���n/bݕ�s�
��T5ص��ir�"�7Zg'6�>\/��)P��<���o9p-6�)��ho�u���Z!إ�N�z��	<�;����:W�4r<�P���I|M+�k%+]�D���֫�/QP�"��4��K�b�t`�U8�k�?��toЉ�D���Fx��{��Ε`�sV�]d=�d 4pӑ��MA�Êa[Q#Ykt�J�H��+���
�%ܾ���ޢ�AEw!js���e�[���_&��hF��O��g����A��0�_L��<;<+��[{�%�o;m�ڔG"�S�.WK��,�!H�z�ԏ�r�J["��5�����C3����Q��
�+3>q��,��]Ւ,�+���'��>�Ugxr��3��R���"�{Y��sG?!������&GwL�Ř��\��
7;pW"#]��Mۂ�K{���Ҷ��\��Ɠ��⓺noj�,�S{�������`3�����gV+����eZ;���)ܤt�K�'mL�ܨ��X\*�>������v��X��#��t��Ԣ���7 �Plrf��bY}w�D 6zzl���ꙣ��{��~�X[�*]HJȆ���H�5�g+���X�-pdmoi�W"К_^^s��*`�p�;�S2	)LKciv��oS������dJ=8�۩��c����6vEׅ�k�@��;b�e�:�I��]fS�x�a�Ŷ��<�e��&��]]^�(]�� �h���5G��®���9n���-�����Y@j�Mf����[y�K:��R���*���9NOhu�|��� ����y�$�YeD���#ݼ`^�u�n䎣*�O�n���i)"�TF�_3�R��u ۵�v^�q���P)����	�����Gp��B���wC��N��e����w0�<�$u��Z��iҸ�.{���n�Y��D��e���̹D肞���E.�N��ʜۨG)<Q�d纺�"	��F��-��U��D��Ug�<�)hY��D��gN�zz��9 S��Nz���,��=@�^B+=<��,ԧ0���ċ��.y;��y;�쫗��d�rs�WE�ZjD�n�Tb�y,� �OY�y��'J<��\I4B����[�����t���C6(��H$�;��&�hG�O$� ��R��)<����ݥ��"Q4*Úx�G�Ћ�*&\�ʳ�s�f�+���Y����"%"��w����RJ�^na�TI!
�Ea!�2T��UJ�X��XQZ�˚�r��ԮZ���XTs���m��(IdF�0YG�f���U��"��2����s8_T��������lDtА�㇤�2��tMt3VlB�gk���F��%���
=\�5��7�Z�m�W5�#$?��c��A-�wx�����㑪_��ڿ3>�2�����������Rދ�q�
in���z3g$�`��/���*��}S+ģ�e������T�|J�LgUB\y���攏f��w	gʳ�\΍�zN���2�L�Wu�<0ӡ�:O��PB@�k���z�����my��x�C�qݎ����qe��fX�x�}u^��}�!�R�.�*��k|�H�w��X�F�^^z=LnD?W�Vz�vA����V%rK!1�#Z	�19��|ld�c޴3�c��Nr"���7�!��V��w>�� �����s�\���ޚ>��V��7�z�C�Oz?��/���ϵ���{�'�����^��=����B�ru|k�?��2�b��Ω���Y yN�%�-ׁ�2�y�k��E?+����#�Ӟ+���o�N��P���Z�1E�=��ۈ��3P�Af����Q��s��7~y֩��y���(�j8(���ͮy���1�=�����'���o�^2)̖����w�������+�Gk����w[���#c�e��f�xY���Go�Ĵ�U.�w���w��Q��
�,��*ﻯUԯ�MB��O���g��Gf�r6c�t%!����y��f`CO8�X��R�ӡ�v������T��.ڙ\d�Z<N>��6���ON�)���;�Tg�WvԌ��������/�b�:����_x�7�� ��[�`��>�3}@�3~�>�<�o��{|�C��Wt.!y׉�x����`~��n�zn��M���~_���g����ԇ#���f���?u�dG����=� ����}���,�5�q�	v�2=s��-C��)D����4u�5[�R�g��s<��h��'�q��R������)��{�+������As7�l�|h䰣N�f��:��:_���n;m\{��>jvz�	���K:�Ԏ�CuK����=q��MC?��7�>;;s>�·UVYѕ*��.�S3Uw<J���א�:~���g����GVq�����E��;�>E��}�]Eq�Ol��^m���{4����4����~21�����^��wHwy<+;*t��Y>Q��~��o��
Ó�i=G�]F��U���y��b}�޲/�/ޞ��W������9\1`ٴ���`kї:���#},��}%��U���E媠Y�������
�I�{�������;E�	��jk�x�}�ܮԥZÎ��Z�)ʳ,����-��[X�'��#R����ͨ�@�1�/V,��'B�4&���i��d	g0h�}7������N��ާs�+jU��ܗ6ā��6�#[�e���$��s{~X��L�����O��u
|	=Q2��U�:����Bv!�~���h��E��MW��]^nϾ]#ǯ�|2��Q��*��B��7�[,f���m��;�% vnl�ZSIF�O�u�Оz�ޑ��3޸;~�f��,��	Q�2[�#gU��F����8�FUf�w��ے����!�}�;c����~��sި8z#�ꉨfK* Ʌ�I=W�.��r�y�����N���u�E��G;ֲF��?;c�H�`��d߽��.=��������#U$��M�w��a9�d[6\�1>�tU#��r�~7�f�n!�~�C����z� �>et�0���{��y��Ul��������eN
��բ�謥��r�ǟ����ӆ:�D������kz�Q4}�/P�U��mG��Z�ʟ���mYw��yě�}�;0i݀귆�Vgw�<ڻF3�ފ���{�rr#K�8t2}a򁵡�T�N�W~[5m��F�rz�[���%�(/v�������ȍ~�����`��.͟��q�U��n�S���ߐ�oRA!�\c���.HOB�3��,9���հ��"���\3�7:>�a�8o__4
+o)�_5�B��Y�q�!oI�"��&��ÏAȅ�<:��� �9IZ��V+��d���������ҮS�X*,Y��J8ˍ�,��DR���1�7]��iW����sʼ:�_3:�KůMӸttg��g�qD�]��5h�>�w������a�b���ȩ�x���� ���쑎���r=u�qy�	Or�\�1�kù�Jz=~��s/�s���<��DB���W�� ;�o��ߜ�p��{��v�]2V
^8��}�H�M�<�7|�Ь��:/���z����o�b�йv|���zk#���x�O�����Ū�ћEi�~�x�S�����:̣L�w��&�,\uҺ��sx{㞹�:伂H��;�B}���z=Lno�3���=�f�aع(�#�J�2�̾>Kw�+tO�}�R�s#���9�>����/�oף"�����P������7�C�%���u�w�	�Qp��.�2�e s��GL����3Q�޿+���yb��~�O�ޢ7���;9}r�l{���c��}2T�̀�h�H�n��-n�u��F�S�6G��l���d{@����;��j�`���=���e�KG`Զl��1/ԅZ�h��e��o����yW�U���w:���ڬ��m|�E��a���2�x�Z��d�+��Y;�X�F�������ۉA< �%��r�8�g��FH��@���;��: ����|�F�v��Z�E��]{�P�"���+)z*wp��g��b�Z]�١�/4��#j�Ufw���ޟ2YϏ�<O�̹̀�	zh����U���xп�.7x��cc֬c�HZ�Z���CJ�;��wF���Q�O�w�`��2M"��HvX/�A�`;^A���㘫%&��z�S�}�ƨ�wzo�T=�Sq�O��U��Dkʐke���n���q�fv�h��8����n��S�>[�W�����2���C�P���x�{&�ͮF�m�w(��#���j��'h����z���A�|O�R�{iW��U^�3��P��=X檺xTf�ơ'���ָ/���^7&����/�N�uYw�*ex�F����~|*���MH�߽gW-��Q�}�;����K"g�?Svg~j�ϛ�P[ó��V����Lo~4��tb�c�7�#���/����u��v�;��#�S��|���
x���>��A5�6��[�5Qy�q]P�\�q�4�>�3��c�{�d}�?s�����
���������ͳ��w����>�7^���NZʂ�)��z�(�	�;�����l{�D��Q���h��op�@v�U�Ї7q�t����]�V��1�m���x�7%+T�ן5T"T�fdS|��6��.�[����cK�����X^�1KǏ�f�3l�Z��wp�U8��j�(_iӹ���U�+!|�V2��p^q�S�U��3�l�Xބ�??U1�= 5,��l��]�����n[�i��s���y��uN�t=��ͣ�y��^!��T���u
@RC����-��ՎG>��q7>��j��k����=����M��>JF���z���=4��9�Y�PB*�}DL�\�X��s��q�Lj;9��zf���X����֙�>ζΟN�7?z��Ǫ�dS�-M���㤌�+�h�ݠ�U{��R�}��n�Rÿ��+����0��ψ�Wo�=��,��߰}���9Op^m\���-tx�N�u��k��9W��;��x_��kμO�z|��	���sWQ��^֭�Kx�W�=3�<�F�ʃ�ñ�����|o���3�utn��u{��8�(���[qe���o���j�z<����]|q���g�\���_9�`�G�N��L���f�zPۭ)�Y��ϡ�*\<�^L��,��±������WM�>ޗ�o�Ρ8����S\9GD�a��J�E�Mw���x��T_~��P��g��n忏�vy�P���С��O������fL0��jWV"�7�J5�@Yy��N^�1ؚ��ފ�q���M㥛vgv�:��p+Ĭ5W�F�r�E)|�Y�҄�q��';�Ժ���e��F�u{A��)$��l��\qva����86_��4����ɉȜ\��U�D����J�:~��g{��ݑ՜c=s:vd��A�y�-�W�=�}��y����g*] �F�����d:~���^��t�1���{Ϸ��*k�h;�k�pU�ڔ{���3}}P��]ѿ��@7��Bz��{e��޹��q^�<;�0_p
33�ݜx���z��#�"�Ğ5��x��Q�Qj"�P,�uP�W����>/|W�ML�Rs���{}�P�M�������n�+�U�OT�G�C�ς�wG���.G8����B٭>95�f��gѽ!q��3���4��liAʌ�&��7e��p�l�G�������'�R<����&��z�ѐ������i��=냷�f���|���Ql_��//j���v#��îgǮH�ޙ���x�X�\4z'�v�g[�?WbR+�+S��95�p8��ϜsN����w<���be�To�Z/���z�H�i��}�D�>��{Ӏ�9b-o��=��
��x�Q �~7��"g�^�p�Z=X����5گQOޤ���W��36.�C�G�"u�&P�s^�<9v�%�0'��H�g�M+���B�A�U$���%��$��!'i�څ�ͪ���X��˥;�**�=ޮ�3���B��+��`5s^k��YˍY�c�c3U���RV7�k�=���sR[�� o�:�L�L������8*"_V���^=g��㟶�Ҽ���ɓpgh�[����4}�z��<�}�%eN��:ǧ��Zt\Ek��r˕nZ4}N�*�(��Kު�}����Uޛ����7���0Ս�p�ϯ�13۰������OdwS�����呑�K����U��
��T���̪p�(S�������ew��E~��TTKS��a�����s��ϫY�Լ^/U�㝳�ſ�%�<��q�rJ�zF�d�z��_��Kn��L��O����#!ܿzNz�5���[��fj��e��[������<�Ӓv�Y?��L�4g��_�7��y���}@;����H�ì�����μ=�Zy�]u	��+��e!�V:j��4�@��xzFLG�āи�i�+˰�ya|�D�w������9�>�Y�w����{�v��e�0�c]�+����x���:s��V�E���������}�3�o�3���=�o���(�>$��M�l��L�A�C"�F�h��{M�����x���<�蛳x��:���{q��sN=��j��xK�� U�s���S���ֵ������=��ʽo� 2f:V��=��#1ága�PD�EB��V�+1:�I�Y3Kκ7˅�.��m� b�Ӑ��g�#�3��#]�]{��Eķ�ѐ���V�z������˘l1��ן9���][�J��F�ޣ> LA^�&����C��o_���O����#�ӣI�|��>��J�<�z�ظ_�je���J�D�I-�q�Z>����h�j~��V$��'�q#ټ���6����{Հw��f�s$�D�Ξ�&"_�
�t�����\5N;yei%_hԮ{���k�����'��<O�:�)�9��= ��W���ϔ���rd1�{��		�͎X���|�>7�T�{ʪ�tB���7�O�w�`��2MB,�����mzsk[��F�9��}9�z2�R�y��_;�c~��=�S~��SbF��4W*3&�-b{޽��{	�Ls��c��a_R���*�ѹY^��#��CƖF��;w�\{'	�yg'!�z���+�=r�e��v�	���P�*�������_��~f}�f�6|=����C5rĨz3���;q�z;���GKN�g �t;�˾9S+Ģ4��1�ǰO�*s3����jڪ�8���J�j{�Ō�������ON0�ݺ�u�Z� �xֺ;5�%�?)��H�����*���yJ��`�f��������<ɼ��ژh���5��ˎXY}�����阶��m٫]"3H�����/��k׬uW����γ����Yƣ�gB�8sbe��]����C�ɱ=7^��e"�-�狥߭���^�^�:~>>�׼{!ڸ��\i�9�U!�?D3���.�s���y�q�w��Fǝ�:7M�e���x=>z=����?W�Vz�p5�5vT��z��8��0M��>���� N�L�&#c�YP]�M�x��z3�p�3����c�v����o���	��N��Β��}ZC>$��0�I��]0�1;��W��q-ߴ�/H�Q�*e��ˌ���5�r�a���ܨ���S�%R���Ib`�^��e溱��S��HC���Ů�h���q���z�=�#o�L�9�YP+g�D�u��~,ogk��5�����ʏ���>�6a�g[g`�wI��\��W���s%��50���'��3J+3��<q���'�o�H΄��1��V|G��Z����k_~[��)e�EOA^n��>\^J
��+�S��5��}�����~x�_}?{��|��� m�o��m���m���1���6���1��P6������m���cm��6���� �6��0`��c���cm��cm�m��6�����m���cm��m�o�l��`�����6��m�o�����)��	Ι�jWl�0(���1$��悪�%E%BUHI����H�T	$�J��RQU@O�H�((��DUJ���*�T�ITU*�
% �J	����eT��
Q$QC�jD������(EWZ�Q)u�(��A֤���R*�*�
P�D(�c(����eI�Ԑ��ATQR$���IT�*�A! P�DvR(�R�$T�R�$�A�R��PB��*�IQIz�������  g�l����L�헛^��)����K
�ۢ��uL��`U:�:����v�z��M+mѷ'8��j��cH�wlU)� ���U�I�c�  �|�U�l���8E]�R��%���Bk�QE��x�QEQE\鸠Ѣ� <���:F�QE�MǣE � ���  ��X   tQGr�)T�kUD�`}�$���   s����E�U�U`ꢻ7s��4����_xgl�y.�]��S]}�Uu���3��Z�����ֈVΠ��]�ܪ�mgiR�%$����klo�  c�*�k�]�����1�%E7S:�������xN�H�6
*�W#9TJ�����r��w:^��
km�R���νsȔ���UJ���w:�|   q����Ӯ�����z������Q��{�Uw�ƹu��tA�(wj흱j����R:޻�Oaힷn�+ǽxS�J�^��eڀz�sҹ�{j�v�u
UH
"*�P�
���   �뮲���{nUg�{^�������@�ҵ����ؽ�]�5%*����W7�����2�^Wn��:ӻ��;m��^�4�J��������l�������R%   �y����Z�wh4�Wv��v��[.�gLƶ��իZz=(Q�Un��]�:O�)��<�+�R�lg�ww�{i����{u��z�$I)(�AHT�U���   �}�M�k��ok�i���+��Nw.�w�g#O`kSk���K���-�:�g��y��RTi[�Tո �{{�m{�z��7m�����ޅl�m*�%%*����   ��}�}cJ\��Jo{�j��:0+F�m��{�=۷��{���۬�y:�[Ȱ����n��U��@�٩[�J\;����ܷ@<���T����z��oG���{`T�!T;aJI�  }ǽ}��zL+Mt�woo{/v�۪佺u��׺�vݶ�5������zz�+
ѧ�Q���vwy=P���ή���!om��PU�xow�w�@-��~BfU%* d ��a%*(� "���T�@ �~%JA� ����D�US@22 I���b�$���fS�~�_��_��B�L����7�b=�a�/(�v^�_z���k~u�}����H@�s_��$ I2B		�H@��	!I�_�@�$�B		�\����W�_�Oٞm;nVn��+��
�F�z�E���Rz3.�Kj��Q��U�ޘ��aX�D�J��(�SU�v�m+c���]^�٤���B���7^�ҭ/XM��D]h��w��u� �GExD٩�G촣.��ŗ{W�1�Q`��E��q�ڙQU�+E�Y��L*E^ݝH0��2T�I�];�tt�5��r�ڴ�'���n���uuv�z��b�V@�����M�jˎ�J��J��/f�u1�wO�6��ʕzQ:m�,i�R�jdX�-�"��O%i��l�$X	KMZzܶ[�^�ʊc��]k��̱��b	
�Q���ky���H����-�L5y���ҋ�a��֡�H�0�6�0��k1�"X+1��rXzk!��� ^m��b̽Q^u�&-e:7x��q���y`H%WD�[EE�dǪ%�Ua�J*�0&2鋵YGM�"�
ջ�ɚ%^�b�.½%J����-�q/���Z���
�!
!{�2�ث$]�L��	,Ӊ��H���^1�{v�4�Z
��kZ-x�4���sr�ZE�2�KWJ��*iۤ6�Gf:{[D�;�t3J�#h�f`���Ee�� �y,R4Ŷ��y���ղ�Wg����uiY�]�6L`�Zƪ�1n��v�Zۘ@j���b�lP����O�:��i�%m�t�k2�3eH�U��͇6�dJ����G�`U�{R�RR�@�7Qk��.�n�mT�dL��� ;*�kk]f`����x�Q�K��[���E�e�Z�;w����J�R����OM�5�~��#V�]�TEG�L�׌��h�;p����T�&�w�9`�v�3E�Qn0�][���J]F�����D��PEC���%��孹��+��]�\E�Z&�CH6�ܣ(�Sǩ"˕��U�6,�3/�Bmh-�Z)֕�l:~���͹�ݻ�r+XoIwbO�+uH~��GU(N�լ��b�٧x������l��b���Ī�66-�3��J�!Y���4M,��
Z���YW�թ��뽺Y��r�
�Dh��p�ѣ���-*[�t�,Q(���xflo17���0�P�;zۭ��e�&ЈT�6�i�@�ʄ��_�ۂ��J�_o�Y�)�C��*S��c��)F컫�ufXPݶU3nK���l�1�6d�(�^�n���H/6�!�pR֝+B��R-]*�U �a�k\�
����p�/.�lFRћF�ٷ�P�)%yc	�zj��Me=�iIVB�u�����6�k��ɨ����30��b�2�rH҉J�R�m���2��i<�`�5��E�SlX©^i���3H�,��V�(�áK�"�;����nF
�X����r�8�����n�j��4�3fZ[m�e=KF�{������7k��.wbQ�1�uZDN�$�D������r$��ol�`[ɮ�޺E �� ���Z�`��#v�����^e��(���ȣ��ۖY�2�]+�~T��AZ����j��Zt�sp��۷�0��!��m�#Q�$dn��v&�m��Y��[������p�"V��X1����*�
X�#�c(6�uM�wx��^8^�B�^�(h���զn�ц�׺.����%8YRUʄ^�;rR�
�������fH�-�Y�;
��X� �4E�է�,*0̀06�]�U��L�EZJk�v�ۉҬg3�f'�f�K;�X�(ųrf�[�K�uݴ��#Y�E�E�F�*blu���'SV�;�ֶd�&kyW Ff�A[�h�ۢ��\#)�;�	n�ZX�vTģn%F�h*��4�2щ�J���Y��Sl-dL���mA�^�ݶ�
!!��LЮ�����սh�t�:cu�u�[P��Kj��A���t�F�ƨ�Pn�8��mϬ���,`7x�&�\�W(��l�.G�չN}�D R�y���ĩ6��n%������t��yw.���#lTC(YU��dY��=�pY
-ЦX�fy�dc*����vub�S6��`h{�b7Or*�ZU��n^�X��,�N�r+9�(����kw,�FP�b��A��Wz�Ʃ�Ʀ(Ru`l8���
��U��2��b��r�V���A͇ ���e5f�c{�f��eaw��I��^-��=����z�X��N�7d+�w��s�S]��E+*�hlTQ���6Z�*�Z�7���EE-yF�5����G"��X��,9q��XN^�Ix�Cvix�W�XN�332R����e�V�	��8�2�͓{�9�]C��ݛJ�aܡN�n���Q0;��\z]h����7�1K1��[�Z4R{GB)����d��ޤ,]�)�������d���7�ɖ�k�z��A�zr:
�Fi
s]�Thnm���e��سSj֜�{��Mkb����<�*��
�h��j��0l	��]^a�j���0%��#p��DV8�^ь�,�N:��ŷ�#��XRѮ�v�7,�va�)]����ޚ(���*�`O2���\j�[��	i�@��i�Ē�V�1��l�5� �Z1�y�v�lF�bɯ$�<i��,&d���ѫ#�Fֺ�M�a��i�m,1#r+n5���0�Q����ll�"�U��+T�ǻA�+^�m��a�//�q���A���4SӍ���A������5^%��lC�J"�	J�,���sr���ɢՄ:t��h'&7F�2�c4�)��ܐ �r�`�����F�+�*Z�l�n�
,f%Z�Nn0f(��Sj �Ê7JK�:���#�J�0��kf*�[����uj�bksN`�B-Š3�֭�bz�}�F�lUM�b���hF�7c��$�� ��A�4��%��3>��<G��ݰ�s&��*��	{+bt�H�V!'��V��jBS��L0U&W�R����Ax��#o3UX�Y)��NS-�����Y6k	 �i(N9u�J�˧�[F���S
MN�{0�{j��ެo!��ηJ��h��/4���S��kX���l`ӻ���r��h:�3�ʲ�M�����
��iU� 30�$�n����Z�8�ɂ#+-֋��t7�lf��T���B+�/���
�,+۵3���o&6�E�ՔuYɅ�j�+,.ͼ�lj��j
�uQ���23a��YSi&"��kb��Ȟ
r*X�5���Oa���[z*/-�Yό�ޙ�w�V8���xfVX��<��a����kY=uN�f�",Vk��M���J�X��e�K7M8�ٵƶ�+,��N@���[�b�� "��Y2�ub�����jn�o쳓�p�vFM���8Qs`��VM�b�GV�t$��P4�P���3 �E5�	�eD!kuՔN�����&���H��H�9$@1�,%�j�aٕ ����9�R���=��8�2�M�v�D��u�2�1:�+ܷ*�R�/6��5�5խSX��H��"S�W�����eӭ~j��X���kv���]�v�ܖ�����ur�`�b5��%�B�}j�Uj�[1�:Xq�U����t>ʄP�ٺ)-еr�f�EZ�:͗ie����J��sU�������̢�!70�Z����Q�`��&nO��,E`��ժڕW��l�����Ӕ)Ű�2�}s9R���H��&��e�w2հi+GW%I"Ձ�,Ҵ�;�t���Y'��]d+s7�+H�=i���`�7S�䷫B����n��b +�)��n��,U5�-������&ݰ��ù���.�G]ElKE�t1\;.���:2P�yW��+o\�i��Sd�"�����毃�*�ſ&��6����GInZ�;�dY�u��U����MkyN�H5X�а�芼IdP���P�����o2#h� wCw-m�]\;���"�HmE����ad�_:� %���\�Y�b�*�5�X���όjj�C.�$�0���0ƐV�n�b�\oZf�ԭe	tu�3(��rKCwcK3^�t��+m@�H&h�l��#uY�B��]4��/cl<�[/ujQ�ˉT�iEʳ�NT��6�7��y�[�*�mE�
.ihnkyxe]�B&�e��]\�i=B�"��7�#)�����ݠ1���ڔ�6��҈��*9��[[�3%btZ��ݛzl0��hZ��n�K���-AI��ٲ�R{�N�Xǚ�)��M^��Яͫ����}���Z�s2��1���jת�x�8q���R���U�H�E�(]�"��KąA6�"̈́0T&�(qT�Zϊ��Q��J��vI��Z�5�Q_:�Aֲbu0�e�m��%�H��)�cb���㡥�Y�iV0��
�W���t�G(b���ZM�E:�6n�kwq
ơjX%)[m�OPP��s3N���R:p�j	�Ȑ�x^�q���V��w�Չ���d�ER}��ihsF6(*)֔^<f�q�́!}xvt�y�v2%�-��˚"<4�BK����ݓ�ŚTz���4M���s�n�,���Eu��Cz���*i5�+�k^�V\{�EҼ�7�l�HG���PX��X�(��Fmhx��@aLj��1�l*�HV�� "�2Q���%
:z��q���n3�wiV�X2JN��vlU	�bh�(��Qn|�2Y�6��A���ϛ��D�&�XX'.������E�M��Y��b�-�I7��R�41؆�����o-����9 ɔ� �o�sV��;va-X�1b<���"�=�(�l*�c˱rVPq~���`�mрP��)9�.˷v�:;�(�R!F�Lц[�0��/��K����Lj�*9)�Ky}�j��T�+l ��H����ܫƚ��9E���.���n�A�6�'n�9Vt֙6��E���@��cp��決sR+�N²�Ò��(d2�c,m,�X2�d˗�DY��٢��A� ��):�J#�Jsv�f��F�ٺ%�����df5V�fRon�0F=�V���K͊V<��(ޤV^Uڋ$�Z�hڂ�Y+E���d����k�!�f�-��vi�JJlaWP�t�r�4n�}z*D�|�ò�Xn܊�[s/�V�j�s)n�C3�H��2�YD䩌���Zt��M[x�g>�ˢ�U��&FV<LP��6�c%�w/HkĆ�4mȉ^݊�{�k��Z*��6�ɬ�0KI]�"+����W0HQ��#w���P �P9fC�V�"��L?hJ��6�S-�S˹SG�7,(n�]��e���0��hݫ2	MƎR��oɗiGgw�Ȯ�eh(��gi�ֵK��&��suY��Mʖ�c��2�i�YJ������b�Q SG.*�D�� ���2��aV�c-eJ�;�$�ݳ�iƝ�gM�� ���fTy�lD�Mݠ�K�6��#l��a�hcf��2�p��+Z�j5,���Q!�6$-�������Ԋ�K�WVRG�0���l1��P�ֳb�J�Lޫg���	V!�ͤƽ����qҽTZ�$�XFI�}��d;�*����a2�oE��xR�wk.�;�GP	�������aZ9e��7,*�q ҺWV�D�!W̆G���+�w��'��*X�-��42��Ad�cԫm]gНӊ���2� .�ل�T���^�1�e�Y��ȣs$T��8˼ʘb;- �F�Z���34�*���R�[�v��hP�x����yO+�V�PBun0V���-T���j��qЀ��;��Q�G�R���ږ�:8�C�[sH�D�rll D��U�Y��Ƴ鶆�"��wo���v��ኗLT�J�M�bl�t�C1^�1���B���trm��O��"ͣoVQ��H/#�K-:T��+֬!�P�&���*)��EY U�cU�F3X�)p����Zhil�@!����+6��eu���I���ۤX	R�*�Rfayzy��Mݴ�yreY�STCj���o�Pfj�l�MQ��l��.�
�5SW);�1�����wQ,0V�LD}�� Z���E/r�ӛ6Y-9�j�mS5�Un���B�%�J�7*�1�r��pUָ�PLb9�x���7jf�.���OM��j��0����ހ�fE{)\��s%�J�1YZ��s(`��S8/9{��(Ȉtr�1����]�-Ԗ.�����զ{��L.�����mC�!�% #��U�^�����#N3S4&�)Y�3��M�m��pis�2�,�d�~	����v�q�6��	�������̢�@�fR!2+vMʶ/[�Z�d�1f�ZsT�R��ϙ�G#N}T��U��`��@����\�
[���u�����0m�%g@r��ڼn3C!��X��D$��Y�u)a�#�����p�w�BibZ9LZ�>�[��5RW{��W[&��>EV]���Wx�Mz>
'O�V54�B�7��[�����R�����Z�]]�˕��l��L�@<�h�M���45���.[֬�Ò��'�jN���b�[ �_a�Nh��Ҁ+���ط�ӈ��h���^�e*�[F����U�ݦ�`P�C0�q�m^&u����r��V˶i���M $:E�L��]ޠ���B.˶5���m+�`�@h��or�@��� �Gbt�ǻ��B���ٽV�9�צp1�oUIs��Q0o�]�ĺq�9w�5V�����W5�Q]JG/�F��<���gIks�"$��j��2�>w��_f�6�%��{�l��B�,��6�閲�0�#�ɱ�K��;�x{�gA�j/����Q�q50D�8��=(�y�؆�X�vB�l]T�WR��6I}��ˢM `�[������cy<[�Vx����p�^�3�t��B�Ϲv�*Q�,S	���r�dY�:g"�ݽ�����i|g*��C]I�ۮE����7��ě�b�H�uk{J��a˖��,�d8����}�����t��B��))�ҷG.}jX3:@on��y�A�d�%Iֲw\���U<)H��}d���\�F����t±Y��K�{	\���͕٘EvS��k����ݸff���%�קln�=.�ߟQ�����˲��O��T�1��pTor'�{�t���p<!�΋Oq=�2Nǳ��wd�g%�;M�	RƯ��"V͋�]��h�h� V�v�����h80'3Ft���8xŏ���{��K;m��Q�㳸���=��%k\�1e�G�����Z/����I�(u����V�����1�WU��n���Y����dz�hzQ�}N�m:F�[K�ߙ��U6vE�����e��<���L�����/�a�X�	Q��
:��S˵�rC	-p��ŝ�wgJ�0�]���9���� [�ʡ��fYk����ƨ:U�U�~ͻ9N���9��l������bI+�7.J�wغ�2�J�N��*Di�#E����l�i�u�]�u�$�r�%Y�Е�[X.��P�N�gi�k���h�V6S2����u5�c���M}Y�Cu��]=.�����ݠW�=T���l%ɾ▫qԝ�uR�囔"�������sڂfKk�R��kx�S[����̯ d�sS{���쵛����֚�B�][Z�j��.�n�E���*ջ(��]L6�YNY��� x�/����-�������W]��WW
���:��<�)�k_���G1��ݭ\�yd{��F�_W-Y�tƛ��˸� 5�1���k��Zo�v�P{��O�_Ew������"�ٽHoO-�	��X�B�w*N���+3k��Wr���hͽ��v��Ď�$x�8�R�LgIjڝ�c]�\����71��R�.볬�]���M�N�Yth��@ß!|5%]�{s�
� x�u��Xí���4���'t7Y��i����WK��f�5���I�$��r[��z{�ւλz��Xf��2��e�Z������[o�򸵼3c��.�;KO/a���i��o�K�;��dX���Ω��9R����X������f_q�s1�O����[9!i��r��������)<����e+ژ9<���ot����KD�Y;�H9/j����V%]P��v��;��	���ݙ����,�D]`U��� ;*�k	5-.���4��j�M7(�Gb����#�;�4�uy�ݫ6����J�D;ʼ�x'})f�6${-���Bvh~�{(q׷wz��m��k�C�xɱ9�)-X���*��r�F�c� ���$�2��H�eh�}w3���U��5�����H���}��		ÍY��T:���͜^E0f���r��#yK.����c1gR�m�7��XC�wc�Ǐ�KA��N��^�Zj�_ڔ���In��j�Q��N�۬�g|	WB���f��oV�k2VZS	<���.�M:D���`c�|V��o[����0�V�!�®�r{r���;Id緤儆�M��=ò����׮m!%�v��2N��B�L]W�Y�^GYٶ7��֞��*�S�	��t����A���V1j�G���¦Xi���.c��(#Ǝ���܋��\��8[���N�b�j;N�O8�₻��w_H��}+���zu��j��%�o�2=����I���+�;����7/�L�J|�0�x
�đ�l�FgaX��gl`�n�s�"��2�f"�j� �ug��Z���޷���cV=2M�:Oj�٠��Ye�Z�&��4��L㨒���MuML�v�:�Y�]�waT��Ɏ����˽]�M���1%@n�=����/���k�q��E6i���7Ƴ{;�w�#ƞ���Ջ�Z.�5�J��m�I���z:.���ֶ�v�e�Z]�W63�On��rfXZ�^ʓ��`���-���NŅ�r�M�5���9��Kfꆴ�����J��5X#��Z��)�A�ك2 K�����;	pK�HL��Q�V&+�{'E�V�xlr���� ��*C;+>�i{�`�鴬G�>����E���P�y�FYP.ɣz�йZ]X�z��z�u�7����Rm��%����6��R��F�\���I����:Ѫ�ʈ���\�v�����B&\8���)-�G]ܮ�Sk:���+����9�]�['�Q뮣se���ܼY�ٌd���Y����E��ħ|��E9f:�f��]7���i���a�����:nݼ������nV,�c�3�<�gt*�͋�[Z^lj5��r��T��t�J�v��]O/�d\�C�h�����m�E��&�v��P:Ϥ�4��5g
��,Ҿ�{e7aj2��R�ۻ{�;��
� �iY�#�+��$�w
�����wC��뢹�a�I��%�(���,Y� 1�;�]��T�̺ѻ�-�^m��cCr��ȍ�̺�Ρ��<O�S���F+k��)��n}��T0�U���q��pF��`�ML�oY���l*�x���,c�Mr���,̫�}+t,��/;��8;��`E��5'x�߈x�0�f�x��\>�
7F��8�m��R��͋�4=%��ε�ZQɧ��x/0���f�{B�܊���XI�S�ؒĦ�"3��FAn���{|9M��ĹT��ttD�嫐�i� �����fH���g x��e�`n�!fh����C4ƌYL�΀���)�7��n�a�D��w��d�j��Ż�u�(�5_u�M�N;T;���#�y�3:���կ�;ʻ��hG"��8�m�4��l�u�m�"̰o��k�a�oP�Y�o�s�nRO�}�9`�]]=����[�@���%� .͕]5��uv��.���ه�-�<g�w���53��{��"@/)��zv0V/�T6r���Wr�m�Ζ-�ڤ�GhE� �R��V�Ь��t��2��ǻ�hMs+2�R�-�i�ܸ��M��mg,�܄WS)T�֜��b��¢@fr�i���N�J��,X��n���NvV�z�R{8������wo�ba� 97hL���OA���`։�%%�/,�j�W~�&�4�U9�	�X-q�����v���/�i���x�)�R�mh���v��{h��&���<�ibk,��`k�E1��A����kc��Q�t��Ղ��(�H��V9���K%�[�n�|����^r�\��5�& ���]ݷK��W;�3o�]>9���f���C{M�V[f�H��7m�O%������oPg�p�Y��Ƈ���[1��V{�*^�xy�prn�;��RE�]�����@����/ ��}iC��
<���d����1�y�}�,�dmE����S��oPH��@o��;���X�\�ç(V��Y��eM�5v�GE^�DMp�0̇kg����ڶ"�k[�otѯ����:H=��Q�rh���������E�T�w�
G�n��o�^��m�6�rAXI�s�(�*m�O��κ<q ^���#�L՝{@2�iR��U{�|��N��� �U�qs]5W}ڪ�š.Й&��J-����YȨ0�ǝ�9}���^�]$4���v	\��
�m��Gw�g=4�Ѐ�t�U�:q�<���z�Ev:�em=ຣ�T��s�*$*GE�k)N��&ӽ�N�Yx���Sp��ٟb���3Z�c���jR�W@��m��m[��84S��=�n����an�f�%G�t���X2�CY�aُm��۷��@����
�O)�4��Z�0�W��-k(fS�)j6���	�v��M!�V+M�
%KOMmv�]n����ރ��{y �(P��3��u���yS�wj'Yu�gj5����A��T���鲕�ޮ�vY��]u����v�w˅-v�:���έĶ�\��ҭʙ���X�3�r�I���jcD.��0nVq#4��L;E��gr��ە�lhŬ�o<�n�Vm���ؼ �-
�7N���:�s��u��7)�p�
�2syV'�2.�I�ڷ�v��=qǚ��p�RL;/mͬr�u���1u㛨�yf�}}w��mF��S&475[��Q]�k�%.5�c���`J�
�N~�x�a�23vjuro�qX3xU��m�v�0.�h.)��&�T�2N��[��y�m��=!^QI�C�5d�.�d/6��f9w��=#r�K�z�V^3�ls+����\s�2)�I�Fr&�%=�f6dް��n��M�:��ҽ�s��z�r�؈��c��m��6�s�ܩ�8��,s�J{�2�^��)QN1	w��.9e�Gi�����z7�H�{�:��;�@+S,eA��
��hY�*_l���:b�Cw�X�u[��>a'�n�Z�}��p����ߋ��N�s`�Σ��uWIu��ejк�����H����J���*i��#F��t�Ҟ<�	9��[�9�� Ax����IR�o!��,�����at��g,� �fܱR�V��n�0�Z�̝R�A�;6��p)��]t�!{Ӳ�.��(foLݑ�2�*Cf���>,3�	����6����)M#%]M�8d8�a�V�V}Ԯ�s�$��T�&V)�:�����k��v��T����[Ңշb.��1N$�{�1�ו{��qtEDo8�c���G��ח���gc�r���9s@Wb�8�%�)d12훩��ܭ,�[V)�G��>o�������CP��wu�MPYڕ0���gZ���9X|�Op�[a�D���ú润�#�dt�d�YѾ�<Ю�5~əOi��jߧ�B��.�����:*v�a�u�k;)A|	��<��z�'�r�4dI�$�X��W�9o	's
勂����2
WE��c$�c� ��}���Z����3�[C4<e<����#o/�w_´�]�����<3K��#`>J�!i�̂�G�Å����(���g+9�\İ:<���o��%l���U�^��aAD��S3�x�g��m�;��>Qe��}�
+���
�S���u���,CW99�j�����#�me�|lw6�7�>})N5��8PpQ�V������E��t���l�w Zl���/����rxou3��ܮn˂�����R�a|9oWe��;tцD�'WQ�W"���zi�	ʔ�.	7x�Fw"�t�K Q���w[�Չma�,��F @���U ���[;r�z�`���$Y��4�w_ot:�cz1�ĚY3u���jWt�wx��.�.;���:Q�qp�P������µ!]�rerOs5�u�gh�3D��X41�,�U�g.�{Bvc��
P��r2�X�b�NA����ob�gp	�U���Q��+YX��]򦻬���pۡ�>U/hsꝕ�'n�[�[㵤Ǧ����������.�j���}���a�P��;��7WLD7��)��ǭν���H{�Y�ՙ1��>呇�f�X�#n��Ȃ�T��δU��ޣLoY֬VF�^VIf>d���l�as����'sd��l�8b�
`ج���~���\�<IȠ�זY=�����o6���1:m�&��sy����Y*�S�M���T��c�qV�3˄��7�Ɛ��M�ͼwNv+6��To���R����T�D����0�7��0�r�,�O����23R��e�QW��r"�[�s�d��dn�ݯn���6����e���V\�k_ĳi���G]��1�{�}G)7J�
��V��N�5vuв�ܢ��*l���ͣX�9N�.T=�rI�{ӓ�⫱l���ct�A���R�66�z�q븕q
L�g+�s�!b�q��MYhK0�O�'_:F�������#3�v���;�!j�ĂH��5�eB�0����2�C��t�CU�,Cwq��A�3�fƢ�Hޚ/z��M���v��݂;:v�]�Ar�=ՔF�cng:ukp ܽ�m��ջ 9sK�_>\�+�MnG���wԸ|<[�7����u۰e�}:�e�v���@mY�K|�{;��Yb��fN��Z�2V�-c�ڡܖZ�Dѝ>�H�R�KML��uȖ�)���A�C=��N�!�v��]2<��m7���ʓ�c�H7b�k��ܻ����o���]f�_Z�;���y�7R�!rf�yv�*A�v���{����]>R=E�'qK��=�c��<�[lg�O�ɩr��:8���v�p=Avou%\�X0��X����v3���r�G�Sa�$F��l��=�a5/��\%pc�N��ЍWNR���45�BpN�C��c����x�f����C�Ayfr��[�mڭ���Vb�w�Zn�\዆{��N�=a(��ѝ�m+��8Vg_�l���w�٤�|�J͠��F|��G/��~X��x��7�ϋV��]�_N�x_9
Y�뽻f\��r�f
��{QM��@VJ��s�OZbr���c��=����b�C�+1�lV�I�Vyd�h���u zs�����[����B		���$�=���<��������^,�Y�pR��X#^&� o>�\;��8�/.1��" �����x���.��cZ�I-�]κ�K"��z��mBj� ��iP��(��@��ms�)72�ʌ��̈n��u��kN��q���D���%�[M��n��w]��J�6��hѴSa���nd �a��QԆtR��C�}�[l^� �g��Xw���B��w��\�%W�z�G/2Ҿ1�5%q	� iW5a4��B���{��c)j'��{�ڽD�� t�8��ë.ufq���g0�+�j�l%	��QI��-�]�
�M�5{� զ'��b
��
;� �u���������ȍ��	r*�UX_�6ƎesOx�nr[�a����a�C0[�}J���&����݈�Ov�ҒoG�,P|-��bp�S/��/�W:G�Y������0�^�>	�ӱ�z��7�}����ټ����^,Ը��%
�_Qs6`t�FS�k~��	��,֑9*�b���GV�b��/,��:%�����|��8�=v��J��qMHb�PѠ闭j�~����A`���]�:n\�/��u�4��7\��#�6<�[�}�KUͷ����+c�����E���gm���1q&��� YF���ъ72�e�� �=;LԹׂ��3��;KJ�ϴ&��O�4uo)7����ߕ��1�����E�c�=�"�T�ַ{}T�Zն�1eZ������W/A_<�M�'}]���ޜl�g@�����������m���E�yq8 =�e�̌S�nT�۷j�rB
�@�4^���9ޠ�cZU1(�f�e-��JR��ys�3���� ��k w�����5et��Qma!��K��B��}�v�ѕ�۝��i}lAғ�Ԇ	��u��A+W^��|�n�"z=���	�h:��B6�ǔ�<^]������Gl��&��oa&�:]�e���s���@p�`X�[��3��4Fn�A ��(�P�d5��Vaз��v�,�˭Gj�B�.�EL�4�8�,��Ok��X���5��2&a�K��TW
�z9�p�a��	�^�ܕ&��
��3p4z���P$�
��wד��Z�sA3#��ޒnf�A>%��v�v��Y�y&������-���<[��quɨ[�r�],]��{5,4���AC�N���I�T{z.�
��O�s>��weګ�5vi*��|X{D�t�϶�N�	�@I�������ܳ�Hڋ���,�5�:Y&�s�]L#�c0�|]�Q>�7���ܛLfiҽ�6��rwL����6.��uh�u*�N�_D�gK���
��l����b�V=z���̥0X��)��r��T�\��$�j��h���#�؀��g�O��U��ȑ"R�v��5��i�ӕi򹊴�ie*G�	`h�'�fJ1W����䲝�u�����v��p{�7�fEL-wZ�5��o&���@��=V6��L��V�1�ت�5�n�@(;���һT&U�o6���^-̽��b;�)��5ĳUX��w�>�Q>�gu���D
(u�5�rҽ��CE�GC��2�����zԺ�5�qs����`��b���#x%C��Wªb�Ef�׷N7'c�fw��sWG����V���B��pwtVv�y��K��P�F�P��,���$�Lir8+2V�%ǔ���W{}�i�A�r#��������e��&^`T���ןv�@uj{C˖@<;�;�ot;��������0��9�Qm�84�}{]W#��{Ȍ�xD���Q�>�������Bp�*��ȟ����Q�Y�������O�5���s_(N.������:ԙ�\�}�����XK(�����&���P}v��'&��\z���H)�\e��,л�;F�����C;��R`ݜ	<�]p�O1��[���-��uP��X�G�,�г<]�I����*��KLF�{1g�CK�U�bv�Ә�1�����;����C_ƛ�s᫱�>Pk��1\��qP��<n�m�u۱s���%��ut(V��d��VuA[�#h�& ����C�X&ڬP9 ��lm��,��E��
�<HD�.�PX"��CV<��Oo�Z���Ae��5w������\�|���9�`�u�tMZ�W	.:�{���W4_�}ǞT6)�9�r]Y�✠��u��.�[6����|�fw43
.U�r��1)�VF>�͡�f�� �鮺���0	н<����H�n�W˚vE�n�{f�դ�΢�K�����������J�Σ���
+���!HK�@^�:w>�v��?7�:��0�X��k��jumk��xgv�'3�v�4��lkp{9N��*L�M�]I*�䀇��f��&���/�c�`�5��`妰v�@��\��9�X;�+eL�{P�Wk�u���R�i��P����{��-p��C�uf,�bW�mZ'���sT�BFW5Ҭ���u�]�若ue��e�޻���m��JU�#J��R��
�v6S�+e=뤳�y�a���H۩�.�o4��A��^U�=��Cm-�r��׬\Q�f2WZ�e,���_e>�8����U��G]���%ٗ����-Φ4hvI	�-J�_JX��/'�rnŗ}˺*��7�3/��ٽ����r4y���+���^�/�I���#�SY,��1",��V ��p��L=�W 6u�Q��u���S���<�A��z�>�X��x�N��+V)v�M�jWN��^����6�*t�P��Gp�5X%<�Gi)
X�4����y{�8b�m�H�ys�w�:Su�\�L;��zzgR2�E��rMˈṚO�����r9��63��'}�3�N�l��qy�w�m�1���s�g��jк����	�Y
ͷ]ڍ�ͳ!���:B�*gū�uX
���Z�G��X�-o�$x�(n���IMy�B��*
�˜���D:J�l�W[��S�Rֈ��f��S��ow{�3$��]��]��C��v�5��zy5.�"G�-ά�)L�μ�z�V�:�Ra[O� �o�Z\K��)�c��k�t
0�k��R�����-�0�t�V��c�)a2��tOU�y6�����K�P�GO��,���%��u0�r��vC039AN��zt<�3x����=`�ö������N�[�A:��(���e�H)9A5��I@��'m)�x����2��`ૺ˰)ۀp�M�b�E�[Nq�Z����l	�g
|;U >E�.X�=�.�Ⱥ�k0\��mbumo ̾G�����빎m�gn݌o�|2���~�ჺ�j��������P�Ҩf�5�K�Hou�m��	�0���d�n)�*���[Frيud�3Dy�j�yR�;���+ 3���``P�J�����c���^k�B���n�P��[5�A*��[��c6r��ww�Gr�e��;�?0�GW
Xyf���\�t5�)V��V���]��\��]%Z���8�3�[U���u0�si�Rޝ˲��0���t��K��e�y9g}ۚ ���ŝ�-nԎ�.����5N�Y�9��hV�w`&��]L�ؠ�ѻ�)xj��p�ey�|��8�Y��ʇ)���[��]�j�nR'���N��[nE-jP���>�'w�ee�ih�f��+��vm�,)^:�ԧQ][�`�Ɉ�Z���3�ҁޮ2�mJ���c��K@^�@�^�v��C.ĭ�\���̙��jeW*.um��:��������߲vt��,��t���2K�pXI�,\�Y\�εc�ot�y�z�vk)��B�wR��]r��cV�	N�LenT-���%��!�N`zfc��L���-]�ѥb��F�5va�L,��w38��e���T)��%�ds�a�t�2�]���|��_ًx�h-)�el�,�>�7�-u��ݡҡ��6��L!��(����4���X��xB�+}N�sٹY��j���r��!�y�xB�ѨFի���AW*x��n'H�~vL;�X�[}нnl�9]uԤ��y��r;D���ح�LY����(�jS[� -���l���,��.R�%1�ugk�8����2\	Pb��Z�O�,��Ū�ٽ����2۲,c��s�5mᒘxs���uJt�/R��)���-{ht�y9�s����]BҮ�lN;�����ԫ����u@��[X:��-�|��OF)���m�p�ҐW��6���/I���c����fC7e�ً�Jx�m���2Xum9���J`�v���ne����jM��lv�k.��Mb��Қ�`r���u�R�Ho�h;����w��{;�-v�0����Fh{��ū[�kY�RYc̽o0[��3��|�L�oº�̽X��7}�b/iGl���M��y��$J��|�*�ޑ�oΦ��i��cW>Ҵ�L]��1���u��z��6hv�Z�\�o1�Z�˨x*l^޲�o(d]HUݪR�����Q(������刧���A�������yPr��|h��rQ|�.Ȥ�L��9�!n%V����5{9�r�b]h�����1�N��&�ty^�u��cv(�;Y� �o0��w�]����Ð(hZ���r�j����N0�D ;(�oFn�lrvlZ���Nl����&O:�qD;���K|`Mu^��6���U�%��\Er1�+��t�rhd�zc%�%���FÝw��6�1YS�9r-}������S!���f�u��UE��sؕ<����81�7�O�uq�٫��>c�t����x�S�Z��q>R�?��
.Ys��݆l/���� �sWT��Uj`���b������wP���+�:E�.&T��8��.T����4�H���m����d��C"7��yˬe_':iˮ���qlŷ������L�4�E�J�=�P�o��R�mI˞�m�oE��Է3���:��!�޽u.��{6Y(�SV����,�n���[ap?M�˦�1����b7G��B�5��,�zt(e %��`s,���[ݠT�&�A�ݝ�7��?�������H�7X۷*�00��f֯�s��fqd<��R�ֻ�N��{�(_.�ѣ�]��FWUҚ�g9'vbE�z��:�j�`[+C�w[��L��:��'�:R4����-�Y�:��8��n�Zh:���ÙV�>س�I�YP�k���,�E9)�|Vk��Oi��5��W`�=��
��̸H�[t{��J]s<FD�.C�7o�u%P�+;�`K)��)g5�56�c{7�	w��o4-w6��s��+Kj��ј6�b�7x�)�R�U�E�H���Ԇ[R���{W��[��WC4��mR�w��u�ܗ�9V_H_c)�h�nt�.G��������$Z��L���xW9���/WR����Uڣ@������hh�$;R2�1���K�MҬ�;�f��NoY%�U��c������0<�U�ډd0W���ҝ��*b��X�w,�d����G֯�He �_0k��M��a�Z}��V�]vov�˒ø���+2���-q��h�B�m٠r4�.51L�#�zч7��@�-ݳ��f�mfRse�1oOcBFd [�+��F�$԰�� !���{"F�^��r	�ͳ��L�h��#�*)�;iڶ�U� gs�؊�ݮT�L#�� y�a\�2gm5�.�T�ԩ����G[b|楴�����,̮j�u�Z�1���Y;7���ʀ�XD��5Ұe��>V[OfHF��F�1���aӗ��*��K�+0N��|�J*�.���x��p��Qx�7t�y�����e���M����l�W���me�)&�s�������߯e�Π�;�3�u*�^;����3�k�bAl��+��Y��+�Un�V-\~6��xW 1 �n���-���'c�1Ƥ�.�Ѳ��V����]��:�3n��U8�8{���-s1�YsUŹ�:l�X��=ѭ����E�ԇ<�G��b}3�a�ѫ͵o�a�ڈkE�:R���Վd�)"�b��	,�`��Y�w^��;_����i�R�g��&�j3(�o
��{r��>C_dJ�N[��R0J���`�JdלN��ۮY��m�và�ՙ4�՗ۻs'4��v@�$ v�%��|����	)�ͬ��W�n�m��:P��m��੻r���QnN�jc�h��P]$�!�Κ��z�T@_sG24��i���M����2BA�]�&�	�ݫ����j��&.
�𙎕�!�m��v�V��u`�j��g	c��gr����~Һ�Q7|M�npW�{�'�a6�(cc�Ȥ�����ʝ�ۄxft�.3�ٸ�$P�[۫��mmҵ�['N�W�>޳����n\D����u��Nr��a�!�gU�����"�k{j�>��R�.k����̷v��VS��y����yt@ /�����6�T؉�ʖ>'Uv�V`�C��P���l�S5�72Yw]��u�j���j�"�L9�LW[*���@�fK�fu�5.���o��tP�hq;N(2�(�gngl�8�|��.��*��}�@B_vj޽1
vol��L"�P�`�	��C�W��N���^�8����5��	����w�zl��{_E��//���4�fxZ\�4�p5!5`�3�v��:�W�f�jf���P�dXo,���>�]�Gz��n�ɋ*,�<��sFU�J��+y�4������$������k�3����t�m�����J����P��^:6����EE�VQ��d<+I��v�K2����
h��۵:���l�K��%>p(J�����޲�Q3���gj7*���A�Ҕ�q2�$�e��W���I4$%4rn���Ǌ��}Bv�ա-[�T���&[��"V�˥�R�����Z+�����ϏnV��]<��mr��a[��6�(�+cG�s�U��+�������MGd�)�����/h���9W���S��nM<yf<���ąfÍV��hT5Y��k��)��f����R6a�mr�*�A�߼i.��"��zBs�'/�tkq9�1�
(�7���~I7.��KaX�dh�+$�o9:�������wҲ�uG�8�+��Lj�W��0��g@��",w+�]f�q���+**�R��v���e�~Z�c�ئ��%n� �p-�k���)ɷ��{.��
����Q�mN�Z8tW��5��#��z�m��]��s��#ܡf�X�IBk���ͫŧ��]y ����M>ʾQ�~`��[���(�HT���]k�o֏&�����ve�Dź��&��_Q������/�ˬ�>���^e�����mਈ.�SS�雄���vfu�PnW��i���̻܄��ux��i�����0gU�u�MuI�`vÂT��xz:N��_�<��X���~�0�wb�0ȱJ�D��L����1�8Z��D��mD�11�L��VKJE�@Rc*��G)q�GQ��*)��J��@S2��U��5Eb�h�Z���(��AQ��,\IQB(�)`5��X�����DH�����bŃ�1�h�e
(�U�IUZc���h���(�b���2T̤0VL�DE"+URTV��X)G+f$b,V�b�E���V5����hĶ��F����F.aJ�)iKl����-j��V,�������J��1�b�Tƙh�+ET"�"1mUX[TX��m�R,c��AKj��EYR�X)J�pdƈ�C(0q�J����U*UQQX�X�������)ǯ����AHN��x���c�W̭y��/r��;�uz�B�|,5Z���)].�>���察)�iB8[Ͼi�wNkt�:X���R��9t4���a�:U�c4j ����Ji���� �8���O2�|�;w�ƻ�wP�����C-p5#D�B;���W%�2�v��}��Iٴ�ٻ�p��Y�q���yY��0)��U�N8)�8�>�Q����,�e<�h����Y`*.�O�_�W�1�V|�⧷�237�
V�j�i�a�OR�&ƐV��o7�7����-]�����!�<Cֲ|��>��9=/�+yt5���pXU�d:7z�d-a�� ͚�P-�T#�o����pV
���`0y����s�����T[�Xtvhk2���K���Z�a9�������y�Jb������o�L}��U�BGӹ�ۚ�L��\lY��0߂�$�b�w8z��c�0�eTLy4�,���}�y�s�-��v/Wړ�7���:x���0I��H��)﨨�w^��4�ʃ�������^��#�ϩf��Ux�X"���=5Y���� �X�)ܬfo��t���#�#3r3º�7�֯�I���s�5N�tqW5��}J�;W�z�w����CX߷s�s�c&P8��yy(�fzmK��˧�6	&}�XŃ�uB1e1�����y�@�n�N1���D�\Vq}id�[���b�+���@�EV^�mr�o4g�Q�a���䱟DUh��J��j%~tb�=0�o�(v�n%�zi᝼4��$���v�eiඓD2-U�ge�u��XYȦ��Iw�/3�.����6ݨY�f��"�n�j�ԋ
��Ϩ&e��y�ޫ�U"f�����?;� ���ޏ_yq���xߧ���/ av�$IT������}��P����j�m�T8lٝ�q�S �~Uqb�â��ff�'���p�:�NU�^��ez�bk��D��x�Jk�dl��o*5�JǦy��3�&\	O��]܅g�����G��Էt�0$�iB���� ���}%&���G���?c�I�os�'�=�bR/49��z�!�u�
�
�]#�<������0u��%f�R%�E�l���-�����ǔEk�`�tZ��>:˸q����f�C,�2�����o}�Yt��b���뤯�pXNP`����c��Y��� �9����U�*o����V&�2�O�9�gf�P� ���p8*�E^a)���r0��W��/ݻ������~(3��M����pQ�t�.�B}��6V�]h��q�<5�]3\U :�k-%[g`z��ָ�j��J6*�/�w5|�6�,�9�޻u��d�Vk��7�BĨ�r���g���*�B�p[�oJ�/j����jD����n!��%�c�ޗ�Z냨^�4c>�pz�c�3��:|�_ޞ�����.��oh�¦pl8i@�1�/ ��X�[�Xd_
���A�L��Z񀸞��'vi�3m&�O\��k���� �%3>�����Sj�ԯ.3��3�����U�9wI淎Ojǝ|bn�}#݀]�"_�f��V�Zi����K�o�]\ ?P@�|s-�.D{�˗��>�w
���a��L�yk�Brf� u`K�H�WU����=\��u����I{.wW_>S��H�Ԫ/R����]s�p���]v|CV��������x����nS�dޓx�}2�+9N\�৮���2m�Vf7xq�(;R�;��^�뽷s8��uٚ�	�@#&E<(P�u�������^�)r��B��i`UƼr��W��w:Q��/l6l'�E�_t�I�8���⿷�l<��Q7b6>R��:���f��`�����Z����+:�cQ�2
�e�x�DsS�z�8r��QZ�-�:k�6�{/��ݡd~��81�sN�K�q�D�~t5^i�C�J��/����z.�\gV�#i]�����775��5�dBk�K�lq-���n�˛�<�Pu9�1�嶶��2YH��I��#�x�v�b�/]&��ͯ9�
��a�}�6�PTɁ��ǋ����%��&
���ItH�^��q��0w�x�N��So{������۞����=~�`�r��jy[˰�w�$͎
yV@���ń��n��gs=3;:�$��u��ޮ:{�Ž*���a5i��2�;�z���KTCm��'�j�1^�e�1O�{�e֟
�)�
��G��U���<G��#=o��R�
܍�w�K7�{�z���m�W��z'���|/k�1�C"�O�5�kK��x>�����.ܦwe5��C~�(�Un�ʦu,��wcr��'��	|���s7�M^��쒲�p�\���W�f���h\��
��5�n[ `�<�K��8k�ېj�Yg�=�Y'i3�a�Է��w�>��F|X����m� ������VĹ�쌵�zT�4��>aH����v	��=�1��R�;e�C<��,�p� #=So�to��*j	|���6�k�)�	�к�"�땧�J�C[��=�J��/+L$5j�H/�*'�A�N���9[�+c�@3�ވh���ȌѲո����3����4��].�i�MY��Ӽ³���|���O)"�qc70]�q/SBwȡݰh�&ZV<�C7�l�e䱭C�[�����7~Z�>�������2�w�2:n���k[k4�~�yO��x��XY��H���`��A~�F-\JV��Δ�.&˹NU��9��&�9f>r!c�2��o{����yB��q�\����Ew�w�H���E�l��ر�l;�}ΔI&cZ(&Enq��܇�#k��rv�U��w{[uí)u�Kr�W��S��\�� �(;-\���u��s\/s�>�������G��g����mw,����]��KA�2���BXyi!u�[�˷X�j�:5�A�zZ�;.�#�w��n���o]�LP����q�O�ϐg�����y��M���~�v�HJ���}����L���CG��=�F`ޘ)[܍Y�-0O)`�ƞe]����c�)���zD5αZ�T��.._�z-��7��J�&ʉ�׸����Lz-�F�>צP4���]�h�ۃAw���
@w�T���i0KUb�C�=T�:�a�e%c��&�(�E�C]����E[��S�18~�a@���3��yVG�Kt�z�s����c�@��N�6Q��5;�KV7��Keu��F��<�ef����Nz
X=F�ǔۺ��3V�%F�o��4�/]<��Oq�i�-7\E���s��p�*�,v�������1gb�2��qF�f�/����֛�f6�����q�ɘ+Jy�/���[ŗ�Ҹ���P=����sfoi�����Ͻ¬�sˋ�m�3��3��S�Q��w^�ll�WۏA�ܥs�s�Q��V�R�B�]C��Z`"���ҡ��bu9Bԡ����$���)�u�/N�+pf�xpϫ�.j�qL�C�Z��5������ÿIk��ԯT����;�����nz�=SpL�x�+���h�\dXUq�e�u��P��+ޜ�=�wt�z�TQ5s�� Y�f}�XdX�hm��֫�,r�Uk\k^��]~�w��<u�A��;�l�����+�D!�`���ͣ({�Պ��{7��[�Y��^�q�8�HΪ�gd�Y�J�>|f"p�S\{����^� ��v{_^��٭�e^�u�9/��zV��������;�i+���G�g�d�W���O��Ȋj��K����(c����X�X�Է��l�\hٶf�֧�p�	����*ҜK��ش���=�����"��Ym\ %�L�rR��3N^���e-a�t���}�;��u����G`ek<h):��~�>l�޶��2>�=m���w/5;��t���u{\�ڙq��ô9���r��W�����ua)����dc{��]�x���>����ܫeg�@O���S%tk��z+�}���.��y���hz�eq�iQM�36U�w�����ұ��S�Zb�N�Z�e>���p������.��󎫊x9Ľ$+�7�)밷Y���$_V��[fmt��8������ժ;���OX�V�ڇ�+Ǡ���5q��/��`�r�r�i�B`�n�f�ήT���xV�>R�
Y�"YB�zי�溞W���x^��Z''w����;���6��^��>FH��y�>�	�<��V�د]fc��,�2�fS[��]�����ڎt4?=��y^����]N��y�ZF����5[A��c�d
AV�8�]tm��x4vP0�Q�@;���@���`�GGTy7ţ#�/>g�[��'�e,+\�n���T�5��7��(��`�J�;�q�2�,�r}�d���k�4�l?k�+sr��H��/$�fNd��U0k��u�};��+(��;�˻'�3m.�����v�v�no:��x���C�P��^�ҋ����_g(����η���fi���8���'溢O��/}jp�wpL�a����\��ss�я}2��si��U��]:��Sq&����?73���d�i��8�~k~;=��L��7�f�����LsǷ��)�to�E]�pV�I�,J��z�<�5w�0)r8�״=Ա�{�Û��x_�$f��X�r�����W6�����z���]�/br�	F/����E�
9��!zo�������[�sF�P��y]��.U2�j/�[�¡{~����U�9ş.��5g���C"w7���vxG6�X�`͛^+3�32�;²5�����f�y�~0�( <]bw�H�;G����ܼPcI��7R�0�En�N�"�m��כA�m(ݵA�3w�^L�N�����\��n��1�Օw.�W`�:����pIҳd�����4oT�9�3��N�>Sh]��]����.�p�R�9e-y�y⫔�`/Z��4��%k�4.�;�;��5.�&U��vj���K�ܮ���1Gf9ڪ����3��P^ݡ��B��{ ɯ^���[^�O�����.g)����`��j̮��A��A�^ֹI�^vz�7y�Օ�N�.��c�Ї���Sǵ�[��RΨ~Ej�&:eW��{��rW���lbu"4�K�$����~��jX����Y}�Dw����Gk��l{r諾͌�˚�eY�v�.#��f���hg�YJ�qp�)�L�+>��r�C�nu���͆�����+�D�m���8�ߣ˩��n���0�\��)+��hΫ�g�Ny��u�\�5�1����s6����.�N�Z��p΋g�k����gS�O��L��C[���ǑW{��d��&	D����	u�Ҷ��L�F駚i2�|w��@͗�u8�Ɵ<��x�57Y�3�B��hYZ���D螦3m�V�|X��^ׂ�&�q�ҧK�؝"�Mv徭h���M7�([�q,�W�Ke�F���.t0W*�Ln��V�`J�A�yV��j��{yK�̏>�����;�u�n&�ge7+՚L�n�n�=P�����8�-���v�k{T{�����t�a�M�C)������;��ώ<91��ݓ��ي������]�},kzD��_'՟8���M��gu�ľ8���3�m������nʜw:���O�jq��h,����$#�r�dv.�]�9�z-&l`���6��R����#���8�Q�v����>u:�o�ց⼍5��YGr���w�]t�	��p϶ܰ�Ų4��v�]���3Пv����{ށY��g���8нb�H7��!����:
!��kϨ���{u���o`�{j����;�z�����`����`y��W�
I�	Ҫ���O�G=����o�Y�>/��-{R���u��V�+�B�mv<�_I,��V��i�f�IfR	&����)xK���U��ukM�'��s%� X�@Q�u-�$��̬��<⷗��m�c=i�f�jƾ�+h�=F�u�[|���P;.RU����[\U��D�B5�������u.��)n?m�'Г�wh���/����E$Zۗ1L��J̺V1���l�[m��F��d4��9��3��^!ۜz���z!��w:9����R�]^�cfs��S��+�ي�ŁQF��{D̳w��<�k�dT�x��L��5f���;&9k��7kef�-�!�Tz;z*i1��LyW�[�v��^0�9�)D���P�ڊ��@�U�&\�އ��Py/h%ۻ��M�Qv�'wE���+�a@�7�Y\����Bm)*�s�l�:�e�#UE/�ع7I��C�7��_l��|ޗ��"��!��( ��6�'=A�e,^eo#��:���Nm�1�S�ז=�|KyDm��U��5�^Mv7ggb�TFvn�MP�\�vul��<��`�ma.D�`�c�ͧ�I�V	nVk�}�g0i}��v<��*�>�SF���E�ӑ�ƺ�ε]�A����mU�0;��֚Y�4P�/!�H���>��:/G`��t���Lx�]Ľh�_%9������>�n�y:�w��=�����:z�qI\�/�>�X�V��"��f��[ۑh��]e�{
t�7J��S�ٻ�b�49���`̳�;��r�>:S&����i����[�8L�4�!��˃]!l��#y�Ѧ�#��i�}o��:�Ӆ�K�$��UI�Y��|J���j.�]���.��{�E������=���U�v�^(�\oug`ͫ�I�Ԭ�OK(7f1�͔�N�:��ǡ>\�X�5\�Bt�?z�]�C��7Y�ղ��Vk����R'*�����4v���	�`�Yn@�7��r`����Ж��Q�J�i�r�Y�qLwi�.W ��v�]��7zuN��ц��/j�2���ԑF�/DCGa�f�x�ܺ}er�S�58��.����v�N�Vy��Ŏ.�e�5l�=�����_"_*@��{�������r�q��/-/�厞z�J���pg�ǎgڰ%�\����u��4n�3�U�����7
q��[��M�Δܟp։�̩vԇ��(�l���jp'��G9��q�J�٠�����������66�q��M{Z���3VŦ9�f��m�������h#t���X�4�[*�xݓ}y��!�Vel�vŌ�}8U5V�7�j���ei��g_Mؠ�����6S�z�N	�՗*Y�/]J�M��DM"�Βnf3N� ��c�7��.��H����(�-����l{���T��m���m%�GC��z\�Z��-u�E�3�3�͠�#��Qf��߻������X*"��,t�)r�DDX9J��DE����(���JbW��PUE2ذS�����ۙTE�EU�����1P�X9eAATm*����q.Ym��S)L��"�*��RU�1AW-QEE��EXʕm���cX��J�ѥK��-(���E��*��%�\�d�VQVҭes2�TVeV�X&f8�JQk*�faZX���E��ʷ-m�
bV0�m���X��4U2�+( �*+dPQKf9���2��D�V�r�Hҕ���6�d\��ċ,eUJ������

(���1+l�+q1�2�6�k1s�X�kE2ڢ�q��3TQX��faKn4�Ub �\���b�j���WՖܹp�\F�5�G�,���Tff��Lf�S���e̹iLqp��2�-(�ե�\G�ʫj�b*[X���i��m~��M�Q�MƘ7,W�v7�!@��n�!���#gt<�8õ�[M��"2�;�t�κ����:�-��|��yx3�?���{�۬u=�V|�y�l�h�qa����ܬ����a:�s*�kWa�2�.%����͚�x�q���W;}��}0�Vs��=��#�u�7Cs��nk�S��N,�HΪ�fv{<�,�{j�R]�V�&���|/h�1�ON��=���3�[�K͏��^tv[�WG#��vph7���_m����(k<h':�SB��6z������@��@��>�oWAO`�+E�6�԰����^���_gf�I���}n�q�5J��)�v�_�伪sc��gD���q�LݶR��$�F���J8q�^�����?9�y��(����=9�k�S���,�S�4o�X�=s�Ǔ=A��w�ZT<�{�_?m>���3�|V��Pə��f�	��X{��gE��Se��ﶤ�7:��ɽ%�g����P��O�b�\��}X�h������5``�/5�90�xP�\�^�-��S(�sm��;t�Nd�5�� �L��R�ؽ�3s����co�4�q���8�R���9w��-���#�������=J�R�vW!w�\�n�o�3a��y�*V�����qy�=6�f��#��Y�풋��w�"9=~a���Z!+z�M}{۷�m��g���[J�Wu�ʺ�v�����X�m�sR����Ov}W�ՙ]����L����o:��W_-/�M�ԨkX�.�Tߣ�)�-��vS���6��p�U�*(�u��S�`-�L�y���Th�IӼs]�9���ۓ�U��=��R�LdwT�1��
=%��k�������s�!`\�u/��+44&%^�?[t��iɇ�6�_o(r��@nu�	��������w��"�d>ہd[��)sI\������yO��Cx�K���}��<��T�lr0{wK��}量zb2L�?d��+�.�\�Bz`�hx�E���(�8��<���\�t��o��w��h�&��u�@gq�OG�m�K�W&db�W��m��������3&�IɌ��v�@��;��B�t{{�V�*8��җ��ΰ�wjq;쎮��)^���5�J�uV�ہ�$��Oe�Z7���]�d�˼S>v�"����>yGN�N&d�Cc��qsds�i�[��Ҳf��e��b4:H�Lk��,9�I�:|�q'soE��{�V2r3)K��~��c��loDh�*�.@���~ϦG6��/.�r�[X2-E岰㿰�Z�N��4s�^��ߴ
r��GGf���ȟ>3A��Z��:ϊ̯32�;²5�����{�LaA�85,���K�kdʓ�qsc(��Y[U���ey,ʯ4/#^�W���W;�gT����S獺���s�1��j�	���aK���Ԩ�d�Qކc���	X+����nXN\��w�s|����t�P�s�TZ}����=Qmqp/�]]gS�(��a�e;��8(0�g)����{+����(�6�}j���-�������$�z	B��<=��RA������h�Ly$/K;A��>,W�;K���.�๳c���3����K�ڃ��鄜�'[۠�lWn�ʈ����M�S-�[O��҈N��lm�����.�G&/�Le+��0�۔tbmɩ#�uf���r��RKBF��y:mvw���铮���N�W,�8��a�f1������Z����CEr�&�{O��s���d�=�6݊��pV�Z{�``ƥb�u�z�3���4�Z溋�ˑ��d�v������ϳ2�0x����eWl�ó�$�$-��>�ë�:�\�bXt�(�]�!X�G��2�ΘΫ�Y��y����*>W{>s�+��S��b�G6��>͉:]+��A�J���u�j�~���o)ȁ ��ZǇ�zZɥ�'��45�:�en[������^}q�㥯��[��p�z:�su����e���%g:hg�G����W�:]-�8����| �'��|I�2�W��� ��Då�~����d����'|ʇ��:��O����N�oVJ�'�[	��N��/��>��Oյ}k���i�W{�����~a;;�f�8�i=>� |�d����O��o���!�)�N%Bo���&�|ʇ�,=d�=�z�q@��ҏ�~?}��RJ]a�ٯ?u���O�Xz�m>gO(i&П�����'X�x{���:��ϵ����;�:��'����u��P�<�q������x����>�t\�����m1�n��g�����糣�A�~����^ ��� �.�r�Q�i��.�t�Tk�.J�5V׵IS%����U�i���A��'���U��aP���W������(���އ{��qS��ZΜ�m������u�s�k�̭j���?+&2~`t�'�I��i��C�q�I����Ԭ���I�'����Mn��d�Vt�X�:���:�d��ϻC���x�>����CS�����_�?}�N}I�y�m�z�3Y%d���=jO�8�L�=O̝J�0�aS�}��I����u�G=�T�I�T׽�����g+\�w�rW�~�q7�=����Y'�:o0�'_Rm�߹�O��y�Y'O�������Z��u��e��?2q*VI�OO�`q���1�����y>ޞ�_�~��:�3���)=I�T��d���r�v�u��3 ��'̞s�$�~d�u�q��k5�T�$?����b�`|�Y8��L?}�!���g�e�����f���|,��?=�0=d�V��`x��N�C߻�'Xk���N2~I��;I�NϺd'�MC��VI�~�쒤�!�ٴ��@'���4��ߗw���8<��>C����$�'�|�u4�?:��2q�����N2w���:ɴ�G�ͼd��'�� ��Oi�s�I��&��|�}��8W�)�U��=��gp���ABtݜB�x��@�N��(�m'�X}l����08���a������g2u��]�u�'�>`{;����3��w�=3�C����Z;��=9o��bq��|�Y'����	�봕��Y?@�N$�(�q���k�\I8�9HW�N���0�$��<3�4���|�]�O�	�W�kz_p���?}�>�d�0�f�6Ş��2jw��q��IR��'VM�d�e':ɿ���a8��y���$�'��2AG�~�j�s(��Z����w�bo��1�0��p�Y'<���'z����?2|��C����&��̓�5�2J�$���
ɷ�L�q��N��� 8�� }�oS�;p��=G���ڿ#�!������t�t�6t���Ibkd��f���%�lq}�����n�t��)`��<>�uj��Q)j��a:<�I,e;Fx{F��\�ep�-x�X�j#���b�ښP��Ե�R���ϋ{o���L#T+.��Ƕ߽����=d����B�I�=�:�1+��a��h�ri'R9܂�=Af��C�=I��bIĞ�$�Y$9�|O�~>#� ��<�}h��g2n�G������ɦ��w�d���k̞>�xé>݁�?2qO��d����ϰ�$�����8������'>J��t�R|���Y?0�d�[h����]�fs���+�I��P�>�q4e�'���̜d?j�'Y4��7���i��_>�|�Xk�è,���ì�J�k���>J����f��u��������o���T�w����l��̒�$�&��,'��4ʇO����8�l���4�ԝI��d�CL�A�}�Ğ����h����P��WAd%\�Z�	^-��������xì�?$����2}��&2q���'�d����XO��4e�d��OƬ:Ì'�l�~I�o$�����q5T�(N�]I�����s�	Ğ���3I'�xoxq��XO��:����́�	��2J��z�La�=�!�?2u4e�d��Oƿd�H��w�D���tT���Y�?u8w��bOP7傓�O������I�9��?0�a��d��	�ް�?2o��M�N��IY:���%d����/�~��Ћ��?�?	��'����ߡ����hz��vk���N%`k�ad�Vjy� �u��2wvI�B��q�&�=�ܒz�&����'���+�w뻇_�?k���{�����VN$�*C�1���SN��k�`q4�?:��8�ĬyH��'_߽���k�w�N2~d�h;d�'{�$�~I���`)���y�����]����:J�>N���V2
m�I�
C�:�ԩXO�q=�C�~I?<3y�s�!��񓌝}C߻�X	��s�l�d��������4�S��6�6.d[}���@ֻ/t� |%��3�k���p�s��Gو��.��,+�5J�$��J��;�ӫ#�Xw���o9:��	�A`�t��.�'�t����T@d;zGR��sap��j�YJu��NE�\�h��]�!�����lDw�� Q����0��w!:�2h9�B�O��?d�	�Y�*N ��l�I�N���M��~>�l�	�xg08��ԇ�����g��r�����~��9��~���ߧꅟ����xs̓��Oi�;�Bm�d��I�?sY%ABa��B�u+'���q�iF�OO��n�'���:֊�1�����y��O�Y|�]}.��o'Y'��3�i��o�s�i��w�'SL�I���p'P�&���RN!�sY%J�d��%d�VO�@��m����Ϳ��{|��};���I+'�Ӟd=�M�u�����&���2q�m�gp�N�Nu�2m������ �G{�:�̚���u'?RVV_��]3�PS/
�����G���݁ܤ���M��G�06��t4���N���W��a���&2�����N�2q!�;�P�OPY�R����[���}Ss��矤���+����T�����d�'_?e'M>3_P�'����O8�۰>N�i�>�u$�T?N}��Y&'���q!��r�G�{�*����n�ޚz�߾��N%C�,�Xz��ް��q[�$�Y'4}�,��$�k��'���(i����0��d�z}�@�4��}���=ޙV�r�Xsڷ�ұϴ�H��'NoY:�	�Y��d�+�Hu�̞���N�zo̒�I�'P�}d���'�SP�q�ה�?2u�=?J����4`�6�Ͼ��iq ��ex��4o�u�����:������Oq�ﬞ��z��'��g�1��M�z�N�u4e	��&�A�q�zʕ�>���<*vr��?��~~~�?Q��'Y<���>Ci:����&�u���u4�=g�y��8��y�q���>�ި0�?��$��`~�Rm����"�O��	w��ϨA�ʍaէj����|1֬�K��������in&e���,-X�Ȁ�0n��1J�R�J���"��� r���6������)eN��|�
��.^��x�I��0���VhTij�F� [ʬ��c�>U=��SU�+G�����=��no\�Z��!�m��YC䓌��_�b�?�06��MO7�m2u*y���:��O�'X|o2u�~�Ow3����_i���>���5��Bn�����~������r�����m
�z���zf�M�S����������J�ל�):�ԩ�;��a����K?}����?����~�����}��w��O�{���ך���z���sY'̓��IR|���z���ÈV�bN3ٗ'�u5��Aa1���8���� �ߏ�~���}�'���_k�\���ws�׿����I��.�=d�O�ʒm�&�u����~�쒰�!��z���,?����5�M��j}��SL���C�8���qu��}�wW��k�o7����d����t�rAB~����l��9�_�4��{�	��&��	RO��s�IX����+'X)��'S�$�3��9�g{�����~�����y���k��3���V���������d���s�m���Ěd�&�w	�q����l&��'�5��'�9�$�(L��B�u+&�L�9����׾��|����N2~N�I����k$�h<�C�����=3�u�z��4��	�w�q�O|�u4ɶ��w$:�I4wX$��Ο~�n��w���ﵽ�}�*
�/�*ORT��'?S����3Ϩuě`q6{̐��:���'RN<a���d��f2m��Nw$�i�h,�v��s�x��/>��z��Z�Bz�w�`,'�?oY%J�d��%I�VO�I�O�:�t~��Ha�ri����a��a
�Hk߲m���v�Iԓ���)�=������g������<�}<d�C���:��59BuY?��'k~d�+	���"ɿ,�I�O�=8ì�d=�����'��a��x��O�x{����}ޚ�Q6�败D��wˁ�	�G�D�s�f��L�dU��`Y�����ʿOuĩ�Ӣo�s�Tv$I��ӷ�hQ�C��:lT�j=�qX�u`��>.��"]�4nn:�Ӓ��-��ۛ�Qի*���� ��+�ݻ9h�x��.^��|�^^`�mȫ��q�宅~�~�ȝa?&�O̜A`s�
d�+Ct�Rz��sX~d�a���W�I�d�'|����C�����写8�w���h�~���5�^��>#�#�#����20�8��o:�m�CG�è,�����M��5��z��>eC��I�'���'Y=ߙ%|I����>�u5ϯ��6\�mG��A������6~��������z�2|é=�́�i��/��0��:�7N������ì�J��i&�zʇd�~�=I8���=}��|��4kN����a���2x����'�=a<M���I�'�5�>f�8���O��'P_>�z�P�y���I�<��u��P�;�@�&����y����?>�����g���>����vd����z�:�״��'�O�Yd>g4�2βOR���`u'P�<�(~d�'��m2u+9>��N��9���I�<������;�;��sv�{��d����t�'>����2N2O]f�J����'�I�'��=O̝ML��&�T��8��=�ف�N��js�%IԝeO;��o߿k}����ۚ��8��3�{�$�Zu���>d���	��&~�m$���+�š�+'Xqd=O̜Me~�� ~#/�@'��#q��������<�y�>������;9�I��eMy̐Y:���p봓�<�`;d���6I��M�Y'M��k$�>H~�=ed����>C��Ny�\�~>9����|<�;���$����&�'�Y�2q+G��������w$N�����d����6�&�9�L��6ɮ�!Y'���쒤�!�s�_��?{���=����>�~�ʅd���<d�50�M��~>�!��$����'��8��hz}�:ɴ�^w6��O̝��i4�N�w	8�d�~>�U{�s���V���Z/�H(ou��B,����!���;F�_}!���r�uf��K���H����ݫ��t/B�9�43��gJ5���6���Հ���br駑N��el����|4�H�DԃO5�����a�y{r����}�W����s���z���������?��|�d�i8�l�0��I�����$�5<�:���/hx�x��̝d���{�x������<}����y߾�?{���Ͼ�6�8�O5I8��;�0I�?5��(O�$��J��P6��6�aa8��~5�C�$�f������4}�8�:�߻�;������ܿxw}ן}���=d�	����&�z��a:�2m�<���2k�`,��~��IR���8²m+'�)8��M����	�O���d>q'Y8����|޲�r��~�>w�������'�:oxu��m���<a�I�;p��Ğ�xs�̟ �]�Hu�;���:��y�T�&^0��|@��d��������31��[.�����}�߷u��?2z���2x���'P���x�L=���bVo�u�XOɮw&�q!���(q��kt�Rz��5��IĚ��$�Y'>yu�9����&s�y~޷���m�O�����ǉ��2u��5�OY<aĞ����L�C���Y&%a��a�I��}�ԜAHh�rz���%a�C�>H�.�fe���/���{�ݿW�{����'Ny�Wē�A�	��'FXu�x��<��'Ƽ���'�8���2��'�O���!����$��<�d�VC~��y�����%��]ݫ��o�~?|�G��r������{�I�Oud��u����Ԛf����u<a��Oۧ����:���d�CL�A��_�=C���׏��x~����pi~�� ~�J�:����p<a�O��{;`z��'߽�c'�I�Y?2q5�ǩ4�e�d��Oڰ�0��a�8���˔�˛���~�ߺy�X���i��a �/�m&��s�I'�y;�:�Ϭ'�~Ì�d��Ou�@����s̒�u������!YY��OL���ԩ�w>����^ܡ�3��1�����z�怱�8���ԭ�{;&�G�>�]Ӻ���)����iEY1��U�1��7�����d�8��rR���%���훙���i>#�T���{l�,��֫�y�j�ݦ��F���f��{�1T;�5h\Ȼ����e\;�$A'��1�I�[�8���ݗ��f X�-���+4C��.��hÎt�8:�j�T�m�N�g%�&��3n�^�i�vp�.[���4��G�p�}ջ�W.� ����� l�kU��e�Ƅ�	� �b�RO6���a�yS�
�'�$ڃL7o+*n5�����ʶ�cJʶ	�B;j���ҤsOq��.��
�Ӆ�.l|	����%&7Fbwa�$]����.��EJ�E���Ŕ�cA rT���^����9�"ƙ��IQ���86}��f���{[�"��-�f�����b�V�|���4Cz=��'��o��	��%C���c�0h�;j��L�5;Y�E��ꖗeb��݊'���:.h�U�]��m��ݶkCt��`��ܖ�T	����ic�^R&r�_W
J]L}Qѥ��!ט�x:��ԍϚ;����#�O2ue���
�S{O-����]o_kH�n��.��*V�ٸ2#���u|�*?w'}l;�ˈ�T�ŶI��uI�f	�=�`91�y�Y�I>���5ե�9;e=�Y
Bv֤�|��PPf��9l��pS�iV�4�2��A���v'�tzuvG�+Mn�ųՏC�bgr�+
W3�'��.7��<���2��5cz�mv�c�]�:��7t/�y߅< ㏣��([��aL�63nQ}���
Um�0��|!�5��	w���0�l	wY띔��E�y\��p�����{o@�ďM�N�Q�܃�M����Y;`�����;���+y�b&����:�*�y�ϫ�����������R���2�G��QͲ�v�9��HXc��8#��P��u���n���f+XͱI}��p=9�V���X���6V��F�����ɣo�|�b��7���N��g/�&�CvK����L���ϕ]���%��3i�I����.���d��m"U��a�@��WhK�}7�A|Ջ�a�;R6�	�@��O-�cx���f��i���X�/Z�%�^���W�֩���R����Q�z��K�n�0F�s��١;�g�e�ir[���-�rM%Ƶ}e�����;}k�9�u
�O<�\%>�w��pu,,6Uh׼9���*��e�����5nj�֛7�PH@w����q�F�����
}.R_�+�F��J����������(����[J���M���j\�;�S%}��j>(�o�՝\�C�R�C.�ޕ�u�?E���}M���iw��B�m]m��İ������2t�"�w =�R�{Iꃣ��f<�ccIL�ۥ�K𫿇�=x����iv.���Wτ�iî��Vׯ'a����BM��
pڀV",EQD�D�iX�S�JZ�%��Tq�ЫU-������j�+[++Uam�R�QFƖ6���ł�ۂڢR�iE��JS�L����+[V����V�ZU�J9aEr"![K\qKKs0Z�%j֕�EkY�ciF��TU�,J��Z�F�Q%�UҖ�*R���T�h�eJ(�kV,E*6�V)m*��J�s.4V����mJ �p��A
؉mV�-�nZ�L�.26�eh�J�mUUm�*V�-[YF�A,��Rm�l����*5��V2څ�������kTZ�[m����˕j�*�U-+(�խU�6D�����m�ZR�h����hU�
�[h�F�6˖\b��R��ER��QKDc-�LjDnR�,Z[J�-�-��*",QmZ�Dm�Kj\�1��)V��JD��m�)��±mPj�oc1ݮ��b��:��X���� e҃^Z%b�'@;�d��`�;Z��#�$.u�)��y!�A�KXS����e��d�o�������>I�9`��'R��ЛI�;��u�a:���ì�}a<�s�'��3��l���5�VN�?n��Y?'�}��+_�s/� ��3���}�`����\d���3�8��{��:���9�Xu��Y�;�������'Xyy�Y8��l����'��k��8�q�=�CX�5&���{����1���~�t�=J��M�S)�����)�'�q��XM2OΌ�C��J��{�"ì�}C����o]�ߩ8�����a��?}�ט;a�6	������މ��{$��M�������d��̇�ӌ*N��R!�N��La6������i$����:��l����N2u�~��?�D���~�Aty:������i��������'�ߘ^�x�I��N3�&���������%ABg�m
��)?ɴ�d�h0�M��~���L$?x
�?}��o���,G�'�������{�m�۶��ORNr��&�?$�|�:�d�&�;�Bm�d��I�,L��D~���Ɠ�П�*�`�=�R���lk�)���ޑ3重OLFI�g�2e;��{X���<�e��3��G_d��3�k}0)q»��$�X��~�/Wdi8�-N����D�A9^s�/]�x싘x�xo�$f�Jb��y�c���)R������+���G^�"Y5����ًg�����/v��1IY��*^#�;��i���NGfN���c9$z����Nu<,�������P�|6j\���jo1w7D+�)M���݀��;C��_���M��"��K�c���'�P�E���:��e�ɜ��K�:�"��VѼ�snjVq�z�>L���x�Ԇ��睊�9YŻ��5�9��>m;�?q�m#2�Xq�aP��r���KHwl��	���Js�ǟp���R�;kok��8�6^ྮG�Nk�|Ʈ7eL玎��ϓ�e^�koqy�BL��g��XT�l��Ϧm|m��l����+�b1�0�;V��H/�`��R�N[K(�E��]�W\(�������y̆�ӑ�q�Չ������b�K����+�i�'��=|61��r��K���i*��Nz����#�s<����=ߕ�1�O��{p*�l�Ԇ�H'����<�%5ײ7FS�I���8�X�v�,a��%��ܺ�%����CI5�~1��s27�+99���L��>�6݊��uq@�+��m��^�h{�U�WM�>�*�8�k��E�/���v��|S+lc8���@�!����KOw�]�{�G�>�sϒ�����51K�3����;��0;�fS�[k���Ju�� ]�}����Bř�n�Jw���Fs�;q��f��<��M�Թ��p���#�)��$�UӾ�x@7	�D=�$�v�v�탹���iK�>����p��T����߆�cs_����a��]Y&u��8���w+O�w�h׍j��D�4�u]=��?3���i��Wz����G�r�۾�Sǵ�us�X�k ތ�rk�S�{+tkϊ�=�.tBϯ �t#7�y��]��ڷ�� j�qU�><t���{��<�o��l����E�u�[���讞[� ����N���>�Ǳ��jSGN���oNZ��S��}6�)c��g����:������.����aͼ+#�V�5#�[�Rq�3�x^�s�w�˾����[ű�-��z\��^}^�^�g�q�+u�qGF���iNu����l>�<��붺.^�Ҳj�$.���B�.L��n��s�mǼ�C@��]f��[�q<ιϦ���o�������L�O|�����(��=�I���O�����ش�5ԬuJZ��3���Ƥ��z�{!��؉���n�]9Ra=��yqO���3���oo�v�S�3�\��c�F������~i��A{F鳗��uqb�s�X�r.�cl@��}�}�.�{z䤳Y�?�}֜逸���TNۇj�n"�e �ʥ�jE
���]Q6���W�����:1���-���tu�t�`���U;:n�{�Ͻ���d��̚�T����O�)�T���i#����v�ּq�+�t��d�C��Uyt~��'X9�K޻5]�{}*����r(�y����h�5�3�6�Og���������w�Q��m�}�]�K�K�6�Jg�)�v�V�	��j�'`c;!v��T��k*&�y������r��%h�.m���x��U�:��V����6oU�r��y�&}�ek~���=m����&��xֱ��>閂�iJ>g^gc����nv����%X[��O:N�y�b�_��<9]%Nƫ���R/*�YE�8��V�d;���*�9:�zAL�2��n�.��O��K�`��i���Cb�'��g�4W�r�U�X$\s��!��_ ��}֟�7�m������b�I.	0-b�	^4K��.ۮ��/�.Uc�+����:��]=/Y�ڷ�$�z��Q]ja�� �_c|:>���}����|�����%m�yo*�eV��̣m}�B֝�Z���� t;�{ �]�oy0��a��2���3�<�g��gnI��+}�X���@M��C�O��Y�;�Q��·����/����;�*f����YM'Y�����xԦ�tw�9����=XRx"([��e3s3ؼ,��/og��/���O��c8Ho�G1��GNFH��t��	�ۄ���euo,}��K��_�I`V�W�ÌHxʗQ·��]8��XT|eozWl]�)��Y�>2O�k�6������<iJ��k�lr��2�Wwu[m[������x�_��~��ѝ�ˋ8�/�Z;Pn,�n�n8���+�;e;��wL;A����p�~ܛ�%W@��U E����2z��.玎q�d���L���	�E�|���֜'��kr,�ɺ��5L�pE�,�<"�e=�m���PP���=�=2�|�G�:������e�r[l+3}ua�?SkH������m��ێ	�&�ڡt�����M�l�մ���'B�hLP��W�*k���֪$$���k񯌻�:I C�������z:����1��d���)~�V�IPK��o�p�C΋��U)��֮�p��0mʾ������v���}w��Z.I��9�a骕�<�oQ}S�۴�v�,B&���C;6OeݏlF�I��~�ݐ��o�_t�'gxD5�u)ŷ��U6|;N��g�J<���i������M��g���hZf��]J��ѕ�]<��Az=si�-м�Ǆ�L@le�z��cK����[��W���p��m�,S8��׊����Տ�&�R�[ֻ�?;�z�ef�J5�f}���F����^j�/L���2�J�g^ΰxJ���ܔVl���y�F8��j��lfV�)_s%\#�a�G��¶�w��PP��;�8>�rӗ8����TouW)^��Ǿ{��`+2��;^�jq�/X�����1!��w �eej!�_��6l��t�v��[��T���N��`�y��}]���� �X�)D�r.��k]"ǽ�z�ڲ'�Q�땽��D�t�V}�eu�T�+v�6�7��c�tz�(X�f�Rp���[��@��YBmNz/��5OѾ�;� ����Ή��6����=�����a��Vv��v��;<6�W͝���Bj�x�31�v�ۤT���	ϲq�gh:;@��Gc��<k�u^��w�-"��Ú��y��x��sV����g�gRS�6݊��ޑo
�¥֬�[���s�]�/!���DC9-s_�z9���)���C��"���*(3H��~΁�Ȝ�
HG=�-���~
K�|�wze������ig�F�+z@���rX��YY�As꿩�f��<�L�>�Ξ��Xz�^o�=]n�3��kD�ۘ%d�<p'���h_�Ѧ��1%H^�����.W{�捷�)�5L[��XM��/��;)=�]\{�k��(-g�A�{wr4u��w3��չl[�����I�݇虫��v�&i�~k{Y�x�nTŇ;&�����ӆ}�P���Վ'��M�X�u�����SLW����筄��,7zf>Ze�Y9aOǥ�i�ڨ�eN���X�j���7܃�k��	�Q=(�OTy���YDC�����Ƿ�ej��C^�rp�-tfRw�%�)��+�嗭_��YC��k�@�b��p?�� �}���کXϻ�̬�9.���q[�׳*�JܪN1�{BE�����8T7��n{�|;�l�����,�52�;���t�d�[�ds7�7�6�\(Z<��p����ºךH[�l�����[�=�v߼cE��۞�&ڞ���7��v�-m�Ec������/�7�%r�HQ�_�:]��R��p9Ө8�*���{���>1����ozI���������>2�hdlm'R�*_��tcy4"w�,+�7"�j��[~[G�z_�G|N��n<��63�̛�������'2~�O�;�����sT��G`��n0Pd��:��]��s�&���Q�����.�����<�,ob�q�n��҈[�
�_�t��.���}��K�7��]O�19{5'Џk]>q�����:�<��;�\��{B�&�+�?a� �	}\Z%X��}=�H�ӧͭ�[f��v`��D%e�t�F��X�����v�X�72�
�[h_F����;�j�{�Rʼ�����_�m(oJ���ptג�}�M���t�Ò0`�yci�mNŹ��k�}��$����| �]�t��9��Ӟ)y���K�&��;��Ɠ�Ug��&��]���^�7�k�FW���Zڎ\|"����$�K�o	��n�y��x=�k��O\��a�܋���xt���u�9MVWE�c�xO����M8�{]�J����ܫee.��^��{���.��~>����<�:.��W��1�3��ʣ��ZӸ�ֽ���\�gt��bv^����?>}�lsǧ8��bx�1��Vey�Ï;nC�$���5�n���<|�n�YS��i��cKbݵ�H����ۓ^^�K�����\h��=�3�,'/��q��9^�dK��n<���۱ڳ����f��Z�t�^��88{�ƥM���d��U�J�2A=xsX��gl�C��@�k���Kyl�8lc�%}�y���E�+UMY)k����!��B�Wrv����+���m�,MZ�Ц�7��M��#��]f]F!C]H�bڽβڬ&�⚤i�i7�ԁ�|҂�Q�h�ԝ�C�'}J���x���C��9�C5g&�.�kE-�}R�p5w:�usbo磌�[�����G|ϟ�{����3��K^V����63��DT����=�Ƴ��;��7;�'�û&��cn�V6@9���G���udz��}St��yݦ�ݔ�Y7����8~q�}������r��i֍�;�]�����?<�d����#B���7ɑ�t=�)���������������A�!�7�=������VԹ.冤��ƇS�WZ��/��4�uS�͋����o�.<�*�c��v�*ǰN�,[bvɾ�e����}[È{/o]�x�ö�xt���e��Tt�˲�OH:ZɩO�mcj�[����n�v�~�%q�x�Y�x��&�W�f��F|�]ы��OP�u��G|;OQގ�Ȇ]O.��H)�X��8�v���}+�E��z:-��gu���7��	w:C�p�_�,���C4L@�C��;��]�[��qtGq���Q܆�v�C�-��hpg+*�L�ǤV�V-��7�Fk�u�Z5VZO�5N���8&��;:P��=���(�)I�]Yke���-�&1����9(�t���5�3r�N��Z+)�Q�逹�<3���f���r=5}��e��vd��d���*��ΛO�C*����ڱ���e������ڢ�s*l�guL�ע�N��x�]�7��չ�ҙc
�����i�ιʒl |�2��f𭵃�|�R,1���U���Jov;�KċN�T�M� V�>V�xN�.NE��������;f��-ז�������a�©���Uۈ9aZ����'5v�ACٓM�:f�)��w�ԋ��.��(�3��A�nՒ�*�-�l^-��i5c��n�Z9��k&k��b|e�<��δ�g}yt�q:�e���[N�]W�]Z�ЛO3�ɶ1�4<Z�5[����]��RȜȭU�E�C<C����T�Z��n�M�9J�n��+���ES�N!q���To ��t�+��:��Uu[˜qc��,���P�ruy�9����u�d3J���f�ü��;ޱ�=����,؇B폫�kc���f<0ofb䫱n%��M�����١�S�Zk�@r�Q���D̤k��+��s�J� �+���4:������������CT7/7sβ��=�j��9!����g8���������X�iг��ǳs����ꈓ$���[�vӉM�
�u.�=*�Ym���v�4p�$�G�D���n�^o�Pf��|�77U��aJ�󖉩��qJ��$�tNW�m�4�n_u��=�H�Λb2� ��h�ϫ)Lj�-��fk���W֍�]�tQ��oo-���~�1����V��*O!�r��}�fe�t7���h��8֠��+��S�Iю�Rb�'c'mL��N���k��V����͐�:=��E�"�]mֆ'TR�����8_Tlm��og��#*IE�Z���h�þ�/�6�f��$��1*����@���!La��M�Ŕ���ǺXd�b"efc�\���'(��ޒ�:W&7HMܾ [F:Ym`Lq�t�a7��Y�4�1�B��C�KO�J�ݨ:���m'F�
1k��q먇a��׶����8���y�,��*X�lANv^T���K�f�݅U���k"�Kq:Er��U�F�����/ @����%j����l����Z�ڽ�f��Tb��J-�޾}�W��);\�}	��
�^IT��g����i�p1�^<Z�n�媄k�f �����=N�U�a5�Z�[]G'<�|e�{RwϷ#FhR]Q��_:7u�l��诨�l�g�y�˜��%�ݟdf���	�4��� 	��b��5F\��+h�Rڶ�յJ1�jU������eKmm�V��J.f8�iZ%j[*�m����Z��eT�D��Un[p0�ԭ�jT���Rۖ�ȱ��������F��0F(bjVW�(�91-,e+ae�(�E�Q*���R�j��Lb��2�e��-PUm��iV���eBګ-*Ɍ�i�EYR�j�j�X�d��*��C��-E��8�,Q��3)�E���h�jPZ�2�����1�0P̦ZT#K�EƪRйb��(dJ[XVEij
��Q���j&Z�Z�Ƞ��3(
ĶU`�Z� �
����#h(V�j��4�A�,[l��
�iX֢Q(�UE*T��`ۖ��QJ�PR�Z"�B�KZ�-���s1E�X�b�r�����5�>�~�i�ϻ�My�7�����G ��v��}2eN׭,tn���eշ�q�k{�I�gp(n�c��q�+�����Š��^�1���/={</z��6�\pm�8���ֶ��y�3㛾ͼ_\�D�F��;�'�/��Ҿ��c�d�倜�j��a�v�sT���Ejv䥽�[*���vfB��yݩ�_]1z#��nZr�WO�v�[=�|t7"K��=nv���j��)�P�=z�|/���1 ��uൽҥ�6Ԗ�!ƵT���
Ώ�������rUs�g���u&�}b5]���K��\Bs�8wL��-�U��)G��3k�-a̗��y�y^��L��ey���L�&�J}�0m��R�x�T��^X�b�>�������}�vE������{˫}�g�q)�hHd�t@9�W���KsX�����ï飯��C:�%����\��d-g�.�WOhf�s4��t��2wx��p�n�=l��Z+7���"�U��n�I���E�Pu5�:k�1}���륹o�E�gfa�¨h29&�Zk�梧%Kjv�x-���7��r�i<�C[��I�y�-����t�|�<[�෭L:��u�d�U_U}_ͯFT�+^~�e<��_\ۘ%d�<q=��b�?Xo�a�����(w���t�`s#ȩ������2���_p���%��/2������ӵ"<b�̝��oc��Lu�Sѕ�;�<Ajd��e�:iI���Wu�s��%�<b���kzq��_?N瞜����<��L^e{^���
Wir�q��Ь8𫏫N�ju>���q�D�����u�Q���V�vRBL��,ϼ�ʣ��+��'Rݕi.c>�S)�淦�w��Cds��<_��xӰ�/Ɣ�3�1��j��T+u�sg�����z�`N_�l�M}5�����%�!o<�g���I�<}�St������ʔ�oVSA��J9��C�q�U��5x�X��B:z!�v�{���ΧD�6��1!�&��t�^��3z[�Y���3D]�G�Ȱ}m��ہ?To�����D�uwՖ�cg�!�*�v���:y�����iU�-��׺ŖeI���1U�԰����b��m��՜֜�%�TT�ò��Ä_·��6�^�a�K6��yݹց{o>�.��k�W�����֫w��������_����ܺ����r{�	@\�u�Ny���䦍�͎��5{ܢ>|���Gh��k���z{/=Ѫx���9=�fn5K5P7����]�M%{��O�y��%��3�}�:nq{�75�${}v0a��������pzeSq�P��0�c4�
�k|�OTAG��/b
��7���o3�SBv���Ɵ�"�ΣW&�L�o �8\ӗ�Z\�J�o�FWsԥ�:���욛��z�[Qˏ���
�bI�.���<A��淤�9�B	��yW��/xKkg�I/\�,8��N�N��n���6JWX��],D�3w�a���Qk���kzx_��W�yY~�YҲ�ͤ��~�5SA��_�`ǺT��̬�㺬*�Ӹ��iKW��?+�/7*Y��#�s�9�A�bkG��<�e}T[��ܭ��A�?H0�#�}Ƿ2�V]
�-�U�����ç2�6��[S����%�yʘ�7Z�
T��%�F*çcLK�}I�<���M�
������Ǜv��`�`��Jۗă��MMƼ ��'��yϱs3��_05���}_}U_D��H4�+�/�S��\��0�����Hy���'�OvK�5��:��+�����rӘ�Tq��Յ'�ip���{^>�NWm9�;P/V�]�_�/Db�����ӳ����X��M� �c����5ys�N�@;R�Χ^l���.����b���jlu<5�Sl�Ln՝��!����r��gX�/���NJǆ;\9�X� s�VI�2q�ghW!�ᣩ|3���ǭk/�5[{u1z�}�����s�o;5q��B6�إ��,Q�)Ԃ�z���/+w�yG�����$DBts;M�p��fS4�������xv-k�\����>O:����4c}��I�)y�"��K�˒덚���\^�l�t֭�s���3Ӫ����s뱭��.<Wx;Wo;X�<��@c���ov�G�{�'J��	'B���΢�cM3x7x1�H:b]�6;��]�k˩��,ע�x��s݊�eJqz�,Y���aQ�[��º}����{[�	S��ܜ�脠/\�wN�V��]�����d���4C�{���P�7��UW�W�l�ȷވs�tޯ��Q��qe�^��͓�tǶ"+GHӒ�s醱�k)�9��9�����K����Wyo��YB�M�mf:��Y��cbcz�>�l�5�{��!zzc�8vw��3�ek����ᔮ�ُ�����O�/��C�p�ҽe���5�o�g�A���]^y�`�������Z�vc�<_aY��tkp��-N1����>>��4���V�{���]�z�?��F�l�kq̯9����=�b��䡩�{+	��E^SAe��ڎ�s�_B�>'��M����e��'� Ӟ��y�+2��;�z��}����p�֪�9{�h��c��:+�}��t4kg��?`۪F;��k�;B���`;d��.�ҡ\1Jq*d��9�û&�v6�s�5䛳�.z,�>�O;Nc��}D��}=�����U��^̧��A�#Xv�vZ��1p;���;��='7��,gCݔ{"�u�w6ze�B��..����Y�,�Q�A2D��%u�va�-�)+��=c.��=��uA��F�[#=Y״����}��U�\��.���fܹty����l;���'fHX�w�6�����:�u��3x@��
��v�:�o>	��.vp�:��<����1r۶�7\�*��J>z�ˡ�B�4���:P����nk���F.7w2��ڭ��J��]1�u�fK�;!k<h.�V)�}�<����0_����_�V�s؛]�K���9/�K�,Od�5�4�ʱM՚�n��-vH�<Җ�딷�2�1��z�c��/�&�ʖ(p�.^���c�U���ǡ��w."�s�{�;���w�&:��}=A�=Y���fL�r�U�]�]���y����<91��d;ӆ}�P��S����ߢP�C�>W�o��v����H;)��a�u�d{��w��c�NJ�#B��M�}��{��{���Z�1!{�g��G�n:4�d��k��,�P�p&�z�˦`±�����3J,_@�V(L���&��Bt���m�g4r
F!��;dK�z�wݘt�u������V.��9�ge��*�S��N�}������Wnl}5��j����}UU��77}�����d��N�5K�9��ºךH[�l̯43�&�'77w�)�یj�Kgw6ܿ���d{5�����_w�;��m+{��f:Vؕ�͆.���d��ZQ�w:5��=~���Vtv��uXT=��s"���|��פ��9���H3�*_�'J{ɡ4��vevy�*�3&H1��Y����׵*�6ly䛰F.v���ic����87c��+q�:ó��ttqc>:�{�w��ѠˈA'r��W2��{�Ş7/���kg�>6Y�8~q�B%Բ�
���C�nqk�Bͯp��>̊����������S���-gUC�otF��ϫ�#h'�oʳ�<���c��} ��1��5��)y���ɝ^�o�)�;<R�G��R��lkׁ��Y�W[�����z��9̏T��
u��y�;�@]��%�A��x�]�X��9r7�_xn�F�'��?)ڲ�R��^�W<�K�Y��s����
�w9�wa{ڂ<���o�[���c=)3�^(P��8]����U�l�1;a���f�.�(p:8�	7�nhU�U�ZQ�ĝ�������5l�G������� y1zl���g����ų�zIx尻w�/������2i�i�A���n��E�Y�C�C��i5���Nu�c<�e�
^DC�6V�?<Q��;��]�}����,ڝm�a��H]YRP�Y�W2���z��(�i�CVq�d�f>���Ξ��������Y�W��z�9�*�^Չ3��UA^[���IH��06���L���|})}�+g��/AU�:U�<�.;v�5Ҫ�M�
0ڊ���_�ɛ/7���V��4��p�"۰�ϩ����z����^z���C�m��ki\s6���y5�+��j�\~�:�K�"��ߗi��R���⎁�}����@5���Y�G��SV�h:�iA��S�|)Ď1R%�D��#���\�N��m��ç�ӛL�f���P̬��XZx1Z�4UgJ�=NfW�����a�훕~�=wM��v ��d��Q�'[����k&R=r�65��י"��թ�!��umu�$���C%q��*meL�ib#�Uм�㛖������]|/�{�*�4�^}��<(���ɢq�}G���y�R[{�X��A��V�J��hJՇ]t��Xt(��D.�L���[};^k���=��V����׊t�� � �Y��S����
�c�M�fp2$2s�FZ��Ε���֏�C�(�(�Y����Q�f?F���,���+���MF,9˅'������0v,�Yw�?X��zOc�� �H�:^J���E�"���a�e��R��LT��d�X�RТ[�B_�WX�� �y�j	������:R-+�P��w_�����;G�`-��*e��
��h��cs����:��<�&��c�B%'�q�k8��r��)��3Mxn�=lwqt���Kь]=�7��l�h�pS�H�D3݄�v4T�E��T����k��t��Q���E�����df��K�܀ѿ���Hi�X:��	�<4k�������(Ṁ��n��ح��x���
�E��4��P����cK"�ή�|tnm�<��:Ӣ+W+�lx�K���G�㞃��a��o�a7<�4�ҽrg|�K�$ ��M����-`��Mk��8Mk���MyX.y�p�|D���{�]l|<|����!U�!���^Mܰۮ&�qޏf�y��*)����f�T���[eM9c��s��{�*u+F�l)M���
�2�f�B�p_z�� �ir��s������:�/&gQ��gQ]���^�Y���c`��{�{BU�%�)�롰޹ǫ��[�U�W��~u��g��b�����B�ۃ�R�-�z�1:��Z�z����W(x�˵�Aw�t����;N�/���3���[�ͦwe��j��[h�/V����X��<�Nq|�^3ԧl�j:��e��̷w9C=��q�wL�GO-5�T�O	ʬ*/��:C���ㅭv8�6�X�Q���ъo�ل�x������hw`���tWy��d����T��F-��؉���e:���-}���q�� t͝�=?{յ�K9�=���Jk�P[�j���H���"�	��wf)Bb�=�B��d�7%�l,�����0]�e'x]$�]2'o��#^�3,w��=*�u���;tV):u/z#���O>�	��hS�@��k���t]yv�_�딜]��=B������4��/!��ov�O�Umi�P�#�eù����$���2~Pm�.�Ҡ�'.]o�;�wY�>��΋\�`��ȃ�WlgGJ퉗f�?Fp�xJ=�l���'�`�Zq'38r�B�޺����3M(y����IY7#�Fn��hG�,�:F�*�g�'J�Z�C�`���qC�o�pK��:����s'iٺ6�ml�4A�k;6ʮ�[���؜�us[wՍ���ØYۥN΁�G�Ű����׆_��r�'+yř��WMjw��H��N��x�m����˲3��t�s�][���ɠY\��BA�ֲ�u���E�O��q2��V�qU�S[��{�.]$��k��P4��:)⚋8��d���u�$i*���F�(��p>�;:�j����.��\���w��j��y.y�T/sl�g'�r�̢�(9a�m�O�F`{ˠn����Ÿ���"�B���Z�
pz��nW��}�o_S�9-ɡf
��j� ��:���%�QP���"��Y.�Ǻ�۸yh���d�#��n�dR�K톻�y����@>Z�r��:���	z�Ij^Iq萅nW-Z��y�t��V㮮�j��t�+�:;�(�b�S�����;T��]�fVv�\B�*�h��3��cV��l�\/5U/:�X�*Zg�i�4��&*}s@x�,��hS��9�[�2�C�X�n|N���;v+bc��Q�ow�ws&>�R�]���^<yl�ޑ>��^YN�XX�8�.f�uoA��wQ��x��Su�5͕}P�;/�Z��LU�ge�H2�3-&��O'!g^�f̛Oi�:a#��>6��D���^Vh�|(�Z��w�����3&Z�z�؛J���{���7]����}\+e�����a�{r�4��[�
Y�k=/ ���Q�7*�.�"�q�Φl�]}�%ɛ�4XȢ(��Y�[��a��c2�R�SƷ7:�����X�o���K!DV��H����՞�jP�1����]�g�n���.��JXN�j�2���SHG6�A��RYYӍ�����5J��u� H7�,��2Q��mJƆ������Y[D�}�K��w
�Ac;�%���6������@/��g�oV�RÙ��n_P(��GիzF�7ˋ�ô�jh#M5ݐ&-:��Ц­vŬ�A��]�w��G�Ă^nS��j�F>���/#.�W;J��/�q��J�W��x�.LM#.�u�Z�,�����7�EP��T�>f����&V���
H��ow�.�������d.�c�5S'8\���9B�r��LĔ�펓^Ts>�`�n�]80 ��J�%$�u��1ʃ��7d]vwu��V�l�ռ�.�+9o#״�Ns8����0���Va	��7�u�7:Nk�e:�R=�8ү��c�[��^�J��AC1CD�Z���Պ�U��:,X�pWχWh����J���oB�o)}]ƥ��t�!�Quӓ�soF���=��׮cם�c���D��Z�7���n�lٟ��_c
�j�����Ym���mF��j�UZYmZ[��Tb�e�m"��(QYF")D������TD+J"��ʀ�*��X�����,D���VU`���ab��DTfZ�����i�r�Thڂʖ"²Q"ʪ�V�)LlX�iJ���`70�TX1W-���XX�����[��VX*�Q�����5�j�6�-jZ(���--։l��
�őAUk%b�E�kE(5���E-mF�b���YE�V�Z�[" �D�i�imj��mQKh�)[TJʖѶƈ��H5l�ª�TV�V+Yej��҈��B�mmX����ƴR�(QcmX���J��F
�
��[J��Bڰ�ʢ��b�j�D�U�m���6�[V`�Kh�"T�"��
V��b���ՕFV1Q�(4�D�Y[V�ZTX�"��YX1D���S�<�F�A3/�1ۨ$���t�*j�x��ǯ(-&1%�&��n�����D�bW��z�Q��k-��h�� �}�vh�w%���}Ku�u�f�3�o_E�s�)+��R]�u�-r�p�;�+�`�����9jv{q遫��=`Q�eP��r�TR��u�g�ޕ�k��~����n�L>��uXޮ�?_�J59X�p�~���ʇ�ӣ�R�&8*r���z���{c)/Vv^�DD't��4��נ
���O�U�76����H��ՊPӠb�����/��I���{QC+Ď�]��wW��8ρRev������E�f�'�9�,��#8,�@��N�q�h��*�Y���fe;����/T�P����K9�2�j�7q�j3�0�����f�j�V�J�b�h�
�8�;���'.j�L�yv��Q�k{s��* �	��/x�e]���w|]t�V�I�:&B��J1_�N�0[�m�knŝ�-��O�����Y�ꠗ����i����ɘm:�#�lYS}��D�5ݷN��N�9볶ZĆA�Xpl�g�����K�`�Z�Aq{޷��S�5#��w��b�GpT������m�=*:�1����D��C>ڐ���쫜�S�T8�t�쮎���ś�@o�Mݶ�x9|�����͝���c��0=�&��36��)�U�(-�ej�}us��1���L�~�+�x��|>����%Ӄ�i��ky�h��{���
�O=��L���("_��ϨP�wȅ��f�Þ���i3�\�����ॏ�y�uE0���&�� �E�u]/����*�=<�?
������
.��Pmd���=@�5���/<�����c�1p�.8&
��6��}^�1H��[PP��Rk]Ǯ�s��4�Y��=0?Ev<p9Fֆ��UdW)3u�xr'j����~[Pf����j.6�km=޵��+C^��ɩ=��JCpy�? ���~N��-u��C�C��i2��y�
Y�Q��s7->8���=}�����q���m��9�I�eIB�dU�t/]��AKEA����#�z�����P�-��Z�ѿ���p1=K��e0R j�o����\��M{���p���B���}���Rӕ��%����徹R�yL :�b�;M�C8b�YX�z
��gR�u��]�sθ�3�,�`ء~Nk�_.�}�eoނm�����*��&~ѩ�b��f�:��=��ؗ	�E�|�o9�<OkqZb�ɤS7!Y�gg���U�-����S�s:V�j���S}!yŬ�Q*A�zs�gl󇫹񌔶�a�#8r�%�ݧ��ݧ���[	ط�9Mo��y��W~��M�=;����v���x*��]���+J�2�c8T���0��ҙ���*�glAs�b�Х�پ�8��P^u��VZ��#H����<�L�+egx+�=�5������E�q�V��t�>�Cx�t���i��֥�b�Z���6I���̘���o��V����j4�¸��k�e��ƵG�o�2�'2���]���L��\Dwah�z�*	��q�b�z|ΓXnB�x��=�"B���k�+89l�Kdhy�]������v�v�ͣ�����!k�W"�vz���XR�W���tW0���=Y��荞��4�;��z�u(��T�k>����>L�ڞ.iK�/�����g��������o�Q��v,�PvZK�E��u�p��u����v�b�k���`֓��ʞ�ն��dYg0l�̃W�4�"PB0��B��k��\e��}=����A����=!�[<�W��#I�}Kި;��N(^J���=GڮHW�\򗬑��3�&��g��pV���������jgHB��e�:���_^�o:)6�j�Cԣ��c� ��b�K'�&q"W�Jˆ|My��A|e8�2���'Z0������.���z��6Ρ/J�������#hQR�7f?�~ڮ��y��\��;Cl��� > +�����5�?���g��ҙ�z`���4v(X6$4�.P��F&�z�uN���<*7+��W��U˩k�G=zS��B(���P����'1��谳�>�O:�{F&=or��N�N�W���!���6�|V�ߏc>�B��J���?z�6J���K�ǳr��M��'����ٷMf�&���m5��sσ���-��[��V|��q�x��d�O٤_uk(E]����S��}'�О=�2kTD�:�ڸ ��zt��z��6�ߋ�6ҏ/�g�3���1�s��ɟwՖ�-�Qm-�,)C��{(G!غ�1SgTپsɽ6��%��S1z�3���������8׏`yl�
�G������˫�\�vN��󳚸*EԂ�<�KG���f��Ī�	Ƈl�GK'�"�%�ko�8L�b�l�@���Ip����Mk�|8N>Ñ�7����9c�[|�c�w��S�@��1DO��ڤ�F��şPL��1J�)�;k~..8>
dEz0�Y�����o0c�M�Lm�-�ZAN=���w��V�=ݫ�l�b������^�zNӏ��u�����"r].�˫�O�w��Y#����[&�QO��h��5V����=l�e�Tڙ/`sM
����[|o�ue�> �W���9A�������zՑԙ$6����D���yB��޶��K�kFd�����"�Ks�W�S��98��.��O\Ň��f��<&�޸�7�B�g�S[��:s��Y�D/��ߔ̅©�a�FL�w'��l$����^��;յU�A�VH"�}j�ٍ]˱d��ԉEp}��Q�+"��q�%v�˳
���a���\��6hg���xpd��C�e�7�{�ґ/�|Uo=��ޣ�ȵ�W���]�S��K��0�l��Fϴ�OpbmH�9w�c�Uk>�Z��(*�\Rº�R�#�M����z�.1�^��,O*I�߇��|���߶��#Uq�]���S�mBz���Ŝ���wz�$w�2���{U�Ͱ��JE��ՙ�Klb���{������ރWw�B}�|:��b?Aa]�K��nf{2!�V`Lt���"�L�F��%�qBԕc���]�8x�Qgۘ��w1i��Փ]�7���g� �5B� ��O���<Хq�αJO��������x�zt�p/q��ͦ=}P炱&��p�)VH����߽���ظ�N�H�c�ڱ�� ��V��En:�7{������#(~�?y9��QD	ʵ;c^�e��F<�ǖ�p��u��Vw着��k>�rR�=��Um�Ϫ��^t/����QeBV��|�5w&G���\�ш�p�QNl�y�U���g�J&��k~��3>�	V1�$��d+�(�$�m߽�N�S��Tt=���O߿���:�%�'W��\[��ӝ��_�טpY�^C#�&�>��i�'9���ho+3`��>�hqDiϒ�$�Qű޷�ϞS���$���4C�����ڳ�%�Nƽ�Os��:]2��.�"�� 4�$�4+Y��2.�d*��e\�p�&N�ڹ�����B���:��{�E�lva�h��]���o�k�'��Q&ΰ�ڬf�3��c[����A�*�▴p�p񒶦:����gM�U|� �U/��Z�9��~k]��Ր�}��Y�uTV����:�'����鳋�}ވs ��w]���A=h��|��1yh��c��l9_٬��~ޙ~���A`[����'tB�"�^��}��N~èو[K*J5�,GQ�(f��^V{��%��b����y6�*J�
Go�b9\��u��!�'W�
ސ�o���qU�׼w�]�{ȣH�Wb�4��fr�<�ǽ�D*�J}�(��v�9�2㕽RZ:d�I�L>*�WY23�wT�����Aws�EN��}���y�2?AO�{W�뢭��i�'~s��89C��Bxw�y��ڢ�3z�����w[7���w~B	��r��n(<gL��\�c�����"�Ŕ�H,���Q3�rwc�ϋ��p�J�s�:��v�Z��X؄�^:����T;��%>��;��94?f�q*3����Zx5�O�G'�-�U�C6eW)P�^�wP�\����-���׽~/T���|`���%a��8T} sizxO ��-���ڹx��׎5ſt8��v�����ܰ^u����_iF�I��-�S�F�8�A��}u��Us��:Q^|+m(ݒ+����{L��3ZԵ��\����?rM5�^v�J��]Y�#�ڦ���R��S3}�	�K�u�/Fi��e#�.��b�x�]\P՞C�(��g�
�b��a5������=�ό�j�����T�0a�Е2�\j�4m��������X�*H#��ԃ]�<��KAw�_��e7G��
8�>��ab���{�N�4=Xy��RF9m�wSit+�D�f��ܜ�z!��z�w�jX������-I�����vLQ<c8�şH�^R9�s�7K��Է=��'5I�)dR��` �qk@��r�3v��9��F����^a���}�7�{�o3����SO㶐;�4���f5�#s����S�T�u�
�~/ϭeoM_^%���%>��x���
8-�œ�Y�ĺ\�9��5޺:z}|��E����=W�j�}=����2�~j�0���*(!�Hh�k��\e�����ov*�8K��%;LB����r�
Eϥ[D��$C��!��]<�j���W���ˁY���9�F㷨A���߹�#3�邕���b(X7!��gT;f�3e����i�5өܩe��Q�J٬���6�U������!�k�9'�P����u!u!�E��5fts�v�F{4��f�O��<Q�2��`���҄�hVt���g�ޚ���&�&7U�G�軖����Lk�V&���vӥ���\2�������"9ޠ��}ES��6�IҮ��3�R�̍�/vl圼S�[�8�4'�}�v#ʮ��;/�:vۻ^���)���
����ܔܶfS��y��0��&}Ֆ�7�f�,���z��dt���]|���Nc��t5k�C�{��\��a��e�H���w�+E�q	��,���,ŗ�ƬL���u	���sj��U+�����g����J�z���^0�DͬX���T��Vy;�����^v8gws�²Ф�º�~�}�,fo��CS��N�*�v��
��3,;��|���^�x�5�w���%?Yow���U�ۨ����\�A��V(G#4К�1M��0�o�SS��J�hd�C��R��rM�6ʯn�|��;y��pp��"ڪfu�^��Xg����&��c��w.�c^��i\�pt}�U�>pX�Xvhm���E�����f_y��*X�C�s��1��m�]P<��_w�I�~\y���c��xbj�h��;�\�J���^P�gz�Q�v&Y&�����W�tGj���_�L�8���&g���1a�C��B�r^=�^��>
=-�w���k�R,�M����Xo�L�_�Umi��z�LX_ T�s�����³!F�f�R9�n�i�77$[%(�yأ��ȃ��+� �xD!�����zߙ�^�G�a��)@���Rg}uQ3�yf�/���{��
J�S"���	������囓���p�'���S�4?�7�И}�j�8Ao�R���gګY����lv���8el���P|��E�@y�	�
���M�n6nKX�/Sw���H����I������R���Vo����J���9�pt�k�p�{�y8��~�kR�������-kSL|���/����G]�U�[i+x���\{���)�;A��[��������|������~�A{�0�lV��asq����:�Ub�����|9nx�/�V7t��[)�M�g�K�c���>�N滄�c&_i^kڶ��ѵ�H�Rz�*X�M��F�fF���|�6��Ը�V���e��u�8�g�ғ+�ʳ�,�:l0kt^�5-�C������YPo�mpӛR����^�x�Q`���N�-<a~Nk�F���Alc?y���w\�����;�X�E�䶓�T�J�x��XB�<�`U^s&���HK[o�[�OmK��?i�CTkN�Q<��m`��3/����&��
�F& ә�s��ܴ���sl���`�sܾ��*?U�H-	y&��ϩW��fϩ܉D��C9��f�m��S�(�d��7欹Ɵ,�a�֨�4�$�'x������(h�ZtAqc��E�z?`��k��E�R�3C�;�2�U(;W2��%�P<D��@��ǳ�T��j�(y�<�:1�������S)
�r4�mE0���&,	��� +��JZڬיmn`^+�G�W�YI�x����L�}��pQ�uxM,���5dT�[f۴�z��j���7�CP�Y�=3xv�E�W��Yw\�Au���c4ͺ:fSvŖ���9ٛ[LJ=�6G�V`�x�|���s��ޚG
����t�� �r��p� c���n�Yì���r�k�Z�1�ib�8�͘��ʊb
�	�Kj��3Pzݽ�V�X6��mv�
("YZ�@�C�Wb50vmJ�E\y��t4^E��8-9|��E��3��w�&_k�`=�`�9����du[��/o�e9�3�H�;�� �{Qr95R�!�s����l�������N���㸴g4�=N�[}�wYv�a�s�p�c"��҃0�n��'�kc5:en���W+���KJ�;��0�����4�G� tݽ�bT��h���U��k����º��ֈ�` PJ��3o��g�����"���:������T�z��b��=�Sׂ��Xv��|�3�EE��#<��p';s��x�!�a�į�2C1K��V�h@P|d�0��ɓ��i�"˩}Y�-���k�k�}5t�Q=L��Zj;ʴ�Ѿ��o�V]���[ksm0X�V�ݾ�or�G����2�uQ�6����P]uԅ�`nl"�r��&-�Y)�\���+l�I����lw5���J�v.���2l��X��ub��y�I]&aAZbDiv�ȕNc
s��S6�����WҰ�srN���:�!D�[2�3e�}��Bl}u�-ftq}y���q��'ض+�*���g��]�#B� �
�/�5���C݈q士.:Ŷ��u}����1���y�1Ė��p�o_ ���ҩ�/m����p��7k;��Cň˰+��75���S=�	�,�u.���͸ U8�nR0�&���;�hYOU�rܧ[6$f�b�:I�yK�2r��ۘ-l!�r����"�R/g\_[�:�ǚt]����1�5�SZ���T#ݼ*lTÌ�ݩn�%�m����Ϝ�Ǧ�CWq���
�n��2���F�e���zV�K�2��o��\;M�W��`/���6�솹'{��u�kY�d�57]��c��3���3QnQMP:m�RVL�ݹx�jJK镗9V�hnKF�g9M�E�ۜD��4ϳ�3s\J�[�ݱy:e�JhҏjTVm��s����"��%�N�*S���{���
'[��%��8e*ۧ����SJ��C�Y�i��.�C�y�(� az[[+�:��1�?w�Syu	�[󄹷-<�r��k37J@J]H�nQ��:�S���R�]����t4����2���+5�j]�]��=ú�`=��n!PDPSȽYV#Ӡ�JTX�V�������:̛M�򧧞q�����gu�#U�G�ƇMW�|��!򩞳�
t�gų�{3��J�ym�o����� ��H�",h�-��*QF*���V��F�Z���R[[iX�E*4,-*��Y[KV�D�@��JҖխ*V�"�ŭjҠ����T�[[R[V֕[h�Q+Y(��"���ұ�TcXU�+*,Kj*��AQ������T�AD��Z�*V*�jؖ��(�R�X��,���EJ�(���,R�Q�(1m��`1R	m��)�*1EPUX*�Q����E���[j5*����V�**�--����EAT�E
�1U��R�5��Q��ZU��k*�+[m�U`�
�E��J�R���#Z0m�ʬ(����Z�QEPV1b!U,A��Z[lDV0�mUE�*�(�`���E�TJ�Q+T�*�mkm�cl���X�AJ2Y��*"��+A�-T�Ŵ������k���/]
�1��b��|�����4M,�[כr0��mnP��i�wA�P�P�ԫs9<�����%�(��ګ꠳;m�v1qD�<�I�� B��y�Xy��R���G�/<��T/��1p#C�ՙ�h{+)��Xz2%ik�1!������i%�^!���Y�I�b��	Ƕ�p�'~mA�W
�I��nk����ќ�NY2�Ԓ���Y�R��I�����!��g��1l��C[�!�7���q��s�`��Q#��A�6���q�Br��I[���k����ڰ�n�{RO�_k��\�x9��\L&�Ѝnz�'(v��b`�Z򮀱�M��L���{�N������3�B��[��&t����u����<�)������y��-��ոF���ї (h����[��Mz�9�*gF�$����-����w�f2-�u6�ox��������Y�I_>K���T8�T|눃j���9�4�݊����3��4�7g5A��/���ό྆�]>J��������'�@j'�|�,�Y�#��7�l�ׁ��oW�A�r�α3��Q_�i�F��H��WP��3lˤ�/Ol�<��S꘶��/]>�V�#Ց����V�ܞ�y�%�i2���7�ݐ�J��%uګ6�2큩ºC�c���z�2n�(���AcR�`�0ޞ4����;�:YķB�#.�B�[�o��n��<B�B����VA)�4iZY��e���==�ZG��E6�K$Ts�O|]G�΁�jZ��G��J-��-d��\MV���`�����ޝ�ج�&ZW���f�l�e��5�2u<S��Re#�%�<k�^�GLɞ�ٹK�tw7���\�%�m�ԁS0�ӓ�0�7��~>����a��e9�9ү��Za�֥��,���&��R��L���mu���o&���R~B�q�	�U���Lj�T��c{��v�õ�B� s�(��3Ϩ(E�6|�}��|��3���w�Ǣ�
y+���xW��.�_�jZx\��&
�$��"Һu��\t�Ѓ��e��'\�磣���M������pP�Z�*bX��ђiVp[f.Z<�w1���6�ܵ�V�����~�j�D�Vl�*Ԋ
��p.�H� uD3vA��.;�ĥ���;��{�=�
ғ+�y�#0oL������,�j��U�v��{�#�+�]��#�>���	g`��#�{E?���!_{j zz�U��1��_����w�h���kV���5�49�u��4G]Ռ~l\�L��B�d��uwg��VZ��N�T^g���I�$N�ή���է=uҩa�}�'���au:��I�v�*�#��v(��I�}��Цb���GԠr��2��MuԮ�.+�N���TLM��W�5:�|��-����w���g>8Fj�U�^��m��2��3�AWB��7N:�s���Ke��j߆���iOJ�3��}���-�.�ꩉ�F�2W�u�Ŧ�5*�H�{���,���X�=<�'�0��3#F=J9���Al�)Q�<zjd֨������=��~��-<���X7-���a����^����x���9�c�<���L��پq�i���S�e�(_q/0����1�NP�����8׏c�g����pm)��y���>t���K�4P�8
�,+�sM+��l�a��jqzUsC�*&�fco{VO.��h����h�;5��[J#�E�US3;.ȫ������yZ��j�K�۞׏K�X�۶�8\Y��E�wh�z�b���Ϩ&e��y�xT�<�q.q��/K$y'R`��ou�'�����\�ֽ��:�$��;���X��^P�d]��BG���6��v�N	����W& �\%<�о����!񡀆� �erO̿e�v��*l6]��U�>�϶[��%*\3�׮��)N��
�J�h��W�b��g��[�ǚ������ٻ�yV�t+^�"��WV{�s!M�Z��y@9�§9�����{��eMܵ4��-�S\u��mzпnz�Q���}Ut�7�)�����w��r���)4:J�3!~�*���j=2���L<¬��gMW^��Rl�#�XR<�^�vͽ��5sy�a�ȃ����L�;�Gˏ�=f�Se:�h ����r���}ϰu��j��׿ X7��6x%S����:��]VaW�I!�H)�>�x��d�t�˸^%�r$_��X'���
z��3C�W�n��ZXp�a��n�����A@��nW�Ը�R�{�<�!=b�ꇲ�5Y�֡趎��Ԭ���yG�o�{D���/�WP��a;��E��}�{潪���x>�ԤH�W��%�==�@���~w��C��X,�׵���3�P�Ӏ'�R]j�g�Y�M���r�K�U���b�Y�E��«®��}B�kQ=�f'R׎���&��o���1�3�/%�NA�}��	d\���i=���c:�P��F(��8�;����TiVs��ò�z��;ڜ�ׂ�26���>J'�Zm���3� x��N��{�*ދ[:\ម����}�*��V���}y	���-�`ۏ�����&�J�x{Q����y��Ρ��ֻB��\3T}5,�Me��M�t�js+����s��������s���PʜN���E�x�sN���+�oﾪ�u���>����A�.��>4'&m��*��A/$����h�/~왆���� =~���+��=����,��/�����D7��8��(�$�L	kS�r�*������v+�U�3�q�Urd�/E�R_l���Nƽ�T\�z��g�d�%W=�B$.�驍�r]R#A�<]���
��Cx��MOX�jX�NF��e����:�f���﷔����|���Q0JD�q�BU�T |���Fe^ �*�w]�gW{�uo��\�mr�Y1���3�E�_JM$�K��v�ud/��5�PeEeymȖ,v���G�ok�OfR�ص��',��p�I/���ϪWV+m��n&��}+���rn���-�-Zg���L�k��#��y[˰�kɜ��c��RR�P�N��Ky�e+���۾�|�{r��]�	��h�s��9����b`�^A��ij�x�%l���U���U3�U����ƽ��n&<��,>���<Gx�<�}��*��8ń;��R����VNu�t�l������u#w��7��O������r����8�L���N�t2�}ckf�Q��pvW���u)�%+��L>��Պ.��Ь]�MZ3��-)��s�x�DK����w^�������Kֻ�����[-;��W3��𥉉�w����9���=y���;k�A���K�9����͸�Wo]x`���o�n���V0*�d�;�Y�J�dK�<|3�ԽC>N�T��)�=-��X�Gv�z|�7FO�q��Mw����k�^WNRV��\�Q�ͥ�Wj!�x���5�t�>D�&7\{9x r��#�j��L���F�MX��O*�h��ߣ+t�ݝ���kH瘧�K$G:���=�c+ܘ�P�ʾ@�B���{��ߵ���Ϫ�o*t�g%̰F�'j����u9ւ;�l;�P�o�(�~�!.TYx��7%@���)^�dK�"9���/ ���e���"B�s�G���g�C%�R��+�S�r��hwDE�}Z�}��S5�!c�W"�F��H�XR��,��+�u�Ƽ�����z26-"�<�؞΀�5ΔJ�S1��L���C���Ya��>3OE0�\��mQ�R�_�x%�`T�(�S}�J��$��G�r���ߢCp���@�0	��o1j����Mh=ٽ�[��5v�2X�:�G��Ea#��m0��Y��a���u���p��-�}��<�:��Ѳr��"\�D�&�`X�����eR�f��R�X)XV�b�O�,�zD�����O��52�ռ�n�����h�X[]T˅�Ev��P4�T"��(GtI��v��s��3K�ޘ��|���^�9x4�Vl�(ȡ}�Um�O|@];�Lnf�ne�1�<�7�X
��U��@T�=\Rҧ���cބR���`EÂ���*X>�.,7ܣ�e�ß{�ꊶ�W����Ls���>B)����z��>��k��W������6s�y(��Uφ���L=��<'�\\�̆hη��h`CX�<���I�n�k�n�]�[L�ǀ4�����;���,a5���WK����|e��Pa���+8��o^�5q�g�S8�~��w3#Q�e�s-���-E~M+�>��[*7-RS�e�ט�/����ld��\dK>ܶfS��y��08�wS�/:٬:/�'�NF���ݮ��v��`Υ)m�au���"�J�^��-��귓� r��u��b��;��+���M�V.���Yh��Zj�Te�J����ුJǝ�K&MN*-�����7��_S��9�(�c8ތN�ל�Y�i��լrі贵�,Exu��WU�L7CU��^,k���箳��� �f�Q˂wR�Y�pv�[�f��:�5Pu�p�w;E�Z����=J��q�cU`�:z���5+:�Q0d�����_�����Ƅ�v4�xk����D?�ڪ��ȫ��V9�{��pP��ǤNz�:&=r��r�GK46ûF��,�Ŕ2�y�WF���X�S�>����B��-���\\o�������Y�L�����J�u2��W�O�ĺJ�@�U+fw��L���U�#���@�<����z�,���j�B�bn�rm�^wͦ]w`�tJϵ${AT�gS��1��B�K�L���֟7��.�5��cd��Gs�ӄ�[�H��D��҅]'���n܋�JMf���ȃ������e�tKK:py^�sޒ���;A�5�<.��!�����R����f��Ip~��ϣL����c؅�lU�d��v���D˸W��uS�_?>�ߥ�閻�s�t�I}�~c-�-=�D��
ܱ��{Jð����V��B���(N{���^HT���zt���z����<c�d�BH����+��j�Ͱ�m"�����
������^�'ӌ0��-�Ŋ*w�� ug��椂��*�d�,�u��^������;U�?]+���0�-���{��U��٤WN���i�G�Tq��d5ݷDl�;�H[0�bձ)e�;3�%]�d]�&u�*�*혭�M�ޗ厸?�zXь�[�����/��|�#��Jǅ�Al��Rz�g ǻBc�%�ϕY���
L���:z8�6�hO�=����C{:��z��:�=����qWh��Vژ*�&��3�΢�J��rR��wy���ڱ�i�w\��t��*����åYh���K�Z=�c�Iǩ����{��j+޽��/SxN�Q�<�:����zlNX��;�� ^�����j���	�v)g��'���n^�䎴&.��e�����J��kM�46¢<h%�p/�9�<����9mH��{5�=�:E���2o�z,���d5�ns�Qs(.�{>��}S��$��[[W��:��E�>JE3�9�Շ�61������e"9T���s��ԓ�+��}SB/h��K3��D�"I@�=���_ٱXy�e�o~
^ysmxW�M����_Aɏs��F�u:�O}0T2�G:Ri]Wڕ8��z,��k��ugTUf	�1RJLi��=�{Mx��^���d�=k�O;��?N��Y╱�����zD��V}w(;��(p���nq��Vʥ�C��x�[Q>�{�l��wo+���:o��Cg�ķ�b=�䨬������u��-�]+�]o��6��0?�ǋ��J�t�����=�΁��
`�Q!{�c��{�$�`(/}&���z�&a�\�`���<�<�;֋7�L[MfmOI<,=�]2NΗ}|6��X�B�ޡ���Q��TW>�M_΄h�<��z��T�J\a�;RI�^�r��֡�V���U�7=�3����ɝ1�@h�h�f'�+W�/�w��;��ĥ���c��ſ���2|�:����۰���Lx��{:�(3��c�7��Ġ}뇻E:|��"<z}I_��p�]O/9�P��Ez��<t������k��~R����.y�=�s�cM�Ͼ��uia�&����N�^Ba�}Q'n\�,�O��p&ǝ32��9OɈ�<lU������4��t�jJc����ī2��f�$1u��(h7m#��T�g��B9� j?W�k&T&��"em���~i3S�i^�,�=K�R��f��e�~b���ɏ%�hd�o����j��OU�����?f��f2jkɗڟuC�)x�hWd�(�\�s��Z��-ݳM��І��W�n�d&|��x-���c.���	��Y�c�m�3��;�:�-�x��,�d�r�c@�hnW�t��:�.c/z����0J��:�'����\(�8��/�\�3�#���*��`��G��a�Su
�帩)x��j��)�J��{��2�VK����ڻ���]@G�\Ώ���"�o^��&��v��51/�8��A�����7�dZf:K��(�a%<��-`��i7�r��]Y 7wm���0ӧۛRwr�4b�(���L�/A;l����o-s�ӯ9�G*������\[ldr��:q���^�� ���Edh��;��6X�b��Pl*,:�|rN�v��Y�F\����}r2-	���ۨ��EQN�=i�7�	��5���`ל(!��V%^fos��la	�>���ht�,u�\�Ҫ�)������݇���U�2ɦ��n#��y��㹃$Zz�Eܒ)Fp���K�t�P�y񮛯�����]� ��V�Z�d�3jQ8�,�e�o��7�2Ƣ2����u;�-<Z�t9m:���b5�][�(��Coi��Y7M�\�|tܫo!
I�n��y�l�� ov7� �0��`4�Q�f,΄�ַ���&��b6pl+���ܟf�V�)�j�rb��V���f�D^am��>������3O�D��6��[gV���3��`�oY0X�����U�Gפ��.�]��ʒS��=�U[w�=+^m�l 
�իo�Mo��z���4eoiDZ���O�%�Zu
ǩ>�������9��nV�iv��SF�ḫ�u�8ɽ7��l5��)NW���l�'p�KˇoYk��BQ1��#YR��b�Mh.�ķ1v�ok��3л�\����ue��]w[��1L�:�.t��Z'k��TˢH�s#H���C܁���q����v'd�Z4��K2��(��["��YQ�V���h8_S�����]�����vN�]S&��
WG=���*�M�m���_EZ.kF�S�7��bh���F�]ٱ�h�����[Ԏ��O���s�]�&� ��n
s̼+�V��e��D�+��S�br�Kk�Ծ�[S�X$(������U�.�0��YGd��k/u[��r�o��9E�����U9��{sn4��:C-'�:�ܤ�;5���`���v&]J.7	��_(5W7:,S� Ly��ʶ�h��cv����eM5{؟;��ī]{����Ќ@վ�^�EI�Jot�jg�r���+%�=������AQ��,P�.���jo^*�3��zS����jF����������i�^�:-۬���_a$v�{Ƴ�d+���jI��ѭ�=I�#9>�����u|(X�RV�11b*6�б�",UEH�YE��Dm(�b*"DZ�Ъ"*�UT-�[*(�jT[eU���%E��-�*�����Z�[*���1�TF6��
�؋���,Qe��*"�m����Um����j-V��Q���L�*`آEDE�Җ("T�(�YQb5���YPY�*�т�%��j���Z��
*EQT��V�������ҭ)ET-J
(�ѭ%���PV��*UU�j«�QE-Xbd�(�*(��D��2�E��DUH�ԷE��U��jҬT��ZV���+�iAQ��(֊�VE��DTD���()KeZQ��F���R�j�V4��D�T�J��E�����6)[��F��h�-�j*�F#Te)A��EF҂�,[h�)iZ����(��V�V�aR�ڣ"��J�]?�]� %�uF�]%|�4�T�,�x��퓷;c��r�#�tt�
ĭ/��:Y��g	�[����D�*:���u�����ݣ�A��	i�H��f�Ma��X;��l3ެ�9����9��텉i�{���M�rK���x�t�n̓����![�U"�(�f�O�L��h^y���y��|ҭ~�$��ؽ��Y3bx���5ΔI&c[���6:s/3;=�����9gqY��W\:תe����~X$��Q����`��疍s�ZWN�w�y���ϛ,g�{4Aӽ��@�arƑ؃�@*e��"�g|%
:�%B.X�,q�yw��r'B{�W�~��~�q_���3�Γ��=�����
��߃�gAg����ؓ�I�|�.��pFn��vClh��>�T�X���E��23zX��r0���˴�8����κ��l�'R�O�xc����k]�ֽ>����ν+�|�Q��ڀy-
�R:���O�|��?>}����:���&? ���,OB�_����o��eDeLUy�{��c�ͭk�A����L��x�;z�<S
�%����p�3�Vfң���P��E��|�[٫%�6������������z6��A�ܱ1(D���6���%���6��d�(��"�\�F�B7^I*ђ���%j]�i��Պ9���������������h,I:�����[��+0Dʹs�zz#�;,I*���2���ڞ/wJ+�bi\T�W���m���;3{H����f�Eq���q&7-����9҇x�{�����jpÙ����w�w���hϘT�>���Ei����Ǧ��6�2���	r�j���=y�¦|���e�3�WJ����~3�~�/+-6��fUQ���g��,+�o(��:1L��`���	�L��]}'Y�-g��W]���{���M�����M��2,T#�ؤ�=�Y[�XU�2�}����-G(��[���AC����v�oR,X+��>��fuW3۩���Vj�8��]y�/Px�|�skK����7r��]��u��@��(rP�*`�9�ލ�έf�
�w��Ħz\#_��#�U�P3�x�
(O�є+���[�kݿu�t�D��J�H�
�z�u�]Ě�򙃙Q��gx	�����7��r���8'���$W��ZU�I�/.�5�n܋�II�͏VD$gxۗ�ʢ��˞N*�.�}6Zwח��8oN���e�А"�>jwv�0(���OwTv�u���4�-�|»WQ�=e��	w��Y�o�� O3w�$`�r��Lq�v�'�[[�B,]�s^��Z��U���+mBV��:���)��I�ٙs7�WL���>8o�%g�Q����c�u�EV"F��YO˃�3u��G��A��o��mJ��$�&�J|�B*�<�(��C��]Ï�l�V�*ab����v�]�[�SM�m����~�w�~;�֙��,�భ��NV�V��a?_����}H�V/��������Zu�*�W�n���a������@�N���v�'��e�s&����
�B�@;���h�
�o�;i�͸`��3>u8ρR�W�K�D��k���˶Fz��D<&`Li<�:����p�2��<z)�LΧs����ũޚ���$�;[:{�:���)JÔF2.Ш��JuT$����p����E��N�Yx����L��5K͐��z���ߖ���T��ح�(�Zi���0����
��gwOmI�)E�v ��D��\�B��C�br�o�몡�d�?�/89%ݤ�2���&� �	�}�nn`�W2Ox�Qx�`L�'&1UK�~ ��*`�ܯX�"�5�ǧrx�ZS��W�c*�P��m���/��R]���t��x��R*2�������E?��g9�n���+Bv�6"�J�k���6�=Na)��*pn\깒��&��;cF�T�|�U��®��F����kru%�]e�j��ڎ���7x�~��5��ʮXϰyˋ��
K�ћ|���̠T�y�{y�7j�>��A�e�L���HΪ@��@p%�<���Xx�c��{sMk_ze!YNF�5�\1��i5�N �wu��"�6P����[q謩�_�������{��a�y;�,�<�.

����N��}r�`�e��D�]�Wڕ��z,��x�}��*��ǥ>���P���Ɂ�Ev<q�6�`���-C�)%])�n_
�`ݫ{���Ż�3<���e�����J�j\�`�H�6Q�\b�}s�;X�ePĭ�ǳ)�YI�����W��9�[�,{)� ^W΄h�$������u��ùw3/�`C���rЅCS�綊+O�iOh��7+qOΙo�F���V��GtB�{0�O��O���:�+,[�����&�:�FxR�5֙�GR����7�`�劽-��ќ�\k8.[�#ʱ�a�iH��~/*�ᄿ����ߨKI�-���	<5OWJݗy0�5����Pou�˙|��{���eN~K2���"^�^9�4�@vuE�6���<E�g�:�7��ϙ�{.�Z�hZ�Q'��3j�f1CV��5. �����1hݬJ�c^yi]���n�@X:m�)Ծ�������n��`ءe�;��h�m�ń3X���7��X�}
b�sm��Q�C�o]�ʫ�9���I�Jf`���.[�gO}O]z(ϋ�����T�hj\T����n�WV������8��<�H�K���5;զ�kY�ʆc���NNU��x�V��p���d0B���p��-+�T3|6a3%ht�o�����1�Znv����Gu���)���7�A@i-!�Do+�0^}]1�Յ��=�H&���
����{�&w�)U��sʂJe��G����G�BA=崇mtɨ���WY:�^�ٶ��2{��>�Gʌ�(ل����f�B�҉_�LưP_M�&��c}SNot���<Ǧ�R��LT��*ŲT�(�ʘ�`��<�hs�ZNq�>�gxp��罾O:���.�~�-�:�ְ��x�9Sٌj�]X�%�YS*�.+ɶ����3=��a[ԐxV,��w�X�W�}Γ���a�3���%����ck�Տ_��w,Z�w{�H�Ӗ^,��6��Wr���F n�S+��d�(���'K���/����Է�J0��-�}ʮԫ�1��Q�2�$�օ���g���U3'U����2�:�Ú�V��<�F
�|��'��z���2mC#�x4� X`��p)�sz�Cm�\9�#3z������-֨��z�F��2���8���:go�f��F���=S.����^�^���d"�]Cy�/DS��IΎ��<����[0������y1�AL !=tW�qp⮰x��n_�;��1����ϋ���]%])K{�J�+Lu���Sy+,���89ř؅�.g9^1��yl�n�t���Gݖ%�%�ϣ���_jb�t���X(���n��n/���� � ȟR�.��j��h�X9����f`� �K�^��'u��f�*ϯ}5�#����]��Di?AR)GB������K� zj�m�e�N�(}�t�T�C{�9pz�Gu�5$���g�VZ<l-5ʪ2�*Eט��o(��1L3myr�z��|bm����"���}8��Ϧ`��>i4l�2,������u��X��F)��G�y_�m�W�?)���o���Y��>�Xd\�C]R9�H�����<Fh�t�k#۽�����i��n��3C[ANw�\�`��z��,*�^e���dqz��&��<<�q�y�*�R0�*+�ު�#���=���;��jR�c���f�D�^3*n���P��Ռup�D�M&(e��6�C9+���$���6�Y(ͱ�]g3+����=	���WDv[�Z\\ruY�/�RϚմHt��1����������<�IuUIi�:��)�c�m)��ֽJήw��ç�ОTY��X����N�^D�עhݡWP ���J�t]�U3םr�EᲓB��,7�3`j�Z}.v�t䮧~��z�v��{������� (ޣ���K۰�ݹ���g�
8)F�1F<k���|��?z���Wp゙�qףc�}�X�GE��O˃�U�5S��[���-����o�RN&Ehs1��Qkp|�6&]Á����H�>��_S�wn�ONkR	�3�iy�\��W���,�V���a`���^@;�
!�l�¶�v�5�b�i�@:��j�h��<e��O���������$;�HS~ɷ��=v:u�H�+R����4��/�f�0{���u�9�"�����V��ː�ǁ�E�ّ��%���0��W2��9�<z)�rٞ��ڮ����z�9�S�ԁ����T�X����k4b��J��W&�4��s��9��9��*z��.7U���q�@��s�o���ڂHp�Z��Φ������-̳nsP38r5�2oq✨�sb���A��[���#2���-�5�k\^�3˼D~�7�� �U�(�eC��i�--�6�h^�c8 �|i�[���[��>�����W�p��o�bd{��dj�B���O*��X*��}O��ZVj�z֦�����hQv�gޔbu	���M��>7�u����wuW���!�����fN��ף���F��{��˨�iKa����\�A��/D��ܥ�_��f���]}�Adq%�`��9U����x��2o�7��ћ|���\��>��,�}��z�ag�MI���@����[� �Eg�,cw5=7�|�����eH��#���:\�N�3�;�El�	�&a�x�M�4��B�Ec6+�i����;˷�q��S{$Í֎���A���▷�ˇ���ن��� ��Zgܗ[����S}י�@���?]t��j{2�.Q��>���*�I*�"��;طF��w�fԾ�ȩ�K]�r��QYcz]%57�lQ#��jy[˰��%Z=Е%�:�l�i�.��T�a5��}���R��a�^�_VS3z'7f�Z�ľ�J�ש�0OB���ц�@3x�����
�b�}m������G���MdN�i�1�/x��v��`�jٗe뽨�>$'s@���;��o��0@��D/ޖ�/+=��|�O��tS�dֺ�\L���`�U�̘�L����u�e���hB�f;���G�Z|+J{FL�"*�&>�B����sr�a�˚�4GBo)�{��	�\�1G^�ſ&ax*��U�/;s;k�1��<��s5.S�4>�IU�{Jv��:ۙJݻ@���8Ю&�F�	����9���V�uѝ�b���.#�۰�N]�h�7���rb�W	�:Zx����ssZ�Xy�P��G��10ʶ�
yPcҙ�)��<\���x�_X�Yj"f�R.�R�j5�=�9)X+����]��e�N$ty��,�����5�K�3Z��i	�º�v���=�?����?�k��+�!_\�8w�^���C7�0�y,k@N�+8��K��x��IF��{@�h��ֶP5x\�ʓ:u�Vy��͓O-�/k���@�󝦬���k�-�g�x�t�n3`��8���Qr,u<��,��F��ֳcs������ݸQ�����r�ɽ������� Y�c�ϟh��oz�E��2����Ђ��;��P�b� uի�)�����(i�3�%B�}`��1�]T�.!F[��@e`wgA}����7n��� �g$��t�6�0`�؇s��SᒡYsbǔ͇���ΔJꙍ��[Pկ{P�rfw@M����~�&[ڞ�p�J]a��,��!B|���JUϣ!P�n#�8:�i�+���0󹈷}�d�`;�n�T˅�Ev���:$�DFQ�S��uf7�Rr�`n����e.���}�Y�3��H�R(^EV�9�G��ʶ�w�z!���	^��]�f��4�S��3����蹮"��5~�����,�Fޝ�!i�8�O��z��ڳDP�m��Fz�}tϷƑ�0��yT�ջ��%�^����c-�ޡ>o�rX5�aX��E��:�,ed��LS�Q,OJ+���y�9��di������m:�2k�e�λ0+�_H,ny�iz,kL���=p�ԃ���ג�G`��Ol�כ�uT���ξ7�M�p{/L��vX���d{#��=��qx�k�Wpmn�W��J��z].�]�ze�c��;�-��cTD���P�|x�����s0�C���	$��/ס��zl˹�����e�^e3��-��]*�S�Ȗ�5�3{9̱��p�T#�w���]��M�Y��N��q�unL}Q�U�%,�ݷ�/�Ŗ=�M���=-U��wJ7���ԚB]���?m
�W��Nl����2��U��B���D2՘N�x�H5�ˮ�K�ZFk��ʳ	�eu��:��hp�&:�d,WP�$�s ��<�����"7�ǻ�a��69���3�j�	�T����cȢ亅v:�{T���uJ��˷l���,��V�ى@�:^�+��r�5CcpZ[.��mU�ne	��t��x���olf@+fDÉ�3F����<���︲�;y`��ԜWu.�F�qH^>*�5q��>���ɛ(p�4��7�EN��v�)�s��C��)��/2�P9�S�ޤ�:�T��m��ܧx��`lu���.��W���\��s�%�ng#��5�^8�n@)3+�8��fٖ�C�1�2�>|IΙ+�X�ȧ#ko�,�F�$�i�I����7 n��&��(��� ��(��|��_�;K��.��,SfS�V��W+y�hz�N>�I(ν3^�7��<�`��(܇���\6�I��w���r��ޥ�Θ�[u��,hɧ��SXPZϒ�\l�v촅�k������Ҫxp��s˔d�U�oy�5m�C�i��u��;��Z�Z�MJh�Ïh g0���	2��f�h��r�Uf�c]��봷��*��(gMZ-���I�����w4d*�^�j�w%8D?-�s-m�N�ڝW�gN�{N7b�$SW/�V��UԶ��(fv��(ؤy6�6{�Y�ҺyK�`	�ڳz��\�;�ݮ�_;�w�*��V�>�.�s1�f�hN��h��[�J�;����:ײ]��P�5��A>άT�3.űՒ����{n�����ݣQz�mw#|01��f��Z��z�P�S�YOa�X����Ӭĳ�+y݆�a�����-�a�Q�CU�08�]�����5�f��Q=��E��}�%E�O�PP�Q��2����0�6����5O�c��M��ۋ��V�\��5�CLĀD�5��;�[�r�8� ��v�/�CR�	�ˡ��@�#�o_:���ܮ2��=�\1�h <#0�t�n�֜��H7�e��E���*I�:ѝ�>�����g����޺ՈC,O!
�E�O�o4��u�kJ��j�4M�S�(�4���,�"�$����,2�&:���;��v���h�i�	�tp�X7;d�@���,�ZުJ��tv�����B�?	t��9�;s���,�r�[�5S�'O=�up�����CÈ�څҥ�����#+����b+�X���/8:�}�����j�j������Z��Ԏ�#��-�]P�,U����[D�����F�n�T��lD���V)XJ��-(��H��+-�"0EEb�[Te���6����DU1TJ��b��*��jUJ�Z�-J���`�5�"�*�����U�J�h�1j-Y���\�-kJ��Z�e��"�V�EE��J�Ue�DR�R����3\J0F�ʕb�q���5X+b�X���Z�c��جL�1Y��Ƣ�b*�Db3-�c��lW0�ZX �+Aa�kS%jJ��+*�
��P�EV��E����̲��V�f��Ir�ER�`����������#e[�T�[�UkKZV,r�E���d�X�ZV�j�%��E��\1(�Q+mcKhڢ�X1[J�.eDS���̅T�mY�c�$b+�F��ʘ��F*�[-̭�j\��28�f,�hQ��2�,��E���B��[��rڵ�-Bա\̘��LLLQF�Rָ�̡cR�LʘfS(�b��.b�R6�30H�R�c�\Lʷ̦-h~B�'�ͦ�>L�!9.Qy��>��A�Z�ѼJ�3zPo��HW}�j�6�٦�@�\�պN�]\���q��gu[<�隄������*��/Z�t5]i�E�.zj��\̉*<w'���{Z�[m=>�9s��uڬd�|6(����^�$��%CH^b���Q)U�n�o�>�����z��呻'��6��U��҄�3�p-�<C�t{ē^q?+�mlȬ���-��k����e�+>,�SV�Oo����� �ȹf���s��E���y`���}r���(�=zzUאyQBN'A��[�Z����������Y�V�!�(�U3��s�{:����C0P�e���3��Ҋ�p�3��9�4/���.xv�������Mu4�f:@���_Թ��T�gT�zR�/[����;.�{Ǘ�K�W[��%�#���ذ
� �.�����9�u�L��x�/���.<l�A�F)ܚ�h�\��֊<մ;�W���(a�eه>~4�I*e��-�/�!�=�w�{rDu� ����oK�)�V�`�r�Z�>;2��<v������Y���&Iy���ƍ�hr)�P����{zhHl�%���]Dq��H�%�䫫m�۶�ܧ\:�V���z�D�2jH��lE��~�j>W�]o�q2�Sp��R�Y��'��t5sj�����qN�o�ㄞ�Ȫ�؆��)
���9�w�HzG�{��]�czX	ʺ�;V�oEiaXv'9��'��ٔ˕����=Z�:�,'C<��yr&t�/�}�HL�Ё�� V|����u��R�U��si]o�(u����9��X/K1�x�^�=W�����ƒ��#�Z�^�����4d~��n���Y2!�}���a�W
��l<z(D߽Y�8Ŭ����y�琕�a��^AZ� �����-e�VډC�]AAW|�wW
KYz�C��0���'R퓮�ɖFl�n�W�a�=�Y�I`|By���b���k-s\r��o삙'&B�ҌW��N�0��-��b5��A�P:�������Λ%+��ؗ���C3�fϩ܉�	�"&L����P��+�e�<���3q����VSŌj[v	>i�J��췊�r��)�{d�^M�j�4v��z��w��)�������P���#���"����5C���0j�ɾU���]��@R�y��v�,��{��q���͍{g
�4(���)��j�Q���j�]z�S�"n�Vj8��o	�ڏn�P�N�u��o{]ۺ�hG/y0����X����X1��� J��mc`
���4�*k����4��{`U��omI�r��l�nf�I�V*�S�'Djc^*,`�`A���� ���U���.���*�[H�M�X�����y��ղ�`���~P�)���29��P��H�I��#�Kq�c>/D�u{߸��q�-5��=��L��C�mh�$�9g�Cbe$�]̴�6����' Q +��=�:��;�v�ý*�fz|e��G����D^��}'���uk�8l��<mY>4����k�|7O��f��]v� ��=�9)���������J.� G�}��Y��g�^�&Rf��
)�o	L�#���;���)؈�3ç;�ت�����7�s]?��� �CWk|M�
Xg�(�&�	���w�`���]����-���"����y*�y�
����]Pq�Hl��`�~�� �Z^d������d�M�G�̧<~�	�_K���5�vb�e��-sgA۷|#�
����C��^��q�2�U��~O���NU���B�]y�%�S.]W��T.�^+T���8�$=�#�M�
���]�y5c���ӻѓ`��� ��kz;��}�"�U�r�VK��(��u������ޭ�^Rk
�Fc�f֛�:�"��ڬH)���v�w(��:2��x�c��(��^�y��Q�¬R��F��K^�z���G>�"^��S�O ]G�ū���w�!%sY[��w�����0VZ�/妃?rOԨl۸��J��C7e�=Fa�t�x{�q��m����a��T�����6��{~�h񿖚���2H��0��|���)��r��,���r�g�cF�<�M�V79Z�*�f��x�߳`᧏�X�*�=�x^�ۣ�SM��>y..��Y��� �x����9�<�/d�FV}sbvS.�ZQ.����"i}eI���gz˴��$�l<L��Ԩ|�2�p�+5xd��Q����`��n�׻s�3�5�@��%u*uP���.O>�z, țYS.S>�JZ����}�]+�צc��"��i!�W%�u�^�hf��\/��^kCҨ��JOj[��_�D����u����ND�s���[b�\�(���K'�S[Y��4Ƨ�[�w�U��כ��޵fi�a��	�j��XC���u�������c��a�RA�^:���,Z#���-�`��_f���.�AEr?�F�؊��Ў'�&2��K�_idq,�ś�i���r�t�v�sO��(�J<��ZO ���p5�\�,�4w���E-�C�η!+vi9Y��)�ω�8Ew]lu���_Ӗ>0�Ǿ�OϷ��K�,+s8XY՝p�d��(AS��-�a`V��o<���ڂeq���q�3��@z/Ϡ�������-?w��+њw <�s�^#V���U�&�+6�����mx��\}���sD��9�3iO#���ݧ��-ֽRw.�����v�����5/������Q/S��x7�yl��aչz=g7X�v����IW��Y��]��1pȣ#�����4�:�V��/��ҡ��u����}*�U�oy��l3�*_�g�Ա�S�XΧo��Q������>�Uh��������H�5�=�.Q��{�Yp@~]��59C�:��1�6]��YZx-�ѰW����}�B�N���Xn˲*�[eag"��6Q6�m��W6��uKU�j�+���`��GWC��6/L����@��]f���ز���̡��?�=O=79Z!B������叄j+�i]ּ�W�`z�k�l3WV���ކ��+_�ňr����݊7�0����+^zN�d�΀��U���*���:�ʵ.;4_ �tlh<ڠj6�N����b����p�g8�?!�C�:��6+FvP�[�(�wp������:�ڝZ:jƋ�uVfu�yɜ��Z,�-^����,ح���n��O�Z�u"��ӏ�O��:�wd�:.g�^Uʅ ���#�vЦ{:�({�J\��n�jӳ�=L�n^�=��x�?g�E]�O�P�#�.��%���$!��b����f�u\�{�q�Ϯ�j�H[�AO������ޯ8*�
v����:�!P�[G�y���}�_X~�U�y�����z���Mf邒���E[��kÝC��˸^%�_��^��	ҋf\���]~�!���R��z:�Z�>ޗI^�,+r�Õ�Pzwm,˺�j�˻؝�k�<Z��(�,�V'��T��ed�G�������$�{�G+�ra������2�kڶ��o�G�)v�ʖ8?���4c>�������z��ÍW[�i�綩��}1L��(`�ɑ��ڕ�ȼ���p�6��%!{do�ԕ_prOEKj�_ϩ�>��y�אV���2=C�]�P�Zqo�3�Rwro�bol`��P�o��P�����t���E�`c���7�Ҵ����f�k����.ǋEê���h�&�R��&Z�/�n����+��$�̼Z��ֈ͜�v����}�&�Ʀ��*!�#�9��XИ�Y��G/K7�r��d�kc�5�,����B���-�Y��
��T�]!�������o^���.��UZ{Ʉ���BM�tL�z#'P����>6#X��:�gv{��.���6��.S���A�<�"^�A�	~��{��ʺ�ƾR��d�� %k�����dW�G��y����
��KJ�-�"��췊�}N\�*�Y%��|$�1{3�]�Wyo_l�(�<�yY��3�"����wh_!�IsS>�C��ԙ�)���d�^u�V2�=����Wt��B���,
��׊���j,�E�u�� �\bP`j�{�u{3k\�7v�9�<��q��za^����xԗ��&W��&F�JM#�����q�#���M�y�ȪP�]d�8�v����Y�L�5C�F֌���,(gvj>^'7��"���܉���uG�c���]<�|v:MYcz]%mC�e��H�f�4ƞ���ߝfK�kt��6�˱��ICk�)�Y+\%>�UF��t��:a�L&��m�^�ؓ9у9��OpLÁ�L�T<�����z�d�Zia��)��q����
�P]�Ws]â'���b.v�,��h�r�$�<ΨZ<Z�M���Փ�C2&"�_LR�e@&$�ooG�f�w9w=������fvJ�W\��G��i�9] ft����,�9��V-荘�W9,�ǫ <��\�Z�7K��J��;��|�u���hC��낮�,�܂�L���_���Y��T̷s��_A�#xݚBq�|�}�+g�������u�(ڹL :��xx�����W�{�\��"�G�O��3y;1����۰�N]�h�iX�wrћC֬�k��Uy�7Pf��m�[*��,�iW���"8<�I�L��g��P�w�h�ԇ^�p�K��zVZ��E4��?T�*��'8ԉA�p�u;ᜭ3�~ꋌק!��G^��S0HkZ������|IإCfnd��L���T3T����.e<�kh��9bE��o��4�ϦR=*��妠$��9�ܙ���s�O���ޤ|y\*� ��mS��<��?.lWǖ��vh�%��]�E�yK���=Ъt��v+��.yzZ����o��{%B2�\�ر�m� e����M3�n/�b	,��F�xeC��j�A�ʮ@���.R�z��O����z(��f�����ڲ��r����� �˱�YY�#Û옥%�Yd^�V���:���X�{����h�3t��o]^�ڍ�hs[X#�Q�t�#��X��z8qk�ɧW}X�B���&�iX�ۃC��wt�6r�.�h'��z�K��Ҳ�V;��˵���H�h>
Q��f#�ZU�'���脉���=Wl�*���b�~�d|��c�0e��.���d�Y�i/��G�^�\7��^kCƨ`�m�{2^��0�<Tv|"����>D�s��͎�h;WyX�Ϫ�$�&{���Ia��y$�gl�}�F��'���i�a�OR���$p�D5�G�̦�^�CC�!�����:t��f�jֺЛ��%�\��t�o�d3N��w��&��s�{]j���r�ono�֠4�K)���ξ���+H���,ny�i`��5�{���
'��E�v�3X�1Z��S<u!���z�E�2�Ŧ�9�2#��zd�b��y����S���rζ����Y�Ca}���x��>GE7G�Y_4�X=¬�pyqq,ܶe*����|u]��3���'8\����'u��4՛F�髋)m�a:����|%�v�cүɞ#7m�x��ϴڀ;z����K��';���g����t�=�RXϥ"�E.��*���t��Z�''Zm_�1�|h82�)��אkg �#�K�Z�+�o��:9[�ĸ����=(�]W;���'���l˳ۓ��ҋ���VP@a5�BQܳC�;�1�&	�
J���cX���_���M���׊t�U�n������-K����L&jr�V�J�&c<s��\l��8�3^���ë�ˇ��p������3S.ȫ��(3qO/DK�q����&�VS�ք_MY��Z�rD��^~M��
�"�(&e��y���0'��փ"㓝���{�}�x{G�R���(��M2H��ݠhji@mu2��ulNV���Jd����9}nN1כxlgM�nWyֶ����xM[ŀ�!ӠAY���\�e
g�딡�J\�x��\�������ܓ16�v�w��U1i�P�#.���%��B��,n�wk�9���F��ؘ%���U�2mQvM�ʇ�N�9q3�W��$��;L�0�~4� Y�{Sm�G��ﻦ�{psk���XxX��g�M邒��B*��`��^C��]����է9��V�ecK���D�j�0��J�F{۞/@�j�T�pXV��^kR��5;v��5���n��i%k����e�gҵU�G�K�����13�w���x��S�z�yE5m�TC�k�*[x�z�Xa�ˇ9�^�E����;Z��>�+������Tn|x���	�S��e�ǵ�X��i*޶�������.��2K8���U��2��ڟlή�� �
@�|�k���w�X8��Zw1��wy��Gb��+�%��Z!��Sx�]D�yވ@ӧ�k��B]f��n�%W��Vy���\6����sB�]�jR��L�B��f8�B�I �o��ZQ�h[�uLO��� �[U�i����J2 U
++{�U��Vx�vJ5��h�n`��I�D�:4ݬ�^d�k/�8��(�m���z�Sdq�SU�
W���b�喩�~k�*^�� �7>�402j�&e�]��N����V�gR�iC�Y2�j�{/��Rls����`���bೣu=��w]��X��gMvhH+��#�w��}f���KAR�f���t:V����ޑm��TSW�N]#}����z�h�ӷs��׈@��8z�WR�7:��*��
Z�ԭGiN�{;�ns�]s��ZaV؎���)ViA,��c?@e֘�R,���l\�jr����ڹf���̎A��3j�&�]�GA�F�LџjƏ;�M'E]we��Y��E�
��_(G)'5�X� �_b���md0�C�ΈaWǝ��r��:����Ƅ�J�I���@[�a�}NWl�ZS��<�6�U�eq����.\�R���]K�Jh���5��y��{w�eS���:�P65��D҅E��N�5��][��O�\
�؏e�f$RΓ(q�h+\2���uN@�oF܍���<�J�w�]RςbE��-��O.�ѻMЫ ��њ�T��&j���PSѝW���IH�F�3�Y�r�4�*Wa�Z��X��U}j�:��6keiz�a*m������]���N_r�D�ͭ��;�d�v�Ay1���"�&��l��e�څ�Y�;)�/��x7���I��r����M[����W�R���*c�Q�I61��K5�C�h�O[��b����X6Ge^s��X'��;/R(��n�e�[;����X�����8�	�K�{#Y��[rIN��j�lJ�9Gʘ:��d�� �@�m��K�s��9šj�w��Dd��M"�AY��s��թ[�h#|�s�(W��Cq�/��'a�|Wv�r�9��Q"{�e4�O��t�%�S�*QY�{�Oo���l����}�wC��[�z��ٔ�]�b���!�`�V��ⵏTvuE�y�m���B�ső*g�-X�W��ϻ��;dtFo
m����6�u��u��^��F��������k�[Ս'��G�DmAG��ui���[�B�V�jY�;%����g0�KVՈ\�U�mܠ�U��Ov�d�������s�t����#:n I�ĕ�H�ٱ��)��lL	�h���^�����ҍ�[k��I��xH��N���yg���b\*%��3
2V�L��U2��*V�"�A[LqQ���Z���Vc��Y��-J�B��\2Z�q�7,p�
�ܶٙ�B�#m�,r�UV1��hc��"��Z��8ܲ�T�m�m��,bcZц\p�R�2".5J���������"�bb8�q���[L���11�Sb�Tb�4�ƌQ��ؘ�֥m)�+m���\anf	�"�".2��Ҙf)���ŉ��Z�n[mD�nfU��U+�Zܶ�p�Q��h�K���+e��L��2����ċl�!Z�b���&YZ�"�[Jb�C.f	�-�)m�e(�5���i(�%��0�K"�K��j�V�Eb�����H�
%LJ+��m��V�kh�m��i`����K� �2�Җ�[`�Vĭ�3)�����E���PR������**�+����"2*����V"�\��Q��Qd�XU���bh�?�(�8]�{<�6*�1Zc̦^ǩn�����H�7�X]�@���y�:�A꾴�Pm���L�X��9�ަ��0Ay�I�P=�n�t3��ZU�~�]c���Y�c�g�ڑnuY�J�w��x�Խ�)9ʵ�ܭpw���4_�^[M�^
޲�_Y�x�|�}p�Z�m`�^���;��]�a�m1�rىԵ�5Փ]�Z������^j�s��&˃�
��3޾���8���b�
��F(��+�d>�.��{����q���+�QP����;��ʹ�Ϫ��,��et�w�I���2�BM��.�{WφT~)�J^�����K��(42����B��'�1jc�+GJ����D�����zQ2�N�7��k|h����tO8�+L�>Xj��A.I�N�6�qy�o���^S���)ݖ�~͹��V�Ȯ���>q�O`��ÎPv�	������Ĺ���9�°��b�P�_�ò?	���w'�@,�ʽ2��q��||Y�̀ĄX<�$�#����ͯH�j��s�{�4-R{U��P�(��
^y�_�	*v/�0a��*��^1^U�e����(p.���p�0�r�:.���
�D㵣��{a�P�O�س5M�(k�#	�����`
��n��	k`i���f�д͢ia�EwS5v`��N ��PWvq��(�I�e�S%_�ָ�z����	7��chUR��h�/��"CC�DsY���3yg��Y�uz,�TɁ�T0��Q��JS��=��sw/�|3��GtE>�= B���QэD��ֲK�`�e�7��V��]�Fz�xTsy#�/�g���L$@x�_��ؙ޴�68)�|i��
�R�p���{7��.��l�M<�-3�\�<6-�8@S9���+�d{=�W->S��𐗟�{-�����z���*>�8��v��xR�ݺ�[b���'��'���P�K�2C<��xr�+�y�5��P1�cbό�i���=l�h������<=��\�Q^�G������%>�L���2�\D6�8���~^K�{���ʖ��<������n�#�q��D�t1j�b���������	;I��S��{�\��4�gY�N��nc�uv�0w�������^#���R���/�����|)Ď}�*D�+��"<���yA��N���eJ�r�~�FkZ�&T<�� t��ړb����@h�&ZY���(�>���L���ڮI��'���;Yy����YP��k��nѮ�V��!/�.�h��'X�m����q����m
ցB�}��%����o��n�y%��-�C�\u9�y�P!@hh�ܨ��:�`0�wXO��˰�-�WD�;���]�3�9��,kP�)��z3M��H��.��t��\C�����%��K�nF�_S�pW�X5afn�$u��q�N�H<��h�f��9҈ο����r�.�6�zo���y�K10��!�<����Z_����ؼ2T#+��J����/o�_N�R�h{y%`UC"�A2+s��Ys���.k¡�nY�*2��Xfm*�v���N�Φ28�y���`�.e�z$Z^�yw_�������dM�2�q�\˭;w��é�;���ڀ�P��X�-�I��pZK\�yϛ�US�\;���#�6K`���<���;>S/ j��p8)�$3�"��Mb
�+����7�=��_H�����G�Ⱦ�cj鑙�0R�����L�8)�\�����U�C\�ZƲz�>�e�܆voc���+�J��vq\�� ��e{>{�/od2��@�B�US��w���l�P�i����d���_b��X}��9�,Ҽ�%��wx�j���C�ب����h�v�}��^�!�ⱪ�%�gG���ɱ��vdh�W��qfK;~5�ҭ���T����h�`���k)�:��-I�O�bu�/�ξ|A�ꄂ����T�JE�A��Z;VL���qn�Y�!V ��s�gP:�Z�f�֎���}Xp��G�.V=mpϡ���k�GV��$��n�5�;�])�'����v�����=��⾣Bx���ƵD��{���åĔ>���\^�qZ�~g`�ه|;P�Gs��f�:�����q<yAr'�¾�z��z�})Ei�G{#�kڨJL[Ʒ)��[�ށ;�K��s��1��xp�h�!�z=wo5LT�����!|\�d�	�\B��>Q����F(��L&jr� w{ޣOE��	c��"�T�W=q�rg�&�wvtD�`�2�a��1EG[en)�艮�_Z`���,23uw���E�~#:�­Ԍ>��#��2$3�ݛb���0'��փ"㓞�C�ˬkͨR�:��l��1N�Đ��h��\��e��)�}�iL�� �~Uqb���z�����y�#���c����'�_E���4)�;�B���J�.k��3�3�R�҂�}�߭6iJ��Zu�M�yy;��~
fx��U1i�P�#�eø'��l�$-t��\SxRn�t@2���p�U�znP+��w�c�`þ{:��,F���à'5��Pɖ�3ö����coU��z����fDU�Bi�/a���~ۗr9���b]��ST!A��i���_@w�l4o%#`Q�}�w>�Og{�,����W����9CHǚ�����0Q��dA�+���
��}�`��/���KP.�z���b�O��|����Y�`�j>/�7ҒV�E_�f0\E��:|5&/B�NT��?;n3���je�+�m\�xg�����ޗIX��a��%꡾����N�g��iu��	]h���Uxhq�w�c��-�����O�\�3t�D\k���ۂv��ܭ$��-�^�r�����h�#گjX㆚�㶤VinW
��vsto<�3�f�]���w��>E���<��6?n���ڞ&��V�2��F������鉺Dރ���}�l��Z�ߚ���5�#j��C��V]��Hr�G[��wl�I���RX8�S�6�x΢�X*�s2ҟ�,��v8��y�k�Z��0;w�n��4D=�b6�V�kUqu���b�&��D�VzC�~}���� ��MV�ܗ袢�ֻW�'6,���A�yFD�򂸼왆�ȑ���"g1���}�&�q�Y�k�v[��3fkĄ0)��˨k�ZkE{�nm#�z6�2�Q3z8�:��&F����ln*�.��8V>��f���+O,i�]J�;]e����
|{v=�߬�n'[Β:���Qtƛ�V��V�@�w7��̮F`ٙr�r}�>���ԯ}U2��ߥ���(�$�L	lS)W���+9N\՚{���+��us������m�#c&�5g���zPv�L�v���!�O5:�~��	���@�Lξq�>~>���}�o�C�iE��u�N�,�g�Ō}�.����C۵��({��o��]D(6�d����p����A��_��Z۹pق`�t��(��{Eǝ6Wo���:�Լ��Ut����g��Y�3�)n�H�ǎ9F���6Ma!���s>������`�6�IW:E�eJ�*�m�ֶ)��v�ý*�桅���m��47��c�JO�T$�*���]��m�O[G�O�;�\7�K:�1�]��'[X-$M��݁�3EO��&�q�Hi�o�P��U��w�!\f4=��-����K�[a�9��\aN�_�P�C����xK�}W����߇��&j��[�^�ż%xdl��P9i�s�y��cr}0�>+I�+WZ����H�9\�L�;��:k�6O��k�>�`S^�Ԗ�66no�2��EZ*k�Cd޶�k��V�%a�IZ���������I��(7���h`ϋ&�Mj��]�B^�V�Jh�x�V����f_)z*_d���S���D�d�)���]heAa�7�c��4 �ϫ_�.���*:!��
��.�'�p�\��;[���Ez�c�sƭ�kT�����P��RxD躭�dŻ^�k�/L_����-���¤G<�Iͺfe9x �I-��:Y-���Ꞟ .����]q[�b`����SV)z�Ϫ_c(0o�q#�b�Jl��ܫM^����M�"	^��u��ֵ�eC��rJ�I�*6�D�n�uVvK�����i(�+�o��3%j�[�O����.��`-5���{������L"�z�LLWFt����_��)�-�`��*w��
e��G��f�^�ħ�Y}�̿rhC�x�Z5��k��p�������z����|e�F�C\}o6��%X>��i��M	"<�P��R�X�f4�d{��6&\�~�ï��������b���Io����X�\�ş�A��t�J��P��wX���;G�&�K)T���7v9�{",�����zP9.
�^��������S�2���6�Pd��ԏOwVd�o]o��0��|d�~y�.���Ϻ�i����"�g>�P&��=�ޯiI^X��_S �����x�=^�	�#���V��+���ֻfT���}�	��"���f]n��e�i�ܕ˥�${�y-�\
C�.���u瘧Խ���S/"�h�z���:���MA]�t��Q�Η�kY����z�
���xO	b���I�Ƭ�6�,�MY�GoH-u;�=ۇ��G�On�9�^�&o��%�G��R���(�綠���e=��3�1���F�{���0���}r	��v�b(�q��>�������ZLOgJ<�=�t�'��/=UsX����o钓�zW��"��ɏ�Äן��R�cҮ>����]i��e雫*�RR�F�[&�w�"�wС���|��;��^-*�"��¬���oh��4����n����^/����9Í�H�]2����'u���-l=5q`��-^�NV	H^e�����zl�����LŃl3���Ա�^���}~�y]#��P��g=#T3t��ua��ݯe�e�r�"�6,+\�J���|=0�Y���U��v+�W��o���/$W1��FOP�l�K�q�$����슺�l����M^�D��k�1� +׽�C8�r� f����9�j���Ju�=�!��ҳ�b��LO�h2�y{WU��Xe�n����(�}w�B�91���jJ�v� ElO�E�?j�8-�6����A�	��5���`��h�s��ɰ��ݻ=*���)�r��ܼ��o0����v˅s�̖I�>R�8��PL��<�yN���shH��o��෮k��:V��E�W,���P�ڸ���O%��e����z�S=.�`��@�w�z_�n��m�q�鶣Xt�O<�9�=o�6�_��D��5�
g�*�Rv��Weַ�������y&��P}������O���s�̢Y�d����vV��;˖����N�1��.�5�U���Y���FÕ�S��Y�(a��Fǀ��:5��}����È���/�x{Z�������|d��JD���V�c�Z�W�kD���]6JW^���h5���;�Vo�@B2�ߊZP{�P�P���J��
��>�l=���t'�����j^i�˸q���Ρ�U��tW�0�
ȼ��^?��S�� �7�4�.�����ӡ�ͥ6�>����0��e�B����;)��@릿{�Sbz�j����#�]��:�0�K�h��4N3�~Qen���a�[��q���G�u���[�Į
}!�k�w;F"�tV����*V��f�KN܊��z1��#�ĥ	����j�˾=]ڋ�+����a�S�.䬊�]���p2�d|6m��6-�T���2����0���y�`(7�Q���)���Vw��s}]�а���Y�>���Ⅸ%�"��.��b��[3)�>Ш9�55���8���[u:js��+Ϊ/�=1�D\��/�ŋ�΢�J����|�[Ы��Jgm5�#Ev��������"�u~���^"�JK�Z=>{��K�h�
�=(�$��ŷyhו�tM�DOU�O����P:�/%�,�e�ԫ���3�;�#�l'��\�ۦ%�s�i��pߛ��5�1T���pN5ܲa�֨�4�$�S@�\^q�}����,pD<mSٓC=���O��8RZ��ό���
�l�T�y��r�dMCƵ8ӜQ�ב�xUs~�����\pT�5yOX�C߹ƖƼTX�1`eB, ���9�Ex�{foLAco�Z���+�R��"y�����A�EB��J����L��{{(L~��u����\��t����G�(��S#�Y�fŜ_��Mf}���08j�!�$�3�����?xq0���P��IWJE�g�+�O參x������D���)B�����F��r�7������R?��f�A,�{��;�|�3L�����!Φ%<%_K���٠W&K�`Vn���M��M�]Yͪr}��t�SL��;P�իS3K��o:�'oV��h��R>�ifov��|����H��[�1M�7�����}Fm�F˰-�K�d�����g��z��$�G�,hO2n��4���N�ض0�a��g;���Z�k�5.�[�yR�:��ۭ�,����+^�e��PF�]�H>�r���u5>�z����ҋ��Ǟ�i8�k�	����/g,�g�8tO_�Z��:�U�)��Z%��B�B�&^V���J���b��>!a
��g_��L4׀�t"c����8�p9(�ci�4-�|!��ƹ�ǅ:�\�'T܆)��.UZ�[a��4*���ǸŜL�l��w��0�B��IvS�"�Av��f��$�ٚp��N	+w�4����%v�hqlYBf@
���9x��`��f��SVfu�*��xT���n��+�HE�����ՙ��n�2�9�
G��%*��ݖL��'U�gyhovMEƎ1y�X��ф�:�n9����7i݇MthD����s�rP@f:qT[��KTys�=�V�w������s��40uS͊���C����w�EXl`�v�+Ryx�%%���b��[&.���E��}j<��$΃�C}��<�Tɔ�֟qEM-��l�\w!�,�\��L8��Ov��+	��M̽2�S�j'p�s����Q7��c9u�ݻ]�s��]�睎�i����Eu��|
}�P��S�O�y���SX��*�ugk1� Wx�������y�Wq���z�kQm蹚ڧ�X��UêJ"�2W'�K�K������3����>�zM�pWƆΓ�rn�qg�[�Ȯ�:�N����+����Ύ0��y!��~/9�rl�'�;(xLd;uWj�q޽�\�Z�,�:s��;�<�.�Fu�r�������}4�p%5�m7�Y��<G���b>��ُ���&nk`�>ݼ��.&�wv�b�N��0�V'mͫ͵��IՐs���l��#S�e�M�Qqb��J�en�ڕ�`�@
R+lbk3)��<\av��!�O�a�՝k;PGK�!�uֹ:���~]եd�-tx��&lc344�X���u-�����GZ�m+�}�/��Jż��L8;x�t�Bн�]��-�u�~`�Ǭ����4�K�(�	fN��>R����[���p�W����@��2�\ki�XA��֏u���\�;B��a���Y��RN��t(�[��t䇊�:�"�����t�D�W�PCk��5�f�a���y�t����*}��]Y��/7��ӈe�<4�#��J7���R:�< ��P�6m.�8wa���]�r��<?qОWs�f�z�BWK�![[���ZQ��_48�݃�vk5�p�&5ƪ�,EQV+�[q�"(���(��bAA�0k0̴D�ƢVUr���Kl�""��6�)-�����cQFE��1KJ�X.f`�X���Af5���QX��Ȫ��ij9�C�X�cqX��KKh
��ƪ6Ԭ���jV�Ym�F#
�ŊF5*b��R)ұ�*���,+L��dR�V
&8����
V��)��rե�(�j�
 �be���VR��X��
�`���X�Er�VLea3E1�Z*
��*��Q�#1�1��C(e�8�˙�"����Z*���X%V��QE������0�!�X#��\eE�m�l�3�PQ�aXnP�E�P0Uam1�㖘�X[QKj�X.U���,EU�Z��D1
&Zc\aE�2�T�1P�46�nW�=y�y!���zb�ݏ��.�{P����^����>Z�]m`��Gk+���r��ݥ�ul�>�MDfV��)�Z�C�^v��:2�&�tH�6����<�ZI����WR�#Sk�4�K:ў�u�v)H�>���c�7�E>�Mjf4M�i�o�>�U���<�L���92�ڡ� Ɨ���Ge���gN�3B��SeIRo�3r98w�lg�Ї�}�]pU��e@j���R�Q�k���׏�>�aq���Y�����0��E�@���iw����0����M��c'��L����i�������Un�ʦu,��2���݇r�ˁ�ۄn�w&�[t5>����b� җ��z�`.�>�?�����a%��f#tH{Ŀ��S�n�jy���i���A���αҋ��SWK֦R���(0h_
q#B���	
-���Q�쎊��[iO��"�N�<����W�9�`���(3��M6m�L]�����_V7������ǒ��)��ل��cZ��)��xFi��L�zĻG��5���pX���g�s�g>"�Df��d���Zl�=�f*��
9�ʝ���
e��e��ʺ�ڶq�|m�G������u�;�f�	a��ם*At�ӽ��y����f�������[��hL� ߖv�Ԓ�Fwq:&��B���Gu׏��6��+\h��2�Q+�W�vԌ��ƻáe�3%�ۯv���ˀ�����ǽ�����>������A_��Z9s˔�������.*���?7��o8o��lSPL4͎�@��J%uLưPL���a�ɗ6��{}o��<uY����o� u.Y
o{$���~�{��
8-��, �<�s�8��xs�M�k��GOO��>
��CM(��^��.t�&��R�\-��}�k��r���B[�I
�rWN��5��t�	����OE��ܔ�-
W�ԞV}��1LP�U�N|�����ئ; �5R�����<�
����o�T�5L�Ƹt���+r5dJLpSԹC��Y��'33�R=�)�S���.�&�e��Ƒ�2�P�����C7��K5�a[ٌp���<%Щ�I��g�4�.k~��bS=�Q�CWd(}p-�F�´�&��>�:y
������^���5�7U�v�������Ä�3��Mr��k�T.����w���:8Wz�e S�e��9 ���=��C �s-�k�51�=���5�"b{����ל+���������]:�Uz�ׯ&�ݻ aW����|+e#��K:tG�k�Ϋ�%�V�k7���z��*܁n�dR׫$�u�����>��(pu�vP�bl&��6��P��Y���d5��2����k;��������X�{M��xU4�i��ոH��L������{��cMY���#�Կ4/�P
m�\��]Z��:��lzj��3����u.�yNy��,c�Y�&�lJI{���gk=n��\1kEb�;�C�l>QgޘL6���V���Bm.��^���ƛK|:l�:���@�:8�F�\dYU\fv]�K�����M^(�rs']��Ճ�ļ%w���f��8!����ݭW��E�+��(&&W&H�V��3�m��%���+[��q<s�Wz׸Jq�CY���P�ڄ�%RGڹ(	��ߨS2�z�S�_�\�����=k;���PWz�9[�A���F��P�UE���4)ۺ��}c��P*ڇt�z�IW<ˮd��.>�r}Bt
fx����O������3��(0
Ȇ�y���f�7���ʂ�����q��R)�s��E�q�+����Vxa�v���'���kbݡ���NB�.���̼���f�/��Qf��Iw�T"����i�TH��E����4C�3z��Z���\�ߎ��W��JN�	DV�Bh����*k|���/���@u����2gY�u���_�C��ox3�짶�h�'��u�:8�k�Gv�KW+]�g�G��uG�W�'����R��眳1wulΨX�/&2d��K��& u�컇�yND�տp�>3 �)iA�]vz�����x�8���OT�������k�汯%��+��L>ʭUxi��R�.���<5�Y1���.�ΘS�)����a;��w��4��t�Bx�w���3�^z �/߿{�[w����>^�]�~�U�4G�, \��0�%�R����i�;�1��P��e/zH_iy��z�(2�@_��A�1u;HJ����yj� ��[=Yޮ[���f�W�g��W`Ll����p�]e�b�p���E���+�d>��An��GjV^Vm�� Mh�r�+E<�L?��=*���ϒZ=)��K���ܥ�����lR�$�7�w�¾yE�َV�E��ǔd`f�|�	m��b����Fs-�T����ϋ���R럈?N���V�(VD�=@��|��ݗ4tj�F݋7c6���Z��_z,���l����o��1�ÎPv�e#���"��Ra�����k.iͬ���0��KB�b�݂.��fj�9��6஛�hp�dt�T��6�k��xy�B��}�Y���g��+=��K�
�d�9��-*�8aK%V\����k�6]ZQ+;DY���I�{��� �wr\����$�\E\���M���R���Y�>]��G���G�X��q��TS�U0a� Ռgpc��]�c���(��0�!"��A�P�)�Sx#��^y��K[y��9��]79��wTn?/]��#\�4�du/��͋8�t���財���b:�;-Q�������]r��i��Z9К�`�ne$��"��T�"��ٿ�bا��k�=��Ӈ�������ߝ%"�T��(��o槕���J�d���.��K�\�f_���~�0Ľ�܋�q<wM����,o�<lզcDؐ�$����b`�Z�V�N�fM��T�u�K��X�u~B��-��[����>�q�8���낯�*���y%ׯF��L��nX=hˀ4fz��
ҙ5ֵ�#���������O[=�P�t�Z#vqN-�������Kr����QP�Y:�ِnW�������3�H�=I��^��.D�7g��gt�jx�\:Z�ly���q�ͥ�#�;fn@L���./̝����W��ͫ�JK_<��O��b�f)�=Ƴ��o,!��";�n�X��i�t�V��\ژ!1��xkK$���z��7��-_H-�ӷ�����M��r"��K4n��Q�����U+z��B�IƇ;f�g�3)j��b�z�ʝx�RިC>���L���VGMX�j`�|U�t�wn�Յ=bs�&��:ċ�]�A�p�u;�u��FkZ�����MlԞ�=�p*!LI2_�	�y{TG_c�T3}�	��K�>S�����k&Q��1��Cce�\}Z༝��I�%�8�^q��\�Vf�f*��
8T�W��S-
ޞJ
�۵�����x�f��%�$��O&��Y�>a|=���9����(��v��ש.���p0n��������5ΔI&c[��h2˞�N�]�w�=����0\*8G�M�B>��mKB�E-I�����5��H��S�� �]����㛻PL��mt��=]4��9�>;��yp�j��(e�ʄX�(K�<���f�+댻�fm��Ҹ��/[���|�Jf���]/��[�F`S.M�
|�|�>�TC=d��1���/x���ݯ
�R��U�����h�L�Ϸ�
V�#Vpi�oԻ	�j�ȱK]N�^�e��Ӓz�\#xe5c(]R�;<Y��q��:i��Tk�]a�B���Q�b��c�2��^��oq�b�S�����s�{!�ً�L�ֹ�B�c�H�]�r�s�iǛ/D��>O]ve�$�eیl<g]k)B;�t@sS��ͫ�EM�y~X��1�{)��zg��Ξ!�zX�\����v8{|��u>�R����>w��N��E�7d(k��m��2	����S�.���e�h�iD5�w�O<ʝo�����p�x�o�^��
�����\�zU���8<_�K�J#$�2`�����==�ɗ��˲7��P���n�S��SSЎ2jd֨QI7Y�Y{�n����C��Q�x.c_'.ϧå��g���Z3i��Yh��������ѾZp�t�H�4�B|����z�;��zj��̱N�(|K�;]ūz�
�{!/��j����r�H�/��[i�C���,+\�Jǝ��L&g({�U��UD�2R�+;K�g5�OLN2x1�ྲྀ�6
�"Iq�;.ȫ���+9�������zm�4���wŬ՞�����,2.Y����au"��WPL��<�yN��&���5���흩s���6�{�>ZfNy�~z��b�ڸ���h�j�6��y�L�3h;�}���Ib��^��X��x�fF����9�󭸺�}eP#����ܡA�y�=��U��d<u���hl�|9g����Y�咮�T=�-8����Ϻ!1;p��
��D-�ʃm�TMUM�U
(@��sV�y�q>��|U�*-L���8�o�ۉ7��=�}S������0Ƭ�𞙜re;B���F��[�g�k�����G�S9SW(T.�\�zR�5���g�x5S���F]C�z�e���U���M;���ow*0m�GZVT����φn��zJMf���ȃ��]�^
��-���pT�pCݽ���sP�CEl-�Vf:�5���H�r�Z��G�Q��]w
cϳ�7F-��tؙwıMD��e�>�P�ؓ*��ʚ=u��S!�|r.f�7����i)'��+�j^�+ܻ��y�S)1Z;(��}|p�|[�gL�O�jf��Jk���Z&S�@�O ���;
�����O,�x�U��~~��s����R`��_����-Ϋ2�-	*���AN3�iE���KXc F�u�Ϊz��pk�ieӐU=Y�S������l���fg��b��\OT�P����/v鮞N�UV�B}������3��a-z�mM�7�E��T!�n�d;2Y'�բ�hm�r�G�vK�� +�;;�냒'�`��;��]5�)�*�n��v�A?��D��)�-{��v����O�]��O+:�Les7�B�G�d�����KE^:Usz���X�6�A��۰FɒՆ�6��tA�J�:�
m�7+�U�%p�9:�]L{�](u֊�����"�J��>2�Z=>{�aBN�d(g�3�-�h�{��V'��︮�=���.�\�TBv@P}��:R+GO�z@��7ʱo�:���;}V��7r%̓���P��fY��տ�(/����i�{βu����;�܅<aJg8����!�Fy�F߫yYy�xr(;V&R;aݠC�7ұ��<��c7�K�Dh1'������Su<���;"���Y��c^+�1��'���,��k�=;�N��4��&����W�������S7�? ��p�X��Ἇ{f��.phs\��Q����\�"�+�&��2:����W��v��A��_Rt��x��-鳝�Ǖ��Wc�>�F֌X�����ؑ�J-"�ն��[�Լ*Pg��t������}�V��]%mC�.�."F���˰�i&o�E�tU�%� &�������$�.�=Yިt��ޕEs�զcD܆��3yP��<�M}_I갬��W,��]�Tƞ����w6S���%�f�̫�d����\�֛S��X�Gvz�J�;�w��hˬ����1���Ճܳg^aN�M��U�����J�54n��6�=��H��S�\����B���F�#�iqI��YQ��]<��=�+�\�;Ԡƫ�ڪk�}�
��Z��ב�m���nV�ťwϮG�l�t�A�ЁT_��{�f[�x?r�v���+Z�,:�|^�
ߊd�Zל|�}�)OA(!�'1���d�p~K}�鋹շ;9Ol^t��sUdڊgR���vd�r��6�tV�2�{ܣ٫����dr-��vK�}��8j+����%c��\���T�^��|�q�Hd��^��V���ے�)��<Է��w��X�Yj+��"�߰-?V{e�.�=����_����
rFy�q,���M���ok���kY=U��-x�e�+��E;����^p�=�f@h�ؙiy���L��Ƶ�
u�^3M��H�׸;�G��{�;xu��xŦ������rf�\��3�6a"���q�N�;6��Y}յ$Mc��-�#�:�_s��
�	q~��A�.yp�+�*c���|#�:���B�q���nI�M_2�]c/`Z�h*��|N����a���B���s���$��H@��H@����$�$�	'��$ I?�	!I��$�	'��$ I?���$��	!I��B����$��$ I,	!I�H@��	!I� IO�H@��	!I� IO�H@�{H@���d�Mg�nU~hAd����v@��������р�Wy��׮�ia�`2
P=�z�j����Ӻɫb��{W�a��f�[��V��U��}Y�l/��M��Ս^�t��/M���kV���������U:ԉ�Ǟ��5��i����H�ޅ��N�^�������{�    1��T�Tdh0#4� ��1%*�       T�L@���& ɀF LA�~%*�?T� 	� L 	�S�J�% h �     $"F##SL)�5=�i�z�xS�I��ҝAS��ԝ-�����p�
Ԣ"� ��-"���%x~��~L?#��n:���`@%D�_΀PS�d�]b7�Q��)�=Y��r�[��~����l��Rib��3��D��2�Sۑ��IF�@����Q�Ԓ�Z
�6��K>n��O��jơXʡx.P�.���wP&Kv�̢�Cpi��݃��Qʂ
�v����]�@�X�VkM)C�-2**M�_fV��H斝f���o ��m�������̭Ȩ���b��LD�%n���e��a��N���7�Z����yx� 'Yl'R�,��C(�S���v�R��V��
�xi,Y�ą=UɈ�]S�l�bD��t�"i�V�tq��u^H�L,3lS���P4��&^+.�hM��t.V;���,��ݍ�0YA��O����$5�Ֆ탭kR������ݭ��eT�)�٥PV�4l`T��e�����N�.ʘ^:�2�(��CB^&�,6��`�ѻkF�a�Va�+َb9�!P7,)l%�V�kw)����wn�j%[��;a���
`�q��H�1�;� )�b��wf\٘!����\�VdV�=B��TBT��-i_\�d�*v�qTG\� $�2�l�/Q�D�^`�J��a���K���8��k�04�3T�c-����ˑcg�7[*n�������N�ke'�T1���˧D��+o*��3�;Tw]� �����E:��Ν�U�:Q�fMx��w{jO6�zt� ��u�I�P?3K|��X������_�gG&q4R�� R��͢�@��W�]M5��*|J� ��*mξ}ԲSBv�}\vVK̾���M^wO���������7�n���J;�����͜�ۙu�	��&>�|H�Ӎ�Gۻ�՜��At\s����\�uLޢ���Ꮾ$�}�N��X�k|�"��Ճ/&�J���2XDXp�𤜺�IX9r��g���d���9�x�kٕ��.��]�p�{�4�}Rnq��\���V��:���SCuոD>�����\T�tI�-æنK4m+�Ae��t�\)w]λqL�}�]�2j���u�����Q�ƛ���Ac�C "�r
���$�����>rPɼ��D��hʎ�����xҫ�z�{G*z&7���fU� �2����E��PPuN�K���K9wt̓���#�6�]0�Z�Ć$�#Wt��N����&V�.�#�>��R>�r]Ǐ9��m�s�{)�EWg99�:�;��S��'s��\�v� �qu���"���uYB󌖵¬ɹ�����/�y���b=j����wl�:�t�:�S��e;i�Y�\9�î�S�I�3�2��c�J[�{�m9R�h������9����J���DF��5N�1r!�ٴ���;T�I}��m�o�o_�Y��rߪ�ߊ�|���!�-�𨪜�k*'�N79=�`P=���g.�	Q�6#i��,^ذ~��ɇ��� ��IZ�.�{u�B(�4�l�&%�CLK�ҙ�/���p%[�&���q6�L��(q\���!��X�EJ�z�Uf��m척Tw)��oT#���E��:�zn �s tSخ��g���9�줸@�{���j$KRW��H.2�K9_D�	kl��ֳ�互Lf�}R1Hd�i̡B�A�	\� 0�Yo\Օ�$N��;u�0�#���Vm�Ӑ~d(!������y�,���)J-
���Iq�C�+�5�a+��ֽhbӕ��!E����@3G�����H$��d3�6��� ���7h*���[�j&���:~�� �t\���D*�}�?]c�to�B0��\�ƻ�v�=�tK�5��l"�`й�@�b��D�p��-�r��)w����5���+�2�?�
a�C����t���&���H�;BiF��I5;�d��N��tzQ}�&3N�t�N������t۹l]/��O[vi�B�aR�/L�`tXt�e���e�%>2L�1t��Cjb���EYc|�l9Y�X�B�X.խ��z�_[����
@��I>hn���%�<��/�^8��v�{�¹w*��3���f��g�k���O�B�	�I�^&�`-V*C��e����q�91%���!�����u�ony��`EjՌ��E�Mr�]b ���}���@�t����;n�6ok����Af�܅�����p0��ş-��f4C������;}����1(���	wf�
�y�:�@|f��y�Il���*r�s(�I��>�+���2��Ovf��$���f$:��V*��:�C��B��L��(@�H�|�I��1U�W�mv�vv��ws�@��n^�i�Gv�q���D&�����>����Or��Pi�_�xny�g��=뱉4�t���7�փ�=���R�o���|0 ۳��K������@a݅�*���f��H`�	��pq�G���TȎ���kp�r��}x��='=f�M��,���oET/�c$��f���o��6��-��'9-l�xV��CU³J9֯J��ӴLM�m�A��F��P�f!Sx��4k{L�Đ*$� ��)DF
H7A�!�,��"�ޅp���٭g�ҹY�[�r3@D|����F��I1QI�{7��b�j5�h�&6(mX �*8�!��k�����/EiFe�y�-�O���F����g��
A,��{"�G��� �>�Lf��4���"^8�e�홬�fj�aom��ϯ^Z�ϽO�����pz �a��dbB�Ś�p�,23����/\�y�U�]#h8�дw֖�4��i�-5�b��l�?KA��$}��Yʏ�D|	��g�dC����=��k�ǲ]��U��8ƃ6G��������Qm)qC:��& ������Z�g�nx���xXy�x��jᑝ�^�ۖ����oLu�r�^Vp����WK5啽w���T{2����hf�����o���f_�>8b[��ܛ������)a�M,��ra���麝���X�R[��R�us����.�D8���p�V�MDn�o�,�:ݻ,s0?ʾ;8'OI+dW�n�5��u�:�]Y��rf��jw(�kČN,�JRp�2��ĥѣr�������xA�#�D���Fq]�߿�^�{�۟R׋�5j�Ι�������<m˵�9W+#�oa/��;A�m��̅b��*���$z���)@�|��-�m�,�dxg<N�s�/nw�dd]<�r�hY� s,I37*��_�o7{�s��S�'/�[���M�kmi���u�w��1���h53��cJ\�
��̀�������}��Sy���k�f	!�4��Hb-�TC2��#�Y�V�0/�r刁'�;���3��ب�:�(��tE��?.vHz�-n����A�`�^ہ�w0RU��+��o滿y�uD��CA���*�ˌ��׿,hv+��AN��]<��(I��Ց�:��\S�e�䕚�P�T|,h��Я=y�Ԙ#V�mDc:���V�~�5�wm+�d�j���Ͼ������w��Bs��ҘCإ�@i-'�G;9C��ÅKv�]�09��ʣ6-�]x�b��DS�VS�O~{lO���Ͷ�s��X�C�X]@��a,!��ꭌ�B�e6�Jr��L_����_��\��[�NHBnlT�TO��ѩ-j�NU�q�lV*xݮ�������x�������h�eO�ii�5�PvW��jDN�A�!��G�Wg���v��nļCG�ge��<�q��4jߵ)l�I*��}�kN����u�9~{��f�����lI�[7k��o?z�u2⨄Y�Wh��j|�j*�Hid�pF6�5�=X�Q��LB�ب0��YT-]Ŏm��昖�<�XwN�W{�N�Ie����VM���I̚V���x�N(p��˄�I&��Y)IP��}���+�;������Bā� �S��bH`$&C�Bf����.9m{^I�O#L�Uk���f��8]�6˫E��N��EG����2�S�(:A���4���D�**b
�-{(����S1o�Y�L���i��o3c�������4����dS�(���K��\kf�i��>)��e�m7��� (5��;�WڒS�5�<��a��G�Qo-vщg��
ĦsպｈT�]��\��qQ9�B�u{[AGpUL�'^�T͙A�3���S����Vҗ4ɰj2�K���^���UX�|�L���(�EW�m&]�[�`EÛ����W���9�����n,�:+�0UYIt��|̏B��s#��l׷�����+�|YK�vu�AuT1�-��׳Rˁ����{3r)�E���v�|��	���o�wMLWJ��U3��Z�����g�o�s�s�Ro��V�����]1�u�&�!�!VqÖ"��Y3a��zkϕ�;�����X���?On-B�p�)uX���P�ӛ5�:����T�=W�lx�>�p"�x%Mk�7n"�T��;���r�p���������ít���V)���M�EL�{3�����(!/�˻нS�OB�u�����)>a@���:��ʙ��WWX��:�A6�*�%JEC���*�S9*�n�������HXFH�e
T>]-��O�m�O�+��s��S���;^����J�^�{�+�4;���vi���NzNh�{B^��7 ]<��YPmd�*oz�y0�TNc� ����;mՎ�˩cow���u�7�v�p|�/���m�o^<2h�ʂuZ�\;�0�>[��y�\k��E�ʶ6�"�!Ot�C8d%6�+5�$�u^�gu�`M���O�0>%�fG��^s�x/t����v-��R�����{��>�q����I2i���;��#2��{�'|�ݦ%�����4r�}��Ps����������h�-hٟ,D�[��`���yK��u#/����PS0if�f���}���"�ͬ7I-���&r}y�Ca4�|SURF�H�P��nw"�[y���`w��u�}f��~s���{�|N���1D���t���C�L�Q�@YŊ�k��}��l�ڠ/+Hzz�٩�ʢ�+���YD{��
�x��RI�N՝��p ���R�k�Z���kw1��"�mp�\{Evm�B�G�J
)�pDs�Z�Eȗ���C�!���!y�-QP��,�2j�saVm��ԙ�	��.wv7fc��Aı[,
T���M�0�B�y�ny��#������
�C��}�����W��/ے&+�3uW�Fc�BE�jVoq�T�N=4U�ST]�����ffg�x4i��v���c�v˩h��r�=`��Z^`��@s�<t?wf�YKUU�{��4|.��!��]C��g+m��۟�������NXlI�Ԕ���y�y�8X2�:]ؽq#�u�T�`c��Na�2�>*;�WAN�������������|{���ޟ�Bc�]TK�hkNM�:X5���LoT���]<����>�������ܨ�ǲ���:^t���X'@g��w�!�j�wA��T�o=-*�V%J�sy��4��P&E�4.�b�U��*lN��0�����˪y��"��-o���}��������Ct�GZ�nyCT?pB�Xl-Zof�֘��x��ud�^,/��o{�?����D�.(�A	���Y@{3�'y�s�
��0E9���ܵ��0�����Lt��g�$X�G�#oX�U�j�f�B(��2�o9h�.�M4��ˋ~���WQ-�{�@qbp���i �f޶����f�Å�
�C�Z��|w�v_Qy��Pt���_Z�x�V�l�;cx��R�*�8
Q�TL���d�	),��B
Rg�e ��ޮ�(w��G�|AE|�H���$J2123Y5j-�e�ћ�s���j�voy�������5�)�D��|�� ��g~�c���#���MR�#�<�So���� C2���+��?{��w�s�8�e���\�ɡդ��d�iX��iW��_7��822���_8�K��@����a�b�>�lP���2�̼Նo���<+=e��"����Z�2�q��	�ٶ�����U�Yb��
�������Ο�S�s�%�7�0��s���U����L¡�Y�y�6�ҳW���k.{�U���*�ܴ�5���LrM��쾚��g�]M���R���G��O�|>o)����K��f���)Vf�w��<��x�>b�}S��/����Nyo���f�	�L�zv�PX;�0tӾ��dKs\_�$j�iө��H�F)�i-�Fg@{Uz����=����}D�p/ͣ�N�����҆�,���rw��vy:����[�)��V�Ɣ��ｾ�?� ����L�U�I%���Z�[K�<�z��+(C�駎�Z2V�K��1�Y�Nf���<>�޵1�Z��ޕ����G���h��A
�ѕ�\C�𕕕lB�E�7��uo�z���%-{�Us��g��Y�`�o{���N>��^Q���,�i;��T�Ħ��w�YIO8eY'/�����%�RT
�J�P��T��P����j"�,�l���<���{V������-�H�!~�������*��lF�B?:ԥ�Yq�o���R�g���֪�2*ʵ�	��QGW��c,R��3�Qt���z�G	OJXZ�EC�w)O�K��eM�L=��7U�m��A��8�
 xm�Ä�L�=1�j���H�d!��i�0������8��v����S���a�,4R0h>+��e�^���X`��Pmঌ�T4\4vm�A�������s�_a����/b���<n8����N�)��ڏjzm�-اʙ�
��r�ע1o9�jd׫e�>���(�Q����^�B/���0�]��j�(��^�	�$Z"�D4����o�+�\�2�Pt�*��H(�79�{����Rp��S�<�'�OtV�#it��]Mi{V�l^:���QT	G�g�TYl��=���O�8��=k�YC�R��)�Ș��|���cr?z�V�Bz��s�{�W�/N7HLb�,2�VhP:��:)�;�����e{nVݥ��K�ô��>9���Wѡ��!��f�=��Jt����N���~��*���bz�j(2C �8wL�o1�n�nj�ߙ��z�չUo,�l-�hv΁Ѯ1,r�[W�ܰۧ�7�l�v��|\[��yW{�ќ�R�T��s[$]�pb�K�BI�ZXqe��J�R����*�$�M�[�F�ԅ�nZ��5n�L�L �V��&j̀ �/������uʌ�y=��j��	~��T)=��&������N��}�	� ����'���n�w�۠j�S�Tn��8�G�{�BC��A��QÕ�2Ƽ�d�ɐ�<�Y��v�j���x4uZ8�����iTҝ�m,a;>�s��Q�&���{EU >��6�:��vG����z��z*r�ZX9x����|a}RV h#T}h��L��V�h��=��r����.��X�^�)@>�6V�u��ؐ�x�9����1�"�"�'R(��Un�YV��-�:x�o�Ti�=�.�{۔D|Tn+�^.{���s"�O �fm6JP��%��0����zMV�o�js�x�c۷�*֙��h+�x�����lu��%��@;�nN�S8�!������zR�ffo���"�#�N�韉�|p?�Y=�;��&���DO�/'%)����d��we^դ*��]� =M�<Z6ݡ|UVԦ2^¥1w�T\�O�/��YS��Q�Xު���P���X���$p�w.��V���{|��tR'���7h@�ؽ�3p�Y�z2ыZ���Gwf��O��k3`�z��!o�ѡ
q�F��T��c̸����w&蹍a��T�k��b�ГI��m�^��ժ��7Zz����=��;��^��٬q�h�B������L��kq2�@�֬b�JJ�K7mլ��
J+�1R�0��j�)L�T����`�d	���Jb�-�F)���0�� ntΎs6�/B�ߌhnxU�"����v��<y��~|�m�HzC�Ik�;�]�N��wMl����T��>33!xdF���V�c�t�恧�A�7h!�������5{�.���N����,�bj���S�Fz|��!|T#��l�v���{}�ɲ�Rv��I&>~��<]���h�����Fx\%k<8]����XK⛏�dx�_��_�>qؽ��wsvNj�p@��dFr����j�V��&w0�k���u��jܽ���v:ooe�m�C;F�(�yQ��Cxi���>m��s�>���$"#*b�D�LC[�hMY�
��pջ�l&B`���M�m:����cMqE��y��"r������=�r]��'T����v���
���x5�g�޻9
G�W&|x������B��w3UO����wM>�Y1��p��<��6c���
��g-T9Ù���g��#sr{��mЌ�1C�[%Rg�9��yʥj7���%>^i�BV]{��k2g��������8����	���Uf���֐�\��F!e�l��ycۓ�՞uV�%J��{�P��T��No:��s��o�s
r���L��>���`u�@^D�Y��ÌU��U)I�i$�vN*�����ixhI�H'������5[*H�[f�ł�FZ��Y]u�Ϯ����L`�2���I�dVC��7�S�[g;A�7�z$m9T#K�|�;2��_����ڣ��1S�l`��x~���M,���?��+ڴ�9Pԣ+�������P�H�������S���O�1���Dd��}�,�Z߆�.]�bCh���)�"%��^��B-Vv����U�y����y�{�f��h�`���uʱ���$tk�v�
��v�4Ć����r�~�r, s<�N���Y�	b��Z��g�b/]�_�:�,B�:��<��H�����{ͮ�h��`4<4!�!ŧ�&TN��=T	x�簂���T(��w� ����A �iy�/w�=v�}�o
}��U�<���*9��*t��M�����Hٵn��6�_Ő�w�{�OK8��]����B��0wrBI\�OFw-d�o��@̫>U�*4�,�l�yPݐdݝ����cnD� p$�B�@���IA!�p]��Y��X��+S?�Ζ]���^��ڭ�]��4��W�~P�U%w���rc^�TZ��51!B.*�':�<z�y���|7Ӳ��Ѕ��������G����
vPN�}#��{�la)/b�fo�b�>=W>�K�֒�C?;%�f� )S<hX����e�2�9E4�JNQ�9����(>�� ��NsH�f��d�;�|��{Rۼp���sA�z\�:)פ��k��Υ����3�)49!0Xx�æ4o�Ȁ)����|v�O{>`04C����2*��z H��<?�\�N����܃�連������~Ǒ��� ���ܠ�� |+�,���A8��C�D,��/��?���\!6�V-+�ƫ�l�������	$ם���)ռH?�
PI����j���$;��ʀ
y��`�^I�E��*�)V�����`|�s�ؠ�����v�����C��o��+t��I��Ӳ�:�Pzu�ˠ�����4)��S̴ӽ3�Q˼#J )�[N��v�9����u2^��Y�;�@Rh��¼��L�=I�I��C
T�N�C��ܐ�3���>)��x� �Q�E�5����}g,.��[jQ���G�����Id�� �����U���/���������M�L
�0���(��v!��K6']� �@�\��t���bۛ��2X}SDL�Y�hF�Z��C/����.�6Wi�=� v�A ������O��N�~���?w�� ?s�~���¾>���������w������"{�܉�u���F��� �����Y�;d�TP���������@.�C@��I�c����o#�O/���'������4��J)=��lA����	��#ύ��b'������3[;n;	�Ԝ� ��tB���gN�-λ�e5!��(�V�ϱN��
"r�N��n�������,�[�%��C�>O��u�z;��@S����$��d{��r��2���ioe�+[W�	�b�<x����rE8P��X�