BZh91AY&SY�R�@ ��_�ryg����ߺ����  `]?}��  ـP6�=� (   �1)T,x�)��=PTQ��.��1P)MM�N�������{�H��� ���')%
 �D�@t�I�@!HD�˰2���m���-�J��Ǽ$
f�
    @�  ��  %OH3�UT�MF�FL�M di�j��D��4�  ��     p�L�i�FL h	�L� @�i�IJ�FCC	�� 	�0 h"DR�OP@���b   
�!4��h4���OL���=
m'���i3�Q������k�Hpl�2e�D���?�"�DU�b��Z����_��$$+���I���?�?���������S.�����8x������YUH�����$F�;<�M��1m�1�O���	��<X$����Ď*Ŷ�m�#��d�Q$I�G�G�������������?����_\y~A�G<�a�/LF}��H��1����R�<�S�=���^��8[Խ��s<g2�� 97qgy:γ��Le��^K�U9���s���a�<þ��zs���Ʃ{T����)�ˏ�����V�<���y�#�1�:��ʣ7QL��dL*�JJ{)�菢>�I����VWY]9�U�"�T�VzDj&rX�#q�e�'nRqeY�ex�K�*�uڕ㛛0�tԤ�r���H�G#�1�u�*�qet� ���:��"m�{n[r��D�J1�u�9���eP�J�����Jw6A��'����%��&2DS�gi����6U�x�����Y�t��t���Z�����nC"d�1=�K/�D�I��dd/%:�+u)6�Rm�I璓JE�X>j�,Ͳ�3ݪ�K�J㒹z�{^��M�������,�5]�i"�e��5Z�+^;���9۪E���U�뒛�sV�nX������7)��%9���2_�%�Iw$��C�O�%O��R~�
���吏x�z{�Wt���<n����
�� ߇};�=�[�-�{uK�W���,�Lf`]�;r��܃��:����N�݉g�OA<�����YNi1��}+�����'f�	�:�PI#D�H2k$���L�J�͔�Jr&���3��#��øɑ���UL����;�*FFFFCc���rǓ
bV5*ڕq*ғy�%ugxw���oM�<燜��'�G��98]1��ꒄ�	�n�VV�{ڧ���l��y6�W.s�p�U�Y�u��g�����/��/d�D����'JG�L�ZL�c,�Y]7q-ew]9ru4ȓ�Dy�G�-��Ypt䤬eY�2�{��<�<<(�}>��^�^zUǁ����v�go���o���:�Ժ�?K�������Hγl$x�g��O\���o�}��G"ͳo��1���y��1j	����+}SN�F��'�;�k4�E�XD��ӡ�2$N<���Hɲx��~D�Gғ��'|_�#�0�rNsl��8����5z���������q1ڏW�s�r&�i�1�Lo��ɢ{�/�5����<�v��Z3��o��>1y��y:�<�/�;�]of��o�C5c��,�]g��$��_[eS$����w&�I�Tq�}{��cg�����.ߝn��7�\%MϜ����V�[u'����y�����8y�����-����ݥQ'�i��ޒFG�S7�c	+�-x�	ën>�A�uPlm93+b�t�[��n:���ra���l�n�R�l�dx������~�ɫ΄�Ttr�����fa��)Ģ�(qs�B�5��Jp<�ɓ�k����� ��Pq�GhV�J�:R�eTZ~6�6?<��u7�Ӂ�����٧��+>Sˤ�}~�[p�Y\��a_=\��y�XE�����(���e�²B�}�Ep�0����%�1ݙ�ᦈ�:��-p�l�!{2r���5X����2<�z��(�}]f��&�l:�|��d��ؗ^Qb��bR"q�� �=<�q��7{Ǌl��	m�[����,�:t��\�R�3�q��z��m�顀��6g���� �gV{��c�_z�Ѱ�'���1%p�nf�YҙM�5�_������/��<���O���8cH[��źբ4���2���`/0�BE�a2��	e2���W�"3=�p�`������I	"\�O�Y�|kD��,��ĳK��!&�M�T���h�G�b��|�a<���6�r�D�����]��+|/���)H��.BM�n�m�T<�
�����4O#	Y*7�ģ�WU�C�4��k��:�F���������B�y@�c�˶dI�q�)+s9))L��������ڡ`�{¬�|�wwu�w�n�m�
	�/�EgLV~�n�ۂp�C�:�df|,Ҍ�ƕ+K�G�����ˌ��7���c�\�%�{��ߣ��>�z=��<Ro:�ǡ.��j���`��[��ANT���5�W��c�2U��f)-D�!d�i���7l�p�c^�{�b2Q1Y4#[�,6(��4��*�Eq�B��8XI祴ì�z/�ޗ圃���%��)Q��_�L�ȿ��~�� }ħͻ��Z�W+��+�����j6{'�����ϲyz��N���|[y�9+�b;�׫����3��D�l�ڧ�ey���h���s��#.��6T�ێkr�5���:	�mR5S���H9YZ���g��f
j'*��*��'� ��� �D�'�5B��M�Aea��7R(.�U*�	���j�U�b�����:�ύ���u6ӕ�B����Q5���|$h!��P2B��P��(���"'�N;��Ndr2Ln�r���L��RP\F˭v�Qj	5R��2Q(Ƅrwq��H�m�)]$<�I�ʭv˚��\�I�6�aH�E�#�"�#h��Z�ǫmq�V�+*`�lL�MN�K"j�d��D9�w�I����֣��:��%�i;�����,W��NMN7����J2+2d�'����8W!3�d�M}�/�~�!��͛c�ȗ��6�{f}*o�b$�v��q�x�nd!�~����b�X�7_K��,���}���z���pz����ኵ'�lgӷ������ݵ�U[ZU���ZUV�v��W����QTV�T$�(&�I��U���w��Uڪ�U��U�b��h��CU��*Tѭʁ�k���TւSض��*��QW{����UꪾWj���5 $�{(��J�jI�T��j�!��I&�&��@�&�ڪ���������W��UU��Uy5�ԀH�0���V�T���*��Ҫ��^m�)UV֕UUU4�֪5�sZ��*+jҪ���U���EUW������2�&�T���ѹ�h�IT�j�;9��W��U^*�U��sh��������{�50�H� D�D��UW��U_+�W��8����UW^9�CD�{��k����-�ӧ���� ���*����g���>�g�C�N^|=��c���|�g�|b'��0N����'M��	N	�6t��gN��<!��:'JbP�%(�O+�%�`�ا���*�	1�j"�"�P�e�ڧ�j׶RV��r8!ૃ��XD�r�V�T�dF�
�:�{�e�+%qQ[��6ӑ��E\r�Y��"��4mQr&�4 ��v((J�M&����K�/W3����8�-��bv6�*ڥ�;1��d�2Ț�R)+R&�L��lv���ջ���^1Ȣ�)`hp�J�ב����탽�{�� ���{ڪ����b!��{�� ����`���{������{� qh��4/?��]����W,��
	ٕ��:�D�t�K.b���\a�%%O�O����a�'ŝr��G<	8`I�vf��7$�UBJ�j��m>�wW��0`���EY&�1ˢ���x��NN�w�TyUQ��{�4�󗳬!n,�f�x�Mf�&�L�h�C.g����j4II�)I�W]dΛ�$
<���Y���x�z��(���B��f�����L�M;u,�y4��/U*�k�����u�G�� n���䚯����Z�;�6|��SN������L޾D[UFu17�u���rI!�!��1f2D7F|���-QER�^���h�T�ra3IӞ���՚�d"m�L���L�,�`�֙y�i�3-8f�������J��*�S�㶓��_?�x�ƈ8�%U���J�����ã,�`���9��yA*�mɍ&��B�eö���;{�ŸamqƜ�0��e�`0�z��0b�UB��:�u�F1�pc��H��MVI�գ[\-���)L��H⑯7��*ם��ۜKVs��UHB���di��>��{7��K��,�8t�FCCē-z�q��:L�1��#�6u2��G���J�X�x�$����e3�1�HkG��ek�w/eӻ6c�f��������a�+LV���i��i�˥�f(�^&I�`�&����+f��5���m�<�L��v4�4�K�,it��e�4��Xl�.�4���َ�1��q��׹�ý�7E���z�Un�"�>�od�sg/Z������{�E6�l���1��=��m�����MkZƵHQF�d�� y"?��]1�����HV=x�T�/��!A�BbIkԍ��� �k�X'R�,h>hM�ӣ���`�Mb^�\)��ނ��LDn(�*��ďO�B��"G�'vSM4'�1��_�� �a�Mm��a>ʰUz�k�P�5r�i�x�qƊ�ci�B
�j&TX7&��m���d$m���T�jY�D��T]��&_�X9��:H�c�Ĩ��Å&�[m�8߾Q:�w�iv�(���9��K�]I$2��/"��h�GC��)L�C���4D
b�>��ޜ�l�I�Fq1x�.\�Q�0��`�K�/X|��C��3$���� � !�NwT2�iÇf�71����LxE�R��v���e:s>$�C����c�9�M�Ԡ��JiB�j��A+�~bb��6@t�J^:h"E�8t�a�$�@by����LV�e��x��L11-��-��`?�)m�1�N
�I0N�2D�e�)x�Z�/?����M�J-ݣyr1Ɠ��c㵽�%MC%N�Ҩh����I ���Ǟ�K>_���bx��GXd%�bZA^M�3�k�b�Ì�m���A�qg�b�p�x�����g
81��2͝�"}&�h�������;���,�v$L&_BG��E�z������$�m�9N�%y�l.�()��D8d�A��R��2�9��'��x4�L�&%�3�$\ypK򫋽�$M��Z��������ֱ�4}.�Jpt�,<�y4d0l�A��v���+�uT�Ou~�V *�
�׋����h [˒XlO%.HI$Kl8y�æ%�R�噮��D!�C�{�K��a��w�צ:iߥ�*��>*jx�x�Sǋ�⬘=RY0+K��v].˕��.�3����e�z^�cwL;��K�iu�q˳4�Q�Ȉ����?�M����%���ީ|�ia�&�u��/��&i@��;� �@6�ޱki��څ<�V��o�AM�/cP{C{#jAܧ��X�bF��7$���q�ڢq�*����6�9�P3v+٪��M����E�c�Vi�U�M� M��7GQT��q>ϒjj+�I�`U�֝�Z�VR�J(�M�$T�m*A����Q�6Ԫ�H��R"'����d�W��+�Z7�^2���}����'ί6�l��m6^m����/6�l�m� m���A��^��Y�5]��[�F1X��,�n�mQ��
��Yo�H�K�in[Ӳ2I�`kJCnL9�T��$�?5Pi�%����`6r}��n�.��|�-4�s���(����D��4�HLI-��훶`5��ä"e�A��vI*���r�Bp������X,�'J,�d���!0XO����rzI&CM�{����5V�lRep�;��B;��~Xѥ��Sf��Þd$zg�螺4�S�l��Q��F9���!�/��߿�+REh� څ��q*��>N9Jv@�t�HVM���|�p�rVR�BBL�˒���ŝ,�ķ8phhLg��e��8�Y	c����l8=�`J��`4��+eMٷY U����~^��V�R�c��hm�Y`sO��p���Kُ�L������qY���Q�ɾ_�뺩]6Q�9~2���o��a'�r�;�ԋ˂j�vK�EJzc�ͅ�iF\�a�I)�צ�>,�A��[@��C���Vɓ��!�����*����T�`��&���ON�"`=��&��`�K��j�J�dh�1S5u�||Μ�s��3[>2Y��48�������ے`:��U5=$��h"|��Ā`��%0���l^�����0�A��m��}^-Qz�k�jvu��kႾ(�����M6�6�T[�j+�+2�2��8�m44d�쀉,R��bJ�ɦK9�h��k�e��e}��|dp�`����!��Rc�|��8�&����"o�4T��E�0Y�OcS�� �/�|Y�)�P�j��1���=�!�Y��YJ�*wH�2a(�=CQ���Vr�݅]���.����.�r΋�,6i���+Li�]4��(�<d��d���Ѣ�!�J5Seiwp�.Ιt��.�a�Lt��b�/}Q����x�����D/��Q��R�YTO�{sP$��D* j���b�3Hf���\FF��xh�1���Nw�>
�����w�=�{�m�؍����a��m��xC2��؉��q��̙���-_��ɲ�����uZ�b�aY��6��ê	�݆N�4`����+�;�#��90`/�p��ݮ"���VĞ.g3ܩp�SJ6�j7Ġ�2hɤ�l�^�!�6��z����:Q��d�N�uUw-��k�5��S����(�֚�k��E"nx�ɛ&�ܲ5�	�RjYYt{\�2H�n���^}�\�����5/�v�l8d͇Ŵ8��	&�i����\J.���W��>��-���NƷ�zfiX��C�t�ssr��}D�f�)�A�7�����چf>��$���*X��Ɩv^('��}��"m4:��ի�oǞ�̑Eo�*�(����7�6���rdd�5$q�A�n!��㍋q�+�:҈S>"���~��J4��s�F��.y�q����]�:�2L��<p�!��m�o4yÔ�x��*�D�y	��Z�"L�^��ՊYP�]Z�{�D��N%}�!���ai��<���Ol�h�A���a\�����'��W%5(�i!��MS�<�|�I����Ο�p����m���&�-QT�-G~��.F*�rY�l�`���$#zP^,&Ὑ1�%�����(�5"B4�����|�7�;dݷx���UYHӧ�B�vC��8�o�RUVA��D�nS�8��N9(�����h�M|I4�0��!m�>'g���x���g͘6�.|e��d2;ɹ5(К5�pGfɡ��-[es��PT�i2y7Kf�ts�<�HFI�����Ĥ�L�d2(��t�Kw���$�2d�,���rن&�Mw�#2Nr`���L�&O�1�ud�	D�m�G���6tΗM9gMb��;4a��1ZcLb��;4�e٦6i�+f�i�+�
ẜ+�ɲ�|W�l���x�G��<^��Ӧ4��9���e�3�f�-�ҳ�F|�Ub>\_�K�=�A���pE���!J-5k�N�����j{SNH�%�ݪ�YR[D�lI��m�hp��$.��M���Q��r5h�Lw譢�|wK�d8�+���i��lV����Ԥ�U[Te�j��l����V�TH���N�D�-U_f���!��+���GZv-�cȵEc)j�$T����ؙ�C��~���{��m��m��m��m��mq�mq�m|!0b�j�v(�u{�s.�e���e%MC6�x�HTl��E,1��_+ap��!*T	�'��M�-��dɓ�.��u��U)��o�rTűs��W�@�*����sV������V+E7v]I!��;]�M6Y��d�bp���!����pK393;�4��?H�~<�2<�*:�Р�9�^/~�Չ��mJ�!|���S���U^N�&p�ŝ�O���D�l��!!��DM��I+�< �k��lm��jd�5�����3a>	6�M����I3V'���p]k����͇����y�k��0��up�ri�~�L�<D֊,�vaӗ�������l����}�2z��*+�� >%B�ڞ�I�J�d�$*J��|��A��]��ψ�l�撖�)2��C^�a�Eݐ�L�o$,�ϡ!
(���x�)lѢ̆�!�bo���'���}E��n�((����nM9"e�p��>a�2��tp��f�!��NUI��]�ؚL|�d!�����u0y�9(�;
�	P��J��h��o�|G��{h͕r�p�S11tJ*k�t��E_��s��\�^�����f�!����|QDɃm4���c��m@�V��A�����<y�iJ'i2CK�2SfM�m���Q���>:YgCa��V��1'&=���Tc����q;X����H���e��Lx�SZ�i��D�h�ĥ�ub�.�7"ug�_�E�a%84|���!���`��q�.�LB's&�ɸc��U4i>Jr[�$��?e�:`�f�!�D���ې��%#��8�&S�q7��~�>�䢡�����E�d�0W$��w]N�u�䬮�a{��vg���vcM9gM1���ugJ�1ZcK�]�٬[���4Ɨei�.�u�/X�xvc���/gL�wcK�Ҵ鎗�Ӧ4��wg��^��չbir�\�k6��c^�/�:>�&�|�x�dsg�P���|�}�m��m��m��m��m��m���0�����%��礝m��߃&
�D�3�I�4`�cI����]��ӆ���,����Ӆ��Nh�`K:V�l'|k�v2��LT�a-��iԇ5G�~>z�4q"|e͟uE�,�f"�~~9y�B��nd7ZT.4F�����bm�R���X�� ϒԇ5�O�M�=������m��O%�o���8�2�C}ʕ$��I�CF^Cg������'lKw��	=g���ʱE���p�Z�ƚe1F.�B�(�^�]<��oh��r%��Kt�x��7��4�1��4>��D����N�'4я\��%]�x�2Rcr%|GXB͛�2D�Б�W[h�֘xl�f�a�z$H�&�,�*�hӃ&t�-8>ӂ�O�ه	�nH[CO&���2�E]���(���c��SJ���I`7�D�)��pҺ�]�b��6��4e�ҍx�܆����|�6}�	ig�M._%�;�GSΒ�br�Ǯ�9�Utb��-�<|h�h0c\�!�x*�,����ɓ�rx�2`���dObnlJ�W���e<��9�i2��ӏR�]�nM��k��&�Y��`�]̉�E<�FӉ��M��4\��.]�	�؜l�O�L�v�r�w����kͧL�du��h�A������s����vK���J�O�q����O�I��&�����~MP<*9cr����p��i�W��ӳY�cN�3��^չ�0�X�p��b��f�٦4�.���ٍײ�9c���/+ӳ�];���t�.�N�Ӧ4��u�����:e�K�ir�.X��L�z;�cֈ@�l�Jz%�|B��UiSP�� ��h�~�羞��Y4e
6
���ЍI,ȇ�5c�LCjȒ��>�R�,r4��Z�Aa]#��� T�Z��!S�DHJ�����Ӆ��8���{9K�%Mi�vJ�@�\��C��W2��:6�eyC1����2��q�'��;�;5T����NV<j�E�QR6V�c���i�j{~��{��m��mv���m��m��m�!0�P ��I%�mvYBQB�4
5bj�f:�r[_E5�m�˝�s�.g߳�&�i���Zw�gIZ�c6}
?B��,����$���Z� ��gƃa������N�:֑�C��k�S�7UR���a�m6�4t�p0Y�*� r:|?<xG�tu:S2yx�s�(a���ޟ3t'E��y�|��E�׆L6�9U2�	'd�~Lzx�m=N������tf��P������M�R���k��Fu�U�r�$�q�FЭh#�5d�Sv�!&=f:B7��FƂ	�����Ѧ�E\��%�%U��pq�0p�W[�܅Qv�}ǖI�ͺs����m��fn�⪌ԕd��N�a���2t:)Jhҙ)�N]��O�s��F�_��8�CMzUI%U��2��;M�M6�����RVx�(K<p��`�`|�_a"�6cɇ=L�u'���⤁��#˳�Sn���}��6�	���#�ZT�u�ae���X�I��N�@���;#VBA��ɠ��G)MF����AchC���7b[�lDӢW(cݓ��h�t峇��:h6u=���?4����1X(bEMfA.	�I�Ab�+K
�� V0K2�����ú=��p�L�`�QڔY��)>0���ap�Kzф����RT�F�C�x����Y��SpbK�K1�@lv�6VՑG�U�Ty[iAA�e��UV$Ӱ�\I=Z֐li6�LO�D�3Ǟ�}�t&�&�����i2���,��B��d�s���/�)�~~tx�d4�8h�a��v����4p���G�1ڝ ۭ9r��n��R]�vQTQ*�0��YrZdѦ�8v7���!ex&��b��q���4��:]4�<.Z1��1ZrΗK�f6k�4ǌ��`�#�&��6b���>&��8|�.���1��t�]+K�Ӧt��c�,r�6a�,:\��+�r�FQʚ%�i���U]Qg��c՚�%D1
��LS����� �7Z����GQ
�!ٸL���Qbu�d$S�y�ۃL���W��m������m��m��m��kZ֝h�d,�'� e�������z�w�.��J�3E�5ə*Q͹9�0�HO��4d4��TźB͇$�x�ʕRB���m:H������K%|��Kє���,�}����g��B��%W6V �U,J�c�M����cpqK^G��F(8�����q�:H]c��dx�ؤ�ƻ'��%�S�Bi) ����Υm��=rFe�=-��C��=��W��3ך6x��Yi���M�NstT��$7��
Smږ�PcUD,������#�rB�T.�c��}�%i-/m��h�h,ͦl��L�4ϙ6GQ7��'���I#$L? `y��U�=}���Ē%�O�|��Æ�gO�^���g�6x����W����ה�H��In�Xf���O«\�rr����t��e������YK�[%Z'�`� iAY����r��̓JLݍHB4I�������/q��ht�"i0��B��}A$�!	��M$~0t���Y�ݬ�f��#���`�>��_�~���Q~����$�������xl�f��iLzd�wq6���v����Ք���5���%úL;u�o���6s��l�·Bϳ*�ö��&�bW�����/������<`�.|���(ӡ��ܻ7	'Ւ�J'&�2b�u��,��-��٦t�i�x\�cHɟ!���STM_�oQW���?���gl�.��wi������c�����1���]�c��t垹^soL��eIe|K>�eO�㙛x[P�$��a$r��4!R�H�٪��b�ť�ȱ���qJ!� �L"�Z�x�0RF���D� �b�@�Yl�w��E�$K���
��"�e4���!��SF_a+�@N3ϫ�Կ��đ��������w�f��)�Sh脟-d�8I��NG1������J���&���vN��f]o�Q�Q'Qm���X�FH�҉�!@Bi ����ӭ5�'��c?f��>wݶ�m��m��m��m��m��m�a@�1�x��.D�"�)��MZY"���c�[!l�+[���:І#XM"."���������E���~6�K2�G$p�N5���*(�$~�=;��S��65���7*J��Wr��ec�N=>#�i�gO�ۆ�ڪ*���Ӯ��$Ө}5OY���/�ӮO�����'�||�;��._�>|������w�e���k�4^����RT�I�Q�S\-/��=��\@�)��o��˱�h�ば�� GVϟ H���b�6��EDf7i�E����]jiZc,�y�$�F�;
�?'����G�p�<f�pe��g��wؼz�,������w��]|�N:,��<���vg��\�]�%����	)ˬ褉�b��h����M��^w�fw�/�:`�p,�`���4�zw�j�稥�U�B>]O7:�����6��mEqAb$�1���<R�K5����G)9�e:`4r���Σ;ܹ�}�. �`jI��}y�BKyC��Ӱ��h�ޕTe��h�����U5⿻G�P���6*��cM�ۣ$ɴ�d#5���IF�c��gq|��}q�qD�L��2y"srBu��+n���d��Oi铅�fHM8i���J��:���㶛垓�{y!��@���B{�VQ�Gɽ1�	!��7���h�Uݧ,4Ӈwwgv��]۩ ����b'؛:l���ۻ�i�f�wiݦ�wwwr��wq�a�1�!�!�!� G��I�\=��Ȩ�N,�泼���;�^ep�9~m��m��m��m��m�m��m�qqER��7���s��T@3p�a!�HI$�m���=kIi�ٓ���a��rHJ����0a�<|B@�q�f�Q	,�i��Iþ8�:pѓ���no��Ď�r�]ZnMjBD�(�vK�$r2�Z�@g��^���ڲ܁6h�O��+I�?rJ>mݖ�$.���?%]`̨B?��w�fq��Rc)���^�WU�#m�B�*�R2��m�q�a3�J�UwM�ѣ��%&�9U�*���FN
6�_]?$��i���1�͗/WNY(Xw"�/�b��|W;�1y��ۋm�$ˇ�0h�f�<G���uwd�q5�II�Q��tۈC�S�6{�<���A~��l6�����8>��%;1-����g� �"�ne��j���M|�g����q�Ӄ.N�MS=������1��.o�x�����	Ƭ��<r���ř����0�i~N&:�Ǝq�,��\!U|:e��̖`0q�O�0�M�Q��w�O[ϱ���K�NO�%�Lh�1��CU䣩��L��',�`޺���u+�%BQWLN�4e�$��޿Y�掜&Ki!�e�ky�t������D���n�jW�T��-[m���*bHep����;?�}�4���������*���ٙ�H3DI��&�,l�|i���-����%A	$D�IH[�`�H�Nl�d��)RRĥ�,)IK
f�	J��)RRȥJXR���)1���JE,�*E)����&�B�B�B��
Y
T)d)d)�LBR�JJY%)%*%,���S�fC%,��JQ)Q)d�Y�R��&$R�*JX���
T)d)bR�S
LI)dRĥ�R�����JT��LRa)T�J��)R�1(5@���c��ٲ�F�j[-[-���1X��Ib�b��8Pġe%�v�*ZUQT�������)1)T,�e3��J��`�I��eKJ����L�%RҨ�EX�I�U%�*��E-ZUZ����f(�-*�U�T1J��R�iT�H��
F��Ie�*�R��I,���U�T�P����*YP���,T,Qb��%U�e*�UR�O��ڶ[mw�¤�T����U�UeUUX�b�eT��b�X�YR�,�YRʖP���K*�K*�*X�b�J�����VT�K,Qe�U�,�eW8bQeB�-R-KRЪ��U��``�)eK)T,��,T��e,T��(YVT�RʱIaE���IRRP��),�KIR)*%%H���m�Q,RJT��J�R�)dRȥE1�	�R��JXR�����L�&"�lclCRĥ�)B�
T)d�T)P�Hs�Q��I����Q���	2��慡4О�X��q/��"��H��B	j�x�i<1��7����o�߷�������#y��~�3�wfLz�����=/�����uW��;:ls�i���\�o"���=>>��;<X�x���>��'�M�L0���[�_��>1���F�1�=�����s���`��!	����9>���������yI�Z$�E:G��X�HY�bU,����?:Oj}�v8|>�~��6=��GL9#؋�<���u��'��_��Q�������K�%�9�����D~'/�$�y?V[g����?�T���,6;ܲ;6M���C`�G���$�D�'�%���?{�bRR�l�md7�h�y�۳~dWoFX�O\y��_k|ɼm[���ߦ��������0�rP~ϱ�ES�s�𨶈l"�(a�B� ���! b*�
��(4@#D��b�	7�ݎ6Z�d�`��Yɉ�i��;��ɺ8O�����M��K�)8Q"b�D��RҨIiUH�$"�!)e	r�>��~6_�=��T�F���z�������O�sZ8Nʖ?5�̵7��'�nfG���f��Ac��Ɇq���O�S�)f �����Y��0��>�r;O����3�O,�̎��������S=���?6�����_��·�0��E��+�ꏄO��ϞG�9�ξ7�����O|H$<Oi��"��x'��q����}g�oN�N����}��0őU�^���$*�{�A!�I�O�"�=��=�t���.s#�ɺ:n�&O$�I�w	G����%�@��?�����.�)S��ۉ�|�$�	F�S$�B�g�n}=ǥ8$�#��d�d�ɜT�#	a��a¿�����%�ژ�NЋdn�͠��2��*��#c�?��$0F�OS�W�>-�����ěp�ĂC�6����U$�Q��'���o�`����O��~���1�{��=o�����7L�"=^����K�O��0=)�?��|���1`l�~(�>籄�s��i��������	I�3g��OI0�%�R���T�������H`=͍��^r���S��sڏ����A�G�O24q�tyr�1e��	eW���ޛ�UR�n��͝2���y'�la�S��D7�=�?��n�(��E&F����9𜣆�;�wr��m�#t�_�������ĂC󿵉�'��~�cp����B=	�bL��1�,I�N�
�_Y��GoqM&��'�����{4�	����O����j$�C�;Ǧ=�B�"M�Rg�O�6�wu�"=�g��9����$I�>���I�N�w�p������ۣ�X}<��~�Ϟ-��F	�RW�X���z:����]��BB�J� 