BZh91AY&SYNW�G��ߔ`q���"� ����  b!                                           y��P  @H P    �
 (          
          s�B(�P��H���d�T�D���
PB����P 	�E%T���"IUJ))	UDI#��BR)wP�T�
�!4P��ї��R�n�r�-��c��QH����H�.`4@4W������ê��q ��@ P��*���������R��,2ם�m��٭O���G�G�����y���ݫme��hy�ڠ���m�y���������`� ����c޳�
 *����6�t�EB�*���JT�("B��Gǰ��������� �}�T�}� n���ް{��}>Z=� >��J� 	`i�P P t��)�+�|� }t\�ǾzI��;�y�@� 9}8���^ �zu�9 �`|@}�  �R�  �}�(;U���ET�%
�'MR)x ��9
� �{ �*�ޒR^ �zz �@ �� o�T!�l<�>�� P��� ��)����� �㪨� &�@=��=��d 4�(��� @�@���( +>�R(���D��QDTE ��I| gc���ru�� �΁T����` m�{<���*\��b�`p ���}*!T�p|�>�#u�t�w��E�l<�=�� $ X z�IJ $ rh�;����    �BB���H�*�
��*J�| l��s�;�Cv s� ���@4��{�P�� lǠ�P � �� ���w0 MT�� -� @�@�� q�I"�R �`�0F{ >     S��T�Ta4`& LF�`�&"���)*� �   @OF�Q�EDm #&��� i�T��IC ��@CA�d	OD�����  1CM 	RdM�m&L��=LF'�ɚi��}W�}f~����::�ɉ;�ߓx���q�"�"��ݿ:��+ʢ 
�DTDW�%q���"����s���?��?�=��*"+?�U_�� Q����� �"������� �AP�����T� H���1�b @�H�D1  �@ Ā!�EC�& C� \J8�qB��q�QĀb@1�q �J H�Āb@1 �q*�Uī�P�+�G�$��W� !�@�bT1*��LH� C& �B )�W�$\@��q��� C�%\B$C��@Ĉ���$C�� � bD1,H$\@��ĉ��*�1 �q�EĀbV LJ$	� Ĉb1
8�C#� B%J��q 
bPD�
��ER%1*�@q *bT� ��C(�% L@
��Ċ�J�'����l�����p��o�?ȖB7u����Ԟ��/�#�k	����	פ�78��4-�4a}�Y=�����ݸojҎ���w�q>C������c�޷�䑛�O����b�߷(��׼0����=����r-q�x�;�"�ӳQ[��\nn�z��(����C
7vML�x��\)gjʎ�nv��{Op!h���wE�7�mz�iw� X�Ƃ�X	�9��1�.���v�����0��y�\��F,B��}�OX@�(C�p\�f�Yܐ~�x���v��ʇ?�2<�߆�;��y$���`]LM� �rv�>%�fk	{V�7$���ԡ��W�Z������1,�s���V�_�;���`iJ�wҁڝ;��L�ҷ%,���w�{�<p�7��v��}4S�H"�)i0ntuS��7��Z�J5C��KoR���&�Bc����9.m)�)�aV�k|�`y�2�W�Ge�9�J��u�E����C{�m�c]i�[c]��D�+i鷴��A��Oa��2qN�3J5����G�xȤ�էy�9앻�H��y��;������N��W_�j�O3s�]	��ٸomڕ[H��tA�[J�s�q0C����!u��k ����X�y�!���83fql��jD��0�i|�/y���cN3���#}�<���8�&�]dqV9F5s
�wP.e�u�k#��#.m�ɸ��#�W���y��Q��Ҷ�(��y��B�T�9�����#˕��&��oQ�7坚&j�����L��%?l�s�B��p�4
��wv27�����P횆�.|�'$�o�l��&μ��R�vkeٰ3���"������;f7�k�(=��7������U�B+�g������n��u@��_axyeМ{��$fh�5���2˓����6�k(H�9��|虩Q��2����4�h!�CI�|!�:u�,��5���0q�}�TYכГ���("+���UP�F�M�T����
�ʆ�0�N䝉=�PV��:�M=�d��y:�Kxom�����{�9���ص�l�zN���}8pT�r�1E�&�,�j����j%bY�ǯ�Y������T�����ϣ�H��cɐ�Zz��C�b��@ͪ!��Ķvh�@��7�����S�"Ň�:�QY���M3��ٳ��Y���"�Ó;׊�vE�9�e�$�gp�fK��r�v\x˔u�@�Vw���w���䵂[��r�^(E��v�C�d`���i��5�j<Jp��^�,NG��44�Z_R:$��u��H�X9hY���MX�\U�.���)�����;p�#���d	�,2����M;F,�A�׺z�OqƤ�`��d�t!V��E����s�[�w_q�#�JD60��N��\����^E�ȾW�B�+���:~�pǺ�o�v��ہ�;r��b�8��*d�6��1���LK+]s÷��/ y�-����tɛ8\�n�{GޭN�0����
q9I�|Ï���ҍ��(�X땼11��޳׶�r���2p������7��r���]szU<؜]S:�xf�Ŝ�7�[��Ԃ���,{a���9�Y�Y�O�f�g\=]��;edpKn�8]c`�r��2�{q�:�܎r5�wp=VG��%� 5���Nnm͑��ɄF�6�*�Y[�:��Nh|;�U�J:YY&��L�{�x63u���i�jr���#ҬF=/v��-23`yK�ݵ��V)h:�Vj앳��l;i�Q|M��ۛt;o)kh�k��ڶ|	�,/lɑC�^�*vv�!��,���]���B`�&��Gj�+�f��kw��Dl�n�ק^�l��ٿg�	��㳇�-)�WY�utwZ�n�F��]�T��F���Ɖ�WϦ��Nnu�;[ñ�E��4�#��(>?�2���!��Ns�e�����<����V�-X~�OSfMb�Q�L�J�٭��.��{��}w)s���i�Y��F���븞��r=��]�n�k����˯�>�%�w|,Ǥ=�.2�����=X�lB+4I��9�b���ge�vKי�<�3�h*pzrg5�h��{�W]�kÝ۫�v$��]Q���f�&��,��sz2<�������~+m� ��9��_
r�u�P��ϱ��r_MZ�p�Q增o;Z�$݌%��s������"��3z)�ΡM'��C�a��IͽČSZ�xkU0h�G�8m�<��L�&���[��*�3J���$�u<��Ή�x{ۇ`c
�(��7m83^�`}Z�od�/LV-�r�H�|��޸3�(�\O�����;��N���钭�ɰ)�{r�%�`�\�Çe�g[�h;v���ԭ|��`��
އ>��j^*��;5����D��.[�w+њBeˆh�3u׋�^mz�P�42W�P�64GwL���b�!�$0�Ŗ�|"��F�eƵ��g.�V���Wm���lM��e� ��Q�	���c �*:w2��7򝩳
(�g`�3Hni����pa��rv��F.v��.�{�v�в#��&�M�u��V�;f�3uC�ˑ�`���5�x3��{�>��?�T�����'�X,-�h)+����Vfo3Þ
t�P@�`�ܫݟ>�!o}f)D#+�N=#Y.�{2��r5g������x�L�HH�l�pA����-�؅(��.QfD���	���cS�vn�cm��t%�G'0�R���):�:�����������&�LA���~�I�I�	��Ǜ�p���8K�[Gr?mt���S��-�U�����8ȅ&旲՛2f��&�ߪ
s��ԗ=w�[\a��;S�N쌨���c_j�ٸ��8j����
E�a�+}��Q3[�ˣ
Z`]�[X�?\�"���u��>��Ź��F�\�g�i�o�]�5���F�t]��cj��J���:�9-k��{���-�ӯ�,�f=u��n���j�:�t�}�"$K����`8�s%`�:��v�Z��Qż����R<������@�H��kqoR�,夤�=ns'@n�z����Z�O���W\O"��3����ռ�m���.0�a !��Hn-��\������ �t�f�;��\¨��UQs����>�|�Px��cMDy���Ţv��fj&>�2=\��@1���� [z�!b��g>r���;P�H�G۸A
�&�Ʋ5���]��ˎEk�5^�kɰwu�x��I�����n�(�׸7^��4VE7�Z�Wt*�&u�3\X�o�\9n�����ϴ�wC��#�ws�!oz�K!^�ܚ��C����P�+��۹�@�E��b��9�Uŵ�
e�ִq�kWq��k�&˴f�8��Gi9���������1=&c0�����Hӝ�Ngy]��X�:���Բ��#�p�rjA���F�nռ���Z:�gP��/���#h�77/���5!�Q� Y����hq�ln�\l�@�>`ϏrXL�M��LJ�
`�(���#F�vt��[U�"�9h��4�E\�Eq|�C)����p��	��ٝT��8ssdpMǢ�L�X솦Z�7�r �]�w�=���CPC�,x���w�|�$�S�E≙�L/�۪r�
Ƭ=��G*���۹r�l�!�B�ޙ�v]�ຸ2� ��$����3�#�����.s���v@���r|8$p�Ѕ��*�L�5�tR7�qm�\T��7ge���[v��9c5�O4ָ�������ѷ����vd&� �O�e��p
xMRw�X���c5����sNڟv;�d�(�4n2��pv ��]���b�ƎqM&Gz�V\7��qÜ��Y1��s�v]<ü�.MB��2���(
]Oc�\E����H-�8��Ś��Y�s�as*ʺ2��AM˓�p�`w�_.{���G���K��mTqK�l�&'�.af��;�!9�7����z{:.*p͖�T�.CP�M�����bZΡ�e��j�s��;�+�G��	��a�
7���ݺ�j\;Mz�A�wv=f����f	2�Q4��û���z6n�{,TF��k�vk��)��.��Ǹ���7�߁st5Щ��#�@t%)C0��k靼og5��^<A|��A�r[�m��0����Ò�1�=���`�:Uk+��u%��8�7�;��~l`w�C���򾁩C�3����MY=��w�ᬸ��qo&��i಻ӵk����5T)�؉�U`=�N�K����h���^���&�*�ղ�Y�P#�q�K�ᄡH�0-@���ݯ��a��sd�7)d�ټyHα<�%����ˈ|o'̼�6>���S
Â�®�����q�c�����������wۓ`}��h�N�����C���f�l'�3-��H�B*�Í�D�
)��b�uH�oq!��7d�k���r�H��89�)ס7�ӗ�^8��u{&�d��R�<6ر�B-Pjk0�1��lL����qT,�8���<=����	0A�����ԑ�op�5^h��c�o1v!Ӏ4��y�n�Մ�'0�}>q���rdh�D'[4���g	�;:N�f�YAZ�P�_wi{�Ǖ��������cq��vns��ay3�"rү}:��Ä��رf�-��`}j6���x��� ݝY�wA*%�ЦU�q���<���h��xy���t���'��'r��Ţ�M�<�3�67��qE���.ot�9zf�j2�s�a}�Z-���۹O<���쥷EkؔM�wd{;;�j��
;�ağ}�+�f�Ny[��Χ�`�n����6�T^XSxUD�ٖ�m���^��3>���U�j"m��]�)�em^_����TB��.�/�m�����p�?�pZ)����3��Gn��ܛt�����nk�z)F��9vޗfX��r�z���{Of�'S��޼܌�{ 6�ݯ,3ˏ]:��h������͂�,�<Ӫ�G&�dk<��swb��[�n���)��0v��gq���oRb���)5�����u<���i���E�0����E*hǓ`��P��H�I�� a��ڻ��q�� Ï���s���0���n2�zf��j�+ܓ罆�f�؂=Gv��8�0���0�zϫ�`*A҆�������϶�˷�V�]��5歘��z�˓��K��%��U#���b��i���ܽ;�WoU�9��p��Q,*�}0�^���T��H����"���o<B�|������'eP㳫ďt�yc����u�S;;����4�,���,ٜ5މ�ÿ�����(ry�<�����e:k�2�t�jI]�;�b
�����q�{}^i���;��s�4H�"��.�V�D��f�6p����X���s�O!.�8ƽz]��>{������%�p�΋�͇#�z!:�Iå��])��]��LP��"c-�UK�X���2%�]�����%�y�M��u.�/�N���N{6�����	7#�Q��'�<yu��]�+�I�W&��{t
�s��m}�R��{xdc��	v��p���m�$�8�/'4^�$�N}�=/�g窊���A�&���3�T�G>CIYχ)��X7d=���
�˵��+lj����.��X�]/{9UsDWrf����Y���
m�ǱYݯOt�ra�z��,=K���凉7l-��S�6�9M�gG׻�Rs���˖��(�Y��<o&��^���݀�ʇE��q�
��p.�r*e�>���"Z#z�v�!��jZ>9z���o1�`ݑ؂R�58�ݛw7g.W1r�I�D�edp�a.0��R��yRn�9. ��u��柆�8��#G>�c��!1���7p�J�xw�鸱cH��MF��c���D&�YZ�2���v!w%����>���tK���*�×��M�&�;u��������\����f���ؾ�#!J��������`O��K�@���oj�G�k���Wj���)͝�wp���l�؈0�6��^Y���7�ܦN��O����(ǲ\�p�fvf�vf��%ȴWoϰoo#ػ��;(�>�=ݍ==�t�2i�x�A��8|@�j���'}݇yn�0�Ӛ�� i�t�x��<K+姺���� D�|�����弙�Ѹ���vڛ���Wr���4[��ݗ��fٻ�!�$e��E�$%c.���ʬ#Vu%�k�y_��{�Ⱦ�;q��1�La ���O6�I"�h�������a��.������]�Gd�Y˷!7b	u�k[gH��W[�1(��'p�snƜأN���>l�K�W*�#��,`��Y�2�H��\g+�R}����ˈ��A}�WV�2�W5���x�a-HNwt��!.|u��7N��h<G.��gv\x ��-�*j�6�9ߞ�m��P�{l��u�Ė�ȧy�����ȘYÿmnze�&3��9���n?�M��q=�q A�Ï�{�pg-�{]W�i<#hc�w�W�s��zp��5�}.q�C��!9d^7��OY��8b��?����M^��n�����w���>;���u��1��i)Q
A��E(!J�P
:E@ h*�!�@t�R��R�H��@ Ђh
A�H�@
P�H���H�B �*�4"� 	J (�@�P�J�Pht �iQJ]*4�*�P��S@%�P�("�B � �H-(� :�	B�ЈiTM(��
4��" �H�R �UЈU]*	B�4����-
�@H�"%
Ѐ�4P"h) �@4����!H�R 4�� 4 R
� - �M"@~b���Л�;x�iB�c]ؾxy
KBP<�x{|��֗���Y�Z�i�Q[�zβN��Z�t5������w|�o����R�[�h�"?���.�����/�����<o�-�n-�~;v�c��U_��Ϸ�UW�׿^y���ʀ +���?�����GϷ���ϳ���.(O�.&��� �!��ٻ���&)09_^#���M}�������ͨ��Ӂ�$\ ͏XL��{����|;���
g������,��4ï�C���^��O^Eú�_�SY3�VIk�*�����o,�R����?�^eG�L��d�;�o`!��s�tk4�||u�aM���H�v%M��{ɮWR�F������wa��;�g��j;h���S�g��j�0�����B�6�;��S�o`����e�2�%�A�ݣ�V��6\�gL�{���/���F�ޝ��O�"{�mÄ��e;��aKs�,�ǧ'�[���Oύ~�b��K�.��D�F�Wؽ^i��3'rv�-��w�����i�_٦?���=C�,�w��7�t)c��<	�y���f��q11（�vj:7������.��	{à`��=�'��^=���Ё��Wt����oQ3��=fW��*ս��'hB����\�P�6�����=׷�HAt����7o{}f�=nzs������!>�y;/z⥎�Wl�}M�Qe�C��WC堬��������O��g�NξY�S���G�O"�	o�㜈��twf�>P���P`xbZn�G��93���� �p4�ӻ�̔�X�<D��_��^1���]$0HJ���V�7���O����͍�,pܘ�b�	X��	0`���0`��(`��0`��F0X�A0`�� @�� `��q����z�[�l�?nM{�ѧ#�O�m����I�l0x<�Xc�E��ד&t��Ԧ�pY~���}���[��G�b��׻(����%��4�7Lޱ'H.OJ)��zyI��Onϐ^���j�I�&M��{k��� ��	t/(����X�p[����l"-D��Î�;	U��EǮ�+()�z�e#8�H���"nDa2���c��g;`��7h�OO�z�n�-<y�Ռ��W4�O-��&2E�(:犗���e���q�K�H���-�/=�M�,�:W����f��\���8t=�^.7�{"���1��>b���ث>X�Sx��tfۛ�:hל,������Do�s�g`�pS:ύ�������{[:�j��>����O����;�/n��}�����O5 �F�vnL;���پ��{���������H\5���ɕ��Kp��8�ŏ���~l跧d��+}�w��FFf�R9M����Ͻ����ٯ�����)sdV!��}�X�F�;��{�sd�̯Ӎ��v+K;��W<qԥ�gt�}������B��cʟ�S�<���}��ˀ�T�޷���=�x}�C^�N��37L}�|`��s}�x��X�v�uk7�.N]����؉$i���Qo�c��Ϧ�T�~���'�����|��5^!��08��9�$�C;�B���O��?{���
3O{X3��������Z�,<��M��io~}�D`����g�F+��g�Y���G���i��:g��<sBO����i=;�u�B7����{}������kϞ�K�q�����'��s�O3Ol���Hy�]�o������g����~����;pr�:�Ǒ�w:Q���.�76��b�/op}�IR@����V���/��Y�<����BH�,��P���~� �l��:�����"�㒞X�5FD���+����_
� ��^���U��ѣ)}����9Ly.�S1�i�ގw�����-��V��x\��>K��T�?w?v��e�w��j�|x�Y��M�Y���a��O7|M��s����Y�e�Ç�ﲘT8!�Γ�.m|=�v�-Q��5{��!��5�f�E�,dԽ��.����>���F8;�^Mf��w���:f�⾓��%���O*�3{:s=���4�q��:)��g�<�����ovy�KL�J�D�M�(���X 0y�e[��u>���Y��{��������2ګ��=�ц�^�.�{����{�q�ׇ���l�-vT����F�7�ym#8�݄�s�w�������'�޹Nzb�/�HQ��V�3�T���J�e�]H�V��nzXO{c�w��x�G��<<�f����-�"m4OO��aY7~Í��������#�0`���0`���0`���0`��� @��`��e�~JbVeD��̥ы��y��X^̩*��s�������7�n81�bܛ���MνΫP��4�Y`�]�z�s}��j\|�uڸ�sow����{kL��v	�:��5����y��秦Բ ~=��핰;e��r���t���b�s}�=���|m��W��ծ�y-W�u\7�>��y7]�W �)׷�#��r]p��"�����sxoa�Z*��i^��=���}|�����{���h�����#���k�O�.���zpL
3�Nr�n�������u;� �4]ǏO�n%Z�,�1��\��_{ ����,_.�8�>=*��k��qýV�[;�s���o����{�~�=��4�{�w]�>��.��>��c�_{7B�ٞ��^�z�\��q�+{ �+��<f5�]N��h�2x���N9�����g�li�wS������,�E�<g]������~����@xȘo�<Wvz����A�^�l )�՘�͎�����=�l���dP��� �vܛ�1Q~�8W��m�`��*�F{f��@��%����;q���4^,�+������ǂ�P^�L�:=���7w+�gnw#껱�y�2����3gb@�?$���^����_`I��g�'��{Gj:�a����:�D�׶{��+��d�w�>A��������wW[�uS�vo���H�����<F<K�h�<'�iBF~w/c�]��^�Pk�5q�֦u|΄`�{M`-����nG�� ��ko��������d��8j(�	,X�Ƭx�>+�G����Qj�8��<��h���{7=.�q���� �yk��7ٲ��yv���T|���07��7���ݻ(� �e�N k]�}�S�2�>��{�x��'\5M�
z�yU�� �+(3�g$w��gw������Jޓ��)�y�)7'H΀�(zº�L�m^P���9mr��<�Z7<��Y����N�����*������,�M;}��>��yO%����sC�',��a��D��������/C��W�ڽ�j�Ǉy�1N��&u�g�C\��tݜ���føBʸ,��C���ַ�B2[��Ȃ�������|;V��ȉ}��^�@��M��R��ٶ�8��܆>��%���s��w���4��ˍ��%��A����z-��}$�����ؑ�к_Oj��e��8{��J�*�^S����Nr#w�f���u�B;?^QC垢���}�.wm�%�6���������(���if��C����8����ܠ7�=n�mu�{��I��a���2��g�ۃ�����6y�����o{w�4���n�Fc4�����wޚ��x���8Q�8^���!?t�ݍw��!=10��8����@g-C��o]�g�����9����7ϸ�w���8�/�����a�^�����#�����H��'bם���r�����$����w���|:y�rZ2�">�~<��ܺ��$�Yd��q�{j�4q�{x�r�M��gQ�=�u�h��"��8�j�=f��f�}�7���꒰g�C6�w-cT�4�R���}#t��<l�9<�|�h�A��n��S��K�x�/5�.�þ�����V�Kˋ>���x�{�����X>ڦ<\Ѻ����U�<��yE����F�xK__L׾�r�ȱ�Y���ǡ�)>NuzVgA��o���udW���jg_�����4���2�˸��n�r!3ٱw�fG�S���=�+ᬙ��.4p���C�G��� N׳۾�^=F�ȸM��y\�כ��9�4��z]K��5�x4��5w���I���a��;<��O�G>�7|��PE�v��Z�.���&��E�����51���¶NW�c��:�~,w�D��ˋ�s�g��XǱ�8�b^$�<��l�-�5o�f����i�މ#��.�^�}���͢r��\������=�l�Fn���ό��.��W�q��^���J����M�ֺ������4r{�����~>�1�9=(��n�o4dW����#�lb�!繾w{���ͺ~c��v?o�#^�%��#�Gk.L>{�{K�9X�yБ�?L��U�B�v����Tx;�G���)�>^����)������4i������{p��;|��]���!/�!�������q�|���k<�m����K��;W��{_W�k�=� bx�*un�s�4t4��{��ξ>�w}�U�_��^ ��x�r��� �[	x*� ���+��4�!�7r�mK=�.xb�s��{_`�{r��b�����'�*�|�@��|3���#;<�W5<���/csY����_�MM������`c����5���^��:���]�|���=��eIwx1C��M���yr��[tgU�<�;=q,�ܫ���ͻ�a[�������p�����Z9	�|�N�Z:�E�}�y�s�����Y�f���4.q��ߺ�,�x���ƙ+^�|�{�;���|!ɞ�.����0HE���:JB�]�<5��씴�˹�����f���V�kE���î�*�,�Q���yc���w4s��ǃ�r�Ӟ�y^Ͷ��}� f���<-�;�Ҳ��i���Κ� ���Qo5}�Ǭ�]c��6k��:��{u���R��еU��p_ ������7%��®M}}���'����G�sSk����{y$�:!�7)^�<�nvI;:,?h��Qa,�'�Õ�����	_p�<��S��6��4�����ch������xz���g��}&ygBm&�HW�*��h�xQzK�Ӿ�~���b�*�ʎW/f�����D��xs��� 4x0���9�<�ޛ�"�����X�Ҿ��37�	4�||0�Y(��ڷoy�{�zM�'gA;���N6@�x�]�⟨�p�}\冯b{��Ӂz(z�� Kڠ��4ՠv{~�XVZ��Hꞯ��ܯ�gc�zm�^�|3�f	�5���${���z[~��O|��[�08���/z�PK3}�k��=�e���x�����g�MV/W��m�٦{x+�f����ْU1w�voܝ�x�
�q���=:7��z����Vі6���2�ó{c� =�v��>���/�f�_���y�HUFh���#'ӗ��B��t�<j����S���[�y���'6�Ό��+�� ��ty-���m��W;]�gg��r��b�����j��;�A<7 ��I�ō>~�U��=��|Y��k��b��	w���Y��ؓ����v�ց8!��QaF���wH��zw?i7��W>WrM�����+5������{�ꖝ���9�F/xy�L�,ދڬL�j9�����h��ȫʡ=8h�:R�pK	�s���;�˂�_�	���n+�hw�	��ٶ������&�S����s}�w�>Κ�m��(ڌ���L�w��{v"���ݓ��|x�xy�u
�\��O�}��vB��pŭ��ww��dqS<S�����]C'Kxg����t��������ۺ}�t�Û�y���te�I�ݒ�}��O�~���~���r��O~գ_�<��}���x�VM�E^<~Jx����B�9U\`.^�/)F�<�I�ÜϼF�/`��)�ZOE��p�ux����f˹{���=�㾋�fZ��s�[�Ǽvu�7��s��5��2đ��[�g1tg�{T�K��އzٛ8�%y��8My��Y�J0`3���Q�0�=gv�`��T&���.���3"xl.i��`�/_t��cއ�g������{8�M��n'F���3��\����/�g�G�z���7����������/p.%Ox�����ָ�'s �^�g�ae}g��P{���m�<�����/{�vM�����_wL&�ك����=�������N?}�}0.]�g~��S�A<�^@�\�ɗ�<8��f��I�0Q����N�$z��Lw'����'�K�߻M���y$G����#��nG���^e����Oy�a�o }�>��}�G���{_�s�"f�e.�G8l��#�E���@�p�v���%�ۭ�{��~�!���7B���I����Z�x�輎.��ڼG��e�g�ڂ�<�@=�(R>�g�|����cc��g�"v�6���r��Rm���k�y@ogQu��A2���83��s�]�|c�9�MZ��'�?w��D���l�j������p=>���bX7���"��V,Rʟ��Õc.-͗�4��6�^�'���}�:T���n�r-D��8��bޙ	jx�:R���8{��ˊ0wW�w�:�����8�>����+��C	$������s�aI_K ܞ)v��!/z��a�G�x."9�c��rT��M�3�g8�����`�v�=m�6��S̜laK����_g�7����;���?q=&�����|n���v����}�-x�n��5t}Ь��hy�ϊ��k�K�����:��{ �^�3�Jm�}jm�w{4����rL��j�0p�g�N����W�LwkKFp���7�)6v�;gm�V{�ue�;��(��|�v�u���gax0�G�+�X�)s��usH����W�tp[���w�PB��g-�_f&����`��=�/co���gmoyG�Mox�F�����J��ۊf��=�.��*k�L)%�ǽw���A��W�����ݍ�]��z�p�:!��P�7���6��p��.�wO`�n�e<�g#��]�c(�+�uپ�������:>�m�˥�t��E�^˜�;�۟=�����Y� ������~O��?����������#'�/��UUUUUUR��2ե��V�e�ٌ�-���7&�M�W��+.�#���.3�9��U�l9M�-&4[�������R�h1x2\ڭ�:aK���`�j*��q(X.Уe�����b�+��:d��ա��ڻ]"(�E�N�KH�[ږ�[�B��(�v�XQ���X��⮨����ĥ�X9{L�顥b����1�(Վ�eB3bʭ�LQɪ4��l�K]+5P���4��	mT+���֎"���ʏ$آj�jA�kդ�f�`Uҷ���,j��Jd�n�`�l@D,�ٱ���Wa�Z�b�]��+�a��lQh�Žr��X��1)�M��Ec��@�W\�."բ���EV�KjR��� GH����vbqjP�&�\�Q���֥�.�M��mHE�d�R6a���[�%�m���kn��Z&,,n��ŔF��4�lk�i6����E(6�f��/6֚V���435�T����Yhc��5-��T�]���1თ�Ń��sf�Hd�wn�8�6�9K��c&�h�]-vC6��`ky����&x���j�d.��bf�i�(�P��Rf�P�in�f��HM�+e���3d+/e�k, ��X���L�ͣe�Ԍ���.+pJ^�6�6��rE���iGi�n���u"R (��4��1a%���U��)aH��n[�e\XLM�p��&�2�
]HW3�FEJV��&�؁@JK��֥���)tK0�lԗ`p�V�e(W5\.5�b����j؁��b.�˭�V\��td ���5����=LD�v��X�e�Fց�Xk�qM��]@�R���-��%�]����)��K����n-¨�;�b5TΘ�ږ��,rFT,�]�Ŵ-U�V"���K�i%6,�,I����Q��jJA��-лWL� ��GMvL&�[s��r	��:�4	6 �5IRt��p�M#�ҽn�RDR�,%��K�]�+� �Ll��i2B�]]H䙃4s	k+�u��Ҧ+�s-3�M!�6j۠ bš.�@�Z͖��@&e��]	���kԖ9SEPq��2
�v%;hD�Ͷt�s\����ee�Қ�An��f�X �G,r�C�J���Y`�͕à�tY�n�;;J]ff��b��Q��Ue�� �L���K��il�Ѝ��v�fІV�v0���y�L:�{m��qE5��Y��B$4��jVc&M��`m�IH��1�]�jsS1Ѽ��9ríڪ�t�l6�闝2�4�³��ɒ\k�4f�e;\B&�
0!�2���4F^�%�����,�6�K�1u�mf�kŖ!*��4�f&���#�c�G]��0�B�ж����������N�`�vv��;]i�ƹڶ(GH���^
Z4�͈�+.\��D��L:p �1�lK���e�T�3��\�X�ޫz��w`-���U`-
�M#,�YF<&f�m-�����g3XK�^��� Dn��ԋ���j�H,��&M��
!;gh�ڢ�--4%��Ƒ���MEk������!�mH�GE�Ab��g�ImE�+w#��!�nXn��ZgjE�(�X����A&.:"��ٙnZA0F�t�Bb��1�2�qus0�S��l ���f�-��s�Tƴ�����"<�����u��/cB�KI����s��5�2��m���blʑ-�����ز�� ���<�.�;'1܈1�im�������4�ɃU��E,����L�Z�f�㱆Q�t�����ЉLa�낭s3w1��
Sr�xK5�8&�[�i�9%NLj��bbʓ��80]�h9�*�N2�Qj筩��JZܹ���nGcU���;�V\jamE5ee3ң��uЃ�VL�Y�kG� ��kL�������Cg���[6�h��u���Q�g]
GmM`"g�P-��`�n��h�n��V�G�.�,����"1�[�k��G����9��qV7:]l�	e�Y��hӝY7@05v��d�+1�m�E���r:f4���LT�](��l&�ٶ�AV�B���8�܊D���h�d�쭰-�(Z�HU�^��ЪZ�gE��Z&���敦��W$�olה�Z���Vhf�fƴK�^�Rl@�szƺU�"�P��u�5��ۡo/hW=�z�Ic�i�	�M�#� �s�$�+st��l	�׍��a�YŲ������� [��4u��&T�!�#��af3p��;Z���]�]Ģ�Mk��1�X6�ҙ-��;=�d�J<eٚǊ�6qV��Y�BK�%��5�Z��6�f��]^�KP��չ���
Jк�3��U��lKR\���0ٮ�6�]0(��2�b���k�"�V5���p:��Ɂ�p2�m���0��ș�va��II�3iLݢ�M��R��ҁ�������a
J��)�Ic+f����f��m)�T��6tu&oS��6�[���r̰4��L��lT��A�6-͵41Flظ@ZK�.����;d4͂��,�`��;�(�K���1���C���lԄa��b���GGlMZ�#��ˉ	u�\�qgKb:�\Ԑ�Y�. #�(sWLM�!Q�Ֆ��s�fݰ�6h+���B5uF��Yz�1u�4���w,�����̈B$&fڮF͘���E̦֛a6�5M�Y�v�,�`�n�#��I�\�.��giV�	%.���:`Θ�5'l��]̸�ܛ-n[�p�`�i[�f���m��iuG��K��;U�5�fdB��0���.V=�rkQ5�b1)y7*�3,ue�е�1�6�PCL���MͳN#Y�Ԯ�`�\�6�i�x*�*ٓvL7#��.E��[���WT�;G:f5�)5չ�1�`��R��m�1r!e�فa��Q� ٲ��Ʊ�ܨ���jM������-Q��A��]��er�
�@�su����v�F�$�U�ٛ[D!�Қ<A���M+0�&FZ:b���&ڔ�n�]@+4/SJ:9��8���RY+YXVV6)r�rp��ε���XK-*tt"�w;��%2`A��hD(&�t�-�V�D�Di4J��B��Z�K��^b�,��Ls�m�a�\�\�f�a��+۳�Ј�K��K������#�Aas�Mk1�"+ck��\������]l��6�	���pպTc���-n-��gjKj�3(�=���K�,E��K�Y�u1���8Ya֐��2a�`��EфÝf(ʳX:d������hS&L��4!r6&��C)fe�qf�
�Ȼ���j���qcc������v�p�\�MLU�Ίq��0"b&E,X��Y�4��!j�.#e1L�풘���F;X�,����Ԇv�U�AV��@����+r2љ�-m�-!�u���6��6e�g��J�Vl�I�4���KT�-�K��s�3Gr�NkHT�YF�AuT�b��)nΚ ]����qj֏KA��\7K1ra��TИ(�ַZƗX�z�	
��6�;f�P�#�Dᘪ��Z$6Ҙ�[FT+�h.��r�� ���gR���n�m.���ɥk��[k�����4�4�Z�-��0�.k���lh)+���ؐFu��{$m�����k�B�%ֺ2͡��h�W)ef��8�-`j���3�e��k���MR��fb���cSX�!��/b�Z���{,�%�ed��Q���uCj� ���y^A�TK��l�V8΍���\�J�F�9�6e-��� �v�3�&����Eש���X�C �je��`ř!�,�l��+�<�ً�����*�av�,�\:%9f�K�Ncs���464��P���.�G�X�H���^f�.��dvm�ff+�JYiU�h�56��6�P)�B* ��Uim���p���u����T�5+�β�L��)�nSV��޳-�.
Z�֦�v�`4���n
��ٱ*"j��aV�)a6sZ�M�K����L,���-hȺu�ַ&DP������P
���tr� ��Ms�z��5��&phč�v��J 5p�1��X�⦘!�Zm�T��������EX�n�lذ�c�gY�b�)Bh�@��GJj:�L�[0k�"�Ya/G����r��&��i�)bX�(��AY
G`�
�M��:�.�؝M�(a5ɒb5D�b�٣JH�B&uɷf[E�݊���0h�@tH���+Z%�i
-�D�d5�Ih�ƪ��ƪ�2A��d�\�,�L�d{%]�'[p�����l"�@��P���)�Ù���5�t�D�ͬ���mp��6�m��r��q�*��Z����v:�	����kBg+[�L:�t��5V����m΍T��6���6�A⹢�ms��-Ƙ�"f�4,ΗiJÝ�Ԥb4�gnF�3H紤��9�)�+���1��:Z༦��&���[-�ۮ&p9))1��+����fa�,Lи�e��aV��2���-�̶j��GA��1�μ��T%S7&�Z��imB�p9�%���b85��
G��,�Bjk7<��a��(!5v�Wa��3)�h�oBP-GR��*r]�R�
77e��r��Y���s���T�feK,��*�Џj�k5L-��Zhasm]k ZK5�뚦�u�"J�@u�&*��S���M)���ۍ�6��\�������uI��%Hf�m�0�qf%�^5����%e0nƩM�[��q�͗F���8M���&�6��j8΂P�q��A��4�I�b���囲���\�fV�+���nܳ;�n��
L2�O�����UD� �E_�MV��8 ��UZ46ɪi�j��"��(�c����',��k�$E��(�ض5��cIQn8x.1��j�`�E1%h��ck�(TQ���Tʤ��(���Y2� ���(�*��`F�����Nb��y��DD�ڢ�(ыm��5����n@TLԊ9�"��fW�O��$�ڦ(����4�Mp�"�"�t͵�i4Q�QF�h��(����I�b��I�G� k�p+�TU���F��ETU�q�MN5�DSj�Q3�;i���-�c�#X�b$���"6F�H���$DN�������)�j��EO�a�ш�AIU���H�)֒����g\Y�����D@��-�*�����!kC��8�"JH�.6��kV�Ί�1kOU��C�i1W�	g� /��5v���6��8��cE����Ġ�.�]n#�ktWG�D�շJ�xЛ%K-�A:���Wv�.�.fQv2B�)K�j�ѶXn�؅�0���
K3��D�N��K�王[�c6�֮n)F���cu��kcF�h�ؚP]0����0��1�R�Mq��
��3 qI�^�K��\�f�i����95���h�]�]\�q���R.���ɶwZ5KSd*٭�Ik��K*��cqM����l�Σ���
�����L:�E[�ݬ�3�!��g�,Z�j��ݗd��,Ќ&,[�Q\�k�ԍ�,ь��4D���-Z�u��\��u�l��C�<�O<�hcD��o%��2�CsKe�M�v�4�������s�w�.��Z�`G8��`�5��j�SF�܄�r�k��r7%��@s� ƒ��tj�w2[�[�iVR�bVV˓�K� %��І�M�l��CV���XVR���[v��Ή�Sr�ʹ�ƅ%�m�G6�'�k+�.�;�+m.��dI�+��U��SBsm�I2�ŚCk�To��&:�%�,��e�V�V�#wd��b�\�PJf4��%�K[ln�� �T;KR����k��[��-Ԉ^r:k���cjMdY�`f��fR�FfY�]u���5��DnY��n�0d[��m�����(.��[N��\�J�lh��ζ{YMm,�X�\���k��6�WQڍ�1MI����5��,6��O��G�m.+�k�T�Fi�h#�1,��*4��5�H�T"�BB[4�[sQ!uQIL�.Q���5��ʐP��qq5HR�9��nХ�`l�ٖa�l�nhQ��	j�BeĻLY�aײ,]�hh����(��&Q�)kd�e �JQ�F���+�˸� �=]�pWF#3k�
8Ф,kM�3�Wt]�Jõ�!R櫐vi�4�*���am��n��1� �lȗ;aH4�N��L��Q,(2VJ1,-Ez��T�l�#i@m�/)l�痋���@KX	H��XZJDF�nXX�4��R����y��!Il ��B�����F!F[l[,VU�Hx�"KhKkkF���J�Ij�!VB��u�X5��D��m%��h�� �T
�a`W�@�^a���e�����ԂRX4 ������M�n[nr���H'㗗"�1�"N�;:��>Ws;����;}�7J#p�:��&��A^�]�e5t�(FMH�$�F�n�H�l�r�V�.w͆t�xW��{��v����4�����\���P�=1�����7t(��4r(�6e@�2"~*�ڟP;RZ>[n�VP�� ���H�N{�Cj���>H����3u��V���sC�~df�?n1��;��9�u`��󲷀`R��I�������㬛�?Ӓ~ZT��Be�[�٥�0L�4&mÆ�]�2�$�B��$�Q/7cfL(`����m}D�yh����&��i���Wźu�+ޞ�b�swAߑ j�˻��0?��\���(�׍6v�+�y�.|�3.^'v�\қ�t\e�/h`'!*��w)����X��/r>5�0l7l�.�>���@��&_�	�{_W���m7O�Fk��c��&n�F�@���+��"	��<�@�k��ِ�7����{:~���hWƆf
dB�H�i�<sG�>n����#iH'��A��W����P�՞��'�ܚ4	(�6e@�2"A)��>�@�H/w�*,FU�j��'�4k�t7}�(�A�m�v>38��¹B ��- � "�ZJd�8��۴#I),h�,�*������{��\�2f���La������?n�]�Pݝ���n���u6Ew��Q��N�zd��T��&_�{n�giM�̛�C�g!��y"�$|sw�(���c�Hd�Y�6	�Eř�*~�A��hF^ТA �g�Q'�&�Q��b�_�<S�E��ȣbv����>S�"�z�N��h���s���f�����o�8'���&~����xzΏ=��J��H?���7w�N�dť!��#Qy_�;��������CB@�y>��~�l�˯G�י���(��4"&&$DP�E��h���
 ���Ǫ������}@�{~{~B���I��Z~<j�RQ��b��1���H.cHƱm*sR��n�u1���e�{���	Y�.���^g��$gM|aT���^�����$���"f����S%Jhj6����ݟ5�!����C���'/=5�?)�-z}�?�!A�ϧs�Œ&v�̕��1"�`��TA{HM�YҠ���]l�3J<0�3/�����<�&���^ԃ�__=�_�k�߳ ���
U���=W��t#A�����J��Xs�c=-���>z.w�����K_�w.��7n��㿕��0`|��kD���WPY��˰~��k9��e��������t�F�����z�0���,9���\-@�~o �{|�~�����:^(9��c>�MDa
`���"��%�D��+�R0l���55AK)^�������s�ܬ�̈�
��6�L]�@��E M��d�W7^R.�~Ֆ��I���	�Eee�P$L��J���	{;~̡�)�0 ��x�?_����p9ޞ_�����/T�1�`�[�%nj�$������E:^���Fk�O��(P$7o�(|H��C�ID)�Q!�x�ؿ�Ԓ�4W��D�N������~��	zp$���!6c�I�?$D��.D�c�{n�9a_���ؗ#1���w="���Cw}>D����xB�"ɑ��%z�{��@+��m2V���>�����0/���/O�����x���s3=����� �@(�i	e���L$l��a��v�=v��[��s�`L������<�(�l�b��.u]�-��i+�Vky-�15͐tzh�(k���-����lF�CJb�`��AMq1kJx�a������j�Rijm���FgDs��vj����b�[G`��+j[����`��fDѶ�XB�$����l�Q�Xf�h��f�5��T�k�R]V�ĵGl\��1��Y��zص�,*��Z-`569%���'|����-щ��ϝ~��zh���m�WĒNT���͡@�w���47�133"�
DW�u���B��=�s���{��w|���T�Y{>����s#��7C�P���	M�uT+�A�uD��e�!��D��O���D�~'w\Щ�930�#&%	 �ԃ�"�ku)6���C׶E H'�~��TA��B�;�[�vh�Z7��(�Ò��2P�l�:��$�٢��#�(nk�f�������[���͡E��N`]Mm�K��iXF]mι"�X�H�)�x�lX��Ů��I�B�-��޻���f�7$M�k;�={Ѱ�O߷��k�����n���㗮��a����!J��6�ȯ��/1�
y�����W���8�ǖ��Bec�ⁿ�w�Z���2�iưV�Mg����^�˒�&sab��x�J'�J�����˼���$�s�'�D>�������e,�J=>������d���XPGqO��9�?�~���=ʹ�M�+�(�IܷB��v� OӴ1����ո���M�uvk =�y��L_�� t [~����kd�~D�yU3f6faJF$LJh�� ��="��غ�ї�r��B$fn�A1�����������.������J���[���8A�����Q����������<��11�$�^r[�aI��Q%���t(�"�&�$�е;�@u��X�~�u�UL_���^�T�S�DJ��_m�P�2��糧ܘ75B.�$��Р	'쭺FY~�Y�'����װP��R$D1*�ٲA'չ"� ��+�uF��/;�y�ehͨˇm�R-���/�F�� ߮�i�tFq�����|��+x�d{Ե@�/X�WJ���᠘˝,0��گ�F*L�Ĉ
)_��4op(v����H�E�ݡ�d��ˡ"�D���n�}6�����D�R����hE�FD���b�*�{�/�yl���"l���n�hP$~;�RAktI�{���\��XlU��6T�sR+7Q��&a3s�7#�i�D����߳ߵZ�f1(I�p��@8��(�H�ڪ=n�p�z7V7jE����
��iV��0�J-�������E,�^��s8A���
$�o��ѷ	��&�>��M\��90q)30BDJ��Q����U�)���DmM|H&��
$�گ���\LL�LJ��^z�"}����*�	�	�_����?s��t�#�=�&�Wv%;���ӆ&�@��_�)H׽m�f��Jz6-�t��V�nr|(�S5���"�+��X�P�ꍊ�4��<�@����O7un,(#��7k�o~oO�W.h�ܲB�t(Iۺ��~���XjN������������!���f�4�l�6�8�RR���ցv�{V�XŌ5e���Bo_���ǳQ���c��C�~�eU~'��ݚ#&q�,�+��}���${n�Q���S2�#&%	?b���P�R���!�'ە4H#ӻ4	 ����}�ςq3�P�an�n���c�~�D�}��N(4�w.�i��mh5���`�	w�_P ��͚ �����I��2TL�"���Y:=��)�� T�$}>��A?kۡ�s��:�I٭�D%ࠢ�d�:t�p1}^f����w�Z�ȗY��������A91�����������z��K��Z��y�7F=���������,�?ב�{�_Q�-l�%���!w����i4�Z�Ǒ��>L��j����
�٪�0�� ������ݢkH�4e�S�y���,Y�l��#HF�HZ��W`F���ŷcM��M�{h�+�źʎ�[�Yin��f*��If�$1�lPҖ2�#����F����z�2δmt8%�[av1U��Х̶��sq]�@j��ғ=[��L�,�X!3rb7�4Q��qi�@��":Q�J2��UcLTY�u����k�j��+�[-�ѫ�\�&%�N^��v͢L�X�i�@P�%�j+�m7��31"�bDi�<���Nʼ���O���W���#\Y�S�#���~�Ln�����dHQ)~�uB� ��f=YN���ڢI��Q
����}��:����=Ω�Ԏ���4g���O��&�fь��_��H'�j�����sǚP[�V��]���/o=�tD��Jͨ$�����|I ����n��w���;���t�#A[��{~�>X{������sD"�K Osǀ`C�ϟ�O��ߕ�m110�z��� MuBĕԡ5Թ�bi��	f�]f�ҿ^��QF�Ɉ"�RkA�O*	��>���AЗ�n��p�5N��z��|m�dQ�8�*$@�&$@[W�?�f3��3�g�ݯ!D�o�l�4��[�/	/��� �EuU�Ҹ{$`��j��$�l���Χ��M�R��d��7ty`�^�箍_��N� �ˑD�����A�#B��.&]謜U�5���#"B�(C9#ĂA�k�(�O���Tz�;YX��]
 �~;��F+�*`�"d�4F�R���K1�w�MVԊ I#o]Wē��N�^ڕV�%��ϗ�k�,LJ�&bJ41�eH77stmj̽$E�P$N]�@�E�ΐ������������L�,�AM+[�#X6�֍�u��T-�\��.�����_F�(fL���B� ��P�H7;Bta�"����w����2�|I?n�Ы�AE�А�wQ� ��@�����~�z-{��Aw�T \��tU�����9s��t�왨�ŉ �y>ﱏ��elid���������n�d�:��1u���	sn��͎=���������y�	�5ڼ�G7Vzͩ���Ӈ,�^��s�	�s��~�YP��b��a!>��}� b	׃������~.��06̲{�����hs'�{H�!�؛h]L��)���>�vԻ9 }Č���]��;٬��i�%ܞ�Ϻ �i�E�Qʵ}���/5�]��IQA�&/0W�.�ǽ������E��>e=G�yg��=�~�"of׊��zh;��2��|�f����q���ʼ�8VCb��
nԬ�����/=��#;�b�k%U����{���f�k��m�[4�{��d�E}K�(|�@u]�v��ý��M�8g�˽��h���T��z��OD>�)��ov{����^<�:�͋����k���˖v�9�rY�}�p>|�\�&����cZ��gQg�n�@�>�Ӎ{q
|_[����_.=��_��!����(��9"b)t�lE�����]]������X�{�����0z��M�U�}ޮ��7�S7��~����5�[j}2x�����yC�e�7EO y��L��?�Ǽ�U�~�yQs�c���ӷ�|�����ɩ���dy�����n{���7ۛ_`荕��_O.�o�o������޸M�Dg���a}_�����@���:\~e0���+ܸ�8�>��A����$[��`R�a�>\캼���1$��)�)�B2V���~,!��b�h�$�M������h)�t�A߃��*5�XT�L�Q)M8p�p:�;�Gb"&��("����2"Vd��/��Ա���D��L"1��L�����HX[Q�F-�q�S�[̮��1I0��$)������s�O�wu��h1"!�TG(���)a	!!l!�-�k�0\��*؉��kG�8�A;$���de�, ��H�F�
RA5kVƪ���a�4N��(�m��gEm�cQ�PQ\Fh��6ccm����.8�T�U�l��4�5�b����t�A�DZ�TQT\EP�-�1�6�ˌ�*I Q���jt�J+�q��ic�S��F
�L�E�I2H���J)�8�q�ZĘ٪*��AZ�JX(��Q3�uh�MUAb�4�8��� ����g!,����Q��IkZ�*E1ʕ
�5����f
a�s	!��׎]e)J�y��>�D%^�6�y)�&+�<G� �����W�g�y�����| D#��y���q8�JO|�����I�4�\�^�y�̽os�w�v�im��/^��r8H�����a��p�{۳j7k���s�����5�$���9�������Nݥ����k��H���"�nx�!���@i���ϮGJR����D��|����KjlO���~"�`���a�<	�(M!Y1�գ6v*6l�����ںX��w�����ȣ�u#�O��g~��,�����N��\���Ϟ޹z	�BbG0S���])�&�|���y~����w��2����'�|�����$"@�w8}!j��m����@�{Η8 G"C��<��'���'���N�^���4:L���>�RiJry3�ۼ�J8q
������_y�`�����Q�{���!}
f���i9�߷�S��S;)�a>w��g��F!�R�<��|]�|�\��x�)!�@i�ߟ~z�h:�A�b3���Η&G	��{?G��v��tᚙ�p��]������z��.`������:C�(N��y��JG��!����PD�ut�x[s�_.��I���)��ձx��y	Ǭ�y��5	��L�m�L��.������[��D'č�{z��b^�<�����?��0C���:1NIIο2~����B����<�����9�9~�/�C?Dל^n�u��?|2j�̤@��뿾�s3�^��~�@��:���ǓR����8F	��A�,� �Sz˴Хb"��b^�`5���D���%+�����٥[��w�9��5��u���R���Ϯ��0�R�!�z��W�2? �ٻ�=B��A3;���s��xe�it��~�u)K�����]6���<q"y��8q����I�]�s�t~��?"8�#��^=��N�1iJ={��������#�!jv��o����1O�$/��|ĵuc6������3�Ҕ]>z��^���"dp�}���8m?���?�z�&)�<u��ne�JR4{��#�����-�~�]�n���p������:��E����R������P:�&�Hhǯ||��:$4�8��>|둠�����\�'����RC��}���#����=���YV�����4v�����'R��K��v��U��~T+ �x�,���?�(L{��~z��Кҙ���|�묡(�E|@��·���$`�zf֊TM0Wՙ}.}�G�E��H���ɧ�/Q�xo3ȃ��=3�g�*��Sܫ]� ���i�c?Og���l	�^��O(��-z�r��&TD���Ǐ�c�|�P�&nKB�%S]�X칛\L�QF�&�M��K#`B���c�K�q����1v�tehJ�Rم�ĘQ�e�6Z��]i[S2��m@�%��	EŊ�FY�D�5�G-so[�&���)`�%�78,&�WL�B.��eq6Fъ�@-�\�d���7��m )8b+��Ie{^�]DV(g�]fi0̦C)mM\/���D��Z����ڑIJ�R�5�E�!nᔭ��K�o;��O��M6-5�`z��{s�\���@h4�=�޻�9�bdDro����p"g��^��<���w��x�t����t��B9��
~�>�`t�s�O�viV�wSy1����C�~�4��z�ɻ���/Y�V�|!Ӫ7P�КR���{�:����ӈ��t>$���G�~���ϧ��sΗD��7|����6�����|h��s�D�K���I��uW���� B?|	�����"):̡:�&-)�c���C���)X��}Ό\�N_�ξbJ:�M�s��9�?k����O����@4]<o���)I�t���~z�hzI4�.g�~=��/�^����z������#����y2pN&���lo�˷mם����\����1�"_|	�v�Q/�>�8�pC�;Hh�����:��4�N���y둠�JPhy���\�tä��ڐ�f��w|�(��L%30O�Dn��[��E�  ���m6##�Z%�sR?�������YV���M�;�9�.`�v���<��C1�1ϫ��Q��u�M�9m�����x���#X��v���<�Hhϲs�2~}X�nm���/��:\� �Ȁ���=�=>2�ƹ�,��{G,K�x�����Km�^�]��L���̟�0�*/�O3�^^�0
 �H�M��6lХ���|}wǲ^��!��'>���#C�I�#�s �_y�:\�D�p>��/v�dW*���d|1�<L����"|�;�N;���)�iLl�	�>��#����~�7��/�����1>��޵��JS��}�둠�A�t}��t�p#�7}���&���>��":�y�6e�0|Vo�o�����A�):���<�v�F��1Ͽ>��#������A!ܻ��/u]���,����9��ъq������$����g�É؁��yΗ8 G0PG��|���}sYQG^}����)<{��F��4�.'�}��	 g�~��]�����d�����B�W����t
M��A�iY�:�SP+��k���4f�&LL��mЙr}{�=A`����i���:��S�қe2l'>�z��L#�(�
O��w08�p#�{t���sk�َ�Y1\ �� ��n�Ā�?|�G2&}��t���ϸ{?rɲ]VU�p�s���c��s'�����u'��F��:�	�}x��T'M�#�O��w0:s�~뾝��7�g���}Ό\�NǮ�g��c�Ź��ӱ��s��brB9�>�}�9��� �G0\������������n���v��Rj���ޛ�s������;sG��x�ky�Ep���|ę�c�y6�"*���r���7��������dҔ��|z��4�A�2N��ߧ���bq0���~���&�u7�00Q�F��|)Y�0J�t��g�?|4$0�s����` A�I�}w0�G�@���·ā/+0Z�?�:B�����\��.#���3�|#]7l.���;qp���8���~������ﯻS��w���~��0��s�a�������{��0�cS��w�teN8E`�.����4��iE�%����:��y��y��u���\M.6VdMe�L`���7ϗ���&�=��>@�}�K�.`��.����门4�LC��y���C�#�~�����fqz�V���1��#@����~�K��B9��A"w�h�a:���-%��7v��0���/ߺ�?���	/�����j����|3'�D��քѤ4o;���Q�!�"r}�Nuw��8�D#��~���*��<>ڏe�G���C�8(J�%)�ӆjg1�&���ÎpԨW2!���g����\J�u��;Gr��$�䒻�0�h��1�Ο�!�qYIFD������At����ʪ���	 ���
a"Q��t�I%^��4��G�N1�_�Ч7��չ�|yt�m����^��g�"�;�JՕ��Yd,�Y� ��\���{��O]��1;�bV$�++/��� �	/�]y�ӑkh��S'�4���� �5��k���Cj�|]�����a���$���t�%^�a��x=#gS��y��(��d2��ʶ+0코%�n�Ѝ�6	Xl)�X[L�B
�x��x""D̡ς]oi��H$#7i��I$+��6�ޠ��T�l��W����_��D�8}<`�	E0�y�1��n��uj�{[��ť�YUO�I����A/	�oR;gj��+�XQt�����v�5���i$K��ZD礂�}}^��3J�`E��B'����/��i��v�BBQ�ZS�u���r���I|���Se�I;�a��D�u�S1�:��h�0F��I�
ZF�d)����! �����{����q�I��w:i �	�s��I��`6�u_�,���^��@{tP.�d�ٰ�	��W��޽�5���?�n���r�+k����v��$�`��E��ly1����ÿ�i������?] �٘�]٬26�tVB5!��!0���r˂�*�@��J�m.�)����m
�u�ز�T�X��c�1�+���V%�V�-�`�S.,"i��I�R�v��e�9n\��͋��g��sf�.�k�h�������B���\P�����ѥ�h��۶�7ckm5��(qJ�1M�Y�MW�TS`�2�E��W4���.p荭3[kS3i�q��`#�����3 ��ɡV���Ͽ�L�%0g�=��ka�PK�ٴH�_o{�l%y��5<}�x�7��1�_/]s5Ry&�"$D�-�%�}L�����u_I�N�o�K��a��5ݞ!�(k�S{>Kh8�	IHIJ��}|�/�_%��O�Ho��]/��s3>���_���+������a��y��D�_���-8tw�H������{�|n$��^L��Y��I/&7�Qc�pq��x|���Pm/���Đ�"A$9`%=�L��D��`�4�j�H��y�����o�l$�Gs�A��	d�ꆖ���ؗ�b��˼��o^}�G�z����(���땻mb��6U�c�Q��mPб������߄�(����*r�w�/�A,�m0ZK�J�&kٹ�z�t]z�J��_��ĥy�b�G#�(0g�4v��H%������^��|�X�xS�y^�e���vͨ"���E����z�~�0��|G��Y�٣����M�lS$�;iK�K�v̊�O#ӘUG}�g�AYUB��Y~�H��Lo8a"f� ��u����lkU$��l""DL��=���ZI|�J�%$�K{ls��jUrg�2�_ �W~�(��Hd�t�,$�1��a$�$����\�0�g��wE_u�I%��9{��C*7Pe��	w�/`�=�WU!=c`�� K�VX�Q�"c�0�~V��r��"k;h0�*.�lר��ZH{Ϙo�J./?��D ���0���\�V�����R��6ԈP�Y��i��4(��]]ƈ��v��i.stf"$�O`9�L�aD��	M��-$��[�� A%^�a���9wuQ�ߧ��mc�a��I!��0���K hF��]�����h�Q�ݭ�F]����A$#.u�_� {y�%���u�9�l;ԛ�hߚ_T�T.A2�S~��
s��	/��ޠ����]����xo�(Gxp5u]�RO�'ޙa�XZŨD�d�c��\�@H�n/VP��0��������$Og	ٻ�CU�Q�ŧV�}�#�G�����%��I������'�a2bd��{�.����DM߽;��$O����D���,$���1P���J���в��m4���zF�B}(�):j���/��g{i�Mo�ޫ��:g���wT�O�E1��i%��-��V3���'��ć�0�����K��L��@\�Cb���)	t:���TO_�'�{�;u\��|g=sD�I'��H$�Hw>a��չ��B�{޺e��I���,sd� ��B+sc���bK��6������{��w�5�$���݌6�	+����h����x���1S�]7������	l�2 @��ࣛa��I%���i$�򋟽�Vq$A;�a��I-��0Nt����A)�?Aml���,�wp�b�A*���R	/�W�Xm$�Ot��	���5�b�9z�Ysg#��3��nj�
9� �z�=o�����=Ś`[�{�����}���EI�1�`��yg�C���X���烿;�s�i�j�"*�>�V�r*��A��@�ӈ�"LL��X	u��ZI�s��Kx��=�˧����zw�В�|�%��1��I(��e��k2u��m��~M�K33YXh0͠�X�Q�i�҃)5��QHjM]�y�}�=�f�$��W���(��_%�_��D��L��_=\j~��%����I�/SiVh���´b;�j�oǧl�I�]��x��\9��TI$���2Z*3�Yi%�>�{Z2c�Uk��04���N|d̓&Hsc�"�*���I-�٦%%P��{}-���8*;G�0"eϹ0)/N��i �jW`P���{�(���	NW3�3�$�T>p�K�o&����}|��vs�� �;�Ȥ����E��*�R'�,�o����.�Q���z��f ����a"WM�2�I$�{|��5?|C�1�)fK����V��t;�3z�E�W"��>�tc��e<t)ŕ5��K7�ۡ�w��~ΟV�z_v�9s�%k�;������{-��0�P�X��H���l]����:7Ԉ��w���^�|��b��g���}�!��3
�[���^/DY�M�8*A�3��[��s��=�h=�ϕ	��-BF�>�y#�`|�L�9��%?��� ՚_�')�Q���|��*+��6�k�`�T��h�~��w�[�3 �j���o���[=�D^\�+�Y�,k�>K�w<��b�'��]���F{�H��n��o��U=Q��!��L��-w���ZOb��ލ��cv����{;Is�`<��v�:���[Ǐ!��i�
y����0�����{�f�3��� H�g���aUc�����\�s��j�aɞם^"��YN��y5 U�Rn�9MHa����m]�W��5>n$���f�M^I_.����k��I�k��F����F�k�-�8	˽飷{5��_2�]^�{/������{�˗�"؜�G�.j�s$U匓Y���$z߽�Y����B�<��x{E>ؒ�PwX��yQ)�FUߍ�
̬�±e,O���L�<��ݹL-Ї�4I|�:t���e~S�8���{5��[�-���o��W}5/���>�5�>�h�V��a}�;[�=��S�U�(@��RR�ޙ��n����$"+s���udS'�����Y땳f�d�Mk�������=m2�Ǘ����ܟ�!��L8��n��3�<���B:6�5z�E��S�\��jeU��B�
b��1�$�EE�p�B���t��.98��DH�28���W��*DlȋfE¥L�*�".W0�b�p\�2."RTs���5*��G��I�V`�P��$`����8M58���9ei�V��#i��Y�ۃ�@�@RJ�&d����K(��a5&��J "Q���i�[&�`�2+��Ģ��dEl������D�� ��hY*k�+dd����F̊�4H�v��&�KmU�\MsPcgĶ�lNYz�:���[i(�����[k��V^[Ji{l:u�rq���$ƹ�WAj��m�,H#h�7H�:7��B)%��lVA]%TVBb�e�$��04�r9� �"��T	�WB���6�e�m�"')�k�fL[E$�8�).:8�J+�浤�J+�)7[18#l�,�:F/﵂15A���� ��6�4e��n(.����ړh�q���6�(CFЛ�X�i�����bb��0��˦TaL�2���l��R`j��,�Y�����q��t3�%�n�L��,
���eWj8�E�q�3V[��.S-��]3B�(G ]-bW&�)` �k��N�����)@�Ý2.sM��B��V	�k�hg���.���cm�]��YzгGcL��W�Ò��@������,7<�sKZZ�BX%�u(f�Р�T��//V
GѬ��t �8��8J��J��c��gR8���Y�X#4���M�&t���[&e�^�"m��L�1�n���H8��V2�I\8��ZFbښ�a���Y+sJ��2�%M��X�9]���Բ���m�jF7a�v�3v!�,�a��T��iDő�.Ѓn�5���X�!:��]�L����6��T�	��[C9�znY��k��av`eт��)	�D(��s�͡.���+F괛X-!p���ik��R�9('j�c��ƹ�C;B�&m2��5��V�̺��9��M��AHt��(�P�v���A�[֚Q9��l*n]���� ]�-	���Υ��,v��ܽ�`����BǬ���530Yp�I�a�!�̍LFE@�:ș�f��ж[���%�ʭ�T��Ű��]��]e�V�	+-�Ñ ��G-��u�-��Д�6��*\�������C]e� R�j�ʖkMm5��%�ґ��	y"]]���@�XB8ӝv��g,
��27�WZ�v�i�	a\4��$W&R�LFS�u�],�"D���y���[����ŷd�.%�����e˶�\��ik��p]$oW[�&���!���δ��V&�Fk�T3�kو��-��s��&ƳKɰ����d*�ьY�Dvu�ѱJB2�������.��m)]�@�U���A��3��ֶ��K]m��������BBG�<���B��Z����ՌQ��rKۊ2��́ۉfz�<�0���e6ڹ]��XTc�Mk5�tq��kX�q\0]s�j��X�[W-�݉��]2LmWCe��$�һ�RX˛�i.����U0݁4��T[�hJm�͔��;\i���I�n"�����1"P"�Bf;��m�/X�J���h[�f>y�cd���P"�]��c��G`7��*��iY\�X�i�v3 U�����┙"d����Kn8d��s����I��������hw�⋛i�+�N�2��B �(�
b�_��a�~�{��{��$�^��e��I'��0�@$�ܰG�wº֫���T}[�!IQ���F`{�!W}T�A$}�A���$�:�bM�@�]�Ւ�B粙i/�I�����s��&D���=q6��/���
�ϒA.���$��{x�%���>I���ǟ�>	,�u2O�:�q`�IH�b�����DB]p�âo����G�W5��J�6�a"POی0���;��0�h������bc�!0	;��zʹ��J���1{K��ee5�I��z��m����2'�:}�x$K����$����~	2�v�@�{���>�2�D�۔Jd�R"��>��K��4ϥ�(:�=��R;���܄��D6�WK����?��C�����Х��nF(��]��;<=8���fo����VΏ׿;����c�"`����W�D�	$����IB���Q$���`θf;&7�;��>�a�D�()��
���$Iv��M$��nw{z�mU����_%����a��Iu���O;��!*>�3*T{�M�K�6��]B�]��]x�8q	 ��k�i�cy�o�y���`I�\���üO
�S2fez��8�b�G�[��l磔��[�'�����6I%���)%��I�u��D��HD��'�
�S"�q��[q�AN�5y�R-iw�P�s�|���۴D�!b�����h��\V��}%�H��p�K32�}9^������� l֦P��$��FD��[+�ؔ��y��A��P ��\�&KI��pI.=3y^ɥ]�uF�r���iD��q)bd��{�,�z����%��i�)�^��>�����G�ly��v��qvO��f��5d>;���ޟ:P��G���ᇶn��-]�g�fs�W�O�瘽�@HfD��~~�����D������s��Ս��n~n�����1���H`�:�P�@&d�O��Y��5P%kj2�e$�Nb��,��Y+:���������Y�����l	)�� �:�{�Q���S�m�I"^d�;�Έ�t{��d�M��	.��p�_$���(�]�/2�J��DR���*3]I��l�����҂1@ʤYn��su��[�k7�A�|�8ur��x��#mS�$��ͧ)$J{��i]�͏71gu+�m2~'����L�ǒ�ؑ'D�j�~�cjers��k�_zc��I$�O�m�ÿD����{;��CD��N
Y�(ȟ�����>��_$�6� �J�5k]�`��zI-��p�I ��i}����	�DLL�3~��Wp���>�~C�[��LJ_$�O��6�I-�>�g�<ڮXN����n�z�r����$�^�e��~��w����?n�,9�:K^���R��1~�=������tm�.����/�Y�(R )���\�>��	&�|�<���U�	�AR�W����H%��hT�e��c�K�q��K�K�������I�X�kr��ꚽ���``Q1)AFjJ�L��F7n�vM�̮l&��sy:�n\�����$J��TĒ�w)��఑�^��<�H�P�a�����?(Vdn���I�����/�:$o�`��"&S��u�?�II�������)}I���)$K�e�I�\����պ{B3�$�?DG�&R @��V�P߃I|�]u��h%�=+4b����.�������~�a�RH.��P�0RωFD���^���*=:�ԒZ��H�]��)�Jɍ�����p�OvW���(�����"��>��]ok�I$�Wm1+k�z�����%��M$K�\�h��V�C	{��g�{�.�_|	~�OSF�
����Șfo��'�<9�&g��i�N�'kZ��x��İ����2ey��F�� �����=��@�D�"% R��y'���PJR.�ʩ]J�1f�8�e����3�f]�kI�L&�AЁ��B�6�acJM\a�Յ����̳C�f �e��s�DMb�q���je��s�t3+��St�ö�+�����L��u��G4����6(���tau�����Bk�гV�b�2ԛF�ee�c6�4`�kB��ܔ3S�g���
%^�h���e"F	��ZЎŮuR��	l�܅��{����+iY�-�_����I$��m18�A1��X��PW���/�޶���X����aPD��L�I({�
o���Dzw����Q���0�H�ek��B3g�%���{�'Ǫ)���]Lg�.d葟J��T��N�U�t)���Κa%�K�ە�,�|�c	/�@.�����IFwS'������T�&*�(�lvR��3�+�H���M$�Joz�a$IWv��.���j��`��v�P��%�����,�&���/yeʓ�^�07��6�I}�Ia$oc�y�ur�Z#�8iߠ�	)L!1	9e��k��B���7n������il�`O�������ebd���#�_��0Y)(���D��wc���6B�M�V����x�h��f�2��/�eY�HF"BA"'���2��=�i��"���s�f�ϥ�ǽ^W�����^{t��]]^n��A��hwp7�q�o�����xL�3�ַ������ �F#V�V�o�π& D�AJP�R��]y�����E�S-$5߲���˿d{�!�����|��w�9A�	�2�vW�Y-$�ݡE��S��?ewT��A%�ɣ�$���a��2tH��DDI��S������7��B�ԐK_�j��Ĕ�Iy�2ZH-��;�c����,$���L���w	}�P*D�j���$�]u0���W�И�I
�t��$��Wf0�?$��a��p������-���?5��*����$M��pڔ�A��]c*�4���R��A�6��� ��ZWK �ۖK�$�Π�K�ޮ�M!�-{���f�H��/��I�om����.�D@��Bg���u��L$�w	؍̿{��$JI
��-%��|�|PHC�1a{<b��8u%�����H�e��_��<�+䲻)�Y(%th�����I�|�G��1�w�<��2=�`KsN�����o����y�z]���%���ط��?\���ZMZ�:�ڃ����b@�%�s��Wͫ]���ZI~���js�1A��2���u�oej�u5�$�K<��h��Kո�`$J�ަH�ۂĹ��]>��Ae瘢ŲtL��DȐ�S��_]
i|�J7�i��L`>x�����"��m"R��a��A%�L�2�ؘV���o�ŏ�z���*�
9e�d�F�d��Ys V,v��VW\!�cX��g�~�}���!Y��V��T9�I�}L�I��ަZ]>���[��}����E|�]�X4��RTgȨR���7�[	 ��W?9��=��D��$��!��$�����'�'z����������}Z(��H�)!"fe	�{�/s�i��_%�4�I$���3wf�ŷNbG��c������a�a{�\x$f_/w�m��K�y��g1�}[�!ǩ~�"z��I����ZI$�����'�)�UI����=�ő-�^gG�8c�a����򾻺��3{��k-}P�ۼvS��Fu7�`�8�f�>������`�������'<����mr�s�׺[I$�J�f�mlp��_�=�?�}��IF_S/�I[|��X�iPVB�]�=.2�������	4���F�&� ��څv�Pe.r�!�R{�>[񈉑!L��K��d��v���$�	*���.�M��-z�-�
!)��e�k�j ��LHB�?��F�P���U���z��$�IG_S$2�5��D��kí��y��hiF�IP1�#�@��
7n[	$�@��:�$�	?���5�x�;I��v�-$AV�0�K�t�2�&fP���qޫj�Q�כI�h�XI}]��%����3��S>g()a���s��$B��F�  �2�W��I$��֘~뜋>�B2��e��(*���N�O+�f�gW�D�g������!w��&T���c��s��JsRX�Ֆ׏Ww�g����S�����!�|�޻�����s�ɏ�V�Ûکg��|����B*D� u�rn:ҥ�օT�(ĩsm#WJ[R�L�-���TK�m��[,l�V]a.��Z25�c��1�ԕ-z��h�l�V-�lu�%6��E�.S7U���bLf����R'f�4�*3\�5I$E�k�3��q�c�)�m4ͪnE�%�h��X�n�+M��R�B�K��eJ��������ui��%����(,at�5�)1w8��	��B��x��3�m�ZhB����V6�k����a�X�r�=}=?��?�I%[�A��A%��W�J�	�ӨQ�ѿ%9�GR%|��a�2vL,��DȐ�S��]��`&����\z</Åi�\c��K�	!]��k�"��ŴRU�s��b�DWNiĒ�h�$F�bB&+�uU�A/WO4�K��yЙ�	\���Ӂ$�U��6�I-��-�E%D��Q���o\��UY������H�{.���	�V��?�L��畂}�=r}�v�]�a���C,�I	3(D�ĸ���&3:i�xb�ye)��x���a�%-��R		��e���O�s���W���E"��������q�h�q6�z�Xh�Z�B+�I���*b��0H@� ���'����W:�`��IFwS,%�j4���F��C�(���x���& ��%���]{���([P;%q-Qx�	X?�;��Wq�������>�"�w�>ns������c\���پa{W"��T$S��v�=������@W�}���� rw�{��Ӻ�r���8KJ3�M!�03z����}�^�1}�`�K�Y;F b&�^K��B�K��nt�I�J)���xW��co�D#u��K����$]�	�@��yG6Ǻ���2���h/�ͺc��	mv�ZI>�bQ඾�]�a!����
�IhA�,A��k�HI��Pmw�DC������[��6��$.b����I�9��)S�vW};�<��t
�)-��vp6���ZWͳm�gFjv�tRډW���z�F��f~o�;��d���i�D��:�?�����b�-A�6z��E|���/\=jZ��# ���Z�g0�i$�u�v�������$��l�k��H$^�Pmb���W�D߽:,4��W!*�OҠ{�Sk���Q$�͡E��π�>� i�t�ڔ��Mvd�M���^���x#u�.\�^;�����=^�����ٻv���U �%��l�ޏ�)7>�_B�n0��6�D���[��[���s���	��������S9p`��W����P��K�r�<��]�h�4�秒�'�a$/g	���t7~�o�_�����(��DF��`Pq�:�[�ܞ��\}�{�Nc�Oa��O����cM�t�|���"4X��z��Q��?)9�ŷzQ�qy-�����������lJ�{Ds�3��7CT�xw�AP��_y���2>i��>p��1�� �m.a]�u<�xb'ݳ:�[�N�39�٧},�����вb���X�ge�{|�b�[�8Ok�w{}i��㮎�swEۻ0�y<�c3$JYD�M���:#,K���O��H֌�����힝�}�&�������]g>��Sŏ�#=w=h�����M��~���:E�'�{�vvFg��g{�՞��{fi����G.��a	�^��-b9����w���=�(e��ٯ���.�{77��?a�{�K���68N�������l�p߼<���������r7���ym�q_get�����������ǝA��@�o]�5e��<��q�J���t�����S!���=B�i^�o�Avw����$������w������]�0d����~�y<H���0:�|�S-�[P=�0�,�z[���q��
�U��竻�5�;��I�G?�x�w�]���
���pS#����h#�a{v͍�����`��1���\@��,E�h�aE�3V�EH1�w&U!4���.u���9�d�ɶR���^H��n6�*tɌLr�������A��"Q0�87&��1�`:��,�T�8e��t��ft$l��@Ĩ��El�!JSN4.�L�!���K����H����[�B�i�NBQzԨÜ�B�� ]�8����ٕ'd�����RD����HX7@l��ԁ5��V�Ic��[������E% Jt����0[��kz��Jt�!���S1x:Xq5�!;%�D$G.jAd��dԎ]�XXZaz�c�.���m���� ��J�mJ�H�vVPZ[�D�d1�E�Զ%Nzب������(�ԉe�M�L�c	���F�(��[:)R
Y���t��ؒ��m����*��a#��*Qh�#@j�U��
�bU  >�t,��\�ꆒ	X��O��-d�Z��Q)�K��Q���l!q�nA.��L%|��$ް������g�sԢ��K2��5�`�F$!a��(��4�_%��^oW�V��|�	��nI|_'۬6�'���m{�#ݽ�uW|�_��v��7It`�0L1��΅;!{s͘6
VS^�<V&��~�����bJ�`�r���H$�w�A��I!�Ws�Շw�$�,j�r��p�I$���Ґ�M�!2be	�{�/Ou?�Ig��j���J��'Ur�	ﶅ0�K�Ws�
&����M���I���I��$HJQ&A"e��o0�%%՛B�I��*�[ٳre�v�$�N�Xm�G���i|�rR��)�TxŪ�v�av�SǣXI�;(6�I|��a��+&;�w��j�>�p��uJ^)�Y�/6�g!nS�X M���F�kaJʑ$�Dạf"/��NT�YW�y�n�p�������"a��$���0�3�@Q�B
%U4�=t�-|�	l��NU������!t��v��I%u����@d�s���~�������R�7�)VJ�Z]�m�2-0���Лr�3+E�(u`R�a3�ٜ�_�%�)����	�U�P�ґ	z{i��_"Pɍ�$-�w���3ٖ�y��E��a��i$d���LBPi��W[r��%�:mW��{�A$]]�6�K%oT4�X0��;4=�=cCK�����*&P�����z�h$��d��r����b�G=����p�H���4RY+z���3��H����DKO�~�c=\�c]ܑB4�I����Hh��N�4K�%�{���b��I'�������FЧ�P=�)��C��@$K���[�������� ����A$��4�H�}��j��g؊�5;���!mSm�]N�y$�{l���U�������*O��)��ߙ�4�����_SpOy�(����?z�uǛh����UH�Qװ���:S4^k+W�R�����J�d���������.U��v5 e�MWb<h�l�߷�%�'�E���� ��b�fY�u�(�]����q�`vN��kG%p��k���h+,�����6b��
��U-Ս�taS[D�U��lk��̉Waf��c����%v�k2c�di,��C�s2�\�qT֥���ř
���.{d.�k��#���	�dԱҮ�j�V����C66k��B?q��(�Q$$bc���ЦA-���!$�I=�a��N\����^��D�.zy�sej"�bB&~QͰ�_%~2uE��۵T*�I�z6�	$�{��h����gM㙟d�M�#���NN�H�{��n�ק���_��I�?u�	 ������uݳ�x$�B=s�4�G������JC�6���J��&}��=��Gp/B�YUr#!%�q���BH�ws��H.�恟N\�ŕ�W}I���>��!)D���W���/�H%՛B����N(��I^��,���a�g���Q�8��?��=�|���.��M�n��sXQ����eS��]����ɠ���`M����+}��n�=G�:��A%�Uٴ(��I/���m-��^[�;}�;��2�H$����Qk;0ThD����D�?P��( !������%�{�IU�(���N�vʕ�%}���PU�o^#��8�wߴq��@mK������<g��7ι�i�8�����ɰ�^(�K�;=ڽ�c3A�!��v��ߎN-��}J��V$[�8�k�I"U_�a��	%��s��Q
�{�hnK�qĪp�DA��HB��9����oS ��@1o��;\Y5ǽo4�H$��xx4Q���b�Ԋ��I�D̥YZ�j��i8��;Pf���=�"o�t�ވ�$C]P�I$����ڣ����䏲��H�����+t�씛���)�����O����N��v{�+�$�Kj��%���u2�ZߙB�/BY�a�4RJ(I�]�M����
��r��%�1H$�^$Մ.�Y���2d%(�G�E����Kkv�-$J�ަZ_w�X��RԔV�r���a�Jk���I熄`�� ��T�{�ew�����b�\�)]�VP�i�]Y�)��S���	 ���v!��mP�������?AB&?�컦Z�$�Κa%�K�Gz�ȍҍΐ�����CQ+q�V�~~�{�߹���^��u/d�f�=���g�l%�y#�:���*݌*�`.��yת&�bǽG���D
J�������lm�ν���PIN~�L��l�$ ��f�0����wD��{�����i!�"\v{��R">�W�4X_$�
�9�_`v;�i%���a��I#��"fR�4�o�[�$�5��(���9P�}	%��θm$4D@��_� ��Vv0�O�9�9��h���gֶ�l�y�**<73M���#�9�y8a�E��Ͱv�!/䨠A�;��}J�(L��^S�X��I%�f��I$��w0�Q^�[��m��ǖ�iǻa�RQ�ɢKhz�L���%�_��{�g�!�#����}��>�+�ZI$�nu2�I$+�����~�\}
���gv=^� ��B0pA��1#��Ꮾ��D�^�m$��9�F�Yٙ�Ӛ_$���I?7�B���1�I*$��Lz��G�׫{=顒7�"o��$�B����K�K_t��sz�v�{�DR3:�����D�[��<���������
)37�X	��^�����&nS����Z��ˣ�P���dJO*]\d��y ���> C�ffg�_���θ�Hu�?Y2���6�=�͇�I$����-�F���U�����3���$K�]z�������[W�|��>)���!OɻS*��Uq��
�qu�a����3L��Kpa �1kM�}~@'��U.R�A�ɮI|�5״I$As�O�T�}2K���d�Oӽ�04���W�G�"T��Bg���N���J��-·Ȣs��_�"W՗�7�I$׽-��Tg3�	��6p`��l^H�O�J?D��Yw�Qa$�'�ĴIzL�dL��F���R� �UޱD���{�E���~��L�x�s��g{+wZ"ɜ'�V��a��7q��~	;}4g}�P���9i �l?�_���ߤ�� ����ˡ �ks���w���0�w�Dd�;N�4�� ��Q-%9�L����C}���~���m�k���V��:F��^�w��{�hm�n�D8i #��nbޣ
�v+��%����x�>�=��o�7��{�?A���a�9��ᙘ���G�l*�ktżZ�.M��M��0�E&]���1��2��]uX˵hA�#�vLTSF�6�K��&ɑe��n�1m���Nka�5j��f�˵��i��k�-�����<h6���`�E�VS@��B�Cfjl�r��f��z��nWd�k�4`��MlĲ)�2U�ɗd�f��v�� f�ff��i[0P�ǐP�mJ�5���۱�����M��T��M����r�t�-��oh�cM��O^�߈s�ȗ?~
+����%����\!����`$*���O�O���K��!��g�HP�1ʔ�cbW�]��È�1���{љZ�����_%�]��H%9�4XI%�qg��7Po5kgBGW� �*TL�3�y/)�KA$��l��DD|�	w�R������	$��݆+�gu2�_j�/$L���%�|���X|w���Uf]#�i$�{1�%%�4ZH$����Wjݓ�$�Uގi>��-��H�Jd{�V���%���t�׼�/�NL��L}љ��H$���ZH/�U�\_�g5{���㯆K�l�S]���&��dn�b�!)L+����"�e\B]
9�ؕq�}���T��؉ �3s�eۖJ	Gf�4����[	tb�����N'�h����ƚK�[	;�0�x{�G:e��K�������:�F6V����c��Yu��z����tj%������� �{=��UZ¿N�j�'V�e�L�Vd�uG%o���5���3��T*^�����|���f?�o�f�I/�_�$X���PH�ʵ���T{��sK�%�����Dn��W��"'	+w������4F�͜bx\�ǉϒQ�8�-$�s�m!#�� � ̘�Bg��^Sܻ���7t��/��p���e$��l?�	/�K�ϣk^A'�M�K�[b���Kٳ�?�@�d��T����KL+��4JK�=b\Wk���fg�Iy���H$�U��6�	%�ϡ�7u�2D��뿀7V[�ʰ�d�$$)���	w.*P57cqŚ^LXCjY@�*{��	p"!)���X�<����U��D������X�رn�ǝK�A$]���O��ߤ���	UL|�/e�%��7�kN�>Y7��^��I*��I$uwz>ml=U����X�V�{�3aO���(��a���/.�9d��f������U�KG�:�y隣�I��]�8��\�_�)Q�#�.�v�8^�8��_��9���؉�7�����>�]n�z��Nܝ|��� '�C��X�I_�~a��'���?�_	�����2��-��}����UO��UP��"W����I$��O5��y�LO��$us��W!d��>����qM"g:6��:�ma��%]ޡL�H��6�Jsc�0�;��T��k=~���ߒ�:�/4�f�#D5l��
chG�kN��@eX��L�k���>�¼�og����У��7�L/�U�I�����=��^��-��8{�PI$4�\?�A�Y!BXH�Jd@���t[D��ѣB9��#��y�%\f�I$���4�I|�<��*:�ny������0��&&~�S���{��	N�u8K��Nk�X-�h�|�I/Gg��iNtu'�HE{b
w�*aB�B���m���ރS��8�F�_�I�܊i ��l�D��ʺ��*��PO�[�8j�5/�����$/a�k�7�%&�Cۘ��Z�3��/m�/�� ��ޞ>�>ق昸�-�)|��>u������ ��p�0��O߂���a�&�E�@���Al(�G4I��C�~���M���;��Ǜ�K	*۞i�J
����Xg;9�Jͦ>gC\�e����uڈ0;et���7J��.ra��![���+j�����z�0�[�϶�w8�XJ��i�J���4�ӽ�o�<ff�>aLM�6�	 +.y�X=^1�`�&_D�¿g1D��y����ǤN�,�o��I$��u�A$u�K#�#�	�Kr(�F8����B��	�����=�7	$�J�6����4n��iں����q���*ܞi���U��6���0��&~�W���?n
��t�FS�~~�I)�G��H$�U��)��"�����]�~�k�����T�M%��C��R�z*#�
5�(��K�_1/;7�8.�P��D?�D�Yz�h�� �5�?�ϝ��;���Y��I�k��pw]䯱1~�ՓH�ײ�ė���;;����I�{_�X�ќ{ތ�ǰ�7Qy�x�P��xx]��T�F���r��=��1�{`Y�ƽ��?n��|=g� M{�S���^�.�m���jʔ����6��ߋ�ߔ��IX���!��d]\89�L��
(co+�c���S��_^����Y�P�[��rQ�מ����Q3�������[��?��NV/\�ĥqK-�1菽�<C��Q���/�	����Nx�.߻&��O!�<��]��J�P���!�K6ʻ	��i|��/t��g/m7���{�����~���Ow��k�$���΅�{l+��a{���U���_]Q��&W�嫢/��=s|_nxm����_B�^/]���@�4L�����]�P[�<o��VAWC��it�
(#M���{N�!{Gf���o�<�.��3݃+�I^�&o��6�bgQ������ ��t �^]�Y�gͼ����������O��\ζs�ߢ������2�^I��d���t����Q�r�ѓ�pBf�޻�g/��ܤ�Jg��=
�u5�}Ͻ|P7a�^o�|��-���Ҳ8���*D{�QNy�"��d�y^]I�}�I��rbl�.��w�<�=�s�_�uٰx�C���:��.�}�Ȏ/zvq�	��ף�|.(+\}IX���iX�V����Y=ӳɚt���a����%r������������O�����w�fj˜ه�x	����d�*!� ��%��ʘ6iu��5���B�lXIK�b���U,�:6�∣a[o��K׬�ZA4���q�u�S�UUD#��5"Qr�B�5D���B��*�&I2 ��9kl&3R�\�5J�G#&! [ώ�jP�(B����'c���䓢֒���Dc����!%��$�P��"5I���$���XD�T��m"B0�����9�V��DU�D�>B�GF�\"�ZAAN��aj��E��tKK(H�	�,��HB� �5�;��B���dE�QQZ�`�R�V�%�lM��b�G5Irલ����-�h9I��) AR0I$p"��qbHV��R�$�
�#�(����*T��v��H2.;mEPe�DUc[�D��rC��E!&;J�$\"H����u8@�o�[�*3J���uoq�V�8k�k�G����]*�h��C�jZ�.�5�Fz���2�Gev���cÂ$.[�G�c����osWh�d�1��:�{&��$�3D���C�.�buU&��!��K(@]5��8��+*M���lLVM��+�e�M34b������畵�Sd�T��yw�������p�;KrJ5��Dgh::k�䃣ܹ�%�lat]�
1e�Ռұ�ˬt��ʔŃR,Â�T�&�,.�6�	t�]v��{F�j��)��r͙�b��m�L�M�R4l�<h�])��Blh�l�k I�*�J���nKZ�׵,�1��-(KQa&H�^.�C��J�DU3��6�d�k���Ȧ��&��6��iN���١����flJZf�,e�F�9`KS�-if���P�-��T6r�Q�a�3A��3H��%�s.6J�.�M�{E�&9���F$mԋH1�$`-��l�A�ؙ*!�1�m#�H����qm2��&4�!�k�j��&Z���3�2&��,�Hݵí�bf7Եz�ɱ��01���̱��a\��Dn�q���5�[�,��W0�g^)h3)�t*����Pf�k��G*Pn2$��2�5�fz�E�v��`�,�XK&�\��!�팋Tj��i�q`�^5� -u�ۘ��G���!��H�S�Ď�b(����5�X�vYc�a@t��[5���TjXK����'�=�� wF嶎f9�l���֙f���5@`K�H��f���O5pѬ�K�j4v��X��f��%tW��(��WjS1kF-�,IxjmF�f*Q�"��ȤF06��`��n���l)Վ��E�m�x���䘬��V�8�R�Iu#���T�Q��i�;�1�%�%kp��Bf��eά{��wM��WHK.�Ѫ�@IkuK�kr=oi���L�����BRhkk�,�ѱF5��s.t#qt�2C#�)5�%��,�ܒ����%U�t�s�v������uZ0#+��=0�N��r��G�� �ͭ��M���l\�1fp�F1���!�[:��tb\�4��ѹ�*ֶ�Vp�u&�e!k3�:4��$ͰcE�֠<e�X���&uȸA�[�Rf˭��q�B�1+���\�nH\qE��]��j�5�R�61X
�f�l�H�y���m1�mJ�b�L-35�,RfThl�ծ"ZE!؍�-�5H���M5L��������&$�{�%���$&��A��	 ��v���Wػ،g�U�v�i��I*��(����7!d��S>��Ob��h%��څ�ݫq�GIW��Q??�D�/���Q��>g�˪��^+�%uxř�f%}}��D�퇪�I�.�F��d����]��$�J�5��D�ݗ��������,d�Fd{�G��O�f��ں�O+a1n��h���*a"W՛<����}s�~9����fD��a�Վ�R�`�&&~��)ׂ�y�[�I*܎��)���ɿT[I�l6_$�ݗɆ�	/�6y��OP�꜉b���_$��beA_DL��*%aqNKk�L�W]t�:��[��0��l�wχ�]gȝHҘ�[�1�K��{!��	 �gGRig�����ܟ=�Tߵ�%��Y��6���!��b$̘1�
=������{�hk����F�%G�<�'���:�0͗U9����d�����5Z��;���ۇ�s �<wy�7���>��?|����z���$_nK��	�_Vt�i���7�߷�;�sK�|l�
Ɂ�}��{ʉ`%YѴ�"PJB�Yʋf�3�<7�$I{��4IA�O4K ���s ����%���1�r���D@K���H�]��?�K䒭�a�D{^�:^�) ��i��ݒ��I���w`��z���$�f�a�?��-�:�*:�?�B"+�6��" $�{\�hd&YW����$�^��1LH�Z!���ف�	bm�tL�ځ��8L4L��/N�)$���eupKm�d��nF��	$�ns�5�⛽�zV��ɪ�O�xR%w���$�?y�~��<&]�I2d$���P���c��}i���I$��y��%��a��A(����N����5;�U<	���"TDE�6�BA$�W��0�"r4z���J�'��)�Vǒ=H�s��d�iڲ!�Ӱ�m�?�Q���n첿k�ލ���"/ޫ�o޳1�c��~|�UB!Eo>;{��g��z�t�W>���6���}pB�2`D��{�"���`�fp���Z�r��'R}��D����a�I/��}4�WX���_�a�^ny�_�|�RL�� /�Za[�a��I�k٭�i�����{T��6�$��;�a�I;�����D�?W�Tl!U��&"2�K��۪Uv.M\JU0��M���YVhY�v�1���)B�W}�
7�2�k��ä{�UٴI/�(���[	MhӠ�&{�q�B���m4�H�nТ��S$���b�M#��b�K!L,�W�*(���*�zk%$�{u��IB][���'#�/J�OE�Ģ�X�k2E|UR�V��Xi|��#u�餉�z�,�uC��`$�IW���I-����h���$�	CaF���uCw«c����J�]�	/�9]�D���tќ�n���vֲ*�-�q����1���9�Jϥ�ڸ{�ŬO����>WF����G��h�j��Ώ��~(�=^�+�̿���?"@F�^��}������˼|�L��&e�|�sߝ2W�N~٦�^`��ck%$+��m"Iʼ�$�9�L���G�f�K����u�����P�!
�Q�y��Yf�`�J4�җ5�e��}���i��P�����/=�i|�	���4&szh��G;6������b����Kܚ.��B�D���M݅��Ka"\H��Tԧ�͡�c�	 ��*��l$��wS$����O��c��K���{ݶ<���b�̒bg�2�o_���$�Κi/�_%��^V��x�L:}у|E"gדD��4p$�����Q -�)_�L~�n�w����k��/�Bs��i$�v�}ב�^�B� ��Q���[��Jf�ahJe	)Cj;�-��H��u�]��m�֡H^�f�I-ǒ�H$����$�H*��O���?��9��{w�T�Ӈc*�<�Ew�8h�EZ*��rf���C��Vޠ?K�{G�.�V��׳z�/q�lF�f��fᙁ���������YF���-��^uSP�Ի;PU-�J+,V��vQk��t.�a���m\U�BZ�b�x��lŘ����,�yg��l��tг�)C���$h�j�v�F��d�4m\�d�����E��Ԇ͠�6�M���x٫Mf�Y2�����\�)��l�v&
�C,7Mcs�RatM�B�`Y��a��ۊ�,����+�t��f��,#���E1���[�:�X;%�<�V�����
d�J?�&���M��Nn�4��"Uvs��]�dǧ������v��'�w���k���be薘V��a��U�t�uh��B�n�s�M$�H}=�L��	 ���m���Ԗ�/22\��yd$�D*(�߂��K%��UٴD���� iΟC�q�\I��_%���K3��2I��&"R�i^ùU_X�w94����}sW4�I%�K����#�+gyZ���^_,<B^�8	�JE�}F�J�+�Q�l0I$��y����]e����~,1L|��0�h���_*>�4�zk��t�~�
_�ᬶiH�(3^����AeCe.��2�нf����w���g���lM6J7���k`B)�v�m �	)��M��$�����*ꆒ$u�攉�|��2f%	�v�F�K�����{�Cf�.T�n�L��Csb�l��kVT����ojs�P����H����?�gg�)D\��t�G+�&D����G��3�h��|�Fa�9���O���b�%9�ݜN2d�O]~/�K���a�{=9���0.$��B�&�V�X��A)�a3�D/���&_]x�ɹ�lbH$���a�PI)�/�>
!F"`DB���p��Bٍ�`Y��$�J溃�S�:i��H��Z&�s9q�iWe�ڽ�bD̒TI(�?�W�m�J!��Ti���O�3��'�}B�H�>���TH{Κ[�y���͐W����1Q���G�j��MD��!�&�ql���Sk�lZʹwS�{t���)L��Nߘ4�IN\�M�HeoU?���}�Bbd��ː�W�mJ{��i
\K 䤦dH�J=���[a���T'Ǧ��n���DG�U��ZK���t�I%��ވ��_�ǃHX�W�d�Lġ3wiC���"FWm6�_%K2�>�*���0WM���Dĺ��`�����O��*bW��ק7q��?����X����k&kӓ/ fe��Y������G������G�| �������$����)$r�~t�B�@W(���>F�z����;���e%�^��`&�I������{�Cr�5g��:�I)�/�������1�x!��:&�Evmf�wiw^�.��%��O�C*������Πڗo{�F�i-�B��R��d�%�/:b�d-ȹ�%��%�;����-е5�ī�>�Z4L�%D�12�Wܕ�i��	��a�RI�s�-��{^�b��{k*��e$@��D��^�N`hE%3� ���m�������DHc�k�2RH��M$>I ��0�$����b��r��%Gە��4�
�%�I3dL�B}�:��$���ݡ�A$[+�n��S�H��;�%�Ck���Z{��H�w�"�3(L�����*��s�6��{)��K��yx�i/�_.�\U�����A���e͸���r����p�s��7^透y��F�7���+̓��W|1���ў�}׶C����q�)��.s��ŗx�����BH�z���^���zv���J32��KO�o�1D��K���Oa�X&���DD�M�	 �OݬH|��.�\_�z���H�d���25�Ȳ�t��[e1�U�f�Ќ	�A��7������q*�~��� ��Ja�|��|�����+䗲��a!q��}Q�lz4-��<z��0�I��4�n+&f	Q$D̓c��%�&�4�օ�wׄw:�>	$�w��a%�(��*��$���s�����)続K�"��C��))����Xi$NeO0A$�\�$�Q�y/VU��Of׾؂az�a��I}UŴ猢A�&bL�����=�x�Vzi��5�A��A$.긶��$m󡺼�N4m�RAow��ȁ9�X�PfL̡3���t�I�m�0�\]:�3K:���/�i��a$����-%�ݾtҌ8#����>���q�D�}�g�7f<˳+���)���l�Bfjs<(�
3}D��n�����F��[�"N,�~�~,,>���7]c��A"P[\�"����.;E�Q�*��0ƹ4*&�. ���t�m�����pVEa0�c-�� �Q2֘v�6X5�`.ٗiIY�.mҨ�fU:�omm�@%��K�A��F�"�������Ee,�h�͗���Q��36��4:Ř��i��W���٭����*	���m�.@�U�[V��jC���A+n�@җ`ֲ�5��Z�X��,� +2���P��\�h�)K�G���y�U�Qi=��E+w����B�'W��0�i|��,�a@p!$�;�ΘI{2Ĩ?_�>sy_1yS��'+Bj�$�BSs�#�ܐ��'2z��I#�S�P$7�͂@>s�{G&�W�=���Xrf`�DL�4�Ody�	7���A9�F��R���H��@�Cy��?���^Ԩ�4������̚�M�B� ��P������d��nN�΁jw��߈�l�%Y�H9$�I�2�ǵ�I}�m�zMߛ����O��5�&��i�O�{��|6i+�O����A!�sk��w1��qJ���#�[e`�-Ҕ���Д���3�`�PfL̡���k�5��L�A�{��9;��r��b�\C>$+o1�H���\ɉ��-�o��|ɊЅ%�y���'����y��b� ɦ>��^wߙ��m���v�z/n��_--�Ԩ�(8��G���s|���U���Nj��|?�����1��~$@�����I�߶�嘱������k�P��?	L;�k�$�=�m�إYwW���d�7�͂@$��l�갘� �bfIl��0���gZ2�;_s�S��j3m�H���ɱD�(��*'��&��D��D���S����>	�s���mI�p}�����${}��~���$��Sƌ8Y���~��򞡺��њ7HD��v��;V&�(�u���5�Xa���f&v�B��~[@�32�I=ʯ��$�6�d����+���{+8!��� �7�t�O��Dɘ�"[�TfA��v������A����l���-�� ��Mj��������OՔ< +�3"B�%�ow��A$v�Т	6<�z�j�eTF���>J*�'/'W�tw {���ں��7��O%�hn
g�n//e��^]��wR��x�	@W����;���{�c���������V������Γ<.�LY�P�5Ӿ���w���,�L:׮{�Ξ�8�1�v٠^�� �!��֯���4���;Y�[���<j�`^�k)�4��3|OQI`��0������1���麦�U<fߒQh+��)M��s`]t�� �(�r
͟	q�*��6��ٔ�I�������}~��w��N�7|�}qٓ�9tۆ�i�x��Y,�f�Jk����{����!��e�u��4L�[�4��?�;�NY�2O�U{리d�3�\���j�';��;;�O�HI���	�_x��z*�N��|9�٧ؽ�!k��F<�z��Б@����|��o�y0HF<}���gw���w�}����n���Y��v��L�-c7�F�#���gca����G�ԜW#�H[O����d//���^��Nyw�ѯ�__n8��4�9��n����z�6�'�*����	�υ��y^�8��cu��'�wa{���F����?�{��y���q z&��-����gM/����zt!ᎌ,1u�{�k���m�C�;��=kc���ڰ������������gF^�����}|�=���7�.�;g��T���I���W޾���w����v�'N2,^��%��|�@�w�lfQ��1�����W9ie�T�z�%ËK�z�ٻ���o�Σ�E�L�B�I��"H�1��$q�a$Č֡^�j�(�LcV2d�	�OGGnJ�.���m5��t���E�J��� �X"&�aE��ڭ�bbM�Z-�F��ŧN+�Fձ��6���͸vu�&ű����H+�#b��T!RA�B�)ã�:FF.)H95�E���
Ē`� �"��$Y�0Ua �$bAC�5QH�dpX�\���1kZ4�mƤ�b���c4h-��km�-j4j�mh��DV��X�LP&H喒0UL��U��
,T0��Qgd�%�"�eR1����cTb����ŭSj�6��AZ�v`�F�ŵA��5XӪ5[fv5iscb����X�1�����)�;c[j���j�Ed�V�g%DӴg����X�v��A���^1��m��XэLF�#�Yմb.DI#	�1��SZM��NأM�l[W��"M�>���.�}���m~�B�hp��!)��/��mg��satx��r��d�Fud�$�/;��'m^�B�1{�w�<���a1*AP$�̒�6�P3��L�E�ƏX']Sl�md�8
�l�2�d��N��1κ��,
S[iV�[�-!��Z�-b���i�7\�WIHB�����Q(h%%3�o	��I?N{��C6�J��7����7Ϧ�"_�#"f%DI0�}V	{��řz$��#^�~d�I���'�~���d�\ϒ��ܯvʮ�d����"d�J/��ٰO�o;h2A���������zc�� �wk$Q3��l��Ĉ��!}!������x2�z�t֊~��Q �g�u�~$]�{Sg���≛�˼`������q	�'��쁛��$]��0%��rΓX��.�MEF�!S��{�.K<~�N���χ ��_~���:$�����?	L{��~�`�+���:�_��ky�	={s@Hט� �]�l1�{���M�$L�S$�%P$V[J&���Y\�n�:�.�l�enQ#�����aL�;�d�D��dH��A���%{!(�����?~��cd����R���
鬦W�o�q�$�r״A?'��O��k{m�@�N�}�@����׳>��x�"p�11 ��k�� ��m�����aP���>���gٜ�$�k{m�I�}ba�*d���k�x�t,�u �
��L�~��6�'ⶺj,)<.S,�}�~l�`�Y�dH���6=]�~`�7kg=$�+rGd O��܆�^�l?�;��F�w��=�3�"��ʳf��S:O��a^ؿk���r����d�����\��/F+�Г�;�[���7*�[w��fa�d�W��߁��3�����ə�����T�p�M������a\Ŧ*�e���h�.W0���@���kh7&��A�p�ҁPŤ�K���`���������n�b�+@Ks�#(J��IY���]�l1���4�]Z*����f�j.��(:�,5%��K��ˑ�ZH������˶�&�iG8�J0+F]Ζ�n,�"�?q�o��jGFX���u��e¹I���5!���3Kaa��Y���,�v=��3�^�%1��;u���}�����)6��t�}�y�Hy���˄���b
�3��.��.+=�.8a�WS<Cݵ���V�ES~ɰ}=Z�W�^���!��Q(`%��`����$���� �a�.�����I �vy�A=�\����&D�)��l{c��T_�eU�gz��B@�y���݊�D����n'G�r��"��&{ٌ:G�E��"D��&_�/Ur����`�pdX�ڋ��sA?���$�خTA���e@��7�0�a��ύ<�����`A��""R���R�m�݁Z7ݭ�ʡ��n6)����������^�Ͽ=�P`���A �9��.9P���J��{1�A7�X��g���b?	L60e�͂L���3˙�Ĵ:I٩�e���θ�a,�W��S�*�~�XϾɗ�����p��F��^��������ʱt�V�^�F�l����|? ����|�����I�U��$'=��d�De��jǯ gזa13""��Ю� ���	'�짎H�$̉�=O$���Qs��L�3@�(��VβXWs��1�k�GĬ�J�]HB'�9����ݗ���#6r��g%�TH�t @�dH�����Wy���o�7�ݽ�)՝	}��(D�g6I���x��XYV|4$�#�"���DP����y&�K��n�y�\���k�JU��y����'�GwSo�ד~�+��~�޹���~�;�i%y��n#iW��L�ްЙ��\H���>�6�|�?U�N�f�|�����vS �k{m�@5Y*�ץu�R�i��`����d1V�$B�ݿ2	/�2����9�>y��k&���\�	�@��ڟ9d7��*��k{�_�f>��i!{�{W���g�CG�*�)]��|>������~��gov�ĂA���Ln�LLL(�ba�=*��UtΚ��/��� �	۶� �خY=�b�So0��/͂@�R/Y�Rt�L�xέ�I�WP�][���:ώ��};t9�\���13�g�y}��:ԶnM+�X�c�͔]3��5n�ڹ��:�(���D��0&e)'�+���Oğ<�l�	Ί�6C�t�����}��]a$y�[d}z��B$�"a����F揬>�r�o}u�I'���$���O�z1��G��O�}5��n�~���lH���W�-�^o�d��Ψ�@�}���!��zv׼��� ��[NuO�����&I*b��;��`w�����y��?^T�A��sጺ�f7�ӊ ]���7�/�~��	{9�����Mn6��q7�iYh���z�G�lӁ~+جM�T��|���.���~��_��A|]n�o?�%J��fa늴I5�����.o/ee;���I��T�H'��w6y^{}��*Г1*D�$in�R�6g\3U���p�0WF�e�iX�4�P��w����@��	Ffb��\�$�TuH��w7�^Ӌ�Y����c��}�:X/����ȑ3%J-����I��͘~���c��m��g��#�ww�;9�=w��H��fDʍ�h�j�v�$�s��tx%[��~Ω�_����L�y"D�̒����|S��u��9>PTeϺ ���kv��$�g�n;ENo�v `߉�s�ƍ{�&��N�(�)�������=�lW�Y�P����ą5>4A�w7X`��������%g<�ڹ�Y���̀�t��n��t��^���y�l45�> ^s�����K�No�k؈,�Ǖ��~�G��V��Fzj�^K��q�P�B#�� U���
h�n��s6���qt^I{ר��,\i���Pg2�aED��
"�؍
BgklA�``Hi���Æ�\�idفnmY�,�*�b2��Z��`k]���7�R(\�6bgE���2�s1�D��tkmI��GW`�sw^�<R�Ѝ
�J��U4���ī�@�ub`�1���;P�9ʘ����%ķKl]K4ME.�(l�X)[A�3-��G
���,Ub�[[�͗@.L5Y����ߩ���S����C�~"}����U��L��T������*x�F���L�3������`>�����=�ֺ��8cbO� ���0A3����a���^UD���o}H��2T��S[��O��cݶ�g�/�z�?�zj�p�H�y��A1��O��z�""A�f�1���'���~���$O���l�~ͩ⳽�8f�?U�c`�5�F��3$��[��?�uF�I���6�z������$�������<k�w�1��˄���R~���M�^�;u��Z�d&@�Y�����0�^�Z�6���=._	�
S���0� ��������gIŉ��A�z���6I&={�����IzLʈ�fa�c��lz�n�J��o�H��C��ڊ�W��S���o�-�l���ց�W�����������L��n������#�5Dב���^�N��!19RIi���
/��~ �r5�~$�~���d�O��_�C=V��OueO0H�z�J_@�ff(����7u?Þ{��}�t�N��� ���$��r;�4d��*Qfgz�E�H]rŃ���7�%�I7�ڢ+}�U[G�{�{�/��3}���"$�&a�t����I���x҂֝^�~o����ӓ_]��d�^�Ȅ d"tI?4	z�r9�қF�ظ%��JD�Pp�։)�XV`���1Q�޴a�3
�g����0~έ�([���1�ܓk����
�kC��}��D��55�1J��0��g�F���P���q���{g&���o6 ��{�*nm��a�c�eD@�0�`��uD�W{�$�g'}ܮ��9�US�+�t?,�(��z�tV�7׷o����k��lor&9@����ἼJ�G���[cp��8 8-9�3���H9ӳD�[��`��9�\!5�
Ffb�\����7���{E7=�(�Mn�S�I�糴w�A��DN��b)��>̕(��W�6 Ϲ�y��[���ǷĂ�t��]��� �g��pTF���p+���(BS
fUb3�,դ��%݆��l�F�� �n+Js�U���A ̉3���A&�;k�?Ws�ą׈/��A�gM|I5٘�Ď]h�9"&$�g��`2g��g�#���
�T������`���{jgs���V�&:��78	dj���0�IL{���6	,��� ���9�wR���g�$�^��	���df�c�eD@�0�dG[Nƚ�[���I$���`����\#��O\���q&��F��g�j�̺����j�FIߓ�������t���j�/޸{ޑ��ύ��ju-�������>}ߩ�O²�Y�TD
Ffb�_�[d�+�
��z���������k/�� �mt�)?��ꜘ<�i$�T��).�����Wa��{hm��m��豳,�c�]�߿F�&fJ������$�^��g�@$�鯌vʩ����{:��$��y��\��'�m]�]�=y�_1��x���x����`�I���?�$�[]����/&6�7}q�>UX��NyG"DDăL���� =[@I$�A��&�������Pd��诹 ��Ox�B�1$�=��z�� ��>�^7[�7kt��o�A?�뢈#�ξu�o�MR�v/�O��610� L��E�����{���c�x�&�/i��"��?-udP$;��Y
Uo�t�QNg�2L�/O&f�Ø��? E@�)d?﷞N�6p�2��#��'�o@/U�/W�
�o�`{w��l�^��e����ܸ�#�P�����c@z*��������w�x"�F��sfyNԞ�0���]w�h_Z������>�c�ĠL<S]C�7��'�s�$~6�֨�/����q����9i����AgkI��t�WJ@͑^F}H콁�M	�˨Y(EMӿMH��|��n����[3����J{�O/l�}tnu݈��s�3b���9�|��aѽ"Y}�v.Ziv4F^E\�9�E��/�`d1�;�3�������.���/{�'=�Lvl�@��k�5��^������}�c��4����/�
�!n�,C/��l\o1G�fs(;�x�{+��\�ÊZ��=����sY{��v��uN��1�"&��A����w�^X{.�.�t��Ey�{7��4D�yճ�x_.w=���	��E���»�v���so�v�^�8ng7�j`׾S�w�w.�����~s� ��^�g�o����lC�s��<��"��3�|ξ{��8�i����8P�@~����ȡ7�Vn�P���7(�.D]��fJy��.f����>��x�����FO�ѻ�O�Lgy(��a:1b��q=�{�;��|�Y�1�2f�'�Ӻ��;��S_Y�$Oq�22�ƾo-�~j�FX�Y������d�u+�_94v���oV�u�Y��..����;�����:�&��BIad]6�BYafq�И�T���$J4��0lX4X��V�'R+�$,��YI�!gN#QC��g����:�3Q���cj���QX�kD[Abf�+Wqfu�Έ*8�Cӵ�E�V��,E�B(*
�������kZ6؈�6����fiSN:�ED���&@\�. �X$R@TX��.28��i�5M��Z��5��mA��N�
�45i6ڂ�i�U�e�j�b�BEF�TX��6ҋ	���ѣmE���#Y�""�|�#FbK��E��#F��������Mb�֋b�lmcY�8
��1�i6��51QkDm��ѭS�X�4S�c7k,\l��b�* �k0��ApDqFM����@c"���H��EEs\�E��VHm�c ̐������ȓ�i4`�M�QG�pS����&�*6Ū�֤�Zj5�:-�vb2Z4�v�Dqm5�Y���m���lf�1�F��""�`�ɋ�L".AF��h�V��SF::<$-�\L�Th˜Q2��.ն�����?�<��:��Q�!e3�*�4�g\�'T,�	�mGW6ݝ)���p7d��n��1Ī������-��շ�$� ذ����c�ˠ����Z�$��,؁�e�Ʈ�A�%�6�9I2�b�`h��|<E�[h`m6!���(`Ը���@Ζ\ GK����֔u����R�S[�봱
�i�H��j�C��&�G8%�a�����#�����n� ����TzYpa�p�],���y��"�lP`�bو�c\	�v��9�Nf�^�u�#fF�.#i���eI����mf��s�sb%U�Z��K)��`M��H���U�<U�l�qJ@J!�v�!2]�unN!�35��*�L"�x��l*�<�V�6��ۅn�53eřIw&)�E�	�446�tMcs���\�.��[�d�s�] gS��"[�&�vB�J�84ao`�k�Z�Il�i�H0���C!`if��D&���%��phfd�[G+v��1���feps5�P��&���m�xj�5H��kMfM�
Yv��v�A�+�gF	-��Q��F*�fY�YcˆY��Ks�B6\�������6V�+�i.�z���jZ��M{Lli�%0u��1ʒ]�aj.�S�Q����\���ml��d���:�#c��*vku�n֍����p��H�-Sc�D�@�9��e��m��v�2�Ck2,
蝳���$��m6fIm ���A�cH�.��M���fi\�:�e��M��m��	eKq�t&�o<���4���E��ZS9lVj�T8MH� �W��H<k��,����h�vș�E�������Z��ڍ�b
��\hG��,4�P\���.�M��q�sA��#,\�4uB�-֒�6��dI���`vpJjJ8n��c4�\@tyh\im��0��W�e��e�v�4#��6��
J"ŷ0�5�7n�g�< X��k6q5��F]�\�jͰ�@P�9�4i5cP��^ Ց���p��\ �ۭ����� 1�kl2��P�:��H�JP�n���b��Ƌc3F�v�.�i�!H�E�m���Z�|�aY�ñ�:�n�̫��C��jl麇bb�Yh!��UЍ�\2�J��r�;u�;4�oF�V�CV���+l�
�tE��8E�q�����e�/+a%�%���E��F:� e;så�u�?��O	=*��0�U~_��&�Xq�I$@����~�ٿ!�Wg��M���:�(!J32TL���I���z������� ���Mg_6H6���B��"$�/#���f~���:}]_I ��n�$KP�B�^�ݯ<Hǫb���󣩂DOyF�`��
>�l������kٟq��4M{ݔ$�v��3|��/$R�诉�l�^@��"#�Jc����H�o_�n<����Oz�5���'�Mom�����u/ʫν����6��%Zu륶WZ�G@�,5b�crm�pk��F�lk{���_M��n��?|����P�ko6�[�m��=P{�'esBK�$�+���5�����TD�3*�]��5�ɂ��o��tZ�.�V<no����|�S���Ϲa��?���c���l���W����Khn��(�"�}���E�1y^Oޘp����$�H'���l�[�o��l�I�zov�����G;��0!8���$��m�I/p7�1&"GW\U�|I4���A ��lК<�����3?Lǽ��츽�"�}/G|j�a'��lAͮ��O�	��1�<W[d����#J0fB��}�?�$��ڦJ��5�^�@��_0�?��a�O�6�ho�[�FC�'nb��n�Sg��:�s���6���� 	*e!0iL�\f"ʀ:��1�%}	Lof_y�I?�����$����4�%9��뤒�^b��� >3w��g;M�L(�"flWTA��;+|�{��<�f�ւI&}���O��s���2=-��G>�z�"nt��a��2*L§�]������P�I�8�j9&�w�)����Z�b��ͬ"x`7�g��t9��y���$�Xo��_!�7y{����xn��ާ(�~x(��$�g/2����h~��$dLɁ
�����ݯD�=�[�)݀I]�o�~'�I��4	��y��y�5(�L��D�W��MF����3?LǇ�?w�L��״b�<���;�S$x$�s�$���sd��m��~z��g�|������-.�cd�ki��-�(Bn�YXU1�ԍ��<5��E���۾݆�Q�������q�O7�6w��T�gw#�����?��x��$�DdH��R�l^_y�@>D{ԢM{�s�H�|�"�w6Fv�Թ�>l2�g�"��)X�O:�$�^���$@E���پ�W5מ�d�<�Q$�y����9t7�1,��&aS ��gTO�FM���H0e�I�Oՙ������"{y_)��?^O�ˉa)
�+ɬ�,���O��]MM,Ӆ����nמ�z�v����a9������sQ������w�P�5?q#��-�E�h�"eJP��3�['�'ݶ�vz� ]�6��>���s`�L�e�����z
V�jҦSEJ�m4�v�q�Fb�MvJKyjظ���F-qB��S��I�11&#����"�7i�I ���m���C�X��ŏ"� �˾l�o��0%3"#�f�o�����2���uo�u��"�w��O���?�'-����޽�ذz�:"2d�})LS���Lvo��𘈲
��ryi ��m2A ����f�0ĩ��0&%/g�yKt;6���xi���HiovS�H&/�͓��U��닌�>�Q�^l�&�?LK"�EI�T�+}V�d⮯�Xu_N_���;��'�~3��l���:#�ޯO'^���͜�?=/��cY�{!��ʹ�j�۾�W�2�_ ��u"�N�~�^{���&��W�y�fp��˶=zL#4�X0e����d7����.ml�sjh��y/���:���&-�	-"�BJ����u��e�L�h�\Ѭ�h�-"B�
K��+kytin�����rD��wa�e4��K��5��\+,M22��+C�Xh@�&��P�Qf��+�SQ�kHˆh(h�Rd �jL�H���u�]��Y�����^P�E̺������Q��=c�S�y�ft�%)��(�F�f��X�\1�Z�G6h36�͔Z�b��|�Y�JR&T��}Y_~��w�g���|����9A�͙�kgs��'��6�&$�6wʺ�F��}oqߺ�$�L��͏�9�\��t|1��uǪ�&���\�RT1L����O�9V�Ik�Y�c<<}n�bk0	3��P`��q�FP#~bL��D�O����'u�+=~�g4�g����ZD
�k����|�	�����|Ȼ�P��S`LM�ۇAI���L�����Vu���sQ�	��o�q3s�3��L{��`�cma���D��l�n�����UB�����[�l��.=���ܼ�}<�#
���l�~9�H�@$�_6r.J��{���� ]��u�ha)H�R�*z���m�A̼���#R��,�_uƞz�Nl�U����L�${Fn�rnE�NdϱT��y��T9�h@�\��7`�Y>n~����<?��f��A� ��?g�_�� �Mi�U����{\���B��`D̘�sp�m��x|q��O���HB:r��Gt{���G�{��$�;�&$��a�m��}��/Α>����=룵��/���v�C��27��oU��Og�h����E����&S`;��`��7�>�9�W��8�D�s�	�ٌ?� �������ʪ�|��������I��Qչ��[�����JлhR���5�lp=ek�������ҟ&nWTL]�Nc�D<ͦ~{��`��?b��������nP��J3"�M
�0�s���}�g��mX�T��O��E��o�~$���`��9����(@�n�Ǟ E&��)B���6H$��0��sgV�wGL�
&��	�Cǝ�+-@Znrl!I���[�d^!~�>QCX�W{����#5^CO�����7����?Ua�;��-�s�H/�}O�ބ�H������w�*PDV0I����$��͂A?����Tq��;_c&�D�
SP�0�������A=�*p��*�EiN𑞯s	/o=A���ޚO�Vox�(\������2 ֛��"��nв����+��܋5�/l�O�J*O�7��)�L��y�l�H/s|À�����Lc���v�dt�}��͒H/s}Lfu�b&�D�3SdO��� ��w~�z�X$���o��N���+Էc"Ɍ�9����Q���Q�T��U�l$ڞ�(�Ot�يȱ>�z�W��$����'㓽5�#��4N
D�2��o�{żF��޸���S��H�ܚ��O����Ȇ�S�R��ؿlB��bj�G��'�����Y;�ہ)�ˀ��1��\k��ņl;������og�$g����,�b�6.�c���P0J#)/T��>��{�﹜n�wa?k�n���C�I�n��w/D�y�H5�� ��}4	�����f6��n��`�Bs�K/V��GVZ��յ)m{S[��)���4%^%���ʈ�!D�̉&$$�	B�q������?�8����U��/s�z����rw��?F�#"�I����|�*"�ϫwn�V�fO�9�@�H��͂Ax��DL���j�[#l��Z�LB���FDI����s@�y�m0N��+h�F�V'^�8��/4p�M��$���;�h�*~u*�¦
�U��*X�����+�,w�-~�$��d�H/��u]�,�;��z��?6p�'	�"eQ�7͒~��r�K��;y��
ǒ+�C{��$=��pbs�k���n��2�"�7 ԫ�-��*'j���~��lթ����o���Vqz�؊d�F����s�Ͳ-ɼ%����HRO�eA�GUSf�z�&�]�p6j3uT���ы�m)�b�����dՔ���K������t�WZ�U�̠iuKf�6e�P�M��[�3��հ�K��1��1��%]�^�m�\��H�*���u"������%�Fl%ljA\W��\l����bd6�4�(iV�)-W6iaæ��-�����V�2
�� �!w6c��k]Wp�8��d]lb,cb,݀r:$�)���^ɩ�6�a��%&$Do�H�W���$�k��NBj��ԍ��GR� ��H�!*�v6H�ܹ�T���(A�o�m����$z��y�=lL����Т���`�Mww�)&�����ά��'�yы�T}&b����$���S �z+v$X�;�]W\�<�+� �wy��l�1
f&`�%�����^�<�N��!�=��?	��lXK�3_L{�����巂��\�>��;�q �߷�Ǎ����|�$�]U(f��������7���}�p�%�W������M;�R�D֒A�O	0�-o(˩.�¤Ơ�]M��=s��v�	�@`�R���/��t�R&Q����z�?W�|� Iή����Z�g}/>}=��H3��6@�/D�(1"!��z�ÍB�\�d/q�ItϘ���7�k����v�Ɂ9�,x'�BO[��7�M�vI��<����2��4�|O߬L�J��M��7n�y}���7�D�g��	9������p�����TE__�1"��q �	L!0 �{��7�0Hέ�(k3l�3�N�������gu�	'n�h�è�1"L��R���9c�{u�����ğd��O��#���$���t����޾�G�oWY��bT�"$�|D�I5{�L��[���h�-=��r�t�C�����Ï^������즷X��;q+�����	c�b-�ɻ0V��s(K�+�ٝ__}z�,�y���O<��{��d�Q ���9��%���{���M�t�'�=h�t�R&B��}U��$�{y�ѯ�p����h�?k���4+.�՜rj|;TT���j��2����;�u�H<�v�?o�}ԵlB�L����(�#�_�Ԋ��9�gw�({���0�Q��>w��|���3���sa�7}ތO ��D�pV5H�\˩���{s�/��^���3�Q�s�t�)~��f9�i��{�\gfC�v���{pK\ᷦ罖��_{|Z�|J݃x��{wG6꾜�^
}�qﹲ5M��P��E�*a��&h^��~����'�����%(�L�[�f���`���x�QI
z@�?���zd��)se�t��>�R�ޓ��I��*Eo�����s�y�P���;����㯻yN��6Ŋ���}|��zx0A�ޤ���Ǒ՚�̇'��7�l/���X3��|R�v^;�ԫ'�x�?!�va�����ϲ�n�z�v�NE'��6g��"o�Q�Ӽn?w��J����{9��Q=�y _�`����^��N�Ɍ��!�r򍒚6�©�L�ڟ��;B�1=JzV'mo�o��[�>Ö���`�p�)�����(�d0�~�3ss���S���}a�%xl{�+�8��'�]�f�њ/��n9U��ug3\8��L�;�C+2W�3��(�x��=��nKt(D�c22n1��f��S��/�/5�w�Rgj�&�=^��{�x�k���I�V�6i�9ޗF�w���ݞ��!��㏼��o���.vk1���{��Yݧ�N_��c{����c����˲�%3NFa72H�!�yI��Ng9��{��M:����cػ�x���{�n��>�9/N��*��r�3!�Am�!d�o����¾gG���ӳ6o�7R~�<y�f.��Q|���Έx������813���X�S�D�PU�5V�Z"
."�A�Q���ь��1�lriHSN���z��kgl\�X��VΘAc$�dX�I H2+#���1E�j�h��)�1��T₪���65Fnָv3k�4l�*	�i��QHB�p�k҉�X�9 �A�K#��dJ�Qd�fD��"��
"�*�@PRc#1����U*"1����MRi�m��L��L �	r��V*1"#6b�X���b�m����-����X3لEU[1�D�
�dLQȐ\YT��h�h��L�UT��c0aTXH"���F*HȖ��9�""6�Dբ�#cE��:1��m�[�f�J��+N��3LDh�EX�
����"'g�[-��[b�����6��hkS\�bk��q�A;k"�5�TADDQkE1�������j��E�*�j�MbtF�Dͧ��UEW��U��S����b�p��N���\��;����I���K���HJa	�a������U��o y\���d�~��$�g�}8UYݤ��˨߰�gM|H��(��$f~��c���?��0��O]�l�y�@.��AﱲI{���7���=������̨Ͷ����@eaCMJMR��!�զ�H٢�S (�cO���G��W5�4��3��~�osi�H$D�o���ݻ��į�{4	_���G�f�*T�>O6���W����K��e�� `�ݍ�t���k�����kf���4	���1"d$b<��M{��̒\�l���d흘�p���;�lL�o�1/�ى� ȉ�����P�&��0�A')����I���`H��ќ��<j6��Έ7��.�)�N��ˠ�������y}��m��1xx�7>���:c�B�c��5�t
����H˾��.mĂ��D��1L�oz�ă��lD�}��}�4L�]��H�gw=A�kk���^X�Q}��g[!����܉�l����&�P��ګe�0CT�eV1a5��4�텿�=���*0��[���~�6Iپa�~"��E�(�CC�E=+'ծ��������/�aL���dD��2z�	e�uƸᎣ�_x�[��l�tP �a�ݱ��w��*f�D�DP<��2�q��"g��{�~��T}b�K�~1ݖ��mmtW����1"$�"ڮ��4ZQKպ�x�Xd���ѯ"�'���<���xk��=ޟ ��~�́l�Ӹ5i[�x�����y�����nlJȝ�=>��$��mlP$�۾lW\�(�׳%������-{u�:�'!�����z[���=��ŭ�w�� �=�G0f>��h�F�͚O��(`����g<K����(������6���,#�m���b�[f��@%؆�.
h�z,A�X��K�Xbm�3�װ�j;;L73\rك:\֑�+����s[F�H�'0���&�.�~د�TYf�f]s5�
/)f�VYGG���r,."h�S7��i���F��
�*�2��H��j�&��-���J�m�Z�l��lV� v%tR��"�̻�.(�:ј�n�����~#<��a�
�h�#+�Y�e5	�N�rjni�D؎q�߿�>�(ɏ�>����o�$��khH ��w͟V�s*�dvh1�Z� 9mtW��j+=L�!O�a`��Ӿa��W�N�}��~$<��(�w��"2�u\GU[���)�
f$B0'�"w*�Nf_S�O����b:�����쬟�f��`���10D��&�"�+�Yҽ�L������?5{$���o�	}�k���s��"~kި���1"$!@luK��$�v���Do�b����n�k#-
���l�A}�u�9LO�w~<$�tZ�Էk]	PG$�
�wfZ0�Z q��X���k��B��S��j��
bTH��߾;i�Ђ�{L� ����=2=��\u���@PڠA~���5\�$�d��D�c�u����obJ�#�f�^=����sf���1�g�W�� �����zN�x1���,;��lL�{�)2ff^aƏFBW[U����S�7�Cܽa�^�[�'�3u5W��|	�I_�L�&�&u۾a�_n�`��[�;5�m����6	�����^����f`8.�55�=��u�u=�q!L�|�e:��>�n��r��|�MQ����u��+;i10D�MU���cj��H8kz�}շ#y9ׯP&:k͒C�ܠ�:k:+��u9U|��c�_,����$\գ�&�lw�J��,�0�r��Q� &�[M�(;������B��

bG%U���۞d�x��P/+���3��/D�؊�����s�}	Y��	L��_*ް(Ɍ�7�[C��_^�`I�ޚ�{��{{��H���A�FL}1�L7���d�ݡG�AcNR9���>����cc�/�L�V�Ȫ8���L(��e��+�B�3h;��9�!�FS ���f%ʫS�F�}�0qD�)㬉�c��N�q kݹA�	3��@�b�Rܓ
`(J~�+��^���m�MP1�	��k�L��h��$���c��� �w����>��RI�"	l�s���Y���"��V�β�{�t�I �_M A��w6�X�7�l*(�3	�"�es�fP^���G��4�̣v]p#�]�_>�>��!;@�DW|Vz���"/6���/s`�z��V^�{=��~�m�I���\'�a` �HBح�͑y��Bx&�����'�Lm��$�Z����6��)�6�$�q�a��A�`%"DM?���4H9��A�H1է�k�f;@Wyu�~�k�ˮw2!I2c�$D�37���`��R�' ����U�yL�O>�\��4�j�ק��Y�]�br����2�p�Uj����6�</�3Q�%��Ɂ7��M\%��Z'a�e�E��H��z�EN�WrJ	O�eh���]a?<�o���3�wH��M	-�d�Oǟv7[��ܱw�dG�I�}|OwBY�(�f��2n�el��+Q#Ch����eR[h�0Qq�{����W\h��8z�E|}���$	�_v17�<�K#n*�ͣM����o;`�;ܑ���>����*ϣ��������~$��<l�~:������^s�Y��M�v�t
���?=���A?}�� ����>��Q�l��I�<l�_v6�M��@���D��gq���`y8�3��$�wO�~#�{)�avtR��3N�LV�����K}��	I2c�$DƏ{�Y=�� x%�۱ә�=5A����J�w����>;[���HD�Ί��>'�t����UQ��
BƖ�Īx���qt��F��u^���u���'ӳP��F���J�=j��Zl��-��q�wz\s�z=*#�-r�Z��M�����L@���0��S��L�/l�Ё��ډ�n!6F5D�њV�bgCM\�$��L�M� Dz!���6��7V.��4�R�[W*;Ku��;hw[��Qn�R��bӕ%�DY�BSp�f�L�k�7<��Uq��-e�c5�#��c#x������B�*V�@e]ex"[S\�1�6�Q͕1�I�K��0�Ih�Kؚl�f��ۆ�
l͆!Lް����))Tͫ�`���2����26�q�A B��}����l���ס�_��6�1�~�7����fB��><ꄐ�F�x�s���(�9�c`�=�PD����DxR��9u�D̈��h)��gcլ2	�T�{�V���z��ǻ�$��y�����D��;0�*dT"�V�p�}�Bw����
�����I"oEc�9�0|D�G�S`2"h.��JD�"%��W�A?�{L��S�{��;���9^�lI��(	�>l�F�j�:/nh�`�aR]E*��Y��mIi^6��^	L&�5�ue4i�eLD���̙	I"c�$��p3��a��nМ�Iپ�&evy{��C�a��"�`T��쀦TT�&Sc��`�#�e�uy�����ڭ����WS��@kN�4[^���|_���9�G �������O4��p��*b�vb+"�<fL�1��9߾���"������ 烲Cد���*�.��9��R
�fb	�]T����,b"v,�t3�ݤ�o���ߵ�0K��J"dD�sBf�S�ձ�H�Á|l��Xh�` ��x��OĞ�v-��s�C���9�|Nɼd�̄J�[��6	����݌8y��p-��H��ȠI/5�d�~=���Gj�@oQؙP`�D��FP�a��q�:ю��Uq\��i�l�Y2j?=C>+$��B����(I ����$�;�����3]	�ܘC�W=O���t�o��%����~o��`^����zLN��A9|�	�wcQ���툱��g��>&�i�?I��w]a$��n6A'�4��R�JKf��Q>�����Ǽ=O#�å-g�ѫ����?m����]p��{c�ؐ���%ȋ�Ȼ��'��=\����������w��ټ��0��fb	cǽ7v���j�/�A�n��O�o�r�$�s�C��U{h&��z�(��a�	��L�z��V������w`�M�2=��o��"�R�˸��:h>�C�x�$�+PL2����Z�;UˇٱYMˠ0���K�eQ@Tlq��{���ss�]O�g��ǭ����l�":3��gN]�n|�w��;۸��&�ߊ�$�H2"[��Yʾ3�"K�$]�t��	${ݘ� �9ɒV�����E�gY"�9zQR���10������A?`S�6��M.��²W9�a�ט�`��tg!M^bT*~�*�o����G�0�
n��Ğ�څ�|���6Ve�B=�me�{c�f��,��&�No��P��t�|Rn{<���)�wl=s�}����l~��r�zm������a��Z��T��" O��� �{����Ϝ�2MQ��L�?w���&<�|A�޾o�u��ވ�uq�ne�dƥ5e��2�p����ѱ8���s-�m�%�Z�:�j����%-����6���ʾ����$��7�9)+��*}����`��vN�='j�D	1$��4�[��1����>�:�Ui$�ӆ� ����'�qs~���O�]�~��
�=���dD�c}h����`������Kk�1�4H$|��0�������S�W��6o}��5�	9�AH$;{��I<��'������.�Q9�4B�5z�P �&UX���s��*��M�s�h�H�V�`���v0�}��ה;;�Y
rUe�8< �ˇkޑ��ܲ�����;"�<����C:[7Ov	P�-/
}7��:�4*]�����E��{ǽ�`�!���zE����m%�N�.9v�b�3΍wz[�޳,כjkV
���ͅ�������{�ދ��ش�=�oH{���:vC�w����\�5��Kr�l����$��5����;ܷ��l|O�[�B":�}��H�|�\%�k���K���ټ�<ُd�޵�{�=.��u�Y�h���0����o�y{������zh�5�����f�^�b�`�����f��D7l������Z��n����G@@)��׏C�8dᡞr�L��}�ʋ�1�3������c��vvkg�7�����ul�gqoA^x-�:���9�t�{|�(~��Y�d�߽h뉟R�ޕۮ����[s654���~j1�ѐ_ܡ0K`{4-�}�9���ЭNyFZ��}�4z��zu���w}vѨkZ
���@��ڟ�t��$�����ݩ��@9��@sx��A�On��Y�i�s[���)t��uǽî�`i�ҟ���ae�ndW %ü}�{����e��~z}�E������ze�c��{.�=�۠��9��;�i���_��7܁C�/z�`���a��n�������Y�ŦOvm���W�k/�_u��G��Y���#X���̾�Eo��B	��^��k�A3r�Z���>W܋ў����+}�v���>��|ǃ+8�i͝[4��y��#5���;�j��а&~뀇Xq���|2����m�![��"<�������g�q���f�Qge�16Ѵ�Q\m4�	J~;?��p�I �pd�Bj�4j���F��[b�ji,X���٣F��m�ki��M$AI�E�Q��N͵L�'��QEZH��"0dR`�"8�aD�8p���c��p�(�d�Z�c6؊���cĕ�t��)�56�5�
�m���)֫X-��M���pn8t�K�c�dDX�J�E��VE\4�kQ1A;m��DQ�����2�4MX�E�1QDTB�؊�1�*9#!F��E�mn-2�CUq)���Z3LEұ�1+��I�6A�'��`(�PZذV�����M1Q��&��Z�`�4�SDX�&�8���6Ɇv0UT[j�l�D�
(��F2-�qG���q����������,�$���@j�(�d���*���9qT�,�<��BǙ���P��� \�r�]�V��L\�՗p��!��b��������U�D��/[)��AC �=P[����T�r��ka�˙utE�tDS�M��be\\뇈Ӗ)Ď� Jf�.��i�S&yuR����a5iE)΍V�HV`���ab�۴k�6֑�K/cam��f����dL`��v%p��J�/\�:�]�d��c�7\��I�&.��t&�*��jmu��d�J0,ʬ`Ҷ�Y�X�a�YI�γLFlYt�j�hۢ��Wi���	��-Ɍ�h�A�X�1b�1n�k��M���Z�*�"XG9���QՎ�ibTȍu�-SR/:i���-+�i��XU�:�˭)v���;Fj[$�-���K4�V�f��� �	�{8Җb"M.��6�]�:�`���ҹe���A���M��5��e����%��u�Dd���,!%
�۱#�d�#����g1Չ�*�������+��(gJn��ܙuQG- lZ*,���9 �1M��Q��d�b)V�F�b8�e��ᆭ-�c�-���^"�m�	��Da�뺆J�9m�����Z*Y�U�4n�L�@����u-�*B�8�2�����G0�5�vBpAhi+�KB1�*v���\��H���l���E�^ewTɥTC2�`.���\6'.�����l�F@�4�v�V�ML	L��e�r�#)6a���� ���&Ԭ�q*�[ؖ�:Q�;4/)#0F]�Ki�M4-D�۪&e�aln+�q!����5�x��c1�D��s+c��Ԋ���n��V,	�Jj�J�-���&��:��T�b1�K(K�4r���LB1&�����jk��^ɥ֣ln��-�p��kR��X8�����2뵼s�r��F.H.f��]ka�sƄ17k�b0ScZŲ�����K�T�A]�t,"���-�"�L˱`��%�U�J��EѦf*�lavb�ƪl��Z+42�:�hZ��f,�0���ٮ�Ұ�V�z��V͈"+����,֩f��n�Mj9������pe]sY��M�����+5�Jb��vƮ�0�IJ�̥�I�&6�	���&�P�]�A\j�u�`ʫi���4*�IM45�M%��;P�L�J��\]T����1�i6��b�:5�pqe�2�Yṷ���4��Xv�2��e�C�[q�۵���DB�P)4�U(`��r�qK4VҺ��c�k_����}˭ͦV���qT �{Y�������a���8���Hܬ�ɫ�ԔL��Њ�T�=�1�����%+���@����i�	_v?��V��ẏW����	���&L�f ��e=l��ϻ̂MK��U���M	��� ���f&��MĢf$-�a�t�v6��=�[�};ީ�Oč��l	�<y�G4�;m�9�����3�^���I���W�~��;]T*�\I�S��� ���v0�$F��=�g�UQ�F�~y�_!!��6gC[FW[qr����1��B��8Ze$ �!����Ϟ��ͬ�>O��y�~�����cv8�B�^˸U4��ǻ͒ ��q��w#�d"b"���� #11�z;M��#�(]f�S>���Ѻ��2�<�/�᫣�~���/M��왩�������x�N�wqh�z0��[3�}��w{n�	$/s*�&>ݎ4	+�ǼDȎqt��7��(�)JsB*�S=�ڢD^�!@A���x�践�,��̡@�c�8�č��b"&��L��y�ʸ��1G��	-���~�H���Ts��1!Ǟ�1�U]��r澉��(��Kfޡ$̮��]t�>�@�@����	1�٠Oć���ǁf��4��&���2��B�ݳ���8�t+YHjeV`���6��ʔ__=}�]��";������_P$������a�2|E?];T	?y�+��]�"�2D�M�y�a��Mm�B�p��)��H$�ݚ������gI��;�S�~�qW���<2��0��ۺ�D�Y��ٛ�w�UVS�r���iӱ5K����Ba��G����x_�_b�x��G���J�aۑ��w�Ś��_�s�Ͻ��t�T>�%�t�$��s`��<ש(�I�P��U�ޫ�WÝ#5>��I+����ws���������s5�9�0Uzh��GkDL!3"`D�5�`�o��e�cp��	=�S@�����'�}@Q{��C(���&��%DIM�t���@l o:7R�K	/��b�\��P�)I����J&L��P����/��_[��`�H�}TD{�v��1M�H緍�W��%D��e	��k���Oo�	W�`��v�$�kz}@��C]N��.�o���o3* ��$�lU����ݚ�8)ֿ�]_xgz�p�F��o�A'�\��~GCA�f@��!��=w�uy�\�`�s��$Nf��I9��0:���_�ڰK�-�5^_�îg��9�W���H����>ɋnn�������Z?�nMN��a�L�w*3�%>�!L2�U�?{�~l�+�ZJ"AP]I��T�����F�u}UUyӹ��3Ӽ�$�Ψ3�����^(����` � �!G�7�,^�����@�s��a�G�a�|�~�z�b̉�{�y�a�I�s�D�':�h�-����Msd�s���l.��L�S$�2���
Y1�UG�{ޯ��+�]Q?mt�ń��[�}�.w	Y��%D�&f�`�u@�E�e}DA�S��Rث��pd���O����D΃���0�	�$�A�o�N3>��#���Q �$��o3��T��{������(���X<��Q}�=�B���u0_�{;����8��7U@��ճ@H��͙���ﵸv�Ϣ!2L����ؘ�P�Oe��vW�5>{�n�f�G��#�F���Z~ʺ��$��0%��P"$/�zwf�}�P���͗4f��I�h�(�"���bJ@��f6�b���vH8h�fJ�\X���u�tڥ��gu�4)��%j8T��6�E�R�MV��e֨)+lY�Q4KR�3`%�c��ػ�� �%ƈ�Sq�(JlaE�Y��Faq4F
[V�	K�S��"�Skv&Ԣ%�aML�e�R���#<x!w�a��L\2�aM�Zgd���x�u�k��]��kѥ�&j���3�ڤ��2��ߟ��ϖ�ҍ�T���_�sճD�3+f��?'�͛�SrV�'��T�\�čg*�(��3"`D�Mw7� a���>��(�I �WM	��͂IDw����Ӓ�]�pFfT��HL�F�vh���	�¥{'OZ�U믉����?S���^�R��`�S�eǥ`��A��@k6�$�/�o�+�|�P�:�
�HJ"e/{�fݶH�" ӷ_S�o�i�l�Λ��:#㞟M�$U�9�'{����;�­�z�c.�Pj�ٹ6)���2��w(gF�	h���f�2�f)"�%O;F$��f@��E�j�����`�w��%U���)�Ϛ��Wē.������Pd��LUB��s�gg�ݳND	��rT�sث��f�e������������V3Zq�ʛ�7�e�|�}�����\ߧ��ޜ�ˌ���ə�ĸ��	 �_u2I=�u���{�Q�'_�|��F9���պP�Z�Ϋ'����_5yu[�~;{ذOӗ��$��Q�D��8�L��HL�V�w�(�RFNw��P"�)�s �؛�D���R#|]��oѿw���Pʘ"&	�0%7�}���	1k���g��f7���hTa��e�� �}}u��1�܄�T���4ǱPFR��(�.�Lj�
��1�»����,3.��E�˵�A� $�6_&L��K��/=@e�Q��do*j�uz�Vug�/83�1���~$޺~�ap�2aFaD	���]P��d��ٯ|k��r�H'��CB`�S��Q&�w5��=Ƣw>$Og2T
!:�P�k����՝_A��/�2�n�G�*O�����s隵yz�5-zR5~7�4a���md=~�������Y�Q�u`� ���bC9�ܪ��އ�k���FnzE�Ɓ�9VLD�* �K���6�:�ȟ��]P �w6k�I��z��9=tu���r}u���Tə�%��+S�@�n�����f�O��E��Ċ��Q$��(�շ̓���}>�D@��GI�ať�W�FjJ)Ҽk�ݞ	L!�]�,,���<����Y�4��"`�3Wp/��"��@$���bg�ht�G���$FFZ�M��}��0 J"e/Nwz��1�w;j#���������?�df* �c�뿉%vS�>]UZ�Y�^��v(�.L#�(�-�yeT	;W�L�"��e���a���-�o'M~$uvc`��wx�&Q�N�������M���Gf��^\z� ��������=�uVW�x�ֳI�P��g%zU\۳��s�>�q�U+e;������y��.>{������=Ԓ�TQ;�[y��u���^^Wݞ��7j���G�/=Á"c��E��TI�12�
M�Ο6Oğw:�/����Q�H[8k�D��'1��;�ꯢ�l�{�Î���� ���"`@�Pe)���fu+��	tـ�2��0 �%�S�QϿ_=���L��)L��ƚ$��L�A#��&�,�+�͊��O��/�`#���SD�0f��>��Pu�����4ͽ���x�_̃�;��P Ӷ���egcwș�$�&R��fm�� �k�G�	|oF;d�Twz���k,,%���o�H��B��$��6�&	�f@��}��*���
5f�ks+�'{�� ������{���k���|+������3Q�N�DԚg�Y5� �,�y�[g͇R����H��s���
��o*��*;�|W�����AH^_sSN{.���W�O��"E�U�Nը��>�l��I�{ݹ�C[ߺ���yO���Ld�8%����67)�����]1LP��؋b\̨�ҎH�:�f��a�6ⰱ5Ъ�Mc3uca*��Z��vH0v�˝%����;V�XM&�S(�p���X��j�E�bT5��&�%B���%�5�!�75t.���_[��Sc3i�uX���0B��5e1z˳oY�iutb1�aN��m��I]���	�c	 ��Vj���A����ff��cGK��D�kS4�)�"�J���m+7�Gߧ�r"b%B)~ʪ����o��&<����ٟT�>l��U��&�T~�yQ
&fd�X8��A�8Z�zh�G9�	/�?P��T	 �a����Wd���b�" )�`�	V+n�a�]�(I:]���)�ɯ)�� ��=@P ������:�(D��JM�w[Q�w�}�8p@�/h
$�H��Z�Aݿs�f��ڜ��וB�{�D0��a�%�5�`A�������c87�QSc"2��&=j��P}m�t}=k|#��O�����@��%�[fK��!�k��"����p�V��&�W�߿a�S�.p������$�o��s%�w\{y�o���E��j�$p��bbT���`$��o�fn���JgkT\]���p�t�NX�ܻ��/q�;�=|����=9)�3[�^�ٚ�q�����ׇ27�]��ʮIǣب���w���f���K�s����"kz�H��)�x�.�A$�w�����;�pq"́D����u������	�0%6_s��J{���g�|��^S�H$lw��I;�i�l�`�ӗ�~'�T�(��l ɉ)�����l� �m������D9s���C��H/�����D�u����מ�����i��]�"�V����XA�`��ĺ��%�+]et�ʴ������4�uVo�t�ڒO��c��$~��1#@IvtQ �s��۬��(�8�
jMX�˭�
�sS�۰�"��ng�H�c�` �u����\��3��\�5Ǆĩ
b`�I��޶	���D���z�I� �=75j^�c���"H�Î�:��ͧ6��Rxh����!�a��\��Rp�=^6`�۾tb��� ��wf�g���y��f�쁆�b�)���,��+vd �W��bhѽ��O�ے�y{���P��?�̞:`�������/��)O�pM�.�a��5��Џw>�]��;ve��G�NSv��!'�_A��nts������*,���{Vl��뗷;}��������2.޾�j�����+�#�ۻ����:��q�}��w4y�5��'���	�A�p3��=5�f.��#p8�y�A�dz�g����ԓ�h ��}��f��}��k�Jq�F�ѻz%��`Bw,��}�2�M�O�ů�98H,�Y�h&�����f�e��7i��g��>DJc����7bGu�S�(��ϥ���%X�|3�����8���b��d-��󢙾��0�����S<�����=N4�6��bNPgNS}�7��;�M��G{���/�+�zn1�-�=꼣����s�H��ssf��B����O��=�ۅ���g��S^��_B�����[�ںHfcb,�u��D��^��~�R�E���.���}��.<�����}�O]~��Յ�H���l��y�g}�{����/V9u�Si����g����g��J������-#�G�K@�೵0�:�vn'�����qvb\t�CV��d%�ө�׳����n?{�n3&P���y��A_��%�jӱc{���H�����.�B�'�p�`V��Zq$1QF�d�$��f�hJ�����G��bQ!N�ώ��^�2��U�ٶ�"�i�����u��$#�Y�Eu ��*��m����UpmF�"�f����V�Q�DT3A
)$\D��Kr�r*��8�r)��4�î�P\#��0m�z3�Z,DE�3�M�EEME[ibv5p���U5El�ՍT9���b"ETB$A�V$UQl15��3S�͠�SPTITQAL��gm1DTTSň"���L�Eq.�Y���ERlb4j��"kgZ�m�4��Vˋ��b��"f���(�*8�$Z��S��F"x㇉��1UL�U�SAm�!��G�kF�j5I�� �fK��LT���Hda$����AB�YdB�3,Ȋ" �W*Q�DP����i*JA1��HQ��%��+1TpqAcU�D��P?d�?~'���g�I��uDD��Q
$L̂�%��o�]��Cx9[S]� fo��Ęoe���:T�f���'��s��&��[�~0}}SuĻأˤ���=~m�	���ȯ���E y�dm\Fz��
j@�MGC)`�
hWCQ\[B]l������eX�QS1�1n@2��Q'������;6�?���b�z�g?�s��'w��z���	F	���T��>�����N{r�A;�s_	���(at��]�����(Ȅ�)�4��V�@0{t�t]�˘�=**����˪��]}�ѥ�%���(c�����Z�v$�9�	���I�����{�wZ]X=�ϳ'�o	3'��r8�݃�M���س�E�3އ�I�����%�g�!ks�q�w#��9� � e,��	��n�s��:1T� F�z���ᨅ&fAS�G��$�K#�P������؉
��$�W�O�}Ϩh�^>���ˇTpZF�\n�@-��� X[V�2�v� �d!nen�Ė����	0�Z\j�L|���}�Xh=��%�����	0}y@I��F�_6���A���H���YW�%&$�IlVvy�ꚯmcYyϞDD+ˊ�3��l��՛�9�>���B2�&l���A'�=� �%�KױC:L���O�+�7�z�!�u�P�N(B��Lޭ������v3�Y�u'�A�}�� �w��x��t�T(z��i Ru�_�J�J3!)��)��z�$�w]
�.��1z���1�~J2��ʼ����{��E�63}Q3�L�xjOٓO|��g�Q�x=Aa��#U���R�nfQHi���Y�ͳ�م�V��)V]E��|o��o\K�V��4� Ε&.֕�Wl���D�̠Ě��_7��]��6��B�����̼��Z��^�(�F2�/:)&լ�X�F+L� �0�-�FSltT�e�7x�`���F�#��Rf��-n���QhZ��6l#ae��E�]��d�����צ8؅!��L�M$���y�����77T�ehR��qD!�tkHl������uEŶ�6:[e�)�+u"��CM���֬DL���������[.b�+����T�~��SO��G����Շ�4	O6+�	��&�J���D0%6_s����Ŗ-��$���w��đ��U �+|�׳4������^ȔL���Q%���6A=�s@�j#|�õ'����̵@�oe� �{���0�"�
&`�����]Y��;���N}+iՐNo�h~%\w,���au�퟉��k���ʔa8�
b�{W�~+Vu}tp����$Vy�d�/��(�
�yQ�����w��s����L%l#��+��M�0�ih�K�Z�L�&��ɰ��>���	Fd%�%s�����uQ$����o��]{�qw�f����P� D��J*$L̂�'���O�A������	�z �Gy��صK6L���K
��w��{�b�>�����n1�^�����[閬����o7d��L�7����E�g��m����{hW�B�*$���G'��k���D" ��)����~*�b�a��2UnOǯ�T�n;���
�D�$L�R�-�Y��k���+��"����� �����{��$�~���_N��m���vH�;t	n]M}����0R�D	�X�,�A?ǝL��:,7a`���U�d{�|H���u�E����
���$.�[�i��j�Ƭf
4�̎s\Y�-�-�BTD�J��ģb�4+�{n��	b͡ ���s�����CHx�=��_�-Q#`���&%�7���� �t�vh����'�WE�I#}���
�Y���k��e�T�^����(�)l�U� �o;�LI>�uΉ9ɱ���ɋ�ާ��l�`��u��=5��˅Լ4ܓ��*�8�����������sY���K��N{J�sxh�o�wk=r�������ߋ���+��>�LBBP��}]��U�W��AP��I�uﹰOă������jU�~:/㶺���"D��$�M:��6?�m}S��CY����TA��͂	��WՈN{�"��ѽ��Jv�v.Z&�3�
�ۃX�dÊ��e��nʇ�	�*bT��$�JQ&J�6ֺ��'����I�������W
o��?���P$���d���11(�u$D�
{uAzz�'�{1(�	���~��S�+��x|�7�g_Do�Su����k�@��(�)���7�$�w�h�V^�#���3����k�x���@=�����RS32�A�`�U݌�x՞��oވ}V>$PH�w;B�\o.�p�u����˶U����dc�#}� �Y��W�w4c"���r{�<�}oO\��<:/#=�~wyd�q��i�r\BHVRC@�Z�y^F8��$U��Q�$%	M���@�U���x���1�����Wo6I?y�D��;��oo�ߕ�����}�opiYu�̓R��̬qĽE�K�����ٻ�&�J���__��)�]9�u��F綐�A.7�|mo�;�wmB��l';m�@>�m}V�G�P�d#`Īg�sTw|�����_/uւI��޽� ��֨�����cw�	��,LJ0�	11B�5ޝ�3�Ahf�6�bNTG��;8{�/z�1{<h��"�Q?uO������/.�����UH�����}β�R�F	��`��ʋ^�R��12� M��O��e��u��ꪠH$F�x�_g�s`�Wtq�e}Ó�w5-��ۃ�d^g^��/.Y�}]�\M͵xv�u�%`E }��G����w�O!����s?Iă�/�"��Ӻ�;$����:�p�*���׉nE. �na3�y�+n4,5��Κ�L�s
Z��`���B��"GLQ�b�)6H^(�Az�Ս��ւ��b��[�JP�&�R$�c���Wqr�c�R���ɖٙ���h�`J��u
�5�m���ɉ,��b�ܓg\j9���ƖV�R^v. �
����ZYv��C7(�e�Kj�f�H�j�m��B:1�+y�4�b^P:�b�4b�M�kytզf����߿�Ң )�HJ��?>�TI1{EGy�6	�y8�{�߶���m�&+B͑ I2J���3�g���D:�q�Kݖ����?gN�@�>�� �{o�!�t͉{�ɓ�P�R�>|���ǝLI�����U�K�7~$�S��2A?������3" K"bU
`�{aSՅ�d���|H.�&�'�@$g=�'��݁SP,�خ��z/k���R�BD�"Q7�>�����B�y���>.}���k?w]U[����[�d��zKn�YW�^fҪ;1a��Y+�qp���,�U�p�篷�[V�X���'�?��>�H'�n2s�O!~P��z���.�x��;�O�{�䮔PԌ!0%6{�Q�,���DM_xuT��ܨi0g�����Q����)�8G���I�}<�ĳ���{�^�
���VM��z���5����/óg��Ŀ<�̈́��+�[�_���w}χU`^�"g�$�D�Wgy�	7�u@�^�|�N��|G��S'�N�]T��rd�20T����Q�u����l��7>$�m�<�I#'��Ldu�39�T�h������`P���L��-�T)�[��I�W��?O�����H���6�nU@�@E�������O���?|t�1k�1ãt`f�p<h��04���m�#2�J.�g���k�F8�kdr�dW�qܨ��u�b���#�n�aw9UP�h(����3M�yY���P��BJ���m�{4	%_O@���x��+}[d�>��Ʌ��0%6z��B��5��\]供��]��`���JW���3<��;|5�L���/�MO&8f]+�;l��+ɐ:ou|��q��>�o��n�HC�������@�}h�/G&~PL����[�r�=ws����GeP�PA��^��s��ޓ]=��&i���'vǤɄd(
`�M�=�E�L_c�$��u_S��@�^>�Έ��z$�zHA�n�Ԗ� ��lҶ�-��Ե�bېR��GK�jŹuL���_Os.4�B&U
��n����i�!��a���j��=n��[�T	^ȳ@��J͘Q���
o���7�1P�:.�]lo��1�<h~�������O�wU�M<3��Oo/��G�q%)���3KeeGG-�S����0p|��1ޱ�;�I!��o�C���Ʌ �`Jl�����,�=��$�S_O���$�_o�5{�^����r�Fe%����*=��6�
��\�����T�f�'�zw������~���J�3�����u�XhpeLŚǙ�2eO�	����0Ⱦ��Qj���dG�Ο'�s��'�{������z+�L4��vD��ٌ�КYy���54��J*h8f�8��7F�e�o]���ݖ:JM�����=��I7�6�?�}VS�=�,l�4^{�f��O�H����;t�0�CB&U
`�m���ٯ���r���pn����@$Ge^7��}B��^z3����W�x|\I^<eD�U1=>�Ad�����^1o��+k��8�$fU�`����5,����ĉ�B[N�yɮ�5�ԩ��/��H �y�TO���ũ��}���P��]׵��=2a@3L��l�� �de ��x=�2�O�sĄ徺j=����G��{�|��?���O;	�"�"���������W�)��
���3��1��(E�EA"��Q �����! 5�% ""T& P"b�ƈ@"bT "&% ""@"   �V.��V	E`�V�b�X$�^y�8Q]��p"�ɀV`��*�1J���`�	Ī!E�X E�DX8���X'���H��H��J(�@��H�,"�
,"�(,��,��,"�@�� A��"�:c��� (�@�@"*�?��y?��]������~������O�q��c�����c珫��x9;8? �N���������~�TDW���������QQ_����+��h~�~��|���������Q_���{��?/����<?���08���~�?a"��R�D����+��ȫ �)�)(� �*�*�@�!(�����B���J��� ��}�""�ߕ�����?�@�Q�(PK�>������<!�����~B������o��S����������c��v>��TDW�=>�����}�� E}��"����������DEg���p�(��s�@g�vNG�;��?�݃��pi��x���G�}��9��Q]��}F���N~����ÿ���}�}��z�������"�x���<4����=�7����q�z|~�WH���!�f<�hH�xA�C��|=��#��ǳ��p�~=�EDEu���������������b��L����.��� � ���fO� �G���                    >�      4        p  �@  	@ QER�$P��� (� u�( P 4 P�@�ɈZ �  (�w�                                             �CS��� dbX  H�`ks2 dӶp ;FB��5:iJ(V��   Y]� �f��L h�T3�����޹��H�* �
R��T�4*��j���+��T���ҨU�% �(p   <         �*�JZ��*�fiT�i�4UK�.c��
�8 $Y�]5*R���fQ=�(U�rԥUNw@:�J�4��ʤ��8W��5��   ��Y�5, LF@��6��  �H���E(Y��i �T�   <         p�t����@; � 6�S!����L��q 80 3p��ŚU����i�  �C��˪TWg ��r��f���ɵ�3�1�����S\ �a5���ʹm�v]�bۈ�S����kf� $ kހ �        �zV�&v������{�ިl��t�B� 䂝��6*.YS��sh�e�A�� ���Q������sp� ր��  ��qoYL���c8 �-����k[�mj�qi�,ۜݥ4�� ]يӝ�-AW6��\̊�Zsj��0�( ����        ުz�����D��M������Zs�j��p -u������Gk5m��Z��ҩ�5� �,�u�T�p  hO�  �re�ۛ��\p .u�S�wzV��59�r�m��/y���p ݆�s�	���l�� 5<����C@ E?	��%QC �D����OP  D�2��IJ�   �=�L�T   $ʔ�S�T�I�b0$Vr�-Rs� U4�#�Dd���6�S�@m�o�7;������c���0m�o��6���@�6Ɍ`x{��o��G��B����*���,�)Q��-,��[�Ǔ��/v=�2Jm�+��:��kʥۄ�]Q�8h�]��ݜjF���4*@�ݲ[�H���	:�Z3���u�x"����fA��,������#}AU�;.6��Vv҉������n���G���<2���	p`jÇ�ڮ��zܽ��4�S��A@��c.��c������>=r�Zz&b�N�WE�oZ��q�׳�H�\�l��	�^,U\��;�L}� �
����w���!t��p1@���	J$��KZ�r��"�mM#��Om�(�x.0�(�?��A�$i���;�0E�N��9��Ֆ�ۨP22❜n���c��:�=�v��EZ���ך�αf� �m4��6��D/������̢�{�$�0��$�j��U�j'��}/K�z��s�8�aK������-�/�5��7rh���tKc\E�[2�IX�R����f�����9L}>j�[Yǲ�#V0�;�h�)Z��Ll@��]2aM���,MeׯJW;9h��.jUh���S��$\���x]�O�@4웛��i�񜞳����2��wzЛO����xjՏ6���IxW�����H��nmE�1����;���*n����7hlp%�����_L���%ȅȩ�ٻ��[��:r�z�6�|`�� ���7��Μ3E�8�8+��v��sӴczu�O�ܘ¼ˤ2ISL��m��n,/h=��ǜ�mȮ;{-8�r��m8~�O%R��F��Նhѐ��k�aOV۲6�|�.���q9��\����Ӹ��¦\��r���^p��sܴq�H���_ϱ���B@�K�E�:�N�\��k�*��k��p��֝��i���l�V%��i�	Lyw�Q;xp}�^�w{��k�1�;�q��2w�m��(��݊��:��ލ�ot3�4�ތ�+�4r0��gL�r#�m�tc�#)tԴ*z!���>�ɎBF'r=.7N]!pi�=j�B�.$�g΋�~�n�]���;�^^1�Ra�ڒ]��ӳ�'pW�d�7����;�]7;{W���z�.�S�R��5�^���&��o"����>W�}�+�N[>��&�^Yo!�a�V�#i;�CczYO%�9�V�vb�ݛ����j;u��+DI��n14�1tŸ�@�����=�vUQqG��4,���yӻ4�=N��D��������.Q��FgwV=Z面cvjbg"�w�:�=1�K���qQ3po|���%�a�C��N�8��ܤa�r)nr�9��ǜa2[�981t8� ��۝��tn.�����o��}9l*I�{'v�C�y����n{�������t4����ش��q��O�a.L<��V�^��3z<᧻&o@̺��]]U,�rM��:����Mu]�Щ�s�DC��ܥQ�u�E\9Z{�c=u���N�t�ĝ�R2wklpc�5)��צ��%�V���[�Y��\���VGL۫��4Ձ��1�Ƹ>LȞ�3��}t���xn�u h��E�Fu�lͺ� _��WTâN/}��6�	��M�OL,b��ۃ"��_n�*�.n�ǃ�swHe>�L�޸�6�X8�{ie�;�E��wQ�S`c��Qv�i]��8M�~G\8V���dӹ4n7s�,����xyJ���Jl�hnMoN<��ks;�.���YH�Yh΃M&�66	o�W�&���ӽ{�$�雐��"X�B挏��bS;Kn'ä���4�kq�U<�T����1�{:���/t�Wdf�x�`{����Ǝ��Zl-���Fj�f���z����/j���g��iJ_N-C�Ώ&ݻ��֣��\*h���;`�F6�>�/f�p}Ă�Vu�9+�V�F��h[��I��bY���PQ�Ջ5���ԑ�:;dN���9r�z�+7�/gq9ۼ,Z��h�muˏ,զ�IV����@��M�f�ѓ������q�����EP��͟��*a�w9n2p�nSY[�`C���B�$�֌Z��� niuэ��k�+]x�f�T���!b�v,�4\� ,]�p��򌘂��j�+A�i��%�X��ww�JB�y���t�yulۖ��n:{z�gn��+9tl�O�S�ސ�n%ٳ�wTt���Rw]�pY5f�k�sn(�*��à|f,�˰v!x��횴ϔ�/<�d�#����b������̓��՝����&�7�r�8.8���xk����)����ً�������X�7��:3�޳��Fw,�-Qk�|6C�,�$98_#�E���t�(�K���hD�qB�<�9��<�ٛ���<��U.b3Wk〡6U����F���s���cF&�:p.֫R�w3��K��۷�w�
L1߯��9�bnv����p,���9��[�$�*�3��:�.����؂[D��HD�\[���D�F6w{&�Q�RG�ٛ�TZ÷�{ڦፈ4�����7n���FtnDIs��a�9�&nR3Wo��@�h�o|�^v�xX�΀r�����ڕ��>e�(�p:�:�͋WpÇn0���\����y�7���wG8M�p�ó�}w��~SW����>�J��Q����j�7S��.����V�F�R�9��J��@ޜa��7��hGynt���up�����13���X7�Ŕt8og<>���͞k$n�����;)4��e���]# UҎ�����ٜp2M����m[e�/KN��Y�i�D�jS]����S�e���(Ȉرs�%M-��� 9n���%;�\6*_۸�w-��wU�7Ή�kM8�sn7Z�}E�wt��l�z-Sz�WX`fķHz��馤��ʼ��7V=z�5�k�BX��݇t�Mᄝ��A�|՛3F����F�͙�s��������7[��&
'p|EXD��;a�fXB���gU�wt��	�q!\�b&\`��U���@������4��6�e�wr���dH)ǉy1��	)]O�M�<�׀�j��o�˸Ѓ��(ʖ���䮒�a*(��$8p^sڗ7#`l"����7��h�c��O=��u��*g�7x�B~�>���(a�&!I7�k
S�o8�>s6-AK�q&��ݶ����n��\=�mx�c	���w�ְ�l�y=C5�<�s7f3����ov�Ż�4N[����H��w"��=8^�ѧ�4c{b�
q�7gs�����P��3�v�$���j��:[�ڡA�W��\1+�����Y.���Z҇�+yIӭ+�Γj�&IϨ��}�'�q��Eȳ��㼹T�z���Z����{V��i�2��!��ɀvUMh���a� w��i��6��\g��1"���BjbYع�@�S�B+Q�w]X:�o&�..y�rǓa�p���V�Ԧn�ॢ����8�nN�I�Wv����#nw�f�e��@4��nz}��;��/N|��Hm���c
\��` [�p$��Ӑ�%�byc/%�.��qi�qC��M���tm�Aſn�=5��錆�gt�sK;;�(JW#�JW@��7�W8�9�����ٺ2K�Z��-��xǡ���;w^#��n��{AXRh�S�h�MM��q�8d�(�J.c ���ܛ�p�u���Y�Q������f��]�j�,�`q
il�8x-J>�Yw(�$wb]��B|ʜ'�I���@���^D�D* �0EɊs�#��v݋ß�;��L8Ԧ�J��7��x�n׵�v倍�'p�3{Z����K7�ٝ����;�(�]�����	�@�=g�xΈv��(n\��; �z��L�dgVM�6vG�ǱI��\����zNo�n��8.��v	��%9��m��&�ld:��tp�{�CIX�i�S7z9�Of���ݛ��0��{�l�2�s�5p��8S:k���wNQ&�1���'G�t����uu8�9D�V����eմʈ{�Q�KͰ�q�jk�,y�Of� ����L�̳z���Ȅn�� �ԮTY�L���i[;�n.ٰM�z��n�՝&�vs�(i�bճ���9��_NK-��J�ӵ��H��d��+,��ъ�/uք�ѕ�K�ul*�c� �87^[_7��Xw����8�lYJ{�	c6)S���,���&�˛ 2�I��'wy�GΫ��E�x�ؼ�-�q���]���ܝ�j�ڳu�C�*:*����\��]n4��a�{v;���hҶQ��>�����Lzg��U%�9w�'�s�8��k�k��<(���l[(�����{SÛ>m�۷.���<{��7H%)ܺ"�VJ�O5�������뽳�[k��K�&�=���3p�+�Ք>���}K�q�����N齺�ɱ�&"��Qӣ�"[��'�e�\[&ii��a?r���A�=ܷrs��ؗ=�ۨw1�t�*���uX$} ��J
�2]_ޖ�XZzbm�;\����ײ䐁"�<���Kՙ��ܪ\���t�����nb��X�9W�A�H�`[>S٧����{�q�0��l�Ա����x�S�l8!0� �V�r �6�i3{wtRe.�Z2�eEܷw��p�##�x5�/��L=S5>�CQ�^+�n��$�N�hC��\�h)�MB�!'e͏�/���a�+9�n[����_SD=��4$�f����=n�'n'w6�UV�����s�%\gw��v ��eKW^`>���v�%��r�M�a9f��{NN宑3K�ʴ�-�UGV���-)%�ͼ�$�9���nL�����f��ig"N��X��KW��{��`b�L36j�취���f��ηK�t����%������p�rl���݇O0l�؂�c ��*�3�<��.�X�U]3�j;��_v�zqX�t�p�,���x�n�l�[�N.ݶbn弓㺨�Ή5���Y�������o@;�4v����p�H�_t���N7��y9e�T�P�V�D�	'�-;�RHw�o����W�t5L3��B��{=vm�`�����.q�n-찕�㻁�wH)�a�d\�������{�ס�q�C7���Y��M��d���&�6�f❩W�����ۨH���5����KV��e<%_DTĠ3l<k#�������M�7.L�2;w.�d/H��<չt&uR�gr�`�@��5��~oh6���٫=�,�	���1�9������%�d������`ɻ4^�W�e�����p��x�{	��=����hQ��v8���Y�)dpR�\�8l�ݭK�r����ME�4���� nh�n�:ss;7c����{&,�wP]���];*@eS<�MR�Xl�sq'�N���\��[�7��k�	�.]��M�\��H��I���}�Ci90a�a����Nɽ���[�,�<�'���Vp!��$/�o�os��-egr�nFt3��`e:v�UZa+�zaU� ^�N�X��z���A&3�9o�x���f:�)j�w���:E���Ykj��PW��!Ӹr�4V���Ѓ�b9.���tiks&ݺ�
��M5��(Q�f�>H�%rc�m�s�<���4�=@;7�Oq�d$2�w��Vgq��������e�ރ�Ȋ�n�����ϵo}�9Oqnn��5���
�`� �3������B9��nM�`�z�!s�Z�2j?-�\B���f����j�^�%]�rf����	Y�C��H���n� ]��7TYϕäl�Y�!�k.�^1��s&O��..M�tV��>�����^�)�7��n�Ԛ�v>u�k�#Hc8��ydܤ�[bFR�.ϯgaN�r��޲��l!�"٦�G�k_Xm��ڷ��ڇ��tc��^������.�A1]�y�L}9I������*��p̽7��=�F!r*�f�^��BB\鱹�Q?v������hb�wT3����{��x�\g;�BPp��!�YƆ��uV�(�@��8A�)�N�b�ې��-*�vR��ӯ�W�ǤaR.��;QA����՜��Ysn��FM�E݃�>;�*	�h����]�CZ�#nb��6Z�=��E�d#.70�X�0�[���2n*2�ǔvE�s�vv5����Z���M������2٠�~Q�3F�m�y��ѩ�Nj�p�c�8�,C�f��ގ��0"[v�N��2����B^n��T��(�kG7G8���\y��5n$���nl�c��Hx7�C[	
�ټ���p�/K�������wB(kKNJ��,F���		����ND"��V2.��i��7w��>L2HG�<{����su>ۑ6Lޏ]A̽�lђm����1�#�tC:�¹[τ��ixN!�o.���1�KO-h9��e��يuwP;�,њ���(���x�c�5��^y�J��>���wi�7E�̻M9�Ԇ�#l�DCy��{��1:�q�q�]ػr���P0�it����1Cܝ$��6Ԋ��)���GM��{S�.+\��vCdԅ2Q���?������{�S�����81�62��
\����e�����.�(apl(�l���Ɛ��aM���v�$�l
`�i�]�P�l)�
l`����`S)�ˍ���P�*�`�;l�  ��2�
m��i�lI��(
���	�v1�P��M�Le���q�� `]�(2�)���( 
N�2�i6ě)��l�Ɯ�lm;lM ���62��\.  p62�`˃`Pe
˰�lHlI�� q�!���
�&��l ���ˍ���1�����m�n�����}�����u����g��yu���ã��E�.:l���d�ft˲6w�9��xwk-�ͭs{�����tAѓ��Ί�����̈́�Y��j1��h~����Y�ӫwS��R,<����d����Fl�C�`���F�=7mUrxm�ʨ��@�u�tȀ�00�T�g�p^ã����u�5G^ܿ_S�ȭ�S��h���{�w����7{��>�3���7uj�X}�]�7q�*�8��v�W��B�u��{�Lxi!�fЏx�6���hZp-]�d�j��W������1��pn�T7g�x{\�t��$���"�ݞ�k웞þ��!��صz�>S�W�O�VS���}T��w��8H+�)M��8�u�#E�ӫ%�4��է�]݌z1�F_z������u��*$��t��pѾ9�A׽}������qOxu~}�\3q_�S�"����w;��-]up�׀>��.�쌂^��W����\k�o��+Ǯ��}@���/dg���}J����<�s"�ӣ��M�廬>��8"+d�B�u~<7�;��7���g�<����j�k�p�G�u_w�x�
�Ël,�����X^��1;�þޙ���(#�(�8;=�� �K�`�����e�]kW�g���5�tqx�����Z:����9�g�=4
�}�ze^q�A8��<;�m�,��Ͻh�'��n��CM�Z!L9���W�uhUѽ�4�[(��"��ՁZ�0�n�N�����1�uJ�ߌz{	ͫ=��%�m>B3���N�۷�:�
��f��~�'�r���߶��!�p{T��]4�{4�ӯ�z��"�J�XX�s�)왾���g$*-F�	��<�I��������Oۓ�7wB��1�d����G60fi�e�%q�E�}��&)�\��][��8��ս�n��N����l����,{�myw�q{5;g���O�8φ��s��o/f�c���"������^������T�S��y:����u�hw��2Y�o����@�~����9�x�J�ENF�5�N�U�W��2�,UvM��)��-3�nw��bPi�=������|}�:MI������-{~h��a�}����C.�xY㸏T6�.�r���9����S�s�}a���=��"{��,��k'$��+Ǵ�xXM��Z�>���ds����<��nr�˸��ڶ��S�yz�8���!�q���M{L�*&;��	� ���!T�;�WRp�w���e��O�p2��� �su%�sT��RȚs��H���n��)�p����P�j/k�ۼ�qԳ�����'�*T�'O�N��/mcwp�`G�<!O{-�φ�X�Y�Q�P/n�v��s38�I�;�zlĞU��ӯ�|�z��b����6�C����Upo���{����w�����ї��,������=����S�bʔ�駼<�:U�~�{�'����������#�M�ݛ�'�<ʛ��q]|�+��$������`���Z0�15-��a*�;����{:xiԶrڒi<������Th������ۃ�ֹ�~�|�	�Opp��ko�4\	n�l2�丝�t��C5��\�κ�I�ٴj��;��OL��ά]�q4�vg��ކ�Y�U'
����܈7��Z�Gg-x}��������<��[DZ�L��S$�U/h��74,��-=W����Ƽ�	����H>���q���������d:9�u�-/N|��ev����ǰC+�ʯ��b�=��F��${�w����53�ؖ�jʶ��tHt���4f�;J(=/�ڂg�����/���n��]�DJұi��!�����rv�mD� B3io/-�f��J�잟��:�M����a^ټ���Nl�׾ov{��T����6\��t�r��%�`������|-/.��D_l�$l�&���W��g��T�u*���'L�M��/�z���x`^&�ը�U�Sٽzl;2ePdMf�
�R�n�>o餕@�r����5{���+��N	,��$��ۊ{�r�;�{D���X��q~$����FJ���K0.�X[S���9�-��f�AB�"+�Ò�Пt�a�&[�'%�g��b����2�ZP��gK=������=�+Br$X~솓�z{qt�O����#��㯇��;�wdȹ/N>=���,���m���m�V�"��|:/��XÊ��d	zg��*�nh|G�L�{S�]W��_6��7|�A�v��ŃF����F��`�ڢ� �A�a{�l���5�Nc����-r��,=��G�@� �Xu��U���z+a^��&���D���8:.�Ӭ�����_�(I�*ѧ�9k�@�r�1��|�������ck/y����l��c2]gQ\��>��X<i�Z�/gki�q�o�_���0�>�f��{F�P'2L��7��3���p��D�	��vj��Vgon���2:koZ�<�xS���u��_{|�Zڝ�Wp'Vޫ�K�z	�ܜ�M�:��@�ѷ�ݹ�����1)ܒ�����>�{�{�`��sX݂�6W�xq&zQ�r����������w�F�V
�u1u@֌�41�ډW�8���{w=�H�ejN����-.�ǆ'gC�O��d��G�n����B$5���*��_`*<��k�iS�Y�oWV۬7<�W���/�5���B�����!����O����c^cվ׳#������N��_-G'`�b��fs�'�����x�g���o�_s�=�yb��]����1�Q��g��XK@��U�sx�[�_����t��1����Ή�:R�]��:��G���6�G�{��Pf�ۥow�[��=����T7�}��qh����d�8�wz�L��FB�;�����,��^��/�j>�Kk}t׳���|0��G�x�or����G��65h��]������
wv4�����JO:��w��D�Mڼ�Şü��'�5�t{s�� S|�l�|xD��^��c��f"�}���E�E�kgD�ag����5V9���f�Y�*���s_mшK��Vo�7�7v6�E�#����16B��B���U�0OeR�ދ��%�~�΃���4Î������Beg�����Ro�{q��S��8?�}�d=O<z�����o؊��{z̑�p�@��U`�w��뻼��f�:�߶y�(w���+���N�4��R�z,�xK:E�Q%����>Вƽ�z继��3���/}N<P��`j���c;�vss�;z���:	5��=�TǼ>�&�X����z�?q;��J�Lě���Էa��;�Qrm�ͭ�����8�h>}<A
���0	���=ki+[b��T���YG(~������<��,W�`��n�@�& ��Y"Bu���wcrġ���{�z{-tgg6<��/��&w���%h[p�d�����jg����W�3�Ʒ�k���Sm��MP��]�z")׫ a��Zs����Z�nP�w�$�挳��Li�t��DCñ�s�
~�c��~���R����#jk>�c���K�a���&OsB�_g����In�gN�^Ҝ�h+�8f��)��=F���j�����Y�N���{sJ�%.u�e4�8��[qm>��P��o=m��!��Y�"��⟍�z6���|;��vu[k�ӟ�x�Y�Y�f���w,Ix�y��[xF>���j>���/4r��²��p�`��s�8m���&������g���lVz���hd8wR�V��(J�6cZa������ograyw���j��Ƿ�/z
��RC�Ӏy�f�����,�	#�x>����:��o�l��v�6��7�δ%A'�5�&	��z��F���L/��S\�^<�����)q(7Y�=�G ��X��}��S���]��w�y�}�{�e��N����}��bn�O�������ۓj�45���û$9����*�N�皽�}�!x�\���I׋s���OhѰ����4]7(ıﻯܜ���<�����8y9h�͜%n{�H�ܖ�!�uX�j�<���(e�U���~����i��f�?-87x�DH;o��k�k���)'H�Ò37o��4.�E�a�A��Fb)�0ش'LX)Auu'M��j���ӱzh8oV;�� ��su�٣����<�u_M��8��тx7��Z���r��|�^'=�w�A�Wx)⮵�Rmb�n:^�ح��*���?Ytǔ�׻={�	٬{r^�(K@[�{&oN|�j�:���z)Ș���g%óe�_Bέ~�ܽɿW�=����ݰ ����)D��Ow��{���趯k���v���=^�o��9�����a|w(�f�;N�Z�Ѩ�vn�GW�e:��9%i�B��[{oqT{'�W�n���;/�o�L�V-�v����ޝ���+���!��}���$[��b��&kc��F�.���<~-��g�x`Y� �w=��s�Ћ�쬎���3��s
�q9�N_M�zz`���\}�ԧ�/��L�㈮V���Ū�Z�Ӹt�mɬ�,[����~]ݞ�w-h�y�9kO$
'���ǭ�=}/�WK��Р�*+V�E͇�{�(L��9ݽ�.�K��;�Y�ɛ���_^��vO�|���?{X��I�fr���֮�l��u�wd��W��3��P��{<!�lH'+�O܈�ZD#uL<���8A�3z���U�v�ǖ���qھI�wF懮n2�ʧ�tw�O��=���g7��Nw\�x�]�U;UzG\Q-k@������g�&���1���\�Qw�s�:1�)�CtƂ�L䧲s���,����7H`c<4�b~w��a��;O����nQ�:hD.���z1�F�7aը=�I��wV��Ǘ�^V
{�7��t��En�==�4�MO7ӂo�cn�ʽr`�9�ڪ+=�n��ޭ���YJ�MP�,n�}?\h��O�{9��iˮ���a����$snV�^<}�����^�8�?�}�+p����+�_r�4��^ӕ��hl߄�왶��������Fr�iō�����[����w���(��{�G�r���z���x�w��b�eUZGQ�WAh0-���Jf�:�p�u��K��-��*�{�G.�'�s`۩n��s�5u
� �%����c���J�xl���
^O͛��P��s�Gz��o�Jw!��{&���}��k=������C�=�����j�- k�۹=���22>+b�Z��z�Q|f2�g�W�a�{kcM2�E�i��G.��w��o��������^B<��~\;�K��&!E�e��b��vʽ�,Q:кT�Kj�w�յba2�2r�����\[�*�'.7j�7A��3�r[��8E�X��	�e���Y���m,� �����=]��~s5��_2��r��>�w+��?��p������ܯ�����ˍ2I��ڌ�]��w�'�C��5�u=�L�J.�r^���:qi��_f��)��@��g�b�"#��Ǽu�P�QC�<6�}�MUҵ�>�(�Z#0���2rcf��V�~]VKw�<�#�&�oaTL���:����4����:�˫Pը�[hd��C�c�	��=��E�Uk}l�Z�\�9ܫ(�6Ŧ��"ܕ��n]gn�ǂ�x��l͈'���I�����C�������|�s��,�ن���n['h)�]��'}b*�����g�ŇB+^��ǰ=|�q2�W���<_۩�U/��&;�}��R��rn{��v����⊯�y��:���\�/n.$���*nh0����42��η�y����ӵ*�I���4�O{�c�x�ۃ����;G�����֥�n;�'y�*��榟�9�,\��޽��;3�}�:N�	��ne�;�6[;}A�a��ӯM�1��=7 z�>�Gd��h�>9���(xJ��Q7��O��ڷ��t�l&��x�n���ݍ>���(�{��.��}볞�`W|1��AVս,Ye�Z֋���ͭïL���D����]8��zr������H��Öz��im8����@�yF�%l��s��z�F�ߊW���� �s����=��T~"h�=D�G�o�뚎��Lw��ܝ���u���@�F�f�c�z��]X���B�b��y�Z��z�$�m�N����z�cq��W_�{{����~��Χ�ăIC�{�ټ�F�ԅ�ͬ}Ïw�"���ξ��˅��g<���gt�� \�6������h���`�r��7����``5�G��)��߇D{��<���#��)'���|���\�"��߷�bEo)[85�N��#�<}�e����w� ��J���oX˺V�77��3����mw��}�ٽ8�R��e��@��1zm�۷͖��˲��(H�wz�>��P�9i]�=� ���;t�r7�8�KH����;޺�������AI������zu�;}�U���@u����$[wnv��\�t��뽠����k�ynݜ� �m{����t��o[W �6Hj0�/��v91B4 ��۞n�v&�q�vH}���H �p|�zo�p�����2e+^�᝵ВH��&x���k^�tj���*�*�hg�Chc�g�_��|1f�ؽ����T]m����n�e�R�2(-z����z6��!����x����z�c]px�g�G�x<��>K�`_�q������`�6ߍ�ן��Wυ�~Q��j������֌�7#�.���kw=��#�Um�Y�!����k�3����:�L��vڶ�7.;k̎�����nMn9�'����g�����Ɏ��������w�s��8��h��+�x�ϫ�\��:3v琷�M�n���ܦnϙ��v.:Ս��q�e����nw��(��u�:;r�ͱ�6s���pt��9��7>��uv�ݞ��uˮ�%�����uӹ:y5�/n�����.�y݆�[v�����볶��)�/f�����&�rk)�<�ܛ�=l��źwQWY}���ÌV�Ik�f�}����j^�[��1�̇;/f��ʝb�9��.ַ����pO�/6N�;t��덆�ԝ��i��׊�E��ș�<�s��M�ԅD�m9���1v:�-<�n�z�Ne�5�"Cݳ�nyqke�4p{�;��*��C���`�nx��谩O=\��M�\���/c�;m�����u�9���q���Y��)�@�蹨{sŞ��'�я]�:)��e6�1���m7-]��(�n��m�nx��[�coIَ�<��a��k-��v=��1�ӹ��À����m8�o\�����هP<�u��]W'����8�u�\�0��]tj�OmAWc�N@q���k^�:�8N�|)�c`�ݪ�nŇ�g��q�X�l���;s�b�Oug�Ǵu��ۛ���k�v��F��W�(��q�q���j�3v`pf����r������r�]�nC���]s�j�m4𝇈�L�����=۶Í�dA��=�&Խ=��k��Qu�As-!_��.�u���OXe�&�v��Y��+n<b� �;ק{B���k��d{qvE�s���'����DS�����1���z6j��n!�;��Vݷ)�vw�(r�ftr���qL�u4pn�\ts�
��ps�
Ϻv��k���f��a�Gm��cvw@�=:ݨ޹]u˛:@�ft���t���=�oG����l�j��q���`��6�w[5�\�<�^5�Mxn����n�Z�֎�c�&�\���m�L��CL�{��Gv�s̴�/Y�]�T�v�疏;���4U�q-^sq��yvܜbŖ�T��]egu\�0�(����xH�����ټn�k��烝՗��ּU�cGm�\����A/Oe<N�qf�n�sV{�N���.�l��'I�<'�N}b�&��7kl3�VG��ѱvݟ]����=+ԝa��lXN�\�F���M=�ݔ��;�i.g��\��t�:cJ�')�Q��Mk�G��Ε�9��6��ֆ�)�or�Q\�[�Z�e���.��=��-�-:�;s�m�	�:��ְ�x;q��
α�y�;;��w����7�Wl��v7&:��^ז1��c���݊�3ъ�3ӎm����ˎ{����X�,��;�;۝7	qtF�<Ŷ�eݺR뎂��tY1�-\og�e�$�c�����ǋ1�H��:�.u7���91�豨-z�8+�����H޹%�=O3���qv͹ܤ�m�Rl�2�B랥+w7]IMu�q)���z3�h�� ��\��\�މ���w�]U٠��''tN�Qkg��Sp�M���;/h!�:ݺ��l+�W^uӓ��1wB:����@�^���++P�q�{����;��W`�$�ΓS-��[�;n5�u�6w������lv`��8LG�=�[����
�&�=����;>�;O�n6�f���[v���U�vݚ1۩��Y}	��f{:��sǎW���܅�p�D[�v��9�5Yݴnk��X�M۞K#��ؐL<s��A��;in�#nO9���Y����sT���۬0G���ض��� ���.�t]�r�&ܜ��<q�یT]8��&us\�[I.�.��=� :��cr��W<�r뮺{5�7,�"� �2ڜ*�D�-��r,��j�㴨n�q�j�Z��G�z���N���`�r-;Ѯ�����v�۪�3�dݗ6�2��!��k�ʎ՚.7��}d������b���X�lk�;u��p���'�|���\+��wm���1��a�V�I��W�ېz�Ҽ�-���#籢-g�@N�u��f�vMmSuڍ�qJ�Y�m��k��!��hs*�ܠx�I^�R��C׵��R�]�g��Хi6��Սx�n�P�a�&��@�+l�k��n�vr\<o`{f�C�'э�x�c���W�^�<v�έ�7�y]WFx���v���v��١��"1(�v���w�C+��0�����3�%��;gm�t5�-��sVg����f�+:�=�G���=s�j{Fu����<u�-�koI��;v�.�e�{^��ݞLv�9�乺nB�p�x�����Y��9�0v|�ú޳ܐv.�^N|�Е��آ�q��2�p�glN{z�WfUL��|&��&o;%�uy񛹼��ٷ6�u�S�\gmb��[{n,�q��G�c%����u��c��q���K�#N�SknSu�]���.B�=mWc�����wƱ1��i-lF��9�tk/�����v+��Pn6:�у/)v�8�Y��w	&��C�ll졸qU�tnc7�=�Ō'.�u5�6Vу��Br�/^n��p�i�;�t�0Z�y睃Yy�<C[�h�r������j�v���9�b��v�v�|<���{V玦c�^'����w8����y�7M��R0�:0sg6��u���Nk��wm.�����u��OR3ԗm�X�����`��[$tn_nnG���x��l���u&�������Gn���{��SI�n�Ɖ���ɦ�76���'����1"��ݎ �]ǭ�b�ܓd1�e=69Ō탗�n.����{���Hsϔ��{p9P��ԢP1�'�y1�u��`iɉn���W;X��;۞qepr]��{u�K�*�xu�m���㖗'W����������/]�۱7h��z($�q��a���u�i7*�r��gx�V����P{/�Z�n[m��U۷D�;
��k������U�q�u�Fu����k��t/��WDpON�;��m�<�������l��]ܽ;v�n]ŭ�s;�lu�ݦ��7��jx]ѽ���Lzݹ���n�7��]�#]fv�v�{:�]� �:��42����	����!6FfHn�Ә4��]ح�����`���ۋK>{WH��F��g�Zw�y*��|� �9�v�5!�㵷'�x�!�>6��<&�����]O���v�'\u���ʽ'nػ7A7)����c�9-x��Q�ro6KNXLM����ǌmE�;�ۂ���d��vPq�x��������%x9����ї�u�����nʠu�Ntm�ch�Kc�љ�N���X:Cu�׷lX����{]sr�y�<-m�g׍^�1��]m�p�mz$7��w.�� ��L��x��^�0�<>�qk�ݚ�ם���r��9F0��@x*��\���#�q��s�긷(��Q݁R�m��剎�k��'2u�����`��<��&ۜWr�>3�C�����۩����W�ǒ�Ց�XB��AȖQ������lu��<��<zK�D/Gf�\1vH��"�[�u��rh�]Ak�"M]���]��Q�1���7k��*��v�{d�3-׳ف�ik���"�]���4kΞ�����3��v7>krk���F���8{{c��V�0ݺ|=���u�وh"�Vў�یH��f�۫����Z<4g�ٮcm�;b�84G-������ےΰ�:^P(�v��g�n�d���u��*��Ŏ�P�܊U��7pwk��J�c���E�)�jۥ�O[u��v�c/�0m��z�Mg���;<��^�;v�v�m���w4[�4��r�뫑���eSr�3ͱ$v�;���cgv����=v���n�d��!��n�I懓q��ٝ�=��#zQ�>2�hA��Su�]�<�nɗ����)=wӗ�����]���vh�n��:ÄB�4��O�v�����Y����8܋rct����<:v��۶OO^ط�c���LU�WS��2�s�nv�ps�k��	x:3���BAD�6�ы*��>^-۞�{�pv�x�C�5hk����:��ۯ��܋���d�͜#�������Q�,��ܶ���l��I�M�����ƺ�l��k;�y6S���q;�/��/���gj9֥�t�v�ks�8N;8-Tv�E�������t��WB��C�,�pK�ã�YNx9��ű8��j��O\�m`j�n��m�]����scm��8��8w<��'�<OOj��/n��uru��P�rn�gu�FB�ۭۘƹ�]6��n;\�$-.���q�]�-�R���.5���4��tm����\	�P{r'&�њ�p�ey�rz�<�Gy�˓���z��`����
��'��qv@�q��s��^/�2�2�"r��OC�nx�^ٍ���؊Fy�յ�x���^y�-8�m��a�E==2���y�m\�=F�[;��V��u]3c;���mr,�ݐ��zoQbmҼ������&�Y;��%T�<�mmwm��Qv��Wk�� v�5�Ƨ��@z�0�����!�<�:��Zz.��!c�Iך�lݭ:���j�"��՝���\[�\�l��q��h�����Q�Wm���Ӫ;j��Vl������깢sU���;X�(��e�T�=e3�nN�Zz���%̓�s;p7c�`1&����su�ѷik��Y7::�R�s�#N�v �7E�Igl�u����뮮Oj��u퇱Ofq4t�{U�pŮ:����^;��(�
4C�Zhh�r.p���i[J�J��6�����<̹jx�����L���	^d��T�º�F�u0��QUg�9<s�*rىXEeDIH��S�@�jF��TD�IX�RG�����,4����e��*�bVlHNK0�CVV
))�3,�E4U"MMa��R�	�Ð�B�)#,.Edn<�2Zi	��RZJ&�]�y%��"s��ZJb�rR�%�¼��s+qT��3KZ�O-g�:����e�U�%J�J�DB�JI��s�]Ƒ�`�%h���������DJ��-R5�`�"͑��U̃3,KH�R��m!d��I^0���˔�Z�LEP�9!��Qv�YJ��BЪ�Z�A"�HE"W:D�JZJHFE�1�8z6�?/�[�|e���JNٵ�x.q9�#6�m���nط>8��p����9�Q�n��;��{�����F>�)�6읶^.L���^��^:��Dm�4%/�҆��Z�nS��c=�6�a
�z<�wa�T�gr���v��S7m�Y�!ݡ������;��	��8�n.5'nڝ������,�[b�N���w\��9��z^�mNy1�z��h�S�[;=��Hzn��l[g��w9m�Q�i<���ĭ�8��OgES��뾈 �G�X��'"��܅��hv�v��#=��x�C�㮠
�n���j�� �o9���9^<N.x�Y�o6x���:�݋����p�猺܏�\�S���'�q�9�m�[e5�7�&]�9W�'��<ִ�a燵����x;]Z�{cF�!{PK��n��
fˍgxx=���]��w�`��b�v���o)���;=d�]�QA�m�����W�N��bݛs�7R޺��;�&<�#$�3����6,'q��C���<�[��^M�9x�k���nb�{N�����[�]u�N�V��}q[=���Y	M��<chx�u�e�2^���=�yI��ʛ��n���r=ǲ���d��z͞w���8�b��xKn�h�\�epXϳ���;;p��)���Lp�k�ez.����ʸ��9�nw,��}X�Fs��j>��^T�3��LӷN�y��Vw\b�d�����k�{m۹��6�C�c�y�7o)���=O��흋��S�T�m��ll��q�#P��<��]�7�P�zu���ՔN�]�3r�wnt��"���������km�:�m\n9�pn;x�w�]�.;:��^�C��Fz�������K�Cy�^mc`��NϷ>=n5�a�3��g�Js�#�=�l�9Ӧ�Y�0n][�{oc��ݬ���^ݞlc�g�ӕ��o]��9��:�;Y������{�g��ݑ�۞S�v�W'a�8��l�d0���q�n�'m��xv�.G�q�&6��݄9(;��n���<��q���`�q���p;�p�=���!��L��%ǐ���7�(&�Wo;��0q�v6܉���a�3�G�>��q�������8�r�nx3��	��y�M��;8�;�3���l�6��{	���<y�����o��� �$R��[��I�n�'��k"��5;�_h�|�I����a.J@�""|�׌����Ř�]��-��k��͒O���H&vE��܌(q�j{�����2��&L�	mF��><r�����ʞ����$���A'�P�jֲ`) �ȑ@�m���&�z���6ﮘ$����3������?����v`��+�&�-�k%M3�++�	���BEP�\v�~'ă�w+��ͫ��{�p�f�8o�� \ۭ�l8'�ve���^!�X�m��g�4�Q^F�^�#�Ȁb%$��v����I�s���V�"qD��v��Y'L�P��hl%L#0	�!��9��w�F������͉���*���s|���S��;;���˰�c}���n�ƼܹM��"��
ؙ�;%��lU�v<V�a�7뿰 O���n��~$��j���s�@7ZK�Q�Q��׍ݡ$��l��Ƅ�s�QL�Qљw`�A�9�>#����>��;L�"I�1Y]λ(ҧTnQ���A6k�zO� ��l@'��{�V9��[X �طȽ�`,H�a(�m�d�{��ɵM���MY$J���n���I׼߁2�V�(G�Om�D�>5�Z�1o�U.+m�;�:�;�����3��\��P��~~9�̺tReN񳗕� �� �H�����TW.RP��O\��]^��`F�!h���Q"���d��[�L���H��x�����b)C�W\G��'�C`�*L	�L)MNua��L����i��1;K:.b����t��Ν�~� �z���)Hש="g<��[��b.\$W]N�loVCa˹�ƍ�/Km���pk^Gx�v���Aټ�$�����"}f���v�d�=y�6�w5�2F�oS'Āp���&�TBΝ�A���`��|�	��I2f Kkg�� 3�S��;�+6����R�s`�n��0��D�P�ٌ�֩-�i/p�_{�<���m0l�+s���u��k�]�r��݌]+p	)3]��T0d��v�� ���0H$��w"��7�:/;y�d����9�1
LJ�2��9yR@7�y�teI��`�F^w6I'�T�Cs�=Q;&{]@!X��2'�[���;�� �ZPU[s.rz�6�$���`�ܡ$C`�(L	@�R�Χ�iէ�2�l[��~$�3��	ͫ簎U�y���sm6r�E�H��=�a\�x\o^mOp8�[|}�.�����+�Z��v �k�<�UB��w{j����c�y͑�01!	DD� �xэآN�^0���j:&�`ü�d���w*A'6������g羇p ~���J/��v[�2=���ۜ]�i�n���Z�%�1y����}��|��շ0Fb���q�L�P�I>�|�#��5~4����['��ٞȣVもf�"�"�;�v��ѨT��u}W�:g�(�m_6D�����37��7<N��*�i-�ԃ���c �~��v�zK$�f��|H��w Q9�|Á�!#�QI��47[�=z���� �l�]	>�'��h2E��9�7o.�;�N۠$��a`�T� �R���r����k��<(at0����E-��$��x�$.�y��Η3�=d7<�4k���=�<�^�����4oū_��,�=i�]��UC��l�.��2T&�6��ld,�Jۥ-B�Ǡ'o�~�E�����y�nS*��G^�<��m���9���v��z�Ε���i��C� �x{K�#��&^�����]:+�c�8�-�=�ZR�;ؗ=�(�F3�aq���n����X�v�N�/�]h{<>�ͤ�:�I���G���]{�GVMi�q�nx���01�rk�ַN7]�d�Ipn��lv�	s�7Z��e�kc#���5u9|��f��7g���{sp�F��[���>5�#,oL;c�?~�wρt���4rz��Nk�a�A���`�#���N�Y���+���޶<m��&J$ɘ�4�w[~����o�VX�gn�Io;�`�H����H5AL�R��f�0�wBH5��P�0d��㽷l2H;{�LA%ި���Nga��{OĒ.�y�O��*��eDC`�{��q�U���ANv� �	{��$�:�9Qz�ڹhh'�oĈ2
�e��Cv�6O� �ב9=�*+��ݍ�O��y�I8u�I����L�'C��"�p<wn�:w55c���\׌=���{IƳ�1�0L�����RIJFp-�e0F_wPd�qkȯ7�c��s�� �u��d�܌f�0�DO�ѣ��2�\V-�G�o`��ӹM�~��@K�}_��{=�9�g���V��fW��7�|C�9I��]Jm^۫�s܈��ղ6�݋�4H�d�7|ψ>�����^T�AS����d��x�}�$�Q&P��4�w[d���P�A����c��17����I����'����B&��%"E����9G���P92�2A$����D��|�
��^F�@	�tɟ��W�A�e�II��pfc�n�c��w.(2���l�O�yS�/s�mD��l=�2QM���SsG�V('���^�A�=d��]�䣶@���{$�H)����>a�Ny	'9�6jm)�!�۫��$�g^P���$����Q�L�Y�̞��s���^��^@��}LM�ܮ[� ������f�0�DH�
h=;BO����� �.��/ޘM��Ḧ́pk�#���{x{{+Nh�]{%ܛ�A[ڔ����/�wC�`�<(�zw�;:#�؍\�eME��-E����OĂA�� P'�]|�>�{� �Q&P��--�U��1�Q 1.���^�I7y��L���r�A%��BI���&$T��H�{5�d��ޠ[�n�c	��(��׍��/3��c�Tq�[�!$����t?V�+�p�1N�g]k���m���q,x���댼�����Q���&f"(3WI$���I"�;�%��o�� k2�	���"l��FR@�HD����?ks:�ɡ;�M��$���������a�����%�ԑq�,J�L$���.^u0I���d�j����q�]�[zy�q$���� �/3y�H�b�d#	DL�0���ӵ'J���[�H5.�	7��Oď�B��yw��3Q�R2fj�l�Ec��G^�ѽ���v�؉0�AF�x��:�f�i �6'7��z��Xኩ�	I�fP̭�gCJ�����d����RO0�4������$����r��pвiQ���d�fo6}��*v
55Ox���0\z�G)�[�ɗ��u��8�!�ۛ���=���[�u����GA3"��"Gx��l0A���`H8z�(Z�s18a���m�I���Sp��J1*
����5��M�WS�J��b�C �M�w6H$=y^	�p�f�<ɥ9�Td�x�@��1%ĄH�ӯ�$�;yBH$���Q3T�)߈9���'��T��Z$��I�L��n�����N��r2l������'��1e�P�|��w�|刏OJ�6�I���H�	�(F�N�7��qMVB�u7� H�� �t��
�#5�6c}DRu�KH'Gt����m.���Ux��G���$�2��NNSTל�O)��=[M7uc5ȷ���&хN(��m-���8�'{�ʣ0(ą"B�)2I!�ۣ��p}}�kG:\8�ԝ9x�;Z��ֺm�^��On�N7��;�iLc���g��n|Q��O4���W��d��>�1����R������x�ul�ƭ�������t��v�-��n2O[�G���=X:���c�9�u��G5�n܌\��Q�ky4���1WM��ƣ����)�w[��9�g�������p�����S��O�vh=�����=���c�~��Rx1��8�bb��&`�q�0��|��l���-tG�[d��ה$�Sp��
BR�"����D#Vfȡ�-�d�ӝ��A:��(�3��d�=|O�>����!2�m����OU@���$�����=����9�I'�^@�Fs�l�Ӧ"�A��A6u�{�IV�TI8H0r�$w��0I7���{�����V��imЕ��8I2��$��i�[���$��u?[����<�ucȯ	��A7���#Ywٳ?���{g$0㵹�ݰC>8�Fnՙ���%q�+[�ջc�w8w`n/������ŵD�$�g	 w]�d��ަQ�2z�ɘ��ک�� ����Re	���t��Kv����n��y�T���V�tx�cy���CGp��٭�����ԟPFi��:�����շwK�ݽ٦�lZ������	����$��l�v�N<�e���IU�p�""BR�vm<� ��ަ	'Ʋ��C��r����$����>$��l�ȯؙ	�l��l���w�/ݣ1�l�w7z�$p�\�8zoL�C�OM��_�K �3���߀��Q��a��hM;�"��[$���oĒp����`�/��.g
A�,i&�8�K�6�v�V���j�x^���n�����z������	F�/���I���`��b�Ȣ�H���B�]�y�l�F�o6j�X���2&`(��NВ�����/r�-�a��f�`�A�Ր(
���=�fvS@ S������>�ܩ �^���1WF�!�]�*���TOL�{%sm�o?f�g��Dfq;oX�s�c=�^�,{�w�c�=5x�=\Ǹ`{IZ�#^�j�L��=��f�/!��<p{��)Of�P>�Mo'�-�s�׀�r)���v�e���6((�j�=C3cPܹ���cvqn
;}�.�������+%�s��A�On_-*"��Wv.�&C>�ۛ�n����aS��Bv��M�$~��q?x���2RM�oOt����?�{�C�Ͼw�wپ_�ܻm�[��~����'5l����{�U���J=��5�q�(Ƭ>��Ɂ��g�(M�X��ΐ��q���㇢�[�N 7Go'8O+lw�}3r�_�]��
��^�f�� �bwe�Ys��S�zX���:�P���Vݛ����*c��'�Gc���J�_-;����� �9M�[������SΡM������C۷����LD�:�9�[�yn�&Oj�d���e��4u��:��2�����yt^u;a����u�9�y�.�SͻZ3q�r�ߪ*�����a�Pa�����6����B1���5��;vI�r��h[i%/!巟.�c���g`Z��~;ᮑ��6F��Χ71ee8����
Sf�+��iJ���Z=�@跴SvxN��`5��b��{qzb�	q���&�zv��[/�׺Nty�>r{fz����s�8B��d^.w{�̓l����l�!��j+ʑn�3z<{�y���e��U9|7Ƕ����{s�����A+�Ya\�S23��`h�"�J�ܡ�;�EDj��Ҭ��;�g�AW����E!fQf��"E"�Z�fG�+��)VU�f�MIB�^R�d�Áɨ�u���J���HG"�H�RY̋
�Z�p��$�AeW*\�8DٙȬ��4H�%$�E"�P�S��DFYfQ�jI�EBR��R�J�A�Z\ҩH�Q5DU.�.�^r��K �"�Idl�8q���Uj��F�兔"T�j�iU�L-�jqP�B�T���IR�Z#5�Er�(����F��rښ"YU1+�$��ͬ�ȭJ�
��1".h�-S҈�e&TD�TabRTQb�*[H̱�hT�D�Xg,͕�aeZ�3��I��.X`V�
$"%,�������� [}�L ������0�E4�!Q��]��s{.�V��n���>յ�D]u�����@ܨ� n�����q2H��.A�Ku�v��x]E�1S�Ӥ������NW_6�����UPR�L0�AJ��oh�^�������HC�q�n��b���=�{����ʉP��s���O��Օ�$�O����]�uA�6{��u����r��p�dRu�4I�$"d�!1J��2X�2�l�����O�udz����Gw�뼵j�d��Z،	p���H�ќ$����~d��o�Qծc�f��l�ʐI]��7A�)�`��eD̆�7�흭��YFyh$5���ܦH&�;�W$o5Ρ���Ǯ������e�zvy=���Nn���߆���{���n~=��l7}=��s�մ��Y
�� M��;Ǳ��M�-����ק�x�v�z�*2����4%U�@�O�Vn6<I7y�F��Y�%��llY�.�n`�����m ������.T����z����R ޵�!4�m�����[�` �gcdE�w6!l��^���Ӿ6n���z�r�>�3��H >"�ݧ͒mI�$�J�ݗ�RI �:���H$]�s`�00iyɽ�o����IY\c��!!%		�5�|I����IG���
���u�~"�;�+ ��xBe<E�N����P��X}���7��I�_o6H$<�<�f���ڪ�&�;�(�*$�P[�{d�8�%<N��u�]2I��w6	� ��2�}ې�)�)D�9��5����	˳wҼ��ZF9�׹޷�R:D;��F80	=s��^{1���;Z\5yIH�P�tB�*`�`J$>B'qS�^j;rs�J���n!��]mlnn1c7������n:�z��=J.�'�6��(k����,�kG\�c�2<�d�Z�-�"][59��Ź�
eJ㇎u��^rk)�킻����lw/h)�V�ѭP񴽴��j�nx7d�塓���I�[60v'�1��c���}�i��`�-ۮ0��u;����6��ݹ�N7�^�d�ݷ��Mם�{B����sc�bu�l�������$%D"x����'�ow��|H���E���
�L��و6���͒	}����G�*b L�R��[�$��6T��*֖�� �w�͟i�>�n�*�7����_�|�"�#�Wm>lO�yR	�*�?,�Y���s�����l�N�y^��l�$"d�!S ���vQ0r`WoD�
��2|I8��P�����R��x�1¹�6Ll��Ĩ�bAS@���H�}���ȇ�X&��7�H� W�#)�6��Upzիc$&� g�2��((�Z�=qFC���K�X�g���ηY��͹+������`��T�P_8���H$8�����L�[40R��*�;a�l��D*��LI�"J�*D�;��� ��y{�P��l�۬�͑=~��ȟ��\�ȁ^��/�uۥ��I�9xٺ�K@�G��R7�]\O�n�e��M�E��3�.�}�I$��@#)��~$7��.�}�~��g��U��-%��\�<7r��	9O9�I$G,��ד��x��$�8�2���	�a��Q0%)DO�V�|�j�&ə$�d�mI�$u�~$�w��s�P��U��;D�c6����ff	�(HM�9�A���e��ۣ\̉i��O�u�d����"$�9�2���J�В#A��!��m</T���[�mE���ɭ�a�f.;D�����w��1$�H�q�$V�6|I7y�ٳsQ<����s��VXg:�A���l���B�
�"��s���u��u��X�ѽ���H����7��I�}�R���vF6�E��/���,�|H;{�L�A����\uv���7"�{�f��vY��u��§Sӣzf�0�Rr�U���ޔ��cET�{���`�Ы�(��QSV;Y���1���xz�&�|OW^�����2F��Q�$��X���~�x���M��4 ��ld�:�H���2�je�b�Uu��GJ��1
�D!��|߉'�VP��j�H�S�~'r��'ǯ;��O�۸��^&+��4cP� �RÃ�u���t-1Rz�k �yn��=�w)Ƹ�?�ɔJB&Jqn{$e�u2I$S�s�\�q�Wb�3������6�y�H���X3�3J�T�4cv�$ƃq�ܷ�N�m^�� �M�o0�	8gr��{`������>��O6o&PP��FQ�M���$��s(I�'�S̭{t]nv?��8����}���n��:v�>]v׀� uk����
J�JC@��}״v���ܽ��O�><Q�/�~���0�F&�	�u�`��D	 @�o�>�}�ëD^����ԎC����V�x���y<���m�}}�s���<t<�C�k���;[XY�I�".��y��z�G'�����B�*��<�{��{�n����w���aq�������>_/�8p����v�_�����&�h #��m>��}���u�]���Y�?����h��	���u��Q�G�>��l �z6���_]�,����j-�����8gSB]UI�x�P."���pl��v�}��?~Y��2�����������v���v����:>�t��L.#�~���v�\{���?���ߺ�&�O�~��Gi�۷Nӧ˯�u�����.��D�be#!1dx�����>x�<>�5Dƨ#��� 7{��#��#g��u�p|O��$�:ߟ�^}`�ȏ@���vd}��5[�@�<���z�>�3$�?
&���tÎ�Bi	��~��GyݻN�,�8~������ο|��z�z��I�3���u�ΰ}�0�18��mx3g�"�;9�((*T�ELC�@>��2'L.<d}9�hO���G��ȴ����ۤ�qw��<���v8�Y�Dy���#��M�*�G~r/@��?:L/˯�u�ܝ X����O�Ϗ/��W����I��=����{pC&"�v�}Aߐ�_uZ�RJ���g������>'�@�'I��|�v�ݤ��v��ǈ�>����~] ��tٿ�Â���uu��Vkq(8wP�|�a�7I-5҆�ٝY3�]J��j�,�׮��Q���e����g����r�lmc8(��tn]�-���/�l�m٦;`x�!������ukǨ�h]�ӧ=���>+PtٲbqڠdYI���>9㛐��WIm�l=��\�����2��wb1x�ǲ���yM��ÖϞ��k��ֲo/Nڎ5cv��!��Q;k�����q=��|�m�{;�1yތ[�w+tfu�8��������iرە�o>��뾬���%πft�q��	pkr���usn�<ރ;�^�У��J�&���[{@0q�i	0��=�wn��0�Y���Y���u���*��Q�O�z���`��ן����&�ν�s�&�?9��>�ߺ���Gi�����u�]��Y�q��X>�i&�u�u��;q&���?{��n��:v���:���z��y�?n����'Hϟ�_�s�%g��/��v��N;����c냱��{�G����0%�nf�'�E��O�H�@�@�Oz��c���󴅐�����v�y4��y�������7�t���|��A�ѳ�S�G�#��N=���t�d�/�<��Ӵ�pL�����=��_�z����b���W�� �W1y��

�fIS��������Ӵ	��&�מt}v�
���ʏ��燤�dy�˯|/��q&���?{��n�'ht�9U�׀� �t{�D\R��� dB<��c���v�s�A�kZ�gv;Uۮ���47R&!)���bBRTBR>G�>{;�\����y�ޏ����0���_�� G�Ǻ-O�TX�s���}w���v�����}���N/β�bT�(B���g���G����QDG���X~��rj1M��W��cB�c4緎��$��v淳�TĨ��o��e��^��8�o����q�N��/�\1O��w�=}w�BO�����<����]�:L(�������8&���N����ϩ�f*�aK���8������Ti��Q&�>s��
}M�����v��N��&˯|��;t�&��i������O���{��8��8�By矽��7y	�;N��|�o��ϝ�y���(�"Q�S@B>7�P[�]Tn���>�����}���������W����H�'�'���g�'|��<t����}v���ן�;C�ӈ����'g���>�o�����~�?~�>��4!&���:;wnߺ���>|������~����;@�'�0�]y�X>&��,u�u����?����~�?���_�A���KX�tCv�qn��&�q��.=���.v�k��v>�����ɉ,k?�i�n�u����]�v��^y��ۤ!4�\G�_���;qۉ�_�u�矹����:��o��I����:��t�ם�?��7+���GHrN?y��a�e�V�����z� +��b10���|����$�:O������Dx]u}�TF�� ��CH?�N/�>�s��x���>q������yߝ�&��Y	ǝy����t@�3��w!���T���y.gn6��e������ww��z=����](���C��uyUo���=S�u�\���w��{��$��0�]{�X>�h�X�����v����|�����FD�����$0G��>�dj���|K��ϝs߷� �0��i���ۤ!4��q����u��;q8���?{��=y�9[C�Ndx�Q�2��^��@��虙$2�LY�8}��g�/G�H���Pdx���6{��6��+����C#>��$� "�'���c���aBC�����v�O��oM��~&�$a&a@ʃ`��0� �u���:�';������n��p��q��;�wμ��o�{��{�O��~�\t�BMN?u��:;wn��I?��~���i8:�'���~�����u�ް~�0��^Vvׅ��"��ΘAA
`�n\����7=�����'NӺ?�_�~�s���������;v�	4�\_�{��v�S
n�����ގ��c�n�?�u����3j���@]#�&bAP�BR(Q�$������vi�1P����G��<�|;�]�+��죲����?�	�Oz��α�aw`�!!����z;C�4����s��/�>W#��?>�>����n�ߝ�ʍ�G����!8������L(H�����v��L.g���:�ϝ�Ls��/�*�8����Z�c<P�z>������-ڛh<Jj�F����DD�p�B6�Z-�rv����n��;l���|Sf��i��� z��C� �3�߿��i��u��|xO��>p�}��{����S�@�gi�;O�^���t{�]��_�����|���;q�q8�i?y�ގ�w���t�_�|�o�� S�\�c>=����!2���N�Ov��[�Z9T��s[ƹ^��������9����s�ϕ^���}���z��&-@~�ޏ����I���׾}�I ����F�����W��~��;wnӬ�!d<�����ؚq\����q�σ|�:L/W�?t�:G����쟺"��q���v� BH����~��v��g�8�{^���+�x)�ϟ�Y���ቅ��~{���"�|�'�r���i�����h�iӴ����G�ۤ$�aq���y���~��>��n=�$�����v�]�&���m�:@���=�T�J�JC@�|;s�0v_ѕs���0�?P���}{�Q��<�����@�|���>��^u����iݎ���<��;N?|�������ϗ9�Ϗα�0��~��<t�SB�>��Ύ�v���~�<����q0�G>{ߟN�;pC8!�/;���<^��k�͟ � n/�'�y�.�=�۾_S��n����|���}��s$���4���3'���ܸ;
��3��䳶��J�Mn���h����٪����uutzgf�1�p\���#����M)�'Wq(͚��,�ɸ÷��bؼs�K��y�:�d^��-��ܠ�Ԙ���s��mܛ�	yf��cH���:��B�]M��Ƒ�qVӬ��8�o�t�w5�� ��y�9c�,�t{�/7�KHF��ӗ*Bh[�⩦n���6����*QJ��[q�{^��7��5M��xu���կ5y̼V<���M�t�o)�s�1F��3�BĽj��X���z��3��t�Ͻ�G�V+�>xu��8����1z�t�r[\ڽ��Y��"�݈S���swD���Z�6n�"Z~}�r���^L�|���r{/v����Ǽ���������{׆��~��`糟��b���=�����-�7n����z4<�٤��ۇ���{��=�[$�{$�n^����J��Ya��s����c���[��z�u;5m�,z]�b�$b�2�6�M�W�T/VRC�ˇ�C����kQx�:�=���_Cs�������P@e��!�w)[���X�PtV��F�hݾF�V����ʽ��=Q�/rT��saw�����^���g�F�1=wݨ<��Ҿ�<n�c	AV��.����
���V��iX�v�Ѹ�5��HӲP��;��sZu�����B-	1+QB��%3J2�T������Tu�#2�5�ZҨԎZ΅GS��r���I�DȺ��ȪTLԠ�!0�3�\CS(hDE�g ��1P���2NV��4��,P�����r
"JRd�d�r�QsU.Y�K��憲��)5UY&�eQ�FD������A"�Y��2���va�J[MJXEDr��x�W��B�fr��r�脑tD
I�b��O!�u�)D���L*�M0��IQY3�.s�i�PB*�8\C��")#D"5%,�,"�P�Jʊ�!]�T�+B��Y���5�YF[\帬P̭j*XR\�S+�&����2#�P�2�q��I�akR�Jd&��tE�s��2��b��2�iB]��IJVB�gI24QHJ��%h��Ԥ45�u���D���p��&m�׫�`�^�ֶ�Gu�!�G1ی]����<n+]rW<�]��9^r=u��`u�m�ɷz�W<<���9m��N�ѳ��ܻ��vg��������-����v;jN��K�ͮa���^6k��ܦ�:�`vmb�x�wnn�:��s�<�vv�r�ۻF6��m��^۠�赸z�<r�n#\��60�{v9�Z���)��;��kgu�mp��Ͳ���n�m7
�,��î�rU��η%��FKv��v��t�v���`��������%=&��E�n�n��eq>/=��a�;\,�{�v���Q�s�fmv٭\=�m�.Vêy�WU�;�6!d����x��F��gdCd]��I�m<8ہk�Xd�ɜ�zk���8�Q���<�7p����/��7�G[sیf��{._
b\иUe�)֣�y軭�[��:O$�G����2d|ܻ�,�ι�`y�[�M�^n��\��ջn^N:��7c�9Mܥ�oa�oq�����9�]��X�Ò��Y2�����p�gn�N�cv�'=vV�a�I��=��vU�ݓ��v]���cu��cג!p�9�p[��ӹb���s�n�/e5v-r*�јn0����`#ou���n�9��Y��q��'�Yzp;A���ek�Ꭓ��nD��H�Q������ٸ\y�מnP�C�!ٮ�b(Ƹ�Y%��;<��Q�-��Kv�{h����-���n�Z՞+���*Ow86��7)[�;c���k۠E�ެ�q`���t\=ׁ��Vݟ=[���]tLl����Ȝ�C< k��Ȼ�ىۮ���i�spGX��3��9�Z�n��^7I�0ke��A�^9��:㭑���s&��;6�*����=jէIc����e����{zN���Å�R���\e�y͋rqS�F�v�gNF.½Z.�mA
\ͫ:v�X����]n��NrM)[�dX)����-Q�WWFY?�w���l��Oi1(v��Vv�v�K`��:.�#���\m�Ł%ݱ�m��>!N`�ud^'�K��G`p��jwk�J��v��v�ufmnų�Y�]�����۶򻉺Smh�S;�������:�i7]b��:�x}p8�t�g���]7\8�8��-�O8˧���`6���7�t�ױ���z���[����\�s�U��}Q�É�p8�Go8RS&������!���[7I��<��U۶���Y.�X�#p����}����Ϝ8_��������?�@��L/������0��ﲼ��|+��(���i_�#�E��������$��:^��X> }�]���>p���ϟ���0��������fO
���2����o���A��W��L��>���S��O>��c���ϼ�}�L�P�a�߸
��B��'Ä���'g���|�}�N>�'����`���i	�����>�v�I�?���{��`�FJU�	��0�4�|(�	���~u���0�b�}��:�on	BF^tBA3HP��"���}�,�޻.�����|�Ӭ�>]��G�ۤ M!iſ���qێ�I�4���}�#ۑ��;|ӥ�z����ex9׿<��|9r���tt�\~������0� �?~��G�����_z�������~����pM�?������	$	ǟ�y�>���u��,!����v�h�>��\�ս�Œp*RTAH�R
G;<��a��M���5m��IbqUO]0v~��D|$�̅0�L��>��'�@0��
k!8�￼��wn��0�_ٿ|Ő������\
��<	������c�����;{�	�}�_>r���8p��S�������0��i�?�߿*�ȗe]ߗ&������!z�46]��Cks�8��U��h�U7�:����
�b�wx/a2u�ٙ��F��ƛ�ЭS5u�#n&�� ��{�em�����BM8����y�>��N'hO�<����n�'ht��}�����Җ�W��Q )�ߢb��*&L���;I�ߟ��u���1����}���b�8'��=>�������>'���?}���c�w��@�!!�~���;M8������Ϝ�7���}q?V����DU}����$�G� #���GyݦI?y��~��w�p@��G}��>�C~ϋʍ��G���1V<���c���=w��9���_�:���=��x�&@�?��<���z�k[d�,�#��,o�~|,�qaĚO��~�����ۧi��}��2(�$D|or���!�Pj&�Au��g�����pH�q�.�w^�t�^v�λ���Q׎�����ڧ�����+������|���A����LT��~���x�PF&pL23�~H�$vE�߷�3�d�������c�aL(v��y����|�ǟ>|>s��|>u����w�΃���z���}���9��í��;��}�|�@��?{����apL�_����!�Px.��+^A�S��]�0�+���\?��_/�|_��Å��p���w�Gi�ݻN�i���Ώ��!d�y =�21�>
�L����QG��YZY�w����݇ww��d/N�g�P�������eݦJ}�_��:�\d��{� #]���|�4�{���v!&ht�{�;��[�D�	D(�&Rb���9���]�k_G�bU�^��
#�$ ��wG����0{�X>�� I N�y׾��;r�]�߽����vw��m��s��{.\�tc����:�{��'�l�e��M��6[��(o��H�u��Ӵ���>y��O��0�<��|���%��+��t��_����o��~���-�|r��m�9^�֤Y��L�,�u��>n�~|��y��9��_�=����~��{�$��;O��<���>��!4���������;����{ߞ�>c��	�z��Gi��I��>y�;�� ��qI�1�!�#��ϳ(����s�������z>�F*13�}��Ϙ:O�B�O:��:�n��t�~w��>}�ޏ�x�q��G	11&b��/�υ��#�} ?}M!&�	ǝy��v�:@� MK쩛Q�C�O ! �>Ͽ߼���}�)�u�u���s��(�2�T��$0�_}�,�q�s���4'��ȏ[ːϼ��$M8���<�����Hy��}M����b�w�i�����2�7�LZ���b�}�kwd�~Ç��چ�UM>�v^�ʖ;�/�^��0��tm����:��|���?�� �v���Ο�����D�:�����9��O9ϟ>_+��aq�>����=������S_?o�����y����O�����X>'�	$	���α�ݎӧiC�<��Ghw�N�D��=Y���w��|�&�! �n\ґ�lt=	�).d�u�ɭ���:aŵ��������;�|�σ��:q��~����}t�SY	ǝ~�α�۱�$�y矽�v�\��������O��\�w�`��~ǂK��wk�͟ ���"	�QX>�`�������0���w?�~_|�����oz���I�	4�޽�α�0��q y����}M�������}�����W�}��q���ζ�'H�ߝ�4|���ϓ�7���Ԝ{���:Ƿ�� �������#���F%�����=WO>��`���$��O�~�αۻ�N������Ghv�q�u��z|y|�1DH��dx����+���^�q7�$Є��?}���ݦ�����}@�I���������>��~|�{���=����&����ϗɾ/�|���@����z>�x;N�i��������@��Q𺍕��{�'�=��k��ۉ�8�B{����v����:v��qe�x	 R(��MF���
�a��`C�������󑡢�ي���ʌoh��d�ͬi��n���F��1;Tm��������B�3O'vUH����  .mx.	Sm����;������{8�=͹���x-���ݵv�˷m���A]Z�%M>�'�$�H�v�����|�<�VL���l���u=�vQv�Δ��sЍ�b}����x��x�$�n�X�F�yp`m�jF���lq7v�� wi�#�[�8j�=:˻l-ͳ�]�����Զ�����n6Ch�k��z,s�����	�6ۑl�����.Ǳ�t�*n��Y���r	wK��Y�y��o���蘀d#
&eB_������Π/��d�����}�1Q��s���p|L)����Ǽ����x�D������awn���~�����E����9�*	O�>����$�G�yz�����9����ݦ$�y��~��v$����_�����a�b����~}<z��=��~��^�m�������)�.}��v&����;N�$_��~t}v�M!&�~����y=���׾��\~N,�M'���ގ�v!;@��t�_���o�t�>���_|>|�QHb����}��̮�쏄��[�^z��ο}�����F&�	���~}��0��	�'���v�߻���>�Et3Nwނ<	�3m X#��/l�D|$��!D�~|,�#����
M!&�'y׾tv;�gǿ�zx���ߩ�x����=���������_����Q��V���^��;{�	���ط\�b�U"�?1#0%*&TFc6�.n��kn�B�e�ͦ�an������~�?�	A��s�ϋ{�Orn�����`�:v�gi����G�v�M!&�G��{��v|/��蟻6}�����{�ٗBɻ�I�0������z����>s��N\���9?N�;I�����A��������dg>H���V*�iUR��2��C�!��G�i��5�@i~��>�%��9a�CݼR�A�ٝێ�(�+�r�1!��~������ ��P�	0�������>�I N�����μ,�����>� <ۿ��L��\3@�w�Ʌǡ{����<��qӏ�'��^�G&��������i�x�@e�;���V�˯��@G�&pL�w�X>�m�ߺ�α�`�=�F��)?dY��yB�o0v}���*���p>�>@yUPc�HI�!4�ߺ���v�S
~���#���F��i��� ��L'�W��@K����&e(��1Dx.=����A�ۂ̘P?y���{#^�c�
�Bޓ|<4�pLos�G�!��:��^��;wnӧiC�߿{���G�Epһ�{���� W�@^�	`�u�'��ɛi:�c�X��pl�v���:���wn&>�ȎLL���D��χ��[�@3��HI����:�Ύ�۴:@�@����z>�v���u�}�ߣ�=��?z���ۿ�u��a��~��|�^������|���ź���ߺ����b�v����?��>������Gn��HI��޿y���q&П����Gi��I���~w�{���ϧϗ���뭿'D �w퉈Q�fbb��G��wPv���LT������db��ÀGh���|���S�Y�Ǔ{�y�[�鼪��rcN����W>iX�p�`܇���"$U����f�/�۩:����9�ӯ�6����� Id	�����c�v�&,�����;C��p;gB8$	��
U�G��Z���j���h���=$G� #�y��,YP!$<��ޏ����g3�}���}ݙDQ���{�x$�}�]xY��^a��Pb	
`�1��dz���d �����>�<�m}� Eu8�Ȫ�y���!ؚq��{��}L.;q&�������ݡ;N��O����X> }?v�vwⓐ��R\P$!H�*EE >��ˢ��-����
��άg�!N��������g����aq�����������~��G��1Dbg��������K�z��~s���ϟ=���;����c�v�:v����~��Gi��g=�������Ϝ�\�|��>�<�r�g�G��f�P���=y�>8���<��ݻ@�I�����;@�'�0�����`�uh�y{�_~8��:�E2>�d�"n|��o��&���{��v N��C��}�����0���ߞ���_�|��n?����M'���{��av�Ӵ:��ߺ��'H���y��䜹���r~��v">��'�x���|Y�����Q	@~�����Ę[�>�{����Dx�F}_mxY��+�FN�ϓ#:�ʟ�`.����z��h���=���t���z�����XT�~����Y��RTjdݼ����=� �{�yB�������&�A{��/��/�s�}�N>�'���z�:MI�	ÿV��}�T��'�" A�����0�;0�_��Ө�h��}��fπD�#���Q��DD�C�2�;63�6����-�y��#cd��;uS����v?�}��B�B�2Dw�� {��2> �giӴ���y��ۤ$�i�u}����'����p*f�a����(�">�����ݡ;C�i�����[}���<��|�<�ύ����t�\~�����Qs��e`�����IP>s���p|O�B�'���v�ݧN�su���睇>���G�&�[��r8I133"
��,�Y�G��W��<�!&���:�Ύ�v��
��7&�;���0�0�|(�
:�=�Ө�h��|��:�i�y��^3$��fIU�	�=չ�#n>���*��=���þ�w�ӧi��������$ӏ��y�X���q&�����ގ�w�����?Ϟ�����Av���?�_���s�}�Ϝ�"��|�'���������Ɉ(�����z1}�]}F6:��ę��>T����O��Oߺ�α�awy�@������dy�C
�2��VC�QV-E��Q#�ג��+m
�wq�UV)�F���{���Tނ�w��I�v�k��ϔ�j�x�_��Z�`��MP������}���>lq���.ƺ7�������p��W����%Ì�.#Ы�D@9]�B��D�X������n��u�cGV\�.�+�/�s�ͳ��-�\���mp�qۮ�3��t��vۍ�;��<��y.[y#4��'fn۵�v`�zy�ᣎ��k���n��ցDր�t������;n1�UZD��j:��dKjی-h'h�9ն�fKs�v�p]l����6�h�2r�mӜnv�;]O��s�8n/������k��Ü�_�t��'�������hBq���}v�t�$�o��߽�v����S�����Ǹ��Q�9u��4b�y�׾u���nϾ��s��7�?����bn����Ӵ	Ӵ��ϯ��u߿9�6��|���n���i�{���}�n;I�4'�~����݂��|��]�ϔ�<��~R��@������s�>?8��}:@���~���:Ƿ�LT����G��F&��tW٭��n�m�ߔe,���I@��:�α���i0�d?���ގ��4���s����ϟ>n|>u��;�'���ߟ=���8������c��P�HN>}�����v�HI�ߟ��v�ؓ�� �GgW�H�j��y��S�\xx>�������c����|<�������ϟ��O�o�}�ގӱt;N��'k:�>� !�o�A���{HG��Y��qێ�aM'��~���ݡ&d�;]��(��&5u�ҭ
	0�Q;�i����]C�Z��2�UKD�����8�Aq����/�>�r|��r}?�=I�}��c�aL(�{�G�H�F&kλ_��<	�e�#:��t ��#�{u�ۻv�;HB�������_�_���s�}�N>��~����&�����pN�!��	��*�m9���,��ri��h���9��3q�������{/y�A���G#ob=�l����������w���s�0c�����}���wn�:@�@�{�{��v�ؓ���'_mx��)��v�}z�|>Nr�4���y�TDA	J�aDW�d�7}~�Ύӱt�:i}��`���@Dy��8�"����>'���߽����	�;N���y��x79�LȈ��aHb��'��2�s�h�Y���H�� �}�}�1DbL,^��ϸ:O������������~W���<���|��0���{���>|�����|�\x�_w�A����hBq����z;wn��}��]��H��{׿��N�;�8&pC/���&�b�{����c����TtmG�!�j��*#ң�L����3e�f,�^�ShяnF�H�b��qs���߿��w�s�>������ߝ�b�v�;K�~���v���HBi������n�>��"~����G�!��dn���'��y�t����������Ϝ�M��>`2h��_1K�֭Ӭ'��	�׉ ��W�?����[������x\% J�* >��tH���|I~�g.���3����^F��h���Ӳ[�Ȍ�k�L޺3��]���nX�#�K� o�oS�ܒ��Վ�}���܆5����yg,��&������<q�+�w4�����h������;�")�
(A�N�m�̭��V4^)��'�b=�>�ͽ���P.�j&b��W�KOvI�lQpV��LN�!-���vv"͕+f�����N����onkz�;y�d�fm����t��ZH�&*ޯX�����!�Dj�°=������a�Hۄ�ޫ�-m� �O|=�8o�z��I�-��I��K�4/.����RE��Os���o��2�CS50�ȉ�VN{�@�9����z4�S��W���x�i�曼G]4���#!WeԖp+��3`�|�����s%{_�+��*5����*��U�#g��+U�m���@���9n��l�q?f�K������7t�b�����wI�J��c�5�����YR�������>�w]؀k&�Yi|���B���
�xa�`��l9E,�D%�wx�]V�����ݷ��f��Se����;M9V�/��M<�rO{�����T|vS�hK���~9�by=���Mݎ������Ǟ��S�{����{Pz;hj�u �Bݤ��s�	w���P�"L�{���<|���lΥ��Q��s� ��e�-�P����KVjl��=���{዁��KBc�8�zt���=���R(�^�^��q�}}� 8.�����~��({��A�=��zpع��jL�hj��@ŇieU�T�9�Q�B����e�����S3	JS5��h�.(�@0�FLEI�ij��JaR��I����B#�(\��2�"(..DF"&\�ԃ\��\�(�jj�(��N*��R98�:,�e�Q&�#6�@R�j,�	��E�-�R�ØZ�#I$�B��Q"'*��MN�qT���
�Qd���G",�ZYږ�!�"SZ4�K�MD�LH�*�ɘ]iZ���K�`��\92�
����(��a��Tӊ�*J�RH�`�$r�䡡rT�4���
�p��X���˕H�E�,,V�bQs��$�D���
��K�G3�ATW.X��"��I$lIAǃ�r�8��H.*Fȓ5�\���r�&�U$���������QTȵq��(I"
+�Ĩ���']�-2,����;r?�`}���}�*��߲�#����X��*"=ʔaDS�{]����1��i\� L7~�A���`�y}�eF�t�uk��H���U7�L�Q&`4s�2��ݽ�`�ר��$�E�*�f�O������c���{�ߔ;�~�O/8�H>�s���ˁ��7>�4��vK�f�����_�������H��D�z�}y/�̂A7���B1����Վ:�1���P$�U����ƓO�7m�eZN��.;��s`�ھ�	��[���x�����C��2�F�17��f�A&��i�	��<�nL�1iuN�	ޛ��7���7G�R��S@Q�D�gp��q�86&{��3;��O���%rprټ��b\�����W|�Icwn�ܞ|c�'��j+������=6�zu����`z[n�ĆW߮��.��p�,��QHȝ�E�+��[�� 
��m���|��*"=��aD6��$GU�T��T}��/��A���$��c�����~�:$��q!�����q��ՃO�2u��m����� ��wnu���S߿7����]!0dO {�2�'s�i�H �آkv����Y���w��'��t�
fbD%�7�BC��V�mZ��{u�}���I �ڐK]�v�}[�N�m�A����
D�LH(WO=l@8n����StwzE��)�� ���l�I�u�&o�L�^B�Doź��/_oOE4��ăѵ�� �آI۞�.�E����p�]6�&���)��d�Jh���� `��l�@�3��1�������$�N����\�P�jh�Ίވs�R�ڟϵ�����i���i�z���F��~�v.�}�>�Ş�3ǥ^��M+nTF;ڪS�-������Б�����N�\tna69]����������Es6�.���oz�\=�#y$6f�ѴY|�b��v'Ń�lg;rX	gE\��:�۞�;��ݳ	����ݏlv�yְ�6�n�k�/b�Ggm��]��\�m�Y�z���f�ۨ������K�m�����`M۶��]�X���mбƴ\��	�nJ3m����j{Nq'��}E�q�j��t�+՘�#�,q�W�$A�p_w��@BD�Q�>���'�m�M	s��ʨ��������VI>#n�����1$L!LG�/d���n�#�{�]6�� �n�E��O��ɾ6���y{�䛈�D�ʑD�l����	 ���� �W5Yn��A����_�>#.��(O���6	1��!H�12!
ާ��:&F�U���X$�5B���Ν�d3{���@��Z�.�P���߷
T����l�]��M�v�Kw+)I+Ƴg $�N�2|Nov�3wKtӼ�s߻�'9�{B9Y�m�-�D�#.[�[�����Ӈp�[X۞??>;���g�M��:�v�@;���';�hv��sd-�>��@���s��¢#Љ�"E?7�l0sƃ��u�VqV��b.rV�r�����/9������r}sCk��c�gv�棿/.F�#=J������
�j�k���ė���z��ޣ�>��	9�v�$��3=U�Sa�V��J˙�R�!LJ23�� �$���H�u�#*=��N�h|K��lA�����Gz&&L�*&K`��������j I���D�v�6��.ޭ[�X�&o��	�\߈����
D���Ws�oĂ|�{'(0�1��/+s�2@9��LH����6Sչ���R
�['f�S�����zN�:&g�������䫰N���r�*m��(�*`�R#8�W�2	�s�2	����D��/n�b�XV��	ξ��$��a)��"L#4Ed�׊
|��
������$�^�d��.�hP �8�3"�0,ޤ�lv�waQ�D̓
!�>���'�����:t���}�a:�5q�w�����X����4d�&%��q|5�gQ�����z��p��;�2>V� 7p[������xggv����0A��hh�y4�,���z?~�������7@���)�$w�^'���{m����ϳ�Q��DJ�Q2[:w.���n�U\-ڬ�S�>����#K��@�7g���p�m"��" �փ��\�P�P���\�d;�v� wj�������0����z�!H�12!
��\O���$��=�*y�L��@�N���pκ�?n�4Y��A&���?Wr��S�W;CS������0�j"D��=A�0���@�&�4c:�$�w�2�&��7g;ƥ�z���$�.�x��=�0(Wf �
d�Q���XJ�$�ɪ�	'6{�y��n�]TD�	"���Y��BR���Nz��Y�{�����Y�}�W��Ŀ�ko�A+�F*f(���P��jDȱVf��s ���{��4��I5Y
d�&D�H��~�/)�F�}��wgJ��W��@�1�+���w)�@&�;���k�N#R f��h 3��Gn���-��76�>����]��6�1tq�ۉ����ʉQ2k�8�$���l�H�����쿕�״1f���-�v|1,��dȘ3&D!Ckz���j�*�5�$��Y��E�o7�|B�[uF%Z̵)zi����AF)fQ�FD15=��{���� ���[P�8Uo8�A묻3 ��~�U<Q-��ǌ"�4F�1����^�y���a�A#w7��M��9�B��tI#2�6hWv �
d�Q�}W͐A��*x�^�
�c�d��l�go!����}"�l�ڻ��M�d�=<n*J�vl�p�9�����T�V�lPqk
ut��R���@o�</�L 9�J���b����������r����rn2�8�v)���s��n:8��ю�^���Wop�#Vq��?\���9��>wl�N�
3��a^�74������أ��3\d��:��`����l�9�<��n�/s������F�]�|k]9���ӹy��n�dc$E��Qж�;��r��5t�:����yə��p[���띝�+�9�����瞸1َ�ֽ�t��7\d�\N��Lmg����k��kˬ\�]Fm�N����^)������0�e$dLL����x�`���H$�Z�ȢL�E�깋��$���1�tJ*$@ED�l��I���D�d
��>u�}ٛ͂����-���3�.��7��"�FD��*dB���� �p�ȠHC9*ff��5\��F�o0�O�yR@��j�"eJ$Cf�gճX� ���0	�5cȢA�w�s�T+kgv�S��`�rj�>�$B2$�m���]�D˩Ϩ�w4�2AÏ*A9�}L��U��,�;߯��瞜����c%��z���6v�7�et�1.LM��b,`�N2���AO)Oَr��I:q�W��#6�;s�;�`����z���������M�C��I����퍞	DTf�5[��Ojt`[R��W�k�]�ﷷ��/u����M���B�n+��8�v)�v-�\8$�
L.��u��K���7���R���|H��"�>'�:���`�\�J��3������&`D���%�Ʒ+�컾lٷ�޷xA�<��w���0wDHR$%!L�B�_[��*��d�p�� ��В ���6 .��S�����a�[ă�hI��*5L�2�!�Yoi�����`뉇uY��=�H$[��� ���������)@����p'�a9�׮8sv��l��۵�K�ܘ�ܛw� �_�?��t��'Ќ�4\�	$k���y�L�������А|u��#k0
��d�6�o�"�&���d�8�I�>�a�n�H#����ԣ\a��`��\LDD�
DLLD��ۡ�o;��IQt1N�j:�q`����
k�k��!l;FWj!��u$�r���"l�Ӽ;<5�zxlz�ۤ'����۟x�{�����~yz����6H�y�f�	�d��v�(A�@�� �nk�|Ono6�����ڳ�+���H���0flD��)�t�:�H$;y^���2z�B����»w� �۝͂H��*P����)uN��e&x{CM��[u��n�i:���j�v�G����� �w
��2ff�"o��ϛ$��ަH �S܊�g�TgVA���`��y2�5���{�B��{?=����[z���ަ ���P�N3%��Ev�4:�(��S&J���a��BO�񌜕�Y�pV�8�y�͒�h݋��I���4�z=��U���9s�Te�H/_:d�I��"�9�|�n��a�����f��.�c�̪�x�ƫ���pd�˃�
}�t����Z��6Fo8�+z�wPZ��V
�l�f:��ddL�n!�3xx �vg����z&$$B��C�{$�W��O�y�'FO��ݠ�H8k2}}W͞��mo}�*;�
������a	�H�����5&uє�.��@��c��t�\��3����|���	HS"�-�A�]� �}W��5gB���9�[M�A'vT���fʉD@�-�Ɲg?3ね�{O�t�uљZ	#�vEH;|߉/�0��V��l��Z�-��'������2��fBI�7v�����uj�vo'L�P��s��Z��	J��Tm>��[�e_W���`��I����	���qBdq;��O�� !=��'�'�x�q4gf?0A����UK3�����q^$������w6hM��W"#f���ų���=o�,�t��F�Z�\m{�֓&���y��������@�`K�V���F���OO�{]�R�g�83��b�Nh���jGTԑk�x)�"���g�[f=��v�3;<SM���|�}N�<4�E������6b�ո�Ft��o�kyvTCo=��}�����g����x�o�ڞM�QA�Y�P��	�URM֣c(U���4j�����wS���}�d:��n�:8���s�������y�u��:�J"_���M�~WC�7rc_��Ne�\���a���S�|6����t��3�����������<N�g�uW�5����H���o��6�o��2q{�-��r�4^��ry�j�o4U�>;�,��5�f���<=�7��?f��CQ�{��y���K��wzIx�
�]\c?g�����:�#yB'3J�Yv�wr�b7;Z��	}���1c>���Yݭ��b���0�B�	e@[/kkv �Lݒ�ӧ5�>��g��O&�Z��W-J(�"siͿNR	3��'Qћ�������i�[�^�vw�i�){�6q׽�U� >)��t�>n�B�[�WoN^�9�c��k_f�y=�l��HeE�Y���l��Ë $S��l>�]`s�Z]ؑ`��}��L�:./�Nz=���G�N`�SS0n��b,fz���o���#�;�>@y��`���N�����^����sb��u{֑$m��G]�.��پ�nڽ�{o]��ȭ a�0D�Yv5Y�زM�->}�G�I�#5�iW�B�E�I�TDEWJ�Z2�RE��%6�:U��"9�R���k�s���J-YЊ��\�1�����+��r�A�&�dʡ2,�$V�Z$D��E" ��RE$�ET��Ӕ(�Il2��
����.A\������"+9(r��\T�s���aJԎ�F�"�r�T���,��-J0Ε!j"���knXF]H�Ab��Ĥ"�4�jiB�W���҂�(�jT��-˃�0�(IN��YZQ��B%0�i��R�0�L��*TE3C��J,��*C�G��D\*�G�t(�5�CJQ�J+*�
g�qTa')1E�ks��'2�!d$�(�:f��BYĳ�*8kJ����KCR��r�E0�5�����vǼ~��ގ�\p��g���n��7�V��~������!�LA<��e�W���m�����C7=�Ժ�A���c�_b����m�!W�m0������|W��V7[&ޗ����t�\b�+���9����Q`�UӍ���NZ�ܱ&���ݭ�;vҮxH���9y-���r�Q���\�xWC= y��oК;on2ܥ�:���mz�R�]�Ŭ��<<3q�<��ܥɡ�Ԥ�T������'=cVۓu�t��Z,���ƙ۱z9^�w���x����F��ח��&G�㇛v��"3�:5���H�ʷ�/�8��rst���9��Ƕ�:���o]9�5iĤ��A�c�+t ���1�͖6sv����sP�f�Ip�����o�J���&.7=s��s_Y�6�sκ����9��5��m��=�VB�7�ף��w]�mn4[��{y�N	F���5��1�;��Ϟ\����-
�>���N������v���v�wn�\��b�:>��m�}Gn5m0�x�� �rnK��ez�.��\��7a���lH�=cj�P���0�cZR��nhk�I*�97m�tbqv�����3��wb�Jlc�:�f��7c���py����X!�ۦ���/;�K&�Y�^���N����67n �J��@ۋ���}5�g��lf�6���۴�6��[�P75���.��;k�,\�=D��a�#�ku�4Fv�q��ꛮ��)��f�xKg�������Z�X�3��n�j&�s�9D��u�l��	���ݞGq&À�p��zr�ˣh+{7;Frv���kc0�`�ڮ[O�����:��Y%���c���r�'ʭ�{^���mr��Ⱥ�k���k���v��c\��&7o5�׬��A��tv���=^c � n���;�vg�n�ͻs�Z3���@;]�fe.�̘��Ux�8^�4��̖n�+`�{������D�9n��l�h���Ħ�����{�����m�m��Ϋ ��6�@U�3��{��7ˆ��Ǝ��<��7[��TY�]t��[�&�<A�v�{k����/} V�'Q�a��]���� 0i�u�ne��v(���C�%���.��"��X�u��
�v�a�66׷���A���:�ݖ�d{Nc�i휶�[������\u�˻kdG�H6��t�ޮɮ��+��d�����mc�\�{8�a��Y8��
�hڜ�fٳ6[[��)��1虒�
fN�6kr��r���H>����Ĳ"PW��=�R���^���)n�2 %!L�B���d���Z%����زA#*��{�͂A�7��C�ֺ��⣦J�ȑ4�j^m0H󻩒Fq�[�\k//��H��^6E�wS6q�12f}1}&�������K|I��#w{��Igc�������<�=Q(�V&�d����'�u��xL	oA�I����$vwsF_9�Qx�Jf��)����n93瓦x����8[���-��.K]`�%����0����萢$@1&f&'�wz�N��S$A ���x�M3Ԇ������w���HT�q��3%"L���{T��<%^�UȚ���Nm���;�p�nHp����!�q�+!��7wb��L��N
�+nu��7�*����/�>u��=�9|��}�
�;���:k�ձQ�tD��~!BK�I� �2!
��`�e�РNP�G�"a]Yd����lI{uG*���J%)ȑ-�Ӯ��3T".��@����A ���@$=�ǝ5ˌQ|[��O�mD12[���ŉ�;�����Ⱦ���w��ë�Mw[lI}u�@}]��al��Fr��Y��J�jTJ� �A�Ӌk���b�q�us�Nn]2�Ϡ�v�b����������0��n���yB�>'�g��M�ko�q�虭l@#��z�U�KŁcl��_��g�e��r,�DW^i�ڮ�F��׉�!��6[/�s�	�觼	
Z��|�d�B���{t(�}�A �h��P1Y���TQ����3��T�ݢ�w{�H�ͭ���N��F��kvɬ�;��;@�*j��fO����;�ω$�{C�	q��L��%�$Ȁf	��{k�5=ٷƍ���I]�� �OE�0�Ngw<Y��bCD��U�¢��Q�"[5/v�7��B���JL'3��$��o���l����m�Q�����.�L+�tκۙ���n�h[���p�Z2�<RDI)'��6Lə�L�&'����Gĝ��`3�|O�;y�z��
��~"����+l�<��D�$,Oi9&���6�|����4Q$2;1�|H��� �&�1Y5��\�J$@(Lʘ�����dnv�2I"N*�T�AV��wt�$���>'3��&%�'�fRI�O�Z����)����z	���7��� �.�
�G����;N��̭-��Dk5{f*s�u���nD���:��R�SS�z��*�ڧՑ�'c�瑚�Jsu�QήQ163AtB_ < ���*]�L`��P����Ie�U,z�}D�uc0f�'�T������.�(Q��;#�7�9�6]�cg��z0n�u��[��͙s�i|��8��j�H�R+^l�&*f&)R�rQt�_���ަH$n�&�ɚw6�գ�k�$;{y�qd�ʙ3 �����"��Q�+fnԉtU�ʻd��� w�@W��8��w�	�w�T�A�3�]u �G^e
$<��ġ�]w̟��͐2�*��R��&aLM�׎Ĺ���I�$��u2A$���H���@�Υ�0v���o��>�j�p
d�)�M�6��9W|�{YYvu�}u/��E�e
����ʋ�svDT�ӓL���B޷�rݙ�I�Tbe�B�3�kD�]k����I=���E�Y�r��u�W#�;�l����{���F�7�1��kŵ7Y�r���t�����S&�L{�`���wZ����(��
;\��ٰg��!��ݠz;ckm�u�-��o���^�ƞ��[b�u����y�;��ᗕvNݭ�%��؇����k�A�:�ĜO2��������; �s�š�zx��玷��G<j���XЉ��nݺ�Zۦ�y���%��+�KvMBz�s'.6�	�(\���r���7m28���H�5*x�;]�������$@��>|��d���^�A7=|�=�sG���3{_np=��R(4�Kf��0όأ^u�{i�x|O�<�	;|߉�{`\(���Sm�=fa����|3_�<�_����t�����vm�A ����9��� H�y �	�"[�m�Д�����z�I"�n���a����}�E��.�>#��ۣڪd��<8�-=����3s���Gg��l4h@=�� ���	7��LZ���S��aP��#����������n^�/A��1��]ˈ�`���QSBc���d$aL�|���|ɻ���o��ͨ9^��#<H���1�h��D	�B����H0l�̝�cX���C��H� \G\<U���0�n���k��o\�~~�q�4j�yU�2U�5j,D kZ��&j�l"����N)��6�^h_�m�}DH����M�o��*�,nZ�g��bl���Sf	�`Լ� �{��� ��gU+{�LU���$���l�	���6 �5�M��������o=	��ô@$f��~$����j.�fGf�m�R�i�d[��J
�S4�m�l	#�ez���=�ܺM۴�����l�����z���c{d�ߣ����صvz�� �^Ŋ�5�#�;��\nWu`X�XD��yy2Z�q�Z�����'s��0O��&��X��S=7��`��ަLIz#�Q&JP�f[���
 ��ֽ*�]g/7<���ۻ͐|F>��u��jq��T���B9$�@�`B��m�H��4H36�,��k/q���s��陾��q���I����`K�i=ݚ����b�.x�QE��I��X�:�mܗO�z���g1�x��v|I=�o����+�2���� �C@9������t����L�A&���"�]٫��7�� �zO��|���x�@7�_�E���~q���*��Ԓ:�� /���O�{������\��pŃ�!@z�'.2�f�.u%�{��y��;M�^MR��$���킡$�	�&_z��['ĝ/2�$	�{��H�J��^�t����~cؼ�ie�^�f0��Գ��K�v۫���/�(�	�����͇V��s1�^��I�(���t�I97����Z�(�B"���޻�	"�ez�'�;��%B;$�@�`B6���n̳7��(���'�=��$^v�Qgo�jd���<[uX�_�����k�s�v��ޙ۵3�m��\�b*�R�'9[��W-�n�xuEFGi2vbsU(:��qU5����<=�W��8�
Ȝ��0��f�5/�a�/w~�Ma"���r�$�VM	{���o7����T������~n6�|]ᓬ\�ݱ׮8r�+����7]�[v�y7n�85���������̹⿸��D���~gĂ}y�̀L���w�x�wu��s��9� ��D�3-����=���،��XȷTA>97�OĂ}{�͒WЧ���3}"'��f!D�%L �v[g����u2I=�btUsS������"�{��/`�$�JL�~#q�k�7�:��[�3�A"����ʫ$§�1`��U�0bDh��"D	�V�w7�A ��TgL�.v�C���$���l���V�?=d�߃�z��L�F~Ŕ|/�ڗ�N�ͅ��A�$�j����e��0����xAq{�&e��W$�zz��w<u��<�C�O�ٙ���	`� �CD�l��-�N�n.��؏�ә�=nS���v�f�6���Żv�Ĝwn�G<��w7ܬ�v��]�=mջm�g�v�&ʽǷ�{v�����ݩ��V��nL����le��F^5�u��Eg�Sm�{Sg����{.-�n�z��Y��e`c�K����7}.��[u�d�;�OV�q��A�(���f㙵�0[$�-��:+r�Z��ƍ��2����Ym�9/7q�y��c��=G�w����U�k
a ͉��� ���	 ��vM0��쳔��{��z�+˷���$��)��<)�V4���ۄ�L��5�ڟ{9��@����?�@$,��l���yU�.w}�� ����
Q�PUU6�ޖ�a����w5-�wU3[���@{�zܐ ��ͤ��d�533U!UIM�{��!�{"��Mz	�m �o��iH �Q��v�D���̽5X{�=��so����WH�Hp���i�	�Y�$�{ݚ��7so1���� �c !m���d�ٹ�s����㲓���A���[���l:��M���)͛��y�8�q�s!�m#�bh�ަ��#<X�#�J��� �@�yͰw=���_�
�;�YE���2!��yͰ���&}4AR��S���f�a���d�k�t�z�a��-;3`���ۅ����g�3�{T{ʁ�2w	7�z�����si`=��LA��v�#���J���6I z��4�@_|���M��VWN�mcN����9���6�ǅ4���+�w� �z�`|
r����\�� ��|� gs��H���!HF�*fa�ί-ɝՙ1=��B[ƛ��s���F�u]oY�f���ښ:<�B�g7���$���%#3)Kk{7.ť䗒��$�&Y(���Av{.��{�����uo�����⬃PR5f�&&�H������A=���RG;bl�V^��c���:��?O�Ǝ�D�Q��c�i� ���ńDF��\4�קܪ|,{Ͳ ���`+��tJDH�`B����崉3�WWe)�Snj����d��39�݄�IyooK$��/�q2�_:[r�����;4@T�5�����H���H$K���e���wX���D�?d��|�|��
�*�ܣ:5�v�V��a�<�""�5l��K�g�K~ȵ�/ ��8���[���Q��asD���ö	{S��s���tl�S8��n0[��{�2o���C��q��-��[b��[P��Wd�-�"�2.��m!�]�#zp-Ep�Z��$g����1���u��ƮL�tm�+�_i�2ief���nvOrV�+}���;�r^�l��>v�eg}�V��ݻ��qkK���&�^�̱WW��.1��v^��)����`26VЫX�.*�I
[[9��,���F�&��\��߷�����_��v�#�7D_R��ȫh�x�S��m�=60]�Eӹ�f����w�����z�ᶝ��O��g5�sz��:�	�Tw�����ؠ��g-B���^13!�Kj�J��5Q�gJ���l�V��[N�D!{�ȼF����_�xf�U��������k�7�垹�>gć��T�y�z��1���f��}՗ޚ|�;o$��sJ8+�{(��z��OOv&Gz2��@�r�k�2q�C�b�l�*�i��,1���Ǳ��W�n	��v��C�g%�w����D�?j	��i?vP�ٱ�eY˩��0�$̬�^���3��Vｚ{[��$���Q�p�#~�5:�
n��pz�ؿSGn_���f�sPvт��u\!f���Or�+��jX[����;D�bk��cN�
�2a=�����M6��w;�dVo�}����&�&���|�i��{H^/|��/�8ϊy�y�I�Dj�jA\�hDr��	��'(�Tʪ2�:�f�VYU�P
�k(Q�"�(��*�"
.r�E%��UI��9*�'P�(�jȒKX�B�$�yˏ^S��q$���A�aTW(U���K2�D��f�2ar$�D�uB��jQ�M&XEQS*T�R@��EG����TC*��O"S����*4��p�H�5����At�*2iJ)j(H����4�(��r��$$��%%�h�I�eR���@�\�*rb\(�Rl���Eȓ���"�iK"��Յb$\��N*yBr"���,�&⨧-":�.�L�X�'
) ˢe$���U�3�x�*�ܠ��ϐJ�� P�|��o���_����I$����8����xS) p��{���W��]�V`H�μv- �	ooU��@,��^[l�b}� 7�;3K�D��*�AUR�}}M� ��͹�o5����gP
������ޫa�+5���?{�ѷn���p�������4F�ɟ<�[��m��B��V'����ƍ͍���;���o�å�;b�?>o���  �ޫ��ef����2����66��k|� ����DG,��& (�&���`Iã�"Iqg������ �]��p�+6�d ���ٗp�����|��(���!
�)��2᣹�7�"�5�ς �6�g���;= }�M��eg6�~�_�^o	x�C^��fo��s�i� ��ޫ�B��]�� �wnc�+���Ue�RH�n��!l�&�s@��f�V��N*�x�p{���4{x{ݳ���<��vq�^m���܌_��?��W�g���M��K=u �|�%y-��]ڹ4�o.o�I��z�$���tK�H���Qs�D/��{�g��62�u��`G����yI`��Yc�k�!HR��A���
#"J��}�S�M� �׼�l� �K׽���+Հ�u��e���,y��D����m ��蒦J��
�E6��ۙ��Ӷ},䊛<��SD��Gg��I����l%{��{ݫ�3Dب'E�		3�������z���` ��2"u��w�9��A"6s)��	ewkv ��'��
�)��2�;���'�Hw79_��]��DC��nf �G��N�wO�u�۶�Ʉ��L�� 2
����k�i$Ngt�H+���x��/�f �k��� 6�w3 H#���h�1��W��sv����MhX%�hUû�8J����LD�W�2�;�����Pbd��Y
�n��η�n"�~���������H`v��v4�q��m�`�5��Ws>P��Ǜ�cvJZ\��Ŏūk��A����v�ޥ�W��U)�[�FnE� �y��k]�kon7^�����s�!Dl�q����ݷE�x6��kn�d�zN�^Zx�9CFG���sqX��g	����<ݹ�R:맲�q�lq=Q��\�/�l(c�zs�)&X�������xRx\���j6ԫ�EItdլ���պ�ݺ��vC��G1��??>wř��M*Uer��l@|}�y�/{���e����^S�A$�Oo�`8I��_���%▄,(��-�&}؄IUF�i�U[$tK�6�D�m^nf =!�LI��}j���Ƚ3�!S�HJ*��}�� H;�=n@ /#}f���h�볮#����ȌH����.b<��TL�5�]��l{�rA�'��� 6���, sg�~H�6{(U��NA�1�]�w~	A�J4D"$H�0"(��X!�C'���-�9�	T��ɴ��f�4K@-��3UuQ�Z�kb<Z�\@L�U���tvݭ֍��ص>���Ks<c�i�'��\���"fz���=�w���` >xަ% %��鄖\�N�y}�v ��0�e�s%M@��eJ�Mo�����am��ȕu�la��5�Qqy�St2u䣢���k�5��/Mj��������*�h-�V4� �k��"QfE���jy3t��U��׾�I+�2;�?$�I��D��#ԛ�2����RJ�?eD�ĉ2�P4}�n2 �m{Ͱ�zd�L��8�y� �;����w�`��:$
T�H��2���q��̓|f��V�D�Wk.��� ��s.�N��F�w�F�[��T��zBeA�2��	Ǎ�I���b�uJ�o*�o/o6�n�=���+����),��n�O�;� �ð��Ģf�4�
���K�xP�[��.9�7h,u�x�J�'�6C	�����g����D�J�؇����>��]� ��nf �f���'���-��l>��	/7��	h8C���~&��-�Fx����Px$�@��:$����J޵u��1��Ψ�;�P}z�QP"h�R��B���l߻^`| Fs�Xj�>\����;���nH�v�M�����[��M��vh�|g(DN$$؝��b+f� ެ���U�A��R�@ž�4�w��2�>�g���x >?�h K����;�D�ĉ2�R����}�c�6�H_z��n�` {�s���������J\�n��<I*T�	��l��f8����c
&H+î�:��&ٳ0��%z��3>���;��v�*-q!S�����[��;C�9 w�.뗍1���t]���8]OkdSBc��|BeAP%I��Cq�Q-,��v-���dw8iV��ݮ�&+c����X��ۻ	/J�*8(
T�`D8����x")�s"�^�o��z��3 @�O2!�N�uY����Z�=�t�R��HZ�v~�w�@����>���cuU��N��]��m�m݄��K�ftsb���щ2R11!S��7�������w�$ m=׋ �]�c�+|��5FB"�r��:���]u��S���#���]��9�co������x�uh%���~d[S��ņ䰑��W��pΑg���)a��S�%U�	/>�ۻ%��H"_�6��_��D�N�v̒sVn�uuf���y�@|=�nH<��;��r�j1�����%{��$��	���B�״;��FW���t���ٔܮ�y��B����H)UDPQ��|�` �D����t�ukJ������M��vt�j@��(�&	UR�@��ͳ����gl��ҳ*}>|� ͞���I!s�ߚ$Ƿm��#�ra�M�~$��+�,�D% ���D�~(\��5䯫{��벜�ʻБ(,܎qI8s���	E�H��H�D� �׭�W� o\�$@�J=]�l�|�[)�JU͕��mH(��dJ�I��%�"�w%y.��ZDCȽ�g��o���>�u�?�!O{ͲHv>˲_u���*�u,󛻤`���'�jM��ʭ�=b3;�#��Q��/���i0K����?�]G��.�9�CXX�؀�pI�I0"&����-݇y�Wg��n2]�C븎��X�x�mt֗^�E��
���ۅ:�V�sV�ܹ�k��s�^or�vsGis��iۗF׳j���V(3/l����k"=��VL�mˢ�#�b�և�cFݛ�F^.��#�	��6^M�:�9h��E�l^�������Vk��� :�Hv�#���[��Y��yΆ^u˞!Fʊ���[�������;������\I=7h ������!J$����_�/�u� ;�6�I$���.��i���i[�+�9�]�"~8��}���!��JL��.�۶I͙��YGb��U�I$^7;�m| u��g���.~�F�T\��ԁj9g$
��&��6��m� �>ן`| z��g��3�rƀ@|,��l�����$ʊ�'��J10�C-q�n��wJ3'n�@$H�x��H�x�n��%䗖�n�ps����Ͻ��rO�$%�*���KA��m�����D��jzj'b<vޤ���v�H���3 Hѝͫ,ˏ~�����ϗBK·�ǟ7�<��>bS%;���ۮ�r����[`�G�/�����[l:^�^��}曈�޽ן`�;����ј�<�q�=��W�������9s��5�T�-��:����gO4�P�!{On6��^��ڄ���r-<�z�/�e>�{,ab퍕�'\�N�ߟ�v^Snm���A�de��S{F�ڥ8!ױ���M�.������u�C'�R���G��r���2Rd8����ŀ�#����� fa�w����u� z��3> ���mX*��Y��&	��M�[��s��}�+7�H ���v�^I{_9a"Ru��D��{��'��wwa%��y0V2Z	��a�~�Ұ�^�����g{����� �67:ݐ ��z�1\@����n��
�B�L��u)m�{uqs���^4�l=���Q���}���S/���i/���=�h����H�P��&�8�ﻻ�3��ۙ���o��^j%PIS(T�!_��&���s�e�v�،�u��I�'�儉"�D��'������$�߅�AËO��r�q{�� [����%O`yV�A��r��f��sZ+.��]�p�̝�n4�ٴm�x��"��܍��~��4o�~��~�s��j�g�oo~�@��o�  Y�[`S�ْ*d�Q3%*m���z�3ҽ�9�� �Lz�mX q�������Y�on�����@\�N6Q)��Bs��2@I���~�D�F�N]���BKл��I| �3�L��V��g�Ы&�qi��z��W�}�w���F�G�[<�k����O>x6�����e�I��������i6�_���!�V"�9��[��|+�uL��t��t^kj���w�+eI;34R������q���-�ȣ3վ�JI��M$[;�vI<L�*���^}`�z��D� ���
�?�?f�� uv�qS�z���ւy�Db39��[ۙ�6=r� #��:��Ud^Cʺ�}��� .��l��Y]�̈���}k�[�2������z��̝�f����l���#�2U��#v#z���0�0H��{X���YW�}��}�j��mӾ�ԍ����H��t�i.�fH���"�B�6w��b� �η��>�4՚��#�����3 ����4���7�Y}wab0��&0��769����"��}�����KB�6�v:�}���䄙�DH�H]�?6JJ�3��$M�t��Uy�&}�������~� +����J�)����%���	z0 C���W�jγ�C��~��ww�|F��6��<�!��ȂWW��L,��$�3SJ`���H�~�Ł����iY/���v/g����� ܬ�	/$t�u1I b�X�e����N�@���=��r�=�7����q?�_��$�N^���-���קBKݗ�w~J���8���O�LLQ��Ք��A!יT�f`�0zh�ҋ�W�>�o�to�ڲ ����cx�u�����/,��DPQxvh�k��P"B�y/��H�" 	�sy��#z�џ/6$/*�ݛ�n����f�, �|R�w�׳��N;r�嗝��?77��[j˹�{t9��ô����7�2N�0����<���{����=D���Q��O%�ϼ׀�7�����,�w:y�҅۲�%�lkE�B$�?�.�yg�8#@˨d>�Vs���q5|;5��M<������u�#��<����u�;�N�)�����SpE;����+gn�F��ZS��}N�6J�3��>)����G
��ޑ��|gg�۝�vR6�.V���͛{!�b��E&3�%n��nm\V�.���(�L���T��s{���:{�&dXD���D�����o�o4y�B�:��*v�bZ��G�Ԧ�^�l�7%��Or��n*����t G�:���{�z��NdH/Y�%7��y�Z���=����uRL���~	��w?�Z�郗��ڷ-�� �p{��k�^�������H޺���u���Ȩ���,8�"O$�K��}�OM�i}ɉ�:��v��>��d�7UA�s���Sû�s�V3�����������9Cq�]7o����Q�^��C�.�������5{|��}����6��P#�^�
~]�o����V-!�^M첲��i麪��C7/]!�LF���$ɖ�$f��^������_��,�t���^�*��͊T�7y'Ĉ(��DR�$���Fd�	6���'v�2�l�ܮ�8y�ck�9\#��5�Z��*q�r�ˊ("'sp�
*��q�K<Q��SU�8�ˁ<W\��ċ���P\��p���+i�^p��pER]āTQQ�#8��ǜ����N'x���ś
�r�Ζx�r%AU+(��9]$�.sqH�9�DA��-QDԨ�^2�E9*����EEfUQ(9���Y�⤹TQ9IT�57��W9QCn$��X�C�$g�r8����s�9N��E�p�$������R^U4+�RKJʍq)nk����.��7eܜ	���=�nO;˽���r���xQ���xqQD^U��QS���pX�<ER(�n??~��v�/��q�I땬,0�����1��u/��)Cl��g�ە�`-�Y���6ɹ�!;g�ʸ��n�s�7.��8������#�}���\����8<\񞍰�1��6R�C�ی%�՛�X�8��8������2��w<���
n{in^���="���<Ji3�Gi:�� �`�4�\=v/.��nuq�y�:��Yw�[�_F���(Ɣ�]]�mS�m�����ݺ���x�wk�xy��:� �I�X.cN�{<7z͜s�շ9��8C m�\��Tv9!��{;��ϭn7�����(d�����ڑ6]�/Zyf��j�ΰ�Z�@�1���uַ�T�����a?�_Sͷ����={;H]�U;#õ�7ym���>{-�����&�j��n{q�p��۟a3���P�Fx�e��=������s�`���Sp���9�������zw<�����;����z�]ۍ��NXz����ޭ��v�zwYn;{c�n����]A���t4k�y�5�^	w<�=`N��Ձv�֪Ů8�h���a���R6K�톨
��۱�0�vE�V�n3��z���������v眧=���ΓK�l�	������ps���?Ap���֧�[�u��Z�j:��n��x릈�t�2soV�sǎv�)��ݛ�7ю�K�s��!�����͈� u���b�����,l�1���{�3�I��h�'�Op �W/[C[<h��}[�'?]�(i7;��qk��[��vsN�RI͎�����f���g��y����Os�W�]�y�b�=g�a�;b7Q��͓���v���v��r�t�9ow=��۞�;)��pXܹ]Ss����֗����Lv����%��m�m��vw���qD�1�8�a���γ����e�,v���8ֹ�l	���<�ը=6��2��-�aNh�ԝfp��g��9������*�=yxqa�cs��mj�gT�;s�.7Z9�@\�mV�/��Fѻ<Ꜷ�f-����;��ʣ�T�=��Mt�:�4m9��sq����8�Y��X�:w5���"=����ͮ��n�$��5;���(e�@O���s���X�E���I�2�|�lg�hLnѷ�>�^��E�&�+��w:!�l�n_g�#n�Qc`���q�gm{^n
Ɯ�d�ԃ!^�G�ʉ�`/�]���$�;}]H�G/q�=د�pe�%�u;+_{3 F��J���z>Q@��R!�{TM�5�y}�2q�ge��y�i��M@/o�� ,�}���~�#��L5��,����{���/o�� �.���c��9��H >6;�ڲ ��������J�)��ـ=w��6{�� ���P�@Gny���{�*y�Ó��;��]�j�<��m�@Ӷ � ��B�L��������7~�M�rd�@Y��O�> Y���Kv���v[d�Tg\#.c;m{��D�S����x��.q��b�O!�L.�u���\[�d�s��DB"'�&&&޶"I��ͤ�ݼ�ɁW���Z{1�R'�/���;��y=2DT�$���M�ws�ŀޝ�*�>~�9d�L9Y���n_���t)5b�q�@;���	��R2{���GuFn��X�f�,X����+b���|�Q�gG?o�$�I��l ��sx�����}x݂E(��H��Rl=�M��g���, x������9Y7��Q{������μ�V���	3��(�C�{=���^g�t@�v������G�w�ߜdFv�K��%lZ!gsm0Ss҂c��R�*�p���� z7zݎ�:��6��?�Qw�� �����ǣw���W8�m�+S�3��<��&W��2A:�֓�θ�wY��,��u�y5��vln�"��(S���y� ��x�> �n�~��Oz��G�t�h�$�m���	'��	9�DD�d��(�u`��D��0!���/0;}�6$@-��f`ѻͫ A>�tZ��f�R��?&=��T�(���)����, tn��4�����z_~9wy-�ѝ��ں����W���jh-���<Oy+k��#nT��<u�Gj��������W��w������G�{��=�n������(�FC$um�d*���\�%��H�}���  �N�t�D�ny����>�W�������$��U1$PL�4q}nK�D���Dռ	��4����IMoeݤJo7H��Xv�)tq������������˝#�B|i�98�dw�t0�(7f�p�-��)�}��mh�r���~��|�]�Xy7[�b�(%���I,$�-�rK�x��3���Z����@ ��7�T�^�C?(��p�=��>�w`��];۾y� ��r�	z7=n� �oZ���ß�����sł����mkD����g��uvۼr���U�����m���ѹ��~��T�(���*��ۙ��O�]���{��6{��""=�t� 3s��{3׵4���9.��L!vC��{����e\�vk�;ý�oD��w6_x��%§9��6�;������|{zKѩF�� �	 ��c~���щ�U*�I��i��v�X5����[���r� ���j��ۙ�zg*z�&�R0B�2"I0J�����6EO7,�ݣ�ץĆ)u�v1��k�}�|��P�b%Elw�1�t�z;<�v >;;s0��zLܙ��{��� ����'�Z������0�fd���8'y�.�n�k���P$�}��?���n"#�qN'׶H��R���'�(R���&v���䷯u���f:�{W�@�=u��@#���� I^�mݤ��� �z'�&fZ��
J2�6gDA�䉓9�Hy"oo���{N�Mۦ��>�[�G�H�kY�<H���MI4QV��ۙ� q�mQ����꫎����?c��u��`�w9����"�j�_(^�m����څK�F�wJo��Nu�-cO�w���~�]���q:asP��!$�OM��&����hx�4ǀ=V��j;q=WX�13��6�n���k\�Y�ON�.��E=��l���gd1�����1x_I��Ѷ��3��Svc#�����Yz��fMv%�r�4WE��9�=Q�]����k�����gH�u�Z�ٹ�8�pe�Br�m �����ƀ��Ϝa��(N��ύ듴=���ί7j�b��M���gq�Q��mv�;��:�;���{lۭ���ϳu�f��X_!3�5p�D�Dʅ2$W�%�0�3ϵ��%��,)�fh[S���e�{[��|�[πۛ����T�J�!2x�u`����z���n��@$���݄�Aa���aO�����(wdz�s�&��L�U*����Wۙ� z7�����N�F���5��[�������P�P�K�l��L�TM��ֲ�՝�` �;��H�FC�|���ˍ��e͙�Jj���$�MЀsЈ��H����mX|�6y����]��*4=� ��{2# ��osj� 239�7��yw���S�o3  � �H�("	#'\��n�.}��A�y0�]�Dz�=������~gq2��&�+9����A�twu�4 fs��}���o;k��ם٘��rZ���BxĘ��!������̨7jc5v���A�k7w(�������Xʹ#x�����-��������2`�uM/g<�=��5>������ x��O� FFg6)�裙;z���/|��TW%
bL�F�	��žrI`%���{�U�c�W�x%.=���#fﮢ��DϠ��ER\y"��rxո�^�ywP�3wa$�;��H����I,���15%V�㥭����fu�a��@�)��Dæ=�t�A�ݯgLlϫ=�Ҁ�s4� 23<ݐJ=�wi���\�<3���� ��F�˦ur����옩r�u�cKe��1��5� [��;��	!�3���[~��K�lfy�b �����{�H��ś��=Ϳ��������$QSJ��"I���n]�K�d���\f��75U�@x��O��>���������.��}�N��d�B�IQ2$6�{oΉ&�;]�I"`
�;�k�fR_�ߕ�����ʭ�hY4������-0���NdK=�H���V��`�ե��Bc�%�(���i�~���y�+��:���L�'�I�PIsݷw�ʎ,�Ę0*,.-�2hS��Z�q�t6�@������j#�lJel��]��H�u%�����UR�*GW��� =�o�(���z�P
��u�o;��đý��nD.��"!���@�A��ˇ��� �;I6�7Gn��W���z.699�Ƹ�r�Ђ�B�*TLz���Ӱy���"PŽ�ZGrr"�o��^7dc����t�G�����USm�ڰJ.�r���*�����` _���@�mY��>�i�w.�*�褼��9&bdĨ�&e�ս�b��twu�4vpX�=Q��i� K���3� G�{��'�o��"1A5J�����1+���O���	A$1os�%��<�N��b��g^���ʅ�3Oið��f�Gg��"�Us.�Gc��q�EV:��j!>e��$�Z�PC0*L��.��n�B6/�UJbQ(�G�w����}������3v9�'C����%yi���C�7�/7�I����1e�5BL�g\���̏�-k�U�][[��&Ҽ�z�w^��E+{�3<"bj&
�#�v�3 =�RXH�=��9~H�
�N��۬;�wi ��ݵ%���<DD��倓/��� ��Xw*y���{i�@b��,�<_e?R$�e�R�5�����:'� �����ș����[~�JK��a�($K�eٺ̈=�:r*��$�67��d ���n��D�MTUJ3,��c%RŽd.��	A���I,ry�I`%v��X�qUɸI&k��It��d��!)DȐ�ӵu$�Wo9ݬ���ξ��Y�u<�	/���PI]��ew�ޱ������*�Y�!l��_��5���}�(�<�_��^�'E�&�AUR��.-_A	�����/�'ՠצ����Y� q�E�k��O񭆍��N�<�F��ӻ�vM	�8���w��(յ������6���w���p���]��q�M��݌��N�#��qķ\�q��ܯjN�i���x����í�=gR�����];�y��^�����͇��\]s�@Dn��'x���%뱟9L�.��.;1۞����Ek�]���}}}kg8����ϮNW̖�z7i�s;=U�6%�;�<��;Rlg�W��"e�w�*&%�$��FC~u�X_eI-+��l�9�J7�j�]^wQ4[�4��'��z����kĥY�p˯>��wNv�vvk��}`�p�΢"Yyݙ� lw+��7�i���Ix�ס"��"& D/�2�[�����y� la��3���纼 X_c~�*n��ɿN� �P��Ȫ�ɍ�wn*W\��ڪq��n�	���I,;��;9�g�L�;1���nȼ��ID�EPMUl���İ A���Y��֫�1�V��<t� �3{3 =�mYO-���j���,O�Qi�p�1b%Ց��e�̗b�tm�]g-�	��2c�������>t�*���-�q�� +3��g�|���I	���Ȼ�&�ՁH������	�|"����38#��6�aNF���9��e�K��,i�٧�����'�D�Q�٣՜�v���q<ך��!44(٬�ͧ6��x0=��ηVD�?fM������ ����� G�s��"L�u�.8������S1�!F��&P-![���@�_�34�~$�>���n<+"��Yu� �7ۙ� ù�K�m�H� ������L�n���*{{�b�x"&��n0 ��ۦ�����ߏ���qc�b u��RNmq`�q?���{�ۤ�I�%��M^,z��*��d�I,;�ߩNٳ�3h=r��s�j�X�D0��g�|<�,��u�q㊞�W�I���mZ�*:�7���8(�Q0bQ�Fe��x�'�\{���x}�L'~��ߟ�T���� ���h�Fr����MR�6���b�rB��������N�:h�}��� �c܈�m���?^�����8,$B@�0�Y3H�&���I+�.��͛�RNVn���c ����=�o	�oy�l�
~���{gР�V�ObT��#nM�=Մ{= <r��@g�y�N[@���ծ/ρ%5�Y����؉�Bo�z�gu����15~�=�M)G��\��}����V�	�#wQy�3U%�v.E��:���	��.�y>�;tw�9%N���:xc�3w��u�V����i?n+9������x��^^��P*ϵ�y�HL�F��}nos�+�-����}�w<�_�ɣ�44w�����
�W!5��#���N���r���}��:���w��!_d@��)�\=�zp�M�=�s��z�[ڎ�f��T]a�vV#3S7 �T�K=�z��;�ޛ���&}�̇�u��_O3f�������(R1�yY��hma"I�`K���Td��u]��T�{���<���	v;^*�,罧j��fh ���}t�}f�D�8�v���غd��n+�6���{5{=�:{%���v �Ozy��h��)ރ�q���7���(��Z2#�_�j@��7t����mJmw�>�� K�d���9ħ�	����&;�WCGDZy��h&yrʧ,d/dt!��^f"�[ܔ��{}��5Mk�{�.9�^�s��T5���ws�@�z�Ȍ�`����?`���M��^��s��l��'�e�Rگ`��݈).��gA����NW�����
�["�D�B�K�nl�P��T�#�rEu��O9�~�<��L�[�cO����pmmv{�>��Cv���vQ{��p��O\Y䤋���D�	�nG8�e�I�(��"Ȍ�� ��p^��#��/�{m�C�p �@��y�7rn\+*�&y�M\\r�Bm�	!D����T x˹@�x��Y���C��EG�rm+�J�8�Nn�r��\������')�.GL(��r!DT��Qy���8��QfTd�U���N�R+���B/^s�'�%�[��[��n$�$�"+2%QS�ZN;��y�J��p����"$�FcC��!�NB�2��'��<E���U�Ȱ����QY��.D#�T����!VKC�U�M"�幐^0�"����-�&�9ǄA�p8p���d�q�����rq9�Z����(�pePfT%BFAA��8ʢ�<�p��8�'+���9�.�)5yi���ÖRd����߿�����v@�	��m+*����U4�&�QaL�u�{���d��ƛ���J��a���0�:��̸��ΚndHV_6�)��Q0��rM���@|}�x����՗=�q��Ql>�v@�oݹ���u>R��e8ﯮ��?7�ro�U�]��u"��n���l� ��`�n�:�o���s��csu���1�����4�@߻[��ܫs�k�]�G-���^I ����H���SE4!2ه��z�g,���e�ڛ=N��I./2���Y�waɉUޥ6ef�{�l�,<�A$�h��I��� W���`6}>�ջ��]�f����$����)�D���o U��QTTL̓(�,h���yMΫׯ��q��; �]ݹ��߮�������)UF��1�*~�}�mE�Y�׍�v�}�ם�M�af*�����4�,�M��>�F���q�15�?a$��M%����MM!O}���~$
=���w~�[��E�|�gn�`D�o�>��1o�w{ܽ����q�'�59�"�u�)�����az��r�m�����n�￾o)A0�Lԓ���q{�'`+{�ݢRXw����rF�;�����Q��w~I<9B�(�$ș��Pw��iP�|�YnggF�q�u:D�������F����:�5�M���c������)�^�nC߿z�p$ twzݑ sPl���u� '�w3#ѽ�j���9R���U*�a����P��v�\o� ��,� �i��L�FE�9��o��A�1 >���A~9�������TD�~�+�Xj���DG.NGwY'��n����Ia�$��Vj��X�лvA��3L��18ug^�0��J��kM��b.�y��{͍��=r�k�f�� ����V4tl-�4��k���,0xX�Gn�f�7nuiG�3���^n;=��uy��p�n�E)ng����>j���<ح��ˍи���;C�8�].|��cx���ۂ���iks��k��������'��g$,��8�mv���/n��z��=sp���q�� v�&�{Bi�k���k�lg!�1zٵ�j4^��2o\뮬*um��8��C���c��z����7��C�6�:�k�䍪2x�v~��"v�D�Ҙ�������@$��)$�J�_9$�����ഽ�׭�� �ocj����
QH�N���ϛ����;r���9�����^ݎ� ���J�h�O(��{�� ��֥FL)�QJ����;���c�� ���<��ѵ�ɉ�^��{�ݨI�ç�4�.���4H�	��h���z��3o���e<@�g[T |����nfٙ;�X�u�������O���Q�<�	���	ۮŮӼԬD��0��R��L �zڲ�Js�s1g�����~:�q��߬r=�up��sk���.t�O��e����V����'gk���|>�W����c���� F>i; 	������W�WF^�ퟑ�M����?F&-C�*�a6�	����=�����ɗ<����Y�f\d<kA�Kwz��}34�
&���Ȉ��zxӯ��['�}b{�"�/I�p˥sqN"��ӗd�Lh�wJ��5���@F?]4 �ۙ��+v�.�i�Z��ꓴ2�$I��rM_y;	���X�|J�s�s� ��n�A%����s�(@9��6�#ߦ�
?V�����VJ��m��)i��vj/o��2`.�˸e{�EUHQ%(*b�����D	F��E�C�齸�6�~���m�������7����C����v?������G�7�����ʀb�`]u�k5�M�a��nŪ�������o�\k;��������g�|۷p�M�uu�J"㚙c3P�x���ۭ�$�:C,��H��%�?�ۚ@�Y���0dY�������hz7��dr�|�hY���W��E4`���6 �om�`�A�Go��D��%�0���oJ��#PS4�\����-󗝁^�<�������$)��e��s���m�]'8#�]m�	��/��_������ G�{n��ĽT�0H�2	��S�c��1lO$�M�UDCA��ۦ Z���J�f�V��b|I�@"��q`�Blc�܅�n�+�w���W_=����	*�m�?�2;��C@^sl��TOBž|H߇�V�)̪���gS��g[`��G[&�dZ��=s�<ӵ�����wi.	���F^sl67vڰ�"��U2{v,��s�R�f�m"R㝮KY5�r�3�*���]��l+��s:������u� Z��<'���7�˻�k�S��%�Y̔d��*ƍ�zڰ�"�sn AK��z%I��mO6�b���j�Z�`���O�PMMI5#���c��Ż��4��m+� �y�� �;���3�#{gt�y�kH��x�i���|jy�����f,���l��M�3�ss|��0=�/Y�8z�eI�+dc�	�B���ܧ�Hzt�� ��1$�X	Y�6�Im�Sk0j|��Y{5��T����@/��5����۰���Ɵ�sZ	���x��9uֺ���;V�Dų�pS�ujx3m�fq���9��)#$H���F.�ĢPHk̪i ��uS�Y��ƚ��3�����A$����>������'A�)��}~`��j�fC�^��9Ң]�+ >	}�M"n���I)2w�B�0�3�<mPd�A�J
&g�UE&�v�l@|���dA�GrwSK5��Z:ݼ� A%��9%�$.��%�G���"`����3lz������WNz8 �k杈 >�����dokQ��ٌ~^��Oᾲ}�0���l2�:!��" �om�dl==y�7����t����H27���V�er�U�ys���LF��'r�M^�J4@��޷.fԆ/�ԗ�9�Y}ا����w�I����9$W]_ R�D�6�Z�e5�[�>��ѻXR��[cN���r����&����KUk���S��������RDC�u�g��k�,Τ;��ɓnƽ�p��r��(o]�x�uup+�l�	nE75Wc��]g0�jz�wWmu�N��y�T�Wn���ts�'b���z��9���l�z8�6�ݛ�{Gɻ��n�i���`�L�
�n;{�"n�lclqκTW���m.5�nH)T�;ǳ���$Ē`d�L��t|��i�@$�{]0���z�T��P�ޓH8I������]ł�R*'�&%�w�g�$��睔vq�I$JﵲIj����H�09�kS�����+�{OTԂ
������o9�� >�ݶ�> /j�E��/�)�>fw6���݂ɬT�h&U0�6㷑y�6q�ٗ�oI'[�P���ۦ�@#a����lt�Vw�#��N=����s%3����E�a���>��;�ۍ^̰<��DB���F��[�f)2��<H�����<�ٖ�m�n�WX�(�ƭ�g\�<�盗��T}>� ���(�"LĉQ2��U�m��!{�m��>�7no��\�+��筿�@���	W�^�(	PdĒ`9a&k����x��ëir�Q�{�Ӕ~g���n�~��v���5��h?�糫S���{F�٣9�+��[�U8�oKB��������&���=f_��0 ��u�l>��"";ӶnEt�Ga,G��D$TO�b[�cl���7`د'����=9[���m�"l>�j��z��UDD̕M�}�o�Z�~��f��@����` G�t� �����̨�Ez^si�˦�5R��&��)6��a��H���`4�ܙ�x���7���� >67<ݐ >��6�Y�Q�WU�#`D�B��&bA^2�T�Fx�g��8�C��Z<j\��y�h�����sn:CT��|,��l> =�; @w�Ϳ�CЎ��ɉ���U�E$t�`RIM��L���$�qefݥdE���Y�3���;�$���e�_�@ng6�I(݂V� �k��B�(�I���5�v w{��� \/��s5�<Ț���2�x�W�U����@�Y��t���&�S�N��71:���K:x�n�+�O�qn֣�$��<�"N���%��3��~�=��)"IO�80��ܯ�Nc��~n� ��6�=�ca�:��7���X]k���NLL$
���������w}w�]|]��Y��� ����� ���6˙�8��)�F�����đ"dL̺�k��zVlby�v�q�Ĺ.qs\9�ۮ������*Q5U_I%-�q~�v ��[L ����@����Yh�w�����~HG-s
%&	S0��Cj��'nX�j!�:zw�PIf�6�I$E�m��L�5�\I�����==�d�:M��QUQD������@���p�������qf�ד�{}ʹ�y�M�t!�R�P$�XI��W��:�8�� ߝ����l�~��0=�3�WT���ڼ���z�pP���!/nckJ�7l�b�lY����t������<�#���OLzg��6c%���-�oj�<�U���q����	��L�hSݍ�	 �t{<�t��&�iWk�i/$E�m0$�=yOԷ�:4Oe���F��R�L�T8C��b��s�n5]V'�8��*�"j;v���c��7��%�������=�L��?4�H$�1u㖖
8*f:w9�ʹ�u�h�T�j����)_���n�����-��sӔ�D�$;;n� $z;<ڲ���w^dC�'�K��*�UƐ��[L Gg�v| S�r��.����uv  ��\��?a��Y4�����a���0�g=y��f᳎I[<Ѕ2Iܺ�� �t���oj}��UNL?`U���L=i�T)	�(�Q$:��`:%%��M�0g1�4�H�n�D�-7�ߩ䯳��� EgEe�bF9�	�� �UA>��ĐX�x.m�&^D����V��x��zt�c{�a��~��j����v�k�^��o���eo1vMp�	��][e�E��)��[�v�q�8���y�}�<`S����^�����پ]�V�޾�y��+�a��N�^�yv<Y��=�W֪�zm1�i���-�������wf�']����u����o=� �/}fIXm��ɣ�aD�f�������	ݸ��Ǧ�+,s�w:�ث�������6�J�|�VLB�o���^�P����O+q� ��B��Pr���վ������O��~5��N�ǒ�F�`���{��xz�B�1�v���oQ�uJ��{�!g�����ɽ�
��8u�cul�����fQ�<?3��G�A�{Pў����8osO8��M������N��μ&=��͞�Í���ލ���v�D5iV��~ӻ���OOS�
�K{p�+�nnu�β{�U��|n��9캷�fv+�Tҳ�d v�T^�ݾ���퍍�G�w�������l�w,�:���2�I=�C�}������qI6�I0���
v�nw{�w۱hݍh���0��D���S/��.���sV�x!z.��q�����Ӏ�	��WE^艨��/#*��	��Ƃ&o�ӛB[��ߊ*��L=�N�ܘ��Gݷ8�9���`4��wpu��ϟ�.~������7˯03�U<�y�+K�й���$o��n��^�|�5�yةX����!���Lt�ǽ^xu�}��K���UWQ�(�G���
�KV�	�k.Wr�U����K�/$�������(� �� �[�7-n'9$�dhG�Z�N3"\�9P�-�UZ�(���	\K���G�����r1;��Q�)Z�q̗.!ÂB��D�{'���Lc���l�S�YD\�*"���V����*�L(����Q�:��x��N�3R���L��+L�9i��$��Yy�F�Q�s���(�*��*J���4�.rQV�S�q�y�^K�(:I\T)Ĝ��$��&�[q�YJx�)	���J����tȊQk'9T�AY-VEQ�9�(�s�ώd��l .CM��Q*%�#�m"YEh�V�IeI����T��+�1�rW9�s����!��ap��;��n\qШ�E�)<���"��-�����έ;�㓚�����EY�Y��d�8<��Ü�q�];{{m�~}���],K�i��۞�n�����㸽��ڃ�'���n\r]9@��K�ˤy�Ob��!�;'��=�qc�RnP<�n�rK.ƃ�Ot���N��ۗ�b���;���k���.��J.	���Β�HN5�1��P�&��i�s����Gf����<��vy�V��tv�s���&'a��8\����d�m�Yz�<�7M�ۛ�EU��ɸ:-�:����6RB����r�9�CW�l�:S=�=h��w�4(g<n���h�ݯq���k�ɻ\v���=��r�s�y�-\o>�v�1�k�ǲ����V�g�n&���[h7=�;%ͻp�v��s�u���h+�w2���Y��olsv��6zǞ.����+b�l�Wj�Ìd�u���d�u��C�:q�P'c�<���;OU�,�^�k���a��N�gN�1�nK�Lny��<Z�l֗{DQ<�v|v�O/�����O�k�����۝=��욳�Ȩ7=Ƴ�J ����X��]���a��7f�>��[g���M�FK��Y::J�"sN�Hn��ײ���n�{�S��&(�ez��kث�y�l��1*[����mZ�x��32��[�۳k�9�yg�y�m���mq��dڼ�r���gfVl�-mF�Ι���Hҹ�ϭ�H�N-�%�;q�ї<��jΰOvi]y׮e�lYp&N��d�/[�;�I��k{s�����Jz��Ҥ���p�d�ȗgF7n �&T�AKЈj�w�0�;t'W���Y�j/n�nK�,(���.՗-����vfۆ���gl��f�xw%;��<\1�n;tU�gƠ�j���-��֢WI��n��縮�^7$vy���W,���̖�'99	���CGۮ�剧�;�:XM�{=B��ۜ�{)&��֏Z�ι�(�7�u۷7Eܼ��'71�kN�%�Kfډ;��r�Eʝ�m�qM��č�(�+�u�n�.7v�,�q��]rp�V�
9�e��sqOJu�i��N�T�8����#0F5��6m�z����sˮ�X��v���n��)^�I�ܸ�=�0�y{>9+�����\t����O
I��2�v��6���-�z�tk>Bʝ�
�]L�5ɜ�S������� ���7�/n��n��v����&vx#��68�|��
u�=r�-�rڰv����u��������͕I(�H���A��%�N�̩i�{�����z*��Ngg#Ո���� t_ct��'�L)D	*�;�� ��LרTt]�� �gy��;���3�bĚ�"����$:.�� �ʙ������o|�� �v��C	�V\����s��@#љ����m��6Z���������b#7��\۬_a'0��`��v�c{�W�z��#?o�#���]�ϴ��k��<A�m$ԆMv�� ��[��ޫŹ��o�&�ےI{���$Ji���JA�Ut�_��X@�R-�Kh� &Z7AUF�F{N����J؈���o]��>G;>-t:2�vsN�ov�L M�:h�>�ɵNӖ��=ݵL$���@���{>����'�@Zz�&�����E���3^�����X�mB
�gc&�K^�YT�&z�ˬ��g??~�xZw�Ḁ�ub_���7Y,�V�D�z���� ���3����7H��L�Gm�2��
K�ӧ�>1�1e���v��"x��I$��Wk����o,�uh	���f`tgy��j�G��*f}*�'K˪�ڽ[yV�̈́�Sٶٴ�^�}�I%�f�;�Ν�/��d$�V�]ߒ@�]D��`*�X���l���'lsW���U;#�P
kss0 ��w�E�|�,�YB̘�d�!($�$BoZ8'޺��[V�nD�C������z�ɹ8�s�߻蝨�1T���29���� �޶�	 ��}RMܳ��]L���]�wd�~9��f��du�_^0��|L��I-.(��{͒w�#��鄉K�l
E%}��%� �w��yuى+���0��14��6�`�Aя�L�?8�9����W*����Np>����'��ج�{?o��u�[߬���N���2c��D�C�d-ȗZ�8ꢕ��y���Y��:�_Vޓ�$����d �|݇�mx�����Q2��:��:kv���� ]?[`�}t�-�ofze��^6�4hy�$'<�H��l��e�	z�8H���Z*�i��0�8PI e޺~I��CH�of`N�z}YY=i���.�/�IA Kx����J8�+x�=���u�;�x,^�	�vn��N�'����~sOhM�Ñ��]C�7b�v�{3 �r[9d]O���rK	6��%�c$Ș�UD�����{��M^S��I$��{R��;���7���L���2����{=2;����"#�����(%ٝ�ť䗒!n����<��� lc�Ր����A�S�	�k�$�e��}��Sҷ�GR��������wf` ���LL1���
�2��*�+�Z�d[�Y�Bz�7Wzu�7T�E�`�f�b6�$^�|��H�%���������;sE	]��$������������T��}�� Aћ��V^z۹�q�e<	Q���_�]��wi ���}m�ID�:{]���[cE�Њ*Dq���K��X�*����m��z{��\���y�v�u��ݴ�g�xe��(��,=�ђN%���ǭ/��}u--5�$�5&�#V��j���^_%D����@D�gmaaPx��۷I����ܻ����� o��3�GFv[�Ȉ������ ���-��2sp���0�M���٘ �mX�We���^� �Y���Ā�ڰ�s�HB<eH��i<W�1V:�����$���l�I.7�RKI,����yFj���Ivn�ݥzvb�J ��|fѓ�w� �~n���P�N��u�۽�� tf�vD@��7Eb��Rޞ���9����R#]�Yz�y�n�X~o�{��yOྣsi�|DZ��w�6��-;.n�'����y���rY`ԡ�ǃ��V	i ��x��&Ci���;Eծ5V��5�8K-��q`�<�r&�9ݸ�
�k'Q��cѥ�j�-v��csxutg���nv ��4�R�퓶�b�/X<s��gm�;,G��Kk�y�{D���kY�9���y�ܢ�K�<�ZM[��o{�hm:���m�q9wkq�$G)X��깜���'.�t�ۛn�6pl�$Ļ&�Sv�
ܺM��v�<v������n�˺�y���������8ScX�'�@�>��!'	=���r��d�qN^�n#� /f��0����xe���I�?��# n���w�Yۯ� �+�/m�/�%��8&�+�U=����I!CWbmaaPjX���`|���: �g��,����;�B f�l��`��5h�Q�g�f"&S'gk���c^U��H ^�˸` d�r�_���ٗ�{n�#l��В�[΋��R�R$�.I�O��H���v-_7�s�-��%�m�����"!�w��1 �MU�_��o��|�ʨY�:�[Su)L�.�\��nb�:�x��V�ݸ>������٣1O����0n����������9Z�z'n�x�Y^�l� ����A�z�<IS���*���|��Q�v���������nr�J���^#Z|8��p�iU�9c98����VK=϶�9�j��ff��
�Փf��Y3*r�»�n�{�^{�i�� �o���@}��vf �6-��3eS�#�kʢ	������l;y�����t���wLS��ˈ��_[� o��0�l⚩ED�LR�B��o�+k[�#���G�%������@ fw]�D�:�E\E7K��Y��W�ݖ������T��T\2�{3��m3��V�^d>=�z9�$�s��H��t�E����u���~�.(<��ػ�}:n�����jԯ�����F"�3�;�)G�I�P�Oy&z�b����|�Gg7m��K�w�vq6;X䖕�o6M��;Q(�(��A�s�JDݣ�/�����$J����I":멆�	qP�c	�$ׄ���stT������{?f}���/m�� ��h��^?5���s�n!��\�]}nm��V��%w��;B��&�%)��rv�6��vUE�W��%WoDb�jŵ��SPs�Y�ڕ��>ˮ@���dF ���kmW$��
�!���/i�.����<� �sv�#я����қ k�I�	��������4��:� ��Xm��nn���'^��Ȍ@s[l��F>o�!z��W��w�_��^�i�EYی�X�m����9�3p��{s���ĉ�>�H�D���4O�LB�Vx7�vͤH��L4JK��ip�j�u���5f:m��$��6�VÜ
B�b�C��ǳ�����L+�l��]��V�߰�>�f�q z1�jȈ�8���t��;�>Ί�r��U��=��` tc�v$ UCS��e_1̽~ !vs��d�}n�*�/T�V&���?-�����Q`!w� ����H�z�oofL~��~ċ��b�g�})����A8r���	��U��UF$c�ך������8ݷ�6|.�'�D~���>z� ��`���"�&�&)D����*I~K7��<���w�t�%�|餀H��H��oo]�J����������;��>��/W#]d�� �)b�y_^�UvOC��ݮ�f�u�������COi�<�������@ ���; H���ςob/'�⢻0��B7y�$�����%H�&|�陂��4V�f8���O�f	���4��1��D�����/�g,�f�F�^cJ�3�$!0&& 'L{5�� ���` ���&��[�;�.�$JXm�t�	!���d�3��(&��W�{�ˆF.#Gh":;�v �=�ݙ� ����Lw��[�������x~��I�ז��Ăh`k*�:�fg� �r��u����r�b5Q�Ο�|��� >]���_$w7׽;�t�Tdv��X��ܧ�s�!Vs�Q�u�B]k�w_GV��^䨐/����@�~��Z3t��o��4cQXi�a��4�C���ڎ(�=W:�ϗ�cWHq٦4V�n�\��!��d�Α;n�bz�nml3p��mq��	�]�n�X�w\������>'��\��p�UDh�jմ�Ucsk	� tXVy^^�u���$�D��']e��q�Ӷ�����8��i��۶-�K�.��]�g:ā�;'
�Wj0=�Y� ��@�wc���y-���8��U��d7#ՙ�I��M�؞�7c;mt���lų[	��պL��RPd��+/��$���w�i$�H��L$z(Q���*��=��ݤ���LL�S
L,�β��QY.H�SoW�\�t�^Iyf�vdF �;Ͳ^�j��n�����XZ+��*�f$��������ϰ �޶�"�~��Y~�έ@ ;7���@$���l5���2������?�}��)��zj�~���-��� ���'�w{�DDg�u��:}D(&���UlOy��a�7�ׯ'���.2�IO���y�@�:�PWi�bT���un؉zO��63E��0��nkpn�a�-q��h��t�`��R@���'Ȼ��D"�"+|�r��z�B�e]� ����v�+����6w_{3vo�`��_DTT�� �Hd�,�RU;aP�Uef�A�q�&̺�3\E�mFs����ɪ�_�U䳹��A��_Y� ��9�j�a-V2�?ZV����ʃ�Z]�hW�'���O_%����w���@#�>n�+�u^�pyי��j���UR�
��c�l A�>n��]7��HǙ;�5݄�����)#��SR&8�`�DRL�d����nzϥ���=��v�� �_��>��޻��w���;;$�>����lE(S�J���]4�u������a޵J�#F�K�I���$姵��wz����v���}�t�:D�" �����qj}�k�!�wS�c���E�;w]Gc����=D(%UDE*}���� pzӡ ����-�%�~�����Wkl�fm�*�a�B��5@��U6��y��w��ͻ"�����&"��/��w�3�>ݧ9+����/.�ZL��QPd��-k1�G��w�,���_N��RusW-��i�f^ۯk���64��� �ݳ�N'��!�L�{�W�܀��c��{ê�wf�\�ٱ�2��i��I����q?u���h�6)�^(����z8��^�h�����m�om<�����x8Ǎ�H򼝿1.�{<����X���}gx��Zsq�ߚ��ŝ��.�!��ޥ ��O]����]�s�K�p<���cFW�v�\���~��,���bl�FW���4SݔA�k� ��ϲ������پ�������*yr�xr���;�4����WA�Oiֻ�[�S���p�j/��fv���#�2ŋ��E��;[�����F6"]׽7,�*�T��[�2SI�=%}��!��������5�����5GT�Ooz�'�P��Mt�z>��,��.̓+٥�N�p����i�0�o=�sG+�{��KP#��ۆ?@��w�yp]䲏6d��/�Z��;>���xw���d��N�mS;4&�owM�u���g$���ǧ�ݢu=��}��ѭ���-'���+�_�s�̌��U����̳}���v	�J��C�ݸ+�E�W��os��¶9�=}�S�'<]�������a�w�O�VY.��$׺������{�)���/�cX}�w+��17��S��������$}{��x��@�N��s���W�n�Ǫ��{�~�H�o��Gs_��ߘ2�Eb�H�W�!��h3��Oi'���[7}�Vɼ2��wf��p�.YX�/d`^=�	�RQ�WP������"(��$��JYʬ��R�5SRD.o��Z���f�%BRNsY8�9ŬE5MY\x<���v�xvvTC��/<.0��:��qQ�4H+.x�8�UZʔ���:��ʹZi�ʪ�H�ǜb���P���N��kAf�iTTC�JV$�H&F�e��F��ÂSJ��ax���BT	�DKP�.���q!��r���#��I"�VgB�dIyH��Eq'�.���#Yb$�L6IR�����!`S�+�B�Bܸ��A�]�224L�"�U��%$�h���S,���!sj�Z���$��r^s��TQ�5��E�\Ќ�UY�[$2�R��0�,L����ّ9�8-�E�R!`��\�(�Mq�QC���S+E*�\��&Bt��4��R"��(i�줚e��i�f̭�W9��ED���4�Q�q�<y�eZ�P������DD ��
5<�K�r���)�A �H$�FN��	$���O�@�ww�ρK/b���5R�*��\��,��W�O��/�XD���3� gy�dʍ���޽"��� �<^�%/P���}b`J�ɍ��Z%��e?4ͩN����2<�Qm�$�vv���"R}��S���FR�v��b&��-;S�8���C4
���-�NcNn�k��מ�^��g:�#��R��$�_T0�	n��H$O�iL�92n3��­Xۢoofb'�=D(%UDE*qq�w� �S*�9�*����ct@�ݽwi$��ٍ�+�a��Sƺ��r^?N�ϕ��=4*�ST
*USf�<��@$�[V  ��^��o��s�[����ۼ� ���y���_DTAT���4�A��f�-n�M9���cՀ�������3�87�јsg�w���WuV7,�่{�F�l�����B��)�!>3�cu^����	o�����G$��DK�@�����N[�{�	?�4��S8B,�-5x䴒Wj��:D*���y�l���o���6��{�ίh��8�)@ �15�c��c�6��Z��qg�v��Lݥ0�r��?����V�h�&29|^_�3 �c��`��s��us�ھ���^\w1�J��2!O�ELC����n����L�_7>�����oy� ��y�@ �3��0#�TnG��u�y =��DJ	UQJ�C���� �3[� �U��fR�O��o����Q��3����[2��f3e��M��n;S�!q�lfu�4 	fNs���n�_��Ny#��jK
�W ��*�3I��o�����<�W��s��{ i�΢G��[� ���x�U�i&u�T�����Þ���ʪ66#��[�%y��ע1�����V���G�������5;�u���]���ϻ�{߶���7'$�	Ăa$�͛Σ��;�ݚѭ4���{vՕ��a��<sƺC&ݞ��'e(u�@y�q�^���k�8d^�9%�9)8�ܶ^�O�\g�mn�Wm�q�&��[g�v��FwFl$;9µ�J�n|����ض6<s��4��������igo�3��`m�]�e�E��Me�ڍ��=mb�n��ͧ�g:�e{���r��8���eݶ+���Gl����@ܼ�j�yqGO��u�5������i7��pa��]���I&a�ӣ�v�7��{�xk��=�mY �3����OG��!D�TA��޻�K#Y���r��b��Rq �2����ۻٙ�FS=sU��{�;=4��A���!�-�2���#����0���U����̎��� ���r@�ݻ��C��O�"PJ��dM0��oF��sK;eѾ	 �܆��I���v�)q�Ɛ��g�z)�:n[���=T*�b�R��_����$���t����}Ne��~K�s�~H�/;z��Kˏn6),L�WLM�u���f������|�uP�>s��O��v`�U�níl۰��p%��Yz��������nӮ��A���Z�����v�����鉖�|��[~�W����ɰb�5L&�I�q8!�7�ba.x���>	��1�E��)�t*���qԴ\H`�j �E�����j3���.� �>�,�^S�!�k񆃇z�V1�;rfFE"�+VY>9u��r�K�.��o>�#��ͥd �GXB���5�P
r%HD�$��Okzٰ�KOfSV �Uu{;��� 	g�{3O�������A���LZ�e=�� ���=1?D��x�7�t�@�9���o�p�'�Su�7��
}�T҈�M�8�m�| v�:g�uT�����������y�C �� ?,,��Hа���%�EaW+r�n�7�:N��r�4鸬7"\�nl������������T��<������ ���r�r��=~����m����:7�u�/�)EM"��4�A��7@u�n�K�/n��[���w��!�{������Uᄏ�=��$'M&�Kq8!�7��@$��ЀA���9��0DD�5�Dtl�-p���3��O�^��c[�sy�;}1�}���|�[R�={=<��5TU�Ea�+p��a;y�O�Zw1�D�����B��2	 ʀp���{��=��f �8�v�> �'5� �w{3L�F���[R_���� �T���r�L������}���^\��U�π�|�0>�w��"�]���=�W��T��vA�K,�.�rg�������\��b��\u]�V�s\.aA!$��k�Rę�A2%�L�sv >��i؀����{���{��N���I8��5�0�	e"�U6������*���a=��u$�ʖ<�=����$O�~���������AZ"���I�2��7��iA4���i� {}���" ��˟Ns�y�ѓN���ԐI����_����$�5ļ�m��@N�;�﷣קW_ N� ���Ȍ�$x��tn+����
7wp��"�k����qV�7��0ImN�Kyw���էu�Go7�q��v�����E��$��u\%*�6�DJ%&Z{����J	i��Hs��%������G{���@|:/��".�`��O���8|�x?>\9��"�9���[��q�1�����ӗp����~���F��'��ݷ�vy�g���� ��΢/�0���p��,���I~���I+�HE�$DB�Ȗ�3�ߩ$��"�xud���x{�٘� GE���iU��\C�ռ��0ڊ�S*�R���u_ff� ���4 w�������ɿ$�]��vM���]�%�m��d�(���$2x��@"�\�q�]=�n1 _k� �|��{m�[�a�'���ws�K�&�K���Ǎ�%%v�?9�w�ӮKO�K�;�=�ݐ|�G�|ڢ���R��j�@ֈ�/*�Xq3��c'wՓze8���n�_.�z��}�{N���0�Gݹ��⽢o �:��?����ߟ���.��-�٤�l�iD�mǋ6�J�[rN�Ƹ^_mg]�Cɞ
7�sr*����vܺU��c]JK�m�9�d�^����J�!�ccZ�M�zz�r;]ûo��a8��vλ+۶�tT�<���92.�ru���:��t�;5ۢ�q�8虓�>���Cf�[l���F�W�S;Jq�����>����bx1R�s�����8�Y�*�m74;t�%�O��5ƺ�.Zn�LAr�A�}�����L��g>�X |�m+�������ab�`lLGk�����[��O=G�0x�!�\�&Sߤg�'�__����w����| i{�� #p|���{$u������"���*S2M(�T�Ê�mX ���t ����=2�� >=�n� F���~��[&H��*Se�)��,���<�ٓ>����Ұ d�r�H�﷮�O��M	,�IžrXWkqE(�QJ*�3I��o�t���y�:s��r�f�;�Q����D ��޻��$�N�\����	t5vv���8R�]�sv�Λ��C]�'$��w�D�/�����)�"eT��rFG�ͫ���N��|�0t����V�v���������� �WR�`�B��
L����� ��%���eD�з=�=���{���yn���ka�>�:^ޝN�ƲV"˘1pp��;]c^B��	<��S���|�����"+�A�;5���V�\BVx��7�[�I"n�m&��1 >r_s���nAV�XmM�B�%*@���<܉�?ws� >	�t�G��3���� �:ڒ�7{3>�"c�I34�Y��G�n��Ј][	%�uo̒O�osd�H<g�DN(��[z#s�Tns��ư�4���KĿ~� �>���D�65D%zd{�����a��׻�~O�;�XR��BH"�<i�%W[���j�'�/>vS]�pM�̺n��K�����|��
�S����C�ަI$�S��o*�éc�&�gmcl�繼�9sq�&T(�!R��� �u�S9��Fv��y�O�!�o6 񞺐A��a΍.r2ﭓB.A�
`�(��g]sd�A�=u'�vr�U}Hl���!YSVg�$Nމ���"�gOo�Xt�ν�t��1���7<»�7a����:���m;�-��\W{�t�����;u�_�gsd�A�=u�qԎ�&�J!%"�/*������.b��g���$�N)܊�$�u�皖�!����v�9�I��a���P�B0&�ݩu��{r�����]�7�I��@�q��f!�^򗃎W����Dɑ �� �g�p�0{u����Π��^m�x-nڣ�{�߿7�Ɩ2ic����@0�` ,�sg&��ꞓ��;���z�#ă�+(	>6ֲd)$#aH���l2su��yq��a�m��u`��Ց@��o��I���s�&���x��n`��QP�-�3��A��>$����hi�u���'*A�� ��0I��JB�ݾn��M�<�������ВH'[�l�	}���Ԗ^A5�D`�'���ї��}E�_=�׸g!"���5;�!jc��rl�X�P��7,7�F�U<q2L؜����ۺGF�tI0�J�����yW���}�O��&7`�J�6+�n@��Xfﻩ�5*��Z(�)7��qL"0��2I�>8-uD�t6x,C����*�����<�ḿ>�?���qvTO�O.v��N���dn���:0\���ɠl����v�雵�d�Pe3%���I�ͪ�m`�g��ܐA>���.���HfN�j,(�U5�"�[&�"|��2(��l������ ��H����۽�]�����y�s�N�����B����3N߬݁FM��q��ov�y�@#OVd�|5�>5s���j^kH��GA�$�J)!Cv�7�I8z�����.�gj�rT��Q5T �;[$��? =�o�0m�o��6����c���0m�������c��|c���m�o� �6��`�6����0m�������l`�X6�����m�P6�����6��l`����m�p6��� m�n��6������)��g�)�1��9,�������_���0�?�� p( QUT   �( P( ( �   ( U$�  PP��o�� {�   )IP@( �JT�EP P   ��� �@H)RUB�J� �   (       GР h  P  @�
�       L   �     C�$��4�E��R;��T\�# �P��J*�JJJ�ܢ�nΊ�� �MR��+���(�  ;��f����B��AC��w�IJ�seJ�d�T��U�p �����DY4�	��'�s�`��J� ;� ��    	 y�]�r��O&)*31)]�6�P��@�V�p��<ډv���T�g&��w �U,������� ��_:   ���Pk�@��� ���� r��=�p� : \��  � � 9 u��@.  |  �>    t ��  H>�� � s��`����cފ�n��K�+�*��K��lu�iUQ� =�O��	B��J�|  ��{ u���T���z�rdfD�`ꪙ��= wB�F@�ڑ͊�fdT% P   � 
    H }�Us1US&�T�K�ͪ�L �U.fE
�"EZ�%]���p ��Psh�C&� ��/�  F��$&X 6�3a*��g��2���;��œ(̈́Td�AaUP� ��  >P      Ϥ��QY�Qf��d�T��Ps����S&�*�jPɤ�t{�T�jQ`�� ��� ��ͪ��s�Q*���QL�Q*�e
���,�	*��;p��r4�L�Q3`���@* P     ���JT�� L���i�#!�4S�b��P�0     T�7���)A��21 hɈ��1ت�<%M(       	2��(J �     �B �LLI�&�
zLF!�=G�ڞQ���~������L�?����x|�n��ա������	$��Q��?X�I$����I"�BI$�rI$��&�R�,�?�q��	$��$����5�ߛG�������?�?~?�?����c��`�hH��Ą$�M�*� �Wp	m����7�?��ԥUpiq�b
 HI�#�������̝��xw����7��p�O�UUUQUUQUUUUUQUUS�������$�0Hl`� �퍂M��plm&62�$ �& ��ؓl`��861;.�0N��Hv�N��m��clH�N6�$60N��� �m��c�
`ؓ`��`��lI�`�c���H�H� (cN0�*����y�I���/\�6���>�Y��H*_�T������������DI�}?~X�	����?�5�L���o)�����h�l��@�-���T]쵡��Nf^^�YSш�±ռcfط�koD�f��+of��7dH�2�&c��3c���Z�Haj��aa�WkcjYՑ���R�������Q�6�I[��;u%뭦��j�Q�n\B�%:]�	X�4Ӻ��M��IRP�/�� ke���fR�[*�D;QVaPT���n��^݆E���Գz�B��t��	���c77�
Zv䙂ѧf��f�U��ő�;�T�X�kg[7�=��{6�2M<���0�`N\834&�:n�Ʈ�2�&,��Y�x"7(\20Z���<bM�j��j$�D6nn���*�]A-.���E]�m<���Zzn�Ǘh���8�����Zk#����fe)�UJ��ݻ�9X�3e%�/u6��v6PE�o����W(b���c0�
��u�d��lT5t���wW�b|-����On�j�M�i��9q�o6��;G4���`���[b�4梈LZ���Б��-w��MɊ���G��d&"$(,DR�3[�,&�;�ݗXQHm�"��h(e��dݲ�J�M�
��4^\N���o�[�:��$�������]��%�;�.�'Qux��k�of�+Ȭ��wi�q���,��':�A�LF\��z�����n�N����A=��2�Z�c�KM���V� �P�!�Q�u�2(q�Q�e�Pf�ٺ�V*t�w�}�l��f&��{�Ɗ�M.��	Acn�chk��������)-�)ȉ��1��a�'��y%�wb���}VU���Qes�t����xX�2�Gnv)cM9��w 	Ҁ:x\z �J��.�-�of�𦈺mj�Ҏ��[f�M���<++5�C*k�ܓgX{I1��\m�Gu�w��7{��d�8TTN�-�� �B:9
b���9m�V忌9��%��*HL{(L��e�YR6�[t*9`66 Y4��p�f�^�G`T�jV�w�ދZS��t7�kfk;CHz�,�	 ����Vw)�)�؊ޘ�N��%�Sb��(^�Ų�7B�� �$0짍�L�6V�˲ סTr�D[ �űY�2ѣ�l���j�ڗU��Y68ڍފ7��w6��P��w�	���pD��.,L^KT�_�1�ZRXRe�f⻰���%�ʹ�+#ۭ��+0l�h*�d# �R�$yG��l��	��q�Ge��o-�eڻ�-��4\TY�v���?C��Nlҳa��.,�ګi�YYq�X��iM����m��{u�
w�����S�f|-��J�1�H��;��p'���fP$�*y���PnKe$�8s1�Vn���L6l�*�υ�w��;��۫�j��Kr�y�ӳ��Z���ڥ��aw��t"���2�`a�e�a��K�31ӗ�`z�]Z��9RCC.�$E�R�Da?jS5 ř�6��B`�f^��������3&���j��sm�H�3�t����,^�o��;�Y� ,����)�Z�"���udͬ�
��ʬ�i�h֜�
x񪣄��;ugsK��)YR!��Y�"���r��EyY�{�l$h	E[���df�U�-�oM�2)@=1�Mݧu�dT]A[i#�T��*�:�d�R�+���QF+Ju��x�̼�7[�T®,��:�^�u��٠�B�nؚ\�+P���X0hA?�n�:���h��b�nig�z��ǂwJ�L�0�
Y7�w{d�J"�J�,��/0M�J���9T|DU��ਝqn<є��,k'�P�Ku�nZkf�X�.,L�k�/Cf�T��#!�w��ɣ���;b��[f6)\�u�&���j��,�%����z2���]KV���晨�4�&Vl�wwЭ/��:����X�3��&E9��ɅM6�o2n�,�GN;�l���%�ˋC��u�D���E�Sp�yhlz@���>�������nKAڵcˋ7~�D��dn�`q"�sDΔ�Yd�f(3���3w=*��{{I���,���\�dڷuq���2�h�H6S�Z`I2�0�6��)�]�֜7B���V��_<�V�`�5n�5-���A�T�M#,R�{q\&�Vp
̵V��۬N�)��fB7P�����EY�y���Q���#zC����v)��+W�2��V�Ճh�����? HW!k#˗e��b���
��R��B�q2�C���x�4X���S�T��S�-6����������x]6։��ӎ�
2����{DԺ㵋,�*��Бw*x�)�m�"���7��<ƨ�`��f!bi��P�-�M��@rD0�I��[�m��*�8�C���cr�Y�����zue;y/���÷m����EPa�JE�Fͼ�<�`���=��.dG���S:6�ӈ+x�Y	�,cv�e�[��hո��kj������*��b���3@�23�CP�,!���iL�jC�3�5;��Uz�f����Y�nKj��7XS33��&P±fP!��T��z��;D�X2������nf�p�͟aTfS{���L�;�+)��s&6�­k«2#%5�Kw���# �_؆ ou3�����ۭI�I�iͤ�.��;x����x�E�u��n�ܐT��X��R��+c6�T�"$���J��,����L�E�p5N'DU�i+ت0ҏkq�%�Z�Ų%��H��6U�ű˽ѹeb{vѦj�n� ,ͻV\"1Z�i"���m��֡BWQ�i�[�R�r�E���*&��y2�Фj0���ͅr�(
X��u�{{�����E�Q͵�VMiVӌUʹkz坙�����0fLU�4�:��f���Ç3���*3# �Lr�""[�Мæ��а_�r��X���*�ռl�5*b�nRcL��yA��*2�U��9��4���ƥ�:��ѕ��1J�j�W�y�r4�XX��"61�:��<9tƧ��(�M�e��z���=lX����p��<۠MK�p�)a2���V`Յˇ0���8��v����*����d�[�++�y��X��Yw[.
vli�P6*�0έ]`�SDڼ3
�V���/+.��Y�@����s+s�1j]ݙ��0��	�� �2ܙBanF��[�
�.n7i�j����1<�<-8�p�(��d&���eZHt+&n<yk�T���
c�i%-9/S
��̷{���Be�7��#�aT��ڀ&�1YF���%��Z&����Wsv^A�(�wt��m��L��eܣuݣ��U���Ŭ��r8%�o�xÕ�Vj"�K
h��CM9y�׺��*ͱ��h���9.Z�<ʆ]��e���rڤv�4Q�+"�(���RD&Qq�,m:ے�I7$ܭL��%`�U���/J	f��x�B�������U��������6�E�͸w"�Z��n¸�lD;J�24�W�ţf��Ѷ�fM?@764l}�F�j�[�yOfeޭ�7B³w�J�	Xi`�c]���ɚ ���Gu\�͚�no�9�ͤ&@��[�)*��F{�����nhV����͵%���r�JQ���Ô�˵,�%i��6*�;��l1/	'fZ�뱫t�@�%�t�J���@N��MĊ�v�V�+�ì� �2{wJ:h�ZN+�2�@ꊥh�bA�6��鼗��ͬU-�&�.�d\	�E���dR�]Y�1zkw-Zafǵ�WM%-�g%Vc�
��Pm�YUxf�5�v]Խ
�i�݈�0�݅Y�2�r��u�9��X5�mշx6�^b*��8��^�;Ot���C"2P���mm��h�V��NR�e�W%�b��[9���өx\f��si^�%�K���<�(��-�jL�Ch�d����Z��.�:Ki���-�޽8'�����Y�E�ƴ<;٢��!�$�z�td5z��yw��1�7TGj5%�xlЩ[�V���1M��`���#LSxt�-Q�YH�ۼ��۠
XL�[�Tp�ui��t1ӛ��3Cj�Y�V���19��B��t�h�H!Z�t,�.�T����ʗJ�Yv�ۓUp��e�Y�U�T�M���PLe��,��Pc����[g�,��*9feGXP��/]j�r�J)����d�	ڼd�"�`bÇ	o�Bbs.j=-���UH���PgKJ�V8@���f�u����rr�a6�"��nX�v�XS��
�Y��K5��Z����wfP*]�#$7��t.f�>�U���R�iu���A�l`W�[���IQбnŬ�V�)�L㼈I�,]Бb��*��Ѐp�?�������6�a�j�sA��Xۂ�c �X��(哹"���'a�#R<ܘr��U��2`Uz`��;�X+�ǖq^e֋�b�TZc�ݳ>ڎ�[�V13�\L�#L���2��cH�B�pڥB���M#�m��~{�PClS$��|�HJ-��f�bP*Lf[�1���8e��d�b�4�)"�=t�S�l,VRw����� d�GE�L*�ܛ���.'k^���5-�q ���^t�rӥ(K5\
�uN�]ҩ�16� �X7V@j���b���r<��w�ܤ�n��l^�!�u�$��fɈ�n�Y�xt��㹺f����@���=P�j�Y���i���U�r��/|�"�T�E��8�ƀ�e��-�r�n�&ݕ�&hZ)�Ӕ�^��P3&�N`��A��wdʑͬ��mlȪ�/m��	�E�ww�u�-�Vl����Kl&;N�@㳾�|[ke�@�b�{f�`ou�܏k�� Y�&�.)�e�w�j-���[�a{K��x/kaS���ww�\Gt���k����Yu7T�!W�h�t�ҧ1�,$�\�h��7k ��������7 rnK������A3�f�쥀�'j*1�wYRaa�[*�Ԟ#S>.8�R�wod��E��'��QF��ܧ�X���K^f�ؤ��cJk�Vhf ����ҥJ�h������#)'6ⷑ�9"2n�.��Ij�d�.S̖��i
ӵ�R�
��Ѽ�-Bv��@��kv&@Q��J˖9���tX���q�` �� �қx� ^d�!������;�s�rE�.�̏,�&�Ė�kiS��n�siUټqT�QX��lfd݅�	��O�m�L���o�[{�dօB\�E��@�[��5�a�����	���S����j��ZyB,�e��l�C��aє��/4��&S��p��ˤͼ+l`�̊^�@t�H�AӶ\�z�3Z3 ��`:��z�Ő*\	�x;�r��$���&�YUq��e�ɇP����ؕ��O]Laf�g �V ��H1�J�c���h�k)�7Uڠ(ڨ5T��5o"#4ء���1Zњő��¼[�3*ݴ�z��e������m��)��n�t4n�ݵ���1S���h}�0Ŗ��^�a�6����g����j^w*̹Tޤ\[��i	 m�����nX�7
͂ۄ��ѻo0�w��١��Z�n����y k4�{w�)�,���5�ͻ�st\2Z�V(����F�٫�n�!�2�Ҧ���4�aqȩ^i�Mɖ�\�7,A�\FC@ō��ԧL₦�ʑJ$6����v*�a�wgĘ�2̋&e��!8��h��n��,��y�6�� l�]aM��0�5��!n�:��nF�r:�[x̈́��V^����]�ǃ.;z�5�K0��Pf��x�FD�kV��oE��r�λecUj؋ǥ�ɩa̰3m��sn\��m��e����	f� i�^ѺiLԶi�.���6dM0�!�@�hñD,�y1L�DN�ʹ��%�B))���b17ӼV��*�.��H��x���b�����
P!@KM�MAP�e���6A�7T�e��n*�j�r(r�kF�KY*��+n\�MF+U����e����VŅG4��XMH�˕n�Uh�y���O�b�*Y���Eˠp,�h]���G3i�[V74��i�-2]�w�on�5��r��� �2�z�Qe�*��FDI%"ez#36õ�1���|��<;�:�]s%� �Oa2���R?���}r����fϧ�r�0��0��}m��3,;M�\"���o�rc=���M�I%�0I&�m�la@ S�ۍ&�2����pc(ˌ�v1���]�` S2�m8���LM�lP�6�`����	��)��M�)�v
؝��v�v�l@6Ӱe�6�P	6'c\m�.� �pm����i�m��Cle�leP�le�lHI�����c�m�0e0m�0�0e��61�.l��]����� �� ��$Ć���)�6 m�v0i�����2�0������.�.]� .64��N�q����(m���81�"4~��'�?����������a����_�� B�;�~��W������s���� K����dB��|�pr8��B�������G���r�ﭺ�'�m�U����u���K�4����`�cq��CK7.�v�Q��۝��hծ� �ـ�蓵y�4�戋�5�l�ɀU԰�ORޱc���@6��N褡ۛp�I�uoW-%5wC�m�����k����:C]���Uݱ�[u�u't�fo;�J)��6� zx6��7B	��yfS8�ř���[�\����t�m����� �˷c:�\�S��v�Tȁ(Kt[�pN!b��6�#6 \Fj����M2wm�j�<Ǻ���F9��9�C�2�LC�@�cј����s����-�QT�xY�:�����f�v�T&�xool���W��r�&���f�x�����`u���`Ե˻sgL.>�wz���a9�������9�{C�Ȳ��K�Z�:U�uL|��=��Q�����/
�v<d;7�xO 9iB�6�]wt�Cl��־[��Dq�WVmKzF`�te���)yLe��V%����K�Ϸ��M��U���繚��fٖR���Ɔ8VP��xRe��m�x[�����Ϯ��dӔ��$�ӫc1��G�v��b�19����󖑗�:C9s]ƴvs��m��60���=���ۧ�nor�����˻��wws��]����w>�뻾��wNZ�U�VV� ��>��u����wnM����HðAy3fof��9*ݖ�W��0SA6�-ѻ�v�Q��U���:7�2�*gY��1ze�^h�L�ዷ���`�R<:=�ǽ �m��]ض<�ˠ2[�0���*�F#�����]Z�tV�6'l۶�v�Ao �mQ�B�cZ	�&�N�'R��J{7ls��H+I����p[�`qk�.\qŻ:�cV�j0i�ɱ���(C�.4�Z����%�,R�f�^5��}NR��_N�6�T��#�����p]i��}�vS9��sSX0V�b�KkYն��x6��6�����M�v���k���<���;��������Wr���z�m���*g,N�@�b�"[6�;���\K��hɸ݆�4�R�p���N�+�=�I|k���2��Λ���W<�QG]��ɰ��$ �cv�u�혻����s.�q��f�weuh̫Z����53��k/i�[B�t�g�Ɲ=��}nnu淯-�H3Y8�Cb�3��j5:�dA��Q�&�ַU�9��XrrW���[f�e�E���:ܸoI�l�p*zr�Cu�Rײ�=բҧ�� G��ъWB�;t���弳Ec�X3e��Z:�9m��\D{��VQ���HS���.�mt�4��(WV%e�� 뱏u�ɵf���5�T�6��CK�V���Xu7�;h��ίO ��+��7�v\���&V(����g`��&qV(8R]F���L�ub�pf��r�k�3lT�q��m�:#8��@���X���]V�s6��ZD��z���K�����n��{ϵ�ֆU�'5���Ȁ�1m��ć�NPy�����yte;Pt�K�t^���*=�Q�f���)}�>W*�����sp�y�\�g>�!�x��E�����#���J]�L��w�o�ۛb����)𺎛�-�9F�3�ᕅ�3���1��,=:7AͶ����T�����㑮����Q;W��8�>�O�튳#̥��B�G�v��}��-�q�AA^S����Oi1�`팅#,�y��Ns���Y�-.����Jݡ��sL���3��m��7��n����a�ɢZ�`
繛�5�sj�p�����U�5�e] �i�+�:�k���J��YǼ�������]�)��xBR��*(D�ME\�Eef��;[(17������敇�y���oNn��������������7wwwwtn��Dh��*���1[x�`8�P�j���[�$�3B��0ri�MA�Ւ*L�n��ful���kpV����om)�4�In��H��]��'IY��하z��dM{���]8�K._[�-���|Xe��&�*�.^o�$�u�vN�t�Rb ���E��d���N�Y��λ�F�\i��pS�թ�,<3��uȦ2�c܅H�7,��YN�\Ac�g�Vu��W�T��pЦ� �����	�4�$ʁ.��M�-�*�c��]*6��s�����A��,�u��y��x��
U�Tj��ьv�K�ja�{�ȩ�\R��>��!l�ʬn�w,��>��v���&j`J��1��g,�C�Aٖ��O�wm�*�AdXp�P����R̜�r&v�Z��3~[vއ1�]S�f!�JoVr�;��۩<���C>Gn�a���(^\X-�
e�^:Ʊ�z��ʱ[�EYd��t��Dt�A^_x�wVT��=��N��Ҹ^�t���g&���;w�I+�|MtB/�5��Ac��;�9�c�K�����i��a���4B���9�˙���Tҏp�54 -�Lp��Ȓ�]���[:�(�]���\�wٓ�=��+y��eH&��ow!$���pt�2�f�l[��5�U��y&�h�z���<P0��tpT�H������k��n�9��u�6t=��ۖ�r���������D������I���sp�7pu���b�����]QPelG�&���ɚ��Ͱ�1mn��m�z)lK#o����M�yN�����1�p��i<y��/���(�9 &]!�W�����wc�Z���[��e2�D1�SPL-�"�ɗ9E`V�c��s&��nb�]�ɶ�lXˀ:{5�v�Ց��J�_*Oi.�Z�m���j6i�ڔ1��ń����7c��\c#Q��ܪ�܍�ٌ��%�B���)�1e�����j^Q�Z�s:�X��v�������~�̽��R�t�Wu>R��ť��k�� ���l�֟I;5p畜�ud��)ޙ���W|/y�O�H`�!`!u���TƜ���ޗ7��ovَt�H�뾛!��F^��/�h��m��{:��,l����&��9������9j黯0�Uؐa�қ�8q�.���(���'W��ܶ{��h��\_[3"�H,��Y��}������,��@�X�@�������U\��y�-Gz���Sz ypKyw�����f���oXy�2�+�C��7,��2NAM��x�ΨnX�t�݋��96�T���[6{�F�#j+�.�uѼn��7�q��I%ޱ��^Svt����;էh�^���Fw�!�2.i��nt�n�np���(^�����㪯@
���e��.I>�t:��9x��Q1rU�us��w-��5n���Y�]��t	m���t��J�3u�҇o�&ъ��k��ra1�b��=w��9,������{}������(���u��\���OI��׽��Ʊ��<\�r�T�ʺ��b2�J��n.1�\v�ZC�-�+*�R�}������;cR��S�I�eFo02(�RS��v�2&j��2\�X1�Keb��)�8̴�kΪ��������T����o��y�;��אWo.�7�*ѐ��^���J��������X���Sk���oK�Lۘ*�|��p����q@�06h�q�Ӻ�S���p�nVӕxK���CZܜ6���/{��F<tf�{-XUc�b˃#u%܂:�ϥ��l��b�V]*o*�1��u���[�u�hj�-�B��gfh�3x�'7r�E;�`��2�r]ٳm�Y��2�Z��1���97�f[��3B�5h�Z�����c�oq]#Y���9���srL0��O;Q�8eәj��,��D���0��3ET�XK$sZF�4�̮���"���΁��]E_\�of"wG|�BI�NLjRV; �`����K{p��&�7ru��]!.ٝ`��!�ǔ�{n��h��qM��h<	׌�L�蒏��1=�1�$��,���q�oiܮ��
�-={yۣ����Z��H�ʤ��-��n	x���3�#���,���4]�R�h�5�	Ö�ͅ�g+s{lReˀ��&�#wr���J���:N�_Iʧ��E�\��/� �9X�v�85�	�y�2�����E�)��4��Ë��f�[Ӕ�����Q['B� ����ۍ;1.��N���O(������C2�Z}[����V�d�U�nV��ek�.�+S�Y$�,LhLYׄXEh�K�n]�V؝�g\"�݀Êj廻u�K�ygPvvo0�ݶR�竫5GՐ�55̍��e�iZT�b^K��C"ٺ�u���y���\�Dm����9{���/t���	�wAS���M��;K ��)^wqR��)�2R��+j��3�m[h����<u�&�ۻ�/7p<$d��lܰ�t����Vef�K�y�Z.X�ڜ��;�F�܀wQVju����Z09�:T�Sv�ό]�ջ��s؏^�
$ �q��������i��U� \��Wi�r�9LvsA�,����K^uh��h�ا-�u�CƘ����N�Kw[/��H�U��{��-=�c��z��*Q������&�cAg��QX��j5�uv8nJj�H� ��5'ұ��F*��k����`v ���Cq�I��<������I�4�/]��C��6$�ƽ���Zp ��E�Qm̵�{nй�^����m}�F%�)��;�6I�U��wܥ�����U���0�[	��.$TMJ6�&��u�%��XtTX�z��m/�^��9ܻl��ʌ%=GjӍ6��),�B�:{�7�owu���j1d���Z��V���R�̹���@���;���y�"[�m��m�wȳKm[L+�V><+��̝��Z�:���[�٫"��w�f�m1�6YV3�@]k;o:*y��N���l��TVԙ����gfq6N�'��n��9����F���Q���WӨ�ƜՎd	Ѭ�˕�dk&֗꺝L]gU�=q����������j���>���]�.�}�^jcq�<�5�]I�������w��'G*5[җ^-JN���]ۈ&n��<iͩ�%�E�us�Cw�Ht'N����KkP���[V�]�q�%EM�<�vӑ�tp^����w0�Z�ww���zU��F�ʽ���(���jĴ�r��%Ap��T�d�3Z����}�ҹv6�*�geMV��[�r�PLZ���X0ǘ设����eӎ�8��j�V�7n`�_*\l�{�.�P��馫	�iA)�I9��݅�^�r��5\�Xő�q��x$�����7���"�(@��#M�|O#h0�l�vɵ�{�X��4V�F~�;��	�F�}��V�a�/�d���L�!��I{ფʝ����[��;���{B#��՚-��ԩ��.�m�	���e��䤘�{���(��*�FCa�<C& c�,�w��e��׳G]�"��h�����GB��au,�ʽ�YS����P;ȇZ��b�z�{��kk�a�TQߨAh�x̗���%{��fa�j��_`Jڸ���v*MG��u&�ZOv�2R�r�Hr��a�X��.��W�{��h��gZ�&�r���}�c`v\��w�W��̔�l�an��6�m���بW� �b��F��p����8���[��,1��&d뵌ƚ��G��Ò�L��j��O6�:�]�#SG)Ҍ�Lc����r���ǂ^�
����x��YL��/c��gnY����73�
��1|���@��{k[�i�M�sY�z�D��®tݝ�wrܩ��{�f[���?��y�nt���yi�m��)§y �w�5{�E�� +��0��͚%f��غ�F�m�夥��e���-+m,��Nb�����^m.���bKj:��w�w�^B!,��V')q�lqwf��6��-#���p����T�i֮�.��b�ZV��l��v��wm�n�8��t�0�d��[#�Wq�y�d�G6�I������XY�� ����B~ݲ@�X����I����u�S[u
.ˠ0aw8m�b7{Z�U�p�Lw7Q�ۺ���xm�f0��;��f7"*D;u[O.��m��[ڲ1W������z�:��2j9Nl�9v�1�����=�e�Ub�E�V���ھqu����Sy�=��~�w֗�BI!4�1��C_��m	%�@�D��؏�H^��:*�꣠���̥>�,&qz�      m�              6�              m�      �4ʷ�%�b�q�+k���mװ��X8ծB��fW��vN��gn�:�/<��n4�F�Wn:�<����j1�u��t�$��a]��:�sv�H/M���'<������7N�t�\i;]�%�*va�'	�툱��@[u&@�^-��HP<�z�aU�]�I�,G=�cd�n���bs�,�ۓ���b�c�l����m���g���cў�wm��Wl\sۭ����;������a����]��p�c t��lv�b�̷�+��	N��ۉ���&�3���Hr��HW<\�v��RWY�Ț�ͻyɞuE�u����Tٯ\�Xl�ͽn��e�^T��X�S�ָx�5^z{��a�{;���ɝ�d��7<ke� ����[�GZ-ڴ�-Pݜ��A��/e����`�����y]`F���h.L�P;vw������kPm��gY�v�H����@����e5;v5�ֺ�ع��(<hћ�c��&��(�u�|�lXմ���Ӟ6���B�L���=sJn&����=�[�v-��u�a��t�%h�.6`m�W���[s� z�moO�����ۓ�L�<�kmi���n�B�v7I��(�ۀ.�a�'6��m[���K�b��8�)���r���v����xD�n��ݗt��2�]<l��S��y�>��7;���l�.%���'�7;�@�s�'c�i��vl곫���8S��69���РL���\���u�햱l��b���n��v�Fz���ݻhn���^�:��N�x�S�G�C�P�'h�=��N�e�R�{��]=�]X�%ڻtWa�=r6�l�Խ�ݢq�sg9����]:^��X��c�����9c��Y�ڑ�ը�=��z�̆
+���q���GV�d9�a׷&��[vm�[��yx ���%̋��!�[)ύ��0D��Y�q���bF*�����[��S���ø�`ڝ�n:��j�G(ڎz�y3f-n�7e��D:)��E����ܜ��˺��a�A����m�t��hٝۮ�u�{u�)�s���p�:�I��v�N�8lS���s�Bۮ�֢<�&��u�ܰ��'
�]=�W^�t�ۛ�Z���<WZG�ִ�{p������v�u��wAVƗ�`:�u��YS<o<����qq�ܙ���A�v7��vE��t��u����E���1/;�s����֌s̝I��r.�y\<�q���.K�O8ɜ1ݚc��n��������ƞx�s����y.ݠ��v�<+����ke(Pݛ���OEɣ:,����}���N���g3B)�JV��kg��Y��p7h<�>8�< n�b{-�x��V䦄%��u�B's��� �ۮ݌n֗\��nK!����"�m6�;����w4\��Mtt�<�� 7����ٻ�8��츻m���(ے2hܽ#�1��ln�S�W�s�e(���۶��V�h�vs����/=�v}r���v�^NKa�ӵ2ݣ��q��R���HX7[<Q0��ny�͸�z;u�x����|⠳����ɶc^����y��wn�x�]��Ɵe�v����ln���8x�=��W�78��O)�������<�흯C9}�v�k��mӏYw����n5vB��8۞4�}V�{%�m�<�\��q��mщ�08;pk�Y�cpc2���۷/8��x���a8q�\v��:�`�8�q��;��뇦� c��]��]=<��=�x�]v���TK.�m�WKt�V�t��ö��K���s�����a
��Ԝ��ƅ�Nӓ�ܲb�M��:��曼U;Ĩz</w�>tH᭎��Pv�b�n�5�Ƽ��;���#�h:����L���z@�ݹ�o���W�F��@f��������
�$x��</^�<���ɶ��np퇷E��wC�׍��p��˛'�c�[.���:�2���u[�j{`RÁʯ7;�����9'�X�ڽ�^kg���lJ���]]���Yx��Fd�E��;\�[:qv�9�8-)[���)g>U�˗5��\F����4m��k�b^e.w�1�'8�[�OkGm�^�tݑ|v��O���t��&�ǚ�4=�=�,[۪�n9�ۍ��}&�5�̶����vt*��ӝ�KQ�Ā�[8A�s�������;�d�����a�N,�7��A'�]�W�g��k2�nL�Ӈ��z]���#F�+)\c���kp]��᫮���h���n����z݆6��.����x4�x�WKx$+� ��=�FM<�+-��^��c�\yci�\[�M�xZ��6�����+y�Sh�gls���K�(�=ks�ѹ���n�0�&�61���3��rWi��)\^n'Ά�&%�p=ql:Nő�����k�g�m�c��T��Qמks�E�y��6L�vz�.^��[��\�Wȥq�m�玫ma������Wd�Ț1۳�;��Y���Hx�Ψ�"ͼݳp��O�\Q��A��{=��V�^v�]=0��8Y
{C�hiLlsv����Y�A5��l[8|��¨���v����ڒ��qӻ��o�%��`����Z�O)5�Wa_..{6h�J��cnn����˽���l&�l;q�͝i&�e�N��=�<u:�|v��Չ
�-��>��GkG���ڣ��;m�G6;q�[��@ܧ,�8ɣ��l�*|�ѻf�O3ٺc�d=��sڵ�fwo+=���^�M��W�=s���\�ٵ�Zny��<��klv�7O[p���vpqC����v'twS�Ɩ���^x�8�fx�t�g���F��e�'U����H2�,�2�z�3��O7&�S>h7-���]�Ξ,ݰ�`]��gF��Yv�=YJ�U�-��2tv���\rgd
��+y�N׺�\��@���c�:�t�<�닡�Fm����Yɬ�D&�\��S�l�n8����:��K����/���Xw����������yɝ�ۭ��6Qn�NN�5q���e��mq����0���Krv�Gf����8l���'�v1�����E�n���/J�"wK;6���6��0�h���:�mn�la��xI�j�&��0��r��EFػ��^�b���� �㧱�9'��p�.�O=�Op��w���ú��-�]�lxWuMp����J۞89�c<[ZG���sM�t�`{;�F�T�t�T\s�lY���:�mgZ�st�Nu�"A]Τ�8����2�0]]��u�NsˡSt�l�YɝŶ��s,�q�:�nίm����@�8��Y�gl�z#7=��J�]�4QӬ�l2�5�㊲�\�u�V�-�;��l�݆���[���Y�ݹ�����wj�N�yy���-cn�|,k�lr�d�{s��lg*SJ�v닞�����ۧp\=���Ȏ%Ө�B�Yu����(4F.vݕ�A���nN9vT���伻oZ�q���K�X��p�q��G��Ã72����U�ګ�<;nʲ�J:Շ��I��V�n���7]��>��x����S�s:��A<7]�z�����8�u��h�w��ѓLpY{	������-��OPe�g�s����+фyՙ�\S��ʱ&y�64-o=Qr���!h�N��'A�dx�����4��l�vڮݧ.Ǎ��Q�*���0Z؝��GN��w�§bpZ2�n��z��dF�v3���T+j�u���W$K��=fR��_3�v뉊���&谯 j�Z;�����M=��_Vc-å����/V�%ۃF:KŮ��Ӕػ[��i7�:{sk����8�mh8z;[&Â�9�ثt�G=���Нuc���g�������b;n�vwm�&3��5�ݡ�b�g�kg���Y��u��!S��g�!�]�"z;F..��]�6v����6�^���䇯=-��z�������c���a)����}qK����Ux����\+[�Gn��1����1��Bg2f������\V�Z&t�y�ӎN#1I�h0^���k�n���\���w�u^6,0`^VYK�sz��X���8�	�y��j��y���NEⓘ�[��MN��n΢���V 9麭��8��uv�g!�۩JŅ	v����=;I�wn����8��0��{[�v[���9v^��I�`M��H��lc.�%�pS��Ŭ�z����W�Y�=����TlvFz�2��۫v�e��.���n�E�ț�Cn���kP�sd`�-֖9�s��oC�Sk�]k��Y"��l�i�P=�\���v���Wa��       �ϟ<z7�N�K�
ad'�G
�QG���&AM�됰����!�ܠ�\�77|������|�D@]βed���:!q�'κ�<��i��O�v�D��촮s���ț�US�"�:�B{��:;�L(%B;#��^2��f���Nn�����؊)�/�C#\�6�;*����<�U®R��Rr9TQW3�N�i��L���i9�q���ȗ�N:�E��z���/]�(�#ԛ�Ip�����ϦUE�w}�	!㴀�S�p��9�r	Aɹ��-D��d�
��Hֹ�U��e2�/8*��Rz��=����*��.A �S.G(yYTʪ��ț���L�I���5�gwY��L8�q�(e$'N�]�P�PQE�3������:E�*#��ȶ��_(]�m����?����`�  �  � �s&'i�7)�]系Q�D棣V�1���|ݾv���jK�W���0z�p\�I�`ܾ�tN�\#���
ov�r��Z���خ8��G6�V�4����a�v��@���a��ݹbM匛s푊w/"gV�u὞:ƏU��{O�8�n9]\ZP7�=�'��W\�L-g	�%��	��^;i-��N�&-���l����{<�Ȕ��	v�vy{��)v��wF����u�m��y�M��.��0֭���j�v��{h�v�s�a9��+�Z��S3���8�1�f����[��NK��zf5�ۯdO<�ˀ��<J+\X.v2�q��4�;p��\�Á�7W]��kZ�<Yf���7E�k������w��E�3��6I��؎�>�k��Wns����si0ۃ�v�l8x)�]���@qۅx�.wΣ�<m�Rm��Uؑ�q㧗c��n7%�-&g����<�t\��p�ۚ��������#�s��5�h��{J��J��/��:}O<�W��͞wl���A�n��t7��	�rJ\k9;8��-Ɵ<��fдͱ�a�m�qۜ�k�`�m������m*2F5$�[;��9\���{��C�x�k=3���tޮL��D����nͣru ���[�d��v݅6��i�̏\\q�1ۜ�σ�w�s�'#ϓ�s�+���.�{h�����8v�u�m�A�l�nBƽn��2&����y)�3��m���K����퓣��FݍqC[j�N�x��h�N��狷!��c\��D���8ƺ4r�i������O�olv]:���OR�^��.Z��q{�t.K�^J� |�'���o�UPO��۞q�l������y��A�;.Ƀ(���;;��v8�N�|vGyE�\�����#�R�;��Y�k���x����/GKے��u��K]��:��.G�x�"�0��1���8^0�<������s� ��t1�\Wn�:�,�q�=ڇL��UL��T�(�\��k���K%Yc�*U���/�mm#۔&�I �	_D*'��8;<��Sр'=�S�Y���7�R�E�F�$ 𛽞v�%uX�\�H=ڜ�I$��I����(�<���A	u �%Ʉ"$�d��٭	$�v�H���2lMJ�}��'�z�ЃTH<�&3�4:�J话ϋ~��"/v�sM ���pTH:d�I$g;���+G�
}	�u�4g��n�7H+�J\$Mă$v�϶X��P�&ɰ�=nf�A$��tK98* j2��D����G�6�ݣ�sn7�ki��H�جjd������W7d6��Ĉ�%8I4H<�2�$�{dw����<'+��M��P���tI���mQ�J��Q2v䐚��52W�(�����q��R�t��E��K^Ugc�X����2���%c��%�QY]�m^��w�5�-�� S{�U�q���i$��Ψ�^3�i��ԨK��wc�X��2|Hމ�h���eX�I6�u��a"P	=ɚI���6��@�	�0DD�n���͑]=z�[�t�ğ�{�I��_gnH)���챎^E�ĳ�Mi��J���Kf%L�S�3Ψ��G;�B����c2cI�rf�K��#_;� �I�v�6�_��b@��w�
6�y(Ͷ�{s�V�y{qq<�J���aoq��M_�����=��A]�]~$9��$�D�� BG�ژ1������ ��ܓ�.��>|R�T.�����8p[z���4J	'��v��I-|扰���F6��y&Jz�֪�R�P(�>=ۑ�I�N���$2*ިP\dTN�ҘYْvf���dT����9lS�Ӷ#m[.�5$��N�j�c��u�l�0ro015 �څ.L9�^I��l	D�'=�S�O�'DUݎ�Ť����a�o�D�����>4I'��RQ(�\���G�2�dr�k�'* �G	�"$�V��ͺ��H�nkԫ�"S��-h	-ͻ�	�K�\ݢJ	s��	,�kow��Cp�:T�L�*�Unjn��}q*��r;6q�[��"-Ӝ�]>�{�����4��G*��v�H$q�&�Isɚ	I�>���>��̒� �ڤ'=s�@����h�5?�$�F��z�
Ӱ�s��$�#;�9�'�M�ę$�A'�v����Mze!�UZ���IA(�d� $����H�VT������H��sD�	 �ɚ	*��q""D���J�v��~�u�ʧ�@${��­�%��&�^]�슜7OE`3�V��xb�u��P�@q����������UZ�}@�wL�2į6�[���J�4�k�i���ÙH//�� ����9�v;��G0�މI�&gk`��6�>�rgQ&�G�BI$��&�Ivs���Ύ���p79lr�������:��"��Tnc��,�<�nӬa׶�sM�:3z �$DI�#��5i$�m�RA$]��ɆM��
8�Ժ��$��&�ؚ>F� RTW�yE�l�	'"����V�yd�p�$�=ړ$�O��$ �B����R�;�9!t�@+)K��9 �$��\��h�N�}��C�I��M�� ��{c�L�<��Ti,H��$}�eF���잻���I$�;��H$�Y��/+ P�!�$	�I�&����Wj��D�|���Iy#��k���-�K$�Ι$�W���Z�	%��6-H�;z�񌁙����#�'9�Z�) ��x�j{(�-�;w��v3�l)��,��^`�)�f�:M���I$�F�UB�k�q��1xΚ��۷V�V8y����޸�v^5�g<�x���S�;)��b!m��X7��������.��;g/G�|~|p��㰯T�gc4p�a�b괁R[s`����k������&�hٕ1�.�m���ζ�s\�[������MukK�����V�+֎*A[�)Q;�Wjмv�kѸ���;m�b����t9����		v�������]�z�ZI�H�D�%ٙ�lO�$�9��"L<�ȪV�wa�*�3A$���Tl*K��_�I
�B��H������4/�6/���J�9I ��J���6Iv� ����!t�b@mig�C�)*+�r�~��$�#7� o5��y���`$�H��ݢa@���o֗��rB���+���$M��m�"u�9�`-��|ߜ��I5G{�HI$�D��U��~��x諻�9P���Hj*�PTM�� ;�Ϝ$�$�M�0{9�ld$��ݒM���شW�Ie��$MM��w���fu��*Ŋ��n����U�k��C�y��<�� Z�:į^��������T]�|�7^]I=ۛV�$���%�n;�M9������$ �ojbV�s�|	B�I�$s�l�'�Y�q��c�����Y�#]��3��T��y�"�}���W��$;ok�zO���ʙ�#Fjzs�Du庯�$�I.�svI �_�$��Ņ�YO�\��(L��c�&H�B���{98I$��tI�n���a�{/��IГ�sD�~K/�i$7"�=%L�S�
�6�m�};�;Ē^>��H%׳4] �s�R����XI#�w���z�@]�A]�, �,d�Oku`Z��z�D�Ө�IyD㛿"'g$�$�;=�}#�]l��F/���i֦�ir�=ظ�:��v �p�[n�\�d۵��8��
�V�ە��UZ����� o�@$�D��
D���.쵼mc�0`{[��s��T �&��NI�ѣ�R�U@�\>��!5D�I��m��-[;��H$�]nf�I$�9݁h��M�CT���u�Bi���w�U�RH��#_'T����r�4I�v���l,�L��<;o`dw2i
䅧F��iZ�4A$������ꁈ'I[:��3�	x0͑�ol�o�I$�>�J*�=<��Ȁ�V�&=�d�� �<�ꘕӻs� �$��9]5H���3�����$x��﷽�~��,��'	��d�,�4hj
�_K�[��}�����Sdς]�3I$��uD�H-��q�m�^����K� >��E+��%�4j����z�u���N�t�#4|�=�>�%�T����'u�ɡH��suv�Ir�qW�"8�c�H���M7ۮBkfREU�I �PO�f{-ω�)�O� �ćQ ��wi �K�y��(%)T��-�[�66y*V��hL���%Cd���̥	 _�N�6�n$�h�}��>�I����'�'���_�$��D�~K/'7�M`I �Suv�^KnEXW�H�^K���8��ѽ4u�������sC4R���8^Ҭ��Ө�o��#z��^v �:�QS-J��"��O!�K�/��֐�\��G��1A�x��}�$�75:fU�L�r�������B@'׽�!�_e��$ɻ��H*��~}ϝ���x�Q��.���K�,v�������>��1�;�zI� �	H�H���hU�R6������N��� $�s<�&u��Ԕ4mI/֊�E���i��2$d����H���ɢNr��35w	�����I$��ݷ!$�3<�$���}m�)�����c�2��UZD��&fE�%��H)�#jf�c�#��u��I=}�r~$��ԟ�I�t��$�A �,����	+BXp+c"!,S�bmy%�|�i$Ks��+��m�Z���߷.C���߂��$��D��H:$�3��3O��bV�/I5��ې���9�Iy$�;.Ū{�ĎXk��]qB�Iv-q��P��mN�K,�yN�_7xN+���������*g��R�h�2����az:�H�[މ��|���I%Q���"����Vא\X�'ogb�<<v<���C�p����z6����}�V��od��t��uI9�[*K�bwn�Y�������(���&�٫�8�x��>��о,�O^��Z'��8;�!=�M�Ol5�VrS�;<��ҕ���������*�\=����"6��aL�g�Z�;5��)Qb�k�����f��0�u­��.�f�<z��7�w�����D�� � ��ޱ6J�Gs�%�˻I�<��9ִ;�[W�I��[�Mn[5ƅY�Fе�^��BIG��m��i$GV��H��eݠh�t=�Z���o/�]/�
�v�
�)`"�gȒ@�n9��f�����!&�{U�I#��ؙ2��*�D���(�}��	�Qٞ�y�4H��h�@����h�����/[�s �I��V�\RA��E��ۑ�D�w�|����r!�[$�O���5G/��*�W��%�g�`�M�X
�C�6�0#��֢�j�ޛ���<Q��g��������q���I#<O����_*W��`}w�{nBu�޺W����}k��$�7��Ф&z @GD�1A�KU�����1�i�����2��|�K8*fz�;����Er��_p���kW_-��^欙�����,��N3,}��*+�@5^�˻H����Ţ�Frm��C�t�IrF�а}H�-}.|[��	�$�:}�A"kLeI�w(gG9�h$��yw�EQ$������>�Pj�+��Ϩ�g!|A�p�^Jf��Z^I�F�$�It71��=����eB%�λ�c&|�֨�I�R�!0�$P �jh�R؅]�I*�wv�	�M��Cs��������bb$�B�I(��B�N;	���f`��������q��}p�'�o'�.�h���;�A$<��&��;��.�U�l�?Oj�3�c�V+��Dд��D��N�4L�����^v�eQ&��nu���@.��	�Ί��ϣ�᱌y��
�m*B�
Q'3]�k0��U=�r��I%X�$a$�����{��~jD�+��/��<w��Q�Al�ںK�n���J�RW�s7fLͬs.�V�`�Zh��y��a�Wd����\�����������	ز���O'�z1+k���	���[�5���̚/:�E��<���-:�pf%wz�$�eSׅ�(d<�,i9tбV�l�U)�Ood�[�3q�����Փzb�bh7N�b������Qkd�q��{i��p{/P�������s#+��l4��v��)]�����T�B'f]��' F�hqfr/[��7� ���8e�8a�8�V������ŵ }��i��Vس��+
�,f�jՓ������(>ӻ�/]��*�8�F�dǞ���w;vް�1
�\4��#3� [�gU�7qdh0����.p�����)�Ocs/l����ٹ0va���b���opSؒ�OV�Ē��me���E��f��Q��:��U�ab�r'��h@w��ʓC�Roo�YDc�s�؇��J��Jcq1��!�����6ᒎ�0r(�/ (�QU����ȁr:Z�d��7�2՛�u�i%-:���}��q���(���
����X��"peӱ�QnP��XsY��R=����A�M�Gu�4�!_])�q�R7ܵ-�f�]���G9��̠yn�|N�k����͝��p�f����� I	�~ ����J�W(��t�ۧ`QE~��t�2"�(�޽|�����b~$��I��yDȜ�U����*��k��w2���Y�CM"�\.��E) �#��Br��;ӷ=�ϯ�A�Dr�� ���9C�:��z�q�=�HH�rS�n:�m�N�w8Z��2�'Ud�I�)�k+��T�uyܝ�Г��1R�������w	��s�7]��5H�Ts��.�\��&hS)���Yp��K��HJ<{���LIP���NEt�f%a�ZThD�g�Qj~��\#W��OW����+�'OD��<��s�wN����W$2I�-��$M�5"����l�5�om�$����jŢ�I}�BT-R� ���Q>��W;��G]΢I��XD�Z�(~�IB��\�V�?�K_�l?Z���HBb&\0�+sR�I�sʱk���3�X�^	 ⷢ���'Or�H�w$���2u��t(*p�q廱�t�Et[�۸+Q�i��H�جf�Gk�8萦R@����J��؛A%�_Gl���	/s�.�%'�]Ҏ��ׁ\f��P�I���U�MP􏍤J�e*(�~ܺv�H���y��7�6��(,��`2Gg��D&��M��w��g��)c�]"��i+xOD�D����T'���.]�s��'�ߌ���I&����d�G���Bh����'�nС'���; K%��B ��XuD�}��O�$��<�]țhm��IM���Y��|�5�(�2T˳��q�`�ɱ����2k�j{=P�s��Jw�����(<�y�ߢa~�Y�@W�B@��]���?�O�$���.e|7+²�OΪ$��e y�� �~3W��J:��q���y[vP)"�C�)QHG�y�����C�bG�<�<� ۘ|�}}}�y�tv=�ߐ�f�����>�����y{L��+_N��a��?Jо�ɊH��w.�~������@�
W�|L��'�p_�S1��sP�<! �O�TM��:y��������ťng��cD��>��nՠI�_v;�M��}�(��K�0s������$����%,��q~�w
��d�bf`���1��1�x%�=��Ќ���티�	���_vG+�_�]��y��P��lo�F�
�ױZ$�hB�W��3���< PNxe��v�	 Ѽ��Rϥ�'C�"�����7i��|��md��|�9\�q2�0�IEnX�|�G6������qDt�v eL	.bK�, �F��>{��<�y>}z|�v<n���o�gt�c����U���&���[	{N�eNک��� ���ν�.��7o�e��y�d�k]�/Yʖ���=v�������]WQ�Sc=�j����`�m�n��U�i}��8�N)7�CN"�rtח[���lEn^Pp��4Ny;k�m�ׄ�qH�j���k&kdR�.:ϟl�ܜ<��y����H�溻&�7=�ձ�.\wn��z1�������1��9�I$��si~�\��vU%5��T�80��쑁	4r�~�bV;�H
�Th+J0�DeQ>��m���f�xw5�  ���M��t�T��:�c����P�>{�_�͍=3�{j�� ���	�t�_�c�_"'�o��~�]�Tv�Q$�z���Nyj.�?s�n����Z�����rhnq[��B�$�(�%(�I��V�$�;=�'��
����c�4]��RR"��$I\�OD�D���� �
�?iI�'��:���D����$�^]��ũ���y*I�IH�Ѻ�>���l�F��6^ՙtІ�&w^W���S��u2��I�$䷣6�גA"�sH�$����(��*j�U#i���V�lŤ�qH%�$�"fb'���nŢL5Q�VA���=M��Pڙ�p�PD�v%&v�]ЗW|�u�O��6Y��D�ǨVވ��S�����$�Bc�"N-u�?{'2���.�!y$�i2Mh�?l�B	6g_uwy~兏����@j۔H���d�~'ݺ��"K�Y���������	Ok��$�G��$&�g��eU�A+�Q2_�/,]s��$�'�Mz�I%�]U��K�:y��������$�N�HY�=��V��bA��6�k���A.�9�_è��1�-�$�;d�I��]�.�y{KfU����m{�y�:	"l��Y@�"���-ٍ�B��um�n�����)��n�r|���w�Վ�Q��m�RA"o9ՋI"W�g��l��2��rĢRԙ&��}��!	4n����'��-�U�&�gz��) �M
I"~��$�Y��Q7�F�=P��Igĝ(�5�W��Wk�p��%BI)7��i"~Bk0���E�O}�oޠ����2�X"2v��*6��f������WC-^Gy�n.Ft���J���xf�yS��7�_]���I$�n��$��_�ʄ��
�
6� �\r�j�79����$��͈n��&�˰�TH g�&^_��F�X�s�IY�3&"QELş�D^Ge��^H��&�pҙ�z�t�pI{wv%�{����IՉ:$�sq��+F�nzs�-B˭��uVu���ۍ��k^ _D�L
�{�(+�nժ��=��Bh�=��  �9�I�OY��:�eC�=?ee�I�q��,ZB�j�����N�S$���#z���'uڍ�8���ʹ(�R(�d�4Rp[gQ��s��J#���*"H7ir�ثH�[ɓ@.�����ޕ&W8��섂GW�8�Z)"_ؓ��^�d�_��RI]����gE��w��^JS��$�I��&�Ky���� ���iX���iǁ�R��ix�F|n8'wT�v�[�\�N0�\�{��*ѤHP�Z���#��'�#Oo\�N�߂��� +W$I�lZH%��:;�v��ey$>��X&�J��Ā�{vHf%o�,���(%h �&�u���'u�ypٞ6��<Q����ݦ���?>��HT	)_��nI}��I)!����}�]�h�߯Jq�*'D�b@?�M�#v��j�"J>��Ī&���H��'��Dֈ��"-Ꙡ�	 {ےB '�r�����q�NLr�޺�&f3П�7I$�K>ܫ�J	v	�/l3C�7�5a ��K7&i%�[�.�%R�� �:%DI���4\����M$�;�5�H$����e���Hܿi�e~�2[�Ā�D�'�$�+ԒWk�p��Q9��3�vO�M�#*X��4L^I�$�G�� J�����0�����>�:#�݈��7Dj�Ôna�wɌ���2���'����ٲvѡ���Jl9YJ�ݰ�S��~?R��~�	���Aggi�է;pM��"�n9�y�0޺��e���9K����#	��򋃋n�vr�\�m\]��v9�����4pH�nd���9�Д�F�ICpr�3q�+��r��z�i\zz��n���,�n�M��s�ِ�w0Rv�	���A�N9�#�����u�\���Y�d�p�k,������\���-�ŷn���0�Mh}���F�>??������-���w����$������I$���]�#�.�ӝ�b+���V�I;ݑ��>W\�]��W ߙ`s���i�o��z�'�O������D���_��A%���
|eX��;���ݫ�V�Z�Hp�{# B{��\$�7
�����"�'�7�HA�������Z����bB&f*�.#~�����5R�{�e�Ym��	 ׹v	?3ר�q��v�쎉4^d��%�+��<%DI��wFm�-$�-74>���`�D�wp$�o.�%䗖���+�$�;�~po��m����}��ڶk�On��w*�t��k?7����[�ؖ*�j�g�`��_���c��w�k��B~$��~���>�n���CS3�M��*�ۣ�g�%�O5b��/���B����p�''T�'����xw�|l�gv�2Uʉpq]�� ��-ɞ��&5n�K�W2���n�1��Sp��b��έ&w�<���x�{�<��j���%��dY6A,��k�/$���~-���Оy��J�P$ڸ!0Η6I$�s&�A'���Gv���mb���;�_���I_�d��W;��*bbD��b��[���r�ry$�*�bl���)2M;�\�/$}�g$�s��B~�:�Yt-Q�i+��I4L��C0,��u���	4�m�I��E��`����7wi���(<������{=�t����i��YbWED���e���hn9���P�A�KV�\�H��sR�I%���;=M��ӽ`W�,Z+�*�׺��l�k�W�R_b
>{�w#��9Y9">�>5���M��Atk�&����TM���t�s^7ZU�}ҡB��<�a��"h�D�ۮ}	��O�rV���iC�HL��d��9A�g{�ݻ!X<3x^r�Q�qi]O�n��:��'e�ӖϵE�s�{�\�����G��> ���$��8�0 ?�������~T� 	6��L3�#���EQ�d��d�I';��D�F��/vSrd�)rN�4��I(�V�$>��!4I'��`Q�g�d�v8��'�Ozf��A��v��I8��j$�������a	B�L�Eh���r�L�;��^�Ć�<0[����M�������+���Gz$ L�lBM~��m���j�TO{�d�OglbQJ��t_R��(ID��t��U��, {�:D�	����"K_|≰��d�P���Ԁb�$x
�E���_� �N��� ���Z��~$�����!$���q`Z@b�وA2A���$n�z�H����Iպ���[}�v��I8��U|xR�6���fߑ0�**�F�RNn.nr�2�6�έ��p}��ᶬ	�݇���u�ר�M^~��OL�Ap�UUr*�l�|$�}�q���Һ=e�X�q`ߒ����$���J}��
�j<*��I$u}�.�^Iyd|�	��1c\~_�������Cm1�f<�g�aq�]�q������f� R?~�HY	ZJ�#W��ݹ��$���͒�Ad|�)-oIY;*���,"h,��v�	�8�i
����*d�bfb�k�\��X�c\�����%{a󋰒�H,�s��ﾌ��F���VQ�'�|&"$�y�Dq��`BF��`J��ն��޿u���ǯݷ*9~�l�'����QI|Ԣߺg�%�]�'�|c��?Iu��'��UR"���:��U�'�/ܮ�)
Z1�&ɢIݺ����Cd��n.�$�nb�H$��;� ��V_��sB�5���hf��l駪��/qCN�u'L����J���1E�i�7�u���z�T��A����W�ٙgYw�:�I��Ek��QA�N�X,-8��μp�]yv{u=s��0���f佮�y�a�7734u�^��+Y��K�w�Y�6V;�
%��o��m}Ry��.���N�)P�xw&��^3v�A��18��l��6V��1�ݗ���/Өl�@���j"ȘcT�%��/2]ci��}-�ճ"ٱ�ӗ��pL�*�����	g)���P7c%�r�!e�kF���\��ܳ/���&X)W��՜­��iy�˵�op��J�������cm��RhL3Q�&	��3y��5�$�}�os��3I̹H�.�rM�x�Cr��ۮ�����[�r�XhD�hș�s�cZ��j��$���8K��  �Z7in�#H�yw��.��o%���,�X�Ӻ��us�Ք�JM�cbN<�]l�;%��v�6�;@�Ֆ��6��.�s�y�Up�Ϋwz27�-��p�Y���Ab���H�l۵�u�]$�Q��.iln��͊�W����H��uh4wyU:	tiGV��d\�6�񸩚k�l�sB���ع]K��*�{X���7��u�5up����{ڥ �^H���u�v͹��
^9��OM����lt�<z�u���ސ�#R(F�lI��Ω�V����O*6�Q�9Ͼ8����>��=;�3I�̥��P�.�өm9����S9t��瓆0�1#F��Bwqq�P�3K����N�Y�ؘ���������*'J ����r�x�K�	Ҳ,ʔ�R�,��<�s�ȶ���wzK�\����w���r�*��B�����Jw�'TS�?;���Q�PC��Q���ͨK��鲢�����VЋ!>$u����z[�字b]ΖHE楅˒JQ9Ĝ�	�d�L�c�	2��<���x�#K��N!<yS�"*�'=��{��4FjW
I ���sC��{�y$�z����        ���6�{X��w��q%��<�N'�C�<8ƹ��^O4c��pthz�{7&�'��u����g
�m巼�n͌;8;a�nN��!�&Řԥ�v6�n�ݺ��=��ѡ��=\n�3u�\f{3��˸U�VǢ.���vxۍY�<A=P�Z���v���wF�qA����͓v���Y�\��v��uF������;&�۰8����ruO5��+��t����b��Z:�Y�[���!Ɗu�ԝ!�ѝ��X��C�OlpY�p=�g��N����/@\5�:��dc��#�.��K�������=��oP������\�g<�랬c=�HŎlY㶺����ҝIa�sO;�z�	ѹ�S]�-�ݞ�*y��n��j9ų�g;=�c�ۚPj� pt�qy���ڦ��v4swbӜ��wn'��p��W`�ۛ��A�]�Ѩ�-v޽'��Ƈ�s&�GLDy������ŎB�:�մp�i�&(�ӧu��z��瓬��um�Y�[�Zwg/�A��r7k��g�#��.����v��p6�ɞk`ϵ�M\��
7/l&�٥���5�z,ی�ӻY�]��[��wd��f��w׃��<G7[��@�z	(���ٰ �˭�p�{s�u�����m�����1��6w-��q��K�m����4���@�5أ#��tPŶ�u�8�vv�m��]��j�����n	�&��:{�-��E��;���k̖���W<biD���eB�p�ڸx7�qPOKu�8J3v9磉�S(�7�uq�..v#k��t:h۳��pa��s��<y蛭<�ƶ6�������mk��9�ڢ��8�\G�����z& �}���'�zz� &��U���9^�:0B۷�8\s���޺w���{�4��yMƎ1�CZlb�O<7^�J�䃝��_��w�>|�j&���J���x����\ܥA������݇K�i�`c�縕��b������6�ָ��R֡��Ŷ��]-h㓇��H���[s�[i��i��- �����4�|~v�|r�g����f2�ܧUƯt��	�|t�=��j����{��v�*�$�����3<�U����ww��J��o�n��VB��{�[Ͷ ���U�$�~حX%$�@�%vd��t���5��m��A$�N5�I �9݋E�lh3���h�o)󩝆-)��]��4H���}�O� ���\� 4���wu�m��H��9�PIx$���O��<n��A]�𒨞3�z��yby�˾$�4���$�g�d�I{�q�^{,�ȀQ^��-��ub����2L�Ν��	5�����BX"ɻ�K�bnb�H�>uE+Y�/֡e�V_kѮ�;۶.���h��J�����Yx��l��ӟ:�<�ۘ{��}{mӧX���׉Z�4%/$Okub�_B-w۳l%�-��~vtH����,$�y���^z#��6�m[���"����֓�Ћ�o�{kd�Okr�]�����\�U�حu6'j\Ա�-K�٠�d�}1I��rVI�Y����tT�%�&Ą�ϳ\���+w�vI6�?~qb�I7tDu���%{D��ފՂRI${2O�	$�o�~I$~�IQ�f	������A�M��RJ6(��)A$����f��6Ft�D�I�z�'�OĚ=��(��ڮ��w�#�u���}�l�����tr
�С�H����?8�&��5��4m/��U���-�Ma$�9���}��6�Azc� ��B�!#��.z8Mc�ѻ1X 8��sun����ϣ�yɿ-a��S���Iۖ:�<�	��RQ�߉����nů�BA.��6-&�F�B�+W&ɢ~'Or�����/?<��*���G7���D�9~�`2fy�`o�/\܄�ϕ�!@m\�#{�`U����#���I`~���Xm�:���M��V����F]*�R���fX�8��H�x����ʱ�^_<��"�V&�,6�j�  �|<<H�� ����%%��ɱh�����	�e��M���H3(�{#W}���ܷI z;�V�A$�9�A~��n� l�?�h~���� �6M�9�O�D�$�f�uL��]bu�:���ω$��Z��I$�۲C��-݇4�^��`n�������OStv�=T�͎����msU�|4�P�3A��� �}�VI'v�"PK%��;=�	���$�	�r���XZ�7hSR���!?��Qe����8~$�Or�@uD�=����K�i���t�2/�b�}�{��Ѣ��&&.�ʮ~���Ik쫴��=���[���t�Kɹ�TI%���Z];7�~E@m^�H�wn�?��_�$�l\�I$��UXI$���-���N��n�����T�1aݚ�V㍃�6^3`_�#X��P7u��{�%=�w�b�\���j�S�A�����{�6Ibv|������x�swu$����@���G��Fw�G�Vn�˿�K6nB��Iy_n]�Ey"s�&�k�z������������ܒ����Us؟o��Q;����m*�����u��A$�x���E$���w��I/�o���*q�g�Ư�w�r��@?Q��$%�+����B��H���ZN���s/��D�{ݜ�p�$��x�B.�+�钥]�����ٺ�P�v�E�щ���߽��o�ͻ>���\��*"�'���cI��)	�=�ŃE|�V�0�[�wv7	]}V-�:�&��I��V�v��ޫs	&{}$&����JV,W�$N��&I#��N��t��Jg�I��H$��R���ڭ�6�wS00Ǖ�@y��im�7����HhJ�4��8�XoK	�d	����`ﻍ���1	险�"���g'�{�{'R�$�� � ���7wwwwePEx�f�g��j�.��m��;N��sx���-�u�u����{����;[!״�=m��/F�@�H��2V���j䠦�[��<��՝��%���x����v�n��\a���8v�l���;S���ϱ��nm��Ɯ�Xu�ۃ�3Z8���綒.7�lp��C�i�Ps�\�+<���e��Y�X*��-+�5�#����� �'����wjïSb�����Q �e"@ǻ2HI �m&I��>�`j���M�}�h��I� D��T��v�Bk�B�M�0?��I/-��z���Z$��󛴒Ids���	�c�1U�rUBi$+�o�,ݡB <��NגC�ۚ��I!��uS]Xyv_$��IE��s5�A�K��!DI&g�GVv�y$�-�2�*�A%�\�$�Ivs�G{���u"z���V*����q��ɢ@�n�G�D\K�~I(깻	/�I󙠒Dv{[t�|\=���%�I*ͪ�#�o����*sc�T���	ܶj^d�3{����{u�&��cO�������H���RI$�>uV�t�m�W�#�(%}4M���Y�P쓻HIY� �21ļ�쩩_�pzb�	#��Ք4u.�;z���yi߹��z<S�&�)|����7oE��/�
�O��C%��������h@"����e��;��I!���I�»��.fOr�y�֒�h���D��H2I3;\�@4L�=����{	�t��"_�3I{�uvM4�~6I�B�� ��˚wK��@�&�$^��!&��Nw�N�cH�Q$���$m�X���7hTR���~��$�ܱWu's\ij~H��$�m�?Z�D$��ش���Ä��tEs�<~?\�»vӷGTV�k�g�i�^�Lg��q��IrJ�tVh/��+����5D�}��6�Y��d���Y�����e��7\�v^|����dڸ'�������,�u`�_\ɠ��K^��H���"�KYq�Bί�ƥU�T���f""Q&��:ܺ6�:�e��PK,G"�{��I</%s�TF�Řz]*674��i{��-}zr��L΅1jY��O�C�W*�D�~�����@�1|��I�o��p�T�S��T�O�0�B��)$d'O��^�!�;o]Ʉ�Q[�b�$��"��$�.s���c���&$�S�$��wv�L����".С'���p�ݑgu:F�:�M(�;v��%�[�k�	��1A'�:x۶�sC�ʫn�[�㲝��V{,Y�����������nM&չW\�"��������E�5��M�� i�e�I�M�j��J�s�y�读2���N>��+��A|���r��g+��еrx��z�UGS˦-��]���$�Y�)$�uJ�b�`d�o1����d�l��V�2����I��	K�3��[ݗ�}	ytol]���k�1U]�&d�H�� 	�6��������(BH$���1^I$w9�U��G���[2���9Vgtx�_\��.w'�'���j�/\�n���_QI���ͭ�q���-����I�d:����{���G���I������yYY�1��c�;.ԻH�'�O�I'�fk������[|{�D@��ػ$Kc�1A%䗗g�辞W ��E&���a�����k7c�V�N��}���^ތ��HW}�}n�_Ό������{�V$��Д�I!��앐2&kuV��9�]�P!/,�s䐴d�,m]ݡQO�~�*�%)���=�Yrt��I$�9�}q$��n������?�~�_���\f���D$c�	#<�f��H$�K)�nn���+�I$��9�P	 ��n�Z��Dh�LȘJf(�J�fOwOT��$�jnkҒH%��������]������c	&Z�l��&� �����@?/���4I'�~˛�X[µ)��%�]1^I ����w�Ey#��"����NZ��etz�D�՛��������52���8x�����?�=}�eӛ�\x�V��JʾʾNI�u�|i Ch@����7wwwu��ہtn�>۪�;ν۞�m���֋hc��qtc�qX=�k\.�ùqm�����%��=8�<�R������gU�N�\���_V;)N�jή=am�k�=d�n��Ӹ�^1Q��Vc��]���/F���nN��kE�9��Q#��#y�J���L� k���/M�Ѷ"V��0�(�z99�\��S�����f,�;�l;v�p�nx`�)�	RK߿_�%�I# ��"I?;u��Ib�ȫ	c�)ޠ�*a����ي	~��]�*d�P�l�""H6N��tM�Zù��L���iͺ��zN7�_�����1��V��P`�whTAy�߿e� q��$�<�?�x�_6*�4$�K�f�wh����ȿZ���n��Q	��K3����>@�$���uF��8�dU�����R�o�үn�������}H��+%+�zLP�h��ښ=���g_�� ��ޒ�I%���FU�K#��$�d(ᵋ�ؖ�[Һp�����+g���-�s���nG����=��ʓ"Q%�u�����r��ͯ$��N>sB}� �6��wv�$�����%F>$�$��D��NR	Bt�xv&������M`�1;x�'�l+;G�����ȯJ���NaV��
+������.����	��Ńo� |b�	 �5�s�䗒_��ȻIy#��'�]�S;���Szc������0(1�L�� ��_u͠�H��ץ �	t���#T^���<H_.�P�D�>�`:�!�b��ڳv�Kϟu�Wvt�'������M�����RD����f`d�Ѹ3�A7~޶<|M�_*!"��\�Iy.�ubЕ=Yй�'���4�I-r��V"	Aw۷~�[	�	(���u�ѭ�Za���4�<�᭚&�v�/#le}{���DZ��)\ 3�z�C�h��^�VRI%���Ҕ��o(K5�gWS��W�ST�s��5L�k̶���wZ��庺r鼢5�i�������Z�i�5L;�s�������S=Yǰm�0�
CT�4S)�h�����j1e�TҪ�}�ޚYj4�Q��{S��9Y�^���5�"��J3X�[3�Yi���Zj4Nz��vҦ���5J�T�{�����z��e4ST�	А�y��Y�랚aSv���|%:�Iv=ְ�gt���4A�`9��)[:�@�Fs�íꊲn�R���A>Ug�'�,hoTR�f����5��չmn	����v+�ޝ����8M�κԑ|@]zVI�Q�i$H/������^��g-��&1�]:�{$9̆�f���]����]���-�]�+6��O*�Pöe[�o�[�iV�Yb6b���"��!l���є�2V��{���C�;��A��U�n4�����}v��*�f���v�fRg]7-J���**�T�s���.,W�l���<�t.�y�r��9�zT[��N��U��a����9�q(��J���ػ~�X2��`��:�f8����a�@^r�}�8��4ys�e-�Cf��0A����OC�*�&G�b���X��F�v��`�Yt{�t%u��E�W�)���Hx��fF#�̕tJ�m�!bu$']n������姞��C��4�f1���<���E�;�\�Xq���Z�e���s�_9h-��<1��X�7[}�7y���H�K��~�],$\�� �de��T��Y��5���/Y�V�����mf6�܊��n���7iH�dΫ�q$`vmf��;/*b�V&i�����^kS����]J5wC�]F�^�E�ʾ�����U��5��F�ਤh���}y�a�z��K� �' D�k-���l�a�oAѫ��t���������(�29��v�V�_׀�����s��ێfU���8��)��CC��ܺ��8f�.*��=� �1�(�8����O=�Ye���'�	�bh��r%Iy}wv��rHQ���;�Hi�h�~���מ��ȉ0��˹��^�����B�aE�!('�'�h�,��5+-�<�֜�!!5eP�B]Ԉ�Vk(�P�vy��T��wq�Q<'c�m��r�,�N�]P���)�V�22MY���2���hw=��'�jGP�����:��*���3Aww5��ӝ�tOt���.z2�Yr��r���K���ºE����uݑ�J��H�/"���u��S�r�]���$3���qԓ�*�
��&SHN��s �֐�_oκ��	1+**�]\�"3�m�Ѐ�HJߵ���Ϡ�MST��2��s��j0��5OLTϟ/w���T�Fq�x��tvU[2F�ŧMS;Z�p��Jn��c�ޚ�J�*iF�D��pc*���Ҏ�M*e���4��h�STҍj��c��)��vsGwx�ڏI�m[����0�3#E5L��1�UJ��U�(�V�&�f}�ޚ�a���ST�����X4յ��́�wp-E��σ"��DMVX��"��b�MSJ���zih�TҍF�t�L߱�`T�3M*c�/��ξ��9�>�Uٮ�m�Syx�����lk�Yy��t%D)��v�/a@3�̮��Y�>
�]
g�m*j��STTJ��뷖�Z�I���P�MS(7�{YE5�hh���Q�N����a���S*����T�-ST���&���zh�4�4R�6u���WR�u�MF�j3>�k��ZiQQSK9���֟et�x�D�߰cJ+iS�SJ��(�g|�����T�t���T7�{X�����A`���:��v6��Т��h�����z�tˎ�t�Q�44S9�z�ֆj�Q������X4յ��5M�j�50k����qOX��g醩��Zt�4�������Z�)���N�L߱�a�3M*ecYl�Y*�N��4��Q�{לf��k��-5J�T�TJ��{w���MS�*j�I��S9����k,��MSJ5����0�0�5����<���(ѝΜ��[�g���-�H�U=�l)�uV�:��P�Q6��E)bEo=+5�1ň�V�9cZ䩃+n��t@/1$�ؐ�F�ҍFT�s^�4i�j�(�q�C��-�#Zb��g�_��4��J���T4M���"��>k���+<���e����s��KL��L�M*j�C��u�SYiF��5N��{��5L��MS^����a�����z)˓��e{�t�A�u��;�N$�����LDj�_[����]�T��yj�ᢙ�ww���MST�e�l-�j��_u�M[ZaCT)��4Ov��SJ5���7�������Q�����騩�**iSQ���XE5��f�Z��eTv���gM,�N�+Z���2�MF�k3-��~��q.38��/�Zj�!���P�MS)o����kL�E5M(�h�����j0��5L%ky��5§�#�����0���8���
�u�MF�j3=�k�mi�U4��=��5M(�iG�SJ��jwG�ΚYfӦ�5Q�*�=�"���J��(�h�����j3&3��L�X�(�i��g���+������<km(�aƩ�fq~�&��0��j�Q��Eo��L5LYt�1Rt�4�=�r���;b�f4�Q�FS3�{xE=3Mu����FkΝYiʻ�4���+��`�
iF�J5�Q*f��^ZYj:�;��1��7��[iF�8��wYE5�i4ST�0���f�|�-S�ST������fϽg���b�9��&n�f�M��wb-,:#�V��l���Ltj[՛�����8�/E�D�5ǭs,��1��j�}w��Y������I+|��<�|��� �N���^�^��s�+��n��ۮ�F���)��Lݸ�	�gq���V ��V�/���v�Dq��{<�b��n'��(=���䱭D�U��م���|��2�)�������k�T�K�[��<\l�SG#;d��6k����n*9A�7E�msڄ��	R�ծ�/�u���k��Y<�kÐ���7%�g`m���8{4����tr�%��9Uc����U�=�}	M��YR���e���gu~�C��Ң���4o��0�4��)�N�M*e��cM-3I�J�ٟo�U�s��K-]C��y�SZZ�SQ�1ST��|�-S2�MS(�<7�U*�J�fQ���h�g~��4�5L)�`��L��Q�3�y�[ZiF�E&ST�K޾`�TҍF�j4�T=�r���Q�4SJ�o�-��ɍ�xE=�L
e�F�ꪎՑ��饖htѭWl�Tҍd*%MUD����yzb�T�b����)�g5��s��1�o���ZQ��ST��o�e�a��5L�,jڶ�3���M,�5�o��Ӳ��Ħb�"=�0}g�� ���>���(�ib�SG�[���T�iF�J2��cM-3N�T�4������յ��W�z�sx��[j<�T�:��̵L�E5L�N�d���9c�#Yf�)�޽zie�kI�5L(j��w��`�V֘V���yx�*��Ն��L�������LYt�1S���AP�{��#F���Q��o����z��37�k�ﻍ����mPX�$u{u�i�ѻ;��u�S�k�K�(HJ�Uc�.��7��*�NUߩ�֣F�Y�SJ5�STTJ�������MSJ5I���o��a�ZQ�Օ̙�;�5Mpg�}�-S�MSJ5���yh�4�4R1�3����Rْ5�-:j��_��Ӷ�ҍF��"����J��!�Y�o/�>�o�_1S�d��eEΆ��g��R���	ö�U��sVT��|�vp�-sVrS�ɛ־�$��@�HZ;�͘�Em*t�iS��iS(��|ƚZf���2�4���o��Z4�ZQ�ҍG����u��6��εM(�fe������R�لe�gF�f}�ޚ��MST)�aMST�{��Mi�0��5M!L�ν瞺���<�xq��1�޽`g0C�H�0�}�F^Z�j�{�:v���d3#s�ٖ4��<s~�|ؒ�c�y�cB=���`i�lA̾l�w�d��GiSQ��1�fŔ̰'o{\�vUԹ%�d��3�jս��� H��ٌ��5���؆��� e��`F��e����D���,�FF�ѿo��e�{�U�d�wc�\�SyyYŕ�D;�Lg����wiïSb�~w���5�t�������k����F�j4w~͙�JQ�F;�sX��\�co���w�#��s`a�y ��s��e堌���څYiʻ�f���j̱���]�/ک�{K,�1�21e&�C�����~cӏyĚ�F{~�ie��6����>��^���;�ݠ�xų���rYRْ4h�}���!�@5�r�1�o)�iSGդ)���w�	��JIXr�ŗ���hэx
�њ�G[D�d�u=���ή:�D�Kw���I�ʻ�~)�ؕÚ���W7�|H@�I m!g�0X��0#G=^�Me�F(�>o�,��5wOS��:�V�#-h�Ϲ��dx��y۽�0ņ�����k�4��ٖ+L���ن!���#��۝ �7!��Jn�G��0ׯ^�)堌��m�x�j��� �2����̳#1�(�o]�,Ya��߹�cz��LCh�oW��і��ڦ*�w�e���ҍF�j1�f���,�-����j��W0�̡%[�tcn��9�0������:�Wx���K�A��=�]�wN��%�x��3�ְv�IE'^��b�4ƴ�L��y�b7�bw��4V+��)�l<��|�,�FSDh�����j�X쬊4e4F{�Fb�#K�c�ܾ�}���;��pm�iA�������Z�Ƃ'��{|�3�!�"?LMQof��q?UxA���qj"<TL�f��]��f��j(�6o|�,��h��4vcl����*vܙ��M#F(����e���&�J5�s�,���0��e�eKf��hq���w��s]�Ѭ1$$X�l�`���G�s��0̰##5k��a�����I����VNo�F�awE��q$�������'R��e>�ZWcc��z���Vo��%_4fo�z��xև�H��Iia���F�}fX�ѕ�b��˺��ṾMh�ϳ�Cidj4s�sXY������b�^��.��T�L	�oX2�eƂ8�I2fr�&��XE<���ϻ��f=S����߯��v��ճz��r$[q�޳V��<��]��e�Qx�co��;�ܺ��0�X��fY�j!��(�oܳ)�, �#Dh����Qm#�{�{�U�aLV3x���K-F��(0��9�Y�c�UʗN�d�A�5=��2<1�ƺv��ʛ�>���h#�Aw��fS20#Q�w�^G� YD�C�;�}��E����LGj�[vV<���va�(0�Ch�ߵ�[K-F�u�v�{��=ά1�2鈊C��l�� ��W}�"�Zɜ`���U������i1s�ՙf��ӭ��6�6�Ҍ߷�2Ŗ�4A�4NW}��؆�6,�]�,�K��8w��y�u����m-5Q��ǵb�2���}>��[2F�#���0�h�U$�o~��G��q+>�쳈#�A���,���Cj3u����Ҍ#ak��h�Db��/2��B����y����S�kw}^y$�U���Q*u_jVW�{Cۺ��S��~v���ü��Yڒ��8�yC�
cu�B}��HBm!	��f�����#�;w-��=[=��ᝡ�ݽ���-��gNt��W=X`��y���6�������J��<�	Pk���y���@�����b�9n�l;��|����vz9���7HK��J�ә�k]Z���	����BU�l���ӯN�Z� �z�	��yQ.��E�k0�ʝA�HJ��cXf�]���uY�\�j:2kq����FtӮ`,V�]v:��~~��`���UIUl�2�6c�݇��X��6�OsXE��5�*e0!��0e�m�a�Zo������\�}��38���׽�"�Zɪ�m�v�v2][�fX��v̱�F�J5���8��J���vu1e�b��4MW����2���;�r̴�5���{�i�{�z��5��š��'���K�wV]U��h4�F���"،�6��Y�a�F�1���{7�{`a�C20#F���"��J0�Q�L;�r̴e4F���}�wm�Vݕ�F��F{=݃��5���t�CLCiX5==�`��Q520'y�`�A���6{�݀�\�<�ob`��V��"؆̙�T}����]�3L^��fX��ZQ�Ҍ׹�;y�9�|أE�F��s�E�� �1A��fX����6{�݋ ̰=v��|�g��c�T{��G]��n��B�ê1��к�ѫ<����ۣ6�h����H]���#A�;3�`2��@�D�oܳ ���頌��o e�`Fj���0Չ��{�E���aao��h�h��#$=�W*J�f�!��,1q�isOk{ǿ]����
ٕ��\���f�:M������EM�][��؞'7y��R�t�k$QC0�LjE��Z�P�6>��&�Bl km=�x<a�������`�A����|��V`�"=�w^���a��;�-����Vcm��ˡ���@�4Ŝ��e��ҍSJ3����1e�b�4F�{~�'ou���Ѣ1F�3��,�K �iF�J5�sv,�e��ݪ�K*�H��a�Q���:k�7f[�g6��") �;�0�7��1�����,�2&h�﵄[^���꽥��FֳfX�ќgl�[�m��쬢4dh��{�����G&��k/{��_�w�;�L���o���!��l�9��0C�F�N�XE������p��̒��NTn՘���-�&����]�{l�"q��yzwM_��y���ӕw�4��s�0�0#4�Q���ve1e�m�4MW����24F.gY�����l)���,��Y�Cg=�ز3-*t�}*u�]���#�91�`8�� �k�۝�=���3��gVa�lCb;�wx,�25�﵁[YQ�lVNs���=:^�h��=�G=�w*J�f�!��,8�,PF����e5�<	 " ӿl?��dL9C����Ϲ>��Uema�Mh�nMa�$L�(�ם]Z�"x��'����A+>��U8��`沧�3����$x� �}�h>1���w`a�y�#F��k���2-Vcm�y]�V��,�ݳ,��n�]����l:4�=�f̱e�b��4MW9���2���{~�iw��%�?f�{�YiP5Pj39�lYfX�;�S��w.ܫ�4�i8љ�o��"H!�=�r�d�#�5�9��= �Md��,�2�f���mdiF!���ܳ-M��/�s&ef�U��ڷ�Ͱ���n.u���n���C�ٹ��e�5�{�ݶ�Y^Di��u`a��#�97�`�XiF�8�L�]练-G�{3w���v�qHcXխ�kPC�Dq4Us��-�lɜc��%�N]�m��i�����2&bY/��ϳ=w��,�c8�0é�4F��پ������6w�Y��Z�(F�y��k�=|�����X�3-Z���.�V̑�m��0xb$[�,�H"8�F!�J����w��x� �8���5r��a�6�û�,��2k�9��w*UU�(�F�#1��«��k����u��Q����pe�1����h28�G�A!�k�W���9��I���c��4�?D��pk���]�
�}��^�g<�V�*��l��z&�C+D�����;�&�!�$ �!�"Dq0��y�[��F|������� �21g>�fFj(1�7��a[�3��.wθ.�dh�՜�(���F(0�Q�߹fZYMF��(�g}�ز̰�&����6��3UN�K�����*�b[���!,�ϋ9gb���?>����V�1��9��� �H��Y���lCd;�o e�Lɋ��7Ҷ�m�����k#J0�aw��,Ch�~�ucn�,�"4m�3���22�F�k3SZ��9=�a��Q�߹f��e�"){��3�!��w��y�a�k��-�4�9�i��%������i��ά�20#Q4�PiFk�݁�b�#G|�k/\P��-��<	�#Ȍ��B#Q��;�nŖe�5�,w��]���#�3=�`;[��cLGI67�Y�!���h#&����,��5C7W�a���\��i-��{~�h�Dh���!6�.�J��eb/��b�#�97�`�Xiv�O��g�k\[bm+7��X���G�!��vV`�	M4j{�Ǆ��"8LC���*�_<3���V�n>T`p��=9� z� w7:�b�ט�T6��%�v��̘֭�fl�\鉤V�+�2¬�G�e3O�6u>�r�9��!͛�w�CJ�7ڻ��D���V��-�x��M��Сjr��]Ժ9�K�Ows ������B��{���v�f������̼ʳ��Q��4z��2ڊM��Y���K-�ެ;[�u�0��;SŊv �]70�Ǜ����3tj=�������mh��SW��V���L��7�c��8�u=͵u�����'G�i���]4�=�˳���n(q�C~[k2�s�����q5��ڱi�0�
ƅpJ��.��ݙl����f`�)��peԖg]����������*�G@v�6m�����.�={K,q�w�������t�I�^ۘ��:�_f𷕚���X.�VF4Gcn=�wh������fwe���7ےwU��7�|
��ٓ�N&�42�G��w+�ή�FC��Ӆ��l�yeQw�+1K�wo!�m7�Dg��sf�X4(�ӥ,(�0(�ɶ��
ܓX̓�-��t6ݼZ�����W@0�ѷ�e.���N���]���{ճ�$XK�Tk9ǖ��7���+I���`9y؍���l��r]�-��j h c�P�/�#����\l�ʼ��t~
��m�~}����ns��u%�%E?N�﮸Vj�M����kRX�TNQi�H��"��=|���]%0H���at�9J��z멕���]�$��*��'*��IBQ9f��DAi�U�WJyN�\#e��JǄ���}y�����"�D��XPf�t�;�܍���ʪ=Ds �%�5CK�wtL�e!	$!�vA')J���'U��.UЎY�I��r�421R�)*4��+"�-J*���(�xQ��rE2�pY]l�<t�PR��j#T��M}[�W�J)o�E�D�r&��*D0Zp1Vjd�rv葙VC�:b�O�̐��J�hp��;���	�R�L�,�#&�](��-2��l�̄�
�[3K�2��<���pI:�:!ƣQƆ�l�r/g'J�/ww`       �ԭ:V�n��:7�Ok��R;�]X,��J�H�\�&t$o/%���z��Q��:�[I�g�
��;��Qb<{�������|r���v���^��a7n5�M���<��݃�qi	$�'�q�r��C��#>�oN�y�U��Sm��ݫ[��zĚ]��r����k)�]<=��<勞nΡ��/����a:�W`�܎���k|�ns�9�4m˞����@�՞�����&�gU����9ݵ�cn�-GKt]�Lq�s�`M�Q
u�����ͺ�m�Om��lF65�u��l�7b�S���!�]��v6z헨Ƿ8nk۸�='�ގ91u�n.��_=��t��iGC���s��[yuŕ�������΀#�v����s�Wm6��#��{�jR:�@/��5�^K�<p�;�y�mΒ�9��f�\FB���Ŭx��56�nx�<Z��C�I{,���K��n����M�o ��������hsɮ�G�9�@v.��>��Kֹ���:��{P��c��Ǌ�۷\c���=+/���N�[i��C�����O�q���-���;���H�%<����x�wr6@�$쫞�'�䗎1�ss�g�i�u.�;[l�����\����n�`�d����^HI���ėv��=]��0�ݰ��"�V��m�׭�:ݢ�ۇ��Ɓ��t��u���Q��=�V#ˮ���n!ä������֦�ǎ����4�[���t�r�\z�\7G����~u�>9�7g�M0�n��1�%�̐)ۢ�{�R����\��`�n��3��\�c�a��=�j�㴰i��B�M[�� ]�^��[���skfz�F�P���@4:+�JKy. �ݓ�?���[<�I��UUU�|o=�ѱ�d��^�M�}��i�n6���b��e,�[��gs'b�ޮ���}s�
���.c��:�������������\3j{l��r֌!��4S]s�s�+���G]�bn2ˆW5�G��M�z���;K�&����֎N�n�tc�8z�oFmm�n�ǉۃuK͐���1�3J�[�5ی<Lg�n��#�;[�t���x��掍�3�������w�m���nۄ���0Ϭb�}�2̌�6!����1�#Dh����Qm#q�u��]��j�b�7�v̱���҃Q��wb�2��Ƕ�rY.�]T��LCh��k�ሒ�}�����&��1�"84�l�����#A��L�w��-����o;�+���<׬�GZ#D+<����$��+H�Cgq�Xb�7=���XiF���e�z�}�~�o�Z�4q��!��vs9GW}�"�Z�g=�>�M�i���3C��Y�>��� �G#TҌ�cVe�4D�&���QlCb��1A�߹fZ^���^�4j���ˈ�ղ���`w��wEB�ul�'�7�a�fA�oܳ ����|�kh8�����8,CfFj�{��-��(�1F���Y����w�7���}������C�.wmg�!�p��愗cҝ��7�9q�v�}����*���m����}`a�m,�97�`�k(�b߹�-G�e����b9!^�l�p�#�W}�"�Z�=�co�zݷ	uo a��g�a�`F�4| �>��B��&��Ub���:�Q�-�����2 ��o;jbĩؔO���t�շV�|��ӏ�I��.�x�54��>	/�6	iy���ω�, � �"�_>k(�!��daLQ���Y��A�҃Q��i����/lo���${@ek�l)2�)��h48щ�o�ሄ�! �yf����Fw>3�����U�s�ʗ{�fFd`F�f��me4���0���2і��y6���ܑ�e��F��F{=݅�3^+�1����-�1��Sz�����C`@׽�h28�G�!�sV����-�6!������6fg>�7�M�I����M.�ڳ,EH�ҍF�f��ٖ,���1|�nw��%g����'�Z�Qmh�Q�b����2��ze4��҃Q��5`a��Û.nNC1�]�Lwr-��8u��9�/-�媥5��6�똬������t�:�x�Ch��y��xb! ���y�1�"8�F!�{�� �����}9�-^��EM�E�a�(�׹�0і��5�9��w.��ٔi�CDf=�Xe0��N��OL��rc���҃Q����bA��"
C�����m��g�[�6xΰ�zh#"�b6�'��#wV��,�ݳ,Ck#J5A��ve�, ��Ѿ�(J����Mf��MN���A���f�VwX�yp3X��w�C���c��N�G7V]�i����(�7�I|h m$�o=�-��Db���>r�4���(5Q�ϟ9��ǶS�U�w)�.�i��8щ�oӎ�{���:�{�b= � �sf3G�A�wv�̌�f���ms5�S��|��a�-0�`^��0�6��+^�rܑ�e��F��Fs>݆S�D�1���������ɇ\��L�	��x2�6�#�Cf���Y� ��W}�"�F�3�כ�����o��������j:�S{B��*�v�5ҢW��RnUc�.���S|��:N��u�b糫2̰#Q��J3^���Ŗ�0�M�5]���h�������;w�.T�k��/8��idj4�Q���y�Y�Ŝ~�v�c�fH�6�Og�M����}�ch�uO >��Q�h#�d߽��e�j�{��-���1F��+Ǳ�{�^�α��m��$��UUl�2�����a�(�4��h�ߵ�[K-F�7�O<��u~�o{醃Íq���7`g0C�Dq����o#A5X����vBV��Ŝ��e��o���sW�)�&�j(�ƹfX��N!�������8�$�dG��g�˽�<��f�M�1y�)�����u�e��Kr��ܵ��弾�VʟNH�NB�c��;/4V)Ү��$`	��Bk�/���6o7b�̰'���UYWpue�M1��}�ǆ"H"���kZ{v��K�>d1�� e�lCk,�{��-�l2�F߹fZ2�;|�w��ϩ�>篟��[ֿ3䍜w!��6�f�q'�Y�3�;	��rc��t�\e�[��.�˒7E�_���c����F���氋idj0"d`w~�h28�f�������9�#��"�� ]�N�܊.�˂yI���S+���J�ڷ���ܙ�N���"�H's�
+��n�zNTB��L6����&A� ׁ���I���A�
�(F��1��F,�@���s$�;AJ՛�*m碉5����� 0w��$���w<	ܨ���xk�"yf8`W� �Th��	.�U�ӝ��[��xI�]�@�7��w<��n���p������Ά!qY�ݳ��D<<�̀��C�����'\�''5�3�*����&�Y$��F���kv@� ��$��	*+;�����ݔ�%�t�v����u�v���96x㋳����ì%^y0�C����Z�v��y->�+g'��ٸ'��Q�9{�b���Lv8�8�4u�]λ��+/�t��.Q���h@`��[68Rے8��m��p��ɖ}�8�ê�v���v�Y,S�H�K4Mm�V����sn��p����լ=2p�3FwTu��wD��۶3��Y��J���+�ݹ�gS�*b3~=�~����M�o�ɧ�D��܊��X�zX�0o~�b�wS	���(�ҥH:}����d�#F� &{S�(
��t(ns+�h����~��ґ�6��6��� �<�$���o��T�%eM7�FvD��H�<�Fvt�3L�2Az���u�rZ]s�+��ʯiy-뉊[k�|ж(�jC+��{AJ՛�*@���@��O<��d�ԓ�G����k��w[8%�i�
�t��Ҟ@�\\�f�qz�p[Q���TnǱ���U%wK=���� �Ay������: �H��q@�۩�����ǓA�kVą��9���Ƞat�F��Y�x+���4/V��V]��N��(�գ{,�"Ft��	�W���o�;�V��}6 Bﯜ�6���D�"�߮+ě���'k{S��>��O�$L	$�;]�(�uפ��Yً�G�� ��}М|˪���7��&�[����A(�1�@%�m*�$��Δs��r/�Mf�$�Y��.z)եeE!A��}����L�^\�b��O��=�TA��H���l+�eq��ew�����R�iR��)��0b�����~lFs/M[�K��W%��������D�+�k�ר�s�����H��T��D֐���(sWR��8WT��o���P�g)l�\m�}���n:Тy�^"�$��f���͡��AN$DI
$LՃ:��^K� ��r|�x����r��������M��:����Kl`�y�jiU���ot}C<��BUw�Ff�� f7��j�7����}6��o��{�|�X>k��;_j�@�T���:o��,� ��I#w�z�{�����	�6�m�"t�D��i)+�q���hOMt���oYPM�[T	'��h���T�<�%}oϟv���_8���7e.�Zn�ٛ������M�N�%*��*Owº�Մ��<����sD�I��TD;��ka�@nGr�|	��\@%eL��)��m�b5��JA#˪��r(��u@�C뙊\���L�<vO����k���N&�آO����$��'�q��A �c���S��DD����̰싃ݣl��QX�I$��B��]J�����@�awp.�}O�:|NX�i���iP������8����l\7����������}���~|hI��K_�����0�_�un� ǜ�t�Cp�7e���������O<ܡ��}b�	i�߆�}=��A�"��8V����x�H�5��X!��Yx�4����Q%(�D��٩�9�j�#9:A�=7����ϲ/6(| ��t�>��Y�!L���v�j��1�w=��^$�m�${J�H$�#��X^.�����h)Z�v�IA�F�3�Yb���-�[WX� ��r(���U�E�D��
'�j�
׹=���L��b���y��Ѷ�I��S�_YW*q ����*ΕbЫ�If�� 7۩�t��w�8H�� ��}j�&����z��,{*$��:��;����9�������r�NY Sޤ36�4�]���'/�T�2���E�����F�d��Ɛ�"�{�����ݔ�%w"�g���n��;��]i����W0�3혧l)���<�K����d���7���|v^j��5ٸ�5أ�)���l(�sp�=l�;bKݹ�ܝ�v�����vާ����ќC����z3�`���;G]�)���c{Z�o]�l��.�c��D�pb׉�k�^\�-o.qL���l]��w%�no4��;>����{��nM�:\]�߿>��2�^��"˝���x��@�{Ψ��n��>���.��	!ڢ@�j�)G�&f�MH`��N#T�,�{�$��6ТE�:�Di���N��v�p�
T�0O���
9��P��ӏ�N1Q5TI#z:РO��ר����L̨�"��V̌�م���C��B'���u^'�w7w8kD�>W�V��I}�|P�&jkv����Tǘ�Xqx��O/[�$���T��
M�o JBW���^�����[ ���o�L�Ŕc�����w���`đ"f�5w�I;��x���ꁅ����m�j�	$fk�&��t0�*A�Cϱ�*OVٖ���5������{9V86J_XH:yq��ʊף	�:�l�Üŵ��Q�U�۔�-�R�\짮cr'f',��W�<?�xM�$o�������n����7����n����9GC��D/��No�t�����K�H��{;;r�%��@�n��|w��S�PR�I��|h�\�P|ډ�O�A콚>����c�4C��6{�VL�vS3*bH�;:�\P.]y΋�0���ϝP ��ޛ"]���w�{��c�m �*ҡWf��'m������ݻ��v��Bۮ���XY�����~~��8���O��C�کН��D�/2l���;�� \ޑ	�"$��6#�,�ӗ1�J�z
�$g9��g}8E\P��2���\�u5�%�2$I�w�(
 ��2���G���L	1sڈ�f"�`,9���0&�2��8L�¶�8wb��(Ԭ�r�H��o�4� �\U��Vƈ��39�}��\%���"M�Yv��ȕ����Tvag�	��A(�x�n���^����<�V�yO��^k�66�`ݹJ��nt�w�x����d�!܉�ג�����4���t�m�on�VQf����5��-�)7MKt➲!z�r�ܮ	�Euu<�ڵ��H���q���nJ'xd�'d��َr����z�.L��M�c����^*ft���T��"��!�ñYSbؘb+T�X�N���n���Psw.T�\ų(ˢ+%�r����B+���kE�"61h�r�SX�otī(��x��ɷV��$c&S��.iAof���kV�0#4�H�$�^ok���ow-�d\eM��`�u�f��SLb{l1FSo��f��-�Pe��Aƣ$ʌ΃�q�<=^��F[|�>��荍��)�yc����/I�N�.-]��w�\��B�lE��2p�1���؈�zl���}7�y�U�(Ne�;�j�����u����r��b��vf�ga�L�nڰ������m�b�0�-|�n��tᴞ�����o[�.�n.I;zqӚF��w��wT^%�D�b̈́�3��
EI��n�m�=w�{��ڍ�gB��y����" /�^=w�K3'��ڂL����p�d�$ß���~�=����(9�$��AeB�}+��_�9܋9�I		�I�(���,ʩ$�Ժ�eH��TT��I
�e��Ϟ�I��9�P�J���ҭ4�U��P��+,��V���b(EVEF�ir᪴$���L� ���,ü�^�uR�Ь�4Y��dIfQ���QQTj*�1J٘i�����(j�(A0čK)2L�CS�5T6p�I"�4T�\�P�d��Fʈ�"�(�2Y�P-5LC��CĂ�A��Pf��%TXh��̫Z��"�*�g�S����DXfT�52�J�SS\Ľ+���%��
S�Ftt��.vC����%5���oѤ�@����_D�>w��<�>���|��uh��I��Y��%Y��랙��V{��F�:�bwLwyH=��[3�HR�I��|h�hy�h�����v��$�ʯ�s�0�:yÚ>.�`Y���-rw���#�GB#��y�X�^gsM)��sƹ��u%	o�t��ʘ�3�j_H���(I$vs�0���Q#�T��Nn�"��H��%*J������՝��/"st
$��4	�;��Q���}��k�3�Quc�-�"$��7fw#kr([V����4kݩ�$�}8E�r"|�D�FD�#�"����9�t���q���νGs���X�b������cGo��&6�V��yd�y[�8�XU�iU��p�3a�8l�*==����X��uE:��7[*Gqժ���C��&���犃��㲭�UWw���3���Ti�I�d�Nx���@ٮh�@;��_�t:���k��+BQ"eN(=��θ^m��g )P@��i@+���֛���j����k�h" �k�D���D��Vzw2J�4kē��Q729(�I�F�JW��(t9�Y��q����8���>$�vUAS}L,�8s�C\"&JT��U�T ��*�$S1V��X|�`	ݩ� �c�*9]d�V�]�J@���ڵ��A�y0(�	m�P�9�8C��w��.�@�͍����5tE�B�0w�:`W�׌�f�2巨Q'�v�A �����ӆ�e����H�d�{7jr7�/�"!���W]����7� (E�0�k��eXa���������}Y/{�L��wZ�I���������ݔ�GC=�v˰�
m�����)L��q�q��do5/^�I��z��U�e���|6��6���sy b�{sx9댋�}�mh�US�mq�M�q�l��K�lX�mi�r�1zv:�iB(^��I��gg���v�8X��6�c�mX�zܜ���t�.�|�x��u�Ɗ��r�;\iKn����|7��8�XXթ4s�N��͗��GY��N���r]��ɱ.�r�������S	�DL��꺢@$���x�t�4���t���U��X�ˮ��"A��ck����Y�U/�l- H�ܯP����W�/:�+��V����J�Hق.���TI9���c&��"�k���r�@�E�v!B.)p�0BR�͊�ں�S�������;#qP$�:�܁�"�t�x��ڢ#j��z�b$L��Wo�A���#�[pz���P$�.�D�F�:�F��7{����*1``D�����M�]727���N�mS��<N�LIS���!
Q�'�wo*� ��B$ns��IЖOE͙���p�
�����/��Rw���
=O�m��,���X*�(�[Pa}34�ε�lovܬ������5�\v��"�LƄR��T�h�1sI������� 7~�'���Q$��Q�@o��oh���"R*'ƏRֽy�,O%kn �
��^$�.�@�O��&�x�̉Rfvjs�Î��j�ߟ�5�B���u@�H=��+!�5�!d_EڠH�K�>L
T���گ��6�8��Q���������Ί$7�ר�_UA���'��'W����%g�vUл�wf��;`-p�f�yj�[q��ybw��5�?�\o��K���Z ��	$���I$�vP̵6�����5��U�GksCąTC��""`�Gl��jõ=�ݮ��*�í@$}�h�Oge
�F��e��8�E�`aT���JM��S=��
V뻭p((K��00ھ��3�sJ;v��������H�)�6=l�azi��Ǟ��gb�±mJ��}�*��;g�G�I?��Q���+�Tv��DH�����8�==����d�r6��>$�&�A���^d�}��v���ʄ9*F��EM�5�lC�-ӡ���7C� �b�@Ua�e�N,�f3���o��(V���Wc�$���K�VO7I����v�v|�q��T�7JL?
�P%}e[��P=��� �{�lh��7$��T�+�`C�؝c�GV�Ut�ڤ�{1���ѓ�՚�g3�  ��ء��˦
&&u9Z=��1唍Yj�T�玨�4�eH �r�����m�
Č>�[�08�J���%'�G ��t/62�.��Q$�\�{3�G�vj�U9+����NN9���lSi���q�����=����T�kw7�;|C�%�ZO:�'���U���_��+����7j���4������g���'��1��]�z9-�`
��˧@{3͋[7�6��=AT-P�]�J=s;uj�.Mw�~|�������O��<�r_Ͽ��!�dJ0���O:�<�$K�:F�.�+�;���E|->ȯZIR����A��7T ��hk�w�X ���M�uP#GOg87=;�h�%`!v�)��h
��L�J�Ҹ���&�u�H^�UB�E�hB ��1"M�Ӹ!`{u=Ѽ	8f����Ϊ>�m�d^�/�<t���}tI� ��i)=��>�On������v�0+6�ۙ́@V��r~�R5o����osۄ�w
z��{����u0/ڝ�e\�[��T35-Z�!��aT���\6艒���Q�Z`=ҝ<v�˧�=�?�� �
MȒI$�Z�9뱣�s��<ln�m�On�k^��{5U�I��'u/7cB�=�5�,[k�W�rrʛrt��Vd�F뛍���&:�g��5'[gl�-�<�/0������=�{p'��5q%ȣ������n�G�i��t7rOld����x�%�yz�K�����f7S���^ܹuƜ�n��8�rS-���y�;�yٴ�bay��3fnǮ:Ǜȝ���v&��7~��1
D�TO��t��H���4��m����y��}�2��$o���d���(D�D^]N��S���َ�$�mI�&�6h|	���AF��]�w�5n�	�K�7��d�M=��{5Т ����cLݸ�A-��|H�{]<p���j�AZ��{3��,�&p�/�W�d�	��TO����r�����U�hQٌ
(�
$I�����Aӝ�鞔���1QN�ĀGḵ`�w�(�t�ƛ˝�+U�K9B��K�e��.@�.vs<��<�����X���GJ���3{�S���ܑGvE�o.�H�[Y|�I�';�qA:R%"�|E�� ��vN�r���*��}{+�[
�V��c/#�� -��#~%f>�c��)����'ץf�H���q_�N�I$}ݕ@H���$��{Qۤ�u�I�"a".�5:�P8y�	>$�sQ��ձ
f�$7�(���"��{�h>��&hU>�����uX�v����A5�"�I=�ԦrdTIPp��NM"0q��d�H'��f4(W�5:�����0
��uP����s:�e���O;���Z���4A�j�mt�
�MۤʷO&*v�7e�٠��;o�ز�7j���� ѝ�胹�PK��C��s["����[H��j��wiOrkh
�9��wG���q@���A��Y�1y+�*���1��Q>!��Ăo3��H$�
R(C����[u���HWh�ι�r����s�X��۾�),�K=uhOa�x���KW���>��/:�w�0�,埇��~�G�����Gٟ����Jq&���vu:��!O�L�����I'�mP$�yt�gA�b|�gы`M�kA����(�c`P��uLލ��1z���
n��P���� ���879GP%!�T'��ջ;v�.+d\�����۰������=}����EZ���S�,vcT���tw�#�|�o�mdP ��uQ;b��pPaL��D�7[t(�L�X�`Ξ�$>Ϊ �s�Ex�t��8�}:K��v�n�]����y5���:v����lOf(r�8󪍔t�DLz<�d�_+��J؇�4�4i�1@{�|I������X�$��*�nY{�!R��
Bd9��[ڎ�5-��OBy�ﯣQq���*�^�M.�2�ɎjL��_��&ݺ6'��D�B&
��5��
���"���r4+��$��r�	;�}f^`�2K��!�_�����[�U˓�.P�p���v۶�8��<�r[ڠm#h$�7o�G�+v�	)�� =���
��
��33����z�/6�>$����މ�eL̩�";2���sw&S�\t�u=!�	��C�~/���V?��]~��>�Lr��vU�JT����G�B�= h>[r1�=�� �k�@
�EO�0=~Wj������5ãd��7s�C�� �A��$����?�x�Ch+��W���%R$��h�<�8��gMx̩s��/0>�	۹	��0B���5��Jl�눓2�Іneh��Í�# �{��Y������N7'dL
�:A`6,����2M�m��:u1H�ŝ��\�rNK7FsZIeJH��K؃7|3��{Bı���I��u���h��ۥ��/�h�$6M�j����ھ�})wv����^ݍs��J7CrL)ݰv�շ�����m>��w�k�޼�A�o'9��#�V]ލ�M���(��۱�ۣs�_[���S��@�{@����=�M�;+GX:NN� �GX��S]�.�,eVz���P/���H�� D��nlQ����ص�T�}�%�'uZʝn�S�aX�C��/'hBBЀ����?i�d~�k��c��<ds:��\{�`�������)j���m40+Zx�g�p
�v.�Bj���J���i�ݥdb�h�1��%K��Y�d̫��d9�������m_l�s�lZ���cm�<w'*�ٟ�]Z{8{n3G�X��iQ����קC��pt�r�pF86����ﺂ���j�{��6"k8m�D{F�i�	gw!��s6�j��H�7hs�gj�a������n�yM�t����剗��ɻ�/q)Q�no>tV�=�˄�Ujx����L�E̫^�v��]��5;a�.�Qʃ_C�(��(�G��o%Z�q��5�W��C�����	���ӽx���*{c�>"�S$�ȫ%iDW>3�O�*<0��BΕI��z�������c�p�6���WAadY4ZQaR�YPY�#TR/��q乪H��W�%��h��A��*�J���wy��/�U�afME�ԋR�ŕbB�PH��JQ2���&��J��h�����6����+.fF"b�RJ3 4NUU'D���͓IT*�"���r��s:D�Ue�fʩ�΄R��wK�+P6K*�P8Z�������PEW'��R��ӡDTE��\�Qs�E�\ �9(�O�z�GZ�Pi\��Bʨ��Da!DDQFZ�J$�GQQ�.Q�
��IQ�<���        y�9�tCt�f�i|G�c��w1Z�un�o����.��>m�G|� ��ݯ%�q��X�]��&���W?ڀ����];��s&ϻm:��3�v�<]n�MwP○fی��<��cS���*�Âʎ�2m76�" ����v0b뮄�N�X�5�h����m�5pt��<|M�wÐ�ѷ�[=�p����e���,�n;7��ۑ^|wD�y�g�s�M�U���xݽ�8�\ڹ3�z]��mv�v��Ͳ�p�Y�9���&٥���3�2��X�n+�ѥi2�%��Y.mu܎�8͔7zT8w<��l�:w
�5�R��-S���hq�c�wbչv�t&�݇��W��s�lm�w�ݕ}]Z+����Ǔ�=A�����wI۶�v�6 -�͖q�:v�#7a퓎ܔ�n=������[KѤ�C'K�1�k�	3���`T��7�n�D����nY�d���s.zm�ӣ4e����շ)�'���,5��]��"'�n:���`�yݹ�-��Rǌ\m۳�NO ��nn;:�=�����׬�.�O6�r&��0qcs%�����6(Yq8�ώR�T9��캭�y˻!�.Θ�^�E��7g����v䮟6��ո'�E��Og��:m8\��vK�#�Ӄt=r�b�Ʊg%�������$�rp�I���'v��8�rg�N���wϝ�g����c����ϋ�����fō�Ov Z�M�su�ň7WW<z��#�E�6:x��j�m-mJ�� �����(�x�km���:��m��4n��!�%׌v�F�R��xnz#��ԋl��^�!{�p�7F��%��������4qT�:���nkS��_��� 
���fwN���W���Ge1n�Aγ��z�c[�j]�8'�SE�����{=\�뇝�m���x�׶�N�ltu��Nfp!�7�7�ѷ�G���	�����vJ͘ӗ�Z�a��m$�P��]��vv���;.��"#��r��;K�q:�q���NL�qm�슷���@�>(����q��5���c�'on�K�=��r�kQ9;u�M�6�;�t��_;��%�E�*�ů�x�;��g���&#�a��yo�3���;��]q�b`���&��Uj�*��p䷱���H'ۊ�H�Ϊ5��G���>��7�"�Wp�WAIZ����I ��4! H3�[�'�u���]�n��P+���*�%/�.yנ�D{�A��U �[Ϊ�$o6��P�xe���g[��^ U��I���T�nd9�Ө� �v@�HǝTA��\߹޹c&��l�"�X�,ZF���yě[��\��NH;\���h������߿�.�IL��:g���Ffl�$;�� �u(��38�Y�(��6���`���(?>t�u�����pK�l/�+Ҵ�ۻ�����u�U��;w>���:��nl�VM�gU�wp坚���z�\n;ћ_��9&�?H'�g�H�����߱.�VLw�C�
5�V*�#I�}B���TA><쓃�y������Mc�Wh�("mZ��Bǳ�e�)�҇/}:I7���=�Su����@���7{H�ER�Q��(�K9�Bc\������d�A{ν@�=�ڊ�2"K7:%�Gd��Y���f��۶]��ʜ.�en�5rWe�6�Y��l�!O�D���$/9����ȠB�f�YCe�W�� �TD@��J�d��p������󑐱ck���`@'[u���(��F]��`k��t�U��*�]Θ�(`�e:@Re{ >�s
�3��~�{Kz5%����9Ok]Ij�5 �Yڟ�=���� �9���k����"D�������Ē�ΨN/߲(k�<BM�I!I-�ٙ���W�_�(�s�� ��P$���8�
��3�|���ܫ#ÍYAjթ���?��(wf����w<? �t�
{.�=�l!��B��v����b��с2���2n�Ft5z�r��s)���h��h��]��Ԉ�/�;cl 8s��	�U�}J�DH�7�N e^o��bǑ@�U)��
�B���ՕD�
,�Z������> ���$�gM[���H�<�1XۧC�ʫWd�����jH"�6E h��{���+�=�k^G��:��<��0D�%���<nF����C��A �͚�>$�vlLDcS�Mȃp�ѧy�P�čo���W�&����X>K0��L���y{n�e���ёf-9�1r�r�������Վp�;>b�!��ۻ�V��c`�5�X���զ1Lz�'�:hN�u������"�x��G�R$ui]��m��OW-�cuu��|,qH�-�~}�������?wE��D{qȠH'y�P7u���[�`ߗ& ����Q�R"�TU�����/f���RË�D�Gvm
#y�
Q�fu�\��%e�r��_]�O�Mx�	�y5�A[Z���Q2�&�uQ ��n6#HǕYF�K�?w��z��{6	�ޚ>�ܟP9�sm�N�jL��D�Yɺyhu��I?HMl}C��JQ���275Y�T ����Q]�#��r�kν�4�׌Bn�6�$QrȄ���)Oq��e4�s��a��բ�z'�z~}#"z��P��ꪪ�ͮ=2`�������=�06y����>�fE��Xx݇[y�HX�d�������爳f:5{8�Df��v�u�Z�:�.$g�;N;+9q���Y�+7�;=4&��.�;mn�q�\���k��nǵ%�@��ŝ;�
[{) >�Ѯ=����݈뇮�mn�Wk=G>�nd�����γu�Whl��k)=�E������x���T=w�I��t�˵_X��m6>뺼fA�ݓ^4��\p��7�UD�A���&h�t�6�Z�U�c�(b�҆�{�*勒I>�ܪ�sk��I�o��Tz���U�g�h"���Ѻ
�=l 3���3;)7`�Iy�@P$���5�ER�"���_]�Sܚ �SwY׏��ʣ�AI<���u^��%��A�N�GҠ�dDS>>�/�^gH�p�<w-��c�ލ:�>��6>}t�}�7�~vnͧd���Q�дYt����tv��y��ҴD�`D�H������HS���B�$fWMI�fu�]f6i����Nh��o�Bc�`T<��@�WA�.��� 9��5���vD�c�胤���nnӈ#p���؉s-S0h�ؔ]T�&��q����s'f��;d���:����$��\���3�Q ̆�r�L���YG��t.�*��%�D_ez����Σ�'�v��o&�$y��N���Q�2�����B^�{����xEK�G���3q�Ggd��ˈ�B��A'�܊S�`10Q�iI�8� *g��@m��N����&$=ΡD���j"���nf'֤D�/!�Ը٠��[-�$��l��h�9ݧ�vk�2_0O(�
!L��k�����@�g�0���2jXz!<�`PW���ҧ�a���?H���F�}�Wu���"s���O?��@��r���g	�N���`3>TV��|{^H�xe���[���-��O��A�ο0��v�z�S�7�� ��_N�K��^O��>G`��M�Mk�o=�����$���P$���5�V��"�S3v��y,v�W�I;�	 �H��+��^�Mϻ8�N@S�6Mj���A�|�o�n������>0S���N�m
�q�P$��E�N���:��ejŋ(�,�AU�
7չ.!�h��vrYyMx�R���$�)9�.��Z �6�;�x^nUJ�@���h�*����q��>7��Q�(��TS>>ޗ,�Ȼ	���ιd��q�$��Q>$��G8�OV����n9�$tX�L��T!vj�j��/��B� �l���ӽ/�@;���	%�dѳ�(��Bg����٬��5�2Vs���I/^M	{ՙqنs�̡�����Y�m�_p��"V��Jgb{��� �q�IQ3F���=��<Xئ����Kw�BWa`�����_������?�޲݅VU��ُ�l�����mī��V�U�&��ﺁn���ўl��wc��Ar�Ue��Mz�>�@�Q���ڧv*�( R"���"�D+_z�zD�۝�������@=4w�
eV�*c�t ��؝P4�]_h�,�RUj�t����^��q��� 
����T��LJVh	���D�~ɯ�[��JLDDώ�����N^t�#R)�7��I�yʱ��>#�nh����5�r�*����/>�+�3;)	�8P���$�z�I �7Kg'�y���ѳ��G���%�k_� ��K����g�u53T	<릀'Ļ�U��suQ����nW�{R�%���Q����hCr��%k���{�3�/�xg��̑���vܛݺNG�U�*P���S����T���KgD�ۼ�����!�_��ݸs���c��^l�N��,]��.�۶ŷg��8.L��˙'�8+�H���=�u���5���J�N��᫴���r�Tݦ�j�Ё�v����V�3U>Y�@�'>���aMvM�x��r�f�(p����<m6�z=/��5�׶B�h9ŭ�n���4��a�c^�l�)tn���E���n9z��>,����h����z�N��r�����{��6H�n��ː�Y�Kn��QB�Q#UX>��A�|ǟED��=\����#;����4	� �7>ۀ��-�Jy�f��4��� �$ٴ�����=�� uަof��KZ�ُnlv���$�70P$�-IQ3���Q[�uC�$��� g<�1/K��׏����ī̯N��FlȘeB�������Qn�20�ﺅߐ�"�%�\ѭS7|�����������.w9:W5�����	���Z;H&�Uwj�AZ�κ��(#I||���I���sF�KG�4ck���V�z�(ٺީ�:.��T�����L`D�3�&��0&���T�[�X��{z^�5�A�3�{@TB<�ķUx�f�C�{9�|�W���3�~��������ȣ$]��U_&k/')��7�R���}>����X�(yżn��6k�`�q �{h
�>w4"��uʑD�f���>q�^u h;�J6���$�H�nk���gM]&�B�[t	�7B�� ��i��"$�Dt�D���4zN�ˆ7)�&�.��|빯H�Ϊ�u�ū���t��?qu�s���mlGB	��*֢��^y����Nd!/O�3 ��J#��4��I#9�Q$�}�T	�a���یG[�@��s]� �,�@�٤�2��t*ՓFnv����s��M����:�t�����9�۴�<�<.��T���ʡW������4I 齈�(d	銅�\n,9{o*�nF�)�dl��d�P��+Xg��:��NN��e'Ô\��yz�W9����G*e,���9�o0����u��2PU�� 1��X��C|vd+�*�`�Ө�l�ъK�61v��P�r��a�1�Qh^m��ᜮ�k:�}���=o��[��iW����i��BM�ބ�4�3�g7���Ǚ.UK=ݣ2!!�'Z�w1:dsݤ:'j&t>�=km^��o�]Zfc�Y��\o��z���)$�H��@p��2Z��W��hN���!הXշ�w�|-��Z��ݜ+
< g=�y͝;���;�����=�FK3��Z�'J��_ћ�2ȇ�U�N�߻��:Na����ɏ\��T/U��v{��}��>O�� ]p��Y[�Wy֡�n�n���P7��<���!r`(OC%��V�&F����� ^�A�`#
W	�X'wUءP*!!�7oj�g�'[�h��R�X��=il��v��2��C-�z�Y͖�Lƶ.X��X��aرM��v�M��lG$��)����%5�ν55FΥn�dJ�����qő�*}Y��'wy;�X�U���N�R��=�.i���hܹH|�S��78�n�`�����D�Y��B�J���%ή�:#��9����5(2b��&4�C:E H �A�JT�5)0���T�\��14��2N�5����_=��֊�B(EEDX��B�4
���at�9!2�J�"�G�y�PAGe�EYbY���7AUg��
9Q9�����߇߲G{�uW�8^�*�,JCAP�*L��"ԱR
T|�v����Ds�W�(y.�瓕��tL��̬�D�ݔ^o�'"PN��ʫ2�t������R�b�q���r�e^(d��35���DUEw%D�L�۝�нܜ�N�
��E���"V�"A���rr��}���P��t��EFdh�Fo�p���i�Uh�(��ʹ@S<ZT"
rr�˕L�H����jQW9�tȫ�ʸTU9�*G!ȹt�[.&K���S�_�����$��A#�g�O��3$@������ۡ^�b��΅|H�͠;��{K���v�7�,*g��*RFͥ's�� '���|]Р��$ݎ�A�(R�r�u��s�P��^{EVx���ω7md��3�I�sźv{M�r��bAZ�� �F���=���
 L�L{�H�Y�=r�s��	�ͪ��h/rJ��D���T�?��"5傔���	%�:�H$�<�
�*��AZ^���WM8��p��	�%g	 ����������5q����BfrtP��o�:.��T�I'Dy͝�^VV�G7�(�1w\Y������md��S��N'�{T��]q�n1����s�;�AT�s��o��_$��]�����v��c�Q�D��$+_1��F�C�GJ2dW=�K�y����l
᝸���=�l5�w5����{��I�E<��]y��4�^pD�T�nG���-oA���Wh�C'm�ʕ+�n�.�o�7_@��ʠG����S׺r��(3b�r�Ē~ǔ(�P	H��
!D�h�yԓ;Q
�LCQ0�t���ɢ|O�wdP'Ǒ�κp26�P�21F�DJ1���Q�H�k����]�2M�gN�A�y"���\D����3�B%�=A:��O������G%Ϝ�'�9ɪ�ßn���Z�jo�Q̼�Zb!B�)LL磪�2��=pb귕C'ӹT���O� �g��J�0�^�mb�U�\�F��`��H�rÞ�E��P~�}�
QU��b�mdj�K��᨜?��/�$�I#��$���vv�iݱ��N�C�����a����(�w Ss�`y��t����<���e\�]VJ�ӣ.�jx����ϯWm����cOT��\j�ݍӞ�6疫�Ɂ��v�re�f��XT\�p��p]�p�7�m���$wF퇭��zzWsۻ'���W��5n����q���N3�[���$���ج6�F����ɺ!;ϛx\�ul.x	��1��/���?����ti�U~�}��TA ��,T,�#�ʥ�?�P�n&5���J��Ks 謯_�Z�«sr� ���@�w3��'���q�WT;\ĂR-�
D�6��@���I�T��>��I;&�����#�9@ȉF#�f������[�m� ����A�Q�gb���jT v�ɁU��.��^��XK����n� {��������P-�b���`P���dY��oyq���,�����W��;u�]7���E��e{�A�����Lr��
D�13�D��
e�r�\���kˣRĠ����ny�6W+�B�Z@�k���Hءsk�w��Yzc��q�]w�\"9��1�&���x�ym�V�
�J���+Ϲ*�Y{�$�V������]q���mU�d��_?�Gu�
|�ͪ ���$Q�x�v:�к��x5�`j�J��I�(��@L�?��`��b�H�\2;3f�'��]���I"p@ػWXk���f!Z�5�]^���P>;ݝ~f��%.�49@'kj��5^7� �.���zJ4M�K� !��0詪�v�����Z���V�G����s�'F�k�l�V�D��ۇ�霗����qc���.�z߿_��&���ί/�����s�`�Z�ȠTr�q��1e��d��>=���d:�1�DR%)��v�) 	W;�ٗȔ�}��3wzT�/�o�(8��/o_�����^!WV�%Z���N8 ���Lu�Md.a�}�2l�I�u�[ءG���սi9�ff�{@�T��i��#�Y�^�I���sV\��!�`P��LO��_��O���W�j��(�]ӸdH�DD�`��/%L����{=�| ��-Ь��7ļso�f�O���,��"��Ґ���h�y�|r�We��"^פ�8�˧@}��l`�*���H��ك^n�$��[�t�?>�ϓ.�7Z��;\�""m���� LJ&#����d�i�W�@#��TU��잪`X$�����W!��0f|�K�"������<���w	'/z�ğp��/F��q�Ff1����DR%37f�^Ex�z��` �b�����}@P_��'y:u�������|ǯ��3���펂���/(I$�Ψ�����L�G�o*���I�Q*hK"f*��G6������3�������pɖ�w�X����ujorTW����z���x�z��Ev�G/��	��P9u���D��M�JfR�7�	ۿ�IMn���@*���>/��$�w_mR�3r�/���'�TH�oWYۮq�/Z#Z��1���btq��LĈUl"�c�!1 ��/��|I�Κ�$�_>��>=���+ăw�h�ty�`�2I��2��X�p����f!פ�.��A�m��=&{8u���Qр��&�B$83DϢĺ�I�����O����l��y�/�i�����u������B�R����Q��9�$�٢I'�b��y�< �_{��_tn��+�ޡJ�B�HT
��ŜH��Kq�ʹ9�}�=B���v-�	+;&�=[����gj��9ua�-1���K#ܩ�M�]��T�R��N��݈�7���e��MnKЧ�O�Si�>}o��v�� :k�u���.�{c�ƹ�nSe��`s<]xnʻ��f�=[ Eޱ�u�UA$�l�v��f�n��*r��ݲ�@�t�Mqkq�:*�\r��y�WW*v�/����6�CM� 5����Ųt���y]��&�Ymgg����������n�k�n�n���G�/V�uV�q%D��@yâSf�Whu�ݧe8�n`r������V+��~�u˰����YTI'���<�����#u�^��>$��b�@H+��Q���h��u� �jmUX��;��F�^q����y� ]	��vY�=aGBL�b=C��hiMAƤu�1��I'��]��K�ɢ}}!��"f}�u�5~s	�$��@P��& 3����'�h���s��&�����J:b =;S�	��a#9Q.{e@>���I u�U���m�7�<��Bfdlv��<��v��;�T�s�L��7��AO��~~1�D��0�d���w��^W�ۏ����S�N���H9�E����fҒ��꩗w�VTK����yT�qV�*����ǹn���4\wؠ�S�%�fƑF���E��DDM����!oҦwk��sɠI>韛� *1]/�߲���#�����U�1 ���(���t�!�U�z�ǭ��$kɢ^uQ"㕃2H��W'���i)�=�Sqj�|{`Y�%�����b��q���d��@�Ԡ�!��"f}�g<H$�ܭ��F��9����&p��ڠI>9�U��2%��������ν�<lkM�^,�Ŗ3�Xm�^���J�����<����E��VI)\�
S�0��?��s_e� 6{�D����ta>&ũd�`DH+]݋�"�*�z+���8�u�B��}�`���ι��Q=	E�q(�����T ��b�87�oZ^��n���
���)�k�k��*of�/7z$�J�ww�+���z�⼹W&���c1�X{��ѡ^��n�Z죍���#i�Q$g?�@.�˫�VHWiPc��{�{���N` {�&�A'��`�Z�h���Y>��`��	L�Tz��_m�$ao"S�ȶL�uQ ��/��9k��O)��ho��	vk69r�G����l�m��<l�m;8ӈ���1/w�B$p��&'�ޜ��3�oE�yd=�u��L��� ��ۖ�sÑ�!#hJA��@Wo�x���b:�]�d��ݻ�dqבD�ʦ.��L��ID�O���YI
tt�P�<�$�z����N�H/7r��9v�խVGZ�j�ٴ�yv;��a��G >����_�m�H���f�z�Yd!�TQ
vLU����넆���T�5͒}ܚ�r��JVե+W�i���D�[W@��r�zxR�����P7'J��H+��̩Fb&A~��	7Y��1�V����	��wd�F�yO�Y�F�_-��jЂF`��(�B1R'ҐJ,r�(�֩�Nvv��>��D+*Ū4�q��R�V���P�;�|p��(�ugU�3+���~7��B���"�o�@�Hb&��*���$��0_Y��f!��$��"�'k:��&LdVȼ�T�9��u�tϠDHI]����̺c˵S���3:�Y��_u��;�l�H��	m��"̐�z�A��N�yY�6{�^�B��
ܧTI�256	>K' LCD�H�`6�ϼ�0(L�d�}��3�RؠI"�:�|H=����U�Q��Ӹ���VS"M	~9�y�&gs��7�"Q��J��dj�v����H`��G�nb�y��5bM�)p�'�6�S�Ȳ��&��4�=�oi�4��WX�NR�l1cK�L�;�ldF!"�L�H�m���cgq��7;�����.���9]������q�$�匭=So��X��9�OI�芭���Y�t��S��x�}H�hl�KFM��x����f���ۦ:�	��5�S���kf�+��i��V�}�
Z^0�m�n�N�Ul#z\+eM�NCW�Vtf��ZY'��\D��-�F���;b��f�f�Q�B4���s��u,ӦKڱ��7�)u��[�D$�%��Yۅ��ݧ*Q�y�e�̆��^�p��o#��\���z�6��i⫬�p*�.�nܸ�1�����8c�i��.�����V���[�	�F�m=�.X�Ta2"��-�sib���%���A��`�s��1-�Ve���{(�n^ef8,�;{ll��G�t�S䍛P�r�գ�d֨=��%һ��s�vi�7������b�0�Gҕ���������%�]�,���R���y-7����\�1�EL�Ҝ��+�Aˀ�[�d ����ksj>Xj5�� ^6��愳)_*ѧV̕��K�;�$��i�����s/������:肊JBwlF�zW�;f����z��.��Xcz����YL4ӄ]H���c��9�|���4#S�PY�,�Sp�����=
V*7���y-D�wVP^�u#��E�����ˇ+�4�-	����A�BT-S���QC$�����Qy��[��|��E���9�
�=�{�^eURR�
d*�A|ep�P�I�ȉ���x�ʪ=�'L(�#D*e�E�C<��udw��mVF�IF�E껧󻻅�f�jb�9��Q$*<���8�
�M�EEQL��"��ZNJ����;�nC���\��Q�6Q�]��E&RTUGS.*܊)Ȏ�*�O��h��#�����Pw3�g�U�R�P0��V'*��	VG�<�y�rԗ��ů���        j�����񎎼��'F�N��٦����؋Cŷnf�Y��{6�]e��T�[�n��2nd�'<���5rY{l^���^��0�I:<{�Gnj�=vW�:��K�w5�l����> l�n�;�����=ÆÙS��l�����#�	��O�ܠt���LM���������<V�4F��Q��w>�p;����5��UYu!��q�I��؍���T�:ܜ&���]n�h�kwa1�,�������lY^A�X7��^z5�b-�sj�s��v�X�ul�zx�7s���%�v�!s�2������ƻh�N��-�m�펷���;{kq�ux6�d�KU]���-kF�8a���I��`mM�nι�ܾgn��M��˻k��vYv���7<��S���s;n�̬ L�n��]���`"����'��X��s��v���9�p65�ۮm�ݣ���:�ϰkj�o��Q��0����Rqu��h�s\!�]l�uYܜn�2��w�{e�#v�K���vD�b�s����YӉmn�a��S;��v�g�';�qͺ16ޠ�.G��k�R�����o>8���=1ي[}�c�[�$����8m��8�C�V���y��!���]]C��7���0�ѕI����{$��n�s"6��.e��4�Z43������:Dy�7��Gi��{����<��W/GH�Mb�{Voq�h���j��I��ơ|�s���L�7��9��tenq��N$����:y-�
3����{5���4�cLmNu��Ǔ��]z���h�'��[����
�<�bX�rv���ԇ<�]��ޝm�k�s�팦b�&w!ѶwV��l��u��ns�9+`�0�,��fxk[:h����"tz� �!ʾ:z6ɲ�qs�
��:�:u�nY�n��g^��j���֪:�؍)�I�n��;�����=xNzi�
��T�\��o^�ѩs���v`%|ZY�{vG�q�v���{��b\][g�:�O�`HDN{a��o�n��r��۩�nW�����sͣ`�l�[��s����a����uD���h�ɸ�:��=��q�ӰRl��4�u�N���]�?~�}����1 ��H&�6EI����R����<T8�H$��@�J�v�� ���� �c�E�͖r��� <�ɂ���k��S�����f��p�
ɀF�$)��ڣ��ܻ ��q�*�S����*.��پ�+fxr"����АS����a��޻�P^�&I������$unL�.��)�H�T�A UYI
c|������{y��Y��8��>'���`�K�ɠDVo9�o����")�u�`���y����u%��z��kz\�\mQHL�9 ��l�]�� 3�ݒ.�&�V��݇�4�ڠO���Y�2\�R��L�`��t(��9�Kj��wр��y.�c�Fq������7�o�d�$^��w����0��T'e��̭�ر�m�G���>���c���'{~w`�h��f��j#}����k'�ʠv�R
�]�5ݶ,��O� f�3��������+᛼�X$���$_B ə�yW�������a ��;G%�A윟W�3�w�B�����y`YG4�bE�v����L=٪:��z�׽�H��� ���scw\q{���m�n��.j�dٝ��S�ƶ��e��8��%M�i�*	��HW�u�
�t�?Q�$�s:��]F�lG��f]�Iv�j���H#`6���x�	�����-�y�(Cg�0(vg� >\m˴����s�O��u�l�
�*W��l
�ϤW�>,Ao�"#�L����`&Z�Db9�_-:�,�� Ȩ�<�ԯ1�єR޾Y��z�I���I�{�������>=��ٟ��<���Q ��a��ݫH�Ҫ��:z+Ǟm
��������>�*9�}X�|�̠��!��6G=�bߜn��¬��y0 ��<�=��"�mj�a�(���[�V�v8��t��s�ף�����)��U��0"H���;�˾��|{qϨ���ݘ�ʫHv� ���x��uP����ʅ�*���A��%A�^�9y; ����A�u@�A�|�X&3����]�َ���Q�H"�6m'ܢ�(پ�  �ɻ��}s���$�|��1b0ʅ0f"dls���D��b�h	����vL\��w��Σ��Ƈ��u�hh[(�m���[Y��t�<��������������{���P#Z�:��l;���~���%��F��H<��@>��m�D��rP0�Q���vM��7�����:|>���G&���Y���wX�˲n��7�u��BfT	��p@��̠��!�� ���Y'ė��?�ϭ迦6���u@�|_�s� �'���j�+�'ϤX4{+�]ܦBU��$-!�:�Y �� �t�fH�<߉�عQ�LH��ex��e�H��>$�nQ1�j/�t΂	��v.�����[[G�Aٵt��/,��=��z�]�$���^'Ď��ہ�f��˧C"�s�R����� ��@C\�hQ�&�:h��ξμ�!�>�$z�&� �ٝTw���:�V�5�ј)l��kWՠ�v++�ʊe��u���jX��[���"¤�������w�|u�� ��5��v��5>�I�<����lZ=uk��)�F��C&�T6��)� :�M�)ٔ�����G�.���M��j�����w\=2F�[s��D��ո�q�w1$\�z1����-���@��J!�K�si�8��.��i�ǭl�}y���vRur
\qc=v�烛���n�j�mϋn�Ũb��"�6ٱy����V�˵�cϏ�>�Wu���oa��i�o������y�"AS�k_�$���
>>#�:����3��3����������!b�2h�ť�l���%�2�TT3=��@{3́T�x2�Qr^�sx��صV��|*vc���{�S  /2ޣЦ5��x�hft�v.Tl�"DDL���n�1�z��.ˡD�q�$�ϞY����R�fdʒb�r��:�wc��Y�� �`̠:��?Зk�h�A�ߝ��A���j����__?�Ψ�ޯOn9�s�v]�W%�k!�V�/#˷i��"I3!U��dDI31Ox���o3��ľ|�Qmdc$������A;9��y�C��7v�%�W��ꂂ�I�t�s��Rnא"My��# �͡�p�]�}�m��m�vT(���QLS�[��ɚ�@�g[��Y_�*;>�A��dP$����`�%T�lJ|z��A����<�����yD=��	��wdw[���5���΂�Ϊ �A|�ݗF�P�bDL�I�"�39�g%'�Mm܊$���݂A%���=kj:u@Vdm������F�%Lt�H�yB�wrF1�TH'��u݃�K�@��\�P"��b����]��.�\�]���c���͌�o=n$u�lW�������&!D��Dv>wd��@X��׭K�ݡ@���vG)��Ȉ�fn�T���/Ƴ��J��t�}��O����/����fI��}�]��T����b}vv��Ő}��
 ����bb�n��\gnv��&2��9[^�վ}w'|���a|��%�">�˦jUV�fVΙX��PԾm_ĒϾt,�����B 11(�Νy�z	��X�ɢI�ά,��;�(�n�H:���*��%v��
���I��0hVј�5A>v���H$��󨟷�`Ez���F�J�����z�S�;+�Z8ջx�6���3�3�W??�����%�EZJ�@�d� +s����uAy\����eJ�����m�_�@$E��s=獊��wv9�dM�� �(N�L���<��|q/�w|���t�w��&f"I��4H7��@O��:'KǊx\�n��/q: ���g��:��DD���z���=����9�ǉLf�x>n���K��5%r�u�Fd��Vٷ.��ϲ��xŋ��_I�Y��B"`Kp�lވ؆k#-��s��f"A��&7���{4H��C���(��0��n���{,d� ���W����v+���1�z�I��v�X��m���{[��Q�gW;7\�O��n���ᏹ	
L��W�#s2�D��r+Ē�v.��-��r9Ƞom��vdǕ��@+V��~��:�������u��6O����`�5��ܢ1<_l׉�L���I��D�}9!���b͓B�a�Q��&���}��v�u�Wh��>�����+z�D�$�N_1=��(
 n{�(wdV�y;��>m:��v����|:Ot�(
�[�����qzp+]�#�T*{�eJ+s�h�
L��g��v�G9R�[��b��M����ʪ�VR��ͼ���a��$��Xک�ʽ'l��˻�6V�駾�������|������>6�m�Z\�2�H��[�h���]h,����u��9q�`e�:��(c]1��)�v�S�f��.6���C{TZ��Ϭ����9}����^��8���ɹ|��Ͳ䪕9W��X!����;OU7EݗX�����y{,pP9��7]Jqz_a޼vxԍ�68n}���(�=�,�[]��f�nK�ۉV�GX�C���|<ќqU]�ܺ�{��C<���ҕY������ �h�Ľ�=��}�?Ux�s;��ӛ�صa+�d�S���Ο�ن^H��9�8�:�	y�4I�;���#&�ΐ1|��E*V�|:6�|+s�MI^OB�,ފ����o]��/;1�����
ȫ�FOy�wL/n�4I������vMOfuL�oI��Q��*
u�𪴨$m�yv��>�3<��z�`��<ܓ�*��f{�^잡�϶�kI3W�"��F�kɓ�{�]<+H�-�ӧq���<���7~}o�ߋ��(��D���U��٠Lt^��ܷ�����$u ���N��5*��t#ʄ��A�nU�P�b.[}���v����̧ ���V)��4gvfܔ�r���*P�fLsu�����:��B��)LA9��]��`�I>?f��}��u����<�rPRh�*-XJ�N�t��f�(PRmʼX�{r�ӳh]��N�fy:�!|Q��r(��j�n��N�A�(z�'ǳ�$���GW�2k$�74je�.d�)��]��$�|�X�,�f�tE���{9����P�����,�Mc�V�6|[��m��{lhIś�����7Yl��_���?�"d3�=�(�/3f�'��������r�wD��~$�wf�x�J�Z��"`�S;W�޲b����;��Q$��A%�s�~��XySי:N�!b	:eD�1��pI����&Ǡwf��\u��}�@�<r���M?�{�Uijt�($�#HQ��{��=z��y����@��^�疮����j��R�TJ���حN���ix�]�4K�|]��I޵��+o�#�
�����Y�a�����O��>ҳ.k�2�/t��-�sv�[��A-��0Կ�y^�Ԭ��O�L˻w]��}�K>yl�l���չZ+��yN^�wqh�� ����ᡎd��'�mn��F��&��B^�*)v��:��}U��Z2��;�p*,�un��u� �Bj]oYr�,�9Z�v�G�2���DG��V�_R���5'3^DX�+.`��[C+*����i���HF�9d�byրX�/sg<�E�鮼᜻�ӻ�GL������k;3�b���k���+��C�j���x���84���B�,w�9;�	t�VE��~�b���:��n���;&^)��-�:�8��z�o@�����Yi�6Jʬ��y9i���y�5(tV��ȫ͊�YՕ5�T��j���Y4:���/����T�Wu�Fcg&�-a�3�-m���Zm�׎�L|�d{�Qq:���]ss1	q\�d	�LAj�u��9x1�؏c��5�!�Vqt�C�A�ٺ� h[n�	y�])	�ٿb}�ge��wH��	�i��Gwy��)�cE�tc&f�K1
w�4?	�#+
�I:���$�f���u�gJU�ww~~{�����]P&�QW($���/�GC���\"A^�f��f�'3#6TM2��'L{�����#Ídm�t��=��*:�Qʇt�IQy�t�*.	��=$y���Q[������)���N�+8$�*���3�YeXRN��tTILMB�
U�\�I;�%EA�`Y!�"'CB�]Q�+%�������AQ@EUT�R���9ˉ!듔\�Z�l��Ga˞��eȯDg�fC�TRpҙ�"(��
>F�,O�t�ʨ(�K��r鑛Ց\��dr;*֕UQ�Awwq�8��s��8A�Y۸�Ģ#�:�8t�r穝LH���t�6Q$Tr�~�}��I?�m|l����w��H�A�*չT*vg�7��%��J�">�� vn��	y�N���j�z/;�@�n����*TQ
ժtt�
v{]1�aOt�ʋ�6���@/;�I9��=�:��s���g�)]HQJ����*��t`P��U�r��YvZރW3uh��}}�}�n������u@�7;�H��k����w/|�l {����xU]�V�:�9�a��[4 ���s;��¯<��,��Yt��4R�����g����
��^�='����46��J |3=���D� j&ҡK��ґ�\���ռ�����^$��Ή��q�� �c��{uyݷ;��ܶ�%H�U��j>d��/yX��n��a�9���+�Uv�n%���cǓ"��0﫼��ɖx�|��U�廼�3<ְ`���˚9��C�q�Hy��	$�sD���zTn����` ���}j��F]�=g��p4�m�:��m=�Bb������߹߽r��)Z�M����g��@]��MD�_��o
�{v#1��ML�'�HR���d�gG��ّ��P�j`P$o7T	*ͳ�"j�][�Y1 �dH�@ �X�oݮ���N� +�1�e�=Et�$�sD��7"�����J&H��]�vo��'�mv��� �E�d�_7TH$����*]���vl׉lX�]D�T/��>n� f��ߩĽ�y� {6'��� ��H���*ŮG����0�,�m��:�nf]��Xn���dgVXT%�6е�~�3T7�r����c��ң*QʮX�����ؚϏ����{נ���[ot;K�m�YMی���v�[�;�Mն�v���O��Y���Gn8�h�;H5E�{H"���Y�a�/F��渡F�m<l��p��[�G�S���I�ݲ��[q�umK٬��kC�\��λr>�\��t�\us��6��g��������=v1ӻZ/[��9���:Ʊa�z�REqY�<j��A;plX:������d�a.^s3��ѳeaZJWw�Pū�PK�|*ne
 ksG��7��+k:"N���M%ƺ�K�2Dp�!B*f'���&�����"s]a#���|C}��m4}Õ�\̭9�*m/X�QD��J��wT'[�b�#�#L>U�¹��+��H�n����Vb�Ȑ�Q12h�7f)w'r�S����k�Gf�ʂ�=���*����<݀���3�ۢ�$<n��ǌ�V�ȇ~'��hQ �n��s9�'U0`Up����\�-n}:�X�y�3�t���7\n����[<E�(xp���d(��&s��A}�m�$�Z���|��"oZb�w*����!ʏ|P�ѤPJ|�M�(I��n��s�j������o�_�o��a��B�ε���u}H縍�3��U���m�*E������Ɏ���dL�F�������#�Iw�vH0s>s`��1T�����ծ�7V$�bD����^+on���Q� ͞���X����  ��t�@3G3�Sie�ʕM]�2V�c���"��M'��}*O�6��M�eS�c_��}�̕��AA]	��+DRV�t*�������.����;�e�5ٛb�$y�h �F����$5��t�Z}j����5�v{Ln�o�q �|�c���k�n[������fa��n����Q'�������7:͏'=*P��ژ�MO��"RTo��/k *u#����ؗ��������s���|-ܸ�W���x/E��$�F�A'��1��� =�o_i`�k!Ȓ=֌��U����zwN]��:o������:���#�>�@�ܦ�ϷVD���J�v�Λ�N���ۜ� ��\�#*đ�!H0�J�0vzuf�Ϯ���U���(7�hH9�υ�u}[�{��I��"�T�R$@2�D��ʖA:�]�bW<�(��W�4	%�]z�gs�4�oq;Uv��%M�ֽ�6���tg���qj2�T�s�;N���i����TH��&fez��
�u��A3���-�7�^κ�s� �bb��U���,��쪁{1�������` ����;q�l�Y"r�̅T&y�A�]�'OG="6n�pO���@���X&�L���A|)�a�^^��x��	�(u���D�׷v	�����V&B����cBԯ�m˸!&£��nϝE����
w(L��m��ǔ����ةfፃ��ȋ��w��Ϫ�*�%̅ �*f$Q[�]X$��]Vq�t��֠"���(=��(Bg�:P��hȅ�.Zx�-�:tf�9�/n:�ݍ��yk�Ӻį^���[��H�eB�Wù�W�$o��  >���f_�	&�tBoq)�n��]��였lFĈ�"ffUx�=��D��X��"U��8H'����v}��E�*�l���׷^$l�G��ԨB&}j��/�Ŗ��2{r�u�6+��H7�����s��B�D��̅W3�T��(@ޝ* (
���{=�'��_�=iЫ̞�S���Dn�E����D���f�����lv��hTN]�>$�nh	��TI��6,V��v��Oz�欐Ҿ��R���ǭ�}ѽh�b:Pـ��Ź�e�sYQ)�Sc��3���g��iu����n����WI���\�n�^��xz.�����f��{�m����%2-v�;d��q�收^y��g���p��[8��LkuP���ۺw1�܅��۬ ]��j�ݍ�Z��]�3s�F��d������ȹp�mPa�����ր�.k�^���<��&�[�;�Y�s���L��`"������luʻ��gA��A�y��nl����j݌�lUh����ߍ�j��mZ��3�|�g��O~��Ng�|�KY����?�3����oo��� +��퍊�*ޱ^W,��H��ŋ.�������u�.�f�,�I$��`��� �b`�5�����D�=�f��E/{&�C����DϪ�پ�P�?5�9WR@$�����1��K+FWW�+ʀ�)$@.R����Gd��No=�n�.��ghTD*��� �ܚ��=}b�y���������s�'��Z]����k�+���u�X}���t�#4{��^�-�ڟ^U���'ĝ�D�A#��=�(o�A.n�T7w���еB�6�S�{����r��G���*,gp=:�x#\��P�-�$���K����I���W�Tz�;��v�3�.���å�Z�)D�~�r��$~��o�?��,�Mv�6ݻ�׭�+}~Wf� �FJ�wT	#[}b�&����꨼�p(/;�(���PP*M��RI/�v��H��D�m��$����w�$�<����o��� �6:���
��*��'��l�	 �/Ф(/���N�նg�$_]�Ay$�cآm"s<���6�A�8�j�J�	F�rt�r�ƴX}����ӝ<����~�����bJ��ߪ���!$��=�BJ&���L�3;3	�<��A2����s�>�7@��$� �,d�>[��^ӥY�ttI%���$�K3�i$���Q@��wО���hZ�dV����BH ny:dM8=FzvG��� 1.�5���P��Vj�pdۣ1���4��^e�7G�[�ڌ�b�����<����~�չ�I�q��,E$���f�27��f�U�V
'2�g�e'ˀ'�'�(h�@���d�9�lz�]����7��P a���b|TtI��!
��2<��$�3ۮT#T�lz���j�&�.�D�$���I$���v-cb�C���z��� ;���k3�[����΍�>���D�Q!�<�"�0�D�s�չ�6JH��d�I ��:�	m3���ƻ���2�  ;<��OӮ]
��IQ_K��~���~T���mdP��w<��I+�wD�\�M8�zn������,��� � ��)p�;�Oā��r�"A'�9''+*���Inl�$�&{�$'r|�mT.�����=��ʙ������g�@[ɲ~$���n%��3�N�g2���&���]W��y�C�O	�S�Μ�ݚ�N�noX�� �:l���ϖ9eu��X�BwT`|KM'D�ie�+��PV
&J=�.�6��ݚ�˗fE.m$�W.dM���h��/�f�dE�+s s2����Bvع�{&�f���]]�;t�L�Q��g��jխ�uj��R�Fx����$��Y�����{�4/�Gp=�D�^���H�m��ZJN�@.L!$$�_mZ�Z��y^���*�ۙ4�I�wv%$��n�Ix��U�u�<�3C�!ʺ@�3O�/ʫv�+I�}��I���I�:����4�I'3�%T �I'}�R��� n�Wt��H��L��#�TU톂D�ͫ�A%��9�I�Y}3��z��^�%yF�]�	�/��%$����#�@���O�,��*�4�K���I$��I4QI��Z�w������(�/�� �ϼ�fUPQ��-�p`6����@�	!W�H�t �1	uH��I��e{�
��TQ��F弧��,3���V����L\:Q�QȌ��B"�(�z��9G�]���w�gy���x �"�r �D��B\&� `c � A�0 ���1���Dclm㍱�������H1�v��nv�	� ���$�&��f��"8�z�1����vĩ��<����1^T�TH%1�-�X�����S��m���6�>�O�k�c����u���H�!��ڰ��!�U�cTŅ��������W�")�U��6��_V����*M�l(+%P���7�ރM��
�Q�k�{� O$$$���=�������P��g��Q%�� BB�0b؏��4���c;��ʙ"౸���~N���D�������Z>ԇ���h�?�}gL�?�
(����>��_�����>����G��HL?:���l�_�Z����CLb�?!���C��@�l�m~ X�qp�o��0�ؖ�J�~�?����i
��lB�JL�4�k�O���>��R7>����d�)�������d�!$&�}fT^LX�Dj?�^F\$�H�$�hJ1I,0&��������b�(@�|Qm����/��>��_W�?�Y�/�!$/���021"�`F$6�*_b�:�?�/��A~'�`|_��������������Qq,���m��>��0x���R_���2��!�X��A����_�.m2����~@1A		$���҈��	�H_R���?����}G��`C�������ZE��u$Q�(��?������+�o&Q��L��H����ϰ<����
>���?O�?�l������B�S8}`��h�K��_���x}�ׄ����4�� �~؇��Bc?����I$&����I$/������CG@f�п;�pGڨV_����K�Y�Ӂ��H�"�Gҁ$!$,��YLm����xT�>�$���3 QB������m�_p~p��N<R>,$Œ�2H����?W�葄�@�&�4A�%ա��6�o��Ұ8d��BhP��?��C����~��B��Y6$!$�� ��a/�I0�ԿI����K��~��?���/��������p����~�����A��H�H�O�?��p�#�c�q��Ay�֏�A�~���IY��Z-�b�M�>�����_�x�BBI����}����pϹ �LhcO��8��?_���@��	I$(���!�S6����/�@�~�>�?7�_�_��&>%��>����X�/��~����`u�C\ aHg���Q�LbjĨ��~���Ţ�rF_�����hi��m|H�����,/�~�_�?G�`\���M�������hHBI!0�f~ �8,d-�C�G�}��0�a�G�����Aч�Р�������,__�>�	P�(,~&H}�L�� Ƀ6�?�#���b!$/��1 ��"�>��G��+���}��>���BH_`�Y���K�C��}A�~?�V0�T@�$gu�#�
�K����g����3�@h�>������Z_���"�(H##� 