BZh91AY&SY���t�|_�`q���#� ����b(_                                          � =�   �
 �@ � 
    (@   �  T             {�EAH�P��H%PJ��A*��TJ� �$��IH� �
��DT*+����   �)!ABAR��H� >z�;���,�ʩ��	��L(�t�q���&��w;�U'8PQ�R�v:P��t}` � 	�   >ܫl���R$�V����R���ޕ	z���I��o.�RE�W�]����� t3�ht��%)`��r 9 נs�=
z;�
��   ����(  Z�@�J�Q@���MU|�՗�����w�:xw/`�yǂ
�҅3�������i�0��Ӡ3�xK�CAt�<��0=x  ((_   <�}���e����(��P�� n�ԅ���n` 僢K(�ঀr���u�ׁT �_   <|TRP�I*U ��R �� 2�݀:�; Y�$V dq ]�@���� n(�0�c�:|�  _ ������9� �T�W �Ð@���r�4�t��X �� [�7X�� z�   � ���RH*($UUJ��> -c� �΂�� q�B;�R��!�v�.`�� 8��E�l: ���@  (�  v���0��P	�N����ݝ�qNu
S�0�� �Šm@ �  �|�%)E(���Q*!$< H�@ 9 d� ��I\ m����;���tP��:dh�>��  �  gO��F� uw(	p ۸�  v�uH���� `9���@         O *T��     ���E @  � 4�j��T��      Od��5E*@4    	OԤ�P�  2 �&& �(���)頌)�0��j'�|����}��m�}����w��wp�Y���y�;}J�(�<<o�AQ^T�(���7�?3Q_���G�����'�������O����(��<���dW���I��ND��}���8Ȃ��Av@ �H��
�
��2
?���YU�D"��D]0��`Pt���tȂ�E�
#� ��(�4�:e2.��L�Q�(�@� `]0��WL0.�L+�U��ydL��@4����t�:e2�L���t��dd4��`2�GL��Q�*i�|`2�L`2�SL)��"i�4eL���M0��L���t�:`_GL��2��L�� �4ʚaOL)��4ঘL�D�*i�t�:`SL��P�WL���t�:a2����/F0��P�*�t��a^� �
�t�� �q�t�� �*�t�:a0��L�ʚad2��L���(�ym2��L��t�:`0�SL��CL)�T�
i�x`2��L�� ��4ʚ`0�S�D�
i�t�:aM0��A�(�4�:dL#�A�*i�7d�*i�t�:a0���A� �t��)�A��t�:eL��t� �t�:d]2��GL��	��� �ʚe�4�:eM2��GL�L�L��T� �8dM2&�SL��ވ�
i�tº`]2��Q� �eM0�L��A�*i�4dQ&�SL���"i�4`M2�2�d0�v�*i�4ʚaM2<2�a2��L��tȺa2��� dCL���"�za]2��L� �
�t��`]2.�WL�i�|`� � i�tȺa]0�� d�L��Q�"�º`L i�t���`L�� 4��@�(3�"�d]2��D�"!� l��2"�����+�ETB<<A�����x;��<^z������~���W�G	��x��T��ㆍڱ���K�8�:��ew'ٳ4�(K��[ۘ;o6��
�M8MM�x��{�"�d�T`�X�]	 �l�\㛊���6���/ݫ�%��R ��g5dH�n=���FI�и�b�UM`ߠx�7��(�3r�PaEJ��V]�%��`�6V"ڊq7�[ĵL�2�3�B����KDi��}�d���|,�׊ӧ��<�;�����PQųb�ʾVF؟Y�iML9(�p�C�Z�sH�h[�iq��'b�9���2'1^�˹�I�gL�M(��Z�%�i��3��n=uv�[�Nq/
ïNS&�{8J��b+ш~�""�]6n��r��=�2�䀜�7����9�����1.h;5cm�˱l��]� @�M�+���BR�ٮ3���X��\������K���oTn;V��l�[��ӑ�9	�'n\3�X1捜vDI ^�h�A��-�N>�W=�nmVq�3�C�ғ�X���N���w>K!҆;����Dݫ{%k����nl����{�u�]��7��vֹ�)'� �������޺eX��y�,烦^P�B��x@�7���Dpv�����@}��=��W*ܮ�S��Ǟp��+rm�k[~���X��f��웫��U�qc[�!1��=|HՅF����N2e�^A�i�U�w��dةOL�ٽ���]'�%D���7G&,4��\��M;�&#
:4���G��7rr�i�th���խ�[m�\�7� .��l�n���(��Zh�.�yV�Я��U�7 �f���_����Z���/�K�Jc\%���obش��ʕ��2\����p�SV�rf��'��C���K=���w7T�[��F)�|X����ZU���lS�c.�Y�\���޽���Gy���kۚ��Yv�i�A��DN�7S2���Ue�~��]�r�Y���1�8R!��wxގ���D���跥����ۧ���-<�N����vU��s���� �ؤ�wl���S�wwZy�7����K��&v��.���cɴ�w6�`V�8��B������&uZ�	S�,!��C�s`�Xy�7�q1m��w���&�m�T*���Z&!L�P��4 9:�S�����4��)��Vݫ_n�>��sj��%�hR#U㺄��8E�-ԝ��wZ׹��<
h�{-�
��h-Von���I],�gu�a��p0L����R��5��1;�lu��0��=~��E%�86>�J9Y���l����x��0�3�2�O�Yl��n�<���{���O	r'���׸wv^��۬ϵ�0AV�[�ޏ^���ٔ2�h{>;+��\z����Ĺ��c �<^s�Z�k�
v��2S�>�d���Y%�x�Hę�6=OJ�ot8Q;�V������ۿ����� pߦv׸7�G[��y ��=�:���̺p��,w�w{�̅��)�	�k泑�CN�.�5�3^�=ıGՠ4�J׉5���1i�lC:i�+Q����<i�ёG�h��5�f�6� o���{'5�v�;�Αe=uc��
�nO@]׳B*�q�w;&�.�W�!�ڷ��m6.�48���wW��BSɳnrÃp��·"�g�����Ӂ�嚉D0���"�����U��!tĲ�a��p�7/۠�ܙ�;�Ҷ`�vC���j˺�ݐ�1�3p�����)2M��ޫ�0b[��N�Cɝl
�Ğ���f�ZN�=�Kњ��r����@5�I��W���H8t�ѧ�A�7b}�K�p�`4ٱ|zL����Y��v����¡RL؛Zbۻo-�c��1�n��
�q��n��v�L���z��d�7j�9WQX���IP)�o+���8"��'}wt��3,��mWe�|���r���{+�2M������a�qMeN��Fd����r��tu��Z+op�On�\%�ww��l�w���2j6-�/&�t���`��ݬ�[������4��k�]��۷LYؙ3"ޛ�u=v��6���J7�ʔ��2�-ä.��v.+���b��GL��������SvKA�V���.=ۆ�����ҙ&n �;��4<nI�h��Ű�os���ަ�������.�s�0�\M3u<�8�`���is^���� ��X�JR{s�O6AP��f��V�kԀ+#�&�Ԝ,�n��j�(�|���tafB..�t��3K�7�ޓ����j(ɼdk�Q>�:�h1⽴���d�k9�Sy76o�h�M�z�ÔR��wec�:b�Gd!3˖t;�KEc������GF�S���;B��tr���5�<�ӐG�GN<���w�^ǝ�,��e�9ې���Y����I��E�=wؠ��4d��O�T�eˊx��rtW���%dX�!�'O�l[P�.vmpq�p�$�J��5k�����B�0f�f�Zy�����b˓#2�#I�ܰ���,(��y��@]��ih� &l�sCa8�<gp�͋�;p�7;����d���ά[z��If�چ���HS�2ԇ\νۂ��뻼�sX㸴`I��E��v��f�֗ ��z�"�3�
d�
�v'�w6��B%Ǘ��;��M�o<B#�R��n
0��qv�nw !�z��ݴ�9�M�LZ�f�>}�o.���@��sut���ӄ�+���tpV9fԆi�a��٠�僫r���XI#���Kv����Ѹt��r�K���ۑsv��Rt��u蓎�[�n\�.���m%{.O����Ӛ2$�B��jNT�]Å������ ��K�{q� �.�������n��ϵ��.�s�~3�W85�R�>�&B.v���OJ]�Qk���Du���	&�9I�<�v�c��)6�<4N�PQR:�l�y<hr؞r�7:+���	p�$GL�����7hj=�Ӽ��w��,w��>���4{����/}�pZ9�loSx�զbNo.�ݻ>S���.��5v^��wU��b�%�i�T�YV\u#����mv���� 4u�P%VF��5�/�`Ug%u�݁i�B+3ynh����!:ȶ�sw�ް+���M����'�5������!�GpVߞ�Er0IR�#ӳ�ݚ	�;Nt&
��W4�ֶmf3���|Ԍk��$�q�0�tke0:��щ����4j�x���gg}��=Ug^W�/wz::�I�fᦡ�>�$�R�]Yz�#MU��S���Ë��}�Ȏ[�8�Fsx�B��:D��c8hm�Z�w`�t���뷖':��������xQ�J��-�<�Q׎S;�K�r�]r����#����k���F�Z^2Xy#ߔ����
ELޠ*My�m�Z��6oMXk�;�;-qn��t�e��M�J�{R1��٫s7	(�>����V����1�х!�o��#&�* Ӆ7�o`cr.gr-�t�"}�:w)��s�l*Aș��P1�w:V�ma�\�ON�\ha��8�L[��;�opwyv�r�]�l��s��� ���{�w��1u�q�d�;��d=�����@���mOGA�KAo6�X���;��ܢT#���Аa$�R��4�pg��Uh��˖�$Xݫ�Ѯ�5���R�$
�,���wq)܇�i6\�!A����g7T��<�Vr���c,���D�Pl�LNrq�B.�3���N�l�e��MZ6�˛��Ncy�n�h7y!�ϹwhQ\�³S
��#����'.e�3���f�5���i��f�.�i|�]���{X�]�n�$o{g�F滅&�v���C/l��/Ww,Cq빩MfM��f�����L�S�L�5mֺ��pRDl��p��9�ȬJ�WE����Bܧ4D�����,�:_q���[���TNF�'<R�ֲC�F��3�<fG3M]�܃�!���@v�#{H�C�y=���6��j���n�e��+d;�>R�K8�%�;��tV��2`��DG6먁{�3@J>���±)�i�B�K�{�[��o!"�u�nj���%�#O�cK��1�硗�8tCd��e��wL9���	�C��`|>�q�voVY�4��H��Md�n5�RVNL�e�D���k�M���&n�/Y�o8;kaMҦ����h�=J�2��ݜ{s^,*f��C�2�}�pzp�iKh}�;�Ų�y���e���"ܽ���l�wg
���*ߨ�l�ͪfm�vcٜ7C�s��z�$p)O��ˆ�w�Zr�+ѶHv�9�/y��Q���_t5����u�˱��)�ӧv�9v��zյ�2��k@'`���iᚖ��C�Du8�2C1u!��T!��'4���+u��m���H� �7�^��钊�}oA�㽃$�XÎZi��#}ӱI��+93���y.�\t��Eʹ��i:���]e�Ԯ$]���'�kK�ෳ�]���P���q�;n�=qÚ0hT�Wt�4-x��%h2��͗�Pല-����mtsv.��x�k����Z ��`׻6ܡ�0}�$�B�N:~��裹)�Ѧ�\���S�%�aMN��7W��
j��]��Ago��9�+�ҳqI���5P:�-k�^�qťaX5���wr`�����I��F�"��=����C�Iu�˩,��iO�\{�#C�n���8�\g9��R��<���Z�#�-oc�Ӹ���We��Rw"謕̹�8�Xi�3��6yP��޼�9:�� ����Q��p����ia�ޏ]����6e�o0N<a���ɻ���Ө׶;�������vrG����E5��r��m�fˤ�׽���e��qM�7�Vx���� z�	��!ۖ�s/gT9��Ǫ�
�����]�{��(�Wݧw�����q��ؕO��=Ӯ�ǀA�Sk��e��v�Ψ��t��W���;����rr1�;��ӳ�����i���ʴ���c�_v��P h�>"d����WԱ��N;|^�OCF�y��͋Vnl�ڹ�Z�c��D2�wp/E�]�LaӸ��&h��٨{`�t$�vtZ;~;��d�û�u��U��C͹�`��Jy���i��
�Xԭۑ �8���Bǳ"��k��2�\�r5u��#�ڷZ�E�:e,m���d���aY&(VǛ��T��������ӝ�TV�V���C0��5oq��0����o�y9�w�s\a�;�"1u`�{�WN�Z	_b�Oh� os�M8�M��޷n�z����G�_t{�Z��hx���gv􉑔��F���ɹ+7;~I��~
e�c�휟�v��k���zv�a�m��p^�a�Jthr�{iع�s����PY^��A�:�·�L��[��\�̟�3�f��zX�nT�Շ{�;�Kr�1i�&����؊�˙a�廽�ٝ/ �o3ub�f��%����{ k��P��2�՚�"�=��D�����2�=s]aJ�G�4t�n0��C:��.��v�d��P�ƹ:��qɧ*:s���B�G92����0�����rg���i���Od�lx�㚏q��mu���ЍX�ǝ��N��/j��w�kw`�T�Z$y����Z��y��G�B81���wNk�c�H)��dwBk�9)���x��P1�{ܜ�HW��<ׅ<�xY���"��զv�Ov��������Ú��x!^��a�4�3q�]�v%�זQݍv��v�N�]�9>�.��ٻm����VqH�7��ï�[؍e�YeȟIn��kvV�w��Y���:��:���nI�*�@z�a8�=ope\�L�TPO�oN�&��p����)Ή>�R@�G:�02x�`u|���3����Wt�dC���G<�#����D���v빻=g"U�2:nS�tٖl�rtfMM�؆'M���u�D�]�J�J�Nf��]�U�^�2�V�ι���7���.8�;�LOB��@�E��B���*�k��|�T7@��s�y��yv):wL���͝ɸ�<��t�(�p%K�N�i	�Aڠ�s�]��9!!�b��c�e��I�ƙ��$�Tro�>�qېe��E���e��6�oM,�h:��Ŏ&\vXt	���Lǖ0�3c���w{z9:n�W�b3����ԋ�3�V����`Y��Y-!]f�\�%���<K&�I�p(W�ä�1�J!�k-nӺoId��'I'p*A$������<Oᚏ��J'��Y�ŢY����l�J{7+&�Ų�0�C+���I4�W`������	�x�%�V��{�"4�'�^�i�I���3J%q�/ĳ�GM%`�}���O��p�n�w�$x����]dഄj+ �x�y�������ѯL�Ē�8=�2��}�瞛޶n�n�W7X��|K&���{d~'��/I�I&I���x�1]�����c%�x�f�T�q�0���^ �$B�y��8S��8��N���?�HzM�ֵ=O�a-�=�-��<��qB�	�<I/�asT��J���?���' �̾'Ē�)��k�.�#^%��}�J��B<g	e��I<H�)�2�I���.��O�G|^���~y�������´�����YLDL%	$�2M��?3���Vf�}��}{�����8��>8 �ʨ(@�J!B4��d"� AH�@�H���ҊR(R��ҠR���@ d &J� ��(��B�BP #B.C��P)Bd(��J-*�@*Rd�(��� �4� &J�P��-"% �R�4-
R�ЩH�H��R�R�B��R���(�J�(4
� "H�� � P	�(d*P�@����!B�"&H�J���P�)B@(�R
҂"�*H" )B%(����*��� *% #@�B��S����<���N���'S�N�G;�P�;���{�{!�@o d�\I@qd<탼�do:��2:�i�|ղs!�%o�x9�ym;N�<��!��o]gp�yO�Bm�u�a�;H�#���+�wq�Gr{ s�%��@e�w���q�|d2<���c��5�!��ְ;��� ������(���Y�_�uQ@���o���A?��?H�*� ����3�������? P,%+��A��p��h�t����y��S˴�@�
QX����8C_M����[������5��^�c�cFq,�I�1�I�󺪈�/�a-׶!�y�k�&��sܒ^��$c7���;�M$!p�~����0��;D>�$��j�t��[˯��5	kꔵ�ܾ���]�.\�/ݲ��)�ۃ��r�aE��C��`�R�C�3��-5�b8᦬`�����'(��>�����s�ܙ��N����{w�����٥x�u8���ʾ<����ou���@�<�U��6�5l<}�n-���G@��{�8����A��?z��<��b�_n�ro�~��&O1�}�8��;�w]�:�8�+�`xɇf��Z9����֡��'Ȉ�]�>��}������ܔ��HIαl�1�F��N�|s�3�������GL�MN|yI�u-�oyr�j����}�LPy5�{w��'Y����j�Hnӱ����\���Q����QK�3���n�'5-�=�,;N��~߮���a��7�ܼ�g��g����{�ͥN�,����v@�[�oYyd 2�����i�,���.e,r����ʷ�����D���=�G3�}����iȢ�q5k�JǺ��*���W���`
�š�a��f������0r������@-Ү��2���^�ܘ틳W��5���5s�A3[샇4�X��C�8Wfu9��1IuL�=�＼�Ѭ
�4�lwI9>L�����X�Zig-�K4v�8f�ؽ`iM����q'����C��[9v��~�{�o��ӑ	U�{�{C�7z��J�lyrzw�
�ܧ���w>�~j�7K���a��4Jv�{7���F]+�f�쿐�Y���S���eԬ��i���5`��M�[a���yd�|��w��[x�~�>	�~���/���#o�)��g���ᩐ�����v1���4/LJG�vG�i?m�a�H�
�{��������:@\S#�zǏ*���>�̛��2�I�g�m��Җ#�CY��&z��N��k��Sw��|	N>>R�Ӟ���ʽ��0�h�8�}���v�����.����;��/5��K����;~��ߐz����>�rDf,�,۽���m�{ƃ�Y�C�o�þ.��3��1���dBu���Ou
x{&}_�`/�����o�[��2�e�^z9*�
��.]\�e��L�y��X�2#����_��=�d'�g�A�(¾�hN���9�<������f���a��|V*^���~���2]�)/�Y19�^�	od���5�*2��2��#yH��}{�^�RO<Ow�����������T���[�%�Gk���;�s�,L�D�h�t#�|H��ݦy���C���vf��7=�s���/��7���2�Q&k�f����{��o�n���Ž _L[@:7	��;��%��<�v��V{{�Ȏ���^;؋�2���jχjd����0)�Ɋ \1��x��-�}�ݯ�p�z���w�Z;�o?fyy�z�����Ez���=�5��E��j6?f��5�"U�� �+��a���:�O���O2�N�f0�f'j�faC�4��zp�lM^5n�Ŝ�
��@�Z$�Ƿ�	�M#d�Y��O�{���O9܆(5%�7�T�w뉢u���	ِ��6�!��%B��狱���|&§	��݇ڔ�܏�����xq����)zLh�Nۤ6��0���k��F��ͻ�H"VS�����U�~vK�`�n)��c����z��^t��ۼ�w�Xg��DK �e��(��+�n��?%�j�Q,�ژ��(�/J��������������Zm��}7,�y��=�HN��\i˒Iv��j�I����凗n� f�����>}{(͞�P�eCu8�n{�/���m�1X�_<�Gpw��y��^�/���ԟ��s��2�;6�k�"gIV��2�H���Ƀ����Fv��8y��k[��0s���=]x-?o|�ťՌ��bG>`A���^����yz�ҳ�FN܉�w�G���9]ˆl���>���7�����C��$$q�8�c��������y\
�p�x��y�w϶4�A�����K��ݍ�]�w/%�P����=���ęޑ6�����D�tx"_�S<����}ܴg,)�{쬾œί-W,z����{}U���Wq�7�3�{lOr�Mx1�p���U��I��X���y^�XT�÷���qyn�7����wX��+v!ˋ=������vL��z2xj�ίo��Gc�Q��Q��u�(�yt�zSy���'��9� �oy��cK.If��Hٛ4z�!%�}�Ú\=����,�](c���;�h�z��rZ����+��x�o_�=��{"�5�Y���6m��nN�y2�'s���a
$p���`Sk� .'�g�n}yh����z�6h�xw��x:.J��^ r9��k��f���CN�~>���k����▍� a���Gx�斑TKw_H�[�+B�v��DQ0��	�;�|�_4��'Rfumg_��F?x�9�w��J�h;��3�W����}�b����N���!7���kt�#5%�԰`:���_nUw{�h�7��}5b�B��ޒ�r۫܏�$sO���<����%���ԉ,��#�f��y,�}�s���!j���g��_�3�������-馷�g���
i��C����U���=���ܹv�*�I�Go��.)�������cT^3���V'$	
�c;�%�d��W�}�>����&p�f�	y��pۚs|�yxP����W����֖�e�"�U�{Μ�s|r/w�Ӡ�U��y��Y���x����Ar��ٞ�,i�������\�������R�^�ҵ����㪁�ğu�������aI�s`�G޺=�;_��8ob�1����?u�D�ÃO<��{w����xf��6|1k����f�5�B՞c~�6O�w�[�2͓Y�Wd�Y��Ǉ���6iȦ�ئ��\4K�j�O� �g�4�2�D���<7����4&9k�76���~qN�y��9>2x�?^�4?K���{NjI{s�;/����܁a���;�g�7�F�zG�n�����3֜�ڃu� v]���\y�c�F����7�I�`��p�x�/��2��u[6U�ū|;B��N���^�"Ϳ<>a�V�Ϧ�A�{���tqgZ{ݳQ|r�D�|�{��=C�9������|�J�8יD�}�f�9�=J��3[g�zlv��s߰���/S�mQ�0����ë���o�z�9|陫I�{݇&n���W�qQ���t����z��=.-'���	��^qG΀��|���y��������}=;]X�.��Mu�o��w��^��m�j���<��՗��.w5�E�ot�����f��*4��a���k�����}�{���y����yw#.�cf*��L2��;���V)c�:�xf�~(�%"����{����w:���.��X;�.�诺3|�`����o��+{�ӦFi��䤻��x;hVO	s+�'��G�i|/���!w��?n1��_RD��=.�rn%��o����F�.\&�]�rzݹWnW��M7}��+���@Z����	�y.��5A�:$Oq�0�K9�p�[�}��zE���]Ѓ!7��<����y��'����(�a]��Fe^��Y$��W� Z�\{�5���͉m&s���
�@���K�{{{�F�����|�.��f����O�A���Y2���4x��[��{,4{�4��_û�{�s�7�=|f]�9Mz��\7�#��yFs��x��˳qK�t
x���\	���I?���w�o�����=�ʊYɟ���	=u}��'ï�#z���9��l){�E���������",�f��}�\����z����'�g�i��2��痐&�������C��j�+^����+ޜ��k�)s�g�S�{w�{ݴ��1�����y{��j�8���X�7<�a���)��%��x9�zv�r����q��g�����
�w�����a��j�c#��o�;D��8L���/@yW�2-���z�7�B.r�\��t�wk,`��fˑh�9�۝�;�ޙs��y����mU�胗2fA��I�8E�l��J���H��>�|{ �4yZ�[�w%�Y=b�h�6��ܙ���	�����-k�{S�<����Om�gy���u� a�g����^�N>O�e��9/�!�=�>�,��K��7-�J�b��o�'��`��B}�;���{S�t�>C����? >��e��֙��Լ��X���Kٶs�7���6�Hg���w�`^��{x�o65�eP����o��$s�*���B�op� ^��Mzw=3��}A� ��J�V=���;xGs�B�91g�
'gBk�X5�(�;�k�3Gb�pG�Wo�y�9�Oc��"��Bx$g������]fOs��C8��7{Fk�2����~^�iF�nw(�������7㳷vxD3��4f�
�ص��{h��9��[�=����\���Y�u�i����#D���yPO������j3��y��;�Z6(��
�7Ǜ�f9{0$�q}ϻ�q9���/v���"i[%8r��wd�>�����<=�=�ݡĂKڞ��� iZ*���1L�.�;_�w��gt+u���PǤK^�)l��<�q��w;��<�X	!Ϟ��.�豵�������x{^<�Mܴ�{��<�{gof����|jτ�u�@�]�w�S�==cm^ې}��w}w4q�۹�IU�6/e�,�]�v�9�������2��ɉ[~�}
�����Lm2L�6Ѻ�v��x�ͧG�����s#��c�0lǼ�Y��C.�*��p(lz�y�m�����s����R��w�6`���W�=s���/���Ofk6���g{q��yN�S�>�9��/�3�מ="��_�������Z�w�����f-:�,u��Y�u3��io5����:!��8fm�z��b���1�-�ko>��Aу�8��wV� 7����;,3�L�Χo��@pZV+���}ޜ��ޞ،�2��3�.�vs�w��w	�x��)����������X=�7P���[��4�ob8n�;ܰ-B�lk������sux`+x1�N�0]�<����ީi�oFpv����-.�`Gu���g�ql�6�����}�xnx̔h*/�)���&v��;����!�wnz�P���V7�W��q:-����:4���hޮ�|J��N�zO^��q�
<�7�|e�7WA3��k�D��f�MIfM�8M�bM�m�{�)���n��9��ta�#���?����}ӏ@�8!�ȑ832�YUdY�$S��л��9.�O�}�u^�|z�ݾ�9��ޅ�k�_Q�<D^÷s��"��4��i��0��=RpiQz,�Tl�ׅ���Vu:	Ys��U�U`@�ɡ|��(-�/8���v��0���}�G����VV>mt�^���
��/���o��1]�Z<�|��,���7�.pѐJ7�č�6<y�Q{rx��n_4zU��`L�m�R5��a�� ����m����.^����=3I��ZG������7�B�r���fz�n��<�{��ky�e;�|�WwS�'{�jx�� ��=���]���.=��N^�"��^�Ocd{�%��:�J�#+����8�Ӕ��K�4yGio��ǆŞa]�o]kF�1�y�4����|�O$����]��w�r�p_��Ö�Q�Gni�C���Ч�k�/=pz�.���w��<3��7.��e��h�~�&��3{���3ݝ*,���/�#<�����;�S޳��׀��;E�;=���7{}㍪@6m�;S���V�!�ڦ[�w=��`����V6��e��i �g=���c�@�Y�ֽ�^x��k�˾�[����37x�Owf��:I�˺c��(n���l�}�5��{'�)��p���/���ī.N>���������r0f܈\���j'�tK==��5P=��>��hZon��̃���==���ɼ-n��R��^{����V';��s�٩G)���h��Ε�v���uʜÌZO�{dU���`]"�mѣ��-!������x�E�������Oj��H������#��a%v2=�!����$�FG�v�wrk������:-K��	ܔ�z��ǡ�ݠ���_3���];Qם���݋��;.���F��#�X2�#)Z�ᢓ�o��� ���ž�fn9��yܢ�;{���Y�{�8��k?Q�`M�G|�S�ϻ϶_{�'/�5��te��RI���*�w�wB�״�]�BW��ؐ����c�)z��3��/e�Wz���^M^���e]+%�p�����Z[�>8�>���u�i�v�N�)s��wzU�w��oχ��}���Rr�L�����ׯ���p�<���f�m��k�1WN���m��C7�{G�N\[����]Ӵ'����<r�5Hf0Z��>���ܹ�*>{�钸��c�W�|p-%Q2����}6l��F�vd�V���:o�c<��z_{zD6q�jQ�v�N�0.������ۃڶ�v�܎�{����×|��l�YY��7��k��+�=Sh�DR��q��h�=Y�U��c���)��~�T����[��a��������E�(?g��������k�G�~��~���3�~�ooooo�o������������>>>>>;��s�N6�n�3 	~ym��������.���.v7/P�Q��
0�x�3�/)���6�q��R�,̤0�w-��?v��w�E�o�5m,��Vk)��Fj���m���<=M�@��s,-�z�L�0��nM�X2���+�se6�m!n㌙��-]*)����j�L8-�v!L�[T,����1��$(Ǚ�n����u��͞"�L�LCe�mi�s���aΗJm��mI�if;�<d�d�Zi\�[u�����4�+V�f�K��m�j����mQ�Ů�K�3W3-���BiPV��mk�t)2�%��/v��f�ت(�5ca\K�KKn��.�V�U���0�b�����-�t^f�sx�.Y��5��2-m��X35�Y���h����l��4t(�&Z
��\����TIe T\�*ӈbV�.�s�B�Q"7�D�6ٰ��.ܕ�K��7j$8�(顢�v�%��kt,���:
J-��H��-ok+\�Na���+t��Jf]��u[����ëxjٓe�T4SL���L��DK-\]��*A��l��-H-�M3�LV�jЉ.���mKF�r���u`�)�\��CͰJV��y.�5ѨR��۰��KZ��%�)�]�	s1�V�mh-���9�4t�n`�Bg�q�g�l���=f��f��*&eکBV��gV]m��`��/^����5���C2�WF$����`��J��6�������3, ��m��\J��q)xB�V:�%�\[`K-�-�l�A�4Õ�s�8a5����m���CX4��$ul!����-�V�������]FXެq.5�Z�-	K��<�0Q����[L��ɳA�(ѤR��0u�9�DdmҴ(0�osm��`0՛XڨTz�.��\�e��m�hl���$.��iMjE��uQ������[���1nep9�ʵ�٬\0��cI�����m[��Is("b](�3P�ˬZ����.+��Z8nV�K�j퓐eB�V�6�ң����v����L�Z�hHš�Хi���l=k���YFY����XFAl!����s٩nژŭes��`Kelx#@��z��*;�َ[t˥��$(IE� !���lJ�E��6΍&%֤��N��3�4�;]6��VQ�eH�r\��bL��5+0����1�Cf@.�nb��)�A(
B�0��`����,b6��-���B�Zg���άՖDE�b�[\Ef��ŻAܛ,M�f��XD��k+[Nd,�&���ɛie�`���f-�8	�1ͬ,,���fQ���&�oa2HSB˱����)W[na��uqCl@V��et[�(Q�"vSC\��e�:9�4��3b˴bf�
b�2j1�g0�W��J����ؔ���Gf3Z���!c�.���)p�q-�l�T�8K[�x%�ڍ�[�fŨً*��X��y,T�٠W���FU�#HR͇ll1a�c���Q4k�a,&ܩxM�s
GYPj`�l����P��,�,b���IB�5`��un�j�%�F�6\m)C96Э��͇QD�250n�k����LL�fZ�F�s���iV�en@u�����l�9Ub���Rfc��j�q"���m���\[���ic�PZ���t5��q�l��8͗&�2¦cW&t͚ K�q�����Ŗh,�tM-T3Ax�yF�hT����em��33yIt(�+�lE�G�f(�l�"��B�1��nf5tl�������ج�#(�:�P����9��3��q�JF\V]���U�cRIa���tc��օ�7c�c������݂�u,#Nq�,�Յ�m��[�J����&ɮr
��XC�#�S�X�^l���eK*4��@�an����i��;:� �4Z�a����S�i�hb�5��D�p�����3J���qMm E��l�+D�f��i�[���]e%�h�$��V�u�Q6�iP@�bmyvf!pi�h�`�M��k]�%y��	v�lu,\��L��\M(���Ŏ���6�.��n�eøKܙG�́i���p�L��fM3�ˡ��5��Y`�LWcnҭ�A�FUISj�˵��rF��\f7F:���\���X�v�]�,M67���q�t�,�ny��m֡#f�TsTo6���l�Fg"�o6k*�´Ic1b�����B��B���2��1y�:�4r�6q���.B�����ێaX0K)�\�:�U�+�ܑ�c@���ՄUҶ�6#�s-�*�LV�l��e	M���b�Ͳf�b:�@�jm��.�F-�J�d��9L2�;�]���+x2�32V�ԛE���`t���t��Y���D��혜q�!�
h��ٶ��R�t�n�ׅ̦��ncCB������5�F8�d�N%�M�*nԁ�������W]cu�#�X��f����6�Kn�Qti���kqB�Va������\7RY��V�<�`��u��nf)��Q�ڐ�X2��jf���f�5�:k\d�f�UF]2)&]+ZG%��$5�R5Gf�cQX►a����1&t8�l�U��-�.Pe��6���X��@D,�.�3�kE,���Ƃ���Ye�7��0�6[؉mA����R�Ќ�KUqƱ�]�-)����f��vR�JktB����M�2�	f�.�
���ai)��k�KMkKy�{6����պU���-�M���t�Fm�@��$�]P�v�Ua��U*�,sZWHe��c2J۝3BRT*ޱc�
۰�%��4�i��#^[Aŏ]f��iɜ$5�hh��m �+l5��b�3�fi�\�p͌4�-.t�чW-dK-��a�����*C`63�ڰB���+�0�k0a��ff.��LL\PA�5�1t!�		�u�a��R�c8�Ef4)-50k�m%]b]��K�S`��!X�ilN;L�� [��i@��3\k4;J�mΑt4f0)�n���u�]rhˆe��a�f�;XX7FX���e�f.�D��Xsk��)H��-���9,48�l�X��X�aj]�6�]��jMd��t,���dIx�0�a�����f�b�;GCi��,�G$&6#-3V�̹��y�U�C �P��6.٢�][-u��t�RZь����۪%F��M�Dٮ�T��\k[d&e��˖f��@jg�n+��`���v��%3�AsHUl5��e3][B&f,HE���eY�	�V6��Ɍ�Y��7hD�v��t����13�f֡J��Z[��:�A�R$6�m�/Wh�Y�Q�Y��us�L��n@��+4��)k[˱���Z$t�J.l��β�u�P7�eұ3s3q�̮�L�c��f��	]�kz���t��ŮWP1�-��u�u�z�ђ�5�,ALH3t�j�3Q�ĉ[`И�(I�\��pp���#���V�Q�وhb6eH�!�C�Żcit�-2�Q(�KMQ��k�P��k��R�+l�K�tqs[+�.	eSpL�Б�#Si���R���Y酘X�5f���nlG�K��VVy���)��m��:�����r����m�2��k٪�W)nn,D1�kcf�р�����!l�6-�� �(n��%t�T1�R�H�6^;�0���T]�v�;0���MBi[2R�h  WJid٨�c$ј��VfKKam�Q35F��ͺ\�� `��
:��B`K�,�B���"��Xj�Y�6V��0r��ֺ�,.4"���$��e�a��%٧6��a�Ů�Ἆ��E��`�(�;7h�f�� ��L�r�.8�Kn!�0�l+kqli*D����,��c\&�)�������,+e��P#��f+r��+�ٕZ�)4�,J��Nѷ.p�Hms�K�5,W:�X�Բ�mY�Re��"blT��ͅ���*�75Eڠ��(K�K��ع)6�!(�Ѳ�+K�Q�u�sb;!��F��B���jK��]���V2���R��+�D�m��r�e��^��ni�-���j���0��gb]��X�*i�v`�+ٱ�d.K[f�Wj�LK��ښ�kX��oD��ЎkF�: Z�,�ۋ�ZR͔��3�V֕1���k/6��+4n�ЋF��t
�k(
݂]U�T��Z�pd�0P�j�S7R�fQ�WJ�q�����x��:�L�zl�ǂa�Te��.Fۆ�j��C`�n���D�ȵ�B�XBT��`dʪb\:gV3v��6[�UuY����+U�i���#NkM.��%�*ڹ�L��뙸ҩ�3����vm�]���-�+�Me�3��q�G�6��m��7\�`��Ċ���̰�fPtu(5m�ЄɖX��ٗZUL����ؚ��$vĦ�E f�lmWYkvˮ�#�Եbr�h�� 1X�u�K2�aH����a�/�JF�1�[�kX�B��D����5�
ˌ3�55L�v;lʶ��U�3c-3�8ոYU�-@k����4��i3kP%͍��b�c���17�l�%.��.�E��v�mtV�L�f���#���e�Gm�[��:�ebŅw,I�Y��M�ڮm��E,�V�LJ��R���&�Dҍ)����!�G�U��E�6ںŘPQ�,f�j5�]r8�F��E8f���[4��f�Es+J�ں�4[�E4�Ff̠)�e�l��A��榵b�s/���X�,��XOm��o�lk	K&�(h`��qvH{4��Jd~fu�W�.�IX�Z[�%��Lŷ��E�$u�^Qk��(t�
h�����0�����(8�$keD��M*p�G� hms%شكj�*XB��Q����(��ST�[jG~z���b�njf.,s�wB:Z4C��[Fg�g��L�(KAn�ex���٧��X5�W��^w4�i�>�-����i�f��۶n#'����c�5�>�"I�a��fݍN2�F��b�Ӓ���RXi#-8m�m� ��kl��S�ِu�f�ad���&5�p��n�6i���{f��	8;���e�;n�jRem�ݶ��0���E�R"@ ��Βt5�M;3q8D������͍�N�Ne��in��me���G9�G*{dD����pq��Y�w��dڊ8��f�n�ݐ�!�f���M��ݠm�A�J6�$��,R.p��՛c�䍵�wd��Yb͖H]�BI��i�O��j;+:�p��'!���vڈK2䓉�Yf�6쓄���8�(8�i���83��:Ӻ8���Y�slh�~���8������X��%����y��۫8k���.�H�C
����q�#�s-��n���iv�f(ؒ��m���F��\r��e���a�5�F-ٗl�b��)e��5e��B�f���Qmqe��� ���ٺ:��0�.�WLL��0"�V)���-Ś�`L�,�h�.���������@�w4�����&6-�Ve,	f�������X�Rîe�Sa���J�9���a"�aʱe�H86���U��e$ˢ1��&%�rMvp���^%����)�����Z��]Mb��j!K5��4RY],ՙI�_!K�xL�V�jʖan��B
k`��՗H(�*��]iIur�Ac���V�+s��Zp�56�ۘ
BS
�ٚ�ƶ�Q� �Yvѓ,CWmqX�˶]���키����4	D�K��t�E�ܤmEε�GM���t��f`�*�"�.��V��J��Ut\[t�	IK�5�mL���(�a��n�7+lJ�W�ɥ��f�k1բ����L�:k���U�<%!h���1nJ��PMŬ8��*�jK,�fB6��3]uEb6���ʁ]���B�&��&�Ri[�sV��;����%�1�l&�32�+�D�g��88�ң����S\�5���h%44�� Ĕd�L�cGm�W!۩2ŷJ-(-+%�v�B�.�-jUMv�
˨k�3n64�E[+rF�H�h�#���	�,º�:e�&�f��5������c˝T�,H��f��#j0n��[M
X�Y5Ef$&��l�C�Mn��	J��:T�	(��:)�����M���LQ��]�3��T^*٘����3��4 ͣbg���S&p�y�x���îЉ�X�k\�4D�g�,�!��e����a��2�Z�\��$ٙ��Ø*a�JKԾ2���L�qb�uìǄ�P��b�.P2������N��XK7L�@򱶖� -d���������H���Ҁ�V�F��ƨ���	mh2�@����)[V�@V1�ڶ),j�����Y[Z��PIW�m	XJ-��i�FW���e�6E�5�1UI�YXն!`$���,H�`"V^T�����akV�j���mE)e[el؊�
�6	��?��?&B�bY�E���V^D�@�|��G��3(��d-\C@��`���?{8��#��^$e����
�6��_�T
5���H$��Nd�-�q �s��� +}��{�A�;�	�b8�x0A�y>x6�?��ci�K%is�9ob�@+3c��n<�`��wr���[4�$Td��ǡG��NDI ,��$����S1�T��}ѡ@�(���lP�A��H�w��Ao� ��wz���y��l݁s_^<gLV6i�D`��X���>(�L�ŝ���)a���X��Jt3j�v�nÜ�N���H?i��I�Afہ�l{x�&��͍x'v��k�]�K��F�Dx��� ��4�,�`����|3�ԫ�=y�$N��;��wF����:7��x�ʲ��Lw��M�����՝ޣ��r(����uSߵ�n��6���RjwH8	纋��B��O���q~�t��Y̾=mm&��A��i��d@�H�5�8I g/�p|�j�냴�x����-�{mp�"|e�^R�bY�41i�	���lG���c �sI��q��u��>���v��@ܲ;;�vwQ ��xUn��j�����f>���U�g��3n�'R�a��{{�&�L�xK��( �R]�H�w	�%a�c6Bi�Hm�:�����/�L�N�#L���1��$����Cy2d̈́H'�Z���6��������h	n�RW���7���6J ��A��x$�M��.��^곥
��6O������k߉�>+o"'��}b/X#Kn̰��w�P2"�ZY����*����c�W~��ٻ��i-�kLoI�Isa����(�K����.BJvJ��P���>Љ��@+wc�{��` %�_��j �湟D�E׉"�m�	>Wx�	'[^�(���_���W0~G�	%�`A�@�𿝀A�M�����ʭn�4��R�H$����:��`o�ͤ#t�я��F�A��M�s+m�f��Ci�P5֤��E�Ys���]��k.]� |�>mf�F*����磝'Đw A�'u��B��U�B����Լ�NO���I�S� AZM�0�Ō�Amc�~k��N-N�$@f�i�[���f4zk����PZ�b?�Ӌ��#ɒ�&���4*��_��ĝ�l0H-4��j��[v��{q`�9� �H�w��/�%A�%��Djj�U��dV՟5N3�@&q����}E����g&w%S�=�g��M�T�Sz��@��q�8���Z���m7��vw���)�eS���2���uf���H6)� AY�S+rX�d��S'Z�H�|y��Dhkh�\؃�O�*7�>![���$�澽����O�(���-jfme��D�fee4iF��J�P�Y���4��T�+p�e��>_�����,�ݑ��F� �Mm��$�׏��ǧǺ�or\@&���}�lF3 �;���� ��x$���!�w`��NC�����I"V�l���{:�b4���)�"���
�l�"}���$��2�{Ԙ6��$mm0O���A���
��d���B�i���S�E�E�Ԓ<Z�� D��x޽��	�[�ml�J��K@��D�0��0`İp� ۾<�|V�@��idnSQ��w� �:���If�z �a�5��q��gF�s�������bi�"ݭ�d�q3B'*�ᮆ[+l��W�����7�(Ⱦ&���{�ѓS�~2o�G�uΫ�g��x$�Na�>m��
�	d(m�Հ�.�Ṟ�H�ŉ1-�.Pw-���kB�Z5�0�[��	�EJA5HZ����e�5�ݚGB�fa,^݁.�v˭A�]ОI�R�����RPE%�ņ�3\ˌ화f`!��m��.�B˦�����٩V؅I���hZ҈�X�l\��C	\��(ّ�7V͐c҄�$̥�a�SiU�j��*��r�f1M+.���iXŢ��cuM�l�Մ�u����[��nؖI��I�\�%�'b��k�G��$^�?����D����;�=6�����?�;��	%X��m�/�fI�ܷ̼U��ں�}J"Z��|O�D�;�|�vy6��;VB&�l��c�ؚ#F��̃�;��L�O�AU���|N^<l�({:���P��fLjj�6O�7o��V�Dm
	�S"�)��ѭ�;~)þ4��jׂH1��[TH'���`�j��F_h:a���x�����a+4��R��/z@�������w�형��ȷ�`��}>�>{��𕿯�J|�z���,#�K���lk�F�.�vX�X̨�A&�fP��뫃K`����{�0^`��#N�ۈ��� �_]��F�AƴD��׀I
s A��	�ؖ.��
d�h0�K볢��zkS��}��ǋ�3(��Թ�F��G����'`���ܘ&o���t�͎���җ�<�?bxu3�b�g<f)��`S<��$����#���_x����6VI��3�[���XK34��;�>�h�^(Z���ck-��>fL$�o'Ă�6 �[[n2A�3���d��q�$�5��z�m5�� ��>�@�{���W �x�U
�B�fD�w��� �ֽx#f5Y����~�$�l|;�$�Sn���X�#I��8���)�3�N�ܳ.4�73f�1��-��=�h�t�3M��K�Y���[��]vf��gAY�p�>$�m׃�9K3ۛ	4��ŵ��^�:�`�r��P`����Dx�>�Ii܁I�-�(kAs�V@�$���|�H1�^	��4uz��fo�)}�R�� �U�i��>��x$�@^7r�x"�H/�3O�q�LOO|���Vx�߿%���o�"�ek�<���I5oh�f�|[	�/�K�K�ꗛ��V��0���N�sؑZ��i	��حZ�6�uy�f>�� �cD �����[�$VmΫ�vK>��I�v� ��P��Ŝ8fw1 ��q��q2��
t���>� �	��q��r=v���Y�s�ɘ�fgB.���j��f�քj���3]��sK�Y�y��|�z�ƴ�q��Eّ)�?�<Լ AkV<�r#�D�hj��S��<I&Z��FQS[gCi+p%��`��^?��W�|��� �����	'�QHJ6&u�P0nl���D0`�H(j1�Ē
���/n�4�L?�N6c�'�-�wx�59!��]�L"�ۆ���A�l�B�vVm �i�IWwg�_[���s�+�z���F�C��ID}OO*�]��C�CV�k���,�s' ��
'H��}ءv����t�0�Ѿ���A>na�Z�XfM.AN���@"u��i���6a�l3}�C;�����$�g���~r�S8��Y{��6u�a�V6#q���6Md,���nq��u3'�=�|�ބ��e�~|�n�W�/čm|0D4S(�K����	���!�2 �,����������04Xu%�7C�w�|J�ȂI�����OO9������7���ac$�����"�[!㌓��S��"�w��� �j�p��$�k�H��KP$ ?��?k��9��ޯ6���-��e���5�>몦ܘ�1��CAo_L�>�|\��C����jL#0 -�{R���
g5�����kSفJRcu������A����o�!MC���[�=&^��/��c[�����B�2B�V[Q����G��݁�� F$���7����o!�e����s1�@����иJ�l�k�lEU�J^n�8&�,!Qh�e5U�.R�B]+ VQ��M6���h�3t���R�I-�6�7��h�P<#�pj�F�����K1�k��(T� ���-�Y�A�6iW7]3�I{L�ױBȺ����ڸV��p���m���kCvƈ���t9���J,��~�=�ϗ⸺lbe�eɳn��cBd@]X�[m�Wr�0�I�����
�i��l*��|>~��� I���~P ۮ�ӵ�z���޾D�6����
lZ��`���ߧ�.��ئ�[�xߨ+�i1��"_u���O�y�E������}�e\D�$���|l��Pk^��A�:ϔ�Aw��w0�	Ʒ� �m׃�(R�`Ν�)4� K�K��'�'H�C �^�p�-|ǒNy&��׳
񭏱e��� �Q	S����x�>��H�دLj;3T�A$k^��	n�]L����jC̓�1��
�nP��Z��aXC7	.�0�V�JԺ���w��e	���|��6~DI�-�A ��n2 �Y�j�M�A�o�����]�)݋��y� �y�/,m�cE&�b7�K��N)��za���4v�d�j|����}F�ZX+.�X6�k�ݗ���V�
Ӊ��"�&�2աA&Z���O�m܁ �S�k���|0ۛ(6؝�����E�r �h��F���I�I4ծ 
���C�JL$��\&	;�&$��c�=+����x� �O�2 G���×:�hѺ1��Dc�<@��X3����J}B^�~^\?S���X���}x�� �j܈']��9����&���Ǜ��޷h݃:m�j�1�iqsIQ�1�J��)le�Q�6��M��}�~~��)�B��y5��O��ȂF�v�
9z}�����A�ּ ��0K� �`a#6!D�kh�"]��ӻ�i���5x�o�t� �x�%�*�)�_Xn��;�S�d2|�<��I�v�<@���>���8�����������:t�����_�{=��g�����%&]��w���ü�M~�o(k[�Q��#�d=�7�,�����1��<@��ֺ��y=��w%x7U�Q�GI�w�<�s/[��>��;C���;�{�{�B	���(]efY�ܙ۞��{H��s�������P|g�8���K�N^}=�k�s�=��Ë��$���2o�C޵��݈$M�v�RON:�����3ހ<;z�7�n-��)v��aB�
���6���+Y:�$7������z�"���8{}ȏM�q�X�G��N�fU}�cq�йf�h�A�p	M�nk��w�O�;���M�-;�����F�
�|��TS�l82���Ji)��z�ma@����޽������8�aG��>���{�7�0(=�ḉ�������ٸz�;�M[���_��K�4�j
��[�;���}�$�]܂b��<��>���1�S>x���k}����2���g���Cݘ�;���Yg�'���w�Қ;u �����ޞ�^MЮ�
Gh=�2�e���qs���н*w��펴sԭL�)����.5�����z��i�-cݮ���۷ݾ>-����;���?x�5�x3޺��6;5iw� 9�<Y�Iqj�<�����N��} �:oi�>���r}��5���=����/|���@^�t�<�˛�=׺u�q�l��r�}��S#��g<eX�3W(Ea��v���]$F?/_u�| 7�O��'�U�D�P%��^�X�jW�;(�N�[��WY�U��!�J4��}G1��m��~O�tsS��**L�ΊkNf Nۻ8��:�i�[k;��s1���w[��%�F[V��-cwi�-e��t";j��Q�YII����N��6�n����N$�Xrm���m�[n��@qE��%ip���fGgf5�*N��2�ge�����D���H��N#$ӑ�
;.����lwf]�B-�#���ݘ] �$�#me��3����tA-2YvM��;0��2�-n�tBrw�1�Іۢ"Fkl'�k��D�e��o=e�m��{ݦv���7'<��2��[k8�)�Ar�q�h�Yi����m�y�מ���٬�t���{[׬�-7���۴�Ӽ�v�7{׭��p��V�E��ye綈�=���y�{;�%�i�zD�2�;vڝBi{m;�� ��|��=�O�d&6Jfa������)\���>��1��|2� �ӻ����D ��܏DŃ͖�}d �����[��̥&C�g�qǜ�C�HDy G�G˻���*Н#+����Ϡ�R��N��5��$s	��q��z	�˥��ïޡ�����Ξ��tx/����sx"�+�����!���������'�}�mGJPrK�a!������@w��<������= ^�,��U�-�8g���ub��SK[����驃9[������S6�6ۃC�>ɑ��r�̸A��I�q��Hr�Hdd&�}�xN����i��tC����)J�L�u��9�dg:�,�,3l�9sNe�� 3�=�{��O]�ـ��lc��އuig��kD?�zH�v��mI�����&C��J�>\��}� " Gȁꬋ�~�$�x�G�"H�%c��D8v!D��@������9����S�/=����d&F'��G;g[��^x��!��I�o� � �\�!�}�}���|2�Z��)݋���}�H�言}�͈Y}���	=��ޠ@G�D|'{8y��0���23�<�xN$�"�L3���y�7�oMxq^�5����l\h������W/���Ҏ��_��l5L�153806x;�ϤOj��u�[9�������}���O @���G��A�"����	vwb��|�N�������x����	r�_�}� xL�Y-M�����=��2�k̀���3Z�q���v���O�����ұ�e�V��͆�*i�K����e6��]i���Om����f� �z�Rm�w��Os��;�[oq	�0�B�"�?,��$H>�����5;Gz�����rR�}�ݸ�����~Ow��L�sv�����Ӣ"#��$�yx	WKQ��{��u'�s�\=��!�d&=���JP�Y)������rs�VBd�w!��{�ǰj܁�D� �Y�T�	�c�9C!3Z�y��� �r6����xI��>�y�gP��6�5��^C�&C�d�O~���JR!���	"H�Cj��Z����P*ϼ	�lw� bo���}�O�Bm�{oq	�Bdd�Fm���1� �� ��#���y{Y�,�z��z��0���xw@����o�k�Q
�v�F��2:�n���ːd�A�s��zA���ƪu���g�O�Dxw߻o	Ő�6I0�a��kty�� �P s�t#�@��خ��xǛ���.�]p���_���]����� O`���ā}Ow���>Bߑx�u�G�E�vp�Y7������9�i�t��|?��s��u�)�L��[�[n�fJ��m&�B� ]	s�c��(��*�RX�� �B���(4���t%����tv����՚��Fl�kͭ���f���K�L�3��u�nΙ�6��ōc�\�l�1��bWhpJ�dV饔��j@{h�cX0Ά�R-+���h��,�T�
ٮ�ZL�;p�Ԏ�8y�atcVԕu-	u���/˔�8F�r�_mA��xm��a�2��f������L�Ļ%#��0Qa�����4��\Uo���?�Iw���$��I)%e�ۿu��/0a.JRy�����<��~>���
���}��f�Ϟ2N�؝�0�#}��p9�a:��f��!ظLg�d�
�~��|����l�D�������L������=�Nc�����:�\{��˄}�}�ʝ״�q�'9��������N�'�����t�P�7o(~N�'~Ì����ә9���2��=���kv 7�c�!4s����r��n��Ȟ�	ݒ��oߜ�'/�[)[�&l�t	b+��"�	V��0�)��� *~w#ܶ�\Z�o���8 2�o�n�/0c.I�&{��{��<ɐ�&BZ�����:7����������8��rC##�5��s�g=w���PH�r�+�Y��>�����^�I����M(>坘m���g�23^{��z��� 2Mq���re�2^�6!�{�}�� 3:߸�|�������Fݱ
&lZ���]vjQ���遌9��d�\�����b��R��]l�}���F��L���[�$�˄.,r��q��i���2M�3��rx�Qc��-�!�ۮ��,$"��'<ൄ&XA�|{Ϝ��ԆFwߚ�?t�W;[��߄�%$���N� ��>ouUwF��Sh]���1N�%������[����nw�����ۉ���hv����o��%�pol�l�A������<$�͇��Ix����rL:��=�rd�p�%�s�}�s�@ #�@�F��7˧oΈ"���ဉ#�XȔd��8Lg�>�|6����)B^����R�y!�y���3�������$_��GȀ�#�`{ �\�	�h6!�{����I��Z����)3�h=g��~� ��k���׽���K�ߜ��,�)Hdd&מq�'vBrY)�a����{5������<@��q�<����	T��0�(��� .}w/9�a.F����̼���[{�[V�{�^�ix�!�:����r��L�';�����2�؝�0����mO��>h��!�6�2d�HHb���6u4.%+*�1p�A̽R� �rL�Q��
D���;�w,��#À(�7c�xI�S3��Z�yJ��J0��z4�
"��Dz&����l������� �\�#�M���}o��0���y�V+�]A�ɧS���^BϞ��@��'�DG�W:��̍UYS�A�ܧ���I���������8,���Ls��mHq)\�dn�d��F*|��`yg�"����'glUo����Iw��D�	%:�II,�r6�ݽ�Yy�����]e��i	��x��M%�$�7Ӓ񞭀�ER���C�`��Mvx
���w>�_\���<fl�������Z�Ӛ���`��tPwd]�����}�9�&C�d�Nk�o��A�9)F�j^H�h��d�8Lg�#�AGê_�y�2��{6��I$Zy�ВI$��je"u���c�_-(4miw��/h,�n�D$:pb�-�8p�:f�wiD4t��$�Y��.#�����G���Kz�$c���*�W�^��D�B�SN��
$:�쭣�Z�� b�Dr���k���� �W1f��_�v�|���iF{ó����@�(�fKI$�Kt)H��nZ�P#�i.�h��Kɀ��Pd	�<N1w	yܲ
��>�����Hm�ً>h׋=�$$�
rՊg� ���RA+��f�l�j5̡���"e�`ɩ˔��vPI�i�i��M�B$ʟ0' k�����N��>F?��@������$�9�-�&vgLS��J�g�7=����lZ�}�A$�cM�iI/��J�$�'��Ǐ��2��I<����6�}t��S�v�`FI����y���M��j��Y�V.�;�U1��(/����[!��Y2�4�����x�t��o��p3IQ!8p�$Π�]��ƙ�I G��r}�U9�z�jǻIx��w�Ox�B3H]��Iy$�w4z�sL��qؾ��ߴ�GB�b4�4�Ԍusvuk]ku�5(�*�%+
4Vy�'��g�*ks]��eO�!���2A-�i��H$�����45�3���ݸ
e�ԁ(����RB�A*�LQL#�T�ϭ�H����N\��T�۷��'�"ޫ��R�	ݯ瀑I ld�ݾ&:l��7Q�QXFaM�q�!�w���_R@-�}��: ��EOi����s� ���S�I-�h�%y�!�&�.S���R'��O��8Zg+���H$ֵĲ$�۬��H��2"2@fY��t�ʐ����Չ&�(����|���}	$��ϥI���X(�)���	.;1�T��@%y��PH����?��D6����O��[�|��2��׊T�^mX����W\�;p'ݐN�v�M�x�ވ�9G�w�iнW��YS1%�߈ >���f%�&vL��b�B1sq-n�lk��#�Yz£t���4�4�v .Sr�B92f:��䩍a6��7m���u�e%`���E�:s)����jc)3��&e��mr5�f��;��g�,MY��!�\K�)�hZ�60��:s60���F`��]xPn��s�fКYDb��[[M���]��6�.�FF˳m�����X.v3�F �1A�mWP23k���RXA�*f�7�g3@v/�{��?��M��������{�o��	 �oq��$�;3%nӗ^]�헙D�I�1�B~,�b�Ν�h$Ϗ����&)��̞~k��dJ�J;��e��%�Q�	$��[yό��ډ��+1E0�)S�y�
E��2ZI^H��r�g����V$J�W��I0���L��#p�����U^\�� F놼7��HݰI�h�$@$��ݠ&|�I{�_�f]�ne]�}��!��>��>��K\��
r�b�PH��n�K+�7Y9�RI=�D��J����)$7e�T�|h��w�:�痗�fnKp���d�&20��f�z�Kt`Z�ai<.��c֡����]]Zm�g}����B$�v͟�>E!�/ҥ#뎬f/�7e{6��˴�$ӵ���
�Jp�0I���~���y/x�<�۳�,�KB���{4�{����{;ⵁ}�f�_�����׾^�\O�hg����ʚ��2�P�s��)�D���������>�Y�g?$��Z����$J�}/��	 �̽[P�ֱ���s""��"ػ�D��hd�����b|Ȕ�eɰ�©.L�i z����!.�l�Mt�L�&H��
��v��#�^.d�J���O�I!�oҥ$^K{Y�4�;�y��(�Np�*})Ea����p�*�[�Z��"I=���G؛���hh��(�$��5�TϒI,�~�)$�[����/Uv�8��d�d��39�326��W\�g��/0��,Ť���jV�$��N`����N�ӕ˒�j�$��9��	 ���;�� %\�W<�l�Z�|�2�*�%O�|������)�ԉ����GЦk�'1���~�d�C�_e!$�^�B(k0)�E�ngS.�t�җ�*AIÆ`�<���m�I$W���J^	G���SA�(����4s�:DTT���EU�Ǔ��$�� �?E�{�9?W�%����M�aϙi9P���j)�&�'��fSE�_��
�B4���H$��q�w�8�0d��>�$�.�Y�~��ΉgN�D�l���v�羶�&�T���H$�U��>I�\u�۾i��	+��EҠ�ءl�L�L�=-^�O���I"y�2ZO�E�-%l?N@��$�-�T��H%�����@����{��1��MT���.�h�������M-`�4�hM�j���u���Ͽc���B��l4�&��a"T��)���C>��L�����I$�^�xBY��Mn\�`�ʕ)u�L������j'a Е��n�dI0�9�Ą�IO�byU-�`L]��,�%�X�^��0L�S��n_��>LE�H�k�늀 ��kN�uX�.4�w)IR9�����󏔏JC�d�!$�ðI��st�Vp�7M�	Y��I )ڹD� �Ids��<}~e�pm��L���8�gqݭ�x��;ǰ����Ρ奮�h�6)�W����gw!ō�ݶ�[:�[��bL��=僸CN�س�G�P�)QB���%��$�߈����t�UI3��!�$��5�%���ֶ�+-5��y$�����K�S�ڂd$���I'�.��#� �������;��aƻh9n.�hG���e<��e��a�6�ˮ�ov��'�E��W$ٯ�$��	k�d��@$�;�L���h
'�M�7k@�PI���D�S�_wrW�� ��,藿Ux2$�Z�udŷ�ܶ	D��;�)��L��~� �I����Z��V����l�����>7S3���}y� o=�u� �@���،c�y��H"��;�)�I��)'��L;��vuB�&�g�i-�N�X��:�+�0��IH�+ѝ�F�K�/%]������# U<��I��Q/V�R�����Ç`�<�0��i/$���ֈGٝ��Тj�a��R%�ȓ)�K{�![��=�oW������g�����ח���:t��ۡӯ�}������+tߢ��*�,c��L�fL����>f���jK��V1<(ܠի#}���v����ӧ"���-�U�w{z�%�f$Ril �Q�s���9�^�FU��O!P/�����;����ww�L��e��=/bX`,�)���zgE�`回��ɀz��6?m{�EI-����݋=-���6�z��r�Ŕ?����=��ý�R��� ϝ��f��gj��_��c�گ ����z�aS�O��y���]6�=8bKn�3:bӃ��h�}�;5v�3���P��˾[�z ��<�,1�n�{�إ���Ѡ��w�_n����e�}t�N�}O3�	4c����wŝ�N��n�]�5���D��K80��̀��쓄�n��v��y�o�*|7��W��{V2Z��S�����(4q�d�=�Z��<=}w���:�/w������vx?�x�D��91jՃ�g��z1���f�7���S�b^5���:���y�8��*�=Qo�������%�>ދڇ�6yw��u��?o�c�r{�MJ�v�X������x_d�W�C���\H	���^�)��;�^N��oި���:�-��^Y�C�f痤�3��]�������<J`����|�X�+�k�u�;8n>��tJ�g���y�j43h���N���-^�z�唱v;�^:*�t����[�埑�q�6��2^�ڳ�_��"� G�>��j�8)ǃ�M��������}:D(Z�nyOY;�ᩧ$��h�@�BG7t���e��gӽ�QE�/�F�`C�1{Ǒ��k{'bq�{zB.������nylӞ��{�1[�f�c�<�ON<��%�J23�����
���
�K=���P�����z������<�v�����ӬO=��^��=���u�)���Ёo^%�Of�f�m��l���ٚw�ye�`T�[c�0,��� YR`^��6m���^z^����F�,�Q�$NX"�(R�(m��{��vu�����N�׽[k���y�8��R�؄ ZƒX���'+˲�휶���Iy�������n�6J�죭m��޽ݜ����On�f^��彻;<�쳼�mm�<���7���^��2�2ɛvߐ��|ɚ����{���n��y��:��(���*Tv��n����^oR���^X^nvo2w��x��4G��[�l���<���n[f��#�2���y��w��Y�Βgnֲ�r�������oZoZ��%۶�tw�b;����ҭ�ҽ�G[n��{۽�y��fܳptEyh%�zډ��f���綼�'��l�),�y����%:��g���myy��Ykn�e瓕�Gy��ۺ�'C���MtX]���5�\������Lf� �]Z�VR�	�:��4Q6(��eLiD���T�Yh1K@Ω��F����t�`΂526�˯R�n��&���͎]6r��#�)��+��1��j�#Wf]rś5��t\g ��o0�\أZi��#5��A\fEmKx@ �R�Ќz�0��[�j�kCv�3SfTh%����WF����.#Iap�N�,��l�L�&l1���ʓF"� ���NV$��+M5
.eT�Kp��Cr�Gl��W\��G1����j
Z��V��-�hE1e�b�k�QJM��c&��uQ��^�f�k
�l�d�uو��Y��#����1/X\�ǇY�X�y��D5�]L��"ULM�\�\�%��-+N)�"�^[���3T�4�٣p:=-���\F�&JM�s3Vp�)S�Z\�S�2��h�&-�ZckL�Q��u	Fa�\�	]n�mki�%]�6tX�H�v�
�˵Y���%��/e�3�(ʑ��;��ƍ"��D��:��n�5�Z�V���n[���c+6����#�#Qs��!���hM'%�.4e��h��.B�X�%e*�ڍ��:�]�L���B�U�.�v��ᙳ����^ ���Ƅ�M/h�6�� r[� RhR�PM�m�[����L����h��ufw4��E���k���B�Y�"��6��!0۱0b�uK2Rceղ�6:�L��FmV�Db3l�+�#Xd���bj�ɶ����Q�X"��n�CXM���x������<����B.1�Mq%�5[��V	0����x���3J��4(�ҙŠ���R7C,��1v*��aZT�Í͘��bT(ZV�8,כCF0�1[ �:غRҮ�΀��16�2D1pͪ�2��-#4�T�J7�a���DƳX m�s(�e�lM�Z��o���-Bۣ˦��X�8-�4�tr7k�]�����p��m���3A�� �ӭҢ��JRl���K�ZZZ�:�>�G�@( ���J ��B �V��8�<�)�W7le��5�s[��n�B$f,0K��\�ف⛛ML-ֆ
�+.�2���Y�v(9�b�.�inQs��eXp+h��j�-�&�4.�{(�l5t]N�+i0d�H[ac\���۰�q1�%�.#eb�
��;�4T\�Xa4e�\c���GȺ�J�G]KhS��i��%]Ik��)����6F˦JMk�u%�X��-pǌZn ;i\��Yv��n �l��%�(D��Mhm�\�9?����b�F8Ͻ�`���-}~iA$���Ą��%��@��֚�@)����Ӎ�;�)�U34ntI�������E��`�S$�nK��D�tuƪi����L�RҒ^Iy�2$�H$�K�Z!@�����V�R��/C;�+��UG9���Iy+]�掖d�H���R��d$�YҬ�� ��{H��ׯ?O��+6��o�=��X�qeyΘ�>����J_a$$�5��$As����A�GF��$7%�T���`�	��r�;:�T綌���Kv_��O��v����6�`����T��H%��$2 ���T� �
�73^O�~H�x�-��l�ф��Cd.��m��v4�BSG\�;]iEs/ZS��o��4�0���_;�-8	��t�� J���ϒ>�hRZi�c�S�z�Nz���������|���=O��?}��>G��������]�Q����HS�R�Z� Q7sG�Y���^ރr�P4�q֞M��`��1�7:��QOc��X�"/���p#�����R�V�(%��(Q�R�'���|o�<�ffffg�sD�?;}�e���u�{/oL�D�[_,�H�b�f��J��u��D�䆒I>�^��ّOќ��$��1�A��Q@$��~�B��g��9(9v,z=U��d��#7T��ai$<����BI ��~�2@$��Џ�n����,���.�h��52I���3p��z���JK��o����ڦ7���X��a�v`�4@I$e��̢�I�_�}�oQ����3xI�$��f����\��WcP���]i4�T�p��[P˼���Ȼ�!�'g\7��e����!�K"�eJ�D��d)}͢��B�i|�`��4E���Eʒ��8��L��v	;���n�l$��㋻e=,����ItDq�H�ٯ�~j�$>l�k�rZ7!��d(�'�����gN�D����PI$�͑,�H��������v|Y����}���߷�6�ESW��f{u�w�,��E=d��F{S�Z&��o�=b򃉈�M���\��l�~ {�� �H$*�%*H P�H� R�B�@�#@�
��<w��~�1I,{��"X�����*BH�t�f��J��ܟ��E����$�j��R�K�/g�:6�4����G���\�צ:j��lZ&	��Ӝ�X@ඝ~V�~J��������"�j��wG��M��Ȓyv��)^Ų{�ჭ�M,1>��d�G��Eƥ4ٗYX����jVm�L�ٓULY�fE41wf`�sr]��}9�D�O���D�$�5�	�b2�F�̭��q�D��j��R^x��l����vur�K�!!�f>=}�ڷ��
q]6d�=r���	5sd"O�Ov������2�\�]���x���h̄�΃XKn��B;0���������C���1�g�w�^�33�>�&BH���BC#�7�����K:P�ݟYQ|�|v�+vm���D�[lHdJ�W�K5�H����x���
�Ķ��tU@�v<a|y?���8��6y���2����w��v��a�]hL�U�ui�"�RI`��A�y��;/?��Fz���� >�

B��P�E&�J�iQ"@)B�%
E���F�'+�3~��\�'����%V0n���@��z� ���o����������KeJK�-�,} �W���r`$�����|��
���Ma:�e�D�Q(�U�4if+�l�R��ѷ�-�*ݚ[p)c�	$�c0�.ΉN��˝l�	su��I~�3 o����o�z�s�����o ^�B@_vE51wf`�YK��6�.�/bkl��/�m�:A$�����BHK1��2�H�޺X:.�"�:޼��g$3$��PI�غ��I+~~0I'��4Ew4ZR%�z�V=��H%}��%������I�
i�kMۆ���s'���z�6�.��H$_y���)��rN'�8��Q)��K�B�즪߲��n�	
/�A���.��U���B�PI�vD�0=Jp�9��ޮ��膈	$����Mz%�$满�>>>�Hx��<c"�\\��b��-jS�{PpFb�}		l�	�W�����9p�^�PLr�E@�Q���6����,���T3���/� }� Х �@	�2�B�)@�"���+!Ht� t��w��K�\ݳ��k�#Zk�1A�+c��^еfŔ��&�g7g`;DD��P�H�rj�qJIH�q^"h֒05qW���ڳM�땲��k�vR�na	Y�ܰ�B�5�6NT�ZV+��U�`n.�q�kV4MF���f.�e�u��f3�U�L�ܘ�^�P�fkk�ۜ[BͩQ���!m"�2鶁�Yv���Kf��bW�$�u����z���jY��+�p�q���2큅����X�E�4�sY�Cw��;����1��w�?��ǩ: 8�o����"\��<�|ݶ��S*�iGcD"�-t� �v�� � [D���~\���$�7�D�<ΰ��blvs@$�	y�#�ϒI1��y	$�e�hv����76B�࿐v&�X�Fe`w�z;��$���,%䗒S5-�|;��D]�pIy%�ّ�%>IY�/!(��e����vu"i&�g�F8dZ��$�9�I&�~1!"PeY�0BI$��5�!q%�����I���ogM�s����%�G��3���;��x�{"��$�[QFd$�K̮�^R@$���r|��l�^Q���ٷ?O:/��uՁ���[�H8�b]��U,͡ ��Z�J����=���|���@�~J"�JI$�/ba!,�7�AosA ōy��z�d(���E��n�#E� ��E��B����H����S������KM�ݣ:�4�e���,ެ�}~9��j�����~�7c�~�^�[���U�{���v���"�v�=��yl��D5���Xm�u�50e�f���K
8�t������#��!� ��1 P�(ĠL�B�2)BP�BR�4��)JBP�%
P�sǾq�s�fff���yI$�﹜� $-��Թ��R�wY��m��.ΉN�cY��c�f($w��@	w��Y!��ng&�f6��N��B37�I/2�ɏD�D����А�clK5wI�9e-)���R8��
-����[�Y�ȘI$=��H�nޟ��x�.:鴰KD��J+�Q`��d��P�I���0k��W�^���j�+z���$|���K��M泒L&�3�@�lz�.�5=A)	ZC�݂�]`�B��F�(9��a5r�E�l�G����C��.�'g~��d�"U3mg0�	 ݱ�I>�i��ٹ������O�f�֏	g
�VӢ]Өv�D?J�O�fOlZ��w�76�T�$�W��$�	�c��)#��\�c�$�j�� g��r�fC"����mb�I&�|�+� �������l��r�4�c��ѬV���5�{�����(�myŖJ����G[P�v��טZE<V�/�s�5x���ג"">>$&(Zi`�X R���)
$��Z %��
@�P"D�Z%B��������gƾ6㌳$���2%/M堸;:%8vtƪ��?L�Yq�䱧��A#�-�A$n0��*d��y�`��j���vu"zq��L��>�WalS�׹�����N���~މ�j��V��zfd�-䗒I���D�_;�'�h�va	��z��nh�Skm�..2(�!.��Kj���ڐ#��k����s�����r�A��D"PI�_L}%"��1>H�\Gr�q+W��1|��E$�mF���	
�;���BvxT����f� 1�!,����¦�D%�H?�*l�$^u���A#ꖥ{��G5HUQ;�V�ˢ]ӫ�I�%JI%;"}	yO�� .�>��-�"P	{�c�i$��~n�i$tU�,��dY?��	s�?�eLY�b�A(�y���S��->H���/m��ێ�\ne,.���*!9���Ӣ%���':���S�{��В�FxJ;��ǳ���Ҕ���ϧמsx-9z�VOd~��s�z���|��4#BP�$*� L-	H4"C*R!$��H%�J0w|3����JO�Ԃ�,�K�vt��m���2 �	����*��dY,���)��IO7t�2^K{Z!U���{
������u�T���Wb�p�;V�sy��B� ����6���-�z��ߓ9��\����g��)%:�b}�/$�J{<�H���sA�X2���(���n�iI{&���$KL�n�?ϓ'��8?�s�,y�fI
�햔�I%]�焊H
��5��\ʃ(�gzi�R:A��e��޿{�x ���S���6��E�N�;Y$��v�>I%���&�ɩ�tK�uUI~�x���$���O�/� Wc90�K;��.#94G�	 ��r��<+`ŊL��T����H�d�I�u�C"��.y2!�R�%����I%���(�����+%�!
1U�h���U,6��[Hr�=M�F�a����x�ϟ�2uw�U�Q�\{C�����z�z�ν2<�����R��J-@�P)��2� $�R$��D�~���^0.J�4%ڍ\�����
٥�V;@�jlF:�P%��շn�
Mc��]��:�Y�jM�ȗ.#�l����!��l7kP�M�c9&s�D�cc�f���$�
M�L�=XG�����	v��&2B㔌ՙ���.`�;Jl��K�Kˊ�kh����U"ؖ�l�bƵ$��+�j��YlCq��[� m��l�ң�Ο�`��������)n�s��;Y�Zэ,\�61h�6�-&5��Ol�l��9Ƴ�,u�2���$wa�ЉIޗ�H���p�)Ѯ����6y ��A,�h�e�ȟتd6
I�j�H�Ӝ���|z�fR����2X�I%�m�h&Iv��o���i���lN�
<���$�ӝ�p���;:�U���$��L���]�p;C�%;#���ZR%+l�p�/;� ���a'��R��]��÷}��:oM�te7 � $�G�"S�����y�%������q�}��Ж�G��ڄ��$�-nC"YӨv�(�h&|�j��u2�UnĜ��M��Iy%���9O����ͽ-  F(��z�������v۟fv�VfjD��ː��l��.v��`��Y]6Yv�ۍ�OߧϷ�1�����|}� ���ԝ��_����S�>�Z�7.���B)$���A����grX2w.j���8 ����'�1��V�����;���K������o���(�.����ю:9	�^�;�}��o\F*�����X�5m�=q�\�[o�
��HB�
P(�*3*4H� }��1��rO�@$;���R[�fwn�Z|�1JR����2�����@�.L��I�T��Sj�����)y.[�-A~l�$�FݻT+Wt1 �N��Ӓ�vuC�vɞ���}�9Z�K��HH��y��d�=����]dz�Iye�ڟJAP�"\33�v!�;�g�9F�	$�v�@	�Ze�l�=�-�w�S $��^w�n�i	 ��U��
�B��i�qT A���3�28θ�%�����M��Ҵ��.j4�\�9:�������X��Sߞ��>�����8�"C�PD�����!�0����Ʊ�b�W4�Q%y�����!��a�L3�R�$���ڍ:V;��j�+�ܻa������ǒ($�Ż�����}���r�XΓ�pYܹ�6�b3ΐIy#٬�I,}��_����{=~_�������������������<9q��#^�����9P��"�<A�nܷ�+OV
zt��HW�'���i��=۪����Q|����w�dʳ�w'ϵ�ϔDR�t�_��o��L�h~���:�kE��K#g����5�ݒ�tY����}�̞��-{�l�H����n-���q�u1�S���;���;{����m~�S��g��.d�@h�T�?5��Gs��$�P���ט��Dy$�ɒݷ]��s��)o�q��]	��S)��G<?9�7��I��7�5��1}��;{''޹��4����ɺut�&��W9�(G�[���׍v�=�Vn�������<]�����۝���&v��ϴ�};�j���u��v53}����7*��ԗ���x��Ǯ�,�q�w7�ٯVOp۽��|S���F�s
R�<!�{l`ыsݗ[��o;�t~G�6}��w�(����w�	t�����#�8�}��� ��9t^�5��ܞAo���"��9nU`��0ɤ�vf���)`�����x�E����\� ��@x掤�
t*e�/*��,��9�ۮ&3V�Ppz����p��Cw��<��M{z<H�����<�)�]��������k�RF>=z2TY�9�N\ihXk�e�
i1�dY��C��ڌ��WK�E�}�r���i�C��e����s˞wv�r�|wV�Q�|u�޶b>��@Bszu�2��8혻ɝ�Ѻ{�	�}��*h�!]ÖY+a�J�� �O�$�?�<�I��e�������+8D�mm�N�3y�;μ�R��s��ε��PD �8���h��m�vy��7q�f��rG�������"!ٶ�A�Y�#;$��3ZF�z�{VB��	�N.Y�.��֙�v�[Zwi�gv�vZHgY���ós�.8��r�3-�DQ[7v�DTYn'�[je�(��(R99m�!����<����B�(��B�u�qD�Ίq�(8��J�'m�]e�Y�ѝ9g�[d�"��vՇN��P�)9lge��GeZ�M����qǇe����e�De�-:I6���N���1[n�Y�NTm�rN.K�hm�ؗ6��:Úݶ;�̳���ӥ�n������w��%��m�Vwht�d�F�L�(��h�QbA()�	��B�"
�rKg$��';=�� ���{����~�'���
�����wwY�s�T��Ȅ5Ϡ�OJ�%�	/$��y�I%��˔HǢZ.tD��s�4�����$�{���̓��^�� w��$�Kt�8�Ӳq���]9��>�>L޿m�u5��)�h�I����-�Ao.�U�Yf<X�p]������:kYXlB�j�5���Z��*M�B���wܿe����]�t���
9FL��+��b�Y�$��ϼ�>J&���}t�٧���i�R$��h�$��L�9	ΝURE�zDI&�CC�TkWdX{�0d�E�Y�$^K_y��&/6���vg�� 7��2f%"���T�&�h�%�<���A+xɃH�?z�ju�%�%x�L���x3우W3��\pk]<D�\�3�l�{q�D��h^I$����3�f�[�������F��pɓ.��zf��7�O�E�=$�1x�b+j������)��g��'�� G��޲�d�34H�j��!9��Ȏy��Pٱ�wP؇� ? ���4�+@�A�Pҋ@�|y������?��&��*ݫwm��7^ru���:%�Wt��9FN:H+�h$	$��	&_�X�#0nf�d�N%����m�m tWJ儤v&�d�d��,s6�jEڬ�D&��L�}��Y�ʉv����?oz�30H�oLJ�3y�K��/�WcB��Ժ)�Q�Z��}c�	�ɝ����d(�2� ��$�2\�U�_�� 7�w}�M�����:ɘ7X����<�x����E�:��$Y��ȉ��e��%�$�Vԓ�!'o[�6X�K�R��x&|�}n�bd2�6�"��S:(��^I�Y�MڙO�MbH%
�e�y$OM�-)$�K�X޺��j$G!�=���X�<��Kf����g.8wUT:��~�"�$lց
�oCP���]�}�j��I�%�$K�okG�7��E��悳�:���ed�<�?�=���t���W�v	b�Ǖ^��zg�>�Є|��vJ��'h��m}��^����ߛ�;��{doO����|H�B�4 �߶�?�8\����Q�k�V�n-�]l��Y��Y�ÐhF�1�L䲍��9kƨ�mr!n�����ͣ��44��mS\�%̆�e6m�h�,��,��˦�/����	N�\[��cZ�lGU��&��� %���=q�{�1�{j�ID�c)n�P\�5X�z������jYu�T�H������e4n%�lԪ���8Hjh��zo]@[T��t�a.��&�3�R�b��L*\�.�	�UF9k�z�����2�+����Օ2�/�v%�  �ݭ�'zmD����U�J)$�vX���[��ɑw4*�n��H$���suD��,�h��A�%��/Ov�[�̝�3���afs/��e�̴����A�d�v��ǽt���$���:I$����q�N��H���!"I��G�O��&jRb�j�$������i��񪆹t��%nD�I$K;�!g����D^P��@�.��7-)/b6m)E�&tQ�)7s@��>�B踉
Ze�Oi�U\��kI�ږ��+�WkD"�^\��&V8�a��|3o�ijkkÓ���lUַP�5-ʗivD��GD���܇)�ʫ	c�Y˂��w+u2�x$I�ց	 +_�DϒU�c�n8�n�uu��U-) ^J�%�h�gb��3��TPK�*'�I`���Қ�w��?Va���W^�'����{M�h�z������+�j�g�Uٞ�1�孬T��쉜��t�*�Z���Q�"��Hs��{����o��>�%yosDy 	Aw��&Q^K+YF�1�h��S��cO�ɑw4*�\��L$o�b|e$��9W����c��OsXI����ra ��tt�O�!W���b��ܱN�*��橀1�5��f��3y��ց	$�J�� Dy$���1;���{�'�3dC9��'�&��b�s��O��#�I �l��%e�������H��<��^Yq� ��f��<ʔ���e������s��Rv�@�E�Ά��1ff�`��Aɶ�[��V8!�29�f`�g��P<��u ��=䛵��H����e$I����O�Z�,.�33U��y��Zz�I=9"�]���L��w��;t#�I���fK�����]L��A%Y"I� ��*RIl޻��;n�mP�v���4E,-��4��lR@����q�H���c=�~އwz]��d�bګ�_OyE��� �w��{�{K��� �]������M�.5]^��'�ٔA� <>�{�{�1� @$A}�}"�^�(��9��)N��l?�&E�τ��M����
vW����U�3 �Iy$)��S�G��I%ݍm��P�@��ې~��d`��������e�$��h�)�D�o]ɘ�9���ޏAΡ3�CeH�30H�{�������u�O�Ñ���84z�!9���TLi�1X�c��Z)B�J�й.� T�����/�6��������tdO���3d[t#I ��	�g��{J=a=�H�(�����RG��2��frQ�J�g ��0�wWt���cL���_%L����	J��m\І�S�p�K/k	N�'r໇u�Mp�(�	{5�Ф 	���O3v���	!O���  ~���A?|��<\�"Ck޷���n��f7�^Ǵ����$J[��	$����G���ЦmBE��-P� �8n��,V�����fN�]�셉p�=�Rl�c%^WP �9�<������n׳Į��n�&b�������?�������E�t�,�sB�K7E��^I%?C�ҩ]nCWk<n�I]k�I$�[����]�dJ�����oG���)]6�έؚg+Gevu�Y��X1+���W�\���ir�a���/߉W-�s���x�dI&�Z!/$37��4��.���sU]O�#"_%HIy"v�B}6�&��s2J�~�))w�b�8��F�D�tg����3f4B�0%�1�	�$�*��h�{�2�󔥾o,�H�,RI��F���m+�u���	/�j*�N�=�U$�I+�g&AoFȂ��:	ܸ.��UR����8>���kl��E��.�3$7fdL�O>�B�#N�c��$�kT$/l���]2d���f�ˊ�M�I.�m��q*'f����3�K�$���A2M��*R>>�/&m1���fۤl�Rᜡu-׻�`V�.xZ���ܽr�0��l��غ{޷���������!�C��0�2�M^;�WJ`���="���I>O=!?5���L�-X$(!m�ѓ(%�l�
��T6k���u�{Z�;9��.�F�n0��˪�mՋ���
@�l�6��,#���\Ѻ+��+()3p;[
��Y��Ɖ�!�FF�Q�k[��lF�ڲ�"JZ�!K-�^�-��×vU ���]J�W; ���\m46��Ɩ`
�#S�Y�p]�{l5�+i�U�V[#�fc��s,HQ��Blc;e���f�H�Kj��.p"�1�d���#X:L����̖sK<��ؓ+�/$��}v�,D���*횋Kq��lۻJ��= "�AuMȑO_��Ke2�i��]����I;?�����*	��9��!�^ݞ�2D���&B*��jym5]��R�Bq�b�� �зp��~�S��$|���\e$��������A���I%7<�L��	76�z��C�� �I��D���4�ؙw�ݲ��MS�"|�+�m�-!$��[|���A������É%="�,c9	ܸ.��@����e��"Ow3���|	s3��I<oH�e$�ٲ��Ik_,��5�k��F�3��K3�G�gM��n��#��f�s�r��,]a��Uf�a����Ox4�2�8?A��m�� �R݉tJ�H�|�{��9�R�;�'RO��-)(��-��Y2.�9S��I���z�U����Թ��nL9=��*�:-#C	���3�z������� ˨���z|,ꤍb�om��_R��o.���]���:�;�S6:it/��=�}��P"��1���(/�>Q��d�J�P���m���ԥ�l�~���ΐ�nG;u������|��$
Y�=	y%�e]��f���q{�DߒQm�-  �I�|�С��o�I&I�
�I��!�U,�Ǚ[F���|�¾�~�3$M�u� $�K��AWs,Z�dcv�2��-)#}H!!�E39(ɐ���B@$�]WQ �+���R��)+�X��K�U�@�PI.��)�l�S[���/�փ�������,��Ye�b�������h1ȡ-@��˭f�cS�=��=�2��p�y5��H$�;���K�H����(���g��
�ִ����K����%��8d�X�s/)t�ă(%-�����6��D`t�I?��4JH"�ܞ�"Q^K:�������]kJJoFe�1%��sB��m�D"I�މ�2I'�/G��3g^��`ήű�6��f�����������$��ۜ��h��.��8/��D�~�NC�1ٗ4љh]�x�Y�Cȯ�����~o��Q�o2ߵ�E�]��dq*����\�:w�
y\�`=��E�6�A#S- BA$��G\��$���t3à�k��NUy$�u��i4-��y�I�qTJm�`T��	F4t1�j�։�$�S<���F���QI ���Ӟf��f�}��շM4Ņ��r��b�9N�3�)3�B�Q���K�m.�VݦfTeY��޽��
I,�L�J=�H��t�Y�I$�We$�O��-)76z��y)�h�PH�NǄ�\�9gw;�uUKGL�%��6/'4'�U�<Z�B%�ܜ�3�;��F�D�$��&5e=g��]��S9�i=��0fE���K�&$��H%�b]/$�W7�׋0�#�|��%䗂"QH����(�U�0,Ļ�A.�d�U+;��r�;$ :���5l!*RH%�!�$y��d7�����mEIx;�K�?;L�<��ز�;�֖���	�.�6�˂G�}���>�����	{7��������/s�qb���QYnUUK�LA���� ��~I �#�H���JB,��S�w�
~]2�I/$k>h^g��]�t1��2&RI=��iH�仵��U^v>���s��Ðz�;A���J�.�b]Hg,0UC�֔M��6:��[s��Ŗ�>_����ԡ��I�:$%$���C�I ���
��p69��c� �����P	/�Ζ��Ź�* �%39(��G��O��g�^M�*�8��>��L��H=�d���H��c�F�]�ç�$��%(۶���;�A�3��ṄI 	=���D���,٩���e�=:2�(���ZBH�K�Z$m�n4�,�
�.˨�hf�<����c��	]���$��AvkDy"O>���"�~�kV����A%��R��c�jO�
b]̉Ĺ휒M��X2\��n�e97���13䉮�B$�}�+G����|��ӧ������O��������x�=��?���*����ɪz���E�? Z9ҽ���qk�U}ǅ��;����2..���Y0�)��N�X�˸n�^��{�ܼR]t|=%���E�P���6O�!���Ɋ�����j�|�9P̮b&y��Ӽnu��C ��+���{�+'Ӽi�4A�LL�I��3���ag��ƥ��1�/��|=�tv�[�,;�_J�3��(��8�[i�Q�l�I8�'1鱚!��ʪ��]�O<�	v
=����S�Ӊ{<}-'��J��7"�/{=���Ĕ>�}oZ�A�?"�s�|ލS��骭H*|:{���2m>zuLOz(��i<WQj�3�v��nv�Ϟ.��Oi����� ]���{b�8��9���/!�\ӣX�k{����:3��,S|��ʷ�c�������/)&�ƶ���k�������xQ����Ô ��4�)FrU<{χ���/i^a���q�6�rMA�E�d<>�K4LE2�{���!c&�w��J*�jkӯ��:��y|A�a��A�������{��tA���:f�p���Vq��p����9����3�p{����DS,���}X�����������p8&����#�z�z{M��>�d�s��{�� ���|=���.u�c`�9�&�Z���������]wF%��3�2�,�%�5�3�rψ�w7j{����ũ>ky�xd@���x�$�/oW�kv�x-�����W��>~�7y�B�^��:�;�W�K�޵I�:�r��@�j�����X�-���b�e!�YYX�jt�����~�cI�7�8����`I�}H�,��":+���҂r�s5Z��٣-#ktէq�E�wf�	�:��{�n���֋+m֑��e�H�7731�!��)Fq���m�t�$�+6�l�w����E'w��ò��k!e��Aaml��a6�y��C����[EÄ���M��ݴiH�m������-���y�ĝ�qȑNzZ'DQrI��O�EF��ݶy�&�qͼ�֯2	KҷB��'fp��}�������� Amn=�fG^Y%�pDv��g��{աA��|>wok�#��A�����H�p|�	�_I�r�B����(㲴�>VW����,[ZQvagi���Ք�:����%/7vu�
^[�9�:�ÚC�F���Ӂ|z�u�%�<�(����5te�@ţ�pCm���$�JD��͡F�q�i�k��..��uT�]���<ǆ4�c�e4ؙ��/`�عc[�qr-�\ǃ�����L�Bl���pQ�M��X�W����V���i�/.v�"�5yx�h.5`C\��R�رɐsc��0��M4(��q�1Z�T[tU�e%�Y�l
�!�p9MI��$Xbk��t��2̰��2�6EM���òXM#4rLXZ	i��l����A���Yc�^Y��10�5G��,�3i���`�qZ��s�r�hMt�MyWR��m�V�-rJ�l��Yc)��5Q��ź_�'<��]y��G#�jŉ+dL��<�ڍ��xu�K�ճ9e�Rk0@��1f#t���Yuo5.c��1�)u�bl6�gU�����o��mɦ��t[ ���[$2�6�s�,`��%L�YQ@�M3k5��*1Ơ�{K��
#jƌV[Z��+�۰*�i��\�Ù��qZ��s.�9�5���� �s֤P-�#hL/!�:4��j-.���d�B<��.�]t�4:����7�l�.K
#j�VY���V����R��u�cT�ѐ���fٶ� �*Զ�h@�l^
�*&-Ѯ*�H�؆b�Sfˍk�ؚ��ִ؉ Ц��)M-E�Pڳ0f�Wk��	e�Y������P����a�Α�f�6�`�K
U3ÃP�	+Yfaڮ�h�"��kT:��Qs����ː�����eme4�#Sl�6$@i�D+�Kt�j��%�gh����,��Që��W"]4���1M��TR5�f�����VQ�a�ڙJ��U٥.Iy�:�XC��G�3$��cT��k��V���5�;]�x�l74�۴Q��s�Y�X:�s���ml8BlAc�P��*��K3j�X�x�����x�A �����n��nc����R���(±��J�>VN�zx�7��1K�ض<	2��2��CclK��st����w�$��L�+l�5��4�u�d&�!�l�XE�5MгlÜ�Ә�ۡLMv8u�#�6B,��;V,E��3� ],�Z�]b�v�i���Լ�*��L	�Bk�`��Ԍm�m�Nڻ�$ �D���n`���fM�Æ.��	�)��-�1��ũ��.�g8�s��ljیS�;Mxkk�+���6�mqv���B�ơ�XCl��&��+YS�J�4�ٞ��͵Z.l�!���4K4`Q6ܫ��49��ڠlU�t[��O���r�mv9��~���>&��H��D$I.}�@-ؕ�c��j���C"����֌�rH$���s��Rp�vE�Q)��F �lC⋳�[���v�klH�I$�^�zd2^�K��zD�QA)畆�3�F"D� ��Ĕ��lֈD��W H/�Q���[PFٯ8M,�Dג@%׍��3x3��R��f�b�� ��Gb�('�IyԒF�! I �]"d$��~��Y�}����f8@%�1�����	8d��s�����bL��I��bYS�����lI�ԗ��W�2I/՗"}(��5�T�(g��vy�0�bHp���1JR2De�su�eYj�e��e�6�e�P;C�nO�Jb]�&���zZ|� �d���}��Dӈ���;��x��B$���"��*ZB,��S�w�S��#�������rVD���iO5������_2ik�x�=������;	%�0s��vӝ��r��j�̗���;//)Ĩ�����]���Vn@�H6��L��gyJ�탈�2�zn89�S,S�.&K7sǉ$�މ�� �knۃ�zz� �N�$���$�]���Ĕ�� H)��>�楬�پ$��<	$[�f���>$�wGgOE��O��c�.{-���gw;�u��bݛ���Z�����K�G��y3�A#Ż�#�L�����z]�S�֌��1�#�a��*L�	���RSf��F��2dP��]:�~�x]0d��s��G��{6'ĐD���eyF�0��KN6��\���|ٽ�&/F�֟ȤȻ�|��y�5x*���(�t�o��O�U�G����m���,�S]m��n
[���"�@��ۙ�����y����Ʒ'���$'aتE��D�fT6UOTF�ӯ�L��r,o��t�-m/_���S�ށ�a�)��;{��/OnX2v�.�}!�y���O�������#}��>��0 �ý ̏���Z�a�&h�K}��JZ�m�ˬ���	񆜨�|	$/5�HI]����ޖN�fz6$δ�����bAZ� A$�ogE�7�gރc�T�oHA�6 ��]�on�\e�<1���.�!�iV$�
�:9���k+.�M��9r#�
�hᭉ�MZ��gA�� ��w���dg���'����SD�:�Z���of�v�ρ ��{��h�Rt��,��",��x�Y��Ƨ||]q�D���'���d��B�"�_(��
m��֜"d]�	�nJ��I.��������I�n������I�6y1vE�:��臗����� �=�I�A!nwH���iѱJ�Z(e��T*�!R�mj�S�^U�:90/%2&B�a}�ڡ'[p�XZ(��.֫1{q�oq� \'Z�u�O�#���{� �ŀ?s�ǟ���.��$����f��I*���!6Ev5#6$?M�x�J����>,ݛ�><ñw3�b��-��� iz��4�J�eWp�j��#���	��y��������z�U߿N�{RZ���xOp �Vݸ�|H[�� ��F�Ǹ-o� ]W<Lu�k3���w�dE>�U���Z��ym� �		ށ�|�7�Io-���V?qn�/�����Rt����I��x�uvĒH:��8eugAf�f�� �$!��x�B�̙�#����!3$�d�&ۭ��5����|�zx�	�꽙'��u�k�t۴�ۺ2�{��P�Ɏ�@�B��&.Ȼ�^�����|O�_l=��V��.S$�=�y��A>Y}� ג �v�X�����j�����������:��n��
g_�=����y�1Fv<�39�{�"UN�I���N�XK(�ٶe3/IU�÷y��iNY����g<��l{VeM5�H�\�j��&Q)C�d�dRKH!q��EHͭ���v�V.Rf�Z�@"]��50h�ĺe�n%ĠA�W��#peBn"�4yf����\�����Ԏ1�f��%֔�^GYIP���YI����e��ΠV��j��W�t��m��5w&ؚ�v�:��%ԣ�eK()��~&������z�]`�\��v�a�t�iL\�KSR�*�vv��AY������O��*��P�tg��+�����S��$��׏��v������ A$��ɒCh�DId33��dݰ �"��nb؇{�x���O |@+3�D�@-ݮ �i9�R����T���3;���R}���H��׈"<�G�y%z�5��M��5o^��$��tD�X���f,X;�����yTq+]�I[wb|A-���n��JyQ�d��L��Ө5���c"A�{q�]�f8����,�މ��_@�A:�� ��̓��)Cd��ff6]r�C3n�5�k��Sk0�tV���dì�X����p�k.fA�׀@>'���#Ǟ���������'�$�׏=j�iwb��vb�d���@�G���n�R���^��``���o9��t��{}���@�_�c�{�g���V��C8P��_���}��v{�sn��Ǽ=�*f> �O���	�����	�=MM�a�c�e�~�-�?�=% Y���3%s��� ��^HAk�Ŋ:�����v���Km� �|����D���V��Y��ԁ4��0�L���;4M������zU�^@Y����-�}8�S:`�ŋs2����$��͉.�����ι\�A mW	$.�������GL������/�,`�@a��(�	��ln�v��!mG0�9H�#ud�/��,�7��$Ȼ ��v��@�f�x�I��ސ'���l��>*yY	Ǿ���Cg��;�S=,׍�7�PE@�N7t� ���>b�>GJ��.)Ud�\�>}Չ��Ӓ�� ��x׷� ������T��퓳S�Y{��;�{�76�֤���t�9po���������J|+��c�j��M�վ�q�2d�n�S��:!��5������ �ݿdH }b��ff�<�۶�S��YlA�G��>޼�$���$�m�������8���X��Y����Z���A ����,���uM�����q ���d��kz#lN=]Be���ϸⵠ��a[	�U���j3E��sc%%J�E�6i�7\k��������EkY��۹0�O�n��I �{�|`^T+�Ν�>�qu��H%�of�NZ��I&b�dI�{�ꇓ�����%[���HD���1'<��1����zz�P䦰i>er$�;�S"r��|H���A����'qE�h�ۛ�>�$����y�N�t鋈�M���u&n�א
&{bI� _�۰#��-���?�Zw��8}e�^&CT�ʧ�}�$���t� x�k_����V�G}������M���߈Y��>�~B��U^��+5L�����U��2	�~��4R��8s�m��H5��z�����'ӕ�"I/ۮ �m���e�1�h��vv��sa���fj+�Mh�j��6���k�b]�r�����"���1frC8g]*�c� ���y/��������e>h�[6�f@'ė�؂h�kvvp�ŋs2\��^Ap��2��ځ��=>��:�m�- @�ז�?Lα�DV4�pa��|LP�,e���v.�D��=Ǡ�H6����fV��֢���j��I�6	�6�z6˅��"��;�S3� <�6zqj��H��A$�j��nwN��7G1|�x.��Z��.�t鋉�PL�Z��$��c���6��� �Z�p#Ē<�]�'�_�Q�k";��2���٢q� ��A;�-����.�:2���g��o����;{�"�X)���gs��"�
C� >�����PJ�Lդ���M�v��R���9�9�Jf�]��[5��]mZմfC��GuP��ԣK��C�M1E��3@����;Y��@(v�e�Yp�B-�����9��l �WJUa�pB�C�%63ʵ��f�� s`�,�+�%��*�^�!�k��Z$��4`4�/E]aM�C�<|4��+k�����H�6;:aƅ#���!˶3�]Xճ0�ىt�����(L�Ý�ّr��A%�7�A��n_^ݸ�A �u��|��Ź�g$3�u3m�R$݉�U7q�̊�	����K�oL�UO�Ի� �:�Yn��3,�ܸ��p�Y�m�D�w������):n��;��_�g�莉$Fi��Y�H�b��O���<�x�_��O�'�7�2I%��w�鱟������x,<��a7���^x��W�̈�فOI�f�U*�:�v3�@$��d~����11���������]��Dߞ6�(��x�`�k`�0�XLYmm�]���Lu���{���#�U�ĒZ�$�A>�����K���o@�O�j�Ȓ��h�Y3bJ�����opy���ШFS��oN#�ho��g�����sf{��i��>$\6l��\��C�z�ۂ�5{�W F�=��1Χ?y���|�mX�!��t>���_^��A$��;���}�8�w-��{V#!��h�#H�;"��v.bO��j$x�O��k��TzP�-.�OF�%���@$./���O��-���;,���������>��}tf�A��n8�@ Nv�H$�	|� �m��M�j���ض�Nρ>Ω��PG�zu1�rJ8p�췧�m���;Vc�f�F]�H��}�� 5��G��_5����T@MΜbɝ�G!�ԥu�F\\́]��Z�#3kF�\�jU��4��~O�cY9wp���ꍑ>$��DH'��� ͦf&��vM�\h_/`/'�`m�,����W��`����5Y��.	���H��z|f'��F�e������`�6��0p�d�~�ۮ����w��1������������ۧ�g�����w����Ǉ������,��y��C��<���_y.t,]T�ƒq�|?�ܟ�1HY�a�D"�7�{������gֶ������MZ���~D�z9(�[���V�T�����K#/j��`Aطq�6�����/�����r�� л��r����X��E��˷�m���`S4{����D�f�Y�sg���#�N����,p^������kɑv?7�%�@Ū|��]�ʠ�K���K����ll����ዸ�%�w�V��ӻ���݆�tG���onX�ë��*�0�� �����u�dMY���'�p�����sn�٩��	V�x�vp��(�&����;u�7*K�b��Z�½Ў�|��-�G����{(c$��<N��*ǳ�7�&�;���=�2�r�)��#N�|9'����l{ۧ���G�r��-��m�K����[�_e�c��� �v�Z���3�X07Y�l��n�6x�箤W_>���/���P�.#I��y��A�<Hg�<^|Vp[P��j-�:�-�?nw��ޛ�}�F��}�xz����B��0F���Ў��z�qn�?:%���4��B�@��ߍ��ݹ)�ty�x���z?e��@�wy������b.�;��y���[F�ҨN�w΋��n??m̙��K�΍N��q���?�Jp��N���!��N��/]q�d���L40��bGF�-A�P|fD���<Z�h�� ��D�`�M(}�a�i!g=��f��A8�.'� �~[�"-�݈$�&�E0c�M$p�g�\^�$�N�3F0F�w�ۂN��8Yn#��''9�Dp9�=���p���*J[%m������ �)8.).N���;�:���ب�
ﵭ��s����'G)�Vw�a嶭���À����t��� �om�u�ɕ�X⼭-��^������<��������
N�����)�,/l$����D��	�k�'	�r2q�-��Y̜��$.��C�㯵�vq�f۳�W�w��۽�%^vq�^ڃ�8(��;W���q�Y��}�qQ�b�c�Bp�٪:{u����p7²M��xg���]u�������ߠA1�d�;"���\��oT�3mMW}:�ס����8�w��$������#�gO�2h��RI�x�Xش���	� �Ή89�2"����H��$�l�>%�;�p�/��6Q�?����߳�E:n�\��mhi���2]���2SS#\�ن4Yb�F+��������B�V!p��Q#ʮ3bA%ڻ�L�޵&�~��Ó��j�N�q�.ȆN]��L�箙#o�՚�ڕ�z	o�h��I>n��@%D����uv�6o��ع.��L\@Ku�؉&���$���_��*n� O�]��I!���=A=� �"�d�9�WXƮ�T�Nۈ�>'���3�A �wW�z<�V����4<�0i٪������b*M�{�:���<�D�g��8���{��{�ox9�
;-��=�{$;�=ۜ�Q���wE� ����O�j�G��/��[]�f�v.fA��uA�[�ع�o8f�rE��zD�	l�ɟIn��݊.9�}?�z=0���:�+��2,�E���+�惠$Ŗ2`3��ͳ9(|���fch�wΩ�g��Ή �m쁊6I,��ՂZ�= ��ٓ&/����J)���E<N$M�!��ZO�'ĂF����I��wG���s[�R�&��z#���LHd�;�i�4�� �Ik� �l�h[��_7U��I$�ݙ �[{�CI�]ӳ��\D��o>艜e��P��Lx�u�Q��ȀI+w�M��o7*Ysd�c�s�Tlb"��d�9�!6���"[���V�H�wf:v������KVd��~�S�n����1&\�z�)��e�%aa�p��0u'%H��L�M��Tu�c{zs=:��Ϸ�h���ã�yr��<jyΚu~xtw-�ϞiI݀A��0�
�-5���$@�B5iK�qX\�ɖ.�t�H�T�����%p,����p��B�,u�
�Bm7Ʈ\�13a��68r���2X���Qu�+B��A��ц4l0Bd���-�hCpP:�
C3&���k��lRgZ�3��7F�-�u�Y�Sl�q-]d%U��H�&��R�]+U%c�ApCv�Ta}��[���,�a�K(��ї5�2�	�0�M�&T�0.�,��&�� �?Z{�V�?�ƶ�H�Kn� ��mށ>/�h�ǎ*�nnfe|�}�_�.Ŝ;�,������<N�ݝ��������,^��@�ށ$��i!B;9�O�p�,��	��O��]B����Ê9����_S���K_l�m�	n�4�"�'t�3�箝��5r��G�6���� �O����$�[��LM+:"��訃�qä��g,���)�^y"U�dO�EJ5y��4�i/�ޙ�H� �S�$�މ�j�23ʿ?۵�9a���[��X>L�43%qT�n���e�[�i�&��������i*,�����d�A]x����M����k�)��a��}�� ]��mM"��`ዱs6��0���a���YU���q�\�a4�mA�i�@z����;��a�Z��]��Ƚ���g>��ϻ��77��=,���~����O�W�C��'���ߦA>3E�4�i��b���v,�òL]�
Ƈ�A ����3b�kue�vȎ��Gz���/�I�!�c��Ki:YK�%���&��:{f��D�I �+�ɒ|H-��ϑ0��e�c��<�K4���'t�D�<�X�Z���ӗ:�%�l�H�H��� �w���2O�n��D��x|����z��y�t�TܬpL�j�tSM	�c �)KK�C9j�ˆi��)|��.�uff.>��v�x�I^�D�H���
�,�{���G@�~^Dnޙ�Q��&`��IM���z�5Ttf��;�$����I ��<n\��v�X�z*�O��
�q�'`�wb�P��"Hj�x$z<޼�ǲ9M3'<�f�TAxu"n	��Mm��z#�����g�	�.VL�Ӭ̜������У!F�gwl;[^�����4&eu��Y�?fz=>�k��xKwgH�Aj���b���fL�òL]ˉMtS�=41��V�	��&"��A$���O�{�*q'VC��	���O��,����ȟQ!zxO���M4\Wte�}��t̂D�/���H]�����}�nve]}�D���6�)5�±�.\T˞�3��b��˥�^]b�h˲������s���o�{�Yek���� �� ��珛�2#��DF�/<�#��wN�X;qh�"b�R������sr�&�CwtA$��� ��vb�RO�٣}���k%�ff������ �o �A�����2S��$7nO�	��� 
�'Y�v�3>
��b�oy���&���Ɉ>^I�7n$��oN�<��j14�9�ueh�W�ע��y�G���^�`�>��m�y㓦��T���^����J�� 022���'M���xj�Xx�q �����d��᭷fN;���̃X��	$�ןD��j�I��^�A>S�<H$cn�g�|Ύ��=3%�7H��?o���ƈ����B�ͦ`ؗ]wi6R�`��5����'�	�'K'tA@�v<ܯb�	*�_H���0<���6�� ���p +af�,�;��Q]3�F�5�7N��U�n�,�^�I .� ߊ�"A<-���sM��r]ӳ�	�8�7�ЏI6���H$�i����
���zQM��$��:M�Xfg%�A5@�wb��i@XhA>:���=�~ͪ�$�[��Zj�\�
`���WfO���rx�`0�bӾ��p�n�v��ו�%�B��/�L�L��)��'�ͽ������J�U�؃[FCs��4ef���3���Vv)�{��� da*��ф3e�9�Ĝq�u"��K�i��!=�I�����S�#��������Z�����J�V�d�^6{]4��U��J<�F3���	�Υ�R*Lh�.pf�bm��
�nQv.��KoQ2qj���3�s�Մ[{�,Ɩ����]5&�L=3.�N�7[fa�[� �@)�uJ��@5(�[���d�� �2��Ma*�Y�].�Y4GMl\Z�K��*m�ܑ؅Ź��g$�vZTR7�x�z��O�-�E�)�U΍��3��W;T���ص�M(��]g}��E)��ц+v������O���ĂI���������}� y��d7č.��G��^���m�WsR�T�ک���K�d�$����z�:�kU+�}���,��gp�Ӵ�O[3�I%��
�E�wȨ����I:�{3�H$�臘6��vr�9g&�A�vJ�2����!��c�H$[w� ����͑��^�4�;hd-D�,��]	�SwG���-�]��E��|�k�&$:!K���o\4��β׭���`~�{���n��W0�MJkUu0m�V!,˝))�˥��a	�~���a���!��I ��Ǡ�>M���g�\��d���fI5w@�zk-�&p�:,]��5�.ޏ"}����]��ujS����F�M?Lc�fsco�T\�/�%@�
�c���klgx.���͵f�c؆Z� a�*��-6[�Xm�$��<>�����I ����w��5wr^�z�12�DӐHp��AA�N!9+|kf#�'�_k�'�[f�'���؂���~@����}Mݎ'��Y��b��;�h��]�_viB���3uq�$�U�;��$<oN
�����z�'g�"�h�����D�mׂJ�v?dO�u�̋��L�W��x��V���H��ޙ���7��	��@�9t%�p6ᡙ�0�.]���&s�ƪ�ẺWE���Կ"��3�c�
|�|IY��I$�>��z�t]��DL�;F%��B$3f��H�ɝ˻�Ř��澩n����ejj8J��A��2���~}���v��T�L�K��3�	�d�fMsˈ \��$��}��x΃;��ӆ%�X��{����l��o�G�:��9߸����ݳ��K���2���Ĝ�+�Jp�H���;���s毽�˿� ��lz =ϿD��$hf�@�ȧ��1N�9F[ 
}���^$u��� �ǋ�v�]5	~�01�#�-����b��;�i����zK_t����%��j���՜�	&z;&A$����w�����~�S�w���Z��j;h�$ʘ�	�sKd�L�[+ r��*��ۜ�N���63�L�k�|I�Ȓ|H-��-�"[AM����q17�}�92$C�٧�fN�����>0�x��6]	g���|� �[�m6�ω6�Ǡ����\���m�Z�P'��P�,�]܆L]	՝1�$[�b$莬���߆x��J��O��[{b�4��38`�&N�d��:؎y}�obw[�I�9��|�����>�?LFH��.�Z�	�4N�l���8u�s��G룯⏹�W�����>I-��-���ڥ�b��n��h��[��mY*��@|>��rD�����f�@�ȧ �����	'q�#���,'�Vx��T	;����B��#�=e�N���ɚ���G��q��3w#6�ۃmD4�F��4*�΃8=wi�;���L��L��ĀC^��?��H+���{��ոث̩��K�tA��cC�wpȺg%lk�$�6���}�QTa30[��"A$��b��~q��(�EHj[�#��k��pȖd������ǐO��ha4������AǼ�=>V���:Y�Ӈ)1t"{�qTL��$�ݷA ������j�m���W�Ί~�K;'���łE�� �^�:$��ܹ.�츬rF�DA$�=��|K�oH�W�����Ǘ�Ƿ������NϏ�������g����{=�og����]{[b��C�����wl��4j����g�=��.jJ���=��Xs^'��5"�Dͽ���{
���7��y\�������z����}Jӌ�g=�I͞��;=���Ҙl9�����ܹ�=�gj�ր_�K7���p�3�ɍs����ൣ�i�]Z�?����m¾���]�,h=�[�ה�$'jxf���Oq<��^h���KWϥ����>oݹn���/(��^�1�XiK
��w�ї���S*�ݧ/�q�^ڕY쿝G��������C�����y��<#D��k��u>�<�lj����gu�)~�#��W��$�NE;���9�-�����3#��
8j�Ho���N{���>�{Y��_`�8ogWs��Y����opum���vհ���۾p.A�\B���o���7|s{۞@y�k�T�NM���/zo�?O�\:��o��$m읹��.�Ƶ�+s��{{�s4>><��6v��#և >�$�m%��	nh]_��#�u; z8}J����=V������S���3�a���ɜ�o��P]�'���qzb���x�YCq��v�F�:���p��z{]����ܴ�:2f���ו��b9�Y�.��\^��b�O�W�L��x_mH��^��$��yA��ܘ��Wڻ��Ue3�-G	s����K.lǔ�8�|ɳ�q�}����o�����j����{,W#y|�umOq]O���Mu�gE7�{����-�b�7���/�ح�b�Ĕ!�?I��)9!W�dE�,�|�!�8�ya�ARO�[���7E������l..��Nq�D�|��ob�ϝ_{4�w�#�n�N!Ϙq����GZEwμﶎ��ʼ�����u�b��:�{w���enG�����kw�twη(�U���o��΃�k̲��׷��|��|���1��֧�onl����ٶ�+�j�3�"����ٻ�����vw���l�Ȇ֙����y�n����ݑ�m���t6��(rj��&6͠����|.�_>�l��-�-�B�qX	� �b<��DB���1
:V�a&˚jꄣ����59�\hB�J�\�3��f��j2�k�6PFl�mɹ@P�G�6f�2Z�lWK���^f6�"��MD�r�3�Z\�(�,�Gf�$��f�@�]aP�B���:�E���i������͕��v�cA�L�IM-3�u��l�,���X]�(�XE�ҖT4Cf�xEҹ��f�F�f!mxJ,�	qUV8e8[խB�]���G(\˚h�0�э̷cL�9����AqhM6����0��],�1^6c�4��z�R���v�'&�HP�)��7.����,E�vj�f!��ѕՖ��D���ֲ��qu�-S@@�b�ˀ(�r,Λ9)�(Gn�L�(��(���d�2�J�uk�,v���EoWVk��Q)��t()[��VVc#s�[qX,�`-��e���T@��TjS��6���TjGK�ƀA��x	pP)�X�V�ڹ%�K�ƚ��ܦӶ��*��KJ0��l�!P� �Z�sC]����a	�c�"�.F���l�6rd�MsL�&�h��^�5+B�0ge ��n!���f�Q53,���:]b��aik@[ (m��ʺX[���l�,�	K��� 3��e[sTۈ��tI�,
@������u�-����*i���ю�l�[���aY�`m6X�g$�������mc�Ę���f�]��n��1-�Z`eІP�T1��ZW�	���̼�-�G�3�a-�:YCi�c��64�����qT���U���gZ.uҘ�<㈪U.��q�Z�(��5L0�%.�t�RW��b+�	tf�s� L�g�T���s,HE�W�mH�Uٖ�%Er����f5�k0�J���ڝ��60���\��Uˢ��1h2G�s�v���-u�*,�m�X`�6KW���YUn�,%h�R�%���҆B�VT֟�K6#hR��3����@.�U��x��͌m�`i��5�%�V�Օݪ��f���2�F˲e�� U�9���FV�.2M{Ce�b��VRcS	e��.��x�)@��%W	u�d�c�4Huۅ�������zK�Y�JKQ[(�٥�!C��T륔+F��6�����ڐ�uզ��Y]D6ұ�ջ9-�[��֑hߚv� ���UZY���ú�vHh�Թ�g5&�e�%��B���1��af�g������NS�� �@/��'�\Mӡ�dEa~������>�5�Pg!��N��ƴ�Y&�w[t�S��I>�}��|O�wzd�1 �7S��ʇ��O�Ƈt��.�$�{�ݑ �A���9�=`�u��O��K�oD��&�2%�'r�d�n�7w��@���$�v�� Z@��2Ŭѫ���}�pu���윤�Љ�� .��W��&�����A ���O�/��2O��M��!,��v�3j��zY������Xd��e�B4TŶ�d�44��C��a¬.�Òz����\�U>Ϗ���:���$	�#{�A|�VȦ��S�h���I>y��Lg5�I@�ȧ'ƹ�=����kh���m�ѹ�dS.�ͫ��2�-��N�.�yVOò�Ɵ?�;w�+�9&��2�:���:Vc�j�vl�2��eS^9#1��f����x��S���̙�D��ij���ϞȈq��k��9d��u2:��d�k� ������'�'��{D�����;�@���e�����ā%l�ԺvEV��Ǥ�ϹI#���7.�߶�(�y����2i�"Y�w,f|a��@z��Uu�7G@�9{�����|��q���H��N�Po��J�d��Iك�� RM�`m�t\k��(��AZ�Z����y���S���윤�Ё�^Lp�5�b����\�J��==�D���� ���- Z6-��:<�4���=�=��6�.�Is�G� O��@��'^�.�b_�����O��12���ȧ�E���$�<+���RmD1�%:g�qx�U����Ĝzm�k�f��;�ɄFa�:��qV��RS����3I���	ny���8���,��}i�X,� b	F��p>�� ����f��,�w	�:�U]3-�?]�[<�$�l�y)��>}���1h��9'���	����`]�H=�	$���H1%�d���Qd�4�()�dA�~q���� �hzC�6�A�����k�"�#n�T���U
)-�Ômy��e4.:v�8u��ᘖd���a��$��I>��n�6���;�5��S1�k2ע�!x��.��)��rΒb�L�v�� �ٓ,ٽ��x��Msۈ$����$`s�s[�N>;� |��0Nŋ��= ��3�J�@�h�=�B�Ce�}�� o-1��O�4����E8�u���ikb4w�8-SO��][���|I��q���nuDY��]Lnv�$������S�����3� ��؊ǆL�]��qy��A��W���Bof`�t��|��^#�U����w���i�p�73 AƼT僲N�3�Q"q�fI"߶ ѣ�k�kgW ���	��{��I�~؈s�%Qg'�l#�{����8J��v[(T�s�0e� l�x&c�"b˳j�0����-rg���o�8{�Ȑ	$��w5��nQ[�q��q�����$���ZӆbY���(O��m�&u�E��Y��Ǩ��A��t�d�[��X�'��nwI	)v)�vvgIr&m��gĒ>lA$�7�Y�KvxH$�m�O��}�7�nŉ�q���v��0�>Jo��×� ���A͛�$ͽY��,����3#�d���cE�A���@�WsSěm�S���=g���m�����y��m��z<�ށ ���oF�A��/��S�O�s�kx{���?ϭ�tU�)zŗ�&����2��'��-���*y9�yHOE;�����G�2`������\3�B��L�PvJ��t��î�n�R�L�/=mb�L�%f]Dq������
b�P���)e���5��F˵�P�X�����s�
T֢]�HA�V�Bݡ`�%�h��v[]jd �m.܅�����!�Mi�d��-�,1m�*�[eԚ!���u؈���wh4�#*j�1�[�챤έ��
A�&�2ʌfWk��>3����*�X�73�[knsЪbX[f*5,���س-WR徆��
����X�t��L��w������{�q I�%�Ѽ��j��輮��� �[s"_�����`]�H/���A���[Ck%glQ> ��r#�	�� u	��A�o�'�g��N�3̝�1"B~��A�x��K�X�=�O�ۤ���x�<N��23�+�wv(3�}m�Q5!	k�b� �zؿJ$���wzfG��P��e���-��K���h�L3�e�<�H����$ƛ�h����q�I>�ہ��s̀^#ֹY��=_�*��j� 3,%�2k0�ˢ��
Ѷ�9��1�]�vt�������0X��q�ȷ�1��A$��w�@=�te�V���`���?\�H$��� ��Z�;I;�Ν!1�=�}��y�����i
�T��7��<��`?/E�R�=-�Z��<(�+�����v�:{�aP?vý���y0��1���l6H:n����B�^$O��$��2$�z+.Z@;��d�t��.�&|Tg<	k�ȐA*^���֪^�U��|O����%���k�.16��1,Y�ә��������[D��|OG=�$�}��I��N�"v{�|.�!@$
v��1g,��3m�S$�������u�cp�t݋�ϛ�&��́��Q��׽Y*�+�(�	�0�W��+�������W��h�ڌL���9qSf��,�K�39u�Z���$�|̀$�^$��� ����fJ��C�V!�/w�$N���(3�D�򮋘 ���=[Ğ-m���C!G���$|[{#� ch�5�vDvfN%sr���T����ggP&��_L�I����=>n�<T��i��n�S��*�`M)���/sΝ��	�-U��~�o�M����Xj�cE�g|�j�:+Qlf���d*���uĞz��$��؃/�Ƈt��.�%,)�Υo*D=hiemô-��	`gtA ���*;���,��3�@�+���fZ��bX���3>���|G2���ovm~��Wp(����<O3g(ow�.���^;�v��=CXD��2	&�.�-��k���\��gc��m-�z�����W�"E��;s	����I#Y��U��*��dDvO���DO�WG��.����I�S�s�P��{Y�(�T���I� ג>�P�K�=��Jj�U<�����>X	Y�tPf)ĉ;oP �'��η��uG5)�F�� ��� �5�9'�ْ��:I�vtޙ��7�y��i�s1Ē)�y'���>���f���҈���܉{Uyn�o9T�2KA���o�ğ��wO}��^O=y;nSӧ��T��w>ں7� �{f��$��^���9w�e{b��.���d]�L�+�xA��ȝ�w�1U�7��I W�VDx�F3f� �u�zd3T�l��d���|&/��k����j�R��Y�sB1��V	M�.X�j�75���~m��3��p*7�	> k*� �	���Ses��F�H/E��Њ�ŀ噃�,����B�~z���O��5���6˭G����H4��6N�X��}�/���<��wd]ٝé�☆>'ǟ3�|}}��j�������ကF�oD�UcB+}I�q>�iC�~3а7h'�n��"|A-��C>�E'��/�c��'_�}��$΋;:�$�����Ι�ͨ3t��`H7 9��$�H-�������ab�2;D���G���6�D������#��ȻkyϗA��ʦ#�Z����
}�^~.B��dö�8� �0	0�'d΄�pB:��S!�R1��U���c� �ӱn������˞-������F0�ͺ
`�4ty5փeD[�q�6%-�q�K�M5������1elX�7JhJF�D�򅲐�͛h�qcA������&e��um�qE;\<Yf�6��f�`�u��b։�M��:Ys�2Ԫ���jE��[-H`k��f����M�pY�ةT�#�S:�Y���,c�0U`M+SV"]����'0��g�ws�
���|	���	 ��؏�0{Ui'���=�!y"@����҂�L�Yvwa2Tv����U�^�<�O��$�KolG���j�h�舼opO
�L]�dЦ����%�q���7�m�A
�LX�H-��D�Am�x�ӈۗN�Γ�u2[��wPs�TgCK��EGFD��@-Y� �H��Wm�u��sC$�w�nd(`Eg�"��N*A�Y��w<~��-4\;���\t��v@o@D�k�@�h3��(�WQD>��wpX��CMQĭnt&E��\�1�F8ͥ��t�l��u�OM�w�gE��p&޲d�
�k͐ �� ��#�憐l��a�fə�Hn�x�NIwN�	`��d��x�ᾏ=�:!i'�򩦫�j�f��2�:x�<����<V�ϗ�}'Y�����F����#5�E�庇�ϻ���b��	�Z�8�I/Y� ���I ���(>���y$�)��ıggv$(��$�͸�	$Ν�Dۄb��P��k�� �؊�@���<H��,_���JBf�:�9��d�����y$k�I!f�M溗u�׭�� �gG�#��6΋�w)�:�-���H+�:'�	�7qۂ�'#����#|���3�nV�����u���|��F�]�e`�ln��+.�ڂ�D���a��F٢�������Ov�lVq�{*"6����	��2u�ی�3�n�e�L��?����޸���fD��M�׊���ܩ���/ӂ$�}��zQ~}�I���L���h��hǚl'd��g�`��e��{����ݐ'�?�Ϯ���Y����������돏�������g����{=��g�ٞ�|ƕY$<х��C�*��	��ŷ|.�^�����r���.���i�x���{QL��k��l��C&����F]-J2��C�#g(]�	�;�+���#w<����'���[��R��)p��/����z?3�,9�О����=�)���=���xt��9/i��WTW���|�AD�Ť��.ק� ���ďZ��]��{ۗr�JzYށ��=�O��[��x��q,�e�u@$���ؐ��|�8���sႦ���\�!�m��k�	��=��؃��o�#���n$�ᗀ��%vU���=�.8�w-��$�У�V�uy�#
$���s�������N���2NΏ��gO��|�d��U滩k��&Y�������þ��jU�'l��+��G�iƀ�;N�G�=�Cܟ�,�ʕ�W�%��,l4��@=�R�f��I�Z�'��t���dv�� ���:�wڵ������g-�߼���t��y�0vn�0a�z{6C�i����Kݷ�R�G^7��}�u��S�t��{	e=����%��&�:��m�ǩ��N�=S��gs�/BԒZ�񺏣/�_@���צ���w�o��
h�9jɏ���x�z����
vĥ��ѯ��u�-��}�*)�(��h�'%�/D/���K��@�lB�oa���\D���噭u���1��y=�l塡r>���La���14dM�,�v-�
s���-윹i���2�p8˹.��H�S�u;$�0�|.��6�-�gu���vW���%m�r������e���m������^{��m��cX�{dQw�M���J٭�3��pwϋ�ӫ�O���ye�y�w�ٗee�!um���zwFf���0Q�u��9.˲���/<{$'ue�+J���n�閶�"nD�(��8��m����ӣ��ml����]��%�mƜDe��-���A���J�8�����2�k,��99l͛����gg�\�GghY�ֶ֝��Yd������xr{�d�S�3E\�γ����싈	 ����'�ґ�fv%�;;��$��0ky�&�$G��ׂA%�7�|O�%�8Vv�Q�χ�����l1gb� [v��>��؋����cmoP���v��C��L�m�{]yWq�,dP[�^�ɓCd]�,�]�b��u4KX�i����63K����\c:,�ܳ8v����>0c��� �|Z�<c��F�q��d�@�Ay����D�Pf)ĉ�\���T@��u��|H�ɐH$��s��n�6�0�r�OS�&[z��gfgt�;�������-y� �@�ۺ���=e���}�W� ��wlD��]����geV�;t�uh欲A|x�Io�mΙ�8���{P����磺���T)A�'܈�w�Z~������H钤��\��;��
jb���w	=:�[���lFz�A��1E�׵>bQ,�ıggv s77�#���ǅ&6(uOLH$���~(�w���1޺H{��C����:�(6���� ����k����MM+��cun�R�g����Fc8I9Y���A�6 ��}��֏*y�d�&���Y@^N��/[�7�Ni,-�2r�Y�;!Rv��	r��������$��A������;�$��:�� ��!c)�q�io=�o��Rh��b����V����= �}��	�̐�����;��i�)�;#��z��r�<@"ںݻ��@����nJ�΢OES���'(��g�"��=π	-��u�f6>��҃�}��@��m�O��woL�Dy�~��#�؁��eɿ�[�~�^޻���#�9м�vs^cKnIe8��2E�3r�9{aՇ�w�W��Q�^K����	�K�$�w�;W�����w\l��h|Ŀî���P��[m�lD����C4&irG3`W\�NX"�؊+b����SR[e��3LY`ׅBV�cK)c�˨�U.]V��KJ[D1�e�e�v�6Q����tK@k�4!L�lح@�q��Vb:L�u���V�8� 5��u�6������F�:\,ic�fˣ���J�YRb�Ͱ�Y�Ŵ,�4쌶gߺ�ך�b���Ӑ�m���v�E!��Һ��74YMr����ϒ����eͬY�݄�TU���\��>$-۽�z��;�y��s��l�*��v)!m�3$��Aٵ�eGG=O���r$ϐE���o��������:�A�U����'.�ô�'na��KvgD��N[�2�P����M�A�/�����w�NN�5�JD��S�k����QQ��V�\�O��k�۝^H���rLsF䀈��R݀S�L�ܳ;��O=l�Ak�|w�WJ�ӕp�C
��Al���Q$;v�w�mOm�"	h_!�|���P���S[sIuP�0������9�����R/��r�:N>�bw�y �[7�$���$6���V�{���z!��Ǭ��}�����4	��[�3���G�ۡV��?c��I�Ɉl��M��ȑ���{-�a�ï�����3���Z��w��>T�}�E/�}������lF��p�d�-&�Dv�-������fn����5�p��I �=�\�$ݼ�O�����H��v(� =�D��Kwl Eh8-:d�ݓ8w���{�Z�2�N���dnoTI;� O���I����I̽s���,�2O���ZR%b�H�Z�	&�yŴ�Y[PJ���Z� @ �l�K�I�R������ׂ����Հf��5q��[��0�P�%vmɐ�ir�'�}��ngs�w���d	-}���Ͻ	�~��.9���MH%�1�_��.����3� ���$�������dh$��H.~�d��o�x�����7N��S��U�T��ؖ,���TZ7c�$�n<�O��~�V&A�[��m�q����S����䷦��bS w�NL�y�R���!�"�fH�o/��׃���<���x��Gc��VAm<�I��^k�Ijވ����@$P�`�8b��$&i�fN�.�S"���o�=��>������n�u�[�׵{��=&A���?gQa�S�����u�(��tIf�WF.����u�1H[9�x�A#���>,�jawW2��"�zeю�i`Z!NJ���e�D�%m�6�1M�K2��u�#X�
�qÁ�z�$�lׂH���rK\�썪�*��W�/�G��2����)�M�s���� ����.yD1��c}!�z� ��[� �tS���{�߉�,�ӆ%3�1�Lݯ���� �Ǳ�J�k5�ӰO����5��d�m�R���1��̃Ͻ9�Z�w��Wad�x��׏	y]�2H$���G��ʎV�(B #g$IDo�{ �M�����sG��MMZ|���;��'�v�flC����}/E��3�ˍˍ�7���G��F�g 9�F�{��hޗ�lde�2)�8���+b�Ĺdؤ�ވ��؀:6��9��`@cc׏�S�l��^Ǆ&����bvx��A�B�� �R�m�N2&ɮ���]�h���mHV]�WD�S��i�T]s������!6gD����4@'6�S`d�<p������`%�vd�r��e�E8�R� �o{�����S��o�dm��$���u'�3�;ke�5�?\�Xe �M�.~׿�/�~� ���.������(}Mٲ�I �v���YӧK3�T�:Y^;'p�x�L����H%�� �9��0]�xn{1�޶���MZ�AM�����w�` �p�֓-z�_�c��x��[�{�9���Gx�ZQ��L�9��~���&�Z����eT�U��SJY ڦ��2ʹ"�%�x��>	Y�E�����9N�ϼ�	�8�E�_�h�nZ�*�Utں�躜4�k�� ��" �3)	��d͵��)]Rb�S���������t4B钸jJ���D��:��3+���%b�l�@ E�����-�nV����.���ë ���e��48&��{*��0m����[I�0D��6�٥�J�t�I��xl.1t7l�,s��e�M\��6��۹٨[��詋�f���6�c��J���9�:Ql� ����O^��B��r�3�Ewx+왐H5��Y��#Ŷ��i�E]�̂$�^�Eh9E;t�ɜ;̞����U��<��i9vِ/���@:ݮ ǎ@�䩅3�Yۋu���gA�F1�D�a�RTm�� �Z��� #�N�u�؎�j���KV��� �z�	9t�]�;�oL�Lt�v���n�':�	��� �nޞ�H�H7�y��VdD�'$��N�g/2a�_�&ۻ )ޖ�c���û��68,�� �9� �N6�H���Ҭ�ށ}mvmsSF\�MIt�mt���5J�6H\��]t�ҵ�u:��'��NQ#���ڪ6=�-�x�%ͻ� ˱���7S1��$����3EX� ��fD�����ׁx�?��7��c����ͫ��폐֓{��ǳ=zv�H�Puk�Q8a�}*|�"{�y����	���X�ʮmTT��D�0�����O�^���@s��� �d3n[��d5f�Nh;e;t�ɝ����x�y�r$��t�j�#v�s�ʺ�A���I#w�|H��t���)�)ĉ����:Ry����秀}Mw�$���S0��|/�7s�ކ&;*$B���0w	��r� ��:��h����L�-�GAع�A���	+��F�n�>���E�=.`�'���+��PP�kn�Z��Dڣ4{�|a���=�h���>�?~>@���ؒ����s�6+w_�`k�@$[U�D���A��0��v,��K���z�|p�ȐO� ��i��w+��ā��U�]2�QFMs�`'ĕٱ�����Jv���2w�l����Fҧ���yl}�2[�`�>.1r���k�P�Ӕةԉ���lA�y��9��@ݢo��5\;���y���I��!�I�,�YӧL�^Es;較���0Y�'��$xډ$Y���wk��9v��Y7:'�� �׺�9\�T_�1E8�>=oO����W���7�����H$M}��˛��o�b�R�.�V�.aڳiv�]��(,����$��f��sF]4+X��H9|��Y�3�N���ڌ��H m���^d	�l-�UM��=��Q]�	:��\�K'ܔ;�I��q �vX�15R�D�}��O�O\A��E#��L��A ]�dm�ɜ;;@�.�� �|T�F�̮�6��UY@ߊ7l@$�wlz ��*�.̃;�Q�Uѳ�xP��nJU�#� HYV�$�wl����1N�+e����H׎��}�kgR����^���\��y����Ώ�˄��c����<GJꉜ2��enػYJ�t1������3��{��� 
��|���h&Ca4�����[;`t��<o;o�j���A�HS{ F7v��)�4w6��A�_gVc�Tv�V5��S!��Wh4��t�k3R�;<n�s�k�3l��ߵ��ܤ@��ܳ��ߜ��\@$��׳$�C(�i�S�ǯ�y����;���?z��$�h�÷��:�I ��(��s�B'<ݑ�@$�����:�����!��[9�N�(2wi���'|�?gG��W��X�^�@�6k�M���u�!�8!�3�goL���K�s������sL"�n�$9���
���S�]\[žq[��=�X�����QFd+�ɐK�#ϛC�{�]�C=>��y�:d��������<6���������������ۦ||||||||z||q������מmO�g�s����h�B��c;_q���h�[�B�=:�M�v��F�%:����x��z���b,���~�V1%���b�dK}܂�:M���j+�= �/jX�E���7Y�ø�@�O��mt�\}=�sw5Oo�^����7/�v]G,f�k�"r�p�ɬln�k^�K�_n�"�g�_�P8���q-ot��S�Rs���np�Psڰ��N`�IO,�h��zi������z�~�Pu�t&��ZWY�^�{��;ws�QC�+�H'v�'��:�jg�����B�x��7;�D����z�X-l���ƞ�Y���e5�A�=$�g�>g�wڳX|�| �3�����5iM^,�S��y�Q}㺽�����~o�t#7nw��Uݘ�}��7m��VN�ȁV���^U�
��%���Op���5z�Ղ^��蚅l,��t읠K�W|� ��r��d<��9��X,ۺs��s�{(�=Z�q��G��z�g?k��*���oV����W�żW:eޤ�v\�Y]ឧ���S����/��4�}ݞ�p��e�5��?d$�Ovzks�����m���}�0<U%�6/e���>���w�S?o�;�/d�8��=�d��������9=NI$��~˓�'�惸���Rw{L'�]ٽ0B��>K6A�y+{���S����iFcUؼ�QYw���w�C)<L\b�ej%��F�oq�}�69����fȇ�ZT@��L�u�tA_�rq9e�Ŵ�}��ͭ���e�M��Y���D٘��"�8-�m�C��ަl�8���3YY��gx�-�����&�m�.m�Xs+C�>�x�O��.&ͻkv�3���klm�l�V6�f��=�<li�gm���{�X�M�l������"Nη�9voh�.�X�8��8���zD�y����kw�ie:>պ$���k�"�{W��ݵ�vu�[k[rKih��qe�˰�-#����<ֲi� ft��3��Mii��S%����m��e�t�ݎ82�[�s��U�����[c ���K���5����f����Ѭ�J�Ŷ[[:�}��#����ۖ�a�ge{`�;n�!8���vՖYH[V��3���s�|��^^�&C�m����\]oL�	֋�AtvZs[�.	n��[sږ�n��ma��V�JHT �V9���Ȫ��SS6J�6ؖYL�bL�8#k�V�!M���un��"&%)h�f^0���-�	���#��5s�d�E�e1�p�g��J��.�倷8^6��� ���0L6ٜMIEM��i]��E�vc)26k�b�*7�i�,+��J�9��í��l3�J$\T�\�C[�l�<k5k��[M�L$�.0�Uv��KG��an2�kÇ�XJL�
��D�6fܪ�L	��Qp2���iθ�4L��#be�Ժl�Q�kYf�U�լ���l�^�v�Z�ټ%��]te�å��9�\�h7!�ku,-�w0���p�F�8bi�m��0\I��35qo2��K��5���j��]��RY�Ä��u]^�з\��].5
���6�WWVWZF��Q�fJͫ���b�e���YL�N:�^gYM.��-W.fc
1l�M����j�ڎ��Eb8!6�%����KF�m�Љ�m�!�e&u�/	G���$�K+13q	�i�+�f��#��h�0�ĬN��,��&�-�,.�4l�I���N	tH`��&nx-��7MQ(�n�IKc`���댉��\XnDul��ˋJcS.��^��f��X��^� 4����&�7�[@�YZ�$]��1w�K�X]QҬ^�eH2�ׯ�F�`�%f�طd\�%ұvFlԔY�4�&��2˛VVff��6��[v�th,��m%h��*목Mc�!��ŮS�5N]\���3��� ݵ)CB6�[l����4��ە��]������m���v�٢��a����Ŗ"�R�"%4��a.�� %y�]� ��(�r�n��(�9�;0	ucP��]�`�GF[��T�[q2�cY�gmb�Z�ע��t^��inWla��u ����b������P�xx�ݩa���l.X�.��$�a�\\�]�.�u�SU�"-��A��Pm2�2��.��3Z�q�������j�e��2�����υ�5!st����H�f��[6��巖=3.�Si�M��u�M3�j(��KR�̼tF]3i����XċQ�d�)l��D�e�4,Ԍ2�#t��$�V�\�CCC8e�n�i���f���U����}��{�ɤ��Z�V�]��TL�ҭ�$�&��&�L��r�~�\Wj����s�F��}����$~��;
�N�R��}�O&��ɔ<���KjtAA�N'�m7�h�2m��]�/�pA���`�7c��d�d����g<H��iL0wt��y]���o� A ��'k���� �H��z�g|�+�ˡ� ���N�(2t�%G75j<յL����]oD��|ױ$��ϥ�m�>ʦW^e3wQ'�a&Ėd���K6s�<�� -�����=4��ސ-wW�	�k���j�'�k&:�ԭ�[Վ1*��c<��3Z�F���&I�f���Z�PL���<3�I?��E�#f@>�[5���`�b�t�M:>��׳$�x��'����N��O[�B W�׭ٱ/�"���W�87�Q}�^�{õ�~��L���ܘkxS�]�F���Z^ޕ<�<���Տo����l=��[�܋���kܡ���H���$�?C��6�-���#^Woф���Ś�"Pd��vޞ<E��@GĒ�*�\������D�vI���B�@��6�Z�0L���N��Dtu�I�pL+�lh5�� ���� �A-��0����u/�8��뉈�9�zY8.����/ͦ�k�ؓ��^�-X G����� �&����d�=]Q�7�/9�)E��Nɋ�)�d���m���p��a��֘	v��s�gߧ�N�Jfg���Y��	<Տ �|���d��ju��k���S�@�@i��S���Q�Ttl��$OV2���l�D{*6D���D��;��d��c�`��d�tYû��^F5�� �����>�y���'�� �U�F���4l�y�ǯ�ǃ����ӳn����z��ǖ��$�ZW�܋|&~��h֧��m��b�V��d��vV�Ʃy~ �y��Nll����'t�f��$�=�ӷ��S�aߪ�$��B ��By��O�����(�F�7Ǣ����Έִ�3wI;��@T��L��H1�z�gbnjD�@�H/=�>$�v�Ep{���IjG����a�o6s%mq.��)q��b��i���,�5]=O����s�AN��VO<w�@�nLH>#������x���!/6^wd�$�e� ��2eh����'h��w��S3z��m{#<��zOoL��M7l@&c�L�c��t)�]�(ċl��$�l�{�mJ���}o�� �^s:g��ߕy�:f{�l[:,��v/3��p뚭�h�&�<��evĐM5���� W�Պ�cĉ3�
nLZ��ZM�Yy��x-�%��r�ESc��k��ws��1����2뿒+�o�#�1qӗ׽K�ꗒ��nډ��,���$�H�zޜ_���s���Srh�E�L̐|y�"6�{�{���|�z}������l3q.0�*��l�4�	��̤m"f9u�.��v^��{9�&�wu��r8q��Ѻ�uJ��<�15ܷvL��'v �r9,�K�)�vy�y�v$�r��+z���.f���A>���I#��0�����*jq�����L�S38d�9��w؁�z�$fJ�g?LF�sj{Fx�5�z$��tz�؊>E?��E�g،�[x���2�7�0 ��H�|� �O�7�{m��u8/�`w:���'3��Μ'r�(s�>A}{��ߪ��Gf�7A6���O���A 7�@ѝ"\���t�5�ݬw%W�75Mօ�G�P�gh��{r�!�c\���˪O�iz.��2������ �����LV�HF��O���>��B�ѵee��&�2�0�-Z*;�,�+meI4�L�cu�"V�͢����i�A�m�Lh�F�-�P�e7	�W��5u�
0kx�kk3��v�6V�����,%�U.iV֑.	�p�^�˭LT�͡F���.�A�B�1-���ݜpR]L���T��6+���h-M����3f�[.��3p��
�ڵ]e9�:�
�D����1,0J�ElSk�+.�����Bevƥ˒y�ϵ��B� i���w�	&�u׌x�B��-�"�0�7$�t@�m�	�k0d�ݒN�U/�� �_��1�.�D[8X�"	 ��5dH$��۽�$��g@O��M�e�k��nи��Ħ)��L�l׀O�8����7������-k���Y>'�6 =ױ��p���%��ˤ� ���u�{F���:�<	 ���$�u�OH���m`����	��^d�0*��:d	 �f�(~���xOnL�D�gL����E��=��s�/P�8��aq��.��*M�J�+6���è�LJh#�vPUi.wIݝ�'r��9��׻$�u�fA���v����� �[nd�9Y��58D��'$��<y��+��J&���fY�V����K�B��O���E�;۹����p*���5߷5cV�?g%�/���.�1�Lڌ�feܞd��I>$[gt�$�n��
���\�]'����pR�]�$��@5��q�	�ƽ�Ă�al��C���=��ol� �k�O6\ �Jb��g�Gs��������Kx�~�I>��������A7̩əغO2�L��>$��x3L�kU�*u��3 n�ԍ���3|���ѓX�O��?y�ì�g�]l�u�(b�m��Z��."=UK[���&4�	v{��p�y�7.D���ْI��͈��ot{�*o�����y�/�PcnD�ғ[靜3�y�k� �V��X".�� h'Ā���
���xݣOV�D��S��K�PLRq"@;oQ �}� ��W���g:���ߖj�w��	ʺ�)+�x�v��w۾�k�@ΝٷM�ݒ�\h��edŵD�Q����/+S�{�WC"̄�z���4��p$�O��q���Kh�K3pX;��枃8^+F��޿.���O��H'˷:[�j϶���s��*��Í P-;pE��H$�����pt��|�\	�qG��#�	Y�� ��"/����:���P�f�J���[6�H�pi�G"�j;Xұ@.�[Z�:����}W�Qspk?{*����l��A$��wkȮhXkF1��O����s�G�gO� S���]�!yp~�ʪ�}� �������dO�|�dKQj�WOs�s�;�M�S�Nᝃ̚���|k�6�tH'���gL\��� �_@�I;:D���Z��(&)8��3�wݺ6�Vh$x�W8�	�K���T �������%�f�0�?��j��7={�T�U����y<Z�g���y�@.l�C�`���z��w�ŷ���n�v�p-���o�e�p�gj�a��ű2Y����ݓ��莙�m�`D�l�9�1�c9ƀ{�퍙�u�`z)�m�^���l���E��+����Ž�Bl5��f�l��4)��H��`��*�"k�N��rS��7|Z[���sr(O?k�ֽ����Y��b�Un��)�?�gb�<�)�^���60;U��Iw�D�A��O�P�}�X�(>��*٧E�c����Θ���5~�詐	$��D{T^���{M;N'������ɒ	��=n�̬3�ft���U����{zg�UB�D��ē�H��؂A!O?�x~��\�3[T���"��1iw����}���B�n/�Ph�>$�����@ ���`�>ߧ��26�c���WpP_�P������v]�A��)�o�̽�&rC�_opNˋ�ρ����;]G���ir�E<`��jx�$g�8�k�˯iG����+���%v��jK�ĸF��6o���PJ����YnE/1���:����< `3��V�]f��ӍSM*r�fC$�#&�3;��Bњ�5���G慆 3r�f�L�����5ᢸ��<F��af �0�idB$�+3���u6k3L���u^�YeU�q6���2��X��7Y�3B\(4sn2ص�)�RĲ�ڡbi�G`&@��ɣ�X�j�u�d�*k����itТ�?�'�a����v]�k�H�D���3g�{�����[p��Uꮙ�>$��Dz�g�Jb���u܁�=[�����ױA��M��$�n��A��|�nC�6��6�&��LY����́\���zl"�z4�6у�^��h�@R����"�?�1A�M�2j,���Y�5�oŌ��B��G�n�D���]�y��rN=\z;��R=���)�w7�3��/ޟ��H2�z"��i��A>\�j	wg@�<�c%�`�KzI�đ*�����ᎺnbڦcEe�����Y������nw*�M�w�v�0%Įl�|O���b	0f�����qx��o:b	ٯ��qL����we3���$��7�����Z�-�z��^�L����wyD�2��������5H'�_.�$��a�s2��r�6�>D8��]���0LwU���q�Z�>�L���D�.๩M7�х�g1vg��N�����H$�՗���r��>�f(���Ι����L�������L�z�z�bǈn���N�a��$^��dH:��wLD�$v6b,t�6�)����gLρ$�|�nʦV3���v4RK_nL���~�u��M�n~w�r�Q��%6�D$k�� K.R:�Lך3&�6 j�ԙ�u-���K�p��N_��g�>$��ؐH$u�`\��s�n�﷚�A��ݻ3>$d�-N���O��l@�j��ū"��s��B�6gĂv��ץ�BΪ�2�v�k/�9Lɝ�`��j,�	�]�������O�C�O�ooooo�����g����z���/g����y������>�٥p9�v�;�^�N�\<6�==�K���.ص�Uw{w7A<}�Eֹ{�t��I&燹�Hs�7����$:�~�]����w�A���lUWݻ��-�~�ܝѾM2�p^�r7} ��/���|y_��;O����b�/u�2z_$�r��\=��BoM�h;������wӸ��N�i��"����sɞ���Xlۨ>v����b�P��8��H������a���8)0w����z��B���꺯����;N=^�A�<3s��P�O�(b͛��|�%���l�/���3Y��S�DS���V�J�Lª鬝��`����{t��d�}����k�6k��޽���=���&�<i����+�C�S;﮾w�4]x��f�Ά����^��7��������d��wY/����p��^�;�������	�=͔��.��цt�s���9�x����2�U��'/�O4I��a�p����+���$X}�۸�Vynk��<21^x4�n�Z�y �9��=OO������!�����B{B��}���BD%�nkF���=�/!p�H^�m}B�;3��e����}��XWӹ�|9�l�ǉ�l��rŽ����������=U�`���t;js}����ŝ��)�������;�G���w�n�����x�8e�ƈc䤽.�.-��X�G�1W[v���!d����A�X3�d�\5멕�\�T��W4s�~��@�������a�ō�޷�>8PI1�}dH@�Q�ĕ�/0ͳnf��Ƕ��fċ�maBض�6֚���%��ힸ�����nf�l���yv�6f[ni��n�6F�kY�+A%�����,�=�s��Nvm��I�9�3o{�6݆�6��d�ޛVm�XƑm��H�hm��ֽ6٦��f�l���۲��#��{��9,/:޴r]�q�v��1�3�6��k-�6m�s�����H��of��N%����YEe�/=�����h�����\��Մ�fG-����f�r{f����M�ݛ�E��kNI#��Z���y�6ݣh�Ng5��8lk2���N��qv�o.�F�Vmf�f��6�osmm�6�2��7�瞵� �N�m�۬@��;Y���Lֻ[���b���[��kkm���i�[�I�)y����a�5�t3�Qso���{N�ֵ��+���؃O���8L]��|S�t�����*������	
��A>���չy�O�g�=�o���1�\_�bMK��g@�I�Ƹ6{:����ݿ&7vgă~I���u���ޔ#��7y�L3k�o1ڱ+t�b�1�"�tR�0Ʋ�B�1�F5�@ƴK�΄3� 9āO�f"`�ᱳ�>$|�M������u��5w�Y��d	�]y�+F�"�32N������`.w2��ǃ�Q ���^�;�@�@��� �C�i�A>��E���5;��C� Z�q�nn�">&�j[�ˬz����$����~}0	jш�fL�vS��PV�W&���\�A$�[��W��� '9���)R��	׋��U\�DeC8�h4��둉2��?E��q�@y��z��}+fK��>�w�K��o�ix��l� �9�>8�v �v(0p��3̂��`"I�{���˨v�@���L��l}1�>@�Dtό]��z}�0�3$t;eH���&������l�*��K�C2�M����-�w�mv2��f���y���$lk�#���Lz��[�6��=?����phl�6Q)���̅�2H9�n�b�� >ڙ܇���d�@�~� ��kK�j�~ɸ�����gL̓�/[�����bA�{*�1��uݲH2��`��ގ�v����r^`�H�Z��s-�AUM��$���Hwn����}�����`�PЄ�L�vQ8��"}K�������.�U�.��ǈ3��2>+�b �^+����N4�����x�ڌ���W�읕�7��{5L��9sƘ���'&�SKJI�B6�)A��Ơ��B�v<s��������X�Q�043Xm-
�a��ɶ4[-�%c�&������w�w�|!�<	���Ȋ�R��/)�l4Ÿ1m1�bD�#5�m����j��-�Ҙ˦-%]h�	���"�Mv�f��lKlt�L� �և9i#��$��/"ulB�r��	�.�k.٥uSq{2ʵ3\�;Y`��e6X �f�ǀ��a@��P,4��:��8B�`U�^�J��!��U�(�*i�,b�`�\��u�W;8L]���|E�B ���� �H'˻byN�@���l[�ɂ�{3�DWC!O�A3�t��A]��~0溩,��O�fͻO|G{�D��@+�\A�'J����!�Ŝl��u�J'`B2rߣ	�!�vl����OA�չ�H=�yI%wlAz1��0d��w��kh�3���CB�O�~I�/"I$ۏ�F�||�e����]S ��\������\K&�*< �H7��Y���\�F��"�΍^fO���̈���`�F�3�D��yޡM.5���ƭ�.�㮙��ݝ@ͫL�R�77E��
l�yvq���m[G�������̀}ĂG����6�*�9�o'+�e<��A��>Q�ؠ��b��d�-��3�άk{�GTg<4
$�X��3�6��+x(���憐qF�I����o����_֣�^iy�����}ަc�UӤ2BI��z��s1/䀏%^�ޙ �;�A���[`��5鰶+�8O�VC!O�A2p�4�fވ�k�I/m[:]�L�W9���b��%��M{� �O����&C�I�������a��Ƚ�R�dx�i���D�/�#��<����s�~H_q�O�]�x/B�^�M�t�2p�A[��<I�~ؐy��*�v�V�LF�%Y�	�q����a���~�;��؎H̹���5!�T�k��T�Z3M��5�k���.\�������RS�t�9�PH;��!��Ύ�㍩*�~6��嗕0�=����2Y;�b��?�G=tϦޢ�C���M<��� Gc�$3��d^�O>Иa�q����5��ؠ��d��d�O<I �=�O��$���0!���&��/wE��<���l��8fP�jMF�++�hլ�W��
�ߵ�'��ťJ�r��ϻ�>eQqm6����B��vx��mÁ�{qg?tJ�Q��Q�d��i��ۖ��DE��:���q����>$ⷳ�i�!\�`��t� '�I����ϗ\t�'�����f*�`p�f~�m�O�^�@�.��d�O��d�5�S^�5p�� �RŊ!�"�'%�ZJ6S;�l�i��ͥ�B���.m�4���׾�(}bp;����-�Sm�A �N�I �c�V"���jr��c��˩	$fWt�>WV��L���\T�G���ů%��a�m���ć�3VWd�$�n�V�d�}.��_;�/��d��;��$-��>�#�A�� �ɢz��p	��H'�չ2	$�v�{i�6;:,���|�~X�5��kj��@ϧ��hI�?l����¼�Rs���ڹ
����y`i^&��.-�SĻ��c��Ʒ�Ӟ2.AUY��+$�nf�����'U��[�k]pq���&w ��x�p�4H)�az ��<��ÚP�yɸ@�|Sw@�*�q�sQ�M������.լ��*�fm��S.���\��b�Ŗ��tࠐ.�I�M��Gu[��>+s^	�Wt ��b�q�)��/��,+��A]�ka�&�9i�N��I11tDw9N{���̸	-�ȟ/$HU�	��?g0�P��£�2�PH�b�Z��1���D	�2� �]e�?�>5�x7��wt �B��J��<F��M�6����u�v)=�,"�� \�� �" $�龝�m���wW�f]��s�2-;pF�<A'�o�N�M4�9�rⷲ���Ov\@'ĭ́�=� ��w�ٯ#������S��u(��K������`&�f�YJ�d������;<�m��/;�
�;���T��s�^��E^�prihe]�M��M��)�5n#G��5:�+
J,kL
�C)�l�L�`��&Rs�KQe��JEDt�&a0�IJ9��T#!&hUZ�cDW:���7�JƌYq*ۈL<l6�)m�u3d93m�ǰt�5$��Aa-�]Φ�E*tR8�Ե��]LGALe��@h6mf�q�� YX�AWEe�v���L&5O<x��mve�5�h�Zit�聦s�@�v��Tl��V�B�V�m����N&��fہ �9�<�>%t�H���)�T�m�1|�ą9� ��KMRo`B3��	�|�~�h:�&c*�ށ
s�@�6�k�$�u�}o�U�{t����z�^&��'E�3N� ��<	7�� ���瘱���������3g�dS�Cg)��q"A�z�\������7�1>0Qo.��$J��w����� �:C_��,���;��];s'�������xIp �H��2H$��A����;5���F��We�	��tk�f�el� �4qtt.#M�,Ҽ�妇ߟ��0��A�ڬ�<����@�9�$�I�7s@��1s�5q�ۘ��Iq�3�D�}�oW�'�HK���#��>���0��G4X�X���0�L�`j����GkLc�D��*�5T���|3�榿(9X*�T�
�j�j�7W����p�Ǹ�K��gc2=>+{�<2�R���@�k	����I&�g%�P�32 ��x$�|�Rc��v��A��I"�/�A>$��>��L�h��b�ò��~sR��2}W�[�d��������������v�t�7H�$��A��ʝ�E �\@���I]���%���!�d����QQ>+�Ȃ��|Hnȁ ��1��,����Z���Mf1	�B6��)����kfo1�A乗B��P���	dp�wgr��wi˙�J���|J��q���r}|jV`�|�I� ��#��dP`]�)�GA�v ��ɒ4A,�5�Q^$I���W�n�q ��xN���:��(}4_�����ä��A�u� H��AFtZ���lk��B��l�UW�L�&��s���v7V)���yp��ww�+"��ȼ3���o�Kr�^5�z��h[5�I� t��^d۝�>[��<W_8�;H锑M��J3#��78��\��㭲��I[�$�����y���� ެ�De�fkE�vd�;(�i����ؐeT�71Ĉ����7�x����x��!�«�_D9ٻ}�y��p�ɣ���G�.���YM��j�B��2���ձ���']wj����)Bf���޽@��J������>1�k�:z������@$����y ��N#D�gw.��So^L�A~�TV��� ��}� {�z$���mc��]y[Z�̊�E;��zBl�x��	fOD�I1���^�ַ��ͣS��<H$v��g���I��I�K7t��Y�Ɔ{���H����$V�p�z<�w��>;�L!D�]�6k"f"\ƣ9�xi�x(�/,��9�3�Zix��g}�_���[�N���d���C봘����Lt��}B�K$Sx���z1�:/؁�" �MPՎLQ$]�t�� �mlH�J���L9���9D�K��LS�����
-����6�LhjFl����Ƨ����]����&p�����A&�k H ��� wѣ��[�:�= *��gƧ80d�a��q|k��<uޚy��p�r��<Hoe�uQ �
��A�y�eA�����-�*@�gw.��N��Y$���=�v����J�%v�Kp����d�I]���kP1�A�v(�y�a��6����@=�}�$��|� �H]����Tr��C��̒k�����I�U~؃�|Wn8C�FL����Bd�r�o�ppM�o�}���_��~j�(�~�TD����G�`���E3�����&ٸ��@�0���
,��2���(,�+2��!*,�+2��(�,0"̨�,!,ʋ2���(,0"�(�,�+!,�+0"̨�(,�+2��(�,ʋ!,�L��L���,�̬�HJ̤��,��,�̬��4�̤�̤��,�̤��4�L��L��̤���́�03032�2�0��03)0�0�0303)q���̬�L�̬���̤�� L�L��L��L��̤��̤���L��̬�L!00ʳ)2�)0�2�0�2��3+0303+2�+2�+2��$��,�̬�̬�L,��,0#032�)2�0�0�)"L��L���!2�+03)2��$�L��(C��s���C"!�2 �
�*�0�� C*�2 `�ʫ�0 � C((2�� C�
�(�����C
��C*�2�� C(��;C��C(0�ȀC(�0�� C�� � C �2����ʫ�2�탴; �2��8©� J��,0��",2��
,9,ʋ0"̨�,0
̨�(,�+����Û����0
�����A�{��������wT�?���?������/�͏��{lԙ����ݿ���䨢�����?�~� @W��QE����� r~��e���ϓ�C�
(�����k��yd����'A����N�>��}밯�
� �
� *�*�$ *ʀ�� (*ʫ� J$(� B$�"J�(H�J��� ��(*���""��"�����'�AhPD�@(
D�g�t߷�}�_�(=���� ��G���QE�?,��ɿ�>_��c~���R>�?�?o����}B�(�����'���;�TQ_�"�+�?Zq�����gf����� ��	EE�~�ژ�u�Ñ�?y�<��|�Mϖě�O��ɱ�p(��>���������qEW��'�m�w��3�ϖ���7�A����	?����>�QE|;����c�?`��+���!����B�GD����;O߁�w����ﰓ���(�	�E'OGޘ���p>}A�ǧk���P~c����������@�>����
�2�̓p)���� ���9�>��.                                       �P  �*� 
�H�
}�B�((P
 �@ %  օ���   +@�                                    �          �F ��� �� �MڃNl
 �@s���d �� 4E<   `y :2 ����!�l<�ɥR�:��(�)t� 8�@e���K1���B��:��e9��R�K�LJZ�N   �        j��2irʥ$\�
N���RY��){x hP�3K�ҩ"�hW��QE�PYW�B�]8 B�Y�E ��(@    tQf�0  �
e��@4��  ���@ $ �@�P�           L�=@8���ٜؐ�˙��. �����*�3Wi�R�j�u�.�4,� :�J�e�hU�R��A��  ���
����t��� vRPͥ"�s�ֳb�Yu��c�WZ��� ��Nm:�jW;��UNl�CF��)֖���
H<  ��      �z,�Z9ڮ��sjf6��Zl� R�17J��:����S�35�R�WW �*��v;[T��u\ 1 	Q� T ;�O;]��Fq4I�n :�qa��\��X�m������tuJˀ �T�mͪ��Xt�]LnZ�8���U'�HU�@          xz��l;KU�vv�a�2gC�38 �K��ڐ���j��N�s�8 :�M\��۶�4$ ��  A�P� =2@` @�tf��� Հ= u!��� �&.�x����Df�����2JT��4 �x�� "{R���� 4 j��&T�A�F�i �)J��F ��|��92	�i*4�w�l�2�\+	�e�@�$�����H@�nB		�@�$��H@��B���D6��R�1|j+��Tz0�7e���:�.���f^�B��vtѝu������p��L�r��u쓮�&�[콗��a���K��wA�{"A��/˷,Ht�((�1���ob=��1�d��L��n��3Y�N=�p{��hW�/[ǇQ�:��x
�N��۰���0��a�խD�J͡���8c�ϗ^$n��R�	�stuq��ߵ�Bڑ0�{�pL�iX"Un!"�eٶݲ=�2c=��CgK�@ˊ꜡Y����"n�Aqv�uCp�{�����B��7P;Ϝ�Wې���C(���C�P0�tU�@
��80�@�6R��GD ��Z�M����9aw��%-��=:µ�������L�0��9ҩ�N	����jX��͍����哯�;#�ۥ�{��P���;�H�D�7�}�#4<F��������7@����,�ɵlKOgs�&�nO$\;��oK���#���E���k&���8AQ8��X2�{dٓ6�pe$u�-(�9���U�ovظdY�wۓwv��11٫�)܍p�q����ś&m�O���5Q_&g�"��[0�oR�YztgT7[}w�ͩ�j8�ҵ�Q���O�:r�6�Ԗrݏ:h"ߖ�zI; aA��1���	�;�X�YlW+>��Ż���U���^wx����x��4L�7ѧ-\_�Myc��]�A;�����sy�w�]�;�DC]�q=5� ��,�Fj�Jc-mK��Vg5ufƨB�Ƌ��	��n:�8�nr�h=@�s
�9V/'0a��yGP)��Tw۸ W�ط����N]��F������uִ�b�V�e��oY��Ε���%s�8,9՗~n=�ϮL��r�h�{"Z�S7;42�{�6�˼r�;�-��N���2E�#+)��KGY��yz�rý�G��v�Bv�*���f�kwuU=�sܻ�9ɜd����V�xC� Z��{�Z0�Hj�Ь^Ә"hqʣW��9\w^��#4Ijv�����o�ap&�/�"*(j����5��~��	�7����s9\vdX[|�:5.���p�)+;��{�c��vp�Ԟp��¦�*�.�n�m�L��a'{�7_|�
�%.�r��xf� ton��������	P�"���4�:L�eZќ�����'ԥ](�Ylɳ���eJ�>�.�;�[��M�6�X�@0�m΃�6I�L��:a��z�H��:���V���^��:�n<�L�M�r�]��n1oUqɄ,/�sk9���G���h8SL[;	��b��{��f����흈W�
����T$�B'd�s�prC��TCOs_={����ŏd*�+��;L4�ۼ�=[Z�4���q��U�='+yn�qɗ�]΢�>��np����t���S�{�R�v�S����;�"��ɰ./6{�hN��A���!Y�k�[qk{q��Uq\�:�Z���ފ9nqܵ��6��/��H�H���s��X ���/4'j۸ŵ+�͛���:=-��w	^�y��i(�y+��E�f;����� xi9Vo,�VoK� �q������,������`�o^3�)�r���'^Hp�46���f�{B��VqIq�Ml�l
����u�������s��D�V�YqL	���Vw������\���#�p�S�ǫ�;�L f�~���$S��>������M�x޼�R���5����Uc�-��#s6�Z��*{:�Ѣv�}��;�5r�ܔu��f��`�],T��)��8��RF����	;�!\��X��\��&p���D�o-;�:O�G-���ˁ��,K�����^�Tpq�u�%�{t.38���x�w[� 3�}�o�S����p�9=n���g�S̲���<�G*�ӷ�<61~�,Y\��V��`��(,�Ƀ�gI_%��{��N�]ak����n��e�E4�.!�6�bG�22���:�P��Č�ȼ`ԛ��mFA�L�o]8{uv�& ��Wm呦���À�aI���:��t�;�ػ�%R�l�k�Z���gv=Ҳ��*�.�!����'F����;��+���n�^:ū�w{��{�ax;��ܣVSGj�]c4�.�Ӄf���4?���=�]�����vD��$�h�xJ��P���Ͱ���Ά�^;�y���r79���dq�F<�K�
�.oQǰ��rA�Nllc���k�m�Y�/���4 �g5֌�p�V���y@��q��'j]3w������{�3z��}���9��X��s�2v���ˉ����9�ob}���Y��B�gN�eVnv�U�n�&nͶ��.��ia��M'f�E=�g��盈�'���*T�Fµt��Ax$��I����75ޑ�Aek��bO;ý��[/oHV-y���"�T��Gn������p�wev��e��;AnT�n�\�^s1�0�+�F���j�'L�!)�WrN���a|�`=Ʀ��(���YP��Q1��k�L�Ѯ�{�t��͢�*�@���\��ZH�u��	ѡ$�)I�]�1�9,[����� �ӎM�����4��9l�J�l�N���V#y��ggI3]�+��[{��GSUՋ���l��9r�4�sF����뒂�v��}Z�,��f�7wvv�X]�do��@�{�^�{< -�o��ٶ��N����;��lcYV��[9�6n��f͘Ʉ��s�j�F� ��t���M<����q�H��F1�;(�n�z�8���^C��������o����Ƒ/��ҳUZu�ۉ+����@*��z14ב;�,"'V3C��r.�h��+��m�SM�4�4l��z��х�q�P/�odo�'�HI�"f�g		Bz�����ä\S���uo��, �o"��wk��N��4��b�2���jۜ`tNSz�ם�~#+�ჰR�͏�oM��Vv�%ɛ�H-�{������4h��߈��E�״9��fk��n�c
k��I��?��6���x���G������� 'ion��^(�j܏�|ZR�4�tr�����7�`ɴnn������h�Л�y�!����j�Xq����H� �[�'&�a���Kɻ�B~8�|7T{���㛯��I&��<t�3F���n9ǳ��8ʛP��+�fl�:�]�7�h���&XR黤����鑑m��#U�#PpKf#��H寣����4Qup��*�w��{;�m�Drj���5��w8��S5�ܷ�ghى���㵭�
�NT	.�ၱ��Ͷn!�qѧ����%���"/]4�ťR�;Y89��U�w1�NO�8hxӋl�t��`n�p޼_<�qԋ�ɳc&�;�oM38��'3��q�6�a�q��K� ��''���<4A��ۚ��:v�a�M���ݙ���`��f[�EjI��q{+(�-�3A(���F��I�+�z�Lߞ�|��C�G�zG�NLv!4f�E�͢��4��ίq��ގ*�|����Ŝ����@p�,H�
adx�Ćtۄ��x�@��S���ݚ�~!�r�x%�������2Sq]([��#��n�X�\��̝1v�ll9�a�;�t�ú�ܴ�2ό����f�3�@mowN�Qnˢ�����3w�޳��װd�{���`�qJ'�:���غ)�\z�<���v��,������Q.����KH�.-*81������ɢ�9���7G�(�9Iֺ=�dA̓x,�츺Q-����
��ř>᪭�g[��`/Go��XV��h��wK�@��3~�z����x�xQ��&�88n�f���M�)��
�����\x�Q@s� �Z|�'�Odq[R/�{��n�����[��Aփ�[�>�׆�eb�-Û�wm�zh�*�����Zy����������N�հ��"x+�+Dr�ȵv=�.U{H�u�r����.j�V�_9�7�Q�_�؎^�BiT����+;m�y�Qnez���2W�9i]��k�.o�l���X۠>�N�ݿ"�A)=�s�1�i/#xn�dp���v���*�v.y4��Á�i���<;���'_FW7ǥ�q2;_�*K�����]�˿mD�NYt捋&�F���OQ�v��x&���Ç��D�.�y�]X�m�e�<Y.6���]Kk��#��9f��鲝�21۽�l�>��vC�[0f����ɝ���\i�U7���A>�ٺ��Y� A����0n氞�H�xŧR��k�A@��
��d٭휯0�2�����!��"����̱�ܧ�^}�Xx�v�h���*z���1�;2���q���3-� ��j�-q�GAo���<�"�
����zչ��1���#�ʛ7'gm-��N��\�.�,�{t����CT<���l3��}��"K{k6o8�sa԰j8q�ܵ��U�f,C-�HCR�}�(u���YL꒍7V�?< ����t�r���;���&�%���c�"�5�u��tj:��@��.0��k�����u�{	�]�'d�b-���
a�v�����<8���=�oi��OlC�J6��U �f���5@ �HG�0g��盯#z�@����wV��v��b�9ǵf8Ci���w@;p�k~�j��z�(-�9j��2n��gN��y��rB{����Pe�i�|��c;9W6tG���Bpt�ƗuL�*>@)vn>	v �/��E��û/M�
vn(8��f��w7-å����wl:j��"�3�v�+op��7�� �+�@;t�S���hvDN���@��|�5�@v�V��,rH����r�/]�[�^�&+���$FWDҔ��4��{��}���o��pu�Agd��:�&�Z���|z�YCZ}����iЫ���sǛ�h;3�����7R$2�o���ە;�ѤI�@�n6(}�s��K�����CGer�Cbr�;&G�E�
˂ '� Е�2M�Ap7��-/�|z�zP�hthJ�j�$6���F�V�.�S�<8ņtq�{�e{���G�w����]0`nn���ew��F����4�5�=����ݰ�m؎+�NR�`=1�G*t�eY�����:k�����"����ٞ��ض)�sh�;+8`ّ�_��]ٳ����� ���=�Wn��O�z�6������M:-�f�9�&�����p*Q�=����{q���aO��N>u0��J&�oB�X�3�ѵ�����2�gd]�c��xGχ:m2�4�E�����t�1�]��u��,��4�!���5ur����D]��[��x�K3q�oS�++�n�~t�u�r���Zwr<O�P�R���gh)\uڈ�b ��h��&��j���;�P��� �W/s��y�vz�"dX��pͧc"z�^o���Q���~�j�2m1exۻ���OT��c&4Ww�1�^9�H��N{��������7KЏc��;�n�R���N���8C�t�]����C����uvj��ʇN��H��Jj32q#t�w&��Tݓ���N���uS����Gv껅#�]���n�����Q�N��Xv�0�%�ñN�\b��j��ʷ���Б�ax�D˱3�3��ۄ��w���S��x؝h��v�7&���!�.E�N��Q�nV�;v��iWS�*�',#wx>e�G�O��g3�sF�cn�gWؤ{���o8\�N����Om+y�]tn��vSږIf���s��-���Z��V���:�-��˸ VsQ�c��7F�����OT����8�㣉���Q��C��l�Otz�sL���]:e�gA��qm�z��6n<3�������r��NP���r�w>��rM���o��ӓ7K߷�v�îQ~�.�.��	ӄh�;9�ix��h2��f��ҔGV��:�	�s	�
�6�.k<%$��͌��ټ冢�s���=��m����v����w����h���w�9[���eC��:��Y&�׷s��Y��7���hx�JuX��S��A� ����"q�b�5���'-f杚N)qP����]E�T�7]ook칿F�vE%�PS�4�� ^�K��h�[ę/Cʭ���s;tb�v�k����b�jhv���k�a[�9�|��������AwL��^����0KGfك�]Ji�jFi<S���K�f>sf��T��͟f�ΐگH^۹�#�ymC;�io��c�qk���&+��<�����ໟ)�	i/���1���׈-ì˝��Ǘ��6�N !qd"�gt5�:kES�I�B��#�]��U��f%�]�eczp[ZQz�wp��a'�:e+=�]��444���W��R�eJ>�0�H���`�^H�8�ݶ�l:���<$<"$���j�w]NO��2��k� ���\�C�e�����m[�`�3�V�:�Y{Vw�X�a6���{az��4��.����K���}&7K]cܺ�s��ߺ��'�o� ���BHE�Y!�� `H����P��E��RB
BH�H@�Z��$�Y$�
`B)  ��"�@$�I	*@�d�E d
BH� (@�P!P	,�
�H	$��$�VBHH( AHI$��`�I!P )	!P$RA`IX�$��XI%B,� �B�J���$+ �*Hd�"�d$���T�T$�	$R �$PV ,�, 
$Y)!P�`�BBVE$��!$X@@	Y  �HaVP �$��)RB�d���$��+
��B		���$�����>�����y��� ��5��^3��{#��V��v�g�����{�e�E�}�I��{a��j@��r�`�1x����yl�#6�6�W�����<����go�x�+���{j�P����)H�[H��Qɒ�c"%�F%�QrBnZ�wY��'�k`�Z�m}�e!�٧:����n�Ӛ(˛JA�0aI0}��h(��w���;#�˴
��`��t���|�޸O���fwH��4�������=.���v0�_�nԡ'��1)7����s�<���{FkWF��~���v��g{�{�7�P�<��K5�Բ��D��OY��A���Ƚ�S�t����oa�6�xi�.K}�{gx̳�d��|���<����M��{V�{��:��"�n諑n����^�}�{ʫ��Cg_!�A����^7�wތ(��be�(���MRwg�"G�<�[�b�M(S�/�n�(���EW�����!�Eo���->#�%���}�׮u����n���N3.���u���hW�k��lZ��|x�'w4}�D��C7� ���������'7����'��}ӛ���I����5P�����?'����C�]��L��xyه}��z�w� ��[祀6-W8$��s��b�;�Eq�`yױnV7���;Fž��Ւp�iq�o]����[�_v��i�[��V�)�L6�ʌY�Em'N���Q����p�J�u�ؽ��\l�b�"^���s��H�_�8�oM��ɤ�މQ��戽"��A���=���Ӟݹ|AG�+4��܉���ҷ�t�Y=js�FR��S�4b��WNs8�os��צ#�u��˻�Bz|
�Y�r�Vy]��K���jmW�v�;�_D���� �^|x<��'�S����!�B\yc���F����Cg!ٯ,��r�X�W��q��+TIO}B!�R��a��-�����hA��x�z�ž�<���ۙJ'ѣ��n-�T�\C7�K7voa���֖�ÌFݜ����:���X� ܞ�%�����K�[�ٓ��閐bxG��F��H6�S�܋�N����x��}۔H<�r7ޢ�Tje1b	̤6�N'���ȱ���W��v��N��͋�F�8�;��$��s�Û��:-����؊0UXK;5ghѮhއV�ܩx�1s`���lŽ���������{�MJ���`P����NI{��'f����cQ�3���*���^�7s�k�<7|mSx}�b��Dּ��u��St�j�ֆ�-X/�dp��������n��^T�ۋ�g\�������&��z�c;�&d���܁��zu����Ė�o���םɓ��ܷ=�����h�drC�ȲC�E9y�A��7(�p>׾�uC��ݍ]���K���>~�"��ow�ѯ=�����1ټtkkg���y=d��|w!����'jy.yV�gp��F�A���%�螔����O��.�O��픗�@=u�jKB[�ο1�ر����&u���S�6Y����7����`�ۨgzy��c�9zuL#�=
�&��o9�����﷎;�ha�*�w���y�s�Ӡ��힅 )��&c����ޙ�/.��J�uMg��sk��@j^΋���-Z��1�z]�υH�o��ٛ������GU�j���e�&��c(n�]Y�������V����=���[�z���S��90q�y���/�pC�h8z������/�y0�U�(E���G�8j�Ԩ�g�8��!�$�^?��:�����R���>�y��������yԦvL�����_]�өm:�n]랖b�r�����[Rwv���(j�6��Xt�0��Q�#�a���k��B�S&,�̀��.`J��
���x�٭`��:�7O�z�{��E���Q�L-����	�n�n�¦r�Q4�D趕=�ӻ�3S��ٔ�-����l�/o_i��g7�e7�G�)�;q;6���r��lL-�ba+,j,Ő�SU���XF��-
���֝	�|RV�������m׼yz�ٰq}����II=b��<����q2�>�3}�H��zx��onˊh�k����v0�-�2e+�Efi0챑Y�=rk��1{�z�߯[nk�vN�Ȼ̼���V���U�0����	P77��/b
]B/ 2��]j��Gt�'/��e8��t]cٺ���.4����G@>����m]�Î,^�������<i�;�$p��;����|������U�|p�|1�D�	��He�b���͋��J�/9�c}y���-���٢o�ù�
 ����Ab-w�p���������E(�1���q�<\=[�w��5���u-�*|7�����~�����<Cyۋ��p^Ҟ�x7�=[~EY}o� M�ǂf!�;�′%ɒwR���u{tj��5���詤�T�̠��8�io�������1��e�5loؖ�ͱ����TG��:v���؟���ۛ�5p�l��v���3����1�w7�	N�p�G�zC����r=���g��s��e� f�7�R�=�r��rИw����S��8���ySD���=�s^�}���Nz����{a
�Ȕ����8�{216�l�{�z}6]w�n����������go�w���򨱎�O-]'�_����O��鳧+��~	+�5	�L�C�&�ST]����� �߼�;�ˁ���
�)��K���Y���X��s�0�}t�5-���E�M�U�%�v���NziH��<]ZS���'���;�\���{�����;�+�16��l���d`�=5{g��G�x"SdY������Ӫ�ޣ��ַ=��dm�Ke��b�N��2�Z���j7]�Z}���\�=��Q�k��Ak�FX�G�%�vJ׽NqWd=�9?z0����+h)��E]>���V�ٲ��E�^������;��^��B��ʅq��]h@&#}62-���f�L��;�c�k�:�bc�T����lomj����;T8�b6	o�����{:��<�:��)ޗi�	Et�j�<�+��nz���R�蘑�cjQt&+'r�|U�S��yJ���eR��Ty���Z(���	3� ݾ�Sg���!V�BX��X�⋬��"d�l��9.��TF�~w�Zk�Й���n��y=�:b�N�!$[��y�Vw�f�/,ﲙ���w�u6��n�{z�tW��ya�{��tca�����������3������ӽ5|�<�t���l'�u��$ׇ��x�V�FRLh�wC�q�����Q�����=u'�����zaڲ̷3q�%�zn!�D5��zȆ��� �\1��l��;��Rß O
��?m+��Vr�[^JI;��1b�,���f�7L7csLd��6d|x���9�_��an��*�}��{�vй��n� �bÐ���(=�/,��;�]��To���gg����n/o�銭���b�T�{�����׎W���ہ���R�R.��z}:j����Ӟ:�?[�� \�_Ox�}�)�b�E�JY����IA��|�y�jC	}��ȳ�o<���oE�-�/s����aLdam���?�;�"��ؼ�9�v6�B3N�.���m'�`�����:ӷ���m���o����{��}�7xuO���ٓ*R��x-�7��,/�[!��6���[@0=��|��r����v��E����<�t>��l�"L�L��>�Fjz ��zz����ڱG�NU��D��r G��r�>�k��F�vZ�@P�]�]�c��^z՛��Fi{�u���e7E����x��?i��>���noz1�J�$���%���9���N�r�f����z�����w��A��#"��f(�lM䶔��k�����z���]�t�&�0��	���;�z/��{4]~*z����-Mz����-3G�Ѫ���œ��3�%`�A���[����z�v�ow^�Oj�}�<囇�
a�G�$�Ț4�kѷ��yL��a�F�{�>�c;�DX�=��,�;~ �<t[w{{�{8�NB�=֡b�ӳ�E~�@��a���xxe��'�k�)�ؘ~=K���I��Ǽ�[��]ٻs�Q���~U�kl[н���ʞ.�}ϱ�^�@����O{x��?]:_zo%�:ũ͊�����F=��ϩ���I�Ќ���P��6��f����:2��7fz��o��b�GMSO����{�:��I�ʚ75�Nn*qha�^�wE�/.7ܻ_�\\	�����	G��{��#w`/����j�a��z���{�q���ű���˞���Dp��r��[=}�B"{���3p�zq�ؘ�<z�3V#��ކq�/�'mw���4��Kk�{p�wNq~ǳPh��(od�i rQ�.3݃}���;�xjӦ���R�&xq����&rV�fmL[v7f�_�nLP�DJ�y�oV�@�n\mH� ��s��ď�s,(ɿ
w��_{w�:W��]���U�iͽ�vyh�|=�d�:����}��T�Ӵ�TdTI��[����5�����������1�	b��w1^?k��V�{_�z7���~�B�@[<c5A��#����>~�w�A��+�M�������l�����c���:M��}�״r��|���s��*���È�ۂȏd����|�82�}��U*�fz��yݑ+gt� ���&�R�r��w�ۙ㩮3�Æ���|<�
��0p[�Ԯ� ����9ݳ�N �2v��>�o� �O���'˂��	����9�7��:ך:f��=g��y��W���;�v�|�kA�M3]>WB�|��)R �/�0wc�r�(�BN�^�q��Cn���u{}4<��rd��b��za��]�T/�"od���x���u���w>j�-ܐ�
�F�͙���R6!�S;9g���I�c�\��:{��;����l����٦n<�m�A�g{��S�W�pwW}�P:�ư�w��T�G�o���g�w�
~�^��X��SD]^^�N���KR#�{�מ���->����i,!�n�\�:By�u�$=�[7�RF�;.�x5�!U|py.��{T9c��<z�9�팿f�	�=4tZ}�ޮ�.�e��B��|�vn$"�()�ks��b��h��4�֏MѾ��������V��3ϴ���`Kh��*��2ֽ��x!V�����pt�!܏��/6�=;|&r��x/1Q��l{p�lB�\`Y�ɥ�o�L�=i&zsX\o�tZ��W��&t�<���q�Ή��knT����f�n����O�=�Ż��j�b��cޙ�ؽ��o��|,�n��V3���͝t��T�AJnD�ծu؝�*����8���q�h��2Հc�E�O��28��z�;����������2'�^VE�s�9�9��EÏ����^�y�I���8�1��i�/x��=�����<����lCx`>�v<���x�HE/���8���3{����"��ѻ<��w9��8+"���m���fju/E��܎A�����bI���}i �� c>��J������g�7�t�dn����e�g���ك���:
|
"�W�w_d�O�������E�'[�;Q����uYy�Kb��r��[��u����Պg ������Y0$^DnM�1-�{B
��vT�F�|��7�z��~η�C ���8G�	��*}��Fm�#�H����s}�1x�(��甗���l�m�h�XÛ���-�$C:Cё�Uєv���4p������v<�X!p��T�K���\A����k��?%�1���ݣ@f�'�V���F�N�׳W(G��K�������.k˔����	�y�4���v��~w�W>�z*;�[V�Ay��7�zi[�Ft�;��[ef�ߪ��j����zL)�j��TL�.��vJHX$ {=���x��A�֎��K*<�^:ޚ�e˗��v���P�}o_�x�����~[=3M�b�70ӭ^�x[��N��c��)3�H�+�W�_9�*�Y�]x�K�;5���  ���|�f�`�o��μ_�!�Y}�U�����9����{�Nv7Ɛ<g�y�;7��I<{z8^�=o�n���{<��{7	�m���痮�8�Ew���{�������z/v�۝y/oiO��wg�)�*e�,�E谆@�{}��UVl�s����r/ ;y�!��{�8/zU
��>(O{�7�zA.��jg��\<���1K����!���'H��۴�E�}�T��O��q�{�7��(�l��D��=�޻y�_wO�P����ƭ�վ����j�y���{A�u�rS������B#�j��:�[�)Cm^�z�����c(��}ޞ��^Ӡe.o1}���ċ��oc0|`@ao�{�u�C$��hs�y�&�gyS�ܩ��K&{�!y�Zwa���|�������w��4����{}�㽡���>f�,�m�j��2�8�置x�����瘽Jl��J� �<:�|��yD�Υ�b��6-K���/f����B�t��K��ؼ�8o��=�J]&�<�LQ�␨t�޸�P�&�[n��Bz�g�*/`>#��<'������͒;����=�Q��|��Jk~<W{�Լ�_�<j�
�`��&�g� �Ib(��^���{z4�c��n�=~h���m㇮�!
q�ŚS��L��n���jq�!�R[Wy�����b�Bfh;�\E��fFwg'��zE���cyh�.p��w�{�w6s,o�}����Q.�N_=���J%�[��I��0	�~�nSN��'��,V\����xx{�;���m���퉫/"�vu�WS�=.ٸ���[Q��]%�As���sl�yxzWY�	.f�n���CYv�ղ��r��6�h��*=�QH;\I�֚�^�<�HF�{s�s�S��tK[[�l�t��1Ϊ��Ȟ�Z�{Y�(<�	j��M��su[`(B)4]�n;��XWk+�aK��0��r�%�Һ�j�cp�C�Î����4�ʜ'k|m�����K���{[\VG\\rv���X������p:7BN���p����Ipb�l�#s���z��H�=�u�z#Ѵkcu���{^y�r������c�Jx�O*{j��jG)���ر�g���1�ݝ�Lp��`�C&���.��s�';���kF�6�tv7Oj�zݽ�\v�n�qۃ1��P�[�c]N�����i:1<��ى��c-�9��V�:�2�N�G��cW]n�s�cE���c��ۍ��Jq�W��,Eaӹy+g=��r�������3M1�ڣn0A����4��sAa��v���7���*�ږ�=��z7t۳B�۵Wn\�a1�ʽ��:�g]��+ �W��Jr��]��\��z�]�Ӹ-��K�	�"]K]=f⇸Q�Ǟ�;fn]�AۇG����V�B�������v-ͫk���\u�W@ې6���lW-�p���^o8��7�`��{b��{cX�ۜ��Aێ��������T�V�����;�vԥ{7<U��r�Ms��n��q�hd{��%,5���˶�x�z�:��`Gp��ڑ��5�=H��D��s�����M�v�T�Z���=`T�kK�n���&l^�p�e�=n����Zm�{=���cu۳͆<�����ݬOn֤�8���.ݭ���ó۞l� ���u�b�f�%�3:�۶ݏQn�]�S�ݎ���nmC�v�(ᤳx��Ū�]��-V0<����m[mo>2�v�Ațr\F��{���Me\lM�R�Nۂ�sN�)�B�^E��6�:V�Ƹ���NE�6b�-%�F�^9v&��^�6�ې�Q��Y8���EED;��y��j�s�s��;fW�jX��3�nw�h�ۃw0OӴI�è���f!���k�^q��R�6��^1�m�����b�{mRS��69v����ۢ+rc���x��{v���ҁ�1q��n֜v�m�G]�Ã���Ჺ^-����O=\^�76ٷsX8�l�jv�h�z��۶4h�#av�ۥ읙n+��[�W,�����ix�̗g�;�':�6�t�p�8�m��e��]��]q��5&N�!=�����o+���'clg�O"<m��,��;oA��{u��n�q�j�,�mq��+�/N!waa�=,��v���{=#�wA�O�XC��ܐ�|��}�nu�{D�շf����9.�[u>x��<vsʇq�=��l��]���sE����3�Ҏ�%�ΞN�7�OZ��Ip�#\��Zطi�g8��pN�D�8$��Om�vv�ktq�6mۊ�8n$N"=��Fn���:�[X6�j���:�Vt��u�6���'&�ݺ�-�Cx�g���/Y%���-�+��c<��{g¸��8qA�qgS�}W��!��b�W�q�V��ʽsJ�;��]�W��ccly��:p�c�g�N�뷠ݝ�B �n���c��֤��=`E�ػ<�t��m�j���:��»�&ԲY{>G���=���rz�7�2M<Z�soOn��LS�6҈�7Y�$觳ջn��ERge��Η��!	�\�tvS�Ͷ��mn��w�P.8�r��Wq�����N-�@ی]���� �q��M��nN��u��c�PrkGZk�S����mT�&���ּ�FלrY�v��=Wl�'[F�}��锵ѷsm��vڲƜ]#;���XP6�>9.9�.�����:�����mҁ�n���{mN����ox�k��8+f�D;ILN�����y�3�eݹu���\����p��U�A��`�s��5m��ۂݺ��s��6Mlwq��N'�3�g]�s���99Q퓧�˻V��Q�;G������I���>ۦ7m[֎-����ݴ��:I�cg��pnCsi��^W��wn��v읗#����W8�t3�l��X���i|��kLr���v�hs�.�G=&���X+���̙Uٴ�!�t��v94z�ntI8{:lX��j냧J��]�-�����t!&-�br'lu�-ŝ�mm�u�Uni��YM[u�2�]��
+#
�"k��؝�#��-�E�u��ђ<�[]�2YG���N�i�[�x��qpuvؼ	���8;n4q�V���r��^�u�3ཹ�k��OgD�A�f݅��JӋ+��HK�N��;u�l��;@sv�.^=c�����z�s�H�qҖ�t�'��Sv-�9�{c�pCmq���q�ոjm��8�=��u��66�Dp����[���IϞ���<�^s���q�)�s5��bIѝ��y���f��#m��7��:�kr�\In��[�M�.-Z���m��z�i칢���c�yU�G�N��]����l��mv��[e3wm�����`�V�1�n�> �^;W�pg��z���tܻ�Cf��.��`�jY�ի��K�6�գ.rG�����˻vu�O��A�6;*����lE/]��{rr�X�gg5͗�l�n�o��O���';܋�ظ �:�7�6u���j8�9y��&��T�x��e�����Vl�n<��0��]�n7=`�Y��9`�5`uݷo�N��JDv��y�Gp��9츫�W;i�ɱ�f��a�q�p�vk�H8Mi�B���\q�u�Q]-��k��m�{S�<���۵�`���#j�`��]��QG��췶��1��ۤ�r��,��'�1�^�q�.j0��F�]�h��}Y8�I�w���8�^ϐ��[�fwq�����rs9�7.�o7.D�^D�5N��.�7�6¯v5��v��Ѹ�a�&�����옄�c:nm<=�є��uuӸ�r��=cg`9Ųsv��@.ַn��n�טb�N����X9�ո� �m�z�r'nۭ������]���cƲ=��� f��nC�-��D<ܥ�Ϟ��^w�7�͞q�3��g��up�]�����s�s�k��^�6<��������;&�b�<o�	t�#�ٍ�=+r�N�^���u��=�+��fy§�.�v��V���狈1���%#��n�;��u��%4ⷣ����ݘv���i�
nƂ�^n�l��1�m�0%�X�n����Gn�8p^����N��pۣB��q��˵�.�l���j�X%�Վg�����Y ��cK�����xp���t7m���ݺ�r8�vy�5O�����w#�jq�Cr�	�����V$�\nv���:����^�=$�)��91�����x�J\7f{e�3������z�oEy�� [vk!c��r5=D��T<�>8����7�-�[�q�Λ��]m�.�=\Y��\�2ջy�o`K\��u����np��֍�S��nɣ� �n�p�n�:R��mpm�h682Ps.�ŭ�{p�۷*���I��ۮ;'��o�;;�vv���1��뎺16\���v�!rB��j�'c[�Iѝn�"�t��0��e�K���47���jT۲k�8y#��ƷoC��9��ۉベ뷞}mod܁x��$��e�k�r��ֻ۶\%�!�v������.4�u�V�����mo;�Dű�ݍ;\ζj�t�g�fX���s/�v�sb�y]��pn�h�kV�3�m�ݔ�����є�x�����iΨk�ܶ|+\��	�!����۝����g{d}��#�����<��c/sˠ�՘���\-�q��:=#�Հp���s��]��g
��;�ܱv���7S���qS����ur���;������e�q��w9���v�pY����vS��4���xl	ͷ�L:2-�NJ.ɂ�����5���Z%��z=��I"����V݀�������;����ŷ9kk�o;�Gu�:�Whȷ]�=sOke��GG
�O;���FN������-[�o��.���S�-���[����=$�]ی:E�.\�lÐ��=����6�ӹ���Ac�'�{&{^w�F�5�m�	�m��n�9�gln���x�l]���<�y�&�\Z�n�vy��v��@M��8��6.5��caN�u��[fx==�q�Μ�ZD�t�:!\�iܽjk�Ѹy�.���#X[����5�����{�'K�ggr��\�.s>����y�.=uۆ��%��[t�:�r�j9S�x3��Z9K9n�8q�s���t��]5�ڶ:�\c�k���糋��ذtWɆ���;l\���:ͬ�����x�����a�y���۶D��g��j�с�7a�$7c���C��%��N1��q�q�����C7	۶��-Z^9��ڦ��]p�m[]��з;h�ewu�&�����qmo�X1��0�s��G.�0pݭ�z;�۱��T9.8�oV��q��L��Wp��L�l]��<6/�X���t�ҝ��:^V�-�6�:킉y#c�G.&Pަ��z�]�V�[�[6�τ⻭pgv�3��:͜=j�a�=Yk�[��7i���[K��Evy��$Gm�,��\���۷.��5�*Rnt-�w�x�]����\ ���;QN{g.��X9�,�Π�Y,GiǦ'z�F���td6�3�n��U�m>4�'<��r�����ՌOn��n�EwJ]�\N �m���k�r����;f���qg�g<�bBi���.���Y��ٶ�귇=t��Im�5l�����UH�V���Ej��J��J��R�f++1̱2˘�Ũ���m�LJ8�1�EƉXR�E�J���ժ��E��JYUe�YXTib�UT��Z��*TkFZ�mE-�Ҫ���Ŷ�-[����iQj�j�K*T���h�r��[l��DKj��q���Աkm����AD*TV��mh��"�Q�l��FV�U��Z��clZ�,ZԴ�QTKT����T�Y[+Pm-�
�m�FT��E�R�X�Q[mF؍jZ4�PYVթUPQ���j��Z5DUKB��֌�EKil*[-jT�����h�����̖(�Q��lYl���(і�ҵ�Q+AI+"�d�Jԭl[J�)Vf\DJ�El�D��b���kh�1�1j�,�m�E@Ql���R��H��`T�KH�
[X+Y�e��,�Z�JJеU���ŵ�bT�I3nq4kO��[w�
6�f�֢f����E�K�sX��ޓή8��g�[�����x���]��mf�䍹�7\q��6[�]ץ݃�t����67"�۱]�x�k9��0n�ۇ����s����'��/|�e�ݼg�ݶ��̝��:RN�eŝm*`9K����`K���aCX8���wl����9��aug��㥆96�.�6�C<!<�[=���;L�5��h�|uٯ6�m
n{���p<�B��j�!�:U�l�]�CĘ;h#vv,sfwj��x1vK�띣���ĕ��7Ck��kmػMv�ml�6�*�a�{t`�u�w`��t��E������*��'z��ǀ�ǭ�q�.����U�l[�����<ƀ�z{v9�i��z������]��gHl��.ǔ��n�Zh���s����m���s�x�<�]������orr������%�u\�EOc�{��;�oZx�i���0Yc�]�M��[��l� L�gqY�6��^�Ib��H�c�҅ W�q�m�ݺF�Ui"��ݽ]$;�N�Ɣ@㸸ε�,/���Ί���=�]C���v9ܲ)[=p���oJ
����y�=�����c�w��ظk���x���D2�۠�v���n�7u��n�G5��;n�n5��e���l{rv�t�5���ID���;	����7fżh������;s�\��q;ٸ�i�C;//Z��ͯ8U8�v9������l�@뉶��v�:��=���M�}'AV|��]���2�`�sTX�6�D��`l<��2k��.���l���َ5�ۗ��������M��Y��08{c�#��q��q��=���C������~r����N<����m���Ǜk�Pn�T+Wv��x\*��m*�v��5.O]ls��WY�M���&<����@.�cO�������F܀����=�yW���N���L��q����y�����;;��v2�c�;dx�n1�&����ɲ=�r����8�<�{g����g6�_.w�l���1˱�۶��w<N��p����)����u�ݼ�'�l���v�<��vTx�Q�cn{�Se���pl�w>97˶�2��c���;og�|�s��B($�a%���K)�؄C�V]̂V^���$�ݦ$�^}�.Y�sUuD o{��q#�
]���� ��әQS�@�B��@�c����b�
�nc�kĊx
ȇ�S����	3��$��=�F8���I+�z��;��XCF
E7@H�7=|t�E���껸�Q �ꪚ$���tD���N�O��j��� ����@-�
X
���'Ȃ�ڥvMVM���&z{(P$܊�%��$�6��������M�g��WV��p���'��m0��.���k���6�ۓ��q��~���Ҝ�Dw�n���I�ȩDo���P�K�x��+�� ��Rt�3d�� �h�Bn����H��qV�Y�3,Or1s�l]�6`K�,������r�,��w�X߷��O�_�������j{����Iɨ��vr����H&7]$|��W�R�ݍ�**:���bǠ(,��b$�!K}�^�|X=yn�|�^���N|||�wUB7!Y�sA��Q���v4E�� ��9�> ��nU[�ջ`O3�n�rto�v��a�4`�8i������
$��{�A��\o0�f�EF\��>$7��D�;����0OI�'X��n#�Q�!�C\��!�;[��ٚ��Aۂ㷶p�����C&3o	�Aa��z6n�	-�mQ$���v��LY�j 7W��	��W�l��D@�Lz����u���ѫ9�>!�������@�e���;��㍺�3d��l4C����@1ٽ5�I3��^�[(H��N\�Y
�f�I62�pMiۺ�[�|���J��`_�=��H�"/"�Y$��{��=���{S�/ԧ���RH�C/L��8Ufm��{>]}Ӡ�"�ǡL��b$Ս��<�/�q�y8�ܙ$���@�����5�MА_o9$`y�%d'�0��nz��gS������^ ��3$��ސt�5]�qU=[��D��D��	¹ص����X=r5WT��P݋�.���W��i��e��p`�8n
G�^�̒G�_n�A+��O�S�jbhM*��<H1ٻ4b�I�Aa��s@�v9�$�=u��J����$���� ���r'.*"���+��L���1��Q""2c���9���'����
�_:�޶qAu��Ȯͪ �I]���83d��,8!���N��m��E�ޑ@�H]["I�[��{���ٺ�UG�T�{DC�Q�[2:f�B;�uZU��Nlly�"���+*б=c�����j��6{zd��#ȢXI�/tt ��\z���i��Vf�P$VֹWoL�y�mY�� ��A�p���ՙ��S��`)9".MX@0�n�us���a뗣�~���\ڄ�w�l�
!ek�I>$�� E�W�d�1N=w���+k��u`�.
%3C����s'�ƘmQ�Ӿ�H+k��	�[��M�N���I�d���|)��"��x�8܂�� �UgL���1ۥYp��!uc�A!n�ρ�c���DDdǧՕ�Jӈ��&x�r'\���|��gĂDWwV��2�('f�ImېN�8j�-�XpC��D�O�WgMs�tiE��b��I ���<DwF�g���50�乼^nF,��%
M�n9��ۑ��ɫc*��D�<��B0�?��f#��5���E�0��b��U%��P�١qo㛓���y��::V�z�:L�R���l���gY��q�&ۗ���w&ּ��lR�A��د�5\�;n��c����Ӟ�K6gAڎͰ�F��^�˼�Cv�ŷb{d�ns�.�@Hb	���j������mM��A�g��mp�����-�§��Y�v�W]��'F�c=Dն0��^�gQ�qm��Fh$����J}����g[V\[]q�������K��QkD%�v�� ~��$�EouQAɃsٸ)��15O\��	�ݑ X}�+���[P���z�ē�:�w�{5N�$�#3fA ��$-nL=5�	Y�7�iK��L���H�/z�H$���|EsJ�yS��1cl.�`��c7��I��T1]��L6�n���7~$����H&;�j���x"=EP=.��ٙ�24�dDC������@��)�G��[�)�L��o4��rDf�MI]��,�[aTD]���ु�0àV7c�tVx��=a��v�wGD5h���`3r&U�<���h0�x�V1 �^t�$WuH��)��2�G7� �s��+rIr�K	"��J�����\�ͷ�Rm��a4��n=�^r��+���svH��q�f�bEbl�oz�BȰ�Fi��T���W��%m̗�uo�/�e�O�7=�T>+�\�A1��|UgE+�Nw��z҄Kd��'46]�
$��s�|H=��|o2�j�פ�EOv�	+�X��tba \"�j
^��G_S��Q �͚��@]�"I ���s�d�x�o�I>��#X�x�܆��ω�Y�<C�W��͂E�v�H+r\�I{�2n��g;2z�F�	�=�\�7.�������u���W�ٽ�^ܫ�v9�I;���1&��_~~��0 0��s�I���z�65���g�OUP�H+v\�i8���h0�.��W9,H�i��sOF����|H�y"|>}}2H=j�r{��d��a�N"#�BA�$b$5�|O�%��Bԑ�X��-VK�L�`}WL�kf��/0QQ�J	���H����{ܵ������hn�k¡�l9K1��dN^�ȭކr;j���E��^�]Vh�l;�$�o����rh=�Z�H�KjsC�o�F��k�㵝&s�ψ �ݲ'Ď�ޤ!���v�4I��rv�ه	�H�`� ��bA��٣1�j��3n�"fzD�g1$��w����������q�"#��tv��;<5���X�[��l���=��8�i�O�d?���3��l��eݿ�$Y�$��~�ު�;<]L�I�����=~�@u�2	�#�������l�������MpyDc�̷@�K�� ��ޚ'Ƶ����dGv�˯ZN*�CM�?7Tn�fI��5�1��у&f����I��wLc�(���H�H.k�˫��E�Wl�A����Y;�D�V����ĭ�v�hwO>]y�r������^�w�%�n+���U]���$��y4I0:}ȵ|�ո9\�� $�ˣU390`��k$M��E���`������\��;8#�(P��z0���];�^$������sG���|�{:����g�q�������Ö�u�u6�u\[�Z{Us�Ɠ����?P��8���'��{;�@�H�}"AM�Ѻ�&aTs�	$]��Q3=��n<����Q��rD�l�a)��S.��H���(���|p����[��b�����	�������P���uݕ@�
��H$��nEl��΍	�>ͪ �����p�m�a������f ���%V�Mx�A+_H�^�9r�wJ�4���=Y=B�
�i��
!�{�@$��D��*to:3�6j� �o��I������qc�)��e������2j}�Wj�5�=wqn��N�4����<�Ӟ��,�_�1�8�Ů�R����չ=�]��5�ɋ��L�Wu���`
��k-ׅ6�sj����<�g�c��qb�ӻv�n��[m�����w�ڵt��9���pr^1���kJ���L]�q�y��u����{7'W�Z�=�^v�V�U�M�7;t���Cw�y:�0��c�m3u�k�J;�Y匰K׃�<ɷ2���u��.�z���緈���v�s?��+����ջ ��Q�;l�[m�t�c�N��(x�1睵�`�GRW���5���٤r�H�%���}��*�>\�ω ���A����Gyu��TA�\��=��Ä�p
�(H/��I�:�����U9�I ��dI�����������aU �}���&�q��l�ꁾ�rH$Y� �ƌ�A�}�+/,X$���ľΙ'؏;��E���~�]�M��"S�q�Ƚ�s�|H.��u���s֧�m��BrGw���t��4��y����I�:h�$��"i>W�,n<�$���zD�}�5�;Rv'(ܹ��{�/�2K,�I j�v��պ`�;9�����ݮ:�c����>���.zTG��|�ْ	� k��WWn�����@$;Ι$Pv8ڈH�%���W7}T	1�aP�f�Y֒���A����mG)��������Ğ24u�A�xU�,����ŗ��^�&,�U|)�"Z/V�k�&r!l�3S6����gN	J�D��|	$��rO��z�������U9�V�{�]��H80l����r$�A�ݳ@��w��K�_��c�	���K��m7PX�n���w�:[��we�$��O����$�V�q��
�	&���:O;��	�M�.�r��IY<��芰���38�$Kڑ �s�ڠO�[<ė�*2���@�QP��:�^z�kF
��]����d��S������8{YB�0��w�T�$�u�t��B��k%gH�g����	'�vС��c%�0B
"|b{�	�e���^�v+:zF�e�u
$��rAihV���6��xڈH���b�ӄ�|
� �k�Cx�DV�լSbe9��޽=����4�%�A��7��B��ai���e=�8��n��j���`��c�:�7s��=��|���$���⽛�qs�ܽ���[z����Jװ��cǰ]�7�ї�@	�yt��oyzL�:G��h��/8�؂� 8-���>�@©�W6�KT�\��.��޽��맇��B�eOGS�}�H�u9_i�|�t	yw%��6/-{t�ɽT�=��ۥcZ�\Ȼ+9{'��ŧ�}��wb��p�o�8DxM�ӹ{ӗ����޴�ׂ��n���rq��/�wx�Ƀ���Ce�W׏����y����^Q7v��՘���.m�ku�L��|�ŵ���ާ��|�G���@�ou��D�<=���=��J'j�gŭ�G�wA��b�����8U�eQ���0�?¿%�s�ӊ�����Ⱥ���"�V{^��<�q�eu�1���ổ���P!�K�=��}⚊�<�Ct�����X��+�Xt��{�[\�������N_�e3/���7˶�_���^ҷԩgt=|˸�|2�g|0N��7�����eo�P6��s=��M��Z��5R�*�1��6������}�	�t8fXHȌEx���Q��ٺ��94���=�b�&e568�^���� q>��Ǹ��Hɽ�)@��GyHr��ܱ����d:I�=Ћ�|���:d؝�ޛ�!�pښU��R.LI҄��2��n��ƷWek�oxM&q��]���u�I=�:ćOec7T~���TY8�F�V�U*�J�j��iEj�DE��-F��E���������iUh�ZҢ���TkkiV�����V�PD*[eU�2�e+%��%�kT+[Z�F�����+"Ŭ��J����Q��TTe���9��4��֕eR�TPZZ�T�ʊQ�k�2()lKq��m*
�Y11ƶ�څ�cbԨ�[A����F�YjR�Km�E��K+J���ZU%V�T���b�T��0`�m1.[S��X��ԶV�Yi`���*�,�j֥e�e)kT�DmU
���m(���(�"�+iDH���#Z[b5`�Kh ���e�j4�� ��Qm�P�Ŵ���-�T("�R���r�Q���0��e���(6��(���#�����"R�jZ��QT���Z-kR���[em�Dr�S�Ĭ�U�����ѕ[[
������=PK�گ%oS�wEه	"�+�պQ8�p�����uK�ݑD����}$���f���慂7cğk�ʢb{���yAbe��o���ޙ��ќymd	��f�j�=�����w����� ���Q�f	F-�fn���,F�k����8Ɍ���^�:��gm�ϻ���;VLBh���˞��Vm9^wt����3����P��17�ᘠ�zQ�κKb�j�n�RsI���$ⷩ� ���T	!�T%O!i��iN��#1�� Ra@q(�'���Ӥ�bl���;3sդ�
̧ �	����#3��J0��.z�͵7ڷa[�U:�ĒK�ު�.��{H�]P+b�Gdd-�Ú-Ӝp��^�.�$dX���%��V"�L���U�9_d�}���9���}S�3^%�Q��j[0�p!�� �Z.�L$ɈC�%�ۡDL��=8*��c�:�>$�Ϊ�'�˽�(M��6�>n���|ku����l�Lk����z:��6�m�c���<<$ᤡAp!�]��0X�ox�^9���� �w�T`fE������s�	!��ЭF���[q��������n][�{�A�:h�	7�T	�UN��2$.=:���LP^������N�y�D��n��`�B3����$_����TA���}��b�)0�8�D��ǹ����M�n�<Iy}�D	���[��.�2	�d�9{�@�X�;iAJJ�Ys�D�A]�����|�#�"�A�]��Q ��ޡ@��ώo^��{u.�I�@֕�M)��G
P�V��̽���Y=���檅<�2�[�C:��ɜ5��:���/z^G_��*�G��8����h]�����y���`A�W� ���\�<Rm�N�٪�=X:�{�k�^�6�Vp�����gp��W<���k��m8��vŨ.&_P���ۙ 磱����Pm��}�q�P9��ݙ�c��X�j -�\�c�L���]s��q� �<�Uu�:��r��˴9���ѣ�X��a��:�����D�'�Np��ղp���ꞎ��W^Mp՗�]��Z�tθ�Ln��r���T���N������`�b�(}���Т	��٣���ZP�d�c�!>�n���J"&��4H]�ڇ0X�n���'����j`pӄ����$D���$-�r&�M2�m�z2;U+�-v"m��@~�͹�A�Y<�'L���Ğ���LNwO���H�E�p+�ꁽ��8n3J�>�	��rD���w�u�3|�_�a�D���^'�̧e�	cH�KB��  s��L��6��>�t�'�t�A.�z}4n�s���
�bj�V�˵ڌsi�z�	$ɍ��t�m�s�- �@j�΅$a��-�-��	l�H���Q
����r�����H+^9 ��*��& 2����sGlMCȍ+�H���ڈv1c���{
עx��-�ҹ��շ�K�q��ۼ�M��m���/n�\{�.^�hL�Nwo��Bv�Q���z���M���/�!��UMY�P��s<�*�P����0X�n���1 �����'cI��V��}��	fK�A�{�B�v"�m� �S�s���v4ܰH7�|O�.�v�	=�O:w�c�B$��$�u)�}zP7�]TI19�4z!�t�qI��bI�y�^�D�u
S��3��54�ҏ�]�ݰq�n�`���[�\�a����<�ڲ���'p`0�x�v~��KG
_�-��@$Y�TI�VuQ�ڡUgg"!9 �m9 ��gM0`���
,���2��m\�5.jL޹ �W�5�uoUH�؈j����zwX-���&BKy�B� �Wl�vu�M�P!M����7�_#8QS�����a��HdwWǃ��SX������V+fU�Iij����|��j�:�����6�����0�uF�1�0�wlf`�����G��G� #�?~��γ��e@�P,׽��@�V�H.{����������ѻ�A�R�ߧ�|(ߏ�E���C`�b
��N���6u:�R+%s����d�:�s�t��I�u%ag�>Xu�H)*k���Τ���VKW=���ݛWۺw̥�r�Ɏ���5��q1r�8d�2���ޮ1
j��_x��!������fk��OP>J�����XjB���l�A�R���w�� DP ��x�q� i��3�˟��� �Pם�ݝH,;���չ\�Y���i��;��a�*&7�aɽQnt|+���������Ȁ*T�{��:��*A`V�����Txx,r/�e�������^��ϏٙisC��� u:	3~~�gS�ed����}�vq�
$�/��h�����V����|8|>�bk���Τ�d���es^����v
�i���)&t	 P!	���>�b� �����Dx$�{Y"����5���
�@�D
ʇ}�O��|�2-�Wl}|u��K儴�8U;o,�Ů�s���ǵ��s:=�t>�������kof�C��'	�`e�����^!W��%�\�Fk����{�ρ��D>����Ԃç;������4iֹ��
�����pa�%�5���t�Nlty�߷���T�����bV��\׺�p8e H�'�����Q�ٝ�q5m��H��~�u҅��]��Y3�.�r��C3���. �n��ϱ�~}���뎆�M�=��)�ϼ�͝N�
�2VQ���>��2T(��D���߽���Aa��y��g��ԝ�����I�+%ed��oϷ�8%@����x~���uè#����Q�Dxtk��h�� ����$%!Z������H,���{���v2VVJ�~��s���:o�r(��#��,�*i b�!���q�u���� ��
�_~�ݝgY(ʐP7�inz{�Ǯ���}=@�D�
5�Z��{��R
A冾��|,�o��lD$"L�N��`�7�>�Ժ���ߞ�7�3����������%B��Q%af���܇Xu�`@�"<�����d{ l����`J�����NFVJ��_{��Ĩ�s��C�̶��kb�Xk�y݇���HR�
���a�p�I2�`�W�Y���>
�������
�+w�>�8Ό����P����C�+��~����q����I����9��Ȭ�f.�gKQ�+�Q��WG�#@>�Vl(���`8���D���a�(M�D��
�� �.̋םu)���<<+����|z}����ۧ��W�j��p��X��Xz��Ð�[�g+�n8��ev���;v(OaxC3����;�F����7C��u�:�<ڝ�k���3x^�!-�y�7vݝۄ���$`ϣn�A�g\dGzs��⇎vH�A�!�-F�;�;6.��f}��s�3k�6Ů(��Ü�����7�#/o�=1i�(�vD��y�18x��Y��޷�f�v|hvRt<�R��=���ɺ��X
�r|�ۯ߿���g��O���a�+��<��)'�5���t�JʁR�_��~���`y��������5���i������߷��Et58�!�[b
��{��vE�`�������L}��}�5�t��2T,IP�+
k��~�:ñ�aF%O��~�ԝ�����|ӿ�ߞ�Ϣ�۞���π$��(ȿApH����J��?}�ã��R�<��g:R ��_��o��W��g�@R
~@��5��}�u����2T,C��߶u��)���i��k2�9$;Ϸ���ϏL���u|�$��+k����gR
�T��~���Xk�s~������?d��W���;�-,9��wp��l�����\+sC��� uY�>���@�����W7�L����;�>��S��@�<���ﶡԂã
��|��8��VJʐX��gޢ |�D�i�]�Qr��D2� D�s��n�c\�ť���<Z�Od��`�v��ٌ���u�����G�>n�@��� �{�{��t�-�+X���π$Q "}��/��}����齘u�d�
!�=��:�Xv�޾V�Ӕֵn�g!�a_߾�{*J���m�)�y�v\*1�ðn�]9'!UK8 �Y��VN}Wݻ:;|�57>��݌1�!��iKcV�,p����]�~s5�I��~�=��βXʁbT�=���Z��\߿۟@$<
C�t\AU@]_;���g��?f��V�Y�.kF�9NO?}�:�@�������>��FJ��
���~���﹟y$�%Oy�}�ԝ���VK\߿orpJ�g��Z��1�-�5è�����k�M��L��&
�/Y�Q$�~�9Ф-)
сZf�y�@S� G�>^!����Y��f�^����5�ߞ��y*}��l�IX~�m�-�k����L9W]��paRG� #������zvvq|�E���<@�����p�R�,k��o�7���e!Xk�<�p�с_�}"ye��I�e�!��$�jQ��cq�Ƴ���2�V�U���N�������7ڷ.���g?~�Ăϙ++%s{����T*J���<���Aa�������xk{�4��5���gR'`��_#�3�Q�����b	-���7�������7ӷ^�]<7�=��
BҐ�����H)�>D>��|,�ϼ��>� `q��*gj{@��#��|��N���!��8�u�A�~���8¤�B��|���J2�T��<�<w�{��yu���x��aɧ��kx���7�}ضr
�C�U��O����tc��P�uq�#Ks;L�M��;h������k�9����X��\ߟop9i���>���ïX���U��X��bxE���F�ϻJ��g��3��R���{8�P�*Aafw��:ì+
*J'���l�N{���9�8d�ed�+�߿orq*:~�)���n��@������l:��^(��;H�C�i!������;���s��J�Ybg�{���td��%B�}�{�Ρԕ��5�?��3f�F�Qjg��T5(��#���)��2X1��`��F�:�c����~��T���4��׿�oa�%B���{��vu�d��*�~��@�S�3��oYP����=_L�
�C��"��y��nz��?u�.T�����rS�7���ΧbH,�=y��|�漑w����P���RVϿ}�!�aXQ�@�~��I�
�YY<�΋��U����g����ϽD" C�NZ#���5�H,5�������HXZ�����aH[
B��_=9��߸��qVz�S�ʞ��G�>�#�~�������~�Ăç{�����r��:�Y�u�`¿�~�{�p���I��*��y��:βQ��P/���xu���F�,k�������p��ĭ����z�Z���%�\���=��D�}�_o<��o�c�v#��r���\�l�|���sKC����Ui�VF�m�J������ ?�B�����{�u����5y��5��n�]/ )�'߾�͝N��2T����3�	n��:>����r�2%a������aR
J���������������@�y������o�)�L�k��"��Dⱈn;fY����k3=9vv��2y�"��X��a8A�� �+߼�݇G�
H(o������h����s���S�o[��Ö�u�3�w����Y�J�2T,C���vu ��=�m��k��K�g!�`E��2��� "=]T��W/ G�>����u���T��w�@�V�`V��~��r��������{���V|�|8��E`������-(qP:��s϶q �����W7����J��#Ȁ��>2�7E���1ٔ����{0�0�(0�*}�{�Τ���VJ����{��P=�s�����:� 9�+�#�?Wd�ݮ����y������?l�e!l�+c�7��^ ��H� Gȇ�o��gܣ+&7�$��%B���s͝C�+
w���ێ�3Y���!�a_����8¤�T��}�H��>����Lc;T️@�k��~���X�
5����H<)K{�Ϸ� |"�}��;���$M�ӊA�I��e�Ă�����>�s���p��j�9���'ue����+�(�y�d�}�_!m/'!�n��$����=:ak�����Ƴ�4���ZN�g����dx�	n?4�Or��غM��V����c��U��
�/���i5��r���8������Z'<t^�#�:H���Y�G��9��޾~�)��N�v�q��\�ښmi���1�'۰�3��|����&�O�Q��yI�@1Ǟ�PԂ�7���m��ޝ�Ϗ��y�m�y՝�x�-/z�1lE����v������[��s��uȤ�����M�n#ϑ�'�j�sˆ�k;�8w�;g=�󄑞�k�N�BR�lۦ�lnn6e@��gu�h�ۏ�
���.�Lf�u�C �Y���Fcٖ�b��
"��S�DB��n\�����U��&�	�{*;�����bQ JQ��M����K�����"��!����E�NC���r�p�ݜN�|w�L��+�/��C��%;y�{�ds|���Z�ס˹K�e"s*K���N-�S��9�_ZmJ1sAVH���d�B�+���o,��כ��%�ݱpm�`a�k����T�>�+�:bo�M(��5c�}Y�Ȇ�F�ko�٠�Mm5y2�Ẹ ��?�q���f�=��X���scH.Go�I;ӽ��_o�E�����.�˴u�	yw��u
,�1v�:��c�񂫛�Ȳ�:ddv�e@�ۛ���7X��!��?�Ҙ��V�%�����V�V���	lm��������-��Xk
�DeA-
��T��U���B�(�Pkb�Kh�*�jhՕ�l�U���fR�ԕYRV�V��jUB���F8�e�m��j�ZQcVŢ���1����(�Q���nfe��D*�lZ��ʣ��*�DT��������0U��X���miVQF
�R�Y\h�-���A�*E���e������1L�KE���ʢ��i�
�E��Z0R�Pˆ�ZŊ���Xʅ�Pm�Eb0B��Km��l*V[E"�+�\lP���E*��[X�V�TT[KDX��QE*�n4Tq��)T��1b"��ª0���ԣm-+mPm�ڵ�lZ�-��m��1e\� �J\���6���*b�H�(�[+m��V����5Qm��eJ�XģP���j-��
ŕR��Z �Ȣ�j(*��J�[[e�F2�VW-r���U5׵\�.�8h�q�ƶ�B�v�°�����f��ݬ��b�l��N7d�[,O&;u�u�Qq]��uk7N�c;%l��%�[�rss��1뙷2��Gvnz;vfo�n{�;I��L��4��lV�hx�^�H�1a�&y\��Ϣu�y�+�q���^g��p6�v��;t���\݊z6�1�fqn�ص��t�v'���Y��k�t��W���mh�k���<[qq�3z˹�3۞��g,�㋕X)���y�J�ϫ*F#�7g���h��l�i6�f ����u�O]�Ih�cp�s���>v��vW��=۳��q=���W�'dsp]���;sjk����k!�Gb%���`�sĮ8����Զ��a��;[�O
= �v�Ú���V2�G�X�]���Ɛ8%8ظy��{GfF�k�y���H��˰]�&��Wq�c�y�Ǎ��6�l4t�Uz��w��-/�:�=����@DY����r'N��-'�[z�;&�tgI��h�ѝ�7u���Q�\���ڲ˻�	�N�vqV��s0��X�v�=�V���@q����7g^J�����i�0��8�ss�Op�.n�Qw���>�b� N��z�ƞ��{x:��9i��#�ݬu�(�(��=�h��	`ݎ�[�� l��lC�S����=n����������;���x��]3E�Vx�4��cf�>q���Tq�����$s���v��`����q�nq���:�8��q�^������W��=�N}�;a�����ܤz]�b���κ���6('�1�ltG=s��u$@u���fŷ�ݹź�<�ڻ+����k��K�>�9vI��u�y�/�S<ͻsN�Vu+2�vy�O6�hڗ��\�wnx���Mh�!n�9^�qx���"�7X�M���)q����&��;K[�`��x�=rs�x�˱�u�C�=�'
���n�9C�=���[±��m��@�^��B����h��qϻ��{�~<L`� ��Nמ���������pW����v���饼���>��=&콨y݇��ڝ���.�œ����9�@�ؙ����+�΍F�7[�n��ܻ#p�%�6S���m��{=؍���u&��OgWYq)/�^9�v�sǳ��<^d�w\r]R�:��6���v��_/�����=J�k���ar맗�[���BR��턽uh��o;g'6�LD�:�͸3�Lg�aw��K��5�K�ﯯ�M7Y�ZӅ� )�	<��<���YFJ�\ߞ�g#%B�*%au��>�:ã
�}�s�����߹��m'����6u'P��� ��|���T
~>�����k�Mp�A����|(�G�e��}����ٽ8����y��� �0+s^}�@S�O|ٿO��H�$
����������!�%a~׷}n�L̺\s90�0���w��
��RT+}��vv3��$ �D1�Q�`;���:8�8�+X5�~�{�����Xk��}�q���y���fZ]hunk9��$���,��nr���O��������fG*AB�+�y�!�T����|��I�kO���ތ�u�l��^s�orpJ�}�s����5na�hJ�s�ۇ
A@�[�ݜH>���5������5��9�
p@�P+(	��{���u���T*o����u%a��;�?yO��t��4%�檥B��\�wks8��{@d�8탶��\\;��\�?�����;Z�]iѫ�=H/���{� �����l�βPe@�T
}�{�����ŽB��G�<	�?L�	iH[a����ïA�[�j���Ӭ��f�/ )�'߿}�ΧD
�YϿp- ������u���˚��6��,���>\�˽�z��w�˯A���O�qW�{�x�{���zڨk�w�݋���3�'R�P��Α��e�!��q׻���(}�
�������%O��߶u'b���{��&�Ϧ��۹� H��U�<5�1ӳ�D�?{�Ϸ$�B�7�H�x"<	@�~�u�����yO
�+*k����u�+,*��~��:$�/����i��D���|+��w������]�����9�������J2�PJ�C��ϸu�V��\׿op�?oEP��M��ϐ�Ixv���Y� �7�k"�+�Y K��E��R,d�k�w���P����%揼�3�1 ����ra��aRPO7߽�ԝ�����W5��ܜ�Pl;[:P��a�>A�pe�()����#�8�u�a��vN�T���W���~�����[�V�@�+��߷0:5 �y�}��t�*Ak�5��� H����ɏC�X ����_O��_����%B�<�>�gP�J���_×h�kNy��a_����T�
��w畾_��y���gYԂ�D�����@�V���kﷸ��R��\2b57�]���i� �����Y��Z��@S�����͝N�����%s_{��d�Q%H,�5�������FX����ڌ�A	��͙�.fP��[4�\{j~6{��F_�u�=l>C#�J���0!�s�C��+
¤��y��ΤN��Q�����@����q����ʳ"�HG�;7�G�}���nm=%�G��ԅ-���ݜ�!iHV�i�����AH,�L���nb��׾p�� �z��ܜds����-�ę�{���"A�y��	?w��x�y���E �z}�9��u+�`V��~j')�B���y��ǣ���̾�|$�� �B�\Cl����p#��uk�P'\B��'Z�w8s�Tnyz?���ߟU�]�u���|�����:�@��� �k~��'�%B�+��{�!��+���{�<]��4����ݝI�+%Y++����q�ǻ��)��4�Æ�(��N���G�YDx=���ɽ� ggf�yH[HV�~������YS?~��é�*y��[��l��%aa�>��u�)�3�u�c
���t#$�%�V�}��:ȏ����s~������/���
���P6�y)K��߷���T���f��]r��^�Ȳ>�ĵ;�}z '�}�|���_�����*J�V��{�q �� ���G��7_=Y���@��
�e;��gsމE�_NX�Ǜ;����^���Qܲ��<o#i�ө�Q�֩����h7�7���&�$������u�����W����p|y��X[`��d`�|3���͟ �Dx$�W�H�����Ӄ��
ӿo�r�S��YD�y���td���
!����:�D��Jw�V�{;��X"LB�0�b	��P��M���Sn.��qu�C�w7{[=������?qpr����4���|���%�*�w�}�8��T
%@���p�D�7��.y�;�}�`�~�{���
A�߽�p�A|<��r�JkC���n��:��E�`����>���T|�n��7��J�IP�J�;��naхH)*o���Τ����<L�;��쮳\��(�o�ӓKti���q+o�n`tjB�����ii
�_?zk}��Wk������R�}�q�2T������C�J�Wݫ1	�
��
>�G3>����j7N;�B��"<	�@G�v����%e@�T���:�X�"�}?L���fc�P�H/ܯ��̓�C[B� ���%׀$Qϳ����R,+�o���%C���9��s�6��J��w��8ì+
0�(���}��:�H,��Ϸ��@�.�G6M?�Q�aC��z�X���E��p��g1��<����7N4m�9lx�g�[[c���:�qGW2%�������̨�?xx{ѓ�	Ɗ�A�$F��sv��.����m��Y������:������ix��ӻ�!�dDI*�D����]��d���=�6����wDi�n��٤�:1�q�;�nۮ���S.W��S��;���\��jӷU�ų����2F������c4g��ǝ����G�ض�`���$+1	��	��=���g�7N�=��nD�P�y�㛞/:��+]��g#vǦ�l7l�oVư��ɻ=d�j�h����}OL0u�L�R|���Ì�Ԃ������!iHV�+s���@S�Ds�&�j���>�9�t�Y��y(�P���}��:	+
{�.��0��-˜��pa]����aRT*K����{��C�7�<�g�:�P(����{èJ������{��H(�3Ρ����g���'to�2"�l]f��:�k�~�gR;++%s����d�T� ��~��ι���s�~����
������I�
�Y(����{��P:k�զ曬t�a�hG§��)��:�ܵ�༐��������h���ןs��������.��_M�ʮ~�K[�J͌�
��w��:�RV�yz.9�0ѕ��Xv+���w��¤�T��=�Ϸ25���^�u�Y�~��@蕁cX��������AxE�}>l ��q}��7�������P�ŢŃ���]�U��K���<nx��3M�:�N�Of���;���:^Z6���O��}���:�@��%e+�}��q��RT($�,���܇Xu�a߶����Y��������ڻ�dz�z��X��_����T>?e�f+�hZc������>�v=`Xԇ�ߞ_GA_F��sid�Q��W�tE���,��^/�CO��N�U\7ټ^==��^�zo��+g��^j� <+(��OI�˯�O6�I	$���<��R���]kϷ�
q�@�3�{��q���D���h���@�<����6u���3Kus��Au�{���%B��V߾�gFu���J����ֿ����*x�@ B>|(��N�p��JB����ۇ�
����b�R-�Ӈ�,� �:߶E�l_ˮ{��x١���W9Ϸ�
�V�߽���Aa�%M}߾���p�V��g+eq�0��������͙��+Y� �^i6Yq��x�|*w�p��HR�5�|�g:R�����c��^�
�?}�rN T��YS;��ngY++%B�k���Ρԕ��N�/�(=W2z�c�D[>p@�FN0\rї�]�ts���NM׋�v5q�Xw?>��ߦ�:�s[�<H/��l>bJ�Ib�}�϶v3��� �S_w�u�#�!f,�~�U[�����u>�R��>��é�t��&.��i���N����:���d��>���<�q�'�{�y��ɈQ%B��)��＇Xv0�+
������H,����V���̫���O�dA /���2��iJcèJ��߼�a׬
ԈHU��֞�	�A$E������>�s�'`dj�cq�٭�ڱ`���B�=��xOi���r���Gާ��W6�UP�;baaY�X�ϲ�!f�&'V��k���No_w�O�X��Ͼ�:βVVJ�C_���C����u;.
�!����g¼|���jw���9��a�AID+kϽ�ѝd��J�u�~��R�X������>��~�{��= �)
ß}߷=`"�þ7��$�0�p��N��(� VVJ�+�y��q�}����y�:�~^�ק����V����Ă�P3�y��$�B�VVK]k�}�8����ZY�ͪ#�Ϧm�C, �P�߉�5'T�v+sv{WvL;����Ep�赞�fL>����z�֝9�~6�Xo�������{�=�ăҐ��Z�rNM{�=:g�~��{�q�FJ�P���{��v$�9�����kE�4en����H��y#��;+��*t4�y��$�@������`Q�
5־�ہR%!w�=�S��5�F���y9>t�V���&.A�\�������ed�־�{82T,IP�$�;���y�׿o�<a�
°�(�߾{����+%eu�����������ʮ��)��u+��϶���~���VcR��y�͜�!hR��5��� )��@��g�{���g��g���nϷ�����,1s��l��	��r�3���^���;���i�eW=ϕ{�}�fm7Fy�-0q�Ѕ��������y����6uĕ����β�p��n��4�]w���~�*J�H,3����}g���f�p3.����� " �����A*A`V���op9- Ҟ	yxG��O���#�ۣg�(�7�3��X��ә��M5pka�p��u�PGN�W9��m6��?���Cp�_�ww|�<�l�AgFJ�2WZ����d�Q%Bĕ��|��C�:°���g�����r��`����l�N�+%ed��[ޙ��(F�(8M��p�I q+}Ͽl:��Z�����x}���|��5����}H[)
с]k�7�
q�@��3�=�p�:2T������ϣ,�:�{�4�|a�DAm�Ʉ���F��|�Ì*J!RPB���|�gY�J2�X��ߟc���yƿs�y|�~? {�,kƺמ�p8ZA�����~�:��[�'�\(��N�"���>�dr=0�j5�f�����>��� �RV���u�XV*���l�M����o^���L����?orr%@��~�qʹ�V�<:�X~�߾�8��jA$ s�t��<���ǅ�>�9U�)�
������w����d�?}�(�dy��s�ҿ�?e�Ċgd������ڼ=���xa�؉82���_׺%^^����Uyf;���@8aU��vQ��9Y3ö|blEJ8��������x��p���۪}h�3�sڪ�n3��=�;[7[�q ��/l�nM����8v�q��\tO4m�?&��� �g��;�K���s�<�&�u�]v�St;!�q��Aq�Sy�KS�^���G)=l��ɞP�ctnՄIH��{��ўxy�+�w[v�P�e,�3��#m�d�g���!У�c�O��v��l�&��]��+�.N.._���헐;u��;�v�"n;J��m�q����J�:,}����i<�����4��a]���a�¤�
������vtgY+*�P)����:�X��ý�����^k�7�- Ґ�5����q�0+g���2�GY���]rP.����'�����*k}���x�����R
�V�}�q ��
�����8�R'�����}y����a��g� ��!!�l���H�<��;����!ms�vq ���_{������?s��@R
p@���}�ۇYђ��T(!���:�RV�z�ژ�Zօ��a�½����W�3f{5����x=�|+f�E�u��T
���8�R�_�~��v��'�p�3���x��^^�y��ף����p�5��kE��(��g��VJ�����d�s]�����_���M���ra��T�7�<�gR'YY++����'" �Ϫ��4��PJ(����og�n���z��/^6�c���=y4�Ӻ}t���������W5������V���vz���h�Ͻ�ă�HV�+~��� )�
���w��S��i�����q ��d�v��Y��>:��aAB!��w0�¿s�����T��|��o��6�҅_:�l`�{�:�ŮQ����̍��؂�������{�GH;����n*�p���Ri8.ej���w/�I$��0��9���O�Q7�?�UH���A�E�O�k�lp��!@����:��;(Q'�$��Xߨ$��U�m>����٢A �>bUV�>l��8a�U^Q�4tj��m�$�̚�I9�$|�s�s�֦�!��U;����6	�j���bI�W{�I����=�kD���l:�	�|�	[��F.ko{d\����� ���]P:�Nwdp謚�F+�9���͊z���g]v�(`��O�L\D@l&3*�x�O�k�'�۝U�WN�ԟ4P��>��ʠ0 �k�3���Њ $� !'���҉�[$����us��gK	&;s��H9�t:Lu�x��C�A���bA}V�	;�f�2/��Ǘ�Bq�G�?/�G����XWX�����튘��Di���> h�s��t����M���_�B����	��=˦�G����^�os3w!�ͅ5gU�S�2s6ٞ�|�|�O,��=� �~�8�'���"tPaՠ��Qئ�r}5�1��C���vY��4��ҟ<���
n�S��Re!흿p�2����ffG�F&�l-F5U�ò���������$6x���uQ(�#�����ޒ8@�q�����[I.V��>��M�c�{�������nTo�7��]�p`q��O�nnY햜�
�;�^�3�j>�ϯmԉ���~�C��=0�!�k�4"tH;0�t�ىyY���J�z�������M<���w=.��{�d������/#~ý�����0�]��{y����������/L�����t�V��od��n=|�*��FX罳<�^��o��p����+|�c��
�Nq�ݱ���7%�f�Ne,�_�F�����m�����#���W�O��.��<���Ty^���x��ŏ�ڴڡ ?A���p��?��+�US��n��Y��A��<s�����|<�@7��+�R��X8(Q�okp�{��dC��zXy�?l�#;d�s۫;�?�~C���M��f�]��>��Rd�E��`��{�vS�����/��sW�t3�.n����凢�u^��}����@:���/.މo��O&���>��٣��hWqI���S�L��޹���k[�y���*#�E-�����UhֶڥD,�ZU�*#m��ZUm���&Z�cb����TT�J�eZR��-�ZYS-���E�+���EK[Z �J��++
��ehV-����fZ�YSQ
b,QDmТ����m��[[V�E-F�(�Yikr��ek*"6���Qm�m��Vb\��6�K+*�E+��mbԨƥm���T��Upj�*
��S ��Z��
e�-h�RTZ�ʬZ"Zmm�[YU�iAE�i���UF֭e�
���ګ)s��ժܱn�Z�F���-R�j4�VڐUA�ָ�(�2�L�m�����Q-l�ʊE�-��m��T��*�T�VE�R�2�KKX	E��b�������Th���jfc1�*ۖ��+r�*P��YiJ�V�Z��f$X��R�j��2�D��i��lk�T��?�H;�����Lw��Lv��F�r������evhB)���>$�� �LWfРK��BUl�Ê�(�]��FV1>l���}�WD�͚����$'�"A ���@���4znwDU�Aគ�~a�KȔ�N
I�:��9�-�.ss��g�3pm�:����ӿ|�5�&�ǯ1�>$���Q$�{hq2D�dZ�˒�םT;�&	." 6+���Āy�12����P���tA�ouQ ���TO���ѩA���牱�0�LCE��_uz�.�h�n�f^�toM�=��I/��g����I�P����&y��1�Bw=^�|O��mP>��yr��Ɩ�ܻ�O)��fu�:}=%E��@���������9��6v�c5WwA���9�;��d߀ʪ��7,�%���� {�>�Ϻ���y�E6'	�y_NA>+�\���u��L]@<g@'�f��C��'Ă��Ɏ���ܭ�<*+���S��Á���x�	/���c�۫Z�e��Żg�svYN���J���������l��⠶�ۻ�(���{f�$��2$fJ�;=g���H$<��H��B��ll�}��i�<�B�6�1�v��A�6h�oK�A,U�3�m�ֽ�푃 �7$�-D(���^� s��O�q�o&]�]7��Hy=�D�I[��`Θ��P�aUu{�F`�8.7f�jEU��H%��Ve����g��r��3?I�L�>���2�É7
	R\�� ���f��q4��'�;�;U�	[���Ϸ:k�lL"	{!�oNF��t���'H�׫��3r�s6��giKU0���v0���Y��5�+��.J�"%l�����{�Y��5�m'g�n�-"�N�V�q�۩�c��8쇵�9�6�^��5�9�I�^L�(+k�g"��uN�Uc:.��]�zg5v�k�kF�:�������5׵M��:y�pj�s��!��y�y����=2��\�6����0��LӬr7[�Y�3S��9��u��S=���	�x�z�-���;r[��Jj�n�m7E�W4NsnʏST[;�d�3Վ��h���u�-�mخu��p �0[$!���	&�I�*��I%f�n�N��-\Gnv�\@�yTI>fK�b���@a��p[f|g��:�&����ڇ��V�ȒA���IK�,��7�&.Ƚ��$N^�~E�6	�j���	.��Q �H}�8o�_r^i�{�$-�~�	oz��� ���6]{���}��750��>$x���"��t�WTT��x{�j�݀�Nqω����P�aP���I.s��V4$��*�$O��כU������S�#������#��;{�ή���-kts�s�۷�[�.n��s�s�3�vz[�_�~���Q疑�����v���j��$C�ꢣ��M8:V;Ù&zi���ސ����D �o-�&>���8#wp4��C%Fy<RnA�y�%w�M�t�C���*{���j>�?^X��0P��,�<�m�4�Q��手���nX�Z7^���{����N?�|^�uyG�Ӡ�┩mP݁ZVOs�|�r�D	���p̃;[t+��vhG�9S��]zk+cH$:��	����i�d�`�Fs��1�ء[e��O����$�k�Vl�Ȭq�d� U�d<�!`PK³d��d�
Ζ:q;�H��S�D�O��6��oK�̰�`�W�naD(`�K>H@�r���z����n�&�v�3��m��Փ�~���������=[�T|O����	!oL�Vϒ=�['�Y�m� ����`�<��%�7
	R\�9 ��8��Q{"#�r�Iw;�^$����k͎1H��zr���!a�I�ꃜ���B�I'�9kov�3��f;�0��:݉��Q��䰚ȩ�a�G�o��{����>#��әBdWE�����Ja�7ݻ��M"m���Q��<���������	+_�I��%����2g��;��*���I5�}4I ��2$�C�Ω]sOH���٩�v�a�"�P��j�o��	w{��� 𓙩�x�ͽ�C����s�$>���G[�W)*�IN�\un�'9���B��X�����	�=l�zˎ-�N��;��(AP
g^eW�$�e���GnuQ���c��r{��'Ă�e�$f3pPLCE�
��ޯPoB|h�}�8�p�gK1۝T	�Fv	��;o,�r�� �Q��nA>$�vm
��c������>�I+2\��H���x9^@@�p�u^s��o�]r�P$��$�|Lgg4��J������7��遭]f��MwVj܉ݝb��+��_ wfh����&BN�U�cP��J���D6�V:"�K��F
c+�����rLh;B
�J0���I~�٠zg4ռ/P9�*��	���	��ڣ��6��_n��+�_KX��H�i�J� ��G\&�݋�;�rpN6^�6�O��ۯ�����b��%#���$W�UH������y�u��R�
�Κ9#rKaA
a@�+�r���=�8H�
�rޒH*��h	}9�@��;S�=s8�qE�:��:k  ��������Gės�4I^�z�j�@Wy�����`�X�����N��-Y<
GĒ���x����%���BA}��@�v�W�0�14�W�n��M�>\��UD�u�+ľy�@��x���%i����ޭ�[����Q�փž���{�݋���)ۣ�rї8����{.oЮs��3�ȮH۫�ٛw�YUmQ��:���Ē����{�ߕv��k��Lt�lY#\u͕v�Z�������Ƚl�����T/;�2�m��pF7��?;a�`<Bu�rgA�y1��N���g�m��*��ӯ\�˲p�}mϋh9;	�-]�㵴���=���1��<�{vi�]:	���m۞���hie}�5�ݙYB�b�g��ug;�6�	��47f�E����Z���۴���I.]\�WV����Q�̚y-�\�:�귎L�9<WSʾ�D�^�����o����st�񝺹�^�٠H$�D�j"��Ḝ�g<H$=y�F�^��ڈa�#4h����ӣ%t5��:�� �K��T	�'�>���$lM[2v���s}]��"�-�(�ko��	�=�A'5�]����g�g�'��ݑ@�i�x�@AA1�n����ޞyz$ź�	�#<B|	]��y1�]�8)����~� ��ED�KMJ��qr��%wn��tW��7u�$PڙʢA �qҁ%v���2��w�Op.�����4mug�hK`�>C9W{k�פz��c<ݴ�2�I�"�Z�L'���u�9�U�G�*�t�A%n���N�H��VT%���'�F�T*��Be�3�=�sF��\�9�]E`��c	���E=��V+���JvF�fں܈ u4/P�oD��3jq~�uٖz��f���{�Q[��c�u��Մ9�7���<���ΒO��|dWo�4	�{�O��n�{��v_�4Y)���'�m_�>D�U�uDx�d����ٞ� 
����{j�2�%����H���Z�S'6��ј ��sj�$�=��8@�S1�Xf$�"�V�9p0�6��7]�T|I�y�@�����-ynk�>$�u
�>�}�@����I�ٓ��l"#�y0a6HF"D��BmϚ�=�T�ݺc��cv&��5��c�����a�3��;7D����|H$G>�
�.�Y�6\M�v�4�'�]۵@��9VB0�P�	�t��Ns�����s�0�%n�У�f�&�m.:�,��	a!p̃9=t(���x�A�+{���t��.C�c�	�#�ٜգ*���=���ר���w���t��d�v��:e��cV��&ҞZ�V� � ��#⳾�H��}�D��z��4���Q���hZ5y�=��G���j�>"#�����fE������!����H�ʢH���r��'�Sy��UH��
$�tt���b�캑8~�?��=�{���v�[7a�[�qbw�����wFۯi�Ӭ��x']���_ϻ�~�Ò��0T��
$�o:hA��=�^�rFq�n��
'���Q:�bT� �pQ*MOE�n�Rf���;�DH��j�>1!xƙ�����D�c�#	5�8����b.:B$�"�����nfv�}���x�tq4����a�6�������'�	G������$	Qo�G�]۴$�賱�F�-c���4w�[Q��5FU��5b��s!�1��qT�����hW���t0Dɰ�M����*�&�E}��< ߉�v��N��R,�iC��f�:|�%_���@Қ�]yh��ު'�(���.�گ�� a��Z��l�%�6[�-��l�rлt�Ɍ�}�w���ݳ�fu�f����4plD`63j���^+�v����ƪ�]7ӧ��l��7-"�(p�0���gP��,ZR!ou��9r0�HO^'ĭ�گN�iԂ��Y��\�_mJ<��T���ROE�@�ٻ4I��V�e�V̱(�TH����@���j�;��,Jj�8qU/�+���T��X�L��(��	�[��D�}�g���DNTL�"o��@�!- �3 ���� ��飔�lŧ��W�UG ��ڢA>��F=*��h��X���հ�Z�˻Ԧ��z�ܙ�:���)l���q3q�Fz�`�[���3�e2m<x�����}½���5���|�]�j����m�xq�E��m���1��
�V(���l�'n���N�2�fL���tBG9��7;���o��yB'KVp'[11%@�XQ��y�2�F���s��يY[kFI��T������&9/�Y�\��y佧}۷�L�8}V���2��K���n�;-�'7����h�}�hr��;Փ�W�x��Aݸu�F��k�S��3��~��G�$��d4�^�w�z�쾃5�e_��f���μ^��/Y�j\�s�偵����h�z�����~���,��m���]8Cۈܞ��"������|{��:m3On��%���dm�T��}0�����z����|�n��y�uCs�\�G #}����`-y�����b�5x�� ߺ�og]�U�Ls�o��))q����w7��i�GwP�w�Gv��n�b}�g{V蚝�l�˽v�$G�L�G�O�m.���w\Ty���U>\~hby'`bY�3chB�K����js+BŬ�9�w�p�����U�;�+���:���bL~�*���{�}e���Bށ�|G��<�M��7AKӰt��pͫ��P{�n��мH�9�f����!��_;CT�~~�P3��'�����r�����q�w(:�n��{�G}�P������ww��%U'"�^�/&���k~�@ uzy�`�����J�X�YAaR�jڊ�J��R�0[j �
�q�Qm(*1�e����*V�YEk
�*UQkkD�EQ�X��Y��ƍ�e&2V#��̥�%KV�j��TE
�ň��Z�kZ���,V��-J�R�JʢXUQ(�iR�[eS,��H�cFVV�V.V�2X��QH�VPKJ�J��-�"�,������,iaP��j5hVB��E���ڴ��5YR֐KX�Z�-��YZ�YE�-T�X�V�PV��Z#
[%�UVڴ��X��EX,D�����eA�[m+%H)UQAKlTQTB�P+*,TX�Kl��)YR���E���mEX�ڶ-�Z��U�mV(��Z�Q`ũF��ZFeE"�1UE�DaR�Q-��[�j("����0EE��J,bł#QT�%�bԨ���f��|;��s��O=ۭ;�v;��YC�<�q	Ϋ-����ɢ�R�v�-B�;v���xyx��tml�80�8ѵcl��@���rB���m�Hэ��X5��sv���ɣ��8��w;��;��m�����s�����c#g�v䛘:v�^�h�}�	�[Y.5�7c+Vs�l	o'O�������j�	6��v؎\�ӻ:`}�h}"*ۂ)(���o���������/n�u�]q��ڎѮyuӕ�}i�'�]��%�mӷ�^���m����g]�����/��-�9+l�s�Z��1�,v^��ֳy�7m���u9:�z���	ں����2��k��aݞv��,|������]�B}�˕�w[���cq�p.G\ܧY�U���-��:h�;�S9U����;y���)v������{-����{q�]�i�Z;��S�x�����-=��8�u;f�u��v��틻}���m��u��\x)M�ؕ�{nr��'��f;z�jØ�'.f�q�a�F��{�^c�#g����vF��ۮ���ݭ<�0�1ۜ&��ۭu�Z�{+�ql�ј8C������Z֫Z�y����n��n������z�U�ȂV���J�d|v����=E޶۵�)�8�iw�q��=c���'7H�+�F#�oU�zgw1��YN;8�8�� �mӮ��G'�lf���[Ѷ���۞y�vr�׃����<��;���Jȝ��kq<�oiyֻ#*hi`x�6�g�����=��5ء�Y���6t�#��<\�{k�^ٻ�	�õ�B�=�l(�o9�	ͬ��H�s�@���]p�m���92۟R��'���ûr���^z��|��(��C��V��혨��Nu�z�!�G/f!�a��q�C�1���y�;b9yw^�E�S�u�k�m>�H�窈��<G&�۲\�s)F���K�gq�q�T�Rr�.9����׷F��i7'A�8���;���yo���b��N��M�V����7\�u��篎�.n�w=���[!m�R��8WSR��"������:��p�x�u�T�n�F�kW4�h�uZ��x�k����W3�ku͋��v�m3����Z�w)��0g�n#���8�6Tx�'��%��n͎���z�;�u�&�v:��)-t۪�@��m�ӭmT�H�3���u��=��۷���ï]�O����<y8�h�7vͭ����O�@eC��u�O���t׈<�z�H��C��,<��H]��@�E����&�1>���5I��;k�&����uz���Q>(���~���[dvZE(P��!H����-��� �
X���{8�B�����U}�Q�0�P���%I�軆*��Lm��Y	&3z�P$��I0�:"*��Ua�$ M]N�;��D����jM�L�7��3�r��R�5���T׈>�U@�]�#����]�q���!��m�0J\{]��;p:BE퇤�sp�KvRq$]�ؼ��{~�CZ(BL4�ٻ�>$}�4	��w)��&���Ձ�;�D���'���b�lG�5F�_N4V��N����_ڟ��rˣ�?f����_lB=�:�hDѫ���s�h`�'�2Y����*A�{˪�hò�N�fnS�}�K�Gn��� W��� Fe}�Mצ��Ӎ՛Y�z��0W�UJe��4�s��`�vv�� ؂5_q�����؎
�[�����ڣ���TEJ�ǝ��s�y�)Z{SWE��W�m����� �J{{�.�B�&Q1��=�w"<怢	�DC��f�ϐ'����x��:�9ԫ���v��vn��)���ă�v�r��Ù��������ݕ�����q��3ͺ����֣[��p[��#�9�շ����}>�[�2�!M�/�EњӠ"	���ς�/���F7��:n�C�/){H�X'�Ƌ%I���=�uD�idVQb�9�\�s�w��dC)���π��kȽ�����7�ɚ�Iz�<X�B�P��7�<��� �'��x����+5#>X"�y�}j�9{�cE�ܤf������F�����s8��j��>ǽ�l)0y��kͅ�æ;��;z)E9��_��x+�ޟ�H$���nH>���٘�[q0���S(�U$�[�9�w�~	��|I'���DI%�޻��H���U��$�O��%���($a�\
�A]^��$���u0:P���Ǥ��DW�����>	�w7����fv�،�ʜ��Rd���+�ןQZװ�^��s��\]]u>gƼ>.�j�Ո��&���'#���ʨ%�w��ϐ G]�va���^��E>�6��	����j���d��MML����;�����N�GN��,���I�+�!��d�H!�=RI0�l�d��<�B^����e��i�3��Yi$�]w�p�!�7�.���ʳ� ��fb .���
�Zz�d���!�y��kWN���d��@ ���0>�z���4 맜V����3��"k�^`=�G��n��t��>��jMԈ����:�{�r�/�-4�[���Mm�s��� e����wi/��PlL�QT��?���6Ȁ~�iώ��Mmڀ�~���  ����D4:��B��Y�7Ƴ�b�A�f	�|�aDD0�v���x�oQYw���I�.��⼘Y8���������"eR�NG>�f,"�}o� �cA��efFV���vo�3� ��ZZV������%�ѕPJ��Bz�=�o��� Q�v�o�e^It^#�Pmb痩/n�0�ԓ/	����%���@$�W� ~�{�,�ǎ5�v��� ��m2�t�	�B����S(�ECh�y�/H��!�Kڽ� V���D�^c�]���^��U����n��z��TL�L(��O7"@ �ws����A���2�w_]�> o'�� >����A_F���Ox�9fK�hU]����%�q���2�2sL��Sy�o\�4��v���}�=����{�+����Z�g��������07;$Y�*&�� ����P�B`2�L�d���}n�2{�c��언�^��Fۮ#"� ����kۃv;�9.zu��I�i�"���{\�p�N{v7H�͞IL4糛�ϛ�Z�p�nU�S\*]��'[���r`�m�UӤ�>%Kg��Cu΍x��Z�N&��z���Mɻn6�K�v�	΋�[�z2Z&��]G],�b�В�g���v��d4�$ok%��Ϯy�w\�j��e�䦫�5�}�����z�L�H���Ǿm��u� ��٘�m�����l��o��ԇ�!o�A5$L�P1��ێ3��:2�~çou��X�˜�A*���� ;�٘����+F�֦g/�#D��Plj),���PJ�Q۽X�DW���ܦ3��M<��@$w��@��^���I�c�D�h0M)�����^��!��ӑ ����π]��[����ڃ<Ը߀����Ԃ��[��� �EEP��?,�@�m���/z-���7�uoP_]k 	�wf` !w[m2��ۛ��S������%r���{u�1��u�I�><��j�uh��(d(��Kd;ᚹ�		� ���r|ӑ ���� ��۶W����O�@u�m�$��7�(z��b!B-���ufT�Jz�A�g-G��,�NV^tn]Nt�e���@Z��w���+D�b�oΕ�S����v��b�-�~���'��k�����=������ O~���b]��@����W���h����.~@�h ��Fnv�` �n�a�S������<���x� �}��Ȍ�w[wF�P�k�XA�I�'+���������Q�8���� @(��w�o�����:��Rd��5U�$7��(p�,�p�B|��"���ӵ�(H;�̈��۸��7����ť�wm�����{R:�C�@�_�A�������2k%:�r�4!$�W�䓫�Ԙ���߿���|QS���sٟa [���C}=dDg.1Gt��m��sz� ^�m��ᒱ�7 ���S�B�y+_�xS�@��מ�Ǐ����@$����D�P��c�D�-��&���츚"x�z�I��$	?/H���a7��:�쁵�L7z�V�ߚ�7��Wa��3��n^;�%��^F���h��꽖���i�~ݢ)����U��Q���ӱG�s�{��n&�� [�ݶA��ӭ�|�B��4���T��v_m��|��ܲh��2��ט� :�y��PR<UBD[����v�"Dd"��MDE��<� =]��j�˷��v�|�g�O��� �{>nH]���+O^u����P�,��& �*L���3�v�rn�e�%3���ŷUn?����~���.w��0@$��Nb"��{3z<��e䙄B}�~I���jBp�$Q�	7bz���I���25ۻ��}ZȈ���o� �7��6���`�ղcDb�b
Bm���	e\m� ����D~�y�i�1��� ��u� A����@}�{"&�I��a:4�veG3:8SmY,%�QR��/���� ��m���brj��K�sdT7�;S���s��+o2���v�W�ʸ]��a�v4�&�Q����u�2R�5��d8j���*�� �O� �����-!_�P �&)@�w�߳0 �ݿ��j-��v�v�P���"V�fb�����90���M��.�w�/lu�U!�\��h�l���
ֱ�jy��q�,~�ݻ��ѵ�ѳ���月 �wsq���ݴ�.�=6�T	��v�Y�NW߿[p��.`Q)�J*jf�g�� +��nlE�Dת	%{�w]�H�&�W\r.VfHؼ�u����i �AUUSe>�c�A���H�{��{x�:�lVz��e{�3 �w\�'��>5��`"��pɘOJ�Mʹ�l�,�w��1��� /m�����mM��8����q�y�MD̨�)��y�?��u����Qέ�8���{3"0{��� d옎���+����x���.<Y[����O.^WD��`ي�쮛.��Ļ�\��$�P�.a�3,f��5$��!�[�e�.����
� DV(|܂��"�m|�n3H��e(I�e� �Ӻ��y��b����c�sԽ=r�����Ϟ91j�z�Cf:{wm����Mjt��=�/h����|���g�gu����v�vE�yiڧ�d���8�yKE>��G�*X��wD�p�P�h��ذt�[k��n���j��v
�mq�h�	ܗma6黲'<�wCC���ض�2K��Ϯ��l��b�n�Ɲn�sY�l�K�����n�!N�ŋ�-���f����69�yq�^m�L������ ��&)A��F���� .��i��}��0��޴�9����f ��۳!?�D<�d2�(L����o"'�,U���~�H���n�덤M��8Ë�Y��r�%�BD�Х%K���~` <���N�&�k�e0�~�@ .�m��d��$00{	��3	�Tuݗ�Z[�Q7u;�y_�'��� �~��D]��g&s�~f��}�m��t�0!�)6�AM%�q�*	Is��Y�~r�ު��V�'w���!�N��)$�޻%.�p�X(sGt3q	J~�u��/�mYۧ�v�ym�Î����rqے��>0�!V���1e�����������^��ND�����Qj'��y�z����l� }��FD+ւhj	R�.�λ�KG����"*�&a��d��9�E��{n�G�ow�<�k��~�۠��V���`z~�¸��m��̳�0{.�������J��R���IV��w�& �V�V���]_��1 �~0"�T���n?���=Zi'�QIe�eT �8�����yV�^���t׮��o�[RA����1j�!)�J*J�b}��}v��6������r|�{�1@.�o�<�I�i O\�#��L��!����{.�h�C�jZa�E9��1� w���� ����	/$��������ș=�v��Ae��v��unݰL[���n4#���`ƀ�� n͙*�^�f8&�),%���BI���ŀ V�L!����e<�A~��ob�I-}�wa$�(�eD3�K�������fj���{#q�~N��>���f ���ݐ �K�*�ү�����<�=���	�F�ʾ�K�>Es������>Uu[1ӣoC��\��T曹�oŔ5ܣ{����<L�8�>�3Ǒ�R�φ痆�������7A�n��=R^9#��2^����K:��-,���T�C[�f��W>z7�*�@C�	�5���殭Ł�;p-�g=\v�ʸt8�Q�y����ص`j��{�>�XY�Ü����;.���}}$��,#x����5�&�x*^��sF�r�Ƒ8��k�l#{ݾ��\��������=n{����S��W�`^���٫ץ�'?eǃ�$���'#��ħ�@���wC�{W��{����ɺ��Z�YB�Y�GH�y&N9��bpH�g\��g[ ǃ.����6���[�BI�o������#��\'���î{����Cw'N:JR��zZ��c�(^��/C	�W�}XU��܋�W0Mo��L69�l����:,�
��1�6�>��fC��1鹻�aQ���ʈ�;��P�kk�4k~")��!��޼��[�K���7Z𢼋���o����f��_'�S�����ڽ��T�L��ۣ���.o
;�vy��|�͓V�;qxvM͋��82���>�}��=�o8������_n�sΨ ��B�>��sR^�$��˹����uW��L���9�8����w���۞�R�6���|0���%�Y���W�e�F=����0U�z��os^��T�^Z�sN���Y����78I������\<g����x)�������1���]���yǞo[�a�3��zʨ�*��	l��$`��"�aFR�Te��J�Em��*+mE�1EX��UV�,��[eJֲ(�)Z%�Zʫm�ZQDV%���Z�R��2�����*�j#R�Z%J"ʔE�Z��Z"��j)Um��TPD����lP��m)m�������JZ�V�TAP�6�Qm+���"
�`�H������(Ķ�"ZZʨ�ֵ���QV*���*�F�*V��I[�b1�*EQq��(�Ĺ��\��DQ[m�F�Ee�2�F#mX��X�j�J%j�AX��Ŋc`,m(V堌����l���j��EF(�)YEQ�A�������61��.AL*�"����Z9j"��0�g������[K}���� > ]Z�L>�\(Nt��&��M���E�w�d�` ���� @G�����|=q6I�:�:)g�8'35�@-�NAB1M
PQChO9������麜�#e=��^vfb !O�-�@�/��b�.f&{�WeO�*�Q�Iܽ���9��t�*s���msۍU9���ĕ��⟣��xN�X�!��嵗�v�$Gm̚�Ix$�=���3��K�5j���fb O�ÞU�TJ��UA����=F�Û�l?_��� O�� ���D�O�S��ۺ���MA3US�\1_g��H�ۖ��L�fԓ	���y�T���G ��m&@ 㞷a�'�A2�#	T��/wLvc�9Ϋ+/;���f[`�@��n��$��뼵]W֡FHt�n`)D�6n�!$�Owzs��{���^�܋�f޾�-������&y��J�Y4VF��r�f��W�b1�����	 �vuW�#���٩�&��M����@ �]���77j��T��@D��Î}U(���������:�䰘��2�C���+�Nz��u�t�5N���΃���:��_�삄j�����	�lD8ǭ������=sS`�Ԟ��k��=�d ��I��<�BCA`7T�:�=�"0�vn2��ҥӿ0 =S��Hs��	$�8���7���ߘ%:�OT�hPQ�l/�� A>�sϰ �ay}���B�}yd�AT�ʠ�I!��v^/@�&QUTE)�\��}nY7jA�w?�� �{��� -���ˋ��M�U7z��E�޹���}�"fJB��F[�{���]��&b�*��A}��u��1����� ��m2*�~��:p7�8�sVi�v�KLVF�9뵶 f�njZ4�;"^w
oN�6�C���E�9�Х7����	/vLj̥g\ӻ"�ݪ��
_Z	0���BGJ��n͵ӱ��ː�.{)ry��3��䓉7m�Ѯ��<�E>M��n2�v-Q.�7n�7]s�[�d�Y�pZg������X�6p&�ۻ]sU͏�OVx�����	�v��I�ux(D���q<˘ݱ\m�o�ה=p�+�\t/cj�'�1f�v����<�EюS�v|A���@�Pt=Bu����ڝ;�s^���S:����p]�mu=�}�k�ɳ@k���}�zj�&$���� z{�:;���%}u4J�#���dd�"�H�޻&���A�	4�7�>���)�����f���� '7{3$F���R$�Wd�$���K݈��	Xc#I�d��P	�v]�H$������c���So�yvx ��fb@|B����U��Q4(
��D:�WWT���fI/�]�e]�RK�+��� "�O:� ͜��vm�ܾ��E��`J����%L�hZ�ͦ �ӭ�:��Ϭ�>��vdF| ���� )��rA�黮�+���"T�q=���{mƣr�\���ڨ����i1ך�S�o:���npH�Ba2�
�˫��� ��K���"")��� n.S��ה�=��v��Dk�4��F8n
�	�ӯ%YѕP���j^赝��'3Zy�:�Q<��5�ږ��u��w���o*�̢s5�O�w��0UBRx�Mp+e�}�i���n��M��'���d}��T~H�c7m �*�O7$D2.eu]���؉v�0�U8��B�P�c�0���i���\z/31_�;ٺ$#���H����u#CҲ$\�ꩴW>�Vt��6w1 �?=��$ }Z��ofUD�U�&����	�\z�L� *�%�c�����{���u,���*���v� |WU���w���x��䍻egS��z�\�筯Vvٸl/����\g���p;bcpl@����2�y]���m���<���I ��'lh���vf h�+ۥ��b�5�jȈ+ru��gϱ$�T�e6_߬	I�8�J�������J�+X�"w��� ���"p���gN��F8nB�~4ɞؼ�I ���` �ܜ�b�O�)ͫV����ޘ��l�,ZR�6վ���^Y7}Vwۀ���~Ð݃tn�H�w���7�9�u�ɴ"��MĿ��Vmm?� >+�O7�� ��vf|��ȑ�B�P���Fǲ7%�h܈���m'1 	O���� =x�gn��Eδd$�٘��HX"Jj�-��*��� ln;iY����kf�_.�7k )���ĀA��u�I�1�s���r�=<N����[o\�`���n�g���V�g����?����?��x��G��O����'��� 㱺��CO��h��e']T!䗣w���@�q�4��J(ׂ�y�BR�v�ʩ����1 ������G�$�H�{�3{�#�[~G/Ӯ	�"*Bƌy��1�Gc�����y�������O$�v�]�~	=sff���>��6�%'�����;��b�ދ��}���` ���=Q�J���1Ep��a�7�8�b������%+�'V������̓q�qiV�EN5w�.p��"[���\�3��H3j
i���G�K�5�wa$pb��D�DAQChq��������c}]��9}�<��o�+�;�����:7Y���jE��x{}�u;���6+�Ӟ�l�O6n�n�V�.�O]k��. 	t�ms�sn[O'��~q��}�s�?J�{��#cq۰� ��'�hU�˕����$�÷R� �3�F6�S�Ch<�zƂ�>�N��\�����;u��I%�n��I}QӐ�	?Z��ʬ�kz߉!���A��`j	��l��D�,��$��!�~om(��� ���m�d��mH(�ϱL�BpAq
�u}י�`�+٨�$N����{��` ����b̼�/�j��'�&��>��A��k����"'���Mś�/s� ���Ԑ=�٘��h����<�E�w���W�w���KC�m�{{پ�i#��a��bר����]�;�8�\��D�^c,��6�t�9^S�B0�nc:1?�c��n�g�cP/[,&�g5��v�n��A6{kc���'i!�v<�Į �ĝ��ڮƴ�D<�h�䱜8t݋<en��QO;�� �#BqtR��OXNgC�J�z7-��\A�n���x�7]N��!���6 'Wm�gv�nζ��J>�9���>ю�[���1���,s�r�n�p�K��=���|��;�P���"4つ�Ɛy�f��k���>@�%];n��^;94omL$s�����w�E��Z��/�� ���� A;����w���j��)��6I�Ϳ�� �{��5�c�,�i���n�uu�HIM��i�k��@ /��� �wf`�����j��K$���K��g1�ӏDҤ"�<�u�1	�o<� .���\�:r�@@#N��� ��{-��7�;$ h6AƠ����/���Nz5�%��"	�ofDg�|z6��������Ͷ�ݏ =�ڐH߯lD���%���vV�%$3������ӯ3�S�l�i ���fb��m3�:�Î�̎����I�D�f����&�|嬾��gƃ9�s�Z��V����0�C���J�(T/$Lvo<X�yv���-���1��=~ʪH�����s�!n`��:��گR'J��3�u�����j^mU���O�.���ʯ|r]�V���;p�W�2���ʙݼb��s�'��KF�u,��n�յɀD	O{�3 �q�A'����"YJ��˟�{
��̑QEU^��;3 �mn]�C@W�Nz.<�z�Ѩ �of`D!z��M	�=ƓqP��K*��?\����R{}�'ל������ U��*gf��U�В�9ܻ���De ԚCs2��+�:�uJ�=�ر�#Wn��0"/V�� ��M�%\�t;�}����6��tY��t��ٕa�Y1ϧ�u��(u�]x�j�����{A�D2�B�wO�I$���f��u����^۱y���4�72# 3��HH�_�LM E�#�N��s!?`C���|�.����ϖ m����U��^	Etv��[T�^��'�@sȩ�JME�]O�တ;Ϋ��p�Y�b��cx�	�ɁQ����Q�50�]�����nFN��9�~nD���׵�e�wY���Ԍ�y�
�eL�#�K��$an�@}-�Y�gh��ཀྵ�o$ [\�d |;��[�j=$�*"A��R}w��N��
ܵ $$=�o�D�� ��߽���#;9�!$�nUP�: �����[�"�{3�����av�^���:����!�u6|�ofDcȘ������7l?}1jH\��<Z��ص��'2c!�q;��pH0��Al�Վ��@!�&�Y�'��a�v�� ��ݙ���'���ǐ���d |;��=��bH"�4�,����r�9�����0A$�nH ��sx�mW���n�ǝ����~ء	0�?t��z�'���b���۷� }��@�
{�٘�U�#�L�_ETQp�{w�Fz�h{+�����6 �w�π
{�먪�VX�br=k��?��s�`>bq�Rn١f�}�{9�P9��C�1��Q}�����nay:�},�m��^^��qǀFg�6��Hu̔**���睙��g\שtےWA��'�q�В	/���ϐ |)���۔����=r
b��	�wk�vg5�c�C�iMY��<��{�{\`7i�J�wY�fi��G;�u�:�}���F >���q']��;s�����s�	�wo]�e��(DBi ���_��[��������L @%>���@ =��!��E��=�5}��+�(DA��8�S���� )��i��L�=~sf�zDfQX�ӽ���
{��������M E�#���4c�q"I;�}�U��@%ݎ����y��C˞�i���������aO�5��١��=�� >��i�q����L�ݠ��٘�H!O�-��.�����8xk��ʉ�����M�e���$��3�]�k|A���:̉o�[�/v�ӻ��ZjGnf5�rF1V�1c*�T��+햘�S�J3R��@��B�1ܾ��4�w#�r��o����<��z��1��t�~=藦���<K���T�,�n1�ַ�����{��7ϛ��#�o�]t���G�H;�9���yز)�h�{��{��>^�)~Y'�!~O7�'i�]S�}6��u�^�؂��s�����&���L9���l���S��^��N�T�Y���c�Sx�m@��N�����!���_Z��x� �ep����r	.��*�z�|a\���]Ds�dAّ��;���{)Z5Xs�<f�s�t�9�]�&���֦����=7��9<=��]s�6��3w�N�vzcZ�/v�Uy���xx�F�Z}+��Q�{%4��4���T��!(H���k��	�[q�)���.j����N"^li;�}=��;�ŝ5pmx�@��[-����š�[5��u�z̙���\��g9��^;���������{���w�5���!��nN�d��'��aլ�ʴ��1N2�3s�I��u��W����}���)�s��4�o��{v��●x3�¾�}�{��3��'���􁮙�=N�^�Z�
�+3u�@�3�AWh�	�L!4�$M���1�#2\�y�!�;Ol�P�d���שY�������ѭ��L�G��5�O��ݷf�1/������N����֟#ǽz���!ۯKY�ALc"�ξ����3_��KW��Z9�Ӵk6�=�r�=�:۾ne;]e�2�U�-��X�r�[F+iY��.	A��"��U�V��DV�p�G�,X�R��RҬLpʕ�.e���&6(�R�V��"Qfe.U�b�Y��V��.Q���̥�Kh�-�1R�P�X��Ƣ�4T�**�Zd��Kc2�ʵPb�s1ڸʬ�eeIm�"�Ab屌1�QEKEX%j��J[A��+--H�*�eh�j�D��F��U�G)Kh*$Q-�V�"�nf�R����2�Q9h1�r�"�QF1�Ԫ*,U1��bfR���1YU2�#��[Z�[j��V+"
�������I`�*1U+*��b(�QE̳1�+V\�(9fa`�S2�%U�R�UfYbV�3̥����sֲ��j5�^�8;�k��X�˺�&��;^��m���|3�c�3vU6c���g�|;vԽ��xNx[a����tj���ڶ,�rq�ji�:���ݏC��6�1gN���9�ʛx�N��q��/Y}��Ol�m�w뫶U�7e���AY�X�Ԙ�L�9�t���ù���'k��V\]���vwk�����N�.6�49�v�f�_�]��՘cJn�bk\!x���v:GK�ލ:��K����W��r�j�p�mn��W����Ջ{j��Vt�\���n�Is�a�x8����\��� �9�@�M:���!�j�n1Ц�\�wkZr��cXx�kQ�q[�M����v�WF�n�g9��0�cf|�3ѹ/�RZ8�l�7V�X���K�s���\��5�=/T��[��;]���I��4�����b3����;����n{A؊8�Z�<��:���r�u�x=iϧv���n���Ӧ���r7f0��r;nC@���v��^8�H�Z<ݫ��۸��ػv��y���rk�#g�ݗ�2Tm��l]`}����pj�+�8ui]W]�v�����.LBrl�nNK��:�!�Cp���n�����ֱev{c�]�f{B[mʣ�1n��xz�
p���c{은�B�Ƌv��[;�`�8�t�td�0�޳7�t�n3-SM�̣��������ٹ��N��,�gv'iӬ��u�����5N-�<�'!�n��K������4r�:�O�]�-�6��y���;/:&8�*���/]���ծ���[���=�q�r�d���.2�[)*��۰s[v㪮-�� ��-�3�� �۶����j��sWEvCR��nEo⹫���V�[j����sT�(3���L;mt�f�ӻA�t�&]�t��=��t��'S塮�����㕭��VT�󭶙ۗv
 w=k�,)�:�=���K�$�L"vHT���8�;����8�l:���.�.�6�;%���ڍ�\����nn�֖Ǩ�K�u3�<�]�����d8�p�h��y�6��|��t��LN��Cp��Gt���sՙ�pT'V9l�Z��.z�$qS��ֱn��M���,=y��
MW��wu��ݞ�Z�\&-�\�^�ۣFB��cT]�͸���T�֝�<s:ɣ����'nD����#f6�8�s�s���p�$q�j��>�n:��d2a�7Pה����nu�8�16��FsS�}�����	��n�'�yv-$�J}�w�J��0ҩg���b��;=m�H�޲C?bWư2�f��ٝM��\��:�_�@�ܻ`|.����*T�d(��?|O/&)*$�C�,�y�4 U����E�Yy���w>@ ~�m0����:��zzP��j`���,�en�����;��u��` *����
{w�.�����HW{L^W��URDL�_E��/:|�r$ Ov�Ň����Ho|����������	��UD�n�]ߒxХ0�v�@��W3�m�.qS����X�y�[#۬mλ�P�B
]c�(�`���j��ړAE^N�� )��̈���w�ˬ]|�7�yW�y��  ���H-���TD&�M�W��H�����f7v�`:�c_S��88^�ڌ1e�}N��]��x5��\]��
k�{��Ŏ<�F#�x�a�Y�Z���=���&*�wɂ@�_��� N�{3I(��H5@��ɺ������d��y��Nb �n�� >��z��=P���-��7�Ne��"���Ғ ���x�<��R(TD�Ȩpŝ�>�����nU۵�Y��9 J}�٘ U��ᙫ�"ӌ��ӌ��=���H�񵉄b��w�i �N>�m�.��˯�wom�D�<鱄@���f`
���s��WX�Ϯ�VA�D���3fɖ�q�/.���i�����6�����92T$^`�n��"b?,�	N�e
�&7�� �|�"����̾���+v6�B($���d��aW�b0C�l��)~��Ez�@���\������$�A�uP�"M��.uԮ�L���>D��ٹ�)"��!~��ܤ@�{wDN����,=�7k|�j�t�~1�}���]k�g���+�ήv'���Y����Y��#��-�dm�MQ[�����ӀH	��( ���Ժ������3A�'��b��w���| 7�kń@W�;a}<�D�s���7���"�DML���f�`���N��\��w��Z��X^wy���)��� A]=d�x��s=K��	�yp[]���X76�]u�ި��gk�K����G7�n�A�tGg�D0�f�.���A%7���]\�.�[�y���9��w�^B'v�:��n1?*��>nb/z23_�������� {�� ]<ڒ"	��=���^dF��H���"b������>�o� �O?�� Z畚n,�"� 	
ovL��%����"}ٴ�0RMjD��~��]и�� ^�v� ^��I��M��t�D�'m��B��sB�A�o��oo	�P�᷹��R3d��Z#AT��8Zʝ]�����tp�
��K��n�i�ˍ���I��M#�(B�q�m��Nڿi�I�'����0ʵP�^4������]U����w~K��J�������(��cVs�� 驝��8ɽӁ.�����L�D�j`���@��8����ʯ�|�UӭȐ=��Ȉ^��~�u�����f7�  ���G�v �e��C0�1]om߭۔�Ɩ�V���� 
���a;��� �=ɥ1^Ք����`g����ha�g��2#�O{y��l�ףG7����ܼ	�{T!䗣s���hb`��	��Z��LGgE^Qѳ��躨 )���� SϚ�^z���[1�I=�H��ٴ�6����'����0 <������}7���_�W��c@$�{�٘�!O>��.	ҽj�LC=�dD��O)�t��d#5;�u���^��T�7�7;{�д����v��t��H���$�6��g������3^l�7�a���0W��h���\��v�bv�@�o8�ܙ؟�V��]��vֹ�y��peص˦�`��{U�ێ޶.9�pu�_6�t�青��prk =vK����I�7n��u�Y�,f7�;rI�c�6.�cۭ������:�cg��dƓ��s��s������0�6���.;pE�<P�l*tƍ8���9�U-۔͚�v(��+֓�7����[�F�=������[�.��Z1=�|>V������ˈ	��ϼ���UBH�ϻ��h�SϮ�-�",.ĉ}<Ȇ���wi/�ч�Ti�ʓ@*�0�=�Ƿy��� DO���  �Sϛd TZ���������"{Pbn3
������a!�5@���gP���ˍ 	����Sݍ�Q���ET �Sr�c�g��p�m�_HI%��u~�I(��@|���}��_z�b�Ɋ������r�s�|D��4P���p�w�O�z�>�f]w���{�5�@| �{L�ﺛ@)�]������GF7�t�=v����ܠ� ��05n�w\8�;��׋9�r}���~��i�g���`|���� �u�ǫ{}��B�<�=��fb Oo���ݔi��e8�٪�Jr�Ф�\եϲnG�N��|�ڤcϢX��Vxi����s�y�yz��vxM8<�I��sa�}L���Bw4/�F�^]��0txz�<���S��� ���m/$��7�Fj���H>� ��7	Qp̎��� Aw�W�t�z�Mm�lo���{� �mY E�u\C^!OF��¨�+��iqW��4���n�� ]�����wf\'���Zຍ�H���(t��4a��->�4��s��,�ɚE�UN-���v�D]����S�ݙ�t���?>@�In	!�RXZm�YM�]Q����8�\�Ïk�ȇ�gr��I����}��p�����<݂ .� |����A �MQwzڲ���������u%QT*���*�;1`��q���d�y�Y+`��f�%L�M	 �9�٘/���뉨'�j��4�� ���ْ^V���^J7{��$3쾝8���!#հ�<"L�׹�������G��_�H�ŷ�4��^��{���u��k]�r��9Pb��M�9x����>$AL�:$�Iz/{�� �`# ��P�&��V{<�^'
g��"+������@)���τJ
vVd�JY�Ȣ�3��h$�8��`�U2��%�Fvv�`$ Lozݙ�Gz�o�g��က�{{3�������Y.�z	lC��OPL�:�-�,�k��p8ؼs:Z86+�����fs�P!l�v�ԒD��uZ���wy�
YA^�S����l 	/Gn��6hb��l�6Cm5E�%`�{w[��wU5o���0Q��Ր|"�Wb��Mzj��ժ��J �l�ٓ0��	,~�l�ɵ��V��Oz9 ��٘��L�eT������l�/+�O�˹���M�^���y����:a}��Jؘ� X��W]<o��uo[��1C7g�rG�
�nkkyKq
Nʛ��ܛ����E!��CR�3�	;*��'�O��X"���M�@jN+=�U�JA$��k�'*��޹��ӽ������ͥd ��{�R@�p��k\@F�hC	C�]1\\�2<���',p4=���ۂ�T_�w~�< �0�`Ů�̼ۣi �;�4� ]�[��J���#6M��sws1�H&{r�J@�%c�����&粼��ݑ�6w�=�z�` �(�y�@ ���o��|i{�틩�]+�/7x�pb��l�0�m5U��j�%$Aw�M��|m���뻺ܮ��$Y��d�Jg��$�ఢ
���m�mU ��e��LI��7RIi��d�����@�;{1W�.tz�Ĥ=��= �ɂ[m���/]R@$L��<�Gf�B�dE� �[��H"�s�H�Q}�wc�p�|ɞP�}3Q]Sό7�>ߗ�7ĕ/��^��[�'�眊O�Hȼ
6��/t��{��؝2z�[�6�	�(�x�E��aG�:7<�Fh�xxww2.��qݸ6�96{n���g���F8y�$�s�g�
�s��u��wd�^��%1=�Ҥ�<��.�qk��9��ܜ��;�o�{;���Q��sN��t���͓�8'Z㞇z�l�^��yv%��[z���0��l8��}7!�܋�uvy;=���;�g���h%�n㒡:�7B�X�7`oTZ�C�.{b���)��J�m��Y0�`�CM0�D��"7xh<`T ���FG�c��v��v�s��1�تkH�}޸��TS�ҴRFg5�4"'A�!��&R�{y��>�^ګ{{�!�VD +��p�����Ā5sU��J�W���ѹy�P�V0�*h)�nvܜ�H"s��,��<�.3��r���D�I���L�̦m��D��qr]�{#�~�.c@\�᠈Q��vI6��eNus�w8$�IL�:�����@)���ƌ�\��nR��;}n����W[��ڞ�g�XƀH	����>�mYU�9D��E�QUry���ѽ:����m��n���u��\����t! a�J�ΏG �Dm���u�P�>��<XD I��Q�WN���Y<ܐ$��oZ���"�2�pё��Ұ�rǳn,��F��<�%��Ӷx��{�����H�:���fj�[�ooR������}�i�ssqw%��7O���Lr!;˿9	�ﻳ"0Lwy� @�s3�8PN`�Ef�HZ"tbJ`�&����� 	��]C�X:����o9�(��H(=�L�ْ0���5!��1��E_�?�nv<� &��D0w���'�R�Fz&ƄΤ��w�v[�������i��0�[��y<��?^^X]<�����@Lwz��@��O2t��O���z}Z���4�E1��e�&w8�6y������<�Q"(sؼ�>��l.����L��)�=��@�Lv��V  .���������|߀ ���o��Fz	d��f�*ˎ�P���L�z�9��@&��D?�.�y�$�,1z팞����В/F��h˙T8��y~�� �������t�U�[��h^���Ş��Z���`�r=�{��O�T7{X�h��G�O5�:�9���f�Q�C}ڪ�q!���{�m���:w㽳���4��A������b緈��#P�)�[@[��@�qf���s��'�:e��A���`�s}��v�9���<���j�}<�Y��������R��!��
v���c@d���]�g�Q��U�����Z�R�@��i����B��]W�ݭ����֞�����e����
��O�d����3p��R��e�2/A"͎��=w]\���ON�^�a��/k�V0љ�Iu�#Sb����F�RAu.F��T�ځ�(�����s��{g��m�x���{Yf
�x������e�bӋT��ܦz(Z��{kݟ�y?u����҇��4���v���	zze���,م,\F��D�=�I�n%
��8V�q�77!�N��`֗g�{����s�`�F���z$D��{�n���O��n�B==;|d�q���w������r_u��Gc�?p��I3I��&���k��`k���	�|�G�b�<_�{/�y@�;K%���Fiw�bx�Ox��Na�Ν��K8��^���qY�ݦ"n�a�`UΥ�V���kтA��nH��a�|�H!���Y�r�rǘ���LΤZ��{sI��R�l�ȑ�*%[10c�Fo��.y����Ϫ�_|��fz����BR�N���`��{�.�{���^w�'r�j�܂�zx Δ�Z�e����1�ՍJ�Ƀ�[�e(���̘mJ"c�Q[JV�˘�\�E��V�[m�8XUE����(��)kFR�WD�m�qUPX�ԮPiEf%,X�q�YUᖙb�&6V��fXV[s0µ���9����U\��%�nfe�̫*�1ZcT�Yl�*�̪�����*�VZZ����6�b%��j��*"�EX�LƂ���Ѡ�),�6�Ijc�0�[ee��U-�U-if%1Ī�m)Q�kRmKm����̹j�a\�\n\f�p�+j��Jy�y�� ���c��ݽ��4L��ndS-��e+ZTs�v�	��e}�����2�Z�1QƆ%�Qh�m�e����˘��q��eD1�R��*)Y[liU����mLh��l��E�J�2��R��3-Tr�ڱ�DƖ�m���Z("W2����%Uq��m+�0����P�Z���Z��$�r�
֪(����nXX�-k�V��k����Z�[i`��s��k*�R�)�V(&61Ź�\�w�y�|��`�d�i$�z:�а�<1� �\��ۘ��=1�:F�L{�ڰ� ����� �7�2��!�_��c%����f��ۣ9<�
a�1O����9>�o<��$�Н8R|޺�h��ͩ A9���z�gD�ߥ��������ߟ\"�&݊	UQb���a)��;ǲ�=����
`�����e�i���&kX�]���>Novf|j�����A�ʡ(���r2�B@GV(��q#����@ۚ7w�i��J>�Q���� {Zƀ�	����	+p5��c8����U��ў�C�m�[@����'�;�� 5E���mT+�3������mIA9���I�	�D2��TiY�ʝ'2Y�M\':���{s�?� �����ݕ<��p!K���w��h=4����	9Fh��]��B~W�6C�'�S�@���<:�Y�`�G��*j��:辽RV�^ٸq��발���H)�����*fa�4���1`| Lozڱo��E�����c9�٘����j�v�)n��Uw��|�����o�nJ�������Y�z� ��.�M���f�e���������C�����A����@﷛�@�v]0DϜ�7ꂪL8Sq�[��h'�����9	�n4��v�J'�C6�4=?{�n:�ݽ���&;�� ���N�ce9��5Q<�D��74������+�;1` �L{��"�oz�="������͌�I%���&�H�޹�JB���_���l�%X�����_B��F> =W�y�A:v\��@"��uU���M2��c@����b�P!�����tq��� �/Om̅��3-=��""1�nH �;�Tk����]v/_A^��/sn5\��/^;=���n�ܶ�|�y��D��,5�<6վ>8�q���ջ�E
����W01�"!�(e�Ra��F��\:9�'��<l�v���l%g���:'����S���������f�qn�4�n�����3�jۍsT��7"���i�}��q�x�x�&�;�دe9<n�m�kq��3�K���%�t�t�8;؇��<m��p`�OY�r�gO;�N��)L��m�]pwܯlm5���'\�k�2<�cK�-�����^.Ǳͻ'W]��j�=v�qvMnw��[l۳��~��S�T)T�v9��`�N[�� *��A������`��7�'�Y3#�}��m,)�p�>&���g0�ѡ]��_������==u�I9]�^h�*7{�{\���;��꫉= ��U54T�8{~� �3�N������͛/%�x 	㱺 ���n�M�2��T�!���}}�'��8!�0N���m���
���h��o�%����]A;��OU�^��_�!�6٪~3��|��y�z�f{øj�r|���- *��tDA=����|�����>=+�Wn��mn�
ڃd�nvٍg��k��z���݈ۖl�m}���~���L�F�l^e��gkN��)�of`=�ʷ�7ue��==4��E�̚,R���!ApDQ�+�λ��J64��=t5\-�M�;��ɘQ�5��ך݉�f�.2q�V���ݖƲ��z%��m�aS����_Eݏu�_;���ǳlqn2x��M���I'��B %;���@ �،꨸gD+&�m߬>����(���*hC��0�4� |��V-L�V�/�Y5l�	/'+��4PI�޻����,�1�[&;5��d �y���W���tv\�	��7� Tocؚe� sk=��[mPM�eI.�
��O>��G�-�#~}3�y<m zw�D��uU��,�\ԭ�LuA�n���^��c�2�7�J݌�뛱��P��'��5�wQ�Ĺ$���ȍ����̐�l��*�~iЀ	���AF�:h<��v�ma&TL�Z%���A4��vo]�HF�&���KM�gD�D��f�.�K��g��: }�������숍ʉ�$�7�Z{V��B��1F���c�Gn[��;�u�R̭�_�&G_�ie�������W^�}��l��׀��f������ .b��eP���y��7훦@��徯t����;�Q{�Ui�gz� �ce���4E��`��,�{��f��	��<�  ���u�	guF���	�.q8�M��ۻIxn�F �`��i�>(~��I�@zo�R~+��H	:����>*;q��� U��C�n	�.��b;��� ?!���a���z���H�:��N�S�^[q'WW'����ʓ�}5S2>En{٘  �����1�QIf�,=�5��}�3��$�I�����$E��$@��4L��BA����U�}�=���ۗQ$\�馉"c�7�:�][e�ܰ��M��'�j��=r�y"\��גA!Q������d�k9��$J	�ۦa�Vw[J�x�r�ML!UH��y�j��j�ϛ�X\�2XKOM	D� ��|�S������b��ѯ5축�Z�ˇ7'e���xBpo-��9��>�����e�U�6������J�1������K��� gP�3���3�@JF�-���hZü� /�s��}�����B��/� ���4�f�Q ����9��*څ��T�� T��kW@���IǇ���rI��n�����>M�%������ܝC.-��r�w�BR�I'*�`�IE���9q9�%YQ�i�d�^NWm@�-�,I% �6�0-��Τ,~ƞ�6MF��I9]��Q}�wa$���ʎ�/4s��Q׹ޔ�W�H����h��[�S^Iy(�ޫ��@��9�+�F^k��gy� Iz/��ɿф�,�SP�Q���c��ͻ���Fg� �Ӗ0��˰�I&w���D��#&l�a$���Xe0���*���]�A"Y��q;=u<�}����k� };��v�+ɝ�zZBs�o2��c�g~�,�?f��{�$�� �}t�ܦ^�{nE���}�,.A�0��th�a�hсL���e�(��TҐR�?���r)�+���g%tֳ�;s�n�x��7<�֎�<ܪ���b�1b|ʳΟ����ҽ]��w<�ۆ���	sƐu6;g]��;A!l�����J'�9�ƹ.���S�n޶.���;����E�Ga�A�]؞�q�y̝��;��sN��Dq�m�0�g���k��u�q����XVgy�n�!� ����&�66�ng\7��fq�R��v��G��/]l�N�1�k�;qۣ���&����Oa,|���ﺴ�:����g��D0����[=�-����F��I�"U�~���ؠF��M2e��3}��O�*��O,��כ���s��0�6�󘈅"Ϩ|u%���J�ĥ�$�&�FL.~���H� ���iP =,�ǒ��d�� ���3�6���A}�q1�UB!�m�U�.:c2X��!�I%nk�ŀDs�r� S��<��:�;��:!'����_���8)���0�]�A�RN�6�Q#�fe�f@pҝ�� z��j���}=d)���w.��[���\Y����Y�$�<�nWr������g<����$��n��0t`Ân��Y���� �:���@�@S��D{��i�t���.���H�ɠ�:�al��I���#NY����a�T�����o4�5�t�
+����Xu��dEµ�m8���FB5p�������Z<�n.Õ��V_տu�ٯ|�eޗ�뷗{���` �w�X�}=H�J���7%mp=m�ø:1d�⪈������5��)���Ȃ �������x������ @�y��[|JXRK@�6�;�u����@��L�C�P| ���A����6������S8IZ�f��� �!���J�㪡�����]3e��o�K�nLMy:�ʡ��no]�E՝�Xs�=q  ��hC-���"<\2�a�n�A��q�u���i��^i�h��>��O"�5�Ւ�]�4JI���B�D���v� v��o��E��U������'�S2Yho���j����JuD�w1�S��"@)�of`~�'11���5s�旎�[.!B��ATRW{>nD	��n3�A;��`�����E
�ݬ8����Fܘ�Vݫ��9�/(B�z������}��p�%{CZlנ�5���^��$��uq�|�$�W��m�O�c�B4�m�������{z� w��Q�I&�V}A%>���� �w��������p���CW]�L��G�U3#h���ŀ��=gz�ea�*ѳ�a޹	 #s���D�-k���t#^��4��g��[���;�X���C�s�[����g��q^�'%�0�%vX������8L��L@|���a ڞ��[��̰5uT)$"���,�M2
j!�Sq���7@;Nv���γ�ߝ ����0h�6���ǪW�:(��̅��羠KKz$���!
�F37;s=i��&�I �ڋ���:��$�y�vI'c��a/y�l�1�mQA�w���f;=՜g� ��s�"����"�w8�N�m��)�s�<�g�V=e�<�s��s}^��MƲQi/��������ɲ�G��e�xN�\�^c"�6m�A��{{����c�$g�Q4��*�t���H��@����v!nR@9���I��є���t����w��"M-{�)�b!���װ�v��wۓvsHr�nZ��J�b�9�^�~��*bT�!S2>)���� ����� 3�堉q�yO����q�nT��&��1�j�U��b��#w=��.��7�/������Id�(��1�����/���A5Ji�����v  �v�B��5�f����z�> b���A�郅�\!b!�J�+�ζ��qm»�قh".7�� Nw\�?�J/w��eʤj�9����XX]m2.}�b�3"��>H3���w<�����6K��Q�r���3v�������-#e5�nclA�=)�ét����ٍn/ʴQ�7bX�u߯�"j��
�v��z����`��j�.��Y�h��ӕ�_L -Z������F�]� ͷp�� vq���+F�3��i�sQ��2Ɯ��=��w��ᢑ�sj��W"�ܝٖ{Fyzo��x�N�-\����Nh%�h�V�̊�̍U��lm2&n	7�ˀu(ֵ���1����w˗����h�\m��v���g���_)}}²���Dz{���\�k�*��Y�g���^RY��O#�ev�d8�{��w��AW�{����t��H:����^y�y��T>[r���z�$Y�#=x/[���q���ފ�Cpص9 ��6�Ji�A����1�}�'����q+�w�_��k����\yg�h�%�mk�߻�L�pM�似�)Į��T��3�ݽ�w�M5a>��g"@�/^���>�y+L�!�<M}|�P:�u�p홼棇�/J���ۡq]��R���o����t�J��f���𦅼U��-�>*������O~;�[̺�刼�F�TV4���6�lJ��\/y�ἓ����&�z��v�(�yh}�{`�%w�Η�K�/��s��C���;$ԯzg{�G�w�b��c$���`����f��\]��{�FRS'W=��zaɚ �rrz���ȇ{IƧr`����������Ν�����UĻu/f���unobba���7�1��[a�3nE֍����w�[Ľ̿^�iA � �Q >�K,B���V��
`�\�v�˼g"��p���Cl���*�ZZ�2�T�
�YS-�T��E�l�k�`"��KJ*�U2�bbjcX(�[a�R�Z&4U+E�W1Ɋ*ܳ���"�j�q�Ħ�Dq�l�k*�ڕ�Q��0�EX֨�(�r�Z��"�m+QiZ��T(����b�2�)mDA��j(�`�T��iYR��S.ab�6Ҋb��YUb��X,�JZZJ�R�Ƣ�J��(�*��EKj�����l�DTU�fPU\�*�i-R�\ʰb5)j�s*1kL�����2��S-�V��(��J"T(�E��AQQ-��aik̆eG2Ԩ��kDYq,T2�jb2�UUeG3 ��9�&%R��-m[X��\�Z�1̣��#LlUTƎV��qG)R2���U�bX�cE��[B�\��Go[�%ۮ����׵#����uoC���v����K�:�m�Z��OA�L�-����[9��GJO��rrݑ1�۳�ζ1q�Q�&-�u�d{%���v��� D����>+��e��#:�Wj�!Í��f$2j��lr������q��(+��Y�Il�m{�zӚVr�v�ތ�\��"2v|�w��#�v뱦����ku����-�c��/��IW���=Qtq�`�n�]�9'����^р��v[e{q�ɡ�6{gv�;Cέǻ2"Gv^�n"�lȮO>�����g��3v2������u�c�i�|��:��ur��(�)\a�.y�v�mݳ�gEz3��of��9s��G\d��Z2r��as�pkh�}Gm��p�\n��9y�rX��Ѵ띹M[��r5�u��1�cxm�-�Fm�厒N�����G��d�+�vOn�5nhn��Qc�슼{=ٶ��1�"�4�mݝo"�Í��;�u�[�2��k��
9^K]3t�ҹH������!�l�ׄ1>t��=��g�i�4n#OM��gF����A;<���{Q)ː���/n;�ݻg!�)dhr������e;��ѹ�ۣ�.�dW���vq؇�R��,��=��yu:�ױZ.�=E+]��r�=��E�=w]\����8�5�8�α�	�0��x�t��7k&��2��v.P���q���Ĵy#�i�{]���K��/=�h�tki��8��0U�ٳ�6��m����^�K�D���;��ˆv�'��\ HYA��q�v-m�3��뭲N'r��[\=�z�1�� .�;�)x�-q�U��z!�+vxv�ۨl���]�'s������\��8ջ޻����Ju�Gbf�s�7����^�vQ��ٮ�<gm�=��<��Zy��'Q���a�4sNdS'9*�)	����N�G��6���ݷBm�\/eե�3ڞ6i��쳎��!:qIv��M[�zd��[[c�v�{����E�ۍ<�#��r��5���d�J�b⋵Ѹ�7�;oq��x��=v�[:��z7:5�=���Yn:䔁t˞S��%���۵ս�5��܌V��q�Aی�J���:�z�yN<mf�͎]MIۗ>{nûu������\��Y��h��gv�n\9��r�:c���v.;2b��H'2��������,��@�ǲ�����]��W��o���&-������t$���$�8W����d��6� S;��+��&TĩUL��O�٘9W�{�<b�5C��|� �>�-��������-f^>�F[7��`؂�bl�3��c A�N��q�CZ{���m@zc��� �):Y�M䗢�z��H0�p��0�C�JM�Vob蕎�8�O%���  ����� ��3��VϡRe�^&��:-�ٯ4��P��-��¥J���$��;�^��gvp�ޘ*�@y=�X9�٘ؾ��bu\�n�31�	�#�l�p�P��N�/=(��z3��u�4W7v.�J"�:������ё��=<��ӡ ����I�A-�}�8U;����O&�D��y.�a$C.
��sK�����S�*v����؇�Ywq�(�-^���B�d:��2�R�2^fѵh�&a��pz���s������w��Fڈ�}��5���:	 ��ofb@ ��t`B_��A�V]Bw�YRVO�� � �O�-��������I'���4�Z�S�{rf�&�ZAO�{2"�GZ�59�LC�Cm�&qWM1yZHS�7�y�@T��4�wJus��ܢ�Y�WU~I�	��}*j&�M8�y�@�AL�i���#��6wYpRNt��� �y�t��?R)��аp߈�ww���zR�'�(Mm�j�d۱ͻ%�]���m�N�l��֯݌ݸ���;D"�l��p�p]��v-�]F��� N{��}�$��:o��ۙ�@$z��j�6��THL���9a޹a�Q>�(^�}s�v�� >z�|�� �w7�|��O{ўY�L"�s3<�h�0��!�Ci����mP 
fst ��D�B.M�
��3�&C��v���Y�V$�zm����ҝN������ܠ�>�U{vBy�xvB4j��� > �7ͪ �����LL��R� ����S��ګ|��*+���
��o�@S�k� )��̋��|��^>�YsA�9�LC�Cm����
d�'�����˝��~����  ,�k�(��$�n4T-C:�q��4��tf� �.`�s.�m�;������/]�ld��N��A0�8��ٕBQ$�v��H"��ݙ��~
����Z|Lz��  �{�a��Ŝ��
��*(r�{ۙ�����t{���~�@|9�r� ��vf HSQ鎋��3�(;:i8;���I�bha�i�ڡ"	�o<� n5��G7�T҂�kP	 �f��COv�f �Sq$z!M�9<]d���S����$���7B�+�(�$�:_Tȝc�ne��¶�f�<g�ѽ�u�=+�;�\z[��h,=�6��qn��%���0f�ʾG^�*Kfp�@��>�PX�Ő5E�$��bΪjY�0�� $ۈSI���K ��W;vC~�;�up��c����}�٘ خm�=�nm������mc��Y���c�1A��2�j���ґ�	����+s��������c\�[��L�u �o�n1 �ZW7O�p� dګ[�:��	(����m�A�a��$�}r�/�=�Rd��ٕ�:c �>��f  6+�j�}���:_��wcz�z��b~RPR*�"��ggn8� tV�X  �{�>�^[��/.tS�ݙ� >:+�j�!�oci$�"��� 3o�	�X���w� ���  >⵺ ��Z�oѦ��q�IOne݄��r`#~��T�h�y����/9�����H��W�1s�o;3>��m�d	;;�2ܫ=�O�z�6�d˪L�'s�t냕������&��2ٸ��ul�v�n�[�+8�j6�3�7�@��T.o4'��������h�#˞uq�<��G7�.�*�Fe�;=(8�$Q�=���ɳ��;��qZǞ�"�>�[̛�"��3͢�����"�օ��>m����m����=�+n��v�l�vA����̸����<n۹�����	m�<˧u��>kt��ɻ{[�w=m>Gnq��&����5�m����=��q�a�z��%VK�aase��8�����f��Dm�x-r3��5^���W�^4���>���������EL8����  �V�X �	��9hU����S�ݙ� �[�P���Щ	���������J��W'��:���~�� ��� C���N���wn&��6k�ڂ3:%�ۜ�I5+���NXt2�u��r�U�@#b�� gs�kŉꚒ)QD�Z3{ۂ�]������ /���T"��y�CH'7���ւ380��H,�=TF�b0AQ����h똈�=��\��}ݾ��sz� vn�D	�w7�^L�R߸��S��b�$\BNfpP�=��ɹ�Q�h��x�0Q�g�Fn���{��=�'6���3<�D;3�N��@|�7�2!�|�T)�4�1�Q�|����st:�ؒaJ�H*��������'�=�t@9���Qj��H8��KZ\͌����ٻ�c0TS��ҙ�۞
e���|��}�U�;�;����y��Ε�kniz��3�1� ��9`��7�%�8f:7�{2�kP��^��&-DР�����9�B��<��"t�*^5ОMA8�U+2��j/���$_&1�fth&�)l�'��W��=7Q Ov�x�]���{�~�^�MTw���tŉꚒ)QD�ZFvv�@ ���g�>�=>�U��	S��- �sw�ϒ^I��S=����e10`�a�#D۬Y�鋶,n��=��@n��Z����\%��6y*	U0�g�>=����  8��꯽.'�m���|�!(�޻�$��r`Y�!� ������j��ݪ��ӴO���N���vY6�\_e2i(UK��;���j� ��8e��	�w]�D�ƻ&	5�Vjr.������m�r�R�Z��{�'�乺��Ц�����q�Oj�w�k�����{IA�6�>�`�G�*|� 	�w7� u�����i	�������7��n���F	��@ �����D ���� C���Uor�����$�V�V��g��Q5*i���;�a���ө7�{}Q���1 6��t@������1�Y�0�ba��h�%ؕͼ��;+�-֎�+V�ۓ�t6�qn���N����h��,¸7yy]�D��5�4�I$'s��-sg��*/�g���0:��[�Q2�U��"�ٮ�v����*�t�__��"ҷΟ� ��o�"#ӯ�Tʏt���ʮ'!Lʨ%ET�S5�0>g��B����Օ3���B GEw���)���@��H�%K�����o�S��Ϙ��O����z݀Ns\� Jo���C�D�i�ÞN"���7��@��r������vE��=:�C�F�`Dm��b��Ԏםw� <���	�v��-�,᭪0҂4�81��6uʸ�$��hNq���$�e�!�~3Zt >	��nY��l'Hfc��L�7�"	�������;�0X��� DEy���D8(�K�p�[j�]�Q��k�i��=u�h�����w���9�*k"{2�� 3u��@|�wf`f�^���{ݻ��h[���d �fsj�x�f��� ��9#7;s H~S
ծ���*s�r� �w]�I$]�.�󺠎�>YO,
C�򈊙RM@)���vy� Nv�İ>�7w9]`�f�� ���Novf/��M��"eT��jb��<�*�"V�����r ;w- �'w�3 �!mw���lS1uӞ���(�7Au���
�T�7�o��>�� �&�\�Եτl��%�v6�	�$Ov�f|�mw���}�O�\���J]!��{_齫{
Oy
}���Z���l7�'}��z+���Rr��,j1'�d��v#��L�N���������qs{;�\�G
���[i�0iyq����'h��v(H��{���v��=�ȝM��;�7Ks�w������Y�E�.�%�g��	oZ�)D���vC��֢N/c��{(<�-ɺ�m���ӺC��_Z�qǊ���h�[sk���s�)waö���[��l�ܜ�{:�		��{mh�c��pu�+��j��!�z���5ź���Z���6-�b��/nj,���)q�\`�DB�%VZ���$�0ࣜ�3�����<�H mw���2�VVU�x$S9��"	���π��蒻aSX����$$�xN^�nۣ� �s�٘ |-��&@�]KO:�����2&9]g������Ey__m�&���,ג^	^.&�qV�Vn�O�"}��� lW�I����"�'S	���6�M��ݤ U���\V� ��+��3m�y��}�����rP\D�<f�sҗ�%�Θ��0�7�f���)��f$6+��d �uSR<�M�6B���܃2��`�f����9����6��j�r�c�-��]+ؼ~~�`DA��)�w�30�N������v�a��U��U�"O�,��f]MO�4��/��Ӡ;2N��EA��>,��>P�;�d\��9Ms�'���a%�a83G6&K�2�ۿx~����7�{�$�]�x�` Z^�i$��U�&��S�rK'Z����W��!�q=t[�4�$��vܿ��:�9��~:����o�#ZΪh��QK���,FM�lCC���7�ێ���EM�e_��݈���T�����ٞW�J���f� �ѷ0�r�y�(��D��1�˟$�9���վ�w�=Ӽ�� EY�n��'7�3VU7v�TzA8ؚ�-��qI�9�C&���`�v�����7⁆�p�04���ۄ��M�ʯ0� �=�,"9�٘�w�8�b��k��ی�	zo�g]>(�-�@qk�k��Ť��<g4k���d-om�A*��9�h	����>+|}�Q�N�s�B��n!�
!��C�ιh"'w�� ����Xܷ�?���^ؔw��9��L�4�Nl
z��Z�>�=Ӯ[�sw�WE� �,.�sss��	Xō(�����h�40ŗ����|��m�
�'ۂ �f�y��ѨS�2�`��3����v+c����Z�� �d˞���UΝ�C�0gg�i�Vo.�Ϟ�f������k�yV��R�紿\�;eQ|"Fj�.����U"yW!�/�{�М}J�����;�f�ar����;ϕt\la��[�o����%������szA�ǘ�)�;Z�"���Ʊ���5/�ɫ�!�)㹹����u�iObH��~�u�!�����S��kc=[Q
�׎�[{����{�����(T]SW�+3wP#����ocȯ����N=Mo^3M��f���o�Kj=���<��e����f��ݓa3�����'D~[�?)�*������mŶ��OM��	Jr���;g0�ҞwD}��3}��a[{��NF��SwE.�r�g���a�F�zh�q��,�^�}�C���)���h[�&K���g���;`6)��jR��`�^���[2��+[⏗g��ZX��0�guK5�X��j�,�.f�E�s'6��Z��n��}ڛe�.�*���N0z1�E���R@�y�{�{^�׿��5h[�c���9���%4�On���B�ܒ��9�fge�Qu�/t�{��������(5t���}�]�<���n���}Ύҭ��ܢ����w�~�;��R�mF�l�j"(�U���
���81��*��1¢���*�A�b����.[�aL�#�LAZ����-DDDjV�*���FQ*5��L�pD�-��[Q�A�PQ��QDq����)j�B�̦��Qr���֫mj�-�m��[h�,�T�b
-)h�-�f�lS1h�5�VԸ�dV���(�m�+kR4���b�Ze�mҮ6ڎQ�Ҷ��j�PeUDBҴ˂h[����8e\m�m-�,�fQ�0�9eˆQ�YiF��X��ib,UF�2�e(��UJ�[h����%Aƀ�Y3
�D�X�+Qr�-V1`���Z5�kE�e�ܡ�,�\̙ZV���܀��1�_ ��x�wg�k-�.`�(��Ƹ)kE[X��b[���"�m�1����",�fbb�b�T����[PT�ffZ)���L����W±kQ��l�X�S+�~"5�w=� |U���s{��$6NQ�mB.�Һ]�B����qxTm� 	�<�	 �Jsw�0 J5vP�X�E�W��\��f��'�y}U�F"��lC!�A��g�p	r˘ȶ�L�勰�5��T ��;����u�+.:b�̹"�����Am��5�
��C��'me���ݨ,WWح��uh/��{��[�
H<�v�2���U���$�Hc�H1@��ئhN;�Isz�}�!�R��Bm�q%�A1Y;#2�:ì��� �f�W���]s�J�+��.��3#���,P�"������'ăp�ԑ�i|���«6�$���^�����ȁP�"h�d���F<\`����뫚GDe�'�'{�Ʒ��\laS���ܠ�)��7�鷔n+΅�ǯe`��y���
[b�SS�4��dtz����3.����8 ��9�s}��Ċ���$oH�J�(����O�V �~��G��⢅@(����;�D	�OwU�.��ˈ�x#SfJ!��0������6��-��;�4�qE�{��^-�p�lo���������!#�ܭʣ텗"��}�U�Q4���m��� ���0wA̠In (i ꁫ�ɯ�'�i��ɨ���I�[jI�>���D�j�3fh�ku���`�`QJPa�Ӂ�,A$���D��h+���uOp�|V,��K}�4H����(��0�UL����l�Q�o�����@$x�7W�@��}�[}չ'�]C(�Fʮ�7X�*p�"$g�篨Q ��{�D�����\<��BI��P �{�U�.�O(j�%<�=[JDN[�:r�=6�/6�#E�h��N��wzY�[��ahK%ˤd�ߠf�2�U^�� �]�Yק�_�pa�Q�NZmv�y[9� ����=�dQ������-��<p#e89�ۅq�t��C�\X�p+�ö�5�ţe�� e-��Ϯ���`��:���g��t[�Z��^ յ7�l�9�[t����n\��Cv�Ƽ��sq�q8��jFq��{y�ۗŷ��cl���P���n#u���R��b��m��\�m2	��s�K��'�Q�Y�C\��H�sou�3����mƸ��<��[�sl�~ﰔw���A��Գ&$�v�J�!��Y�R����9��DHn��V"��lC!D$d
��VTgV(�|��I��z��uP'ǸYk^W��E�Q��CqCI"j���G�*�zhI�˳����^3��mP$�}�B�I�E!������8���+]�$��e
 ��w�� �b�WM�+a�#'��QkT$I��" '����B�9ӑ#�5;��,}�mDAW��^ٰ�-1��[ �dGTe�yu���\\q��i�Mٺ��DPΝ�">3,�Ͼ�YL�!�!�N�P�H+�ޑ@�Lw;"�͆of�Y��W{{ו��ު�3��g���A��n�2@G���h����]������чw���<	�.\�Η����tzY����d�m���8.�:�	5y��.��*�\^w�J����r�a��
�]��M̀N��YlC��Dg��}T	$�fI�u՛N���8I*�z�	�]�R��AɶP%�a�����YUp��uS���ؑg;3�����>��wMT��(]F4	]}�(^�f,��2"��O�ڌ�"	�Ϊ��4�ͰM7�TO�_E$���"��]�R������A�6���8cp�3ꗰ��d.ںP}��ݫO]]>��o��0`$��;����b�A-�uQ��ޅ��60�˪ ����;X�SA2�@�E���K%����)����H ��j} ���Aۂ�Ԩ��Sy�H�d%�.p�n��v9 �Ku�T�孨�H��f�*�$��٬r�N�ۥ�W��F�E�Y��6�GW��o��N�QN�=���H���,߸R2�!����VNY�'5��j�G���>$��~�O�}�TN"�Zl6Km�(Ϫw�����50�v�ĝ��2O��y�TA]��QB�:��;}du�\��zm�	hi �]�UWf��,]i��/>]O�����U�B��<�sH��L�����w��q�۱��$76S���Has�%q�ε"`��ݛ�9�����߃�p���8����:E N�wU:w�Yk��r����za E���8�W]U�|uYt��J��f9� �D>���;��vۊ���EM�ƻ'�Z[H�	�l��d���$���>�a��I��*����4q>&^UN�wU�|.���p�n��[ޘ�1��}]5V/6���ު�$��L�z�wU��_L���=�z27���l�8�Y<Z���֛�=a�Ҭӆ�پ�_�x\s�����w*-��U�R��a�m
ț�Շ�:�D��jh�ȼ�M�a6Yq�vP�H_S����v�o'���Vwu w��1���~�?]e�	#�l���p����W"�oW�Cň�:��L$�
*x���Z�H=�k�2kĀWf��$���� ȶ4U�X$�v���m� B��^܂�Y
 
m8����wỎ��(�@+;zhI[��jc`�D�,�ΝЌҒ�p�	�T��P�^�A
�z��w@J�2�+���@$�NIXSJ%�p`B2�_oL�rʝ:�/WT��$�|�j}>$7��P�<��q:��H�}t6:�&Km���"�r�+��\2r���	nS�A-�uQ�\"F�l���8��B!���/b/{��9��d���e=x��4����r���3��ʹ�w6�յj�Q~M·�{&��Y�'����M��3�nVN˽qnv�1�lP���/oD�X�!�ֺ%7=oc{O���j9㔻+d=��m��^WWF	6�[�<��x�Ի@I�p�o"���;/G0"��PD���uѬu{u7�s����r��kChx�]>�x�Mv{n^U+�����.��ћsZ�Bƙ���`�׮nM�p�K���[�m���a�U`�/O<t�d�p�d1v����<��d��2��e���;r9d�=x��n�;��m�\AF�e��
� �"wUB�ч�':b�Nx��9�>��ő	�����H��ʔ��\�q���ٲ	[�Ē=�@���,�]��tn�ނ�-�	5N$��~���������X>7�N6��AY��=�2"�����8Bq5=u�u&2�C�������@&fP�	s��>;y7�q�����)�	�80!.���D���5�j��)�t���H$zv�gt�5�Rxw%���"#��L�"��A,��KŲ\MG��A�ǅ�l�Ѫ�7'��������zꎬ�v��|O�:ݚ$��4{\(&9�(�Y�L��> �D<Ϊ�}��CE�Xi6o�t���nV,��JKl.k&���fZ2�v
���U2���~x�Ħ�B�^��`
Խ����ք[��lq{<d⯼���'o­��p��1�B�o�	�U	{z��4�TTVDS��ޒ/��V��&R���d�$��5�|H5��q�s�$�H�}�D����B�dJ�ӈtLڊ���~|�<�#[�q#7y�+z_�+�k=�Q� ��Ρ^��$-����/��Q%gK��OE��,�)'ӎz��H�z�;��q�x�)⨹.~��P��2V&Y)�L`A�7۫��w^��v�����u�"vbǳ�|���h�p�(��ھ�B��$�|��}�����:���9�D��w�P��0b,��mꁺ�bA���Ը�1��n.{�Q �{�TI �/�]n'�:z1���4�3��Q�����%ω���r�Z+cf�l�m�w�X�W#�軽�����{�ȿ�r��\c�Đ�;�Hv�ɋ�Ȼ��ry\�7)>&���Pv]4a���$.��AzX��vU�L��Q��ˉP�S�xH/^t� ��2�7��J��.�\
�ښ=����Ai'
"K�$[���75=rH���H$��r>-�tёH�ݶD�tG�����pZ�c�zn�N�=��t�)A�); �N��^���?���!�H@N+�����
Ζ'Ē��U+5�vD��7�YU�I+�\�6�:��JmB�ύ�_W���&��9�.7�o���|�fD�o���'"kk�y��u�/�ۅ� 0�A����$�[��I�1�B�͸�ިȫ���.H �7��@�	�2�h6`#]=r�U�qN�0����'Ă��MB�ޫ�v��W7*o\m�ޘf=�3k669��.��mד��i��wڻ�n'�o���ǳ~�'�4{O!���w��;Ȃd:O�����>Nz'��� e2�sF��&�%goH���I�2�#&�D�Ku�T	�ݽT�"/����/����o�'�%�	9r���ۙ.|N�!���a���Q�[���c������|��^~|�|I�l�%ooU����V"Q��~��EVg7���`���I-����d��g�&�jt7�$�w�B���$�j+�!;�K������p�$x��� ��{�P$�����#U�=��Cy�TO�]��*3��Q`(6�n��v7�19grj3�5uU
$�|����%wSv�UtH��"f{��>��[)D4�!�"EN�U H��ƈ��ŵ��pW��Hsv�y�m�	!I��B���	!I��	!I`IO��$ I?�	!I�xB���IO�$ I?�H@��	!I��IO`IKH@�r$ I?�	!I��IO�H@��B����$���$ I;H@���d�Mg�\��?f�A@��̟\���                }                  ���  �Gf�P
��V�5��%a��7��(�:�@v�];1�`Y�����6��En��5@����ZeM�{�                                              
�7 ����yt��@O,rh
�  	5 �k����0=�\�:;g  	 ��Ѡ$�	>   ��ٸà8� 4 ��`4��#@���� h�����r�� ^�� (jA�|    �      P ��#�m r2�}��=�7� � ���{�^@wX]=}� ��� ` �ǔ�$.f�'�JlV�n    O�gAA+ϸ��JM�]� OJ*������y�z{>�E�Р0=� �}�� )@�77��AAW�җm��Px��)JO��ҽ4����ej��Δֻ�  >        ��ZҮw��P���W=ϧ��aҕ�}�z�|��*��p <�3�j)́�T�u��څ}� {�T�m{R���'��� �:w� �|ڕ^�;u�L� ::����떇��73EQ� t��#��ODA����y�Q'� z��    P      �>�y��E8�]
rtWRq�
;� �(�-w�q>ç�}|@�k����U(d���R�Z}�ݰ�E^��H��  �6%_*s�E/�� ;��W�@��X�\��m��k����]��GNv�ѹ�Uu��R*u�[m��kJ  �        �}
�k��q5�E9��l�b��� ]��9��j�ا��6�A6sb��>�z���v`��]d|��_   ��^�r �;�� v r>�����@;W à=�x��z���r| ��4�* �S�0�)P   �=�3U*I�@ ت��R�  T��*R�  $�D�J�  b_��?�?ؗ����߾ }��L����'�˒���$��3?�HH@�j ̐��$��!!I� �$�  >�}��/��x���������-��G��"���ɫ&�O(2m��e��3n���7"�ܐ�=���f��=7�]7��=���i����U5X�cF��c���C��h���mv-����njᕏ����:�Ѻf���7΢0���i�7��@��Bc�8l�Սs�sWX@�]��
8oR�,Xw���6�7��[��͖j�*4�L����S�F�0�ɩ"�Y��j֒���.��#�]p��av�|�ܓ�z�����l	5�n��$�w0ױ*��õ���2T�d�bS������w�
��<{5��B{��`.Wu���r-s���^݈���Y��We]٣������r=3�#tb���:���j*���/�w�,úpm܍\6J��X������������ݾJ�5�(J9�I�rM�s%+GM��v�6��P��0oeyOiX�|\E��H
���Cj|`�ڃ��-���Z�YgaN�wz�f��rټ&��i;)�4��&�\�$[p�������ي��.���8%���M�کH6�	���;��U!`�Үm�Y�m&�1�崶��[��֞� ��,�D�N����w�����֣�Ρ[�\�h��C�Ϋ���9�'��TP=�H�b%ۊ&��t���:�O��ʝ�j�w��<��e�Z�f��E���l���@6��s��ht�N�2麅S�%XÂ@(XVb�uv�����"�n�������r�uә��y�n#8`}��I靋��k�99c9���º��nW��T�fN쫰�G@λ�Pga�'�7������;�X�\�[	Sk��+�{�}��X�%f�dr��V�,Ȟ�f���t^�l+������KpR���Oii�H��3Õ�,�W�\�úu#�bē\���;;�3��P�k�t3�ų�"ly��U�1!����ҫFn�g`���W�97n�Z�d`S{��������r"۷vDs��7f�p��
�Y��v�ݚ���*ŗ�ܣp�N���y�9�Ү�q�>�%��{����Ai�H�섰q^�8�9��)2q����:7yv�5&-z֛A�d��xQ�|��� @*	6��@��pu��6N��7�c��"�Mm�{[��:�M7���ƻ�n:i�i�Q����8�Ռ�P-;;9�{:=;�mܹ �ͧY/r�;rTWW;���ڵk1�38�/l�c��+��p��z����W�%Y��śäӗn��!��3�q�nl.�#�!��x�-8�m(��[0u�h�PsH��:��	�������$�m+����
�r�0��k(]y�oXr�D
w^�c-;{-�ݧLV=>T��p�N�g+;N��[�}��$��e����v�'�l��}�{xM>�&���;����Z(g'"_G΍�w��[��%Jۗ�o����#���z1>W���zl�O�9�;r�:�-��������E�P#g��c{���^.�y�yp�2f�gXg�r@��C����2��"�k����q�`��;�^ȴ�ebQ�w�Z���;ze9٬	��*Osuao똝�bZ���������ޘ��)9ܦn��E��d��������D:~� \'n�x�z*���4l�*��v���1`̪.�g~�y���5f�9�=�DpT��0�7@89P�u�1N�*�]Q`ʺn�w^�����V��Z���,ղb�nKw�m�өnjh�����Mյ�ٵ�1et�{*LU-�p�9/
��]�]�����Pޙ�KSW�P;V̕�Fїk-�]{7+)�1�l3we�Qɐ�:�N�X�a|��8�ڛ}LnjZ����״�0�g'���_|��6�mD�/N�����gP�����܀�u9);����V���bv�na.Ïdd��\ldWh�Ey���K\96�iĳ�� ��֭%或�E�]Bvd��f���uf�����W:��(�s7;�R��B�\�n�n���응�q��6P'lÜ�Mh>e�ݻ�c��b t��&S.��ͽ�qŬ���ج��V�f�.L%4�i�ۋ\��r�Wbp�w6�X�7wasiH=]����^�=�Wo֮���n�V@*��T�5 4e�>{gq"�7@xy��~,˛i]�/<ou��K.��8\D�뉌;C|�{� n5%�s5�R���ʹB�/��m�!��k�yo�ᄗ��(��2���U���6���N��	��x�Evn ó����x���hף��6WzP�g��\����$�azey(9���}�B�n� ��Ȃ7%W6��Qq��8��<c�Df��'U�pdwh�)w�d��������ȴ�}�9�U�w�\э���o�7q��	�\�]��d�9$�\�VnoGf�V�e��G�D&hI�Z���8���v4�i�..n���(7��#{���[�rN�ge� �
��Š��:�[�PzNXC��W�=�c��:�_����D�0ݸaSt	���YG3q���"ץ�&#ϞjqiW�{��CFs�K5�X�)ޗ_[�wG�7R�G8ϯgnԠ!�
�p����9oמ��ը�S�.���7/v��"ޒn0o�v1^�2��Vw(Q|62T���b�`?i���U����[JAKɭzL�7�X�]�M횩w��u3�->	곏bذP�fJL7Y�{�F[����,Gqn���W�^�,Քd#��v�AB�:�k;ji6n����wk��a�N\p��A���W�B�FֻTƳс���&f�N�z4�"($͙��X�7�P4n�e�C�������t�v�p@��kANj�1����u`Ǧt�S�����ͰV����:Qɯ']z˕ཧ{���gm���p�@Z�-�s����}OsL��J���ӣfN�\��w�۶J��k'g1S�x�hve���r}��;N� �S��L-R�G7L�4]:hg~ћ�g'���YW=��DqQ��ʱ��afh*���yr[Ә�����k[���l<���!��-C�C5��D��4�/&�v,�:�)a�4��"�ܩ楼�n:A�Ѻ]{6�,՝�"�>\�6�=�s����x�-��q�k@/9�p��y%;�U��[�D�ۼR����y�p�^3DX;�
�[E�.�;�6u��u�T�SJû�3,�v޴`���j�уnl�c����;x���{7�vm�Y��?ct=Jl�w;/�l/=0ܯ=�un$�v�6p o[�ݯA*��plKY�f���\��{t�'Zʷ�d�Q�hWsQ�;U�:Hn��D-�鋓�A#��~�c%�7�|�cq�Y'��({9���Ŝ�{Ip�읇�DV����b��à򦒔������{�{�k��)�9���������8�V�:+��s��d�0ԞU�-�c��� }r��ݏOw.s8��Gt����Sx+[T�߮�ذѼ��\:��hynYJaF�'$�縫Ž���wz�{n��N�=7��wi�i?,;�6��U姂�r���Bg'1VM�b 2f�Qj�u��%�0CV�y�wBK�.�=ے�j	�Q�]m��%�r>=x�A�r>ͭ�XC
�Yݮ�+���t�q曦�\�Y���2�]A6M��h!���=Ie��y��.B�^�n���_;{R�a��N�q�i/7��8���O)�ٮ#�V>t(F���U��(9x�v�sc��"���Wn�h��A�=��h���qӑ�jZffI��H�w7�r����
v�ĉ��~���21�~n�3���N��g��-�^�������rk[z>r����w��rE�k�����J�p՜��$��;inmѧ+1��,���'������b���`�E���P����Y0L�r�]���|R��ГR7z�ޱ�^4q��B���y�ݛpK���
�9�,�������� ��\�m�yf�3�(�b�l ��^�D�e��q v�]���K�A_oa\tt34���c
w�ģZ�f��g��-j�gV����+�&>5 Χ���X���&�$歳����>��4��8�����ni�-��d�ob�Õ˝�3��<�,��b�\�#|n�uu��&6I����>K��1 !�1&��#y�/V=qnG�w2��yTA�t���&��ْ�D������L�ct�e��i��<p���'_f���ă�&�T�ͳ����C����UƨKR�*sČ!ս��a�n;b�R\��g���ru�p?Sۈ�2+%ss^r�p��U�l�����pw���^q9�up�5�R���I�}o�V�W$Ŝ���wD���:,ۗF�JC�`ü�3{{y�X��˰�n ޸�j't�:�<�X�*�r0V8I�g&�̤w;-g�,l�^���aS���&��"�����'�����\��R$�k�>F�6]�N�&ӗ@�����4Du\{��N7�SN0��ɡܯu6;�8+��$˸ļ5waQ�t��n�y�x�uH��0��ڙ� �C�sz�@�74U'�؇��x싙��������n�4KtU�!�fPf�/7y�]eٜn�/���+myv�kBԲC��՜�T`�
��&��uyV�u�^�w�QC\i�5]3'E�YG.�^p՗�׽�2B��V�i����lq#gj/��ls��M�X/+���A�<�9��j��	v.�^-��F���.%3J����a{4�ܽk���82��,bY�U��{W��$j㰯��'N��Xg�5�f�	KΌ�r�K����51�b�^��ñh	��y�Z��יniЭo�}Թ�p�m�������C�8���%u�yC�4���PFc�]�{��׉��6���%gt���r�\Lc;e������ݻ��#6��'�ױ����{�k��V��ӝ����Th��C8 �ӻ���0a�o9�"m��=5��bItbނoJw�1�L1,�m�+��	5}�K�����yGu�]S�UI�\W���݋�,Ц�+bÚ��Ժ��z�t�S���6��FY��>/7��p�M۱���vޜ��[d�v��)ٯṵ
�ntg26e���´�$n�-�(��gV��P͊<0��N	o5|������񛛓��$Nv���vd�ۧ{).bN xb�ݹ*�������Q�6�W�{�6�/�k�z˚�!�"%osGhם�K���ΐR�;���L�}}�`Z ��#�̥��
zܜ�&���5�n��N��o�\Ċ\�ݛ/m�l�'�jW�,�x�N��dӶ�齚�M�T�4%��ө�\�w�,�sx=-�=!�p����dկ^���T;:��vp[��=o� �(���3Oʑ�V_{�>�S��!޲U����\d��c���ГnȐH��80I;��[���&J�
4Z4őᗤa^�;]LN�#E=�w�^}�1od����k�L<���8��˻��B9]�ӓHm�;�^+�pg)����;v�ϑ<IМMn�z�����)h�W;Qr�5wL�I9c<����x���{�6��ʈ��HM���A�тq�n�/x��86�:tW���h��p�3o,[�:7z$0��BL؞�z]gI2����ҹh��5�����K��3�,ݥ�Ԓ��o-n&S��{o��潯�X�;��z�U�3�ٳ /.W�d}�mސe��ͷ#�E9���i�Zbcҋ����A7G�!��,Չ��G_��t*��J�v����K�	뽝�B7�3l��#�>�֭AN}����L�fq<�Cw�ܒ��ғ�rn�\�5^��;���ټor:Q��l��'s{�l\p0]����vAl��L�Ac�P}�ܩ��ƅ�i�;gG�CC(hsn��K����3�	�t��v�sE�io/oA�|h�,Z�ֲ���]���`y.��K�Q�8��l�؈Y7�E5��w�P��&���$�7�*����2�kQo ���7��ag�jŎs���>��dc_�C�E(�r1��c��G{�ٸ5p�X�9q��,ۗ7�A�:�C�I'T�{;.�^<	�N6m��9s$A��C:"�N�u�]���9��Iۢ�a�' ����bU�v��Ly75;_#����>B�=oq��e��9�5FK;��!K���5!e�,�D���]��b�˛�LVcK�,��&���LcRn�.:��8\]c�^Z��Y,ɸVdۄ6�99�˖Lہ�^�/�wC۫��x���ѷ=g�����;cFr7u�wMT���y�dyt;u�d�uJaݘ�+޷YݖǤmO�|��Z�C�BN�m6yh݊v��<䒻�����v�]\�J��=�}�@]L�)���8���ܩTv$E�{E]6ֺ��f�;U��FM�Oӕ�[�.T9n�ǫ�L)����E������m\t�r&��zf�څ�q!�t6'
� ����7�Eˇ�sI4$��w,���@{1[ّ4��ª�V�v�Uw&��dSd}���Z����;S�ZM#�g2����<<?i����	+!�T�
�H,
�� �$�� (�)*�$"�P�,!��R��� �H)!+HVI�
� VB,	�@XH@Y�AI X!!R� THHE �I%d ,!*
�!	 YI, )$X,�
H ,$�	$"�, �d� �$� E��H����$ ���`V �X @����P$�J�E$a,  P���I T� ��
��,XI"�I$�$�R (I	R IH��"�
��R@
���d ),
,�I �� ��V�BC��$����?\�3���<����gN��[̃��n���Ӕy��8�����Z�~Ą���^��G������9�/���@^"]l�d���a.���i��FOw}��>�X��И�<v�h�w���g�yd㣦�{��u�W<�U���۸}���n�˳+tp0?7�[�Ùmi�t{;�|BH�b�Wֺ�;�@�֭�:��9�F���Qv�ӯ�Rw�+騋�6���5}��ַ�����f��n��w^�����m�}��o���<����f�>gw-�>�uz��W`��h���h�4�3��z8vI�f�0[������Q�&B�G���ͼ�9{#Wjw�������t��$��q�[o|���N��R���Ɨh�slH���D�S��Y�o�~��g	��j���彬���,a����W�9weVS$����.}���:�\N��(��h͉`�/f�#�>��]��6r9�D�\[����og��9�t�.�:�EX5��n\�ǜ�[�n���&3���{�u��{3ћ���*��?"0_g4F�.�`oȲ,wJ]7:��gf��uE���8'Q�3��	���e�P���3D�-g=d:N��k����I���ܑ�қ��&��,��E2ݘ\�������l�����ȷ{W��t4��r�N��j>�=S�἟W�ᴻׅ�ٹ��������й"��"嚽�-CqǊ�ˉ�{�J|�[.2�d������������z5�@n���	<�����V`ol��5�|�M��Lt[N��xzvg7��3C��0�}~|fH����gNr�x<�����$���:V�ޛ����v'��N�q�-���2������vc{}M^冤*
ɬ���콯>��l��^G~2�j_77pl6��aϒ��ג ��r�G��d6f�(�u�l�/<�7{%s�k�<��0������`n�z5�]���Ng��QZ ��z��X����tf�J��o�EH�n���;]Xx�{�.�5f���k��Vs�]����\
W�N�s<9h��
x+�f-��������ObQ-��Qd��%���<|	fj[3�a��C�o��vCu���I��!ag*D�p%�B�VY�0�4�=s�u"L�%�"��8u�^�Q"���G�uǊ�9w��C���i��a��T~C��[�Y{^���bT\\gwh����n��w�>��
�X�/Y��|�L�c�]K��{�f��cջ�n]�;�`�x���#A۷sܯp�J眞v��n�ț���x�R��
��fLQ�cU1}��X����O]���~�>��e��oED6��T�"�&��6���b�������D}񊁺|G{W[U�25��l������<�0�H�ͯ�F�Բ��"\缟N��^2��]���V�`�<*nB��eo$�*#����;�5��T�$g,�;T"�a�*����΅3�C3��ڥAI5F��T��аЅ��Z9��L������R�~O�ԀZ�K8=�*�s������X�×�/eK����U�p���Uo���Ὕ�6�௶LoNS���kRJ�!h�ۮAf�>�0����q���?R@Ik}7iB�s���+ F��.�>�yU�\6-^&�.�wq�sy1�� v=dt9�7{V�6��d91l#�ޠ�7��K�`��0|^��A���Tt�0�,��ƃ1�0_xC�3͛�KcM N�FS׷v��#�oA=���2�Q�N6l���Ŵu�HCT�i7rbź��YNɪȖ8*�`EкT�xp��|=�gq��g�5�
]<�5G��N���.���r�����������C���cYd~\����r����S�&���w<�L=�V�M!{j�Qā�M�^�D�ݠ��j\�QcDܭy={���U�Q�m�Q�	�yANɁT3�2�NOL�ᚷ�=Zy��_�;(mi�7��N{��yz\�*��*H�UPuJH{��p#8nd�}ڼ]�<{;OM�]����sR��h�{(����-zzW�8x����O_Fw%{��O���1����p�N�#y��Ie�$�}�
6�jB�B�����l�CA:��$J�nk��P��9����B�
p�9P�{��R�����77���A���S�7y�ұ�����h}�îQȠ�%��s�\WI.�×���4N�}���H�\�G�v�x�Z��fc�V�7���Y�K]9��K<��k�JiǿL<ޫQ���;��_<6�ƒl��y&�K}�r��_�*���|�c��w(Z����w��{����_?�Yǲ�s�Pt��>�n�s�=֏-'������{���[�|�����t�n����,Qf�YM�*��p���(�ߒ��#��O�İ�!�dtOa�yHF�"�&lh4	�'����15b�eʹ�ԭ�u8�|lX����H9˨��dQ!���������8'ݩ�Ci�����]5D.�ه����[${���B����b�����b��N)��W�z����a�e��7���O.
�P�r:�gW�����m䔨�d[����������uP��{8T�)$�\�@���}8T=����Wib�v�b��s^<po��|0��mH���Kwn/eÿ_�[~w\�\צ�۱�l�8]�7!�(�_�~�/O����ʍ�,���TLN�r��UFK��T��U,l[����o�d^�l���k���-ۼs�6L�I�Ƕ���7�!q����v4}!*��sy��.��J~\2rk����{v��r]��ִ������R�3j1��i�#�^0sл��9$|L?-@�ZE�S���m�n���%z�"���b9ݽ'�s��\�>��H�7~XL3I�^Xm����*��^��,����&W��}���of�N|3���.;�,h��J�֥����O.q�:�i+]�6����cn�O	�3}L
�I�1���Gz��؍��h��7+����p���CZ&E��U~į[�l��{���77[�',��,�h�ξ٤���Hr1�/{×l<ur�{��`�/k[��v�Ӷ�;e8JP٨����@=7~�(��^��MV�U`:��y��)<��ug�{"��(z�Gp��Q�7B�S��"��]�:�[�Y�Mn]�K�|�f���-k��/+{^V:jӽ���˩dd4�Z����
�t��]3)錊ؔ��Q�H��M7ǵQ�&g���7�w�$I�G'L4s���1��gے�p�y��2^U�Q�`�m995�a��"y	�I�SvĴ���w�����<��|BY�$�a�n���������e�w�ߝ�8]�oH�gY�Px�S�1���v\\-Z����zG)nͼr��T$�{"W����}��'��:r"\�ڠ�3����z6'Buh6p.x�lJ��/^��CJ{qנ�p���٫ � n�E�9�i�Ś����U{�u�z�����k���~���7H���[��r�Y[�zC�l����j��L��(��g��=��uI�o	��YsI��cQ�������2�^0@��=�O�ID�u��="a�~���Ϸ*�����:f�Υ)�ss��,�8ќ�SY���c_d��St��λ�9��^���c�m���MϞ۱-��Va�VI�����[ĹsG����4GO�t�����c���엯�����wH��ٹ��*
��྽��.�l-�F�k��-�S�
�e=cKR�p�^ё�f��J�sB�j^��r0j���"�%("2�P�2O�S��U��_o�,<K�ؔ=�oV� ���)��'�{������N���Xu�
��	��E����w��6p"�kr_''��I�t�4t����� v�.ۥ�G��76�����O&Atj$B7��;tg��`b���`��c�s|=;|!~���oc�:S�=1�'|��v���7GzVH�{���v���FEޅ-Yr�n��yL�¬�.����-�`s�o����������)s�zz��S<�]�ViӅ䟍#CWq=�u�⽍��m���Fm�7&UF�����:���npRR�e��84RI��q��*�>7���vհn����7�s���$	�a����/	 �^\��`#��כּƬ���۝����yx��7P����)����1P�dH��Bf��N
E	��
�)�cyK,NmSyͽ�S��\L�nٔQi�ĵ�ՓGbn�������%F7��Ǿk�Z���bhf:ګ���A�B�u��8��|�fa�`!h���,����<bh����@�o.��"w�x�l�ؖ��`d�rm�VVsj؅�A���sA��w��2Ḓ�<�痽J~�3d|��;ws|_W}�t���Y��um�yU�<��P���e[�$�m9�h���j��]�Ӱdx.�E�=����%6�ś6fʤ��n���ݓ�����[{�(�����6�o�V��IY1���4t�fǾ�9AzT�˽��CO���DO��C�'���'#��]z���z�>�Щ��}u���Ox�S.�0���h����rm�ۊ��?x�di���>���l6��
�O����trğ:ȝ��5�y����w{�ڦO ��t�G�f��Y
�T	�b���n's�T����r��qrH��yqS�`=Nrw�J7Ԟ�vij�[��}�30�$�Bf�Li��9f��#�*]�N.G�c�YY�Bs^������.��_��5WN��j��Ir*с*�VL�v���&֙�wR��R����\�N��<J��6nu��*(>�y����љ��r7h��3Ud�&$���h8��u����Q��L��y�Y3��׷��1ܾ�=@&�m�['ϯ��8�A�Mǣ��]�Og-��T:�p2^^���jk�@ةX�������_�֒�gn��x���2A=��"��C�V<ȝ;x5��$tyi�w}
��Md
�-���f�E��Z+]x���;4i�B9�|]��C��A���t�k7Ar��o�4�L;u�a�Nݫ�4.�;�]՞��.������Ǆ-��0;Z����),Hw,������勥�`���x�� ��Qv��4 �t�η��p�L��l�̦ܽ-�{1T�k['
z�*���_!	˒ŷ"��&r���|sH#}���4�L��>4���`ky��,�+����5dB��ɜipݙֶ�� 6��_�b�^�Qt�& ���@����-n7�Ӥ�}����gsuT���Ӭy�	�x�{�JR�u�*�9?1,�{\vs��K��`ǎh����7?��X��/�^�T�*��甜%}��F�!f�Y6L8�j�:\��e�j��o���ǑF����J@�t��C��r��(-�b���1�E=Ul�#j�T,�n�pB�2rL�CD�Op�;#f�X���z=&��sý0��	�FhF�������;�ɦ	�0-��9s�8�^��gm3�W#fn�P<}�;��n��R�;��(�)�����s�e�������/`��6�u}��n�;�=˼�GbSßd7]���U骼��t����y�:{F��"�����;ۍ6fq��򍍷ݓߖ�^�{���<=��'�鶽/)a��R�R���a�)������꧜FC!���L1�ŝ�N^tw��!���<s*6�,��fN8|�)��y���{�|�8Q�'�oE|��d�+�]G�u��gg\9�d�@����+�����&�{��W7����
]�cַz��������T����y;a��<��@�~����:H��i7DSz�˂��)�������]y��#-��U\��L�����v���E[�����;BǨ���y�sTd
����Cȵhjv���5j�$�J�(��D&��/��%هICb��;|��o���.�R5�>����뽢��v�ٺ�0'T8�C���,��Y�s���"F�s���.1��^~�����s���za�µ�'��}5��ރ-b)욎\�V)���R���W��-�D��1a�W	�^���>�j�*���vJ���o�{Gj|7�z��_���It"tZt"�*4QV԰��c/E�x��}ݹϣsz��PW�-���w�.Lܑ���_ZO�n�(�z�ܻ>�1����d��t�u����!�9ǻ*)2�7Nc'6h�׀ہ�(a�E6�m����Skb���n�3u���s���Y6��I���f�W���k��J��9f�=������ӹ�L��+N���gn`YKo��T9.�F�m�����[ۄ�NҔ^zM�>���njI���]@>^Z	���/�̰T�"L�]at�Rc�=��3��{��77��=�9u���i,)V���M�'1umR�ܓS���V;����ӫ��}��Ƴ�_�)��Ut�O�w�����~,�8�V.q�K����|���XQ���Ӧj=��J؝�ё�蚬ZӓM�d�lD*����x��^۩CuR�MC�96jp���֖n�<N�}�M��解�&�E��c*���]��^�2���q~U�<'�ؤ�s��7Zͯ��$�֡�~�j�vl)�z����+h���˪NyW���5o�nm����[TC%(�5$�ӌ��k]{�dyc[��evmy�᝝v�!F��89����q-�v�/��R㹳���{�2�gG=~�"n�}��S٭*��F��x��Ѱ��׷h��t��!!I�$�̼��4�.��kZ�˨$g[�l���i�c�[��Z:6z���y�%�:�q�fa�K�*l�'V�����g�t�2�We0]�������9�YY�q����k����zy5qܦ��z�[qvLm����h;S	���[�.ۧ(�W
��.W��r�m�e��c:�������2�nMdۄ,�Fh[gqՃA����ݗb���Jvtx.z�Œўԝ���\t���ڻ �{s�ԶB�ݻg�٥9�&���K^�Inbz:�K풹n�l����svc�;���c���۷)z덭�=���[�]=���pk�����g��6��ۭz��bs���t���=\�:�5���b����E�{B;����c�=�mչ��"=$�[wI�n�[
Ҷ�ݷkV;��m����uה�q���;[۬�&�2y#�eɣo:7	�	X���7<�N��&퐸�]�+���+,a8j��S��]���ý��oWa��NLg*u��-�=�#�v�<�D�@�Ynˇ�3/�X����\��76�Yч��5��b�xi�v���'���u��c�,/h6뮰����C�=��ca���6@����s�8ݨ��Y3�/6���a�t�>��f�k���YR��H�n��>S�9��S�ι]���l��]�6�;���7m�v�Ńv�8v�"k�8�Op�1�����m�rp����.ն�ܛ�T�����Ӟ�ck[����q��/F��3lO<!�\[��m��7�Իl�u�6��k��=���S5��8����s.���W�Z��7<��O�m�73��.���¯'C��,xLֵ�&�<l�&�ִqe�Lk�k���v�Qj�-�[����}6�q������n���Pts�I�G �=���r��=p���������y{�}�ȁ�!�jPI=��Kv��@��+���b�����nP���p>�"v;��X;'aCu��ɸ�$��\pq���٩6Kq"cZ�B෱�ݫ���W1�m�`;1�On<13�gv��n7vv�|�#�:��k(Og�'']�{\�Wh�X1[r׎w[��3�{��6��v��2F���q�����=���b��\��9�Ig���n�������j�8��	���堇X��靮�=g�ݧ v���u<���toj;8�f2���Z��s�76��۞�Z�4��0��m�7n�n�y�.�.6;�Q���9��.ド9�m�;>���%����<���\.��/[�ۨ�'�q4�t���˯g��g0��Q�㵽��
�ET�8q��lp�/��h;q�zcSӸ���&u��s��;s���m��3{l���O)��:7k���b��`�ѹiۮN�I��P�\��=��L��={���I�N��zA�E�W\K�7��s���K��G�a�NpM�,NB}trk�����ڧ�e\縺� -��+��$`�1��Mg�/ f�/l��
f��6ml&�����]�Ԓ�@��ݶH#�ۇ�&�敠�:����.�p�e�=[4����nlV��c2�y���+o-{���:6�Gk��X*趨��۫Z<	��=��붷'k�^�s����н�r2�:N9/2\g��6�V��Eʪtn�7&�z1 �L��s�9�4��]�����1tƞn;=g�7Z��d�ugg���4\�L7[�N�Mb�,�m�3�E�e�:{@�Z1�K%�e��1�5�=p����w[�����7'rp��1�z���n3\� �;>o<�r�,�1L Fk�8�r��'um��b�f7�i�l^:���x�{7n�jM���X�}���c�c�p�$�Wa"/{=��*�k�9�3���E�6�1��68��k�[yyϞK���zn�]�%�;m��wcV޽^9)�m۬	�:�z�9\����)i֗rwn��cgʆi�<�9�ź�Ó�x����n���ز[h��rk�	��d�ƶ��֓��R$��GI�e;���'��-�Zaa5s[q����^�2�(��p�e��^f�4/cl��=S�Kv-=�uX��v�\�8��yî�ג����v8Ca���R��t�vx�n��p�p:�b ۮ-۷f˞�e��֭t�q��u��	��Ϝ�o58�4kF����^M��n�v⛧d�iM��c��s�9���,�wb��f��L���N]C�r�q]��Üu�K[�{Bκ��؞kd���uAeގƎ:Xs�z�v{�[uǶ�z��Q�cN�����ץm�Z���N��6�����=Q��mv��������Р`K�ܜ�ո�w�����֎�5�O��1� \�x�9cOd[��γ�h<�s�hݠ{nWGn��7Hy��u��6X��lD`5Y�En���z�ϗq�W�=�ΫNr��\������:ֳ�qg�h{>ŮU�+m�����/nn�Ո�6.��ݎ���۱�ݶ�&���ӓ]�"�;=�v��cnd둽[�����ۃc	�=�J�[W��7h׶�B����Rk+p�Ǯ�<ݻf��n��u%�ˈ���%%�v�$Dóz�a��j=��5�u�q[k�sh�q�ڸzݮ��S��ִ�GdʽF�s�e����Ѳ��iħ-�-���k�� ��c
nY�y˖��&m����9s��^.��x��W�>��;1�-	�\�٥���n��.7�{8���]�u�`��ܧ��aݹÖlk�q��8i{J�d��3x�(d��p�dK@FI��iB�݊�q����K����Sg�ir�m�۩ƌ��6Q�G�;*y�g�5���m�6k@�z����@eK�n@�>v�ܞ���ݻ1:2u�n�qt��T�:��5nz��k[.�Ժu�!�<v���������s�&�nu�ƓbD�[c;5��n��k��4��a:VPO#=�N�f���rlP:��$3͝��nHW����s�ne���@����ۋnɽ��[uF��ͻ8@�
j�:�E�4k�g�>�*[/�V�1�M�_���oQ���X'J���O�&��gt��svc��q�n��Jw=�m�S�tzc�I�S�:�[<�C���U<WC�.����<�q���A"�`��am��oB����ln7���,�8�v޶ظ�<BS �-\��#ۻ{T/���C�M��fE����޼Hk*��P<Ѡ�]+�V_Z��;�����J�6�v�C��JO8�]�z�آ*ꭻWJT���n�b��n�h�x��[�i�,��S����c�G��V{1�{��rwg��հ��؋c���	w��u�ӻ)��.�W�&�k��s�1�r�JƝ��V��x.3��Ga�$�&P'W��sۜWC��n��m�n}u�]ܺ����v�)͎ݦ�C�Y�[��<�r��=d����۷��6�CǞ5�OU�x���26���eK�5l�\u�wm��v�M=k���Jnnǵr[]sݔ��rr�u���=��%%���85�('BNs�{n��8��9�n��-u-`���5�&���\��v��N��=���|��	նݷm��%<��0u�'̅sn�Wz8u��sq�h�\��1��5���}��M8�y�/Yofu]��CXuw�.���W���[aT���cj{YʄH�"�-g2q�]���;2�g�"�<�x�^n�,qssx�X�g]���p���/��S�J��2=bt����'�*)��e7P�\&q�W^;n���v�9Ҩ6�mN��l�N�ݞ��l��=n�]�3����m/og��X�v��۰��o9�S�u��$�Q]�u�c5ѷKN{O���<����F�cX2��ڹ$���y˺0�In�/8�����]��u�rGlh�ۡ��볱�ۍ�v��g��M�Ǖ�-p��{]�T ����"l��6�nrnp����Z�n:�s�l�
�4��7%���=�v�şX���l�L�qc;v�`)��\�[����V��W��{1�bݖ���vNʫ�$��*�c�78�]� u��.��GZ;Zn_)6��4�'<�>y���=�ɴk���[u��$���{���w��K�[Y(����σ�R��t'OU�^K;���s�tܙ�8<���r���ȼpŻvF�ƣF�T�Zյ��mHݻ��!s��oDq���<���v"G�Gm����-��Z'�ն�l�crf�^�k�p�Z�G�<TN=��xm����˝q�S���{@g9��т��X�$#�N1yݭ����+��� �a��9m�n-u�;b�6�v�8أ���n;��nQ���.Rt�6���9]�+�>�v�U�=�o[
���k�ub�f1r��u��-��m��]��:����+�O#�nl�B�11�Wa�&R䱜���v�	ś\[����q�ϟf�:���� �U;�ܾ�aN�]m�y�/1�s�󚚷9xd�ގ��8�P��r!㚵��4�qM�ݻW����mm٧FdMú�]�9#q�&��/hmã�LqӶ�wcY��H��/Ndz�^�;E�N��Ey.ޮz1/gpų��1����v�\��yf;�n9�c�q�[�(�w<��m���<�G��k��d��m��n�\���ո��%v�G��[�䋀 �Hi	�h��՞���䍸��	��K�l*��&5G��XCv����j�G;�{FYx�fc�q�5��m&�6���Z۩y��w6烒Z6�ηb�Ku�n�����7n��6Ӟ77[�c�zۮ���3㍑�d����r�t��'s��\���Y�`���]"��F�kGugv�t���N'�����x5�=m1	�a�Z��UZ�A\ij��*%���a�pG��۔�̢%Qcm�[Z�e)Z�QE-��V��-������km��h�*��7(�(���.\���ҔmKB� ���Z�Z����E"9�dkZ�ڶ�4�P��.\��b�U�k����-�*6�T���Z6�m�����B��!E[eZڍ%��m��J��"%
�aZZ�X��Qm��E�Dke�JT�J�m�((�[E��mZ�iK+Z1�Ѷ�,��e�R�Qm�E�l�bQ�Т���ҍJԢ��lh���U[T�Z�آ����-h�*�h�F�F�j�c���[-�R�EJ�(U�[cT���mR�m���-KF��6ѫU��`���*�lEbV���Z�ikT����)[���"YZ%�����-F4b�Ԫ���5ih�����jV)KZ+T����Km��l�ԥLB���,T
�FԢ�U�8�Uie[j6�Yb$ch������TQ���m���Z"5��Z��Z�(�j,m�JZ��)s
*��e*V�maKaQXĻ$�u�ަSuf.,�Ŷy������{qm�@���m��l ��D]�sg�v�2AN����uS��Q�����]��q��*�b#�NG����<Yۊ��2��ᧃ��N�=`x;lk�%y:����h:�cMv�Kks�<����v�m�Z��N���#��Gg��y���>�攜ӻG�v�c��7J�=����hm��6�9��Fm!��v[��6M��r�ɂL�q�sr�ն V3�\�^����p�`�f{r�m�񶹬�ն�{6�pr�v:�%s�tz���.8�A�බ���n�4���rv����ۮ��9�����돬��l�9�NO���k�c�hÛ����=�{p�bV�Q����K�{q�v�.䭎�v��`Җz��	�.8��9�CQ�φ�����gq���;���y^�Ǳ�8�ڱ{.�;m�q�=ƭ����nǣ�v�<�s�*���&�)�tC;n%N3��Ѷ��q���g^�; n���ݞw4���W�&p�f�#��g���)�ڮn0�2r$���C��nĆܝ=�Nݶ+u��;�?M��ޝ�x�P���<�a�c�\�v��yؼ�ێ^�Z6݇�ݶ��c��	s��v��s�ax�;Vq4g�\�7[���X7	�����﫭�ns� ���/u��}<���N�M��;�WZ�֌��v��g������v5��:�j���;����W���֪ez}/�@j宬�h�XJpv�'f��[V!#�����!�u��������9���%ۣ6ڞ��h���qы�O��y9�nL]�f�M-F�;u����b��nl]���;3 �ѫ�m*8�6�@m�&Mq�ݻC�g�B�y�����ە���n��gN8�ٵ�\��q�Ҝ��]�|c�=�'7�Z��g��3�m��q,�7̥ָ��n#�;lk-ݰE��ˮ�uN��w��y�������c.{�M� v�Crq����{��YjڎƮb�R�K\�R���(g��v1�c+�ɳ�p̋�.-�)p\�cE1j���8rgÇ�p;q��T�Þ��<���ʉ��Ȫ	��y28��r�e����G>y�v���T�m��+��xW���3��v�=��9�p��;r����C�w��p<g�������v��	 OU�ȒI"o������Siһ��|{�.��{�o�`E�A�r�ʑJwb�_@�3Y�!�d�Z�� on��6|�3���A�$�Ow���츂���l!l��\�B&"R���j���4��H
s�{|�ئ}_d]X ���4ݤ��&��s4������PE��O^�x^���mw�|�=ug� ��_b/������~;]�{>ٻ+�=�pL0�YQ
#l��=�꿬}����=�\VT��G�:n� ��i �/��iY�;{s�tǺ�_��&�Q2�C���0���Z��딼[�kd�ۮa�۱����+����q���\��������8�����wh�v.ޝȵ�ղ�krmX�^3I���rC�������B#��'��d�f�qz2hCh��ł���rF¥�-\l�U�s������ߋ�r�-޹�,9���Bz��k�,C��s���{;t�P�3�g/ɒN'��MbE�z��++��`��ٟ{��z�E�ܵ�R����_* gg��� 2�(ޝo_��g8�O#8�� {�w���(�3$"a�%+�o��+	��Kܳi��� 6}�ͻ� ���s����\cԀY��._w%SX¼�[��$|�v��r�����W�yķ_ {���b����:�8����}��ka�s<MϏ+zƬc�s�{��c�g�.�ڃ3a��D����}-�0L�2���%�� �Oɲ ���<'n��;[<���{��j��R�q��8��m�u���]�&=~�Vr�{�ga.�H�u݀wlڱ�ox��G�3l��%��
'
�Yv���`����V�J��=^��.H���~���YR�h��Ogn�PX-P�	�
����6��m=�qSb�D^Ci��W7��;;��2OJ~�fn�7d�6�{�y�lA��6�>"�8�m�jeȥ;�/E�/J�4�Fs�y{�Q� �t��  >Gf�ݤ�����Y�$u]�x> ���ńۍQ�e�'0��_�������i�R�V��ݚWq�y��@%u]������4�v��8�H.���b��U���HY��%
X����HI��Rۢ�7n^�1;ys؁���������D�S��F�w��|��۷V�@;9�VG.�K^���1��D�%�lڰ����[�\L��\ZB��*��EN�F��v��ʽ��� ��5`|�OќM o;�ż�L�.�o���P�H%6	ħ%E�q�v�Y��g۠¦��qwiO\t{݀�~���v��P�*�9P�8��r�g���<���! ;=u` }�g���ѹ�����V�n]j9-�v�FN3 �a�@������N�� ��-��b��Oێ+<ݨ��w~�<ڄ��r�� 0sZ��%��7�{�5�0��i�D/�����̢I�F��Jw!l_����Xi~�w4b �͛��fq��}ىa���ʭ�P�����6�Y$�Bi!A�����ͦ�4H `�bυ-������|��6�Ӹe+���u`��+�l�o�3>�V�݈'���g�,#<E$�s6"��15$T��%�v&2	/���t�[�o�nvU�b�3�R�{7ݖ�v<�Yۘ��M����7��N������.6�t���|�3Ӿ�J�9f���{����Fx�@ >=���y�ܥ*8���7��6�3��+Tkb	faIH l[���b �}�=�\M�\�
�%��&��2�u�ʇ#�F���r	�^�^���ˎc1M=�\ܿSc#���{�x�m��훸b�����ؽ[�	�-.�phQ�D_���xG(Ms�3����e��h�gUC�`�ce��;�����"�z���_�����r�ڎyR7N���v]���ڶ�p�}���=z�ݛ՞���4�)�L�Z������+�Em��w=	����ֶ��9��8�n�:�ɓ���9��;c����[�lc<�n���g��^��Mj�����n탥Q��K��Y����ux�x�GOa�)v���[0�V{b,T6�.�c[��j2���;�&��!�	Գ��җY�E�8;��NI�/YƋ����tq�q1SgiI�ԑ��lcE������n��I"���/Hu�7��X |�훴�]��w�}��H�ȼ"�Hf��3�	�<�K%�PȔ���ݿU���!����d�r  /��fg���zo�c>��=Z�=2F �wH�8�j`"��]�m���}ug�$�q��˼�:N��	��m��3��w��:�.Jp���"B��.6��_����� 3}�^,  G��7 ���o�mFz+�l�/{��Xt�]�P&�S��������3��������]̀�s=��m�o�Ռ@%�3�n&.�u�;6��8�c�9�(%��m��հd���j�s�l�J���J��׮�:����s�Bd|J�S����X��w��π��REw���'׻�u��S^x�Ȃ^vՕ蕄̢�F��P)xF��)H ��c����o2�w��2S�����QQ��+R�TRJ�Cy�,f���3TݑG��]k�
 feVl��Mժ��T3f#J�^����	��݁��O8� ��r�|F�v��⛓�b�	�dJWh�uՉ �5�� ���_�z�螊�o�@��i��O8��i�
&�d\Z'{���ӽO}p����~�Um��#�R پ�f�1R�˽�krJ׀_\ڰ�t�ZQ(��&H������DD�w�'������v�16" F�lݠd���g{�>�ݸA�v���[���&�"b%�MK�1Z B=d��㜅c�8g��+l��:q�������;fS���FW)�|��#�){���ςfw!w��śRLul]�.2|�e�듟��*\U�l�vb���Ng�����d� k���?{7�0`c�.M��Wt�
S�3�MA�"�K���]} �3s��;�>�]�z�%���.�A��[�<PGٻ�xw[~ې������=�����g*5d��'a�+^Z�ɳ�*�j��=�7��#<Cu��7���rh�Ƿ��w�'�ߩ�[�5�`Ws��zC��_�{3 ��lz<�>ɞ5H��:�n��i�dB��9N.-"{{٘ �۱[N��~���u�c+�P |_f�f@#cݱj�	�ԩÄ��� �x[�#+�W"��B��'dcM��Zw��װ]3\p�_���O��ܴ��.:ʑ�;��m����b�^,+]�lצ��R �����g̞p�����Mm��|�\
�譜"�y���A ����f l6=ދ��$�)�"ֲ8�A��W'?D'
T��H�U�b�� ���S`��t��/����|���m���ЃǮh݃p�{�v�>�߬VJ�_�s�~��^`$ ���[v�H�#
[{]�CȒ����{����ّ�Tlsjû�����0<?A������o��;ǰ������&m2�D�xky��&�o�� ȏ)Q���1#�L��Í�\ؐ�4�"�ۛ}�cl�G��ŭ"I;��K=�gA��׈�����'銈�C������ٺ^�-�-g	ymk�����������G�"!�@�8�q~ܿ�6 �F��� �H�"�]�{�Q��l������|Z����D� Q.f$./�\n�g�ҫ'���w���}=�ۿ�Y�E|nnM�#.���ښ���29Øj�JrT_��J,@�8� �
"�Ulz�ښ9d�ky 7��)�@i�7WnUrr��!��K��r��6���*��v\[`k3����+���K�xu��'N�J���Xڙ2ԧvy��_H {�y�����S���#!��{�Z@ظ��(ǯ7�ª�x�=��t"�l�Q1��UK�+�;I%07�N�'���nQyY��rb��۷yǚ��cvW�酞��"ܯ>��65�T�~+v�Ǯx���	ȡ2X�O�h9{ns��.��6�1�6Ӭ���==��t7;�;sݘ���Օ�B�l�7e�:�j�p��T4��<�.�gq/�|�;���q×`;%q������7+����ì����J�g��s�.DK�\�l<fg]�7X���M���:8��}�]4Sͻt�=Zb�gui���ןc�gEm�Ⳅ���-,룡ۗ>�[+^�^�I[d�Z`v{*�t>1�L�]�7��|�ڣ8�{�7�iM� �f���7�1��'y]Qz���ϕ��x��Ҝ��JDC��[qqi��f`���n�g���ۛl@a�R ����Ń�R��st���q��Fp��Q(�	�\Y.6�m��{�0 A	�1F���k��� ���������4s�?8MD�%Ť&�K�Β����r����vf 7�힤M� ����̢) \��9P�n!�R�����x =�m��Ҫ���QoT�ȟ�TGa���7s>�� �v�<�tN*���E��"z��$��]���!nznG��H�b��x9��e�*[�S\������9��:x���H؃;;o0l@�ٻ�9.9����+�8F��g�1`|R�,��s28sZ�@�{�V�~��#
��2Q1.�Og�q�Gм��$s�9��^��B�T����F/ot��������S�V�>�JF�<nT�Yt��ٝ�m��7ݳv1�q][מQY8G��{|T� na�l��{{٘  {�۫> vFf<��/�4U�����ϰm��훲=���!�d&YP�E��{'���	�{�0 �l��H�"�tW}ȳ!���ٙ�`}��C'�	��丿����[g���+�B��q�_NY�נ(���0��6�bi�6U�T���b�K����.���gԏ]x��ͽ����m9)���Zak�.Z�b���NT8�jT����������� �gH.���u\��M���f}�lA�v��%v򛅉�N\�P�ٮ3��C੕�'J����������ݠl�3��n�/ٙ�TVo^y`oV}.bB��]��޵�ؾ�4�@/���<����ɼ�z�+.�CJ\�M=�f���Z��߳N�3ω�=ۛ����9��'��9�,���<�wL�I�����r��i��Uwr���wU�o��o*�r)�r����	�;�]�xz��xQ��K�塂�c}5�J���=S�x��.iMwh��WkD��o�܋�=����qf�ǿ���C�ڦ=��`��7Eհ�Nu<QB��#S�a�xCF躽	�8�M۽���'�N=�\��^�`��|��`fΨ[pYQپ�֗1O�������Tq��o���ww����i���-�����ѸΫQ�uX��!�Zp��%��;����#y��*���V�K��y�N�?P⽧&s{m��}�y<�ͳO9e�z��|	ӝD)a����=^6 �lڏzn8D��,�9��������MA������������
�g��ޔ�t�>��!�;�ݸH�>@�g�C}�ձ�{�Vr��J�Җo��V��y۞�P�W�JuSq���H�'b�{�f�ŦpUc�&xSB=5���5u./��M��v6����b����e
4�&rA���ž{�=i�>��@}�5}��oc>Sޒ뮏g�Ü�kԴ9M;�^��ZS�מ�.�'�C{��ϭ�����ݯtѾʈ+8��F���ڍ� "�������z��u��(S�)�"���{cW3������&�KLL6��0w¾�!4��-�NQyg�㭍N�s�J�G��jQmޱd����:\��(g��)���`��5�dDD�	[hѶ[P��խ��6�AJ�PU��Z�me�UamjQ�)e�5�µ��������d��-��m,Dm(��%���m�DUiZ�UAQ
�Q`�[KZ��A�Tb&QZQQiKڢ�����Tl�hUh�Z��ei-�q�a��U��U��4�X�*5%E*Q���J2�E�6�ڣDK��V�ʃT�F�TV2���R���-kZ��V�+YESe�k�fU�E�����Y(�lXѵ�DZZ���h%��W-G��V(��Ub[Z�UJ�X��*���H��iV�E-*f\�m���jֱK�����*�A��EP[h�����
�Z)QbF�ڴ�R�
-iF�T�X�c%H������b��eQE��Q-��Z�Aa��DTE[)R�X()R�DE���Q��D���-J[k*
��F�0m���RҢ�UJ�-�#mJ�b����b#mq�������+Z�KmK#X�Z&��}u�m-�����u:��FqӞډ "!�0�\Z'w�6J2�>�H���\�I>6���$��;8�@|=�ݎ�7D��<�vy�@""��j�F�:�r�&Be��.6ʐ 6��ml,�o<Ό�o��s�v #<E �G�;�>Xx=n}����:9����s+��C���=����u�
^m�mvlu�l[��mjP+�����b�{sv���MlU�|������@��&�Q}��ۑv6ϼFi���GZ��p7ԩsvnU�fǺ&s�d<�����ba�R߯7����)E�T�j��H�����B���q��|����o��~�n���}Q� Fi� ���g��~Y�D��"��[ow�5���k/JR �߷�1 ��N����a6J����f�S�r;��ܴ�ً��rc��y��2�7:��"��/q:��U�2&��t�(ඊ*AfaU�2���=�P}�I C���ˋ'�ۙ�  ���_>]U3��<� �g{�Na$�k@ �Vc:��?��������v��۪Z�7V��O�M�n8Г���p����3c�{p������|�.�X�r%Ǭ� ���v���w����#7�w)��x���!�}ݙ��5Hd��
%9.dO�����,��5�E\20� ^�fb@���/(1ucj~Q�.�'}ʠ����sv{*�3  {��Ո�=�~��GeE@ �_�r��}ޛ�WxQ9D�R�;z��=�"'/�A{�e�� �ޛ��H�!S���x7|ߤmv^,��ψs13-�+���iU� �Ҕ�������j��n�0���ٴ�`H�!����1zz/h��g~��Z埘���p�J����^�L�Oh�{����^��nU���-XnA�ñ��/�X�ص$��m4�up�<�%n=>�$7m���9��y6�F�՚ۇ�˶��s�9��丣�2���u�n�3�;usA��Ϥ'�.��-ϣm�N}��^��/X"�9��W`�s�:ֺS��mm�m������I��s��r��ɋ����æ3o$����,5�{]{ m�뷧���A��kv�]n�Q��!�DT\�띗�}ywi��dl�2%4��S���'ohxc����蘇ӻZێ��{,��vƇ�&e��n�@�I�̎'�ۙ�� ��Ո ��EC.%_����������� ���7e{���r��4*�\�"���$�����f�}��V��v�7`i�7@	�^z{�VўF�)�D9D����ګ��+� h�.3�L߯l���� �vͫ�H�H\������C�䛿�����}�Qk�4ݠs~� }�o�� �f�[u~���L�%� :�&��s�XӔK��vs��JA|�������|攞;��Y��sv��H�@ _��3UC��t���6-�d���� ����`t]�u��8u�y�g�������������l�_��ګm�f��@ >�f�c|���/i���AS�M����(��$���b	m�N�nf )�а�^P�bs����zgV��	^�j�T���t8o��O�7��n v�T$�;�P����'�Ua�+VG�zIk�u�U�|��"�����٘1w��:s=[ݝ=`�86�r�J�%�K�� ���u�� У$�����@�w����_�{-�O��C%��*`��8۲î/�Rqwf��ٖRRf{;s3�=���Jki�φ��I�PnG� Cp�Ga�<ٽ���p������\���`�@x��(=���`�>glݔ�ec;�ϪC�ט��Cc�K3���A��+��0�<����]9��h8�`�
����?�tb\�0��k��R �7;o0l�����}Q���^�:��'0�/�-v4(�"fe
����Z�>	�
�x��ކU�� 7;�3� gl�w�V+~���׷=D7�;v�! 8�	m�Oong� �ݵ�X��~wθ_[��������M���ټ<��dפҁ��A	V4�5=;��1��B��j`����C�w����1n.�ʚy!�@#��v[y��티�pOBr�hQ*T�_ĸ�'���D+�8u���>�;�޼X6���7b���#(�ɒԨ{q��vf`}��@9�T�e��n�M�$��3O��ؔ����31 63v)�A��H'��O�[
��25�Bn\��L�p�ە�sQ�%�]����g��h������Ͽ���,!�8�"���zr�3�q��V�H�w�nG�4ʿw���	���򊌘b��g�v�q�)H몇ѷ�Mz4��[Y�I0��R�D���"���T'y�|w7�Ϊ��E�<L�D�( Wa�gZ�lf�� >���Ɋ���5[���|to�)��}�w��^Ω c�1JeÍ������>�-�����jl@��Hy�����_��3e��3H��=�ŉ�Ϯ��K|t�:�ov�Q�
A�K���Ӽ2��_�1��3���*	țZ�mj��+2@��=�>@Wa9����@ТT�,�K�Ҥ�{=�ml�'f�Ϡn����@ �g@ >/3�-�S��^�~��u)��=��{ [ZWA�w��Xl�m*�����nx���}��-����L8 �]͈��e�wf`E�K"�6�
���#c�"�n��)\�XCbq)˘�Z�ع�#��Q��V�%�{�$��E|��3z�Qѝ.�v)ڿQQ����D[�/�m����y���Tp�9UOF�`-#<E��of`|]��ТI���
��vv��u�$�	�ĀA��))ff��y��n�)�*�Q[}�d�=H��aҟd�I�a�S.,���ŀ i�����{�Uk���"�@�����$lv�Z�1o�J�
	�&�s��V^/Q���(ֈ��C�7��b2w�`����x{���z3N*>{��V�اq�s�z���=�s�.~!L#rU��q��C���,�')7�3���YeN���C<6E��p���b�7H����  ���u��NwzYN��.��9O��X��;�;+��G�J��<��!��Ob�x'azvtڲ8�L�z�t ոv�ukQ=���{���ϫ���|ڂ�Q&�4��F��S�v^�s�[��d�v^��*ڮ�&�,�IWn*v4���]{�/��W��k�NpŨ�7S��pk�.��x���ߡ9P4)�*M?���)H ��^`$���-��sw�.μ�gi� �f�b����-����LZ��� �vR�]E��S7��  �w=٘�6��t��"�e�)���قk��}t���b�_�ѻj,@ �K;Dq ?fvݷ�|oN�j��	���~��8�&�� #o��� v��v��"���M��ۆ���٘;�`Q$�0( Ua���E���R���:.P	M_fcm�;��݌b/�)�K�ʇ�Y�������"&%K�&! ݨ�ųt��Xdgd�����[�Ϗ3��"F�~~���LcR�)��;��İ A�l� ����.'n[����w�0b#����>�pOBr�hS.e�.2@3����Bj�+�����*6&(o����!Y&�ڞ��ϴ��匔�c놣e���#��6ֆ˅��阷��Z��
�4���Y����o[6݀�*AH ��՛��CS^�t��1a��[*!�$�����H�zTt�@�!�t���x��NUM߀��.� ң�n�����ln%51ob�����ZeQ�F�fGe����=�?fw]Vjkgpi���������`��d�c�&~�h�dtW�6$��x��r>�����x���7�� �������g>���S�ȿ`�(��|��Jd{{M�[
�ĽS[g�]���G�j�u|�����Ǚ�)����\�`iQ�I@ >�|�xDg+$!g/$�T�r�cf려�l�1���\Y;����Vŝ�>|�0�gM� =;|���of1�U����#�بQ*�2�Yqdǣ t�A��u�� $�O ���s�M�������$��w����͓��niz5��9u�%k���Z8��k:�Ӷ�̱���U'S��*��F��b��Ydp���&O�_}��[]� ߢ������߯����-����\7N�����;g�j��o�E��g�=����{b�h��p�Kc'�n�����ln%51vl��g� ��횽�<�0{��ȩ��OA@���Ń> 3{fՃ�}��ϟ��*w�.��2�<��ݬ��u�kA��8�`K��N\��pMW[__����4�d��"��P vv�`|���w�_�w8 =���g�N�@|���İ�c}�NH����Z�m�n�Ƕ�����I1q�l@g�ݙ� �o�fՌ-���+o)ϲ`��5��) c�1JeC��������v�X���TՑ�x>3�ۙ�> 7ݳj�G��S.�2�YqS�I�ׂ-�$�?9��s	��&H2zb��U[}�BŸ*�"�Y�Brf�����S�^MoM�'Vb�=F���ۼ�꣝��Gi0��-^Ij��͟B�ҽ{�{��[��ٵ���#�q`�kmU�$d~��1ҕ)�(��vf ����3��#�l�S��{��?y���`" S��dJDK�>1�3om���\�:h�e��Wk��խb?���ќ	̶�"k�F���` �n�_� 62z
�6��Ƿ��m�7��N���2�	��Eٱq�I@�F򅼮;.au��{}뷠 ~��Հ�OAI ��<�g���oy`|W� O�"rD@���w���dlW�6 ���qӝ�3����c~@n�mX��OAH	��r@�S*)�œ���ދ�̿}�[��`篦���	td����#>�W��N����q'b6��
;�EB�p�K�e������ ��9�7ۿ�yt��(^<�%�����'�6�$e��b�>J�:X����P����T���c��ĜąiM���8tW#�p�0���̄��6�NO�Ly�Vf-o�l+T^�ha>e����m;����E��$�[���+^Z�S8v#�� |,[�3�u[��W4c��Oӻ�(fh�azpSv�
O�ΠHU��Z�Rl��*�����#Ժ��X&�;/�/�:ΔpLi��M��0gC{�\b�Z�w�s�>��Z�gsLЛ葭���w=}ժ4�b|o�W�9���ߛgzNj�'{{��������s����Oy!!\)\3WF�����s�<{�VǶ١�R�p�Bv�y��+���xs~,�ew_����U׎T���o�ʤ�;��w�D;)ݼF��y��Z���kw=L���\��Β����edѾ����>��ɓ���`�����W�k��ն�X�8�n���jz�)�r\�UK�Ue��ii՛qxW=>�DC���C[���e(�9t��/]X�MD;��0�j��CM�T��ޤC/`��Q�HT�y�S׆s�۸���Ī�ټ�g�ڞ�UDȼ��4 ;�s�;���DC�>P���^M툭(;j�9t��&{޽��=z��r�]e��94d��tW��7_���^>Y����7}�O��W��0e���N(V��%�2���{����1LpJY�zvҷ��N'��֫��*��sw��Y�7F�Sմ| ���C���gk���ʧ�·mxE���nq�{{íҷ�ns[�3h��Tb��*+�+Z*���AYl��ʢ���A��t��V**e�Kj��ĮR��iYUkm�ʍ%Z«D��T+UF* �����ʖѭY�T��S2��TX6��YD�X�e30��Q��AQ[h��b���QQ6�-��V1H�2���������Eb* �"��*�R�1��*�F,b�T�0������[E��"ܷ
DEE-(��1U���KUJ%����X�*����A�[*����-��*
�R���hʊUJ$V(0��T[j)�Z��%*��+EB҉m�b�*U*[
Ŷ�1��Q��"�Qbȩl��mK-X��F,Q��ҕEBԣj��J�J��X6�Vڕ
�*TX(��kaR���U�cPX�j���4�r�EC-`���b�*UjQ��K*5-j�k����X֩e-�PYU+(�Z�[QUEb(�Z�A�(�j�ee�RҨ"+kV(�ª*�#TUD`)(�-,�eee�dA�QlX�F�V����%�eh�TQTE-j(��1e�1�Ki�bUX�
,�Z���*+
�)-%�-dK@��h��fLK�Z�~g}hn�5�TL�H�%��r)��]�vx����ã���j���<sڐ�w�,g�>�rU���X�.��!�e�V6�����/�;\c�v����^7Z]�t��\���z�v��:];c���{Vnݎqǎcuq����A�3���<RJr7�0���_a�贕#^�Ȫ]=s�9� m��"y��h���:��u���v���os�����g�S��a�vӥ��y��_c�潋��I���N�w@n��v�t���s�u#��j�x���]��8l���/��v�>�0��V����GQ�v���炣6�;-3:p�q��
�vj틫1Z{��ʙs�c;�i�ݐ��x�x\�zŭl�z��K]��t�;k]�Nؘ��i˞;��'.��N�{U���ڔ;�5�&�klN�6��范����g�{M]�>,�қ=�s:q̇=�����F6�+��u�=G��Hz��vm�\������e���+��!�*OoY:x��̾�t�2����ݹ�y���t�n�Z�u�Xn5#��7c�n���Ox��vZ���'P�v��
]�����s���og�:�u�]��7F�z��3�Iޭ��Lt��s#��b�3�D�Ogtv��8$�&	�0t78�����ݐ-A�	�Л�%�5��\��6�{w&���J=v68�p����˜�ŭ�����Oj�yU�mhm�8C6�1�I��P@\/-c-��<���/M������m��m�����D�O!�����Me�����=��듵���v�6 ��w�(����u��I�a:�9�h�wg�\�:ٴ\���]'`��Ѭ���u՜n���w�t�I	p�C��;v�[�k�Ɋzݛj����<^�MCǌg��k�vC]��7��=sv�r��-��Ƚ���b��[�ե,D�Q�GN����z�,ks�4Ls���j�bP�t'W<�$|7��={3<��b�v��z ��ԗ������X�{��ng��b8ȱ�rf�g�>�r����i���vD�6.k�llc�ջ���۱�=@�JH�荓q�y범��g�y�7�Y�"�q�vb.yI�/T��kRl��#�k���d��g�ϳ���k{-Ѹ|�92Q���8�-4l�۴c��n$�2��n�]Xػ���tq��6[��5�,�4R\ӫ+\u,9x�I��,Q�=V:��mף[��^5�z�ԠW����?���CqG/c���V�[`q��P ٗ�٘�=#�.wbj�z�orrs����(�彵#�	̶�"n�M�f`|c�$�8}]�H�N�@ ������9_�w�7X�d�{f����2�	��E��3s�� >��_�'�'u �'�7@�3z����%H��@���ޮ�Z�T�\��G�t��wf�cm����37J�/g�<ߒ���l� `*�0(�B+�<GDD�V�+�^����� ���ŃlA��4�ou�۹���k9��%�Lʒ&�(�'��Ɣ2^M�c��n���x����t���>�o���՞1h�g��0{"�����u��m�n�Z��f�x�z"�"�{3ݘ����R6�Cp�[�P�&vk��97~�Auۡ��j���'|C�Q�p�D��>ޱۚ55b�ȃ��U�'�U<��݄(y�9�|v��Ca���n/�	��l��>K��|_�n?|� @}���0�In��+u�y�V�f9mV̸^��\�(���w���ϖ���nګ> .J�מ��z��\�G� o�ݘ��7�fҲі�"`��3��6轋��r����Q�{�x ��e�Xǻvn� �Έ��*rrres��z�����[�mD��D
�wz����R���U�z�<��P6���i�@-�Έ����^,���[���K��a�ܩDJ��9�h㞍�c����ß#��D<�����qQ������"c�
S��D��s>������@-�Έ��߳վpۿ@KߏV��>X0 �劣Ǹ�S.�2�Yqh�7"��)��ϯz�`���M� �#:"��Q?W;��[��L�	n�l��U� �Ί�@���b����@�'h(ټ�X��lDBwG`�s�α�`l��Hl���&EA��'$85�]�So>[|gK������2ݬ�����gZ�0u���x{�d��g�����i��������뛟�j%8rDݣ�W�څ�6����E,�� m�ն >�d�@��z��o1�O��>yuL>���I�|ӧ��@�~��Z�3=QQ�v�+@=��vA�#`�l����ł�.����?~���חwݶ��7.��f���z�n]њ��瑃k�4�H�"-���ڙr)���������4��� ,����1��篬��K��l�m�FN�_ �Wm8 h	��������X7ʝ;٩�p������]; ����u�N=��Μ����"��S.T�Y1��P	~�{� ��=��TU*;�}������Ł�RX�dM%J�3v��,U!l]����z:)@| =�����{v}���5�pbzw�z_D�5���2`�f�=���.B�'�=3w�E�,-ID�o%��K߶M�Az�-�Kｯ�~����������8r�rDݤ~���K�=��uu��{=����~mעg`n�fn�,���7���W/_�j����@��(�IK�)�ú�9�����C=��dۮ�[b��Ҝۣ�[����㉈�󘟢|l\lRP6�nvݼ� �n��\��xmw��nDT� �we�E�0ڙr)���vl�\���cy&�E|�ϯ3�3��PPIe_V��
�L�޻���芠ۋ����ܷ�|�Mݹ��zk��:�6�'��� ����0��f��C��2�IE��{�A�x�"NxDGKnQ(D@�����K\չF�#����Nܾ�����hz L�%6~2:�5q����yw� ~7v-X�== ����=�#�Y{��Qs	8I�k�ڡ9�뛞����t#4�����t��M�0W�!n���U�����HY<ɨ�*���J['�p����R����{���^��8�:��^2�k�8W��\�}��Aq�}���P�Gu�r*v�p=��h�n\�<ۂ��l�#Wl/�}m��;���e�vx��K���� ��(�:OĤ��l��.���-�Ë��"i������^�*�/��0!�@vM��ݍ��ywW�������#���5r�;+���u���Q��+][Vm=8�E%�<t�»e�.;(���.�}�����t*X�v���h+ی-������ב:2C}����b����݊��}���{*a��ô�rb{ѐI�-�J
a1��'�V�E�E%}y�gW��ѧ��}����z�tv�[v�����s�{b2Tՙ]���E���2�R+o��ٰdz*�Y�������{ڐ #c�b���FOA_��P��D����N�ny>�T��7%v\�� 0���	���F��f�yy�#�����D9;���Y}�g�I [o�>�@Â��Y>@}�qv�#:�� #3�ٞg�Zx�m`֭�Aq&�P&�ڎɤ:�<1��k�9�zk¨ۍ痧rnx�Μ|�^��!B��n���Ȯ@|gLP6����A隍�^�Y�c���]�t�q��c K#6��IU�u�F� S	"n����wvl��F�D�7��M�i\F!��b�Gy�nx�q���A=�*,��,g�3���eP�I}Ug�p��]��3������ �qZ�)��>�g�H3;�����z�1+ד�$���g�v���� f�m�� y�U,�Ӻ�3�>ћP� ��ً~ǃm̄ı�@��;��u�GvM�� z�) �A����6;v8��v���چ�z�ܨ�DL�6����}�������-n�t���)%�KB$�z~�x��ا
^�ʎu�����m�6�3vێ�u�ȏany�r�e#��sV�ܝ)�]f��n��C��2�Y����{=ט6 6=�aחFƩnQ�=�"��� }���
5{���!�Kp�/��knl	����N�$&T�||��vf �6=�cmWv �ͩ�h�%:�#S)��7hٻ�ϰl=�sb 0�6�s�N	R�y���"�K�J0
�����Dt��qY��,�d����ڳ�^<�>� ����3 ���Fl�NU`��h�<=��'sT?�?nw��c߶.��;�Ho�"Z!f���Z�D�k��@u_�� >t{v.�lgT>�$��z����"�ۙ�`�q��s!1,dCU��sm��za���P�Uj}:Ӕ޾�fb@ t{�ci�0�;��nv�:+�o��a�S
fIp�̎`c!7n5�t]�R�V�{S�����v���xL�~|������c;f��;��ŀ������ �c:��~a�E~�␲��B ?��_̛��j��!�$�.,�ܘm�~���p�;�Mum�m�  =�E�7�tà>7�7e��{�iu���!Qߔ'K1%��Z'nқl3�m��ʹ�f�LEw�� ���.� �3�|��s���)ĸ��f�����@�ފ� �� ����|���b��%w�,�켵Sc�ws�o��4�<�j�}�8���38\de��bVl�MA:wҗ�rW��7���~�U�㟤� {��m/3Ϲ�uiz;��ঢ$D"ޕ�  ���v�ܔ���ߜf�t�F��۴�mC� ���1,;57O��y�w)P�
N �i�L��B�`.&�e�	�J�[Yz��z�ݜ=z+�W������h�LK׻��s���3�  /{7�1 ���W����tt�b���za��~n�D8�LME��N�n[��w;ֺ���'���l ў�u� #ٟٝ`����K6{\]������e��ծ�!I(d�&Yqi�� �=׋ 9����W#�*똻�g�u��ם٘��Sl'�`�-^x��֦��-poLP ����3  ��z=��ܒ>|�Y�0�^����K���5��Iq��ԅ-���*q��D�s��"_wf,�6=ދ�Ź�g*�&�˼�X�{�-���,�U��ô�C�b�Ž.2w�̕�1Nv:z�71��vp��D����Ð�E��{���Ԕ0��=��\�=!{��q�r��q�`���\/nر���Ų=���;z�A�&6�vz��m�ی��[{.6÷����zey�En�x��n�w["[3����v��b�����õ��p�	��8�����۴��#	�n=�P��g.��ܼ�um]���tssy��\���ٻca�v��@۫��vcL�k��+�(��M�te��:���A`�kmX�`B�n�5N,��*"�L�7��NnaLD��W��q�:����,  [�E�q7ֽ�W��.n
@���u�s�v��DL��{��{�M��A�^C�c�@|�{ۙ�z{��b�+mt�\���t�?fP&����v�|�l=���t�>�{}� ={�����z/��u1
IC%�ą��Lld^��۩�@ ��۶�${}h�[=��Ew�q��ܐ8޿^}�����l'�`�-^�6��i��J	����bU�vf ����-X��OAH)����_*ޭ���栂��YW�Qrm�lM�v��r�F�c	����p�\��	7�>�#D�D��k����y�4�z��-����6�H�W�����@�E��b��C�"%�����s~�w�F�R��?uĔf\�e
�F�����Q�wP�r˝"�j��z�q���U�݌�� rg�F�N�Z{a�[{y�:T�y5d��=�u��ם}�a��������ϼ�g�1��C�=���f�������@�E�S�s��E���σi��	׽��u�]kEncг�9f'���ngL��f2fY�=����uf�1Ș�&@"O�$U:쿒�fg�X2w*�����O11�Lfe=ןy�i��\c1��޾٦bt0�bd��z��+SQ R���# >E���O�k{鯤�~|3�vc1���w�{���%ea�Lf0������1����8�g���?��i}�^ʆ��7��'ޅ��I�D���/0��D��%T��b�Vj޸ɤ�8�z�]��1���,���&'��ϷǴ��η�y��k=��ed���޻��CL�q�3��3�y����3+*3�`�O9��o�N2��l�}W3��{��d�H���&&jA����wH��o7Rf�n�jk;�uu��/[Z�
������-�4�|z�$��bk7�73�Ne�ɆY�>����uf�1�1��ޒ%�����i�z����v6:d}�}�J�r��9�i�2VVJ��C�w��i��f&u�ǯ�T�ĺӝCl�q�'��>�l�C�c2!��<�y�מ)��s�T�;�[=m�C �f0�1��u����1'N3c��L�yϽ�}�vٌ�,�LwϺ��~�;3^�˿O�}u�w>�10��^�XWNf�tu��N8��g>٤��c0�&32ɉ�>����'l�c10a�Ĳ|}���\���lZ���.r��&X�����Mib5-��S��`�d��Z��t�F�+�����rdS��L���YZ.�͜ �ذ�v�mc�+���,\/f��#^��x{��q�'��֥:G^��{���)~у����㻊��s����rٵ�������/z��
�c��l�˕Y�q��a�^fQ܌uA�Y�QN�FP���ke��77gvMɕ��4�u����Ȩ��u������?d~��c`��ԙ�3��fe�mTL݋�T�ޘ�.�꒸�v��=K]%?n�B^��1����.��5N��T��=�rvv�N��Jƻd{֦�����np�#���,g�w<��b���A����>@6��
�u�O
d^M_gftU�AB��ОˑI�/U���wB]���uTPUc�em�߼�~v�#˗1�p){P��-�kMz�N�HB��g-l��o�T��(w����jS7V���]��e6�SwC]q$wSɏg{^{a]�<"Y<p�"���Ts���{;�:��{,���{6_N�J��	��ER���CD	�U-�t�
�\��J�ԡ1	hý�r=�U�Ey�^
_�~�[']v=��F�"*!�CC�͈��'q5E��~�{�7;;�f�[̮÷if�i��w]�� �^��]����G�{��p��W'�S���
K�_&4]y�x:w�������x�[��Hx[�%èc�~�|:�ک6��~����^�^����;Ǻ֎� �C6Y�r����Κ�XB�f�H+T�F��{J�'�&@O��>m�ZQJ�X�Z����c+E(���,b�[,�X
QV��KETEU�UJ�DX���kT��J+�UUjQڨ"����JP�U�m��1�QF���UjQ�(���Z��	�LQ���+YPR�[E��R�Qi����e�*�����E��Qb
e*�,db��[��ʣl�V�KDAU`��)�F+Y�#c����FTmX�X����-A��[JbDVڕ��[A��֪�,�UX�TB�.5����b��Us-j�,`�EA��5�,E-��J��-�DPUUE��*��B��l(�UJR�����b��Qb���Z��b�"1J�*�Y�LDQT�UE[lU��&5r�U#��h��QUV(�TE�R�A���J�Pm�Tl*" �����EX�"��bc�`�5��r��ATV�Z���
�j��UA�Z���(�,S�#�E�r�E�A�1bV��Qjb~�@��Z�݆��J��YY�O���i��C1��YY*yϽ��0�Nٌ37�oe]j�Z�m�zq�����_l>�y��z��k�~g��f2VVε��uf�1��Lq1�9�����;N�1������>�4ϧ���w\�uܚepc1�>���f���f&����u�usYiMu3I���߽�l�C�c1f2W�GKα��ϰ�S����qrt?Q�Lf0�{��i����������߷�N���K�c&8&'��nx'1_���������UM��s�I*&\�ݛ�W�]����y�ssͬ�z[��F���������տzɤ�q���٤��&2�Va�LOyߟo�bNَ	1�������/
>�0�I��r>�w�v⡛�&���q��'���٦c%eC���C��;���ø��f�<��K\.���i'f&�}�a�l�&f2o�.�;��ν=���=���7��i��_�LpLd��}�����d��1�2���}�i�>�A�G��K���~Bf��}���2�VT�u�޻uR��t\ӝCl�pa��9�w�;C�c0C�c1����g�g++Lf0������}�;^�ߺ禙Rwf$�����>�����vc%�1��yϷ<����;
4��f�E'��0���Ϯ�ן:�wm�'��Q����=�>�L{�C�μ>�2��1��c13�y߽CL�%ed��}�u|Պ>����󧎶.s*���Z�'{���Ց�>�0����7��R7�$6��r�^��7j�|_X��aqP�p�7�]��Y��_��N��?Fc1������a�Nٌ0οq��Zr�8��3�{��;g3,�J�������Vc&<뾔��1y�!�}�6��I>��է��v�&&2c3)�����L�,���YH_5b�����'�F�d�0%f������v���bqպ�uV㞹zsmb�۰�ͅیq䎍�����ݾv��2u��~�I�boϾ�}��;f31��3��y߻83l��f0��cs�7�L�:q��G�}�֯�q��ٔ�}s����VK�f2c������O�����z�5�F�Y��z�&�Xk7��i����,�}��^�T��V��D��� �i��#�}��1��{�;��i�N0�c0C�Ȟ��:٦VJʇC1���9�o���Y�Bת��0F�I��;��"��dj�G��f&�~sa��d���2�a�}��i���&2c�Ld���w׻k�|}���{�'�󌘙d�d�{�;�p�9�&2���D=��u�L���V����T�%���5��v^~�3����i�>�g�І3���O��=��f��1��d��=�<��2����G��O���0?��>�s��%3c���w��%�1�9���ᧉ�LL�S�麸��tu��ea�}���x2c0�&2�T������W�{�^򩙿:�ײq��1������t��1���c0Ou�l�*3�c1���}$<}����4�O�_~.y�S�$s?rW���4������n��R'��K�O��F�ۛ��x�؎�ד�߅���<�r�;7=7,���Y�Iu�m�p�7KWZ���T�����Gv2�����l���`��k�gpy=;�@��lv<����P��
YvKY��8ۗs�N��gAk�����J�h�nܸ�c�f�Իn�n�:���B�Ţcv�=j��d���I��m�ݭ�0v1nn��q�4ps��Ȗ1t��ۑx�YIj1�"�ă�ۇ�[����k���U��KSvb�x�DE�����g<&�,t6��i
N��<�]����]�t������պMkF�b��2VT�;�͇��d̳++s�7�]c&8&2c+%"C��->���O�$}����UL.��2}=f�k���i��\c1�5�l�+%eN�����%��e�5�8�'��o���� i��H I��&6�mqf���z��y͟3l��f0��c�^y�F�Y+*N�f2T����|d�wf2\�c&;����{�Iw��{N2b`7��Ub��j!a���O���Dt�&32Ɍ�,���ߟo�i;f8�$I��"x�?WQrf�}��|���f!��bw�<�f�P��C��23�;�����V����}R�NQ�F=f�r8�Mf����6y}�oy�o{7���=2�d�,�ϻ��2�W��Lq1��;����q�1�C��_�t�Jf�4��}���I��<�f�S��L�ͼ��K�)�sM�g�1<�9��gb��f2VTt���(�.�{���}�>�����b��O����&S�������vc%�f2c*y�}�ᧂq���:�|eOq����N�S0.2u�h�\���
'g��cY�u�-�ؼ[d)o�������R=�����=׽�f���&3&Y1��LN���wǴ��I����L�^}�P�8�a��}���M�
�MgeGG�} ��S*�b�f!������}���c�x�]]dִjf.ŝ$�q���m�Q�>�LzO��Z�~�>�\غY��M�Q��]P��f�g^2nI���4�	N�X��mWQh�A���R�A�/C�Ֆb���E+A�Q�������>=�}��ed���Lp13߻����;N�11�LeO<���9�&2��I��IL>��6���v(���F{up=̥��e�5�8�2T׾����P��YP�c1=��tq�g���a���a�=����c��>�wߞ�ed��>q�ɆS����퓳�1��,�LpLO>��C�钧���ީ�h[�k3V�M'��7����#!w�9���Ts5��x��H,{׽��)����<�'H!�?��{�?&��ڼ���zI6wO��%eC�bkλ�}��;f0�w����WNQ�F=f�q�bk���:gL��1�&Y�=ϼ��u,�Ls{����G4�1�=��}�NӸ8Ɍ���=��u�ÖLepc1�u��l�+!ώY#�N!�_��,&�Đ��ػ<�WM5j
��h��N����x�l�ֺ&ۏe��>o��FSX��4Γ��o��}��ٌ�f!��b}���3�8�f0�1��u��ti�'N3{z�c���՞\�}�d��:�{�'gvc%�f2c*{���<N2bfp�;0֜��:Ǫ���=���f��1�e�����>�\��=�J��������I����3�=�P�2VVr!��dOu��l�*��O��@��3��|�ߖ;���f0���ur��j�b�Y�NA�b}���8<g02�dɖcs�7�]K1�$�?�����k}���E;�[I�UA�Q��]_X�Ri`%+�Í�L��y�`��6v��³&�.�˅�O' =ns7ބa�����=�{|���H�}���OS󌘘8Ɍ�e>ן��4�rɌ���������+%eN���/F�)usYiMu3I��~��^�S��B�+�>��@��>�A<���L�3�2&3gz�κ4ʓ��1&8�d�)�}���d���}{���p�׻מ�Y.Y���bu����t�S�{����U@��������F>K����1��Lfe��;����v�]��u��y�u�=xO�v���}�{���%eg"�fA<׾u�L����c1f�{���i����ӽ���x}�<���kp�����e�����v��.�F|��0��u�E]e�7������]e��F?3I>q�����Î��J��YX{�y����d��Lq1�<￾�NӸ8ɉ�g�o�OWγ뙙��������U�����2�$�c�}�|�f�S��L:��z���sM�g�1=�9��ghv�d��s��G5Χ��<��<�qf3++�k�:��*N�f$��1��{�}z}�>��FǤ��g�#?UC�b�z�n}�����iن�\r�W.�'L�<Ϲ��ed���&3�bw�{�=���I��������^o�us^}����w޽���}c1��3�޽�eC�c1���T���|d�+��{���f���г���=�~�Ç�^��b߽�6���c&e�ÙϷ�]K1�Y+�1�'���v��v�&&8��}>���~}�Tn}t�	1�7v�~����;�{j���-r��
3EP��!O�#��'�HN�%�|�E�@��[��wi�1篜��s:�~_�	 I�W��y�=�f�S�a������z5�K���Jk�q�N0�����}���l�JʆFc1=�=�gm�C޽���eל�Vx��1��Y�{٦T�8�I��c&e>�=�l��f2\�c&9�y���&���45�I�6��|&�.d_*X�cӕ���N��'��c:��ZA�.�W\6,��4I����?q������t��GN2c3,���S�;����$��Lf&F�L<ן{�4�'#f2��<����³�z'�ﾶi��1��Fc1��~������]�o�i��Z\4c��i'���^�gL�&Y�����/���f���r�d��Lq1��{���ی��8Ɍɔ�^}��s�Ler	1�󮾱��}�x{מ��*}c10����JhsX�7�i�NF�o��}�q���1��A��K�{��Ι�J��1���\ߓ����������eI��1&8�d�e;�}�l��ٌ�,�LpLL�Ͻ�6�8ɉ�þ4�F�e����q����7�DR�sJCߧEO݇�G�1�I��{�F_s�񓌯pI����3����gI��fc1�'��ζi��^�z�zʞ�o4Wzϰ��}>�9���>�1�g<��kY��]S*�,�N8�K��w�m�2s,�L2�a�y��k��d�ý���C�Gl��Ld��s�}�l��c���d�a��|���l�rɌ�$�cO��Q���� � �)���[��3Vu�of�uc9�3<z�L�֟&<p��3����Z���pg��9���N��5�7����V�2��f���  y����cs�˧K�"��t]H���:�C�tz9l����]k�.Nڞ�kr%���۞ױ�X�5k��Xp��x��*�����n,����0��k�8�v��nyz���#��g��>�<Gl=�(��q�A��$Ū��	��q]m�mۮwY�O'j���=\qȈ�#]v-���,�,����}V�Li��������]��[��WGD]�]!N�mkn��y�n`��Z�kn�'<q�:��ly�ɛo��ߎ��m�j�)���4����Ͻ�l�egb�Cc1/�{���Cc1�D�cu��ti������<��o�.��y�8ɳ)��������d�Y��ʗ��~p0��D���U@��LUUU��L�5��{4��YٖLg.<��w�<��޻��񓌯i1��YS3�>��m�N1���c0Ou��l�*Fc1��� X^�űG��Gf���{��Hݧ6������3I>f%���a���2VVL2�a�}��i����W���IU箎�P�E���|}�#A��Ie��)�yﻆ�ÖLeq&3C�}�[4ʝ1���6��U)��ctޡ�q9��w�ٿG[O��_v3�b�C�ľ��vq�3�c1��YXd�^��F�Rt�1&8�ḑ������|�߳Z�t�YY+�13_u�᷂q�1~�/C��$�?����_���KZ8Ɍ̲c3,����o�q'l��u�Oy���	�v�1�����}Cl�r0�c1f0�=�{4ʇC1��3�`}$=�������|E\}F���8��9xwnu��n-�����)����<ͳ��u:[�vQ"'�b�����|3/lL�m��{����~�����Nf2a�cs�7�]c&8&2c+%L����;N�19�r׻׽{�6�2�����l钲��1��C�}�[4ʝF�L��y�Zr�]f�R��f��17�~���8��YPc���zh��>�gq֫!�����er9�.�$V}�G�?���EUF1�(�ZL,Q�R���-=�����x�����$���/\�6xΙ�1��a���>��uѦT�3`�1�2�y���퓰��d�,�L{����i.�����~p�>��=�|
�4I���iz�&���7����'C���2Ɍ��=��=��Nَ	1��YR�[0���ƹ�zߐ�;N��fD1�������*3�`�f!��O<�Ϸ��;f0����2������3I88�H����T��5Ӷ}������L�Y�9�����Y����Ɍ��3��޻d�;d�VJ��g�y��y�Kw�yM�Rq��&3ַ�[4ʝF�L���]T��5]az���J���s|g���c1�����>���3�iy}�덡Zo��a�`�>��?V|��+%eI��1��y��퓌���1���D���>Gނ>��K�N]���;���8e���6<�ٔѶ�����;lf�8��K1��҆�=~~w����ݬ&�?������5�{٤�8Ɍ�,�̙d���<�|{v�r$�b`���<�Ϻ���0	>����mA�J7@��>~"�qX�+%eC��f!������}��'l�9���.�p\�SX�B�$�ľ�Ϸ�g���}����u&��,#�_��ç�}�L�J��_�LL<��=�NӸ�&&2c3)�y�ۆ��%ex$�c���6dn�dc�s��v(�H��I����!��P2e��5�����W{�W��eghc1�ľ�细��f2O���>��М^Ə���E��O�wY�x��~�w�e��=1������O8F'��%���sm��6���[&��T3y����9%���{�����Q�$��1&��L2�����퓳�1��1Ș��~�6Ι*s�9�����LMUT����Fx��U�(��;�?_M��{����Y�Y17�;�|d�+�Lf2VT��y�CL�q�3�f3u��}$	�����I���I|���v�a����2�����.=f�+*fk޶���L�1��{�k͚�,�&7Y����������Lv&2b`u�y�]�v��11�Lfe>מ}�i�9d�VJ����^l�1�����׏�������ߟ�J�%���9�ѱ���g���6�z����Y�-6K�������n:�m<����|1=߽���؇l�b�C���<��f��1��a�1����^l�1'Q�bL7ѯO�f�y�4��e>���l��f2\,�Lq1=מ}�i��d�Dg;c�NY�$���5���t��R�4}�>��A�9J&���~��A�r��$��I����L���>�g�f3f3�_o͚f!�3�}'�@��_9<G����!V,�>F�c9���.�qL�SX�B�$��1>�y�À�d���e����^l�1��'ޓ>"O�$l��Ue(�W�}\ϼ̬�;d�d�y�<�p�9�&2���y����3��L���cz2�[�3/>�0�I��^�T}f-�ȉ�]�������bu����3l��c%ea�z�~ti����0q�ə��O�~�<�c���Ry�%*,���b�WZ&��W��|�E�q͘��d�[�tQ.�N����5��<К�5�LV�WT�Ј��n�� $���/�c&8��k��ny�����z�]j��kZ�댚N0޺׻4�d����e��;����v�{���]���4����}�4�'c1�!��b}�|�f�Y+*3�$�Ho{��᠍>��9j _�>6�UQ���ed�w�uu`�v�ыm��1Y0Q�=!��֥�;����GF�a�w������35�[�l�&f2a�c��7�]Y����\13�;��d�;q��5��+��c�M)�>��A
_�_�#�A��1��k�:٦T�3�m�ΪSN].��CL�r0��|������� I��'��y����d��|ENf_�3�8�@�*=�<�L��R�{��If��/��d��2Vb]��4�0*S�v�zu][��]^����u�I��YY+,d�߽���N A�� �A�߷������}3xRAI�%Os��٤���+%���}����~���W�e.�ؤ��t���O�G��7j}-|��|�	(3�ٮ�
с[#��w����J�Yby����LN�u���{���$Ă��5���H,:��9����i�W]C�8*{�|�a�8�Y++o<�aY��\��jG}�d@� �OP��t��H)�����)��y��߅�H�����??�髬�܆�S�����������g�#�)�ǥ�珍�P�|�s7=�֥<s��#Z���O�<�F���oo��U�rx�9�Sǟ �e;v�)��v=����s�
�pP%�/{*��ڮ�P���\/ڋ�� �X�w��+���c��`8:{.��+��r�b镚u귏;=ْ�pcGP�a�6(ٱ1I6��"�ZneR�쑼�p��9���^�`)�d3���׸�{�:3�7���\��S��[�6|�ЁPc��a�Ξ�o�<v��Ƕ5o��u���T~���hlX"�V>#=��x��-����f�r���o�}�ۓ���=w��)�T�G$�����[�X����|���N�%��2�DA��*���I���n�=�n�=��>���.[���x�a��O����m��ϴ�<��;s���J��]��G���$ls-����J���3r���w1�彔w�p��{���q��M���;2z������/b���>=<�����OFzdF�E)zꩈ��Ջ���d�Z���^Xs{Xmx�I��묞��Ma�^dDb�����,3�y�{��o��*�тч8.�[B�S���}n��*e�U}�$�L��L�[�g�<{y���f����<�c�YvD\ݺ<}:�ۜ�j|�g���������e8V�:��	a����CE���v�;�R£T�
��X�P��q
��)���^F�4v�52.{9����,
�2K�=t���;MΩm���M6�i�YeLV(�"Z-"�*��UQDV"�e2�+TXň,�*�,r��V1Y�V�D�*U"
�-B��e��\����X"1�԰b#�̦ �
�[R"�X�K��AR�Q*�X�#[[F((��mmX[i��R�K-�Z	���E�J�Am����1+H�A�F��-J¦���*�"�-(����QU(��(��V��QA���$��L����Db�6�jS���FciaW���#EX�U�*��PPDX��,F�E�m�[D-m�)[m�0f2��d��*([Q.a�-�V�*"%*Ո�%��؊��F�1KiP��U�QTTV�EQU�Z��j*1b1�E��X�L�,Qh�mDb�J�R�~����k��5��M��r^M��{g�۝�9y�Ǡ6�m�|�g��˶��v����1�.��'lq�lp���3��C�^�>xi��]������m�i�r�S�;JLWJv�c�\���\���է��q��;���lvW��q�]���:4si��ct�;ٗ����q��l�sN�v,n=nA�v��':v��W]��v��D�vz�r��.53��Y����[ُiR��y8�;lt�.:w����&��q���f����<px͜sp�4;q��u�w;�v���]<k�P�u�7Gh�eq�Cu��]���¹Unn�<dӤ��s����ۗ���s�u�ˁ�]ﯣn|�����D�ctns�����H8˹Ԝ��c��u�"�Fwt�깸�l�]�a�G���7}>��ܽU��m���=���rt���c����6�.E��WzS��6��s�ƍ��狵E����u��|�cq���r��:S�vX���8�c�ʸ9�6� w[]u�s�nk�N%�^q�l=�\st�9�r�S�[����|��d�M��dNB|�lkN:�`,�s7=�@]�C ���/:��5;<����ŷGc�]����iF��/��ox���M���a���;���\�k�5>��a���{0����AS���D�Ś4޻x�.��iM<��1'Ac�\����h��V���os�6E�0���W\��c��o5^=�ɳ�9�����ӊ�\��#����h�˰۱��#93���˦��I]W��gt�lÛuA�vcq�n��g�]���x��^�,�9y�Ϻ��n�{9#�Tx�lmyzR�6%F]a��n\Ӆ��c�Kjb��n[F�/nﳆ��&����m;Vk��/e��+��I�yz���Z<�����{"���9;x��˶�=sې����g����Rn���<n6��sJ۶,���l���@�Xj��E�pv�S�Ƈ����=�9ܯV�D�V�{��sV������z���._����0=l�ŎGr%q�p����H�`\�S�B�����{&��2ƌ��G%4��m�[q��=�OL�l"s�+�4�C�۷0���q�c��խ�K��n��a����N��s�Vy&+��ɫ�9��3�	�����
Z�ۙxv�Nv�<��l$\k��y�ƺ��ۊ��l��e끎�uq�`;$��(�^���m�j��9��bx�շl ��s��O;I�z�0�?�����N+�4����ȓY��٤�+(�Yc%N���vpIĂ°�)�s�:��t¤޹�ϵ�]p8���_l�'���ed���u/�5�%+w��B�ʀ"[�Jڂ��߻㴅����}����w�}������ץ!Z��(}�~{�N,@�<����L�d�Q%A��������N����
ϯlQ�g��,�y몔�.�X^�������a؇X�d��=���ᤂ�Е��9���9F���xQ���A�< D����HV���ᷦK׾S���G!ē�Ʊ��?{)KQ2��� �A�:d�����s��q'�J�XX���#���H�!�o�(��[����v�Y4ʛ����q8�׹�u�jf��B�X`���t=$,�����~�K�< ���7����� D|�R��/����u*AB����b�����Pٌ|n���\�0M���^�ѷf�n�0��U��^U�u������ݱL���͆~P(2���/?���CS���a�$�
�FV���Σ:d�*�P<�}��0:���n�����!�i�<����e!Z��<�6�S�;���au���f/@bt$�o�v(�|����X���[B~��"f��4�X���h��~K����"��{��~���q�gA��32/r�q�P��z���E'Zdх��dm�&E�0!��\�!!?I�y�<�`t�� �����:��t0�*%��}�͚d�eH'��w�����#�,y�0� V���dj�2��W�$���v;H)
Z��<٤��0+X:��|����4}UV�> |F�O�F�
>@2T*J��=�͚a�°�Y���U)�].��CL:aS�u�6�s�']���>I�
�c+���p�'C*J�{���L��R������<��ɭ���#�p��D�����%�x���un.j�6H߷͚Obe���F��� ��-��Ơ;�����Xr��[��t0�*%���6i �t2�Q�<�~�8�@�����^��_��0�"uշ�*p>Y��\s��t�Pu&��˶ntH�����|�S�:R�ݴ�����7$������k��
�����8�S�{�����k�h��@�:���4ΆJ�T*���L:aXS�:�-�㕺Ӗ���r0��}��"Ib�\�����w�;���9ߓ�2����H(*���٤��RKO;�߶9H4�+���g���a�W�+�|~��S"*�I��e^���I�ߞ��AgL��d������a�@��9��=7k��}Nq�OsT��\ܪ�ʠ_n�
'!����{^q�	�rdj�N�{j�r|( YF-����z��3fz-3i�wß�@�u�;�a�aRQ
���9��4�Y:R
y�~� _|�y�.G*&B+%�(&����j���˞g<�!Դ�-���ٮ�!Z��/�w����R�VT�;���L������\O{�@��= �X����XS��|ᢴ�5��/P��<�]{��ID*Aa���72w�����u��bT�����AH)�������R�s���4�����ּ��W��U3o��S � �}(�q̖�3�aw�;�-'ZW��[��{n�%�?��ո����'�Os��f��
��YFJ������N!RV�a}���i ����}���9�}��2t��A� �����'��θe֩�N�.���'á���<" xX����a��{�y��k�B��[)���ހ�p@�P+*{����t�P�*T_�:I��Z�ݼ�G�@>| }�}��q��k-W]C�8¦���v�K��X{{�͝�%P(� T��ɪ�T+����|>��<�϶9H)�{���᧡�R�m~n�2��$��ICIA�����ii�����g�,�%H)���6Hp�+
°��~��4æ%�^}��yܞj�K����&[����BȂ�f=Bdt��}s�:��g9�V�!I�3Ԅ��W��ץ~ü�s\�?��G[���z�kO�[��$�~����������}�5�$G�$�D��%��8�˭����AH[@����5�!�!���p>�j����q�� �կ����+*}����t�R
��X�����������	�u3r`H�6�,Bw-S���=5nY�����7��Aɑ�ןx>zh��`�E�a�aS�u�6C�,��ea���7$��Xy���0:�ι�_xo��7i�w϶9H6�h���<�4�S��r��WF���]g@q8	=�}͚H,���|���ծ�(�,_e���>aXS��u0�0�(�ID�9��4��2�Q���-��:]}����^LN��:� s���u�hӬ˨�T�����l<�����l�T�k��������-��=��@�P+*y����t�R
C��l��V�ϲ�9[�e��p�#
���>�7�k4k��${}���+��#*J�g9�>��MH)
�w��X|�gݕ�V-k��.m��i�S�o����Ffeӕv'BMy��ىЁYY+(�S�;�ݜ�8�}Qb�_EԮ����`>|!Mޯ
> �C�@��w������<2B���6O�B�V��0齱�Vg�i4b��s7�)0_:(UI�fᚎ��bnU�0ƫGU��¢ث�����<ݿ#֍i�洕�p��!�a�nGiv݋<���M����7mX�i���.65{>FI���8�� �u�n[v��ώ]N����ⶓ�0�y�<rG=�JNqg9�s;�&㜛����nJ�s�6˞�ρ��a�:ȕ΃�6�1U�c���ͫ<�[�g� �.�w�g���\���.{���>���9ݾ�3���I��<;���Qq]�b۵&�xu�^kqS�y�n���l���qoa{N��gn�N?�����J�"[�<�#?��i��oٛ��ƪ���8�C����n�3�t�>�(	�5"�����^Dk^B��m�v����H	K�@$�gr@��gM�7-Wn�N����U�DI2j��IǛր$�`l13U>�Ó�"�8��	�Ļ����T	jf+��:u�7�cJ��Q����Y�A ���� K��|�f�R�� ����F�.
L����$�^3�yA>,���;[#bul��j�W�&�[ٽiZm�3:)0x��~�S��{�%̒�Sd8��)����x�n�f�gx���w�m�t"d��])}��|���\"X�c���E��N<漉 �����Z�GI�`靸�F�oZu�SF�P���;Kx�%���W����''�y)��'|��^9<��|�5�6Z�죏M�n�e�6�E���By��N�/R�ye\�Cyq
6'�����&�ɦ��<��%�Ϧ�$(@۬�u5�M��Z�����Rf�]�m=w�JZ!��4�@.�8�O�y�y	p��]����"�$�5R��
Z!�Ie�3�We=ā�Y�d�}�{�nmE�VQ-�EwZ�a7�)dß���m߯ڣ:,��6�{_���qV� I ����j��$v��ʪ����H��I��F���\�`h��4��]n��1�����d��K���'L�6��=�{��Mjͫ$����P�r�T��kA��k���Ւ��3rMT3b	���U]���Wz9���DA%�u���3�M�v����y=ѵ5Pb���&��.�� ��c��V����XLev���F�NB�3Y�UO��"I��� <N�yÄ�Z�r�!8��b6��t�^���{�gZ��w#��ޭʽ�ĂGб͂A#ڧ��M�B�֥$9�d�S6���g�o�f8ֱ E���$�Z�زA �����Ou���(o���mW׎�dp�!�5R�\�	��9�(K�Gd�DUFǌ�͟X�9�d�A������1Yx�����?ݕ�+�;y�;n-�6��-�m/[]Oa�usR�V켴��j�����s�'^����w@�Q��7Z+�ON¼��W��s���S��pP2dDT�$]�iDOwNdݞ����9eAj3b�$����Z�ԫ��v��S~$uoA��w��� ��W�d���*�Z�j��J$�%-Œ	7 ���٪��T8�*d�ٳ����F36����>=��,�	��i Ap��4L�dF��ٹ�p\����Y;�DB�{ܻwrl��]�Ԙ�b+��s,7X�ca ���qn\�a26�^.wo�"��ff��Aɏo��K��#����k�nHs�N꯳ȒYY��*lm<��lT��;�d�vkH|,�o�n�9�o�`N��ۆ2�6=��M;.��r�,Ĝ��M�[t�4B�#�	�B����fH�f+��Z��$�ۜ�Ip���S��qS�	Dq����U�o37��o�p"�,%O��v����A��kI�R8O�cix�YY�d���6*��ޜ'ˑpP30b*j	��v�����t|O��Б�.i�5���k�&��6�\,��q0���C��ʃ��9yQ��-��3:�>$d,�I���,���Փ��}����E�gfj �zfE	�H2��]��1�n�!C�[~&j��G�Λ��EVᙎ���&�dNJ����ҷ*��A�r^Ȼr'U9�'*��� Zx`ᚍͣ6]�&ͭkݨ1L�ox����W�� >t���Xx�S[��]��j�0���A�n��L�j����7;��	���5�C�4�q6+��&z�7�Z�h��=p� �x���ۮ^�N�xWr��ƹd6=��sՎ���>	�&N��=v N��Cճv��y�Ӎ�2T���m;�	G<�λu۷p�u�{c��1��K������7N��%�F�Mv1k�<A;Yz|Qp���xf�ܔ5C[c��Y�q�O+���D/�7#U��w.��)P(&B?��[v����y�(�I	�ٓ�fC��⹬HVtSu�k�� r�9��Һ��7�X:8�|�4@$���>�����=i���gN��^��}��ȡH�������	8Vt�$X�[��E� �^�ͷ��E&��{�I��ô� �I��f���X�g�ă'v��'�͛�3q�2�����Pj��}�ױM�W�˟��&R���I��nv߂Y�3l����;]7�I�Z�������S�F�37UR*��Sx�X�l�z:�S�#tk�1�*�b����L�+�����,q-DB�o|�U-����I��>�{�x�yÅ��YS��6	���+R�$PL�&W�޻���S�F���8?i��׋-nx�n����탟H`���-�f��Z�f �y5�����؟5�}�ܓc�·���a��`(ԊǑ��<����u"�_� F���$�}��7�� |b6�X{P��#�V�}j3�����[�W�������:����nK�NBݛ�Noo$F��\�*P�~,��Wݎ�"'bI�f������ I.t���q�.��ͯ"���(�b��M$^>H�H,��7�M�E��Gk��$���  �:l����'�ر�m8%Ja̹����~�U�.]u�o`�a뮶�pkM;�u�1�����?�yu��8Le��>���@�|�gHw�,�I'�чeȲJ��i�1�4DM"��l�K�H�Ų&���  c����<Hp����Gc�U}��`�W,dn(�5"b�"A�1�$���I(E� #�'��_�r?oL��s�������/�h�׽��z��sn��w�
m�NǼ�;2�T=�&OIzx�쥦�]>����k'����&���=�]֞ď{l�-uU���y�ַz��-��p��:w�r���o;�l�s��j�M�:�k������)��znՔ�V ��gw�yT�]�tWӻ.�'zP2��g��<��u�6���y�I��؛״����܌�വ�p	�4LX7h�q�ŗz9�F%�\�Ō;�e�0��/'�~��O��c�`o��v�=:�؎���EN΀���C�^�t�Ë�znX|����i� ����p��۾Ўuкȴj·T����J�_E���=c�hs���`xx�'z�ҵVoB��������/Y�WI�y�1znq�`�<u%x�~�Wv>���q$z��r�x��('�<6��^��05I���N~L6l��x=�MR'�]���������\��G�]~~p�������s�0�j�)���+/C �/'{�&����7��?LVgaW)ō���Z ���-�'|7wwΞ���O�/4|�~�p��]���o��}Q8��2��[%G��V�ND{��i��y��E��^�a�w�����R�����׶�3n�hz��	�ׄK"*X�)֍�.������-I�-+��Hj�b���+g���p�NDR����۾sǳR��5���U�z�{=B��Bu%(I��n��#F0Z�X��,X��R ���Qm��������F1�B�ʔ�*������TPQ-�`�(Ε,Q�lX
+F*"2�)Z$X8�m+ʴU�P`�cH�k1(�X$��1�Uij�RS�E������1��1����D��*0�UJ�`���V���X��Z«i\�1��Eb"���P�1j�EQA�T*�eUIU*��V��*(5��"5�V[j"�EU)h�,W
�YX(1+VbY�ő���* ������Q,QZ�E�1X(�q�
Eb�Q��U�j�)S�Cy�y������ݝx���/��&�hA��2j�3]r�l�Ƀ��Vx�k�H��gH�H�O�1��4O(6��yUyi[K2䨒Z�����,��F�#5J>ʔ6n�#';�@�6l�wHjon#�5]_*���L|��ݻ<��u书�@�u�k<�r��r�]�2ѻb&FL�/k|�2�nql�7���ҳn� ���68�ޔ��U^*�����3�_7�Z�&!ˏ��&T����D��N�w���v����H#3:��N�}6Iʗ�gm�ܻZ>;fZ"Z"���4F��m=wފm�ў�VRx^^��H�uX$+�lMo��nd!2�����yu(�H�1��� ���l^���>�#b�h-yޫ��21���צ�sۣn��k����冕]�0xe��.��d���R2��w?{�@�����#o*�hA��2j�/}��A�{��X���Ĕ\�As]VA�B}"�"�{����w)�f8{�^܅,�׹3�|%��v[�k�(a�s��u<�n%C�\e<��Ij��?7�]{��|p�sd��ow�-t��GcRgK�@�,���� ��W^��zesCr�	\����� �{�֭4���&�C����s���.>�r���s`A���@�lt桍u�}uĀHv}f�_Z����4DL�P�ck�)r����¹�����|H��� ��ꃘ�1[/N	�&8�E:kqZ��HQ!	��s��^D�_�e�N"&�E��׭y�KK��޾׎���3�9a^�X�A�Ҁs�{�{�4�B�%f�i���K�0z\Y�2M��eDx���W�Ӭ��|����$c��=[l�Ŋ8�O
�Z�.��&��վ��g��ٸ۳�����a\ݰ�M�������}}_V6>��x�c]���Z�βhܻ�L���mr����V��I�� G!��:�籸Z{Rqջ�a�nt<wX�ه6綶k[^�g�\{p�Aq����Sݵ7c�|\��x�pW75��3&�@��Kh^�\6����+�t{+�:`�/BoV��s�棭��8�e�:��&�LW�G}�USB	���W�[Sd���AA-.�3�2`oh\c��l�M�my����1F"�׉�C��f�Y�}F�~f��m� I7�K�� ֳW�s]�md��!�\J��	0��]a�[vA>=�o���IAoU�~$y��K��J��f���)�)A������"��o�X��:�A#awMb{��..����ϒH��6&�D�2(MB@���,�ٰxF�U�w�P�H��IHĶ��@�O��c�ܹU�2��"j�ø��\�<�)�ۙ��urۖ�F�2��۵tOm��Ctp�f�d�TErv�I�]�F�}6�}�:wE�h��78�x�K�����f�Q"T���"�6���Z�sZLf����Z�$P�������.����y�-��#�Ai��z�&q9\�ׯ�g�f����[���DƆ\b����¶o�ȂI/�� �����r쩛Ϝ�8[�'{��ڷ2(	a#���׽}J�`�Y�,�L�`��\mU����K��/�J}6N�\T�ύQ�H��Sp�����uC<Dkʰ	<Wt���Z�Q�뺺a������H��@�J��W�_ �<��߻V]��,�I�]VA
l� �[܂��&�f��=����/i���h<�ƛr�ݺ᭗ˋb�ݪ�-�;g��q����������~�v�ۻ��g�Hս���C8n���
���O�ewM��Bf(ĉ���b�]��fw�u��[�:RI$t,ٰI'V�$	�ͻ�& ���Y�����٧$L��!f.�����o/{n�k9NF�M�GFF[<a����k,l�y՗^o�UsG����^�0��7&��Gw��r���vTq�H�w���#jg�{�c����	�B�6H$[�ֶћ������k}|GW�<�5lcM�.�� �Z�����"�F�f�V��`�q=�~'�ZTD3�TA3�ڂ>$�m�N`plodn&�nH�-m��겐��.DX�[����c�溛v(ݵ0N�������JgQ��i���VV������������w�����n�D�Ax��_n'2�,ӣ�o=q8��#��A>�M@��dP��DD��M�mm
�d�P*)��WsH��}4�M��D?�b���N��W-A,�5U3/�n��$������th���d���7������.ѧQUQ ё�S5�-D�R<�Z��	ufZ �ŵa���ގ��O��}��+�2��xM���WT8�e�i��|��W�1ۢT�ݼ�ڛúva��i�gh�w���5C�[�&	�S�I�+�<7��ǟ}k�UP��LEx�!����H8V}#28�ꨲi�bD�Nbu`�H�O����ٗ���i#�B��̲%�d�'�²�7��*-XŴ�q�tY�=����6�������5Da|g7�"O�x��� ����^<���F�36ǝ�	=���#:����S8R��A�����~��v��A$��-��)��$e9���Fa�ڽu�bj�@3"��/��d�t��`�E�=�lY"�5�Z�$�͡gJ�J�ڮZ�Y
f$�e$�*���<IłHͫ�Y�v�߁$f�����B}޷��?53Y4�s��S1#N!�JAŵ6 y�ϓqS}�,�evU�|H�Z�� ���I��ݚj.��£����.˄���5k�[�͏�l{¦��t��'S�}��3l Ոv�����U��(ը"������|���uoU^�l]�v�|,�\��ۇl���]�\=kmf{��\f7n��獦%v�st��ۓsa��ych�1�m��1����gT���L�g��[m��cX����G���y'f�����n��^q�NwX5�/k�ϰ��%6�nTqd��T��馫c��������L�=������=y��{X���8��L9�6�ۭ�o�.:{k�����\��x�2�[���s݋��������Y�^'�GV��'
Λ'ē����JLA����P�꺚I�ߋ�E&��V���#ƨ�$e�jUM��u�@۫�	:Vt߈>9��aq�!�ޖ�v&�f�<�S�1?L|�X T��I��{�{�[@��ȩ��6.�kk@$���ȰO�v�ڶ��V�"��A
Q%�G��c�Vt���M�]6	 ��m/�@.�e��|���O�72*�j	d)��$���SV�$;λ��	Ѹ�Հhڹ�A ��h |Iw�VΙ{q�jE�����b�۞�����N���,�\��(9��Ӧl��z�����멍�<j~�bڛ$A���D�y�g��t��C+�yQ+�X$��v��ԪI�4f+�����A�qd�Ǐ���gu1+ԏ����
�46��/5���ó	B�n�<yuG��P�� d�r�~�m�
�6�E���Q�[\� ��U�Ӟ����	!�}V	��7���֩�D�Ї"gƤ�$e�u�C�ڰI�#r\�vqm)�H$���^%�uX;�N�Mz��DDA��гi�"-�{"� 	;y�~$����ԳbW9:�Ͼm�W������"��DH��f�>:Wl�:A���Ͱ�2�ԁ$���	%B�[y��/���������s��[[����<xM��ڴ�����Y�*���
|�ϛ幞�ˎ�_Ϯ@��:�d��	������L�/f.�S�aWjz�ՀlN5Bjj	��;�?�_����rq.~�r�0՝VH�	���c�y�Y���U(њ3�l��ud��gH�H!a(CE�Q.��"��Br��T�s7���p=�{��l�6�ל�;�N��W[�F/�=O����7��H��ᝌm�c�g;�s� ?9y|`EwM�}��eD�� �C��n�lmL��	.7�	#z�����H����	�f\�(�i.���6���>��b""�6܋$��yHWPIM���*E�����n͂I5�@(��&����)��nz���p������qsy�lL��h1)��h1_��;��4r=q?����Y#��`�s{����)�͹�����T/s�j&��C�՟X�ȼ5O��7t�O�#cs������1�w죹{R옴U7;��'sGv���M�A��$���MjD��ܻ��I 8���������訚5�p�x(�m6�5�q�I$���$��:�#�X�|�9J."�)Mj��7=�<8˻֩�i��wo��]k�t����K�n�<.�]�Z��D�����ox�N,�Y,��>5$�b�3ݝh�ͿY�*�<�����E�Iv�aA՝@��A���gu�%�7�ڱ{�n���콮h;0n�N����u��V���s?8D���.���c����&3�o�K��$���A��c��e��r��ϸ��[�É�UbE
���"�زqZf�:���ñ�7��O�����t�h��i�{C:Ŵ+�r�LUF(ŀzi�� ���d��g]M_tl�ԍ�5:�*3Ē�my �:�����UQ��"MT��<�G�cј�
1�q[m=��T���7�Q�3`{�C��Bm8��ڼ�LX� Q.I��I��mSkg@����uݹzb�h��Ϋ'Ą��,��uv�d��F���oe�y�u��~=��)��վ�S���f=�+�w{����|�@�n���ƽVS3z��F3ss�ql�{2]	w���iJ{e�=�x�K٫��;2'����57Ǽ��o�ʺ�[<F���eA��!B�\�.��@αb��	/�^�����`:9��i+C�j4�/�}+Anq�w�K��֧�>��{	�諄�;��Q#���Lc�����Z��m�5t��D�/G��t�$�dXwk��@��{���kh�>����ا3'f�^����ʀcد�sz�^N��g��S���4�/o{fA+���=���.j�3׹n��1Wq� ��v}�����%��^�;��t¯*��EFe�$n�6��^�An��{�7.n��^�6�d¯|�k��YҴp�^+�97�@M�T�l�E�9]��J�+m�۫�3j�-Bq����c���k�2)�wm�����5�C�60����۬Q�����|��eڽ�zJ�_Zhj���&�f����
�Sˈ����B��J#��H^.���g�|)���=;w���{��W�2����i>�`ӳ����t������G;_,�<�.n��n2Mq���b��ʴs峊�?]�1�n#;}����5��\q��w����'�]
���ʌ� �I�[�;R�I� <�@���l���
f%�Z{�ķo����s����o�vhd����3^��4�p��3ީ��#�j�ط��j3GK$p0�7���V���{��v��/T��*�m��)�b$�QE�����Z����DF"��L��TCX�Jږ1H�(�E@PU�1H��EPX�b�R"���
��ck ��EU���DTF�E�F�����"Eb�bbX�AQ$UE\�eiA��"1U��"1b�*��*���Jь�EX�V1E�F0DV*��DV1X�"�DE��B�UT���PU��TQ�����eȋZT�F�F,DQBШ��b�D���� �lQ��b�b���N��h��<E�Mn��W[�;rn�DL=oIt�Gy�V���v�r�&#r�&�d��0^c�+�wqvٍ�tvx���-H=�C���`-ϳ�q˭�c���u���6dش����Nc��u�E�<h��`Nl��=s����ݛ�V��Hi��g�{v�I��m�2�z}���]�Wn,3i��wdݴnz��L����ơΑ��l����O^��g�n2��:z3�C�YHG��z�32��lơ5�Cn:\���b�;��f�Wv ���[�~�S�0o�W��q#�ZjoY�1��fiA
kM��V|�N�=�i��p�	|]Q��ruZ�os%�<tvxM�\`4tP)�7j�;th'��H#9S��r��t\�\� ���ݷl<�;���<L�hv�W���G�5r�ۏ
�WL펢v�W�=sНq���&%�6�Uf75��^n����`|�uϵbO��C�7��t���q�]-��;r��=s�a9h��Փ%L��Ʊr�Q:Ѭ�s�'k:�V�L^��z�m]���y�q=N^��gt\�nu��n5�N˩x�g�]��f1,�����cA�1v*�3�ԂC�Ӊ�іX��՜s�(c�
��=&�;9x��.�67Rl�0��R��hc7I��瞽<u��Mmy�Cd���/vs�����. ��v�}����+gv���r���0�O������v�s���i�h��N��S�v��r�CnG�#�-����z�����j&9�gn�[<��ڷ���t[�9���mc�!�zٞDy{spw������b7lk������5����,�t�n7g܆�#��h,��Vni��[˦oN���vvKݞ�b��Y�m�e:uV�-v��8�8ڇAǣ&.�F^s͏9�N���d��۬���S�uںi�b�Ů]��u�=ǵ�mNn�9���Ʊl9P�|r�m�<��`���r�V��{���L��72�s��=�U���Y��3�1"j�uF���[��3ӹ�q�i�=�Q���w�(v�l�'K���BU��'�=����c 񧳲�q�h���$<�v�Hvt�[pb�nz�չ��n�ۀ��g��;/G�3�tv��2U\Bnx���m׸�j�ml uܞ�q�]Kp�{
��N�'�[�s��j���څ����6nCnݮz���Zk۵�5���,�L����3պ:���8:�q�<Qp�g���yX82��\b�+�nS��Ng�cp�]��4���LW�����2:���s�y�]1S�s��PS���,�;R��w1��U`���>$%���Y{{����vI4��0H��Z��J�q<�#�A>;��,���~$�:oco���j#���ME�PB�0]�N�Sm|�gxT�i�ʐM�6�>�Ϋ ���Y�3�1S&`�Q�0O]�$]oa݅D�/.�䧶,�7{�jZ�r�#�b���׽U�j�K��ˀp����B�m����L�wK�Y�s�M⺲A#T�>�|הL�P�n���e*���7Rd������3��qtnm9z6�e֮����ss\&3y��L��{��4@�\��|ײ��4�yf��A$���	��9T����x�Q�,��O0bgƤ�D!���=�����"�U���zLAr���&��ݻ�����nUӴ�{��Of�{�o'X�o� Ě¨��{}����WJ�>m�_$���E�A'y�HZ㘼�7$��W����?L)b�
�=e�K�ݢO��ȉ��
��4�S����}��f�TT���jb�")��5�\�ƫdk������ �^.���s��n�7J���YΔ�13,�\��$�u����9�j�5y40J���N7��x����J�y]|n'+���𽃛���8�m[�a�[�n�ԅ�U��:3�ZK������Z;����6��I�z��Πk6&wխ���Si��{m+k-�T�D�~n������sn���=	E�A ��w�.���º�nt�fq�7�oE��I(lBF[�^Dy�W�O��8'a9�o����M����&�	̯�ɾW�yw�������L�҈�������U��l(�.*MJ��;x#jylq>'��|� H/U�]�SU�F	1s��Ǭ��$��	�؝X��_Bٱ}�U{Eֿ 9J��߯���ۄ��[�vAFtYr�ԇ����"s/�u_�'T��*��i�*NP1S[Yy�%8uv��홏c��Ջ���V���q͠�I�����S2fU�ۦ���$v.�����q��(��.���&�e��ͥY%�ff%�9��b�I�̐�&�X[go9�@$�.��$��d���e�22��K���1k��U�l��wd�3��c�[/yfFe�U&�q�Sk�oEm�
Y*E��<�cc"j��s�dA:�v,Iկ�?�Ll�ߧ7�Z59�ak��hgn��W�T�����tޥ�uK3�f1���r�)��v�r�yם�"�^�d�7
\8iD��0����k������(ԉ&�0b������� �݀��c�|I��B�>�;�d��wY�c��W�w�'��L��z)���y��u��ۣ��[7�T�ݞ4������1���ݑ>����l�6߽��;#�k)�"ns柮;�-b�R��eıi3�38���:cH��v|H$5<�� ����^�|F���neY��F2���D�*�٪��<Iǜ� B(s|�.��o+� �]�`�wq��x&-x�"���M���˶-N���q+vY$])�O��;��"|	 �΢5V�ˮ����S�I��z,l R�P�-������CzK���ywz-����_��[�א ���ev���Nnع�;W5�\�ڬu��&.��kJ���js'i�"���;`��Dy7����v�����߾�:�w�2��`���v��{��ƞ���W7�(�����.�r��0�7�V�H�����:v�K�qy�s�o&�ؗ�]s��4�:�gn��㥘�͚��9�}��ӻ';͝�m�
l<��:��qe�=���m�6�m�g�;�v�$�]��0
�r��Z����zV�g�v�s�]b�L�y��<XG=�l��S�NY�k��#���٨�{��3Y�;��e�l�ڝ���+}��~�ʮa��A�)��$��7�H/3�����
֪�'�4E��n���"%Ē ��")�Yw�k��V�5@�33]�|�:��1���U��wC �q�劈��	���Ob�mZi���T�nfI��y�+�O�<y�W�E����jEQ�RET�Q]�(��ƼH79�|H$��~$�S���1�{J�#F����m*�_Ͳ3$��&�յM5�w� ���ڇ:�]�'�Y|��#3:�F�o��9����8�����)`�"�0��%��&3�V��S���g�}\��������l)d�m�����ۙ���i��x��م�2�Y�.`��^@��:�@ΛfbaD�19�a���o���qQ�}�V�Ѯ}�6�� ��5Yصg/%�4������$�ce�T`���\��w�����)\ �^��Mg៦uX$�R���6:�a���zN��q$�&S�.��j�4���՚�j}��V=�����3:U6��;�n�o�HLDĩ�p���~�^�5ʨm��ʧ�R�X$wq�:֪8k���#I98�_�����FI�R��6��$q�4�¨�!R$��u_��qd�A���W,�Ox�CÕ2D��A�E{;�ƺ��h[dZ�и��.�×�=رj��߇~\������=�~oh(��wk	��#�b�In�~�u�%)��p0��FhI"��m��&�qL�������8�������;l��:�1���ʻ3lG=�%�ޚ��1R`���*=b���=�i��������KN���fs8�-k����ɡYM��S�\��vKxR�y��2��S��sV��|���,G˞�}�g�&gVVˮ ���X$���.{xDњ��ʒ�D�+�w=�^���7
M���sHH/3���{��b�(����p�:<8�D��l!Kvo٘.���.���~~$k���I��A	�uX��߿����;�a?]�=@���q�9�{g���6`9��oZ;Rr�S3c������Ï��O6�Rh��j�qd�|vs�	!�uY����X�S5�d�㽍��a"	1P*���|��E��*�&Ow�'�`�^�;^d׉�+z2�<�Vb�;�p0�"�ВB���A$<�VH7'X�֙z�z8	���� A �Ϋ�'V���(n'��Q��ނ���ҩ�����޵o�y��T�����D�eΥ��W�2g����q�:nN�O*��|� �d�41�ln�����8x�eo����y>�x����E�튥�A�#o�ml�3Q5S �P����R��i��Ⓟ��=��nl,�'�K;t�D����H�=�d�Vra\�1���o�����:��izI�kv6����Yp��n�%֑�n��+�!������T&��.v�� �gX��AJ;��sbmh��BfY�����`�zj!�	�4`Ԛ5)�o�� �e䨉��J��'ė����!)��'����UV�����&*�$�@���	��nŐO�(�_�m�T:�j�z�-	9��o���w߲ދ����ݳ{;rj��b���|E:����`�F�����#�H7֪��szjjD��Lԑ3'e����y�G	����l�"IJ{�� �iVgob7}�.�8Ά*�.�M���k�i��<��YLC5Oq�&�B7#�pJ=�Y+���o�d��N�㟱��ϒhH�v��V��YN��Κ�8T�̗\�A:ܽ�m��Ϥ^��8ݝ�uv��O3��T�7+�]fM����r�s����kQ�z�g��M;6�8g����٩����t�9�\M���ɝ�BT皇�V^[�=��[42�z�kǮ �hx��z�e��<���c�8�����c�oXy.-9l'd:�J�ے�NX�+9�b;tVBqÜ+<�+q�7׍��Z�C�۰֢���w{�D�2eI~q���M��8���7{�^1�(�nk��uՒ	j^���}�1�eB�:�[��:�vn�i�s1�!]�	�v,	;����=B�;2+_��HtL�&��nO�W���L�槔_�����I�+�`��D�eh$�p/�n�h"/D�"d
ffo���U]>D�Vb���Ig����v�O��y�N'��x��� ㍸�Nj;3��L�0�9y|�6&�p�+���Kq~ �������곐�[Y�mw�g�EDT���i�ov-�9�L\�6Ok3;N�,�۳��l>~~��5"MI&jH���7�`���h	�y�V���m�d9��%tX ����.�ڢ$��i�*Hwm�T���]u�.<������P@���4S�`�q�;ݷ�y�����2_�
���{`g�"n,Y�{�vS��j=V���@5��>%gsH�gP�r���e�df�ҧ6E�9��C��	�S�~��`�g]�AN��{3Wt�.�O�����ΕJ�zb�S?2(/�uEt�
���M�_$A �X��'��Os*3�=���ȩ��{Zk��p���& S30�t��WRT�i��|�N}~�HH���D5�V	�#���i%Y���������֡���b����5�B��y.���o�cv3��~���㿻)��������m�ͱD�qOtY�#|`�J�or��ޗ���El�"�0Ӊ������CM��\������f���P�/ăQ^�}ggo��"�13Q�G5�W�k�7�N���wX8�q��Γ�f�zH��Z�/bps����÷u�@S|'@�W
��y�y�B�Q�%=F�Zم<˷�{̞�07
�@b�p�"SK�ڱ��ֈf|�,Wv�ʼ�t�cA5���/~�X���U�|�T�hTf�ߕzw4���/��T����%�e���'���������nl���D�h��Oe݈ջ�r�C..�E-����G����;�PG�zy�z���oK�y.�Z��8��#�0Nf�D�⋷է�1�{��.�^�y y�(�W�$�{@��7tO�!�S��y+G�K/8bkݓ~՞%��Ä��]]�'�ND��K�����Чno8GlcJ�{��K�;A�y���Pg�����_p/.wNE=iZ�ֲ�z�~Y�R������$+P�o�G��iԞ��`��ڠ3Q�I�Lg�E�.�a�п˰�Ά~�*�zHC�g�js)�֕m{VV^̹���P��[tgE��SK�ݻ�$�\�kw����|_oض��f ��G���3-�n��8B_B���{�By�1Vr��8�����-���碙�N�7c�=6x�}�&�f���.�<���$�^KF�4�PF�rks����s1���:��+wx�N�wo.���)h�*�oP�_�V��l�8��A��ZNH����VS�{�ۻ>D�z��Z�
�1N�pv{j�ʕ9�Us�y}�f�I�v!�S�t[g���m�Y�6��Kxh�)�xl|J�mK�f�t^*�򭗘���@c	���TU���h�+b�AUE�5l�#F��j�����UPb�Q�U�Ab"()���T��1Q�+D�Y�U���%F8�EEX�*,f[hQE��������Tb+F�1�TUEV ��
"$A�PTU�3�Tf9hc+D�"��B��iTTR+"�TEA�r)�A�B�Z�U�PG-ED��-���Z��̢�Em*1V(�̴��V($�(�(����UQ��Q��\��Q��-�*媌UX��"���b(���Qq*(�Z����f�".Z�b��DF&Z�����n[F�[�����U�Z"
�
ڕ�E̔bn�]o�/\�6(�:��j�o����73.b\S6k�	��u]�����A�8���>9��uE�[����#!>�'Q4^I�^���0�jZ����i	�G5���\a
�ޛ'Ć��,H5� ��C�`L����jU�n����K�g�����2[vk��L��K��O�a�ɧ)��|��mK$Q�,�k�H�Њ޺E��$��E�F�=3��L���H����q��T0�.�I-K�Foo ��{3�nvO��Lgͮ�z�Ċ�N% <O�M��}�i�&.�e���f78AT�$A���.{����!�ʒ��.R8��USi���m�{�� �:^�	v�r��������N����/�dr���"p(�"�ek��d�5ժ�'~�����n��᣺��:�ВVCDf��P���?g=����F�u�7@����o�:���$Vt�w1^�Ohv�:���ח�p������Ԧ�[W&�c�҆[�=O���;�=�n��^��tF���IN�B��}��ނ!L�LȠ�Z^�SL��h|H��#N�앑ے/Ă��$V��f`T�L�C;]��,�=r��[��@ ���D�gM�H��V���2%�I�����߁ZNE���\�u�YY�(��2+�c֮l	/wz����#zњ�MI	����RXګ�|2�B�R�&g�$I$8Y�)�/�;�ӗ�c��h�x/�jwj�M�&j"b�f�TI�w~�iY�`�����cO.�O�y��t,sd�FB}6���وy����/w���:9���?�*�3F���mQ�:g<2�u�S��������fC�vǏy٫R��ɋ�ŲNSܾ"2ws{��v��n0�u�p+�^2�ɫg�N=�.8�Ü�	u�7\7n�Gb��R�*��"o,љL�$m��V�	�q����Fp�A=˅�^�r<�7[<�Ɨ�M[�^og����Q��	�p.j츹���㞤��6m��	�WL��81���]8Q �ڷp�qݺu۹���v�#�io�����y�kc�M%��U����f-m��=79��Tq'Z�m\k�Q��(�������|HBs2ɒ?|�Um�>w�J[Oл�sۀf�cș�=@ |H�Y�d�"h�12*�SU"a'
�l�*�5 �\�����6	�'�	�߉2�D������&��ڿ(-Zi���t�
��  ���p�gM�l�c36?;͊m��
��^��(j%Kw�r�r��Z����D���͒	7;�[㧲3���<Նv=��6KޥF$�&	M��Tci6�s�vsY��Xg�E�@��S`�|-�	�����k����ߧ�"]���v��n#]nq[�ν�=��:�yn�](K�/'Y������[���I��͐�Α`�3s�/�����ܮ��V��i�/v)�F7�-�w�u�_�0s���WgK����7���ˇ�|b
��-�ӻ�91l+H���͌d-U��}� ��u)�.5B�R���Ț�CE���GmV�\O�FBޛ�㛏����L���NvoČDҍ��^���0��t�$��iA�#�7z�E�7W8IEv���nwZX&@�3j�(��3B^��r��@�.�lH��iK��:�*�B��R�$3!�͂�t@�4	B�@�r� Ief߅'7��*���ރǯf�$x�grHt�3.�N���mr�`6��f!�	�$G�.L\�:���y�lu�[m�<��J�o�ߟ��G��.�&:c9H�HsH�	p��X]�̗��%��8]�,���D]�&hĞ�ow����g�����\�e?ڈ �7��@O�,�3���j'�z�"�t�����!8��+�t�ݦ��u�� �R�o���Эh���E3�0Օ�'{U��Έy<�g[�j!���=�l�F�W�������y^��|w��ˇ_l������ %���M�y�I��ۺD
%˙�Az�z!�ɋ7��($5ͤ$8Y�~$����"��t�j֤	Ʉ,jbUT�G��>#
�1�γ����	�\�$@�Y�d�6�VfP�|����P�R�k*a��A.!�" �i��a�I�n�6W;��9��ϲ6����w���(����䏉�ef�A	��:�z�]E^�ʥ� I�Y�d���EG�������o)�AzL�QX��n���|H�Y�/��.�HG>1__%��oi��k�Tb�F�� �YY�,�v7��J!E]C��|	,�ٰH$i{�N�7Zԓ'!E&l�������q�c�H6w�߉$8[�d������>ۦG��w6�ài�ѡk��T+�)�\`�l�Q[[�N�F�GW.���RvJ���E�ܻ�QUU5c_M>�����-��&���C�7*&����USUB"��r�$��9�%�W=��{$�m���;�6O���ו��Nqa��l;	�pɈj`d6
C,��%���vp�,-r�j�;t�P�Ũ��ߘ����LA���ۿQ �Α`sq��i���՜����f�>:{6F�p*S)�J�
����m��$w���{�NWp�A dv9�A7;� u�D)8S�͙�@�U��x��������צ�$���'�i��83c�[JG=�"�'�%����^���m��a���Ġ��R	Nc�d�56��"�?lF�d�/�"z��X(���L�I�#�֭?��Υ=s0�A��F�͂Hk���$��#��2�K�N�Mn��Ӕ7���T|��x�&���+��~�T��]�Jz}˯�q�9a>w�����+��{���>��T���}E�w��BfX���L���1���5E�2H�n�#�h�O��7:��&X����Rq	��y3kn����1Յkq���W"��[��;!�^x�z\�s{'X.��ٻR{ۀ�c�l�:�X�n���gjc=�9_)ڼa/������m��ێ7�=u�ֻ]ɮI���v5k��^�W�c��4淘��ṭB�M�j����)�l���1nmt���p�<M��Aᴴ�A!��������ꢦ�E�U���I��x�O�^t�2��*Njrl�)`�Iż�,�� ���� �,�������:�d�d�$�o�$If�H�	��;q�6�qML�$L5#T�c�~���Y��Zm&���Nn� $����b���n�b��Z=�+O�=hU}����z}m� �f�"	�^l�$�gI��p#�8w8^�%�<A���f�I�LUQ�N�Q��t�56{;�B!�4�jo����o�gB��)�[����D����]�_c�n�.�s֓W�<mh9����� :��Z�b nfB&#�^�5���
>$���~7����O줗� �+=��N�{I��q}o�$;�/C��(�O�k�UP�SW:j���	uR��%��W�u
��*��fHܞ���h���:����P�{�n�b]�� ��'b�͂I���n^��diM�r�����S8��'Dnۻ>$��ٰ ²�'��d֝Y$���nS�D��EI^��/�)�MH*��3yU�A#��f��l��>���'�=9r�Wi����|v.c�����AdC&b��0)m�Y �27�$�|��Y�r�Y�WU�[�Cuq�;��ūj۲�ڭ�v5i�iS��nƙs$K3��]1,�?A32B�h��T�<s:E�|��X��v1�1��L�l��!�8�.� ������źŦ�ݿYay�d�ou���I1������/�"����Z��gM�@$�>v�4ʉ�RfkwT"����-�ݔ�%H�R/jT��\�wm��e��,�l��{�	}���{{l�i�ƍ��C2ܬ=wĄ�n�S���\tܵVI>��r/Āou��&#-���&e	�^�tB�{J[o�H6i��>&���$x��uc�˹;��^|�sd_��q����"d���=�"	,�۩u[�.��O�-��$�v����R��C���?�s('I�Ə��v9�9�g��n;;����YWv��ջrn{qm�2�7;�d���%�������f��Iص�`�w7����Tc6E�E��^Q��rh�񚨨�k�j�m�ّ�jީ¦�|H$���^Cb�M�o���>n�r<s173$D���s�L��D���-r��I ��k�v*�+��Ք�D1������C7͹�*x��4�$�b�M�v;:wb�JZ�n��3�T����br3�������sELR�f2i�U�<&/1۱�t���m��;0�J����S����(�������Qɿ��vU�Z�[m��UP�F���P ���uWfyN��4wשI�Ů��/:F�vl4cVAQ�9֗��l͑��]n7V�䎁���3+�=�Ϧ�"`	���RL�D5#^{�i�ͭ�$�/:l����j�	�~/uݫM7�{�k'v�I>q)���Njl�!�M�ޮx�>�]6I;�6	��7�1�g��י�Dn�3F��d���s��^gBR̮G���tf�e���/�M5�s��mQ�G�f"$�DL���M��ڦg��14��	��{�7�{ʣ�>%E����_��L0���΅_&���ۻ���2Kjl�!7>�dvt�$����=�xS�+��Įx�Z[oS�0SoZі1������S����<7 ��dz����6jˎ5�UVJ
T&n�bj��Ce��a	x�Dz�x�,�W��Q���RC�Vm���3R_n���U�
��4L�,@�5��f��i��������r�M���[�6� S����z�޼N�w�Ԗj��g��D�P2w�u*�Şʹ���}��ni��ƜK��C0�iOh��y�ڽ�4�`�O?A�	58,���������MD���N�ٮ����ڷ.44'�p�r&Xtov��NS�2D[��r��J���!�G �҇��u���t�A�F;�%�sL)�|&�0}�\I���m���t0�3I�0��<1��N~��so4���A�7�"^�8y44��qNO/c*˵�����1ݓ��7��H8œ��Oa��W/h�y� G��t�X�p�3���ٱ���B�!�%�����4.z%x�"��3Ϛѯ�K�ׁ>�x���֯�xh�,�f+'BT�bٌ6}Me=��6��(q�O�׫�<�̄�3|����D�����7=̰��쎪<��Q���.Ǆ���|��Hw[�qIG�0�C�x�*��^�$�Y���:<D�0�,��,X�J��Q��o�}ӽ{A쪬�Dhc���/ʏ����مs;�g
,IH`ӗ�kέ��}�h�0	��]�V�adO;�%��Mo?%�}V�p�Tx=�����٘��d��+�s�M^F�����ג�����i�n�aw������^�C�ň\��Um(�X11
���*�D�Q�r�#Qe\J[��q*��U"ZW���UE(6�����h�1�)�h�Dr�iV�hڦ5E��-e�b�
���DZ�c)e�A�����Z���%eJ%�T`��H(��Q�TVU�R1UUX�U-(��S�DQ��̢�j��5QB�Թa[��TX��EUE��UAb332�F"�ب�EdkVF+
ܵ��L`�V�br�*�.fAQ�(��*�"��(���FceKm���AV[-B��
R�6�J�k��(�`�J4q���+�Q\K-(�Q��E���ZU��F�TQD��ª��U8�~_�p;t�Ҽ����":�2��ղ�ݧn��y�ܽ�t��8�7�gg��=w!.!q�9V���`*(�vnS�����n�m!s�XMTˮ�#�ή�ڜK���:���cmk���wiU��=�D�q�Qz��`�h����t�9C�l��b��l"����8׷W�f�Dd�XU.��ݹ�(�Yӻ{s��ي�U�d9���8�0���N����g��臷ch����;�t�PW�&�z,�:.x��on�ݐH�vc�]]�z�e*mSn�9ANr��'eLi���=b,�k����	ӷYz�m��ӧ��Y8<�Ɯ��[�&ev�W��OT;��9�ұ�ܐ�Zs��9Z�{<����ΜZ\���w����9F��V��=v㶈��r�ܾx2
��7n���ڸ��Ζ��wL�\b5����0��Ŗ{\��7\\u��^G݃�Na�:�s��wN-�ycr����w
�zT{Qɷ#���v\{ll����7'=�nz�8�v�Jݹ�nۚ�˅q� ���:�;׭���ۻn3ƻ�aύ�W]�'q���nLZ�,g��,���z��<��˨uE.�R{m�n��E�m�{c[p�GGpuœd��Ӯ�x�J6B[�mu#�Ÿ�k<�mK�S6a�88�ѷ=��]�U�d]�Ge���sۅ�0�ޠ����n��.B�x��ε۶�]F���-���p��&G����z�u�u�_<������v�pr٧c�Wv9�8�jݱ���ŇԧN�鶭���h}�[����^�v[y:��r�v����tsSo/��u����.����\���۲�p1nν��<[6�Ϯ�ͪ��1j�
�x�ȃ�捍�^�]��gd;*��nsSu솓uƍ�<�n=����n^�7Y��{<�1���7[�qѼ8o]�۶0n�m[��Y�q�|��q\s;0�L8�������Ǜ(8�[�iU�ƺ4�]Y��Չ�����vGvN�%�m˷g����ɑ�χl��lWk�/��Ze�x�i󎋺�ķd�M�C���G+��i�jm�=n�=���^�k��2s8�rY�2!ε˕0u��v�z�E�u�t+ԗ��m�R�'>�&���yt)�q���k�s��l(�3��nN��N��__GOH#�t��0�N�uI�0�A�d.dM�]7�:�<��ntn�j��2p�Me��pW��ק�
�������F���[�Gă��͒	���ӂ6*=�E̵�V�f3e�G�s���Z ƾԃ�2z����O]�O�3:l�O��|� ���K[��d��Ro'ި�c��Ja�F$� �����M��}SF��u���3��H$Z�"#{�è�U�5FBFj��2!���'v.�p�&��M�A �j��$�����X0еM�n4�����f"&
O�5���~y}Jr|�=��\1�s~$�qv���.��9���|z9m\�n���0�0�˄���5�x��ܼe�xE��F�n.�[�:��ZK�����@�,�a}���|�m<��i��/���uyךA�^�����}�ȃX
D�!3(N���u)iպn��+�r�x%^�o���O����1I�	5��w�R�s��-�ۻQ�H�W?o�x݃�C����)鹃�(Wp3V�7w�S���ٹ�A ��4�.���.;�����D�/��m,�8�$L����H��j�$��-�D��3HqFr�X�<O�ջ��r1t�#+��EO��1D��Es��n��pG5�A ��l�@ޞ�Yڧ��3�<I��iN��MW�h�;yD�݋���ۊ� �9��^$���X�\�őYB�g��?�?��ۂ�k��ڥ���c���qa��}c����[�tnVݔ�lW����70���8�SV�.��5�lY�5Z��G�I�k��$�db�"�I�0e�.���Sny��x9F����:+�P>'#� ��{b�B���d��߇L$n��v�E^_p��(O�.h��7�a�
2��:�xq��v��-=���y]�����fQ�"�yõQȼX�LSP�$^����t�-axi�� lb�	�=�emA�U��*�u���)Oc�\�wr��	'�%�z����J�N�vr���o��\oE&�}�*\!ħ����)4�^�4���mF��H5W�d��s����>AS���!a���2�Uy�1�t�����y|�[GV����c[�Z����g�.�,�	&���$�8���߆���3d�H'w%�|�-ٵZ&6�A$�d�`�k�b�̑�؞�B��ypsr]Պ$����,�A��������;�������7�0��&U��V,IǛ�A���]Wٯ+mNT� �y�,�|ws�Ѷ
F	335T ����E�b)���A$��D���3��tP��nz��wu�\e7���GB<i�U\�{��mj�|���(.ɪar'u�o�T�����}6l)��m�7	��O��c2�b�6Fu��PZ����D� y�a��fخ��{Wd�&%���V,�O�nw/$�oLΏ���%�fQ�r�)�r�o�a��+r��\d\s���T&7�����𛧑��R�'�8��Q)�)�8��\�O}�����6��1�ܓ�������	�#�^kH�{�LK�5>�5UR��j��5%�i���\��	���Hu�tSo��cBy�E�mW�X.��SQS5g��D��gX�8���;;��LDs�"K�ް�Y��qbGL��F*LE���M	={P�]�P	3:E��O��B�y��$�^$7���$�33UB�;n�A՝B����YI�-�{��O���s`���{������ͣ����y	�1=X�F�0��^�S������w\:7}�=��3B�&�$�[�����k���{�w��s.�\鍱®��mU��:8۶���k��-�H��;���s��ӫ�l/%��ػ��9Ϣ�n�Ж�y�t��6�q�n�퇃��m�C�'g.n�p�!ȝ-N��w��k��Y{;F�lhI��EN�\�)�g�ݷ0�����Y�,�	�����]�g�w���{�}wЩ�6���a�pr���1n8[]r�]�Ar۶﫟�o��3��� �������mvt]Eu٪y��C��8��F�������Zv��PB���H�C9�>�O�Y�6�9u��Y}>���]�M�3:)���*\Gf��4�Y�5�����ʬ���f.��FfȲF�����!vc�|f+y��k�H�������MM�Ρd��-�+�y�3�	,�t�$j�a���[2����!I�Oe�_{�T�CJ�Hŝb�	 �����Em�F�R��~m�E'��.��I#
��nŒF<�@!f�7�����h���$rޱ`A���*��w��ǔ���g������ v��X��[��g5���g7\�,A2�9&I��]��l���B}���ۢF��I ���H�S�z��ot�V�S�"�ջb�'���ɩ��$D�PB@�y�w'��F��3B�T�r�8p��|.�v����Yi�r��t�6Cw�\�i1��f��
fl)NL��v�S�\�طN-�7Gwz� �Y�,	;��� ��V���J�fuޝk�&��5&1&u��9�A>:�fr��U�d���B� ����\v�	�LL@�����b�e���Z�V5CA>$���%�A.3:bFL9�ە��RM�\Ï,��s0HR}.� K9�b���Gb�ٗ<�����nŒ	9�Z^g3��YJ�EӒfj�۪��q���l�s<���7Fӳ]�GOV0��2@H�qk��P�@�� V\�W6�G;w���%�Λ�`��2�rj�o(0A �{�"๛	135T ,���1�D.���N�R���� �B�֐-����~�G����z���{	���DI$4�y|9�tA&�o#�</r1�f��Jr ^��s��]�{�,zA�|e۫��dul1uBt�sO���\��+����'�`~�.؞%�㸌�ó�ϸ��w��3��O�3�tdj	C���J}�o)n�"g���7��A:�yI�Ff���N.�#%�D��#\��5ό�È��&��`�L�����ʽb#�t�/V�c�>��R� ��ٲ'\l�'�Kw�@��-Df*����y�ˤ�v�D����6�x1ը�X ��^�[������I�@Թ�$���m�y�R�b��g"�8������{� N��E7�wKeCaS0w��O:m?9]4RWL�U�$�:36o�����'��nt���=Z��/�N�  OMEq���I�Ӧ�&�Lk�g-\er^$23:l�1uq�@W�3�����EA	x�O�����x�*#K� �6���Z��~$�w{yƛ�O�]�j*i���bBcC�;,1v��z5m���Q�:}�9���3b;�������o�kݰh7�{V�i8�b�����i���n~�F�8!Ƕ)�l�^���֫d�[�%�
��I�,�"�>;�yys=뽤S�ͣzj��k��5�X6�v��S�D^ͺ|5���ix��ݸ��������	�p�& {��5�]�鿉��{ּޫ�2fMc�{����Rz����Q����.z�y�aH+��˩�uB���^c�`�H;��~�n�]�
�������Lp53��αd�N=�^�w��WE��&��>=���H;�yy��7D�b*j�@6F��F�E�>�&�]��{��$��Γ#B���2���]�$r�b̽q8f��I$Thi��K9�Z�y��\�:O��X�H�u� AÙ�g@�z���s|�C��.�TA73{�E�D�$����+"�\P��z�u�=8�{���$�(���mLy'<��Y5g\<=f9@�\�n�ۍ;�C�s6/I�^�%���,sV߷�n�-We�������j�緳�T��`�.sgc]Q瓤�cl�"�y��72�)�\:�����|`��-��nCWJ�p���1�pv�z�o,�r�v��xܝ�Y[yÃ4z0mg����Z��oDt��N��j[��!<mk�'c�J�������͡-���u��eҝm�z���K��ù��Թ]��t&�dۋnpfh�,�I5�4H�f$˥C�A{�����3�h�\m�w�����>�|fe���&��`�`�W�'e	9��r����$���H	�FgM�S�=�������?L@|+Z/�#�;��%}�e� �>:s:l���5�C�jJm�{�j�a��I��wK�Bc��%I�m�kJ��fm�D����d�=�ޥҍ�g�+H��g:մ�O(�m��ۇ�^Y��v������x+����@�63�$�3���=�EN���
��UF���f9n `�C�%p᭮c��s�������O;=ۇ��k�W���|ʽ��#&/� P������^쁯z�OU��<�j@�63�%P훒k�h�@�I�]t͂L�ٽ�Vi�r�+��7^99� jVN�W����d2��B'���z��=�wҜu@�%gn��#��}�9��w����,����2]��դYl�1Q�4��5��ɖb�L������MX�yӦ� ����#'jŧ���fl�$�}Zo�b�,�צ���5~.z�+q���[�W�`�
{�����c1�hu���J�6	���� ��"��AHu=�d��w���I�;�Nr���E�]���ݛB�O�u�$������歯,��d�H���u�%�iL�Z祬ݭ�A��q\sd]�Ί���p�D�"*j�@=�-͂AכB�H$�n��-�o^����G^͒H�b�"^38j���I�$$4�yuN�ɑ�*�+6�D���_���ް�E�s��:�Μ����$P&f/��X�I>/{Z� �a!��8	�����piq+��ͅ >Ё�'��0�lym���Hבmf�yiކE�+�}�g��#]�oR)�������.j~X����<f�]{��d����&�s�X�w��P��ڪ�NzY�5��8sF?p���rշ��˦*.!�v9�D�&т�_���S3s��R>3/sɓ&�Y5��P9��sy����Z�R6��J�ų4�e������f�V�%�U�ÙWN���&�,�:V���ݫ���ݹ�]��s����:X�Ÿn��?�"���>�zk���!�٬r�P�3��w���J����5�a��c�[��pŸ�;�r�_*b���ӎ_.~�Q�FWm}��9"�sf�/1�<�r�d=|�>�w��!='7q�ƃ1�۾�
$��)� �J;|G#4)�'�"V=6n-k(M�����I�h���Y�j�đ@��B����֕M�6�Gjj1	��E/-��=��2����<|�Rr}�j��uo5/v7��%��q����r���{4h6�%FV��Ȫ��z���<���Ŵ�
�^MdM�ۯ�T��/5Q�{�2 ���ޮw��g�nX�=�%�=�>��4A�=)o=>�G�d�O��MҼ��Z�Y!�2!��!�[V�A�.��w5t.�={3U��~�34�����E�ԋ��d-��8Y����U&��E�ٿ�Z��Cs
��7���7��6uZ#2Q�ɵx�Y�wF
��;o�V��ۉ��l�!��H�a��ê:�Ib*+�Qƣ�m�h�X�����ie���ډm2�U`���V��kR�YDm��9�����b�ڔJ���2�q�W�p����(�Q5b*2�iJ6�lERб�D�hP����J���r�ʔ��[F[F\q�`�Z�s0UT3)U\X����8��T�mJ	�e�L��-��q��"�h�R�DJ�-�ETD�e����֭m�PW
(��D"��kQ`�iQ���ԥ��%�(�e�H��R9j6���\���J�R��m������h��Am��e�-im��إQ(R����J�ZTZ0UVږ�jV�Q��m���E�JEF�A*����DV�[
�4��������#KYj�B�k[J�J-��F�J��-Q��j�J�iV�0�ciQ���
*��QKh5m-�lUYE�kk-�Uj%�֪*,��ke)m(�)km��ѣR�h�4mЪ�[FگYw�OC�s��Gw��DV�3&Y��"b��
C�5����$�S�Y$��i	�0e�zP�d��ת��fE7�b~�I#���8�˫ ���Ci��<��݈��>[5\�����7cl^#8�A��ޜW��{��s�d�[�r��d�ݱ�^�=���8t���Tkn�s��t�~�g�ˁ�%/����Ս���5`|fq�~��Օ�\�H�w{fՁtb���A13N�q\T��^}H���l��>38�Hf�����_�'�N2I��!�}{�V|fiR ��	���l�|�3��X�>��R�o��k�h�@��(���ݺx�����tl@��wV �#4� 6s�[P,s�3����'m�;�C��|�ٵ�L�V�嵽�����М�!�(U����:���o�k��ɜ��lG��?U�E�����gd݅n�qA05̃��C����@ ܌�՞;ǫ�گ �g�m���"�Hf�qvN�^�[<�y�7�̘dȜ�"A�duO<�s����qaz�n�+%�u�W-��-�4�b�|���\��*Z�G&G���n�s3��@tga"29��.��@w��Ռ�2u� >^W5�'���6�8�h=����},�۫l�2y� 3g8��`Y;��>��>���l�"�M��!;�y��  {�<_�s�=G�ygOOr��'�R�tg`��N2I��H�D����ިȾ�.�>��o�����>@�lg$���p������ ��gWĜi{a�s�MJn"��+�p�`���_E�D��p ��Q�?tg�`��M6׸��n�"�/˶���oOD[����W��S;*��l�p��61s���=�k3��K5.�/>���BǼ�fj�Rܩ�;AP��n��E��kd=��nE�mt��E�3ɑ�������B�m�'m�y�%���9|#��:Ʀ$/^��msq���뎷}p\��G=�D�j�ٳ]�`�&��t틃�����٫�l�\�ۑ��hyfњ\�Wm��S{\- �mյ[��\z��gm� �J���] �v��\�Ws�]g�ܓ��˴6����燩���Ж����g��%�O8�j�3����tu�[TOp'']nb&���p
	�!��C�YR6͟� 2N���'�����S_���"� �7'<S�
y���~�$�J� q՗V$�A�ƚ��Y�CπvsK����M�c
t�r����o�y\ָ��P5$�e�6�8� =��j��v����,��q�L^���j�~�tڰ��1i��bIbwh����ˇ{0݇\u�` o�n�6x��2��=�[�������8�&&b�}{��X�fi<�D�����=X�U��]� {�7c>�g�[�:�f2Q���OY'�`��b��(ku�G �^D�%��(Q�ƩN�oC���2���FG"�w�߻�ub�<Fq�tߦ�ҾMN�iXϐ�{�����qL&H\(�-E��=��9dev��y�"�Jۭ���{)���,��Kj�G��t�]��cbkd�aZ����nb(�f�l�w�Oz_B6m�Y㚞�o��� ��7��gI ����Ò[g]zz�t�a��*\�'��\�9.-����y��H$ê��QNt��v 7����|�^#8��+���CNe1�h�����zc�� ���MZ��"��ޥ�����܂�s�A[����1m�����'vk�┍�=��+Vu'�]��LC��mw��4��) 3{֭X�W5s�Uw��5���P}>�&�g�!B��:|���b��B���]i���t�썷������D��3������V�k3J�F�oz���;n��H�6>�ɻg��"��y��9�Ķ�6EŢ��ի ���37bB�S�[U4݁�f�H���Z��`V�]�gu�m+;�D8��e�\Y6�R�nw�]�6���\��F'�Kh��)�e����	$M�t�+!�٩ɄA!"�"�Q�%�~�ZQ��y	�㸡�h�����y$�E-�8q����X5u��@�3�P��J����'���9.,Og�K�F^�t x�*�;���>f���n�v<\�����K��y�8әLeٵ޻����$z_����}�dGޒo��J|�O"�M ����������mY�uu2�i_�'�����c$�ˁ2b6�pIp1�8�{.���:�7k� �\cE��������0L̸N�b�������Ս����W�l�P����ś��&��w�W��Q���� ��%KWh�u���e�s]���ߨ ��z��6��n� �s�H����]��k��݂���Kr�d\�Eum�V��;o� �l�oM��X��N��o��V0���6��JwϢL&��^���gL����8��(6IQT�> n{�� ��'j���3x���C�*��Y"%�w�����q��������{d2��[���ǟ�G���Du��v����=�T���r �ݻ�K�-�%Kj�9./�'���>38��s1��>����^]�����M�k�g@T��S�[�ʊ*J��ġ9�$��i�q ��f����eE�Z���hِ��@uݗ_]����.C�m\�ǫ6�+ >�~��k����lGz��q�Dneݫf��V
��d[m��f)ݣ�+��	�Dت:;�S�������w�6�g_�]Gm2	^q=~�S��#	&��J�����]Y�6��)P j�ݏn�0�Yyl��� {;f�m���M��%9�ĹL��+��_��Yt]z�m�qw֦�'��M DF����yu��I:"g��E6\()8��Yp�m���Wg`΃��@�3"��Oc8�ۥ���m������B4��ܜ����G_^L����8FQ��2n�m��3��F�����d9�yI�U��"�u��)SVh���BX�a��P1���|���6��ٽwm��>\�=6x�.��m��;�3��4�Ÿk�K���p�rs]Yy��P�16�n�tm���2��={</+��[<�%.��S�N2�b��3ޗ8Ӹ���X⻥+$��Í۶�^9�rk=�&�e�WC���[�61۰��7�v������[+C�.֧nj�����u�ps�ţ,����˵�z��KٻX�V:���Jv;8���4��H0Z�XW���na����������w� �e����3�T	 �g]�V��X(��Q�vu�_�0њM 1\�8��M̧�6���D�}�S�Dnl� ,3���${s��gĿ��~B�Rɭ��\ � �=�Gc�Bح*��� l�]�ʩꙘ� >�g@�gU�`���&�5/��s���n��4@��� �λ��ޏG�s�Y���� >yD��N����&�.{j����;no��l�WS�&�D���I�w@ f��7����<�0�G�|Ģrx�0���4��ڛ�LWlθ	��k�W&�8-��������<�Kq$(%L�a��9P ��:�X�ћ�v����#އ�&�@��v��i�I��	�6=����d�ed�Q��\X����ζ�.��1��+dU�uZ9я��ByMtk':��"���Eւ�E�os6��Q-f�o�=�E����ʃd�vg�������/Ū��"�QD��}j湲c�����o�� L�ZS`~cu����gU�c�f�_�Qx2-��˙��ub�W���2P:���>@ >��ػ ��q�ݩ��}�|׹w���s�2d�0�D�v��ι��Zf��5U��R�T�Q����FwE�c�3�o��G����ܫmf(d:s3(p�Uuۏ=G&���y+�Ԝ�׶�C9�Onq�����ƧA3"�+�wN���M� �gH&<�Tu��iZ��z���ފw��q�n$���\X�6�t�ܹV�R.}u�6[����g|I��Vڼ��.�ǀ_���B���e�ޡ~�]�dSq��9$r\_��_�`��m�eN�����O���~���8�<�3��0��
虪����Vz�gm[�Nbr����i˺����֮_)���v��o�E��]�Z�N�o� ѝ�j�؟�8��Qu��&����f�u���vˢ�c���k�;2���c4���~���^2�0�6J�tntZ����[m˗2�Jwbح*��gg��w;�멨����Ȼ@�8��ݝv��u*�
��O�+��s�ێ;s���جζ�B[�5�U�9%�8{��Q ���#��~�2L�j"R�|��ι�Lҕ =��V�����/o��}1���N�r6:�-}c	?Fq4�lDRq�0МE͕ۗj�=��î���spO��M� �3�� �nuڱ���C۞���F�9�B*[�`�T�.� 7��V�> ##�^z+ ̩ތ�@'њKt�=��O�Kq���9�������~�u{��$�¨ Hy�wh {7�vb�����rwq���8�Q0.Zd¬Ȩ7��fEW[]�&��Y�(��$�s*�ŎhQ�Ӈj^��f.�j���i蘱Rt�=o�'��M��w ��v����$z_�7�[��};W�@q�[�ٞ��� �wM5r�{/�i��	�KQ31�T��X�\���g����Mi5�vlsl�2��u��(#�n\��
S�����7=V�lH��7aR�ïUs�S���<��4@#3:��Vχ�$@��������][x�V�4�=��PmT  ��l�	7��6A&���������%���*��"a�PE��N�]��@��٫⽟PT�<N| �:� =��v���n	�&�.,Qefʬ�LҿY��H:���l@�۳V�@�g_��5]��<�:���X}��z ��'2������ګ �:(�i��X.q���D��Gń��ӗ�4[�_���	#$$ I?�I	O��$�HH@�`$�	'�H@�̐��$��BB����$��$$ I?�	!I�@�$��HH@�d���$�HH@�@$�	'�H@�@$�	'�H@�`$�	'�$$ I8��$���e5���Q�k�u� ?�s2}p"q�� k� �F�   
(  ��      @   P(  
 �   4   1TJJ�t����T���k�j	+LKm�;�	�4�M�V���Q�M���d"m�Q�-ikRUM�Z�`P��                                       @      
)'�=ˮ�Ash 2 hdK��J2>�p�4\��r ` ] 2 diؒ�i���   = q,�]� ���������@�� ]�� �#C��`_DAf��� J��QE'�  �        �doZ�r�{ q�K   �� dd  Y u�BtE"����x  @;9 }�=� �!��G j��}�ˮ���  둽� �tz�� }B��f��	/�           =�}��͟0kM�U^�t/-B��\�*�|�� ���	A�AsRO�E)r�(�\�U(H�� p� *��)r�

\�Q'�W��`(P��  Ȫ_,$���Qr�J )��� *�
R�����ХU<�@����
Q٪�@��� yRR�����L� ��R���U^YA*����q����4%m@�  �        �Mi�w>�ԡz�9���e+���P�� \*�35��=��w��{�*��� u(S6<�T�F�)L�lU7�  =�_3J���R�o�� tJ�gL��nگX��ziM�r©N�� ��JU�<��UfʥNڹ�E.�%���|   >         {�Y(\����G�;kf�͕J�u:�©O7 :�C�oZT��޸�yjU�s͝jT�x ��H��{�y=%((���   ��dX !�e
���4l� {ۀ 	��9u�� 
  5O�&*J�2�E?&��%T�@h2d0�7�5R�d� =��L"�  E=���U4��$�D�=T��� ��?����k����������+�9}�z���W�@�$��M��H@�nB		���$�hB��@�$�@$$;�=�_�����������w��s�E
t���v�2�8Q�����kaAdY�2@SܜH�>j������̄�.WxN���W�樍��\�k=�;� ŗ�jpa-�7��m�E�Mj��f�q�)�8F+���Iıv��T֛�X˃l�ׅG�ln,aYl�q#��lhћ�R�<��$��4.K]ۖ�Y�ݶݫ5Tѹ:K0Xs.���۩ل���	���c3����P�^��t�z�ٛ�.Kw]Y7r�m���ȷ�RN�p�y�g�sC�
���\P���p�#�͇ ��y�>���� sG��ԭ��9�� :�3�!���ֈһI��s���O7�)��tiI�e����wTp� ��YN=���X�-��;|g��w��隵���w�b��˸�kNA��.=�ٝ;&G��7cν:Iv|8"r�M��+&�a�V�ѯ0d�X2�S)�u�VA�Ҙ#Rnp>��s9Z��2�B͗V��^���`�.���4�S$p-B��)g5�q��h���1o.Ơ�8VML`K��orіt]�{-?Q)��Z���1Ms��w`c�&:ub���)kz�[��"�j
5�e�]�+�Д�)gf>y�́Ņ��:p�K�-8���Gt�)��jnj]�N)�'Mˋ���,=�j��^�tϪ���L��
�'O��Cv�Bn@���I�k�#�8�Mɕ�;�����E�պ��x�s�r��k��bz���[ث[��8XΒ��2c�6H�u�l+��ɺ��⫭&�.�؜�Dӯ�����L���ZS=�z���\ �ggt#4����;�Gze�&��i{��X�M�k;:�ʶ��y~kEї��-��Q�1n��\�����8́��ps�>]O\}��(70�����=��U�Zv�����1ۦ'�Q�}fqqV<ۋ-D�8��8(\=�td�f�9��������iC�Û�d���s&�x}d���p�,�d�v.�A��-�����^ӯ�yF����Z���c��_j*�+D�}��yH�'V�N[xV8o�]z�{/S���(��U��"�^ovit��ͤ�<3z�9b�1ADک�E�r�5�ȄYY�cf�R��r��G&�u׼�RD�՟���i�G���';�G�v>���'i�']P��^kO^�ɕwW#F�(��T���齐��9��]��h:��;�	w��ܸ:��p�T�}N����Bq�@�IٍI{�c��$vhT$�����a�L�n�nk�j8ݺoa笳��qD,�#ƫ����S��h�'�J��R��ުH&�[��`edX�ͱ��x�����.�+'K-ȫ�1�w�᳅X	 ���	sG]�v+{-8��Xͤ�� ��i"&��߁���X�d���DZP�]��Xk���
"a׼�.�뙬ܽ���/!V3:�w�"���)%*^�魽�C��a�a>�)�ٙFvvP4����ݬ8V5��4�;ۣ\k	2�2`�V��wkoU2"�o����ʴ�ȸu0�\s!������u����^��UZ�uf��w�烓��%�1؇��A����q�g�Ą���T�%�8��sP��:�=ܨʹ�[6	\V#�f=��b�� �Xq �d����v��
c��8>Fr=�;��z̃4zn�u9�?i�S�^y�GP�Y�
/5Q<��`�å}��$b�4�;&�̯�z�l ��ɛ�A3�^�>}��^�v63��OT�8Z��ѵ,���:�ͼ�M��1@H[�<�ۏFF2D��ЈoX7{��C�G�슡��i��wZ�b���i�M�x{��7��6�0����8��3G.L;�r�ͽk��h� �ppR�S1���3�N��FB�������ؔ^��G�b=�!N�'Ҧ��}ح�f��.�o6�<:+�q1�v}γze�X�aH*�T��۝���E��Z�h�{@ü��h	|D:�ֱb��WV� �t�z��������� .�W;�J��о������-w%\z�Sgq��p�w���<��/�ñȷV�F���Pk��Kk~In���7�.�ͺ0=a<#jj;���` �'F�Y�F���#�[���3��CqZ0��Ϩ���۷od����u�,���[M9Bɇ4w��+xs���~�`c�Q���YgSX2��0a�;@ݕqwrW�"�����5��B ���KYI�*�׏yOl-�8��.�*
\�v�\�*K�ǟkx�����V�$y��X�w	0(M��j��d���!�ML�`x%@l�U����fJ�o^v���2P�I&�"Ih6H2���3;���v�|�ɬvv����@u��2�22����������װ��n1WN!�y�����irN�C���.�S#{�e�)Ĭ���\�6�:�J�؅D1������kNL1��ǤK���WunH^�w:>��5��ͷ]���2�Y����6.��u��4���#:��ixyplPM;���� ���q.������(���y.�i���l��h+��֪1���ɍI����w���t���!���x7�v��u��l�ƞ̯"n؍��T�����K�zeG[
�7
 �.N{����M�A������x8r��)�=����DS�!3�]��f�R3���%�z#�(�X"���9�s��Lٌ:Z�]�uHz��flcq����V�Ü7��fEs ��'��
�Lb��v���������P�qW�vǮ�0`���[ӱ����vw,T���'%��=m-��+���M�͘��.�7,y�p�O	!}�<�y�!X5|�U�UKn�����x�qh҉Z��#}Lo��mr��Hf��,��;�r�r-�� n8aG����s>&�"�2��aIߥ�#�	�G&t���xv;��19;�bi!�1�TM���r�tr�g��磷q�{:�p����J0u��2�-�L��g�;3��EͻT%Q�q�q��+��{CԱ����sA=��%�`���7�V����"�U��M�m�u�Ǉ>b�H��
׫��]m��`L@�h����w���	�����br&a�nv���on��MJ�fE*�l�.��%v�v�?s�cQgqH�yu�yo�vt�
���.�x����c_V�������ǻ)�����`,�� e���Ѓ�{p5sx�E�.�q%@���C�p�D�v6�� �f7٬6�$Z�oɫKFb|�هw.��~g�����RR��x�z��8�}�7��v���|�=�OM�.���Tukrl��MH�pM(��Ԗ	��Edx3�1�h}Q����}�>իw�UL݂�&w��݃@U�m����:��}�ғ;Qz�c�wJ����fQ��/6��e`G��Q{n������v�-�B9�Z�����kK���X�R�ob��偽�,���=�ȑ�oRN;~��;��pm	�	R�.��������ݓ&,�	�����!���+7
�		���'8��v:�Lv;x&�y��u�Ջ�J���}�-}]��U�񵼟B;[�^���N��Y�cS�+�w�M��i����U�z�F&R�C��M/4�D�4{�4��R&��9BW���m�{��;9P+��,�7'``�����#78����芕d,Aϲ��'p�6Ҏ@�k���T��;&�]�Q��!pɈ�:�i� �OxN�Vq���wm6u�Z�n�W�z�4\�ʐ"y8zg��2T��?���رh�I����Glꝝrм�=��n��Y6�Ł�=} р��%� �	hq�����OU.��
z.wUicw�N�e�v����m#�L�f���ޙ��vv�_ {Q��}yq�uI�1��F,29��B��y1�Ǵ�H$�w��"q��_�a$�y�t�]�H(]l���;����yg	�g�>zx�=B�&�(��.�����,��Xĭ(�ף{T;z�"��vv�SƖ��`��D�Wf({�t��ۛ�2�W�xL�Ci��f�Ry��T�B�$Ɖ�4������p�դ��fQ�0�K�v֜[7L�u�Fl���@֡'C�2|8���5J4o�^p�e�Gt���{Js�\�*�<�r���'4�7��WFov(������5o N:�M��CrV�s�9C+@P;��F�V�M��J��I�	���ƕ�3���\<5���[9':v\�wn���s�n�޺tR�\'�:6��c���݊v��4����6�5ι���t�e;�3Wp�$��K:U�y!�w-s@XK��:��Fw]fuf���e`e�;G�&ͤV�T�(y���ɧ�v΅����䘒�j���Q�i��wF�:�{.�z�]V��q�2�����\�۳�ri�T 3h�ENM�^R�=�)L�'��!!wl�b���iLppa�s� �����s��a~�������4�#z���]���(-'*3�u�8lz�®�x�ְ�ɗu�y�q鸩�h��D�t���h�a�7 j�im�;��Ӻ�/�p�<���8���(_x�;
ȵ�F�f@��]������W���ۖx`붩�j���¶�萃V���Ű�(���.�u��;ܣ��	�l�a��f�ᄲ��3��"=bu9j�q�WIz�t�ѿ;А3��:z��T���tq�.Ge7�^T�Gt�O�k�rU�kǣq�vȹ0��.�# ���;�vLՕ謱n0j�xoT����Dr�(	9�:v��8�g�0�=G_i�'X��Ķw'�/h��L��u��)��os����p�S�!٫�j7tby���y#�4�LF���7	��u��f��+���q!+�1�ӝ�P�i�[�(��ķ�%�Io�[:�t��JI��g5�;��#��B���z�Cw^=�e���1���4G|/n@�h�ti��ێC>�5Yp#���Ãsb�I{.rY6����ˢ����9&���@�~�����%�x5����c%��ǘ�!�m��j��)"�$ίf�m��?��P��nkT�e�~�e�V'f���� �2t5��}�F�@��(�F��uc�$�>�z!$�B5jݽf�[%H#{vK̖R׬��G��Y�8��dq�ʄ���U	B��{�n������B�m�s�!��L ��ͬZzeNn��/T�v�r=)v���/n@n�XW%1K�E���.a� l��@S�p�ra�0ɾ�Y�!�h�hꌅ�!8a�d�N.�f��θq�=n�ڭ�R�}P�N��6�F�r��CM���"A2]��4�|�lr����va����`M;+;����q�[�`:NsAv,�2�f���.�6�u�Vc�è�.��vty;#W,�9��(T���Nr�����.;v�֑8K3�����g	���f�&�����H6���!	$�GL�޼0Tb������w�,�9�]��ԺZ��7��Ew��r �7��Ս��y�����f�l�$�b}F�/��5ߩʡ�^&,2ߪ�R��x�s�~��Jx֫�x}GA���1i���.��gl7���d`��� �B��z1e���<�I^ܽ;;"�44�A�0X7h�U��wr�+�����%c7���,`zc���I�I���~��+�v:�Ԏ/�l�p]�q��Ǜ�S�<1vC�GQ�;�nm��'d�6��7!���-�"ld�:�0�a�$���b՛�l�czU�k��#��vhZ!ܬ��
�nhz�)A�(�x��Xùa��|��������[l�Z�a�^��rg\�b빲��E3H�8Ab�n��W��&(��>��oL���� ��΃D}q����27���z�x%�0�'ezZ����ru״��l���'�4�i�7Z^����x╉�b���%$l���OT=�r�[0r���ɣX7Vދ���@��^z> 	(7�����[� 9���m�s���9��.�Au��N�=qܳ�V5���{Q2[�%����0o˻�ʾ���V6!�,��ۼ��ֵֶ4�
-'�s7��,j��G����O{`�N���<��ػ���Ȫ՜MJ����f��_A͛Exv����Jp#SM#�2Hi�\<���(�w4H��Ag!��7#�mה�O��ؕ���W�轈����l+P�w;����)�I;׶��������jٌ�uƱ�s�I���B���{Mk�3C��jZĈk�8���L�x������T��a��ǚ�`1�t;���_+t�\��\X,ݣb���Ӈ,�"$u�������o7�袅�a�@�r<J�{����Q�SȌ�����gp�h�owS�NGqXz�ܕ���!��.O<&�R�F�Gp����^��.�ո�N�ݖor��v��j�6��;#���;�g:K�p�37n���F~��F��bk;3�)�s3��D7��ݧ;�Z(�u���D��
�Ԥ٣A`^��>8�+�ny��}��֍���B~`H�!
�+$ �BJ���(H��I$*H
��Y 
�� �RH�$��THVH
B
�I!RI�I
� ,� �d���!BH�$Y$ �!�I��H�H(@�T����a
�Y$�H��$�P�� �B
@$��RBE��,	$Xd�RB)!$ �� d�"��* V�RHE��$P�)`�$P�����X@P �BH��!� V Aa�!�$�R
��I!@!X	XAa RI�$��T��@�V�$���@��"��E�E�� O���BC�@�$���{���]�y���3r��-yе=�6A�Gl�923WC2`Y�Ӄ3z4���rNԻS��K��2�������pi\n�LŊ�b���a���അ���W�y��+^����]�����H<��|���Z��Adߖ8�o�/�A�N��X� ܛ|���ig.=}�4o!����çJs���Sΐj+n#Z{�6TtL��)�Ͷ�s֩�W���䟘���1L}��`��[zYgfY�{��ں�Y��8'���^�E�z\y]�:�q�����3VV����#�ܤGthWt����6�l�_G�aȯ0��h����N�ߩۣ�6Y�����z2OzI8\�i�2>�Ԫ�0d��S���Μ;h�$xxp2\Y"���i��$��p�#�ɯGpͮ�.���n<{�����F�p�� ���U�6\w;U[t��=����o	T�����j�m�6�}�3��#/��K���W�U��R#$~�j][)Y ���;<��8ᚨ�g�tM�kf|p<l�}�x����4z����=�=޹���yN��J�nC���`��/��;��y'��ț��|5���f�ڽ-�KgAg�޽!��;��!o���6�d��Y�#��Z���_YH��w'58��>�]���=Ҏ�a{��M��4��M\�u��ɚd'wI�9��[��<��{dYǞ����e�0��_#�,݉u�]�%��;����vU�*�)	�a�q2���Xۻ�M��NI0;7���_oa"e��1�D�_h�<T,�{]�8�F��q7��spp,�x7��[գO��z�Ƃ�gO0wg:Nx�2'��#{V�p��7�z��͛&(�iт�}��)9ǅ:<&k�6}��Vv@,�b3v/zx<!�2�	��@��uY��^����T���ru��Jf��<�z躝�|e�}���5�<q��W�v��{z���y� �{*��A�}�p^+��٧�,�]���E�b�=hd�9V��}e�ޕ	ӵ�ő�[�ge�]��Z�F ���+���<g�ŗ�3�ݺڛaũ꽯��#f`��E��Rx�(�h��e�_O'�����<Υh�Y�*��t`�uy�m�x��P�y��$'cޯ�Od���w��>�+�؃F��7�Ys|��E4�/t������l�k\N���[�C~NX2�q����j���p��v9`�\ƌ�h͂�t]�+�7�q��� K�b	]Z�.�t�6v{:\ ����}m����:��ɢ请y�XÜ�ËU�� $i�W;^��~e1��o����箜���\0�!�&gcҭ���?.�[��y`��{�5��//'E�m�P�9�HH��3�{��=��"�t�1ya���ۥj�x����-}�<��4�L�������R}��L�o�)�q&B�	(fe^����ڵ,ԍ��d4p���-aH�k�W�_1�Vֽ���RO�A9����-3�N����h��Ďzf���\�E���ix<n���ENtTe�e��i����'��WB�4{�#��n�_v_y��\e5ޭ��sWH����C=rU;���F�n��Nמ{A锖�Z���`E�K�������k���!��H̺�X5)�7
⬔lLm�)��i�@�/��3��kĚ��鲡z���5v{��m�K��|+��d�u�����R���c7���γ�V��G֛�p�	y��:.S��Ӿ�..!Ʃ�9`�!l��u��#7*=ޢg�|+[|K�m��#�>^�����i�/z9O^����p�����,KyO���)�;�Z�ՠ�?G��Ӌy'��jRSd
'�n�I<	!��m��\ks�f�t������(���轋X{�H��W����U0�w���狻��dS�D��o)�~;m�-�ȡ42��)�~��x]�~;��S��:&g��a`On�ӽ�<���X��������7�\���z{��ަt��'o��	�������bwAW=����uc>�,Mhn�Gf��+vz.��ә�G<s��~�y1�����m_.}��F�k�4Wd]�"Rx���g���#���N��d��+�n�C���+���C�/
sn~N�ձ_";.O@[��*x��ȇ��Y~巙���C(��m��2����Ƕj�-��B�{�B�W"��JPLj�{��Z�����
#jt@�0����c�sW���Or+Gx���ד]�+���u,�нn#pm��ޜ�o`�<L=���|�Ȉa��{kw�^�r��>N�kZ7�{����[�,f�C�<@d_e~xY~^U��W�j�^��J�yB�ޣ"��T�����g�KS|�~z��kG��e^2�w��:����n��-��r�]�/E�¬��	�dŎ�-e�;��cx���]W|����jC-�1+/X�g���k�yz>���mz����7
�QƋ�^�P�"��}�ͣ��|���ו��?|ŵ���nYnq�lɬ>p�׹�D�o.M� Ts$��]懘Z ���<�D�" ��z�=�MA]6�9<�*�
jxխ>C;'�}ݔ�$t�/vAF�L�Q����?��g��%�Ƞ����w&�\��؟�d��>��|wzSMIB���[���6��v� �8y�� ���T^1V������t��v���ݣӠ�eZ�"�I���c ]�F�y��\%�>R�u�Τ�J�AƯ���z�9����3L��}�rbx��l^�P��abk��HO8���
�׼�m�,�/=�ҷ��3��B�N��/r�z�ϊ����%�DG"ߧ��٨�O&h���5���Tw�X�L/h_y����{V���B��/�ģ���ڧ�a�E#�xL�8{-M��ѳ����]|<��;�VJ(�C�=���}�Ȝ�\��I�K�;��X�F��p���-�����ɷ.�#x*Q�~06�� �:F���d���v�a��ŝ��ga�o�Ng'�����!ٛ�7ݻ��a�`s�؁C�yv/��s���V�M�>�SkVq�3O����j�I�|<7@Zyq~^י5�*}:'�����fzgF���=W��9lQ�D�����Sn��Iw��V�{�~��;���;���e�)�ؙu��߲>W�����$��rH��tV��8��:��x��4b�������T��A��
DSyc*F��_�k�|Oj{?b�R��O�^h\��*| fˎ)� {_^�Z�3�!��eR�tg�P��~�l�['�$1�|ﲓ��w���z���,Pca�W����X���JA����tA��Q�7�{��i;j���Y�̉w4\�RK{�=����׊;���3&b�j�u���]�O�W�4����B��S�s�<t�nݡ�8��S^�mg#�y�J�<����cuqU[�������<or��Y�E��k��:p���A���+O���د�~�z/i������
���"�����g���ly���m�%�`���
�;��zd"o�?@�!��~�+ƞ�7���f��%�#6y�<P�BV��ߤ�ÞL;l������ޗ:���&{+��&5t�G�����Un!�����ǖ��q�{���k<�N
E�\/�U�ǡ�޺
�p:�q���"���-9�Ί�]��,�a�5���*��x�5�&Z}$��%;��j�a�}��U�e>Δ9���3�L{
�W�����Qc�B�ĳ~N�f�L�E�2��1���5=�Vt���q��Aet�w�e��壤��)�-� �GW��9X����� or#���~j=���m���L��{9b�b>��ǉ��T����p���)���Jm��]�������@f���6͎6*���F,/������ӈ�-�5��@�����=�d�a�k��>��\�ya(��\+W�}�M'y��B�wH٨hɭ��l���j�n���C��y��*(� ƪ�m	���JI�C��ՠ��aFVw��E������Z�̜���{wp\�lH�������}�o&��9yj��@��G��~`��I�=��gv���/��h8w���xA g��DH*���j`��za�Nv౹��ؤ�c^��'��C_u|=3���N/r����B�8���o�պ�� �5�#^Z��z2�j,?���u�}��K��۝@���8���3o/Q*T�<h�|��1�E�D?z�V����k��{��yR�<�Ὑs���M���Z���+�*��G���,:�:�|��I�-9�V�����Ҍ�1{\@i��ݒf��e��Fm��0�����6�Ś"K���=�}��z�Y��BEn��������C�d�#ދ
f���~Qv8gT0KB�]�;C0��0��l�vl��'m~ɦ��%m��dM��:0eŸ���y��|{���`s�b�<����z�7��b/H���;;���	kpI���*-�������D�:�R���Pg��p�{W�{Ptm:�I�3�b�ߛ���ۘi/�,ʆ͈�w�p�Q�ߙ��30QYGT7p{�y��	��o�0�Y=�=A���&������s|��r<�k��{����OcR;NF'_v!�w�?i�ʌn����i�W���߲1w<��;�C�^lAfm��Ҟ�p�߃s��M���CwF<���v:%�¿Z�:��� Y�\�-	�?{_<�{v]�	{ڱ�7�+	4:�7����X��ɕ��^�Z˃��yj
�*��$��W��hs8�||H��3��P;
�OJ�ؓӴ��H��u�䧞��ܝ�Y�_xz�������D�g���\�0�p}�z5�d���|�u:�2xU�Ə��⅒v� ��7	��==�'`�ë���;B���jհ,��������0�[��7��H^{}`-�z8Ӿ�f/5���ru�F{i�#�zf<�.�b�9r��v@�MÝ�^Pf�eo���@��;� ���ٺ�Xt9|/}؆�aޖI{���l�Jp`����������9��;_�f=�C������8�鳞��o��En@��Yý�������%'=���R���Bz`+|G7�MąG	���A�w�L�͘�x�'�p�ְ�a��xn�,�OaC����F7X<�8��)�7w ~"�O��Y8�����8G����7��h�u�j�Ľ�������z_ue����/��y��,���+D����zd����qlUo�˭]һ�;�G��8EG�� w���C���V��뾂ݾ���R��xe����ו��{�MU�0��Ъ�7�7{��:nn%�{8�=�(���[�ˣwY��K�-�TU������9�kC+FdA�>\���z��v̟J^��<���ŭ��|������6.��I��_k��Ky�y^[�==&]�*{)K�h���P����x�\c6]R�SW&�Hwv	�uv>�O�h�9^�3�<���z�֜�n�9�ݷ(��H=M�1qgx.}�'ٯ+M��y};8KQ5W�0�{��A/Dm�Ȳy��]JY}GL���Cg�����R�\Q+�F��}��X�|��#z	f����Ӌ����U��@W�֕�����z-azD���ܯ����{��E�~�˃
�1�=�R����q~�O�ǹ��8���� �k���U���Q�8ߑw��U��74y�dˬy�"�ө��sKW�x��p�G�6Ǘ����=��Ҿ��x0��� ���{\~��`��(v��]�)�d���^��|
��-�w��:/�ꁆ�M;:zAa���:�{ё`!og���U���;/�;`��K<q/.�_��&9��ջ.���Nz�Ly =9��z���y�<,$]j�1X��캧���*��ɉ�>M�R1�I:����Xg\�Gtk�g����'׋m�x�cfO�+��O�Ӷ	{«ZEb�'U���S��Xe��7r,��zs�+N⓽q��#^�mRq���<ǃ�M�4�'D�'��˕ٳ4gT�k<�r�k��/��9�y �.o_i�"8Й��>W9b����eX��}��=�o���S�4nz��§�V�2�p�L��q�*7}��r<�j�4�Q���h�9�f��hY��qǳɏA1�<��m׾G��^壁��\�K���l�I�9�ӛ/�
z�noA�M 4��[ö���n�h�ɷ��[�N�.��6-b�dUy���.d������, K��z3�,�r�u�d�W��-v⾟z0$��%/vMC{gUW=������$~.=֌ż�9����id{�	����c��2��؁z���ݻ��l [�/�?gP������f���3f(�특�H�
�hȼ��~����b�<��Ʃ�����`�|� ��nN�ۇ����x���O�\���4Y�P��Ci6SJ�Ɩ6��5����2���ZwE��=�P�vgI�y	��G/�{k�^F-֞�X��%�=�J{ J��N�$"~�N�{�3No��X����v=�X����0����tz�;��&lZ��+��z��l	�� Ѥ�p�����]����[.��� �|�~��;!8��yf�;K��y7�w!Â���Pza�-�|�D�}�=ή�
k^�>!)�#��&0�QTPڲw&T��o��R�zpܞbo��Z^�y!�=�U�gS��o���}������S ��e;���*=䩾��u�wo��Nr�dbjt���c�u�������3�w�_�H@�zI$����Uعg^��x�q��*���pM����:|��6[�X����A�7:Ǟݣ\�S��X�Z#h1��QS��3��k�wN���˼��]���+g�2�A���=p�w�r�+�q�8�x	��<����<��4[eSם�&�n+� ���|��^�қ���f�6Mjۂ�q&���+��s�Bc]�T/Y'<����%�ے1��ɰ��1�o]J�{Mm��n��K�l��cA�M�[v(���W6�'۬�h��˫ϋ��a9��:uv7t�r5����a���65�Aq���mt�уv��kf��v��؛�=����p>�;@��8��'=w�G6�m��eӷl\;��V�	�=��;��v�����˜�u�b�s��fsg�-M�`�g�͸9wF(��Q��eG��'�T\k�v�%�]v�l���5
q�Y���X�{��e�9�q�e���]�B4���4c�O]S��;��Į��v�rܽpOhf��m��k����<q�%����v�4nv�u�[����W��3�q8��ݍ�3n���B뢵��z���85Ȏ�����r��n㷮z1X=&��݋pI��V|��P�-;��V�H9�w"	M�t)�s��\�c�"P��8��v��3�1��W\v�����j���yӠ�.P- �%��c���m�؆L���x�t{!���vn�/Pc���`Ղ�4��g=�2�0W[�8�Zع��7���F���9�&cN�z�N�#��cj#�׫�Uvؚ:w@Ic��&�͇7a�ƹQ�g:�wd��;��꽈����nۇPv1ײ��r��ц޷1����2�Á�dҙ�g�e;oU�;Vg(C�����],)�������nی>^��z:F�N+us�z��6x�y�8��ufTH'���4a}��cG6�GB^��8ӛv9x��Ɖ�:�<s�]�¬s=��#ͱ�
σO��c�Cn�uc�;�2kY��Ol<]ϝ7N����Єm�"�l�i;=,s�Vە����n.s�\��×�b�cK.����5L/����˟]��
vb�iq��-��Ճ��;=s�k�s��n�ck;��'cN��f�R^��n�u��v]�S�{-���of�l;qp��by93u�a:�}ls. �kl�Nz!�S[�X�H.�d��Oux��yǛ�;q��-��c�,���\h_���� 枲:y]=���[��m� ��ygs�vגՙv�����Ѯ��^ն����f�pmՎނ��h�l�:N�Xrx�m���Î{\�H�ci�n4�x ���j�5�r-����.�g�;qm�e3mqm�n|C�kɍ�;K!����9����x��C�J�c�㳦�vδ��:���ƫTU�lj�b���W
���k�p������7-g��U�z�l�Ϻ�s�+%��y�k��a�ÁnY�k�=�;�ּn7=��7p���c�l�L��+�|rZhzu���2n(�\έ�v���Ȼ�OYyMq�:��d�v��9��f��=ۮ� ��:ث[��]���Z�d�D�� �.��[���컭br��M����R�Y�Gs��wfx��n�C�1Jx��z6rn�����q�E��zv.�o-�qn7E�r�p��v�
�����Ψ��q8G+&=���t�i��n����E���Ʈ�r΋x�T�n�xm�㶨[���>`�Ng����iڝ^us�.ӮƗ�Ѭ�;"v�m/4�î�s�r��g�ޒۭs�vô�;1G���F�f�˟��<V"z�{ns�%�N�<WF.8y�v�G7��2�ݘ��&�;�ۓu���{x�����X�bn/n_;��Dz-F:��p�;s�Y��,�݃Q�ۛnK��Z�è6�ܻ��[z�l�I��!�S>H<]p/i�,I=ѻ[^9��Y׶D���v��R�.Ã�[I�d;=�r�NM�st�u�յ�y�-v;Q����<LdB�u���ێvs�t�W��3�{n6ʯS�0=]��v,a܇t�%��9���#����sv�\"'΢%��N��S��������^��ѹ��f�.��;�����U�dZ�������V�=ɱ��*� ��v�O=�M�<n:v��ilL眃]���N'�����n^�7*�8��m���k�6���m5������ug�0��z&N�$�I�e�%���s���;%e=��k����3�pv��Ga�v{Wm�C�a��NPC�lT�v�s���m�z5d��y���xL{vg	�N� ���M�%9	Mm��f���^��Gn��5�p�����6O>�vwu�08�Y�g�]v9��Ӕ��H�m��x�\����rwO]z��:�us�1�NN����'�8���Luk2]X������x(�1cf�"��v�E�f��ӷn�'x�S���]�u�N�p�ѫ��Н�cu�fm ���)�ƭ��.9�����CQ�3���@뷓c��qhW��\l{���8�-�SR��q�<�Z�<W:��x��^��y�u��El]��㗃6�<Ts� ����b�u�e�����q�oj�lf�q�ힹ4;s�:.y�]![O9�N��]�j��%%�g�wE�wd�z�G@�Lm�9$�J�ɸd�*��7�c�ws�<v����n�k��.��1�%�͎T2r���R���� V뱝�����۝v �]�1����;\�*�� ���ڍ!ؗ�r�7;��ݐ}���1�[����;"�&����Wn��Gk=t:{�������a]ge��I=K�����ܻ�3����õ�e�����v��I�x�杭>�r;��4�m����j��n����י3���2��a�ܬv�$qu�׺9��y����tc�m�E��[���p�#��ۋ�pK�3��jr��m�g{Rm��/\�gNBÎ�g�Cw"�[(�t�/�+#�[���'%�3l�����xۏyы�������s۴�	ǯ	+q6�u	1ۓ��d.�|��r�J�ӫO����<ۃ@�wV4u�-��rU���������;%�x��u�\�0��v�er�3����mr�X�%����v����]����z[��x����7tk��ގ�v�8&��	"9�ˁ�y�kYg�\���mΉ�5�Q��v4py�=h� g�y݇g��8�`�<�b:��<�8{vJ��]��C@a����綆�[4ݷ6���cz��r��h�t�:�Ws�{�[�0���佇h���#�vݰ��)�L\�Z���!���ر;�ׅ��z�F�v�@#R�3]��cZX�R���h⻝���ݮ��pn|�"����;d���,��kv7j��
�R���.y�gY��I��<�N�|��˪#���Y�CW4�G-�Lb�}�+��UmX$. q���n������ܑ��q<n�C�q�荶.:'�,ܙ����\v\��)�Y�9ݻ;uy����%�ެZ��.�q�{t����F�cۛ�;uyٵɒ,��ʤ�8��3���r4[�ꝸ����k۞uDs�u����rb�4Fw[p�����*��ٷh���@���˴<y�x[w6�nZ+�ۙ� ��P��v띝��nPe�nw8��Y�i;7��>�� �ˮ����+!��z'���H��m��k�������Ň �u>{"g���nI˟O�a�7n{�h��::����qp��m7V���u�m!���m�7k��V��&�OLQq�Q�yâ�N�Y��]�gq m�ƌDr�P�y��_nz+�����q��s=!�5<�;k�αQ��\��qnM@.���a���n��a�i�M�"�����[#[b�	�:۔�cawX�����gv�TQ��.lY�.�JE�y6	ƶ㴡��v��z��<��6��)طU�|˟T����c�q�B+3&�SZ6�v������.2q�)u���z6�n��֮�nC�\m�n��J�����ۈ��V����{vtcZ���a��x��ָ�@�����6�N�x�<X��L��]v�[��۠���N�qػ���K�ۮ��� ��!�ӽ))��Ν�=�-�;	պ����k�6������]��l��n�ٻs���v;��۔=��q��9��0kuNd�6;8�X�{pm��Oi�ݹݶ1e��y+�.�%t4��8m�ry��m�=��m\�	��B�p�%[q�{p[��{!��Km�v�Qf"�ܻtWv��^��cm�<c�vGT�n!;).���YvΎԽc�mz)x�ܧn#:�wܛ�1&����Q�^׹���@a+D˜9|<z����L,�uqn���iE�`6�n�T�����{[T����3��Omۮ���aws�60���hxq�e���=�=V\�mH-� lTr�y�D����2�˚�RI��J#r�un�<=���n#�J���h8)��֢�3uz�`��+m=��$��7Pr������\�q�r�����]W�PvPZ=�ۮ���\��՝�[fūgk�+��y8+=<��v�6�g&�ا��n�u�K��%���G��/`껢nu�l\I؄�G�<�2n����Ѵ���W�9�7#�q��n�=�vw���� ��%1�<�Ǳ磖:r;vnm��v���{A��4QJ�n�v�g�Y�8γs����$ǘ턹�d ]n���n���`����1;��)���s�.�^���
ˮw6������A��V"=��]Ao2��Ё72�]'\h�ٺ�wC�ڮ�g��\������c�T��fc��B�سӒ�͵�y��g����b��.ź����5�f2��QX�b*(0ADV0UUDc[���*��J�mX�� ��F0b�EQ
5dTm�5��UdQb�QI,�mVA-��EUQc���-�VDV������e��+V(���V1Kh�,aQ`�"�F1F*�D(����Ec�e��""��5�UJ�`�QE�F���DQm,UUEEҶ���eJ*,"-eQb���F*�QUH�UR҉[TX�UX�VUcUA���#JQb��UU�,T������*�b�V1mib�0��V�Um�����e�F%J�1b�EH���H�TX�� ���i`���Ԩ[TTH�2,E��Tm*����("
�e�KA���A�hTE�P��UKmJ$�k{_��Y�	�s��������@��;���;���Yó[u���>��y�۶�K=iqZ��M������n�7Gv���g��dC��U�3̬]�wd˹�.�T����ۆn7Vӷ0g�Ê,x�Z��F۷9zK��cͶz��K��;{�v��n�[s̭��k��N4��F��`�ۙ�E�wnn���V�S�8�{s���飐�&�<H��Yٹ�\U/����hۭs��qf����W�w\˕Gg���M���;7j��u�;J�)�<�yy�lv��F�s<m�^��ݷ���7	g�q�s�..�+v���.F*��xݵY�/=�Aiz�f��ZGP]��z�\<ZzͭЯ<��u�V��5��3&�ZX7�.���o��O/|�CS���X����9�G ۇq�<v�8l�;g��춲�D�\�	�4{bnb�m���n\c�aU��;�ú�j<u� ����'�K����N�:ҽ�C�3� �X�u=���Vi�G10�g׭ϖ��ӝ��TD����Z܈F#tC��)ڣz�S��tM��"�m8(������;{,hy3�m�뢔���n2��8X�Z��:�\�A��������U.���Mףb_b3Mu�Z�nk��Wu���^v0]���b��y<녻�]�Y��>m7��g�s�]�;&�;uh���E��'.v�n��j#��0p
��ٍ䭲6{;�K���m�p�4��ۭӳ��:63�����Ony2k�y�in�q���M�(��ޮ�:�f��H�o|��|��N:�Lv�����,��N��Wm`6,q�x:s��t�sڪ 
�t9B�Ƨ��:����cUv��8n��z��Oq��u��\�b��r��Y���wN���A�.���������:wF�L5n�❞tx��k��{#��:�B.���{��E����%��-Ǝ8�d���eE�����9w'9Ï(�wێ�8^�q�?
ۺ�d�wcÌ���N62�*�Qr%
f-��
eS-�9糐�3���U��m헌l���ly�c���#\���֔s-�h�V&Z�B�`����W��0�x�0������99۸�NS&=��l/��g ����;<��~���$[,E#
)"Y��`O�K�����;��-���huL��q�)}�U��1������4ެ�˜��	'�O1���d���|t�ӓ�勒-��a$�S�$�}�����{*�V����']�$���1@��	%>�!�Idݜ�g�B}�u����:�����W�M�{��e�Oc����<ٞ)"������݂� �w������]}���'�W���A �nO��}��-����q<������>�RF��0E�#7][^�N�%�y�<q�S�"N�m�u�q�_����Uz\�_����̔A����u��?.��(���R���`�/����$n�$q���o��Y5Y�պ}��/�p����ͬy]i��k��i�gb ��P� �zJբc�-]e�`5��8�gi[�5�ĐC5;���]�R�)�ĒOoeC���}Ky��;�S����ߴ#�V(f���}G{}��@5ٱ�g����'�O��(A?{{�c�+�JH�p(�k ��m�K�w�0I�6
$���A�~�G!�;<	�]�a ���_'J~�"�Id݀{s=X'����x߭�>��0���|��~@_�Y~�(��O@nH{�:�q�����n�n-\Y�!�n;/q�7t<���	���)"q�Ґ���OM���� ��xC��vw����9�_ۻ� ���vci�g�87`Z��@�{�R��FeJ{a	��'�:�~��Q�W|��"=�1$[,I#'%��]�I����$�����~�Ǐ�6zg�?rB3�	�O�e�T�8C�K�q��Mþ̼"�>j�)�G���L�yq��r]�C��߱��~��u�>/���E�ϙ�
������'�]+y�	��o]�d�#��|H$�<�{��Nvz?c�˿��/dJH�p(�j���n��}��{���c�*�X����e�~O��H;�yI1�Is��s�{�,�a�E�*��n���㗷��c���e�q��g���k������M��w����� ��k�A'���,�|Ǩs>����A<���8ٜ�R�p�!t�{_"fX��>}���+�H�:�g<��]�Q����<�]�컳L�1����yξ${�� s<��Vt��`�����$���){�$�����wA�2Rtk�Ad�x���~�لP'�}�~��+��븫���=X����7|;����Kh�ʱt=꩖�h���v�?hk,��2��l�&��Xt�YZ���_�Q�չ�-#�I��OrP'�X���	p ���?R$��{�˯ʖ2��d
�ԯ����<�ā��|7�+�\9��9���	e�]�O[�7=��4�X�;pܓǥ�c�=���;a7}�qމIl�ڌ��@�O�ٯ)E��U�s���x���2�M�~T	�{�R3%=�"�Id�ο^X^+�G�WAR�V	����Ɓ �_uY �꽞���T��d�
�8J����׵�$���d�o�]�]�]�m��~�0{^R����.���(@�q��[�G�n�ݐ��?���A##�� �7�>]��h~��/���wA07r��{�b�Z� N�Zʤ��	�x���o��v	������ܟ����ieC�!'�L���$�2��m�2��U��s\����/���U�cN��Ղ���<��~����SH�0+78>ê��+H)̯ä���ל=�lz^h�.�qZQv�mh��o]7g=<�un�3�����+��)�']���ڵ��=��7���f����kw3��[r�6�3�i���������{R�٧';�n�"b㸝G$\rn��j�9��=/=�"7@͸;u��ȉ�N|�>��i=�s�ۖ�G�����d���ǩ�ԣq���v�s�tǴ�A{�u���n�U�;Gc=-�U���������ߙ"0�z��"��m���J��U��u�I��}<��ηԁ'{}�`��}�) m�Q��I�ɯ�w��{��W�$��
������W��j��1��n�vdl�S�`7q��;h�L���w��'��{n�$�����	̕!PGRv��s�t]�f+�.�� �Hv����P�����<�ζ�]��e��"�ݫ�t	���d��n��An�'�;�.���O��A�vJ"�o�>����#i��$SPC.\�:+��"�Ś��3Ϝ���:-ӷ�<8�����C\�28\�N1߶ŐH:_�� �wݔ(6��46J�L�N'�t	�X��W`���Q�����|Ӕ+�^��ݸ�=�*m߈�W68΃���u+���T�����C����\k��W�l;==��g��A��ŝv,�Oڟ��$�{ݓ�+Bzg�C^s�p��I�j�g5z[�I��;%C��o�n!�=��O_{�~$r~�(��vJ&eS��r)�FM��{3���\јf�ń�C�A�vAD=���ͼ��	������b�1�J�*B���� �g��M�#r�����'���_	��+������׾����z�C���HAD?�5�܊�؃\��{V痨����.��p�@�����Ўm�0Z��}���{ْ��=��J&�3>%��W��~>��@���1�`n.G |���$u�Ǟ��
{���7���~'�E��}@�=��_��{�ow�w]c��;��`�0�»=~���$��݂�B�0���}oGW�wf���� ����&5�7����ɻ�_o�D�2��{�q^z
�:�?6+E3WQ�~�r��2���T��A'��(����]�ï"N@ہ6�45?[滻<9�����q���A��u_ē���?f�"�ڽa �g�|	�]S��rG�FM�ǽ��	���GeN	��v��~'+r���m� ��s�#����?A'�t���D�	@"f�^��Ѷ�]:�
+s�J���h���"PE )��U� ~��` !����S��e�N���ʻ 秹�z0��҉8�I���g��q�'m\�$�{��'�����"�;rQ9�1�`n�G%�zŐI���P���x�h���YC��7�b�$y?s��"�X��� d�c
����KeU(6�%����7׻Y$F'�u�?��t�x&��{��R<����9.���[�gOf{7�WY��f�/M^�{�z<yϱ�'T<�[���iCd���K��c��������xbq������Ku�gd��؟�0���]�A#W�:'�N��WƁj��r4����~w���Fǝ�:�f�������Gr�:1��F�d��k��rI�(�z� MtA��e
>��������zW]�I������-H�@T�W���	4 ���OW�{��m��?	�W�1_��~�j4���=u�$f׬��q����n�g��$�}�(�I�k���;��$5zk���d�sry�`r��G%]7�����m��|Iò� A��W�Nog_�5��i?5�N���
�2Dd�a]�[�J$��ٷc*��o��:!!/z�A'32W����f�T`�x{J�Fx��i�V�u�����=��J�������-�:�#�'�idX�욟!�2���Rf��oMe��jv6^H���<6��9;�ϳ�vA��`��6"7m�^!q�ŷA[8�S��ې���v����nǄ@�ͅ7��A�;r�c��8��99��[�6�#�mԆ����e��K�KНG\G��WG����c�(�7u��cI��ی�f�x���e�"&(��2=9I��\�c;���M������d���	;no6��|���.�Z��=�MTtt^S	Kc��ɝ��v�
I��)���θ�!m��P���bj�������@�}W}�|�����Rִc�a���t�ے�"�T�8��B�Jvwݞ�%���]i��_O��{��	���A�V��j�K=�h�v<'�&)a*D���*�97e~"�3��?_�����U�_��(�	��v}��F4�L�$)���rs9;�7�ҁ �H�fu�#ޝ8L�^`����qH7]PW��iDc��!��_�`Y����(�p��.�,�T	.�P����~'��N�i�fm+�g��$[&�IihZ7Z�n|ͳ�7՛uWn��ץ���w��}����Z#W�׽�_H���G�?J/k�P�ł�^��	?wfm�'�^��7i�(~�DvW,��3��^��y2���P~��u#�^�Zf邧����gf�g�;COz�Ŏ�������r�-����7�G;�gx:��گ^�Y�2�rK������A���@��VR>���k��}�*�V��H�m@n��vz����΁$���X�o� �˱@�~�nm��zs��b��M��*B��햍c�^h�zm��vݐA���@~��w��G�o�o]�:`���;�j� w]�"3��L݋Yz�~7ِW*�~J�d���'�o]�~$r��_E�d�Z65{�i�?�֭[�n���s�/f�7��Fzm�����D�
&}��Q��c.C��4��vI��:'�I�����~��RR��]�e�'O�:'��^ă(�IFٮ�]�`(gxb�w�s�
"���|1��@%z�s��i�U{�{�[� ��a1�P2ق�'�u��vJ'�M�>���;�����������eA�廳�.t��X6��>}�^��&,~�c�E��u�y��9׷�_t&O�#��H�����,����^g=;��]�oW����f.S��{��RDC>hqC�=t.�K�g���G��)�O�����o ��	������ҽ�:A�7�).�3fr���ou;���ewfp��q�{�ΐJqjыp�|dɬ�a�,���޵d��dQQVzZ21��=;����qr��ө���qB'f�(DȚ��m��������6��{<`�������ub�(�
w��m�Cb@�� k�Rߖk^�Q�Zv�GA��9��x��{�N[�3r��E��=���
N���������a��%齯���,�>�f��ݔI����G�w~5�{�(�?6i/CЁ=t�;����$�8��vQxW��r%�<�]ii����oM�oҍ��y\�d���ě�g�ס�+dK�Aヱ��s���LW�<8��MN�"m�fs\3��}6{&;6-��5���g�;	Ы_�ɠ;�U���{��Nۑ�Ő�Ӗ��wʼ�bd���s��g9*��e7��^L.�_g�sYO����$�Ǫ2 ŧ��w8o�GB�ʳ�&ߚ���|�� /�.� �r.��˦�����.f�m^��o��1Nl�oP��~��L�a�+n��
��Ď�r�F*S�W~dy�5?2ش��:z8w7���f���~tV�Ex-{ɽ}8�"��8sO��A�����_��b�o��[�@�r���}�/�{^��u���|�����k��a%	j1�*(�Z
V�`���-*1b%J���`����A-�DQ+EUV���YR*E��#m�� �mKE�ej�Eb��EIPZ�ժ�X�$Q�,e�Qm��QH��X(���TX-���EaXT��ZԂ��l��
QT�T�*6Ղ[F1Z�TR�*��*
�EAD�
J�PEZ�)R�UDYV�b��UX���	R���V¥�UҥJ�UA�YZ#J�a[h�´`��b�(�Z"""+DE�PPTA"1������Dm�6�X6�KJ�b�U�H��"��YR�U����TQA
�E%�b���1TV �A�E��,F�ADb��¶����*��(�i�Q�6���j�U
���m��Qb11���-�(�*�"
�� �b5��Q���QQ�,Tm��*�1F#Q�b�Ydb#-��ֱJ���b�ZX�b%j��T]�y�O�{y��h&��Q"�j�(�rEnc{޳={��I�w���a��@$���B� ����My��{���{���)<�)"l�RG&�I�vu�nTrϦVTҹΉ$�fJ�3{:�f��8*�NʿkQ�%$RBQ�ٌ�M����M)Xu�����1�M"Y�P4 �n�" �C �4���x�H7���$����+Å=|�V��<~$�v�3r/#��T�7%}�Y'֨�U��"��H=��(��Ϋ'�h���HS��nʃ&��/�%U��ޔA��nm� �s����|��ǉ�߳%IݝvH<;�LdD��`�����g�:��'�%~�Gn�ݐG��2�,��G�F���R��K�v�:�>n� Ǖ�cݫ�Oh�O]�<�ML�vxE��v��bTm]�>�}/�e/dQ�fa��|�No��N��6ӄׁ�v]�d|}9�ugpeW��{8`������1/j�������� �t��z�X��.���{v�k1c;��m���:�Zl'[��СP�JB��gJ ���=�,���ӝ҇+�(����Q�پ۰H�]�d"E �4��ֲ��$Τ���M6�$gg����Ή6zA�.b�����2�1�罖~$/��}���9o���s3\� ���m�$�t	���21��+Wr�\k����W��H9���?�~�(��vIV�^!�п�����ᗄ�A�ϛP���G���F���X��ľ$��vH$j~�D�H=��G�R�7����m{�z̙pכ?u\?/w��7ݿk$Z��=�\�S�u���m�	S�ķ��8<��i���[�N#5�:^\�/6��{u���Ń���B��:�v6�m���v�/�v��*-=[�+�2��m�܄�iŲ����\�������bE.rΝ�;!Ӟ+��=�x�d�=�n�0��ݼ�v�tg�;<j7��k��q�tt��N�u��y�������V��<n=�kE�R;O�w��d��q�����;�IH��=$v�6�5�۳�1�7�ۜ��r�{F9�y��˹��Mf��w�����fb;�{r��z� H=��(��X�W	�k.���*�쓥�] |X�r �Ќ%!U�/;e|	R�{I�H�H����O��G{�P �=�	����9��{�'>�H$3Wj�] A�d�H$�������^$�u��%G�"�b��ʐ��v��on�gS�o-4��A$w�(Q?o{�{��)l�d��Ή���ЈbJ0�����|I���z u�O�����$��l�	��������YG6�O�H�����\n{kOu�����43�^ǫ��B7G�I���6�-zS�~$���$�ogU�֋����Ϲ\#;z��I��AB��h&H�f2�F��eeX��Tz��ם=�Vu��s�ឳ/-5���f���+n�����<E-.��}�݃E%��^5S�ʺu��� 	ǳ_߉�������˿��^^]�ڏA����%��a)
sfA�oe���u�w\|�%�������o=Ҿ?��˲~ɗd9Q8\v-Vs�3�~~�A�UJ'�I7��b�?b�s��}̪ͮ��s[�z�$7%{�MF\�7 �{��d���:>�j�fe%���o{��qW���+7{�=���B����m��ql���%�ݷ;��-Ɛ�s:���śsɄKW���j0�[�.�(�H=�ܯ���K��u@|���(~$owe�ë�Ϙ�"f8��=�}�J�غ�Ʋ��	��gvX���~�@�����X��y�$�?A���N3n#c{�d�|o��~8=����*(uA*%��`m���f�����Nxd�L��Cpg�>��B�9��㬺}����pi�2��E�ryT�g����*�����<|�sk=�:UL��.f�`���T���]ת�����Wă��]/�z�>��mv7�}繩+v'A�ڬ�Dٙ(��ZzYX�=���'}[�`�u_��'�A�vJ/gd���nx��[E����1B�lo��\p=h��Ҁ�8��R��n�D�������š.Z���=̿��I�^�_	�(Q#+_o-���5s�����K����:P8a��Y���ߥO���k���Gz_��qW��?w�ҏ�1]eS�{����g�7�}�%:$�WĒF
�����+׹`O�S�����(A�\Hr'��!�nv������?k5�$��=�޼��w��v�1K{9q�hz��sHF���~��On*��9jMgu��)�f���[��7'�^�XsW��U��6����{6]��������<�0�$�>0��4zg�@�o��l]���ڇg��%,�b�>��P �����!\�}ƿ������aVwhxMƻM�n�[:����X���nL9H��L�ٙ�9QȜ|-Wk�	�{%A��u�B�T�^9�$�}ْ�${r/"m����%|ww�? ߁�����8�c�I$��P�������O�gO�<�������bn06']�H;�λ$�4�]f�O���tAٙ+�	 {�:���#>a�m�+VJvg{��ycK��
�\�H$�n�Y'ƽ�h�J�ZzH.{%|L:�D�1�7`��˲G�{��V�W��<�`l���o��<����� ���!�꾜ǎzfe�N�xޯ%��_j�]���{�����]wI�/��z�^�OzxI�ڏ��~0���Na�9��f��-O�����sZk�u�%m�V�qq]T��&Ck�ێ�*�u*�{k��^�F����d�u�2m��ݽbL��.��n岘�&�=�Ll�M�n:����6����_<I���X��u���\��V�P5۟C�n��W�՝b��׹�8�m�ӭ�G�U�����6�g�Yۚ�۟gp�Q�����.	^1�w]ubs�=q��sps�y:Ć�nѼ�v�q�m#r]� ;+&�0���F�G��<"Hs�n����}��`�|���QV�sA��)*� ��������5 B�Ӏ���Vs�ATk��b�l�d�F�;*���:$�݉A�_�ϺA���H�nC�G����H:k���U�D���������vU�H'�+�:7��14��A`(h�?9yv="J ��cc� �˼ ?O�l]�OYq	ߧ��@<+1�e��a�_jڧDy�(`���:>�O�Y�vH$j�k�Oă��z���B����Z%|�S�L��9K��T<�ӷ1��1�6
AH�,0���L�Cw��N3n	�~��~$�׵�$��vA_=����*X�L��'�N��:'j(��4��gl�A���_e[�?h�g�z蘶֎L��͆�&zf,�pX۽܄^�=�s1�8��;-��]�-�bl^-.���*�����y��~�E����7��msr���x�=ܕ{/�G��r[�8.��׀	��fJ��fͭ��~���#�{I}�vE�H�p7!�H$��wGM��6fS�I'w���}�eu���t�7V�z/�Qq ��(��=~��A �o���q��`�����I��;����ݾ뿎�Y�/aU3�T�L���E
��S�7Z7;;�[���
źWϭ���a�2�W���~�~��,&����$��H${w�w���'vڼr�o` ��\�NՄ$��b-�,oO{,ݷ��S�&��� H'�v�]�F�=Y|K�zDM�e:����Z�9�9	]�f ����꟎��L����E�{Ù��?@}?t��;힆MQ���ћ&M�R���ׇ�8Xzu�n�Y�ob�g+����}�<����+�	�ٟ�� z�!nB�q��ݛ��ݿSY�.��{�M�:Q$�}��vA���U�u�8�|IrT�Fv���8#�I��m�]��o� �1vm[\SUM9���	������\<~#��v~;������Y�lT�]�v�o�ݻB]{Tz�<����,���q	Ƃ�f���(�����I{��(b��>����(Iٝv	�^>m�XL9����������2<w-���D�	��v~��ҁ&�VhV��@Vv�!$N8�nCc{Մ�=~�D�I�ʍ�X����r^�Ē�sn�_�P'r(g�4�&�;}���;����A۹����U�	��F����_|$S:MW|����������av����-ov�xv��f������`[� ����n�Fep���so0�o��P�3o?��}����$^αc.j�i9peٺΔH$�ِ{W�{U�N��*�� 5:�` |<�\��Uè��er���xt��F�DۂDKA$Q0��oRE�$!�`�ues��w'h�|�����y�n�	$s�g{lY�:���'�Noe
���>|w����u�v,z�ҁ9��0�H
���]�J�R��f�������~9~�@�Nwd�łfz�y}&g��m�'�6�L��vI�I��'��a�ϞV������'���A7�
�;V��'I'!�����u��=/��̢AL�I?;7(P$=��"{���l�^�J'�&АLϒ��M|r�e~$��:�ӫs"���Y?^o��$��@�	����p��/_�\�k�nĮ�:]s��H�튰����'�8���a�Mc�r�E�B���q���ʉ���}�������վj�t��X\播v��n�V�׸b]�۳����|���h��}Mq7p�!i<oc{�t-�7���9�G29}Jw��9��]�\�!�uOn��x��˸)S�Vy��Ӥ�z�˲�-*F��^�y$x7U�o�%�i����-��s��V`BlGA�us[���i|\�,�x��d��i1�×�j�:��#��[$�}��5���b;��}'�����8�T�@�ȿ[S]n/N�H\>s=�L�W&���!�������q�Nn��v[����|��&xU�}֌	{š96�t#f��T;��6�4G�}��c�z��8��=ƅ�L�A�qBOE6zf��OB3{��ۜ�M7��?+�r��� ^?qx{G:L�o�t0!�Z�l>�&Μ8���9.�6�/����N�H�u-sZ��Y�}��F��V����G�s��߬�sE��A�wy��#���^~5��w����=�P	�.�d�m���Gѥ�s��M�i0E;GG��GA���wJv�˱�K���;�Gw�t W�T2�!k?]��������,�f>Dɧ��VF�4�f�6bX}�bb���S�;.<�]B�܃��ˤ#���r��z�����xQJ���3��zv�^�*����۽&V�{���3\��J�*��TPm*�����h�mF��Y�,m�k-h��1��X���H�DEQ�A��F1
¨��U""�*�1-��,TbȨ��Ԩ�Q(�5*�ab�EE)+A-���Qڊ,b�*E�[mj�[*UUD� �
�+�VTU��[j�#�eAQb
�"�
��"��X�AeT�V���V����T-�)F����Qj��[JZX��i*�m*0�V*"(*�բ*$DDX�(�����+X�-�TT�+*������*+���Z
1Q��Tk`�����F�%k���� !l����gԪ(��TFڪ��UQE�QVje(�QQ�(�kTU�1b�����F*� ��*���"��UQDA�(��`���(��h��U��V1TAb��QX��A��*#�+UdQR��iV*�EDb~(��HB'��4�jC1�N+��9�.nfǜ�͂;D�iŎݩ��p���N�Z
I<�Ets����k�3�[̢����8��Ň��w+�{8�da��>z�x�	Ƹ�B�<�mIɵ���Ca�l��E0�=��g�cDl ����7���׸M׮n��|�ca\��]�}�NƠu��Փ�8��ףcv����ݹ���]�ϰ�=�2�hcm���M�u�Ƭ�펎�ú�ƍ��F�fMg�mFv�Fs�v.�TF�U��=�+������N��#ۻ��_h\v�޷���n�*��B����3v[��]utO<��8G��^����y'i�d�Y��qA�;uA�klX;	۵��zâ����;l9Q�y7##��<qn�3�+��G���nڷ��Z�ю^�\�mv���Z��I�͸_l{`K�zۮ4��qE��ݛ.��p=*�x�e!k��XKM����yGl��s�n�[c��� ]˱��q�.��.a���WwVSp=p���=m��*G�7����-{F۶��$��s�� }I�D�Q���l�u�ڮmx��h��c�ܻy�e�Vܭ�t��+ݥ�n�[��N��a�p#��+�����n�]gG��Wc���n�]=����/GP�pƹ�v;Xsӷe�Î�^^��3����ԷQ�����ǃ�6�WV�kWi�Z�ݺ��od"�n,muדngt'�iN3Gc���՘�Q=f9*��m��c1c�ջz��-��%n2��ۂ��7c��;W�۳���p�[�NL��qm�L�g�[�Hy���ύk����8�=�<�&�u�-ێ.������.�ې��Y�qwF(n6��츋��Pzy�ӟ@�
��m�������8� ��;b�{[c
���q��|v�v:n�f\�+�����������m��Ӽ���ۢ#�f9��qj&��c'W[�ȜR�"�I1�M���ج��'��˞� b����)۳A�s��)d��գ��w��wKǎ5�&7�*�����N��ɫ���"�g�����e T�\k�%������e�M�=��[�۸
ޢ�W�����`�ۧd8z������<n�۞n�|���<?t�!��;���\�m۵خ�.��Q�ͷb��j�.B9�tSOv����z���a�Wl�v0����m���s�i�2�۶��������ky��st6���z��
ܹ���՘N����!-�%@�����$$F;re���#*��׶}_nd�I$���u�5��ua[�A�8{4a��OĜ��D��'��M���{��c�\V���������$�g��X*���D�^낆�-��f���	��lnP����L ���`���`����O�q�b
v�p��=��I���	$�{�ۿ�?A��Eưߪ��B@-���+���8�I9Y����d�G��P;F�����*�B�?�wP�=}��7d��	�jilm�0Iє��t�.��m���w$�əT�9M��ŞU�	�4ҐLϒ��O�΂� ��:��A��J>�ߖ�X��`}�+�	7���똙~����7]�P#���p7�ѫ���ٓ����7��a�`�{5��D��֮����~۽D���^���<m�$w����t�/p��~��T�m�_� >�|���� ��=��� ��������k��}���7����lO�ț�8#���o�ay������]N����Ĝ�nвO��Q?f�x�n6��7`�����֥ㅂ7Ӳş�$�� �	;�e_����^՚��k?W�]`�xOjP2�F��n�<H$��_�������v	����I;�P2T�����˕6�?���L%jB6�\��;g7u�{]�l`�NyL�gi+���o��TU9'!�8�޻���O��vP���h��v(�������:��R	��Q8ɣ��>��g!��W}u�d�Oد1�$��od�	��)^�['>��wt�12�q�"&v��u�?�̕����t�<�-_ۄ[�yU��9���溤Ef�`θږ��(ـ�C/�M)�'�B_=[�7�ί]"i��I��? >��Vn��{������(~�Ȟ�j��)+�7}�1�&�_�5��I?v�P���^ �����$E]�V]�	������ �չK6nV5(V�b�y�$s{%	?^_uٕy��_�Թ�`���xQ(պ�.4d�f��u�u�s�ۡ[v�9���\`�&JL��3��N#NF�|H$�7%I�.�z�F�#�5{�tA��D��n�r�%��˝�tK�oZ>�=ד�����_P&�;��Ě�^xzq��O�<�$� �q�@�n����?u��,�O���ٛuU���H=�����/;��>����I�"a�f�{��{�Yp�����	;�D�~&vgX�H>��5T����r�������ާa�C�Jovf6%J^��ߨ�و�<�û�=��N�,��J�ۛ�d���~Ie>�f%�]͝���{=�����o�OJ�(|NwD�7PGqI@�~��	#k}({\����5�����_Q3w��O��(�)e}�ky퍹�CX�u�5������=�[�s��06��qa�F���!���j��kx�zP$�gf�����J4j����_OJ���뿉���S������'�S�Y��w��mK͂�'�D�޻$�w��t�f��{�d�'���7[�H�H7���~�� nx`�Y����L�o_�3��#��J�	�R1�ɣ[�<��&K��O[�u��� �Wy� �{{%^:�������{+O�cl�) ��%]��u���2WƟ�T�;��$uM�H�Y�@����w2�r���Fc4�Q�Z�Ej��呌�ʖRK��,����?{����C�K>�/�U�kR������Ǭ����\ ���<w=S�e�3F��  ���%y��h���������wgl=�k#wJ�u{O	���s�d�/\�i썳��7s����d|iHDzYˬGb\s�&���ۺ��)�av{&�GR=K�7r{ۀ��:���m��shup �ny�������xnk/%]�m@�|�ܹ�m<�t�m�:��sc>;�n��5m=c[�eў��SlݷZ��ng[��a��]r��ӗ����.um[�u.�౛1�f�X�)���5>�
E$R~7{� �t���Ă7{'ޛL��{�˰H$yV��#8{؃q����ڱ��{�@<W��}lc+�w}d���<�|F�d�ƅ��7�OCc���'	�?A��J��~���ܺ������߁k���~$��@7M�M�cq�܆��;��	o�DaG;	����(P$��o]��v�_��s#���@��H��&�5��Q&�s�&��}w��6�>���ܧ@�A�̔A��f�X�͒l��°���
�
[m	�06��$��Ҿ�j������gm����1�'���أ����Z��g: �H=���$�M��X�y�|�J�A?��+�}�d,��)��RP5��?�c��Z;�<2b�|�>+��S�ޫ~�S�2BE=��;��l�������{%`�ob� ���<P�<)���w�/�������s_��we
$��������{����,;�tH�� �n#&6�l���}�,׫D�y�����_H;ْ�?�/z��A�|9�BqD�p����(�y�$6t�I$�_u� �W��A����������=Ƌ��-��nCv����7��u��e����m���;��d�1_c��l�c����$O����=�x��仱�s�ς$��N�k�['c�ņ���4�;��^�T��cQ���{e I&�=�d�@�}��7�����<���	��u�siّIE�.Ū�b�v���O��ou�o�/�A��$��@>[����d%U.x���d,��MƤRQ�����'��:��w��d��jt��>��,󅹒�XG���OA=^,7U5��~V-�b]�8rr�YD��w|��;57�v�3�ݶ���}���?3�{�X8o�:�=�8\LFm��z��Gfg��D?���w`�H�y��v{���6ܘ/�e�z����,���5�n�A ���2�mo_`�("���O��07o��O	=	AAx6�	�W�eTu.��h��7X��{t�y�!K�竍��;o����~Μ��M�|-W���I��@�	$v��W�ӝ��{�o�t���ă����*�"������J$I��mf�/L.{�Y��|�1� ���Q������"k=�	˜Sh��$���]���d	+���u�C�T�j�^�Oگ��$�����$�8��I@����$�Ão�AG��� ��e}_o7�hp��{�;}�3q^S��mqj]��r�������S[}�$�oG�����Wøp�9������� �����h����q��17v =/�Q?��m��w���U8��q"'�u�$�s���|o;�W�9���p/���H���r�s�8�l{�n{�[�|c-�t�\n2ì�XCr1��:	�pĊp��ˮ��/���^o������^]z�ou�$�}��"h��Cm�R�>�������_{�a ��m}_o;:쟎e{ޕWG:�����P.�*BP��ɠz�A ��u�$� }������;� ��uh��0�ʷ��Z��z����vob����A�vm������8A�h��zQ n�&�1��2J5սY$7���餮���:8��M�D�N{sn���E9G29НK�E2]�w�|���K��{�v{��^H(b�."��v��[5�kѢ�g0:��Y���wҾ�>��i�����}�����}Y�<�csÁ�Q�}lom��x�b�.��6�zx{j�'z��֕� p��e�;vv�]���찒�/����WB�]ݖ�o<�t����`;n㭆:��#���q��{'�Ǿo��v��H��ͨ�1�rX�]\�.�]�i�nppW烹k�����Ȗ��֛��h��j ���;<�:1x9�\�u��u��n���-��EZj���n��;n;��b��WI�4���ų���������ᰨAB��|_��(�s�6Œ�����Uط�����i�� ԛ>�sٝv	��.� �$�49mS�	��qR���A`�}ݛb�8k�� ��Õa���zk�4���!l��1��X;�޻ �]�W��{����X�g �vm� ��_;]�"�%F���o:U{Ο>�o,�No�lY<�1�o�)Z�g��a"�Vر�ʹ������{�� ���p���Jr���Wc�H�{�|vY�!��U�s���X[��w��hO!���:QŔ�&\n�' 0 �͜�=�$�&8�H�����:�@${}8�T��^y��/.U{�I�y����x���q�cu`�����^���g����{V��2�J91]�}k��n;���H�yd���GA����\O
�zl��P65���+�m�.�أL��~�VY1��Po��y�� ���ݾ��������A'ߗ�PH�^��������GQ�\'�AI�k�[T��{��A��u�,fvg���t	$r�Pf����l��JB���{ӯ-A��vW��\�{-��	�ܨ��R�5�A��r��(�@�� Q�)³�v�����=�+=s��4η_� ���λ'�庺������jk."6��,njml�c��ͺ�7+0IE��e�Й[#��bgZ���|'��� ����<�؁�F�~���6�#|�)��>�L�L�$����kcy��W_ּ��~��Ob�U���$�m�Ew<�mr�ۏ��{Ĝp����+�����b� ���.Ud�y�ߍ�������冹�ӧ��́y��Gu��7�������B>�㘍j��as��馝�9�'.�!�dX�ev#O�}���[9�%���?/8�#K�o'��ڴ����'�����>�i�܏��g{� S9�쉗ؠS)5�t��}�J;'�'6z����)�r�|��>�AK��+�ۨMZ��vX7vC�ҾT��u�Q*�n�wR<����iNeT{��r�T�"�K���y#�Gv�f���@����C�c{���\�N#B���)ܷ�p�v�\�S:�l4����z�ա�xy��rLVM9B�x ��D�ɗ؏1.�3�n�{���7:���<�v��˛����Ӄs}�w�v�C�toVBG�H7޳o��(m�w���sd�Fq�z��qU=��e=x�ǩ�|ǳׯ��E�Ϲ��C����{E�ܷ}�f��}��="�8��W6���$i+8p;<���w�yo�f*�,*��g�u��|�ޑ�a����/���m��K<w Dn��\b �^����b�s�]�P�Xݳ��~���cz:<����uw��c��>&����]��"�=��Z�*U]���尩`�`�eA��z�;P��M��׵������"]�Ww��,�D�ޤJj1ڪ�:^�VN�%�:=��W�63V'�!��b,%)^�#�l��1�G4��ݰ��y�R,l�Y�6��^)�h�0��FU��1zf�u���v��9��8����v!�~uP��cì��,~3_y^s<��3zO?.�X�DEH��D��񨊢�+�U��Q��ڂ)��*�ZTV*�Q��֊��E�E۔�"����PDm�%�QE��b��DUeQ"��H�
�9B���b�IP��U�0b�H�`��V��TTPQ����V*�j�Q"(,ʴb
�R�Q�[mC2V��,EV*�ETX��*�1X�"�`����PQA�����V�kF-�EX�����*���(�A��QUQb
��1��U�0KjV)mb*��
 �eEPUADPTQUQ�&%��QEb��Bҕ(�mȭIQ���U�4(�J�U��BҨ�DF"��0ĬX�Qa�TDzB���?��H;˲� �{�U�OC�O��DS����F˘�ܧ*���mX#���^Q+|��o�uEM��[%4����q�����'����z���)����8�$�{��~��'������y��3|�!��.Ԍ����'lܭq�OK���z4Q�A��
��,~�	�EAl�!<}x��?�gU�G��:����GF�ߒ.�r	��۷���	��$��[�Z��_�aF���-��d�o}�vH>7��y�X��1^-��%����1$�FRM�o�X ��@�II��UK�h�!ޚ�A{۶,<���#4{�p��5�r��y�4Z}w��c���u�����W�;�_
gѼo�����{�,zk��s��=#�Z��衁$Y�|�<����ۖ�y��~���Υ{xEc�{�m����BI'��;�x��O��kZ.����j�|Ho�<�U~ꕼ+�u�ޟ�*�v	���@�$���JdT/~d?y\;uul�:�w�����털�y��1= 3٦ME�&����-��E��w����7������|{��~4��~�]��c�:��	�EHLl�!4v��"�=<5E^���o��ŐO���w��$��y_ J���)j:y��}u�F�Ԑi�H�%ص׮��ݏ)AlL�Gw��|t籁��؍��Q���*0�WƷo��ZoT�Z,�>�tH$���0��oP�\��s��.�8f[��=��bqPP��T���|��?N{ݭ�E>,�C�s�&��`���ќ9=�����R%���S�d4��{f^���V�s�<�~��rd�=���:�]�aR��9v��x$�^s�y��ދ����	,��n�k��ҙ�&+���8��k�<�u۝�Vt�tk<�6��^�.�k�䞞j��u�;h݃u��J�X��MQ�s�����9��Iق�F�&�S����ok�^|�(�cI�4NNUx����{uâ�ܥs���ãB��;2m:9��W;�Cpv��(�����X��,�b�0�Δ�(xWn����u3���.󬗭j���;<��Я�g�l;d��;��sط?6�*2	������D?��h�g�@�M�?jz��k�D�~�u�zO�n�z��Gʻǻ�PD	;�n�l��j�g;���]O�Eu�⟞A?{���םvH(;��ޙ.,�)|ƛ���M��'g=�$�{z��	3
�7���))��ڕ��đ~ׄP7]�V	�?IP�Ļ����yY� z[�@��f��I���}v��g_�v���F8J��$�Y[�,���tͨ��Ϩ��H^���z��b�#˫rsAP������өwY#�ɍ����;G�]y��ȉ%��3�۝�CW�4��#�D�[���(�nm�$��c�eޫ>�?zm�9��	���
��g�Am�(S)�7����QJ���n�6�/+����U��MTkӰq�o�٦e�{E��J�f�?5���A������SL�f�}[�ه<�߹� �{���d���<�V:��Gs5E����[��I�sv`��P7W���z���z�� �3�U���ä�u�݂I���@�)�E9eGy����6i���i�����c7��`?_m�D@��(�.}���U`1�I���1Ļ��^�$�{1�)Z�}�8U���ՀH���@�Oǳ�R��*���-����l8zq����^]��f	�b䓱�s�h�ְ�%ͣ�ڢ!G	M8���{�`�;X�I�s�'�ϓ@~���`�H�Վ�>�� ���"Q9X���G�x�!�|mx{m�q8��,�I>[X蟉;������I{{�߰U�F}$����蟉>�yAs��P�n��n�]��K��c8w�x��M�������H�\�Ы���D�T=KJʾ��wAA�E�JK'@!�0�u~��E��F�ͻ� ��ڬ�zH'�_��'���DI�,v`���w���z���r��@>2��$���Q��u*}�Wy���!�ʽ�Wڨ�t!R�J8����?o���=y���P+����f?��-����{�Jn�!���l�D+���Fr]��M�ޥ5��K���Ʀ���abvxv���I�D�1ľ��΀'�A�Y�����{�Κ�6����csǮ>���'1vP���5	
8
m�$�f���d���[���B�1R���c	${�I��]�E`�}���Q2����W�Ka)8�NEv5��=��I��E��u^���I�]����U�
��g�Aa8(j�o*��[��T��v� �-�͌��aӐvas3ĉ!k��6w����CZ
��-d��E��N�i'�UN��[�M������y'��J��l���y/?��3>�2����W�ɟ/��L�p���:�޻���:��WR��yO�s������Y>]�u���+w�U"�,
*�v�w����g�[���-��Q�.��<k����ߟ���"M%G���U�{��yw��oyXu_��;���������j�I���̪=Z�]h��Rw\���� |��o� �K������=��E��ߙ�{MBDN�28��6��$�;�tI�md~�C��{�`�~��c�����JN$c�]�j�·�W��j���]��?H��D�wWe���ﶪ�w;�v	���$,'��ǉڻ(:�3���O��E�ggU�I�U�:�H=���p*�A\��o�hh��ef䐛�.�tj,w��E�5���9�ǥn/7(��8ir���ז�f��DN7Њ"�{���Ko.�Z׬ϯ�<�UzI	��y�\��/a�xh\Jnm��c��%í`�85�8�:��h�o�9>n��n]�[�8
d�<L�.�%���n���7K��|jF��v�cb87s[�G�lw�`���p*v�ˣm.Wum�X�����ln�n�e��ݹ��u^]v6w]�q����5(/\�C/��J�X���m��m�s�`��l�k]yv�v��gu�\\��9�a��<Qz��ۗ��s]i��E�Y�!̪<�	��}�{�31L.is9�y�����n:$�Oݯ�	/���^�m؞��4��G!0�0�"M%F���L�]�kݵyUՖ~'�ƻI;���`�iovt�����㗽�O��A'��`���v�u� �س|I��:���������]�HL)���I�]^�����P&%��A �.�_�?��ފ��qgc����X�V���ȶ{ ��6V��eڠӽo�$��B����rK��ۘ�ﯳ�}Y�k��&]:;�;�u�9���ǂ�>R�\@�����]�x�R\1@�����#ܷ�u��-_���ˣ���$�w��3'|��i�N��9S�Va�_L���|M��u1Վ?�v���/G��6����.��3%�+e�`�d՚e&ڦ��"i���fl�}��!{���:��?w?{v�_+���f�Ӽ���](��8Ex�0��L�D>]��'�u��/�� ������&���c���]�������?y�$�O#a�f]�~���t�8j���f��_Ē<���^��r��wL燆T1�)G$������Nռ?_�%�]Y$�O�
f�ՀH$yu��7�4�ڂ�2�^��D!Q��f�{v��|`�rI�ƏZK�[�]m;�xO��}�yВ�����+�L�mX'�G���zՔ�X��W�~��۰GY���	�XI�K�B{|u��{9]<� �n�Y$��׎� �ɗ�ȟR��ro�e��!��-��r��ŐG�^1@�z}���Kv�G/��+�}�I2�����f4�����DojQ:]�^îY�F��4(�7�|��T��}�#}~ŘVN����\-����/oV�H���vI>_�y
�P£�2�q3Wo��ϵp�<�_��^: �ڻ^uN����̡cjqH$�2�Z��({e�e�k��b�kf��V��$��y(	;�������{=��mrB�8ɉ��۹:���B�t�.�[Ye�+���.���~���}�3�)G$�=ɕ������!ݗ�p�m��ݻ��yh�Y	!ȜpJ��]�d�OOZU������n{=�u�g�I���J$�����W�ŕΌ��=����Q�Q���D�]�� �>[e����i$��d������)ɿ%XZd����V:�NW�l��Χp�Po�n-�@�����±�ч�\�!��k���P��`b�Z&2o��{}��S'ݽ7/[�^���e�E���B���TCM�	�8M��������\��!_��
�"�Q�k�5~�@�oo?V�<g~�⯁^�D�7�o��;8��0bi���z�7V���{+L���`M`rc�n�f�����I�l0`L��oo%�'qf* ��{��OJ��ITvd�@'㚻(3z<&�>h���6�׽��%U�+�$Cgw	��>%�P�{���^{�vM���Q�ˣ�V�W�-�<[	!�PAv��N.�tIД/�ԝTlnl�]>����n(�-�'2��p.���m-�s�����Vb|��d�=c�G�@]�M� �eR�g1��Xv7��|�R&E',����0}�(���W�S1��=��ɗ b�rl��,�D�>��f�*�����#���Ǜ��+7y���^��J��[�=��yw�q��"�Eh`\xv���%��2mY�)��[�=�'o�{��8s���d�aI	���q��;&��"�Q;��
��_;�-g�b����­L��'�t�_L�Q5��҆H'�X�t��$���#˞u���y�p�{A���\I����9��u8�b�-'�
f<��l�C3���q��zM1����NzK?y*���i�SO.�_Ol��9���7��ݶ�i�s\܃�{z�^u�P��ƞ�칞F5vW�g&4��x�e����LoM�U�[���r��=���&}�Kyغ\^;���|=��g�W�'�|'��1�?Mf�O��A��"�#C1��~Xt��涎�̻7x �zp9����Y��ƽo�-v�p"�;t�>~ػ��M�P�ǽ����Gm�:`�\(�}i�-��v�.��9�����;�4��j�k�Q[�/��Ht`_&�>������T�N��S�M�WDL����CL��p� JBRy7��%>�p�V"�+z���%�ݑ���GG_\e-��Z�B������i��mTu����KBZL�T��Q�^� 5��>���M��z\᧤�͎�wk0��Κ�<zK��iD�Y����U�/\�C����2�c�>T�/W�����a�.��+��:]L�����1�}۵�X���������o���J�b�"wA;:tiI(�{���	,(�4�Y�Z���N�c|�g����Ub�Q��Uwh�s. �A"�TF1H�c��,U�R��*Q�)�b
���V�b1ڈ�,**��b�(���V*�QEUDX����Ar�e,E`���VF()Z������"��TQF"�Lk���
�V��Ƃ��bۙX�����Ċ��Tb�J"�h�1EEX5l�1VV�AQ"���(.P��������LJ����A`�(VQEQE�*����m�Q��X��+Q��(��E.%b��UU�$QE�UE�5V�UGffR�����U(��e��J�W0��\B�"$c�b"��e�S-Z4TQ�QaDA��-U�JնEV0QF�iX���*�*����*��U�m(���s~w5��.i�X^t6I\u�9�0y�*��OZ�'tim�'��|���9+"v���vj�I�4D��zi6	�cz���Y�n��>���?���UÌ�]lu���0?�N̜�F��==����:��e�\�Q��=3��r$cc>{�Z�n���=rqY9�[�o8��l�pYp��;���G=k8����v�::g.P\F����s�5��S���]��Z��n��J�� h�۲k\ױנ9v���f�z�㓫<юOnA��qZ$S���3�tcPft&#u��dݎ��)��{N���t��Ou�y��\m�x}����nol�{whtܺ�m;{v�ݟy�l<]{@&m��d���<�"�p�4�]tWl�c��cuG�-�;�^^{w:�A�t�G6��b��b3�Y|�f���6y��8��s�dgV�q��4õا��������MϬ��5&��v$�C�d�����8̕ي�O�k�w����ޞ`1z��ݶٓ1c��Fō�]���9^4�dgc��9�ӱ�ۉ�vͷ�,��y4\�װ�N�y�"6A��&�U�&{5̜6��v7;6� rF\��x����M��l���ƶ=А=��n@8v#M���ŗ���g\�N��m�=��vlV�S�S�k5���\E�׌�����Q;^��^��Oc�����Ʉ�3�e.��<G;<��[�z�Go
qk��Mmj�I�pi{u�YŎƲ��Q�_e^.R�ہ��Ƶݽuzқ^	��8���NGk�q�\C�]���\���v&-ٺx�Q��ĭx��y�A�瘳��Ԟ��.#�:�ȶ,����U�v[cW]�kW\[�t!�q�{0擅��Z-��l=]��t����&{��ܰ�u�5mێA�e�m��t˦^(����M��b^Թ�Kڛr��F�8�0'n]���*��Ov��kx��v*v�$�s��@��:r]ʓ�9�.�q-O>-����3bug���������9���2۞��t�s�W:���E��v�����'Ap��i�:���,N���:.��p{��k.��L��;s��gx
6�����d5���*�����}��q�Q�Ck%�16-�1ȧm��n�h���2!�.3�N�j����!�}��p�����]W\���T�|<�D�Gaݑ�x3:P�Jt�]T��Z�H���B���\���n�{l�w��<y�m��0eR�A�߆��*8�EG�c��	��M���. 2⺯������$V��`}�Q�ĉ�(Q5�����D�ʠ̾�9���}�� ��d�I ���)*9=Ԙ�*�I׏���n"F��T_��?�H��O��:nR��&OB�nU{C��Y� �=ɸ� ��e_��� �IH�b����+:��Sa|@�� � ŹJ��q��v{G�o�谒�-݀��}��!@TY���w��	n.˹\;��`O�6 nU�D��N�qG�K��:�iPm�RB�e(#Q��v��^@6��^�z������jcv��~���͇��d�A����e��ܫ�dܻp�)�N3܂�b:�;��I �,��u:��%�T��[��b��!�[+�[�;NWsvcҎ�Τ�:�(�˹�/G�Kg����u��\��p�{%�B_?M0���m�~g�f��^3��}����� �� ���n�ߕ��詿�~�#F:�!D�
hn �W��D��n�����>X��z�g��� r7� r�}��֧�#
R6�j�7�[�[O�·��� j�je�79\��'ℓI8}���9<��IP����m���f�Χˍ����%M+ ��f7D�;9[��K�������QH&"m��L&�<�����v�[�-�Ͷ" B�&�EH��Zd��gG����7-0>���$��5hH�"� �;�w�1S)��1����W�ow��a�%��H]3�fZ`�ɰ1I�ky˼�m�7��z��*<��Tq�iP��7m8 <frl� 3��U����U��;�Q���.Ṱma&=��S����Q��Zk�,�+��v������Ȅ���r����W�?m��P�qw�>�>�۽i~�&Cp�n� �����^Pb ے(I�3_���ww������"�Ϡ �-�D�[��� �;]v�8̟f�� tcn��dz/U)��@U$��U��X���'����_�b���3�kL #Wg'32�%��%O�nr�e����� �bBF��i��`W&"�X�o<�;��y�PD�\����ە~9��В�q��J��.�\�5\�>bV�c��nU�TGsqAIyvk��$Y���PH��ֽ�ttn���3ў�<;�t ,�M��v+�fr=��.����V�_*����Vߓ`>�q@����;=��w�$b�jn 	��*:����N;V����/�Y}.�;�\̸��J���X��v�������׮�����d�
a��D�z�:��Dv���Y��tjơ~?SɞG�:�
#ٲ)٘%%=nߗ��}�C'�n�l4��I������%��ϒ'�c���ꋵ�5�%-���Z�7 @��2h$�g<�kMy��%ח��L��6�^&��!���Q���J��z�G���g0p����D���*�Fqj��� Cq\P��,�����JG�������I#�f:��<Y	(A�o��i��=ʟNNd^��  �K�+ s�6�}I���9��}���k��\	Hc�kZ���I!�,m �*��{�{Ù`A��V"($w9�[J�~�J"�r�vNs�����bWܽfú�a`���L����`@�p�*�����ۍ��s�	΀�Tu\"#%��v�%y�l[D�.���$E�'���t��I��x��b������&!rRb���߽�!ĕ
�K��~��~���9����s������^��,*��到������ҡ~y_PN��~��E�rz��Oɤ�ky�cC�k����^|�Ձ���Z}����
4�A�B�mPQ�
p�{$�m��$�T��*�h���m�ٰ����Z���E%�4�f:.w��qk�������ۏml��n����Xݑp������؍a���ֺ�r��MFىw��-!�p�v�O���w\<	���ю;<��;�ЬSu��ެ�c�w��;Z쬽c<��c��xTro�)�ݴ�{;E�0�:�zw�9�.u�Īh��m���jgy���z<v{Jg�ey��}�?|�>.���C�������x���`�C���=��}���Cĕ
�'����a���{�R�����P���37�f�i
����1�c����É��LL=�|~�h�K�n��<1'�c<��q��c0I�s�ߟ����˭�|LM�o�����&!�0�1���w�!�4�Cĕ
����\C���C�1C��|�?:��y�o�<�hB�(����������35�r!�|�saǈm&eI�C}�kǑ�I�Ę�b0����}׼;����1 �:5�c_߳�w�XD����ڇ��������		.����B,��T�+���I����H|��RT+��]�ќCHbb�b�����IP�8�������I0����\�8��RWlǼ�nN&�bd<�����ɚӬ��J���?w�u�r<I��Ę��C�F7�hKC� >k�i��>�x>�_�8k�w�����10C�����<IP��1C��YߨB>�~Z��˻�ۻ�|��,»u�箳�6��E�5��ў�=A�+�GʴnЈ�0#q��?�@g���Aǈi&CfP���u�$��1
���]��I4�	�1��sY���$�+��_�ĕ�&!�?}�u�<b�����N���qא�8������I���f!�����|!��˵����r�ʉ8Qk'TL��r�q^�o��� ��f����f���WE�2���,�!82Ru���*mЎ]�S�v|?��{����!��1�����͡�qa�!�3)����$���+��I�~�~f7_"����4�Ġ����1:�\�ĜN&0�<���x��$�3)1?f~�f������81}�����߼;�/�����C�1����w{C�*�f!�bb{���4���1��z9~Һi.�[P�%L!�4�1Ag�οո���g�����C^��oĘ�f$��Ę��>�f�i<LI��c0q��u���<�b��c^U~�Qx!� 3�W]�D"T+�����i�#�-֮��q�����͚I�+<f!��b����gq!�׃���v}y�_
����0���ohxÐqIP�02�k;��$�n�$�Ę��}��}�q8&�b_vg��*��sb�p~��"�0D_0UǤ�wnP�fW�K	�G�y�벌��HϮy{w���ߦ��ɭ:���J����{���Ę̎$�0�LOs?}�^Rm�b����C��&y�ys�y{���k�uY�3�=����b�f!�dLN�?}�Hx�Cd�~y��k3Y�ĕ
��u�a��I�C�������n�?y��:~�2�̏�bbLL����xi&��&$�`�Lc,���k���2!� 1[�=��;"}]���T@������-i.!"�qא�8�C���٤�����C��C�����3�iLCT~�������*���Uz~W���7���@�}>�(�$�Z�\)?mx��O*�����-�m�n\�s}��xo�)��5� ���@�~Ő�0qI�)�Y��f�x��+�1&8�o���x�!2~;�_���Iى8�La���w�~�ߟ���bOP�*�I��Ϲ�^�C2���!�s���!�18!�bb�0���w�~��Y_���W}�~`����߶���M��2w��?]Q�u���x��C��\�r<CI*&C^�Ϊ>?x��놻͕��o�G�E�ba�Z��$�x&$�*J�q��k�Èp�&!RT.��������!����_hw�g��ċ9"�l�y�vP�g���M�`qSXն!�uX��Kj������� Q��(����G�����C�1}��}���C�1LCa��{�4�T+���t�Y{���w�C�<�sY϶i'���+���f=����8�I10��ӕ�&�kTo�T�c�ߞ���LB��&�Zx���m=���5���&!�0�1�����8�'�11C}�^�x����C�1C?f�}s�=�#�����Q��!z|#�9	a�k7�Î!�;�~�px��fPĘea����Ǒ�I�Ę�	�1�w޳i���7�Oɉ1�I�����ۇ�j��*o������=��o�uM]%єא�8�C���٤����w��g�1f�1���l�8����1�������q�1�!�2e=�w�I��߂�	�`��ؕxd�O"��TX�>E�`�6F��J���V1�6SW��u2�;ó�l�tO�;������Z9�k�>��&��<�g���:������~���'"i&'��4W%t]i����8���7���g#Ę�b���o�����@|Z_��_#[�S�/��@��1s�s~�!�*%B���{�x����c0f!�*{�߶i&���]^��>�~B��k<�Р�EF�2��Y�h�}�s�t��A4k���3�O�e?ߛ�Oں��u5u��T8�����k���bNCfP�w_~�<��Lr3ba��d��b�"����u�}���g�$�{��wp��&!rRb�zo�d>?@e����!!@c�?!�6�����͚O���c%�W�L[��n��@���C�� B�1��c�����!�Cc�bL�Ou��f�i
��FbLa�<��]�}f��WÈ�!2��N�@��o�T�La�����$���LC)1=���5����\b��<��<�?{�{�y��uIP�؆!��>����C��1f3�0LOu��� X"��ߘ��.B`m�~ 3��d{?N���*&������B��P��_��x�$�*J�&$�ɝ��6�HT��$�`��{��!߻����~��B��,<�}�x�0�1����z�du�]MyC��13���ͧ�C��1��c�~��83�i�o��{��y��!�|��0�����ba���CfS?g�m'��bJ�I\����8��|�[��O�J�"��B�s�=n�i��ǥ��˃�ڠ+��R>��S��B�Z{�ܳ��)���>�^�W��aXw��kj�}��:HL���2K(F���nv�^�ۇ�8;.�r\�i�Σ�l�\sΪ�v����6��<�:����c\i�=�9-�S�چw�;���r)���Xǋn�\����ٞA��Z�3��kW:��W"�`9uny6S�[��wWc��*�V�,t�w��I�2��q��M�
E�۞�R2�E��<�m��d���a�u�g �7�sջ6�^�̧��o;6���X�wZ^7�k�c�Ʒ��N�ϗ������>4js?�I�y���x��+9I�d�LK���ͤ�%B�F�9����!�18!�bwy��3������P��s����3��1�3�0LL���ٲ�E�>�C�0@�n;��Cw��À�$�eIߗ��}�i���k�Ck�o����$�*J�&$��;����M'�bLfGb���_ {�̀�2�7w���y������S a�?@e��3DA�"��Ӭ�Ci*^�7�i4�g���$�W���ۇ�b��bJ�a��:w�y��t�Ϸ�w�%B��bL�{�}�i<�ĕ�������<CT��ksc�&]i��J��1��ߞ���m��~�9Rz��b%K��6o�I�3)1q�!�=�_n!�*������2�����=��=�jf3�113��6m��=����q!07#�!�{����Ө!��
���=�_wx�Ę������7�����d|�m��D}DX!�c1Ę�q�~�ۇĕ���7�2�|�������9�^�,E�]�.�ٞ:�u��H�]��NP;>3ƍ��Nݻ)9�F!ۚW�D�����GȖ���6�C�1�3�`�C}��q�CHbb��Xa߷�|�8Ã�~�X��BoT�8��	VU
#��1%q���ǟ���!�*s�ޯ�f��c�Zs<*N!Xoz���$�����8�?k^~�}Z��Fj��2���?�?ڋ6��F�ݥ�Y&�I�L�G妇�Q]ܣ{|�;pg�I���|}�+���|�I���}d�&!�0�1������18!�bb�3�����8�3�c1C���{��x��<��P�>�?f:-`�K��j��8Î!�;�sp�I�(bL�Cw����x3�1
��	�1=;�����=�鴛N	�1
��w���8�$�^��aa�����IP��3�f��֗ZѬ�<Ci�C]�B���u���]�ˀD?i���c1|����3�i%B���c~�߷�x��Xq�1&L�_{�ͤ��'(o�߾�+�3b��k���bJ����ZL�Ӎ��M!Xw��7�x���b����߶m&л�����__�+�h=��|�<~��ۯ|����!���!�������8��Y���!�be��l�	��?<��o~f�#H0����%�b�>����7G;c���+�x�Df��2}~���~t�kj���~�a��1�ߵ݇�i&Ca�1��k��3�1
��	�0��~�G�E�3����_mA-/����?3���nC��1���e���}H��>D}���*?��������&^w�ͧ�x�3�c4a�\����?{Ϧ���y�6z�C�1�w��uq�1%B�ɔk?m
#�#�@D|�	�r����������0��������	v���y��c0q&!RT���o�I��&!�0�1d;�ǟ��J����Q���ք�y���9��Ȳ��=��pu�~}YC��{�9�Њ=��O4���`�K�p�ax8��ײ�=�ݑ��>ب+v�qg�{��%wj���}�����U6��~��8MC��+�4c)�<����LyS��=�a����iOsܴ��[:�D��.��}��N�zf��&���U'��~X=#�dA�X��!|�n���.@�yK�N�	e���V�G��C���8�ҡ.R��_�[i�w}�7z�h����3h~��Dv���"������]�����M�z���#�McP}�OZpu2�.[w����)��~r-�y�~Hi˺��|�w}���/3����XrA�@�Fަc]�s<7���h�N�.��x��[͈�sd8%��0�.�c���_W3}��\��+��1;�yK�;�}��>�Sy��[u����~�:Ƌ�xx{������a�1p���F�X$φ���\IT��3}<��{X�zLf7~ֆ��Ҝ-��R�⋃`�*Y����y,�|���eɊ��U݊�"﯏X.U�9<+�f=M&��pgG�F�Z�z���ՎM�)�:ğ����~J ��%�7�x�ݔ�@qN�M�oN�Iy�ןt��;��e*��b�5K��,��z�em���y���.�C�ޅ,��.��mǏ�NKǰz>�5,a�we�҇����l%|�&|)Y� �#���i�a�&{2͸�fS���E�)�ٽ�����2���}��
�%�QEKj�`��j�Z��"���)`�V �,T
���*+iAH�(��%"��+j�����kF��J�QQQEe�D[kiAEb��j�"("�YAU�-e��AX�*�DDX�dV"e*ơkFKQ"
�E@���Ċ(����b��������2�X�Q6�Z�TH��TW)AE��V�d-��Z6��Ee�+db[U���J��R�V��H���)h�*U-,H��҈ւ"�Dc��[J�A�ұF�U���Դ��ecK�Y�X����%�Q�*V�EZ�����VVP�ETQ�T�)Z����+*��Z�F,(֡QjR���UEXV(�e*���4qV�őV����E[)mmF*#mTUU��Ub���"�)DF`�R��*"(*եD�g��P���&!�c1?}���C��1f�1%K}��@�,����;i�`�J8��?@g߽=@b��&���o�	̀���eI�C{������I�Ę�������i4�&$�*J�q��u���;���|��?k�|���̖��2���� 2���Dd�;�y��g7�i���c1f3���m����~+q������Y`��0��?y�*a���#�bL�g���ͤ��I\f$������������Ty�����C�6��VC8�$��ڮ�N��N��8G�����`5�2)=��q!HY_��� #�Ϊ��:�&3I�a��������I�3)1q�!�{���!�18b������{��^�!�~O|��C�*�f!�bbg�߶m"ma���ZL�@[�߈�<d{?N�=���hGѺ��zo��O�}��H���|�f$��Ę�3�����i<LI��b��u���5I�\���s\?s95��>�r�<s��d_�*���kT�2��������I�+<f!��b�k�g�&!�`��0��=ﳉ��k]�P����1%B�̦w>�f�y����I�3w_nN	���{�W�3Er�֝[ᤜO�]���~��W�z�����}�� ZLC2���}�~Rm�#C��_n!��C��1f	���"��������>��~�r���z�rŬ*�o��f�P���C�pM	�P4�Gm��HOxF�����:�I[���c�.����`��0��f!�`�����C�6�0�����C .Z�+�����t!d��2�0��o���q&?w>�z{|����=M&$�����i4�DĘ̎$�`��~�ۇ�LB��\���y�D�do�f���z��0|
I��g���)�[=�l�wn[q���={a��E��v�t��Ţ=�٤�!@����x�D~C��͛O"C��1��C����q�CHbb��X{�_wx��8�����k����!��/��vm't1%B��3߻��'I13�w��f��]k-|8�HVw^sxϞ$�*J�W���s}U����Я!�"80�1Ý�y!��C1f'����!�pf!�*+�g����"s�B��?1���1E4�5���J�s����<CI*&L��=Ͼ���3�1�bLB���������{�5Ͼ��y��M'�bLB����߿k�ÈsT���LC{����$�W�����u�]�C�pC9���i���y�;��m3�1IP���\���!�0�11a�����$�VqI��g�߶m&ϳYN��~�σ�*%A���u�É�M$���ޯ�f�91����N'�k�;�3��&!RT0�LK�?}�~Rl��~���F��Q�Gā� 2����18b��Y�~׿��!�q��3�b&&{��f��&���ѝ��{�BV���c��S5�A=z?�Ō��_��ͱ�8����3� Df{���E=u�4��EǤm�g�B�}-�R�K�&]6�2i�ƹ�]�����Ѻ���ܛ�28ޮ���oL5����u�m����^���MGR�����b�t����ݶ^x�v/7bSc����]������]Z�0svh�*�0�9�=5;��ɷ3č�[��n�*��n�z�1�%\YuG<v�m�7D��k�&.,�9ݽ[�!�msI�s��p<[��m�N&���g��N���SƠN�:y*b�i��\ΞN,��@��qj���Hj(�Q���qy�����%B��1�s�߷���$�*J������f�i<�~�ڹ�ovW���?x��{�W��|�1���3��߷�8��^o��?	$!��(������
 �c1g����=����OӚ�7��C�1C�1�O�����a��1�8�$�)��~ٴ�B��T��Y�O���
u�_#�!��!���Yq����Yk�ĚN&0����x�c1Ę�IR���f���C2�ĕ
������~�������C��1a����<g�c0f!�bbg�߶mhc�����sF��iu���C��d{?uP��x���~威d}�2�$̡�;�}��$�bLB�������I�*J�I�������Ä	���#�ۺ>d�����fS x�b�{��:̗Zi�u��i'��g��6�mIP����<��W���c"��'�������)��!�*&L�;�ͤ�n�$�3b���{���Ę���9����<?mx�DB����8Kd��E�m�l���qי����v��`Ip�ۈ��9�Nk���a�6��+�^{�gG�1��LB��g�o�I�1%B��W���{��T� 2;����_K�������VW�@�8�C��C����߶mh3��kz!p	De����Y�~�7�x�I�(bK����;�;�l��}�_���r��rѸUh�ˍ�\�u���z�ҮIU<��&�]�wM%ƻ.��C�%�5{j���5�7߹矃y��x�3�1���Ę�g�����i<LI��c1����{�ᔘ��LC?y��s�/���ߙ�� q"3�~$��#.DU|,�dJ�����~�mf�1%B������qC�1%B���7�����5���Xtqa�!�3)�Ͼٴ�M�ĕ�bLq���{�É�Ę���e�Q��EG4,��!���~�g�gS����b%CfRb_3���M!|��1��9w߼�B�"�# ����̯ߩ�<~�	�?3R_��~�C���CȘ���͛C��������7#1ȯ�~,�����A��I�Pę2�0��}���q&?��+[�Trt��>�4�G̅������Ę�q&3w߷�q
��yI�f���x�F�>��������;�}wӍ�D.tWl*X��]����������G���	�%���Ø���(Fd����C9�wf��6�$�T�
�������&!�bb�=�}�Ő�~Y��ߟ���_x����hdu��$��I\�1
�����<NDĘ�����h���.�;4���c~�;�g#Ę�I�}���^��|���S��{�\�����80�1������q
�C��C�����g�c0f!�\��ǝ�ۃ���;�9ݚC��1�s߳>�����]c��q�1�y��!RT*Nea����׌�LB����1>������|�ty�y�<���ZyԅЧ�ޣ���}7�b�j����0����o�U��=�����O>;��	��u���}��<浬��j���I�蘓�+0q�����8e&!RT.X{��;��0������$!�ˑ,��ˡi�S7�{2^xHF��~�~d�f!����p�
��11a��wP�CT*L�O���f�n���f�~�ǿ|I_ј�f?��w�q8&$��s���]b���U��M!Xw}�7P�%B��|e&'���f���{���]�q%B�����!�*p�11C�?{���C��3�c1C��Y߶ihcu���������m�,&R��m&
�2���ֻ��-�C��]/0a�y��.�������?8��N�kW�����?����8<Cd��2�0�߷�׃8��*`����؄}������?p�=����C������!RT/)1a�~�wP�%B�>�<>�W�M5��y!����u�f��4�3#1g�{�;����?!��w��|3�b�11a���y�*a�������٤��I_�1�����ֹ=|�^�p�>��1?}����R�4��O�1�?s�c28�ɔ�����f�
M",� 3�}�{Ɣꮥ���C�*|!�bb�3�����8��1�3�11>�u��!�M!�L���6��ˢ����u@~������߻������&���0���w}�x�$�*J�bw;��i&'��1�8������<B�~����?軜�vOdK_����x�����T�Ku}�坃����>�7��BΡw�5J��;�|�|����>����zO��LC0���u<a�2�p���F\���x�d|���*��؆��c1f3����Gq N��,�@�!��9�~�@�����Ca��]��4��T1%pf$����{�q8�I����'��]�~)�5җ��r�u�K3-˸_o<��"�@Z}���^���=`�۾~~~'���Ɩs�ԚN�0�ϼ�u�x��*e&'��_lׅ&�ĕ
������C��C��{����;ך}!�k{�u�b�f!�`����f��Hc�y���Z.j�毜CL88�?�����x��C}���_;��z��w��7_�gc���b}����$��LI�T�
���P�r��Rb~���~�w_C�k{�H	�p�t?1!H���/���z��lC
Aa矽���*T
%`_~򿾿o����c�o�X~��1�8�$��~��4��T1%B����~����10�ܯ��k�M|4��Vo����]o��g{�w��ƿ��l�I�d�LM�5��x�C2�ĕ
��=�p�Nb��Y�{��<~9�^�a�k�O��}�?C�C�19��ݚC�M!�3�v~�IK��ʺ�^i0�����A�x�T*J�a�u����q&<�}�'}����I=B����}�I19c1Ę�q���P�$�^Rb��wx�� "�ǟ~�!��Wu���d/G�G)�?ф��YQ$�>�a^��3�[6�6��+N�F^�G_M�A�h�G\�_b-VG-�dH8�	B�Bv�Cv�:v�����V�LcF�m�ɋl���ܞ|����	�87kO�;a�8cD[n ��lӬ�6�i-M��pu�I�ކ��Òu� ����6���6��g����06�2n
��u���o�|�|"ޗ���Vz�	�K��1p��k��Hq����W@�t�1��onL�i'��܁�ɷo���I�p�n�C��шy��S��^8�k�>�La>g�臻\����F��v�I"�xoq2@�2+���#����{�6i<�if�1��C�����qC�1������@g�!��r��+�5{dG�4&�}٤�n�$�T�
�~���q1>d:�cV�h�����#��~��)������d|�Y·��l����m5��l�ғhfJLCa�c����q
�C��C{�}��3�dGȀ���?�3��G�����6�0��u�u�nt���CL8���oaǈbL2�$̡�=�_wx�G̳�#�@D|��U�9��IeO�.��NH����1�8�����8e&!rRb�������8�0�1���L�"EA �� x�#���<����������?3��c1��<����	�bJ�a������J@G���������~����:���^��C�*%x�}�op�%N��kHۅM|4���La�7���px��*2��g�khg���_w�_=��T+�C����%B��1���wx��b�f 2>Dk�� X"��:V�ߏ�o1�������4�1D
Q)
*B[L��o�����s�]m�v�X:��vW^���������hH]�IP���7���1&eI�C}����!�J�b}�߶i&��+5�5��h��Ԛf��s��8�IP��&!�=Ͼ���8y�n����Q������@dtyt!mIP���~�9�����&�W�lvז(u�_<��v����+�	cGܷPm~c���p�6o��3�^y��U���n�+�������fQ���g�3�bJ�IP�3�����C�88�0��1&e>�w�I��bJ�f$Þ��K�z�\��ɯW|ON�W�H�!��"���8�*dq�B����!���כ�8�&3b����w��)6�#�@E�~�ɩ��[����W^知��u
��CC������gb��P�1>�w�C���1||p�ʊ'����Ő���@Uv�Y����Ys��d}�� &g?}�<gc�Ę�&$��g�i&��+<c0q���{��_�����������'�^�b�����<a�c�5�Zk1.�[tk�hx������I4�gј�3b��{��g�	߷���@���ɾۄ�!�0qI�S�g�l�O�ĕ�3c������N&$��s�����s��~�TI�$B�l@�F4#�t�6�u+�\�l��)l6?@S��$�_��#���$AM$�;s^w���<I�T��I����lג�hbJ�IP�{�{��%B����|��믃��D�_~���f!��b�&'���l�M!Xx;(n�H�.<GȀ���T�#��@2>��w�z0?�v��Lpf$��1&&{�~��I4�	�1
��}����8e&!r�̟���z�_�0��do�}��>M�7Y[�x���C��|٤�!�1�3�`�C������!�*" #�3n����2��_g���l�|����2d;���9�U=7�8ǈ$hTa��82^�f��)AuI�{�F�F"�u�7�:aN�����Hzñ�1�!�2e=�}��$�t1%B��3{��NDĘ�y�f�L��9�d}Dx�~?g�����?z��ew��̏���G̀�2#}������9b���<��*8!�c0Ou����8˭��^�ߟg�q���b&'u��f�i
�ϲ�/i0��~ 3��dwuW��T�2�$�(cs��ޞ�Ls��<�\��<���2>d?�L��#�E�c28��;�w�x���.Rb?�uB�� 3Y�3ߠw�E*<q����$sۧɷJX+J���Tv7N�omq�q��e's( ������Q�1�
 i�bg3��6�mf�1��C{�����!�*LCa�w��b`�d~z���iFV$G��~~����I\f$�cϽ�{��bLN��xkJ���٤�!Xy�w��|<I���LC��<?\�s3��Iy����Rm�b����y�8�N!�b`�!��=���x�T+8~d@��;O)�6��#�?�B���{�e�Q1�$�������]T�Ca�1%B�����x�3�1��Ġ���U{����}�3�~G�:	�1�I��8��{��*���>���Ǽ��_J��%ۀ��_�f<��٨J�ޙA���� @-�ڮ�I$N.���g�ݲ���_�2�g�g���~偭4�R >�V�]dYy��]�2gʛu�Y�����;�N7��<��s�f��*��uM{�,�$�[���ɖ�G�&�l8��pഀH���(Dխ�y�#4(��-�}H�s^�	�X�%Eӽ�<���|����Q���v�y;[woWnڞw�ɏe]҇Xw;ct�D"!#7'��Jh�
���r�3�]�d�����B�^��w%�<�z�'��t�U��!DQPTEC.�V�c$�=����:|:�m[��� �:�F��"ʺ$�<��w9�_;��؝��'�T�/�f�6:���Iչ*"W�-ǇE�7+�|�'3f�H�qvJ����P1���QlZ�u��I��.	�2��mcC ��;)L��|=��^�7��og�{2p����^B�UD�$v�O]\P} }���s��-�fD���� � �r�(���\����]Q�J���AeY��IL4;�y?{�å�L�_�*w��~6���S������˼��K��;�-��!��]1�V]�=(�;y�X�&0�P�y�u��Uy�1��Ĳ��6.��ۖ�f�y�HH}�@W���s��5��ՠ��6��4�:=�!�v�=�In�yZ5��h��Q{=��#a�m;��0QϪ<�))���=�F����1ݾ���:	��|3��Nx?yLx��{��$�bZ4�IY�I�/]W��2��7B$���tw-ྯ�k���:����%���޷T"�:�9�!�jQ���V�����^g������.����\
��'��`�;����@򙻝f��\k���ѧ��Ӗ�}]�:��zN�����n�����Ւ;��N����+�b�����֯wC&��&w�|���
����묾W��5O�d{�L�N��y�^�C(Fs\T�۷���mn嚽q[��w �+��E�k�u^W�X��}���M���{�n���1 #�ݬ�~�Y�lx���>9OoR�?��C�^8ޮ�/���߿^b�+`�ϩe�d��Œ[��^���8����+�s�՛�rK!'��8�wA��}2PNh��x��"1��ɱÄ�_����� �>���b��s�b(���j|���k�3O���fY᦯Q�	���`s�3�^o��H���_2�F΍J�iӒ��i�C�!�%��/{���տ4*��u��	�qg��5�]g�חǔ�U���j��RU����TQKh��TR0ER��#V�F
��
���m(��ĕ��Kkm�����T~���\��m(�m���Z���ե[ZZ���V�kD�V�B��D��ҕ�֬R����

[Tm("�JT1�YdRV�hQV�T���**�ҩh����m�KAe������V����UPƢ!�UcX����j��RT���X--[+m�����T��Tm�[J ���R�Z�",-��*��B�(6ѭ�b%ie�R�
m�h,�H�"0Z�+YZƴ
���`fZ�bc&U����Z�Ȍ+eZګ���dkTX4jZh�K����j赺4�H׮�@�].s=�nC\�s��S�뙺�u���s֝)����Y�9�ۛ`�4�Nu*Y��pf�q��lK�kvm�^�^��ݻrcN����7Zs�Ohlp�A'V`�<��Z	Ζ'qS��Z#�9��9��x:��v�-���!�|�~O:7llU�p������-���3����m`��N�x,����c��>���gۃ���:7ob���ڪ--\����wc|W9��׷�j�3F:Ǉ Gd��y�x1���!x8�Z�.D��n��ڐ��ܽ]��m��������	�v���^�U��ϙ���#���ۉ��n�d�c
��)���*��ApWK�-���`������ɝ�;Rn3�v�s�O	Gn@-Z�n��<�D�;S�n�'F=�]ڳ�I�p�H\<s���@�zƌ�\�@���i�q�y{p����g��]]�\]�Kpⶅ��H��I�mmƃrv���2���+����0
qm�esƃ�f�mn�1��OZ���=�V��㸸FU6�nDh��m��K�lu�z����e��@�F�Ӷ�st�ӝ�xh�vu�,a�w�w�m�R�ܪ��{��',UB�U�'�pk�������p�s�=��X.�F��7�g��<Ů�*��>|���ˮÄ��ڹ���۶Bz�zX�LO3ԛ�d����r��!��pl|�|�.�Mu#EAm��>���7�+�9�&�gW�ێ�<ƥ����U8��x����pk==[����]���k�x� �5Z�M���kq�����<j�7�飓�Pz���ȺN�:��"��[g����;k�8�;���B/@Gl��t���ػ^��/C�y{K�g�bێm�eg�0�l��vKs#G]vnyѷ��.:vyM���
r����ግn�s����b=�u���gg&L֖�>k�w�8��\����6�''ZnĤU<7a���[�:�g����n�'[.�+Dn�=���v�;Z;]�㧍���0�����z�5o[��}�7 ��)غ��.ø{�wc�L:�c�]����N�P{[�(x5�������8�wcU���mM	�t�]�k5��7mō�F�����o`O.���i�x��p\r��N��< �!�<�6;k0v{#=K�ru&z��Ƿon\[��9;5v�v�ԫ��O���:���*��A!�Kv�p���9Y�ds
WE852�Ow~��0�q��?�Y��6�>7)L̀���q颧f�Ol7�]>	��ʺ.tpT��P���X�3�k��l��/���e��=uks�2A���� @�˛D�=1N�>z��r�u�"�IE7�3����\� ��U��aШک�m2� �r�(�=�\��-�H ��ƍ��yVW�v������6�( g�X������;���Hm������.�O���*QP�Cp�m�.�M�N��^No��Ut��\�&d���v�b�X��|g��a�(��`�񝴭��mvywn:�Õ�N�L����8���g����{�F8�h��m\�"_$No�R��l��`6��7����=Wb �.m��YT�aT"�Tӷ*�'���5p��|]wF�m��/;g�;n����A��0z����p*|�R���3��T�� d��{���'7l�Qp��E��Lo��c��:��>;լp^�M����5=�yf5y6+4uXP�&�4��՚��=��C =��z]��g��s}J���>7�X�$���rn��R���P��	Z풃�����($�]�󆈀�#���`|vU[�T=��� .��h;��j�Q1Q4��Z�8a ��-ďm�DU\�y�^'c 8�� #�]5h�2�J�����>.$�ϡ���Ay7M;��ۀ�-tH��d��L6KH�,��;��cT!Q��m� ��۩� �"1.��͵��{��B޷�a�J���I|'}���1ģE]XZ�:$�'cܹ��W.W�� ����8�L�@'歷z���Os�A~~Sj��U�4����ɰ	�b�	n=���ߝ�y���^�E�q��VM��uƹ�ΗV��h�ݧ��'|�3�Y^ͻ�M�Y�N��:�Sy�6�S��Jw��SԺ.?�$�0��l&Cخ�K�%*��P��c��ժ���YE�����6 BHk}��H�o�Y���bf�t���T�Ne�pLҩ���E9��X"I$��}`[�=������!�K�d�Ik]��M/w�Z>��k,3�M��jzn�ek�4�ySqm�d�Ә���<�֝��٢!2%�H�j=�JL3���;�Ij[��@$O�ϩ}{sF�gYvr�VۢI�Ʒ|"_~9� R�!T7 ��8�����ɵ�������0 �,Į � ��sp�A.�|k<n���HW|�t1�R$w<��@L�ych� 4�Mv�}���/o�3>�qD� D�.�i|+o�ӈ�j"�W�X�����{�6�܍wo���S {}\ə��{�Ηkտ�npm����c����<�۝�Mӣߥ�2~����}�͚���j���k�����ܡ��}�X;/ON7r?/I�L���>�Ȝ�xxd�T%
�J��3���H����:K�Y~��� &H��.d�ϗ{�jU޷ك%�x41L�%&�3�5�B��n����`������ X)�A��e��w�)���ME��|4g%7��sh �.�M���/=�v����w��BIz���� ;)�
��͚Syc&Z��aͩY{�m)��kՖ8�>�>����L��-R�s��%:ק2(��H�T���ݭ4 vjpɐ
g�]Z�'~�]��& y��� [���/�L�r��(��Gs��b�MK��5�ff�,m�j���X��L{픤������"����BD\R��Z����D�.�Q��;�~π�}X� @噩� 'C��#���x���� �*Po����幷��M��� ]�\��|��+�&I=���yֆ6t��4���7�U��Gg]y�m�7}�j�v����Z��<��Z��s�qc�/7f�7��+v����Wø3�l;�gOc�;+=GV[rx�bm���[vN.Ey�l4��۷�,��ap+��c����\��z����s�wK%�u��5=���ꃭ��3���5��̷���N�jW1����s-��n˲���e��{h덮�s�7q���N{`t[v�,�����͸�c�h�nyye�7^��wnz���	[p����*+�����"܉��è��y��d�3963�ؔ�������M\X'��&�"O���V�6�n�U�&��H�cGj�
νmo�M�r-[f@L���S`@��)���0㜒E�jU�� ���܅��cf��n���_�⸠� �4�����=;|����V�)k]��\�fB�nˀ�I�wk�Q�ѾwxNK��/y\� Ļ� ��D����L�,�g�-}\��I
���k�p�H��r=j�(� 5���>gv���w�i ��d�I�v6I'�ϫ j�z�.�u�;��D��A�A�4QN"H�9@�a��1�ljv��6�S��� v����}xy.W����C����( �{\��V�ӗ/M������_�A��V>�TqZ-�*(�6�%��n�;篳�;��&�9�����}������:��6���m��]��i��M�$n$=�%홹跲�y��7B]�F�|z�mt0 K1+��|��D��7��_�f�7`����O*
����E7F꿨 ��.p� |�[�������� b;���"|��A�N�RD��5IKcZ�j誻�p�xs7� ���fd�{�������z�\,9?G���v���%*�J��R�w��`���S�f߾�Wz�m�s����R��� ��M�����۟Y�|{ͮ��=r��k<�Gg����|�ݰ��\����:jюnba$�_�`'��K�(�Em~�c^�����M�@����G>��~x��"��Z7���m7 Es���QD�T혫�� �܉��=jmm��.����#_u�p$y{y7 V�x�{p���YA��:2R�&�h��Y3��Z��O� @\F�_.�AG�v/�#(�9I0e#;/b�9La{����V,Ƶ�`чE��Z�,^oP�צ��`R,�z�Y��X��@?m6|����������QM��ڥW�=&ns��=�8` �٩��Gb���+I'�I��Y6��S�d��EPM%-�k���|���S��k�w�ϳTU~�. W�� ��u��qo�P�b����#p"ۅZx�G'g�ƽd^�n,i�#�n�W����~}w���	UP�*�'3uN�|� =ڮX����R�/,���Ԝ۔���^�M�Тg�	�T�$v�G�]���^v���+U7�;
� 1�qD��y���n�@��Ɋ�QE�S�*�&� b� "3��&ny�������Gc���ۅ�I��-Z[��6��皥Q� =��&O��[�L�>�}��e��Z������/9r�Z�!�����8��x�Yŵ0�V.��ko\v5��]Ρӻ��/� w�E���"����Znk۩����QB(��՟Q2D~�2ꚜ�os'*��ح�L�r;��ޫp���!g��8I6'����?!+s�{[�x�9ޝ�2[]�O�!�RB�R��V�P������p�=M� ��&H��n_��_�n�[[�%�q ���(#���$�68��J�X��J!^��я���E>[ &Hĳ���t�M����e���BVg������a3U@*�GnG�]���l>��/s�o#-o��ygA��WR�ޗa$���1��.�,r�ubȒj���u @ �WA �nX���븩��R�Ѣ������P�	28ū.��b�)//v��t��{t��^�]xī�X @߶��$�/w'3w*�k��R^~q��*ǟcܹ�>e�N�r{=���q�jq���>��!�{=hS�r�n�E��_/y���=�Y�o\����v8�]��6��ω�eױ4��vn�s��\�r�x�S�.ݶ������ݕzw��Ζ�zi2g���T�g�@c����oo\\�,�%q�\ �C��#sd�ˤ�ę���utW�� �:m�A��3lku�Sru[������[p�ɶ|p�H���v�\I�8�m��O8���ō���|#(���;9�;i�l��::�O��jW�m�t��!����Wr�.v�Adf��1)!E1QL����B%� ߶�0 ���ɰv�ڳR��k�v6M|��ܕa.�EM(@��RSn����;]���G��bS��?e�`�w+p #r%�tJ���m�m��=��MN;���c� |{98`��v5���U��2|c�Sa'�����.��MU*����r=j`�;Ǫe{��u�i� g+p ��*��ξ³cI�>^��d��p(�LDc1ʞZ��-  x;�z��Ң��[��A������V��Gb�1l^�;dJ�9��J�mc׎�j۳��n:L���q���A�"�����Q5	2Hǟ ��v]��x�j0 4;��.��T��z���Aw~��@#W��aZ�\PR�`QEU�v���+���������� f{?͙�8�oy��a�!����9y��et"�p�7g�E�M���➾R󲛠E
�ײ�vu�T@������Ӳ��GE�+��W�u{^�;��QP
*PRR�oy8a@O�tL��`t�i�.���Ϡ "<���� ;*��Q�ؐI��p��+���z�'Me���]7�gy\̰ ��J��<��Û��[�A$;�;&��Ǌ{�F�˫KW�P� �	e�K�eJ�=��s��l^�Ne�㲔́��,�S�웳:�X�e��r!�7N��S[�ѓ�s��r��m5��
7l��E}}l�
"(̓'|��s�I%�G�rTD��ޔI]��������w��M��2P�j��m��p�$�[��;e�h���4tǧi[0*�\� 'M�V��U��O�E�ӹ\�ib��|�PS0(��)�f�\P ���� }��k���J׉���6Y��Rn��G��X�>�G���׮�����x�A�ި��:��x����DwO{����I
�����A�h��v����F\ˮ�r�������N�#���8����:��_Jgz9�F�R�oxY�ݻ'{ܣ3G�ZF�ϗj��q ����ӁZr?F�@�������ۼ^8r9s��r���]Z;��O��k$�W���<V,j.�n��ڲX�n��B������Ʒ�O�H��}���ҧ�盌�0G�c����O6�;�f��+��=�WY�iu�h��|.��gB�Sq��v sQ�YG'����V��4�9��>f�T�:���&OiY췢y7M�N���`��:	��~�1����˸,�ʼ+=��D�K#O
� w��E^������fOڲ����6~��4�$�H�~n��ɮ�^xn�W�z��֚���.�o�6���_:F��Ӭ͉��@�Y.�ӽd��윃&:v򖹐��̓4��y>K|gk��x�T��RicQ8hզ`�ډJʼ3�����tf�s�q�"49�}�������hF*Og�]�VI�����/Rۗ؄B�|Vb�|���_J6�\cs\&�6e��N՝��y�<�^sdT2�*O�G%1��D���f���6�!!>��F��Ν��u�N1��׺m�l'2Z���b�ɴ�B�]�s��A�Mt�z�*��#�����tv�H�{F��3Q�4,3��C�k�I��Q桇ĶP%Y�RԬ��kIce��R����B�+l�D�X"-�-���le����k
[��Ԫ[V �h�E�ekm,�Qe-*���U�V�UE�J�-PmX�F�V5�iJZ���U�m�[e-mkm��mU%J1EYF�*��l5im��e(���iikڣe��F*�h(U�J��P��ض*T���R���k(�*6֌*,Z$*-��aF�A�J��UJ���m�Z�m�ZYT�Jֶ)X�mb�UZ��"�[e+Am��B�Uj,��J֪�ƔYYF"��j�j�1���F��[[IQ��KQA�P�J�Ɣ�
V*�X�eZ�֪
*�bZ���X��V�l�ֱk(�)kP��Ҩ��UX��Rգ6�Q�Q+
4��*�#m��ҢU�P�� �d&��׺ 	�7*�<���HnQJ��LB����o������M3<wR�� ��, ��ʞvX����'V��D��{aE'p�$T���Sa @a������[4���{ �t����}�o��-�N�`�g8p5��I���&2L���	���������K�ۚv8��g���ߝ��S��$�&i�@x�қ�{�r��.�M��x�:Y1�����vU� u�˰�}�D( Q�%3��<��w�J���jy�$9ҙ��>o�ܸ �����{�o�=Ҿ���'�D�;	nn��� �٩� �}�Z٨�y���J� ��6|G��'2���q@UL���(������t��<"0� V�)�	�˳Sp L��Y\�ӹ>�2�ӫ~�^���[����b�Y���{��+ �kV�~�*�x�/�)���􋷼s��w�[�cѱjVx�Q�嘡����lι�&�E RR��]�N@<nR���T?sJfMݫ� ՙɸ �]��9���e|XĜQGfT��dծ���Y�J�O4n�Zy�h����?l`T��Q"���i�� ��3�� j�a�tO]��{��n@#g;����<�D�m�I�,%��(�6<;~.���η��N�V��>]��E$xe�K����ީ�n �C޸(�**
TU4���S��㲔�.���̷[�s�$b����|�KWd����i8DR&)��fvĵ(]�v{��^����@q��r� ��J�  �ާ��N@��l��S%!(��˴�vʉ �	]����Yl�7�W�3�K����'�@���Q$ cަ��g\�Z�GEc�~�Lf�]ʫ��ߨ�[�{�!�57�h�y�R��D,�f����=]��l;�K?H�
�ȔRd9K����L�5޲E�Z(��%"C�#P�b��z�S��N����x�m!����;XL��T��b ��n6��^�&3��R�g�Bxqq����ۮ@��qkk�x�afSkF�q�$*�vb�g�n��zg��S��r�n��Q������<�@lnݧZ^���+�q�n2	�%��7�얍���Yb[���!��Ov��˹C�g����{��6R8N�F���V��h��]�q�D�L܅]i�N�&��m�g֋C|�}�����zi)ٱ��a �WL�c�,�����%ꉹKɳ��o	 ���j�Փ�$*�P�$T��w}M���
�g��~Ɗ�^d��jܥp N>�@1Ov�.��j3wZހ>Y
1eMP�R)L�:f�֮� }�� g��<K_�צf|y���PI��.�I�~�b!A�G-N�u�;):�j Ħf����̸���*��ʕ��iO`.k)�Vh�e8DN&)���4ZI ��f���\*�Ի� �	 .�+��Vĳ�J�d��vIk�D6�?'^�]!7����.Ƌq�қOq�0���󓜿>��_ΌUBSU4��9_�o�N 7ܭ��Po�e#���" ���Wi.�*��8La�v�ێ���HB3�C�`�0>}�c��{��=Z/��3��;�������=���@$�y�2�S�Um�ݚ����(����tgB6�yܔӡa���6$�	/��-��"<�ܛ� */c��Z���A���$�HP�%*M���l> 0�s�$���zp�h��v�<	$�^��	����_� �</��1�e�=u͢5t��Y�)�ӆ��}ɰgNʟ�:jo՛�� v��n=�
���R�3��W, ��tCO�6'}ykah�[��w�Y$�Z�Ң�ցw$���ƥ��ɣ&��\�Սα�w���LgH�]5�-$�eܚI�ލ�*
p��Lk���h���N�j�R��e�e������]�gϚo	 �{X���-1!p˰���Q ��������r���s&@�=�������$�'����/_�ީ(��i��p��f�5ۉ�ɓ��7*��&�3�Hr7T��H��ґuvg�I�U^o�dӊ���m���L9�'�-��ʾ]5���f�b�1u��+����zY'�ݯh� @i�Jo�϶���!B���6艹����"��� >�˲���A~���9���J=-�C�=����֖�P�&\�z�≓���O�n�;��lUe�R�TI6���ɠ���J$KC�g_`5s������L#d$�$�|�D��ɣ$V�S+l�nj8��p�LE&H��"H( Q��/:�0����qD��W377Y��8*���@8L6�D�x�t!�)��P���fv�a�]�fu�\g�.�qs� A��J�d��z���@qx�SB�r���|�>J��Ќ�	�
��`�ڸ� >��� ��z��c��  �2�(���ަ��(�{$0�1���
�v.,�w��syL��	Ү�� 1�-ˈ�=՜=���N��3}��o!U�H����8�^�<{����c?s�A�ۤ�oo�ıUzd����mS9�������w�ӗ=��.�(1d�jI)R*�J�p�S` a���)X��k>� |r�� ��p]���dH�ׯ��0�1/�!�d�"+�������Q�vVՒ�\�N��A�V��`2}�w���F"$͟����I|�^�a#'�]��	�ί$m��%��8{*� �^e6�p�q@AQPR�T����l��X�u�����>	�#�u�`��V��9��O
�&̒�kh�5G�RQ8��a-��F�Iyv뿾d�쌫�ێ[>=E��r[ޫ`$W�%��v���&�
�����i���Lʵ�
�Q�}y� {�ӈa �u6!��D�����	S,v�I*�r�%�3�@�.l����p�| pn%)UB���9۾�r� 7kto� �Gb��B���	����7�N�7U����a�ۯk����;�ܓs�\��_�C�����(�0�t�h��#��H��ͽ��v;�-��ˡ���
���Ô�ܩ�[���2ˊz���j���rP�V{��p�.73s��j�9M+θ8y^ms�6�1�(x�]�ܼ�v6�Zَ�ܮ��\�-�;��3�X^`v�Z��Z�t//\�[����Y�ɮ9w��ۃqe�v���9�8`|��-ٸ�֗�j��A��������Nx6<�K���;�D�q�k:��*O\k�x����n5�L��!���_��35t,��L8q_��S���r��5/ؕ�8���VW��7��l$3u\���0�`� c]���: ��U�ws�F��Z���L�.�M���\E|�����06�Ω�tz���E��UT���WcN!���WA�**��r!\����� ����L�j]��H4+arD\QH��`%��*�ׂ&ˀ (�������������s�Wo��xm�`TWs���R��[]��Iw�k�
/���w���e}��ɸ ��WD� �u]���[��ӽ����- ��㷭��y��.-��&�-��F�s��ݷ�p}}}����&Bd	�w���;��I.Kq� @�[��+���GXtW��=���7  y���7}�B��!ERC��0��~��뭔�{)�z�(�S��R�r%ksw@�3:�*��{�$n��.���l=Z��N�C����?;)�A᷊iLm��W<��ؕ� @��6��+|�j씢�}o5)�SG�����L�Wo�L������Z�K��w��]�0 ��WI }}��_[����B*�*c1{���+���	�^t?o� �=�S ��mˀ ����]E�M�8�,�Q })�������1r���� <v�p�Y~�uc�^.���[F�����O��-�M�{�%w��N{�¸6�#���b	Nෳ׷V�J�Ƹ/l��9�$��1��}�*)�b��V��@��i� ��s�pｷ�{��_%P@��l2�q(!)B�Sv�W+���4s^^�� @}��79[����6�Dì��\G�.�t��-�#N+��]t�`$��M��4�����{Q�y{;7U�������B�P�[�k��y��=�����"�L���:�z&l�w M,4�Y.ר��^e6@���$�b��0��]�	_:��u2/=��B	���q @�572|�y����ŝ.i%�*�]����]I(��E*J��N�8��ObʸQ��=�0���K�%�ݫ6�	!�3�� �eZ5�T�o/�j�i�@B��$Fݧ��q�[N��c�g��;�cR<$q��i_�C|p�R&=8�۲��LϹf���ue%�S��or�u�]w	�ә��n�p�w��(��͈$�]���W� �w[3��M�p=�̺� @��6 ܲ���#��ng<��I.�H�p���No�x��,�l&Pr�n3=y�wד��Y�`�q�W��j�*8[�F�VL��=X�c��g�c	ڳ�`��)_�2|z���t<ehJ_�l�^�swI2��u��3h�^ʭ�G��W�*z�W�mה�vx:���tɼǽ#�����=���u�ד"��k����Q93�FIw	5�z�I��%��6�_�̸�h�X>̫�@^�6���-��z5/�L�\nBHq�К+�Mֈ���
� ��絍��֒�[���������MT �Ea�:�.\| L�eT�z����=UU{�P�ͥ�v��耙>	�ʿ�'i�^�*�QB�CN3��0�y�蚊kmz̆ ەV$��n@ܬ][=�Һ�cZ{�.�m2�f|؁�eXH�l��I�����3�{��ka��� N�UL����� ����HU@��C��j;3e=W�334�� _���a%������_.�c��"NL��X�*�%(��j���-��a3�����ny�
�hvUL�@_�]��%{�r�w��8�D+R/��/p�@����d����>��1��k��2L@������q� q`>�s�/{=���R�V{�a�㧺Q/u>~	=�xj����y̐�iVv@���u�сa�zZ��t<2��-��:�����/w��� %(^z�;PԀ�^��,m�$ֿ���˾3-��"���SW�{�^g*^`Q*:�w�����������g\��Ľ��4C���7�)��/w6}˶�F[D�
 �h�Ⳡbg9�>�V=	=��y۷&w�j+�M�7�9�ag�%u55���Oʅ�);u[nX=�v���L�=f�QL=Fv����q[z��,�����]޵�	)�f{2���Z��[�_Sw���:����]AgS�r�T�g��cf�E��F˃�s���7�[R�[_t�Nfyek��j�;MC�ڷJ�S���D�x65��`ɷ��^�.��国  �i�Z�S�V��κ� �~�y s�I	�[�7�]�������͏gv}:T�,{������-�A��*]�+��ٳ�'VI�,L�����Ѻ^�5v���1��B�o�����I]:�s�h��Ą����p�JZNwu�>^�4�<jMLx���x�rMg�-o5���\����V��g./�����]k޽ a��۰]Cȥ�F��f�*ɻ��/�
x?A�	�����+�D�c	�Q��D
V8{+	://?%�;�=��{=�;,�ck˷�c�,y��� m����TE*�ыh�R��h�j[A��YU)lZ��-B�Q����FZ�D��e[E�JաJ�X��ѕ��Qj��,YZ�VQmXѬD��R�Kl��j%�Tmb[R��
֊������Z-��m�2���J�,D�h�kQ�����j��Q�[[jTZ[�-*�F�b-j�YmF�h1UB��QJմ��ȤP��J���-kQ��+Q�`��
4�KV
R�JZ�J,b#-�ZTE�cK
�)l)l��aUE-��4X������"�ZUQ�
ш-VJ*�V1���(�R���**�V��[J�ڠ�k[[)j�m��(�AUjڶ��Z-X�X��1�UJQ���T
��[[-YX�Z�-�J�UR�hʖ���UT��*Pj[`�R6�b�bJ)U�YYR�TF����+m�m+Z5-��
�QZ�ڊJ�A���kB���E�=���N��fk5����4q�&+�smu��nՇȐ�^�z\[@4ü�ƛOL��[muuH݃��
S��v��m@���h����Og�9n���p���99ֵ�����˛F�'Wd�{pl���+�k�=�6�z��#�&w<�`�XvY6^8��ې븹�K��Y�hR6ݑq����SB۵�]�+��۵��	�Sm�=�ru=���m�Z���l�
!F��dC��ƌmNr��L�6�Sm<�����������j	��e��!K�nO;E��X���F�n{ms/3oc\�îOokj�|' G]u��Uۛ���O0�l\'s���ϵT�:�"vN^������ؗ�m�{57%��Z�}�����i���^89!�ws�;Tu������̴u�C�7�CQ����nr����[1�Y��]��],�l�����kc��V�ڋ�維���	�=�;qv��9���^����bx�ɻQ�Wj����$併�ۃnf�;ePcyf�@�g�!.�<Nu�c%�t������Q�����Z������0\�h�0�ur�Q�eg*1��|���Ύy�؄;}���v�8�N9�����A�FضѸ���\����,��Ŝr�=L\<��=2m�L[�[E�&�l��=vx�F����F�Y�C�il����(��-ڧk��k�8�]&�qm0�5�MC�m�1�ؐ꺤�F�8��*�[ڋ�`�z���y����Qۭ�ݭ�Iʄ;��E�i��⨸o]R۴�{
���s�v�:�e�;�f�'\���z-.����\�v����;\��M۠�bMU��M�x���z����R����v0���xNnݦ��w.&�u��nyۡzvՐ��i	�ݖ;-������8+�\�.�&5��/k�͵����y��yy�{��<�1�kO�[�u��=yS�F7*6��[��{]�k]`sŻmhd�S<�v�64�������r��[�Ri뜯 ��vU�l��Vn�v�G/�g���风�ym�Ʒ�]��<q��9��.�Wu��z튦x93ׅk�n۸�y��n�t$�N�ad..s�8��;�Fw*�v.۫n0o7(��=��������4c[�f3)=d}���ժ��M�X���p��]]qۮۖd���<���V�\�l��:�s��N����x����=�S��=c\q#Ƹ72�)�`&ɱ8��{nu�2�n�����t=�m��8]�v��<�jO�b2K���J��A,��a�@ G����	᷻�н3�XJ��� '�*o	?/�(:BX4�z��W��
ܨ�{�g�u�`@���̈́��g+$�_g�����}�ĵ:dK��l�H�9,%��,H$O�f�| jյ<�����nכ�33���nH=��7��ޚ��%5�(��e�\�a�<3H�3�K佹��  �Y��p q�S��l�k��`����d�T*�*�Hl}]�` Nrʸ�d�V�b3^��S;�ܸ �v���  7�U�+s�54��*�C�/���(�24�(��-<�{\���"U�ܺ$H^���Ny�����be�JU��j��b�._�@�e~�U���p���e�6Df�qw�O�"��	�1!Դ�Υ4��K�2�#j���^��㱸"|2����W�&��4wXb{���ع
'�t��R�x�Mvw|�<O�ݪ٢ݏ2�Oc����g~q>�c�_�t0� �r�F� �L�Gt9��9�U%�bHN<bQjC%���,�J>�p��:��b^��˗ ���� ye\"jD�P��UB���nv�z�&}��&�  �VQp=�n���\�O�ʙ�"�����]lȘ�F nw�S^��W~�Z̊X�Ǟ�ݻ/��][�I'9�cE��ޗiUP5+�nx"����,�Ŵ���>�q�U�-�����,��F�mQ>�ZS�!n@��K���i$�:fU�| y�U����?,�����.�Ne�nU�@s�TR�����RP�[���'�-(�������yv-�@���H?.W�ȋ=���O�q݄�}�,��$F�dp�W'�B ���N!�@��.yu_���U�_i�Ag&%��nW*�7���p�y�U��&n5��Cۙó�	�׵���}�]��㼂�R}����'Ǘ'�|��Q y�S`}\��"&�����c����z��O�"Z�$M%5\P@��r�����g�����d�V׼��..G�n��D��{;+X@�S�[�[d�2g��#R����d�5�S���[ڛ�	{��Z�7������C��y��ANf����f�ܖۇf�i�{4Qp0�a��-���b}��e�H�W |���� �{S��Jj���f�7U� O�e\˃��'B܁5f�_<��o��l�����W @y�����[ڜ�I_�~��R�t"K�ClI$Q�Can��\ gjl ����Qy;��OeI8	��_u9�p�������c��$F�dr�5�~��z\��=�|�2d�7S`|A��Fw�Ȑ8��j}@#�7E^��o���휽���^�o�+Ӻ�G��v�B뢭+�E��yo:�X}�7�,ǋ�����<��8ţ��u����oA|��ɻ���ݿM��Q<%h�Ц��!r��]o-$�^K��x����\�`�<�3,Y����Gb���yVA$�Vg;1%3��)���@��1�܍��.wK���b�uS��>]��������Ȩ�Ll�{el%�ۮ���+[�n�N�7���s�7��t�I��7S`}u��4��P�M9Aڳ� #���˫�oYլ� �[�� 5��T�JY�r�Ts��Aݔ��՜Xj̅9j�+}�v-/�'��t"��"���˷� �y��ɫ�U�`$u.��׫!�6$�(ʊ�*w��vz+#/i�����J��%��ҽԢ��s���M���+|�"6c ����S�	$�����-����S��v+�`A��WD��S����/A{���Ԃ�F�U�b!�)=�2-��$����=~غp��ypG�K��1㰜��A�1�ְN���_������Q��FD��6�Ek:�&�:뷷[�]bgq)�nS�^mۃFݹ!:��
񄜃W�`󓚮i�O��P���#��g�Won�����LݸH�ۗUq��N�+��\y�n%�L�	��ru�ڑg
��y�m�l�I��t���؃��v�PI�Nx����Nvw��?7B�ٰ3�㍵�Hg2=�{u���xl����rI�=G�ϗ��]ɳs�U�q��`�ۛ����E<�z�Fa��GB�(!��/��=�v�� ���tI"U�uY����3(x��w[�p$u-�Qg�9E�b���3��d�on@M urϘ@ y,Ħn]�J$�����Q6u{����t�i�AAP*��J�.�&[����!b���#�	 ��T"$���D�S;I��)"0٥��S�����+E��0 @�1�'	9�0� �����|8��_$�n�CK�ClI!���Uz�$�׶��L���e����	��9z�J���}�5&0בGW��!��Gl"|�v���T�o\�:�5d�۩��C'�����n�N��~#��  9��� ����C��vwZb���� �Xˋ$�x���
�*=%5EM%Lf+|�0'Κk����I=��U�M�W������ȹWQ��vO-�8ת��uݝ;<#.R�c��i&u�Q��6�>��q��6�DΏ� ��yX� ^�VM�z�{����Z��EB$\^GdqF�4��s<�~�JK�ݮ�/�':zԔ㺌~�hެ�� ��rl�V�,@�P'�
ڽ��]�l�S1� 5��� @y{y6 N��oW���z�M��7 }�����٘	ER$��j[��r� ���WD�3�x�y�>���`@���� D��tm�'�Qw1U:zW�* ��^[�a�;� v�V���϶u�8��xs��O���Oꔩ(�UI/��&� ����� ԿbW��^���^X�ș��]��>ұ��DF�dR�5�u�3�1��{xSOivCS3<{�[� ����DPK��_i�r���UT�T�%L��0	�bSp=U�|�ŮU�=A�)q�;�]���0s�s���b�H��q�۝�ra���ǃ�s	ۃC���.�h&=Ԉݘ$�F��a�N�/��߳������`@j;��Tq>�TR�T(i����j�{�7���2�p� �#�J�d1��/����ګ!���(�m�7����6X���J�oࣶ��� ��j,^�]{�yoy6 �e)�	ǫ��.�����u��Q��)����
�6�rk��P�zẔ�7m�g��_���d�EH`�Ɩ�Z@$�G�d�"A%���\�=��j��՞���@�rW�o���lD�5XJ�TT"��8�VE`�O�^��>;)X�u�"H�����%r�=��7'�VHQ�����XK��P���]q��o̙͋]���2@a�UA$�]H��ŉ��>��^c��;�b����ױu� ��] <[e� �ܯճ�]�V��Շb���$\���D��]�V�[��oʮ����V�\w�O9�$9�FsB��z\�����㟵9�a������xݕŋT�%	q(��ig�P�Jc�W:��)�oW�rfp��p�m�$������^�V�gK�)���>[�5�����F����s�8��'&7k�5��ck.��ޅ�،£.9��%䯢P��r����Oy6�C�tװ�(H��˺�s�$%H��V ���׌��?�ޜ��	�r !�֯� �rn 
�(�޵
��q�Y�/�q��H�7%Gj�DH����� �u���}���Խ� |x�U_%j��XI=Ҳ�P4
�"�a.^�.�z�W	+|'yRH%�2�C$���`�eM|����w(�jhIxΪ �In}�����` O�ʿ�ѵ�=��xG��`�S6'�M����������Z�"��u�!�7wC��]���aO+PJ�ox��5���ы�ްqk�-�J9K��3��X�-S�|up���W6Z�t�
�p�sΊN�+�;\�5�pn�v̓����
���\ 㝻��d�#��ڍ�y*�uu�����CرtO3cM5�3O=qڸ�wK�m5��cqh��'$%�93D��5�����c0�7/���֝��ŞQ��� vc5�����ۮ��k�nV�y�|�d�s�ܸ|S�=�Z�O[<nI5��냲v��K���� gq���xB�q�v���@_D�L���T�$ q(�������� D��O���.��㏵�ftȊIy�c�IO]>�тq˿���P�%Y͵J��}Y����@ F'��� �㲮(��!���pxI�����b%��Z����In���0��x̫�<��ǭ��ì]�`5>����e)�-�ZPD�E�P�K�|Εu�� ����2d	ò��L�Ou�/x��-��ٰ!��M�vL��R)��Dbj��;y�X؊����g�l�a������Y� ���>
C�����kO�L��IjC�9��t�'<�Tys1Mn�Ǜ����n�G��W������@|�m�5�'�AӞ��Hջf|�ӄ%n!�ձD��̠����EH�LU�v�ҁ��v��Xq��3`�}����"U�s�v_ 9��RN?Ks���_�z�N��O���5�S)�1�����L����߽��~yf*���^�
��8�����W΀$=t�&p�\n7(Էh3� ��ТA�-J��:瀐G�nS��T?Onx��q�A.����3��uq�~9�2������r��m^�o�٪��$��m ��e��I�"����}��΁˼������H�}j�$6�*� �j��3�A˹�J)��6:�J�xM�l��7�p�n�zn7�z�9v�۳���[��aE_^^��^m
�@�}�Wo-[�4�:�ۥ�*�`�H��U��H�s�5�W:'�納�sWu0A#/�B�$Z��D�|����C��J�N,�R&�� bb��{�
7��	�����0U[�uy��]�~�\�zG9M���g�rz��ʊ�%)����z��L���1��u�y�  ��f+I�a�If>��72@E�[�
¶��X���8]�tU.�&E#r���>��G{l�4N�{�O�}!=��KUI�+�d���ˮ��{�l�m�(��P�cƳf�m�j�)Q|V���F��=w���P��n{UVJɝ���0x��w����(�f-��N�\��0�<�,�:�C�f�����p�M�A�f��١����>/#�`�޽����ǽE�{ygJ�����I9�{aw)���x������:�u���Ң]�0T�N�,�����R��{W+�֠8=�mg|F
V|#x�ݏ�D����uvi�-����o�ѝ�%(���0Żc;Á?��
I�d>}�Jr�pbW�S��[�y�~�Y�^E�<(th�X�)������]�aػ.�d:O��F�V�}=3}�}�8v�VS�� �!t�o���x�Fe�X�_�'"{��n��f����
l���o=1����r��{���w��4�/��֫�"bmm{6�~%��̯*����~lL�$�~��1#h�jd�݋Fޞa��^4�<�3��Z^��X�V�cj��ݽpQN%=܀f�/��ū{�O	1g����DW��!�s�4��'�����N}���v��l`F�oX���zD}��[�ڎ��G53�&ɛ�l�����A�#�z{�ȸ������^��w�\߶�ۂ��,Q�B�,��QX���Ub0Fej1iA-V��Ь���E*UV"�ڣYT�lD�*
1U�R��Eb�
"Ĕ�eJ$�[K6�ҴEkVJ�kU-���h,PE,�����Z��+"ʕ�Tk)e,BڌZ��������V�����Z���X(�+H����cl�hT�m� ��j�j%�V(1AF����ETU��VV��b�V(����* �V��"�bZQ�����TU-,U�A������E��"
��EQj�֢E�´����!mZ�+E[h���
���U�*Tʔb21m�V)X��
VV,��Q�(���*��DH�"
�KJ)��AUDUT�X�*+�F"�,DT��"�J�e�H��* �4J��jUQATUEb���DU����,V*���R�QQEg�����H'�ʢI7}҇ćn��2�F���.�%���vH;��I#o6P'�Nr��qY&���jt�u��E�
C!���vJ�o�b�6��޾���ω��U;y��?sWe^��t�ҹ̎m|�ْ6�pC#g�'�vMs���{H0���p�ƅ�8������߮]26����ڪ$�G_�W��I9��z�b��u���<A=��_�
��Tm�DEVk���d�m�w�՞��Q�/�����)��m�P!�g��]�h$�=@�$m��N�W:��A�.����.�q�/�yV���X$Z�kH9vẂN+�a��$@����+�/M�*Z�2�� 	��b�H$z�������+	�OJߴ6 �Ӳ/Vj�V+r��������E'9�`˞9�=���k�ɸ ������@����+���Ԗ���+���1�ИqDbq��Kuﶀ�1��]n���|G�A<������L}{�D���U��%$rDȉ�"k�kÓ붖x��]2�:@�]�q���߿� %'���tH�՘��O�z����W��C�8�׀�~=師Y�[)��1��^uU�ޭ�~��L` �=�(�={�(��dK^�,�|�cW��l8�"*�ט'/:�� �����E��w� S�s����� ���$�7>I�C�M��7k}/Q'�NB�'�����֯��ߖv/@O�EާNk�al�AF���~$7�ő<_�}�������;}�D�m^�|�5�W���$:��l����;�~���bu���?_WVa%���Iy+}�(�
?(桋���(B��6�����0�g��o.���A���܆$���S��j�8�� N��>8׵1���w0�N���qUgsуi���� K��u�jtiz�˝�qFŵ�q͋\���u��:��g�mع�z5Ӱ���v�,���QP�e���l���[^͗��=�����p�7d�|�]sc����h�y.N�y�f�E�޷l�u����u�o^�;�Z���M��wn�o-��uv�󡂛��c��8��'&n6��n��粼�_�_n�Ê#�F�|}k:�$_{e|I�{��o=w��mw`5k*�3}�+�px$SRT�Cts��|w7�|&����+�(��yU� 7��-��=���a��k#Wx�-�ґQ{�B�o��{o+����혷�I��P ھ�@���^b*0�h��u+��*��>{v�����2���:���|	��0yg���~���x=�H�s��u�@oe|�ƥ<���2��"veP$�+�b��.���o�����)<=�A�Mn:%�ͷ^����sϒ�>��l-vNkF v�&H#Q��=f��l�|s��@����~�>�=�ێ�ա�i�~��0�+�tH�t�&�(�r7(�.���p���N��'7�Xܞ���e
v���s�T��k.:/�k�c��wmꬥ���� Luo0�h�_w,t�z��(����1`͙�w�m�$y_k��?��B��N�NE��g���|/JA�H7���� �{�N��YG;]W�{|$�^믈'|�(mo�4�L$L�\�D�1�)eo��ǥ1@�ڻ|OČ��Vz�q�>WcȖ�<蟟��������;���Q�n��s�s�5�c���i��� ���)�	�;�U�<��쭮�	��ɞs��W�w==n����-b��棷j���=xd���3�rH�s�jz�	�ŹL�I��U��f=}����?wVe2#�|M�P�ٻ}ޡ@���'y��_1��O��1P�Nwz�N�a{��7��1z<$st�&�(�m�+��v�����
$�w=�Эiz�����;z�����	H�MY��_��g��z}f��~������x�"����zߓY�'�fFx"�'�ۋ+�lQ��{�`p�s�����&�>	Ԇ!���h�֦5^ӊ|A�[t�'w�T	'�W��Ϭa�o^�$՘����6�m���#�^����?>��@��=	n�P$w;:�1~���\������θ���<搜֮���ՃO	��6���\T<=+�Ӕ��Dn�4KI��k�oM�G��Z�� �پ�������΁�[�ܭ>���^��g{��\2�rH�s�5O[�gg���{��H&�}�d/u:$٬�=ݪ�f��yo���~��lǚP+t6,�����ـ����sۙۛ�i7��]�	^�t}.E�J)q�/9��T!��Z=Y�G������N�${�X�����,z�;�hS�]�L�*��~�ʓ�ͫv,���x�|�z�mx����'���������O��ʻ�}:����ի={��s��t����	��А@��g�|O���Ǖ������ݳ���Ml�]�@���D�{��U�ͭW�K�#��m��z���+��[v��\nm��;n��4�I���fo6�m���#���b�?>�t���醀<�vQѤ{��3�:VݐF[�B���!I�`,B��_��"{���T�{�Tw׀X$���@�N��R�~>���;w�}@�$-��Nk){�A �yH�O�\6lB�������O�n�
��<4#�>
&�a�hح���V��h��U/yW��I�醁?���4����`���B��^E�.q�/y�I ��������~<Z�'��*�OǳR�ݎ/��(ٟ�Sn�׋��4g,��U��F�ۑf��Ǥ��{�y��v6�f��`����<󾩼r_����1�m�;�س�]Z=�Cu��wnD��b�1W]�[0�!��/��s��8נ	��[n��&��LfM���>|���Y����\��\�I��,a�t7V�nc���i]�;�TKqr���|Ə<8�⺲dۨ��"Wr;E���=�/I����c�j���Gkl�6�:;���< Ǘy�:�r�,�gݓy����7n������P�=�k��ƴ��q�!��"���l��l�������-%��<i�)�b���ڨ�{��$�7{����ë���vTO��I�ǔ���m�L����I�Y9�,[WW��ԩV+�	9�����N�v]�x�x��o��Vdՠ����Ж�0!wgo������nX�	K�.w���ε�Z$^��@�H��˰{�d�mO�pVǖ��u����'�Ω~&�{.�$G���6/'��'��H��PG����1��nF�7g���,�|}\��+Q�~>�� Hw�Ɓ$��s��<}\���F�Y�f���J���n��v�k۵�N�;�g.������Wj�g������6F���Z�3 ����^WȂA��ʲA#��Έ��}WaY��DW�s�*�<���l(!NC]��1@�/w�����M����m�:��|O�L���"1����{݂Oa��ϔ�l�5���>Ww�k��2�@8��Mɓ��t�\&ŗӞ&Q�j�U�G���ܻ$���\蓻zG;|Ǯ�����~[���d�mH轝�,��Վ���p�n�>}�����Oݙ�vA����V���&2��]��w<E�ĞQ��6O�VW}�z��ĂA�s�sn����3�D}�vH�ڟ6�O)�$��yI�p�!�״	���	�S��Oǽ��OH�N���iqj�nNY�9\�QA�{��F�k��j��c{[�8�����r(��N�W���x�k�I=�xk�G����,�>���~'�������\2F\24�^s����u���c��^_ �F)�tH$�<"�z��<�˺��t7�{^E��PB��+��^sH7�� ��s:Q�2��}�� ��Ł�Ѓ�w�tf`���x�s�:��=��b��IєI;�����ܼru�s��G�*;��'�R���G)�u�����{��6�d�mH辝�ci:��y	>35��H�t�@����m�ԸټP8}9�7G�3�Li��k��h��۶/�����%	�x�
/����s��ovՀkv����2���Pa� �'s��Ըָ�2��v�j�v��l�B+͋O�����-In2�pY��~����۰b����nC���k�H'㽯
yOB1ȠNF�7g}ז�����-��Q�Y[Ez� H$���h�~��m���ž6+iXL?o?9��0䑨�i�(�צ� �gm���lT[n��6K礒o3%'�wvݒ1�&�AO�q���g;w�s��.V�E�gX�G��<ñ��^Q�G]�	f��8\�u����|�ا�k��~�7����������:�����YXso�je��	�Bŕƴ�~��wV.�}mk��8�*Q�k�I��2DR@��e�	K�:���&��x'u
$~��A>O��պT��AG�Fa)&�@�MI N��kӌ8���3��5�m�	�2DF�PG�������5�zP$~9��b��<�����[}8yҾ �Oٛ�w�'��q�jHq�ӃO�?�����~�'D{�+�T�$�@�nu�$~O����/c�K��L&�)�"��m�w��vz���_��Ēz��M;����?ٙ�����=�RH�R%!���W��*�뾚?�~���OĎO1�$��vA�Sx��7�*��D�v��H;֓m�gѸ7v���đ�̃f՝]���y���O<�O�=���$���$ I?� �$���$ I,	!I���$����$��	!I��IO�$ I?���$��	!I�`IO�$�	%�$ I<�IO�H@��B��@�$����$�P$�	'�@�BBu$Hz��$���
�2��Oo9(��� ���9�>���ր*� � � 5�AA@
��J�P*�@h  iEV����B�E&�m@)��� k��)w�J�A%  ( SF@*�IlP(�J�$���@ 4�( � �T*�hQ ���R��      @                             �          T#z�ڕ��N�ڎ]K��t�PI�Wm[f� �aIswa����Z�Ԫ6�m�r%S6�i��J d   ��
��9��]�� �U:]ή�W;�\�Xv�fˬ�R�p 9�+���b��ԧ}ܗ�zj��u���
���TT�   w�� @   P ^�R����c��N��t�jU��ʒ�. u*�́�wJ�l�6n��C���jUzT� w�6S�g�wM ��)O�  ��/�*��nf�v֮ :�R�Q�׶�wP�{r�mJ�͜��5��� ��yg1��9�<�zt�zE��]S(%A  ��  �        �%6]p�Zk��ʇ-:2S����p ,�nM�;S���������7 ��w3q���L J���  ���}�h��Mn ��@��ӈ�s��K;�ƫi� �@��wj��6D����0w� ^�^Q%:�
�  �    �   /�>�����@����y� {�/0 �S����= ��÷�(F��y`)�a�)�m�:��x � ��'E���:
^�R�'{� _�͇���<�(
��x 
;��hP�8x����j��M�s�P�� M
�vJ�(B�(>  =�       �^���i���� 'u��àWMS�Q ����G$�N���: ���lT��� ��)�   v*��Ҩ)s4�K�� �Ur��vj�ӛS������i��.���� ��Ue�:d�jP�j��H���D����CE)" �"������hL�"~�U(mIH  �~�M)P  ��JT�Ph  ����`<Oǿ�G��֜t�G��z���#����~hB� ]�����%I@$$~$�	/�H@���$�	&	�xw��?n����\T~�$˜X1'yjL���"ޝ�uЫ��heJ�e����X�Ee� �Tu:�05kjڂU���ui���0�V#3W��GB��f�˄��Տh���&n��2��u&.a�P�HYW��k)^j�eT*2r�#z�N�հ�T)B[�v��[[H���7c�8��C!�l��Yp|�PQ��P�����a�r�un=���B�m�
ܬq�����f
���It*�N�ۭ��:l�͙ Ԫ����,��$v���	9zK�� ����8�E]l�b�w��5���	�������[��w�j�sS�=z��U�XY 쏦ꔄ:�-Uܛ�Y�m��X�KL���u��2�Wf�z�wf��y A��d���҆n��2�<j쩼Ǒ�sLT��@���Ќh��	�f㹢�e�N�����X%6�-GS�[v�o[�������Aڱw��S)�2�Y�s
T�t]ӱqi&��n�ݼ���Ȓa����q<�wy�WH�U�o3%�&e�t��au����v��: òP�o��U�X��*nҘ3)�R�
��
3qija�0$QW`qQG�6Ƈl��^,�N�y��iȈ�&�M���Y�>S;
�g�5{%������7@Y`�Ib�Ai�,a�:��xr�I�c]��朕�l�ڐb+(��Զ)-��Z�O�Wug5��qXL�՚3s�-"6B32�V��J����1��{�݋U�62\
�n�D�:r����:�+yU��h�ȐM�)U�n�ҢR��jZ�
`��kUm-�-f`����Ib�[+l�q$㰃������+F�U0k�s
srЎ�XUr�6��U�A�Q�����r�}�b\@w��d-66�b;/NJ�@ܚdQ]�p5�[k]9����)�O^U����m���t&���M��-fb�[r;5�*ٺ#�5��f�a���(p֣.���T:�1�����%��Nic;q������7�RM��;9��c���7wOq헔�=a��e@j�cz죒5y��Qz�V:v7r�a۴L��U��;o.��.=��Ţ��/Z��R��ol����wD�`A����GSl,U���gإn��=���,nR.�<�wi�4��9�m��������3U`�P�3U6�k76�Nc�b\(�A�cn��=r��f���;DJ������9�)�O�=������^Y�(�FY�`)�rK�[r͗bn���j�{Vu�lV)V�%h�v�1�jĠ�2�<�n��F�.���٣h[��S�z*��P_jI�J��Uw�om8)��q�֥sz�5���jV�(H����_+�ͥoVEF��K��xNPc���M�M
�4�Ws��
����S�b�LJ#�<N��H[�1����ظY{vI�݂m�MPx>͐����>,���Z��Ej��+l#�ƀ
����k�Q��F��Q� Lz�۫Т���;Z5���v�@���EGk%̼(CYT�"������Q����ݫHZ��	b2Q��e<�����4nYܢ�'pj!�+�а�Ȱ��U�F�켛��j�(J�kvz�*T*|֡���1�fa�3oc��[Fh�߮m7��z���a��thr-Uҩ"S��u�7�T���:^�.K�v�vµ"��)��7T���+�����p��!Z޿�t�[��v���p�FL��l���N!��ö�AB��?�fZY��ॿl.⼊�2��F��x�<O2l�2)c)V,yv@��O��X�c˓Iۑ)үS ĉ�g$չ
L;�F���65;ݷ�j���307U�Y1jҳ%���sA��{�!�(Z���V�7r���ĒbU��L�q\�mc9�j��7�Z*h7�n�\��k���4��K.Du+r!�O(7T�o�G�5A�#/��*�wegd{V��8E��-"LjX��#VS�䣹tS�)���y�K+E2ތ���ZutTa��&λ�V`x��Z����V�z��
yj,�T�b�[����V��e�Sw.]��l��u`6(�Y�I�&g+u'��Rw�Xm\j��;h�+iD��Y���B�k�+Ы��ln�S�T�fa�Lb�{��k��/v2̗��jPc,��!!1y%�n	^�A�d<sa)	�2�b.�]����){Z�S��:�S.�YV�Y!l��jF42e�!XyF�cyi�TѸu6�U�\n�t�7Ne:o,�%ej��PЩ��!Z���y��,���N�ޖm�W,Wj�ة,{Fd��~�s1�SZ����Ic;ǈ���,�P��8�HS�E���K�˛0���5jqX�O��ͥ*s-���HC*\�1��p�)	&B��"�*���٘�2�w&���jd��
�72R��%pw6�&V�&��ɔV��x�o2�ݬ֥�ٺ�bV��33,� 6]D�ݻ�ib�h�Ū���r�3V+G'��DͣV�sIͧfe��M�W)��?��ص�Y��l=)x����Zw��@Xs2��5�X7.RF<Ǒ;Y�fh��ȅ�v�*f�����!K��r;�7�q�a�;qش���h�ܲ�<�m�j�f��V�]�Av�R�ܻdPI���e���y1ɸ��ѧ��|�����9����-8f��U��MY,��8�+5�0JH[ȋ"�PY��lӐK��rE3�������2�/�̻X\ڃ`ч`	�i=�T(�雉�y�3�n��%�j�}��,[��v��n6�j��&�Pl�bAtVJۀk�\6� �f �N�n]��W9(5qT�S��c(S�����HMc2�ٺ�7z��	gD"Z�-e�]��f���;���Ҳ��6�[Lvfev�ڌ�n�[b���\��U�wg�W6q ��jH7*(��s7�A��D�K�G��\��c[gVV*Ճocչ&E��ŷ�w+*�VV9n<e⑀��r�B4)��1+
��/�J�,� b�S��r���)B٬�
-^���(4�Ԯu/&����ڭ�V/)Ҧ7,]%�����[ll���u��2Ͱ2A��3�X�l]��H.m�6&��bp(Vd�:��4Z[#'�Z�4��2U��n��C�I�W6᨜�.�FD��~:ָ�JKkJ]2(⩈�R��wԙn�"2�͔j^�Ȱ�,ҫ��	 U��Ab�ot^�l(lTWN�nv�v}2�k�[�Uᷬ���W�T�9�P�E�7�=2F;951Ic�m���8*jW�'&+"�C0�,G.�ͺ�[�kqgɜ�1�̫���b��-���������,e蹭�hVØ ����!t�eԙE9"����
���e��P���Mi-PE^Ļ�X�t$���+5ba̬�L�L'Ov��uޫ+ԳAƘ���+�3� j�n��J�coUm��cq��6��@S*��%�Q���ka�%�0?�W��f�˻�Z��e�yF3��7nfc[j��ުl��.*Ց��G�Cn�̀�ׂ��3F�����qVЬ�w 4v���B^]���B8bd�93v 4꟔���	��>��f^8v���6��[׻�KSz%��%���&n�Kmm�:0Ҩ�j�0�2��fmj�(��N���!�ka8�qcO�xm��'��Y�=Ia��s[EMm]�yR��x�hQ˺x¦��FRA�0��6�	i��{���j໶��6Xc
�KYT�����ֵ*�]Յ��q��`.;�F&�qb!ǀnX���n� \u{���yW��S�f����'JEf�.�=j[S|]&�A����P����ɬ��u%v"�mne�;J=ٴUȓ�5{R��TA.��b��1���F���t�����̔n�qc�,�:zt�F�e�:���O
����iֽ�� T�桻M�7���G�1����X=����l	�]��<��+ӡ<��/6���)=�GM��Z���\�h� n�:�=ݜ�G�2�5��J�^��Y���`+d�+o$��gs~�U�p�.e-����FS���%5��)Ե�EM�o��GJhH	�MCGr�dG~�Izq���n왴�R9�;�m�ӻ4��H��Q*��f�%V6@� @�����1]7l����{��2���3�b�:���Rf�74�r�0oE���5��CO5��X�-S)nQҞ�����U�(&�X�ٴ*�:�d��q��0���)��&�ŹXnaa�rŦ�8ִ��B�+C�n���P� �1D�v�w*�f�5�`*vx�/�E.n�3�/��x˛ڙ��3Zb�\��7���,A�r�]D�sMħ����]��ޑom@N�l�hGrZ��������"w!Yv���ϠL^a�܇�$��o=bj�&0�6��0�m�����)�P�aV�3`2�Ɯmm�V
{���Wd��UګH��U�6owJ��n�����ĘJ�i���l($)B�y�hU\)S�4J���u��TR����b���	N��n�U̻�&��Z򩈉̼"#��j�{j��h-!�XĉV��Eš���M+ܱ�cSx�ɨ��Cm�cQ�Ո
U�fͽ�ȴ��VX���nl;/#n���Y.���km�w�'1]c�ٕŜ��e��*aNA�Q�&j�8�L�&���̫����R"��dcv��涁��^�W��鱍������E�*_�$�b�sm��6�N`��3�eݻv�mJqe ڛa�o`��f�r���1���(�7�n��\��+,ָ3Jx�R�{����V�-��aJ���ͦ��ãcR^�.]�xthKe'�� �ܸ��X]�7�Z��$*��6��Ɲ8�Ku�7��k��1�a�pA�I�����R���檠��Y�yi�kSC\E�Qq�m�=��
�fյ�IMn��74��[B���3�����C-��7��U'��f6NZO�՘�n���RQ�uj�P�,��ㆱ؝a���$3匦��6-:3�M�� �fܢ�ͽ��;�a���8�z ����7�`��T��oZ���tXӵZqe�JV\��P�4i��m���2���d�1j�`���#0�!�a�[CaZf^�2���Z��T6��CT���[8j��m�Җ#U���>�r�)��^�&��e0@8GF��n��Q�R)�N��y�c`�e��Z�i:�j�7�S3�R�iͧn��o�z�\:	�V�41Q6�R���F�� ���Z�eK��bRjf�䮯	�����	*Ʉ��K=F��Mc��wqۈ2���-�6�� ���ϰ��`�Ș��L�i�s>����Y����KM�#F�촴���/cx��Z�Avm�:b�u���&^Zc"X��f��v�U�kɢ*䐋�Ǝ�-ڷt�k%��E1Ln�́!�b%�L�a/\��D�laǇP[��4N��ݶ2(ʬ�B�'֚�E��N�3>�!,,{��k��SA���S��BqD��d�)��aL�5�֝b��\�!Cb����
�J����90��V��٩�*\�6��w&��kv�e���ԅ^��:1�Ұ[���
������<bC��1Mȋ�`[� �.���&����w327&R�n �mD/4Yf�#AD���͂`b8��d�]��!
��LV$��be:̑+�r�҈9-�FRC �I!��:ri�kzP0j�ks��Ԇ�-h/N�s7L���'*���Z�����1ͳ.FM��L���2�$l�2�j��O�Ȃ
\C��Q�F��6�� �ϛ�a�Ħ���ں�����Cm�t�m]�?,ȹV����J�d7-�5�6g����"�Yqe�x��VU�Ŗ}FK�*��;�FR��������	c�5b� ��
���� �l`�^�u2� F]�.�[��D /o$�L$�ԣ���D�O.�0��md�W%�3�nfl�n�42���tm��i�Ie�S&c�6	�	 �Z9��/ww���:��ʡ+&�P�wE�'Z��Y��![/�3k2һw[���ܹ2Ѩ2�0��k5Y5{���9oJ���'eN8�*55Ӷ6�j�3iPw�,k&b�fQ�N*P�ǧkf\�Gom�"�c�2a��)�6)���2L�q�Ö��
n7*;��m'�f]�k�M�ӓ���j�H4]�`��o�#|w�欜�na|��Ȧ--�,IB�Mڬ�b��K���U�Ϧ��x�4bh0j�2C���z�AV�\0\ܻ�cd׻b�V���X	��4���"^��9�B�Ď�̄�m��\7��fMoX◄���7-�Z8�6����nnM����f�n�Z@0D-^Z� ���G*���H��9Uh7t%��in�	�1� c��n�6��u��ۅ�$�rdR�.�	ؚ9�͈�����i�șP�F,�6ۘRDT��!V�2��H�-Zr�9�1��7Vf2ZD�ӵ�tÕ�˄�PaJU#�AK�r���I;�[k>w����GYe:�Ǘ( ���20E� �ÃA�!��E��˼��˧%��6ӓ��wSFIhE�t��-�)�zl�q��wpF7�>�Lx�<�݉����J�On]^i%��K1�k�{nl��� �}�2�Na�-EQ��i�]����wYW�襡n+O2m�0Y,�{�A<{���!7.6~�ϙs]����[k��.�f%l���B՚�����;�m��&��6�-a�i�JYʥ2����m}�h=;b2vD�$5t.��hQnD�BE��Ê��V�ļ��eaݒ(���Lxr��0ݎ�]on���HG���~�IF 6	!����γ��������쮻�:��ꬮ����+��������;���곻���������+�;��⮊����ή��;��������ꢮ닺���*������9	!��$�HBm	(�@�J>�����.�����넣$�	��ĒQ�H����ꨮ븮첮����ˢ�����;��ꎺ������;�:�+�����;���;�������I�"0HBm ��$�]]wW�EGwY�U]�UY�uE�U�Q�����tb� �@H@$$~hB�����{�	�\�~)�j�~���Sy��佭O�j67p� �d=�9�y>��`V-�sx�I�[;j����P`����ηnr��Z����-�=�hS4���l�r�+��I��͕�a4�b�!u�C0B��v!�Qi���=.�_�!�+CJ�Ǫnŷ�&�w��WBA��Y&�${^���G�(U�ؓ��{�pIF"�e��@X��G�gY��7`n�w'6�E���F'w���-ˠ3��58?�G��^��+UI2�+�P͹�{[&��Kp���ͨK 7��>��bІ�gE���~X$0d��+*�-��y)�{�n��;gr�2�&I5��npF�	j+�@��K��%$7S̥R�Z���:ّ�B��w2����o3]u>�B
}�+J�t�Q���ص:�)O��S���jw%!�g�����w�J��o]���MW�֫f��[ە��y��GQP��/M��I��X�s�9Y7o1g_N�2����g]`c��d�y����1�0��k��n@.�����]ڂ�c-X8�s2s[���,�kC�5Ј����j�K���4���.�CR�~ʛ{���+���RzjďN��n	]ÎI|�ПK���IK�҉}�k�X��ȼx�z�=��@�C���9�X�T޽X,�˼O�-А=��7-V?��aEH,���W�K���٧h0���X�ʢ���Oɼ�tt-����m2�N+рP�}m�d��U╹�m��[�Zr��p��W�b��;��_j�Nq�r����ذ�
�6�ʫ?v�B�'���wDwp+��d౏4�J�n��x�E_h�R"AY�} ׫�s%�8��WIQ�T���b����jm�8�HC0��,紳5|UNU|�9��5����{���X���Q�������>�ָ��JQ�v��v�qg��P�V+M^��x��ܚ���;�)�fv%:`�{/�)��3A�����*�^��ڀS����c��\�֕kI�-xN��ٗO���{c�jC{m8�P_B��)m�iۼX�\��07S06��hRb؉Cv�l��0���Z��ܦ�Z�"f��X�n���ә�9��*��:owL��\���m�:���ݽE���x��V!��ּOԔ��vhU�uЫ9 -о�zm��yPɰp�{qw+�/�O��p�����VM��	S�o�o7��D;gs\�.�✀��g^��I�[Q��r��E��ۄ�nM�O��[��H �ۀ���{{�����u8v���A�q�����%�a�хP����hf��Qʽ�������{��^�m­��f�FWGN�[S
�"2�]�c��oI�7�^�b��X��p��UL��B�3���eu!���7�QK�}k�磌�(�ʮ:�6�E���[��ݐ���ZV��)w�W ��B^�y�s����˕��Wn$*+_1C�fs�#�� �F'q&�z���d8~�I���Z�z��u>�@N�+��t�Jm�Z6��UVkiKK`�p�,�$���,�m�-��+p�ngN�0�B�u�L�x��=��[չК����#�Y
�"��u�@&h���:������M�T�
C�u��m�,�m\6����Tn�XT"{�vq�B�����ƫA�W����ת��5��������0�:���=��]�.�o=Z�Z�]{`R/p�]8Cw}������A&m�C�P�Y�r�������ʘ�X��^Xb�Z��E�7�e�+P�5�=��(t��v_T6�tPŗݚ�䡲���V�1Ci��E�¹�`w]�*#:�����Xw�_�8�ުKx�#g�}g�jI(3yt3Ma�����J��;���t�t��J_)�� 2i�[��{���=[�(��[�ؕ��)mb]eg:��h�hrrb"�]Vm��F�ju��+bW���t�
��K,�Lu�#w&G�O�2v� ������G�B�Y�bp�'j$�p9�Z��nލ�յ��)��P�C�f���Hw�`zv�$�J���r�3˅����5�2�(zZ�)鷉(�x�k9�go{���u�e���qu�A#e����1�ΑF�:e)��8������ǅ�=����"�h�b�v��"i�7M�.3Y[�U��b�B�6m��d6��&t�Y���/H��#7Gf�ӫ����X��p��8��i*�����[�Zs	�f��Q-�W�8�ݖth0������]�tkm^]��.V�e��1ă�����XJ����tV�;�'Q�3�Bs�V��CS"�j��d���=�5�o.��iؼM�j�&���g)d���7���tj�0�V��S��Nໝ0�\���c���4���Z���>t�M��4�	��E���4�g8w�2���7��R	G��M���յs�
����t�n��}�le�uk��Y�lQ;Ԗջ�]w;�w;���S8[׻5�X�1��buB����f�;�n:�N|d��;��v�������yќ��ݱ|1X�{,�f�j5�����bh�cZU�;A��hd8jNd�ŻB���l0�pm*�C3�Ikt�[����M�YK��)
����j��Z�ݣ��]��u��ßgk]N�tj#f�"F��z�-!i�vh&�&���r��WY5r]v��[�3ط��ƄZJ�`.�Zp
KU�%Ys��'���2�:�R؋Uq��]���v�q}��wr<��nb#Qr<��DQ�S����M���L�,˽g]	�x��ɻ�r�W8���e�V�o.<�i4v�=!{��^Ik�il��턦obثS�v�M�o{t�Y�Z^ޮד2r�
�@��n'�6�V8Ήel:2�;��B2�K0^�y:�bU���[���G��r��'�JIB=��f�4#Ww��Q��.Cw`�VT6��C"%&��cnk/]��8�:�����Y���{{%03ٲ
��2��zNr��b�:gg���dl\��gm��γ� �9���'f-��g%�X+r3%XCO��Af��NG;I|�ʳu�j���M�Lu�C
>�����F�.�#j���["%�j��NCL�J�۝��(ix�d�,͵�����UfɄW�Hw��m(��}�]{�T��kMt��J�V]��X�GW�Oz�Y�"��>�X�彵*r�t��wf����k����뇖�"�T�;��&�#��%:������/w�Z|Y��Δ��h5;z�xi@�H�E��+|u3˙�γ7:�S��4�#VZ�������H�lpm!X�����#���'��q[r��F`�.���
f��K��*q8����mb
�ݚƷ׶k�T�-��T��mmr���W�L�Ŏ]o(�+�5+�{J��Q��}�SVan��s��˷A�|�wk8ͼDj}7����f�ֆ�D*��z���a��j�^�*��kw5e���Z"���,�iq��{�0,S-]d��P��hY��5kL���+��S֓�mS��y=�{kc�d�����$dv����'�3tM�7�H�rG)SM^�."[����L�7�[���iVX�Ȧd\�w���P�w����V���9����GX�tԎMm�_c�k���ں�{�=������Yô��1��!�X# �o���JQ��[��U���j�.s1ef�`��w�3�x�[P������m�m����t����vX�bB�i��������/� ��vei�jM��]D�+wt�}Jԯ{�f���٥S��BP�x5VvQ��cS(�Hq��G^w��;zEw�p��=d�=�}׍v>1�)]�w(/uh/"|*��	��VL�vF��̌9%.3Q�un�ׂ�.t;3��\���Ν�2�6�V���go��(�Z�cy)��{kBZ�"�����S�GR���IE����-��[z*�i��.<�s�5i�.��
U�2m��3���鏁�\fnO���b�}���C�a6H��PІ@��V��Wf�B�d�9n2�ݛ�1f��31�Q����o0�I�0|r���9Ps�d�,)Ӎ_>��ˮ뱸��e��AfۓQ9�.l�ll��<O.]|�m|c����Ǚ���b]�Q�t`��[�c�z䪲���X�ID��$y�([��,,}r�e����u���|rί��c� ��y�M�Vi�ˢ��{���N����Ŵ F��bP+�`��D��U^Q�Z�����\���n@�R��,�)q��5 �r��U�_gJU0f�9�����u8��&��ty�+I��Z
x�ü���Vs�C��:�&S�IZ�u��� ��9�S��Y��ޡ�N����܃WW+.q��S����ju]�9K.&9L�Z��e�{6�K����"v�^��n]�{ؒ�[}0���1O�>�k��!=�z���c��f�1�F�nAˁT�Ww)]�L�V~N:�ޜۛrޛ���`aʻhkK�u���nz��-I���YqEF����y�tv���NA���"�г��������e��M�4�yF�L7x����N�o$���h^�,��r��Q�i7�n]Kß)f�o�D��nd���p1���uۣ�%�sr԰�rfL<����n]U�9�fg�0�4���N.f)��"�H���
�U�V�_�K��1r�\x&�G��U�u�I뉔w�9Kq���o0U��Ĳz���weseZv���:+�BC�Ta�[S9XۥY�UN˗u�PQ7�`Z4b�.�*ڙ^�*1�#���M��`ݺ�qR����M��a�S�f��7���f��wq��B9j�ӕ-y��Tx]ϭ���Q��1r����;-Vh�Eؔ0:)�y�ҮRu���P=��{�q�M����[O_S5���P�*�V��*L�vG9I,�O=�̦&e)���J5���,�)h<I#r<;�vz��r�NP�&�lҚaYn��3����Ƶf)y��(q�f�z�p����Wrt۽|6�ͻ������^�6�Ȓ�K5|�=�л���;:T�^F(wr�PQ"[�CNn�uYC	+nb3L�E6�ДT!�B�a�۔n���<�6��ab.nm=�E,�¡7�mꆑ\ɜ:�a�Q8����{E���&�}\��[]�x��V�ӭghNj��G	�q2�c.�(32��2oj0�pq�C{3����Ls���!����q�W#-�V$ejQ�ރ~EhT�(t�H�rvo �	��qDV-�|sYwjc�WnF]8�0#W�nu�`��޽SXĺ��a�NCru]yܜ�Ͱ6s�*!��Ǧ��R�]Ҫl�9�hd��Ֆ�Ն�T5EB4pϜ�
��-(0�S��P��6ċSZ�����Cr���
ͥ5-�9���������^B�a��#���8�Z*��CX�-�Kwr��㹩`&wh(7I%�0>�����v�J���tW՝b��[N�*@�^k�i�w�����;�*|WoIjevm8f-����Hɜ��[��C-9�}�If��s;+F̱��Nu��i�%�2�`P662��nR:j���3U�f�õ�,��v��R����XZ�YA[���D�p����%S�!�`{��L�W�T1�2��o�Ҝ��yt�2�*1+�K��2]�k�����K�#3^A�'H���]�S�" ��}z�F�e$8S
��c�VCX-��ͱI��+������8���3�y����w1����L�9wCD�^�e	���)��^���Ȳ2lJ�)T��P�r)��eΫ�PV�, u���K�/,n�nfp��x�(GE=�х{���4c�靵w]R��m���wl!�:��ꊪʾx�\4^�:V����7V�A���h%�e@yc��X��ii7@��,� �z|�f�6��P��{+�ś���=z�qw6\1�:��F��|��Ϋ�tU� լ5�\*�_'L�L������z��h�޷��u�$ՋU��8a�]�*�T+�qhv����EN��VnG�,$}�4��Q��#�ǒ���>��L�/5I-��؊˿^�s8��'4��L\�VԡS"����s�v�{1�I��z/���F��V/gG+l"���3�ۗ�Hkk��i�k
S=��|��k��F��TQ����+�'-��n�_M�A���V�c�B�������P�0�3�U��m�^��z�)����z,��G<��L�_[�'b+��j��켠&�ը��B�[c�E���-nBfSF�j�i:��ڝ�T�
�GE)�%���ξ��Aj��[���=�|���Wt����[[�u�Qun�Jڶ���s�8���"V��˲��6�N� ql�)�	]�����0��l��%��v��^�/�\�x������	+���Q���׏��ʅ��M#d8藝��\i��`m��n�;l��鸊.�Q�Bֲ%c��ڤmX���G|��k�n^�<�-�X�r�� w ɲºm�s�mROf6��K!�E�[p��5��V�$LX�fw٥��I7 ���1b�+."���>�#յ���M<��o��K���fp� 5*:�}U��=9�k]Lx�,�؍іl��]��m!���b�0Ǖ\��u1�����J���jҸ+wr�e]yo�q�Xn8�Q`�f��Co��ئk;S���sԔvs*�T��ǹt�V�֝2�R�����Ԝ�d@���V�"���V������/7���f�����dX����Y�_e������J���Z�9cͺ�lݱPL�yx)e%�R�� G��S *+��ⷪvo/-��i}���J�
ٸ��3c6�j��(�D��,�r��1�=������W��V�Y.e�5Fvll§�V�Bb��̺͜¯�i�2�e�1d����K�+Gs�k�����v�����P$�	/��[Կ��2rݸ�*긆Km��Z��o;Q�(�/(��j�zez�7Q&�9�wg��Q;�4c�\���9��#�v��ϱ�-���5�L�,�Pm�i7'=q����B�JK�$4�rs�{h�7`{47Ocm�1݁�Vغ� ynN�z�8��gz�h]sk��j��u��v�,wI��6}���ѝ��<	<R:��=g=u��ٱ6��/fw�[��hf��o2�-���:T��cFȎi�k:^_fz-]:N��r�� Nδ9Q���GH�ns�Ş�e"ڷs7�[׷-�;x�[y���|��IO=Z{����1�w��5�I���(�v��_uuX�Gm,��D�nZ@�q��d�w��sv�k��e8&zI�Q<s�n�/I�f2���)��k�K6��N���EGa�=�d��y����y8����|=��Chm�R��q�.�ܙv�l� Ss;��g�ȝ��\�����y6���/5�uӰa8x�a�Fw5��@ݍ�\rPtI��h�=�kHF�Ŭ�\�Vsu��^�a���)c�l/Y՝燮�n��l�Aϖ�=������h�.=.�gn�'\vn�5�N\{a۴��Y������lo`����[nL,x�7#���lZ���h,��D::����z뎚^ɬ�c�ldI�Rٸ���7u]=a1[L�4���=@.�s��	�x8#��e[(ۀ�p3��{�hۍ��f�7��7��.�F��U����: �V���.'(����\f����.*�N۲ت�����C�s������E n�x����/]ϯ k��`�ݛۤ#u҅�N���E�;{��۝y74c�bm��Z���fӮ��tbNG�D1��z�zn�OU�%����$D�nu�v�m�J�ouN[�v-Dmq�b�m��1�7��/6J��2�V��J9��U��sɞ�gMk,�\u���;uJ�g�����:*VQ�-`��tNT��C��9�>�/���oc���F)��J�R>��;�GT�s�GSm���j��m��c�lc��Ѳ�آB��\�٦��՝e�:�����-�����7����ޘwDԲ��nu穹�Dܜ<'v�>m�b8�[���n�d�Iqֻ)�W�7m���y���.��'r�\�nݬ�x��C[j^;h&�t�$Gf�t�L �㈥ �������WG9�m�'g��D�f�X�稴[�|��.�\��su�7\L��i�ͣ�r`m�Ҕ����훗�s�\]��v��^��l�gv�ش�'���t\a�U�Z#ݢQ�
��x�]lA�ݹj�^tz5��s!QU���u�荴��F�����s>[���8�:�.�zN�s�ş"�olk��I���8u��*��+:����v{�;p.�7��p�7d��FY�^�p�Ω,:^�n�i�㣦�mV..����7e<sçh��yN�Ί�<���kx�\�������=�M��YK���f�Z�8�� 5�\{J@�׍���q��ۀA�p^�ƒ�6�\���;{$v"@�&�g�u�tX	orlkv��v�1ɵ�^�9�[�&g[p�z�z�Zg��g'6�g˸w���nݮ)y�Mh�bs�G��j{d�b�j�v�q�=Y�� ���]�����3��=��2�N�ml�����n��\S�nu$��̻���:�u�<�V�˯7O:}�Ļp��ҽO:-K��N�z�rv�q��'���u�n�6��q;������k����`�<��[��j�o��q�]E
YS�N����ƶ���hv���rx����Z�b��OoƋ�L���z�6�^H�'���]���`��PR�[��6���j��]z��g �.X��7]�W� E�,��clb;��ŋ�K�����x��c<����ng�=L��us5v���n�.}BK���:��v� �����%j�8����jd�W>��"�M7�[L�Ocn����Q躠�e.3�6��;s�y絵�q�z�X�t���v�lAm3��m�g��S�v����n^"�*���\/NX���v��M�FS�����팫�n���;�����NݮV屼Z���b���}`B|g	���������k^*��0�sF��ӗ�ܜ7n��s�p����ct{b��TY��Y������V��=#/5�<�Hld7�4$v��*g��s��cHZ:���˻m��ٞ-�G'H�g�r�A�'OfK�;X�`��v�Y0޺;�lv�u�P������pZ6��W$m-ۏ6�z�9�f7�Rk��z����l��[����t�k�ۉ�b�hw�Ce%@�"[���m�k����۞�ފ���v�<`7쬀�u����s>"����YW��b*�꺀3�b�8�]8Q���Xɘ�[Q�l:3�����+�А^�K���6;vݱ��D�Q�z<&�yƮ�vֵs��v1��5۳\�	Z����ۧ����u�w��r���2�/]�Gc�������};��[�w:h���ݡ�z�C��� �=�ً=�EW[��L���]tx}n����m�'.$�C �9��.M�6�mL���l�W���1̾ݻn�#U���!��˙���R��y�<��ٽ���](�dN\��n�G�i�r�Z�:�Q��{v�2C֍v�w;s���te�Xm�^�<�\���o*�͎�Gpr%�Z�q�.�O���<o�]�.w��d���5���tdՏ)1w��W'*]�\�]�a�L0u��txݷ�	K���&�F�U�n����e�#E��;��pd��m��G��l��oC��=t���v�9�-]t�np�u���3v۰ls�Ij�ؼ>���Ѹ�q��0�[<<v�̏@y�z��<pn����s�\P�;v_ixv0�0pnx����CL;�mm����������(�F���r�8��m��YOd�7���63���+m4(8Z;���;��{#�z�s۟&c��M��Og��ΩGE���S��m6h��m̛[�-�C����lk��-p�%�y�woP�عw	�;�G�P��ύ��j^;k������y��-n-\��M�v3�Y��%�m��>^q�'v�<����N.�b�Ý��g�pt�4��V;s�U�Z���M��^��<nw;b��]6=�=�lȎ�"u�s�[�ݞ8�0Y��y�hBn�yѪ��wkE�v^�.m���mU�4\�xlz�;TK�y͸����z�'n.7F�ܴ��N�.�+��#Grk�NL8���R��ۛ�pN{g
��s/iK�l5�c͓�ۭ�;1�q�$�x�ö�޴4�=z��%�hhCrƎal����Ol�܉��8듷�u���ݙq���QY���N���.���#�r����谁ü���ϵ���ē����ʹ6���C�.�=�Z�n�l�u�݉3�\�y�r�WcI�]t���ȗ [X�X����m��.���Of8���g��ǆ���s�Ƿ�]�9���x��ݳ���xk:.�X�5>�Z�I�w<��)o)�s���%ђՆ��̳T�`��]s��w(��ӎ3�{�����s�O"9}sΌ���{Z���nӮ���_gs㳋=Cv���g��V�u��uu=��]��I������z��Nh��Nn6f݀��Qi���u!r��s���݌���q�����6��#����:�Cn�u��s��lэ�-�u�ym���ع�����}�����s>2u���o8�n������b����v��	�d�#��qѣ�LvL�=�������m�r�Òr���<z.�4��xݸ6�}��z7,pkk�m���)���x���>��@%:��c�v�-�v��[�89]�c��uٞv��l��h�7�sŚ���U����ln6<{JyQ��'`5����k�F��7��4v:(�<�\�0��'94]�zT7N'sD��r�λz�dy���� iOu=���ÎܹK6���;�g\��\�vfܖ�r�ٞ0c�in^�m>'��zrmxE"r�ܻ�6�vF��U.�D��u�F{��m�P��fyg����퓷ˑ�oE�Rv�;ro<��8ޏ!�/v��V;[=��z��^��|Qӄjݔp�k6�q�#��Gm\����Prn��Яi]�c��(>Pyv#����#���!�F��8����a�m��g��1�^0��ɱ�ms���n���X;vGF�i-�]\z7��ۛ�kW�ђ3��[�v����=E7]� l,�0c��1�����c�b�ln�)�#�:�c�v� +���:ݗ�aKpJ�:�j�n� �u�S�r7t�z��h�n��X��Ց���z����=bFvp'Nmv=u�ڻ��[���fAS��	������Gm�����v6J�v�lu���<�۝�ǻ/h��S�_k=�x]��[	j�6�uժ�����z����<�ۗ�kCq��q�]�˓ae9	�{`�nM�E�� M��N7Zi󼚼��N��H��(��+��{�u���ėm��.�h���q�vm۵���re%8�<m���v�t�nl�szH����bz˛o�`�8z�G�mu�<eKt���������n.շ��+s�-�mcۀ�&�t�`�i6��7H���Z��v0���ܧ=�j��:��@l�5��<�m�R�c���=頹����J�6pDa�Q*�[kɍ�K:�o]U���1ݩ�9�2tj��L���ƹ0�[�5n�jx���Hk^CM�����p�6�Lۮt�jn\yxoO�QGny���wn���t��Ck���xoJݸ�'��)a�E,�z�E�b���:�5��l���3��ߝ�7px�e�����9�p^�g�m�C�m��y�͆�Y�6�:2�l�h�H�v��,Յh�NV�d�t�l�r,�����y�ٶ�;%�ZND���/3f��[X([nƒ�6݈�i���E���m;�6]��$��������p���$C6������Nq�������=�2N2��8�۷i��t�pq����R��8�$����(8���v�`v��kCl֭�+	�u��gv��m���M�A���h�+n�[��r�k:GC���H�ݯ;^�v��!(�r��8[U�D�f��,�9;���GE)@dՀ�3�i$�m֓kmm��M���XrD��;j��"�I'	�I,�!�e�qm�N�6�6�$I@,�[u�Nt�[[L@EGI��՝8MY9f�����9ծ[[�Vi�hj˻���>�/|��f�t��;��9M�s�O]ld;t�{i㥏;vm�ݴ�wF��+`�ό�a7��n�F8�W�� ��Jø(��n�<�x63��w+�ƻ�Uە7]�ґ�W\v�1����;�pE֝+]����l]OW���T�g$kcmpN�j��^m,.�On"D`�k�������w�|�����o[fvӺwr�;����g ����/c�\b�c�Ϯv���vƷd�G�K�{^�]�\,Y�q�^<�8�m��lE���'F��D9�닪H|�ͣM�`�Ż.�X��;�88{nC�.���!�;;t��3lknI#N�����'�ewf7au������!�]a^
Ƚx}Qیqd.��۫�W_7ϔnƝmq�U�.�����.R�͈��b{7�צ8t�X7/ɺ�7�㣳���/
�6^L��hc��]6����%�
�<H�]a�N�b�^��Pk���`ݭ�]v�ʩ��λg��X�Rn�u�>�z6��9����-��T��(	��ks���jGe1ǈJ���z�ۓd7>E�c���b�<�2��k�|;O	h���d1p�A�wEk���y�캶�q�8]=/��؎��S�^3���i��ѓ�瓞�	���񍳻t%��mX<��u<�\�N1Oo\�v:�^��c/;98Nv���8N�Ca���[h�Ά6��C<�=���;��Z���w�������ܝOi��8�1x��M��^[��`Xӷ]su�u��c�m�]�bq9�Skq�z��O\u�kMVí��n��4�(��x��F���g��n!��3�����]���������lR v�>���@���@v����8�ix9�魟]ucq�lv`��ѵ���:6��u�ۍH��x��q�4u���ڎ�vT6���n�w<v�l��:7:KnP�<<�S�{E�g����S�7www��|��2�p���x�����;�|rrq�*�ϲ�=�m{׭���3��זW��������g�qˇ;���n}�Do{����/=�^z�g�y{Lm=�yyo=mދY�zǼ����9�筷�Ǵ��L��hs{۱������k�a1��!�'a�Ȏa=�	�w���6�_۝�*n�q���7//d;���c��G@=�����G*��G�s[��� G5UZ$�a�Q3���&2�	��mlb ��?L����en�������H�ݺ��b�H���$��oZ��`8]��""i�yʕk��$$�{�a�7�+�"V�3Xg�5�� ě�m����|��G(�TH���i�������I����-E3��w"k��^�!<q7�2HJ���&�4}�ޝ�x@�$ї�փ���8KE	�W0���1hm�{��mlʩn�p�W{����X�4I����fG9HC�=��)�3�Q"%x������ɨ�;�y-�6������KX���]���'�U�E/|����W=wz�>����BzyM����O����̂I�tx��;9�T;/̏�9��`�z�{=	]���.:Q�KE�A�ztm�3��o)���st�� ��M�Ϭ���\k���wfÒ&h����E�VE�Z]g�6�^�\����9�o{ON�n�'��ٿM?wQ��[�"�D�<G��@�A�s��� H3��{��:�$�~ti�&�?����X
m�H(�b��E����luK�ĝ�.]f���A�s��� I�r]���5�#���� �u�\E>S3��BRF�#3���� ��&���w7߀��{٬ώ�������'=ɘ1����|��5S�H����41�e�v;bx�-^Z{m��b{P�.ux��瞺�>����yϪ��,�y�� A�s�ͭ��$�N{m������-�F��}(y���?{{���j{�d}v�K��g�ɬzqg�f�K9)L�$�I��zID�O���q�	2
K};u���j�Iܾ��b�(v֙7�o{�l�9��@d����-{V=:��;3�n�{9C,�V�IË��Q���	��jW�x�w��Op3/����,7m����k���-&��F��́(�M�2k����Ta ����e����}�{��Ēwy����o���Ě$�5z4�1����u��M>�$&���࿍��0�Q!��I�h��������톶�;D��͒h�M� 1�{y�A�9��7����u�'A��]v+Ul�ݞ5�۝��5~� ��$��
�h^�}�.���KQQ������ ��w���8��/k������} ��t��9ǣ���I>��9�f`�x޷ږ�~Z�I������Iz4��$�D�]|��]��S|��*����Â��D�֘���6@4J띮l�:�s���s�| ^{��� ���:$�ι��^Q�(�,3�I���۞�a�ĒG-��4I$�3�4�$�H��s�Oz���85p��/��	\�FU�k�c���y
� �� �_���?&�V�(:h��&��}�+�x��9�/eq�Il�ʣ���tqm������5��Ta��Lmk��s"@���!g¦׭��� !^[��H��&I�$���tb�[9�\�+@b�]Xg�<�E���)�F7rz�ݸ���j��u��]�g�6quw��|D�[�޼3��o>y�~$�^��I>%�䝏}�ʀ�D=�z�;��5�w�H�ڪ��R��Qo�����c֑F�X��  ��i8��D��0d������涧s�%�y��@v�$���B���ŀ��w��I h���r�M�@?�F�$��w��<F{��7i\��}��{Ğ���h���t��$��{���DE>k]�L[+�z����.���T;Uax{پol A���\��t����W�!5}蓢Oď{��T �&����f�/��7�b/M���b�Ÿu*щ�k�I9O�<��Pf�־ۀ����ݠ��Qj�	���U��U��6�7�9N"��+~�9��6n�oX ��V�G�h1�ݗu��C���槓i��y��m��{nYyv.7��TF�����S{o��9��ۺ�{t�u�đ�n<�vc�];�����8�q�E����Wru��v�v���h=k�U��*'��<��t����� X%�.Gln�6uy$vX,l�[�y����ql	��!H������b���zIݻk��x��̺Ki3�v����M=[nq�h䤔�����0���&��,����'�f��ʄIW��`neͫ�i��a<����ݹgB��"�/ �ZtK/��Z�أ�7��7;�>� ����� g=ɋ��o��oW�� 3�ԑm�U*�ʌ�3���=�e�� .;; ����� �=��kc�=ɘ�惑��o�w�V6kg���B����O�lr	&�{ɘ��w���{^�N����+�[����{[�7΄ qҺ�w1|O=��+;�l�2�{���� ה$����J��L�D�OD��ׯ36�[Nnl��n�$�*�(FܟY�ۮ[H��;v�u�oc�gqv��{~�?>�gy��&���l�%�<`pOE�<Tg�����KЯ�'=*_l���(�*�;$�����>Z��^��9%����@�����o��,�p�}ux��}(��~��,��X�uy�/wveR�";����;�L���ٖ���5�h�!sy�=D����2M~�=` u�-��}7�s`�[˕�8�����z5���A_=�f� �
���z�ki����� z=����*o�ˈ|�fF�Q(�"�*��%��©ey�����\ �N�yq�߻��]�}�{��ǀ�!�d�iP�Ș	yL�d;�. D�����U�o.D��o�m�I#7�O�I&��{��٭�������ⴰ�F!V��n��UA��ێ���2(N��%��J�S"�B�!���ă(W]�����ɦ�S��q`/�@.������lU��foz�G'��`����X�)���T;Uao�N=�
ҕ�f���d�D�^�:$�$���$ �S�e���V����n��q;$ǟ��3�@��{7��$���{K�vGu�E+��e��)�)��w}gm!�`�Fez/N�}�'X�̇��u���2���h�h̴��\����t��i�r�؈ا��π;�����4櫨q'+u��>A�{P��=����M*��L�`�>����H�����=io����I�5�$��I6�UB��Q���{{[ h�y�Wbd7\����2.m��}�y�[��rb��{]���ɮ:5��:凣;ss��۲�Hm��,]U:6yŋR���o}~ ����W^1��� =�����I$��}��<�xz����'	���{.| 9�{x��M�ă-�Q�1���펱��[z���VB>\�$_N�zID����%f��uM]����>�^��j���<��l�T  ��2I+��Wd|<��W�I����ilm���`}���~���ݰ�<$�~�ޥ˅����TH
y�*Ě�~�[tH�y~u���G�4��H�3�e1�qjU��G�k	`*�t�ڼ����NL�����nˇ1���e���أ�=���q�p����B}��x2���x���^�g�O���D�E�����Bs�mP	]������j{���m�e���^�ѵcM^et��;X4��PFI �^m�v�{n�I��m[u��d�jTE��X(�B��7�I:�UK	\��#Y��x��q+�$�P��K�=�ˮ�Ϊ;�t`BISٳb�1�E���	yL�f�vR."��,�j� Y�w9	�OĚW����z<I�/�Ӟʞ�;jR�{����dU��g����� ��z� �T��VY>�s��� 9{:� 8s��@pٮ�~�WXC��;E5x��= D��x�Q$�z<�#��y������9���$�}r;l��W[n��"��ݰ�	5�OĒf��lB����o;޿�~�� ½?�4I=����yevp���f����_�.^퀐\��R���*�zHNQy;H�6�
�X��`y96�����bsL\��X���g�gc
Ӭ���D:�w\	�AM箶��öZzؗ�����.���񞻝v�xU'�Gmٰ�8t>xۧ������{���͊�޽�p%�(�/A���k�]�3�+v�,R��q;��+�`ݷ;ƻ/98�g�gr���rU�lK�N3m)��6�i��5m'\���z.0
����9Ŕ���x���x��ȶ��x�*ț�b�3��[�N˺�Y��U��h����\
;a7�k����P`:�D��α��I:�h�h�����!4ۓۆ߻����@?��,�r��MX쒹Q�5�����~7���9�}W ƻ���#}����`>/C�����\4C�����4�Q�[���l����	=�{̀'���z�V\�;m���TI�������I��g��F&)�zH�9l�җ��mz�ɾ�o�_'�$�N���`(��թ�B�߀T�̹�.5��֍J�c�w�l��$�N�<o��-�^�kw�2MO���� ���Zx7��B��J��@vM�ιC���Wh�%�Vn�ț�B�����UTͮ����n�I1��{�W�Q&���yϡ4I$��ۢ|����wr4�v�d�L����֠���d}yd�-:�Y~��3�=�+��LU�13�l}Y���[R������ m�}ԃ�9Q�kyw�l��?A�/޻>ew�'E�P*j�s"����"4�Y.k�%�DI��z@'Č;�� �����>����2J�+���8n����>���D��u�I'+;��}�[�w\�� �{��IP�Hþ�3+w	h����I*���ۚ8�s��Q���o�}�5���l�I��z<⳼vm3!�@|w��ok`�M�����e���|����I�&�:�]crl�.E�j��:I�$�G/��@2OЮ�WlcΝyv��l���D����AL�Ln��u&�v ϶�y$Ƶ &�̽r�� �g�L����W~�����w{��� �=٬"`^�7`켊�1�w���{�,iz���G��Lx�׽�1hm��y/j�u��lm~$�_w[tI$�
�x�$�i<=���{7��s�X�*�vB�Z�g{� �^ޱh_�7I�C^�P��1���7������۾1|�n�OgRy����끬EJW�Vg`v��n\*����+���ܒ�]�9㕒$ʵ��wD%kfͳ����E�Y�Y��A\�'3]v��,��v��
G.�С�vr�\�����Q��E��m+Z"KC��TB
�.��xáyu�E�׺�)Z��b�f�(�[͡�������$ÈUIX���U7y����oCdBnq�Ӊ��
ջt�����B��J�/��c+V7��0��a;tl&��i��av��s�����5e��~ur�R�,S�ܬ�ϳs{�����<�����Q�F���]�^�^w ��.��}�hKw��EJ�']Ϲ�'l�g%k�q0���4�*�ɓ�7{�\M]�pay����[�]�Nc&�T0�[:����ǕC��_p�7s�Al��;9]8j6�T����2Al�Ю��u��x�%c��ݰ��pj{(E���˄K���}>�c-�k�[O���y%^�`�v�p�'dY-��� }�m�ʴ���u��WeQ((i���"��nЧ�2��"]K:�p�c&�Rr��٩���J�9����E��//���^�A�#3kV��h���)�x�5XN��`���N�ۓ-�jN���Iz��u�ҝ�߆7r���Z�˔�M���8�s2��J�Hd��Z�LG�,�Y8��wX4@94F�V�%�Ue����[�jf_S��B�\�ɵ�o\4��_'�)05���FJ����im�7ٍ � �C�Ƈ��B�';���G(�Ims`��֜I[Z�8�fb�,*ά�[n$����Ƒ��k-2+E�ۣ�&d�e�q;k$Y���Z'8E%�r��n�nr\��F���n���m�;��gf�c����lS�E�i�Pڬ+kf��Vi(����q���\H$'Kn�P��	9��m�kt��6ܶ�mn�ڱ8�E]�Qͬ�tp���ֆh%���9�)¶����l�S��i�'*Y����GQBDr\�		 t��fNmp�6�P(�m�%9��2j����
��6�N�N�6�GK�C��9#�"K4A
"R�v����4�5�[n�K�6��I�[u�6�eI;kN�HK4�����9�@"�{���=���`��i�,!YQ��5���:����n~ !��|�>k��` �����@�Y�>��z@#s^ɋ�����+Se�W�;�pLz#w��=����ڵk��<��D�$���i�h���z1�QW��O�t=�_�/��D�uWTq���V��*4q;�>Ÿ�lz�J*[)�±WJ����y� �W]/|����� ����b�@ ��zHN�L�g�_�Ͻ3���@ �-�2O�`�3>��f�a���%BI�A]��I�Bs�`O�/F�d��=�zJ��C��؏�/'8;ɼ7m�ߘ/kΩ�}G��Lx��`{��*�$�ei�W��{\�,���sz� lF��{{�^-W��`(�fi��c��wt�`ޫ���M�@I��{�BI$��vO�a�]X�R琇2?^��7������?yIf���Q�!J�3Zu��sԓn`^`#f��G�=g<g5P��s%���m�
f��7�w/Hm�\�GYQ�k=�o{�w4��+��F�B!	&��,Q&���l�I&�n?����m�����t��V���k�]m��û,���M1��׳]Y�����*��Ώո+[E���B���İ;�{ٿ�  ��v� ��s��x;n͎
��kL�D�;��>�ӫ�W[@9l��K��>{9�X$�3�����S��S&�}��`J$����L�$oz]��:���L׵���1����(;,:=�6J��D�$f��&I5D��ݣ�o���lH�{�o{b	�v����4��q�$�໽�':�����]�%h�ټ�B �݉�I�O�/F��\��|�.�/��"<"����Ḧ́���f�g�u������٘��-��0��l��4M�݈D��N�lz �[�y���(�ikWu��V����u
���:������=&%��˭D�q��T���7
z��Z�޾�\�(��&�ԏA[�5j�v5u�/�C���.��\�˹ɵU�r��w8�ȎgNF�6λ!˷nsHrˎ��d�-�>;n�]���q�CGi�\[�1�[Bu�!��sǭ�����c� Li�K]��ˉy���Z�햃��ǭ�s�e���=]�]\�WW5/lZ�s;�ݱ����ݡ��8�A؍ur��/Z���V�mҾͭ���v�=��Z2������M[�lWf��l\7�t+ʪƹ�B�}�����*5�g}�������$�Bg�N����Ue�~��ilb��mo�G+`��*���)�n�$�m{F��(??srH緱��OĚ=h�����A��Ȼ�g>�b���c��u�� |�7�&I$�gD��&���!�2�K���{i ��/9�`�>{��k O�}c/�X0�e���I����|�����	4H�����O���D�tH����g;<w��)�n �t��F:M��$e�wl3]&�L��M7��	J2��p+�񿨓D����~3����Y%�mV�|O�2L�B��JDA0�n��͎����Vu�e�E�R�BEG􉒕�N��,�ꪸF��#z����� ._oY�� g��I*����X�l���؀tI����`?gm�(���#N��w`��z�<�E���lȶ�D&#K1�z��'�J�ѹZ�g���E���$%���Zg
,����t��ZS���[�i�`3;ԙ$�GfƀtH��yϡ ������X���2��V·~,U]g����� w���{�a��nnj� \�޵� ������J{��ݥ+�}��E{���l�5�����+u��4H��� �	��dq6�eI�I���\D�T�P
N����LDo�7tU�~+�g�$����I$�����h��3_*<�F[�i��Ҡ�D�J>�3iq�k;��эit��an{s�4�f�H�k�bmw=��)�n�I6���3� w����Ě3w���u�n|%r���?$���{�o{.j����,���|����-���_���	`!�"���5D����$�3w���b�7���{3]��m�(���#0���ok`�$�����<]^�����N��^r]q3	TT�Z��EMB�+��m����}��z{�yO�B���E�E��<��Qg�vˏh2�s�FH�I��F{�������q`-��Jr���b��J{Z٪�D�M��}��E��o�MD�F�Zǅ׊���j�����Oү��(��p��g�G{c��'�k��t��1^����I��ޒ~$��v?��~$Й���~�	�jk|�G-�#*����ϩ!�I���x�n���X�2'F�VҪDs���V�����|ut�ĢM�b�D�=�ӦΙ梔T�z0!'�_N�T���]_�E��ݰ�t��d���K1rx&�+��li&�%z{�@4&z4��:)�G��{#�Wf����3af���4�ַ�k ���0���;���3�~�$ ��L�D�=d��L]fX�n�t[�z0K��q]xz�@���g�X$?_o5�Q&����yܗ~���c���Crs��ĀyЫ����]|��6��RujF=�L-r�d��.�2�X�z^�.2t�fU�EKr�)Z��<=6~@|��ϰv�\�Nȋ�b��[�� ~�{͉^����Sit��$�Yݍ�~&��d�I����T�Xn���v�{|Y���X;[c���U�NWBWn�{����[n�E��J�S"�B�!��>vA	��s@��ɒI5��&� �����M\ʘ*y�M��3�q� �'ṱ�I��v*�V�*�<;��7����f��`��|�4I����F�I&{��!��k^*h�{t�u��>z���a����g5ϰ�w����  Zܓ˛]C�+}$Ǥ��"/F������,�sU�JYj3M�kݓg�T\�yN�$
��6I$������4I����^���C�7#��4;����J&���"3�o��6��w��M�d��{���P�w4�4H����B~.��hu;��κ�S�h�#n�v����c7�3�Th������T���$�툩a�]{E϶Df�+]綫!XP�˽GYH<X�<<=t	�!W�L�{j��������oh�q�����Ӡ�iy��pss�q��kr�٨�z�x�Ax�m<�\�����+l�MEҼ�@D��ۛ�AN�� 9�a

�̒v��|d�e��w]n-ڳ�]�5��ݱ���=�R��G<kW"���;j��ZE\���O:����v7��xV�f󱺹��{\��mo%�y+r�c6��Å���XHĎ�Oi�]F2	���\v��Y]�ee�_|��*H��+���i���؃����[ d�3>�����+�$�co~g=�:$���I
�U��� ̱xp��O=u�N�7�w��y�R����o{ ���f,x�^0�8��Ÿf���v���Z��V8XtyzlbQ'�Y�s�h�� M����q���ݎ�$�;��I4I.��h:�~U�n�Bc�u�|�2X���� �y/y�M~$�+�m�I$���V\.�j��X3w�,�JL�A�)L�QY���$�5��!�wg�u�T?���h��W���tI�4ɻ�^��s��>��ʛ��;��	f��di$�#I�Q�3f��h�"�U֛��b�w��u�+c���$fw��=�G=�W -�D���Y����ל�9�M9��XonqɵB9~e*��-s���Q�̥�p�:fE�>��S2b�y��Ҷb�gQwr�T](�j�3%Hiǯ+v앣G�m�ͻ��5`q'Dy��ȕO���b$�������Y}��`���s1�	�?o5�|���/|��^]��ھ�d�3.��d�^�X�s�$�TM%߼ۺ!l3��>$�N_�- �?�d����ʍUhWc����{
�멼��0�{�c4I$�{d�O���zU�#�+�:4ލ<�{�0���⊁��M7^oV�h�L�{�T#����A^h���{m�� ���ӢI'�=�zHsg�w�'|�����% �j�3������F蓴��;�n>����ſ.Ϋ����r�0�����	�{zŀ�����`����QG���;{�hI��O�$��L۬Q[(���Y�{x��vi{����L�Z|�q�~$�~�?�4I�=�zO����o�O��[K;V����_�ܬ&�ߙJ��!k��b�}�{6� ��yy@y��u��k��ҝ"p�^)�e5V��ٽ�����gkgoUj�6ä��/.;���FKq(�����k�5�@%w��W��I���  o��{{[1yOvD&퐮��o��>�	��f� �ڧ̒MQ'����Q$��؁�{*p��V07�Hɿf�y̒����i�����o{
s��r9�Ҩ������{ޒ��4r��hw�z����g�l���`��g8�Mں�BA�i��t���N�mj�QL�ׇ�7U����1`h��{͉�'�N^���^6U-[�������m��@�:���"����%�s(�d���2K��Y ��R��W� �>����H��v:d&*�N{�.�kz�>��6�V�"#׽��'�MQ#=݈Nqn��<�d����$ �{�o�7y��<���N*��E���F�}�&LWYݨB��$���!$������ME�j����I�<{���n�֨�Uf!���R�yV3���4Y��u9.7�1PJا"v+�ud`.H��u�sf�N,��������o�?o�������!7l�u�� ��]&I4Mr�̝������5=��%I$���h�"�h�
|���_q���ii�k(7o�Nѽ���g�j����rnފ�gi�8�dl�����-CV��P�@�n?К�I#7��3D�$ЋѧD����R�M
X$z�=�o` ��n�t���E@��G&<w�f` ��έ��?s�C��s<�  }��π@|��F� 
]���;���;�?ub9n�:�lr�2����`5��O k7�<�wCP��� ��{���$��� {��6�V�"#N���z�%Una4����D�]12M~�4� ��{��v�
��j㤒J��\@�Q�2�Zh�\�^{y�`| w�����7Õ�l��������I#�ѠL���*_x���8��!� ��c��^�w�fi�m���9]{`�F�Y8U�9���!my�aJ��fR0��Y��)q�;]��s��n�)6Y�]� �\��,Z�|:1� s^�s�T��hwK��s��]F[�2}xz��(Z���k���)	E=���d�a@��Scj�5�d`�r��R��U�Y\p^jΣ�����54DI�Y^�F��x�qU��f�LՉm����78+UpT��� ��ea�G(u��]�Ua
P�g�����ǽ�M`�,J�+]F�/n�ɆN��]�t��v��t6���wP�vi�k)��3F�]+Z�Ƌ��4����R��K��RlR �m,�!x����
�:��8ri��cB�Wm�.�;oH:�%~��O���^U�N$^j�B2�m����0	ء�fF�ne,��'�0l&�����P�� �M�$j�CDTu�7_����
��>�*x����)n�ɦb�����y��H�b���̬.�1G�j�s�B�Z;X���.����y�z�#l&�ۇ�#�	��D,���r%�U�&�D+X:57���{�jV�J��&�H�eӺ�ĭn�*&UÆ�`M�Ҧ0�(O���I�dN���f	�0S,5�����$f-8&n�JQ@�s �����n.��.�+�s��J�5*6����WsQ,�9�{��0N�0W�;�KS�Yl��&��<�}� ��VΆ���8��k+5m���BgTw�t�V���=��4 	�O�$�H'Hr,L�:��k(�D�;lvVV�m'Y��2Ҁ̌��m���s���I8�gbQN�;6�N"�)(Yif�������D�7Y�tr���mb�f������93&��	���ܗ%�kb��-���+�I%kZ9,��)�gm�6�Ym��K16�5sl��³-������QM��H�h(��8�.N��9 �kR9[Kf���âm�m������D$��6�(��L-˓�K��v 'GS�a�I(A8�GH;-'Gĥ�ͻ	��(�ٵ�ؓ�;0�q9�FݫlQ��!$��:mA��Ҷ���snnm�#�)i�5�q#�F�`�4��l+t�[k����2�Sr�-�n�}cK&�K'a+����������nN;\�prD�۟A[��q�n���L]�1�B�Յ���h�+��+�\u�v��;NN����v]X���ۙ񎞇\�rɅ�]���u��9��"4�Q��IiF
T�Q�s��g��z�]�Hv�/uB&Q��c�Dny���^�ZzLrScl��r��뵺Ob��{ٝd�6R�����>о/I3��Z2��59�z�\-oG���[8�EJ'���R����.{�W��k��\�c��a��� Q��p�p�:n����B�vs=f�۴Q��4X�I��7u��wM5�ۗ�<q×v���i�X!�e8ʡ�;�,`ū�cQ�ӗn84��\e�qƵ�����:-�^2���*]�[��c�c�<�y�&Q������<"�]�y��6����SaNyy����}��lp��a:Dp�G9��ȡ�>�
�v�6�TP�RD�UZ�����l�p����n�liՔ!v��^.���s�sT���zޮz^��p��YG�'�pt[k'<�B�V��^B��n}�yl!����F���m����F1e�
2��!�nB��[�é��'O�ݟn:ƻv�\�km�`}�C�ݏ]��c/m����nGsVέq�`!��0=�9s�u�[�\&��gl&3t�Y�vM���1��6�md����o!�v�^��狣�(6\�0����^A3�e��Z{d��G��ڸ:�j����z����`f9����s�kY#/	�ǆ%��2�u�v����1�u������r���ɝv:�!ݩ�c�Q��ͮ<fN6�X��ֹG�t\t�<�Z��m�%�-nvgq�67I�	�=���7f`q�]r��y�ظ�s΅��lm��k�h�R��z��8ͻ[�8�x�.��]v����ۣxם���7��^��M\���s�N+%ڵ�qR�Wsh��[4-��)У����ww��t����hzl,��O�\4��h����g+z�;`�r�v�wMnV�q���V�1�9 �=�����{F��(m�<f5C��ү��Ѳn!ԝ��y6�E� ��˪�t2��l�eKUϕƠ{6�y��Gw\p���&^�՜n8��y�%k�V6�;�]���t\��={k.N�\��q������ݱ���sn���ͮG�"v{����B���;���t��cfv��������e�ޯ���t��@�m���� ^Ή��Oӽ�I	��k�<�l	k�x6�/7�g�'���6�v�Ixw��Ģ|�?�RG�՚�i�I4764�$�L���*h��,DtwH��5��]��dttrc�{{�b���{�Bh��|��[�����5{#�I%'=����߽��ka�tY��X���U�tHo}�a�D}���Q4��2h�I�{��(�D��X�d�3u��9�{5� w�L۬Q[(���Y�{r��&���I��ߓ�!�I�,~k H9�w7�� �󞹆�=9�m�k{Z{��,����:�T�@vG^�V�:^���sI˴��/�5TqEU�:zI�B�Zjʮx[��1`$��{�ͭ� ����<6�Pz�,�z�O�Oč�{���4�Ϣ�	P���!Y%�cd�C簮���V�P��UW9.��tl��J���K#�Eu9���\n:�t7#�����&�u�^�ʝw]�u!��z����{�G��}�!SF{��|$����3=Lz!7����"$�����.\�= �iH$$�3l��T&��n��g�@u8�/z)V.����H���I����cd���W����.�f��z��10:�I'zf=�Vs����s��k�NI�=�fqX�7�s���.+��+br�b�00�{.
{��`���7��� ��}��h,�vb��9�o5�.��)�.�e�}DS�r� ��7#T�/[1�$,n���H�$+�D�K���}��b��DDk�����`�
{;�>9�|:���u%;�=F�ޓ�A�M;�����N�8�WUM�����f��|��Z���3kc`Y���� S�*���W����=�cs��	Q�0#}%�$�W��@4L��Zx&����_E�e��s��m��x��v�6�͔WCr�iZ��Q�۾(�36;�u�ؔ�F��OLҜ����s��a$�O���[�mǬ��Hs��H�$�3n+�\W��\� #$c$�H�ti� ����Ṣ�3�x��OP��$���M�{�o 	=�V��¸CD����$�I�sѠO{��}yk���r����W��m�\����Vpn��^�\t����J\������3k�;<�u���ny��j{�t� �w�I�5㘳��(L�v.Q���Ń�sy���
*Z�tX�~�c��rjGm�^��9�+�@?P�ѦI�M{��T �M�ׇ,Rw��y�Ӱ�E+�&��-�9��N���!4I�Q*��9��۶��@'7���w�ͭ������n�XQ��'O�W���� SS��Mh�����'ĒM�~�h>���/�3,�RNm:�X���y�9���9CJ��p�-gW�r�ܭw86q	�M���Qxx���	�﹬@'�����֫H�s5��� a��!Az�t�h��5&H�{�$ �0������6�>_<�3c�vV�:d{\�ƴ�ҥ]���6�E�v�I]�����uJ�WGG&?3��� �}��� >
s=4������.��:$�&���l���������9�wE���\��I*U�`V�v9�r�k����w����3�M��?n�ӹ��&_���
5tr��h����߶ �w� ;;��=��������[��M<K{��s�YT@����O=an�xH	�@�պ�Bh�D�����H�~�։�>0�����fp�gw��a�����M�AUh�'�Zf�?W:&�� ���z%��!��Ě��$���?z��/��M���AA�M��ȼk�8ø�'S^~�r�Z�n��2�D� ����P;�x�ٙ�3;;�{����f#eP�&{���>�����b8�$��S�s��).���n���6�};�]�lc`7G���t�d-ss�3q^�wf�:ፋ9���׎y��2�uN.��У��M��'K�v��m�<� {���XCoi�	D�Ŷ��܏���-��h���Ӝ�W���ws�1q��n�V�mΕ����.t�Sz棎�E��<��0\Nw:�.�u;���i�0�:;n٥�;W=r���n}��/n�æ�3��8��x���1�r�7Z������Z�֫H��O�#��s{[m�g�k��&�_�4ꉹ�NVs���>��E���v�����*]���kl�G��ry��hwR�ߟ}	$�M��0$_�4�$ ��媖���ӛǿ�U�M�h�����ַ�k׳�tɢOĭ��������gĆ��z������6{i�օe��S��;�5��x9�$�H�ى���Q�D�M{��-ݞܴ�����Ik������ʢaj����İ D���r��[�U�JӇh�k�� �Q��$����CNޝ�Ϸ�,��[]\m�F�
f93di���ݮv3$�k]�T�e���zy�q�*�Nx=�bg�I5�Q6OĚ$���zHJ��|����9�c�A�M	�4ɭ�3 �2�Ѻ�G��loļ�7vx�d��;�[�4R8���|���r^g��v�꙼k��M[gn:��wc�4Td�;��4����L�./��,�`bT�ɷ[�x��A�u���ܒG���7�D@�wvY9�s�����㴙��k>�Q�1J�WGG&<��f�{��͈I'~<=<N�����ɏā^�5��w��w����XmZ�RWa��o��{�{=��;����5�`| ��I(�Hzf�;+ޙo�]�	4&{y��rk��օe���3�緵�@I�c=�X��WZ��M�֝I4w��IP�	+zcf���VA�t�����Zܖ��.5��h�R뭲�X[�o�m�(n���v��v?�ʢaj�������M��s��I&�ޘ�|{4z�,,kO*������2�а(�]!&���;�E?�\�5oqm-DI��t��4Hzcd����<lwk*��3�<tI������6Eղ��?l��� -��3�'�X��M������c{�N��ћ�YٚeF����9Cp�-lC^���T��&F�'�7�ih"�c0+u��F�� �w�)��$������ j�[�u��x�C#�������{��V�rOoՐ�w��o`�|k���@�㙼�`�7����"=��g�DJcJ=2�Y�.���� xs��%�������u�zHI$�J����<d�W}�||���/Fr�ȩJ+U�+�f���"2�u��3`�beQX����	���kQDI���5�� �!{��3�&�5�<d��*&���>��$���Tɩ{	ωeQ0�\�/k��X7����ߓɣ��p�k�Ͼ��h��]��D��?P�����D�j�)��������V�m{�|&�
�3>@����
�$����D�'��_sX��=�{� o^��`π~�o5�|��䶷���d]��~�W�;fI��t#��H���3D�$�=�4��I#��s������+�X�w��Q�T�J.*~����Z �+��ۛf���ܸ%�s��]W�m��m!��Of��Y�fogr��W�g��HI�=I*��l܋�k�b����1௷�İ���sj�
��ea$*$�W=��k��N��I����HDv��SV��WX�,�u�n�]a�t{\�ü��*�'�]�_+��v�C�T&�������#����sX��/s�I��^���Bko�OӸ�Y߰`|�� �5��֤l������B}�L޹��5>��۸�h���L�I����HA�����Uuɚ��+nl}'>%�D�f��30���9	$�s�R��O$��8����"��������>q�u���d�OW�H��5��M�TI��{���M{�]X���:��+��mU��r�'���6l�A��~�! ��i�x��ק��X��RlI�I��l	D�%n⻎Zw�.8���+�U�%$6У���#`��9���Ս�n S��5x��ؑw�3{������H��vR�z�"6k49�&Y1hV^G�� Rd\�C-㳷���lv�u]��c!�v�Wk��q��՝�+�ֳ��Y���pn9:���N��`}��LNN�훱�!Nn�%Dm�N�X�F��2n݃�887#u�8��Ѝ���e4�n7\wnԯ�<qu��ҽ�g�y��\���;E��x�,�z=e��D��e��w;]�0s�\>�x�;��a�÷i�@U��kvݳTP��@�`z�V�0��wm�v�I纬��ubR]<��\�痼甿�E$��
w|�� 7�{�BI$��1 =���x�nZ�{� �'�;�щZ��,f3+0�n����y-;Y˦U����\�?�$���{� 	D��D��ܺ3��Nm]��^oנrk���82GX#0�{���6 z�wt�r��!N�����/������b 5����sc�9�-� -�o�^]�Y�����v0,�d�9	$�J�Lo�@4=�5��t�#��8��$�/t��^�i�h�h�d��֘ T�(tELJ��=��I	$�%wLl�TI�{\i�g��r����h��O��=�>Cl�p�7gk
v����ж�tz�,�������sޖ���[�8����Q$����=�4ɨkӍu�ʿr��ӱI%B�I%{�'ʯ��^Qe�*�c�N{�ߦ+��rx�Q̱ӋyS��gc�^�&�Y�_[����^ȭ��������n�*{4�3�{qH[Ѻvkpᕱ������{���$u쿩����7{�����".e��5or!٥%"���Q4]��ߓ4I&��'L�_�=���0��{e%oLl�D��uD����Z�"�f�s۷~�Fn���y���s3��� ���k ��ݞ���e�߸�����9q`vl}9Z-��T�B��ŀ�w��c����xm��o-�߻����f�X ��ܳ�]��E����#3%����=ms���f�'bxqv[9�=��Ǝ :�k����p��-@��>�|��moٽf@ ���nQ3����+�-�Y9�q� �A}yu~������J	I�2l�r�y�	'o5���g��VK��&I4I��q��$�{��I4O���lu���<�}�t?�euRi�w�ŀ���9 oپ�/��<K�ٲK-�ۼ�g�O8ی�w����7�ۄ�L#�=����,:'�t>����J4�q�Ua'{�Φ��2�s�ob��RЦl�f��Д�ܮn"m�j.���O7�X7B��aʰ�6ka=@jѫ��7> ��\�rS���� ���Ā�j��"Y��cmeZl��YɹY�r���������[���^������d����`k6f��|/2�p��d9��-�S�k+��"���*��cB�;��ޜ���EʰU���1TVV�6��jj��W�e�x�����"��� /��KIgQ�/8u@��epW}��Q�m���M<����<.am�h�
wF�[
�I��"CV�o+Ε�̃;`Z�h��E3��kke�Të�)������s<�&�{���qN�}�}o��zo��K��z�����C1�av:�x�ۥ-uX���Hh9	�J�e��}����R�w��v���9#�Ew��8�%�$Tc Kwz��Wv'β>v*�[�ǳ�-�ކ�6�\Rk���姺� �:ӫ�`��&���q<�/+��i���³���7off�A�a��)e*�Ѕ6Ntm�4�@��'f�
�|;U0YZir�Q����^�t�-gy���҅�i�"�k���g=b��^օQ����v�X�wIT\��Fu��ۙ����^ָz�7�/�=�.P}�=Y�)�H<T*�E���v1c�l�#,V�׊u o5ʡ����b�R�f�k�I����L�ni������䜑BrO�����i�c��D�p�wD�r&֩G$	��mc��;L�嵥���	��#���9F�N:NCl6�(�D�����;Q$e�ȳa�X�qґ6��6�
PBI$��N���lIbE�
��h9��qˉ,�NmZ�I�-˜�RA�r"Hی�7(���D��J#l� Nv��D�6-��R�VA+1��T�cm2w��+��"u���N��N��m!�֛[������,�%N�����R�j%����m9��۬j�6�N�!�5�"6�RY�GH��"Hv�Y��e���:��L��9�P���bmۑG㍧$�m� �=�r��$l���o5��?~�����a��i����C}���f�o�ޢI5��l��w���$�I[�!w��؃���B�ݚĀ7�>��ȥ�{���� !{��1[������"Z��2I#��s����?���7^�'�Y.'�n.�Y��U8�*�N�+PF�z����k��L�;+"��X�⊫�p};Z,���+��l���͉D��%oLo�w�5�����n�ލ:$�~;���DhQ�,�Dд �9�&��ׅ��jS���M����@7�?� w��glZ�g�]��Z�R�H<o�ټ����#7���h�������G��@B���m�/;����~&*��ʡaѫ�K�{ל�H	��b|I��F�۹� ?s7�Ձ��yGc>�7�v�oܰ��<��z۞���&{'	h�;�ovr�檕"�;�Q�	K�(��ooh�6���Lb8����;������ۻ����X%	JBH�".�|HO��4I����S�V�_CyH+s�|���$�'�szb�j��ƀۺ#����7����e���M��cn���ʣнTlĘ���3���[?Ͽ���a(�j(-}��h����2H�{\h����+Q�!O{�o�쐃� g�1�&�6>��T�B���İ>�^kV�=��D��4yzctH���O�MV�~��/:�x�l����(Q�e��D�6���� @����_? �������<�b�j���N�?t�Kh��2)���o�~��p�M$�*TI<yۺ&�D�����D(��sD�I�{z����Ւq�ʡ�=��, s��ska��{���L�<`2H�z�$�D�����!9�,�)�*���(������SB��}�v�3L=��Y4Hɂ�R�PfQ٧b�52q6M�^����w~�����g�Ǵ�_>��4{ t��vܘ�sn)۶^'���05�����׮z��`��ֻ��q�A϶m�s���(G5˵ h�Y8/'t��5۟Z�=s���ŭ�%-;��ع�v��{4��ogq<K��l��:2r"UǍ]���Лv�<a�G�|��{j�p\�޶-�u6����\��۶�T���9��olu8wmK�v���dٜ[�G7�8zZ%��8F^��͹���J�͙e��g��]=������7T�]���t���=M�H���I	����L����g���������\pr9@F��o��=���'ȭ�!���`$��z���w�� U<��e���W�ž�[`�Z��.���$w��UB~$�L̢��3Y�-�p����b@ >=�����mz�� pl�Q9�����ܻ����a�)� �����'�I'}�� �Q&���۸�6wn|��u��i��F�V�����j� ގ�T=6��乬=�!�sN�5D���t`BM����޹�[ދ�����	�i�-_�+�а��tH�l�E�+;g�b����X�mV�}�]'���ʡ��30����=�����+<<����sL��&���щ�iݩU�+j�#&��3�k�)�[��0��0�M��:Y6-K�7��.i���ɶ{%�s;�9�D^����&!h�Xε��c
}��`���u}7mϏ�F����nI$�{ٝ�Q'�@�}�N��y�����Ƹ�ּ4�Eر�Ql�Oz1	 g�?� ��,��6)D�$o����3_cXq�l���Q���s���\�\�WR���$I#����D��m"MOeRv�n3�77KӸ#X��#����`��w�����'3?w�ϵ�*rԃ��i���6�����I'��w�<��
�>������R���pUH�닑�I�Z�t�Gu�޻@Wn�W5U*3�^�Ki ��{����c`=O�2I&��RtIþ��"{��_���c A�g�|�=b�1
h�j������</+sk�v�#}U	��Ǔ�0${V��?��7��7��П��*�2�.�.�Ć�?� �^��  n����R������6P�4D��!E�U�;��
,�Bs���������\ԕv`rI��5*��F�˨J��,�|�.��W2���` �s���xI��}�q�"y����-�b�k��R+3����mś\���Do�:$=�2@4}��G�y�6�_-�.�"�6L��8/.ր-F5���O� ���[=���:�nv=�\���l��${�Zd�$�{��C�Q�f;,��VQ���'�H�A�y�#I�;���r�I���Q�nں��D*I�[�W����j�s��󘵇�ߵ��D���w��<������Q7��������i�^:��h����d~���j&�{}�+Og�X�:$�G��N�$�>�{��A' �{�{�L%�+=��.j.���CG�������T$�D�Uk��; �$Mz�$0����k`���v�Vإ��3�z��U�Cµ��OI���l��o{���MQ:�b^Oy����-�6t�}��I<��"��v�^�v-�Sw�ѹ�!��Q�j�4�j����omU]���vF,/.�#�L��Tq�  	g��7�b��'�QDGcFa�������]'����Wsr=��CusN�4I�=�t�$���6v����<����]���ks�m��5��)]q���x���"�5��U%uKa{���J�Vj5�˵�d�I�}��6!&�'WLn�T��B�����N�$���t�	���4b&	���f�=������s�U�˵1؇��r�@4I���t�� ��2	)��������Dۍ�(�E�/g���&�4H�ѦI$Ӟ���������%ĀN�{��I4N���>4�LB�Z6X�x+��7����j���I�\�9	��]1�MQ&����u��
�n4����Du+���-U�ɀ���5� ��k0:?�,���*$�o��I5D�9��A�Ml֯�9����NZ��������V��U���n�V�H����T۬9,��볨m�w-"��t^{��E2�;������ߙ�5���l�Ͷ�7p�\Y���͍Od1�,[�3�����&���ü�k�Nҝ=y.��U����q�u�;�^l��%�<���#��,�9#:^mi8��w E��m�ᵵ�-�($���N��+�5�nz�p��]q�3�{q�pDk�����l�ѫ)Z�7ݤ$�X��-�406.3g�y*�;�psX:뮋�۞q���ث�t6�h��1�':�vON]=�닐ճ�n4����y�������B�џ�����l>�~�o����5��3�.��{P*�훱������}���p�YU`���[L���{Y�Ү{��c��H�9��I$�=�ZuD�r^^a9�rԽm��-�]��0�d�	����g���[���ĉ�)1�@V߳6w>$�Os���7��ӫ[V��iYL��uu�BT�Q��wb �αW D ��u`DDD�ݔ���k��hD@�k���ޟI�PF£O�o�� ��s�L��`���TI){��ĀD�2M~>�{�}*�U3b�
�갛��뷭��p݄��Wm策�P���/9wA�<�􎔞Ƿ�)k�R�A��@���� ms��b�����fm�9�Oyx�����\����浀}��չT���(�_��%Bh���焼ܞZn���_����g.�{�Q=�;�:�Z���R�;�Z�Twz��k���c����HsD^�Y2Q���lp���~I$�?��·�C��UmI�fw޹P�4�!�
>mެ��
�Y��y��"�f��[�Oā����|O�td�����$�]�Rd�M�{�C+�<@�A2W����F'���o��6�
s]�}��H;��ٛ� s���=Ǝ��_��P4I����$�m-�0e��v	���� oč�}@��f
��A�a�\{HD�=��`J$�;ٻ�\u��]]�^i�P�,��(���������s�V{�ӲGj�8;ab��T)����B�Z6ʞ?!w[�g�  ��f=��'y�l�W����-�7ZQ$���w�$:�*��ˬ$n����2^�Gm�ñ*��Hq&�����  ��m�x�"�&$��̐�7m�����&bfDIRD��L�5ա@�t^U�\6�=G���Պ��œy�*���h��9QÛWۉ_�<�N�]mwx���U��]�0��:���H^�R�Кi���o @�{}�bm�����m1�+j��41�"�R ��XK�٩�b����,h/��� �N�Z�79���}[6�Tk�m=��y��[��&J���!k��יL[du��&�w}w���V�x�n���lت���T4|W����>?:Z��ŝq۳�sˬ�E�؇z*�=N�\��!FMh߽*R�L�/��S�>'�s��DI��7vy��V�2^5J��`�A|�R�=�F���@(W�- }�m��ŝO7,�IͫTI����DV�,-3]�JY�Ò��%#*�
 ��j����7V$���g*"�pJV�O�9�j�O����^B.P���%I���/�&���U�X�
�ۺ� ���"ųMt�u��x��	ћ��ք�)_Ql-�g�Ob��.ϫJV35XkB�u�:�bX��qH둈#b����K`dZ��f��� c�|V֡�(W����&�O�v��Aow:�V����gq�`�b� ��_�{���J�w���m�+��l����Q����`�ì=T�] ���8��O��~~}� �(�>��q �6�Y���vlo.�#r���+��I������`�ÖE�i�g��cH'�E��X5�F�A[z(����'��om{j2z��ko��_l��4�@�m�5���}�~$��b� �]�V�3�\����o�ﻟcܢ��J)b��ƻ��Ts�ǲj��/-�V�wvՓ�|[�X�`�i�B�F__]��1w�,]�b����Θ T�ҫ T�����K��{}�:����r}o��ꡫs�Y����#Z˙�SX�a�����U�3�EZu��o(�%njת��*Ϻ�Uבe����S2�8/�ٚ��ק�����*DR���.�Lf��od�-��o;o`������|w,u(��$��d��$Q�'\��D(6U�WlLe��'Z$\T+ǩ-�Q0rC��s�me�{���+�����k]pc�r�s�ł�^2�������K������d�[�_c��\����L]LA��܈��Ώgv�<4�`�[To��3�GG�pA���[��}z3��j5e��vL�'$J'\f]*3'ۭŔ\��l�)c��	s�N�IVT��0�vf�ٷ�m�I�ˍ���cS�ތ ڑ���2ܭȈі��t�CVg��egY���i�����EJ��(�I+��BeX�x�e<��˻�)�����#���1t#��u�s���h�#�0����U�6���������ɢ�����n0A�"��v�V���T�y/��Ni�����c������Ys�9�&���������I5D7�������Վ&�ZzdϻD|*�L���1V��
'��wi3����k.�Q�����3ᯍ#L�ъ`����Q���%���q�������%C)�l��f����ŃL!̬��׌x/Slj�VŁs��ڌ��]��t��Je�9s*%LT�N��h��&�81:�"LWopBa��ʊue^w2�n��w��n�1�TI�Q�d�`a�y�=a��(,�-Ȭ�ê"��|�&�Am��BK;��)9)m�:p�tP:r�RqN�b�Z�N���gjH�8f��$��"��%m�9	�[�"��ZI�R%���6�Xq�Hvu��%��pRQ�whr���pe��pPpN�H���#��� �N��G(r�]�DRc�s�� �H�vg#�Jq���8�;-�p�ӇJ8.	�A$����9��m��Zq Vv�B$%��!�Bq
"�D$B�#�'$@�M0�\pN$ڍ�$��'�4#�rI�p�(u6�"��q0���s�2s�����˫��{m3v�u]��"c`콭��k��ny��&��^	����#g#��DZ��ڨ�vuy���<.wf;c���#jݡ����Jm��p�۲v��[y�շ3n�}���r��g]�ɆB�ɪ�[u黎����N٭�۷3�ᡣ�z+�����]��v��p�僵�;7�<�1�Mӡ92��M�WtY+X�F]�m�;��G�۝�5\�z�wW\l���̊F���>�3'ly$�]Ϋ�wn���b�d��n��\f��24;f�z�9�$�f���U�_��㰼�v���n�!�/Iu3��׋���6XScM���.7om���\�أ3`��8�q�m���M�w:���f�zp�]�=`X�nt��8�g����{��科�P^_W[j�{hѪ�[�sY�C��12{i5���p؋s�.�E�b��nS���n����jp�6(�k�����9�8���籵�狐�ɶ�aN��`�@�&�,4�ݨ�Ǿ v=�t��yC��t]��;4-��vV�`{ne_A�\�����сu[�v�q�vYO\����&ƙ�t͗��:ư��V;��OqȆ�vwE��Í��<m�-m�m¦ywF9���v�s�y�c�iRܝ�N�C���L�os��v���f:;��;�'�]�b����ˍ�Mc{N�<P�b���w�Y㷜u��d^s�a�R��l��z����������9��ˍ0Ÿ#���mq�7s��nOr[�:ے���b�cX������c4E�<:�^q��z�ˋ��M��\
uvɷg�n�s��ۍ���n3�w8�a%ٸ��xs���׋q��[�q�e�-+t'nq���q���c����R�uiK��;c��� ��a���ϵ��ۦ��ts���`,�G=<�`HěL�W�kڮ��N�QU��J�\yή�.9n(��/<3vBقwA�d|=�ؘ�Z�ѼYD�f�D����:v�a���.�P]��5b�&�N�I�c�����c�|�<�mU���HŎ@����k�q̬g]��ٻn#��K4�X-���c�v�"�h�Mz�9�\�A���Sӱ:���]�k�����l�a��<ax��g�3�cx�+��l���۞�k 9����
��w���n(�g���Epݒy�u�<ܹ]ֱF�``y7�Dnk��[��d79�g]p>ݞ#Q���rNvٮm�[�{gu�ń��4ᝑB�t�qs�Apq�YX�8������!]�"H�(_�%�ؿ{{�Œ	�V��ua���u珛�o�ܛ��$8I�е�[1P�v��7��ߦf?.�:���A�V��U4�]�+�O5��Z	���	$��0f��]N��6��V�^�k̨� >��/�	�b�6��
" E�Ͷ�K���vv}@K���X������;�SչɩSm�{�3ۍ^`풊X�314��R�7|�:B��;��%w�,�F����*+�����V�=d�mk[e> ��C��u���U���'/Fq��69�x뙻rۃ���#rК�_�ҡ�<���qY$��Q$����K��q ��!�R�3�vłO���@��c�0� }!s=�A�-����ŵ޷��5�p�h�z͕�Z�F�w9����6�kl�6U,M���f|�[綇=c�[V�<���u6/��=���|Z�HP������$��}����8I��k�^� w=N�
 K�K�R�G�q�I;TA�n�z]�$�VX�Nf'��s�ݛ!&�5�����d�ٶ�_�����k�;�7��4�nA�B�0�7�6�|H/��ٻ�u�43<����[5�H=��b�u�s�[*_v�q
�*-���-�s�mxә�[v �G�2��ѝf�������P�	RA��D}n�A��۰T�0�Y�{P����D�@��w�����(Ԑp��O^�w1��Þ�`�[�1�I �om������Yñ�x���������[��H=��vA ��ǻ|Lz�vl7^��OCdkdn+LT*��K�݇;X�]\j�.o^����"1�����ڜ����(m�]�rt��l��߼�X������ ���۳zm�A����M_
�r=�Wp�=�g|��VH'����~����˳v�N���2��$���D�7`��wg���[uI\�b
ˊ�ҪA���I{��c��wlD�7�o8 ȓ �T�G�tuځ����6n��6�$��\/hu�S�͘o��ۃ��Q
P �w��;�I>/�����x��}���(���(
�{ΪϲH\q0�J��]���j����s�H[99�Ē	�u�$�8�P"M_e2.���:�����A�Ǝ��g�b�>�v��J��$5F{��H����A�v�׀�F��$*�v���(�^OX�LooX�>Nm����~�ma�9��f\�ux��Z�y�{�ZT���=藍͏y�ڝ��eX��4Z��c�}kv��DL��Ԯ"�_o�DN��U��F����<�| ջ�S���M$�hZ?8���A;ʰ\t�:��`��7Ω�A&u�	��v]�������>��	�J��0�s�1u�}��kt�m�mm������k �=���P;�_$��I�gx����A��]U����磵���(7���~׈
�"����IRH��-݂A�,w.�R��ng��'ă9��}}]�d��ίz�m�鏶�f��,�ˬ$�\آHvP�E�tHPT�F3�/�z[i��*�o;�o1�C�0w�!�N���w������$����I̮ʱ��v�g+��6B*�o�$׈mh7��JB����|H�{�]*p5^�I �T	�$���;������>#{�x��x����V��Ӷ��
�*Z�Aœ,v�󨪆����\�wf)M	k3^�1��U�����*F�8t+y�u�_|��:�1�uP���nw<u�oF����&�v�N���j��4[d�a�%�,�Ax7��u�"�f��*���ޣ�k��}��In9V,J���_���=�]�[ǎ�mhړ��ɲ�F|�n��m�r�ALm�9��9v͎�D�˻K��](�q�ݮ�:{#a�������*�2@�+tM!����x����b�(�t�+3s���k=��fY:�Z��cy�NC���/,�y��7f��Xڸ˱����Gkߟ�~l���������i���yV	$����f�J��S��k :�@�/6��xv��R�	!&,tOc�X��٫�<(^+/�� �ݷ�d����g�4lUZ
�����!H@̒(=�w`>��;=����g]��TH6�
��wl�"��0�J��U�E޳1]�1�`�صаO��wU�HX�Bރ|V0vsn�椵�/Ď4��o�X���k�f�eB�=[�_wO��wV$���V;T��{ػ̋5o��u�DPuX�]>�.�3���.ɗ��lD�'X6��� ;%uKas{O݅�R� �+�n��|H=��vH>+�P������z�&o7@ '{�m�W�M�@�*s��C���eO�����ɬ�N�Ayc|���c�����kA{QvS����H�yg���xR���1���.�f����Q;1����{�z����}�d�J�j� ښ(�6%uU`�S÷>R��IA�3v�\�Y�+'<T ��Y���
���u ����`�V;T	B)DB�H3$����:�0D��%�LO������f��圇;�y���ֹ�P� -�ny*&�t=/�>ɴ��v�W!D��v]���HM�(�+��H�2���V���;\s��\�qZ��ؒ}�{	JQ>w��_���z�w�ƛj�u@��/�]�<��s��ݙwN�ī�կ��;
X3�՘�߹����+�_p��r�|H����,�1����	s����0��b	^��C<w��0*�X�η�^ˈ�!v���b��.�b�ͷ��6�h�IK+p΂����iv�csXڰ���5}w5��*V�f��Y�<��wFN��]#qv���x�����'�-�@�/�����>R������Y�\�+	7�	#-�A>�N��I'{��仛���&mRrDR2��(�fI��1ز;{zźo4E�϶���|b�P�H�]wd�{�z�qZ�l�����mc/��T�F곞��I�luђ���,�#P�*&�D�))6����t���Lg�/z�'���w�z���GGm7\h)zb�@�o�]߉
28Z�Dܱ������b�s;}_^�i�I�]w`�N�oX�J�Y����I*���aD)S=	�+9����w��9!Ndԫ"�;�� ��;�$A�{�ōk��M@���w��g{�RjjӲLs˫�$�s�z�ĂG��մ9��ER\�N[ا]�fwL۠绽0[5o�(W�qF����c����:^�9�s��g+�U�K,Mz2�ل[�]\Qsra�8����wE|���_om߉�ލ�!JRe%*̓���Y$�:��H"tϧ�4�V,w`�@:�y�|��B�n�^�X���0��Hh쭥+��:롮&����eǗշ3Gmڝ��9�@���f9DD%�G����ޱ~ �Z��ޘ�ǯ+h2�볁Ttܡ��X�$ئ�V�߅y܎���F>޻ �BŪ�H.^����T���!i�j�>2�����~� VvjB�X.��-g��t ;��?����O^�7�P����~ަE��W��D�'�o-�I��U A�]�[;xa��6��9�K5�O'��F!S�b��:'B��X.�g6q��s�$�V��/�e��faJP2�*�]�5���30���)דb�F��JۚL�׺��)�'�����[}�`�'$�k~[�|�v��H����?}T��qh�tiʥ�U	�7�[t:5��5��m�c	!x����g�u���q���:�ǵYSL=G��K�GmmW2�ɺश�j�u����H�ۈ���vv0���qx6ͳҖ1�=qD
���r���d�:§51�K�N��s�u��j.vM�ll]vk@a��7=���V�<m�hQ��N}�!�%{'���x�t8�	�fM���$|>]��Ui�j�絣����FS�T=g��Rl��e(ɿ�����Y�VM��I:��ok����7�!��M߬Wu* ��A�3$DIP"d�A�7vI�I��D9�v�ذ|I[���|�~n��<���-y]����}���[30� ��_c�W���X$E�����C��n�Foh$
{J�>�{w��S�a��M�/�C���W�9&��D�$Us���w�`OwwS�U1�4�w�V�Tt#*R���?Jy�,�۽�n�ZU/�b�A6�Ne_XϚ��bͿ�)L��n�����R;i��v���F�'g]��F�e���ۮ-��iS��Lg�*" �c��P>;�{W�I{������M#����m_]�}ov�壶����Oo�{�e���x׭�"��f��=��%��!�3ig�_�ӛ�{WN٭��p����ؤ����I�͢���^M�Ea�Փ��E���L�~�� x@��_x�Or���w��b�/���ԛ˭<�Z��g�4�IJ12H޻t� ��W�AJ	w�f�Un�&O��ܻ�ww_����9�3�7퓳�y��ui��,ڰI$���	YZ�ʄ����ӳKh���>(wR&b"|eA@��s�(Y�UR����@��19������'�ej�ec�U�1�D( ��ۮH�6,Ӝ�k�w� s��)Fݶ�	�گlqs�OX���eJPcА��]߉�۽�,P�.�1�y�wEU���n#}B�/�xI#��$>7��3��߻�ư)Ju[�|H%��S�B�b/��oK\��>���my{{l�Z;BГ�v? �Y]^�	<'F��x�=��&wHxơwhD��j��[�)Mfbl0�:,�@�<y+/$9�`64��u��ۜ�_#��r�u�1���������v]��Q�^+�8�e���ݫ�؆�s�N��� �aC6+:`�:��{ݹop���6��x���	�ZZZ�n˺�$��낞��Vw�:ح��>6bpo֮��v���OT�\�?�d��Fd����O��\�-�{.r�X6]p�'���\��պ�DÖ�h�W�l��7��w7H�����2�),Yjp�����1�]��W-(��ZK�����9vp�n��{r�;u��X��'ڸ����,1msY��@Y�Y��r������[܄2j<�C�w��n;�(u�RHF#%��M�չ��o�o1+Vȳ�g�j�C�M�7+,2�B�&������C��×��أ�ËvA��CC/�߷2�ٓ{j�(5��XcX#m��Dz�����oimΨ��I��)Y׀�|D�p���v��ms$�[*�R�T��~@o*�q:�ڶs"&�E7>r�#{ED]j�A"�ׂ��0��
Z����&&�PVs%�;�S9g&��Dk�#ut��_Y/5_#�-<F�F���7y���\iB�̹z�xjT�#Tߦ2�j���z��\t�7%�#���ڛ,w9�9uiꇐE���8�R�.����kvs����kf|�M�ΥFۣ�L�f[����֐%�� {�����&-�C�f���^�J�7]ӎ�v��᮴K��tWB�	�.p���'q|iΜt�:
B�(�7H�3�F�۲�ʎD��82�8��4ڳl��0NI�j;�%����
�l�qmnij��-�v蜊"��qö�Y�8�gbIhV$S�nlpN9�II9�s��	4�Fr9P�K4rq0�m���gk��'�e�9	I�K����fg��m��6�-��0w �p
'�p@/{׎�;e����y����y����^�����Yff��^�klm�v^�kkv�L��y�D���I"����Yy��{ݬ������$�	7���&@m�`�{�o��{���-�Tt��Hđ$#$�|۵ǳ\�Wt��X�	$�\����뵹�1��+�A �ǖ/��\�2D��b)Ц�b5���+����c^��c@)֯U�����=Xܭ��Lb �	�%�0�u׵�����#�㵊��vۜtnT�'|���Y O��S�]�������4��|��tr���hy/r�@|3'n��m<8+)hϋVd��f6���)�=��wY�Rz�ok��㑑yږ4�{Jb��9�,���$�T_eQ��n�Y>5% ��N�1ݖI ��W�&����^�Č�(�Pfj�Ms�>��vz��A*�Qvu݋5���Iw�"��g�M�H��ܭX�vAW&y���[��z���K�#*5Dk�3��M�&�����疐�Վ�&�+��b5DE����t�� ���G��r�$��!�$P޶��I �����op�Z�U�I9�ww�I����ˇR{n�T�%ڝt��(32!�5ɵ���1s�3pF��i݈��#fV��1Rm�~�Ӡ�Q�&/�v�@8��I���n�g@91X�;��(��Wo6� ׸3Ywd������<�y�!�^Xx��}m�ؿ�ݽ�,;�Z�cq��`����l*�����d{w��g@&��4S�j� �7]]��v�X��2�����2�@Y{�qj�,�A ��ʲ@'���u߉JƯ��
Ȕ����DI��n엃#��-�+rf?M{���ڗ�֧!x�Ώeh�c�r��N���Jƫ�U\˅$΋��\q�aBAI���2����l�w9���j�xz��my���31aas���_�N�%�}#)�+�g:T˯W,�(k����N������<G|��2�Z��,�s<�ɓ6�:hWv!{A��.�&�<���՛��Æ�%�i��2�,�]Aw/]];4�v��n��\��r�Zu�qm�T�����.�A�\<'�d��3c� �ܯ5��m�@�X ��b�k��煺�lƺ=����+&ڳ�ݵf����]2�X2�[��\GX���b��_>�[��t�V����ϊ\x���`��λ8ᓎ��]y b�m��d��t�rF0�!�s�tJmk�BY+�7�z;EX)� ������̒_wu�>�+*xJ�b�fڀ�C��v	$������zp"`�1��fk�D�c�ME�6��:�I��v�m9wʴ�}�˽����B|R�@�vm� �D�ڣ�Iw/0��6���H���v�2��$u`5������]�ż��y23���]�,��Yʉ�>��[כ�,u_q�m/A��v��)��eL
�Ee� ��ɧC�jߔR�,�&�lP��@�H�껰��g#a��p0�
Q��N'��j2��Kk�O>��nD2����v���LwB2��%�\�:�H�Ϋ�s���-e��R����r{�Ń�L�j�t�ܔQF O�L(v�wd�]C
���&NNB��.Jʾ������KAQ��]�l�e>(ںs���n�g�׼he[ dÅ��Ys�י�P��js T/;qP��ɷ���w�O7������,�(�H���1vFg:�	-�]_��׉��^�} ���$�[��#s���i6b�ϊQh�vn���S���]'T@'ā�՗dݽ�yT��u��kcA'w-P&փQ����	���$�����
��e�մk��@>�+��w�NO-���5��-�6 G.���lH��9@z�(Y+�iWwl�<��A�>���& �dD0x���(�W�I�;��B�䫮&�is(\�7N�Y�.��h�U[&/��ƝZ���w��ڂ�դ���u~����~��&�J���f�0"�1|�Dz�ݶ��O��o��t� ,y3<]�{x�&x�V��υ_���Z���f���j�;%�C�Q�%�|7F����>q��V�C&�횬nx���4C۬y��q"�ӱ`�ݽ�d:(��`H�D�1v�lNV�Kw�i�Ο,����H�{�w����{���͖rOw��(�Pd13�����X�ͻ�W$�x��Π/���
���:�@5�T
j=sN3\�n���W����n�
���]���뛞ݳ�on��<���Z�WI�Ն�~~�g�~(PRSD$+�[�v��d�wj������Q E8O:�:��Ő7(�& �H2�D�T�x�ƥ8��us\�>����1ݪ�(Gk�V*qM���"��2�0�%M��\��$�whPq���7��$�w{���| ��*��j��t~^���y�w�7�H2����D�Ggc�𧼣{�ٝ�'��٥�������rR��f��s��3f�EoAϸ_e讐s��浵�om����.P#V;Ƕm'B6����W��v������r2`H�D�v�У��Օmj��v�E�}ɿ6(^x�<�?�]��\��s�����2��ݮwmA��`J�Wj7	����m���w8.e1���q=c�����y��4,����O�g[��G������9\��?�O��]&��y�"���h�f+}��Q��]�X�l/K���9k�@�ηW�O�xD-r�Wf��
>t]0�d�����Ǌ�'���1O�Ω9��xu�ՂA[hQ#s�݃Ol^����U[�Y�׸M�U\G��J��$MoP�I��wdw��M�׵՜��u1m�^v�%��]u�����%ݶ�����h��l�k� ��^�j-�
 {���着I�ڶ=��&���'ڛs��D������^{�<`Xǚ\�:�6�6��3f�5Ò��%���)��^�5o�i�X�m�fz$�mvgpKW\��	ؗr�m%d��=;śMḾ_m�է����Q^0����Z�lm�HV�z�y������a=�k�A���ilz:뗝���Ak��u���Ix��݋6^�xy�|�� Gc����/U�G�OumOٱ�q�k�Z�<s�OmF�6�W��ꐹ�K��=�.x8�4�����^��s�7�b�g0� �x�&'Gq�׉�v�7m��#��[��
���1�>E�jj#~I�o}��m��[��#����J�]9�!ͫ������Lo�O:C�V(���ss�d����<(�N=�w�O��{���Y��i#]�ɘ
&���v[�v>$��,�웅�j�H��B�$k�v/ă���,�Ytd�
D�S!PNnQ<e�]h�+̫�A<���'i�o 8ک�g�;���$&��0�2��ǳ�[
��e�U5�0-�f9*wd����X�> L׋��\f�dB�;�>�͛���Sk��']v��-���ݦ�۲E�R�7g�k/an77��|��!D���v���K��$�N�K4�.�e0O�_wXӨ<mAEeB��&����>�ou�K�o�uumnx���MkaG�;ӱu]VU�y�E�3e[bР�ۅ���z��,\c�5�X��z���w���3���6e�:�|C{�VO� Ÿ���v��8��Ʃ�"m2�(FѮ��H#m@��Z�=��E抽����i}��,H9T��E��#)DAFP��6��NIe� ����t��nR����4��� � ?'͇�v��@�
bd* ���|O�nӫ'b��y�d�ҷw�I9U��$�u;aߗ��j�`@麕������K�V�8��V������9pq0w<���vP���������D%TK���u~>�^�	�ΧbV�ϗ��O��7@W�� 8�s�	5d`7*�>�� ���]ڮv���
)�B��yv�ᗻ4�Mcʱ�K�1�9�d�R�	~μtI8��Im����=ͧc��z�N�]SW��t����Cd�5�|���F+r�ٻ7Tׯ=m�_r^�x}�����3/%�|���V�&�,5Λ��'<_���7�=���>Àկ���5��x�BWx�ʀP�2/� �y�N��ڰ�y�bA ��T	�n&���(�.�5���ov߯�N�X�]��+H�ז,�w���s6�{�0�7���i��5��Wck�\F�	�����`�n�H�8�[��^^p��I\r+���u��'�o*��'{�jʚe��Gx��W�ӜL9 �VVk0VLyy���q�Q�|¬�d��yVI ��}�=hc��]���R}��&��&�����vH$�om�� �y�/�F��ԗM�^X�H=����a@�M�X2d)B���x�{q�ڻ��F��#��A@7y�Q� ��4��FC�����[2&j2s{�"����s���V�Rjm���"�^��7��!Uգ4+)���C!���ʼ�)Q�φP��S���}�r��9W5��.Cng1.���07�^Q��M�-i�$���|�|Ѵ��^z����D�4�Q��{�"�]=���}���m|�����f�6[AiƂ'��w�����"8�s{�"��AS��|��޻�VP芚��(���Xuͮ;��M��m��8qc�R�4�UW��t�r[Yr� �bb�｢�`��A��J3=��-�؆���9��h��������֏��a�-39yt[Jڍ(�iF�3=��6�����ޚ�G�|���e4N4?��Pl{b��M�[��S�w���Mq���{=@m�l����ߩ�6b�5Zީ�k��߸v�(�GF�����#����}	���-�3ח�alPaQ5o}�c[iF�#�rf��}s7jj�h"q��C;���r�Gs=���?�>���>�����������G���(��;�| ����PiF{�稱�؆�Dh����Ѷ���=�^Qm.���糵����9��ixj4�j2������FMpq��_G���h,h~�;A��lC`s���wG�{��^�?���O�A}�e�X����d��t�ki���=�^Qm��z��	�����~���ˌp��pT۔�͙1��5�#��u�<�8�6�1�4�3�e�z�Cw!Ga�ƅ,�D��@©U21kV��Ҧ�)��
�x�kK�-���ؽ��V-v,��3]e����Ԣ��6�v�9x��㊖�6�@]���5tw:���A�% X9����T��s��7x嚍��ҩ�l��Q�aNrun��	�&#2�A�e��Mち�NKF�x�6~�xx��6��=s{\�$q��G-`�ܫ�2�R��yM��b�ƝhN=�Qk^��L�{(É�,`z:�5��N#I����@VB�P�.Z.o��Y_b3��x���6�����Y"B�ý/r����}�Y��4Y��wx�����c	jђ"8�*�{u7��^Nfʷ��z�yr�c���^[s���,3���]��ۃ:i�j>���wv�(��U�a������Pf\���
�^aµ�kC��Vۋ�lj-�Lob�����f�T�JZZw���D30�@ʀ]ŭvj��]�x+��MC��e��5C����ذb�56L����gjҹ%m�^Y]��T[+��'[o�^na�(+�e��@�).�o,V�W�������fbu۸�[�὇�R�ع�Y1��,���\����"��n!!
kb�"�v��_"!�Qsַ���<����[����P*&m�C],�j�	�u `�<�Yf�����:ԣHmM���(|�tA9������X-���ْO2�'�n���ej'����"��z�t��C�,��6�I�9r:�D�QS��;�Nv�-m��R�-��s�,f��	�"Slol�����9N�\�v�
��{v�'��R�����kӜ��m�P
� �̏kG���h��Q�y�k[F�N\����kP�b����w�bB����m�E=����%�<vHy�=�-,��Y���He��,���󽝡�vq4lvYٜ�m�מ)�',�׻C�i�ӛn8����Y��m�w��k{e�hMd�3Yu��Y�։3�z���6�A���Zūo,�[���֍���~o�Б73y��I]�s�ٮ]q��nv<Ֆaݸfn۰�8,���`,���^n��/�<��`��j�6��n��ݱ����ɹt�m��*ɹ�����n����"�\�֖77c���棚:�]���.�-���w"5��5�7TlD��0�xn��NKd��m۳�dK.����C��T(vu��u�w�v�N�;nn�q�2�uZ���/�����k8ܛ�r�L��ZC,)ڎy�y�t�=�Eѡz{rZ@�{q됧]�c�0�*.�g�=��gj�=
l�	,Zp�sm�v^�{k��v9���m��Z�84�(G'���㺱��t�;n�7[�ն���c�{��o]�ϲ@APq�9��2i7kgy�@>��砎g��ռ��<uvֺ�F�pלf9W��;gˆ���[z������t:1�9�z��gB[%Ի�ĮC�G^gY�|��8����ӎ,V�E�)0;g����Uٗ����������2s��NM�]��l�0苝���v=��[OK�]ՙG��'�A�<GXKvNk���<Y�(v��v�9��Ɋ��\-\Q��{:�Eˊ	���eK�^�g��7�c l��;\-Øz-��t�6]��8��.�k�56�]��'����-�m�S�-���wkpӑwhu�����Uv�<�Cط8�������1�v&{V�<��3b�+���۶��7t�碧��H�f��][Q�]�O���l�KZ�HA9`ȧ�r{W��=�r�veMc�y�9���n�ܘ���<;Ok�t�rP���t�:��Eθ9�6:�m�<��x�s�'V�Rd�9ݸ�mnu����r�ι�[���9����o�{q��Q��<M�ؔ0[����N�6q���f=tr&&� �[:;�������۬���{�c1�����ݸoeW]X}��v��]˹��ݞrW�1��u���{uN��%��;�$�{4nw��Kl���7ks��W{,�]3v�v&�a�X^�5�*/.3ˤ��ù�8�JcL�P-�]��:��g�`u���h으�����<��[��������ٻ9�!��tT����p�B�t�_e�j���s|w�ۭ��|���ڞ.<s��]�Y�SWQ�u��id�^�]n۞7n7a�nKi\=���z���{.��#�Ë��ζ-G=;nꔉ�M�qcgqf�{ŵ�7k���pt���i���]E��RU�)hO.���k��EE��V�+���~L-�&���ˣc[i@j0##�^l�!�=Z�[����b>�ϫ;@]��n0���E<$4o��vB�-��X��[k�����ҍ{\��v{����%�3�^�ح��D#D��oh���F(0�Q39��ұ5Q�������h����������0�!���>QeLѲ�����m=�����F��4��F}�}�}�����ߪ����80#�o�H��4�1F0�s9E�Zh��S�������������>͠o϶b쩻
��H��4�j4=z�H��ڌ����3�-���A�!��������L�<!�a=��H���������s��hMC`6l�ܿQl�`F�ҌCg3��,��o7ZT(ѱ�4@����LCb��1D�����6!��j333�+L��������eU�s�۲�H�����>Vn����VG,�U�=L��"������x�LqX�?-������)��H"H;���"1Ƃ333��l�w�{�r�X9��\~5��Y~�S[Q�b�"a�s9E�[Dh��nA�a�>����YY�l]�̮����~�sM�y4��]��Hl��.r�:��pŶt�#)bӣ��*���e���7@�>���Sy3A\�Vt,����o�����H��F�9��m��q���fg�.qA�凞��Ԍ��[^p�" ck�)�_jkSN|l`k}�(�؆�6gsݣ��h�Dh��4�k��c��sY~E4u�1F��sܢ�V��(��JFffz�����Czi�&����)�mU��W��[�6�#��lFH}���"1Ƃ2���h`F@`F�������Wy7�f���m�l,aW��-��#D/)�s�CZ�Mm�m����X�أҍF���Ѱkm-v�9Y���Ü�y^-0 ������Ac�b9�g�.r�	���)������64!~l8�q֨�X:v���/\E�����t\�5�M��K�b������k�C�jf1s9}��c5J5�g33�X�l �#Dh����)��| �O؛�S����r�@�=�J��0�hj1����g�V�[sc�s\�֜�m��;��m�lG�y�Oy��`Mz�F�A�h#�A���c2�=]�E1��a2�y�9��G�t'��G-�4Q���Zk�}
G�#7�~����D�4��h|�]"���6��o��f��E�1����H>���hn�f*0����ކ��;���YQf�m��y���3P6��P����Un���1��fz�����?����|����ѵ�]�K	l�5
le�/���-�����wO�9*t5���J2��t�[bC�e�)�cDb��b��s9E��팭�m[K�Q��3��V2���t����M}���)��q���v�LCb6�=�r���\�_F���4�6w�Pb8��2z�t�kcJ0��0������6�˱󽕧��&���s����-�n�v^�$K�1�k����u�˝=S��pյ��9�߹҂���O�/?�����v�����+�F��JFF���h-ƃ���kG	��9ܼvoYlF�7��h.lCq��n���F@�y��>�7��5�ٴŞ���e�#PQ���&��vfn�ԣ>�{�<1[؆�'���)�l[F(&{���m+j4�j4�w����*��٬Zeg=�.�-�lu�k��G�i͖�[�/���{b H"H{���"1�l�d�_��WU��6�&d`F�����Ɣa(�&�gh��h�g��Q�}�H��cDf�/(/�w^�}�7�\�i�m/�Q����"�[�����F�h#�Cg�ٔ���=��c���؇Di<�=���G;n��˦k*-l7��^Yv�Z����fSی��)��ɍS2&т�1l���i޻�{� ��N��H���FN.�-"��#P�[i,��������iF�4�3�̢�+`�����{�o�{Ch�]���6���1A��{�[�V5Pj3����[W�ys������zi��
�p �S�[�\Y�mї��dk:�iWm���G���=G����?�&��L֌)��Ƈ��{b! ���sܣvAƂ1��{3`[-��������Ox�&M���S[iFb�"a��9E���������CZ�Mm�cDf�y�alQ�i]ߦ��u��Ej�����km(5���;͖�[�b3=�@m�wG�l�˯�w��k7��S��2�;��ω#�����le��m��ҍA����-V�6�4F������������b)�m�0�Q3��r�i[Q�lCg�ٔ+e�'6T�5��ABP�1c��>�{@KH���"�w[��}����A���&�2.wٛ�c2�d�v��/���f�e�������Q���Q�[rm�C�m1������؁#��벅�}gޘ�<����:�p�y��������h,q���$=�fPpC��'��H��h#7�O�=���~]���V����P��I�r������=m��9�p����SOF��h+:��{��C��K��S��f
b߸��_w��Y�'m*	UQ�qU[�w.�:��.�&�]�J�:Aw\���n��[�̈́����B��-�>���/����N܅��v������G�:�M�Gv[��n��;f���8t ���	s��͋��MǭGc��WSz��{qֱ��u�nڟ`E�R;e{q�s�ڱ���WY3�֍Ҫ�Z��u���bqug&�ͺ)by�:60�mt�:���":ڮ3�k�8�u�v�goX�]����i�����%'kZc�ǀ�1���r�e�#PiF�Ҍ�{2����D#C�v�Ѱh�Y�8Ur+v�c>���lCiZj1��fP����������s_}�kF�h6�C�~��؈H#��ھ���F�r��7��Cq4�gs3`[,`F!�OWn�LCa������Gi��v��a�e�~闯�5	����m���v��[aPj4<��km(�b{-���ٽx��U��h-Ƃ8�BC�����("4?Wn�OcAk���s�H�?���6�.�/�[0��O�5��}�汥�iFw�~����m+�H���F(0�Pe�3�[K+����w/Y���cK�Q����s(V2�>�� �T3&,a�`�״�lD$@;�g(�߉�`��-��FE�g3`[-����t�km(�Q�aw���m�T���g����1��N��E����9i����a���p����iDV���������vL�C�F&�����alPaP���Fƶ҃Q�#]�se��ϝ�z��}z�L�}Y�#Rs��˂�#�	���)�Ɂwd��J���B�F=��:F�����@=����J�{5�wϷ��%	׺;�k��v�c�5�FWi�4�9ɧ1��ly2$SC&j�ǲ+N�Bs��>M�^f��n���m�4<�]"�6�����r���j4��~�+�-�����G'N�@�$�D�}��4QMG���m툒���r��A�h#�er�������=�7�G���e����վ�)���aa]�.�h��4J�Ś���4ᯓ�E�����֝Sֺ<��{���b�����ѱ���Q�lr���m�4�!�3ٔ����;��5F��PDhu�n�Omh]��8�EL� �$�K��;��u��A��J3;���o��I͒�����K�M�>�mѱ�1F����E���ҍF���{2�l� �Z�X��9X< �A�%b�T�����]��v�c��c���
��f�����ېgAJ!�ɏ�>����h���@;}�Q� ��7�3��� �0� ��ߎ�v�]X(,�>^"��S[�b��6�m�gOq�
��>�Ф|Ѷ�̼�����A�iv�G>������~T�����C[b20=}�(��q����ٔ��G��m��zMk�ϽUH���"��1B�*fb|a a�=��t[ڱ��(���(���"~|��3 ���X�'T+��݃nޔ/�� �V�r�Nh����Y-l��w��2�{E��ƕ¯&�D���p�2E��`�������O�h�Pa��{��ұ�ҍF!�������gt��c9��i�F�h68���߂k�������q��D�{��7d��Fw=�@m���0#Pg�����g5^�})�Υ�!�%g���q�4E]8�R��SO�&�m���v����@aP~���b��>�>�f~�2���U� `20!��͖�[�Cb$�g�(������v�F�����}3_5�ף���Zw���ܧ���s\��d-vwl��v���]d��BJ�����δV�#t���m`���;E����Q�Ҍ�fe��#Dh��v�h�Db�n�����|�/��Q��Q�m(�fg�(V�ls~{�s���|}�G���N4>@X6G�D=�f�=G����B�Cb�{���M!�W\�
Cb>�f��{׸��(�E����d�	�}�H��m��^P[b�҉����ߑM-��ׯg�z���s���_/=�Zh#�DR�̠6�;�#��������;���L�S3>0� ,�#�k��o�U�s�Q��Mx5��j(����,b�b�4F��w���lh�Cb����(���߫<�o\w��ܹ���v!}�7M��z�`����<P�>���9-J����T|�U�=Ve�uA�)��
�u}ot�_guϻ��b�,j4��g)��=�#kvI�A(�JH�(�|:��lD���7pDsG��Z�?��oe��A+3���`F!�>��H��Ҍ#a��Qm-���F�o���{�>�W`�U�����ٺʄGn�9�Xk��|յ�Ԏ�-eA9c7�~��]��3��֌#;��h-0�(�1�����J5d`E�f݌#����7n�]�N�[�G��w�t��A�����"��͞��q���q�M�5�ٱ�=�z�e�#Q�����e�z�>�{�u.�{��@m���Dh�}���M#L#fs7�-�`�iA���}u�>�5����_~�[��/���I��#"�UG	1[�7yH�#���w��Q� ��h#���|��5�k�l��hs}�S[iF�0��o�[E�F�������	�}��|Ѵ������W�U3��X��iA������i���Q��o�m�m�1H{=��5������ǆlChw���>X;�iL���(da��yE��j4�Q���z��{Y\���g���Tэ����"�64F(�0;�o�m�mF��(����z�t*
��y�~�ˈ-&����]��t����'�r�Ԛ�d/-�3�ƪE��[ʹje���-���Wք��ӳ�m�̥M��y���c��jVJ[����m��{q�Q׆��w��y� ��*�Cmk�8�&˻g��F�3�˓c�Q��έvn�c���sVx猑���l�)����U�qQ��vM��x��׮�۝�F������nx�Ύ-7Ad&�C]n��Gcl���.g�)�:���mvl�ޑ9�ɍî�=������{�/�1��ّή�.K8���bb��7$h�Fcv{k�ޮ4���[7Q��gO[��[W-��	�J�D���'Q�	)"$|(��`����	B@3=�Q��#���d=��le�f��w��w��Y�c\>��"��Ҍ#a�o�[E�F�����\>��i���-�lˬ�F��vY��=Ŧ���T[[iF�&F�|�lCh-�"Hf{=@YpCbߌ��}�ӛg�g�|��|�Hh�j�j��#t�ēf�,���-�mXҍA����1[Q�Dh�v��}�&9��~�SG#a�/;�Qm+j4�Q����z�l����NsN|�>>�SZ�m�4>_=A�s~oZ���Y�1H"H�}��G��Fffz��-������ME�{����3&%�b�#o�t[�-7�snL�Ch��cDf�/��أҍF����6����\��f?,b�+;��q���D$;�g��!�"80��k�|2Qџ���3i#(����`��l�>�W:{����q��n�۵�ۉy�����S30���� 0����t-�0#PiF�Ҍ������؆�	��Bw��Dx=�l������0��gn�i[Q�Q��g����� ���&����b���>�r��dxD@��ۿ��	�KY���w�l���C���p.��FA�@�����ѰT����6f�f3a�n����ɘ��g�hŗ���u��׮& ��O������ph#'33��c1�����MliF�0}�o;�|����"�Y����!���q/�b��Rm�m���h�X�4��hs~�mm����}z���Fw;�q���D��{=@]�("8�/3��i�O䆏�괹Eca#t��"�G��}C���?j_^<=�� Ȇ׆�g���E�[� �$��͢�64F(�0=��(�K�}��s�}km-F�j3+����;�{Ԝ�����74����[��̠�{b$� � n�n���N�t�.+�اb���	0�FB�=́l��j�{~�S[iF��g3|��-4F����35v���ߠ&��
�j��mכ��dpz]c��1A�j�������E-	Ջ�Mb4ϡ�14bh�߲�@m��F��+}�i���Q�l	���e�?SB���ُ�T�~�<0D��@9G	��R)�d>�>��Z֧�kJk�`[,b���e��iF��ɜ骭���k3ޣ����#Dh}��LCb��1D�s7�-�mF�MF�z�+��L����=�ח��e`��vI�AP��,Q��`��w��lDR�������Ab���f���T��m�v��_ܐ⢥��0�9XLw/2��%�oC��731<ک
�p�ŽrF��Y�r�D��啡�'jF�U�N��ݘ��M�w��f�:�N�^���M�l�>�*�4gR�Uh����z��<�+n�r2�1N���\u�Q���9���۾�Ү���gI��i�a ?��`emF��1�pj,�����uk���-��2����;�Tls_<h}2�;^$J�Z�f<�Yq\�K�F����9wX1��L��PqgI`$;F�]���d�u&sH����hېm�e�N�ni�c�Kgnn��˵ݹ*�s4-��N�-��.�ݹ���9��ʪ���n�'���^j<`�&.�����i�@�[2���`Сp�K@�='4J���7,]\��]��LW�s�z;n���Lgb�}&MQ�a�|��nm���x�n#k�F�r1b�ż�w��4����m�sup�]w(� ���`^��FX��ngW+��'�^876���os�9jr��ʺٛe֌��\�б��2^�Ӣ]u��2؁^Y
�юq\jj����k7�w])� ��K����]l��9�����V8^�2��q�! �.W]��o4+{��q�e�_�-|��Z��Dڵ"Y��ֳ��,�@Fؚ)��ۛʁ�Z �9h��Ws�#�oR\:&pC�i]���@��6ѱ�Z�ܒ�N��ՙ�ɜie*�4j�ȺLE�/9�@�tB&�������[��"�"�*��T'lN���P�qN�H鮵*6{t�T:�h-��mI�%bߖ�8�M���C��48��1���ۀ;�_'��;��OkYa(�D���I'5��X	Dv�$���[7{ݯ-���m��v���f�#6[��V����Qy�fH;�e��z7������Ͷ�ۭ��7m��m圽�r���<��m֘Y�v{��:������p�㰑���1��/7^ZR2�0J�!姖gi��p�i��2-�� ����f�����4�.�J����͜Ι��I��q�:�m�ڐ��v�����ʹ�[����m9f��6�{�y�����gA��ɶ�4'���3�ݜo/mb�[[I����)�5������y��m���l�m�og'c�0�������m���[ݘ���<�! �G"�#z�����%�u���FN�.�MliF�0�3��Qm�!}�k���E�5�sh�!�.��g���{^�/��F�j4=�n���ҍF!�"�g{�؆�6"�=���/=��}8���=��!��f����?�=�񼢱��БbI�l]���-�0#PiF�J3���-��z|k�
���DM��s�E4m�1A�b��}��V5Pj4��g�3�+e�/�M����|f�c�����7#=�ځ�Hs�Q��H;��w��fd��Y{R��?{���'U����m���?��������@;��h�ݴƂ2ff{`[-��Ӗ��{�o��q���S[iF�0������6�֟1�	�4����>b+3~��g�>��O9��Y�������8��|_�F&��6d`K�s�-��Ƃ'�H{3=@YpC�D|�Y�}��Ϲ����ׅ�Hs��fbTDϦP�ت�~��i��(�6g���ح�b�Ch�٭�^�gMo{�)�lCb���y�-�mF!���fg��+l��&o�@R��H�G�X0|
���{�z�]�]t�T�$�e�.�ڂ#��2{3=�-����ü�������5��ql~hߺ_eeVoF�ewf�mA\2����O��<�=�V}�w���f�_b����Fov�뮷|�i
B�0��鵹��$�B� 0�=��m�/8��Ni��}��m�ƈ�sy�alPF��C�wtlkm'�6F�5fwV��l��춂Ӎq�l����!�NwwH���Fh��gN��u���y���?�㩺g��A�=zs��]d�Ӻ��2s�4ui�7Y*���l�=�7�+*/�&�1s7��l���F�b9����+bDh�';w�SFƈ���t�j���.�7��[�V�b9��P�m�������#v�2�1m����O��i�6"}��o���]>�}ۺ7d�A�fle����D����)�����o�s�翺}a3Uh�������O�!��>����^��F�F��C����Q��/�����}�2��am�q��!��ew9G��z�i�$5w���䄡'�U��2�+�_��f���5�����s�i�iF�J3ﳝ��+a(�#C�]�)�l[a�/3���_s\.e]*��.4���(�g37t+L�+��z�����)��h68����olD�D$��v��G���]�s^�u;h#"�yw�-��0#Pd�n���Q�LQ�_���؆�F��ޛ�>���X�&�Wm�6+E���z�h��j��7X�H���hJ�@�ڙV�J�GUTm��w����υD�����e�5w��,3D��LB�ȣ����c�n;g�;�[tv˭o=�O�|����9[���ڍ����Eqn���mKn�^ۣ��C]y��\V�ݸ6�3z6]����zw7l�ۗ��rF77F�U7nm�<:��S��p��d���١[�U��i��s��Ֆݱ�ݮ�3c����=�;9��7'�V��D�����77T�h���m�l'Cڮ�k�N�s�O�����Æ���$B���On#ls`RH�-%N"�T�������=�M?�c��<�6r�ܠ��[L#JF����)�����#�춂���7ݽs���!y��˂ ���{~�E=�������>�rMI��l]���[-��J5�w�z����������1�7��SF�Db�#e�/�[JƣJ5Y�O��[f�3�.��=��ˎkM���9�ֶ[An4?s���{b$������b>���g�k5���2&j2s~�E5��b���6�cDh�Z|�d'���Ch��m�̼��sw�>ݽ�t-��#J&�C��Ԋim��6����h,h ��ffP�_N�N��5����F���妾M����p��P��>6�7Y�Q�u0#PiF�Ҍ�{2�LV�������
� �"����LCb���2�F�V��(�iF�}��P�� �'�c�nZ"`�Ew)��Zh�q�Y^�-�Fq8\���L݀I$	�sx�R��H�Q�>>t�b6���_h���4Ƃ2{33`[-�]��9�o&׀ƣ&�2�LCa�(�0�{}��-4F����Ӝ>Қ|۔���{�Pu0�(
�>�S��g/ڡsT��?�vi�L� ݓ�qz�|���9��b�j;�4����[����h����~{�[�}>�m�(����"�X5���{��lCh-�"��@m�lC|��nUx��)wuxQ�|��
I��
&�P�b�߻E����Q�Ҍ�g��b��Dh��*����z�������Sض�F(���;E��`�b33�B�[wy9�75����p�͌>��{���z����o���j@5�ߨ�ݴƂ3��e�[1�2s��E5u�R�7����acan�}�؆�a4{��8CO�}�捍���Pb��iF�C�tlkm*]�o]g^���u�ᑁ�{���Zq�lD��g����!����ot�{h#'=ɫ��tɷ�wP� Ói#���*V՜U�z��kv�L/&ػ���RZ��-��	���Г�*��ƿ&+߯�[-��J5Q��{(��m9���Mh�W_'ڲkW=\
b�����[Jڍ(�iF�=��P�e�O�׊���B��'���
 ��{�U��Q�)�[�H>��_��^�Sɽ�4^|��xHbrT/)b��^u�$5�*$�E�@,��B�.S���gr�|���Y�v�4�@sI�b�د&r�/�('����US%���o<�]��-"7�u�N�����-�%J��woP�|q�*��JB�	7XM�ʷ�sK�y[�B�����n�Q&�����xE>"����Ս��Q��yXA�vخsRB��u?��ZPV��=��-�˲	�T /y�*﮵휉��D8H�P	
�V��,�����7]d�yu�����cp��⊨������Tx{n�dFu�Q�$�_sweҰv�:�R�����*��vnJ����K��X��rj��wn��7VA��멳�a��,���3^*�W�B�'�P|C�n������bs0\���s��>λT	��n�āO:&�B�".��j�V�6����A�x�Nsn������=H���I[4e��#���ͱG �}W-)�Η�f	
b�b�F���:�YY���.�jw#y;�����}:b0��ư'i��x�ըV��i
�����w�;�&�i����g�^��f�0�?�j�7�_� ��wPq]ʵf��b�	Ӳ���c�M����[��]��v�R�<�l�H�N7-!,�����]D�ʨbL�p"�5
8�_�wwuY���N�����j�@@�x��'�Fi�Q��%@P&���공�O#�gX�׾�	'�q݀A����̡����\��9��U~�7��݁�X������$���df���/�z�H|�ݒ�������d�x�
Q^�
���UO���K�'ܫ$O��u� ���Z<��9ꓗU�� �V�m�e�E���vIf�ЭN�ש�|�� I{��`����Q�\��vb�Ҡ�T�w�̄�e�SF-�Εk6��S�|xw2��7r�;:�f�y@%�nsn<�\�4@Uі)Y�׎aÞ{u�=s���{ƴq�7qE٣t�QTա�7������z����]q�8��E���|�j�pn�E�t��2�����9ďv�ևsn�	m�gC=�9�;�=�Ҧ�Y�n:b�ռ�<k��j03���&�g�NGY�W"O=��7m�9<܅���2yF�䛊G�-���8�E��ݰ�ڌ�V��59�`׮6�����nju���vfG��7�j�7/�T�;��}�n "���n�ݒ	9۽b�$���P;یj�z��&�݀H�ݻ�,��ђ,D�2��j�۪�����wE޺�wG��>��|H���H'�Ң�N�uK�[�w���x�Td�z��XI#]�QZ!�"S��={y~$��gؚM��f�����GTq�*����w���b��m+�H$��B� ^�;�[��C+�f����;��&k�@R��H^٬�D_n:�f'���.������$��HQ7���E���cU��V��P��z#��H��U����+�ܘM��^�ൣM�P��3����)Rʄs�|�7vI��T(�I��w`��v���@1���`��wHn�IH2""B13��9��(*�n�Sa�@J�B�ަ":�4I\����Ffj�ʴ�]{�a�"�T�����:J̜�9J�yի�W��w������A'v�P$}��˝Ě��W��,��n�,��d�2
EA�37d.n�}��A ��!oei��C���* ���ݒ�:���
�4k�z�6�b�>\I���|A��v/�ov�[�QK;yya�V���̲"B�2�Rݺ�{{z�m!1�^CǴ���O����b� �v���֛���! ���PH�L�(1I�u��=]d�m]an���Lk�����B�� ��j��$on:�A��ޱ����/=U��z��A�x�����LH(r����v��H�q��� �w?kQ �w���(�YR�w��	�t�4��""d�>����d�s����h�]��C�-Ҩy&Y�u�ż�;X2��Ss��Z��AY���9`�r[�=��st��Ӷqɥ�޵���'J���١u�p'z�ݒI�����ň�;]���_o�;���޺���N����w��IͫQ�C3���y�|;]m�'����0B�@P&�u{��@Wjiw�
��'X'z�?PyU`���b��'6�@�C�\���)1sr\nu{<]so$S�c���(�6���,񧵩�w�잢�7QE%Y������ͧ���A$�ڵ@�ےNFr/���[b���볹{2f�(�(�BѮ�Q�6�r�1��L�I>o{��>'�]Z��˸�ܩ9/�:��M�*"T�,m��H#�]Q$���qq��M��� [��A>:��@ݑ�R�dDL�b���y)v?��J� w��L�y<��uf#pm�+��TR�TUt�p����9�S4�Zr���H���fs\��mr|��̔ho=��!���b�ȧ���	�2���O�X���$�ۻ-8�"d��fn�X�
 �q�*���)	]]]L��-�]�$έP${���i�D�r�9&w=]������ �\���t��nkC[!�FT�'1yw��Q�TTS�]׻�coM �?O%C�fZ&\Z�0|��t+��]6���I�+E%Y�5�kM��ȹɒ#^s���`�N�Z�|M�u
�!q���^p����4		D��*N�TO�}���8i���0����qա@�{�THڶ�"��$Ŏ��ۃ�9�j�N��>$���x���<��Pd����+P����L���*�$_=��H��qOĂ�
%�rU���?���q�۽N9��^��NY�ޭ�R��S�#���bx�����M�Z�Z�ԾeU�R� �S8b�HT�F��|��1�=��������`��N|L���YS5�j7����S��8osey�Y(5���w]��a��w]cVm�����iek�\@�w� `�dj�ݚxuZc$Qq�Q�unl-p5��emq��|�Tb���|�N�v�g0ѾZ ]HtYޮ��Uq�iRڼ̭�wGb����K%E�&s���+�oo[�+u�i�k��Kv�oJ��B�v��Vn�����&��S�Vv[2�o�M��&'Q�Qj�i�+B6�&�L3��A�f�Lk�M��cU3d��nÄBWyH����o*52suu#e+�O���R�X�Ѯ�*������$�;�jq<��^G3�1A��h�;Fm�&��lkk+IV�AnhX��oD������ ��#蛇�[�3WBذ�LGݐ-�C�.����М��8��74h��c�X����Z:t����T�e��I���[2huT��$;�%7���cf\\��&��2VZ�c1D�Ȟ�̥��Q+X��M�Z����e��Ģ��]Ǉ�U9�豠�mrx5fَ�7Y�r��=�:��d�ʓ��n��t!b �vB�cIY¤�j�'A�4 ���2����Ms�|��.�/%��m������'�z�����A-ȯ(���Va(������kc]\l(z��KW%�S���hؾ����N�C+S޲�q������gF���y��^��f�i�6��[[b�m�#\�[��{z61��l�7&���Y�8m�=��z���ǽ佷(��y���-hٶ�P�k47�M�G���u�m��h�Z�����H͎��y�{7mn֤�mCn��Y�痻ls�[��'+8��7kt�imn�O<��mkbՆgy�������X����mb'��7��m�FKd�[[lجsk8M#^ם�kf�f���[hf������0�����^Y�Lٴ�K��k1�����K5�Ӓm�v�:��b�`��CY�����ݎp�7 cm���m혷$m�Y�fE�9m��G'N�'�od�(��qk�/M��˓l�������eX����{v�������{s��͹��a���a������<����mch>|�M���d�	�b4����ܰcs�k˼ɼN�W.��ݳ���dG8�u�8t[;u� Hv�;4��ۣ�&�fd6B�a#�b���u��n�	р��2֍���\�ێy��Fܫۇtm66�-�ۆ�K�炷l�d��8�=+�wb��h�^2�Y�n�/�Λ�F8یԀ콓�����tB�н���K��m���5���n�uv�r�����Y��W�����k7I�6N&�¼n2qs�����fn��[m$rY���c	��<c��v6/>n�v<�L���l��n]�k�)�%cC�㞴�UȄ�ۈC�Ov���Y����㱓/S��˺C��]�qnt�k�mg�x��b���j�h➹{u��\�y��;7W<���٥�Y�v�k10&�9��:����@�� v��T�%��s�wEA*
#;l���ωu�&����Dn�zW���{mc�\�e�eN����e��κ�����5fѭ%��mó�C�y��IZᗧ��nv޸����U���L��i۰�n^<p�܂���>��hո���@�k&ݺ�qj�� ��I�9����srmخ��e�h�u�V^�]h�Y�ӕ���j��S��N̺��;
�S��"Z�������C�g��pdӌ�cφ�-�q�@�X�nMn3��e&w
�듶ˎ��1ɶ�օ1��0X���;��+mlpE��vȱ��v7n�H88c��n��Z���mu�Q���ƺ�vøQ����e8ꮣ���.n��u�,�	��ջg�S�k��6���ǂ�'<t퍶1B>�Ha�uo=���ì�'��� @��7K�Q^.�]�5�x�|�6R�c�s��Z�6�ڲC�FC�ܝ��;
��5�6�;�p��-��n��[B���t��]��m.�nN�qܙŋ[4��9�]]xQNreR��ZxE;tU���%S��g�N�����xֻ��h6w#����Rܷ/I�c��n�d�M\K��5Л�y�ݓH�{lv��Ʈ�����+�L`�n�%��6���g����g������d�֌v��GG�3��0�[��9 	S�V�(N�,T5n}�f��a��$<��������ݶ���gk���=�͇�ۙs���ո�Pm�%���$�a�vU۵؊�%���A����ݵt���+h�98ý�e��]ٸ7]�۷%�LPkl=Un��݌Ya�cs�PՊ4Yl⪨o�?"EJ������mf�H8������E��eݜ�ك,�4�*$�3���&E�8A
L@���ؿmC��f�&�>8�@�{�۰H�O��]��$�L��$؂R*�Yy�-6��s���۠���/�P���9�ʁ��߬�幓4O��P�* ��ɬ�q��qn��$���n�	>V��I+�r�/�����"��$�X=����9��n��TS����].�$o�����yN\�ӶI&��!JFmӌ=l���0i9�z���0�Z��L�=��OT̷���dDL�bg�9�UI�o�Y%�@��\�eQ���ۻU�|E�>�����H�J1I3�\���mTΨ�s�m�n��Y�o��u�*��>L,L�xKW'`�.����H/li��bb���V�)�͸R脣����#f)�ݷ�r�Z�d�A#s^ݒO��hW���{�d����^CN�
��i�{VH#9]
$=ۃ(�3����f���|���m>z�ZS=�&���DB�_*�/Y��S�Ҽ��Y�� �槊�����yFc��B���1���O��P�*"{1y��`Õ�+�A�)`�HW��~$���o�� l�Ƙ�����￱?;!.��{-���gs��p�M�q�:6�zڴ��Z����y>ºTհ������X$sV��{�TrL�ɧ8�r�,j�x��P���&}A�e �w�gQڃ�w?���<@O����՚.����zx6�*R���߈��B����B� ��t�l�!q>7y��9N��icy���$.q���rX����P�u�2�!d���0��4���ݴ��;@�ݫ��^�.�@�ΪH�� �@(��{�qO�&�)�{7��C��^^�*w��P����1w��H@�{ˤ��vI�vZGDJ�S��M���|�� �=���w��H;�ʁ'39Q$�����Q�UL�n�OQbc��)L<3����������I5���H�թ�%�!}��#I����Az�
��j�I>'y����aŨ����Ky�@��`��)I!)�L]��s�����ڜ�B��t�$��Q ��ذ@3�M,�0*�R`�X�dDJPϟ]�>�on���)6+jO.�}��TA;��_H�sb&B���33w�GV=�D�O_��:�so�|su�Y ����~�5#���;�i�+�+h��:͋bS���P�VU����>��{v�B�#�Vh��K��%^q�*e���s���gs��9�tv�R˜��Y�T�xJ ��L �5�]��I#9]U�OL��
�`:�-�U@Nv��X �_\��s{��]J��bg�i�O���l���i�=aB�كnx�T�( ��'$��*�н�$�)�R��	
�OhQ>/�v�A}V��zJ�Q#y��}�wo�]�Ɉ�}*eD�U�'�U�[}��pT�M$�$�^n��$���
���E��L�Z		�HE)$%0���{�� �9��I'nb�aNE_W��{�,}V�����&g��2��1��d��Q���s˛ | ���@ �<��h^L '=��5�rb$UYH9&bk��.�l�!|Nu��Xyy�(T��P|�<���D)?���;�����y�0�!��=�4[��8�+E]F�u�5v���d�8��ػ���J5�3�Cw&�>�Q-�鉋�)+��U��J����G��=�t5]v0��f�O/8�F:�c=���������m�2cv���Z5��	�]�SqBB0�W@H�+Wu���&�����<�vۭx%�Qp���z��v�[�純�|tp�4���ͼG.`�J��H�Γ�4�˽/m���k�ĖHݖy�mPs�u�Ue�k���]��)��4Za�����]�������k���tp�S=�k�9	u�ó�dtq����uTN��>f��X�$gUТI��T\g!��OL�Y�����k.����6IetE�1e絠O���q[-Wov��b��ڵ@� �y ��4�&�����z��?d�}*eD�T�y^�%�j�	8�Qm�1�7g:�X#Z�I�Ϊ$.xv�]��I+fc׽���wʚ'��/1{�T@$��ڠO�=Ϸ*�\y��u�ק��s���m'��jQ��'��{2�|{:<Q�5�ۻpH=��A!�mQ�Δ!�{OX��&&}>(Siݧgۡ��m�����S�-plqpֳ*�V�<"e�D����;-�Kyʉ�>�����^�}d*<�b� �ӨA�8IA����v,�J놤�f�࣮�3 "�|~�㫦9��_�c˧�+.ic ����y�rt�΢�/�v�P=��t[��R���W#��!�E���$c͡D���݂lw!InR�q��{U4�i>V�̌�2����o�P$��u~$���7&�x�{1����>wd�2TJ�Q>�9�i�ݼ����D�H7ݮ��H-u��eE\ω�5�@�+���$�(��5�n���9;�K�����Y��H$��t,x�Z�TcU�����?u����h�����;�����{Lo=v�&#W�kV��l產"	Z�O�y�q �ά�K]j��+(L���d_>��A-�m�>�n�eB�37~#��Pp6���K�~$Of�X�C��^$�Y���e���3B'�A�����œ잺|IS�2�nj�tȞ��o��nX���vg�LH���T9=HV���x3q��H��F�SN�2\9�\ۮ��ܫ�6����]���6�`��=hPW�3 �S1(̈H]�m�R�뵕�4��b��FK�@��峘1��]&����q�b��*aD�(*!_eQ$��km�:n�=$)ݻ�H#'mP'��s:�ŕg&i�J�3�?�;�w���M�&�V�cnG�	Ȋ�IՋ�^���Ual���~��R������sʿGK��	�u�� �\������\rk~����r�'�ٵ(��W[��ӹ�~$���!�U�߬�s������	;���#.�9w7������-DJD̨Pff��M� �޾��>���r#�Z��.� �m��(?v��*僈Y�a��-|��Ӌ^ԈU@G�T$_k�|I\�f�;�E7Kb{�T�s�V��c�ldL���{;y��i[M)�8c�yiv�ź����C��
SjB�z?e(�����-��SmQ>]�3�PfQ����z�H[�lZr�D�ɘu�P"�_U�H$�o�\Cڽ׵�$��h�^�e	;k������r�uhp۩�Xu��nt;����S/I��$�� ���(Q����.o�˛-��hW��{W�Mw7=v(�![3�{�ō5��Z9��`�B򮨂I�Ϯ�I �o�X �������*qM���)�D!(�&}^|�.�$�o�X,utl�4�V��O�5��$�W7�,􎌵))B�37`�o�Gr�6nJ�	��|�� ��_6 o�4�EB�zZ�+�7́W,e�1�c�Fht�şFOZ�y�>�A�f"A.�e�$x����Z�_��l���e�cN�G�H�2�Th�Ϲ#{u��εג��Aa�}5����ۖ�-�ZR����"��ŕ����8�^ܛ�ֹ�0�n�4�yyrd�3n���C�<Im��Luغ��8��K��`���]d9���K#�]�cxm�=�n-es�=[X�v��z�PQ0�!KZ	���y��Uɤ���cuDf�WOR��ge[����;J���7a�i�^�r���e�%��3�����n�G�R ��yg\pb��I7q,˷vֲ�\�V��8���bM���]soD-�m���0hyG^K]s��������3���:��`����P9�#%�nh+����H[ϯ�ٶaA�>Azo�]��u���u�U��	��	�s֨�DY�=Q�2%�[�6��;!"D��D�ߋ�y~�	#��W��wrg M^�I� �����\��$�݅h�%j�>�f�ws$�v�uȯU��d�KN��}}��v�b�=59��/��X�W�㤱�ic�c�/m�A�h���r�Wy��G.�7s�m��j�i�I4f��%T/�ޚ�Ǉ{��@㔭��㉚zyC��;c�ʦ���38�h�x���Y�&������w��ut�����MQ$�;y�M�k�}�Eݴv�m�A$��tI�L��Vw����ӽ�L�v/773e6�����],8F{fYw��/�Uc�Kiʽ��<�v��v�*Ƽ��|èpun�yhûYM�ob����F�Yfo��'�H�ѧD�$��ޒ >Fo_'̙OU�KBT�dX���o�n�)�m�D�{}�lB@��^[��g͢I&���$�7��}
>�>��$n;l�����7Vf�]���7��&�$�{��$�Mj���^�^��ϻ[��=�ˀ��r´T�9����쐚$�,��6{�n�z.�#�6,=�eπ@����{� ���f}��k��wG�,㏟r���-t��c1#Ʃ����ë�ۅ�Q��YJ6�EUS�\�=]�r��$��3���{�f�� l��vf|�Yw�fy�x}�p7�щU�V�� �X@����<f�Ѿj�=��dK~DI��zID��O����� �LE����y7�J����JX��;�ﳻ ow�X�
�gj'Y\��8Mh��R��+{3A�\�ꄣ�V���-�dw�!�%��y'���0�s��w]hʝ�D4gͥ7�����.��v�[ź]IIF���KۘI���L���힝{���RX&X��+$]X�W���*��K-��o�6R'g^��4�ܑ�јt[x7�L�*�Mq�ǝ�Fx���޾�.�;�`���n�`��IR�sЉ;I���t�V���z��e���)�Sou������(o+�O���	wR�,��I���3��UFl�-��kJXq��Y[6�+[�]���-:ΨhZ�3��S����;��2u֢��5vV�ƀ7B��l��+-���òu��,Ӹ��|F��k��yi{����[{Ա��(m�z�eX�k{�2ѯ�����L�*v���H�tn���a�W97��VP�/.���:��\�5Cn��v�-���wrش�۫���p�זn&$�����{��q6�����Wa�8~��w�KKn���;kl�
��p�Z���[���c�u�%����[b�l���<��Q*k2����`������L�[B�Ɉq0��P�,6�ŨV�ӭ�����'S���u;=]C���QN'�9�V�F��	�л��೛�v��t�+^]Aݎ��S�'��Ǉ��7���p#�%H���J�O�3�6K�7�üa�v^Zzg�:0_
���=�h�������j#K*%c��,�N�W�D�0:�G'y�3�)�t���
X��m��8]]F�0u�P�i�o����ɷ�Y�~��r�۽�=�R͵�{�^6e��+8๵����:�{oi%����m"ɵ��y��ұm�;F�6��#��v�pm�d�nf۱��oL�"q8y��s�e��e3M�ˊ��n��k�a��o^����"��׷��G�[ef�fI��4�Z�8;2��i��贰�#I������yi8�;��^�;ۭz��k�a�k"6���!/&3��v͖�[k�;ͱkC,��ͬ2�������4��7�w�kM6ݛ5�%�[��5�)�����/fm݉�h�$����3Q�f�v�ݳm.r�޵��3�:\[NM�[X��v�+/<�3�n�9�nЭ�5�Ԝ�Ƕ֋mŻv۷'E{{֢�(��ɲ�;9�X�Xv76'3Iق15�glmm���[I�,�L'-�u��jHtN۬S-yڼa��i��m������ }����Hg}����E���&�����xB�񽵀o����*D�'{�:$�&��G��z��#jU~/϶Htw��U�V¶]7���.	 z���J�c���n(��L��$$����6Κ�����"�Ow~g�m��4[L�C��E��9,g�����3��B'3�s��L��3;y�
�BH�2���y��$���?I<W��M
�^�t��<�c|g}٘{Jv]+��BI��湪 �	��h�{���3�q.oЀ�/}��$�\W��H���м�η�1�SYKu���\�0�{5�޽�DJ��X/��I�9D�h��u�e�t׷�>kw�c�����;�
�i5Hgd�MQ:}�f�?k�lx�$�'w����Vu�(>�z������	�YL�$�.�)��+N���=�:sV�]�ܥ��Jt��	2���p�ũo_f��T�Yl��{�E=�
����U��.�4�w��o# K�걺(okh�$��9P׻��f�@?_�[d�$�
�x�$�2wzO��=Z�����ؽE�Fݍ���%��ߥ���sz��Ƭq�M���#��URn��������M�y^
t��t���h��>bt�$�&N�I	����y,��-�w��t�5D�WG����+R������y϶εt����b�wd�f��z,d��O�N�I_B	,���z�)i^�j�����	-$�Lx.�|������7�� �׷���ٽ���{�D�&�~I�I$7�w�ǵ��\-��ڮ��. �^�maq۵���j~Z�����%h����u�O�.�� AgkN�4�z��.�K,DFgƳ�������J��J;βf�&���f� �9�o{$���u�gwǷ��d(�z^틱Q���%Ў�a�L��X��V�ٷSj;���G����?,X�Ȃ��u7ڻ�l�ẕj��>c�	Wd��ۇ���x�k��v�s������sn�Pp�b��s�6�(8���5�f��7�8�'x�;mrs�����=jػ&�(2,Vu���녙K��͞q�<�;�� uۖ}�&��6pR�3�{T�.����m����#]4�SR�>���j�x��Ӟ�v^����ƸP��m'�fc������ٮ=��c�ҵ7%j��:�cMܱ���<s`����������%�"\]~����y̒�$���k3��� ��f�  ��$Ӵ��K���uՁLGs﷏d�'IDH����$=��o�w��K�ˋ�����;��` t�lظ0"[x�(Et�����'���iZ���E�����6 9���������Vw,p�=�u��k}ك �"���>����2�+%��I��g7���mӗ�~�*;�I1t�B~$�r��ۢI$j~jJ���2�4fw�HWV��jn���������moY�e2r�L��ݳWL���~$�h���� �CS�N�'�.��}C�۞p�b���m'WV�]����.^�Ƿ����w��ʋk/��B.��X��y�w����7���+�@�|�{5�%ؐ5���yzú;'I!��u�Mo(I%�I�W19�f`|��$ nB�SQ��`nB�IY����a��}���W4i�ӷcc�!*��Y��Md������k,>[�����2irb�oun}��������٘�6hj~i�'�m
l)\3�E~�v��P���N���7l+e�_Og1\��f�ɢ@J��[�z7塚{�L��_UX���B"P��x̊7����9w�_�u|Hwc��I �5>i�&�?�ޛ��/U�I.޻2~�?I��Y,$�Lx���{�{��;�W��]/����'�~��$�hD���&{��C2Nu6����]C��:���h��Cn���h�s��nK8�[��w]���}�Z�����n�0���&��&��TI�����k�yWt��k��g����eĀ���E������}ޓ�@��=�=�,�S�f� <tI$ѝ��*�����Ѽ7΃/:���>,1bbfeH�� ��w��D�{��s�Mh�����k�)N����CTr��*�f��G/"6#���)��3�F�U3p�:2����k��K�l�=�)E����	�h��E�ܜr:3�yz �=x�	���`�x�T�$��X�s���ͽ���"��I�X�&��M|I�{��BI'⯽��v}�����If&��x�na���cώ�9��`�A���/�,��������;�J9<�h�G����� �N��0�Ww6��B���������۵�>'�&��g�^#���Mt��ݶ�ٔ��?I��(I$�o�7�{@ o����MI*��l�hv�%��9y` ������ՙijn�ԭ���g���Gfq9mNw;���Xh�o{�	ȈS��D�Lu�@-����r��w���`Yb"4���?z=��W k[�9��\�/R w��������vf��曄�X��Ut����髰U���I>m�bQ'�$��u�D�$�)��eĝ���|Xw��uj���M�����K�#a��l-�����Z�2��˫�.����`�������S�inj�������C�����Y8{�Q|�'.`t�rk(�O�`��wq@:g��|I��U�u�&�O� {�=EC����N��H�D���[!]�[�F3��{y#v+��x��\��Z$V;,�s��l#R��~r.�#�ɲ}	�I(��3D�$��ۦ�����h���!�O�_{��&��z���G/	���a�xM��W�N�s��sk`�-Nw�3�@l�{. D�M�kaɺ}��"t�*I	�����y� >�g��h> =s����GN�`�g��$��wZ �)����je��k���~�OS��۾�m�;�˂���sU�#|���iS#�>�A[z����9m��6��	$�I>��#7�;�{ٿ�}f�}}m� }�D�N����7��^�����p���ﭚ���w�T$4����N��h�]VH뻬
럻(�s�0��ݛ�v-OZ^_�}t�9����6�"ȆJ6�#���nF�'rH��	�z���q�lv��r����cn
;ah2g�N�9y�Y�6���7�뭠1����k�G)>�ݟR�=k�n�'mk��v��tE-��۫cIֲ�`�ezϒ�Νt����˯Y-V]k�tZ�6�g4�RE��f�wj�qn��5um��N�&��`'�g��[�瞎:'��wU�NT�hI�ӳ�V���X��8�k��j͜ݼl�P�s��v��.z�=+�]����~�d�]�B񽝻�� z�j�������kͿ7���9�{L�C����={b�^Qy�^��O)�5M{�J������>��� TqWl~V�[��챷o9xBLx/o���  �{�f���o\�y띞�s�$&>hI�7��`�j�5jV�j�0�{�����%���� ���X������� ��zBl�[�ݕ	���49ti�%{U�b��,���w�okcg����W6Ofn�x]��� �q&�4w����$�}�L���{_q����8�Ec���v}].�n�Df�k9޲oX��n.���N �Ʊ}�߾���b�}Uב���b� ����  ���n��BO*ˠ���5j��$�G�����S�z�(�v�����ɬ�.��sJc�{���p|���s�m����9�����ts$�����7/t��O��s��_�-iݹ�]�RɗI�C��Nc���H��nI4]���̂N�x���䳧`��^رV�+�dY<�2߲	�D\>٢I]ew���N���� ;�|��C=�=�z�`�G/	��v��	����׸|N�{�o` '�٘��k=�ͪ�N��%�}����{�\�7+t/Ĳ��c?Q&��?&�B�1Z���ܗ,�7ټ���D�{�� �t��\�>,koj7�lv5*�����NJ.�y�e�\��Z��4] �cu��Ah�u%�?_y�����#<k;��k`���f�$�O�73%@�wc�G}�d�A$�9���[����X��Us|�3�9eRo�;#�3y��>��I�%wZҽ ��=�݌������d~�QD
7]�2�Ok�� �]I'�8ś6��ӷ��R/�CV�K}dN�xŤ�:E�ۧJ�mW[����WM״�����s�w8؝w�v9�Y��m�9\
kc���g8�^���l5;��7�p׷�>�vr5�jW�ȳb7������p���Dſ?�����&���aپ#�*`PH�L��,�G�2�"�9&<:#��D�&����	�^��r�r��M�נ��f� �������@#~ｽ�n�vrNԼά���R|}"R2d����L��;XӶt�d	 *�bmx���g����Ͽ��NV�s^3��p������3��7	�;��B�>�s��o��ۛ/ƹ���k~�&�h��j"3�ތBT�]�t����%E+�O��$�h��zHA'*��2ׯ�z��s'~��x޸�!%��b1���� �}���Þ��W8s���$l�7����}�����"�n�H��Px�l�l���;י��I%8�" ��{�	%^���C���ߛ�'m"��lu�Au=�tegM6�!`k3���X��nE_(��9����w7'ݼ<��2�=�YGS�W =ǵ������r��~dx�}��sa����X�ym��&���m�$��sx��}���@��f/��s�)���F��cu3�^6����or݄f����/%�2é�UT���'�u�T����u�5�d�w{�r G}֙4g�R����e� 7�����sM���I��%�K/��wn^�um��|&��I%�{��{oi ���vb��-�{�����k��5	����Z�c��}�[ h�;��{�y<҂�əٚH�{�$ �&���u�dɴ�ѳf�Y����7�u��^ܗ���L���`���;����ǯoU�Y��Wki��g9��`�>{��E]�R�|>Z�$��,^��{�x�l��ql�����J��+��i�@�$����%���%�P$�	(�$ IB��$ I�	!K�@�$���B��@�$����%��I^@�$���%b��%� I_���%� I_���%� I_�	!J�$�	/�b��L��̋���� � ����{λ �����           @                    ��      @ t   P   ��                          �     i��^�>��k��<��ur{7�Ϊ<�q*��%�ý��c��s�ܭ�� �zzn�7��{��z�  o� �y=z�������U/{��w�s���m�x�ę��g���q��ޅz��4�  � �  @  �U/#�{��֫��!n��^� ��l���Z�>Ǿ����8>�����������W�  �  �^�t>�sm�׀�������=��Fݹ�W��<���������z۹튥x  � x      {�Ej�wϸz}�_��_x{��k���l�۽2]��\{�{nm[׀�miamn��x  >  �{�ݛ|�;m�� =�˻������n��_G�Sͽx��5��h�u�u��6�w�/�    >      =�m۟Z��wZ���zk۞�sLn ��۷=P�5u�ʶ���y+� =�4����v��^  � {��ˏ�T+;��h�n�,�[�j����;� ^w�^  �{ t{c��@����}� �    �      ��vOE��
=��{}ǐ�S� ��ǻ{o��^������/;���x����:w��� � ���9_6�49� ����{��ͫ��%��ii� wx�כ�8���+ֹ���    ��T�D#F�S��ѠhO���SM= L#&4��TR�@       D�*� �P      ���h�R��` 	�	�4�M$@�IOA24='�ѐ������?u�ߡ �5���?�;����$$!a��a0�p��!�?�Id&�  ��H�HB�7�G������:B+&����8D	!C��d?�0��!��.��������?��}�!2u��oR���(���������y��Q��l�"/��o�f��vO�Η$�e���ٷ���t�xh�i*�+����zh$�k��u��k��v�.y� ����7:�8���o5�Z��L@�[cC�)a|�K��m��fL����*f�.CFe];��nCA�.��D&�;�C�.���xKqMٚ��.�x>��U��Ovl՝;b>�]\Sۮv��1�1Hx�3�yՕ֎�-S���q��wn�i�ٽK�Ž�e{����[cmѸ�i!Ү�`�sD�:�t�3��3xCtM�U�;&�0Y-�2���cױգ�i�;��V�tb��Չ]�����v��ء@�K�.��������q�piZ���a�9؈Ssx���"1�]mn�ގ��$��g뻯�v�O2��t����w�;Gzܥ�����L`����wg`.ܚ����N�@�χõ�GA`�n�͵���4�F�\9v�K�Aܲ^TKo=6��x૷W7�L9�s��HЭdڢ���ɀ�y��*'�r�S��%� �=K�����UY��WL���!�=-��	�,�q)�n�$\��H�?Kzp�<��⮍�e���_ou�&�3fRq��g4�K����nin<�#�{i�,�1Bt�0G�$ޜ�|1,�L��+����[�5����r��6I��z���!�R��;���c��e�0^�VnZ�uέ�7{��f��|Z�P�m�g���Ϲ>��l1>7�bp����s��l�FZWۃWe��WN�&ݍ#{X��kwv`m)#'��o����V6�@|���n���ڋ�;�u����K���lv%G<on����y�.��8��0n7�otݣ&t"�%���D�&�%h��i�H�}L��)�V	S[$-�K-��q�h�q�:��9hxI�p���|�F�/��_1��zc�,u�gd�
:X��
�����6���]�]��;�h�n�ZBEw��]v��͢��������U��w��7�<o�3��U��睹�.ZaE�A��,\��p6u�J��,���6���i���� ��ńv�$�
��L���Ӆ<�0L.l����la=.^��nX�Ӽ�]���yM��{�ݝ�ɒD��kՎ��gf���rjP�]�|j+�����h��*������ɉ���7W=��k�m�7�n��x�ʜ�L�*�d��
%��bɝ�s��v賷�,��iqW,*�0�k�/	�`�rȲ���ե�#�e��BbG��Ӡ^�&S��%����l�Wp�1��,ӭ����N�p�u�F�rqy�a+s�`��0���5�-��x����v$Fn�-��k� �?�FQ�L]�c$k�Ө��X89\}��/Zu��iVN�yCǳ�-�~<ܗ����:]�x�c$�ېut��mt7P9xw<���vp��7�'ֳ!ͭf�w�b۱0�ϰv^3���K%��z{e��渭���=6ٽ�!)�C%kOzY�g]�r��qDS�%Jnojh}ٴ7�L�54��^�{u<��Y-��urU���g^M�	px��id@�jҤ�r8V$�[$���x%���ww�[�����Ʌ�f��i�HI�@���>SF��9��q�	U4L�4��G�6����s�ww]�!�dT���(��PŋqAq�!���CT�l&,	˯r<K6ˆ�F�-x�:N�T��䷜(a���{1N��5�{��.�>X>睩" �,��PF��\�V��sWC��9\�i$����8� XP�(L�J��8�'\�W 78�jỌ�i11�'>�f�_oE�P���@"��m���fA��d�w)�V �2�v�M�kW��N|�]um珊� q<$+
vVF t���&��Y�u8�)�|p��S�NȦ�iaTOgr�9a͛�պ~�9�u��m�UCpo-��i�ڙ��)�w�.m���4�g+�&��ȼw�$�����z'C�	�c�{wL�;��s�ٳ9�Ѽ�q%��Nݺ��b�c��6��V��ۨ����HzV�Z�+�i�,%pu�5c%
������s���r��+�O`�]Rs�&B�h�JN��m�:�ѣ��������v������H�挤gS�o��WX,�6��ө�74�(�6H=ĹB��+HDq���96e��{�I=y�T��+O�wGr��(2�"=�'t���6n.�����\�����2�4��{L�3���W���w�p�f���ĭ�)�KC���t��n8����|@�Z�K����;�^�a�nM\9�ȹv^��NN���H�;�w�i�����Q���YD�.�N��h���!����7h]a�ר�)��{����Ui�.�w�P�Ds���Xv�A�z�����g`���' ��P��@�M��ʞ��W�fvv�<���I޳{�z����p��[�'ꂯ�a��{{�cW#��ŭ����3�{F���*��o}�^������������( 0\^hj���3�'��̵8n^ӡgp�B��������T��7�,콌oq9��\�:�NA~4��m���t�34�m,1��]��^�m}q"m�3�A����١:7^���;�,v��"�r*�Mx�-��ʭӎX�'A�^��!�̟>D+��vb�F�GeG
OV�eٜ^5ۮ$��9�v杰��#.UvW�hї{���d�3�ܰcD��sgl���È���+��mz�hh��VmjNé-�Oh�O9a�,�� �	�N�YE%n[�����3�� �L՚�hl����w��{e!��ނ9r�Ő�&Sp���.V��2'kL���;�!{%��ǗsHZ�J��y��N靸�(����Z�ѽ�]�\��HΖ�XԴJ��kZ'yh�y��j����KF�;b���3�՜�avE�V�3Ѽĩ8��݋5 ��p,��<�A�5K�7��n�̼Y���gd�Nл7� ���ɖ;	��-��*��Ц�9n@~��[}�rO��9Ϳ�Z�� y�A�f,8�$�n5��!�It tJڽw��.��ǚ4.]e�Z�M��r<��<����NZ����P�2�Mk����ɬ��Ցe{s��ssB�N���T�Ȓ,��� `,en�S���6�#dG9�&�у�[�6��!<o�]X�H�*��y��ǹ �@	-qMX �.���Y�{FE���6���44w���8A�����N̙JT^�mG��z`Z�ћ��ѬXq�j:�4s��"�W��X�E��A�1sĮ���8��·'K�qTQ���ؐٶ���ˉ�` �N�j=�X��4�C�7�nٚ�9�� �@�&��X�N�n�����RD�J�]�I9-J����F���SB=�j4t݉���G*s�����P-��V�n���7@)�����>�iS��A�����u��xF�v��:�su��PD],�AFة�6nR��(�j,e��y�6���(;s�K�6Ŗ��ojsGq�9�SΫz^�c7U�S���uZ�M�����d秸��w���٦�F�v�3�W�u��X�`����7�h�r��8˱��]�ǣy�NΒ�w8�PY�vEy%�b���~f��wtd��;T
��L�w�H;;y=�������ۨ5� W��2s r�n]Օe�m˱
�hs�i�j<#�;9�@���F�Vg��7*���Xޮб��&��;q�^�z�ћ6��r�>Y���[�o^�Xy��:@�G�oH.m5v)fB0��
��Q��B���l�Ը�O�w7/}~C�W�B���O�u+o=O����X/b�DS�?�bp�9A��K>��ch��Yj�:aɁ.⎴zX7V5owM�����.ٶ��8�����# Q�t뮞WB���%㚟lɋe����[9��M�w`�'A:J2�(��ls�X��`���6@axE����K��艜85����
��$�8=���/��h�nǼ��8Ѫ;fǴ8�\9�[�$� �Ц8����GM��Yr`죶�s�$���k�y���ν����sT�/��t�׸C'�9	G�t9nn<���d
��u��^7��7 �{�`�xa�v�&i��s%.�8�۽�wN���h/v��Ӂ��8)��/Ru+4}�Z�-����VD��B؞�Q���'�d���&�Vq��U�`��G�E��#�nN�g�8�[
'�ܿ�]�n�e�2��_&���M�E�;��SwF�P|�o�,���f�Q�;�cGd��3B��y�����\�vĸ���''��\��j5!�K��-Uo`9vn�@[�r5>3[��xo?�W��Q�­�[�x$w<�� z$�K9|����]��,ќ��J`������7���[�=��R�>��X.*1n����l3���3������Y���� ���/Nׯ%�J�˦���8hu\�ݺS�C����<k��n,,ӑ�nL��ڂ�ON��i�H��XYc.<�}8��6v, ]�/t�H�]��;��9�ʶ�,�.�(aA�r#�su����}�^Ţ�n�X��C.Èa�"�;LY&����-�c�&4j��?��_
�D��1����x��l��˨f�B{ʨ�'I��������,����]'�~O^է���0���	?4�B �XR@!�J�$$��E T"�HT) V� "� �((�P� ��d�IY	� P�
YA`E B)$��Ad	`E�I �H)	
�"��$P @�@P��*I	U�$�$�J��RH(� �@�Y	"� Y�d,��`E II	� �HB�$%B�$�� + , ������������^��B���g{  ��:�! ��������!����������/���9%��Wu{��@w����K=�I��_/Y�"��ס晤	�^��b�o�t�J��f�4^���x[�I�ӊ�F��O�+�3�cr��?D;<��6�L��mѹt�[B �l�׊nsC6�\x��
f̓�<�e��#���/���Zؾ�����t��^��}����X�����|f�����w�u�����"p�������+���y%�sۦ��E޸Vq��w����{}��<�@��ŷ_���W���t?c!ݏJ�7	�ޞ����\�&�\���7\���s�Ӧ�l��:<�����c��X��-�ɞp�k����=�:aw�KV��/"��*[�s�'G-,{'�Z`�P���|���{���lP��{����F���"/w�><���"�{�yz�E�L�p�}�H����!\�x��]^�'�%kcOt~�h�M�ֈ�{�w��N]-z��M����{9-��%��= \V�D`cf��$�?W�yG�;O�e!�����W��^�6]����Ɏ��enx}o ���:��xoz�q���'U�뽭v-��-~�;�+��s�r��d�WZ 	k�|��X(l��;0ܻ�p�xK��{fqc��ΟqJg&�Z�BĢ{˳=ں\�lҽ�}��F�ϱ��P�>�>�R�;����0}�o{�V.��ۻ���B�Q�xꤗ�c��>�8x	��0ԟ�e��^�r,���	Ǿ9���z������y�FE��=�SJRз�Y���{_�-�ڛ��'�����D�o���B~�Ƞ5:J���@���Μ<xÄ�=罖6t�]>������sW��W�U�V.9�m^��P˝T���]z��#l𻼽�=��ws�{�'��s�UL,�.y�\�h1w{���x<5G�TyN׳7}���@;�RZoa�i�x��g�Q:5jX���z�|���� B|���y��u��\&
�o����
؎5���ԲP~�����c�x���[�M� �>;���m�lVy��O
4�^��z����^��N�8�ۜ�2�>��E1�=��Q�(
�p{R옞[lw���FFx��������^8yc�X笫"�W��x�Ьx�z��~�{��|� �0��;$B.�;F������TB���D�꺼�="�r!7T���9�/���O��ڮ�{%�]���5�'�@��������s!*�=������f.�,;#=�w5|xA������ǽ�����S='`K�ǽ_w���G<|7� +|������.������M�W��-ͬ;�mˇ#Bǝ��k�4�OP�M���	�|�� +��l���v���W� l[�uT�F��G���g�M�[�\ص�=ќcm��[��iӾS@�x	�8���3���r�~3�"l�ƞ���þ�q��}���D���I/�������BH����ۙ�s�3�T�Rťk�ՠ�\�Ć)t��gҽ\��k{���AX�{�Lq����;�p�ڐ�_��Bz�C1�������}4С��^�}�pLV��[S��$�.�{\�"/�C����B��R|F�FpcTy쪋�ٴ��2歙a��	�;H��Xq�Wyܹv�U�����ڍ&�0O\wE�/�K�{7;G��&n��{���Y���x��أ�;]}�h�uw �` �����s��/f���eB��=�3x��W�vi���Yž2t�|^�7���i��xo�3<#�%�g��y��i*��`C�G��~��RJ��9k^`�_0�d:�i���?z_V=8<p����u��k:d�����ǣ�`2ļ��.��f����+#��5>^7�o������w�����پ�+�53q������ɱ������*�K�s��>w����@S<�߆��0����_Kp���}=������d*����ox	~MR�4Ӳ����5�n�(�:��=^�2�LO[�q��ǩ���{.��9S����r�z,���Z��glǋxy�E];դ:��=����S�$��-�S+��-s{=	d��=��Y����u�7Ӻ��W)e~�O��\���L���6���CWw�� r|=���i'R�H��{���S��t5q�G|d龾�r���<;F{��N��N�>��=���ň�������t��Uf�u?Hߖ��C���d~����p�����/=d�@zA78��������3s�^쫼�vx�/�=�@ex�c���oRkx�u@G�2��y���[�U��:DO�yX�üNkܣ�)\�D�.�A�=���z�\�vm,y>{�/�>�wÍ޺��,�|'����M��])�܅�M>[V�û=�y7,L�dL!�T����+f�W59<����b;�WB�����Z�-H�{�'㚖zjƺ�g�$�>�C�=���z�{t�M���}}B�{A���L�z���W�{���*S��':�,ۻ���{���m�����;�����іW��4���׹d_��$������-�/��|�����Ȏm~���>=M���nu��}��k�k�o�>����ɾ/̽��,�z��M���j:��J���ɲc��=ֹ)����}��{�H�˞(��D�ضn3-���Y�1���;��;\����H 3u��+�ޔ�|2����Ϯq��/���lsW�ח��<�QI�x?KI�z�o�v++�6L�hd����X�u��r��*�G�ڴ�Q�*w�s�5�B���>3��!Ü���#,G��ᎊc>�6�w��'��~�8�C��������j�Υ��.���k���,���N����$��a�wۓ�퓃�s��VNy���-�|�>�Փ�SwD9}q=�#�Ւ���^���`�8��%g�+��'v"�V1���0W=M'wQb�X��/�hy�4��=�;�ל�sy��z���oӐ(oI�7CR������	�V�o�=�)��K�"d���bǾn��=�����ѨN���ug�a�]=��i���Ώ*=��0 �[y}�|�(���}�O��2ѭ�=�=훗4:i��V	ڐ�h���w�z���NN��)l�w��<�ל�Ξ�!ᾢ�G�yۺoc>!o����Y�X�{����}V��rA�}��>ٜ{���}\�~��f�n��P�L���E��� �/"��k�\��kR94���s}d�s�I�q<ܛ"�.ѩ������@:������{4rdk�\�rr	��Pd�|_������]D�hK�_�ݜ��Н]π<�ֺZe,�_��~�T�G�vz��@��e�>���W�����4{��ߙ/��޷�H�7lˈ��T��r>K|ʰ��;�J��{ϻ��ڰ9�
�yc�_��8��{+�O�[�f�˲c����˾�Z�nL�u5��a��tn�9����x-���z.��j��{�h��F�g*܁��W��1�{����V�;��{��5��SG�{�W��Y�[W=���C*>jJl�����:V���>��Fg����އ���c/�����O,�{�	�N��S4o<�Ggo����*1`� l9疏]��}۞�#��-�8���]�G:���2k�s���+��)��	�^�y��;��>��M�
rv+�_x��2�
6`�9F�m���zd����{;��r����p˝�m��{W���xI�v<���k��'�I����S��8w_o��HyiB����8����D�$:�vq/�u��=��_R��X�˭�}����A�<�~��si>��VA��4^�&���\5�/���B�;ۜ��/�d%t����i��t_{�s��s6�y�>盜����-�2v���F�i�77�̽X[�����;�l�V_o�2j���pl��^<,����3���w���>�WG���K7#mU%�yuP����Fw�M�=g���x�����ċc��O��[����;�G���oN+�O`�E|�]i��򯻳H��8�q�Եo#�u]=�qUiH�5=�L�����m�0�w���o1C�F:L�3_{| ]�!ؽ��]5ֆ�%<q_J�:lꘉ���^b]�<��o����l�P0��ݞK;�{�����������V;8׏=��y�H�S��<ojɕ��O�^��mL]�s��]�zE��M������
Pwm��85F�5�� �{h�ՓF����&�e�����e}۞����;��W+�S��s���ǁ�n����8zj��y}5y��s�;|�	�h���I������M�;�}}�^ٰLN-�P�M������ݗ��Zqa��<�w�N��m,П��-�pS���s��^t��o����0j��P����J���� ��HL>��`7�>M�O|�=��^�u)���A�c���I�zz�c�:���(cY���Z�C��}���	���4��K�,{��'�͌�|pG��T`��q��/`��X��=�����p�e���ﷄ�=��Ϭ��=���cɾ��S���<&,��e%�?#�,sۋ�҉��绦��i��x����}��˦�z�ӽ��_����K���s}8��U�� �o���i�k���%�3D|�3��M�����O9-9��y3�/��S|��.Ӛ�n�q�c}*�L�:_{y5�����j���OY�iݾ�=����zwyS�j�@�Y�	����eg����
��R�Ё��~:|����OAnY��s�a�\Tv�^�=�]-��W��klʎ�=�z��1y΢�y������OO/v�v;�yּ/�����B! ���||���o��˝�|��=6�N ʊ�uu��={pN+`z�u��k��p�Ӳ���b������\{v�O[�Z�;c�m�n+�k�'�6y5��[WSְ�8�:���'���f������x���Y�m�;��g���]��m� Э�ҍ��f�R�6l��m���n�T�(�qz:*G%��\<@�f뵫3t.N��Ƈ�Tֆ����:�8��xK��|�ëv�=l�[<�9L�;�\��e]��kJ3���O�D�Z�h�;�zݘ썃s���k;���|WU�ŗQ�f����/M���Ɇu�O\�8�w@]��kq���䮞wV�i����3����y*�c�g���C��[���u��i9��>{$��ss�`��.T���v.�-ι�p���U��@���*QF 6�q��5�nl�l�3�����һC�
��n�׸��s�Ÿ
���{+7I�ۃ�ѵ��eQ�'�'���q˭�Gv�.biC�
ؼ�F�l�	{���o\��˪��6�b�/m�t�ӏl��؞���g��S� ��=�ypy�փ�nf�g(��b�=�Y}�����vOl�^t�93�qu��Xɭ�c��k0��������g�l�͛�r���-�m����1�X�=���[��<3����]�����zҷB��t�v��O������ndŮ��[]�b�	�U�Xx7\ػs�K���6Sw�6�s{ΥCQ>L]��&��x�-��Zʮ��'7����9ڶ��G�fN(�5�tvq��#p���6+8�'[�1[b�ɸb�y뎶�).��h.ֱٝ��6�1^yӆC�qs����\n{9y^����z� S�]�`�q��W���
z۴�j|�v��+�5��z;wg�٪8�4V�1�˸.Q�r��ڷ\cJu�3�>�8�F��:�5�u�%�{��n&{.�	8�'����Ӊ9��Z7[�ލ�v6��5TK��9D*�;by��W�0��m��M݀��ۡ�um��ۡ��5����2I`�>8�mˮk���:�E��̕��<4i��������0 �Վ0�oX{�{`����Y�#s]��i4�7S���!��7n�إ����l��; �`�[�r[�����G
�Wn��9y2�ݻNoX�']�.��Cq�s�x8A���ùg۶�]�����4<�bj�t��ǖ�qǶm\q��q���=�������3n����n��Nڤn73�cuj5��M�Zθ�զ��f<܉��O�j�C��N�����n͸Y�r��/=Wu�<j%{k�۴h�s�y�c��A\p4aL�a{N2+k���&�3ۃ�VDn���T�:T�n�y���G^�.�b㲋�q�օ�v��x�i�L.�b̍rl����B�f���h�w"��]\q���p��eM��8�69�r�g��Vx�8ێNE�/�Kq��� �ՓuHً��U��F�h�1���u�0d�;r\��%��<���{n�a�MQ'k���]&�\sĽ���y�n�E��:�D��x�o=p�Gnӷ$'C�v�<�J��xw�O�S����	����]q�n8��R�� s�-+���Q�w6TW�ٰ�θ��).���F���ё1n�ve{���ɷG�	+�n��v;��8ƖM���;lS<c��K�:�t�퍛pn��s�hLZ=����<pOn��]j6�:��A##9�q9m̉��Fq��η�8�6�.C������v{\�@�Ǩ-iI�]��]��׊�MF��ÇJ��W������4�l�e^6c���/:�ϵ�.��$bF�Gk��wQX�l��Y��js�u��%�;�g��Y���GaK�R˶����p@ތ^x�Lݵ{$Υ]�Y�;z-k���í���k<l��Yw��W[��ơ��Y�&���.��V+��A��Ǝ���ɨ���mһ]�K����yzh�E��ݡ���vӦ��ۚuf����ٓ�]\��2�a�����n$�]�6<�;=�6/Z�9$�\]Y.����,a�v��u�n��+��"��l�f�<�aݏO�x�:5�R�)���ǳ�2v�cvrun8�����%��=d�s�,�j�.ݣ��e�<�����ieڽ�BŔ9�
.ͱюq�bn��j�HS�4�7.���u����8�zz���nN��یc�j�Kڌ���/��7F�F�<-.��ِ㡸���&��[��Ƀ�t�zy��x��>:�D�u�hgqwK�8�,��.��G`�0c��9�:��.:�G->�@.X�[A8h�m\��9�^��I�1z��EY_U��r6��>���!���u�v��/����j{]���ŷ5��]j8�#]v��^�痨�,�u�듺�s�g��E�˱�Y��!�T�s׮��K��j:S�p��F�۝�-nK6ǧ� e-�v��]Tljz�v�U��㍊⢎N�5gǷNK��&�'gj�v��kc���G��-m���l�3����&��Ѹ9ݎ�pV�9��l�x��D9q�=�6�	��:�����3�b�탍���Viހ4��3�v�c�:�}�(K�� �����nN��mی�6р�#i���Ƹy�(j'���웥Iv��)�-���<�z�C���B�q��KTJU3�5�M;]��nY��>x��l0�ú6��r[�jX^�;��3�)���Få��=�CHj�c=7�/.��ûVz �vN^�O<��q�P�8��:������Ckv�1�Z���i��V����s&�`���5�M�n�a�X�v�p���׭��Ǟ�Zi�v�\{gS�K\Z����nlcC�@��s�K�v{Z]�j,9	���vP���1�ر�Abx�9東ƞ#<xݰ�\cqι�8��ܨ	��K;)��[��Ŋ�u�_b�;>�h��<��3G�P*x�5������}
�4�4�v��F�*��Lr]�Rw.�������k�{'����7V�M��Oq��5�x���]a\r^[l��+gP�u�5��m퓮@cv�U�v
�X�^�i͓z��n�l0�s���k�Z<�s�G=!�Ʒm��z�<��Kp�c���8�:�Gˍ�K��܄vڰm0��72���]�m΋���]ڽ:�)rt\3�f9qP�d��s+]s%5MP�;�P�K,�x3x[+��5���s���q鋎�z�ڍn��ԫ\j{q�Z�l��eݱ�����ϮEv�t���Ny�����9Î��׮my3���鮊'��zt�u�v�%��d�nm"�-�9yn��OO=�v�gt �������ٖj́�8�A���8u�E��p�&¤=u�[pq����n�^M��n$�#�� �ۄ�.=�f�[v.�pwn80��w+Gc9���u��8%�G]RR��K�eu�Nf��f�1��g㥋 �0�ADb������ER,Q ����
"
E-,h�*,F*�#��`���e�UUX����*"��U"1X�(�R*�(�*��DA`��b�b�ieH����,F""�T���Qf5X��Q�"��,EX�dF(�(��*,AX��[T*Őb�
E��X�(Ԫ��*��D(��#`���ATDUH�E��Qb��ED��Q*�#PX��H�Y�,PG���z����
�#�©�D�j6i3�E�<zyc�7�����v��ͧk�����oA9�\Wk�ه6���a��<8��m �������/4-��z�g�[j�.����Lp�1e�|s�{�q�<�Ò�a���Y����%��6�m[<L<!��s=G���6�el�ښ�2��c�Z=��M��܀17�q���ۀ��nw)�7��ʢ\�^{M�aMϭqU�v׋��=8ytcܮ�,�8��.��)��^��K#3美�qq��7[��j�G�>�[v�<���h�!ݳm�1�wM�϶d	)�2c�kce��\��n�=F�` o77� �BG�Bf��66��[4��uAZ{y.���o�~�vޫ��N�+!��v��}�6�m�-۝����]��۵wU�6��eɶ���wy;v\c�d�W[t�q�ݻ`�O[�2=1�NݳN���x.�kR��<%��6|��5������㭙P��Ż���e���v<\aڧ�#��k�u��5F�(t�칝��Ít%��`I�1rO�Xyݜ����^맞���[q�3g�vڍ��ꮻ&6-�����uɳ�U���q�s����F���7�¥���ͮ�ڴXM���h�0�b:�3�u�L�غ�҆n�e�M���<�pY�t�2�g��[�<��%�w��9�X��E7Q���7	�^�r*��vݓw;ǀ]�p!������Sv�_m��s���n{aW��l�rnPG�m�χs�n^0�<�)��9*�L1�p�lm¶����"�Wc�L��
���v�.p�ˍ�1���_�~��}� ��R
��ᜱ�9p�A�4���ݨ���j�,�@@�T��M�RE�7��p�LV�M��wdG��X2����a�����myJ*�~�w]aSw�#� ݐMߛ�
��N��o��1q:����i�8 ��@H/�۾Wf����9�ET�B�ޔI�}B�e]B�Y�K7Po�����4��moO�&(��$Vʘ�v���o��|=������-���"����(�2����ͦ��9D֟5^8�r���UB���Et/McH���feH*�C�?nc�f˚���ϭ1�n;�t��!V��R�@�F���];�U텼�mMv]W�,.��͝t�-�<�ھD�[�!�����1^�s�z��ބm���gjE籪^Lڨ���h>m�&��
\ر%pT�q������NM�8!����@^��Օ�����T�ɉ�u-� �]�'T���N�S(�Ns}j�k�8���U��>�	Q^Cv�sL:L�>I��K�t+v����0^Oܫ3<}�L�T� �g�6�Y�|��,��R��T�e��+��ݚ�VC�nw�� ׶� ]��&)�H���H�� ���W��@D��]�
�Mʺ���K#f�.�E��44�����`���ƅ�;��پ��5��\�=�:1z���گ�`�������Q8��4\�;���ulP".�@�=P�A[��7*ݵ@��ň�����19N6��l����K99:�1��.����o�T��0\U�;c��#p�\oQh5)-pn8�ep�!%^���O�=P��m�W��]�UuB���Eo{�� `�Ϝ�>j�ߧ7=K�)B��n�$e@� Jt�Gpp�ʶR�$R5�x�>�̐��)�o*s�Ƕ���gЙ��
��"r�7�UN왽u���x��P@����]�>�}�{�6t0�b��
v	���r�X�<B����s��0Ѽ�=py�\*�ȫ�uy_0���ָt�L �9V��*�fݮW�>u�� ����Tb�)T���M�LL�����ש/:�b����*�A��/+jb���e�Bk��@{smm�9�����쌽��B��=Se��ʍ<j�]� �B;�u@��e�k�������a ��.���f��.߫��(�f3"�oP+(�R�#$Ssfw�Le�β����ۿ� �Վ�b�m�ҽ�K���z�PWѺH�� ���P&�(�3i���0n9}�B�<��ѣ���=���J|.�+)GVrK������������dUA��:ʯ��js��g��_�����ۍ�3V$����x0*�S�#��n;v� Z�米g�n:�	��ړ��۹�ݞ���٤�Fͧ�����s�v����a��AC��X����r-�� ���W
$p�]vyy�v$;c�>sx�^�O5zss<]������]�S�Z����6܊��a�us;� �CTF'M���z�? �9Z���� ���	�4P6r�FVv����A7¤ē()�ٙ%�ȵի�����(�N�ڂ�hDDv�AR���f =�Ȅ#��>��l����n��d	=�"�T\����*棲O��TF����:L'{Qph�����]�'l�I*T�
��p���IQc6�9�TI7�E��.ș�Y鲷#���4���(����h�Ujv�40!k��zwͅ2�@�ۢE�Q��Ю93���u>��V)ǲ�? �9V=�A~�'ёV�NgU���+f:�ݛY%n�h4�)�B�m�M�]#���mv"�E�u�آ7�ϋ�7�=X6�z�N���Uq�� �j G/���\׳�s�d@���ڍ߇�"H6�Syyy+1-��sB#��	��:u�.l���&!!e��H��C�qպ�ڭB�v��fΏ�/W���BVk����m5�C�"��N�Q�U��y���>ſ]��M�K��:�B�kN��S�I���Bo#�!L�]�o m���PxΨ�8	�iOv5����!�%�'�ҢI�	AB�0ԯ]�^�w<8uO/y�.P9�gVR�'s:.<w�u���M��;�<=��y����6?{��m�M��Y�E�A�h/wcT� �|#"bfPP�"4���Ni� wn}�9iv�[�Y׎V���䌽� �TrV���X��䖚^ ��U�ײ�ڙ�yyBj�]��m�5��sbx�q���\��x���)Vss��2��-y1��D��h�Fv����ƻ��N�ɥ	J��W9���d���fdY7��I<��ﾧ�%�>b��<�R�R%�w-X��d 9�)+'o^� ���_��byy]n�6"N`k&��uڪ{� �qD/��^m���^�e��ڛ.|�W�&���:�&�洅�f�>A�Jޑ ���VU���ko���+9����s��0ݟJ�wvs19~��w]� �ئ+h3��yv��,n�=���K���r�[���*�Z�U�,a�w����}� ����s��g���۴݊(�rb&P�=.C�}w�hs�>@�r���;�{���VQsE%Q�|��}�Ƞ�~�}�\G5ؠ�����H�� ��c�_��ѥ�y~o3K�W�Ǌv�I2���^���ȣ�c���ͻ��F��〪WH ݴ �|�_���E�\�����Cnl ��$���0ʿ4X���=���$\�e�t]��w/?\Hh����.V�Y6�ݐ3����d���E�!����N��N���=n���|f��_8*�rRr�5/\�9x�.ƭ�c>�z7�ݼ[v�0�<n$��wvC�\:`��"����pk���1��&n[sӻ)��z�9nkR�JY��0PbNPkL��n�Rkʊ��$�	�DZ[�����`�0��3<Bn�Du�Tq�\V�/�B�l���D�mŵ[1���Kkq���Ȣ,�O�� C�hQ6/�[&/M����)	�(Pp� Ns��x��Oa7��/Ҍ``s��t����IDL�Pnl��Un��$�|O��n�qg/4�vyŴf�g���R
�˱�|�]}!�WxM��wo�Y�l}!�/����q�/��B�<�<w/Pgt#�F�&�C���W�E�Ingnπ=��qw{��ix?vD�z��|���ENq��b:�E_�6��#&�wݙ�7�,�t�뷽��k�Sj��4��s9��x.�r�j<m�Xb�;ٱ_��
#���m7v�������YU���|A�O���j�ѭȸ�y��[�(����)	�(]��EeپS얰W�9��$s}��nPu�@�gy��qƒH�����I�./���{��j��(A�Ҏ��5�W2U7��x^y��v���in͂*��G�#�IN{ݹ��3��[�E�Y@�	��]�<f�R2�D	=�b+PE�l�v��
��I�M�A���65�M�s���}��\Tȩ�qUWH��E���}�φ����/��}"���q�B�-��w����������<Ү�/�{�7B�RM�H�q#�mcE����v�ٻ���:�!��uc�����?4�;;q�#P���|"v��<���vjo����{����������}�ņdKz[o�pw�
�&n)ı�؟�ۥ��ظ��% n��s��"d���V��L	=�v��<M�㽸�/{�q�=�1���v�:�q�b�
�$�����ڻ8}t���=��:��������{y8��_r�#.�'|p��n%�|a��j��&�0yֻ�vv�<��^�5��^�:h#޲[Ĝ��}Rz��×�Kq�Y�r�Y[��3r=�wh���_q���a��״�ۋ������3��a�������U�i���L��>�f��w��x�$��<�Y|������	��f��/z�o��Έ�sP�g<��;��4�4s���[9��!���lqٳ���!7a�m��L� �3�<e���
��j=��׼ZV�A��=�x�H"��7EZu�Kĩò,�=fpl�@���h���������D�" 1U$�%Q`�R(�TUE���	mX����b����DT�TR"
"*+3.�n$�X�P�*Q�Y*,+Q"��U�q��m��ˌ�R(�Ԙ�0PEQ�L�������eU��JE+YVڈ�`�bbbWZ��b(�Q*Fcq!��L`Rڨ(J�b�-k1��E�ҷ00EUV���eTb( ��KQQp¨#�e�I���QX��V�2ۆIV��=�ߐ!g�(/~O���r��Q6��6M'6�uv�oK�"fDN�H}����eV�X"��P$}�y'�BdJ�F?��r�Je2H�8Q�r!�u���w{����֨YZ��/��i�M;(�WV��-T)���$�L�wB?E�����d>㼶Q@�k��-,A�� ���Vv�ދQtA|׺�^�<�c�����cX�(�_í����-|�i�S!T. F�R��ݻ�>�i�W1�»�!�M�`�u�^=TH$t;���ҋ��Oc�͑�05f�*l��p���^�"�9����_�7���f{8�]e��9���A��Q��"��e����ۛy�sslX��WC��^SP�]�R�D����z(��n���o}�������O1Z�_bp��Zt��Q��7����Q{Ԃ$����I��:� /^\m
�w>O1�;GdRHĉ"�:�F_X���r�?vb��������y�o^�S;<jd���|�]�3�@D}|�/OC�{^�Y���x�8�'��
�SS@ļ��TM���hQ.6�>k�!�g���^ڻ�I�Nq������6�h����>p��$�k��r%j�<��pڎ�4�MS��iR��Z��3*z�K���a�z$[������V��L��k~��҇�g�d�~�����i�Ƿk*�/A\Z��r�1��[���w[P���m�ܚ֭�=�����k�oWB;���wk��T6�v�3�^�{-�캌�p�������<�x�u��[������Ӝ:��v��@IqjY���&+���!�\ܛN	�X��\ti��ͨ0����Gj�q��{�(0�*'�Z\��z�"I�iN5�Gf��n��q����F*�Us���k�Y�ɜ�|��::�"O7!��ݒz'���}Y�ԮHU.��͐�HZί<�iu@�܄�����b
����#ոFQ����j /}��W��k�]���� �A9W�Z�D�x�����_NR�I��(�K�^X }����^���;�+�I�F$R� ��Iu�m�q�N�z,��QETI{����"r���@@w�� ���vK�w�^�<�@��Q޶Zc�������r��y=��6�|]B�}!���;����僗	��d�./=(��t]�ӱ3{s9�4�����/M7�Q��qy��US%�(S=-�kگn,Ug������"@�Ψ���	JHn$���K�x�i"F�j�I�ɉ��!RJ���L�P�w����_I���C�Kē���|���Y:'��1jbEN9�;F����l��8�#R�)��]��6+��o���A$��
Í֧;l��Hi�$��"�*�#H���iOV娹���ku�@���$��)��Q�-�sRE2U��\~ɶ7�mY|G���U��L����K�g&k���>��㨉��n�cې+<��W��دv�~��$�ߐ�~�l�նg��J:*�h����A��Mz��+���)P���t8O�trE)Rb$��|�<ANp�DuD�$>��$�[�(��.����|�>v�,��$��h���Ek�T�V�lg�)������*�"Z=��bs� A��Ga�N�Я/&�[3=,�m�}�ͻ2�@A�D|~��fk4�,�"�V&gJݭ9��e{�\��\۵V�4O�-����fߧ����| ��.����>94^<��b�S���:�g`�W9l�u��՘G��<Nj$L��������[�?����e2P�.\�s���t�8�I�:Q$��/m��쌽����rL��j�("ѱ�$`�J�@��R�Q�U�����,D���(�	S�D;���{5uϻSEײ�6ÂʐUَy^��n	�Qd`!�����0$l@-�L@�N��S@�S��Ӎ���.��/���nݢ�����8�|���YGX����͗� [��i������]���`�*�s�&�y�mUo=��{�*�P$��u��qN'�P������a��w�ޗ6<���+Ƿ,æ�GŤ���:,5Ҩ^Ӂ�A�9��/�pw�D5
l���v��ۤ��v�.f����~;u�ܕa�N��\lq���q��}��i�=eш.і�;��:�n���WO�lSg�^<C����c���nuڸɛ#�1oe��n�խ<	�׵l�#ũf�e����CG<�ph�;�/I����,�b�0���c���<��cc��	��{B�$�(�pu���h���!�o��W,�+��n�{���o�꯷��{����P���eB��g;Ŭ�T�����-�| ǳ{;��ck�����l��03��J��@:��]W����$�rVZ�%��e�z��ϜD�}U]���u��aS,={wh}�\"w��Yq�{�5�c]D�+TҹQ�Դ�����8�9c�<���Hͤ�$�E�/�m#/ר]���{�a��|!=�c�Pr�V��,�^]��1��>�I׬���˞����$D�<Ťa<"����
�Z���Q���l�A����_�7b5�*JF��B"�J$�;���>:�s��{"����"�l8P&R]���|�TşS�,�n�|���O�l�:q��﫠��)>�`�����in�<���Y�J ]���)a��=�~p��q9�m�ݭ�*�mD9T��18�Ib�8�z7"Ϡ
�&g���!F�t8�޺Wo�7��^j�	�l�v�ӝ�Q����ڀ�s�,�n�}�Q��oi��&����R��7v��j?����������&A����V�g�֧��=(��yǗ�g,k��w��g,�O����ւD��1A�Cq%��ū�"r|Iݴ���$�x�Z�M��G>H�{bzH�Hvv�G1�F��'\�?l�
��j��c�έ�y+�r^�h�VZ|Q�v;u�u���!:I���5��b���+%(����|��^P]|*�f6�^�P&��& _���$�@`ցhK�����{מ0>�6B<��(]\73q�:I*�
�i:�In,�E�H�Q�ߴ;ͯPnl��˙�F&a
K��zb��I�D�����lL��S�!ho��#0���&hďfě�(y�޼u���7�s��oI�pH�1n�ޞ[J��<�q5���!��^���UyB�q����-;_�w�zyM������v5���D����#)�Jg;���@l�|��i�N�D��v�8����d3��kb���6I�n���\ۗ�o{v(�:��U�vn�No������u�=� ]s����{]��2{p����)���d �ܖLг���8\q�7r@�v��~�%�:����(�����@3�۹U���̭�!���8�/m�C<>�����s�~gP�m�_"*I���w���0g��xu�����w��ϼn/v�;3��_�3�\C�}��Ԟ�����_��@^�tzi��=<�����y{9�篻�lٿKtd+�|Y�� ���:�����/�d���eC+sx�6׸g�z�3���+U�ݲ�$엥E�<��;��|��zC�i��վ|'_���e\r��b��6B�ONc�ݗ�+���2ӫd
c�TN��D�O:�O4�>�Y��!晩q��M>7���-�'������|����믛ے�#���A�۾���ۛ��>�=C����h�tM��� �Y�,~�=tzT&��sK��V�K>���[�0�ǰ�W�]����������䢋uk�})�:5L��{'��2��U��`v��1�ڴyla��>yKD56�z�~�ٳ޻�^;��3���O6 [<���J}��	��~�4��>O)\�+���4���=�X��hE|�%��ҷ�����9p�tow���g��%zO~Փҥ�q��gS�]�H���z
<ư�Q����w����_Q9�gۏV��eE�ԥZ���*�G��P�3!S��Qh�T�l�HڤQAV���@�r�5ĭʬ��*�+�AB,Qj��+
Ԃ�j���j��`��"���)-��0�r�)iG.c#Z��fRQ��V�Z�ҍl��
+*m�*"�r��1*LLL`"E\a[[��QLIX�Dd�ѵL���X*0-*�YF.2e��e�ʘ���\�1*���rʩ
$�+��-���P�
��̶��QVc"�e	�U�*�Q1�����B�10a�G�j�[��뢒�����;n!��e��]��fw>^�	�k��ۮ>�c������r��i4��=:�v:��]�ܚ�V[:��C�v�hy�l�m�T�w,��&c���c��Y�d췷�n{6.6-��W���;r��Hq�S�]�G�n�ϗI��x�1�qքwA�	|;��[m���H�d:�N�=�\R.��6�\F6v��X��:������e��^�I#�8v㰡jѸ`l2��f3��@�n1jp�x��O��3rF��l��P�y����;\�7ku^G��ƹv����3�vy��۶�E�z74.�}��On�Uݞ���au���c��:|��r��Ө�a=��8�Eŧ��
�ӱֻP�q�ٝ= Tf�<�#ۉ{<��)TM8�e4:4��sE4��S�7g�yށ�Ķ�H���أ����Խ�)�]���v]�^�ۮ�Nv�c�e�ҹڹf�M���N{ob�i���Ar�g9b��ϐ����v�v�uЖ!:i:Y����IW����On���{=�Wd
|��:���v�A.��<[9N����l�u��v�ԅ�Lg���;U0�������\�m�Q۶-���Nylzfڃ�!6^y�����2��Vצ&�g��n�^!�֦��W7n����6�M����˦�z�S�]�6K�ۥ*;<ӌ���'�����V�nu��N;���^ͥ�y�v�$�n�����>�^6W�3ֽ��}��k�/m��S���zK˥���ٳ�9�nwZ��ن�m>z֙�m���pWV��A�{�kx�v㧶,=�]m�gjU�.ϩ.\^-MU�E��4IR1������[�ﻮ|}��H��e�x����=����s�jQ��� }��~̭?>1��?[P>3�Nf�OɎ@�G����7���5�2����@���ѱ!�ne{��]m��12*r�:��fm�`$�Zf�U��C͐�#m��k���B����%���svDfm���m����(���ڏiu��B'���|��=U��|�d��:��9���3tN����ZU6�j���-���(DK��+�֝ePv;d�v!�*&!���{T	�W������$���L���2��>ng��G���Y���3}�9</��"��N�����R�)�SS�峑������:�#eG~��l�ȑ�����F��o�e��}P���}Lrs�!��V��ʀ�>4��\�n�F����Q=3�P�2���@�d[U^I��+ĂKm�Ȏ�ޭ�	�uAnlA��B�U��i�h!����$5WU�H�s�K*d�r�f��,`����QNtQ��[��L���c�*�K+#�9�z�1R����d>�D�Km#�2���9�XH'�]�'�����鸹��ȟ_�>�X ��۟f#���Z�1�\�1*L�(��A ���x]�gLl���b�0� ���Τ��C�W��R��Y�i��핣c��Ԩ����������AϮb>���}Y�F�:�\G�QO/]4���� �M�.��<*ۖ�S�7�NDI�L��T��H=�d��v��e}��	ײ m�^|7�can�ɋ5�32"��꼖չ�y�����4����ho|��M�X������9ܑ��hZՓFzʢ��"N<H��"�D!*&�N�QZ���y�:�h�d� %�ݵg��8��� +9P��d��7�{��=�v +^5�-�W��^�(��vX>Y�r�9Dj�-�e�2����iKm�$�[����Qw�Of�UTLa�!Ҹ���J^tjt��f���U1{d���p�v��ZzZ��gA�Ծ�h6�"�}�b�s��~%�3��)լ��쀛Z��ZO��Ѽ�s���wv��-��9½��;�B������F��S7��G�.< M<续6I-ܣ���Ɲ�'+R�f�B�32���o��UŸ�o�\��W��X|Cw(�ׇ{\F��F���R�B�GN��A�B$��ħ,n��6H'��Т�nڙ��b�0ݲ��d�<r��P"�ܿ��*��:eo]��}��΃�W)�*6��](�"��kL���H8�B� �9�}|�q�;��>��;��㣷�חg�^���>�ԑ0c��p:t����[�C6�;��㹻���#/ �=�E���	SI�1 ���n��J���ĭ�\^ѫ�Δl�S�=�9�r�z�6�۴��X�q�gƓ\�ʘ9� F���P	�h�����E۴�׋#t�6��7m�=Ebscn:0`�뭽���Zw'ɺ�l�q����g�S]$S�k�hG�[����*�2�w�K*�*!�HEe6���F���7�(���D�A�G���ӧ:�y�ZM���T/[�����Ӹh�^\���T�lsr� F�b�^*9���j��[�3��)ʚ+f��� �h"I�6�6j����}�8{�P��K�>�Q�GKkg3����<��[t����|�ݼ�k|ۿ[u eSj"ARa�Q$�cK�kp�! �S��ܯ��=��%o'��f��>&9�vUtrj�k�n\B�rUe7����,Y��uD�y����m�I�B����� ^9@c;��@�D��1�ꉜ]�q\^XN�pc�׎ޕ莆_C��(LL�3V{�nc5b�����T�i�5N���   �۟|H�ix�z��@�����۬�ufS�"�������� ����~���dN}��n��|��)%]����*��>�AM$A6���y�ʩd�vMz�hF���RQ�%D�k�W��ܠr`wz��wKʳ
!���{���*ƾ���;UQ��;$p�>�b��ϣ���Y�Vʝ�����%L�!l�(���Q�r�5����M��w�9�۴�L��%Jj�ۨ.a˻ye�V� Iٵ@�|[���#�rmKP�͍4�Eq��.g)DO�c��k���]����
����a������>�=`���|�9�	���i�{�r��v�cz̾kG=���1
�=�$	#���>s�lڃ�u��3:��Kn��gZ�7�6�<���C됁'�ͻڪ�w`�c��j�rRJ��1;(I��[1SL.���eU�w+Ķ���������U�V�Q��K���볂Zr��B�&�S�(�qҺ�m��r�| >i�U�����	;�!5[�D���.�6�7���gEK�H&��Aݑ�Ҿ�ԼۼEr��G	*T{Z�����xŢ뢲��>/n|���:�n�s�h�V��"\I N]���m��i���"����I9�$lj6���7+���ٔF������TF��ק6�dDc�;?zB �O��.��`煷F]f�kZ�(^g�*	�q�E���V�@����1c5	�u�;T��Z�8ۈ����f�ץ�[h�z7	���Lѱ�#������ob�H�ݗ�����G)Ђ_$=)5�GI�Vl�v�-�fl���^4�'��P$f6�5M8�Hi>)I)B��t�ՠ��wH�z���S*"�  ��K�[U�7�JT���j��m�.S��kI ��C�/kF��(n��������P� �_+*yk���UCq%z�,w�߹A��P��{�i�Wu;��5��������o>E���]�� �B�9�
�E�f9]e�؎�f'X�{s�ۛ=^|��"QF��qn�.�=�yx�*�T2q�[8x|�����2S&f��^�;��Yu���s�ihW���\�G]j
{p>v�uړ��Ɏ�wCv�qj��^��,�݉�Cm�]�"�ݮs��]����-��Zƥ�{t����n�iI�-E� �����'`�*���"H/3P�oI�z*�x��� <�v
��d�\Fۻ�8�Lء#[��-�!��bx�R ]I�q��V���  +$�L����v��[�<��%H���v\�nn�wH$�UU��	6�+}=�d���t!S�*c��I�sr]E�;#����h�n��@��m]g<���������ی9t���׮��V��	ZԈ�r�)��{ⴎ�>{s~>�t �����w�{8	7Ҷ�������ӸM�uz�8+z��Uo.=܉�2�(�=�N�{C�GWc����;h��*5_):�pW�R�����ѯ�$ .{��6�~�����O���E��:��;�I6�����G���
^�#�[�^@���d:�@�H�E��;XްIQ ��LHG����Z���Z�2�~t��*.|�%�ڨ�ꘉ�Bp��Xm���Y�Nn�7��p�T2J��s���ݟ�\�s��JD����?���a	L��>�$n�����T���j�]i��!��8�<A�����w�0uj|� G<� �:��8�5�׵�
�)�ܫ;%(ssmY�#���ޖ~��7�Wu3p`v�4#��c��$���y�+9ɝ���K�b{����n��|(����L ����@��w�����7��lH~��!�!oԟn5N�<qfY����>��t�����ٛ�7�H�wz�� ��������˼�/A�;X�� 3�|�F c��}��ٰ�=֬؍����v���7�t7��h����[��l�8���4��Căz\^p��x��$[�^^\o��2�.�[��ѽ���v��e9}��/�<��jͦA�]�y�`Bn�ixt��|q���]�[�Ǽ�:�<�A��=�*���{�vj:���=U�
�t��A븯
T>>�r������.{:�	ؤ\`��{8U{'vө��ܻ��2P�]�&��G��w��o{.9�u���Vo�ݥe����8�K�7��\�7��
/���,�vv��<����ny{�d�՗6���M����ʫ͗voM'�zz��t�	8ݫ�s��o|z��	�xʳ�j�&5e���끛���z��Q1-iDKB�Ķʘ�R����EU����e�e���C-��b"0(�����L�+1������U�b�ԱV�kb�W2̩[h����`�☕���"�U)`�2(Ujb@PȭJ�UB�"�Ƹ����
���C��
Q�#�Ĭ�Qb"�X6�j[B��!�dX�b
&��rҴjAaZ	P�Z��e�bVE��`�FQ1�HUG,���jQR(�kT(��,Zږ�����c�+Q@�����	L�KmX��@$!����W�{�������	�-M�N8�������(�Z���H�k5��$���뛎���#jD�t�uel�`��tn�+��`%7���4���H;��;+���� �&N�ݒS�}�ۙ�wnr\�Pv9cw��b 0]��0B'��ТA �5���j�0r������>p�N�U���$c�"�@��$ �N��@�q ��J�z��Q�)DM�r���C��f�-�B�%����1D)��o^�-���nm� ��$�[}�UĹ��E��=�7zA(zfL[޴�/o�>�PyZ<�U�
�j�ea�'O^��́�x{�>&��T	M��AWff$[�+�QT�`M��>�I�LNB���M����U*l��9���T���+t�)UEu��3�/z�J�u��=v��>�l��^�o
��O��`��t�k��MG!"�V�5/�u�c-[�A��-�'y´����.+9����-ZO2*�\�߸뎜o��nX!f:>�ؔqg4��D�-��K�#�"TzA�r��z�G�L�g�R[�)��NI:���B�\�nf�\����iD�@.o�������ַ (UQQ�7qh��J�D�.��Ƀ'�M�c�+��qȷ��ʡݛ}���$f�#�>�����v��:��7oG#P:�f���I��3�������յ��^{qt��Py8�g�=�T�&{v�7\@�ϯ]���4gi�Hng��Ir4u���o\��m\F��m�7���ܻѫ���`��E57n�'�r����W�-��dL��Kjη��vk.��y���Z��8�%�
�B��>���\n>Q���$��i-�GEyD�Q4y&�q���n�	1D��"{[�@����^�����@�\�:j9���h"	8����܂��h\�� n����1tuL"RQ"�q-mv՗c�����$�-�Q$�pWu���1-���DL%14w�IfD�{K�f�Z��3�"[Ϊ �[�w��$s������k�viF��@��$�A�)T��}��	�)
#e�Iy�U��[����r���e��þ�lV�	�N����O%���[��_���gt;��sA
�w�aW�GՖ�;RyUA�Kw:v�r>���=�۝#�~ﺨ�	/�D[��z/g�Rɵ�q^Q"H藔||�	 �}���v�� �Ǵ(��I=;WBFEߋ���[����A{� Iz$��P��M	8���JJ'�a�I�s���3�B}��s]| {�Ke.�x'�V�U*7[A�Y�[n^�t�֕WM�*���S^��2.�9�pZk��I/�^<��k��"z��*�#6�u�DM�Ok�>�ʅw�ۻ�j��wdAa~�[7y��t�>�2q8�:ހ���F���{{��0��&vP6�9����{�!�)Y��r�cH[{pc+7�q}� �ݞ��?�I ��J[ ����h�M���}\����m�@����ƨ�Q�NO
�*:���6�7{j���/�q��@nl� 3����r��c7@i��7�vrp�U�8摝V���5�y�T�	V'���M�6 ��u@کY���.�A�ԏ^eJ����˴���]mZB7r@��P"�v��_F�:��B!H����B�B�I�է���y�FkuD��W&㌜��S}v?�5�>���׉$p���W/�����P3ӓQY����~k���.Y�1<g����)M	߲9y��']T���=�Ju5ٯ�T%O�6��ҵ���f�֨@�m�>�u�I�얚�m:�HW�v9�z��p�q{%J��c���̱����}����2|I�Q�`�g��i�@���͉�(BJ��I,M���ΥA��Dn�_�w/1�y�/��T���U�z�Q�dzJ�ucs���j��86�(68��h����n{��Gz�係E�	� �uPUvޔ,���47d���{6��f�_�Wb�/mQ'\I�7,d���R�����F�V���JF�ל
���8@�Ȳ�|�{��D��^@�+#!�p}��w1����9���i�|���v�����BR M�b�Q=V�r�ܛW=���h�r���ێ��Ѻg���<{<��m���Q�;\��˹絚�Q���$����]�Ͷ��ݝ�4��uR����9m��k�F��q��������M��O[NGl��ː��;�Ǟ�
��5��{b͘�<j�0��	}߀�yD�Q"�{�P�I��Gvм��7溨Q%��SL�HU�堉�p�\�{���$Cm @;7ѻ{��/b����f��Y��D#o�Ny�kb˜�� Fk�wv�f.x�R:���krV+��>�� ��P3���'ʿR�n:6�Pv8��h�����J�iz�K��*G1��n|�7Tz�u*��31 ��� n�3۳g2�GO8glr�5,p=ο/Z�!�v�Si�:!�C��Ψc^�W
��H$����_�Vj����S5���'}�Ŧg庲ʺ8�ƾ� V�eeE��YՅL�fa���1�vd�����Y�wG���K��E�g^nU�{�ʥ~{���<��H�Ax���
N�r^uS����rh;�FeD�vzyy^��Dlor����;����)M�А��!@�I��Q܉ ��hQ'�iPڃ]4�ă6���/L�J%)�.^U�.c�{2v����j�wn���3��K��V���e,�����0�8��u�n��?ǽ[�+!Tݫ�s��M{"ҏ��t���_;��5q�n8���!b���u:⽻��s�h �k�7A[���_qjk�>9��(K��f둃M��e�Nљ�c~�)��s�Y�qg�Ъ���t�m������AdCS1Wbq粑E)15�
�����{��W�O�">��D@���� ��E��3*%	�\��Do7��ֈo���p�����'ʹ�O���pk��X�ے�l#��(CO�{�H�H�����U�^�VWkx��lM�\Dmϧ}����wv�%�Y�Q��q�V����5�Kt��r�)�οK �/�)ۜ�oR=����l������UU���m�8�~�qذ�7T@� $Վ��"�wzkV�m���96�����ƛ�gr���Wͧ���OpuC�8�G`���Wm��e)��{)�6�#l��
���q�(B���)�s傜�z]���0m��;�=�9.g�Y�`��C�?>Z �z?{���m���T��ܴ��F����4���EbUU�w�ZՕ��/��/���I�Y�Ui(��of��4���:�߶�,�{r�l�t�����o����Y�WA�}��fQ��!Z�wc��\g��u��Zc�X:QAB��׋)i?��l;�������{c�n]�Z�`7��ݷ�󨺧#rW?V�m�ݻ��8���;���?�{wi���{]��6U�#2h�]���+�ٹֵ��m��v���M�����^�8�M���5�G���ԓ��X��!7�n�{ݺ���9�=�n�.�}�m�ߵ��ǖ��l�0�6�v�շ{�6�EIv콜�nH�%}�95��9#Sv�/����]�`�#�����{��G��ު�T��a��.�Z��v�vW����o�q��ޞ�@���ɶ��9g��͉�7��s�-ח�ɱ��1��j�鯷Ϊ_�K�DWj�~/{��ױ�2��d��v�6��\����c����߯�ov9D�5�ӛ����?@Pu^�����V�R�G���~h�k�;��ucO;������e;�Y�	wo�T7����jb>������y�ct|����ߺ��ڻl$�3\���Z����w�!=ۮI9�v��̹ݚ�2��,�<�Y��i#�������fXJ맹��ṽ����9OE���z.�]<���v��&����%�R+��*����d'�n_X���i�`��N���eb�[C6�Ѧ�;4qo����^����]�gގ���=A���� �욦�;�����E�\۬�l�o�m>��0���Q��{���nY>��,�.i�w�/;|t�͝�[��7�2{y?,�-�ܛbE�-9j�2�p w�5v1Ր��3���ƺ�B�������G�g��J��m�I\`-LJ8�&+XT���`�Pm�ā��*J��
�����[J��RԵ��QVc3-2�Ҳ,�s,�T���!11�kh��.6-J2)���cQ@��dU��\�),b�$̡RV���a��VA@�a\̹+���)�dRV����c��ˌ`T+�rⲰ��h��$S�Ls
CcP�LaZȱ�!X���E1���b���R���,*J���P� �����U��(.&7R[k�ν��7��w���=��:ܗ*���۸_ [���d�Pt�@�r�ƃ��vc�Ltz�5���6�K�7	�[kun��mp����dy�#��w'�vm'3WJmF�-�g�=����+j��r]��}�F��~�]���lu�.�N�Om����l.�Z	�"�]On롸���ZM��s�c��E{���zz��$ݖ�h86���tqk���� ��'{N�����ӛ��l:w��F�lE��O;7m���'%77;5��m�Ăva�`�ש�\�۫m�OV�x�\z�ƻb&�c�VC��{��TB����:����NC��Gf�cg��n5�9�:�ѣǋQ�=�����"t�d���v D�j�s�z��ɸ�g���+���g���v��j�����0bx �M�������,�(���p�PN��mcd�[l���7f�q�S��ےW���G�q���ٍ';�؝�;���q��n�p�-D�1K�k��s�bqa^��ںlY1u���l]<�3�+�g����I����=�{o-�qƛ�<���S�mlv����t��7��G�.Ę:؃�^Mƻ�� �gvL�m�u��=vu/�QG�p��nη�gq��civC��;q�v���U��䴹�b�썌�mq<E!CVӣR����9��x�=]8y�D�؇3����o�6���	Qn%܇%�,VƳ�{��{�����|h1����|��Y�j���s�ƛh�m��3w9��AI�X��w���ն�i�n��;��3���ns5ۭuҨn��52uO �p7k%ҥ8��6J����R�)t=�e�m�X��XWC���A{@�M��A�k� 7cy�۹�qIzs�'g=�M��r^k�1�P~����Ui(����ikM�'�v��m�\t��[�ޜ�d���u�n�E�
DL�TIn5A9�]��s:;�w;v�m7Ǟr�i��qF;��=�8���]w�����tHܕÏkq���m�1�M��ʶz��m�ɍ�����Jݝ�XBP�*Ո��3���ݪ&���v��{D�m��v���{L�s2g��n��M��<��!4ݧG~l=�w{���s�W*�ݦ�m�y��'�����5Lݓ+����[klr6�t�Xó���.�8�sx���*K�=5��rG�tM��ۻl�J�s�5���m�k�y�.�H��PW~�i�Q*)�ƅJ80�/�zg{A�0�''����Ƽ��%�������˻�ju�?t����{ֻ�8I.��n�v�����E��~���lm拞�);���C�j���'U���u����� �w���r�_q������{�_{Φ�M�\8���mx��f6{Έ�m���ݦïu��ɮ�����I�����o�TV3f䞻�i��<��qm&�:�m��.��ݭ%����^�mg�]T"�l��jR�\kq���'g�صv���UP�vg���,&�)V��g���͵�]��������'^�]:�Oy녫�A��	G\*�Hcy|���Y���o��;s.���o��%�ۛS�o����9<�47J�J#m��um6�~��[m��ў��]�ڷ�x����%m5�6੿DS�Sk���^J�PZ	Ef���'�eNYΛ�����m�'�ۤMz#����T.N�F&S���R���m��-���riv�m��~=�P mܻo��SwD�����.�l�#˧T�Q���vk�4�m��{]�q̼*�{�ct�k�@y7/����rZu՚�n��QIZR�)�{ռB���2C4�3+��6�ouț����|��ˀޖt�־�._Mb�����v͒I�}Jn�;9�^�݀f׈�m�];ܙT
n������
����!����{�� ���F�t���/U.;pa(���W�ӵ6�hk��5��c��~�C���j�Eg�$����}Ę�=qUZ��B�z��X"��mV�A�Tʞ�VB�����#a� JB�<!�EX=��>�
��������\h$���>�i�ܩ���d�ĉ� ��b���۞@�7�^�)�+��Χ=XHg�w����pBl�i b�Fy�	/�XBP�*�-H�/"�����N�>˽��-�ksm�rR�i4��mg2(��/�s2�Ǻ��+�Ģ�m��Y���*.�%�o�܌/k3nB�ԉ��6RȲL�At�٨8��y||����C�S:�_;���H�o%N�p$Z܁.k�$6�`����ަ�}�r�g��Nϯ��T�NV
Hw��n�2�S�&2	7�|�ů9��Y 䕃P���:F�K���:k2n�jH�y�\l��z�]p�c;v�	����U;m<U�|�=j����g���F1�哞�X�ӓLY�]G��㘺��nֶn�v<�r^Zv=�"�c2����M6�Q���n[�v۲��'���.)�#H�#��{����$�9���CM����$��n���v��Hv���%(��c�p�z���u8or*Gx��A|���1�r�MUd��B`��.H�5�D_;�ν����!����/c��%&��#�ӫZ]�m?p@"I.7a>t���"7��R-�fsҌ��Ѐ>��K�SX	j��7v�=��o#��Ӳ�'S�s�1�\���m:�ݒ�%��c��b�X:�ϟ�>o�ל� A��
��r�9�l�ݐ,y�D��DJ*�oQk�vr�7�j���%���W�[��IBb_ɯ0�p�f�\��x+����7Lg�cbI�_{�*w��#t"|H���&�)DE6�N�P�#]=o>�E2k�9{�� ��� F�d�y�F��T�B��Ӌ�p7�,�'�
��i�D��=���}�N��=�̘ID�ύ�D#ٱN��̼�#޸���0]�m3��#�F쑦��
;nk=d�C��tU�a♝���BG{N��wd>��Ù����չ�A��7��jެE���&$�Q{7��y}�҉$6�$�Q�e�q���8(��U�5�Hג�H=ۖQ[Z0�^��1x��v��3�;�36g��\���8q3J�	��`�ed��]��ToG��O�gH@��������H�P(}\|���Y�L�^D���D���pE�Q=s9˸/}4�$l�%V�j}��`3{8E_�=i�;D�y=�gw53˺��Yal����m�pg�����[��h�Kw���/[�m�:|�$���oQ�͒�V��N����L_���LK��NW��ON���;����N�z��w��H�X���� 4�j _�:����. �� �u�RXjꍺ��7n�n����d@/?k� ����拐R���[PjI�l� ������2�;�d�@�i5UQ��߀s9����)Jy� H�fE�{a½��{�|g�;����ߓ��K/�V����3������7[�æ&����"��'��Ȕ Ýp#��>~����e�wa�m�s �׌�� ��9�A�غ�k�"I.5�^$�h AU��g/n���[ ���QJ.�'��ڀsK}����z�+}� ;퇬F�eY1�4�ǝ�ͤ�gl@���m�ruqqS�j��Ŋ6������Z����.��Y)����A	� Gy n���^O8��\��U�%��m�]���GsG�s�חxP\o��(=�4,,�8��c-}��~����#�l����W|A=�!�'k٫m�쌨�/q�wvh�998��96�'��z����e4c{dn���A92��(���;[qWt��7\�ga�1b���ݖj��l��-��r溝ͨȝ�>�ف���u��z�ou�=v식p�%��r�W]5����z��v�M��%RS��~n~�D����i�����n�|T-�;�^ݸ�ࠄɏ���}��{�U����gj�wd]�3M�.�M~צ*��$r5ڮ@f� 7��&�C�͏�Ffτ�fQ6ss&��	��ryſY�'�ϳvpC��b���Ա��ב�Q�Xi��מrZ�M�S*�7r@��\/o�-�.�\�j���6������j��]��c�X:QAB�����J;������p>>���9�T���"}��.��:����WC�^$�����އ9�e�j�P��tg�'ۜA��WN�bK$����/�,�ݸ�s]\ f���xx*��> �ߗ���/MԱ�f�Es�Md�TG�!쯰浈~�]�5�K��x!>��5���[h&��ݣ_�(`5� A��� �}���.iVuy'<T#�i���{V\�m���Q}�\EV҈�q� ���'a�U�����m�u�g����`i X�v�}Q��3}��IA�'�r�#�� �(��/q�C,䪴#_q��K]PuQ�8��|�2�y7W�#�AÙ 6� M�i������99�;dU*Ǹ� ܑ��9Q�dg��}�j9�{s��d��P�$����
w������΃��v���*�t�׳�Χv.�΄2*]v]����(<#^��S�����-7M �g���/�*�{uv��2�}QS��^|9��C�E�Fc]��>������Κ2��J��p�@0�ȝ����1���,�\"�nq���쓽G�p���N«�gd��vrH#8=����)�֍��5�5�&	�Ul��Ί<���z�"����֏I3D7�><��M�|&^û�9:߭����zts��0>����l,O�=��c����T'���F�_g��.c�O���td�Q��(�O<���;���܊�������w������:�w��.I}�<��3�w�1/eWpt��wN�=�Y����{�R[�}���=�=�r��k�ٴe�7�G�e����*Gő=v���
˻���ԧ������Uw�3����7�ʕ�C�*d<���'�O`'\�О������GvAˉLL�r�0�-J�Ir³--���V�

�l3)R̹q����G)EACDX��LE��)6�V�&Z�ɉYC- ʶV�1�r�,R�pCV*����[#��0E"�(�R�I� �E���*5�c�Ę����-b0���R�B�1q�B)�J�0��9�cm���K�QIP.XV�ʊ�mm"�[m�$�֥Adb-�(����`��Im��"B��EXVTVe����S0��$�[Z�VJ�iZ��dF�YU�*b(-��}6��D~3���YQDw���������С�ifmb�l�Gݕ����f�ճ̪t����Ԓ$�Ƃ3WK*�-Ő|oy	��{��\����XWKRe�G(�.����1/l�i��&wD=~��G�^p#����{�,��m�O4�w�$�j���VzZD��Y=�_G���� �r�/)���O[�}'(:��C����H E�m��9V� ��Q��.��sQ���joޤF��M��o�l��D���yk��b��q�Q�\9�x�_p��r��/�-	�����oݸW�4]����� p��Y���3>��L:|��ߢ��V�Mm��?�|{�vw�M�DRH�y+��A�]����m��ځhv7IG
�'Ѫ|5lR�~j�VR��5���u�Z��}�&��̃������$����&h���8H�Z�J�]�}/&)I�'[H�v9�'�n���v�T���y{P���8[�潮�\��vD�Ԓ�WTQ+�Co_Ufr$��@����A�yOyF\nHl�c��9���@����'�uڲyR�̀�/��.�1^Cj�����͒(6�J��z�'��9B.�q��{.�"�.��36>�����l��X=Fw7k0Dt�^v-ً<�]��kzw/6z=4��L����6�:����Cr&�p�����ka6v���
m��q���N�I�7t��n'�D��5�ѝ��mr��m�R`�p��n-+=�M=]�w\��;e�g���b팽��[vN^�ں����=�B�Jo;�e�V�O~N`|6�|{�wi{����[^ ǽp.�2�� E�ݧ{�d��Ρ��^z	��myb\e�oxvA���"�U�K��sv} ��D��A��k��R��
Ti��9��oQu� |CƑ'yɣ=��E�d�V�A+'bd��1� N���hڹXp��-��k������z���k����3��o3�]nu�.t���P��S��c�%F�e�A��H�|�Z�]y9����`$y��w�,k&���]l�}#��Z�,��]�So�Q|�v,Z;�I���&q�.<;��/�oHȊ��*��Tg�"V�"^+����� ���(��y��Ә��3A�ּ�rX�!i'���7���&ݙ���*ķ	�%�![i28�B)E��"���u�ԁ;{D�x�&��Òr�(�I��[R����6��}ԿW�2���i^�G�2y������$n&UTьp����ף� ��I+�)S�~�uj��%b3���b�@�����6��RW$&���̃
2�qd��|�^�p����Wf��o$��C��9�9�=�yK�}y}&KZɽ���Ǽ����e��9������ꡳ�Tz�>��M"�k�,��XFzz�)ѡ�6�1D�����m{�356�K���6��?V�!i���]oj =���N�H�+v����s�	9N��7kė9��ix���H;�{�pЍ9�&B��wy�=�����\���*�S���=�IAڌO�}�܂h�4�R�}ӅwRQ��D�ЌD�5`�h"
ؚܛ�x��N�h$���gs��U�^v�(r?��X��>�f&�(�V�$�i�@�y�>w}�m��ٵ2�~�BG��m����]�Im��;����Ҩ!Bc\kX�K;N;Fi=8�!��;+���1]��혈������>/6Q ��\�2�BQ^<�D��y��`��ɋ�z�A�	|��uDC���ȁ����ծ��k'@�u2�:�B�T����@�ғ�"��"A��5�������)ԠA�Ć��m�--F��<z��*-^��I�r�$w4���Pn�L�6,#!Mi�Aǉn4n*������b
�e�9�w+�w瀍�T�iO���{��X�F�Խ�UUHJ	�=x����r�
�߬fm���Ϝ��L�&q��Y��X��d/;��2��^/P�����Ӟ^��N������|=��@�#O)AO����١�=�g���Gm��a���h����[�ϧ��pq��ޭ���P��+��u3�u��lt���:��ݶ�6���?/{:,['��봻-朙���H!W��K�v�Y��n������*�U��l;��-��U�W+���ٞ�64�:��i~�D�h�Kb����J@�����y�Ѷ�2��Wn�\Ƭ�l�@�� L�܂r8s�V� ��=�ܜ�ԁ'u� w��I�V���&oȸ\rF���Bm{9~>{�ޗ����7�"Am�IQ,hF"B���]>*'IH@�s�K�8�>L�U�ܑ{�-ENG�w���/,AK��sH�H8܀��\jyn]'���+-C�J�E"#�U&�5E��E%`B�sݙ-�ems3�@���5�6�3���դ	k=�6��ߦ�t�	�� ,�\�N�_~�Q�ɾ�Ξ���W�m���;�Ş���:���،�D��Z}�j����S�#�>ݔ	#���r��[��	�$�JD��3.Qm/m�4wV{{�^M������0�m��h.F��
FU��@�inxw�	���'Ʈ����B1���r�d�˪��[�D�N6���hg:���PrB݈U:� lFUI)Q)�:���8K`Y%R�&}1!�o�B$�(	|�ʫo��M�g��{��m�el�ӸQ'�8J����������(OsHxP9�ooT�U���r;��$B=Ɛ �ZY��c)ʻ�9�
nWv����zM�H�~``@穳�
�åv��(�MF�3�Tܙ���S�^�^=����M)���V˗����z��� �o2(��7ܯPK�f�$^nA�
��8��������!�mC=���t�Ց���wV����s�ܿ,��rZ;22��7�~�����&�w�yI�r�
� �#I�{�!/|�D9+��V � K���Ȅo� I%�	;V2&oip�s+��t�ʒ��b:p"	]��<�z&�.܏��_����!q<��j�T��j��\ 7�_rKT�]��묮^e��ý[ފ���Ww�������<�׺��RȻO2�xav��J���&;䏵w&����~)JQ�9�Ɵϙ����v�Z�� �z��/�Im�z߾�{n�ó(�1�p0�%9� ��i,L�:���yȊ���it�@>i8&���-��n!*%�DDHSw��K[�3'�_*�6G��ח�7FU썦�t�ܙ���V���A���>m�ۭ��5%��Z� @{�S;�{UU*:d�{D��r܀�9�#��d ��=�����k���mr5�@sim�WψH�n Ǹ�'ʹ�(c�p95��C�����ny/��x[gu�ᗤwF���ޘo�?G)���ڵz���
���4�t�.��/;^}��N�~�xO%⟯?e]��Dr���qIw7j���k:<�~��Gr���Ʃ��w�!�Ƌ�t���c�	�A8j>랺��l��=A��N�g����\��|Ư`ګ$�*���<;�V�>rs�4̔E���ն^�\z_�_g�\Z�_m��R���j�w�
y��&hxC^��D�wH�q�i��B-�,�[g�����6���{ ���s����x��N���c��>�TyN�>�>y<�S	�'�z�ǋ�v�$ߔ]}p��B������&���N�ujw�Cər��^�U��q0/�H�"zj�y2���УH�MM�'w��Ą�p������v��1
��x#����u)��u{�0-���\��(;fMP�^�;�Z%ܓ���oie�yq?5������3�x�y���|�Nv���G�����/v뾣9N����8���ݝ˫��R��;�̞^׫�Y�}TK��^�f��������Z�1+&1q
˕f2�IP�f8�J��E"�(�m-`-IZ��ER�m���ʕ�ZjH�Ɉ�D�j�`Ql*(V@�V�TbŨQDE,H��%��,�Z�X%���T�Ņeը��Z,R��ib��TS-ĬP��R���U��*Ĵ�����c�Kl��jV�ܢ��mJ�"Ls-V��Y�X�*
ۉ����Q����+Z��.8�W)��%�
c�Җ��������9aET��ZKlF[A���D-��m��� �e%"cU�ZҰ��PYX�A�u΍i�u�kN���4WHݶ�m�����@΍/��5��Ǐv;�tsj����и3��<�K�l���=������8v��:�ь7p�˓n��`�9���uEn��c��bݛ�ZB��aj�α�tv{m8�#[Wmm�����ƍ{���%�M�ۣJ�N=�{�i윗R�!n��n;g���y��ی�#�cm��������'k�����7�B��̝�f
�������U�;,�R�UZ魩���ހ�v5�]�xV�y��9�L�꬇h�6'�L:����]��#�$?�ﾶ��`�G�ryش[Pma��6�<��S#ϷO�#z��3�m���n眻�f�l�`�.�5c<�m�ɭT�[k��Mۉ�rK���!����7۟���]HX�O�H�9ݫ�a�Cgvzs<�F��C���;�q��m��˦;\vn��:��m�#uɹ��SY�-�l<ζ�����7�c;����]����}�:_\����͜�)�+�g::�[�{�N�'c�4S�y�=f۫<v�4kq�x�,��rg����}�ݧvv{��qX�=�=���{u��n9��pcu��.�a1n�g��y������whcY#�v�ہzc��&�n�h�Y����q�M���3rvVsaz����s沽�N�./sƋؕ�����eɰ�a�:r�=n>���:�X��땭Err����ūpv���.�"�z&���/��[�'����=��$�Nr���λA�َ���wi��D.u�=u�ւ;HG\[�.��ct��볋t�_I^:u���s�s5u]+�TuV�u���㱙9Z�sCݺ��Oc����d�2s�!�~���o'�H?/`�o�����}��7��4��m5����zn�T/L���ס)"���H9m�N��#-�t����9����ՐMҕ�!���������u��=v o2O�v�]��BJC.��\���qTȧH |kvP#Kq1N�'�K}��qd�;F�̠�3{��koy�Q�w٭�R���҈��j�M|^�0��X�)@���ҁQ�������M�Н*P@o�y'�t��n6��d��#{�����֤	>�h%�j!����p0À���!���˳�"��7v_\S��^�N�g����d�s򠮢gg��Ɋ*7�4A$����3 �\�ry���gP��u2Щ ����#��@�{�w:�������{�^~֪�5v	�R����Wc~���ڈF=�����^V\�����|�D9)x�5���$�v�e�U�G^�>=풽&�e���R秷vr�v�9L�OP��hQ8Ѕ*�����m��g��(I�}N�"McX�7kH���+�<��*8�vl�@~���Z��ns7�i)�|M�l"/��U�Y�;�D�+�Ԏ�
{ڲ�	��|�oF��]����5�f��d�o=[��Oz��׽x�$�����7��������Ludl������>h#<��*`�yr�6t減���!4�����s�|�[��Uĸ^��� DHSv6���R�)�ӵ��	4�4��`'�{7vrkUf��TW~�����A�clځ�]"��̙���/>�cm���Mg���z�	.��P��Ԉ�܇d�J'9�[$��E(�N�菁q����$|���Ƃ9����J(�II�r��v˨	;�|�f9������0���3r�i�ؐ �ϗ��q/g̨P��02�+�G<߲���碋H�G������zr�M�O�'�M��6�)xU�QK6�">4�p���xy#��ă9$B�E^�L��ϼ~<�h�]�V��$��r�׬q�$�[�e7�7�2)k/1�����׫�<�fk�-���Sԁ�J&oc=4*R���X������+�{�DiK�l�{w3�ǩ�R�D���aÚ� AK��ŪWz	[ܓ�����}&�V��[�{���ܞ��H|�뀀���w�B�Cy�K�lu�*�G8UmD�أn��}�c:��H�7�W�$�rw�s��7�ʤ���0Lf��
�[�}�H8�� �WNg+�4e�Q��ʲ�4�����^�[�.��۰T��
�R.z�]��]�T�g����9�	�G ��h�=��<=�����7���x�*n�eƊQ�nz��D�[�آ����u�&�w<kn��cՒ���G��U��o�n�.-��=]TثUU�9��g��j�y͗����u�d�����:��5t���$��fb��r���pm��*����N���g��e@RZ;�0�aM�ޢM�OǚʬY ]��kk��	坺5�ɉFs�=("T���ndJ 4����r��ʂ����܆"$)*J�Z��t�N��t.�$�+ZD���!&q��LʔF��T�Ѱ.���S&�s2�����;�"���~���^#�uM5M�2�NR4�F^N��:�v3��-�Pw��x���JNՍs���ʫ6�p��!���A&��-Z�
Q1(*H�c?<޵7�K�����*Zͺ%����#y.ɽ5�f_�J�x:�T�W�2gV��Ų�"۔	%�H�dӮ�;�{񅀔�x-�N�&n}�p"Dmd\W':H$�r$w4���zPD�HW�y. '������^��@�y���3x��;.4H�PR*��>"�ȷ�ӂț�춑 �ւm�2�������-�%��uD�M���[�̎F)��i�8�;�qc����zUh�z�Y��6��ʍ�k��.��y�G�^�s����rn�˔	#|�oOs�o���s������/���Q�Di<���r����ځ9����q����XŅ1��Տ������I�d͖1�3o�i��p�^Ӭo�;	���<ܢ���J*U�{���2�v�7$�7��{���ԼH���MJ����$���)f*�f
�h C��7�����9�7Ϥ����	�5X����D�����ے�!@s��*r�H�`�$�$���|F�����e��A��9�&��I�U�`]< X�`����BA!��D�ې���m�L(��[m��8Q�?<�ݯ�6�u��!ϛo&v|'����z� ��4�]��W����ۀ��m@��V�3����l��¼n�=���t_Y	��Ww�a�D�o�?�8#�D��fI����QLP�KAz��*h�4���ڳRl��Amϐm�^�r^���UlV�" ����yR8r,*[��T�_���~n���R�~�� ^bD�4:��	+-y¨�/5s;�Q)w�-J(�[&��&�F���!U�j�2����g:ݺUQH��p�ȁ��w\6���sԁ:܄:����F�f�i�D�^�	9�ߊ۶pOv�ve�RD:�#v��㈈�9vj}�
�F��7<F���W��y^�ͅ���YK�ww!{w=�H27�����]�\��:�b�����d�K��]�8��:n�)s��mLy�qu�I��|��5�Ľ���r�{]N�6#]N�6�M��^@}!�m�b�[�=N�a:����7k��[\������kp��rd��.Gp��&�cwCC6��C��W6���g�E��um�#���������K��ȴ�WkN{��":^'�~Cm���~��84�.�o<�����D���j�w}YmT�D�\��$��H�OG8��[�z�׍y�"A�JE]��^@�v�x�
1�l�uhI�������[U�O[���-6��/y(�u���̡<�-d�e�r�������	�ȋ�n��|mr�0�q ݊{��Wg����=i#<�]����vv��n�a��Q������dS�F9̣i��G���(/��-Z@�\f���^(�b%Ma�� ��5� ��&=������1�ӆ�7�y�b7�w�=�����&GvX7�*�<f���=\j��@{�A{v�A��;W�Ǚ�	~�ʁ
R����H���s�k-�mE�	��i�� �A#a���L֢�{��HU� �v��{�C�D�x�	�w�=T���ײ�������=�	$�� ��a�۪���+�Y.�7��l�݀��thn�r+�$����'�X8����#�}(�[i}��ܥ4r!�/A���*�2��"v{f�P��$~@ ��  ��P6�|[Sv��1X�7R�����EI/����K���%�bcM
����uW��{s/3���L~�]�>�௷�U��ó�=�B>����|���sd�鷽�.n�U�8;b��_nwy����ޞmw��[�C�Q�8���S�ga��;����|���V�U?7D��<��l��\�Z�T�G}�zx=<XG�U�ˇ�
���m�XB�}����'�����WT#����ݓx�f�e�]�lfV=�Og��+���?z�g!�8���H�w�UJ�.-�v�Z�Wp$�dz������$���/v"WI�4`e����'������᎐���Íw{s5��R�}W�ޓtْ)�	����>ݻ��;_>�^�������]������t�M��^tD#�Sԁ�x�F��H�����v���s��kd40d4��}�{����t�)g��a�G	��CMs֏+�x��K5	;�L�̫����7L�V.Ӻ���a���}9(�ѡ_v��c'�s��=§�p�y���6'vf�Ɯ�y�|ךu�k�f�z�����{ܶ�G;����2(Jp�,Ƿ�O�Wf�j�����;lZ�Ab�%[*���b�[[T��AQU��E�*\W��c�k �V�I�Ec*1GPZ�Tj��R�Q(�*��`()U*!P������Vեb�*Զ�-�YQ���l�`������j�RQQ+�Q�
�V�Q-���1#[EIUYX��"��T�F#�D��J��
�Ƙ�m��j��`���֢��"�-h1,QV�TeH�PQ��Q�hZXT�"-�TUb�B��UdQ�[Z"��A-*("���v�Ͷ�w�I��h�yZ�Q�R���>�o�]z�!��j ���]-�9}6v��i�m� �A#v�Az͸F�wufO �Ff ��p��9�����Dc����o6�[�Wv1:�3s�}�d��:(�t�k]�4���2+�'Y�ߍ�$B�r@��Й�S�8ǯ�5��fNo; 7}P�="@{s���9sd��@��Di��&�d��^�:{�K��Z^�v�D���p�T<DD��[\"tv��G-D� �iI���I|��N�׼8��`����<���rg��>�~g��&HELfWS��(%�	^l�3PT�����KQ���܊��m�xQ���[��R5kN��q� :�H�V��Q��*���;���e�J�&��yF�H����ݼw����k��MT��v����z߆�U�Q�H����L��"Ba7fe���B:P�+K���}(�[����JLL�����O�x�̟#�d"ۖ%t��;��J�--��%.��pG��㶵���35��
4��Hi *�����f3� L��K{�{�.��g:�8�B��u�:[��[��\��{<^z|s��@�P�>(@J�L����qù�ev.GWcY��C�M�ltI`Էg�6�.����9�+�ܶ�wg��9X63\��x�1����,ݷC��܆@Tp8������ؤ��]oa5��eU-I�l4k����p�q\�;q�r��^x׌�Ab��%-U�"+i�sժ�2by�Q6�}��u��S�6��ĀqܠAm����4R�C�_)a��޻�^������m�w�0Ժ&�{�"���@#jD�+ݐ=]���������o��
��Lة���Z�.���v��h䔢��x���n꿞�g�m�lC�=� �Z#I��6�<���C=7h {(�}�����������v���$n��,/M�hQH:�-(���w�Ng�$u+��l�E �=�vR.��wX����	o$%��D�EB�^p�<�ct��������h����i��M�ٮ�����9u�
��b�d��gk]�@��m{�8l�˔~�-�W��$	�����5��>G��\�UP�7+[�" �����i�C��&"�*���l�m�'��^�Ϝ�Y�1�}��ĉ�7�Z��1��K��#��L�]IE�"A�U�	��MyU��+T�R@#g�ț��W�Rm2�Z۠)+eRIy���W( w�@�{!A-��
{�d`>�r k��Ii�Ѹ�#��_��}���t����H(	X����ư+R��s �Av0+�h��o�żi�K���)�Zuu� �9yޱ�����RT�~a�$�%aO��<�w�ۂs~�[#t_�̩2��'��7e���ڈT�N�w3 �s3o�%b9�r�t_PY_xQ�|@�%N��5��ed��J�}�&�l��`�)��>�����|��7��!ܶ^oX�]�*AN�� �Af�+('�s!�7z>/:��7��t��*�����60�)}�Խ`�Z�P�N���6�Y++w̆�9��}\�ۭ�z��O3��
AHnӮ}�l���
�=�2V�i(׮�t����-��ۊ�,@Q��\`�y:�v3f����Z���%y�.���s�bAgJ�ISϾ�4��V�a~�5�؅In�����a�&	��z�M�VJ2��=�m6�����3Z�73G[`t5���㴂���o]���}���u�c��9�`M�
�YS�>G� Q���&;��CƤ�q�Xo}{�fj�Z��I;�TϹ���Q� ���d4�P7��t}�>�ۣ�u�0;��HRӮ��4�]�
�=�2H)�{�qzӫ��:d�s�c=�w���ֻ�Ă�BJ���n$�AaXV�솒m
�Y*{��I���G�����`�U���*���4�K�<q�=�ޒ�`��2����WN�K�6�Nk��H�=� #�no��K�.������y��Ce�w�k�+�}|���I���Ԃ�sh����s!�<�*%`r��aXu��}�7�Y�˖��hs#���ӳ��]M���q��F�����s�n
����_&�I	 ���p�ͤ
��Ng9�`m���n����R����f��
�9���*Xo���F]5�ӱ�Y�k����T5�i�z��:Mu�6�hQ%aXVs�$�B�T�>汓q����S}���15��8�>�]̤���G�Y����il�<�;`V�*X�Sη����k�x���YY+{�CI��X���5�6°��G=Ӭ�7Z�C������:��q�ô��Xu�0�3i�X���H,�H[N}�������[��zAH,9�Y$���]���l>9�y�f�*AB�*s�0ؓhy�O~��'�=aX]��Ci7�(�d��w���l��� ���=@�>s����o��P
��=��W,����ػW�)�:\��3٣��x4q}����xz$�i�w���6�%`�q�)(7Ud�R�������k�n�I/q��r<zL���ۣvkXU�����e�C�l.���v�\�n��^8c�y�F��]oS;����^��=�f�<�8]ػ[�N��qv]Y��Rc�����k�l�v`�{=��ug%�6�'�V'P�u�h�{�֝]_�H,/��pv���,�w�u����*K���H,���՝I��C�%B��V�sX�l+�^7�[�u��4��*s{��d�+'��z���L9�0�3iĬ
u��x����R
}�0����y��˚΃��!�v T���w+�tנ;`e�k�%ed�<�0ؓhT���+�맮���_5��Ԃ��
�D�9l��eH)�s	��>��ֵ�s4oL�Ú���ٜ�����˿u��k���i �i�9��u��:�A`[�k�ӿ��5�֯P� �������YX{ϰ�6��[�z��k^ t��o|�zH,Ƥ�`� ��Z�9̆�h;3�睻~�����]a�<a�mr�*���`J����+�B�NFK��kL��R
%Nw��6�� ����i&�*M��~�[�6%湭2m����T��9��M�7����ӫ����a��!�������ݩ��`��I���Ǫ%mK{'��>�r���z� b��џ�م#����R
^��@m6�YFJ��s!�7T(��|=���r�6ö��q9z�u��]CI:B�����%eH,9�2@�T
%`>��:�^����Ѭ
5!KN{���Fh��s!�؁S|�켺34�`t��k\ͳ޷�{�^o$���T�ᴛB�+V߹�m&Щ*����2y�������
�*�ou$?���(��C�.'���������4�W�5��|�Op4�S����6�++%e�9��ACi*�9��Aay���3��-��5V�nݭ�]��o=�i��p�+`��^�:���&|���4�W?T��Y6��߾�c6�R�T���i �'�����$6'{� �"�&����nb�9�d���&�C�n��7x=���`�Q��O�oj񴂐Y6'��m�l����Ng+��U
��N��r�|�>/;���AH,��i�`V�
�H['�wD�GG���l,9}{���J���\_oCc�n�Fh��X�]��fUM�wٹ���s�����w��ێ����������H(m%B�/9�i��V���^�ۣY����T淁�O=������
Aa�|�i�*A`<��i���,jAO�����[o�d��9�2M�T�~l�^]5k��c%־֙�J�2T*J�}�6$��I�+
���jI�*J!Y*^w�i�l��2�T��s ��s�6k�~���e���BY(�Ptu��I%ݒ��:~�?zP֭���$�����}��i ������H,�]���k}}�3Bs�rCbJ�T+�>֘m�a���k�f�n�w�
^s�6�FVO�ߝv����>� m*J���߷�Ƥ���9�i �k�~��?�\P�b�_J��G*�@t�}��6�YFJ�T�`H)���z���5�>H)>B�T���i �m� ��s	��~y��ZTLU��0|'>�)}�dDus��Dx �����
�S�������G=�xYt�ۯ�A��0:&�T��F�U<���w
�F�zF^��9�g{�{|b�n��-�F�->���N��J�w�5�V��yҶ��k�i'B=��2m�����=�P�����y�{<@�V����XjAO<� ٺAk�s�j5��Q�~�~N�\��-�t�	�M�K�x�v��،�Ucc$b n�ν<��љ�_��8�u����ͲT*J�s�6�hX�������N��/}s��y�v�ؗZ�Zd�+%eRQ���v���ZG���%���ɿ�5��<zH[Hws��&���}�$���,��4�h�d�9�9�m�� ��ם�Ρ��z�V����e��[�^��NЩ����%ed���߾桴��+�s���:��s�����F�-�}�l7H-�
؇;�5��
���2�w�WY���kLo�߽�����"�R
w��v�i ���=�:I�%B�T��z�#�&��YP*T�9��m�w�pn��j�봂���5�=-!K`>y޴�]���=oP;O
�>�4�q����>��u��%B�� bG��+^����P���;�~ȑ㇭j^#���;Ktf�҆�S_���s��{6iW}�Ӹ��`�J��&�aO���N�aݳ$��;���3����An�����X�3�ӲO
�����ת�;�ݯ͸�٭O9�0l����(�uj�#��<~�}L�v�z�xn�šhG����χ+�����3�W<,l�..�9����w<�M�Wh͒E�_�/f�b.^�_������]�0%�|��G[\֎��_f�^=C��>�pM���zr"K��x�}�y-�n�7P#�y����&PP	�A/5s�Mc���ϳ��{p�AG�_��ūtA+�^>����x=cl|ņ{�{�io�b�a�ZK�d��7v��X���{u�Q�t�77=��z�ݯR��������g�P���3O����'rs��b��+�7��#�~Ww�����%�>��q*2sʀ�,��nB��
�vM�x[O=n9���xc��� C�yX8�sѹ���U����|�v��{��=ߺ�^�m-���Җ�(�-,dm+��#k[Tkb%��znذ�X�*U�B�`(�l��VV��*�h�EƊ��1r�"��e*)P���`Ċ$TQDH�APU�W-DQH�b�[QA���QdLJ5���
*�e1�QLB��(�)j�Q�A+QDa�*����\KX#\Lk(ŋQJ��jV�V�"��UAEE�*��EUX��Bڠ��b�Q`�����Y��b(���,1��m��Ub(+��cg�}���Kɬ�+i�wT�\�'��m�sF�vg���ª��
��.,��-S�nۮ'ܦ��L�U�N�86�w5�֜Un�姞�Y�v���F�Y����dƺ���lZ��&1ѥ���8��cv�yǡ;/��-�����`��-�ny1��S�S!<�u���uq��+�.����#4pv�vx�σ��7[���mmS&�w$�t\�g����wQ�Nxv�]��0lN��Snx��X���M��:�� �s�����.(L��"X�nq]�tBGm��Pc(��St��Tq�6��O0sӸ9PEM����@�y��.An�m���Cp^������v۔��l=��J�2�'�8���;�$�W'a8y5ս��k�d�������l�`��݀��n��X���c���%A������gי�+XǺ�e�<m��fM�8�H�m��F����&��ٰ=�bn�:�dpk������Oy�ݧns���t���g@-�f2�Q�;9D�m�m��k�7;����jCZ��9ݛq�ڶ{ul���x6��t�)�rE�Nu�[���Zۮ�m�u�^�v�x:WJ�m��v�]���Vi�`E:�x��:����|.�[���'�,�v�z����+��2v���\3v���h��ʥ��R�9�k�l\�֭s�q���;Fۣi+���ۍ5qM��ȦڢHP;v;l�k��8\@&���I"y�q�����n�Yx�z;sÅ�]�!�^2�`n�=��&خw�A�^����;�ŷ������v�;<x|8ѹ��s����{hg��g�]��׏\gn6|���U����Ѯ�;�D���ҽ����8����k�Ƅ���l[��ܯ�n�Ta�ƞcnA�!��kt�!�������>�GC:H(+߹����X���Z��뭤-�����`��9�9�m:�/\��㎌�Z�l3�i�� �٬��gI�}��	��u�i6�IXQ�a��P�AIЅ`?s�i�l���G��^|^xz�\��"����]Ĥ�D���'��H6D���;֝�+X*O3�u�����h ������$�^s�i��V���˫��5z�i;B�s����6 �m����h��A@�X|�Z`l��H[Ns���}Q�ݞ_�j��j$��]s.^��WY�
t2_~�Zf�++%B���<�bM�u��{޻%H,;��n$�B�J���Zd�ʐP(�>�0�M�;�U:r�����aM˹��`�$����n�U%=����Kfc�/�?���H)�`=�޴�R
X�R��i�������ޤ����Cԕ
$�X�����aXY{�?t��ֺ��u��o �&�VM��{�5��}��v�7����A�H!��b�E��6�8�;=��73�NYs�+������g�y���uy;a�y����@�V�;֒cR
s��7�Ak�]}���ˤ/@Wv�8� "/�1��X沽�w.k�i�++%B�����i6�R{z��>��k7�>H)<��z֒
AH)�s	��`Byw	)()B��}+��5|f��AHwl�sZv��`T��s�I�d���<��o�{��T��C�%B���z���5�����.f�ä���`{�%ed�+y�h���ߧZ�]�lJ�{��q� �>��t�с[��sP� ��=�]��X��(�*��ѐ��YX��+��`�L*��(���~��ٕ�WY����L��R
%O|� �T���n$�B����N�0u�i�`��FT
�:�M���=曋�k2�����s�C�B�C}}���^}�=��޵����;��I������y�Cht$�T����yίp����a�°z�>���ַ$�!S��bd���;�:�J�R�5�Ͼ��ބ�E�]�V��)Q���J���;G�&9?j�{�}�����=ɏp��:n*�/t�:J�	����H��@i �`V�9���:H)��|q�X治���3^k־��No��O���D�;��6�i�V�ϵ��
��X�ޱ�����Υd�T���0z�|O�]�HJ	I�|�>����ZB����;`W��������$�{�4�Y�%a�9�ChuT,IP�g7�a��}}u3s��=�Kv�i&yd{{]�@�@�#���3��Yh���J_|��H,������:gI�`r�z���������ﴇ���0�[�s�j'Q���̹]�uu�N�>�y�f�J��P�z�>�{ӷ�i3��&Щ+
°��{�m ��
�A9�ޱ �m�\���;�?0�"��y��>*��b$���^cXg<惧��-!K`y|ޱ���`T�L��y�s�6� VQ��������$�������tLAB�G�#�R���D�8�8
�R7ϵ�z� �)�{��m`XԂ���o��j����O}�x�q��s�z�;<U��oe+h�e�mEUOF�f�:b<�Gk�|%3��.�I�����D�r��K�&f��$m��RT��a��C~��}��I��V5�7�
Ad�'y����eH(J�}�L���5�}��=~V�E#�F&&ԍ:�$�Q���kn��������Q�kX�L5�}δIi
[���
AM�T���4�Y�vw{�z�:�M�bu�:�:C�IP�*a���������Yuu����;H)y�L����fyקy��דs[掆t�D�+����� �-�9�{��w�:�v��5�v��
��]߮cѧWY�
t����bAf�J�IS�y�ěB�����<9Ö��=I�%B�>��XɶVJʁR���p�>�zX�%%3dx����
õ�wϻ�5�ZB�����bAw ��s �m��VT���P��ןt��v��}'�z$�XÙ��Ă�w�����ѭgP�AO����%ed�)���D[v[k�"��>��A�m�
5 ��{�nn�Z0+D9�ܼ,� !i�����J ��yX�Ev}�E��@��u� �������'����r��Yguy�>'�O"���uQq����!b�;n��WY#�bf�ɰt��]�����;-���	ک#qi^�?f��{��i�\k�<�oc
b���g���u;Wa�\�����b��ӻ/���N%`�:�qv^�n��p�q�Em���
�ݜ�S�CI>��V���
�GGB�(�A��ō[��1���{���%e*%O>�ěH)�9�u��:�y�|�gZ�=`s�ުAH)7��O"m�L�}uu��F���X_��Ci!�9��p5��U��`T�/���<	�x��G���R�ȇ�'x�2��L(S2��1�J$��A�'��!��f�!� ��������*�npێp��3쪵 {��u�a���@���u��MD�{O/0����ࢾD�}TA�#�K� ҙ�17(@���8�`4vz�����x4nV��$����9Z�.!��uݪ�'��:�����2���Ф�p�0�Љwh�8�h�k��6z~w��I�,�{p�o��;{�e��z.�c#lk��F�桱b�Y��� ,�,`s�|E\��II�7�P�)AL���THnD�2}swڢ%����:��17�k8XB�{s3��\\k7�֟�%䢁 |ϒWv�	�Kx��xꈡ�{��| ���;��k>{�U�A/e}ͯ#gz�F֙���s�%ܝO�㚧�����:��l�I~#C�Y��j*ͮ�����pP]ݨoh�q]o�Z�j��1Jf����ev�=��Њ>|��{o�FI�U�բ�*�m���m|I��/S�}j�Ot*������/N�,`���薍~�{���wߔoz2����]]�꺭숃ѩ�I҅#wg�AV���NEcݷ��� �p��6���ۚ�O�6�Js�T)�HX-���k��T�5���b@�=�8-�]���x�2��X�z��8x5�z��c����`J��'���d*�}8Q��K�k{T��r��u|��p�F�I�����Pqoh�����zf����^|�i��}�\�a�>� �A�E%R�]E���@�y
g�� ��76D/�۽�&߃J�U���9����s-&��P$p���R�H���3���eO�״�4�.�MFt�8����M^���+؂s�K�����-37�b�p��3��]W٭H9F�:G}2�7\�(+v9���Ȁ�g����>b�Z籬��� 9j�z�_�|t㟰k]=�k����`s��'������	��s_i���pCe���l�O��s�a����Z�B�^np�X2��;&�x����H}�^�s�W�ȹ�����u�"�X"�T�w��`��mk���|�gmP��Q��O
	L�r�1y��]hQ#�� �u���� �U�7L�"`��Ml���8ܺ��Wp�st��e
�9��'�o9�US��n7y|���tz���I�qR�1��N)���E�{��T܃���O7F05��q]v�e����h��Y⓱)]O&{!۵�;5.��Bg����.4o=���n�=q:ݸD
����7%g�rhj�c]�qP�v�clY��wo+��ä|��nՎ݃��F!��:l:��ηb�d��{]��c]��u�X�Z�O#�Z<ݍ����Yy�l�w�a�J��z���w��%�2��>ϭ$(���!J��%3	�c���ٴ��w�����iD��7n��׈�G��$�V������D|Iиv�:���$��+Ē�
����n�%���U�n
 .n�w{|�����@3���W�$7�U�r��QDې����}�k=��]v̬��Ń�j}TT�
 ��	���RG7���V��J��&��m���y��=��Z�Z�>�֬�L��e����/�R~��}&]#e��_w���'�S}w��x'37�=�����Ӎ�C"��˛ڢA0�2^�b����O�pID�B������P&���b�NA����I�Q��EB�^np���]Þ�X�� ���h7jw��l�oR�y�)L�\��o!Cx�=�����HnQ^=�zmw�<��1��]ѐg�H�e�8����;�;�I��M����B"��P�*���`#�����ׇϲ���]zK2bS&�ft�g��]׹�gv�mY�6���u7b��ˢ��N��]݈>7]�#_�����_ײ����_E��!^���,�j{*���yG_������''�_�U�qj�&��s�]�:��!����;�hʎ��;'I˸�^�WBIm�Χ��o��� �"�<f�)�ݛ��0�8gU�� �H��h�g`D�3�������3�V�i��<�9_GW���9������WM���y9�M�ܘ9ۚ2�Ysݴ9��y�^?�J<��ŏ��t(xS��^��R�_��T��g����X��MtV��4��<�l���bf0�ҡD�"Q�pFU�v�΋�Ÿ������U:����=P9s˵?lF�f]���N�׭�w:�$��#t��ˌ�Q�T���y�^P:�mw�t�@��z�ѵ��d��-Em�H3Z��ֵ{w_B������u�i���n�s��t���*Vt�S�AxY�$;�wv���!`�:|gd�[�S�������x�����Sg���た{���O7s���;�kK��X��y<NY�Of��B��Blh y����=��j��=׬,�;���շ�{8�Yu|/�w̓{�m��OO��*�wJ����QP�X�EQ�E"Ȋ �EET`�EDUX�1��J��+��U��-
���X��X�bVA�pQEA���E2�QE`��9h�V�UEH�E�b"�H�Y[TcmEDAQAX�1E��A����TUV"1Q�DTTFF(�G)V"**��F+
�EQb�b���*�8�EF"��DEQ`��*2�PUEKaQ�0X�DJ�
#ATX�U��*�QEAQ�"�b1dU��A�#IZ.yלD�}����ۡ�{�4$�a!V���P_:j�	f*����tϽF���K���9#�w
Es�x�-��Fu��Ձ�����L����e����Ž�G9wЪ����n݃���<�N��[q�Tc��O,��I)�+y����~�g��m˻u�}��IUc� nsW�4��+��b@�d�>@���8���۾�+{�&!2n"4�$=h"H.�+\�Pu{x	 ۊ+��jK� ����۾Q�����gx�(�A/5Ov:�U3ޮ��7v�S&�KdA��4��i3�x��/U��s)�:lj���(�^�r��f��BQ"�;^�3�۾�����.8�36P$��Hv��`��{5��Qs}M:XKkQ�j�X��4� ��ac��G@@")i���
Cnp�&�%	w΃�X��Ο#�����&!BQVs�����vz"��I϶�CJ1�����I��E%R�T������S���2lZp�ޟ'|���fLB
d��Δ�7+hW�[A�[�Ksg�h�Y1X	/\�梼�Bff�u.� �Y�p���w����_=^���^;��G{s��H�Ю'y���{�;���_]��)�F��6N:Xd�w����<.��nl��|w�'QB`��qn�w��cvc���F�îNr��m�x����wV���ASv�wFN:�쭮F�0��c���v{v�tj�i�oi[��0�����(z�w)���Fv�r�j��I���c�⎻1:�+78�m������n�yθķm����wk�/l�J�
�]��w�Ճ+�Ns�Fv���C�2A�>�;n�t�"�J!@��F�o�GRӷ�I�f:���p�q���כ�����㑷va�� ��YD�H<���.�������ݮ\���K]V�tݮ�#2l�I�ufd��5F�P,ɈAL���8��[�����kj�݋(�H:�Vؗ�;za�,��)c��[{���nn.�Zl����� k���ĨN�s灇��0��Htx�`��u��+�V�I��R*�7(��s��dp��0E��ˎ�gl���g��F����t�0x?�XY�Fp��}8r�0�6yw�@�|�l��Km !��X�Y��6�6*P���ϰ���H}��ln���^'Ğ漊�ɈJQ��=/vn�T�Q$���S��/��$d��PJf��(ok6s'�������>�{e��u���"㪪U�;����q�����j$��T�b~u�"׬����{�Esu@+6.cdI�7L��D�_l�{�(�����.��ʳ�t��vA ��^^��B�e���M&���n0B
d�f;�#����O-����]Sc�ay��e�8�q����{N���ݿ�.O�s���~	�,-�Y����H�76D�v�>�[�u������\�f�{3w9��H��K��@�[�'�lړ�}��J�|����g1�7��d��i��Q>-��y7V2��ϫ�U�۷e�C=Z�,,Q���5,���6�|�ER�M�D#��ZV A�X,u�v	��E�uEwP.`D �MX��(lT{P���#�9
�(q7;�-��������͙k�|y�A�k�Ҵ';�K����V��u�x�R���>�k^zb�ܵ`Ǆ����؋B4��!ݮ��3�yo��$�٬2��b��G�!>�L��\vt)�b�������J�B�A��G��s0�E;j�R��#2p�Hm���8B�p�|���iDd�AGjPq��+v�j#C���cvR��j=^���x@�ڈw~�/��Y|��������UZ6J�+q��OEx�>E�A4�0��O���t_*��g��_��������C�1�}���S�����ٸ����#DN,�X�$Z�^<��'Nj�i���4S�:�;X-��xC@����8��ӛ�z+��_rH�Ψ�(�3+��x�LuQ��5�+|OK�Ol>��wyC�l��k��}a`�%��]�i��+��e���Hߖ��uF�쫀�[=��\������ݣ�8��7�'���ܞN��Tqt'f�]�z��Z�<ݛ��3e�gl�e�����s��ݷi���h�t�t����ͧ=��=�km�y��]c%������g�]��Z�<��<ƻw�m���9�)��.6,:2�rȤ"����@rUJo==\�	D(_N�w�Ew5@�;G���2:��!�fԙ�|�T�������/��q�H����}�\�~��9E�=�Q��*r��J��V B��z�������d�/}��M���QGG9U]>v�b��s3�^� ����[��t{�V�z�
U@���:��A�}8X�ݒ3M�(�F��� �v����|�b����T)F}���A�}=�wo����g�̩���~�?(������s��I�y�C���ܼ�a�����q�R�	��x���o���������T��W��OQ>���&l�b�=݃�)�/*�md������<L����5��2;��$��� �(����7Yo:��y�RDݭ{��Ўc�D,�vX]9n0����D�!�Q��JT�-uE�0��{�`ׄ���)>=<�U:B�k&�I���(�Fs^K��m��rp�I'[K0h��97��mi>�m��Q��BU�KO�#���|@�uK9����h�eSw�&�}8���ʸ.fa��XD7���$\F�b�:��ܯ��K� ���ܺ7��m�()ELqd2K�ADV�]7u��n"if���51*w���ƞ��g]9�<&�GX���h]�5�l�A���y#���nŞ�%���2�1C�⪣���`$��(�A�r"��,�m��3�Hq�;�FߐENR�\������ƊŦ^��Δ}v�ʷ�Qک��wO߇9K��=���/X�d��j����cq����o9Պ�`�ODF��9�/\����;�(�v�N�]�Q��Y^�v|X�%W7^�|� �s�$�bB�s�6ȉ��1(L��i�ב �ϹQ �'c�c�J(>��D|_�e��2�E*��|����$�ԉn�s�6�[>�Q�?p�4rrg��WKړ�r�.7����a�>��<��΁�v�+55\�A�'�S<��DNp�oe�9�l��Dc�ر�s����(��O�k{�z]����w��I~g�&�ګ�?��mև�Z��,(�f���? �9J�V��=�����q�k��d���ws��{uq6��*�1���sdR'H�4��n�GC��9������|��B�nS�+&ݠ�����^c�7�_=TI�����BPHP-��kv�"	�����	-�:�MKso�뜻
����BSW���s+�g�<���aN$A�ۏ#���c����`~���T��V�*���!Cw�I�?��Ig��B����O��K3
�w)���Z0���6�nӻG�, B�T,�$��>g���K%������!f��=���O���������~s9��Kà��f��Fi�a;����o�Ǔ����$tz���}��� B������������@
I�I$�$�ɐ����A'�!B�a�B,,�I��{�p�:�?�&��d�?��u�|��3������)���B������R{�g_�2d!���S��}	�>�����ֲ[�����d��������Y���'���) B�ޟP�7�����;��OP�B��t�͒�]�/̗3�tt�h����z>?А!C��t�����'럙�����	���,�2~?����=?,$����� ���������ͧ?h2�!�+�~����u��?�~���6e�'��g��Y�'������?I����{�I�������I�������𝟬�0�B�~�1��?i���~�y��������?$�!��Ȑ!C���?�?c��a��,��	�O�/�A�3��aI�ܟ�u�d!!C����Tc�2`����xO��HBc&�6v2O�D�6Mx{��,O�z nzL����`��?ǳF��
��!z`O����$����@�!�� �2��������?������O�����	������O���~�?N	�x�|?�@����?��?����Ρ�?C��_��_�$?������?l��������O�<��?�<�	��	���7��$pO쟻F!������r~����_���_�����'t�y�~���5�!�������������C��]ʟ������3�ۻ��f�D�?�7$�?$�!B��a?�?��~��������~���!П��a�t�S��):���,�	7�Y�.���	�`��I���������)��;�@