BZh91AY&SY��T߀`qg�����*?���b _     �                                    @  ;�ع�   T  �   -`   &�       �@       �      7�J�
��
���) ��@(�TT��
$(�JRR�T�AEE�BBU
DQU	PP C�DH�RTJ�D���J)JJ�y�I͒�����:�NF�U�I)W 3���PI������������I��   ���R�*��� �  k�*�� �� w`9wp�w` q�D)���@��v ;�=�  	  �a��*|
$�QU��*�| a�� �`{� �w� 9{��)p -�/@���7{�y@ �z�k=�@u P ;|��(E�� /G�` ��x���z�r�0�v��ף� wzAJ� mc���`�y�� 9�y :    ��� j�@�RH�(�)Aww*H� l||� 9�z�^G{ ��{���C��ްx�� �������N ��k��`x   (�� >�>@��  s��T��N�t� ��F�{��@ �{���C�`�;��A�    w|�(�(� �*� �"� �<��@7`�f � �X -� v� ���.�H�� �Ѐ � w� ��{ >A� �U� 6��vE2	� f�"�pv9 ��ħ �     8�� zU"�(��B@�@x���e� ��� �$�������D��� 9n�*� ��A�0  �J@���<���:
n���v���t��(��@;�9@d2>�     ���)T� �    ��bJJ�  h     "~�U)3D� 2h     y"i�*F�& #M4�CFL#A)�J��14�`&&&�  ���2jmQ4ѥ<&�S�Oj�xP���i�a'�������~��O?V�����~���O�����>~o�O||����J����t��]���T����IR�g���W�/��������?��{G�/��JU��]m����J��_k��ٔ*U�������0~�WmW�j���W�1ƫ���8�q��W8��'�48��.��`�C�G8��C��28��C�\d̎5\iq�ƫ��1q��K��358��+�L�2���+�`�+�W`�C�v�ƫ���W\eq��UƓ�W\l��+�W�2��q��K��2����Uq��Ɨ\iq�Ɨ\eq��:a�GN�dq�Ƈ8��GL8��+��8�q�ƣ�G8��G:j8��C�j��q�Ƨl�2�4hq�ƇWY��5H�R��q�S�*8�N4QƕiT�J.5$�8ԫ�K�J8�N�ƥeQƊ�d��JN0G���锎1#�Dq�N5�T8�G��T�5ƪ:b�4I�*;j#�R8�GTq��5(�P�j��J�j�5Rq�'T�8�e#� �"8�b��%q�.�N5Ut����WAƕ\d��R�Ȯ2U��(8ԗmUƀ�\h��%q�8ԫ�
�D8�0���q��5Uq���8��+�W\eq���2��q��Glq��U�5\eq���2���W\a�.0t��K�.2���\b�UƗ�b�f8�Ƨ\d��n��������������m>�Rf���vƛA���ŕ��'��t>��	���;F�)z��'%��wq~]�z'�Ç,لom��#~Ց��0-K������Wr7|�6�{�m�@z��E�v�9��t�ǩ�b�&V!��]�yt���l蠶l��#��v}�WbZrc�J�B��=��o��̎��Q��F�Vk������
aU�8W&�¥�TX��2)Ga��{��M����qYz�O[�`,� ���]Ĳ�'n*fu8֭�����^ӝ�n��/�e|��V9i��ʩ�����B޷��7]��yK2+;wsb��{Yd�xw�Z�1�UZ�gwRŖ�-��ŕ
ƌ�'�Bݓ�A�_�@����v��;;5lw7�μߍ*�4��bԟd5�mg���*�;��x�<Ha��� �tըv�����r�n�r[��ܔ��
����,{<��'Bʋ����_�\� d�*n��^�����r��F����:�����'P���z��wq!�|Y��6��Vn��㈌]�!���7�t��:�X�;DYǶ9�8vW�a'����,ǯ;1�fZ�������G�Gv�����jq &�y&\�fL|^�δp�� n�._s�ɀ�9϶r���ť�<3��&��i�j��uqf�K	=���@���6 �� ��|�g;>�m��j���g��c��tn�q��r%��vf��pm0N'vj�رn�$�=�8c�&��s��{���8�b��u.�+��S.���Eg.4��nL�2ň���bS8�8�6���dð.��ǤJ6�2ov��Ϛ�{N��IkX��nU�/c7:�V�"�ڞ��-�}gH9�ag����r�M��`Ʈ���yغ��{ANWٛ ��	��M��|ť B7'(Yz�)^lۗM��v[��+q��t��7|X�	�q?q�}��gT�9��	]��a�6ܒ�{���n�2 ��Q"[���=}�����-�]<W�n뽰\}T�x��Y�c�cg��n�gv�ayu�wV����8;�q�,�*��w��u�=���3��-�+����Oȇg۽����8ǹ�G�%8���X�z����O�Ż�%s�ܸ�F�ͣ�j��FS�r�oeŊv�p�[��r��F���^oF��҇4L�O��Y�P;�}��Q���^̓�Ʀ�qc�v�f�M�3�E�uC;5`�������&��V���0�k���C=:����F�eZ;'u�:2�� ЄԘ8�[��<w����cB,*,�g���F�)��rf�	jPظ�U��������n�E����͝���ǆib��/mw&vnv�5\9�E�b�:m������[ ˔���/�L�	wz���{�jf��=�;r���f����rI���k�Z�f�˗I7ȍ梚:榙Y���ȯ�6�x���Nŷ� ������F�b�J'�n�;�{���xi�\uף�i��չp%�j�o=�+u��q�qhȲ��4h�Қ� ��k��ȃߟ�2	G�sx���I>�F�f�Έ�ۼ�ޜ	)\�Ը�x;�7b�f���p�~��������]&,���uk�v5���Y5�IPd�q�V�;�t����!z6	�)D��l���t����Gvj��<ܨQF���ǻi�m���d{6e�|eõ�9�L��vk�ٍ�n�uf���'�P�V�k79#��'����<ܽ�NYw,�Ն�!_|���A|$4����V��������-W:k��'��`ف���&����68q"���V�5s�CcI��a\��F�t�Zқ�˽��9��\=֣ϣX7��K.�K�,u�FAT�yoGswK�'s{�ۊ44�ewj�J꒰{���jï�Yd:��dGZ��\�qgB���
�l��1Üyww=Ⱥ����ުW��TsVt�%�U,G��Yۛ�M,�2�|geZ��͘�JD��o8��8��V�𑄠�h��{�s�23��	�I�uH_#~�wC�JN���v��j�����{V$�]*� ���rt����>큁N��wz,�fAb.����;9��8��nr�]Kеt�Q���dt�����li�h�d�nգ�d�	��ôl��+��Yש���Y��A�s]��M��w��d�H�@��r>*����xi�������ݧbB%�g���[���K�l�g�Zqa���`�w�=�NF�{���َN�W�tB~</RYYL�K�&v��X\f+{Y��ަk�z�i�^�q2u ����駴Tk'&KtNR$�d]�wN|�c��Ѻ0B4�SX}����Y��>��Rc��v� � "����˦��ۅc�H�b��Wq��ɧ�#��i8GwN�zބ�@B��,�s���v��9��D�*`�l��(�Tۘ���6����&H�nuVc�<Ļ��n�~�Ӌp=�:�ɣ�ڦ]�0�+Ǉc��8��8��y�o8���K�.R�Wy���2m��ւW�;M=��"�ݦ�b�O��&�ׁUD�g%7��Ym�PKwc;[�¤y�w9d8��ܼ�;��t�2;n{<�`�vj�ښ����N4ecw�*N�<�W7��ҳE�ٽ�tgg2-k����'>\��	�5��淥"2���ہ�����:i��T�pup�z$<��P�;�|�MF�e���6(�p�$nn6�ʯ7��;�����]��;���g�Yk����n/�2�,��E�z�q�9��w%����g�C���>n���\��U�ǜ�R�ی[:�����0�͂��V�tƳB;̆�	��T�wp'��`Y1)C}ۥ�QGѮ�XΠ�"��х˰W�)%�ݶ��[�Ö�}�	;�0g �����W>��?�w����3���ŤH�v�;%ym�eP�D͕f��5�E�ܖ��Ky�rr�a�|eWips�0��̀�Y2d�6`�td�M���l]����]9�ZƋ2d��ŋ���vp�~�V�;�ܸ��Uf�\|/p�$�V���ܷ��#jű)�Ug�Y��}��mĿ�IvG���t�$��y���=
�#��;�6�0�Ռ]���!O&����<�H����^I��-=��������}c�e���z�V�`��	�q���W ��ޑÜ��t4~7A�9��_9Q��~%�S���F����㛯iS]�i��˴��)<���K��:z��k�
N�����`�s���8��-Mn�%q�V�-
���qe=v��������9EnPB��&���Q�B�kJ��%_u�_9�Q*(����r���7�l��*���7;X&������Or*��&��>��V ��\�g-+��_1��}�w�^/4�#y66 �ĘNM}���yG7�N�b�A���
�5� s�"��uɕ���X������I�83j��6���*]�M��{����/p|q۱��]k��N��;8$��f�V���\��mHH�͵���qxJ��sjo�m��U]� ���{���-�i9-ݕ���:3��:�b���M_\�o&� ��D˘wt�Wa�'\�[ �h@���x7�8�Y�P���a&��sA9ƃ�kV�2�e�up�ww�q�Fv���*�ro%s{8nn���?MGw�{[osl�)X���]�w1��uw�����R�-��1�Ⱥ�-T���;F$:�X�9ٔ]j��s�t|Vϟ.�)ӂs����_>���L6�C[I��Em�]�;�Vqt�+�fv��R�uZAZ�.۷+�"Qa\2����w"(Ow���oL�{,����f;'@��1l�V@�4��&3N]ٰ��t<�[<팔��pKKӯL�t��9�8�X3�(@�f]/r�#qG�7��������&�(.�ӱZқ��c�d�;�;*����9�r��XGr(t�7T;���0Օn�d��@r���%����Q���ǢaӤ��{��L�fA�H86t�xn��#�L�R�V�r5.�T<�6�øB�lx�ޮ���Y�.DY4C�ǻ,���h�og;�����b�\O=�ꟗ�>38Q�ʣ�ろ'{�vǋ�r����7;l��M�{:wY����d�`y{r���sO�H��"�m	#��"�n6���X	��K��8�퇪�����5a�yC���t�D�S<(f�u0Y[ɞN�.ӫ��i���9�i馡r'����m	`�Y<�姆�x`ù9����r�k}!���&���'!s�,��\��{.*7�ڕ	�T�6��Y�T�"�V�݄�n{Eܩ�݁p#&@!+pY�hA/�*�Yu|�d���;����E��Q��c�v�ٶ��)ܶBh���+�Y�.v�Uv-}�s~ם��p��F���L�2%^kN�`/+��c��p�i�2��H�7�;I�>o�U�\�Y�d3Qwx�^9��˳���Y�4�97Z�vӱ9�{��� ˗n-�i�n����r�ω:��V� ���"N��at|uv�]��gz�{�	K�zs~c�Y�"�+E�2����T�;:m�����S<�t�ᇹ��cX3�,��f�J�w��;ȑ|c��Ɠ �_j®�a�\-nQDG�mc�Hm�Mc��9�n��l�\�A{�5,u�����F�&�8yţ�+�6n�W���r���]y����\�z�㽜X<R��G��������\��P ���Taǚ��>h��F��I�����
1���>��w�Y�/#�I�gE��5NG֫q\m�P���05�`�ٽ�#	�p�vR�WjX�l�#DPO��w�KA8�3�=�H겐������\�9bb�Q^t�ŉ���;x����U�B���sc<�]p�{`"�Ȑ�jY�ٮur��3{�(�0�V�B�l��\��5�E�;5�@뽼��*�jֵv�eK�;rgs����LB���w+V���kX�87�Y��Tzd������Z�������<\Ψ�&�M�۸���&�e\B,�%eGypw��;V��6s;j���4=�4s\���W�W ��ɰbћ���e\�>��G�]�l�YfN����J�n̑iX3�aS�᭡�u�@��+*�S�A��8���)����{Au�����$�@孧q�XqS-�.`/���|�R�yvs�w(�;�!�x�x�=�=�9��M.M
�'hb�J�4���Or�����i��3��4t��P��"�Ӭ&�v��x֤9!��b�G;�d=�ool��S���M���T �p�*e���pt�9���#4�U�.�g	�T<9eƴ���8��.��R�{%�C��]��BD�H�y�)�p^/�b㹨f%��Ӌ*�N��M��J,M7�1�qg*�j5�[p9�X�����W�#{VD��݋F��رN�׳m�a!�Q���"pR�^G�l���d�5�H�/��@�-m��8�z`��W��	�y��'U��m3ARonQ�����5N��m���J�{.�8��v�U��y��OF��˔pj�n3�Jc�y�5��n��L�W[_}4�c�	6��:5��q�e�3�J�I�����S��v�㧦n�q�*0WeǱ\$f�KݺN:p,y�Գt
np���<�KF-��bՖ���s�4�i��H�̈́����D0R��>�A�p��8s��"-u���^�q�h�)1v�ILC�7,�l啍8�i�D�7D�y���f�yԌP*G5�1�6�[!'�eǓ9&����Vla&qc��L�k�ū�wAO^X��>p^zBi:>�,�¸� 3{�8n���wE�z�����j�]M^Y���4�!�����(�������ޜ�܋�T׺�� 4�.[���T6����H�K����B\ak�E�f�>o�(g
���x>믕���oV�ؤ����u�Ć�=�P�	�˞ɺ�4�9Ҷi<ҕ���ah�t�6\����{�pTQjɶn�/c�#�Y��T�$�U���0h�ós��w��J5��^��w8���C\+��gK�f��s�@�z1n���O�P����w�S��g077++L����E��\8pZ�Lt�F�%%����8;HewbÎ��uT]R&I-����mO^��	�e!W{{�Z���睊��͚��yCud�;���qI�s���4qt޽lm�2����ǶU2�g'��I�6�󆬌n��[d�"u�{�i,�5h2b9'f��!�P&����ߒW4^�
�@{L竱�a�-�d�}^U�^q���7�i�@s��{[P`yv�bݯ6ţU;4�)C�-�p�b�4L8z���J�2z��
�PB���#ٛ;$�	�It1�nѸX�X�{��/���9�y�����c�<sy-�35�"��_�a�l������2䜡p�nE/O��X,8�5�}�g�s�ܷ+;��26��lոNw;V4�QF�p�u��7րo�h�vpf��a���盾��Q�Ai5�y.�Z"9��R��1x�9�f�;P���q��h��ɨ$��E���y��g��B�.o�2.���e��P>f��}�x]Ah8��B7��D��5�`��t�Lsago.3Aײ��<" ���69���������>>����O�����T�2��[UD���������-�l�m	�T��M�6��&�ڨ�(�[*� ؍�[(����#dʍ�T�ڥ��ڕ�+dM�6R[D�%m#e-�&�(ڶ�mFғdF�m6���ڥ[l�lبڪ�+j���6I�Il�j�m&�[R��l��CiPڕ�����b�Rm�#e[*lإ�+`أiM��ڦ�Q�6���V�iSd��څl%�-�m+iFԩl��U�#h6�� ̪��6R}����\��>>�s��~7���L��lS_�:��?5�M��M[t";/���ޟ^�B���X�X[cml��~>y����o�|폂n����e�<��+E�����:�w�8w�;oK���
���wYO5`�Z��F�bŅ���[��g枻���}h�5�e��D�maϲO	���Ma���j?����2����H�6q�3��f�&�C}�����7wͳ����w�>'|������R����� ���_w�¿���������+��������S��w������?-�� ��C�ϊ"��]��|�����øy-���Sc����ɛ���W���ċ&��j
uV<�e�:]ٽң�����/V�������=�69������ ��>�\���&�>���� �ծ ot]ϻR[������@���F�ys}�i�n �g�{�I���J߼���;��S8�~'zpg�κ��V�h�θ�������&�^��������bzo��gjZ>�_���g=������������{�QD䈽�Ѝ����e|�G��>�wyp3F[F��x��'7I$*o����O�w�Β.;����^窽4��WIG��\������
tG�_/,#��c� ����yU�������2g������Vo��5�/�]�,U�o��e��x���cX�{sx73��j��4a?d�Q�[�"�,���;66���h��;��1l���=����.����}���R�YY_��M��ֽ�ۅv� s�NPs�y��&������:�����E<���x�4�����ð��3WAq;��98���h{7r�i���wm�^���{��}%�ܚ��έ��yYZ]&N5�W.���mŤ����GF3q���ՌysP�� d�S�xo�ӳ�Y��b�#(���.�\����t���[,�g�&j�.l��|�9E�eC8�BĆ0P����`��0`���0`A��`��0`���0`�0`�ُX��6����9��my�$b$Wׂ�>��ӞM��;��gz�z:�������@{��N��x[��Xxb�J�v��ѓ��������POY�V�����r>9��.bY�5�)��к_E琟.�W�����g��4�ӣ�f�%��4�ż��#Ci�w�����[8ў��OS�ڄ�s�[P�q�F��nM��t��h�y{-+�w{���'����9x��{L3�xkQ�����~!wޝ��z���K;�}3�ˢ�q�LՍ��Sɞ�.�H�WcC��Q��ص��55�1��^�e�o��rp��܄c�������O#����{�̠=��ヲs���#%�z/�$���;n���&��)�K�N�U�y{1��Y4FfG�s���]���Vͮ�o��O'�����trOv�׍7X
����έx������C%��^<U9�xc�2�%e�l�Ȣ��,Ձ����QG�8W���}�/�����)#�<:��'�(�F�n2F������L7��!T��~ ��6����c���\{i0�0��@'������=��\rɧv���m��}�s,��IE��G�n��d�û�E|ۆx��ܯ�&��M�������7M��;�L���=����ݫ#Z�=A���q\빠nrؽ�OV
��v�G�g��Ȁ�C�p���VD;\ɫ�,,H��@��0`��`��0`��`��8p�0`�`��0P���0{=����;Wz��~���X����Y�����\������ �v����N��[���f�ݭ0�L�f����\���"�l�H��=�ۂ?f�1v��*r�(�^FS��z,�߻a�!����~ܪ׷�Qf��������<m޽�g]�\'{�^x��7�W�p�)h��)�	��ۏ4h�a��3�OI��w�#�}�r�0���9����#��.L0��?O�=�ޤ
}[�W��`�����������2���.��TDLe�8 |X���a��X�9��}�C��hi�}�<6{p등����w��r��7=���k�T����W�����x��v+��7�)g9��=�zL�}�g�g������z??H7�1OU�ݷᗼ0�7��u�G׽�R6	xo����r��_j�����f7@;�0[AT	����A�N��s<����"=�I�ƞ�YZ]˻���|$�<��N���ƘVMK�<�/3��J�s�֎�i�dTy��G��}W��1�Tu����Brb��������ע�ʱ�4���2&�����m���)��|�d\�h���'ԫ��6���	�u�{�4��8�>p�"����K#Ƨ7[�y��q+�bG*���}�&�X��{=wh����?+��{}7>�|nܙ{|Љ��l�����5��y�oHAǭ�w_��"�츺O<M�4V�u�}j��
i�<�r�0X��0`��0`��FON���q�ӌ����������zg��0`���3��n�ja
��~�7�Ͻ�{��7_ᛴ���<m�p���M��1�P���i磷,�#�Y:�h�`�'\N7г��,�v����w�@2k��gC�G��=u"��z���(8��Ap��wm�ϣ�g��� ���晋XT��3���"��E�N��2l��jȧ��fw����gL���7CTy�-�W��Eӽ��{���I�D�{p��]I{8��_C=�9k@�b�j��m^ƽ9�Do��7J��<��Y�[�j�0�=~�Z��@7#/�(�i_Y�����T���KVu]/�t��#��38��yT�3����y���1��Ǚ�_K����K�ҏg�q:H���C]�Ye;�A�.�h�(�<n�%��7�F�D{�.�-V{�ɟq�=��o�V�(�螄��r�i^��:���:��g`����Sk|�n�	���7���z������kG�2 y���I�������q����}�'�Usx��:r_Lյ��#ا�PhF��l��V�8�c�Է׽us�5��~�����{ǎ6u�||��$�/�<n�C���;���I���Q�ӄx��'3���DC��l� "����C��`�f8$�^,{��L^�����^%��^P|g,����rN�Ksχ@��p�Ȗ��+�n*�>��GI��� ���� [�tG̯Q]����P����n�J��J��^�w��(`��	0`C0`�#`��8�������������鞞�������/C`�����$�=b�lƊI���ב�l�ut�j��N�o���P��#�{�M��x�ǸL4�s��h'v�a����k�7㳕�ˇ:��=!��[ͷ�>��U$�fx�����e^��Ѻ��#�P�]	v�>¸����qv�WeA�u�ٵy��S�Zό�6��F:�0�����{�o]f6Nܗ8��}<��2g�-�dJ�;v������j�1ц����=��X1_:W�q��ר|w���W5�1��8 $���p�y�27����s=�#���=s@{�oe�&f�q���#|D�A!��;��;�;@pK�+��KbV����;���El�S����w���-	�ӱ��v\����{Tծ�b�xF�����v%�8���*�����{vg��}��s۞?z#���n\\p�W���i�^{��=��I���x�9}��FX�\�F�ٳN��t��Ү��<��<;:�ʨ٥J8�{wc��7�����Y�v�n*�=��\�=�8��^���O���W��^FX*~�"�����ݠ���7�4uSӏv��/>~��n)]������q+��7�@���'r�ks(��>H�[_$�f�J��ɓ �M�&
2`�q|;�My���v���nӏ}��<�d}��YrA�I8O��x��`�������u3�����Mw���i�Ny����{�'���}��{ik��㣳�g��F6Gg�#��/�Cj��ue��u:�e�=r��5{uɖy/����з����ט�Ip/7h��8��g�F�2��u�5��U����e�XR%s�"D��7��S�g����;̙��~Բ��L�>|қL��;K�5{Ü�<�+��b��_}���j{�)��9���r�!�8}��S,q{���7�XQ����r��on����:R�z����6�x��ߏ����8+��ygf�ʛ��K4��M�4)L���<I��q�G�e��E�vypp�X�(��͎���a���?v{���ճ�U\��F����1AӜ$����<�V4+��)�༂��}�i���4ķ����w��7�;�<�swо�$��'����b����:o�KF�N���,��g_&'�<�a�>�꥓�{}�FJK��BI�ɕ�sֽ�}r>*y�s����Ǖ�y��s��M�c�����%-t��{�(K�~X%N����fy�KON�v2��>l/5�h��Ṧ{6#(���0nR��r d�y=}8'R��3��_��f��5�Az-��'���7l^G��/h"SsJ�;3VԦ�gn{��s�4=��O���ew��g���g�.Uv�w���9rޘ�-�n2s-�;�i��j�4>d͡�p4��7 �zw�V~y䶚��=,yt#�7����?��;�*�웥�o��y-��a�$�xq��^0{}�W��mm��3�/����˞V`�_��G�����M�*P2�j-�	���fø����[�{נ�daN���}�Ķs!"�q)s��˝^s������7Uķ	?#�2�Y�֯f����ۙ;�Ju�"ݎr�!�ݡ&�����W��(��j�Z�vo���u����p�E���N��ٹ�ܫ�,�{�o�z�>�/�ס<��wI�G�7;�ǳs9�û@��vQ$ j6�+����v���3)�Ǯ��7��O!_>A��K��\ \�����3�z�~h�
�v��Z�Nn�p����<q���2�(j�=���`չ�����.�Y.!�۸���EZԽ�ڍ����e�5����������-�E^��b~�{h0t)�:z�1�^c%��Vk�9����>Ƙr������܇����2���*���R�b򁧹S�FW���7���4Z�/*�V�O�:}��ĩ�G��e�e���;���=٬)���|�x�OO�ŵD$���z�Λ�{{tK��#/)}������h>ʀ!pk��K�x�*<��ס�� /����a�I��x.�3\���͒o��~�Xt�p\��{:Ͻ��γi��L�gc��w����Ӳ�8����T-ӵ����Y+�G�~�'{��0�~]����c�����w��qCH��Ox���R���c50sy�m���|:a�Z_z��c�'�6��΃���-���V��zG��@<<�xGN����\Y݋tu�}�-xq�wu��{.nx���x��q��f̕>��8w�K¾�(F��#Hy��fw��3�A��?5�n�,�j{b�^7��o]�B	����n�tϑ����t�uxo�;��=�)�Z��9k�Z���9}Z[���2=���j�kt�!{w�G8��ol��v��6��8+,t��3I�QY��ۣo�/��^�d�ty�S{P�w^�+�}�s���l���9��F; 4K̾�V,����I{Ե����{=�k�ܶ������x�=1!�<�e��NΛ��ah�}�G����&i�����ƃ�w�%��3=���tz���^�7}'���!۞�� 0{���r�o����ٜ|�^�](������d_S٥d��ݹ�]�Mp��z�e��e��|.s}�ں�� }{޷e��M{���\��c�Rǋ���EӜ���F_4���<c���<j�07�w�0/%<�����������=��@��˼}_qIW4��>oޝϽw�v�_v"�r���3�]�����s���j:��7z���㺧P��q�o���7w���dC��W�ޜ� ����	/��7<��cB��+^��Jy����o-�Z0w�>
{��5�����O�G�_e������(=�5���x��*y���k<6�}��p�h��6S� ԰�"�YB�,m!ĉl�c2�񲱳Ke�gK�wS���M�<���ڥz�؟u�@yn���/R�W{�͊�0�ɗ]��������=����5A��ۻ��3������R'��U}I[����1�}٩Ny�۵Bs�h(I��p����]��e���CyN(�K�G�d���Z�������p�T��퇄�__%��^� 88���@{�]�5���\��g��_��ʞTĜ>)�0g_>�3�{���&Hnx��+ڇ.�<=V>QG�v�j�i�B���"�~�&sN�7�Z�;�,|�"2�hGO��~�̸� �ɽ����7���3���@���s�{=�ˉG�/_/n����'Rfq�'�O�Nã�KX� ��ʶoYP�S$MZ}�׀�����t����ǒ*��l'�����i-���0�w=���k=�,Ӝ�=7}�go��l����T|�/�u�S�>����Oo�͋������|�U WF�&)�U���k��mt@Q�p�d��@ֲ,�&�'9i�oE�����u��� /G��q�<�Ǎ5ZV��=��ޗ=��;��P�<u�h t�toj��s���L�h��]�}�<���É����K<�xi�byu*ro���V��̛{���<����~��n�w��o�u� 1pw��8����9	o��ww��#�Ǐ���2�Ǧ�Ce��|�6����ly�6�j/=Q:7d�;�8��3ۖP�5a���sy#��f��ͶMO^n��зp�W������]�R�{|�}�֝���|/z�����=,W}�����|c^^띴�o>;zg�&7�!J� �>/�\�k��e��=��̭t���	J9���;���������Y��K��!�};�?�O�u惩0���8oU��`�_�TyW{��88gc������}s�~�w�s9�q���"��'*��������q��Y�,��4��H��q<�y��3e���"����BC����$�_G���of�q��<���A�"�ás>�F�����ns��I�s@^
��� �Ӿ�x}}V���5�xOH=�r1\`[1��\8�u���~��u����wbb��L�87sS��0�ygzv�
���-��'M�����S�M���Q2��A���������ĸ���3�Z��^xv-��˳˵z��s����q�l[s�G����������ǹ�!��{4\��q��{�\p_[����J��������🔪������ǿ���v�t<]������f�e�a�4[�W]��7��.|��W�I��uh�䲺�d�k�G����k7i[\�s��v-��{e	�Z;]���{=U"��v݌A�m-���da.+�e�HK�ޮ0=�y��;OL�9ص`T�m���p^t�Ȑ�b6�c��i��-n�J�:�֙�g��yc�Ye�Sr���3�g*��<<0{]�����,ts����W1�/H�i�J�mb�=���DΤ��!R�#-VRR7d���-`�+m�W�Z^%γej�%(�eֳ6�"^.䎭��V;-��.qmp�7=�遁��ˍ�]i�: 舖t0l{kG���͸�9�i��i�M0��f	��Ľ��U����1��v�2�B4�]�[#,���TƯd� 	�;m�IՓ���^k��s�G[wZ����m0=��\��K�5���u�RT(���vl]*���.��v��p1ܢ^z7Z��n��܆N� ��ڞ��"�{�^�I�̛iW��i�99��!�y�P����.� �5�E��V$����͒��N�9��v�;X�]�b�͸�]�5k;g�=�4n�*�a�ݕ`�j2ڰ8-qў�2�2�!lq����l�e޺����Bse67���׳�i��Ph�ѱ-�
Y�M�:��a�T;��a�WD�e�k�̚ص�̫�f��[h��th44lu"�M�M��V���D�W:�Mn9������n�뮉br6X1r7��í�;��zq�+�Vu{oG:���mE]��GHvE�gU[u�fM��9���ӹ�u�{�����W`��l��7�d�ۡN�^��ϝ�P6�X���7�Kaci��T�O�=�*�r7v��] m�d�����z�F���ke8i&C�K.�1a�c�ME����Z�X�#]nۧ)5����GY絧3���GQ����t'N���9b']�wud����=��{���wn�:(����YHՔ�z�½�D͵%u�������o=���n��,Q���ԫ1�`Hv����@���(�K]N+�#�6��ũe��g"n;A��l��%�>;q��k\�+[��|��s����p庮`Z�ܩ����6R��7b��ݛt�#�Of}�s��.�5�.vV�ޏ^ѳ�L�%]�@csx�[��jݺ��|��q�{.�Ftq�G K,H��d�`�*�i]/^�v����:ݩX:{]�����5���I��^52!&Ր��Fme�&@0�g�x_;��cvzwV��\6E��n��t�ْ��2�-���s�<�l�-um�����(]ͳ��\<�]�C�׉��\Z�\m6M�b�������S��-1-�޸сhrh[�B%�5�VyL�Jԛu�V�+r�h;M�i��Ҫ��F�&(�۱�]��u�-���;!��t�;-����M�kl�%�nL�/7Yc�WjT�
c.!A�Q�0�+/b�zl�3�,���n��ت�]���,P���\���Y����{n��z�s>��:]���\�m�HD^��\/��S�y�=����r�Q[˨�cq�e����N�q�g�*�9��g��x����(s�V�!	�f��D��q����Ǟ;�O<��s�û#M��Yd�S������\��d�̤�ݵ���Hg�zy����|b�|�c���7[�{�tvY�Zz���ڇn=m>#JNZ�d��nCȔ�m�I�nָr�.|�^㇮��9���[�v�2`�q�I�cA`�X�2qgև/iX؋R=����8��F��&��X���U��ZL3WG=�d�7j���3�ۍ[`�+�7\pN^d��s��B˲�6���ֺ���<����h�V֩�@�Wgbxb̨x4<uu<���p��X���0�e��ɞT�YZ�d{V�A����'���ۙ�Z���p�l�!<��9ms���;�M�n[c�4u��|�Ьjݘ�m0��3֬<�u��k�R;���.�Zha���FԵ�+1qqD́mYFҶ�3.lr���7�7uӲ�>u�c�=�z�@���h��$P�4��O3Ǌ�Ey��,n�+y�l�ʻM,+/`1��ɷ�5�rg,<�٫B\��V-(�K��c�;]4U���m֫�-vj2�l�,b$�u1H�aQ��hP����b�XP�u^[�39qa����6m=��bz����]������S7f����<�M�Y�n��|3 �p�bб�]���X�����3���'g�m� W'�[<���#`�3��#�h�ۈ����Ʌ2�^��l��2��ѧ'����4�jUXY�0˻s]��b����V �%��5v�AX7�Ɏq:'�la�c��\q؉B�n#���I��k��[#�]pC��$�u��sp����M�myaT���Q�Pԩ%R��ޗ�q�S�� 	�{�ݧj�僫z��̓EixS�%IەͻvI�|{|�=u.�qΎYٳ�����3;���"��u`�<�q�`b�Ѽ�4�d5k���OK�k����0N�܀�{X���J�Q�Ü�X;jUѺ�Q�Tl��W��FLa�R��l��>Ct$��μ��gkc�͆Y������i+���Ky,s�#nj<���M3)��gu�q�����-
���9��}�cF�1�+��7#�Ft��8�q���fi\݋utlaaB��;f�L���qz����XJ���u��%��ϞE�.���`v{a���L�e����[�ODn	!&�^��ʓu�m��O]��۷k�u���1ܖZ�[e�n+����UfnFj�f�a��nN�A8l۸۪���X�0s-89@{&�f�9�ev73M�yZK�¸����痜L�Aر��3,�$� �hGp�m��T�&�4���������9�^���gg�����sUee��<�@�	5����wsb�#o3�]a�Cp�n̫R;S5t73M�0� V���fNzįsk]�����;L���3!X��r4���e�@]�����<�3��l�]Z��=��=��^tx���tn1�ɲ��W�a�Mh��0Ӱ�(�N���3QZ��m)a��(��˙Yv�Z�����5������؎x�<���`S\xZ�Ä�hT.�kݮ�a�vn0�{c�d��#ۮ{c�\�^�H}-�e�pQ��ݑ��V�q����ܱm.�j��P�t[�N���ozXd8��:��l8�^�\��D�:щ�=V���!��+V��yյ

ƣ��J�e6���&kλX�ui�8��3���L���L����"��Qf	�aXh�ݴ� #�Ҫ��ib�ێ�GV|[�2;��R�KH�õW#�ͫ-�k�eXݍ.��LE�\�bAʰ� ��͕��(BF³6�6�vև�mi���Cl+p��=B�`.���c���v����k1��hEf�SB���W]ð�����m[�h�B�03@��M	";kΎ�y���nU@P��smeC9�v�-U��p��a�^V�h+m�V���fU=�F��omrv�8�RWN��Ş@�]=
�I6�+��Wg��C����Ou$�ֳ<n��*��U�2<����ͷhKnՂR�y᧌g�f��P�l,�u���H�kZ�����Շ�;�!C]�����^p�n��mѪ�ݤx�N��a�^�/]�TNc��;��Lh��4)���$"k����Uę[��JieL 2S�x��5i�����=��&nF�'�h�_&m�%��fv'�m�L[��:�H�*ɘQ�[3��܋1��:]5с
�v%��6�ޱ*�rE�ҫ��3���(c1f�떤�{��Ob��i��'k��3g1Ƃ�te�1�ʼ�� ϐ�v�nB�NY�v<��̻�S�n�0�8k=<�n���`�����:zX�2q؇:�uۜb�N��%,<vMX��9��<�r)�lNn٤�%��3��a�H��X�\y��H����imZ�,.5�ul�m��%vn��l��s�Ӽ�
�oW[�'N�m4BT��N̕f��lF�������ŤkEԕk �-ݓaJ�m�t�Zd{#�sIYWh�$mu�G7)n�y���]��<��n&��'\�;�ܗ��5�{[ir��� ∔�f��aH��&�,���R+v�B�
C�Ա��iuk��4�^e�	Y{rD%�t�mf�U��\��ַdqy�ɼH����Yc3&�kZbЕJdR���&�,گ��'��@��#uv��8�B�4v�y:,�M�d�ڹVzYfB����ژƅ�ΙdS��c-�w*��895�u����cK(c]��:��@��&Gz:���ϑy����ҝr�S�\�v+k`�c��)n���Z��i=���&o4���抃a�0�b�l�[���6��������&f��T�W����m�r�۳n�����Gm�ĭU�4�.�c-uړ2�$2���'GR[gu�;�1�E�Ɠ�����ϕ;�Kq��n�=Z��xļ]� 7\����`k	����q��j��[�ꮶ���t�;^�4�28J8�2��L��x��t���䲈p�ј���t�!��l.��x7�p崛�����v��\��7M�n�tI�E�u¡�E�q���Q-g9�/`ۓq)	h��q�ٺ���=��"i�sSC�k���Z���m]<�ɉtnmU�B-t�:����fX�7VuEY�EMs�UAj���e��e�����n�gT�\f훍V���Vz��l�ˀr똩M����{e�t͕�6��lFT���7�8�攁Q���G�<_=a|dY�o	[b�e�K~>y3M�^��7<�M�U����^].�)nԃ0~�WƐ��Vy%�md��d,BL�#4�D�=I=>�����/�����KS��1JC�Ɏ�:���<zQ=C&��xz|||w��l8��)�GG�{��ʪ3ȈGcx�jB�_���4�z�OP!�3�}̓.%;�����.[��@�F
f�e�d�F�N�]S��B
<�S�2)���������ʍ��g,Ylh�B$2!T��D�J��T	���(�d� J�
�a�Lz o�-:�;b�H��3���r5��Ag9��)�����B�N�V�8l����Ju�Jq)Z�Ij�4�iD�S\���½��˚�������A`���_�,�d-�������F��r�0H��y��w(�
F�˝H���U�6��e���Xh��Uy��g$� �9U`�P�c:^!� u Zr:����i��/�!��i<X�RX1�	}WA����:I'�~���qu��sWd�(݆wt3t�xZ����<L7;�]MSp��ɶ2fyz�LcV��d5%���u����O����tͲ=5F�E���뇩l����1�m���n�Y��&�I��S�F�ϭ����]�]� M���=ss�cp'I����[؎�N�e�u���ܡ�&��f�U����u�J��j9�<n�fŌhh�Je��5KT�����3�e��p�i��]�呁.P��������3��#b	�سM��hٙl�h��V��Y���tW<rH�G�[��TWK�/8��mє�iv�|�.&�\n���$>ݕiP�]ݵ�����r�-�v�U�JjG�h�nM�"%�fҺ�B$�JƑ���6����9Am�=��:�7볨�]��7y��
��et��e���T��@g��Pe����qR�+R�2��Mƥ�Ѳsx��^+�dJܙ���Q�Ю؊��91a*ѵ�*qbj6�ʴ͓X7���v�
��>���V<oe���u#��I��&vUη�D�e�lju�]n�n+)a��&4��!�b1���p���3g��9���2�iq#,n�eZ�ڌٶc31l!]	lı��RS
���!1�;Y�BӬ.{q�R�ڰ������kɍm�n`U�:�]��q�-)^p��`Ȱ��lvx9��';�WL�!�����lzN���(�6�����a�cdm��i�8�o(m6�4��-m˴����H�{qV��lu�)mp�
���c�|�I�KD=Lk��I��ت9ut�pr��-�\�����:!o"�>,��mz�-��6ݞ�ֳ�%-�[A����(,\�U����KU�v,'7n38��6�a[��^ˢn^�n�҂��v���)	��B[��HQ%�cu#�1��f|����^�x��kDsp�se������ 7N��LlF�Yl�-%eږ��aicaHP��� ��
4ĴTiѠy�%��Ĕ#Ke�i)+e!�T�V��^l�e@e,G�-�`��"�0��r������ڬ�
�,ci�"�V,(�ժ�j2cB��^cS�
F5�B��Я<�*K-�V�Jش� ���~���_�)3n�+l޼9.wK��v:9��8=�Wu�Mҵ��w�[��|���7wSmYi�JGyؤ��r��-�2�yM���>��ڭ6�E�Ϊ�9JY�l*9Z��U��6)�X1-����;�o7�P�۟~ӝ����O�m�D�`�s�3�N�Y3x.�෸ZAn/�%i�-9mG�ߩ�|uK���s�d��߶uv�C쿲Z��}���S6�5��E�whUf>���e�n�]�*�Qtf�>��ުoUR�|��i��O?4��=O٥��FSfT�����s챂2�g6
iN�#�f�;�V����|m?[V`��F��Ӹ.�跸E�l���E�+��"�xU0�0}��L[�Rk�X���}�m�s;�f�������(�ڥf^�{����B�o�w���yҚJ�U�5۶���Fb���#�,��d��~޶[���̖��X���4F��3��VZs;;�o{/���/O�]i�\�ߴj�w�f���j��w"�ZcQ�d����0����[sN�w��n�v6�r��ۏ�]U@�aTª�����l�43*��Z�U5[�vQ����]�-��t~?�p�1g������w*X���0.�p�>��NƮ�7n��!w$�p���31v{����
��Q�3�u<NF�F�S��71o	DL�����@Zs-6ԗ��P����їW��_��[sN�w��nځ��v�U��z��C����O��]�����Y#�e��C���8�{��A���%��}G�����v6���z��������>µ˖绯��\��o�su�����;����U�l��'e�-Y�j�rڲ��"�#Y�
����1	���eK`ů���ɪ�>���y�+.��i�}�scDf��ј���v�P��fe���������m��M�>��s�Nދ�ER������ǋ��pt�WY�0f�$,: [�]�[�m���i�Y�Z�n�D5��5r���'��~~����`pT��[�U/Z�lTʹq�ǕC��T��e�T�ww Ff�h��n��[Jы^'uݓU�}xa�ٙ��l�U�`���O�.��9f[n崱�.�"���Sj�-qBUaWO�U�����_Z~��V{/2_����۫�߬����N��}k��j�3b�UR��K�ϒQ%(ʭ[a�Hw�tN(�L���5'������=k��ɍ��G�yc����3=3� #�tʤ�܃F���f�͘zz�p��b�����jӖ�j�q���U�D`wv�Z�D��wd�b�\NU!T6��)���c�2�mcv�1�MnSfY����xn�M/K�֠Ru�,�-`Q]���
�Ӓ[s���O�U����u��b
JbkP�oU0��T���Cq8�������'�����s4/}UW�i��*?W��>lS�f{/�ϻ�v��Y�B����՗Uo��)��Tª���iX8�']����V̖�@m��o
�Z�%�0M��j�E\P�x��i%߲QߞZs?SmY��N[r~x�-�É�!�o�-�]���.w�ڲSi��[�z�/�%-�M�i*iS4��2��4o{سs���/-�����{sTA� ��|��F���I�i�S�m\���n�|~����׾��8�<��A�H�_����g;��1��y,Lr؝{uue�s=q���	6�8e�V��m4ˊk1Y�;�8�vM�N98ݞ7>,������ ��BU�������PՆe�ݶ��K��α����Jۜ�r�[�^�Rp4[]j�Yn�.:티Z�!΍�Xh0��Q"�S�4εm�*zāy:r�r�Ɇ�NY6B{uN����.�U����={�F&XML��[���G6��v�e��K.�0��cr�e���}ϗ��}�QP�o��P��c�V�zgl�O�6oM�Q7�[�Z�T�*�k��֊L�P�h�����Mbс�pM��oM:,N�<7���b�E�f�"W�;��o
���Vb�"�c��>]Fn;Ƶ�	�//EܯM8B��=$*�+�^@W<�­�Sb�X��6�V���P��(����F��ҧӠm���j��U)�R4e��Mg[�<�[06n�����E�צ���*��S��MH�A�svY-bIt��!����*\[-�@��]Y�ݵ��23^Gu�����;����M�fZsś����/�s��gL����>_?�����M�]����z�pɥ
%��7��^z� XWt�/�7s�����iW�vx�)�z����1N4kFBW,�a�)�;=�B�d�mF�?�.Q���cU+��Fukl[;e
}ꪪ�X�6���_\d���Sz��\8--�,�oQ�Qbv�JO���1G�v�V��8�R��Z��Ng^ܷ�=�ߦ�[�yl�߳�i��i����S�)̶���x�2u��?5�{%>U����{��<t�go�Y̹m�`���2�<���|��λZ4�@��L/N4 T��i�3\�p��Z��3t�ѫN��^����M�h�ۘ"w)��&��E���.����/����_֜��Y������w3�s1��j�^mV���"��P�oU)�hj��zb����[U�-��p���o�*����V�3��M������v�߅�}�~���?v��,�}C�)w�FN[�$�{SQ]��.y�(��#:�Q�uf��|������o��_��`z��b�{_o=��8������Im��N�4�֋��SO��޴����́T_�i̴�d����3�&{s?2�#ӽ�ؿ��/-�;�tV�N��FQ���?�(-���??���MtV�v���\'hۋ�kv2�	�z���.�r�`2$�>>�\7��TުkU;P�!�t����N\��S��)�f�ꪧ�U!��Vf�	��7���E�2magSZ.N�-���/UFe\��FƂYk7����SUU聙C���ｺU�������g~�׊Ә�@��(L�'Bf3i��ڽ��U7�T�BxQ��g�HŠ<7��<�g%�����)ӻ������x<�|�l\��W��mx�T��ў�qξ׺ow�e�iJ���W@��VtG�`��X��NZ~���Ӗ�����M�U@ju�1�]�0��즴[�m�V��ǵ~��T0�B��3V��.���Ru�ct����v��e�R�٦b�������I��ݻ�l6nU�Dڡ�l�"��ֽCj���խ�B��T������2X��s����;�g�V��3z�ª��5.a�i�Sy[	�D��`*�Q&���!���7�iQO8��<֋s����*�Ne�י҃ީ�����|��E��+.�v ���i�Z-�e'wu��7�dæ��z6ת��L����f�����zkj|�a��kl���´<0�"���G+J"�lMZ�\�FG�s���t?�HC���k�cc��O����Y��;��gns>/#cB��xD��S¦f�Mb��i�'H#C���[e%[�#��sbفm�<Y��IM-�$�٣+S�Y���ս.����a�v���5�潒z����yJ��͕v6ڕ�w4WZ�a�6��Z4!�rU���Y��m�rG:��Py6nyt	6*ѧ�ɇ��ݴ��oN�b��]�ܜoBb��Y��ng��n:�sv9��]+!��7gL��2��5���e��:9rR:6i]�������q[������ٷ*�#/=t>�v��bŶ�n�N�ɛ�� .�U7��nIU����}���{���Q�~�R���gwwN�n�;�&	�z��[w�j(m[DH�p�*��Ov��0���8l�w0T���������ыvwkG�3��܉��xӋ����Y����~��[U�~ �M�=Z�}z����ުoUR;�UnƸ�r�;f�����2��#��q��UU 
���U^�Q�R����z�-�����QC*����Nk2����o/a�g�؃���z���U��^]��k�-��c�q�W]�f��'���`��ᓤ�v���ު���ܚ�V����*��I�ޗ�u���ܴ��j�9��1����]����>|�z���L0��WN��ZS�-���������57�?��sop�ZA�s?��n�Ծ;�!�2�p�&ձ@��G6��ݗ�B��pte��M*���ҕ�i:?����̴�m_Z�p�?�5 u�v�������߱�_}i��m_<�{G�U�6TX�Z5�}�yl�ɡ
�n�lc��Hi�h<�tӑ�����U5U!`ݐ޻��c�H�X�Z��Ҫ�e��3��7G@�l�B��P���u/�p>�=~��!]mae�74����"��{t��x9���R��/&.Y2r��hl���	����$���}�ڊ*�$^�oUJ	�n�LA�7\?)�2֭?Zp:f����|����dЋy[���/1-��U4�5a�73ke�ݽwL%�·j��M�{� ~�&kM˩.�B��垙��Q4�I��AnOdC�<�3qn�H���ճ|.�K�a����s�+�x�g���41�k��_ͼ������=5�DZp�[�j�@!�7��E6N���{�9ɿN
��F�/s��mID�6�cx�{�9Ɱ.��5�!��:/�:�:k�#�#}O�ݾ=��H����g��x_)��~�Y�+>����y�v{��'��y.eq��9];��M���Q�`>��7��jg���Y�j��p|�_f�oz^*U�ź��W�
i��wA���3��ĿI<�f���r^��;�X-�>���ˌ�|��P�S�;F	$�[Ǹ�����yn�L���/�t���Z���S;�z����wb\�Q�a�<=����O|rK{�-��&���V@<ϊܩ{�������6=DeN� 3ç���g��n�{��G��!�m�Ch��'�|�ˬ�C���vӊ�gu�Su�����b������w7�f�"x�s7�w����f�����+v�LRNz�KZ�6u�j{�b¼�����y��z���}���A�����OΆr��������d�<yQ�뾳�dk�\�������4��y�b�sg��w����rDC��ټ=��>�:N'㓧%���;Wn{���f�BOE�|�M�v�rw��瞙�oaٮ��q�Bf�E���ҙ�-�4�����Yӂa��e��/��-���ż=b��3�L���z[�����1��s@�ud^ k�X緎���_
��^.C�����ͧ|!���i,�x�G�(�	�"��8=��N�%�.I)��dA>.}�gB Lp�Rg7��Ӂ<�;.d�v�b*$�L�c���^5a���11OS��=Oq}��g�O<C�<@�N˗�"M��2�����eHBф:�і&"c�19&�YFh�w%�9��<����N�{�}"�[�ob<{�<�1<d�����P�'�i3�9�[��B�hX��X�g�Ob����=C�5"zW��>1����)R�w�O�~����{r�ke%YgB'����$�����rdU��mP{��\���]f%��f˽d<��.�x K8�������G��x�4]ۇ<����=g��ZtQi[�f�"�
%`DC��t`�^S�d��V�(�s:�3�aԔ@�B�oD]i�g�Ȕ'��[���d����dH�@S�^$���;��f�ƚMp��&%�\k� `�d\�D�QRb���3�=���/	���
I<�H��i'���gd�UI����Q��h2D�F+��8i�nГW��I�n^5t"<����Qm�\�T���^cjxʙ�H���^2	u�W�bZ��ǃ��*RK��ZQ���"�?&{^l�JbzR��^iK�s܋e�5gR@N���kԍ*%\�\�� x���*�.\-��;f�[7|w >ڷ�n� �`���R�3tg�eu̜�`(E��m��ݯ.�x�������Oo ��p���E�c��{|jA���]�>�`v���{�뾳\�2�pU�u�ס�J޶�Ɔ��l:���hz�צ�z�.��4nxr�O�X�WQk	�+�X��Mz��և�<��h Mb�;�;�N�:y�	����k��^wh�Rk��w;e�k�f�w]?ɓ���<�Y����a$���C3$8')�"�`�����h�~""\�"�y�x������Oow����"Z�j����݈E�``yJpGc A=�<�~�]��7h6P����S�*�u��45��a����B��_��vѡ�Y�xu�r����bY�Z�'�#�O��jk���ir�W�c7Iu�� ��Giָ����]ʘh4�Uą��5�^1y�a��a�vHݯ��zaR��Vu8G��o>�#o�6]Ȝ[	����
�4������˦� 6j��A���������^]���3P�23[���7��3l�eQ��|A/,� ����dA���[P<"���O�6��P,ɖ,Me둫ַ\[�]m�:�����e=�=HlGd?]����%��p�퀻` .٭8�[�ۣ���&��xD�SS�k ������v�F�7v������������ ��Gu��7��kKT�h�n� ���FW8p}v���[E��,#��"2������]��ݯf�u��+j,��˦us:��&&S�E��F�>������U��Y�e���w1Û��v�[�Cq�[�ۣ!5�{e�?�KŇ�6'-�kD�s��ڼ��#�wi�>�^@ݴ�v���y�4���p������*�[7�lÈ#+��l$�,-!Xe��L��d:�8qT��`i�M�.�yFKlM��9Y�X^w�לfB�X+��y��G�k�b��R͎LI|�݈�a�tP&˦`Ė�LJ��X��#�V.�"mqf�x(�<g;����/Fy�Y[]QT����@�������45��L���p��p��ˢ}pe+���՗rE�N��g��H�g�t�����.��46�#5�Ԗ^�LE��66Y<�av$�,Zn���������E������5�Er`+n���K*����2�0��L76���V�`���v�]�;����-�7��E.wHc�qvպ�=0F��8��]靷�,xް� wn�"�x-�j�8�Tu�:��kn#��P�1�ge�8v������;R ��@�ݯ9l� ݷ���kBhU
�fa�H�`���s-�mѐ�3���p%� �v� ��q����w���~�n��Nܯ=��@ݷ�����E�5�����+�z1���� �n�?��Ahz���\r�=jz[10���'���.��El5^G��N�g�ۈ>12�o�	5z��{�o���d}W����y��`n��l:����D�wAӕ��J޾P��3�6_�vD�pA�Eݸ�vޑp�V6O	�b1ʃ�3�[��s��{!<��&[n���k=��8���v�����:W��x#�@�滴{Z�3�6�[�)�����lj�'b�0�GM 湂]����pA�`'��zm�m�#b�����H1B�Y/�7jBLc�v@���)��yN��Lfc=��?0z�j��f�g���l��>�����Z�=b�Ẽ�WCU�qn����s<���ey�'��y n� vR}�ϛ��hs�I��=�� ]ۇ7l v�Ï�;k�d���m6��ğ�w���bX.���p�7k�0k���j,�z�C�q�X�i`����Y��f'�:���n��2�c7x�c �o�ʶ��3��2z���#3<����:f �#3:*��;����M�T#a�64�WT�v��k`A�)� ݯ n� @ ���n��״xyZ�dϴ�"�X�X8!��F]3Mv�e��8͋f.��=u8pt����:���>/l��� �7h6�զ���ڙ��f�i�8��Kk'���oF�a���fC�v���o#wk�Cf�C����i��<�Ky�N9���9u,t�|1���/v��vå�kS�kkʣ�����o� E�Eݿ�ă��ޫ\JhTm��D��(h��*��5�	�o�a�R�M҇�n?z����{����|�;�n�_�� ��O��]�n��;��OJ�.�� ~kތm]u4�,o}�1+��א� ���pE�x+�;k����7���5N�9��ޚ����w&|s��O�!������ˀs�E7u��^7��g���9��ݴRc��ѵ��`��k��U��+���Le��op9��v���8�`�X�_�t�V�m ��	T|>KP�A-�*��Y��j7�6i�h@�v��ϵSs���4lS��kL �"����v���B�ΞM�SA��y������*��J��2�����N@�o#v�s�gL�qZ�+1����y���r-;]ɟ�w����,- �����z���K�!��@9����.ב�d��z(ԙ�.'�v&�w�f2�c71� �n��l$n�^ ]����ƣ�S�0���J]H9�k˨�*����u4����e9�XM=.�	��͛"�{�w��a 3��Qi�`�� ]��y60�S<�Ɨx�S�˱`��핗x�y8����I}�[ �,T+@���p ����PC1�	|`�I���ݰ�]3�ԑNmV�C�Lm��M;]ɟ�w���bX���?�k�[@��7p�9�*ܗ/���	�d�����{QMJ�v
��q�Pp&�lV�L�:Y��_98z��d>7v�b�M���4��|�����0�%&��H ��q�"���fd8'1�!�8���V��)��O�����o?��»ΞM�SA��y���.W��v�{��t9qJ���햒�`�Av����h��U��ƉI��x'������)� �� ��v��"�y n�{0K��!�޵X ��@>����śܓO>K����9�>-l#0�ΥQ��S�p���Fb	�wq���>b��}�Y���Zח�aƻގM�=A��;͍�)�]�/�Dn�b��k���]Jq�"�f�L���q�����af�vﯷOE�C��:=���Ov[��pM����Z��-���y�_�����|'q(A8�j٘1�c���pg0�
�l�Z��#�������Ŏ��N�5�ez��	vm�eBTb2&4�䪦闎K�ud�2s+,R��F�Ճ-����c����&�B,�*�\���/(��׍lz+4�s;Ϋ���K�=;�ɮ�H<��ۅ�{q�׷n�s8�n��9l<)�ۮ���a����ן<Z�X��2�Bk�2��s����������h��	f��n�h44���{kr�x��e%��	���%��V��턐n��V�Ri��	�>g{-�8/�E�m��k �����E��7m��	���;��:�/xzñ�G�v�\k�s&�|�������,�	��ݰ����ml�vP�44 �@���r�.�@��w��xNY7xΓl�g���1���[\&-���v���"�����p}|G5������M޸p}��!v�[�J�&�����w�b�������D��XѺ�`��A ��O���� ݶk�w��zf�\�����ɥvKd>p�n>�`/q	�$]�@E�2<o�>���Z_iJB`���ѻ�Q���rX�d���Ö���j:��������?}�����^�olk4�wR:�:]��[�F��v�D���b�m� ��X�Dcz(n����6��.�)VVg�:i>��j��N<�9�+��e�?hܜ�?^�93�6x�ɷ��M����;.�Z�������WoB���	�C�S���	lm+�M==�d��
��pLS<A�Bö��.u�e�i��[�}^^�ޭgW)Ȼ`.�  �wk�[��ÿ0�Zj�4Uޤ�ه*�c7�Kf��`�Fc ���2����wɃ���	��z������2y��w��)��n��A���,�����e�@'6�'�l�&� �ۇ�`g^������ѕ��j�dӳ�VA���Z���ڭ����wn�]�&�--]k�ۮ�x�6 J\39>N|���㞮�ώ��4�b�hnK�����T�VˇW��~B��91yx�� �wiƭ4ٻ����ƨ{��z��L/'[��ه A��i��l`���?����OCF�-��}����G��_x�(�x]�67 A�1R���1��j�!�\�P'�W�3�x��{� Av�9�`�lh_V�������'�oI�U����4���X�z�ْ��ֵnު�9"�4�KQ;bb����0'��@�e�Ӷu��Ĵ��zx�J&b��BgY�p���kqu�S�\�����_8&i�v�D]��y� .����ooa�m�R
����@Nf-n4ٻ����ƨ{ь��rX$�fo0**�y�'��[]�n�yz�Eݳ�pR�{����)o^@�[��[��q͍�LT�v���e�뻀��g�U>�k-��Ɖ�٘^)��Qkl����6-�M-�9ڡ@�(͈����/�� ��0}���E��ԯX��V�<��o��8yG(�������/�Dm���nӂ�0#���I���.ב���Y�e�<Oo'妛7u�)n�i����rX_�5k�]��Y��C|��+eÂ� �v��v�v����ppkT����v�&�u��s�'���{�����\fn5�GY��ζa�p浂 ݠ�Fҽc/�\�����]��� �y�y�٦�}"�o;p�8')l�7�Nx�va=����w��-:�#E�q��Ԯ�3���x��:��s�����OmS0fViM����Ǽ��㜳�ﻶ���m���ۚ��yv�d���@�Rfv���ōd���46�4�ތf�'%�@nk����v�Ȏ/J��� �YQ�ɝ�o�A�������Mmim���պ^u�i�X��ؿ#�׹��[h Eݯ8�^Bw��|�+��q�����$[ǌf�U���������o�w)�l� �,r�]�5�W ���[�)��۞�_;�k��f� E�fc0q.�Y��}^�^@�2���p�o/Xcl���S��j�#9��k;MZhl�i�������x���ݰ^ ݠ���$qq[dk+L��>�A;�䋶�6q�w��;�S5�67MT�\��f���f;X�v���H!��Àn�f*�s�Cr�Z�ZS�U�zy|�e� ��x�.�^]���v���!�x ~m�iCw��s��^*�YC�]�<�N>�OÖr���7N����RntZ3�{���������Z��o��~=��z�v^o�
� �� ���+�!�h'��^y��b}ugN�ȿ�ݼ�>��!�-A7t盃et��y�+3�<}�<>�~�c�t���rƫ�6��=S����wf���?z��84�	f��}T�"�o�k�����|'�	w.��{����`p^���i������Ϸ�V��"y��۾����rM��礭Cn'���ؐ�w7l����YwQ���y{;�f�aR��.=�.K�Y3����4���By�3BdT��m�'A�'��ǜ�R�y^�}}6w�#t�罜:j^V�M����iY�Y���X�W����ׇd�wxe�*����[��G�w�N����ԏY�ⱒq<є����{��'�%�}+Xc홊z41j���Wz|����|�]|�Ƶ��|��x�m��������&o.��'�Ǉ_W��qǴg{ ��@R�H���e�3tˈB���m�e~�;��w�9c��bQ��;$~���JC��}��և3N����p�Ź�ZL����n���w^��v��*���m�c�{^���*�Ɛ�}��F���/EY'��	OWk8;s��.� x�k"t��Y�z��Sc�����Grzy�ގ���c����#�\W0jh��_h/��Bi����d��e�c��KoO��>�sݐ��4�ؘ��㫋�p>gw�p�~5.�y�:��Jw������so@�6Y��j:iL��5�7y�D����וA�+Џ�֧�No��2̴��v&d�z^閃�X�1��~>>�g�y[�wZ�F�d3ܑI-g����Ir�v9%cJ� =�Eu=�������d��'��������7yl���{�a{������I��+L���IDc������I��]$��.K\�$JB��39�������	�؎U�LL]5�X��*�C2%�C�e9�yt�������y��9պͮ��v��ݑzTu"������7s1*�1K���GĤ�!�!!�09$�����{3�R�M�53�JEiob0��x�Z4�)�;-Y$� �5'�+Pg�UDT��D-�g&C-7'ɔ��;�5B+AWH��%-��I���"��[�|�8QA���%s�*�]�Pc���I�x;C���j��BV5�4�"� ����'ȑ�Cg�*�<��G��lx=fm:� �I�Zc/�yIH��Z؝%,,�t>�����I舄�S��H���Q�\���\�2�'*ԯ���^VjC�!JP8�S��~Z��5���d���'��֙����d�2�����sDdNW+>!ٮܳ��']8ܻc����]vׇΰ���d���Nx�j�s��w�%�g�q�gs������L�P��E��N2��U��݊�6���ܳ�y�6���p���\���a�׊���jkQ�m#�H���7n��<��\�1�;�ڸ�zbp��=�i��<��4V�Å��v�f�n�B�nF4��������ȋ�,lH�� �����.M�9�&�x��V,u�'zG�J�5���0��]����{c��T�F��Vѹeo>W��\E�8$���\nM�؜k��Q��+���GvG� u����Q�V2�8�z V�[�:�r�lղ�ye4���Ć��<�h�ė��qyì-�Un�k4qY��W�dT��;s�m)����=��-ˡ��������5��&^e�[�75�u"�^t �vX�$�d�C������5�uj��hL���ۂ̻�G���f�ܦ�V�)�hh�:�v�5Z6"�/R!O�ѕm�{]{K�Xq�9��	\�8�Kۛ��90p�g�M��2�զ3�:�Z؄�Vc[v {B�u&�$�j=��cp��x���n�k�v��V�M�z������&�Ge%Yiۂ�YlUEG�x�Grt�ۛ���]vkۖ�\k�Y��d\�L�ID��wO#ӓ��.͍)m�N1������;r��R�TF2Zr�]6H蹝(v���t<�[=mr��[�ڻ{{��[��sm馡�.C-��&��cA�����C,.c���٢������p+l�GmZ��N��[u��!y.�/�m�������M��H�)z�Y�v�t:h�ݔ�fZ���[6q���f�-�"��p�s\Y�������mitTv�����P�Iq�m\�U�;�xI;�T���Ƴ�G�Yx8�͝׭k�/K�y����>M�!�����W	>j:�^^dꕳ:���!��:O�N���'w�Ӻy,<�����[�U���Xue�]<8��r����XY���2�����rE�a �ש�[%�t���F�:l�;"k��]�[���R��Kf3].2H7��M��nã�p�+%��@�X��lm��je�Z�[���֪���K�H�/l
������s���b�]E[��k����z��׳����Ɯ�ƛ����֮������Ғl[S�w u�tdf�tm%�VX�l,*K6 �n��˱�}O�����W�����ӌ\Mf�%ٍ0���`��αs]�,�Ab�7XO��j��([Dݱx�������j�X"�������';[�x���͍͑��R�|+l�ᨶ��(@;Z���I���� ]ۇ5l�ht�7Ϣ,<:w�Ҳ2��җ��Z���`�Ah�^��������)��pM�Ku 7D��w�����rPݘ�z7�KF�ǠcԎMמ�`2� 0��pH�o+��v�m�U�kCF��Ly�mu�̸'��l�嬁�JpA��`��`.�t62��o@�i�	`�hk@�vl�p�p���A��b�5�s���"���/;��;-�FyK	?�1Ñ��Y�b��Ӓ�:���*��k�FS�a�7��ա���]���)[���`�5�  ��pG_
״X����_�'�+^�n�Eތ/��������'�awg)�vK�y���Vh�d�"�u���
���Y����>�<�|u�9��y�q{j���f�[�秶���fky����~�����{�a�1��������`�#s\��Cx�k��o��A؄x��DU�w!�|n�L�F�B�޻���޶\���ln�`j�y��`��dA7v��� �{�<�A����(ƒ�c����[I���_{-p� D�b���x��;�y��`�7l����vŖT�����r�r�Gr0���}�f��nj�p��v���4�q�;{��?|����o��ֳ%�1��G�2�j��&�F.�%]�oE��.��h���e��A.���v�M��v���)�y�G67�ު����F�U���7�7v��1׳�m�WɠBn걢�pA�As�W@�]3���C_{-s�,�d"����Uo��o]�x�w59`Xݰ^��S��2��U-\���3��Sp5`Br��`��	���C��vv�y��;�G�lPe�R�S9�	�3�??Ԕ��z	=5�����W��̫4���W�f���?e�C�z��!!��Ls\8#1��wr!WV�7=��7Xp5���r��ݰ�i����y�cѭ��>R�����i�a��oMv�Q���!��)S���/�W�&5�!n��Ev�i�F���������`.�|� [Y3�[�9�Y�I;:.��9��g7Eq�Q�vi^�B'4)�3t�i^cN�����<�=I��Ϯ�>7v�ܴ���?e҇�[���*	����Q���p������N!D��twv���|FU/?6�<:�gn�d�:ǣ�����怀�C�ݴ
.��5��
���(%7��V��ٲ�7hpW1�2gO[�旻��Ff�����\��Ex�.�D]���fυ�X"�b�Z]���9��^�k!�F�b�k�A�������+�E�7�X/�+W68.�W<�e��R�b�I����?K������fs�{����{�l��]~�h�k��6Vdܾ�&j�P��5*߅��3U3�
|����~?�PD]���7lpn�8"�uWϭ1q�:���i�`�^�Ѻ��9�'��r5���j�y�׬?������c�WkH�����=�&��>�5a �#|S��C[��b-FirR\��ja�f;:�O�_�c#s��lݡ�:�5�i�x=�/[���3:�kfל�	{A}����n�A����+Z�:��"<fY	���j�k7F�4;�cC_
-��;,�;x���g�;5K5�� ��<���D�v�"�ל[Y1��{SN��#��y���'	����5R��2ב�dA��]��G��ȽL�S����8{15�c[U<O�ｸ��%�#���M���E�Oh�9���b��7m�ݧ"퀻f���ע[K='�);�o3ÿa�W�ٸ���A���a �v�hUݮ�ʃL8z���߫����Y���ٽ����Ji�����B��(��ڇ���U|<9:��^������:��o};��3B%�0�w�픳J�*�I��x�l�l��&�Y�\���n�۬>�tt��BM��8�',�� �D�]��5ڋ�n�n[�ʝ&�v�1!�[�9�֭1�t�1��=���٨����J�RW�ZY`h�Y����bݨ��wR̆,��͇�Ƚ�P�m)��{K�-��%���.���3@m��e��B�	l�nź����l8�l\ʍ�3��,�оygϟ!���f4�8�$��X7�6�N�r�nx5d`NN�*r��ܰ@�ᖂ"�����yTw}|�vt�<NG67x��bEοN���u`��d#Z��ݧp�͐����s�BYn�p�t�D��ǉ�m�y�|_{q!ń4��]��E����B� �����@�7�3X�,�v˘7�f-���NH�@�Mѳ�n��w��A��͛+�]��Eݻ�Y�^٠V�a�� D�?�ƚț��q����t��lop5R���dM�ӓ�G�m ��'"��!� �0^#38p�t3oS���S��[�Vt��y�1|_{u!���`���網-N�,��b5E'f.��f�wd�ѷ6���vM&Y�µ��Ԗ��v���|����<�\�<მ�@��S��wst�w�9
�Yn5�f`r����\9�(�.ФkBM�>ԹU�ѭ�7%mn)CE'<�5���K`t?\ �t���K�hˊ�Y�eZ��]KwA�I��7���z��]4��c�� {�@2Fj$���~��z�u��w����>�|9�x�''�ۈ �J�Z�7m|��{L���nzn_'xib�0^ �Mۇ ٲ��hl;H�-�Q;i���1]�ԇx���7h".���[Y�@��y(���������ͬȂn�X�~%�7OC;�a�W���@o6�1�c#[*��^��m�����P@wn�l�Eݰ��s�3�V��o��p^��c��r�'����	���^@ݲ ��K���4N�T�C��~�jiF�L���ir�16׷'i%��:ǃ��m�F��$�;,�rX"��Ãv�x�v�ɉ܍k���1=����q(��t�n�����v� ݷ��i�E�f�҆mh���6ԍZN�n��w]�!_f���㹎ݰ�����>�l,��׬$E�wn�"�zQ4��+���LJ=�fy��-��Й]���j�ݭͰ�F����dN��S(�ݒ"&7\lT�ۧq"D啐�^~y׏]w�z�^���ȳ$fP� ��#�  �`c�l��'�����r�y�v�������Oa�3 ��-�1oz.�L�R��փ���.�,��͖h[�;	y�f�1,)����5�X��㒼��v�A�לU�.�2&M�i:,"ѩ�+����<]�a�W���vX71�v�]���mV�m����\x�N��Ӏ��P��Ehsn�t8�n�����[P�V����l��B~k�w��K�?l^"��?��^AN�lOQ~�<NO5���w���W��-��׬�'3A8��	�`��;�]�4$�0D�:^w6Y�lW�%�A5w�bX+��Z��/�R_[��r� ��ǵ�9�/ܜnא7m��wk3���5-�qb�k��;�Í��}��F�8v�x�.РE�ϜL!ɖ���
y�	�\?����kf�e3����ru���r�8#{�*ӴCK�6��q6����У �}t���|l緟Q^ol�G�{ْ*�N<c�1] 꺕�ز�'MK�Iמ�w�^�;��񽪽�U�VdY��JNz����z�}������3|��v���s�ڄ�څ�MK�`� �����2��5�;	y�f�pA�`�>�@]܇����ێCC�HxsLe�f��ve��w`�3zm���T�8��`wP��.[�L��:jN�E�[i�;�Ƒ,�ۣ�F�Z�!�nh���Ne���{m�5��$�W~}a$.аA����H.���:��S��G*ux=��������(��'�ۼ}�)��y��n3�5�&��n'n2 ����p��.Ѝ��X�3Y��0L������R�`��Eݯ]��ݲvE�k�kv��d/�@Mݧl:7s���E�����v!�]se:��Q�>�a �7i�eE�n��G�f����^��m��4�!D�<���+�����������]iw��"X�x}u0�ed]�5��L��o���{��kiԎ;�`��W�����}�@o��wwz��>�=5�Z9�|�dkD�<<��ϟW�o^>s�]�ߗ\�s�{jj&hL�J��n>6�w���9��y+m��eal�-��s2u������_ ����7nf�.���s�%+<�!�	u���e`���j@Z�m.�M�ź
�T�B�P)M+��:E�GZ�F4�fr]3���t:�Mr\�j�a�8r�\�6� �����(��,�cq$�Tu�a\f��#��^�)ن֭��D.�B6V�M�4�Ҹa����3���X�2��&˂��CK��X�,�ƸnN�Jʖէ�����;�D~q� �;9Â.����~�Dmp��^7٫��)^�8Bn��u�SQm�.����v�x�@A�������������U�����żC��8�}�nv/w1��X]�*ݫz�Ro��dv�]ۀ� ݰ��J�cF���ED)��O�P�9�5��+��n�MݯY�!ŏ�����_0�a��A�t�^0�׮�:"`�p��^;٫�`��
3�%'��lg����:B�>���Y���綣���$�O�X{q��w���/�����`����6h|��^W1ܔ�����~����1	����0.��Q�	�S'�=ԐF�8�W6��u�~O�_^�@�z/��,"���@��'�qlp�~�C`�kn��S/�����j#���N���p40Î���0^��^��3l�4�C���}d1�Z�LÌ�v��f�Dz��%��[��خ���r~�9�K�n��߁ ԧeݗj��=R��5���r�ұ���s:�}Ğڅ�2&h���N>2~(}�!�΅6��K��5w�2W�]�.�2{�6�����N���e�&nל���wie��]�#s��iǬ!��(�������8sv�v�]����Lwv���G��V[[����Nn���ʹE'n��m��ʤ�E���B�6Aҩ������x��`m������]�k�W�i�޴�]y���dup{�^;׫��bX"఻Aw.��o(����H&r���c��wJh�(jh�@��7�����܋a�fwd���0���/W�7l����p�{u�x�{�8�8c71�7��r�F��^ �Ӈ5�]��"��8&�j�i�/�8(��?�����ޭ��O�r�߆q���M' ����!o$L�t�'�Ѧ_�Ά���P`֭Ãv��C��� >�o��}�G�&躉a�	�`�p�:�ط7�6��T���=V�UK��k*���Q���M`��q�=����>�A LD����i���=1V}����%>z�n���O���H8�o�����̓���Ga�]6���g����'-�=Ξ�'듷���^��xt_6J �=��>���v���S0�v�>�.�I�p���*]��e�[4�}W_y畦���cw"��	�X!��JLh<�8�ͺ�9�v*5�bfD7��XA��s����$pG���@�k�q�r�,�{�fzwo,�gV��w|�o�� �}���S���4M�=�/wy��.���ƽ1ࢩ��h����a����;�~l+���n�+��>y��5��{���{}������OB�:hgV�7�k&v�Z��Y9:-�\9[1v��{e۷{��<=�tN]��-#�#/�~�t�D�۾��;���~��}�pD�ɾsvy�6N���[�c.�4o�}�%�Y����J^	���^FW�͘��"}�
�|G�`��i����o���i���A���/8U(u�v�y
�O�-#����T������\��n��5��֟u�J4G��f{H�UOd�Q�&���=���y�F�"�!�*i�Y��94�h��ג�瞼+]2:���Y>2��io�ܟ?���zl�%�{���&��T%>�9~s�A9�����zw��=�@��}�q��}Ϸs��t��η{Ο>:6��U�u��m<�׼�s�.G��yȯ��P���`Y6�bOƻ�Qԏ/<�ia4��@�ҿ��(b��f�:ΰ�����<<��7l��k����g�����J��9��2nF��[`0�׏g������|_S=%1�qR����2)rv(&Ay�[0&a�`�$W�KVz���<���*G������G߱�x���cn�M��ҫȯ�/�\�B����J���H�^RyfByTF=<?�����y� BcIe���$-U����J�z*W��:��D2�I%+r�/
)P�o/2�a	��{<l����D&x��]�'����msωez��ù��K+Mڳȵ�B&`E�1zτ��@F$D �oJR��9�0�Dih��ñ�U�WdQa�PTz��&�$9 GԐOi��G��r�|{/���fb�!�����)1�f,+Iz��c��X�G�Ֆ!�aL�p[-�@�5����(�3�3�=��8���LʌԦi&¦�'=_U�J$�s��^;׫�8&%��-p.����1��6c8 hnT��-^���O��������}�;�9�������z�N�O�/tY�`�A�b�̇�c@��^"��f��������Y]�������O�8�{�M/>Z��d&��n9v��o4��X��3�[70t�Ch���t�D��sv31���ӳ����C��P��	�d|En8pn�".�6Of�l�3��4���A�6OP��A�DE�8�^@ݲ>���h���(���$�Na��כ�e|�gf�26PpAܗn�;��v�� �+PDL[�ְ\z2��pn��?���1���{_a��MK�Q�8�p>ɤ�2׸8l��3�A�'[!���6ʦ֖C��pw >�A �w5��$���b;׋�p|bX"#	Q4.9V�C��Fc�1�6��Xәn�q��X^6P~�,�_b�ڢ<'G<7��G�]��Kc����ß��}&	����l��Ƭxo���eq�[��h-� -�l��Y��b���v> ��w������$��N9����Rp���"b-�7��'h;���9+�8�8c7��0@��^�a>"���5����O�����e��#�o;Yv��殃��h{n���#�h�腭K�6���	�~�����/��x��w��yOu�oI�x��xgo%w�^Z�O�#uy���Y0`��S�C����0��(�k���a��3K�p��3��8��\��`� �-we��Ll)�X/�	z�hV' ���@ ���BN;[�E�KMSJ��'���;"� Ѣ�LA�S�
����g���6xW9�> �8�#9��MD!��ٱ�4����x_np��j[���na���d�-�����0�H"�5LD0F��BY_��]��V�lh�=��p��o#�5H/T��Ձ�i��Yr��u�ow��8��5R2�{���W\�{�Ė#ޗ}Db�m��N�u�;��D0�6��I���y���x�t�i�����1g��71,�}��=���E��j&b\ӧ@�'w_�'��tP�/;�6��2Ҳ��[��#(�aPV9��ܶ��;h��%�}Ǯx�k��7��0Q���ū�U��a�A��]��v����$-V8q���`�z.ɴ1�HX��ZA��u�^�n��������!{k��tZ2���8�^.c��Ȗٺ����&�f�����z$���W����!�J�,lfzٞE�����Up����vߟ��em���my����ɸ�]����^��˵Ӈ�W�����ߣ���$�l!���d��-�����O�0�-�;&�m����(}T�����>���<�_B9���������Ƴcz)��CD���A5(H"ڈ^5M��P�@�=́q0 �D��ER�>X��{�D�]���c�s��.d�ERT���2�>���ï˶kk��^\8I��e�	�d��-���+᎟8an�r
�����ց�Ic$�T�4P � *���Q��ݾ��tY���ix��:/M�A�dA���S"5L]51jmmc�=��A%��j-���rS5GB=��v��uk��nK�F뛴����^mY���̰
mz�"����_#-�F��x��60��:|�Z����4F�v�}v�C��f�A5a����[��?X9{V��2&���ü$�/:���ݬ����f�^���WW����\���	�ɱ:�n���R&�Žc�fC�>�\�����RX����߮s�M��T�ԦjF��U3Pl	���ם}�u�6�{�~��Ά����|1��-�	�`�F��7:���Ӊ��� ���(T�x��Xamdݱ��Gz�����KL�6�&��"��5L��j�z�`�=휩����}n�8h��gPc ��Ay\N�b��D>���/9EEA��-���Э�U��1��05�9v�M���S3�.݈���p�h7X7KqW�a>h��p9 �1�h�DU!�{���zЩʃ��>�y�c�4BiM6T�4�n���mh��v�Y���(}ւ"��)��/x�loT��Ii����i�����P���" 9�SAh����U��ĺb0#J ��W5�y�m�1�c�s�%͔`�@=E7R�ʪ᯾�l>�h����d&��)���:q��]�v��`��h����<û��p>��vܦ�rX��C]�h���A����ns��t�<t�؏mP̪�5x��{����LƆ��d�O�0���CA��pl�@.� �d�7\�UL>��c	���@m����f�3�Z_d�΋�m���S�����n;/Q�dA��"�&�0©<h��1،R����%��������c�o�>.l��AT������m��٭�'�!�~/�vrM��ra9�f\xP���9�vx��B)8wE�wvw]�'��G��@��d��pm��*�a��ᅨpA�p�E6l5=�0�A~^�aU *�5LRF���]�w,¦�6��^@f��ީi~��</��A�d+����x�1�lM�ڈ)�86�F� A�����-L�R��cž���jk��6L��l=��A����A3��c E��4ō촷j��r�7�� �3q��۽��2^3F3q�/hB�_�h���]Р�o-(�L�*��<��q�US��~����:~g����zl���^5�+gǖ)�>^�6��=�|��-jVjMef�F`(|�0v �0�p �0@�T�"��5��c/Ř�6��ח�f�3�U�Zc���%���7K��2 ��x#pz'�<����[5-o����,��n-�.�Sr���h*M���:t�1t������r��#T�x�-�*�Έy�;�cC�����L��I���@ Fbx�k (T�>5�vۧх��82�1�0C�	�dMކ��hp�y�[���x�1�F���ơ�s��$���)U^^&i�Rɼsy�MԶ���2KK�6��1�^ ���SG�&���7�� W�Om�{.` Ġ��dAH/,��/��^t��s=�~�x�|��aMI�+ ��/� �L��A� D��k��Xq�$��X4�d�΋]�����n^�`bT�U!��Ǝ/�<y�T
��"�b�u;J{�%�2��sm���}�hȹ�,n�^)��R�;/���x�ry���,�l�����n�0�	�������J ��Q�5K5+6iL�#'GׯG�4!�5	�v���ݳ�2���\�ϋ���.ݹ�SVhM�aqu�qtf�32�cQ�%Ȕ\�쉫����_q]�xI3ո�u��^��6F랞Br��Z�U�`⫬�l�'=u��
:�vƎ�ۥW�c�qmg�7����\!�Ч���VB���E�is(���\]c��J��.z�˭�c�=�j�-��c=�hun��}���Z^�I��z�:��1v]�}u�M�\k�rڴ��B% Ɋt]�ۼ���>"����`��Ax���k�z�Fɔ�/M�2��4�p[sY A5L��T��`!�DKc�ŀd7���M���3�#��z߇�>=��R�"����\�<�Cc�	�e�3U0@�2�T�s"ґ��3��D 8ڼ+kCZ2�s���r A�"*�x�*�^"�x ���`�Y�ޤ��k����n��ު�Q�T��m�@4̍��R���
N�f�	7��>5�=Uj� A�@U3R9�42��hp,G8uWy��<��.�g�o���AT��A�g����7߿}x�稘sr)��q�k��)�5�0�-�Fp��3��Z�l�[f����>|��w�2 ���DT��fﴮ�hp�y��7 �H���c/m��[a9l8��H�k�-m�M�,�d�N{]3����D���8^=��;f����:5Oi��{vf��K��byK���yUϢYL��*�������>�� ����Y�fC�X��b�^^'1�Ͼ��oUB��*_����^>�oU5��dׂ���m���P���y�p.l�Dv��w<Գ�S���sa�fu�F9����"��,U:4@`k���Y\f9L��o���M$ ����w�Wo3Z2�3�>�a����t�ô,���<h�2�AN�F��^iz��7�+�K@��SqoV.��U=%K�6� �2�ڈ@�DT�>wc`p���v�����iV�K��P�멷��N�����<�v"�Vl���e>�=猼O���{=�}T���h��3:�#��y_ �P~,_�����FZ�^"�yx�7��d�}��`\� A���q]��hh�x��� ���Hj�t̪ ;$�z�R��K�t�S6ӈ��h��u3���N��V�vG=�	���1��[���W�%�&w�աn�^�����+a������^~w���x���hY��#3J�*�CeF�Kj�_o����R�jYOA�6�x�S A�^CƩ���H���@�UU��F9ߕ����AxְU ��]���ο\'����퀼�־��M�фv//U���S A�o*��j��.2�ذA�d��v���mo���!�^ �j�"HK!9�:vk��ݬ�R僃y�y��<m�6�9���D��8��n��[�e���=��'a� ���"��T���ϝ�R�jYN����C�d
�S�8�G6��:��s A5M����A��髻u5k�	]��/�&�h��3;�ap��xŰ^��wӮq�hY�}���� O2 ��T�}T�ƴs>扒���z��2�3�3p��`�AT��A*�@��-h6�q#�\�<A�A�ުo@�����~�����n ��D ���h�����u�
��Ɩ�X��jaK3�[�*)�!�6h��@g�����ɺb>���n�_�HY�/���/��͞�N׹��e{��ԙ��-a3P�J�Tf�w�w��>z�0�����A1lh j�TlG�C����]��V�1�壄w��p,Ё�H C�ySQf'�dD<��(��|�Gn�g]eH���]��Y�Gh򘄵h��L,��K��ݝ�ƶd2M� j��T�+7٬�����-�8an��ِ�bmW�Z���0pA�A�
U0PM:4PVcd�f����*Ί�.�E�����f�<�M�Q�/��@�7,�>v�5L�Q�e���TM�8숓����x�*�@��@�����̔�T
b'��F�\p@���ER0�^^>�7m��~7�Z���x`��0��@�j�yq��e���33���{!�":�G��<�r��6��9�U�!�>��U8�|�f�wx�h!٥�ܪ_��(��ۈ%�[QƩ��c�� U�quI��ૅtӏ��j���Q���x�4������^-_E��,��Eo��,����p��7��j�=��I�l�rYox��5=�"�zz��ߠ~�&=U��s�{�6&P5x{�|s�.巉��={�^B�'x��P��)��D&���۬.����=U#x�4�y�=�/=����)����e��=�	�S$m��d���9L�8z�#R���`z����%.�n݋~|s��>�o,1Oi��&�ungtE���^;����o���v����4o�����}��}i�_\�c&�������۱9��W���\:�T��q����l�{�\�nR��x袸6\�٢v��<��x_V��
�cP�.c���ү�ܸ�Kf=�C�������r���/%��Q�{Ɩ��U@�{�n��: "�=p����nN�wZ��yw��}`s.�Ը��g\�<���q&��X��H�_� X���?x��q�I�A����D�eix��TU\Vx�|��7���$c��9'�㹁�ך��y���{pt�ra�����'�6p����Mgޚ��o��=G�[�}Ozz�c��[��:y��W2xu��qc$���v�n��8l�E�U�5�#8P)��n���
�|���v�@Pչ�=��oy�R��{x��o5F��{ư;�_c�:R��*���D�Y=rd�Pk����>gI[x]���1gz{�JÁYR�_7̞��?�|/9�V�ȟ��޳Fv�jǷ�L�X��M)�@��J��Ai]���@ n&sttj[�5��	�Gʾ����$<#��i�#������y�! p�Z�8'�����[c;k/<|���AK������yGژ�XO{"@���B�k��� H�2�1`��z��m��Ȃ����<���z�C�ܭϻ�!�E���;J�H�"3r���#tK±�Uuu��O�����(ҝt���D���ќ���D{]m�(�=39���v������Ͷ��Ͷ�ٲ��R���"����_hPuĢ������ȯfQT{ey�ʊ�Ip��(�"(��d��B�Br��(���]O/(��ٙG��g��D����*k�TyQDQ���\��<��*�+SƂ_k�hG�PxDW�dJ�A��z4�,(�<����<�ܜ��3��`�)�5=^VA�T��$��(���B���GR�ȳ�"�g�U䢝�DE��*� P)B�<l�ʄ�E^���=�UA$:���b뉜����+Cn ��L�n��7\{lW���U��eLMM��B�׬�A�m05�[P�f�LGA�:��L�Ön�8���m����f.�wi�\���T7eM�汈�69��.&�̩�]����',o[��ymsɽ�6�.����t�Ŧ���դ 
B��X�V�LîVimc-ذ�]2�e��%�hm/���R]�ksu��"O=��5Ƈ�%��lu�Yݰ7ny��\����S�lM�����$�����Zl����ưuBf4�6��%4Y���`��[d�=V[{g�d�)��c��;���㵈��f���\ �[q#y<Z9J�!3����Im��6'��jnŋuw,n*�p�ta-&6Á�]Ɖ��ŗ�W�y�6�m�����^d��MM�;(��&�*#��u�e�1i��n�ŗb\�J/<B@�66�;��ۭ�WCJ\�зYeV3-]ni3��Ǩp�k�4k��7�E:�Q�:h��ט�b����@��\����l#�ܧ	�H]hp;/\��ێX�ŗF�*���;�͢���ַ�#�mf}"�-�GM�pg/-�e�r�Bl�ȊV�
���Aa����[\��8�V�{Z�v�8�����$5�:�x��]��h,X��#�c�a{ķ0���`.�5���p�����׋�@OW5L�pvjg����<�/�qoK`�1�,r�ژ��6nWv[e����J�]q-8�[�����s�,ޓ1c���g9��<�n�2{VŰbsK���o6*L]��2˘r�k�ㅝ�kz�u��=���m��:�O/Gm�x� i��M)�[	�&kt�a��[�mt�Q[8W��tc�uu��Oh�K׫t�:[官e�c6,�yA4iƩ��QJi[�����,�]���qU�D��Y�a�&N{q�e�i5�Z�`on]
g��z���3�0C���k���K����Z\fk�,lݭ5^j����g���}83*�3J�)��#B r�y��~������(M�5�r�L�6�p���2l�8&m�#s6r�u���M�,��ɲDpX��n�K0;X��$�ͺ�f��z.wJL��H�t��!z���,�rG�0�EGb�Ñ���ݒug;i6ݻy��J�-ד�4��E�Z`��eQ�ܒ��eX2�`�]1J���Mq����ҙ���l7�b{lݚ&�&���b
5���~N�}~��q��\+$�Xk5����E�/"�:�]qlζ1չ�g��,��I��P�>�a\N+mc3�壄w�9���C�(�Df ���5L�TȊC���YT������	�d��v���l�Ȍᅻ������f�D
�	��1�M�
�a���p�.�"*�^(R�)o~�΃ma�i8���v�_n�(��ۈ&1� �k#��5�"	�e�,��G*����A�K�U0Adu+\�f'y٣�w�8 K�+�5�Ӯ���s<�<V���x�a@�SO�>5��md��ݵ�G5qv��<�F��L��-�6�ḧ�[���4���CZ��1� �랰�H��02&m��:dC�X�NX ���Z}9��n�5ۗngg!�q���4��.��?{�g�=�b���*��K۳�ۼ�vn�<h��m�t��sF�Y�A�^G-��@��DT���kc�2�0�I
���o�zg7{c,v�o�[ϛl�������!�PE�z}w�����Mo���#�A&�����9����<�+w�=|o㞳�_VVh�A��f��6��/�]���}��e��斉��3O�FrF0q��c#3bNV����j,�}����2 ��D���T�MS ��pG;[L�x[!�#8c7x�d0@�x��`�"��U$)�D�O[WW^�0��BH7x�T���[�yT��x��ہ�ȅQ�݇���[��D�@4�5L�R�S
�c�N��2r,E�-խ����3���o�8 A���a ���|*��m��H�o]��܆��Xكf�jI�Ndg^����l�ƴ2����V�gM�RXA�#�y�@�S ������l�|���E@�#n�����*�AN��l��&�	�De �FR�6u���OM�Q"�ٸ���^)yT��.vc���M���X��ת�G�"�	�9�wd[WO��e�lͶ�n:��5�)%A�	���Oup�/�L3E�}/���Lү��{sC܂��u�+.�륾>>w�u��^�,���f��j���dx������Ϯ�u�����}u�w�>\ c"Zvުo@ ����	�ݫ�T�g���`d/ z�5L�o����l��|�ь��")�NVy�W�Cz�{H"*�	��0^:z��*�;AGX�,����Y5�x�OU�h�]l�*n �/ j�x�j�E#�:�v��?3��ňZM*�ҕ��\h��/mz��n=L�4�O1T[��m����~����R�Ya�� � �oKV?4�N�r3�;�,��Dv�y�y` ��.�K��2��S Eֵh�~f~���E�`{� �o4���,�����|��,ŀ��a�nz�v���D�@��U �K�ƚ����-Ք�lu-}wgMT��%�+����2 ��G�M�j�Xaf�0��ʱ�A�u��9�����x8W��6Z����t�)n���	seZ.��L�6R��l���lX��)�V]��U9�ν5?sWyw�(�b=�,˻wJ𘖛�"U
�c)��U���}5��3U��ضF�66�_n�O}>����������S/|0�}v��q ��r��Bb�3œ&���u��t��C����p1�f0F� �N/���aa�����>{��2䌵��
�f��]�������sZݧ��KffL�:x �r�>W� ER�SQ��=��z���痖lN��x�s/HF��>�d�D#T�*�j����.p�A� ْՏ�f'OZ����,8ph8\k@��h50���[���o���Z �2� �R`MS"�SODi�t�E�Ɏs:���,��sz1� ���Ex�*�@���@xj,�YE��$n�^#q/SQ��=��zp��f�T2!DX���ȷ�"�!�YϞ�(�ST�<h�ގ=q�s����n�63���^�|1#z��E��%͔D�Ux�Q�v꒕�qȮ�	ۋA���yOV^á��w�e�#E>�Ѹ�T^}L�\u�<�xj�����3�`E�5�t��~����~��w�3��3�Z��2�{3D��|w�"p"w'"=��l�2[>9���:�m�����ܜ&���0d�$v�a�Ӵ̻,� D���-�#�t�#@��#͖K,5nqZm��[��ΓP5#7*�1��m�M45�S-�!����XIV��;�mͺ�Q�:���]���t�v�vc��9&�TfG�\m�g.�Fv�:,�swM�ܡ��]sW�k�x=�K�t��	mxBm���]�/v:�`�"<np:;��}�g�I��\X�2;����u�a�v�C�6�^]2�E�mv������0����{��^5L���Xrt�?7YK�#/�3y�u�:�SL��D���U ��^@��E���N�p�M%����Ӝ:�����W[4��f�����kN/�2�Ȍ�Dn�/@�AT� ����y�e���R��
D<���?y�0%S8>E ��o	���T�IV�\��D�of�u����\o�9�˓��f���+9��;U����������D.� A�`�]����O�I��CG
l�c:�������S����n�L�E�T�}Tƣ�`wm�����D[$��̼Hwp��+G1уue�%w6�K�d��E9�.�����?g����5� � �j�"*�&̓v�Ď�\��Ĭ�s��6*%���"�@����^@�2���v��;�m�q��m��U��F�I[�"��>�%�7o\�O#���x9�)z�!=�HG�_�(-��Y,�U4�V��`�nj���wkRz��Uji^_ 3���>�> �Lk1�l���i���ᔼ��6���_Y ���GYO�>]��n ��@��A�71T���3nm�,�o?� �
�ESyxU/JO�����+{��L��zj��VD�W[7��鼁M��j�|j�T��_V���y�
S����E�
Ƭ�9�&�č�\���{`�E]ok�U�r<�v��5L�&�� � *��E�6=D�U��o�ǲ�p��i���_f��"b�z�͋�w�Բ2��_�̦�9��z�k+)�N��1�{<��]������X˱������`{�� ��b!�/���9���n�lKEm�y��V��xB�ۈ5K��2 ��@T�@�0C�5�l,��A�r���n�7o�^'��WA~�߻����S�ˎ����`
W���/A�dA�^@�D����=��8�a��0��7�w}�����\��my���6v�S%�O�,��D�[};>�Ļ5H���cC_�ώ�g�>~]���<u�=�o��f�&�5Y��Z�ړ,�h��x���~�G�O�|1�� ��`�!�p.�E�E���=d�gT�Y���E�yx�%�T����8?V�;̴V�7K� F^[!�����/�� �o/�P`i���������:42@�Sr��=ԧ^7�|%� ͠�H����~~��:�	�%��1���vm���Me�C5�+�ps�,;:��2Φ���r�i�D�ύ�3-@����,� �����/�>e��oTuk�f�)q�6Y�����AU *�>�.*�R�RS5�FJ����Ӝ�m��fZ*�n ����%������~�=I�=rY;9|�/f�8�G�RѢ�L*����zm�3��1WKj!F��6P �6�	�Sy
j!K������l��oX֢��� �3Y�ӹǤ޼:|�х�0&�����([�f�Lnz�|��e=y~���?��uy�
�q6&���q���RX�
ӽG'�2������D��\f/y����>>~3�[ϵ�,ɘf���F0�{{����o�}��>{��yݳϞ���Sgx�B�������B5�3��]o6�2�]L���h!�Dj�����-;���{WA�[T�ĤC�3?�v�!a	�GRf��T:��v���+�w�??�0 ���H=��hׁ�.�;v�b����Q
;�L2�a��n��,k���|)�O��`�N9tfƻ	� �2>�d��i��i�焟2�an�`A�`��5� �$3�Pt�;�#�Ax��$?��DT��H/Q�7�0�e��"r+��~���~�h��n���Y��o#T�paf�0ދ�]ݢ�dC�y㦊 � �6Z�𘍮��Q�z��.l�[��qp��0�����F��0�W��O�����iXu����-d��9��o���_f�}z�x@�z���7i��`����֭�S"�A/��|���������H;���z������eu�w"6"+�Ʒ���Ά��Hy�N�b0kW7���u�]w�f��2��$�����=� �Zmn��P���\���v[���Z�c��� �k���M�K^:�q�_��
|�5�:;A\v�휺"��#��F��[�Z3kV�Cn8ޜ`wOL�i�٠ʩ�mg�j�����o`\[���/Y�CGj�{��nwٝͲ��t�מ��ri�'>K�ÁƖ����wU��Y�-��0%�XmYv�#�k�	;h&�-���~�ߟ՘*�y]��6�:��f�2�e���:�ct�mub�7��w���X��}Z�Am��^@mV��/���ߦ+����S���-U�����@�jd�`*�@h�9��;L�g���� ��咭_	���n����<Ah"*�M�|C+Q�n��7l�AM�Sy����L��,n/Rr�e�%C;�_fx�`�A�z��n�"��A�
�B�b���o����Du7��R�̜��c��ͿL4WS7Aye�D<�_^7z)���a�>�P�J�`��T�5L�z�� �˥r5���;�\��� A��Tުo?u!�P���O��=B� �z�i+�][��#jͮ�/�soWS�pub�Wck-ct,��]���O���X5��a��zc A1����m�F�/F3q�۬jL�s�M��+���`E[�B�нT����7�黫E�<M�����]�pU�5��>�8��]~~.nB��3� ��*�^H����[��~;���z�������G��jl�5cY�f�6m�Q�뷼�竿_=�{c�����n�����������ꦼ���6�-"24o��0#q��<wX/f��RU �-K�k�C�+rq���^�;�\��/l M�M��yx�2=��lA��f�M�����V$�ղ�;�v���c	�/�3p>�`�h�ܞ���tp��T���ϐ>7l��L��	M�^����_��.�˴V�73���^F�� ���O�j�H�#k�H8,�Ĺ	˰,�v����[�-=H�f�k��d�pܿg���<f�|�T�5H+Y*���MT�=[�w��!m�s��&���#�H"���@U45M���}5~��D��_h�ޞ|�0�2�c7f�DU��S
C�Q� ؁|� ����'y��LIx�
��xZ��g��%�ѕ��n�ݣ��#���8Hħ�Rtww���;�]�튲��,���wC��g#n>{^L��~�>���wq��k`����;W�}�|�x����y�Y�Q3v�gt0�}��C������l_����~��<E�񇘗N�������r��}�۴{����.ʮ�,��x���jf�>��%÷��f�0�|s±��z�_�{1���~��� 9�3��w����nr��$���Rx������#�h(��	��n��s��k�o-��e�oo}]�<�;�"v@kN{��[(
�����C�W�w�\�k3+�y�����;�_��!��?-��n�=�\���.��{�ΣL�Q{^��������xtgwz'_}��*�t��a7��;|��F_L[�r_-^�YJ�K�X0�Jk�lX'�_0�O�;����!xܽ�n�_q�����y�vW��}����/��cr���3:�H����&x��=���ׅV��e;�f�-&N���*$�x#���kO%n�`&����n�~�=t��y��Hsh���j��}�מy�����_��$���7ٻ=��cXr?dsF�=T̘x{'ƞ��nW�E��z������ �'XO޽FU���h��S��r�a�;��9H��z>�>�U��B����u���Ivb� F�[����X	�{r�Op[���HG1/N�n����!��HƳ�V�Ui�H��^������NTu� �7~#��7��?{�H3 �b��\D�%OM.q�tz����Ȯ^��j�U'�I.	Z�G��(���L=+2�+1_8̊������O��E^TWD����G�yK��ȋ��t<�c�,�<CΥq��O�O���&��dI%UDi.�iʤʈ�Ȉڶ��&ZHʡ %��ؑ:�=OO�O���a�>afԬ���\ԓ<�\���<���ur����V��0�я���O���Y!xO��J���+�P̦��*����"���x����rd�EG�$(�^I�(����i<��+E�0d��af$yBE$G��E�jL�U��l��OL
�P�y\�(��	/ �"���R�J�;P�"�w"�9�{$�##R\2<:�rg��U[@�sQ(��MOT��.��+Đ�jrC�.�-6�L�q��E�J��L�����2�8$!*�;M��zP��V�S�Q���"�F]��I=F�G���{�6l�4f��6�ǯ>�_[���E��v��f��b�2�����L�@Û��*5�a ���["���.�j�i��k��Dw�� |^���)6��*t��|EZ{y��h>�d�o/�Bf�s�wQ-�JL��9C�z{&A���������x�*ӂ�5L"���\�v��	ې�:�6M�fs���X��Rq]�����<�!�9��	a͆˞��U�?��a��0�H�4Bؼ��y��]���]L�C�������֒�dA5L�j�A�`9KU6�^|�'Ӕ��ҭ^m���S���0�@Tc�T-��3����{��s��~"�U4���i�6�;�w���.s&A����p`|sX"Zƍ�*�"*�C��f|�7���5>BuD�ySQ
��wi�G���K�t�w� �2�!N�y�}�R|�I����n�͕��ˇ�y3zw�</|�;3�y�;�
��י;���;��;ǋ4-nv;{�����-����χ~z��{�5�Y�٦���R���ƾ�����^��(�`A�`�"��4h�٘��d��z$BAJ�T�tUV��K\�yWx Asex�����i�pT��ћg�,�!���-�Sf���
�5����ݹ�7=H4]��ܐt鋦���|A ��f *�<A �2������T�	�/�[��!�Tΰ�A�J�j� ©�&��k[�̆e���>"!���W�����*�A��-��� ���$]7�5My���6��{u���c"��5L<�l:K�
�d4ub��o�Z�{ʻ���x�&�M�^T� B�����e�7���v�]h
��/z���rhO�z1��Bf�@������ۮ�l���0@�x�`ԗ��"*�/T&1��Y��=��ѝ�ٝ�Q�7}%��Y�<2 �/ j�ꦶ��nl]U��ل�Ė,링)\f�m��Wn+n��+����o���@fs���������\��q����/��d��-#��ھ�ݷOofmf��j�ڶ.z�x����f␧@3��'GFy���]�۬�4���+˓�D���e��Q&l�V ۶���٢�lD���Q�
v�Ii�dK[��m0�m���N�R^�����c�WI�,����,��j�ȳ].@�c0�ݵ�;�3��4�˨�׉����tx��R&eIQp���˵�Ǔٯc8�w1d��)��u֨�oS� B
�m�_����{t�'./=�Ь�Z�uڱy#]M��70�Cn�q	ܷ�����!�������ͬ�5���g����J�����3�/z�^>�^�n�H>7l��Qy�0F�c{�%��Sj�x�ӹ4VF^�fq����W�L/���q݂��^�
��sDU �j���avB��k�{Qض��}L�AἽv��S Ei���휉�PF�Ɗ�a�"1�;���]����,�U�ђ�g�.�TÈg���܊������/�?,8m:>����fZf�|{�?X������go<��+#3F3{�kX"Z�S ��-���<���D��f�vx�E�<�����j�n���-+!��X�:���U�9wr8\�&� ��T/��{�ם��趾�}L��E�w٭��]�jv�A�r�3l�>5L�0�dA����Z��w���Ǵ;��� z>�.3	���؇{N�X����e�^
�O8ڻ����L]d5��M��{FŃ����}ZfY��kd9���y�ӹ����A�L���D֨�\�z_�`C� �M ���<ͻX��T�������)��{Yz��%�j����������\�u�W[��PR�38c7�Ƶ���z��}T�U:�(�Y#����,a$l�Pm7����J�x=��Z/����"&��>�s�g�Ʋ��"��S �T��`^���B2��I��3����+�®����|^�4�	�RBAoR^�yV���<,_��n��il��c��Y�u�g�q�֗������77���nft�갞4�P,rX0+�k�[H>�e�q�����!J���q���v���=cC �� ��`�AzA0~%��	 ܰ@��muli�l9�@�9M�^@OcU��5�r����S7x�^}V��S\�_c��ףL�z��m�0@ER�ER�ҞS����hlk�y���~${�n�=��E:�ft��违��f��מ��@`��l��<��F�*��Yq7-9�����s�罶j��36l�}�|���ۿ��oa{��)a�`�M ��Ax�����dE��c��;���F�j ���������q�����!J���q��a��,�_���>@������ f��ST�W6�j�i���zR�+[3���k��e�����@����`�Zo�g/{O��;�c��vu0�t۬R����������K�ī�=�5�K�س)ٴ6��`��`�j� AH&�6٘tm[�a{��)�:�3�2��^��L8sP^#�/U/#T�U4��o0�$Vy����^�y�{�9K�Y�1��A����v��CXD�/}�( F�@����I G�U/	��,��{�jڹM�e}L���^ ݯ j�x���L��|�y祅��A o�"R��f`ѕo��|���/l�^kD�L;����f��@��^f�p�ʖ�16*�!Ì��ĭ��7z�4��l��u?Ұ{#]�˻9��i��;�t�4Y:��]y�{mfa�m���/>;{g�^^�o#TȂj�ʩyx�2K�w}�_��A�-��WWcw\j�0�34c7�ްpA�N���*wǇ��+C
�^�h�6���V�
�GGh��0[��֝�J�/;���g�0�Z�@�@U7�U/,�7{�ζ�ye}L��*�͞��Y����f4|j��ݴ�ot��i��C,ۼOh�\�r7p����j�xc�����^�	���l��XN̛���, �2&Q/,l5Lcvt1�v��2�7�q�D�y���=A��@�.�F��UH(*��-:����I-�㘼�}T����v�s�Ĳ��n>xdE�Y1�c��H��'X	��Sy�z`��`��m1����]�� �d
�|n���/����=�r&� D��U/kV/j*5��#u���idX��h�|�DcKa@��lz�2K1�h�;x��~ɞ`g+��51n���M{�}��μ;���7|���|�^�L��5f�ޯ�D����\ScH�a���r[��m�2p�t����u���)�:8.z�(p�ϣb�����M�5�aS�[gV�qGTo���kL�pv˹�v�:�.��^ t����{v� yrqq�v�Y��Si��m�̳j-�G�.�&��f�����M燪��&x�9�a���!�K���|���.<e�x�nS�:�:�����j�n��ߣ�۷��}R+s�H�N�P�n��v���6��e�;Ck�î���������?~Y=�|�8�2⻴�u�%q��3p!�(�4���U0�i��T5L�SֻH�Q}�#Ӡ>�^#iz��fw��o7�����^nא5MP�{�[��p ��EBT�ERS�E�l�8�Ƿ���yrX47�0��AT��^F���P�ݳJ�Z�n�/�@��f�³F��v�8�y���L�D#C��1�5L�7h ER��������.���ԯ(��y��_=�\K+�f;{��^@�7�5M��:�-����<KU_c���L!'q���V�Y�ء psv�r^n�m��fg!'�����0iS�`w��>G����[������ֳNY�E밐A�"3[�U/#TȂj�9W)�P���HEK��쫱�!�$�8<_���A����������x����OM��ǻ|�௓�&�ߝ��]�=|>_z������33�x���~�D[/�W�77�|��1��3p �Ͱ@�.��0`ʢP;���mC�@��0
�Tފ�霖�oV;����2�.�Y_[7��/E����TȊ�Dc���x����v0���^�7s�v�[�Gq�~��ϖ�Gy�����2ˬa$g�T�����S/U2U7���6��I2�,�2�\;w���ǋ���m�����䕏�xHp��n�!j�
X3R�&bk6�1�[f75����j]�k�#����={���,"�U7�R��a����{-��e��K�w{ɹf�74x�&ב�d���M ��0B�wN�<�{K=H&̚�|��J;'9�-�G A|`�A�AT����l�k��LS5������2>�dA�R�������n۪��2Ռ��x�8���J����&K^]M�e��RϽ��*�����J*���ݢ��O_&=������*��������e����^�ff3L����^�����_?\���������`�@ U ��`F=�Ɖ������on�7[�4�3Efg�OS,�M�K�{k2���RW�=́ƹ�L�>5L�>�Ax���L�
���m^>DoS'��|��/G��M��M�s������߃�|Д��]�l�F���q.�v^�\�<����ä' ��gu�m���EcyT��,Z����;9���s'����1�����2�/�U{�ޠ��ES�*��>5L���j�P|�Z�ٝ������A�U�p�8�u0��ټ�.��0l�Cvz,6��EڙHa,�`�u��"���� ���Ú��O=�7I=l��p�� K�U �K���J�SI���2��cQ� �V��2�/Z�����1��3y�3[�;
4;�c�Cf[�1q��ظje-`�N�Z�o�Uh�{�i[����}9y���M�
��w"�������eL�Fv�H�d��p������>5L]���HT�}T�"��ߣ4^���"E�f���q�����q�22���o S6f#��v���e+a�4"��\�;:h�[5A#5��q*�#\-t-�vn���Z�$5����Al�2Z��K�vs6c��G2&�j�`+uxށT��j����2#�.k��:���y���!��{�h��1Ǽь�A1L�5k�L#��fmuQ�&�\F8^~`*�@"���V¹���Lg9�ۚg.ޙ_[7��e��� �2"���4���]p���,�����6���OL�y��l���	{`��׺�/�8�^ N�����5L�>z@�*�;_�.��SH��@���gZ���nxlg���A İ^ ��5L��a�6K�˸�͜��S�a��UFM�zŐ'3(V>S��&�f��7�XTbvٍ�������+�[�X^<�Z�b��[�({=�Er� B���D�t����og�0+)�\��l�q��6�w��Ş;��pEf�z（��>[�*�Pg/43f>{��иF�u�xL}E��xM���~�X��u�����[�;���oM��w��k��y]��s�*��&��lf�H|/{���O������5��&�p��4�]������ �r�o{��%��For����/�f>�a����f�o�N�;;_��v����KNgv�!�y��cG<Y9�5��}}�ǻH���z�S���|�x�'��s�bfG�rB�����Y;h� ��Z�Z�QǙ�Ohp#�A>��p�Ax ����y�;��������%�e
	w���;@��F�lg��ӿ:�-~��h��p�7f?z��j<�ӣj���y|��2<��(�.�tBz��0Oo�3�-X���N����.i�=�s{׷w=u\{���.���w�齶Mӆ���X��A��3}������k��$���u�vMOf��d�s2r;��{�����G�C_�CE�7W:�\3Ӈ�iG��rM�2/x�{�b���m�NEp��ڗ���2�3U�}7��q���3j����;�ţͨu{�\��_{Nv[��y�����g[��9�׳A[�}�.��\@����5�^�<7|{M�����n�''��A��BR�N0�Z��E�l3U��mc.-�Lxp3�n�{�@(H_����I���Z���%����l�<�y�@�i�߳��>!��\u"�9T��J
�5p���v%x�W���3rF?���������3I��"��hYD��%Z%�IA�����$��+���1�����	�*�r%tr�?Y)ҏj�(򂫋8�P���� �ZݸUy5q�|||z|'}IOD�c��ĵ@H���љT֣s�jT�")�W�И������~nD&T(�V�y皞S�izdQU��%h��;������a�b%D*��ͰL�T�(*:n��iDFy�C�g�EUV��H��44��IT �¢*��Mm��2
��
\�B�+�Q�#bk���(�)�eE�&�DQs*�+�<<�%t�ԅd��L��WH#0̳H��yP��@��"��/mf"���r�2�mx���ay�QTA`v�_���V6XC��a! X �'bx�Ͷ��;Qșk6ɮ5,ef�d�ч>�U8+����=	�ꬒq)V޶�n����Q��܇6��<aw����A�Bm�A�J��l/]x�b��h&�0�h�Ƶ�+Z�E��,��s-%x�]��Ze�dܡ��!�kr�)E��Q�Ua�hf��Y��;E�J�)[�a��ʻ�4�e�T���GX9Ǟq�$]E�GX�v+Ջm���LC�F���a�+��N��9�=Z�`��<q��5�1q"�y�eß.�n��Ys�'WV+��6�t:�q1��ܼ-�k��"�%��,E�wk3��msΛGa��Aj\L21)�pn��^X�6���
E��!RL�C:٥�ʠ�-�e34*q�:Ŧ%uM�a�e��F�Ь�eԮR,f���7Vry6��Ep`�����:�������.{n��Np�AzʩQ��B;n�4nl\�>�d�Y�q�Y�ƛGI�N�ۄ��܎4���W��j��hNɁ�gu����s�ɫ�b��j�h�L*�jg:,p ;k�=WK��z�+)��ݴ��	���Yi�D��8�^	��C*M++�t!��â@���%#KG-�M�r�&�Ux�,Y�u4�*ū+)�
�����m��Z	y��ڴ!��� 8�2!^�-�u�EaZ�\,|��Ź�v~9}�����6�43յqut�<qx*�X�מ�uOm�:��ݕ��3�u��i��Jv�����㜽#v��:����p\�s��W2�عg��>��GEϚsh�;���&�n4F�䦂�/c���X��t�r�9�Б׶�xt��L�4�6��3u6�v6�[��n�ʍ�=Ae�v�#/3�qn���wnuܘ�+�ѯm�]�N�z�e��[9��h3̺��l��p�1��KkcJ�c��==��om�;02���\�On��:���SRkmFS�]G	i�X���g����ÿ<q�N}y< ��f�M3 i�v�����nn;��%�F���t��K�ڱ!���ܢVL��y���{��;'B���&�����N��m�414��1�6k�:/v���ާ�U�nrK�V��65�ww���ٺ6����V�ta�#�Y�0�,��W"�K�{6ŕMV�C6;�T��A�6�lp�K���:��w������W��[�f˘(Z9�[���ֈ�1ζ�I�q�!���ݻڿ`�����&�^�o!�+w5oq�x�ze}l��`�ޝ�$oTΥ���"aT����-@����8�lٹk��0D�k�k�Ξ�t����n8/=�@�T�Uz�.�Ń91B��'9�e���^ ��=T�Ʃ�.��&���UJh�ӹ��k�c\gf��j�@�0DT��)��������>�A���xU/g���᳏5o)^�7/�!�ӥ�u�Q��l����l"���0DT�T��=�ሀU07P��ݎ�����d�l�綀d@`E$�z^^>�^�w3�˦7z��_�
�~��'��[��[u4u\�e�I�Kv�o=���8���;6��W]����~����t����Dj��o����nsn3�3qO`�Z&��"���h� ��a�[��5l�Nk'��*Y�ɓ����4#��e�ܼ��^zS���0��U��N�WJ�g@ay�z[�vZq�cd[fR�#�p�>�H}�'�n�-�=�۟�y�xJ�ٸ����FR���ȻPɵ�!�d�����l �T��`R��G�*OX�#��$�̛�|��q{`� � ��K�U/#T��F#�9�����  �iy	�-M���Y�ƽ޴W9�9�����^"����+�Iƶ��!� �T��K���U0^ U^�$��=y����n�j�|�Op�����2e7��d>5M1l_u?: �~��ĄK�\�I�l�'�7u�q����4�т���EC��5	��z"'� SA�A�V���^{&��%�.0��r��;��gM?\��A�@g7�U/+v���/Y���k(�M����["��q�ƽ޴R����	x`H#T�2-�9��*�@�A D��������Sx�1��طi�$������P̥��6lk����y�=9sR���w2�5�6>�TM[LŚ�E¼�R'Rb�5r@�> <cp��p�y��M}��1��)z��i��^"허�ޡ�O/��s0�X#��*�&�V��{&��%�gy��]#9��!'��V����5L�}T����<j�c�4���+cC��Z����z�K����vAh#T�x���{Щ�y?��?/�~�ƻ�GK��V� pmYL&#un;2���]@9t�`�')���rX".�#�ݷ��yv����/�i�_c7ӆ&e��}UmD2W�>�d �7��  �T��'D�m�Mj9�_E��,���.��^8<�Oc�LZ�@"1��O�h��ϰY[������P`��o*�S@>�k�˽��aY&m8Nj��%�g_f�	x`�3H/��T�U0���\$��C� 6ل A~A����k˸�����|�Op�������V�m�܂���
��.�ig=�߂���N��!ؑ����0��z��<.��!���ra��xv.FUMvS� �����5��LST�aUBr�3Ͽ	q�+�kV���"/��>T���R*�_Z~��z�?�S�``�=�� `դ�gy��c�m�Xێ��䱝�:y�=*��w���~8�^��V/ 5S8����/:�/w��]fp���oG�6熳uLg[
�� ����a5L"��$`�l*� �����5�wN�Sw��3 ���e *��#1�"��o<4 A�a�T����,
�Vxd��9Z��C!E�����O�/l�RT�^�@U4O�����-1;IM��dA5L��y���.�8b�c7x���<�u�9�$�H5l#9��I�`�@��p�UD�/�'���K��hnq������`���F���\U'��a���jޏ6n����_��U+c���w\����=5�[�T��;�:�:����Y�������~voG�~}��z`94Ā��,� ��<1��{w`hxy!�ٳ��>cE���������kن�l12`kA���rp�.&��t���ʌw'c�sd獉K���8�k����F��o�Hx��B0��s�{:�.ȼ���i�c؍�a1��I�u+mļ3s��V^�j⭀��5�lK���Ƹ�ժ�n������-����:�fe���7���������u��m��f;qa�N���R�؊0�f�$k��bڮn_^���<o�}���AT�R�x1��Tpx����P��r|׭��6��2�x���m ��@U0MD.W�Xw\t�=̈'���;M�o�鱢�c7x����5LՈO�+���A�HA����^ ���K�
��!�߹�Us��F0T����q	^�7D7�H
��T��U2�[0�\���X �e�`�A6n��i�1}=���b���.�����Ì����v/!��� �y��Sg`h[9{�"4W��!hosooZ2�鱢���&�A%�� ݠ��`� U �Z�=#8�����|������m���bۨD2F�jv1mn�ri�[$�����!��;�w�[Ѭ0�7Q���q�7�s�ν�3��f��0E�]�$񁏯SY�sYU@NES"/L��zffƼt��P6�r��Y,(�suY��="�$콺�f���{����o�V��g�r�-��7�{W@�X��=��Hu�}� �����O�맱FdL8��U �EE�C7�1�Do ��R�5M���5�է��N���\S�u�bj[t��|1��� �*���@ � �N�YgKm?P2�@ 
��s%�*��=f�u�\�]�%}��A�jY F>X��\B������ ��DU2j�/ERƩ���[�ȺR��3׬������ި�q����� ©/
��`�ή��ة�@��D�҂-v̺�q�#Vn��k)vܖ]��X�0v�ֹ�65]��h�́�a�!n *��2�6��v�5.�lh�����6�[�,��"e�q�A�M ��K�L�[���u-�#ǁ�u�м��Y��nU]�����@�E�����+^�^;���?�-�v�8!�@�0^(8j�<�47ih��<�<���r��<��*n�1�T֠|,��x(w��{}w�tyW�>�� �5tY_�r�xW��"a-�cG�A��N�xwd��g4f8��@����H/U//Xk�pB�����\ޑ2���/A�na�v�i����E��n ��0�m�qu5!,��@հ@j��E�	7lh ES���WN63��y��s7[��E?AW����� �/#Tȇ�M��geo�;A$"\&fܙ��.���l����K�X�&���� ��F�,ź?#�D�
B �z��j�;ݩ^��6����1pA��5�'���0��^#yyz���5L�d4�⇍g_f��[�/���i��Q���-�6�+>ҝ���4E����P�H�8`�Y��l��"� �5�SU �ER�B-,n���禔�V�&�*��n� �P�E��5L���v��i<@�'�0���H oX >�R5��W�c���sFc�]�����7�π���\q$E�=�Q�f�s(�T�n�T廝����"���Z�|e�;<9�)���vI�}����{:�py�����l'��̷9�����\�T�&;Q,a��> �A�(��"�o^��O�Z~V��J[ �����*P�Nf�7�M�X�/�3q�0DM �5L��s�S}��B���̙â�\����⃬�B��qm�m��uk��膣�e�wѣk���=,�A*�ƩyokZ���v��������\��1G3�l �E//�Dq�o]��|n�"����� �3&��K3KG{���1r�0@}T�"��+�6�E�:��7���ުoG��e��SF��JI잭/W~����SkSeV&���A/"i����8.�r'�X��؝�� Z�N���I7�\�.縪��ss؛��S"랝d��W��Y�d}v˃�r��>�^�`h]٣"�U w��f�g�qW�c1�.@��0^ �nv���{��$�ᷰ�8�P��z���&�ۚ{������d�W��I�x���D�{���^�^��ϱ��)b�YBj��pU��f�p��M4={�U��W,eWMn��q�Ǯ:A�tfm�6�s���$�Y�B���*KF�XK�ҳ]3f�
�m�&qv�2�͈::�b:�%���77h�Ǒ��{Dѹ@��blŲ-�ʒ2q6vՓ&��vt@�Q�қ;f�`(�F1,5%l�F���+d֏]k!���X��f�Żj��㓎n�k��ZC��&�\[���~|�����U���l)]F�h�un�c�Ř�e��Cf�a,�۳�|{�7���^@�2 ��B��;{��Y��M��og�"M��>-a��q� ��H	�`#6)+)`��$q��+׭�ݡ����UK�9�8���"���5L�+��f�����V�L�ES�T�p^��i�Mf�֚�H�}s{��b��/l�H"*��^B,v��2��\���7�ܭ�2X
��	�ka�z�Mt�mV7���,jX M��m��p^7�#��U%��Z�ERj7ǚ0�o�yb��ٽ�W\UK��\q���D] *��3)�u>����'��j:�������{rp�^��$� �ݠ=��Tm�깹~ϳ�~7�)�,^��l"�[�ifg�77�_1�.A��������ks�'���a�GrƩy	i���e�$6W�Q;��ϖ��D��kP/&/�D�1�2�6'u*b�DX:��hla�W^]�ޒD֖���)���M�>�@$��x|�����_^�7қ�����q7A�`�A�A���v6#WU�嶃�#�y�T�<ER�a��Z�!/�p9s�=Mer�wR��Wc7|f[��TރTȊ��O[��ʛL��aB�l�5c ����u����/�� }a��"���e�l6tX!���k�ݲvȂ*��5M�)��D>;����yeˉ�ܓ�.�5���c7�����`���ZUk�n��������P�q�0�Kn�8ԱY��VW���S�n,����h�Mn���,_��?~Y`*����R�i����닩z\+��Ʈ\���%�φ>?/����iX2Ҿ���I{9Ժݔ{/��z�q܌����s>c�\%� ��EUlKn�`0h�U������A;��LS	M&�1/�̘�p�X�	�uJ�Òh�]U��� ���lCעeyzf�۔�������nn���(l7��.�ڝ�P^�ϫBvW�3^�;;R���\�f�2�7$p�c�a�p�z���������O]�}C9�x�G��5<�8mѦu�{uwo�yû��ev��.�y��{�N	x�J�oʮ��wurA��3���{��n���"���q��o[_�E1��{�*�`؟�{��}<�x�'�����|a��ٞ��,W�+	h��<���[ؼ���g{��@߄4Uץ� ����褺��]k��q�W�;�զ���4o�<qJY��\[�oq�jf������k�)*�_�En�Y��96o,���2�Eٵ&����YbK[�o�]:,��n���~-��פ��#�h���AE��	�=���{v��#�� ��8�g�o�7�KۣP����/d���(�νyy�?�ۻ�2�T���?J���=�����@P�Ԟ�F���\V��;�|G	�=�7��ͽ$�f?&,>[�	wO�����;u�vx��'�?"��w��E{��#�{�.>�`c����rwSˏ��{���se����#Oޤ���'_i�M>�n��a\���9��LT���x�����z�7��t>:�ZB� }�?)�^j��ev73���R���*i����a�VMc��C5n���_���k(�_��*�	��=����� x��6R1�\ӭ�uן��S�|�����z��0| D����ߖ���B�<����C�/<�f��[0؝�d�U�^���1������	&@����R��<�����yJ���j����Ǉ����<��WH�"�}A$)����TJ�W���Y/��������{|�W!��W�%.%QJ�DHa�ɰ����xa<>>>>^Q~�iF���X���3*�����I���PJf-�U^2���'���[�)B��U�$�
�	�`Ek`F(^D�ↇ�"<8!K"]9�^G\C���K�"�gh��hY�U�%2J�TTW����2u�b�P^�3�^�N���QTG�T�bLA(�)Iխ�z5�#�
�Ĩ���<��"��1���(���*������7}�����ӏg���h�O_?[|��,ts���U\1��/,H#T�T�hav�U����n�İ�C�:����݃l�k�뉹������A�oWLl�lM��k��>7�A��oU4 A5L�AH/���_;郸,=����k��k��g�q����  U �Iz���*2�C����F֑�H�nSh�����)	��Ռ�e�T�3b��GkuZ��Aa��>�A�M ��P�r�k���t?N[*���#g*�1��0@�*�G1�T��K�T�6��]ը���5>�/kӍ��6�v�������]��A�A�yxU3n�y?5NU$9��d��oA�`��S>�A[���ƃ����s+��p/l�TށT��P
4��0��o}M���[I�66\���жr�]h�n��9-}��Z��\[sp���8�l�)�g�S6#��Axq{�w�r�n�K�;\<}:�����4�SVAe�>��7V�0��;���U�˳FTL���1�����t>1��#��ASz�4�x��֧O��s�O5��2�B4���ۋ�����op7L��7h
���7Oy{Z��kR;,(�Ap��#z{vЫ��d�s�\�m���.[\l��B��pT��e�����H!˸�Ɔ��1}����&��X��I�j�DM!��*����l�H��U[!��fm�ń�=��~]9l�xc7	�`�AT��sz��X����õ���T�U �T�`��d!I��٩�#�Ϫ�4WnnY���T�|j�T�n#�'��_s	"9�5�<�R
�x������s*��� ���m�9��ix���S }TȂ*�`P5M(�WE;���8��Ok��g���es��L0@��aT��T�N�ӗ9���|�\@���Ub��b�A@Q��VI��VuӬU���2�wd|�|}��Q<G�����]Ӓ��{{�jᢆ�a�����g��VЍ;���<�o�m��ei���]�:��'f=�Ṭ.ݤ���)��N�vn9�`��WC<]e�]Z�zmL�]�Z�睺��SGM�k������z�L1F��7t�qi[�W@�X��X�m�e3�	[z���x�[;�7^űr�z�V�G���7W�9s�W����3�������d�.l����ffq�E����ح�b1٥�gh_��h>���eҦv/#nQF$ɻYveÂ�N�ȣi��=��DU;�ݔ�������n22�Q��*����=���ީ�q��DEV�מ�{�����ֲ���d&��T�<}T�@���4�qk�S�4�7�A�AoG5�`KxL_g2�p�Á{a���@��U��Vz����5�9�C A�@U4 �)�L�s�ͦ��ӹ����l�xc7 E�j����p桂�LL>�"�hL��<[�]x�v���4Wn�u�oR�F��q@��dMc�G*�P��q3#�w��ȂS!a��8>�`�0av���U�8���K��l{Лx�_g2�p��X.hv�4�M7����������>��a�&�c}L �5�Sn++	i!�y�Q&\�q��AL�h�������4�{�z�TȂj�}&uۻK��M�s�����Ǳ���x�;PG5� ��"�/U0@�{���mi&�����I7�Ѣ*���O�J;<Wa�	A�a��։�2:o�}L�v[����,W?��K�ر�56
fy8�5/e�}� 1�_%��^�
�t㮻z��5���c"�^^5M٢�7���^����	:��&��ݷ�U
���"�1|��s'���b�9�a�8=�zg�B���z�e���t��E�fw9#��'݈P!�6���1��"ʹ��&o#/r�5�k�Mm�rm�*��T/UPF���<	�s�/���q�U��1�h_ �ީ�N��9��ǩ�I���hjv�-0ֆ�y�qe�74<ݻ@v:,̙ٙ�gd��9wz�}UQ��\���旽�eXs���^'	��"[���@U5U78w�;�v�[�i�!�y�r9ϸ����@�7��UUf9���t�s�ޡԼ2�=ڧj���6�v ;�ĜJ�!��v���Y��O$��-p҇�]�=��N��x��r��0�ޑ�dݢZ���ly�0H#��e��U��ch՟���T��T�MpM�Ƈ�C��n
f��2"Z�W���s+�c˚^�9�a��u+5��2��oyef����ۥ�l�jjmC�{4���v7Z���ՄUTUV_y��ֻk��/����N��"ӳ��N������3��絗�tЎ.�,��~��S��oU7��{�h��me]j�:�Y�6;���v��l���	�^�`*�o���ѝ��(�	w܀�A�W�Ǘ4�vs*����A뺭N�(ݵ(��e��^ayw��Sz���ިA�UR��U��w�Z�aM���骪�,]�R�ިi[���V���th��le]i�қ����]����b�
��}�=��{q�|�����Ł�:W�ד%�����x{��w��, )�Pŏ���!��ۂ�In��Z�������.�}v޻j�;Y��l:��-2��ԛe��9�WK���LU[�Z-�~O����E>�xq��d]��]�ٯ\�جhە��;�$���E�wgto|��_".ׅ�0�M��ö3�s"��j�-��`������Sz��U/s�哧8�r�����!�4wa�*��WM5Y��z痪���$��>?gG��p����t�n\��j4"�;-�ke	��8�Ü�UUN�T�����3�ܽE��?/n���aқy߇l�!j�pzjJ^�.Y9ӃZ�a5�Ռ�R*�Ǫ�kr'6m6�"{C�'ѣr�x�u�Uʪ��+a�UM�U/�J}���2��v�ʗu'����A��\�`�P�H�/�C�s6g4�jS�y��dېf�Y��1�٢c��yΌ�����A_g���s��< F��e����0�������4&y#���+��^��|����ѓ�\-�]q�{<;�:8�;^�"ǧOS`۷l�å[����,%���f���[t��<TmIn�DR��9��01.	��[V�]��b��u�ۤU�}'۷I	� 瞲#�m��St�9�f�`�[��M��:�b�fc��L�k�'X����9�������"�~3��P��1AsR:Ju��O45<v˦ʁR%�Մ��Kp����}�m��O������R����>�P�e��y�;�5��UK�.ׅ�yyt�y
Y�b����M���vw�uG�=7��UT\�_7��*E.�e�zj��UZ'V��!��|i��U��Э�sʩ�����]Jh����h������L�Y�x�+j��>�,��P'TCo�UM�𪪬;}^Ѱ��P�-6S�a��B���ꪢ���#ch�f��8L��4[eՋ�WLYu%�SwZ����18�1ծ�-��}��m�S!UO|8W[n��|�r�B�B��<պ��^�a�����`�ݎ�R�jOU��kr����\l��h�زp����Q�A�w�EP��
��v
���n���_�I���]���
��p��y3�ƹ�G���㡛T0Y2���׭�UK�L*�����"_;�4�Z�66��z���.�^��T�Sz����|�;y�O��s�m�ݰ��2��m\��w/T/|��ʄ2���j�ʜY�[
���*��MUT������"�2�M��.9��FhmC�vׅ�
���ȘU͸��! p�
�(ѻ��	XK&ˊh�����6��^����f�v�dS�.��g*��SCar���x��]��lF�mw�U0��R
����&���f{�y�:m�۷����Z6���z�z���^�0}�)2�������L*�U\7u�������l��y{�K��]��4@s	����\)Coy�!���IF��JSϷZ���Կ�R��(����O�{t�:�����n�yɧp
�
��SxUUTx�:��6�lz��B��'r���=�-�r�����ܚr}�{��>���mIٺdb'���N�_8ʗ��+as���{p><kY�V�D�"��rK�|�bX�JЙ%o�%� �65 1�M+ֺTpk\ܺ%6����U!@�o^i�v{C�;M�&�8JMn׫b�s��X⪐�aU*��=Eݠt�W8���\�c���!uG�T�^`@�ު�`�	zj�;����m�~UUO�UIuে��$1�1�*�eK��/m�~UM����Fct�{�_S��Ckg�]�n�J�����y�p� ���7k
Kc�����
f������p^K:�+���n���n��U�릴�!��E��!�kE:ۭ�u���};�A��D�����[n�m���J���j+�ld��8n���T���UR���Ki�3%�ZZa��``;�!ܼ[��ϣ��fx�#R��;���%밴#��M�_��ѯb��T�UR4�����2��껫Y��/y{���UR��Sbe���ݯ^��uv{B~uu��8s��@UUIQ�v��Eey���a����U �ª����Uڧ����5"�r��x/�.�@�U8@]��@#�L4=�.�L�e�]��n碲�UR�����q�/T/@V�^�D
X3�e���U�*��31�澢�;%j�������y�p���E0�`*�=��s��R�م�L�A�A�.G�kW��Ry*��N�Ǧ�y_{J�Ԟs��!��{	|4���}>��rH,�4L�1t�\i��&�vZ;Ɏ���C�}��j/�}0�f��e%͝����G���6X�.�Ó�cc���~�O��q�|�a>C�w��bКg:u�U�wݑ��>���=�����Pɗ�����ot��d��N�JR3Z�sNi�w%��\7��1[O:�f.�n�^�c��'��>���_x����g��{wB�"������w{��"���~��p������l�}-B*�Q���9��4w�O
�������;��ǹ�y�{�s�J𾝾ѓ��S�����ģ�R���Z��}�F�l(k�i�ޫ\;����x�i/c��pqF�>�j�f�y���3�ʸ���t�];��mW���ۘӚ��|{Ǟ��_=Ë^k��W�9�O5^Os���Xa����N����cw������V�P����o&�.�^�N�z{q�q	��������DΜ��~"�uy��{�`�s��a�r�=<*��\4�:��+��ot��g!o���f�Y`Ǘ�'�r�u[�g��k{|nM��훃u�aܰA4[���L�&�{��]~��tq���ɞ$�N�|�^�,�c��:Oy�훝�\�y!�us����k#׊�����]f^t�SbA��Yw{%	��ǳ��M�b	�?+����/gd���ˮw���X��b��u��f'!�[G��a{.>�c�tQ�iK��?ز�Fn� �z[�_R�D�Uani����
]�)��y7�_ؾ��kҍiֳ�T����E���U�٧��t�.Ş�9���B�4�>O'��t}1xS��ErB�s!��F�^	Y�EghRE�y��c��/}BI?$#��<��+��E�W���(��x����r���Ǉ�ǧ܊/�t}p�+=+�*�TY.��yE�*���u7qF<>>>>y羉E��ZG�yPU���2@�4eDEPyE�5Ԟnb5r�Q ��+���Y|!�7�����UW¹QFF��xS=<��z^<Ő^S"����POOJM�<$����$�{��b{׬�0܈��<^�t���sʼ�OG{J���$���g�z���Ry<r)�2�ّC��(AE�]�.x�+���L"
-��fUE�dP��ڽ $,��FS�H_�z�b[+�����4�1�aЛ��I^�t;n�8�R�{ZJL�h#Q�����[�с2v�6e�%�9�T�j�%���e�(6˫�A�4v�${gJFK��p��͚�8�{5In,Ջ�\�м�\�]��ؼ;;q]�����[���y�1��Y�0��p�9i�s�ٷoN{�cF�3���p���Lf��h��-�l�U۵&I痍���;
��-ȱ&klql��|�S��8���Y��2�9�f�o<��/��,�n�5�=�y����5Y�����W�.�E�{F5�.3�l5u��%���]�[��0j��Y`k7XXK�C]e.I9��W=�aVu��Z��:�Q�ރX*�(-�nƗ3k5�ڹ`���0�H�n��;OK���:�wD�[c\��bh�W0ڍ��e�
�f�x�f��Og����ts6�W���vٗYz�5l��2�R2����0n3I):lMڙ����V/Pҕ-6��;�.��Ǎ��j��@^�ƹ�j�]��H|uzRw-흜�pJ9%=`��GI'U�`B<�!�8�n�(�u�ݍ�[�L�H��U&�-�E���\���@W*��+��;���\�a���<��F��v�a�2�DOhā�v�0�s��E<!��%z7g�4x/h������7(ֳYn��B
�	��[��޲�'2�ۣ�u̕��5>9r�v�ns�b4l��BhY�v�8v�9���/]\�6/;���J��ˋ\u�;�=������Ɇm��rg��p�ݗ��Ėv���c�8�8G�<�a5[�I���&��e9��8���	�66��7n�ׇ�ƵZ�sr1��+�n�����kay�s�����¨�t��^�8vؖ�{	�K(X�n�clV�S�ba�@��؀�x����.�k�56��eQ�G+8躹�8�.��\l�gb���H��j�Iײm�{MիA=��#-�]G	h��;����&�>kn�sڮ�l;���0�ņ��SXk
eE@6��+jB[tE�I�]]<����ez<1p���2�v�h�Z)��# �eo#�m#�ˑ�A��P�ڵ����4��E�-�scĺF�)nX�z�O\�m!gq�z�]������;7gGe�랮.� �nW��Y:�'i6��-��+�u��o\:���)s��{����6�p�����lAum��>�=vNȬ9�+e�w$Y'vwR߂����"*����Ͻ&�^5\]�b���÷��z��]�ܴ���ia�r�������:3��_8ʗ���٤��Yi��ҝ��s0��?�=NU7��z���<O\	}���f���Tk���Ӈ���UU8��S�
�=ˆn4`,�#P�j��2W.~�l�x�qt{�&�5,]`q��!�;��Z@�ު�"�z�!# ̛/�����E�c8�u�z�:�k����
�$Qt=w#�Av��ۋy�uϴ�<�Zf�א=�h�x鳗�F�]�Rp�������=Tû����&�w��-8s��Or��N����a�CE�� �;�������M�"%��ɧ�S7x0�I��1)wT��<<����i�I]qq����dvك鯿~���Z�6qC����^[�˟�u�Uqt{�4��M%9e�7�c�f���&��z�����D78h07�U�8��������STª�w0$vXꮔɢ�$=��n�����g�;�5�Vஐ�@���Q:_��3�UB�
�^��:��p�53q�R��6��ʋ����Ut����ƹڍd&!�F5�qt,[#!�2C̞R�G!����6��x�K���:.���>�֪`*�z�t��k��NK���~=Zd�f�\��Js-9mYo�J���k�����k{��:V�Ҫj�>e�9l�1����[UR�aT�����ƽ��!�Vzj��${p�Y>�OQͼ�\x�үa\#���y�}ٵom��^�4���,��9�s=Ku_����a�j��}ԯ{���?��M6S
�UM^�7]�"�����m0��;Dh��v��Kd�P�#����Ǖ�'�l=�ު�4��UU��s.	�� �/L��!�]o�7���UT�U�_�����J7�״������C"���{';����&�JMu�<�B�n��E��a���/�{���aTl�\��L�2����U޴��xPu����n�@U0�oUUۊ0��7��f�l4W/_Ѹy���Kd�U�S�EO*�-��'�j�`{)�*�������e���L�-��٫w��%u�Z��_y�����U!T�`��l��#��1P6�*���˟���fT\]�U0�'�kz��c��B�%<#a;XY;��c��Wʎ++;F������w翍�eo]i�	�	���ay֧�Ӄ����z�����w��+�b��Sz/�@�ǹW[��K�Y�0��Tު۵���韄��4T�ŋ���X;��_���>8��4��Zى[e.J�k�g�����Ϭ����U6�\^'��-u�Z��S��.�{V�5�"����UX.�z�[uB��H��9��J�o�ƕ�T���
�������*xv=X�֨K�k\��`&�����������Cb�5r����/UgT�<��������:�S��<5U�U7�5���>��n��V�u������E�ϟ[oV��=waxݯUlOl�c�!\H�f�:�c��{�6�G��.וUTz� ���2M�Kp�O'u�i���[�}?xO��N�N
z�g$NU��5�I{��m =�������_{��ozK�<��ܨ �����[,6��������s���&�D�\��t]R��*�X�mq�n�5�ԧ:޷�2��F�Gv�� v����u�y���{�7k���&nqU�3�4�k��糍�H����rǻCin��r������5ȣ�K���[3�?��4���6�<S��l`�����K���\�[\�ж�\��p�3t��k�l�b���=�O���ɴ�be�E31+v��6-"t1½�3e�Y3�,:	/��������m ݥz#4cv���N*z�;�����ɪU����[�ꦪ�T�Z^��w�"l2������q��]���Ն����Tʉ�C�d��ǿ}��Χ-��M���������6*�j��x6��U[��U7�UU@L*��wrbh3����Lso�{�P�`*�z�Fp9�K��r���P�	��z��]sm������l.�u��]L�9��2[��+VC��u�Z��_=�D7����yK�Y���|������/�X?�<7Fk3�AZ7@�+��-odwP�bd�=�m�s�Sv��w_[���SU0�����'���Z���)�Uw�D���֪�*�
�Inӻ;��	�&Sh<���4���/*�(��%S�3�4(�G�IgC9ض��yjj,�z�ӊ��Њ�gm�q+cJZ"�h/c��y���m.���w���P§��?�1q���Ν�?w��<�jՖ���k��h���ͧ�|�x�a�
�ޭ�v�v�����Ⱥ��3�mj�`*������<��*-U�చB�b]r9E�g/�*�U5F�v5%���㐜|OoR뎜�z�z>�aS�U0B�
�~�W�|�>O��a��E̖+dHe��;G������C�۵`�N�wsq$�Kp�3�c��N[W�L7�5��:�j��f[p�ђ\���;u�/:C@�AUU@�j�я^��腘�
��a�6.{��U{Oj��zi��ڪ�i2j�p�L��g?9�2Ӗ���c��3�taj��)#v����ҙ	
�7�L��K�u{D�s徛���I�/i�>�B�f������2v��~��
oM��s�w�8z�u����ݔ/@�op"�U@�o0���;���S.�rv�oOr�Sn�5�n�%�������8�mC_�f6s��+M�a̶�No�p�k���R�:u�^�گW7xM0��UHUC��xȜ�H��K��d�]�^qb��h��1�h �`�#�&��i��ݲ�k����~�>~{������s;��:r]�o��Va9r�CO�y_0�a�����{-�65�����6�vs��xK���ְ_�A��q�.��u��@���g!��H������ULSg;>��e-w���k�M�M�UG�M0MUP�L0�Y�L�,��	�ꪫ���w[�t䧚�;����������ш�n��������Gg|��9,ݹ��{Ɓ��|5�9n{86m�x���p�[�����4l���(R|������UPSz���\ui�<�{�-=W�F�Zڲ�!�C\��YgGFR���h����b��֝��-��30��ǹBV%�1u����fcJ��{L=C퉪��l8�vu��E3;�V������`�������omR�=�狣�<�`�4�]���znj���v���њ#p���{~ɔ�B����/Ul��-O��=�*���UU�����T.��55J٧vX�Er�,:.W����UJ��ƃ��������C1�sӾ�5]e�*��=4��f{b�lv�Y��ʧT��
��'rS�o��X�y�j߲e<н�����۽�� �n�Zɋv�~y*�=cNML��t�7,��-���w�q'�[�$�m���������,��=̞�����v����m���T�))Ȳ��s��)�|�^�&�^2K���J*L�e�k�L�8e��ƞx`٤��(������@	�����,e��R�d�$����uѳ�^��D�]nx&�c���7Z�9jc��u�]Xѹ����ۗ2�j�vG�G������L�o���O>�m�<�Qr����"j���<G�K�;*a�l�{6�+u^���,6.�u���?k�6&��Y��oYw-q���4���m�kk0)�5�i�W����g��~�=U����v���\��������/O[�t������A��E�w�Nf����)�M���d����Mƚ�4{�T�mUW�f�cv��ɲ�� V���v
����w�"GH��V��)����\��Szh�7w>��GV��N`>�����w"vs���\�_Eʩ�Rk��aw��i�ULS
�UUE��@�R�;a�B��d����ƚ�4zat�T�U�����bX+�y�f��2A3�%�F���ch !`,%l,�2L���3u���T���L*�{0E��z}���vptJ�<�#3�9
��o!UN*Mw`.z��hH3�g3;��� ���`�\���L|!��٦2g"����2#T:�S������������U�4;�=�7�qXv���3�i�v�b��v�-u�yh���Tު�Ø�c�X��z���g쵯�?[��?�}��?��~�Mt{���mUJ��Xfai�U�2�/�E�wk�td��;����,��'f���L)�RHwMװo ���`.ڪ�姍�sܵ�hWYx��-�չM�H7�bׄ�
�U�3�������F?���X��%��Ξ�RY!�p��#��)��ꖜ�l1nҙݓ��B�����US��d���tm�i���δ��|n�nq��օS*�5/+䵻��YPs}[�6N�[�VL�������*�;�Y|Z�2�GZ������1�S�Z����2���1%�:=��]0W��=vXj��ȁ x�{o�O<����Rrw����Ǟo���
���2�P�ߖyOR_�پ�{Z�cx�l�o�w��z������~�D��{f{�F�nG��E������ɕ��=�{ݾ�������qq�������7�}���ó��� w�ǛVW�W��Ta�&�,�d)�z���sQq�{�.��y��ɂL�b%���'��<�O���a�;�|�E��Q����dn��|�`�O{E��m��~X�D~ۻ�u^<�+dƼs�_o����a`��o��3�X8>�}�O�vAls���#�g��ۉyǷ6�=g�Ǔ{9�K���}@��dr��9�X�u�����ˀo����>:�$�f�ۙ�`�
��DN�^ �o}�T�!��x���ξc}]�;�ǉp�%��{r��ȧ-����>����x`Y*io�֒Ԃ��A>�bK�ܞ����8��t��̶է��m+}���;���G��߆��؟5��������.D�.�U؅9�u?=9�Z=��s��Ҟ��z�]�y��r�7�O�k@���v���͝�N��p}ø������0���v�0,��{7��ޝ2{_i�ϖ{ڧH-��;�Ó�H��ͣ�O��Y�[�/����q��S�Oj�;%}�u����^�<n�g��e����zy�h�WJ���t�|����xc�R{�x��0A<�i�3
�Z7�^�o����P�D8C��IF9���Rn��Oz����Eqʂ�<�W0������O�8f�G��%x��<���z�O<�\�#��G�i9��"@�xܳ�h��I������³��eRH �fn%ʏ'q�x���6n܎v�센���r���9)Ǉ�ǧ���m�_n��P�ֽ%km�BK �z���Dr7/Ss�]O*�,�S"�c�����>�[�E~M�
�
��\��b	�d�D��N��5� x�gbbh32Z�e��*�(���hQ��"��)�Մű&�Q�ɆFT�%��QD����a&P�ۛYyB�0�rs�ޖ��C�Ij-��Ǯ<��Os��+&�@E;�e�U�n��R�n-� M��Km,D/��@���G[�ؠ�ԪJ@���*��V�n�H9�]o+ނ1�CL�@s`f�����@83)�mx���8:$�ǠC4�(Bmc��y癏�Y�9������N��l���E���z���U4�ˉ{��q����"� �l[�6ŷF��51\�;���t�q�J酋�.��J�1/�4�v��������K>Q�	ۆ^�aT�΂O�^w���wGEu=�8�|q�u��e�S�m�KXj���+�g)8j�W7 |#�⪼*��n欧I���R��}�d�I-�64��UU��f����|ͅ�iD7�m�Y.m�n���jb��z(⪝K���g�0�M��^��
��k����9ي��"hL�]�\Lଊ��p]����8m�v�]��Y
yO7<�*��7sVS��rqs��F,h���^�WCn�t��a���ѧt��l�����m��緻M{�Aɾso2��ѨѷV x���t�Uk�#zXN�k�[2�Od
���U/Uu]�k��ȝ�ace$�d���*+��yo]���xUE���� ���G���Vշt�v��z��i�]!��Rh�
�[�U�����;����YM�UR��7w�"�gEcݭ����OOB�4�P$�C�ն�c]��l��ዱ�;�0���'�wXw&��YP����Ϣ���T�Ub%��>q������{����T�V9���!���Ki��QQ1�~�ǎ�̢���UU#s�3s��}�����j�������{��X�kBv��ڜ�+'�sgW�TxU0�j���b��	�>8�Zf�1T�����h����퀻������}���°���O��i.f�l����6�|��N<��ݾ �)����,o�������'v���ܴ��φ9�y#hI��� ��Ը$�ffe^:N��r�vM�Kq>�*�݋��6�헧x^�a�s�6�tXƱ�����gu��k�U�V��]���Nݞ�����N�\5�ㄳXڄ�:�1�հ�76�!- �&����[˱�̑�;&�2@nbݣ�����[�i�]]��nT���j�|��7w]G��d{u�*�}@;���"N�7f��%���W3����~��[�;@
�O�獣��Wj�fd!|�ҥ����/�}[�����r�*�kC���e�UX��"�Y)��V���m���Y���߲:�����3{^��gD��"8'o�Bj��țc2!�y�
|��*�UT�V�ts�/\�wɧ�e�ј��_z�P��UR�j�j]
'�����v5S])�n�n��(=E�[<v�L�౴��aU!z���j�����0bDn�t3�ow=����{.�ݲ�U0�S�-Y'Du���R"�y�_q�4����Bm�n³]���d@.u���a���K�]&.��?e���T�T�kN���IQͭ��l�����)��y��۾{j̴�qw$���6����bk\Z}�y����t^���r�{�->P�.,>��.w�������A��e���p�b����͠��yLVt3_v�p�{����UXϽϱ�7�tݵ
oUW�=5(=��t�
�v�s:#�o� o��������T�!�EtRh�*�`@����}���:��1�h���u�h��;Uᗩ�R�*����0���[%	����E8z�=�-�V�T�T.dS��7�|nӌ��	|>O�T��� ��.,�jm@�"���.ꍝ��7��ɓ8.��K��>B�eS�����^oV�s�2*��}�,3u�@�R;d]���T���s�<�vx@���^�o���זi�w'>��z�PM�U[�C0Q�:*z�<:��T��ާbϝ�oWϏ�G��������F�&����i�a��0ǋʱ3oe�c:Pj�Vʂ��c[Zյr��%:���0g��X,e��e�����!,��N��(���T�L*���J��!�]�q���MUTf��{�9���dT-N�_T֚gp�-+�W����j̴�Zm�n��ߦ�7ۃ��s湖�vܜ\���xVB�j���R�_�7��$4���A�ٞSM��9��Zɣ/U��c��L�,��r<F\f.���������ϷߴH#�ͫ%bm��{�)ј��VT���{���]?d��%9i�>���.<��đ)ڧ��9�Ú�.xFE4%��]r�We�?5�����(Ms�]���
��O��!wNfGJ%��e;nNs�Y�+)	�
����]��w,>Au�~�aT��[%s�C���tf(���EЃ,�7f���T���&_$��-�=�w���˫�~�o �����q�l1�p�ٌK�y6��m�����j�l�#w�Jq3�yƹu�0����T�T�Mꪆͥ���Nd�^��^�=g{xs[E�Ȧ����UM�5��ݷ��h� ��]���n�����\�J���Wkc�YK��h�����s���z�m������
O*kɾO�y���.ۺ�G�X]�TT��5���Mt��\�|u�W<B���I�=�D0��US�f��mNvLd
�,UG��/
��oUU�n�OA��C�sk��k�����ݽuʩ����Mm�FN��Q�Sb���PͶviRyS^��|�ެ�枊��vZ��
�T��X�v;��.g;�<�`���f�<0����^�9Km󤶅�=Gy��u6�x1�n��><����]r�=� ���E��=�v��@�����,��lT��S<�w�Zxy��H�msl(��!�s4c6uK�O-��8K57��qp�K��ߪ��]�Aޒ�wgev�0��k�R�	���]�!f�7f-�<n�� �r��m�*����Ƴ�٣�\���I	�r�6\p�=�27g���ힼj��ʸ�S���cm���kh��f�Z�zt�nx�2Z�g`n����k�� {�?g���lal��%V���1ڳER;����xx���Γ�j&�~�����ꦪ����3;��73�-���4�[-^�Y�g�n�<���Ç��2����&�w�n��|і{Å�m����B8Z��؈f�4��L*�U7���4t�����z�i��/Sx!�y���U�P�*��R�ޖmjr�6����:ª�qљ��u����@Nް��
�q�ku�ݯU5Sz����4�P�:u����t�Vcu\���Ք�P࿪�ʡ=����=҈�%3X~:���ugr�e�����"��^:˭:y��!�"����|.':ST�����>�d��t^h�{�Mw<�<.[��J���
���*9�9���q/��΍0����o�p��N��fv]>�&����X��-}�J���Y/�C�:x?���jEM͜�qn�e���3;��73�-��;u�U��|���F!��V�����.ک��
��v.CLúZ^'5���ŕr�o�p_
�B��SUS���؋��v!M���%��V�Lٸ�׏=��=��a��}���Ξ�V7�Uy *�U*�����֪�c{��W���Bv]� �-�pӒ����ߚy���-Lk��M]Kj�u7�s�{q�W�͗��ӳ,K��.�ڗh�}UP*��.�&5u\����V���\+��{xy�svXB��l�.�����9�T�y��z�1��!�{����`*�Ũ�{0�����T©�*��F�[��~4`�w�v\Υ�.+UB2���D�W"�6/��8�{�s�gֻ��~�[���E]{웦~��Dw��j�s8"��@�����SU5U �'�ۋ��͵6y
��K�`�S�-;|ӂ�Ք�jX�[��^���UL=Tު�UZ��gA�z�0��<�7_<Ld�t^��{,㋻�y���Ϗ �9�$�Jo��7M���xyC��5�ܔ&:�eS^a�K����Y͡��T�U{�k3�5h��op�vde����zQ{���𪪨���aq�~�܀��T���=pӗ�8/��w-a��l�sWZ��U����mwk�L*�wWt�B	��ôb�����������p����fke����-�n�:��t��j��p�~op�힠��^��		%��>jw��z9�ˈ���0���×���h�Oes{/�[T�޺�R��1�N�g�`gc"F�,�\*���i�ܳ�x�Eݿ���l*���N嶥}�԰�/���r�[�p_xeR��Lު`*��t�iCA��֠�Cgm���c�u=>�Q5��u�6�훩3/��6�cOE�'Zl�|�SM��Z��&��(F.�p�xj��rV5�sW���-`#3�ikި�:���Ϋ�n��p�~o|%���US�k�D����,�.��p�U0T�VB��b6J;��������{���}i�O��i�~��遪�ʊ��B퇪������]�:1t{�������K�bi�U ��.��=�96Ё!��<Mn�/�i�㿷ٟ^=|v��ý������c�>'���~4�J��b+�7�<��tB�o�����O�w�܈qȝ�"A��0���0� �P @@0��@ ���{|\s63���+)Xd��:I]R��+R��+��^:�+3-IYl�+����Vf5�*�cRVl�4�c�U��B�s��c64�e���cEV4�X��Xٌ«2�T��EXd��f3IW]S��2�f�f�
�e��4�a��mR�ٳJV3���ҕ�
���W]���2J�$��:uIXiJ�JV�a�VJ����Vj)0��?�x�,������bPVh�Q�/^�������~w�~�������>?��=�e�����t��=�����������w��~�߿�U)W����������)W����W����/��8�>�y}������?5���JU��W�}�vl�[�F_W��3���������]��ͺ�*��
�إcV�+j�M�V�SX�f��a+Z%lR�iJ�IX�J��VV��-IZZ��1J��VF��J�d��RV��:�]U�VZ��h��)Z�+VT�Z���V5%fT�Ԓ����+7G������!R�
l������~��ݵ��?5��s�����_���R��~ޯ�_���:w�\����_���Gu�iR���+�����9U)W�*R���W�c�K�x}:*��￡z;��*�Yu~�u�'��gW��m���8�����Ú��./��J���g��g�~��o��R�*����^?W����>�����������/��꿝��)W��~O)Wk�W+�c���߂��M��_���������x�JU�~���f�_���]�������������T�_���:�����JU�������_��]/����e5�[D�T\� ?�s2}p!���                                     0�� )@�$@�*�JT��*�T( � �P *@�PIU@�B�Q@��
UH/>��J
����E )R)Q
(��P*����U(�*)U@(�
U�)%�@H$��J�� (�����R
 �hk�L%��ꏫ�w� �� �EE\ݎ%���zw��{ :��B�� g�=)C��׊�E���  �=�����|���oЧ�  @oMA@
<�h.� i�aР�!�g�)\C�� ��� �9��B�P(IA� } |(�"%AB�(

 � [���z(�"����t��u���
����=�A��N�)EX Z�B�4���Z�TR@T��   `=��(}4w��n J�kz ���]� ��� ��� ��G�;�נ�X�;���(AU
���  �ĩBURUP��E*$G � ��:u��o{�������� {����w`�A�@�� $R��/�  �>@ ���
� �: w` � �����(��-��2@݀�]��AR �  ���T�����	*� m�@.� �:;���Xlt��:�� n�+�r ���

$>�  ���o����9 {y�d S��ռ�	\��z @g�{� '@(���� �)C�$��T�H��)I(��=�� ��-^�T� ���[�<��{��;�z�� =;�JX >� ����A@"P|  G�`�ݟK�{�Up ���zw��<��  =�E��� ��C� 	���� jzh4RU	� ��E?RUC� h'�J���@  M�����  ��IUM��   �Q)��T��(<S����������P�FHc���n�&����7ti1>��BI�����	 ���!$$?�$O�	 ���� �$�BHHs��U��ԣ�ƿ����Z�����:9��^ܐzt�l�%�[�5b�"�y�M��z
�
��x��6��\��8�mYhꝙӱ��j���:w,���B��2%�81���m.,ߴ�����ӁƱ�$�f2�w�*'�������o[ҕ^�Z ��%3xww9���ӧ8���˕3�v-6�A��`K/l7�b;;5��MZ�k�i��!�ԣ{:�N�7g:�Ś��3���g��Y��@��f7���@7����%]���T�X���v��mv��o6��x�p9ӡ]�q���V0��Ń��!��v�
Ր����[-0b�fvU1�ލߖ�w��h�<rrL{���R�Q�S�ӲT�$9זu�(7�,�ou�{p�U���^�*���z䰽�׶[�U�z񫆮κ9�@�Xs�gNE�`Z�0r�B4���v��ɼ�v��o�^K��sXd"'���x�em��Z1�BG*�ƁY��7����[WL���fo}�xgM]�XgA]�Cs�t�m�������ۮN�+��xM�N0(n�Xc��n�<5l��9Q����C);�X]���v�qyNNF�<u*+i漹����d�ߌe>�D�U�uWnn��l`Tq.�+��OA<��`��z�,��+�X}ȘO6���pv�໴���>��`f��wt��/L�&��G>�x1�Z;�ܮ:��v��A�1�wU��@��f��~�7ol!�,�ӹ�$�چ��b;ȹ��'oA]�.����(�1R��غ�D��ɲ�����f�q]$T9��{v��ǌ�5v^s�&�Ƈ��Ҏ�5&&�.C�[���6n��V���bxPz7�K���Z��k���c@��a��3�s���^6�?w�d�� �;�*5-A�{sL��y%�e���vW1#�E�yзг�T���h�v�����ܚ\b�Y�!# �+y�.{t�A~�'�r�pb�7-=��3�=�77��c-q;�([Ǚ����ٳ�B��N��vUWE������`;���r�P�Tz��0'ٷ�rِ��4����*�#邙�l������j*\ܳ�j姧�u���;'{w�	�7����Kv�r�����A��J堜��L�= ����g���im9��&Au����J��_<1p{G%�M9w8y��F�2H7nY�9׸���E޼xC�ĵ�i=8��X�����cl��nv=�K�;c�'oL��z�������;�ua����z,�#�jw�n,7���р���^m�2i/�<{�Lic�f� ww:%/�[m=6������B2��%3>4[V����'W�G�e��4�ݥ�3��*�*�4΋��Q3����R)�N���L�Q�8��j#�:JGd�9@΅�G��7Y1@GWe��1��[�:������͌!5$L<\{;yT8���e�7�̈́p��i��~�Q�od!\z:�X�ޤ�7�e�K�a�FMYFC!;0�a6p���-7w�T��XKmew�+I�YgL�����ɻ�;�����x�	m��߻8a��^����:�M=���gۚ�8�
���PC��8tsH��JV�|�r�O��W�r]w�ň\Ol��Z+H��E��&�!rP9���ٸ�@�`/8L��X���뫴��VS���8mV#zF�A����3��d-~}��0sG�����+�]�D�e�Z���'l�3K��H	�.SJ8
皻%��vԃ��}��S;&nw<ٌ☺$�k�ӱkx]|om�a��k;$S������K���;��C��QF���9��Žޑ��C�)�j\�C2PDx��_=�h�ۜ����3[��l&� �{����&w��Q`�n�R\����W4oH����u��>�p`-lLuo�1lW�wDnZwy|NQj��f���ˋru��z���s�.�XHmjH��t����:T�Wܗt4u�W�J8\q�Z"��cϽ�X�i�f��L�Hp�$�2�̔Yf����̌B���N
Q�$VZ�SY�X�֯W�N�:����<��K�쑼�0lj��7�f�n�X۫J��ΊĞ!rHz�c*��InZ�uV��Q�z�D��dĞ�58s�h��w��F�G ��}�*;�t��v�D6��q:s��2��q)�l�(г�вP�����ɋ.��)�}r@
ִ�zh��s�.
��vq�w��v,��A�%��/$~`�I�;����. �	��S�t�Oj�[�od|��Jq]�${(x���9RU#�GB�A�.����&b��IԏQ�逎���Q�f������l�n�KC���&�Y�k�(���KUl��wLo+;Fbʢ �e�L��9L��N��ӛ9	�Qb��[ܻ��-����^��ar����ݜ��'y��_�#��Z9��/jo��v��r�7-��q�׋B��u|B��@���wD�n�����=N�t�׷�[��t1��b���jٛ��[2�4C�N�p&>�@�!��w��R����U��v�n�V�����"8��N�;ܧ�0ͬ�øV���k��O�Βû��T��{.4��;�\ٚ��{�j�⊁87�x�o4���&U�h���2pAEӰ�Ά���;x.{�e�Kc��3��0��q��)�7H����/�&O��x؛C{o<��f��qD��%\Ӿ�W+�.=�%;p N�{tu��"r�� �^(��	
LXFDԳ���'Y�^򸃄a��gn�p�v���rp*�BqO��B	 x�!�he\P��mI�7;�\�#�s[�'�Ԑ�Zn�2J7Frѱ�4��z�o��'��^,J�%_ P��fo,��=r=36�yejoF���@Z3]�D�r�<-F�l�K�ǖ�gd���j��ӥ���-]Qg^��7�.��^iس��<��i�i���N �-�vqgd�㱥�dv�9�H�5�����B�gj�z3�p��sJT�i��쳷[�'s�'�S�nȜ�w���!W�o)3bɣuȘ���n)a�6�������}9�_q8�ѳ�E^Q6�w
��8���2> ̓��E�i���yv�å|[�Ū@���Pd�짫�/4w��F��1X��wt]�D��I�f��TV	�O��]�ΌZXl��[����ƛ��μ�r��:N�rf��χC�)�3fY�x�|o�%�a�c�5n�J����g��]���Ѵ��Qr�!�Ɔ��oL��gzp�{F�؎�\n�֩vt�����>Q'YͲ���*o,�u�ae�}��'��gXTA��ww���k���WG,�5R<�/��s��s5(��v-�4ͳs�qW�����:�mkK�Ð�z���	���,�Ê��9�|�Ԓ�Z���c�C����-ÜuA�e�|EMܔ�g\�n8v�C�� ��{��.���fU�J.aѓ�q�i�xvU��ѕ �[н;2������=�E����[�v���z�	Nu���D:�+ �x齊���W%X�IyRr��a)���8�����T�ı�d�$���:��)J���{AS�K��0�pќMX��tZ@kWvjÜ��%����Oc��ڛۼĞۜO]9�$���*[��ե�E��u!QVi:��A��g5>z�Ut�)Wj��Y%A����J��싐Y�7O^�p�<+�˵���4�[��g^�E:z��ɛ�c����3_p�t��^h��UR��e�������^�۲�()�z{9���-��f���ם�/N�>!�m��8[�6W������<�F��T[��
8 ��"Y����o\��a=� 6�wQɥ���{{�X���^#.��f�ۋ;���}˓₤qXg-�32nG"�s��Ӛh����=}�t�'�-\!��3�ל��[��坽JS����M]�/����%5b�$���������7X�n3իuJ9e��M�ռ��7�����]�[M���Fv��3��x���և�B#8C"�]Mz�k�h���^�_p��%� ;6s�)��3��oq��<4��	�.�N<�3�s�4-.�N�i-��2��۸1�U�(�<�U���8w6��Rq�ř�p���;C��>��N{u��T3{	;��8��@��c�=��7pE6�l��dȴ̀�ܩ:�"wM3�fv����i�{���%<}�&=���〳���{�����#��(A��wqT�\$nR�rG���`ۏ��]ٛ�h�͜�@.����,�t�Ҙ�:�r�"m�5�t,7�ܚ�h˩�ۂq+�I�i��{D��(K9�d�{v�a�3In���{D�o֞܎�u��`�Ջ��'�����:oQ]���s*��@�!�\��oQ����"��11ݠ�#�e0���y���x�ִ�7`U�AdOp�A�$Fh�hF,\:Y8!m����{zK�T�֞:
y�퉥��7@�k����F��O$��s�9����\�ed�������'�Y����u���띚4@��vh��� �[�1���4;�ڗ7�:�ys[�{ ��2l��YwZ�˗��<e��f���v�G��������t��U�B�#�gN���� �#��{�&�-���v��ow|r5ZD��DѵAr��ײw�v�{:/e�˙sn���n�,��c��߫��	�2���
JX5��A�����,�P�ݗ��9�R�5Q�����
��x�yd��2k��C�Y���- %�qΔJ�g�뀊���|;x�H�_��نpE �f�)ܝ[��to5�w���8�o��#���qmˋ{�ד��3J�r�#�����v�aW���kŃ�]��k�V��L��Gv]�JJղ\3� ���
s�R��NNC]D��\�F���y擡�Ö�fS�<	�[b�8a,Ƕ u��hƯ	U�n�xꩥG9W��v�II��*��c��%���2��:�v���A�m��`�����n������y�wg)��j�懃�)i��˷&��5���a��tb�Æn���!�y�ӝ��w|���X��ݚ�Gn _��^XZZn���i6k۽&ZN�%�i���|��y���!
rXJ��oC�z>2iPj?u�ɕ��c�Ԍ�C����q��L��~�]\Y�fNCwgY�S��e���>��C�i����#���xvܸ�L8t�G=���W)x��Aɝ-�ɛ�=`S���	3� ���z��TNp
�ws���%�����tDrN������bԀ�1q*־U����|�e�r��`ѡ�P��s�N]���ZsN�0f�Q{F���ho }ֱZ'gqd��G�W7(�z'���}�.����ϡ+�'ΐ+۩�{t��[�u�/+=�-O~���LW^��sYW��t��T8�YC9��}�'�ɯ�����бİ��V�@�>�ຩ�ڮ��0Њ���員���0��;�:�Տ����B��j��ېRV���ölt^cg]��eZ+��#n������Þ!_-��B%�4'�˰n����u2�k4�:���9��z��k,w@�PD�4��6u}�0[�v[��K�7����Z����{E����Ο,x@��2x�9���C����W�$�c�	�$�W�����/b9�C��ת�����4�c�_Mݕt�F8��Z��v7��-|���)�GbWWt`wo3��wg;�glW��z�L��Z�zøM[ۧ��n�yi���S��y��u�m��9�ga7���(L�Q�ǲ�U.8��AlD.�EC.���pB�S��5�8�|^��+L�h�K:��NDD�~����pa/^�9,R��][��܅m��*����V��w��4�T�a����~3v�_u2�F�8�6�5�P
��.����W,*I�.���F��}��j�n6�׋�ud<C�x����ڕ���:�t8]����w.�2�h�2M���.��c��nGkszj��M��c�:�}���Y�;�9�y�b<[�:Ր\^Ÿ�Agm�t�ى�^�[�&\`,C�3�HoE+y(�:`�:`r�`ゃ٤p9���2��R��@nk��qi%٥Mǀ��\-�Z��+/=��!莵�`Ν�4��nE�T�6��-א�1;�F�CS����_��d��.طIO���St+Q+����f!7M��N��9�d�*���l�җ����{#]fDP���!�a�c�|i;�R����Pd�qvi�0+��zv��Y(����'��I���L���B�Xi	�����@��ܣ�n�T������YƋ��f�(eb7zn^]�C�Z �Г,�2]t�{h<���B�=��W��7��ϱ�QikUwE�d�p:��+��u�<�o12�E/^Z�]�t�T��(݆��ŝ�;4���7Xn7��m�s����lkz�[�6��\ϲ9jjԨ(�,i�`�+X��j+7+
@m�L-;w�r�O5�&��e��W��D7ׁ��� ɶ��}2fD�W�׍���u!Y "�$"�B,�	BU�	�$X� )	I	@RYI R��X((�I$�P�a)E ,�"�EE�"�I�,��P	�"�	@���`AI,$�:��*�껊���*�H@�� 
@�P��!$�E��
(�Y a ) ,�HH�a$RI�H
I$Y!�d$Qd��B,�d�RE�� I@aI$X@�,�� � XI$�"� 	BH� P (HA`Ad A`@���)� �@PaE���@�HC�$�BH=��������Ị!�¿NX�d��D��%@�Gs���<�tMmN�&���o��G��z	w���z�wF{�4s��2o?#�����#s�ٴ��&�ԽO��]��"�~��\�.��[f��nq��k<�yo��'�^1�Ⱦx{�O^�vΦ��+���v?{�t`���95��������{�Ó�({r�J���=}�eЇ�1�����w��N��ݞ��|9�3ǃ����{��gOG;
W<�[���LA����Eչ�w'}���n5���~��D~��0o���v/y|w�Q寧����i��摇ؐ�Wu�O =���W�ZFt�iRN,^l��rPs��;��ǽ�����{�N����圷#��$޵nžy}�q��O�E�VR�89�ufXGѬ8��f��M�h�흞�]עbu-{��K���z�A��3��S�o�Y#�:\\P[	���Rn]������c���uoMd����ˉ�_�#��}�!Ӭ�M�
�ns�����ټ�޾Cm,mx���3�,��OBI^U��9�̏H5/9�ڪs�<�xv����&�#�mw��<�Ʒ�g�w�~Nź��N���b\�K�	���3ǧ�ko���4��T�̊�ͽ�^�0q}ws٤o�1�ٮTO��H�w��;q4�A���4��UlXZm��m�ڶ2�N
Ӻ.2�V��aΘ����b�&�H���Ч�uw�(�_\��O�YVi�kM�R�Nm܉�iȋ!b;2ߴ���z���7���ֆ4���0&6�ȸ�^^��aEʬr��h�?`����l����ϳίL��f+�d�Z������	�mj<�ׅ�q͙�xK��o������K���A8q� �Q�0Y�S�v�)�	;�(�ay�2��^��֤c�N`�:}٤x�c�����{���%�`�Kw0�xj��y��a���Gg}��@	��H�g���ٻ�g\�nj��M;;^������#��ń�^��:%�m����OO��:���֯�օ�7���u}���)�i�!��s���1{׷�3ξ�w�v���Z�{�w̧���B0�22�Y�"�kf�L�6��4$E:���F�n��6r�!�[�K�T�\�N�L��r��/2;�E�{�;��s^3�Đs���I���ǌ��Bu�}���Wf�
�>;�F�~�M����Rڷ�I��y/���'��=���p<�4A�Yr3��m�z3j�.�s����=�6gh|N�ͬ4Vc[ɔј�d�Qw�bL���s�E�Elo�NB�,����U�,���!�.E+�=��d����fm�i�}�u�|��T�"̩����8��I�A���#������OW���`������/Ocy��3���jI�3ڧo���9�
�W��P�C�2\l�w-7kUŨ�B(3����횀<]Ɂ��}b2BRQ����nrq�P�v$�{�؋�"u����~6�l��ohn=��P��7=j����2�\��m�v���7ȩ��p��sQ�^�F���+��;�{�w>M���_�%����w�j�9���o;L?s\�} g�<Jn�m�<�U��U֓�O�٧F�l�Y��\�ܹ�F�N���{"^����{�D��G雵�3ʰ�j fomgnRN��?G:/D�/y�ċA	ܻ"�f�e[dj݁*���ma,���{�����ܧ��O��6x��)ͪz��{â����F_)�z4�:�egp��=�gO9�A�����傑t�{���	/����������-i�N{O��̍_`Y�=��v�:_3��8��_X}�����8A����ٽ��]��	iY�`\�n!Ӟ�wy��9��3� ��#r&Z׊�m��yF-ŷx"_A����<��Oyn�:z��c>�Z�X�+ե��ڒ	�5-�]V���a	9W�#�l
*/
�Mf/o�K{{F�m���}����Z�5[�a��ᓢ���`̆iz-���f�v��Tw�wp5��0y���J��-�˝������y;ݯ�m�u�������ޛ�F�]o���͹s���Aʍ�R����P&2#��O/Qܻ0�ْ�{�s�- ;�{�����UV������r�ҋ(UF�y�D~�g�t�v���-�&�;��n��ρ��1�K<����v�a5ư�>�/R/Q��˷��]�R㫛N�3�"���}�����c�ˇV�Ww��xû̈́��==�f��w9N�ϧa=�է&�m�D�n��G;�r�Vi!��d�S�⁐<�M�9�5{���~ӛE[��i�9e���7,9Z�Ws�{:ov�z�w�����2GH)q�{�{x�Q<�a��<�_x��>1�Sck�z��p�ۇGU�ɻ��xbx��M7���aW�g���a[ؽ�'،��U���A���!�^Rtጾ���.�f�ko3Ӏ�y�M<^���d���;�}�ۄ�W�����0��i�Vk]�M1���d�o�>��zp��v��W�ؼ�q�t�X���ު�F���r�y��4G�3��O{ޒ�}�,k��='�d�d����kc�g���LY��|Q�n]=���o{��=Ք�s�}�1��:�<0i��"���0�ٛI�׶����u%���Wx��=5c���vM�Z�kե0䰤��,�4n�إ-l^1Nh2���Ð[�����n��Ӹ�{�wۊoH�1���J�=�|Wi�yPƌ�eń��4�#�)�\v�z:��e���}�56zp�>�\w��x#f�l=�Ose*;e4r�QM��0F�w�����x�����N�7�9��m�<C��z{�xc��,�3M{��<w���=WT��ƽ�'}u�4�p03Ɲ��4S�sЬ}e�4{o�A/����͘.��mwi�������Y\{���<Ը��u|��?�����[�����{����fА��o��B�=6�:=�����mՓG�u��]��_m��{�����11�{��kP�٪)�>�{΂�+�%S�v
���Ȟ�Bt*m�7�_t�"���/B1�b�P��f��j�
�yG��>�u�b]��nn	�{�-��q���_{��V�����Ŏ�|�U��{�&�e
]}�}�0��HAe����>ʽ���7����=�N=X5���*e�]*.:��U�@�͝0�DHB� �L���u���x��9�˹-�,'�ʣek�5r�hJ.�������v�vN��`�f:��KX� Nl\�-2��"G������h�ɮ�>>��l�l��s�SQ�YT�����{3�2�l� t`<���uw�>|��^M��/y ��{�<��iL�˄yi�P=���{�{Ďޢ������ݞMj�[1?�oN���=k�z�2Bv�O��ݸ�]rp�{��&Θ\��-�i��3��fu���U�.�=�~b���[���Č}�3��j?#�)�2��=��U���a����{[�eDY�_f�ς��1T�����'j�Ք��e�nxK������������X��G:%���&E�,)�3��C���|�V��c'��/i�~[��Ԭ��U}���Ar��N���&�ݶ>��"h]����8ޢ���p���T�bb�C`^m�żv'P��0��S��+�HگM�I^�|����a�$��Ŵ���?�G������osQ�{�+<�h=����Wmg�r�<�&�|f�f�,7�}/=��X�2�,�����������/Xy6�h��S�h��S�ډ�J�g^�"b�#A�{*S]�坪�z��ox���
O%�{�_a�敾��8�y�%�����kW�=o_u���lx����'�}u�w��������݂$�m�+9M��y�!�� �=9����fd�ޫ�|��mK��{���B�4��s�[1F��7�:��=�BV�|W��&C�SznzJ:S�ׇ���w��5��NiьM^)$�z{�>���\'�F�ůh2���}���q����{�Ǟ��n�m�o��
FS��ǝ ,��\�����sa����(�ּ{w9�fw�XS�/�Mo}�z=$v/kL�s�qKraf"�1�U��J��S3zЙx��k{�i�����E{K^��}s���uh�v�b"�ɨ��B:�k(F��B��ځ/7&`�j�2s4C���Ɵ�x�b���oS�sT���ݕA��{��_I�%�E�5.ҠL�jސ�pn?c��܋/]��9<�0=��ݸ��w�w���\^Q�YL�u,?G�r���#���6k�6����vv&�r�.�7�}A�蟻��<G���Ӯ�V�6d+-�t����kq�Gm��;�ޚG��P��M]9Y��Zq���ҵW�}rǹ�S��2����MsX�x/oih�p$x3��UЭ��f�L�}�&�\/:���/z{/�m[�(�7�L5!m�$�v���ݥ��g #�ɶ=����%���[5#��;�x;ӽ`��V�橂����<�����'e�IJ��m�v64CFAsm�/jk�4�g^��WV#`�_o'���tf�d�H��{�Ĳw�2m��쒍�/A����sA��Q����U�wVC��.2��!�[�0un��ǹ�v��Z�=�ʱ��IV��jN�9�_0�|w�c^��,�E֘�Pk�D(��ݞ�&�-w���$����kt�f�ߓǂy�8:����gDA�a���vћ��變�7;Y�md�����F����e6��[SbN�]�e�1��ڤ��n�m��i4B��1kힶSOXa�7���oQ���n��{M�U��ʇ)�ê�g�t�0ԋ��C6��ۣJ�YGyr�x@��wȍ�A'��`q���	s�h-�(�k_�e�E(��Gt��E]G�n��l}n�j���j{�Ӳ�&N��廉D8H���!�S���R�/ӷӰ�'7��m.`����~�Y��aU)ax�g����i���xA"�wF�k(�[�x{t	���I����f[�Y�m��̙��:{;�5ggz4|`�Ǟ߅��OC����̽x�J�L]���7�R>^��
�=
}����-��L8R�?�_GC��#������gg��n�`^{�ᾙއ��� �'�4}��O.�;�mn�1zW�{��*� 2q��]�Dc�r����:�I�9AQt��#v�C�b�dۖ��4@���m��0Y�}�A~~ˁ���^��G`�:�F��A�7�'�r�+�peo5O?,�w���V�f6�Q�;�Z
r���[V��y@�n�Mh\���{��7���� �w�:�{�v����9�������^�l홦To��7T"����{��A�����ܤ�goJ�UN;�x�T	�^ؘ�Y�2��kL� ۱>É���zn2�� ]��)��s*D���W*��6w\��P�O˧�&�W��،�9f�Yw�e٤	����{�T(r�Z�ͻn����.W��T���&R�ڧ>Y�-o�����o{����e�L��w}o���v�2��՚HB�H�Yqr��(�vÝ�a�;4l������(�8�)�}�o�!�{g�����~��t����e�JZ�D�Pf�	�S�H��<+�K�:��g��=|���[��p� A=ڻӚ�Vdڠ��Qs��OE;Î�,\�gB�����ѐE ��j��u	�kF����d?`�!���m=Љ;3.�������;��PC�39�A��<�p�w}c��h5�Iܹ�e�<�t?Y�n�toՙ���� ����i��v��|$��׼�I��{e��bw4��j��s$cs�Y����&iЄ[�m^�����@rK������I.�D�g�e5��u��ջ�1����n�C�+u.���CǓ���Eޯkփ�;���r䃰U�<F{2�J��{�K��RU�s�ba�b��Qq���K��H��z���'��{�����K���cǅ`�Ro��^1�K�E�'�C8I�U����/I�.��6f׳�wOS��G��WU��J��
�l�xk���f8�d���Y~���Zw������X��W�#�z5����Oo>�����#�⯭kC2��ۀ�LN@�[��,ȧQ9��x>�G�G~�9u�|쀉}�~Z��ܽ���뀮L]���X����NoT@�;;XwWi�_a�������9B\�D�z0nf��اZ,Nn�d��F�<*n31��[(A@JC�6�V60�M�b[�������kL�׽����q];��xX��#r����d6��}��ί\p+�W�C��X��gVl�Tѫ�q���֭^�bkfd���0@&�{K�4�wz�O�3>�s��-\��û�.����;�z�4�"o�{�ݜ1e׈]���j�w��2���c��*ͪ� �j�������WF��=�`!�|��<�_tw_�K�	�rw��x�
�v��SI�9��]K�vO���{�P��Y��gS�S��W�#S�]/��g��Q�]�`A�_f�aׂ~�����wg�G<F�����}��}�G]J�F��z{�Y����/%��5D�꯵v*��i���{s����
�ީ���T�5.fgYqq6&2�����#jN�m�9��NB���XFw�y8H��g=�D<��nmn�zh�4�o/�*ܛG����0�D�`�*$�vH�wh�pjK�u�6p����8V@�'O�'�u�����g�s]�{X�;���3b��/[�&��0�:��!?,�3�٥��u�Sr�݄Ɲ�������[���J�ͳV�޼ϯ����&���מ�n�o���͞�,�OAle^��8Of�q��~��^�����| ��M�2fK�;�,;��M&�����PY�p�"��m��E։��ܦ��+� =����  ���ݨ5bn5yβ�j�R���ѷO]W'm�4��.c,f�`.�SiG�&&�S5�kW �`���κ,vuq�'Y�4`e6�� ��'�w+D�<�\��4��6����+e�:�oZ˭��*�=����DK�f�kf.*ZKh$`�Mͫ]��n�V|ۭ]	v`��j͸����cf-WU��M�@����u�\h���[�LF�ģL��;P��atq���dmfF��� 듺z뱣�������s��ڮBqu����gi�,c$mE���8�fnq��:g>��Mn�0r�c�5������b^���{�<q�1��/B\s���՛�w`�gu�Y��d�͞3ǵx�'�7����4��ke�Xe)�/��6��*��V�S��ێb)^�M�m�z��=Q�aۨmQ��s&���DB��n*0��Rv�ݚ`�+0L�6b+��`�E����7���:y�a%�M�ݮ9���b�7A.��G�#aDi��R`.w����Q�<W��5M�yy'��7���ֹg��Nɮ��.�(������	9�K�b��Y�jF�gƺp�����M�<�$[mXgb���hGL�
v$��ފ{m�9�t�k��[֙�c]&���Y`8�ty3m�h�9�Aȼ�,���-�%i�v ���q�>P$ӹ*�A��[��pwE�X�Y�21�=�^�/A�-���t_w��Bw!�G7:n��Aֶ0���#�[ǂ���@�w��5mv��e���4J�.-���s�#H��jιc�c=�Q�msN���".C]��Ѷ�sn8I)��x-�.����FM=:�e�z���Ԯ�ʜ�ٴ��5��+�݆���3�k��Vݹ�H��M�I���a�s�Grp+b�A(�����I]5��D,���TN�uQ���'#��E�	�1-��v�)w �ZB���r���(��C:��'���8���Շ���N�]l��\;l..ghV���g)Y�-=�-+p�\J�4�t��$g� ��q�#�\����r�nۋ5��8��`z�d[����)]�Sfdq�S��I�iM3s��F��%љ��3u�u�&���<j}��\��h��m��Lv�Q ������%��n�`άc�	���V�X�\�j-I�fմp�$��!n��M����䭴Ω%9�{�0���8�t˸V�=��ֽf{A[b��K]��XFw8��������ۋgg�0�y;��MGY��&��e�88Ƌ�<v��-�vwk73�ۍX֐w@�����O�}|���x���l"���'1۱TpE�ձ��}Ԃm1�n�GgS�:K��!�v8�469����^͆������RD6��MI�e�N�	�&-6e��ѹ)��m��8v8�h:�#]؆�����>�s\��_iurv��9�'��Dv��A�� ��"�q��}����6�	Su�m֦i�K`0C�ûZW�P����a�k���.��5��4��]���r%	S��Σ`��.L����yl�K�'�"[Q`ձ���b[��tl���M�[6���G
LK�X����t5޺cl�ƳEn�
�)�c�d�gm�e�Xz4n:�\v��X�1۷:��@+ό��6�23W�6�e.��C�m��c��k�����		5�N:T�wUz���l���cD}�ױ�˘��5��eID���������f�a����vzt.-n��,�Jqm,�sAFr�4j�N���1�oWc[ҁr�6�v��sڒ^v��֫�+%㍰�!'m�+��W,�8�P�m�v��2�S2��(89���v����g����=&�Ӻ��ח�'���$(r��uh��n��\����JA�[�`N�m]��m�\8��f;l��Ԥ��1ۆ�z(��76�N�mڇgv�uj��ۜ������㮶�S�{P��Y��(��
h���2��Mk4�,�;:a�Ź�fn���Mt�����l��T2䫢�.h�[��vu������@9�Iƍ2���v�q�G�<�v�y��`l[���V�v���x��xy��Wh�8���Nv�Qڦ�k���|�:-�l������&���u�'e���h�'jO]���we�)]�n����V�x;h��P�x���F{b�jY�#h0V[,�ӈ.����BӃ6�L�F�=R,�d�v�K�
YZ�g�Y�ɖ�i:�C�^v�8R`�z��u��ʄ^��MDv�K�u�L:
$l���b�Rj�*u��XK��b��l6��g�ɻ4�*���]Sn(�����>9u}�]g����L6�x���:��Ld7 �C<�v�nk�M�ɴh0Sv�^-�v���^���>����dl>Q݊��n�N]ZS��S@�j�������.N:)�!�N��v�N닛�99��F����c�lmz�+���q��1�v���i�K%`i�λFFZ�wg-�m�pAo�mX+�D@in�w��κ���@������Q&��:1�q��q�q&n��dwg�v����&������ǭ�{�M���H�b����CKn���u�۵��нvN���@V�6�	���۬�6�f�B9���l6�/]MFZi���a�����-fL=�݌��x�U����oT�!�d�:;��
G���W4e�0Q��<�Sۺ���#Vݷ`�p�	V�-� nm4,eT��Q�Wn4v���|��}��/�W���:�8�lc%Ŗ�p��Mu1�C�a�Qƺqv0M�\��f�k�.��t���]h����+z��[vV�p�j�����u�v����7.N�p����<�܄^ڸ۔ݻByU���'۾>��n��,�f��S@�ƥ!,.��XLmQI�)��۠�\���b�S�~>��OAϫC]It��n3^���@��K�ruĻq��s�Ht�v���[��@�XQ�XmH�	�tml+�m��1�!.MH�J�DLFX$�)4(Lm([+Y��(ka�B����rP��JWmv}��"�u��v-J���Y�5�AΊ��L���h���J�5�^�D�B�c���n�^���e�n��>�RUڲDY�gg�d��A�sĠ�bY�ms�����7Z;�5ä����kEד�l=�v�ycsM:�%i�Y�1����4DM�R̯Z�B��$^���l�V��d���C���&�5
c��t�w2�X�C���{x���k�0�p�4bZ�5#^Rl4��5�A���k7P3���%��v(�4!-��t�,����|t��-�V=����Zn�v���А�t5,Ѭ��:��uH&�v�+�0fj�[�nJR1���-meԑ��vV܅e�;�sZ�������m�ְ�9�c��s�FIK��Mˬk��@��t��"�W�2}�n>�7���I\�9���j��h춹�ϛǢ�$�K�,�� ˮ��r7Cp�ɥ0�%׌,nU6�b#E�[l�`��:FG����x�)ܛY�@p���NA��I��8:�u���wT�)���tl�8�iz�x�\<�7l۳I��8�X��8K�[dya��g�{tlp��K�1KFK5�3f��p�dӣG[X�:��t`�r�N���0�p��X�8��Iܛk�W9��c�1�r�+׮�v���D1=�LP4^�.e��k+�aKC��vc�n� =�ශ���s���@��tB��Дi%���6RŶ5�9��;z�F����#���e�F4ҕ�����qae+rY����:���]ەؔph���`��r7m[�=[�خے��zq� ���l�*����MK����n�lƄj49e�P��:�+�/T^���l�ݎ�&a.1�v���T�.
��w�);+�]� �lzn�@�m�fM��fM7][m�#`9��6�u��ۍG�F\kD��=v���OJnzƨ�7u0m�bv�M����Җs�c�sٱ�_o��ۻOTa�7j�n��1٫D��͸ĵU�����������.��h�ֽ8�wn��W��9@��yQ�f�:���31��K+���\!-�Y�q�2���lp������>��R&���Ar���c��:lE�S��A׌k+yi���N����p��pқ8+�Ԝ�ޮ�ͷe��{O`�Q�&�A�7}s՟�ms.&`eB�Lڒ&�M�O��M���z܏3V%����x�t
r��֍I�4\Y���* ̷ ݸ��m�C�')yz�pV{�G�+my�M
r�J]��;d�����>�gU�vخR�x�ݵI����ǔ�	�ѳ�k�MvՁFj�Z�3]�����1/g=3�M�3O6�.������zf�����|Qʺ�a�(���.9��h�.��-Ӝ��������]ȂӸ7�ݦ��i�$�ٰ���.㭷8h0z�¼ݺ����/:��#{-��d���k�4�$��0����[��'��}w?m��d6�F�Z$<�y�nW ���z�L3�Kt7o^Dܞ�i��8�kn��	Z��cz�]z�`0%��֭��^���u��-�����&,l�Zv�7t2t�4-f��CZm�-��砗[��̧9w�;�	�3������������4��@�����U	\J�+7@xjM�js�[,In�[Ħ)i�[f#
)�vW������q�S��@�)�!y���VX6%vz��<�E�p�k�u��������2�Ǧ�t�ւ�+��pi�Q��]�L" ]nN�<�vk�q�i��XlEpV�"�n`��3�p���&���'Y��иpUCYB��)�$9톚��ΗKW��&#14�B{o3�&��N@/3�Vl�e��æ���T���x37#���T��vN�n�٢˙����H�ƺ\Wh�M����!4[-�Ka�έ��JlU����[e��J��~e�4������Ή{M���z�i��[VD\[h��ud{�f�gggi�du�Eg�������鱺-�w[n�0��!�{=Z\�M��k[#�ѷ�x3m��%���w����h�gf�b�v���ͭ��d��bvT�:͖ܲ6i-��M���	���m�4-�vK.l�޷�	*� ��oR��mmv�i����ݶg��!$ll�T�RC�l�G����	�5�a�3���޷��;3&n�f�:8���絗��[bNY�8���B���K6���k�����s��ݙ�\s/{��-�48��	m�e�[����{Y�^�BF�am��6ݭ����.�J��=�$�����9�3�r��i��ٸ��jɮ^�3-hEЊv�+�6�=��Y0MF�	�Q�����X[��۶��3b���̚�%�vݚ�jE�3%$]�Ev�+�#��Kk�y5�����#�s����q)q.�w���кSa�k��" ��"ʰu�a*l۝vj�$a�Q*vϜ{��w5m��M�ɆggZfKƃf�iM��k�x�j�^N�7m\��A�ӺK��<�i:z�v�ol���!F�{O�ZaJ���E�룅��,�q��8o'bktx�=�p����x�I�[Kv���9r]�ڷ`riu�Kgd,bI`�X۞���u��s�: ��I��ԃj�!o7�YbrA�Fe.]�n���<c��4�O]h�@��Y�猃cR�<��OXx�\s�p�=kț����9���ߝc}�<v����uÆ���H`W��\p��M���p�FcmKv��f17c�7c������E�/c���p�e8�a�M�0j�Jq�sq����è�,\O��&hlۥ�D#�m!-p�BƳFk*ڄ�iiX�z�wX�[��2��R��:K&N�f�^^�����ך�ز�t��M�xL=�Ǎ�����m�pB�5����`���om�x�Ś�Nca�&�h����pq<�0%��&=vq6�-gQ�!:ڼ��na�gns��&G<�-��3��`�:8��<r�����[�V ��ݢx9z旝cu���1���3���B1�]�������mܻ^�&ݮ;s��d�ź�:+^(�/4k<Iťz�m�s��v{���-��-��S��=V�=9��]	t���=kk'=`��l*���SaP�a��uԺD������E\�.�&�1�b��i����aihB��ݣ.�%�46�,�Ӓ�6î��nc8,�#B�ۮ�ӓ�k�C(�a��h��H;XÔc��FU�k"��JH�X���6<��Q�)B���"*����6��ic⥐�ah-��-��E�iTe������07缉���x{M���x[)d��+�maF�(�V�ehR�5�ë%#AHW���iRn"� T�)*���c�_�����:�6�r&�-;cm�I�ZL�s�ہ�� �6��E�Y6�o���}|#e�>A���R�����^�!��Z�m�Ӫ>��ӈ/Ũ�1��p������}����Dp�.S�.I�#��+�^�Ƽ�d�㳊��"��@�p��� �����}i�O�W�:�?��ɡ7�y���kD��=�� ���Nd�H;/7��4V���8�}��k�9}|���Te]�� �Bl����\7����3`m{2(���G2&��ب�C��6��d��j��j��^#�9��9�M��ʋ".L3!B�bR��f�aW�q�\ň�4ԍz��:�feհ��f��Sν}��̄��/Lu錨\'x��N���#�,�̽~��*��#�P��-8�Z�}i�3Ԗ�㖟f��=�{}%'��G�!���1������+���-I=��Ӝλ�9�o'��O�B���rwV�8�>�h��{o$DF��M�|��v59ήU�f�e]��A;Ј"������ݛ1�t)�Vr|+ߎ,ił҇֜�����Rt�9��j���Aב̄#1�C����{��J�<A�"3a����^���ç���4MLw� ���F�y��s�ݱR(�B��� NdA��ȥϙ11��+kEt�u9쮊�3b���Z� ���#2��m��xv+�������{��q�h\�چZF�r�(��y:GXܷBggN�(��`��	\S��I��~���e��^ �s !:.��;�l!�f��A;��X���yy��� Fd"�d"*�o�����`����br�L���jc��@@�A��1CMA�w "7P@���3�̄A�bq�!�2��T��[PO^��6jEB=U����l���k����|{�~�*��&�s��R	Vެ��fy�/��i���w�ϫ�G�ݿ�����jȸ��@�m�}�̊"4��O.o��Jx���yx�@@O��z�m��`�\�;���W�S5u�8;�X����X�w��f�a��kF�#g�J�h�A�x`M��C�#B���c��`�3,��ub.�F���r�W�䤰�-�R؝�)s6Ԥ���;wh�یv�i�X�eMYXRܿ|e��#e����D3B��[<�E��5�d\G��`�1l��Y�"�3ԡ��V,�0N,#ZH�]�O��?*}���v��p]�n-����1)w� �@�9��\6lO��@;�{!x�3�@��1��}[.�uf�;����87L���&�8���[A�@��x�����'Y�z:�����s!�^��g���&�eY���+9�'<=�j[�/��^9��$�a� �}���Dwp��v=������`ۥ��l^q=��s�= �9أ�8k���VAp��1¾_X-(}i�Yj�-1��j�~�T~/.̄��G^odNً�`�\�z Xב̄A�BYqx����/�s����V�:2���3`�K&Ce�wN�#�F:yɃ�Y�~^�c����h"3 ��ip����;�.L��EɻQ�!Lf�d"\��"	̀��s P\^�e����������/���7VEDq��/wDfFć$å�hR�I�";��#�ÁQ2}W�BD���F#��OY��`�\��ހ�8ב̅�b��V��n��EF7`//ax������=9<;��\�5S}�T>"�A��7z u
v ��3�s�Ux�3�! �w�u5�|8�e�Y��ւ#2��`��#�rE
$c�}Vv5�E3:E�F��q��(�bm`1S;DD�t1�c�;�렛�1�w��vē4������0W�<�h@��6!��� [���$�q�e�6n���ѵ5f��fCe��lO����y�#�q�sn���f��6����&N.�ٗ�
d�5�V���C ��JJS�+Qn��ئ�e,�])R6��u�U]`��Fs����'���,�C��Qbݰd{JB\�u��S����ڇ�ݺ��1<Îz�>Zʉѹ��Y��-m�uE�ʡ�]�͹������\U掴�ݳƺ1=z�i�۬����v�%f���;�w��K� ���G�̀�;f!�w�eX�3R� ��$�NU�:�Yiy wab��s#�F^������Wh�F�^>6К��vmpf��Lp �����Ge��^ZpiYt� __Z�-,`�Տ�����#w9W�yqVEDpw�G���̄�b�B>'��p;�r.�5ոCh sax�s /OY�y��3l��`�\��ހ����)�\pW[�W~������'2<�@��!֞��U���d�LwKIgx�Tw�'� A�2>́H��Ԟ\�T��]c^ZLm��81)�qNA�.�b2ͥ�k@�(����@�� ]���2f �5ѝ=N:/��yqVEDx�b�-������A s!9��3�}��-'}����d9�2� �s�kY
SZ����?�^I�A|b��5�4��P�K^-l�J����{?`�#yzv�E�ރ�Flv�)r���y���P����#6�B�`�V!����j�-^�ݛ�����OK|��8�{� Cp̏ s �]cZM,�Օ��G�f ���t�8��%�Ҹ���2�DX���@�B��@�G��d ��!\#C;�hq�|b.�ƌ�S|r*���1��D���'+��P�rv�7P�����%l�N�Z3�Z��kgv9z�K\/<b�Z���e��e������>#1	5���6��!o����F-�n����V@�A�A�^ �����s��7N��mC����S���"^]+�Q �B�Z2)��O��/.A��� C1{2+���wQ�;���3E�G#^ͽ~��[�{7�;��o�ǯ��
<��ЂU�����3t�^?b;
�V�m׵�!'��	��v-����h��9R�	Aב̄A�A3!Q��Te�{1� ���Q��bM.�w�����ޛ��w�t�+f�/1�6hy�b1��X����{��;��̏dݮ���Kz�ᲄ�kgk#�7H�wQp*#�'zZ��� ��D��}��-��PK!��"���U3�ő.�]���n4�f�ꋰMz�6i��;�_�H���~|�d*�D]��ʛ�PE.�[s��d��HΏ �y���>9��i�o{���Ȟ�8-��Rh�sjkG	�M�G@=� ��@�E��cv�:�Ր���@�G��{��3�LG�8B�ڦ����͝�>��h ̄�  o!x��cx������}|��=G%و�Ӽ5�7�"��\ �@@�wz9�a^����@�I�E<@E{|���;Ȯf5y�p�6�luܚS	I���P���cEB����PqK.�_B�T��f@Da��v���~聛��˛���V���8O(�p�d"	Æ�-�zt½�.�
`�0 wF��M��mf�{��"�b�mt,<�{8ۉ�h��ۜ����eˎ�V"ݗ��=;��u�8���X�h��ˇuA� Fl �b�B �� W%]}��D�{z,��6�".���e]tdT�@���<�̈�۵��w]�0$YM�"�@fE�,蕄vc7���Z��;-�eTw� �@@��h s!9�eG��:٭���W����@�M[����s{�nn-
��}�3��z�nb�dV@cAx�^ ��sF�2{HK���f�I���r3�5ik�'����x�B�&�x]��#5�Y�#�4|�������b�҈c�?]�p�?C����=
�W�]9��XY-U�)$6j����Ƭ�a�N1E�{�����ܼ�;���q���O�`7k����v�E��!�j���#�Z�rU!]�s�k�(\C�Yӂ�;(�8���շ&���NWqR��.N.۶7l	�g�ko`��B�שUm�y��.yDGi�>et3Ĳ�m�\b8֦G�w]^wEi�t��c��7���r�m�'sq���tc.x��M�c�����X�a���4s����g�&�4θ�� :Og�v�H�j�� ��f#N���g���� �D�� W�^�\���]�M���"�n=g��s��O�
 �h#��2 ̤9�"���(�Q�����@�4&�����{�7�Dq�B#\Fdk��uچ�A]�� � ��d '2��;�(GDGullۈ�$Er�t �����^fB �b�Y.1�7��2(����K���˞W�'�sq�Ot ��;�
�����A퀁�dA�@fEm&�"��u��5����m�šQ�A=��p(y fG�tv8�<����l瓞��;f�/^m4�ɹ����v_A�:oUZ��uǕ:�E��7e��Kw�U����m�7��$��t�-H��v�����&�R�n�#��q7��;�Z}8M��[�`�A��7lU�U��R��թ;���}s��F�ۀ���"���8?,&����̘� .���ٕ4:7b+e���m�n �z�����:k:�8ew���p �����de�}�Rs0Dq�8���0}j�`���B���6z�2nM���&��Z��B#\Fd }�̊E,ên/�T���O�T�L��`���֜_� �g{���(��tGs��[7'^�ƥ�:<�r��@�2f@DfE<�Οv�ƀ�d;�+j�Ƴu��sq�;��n=� f@jOqћ\�T�&UF,�j�n]q\͞v�vT&��`�2��l���)� À����̄̀������m�Šn8\����$��3��s� F�Gِ̄A�̀�D��/�p�k��j�	�q]�M�َWD������^9�z��b�e}F���D�eZ!��i�Ռw���H0k��R\��x�u�4R	�V���A�,�tj�u/y�
ܞ|�9^x���Im@i&A�����=)!�dK��kLS�G{���꽔�~}`�f2�N�;5��$���l�/���'�	�[8ۥh��+��gM��w7\�6-�*͘u{b���駠�����U�
�f�0�>봻r���rx�������o���?n�1M���ӗ��/%Լ�3�%����n�6�N�j&�����$ه��4��zcYZң3��/�e74W5�0y�5��ӯ�*�����z��!�ZemFM�wv"4���漽[Y�bW}#0�����9zy.C��/<1�_l�6@��#X������jݛx����8����7S�d��v�>7�t��ՊA��8u��y{���&�A��;�7W���@`�s�v�n�ar�y��0}�kj����2�C���u��q��?mE\�����`D�v�+u�o���zB�Fi����G�L�Oez�{vP��v�P�s��0V��{�	�f؃��Xf������ ��x�-��Y<���nÈy��Ʈ����P�h3��_v���<���x����qs(�h;����6rU�nu-NL�2��s8��п8��������{(��O��<}�{�)��Qi�<�&���U�]��[���w��-�Z�C}�N�z���)�@��:����J�{Z8���Mۻ�t�iujZܜ�2�L���)�u��=d�`�4�;�՞ƽ/�nfQ������h��H�Q(F����N�������/m�yךB�V�(,oV�	e���vQ�ִL����Y�g�v]���剄6�ki���ܶ�,�;�l�0���[<�'���s46ۭ���ՓX��i�[��mm���[,���s��=7fC-,�<���8�Gsnk!m�)��[��ֶs,�l�m�ڛQD��[V�Ngk7e�m��IͳB�h������іF���{ix���+n�Xnmml֯;^[[ ���vfZڵ�Y�-��[8�N�lrm�m�L۷�$۶�����l�g-�mF��y�[��[i@AX�n͙�bf��8'۱�em��[vr�M�V���vJ�6����;4�l�nG[W�,@�0�#	8N@��:�}Y�<��~��@���i �ђ�����%$9ˆ�
A@̢�|!I ��p	I�e�� �?Z�~�̯k ��ZA�Q
H.�wH)��s�f�%$�- �����_���Ɲ澯�$�vaI%Sz�l�I��}?[ԫ3�>�?	#���<	�K�R
A�C=P�At0)2�M$P2S�wCBJH,+2ᤂ�L)2�I�����M�=��Ad��~���k��U�g���ϵ^�$��I!R���H:
!I�]�R
h@��f�JH	 7�O�MR���fxը����0Z��s6��['7M�z; �\d�e���Mih�C��wa�aI%SeB�
A@��i��i ��p4URʆ���k��G�g�W�տ���@���i�
H,wg�?����y'����R�rᤂ�L);E�Ѕ$JNe�II�e�$���E�Q
H-����{�y�����R�l�%$*{�i �����w����n���_�������
H)��P�M2�
�H) ��py�g߹�7[=�)�Cܨi �`R2�H)�����p4$��³.H,4F��E���Y(}�� 9��f:�C� ��WL߾yZ�{<|�X_�:H)�����$��� ��
a�P���P�C2�$aI̻F�Ro��~�}[��ߴS^���?n�l��RA@�贂��I���jU<G�q�$x5s��?W/���5��~��@���^���R	�>�Y͊_B��0�}v�'�	4Np�����ó��@�u����]�ޗG�����T&�^�o�gn�eu�'t�e�s&�>N���rA"4��I6U����C�)�E��B�%2�e@���XfP|�
B��̢��!I̨�S@�L3*���]w����k}�6&�T�c���S�b�\ q�=�>� � �˄-	��`M����׿��pg� \̐a� �P�@ `��6�0�Q�����&�#�Φ�Ya6��ΓY'�FΖ΋82S�TCBJH,(7ۆ�0��-&�) �2�Z������o�>�߯gO��A��AHkY�8��o�~��pڢ�h�$��p4�R�l���
e�Xi�$2�Q��
JB�fT- ��r����~H,i �ʁi ��T- �~�\|k��羿q����@��-=) ��J{�hhII�Ne�I��Re�~�����3������>�|�Y9Nv�Z������ �r�H:��Z̸H)�
a�P�i��@�p$�|:�wp�EGd���9�W����]����<�I%!L=څ����r�$���P- �T3*H.��3(��$]}�����~���'z�ZRAaF�p�Aa�� g���) �2�Z��m���㵾���~��>H,/��I!EP��uD) ������{��`q ��)�7P�i��
�}F�) ��a������d�e$�- �44�\ʁ��_�꯿w���)EC]�I�t�xO{��;�M}�8�+ ">) ��J{�hi%$ʅ��)2�H)�C)̨��/��|{�����M�RN��3�Gi���������(��7JU��n���.���&�K��ioɃ��=�6���1��L�Td���&�;v��W%�{���d@�M�]��;���/��1K�]J���2��It8��Ʀ�zm��:p��k��N��UƧZC����9����l�k%�M��ûv�hv�֨6���l%-�������[pu ,��ftŹ΁�ld;[�9�w���ps����|��݀�
+��.��1i�ttC[�����S��[S��mg:��MpwJFT6��k�Vi���E��c�bAa����AHUP��u(�$��� ��g̔�P�"<	�y��M��尞+�����-��<
K�~~�~3a�7څ�����i�Ѥ��.�j���h*�$L
@̢�Q�*2S�wCI) �����ug�솒���Qi4!I��O{w@���j��x�o�z�������_��R�ޢ���$��� ��
a�P�]v���s�<�$� �{tZAH)��c
H))
aܨ[&�RA@̢�M$2��Rʅ����~����~���ߩ|Lѯ��[�M}�8�2�"<	��J{�
RAaG2ᤂ�Q� fQi �i��]�P4%$�I!�����[�^N�<�E���\�kP��)�9P�i��
!�F�~���������ϯ���>H-���Rx�Sv�l�e$�ٿ�<��w���xm �:�A{�
AH:
��P�At0)2�M�R�wCQ%$3.H,43(���ݽӣ�~���}��Ad��owpO��U�s��}��_���$�A�I!EP��R
At�j�Rʅ��JH(P�eH,=bw��������g�WF�Ͳ�
B����.�H���[��z�2�ԸKjUT�i֮� �n��Ru
a��d�I~��Q���]��TAH5P̨i �?}��]y��w�_+?|k��uQi �=yV�9�����]��������XW�p�Aa���E�Ѕ$��]�P4��XfPht�RTe�tQ�M⏃��/�(\�rڅU|$�{��5�k᱂��N*/f��V}�(m��#�3F�aDT�=�V�m�u�U꜍�5��ΐ��Q��Ol@s� ��
a��[5) �Hs�$�|'�o��]|�|6�T��dx�\ ���ݨ[&�I���Q���]������ίZ���w%CT4�]
@��ZAH,�%;˸
AH,4f\4�XhaH�ZMD) �S)̻��wh|k��P���C���c���X>G�>Q��!�=�- ��Z�kP��XfT-�2RAB�̣I��RAs.�@
K���i��~�����z�l�I��4�R
Aw�URT3*H.�}��]y������������H)�����p5��XQ���v����R��i4!I��S�]�P4��XfPi�AHUP�ZAH)��֠) �̨[>�e[���[��N�H����O��g���j����wU�C�����
H)(��B�42�
�H,4�\˸� ��fT4�\�D���ݿY��{����UNz�ru�������]"�V�nu�ԛ��t���UkSM�`mwE�) ��)̻�����XW�ᤂ�P3(���Y>e9�p{m}~�u���u_~������:H)�=��n��~�� ��ZA�D) ���P��Xw�g̔�P��4�R
As.��
Aa�P�M���\�¾�k�����H,�$���S���dG�lxI���h��/�����/ށ��E��
H,���z�����XQ̸i ��
@̢�_17wU��z}z�u �|2���II�n�Q�AHQT9E�J!I��j�SQ�fT-�JH n#�������E�9T�u�c�9==c�xs���d>眰q�������fCCs���4!btݹ�����W��~CJ�����b����]镟~��^���݇�0����)��P�M) �s�ZA`i���]��Q �̨ZAt���-4�I������o��{���$��½��I�����i4�$��]�P5�6���{�~�z������ߨ=$�U�QiTB�f}��}�k}u��R
~@��B٨�I}��0���]��RAIHSʅ�i��P*fY�����As.�W:?[���)��{P�<	�϶�FԾ��N�������R<�O�wH)��ˆ�
A@̢�}) �2��]���=y����?��;L,ML�Ck)j+�۵�uG5�s������T����i�N��Z���Aa�A����P>��R
Atw�� ��g̔�P�3(�Aa��竾�߾�}�~��^���݇�RAOw}��O�Q�Uq�q�� �]ǂ>�����S���AH)�]�����h�fT4�]0)2�M�R�wCI) �j�����k��15��I�����-&����C)�Z��/��vW�Z��Lp�<	�>$�J�=�- ��Z�kP��@��g?;������\��
��H,40���n�)&��9P�M) �fQi����wH)�eB�[���N����d^(���-�F����\G���W�Ạ��U�;��ݖe}��+[��>�� �/ oa�	��ޭ�ස�uU4"��t }�s�xq	]\wˠT�AS��dJ�E0Z��3�+V9�S;����㞲�F���-�g���%���#`FnSW#jb��:of��a{������{i��{ !�dy�Fb�Ds��¾=�Ӯy�)�o�}LP���=� �hȢ�B�-�әR�zTDj2�JIF�5qs@�f��Ɨа�����#Ō�)�y�!��u��'r�-��Fd �UOiDuf��Tk�
��;��n�3��+#��>2���d��-�\o�#1	���N��zyJ����=��@fA�?��̬����������8�e��K�}r���\FV���1YT�esب�b��/w@@�1�3"�̀3"�GI���;�����p���AUn҈�ͻ�=�0�ۨ�OtN�&b�y��8�Dw`"3 /�����̌���<T�t葠U ��@{[W�w�R���8���̀b���L9vo-������"�ѯR� �fȼByO3�7q���w<!;����Mm:8V�ZӇ6�A�|��^��$��x"{=��s�܃��\��`t~��:�Ĵ�'tf�;�u slg��U7]���\n����۔�F����v�D,[0F0&лk��6���N�xݺ�
Y�i����Q�)]��b�E&2ۓ��h����	�I�׷0�������lK2�'MX��m46	[KF��&M�v,l(]�X���W����L>����º(������v	Zn�X��6c��t5��矹�k�os`<�<n̈́�iH��dt�k��P6�,k�ީ�����> ��̄>9�+l���-���7lP���]8�O@�b��yf �������$h�x"�T�`��@�Wuٵ|'�cN�GOt/�"�#o`�y�D<AtA�b2(����{{�����f⪘���O�Ǖ4�8�B ���K�f �d F5�/ڙ�ǥ�����i_7�>�~�V��jر3���Փ2R��:����^ّ�Ȣb�2m��T�*��"Py�%D�ھ���'n��>#z���DFdoc�Vs��z6���~S����*2���X�/�;�m؟m��WT��D*�N�H��v��{�"��X�u,��/O^��[Wç����k�P��1���o���DM ����㘽�����{� ��^L�و�z臏�p3eڠ�h�ee�l0�4(ċs��}s�X��lTڑxP��lDƷ�7�rwJ�;[�xmп��#�W����Z;r*ر3�{� |�̉\fcrzC�܂�>�Az�y{1�*<Fb8��Lʎ�͢�k6�
����Q��OC��B���@��dP�پ�d�y}�3���m:�����uAzֻ"��B���El/���̄'2 ��̅N�:N��z�_f�h�Ȭb��x�K��V"݊oF������i�&�[�!�6��d�'*F.oNN�Wc.��c�����A�ڄE�� P�AMwQR��v�;�1�1vꑺ0(� p�΄'2#1	̀�E1�rUSoL�x�Ǔ����۾��U�53B�;�w��A Fd<Q�m�m{j(x�6��d� �r��1#3�&e��F�=/����Q���O�;��3�`�N��+R���
\fCv2�=jI�Z�U�������4u��ۑXŅ? AAmy�^�A�0z��N�s]�@�������MF��ِ�F��w1�;�I?.o��(��i��|��^@������̇7��07�lXhMfyo:�ӴU嚙�uA�ބ>m���^�צn���;m�-�3(�0�A�Q���8��/&�9{nS�m��o:�&��b3sq���{�E��dQ�@B�l��=�;r/����t�q�[>�V���^G2�9�"3!Nd"�v<q9����p�>#u4������|4�K�� ��E�̊yvj�-��;�:F�]@^� ^�@fE}����ͪe*�H��+��7��^Y��P��Cp�̀��B!2"*�Ƙ���}�݄A9��tzrOi��k4XS�{`"3��6&��(���JӛM)1+�˫R��%h��ؼ5Qu�1�b�Թ��M4��)<����N巻��1;۵o'(Ū�u=��έ�B�[X��}���W/|p�#u�3!Ndy{1�m,��רcAzig(��;�"o��e��Ol��"�'2�\m;[��k���]vϮ�vstf����ue�B.j:es��=7N��:���K�Q`��Kw�����ny>޼�J���Л�n�1+;��r/���Q��b�Bo#�K��!�Qͨ�=}�
�cg����v�E�<�=�k��D�oO�܉��8Ā̀/"��b�6c҈��td��Q9��y{�f]�q����R�`��Zͣ��p�@^8�`�y�@�3����}y�&�r̩�7�{��EZ��o1�e@�2�@^ �/fDD^�Qڣ��N��c��7e��f�wk4XS�}��!�Ұ`�V�ｯ�x�G#{��׎~�\ U�ULq�&�M4���k�m�4J�����Umⵅ�lE��o��ݞkbB�+h��-{������~�߻^�rv���QZ��6����t.9����D=��5�l�eP�'�X��gu���ӈح�q���e��f6/)S�!~	����o��A3�����B�퍘�*�B��5��kq\ʎv�O�����ܸ��dSޭ�0a��Ǩ.ʖq�{��Y����VX����I��lèo%�L]���G_n2w�)��ǁN�;���ӯ4�*L3�$���MH�s%C�ڝ���資wf���r�1QT����޾Ӷrg}�����I���x���;!�{�|(>��ɥ��k���h�}x�d�'�6\�{�^��hl��זp��<���ѽX�/B��>+�^�m���1{��}�<]��m��1�w���b%�.;hZٸ�q��ev�՞ũ^�?rX�=��g<�/��%�\5��t^�ܘV1=�L*xr"��kL�����מ�{͟EȎ�)�!?E/�3�=�j�Nzb�75C���akU{��gBE��2j��^��f];5�ɵr,)���Z�w�dKLo  r�5�^��3ѿz�{ڗN�]�q�||@p[��	���\%"�K��õ �^��2[��gdC(��*Y+$��9`c=�fz��<��w�e:�����Vk�'����^'���R~ո"�s��o\�.P`�������\��uZ�=�����V�28�oW#��>@  N|pa5�@�kK�gb� ����kT�۰�a�P�ˎ�1h��l�vi��z�!mdF�,������y�ms�ٶp���)�{��s�����3�4ֶ[��m�36�rY�Z��v�L�3X���@������m��k�z�֜[ck(��Mamv�-�^a�Y������u�m{�qM�+-/m����%���b�T̷��	, K��
fݎݩ��#;��s�v��]����YZ[g=�=�h�E��É�6m$�l�ͱi������i��-km,ɶok<��sl�3h+�̬�[c4��:��ݜ[`�/k�ͫt��ޖ�t��Im��5i���)��;2�ó�f��ᴼ���ݹ�is۳̭8�Z��ۍ���f]�0M�����YѶ�-�Y^����%���`��uikbq��s�v�8�l�kJ��»)�kT�ilM��P�Ye"��pl�(U��dޞvL� N��M�G\��
�A�s�E�z�Jrǁ�dx�ֳ���ꋪ�Uƌn�sI�z�0Il�ڸd^7;���#ɪ��%���Pu2odm�j�ӎ����� ��r�w:{�6��<DY����K�m��B��qqp6�/޻f�3qP�F�C�En�d搷ЇoY\�Pm��2{m�C� us'[�0{-�F��d�BH�����۵n9�89��cVԳE]ed%�8M0W)Z1�S#�mڰq�Ф2ީ���˶q,��hJ�;��]�;]\�۪��5ӶM�5]��S�d�k;���ps�MY���N�zF��.�Y�Kn��KeA�--ێ���:�,S�{pǞ�[`F`��nJ�B2�l̶_���KG�f�,�BrmX��M��m.�ۮ�g��<ky�X4Y�������9q<�#�n�z4%=!��֝r���Wj�h�ƞs<n��auu�cs9-��u@����׌��sM�n��L\�8�厹[�����o��ۉ��qv��O�n��q�xz9�`H�'��lk(sS���4P��d�.ڈ*6�t'�-;q�c���.���N9�4���Ѵ�=cr��v<�B�/]�$=��8g�h��s%:ǵn��0�h���:�L���91��y�9�$�m��3����s���Z�CE�@��)kJ�@�]G[�uv��z�����gt�9�7g�j��6ɣ��{ﭶ��㚹�#ӹ�b���L���=u�fKn�f��[���W��]tsҜ��:��n;"d&�}�.��k�ܘ��4�k��5��xШ�ܔ�����L�;:�grZ�y��%�I�b�V�r �J�f�Pu՘܎�1���d<�st>#���Kt(��:�	c=ǆ��b�O@�f��R^��1#����']�k'#�r�g�C�6�;-�u[P���������sQ�U�]�>#n��s��e��Ǜ�n;<t�u��������sW��҆���j��9M�8�[����ﻢ�F8��b����[y��T��.���'���n���1f�͗V�E�c�����X�҉���Ńt@�;(%�;I� ���o^֮ɸE���B&��[v9��e����-{\`�6j5���A���G>}��_�V��kcq��`�,Lk ��zcB������n��Z��QBb?A�,�#2>#1
5�=}��*�ٲZ��;"1uM[7�;���A��2f%���L#W��Ӫ�n#<�9��F�'wϯ;���Y�6&�Az�F�v,o\(��5�ᴂ�/�ç�f �d"#219��'B��F�:'4s:]\�
�p�As!3 #�Ć�ʧeǭ���{2�EoDOgs�ʾ�l��;��@��tv;Y�o�v����"#�"3y�+�27��7G�V���Dn�^w	���*o�}���D�@�1㘆Q��ۋE���\��l�4/��9���y��hюs�v%�v���L^����ǌG@`2��dQ�UV��k<]\�
��ޏk5�� A�^@�B��#2���Z�[[�za੢�����ٛ�8af���x��e�ع���z�it3��m�:���`�=V��o�w��fn������< ��[ﾀ�+~���y�N_{6�ɎϠ"h s#��k���l-L�/ Kp�^@�B �1y�dA���4o�3�Mܼ)M�~���h��Zouq��;�\L�'1fN@�3Fv �H ^� ���S�2���w9�¾{` EOv�Βm��ڥ�7��"�fBs!}��#2,��ͫ(:��=�<Ay�툝��.k8a�7��y�@�^̊��g'6Wu[ɓ]���x b'Ȓ��F �Be,�N�B�O[������x&ZҔ��Jw��O%�p���A	{������6��6&�E�伇1+'��3�/��d�0Zq`��rj[�v���QР �UOp�N�h}N^�
� OlA�j��̅�qv��	H˔"r���2 ����Glqq�/�YTc;�����z����2Us��X��50�Te�b7{7���MD4��}��F^�*������N�i��uC�}1�(T�CFB���Y��� ]U7ݴ���m�� n@��A�@�s �AU^Ȩˮ鬣��q���n �!;|�}��u
�WBn8�ޅ�3»8�ѹ����B�p� �n�.�F�F9�ظ�G=w�]/
�ѡ�U9z,+��f� s#�f �.��īi�
=����F�!A*$(]n�Z�� �����Q�ê�%,�fl�������|3�fB>>�!Q]�D���/;ۆq���Úk�U���D��}�3���k):�T:��1d�%�(�ov��WBn8��"�Ax�����˂}^}h#]�2 � �d A2��ݽ�<1�wC�/+�
�ѡ�U9z,+��� ���d/|3�G�}7]i�[w/ax�2�����R�f�{�y����;���ދ��������T��xm5!�|�g�}=�����m�}<RE����n�Ov7��ϭ����q\#Ee�J�A��lPg�� ߯��A�����f/ s#b��r���)�(9ZݥSآꂸ���^ �X�e�`�Z�A:�@�3�x�"u�����Sqfִº$ |\R	9-q��pLd	�cz!��dC��B ��Ump�.xhg������w[�/j�0v�b�2وȢ9����Q�[�������݈���6�fÉʏw�8�A�Diq�"��k`��q����-Y�wX>`1�D��*��ʙ�QuA\q�@�mr҇�2Ջ�iC=�z�"[o������F�À��n�e�ta�v�E�p8�������o�p���و Ȁ 3@�3f�(ι���}�d]�D�ފSo�l8�����!�2�2|⦔G�r�@�14�N�����f0M�\V�3�dd�*��x�nE�x�͇���<-|�.
{y�6Ͱf+�i������+.7]��m����\tV4!n���=Y�d{pn��Mnw\��s�k��6��.�:ǧ��.w����^�}v��݁�>z��8�����tr��nS.`�s+<����#�xvz������ޭm���Fu�Y���{yh�B� -�[Q3���:�z�i�RY9}]����&\�� J,�a�u ���#-3p�5�E�F�����ߥ����GB�h��MGv��[n���3��5Ý���
�!v,t����~�-��2��4����+^����(��+��:���'l>��A�^���1s!H��A��:7i����xnC���_V����f�
� A퀈 �̉��M�A���f@^>�Ax� � �8m1���ӡ:N��Z�����k?�`�e��A�G�p�2��@��Y[=����@�8}�A�)wr�ݨ���t,�@ �DK���e�`�6�#�d/f@^ ��̉,<u��Ց#�.%V�/ !���poV����f�
�{`"my���F��ƍ��O_3�ڵ�4
7@#]���i����Н��dVW۝q�e٪3���.<��������LȠ}�zb�b'��R��7��r��u���������3�	�6�Nd�Hs  C�&������`�Kc2��L ��I݀��4<�O+'��X�4ݕ��K�
ʡ�ɺK�U�v�ʋ>�;e����ڸ�mU��N�fm��~���&��7� F�	ێ��\ۨS=�t.c��B���ȋ쾐�_��V!_;��_O�Zsk��w{��K)��}w�®���@���9��1Fd B��7�ٮȍ� ���΀�BMwDO_�7�oS�ʎ ��Ԫ�/!��f�� ̤�dFdy��t^�������������7r.c�AzqFd#㘽�&�ɂ�e�e��	]11bB(�2$�i`�q����Բ����l�\�Z]�M4�\c�|>Y`��,<~���Zq|�z�ߟ�t���r�L�+���܀�9� Fd/A̅�FL�(��O�`���jkz"z��Lލ�N&�=�: ��2#��B��{pQ�+ #n C1|��`�j���W�wߵ���	��b[��Յi�n|Ҽl�K4��!{�z������y�o�r=��o����y�yo�3��/W��r<K��?�>ϰ��y��O;����D��#2>9� s#�vϮ�uOd �3�@�B ��@^��WmE,5�sE\ 󀈘ؤvm���{c��W�̄A�iC��-8wT�����/��R�Q=�z���ާU f���fG��9�{۾�JNθY��a'~At���x��<	:1ӝ/OcY��s�eB�h�0�s�w� h��̊����{�n�L�;��j8ª�hw9�=��/7!f ���9�e�ٻ_�߼�>�����۵R��Y�w� �c@fG2L@�q#HT�D=�'6 � ���|s�A�����E҉}�z�mjq5Q� ���@�� s#��@@���;j�?Dө�;�1H7KȽ���AK;� v�ݘ��w".8A}�v�/�ﯸ�;͇��;�]��F��vχ�����Ք۶ߍ���%���e�{�#ف�(���{��RcJ�N����}E��Xo+�N�˃�ճ{��̀�s#l���T�e�W�b��ymTa��w���D�y�@s̙{e��?42,bEֶ�鈶]*���]͘M�u�¼�bl�����e���Y~ �̅�㘅Tw�W�˕�h�Ր���8�6^��­�W�7#�{!	������[�PSSLj�늘g#˹�㸢n�ى��fע��D�#���6x�59�&PGn �Fl"Z����e�E�j��.���k��W�>ڨôj�P����A 〼s#��1xfPCf���O� �Ax��� *���vr�u\+ud*��lzK�ʹ��\1̫9ʸ���Ac��n�O2;Aάs�h/[Az�zT2��Е3�u|_�w��������5B{^�ߗ���({�{�'�,��*/ͪT������1$.X�diP�6��L4��U�RU�.#l�zP\�{�g��� ��|��D�4a�	l����ݮ�ݘ�X��9�u��E�Bl�ƛ0R4���ma c�;i�t7�2;��	�>�\U��H�
�'��JA�n�$3[.�)���n'�ϋԁΗ�dzs<�M�ZQ q�W�Cd��W ��C=��Z@:�ZGm��=^z�:�n�������8�Hè7/N��c�Tr�n��+O�6玮�q�G�w����|���T�k����.�]�\�F�`ãv��� �4��v�a3�f=���|�6~�F�@�̅[خFqݩ�訫�Bk�B�w�mD ���/s@�1�d"73"��\1£��͵�!U�W\w+��OV%U�Gl"ms#��a���r�R݁�b "6#@�p�'2 �B ���닶N��E��*P�7�;�W���_B �A����x��#9Z��v��s""=y���D3!
}�Ύ٘Υz$Uw�><�"��@�
�8YjY}����^��9�嘂>�2`�E��y���KM��W8���/U�UA�#� ��{2(3"�����={�mo�Z��K�V��s��n0��t! �
�]�L��� Х������ ���́B�F%�5��3�ez/�W���b1(`D��{K�ًّ@�Fd D�l��"�jc��^pqR����f���r}�g�8ߨ��8�庫f�ȖS,VM�����z*�H��1�#u�]�H���6�< ���P�x�Ѐ ��B�bC3�홌�QW�ET�Adnb��!���^�`�X0e��K�O�s�o����JWl���^�J�8|GtycA�
"&�S���U_q^j��E��q���́=щr�rf{�E��_BJ�͛�u|b9H�w%��fEx�Fd Fałӱ�����v�����<�[���9Ԣ�D��^�x���d A�NK��7P�ݼ���"!B�	2f4����:ݗq���L�Wkfk+q�-P�Gv@����[���͠�}���}���[�Wd���^ܥUzc�=�YL�����: ��iǂӋ{��|�?\pSl??F�'z1.D��6��a� �z/���۳e_95�~7�S
�r�##�jf@^9��8<���|��8}��~�+�o��tZʅ�<����b
�8؉+n�K�̍GX+w2&��(��*ٓ=�2$5J2{={�9}�9����=WC��R�J���{gH58j����8�eg�="���>��>���V�65�����=&q^��i��}ȮگsK��P��v-c'��ٽ�V��?5����\Z^��V�IOf0��ה�q���ЗbUdo�b����R���u�+��]6�ї�]V]`ʭٲRJ]����;!��W�J�N{/nݙ�隴˄�cm��u/���{ܽw�����/r��w|�D�6úQ�$����k�;b�ae������Y+oOS�u��\p�L�Yx8@��K_#����7���ΰ3�{���vr����r��i��6mj&T��q=�[K1Py�}��ji�sf�4@�5�q��sa�˞����<|^�4���;��I��	�)�O-�B_t����| �/Z���eݙ��}��f�і������r��,�͛t,���!�<+ފ_"y��ug�����<�b�<�e����,��͞��޶��`*���I����
W��v�^�{7���k��Kv���`�4���ot]��Vu�܃�V,���2Ž�z}�{��oYG^Nة;:���Jvv�l&���w0n��A�;�y1��h�V��ר���3��=��N�i4{��È8�h��W�{���P���=$qL�u{�"x6W��������=��ü�u�ع�Nu���s�{J���Me��Ooc7ﱊO� a@��Af���Ί�L��w)�Ft؜��h�����q�Kj#)�Y-�m�c#��%;4�#�3��=�u!99�7�nŖl�a�̂�k;2�:6�(BC�1�ܭ�Aݵ��3����;kE9$A�Dv՛tGv[l5�{ΖZ���gY�u�6����c�Yp�Z�a!dvDM�l�;6��78I�����m�PE{{�Zu6���:��g�������m��v�m��L3�:C�3�e�:�'-��p6�q�[�֒I�m�6�)e��Y�8��Ea���+�\S�BVY��D���lr'4�Z)"qJ$x�ڱ�tN��nFբta�m�Iō��$��jV�Ռ��f;���v؈�5�� ����i@S��rrFsk���"��p�: �e���o{/nΒ8�#�/uw��ӊC����줮�H��y�^ ��!�|3Da� �/�B��7> ��#�B<o���'�r��^ܥU i��1W{F�ָ5�my8�Y��HdF!ȱ ة����I����iʂ�p�=�P�}����Ç�f v&���4`9��-_k���:���k�F�ˍq0����1ն-����,�L��]ޫU�����Fsv[�Ո �«t�F}���-M�3���[��2�w��` ��!p�9�8E�������JEQ�;����ON�+D�و��q���ͯfEKme��ꙿ��;�.";��W{�\�P��1Q��1�P�='B��+�\>=����ļFb�@�T��7D��ޭ"�뀼{!A�]�2���
'��ވ
x Od�c7����:yN�Q���u�2W}�Db���3/�c�8��с"5��5y��W��rЧ�1��n�+T�Na�	həh(�����Q��j�z��݋�Խ�ˌ��SS�3L��A˪��$�Wg�}�<�������/@md"#2W]\n�ҴS#\uYa�(�2& կQ�sؗk<[���m��6�Y�V�Jhf0�r��e�P�  d"�B��r2�Y�,)���c,�sH�����lIg/��O���J�kܧ�I+���u>����+�Z�w��  }��̋z��ՠ������yf/���c^�ۖ�U�)%eM�F��R�b*��>#���7A�Ǜw!V����8$>�Ǎ@~���~ ����r2�_EC
o��R�/v�B���5�J�rF����z�H-��Cmy��c9Mf�W=:8qP�����R���ք.����>xׯ͡��.����]�6�SʽK^��A=�la�c{��r��Ywю}���.��w�,pj/D3G�A�Mf�I��|�Qy<�����33�o����4�Ů�#���m1��)�j�nF�0h�i'���Y- ��U��:��ƽ��˹d��
bv������6�Zc��gv�HÎG����s��GFq=t�|�u��T������m2�-�ca{;�����y�k��x�G�#\���۷c��mq�.�6�6N�@�nq-���cuF��d�6h��,�\i��_߿y|P�԰�Ib��3���X�f�Lb���zs�s��m�$�	�f7�{����YwZ������r&�*�}R�#��̽������T0��f�nD�p��s ��x�A���n�z�[S�5�W���:�h���(�����h Cq�ȓ�y����!>;p��@������;��y�����dj����B
){n� 6ׯ͠�Cp��'�di�1/, �A����"|*­]R�#��D�Q1��!j��l�]j��c@.��p�$�"k���L�X�d4��hĜ���3|%
Q��S���ʹ;):L��VlZʘР���q�m�][i�v�O�������u�aq�f=����/�?i����[�\�GFt5<���(�'`m���3���/5Y�@� A�m��"�TGd�Їe�����ʂ����L���H�K��ۧOH��7��0Y%I���|�8�R��\�*�]��ε_Wu��O��o��$$����[���XU���ܪ�3�� A�}�$�f��:�Uw /9A��^@�Ԃm	���e)ձ��M��D։B�q�^�h⏋nD���<��ZH+s�k@�@�'�Ү�íTa�a7�n�1pר�r��A�%�RA��nGN`�2f3թ�<������D)� ��@@���Ȓ� A�n]�q^ܓ�����]E��d�1eݴj7B+qsr�xLZhVl�$DyL@�	z�#v<�mH ��������z$Mp�-G7^�vF:�TEl �(܉�D[� �Z��O`��<��
�į���\V�AR��df�"�V�H���m�����z�Ed  ��$7�|CnA.2,�%�����p������*�������@~��u��b��u��ǻ���lqn�9&״l	��Wuq#[�������=�G���:aw#�D)��>=� ��$��p��8-��@�R��7�{x�$%��"k��j8A}�A�����M�)r������7�p���U�� �VC£9���*�9�rq�P�]>쀈>�^@�jHn��o5u�ѷY��ˋp$���Jz��rn�+<��93Ѡ�M�mcZ��(�=�+�\}��קۨ"�||ۑ"�+���%l�*ި�1�8��;���@���t"	n ���A�n<+'z���j:��{�A���LB�ّ5�P��G�yI����[���\P�O��D�����"|[����׻o+4g��in9�+����������ԐCh |�
�_h�P �����^!�"��j�̹r�
��"f<7c���G��eT�UNS�.���Tچh_����sJ샐�PA�����i������!��ճ�Uk���Ц8VFj�"�t��]F\�ɂ1� �����y��� ��X&f\̣�c�E�f+���Z�H,ןLD�y�EȚ�Kָ N�) �Z�Z�nC��Ɋ��_������'�i�.7b(�r�on.�z���@��2Q�������%�>��,�,��n�=�iruh�T�:��.��p�"�zפ6�e�^-�$eE9��es�ѷ`Y��܉�*�w<��G���!Lpx�@�z���
��s���w�pv�O�;�"ebm� ��3:ܬ�B����"D��Ѹ��HZ� ��RF������� F�R��ϗ=�`�5 H�"|s�7V�+����O'P��JdD�xlR����;`� �ץ�!�a�׳lօ�۩�|�<��G���!L{���"An[���eT�R8��[0�I,���)��c��Hw�n)!�zw�s�O](
���Ϋ�ڈ��xG?
��7;�c��oϿ=wI;�l�T�݀%W"JM�f�R��i��n�����a�fv$�Z�cZ�mK���=���� �ێ��[;��n�R�u�N%�l�*0�
�ͪ�6/Q��q�����\��ٙ	zgqs�F��C�q��jp�K��C#-t-��J�U�!j)�F f�\ݦĤ�Pշ)7�kFש��79ͥ��Y���������* i"�J�m�Yӗ�}+1(\A���9) iK�{�����A�ڿ�7���2�h���HZ� �k�T�EN�&E��5�>>mȟ�An"��kcwr�o��[���+�����C�٨AD�|{ "�^^-��^�Ť@���DWB�T�AmCp��mȧ����������J=&��B��	����/KpnĈj�楼�F�y�RA��������\��2.#��� ���(M�^��QbD_D� |F�H�[�%�܉�nVAܷ�t��
���rt�]����������ȶ����tV�N�{=��߾����P��X�Zh69����5�G�%��5����@��c���߯�ߝe��!�^>m�vaG�u�K�E��B��;��z�V�yX܀��hH9�pm��F���R�AZ`��jܝ���>Hug�g��U���p�~��ypޛ�!��(#�����Xv���Nl�41JD�P����G��<<��|��$>����%9����WQ�q�/�H �h�Ds5���龑#�բ9�."ff�9�h�2��uܫ�x�cY'Kvy�ؚH(��|dA9 �VCp!�@��(��U�E��A� ͅ��ۑvbc����GJ�͸�1����	��0r����6�Yw��{`"s �����m�y^�!|�h�3W���U<$\G |���|5��n���&2rq)}W�rr�}6}��-IX����˗2�GQ��q�z_Z3�خ��D��.1{}�^������_�a@-�^�x�O��KS�T�Q<$2�A�z��@�G8�+��@��Am�[bsN�`�FT#��Bnʨ�맵Ң�n!Lq�@Df���Q�0n�݀�F�H�n�	�mz�CQit=}*'0'��'e�;P�.0��1�XP�{V���,���^�J*b����wD���w�^C8%U����y7��� <Tof�8Wzf���Uz"9�ބw�,2��ffhәH��6�60��v3 �^܎���z��Wĸ[}�gbe �xH'�#$V�s�{I�d�z����j�m�!��2Bb�%�/d��UF=�{Q%fm�U�<W���$�2�����>������c��t�
��q����=h�<� �ؒ�`c�W�iO_����2Ϸ��m�Kh/Ol�9·�5<��&w�F���E�L� �-G�nD�� A,��F��^cKrla��A8t��_I�g{�e	�AD�n��F��m�hn�b���9B={�A��x�܌�{*�OX{��)V���Dh��ۘWA<x�3u	-Ǒe�6�C�=xoDE��D��^9��ChOl�E]p��5<��RF՝��ђ�����ޮ���:u�]�N�8>�����uv�J+#�/[�ّ<*nU���)6v4):��RM�E���gb��Pɚ{��V>"���f�-�>n��������噯�fF�p%�%d���&e�A=� �f�"�RA�+��ޕ�v]�ˣ��	%t<tjW�;p�� ��a�gV�6(fj0YV��Ux:��\�^�g9e�eX���>�ou��+���v��!ōّ/�Y ?S�}7�BKp�4.譽����3Y����RA�jǱ����US��{��RA�A��5��Y�;زD��D��۟7��
����3)J+��\���2����@@����mI6�!����ގ᝘����^�h GQ�ۑ6-R��{�
�m˻�p�<Drڙ����������x���� A�>m���3�6���A�
����++F�
�x@�#ݼ�9�]z<�B����Ү8�����'z���x�� ���w��x����_n�{e5���M�uc��|�klc"�f�/�؝M��?%�)����)�?ӄ^2��c�be�g{l�3	p���[�X_8PS<��{�\���3#��y#��-��SW}�����]��d�]�c׫(�=�[�gh3(
ox�0b�:wcԨ�r(�{ޖ�1��A�����m	8 �i�~��;�aL.�rSL��l�ѫ(�t���S]熥�O�������������9;���f��7u�s��w�[�ss},>���Ni�#R<�`C1x���M�iޓ
r�AC�\f�2F՛�
���s+]�׃U�3�u���ơ3Z�(��G�����Ea��*�
����i��A��6&��ؙ�����A��jhkŕN'C ㅲb4L���d\f�2����;v��w@[�x�����	�m�n�5+��74�7O�"F�؆5Z�2	�${���Vo7�H��r�^����5�1k5U��&lK�y�)�,���^4����Լ+�I7Hzv3���� �h�;%�1�V<����у�j��_g��M��&����t�_c�����J�iyN7EX�PT��/��J�F=�n������ElH9[#[C;9U�zKM���b�i:�Dd����ݱS}�Y�9�7�g���b8d��Eڣ8��A���j~^��h��֦�P"��@'�U���u@[ݑ�ʂ����!.��"(��"*F5-�S��=��'W��ݓ�0�w�Տ&#e��\A��Fi�v�h$|A$��~5�lF��;���d�{�:����(��vۋL��dڡ{��ڴ���3{X�%�e���"qOZ�R�m٧'8�'v�N�������""9"8y��`��t��H8u�k'+�9�j̹K����I݄�(��Y(��<�W�H������@�^�H���� ��6e$"(�<ʓ�J$�"jȈM�9�؞�I���q6ӆ������I�[h3�p����МG�bG��}�S�N��mk��;�9��{�>Ճ�XQ揳Q�gd��lw9��8����ν�ݞ���u��6�m��C���))�����8���x��pB>���m��7h��اqə'8�v��n�[�y��o�@OJ��P��ݝ�۳���ރ�����6��p�2GNm�kv�e�������%��������)���n�Y�.��-E�!�y�c��v�v��[��Sn(Ջ���i:R�T'VSXN�mTbz�]����1ôH�:�ћ :K��̴�KF��V�նذ*��l�&m���p��ޥ�X�fT#`��#�PΤ�AGA�р���o;f"z�k�1�!/n�3�\R�^B���7]e+q��m;u[<YV�n�y:�ؼ���ͷc��iS�=�X�۩�(x�4�=���f�8u�@���n�"#�썦�rdj0�.惱���+VZk,]3֚l
Ŷ�$YO[I�8�Y\;�a�-ёzؗ`�T٬Ka�c��ɵ��S��϶�j�u)HG��/b�IZ���F��ۅ��Yֺ��2�D`+Bh@���Z���(����t��ك�SW=���9s	T<�{m.��p�^��=t�6rH���V�� ���Q-\b�3+(�����]R�X�,P�f���QŌ��YT���4 ޞ�7].-�c�`Y�WL�4ͬHj5����U�7L�wW�.�����l#��v�F�qw\8�ε�X�5�Ÿ�i���k��y�,�
Xvذ �b��0(�,7V;g:ek��u��7,Ʀv�v��U3H�ZY�`]�F�	A:8q���:�g��HK6ZU�&�Ɓ�R$`�b4�4\[4��]A`��y�w:�V�r�;L@�Z.�2�EdN���5���I�
z�S�[��Wk��sz��}��؝荷u�7��lڲ4)�\\��h�`��rΛ�5u��$Z�ч�^9���mQW����ԉ(
ڄ�(.݀��ee�q����	�v�ն���K)�88S�v��a�h�(󕇖3`�)�i̯h�A T����q��;GY��1��B[m�6yN��=8�U����k�iٷE5��u3�fZ�8�b��Ǳ�/;P�f.�b��R�c���tu�el�4����t���Ě�.�^��Tq����Q���:]������;�=M��i�DΠ�ZlL\F��b�0�p�(lxg�^_�M]r��o2*F�	-�	������95����ss�9�;{/K٥d(�N���G<1���ԗ��+���z�Kv��5�!}��x/���Fh����%��KضV�}��<�F�ol�&�z^G�&u�!���^�.ڕy�!�n;gF�R�6�3L�폿߼�Y��c��G.�Э��b[IItlXL��i��k4� ��C����:Q�Ȓ�"	e����Wa,��V�2���V膦Nl끾 �Y�r�me� ���C��֜�e��Z�l�-J���ʄ󅺺���x��7�$�\�V۾����e]Tϸ��FnϤ� ᐋƧ���G\8�oxۑ�+���*�����r�3�/�Q��[�@�O����t�f���}���s�WX9յ����3= ��@DY2:-��\pD�� ���P-�$6�2��'���˼��r'+Z��rZ��mU\�p �<W�;�"Kp�%�r��Q컾2����?��4��醌�-&Ċ��Xks+-�/s@ՃejŭX͙�s���cı�˘�-7�1E�xDMO`���)�|�#�)�#O(�mϛ���,��b�R*i>�I��yI39��%�ӌ��<��ypA�9���m�"������(4���K�ò��Pz���?����p����]��}`�o^�ң3 �� ���ᑤ [iVUb;b�mUt���f��r�h]G�mȝ�n���A�\�+s����mUd�w�����B�-Ǒe�m��n,�n**����� o���S�9��/��D���p�n�E���,�օ,�#yȒ� A�e� ۑ �t��t��n���ģl����Tf`=>#H@�ԐCheԫ�WeS�2{+�4 R� �)!��ݎ�4�R�.�<��hmf�hSgY��{����9H ��^!��-��V���޹���VM�Qi6o4��ǨI�	�!���"��W;�=�ꃕ�%��� ������a��Ṇ�Q�\w� ���A7�1����[>ˏY��A�"An�x��uE�l�шL�y곢7�Q3�)��P[�SB�pE#"�ݘQ;,;Je�J1�E�eLTK�>������P��������^2CE��B1�_�=��e_B�����[SFfS��� /��Ԑ[A��C%��ݕ����gia¹}�yx��H�j�l�=j.z���5A�Ј�,�L����� A ��^!�2-�C�[�6֥G2����Av��-F_
�Mu�� A���Ƃ�ǐ��y������[�Ƶ�Jn`CS����u��x5t/B�wl����mL[�^��a���{�=e��Ȓ�y�v�]!��{wT�*{�7g\M�N�$�椂A��͵dS4��ڪ�v��>y^�EفQӽ�
��6��j8��;����n/^�1���'�Ѱ�o\�A �@Dpm�!�.��yn&�rN;#_	�Mm�� K�R>Ƃ͠�CnD���n{d�Ô�eG�ג$��A!��Ӌ����kۺ��S�A;���1Wlt��sʧK;#o�"`E�gM�X�s�{p~�sUu��N�T��Ƨ.�mH歾���;r�jK���:j�n����B����~��Q��˖1�jHn>o�[��񘗆= s��e���p���7�Q���!���Ǭ�ǋ��gݞ�t�Å�i�w:Po*�1ٍr�W7l�MK�6\ݩbW �����C�Ͻs "��q�>!�
��q��N�2k�Ǯ9��X v&��ǆ��^!�"Kp���x��U|_lF�AY����H}���*9��sAL	���l �̀�mk�k*V	(/n�	�� �� ��&܇΢�B�M�V�.]�������G�� Cּ�X� Cnd>ӧ2�Rn W�>/�/�RA�������;�ɮ���Ƿ�����.��:0(��yx�9qǑ�۟7��&nbc��z-�u1����mZ����} #�m� ����'Q���K�ͻ�ޕ�.�à�	�#&p�O���E�oM�~��f̲ds��{4�lW�ʨz1{O�����P�e���\`�E�D_�{��i�O�з$�&�&�&�z�0G�=�9tXu���Z:6�6� �@���4y�f�,f��8w@��.i:,<Nӱ��z}�q�դ
���Hƻ]4��F�5eW�m��7�z��%���&K�mv�r�X�M
Efvګ�I/�ͼ[Dlދ���u�<v��M��zOn��L4�����p�a��څMCE�u�݌fy�$�&����|��]�n����A��dS��0fŁcb�amaH��%����O� ��^^8܉���\d��������GG�����NUHʍ��'6�$7m�`� Z�{5�zˈ���j�A�P�����	�L��1�������};}%�5&7�t�Y�wG�mȒ�yx�� v�"�rI������w�̄AK�sc��'3�3#�'� 0o{�l<��VF\xk�Pmȟ\\E�NwnJ{]l�q� ��z6����Σ��p�m̂[��>-�@��r����gr1��r':�^�1]F=q� A}�H-���C�ʹ7�tUYF��ˡ��10G0]�4.CRhX������=�4ר絻��Xtk�\�1;�bgr�A̫��3+\㋅���>�"�����^��o��������;z̲ٙe��e�J�|$��6�!Ul$�n��!қ5��@Q(�ݷ��ث�:v�$٪�����&�ܘ�OLP}v�wd����;U+%
��&��{�}�^!�H�\Y�99�ۆ�˅Z�=�wB �{"Kp͊�����͋n���[��m�7L��j'u�
w�f���Vя\p@������q������2+��`�X���.}���n't��=���AL3�A�B���p�ɝ�x���^͠��RA���q���#}|�2�D�i�=���aB���c���D�D����7[u:w�kϓ��_~�˿X ��B]v �4�����@�n�TN���4���\�^\K�Og�&�__��-���xԐ�&�5vEgY��0k�Ǯ8/n�V�bgw6��G�myx�܉-� ����1q׽S�#���� �;a	�8���n9�4�*zA/� A6��5�N�mxV�� �� |�^ 6�`�^<�֞\���Rj&�r���3V����w�:��nx�>�=�a�N_{���f ZG�G����ͳ3f��j�60˙�Bf5�=�<�\Y�=݆
W�ej������y����%�|۹0�����܉��q��� [AUn%����d����t����0�M���a��(���[�ŖP6Г��;�ֺU��U��J�����ӷ����0�	�0�[jHn­OVקW�a$�B�PKsԫF�OssٻD����Q������c��~y	K֧�>@2�<[r$\�6��Q���J٘�a؛��J�ц�s�qd�>mؐ|[�� vD甈�y�A�B�q.�W�jܑ�`Y��or�3`]p�&�������"K�@��>M�p� ���W
�7y�\��n��m������ �p �i�-� �A�"6�4Up�#*�- � ��ףʹ$\�/'{D�K�D���>!�Ǘ!q��*��oV�R�j���p,LAyE�ONx�Z�}t��ؔ'9<�R&�n)��Mk��I�
��sۇ�{��=�(�B�tCn|$� �^^/ᙹWT�#�u$U�\�ga��(�Q�q�;���1��ŷ#T�wt�7"ز���H�L#�!j�^�V���)5���s�d�A�MMu&����<���F� �E�WnB�a��%\���3ZtӮ�.�C���KȽk�����%���n򁄷i��u�ip���"�8��bL.��N��=��Ȑ[������Rr�ZL������̩nf^��Ɔ�\+%^ҩvfWM�k�v�]F�N��v�"o,�3*ؙ��C�V��q���c��\� ���s���!]{
�l=ŉ�a3�
�	쀈�sIm-�i2"_�����Ax��Am�Hm�CqQ�A���`��FBعzĨ]-������{�'Ÿ�-���R�֬�f ���U�D�kB���2���Ć��9&�sx��>�+��a�ػ;;�����t�;=�l�V4loݑ�������ӷ��|M+5+��5�q�l햻i�Ӹ��=,sL<�f0H�uZ,k�,4���;v�S��	"�V����غ+tއ��`MF�-�zvײt�x�f1��S���1�d�2�����A0��mk�<Ӷ׮Xc��n �kXC�ܡs�Ѫ�`��Mg���sb�ק�:�1\���/���)�~�~/������m��[s�j��0��W7Fm�����9��ó�K#y{]��\g�d*����Rk'��4��uv���H&�;����Ԑ@m5غ\�v���u�����We��Y�����F8^>!�"Kq�p�����-�P�P~<�q��ة�-��w�c� vFk@6�ozh�L�>S�ݼ����A�x(�&w�;x��N��JKj%.w������6��"&8����ٸ���ʶ�NL>�w�B��ep�޹�f��d%:jj�����w�[�뛡��8�����ެ�w�c��=��m�іfy#r�Q�fm'n���/W$����Ĭ�J$Y�QH�$W��k�a��m��19\����ډ��4V���IFOn��pm�m�`�"�37�[KU�����ݝ^��F�kn�8�q���8,a;qq�J�zr3:��'J�a{/L^��;vs��:$�X�k���e����u���{�]���]G/`ᮣf��y�3����4l��3�����m��﷮���ў���MM��{��	�F{��cM�p�E��ޭ�b�|-�:��ݘ����
as�����BXˬ��V�盁m���8�n���(���T�qr��:2�5�n�����a��k�OL�!�����YOV�R�%f��Bb�:�ci ��`24�%��>�	A��Q�{�tׅ�n�m�Ul����S��p�YOc�T\s��my�m�1��/lS�\�N�;�o �wva8��bf'��S�7�y�6�"#c�C�[�3��y��h�2{	���c��P�~��b�	}F�0ɓO\�:c���������
�>�뫠�����M��x>{�*�w/n�axd(J�b�Ћ�*���N������wP�_s�y�*l�-���lz���R�흢�؛�{5O�Bg�d�䅕���Dc�� �sf%n�n����������e��-�6��yQ
�Ά�n3���Ψ�v�n�X.�^<c���n�{�ܧZ�����3"��2pm��K��^"m���ջ��d��d�w���)��NaT��xo�׮ɽ��V>>er�M[G��@��}�y���a߹�������g��6���Ӻ�2��9�s�_Si�m�g�����,=�'])zJyإ���O�U�C����ᜌ�94m��x�U���D(""��c.��n��!m7Lѻ/4N]KFx������ז_&��5�eA��)?8�\|�|��e�=2/,OZ>[W��
�[nk䄣%ajEV�jn�.�v��3�XSӥ]ࣞ���5�����VS�DΜwB�������-=�O��9}�v����^0?y�K\�v�ｄ_+2h^�����oE:��7��y��^�S/	=;Ǩ���M��xm�b[�^+�;��f�xe[��u��輱�|+^�Ĝ����~��.��hɚ��NH�Y\J:<9�3wC���T=��Ŏ�Z>�R\�����ߔQ FmJqR`]\�Q�vC71�Cw]:íܸ#͍cE����ڡZb�ƍ�.+�Iㇷ�p��=<>j�=weY�d��9ge)��$��%�6�GG6��vq��=�N��2�ٓn�v>��6Ś����Z��hGw���{i�q	��l9A
*Ӧ�'98q�v��.�Z�wDr@�ֵ�X���Y�-�%%���Nr{`�,��drHsk� fw��ݭ۶�۳���B�m�#l��=�s�g�M�l��bd���:�YMbm���Zgm-܅Ig�D���ƚX}�����m�6�rq�jJ]��t_lB^l쓧$��f[v;�l�Ӊ�l�;s����3n�+S�&�{Yz��z^֧{l�ְO,'�yyμ��f�Lm1���J�8��kD����ق�gln���[�Fl��q�5���Y�m5��ݹ";*[w���S���$�I��[J�m`p�;�
i*�i���s��y��:2��7Q��yf�m�6�n
��tL�C�`:��x6�[.۽¥�
Ģ��=*�-�R;�N���A���<۹�6�����V�NGk��y�50�ۼ�u �6�D잓��fa��;���|d�̞8�)���ٷ8�f��v�j��֖EAD�)L�ި�ͻ�nծ��O������w�dGc�޷����h7�m_\\��v_l{{P��ipͻ�*]�J+�� ckͽ�|]#��sw*u!�mᶼ{(`�ǖ������:���a(�sL.w�����M��{79���w���l�uZ�n����7k���q�4��]�v������y���sxFлZ��h3�3�ӻ�-{j�N��p�������t����
Z��HV�L��G���3�^�����MT�(eb��T|�F�귆%���p�1�h6h�b̀s]�x��H�I6{�ۙ-���F�P����n���v���3�Y�%�G��@>����j�̦~�愢y�50�E�"�|��Y�m�A��k�������Jk�T_8u�+Dg)����{�h۷Y��#r E������n�o���q����Ꞧ���'{��*�� ci���m�8X��j��^jm�YI�����)��������Lݫo6�pk;�_��?nΝ���4��=?���-6���A�y��m�"�y�ّ�98V�\?�ɪ��=ª���;ێ��/�loz��r?�Ny���r$��7ҹ��{٥��2PS")LL\��W:�s�`]����2!���i�j�5��1擇��׻ssq�BI��,�i[-����/aƢiwtq�q���ë��78���q��MI��Y���	X����
٣�n����m2V�X69�ڗ�9�e�Մ`#���l̷�����N�s���2.j�u�5Mn���߳�m�ci�on�R��0�.qv)5�i4&�2B8�ƚ�M1��z���h7 6�=`�����jX�q4.bu��I$P�hgr����A��RCu%��MGOz��܅�� ��hJ:�V)��n����d��͙쑻bi���7�y�۰��댗yiTvas*]�w�y �h6�q;�69�l��mm�e�f�mD탼n��R��U���w]:m���m��(�l�t��׏'iB�񄣫eb�]�n�u��x�<n��G��R�`(:j�t��T��F��q���˙��5���9"�4%s[�	'�հ=A�^������vи5.�1��;�m�5$���6�p<�C֘}ɯb��w�3�z+�z�X[R�ˉ�b���憐5y���@�΃s[���Yl��[���6�`��ב��4r�Tj��d�¾�}�/��߁���)�ۉ�]���i�}�������y|����m��3�X5���y�(��X������pm6Ў	�T4T��w��z��ZF�h\˹��{I����A�u���[�6כi���i��#��C]yQ���cwP���&iw\{1�6���3Ц*����$�EL̢x�����s�Pp���4p��X3L�V*�������\ᶀm�wt�{ۚ����a����$�������mx7yn0f|��cjWv �=;q}��WeF��Ի���vg��	�ss�᜻��3�m�7m�*����z����DzQ��J}�/C���7Vi��:��ChʑP3TہP����4jʨ��⵶f�]��~���j��oc~�������UuSS�p3��������\aP�X�5�ww(9�x�ղ��]��ĥr�1ʤ���V@����@7 6�f���0]u7����\5�Q�pu.�>�����m���i1e-� ��������Ѷ�\1�*Fn�EiGi|���^��q\a*<N�nמ�p<�Q;`�8��쪮��jz�0��Y�������6����J:�'F=��jWH>���Qƶe�������y�0����{9���m���Fj����3[8���O*8.��Wx>������qI8ۂj���F�
��m���{:�WQ�5=�o;�b��,�[���sv4�q5�0Ͱ���6za�͍*����T����z���"�ʸ¢�۞r��2�r'r�f+|n�wX>���{��y��mx7�3/����EFfþ�/�qQ������;y��ڢ�>�/���'�wa�Gsl�ʓqf���n���k�z�)
b ���%'�q��Q��!��nv��<�]�p�R��T��o��t^
��w �A�����yYNȭ��T�T�"v���/��T�������ckͳ�\ޓ8K���Skʹ���n�u���7�
ܼ�oj\�.��y��m���j�ԥ�_��z�W�q���U}'��t��w�r�k2��m�kh[i�����Q�:s�D=-n\�郹�_M0�x^���� cm�o�{��(��e'�S3��;�6�V�-���#1D�Tn;F�b�9�x�ZAnQ��i�sE�4�����r�1�mKfO;��K�ӷ������=5F�0�+���;'FC���7*Bu����=[y.7<�z��
f�5
Kc5�5��d.,`�aŗ@�Wa�f�YHƶ��%msc�ѳˎ݊L�Or��5m�}�@2%۩�͜�݁_^q�և��� �&�%�0�[,�6�3t�ʡr1��uݠ�۲Pd��6�)��I��l����"��{�jgL��h�Z������g�D�k/�
��9�I�=�<\�;:�^�fk���6�o1����߿2|�h6л�A�չ�\��K��q��^�|�S�ƃ��m76�*;]Ϸ|�W\X�Z���<)�wu���=��/���̍���=�.�!���m��z֐۝�-�9�L%\/ML��\ckʹ<� �MtR�BWgt|�n���OW-ȩsP�÷�L$��9�V�����^n<�A�an��U��	��˹���n�������m�Νʴ��v�X&ߢ��"�B��a-jX�ʗ[2h�؈q����dL�I(��/�؅�A��m��}���b&�V���;讜؝5+B���3nmx6�k�if�@L��b���>`�WO�
��֌�wb�L�/4�5�',�ݴ+k��bp�G)�;7��.q5P4���9M_�xd0�PǷWH?���+��)sP�wr�PlY�z*M`�ec���W�m��{�~1Uu���.���#���s|;y�ۯ�t0玼HF��>���h�t�&k=f���{�.2���=%M�ӳ��{:<�^���Oc��\��)�������[8�UB�;��M���Y�}=׆;��E�z�V���J�]����k�kL�
���𧁫m���Q�&�D��_/6�ǫ�,v�9�蘾a��z#��s�|���n5��M��2jd���Uu���܏�@TV�}�=�E���S=�1��9�dR$��:�ᵓ�z����6כgp�Y_CW9�6UM_��Կ��r�q_g�Jo��>�x�>���pY"��0�j�3N�֯^��Ƞ^�%����V��C��egD��ym��0����{���my�w�,k���}1���n�z�nuţ�^��a��{���"���'*��כ���m��m�6o&�rĽ^��q���b/�֚��uǱ���Ľ�d�4lA��D"�̈%[��+k�s<��{h�-c)��lW:�v c����!�my�����O�Vٵ�'�89�Ц9�MZޏ6�v�_ODY<�om(xc��c�눱̽�q3�û�{���6�X�����B�A���m�m�3C��[�e�T�J�c�EV������vpkD��}z��,���F� j��v�;�X{f�j����y������~uտ�����޽2��k���ZC���م��in��*Uj�`�.q ����US��o��5_ ��}��A����������bñ_F�\/b��p��y�L��wu�or��y��������АAù��Dh+J�.6-�us�3��(��R�5l�[^��@n����'�����y��
[ev��vLUi�=u�v���*`wk�/�6�m��	[�
}6������]nЬ�hgmR:�'�o!}���.V.�рK����m�������7M�;8�H���Y�|2a��or���k��L�]m&�n���@OM��*;X옪�<+�V*�a�"��;5��A���� ��d��C��ڹ�U��gmR:�Wv�f��m�/���e����������N-��WU[�V��L}�쾋���S����	k��v�����2������ڤ��N���m{6�Y�<Q۫_��vڔ6�+̟8���u��wW����4"vJ�9t��W3��&Ű�n�e�_��w�@��.�:*�=\�A�z| �rP=+�<$o�>R�i?p>����U�J��(2������W���7��8;�uY���Y},v�ن�yp����xn+{��9�_w]����Ԉ݁D�jv"$�#n-lP�&N���\
�rh�'ҋx�q�Fp鬭5EUesDUF�z�
�Ȧ���=a��@��ݘ��M�"0nӪ�/ٺ�;�^��,����y}�Ƣ�\^���o��������Z,^�q�%���2/w����%�f/D^[ǻݴ���E��zv�]��lo7Ψ|oNٞ���݅����N���J�
e���9��<�5�8��С ܜ��Ignj۫O^=�o�/�SL�����Q�x����Ǧw�������"v�kξl=�w�n[���`�Gg�{����1�2u)�;���ol���ͭ�3�c�KO� w>�$5viEu�GŘA��FU��^� �6m��ț:��D"��_�{-{y.��� �p׹j|k*���?V��{5M���B�J.x�aS�ڮ��O��Q&Q�{�!�5yy��ݸS��wvص���WV�x���0��v���E��y�>~����;�B�y���dw7u�ڦ��fx�(�ַ;G��*���x'�+��Yy[pF�TdƠczą YA�^8��m
���R[l����k��]�۲�+kt�8B/l�(�{v�Q�$�tn����Xtr{Zy���Ys��q�p��ĜD!3	'#08.�K9�#���$Sn���' B��A�\�H���=�f�[Q�A�NIϵ��th�f���{��R��h�:�N�ΆEaN�����0�8���.r�s�nӉ"�њ\\�F�[]�t,-'p�҈RNN��Ӣ;,�mZ�m�噵ч!�m)Ѕ"e��鈢ҲfNq�l�m��+l'Q��ɖ��:ma��5�9�k-	:m���ʹ܌�݁g$��-���G��4�ݥ�ͭH�^ݝmX��k���Esv�"v�����!���k��I���.�膍��ˠm/2�T&ׂ3Mn�wg�؜u`�kzy.�.m�E��L֋�����E���]�q�'�kP
kuaͨ)�!�]�ꗷL��lm��Ǫ���n�S8xȨ��S�����8�F��"���	Ms����M%��.��a).%�y �RW[�%o�0�z����g������v���%����$`�Q�\k�ӫPZ���}�]x�s�ƫ/4�.����ۓ`����s�IaE�F�Fi�A�������䔮]�<���� �У-�M6�Ћ�*�R��vMط:^��c��M���'a�h�A���v�<79���
�vׇ���*Gqu�;G������n3U�:�=���[��ƅ��zѝ�sy�!���׬���b��Ě6bJh�^�eqQ�k�)^]bOch#��㫭��{k�W6b	�ڹs��������\���.��N�1i���������u��ici!4áMQMc
MBb \M.P��P�..���<\Ƅ܇wQ���P��I�ٟWj�wm�V^�lu��e�Ƹ�!�.�(�7n�n�k��stVB�朝<�1l���� ��M�c�Y���Q�� ��b6^:�W	�N9�mm6��V��Cq&�����7^�-[v/7&�c�j��h��g��	J =^�qkp�0Ѣl6�9�َ�mWi76�z�1�N;	ں�R7iظ`�n�n�ڧ�}�󣍸sgr���5�����[miF�����[g��ZQ ��g���Vn5{���8.�����O1!ѳWJ�Z`�CK(j�p�0ZD�t�1�Jłj���»g=��zWx��'�@g���'&�N�gm��k �L��`��Ocp�t��ځ��n��e��f��2"X��u� ���+�T&�{LKs��A%-ݩ]+^�r��]���&p�a⎅e�O1��T�:�9���01&�)����� ���0竣��|ex�tq��vD��t"���ֶ �M������^k[���>5��vƸX�s�G=��*tp3���Qa�ĳD5ұ0B�
��ҙ�ҐpZ[m�[�vQwð�7K]�D��۲��'XMs�e؞"/c�!�j�
��[��{k{	���8^o]��v�q�ܴ�0�5������/��Qt���r]ظ\7V�ĵ�ܣ�Dn3X�vi. C7[�o��� 7�͵���v�X��s�̾0���A��Q��]����A��myh0��N�Bۀ35���J��;&&�"g�]����*j��9��q�վ@6ۯ6����jb�ҝ�5��3v�S+���;5�<i���j�uo�^{ɸ�������YR�dû����P�����S��s��n��@6��17�m����^WP���pvT�����6�m��{�anaͭP1O�""$2��p�B�+k�����a,�FX�����v�o�}?������6��mM�s�/��9�ԝS+j��2"���-7ʹ�^�q�S���FiU�}�.{�I��	��+{�-�k,h��7}���%�>^^b,y�_{B��[Q��D$gcW"�|�S��	�1c�ל-K�\�{���m��4f8�u�3��B�=���m���D�Q��¶9,[��R��3ޞ��my��n m�*´���WsC�7��`M�k�=��9�ԝS+w{��㲜W_M�Ϯ���my���n�t�}3�K���xN����Y.xor`y��m���pyD�<R�>�`�+RsHKp"tn�`b���w7Nd�;tk�B$�4�u��+u'�z���~���꺅�#�F��T�lL����v��
�f��m���}C^�{p�*i����w\�Onl{u'T����vj�Z%X�L�����m6��E���2��{j���Ze�9�{Y����ĩ�OC�u2���Z�v���T�UԞ�V5(�ynG��$I�%��G&D�uV��s�;�K��n%�X�\�ܽ�m����6)�y�Y�#i�k�6׺�v�ֶ;*[=�uG����ßdS�%<���{:<�A��nwt9�La�� r�u3:ہ�n�aJ��w/vj�q�ں�絚�f�����bfdD�Ny������k��^��<�ݑmq��h� Z�8!�xV@��m���W����e�X�\��x�k���6P���^�m�m���ΪgUo�e�Tc�]�yW-]IV����כn�u�(c}���/57m��ۊ�'&+c.����^��=��{�Pn m��K��1�5廸����K�{�+��w=��ܐoI�qݢ.wEj2-�H�7[p�^бb؅�f���e�"�N��;?M��Y�f�ޙ�Ng��F�M$^V_E�g���@�5Z���q��m���U\��\�&��W���:���J�����^m�����q��O�
��*#���M,��6ζx����.ՀϷg��ĉe0W���X�{\6�nn疛�l�{y;*H��|v����ǭ��~n��ڕj2��8���\�ޓ�'8,k.xy�/k�����̬��Q��[q��^m��6��{i=�P�]��e�ۊ54�\T���Ͷ��w*��<&j�@����黨݌��^�Vʕ=��
�Y��ayk}�����۽b�̞�\ʁ�Qy1�FhY�cYs�ϹfǛh6�7��֨NL]��Ԃw�&�[(
Q��zz8EDƍ�F�o�p���n��S�<���W�Gw�zDUu���U祢4��Ue�f H@ϒ��I�cwrv��V�\hɮ�����QZ�]a�3�`n�gF础���I�����\%����28n������f��97'g��o��{tp�-��r�ź��]����s�Μ�1�s[(�ΧL-K�A��a9��a�9r�²������WPn˓��hL:��4�IWK�'1���6��CK�4�ұ�dCL������Z~�E-��2��֐���F�ԫ��Y�)�.�=r���s�<���͵�t�#�g��Ъ�e.ˍWz���x]j��^n<�^�U�%�8�+s8؛�o)�������T��w/{�W�s��*�l�r��5���^n�F�����W;y��9c#C��\�C�ᶼ�@7]\.���}=����<hm���3=�n⪩��u���B��t5���� �@7m�f����spbTӨ͌��8����*x�^�Pn<�s.� $,�z��)W�c�����7gDh�c�R�@�[H�
6�Y2ں[>�7� ���M��vI��w�:3"�w�t7t��gF/{�sh6�n m�F{cpj��Ԯ�)F�Q'=]�oVT��ԉ#Q9��:��"��(U�ݐw��cV7*e���Q������&3Zl�y��hu����/����R�����fPwg5��z�*Z� ���mڱ��\����g���Z�'����ۨ7��o^���RLg����ۉ��#��O{ȹ]���Gx뉩�Y����m�G=�ƍzV�������Jۈs��SF�����P-�ݷ��CiI��������5,X4u��3���i�K�ѫl4`[	(�z�J�"}?L}���j>���m�ut�c+�g���Z�'��Sy�y�o��k�<�A���xj��7��V�]�[z�Ή���G-����r�Ϲpw�)=+)�d�xfj�m��;�g��]�W���&���\h�{1UGc.��A��(x��@�(�i�%����vy?R�#��L�^�.���W�ɼʿ7�7�a��ףD��������4jj�K���@6�nn�k`�`n��͆� �WWK�2�Y�������wr��]Q��9;�o�v:� �i����6�v`�貵n%o���kB;]kx��qr�w��<�^�nHQ�k��tS7��D�*eL��L�ebη=<�m��
]=��֓�/2&�T�(�*�W���M��J�1ӛ}SFf���V\�߮"ynPoS�A�����ޓ���̑^\���.��e�:q��Eh��5������L����6�m���)����^n+��_?bZ,�Y���ti��M�wI�7���O��mW��c���U4�J����Ac�
f�0�k=!*��:�yoa7�.n�u�{tf�-��b��>�Ytz��^�A>�w���٘����UP�M7����A�m��^�*ɝ���*�gk<^���1<=��v����Y1����ĩ�������B�[�@�e��-a�r\kK��"�N���{w[v������{�.m.tł���T�מ6�u�:�GA��p;��i�]�:__UE	�b+��[m��g(I��	�əȨ�U���� �M��;zic��2'c�*�g\m����ܽ�Sp<�m�uf&Z{��V��C3W��
������tF.m,{�fr+�Vf���y��m7r�*���(c,�.�/�r�����T[h6�m��s��·�άU��NKQ5�1�R�j�q���w�n&�ˊ�f�"'���SN�@T`��<�*-���
�H�jLA�7�#nl�@�	����RXPZ�z}�����n�F���)s��9J6�G�V��	cv�������
��-J؊���+����:��q��Bvk��3]�3��lЙ�«e�m{Y0A	���֍��G;c�u�u�èP �.GB�f���<���*0I^���u���usuL(��h�6ȴ�uX��	ƈY����ikGB51[4\;��)������1���Y�Wd��٣��j�儺M��[���tұ�ZP��*���{�ᶀm�U��m,�g�h��*q�[j�P���o,p<�M���[yx�Tf�7����;у��[��Z�F��������5�їζ�(z�m��y�W[�����]F7���K���Q፶���m�XQ8^Z��&�iw�%��=��Uw1�����4\�*����)��<�.�=�[w��ͷ�h7۶btT��q��U:������}�{�6כz��l�|"	&(	�(D�4��Ѹ��0$]M�Ֆ�x2uM��;]t�S������Ϻ۠�^�K��n�Lpb�И��0�1S�Gos7W���m�b��Ú�s�-{��zp��t��\7���
�$��I��!���i��{��բN���&�k����W�n��b�b���B����B��t��y�76ʅ�or{�7�:OT߶�t�Wk:m��wFN���F0���T��n�
6��\�u��MǳeEI��l9��^���m��t�dN��0pH��8 �BO"�U�T�;Z�8�h7 6�:�|�'��K��ce�J��P�or��gU��Ī��Ăk�"�)T wd6p6�qOk�n�'8��.��d!B��>��D���͵��zk�0q�U�8�_
9+��Y8T��}٣/6�ǃm0u��+�Q��3�R]p;�m٥�qn��M�*��{�1�۲F�l��}]���6ۯ6ϟG11H9RU#��Z:bnαQf��]�ɹ�#b�N&�\Tݝoe��>���_l{8�Do��F��3}GvͷV�����Z��;ӱ:4����ܨ����K�ޛ7�L۾Y����!����������� �{f�U����y1�;�6C�^��C���������+�7��͞��Ւ!�U�pL;������Dy�D��8�)� -ݺ>����~�n���S�|4�Z�S龓����j�i����/&fclu Q�]�H�9��3�z��{�Pt׸�k�������5�0b��.[�z��8�H79s@=XH躒����uy�~��8���n����md*�����Y��H��}��;Q�@;<|�S��1p
ww>��CSzxe3vD�^��d\ޫ]G	���h�Lv=(y��.7��lݙ�#���z�ׂ��g����I�q��Ԃ8��ԝ�<S����ߏ�d�ټ���O����1���ٷ�n����,��f��z��7�詓AF��,�q3�(���4a���;��UOY�ܢ��_n��g���&M�{�}�7ܞ�D��gKВ�0�0>�×���pL����W�zMf��\1:��D�	�A拰Bq�6�)�M֌Y��v���7�B7z�ޝ��) �����+�x#7�����:{W�u�C�=W�j��5�Y�7�{�5n���Y�&�����J�}���Bx1J��m7�;��h;���}Ϸ�k'�4,��i��
ͷeo�^�K[Z�GY�q�n�N����g~=��3��}�|���;0�����&�$$����VYם�ÑB9J^ۣ��of_k��`r"�m���w��Ay��(�m����s�p|�y6�gMh��[�.�"C�p>���9��γ��ϖu$�DE���q��D^^��.�;���e��w��$����)��������r���#�}�=$[nv�+��D��!K�ѶQ)�������L/=2��y��i{_{Hv"HX��)-��W�$�{ס�g���y����ܳ�d�$�+r}�S�R�q#·y�h��9�� G������fח�N�^su�����i)Di*))�[B��o�����8֖M�P�orwSpm6��5�"�<W=;]ޥ���ǧ��3[���Q��÷�2�_dh�r��cM�my����7�Cv���Ipź{YQTc�tm��8��aÕ!^�#		�㶃�K7g�&ݳ$X5ڤ�v��@$�7oe���7�T��~��t �@6ת���C��i9�*�hF����<�~�m���m���'oT�.X�n��X�<L�`ޅ.�%w�o 9�l�:$,�/������n�z��tM�P�n��AUTc����cmߛ��C"\R�=<n���skʹ]Zޡ���i9�*��*��l�Awa������95��������z�5�{�H��ML`���<urn�C�G�Ȧ���T˫��h����m�n<kͱt���|2�+�g�3Tƞ]�2Wv�����Լꖆ��=b�ܺ�W��LJ��	)���N��E�FeKۘ�M�ym�:�]��0�|����ɸ��]�K��i�7M
��2��\�t��A�m��CeBS3�7�����B������������^}��"���\�^'���m�(d�ё�7�1[�܁��dj�6k&8y�/s��m�n ��4��.nN���{m�\]f;Mp��DЪ�w@����G�����C��͵�����)����I��zD�����.��/��y�1��!;�
[���J���p�Z�6�L-5IO�����f7�G>x�o����-�p#���Ǽ��A�2������OtE�n��d1�].�й�@�5��MM��f��Z��.�y�m���ܦ1:!�n�C�7mr�Z�8ɣ����e�A��q��0���4ێ�2K���;�x��ή�����5���r[EoN:�n�fOg;�q����R!�L��=���v�ՙ�y�b�q����X:<�>��po���!ڮr6���5��1��~�_�Z8*�����(=��/��q"o=T���J��e(*a&��t����q[]��N�.�f��sfv6�k�﫮@��i��pkԘ��ɢ�f�w�����.���\��hUpޏf6�E��w&�=P.�{sSpk����Wݷ����������.� �Pn=��m��N@U�M�o�M��`�2k7 �pӘ�>��4![ƫm�8�WK@vku���m��`.�Y»N�D�f;�m��LЪ�7�^6�����j����9ߎWl�7	]��7E��Bn�e�[u����d�%"b`L([�\6��*��ޡ�C�k*�.��pk�/w���/u׃m��n��9HsѷlI�Q���i�q��a����/m�m���ez��Q��O�[��V�hl7�?~�d���ʘ7�݊�Eܘ�X�کFr���o/f��N�UN�H�s��[�۽�P�b�}w�]G�k_čݑ>;��wd|�m�j�:�{�D%�b�Uh���p7	�ЁȒ7v}>#u{wU�5}�#�>��?�vjL]�W��wU�_}C�>�YUp�)����! M��b(\h�ч2s�F�̂wa�vD���4,[t~�b؊����A|�xh���v��/߽��~��}�Ќ�ns���A�y{5��7�� �� �4� ��Ấ��і��t؋	\s�c.�]��Pq1��=��~�� �l�;��A��=W��f7�5�������$w�wmߘ�P/:*=�WHݓ㺂wP����&�mX���Z'_*�������ZYUp�)�w�@OwH���u_BU����fH�3�dwa��Ȓ7vg�u�&�ꑴ8����[��n!��D�e�{Tѯ��dD��g9� H��Ӳyx�
�G�c>�i��$L{�p^��7%�݃O�4{E���B�}���M��O'%�j�*�vI���_��� �܂;�����H݁�"���y���Ć E|Аw�F�ț��Z��߄��~����{�D-�����`�������� ��g���wT�n�����~P>ى�ۜ0���,�D_�P��ZYUp�
~��wH�wc�ۻ ��f�����[(_�;����������IC`k���jm.l�2]աuV॒�t,��Ǟv�_=��-�"A����u�|~��j�������s裂'~���nb��+��|F�@��@C���3Yz~����:<����ů���������^ޏ|3vD�������G}~V�9ڧ�|� n����$�S_}����Do�C^�W%�7��	��	 ���$�@��@n�	$�n����켑$7�'۰��>?U5}��W�R�A�RDo�鍜_����S�����<���+�G���F)�F������X7�J����k;]�eN���^Y.?a�����`���Oϔ����,}��$����QQ����� 9�ވ����M|>��������q|�'9�j!�Y�]<W������R.[)t�mRKfp;&h&�af^i0�hYP���L�33��H��%����H�ۺ��㻪E^D~�֝�M|�d�_? ���=ŋۋW�>@?�g�lXݐ7w �n�#e�]��]�����H!��'�}�/]}���7}��W�R�Ǿ�I��/�K0s_m�u�����D(�7*H΀���$��ݑ>;��n�_flW}_H����-_�	��S�7H ��y �dI�"|F��R����у]�*���V'wT��">���|��J�m/���'{�$�����/�)����yǐǲ$��$��7vD���s7
I5=>�W��<����5pG���e|�{�GwT�n�=0 ���g�+T�ɚ�d�Sp�}�z�U��~_ޜx�:�W9�RZ�	ӽ�*v�z��6_N=�m��6��������0����ci�?����h�Jh$���t�Lv�<h9�4�n��:`68��X�á�O�R�g3%�K2K!��ɮ�h k���B�����uq��Ĳ�m�4�,�Yr�s��� vN�}N�zí	�׊��1��z�m۷3��in����6X�A{t]�u�9�!�q�ƥӴ�W;1�:g�W4%�c��񮫄ax0%��v.��ffs]o�6��z�|�߻�MtL��8@��j8Е��X6k�����Ʀ�Isf�c������Y}f� ���$�@wvE���õ�߅��Ww􉡟}����7`#����O��Ax�R'wT�Y�u1usg0da�,�� �ڪ�>_N6�S��W���>;�! �|��ؗR��p�hp��4hG���9�Bs�Ѩ�9c}���8?UK�L۫F�ς:���̯���RA�A�^�wuI������6��(����vt� �B �wdM���=���Z������Ё_}�5[QmF}���>>ߐ@��'wW�n����_i���k&Lh������﹥��k�.>W��pS��|��}ϤI݄wd}5ü�����|�����Ԙ�Y��b@3ʷM�e7h�Z�`:�aY�Kp�2]�'�����e���i �ݙ��*�ώ}W�9���2�����Q�����紸�+PGwT��wuI� |wu��a��ڶR.�e���7�\M��}���L�th�)S�%�@�๬�E7�M����qUm����\C�DDge�<����Ј?}��b����ڙ�����Ёu	#wF��F:z�P@�r���Ӻ� �����K띈�х)ȱs]�W5�7.9^+��S�@���A��$�ǐ���2��*���Qܡ�vH�G}�>݀����\�j�����A��I�����::����?9�) ���7W��u	ݑ'v��tP��x�[���Z��5h|~� �ݑ$n�ψ�A�8>��7�����QS	(�bg�a+3	5[��;��n�ŭ`ꄞ�ك��x�%��������j���� �wT�|��c��\|���)�!���=��,(ԥ �1�"hH!����ue�#�*�X�.�}>!�U��zɞ�,����9_Ow��܂wU���S�li��Hw��@N�Ϸcۺ���X��^��3V�5��mц2���Sa^��Ы�.�'f0Wޱ������z6|�>�,�[�ƕ'}*���C��@���։�e�Q���}�y�hМ�.k���s��F�uˆ�����>^���}�H'wT�sI��W�N>�˘����{�BA���J����7w�v ��#w~���l����7'l�w��O����{�^����VA��Ԣ�����?��v~��R��P��CBk�g��)�ܹ�&��5t)����Cq1��{�������}�wa��M��%��.>e�(����E����f��Dݡ ��^���;����>m����s2.{w���]��ϔ��i5�j����9s�����<�D��H�M��0��r'�����	�F������#�_�e�ϵTnK�1�0i|�W����ܽ��� ��R�A
��J4�\͇����#w��{��wd_�c�]�\|;.)Ep5H ��"'��Mv��\e�1S*�Y_\!:&��^��C��,^1���y9�y��:]W������J7��⨛fj�D]�12�b#����Nfώ�����H;� wulh�]�s�cN��֜��W�N>�˘������	�>� �� �ݑ���f>^Bʱ*�`%A�
%<^�b�Ju�d�<mV%7F�w�`:���g������ǐo�F�n��U_��O�gza����_�6[K����ݛ\F�w�"9˜��9�Xx�~���l�n�}�}�>�k~�����W������/|�dH#wk����|�@�b�AתH;�ۺ������_|���1;�s�1<&~����'�vn쁻�$*��I.��}��r����j�>����L��6"�Υ}�	�RGu|"�+�@� >ߖx�Խ��H �ݑ>;��it�9��d��W�G�qw_�?}�ޫ���h�s���g9f�ޖ��*���Qb6334�=m,�#$�	5����ԛ����E'�EY�B�3WqQ��:[�� ��Σ�!IV�Y��	{�@��M��}F�Ɠ�r���y����e��0\�Yv�=���d�Tƥ��kQ�����n��wr��<w}�3I�vv������Z3T����_a��^"�o�Xq㽱�)��o`w��/j=�/x��yo`��+rK��?f�/(C]�$M&/�`��,��y>��z˹�s��s`l��$Ǉ��p�R��<�q�pV��R����.\]��kO=�Wއ��e�r�PB�[@��+��=]�g)�9��R]f�w����4�OO��C*K�N�˻�kC'�ɮ���.��5{�gOp�K�m�l���e^���xH�F�.�VDDcSL;��q����$�܅�묺3Z���u�I3�T���|�"���79=�L�4��<'3�{�O� t<}�(֤FR�Ǥ�"of��ǯ�W{Nu��m�sb�$nl���ňɞwV�=���92O��k�&8� #۾�N�Ep��d�yu�7x�;l��N�C��F�tj�Pf3{WXfx⟳�^bL�*Vњ�Xo�e�D����/o92��ٳ�H^�Z����r�D�L������禚Pl���{ޙ��w�*�#�l
 �[�3v�3���^ކ�x�������j���}��y5n�0��^�Ol�\=��?u�[UI�z�p�w����,��������ڤs�ܧwl�UQ�U�[h��B��8�'|������Y�t�;�{v��-ҝ9m�q\��ڛ�Idbm[��y�G ��y�:3D�mi7���Lܗ����l����L���{np��i�������{�ϽbAfJr��б�y�w�e�����Om����6��gy��ǖ���������5��}2Z���J��X[-@^ZK%��B��� �k��k�ͷ#�+���s�BN:�^���[n����L�寗�=�<ז��֢�n��޵��m�jJ�@�%��^e�[ L2�m�Ck޷��#-�jɵ�`�����O1!�I�i�K#IkKQH��u�'3�kr�g|k-��.;t%�����g{����"��1D��׽�7�^��D�u6ӣ;/+{v����������q	��۟���S�=`�DJ<.3ޚaE\�v��&k��@t�l!k��FZY`�	�m5�3��Rֵ�`(�͛NV����k�ݖ�8�f�C�E\v�s%��<��uwc���t�nR�]b�	�E�YlT����r��w.�S]�Kہ��z۾��c�I�;nէ��n���^�It򖛙�,`:62k[���7�P��pciu��C�j���:u��L�u�k[4-� ��uPW�c�,��.��aɉ�V�
���9�\��L�敬�y4b��[IW�n�קnt��L�Z������\k��Yq�:ڽk��:^0	�mj;(�q =��;[�m�..74����qҙ����r9'�� q�ee2�:��t�"�7&�OZܦ�69m�nppm\�#��K*�K/k�A%�A�vU0�����-�[�R�L����cs,�kb��Jb�K�M�	�ܐ������b�j�]�ݶ�k��õ^�5�v�s*pJ�A�YWXivz���d��������PvP��!���l�>"��-�uk��@�q�-��ۉ�fh&�\�e�Ev�5�3��e3���IF�a�6 �ݻl�l</(�\��H��^ޞ����/^8X�;���7i�:��cb5�+-��ňT���mu����x�c�w��3��ѫ�$n�u�����l�h��l��/W8z�r/���u��\��8TE����l�y���]��Z�4.��Ғ(c�*F0�3F/d�0��Uj�ݭ��kݍ��z�ݚ���n^�9��+	��*�.���V:^�:4����Gl
.�Xݝ��.l�6�D���r\N���p��WZfQ���a��%����JL�#�v���e
��e*�z�.X-����ćm��3����Jl��m����#�6�GM���{uF$�P6�rj��X��M0��Ē�䍭��q�5Z���NK��\I�ok�l�&4k��b��fi����w:���i�6�����A&��5:�`)K��Ys�+4����M��+s��*�ͱ*ؒh�UڪѮN�ێ�h	�#O&����5�2�l�T�e��"�\�+��,�L�nͻgTz�WcW����.�C^��n�E��;�D6����v�㍵�6��#ku.��\ߟ|���G0!l����sחZ�\mq��◲��ic�KY�����^�����:�v� ���wT�	��>�朧�W�O�sYF~? ����;���QYB�}�O�ϐg� 7vD�7u	v9�"���埖ε�H����SW�Jϯo�fOױ�u+�Ow�A�wu}w!
��ծ꿳j>ƭ�_��!$ݑ �ǐ��S/�3��wM��m.ˋQ_W��_z�#3�ѡ9�h5�Y`�D�5�s�w\��/P@��O�'wT����s�_M���T|)| �KP����A��$��BN� F�>#wFjG{�l�����]�o~�V}{L̟�b1|�W���$��� �wT����쫩�* �311*"f$�A��-�ի8����\˲�%4.�1s����e�� ;�C� A��ȿ���8�ﭥ�qj+���E�G�NǠ\��n�D��g�㺂wT��wT�S�� %Uw#�M��"1�	����D��".����1�/rv���C��;�(����]�xK��{�0o�����y۬O��'�� AǪj�����?M����Q�R��w�@O���$���wՙ_dE�[R'�}�/w�~ �쁻�>#u��G�p��闗��fN����R���)w �� ���|F�}]reH����ڄ��<��ț�}��}���ˋQ_W�@?}�;��s�o쎔�����D�� ���H;�/�Q�#a������ӈ�OO�F�jjs�z^|lV]G�Ty�!� ��'vۻ#t_�K���)��HR]��®�ҕ!1��B�A��qj����.i.�R��d��o���H�����7}���r��ɯ��?:��3���ٱ�������wV��'wP�6�M]8<����D=�$_a��Z���_eŨ����A?}x���@�ؼ�b~�+�a�s�ݠ���$��Ӻ��;���wu;[���1�D��w����r�Mj����f]��Nb'ꊞ*����eβ$S;/t�ӎ�mn����ap�{7� �^a�e�KX����6��]G�W�@��|���;�D��^ �wdO���&&#0�S�wEx�Ꮴݞ��&ﾙ�_Ԧj>�y�_=�)L|e��r�핫+�]�A�ܤ���-�^ ��O�q�C��	�������f�ۖ����.-E��Y�ޫM򋉙��L�+���/���w�����َ��-=��H8��Ɯ]�5]>,�y�j]��QM�jŮz�_w��}�\s!�mM�|S��mg�_D,�����CD��=���q��`�_��Ax���qdj�B���t�Ϗ�PWW��~������?D��>��zwPE�p����ڷ״��cH�ۑ �M������]Bfi}�r��_��� ��Ј#5�k����qDGM�ȼ<�'��� �u{z=E��]����W�.��+�� Gn娉�����W�0_W�&�v��=�#{�.�7��O��'Y�ݾj�z����O�W���qt�8A�25i�9(o����ݑ��g�ˉ��ЎeZ!�e���er�y�h���"�����ܿ�)�����Ly���rˎeX"f_���{�o߼}P�L����B����
L��
�b��0[tlD�>)AQ0&<tC��5��|�X ��B�h����}g�n�����	�0{:0��2ߐ@����m[�"�"�u-q���Q1?4�o��/K�����s?=�ϝ|ae�|%|��"��%�z�}�h��W��ݖ	���C���f4���[�o3��>7�^)�ܽ����\���xDs޹�rˎeZ#�����;�g����O��?�Fo�$�n�
�k��}F>yw3𬯄�~�=��J�Y�wG��}�n(�ڟ[A���bD?�J�8�T��\ν9���2��+�ﾀ�ȟ��k"�q+9��g���#�b�s12o����N��˄*��9���w����B�5�/{�̈o]�䞾9���0d�t`Df��$�Ј�,Ix���L.� ��Z0y���Ktf
�ib��df�����eŉ	e�i�QUH��֩�2�:Z���+�t���ó��䡛S�}��n�s[ku�n�n�J� �zۉӻ���>m��2��]d�`��E�>��;�)J:N�Fz{n�c�l٣��Ag��8�Jf�ܵZ�X}V�Ti�q.��h�Sk������CF�P���<�c���vC<�.ƃ���"@p[!H�O��	ۄA�6�	�p���R�ܿ�)�ɍ��T|D]�q���a��������ڟ�@������R���h�x�G�悡C�_}�w£��˹��V!�z�#�Yq32���ߵ��Yq��+/7n>m��~��-"~S?�9�3�)fTp��� �� �vD�[�A�h"r$uۅ��eҏ.h F��O���U��/��_D��Lm����9������}9��xw78qޏ �5 ���[r$�.�\
cw��+;���fV�}�x��~�>�\M�L���L�5���?���?�^͟���R�H�'X�M����:�W1å�@���f�_[׭5���Yo���F~��[�ڛ��d��љ��Y�
_2�����Ҡ��}|�ۙ� ���#~�J>�jۧ��=�u�>�^~Hpw�g�o`3�J��Å�7�kڽI�sF����X����K�Ƌӂ.M��g�{!:��7�K��|����_t������V#g���>�In�70X�W���~Uj�|�%� �r$� Cp%O�s��E�A�_F�F722�g�U�	�� A� CnD���^-�!��uv����ug����/�S�Oۣ+��Y�
_ @=��v}V�?;�m�ve\Fo�X!�2	n��������⍱{�P0:o�u��_��Em��G� ��)#v��Am����B���˗^�AIH����T
E���z�۷��nM+($&-�l`v�&J�GF/n@D� ���*�~�}}Q^FU��*��#����ȧ�s��#�Gl�;\�|Ch [���mO��_nv/��W�/��?G�9�+�_O͌����fLp��@��� �wg���ٙ6lV���"A�D�ۑ>>m��2p:_?}����'����5s]JD�2�4�7�	��l���!������H�g�vd0d�.q�b�WB��Y�&�������s 
:^������l��J6��Q���) ����|[jHnͭ�o�Gѳ�0}�9}nU���ԣ��ʺ��e� ���FI�m��᠇N@�f�E��-�$��q��ݳW��,~m,��W�ۣ*���dd|*`}���^Ȓ�/�
��\e7N&#v�v�&��@N��i��0���J�����
�HvL�|����Y}�g��d��3��[��S�v;�NvU.���E�ѻ�)�n�nǨڒH[����/k�.�����w�O	9��>AU��~_T�}�*�~��A��Df��Cnj�=߯��Oe���n���B&e��T��G��j�ު?A�;�.�hY
����@D{"An��܉�������@�ݑ>-����uK�Z{�NvjWʣ�N}��0ws:&e��UD�2�?�D��g�3?\��z�dE�Ъ!�"��^��Gj%f��D�QS���fs���iba.tGgFD'Y�w�ع��x��ʱ��/Bf\��e�����m�W����}��ː^��tVn�}S����Mg�A?}���!��-�O`I��~{ߧ��1�3]����5դ؎]&�*u�rݴ�W 2JcQ�f��������/���t �A� A-�7}���EU�D�N2>?-�Y�a_Jރ���$
ܟw�~ ���܉�p�N�!敚���
}�"|@z���n�O��}�j�}5����,�)}�b�2g��ϗ�v���ۑ>-��ڙ��?���{�7�3W�]��&����"j�^��E�@p�~�F�z�܂<�KmM��}OMU�D�N2>? �?}�1�2u?X�cA��'���A�D7 6Ȋ��I��4z>��G�!_f|�T�=�s;SM@ܾ���|[j���m^ֿ�w�X�>[��c������s_]6�+�n�n���mrGdn`�s��ȫ�[�of�M�t�|r����w���o�w���.˶��Dh��kW�m�ao+��̪f���`k^�u�j#�v�^��H��P�Q�X�٥6V{s#u�6�mڵȼ�z��5�5�,����.��x2��I<c]Z�1�[��s��[�����|��lƄ�#v2(魹8�����f�%3�K@2"�Su�d��WO7C�����tK�&�\,�mk���� )��RZ��)��B�@ln͆��"0F�g�4B$ę1��# Ml6��%���h*4W}���f��\�&���{�
�A�"/:}>>m[�A-� &~4b���s�dq�57gE��=5W��8��\�'� A�"Kp]�k����:��k�$�q�����h�y<�fD�5=�U7'>3�;SUG��Ͼ^���n>m�!��R�@��w�p��!��C���G�Q���Z��Mg�	���P�W}Qjm/�d}_/g�,�6ԀA��n>��Ý��r�H�ؿ�^���&~g#�s�@��ݑ>-Ǔh@�t�3��ĕ�Q	�/H����i��-�/i��h��]4��t-�Jp�_�.}V#���x�����WQ�5�ʎ����v�R�>Ӹ���p� �ڒ^@��D��ܪ]W��8e�D2b0�Kܜ���V³�ў�s��>������I�7�����T��mO.��hY.(n�����4�<>�n�B���}���m\�Ϥ������_^=�.Y�[��Rq�wZ�h/�"�m���ځpM�7�b�s9�� ��wdH���h Cn}#�4g������ Gs^��U]�n�����6�v�>��|s�:w�.XM[��i�r�H�m� ��Y�����R��'%b�����u�s�U���b&e�����̣f{s~{�u�s-`K75p�����(D)�v^ݹ��1QP�P���&�T�}�/7%������kbo�"�g#�s��{�f�V�~�`��������3(�L�ѡ�eX�pX�?V�������>��_qyQ_Wѿu;SU@9��|C��qyN�f��ƽ���@������������Y�?�,���֋���=W]�!�o���-ك/���>�[�d�~���Q�?{6y���U.��x6oG�_�;�ưlmC4ƹ�Prr�lF�4��5ӓ�����G����}ӹ����߷a͘��A��������Q���{�m����X�cł�\f���V�[k�;�����Q��<��͝�#i�'8h��Z��c8k)f7u^=��Ua�c6E�[8�27=[q���˥n��9o�E3`Y��>�����pР�Ǔ��/��}N7����i}$�{���۾�>����v3�C6���'��7����`g��Д䉄Tc�{ue^,�ؽ���{����mta�!�MM��J����8_-��{!�_Vx��Nz�[�X�o&-���㻼#�w�A��V��/VԠ��M3�C�7f�jbUl��2kiC�r5TN����mN�<�Ѭ��bC$Q���N*ݫ!{4������K���+ꨇrΡ�M��w��7j�}�F4���v�Or��q��(MR��
o0��U���������g�'�,�-�$,�}���7/�#�1��|��قѷ��Q&nm��k�]9>:�H4����lȈ�.�l�W&^$_���'�^F���]�/a�~T�Jl����צ3�����tL�x�֎�=�kz�����s� �	�GXy"�WtHDt�������X��*�{�/[��m{�.�}�����I����1?}�W;��I��s_�L�wW���+a�}Onq�Ҝ�{��M��t���f,Q�Y�%g�x�u�W���9�<�G�N���n�B\f�=//<��n�G�l�)I瞯��3��e{5�{ݨ���+h��v�4Iŕ�ާG�&�um�=��"Z������n�m���y�my��N�!�z������,���G<��	�KnӸ��j��ä��u�O���ã��y���6��7'Ͻ�Ok8��C�"Dr���������gv��|�:���GG=�����F�����ݝ|�:m�_m���$�>X���{ɶ��
�[w�h�ٺ �kޚ��I3emx�����y�ҽ:Ӷ�Y��{יns6h#l��pY��J�SU�Z��״���Vr�H��7��!$�����-М!g7l�#�ڶ�����P.8��P��U�h�s�UzA?}[Aې'�6�-�"T��	�TM�e��n �q�>m����}0���$W��|.c��>W}�sU��ϸW��^ �kAۑ ��x�Ax��Q����w�|�Bs��W��w�ڭ�����g�/O���p�گ��/��)3�{$�)Lݵ�����g'۱W=u��ZcJ���j ���l���x8���{���qd7
>�����N#Y?���6�kѿ}A�/7\ϋh"� A����w��JigF���D�Ԋ��釦o�T>g#�s��=�$�S���P�7�@��� ���p(�܉�m�`�G�v����Q�x�M�[SUx�s���y�Rmx!���PQ������"}� ���CEv������(�O�&��|~�MFgΠ@�������`��Pj�C��n$2��Wz��|����D�!���>���h������Bɳ��Y.λN��Y�n\.{����@@�@ڐ-��q��������C�`�J�W�cs釦�P������ O�@@^���m����>���
��Ne����q���HLB��l4k<m�b�.u�o@�I�<
�|o�� ��������yQ��-��U����F۶7~�|����=V#̽D̲�9�\M�ߺw)nsĴp/!��������Y<"��H>?}�1��m�����(I]��Gwe�ܫDy�^�C2ˎeX�s2��h�������S��1h-�c�8����>?} /?�D��/�CnD��SU�y�ןl^ul{����/Kh*�9Η�q��'G�Q���雷y���>xԐ�y���܉�n.��ﾬ�P?J�)���>��Gʯ�pMd�"���� AƂ6ק͡k�|6�[�U�k��nV3���k"-+�XG{ςM�e}X;��L�NBQ�Ǧi�ɸs�:��e:7L�d+=�K��8&��_���o�������=d-�Slٍ�Eض����ȹOl�Ÿ�p�'&��Yt���HJ���@��#b{u%�\���#Է��%E�n�lZѓi�򑙰�(:բݻr�x���W9����b�\�粖�We����s�Ơ�;�@	�1#4�6�l6�sr{d)bw]="c�r�M-���yeƕt2v�V��<չ�7�k�f	���S矬3 �5i6i2��tH�Y�c먩��&�BcQ�4������K,�~����7�	m����T3�U🋋��O�[W�}����fc����W�! �B�^!�"A-�����g�s4�^�>A}w��O�o��m�T�����|A���s?}�B~���R�}k��x6�In��̓3j}CD��8����k+�?H>?}X�D6�O�h p�N���Y]#^�����|�R�G�>�j>�?
������n&l��;p�9mȟ7�Ax�ܮ>;��W��K��5��Ώ�c��/O�P@��m�q��˾��7�J@=���&��S7L��y��[��D��-9)��nC]N?C��޿�_}�{ ���CFv}M�%`���S����o����@]ٱ��ր�����p��mI׹;��|҉�d�N��û+r����L�F1d�u����M~�L����P�eTJ�+&��9�S	;.꨻1��.%�{0�#
��'x�o��":��[�_
�����C!>-��������2	{�� Cng�6��Ԭ���}X>��u8&�t[
gGL����RA� [�%���4/O*�Jr��e9��M��W�>_G�/�8*��
~	��D}�G��kfyZs=�q7�֢{,�̫�f^�3, [�8��d$��trw��ڀ���Q�q1�� O�@D�ȟ�ɴ7����~��[/�r���,e���;/���,�#{�v֩�R���M]��=y4/��e����	��m�ϧ*~�}��L���&B����g\��ޅ����[�.�,�0�s����>|��_/y�_��<o[?}��k^Џ�V���Ln>1q�A����]�����|��I�-� ��Y=�C������q/��ts�o��hn��Ǚ�|�G�����{�茧���V L����\���������za��`ykz����B�d�,�ˉ��9ZmDiq1����.	�嚎e\D3,32�Yf~�#��A�"7yz@m�ϧ*W���
���1� ��ڤ���ݛ��F m��E�z2�be��s+U����q��4�v��_��u������B �9Cng�6��i��j�ʾ��^�Cn:��0l�y������m��;m[�Ӝ
�mn�JfH���gן) ��n>m����?�O�������T��ĕ�>-L �w>ݏ7�ۑ ��"�~�Ŷ&~��CϦ|Fr��r�/�g��T��f>�j��n#�ʋ�����}aQ�h.�I���r$�ɴ!��3��N�%��X*��?O��9Cn}>n-� �x����W�A���}y���h#�|[j��?+G�~zb>.&8T�'� C���|\M�Tپ�4d�G�N�I��毎g`mw)��*&�	�,,z�mP�Ԟi�Z1U>�bڱ�Ժ�uJl�ld�9VD�>"j�s��@mCo�b��
��{i��kr�/�g�eT��f> �;T��^n(�m�ϟ�����ˮ]n�4�`��&T�u�3�jS�R��a6QE�������F[����~��H-ǐm
��n}G�>�<�7_���/�.f�}�TH �����'�6��QŶ��1Գ��~P~�W�d/A���D|���������S�@����/vD�q�*���D�Ҡ��į��� ��@��ۙ��h}�n�dӝ��]�4�<�C�t}3	��$�����˙�^�:����eD���O����+xF��~C�Ӊ��D��}�B ���y-�o%��;:D��A��m�!�Ÿ�CՑ�4�r��"#��{\�t{�U��x���E�fs�����e�C�������뱟a.�f��6�As^o!B��Q�J/op��{4Y�J�M:����ĵ��S�W����f`���7�^��G�JC,��M�&��Z'��a^u�b�ci�v�8;tl�A���xp�R�g��ˮ^6�+�V��q8�C����SH��kYGaF�i1\\ME�6��R�v�4�\6]��K5�p�G͊��dI��� �6N��loz�t��ۇ����I!m��5f��+��5����Ɠ_���}���˵��v��s�e��i�W]�_"y4�[P��3�f�[ۭZ6��(��p��V.q>=p�=u���=�;!�mz�����_ϳ�p�t}3 Gݟ.���d��m�o|���jHm	n!�٫c���]��>�/H����}}�r����H'��΀�m��AjʛO�6�@��o9I��p�Ŷ�2�����1��Ȉ��އ
٘�T�� ��>{�$����&6���m(G�kȲ/� GoH��Э�he/�g�]Th����� ���:o�E�>�k���/9������۟7�N���G��pnӌoo��d�W\"g���B ���mȟЎ�o�&z:�ʔr����2a.�!�2-�h����q�"���Y�R�r{n�(�M����A� |�W|"#���i�P>�1§��Woݻg�|����\�/a[Ax���qd1ټ�����c�Ȍ����ܺ�~�r�p6��4�O����$<�UY���񝇶���Q����˜��'i�gD=�X���}�2�g���}�_����Q��Ly��n�7MĔ"E��)[��8CnD��"m	�\b�p����}{n��75�L����A�A C�3����'z	k������m���A�;Ё��^��UWw����u^?k��{�,EL�������5��>z�6�H%�@����=��ʧ�hmo��)p�V|
::�> ��T�����Gʹ�GB��*L��Y1*I�B�LA�i�ַni2vB;�Gb9�*n1����n"7c����h&�"��H-��6�_r;9��W�	w5_	S���Y��i}�">{"|���"����ijV#/n��h�ʄA=���DD_|>ZO">�1���}{�'Ÿ�9�&��Z: 
۹�p�!����f���D�ԏ����n��sN�dۗ;Nk��� ��aI�67j�Ҝ�$�T=���
���ŹJ�w��nìr�١6��o��٪;�K���1����D�T�� �w�H#v������zݵ;f^��dnbs�|�
�y����]D������O��C��5٧��O�X���-�͵ ��Ÿ�70G�EV��R��"+��d����? � ���� ��B\�{4R&6��>�њ9mO��r� :N]<Nk=VM�݅��]d`�%B����c{�5���Cng�6���кC�{�g��S6��W�)��jmp �h/��>-�����߂�F$|9��H� A�5�����U��uw�> �Ј>�A۫��"~��������#�������� �mfP�05p��"!}vV�䏮b8Ez�}E��˛��"fYq33Z.��路�+������uψm	��h���?|�xI��1�������{å+�5+3ꈟNKPL�[��hL����[�!b>���%�ޗ�6=={}�\��/����q»jۇ���f�0���������p�"@-�	_/j��PU��e�|�{�*�]�*g� ��Ј��^n�=�����ͪW�"
AH(�hsE��/64Iu��6�ћ��=��߷�,�foDGߢoZ�A�rŸ@��S��E�~+I�#�3
����?n�C8WI���yl ���lY�����Y�%Ϫ]���c ��:7�uj�p.���/���+�� �j�A�A�`��N%e�o�Z���q�D܉-� ��fR0�����w3y|��bj]]�.e��B�Cn}>!�-�eO�39UNkj�A� u�͵>���|6I�#�5
�����S����]�cN3��=W=�-33Z��,3,�����y��)����������	��8"�*��.je;�X��w� ��	 ������BI��H$�$ ��! ��� ����BI�d�O� �� BHْ���	'�@!$�	%I$��B	'�@!$� H$��	 ��� ��$O�H@!$ܐ�BI���e5�\�=�H��!����}٫���u�@�                     +  a� H �D���UDUPR�($*�R� P� QT���H�%(%�RJJ�P�U��H�QTP*B�$J���Uf��T
I �4|��Y)�)6��Hܦ�Th���rVtkv}�H����*� ���D`S�h���t7�4=�K��c݀Z� �ށ�
 w�Ң�UJB�*Qm��}����Aݽ�{�)w��zj��Z�5�@��9�v=:�`J�'����:5�J�} ��8z齇���W^�Ws��Ѭ��;o6������,�}mj�5*ATEkU8��j�ݎ�:oI8��`[hu�U]�B�^����� � ���Ӡ�;�J\'���h��>���)��:�]>�} j	*p ʑRT)B�(��h}����@<���x�l��(�U�I��@���� 3��F� v��4CA�E.��H΃@C��d��� z �"UEI {� 6�A�4t.u�4CA��� � � :D�$� ���(�yJ���B�16�Z�7U���Uv�      ����%OS&������`���LS��I*TP�M�d2 ����i��PSR 2h      4�*D�ST  �     �J�(SP        "HҦ�F�&��F�i����&i=~������� q��tcF6f�۟E U�����@QP=��d�K�
(��DU@�'��U�T	�I�[_���:?��?���������y�^���O`EH�A��T
-�}G��*��=(SHE�@���D@�)���u�^����-?�����?_������EUU�*��UUb�UUQ���U_�ӻ��r���
�R�� -V�o V�QoV�o� �@/�J�!x %� 6��^
	x*���^�x*�A�� �o ���/D�B�Q- B�
��^)x��(��^ x��� �(�x�AQ�/P�AB�P�d@or�����U���EUV*��5UUQ����UUTj���UUUX��~���N���U~�l%��{��
��P���d�!��^�>�˅�2\������ۊ�����[�s��)�E�]��f#���(�Wm)�i{3��:-;�f�&�q{��{4k���9�E\����� j�E�=1�"q�/�&-�	�9ӽn�	gxs��#
�z�W��"�{2{��3��=�nU5=�x+4%��6o,8��DgwK�� �/�q�������E���}uE Yw���D�+�S���Byǌ�i�DWMU��5���drq�����.�%9��ա��6����G �!�ԛ��q� 77U�^�Ji��9f�Κ�#`���L|�O�75hO_gp���*q[!�3cY{��{{G�xn�"���ؑ<҇^�ka⚢,a�][�<�N)FM�FZ�ɥc���٣�N��cR�$u�{��a����p��
�Y4#�m:6rOw�.X��W�x��1�w�.GG`�r��� �͛�f�A��.��',�U5�
0`�ܒm� YNp�v�����16��~�]�5j�fs�d�H=p�#KA-�a��5��;Pxj]���S�iB�t�x{������i�g-hi�R�ō��Y7�
��V.dv#u�(�Y�mѸ�a%�7��;�0�A�lI�G����կE�z5����7�*�w��JѹƓ&��y��b]���ӹ���Ȥ�e+�Z�N@����=��:�]�8;cX��@[ۢ]5��ʯob��۰�z9vl�M��? OC���Z���;M�I� �'�fC�P�u���,zޙ��.�Mc�S��&��Ι֙�-N�T^�q\ !���7�wt�;b�.� ����S�N��<����2���!1�ɏya�+�sGjɔ7���towf�.y�gp0�pV�b6>�LbhFH��7�\IޘI:s^�}w�5��h9��9
(Ay�	�V�{���m�b3��˳x�u��æ'�.���	6n�G�ۦ��$)9��Mh�#;�[On=�\|O<"B.��GW�=h���u��P�w��삌V~u�2�I�%�k+�\xʣ��&���7�uR�tQ`���a����̻�b�a��s{|�ʰM9��:F�w�ʑ�yc���ŧ��A߈��=D���>ю�YK��!T��tK���՗N��0��>�r���^�E�̰gcr�8,�8c�SM�.�gf��}��M<�,i��һ�M�}�3�uK|��i�����VQ��r���v<Dպ�s�r�ٚ�5'4f���K�b�LQ�_>�qL:�	��t�����Tj�s/lJa���ƾ�iWW��&�Q5=��6���h���^���fl�]h⃫÷ [�r-e�v���-[����yQ�sn�C�j؛ۛl��K$�r���\��Nt&m���o^�i�>�D�ۺ��9���T�6;;A�񉜲C�\���!�-Ŧ<[�&3p�0�6]g�r|��u�\z�5쨷0�,��q���\�d�3��5<�����H�L[����㧓�k�O��f�1�΀�i�O1��T(r����l���;1�oh
Nù���8�,�t�RZ��q���PvDӗ6�8�p��!�6�����:������a}�{�fѤ��C�p����D*���	E���^���#6����=Ѽ�]�f�&�5�������H��'e�7�R��{N�ͤ�\U��N�'p
3�Q�n�5�~�*_t�_i�l;�¥��?h&@��6�O C���{���n>B�UѧT�C���"�� ׏[�Rv� x�T�$��;�6�\C��K\������'5��fM������1��^z�������.���X�Or�}^]9�S%����1^I%���R%]lΏ�gfh��H��.j�طA��:�ӑ����ٛd��u{�h^���Ξ��K�w�-�^0��+ե��H]���թݲ�R<�,�. p;��Kb<��l]Y_V�pՆ꺧/nouE��A�oO^k�_QW=��)�Nw7�ټ��j�����v�F,-s�q`f���b�d#p.��$�5Tu����1>E�K��3r���J[F�vj�Z��&��1�o�mqdԑ�\1u���)ݽ2� �6�`�G]��:0�ď�\@��2�O�K@G�������(�P_���n\��==����Ṵ��{��(N���&���78�c�C�[�q��\�W���胖^�N�ѽ���0���P�0�5sʧe��״���qC6:��(���i�F�����{�`��-Ǔ;h�s��&NO�a�:AC�Ɓp�_��;��X"��ݛ�:��b\"�<�D{{��lպ9��y�m�\�a6h3w�&�Ɨ#�FK�S�����������؆�f�pٛq.�F��㵑�;u[��ulyX�q��r �K}4eǒ��[9����;6q�'�1n�&����Ћ]��/me��Љ8�)�N\:�����nW\ܣ���u�@N�=ɦw�0%����^�wr�U�u�gs������[�v�wyJ��� ӛ?+����Ҕ`��+��Ÿ��u>Z�Ü�t9�1j7�H��a}{�U����1c�.����|�Z<��.ठ��s��9��j�N[��nԞ���[��ŗ�:���6����bWc�Z.oh�f��p�]U�W	6SU �k��6��uk��r�F���vu@�qX��ոٔ����8��e�Q���'��Z��b�Eo f�[�����-�r�߸���w�2�ۓ��/3[(E��!R�]���(k46F�yb�#Ŏ3�����1m+;�i�k�0;FI@�LQōz:nA�˜�.[4��N�|�a���J�x�L�����G^te	R{<��������[����p!��wh:�w*�Ϋc���b3bēyu]l��7 
���{��s�iX[���M�+fKp�P�m�ۦnC<��IN=��>y�Y5�k�^�fvSz�
�erMp��7;	�sV�{T�.)�'��+�.����7Z����3�r��&�6;(=�a��� �g�e��Bc�v�s+D`Lzf�ҵ8HTҨ��2W,�,7rG�����@�H�ߝ݈�;��)�͏:!�8�ԑ߻^'���׸&�)��/a�O�� .7�!V>��Z�ݺ�GL��Y�ܺDekq�\�7�SlB����w6*�G1������y��o At������O~2Ы�Jv�$[�'���ȉ��qԳ@ظ!��!c�q��#��u�^we|{���n���|�m���⽗k/������yW#zbPoO �8E�7�sK"Fj���S]Aj3��}��:]*��j�d:�zq�Z4����Õ`ĸ�5��ݝ�콎��Ʋ��/�;Qk��2Ԭ��ש_ܲ����(��<�V]�R,A].o"r��.������uR�l5hO�W≝�걑��Ť?�=��ݙ���	n֧>,NԲ6��nlgI�EKD�Bx���� ��XR���x�vf��(.�9p���&�!ߖ�E�+cZ��q��\�m�:c��e��n��V;�>�ۓ���J���D��pݛ����{�1�5a��r��Ʈ�(�we��'����x���kǹ�6b�L#�j[|�1܀
v�غ	�mO����j{��9cO�o&UzsR��p�Wmc�ZA�!�ݗ=9�q�%�2�;�0�C���IP�K�SKOw�׽��L=��H^�f��f��7^`�&�À|| �g��啉!h�<��.OZ���i~���bXK
�ٖ��b�&�5����V`��7[s%|K�cס-48�/�������]�v6[���;����5ŞG���ES�o'�T��>���t�#g灯C��oLN�B��l�I�'�˞�_Y;=Ō� �����   2 "�� �$� H�,���2 ��� ��*! (��H��H������  ��#"� (�H* �"� ���H("� � � ($�� �"H��"
�+"�2� �H���"�� �(ȣ"� (2��2  H����"����V���+"�W���������z[��g��`���UD$�Ek_����"�����AW���UIS�Qpqo﵁DY�y迢{��zz�9�폂L^��k:�}����j������ռj���������w���'ѯGM�R>��}�EO�
��e�ŗ'�5oO1B�������%r����-C�g��*����)�U�5��RU0�ЄhT7N���S{�	���\�Տ���8{=�K�&|^�ؼ�s�U�Ò�.���(Pd%*��;���/]������v��Ҭ��1�̚;/���L�gv[��{:x���_K��R�'��{���G<T':k�wb�M�h�o��D�%������kYC���	ܫDiN�oh=�R�������97��Ǩ�{eĥ�9,z����q�|}��~�	�7�����h����m��s�v�3���؝���˹ܡsŶ6`�s�m5O{�����Z����[m�޲�q��۶�r�n�m��%����	���mdȍ��J��x�)i�ػ�\�o��^�ʿ�r�Z�T�qv�nQ�{����3�/���[-��+u��� o۱�9���yØ�#DԼ�%�x�[�i&[؝k���r�+'�2v�wC�?7@�4a�T�aX����Sш{�v�=�w�wBἓ�yc��od{G�9���x�]�o 3`��ߢ1���.xͯ���{^�qd��/c�k�C�K��i5�oO)���F����;n�|�����=�æ��sO�F�k>kh�`�Ȭ��L;�y��8��~�޸�;�������Ѿ۽���$m�F��bӭѶ{�,xnP�����0�A��k4�È�*g2��PqoÐY!ib��X��ϣ;oM���9H������~�>9����jj�Y�y�Vf�ܱ���m��m���fa�ۦۖ�m�m6�zƑ5�	����#�[�w���{���E2�}r��f�@���n<����E�^6Q�n���S�"���Wy��8lk�f��k
{T�y������wlyAȧ�c6JݺMPr��^�7N�a�#5��{;��T4F�w8��q9���X���ђ��v�|�S;nY�o.��t���M:�ԩp���3�sR"���1(�l�N"F�*k[�� ��w�;	�2}y�r�^�_?RQ�l9�_"��^�����"a�{��Δ�Ό�oa}����N�|k�7�@��B�-<��ǁ�>�A��IN�S�6F���8����c���3��Z�0-���/u�Fu=f^�RA��ͽ4�l*��/��T��~S������{|�Gf�����۶�nf��m����m��m�\�݁�p��h����Ơ��p*��tj�k�l}���9��/a���nQ�lg�և��|��ib0�恼J�� q�{.+��Kٶh��C
	f�̻N��	���nN�S)cu;*��Dd�z�6n,��sb�D�9�p�=���	i��W���Q��8C��v������B3���wپ�:�{٣����%�W<�b��f�C�F�TC.��P�������s*� �ZP4�)I��Kh7d�>��J��"$c��Z�ډp�)ΧP#!��mH�ۺ����w�.Y<�Mn"��؍��d�Z�Y$��b���zw=݌��C��1o� .
��hmȘ�P�湪�,���ajEE)����PH`�@o)�0R�(���S�z�%D�����/3[�v��ݶ��vۆ�s32�m��m��m�m�/CRL[(��c%�F:�qqT���]���h��������g��|��3���{5���1���y����䯔�l�&��Y�O9�$g
��7��dB����v�>��*r�ۛ��vjڔ����m^�M����9���#c���ۭb�Θ������ Q��_�e��	���(L�i��Ʈ�E��sm`��8���7G����ts��O)}�j���f�I�u��%�Oێwe;蚾{�c�Q�=����W{Ñ�G���|�\�$�����h�Ò����;@za�pZyh�4���w�~��O]�y♢�ہ�~%�n����Nv�n��n��h���V��p��W5��}����z�o�Z��1���س�?^����	5x�i�$���/L��t��r�>ǉ{��귗aZ�,�B
k�j���3Սm�L �7�Y�4D�;[N��sO�7w)�.@=<T�ˠۊ��h�b��y�����������/b܁{��ߑ��P���jŤ^��6���.�|#���܇7�gtJzYr]�Ж���L:�\���.'�_��Y�������n��(�.��0dBg�_��U{���,������'����Q�K<F�YM�c��'PÃޗ��8G�=!�ur�\�0�s����a�})�q��n�Ӟm�&^�z{gj7�޴� B^A�^H���Z�X���"���v`l�ñ`AC6kk^���EZ(�Z�N��T��k��ιǓs�'�S�
�z<"��w���B�Vo(��K�N�p7��pn���6�=�� ����ݨUn����n�f�h�o������6�Ӝ��S&1��>�6�UZs�.��Z��R��l������aa'���{uVњ����rlȐЗ/iV���2z�)�/���j'�깗�v�^i�S�;�����]�1��2�2M�}���y]�c��{��"�`aBO<�C�$~w�v]oȑb�{}�JX���Ml!��(���bt�m�����K�7=�������|�K=����Nw%�ҫjѶb��DT;���pUa�̎�/���%sj*������:`��w�Ţ�� !�C���S2mb�^7�?',G��(U졺ǟ� �n;�Ë��jz�����=!?[�ݢ#ɟIհ��c7y��A���*����EOU�%��׎,Y��n�
s�lm�1A=��|���L�������{��r��=+H.l�u�Y��v�|VzE��}Ў[�����q�Ƈ���z�z��$>�C����?nsTԧo�;�z!�{�����{<t{�}P���H����%������o?1]�@���[�=ė��8��Q!#~X�x����\Y>+P>B_�dlXw-f{�������_'yT�^"�E�r{�gp���D���|϶{���S�g��-l�H,�G%3/F������8Ɂ��Go?�;=?z�zc�.����1䗩��v�w�8�2@u��Qn��y�f���Gz�����G=���zy��w�B	3w��z�pU�*�זyn�g���s*���(�t$�I�m*��6`|Gg�\�<]8�z6y_v�lH�q�w�z�����:\Ӂ!�Om�mD=4ʹ���fI�w+0H*K�N���P���n=Q�l�X���1��t��d�?r�q/@߫�)�0a�nպ��x�9�?�q�OI[�*����G�ـ�k��������Z�[�� Gdv���1�Z�&M�9O)��U�b����%O֎�j�e�Mw�fyg�;{Q��gy��,� `���獥�.J���9�B��f�\SP�ހ�w�)�=��/33yd���8��V�X�s��.��{$:��"�a�?yR}�L�W�o����<��!e���=FvQޞ�*���Q|�ɜ��M��/�m�1]Z���5?o囼q{�y�eq!�:����O��#�E)�^����=ɑ��{����7B��O;��t��}���XT��ʣ�Ɔ������1�f{����=<�W��!���;��X���ݜ�2���������}��=Y�E�H�k81����"M�7�z���w��56�d�<�dЁ�lD(�7��z�)��_K �z�X@}n�o�"]�(��	��=�Wv�WP���0F(Τ��&')�v�HCu:>ʵg�&v%'�(�Au� ��zc]e���+X/��W���,��c�~��j�j[|_�/l�ڍ(=�q��p�f�nvm��=����I8��3X����ƽ���7
8�w�/c����p	�<��'�
�;��N�M-�C$�NorIQg�,��]c�˝��Ǟk�o1� ��\q���7|���g5v��|���E@�Ad��R�b;�x!��w������}x{�\�z�.��a`�O�����7��<�'�k<�i��CV��-SU��A�u�����9�L��B�nb8�p�Pk.&M���U��.�uL�m3�W��"K0k�6(ؖ�ˣ��v����� �R�������/����;7\�f�hM�M`�řb�(P�+p��ذ�����B���uԺ�,�.֨�D�)Qɥ�]��r�d�RSU%�T�l\��ܥ�K4�DS��l���0��e�y5�e���a��/k<oo��9t�BІJ͒�QcdԆw[���;(�8�С`��n5��)�J�t7\�05az56�h5Y\Q*gi�b4e6PTn	���eԎ,��	^��a���ҍT�qTh�Ս���	m��%��W2�J�@qa��рK�#��V&&c�`B�%�.JgS\�k�5�B�镫vS-�
f	{^���e.��f���VhZ��0aQ������\B�:84lf:h��܂�%���L�U�Q��M]�Y�44%b�v�����L�q+�Gq�f��^�B����|:����#	�L�M��������:�[I�-��5��sn�h$!�CP���#c�ڷB��M]"i�	�0�q��x��@�K��f����']. ���\�y�l3P��f��V֕ɶڳL6���ֻX���ut��)��ؔt\6S"�LP��A�[t`Xl�P�D\�Sl�����d�ٙ��b�d+.ѶT���G]�*���ȅ:�\�,-Fs�\�dX/��$�2�����uR�K��7`[�K�-*�\�fM0�%�P�fS�RZ�tW��+ji,ir4a��˯2�`��D�5���9T+q�ܷ)X��[0s4WY2�K�0i�բ��(a�I��v�qE�:c1`╁��r���d�p ��N�qL��c��;�%�k3l�!�X��۫"�Q��d��ʣ���m�pekHKL�����6[2!f����j�V��9^��Q�̗Y�Zh��Xx�yu�����yЅ3nVۺ�F9��vsc�ॲ�����LƱ��n`Z�[Vݱ5��-��Zm��[�c�b��6r��j�m�Ԯ���8�l:��መ��Y��[��� �1�!n*�����Z]7Vf+r��3@�j�Z�ef�W�X"7Cr����ř���]�4n�F���vB�v����<e��6;Kx�yKs�*�c-�`bW��%n��B!#�,С�<J�&��fְ�Mm�n�f��{L�c�zU+(ݖT�JV_(���&)]��1�f��W5�(�2ٖ&��.�Xʳdu�0uZG6`��mvt+\�K���븭u���۝P(�0ل��[��lA�K��U�,\mD��i�����('ɑ����16ѹbK��%r�
	�]��9�&���%�6@M/�Z鳬��F��b�#�ٺꡰ�&�I��g*`�)ֶ�JL��k.f̦�)����@dN��F��q����G�0S�is�<��x�[A��4`u�^�d1�`��mkM.c�L�R-0�U�#�D���4��/]�.�&k��\P�xm�X�۝Ɋ�U�Z��3GX�֐-P���qK���MWB�F��٬D�t%���5v̥E���%Զi�����"L�$.b��V�UÞ[�c[3���ihD�
鰑��
�-Uu�b���عk�4�%�уu������y���
�Dn�hX�nn�&��0�ԫ�qfu�gXA���!��b�K��1Z��GB�,]p���9�Iz��Ti���a�����Z\m5��� �v\��R \!j�Y�`P�3���A̲6�;0� �x#j�E��v�Ydm���,c�bMvJ��MĬ��1��c���ƼP��92k^QUl�ʍI�M�v��Z�l�ݜKx3k^Ŭ��*��ڰ-�uٶ�em�i+m��53�Ѭ�4j�@fR[2ڑm"�2�v�̻`N)(�7EKV��1���؅9ٲW�MM^Ê�
M����QJ�H\&n�a��'�6�f::+P�s�iJ�p�:�a��Ekn������l�F�b�bRK���\�F�)(Lr]�4![��m6j�M�t�Aҭ�W�T����h��a1%�*#�8]��v�"�AZ8�cc,h�YZD��rQv)%�0E�[+��W��Z�c+3B���Ѯ�]���a�Pf\[)U�7�� ���XR�Ħ
e�3J0%�k���eێ��fM
�qi���Ƒq�ɳ.s�^bZK��z������ұ�x�%��%!��*X�]�0<,ْ�5��1FiT��i����Wm�bKY]2�
2�\]��7||�@�9��mW���]��k5t�T��9�D�tKu�l1ҦF5���b�RlLԵEy�2��mm�qn���n�l5�5����@�b]q5v�ћCh(��z�F[�`fS�I����20ff��2�&	a���tj�����X�L�v��+�v�Q�U��Rݡ�;#���pRW�ۈ�)U6��
ڹf�h��z�"�t�om�n�����.u�m�Dz�-�����21��͒#�+.��ie�a-;���]c,�Wa�2Ui��ۘ0���\��UW"�Y�W�r���2�3�۔��#3d���Z�(E�z�:0�	�J9n-6���n���яtvu��ʠᣐ��Q�*�UUUUU*UUUUUUT.x���8b�b[)�1����"���4k�6�M�v����^F`�an��f�'h-#�-���h��n�c3C+J�e�����`+��b�1`��"�!�b�K.�g��7����{�{�%��=ԋ�R
H�~��$y�x��̭�o=������bEDU��	e��b^�>Y�>���{Xu�J*%NCj�MW#9�#�n�6��LB ��ϟD�zh��6 �
������d��Q7��}��*��3�����ԊՖk]�������L��x��t���XE���R����2��Ԋ��Z�O-	Uц���\��F^��1O��yu�+���Z��YcaK�2�F8YR���#˒2H"+ˮ�Vv f�t{�x���#�� �;���ſ���=���b;\�F�9�+�
9cf��7
�C�i"¡�(�t���т�U-�qNB�nm�Z�0sf�S)�۬�ʬ���щ����v�e1R�`�t֦u]���lc���+��u��VT�R��#E.�KQu�v��є��#�nu�b��M�Q�`�q����i.|�[l)e�4���A�t!-�J���qn���c9]��i��SQ���7jܕ�b�Ԫ�m���s�����c�U#6�`�h���.�u�]�4\�L����Wi�J��YZK�R�ŦJ���[��j˫Ps1���J)Z���G5�2#�*���3k�R��u��M�4��S����ō��g\�h�bǀ���r�B�q���A�Ûf�sJbZ�.�P�aJ�fȨ�[eq��^���Q���ڴ6#6 mW���(#tk�eQ!Yu�eF�e�Y�s�]��ֵ-D�dc�Gk�n�.�Z\��	�*5T�(&�[�y�u�[���+LV!��jʭ�t*�Zd���*��SgK��J�;��)5q7�:�t�F�m��Eek��*��%�[-[iP-acW��V�@�A��A�,��,VJ���3e��1B2��bl�F
�+Җ�e��J��Z,F�^��/��?��ECa�a���Dc���w�~��ڝ������SU����։��㼌��3J�Q�<b��L_��<�Ǽ�:�ᥤ�V�n�F�lMS�}�rW���n�>���r�j��g�Mdn�5US5[�����ٿM^X����,ce���p3��[��z�gZ<p*����^�B�6ܼXpD%�NbƑ˦��k��|*������1H���\���'��)�s�ߟ۞c�7&��#��(��\a�`�j>������\q㝑ODE��1ۈg!5W��s��z�Ǯ�t�wSwL\�j���kR�'�v_?~�ww͟�ْ����{���Vެ����f���B���uz�R�B�C��5��ɼ�E����{��V@��<��/��g�|s�4ZB�3��tX+P��A܃>�?��};���G�� F>���;���R�D�Bw�7��Bn�w��|�f��#H�Wx�C���6�UEQ�K&"��莎�y]�2ј�Wsuwצ��e쥽��:�Bх�1��V��;ӽը���<;��UU���D�� f!T�]6�:*���y�a9�:tV,�E��>�uӣ�;��ܓ#��&�Y�|;��\����BA+��Uef��u�Z���ꪪBf�4_>�=�"ku�mR�̟a�Ȫ�95�97�ۮ*����� Ui���UQ��E��k��Q�[�خ�ǝ��SH��ݪ�*�m���;��e�l��Ow۽��4:㢣!lC��p��%�z����h�_�A�c;�8�O_���n>�*����:��[^g�H
��_��#l�S1��(�8�ƵNE��r��tH�k��*��n�sښD�[�5�G�f�����wn���]�[ג{��U֒�j�Ӄ�`�FT���΂��췱V�ݙ}�p��������_=��{OCO#�瞯3�Rj����_bʞv���'��]EU`��p��Va�Qy,�iX��>Er�c�f��5Ȱ��/cr^�N�F�v-CF������Z�V�i��0�Һ�c��b�i�5�ű����"�9�kP�H-�4�k�`�p.l�ڊ�Vm�)g�_k�K�v���vr%�s��㊶�зR���ljW1�u�g�w��+���4q�6�����3�V9�g���l�ٓ�z}���Џ����O)��Yv��zc��綖']��mU#�v��pSq�+!i�F��kz�"v���}�xwq��g�{2_�ޛܱ�����ϡx6��)�`�[uU318jD�3�n^�wmU#�a�UJ���ӯ�3:I�q=]�u�Z:���b�9��ԩ�_���R{�>��P���jn^�
�W�n����/b����XsD�nNC����~?>�=�5~�m�{�Z��@I��p䩂��2�ۆ���.�_��{�Z<L��%W54B���C��)��}�-���#�2߭��jƬ��9��5�]���p_>�=���MH���J�=SQT�A].���6*ݣ���!�]��u�w-Yٜ��&`�ϒc��ZK
�h�*�;>~���&�R3�[�uT��
B����.n�ު��FN�_N��Y�f�6��%���t�N���U*�M��b������v�����q�U����ziW�g>� ��v�˽�ثv��-��C�.�ڻ�:����ՑT������U#���z�Wm�,˹j�U�4��V�[�O�\��u^��S��$�g9@��X陏ABQ��:���F�a�����)���ۚ�}o�ϡ{�N$�����;���a��o���{�j�6ky2�AP�B�R��Q�Ы���U����3YUCn�q�m@�BNMe��}k�u�QS�#39	��')����r���"^�oq(��g$U�ۉn.f��|�`	32(N��w<��uT�xa��mO)�r=\>@��b�Af��	,�`-77�ۭSǏR|U�����o�{�����0$�m�+�)v������_Z�������7cv6EUP*��O��UH�9U@�:/��@�C*�_>q��'��_oF��|���I��W[��wq�D����ڣ�7IuN�1�Ll��)"����s
&X�ވ�,5�����u�L����,�2��)��� i��],]E��E��(ˊ.�(\͊��[�4XG1��5��r#�.Gf0
)p��e�D�RRm�ɋu�s�fФibW:\���^͵�sp �VS0J����]��ˣv|�>�e����6�spl[*��L	����B���ϩ�	8����uT�\uf����UE�<(�mK1W����G�{���z�x%�|�
s"Z�����V���֜��+�H"�a�DoW; M^u�n���\�P��bL���Oݼ������f�Lӊ�x�f-hS	T㳮#+M]�(�dD���9��`N�V���d�f��a
��[�}��<ѹ�������ָ{��mǫ�.���|��X��C������z&G�dH��W���$R�y��fw\��T��IuE�=��Gb��u�^Y5�K�[�r&#H�����E��v5y��7sH��.f����(J�>?o�9�7t�Ҵ��w
[�f:���wߟw����3���v#���փs�m3陁&,�u�{6���鼳�י�yȴY�k����=hiP3@I�|�v���T����5k���I�1�3�!��!]���K\=*�D5?v��iJ��ĺ_�l���H�&e0K4mjQ蛈�P�h0�]���^_W����oE�^�l��3�T���uW�]N��Ȱ�Vu�V���rqM��B�:�AR1�7n��������*,��ҫ�P���)ӽ�bB�{<0^��Cy{h���fXO%��������V��A�жl�*\�*�[3�
�E�^�G�m\N��힜%wT�.k��]���_�K7n^�Z����"��p�����L=�q�h�;w�>j���P�Z�Cw[.X��1B�.m�Ai(N��#�L�G��j�.�LhcP ��DTu��rb(�B�T�y�1)؂\+η峮?�=����~�v�,k��ܫ��U��V�`}���D��V��2{�&��"�Oz���"�U(/\}��z���E}E�>K����қ]޺:k}����'���ϣ�*+ɹ��V�>�%ˌ�7`�3/Z������~#0��r���O�7�����O��%����?5�Xyt�n��*;���`ƶ��{��{4�f�}�y:|L�a��W��.nJ�'̲c�Xy6�L*���N���J�2��l�X�5;X;�.��ִF�j�a�e]J�	CD�Nh�nJZXu;T6��K�y`��a�=2+0�Y��ov�:�L�Í.�(Md���
J�"���E������|~߽��}��M#�aϐ�^�*	G~Vr���S���#�n��>���	��������������Y_wݿ}7�xkA�PV��2��~>�Ｘ3���b��G�	�"$��1�#��T
=�����B�/�e<)��W���X`��΄�F5��q}�rw���U�6[������C�xH��t�Y��*��#.�
�L���2]�gk<���Ӏ'���t������+{��w'{�*���!Χ;�t�Sۮ�Ñ."�rӉ˄~��'���&x%�Z����W�wT�4��fL^}:.��'����y!�L�a��k�֋U�m��|���8��=4��f7���Y�9:����p���*��S�`�Y������~y8�a}�S��\�zy
"�#u|�G}������ꚪ�|�m2�}��Ne����l1�#(eg1��%����^������~_{N��$n��|2}+ �ic�ʊ̀�l+f�2��\9X��͌�ö����؍����<D|<ԪT�4�#m�1�\�]�sQ7�_z���ae��bBe��Q�+WD��ڮ���Ep�C$�H��SZE14% �%�r��Ƅ9�]��4e��wl.۰@��[�J�d���<�플������Q�à�kT2��L۹���n�u}߇4,�7�sq�}rq�6��`dO�U/T�t�r3��s����Y��>�-�?4�hq���VT@���oͻ�G�妩Q�B�O�D�l{q��y�q��Ï���2bU_�Gت��HQ���H}æ�^޿��Ne�����ƈj�k��C��=w��ם�6���:��)	�1!D(�i�¦ik�m���s���ƺ �9�NT
���Lt��r6��A�757r����
��w�����"ho��T�騬�����77~��_xN�g|�>�]�|j�P�~����qET����fZQ�=ٻ�Ne���~�"�n@���ZY�0i���}N2�t]8:�޴,�΁v�q
2UU�gs����'��)?W�?_wE֡k����A�&Ec��uCkuv�b͝6|�����T�/3���9�xN�G��^ҍ��U�wRX���>��Ͼ�ｧH��g>��KU*��d���[+�>�ɞo=�.3R���z��~����wn�dյ��G[g�v�8�E�u����4����4fj�e|
,q����u'c��s�̿�>�d	�9��j�˟Y�R�O@�ֽV�Ͼ��&g���(�~$��8����L��[��`���p"'�'�b^�*�f��#���OI��T}�c^��5U����~I��������������v>�y��|�
��Fw��h��f}�umZq�G�n�b��q@�Q^�������R�u :��Z"BsH�Z�:�����P9y�)�s�y\�y���>g�c{į*u�~�v�8@�t�`O���2���ޑ;ox�����R�Z� T �!��L�
�,��P\ ��f�1@j������QCG/�k���/���D���m&��� !� �s]�u��-2��S2B^2%d����4bʬ���$�I���$B� ިR�@� �[�����:��@�R�j��{���q0��[����9�pDLU�η��4Dm �!��@�t��w�����;�� �����1�@1�uZ�Z�hdKD��w���	G��H �Q�����FwЦ�5ֳ��*"/]�6"'PR�<��Z"H� X��9��:��;�肛�-�"�L@w�o}o�c�k��Z<`�Q��5&w����i � Z^H�lPH�& �D���˾�=|� �^�k����?x ����DƩ�D(�8��/���QӰ������Z4��c�
�-K�0�6A��p�_I�\�n�ҏÏg���#e5^M�]��\5ݗ��ͬv4�4��4ٌ�b�q1�m"��T�m�Wi�d���7:�f�4k��
�u�P�i6Ү91l�f�\�j�#Z\V�R�B˜M+�s�6�7Ͽ'�����Fl�݊�q��E����t�ݓ�ӠI=��N�c� bqKk�}w���g<@� ��G}o�5&���DI�;�1H`"TD�C�-ʭ���:+h� 8�TA� uε���[]�^�G��5:�1@w�%V�U����Z ���6"$�"Q�����$
�<�*��TE:蛈�γ~�*j<`� 53�@3o�R1Ax�����l��GdD��J���A�@���=���k9��D��m;�u�/��Α)��DA��b bAHD1���R%�8�tk��uZA�@������c�k��@7�DN���P�@��)��v�e�L�BT��d�L��+���c�55��m󤅆ȋ�P6���D[@�)��;��}��ۀ������&����'[�� b jc".b5�3>~�h��X�Gӕ���MU���o�Z^N8�q�9�j�P��17�8եnwk�|���i������9��<�"$ w@�"Ct��qu �/��e�R�`j
� �� �E���x�ևv��ַα����y �#L�Sȁh�sHb�����w���T�l�A�ߝ�j�뚷`�D9�Td4u} ��TS1�@/
1@�Dq�6��b�c����3�k���x�s�D��m&�@���)��3��:u\�����F��vuzdYs�j��ֿ@QD7�B �$ +~������>�R���[+;P@�:��@d��b���D�ؠm1��\�U���/Q�u�	�[ֳ���;��
��+���7�dKD1���w�D�{��D�A�B1H�� Y��ѸOBP�-WDEW�+�>��Ѽ��繾�{�yz�ķ���sT��S�M��Y��n�r�?��gw�}�m���xDH��ۥDI���e���:z��Q�5 ;�5���sc]�^�8DH@:�����W� �@�tdA��6 �b
b�w�u�:ќu�N�uj@�;�:��;��
�<�w�.@q�����$��{)>�}���[��(-+v��QTΨ�gM��$�oI'�;��:�TG�-$D
9�3��s�x�P8�Nru���9�dD�D��p
��1Op[�݀7��@%��u�QWDM@
����\�:Ƹ�z�qDI�"Q�(	�W�*�w�ch=��Q �h�Hb�(��Q1���V{�7~w֭�@�D�C��gt��".��1Ar"o=�c�������q� ���}�u�}s;�{@��� �x ;F��ם��XT�S�a���?p�����iɾ�/vv�綟;�ٝQ|�gW��$��{͑<�� ��甁b b�X1�Nw�*n��Lg��k�]d�2���B��D�{10}������a����39Ĉ�~�@\���y�s��Aej�|5�{��7r,����V2��v�׿^՞�׵Sqw���i3ҧǅ��uֽ��upxi32&�Fݏm�37����od�';���ʹ��L��8�V[}s��y����ڳ�jf~���� �����!T'��[L����<�~�x��'/`���F�S���ܠ���9n�-���,��Ś*�&$_��UVq�1S���R�&9Z��4���)I18ΩE�쮀&Y�+��ϧw<�r���.ck�E����U�p���+���Y��|�O���͒��ʾ�-M%�枲H�T�Aq-ƿ�i��ɽ�۰n��gi�P�δ�jb�1�-n�	��@3bۂ�|ð�������ٌ�ǹByd���su�7�/��K�=�I�_��}��/V�0ľ�;�sߺj�����@"�ַ�똗+��@����c��_I��/�ї����Ա���S����@>��Qo8����pٗ�f�ݩ͌j�p�rƗ��Ze}�ܾ҃�D{�!�<�c�o�����s�9b�������=^#��n��;��:m4�����w�n�e�;n��~˸�X�E^QR�Z^�rw����gd�!E	O͹.v 郩��1L؃�b��+��?~����cW(-gD�h�]����T��Y��Ͼ� �ZŞ��ёQB��t�*�+�=p�<�~~~~~	�ݗP0L�%�g:V%��M����}�=�����M�8�M�Rf#cai.R��	�2�%��(d^$N\��ǃ�	�t٨b5k5��#[+l�-!�� �\QA�A�7W^����yѯ_ �0nݳf�X�9�겊���հ��jPKW��kC�[7��	.c�Z�p2Ƽ/0���p��j3��m�k���Ka���141�x��n���J^�a�r�	)-��k<�<�rh)bt5�)�6��^Վ�����X�Ƴ-����c�	F�v�p\�&pZ�ƞ0�jbU,�)j	�ţV�m��J��F�g�Tm�g!E�GB2� �t� ��CT
�+6�����GGGA��ά�s
���)k��&�2�=�R1{�;*$����]�fJ�)Cf�bD�MX��k��YW)��mbL��������@`Ssb�V�[{L0�32c15�wQ5��e�`�
ĉf#����m۶�]1f8e�sI���ɛ)Tz��\.�M�fe�%�ѳV0��a6�It�2�gJ��L�GmSY[E�l�$�m��e�tY�Vi��6���yMp=K\��뀴X��Z�)���	�h9c�l"5q5H�׀�Pé*�f�Ka�e�Q�q��3��XAF�XiIc�kFi���u��{RFJ�h��q�4a\�
���6[cdՅSAe��b6�Z�+�j4u� [���+�9�v1�����J�K6��hgE�7=�h����km�u�૴UL�3r7%�0�HS0ʪ���.n�"J�+�%1ZW
.ͯ/?��r���q����})k"^�vv����m��5D%Ѭu ���U�B髪e����*À����M0��f�5�#��`����ژB��j�kk]�uƭ�*�Ma�����hk���6�3s�ͺ9�W���{�������z������ы*�;>�i�ܺW�[������Qvi��j0Kё�s=�ە���q�FoV�U�odd
�雃��pOt1=�$̡(f,�+{z�����f`D���'s���}����{���� �eݣ��P�P*����;�w2�+�����f��9�a:;�a:g�!��̵R�<�r:�Z�p��bd��HQ�;{���Y�IEf���*�@�8\�Nj��Q:gRh�F�y/\����
��c�z�:��s��u]X�<RDd@�Y �/���}O3�~�9�W�b��;�°x]*"fn�J�7ܲ���x�2+��35f��g2��ڒ�r�[�ڳ���-��q�zff����~���}���S��Î�3�I;*M��z��~������J�FR%���%IX��T�=y�����S͜�}��7$�Z��1&g��Jn�s�J�]��oo^՞��EdI��e��q[ԑ_-��t��>�o�]J�a��\�"�~�\$���)�L�l[r�x"��*H(�zuz�}Nr��j���;T#-��kO���v9ͮ�G�&˸��qL�MT
�R���>{����kCL����������]��v�%���`,�MZ¦$B�QNej�'#j�9��Nħ��"�u,�.�Aв��:Fe��-�Vm}�#��x�l���`�gnfD�R?k���׷g���&@���ρ���"\]_׽���q�l���bpr�U�YJ.�A�-�ux�+��>�{q☨�M6sԀH�H# " 8�3�9����U�/�j���YO�#�g׎*�#���O�>~��5GC0�t�2�n����3Vl���'�ȶ'�o�>�]vݞ�6���2��NGL��П�x|�2�m�;�G���jaao��P���}�h��3�U�����$I�\ƴ��g�wF�F�]�k�۳�Zڽ��`�B��H��W4�1v�_;�E�������po��<y0&�����7&�����/{Bw��{�u�MM�%u�7�g�_ �"$�2
>w�K�,e�E�K���X�ݬ3�������B�����1M��dM+��Vkv�e�iX�q�#�s@.�MA�XvX�"�i�,��\ܭ��+6Ur�l�/&�]U�2W9�~�<3�5���~���՛H�R;,�R8�X(Kq%�����������O���t�ĩ���.�쫿��̮�{������|i�p�I�2�̂�F\�]������fbeVݲ�f>DL���c�n�	��5ћzt�TQ�FLMw]��J�u�c�ܳ�Zr�s'ڲ�"�KRT���-/Z� ��Pf��0Vgg�:4z2�q�;�G�D6
c�N�x!�6C�`�{p!�����Uҗ���3���9mcbbyq�s]�E��(F��N���E���k�B��VDBA�x@����/��~�V�������A�����q9�����:{�{Zfff}J�שGn�˽'N�ު������ˆ�t�T�L7�:FM�Fv�]��'�JO��o�\��ЬҖ"-�o�A*�%�6�V卛je=��O��O's3z�r�V'T&���&d@�c��C�y�wIz2�s_<�E���u@����������Ľ�'�O����'#R��U/<���X{���5��t��ݭY��X�V�z���dǊ>Ad'����{?7w�����X����*�r�U����|������;f%�ׄ�~p=
�酔ʬ4���w<�Gxi�S"s��������v.h�=c�֙Ni(D�2T��J*�嗐�2�]>�vﬞ�b�odW��N'��Y��ѤgM�g9��k���}�������S�ffe�m��{��f�� L�u�����)�[��n���ϔV=�ot�G�	�GnQ���(w/�^�`q�.<r�ޔ�3��������߈�"��$���|<���{�]vNᙧ��*����~��3$	���؁,�����'�9�v��f�Tk�m�L�HJbD��#4�MzmVmfu�s��xe�X$�v���4%zfc���\��g�������o�'��&�ji�VD��n�9��
2���5�Q�փ����U˕��F��w�Ϝf��*�)��t�Ⳕ��p�����l��n�o����ڊ���rCI��"��ڴ��8��ğ,�2=5{M�3�c6J��e��tƓaO�x~*��$�������eU�U��f�����ۛX��ܘ�/e��2 ��eٛXi��-�mP+[�]Jl�b����ET���X�J�X�3�����ڃC��H�!vf�D"��+��m
�����3���*l,.��ߟ��ms-�f�P��]+kf���f{?E���+�Y�t�}Q���\F)��7�z�s���뛼��q�O}�d�Ii�1H�����I����#�fJP� � �K%W�}�ߚ�;����,�� �6�(��.�ș��}�3	��>�/ς}ߥ�h#�!�hG4���b8D:�[�6�#���������kk�$t��r�S�uMb����u�fז���+Mt��04�fj#��@���ڨ���E�F7��2cW�{��}��P		 AϜ�=C\�{ֻ�ח�{�/�]L�ދ"eI�o"�*�s��y�4̡2�������:��NG=����w��}wW�}86�����(������t�k\GR���*}g��% ��!x�CQ��j��`�gg�ɏe�2]��f�q�O��m����&f(I�t�_y�=������fzY!@���HW�}��=�ڕ��1�,��a����n[���J��ل�;b�܉f�il��G��D*�X����#�{9�p�>k}�E�L$R̈�}?x'�8P��ow��m�]�{�P���9������
�Ġ���F���D_f�i��Y�f�iQ�=�|7޷;k�9�,�E4PO&Έ�
v&��Gh¤�jʚ���S�%���ܪ���ܪ؁m!�����sؽ6�����#������N٩QRu�#�+ �7W*�9P!Êi@;�7nkAq �J姶��;�7c��D�R�dާ݋0�c=��R��!���e��C;9��p�rs��m;�Bmǝ�����8�v쪳V3R��}y=���$��ZS�%���$E���wN�U\�x�v�����˗
@�{�konm�΂l�2�!�i�[��o�8�:���Z]ICtS�s`���W�((E`�5ق7=9��^����$�@}+Tm+�l^�~���[�����R��[l��-ے;����HCz4%6&��fW�α���+�Ra��D��x��;��9��O??=��쬪�w��ZƶJ�ظ��tK���FԂ��w
n5����EF a8.��&�bˮ������r%.��%O.�<��������lИE!4�'Z[�i��l{�r�O7#�BX�����̈�[=mY���Uh&F�Ho`����RضrZ�N�(^�rM�'��\�̬�����z�|O/�zRŃ�-��f�7��-�0�G�>s�#d܎���h��z���Ǥדw��<����r�h"�L�ȅҫ\JJ`4��KKIB{Cj�%�~�8?�^������������*����מTU;�󗳥��]7}z�q�OSB��fd@��6˪��KU/9���s��Ӯ�y�+f<$êYr����ϟ~f���1@�;b���
L��ɮ}�1%���s�ޙ������O�vnq+C=�Z(���o�f��ڣP�vN����&�|�/fw��Nng�GVӲx}�&��u���׬�b��y��+�g>D����2|~���q�xGj�my��`݌BU�N���F^�j�*h�[y׀�P�D�FE ������Q�����Zþ�������x3�0&"g���6� �`L'�I��j��,s]*Q��j��~l������cn_Y<,IU�����3X�}F���^_��ݛ�����_�3:9�c��n\�&~�����\n���9�����5Qкv"�8��{L��G=ɹ�s��2"�h��Y����wL�!�7����zg��4ə�+)�N�ܫ��a�k���1��P픕�0d�K2mQa{<V�	w�D�����@K����		$TR��Y��5b�Rҭ�a�a-Kq��AuW\���3���ťRVc��!�4׌�	�m���bTڔ*ꖗP ��)����ckq�1@��
��FV�T�VלJ��j�̥����s0�]*���p?�������F��ٕsZ�����vc�6g��+%�oVfv�s�O
�:���פ]G�T����.#r7jo{f���}�͡0��j"��&eI������N�����>�T�ӣ#�z�y�$WM���9�'�� �3�5�~H�H#՝��w�wvͺ�'��BHy�؞Z����2����5�U���.b�Z�3"v��t����GG'șA�~�C�OG<5X�*tQ��*�:����_H�	Xf���˧a�s_��	d$9���r��^o��r���2�(�3u�2�z��)�Gm0�f���<'{u	.�T�|��Y��#*�(�ڬ�gD?n�w#���>mH2}3'"��u����n���L��{�|��(ة+J���m������[�-G5.߲1#��w9��O�;߻�ϦP��+f��8٬�s:�{Ú��e��r�W��(I��V�k�(up��Cvl�� �P�j��
���.�YP��n�	n�ϐBDI dA;�]��{�:�s'�q�R��P������T<���ƪ�r���Ox2s�HY�2Dʒ��p�w7ї���;�=���I�̭���f&F֏]��/ �jZ�Cff"s}�H������.ɾ/!Ζ�j��y��7v5�^vݺ�'����=��ʹ�ϖ�س�j��.�^�s,mT@�n���!D	*��5�ث'�Ⱦ�G�>[��\/�-�5v�^4gMҷj�r��ou��4��R�P? ? !",� �w����,_��~U�n�s���W�&��r���d^-�&ckS���7Y��[{1�5�12k@��f\
3W��g:g�,tc3ÿt�Uw�����1�٭��*���d��7�li!�P<R�2�5��S�x26�$ȕu�fv�v!N�<ΙΙ�a�'����uF�>�qC1M^���T��fWƅV��.��C��=�;���6���m}�n��}�<4�o|��"H�"�7���fѴ˅e 0dU�[��Z���m���\ֶ��� -��vQ#�Е�Z�8K�kX��v�Gf� �i��͸��R�4Ă���i
�.��+���LZ`���
˫��6[�������5E�e	X�����3�llQ�Z����>���e���w
V���\zL�^�Kmi�I����ھy�9�=�i���l"��1b[�o8��W�߻ީ�>�fL����p��nZ0d���U��2�	�N[�3N����Dg�T��Q8�EGL���fn�3�L�潦H�y�s�g;�Á�\.J�-3��rde�&"D�~�eyn����5d�pWb�\�l�Lt2vz_����-?)_O#�^�����*'��Y����#������⏐ �@�VDo߀����>̯�Oy��,8�8�b�C�.��܋�ʡ����2����U�33/�T6U	]���~ɻ%�����;�}��T���m������'�ڙ���97��w��/��lj�vȱ�PƵaGuh%�Y��7S}��%w����w�!;ɍ�T�2��H�i�<ɒ��wُ��n��v�Uk�#��h�ə3;3M�ћ�Vm�l��Pz i8�PP�z�-ƬH�Nf3v*]M�Ʌ2�8�ͯ�����"��� ֻǝ����Ry�w�ؼĵ��N0���K�t�_���>�ze��x��>33q��R�{��ɻ'�>��$���Z�}�A�C&+Ih�ٚ:�]��\ٗ����G1"�׾��B?bX\�������s�X[�������;��y!�rS�
J����m���>����R�����"oi��9�Y�mU�}�����h�9l]��l2�!��t�^.v�ǖ�<Ż8"�V�UA=�[�[�O�=��EYdR�xw��g93���V��m��c��gzg����j�&��N��tc���40E�[,�b$D�Ml����ѹ�7_�vNY5:;�BL��8�7k��qW��ӝ��:R��ݱ�fb\��.v�������m��U�e�f��gm���練��Z/A�N�e�4fW�U7�d�⽋��o�>�{̺RD�nG� V�E�D��������t��7��f�[Ai�[Ya]Lc��s��q�a�#����E���sO6v��@����k�py'ǂ���75�%�k~"�'#t�5����8�`8m���~����6{7'YfՠҐ�%���9
=V�.��]7yA�e���B&�#S��)�e:|�{���x�i+�4[�_m�۝ =��S}{�G����(\������裦��o�ugxp��p{E۠�֨'�OY�dV��{(�m(~�t�N��A J�zw6��1��E�R�G�pP���q����ɞEg� (�O!�t��zs�e��wDU�Q��\U3�sYPv�����.S�w���-�=,��f���N��Ɲ<N��w���A���l�a��^�_]/�'cގ�u��Z�n���<&�n�����l�/�m�|ߨ�v�����O�';�xf��<�,h���C���h�R(�q���+��Yu��k���uc� �8����=y�,��x�l"�l#+utC�s%�v4�N;[�-z��ׯ~zޡ=�f�n��%%N/�c7��,�f����ڼo0��=��ߞ��V=��v��hz�ܛ�,u���.�6X�������>[�߿>���fb~I��V��!\���*�̴�(�(4�f4��(J�y�iJR�J{%&�ok�&�������8ð�v�:�1��Ա%��ať�Ś敍��-6ؠc�1&l[԰� YZV�m���S-�a�1{ŚN}�/!��:	�Y^�L3ݛL$��EB�\��V�L��D7y��dj[��<�z�������D���0��D�2��96�r@�J�j����ld��S��Q��m�V�ns�vw`�c��������u��H�1 LP����I���-)YE�WZݵa.jH�TYk��Kn�4�M��יL��c*�n�X���5n�o��b��lcT�U�F�L���[��F�`!-�wa�T�#ba���q-5�Ѐ�[�M��ơ6�a�,AFk�\i�.�)Kh^���TM���֜�s4F�g`��5����ט䴅�����l�%�W9�-�M�̸MÚ�M4��4�&]�$-YM�Ѕ�2i�(�J�M�K�	u���T+c]#s]�e�
A�.,K��8�ڌ�*�ť%��Ja�F���hMa]\�VS;��s�����)M�^cK*1�M3$"�f��+�8Ek6+3A��"��V��`�Q-6P8�ݶp�rШ[��9�û:9lp���M5V�7���8�+A��4�Zf�Ĺ!�E�G�2����7;f��8C��SR����մUuQ�E�knE �)��m��mm��EvQ�kE�Cg�Iމ'� N�S��<y_[�M�
��2xj1`�K,�a �֕BX֖b�B���%������9���[�)�o8�;[evcƱ`�E�!�M�K[j1P���mvʄ���[\(�0��՛j;B�������̺!�]�b����2��&J��&K�@\�U*q7����L�&n5OXg�D��.4��"NC���윲x�ff��up���z�8��ν��$p�
L���]��#�~^�^��9��t��<�U���1��1��-lUA���2m�}�9d�g�ffZz��z����i]3� �I�)�Z'qi�Ă'IH}�,:(#�����<�'�G
�p��	#���ڣ���11D5_*OD��5���=�x^uT�8�����&&ځ�6.��,���<H$�� !�|�����\�sx�����lc��e�-�� ����/��+ �߹��2� ���eL�ڞǷ��b;\�V�a�C������y��`꟭��Ӊ�9{e	����#z)��fd)�e����=22ݘ퍚1�ºbwfﻹ���"�x
9�TL+�Y�m�Mlޯc��{n�1;�A�������T8��c�S�SM_g�䓨������I9�`z^흒��g���� $��"H���]���}��&�>Pd��+��1,���7k���7o���a<�U�V�e�M�(�[��-OS��׹}]��3��3}��{>����1��0uf�<��Gu!jE,�[���|2�#WOu߭tO�J���H�T��I|]��]��Y�o>s�O}���ڵ' �RḒO^D%Z�۞�G�dm}SWwJ�B�,L�7jU�^���~�Ὄ]n�]��lB�vr�_F!vK9p�A�	m�Ǎ;�r�T�5�f�w����1l�	<=�@Bk��9UQ=�ߙ�ً؈�x�o<�G��3�ޫ�����K#d�9[%l�cl�i.�lY�B&Mo�����ɿ���̂\[��Φ&f%�g��ux�OD��yN]ښ��ũ�Fe	3-���y����ezH��g���0�L�F��{]ՙ���̝������Q�&rb���n�����'�3,eDS�9U��5�EF�K#��ؼ���`ش�:�F�N�l���Υ��]uP���$@�E���i4�1k�[�%��FhEJg��3ul�%�Ye���\�K��q��d�%��²`E�`�����3jФ
�4��L�1��]�Z҆yG0�,!��Pe������XK������&��j�m�����,�b$D�K� �.�]���k���j'�ku`���31�(���w�Њپ{O�2>ۭOq�����2��)�f�媛v��D�n"����%�F
l_��>�)�^w>{X��e����_\��S��n/��ެ�<8�/I�[X&;Xe���LU[,5՗Th��ΙQ ����!�Ĕ��=�s�ab��K��j�{���� ��$ҁK�����w��vA�,����a���<7mg��l�귝W�y�DdKs������������j�eN��Dz��D�B���q���+]fI�ߓ�� T�tW��N�蒺�3���<r==݋(�)�&T�wI�C���>{x� �f}"�����׹�oݥtXg�*���L���!��D�)}>����_�v���s�g��H�;Ǡ���ixIU��v��(���:�bî�GL����41lT����| 3bY�RʻBj�ʋ�Ke�8a@�ak2+r*5���� ��O�����=��yx��hf+��>͎}�&��q�����fQ�wR��uTd̡%�Y��m��_]tGg!�RM��{`v}��աjŋ� 5*)Vg�M-َ���|���O���fn���b<�3qQ���D�3�n�p�9�N�ώoܧ{���k����T�0�3R��y�ۮ��g/m�U!ց���b�ۗ���>ܻG��ͪV�h�x0�����](Ňb���8`c�}7R��(�:#E�z�Y���{� }�D$P
��Or�/z����8ź�������=� m!$	�v����DF�����g��&�ÁȬ��g�Li�2���^��]}�`�r+���bKP��#���������w�im�4��'X����w�v:Ƿ�yG��aAj�C�dsq:��7���ﴯ_�.�"`O�MT{��O���}��^]��υ8�ż;~�@�zU�Bwm��=��/�N����HBg���apsuY��F�w J��� � H���}Kg�	��VZm٘����c�Y-sU�s�*Ѳf,mؼڹ�ւ5�X&����I]��;�;+�gMfY��5и3,IK-0EVV�"F0ډr�n�Z��[cв����SG%s
�=O���Pj�e����v��,�%b�(L�13]�@&OJ�8�>�����x�Nㄅ
�t�R���j�^�*.3������F�u��TP��0(��O�
ngn�Yw�5�]̥҂<Q�A�P �dY�z�A�|�G~PA���'>�����A�<P"k���B5KǐF�A�DH#T�`�]����׻n��D�cC�����Ͽ><������z�K2�w6��P��ltG�ٙ��=|���S����]/YFfw>�H
QƘ��\}$	L��0|ri��C��;��K��uC�;���f�f�_�T�ͅq�(C�9�!�jD��T�1�Fԫ���� �#" c�2�����k�s���ˠ�{�����^�zKH'
 �Ʃz��Ó9[�}N�D��;�ߏF�]�*Pi��34�M�!i
П�����]̥��� w`:�X-���(�q�@E�Q4�X�.(h�ؗ���/.�#�A[�$�K�R�v��d��}�c5Ւ�*�x�ej4G�1��m/�O/�e�;�{�s���k_]ƈ# ��.n�] 9�"���w Y�C3�7�ފ#^-3���˹��q���N�MT^@^6}� �6��R�����#��4���������w(�'ϸ�Q�9����<��/zj�`Bp���ִ��(�C�"-��I:�3�{�O��d�4����wh�Z�
�Њ��l�{�k��von��˺�}�^� -���B�O��{�[��1�����v�{�H�޷Vp�z���c�8|�z�*��	���Pfj�f�� ��yqa�yFa`��nEcj��5��Vř�����Q��lx��!���ˉ��E���b��y�$�,�dvT��?~���c�Lm/&�z�Ft�3�fr�4A����w��w�	���>��^2G�jz���cj ��ܞɺnC)0st�ꔳ8�Y�_>�O�Uo�w3����3^/PYB� �O{�^5�7/r��=��x���џ�x��q:�n����q��F�C��$��͗�Q�1s�3��Vf���>��A�
��a�Ե3"<�̍J"��}�o�ߎ|O��̋�����*���>��~QS�r�uS+-0�Jr��%C�,JF���D�)�"�J��Ϭ���%DR�^o>��Z%&>W;���T��b���KV�v�aX^�5�ȯT<��9��*:�k&��-5/"(�1"URIE"�+T/-���Jig��zK��"ja�dH��y*�'�r��U-R�T(��1
	*T(�碻�H$�"��u^�W{�����AO�,��"���R��)�F�oQDAT�4c���^�Z� � !���hg��/P�)/Q@�U P1���g�����˹��|��Di1z��wv�T����0ϥ J����^���G�����ZO����G*�z�v^]��L���o=�O������\����a��̈���=���F?�����G/o 0����t�5� Il��	"�C��3.}ȹ�ۮ��e.��5H
2E�x13�14$�!}T���o��uf]G��]�4��{��];�]�����u�5�h<�=2����v��������,�H��&���9>�_�&�"�����e��^Y�ɷ�{�kDr�r��� �+MN�����[�ٛ(�M@�l3���0�4�D���(�%�V� G�DGnk}�yw9QÕϫ1A�F�;k�k�D] LZCQ�%3{W��C�W/��yt,�ۀ*iE�0%v�K-F�"�F�`ђ�p�5����-h� �ͧc�g�?r+�Zm��CFL@Y�H(��o��.�RC>\2�W[�~���Y����D#G�ɗd���W�Ai�6�+Ɛ���6oq�W���Q�݊,��z�٨����U��ƥ����k�7�<�2� g���m��ʗ\�j��m��`umC,։�p�X�jI�,4ڇ*�ͪ݅�WS<:1�j�ku��**�Ea^R ��4�[じ�5�Q����E�ԻH�KqR����(��#cR��˯��>��M���](70%�Eȅ�2�lWw���K-���݄�xs/�5_kw���A��^�ހ��|��y{T�Z^��0�+�r��dJ^�Of��˸����A�v���� A�B6�F5P��xz)�����W�ArQ�p � !H+Wk�[F�vWu��R�@��r����b��9�A	�(0v�F�U���Y�� ��&�ω^�=�yw�|YDAx�( <���^���{��S�7XQm�)Y`i���eg�V�f'��U!V�m�y՛t�,���\f�}������9]�e@�f4�J�g�\��kMOSl9Μ&(oh�܊�S�4�ڵZ���N6��{�$x�O����N#b���o�b���B<2�!�Ci��=��0�i�2��Ё��:{���e 4����P&�hY�qj#uBP@��UR,�Ws��ͺ�O&h�s�h�5�-R��E �R+(.j��1gv���Z#���� ���!��+����E����3IP��B/6Q�gXb$L�N�Qd{�ח��Mgs|��j'�W-�'�<P�
�<��� ܠ
�Ԗ���L�P�q|��Vm�G�x��t�v��F5z�����0�qj�� �K�� ~�ثW۳n�Ɖ��;� ��p�ɗT>��|	 � �����ՋB��9�"MA���Y�=�(爬B��~�Wo���캉K��YDb���ɾ��* ��}T��(*�Ub�|����m��ͺ�O��)/Cdg[ٛ�_4��^�ȭ���Z�lt��1AS ���� �@� (�W϶���D�>J�e�\��p�*��EQ�'�6�Ƞ ���1�}]�Q)q��"Rw�T�"�Gu"�@(���B.�L,)����:ͺ��,���
>�A� �}[�娬f�-k�0��s��áw����#�P�Sf����Mc�8�l6�*E�[c7��b����p�q�S$^�ˏ��$�D����9�iĨLbš��{��f<���y�;���%!$i�jY�><{~S翬�/�\�j�@&���␎���6�����/��U �Ž{�Y�ApA������ i���2�%?�F�!a�����4��l���[�߰�\����AxѯeԞ��y~D/��y|��������k~�ӓ[���%/#��Gx�( �*�$tmΝ��gO���qO^�Vm�\�ϻE���݁'�ТiG�}2��k�Px,�[Q]��aл�Fr-h�AP+6��!mfc����**١	_ډ���ՠl�gJ�r\b�x�I�5���ܾ�W�� $	�M�ǐ'��zZ9�
��G!��å�5������e&�=m�+ m��
���j˴p�6:��˙a�y�,	��7X�l�\��m4k-�
�PM���P�)�$�e�crT(	h�Ѝ��%r���>�~~VZ��k�\�*�$t�uf�+�	��}������_��u�6:f��$A�ED j����ϻ�p����񷝗�Arş-��Es�U�`Kiq�6A�� ��u��8�áSC�6�F�B��JQgta>�CH��>��ǜ��*�R���T'��^�h��j��A��?;���Bˀ�@�N~}��yt�� �@+�Rk�V��pjΞDC��� �R����i�vJ�͙~zˈ'J#F�z�۷/��\�C�%�=�@A�<AP Ih���-����\�^B�R߽�Nk/��Ncqh�""��D�T�E;�������H1�W��k�G��\םy���Z�Os���RB����L�1 A�@@�4QU@��;=��׮��ˠ��϶�K�R�R�G+��Usf�>��@Q���}n_aи/_ !��!�O�jIh�*����{CB��^�Sʨ��K(�5j�4V�����Jbd�2��)J�M�h�T��#A�z�� l�
��u]�9��.��҈�1�y5��n!�Z
>�R&�#%�'т��.�w�]�B>����=���Ϭ�"�"���D�*����%�����{�=:�b�r&��E�!GGQ��{�`TBʁu�����^�d	$P/�7����c�W�Y��5J? ��E��}9����0Q�M:���?Ve�\����;�,�K�}T���H#T���Nl�mV�[��: M��5P2s25�K�ݽGD	Bf$�L�&D��J�Q63�2���|;�͟	��<�;��<�����:!l�Mi{1G�G�h�f����&��;�y|��#��ہTВ8S"��گ�R]jW��O����w�_aЏ����I����ۓԽ���<r?{��Eϱ9�o_Wd�L ���^�%پ��=M�s������V��N�t�Tk������`�Y&D��� �@��x��∤�T��^���,�V M@��n���f]�>Cn ����U.f2�~��}�=�Gk�v6a�s\GL@�"J�����Z`��^���@���[u�t/�@�B�? 8� �D�E����)��>�&�/����7�>CW���DpB���'1�4P"�����ox���Ve�\�`�@�-/AT�.v$a�DV)>��b�ۮáSC��u+�(��l|dRQ�.�����Wo���7s��M����ij�a�}���}�?��J���V�}9Fs%�7Ŭ4�
v��u�B���7�����g t�߁�2=�Ν��E���x�nt �2.L!��=()���c�K˫��򑋾9K�/`���%|�^����{0�y���t㨑����R�l�gݧ����E�ʼ�͐E��X�Z�Շ6n��t���^�m�U���0���x�2D�F�kg���u����*�_��^ةJo�6w���%�������f��K���%����ХIb�+s\�4�t�n��;�>7�g�yN�3�ZνG��$e�����"���̨1�g0���~.ַEAmQPow`��pY�bn��5R��åY!�r'�O A��2cj��1z�Y-6�I�rr�r�㽇���c6�	��`Ϋ=�S��v�G��fxz��Z��;��x9\��v�7��,ɬ�C���f��|q'��B��Iʋ]5����	]F������庡�dUU�d������O>y��|+�L|�:H!���(��{��q�凢n^f'ZhV���}��W*��'\H��\��,3k�/�QL���QUL2�����W(�+�Z�
���d	&y�FҨ��J����H����X�G�(S���(oY�r��,�F��e2C�2�=���a���ԍ-�i�ysҋ�m˫�3�DQ6�RS��MrH�~���/������s�eUb�n��k3nn��3��2�ԫe��ᣂY�h�GSf�56ce�ғ%�)6::�B!tA�j��l��R��n�L�ۆ�2�4l��nܶ�J��l#�(�Q!�	�&Jk�M�������P�fr�����+�R�)�GLa�l����q�*��4��7��fN�okݣ��m��kx#�l�i��n��2��L~���غ��i�%tJ^[��ؗ4�"�.$f)� YYvZJ9�Q�DҒ�oh	t%Ļ#�ۮ��Y���6m�E�KMb��F	�n�i�6"8U�I[v�
9����ZMNv�K�G.TF�*(��V��˜*@f��m0h�4�ɶ)`�-e^tR�-�ZJ(ҵ6���\XmH7kJ Wm)�j�3D�e9��:����B˖�hQ��]ƌ�f#v҄u�Т�B�x]�S�\͙�e����&�u`�F�2�� ��Zk�[�ȹK�u5��E5`Ķ��A�9f�It�U]X��	rc��ٍ@��Q�]�n
���f�63�����hb�ZP�*������V�/]���S(A^�V�s���@�y��*�J��GZ�6�Y�f�Di6��M�IbxrY���l4��:3b��h�aA���9s���;(�2����f�t1c�XĚrg3S�5�{-�W�hJS7CR���Z�;g����~�'�/�i�gsiXc&�\��@���!{������_/�;��O[��ˠ�;K��Bk�x�.����]�Pω1T�E�i{²b�n��G�b��`n�}��:}T��E�]�[M�D}ov�ͩ�<A��PA�#:�m��l�ut�nМ���Ϋ2�.@�(��Z�Wp���"�^�E(��=�cb_�,ȍ���ޮáKA�p�����=����.��>0��c-��P,�r�\6F�Ȉ�1��8}X��^�n�}W�ja�f.g��^�>�e$.�ЀC�/��3�H#�����8�]�c�����7�ev��u�����q�Ѹ^���5�Q�!�g��џ,X�w�<��;�fT�G(�����^� ��PA4Q�����hёL(��{��t.^�@@��05P �HTݷ���٨	��HFf>��nmL/p<}�X�ߦ�}$i�B"��l��t�52��oUfL���\G�)}� �P�RF�0x"�4�����kZ 
eԚDJ3�{�a�( �+f-����\�J؅���%{O��$*�BT�e�Q���5}���[�S�x���R��z$a҈��@E �6qL���R�U�Ϸ~>��w��ԡ������6��߄�v4�s�oa3�7*����Ĝk��荒&B#�����B�'�)j��g�!��G
AJ�혿��^-�Z���0�n��AU��E���5P;�n=��An�s�꾜S�!��JO�ʛ;�N�߻�`ˤK���J�@Ѷ3a�U�2���|�n�g��ϟ:gӕ��zs"BཔH<w�n�Á}q6�v���E���_c�fDN�R��Y���e�u�й�C!+M}pD��4��� ��E��H���马Ϋs�aq>Z�T��DQ�l�e�B,�t�w��s{g��$.@�>�32y	�N�]>Qw3�t�s���h�S�fʙZ ���Uӯ�Ś�q:�0kUy焄W�`��e�EL�G2�(�j���W�M��eV����Z MrAh#EP��ʙ�J�&fH��e����jirXeg!�'�rQ�"�S}���_N)��ԣ�,�@Q��@�� �Y�i�7P�����鬉��AˁQ���O��f�Ie�V�v�4p�}��tOkx��йs��@�D������وI�����x���)�����;�E>���>��*PT��Bu&�F��ݻ�q�Y�>�!x�q7o�ɿlZ��}��d,�odx�ˠ緺�<?/ّ�����A>�&��_��܂���~��eίU�Z�W7�hh�,[3�4�e!1�R�lڶ��f���i[r��Q�nv�&�8��.5.2	t� �m-�6�[b��H�e�6��n&�m�Lbn3
miP���@��emխ�������W6AS:^�W:,m����.ظ�W� |l��( ��]1z�s��o�Ky+[i�����.�G���gκr(_�ļi!�|��_N)���QW���P,.�W�P��Q�U@�;F�Nfo8��R A�9p �>���ثRdT�^�R}Gevv�>�Z/o :ob^� �@��"иd"�Jٹ�,
�v���s��_	���yᬷ�O<{�����<k}̡��K"d�t��Z�e�a~��A>UP#��ʽ�+�ԅ�{{X�� ]� �� g�)Q��@>���H�s��8���=	��/[YlL	���ԉ�s��X5� �������H����>¿L}�n��ّ�p@�� ��DgF�:cp 42%�t�!$_�� �8�u��mkuo)J\}��j�( �6E�<�X�|��aDw%�U�f~�P$3�p�"1S�E�!��J@>�����+<-P@�r�{��Z!�! ��Ryƞ	�����2�0�mZ��ԓ��j�C��ZƐQ��z���)qպ����BO����0D �5H跳y*Hf��.�3�j����E�ѫz|��ւ:~"���BH�f �?M�aGv�q7�Q�����\B���n���?�R'U]�u3����:;�w�oו���@2$��в&"1����2�A�������6�T��<P"�3�*��%���ҭ�	�@E�������^��"u�c�=V�&���.IP�����ӧ����O���5��v�c���B%�kf�������)�>�_~�0�l_f�μ���+!�f����}PH^&�#`��;n�g�B�����J^e�̦�bL�p7~���Js���/���+(\��#�9pO���4�ɬ�5�>�����7�|���Ј�� ��~�wU�+ �[����X=�ca�y��=��;4Aڼ�,�/m4�&�
����Y=�R��*�E}Eح�o�m<���R��>��@(�S��z��Y�\�iL�a����`�l8�H��ϼp`�9�(�#9���sz�@DS�|��Äu ,���T���������C ���yO��Yxy_!i"՝tA���4�YDU@}4��7x�����1) �� j��8�@���M��A(���{�\��U����>�ȱ$N��Z^#P�p���͙��f.����v\?y{��Y��Y�.�K
`�<���V�$\������1/�s\��}*�aw��m��Mͫ;T}��	>��E�R�X��
���խp�85є�Fa롸�1��Żh!����wj��L�t����Z���Z�47 B�g$f�3��k�-Vii�,5,�%��&D�:�Җ�sPy)%p��7=�ۣ�5~��_�o�[n�L�Й �;%�LD��������y��D(��|�{.bR�%Lh��>!�k^�ED#T�JM54��"調����{����U�y�Ϭ�7*>:Q�@�  0��&b�Q��ٚ��/>m�p4P ����a3EB�Y�vВ0��]�o}�.�bR$p<Q�R�"(@9N���a���13�GH��8���5�Y �Ǐ���A}DV<[���>���3yك�L�s�ģB�T�QT2 (��T��(�����V^�/�b�}�|ER����x���A��E���Ut�J#�O�.H^Z� ��k�V�	�n�>q{+>�I$�޾�O���~���~O]�	K�'� �A�]Ņ�LP�E(/e�K�`�pEC��:Ƚ�:���n�
��iz�zUgmɺAA��&r�S��������f
|���f@(l�ER�J�Y�v�Ws2��Pa�/@4~y��?�z��X��+S2W�ё��\�;5Zm��%��2��;��<��	뮽�� 8⺜zc����iz�G�'cv^�-�A�3�9η�/�	�@ih��#dF!�P� �.ЀE$� |,Y�FX_�yc }�;ia���<��7�����m�Ӓ"#VH�[t1�R]l{/JuS����Z;vGvŲ���Wl���c��{g��:��m/�I<��\�t�<�w��&��>��]8q�l�V(�N�q0�k��לL��$F�e�U�z�	l�>�1�)�P [߫"l�۠�;W
��й{�{!���q�˃}�����{�&�
`ΰOipl�|�m���~�0�}�$:kX��7�Ы��C뛯=���<<bm�W������iN�M��#�&Hx��,��y�9���{bK$7i���璲S��X��!��ݫjj[�;B��1��Z2�SA�\�������<tt�DC����;����3��Po��r5��?o\x������c^Y��ߗP�����>X��|�ݟ�끵����f�Į��K�hdZ��1��'sq!���?Uhf��Kʺ6�es4QOC�[�~��q�%���u���#�<b��y�z��}��{��2�
�7QB����"K����W䨗�Z��S�ʭ\����j��}��z��������j��I�QW�,�� �T/)]L<�
""$�3�&��G��B5r��@�	��C-M
��uK�¨)E�jQy�9GS�ܭH�˪�U\�\�2*���h{��h�)xQyTT�nAfeQ�Ж�cr�f֣&X�t�!����$���Sʯb���H$���m�����K���� �R�*�;j2Ђ��5P&�]66:���3��ޭ�+�y���S�(��ZbP ��-�Ӕ�ԋ0W��X��V^�{��A��>�@\�QǻM8TD��4�G]*���Eq&b��"P4%��= �>^�ާ�Ϻ��e.�#���c�D���P �@�!��t��
���2���:��	en�G����$�h"��(�H#T�Q����V��������'� �Ex��"��ʱ}�{�A�\xd�x�oV���Ws2���D]��V��ߦ�P�PQ�U�v�=�=�w�P�nmm��26��)�כ���������T�4Q�EM}��02 @��_�XqאI#�>�@U/@�:/�-뻓}_�O�<⎰�]�m��s],Y���m���|!���5���w]�������gzX���B�#�ǁ�$(�4Q{ч��tΆ��"�{����fR�}��@�.mY; *��{u �^�誀�s�o�:k������g�]@dY�Zݨ �2��9�:�;��Y���}O�����܄�����<�̟!� Q�L�4��y��P|�ͺ���Ws2�	��
�$h�P����r�e�bz��0�>󉑯Nn�J#��fD���	0r�=��~�N�N�u�Ś�͙Re]��fl;���ɣH�h�\h��@̴�Cij`�g�bQ���Yi��6J4�%6/Y�l`�
�{�ҳK��k�4ʔְf�FXm	du.��`�߻>+<f����|�~F쫈S5�6L=f�0M��V&L�����G혞�M�U!9WU�Þ��x �w��>��������#-x�IHÈ&h`���ާ՗�p^�Zd�G�M���"�s�u=�a��B���#�o�Ӵ��e�<���fR��,^�^�h�(����@��A�҈"�eM�kf{26xQ�:�ɼ��"M%�4P�,�7k��Z��=ε�^�I�>�`�UV��A\%&LʔTyI4�-	�d,��ً��}�/ID���
AfS���]���>"(u̧p�>�R��B� :�Cx�7�MQoo��K����w��{����γ�ȳ"(M*��?ǀ����x�NuM��f~̀yy�FREa�[��0ίP8Qת��QDD�X碢���+�e�Dg.� �@�D�E�����D���*A���o��&R�>���;B��P}e��G���^@ў?[Ϫ�8B����ٞ̀H���HA|�Y����|~�~=q����s]%��m����}�y)=��J�̻��[՗�پ
N��ܠ(�:}T��@�����)�@i��7Y��뻉����1z�o�X��*��^�B�4P ��GIk�yA�DT�����Oq���a:�P�^��N��;��;�{��4�̐O��FW�Ϭ���jH�ff��9�����o՗�r�!4;��L�9��	���^�*��8��Y�Hw;��޻��K�'H@���JAGlٷc��2��DJ&tAHV�,��Ll���&p.��b9h�U@ꋞ��]� ��FoT�A��b^��ZR �^#N^���z�i����+~�V^�@���!�~�z�;��A�	�$9���V�12��=뻇U��>���4x� �VR-n� ��#�ʪ�_W=�ْ	YG�cN�p;8��
�#ؘ�"��T"�n>����|���Q���_n�{Ny��C�k��؂�*�$%i�I���iYw8���^�܄����}^+�w��a�HH�Q+�̬p�;V(�\�\Kg��cb�=����������&R�FmNyub�8A㖠Q@�!T�&U��P�g׈Hu6�6�fH< ���P;k	5��D�\�]� �=�2�=N5��R��moV^|������?�C1@\a�(�>T�}Y�|�]�L��i��Om�,�5zG�@h��?GfZ�u�E������4�2A>����z���h���2�OFչV�@<��t�t{���%�>d }I�w�0L�xD;@EP�=��eD��<�x����2��KR�\4
��lV2�J�fF\�V3`����@\f�hǜ��`��#c�ƍ�6-[1f�P���B[�[Y�f2�k���IMo$]��f1�#��v�a�����~T
�0r�MA�Vn�+�����w�~�=��x�� L��wS�����Y@�hqB,��EW���U��(�F�Խ�,�����jD�0~������@�ܢ���^�@E/Q�U@y��e��˳(��)	"������k�Al�A��$�������}yx{��"��Jm! �Az����EA�^�A^n�s}wq2�OF�R��8�TL���'�.΅����Y�]�H�Fص�l&���Ma�#؂4P"�!Sy��]�@��32P�F*^�@Q��֘s��t�TXT�ިu���d�i�-ʡV��Ν8�a'%��\Y�R�*f�m�u]XMy� yh�yY��m�"H� �D�E%�H9�J{�fw]�̥��! F��Q��>�*rfm
Y�@�U�76���t/2�"���C���z<h�%
�E,��C�!�Ooz����@��#�H#Ej�G9���Z�!L	2dHP$�T�-	�s3\�W��u4�G�Ez/3�>뻙���,��nC^�^��DQ� /��FM+�d�M@���y�k��'J��Ɋ���h#x���4�5J��ѻ5DH&��B�'�o߄�<'�)p��0�g��Op�D����K��^���s+]��\'� ��ET"�q����>�p �>@�
3s�>뻙��g�>��|Lذv�g�R@�� "�F�%
u��C+�os�]W@�^�����={�����}��03Y]��V9������b��,�N�O�ǋ?�U_g_7^^��Q3[]haJ�D���������a�jٝݼ��fR�	���$ݡwBLO�j��$�k�`�*�v�NTs���-:���P�) �iz�I��>�*���3v��^^�� ��=rط�3T���2���h�f��7��&n	ݴ�x`�P�7��څRj������z��Ϸ�u���^��F �R�#�ܪ��}ޥ��:0RՔK��-�7h�&���{>z�{#ǂ���M��73�]7@�B��o��d�� a���R�}Ef�Ι��wTN�����}yx{�ר�V�34&* �@�#��E�Y	ͨ��Zﳜ���\+ǾPAs,�B�����"Ђ,�t�
���ng4�jA#�D^]�*�i��FJ�r�E��ZA�FE^W��K�׵ח�r�#��IH �Pݑ
�ƆX�r�g�n�M8rV1=�dAyEbY���b=r�}p�+x,��cM�v��0�*�w#D:0:=ź�Ս|��
�N���`�_f�I��;�Oi+�-�icrs�3��e����|燶s�pwf���ׁs�8�������{a��)��^~���d���l��R576�1�0)yb�ؑ�JL�+S�ӱY ��ܩXuSW��A��e��n�6,�1�\:���2�H����k�}B�=�����Т�[�>�&=��u��4_�<�;��wBd�����qÚw|i���<> �7Ն0onx\�@P�C\��=���v�Z걄n]8U
D�]��nF�;0����:��ꩍ��<4�;���[w�	x�����`=�p�������t;|�wz�н�0hhq��W����&=#[�N#�O$���ߧ�q���~3H8�<D�cю�6��j�$,�����z��?K����7�Ģ5"������t�Q�D���M�ÿ?{�~=�}�J��R5�h^�r*�KÐ����
�#�j�}��?R�p�*�s'�j�����Wls��}����`�͜�Oa��ؼ�<�.Ɋn�lQSS9�B-�o>�ߕ�_O��vHX�%,XbL�8噥�����O3sD���(�t�/'��KP�(�Vֳ���^!z��M�0��/���J*�����/k9QEEDU�Mv��[�|Z�^��UW��i��D�H�ƺ%#�*�̋u$�U^^cȜ�2���[�ah`�^���|���پh��m�P°GK��6��U`�x[����NR�`�֊�v�uD����*��9��QSM�-��lp��(f�XYrDN\����8׫��s1�e�v@!-�0��T�v�z����qv-Xm�]���L�3����.AeD���	3rU�܍��R=nu�"Y�\̚2�bi���ɋJ���vȶ�Y\�B���u�T͡�1γ@9���a56�`�R�+�rZ[��A.���c\	M�t �#�)-K.77bmb�v�QK�I��]X�0v�]�Z���*2A��U�ʷ`1cV�0��
�ka�Gk���D���oJ��FP���V5�c^�э)�J�J�1*fˍ�X�6��Pз2�Ҥթ4IsvxK,��9��/;W�5�%�H �R�d��K����4�k�G\+MDƌh0ʃ�궍^�5��Sۈ��-o7\6;٘L��з)k їW�ZcJ��үh��WMH�.�V+lUa��l��U�+�UW�aG\�3�W��z���n�b�P�e�S!���[��W;ˁ\�M�0.UUU�l��t�&P�\���f�Y�>4zo3�T<Ķh�[������[��T�h*�lf�q�P� K6�׶�W6˫�-h�֗��J0���K��DԵ��iR���@�l!k+���1@a��c���-�̢�lʛ��>|��K�2�2�4�&׌��H� �D�@�����h<E�}�g�ڑ-'�3�m��A�3�*t`rB����](ig�#�}���sK��8P#-so+X�h��Ԃ	¼EU)>�7����ʗZ�;��.@�܀g�h��J[�h����v�}��wS	q�e�S��80!p�v��q��p=�"�����]�$q�������1�s`��z%�V��Pcpu!첲bP��i�|p��0}eL����_^^��1�Y}F�@�G�}P������٘�vrÕN3��ChA%��a����k3�w�UB:� C>CP�yϹ������}W���Ս,���Ȑc���0ER�./�ij���K��^* ��>�^j72; �P@� ��F&�����%����}�Ae
Af�D��]�D\��`����v����K�'� ��e�Ǯ֗�>�+A_� ��]`F:6�L���;i��	a��y=������ݺtϭ��^�R}P�G���^�^����κ��.@��@!��U]B�|E�G
"�R��~4��ɯ����A�g^W`~��@��5��D�����M����0���ٷz���B\A���R��Q4�V�ZE�Y�Tq���+�L��L���}J�
q�"R�>��~�
�y�o�u��G����}�p�[��F��	0`HQ5�f���t�t��~C�G��A� v��Q���tu�D%�Z��A7�j���k�n�g�h
!�ܛ�7�:;p#!��m,�+�p�3}�wж�-�3���4�mn�x�nЖ�{*���������G���7�@6|��Ah}9P|�]�zȏ�9��;��K����w@z�V�j��Q'���b�˿3&�8��_�7d^�������%B8o)z9w���Z�ݡ]�2��6k�k#�D%�>���� �u`b��J�*`ʓ(�(�Qsf@G���b�<��|�|ȓv��Q6�<�w��r-eGa��0����^��#A�2q¯����<u[�w�Wp���#v���W_�U�����e��J��퉺���"G���E�G������ɳn� �A�ډ����^}�"W�Te�X�ϷP�����(�� ������þ$8�yϹu]�K���C�!�&�Rk��ͺT9��7�}��;;���֎=��U|G��8�ک��P�D>(�0�A��BF�A�X�D.��ZW\7u�v�u��&���$��ڱso�R�j�X�,#M�ͦnÓ4��n��Jh�6�!Ք���(�9n�e59ű��-0McfmTÔt��-���=�6�.����VQ�a��jۅ!6�Ϩ���w�|�8G�u�}��VG�"�&V!� �O�����k��t:?^;�I�}�]{x_/΁6T�N�{Q�(n�Ak�hg&����|��uw	.�����jH&�A���ڜ��H"�z̑v��y��":�B�>���[ee�]Ǵ��*�Z�����%x��z볩���� ���A�,�hu|`��f��?���"d�� ��2K�WIf�b��eb�?^����{ ]�U���=���v�!q�=|�sn�� ��@]�"�Z|��q��*��@�4�ߓ��==�{�\����˪bg5����O��`@�痭����8}���B%�\n�HF�J�'qAF�v�Z�6��7�n��";��A�A��hF!��*�=�ܩG4��hF�v�4��\�򏗾&g��{�q�+�1��f8\]�2Pi�W=��	/p8Q�Ak�D~�'� �~,V��7Pa�	���vX�q3��,�|=�_^��ݨ��w��o����.B�n�g���g�\��;뺕��^�'g-��]Yp�5w���W����A���!�"�z̑v��$�Lճ�RxEݡb�_n	ǟ>��6��9����k�`��|�n{�rzjHq�>1�́��]�Mu�����;�&�]fu}�n��Di-"���͙��� �h@"�= �gȃw�.	yW��":���r�ˋ��>֠�}v���E�h��ߟ'�J{�
�dI���魃!��2عY�偽Y>{��N�w[�{��PA�ut%|}��G����A;�je��jti�� ����k�}N�.ϐ�A���sx��BL�1ȏI@�.�����4��uϓ��I��CAxݠ ݨ"�BL�o`�#2(v�8ۧ��t��O��oh8�;��1/d�ԣ�����r�
ŷ�오Ԣ�m���vk�E���k��Av���Ben���o��:���O�HQ�G!8��\�Ϻ}�ڷq��p�ҵB��h�fjd̮�/�>��HN���� ��7���˄�:`�>^��/�k� �������F'�#�A��F��=o+�	*#���#f�"����� ݯ@7i�Ur"**�9O��:��í#y8Q�p ��'y\� ����^�Al��˧.\A:���uכV�^����A����6SW��ͼ��K�{J#1�3" 8���76lV��'J�:Dg�,D��3�2���̇9��ب73��0�(!�Հqqu�c`X[���M)Ef��PIl)�0��J�Y�`GVk��Rfk�1��I��(L�kYt�u�.[,L@��SZh�c���̫-0MR���u6\�篓�ֱ�f��E͙��Wku��O^o�C��'�jӗ���hG�P�J_!�O@���"�v��e�G�ӓS�O^"�����u�����m{���ڕ0��5\!�'i"�6PM�MJ���u� �t�f@k�Gv���He���@���T'1et?��r�hDp;�-�)�Z]���]��.׬�"�"�
�[u�H���w�(�&�G�֠��@ՠ.� �Ǻ��K����-@k`4G��[?/�O_A&�Y�7D����iel�dfn�m9��2�/�<����[��M���a��T�|��d��!��u�;Es�}M�u�����`Dp;�hQ����Zp ��>(>�@f/Q��7�|�Q�i%����D�� �v�g���!�݁��C!�+���jv{�E�	/i�;.�IQ/H�*�G�G1Q� ��#v���^:��'6{e��0G�@ ��"�[F�M�M�=|�����	��ifM�^���Q"D�@��5?G�����"�*�����\ݷP�'2Ց$"���DY�ߌ�N�%�3^�^ ��2)����!.�Ae��ws��s�����BJuQ��z-z�zM����۾����6SK�FJ}�W��w�C�Յ��[7� �@iN�z��73�'jl��z*xϳՁ��ޙކ��Uk�y��՟E�^����;��g���AZ֟?M>��ǯ���^�^����ɩJ.�tn��f��b0664mC�:�B�j�mۋN��i� �o3F���ϳ���qĶ� ����w�Ywr�cKӷZ������w���6Wzc`e�3}����v54a���ʚ���0����!���"��m$�R�+`�C=]H�s�ޚ8�U�jѻ�Vk�d�m"�c
v��Ҡ���;��� Έp�˃��Y4���9N�ȋ;u)�/&fY�Oa��e�5��LdD�3p$9/Ϊ�l���Ǣ���fMW�[.�9/������t�{�Y�I彉-ՅcUn_��;5`d�N���[P0�P����$���B
�-T��R%K�=�߻�g닰�0�yhK�1���{���/<a![�~�ߞNS�ګ�^3*/f뾌�JcԱ�}���D�%(*�|ǝK/G���P��+�Z���>D���E��xL�UT��+�b�q��DQT���Eʬ�L
>^iK�sQ�R��H)�+��KU�로� QDy*U/Jכ�<��{L���8A_R�4-)
+Ƞ��3�*"���&dh�^�=�9��£�׫�����+���|�o@�/�g�]�hU�gq
�h�hAנZ�y�������,Pm߫UMj��as�ȀY��u��nt]���?� f/a�뛺ſ
5����"BFb�L*:��JE��a�����}�Ы��J� �ڋ���g�8��ɠ��\�4���hX"�l�)Қȱ ���C��;��=����j<||��;�;�:��}܀������~싧��E�<Y��U@�����.E����~���Yq6&�fgL��W��*"��n�8mN>��-tڮ�yv�Z�{-��&��΅�g���l6��ˁq�g��t��j��s��e���qJ�HH$35	���f �(��W�����[0�������qw��-�L=mb�Rool������������2R��M��4��T�U
Y�׻�>�#���������vĮ�n{��ld|<����v�*���S���i��͵���������DU^f=�s4q��Dd�XW�0V�N�T"1^[&<Hv��~��=�~���i�J��|>x���h,���
�#�X��[1a���k��֩�$L-Ƌ�+Pfg���a�ݳ��Hat]�A��4�и&b4��`
�31�*��i��!�4	�P���]�;�R�\�^��|u��E�v�`s4��]3u�����z�ߢy���u�ߺ	�7Η���U����Ϫ�udN�\x�����H����U}�%�_	����T* �M�g���1ۭ���U�UUN��p�.���j�u��xo�}�S�\���y}�M�nHc�$��F���z.��FeT����yuͲa1kYtd�[�j� #5(��J��]�uQ�*_s0���,N�~ͦ����2/������(�*R�瞵�q$�z�����G����5��d���Q���֙[f���"��v�v��}?z�KSgٽ�.��fE����92Q�{��9B�jq�a�sG�\��t���d�x�6����D��Yӻ9Fv#�kA�@O���Ix�L�DW�rTn�D4�]\�΄�������F�g=މ�xJ9"b�����+�H]i�m��S��P�����U�
��|�dt٪�����
*��%����B��Z�g�ydQM��]�����;�c�r�L�#���'w-�ǒ��;}H��66X�q�D��Ƞ��o>�m�{����+ud��H
�*�u�î�&v=ڮj�Q�����!yP*�|�����O���Ά��ٺ#���ËwsN�)bչ��=ᗋa�"�}�Nv#ÉڱN�וSFϮ��͸��~�׸Chî�}�&�|.ЪP�`�QΛ�uUX&6rw4��Q|����W�d]�۳�u�>�:��ǭV}���\�]�=Ě��z/�󚫹��-�BU>!>�&w��!/������g,~��R��H{����}�&�}�*��,����_���P4vS)G,#%Y
d��11(DM�\�UTgs[=���gW�o�?�q�9��I��d1��ҼϷ�y؏{Z�dUl.���(�3>�B�Q��֑wyj��o54�{�ڪB���*&��
'⪩׼�{[��ƩeNX̸�B������
���ٻ���_>^�U�J��f�����oٌ�u�fؠÙҸQ%�7:�3i��r���-�ڑ|B�ԙ6)�V:!���=��*VཋaQ�e�Eִu�V�1���٬�a^�X3Z�*͕�4Wa�:^Te`pZ��#-�,�VԻJ�v�I[�� k��#vs�h�B��{�>��k�@��j1	f�@��gg�����՞	��<�w;���G�����XQuv!F��z�V�D��bU<��OkpxNtz�e��5�j�5Ōce�����^���}�Y�q�z�6�#��W}r:~��p�`
�s��ڊG�"О�������*��9dݫ���'�8=����"����}�꿡܋��RcF��t�c{#k�j�E5aԃ�'�m��޿~�*g��χZ��qg�n����u�_dQW3$t�+��!�_1[�n�2f���s�ݝ9&�r��(�Ӳ#r�ow5�3�*�'/E���m
��*�:�����%�p{��
�(����7Y�t�+#oo1�W����r���V�UU���s�_|�\m��ʯ���$��wwB�8WY�Wn��2Qu�2k��5f�J;"�%2k���HT���|�������B�T�Q�tքYu��n�;y^v#ͺ�x�3���������SP�w�t���\^��$�|Od>��{7{6e1p���Bo%eu�}������z��@}���q��Dq�p��:�ƽ��)��>��j�;F�ݺUK�G����_��gi�G/w��R/_q����o'�s�����<j]4�s`"j\f3 ��"��tU�^�7$����3~:���U,B3�PmT����|����sG��vgQN��2R���٘�o�U�b<^t��R�*�F
�G�fd��ϱ��8�'��2_0��X*Q�9�f߭�61����~{ak�"��B��̀�ՙ1�w!Du��f��pY����Y�����>UhQ�����*�XQ2���ȅ(�"j�C\�GCi���o��{��燜��;��G��Tx�~쨪ok1U�����ӗ{��&uu�Ϲ����}�U����d���"�U���Ö�]����
�G�J��(挫X��Cyw��fu�͠v��hZ�My��R�v�E�Ub�Z����DR/��e���7����?�?���L@v�?�]�?�A2������T	j(�Ԋ ~_�',0T@�^���!���l`.ر��ctd��&k��v߮�8ɋ�vX셂G1[�(Z((B�(B$��Pł� �
@P�( A*(�2��@��F�X !�����Ш"�AAPDAPA�T=�APD���DRAy@DAAAPD9���d�Wņ`����h8��Z$�U�(Z�-ZJO���[�PEAD�J�IQ5�����W�g���ߴJC����2�BΗ�4�����.%�#ή��@�4k��UD�D�Ԑ��&��C��É��1�c���"��O?��:~W�@��Ah]�}"�"�t!*?��"������c��z����b'�������g�����{O�~�A��>�YG���T��~e?e���\>`�����'��d?PE5uSG��&&�#D����T�"ļO���pO�����:/h���U�Ɛ c�}� ��Hu^���d���V��a�X�'v(���LvX��!i���@P.�Y�/`	/��J /�j Az�	ZlP`<(�R�`����xcq=��=<�`��Q@D@)J�$(��@R�P
@���c��z�Op?#�g����`����hF��~�������H�>�c�{T�!�}v+/���p�O�@�����*գ��W�����`�����Z=�C�5���2}X?G�OY��2\(��z}�X��ﺗ˱O�}%w��M>��>L����'�A?�>���pO�=acց�:?�>��������"�q�:���`e���?�����`6!�����(#T���AU,0����p}c��"v3'�|!L�'�������z�f�N�I`R�P? tz��" dr��� H�"�5`��B���a�%"�����`{l�>�t�vr�xL�(�U���!�[����E�����	�h�����(�'a�K�ѕAX=���c�.Y����9�����Y��a`s��gB�/c@\�?����=�����_������d����>a.
|O�>e�/@O�r,O��\
�z��N(�j�z�-ϭ,�����������?yH�*��>�g�{��@��D�h@�?���܈"�R?,��m�������=���?`}�� ���}��=���]����ā�� ~Qv�,w�>s��\(� ��� Q����)���)�N�g�L�߬�����s��=. �� ��c���|��΂^��K��z�]?9��D: }�
!?hp=�<�xH>|hl@�I���G������?)�����{b0Q@��b�l��,����)�!�_��O{�ߡ�{EDr���>�=�C��'��C��9f��:bݾ�	�����I~4��H�� ����z:�.�p� �[7�