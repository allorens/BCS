BZh91AY&SY^~u��`_�`qc���"� ����bD��          ��R���HUB ��j%
ڵB��J��T) �
��)D�����A�ThVH��JR*�-!�  �ov���VĊ �	)U"H�T�*�PP�ld
��$l0TTU�T�2J��Q%UT���Mi
mf� ��
B��W �@��t�������%p�ԆFBJ��D*�iR���%UP��Zd�6dT*-j��R�
T�QY�t 0�хD�  8    !�J���kK`�Mf�U�
 `کTb1(��T�T����i���֦�����Dm֫��)J��UIURU�  < ��GiV�(+l4��
3P�P�3V���T��� (*� P��& h�
1� �6�j{�� I 	�m�%R��x  bx
Pv��UAG4��N@PmWwT\�z�ON
��� �N�U(��5H5Ӆ �oks�t:tj�m��H )@��  1x���;�  ;IӔ�(���Pv�pA@87q�@p���
���.���P��P ��+��ڢ�����MB���x  d<(P��B�Pʺ�ښ�Wp�R��'G��y{� *��p5�Jw����0U�L��P��%/l*�(P�x  m� �� �9B�B��` �1�B�d*4��F��� �JM+U� Ƙ���.I�@I@$I� m�J��  :�zZij � ��� �0 (�V 4
��Ř�`  �MBR��*D"�H
�g�  k�P�`(UTiP �0�#S *��0P46��Bh�,  �IH)${	J*��  q�(3 4����(�L �  �X
�� ݃�h4�� ֆaP�%��UT)U^  3p
!�T �p u]��@a� �` 	�  7�r�@��P�N�p 4�        S eJU!�L` 2bOh�JR���4��`�F&��0	�2 	�`  5< TԥTbi� FFC	��T��4�A���     JJ�
~�Oh&CS&ji�z���G�}��!�%�J�L|/��|G�c�r=m���{���g���{�󿠢 ��~z���"�
��T��"��@�h'���_��S�Ȉ��U�@P_�T�\ ����G��_O�e�[��3�d1��<d���'2q�a�a�`�M`�MgZgY5�Y5�X5�X5�X5��d�d�M`�M`�`�&5�Y5�X5�X5�Xu�Za�a�Ma�d�l`�L`�M`�M`�a�&5�X5�Y5�Y5�X5�Y�Xu�Y5�X5�X5�Y֘u�Y5�Y5�X5�md��d�M`�d�Ma�c�`�`�M`�M`֙5�X5�X5�Xu�X�u�5�Y5�Y5�d�f5�Y5�Xu�X5�Y5�X��d�]d�d�Md�5�X5�X5�X5�X5�X5�cX1�X5�Y5�X5�X5�X5�u�Y�d�u�X5�X5�md�Ma�u�md�d�5��d�d�d�MgX5�X5�X1�Y5�Xu�Xu�X5�gY1�Xu�Y5�Y5�Y5��Xq�Y5�Xu�Y1�a�Yu�q�aSYP�FeGXU�Q5�M`XT�u�MeSYXdSY�U5�MeX�@u�`SXSYRdXA�Tu�M`XT�5�`CX@1�`X�u�MeYT�E&u�M`SX�E5�MaSX�Tu�5�fE5�M`SX�Au�d �U&5�MaY�5�M`SY�5�MdgYD�5�`X�E5�MdXP�5��5�LaSYP�5�MaYP�5�MdaeC�Q5�MaX�5�MdYD�CYT�Q5�MaSX�5�MdYD��P�1�MdSXD�5�MeX�Q5�1�5�LeXT�E5�eX�5�M`LaaGU� u�aSXT�u�M`��E�GY�u�dX��WYQ�dP�DX1��C@5�CY5�XI�SX5�X@5�X@5�ed �Uu�]e �d�XE�U�PeX@5�u�T�PeT�`�a�@aU�]`CY&I�CYP5�YP5��5�X@5�Y@5�XA�U�5�]a �5�Y�YP5�5�Y�]`@� a �Dd �u�a�Yu�Yd�`q��Xu�Ze�Yu�Xu�Xtd5�Yu�Yu�X5�e�Yu�Yu�X�I�Yu�Yu�YcXd5�Yu��Me��e�Xu��]e�u�d5�Yu�Yu��]a��1��d5�Ye�d5��a��\e�Xa�]e����CXu��e�u�e�]`5�Xa�5��XMa5�X&u�Xa�Yu�d�u��]e�]`�u�u��Yu��pa�]`5�X`'\]d5��d���&�J!˘��W�詝�����.n�SRz���|�;-/�P����K&��s�8�s�.mef��8�Ѱ��,8mG����������]��4M�Q�4��B�xD[sn���a=��x�	A��K��̹5ł-5�	�D�l�E if��j��O2�뭶���h���gtS܆�n��4D���Uy���d�d 5?�Sm�[�Y�� ���`�5�ǌ%��Ii�ŌЦu�Y!#�(��0�Wxub��V�D�롢l�ȪƚhfU�!���/5Ӧθ�扸V�U���J��.�筡 �!���c�xәY�nV�	V:�"��aD�v�Y�j�%4�Q�2�X1=��/�=B�ݼ-h�T:S�n̂S�j%�p�թ�:�N0�9�(��9BS��R��cǡi�Sߍ8���$1Cp ��qn�$��5��Y�I�1�FX�FT�kO��V1�d�v&�@��KZq�+
�o^�������iYw�u�����i�a� ^
�m=H�oa�Ћ�M��+1چ�Ud��2򭀊F�7g.*�uO/,�U���2�G1d��'�X�u��V�4nl��� ʰjGL�zEXT�㲃�^�/��6���x�е�Y�2��X�����n�CS
����t�Od-���*�-,`63S��]�3h���%�j1x�������c�28ik���h�O`��w�z(�on稃,A��.�wm��S��&�C���5��(�Y�����3jn���Z2��7o��խ��d��Q\��[f�*�r���&S����0��:*�6���c��%��t�"��Q9N-��▤��x�U[L�6N��Y�������BK��SN� :ڷN�������ܳh5�&D�@q�E������B�ӬZ��K�-�k��*��K9n�ͭ'n�[A�iZ֍j�!,�G-^C��(�"馭�ɹ���i�z�@ZN#�ђ,F�غ5l,x�a�A}bU�
dڷBYن� �L��:l�@�*�14�Zj�H�j�y����#AC����M��d�~�)�*��4�ܱv��)�(e��#�AeEUW�:�;e��[�*H�̀n�lYO$��7mP�LQqHP&*[I����t�U.K�] ӢrLʨ��d�m�)W�Yz���CB�2�	�nTFKzD[D�h�Բ����շ,�d:�>Q�tK����1�JA��	/u<#˺9�eL��l8�0&�L�7�9�A�b��]�Y7fDm]9����P�0\�Z��hZV��t�*�͸�6]�+�v��MYzv��$,�Z�v���,.Z���j�Y���X�j����0m�Y6��t���"�Kp���E��p�b۽7+`b��K��h�\P5V,���;&���Mn%��i�xQ��r���5`�^R�[�[�ܥ�Oq�q���ǅiɔ"sh��ԫ^�T'(ٰ��g]U����;ga��2�Jz�+)R.��'`��U�_Z%R�-��f��ʴMk)�*T��!��mؕB�Ȏ�Zj"i��r�r�zc���mwKS��@��h�-Mv�{V���!��T���<�%ư$fT���'I��Ԑ�!�U�);��l��z[.3e�2�wuAk�XH}P�cvW!%�ڑnQnf�:�a?��
1=X�ɛ
*�"��'&��^�+F˗��X1Y.=Q�c-���7�rHijt�y�!Y��e�l��B4���#Mo�0��uLĨ�˖�"惧4h͕�r�;Ad��C��H)�e����P4����#�r���7+X�!�jn��&��y-�ߚ�lUe�"<,�n�i�2�{4���=d-�+*亹���Im����ޤ�bo76��H!,&�t�p�%)ݛ��4H�����V�&弘i�Ĝ)�(T��r��T6@7�ҧu�+M�b�uae����h���h�8���/�n��4��Lv�c��;R�pV+(fF� �h�٤R93+�([�A.�`D�JjF�Y3M�*Ѹ5��뭶E�9n��6�<z��I�)�5���"6&kh5�vXί*��Wм�ې!w-�&l'��������^R��b7
����"m��^�jl�4Lf�*,�wnLEXcFTMЂc2MT�V�Y�7�i�sn4�*�V��̋%���$Y�$�h���	����v�(A���'���li˺l�b����]*���wt�Ɋ�)3UKkj�!��/K��k\R��q�[nm���/l�������ҵW�&$a�]���ۙ,Z�7X�eAG ��b�T�QÔ�]��N���W[����d�͍��=ʂ#s0emj".��#��5�p���:d�U�u��(쬺2��L��`��^jS�e��f�Z����{�I��\�$Xlm�Ec�]�(���i$�U��*�n�u:Xʺ�NY������.����K�i4ZJ���E���1��cWz���c���mw���3e`�ʏ�nu���VIj�����k���dV�i��]�z��{`i�kudO[�	V�W��}(���h<�OZ��z�U���r�� �1�V+
���n�����*�`���uAVT�te�~4�Alٶ�y!gF[YR����Tѱ�+�޾�V^a�z��v�*�e[a�2r�l��*µ��6I���"���-,�T!��;��%��-Z�R��j�*Z�{s����@r�6��&����V]aef#��
�)Z/%[�bIݱQ�$��VO��@�On��3t�Jj.�Z������V��TH�Ϯ��ӡ"˨N�YCu��P��cq��4�^�4�Iaش;M��Ff0�U��al˚�]X-�9�iPN©vU�������S��w{hKn`tf�xa��V�X�4�Gd�&
��i-bڻAՆX�܌m
8)�
T�)И�#�19EԔ,dͭ8��{w�M=��Za�lb�dJ�w�㔠���F�a�Oq3�
)1D�ݡkV�,�M�5��򡭍�&�56��ܠ�Cx&\����]	I���A�F�JZ7"tMAa]<B���+S{Dk��5T�n�w#4-ܭ�ݽM�{%�MC4V+�,uyt�@�q=1L�zYf�o
]O��o�/ۛB�:����r�-����zl�v�`�Bʂ������Q�RbH����� �F��l�&`߅�̵9��(53��I�݇l��<dB �wP�Z�'J{/j7/�d�Q-�"3p�X�+��b�R�YVhm�wl��:�m�v$�L;W��z����[{��L־��6+F����Ld�TklVh�i�D�e)C�(l����h�Nw���d��`X"ݥ��6),����P�or��w{.��e�G6ل
6մ��Tdlv(���g,7�������F#@����>`�՜<�I?�p6p�[�%lJyLE7p�MF�
sV^8s�+֠���+�ȘT�LGr�v,��q��"�9�$K�V	�� �A����t�k[�$YZj;�ke�(�Gb#m:�Q=d��1�O�ݬ�rK�u.�תf���	p�iX�w{�C�=;�Óv&��`9���3)!�u�j��Ԃ�$K�)����úӷ�������}��i|{Hr��,�u��&2�[J�Sj��IR�7 ����h��.�S@�w����tu�v�0��E�d�!%���dF�W.��%��
��V��µ)BA@,�,L
�A%�E�����-Мw�˥-PҢ���n+���e������2�7`�g,��Ci`b�+�r�_�	��� ���I�c�.��R�`��y{SmU��.�%��%�m*x�k�ǲ�[�f�V���a�P�
�+t�DИܧ�Y��'rAh������a���w<wbU���CXѷ���vu�qM��h�׳a�3M+�t���S����@���&��8����Ѭ;D]��m9f	�ne7x݋āy&��3E�y��x.�ٷR���7S�j��f�3H�уH��goFm�Y�Zn�G7��*���ZYi:^O�eՁ�H|���4���������w��%j�L�u#��)�4C�<�z"�5�6��u.�4���,����.CW�O��6� Lt #(��`�J"�#N�~��Svf�a*��Vf=.����7[ݒ�э�ǥ8����S�D���{���/S��W�cl�T�i蒦བlH�*� ��[X԰�n��A�1�*�9����V����Gx}�.hM a�[�e�Ȧ���4��e��Sbe<����3Q��5yB���Ъ5�4��E�F[����4hܲ�ص��e�1]�fɗ{BVK���.m-ٹ�f#X��i������HZ��k�6�%.��`<���� �p-ɀC2���Ӓ���2���T��v�E����n�LN$�Adcŀ�z�f\}�r�Ƭ5)jSq�z��7E�*n��T�GVv��Q�YR^`�Za�BXN�z}N��x�v����Ԯ]�cu�Ә���)a���*Qʳs
ߐZ@�Sİ��ǿ�m�� �1A`V�ش��"

�*�4���H]u�ׁ��P�UqFBj�f�-a�V�N�4i*ތQ@���,Ӊ�V����9\Uu��V,oo��/_@���x� �+�Vq;XkK�V���֬#�i�2�fƬ�[�vi��ˋsZ������F�׫r�WTKs �R�fl�	E�-'R��vT�D��Y�ml��ާ"�,Ѫ��Ef悔Q��9�A�7QM�1�un�c7w$�Tbͭ�4���T�j�i�<�9lmT�c�U��V��&��݈+$���e�7�k*�=��B�a$�ʹ�W��lI+-�B����X�k6.$n�7ysp�V�B;�y5� R��b�����5�W�+�tn�sR7U�T��k��v4��t�ZW���E�̙��e�Sp�t�C�Y!\ݩZ���%3k�u�gT�S,��:��ܻ�ܣ�V��5Z5�Ȁ�cJdޝCY�Rn�x�XKkwrcS��%�%�WXC�eo+-�5p�'��F�;�]���x��'������/1e��AQ�63m�c%�ل=D3��������5-�w#!�	z*�tT��JolG[��͵����wY�"F�q�:6�$�FK�*��u�̗�-j�-�v��b.��Pɀfb-+,�F��t*d��*��;�ٰ�ƴ��F-� #���h�J��Y(�h �7�n1�-� щ�|7]JʩĶ��nH��V~j�=��ՋtjI��F۫ۄ�v�6	���T�dSlf��A�"+�ͽ�K�D"iЙr�p!��h�3Notm����%eT�j�{d8��$����H`��a�QӔЪ˱��G�D�h�5�붚(�y�tjβx��,)��,�*8.��1�fKF!uޒV,�{-�b����%��M#N�%ొ�	�.K�C��kUa��
ZV֣Z삛�e�]T�Ȳ�Ժ�=h[G"�uz ���)�
x���
օ��K5������$�Y�[N�J�;q*���J��!��/#́%�Kf�i`%�j76��wYѶ����;��<��X��S&Oe腬�A@�̥�7��weeW�[ ��r�V)O�0��ʒ�]�4ݻ�ޑR���.]�i�#�d �X[E	��F�e�r[�ͳ�ovu7F��Ҳ-���LcC���2���E�	d�d�,�zr�APÂ�&�e�P���I9��nm7s��
��VB{z�m���Ǣ����4Փ�0�er�T��t��a�*��<�3�$0�jA�v7V�{����u��Э��%��I�$1\�j�6�"���nOi��0�mL��h��"hǴv�*%��x��hٰ� c���g%(��-�J�EcWV�(�Pe�"�����o])//XR��8�;AJc��-=&Bκ�`��H��)�F�HD��$�ܽXꅫܑ���Ra�I&�4��$�G��^n(���Z䢓��JnĽ�P�#v�Yn�*�xs[b͚vm�F��i�;/4��Q@SOD
�	�Cx�Z6��F9Z��0�1f��Yv=,*�Ґ�*�ac�6��d�Ac��Z��贬44��Vv�
Ӑ�`�Q5��W���b_���H	W�D��	ص�v���2x"J,���f�˱ �aQ/��(�.�s��h+IӨ�x�[j��j��8"FhX19��ر�3b@�7TD�.�d�.鮣0H��gXD� bh/�KC��h��-���n��\J:ɣ|��sT2�@��Z&r��e��P+1�a�w��'r�'��g
5]LXZ;�P�T>2ړo����<Gq\�Ћ�x�
��Q�,W\J:�A�h�p��B�0�1�V���6N�0�'Ϭʠ"|�]T�il�2���tO�\k$�nXD�\�nJ5����XH8��z�N���İV؞�A�zS��4s&�Ӵ�%��b{F�tLJ��p0��do��.��a����|9��)�Y@���\M��E���Qvr&��T(�u��((�+��"P;Ε�k�:���2�����-�@��̤TO!1��;8&���l�w��<Z9�� g1���D�6��8�Je7��FQ(��^yO�<'���4<�qȶv}��7���(����13���z*.���)�1�f�ɳ+�h@��'M|ʴd\�TL4�l�,���QX2�,�A��.��#JC��UD�+
�\e���0�x�.6����x�(<;��㰤����)EeoF�D�P(ꕜ��0�R9�'Gf�*�E��Ĕ���\R���J�L�|+�F�\8�3��B��4~����`[���ބ}+�q��Awc?���>�c;�_u�4Ks�XYL�G�;����(��ە��ø�pܷ�U����+�㍼з��i���ʔ���b�Z�w
�&��/�(	8_ƪѾ�|u-_��^.���و*�4�Ҩ�"�j��%*ź����t7Qx�eR�j�G�I�~��ss!��YV8K�M{R�AͶ��� �IE��x�=j��z���j���+գR�Lm;���P��{�r" �]�j)��s�:k�.�����Khp�e��uiݺ�Q��V�;�MM8�ܾ�#3�t3�r�I:�.W��˞u'���P4]��ޝU\RQR�.�:�U�g���=��f�(Q@�������4jF��g8�xL���Ǻ�5�ڬXGr��-�ECIy�]���8�:f����3fa�w�us���!7�Ⱥ���Fm �J�+���T�NYG���6����5�G�W7�8]L�4t$�X`�����w�M��H�n���>ݳ3
�����-V=� ��3�:@c4(�V���	͛f���ub4,�+awk9ˤi�H�29�]y9\�y�N\{f;:);"���MG��_p�S��U�9t5����u��T��;�S�_UjJ�J����K5^×�[��a�s6�n8t����5�����W���DI��:����
���/�Ʃ\�Q��Sx��}z�ܩ�V��<b_sK�c^@�9O�;1L=��VG��Wg��7�Agq�*t��u9ieݞ�%�k�*�n��5����Ɨgvv�s2Z�v+A�kv+l'�h�2�����pW}}�ܥxy��k�%q�wD�+�IKO� k�V!�2w+��g�c����Ќ���R���f��z��׵m��|�,̡ڔ��b���O�sE��77�˥������$��w�:�ݴ7�{��H-�k���=�L��3b��	}�o�Y/9�(�b�mj#/h#��9�]��z��g&m6��unw9H���gQ�BP��A��\��7:
O������6�4�Ūvi���w�6gj;��!�I�.`��gem�q�f+�5_]l�*��y�P�q��lvn��)�>ہ�L�qf5�R�돮��\������Ōu̶l������C��fD]�[qN�[벭�)��>�����p4��J�t0�usrN�j�)�H��y����z�wkx1L2�]��Y�Z��P �]��@��H�2(ND�F�����Y�о�;9���\���SW_C59�V�a�|2Ӭ�]�I�;��\�G:�nd�ܶ��6J������7��M[5C�c��k{�F[|ي�Z�2�5�:���f���	ò�܍X��������ud���V���}���$����`�.!�¹K��(�YB�m-��7͕���8�Ρ�ǵlO�\��/�c�a�řyxnN�����cM拢�*���(YU���s����8���n�����:]�r���~��`�;������=Y��{9P]g_��{��Ժ��$յ��<��4Jwy�V�Ar�2�d���.kG��U�f�p�2*=������[k,�J�eN�@��%k�lI������m���Sk
�ڊ����,玖�R��U`ޙ��p��|q����Z�ٝ2ېb�'u�wQ��QT�cG$R�P�ogm�|���u,Bs1��4���Y�2D�q��ϯm,�݌���]�\J*�*'��Zv�������q��ؔ��,U
���r�9��L��zd���@}��oi6��_Y���g(�w=Ff;�3���6`��I�<�p|��4�n�l�SD�ܬ������wf�HuF��g:��Qr���}�)qĮ�U�8��K��]�Vo)0��n�C1�U�<'�bV�v�>�
z�P�8�(��V̪3H���I�ӧZ#��7y�������-�r�!}���VsU�a~3�J��K;��VG����|��N��d��ވN��,w���ʑ�����Ù�j�l[����6�:5�Cz�[�/PF�����s#���1��m#W��U%6�;՝إhu��9
"��3r��Hǆ��+nC�%4��Ί�^��8��ї��o%vJK�a*^rj+�{�HC.�ttv�l�w
���l�S"�іo�6�t��E��]y�u8W]l`Bò�rU�x޺鷀!�w��ٚ��:�캙܍C��N����gm8�s��{�E�e]�v���B�hا�*�WV�>=�HD�S�w�����dN�f�"\u<��e�)�s�(�/xڴ5d������x�go�~�Lm�;�5��H��1�����Hڑ�O��ʮ��TY+b�&u�w����S�6�7M=սn,yZ.s2o:i�+�v�9��9�k��bmi�md���;44����T���]}��
5��w��gQ宄�jd2���5�n#�d��̻�L��6}����ĥ�>��m>��X�R9W�u�;�<c�/��7���W�q�+��.�u��Qڊ�)\X��IU^ݱg��d�{; �V��	�$_Sc�_X�,�V���#�b��d��oo{Hv9ǺDw(��r��t�ì�(��I��:�f8J��m��X�ɂ�ڂ@f���Fg9ݸhu��2�Z��U�eؠ����v�ἤx�"'�nV��o:̠�9YO��/��C���I�4Gs��/\���x�x_ƣt�з��+^!���.k�P�s�}ɻȽ1�'l��N��*1�P���7�:�����_3�Wi��it=��ѵRXS˦���v�����um�O��@��ђ�a�F�)�-@�X�qD�.꾤�W]wswOUL��K9��qM�r�c�T9���u�l9ܨtu6��e������xh��Ք8�Xw�� 8��������5b�9uZ׆\x�3 ki�kBYҡ�q���g���M,�Jpfb�0���6{�r�����L��V[=|ȩ�4L�����X��}{��jr$i�A�Ǥ�Okr���:��Ú/�FƢ8]�S="ذVpy#����K`~PQ,xI�&����[`�VM�6�b��VMz̺�q�帳��6Z�g����e��J�<j��Y��t��fH�幏�ٔ�]����m�1���}l_"��f�3�P��D��I�o.��#ð�g7���M,�ֺ�*�>Q��>�[��db�pt-	Jѹv�-a
F+{���*��BV����w̍���{b�l�NU�Q���xk�a������Wf]u\_u���l��[nɇ)�(�uOlJ�n�u<�'���Fl/��B��qMd�V�J�ӵl��sc9�Y����Oq�5D�(<�dIV�R�z����Y�\��:�u���}{����'�2(����*�	봥���K�4� B�����5�T0ȓ�\u��*�{���wPBK��E$�_R&ыz�A��۫���٣��,ڬ��p�{��TS�ȂŞ6�]1�+v�;y�(�ֺ:z��}�P1k�R�mc
Ia��	w/������{��Ϋ�ڃ;c�:�@���,V��\�q������,����L�c:�����'qck7AU�Z�J��j��h氭%�X}'��m>j�Uc�TN���z�K�Xze�EX��b[D������m+wE[ڊ�wf���Zn���P���u�ч�}r����uc��/����W..���{�݀�5Usuv�B1�rvLt�]�t���{M1z߬6�p�c��5�)䥼�h�����.�؞h��(�*<��	�*������ebnݙjδ���-�/�*��5Bp�
<ӂlR�ވ�<���4#�zu���8�����q�tѺ�y����;y�m�
��s��Cc����z1]A%h�;3B,�`�ŵӄ�8^f�"��w^��F���v��W��1�Mȑ.qӖ.i���ͅ�Ɋ	�J�����^{��&/{i���rUd�2��A3���`��fea�;�z�������1f3�N�^
�f���C�Q=x6�yP�U��ո�Q����;�ܐ*�b��Ԟ.����Ȫ�f�TB�]�>��o��U�ȇ���[t��X��*���a�{㱂�:rރ\�ug):�W�CqnH�S�܁"N#c�jzWUd�fK�1��vU��[0c���g)M5;�]B�����[��r������� j��f���jk9���p�L�]9R� 5�T_q�#�-<״�)gWf�;�a�ܨ�n���g2^�+�ʐ0N�[4�\�WީՎ�r�q��-X�Q�n�5T�K\n:�q��E8���ju5�@C8��:
��V;e 77����Q~���3s�T��xFr��r��QNf�Փ�][ϫ�<��܅ �g<�v�gN�m,R�t���[�'��M�K�ϏK7�ykܦj�Ŷ��Vm5r�CD-B�%�l������t��]�sv�lͦt%uGcr=崀g٢���M��\x��K{�9E.�NNv�sUP	�O%�*��,e;�r�i�n�J�n����F$��d�^�w�cMvYY]v�h�ٕ�[4˘yQ���oE
�����Ρ@�A
�H�D��l�L�;(����Hə�'�n#�`��d�HteϦoit�|wz�voWU������
��Ƚ��P��袵��]c�����昳��nߔ:�ӻ�*���6�jA�L-ة�\�֌�GzV��)*Gs�e2�����|��t���*��$r��\��p�W%�EnPs.h{]yKn�۔���ҍ��"����͝��=�2�������!�UN����/:w)��K��`	�hWR� Z�|3,hS�lnf,�hڛ�6{�>���'a�J)��0k��E�;���j�Q�WK�6��4�4*fa鼓B��XUsl�˒֥��ST74��C@����<qr�����*w�"[�:�[#(`3��Z˫z�;��d�{��֬�B̓�T)+[Ht�Kb��G!Q������4תv�ξ��b��f��.Z�b�v��ڨx\b�`�c;��}Y�6�5�0YM�[WwM�.4v
*��}*&1��8�:���T�����2��G	3�ERɝz������� �V ��X�{�\|���	b�^v� ��qp�J�R�%�P�&��j����-	�45�ާ�rέ�6�a+�����-��3v�~�zq66��8Q®�f���z�X�Up�-h�l��)��i������[!�z�)�ˊ����Uݎ�7\@䬂V�Z�Zp3��r��Wj�.r�z�]4�Ŧ	�=ν���+]�zǻ�+�"t��m$�f�)0G�ֲVR��żZ�[9u=U}lf[vS�Ή_L��p5o��xu	e���$!��D��4&j[Xt�x��عB�7V�+7��T�qn�&��I�e��߫&{�\$DÊ�2i��;�k��]�SN���>omO>�X�t�-X�����3���A��{�b�����|�E�zo\�%�3f�T�\��E3�v�J?�oZ���y݉g����{��:��gM4����녮K�G���6�3�E���%G���;�Jq��_ãh�>,�m�#]��gIgg�ZS��<sM�(�H���RCΘ�m���A�g�cS��-Ҵk��Vv�:���f��EE��(;��]!�[u�v���.pi�j$�˒�� �Y�8ݍ�}ջ������{�U���٧���ݮ��;�c�F�;�{D�;o�ǚ�]��W/�ck%�ɓWU�F!t	�oP1^���&�bƈ\��6��K&6�d��ES�����Sx�y����Q�D�� :t`�^�x:�[�]���@�c�x�fK�����p�^j9�:9�ۮp�`��aZvAZ�N�בz��X���D\�3|Vl63�����������+�ʺ�tA�K�Z��V��&쨤d��@�Q���Fb��.��, �︎�f��wƻ5��.eՑ��Tܳ�+���7��]e"��WeB��'��-��7���'�L�2���Ww\+��;����v�t[[��z���a��sĺ0.�7�wO��[���|ɝܸ��$6)�N�z#7-v�iH ��g^wXeq����1��̗����}һ{���W����"_ח'[�t��O�\7���ӻ;�/+s;���^�<�3�u�pO����<�>�b�������=꜎J~!~��}��
s�C�Ce�<��ġ��(��QF��z�`�O�~=`�c�>��|�����D��eB|�����~�K��0�Hv�"z��+� �|��rS솟wS�~}�~g���u �`�CG�O��e����W!M��d��{��	@z���b{��@!��W3ց��T�@�T�~����C�����>�?����� ������������/����>J���.n��w6�R�&n��ӯ�����!o4�[�iLIM����Y�S3�*����k�à9��Fb�Y�g`�z�\0*ݗXSus\d�I��t��N�꧊���5pW�+m���r�*dp���;��.�֞鴝�6B _,Y;F�q�aq�ݡ�Mڝk\� i_eʕ[o�2����R�̐�P��y��E�)ڧ3����y:0&P�G�q��4 �|W{�V��6�������B8f�s�e�M΂�,�Z%�GT��`�4}P=+9k��h;Ǟ��^�R�X<3�'���<p%�gnf˽���ȝ��
K(�ۤg�c�H��O�7��L�,�������,�\M��s}�����oʣ:��8Vݟ�EXZv��_6����(7Ɨ�'C5�h0e�
�9!�E��X�]g�Uo(D�s3+A2���x�W�,�ٽ��%��m��]!��F+Mg+Md�K6�}��[f�]=�p�N�P؅FOn�W"�����"���,=�{��\�+!�X�k�N��m^6�KU]+d�P�����3ݕ���qb��� �+)t��i}c�s�'��m��4�p*�ё��O�n�V�ykx�P�e�{ʂ�)��F�r�֯��t��n���zp
<2c�/h3/������}>��u����������ׯ^=z����ׯ\z��ׯ_�_�^�z��ׯ_�Y�ׯ^�z����^�z����ׯ]z��ׯ^�޽z�ׯ^��q�ׯ^�z�z��^�z��ׯ^�}=z��^�z����׮=z��ׯ^�Y�ׯ]z��ׯׯ��z��z��ׯ^��ׯ^�z��ׯ��ׯ^�_���������{����{���w�����{��S��0Vfݾ���
	R;�Z�kxV�s�]j�'32WJ��V>��r_*�\����Fn�+4$7E�{܍j���>�P�����:ܳ��H�?JK�Î��tp���Vu	(l�$.��՘Lnm����ù�qx&�Kc��m�3v��JC��U�{	JL��(W\��E`j��\x�C�"4�N���=�ڢ}DaYw5F���"p����y����u�UE�1�WKh�\�ƥ�ȝ3�mĠ�&pq�p\M��S��QS&��"���(�j�38� ٹr>�C���U!�}�N�nr�v��	��`���*��Kp;�qO����Q��kF�);�{� �x�ݽ���Z��E�ۼ��xj�94v�|n���u�L��v�7A�P9-k�Z�р��Stl��8WW���6��o*�|f�W���Ta���Ur&swB�iز�j�2�7�v%%��*u���3)>ͭ"��m��¯.M�5k4��!3�Wx��ٺ˘T5��E�噱�b'�ݻ)F�a���@��NM*	�Uw�J�Vc�l�6����[���i�7�:o���)m����J�.��0�g�,��$'Ø�)k.q�I��E^�{���S�]z�����^�z����ׯ]z��ׯ�z����׮=z��ׯ_�^�ׯ^�z�����z��ׯ׬���z��ׯ^�z�z��ׯ^��^�z��ׯ׬��ׯ^�z�z�ǯ^�z����׮�z��׏^�z���z��ׯ_O^�u�?_������~�z����ׯ^�z�z��^�z������������ׯ_O^��ޞ���{�ޯMw�ij�oCܰMƶ3���t%&�o��� �;Y�e0��{
�.���ĺ���q	Q�Q^�D�!ٕR�;�G�49ok��^�s@hڳe���a�5�a3'N��N��_@�tbX��������Ӽ�Js.���kjQ���_R�vr�)d|Tt�+^�x<V���u{�X��U�G[��Ǜ��gv*����qaۛe�Rt�Z(g)ƅ�3�l��]��(�2X�Z�U�#ۋk��������6�!f�^�sB��}�k�ͦ�㮝"fHcTL���dI�:�3��[MtM���D��)�\ngfpX��S70�7���͊�t����g&�	toR�;��g�d��᠓�c5;��<8��N��A��.�ʹ8��h"ʤ��/���o_�:.�E0_�9q����Knŝ��Q�,;.Mͽ�r�fYA��A��ҫsl44MRf8e����W*��i��F-I5�Cs�M��o�������y�f�u�N��3�7�[d���wRl9���J��]N��VeXt���J��af���g�M�-]�/���D��U��W�:QRul�ڞ]uZ�k�|�����FbFD�`��8�ʍ�n�_�������{}��o�����=z��ׯףׯ^�z������z����ׯ^�z���^�z����ׯ^�x��ׯ_O^�z�ׯ^�z�z��ׯ^���z�ׯ^�z����=z��ׯ^�^�^�z��ׯ^��z����~=z�׬�z��ׯǯ\~�Y��~�_�ׯׯ\z��^�z��ׯ�z��ׯ����������ׯ^��z�ׯ\z����t�l��cw�$Œ���N�t;]؃Mo�&����� �eu��0Y�ִ�e���.GZmexb&6UF�&<[R�C�m'�Q�34[B���Xzޝ��
�ӑ`F<�3�j+���k._.���	V���mj����S^iv��s"m�Ԏ��ō�g:�ɧc{��l��t��KK�*�VP�,RZ���:�*�]�r-�m�g<ܷJ�R3¯x�tđf���7�{���`�zn��u5���U�����`]��
���m\���F][��h�Gi�j.[�)t�+��8��%��N�C����: ��M�L��DDw^ж��Օ�LH�#o�;;���IS�+��A���z7z���YiUk��vF�B���M�d�w��ъ�`�O�5��ܪ\;.80�_,t=�N����L�:6��	n�ݘw!�Ӿ�|ޢ7B�|����*.:|���ĢD{�SCvAν�Ŝ/B|E9��ԱV:�[@̭�d�y�T�A���񞍻���%�Uh��z�ۗy9��v�ܳ��8��e-�i��G�RX���NvTxFnz���I�NPʼxk�+Q�J5�}њy�soT�eܧ?W�U9��q3�(w!j���t�u����<�����	a։�Γ�e��y��n��P������Ϩ��T�F��I`J�zRW�:B�s���a�P)�oK����%������� ��B�I7g���K��;�K{hDb��WP�&A=��a��Fek�� f�/:�7n1�V5}�u��B|�J���<Cu�L��)"aU��9G�G��k�����X��Cy�A��BM[�w����8&�%m�I�UU��K�\}�g;���X�B�s�S�8��ެ��.�]�&Ԇ��U�&��L٬]ծ'*�Tt�3��LQi�Qy=;:�P�޽~���V�A�r�eowY�t6Uo��C��vn10b�����hZ��e��K3�9!ֽ�1l�Su���嚦A�7\�eRr;�ld��"��\+F����1���<�&ˋ	�4�� *<�|�P�:�v%�����`�e	����}ȹy�bǌ�ܞ�*��Y�od��h�x!B���P}�4�Hu�MwT�������&'C+����;�� �%*mҫ��ݘ���ru1-a���֪��M�z/��:�`9�xs4��N<̺��%7��S���ӯ`��XC�;v��� 2a{W�Y!�{@=���.�Z�����熵�����C.X�؟^V��M��Ӑ��\A���B���$T:�a�m��3|z`��ʷ��m��Jfǎ��Z}�N2�\��aT��q�&F��5]�5���t�]/�]�&�zp"�W%]#,�E�i�}Qs�]V�{��R{7���&iʑ
.���4��*��f
4J`V��k�S#_*���4�	]��ގM�X��})BQ��wUl2��'=;F���⵸��sٞ���epݓ*��fV�1�A�u��7{#}�vh��L��������x����eb=��**�|4�G
nk�kE�vh,|:�k���B_:�r���!��K���,1� ްm+��%��Y5�o$�X(���\�k.@�:�]��0���F�f2�_	���8���'���K�*{i�ok���ou]�#/,�j�Q�fat�weN�ή��ς��#yd���i�X�M�mڻ�cn���X��νj��Jћ̺��P�{%�4��Î��;R�d�adǶ=��g��gM��@�;������&;����~��e�rs�wҵ�ɻ`7Ө>�F���H��Y�UU����?lZk8��v^��}��YF;�2耄e֫�E^��s칆ÅV#v�f.�v!���Q-}ZB���Y�����f��u�M�P5��a����&�3��yV1kڮ��S��6�+��L��t᫧xrqJΉHi4�*9vq�7��'@˗�Wqj�ft�m�I��s�#'6>����m�}�2L�zV���|��a�n��R�+�؃R�����5����c~��y��U�@f�9ou�K �՛���͝[���ڧo�P�Y������_!�����I�|�' P
��)u��}���+ָn-��z��A \TORi-b���	�[�[ʭK�����ݼ��23��v�1Q�+6n��ZfuW����T�^fH����A1�;Q���k�q����:rD	6+d����߃ݩs��X���CD�`�~f�h��U���=ض��^��md��S��oJ�} )歩ե���1ŷ�R[��A��(���^Z�sx-u]�s1PG�N5����ӄ�1C�q���m�tp|�L.�J%V3:�g�Y��0�y���ݘ=`�͜9���������н�N�� N���^R�Y�X��=�ѥf�F0Ի������$A��S�d�B*��FLŹ@]��b��m�����l��Ӯ��Z�,��Y���WA�Tw���a��HV�f
����2���ʄ֬�_����]�tl�WXxC���v�Ss"�֘d+�Z�˨O
ٕW�%�|ҹR����A/���f��^�r�Rޫ�[a��&�*s7�$�\Xy�D�l�EJ�������1r��N�+R��>]}�{�;�C����rC�QVwiB�}?b�}��ڻд�PP�)�F�;Jج�9�Cʭ�f�}Z�b�)�wu�.�Xy�k��ӫ:F����������>��B�wB*@��)8�WoJ�R2��/�V��7�]W*�	2y`�����_z	�`su��W��&ڔFnJ\M�W��e�U�W7��c��8�f�n��� �7a�[�]��7e��''v��n�91�Z����x�|������>��QwJ��w�}UL
�Y����i�G>�ۄNz�E�Θc�5D��;�v^_\�N�N�)M�[.u�vͽtd�m�J�N���uOu �V.$^(��+�.	��άl\�}| j�*�C�t�8f:��+1W\�l��8(�Kg,�^uQ�,�YO���'�C3]U�:O�7�X�tN�U%�ܭ�܋ǤX��b���j����ym խܷySJ��Ԩ�ޮ�Dt,�U�M��j��m�rM��ŷn�]q �u{�Ay�]�Gvu�P:^�q�! ^>�óF��9ݦ�f�e��l��K�BoVY��Ѝ����A�\��r���˜��C@�s��IN��Kݭb���{��C7�^����ٝ����^r���oyo%�C�w7�]����v��/�}�
���aX�/t��6b{3��z�_'��G��d�8p�}d�]�Wkgmh� ]��營\]B4U�j��1#�rI��\�i�u��E	*����Ym��Q;.r�R՚�Y�uu�!�֥X��{�U��{�jR̠��M�pN�u����7���+8>���yGJF̬i��.80�n�����w�=���9�"�Ccm�-ٜ#���-�36��(�]<���������bWVӬ�uB�P����� �]�2�ía�P�7,�m��YA��iNz$n�9��6��*V�SY�Z�oJ�5��x�7I��.���o\�;�0�����q�-��2�`BeLd�z����[ű��֙��N�۝����U�P���Q�_D����<x:d!����G���7��{v,���ݦ�uɂ�Nꡌ^=����YK
�f�n}4Q=*ı5���;�=�r�M\�/��]�Kɪ��=�,x2k;Z]�)��7�܍R�lUqZ�>�I��ޱ���#�^�HVs7�4hFM0�y���o�׃�[Ƌ�G1�4��f�I��72�NjB�c�*��P*�̧��U�瘜��h�J�&�aW��)!g�4pG^�׺;uS��<��ú�R�X�yq�|v	�q�4�c,.���T9:����]�cW;U;�k�ճ;�I�$���`���]��J*atuM�:�Uә�9�Ok����Sm�����B�T�����<�}�I^0^�3��q�d�鶺���:�VU�N��s�/擹}{1���Ks�*䲀��K��4���Wb��Y�$j��\��wmg�b��\h=�_gL��^�K�[��S�gIpX�}�0;���g^��gk���=ւ��򹹚v棪�}vTN�n��e�o���{�veZ�����ք�r��fT�}x�Ҷ�+�vQ�ȥ���$��]�;mpA��
���ei�9X�$�60SbF�	g�CP�MnUB5��O}tO�A��z�=k+&�)u��V�u^"
� �
3q�$�z��(��C��V9,+��gAëo�eM�1�g'����O;���4{9Vm�
G�`��˜�zވ��qP�媂��̭�J��F��Y�p��N<�&�!�z5bOj�40�v3e�.�Bu�XԪ*�c)V�W*�;���VM��Z9�sS+�6'���xo���ԂԻ��4�U_J얒+O��eLS����Δ�Vm.���姀�sٌ�cK��un_W>w�yv�:M�o"��V�D�P_+��*�� .0��)�8E��2&'
n�V���,�>�9N�����`�����7�ײ讝g.���%��q9���Gc�8m��C�meZ�s1SPSX�G���R�+����&�F�mQۭ�e�������������?��������z�����?\���T+��H�!YE$�i�|ӟ�!*���H��Q�ӌ2
&y�5D		!��a�j���
��#��B�aB��4�	�Th�g��Q3#r4>!��D���,�[E�-�$��" �	��)C�R/2����(���f"Ȁ��p�b���&㐔�QR(�A�F�e����Li��!
��X���hPL��AxF�MHH$�HJ���S�(���*{�\�V��k��cEx7��.:���r�J��ȏ1�{��n۰���gY�7xRv�b�����s��嚵F�+��2���[�53Wk9-ϧ^q<�jG�����d�Kx�Yۘo���::]Pe�!�V(/��g6F��F�Ӻ�˻2Ko-:"V8���]Eu�#��^�f�n]&kCmms�M�Y���!6�%���D1�̃/��v��O^	Ȥ��I��j��9^�o��t�Ci�y�Dt���5��U�j�y�z+]�L��w9عBJ'��]_���Dx�n��Ǜ�9Y�r�U�f�(�8�2����\���s9/�1��vMPeR/��gN6r�J-�ʬ�F�f��ܜOq�j��Z(�9��7{ꂆF�l�6�CR�dJ���,�{�C���N1|-��čB:�hzG��5�wF�/�>��i�:u��fR�w�5�:�nm�aC�^b�ٶhk#J*K�{��8�mh�����$^�5y��9j�=] �TF���K%�j��hmvn�r]	݅j;�Eq�)-��uUL��K穋��,�5m�͑��\I�*s�:�����qÚa���hͽ�((�-��PH�-�]��b�����O�՘L	=���ow2�X(i��ap�P(��	/2~1���7!E�"IhI	'B�mБ�dp)"ə �@\@8̑�BR)Ex��0������e�ߒf"�$眉�<��$�j5rbq9<� &#L�C�Cq�) p�!EERH�Bq"����i��m&�M� 1��Q3H��e"�f!!l���(�Zm�R5MIS����Q�B�ImQ�^EPEĉ%���**�x�
E��qE6SpDA.��	Lba��a?$�ă�HJE�I���ah���&!HF���ˑ� F��z&A$�2E	/�0Ԓ
IG�	rB7�"�A,!��N	$�m��GB' R6FE=E$�đM���7��`�!�ɍ�YBѐ$RHӁ�1I��at���1EJAf�aƜ�$�ߙ`"U8�z#i�>E���p���F��Ӗ�z)�S@wZv��͍�`�2���pJ��3�c#)�룮�~?^<x�����^�:�;=�#3�lC��Ƞ���r����&���-�7q�33&�����x��ǏG���3�~�.�a����FFn��r0�̥�Ī}z�`��FBe�Q�p�������������Ǐ<~?G���3�Cʛ��j"�$671�E�>��cq17
wv�sj�9��.��I��W22\,�1��e�+��Y��;el!�B�Q�a%�� �@�s31���B%��U��Y��K r*�2��2ȷw7sm�1��7,�0,2$�$�7�n��74&M�1�g.G76#1�2�61�p�u�m�:k��m���Ƞ�&��b��-���Y�7�w���E�c�ÙfX`a�a�l��2 �"Z6�6L�2�l,����nq��7,7�����'�̳w13sL�+����gXW3(2�7�1��H5�p�
�����	A���GK�B!�M$��D$�E JQ���̃(�
lȲ-�7�.k��-��-��3sr��(�6�͖�m�m,��0�6�-��sK���s3#7���r/\��
r=NA�G�'��:��p�`��Lp�\��`����ld�ف�4QV�nf�9�n�aV�dEET�aeT��*#*"K�p�yn�f뛶��7xF�r �C�cM����L�a����Z/(X_Wqa#ɝy�:J��J|L��F�'��sM竷�R��0�G�IinOV��e��\9��	#�q�d�&��A�����P��Lq���Ԏ2#d6�e�h�\�(ג
\B ,��l��2\l L("�E�Sh�D�cj>^��"�d����%�"	e�(��DA\�W�[ǻEfW�O�,k7�;�̿�c^�N�B����ù��NR��o�w��U������n�~�V2�ښ�\m��_},{�q��y�����4�=�O�ݣ��>�m�����:.?Sk�fs����ϯ��g�܆��&��1Y���3�k��w{���zgu�c1��&w�}]��Z+��i�*�CwW�[�����{�׋oy�}��e�q)�v6�����Ԇ��;Y޷�d�K�{�;fu��SL�w���>�c����N�w'�ͨ<�FWk7�hh�������f+y�;�+����|s�E������h:�7�;��
�̈뚼��#�=n��f�{@e�Y��h6���2oL�ޑ׎dq�9f:<q�+E���Q�z:FKm�t>`-|��L�awƵu-�{��˔4`^�<6��pv<��W�.9��:Er�Rz(.�}�I����1l��p�������"ȋ��πJ�Mz��o��~���}��CE�J/bЭ;�9�������N4L�Rw�8_�]E���n��}��j�_+|T�ʱU�ӄ&K�˅ϸ�7O��͒���� m�����M�I�-.�;bY�5��&�OWT;N�?�O��zC߶���4��� �O�Y=$3��}�51�y��׏���{k��ɾ�-x����},1���V���\y�m���^�����9}$�O�z���V���0�-�\�18#x�s�GWO�l٥�(�����*s���w�<G��P^�u/+��u��]�^��{�=S4M�F�Aj��^��FO�jy��f�Y�5�2�鿻;|�av $�Lx�J���l�BU;_������|UWE�� �B���bSO��Z��k��>�?E~�$}kV��w�>vz��Tרe�IC�+������c��U�|��^�;�K"w�]��;��[{�2�*��;���p��6�t17��8g$���ce6oUJ��i�-�~��G]|>��q�f�W;�ˡ�֬|$�����4��dzk7����.M�w9����U��wu��0�E���`�9M��<#�F��}vx[2���h=�����e�΀���ܘ�sZ�F�h$�xȓ)�U�I_9���Z�=��=�XN���ѽC�Ne�I=f���i�ut�[=XU���jz��ʭ��"=�%�����z�y�#�<휿_O��l�������z���#u���	^���'�s��#���=�zx�.��K�X{�������Ev�?������+3��2����5��~^�}���O2��[�ya&�D	'r���j��2���؞84���<0��o�a�����T���r�휮�~�Noo�G`�`�6O�D�\��&����eQ8kӽ����L\鿹�Z��z<���Л�v[��������^N���\��;�R^�=�]1�کom+��f��w��%�q��e����7�Yo�c��k9�3�T�j|��5Y�S�	����k�������
�^��l��W>����#����f��Ḍ�h��Ψ4�*�`���e��s��dk/�Vs�I7�\��}��c:1���^�z����6��H'&g^1��V��� ��^������c�vq��J�sw��zR�f��SWk[ƒ���ݽi�rÍu��O����»�W]2�I�3{1��
��m��X٢�pa�2͠�3�M��@�����+a��FM4�����3w����/���a�-P�����c���l��i�4������U�����.����,�U���{����y����ͤ�z�kxC7={D$�w0v+߹��o�w#���5U��w��|S��5u�h2*����<N'xl�䇫�WP=B���[��\7�Y���8�����4����P�5Z�ⵝ�Ω7��=׉q��9|4Fs�4�1=����L
��%�t�#����A�,Շ�X=76���N?S�n-���2x��sB)ӽ�}{�޾����� _yJ�nN��6_�E��L�o�sw�ә�}�g�h\]��z��[�;���r׫���z����y�2����T�y1�{��~��J#]�۽ӽ�bw�z�Oަ*{H�;9�/��{��t4;���b6ܔ	�3�'|/2���M�[WK�a�4�N]�e�/�7@3���ݛv~v���̥�.�$ś��A�۱*J��ޭ��W���UE���O戗\U����4���3��D0�i��d&���ôXӼ�&���H�P�\-�DM"W�ϼ�/�X;������v���y����C�!놓��_n8�Pc#�q~��dh_��ŵG,������7�π1����=��n�t؍ަ�l^�9�|�<xb�*Y�a:6��z:0�d��_Bf�kǴ]l8ЏwS��%��g�5�ۙT�ԯ{��'�yd���q(�!��ާ�`�~W��7�Um�Yrl��+Ƹ�di��74�2�g a3t30�\\���-B�k�w����{�PY����%��~�k�5�H~��u��wg���Cֽ\���Я6EtU��#����m�>�v2��s6�߆P�>�>������gL������gL3n��L�����=^I]2�����E^��q������y�vܻ>��#��.���]zs�s��zN�2I�;�v�����my|v*㓔���@���+�v�M�$g��>��݉f�A��)���pgu`0�-˾�s����w�x{�/v�(��/���b�-t@6@ƻwwNMkLܺ���S���V�9�;�^���y�0�ۇy����T���G1�w�u�GEg-j鍥|��6�*}_U�H�aےY���9/9�����2Vz�.k��)7�#�V����<�{���_m�f�Ɋ<\�����1��v���ť�i`w,X�.d���@n����9����Q�;�:����;y�Ӹ[z�Ou1]j�)�^�緻�����_N���ǟ7���)�9�.�0S��#�ma���������b=�a��7_�W��M#�A)7�;�ffg��;�B�>�~�ߏK{�'m	>\�1����|kh.���*���E���J<��/*�.ѕg_����=<���U�1���*���<MB�J��E�"��vم7>��_~�뷗�`^6������{��y�a�U�3��8W#�D�ר�py����飳�[�r`��'z*;��oC~ U�u
�����|t���{�o�y�>���\�	����w�����e�˂�)��o�[����s}2i���YEiMo2�N���z��"m��h�^
�³���Uӥ�Iv�[�/��$e�p73��k��S����gU�Kr�>5�j�����+�S+����b�_�[���V����JU�{���;�fk �p��{�=gpyY�����y2j��^����M;��m]g�sS�=�x����ݾ�W�����x�]��S����I��f�3\����m��0"={�7�G�`��{�+ܗ�����ڮz�\v�Q�|�����X�����a3O�;�ɢV�@~�۝8��k��}�9%qހ�ڞ���)�+Օ��U�D��uC~:��yIOvz,q� �zoY�r�}�b/p�'$}^��k*��ʾ}�$߳=;G=>&���`s�{g��Y��}���O�����N����.ޞo3ߺN�[��ȭs��,^��n.�r�B���;;]�>�w�{��sK=��>�s�%O��~�%u�A���z�|}jp��wE�z[�s�������Z�u3�c����?֥ �ͼ��(�Օc�J .����X�VM�����]l݄Z����|ױS������,�u� �e�tw;��<��S��\m�iO�������6Ha��e�滮���ns�&�¯��x��A�ޓ�ځ�ѺC޶|<�U�\7+�DU�^?(h75��q3Pqڝ�f��4!��p�n�t�떨.8[C����ߩR�͞g�]Vε��54u����v��g��kb(�m߁�9=�
�{c�]�W�<�@M��l��r�|��j|�Y�^��}8�mJ~��,��^���dUw^�8`�����'K�vh�@=��w��=�Y�ǩ�=���B�-�"�<��ڙ������-~��I]^{|���誇���e�*��y�-Cyb�\���}���29���;@�����u��wv�b�0.��鳛���L�m��8|p$�Ϯ�_;���-�|�{��̮(p��b}�w�х;��;�j{���^c�����p��a�4�{�ӹg�\=�8���̧��T�GΔ�Q>�>��T���G��4J�M����=����X˶��ƺ��;F�F�[{룰����]�g}}(OK���Z���}&6�v�1<�wVt��V�A�ۮ� b��l]{Q��w\�y4:*O���(�F��a�ī��QR�^wW�TY�X(��1!5n����kŁBd�Ɉ"	���XDU�A>_�~���n/�`}�M��� \���D9ك:��/ziB���������w�};�N��o����PU��ܤKy����.K�Yv�k:+�ٮd�QzƜ���l�U�ջ���x�Fq㱣�(U�=̞��*���y|�vDz^�ο�*�������]�����K��6߰Q3L7^���:2W�Uv�G�}��t��n��j&f��cz3�d�����4f%�=�W���-�я�^�w�^N��^�� ;�e���@ �A��s;�b�x����Z��S��cc'{Ca�F�qy�({\��w5��^���϶>��v�쪠B��I���� BI�f�s���%a'����X�����o>�k�H���茷�rpoi'�ܐ��lt�ĝ�;;�M%ﺯ6�y�x���MW�;���(-7c=}�E��^���x��Kl��-���d�����C_`}��Zz���@%]����]����Ͷ��eJ
�u������@H��2���u�Ӆ6e!��8���x��0����5.�2\JTɉk��D�b��	���`)�ZIvfQ�mt��}����Y�2�ܶ
�l5!�Ԏ��Ft�_�d��8��+�NrY��#w��%�Wus5�߻�[y����;�P�O��	K)�<�q��zw�OQ'b�Mi/U�;hS�{�WV�����UU7a���7�K����w�zoH��6���ڐ�;�Z;����a������{j-�:����>i`t߇<�װ�jwF�v����р�l�3����N���9�d�w��9�GݕD��{���~���}F�Y
������B���g�7���p�3����N5�����dT�C<��1y�&����kk�D��x������;��2".<��"�{�ƛ �^�t�9�=�i�ޮu��y����St��l�w�9��������l���p8k�l��X��8�W��]ߣ��|g�����v��<<χ���'���>[��"��_~X��� �v���rُ&ݮs�.E2|]U(��}��iI?]�c�;/�)�f�������G'֞YS��gi�U`���t��4�~I�B@K��E��m]��'/y;g��ԃ�f.T��r�S�U˫��r��1e�6U��&caZ��զ#cN�4�[��39WeDx�����-�r@iun�s�}S�NH3�4_$��5���SF͒q9}��9�pf�}c�^��l���O��8Nۼ"��oq�I�lȬu�R�wwP��e�>��E��N�w�rZD�iu���fù]���^tb�ȍ�"�[l�\�2�Y�i���4N�{r���F3�'�;��fdw5��� �#���2D�q��fe��y�r��Z\�y/�1�J��c�����>�yf-��eֽ�����Fo2�MB�!P���N�gV۵+��0C��x���< Ee���u�9Upq�1A�,<����M��{\�40F����U�5��;��}՗ƻj�Q@_e��+���;Y�0#Pvv��t�=N�������;�M��<(v�tk2=Ɯ!��(���;/�U��V�y�RKN�f[-�5WN�Z0n�ܠ�"��]:�w�]�j������[��\�N��[���9̮���!�N��n�X�����*UK�غ3��UN�d�3���ؤɠ���Y�%�5����5g�F�F���"�$�L~L���M��/5��BH-��V>����/���\�^�՜�W(���WN�I����X⍮�(�%e�q��ysF'M��	9_l@Z����δ+����q�ˬ�v�J���{	�"��VR�k�_*0��N)w��s�vfI#����*ViɗR(S�Y���ND�e�wF�.nB��J�E����nIvI�� ��p��wy\���@��n��X��ҋv��[�E�Y�\pr���f	��n�]+,+�Q��|������>��'�N�\�vä�:�md���z�q�,`��K����I.d|
؟T��u+���v3$�T(�]��K�YР��]��k�Z�d���?��P�7�cs���܃�o7X��wϭ2����W�����ݖB��v�VR��F%9ؕ�|�RIQ�f�"�N�3�X����wap�rV�f�f�8�����W ��!�ĥN�2���F�����Å�@����h�6�;	����
zh#���3�-�4�p�u+�&n䵣�$Û�=�Y�6��N�oD\$�4��'Mت�
4NA�ؽ���D�Y�.9�C��+qg�Ϲ���e�
���S�u�|�Q�)�'
����5:�l�gd���6�Y�"[���&T��V���V]�t����ML���q|H1��O���7L37r+�dE �,���s1�����eU5LU���"�����������Ǐ���������3a��Y��U�d�XU9�g5ݱ�r<ܷ�3,���c*��6�8\�}�<x�||x��Ǐ������{��a��cIa�TSr0�|�M!�P��nem�e���X��1S������3��O��<x��~>>3=��ƈ(��䛖li;�Mf5�����9e�9E茨"��M���囏�Cʲ���bZ+32��,̆*"������;|�)�Ɉ+0Ʀ��vf&�U%9P�U�e6�Q�fc�NY1��I6tؘ�NYz���CdX�����-�*��0*	�s0f���"�� ��h�"���l�Ct����@�cp��3>��fE<�60�C#"&���	0�"�!�i�(���+,��J�j�o�W��l���4RD%�g�"��,�̈���f-�7 �"i���()�����������y�;;��8��/z.}�����_U�w%��X�,��X�|�*6b�&�s%N���z�G�x��r�*u�<=v�n�vo&3�#d7t�mk�-�Z��&Kz4k��;0���oV��({��_��d{[�j1��f�>̠�f���9��%��QE���NVe?RA����i0��7;���6;�2x`s×S��}���${��ݫ׷�6�V�����u��U=,�SWtsi+0��;e�:��_��ߕ<xO<�������p��\�xrQ�2����5�����\������x75;c����M"q|>����m���`Oʒ����L�� �y(�]Ϗ~P]?E���m�Z;+��-n�^O��%�f�zf�Λ[�Ȗ�+)0z1�n���|��KE��Po�xX��yߏ�^������SK����7q�ϴ�wE's�yO�ا<�[=�1���!�6�T�bz"R���f�>,3��mo,��}�9�'ܡ�*�Z��Zp#�罪�3�M�� ���q�8k�Q8�ۣ&#Vog!�
��M�Q���?-�[�o�k~~�ä~�`rω&[��2{���k�6x��:�pԝ��������»1���{���!��vMu� t=dߕ��2O�{����L2��X�����`3�R%�ҕ`���ץy[� 8��8z��0V��K���w�k����(Sj�v�S��<�G�G��7�3�u�ݫn9�']%����w ��^��.��J�ʅ�b`YZ�E��\Iw#z�M�����v9�ݔn�Dŝ]W���x��<@��kxv�>���u¹Rm�rzc�{�zI&i@���1���Y.��T���Cp�����9��i��gT��/[v�{�Lk�= s p�x�<5��va����4��s���J�~9��O�0M9Con�>�E憖j�����=1.�
<���[����:�B~����g�kV��?qrTI�-|@W�9Sn��W=���C=����#kd����[H�}��F�ZG�ކ,O��sDxe�Y���׀��Pg�w`$9R��:ocĨ�h�����޶oP&y�׌�7�vhDd7�׿�_�n��/��"Y����Et�����H��s'я���^׎.�1qz��������5����"b����o��Ԙ���X���'�H�0,����c�	�V@�Z��(���X�[�������Aʞf׳p3R��b��˺<ڢa彭φg�y[ Rz���2����I��@}*ߎ��@U�xJ1L��o3t=�A�I|%�j�s��S��hc.�����22/7�x3�$��f[tl��&�����OE�'�ۡn�z��M�VP��ʱ�)�tD8��k�L"Ai2z/V�.��̱4���{��3���t=�G�[�+7�.�u����i�J��=��ݕ�b�k_鿍��0�#"���(N0���]\�)r9��=][�(�Vbu�b�{���u�ٮ=�2D�*>*�^��{W�\*��f�к���<@ܭ)���E��~��v�t9[m�J$CR8\l��L���)�	/(��΋����x9� qzɍn��mk.�s�K"��;B�ڔf8�n/D�vK�t&�S��ܷ���oC7�a� [{z���u�fSG����t����z��y7�j�!��B}6Ϛ��|���W���#���۾��CNd�k�!�P��!��7y�j�'^,��%t�J��6řxV7�:=���-��p"�{�Y�@Ծ@�Z�q�D����ʢ�ʽ�SǭIM]5������5mY'c���0�06��L�<͜T�qP�hf{٨{���t����[H�d��X/ �mꂨ�^ӎ���i�3�O�����)�����Jg��V���Q}w=1�.��s'8�v�X��Jb5�P����2���ׅV���`�T'�Z�~��)��Z��$�����~y��n��|5�C������
.��TL�2KH�J�Y3�qe��B����SoS��9�Ǳ���gx�`��hN������|u|E��>�D���X	���@���ǃF�����=��-���ώ������	M�v�6vf��(0`�Ltjp4K�����5�5�=V��}��U��{�n8����._l�ʉ�h��#��v�m)��f�y,CMm����k��@�v߀D!�oM�ӷ����TK�:Pʼ�����N��X|rQ���5pY#T�b���P;dݴZ�Y�v��1�ͬ{��x���7��o�wD��>ŷ���T��tH��-�
�,t\�:��Y�{YTG�a��*p�y��mN���#� Ȑ]��|Cm���7�>���1cS���@�Ƌz3��5-��m�����-SK��5F�^��r�C��xD���k`;s$;@���~Ny���ўj��*�p7�4�C���No=�y{�N7��'��,�eb�@28ȡ��4���šz��&TUЬ{�z�W�����G6�M��Qvz��������l4�3mP�N�?�[��l*���b�s�U�����H�r�0c��_8OhU�=ֲ�Rː�;�p��X
l�%�x�kd�t�+�x���׏���>j�h��t_�þ���NULK��>0�B��0��c{!כ5�*5�70D�.y�X���Gz���<���ᖭ��a���k�Ky2aa��w%4�����8~58��-�M6U�?_���`��q��|��/C��@���>�%^Wʶ\W?�qr�)����J�n2�·0\��[N��o��xg}�����	5G�.#H�*E)���hA1�ܜ���s>��mR���))���� Xz����}�a����]_o����k�Nq̹\s^7{K�Q��I�NA9,���ڧ��݀蚽�������K�6B����x�`dN��M����}p���i�LLͣVM�6	�Ph��|-���Dkv7�02N�nH��x� (�?/�y�O�!_j�D�� m�w��R�o��W�Z/������u҄�ӷYݰ|��V� �<; e���lLh,k���^}��^�r��B !��{��{��-�w��~*B��wy[�^��HRZy�`���	�`'�wϔ�E�6�H��և���0�ŨK�a}�V����t���yF4��!�[[x��(��y;�r�;;'�:�=����q0��N3��6f�������~B{������}����a��\;���R���MUÁ@��v{2����VJ	���=:U��ri��z׉���N��Ydvwӵ���/�x�;�|d}��`/	i6	MjN
��Va�gd
�oW}���+����L��W�� �	��&-�^O��7}ꆯt�vE�k�v�3�7�1��VZ��u�=x���Y�n��g2W�-��VA�H��|�Tz��|�-��y�Wsb�p�5+m/k�Ά��Ӭ���M6_�T�	�������{�m?V��:Q~��><V�o<�~�ͬSK-�+�=�~ݙ��|�콛d�eeSm��)ln��3�2��{g�^W����ނUm.�0��NγN�1�^��qR���5���pO
��N�
|Ά�N�5����:��J���5�^�=��Ss6�[�V�]���˽�%�3�*�@����e�م۶�7�:yN�y9�Y�x]jK�:�o�x�rY�ev ��8�Y�wE�s�Z�K��Se T�=ߊ�hi���h��b(����b�W���=���E�v�o��R�`)�w8��T��(LM�T/hZ�a��a�'~���kf㌹�����6TC�?�c���^.��n9��lJ5���!��"�j �4l����vu��c�4���["�(wM˰�n�}M�]s�����,�c
2�nC����r�RW��;%{��~�����/�d��D8�x�>0�e��n֦�OL����O<G3�����ks�'^3q*��^���z���(�dq��Ɗl���p%���xD=�z�g�^[�d?<��U9�B�4ޑU��L�+�u�=Y���&y��=����������'�e�]qy��͕�2�2g�r�%��ҟ#L�7s�qd�j��MV��h//��6f��ڮ��d�����f�;�g�wh��#���t�K���P�T��N�i����Wi��OժY{ñ����L���"{b`�?�F��T�_V2p�����-�0��$�X�@��P�J�^����S^m���u�9��%��K�R�X��i3�kK9��6#:$ἔ��ù't!����t���л���Y���TY�c��ʷ!Kwv�ۗ�9�O�-����r���<��yp?QK�&[Ϯ��}�B�|m2�i7,(AH�>������z�~�Y!0H�^7�H�ӆ����-�|����M<h|2"D���~O�C�L6�,�M�u�r"󯆦d2z_א,s�ly%��IWA�q��L&�����&y�����Ԏe�1E�^�v}qw�jq�^˴z�z�0�mdK]j�wyͻ��L>9�D{�q]�DJ�60J�g���yP1Df\
��,S���҅nc����ET��Sl%�,���M����n�CQ��b�� Ϭ�-��󘖪PS�*GH���;�2�v�7>Q�5]�=������5�M��z�|>���H�H�o�Ϙ�vo��Nn�8ɨ�#����;�e������X��x�}yB�NNC�c��Ǹ���o�2;�g��f���:��ǉ��Iv�v���v1��C�S.~���l�9co�L��aҁ+,����������/��3O�ﾗ��jN��e��$ʨ��x����娘��X!����b�'�5G6�R��P��_b���'�ً��0�]�����x~p�ތq���r��F�n.7�ڭa}IyZhL��[�[a����@��~I�(<�{�������E�9݆�n���G+��D��Z������j�qX���:�Όf�~��_J�� �}�;���`��Z���Yҝ�2���������x雊�]�6��7��iN(A����K��fWL��k���5=����<�<��`Ql���1�s�o��H��.���hػ�)0�M��z�(��0� ����l�K\N�T�Ua/J�S/f&^�gL�9�/�j|��R"���A"��Ȥ�}���<יgf�Q|1Վ��@�禄�0� ����8q����#<��}B�3�������in�q��u���Ak�3���j�H&�����f��ͯAё1���K�|`T�4E�J�^r�j9������-b�W��+���䩚����-r���ؖxsYgd#>�}�L.+��5<��W��/@c�=4��v�~O����K@���� q�hO]0 sH?� ?x��v��V3�]�߅���D#?~c�NϾ�c������ܡ�%�c�i�p厜1w%���}W��mі;P���a0�[bY�(N��Sȗ�k�6�%L���	�A2W��jڮ�f����l�����U�#�֑7�)� �󶙀%f���Q�ϼO�~�s��4��Z��
Y˻�J��]yz�ܗ��=8���Ve����qٳ������m!���	��樼�����4+���`ůq�u��n��ں��Wዐ����˧?"�O[I^��u��G�EYE�"����A���+~7��|�v�[ui�>��`������{���b����-�u�QK�SG�cY2�1U��XuQsoq����{AC�x���;Rsc��f)��`~/�I�,�
�d^�z�� [8�|�Y�yn�i����t��{�*�yn�X�4ݑ#z �(�W@:a����SM��Sm~�3�����m�y'u,d:g��2yy� 5�=.�}O�[o�4]g;��c���맓��O͉���V��u����\;�Zʮh�}}hN���˩O5y�xaJ�"�ݮN��� ժz�z'���wv��ܙ��F����Z�.�������^c�+�����]Hv_�C}��:;�LV�bW�7����Y(i��:6����kϣale�`�ؘ�XXoĢ������[e�j�L;k'�����f����ͳq
��{ѭ�c[UY�3Q=���-r��v����}�1�]�uT�L���L^'<��0�|�~��~���3����oFO��c�8�D�f��M��)��DvY�P�C��
��2�.޶���j���[����=#L0�f�E��Pha96���6*��=w�3ɚ5�3��ӶJ>�c-��O5Kי5�f�#2��fF��eŦ���Ƞ��]���}u�4�;� ��=�W��!=vyl�Oq�8
ɢ�4�V��<�t�pW�4A:���&�B�\/a�e�g�-��nS���]Wi���B镣�L|�.����G%WχO^��|����w>���ea��TA�` ���))ˍ�%��:�|z��g'���&g���yT�g����]�E�gv�+Q�������E�BJ]�i�g���]?�r'~�15ElQ����qz%�t�OK��Z8��߲����^ޒͮK�V��a����zw��ba��7����SX};hkHcfS��=�C��^�&��M��bY2*�[
�V�;�yك.�j�Y�N�w���k0�J	�K���1���A�>�E�ZfӜ[$��{�U��I��J��f~Ӯ��C�K�S(F]�\z85B�`���?J�]'�'�>�B��&	S������|Ѹ��2K'!�lz�[
�S�s�h�f����5)��kw�7�n��^/uw?N�[Z���9P֑D�z�6�쁖!��>p�`�k� ���ŧ��Ұ��0Ț[	ﻏ�/l��6�����C���Ý�XkH|�e�xV�C&�+wW��.��E��DϠ���닝羨L��]=α��,g�θ;;�v�>0oz�{� x@tsD�))�J��(���&��Z���e2���3z����q���"��pa�Y��9�YB�P.���,�m&+%jC����|�/n�N�bY|��<�ɗ|�K,gצo'�	w�R{�r|�a����'Z�|��cRm�ɾ$T�{�h�{};-4	��ti�D�TGQ�`�:�r�����,���]WhEƠ9�l��
Ff��v�W�H��WP	uݑ5�"Բ�0�[W�{/u_v
|ii�{-7[���w�! ^up���Y�,1�{�ue�y�Vue�]J|7��Uo�L%���ﶶ��ݳz1�ə�U�]�,�3a���`��0]Ojh��Ti.��P�J�B3�^�,��w�w�bV�4զ�!l쇸a��R�؂�j�&�`av�W�Q�k]]��[��MÜǒf���S��ɵ��[�OS�о��d�i��\t���h�v{��`\�k��l1)����l<y��N��m�j��|�ሑ{��{�"�k��gL���G�v����2S���6�30n˗�ݑG9�[W��	na�+�$�~l['˦[�s�k���"��	�[�<�g��]���vCXj���o7�y�xvP޶:�ɕ��o�q+W.��������/�b4uNt`�;.��j��-wC麚�7��x�{��v�}Ԗ�L��z+�e#��n���7!	
�4O�n���Ici8r-�6�LK��J����#��H�z�G/"���] G��lc�a]�?y�/�_��������V.޺��L(���K}r)� f���ж�*"x*�[g�&�+k36\�3� �ɍ�P���FUʮUR�Q��յ��:bU��or�]�FB%>�i1׉��%]���r�w �.�m�|��å��gMDG�� �U��T+.����g�]ʻy�ҳ��N�}ץ	I��F�B�]K�pT���W�O�,��J��B?��Y�Q�]���t<�'�S[U���2!�]hE���q�����&R���:�|g�S]�Ը��]۽�Km7����(�`{�9�5&6QM���W}اrn��̝U}1],�U�嶻61��o����WfWX(�������YF�@�BI1�_dT���.�]�f���l�o���Ġ�X+:&	��;�cN\ �+r��;�dV��5�]H���·+����ݸ���B;tP��Wv�\wEQ�o��$��nrCՏ)]��10�{
�n�\������\<n%�.���k'#۳gMݾp˻k�v�Y�U�,WJܬ{����8���E�F�7��ʌ���S[Y�ة ݋;U����* Ұmբ�rt�q�󩕀v
���8�V��.�v��B�Xh���7c1p�[W:��ѷ��jul��o�]e��z�9*���n��Ur��X�I�� �	��C.32'3������AAF�1��L"�arNs)��h�7��q�Oׯ��<|����ӽ����AQ�.A�DC5&VfY?g7�1�*2�F�EQf/��x�<~��������ǣׯ�3��yW���Y�1(��*`��0����z������w��6�
��3�������}��O���z���~��}̨��V�f.[m���UfM5��9da6b��|��=�f��c��2���f�PT�SQ7p�b�j�,�*�g$�$���#ȩ*���cPl��PUUG�ɪ�pt�"�h��(�m� *�0ʒ"�&
Jb2p2$���()���̤ṶTRRQNYRS��DE7��s�l��*�2Zr�̬��0����0
��J���,��U�a�Ctl
�¢
(��(�%�0�3&�H�*�*�����G�,#��bg��	��H`b0�i�)��>�$@�B8�p�����^�bi|�������Z�w�����tˡ�o��]��1�T��z����ї���=2,u�����`��t�'�e@P&y�Qa¢q�D�DI�£n4�jI
d"� �l��a�jH�NH�L�r[IE��qG�$��9"$[�!3s�6�� ~@�U�A��xx�x{ƄA)��a[��U��$��E~i�%d���O�J�yO��)�@�2*���@ok������g�	!����R�&_�ԙ��M.�u��3w�:g���2�@�cZS�r�;�Qq�	��,���Z*��ʡ&'y�D��TZ�R��t5�74dC3�b�Հ��u`?7����*��r��C�;�N�6u\�O%L�Zb�ah��־�?�_�[`�O�(T0�x�@�*E�'�5�>�g7�b�w�h�^J��KFk��#0X�t�9��M�� ���|(#�@<?�G�O��&���҃���T;O�vx��Y�͎K=�g���*g�<��S^��y{2(��ԼgȘM���J8�^��koS�e�dP�J�k����w�{�A�F��
��q"�q��^�^��ȧ}����zaa[���
�қ�D���Uk
n�ڛ�}Yt��w\�hg����җé��f�]�z/��~�J.w�y޵�5��Lyμ����,���¬{�7ڑy�5qhY1v���ۆ�ǩ��ѵ��]ħ,�*q�V�H�w��v�n�����A�3HVE��]&�*ã��2_higx�X%�����Q�D���g�#�,K�q,�łY^$"<O�+����pug��{v��Q�G���֞�l�!)�[ԁ��'Pc]:ι/�GG˖_{N�e͋����� #
�Ȥ0 ���Ue��}�)�&��5�׭fP��NCվ8)�=���8�!�~��C5{�rjZ�*�z��۾C�oeZ�e��<���"��=���f�2#�T�55�t�]�O!�6�����}��Ն�t-�_z�z�'&ۋ>{��7d��:�G4�ػ|��kiҰ�wS��c�an�ͨL��CKȴdH�\Jy�d�Lc�rضֈ�~���V��7�{5�D>�#���	k�{(?k��
�j�/�Xzc���K�[�koog�#^O��z�ȍ�|j|hD������:�/��%唈���x�����}5~����}ү�ԕII$�m�}�@fuP֒b��v�/Z��<��`ᵯ��'��M�V�<�d��tY��8A(Mt��>�U"A6%ۻ�30��������	Sy�^�U�|�b�}=����i�����f��]�;^���zy�'���?;�����d�?g�?A����N��h�d��C��B������]��4�fG���-�`X��4�3mr�}�C;SY5�z�[\3T�������_���x�[��L�GQ��[��Q
�Iaw�೺��X(;��~�~����4��p}����Yy��4n�$zu%�uךka�#���I,�}�kT�6u�K۱�&FSs.���rE�S�o�Xҵ
���� G�A:��<�\>�<�����?9��s���SQg#%�:�Ch��,a�'A���Zf���~�97�U�scø}50��ϡ�m��Z�b��ﮠs\�Sm�-L��"`��CD|8�G<�*�>�y�,!+)m7� ��o,՛7�gŭ�C�j�`tT{[�1x�~��.��<K 9Csϩ��JobWt(���C�۳.P%v��Tl���W�u���Y�_@���ƾ��2�8I?
�}�1�2|D1�%2ɽ��T��X½�g# _�"���6E�2��Wmu�oKG2@�De���������ѡ�$�aig���QUm�#%���1��o����=�ۅ-���m����x��F]�&��W�/�C��+�7���b�I񗊂���&Rw�N������A��x���]/̂�	����R~�AG��{��&J�q��F�����V��Puv����V�����`9�s���u�	�a LBm��m�jD��a[�r�͍�x����j���E@��T'c� e�l�������n.�4�=��qډ����m�L��y�M��i��
=t��O*Y,<�H��O���w�x�:�W|��^�^�	!�5ɯ/W���=�����k��#&�&�_v�6��I��v�����osK9���#*�$0+� Tc�{����fja(
ho�#4�7zFvF�*7��C�����FD=~Ky��}�_N����S"v �:ie��,��=s�li��+�O�tv��{���h7�]u�wxc���<�=۲I�Ѳ����C:��'�.(*0�|d�dh�m�����.0�3Eۖ��`���0�ysU(>�?���8��"�\�^�}��Y�h������=�8?��pˁ����U�e�?�-W�U����(��xu��_f�|�Н6����r���a� fC�Sv��}�I{j�u;$�CmyS0v���)�] �U�D��15O+b��|�^��޹�O��ڴ����a
5P�4�:<I5�gN�R�}��0���J����u���^�y�}�7�b��$f���&'�.��=�M�fB�-y1,�,��m��Fڛ����/�����8��9q$m���W��^w�qZ�[#�s�Ǯ�M^]E''5P��jٛz�/��{������Z-��c��T�2&�?��[�MmP��H�M�0��;�W��R�)�wf�lc���ߙY}��Y�Iv���?�4����.H�+����~�Wg�H�5Z/N[�}�i�5�VH��G}Z��bځ�;K-��gN���Q-���V⃆��X�	B������y]�`*��<���ȴ��|�U�Y����?{��H`F��U>���_5�<���o���-m�ծ���I	Bx��iE	F�>l�
���$~
��>�a�\�_����Tь"��Hs�h\s4_Hf�Je���Kj��1ڰ����4�V�
"���45�����5����/��@���.CsH�ɛ���0{3s��vk�v@��>�S���1�)���GF����S�b�k��TO�N��1Ng�4D$H/�aCC$J{��5�� �~ʂɸ$d�X�|��[9��ٚ�B����T�d/�հ^q���_�EJ��r�|���zy�Wd���=;>��9�,�,�o�*�s{��v�Ey�����@�1�HeŨ��+�ϣL�݄�gx�M4vA��aT�h�*7a�ow��?3ߕ��~�4�I� *�>�0��UǑ�x�CHӒ3Z�A�U�Nv�l��@�t9F��fja�Ϝ��pz���"�_+�|~�M��Q��ai�u�Ʌ��uV��<�r�ֽ�]�@��L.b���<�駈�k �`EʛaX���m��L��q�ZpsM�ޞ�vX�N��U.�1���PY�����P!�q��U�>gQ:���e�U�Ahds�7]>!����wu���,��mC��= ]�gU�[K��<��������=����6�����B�IG�#f�P�I�B��	�?f�'o
��b#.�n��t�%�n��jz�U��d�jߧ�}��P_��� XT &��D�^��sx��z��븖��K�]�1��a�&D�֩�o;HFm��zN̾*�r�ױ �ǎ4�4�����:�`Lgd
��SȨ�S	�P���P��fmt+�R��
/ݗ#����
e�Y0���.S��|�����u�~���Lv��٦"�LӜ��&����)�i�մ��+hj1v��[��&��3�{d�v%�nf���VT�elCݸ
�h���u:������P#̻�P�z5r\\:��v�SO�2B,��2����/�j2�����g�@e�P��7^���O|b�s�Q��G,m�S���*��Q����Ƹ���V_C�C�Bƒ���6��r�d�y�)����_T�����m�+\9~hl,�Q؟T��3��M��O��������yǑhȾ~.6	qj���d���
��ڞ`�1���\�4x�_���?=?�\���}ʮ���ߨw���q�6a?\5���M��[�Ǩcծܻ7��)Ťd����i�,ͽ�|����{�@H�ߕ�����vs�B����u��ukU�P���`��?��y�y���/`3���0�@���Qn�Y��df.���f��u��4�y�	���s�Ӧ����{=0mG��&��ա%�0J��j�Q��.�SJ'+tܬ���},�5N��|!? � ~�
�0
C��;���w�w�~f}B�
�,�j�hkO���_��掖q�o�u����:abC�_-��QW{	�S^s\oYƖP����������6Ù��lK�W�@f��ͯN��գo��{r�C������#��%��'e��ۗWv����p�������^�,1ݭ��	w����W�?ke��A��D?�$��r|fǖ�f�����Ŭ�ZA
�`�ձ���]� z��l7dD�	��~Ӕ�����	gl�'�_}�&��E��:܇h��0�9B����R�MΞ�fNΛy�#Sn��ja������ |h���TB�]z����
�UL��,vM�o���i�rp^�M�\~�;�X�o�`Ϗ����%f�� ܢ��ĵ'w5�0�L��=��ڮ��ˢ���a��Ȗ[iV���Y�-Ț>�d�� �ڞ	Q���x�����0f�u#��h�����En�49�0���_�
�d_ש�R���ٙ�"`U�En�|�H@7���v�*�/DۯX�4["F���{�%�J�����-����y�v\<(F�x�eڶ^]t��A-�p]	�3s%j�QS���&�3x/���B���5���z��Xw�;z.�3{��[��Pm>>9z+�e�����(��/�tgv�'�oP�3��#���c#�0�3i�\�.p�h�ר�gv�U+�o�*�=�����2�� ��OǞ�_���ǷJ�S\?��ڃ[BqK���!.�W5�@z�*\w��.�Y�.c��-����c��V6"�q�X5�@��4x�����{���Mı�T������Ȃ)څ9w�V��9,��6;�{��B���e�۔���8����Ѱ2ָ4��$DBm멖�f���%tʫ�Y�o�dAi�8�eE�^��68б�|3U�f����@{"aG�P���6�Y�[wG�顡�<�M2~��C���2�t����2�� ��1�r���{�.����F��`�<D&��z�M��zoz��Py��U]��zy�x��q��͋�C�5��OՇd2��yݹ��9�í0 '�����W��[�u�5���1ǣ��'�uk�y	�Es�6��m�%�@�X,�/�W�B���!��b'���f�졳7J����c����-�{�����!K���Q-3�3���2%)�x{nY����5�5K�ToJ�D^�̆��p�t�^&]�����=x�|�"s��
jXB���۔]�8���B��w���Z�]6K��H+��V�_=d���c�{%�7T����A������+���ܲ*P�N#�+��.]q��򶸌�u㊴��=vf+��	])fn��X�C�扼{z�!�bysk{��� {��x���`*�~<�{�gs�<}�|���h�����@�)�HH"$�H�M�R	}��-�������a3c�ĵ��T<��c"y���<zݝ����l�#i�S��C��L��p�P9�p!l+|�A�R�D�lEmSu�r�b���Sk�齬��6�3���H=)b��Ԅ��?_lC����2簴��c�l�/Y�ڦc��3cs�a��B�Cږ�ي)��].��~��1Gs��R��n{�Uq稛���0�/���!yH���a��������l+�T�C�d�^���%���W\�g(
����5c ����u@�2�׆t܇l=�>0�P��K�g权�7��elF���]
Z#�+6D�ԮrY��ڥ��܄�Шp�k�w���$vd;= ���+U�7��r˨�	�j���7��.U��b�Ί�g�xm�`�D��q�����Gsh�m��L������T��E?/�WK��E^���#kϩ�a��� sF)\z��3�F�o<7���>�������@hg��\j1^��z]=�;�S���4�ÙKo}�,�ވ���ۜ`�+n¤<E����:�ԓ�J�#[]b�y���-F��ȓ`�۝U��O0��i眻ǞLd�3'�*R_	u���9�+�o^�F�a�*���%ʳƦ{w_r*$^�$f�E�հ�gUL|��sPK��Fi��� ���� O���=���<=�y��xx{_)�֥L_ ���`�	f|�A�J�W�o�1g�AտW�<���c��msЦ�o����}!{�+zF9�љ�⃛���ͥ�6Ǣ�@v|z�ɕ۷��"�:����ө�EO����g��x���U�_��r{:Po��,��e���Y�{7++�X� �f���Gva�ͥ�7�T;@��E���f�%�̓
˟3���XE���d �3�Һ�.�T�'ۑ>��^�/V�����fqY�=P�j0"ӟ� �����!�?/		3��_���_(D{#ͪETE��
��zi`�Ey\l����a2t�mn�7ǘu*��g}c{UB�A"Y`g�g��qk��S�4t5��?'�薪PS�eH�gMLي95-�C��*���onD�x���uI���ݑ�
�..���0��L��i��z}�>�j����&���E�d��[1��������	2o����Oΰ��&�ؼz�(W���z��)�=Ǆ�8� �	xT�N��5�=M6A��@��$3^�/SS�� �����S�n���؇`�� ��x
��n%�Do4n����YI/d�;۳^8�i���gS�X�z&��M
ȟl�E:���3Ů�o��7�̽$����ζL�`�y3Ɩ��T.�Pk�����v��ڝ�%޴X�:��wr��ת��#�i<͹D,G8���c4�F����Cs��}��a����[��m+����(ɸ.��XhU@2�Yf�WM��׹�R��ׄ�g'2W3u0���F^�͹�݉�D�x;���7J�[V+�*�����[wa-�t�]����-b:MwI�����vЮ�dM�[ݙPi5��!��I4��]0��e�w�y��F�e�]	�ٵܫ�Y�Ɵ�dSG�o^�p��X8^<zq�'��5�\�%��*�j�O`U�H�U���\�Ѩs\�Oe���ԝV�U���ξ\��˰���<2c�L�v�Z�f@E]:��J�;{
-�c������+=��q���.��ҴvT��yA�n�7������i�e͆_U�U��7���wv.��gZ/��{/����|�v9�5g��k���S9WA���w,<����q[K�j�2-f�]n����I�uW��К���%=�8�s���bb�sh3��1���{�{�n�Dr�;X0V�i���s���VO'�v�+)�M�d+�+�Y���3{l���$7SV�zW[�׻VǆH�5r�/���'�s-W/!S2<��X���ψMeĲ紾^�&�t�<��e+�����R4��w�r!c9>˧��+YɌ����|���.և���Z���I⳷H�SC�X�S��6�VMw����5�l��]�)�5��Q*ef��ξ�ʎ�>�O�1�٩x��3v�7�b4 ���mf;�U됎F��ɵ��Ρ�Q�!�g�*ʥm�����%tR+4��>�Vh�N��A��@#�~sjR��f�)�D������U�^��uLK�ܸG��W{{D�f�Ʌ�A��[�qsq�P!s�8��'�P��Հ����Hi�O�3�۽}{Z�Y��'�!�&���m\�-�J}�M�@�٘�ޙ���_d���+�ЦN3�]�&U��'fj�D�Ծ��l�z�������L�Jd�t7�H.�&�Rݤ.3f��C�4޲x)�:�p a�e���.���6��}%�GՔys+����R\gggG�_vj� �f����mm��Ue	�f1����]-�s;;��˃כ�n��=ָ�SxH�A	z&]�+_��I�xUX���到n�G���&��S�%6n�n��V$���.��4���!�	h�X�m�O��skV����u�;���a<��6$9X�[��R���_q��I�zĳr]��$���K�����3	��E��UFa�ՖIQ=�����/��q�x�||~>�O��������~��
J�*��c����,�1���Ȫ�3,(#��8��O�������}?Gǯ�3�C4Q@vʚr�*���*"�2�r���>3��q�����}��O��������Eaa�PL��S5UL���!B�Y��FYVDddzp65!�I���LQ9d��I�YdQT=��a�� �dnd�MSQ��[!��p��«0ʒ+X���3&� �h(j��³2f� �))*�����Ĉ��˔�eFES�LYc�SKMeՃJ����RSL���$V!bQ0P3*v�r�)�(2L��f>f:{ͭ���fe��T�M[����M&��9Y�M|��rL�1�+/�>�]G:��OIj�{�%_��^k<��ֲ��7���Ƈǐ)����h�Hv:ܩ�w�݅S�'e������~FDe=���0A� ���{Y��rz��z��L�<��I��-���M�_��m)\��S���t��j{-SDyקbu��+�<kmL��^ǔ򱌋�\p4��Q]<ܸ���J]8��'�j���iv�@[�-�R�wQ#33�~i��~������g���
��x�ͬ�T��ꬸ���5F�J;�q�T��S�Y�{^�������j��OYQL�uKꉚ{�|�6�E���6hT��"_���c�\���1������g�׀�|_�$h��oD����f2��Ɂ�1�㬛VՋ&�3��X|��P�]q�gׯU ��λ*�xn��˄)�o=Gh��_�s_�y�x�?����g��0�Bߑ�f�/���c6���\�8�Ȅ�i�nk����WA�xǤ"<m��q2 �#]��]ö�}nz��	i;;3����,=]ww[�)`˔�@��^]�Z�H�%@�{o|���k�cQ����S��_=��يCQ���6��~�dM��IÁy|a�u��qx(�<�P����;������NŮf7>�S�b�^�1�ԵͰ��t��[�;����ndQ�3]	�j�}uN�s2N1t��P��=�Ֆ
c�J/����=]�(ud���6�l7����o����38�_����� {�����)�Р��9�|�����|�s:"�3zAm�$Kz�U�U����+6g�},ך����=�*����w̍��^��}�;�V�;T�w�Ȗ�ԫw��Ve���i��[�.vk��鶳|�B�3z�w�g��0������d*��{�S-Je�9��Iec�����M�7�*�um�{�A�<��d[��Z����l�S8j-�k�/4�S	�J�m�1S�&�xھ8�j���l���ڤ3�@�R�$�	���M}�T-q���<^�5CWx���),�V���=�[j�_�u��^U�/`���.���z^E�1�R�o)���<�,K��:�W1�n�#ON�J#�u����TcsP/��2�ָ4&�0i��=	���ʹ�f4�b�	��s�ҡ�R%�69��P��m��j��Q�X�ٲ��[!��t�u%�66�z`ݼ4s�R�����������ޠ,��yި��-r�^����mtә�=&�Mw��ed��\�%�azǤ�S�r|����v�{Ϊ���X��j���Q�i�qdw�)zg��u�Y㷔xJ�:Rr�����p�·Bqn��Ur�bm����#��z)v�S�;��-Q.��F9���xPɒ�Cgb��?��k���r7�ux�Q*��x6'!���N�+n�ح㼖.j8���;�<<=�H�$��@�y�g�-�"o�U��7�ƊEF·0��,��R(�m`��L���:��3t�����
3��>1���p�������}̂�q�o���a�E�h�PL�g������|�l h>�0�d8���[�x�l�i̭@�� �ٹ
�.1��TC�<���^J������;?��@����Nz�U��ח������g||V�m=�&]�M�ܮ�?3��V�	ן=�����[xĳ罪�N4�.�멨�Mt�A^+�b�Ǻe3k׹D��v�ND�oV�]��(;�P��:���e1zGTd�x]z`7��P O)X��1n�ɳ�̶hK(W�gD�f�Yf'�"�㶿F��?|�K��+�\n�(�_���M��vD�{�L��dR}��صWY�M�s�]����L]�2][r��/v1y�z<ZZ��C�z߃R|a~��+X5[�13����ٛW�=�[�ff�fgպ�n7ƅ��N0�F���Ǩ5��aQ~`����1��*�CN���iU9�A�̄��['�� ]�>bR1����k}�!���#&�:	� Kq;x�[�_�[w)t��4��Fqo%ʡ�clT���J��OM���*ݮ�����vC��M�i�r��릵G9��^9��52vJ@��r�={������+*[ũB�t�r�O��:�����d �D|XW�#�^�������M"�K��}�$wT�s�/Hň���H�Ϛ���x�i��^,_Y[۔�9l�h*�M��2��N1YR$����ϼ��˔Ɋ0Y�|ޏ,i��u�˖B�+�l��*�vN�=�ИHy�4'E�S�@�2*��y�Wgs0kv��X����V�REѓnn���s�����䬖0Xw��B\y���q@fG%�O�+�z�uWd��ˠ>O�V6��~c>w���d}.�!�W�
�����ǊS�b&DP{׾��кN Y:WAr�o�ǣ�m3e���噴��mx��#"�ɂ٣(�͑:]�mgk�<C;ϥsj�fMױ���x�6����<dXi*��y�[:z��P�l<f��l��+�z�?a��~�Y(��R��c�J�����}%�\�=�`*���<�3p�So3kDø���^k0��L##��^�ŵ�ϛreS��0��cDȖ���mǍ�R��YGNnʇwA�q8m���u��G�#]���������oB�e%U���������G���@�h��w;��B�f�8GY�Չb�S�R���f���S�(|���*صy��]��slϪA��˶�NM]���ݱ�}%�ᇷ�Ҙq��h&1�*��j�E�27z��t�������G�Gr����߾�w��?#"�0� ��oxxa� �7� 6X��Q�����0f�"�CQ��r:��٭�7'���U>C����'nj�ǽR�V!���K�n��ؤ�x�����.��;�v�[z�[L?f�OT҈��q�V٩ܟ(f+�Z۟�wD�O�W�Y�b��ֳ(R9/�V��%�=ǃ�N�M�̹�wq�R��L���VH������&_a�>�:���S�V���b�"g��|#�����[�[P��t=�g/�yh��Z�%�2��-��d<�2�Ky��R[��T��t�����:Mj.��핦8�uV��p�
1�]�O��>������M��پ�OXn|$Y�.(j���r���|�;Y�t��5���u)��vt��6�,���~�r��|��_��8�
���	�p�ƻ�R�(a��y���)�Yݝ����R�H�S�^�m~�D����iz��N�;�/���~Yg�bs�R��5�0^��V7<8�9��g&F�1m�0m:Xfj�����<4U��x^'"��������]�/Oͱ�]�\��t�g�����lK�Pΐ���M)����l8ֿ�jmIضS��v�̇`ߗe5��h���v2j����lGRW����s(�zÎ��Jr�_{�u��}�V����.��a	t�CAm�4u���uZ���\�t�2�5��X����!��Tׂ�=��0��<#��>��!�XaE��ZUB�������;^��O�DT����Ի�g���)�5�6k8�{���T�۾�\ =.��R�����M���#���c�f
/�ʆ,�(?]\f]�i�c��ު�Fj���IS�=՜��E�p����A�3�_ʳ�&�(S��s!~_1bS����w5/(�����}��a��.k�@�����i��4��}u~�VSF�Rp�+���&o�U�\�jV��h;AM�v��OY��5L��
��(�	���m�וm}��!�ݑp��n3�y�K6n]��H�R ۶&��F7.�j�ff�̀j�R��<-��p��{h���%��ݛS�[y�!���ur�vnke��8-��@�1�s�a 2�wUL��)��m������4����kKe�n0��5�uq["y�\��<��k]��=y�$�aa*����r�S�8,�'/���d-kEN0\�;�֔j�s�.��:m�p_t��W8�t*s��L��]�w�j#/U�+^���r�m�+���4�+h��L:Zx�YꌐL?���܌�7��eMs�:�~�{t5��1�����5����/0R��1��Hi��k�ǹoKZ�<���]mпf�ϳ�� �P�ɹ[�,���m���L�տ�I�{x{������X��]��r�y�x��M��9gB�nc�T
�< � x<}�2X
DJ/�����g8�~���}��/��'��ȉ'qD�,��0%�e�"���YB($k�߂��]j�ox'�E�={�$F�2ϸ�����U]��ao�\��a�R���^Ș�Ϩ��P�(�Tr���5��R+\3fk�����ɥ��S��6�J�����ʢ���t�Δhg��
�u�U��5I.=:�8�˳�Ĝ#D�;\���?oƠ$�G�~[xJIo`X~t}d���5n*�O=cߕ�t��푑9J3y��2��w*�8��/U-��vǀ�͐lslFzB�/X��Vð������V�W=6��ǰ��e�7������ɚO��l40��v�^L� �s�]q�"~��"r�U�=�)���;7ck��-ne��pZ䖐D�7�׼����Q-3�3��%|���?�{���y��o����/�a7t�ֵb�ϱ��ڷ8ӵ{� �@�v�Q�=����9ٵ3�נ���l������2�7�6�D Q�M|0����?T�Dtzk�3�����b�8ĵ֠.�����̊�$:ju��ն��j��N��˻^:
��
7Q��.�a� �6�j��651,�,����l�1J[�PQX+WU��fo	�K����i4�nl��z�g<�=���Ż�%ޖ��v��� �}T���U��0�k�d���z�1��'En�4l�mĵIu��}��=G@p�a�x�D�{�ߛ����~G�+���)���{������N���nS�����9	���M�>���]~�/�>3�c;Å�ܽϾ<�g���u�ʊ����.U�i� T�l�g1���"�];���l��)f�[�jO� =��O��wf��Dh�u~���:����黏�W��U�/��������Hg�����W���2~�Q�������=�]�T�h��R�5�F���JF4��� 5��;�W`h�ahg=>𘽼�u;΄��Ml�0c���vK�;��fro�z�<�A�ֹH�� �;�v�<0{=|��gz̰���s�������Ld���x�-�L��,�y������|k�oz���h��Q���}�%;I������F�Լ��~�<��40'��tc:��早w�y��ɴh|�n�Hj�i��/��Yk`�(k���~6C��='��(N
�-A���v��s�C���VzW�:��M��q�=�3�>r�����~�=�����$?K��;C�}t�����>�CUר�Y�^�O��-���Xj/�̕�XiW�33�.����#��l��<ʻ��:\����'�u���7��D͗I������woVt꛸���<�~���W_^�j�+���F`�=��K ���n��bMqf��B�w_�v�!Dg_2J�{]w�m��N�>��^��>�9Q�Q��� ��������{��������P�3[f��n����.�`Xl*���t�У����5�����E安a�$����>"y�g+��2Uc�B��,��-��f�Q����U�
s�[9�[��;�2<ّ �T<�e#ZSܽۋj���[��u�X���6��Qhiȣ�=��]Q�KE!-|b��:)D��T"=���B�De�
��y���o��:�8�ʬ'/�d]��.�� ��PK��VF�써:�,xi*�����疩PS�P�7._��m�����K+��\��b���]c8��qU��aӐ��ƚ-�O�
a��8p�ZmF8Z���sP�R;��lҍy_�yl��y�{B���{lw�]��Ҥ�]9,�݅�Lz�Cw�ڄ:n�!�f4b������M�.u�{dJ7b��n-o�:�x���O>v���?��mס.�z�5��e0�Nz�[���-|~.�e[<|��UjƴT�8��~yg׻ȷq�%�7F4�_��8�hȟY�.?\���j��2�����X����.,]�����ŝ0�v"���ΣY�9*vJ���T��X&v����f�(�e�d�8S�Y]�a������_d��}E3�+U]��4-l��Q�6�Ap�K�֮[�#᎟9R��-N\�\�����W}|�����f=�X����d��f9�׶ֲ����?{Q>�ޚij�]t������6���P���-���B���qqc65=���X*K	Z�Z�.ͼ�7��~��<4y�iu�aYܱS��м�\5�Űy�<���R�)�l�􁋍�L�z1���&�����]�oK���m=/�
[:;k����@t�n.��Q�/���xwo��\��󶹛��Й��g�$�kS��9�����m"u|���眨D~XD�U�c������ƞ��1_�o@�vT���Ah��k��a$u�vS��-���jL�_��Y��x b�?{J�3߃�b�X,���ֶm�y�07�Q���%KA- �ئ�C�c	����T<�Hj��إ"%�U��a]p��cM�_�2����C2Ş�l��r{�H��������"����'O�<��~uا�+�3���媔[y'��&E��Bh�d&5�*Z��jƑ���e��!����	�j��Fm�n_4Λ���q-S�;g֫ɥ�T��,^�t�.��[�%Y�wබ�]=�1j[��Z��܊Ŏ�+�`�Z%�Vj�9��,�;��Y7X�[�|����,�JP>��:���a������/
��dR������)h�'j�]��G)����F����{\ik�[��'��x���Ol��i�&��H���0������N�m/������a�s����V��+iR+]5dݠ�튠
cReX���G*� �E�ڻ�G��ȉ�����	m�~Ok��w-�BU$�5�mR%��Op��\]�Q�ՙ��t�Ci�t���+^]�u"gJ8@��55e�ǆ*��CH���e��z`�+Q�J�p��j�֮��#�@��"7�vt��m���I=��10��"()�V��|ŭ�犳w6,Mu�t��{r�f�%���Iح�H4ruWT5Ҷ�%��4i��-.T��X�27q��u�P����3��Ӯ=g;y�#�1$����CNRAy\��]�:������iR�����@�:Eo�ɻ2{F�X�7(��t��H>�CWc��\+R��7 ���N孮�ȽxR�6�½C��2����4�[f�v�1����4;�=��}�]]ݴ��H���Y�@����Yj�F���p��{ז���4���J]�ϡ�#�=�[.�U��&L�Au�:I�J=��n�O<qSf�XT��/+%=�}Z`�]5�W*��N䜑޶'U��eМE�J�"�v_.9s��m]�dHM�lAʄp#���e����
%^M���Ը���z(d枚j�C}kZ_sI�%���.�v�h���2��E�P��M.�N@���P����:ƍ9lL����Ws�{��t�xg&h�a����庮���;�Ӷ9�' oJ��®�����|�l��s�8u۽�w�7�BHi���7:S֦�kEO�r��䧵�4�  �n�lݺMP��j4n�!��c�x�Yy�Ȭ��t;W4��X+�U-�|��l��r�4��s4��A����&F�
�7J뽾��;{�����d�ֳ��N��n;����|֎��I��g%�R�/
�a��5^SW�!Y�D�,\�'5T�7M|�At��K3c��Ll:I�Y|e��R���e�|f;�C�W6���J�U��-%�˓8kRDx	x�Çt�H�y�V�v�s���Hԥ��osWo!�]͐ѾW���;4�[����z�vF�7ƺ-y��*r�u��K;ǁyS��'5dX�P�-�9�X��G"�B��X�Pы�p�r4��ѫ����զ]����ֻ{�Ӻ�������9��:z=��B֜�4E�@��3���ፌ��֩u#Ƿ"e�楌�[�6����+��{ْ,����Ƒ���j�1R'S끔T�̫�dQT��e�Y�Q�m�,0ȡ��d��4ddf�=?�x�������~>�O��������=���.ٙ�E4����aSE4�������κ�~:��}?o����>>>8��W����QPUG�Ƴ0(��*���3"&�"���~:��ۯ�������}>_q�ڼ�0��i�Q1EAQF���(�����*�(�&#0�YTL�E�dTn4n�-LQ�Q_00`��Ȩ��T��&�`�"hna��Y5�3c"	����9��O,���AYD�ʶ��3	�a���)��3 ��UAUUs�&�� ���D�^�&�UED�fDPLPG,��2�,�2�=��QUP�,"(�j�=ޭ�Ȫf"�"*��*�
�
�0�"""��3��I�$�@�A!sE�TI�d)��0����)8�(�Bх%	 h6Q��<�ɷ��¬�D�73q+�:\�C3;��:�u;Դ>��*ԃ[����{B��<yM���3ו�A��9��-���S1��(��.%)�$	H�6��2@A%�؉��q�D"���l���Q�ȣ��@Ɖ��I�Ay&� C$Q��s�~����S%R� ��d7�H[p"W��Ʀ48�d��EIC$!��"a%  �����W���E�����~,]�m��|L�j[䪙��)�T��馎���d�뭾�����1�/��]�@�s-�@�Z��=�3O��W�P��x.�O8VѼ��I����V���Um�fq����ӯ�� ��)��zG���v[���v��L�!hl�]���G�6>F)>4�m���~kU� �-:އ���'֎v׃��DO+��9���{��B�&<��.7�����N�ִ7Inװ���C�0N�0�����uߣ?q�Op�cK�s#
�(���,���dKO�-���p�BO�� �0 ,i���!����m�T�aձ�7�}:vP���Ș0��߽�	����3�����Ƅ��3I&u�Uϵ���W̱�ZPC]�s&C�	�׈��@nl/6��}��W��wO���(�m�t�����)��&:g�mKC����ٰ',(C�0*B��Xw����乒�n礎�2��]e�Q�H�3E��,�؇l,��c�8y^zY�]y�DP n��B���.������sN1�F3�,Q�R&�˭�ᢝ�וPǶ#��y��b�Cɝ�(
��<ha�@���3�N鸶����tT�+v3������PT�t���a�;>#x)Y��8K~��6���m�=� dx�<U�I��|��;ߦ|������|�>��o�m��M�8���ӊ�O��Ӂ&r U�+�,��J�_]_�Nj|Yu�-��H�k�v�JE�Q�a�>*�ey�
ʋz�ڲI��2��y:�y��k�^~�l��MG�EE0�1�Ά/u&mt^�r�v|t%԰[��]��~���~��?S{��Փ�1�j�^o|���zV�Dhb�f�鲙���5=o5�k���=ʦ��T�8Μ�����>$���퐀R���>.����9
�KYO4��B��w��Ӱ�k�5גx���0%��9�m�aڭݗg�<�SmPT���pm�U��2����o�CJ B��i��qUt���>ײ�161T5����\?x�j3�*=0:��6��8h�Ͱ�Ud�Zk}Y	�</�<;8�gZ�`r1f")F��|Y��v!�r&jge������ڍ@�����S���-�MoK��_);�W9�ǒ1b:5��;b�lnlsTIGe���΄=�����K�w<K���"c}(�.�y��2b�u~��,Ix��g�c�c�A����3x�ssb�����M�w����z����3S�=�̺��|X�lYֻV�ĝ���J�s�I{�8�E-����u�05.�Rs��N�>6��6b\�-E�_`uo�t���jsy*n��L���]���싱�x���<|!B>}�����<�~3�~}�������U��"���?������O�g��` �S��W0�7[���Q�p�]:��t<�O��Jz]�C��x;>F���a�1NW�ѣ@�1�)����s�ѥj��������o/؅�����a�x�����cA|f����́����"7�^����Fg*��z&<��P֐�r�{����f��-�9�/OC��ۛʢ*�{���X��3T���'�����~��o�W�Xz�F����G�Kl�}�.XXlT��9�gO���<�˃D��kV�� M)g@��MQ��}���-7���S�krY�2�F�;�1�<��`��A�)�|���`�b���"M���?Z
��[P�/j��=~`�0ˁi:\ѽ�9?7JJFD�R�w�L۸�ꗇ4��T������^}OL4���(l(����˶I�A9�?s͘M�WB��7�SV+����v�Y�s�$��/Z��V_��w&~|oQ3�h˯c�t&'Z���-z�Ȥ�c�߾whV��������6a��ls�(�[~�O�0�~Q�W�X�wَ� 7�%�ˠ� u~־���ݶw:���h��^�e��v�[Zտg�������s�O���e>�s��z�wG�jp��)ް���rfn�S��2������|3�o����s]��x���0�9R��w���7jwJ{Υ����c�;<��M�7�� ��O�T�~İf����)+�+'y�b�	�"q	���F�e��c;r}�1��(:��3��^�s��>��_|>���+�s���b=�J<����~ky�>����P7�fD��x�?j��_;ҘO��Kq��M���g=Ky��)S_�ڭJ�5:�hg��wa�+�.�O����"n+�wj<CJ[հx��<� U��`�(9�"}�Κ���вG�a�M�/���h�k��*,S���{�]'҅�B�n�<\P9�*��1Q���PX-j�l.ͽ#ɍ��v��-C�Wp]����;�-��LG'��~x�O���7�˚��,0CK{=��Y�y��Tk�<�bc�p�L��C�	��k칦I�	g�z��N/ݝ%��3�����m>�]>�����F����L�ɯ����?, �������Y�(K��?�r����K{��M�yfr�Ʈ����xg���@bdD�T�qS�S�;c���vq�z;�8����z�Z�V��c緩����/F;�v�.L��F���V \�s�/ԩ�yc��˽���E�X��k�������3w'�\m�Ba�(�M�6Q*9GA��q�>���߾��#�3��SM O���}Eb��J?M��|7���y.O�q��",`CS-�K��Y���?qc��%�g~�_ʇ@�m��H�E@����������q����q{νZ���q��K�A�x����m�<��e�
هc=�,驛I����4]�v��D�yЗӑQum$��gM	��y,�kׁג�i�b�]�c���:�k�l=�X��(q-I�Ys�h�4ۊ��,�ʭoiUt(�{Ǜ�9H�W�k����xL��$l^��sOt_�?��?0݂�NÝ�q�nj�\T�K]��=Z�YXµF>@�y���ZfEЈ	��xc�h��'תL�Zm�g�{ל��M�V�,ԧ���W<�iLS�Zy�1��X�@������J�aȅ^~����+&^.�U���g����'\S�<\��|m�QʹR���*��>��/C���'�!@��+���|��ZCr�"�TYj8C?�~���^�
���`�B(�\�MaDs.cm�{mnmw ����gݬ�g�@k��0R�e�����$DBm6*e�mH��Kg��}G)�1��c<f 4��0���Q�
��6�wj�C�ȳG���?q�nu${FLs]=5[��F�e������n��	@��m��1�~���;<~�ыw��V��ͧ�.�"������<���=Ŗ�%��V3���]:N�)9Iюl�[�peDv>_)�?#�0d80	��g�8�|��������>xK�:hhmk�馡x��dkj�a�S��˘��hM��fo$g#��0�J��N���?4��f����~�\s��U��d�+V��WTS�랊��w��n+���-��@�{L�C�W`�?�!��
0�62X��Y<�+�ov�n�����O^G�m3E�$�]�ya��Y��l���W<������͇u�z��j�C�!s�b���i��൝-#����/L;�<��[C=�iO�U@�{��ʙ���5�fBzH��e���hp��FP�m.�	(���E������R�t�[���0̳;L�z3(k,�������z��利gC�:���$����Qaڍ�O@�oz�2��Y�%ӰApy�X�'�g��|X�-�7�@�<��	(���1g,����C��3˵��Z�=o��2؂9B�E����y����a��ń�!U� _��xqp�����v��ƻ�ew:G7s���R~�[4��z�*u���v�y�I�kb�T<_(\_"أY��<��X��U���?�[�:��^ ��d��~��P')��c��^�y0ڥ�'���Mn�ζ`ژ���'�ڎԱK�^�8�0� ��������Rʪ�9r7���g#'e�H�9+���R����`4N��`Q��ݨ5�0�m�G6������� ��O�}sϞo���ǿ^P�:9���q�ҩk��	��T/(Z�a�H��@Cx�zd3�l6e"���
g6dé�q�ϰ���q��`3W�)֠���1�w��4�P�9"��ݼ�zﺚ&��wmG���Ѭ hE��w��v���D���K?��!I����B���,�>��A��h����~nj�GC9ǆL�'�ӈi��}�����O�[�A��]�s�wF���(U�$���?i�+�~��Kߛ ka�c/��/%�{�ѵ�hX��'EP��g�5|<wvZ���1�ah��^K�^�]{���~ƭzpG��$�׎�`1�ū��ES[�?8UQ�;ֲ]	O�N��/���mB�Hؠj���Y�ȃ��N2��&`Z|�o�[ϰueh��|��>'5��O��Mi~ܡC��{��4�Iq�lK��;6�,�8��̚3w�[�Xk.e���;��]S��R.��ˏ0��X���'�1S�9�Y�X�eՎ{��X�樂kag�9?L"��`>�*�9kyߟ���޸3W�7���C.�gM�%�@�\),ܓ���eA�_>���e>�:^�T���fR����gtww���"���4sgmi7�U/V�z;�o�m��g$G�]�y����a�m�Q�e��S�O���Z��!�z�/�� J���V]f�,����� �_򟁃�8�ʘ�(Q��w�~?�+|��|��YA���}��6��:�ّ"2
z��qmt�r,ӷV��7ɜMK�D��w-sT>���dKej�wyͻ��|s� ?�`*;٨��/��3 B��%��?ϳUu���$O�#�<ǫ���˦ªD��SW�d�<�C�σ=������M���zг��֗V��iз𚚽�	�=��O׋��:�S ��HE�s2��/ݾ��h��4�+k�;����A1� C�q#��&h�8ū�"}�2��Q��F+f�z�B/߮�t��zB�=���1-�����oBʁ������d}f4V)�z1��q�e��m��j�M�+��鬞�� ��`�+���y,0�sVz.�U��w���0���p��6Wv�i�]�p���su�أ�$�X┩���zǐ�:Y�e���y�K�=��"�֖��y:BO��T�Xo#%��9�S`+�"�Z�뻰�i�(�ꘈ��w7��A"�^n+�6��G�w�b�1�/�q�>��c��Zc[0�3��`�V![�*�m��G�f�jua}tb�pqɓ�Q&��圉d�*q��\9�f�8&4��Y�����M�&'w|��r�b���w:=Y.��E��ś�>Fl�ƃY.�G���n�vu]7�h.(�j��S���⮬|<@#�QC���O����Hq���axM�f��Ϭq.� �N8��H"I$�y���I��'�-�T��U���|}=��`=Vd5�^�͠i�h/�MÐ�(Z���]��W �^ni|��4���̸�M��C�;���f����^�<�TsMiS��g�c\�b�X�}��zD;�fC3�ևz�`@��.�터����0ŬY�㦾~N��y�Zd���[���l�8�Z�����E���C��eb�O�=��&^���A���ш⣹f�e��n�W����L�Qv��: ���,QFc�AN��όÁ����WP3�o�J�nv�O3o�?.&����w�
�X����%�0�SN��r���v�^x�ʳ��س�r�A�rg�S[(���a.T�St��ՄBh&l=�(V+�&}q���G,�'��1{{�N��}bӱ�6ލ�ՅL��� P��z�ک����}��Um��Ob;!T\�+ʕ����a婆Q_z�	��M@-ܧ��Q*6`h�~w��1����"��T�Ǩ��8��k���O9�qs^9hkH��fD5�f�Zz�>M� i�k̍��������o��q����nރ�|\E⹓�F���L]�:���M�b��n�<�=��m���yBZ�P��T�Vn��m�.���&i`I�g;�:�,�XC��ЇĂf���2v�Gz���A��"��>��*b�'�(�-�K)�|�V���:�%�Q�˲��WʞѵcU=������7�y��oxxn���c��'_XX��I�Ц�g�ei�l� �y����IS��� ���1� ڷ՛�S'�l=֝�vk0ኂ����ְ�sm+_�¨�@��4x�V�WGI�x�Q=:�N�2sM,���iO7�_B(���v�:�dn=��3V�5��{���k��]Y�R�9����b!6�Կ��#�ih��1��	?7,��Ύ�cj������ӶZP�p�ܼ�43�-`([�#��At����#:i��k��քe�v�6:5e��]#}�8��zc��pAȃ�cc	�~
����g�~[�U��ll�F�iG9_r=����^V^�g��+v��^~ިZ�@pGZY��a"R�^�х��3y�ے��F�7o>$%��l#���zh34^�����F�;agf��;C��:hu��lK�/���������f����{�m��p[8�0�ˊn] ���s�n��������׵,��x3ݼ4w���*1��_�}%����T9:x�Q�a�J�� Fjz�L5;�mQ�]ӍVC5��UyV���T}��D������*V@l3W��,��kob��%U��3N���t�d��gP8>lb��<WL�f�}׻
���uX�}p��/��6C��F��� ����ǹNwt�q���D޺ǩ����4hx������6���YiU �
Ώ�j����:�G��ֳ���8��D�P�7���+�\8�Ɍ��k�w���\��6\5Sf�c[�3+m�T�w/�Ьc1t��H�9SЙ���F������*(��l�ŧ;h�X0��E���h3�����v<waU�/YԷ�el�.eA�����7X+��i��`����q��"u&��N6�2��n� ����
$�vpwL���@>��{6�,�]��jk뒎8�`׎�%�Q�$�ԅp��u�{%Ī�b�:u<�=maS5,��R�Ҋ���Jb�lu�t8��i ھV;)��0���[ב�۷AL�ۍ�8��<<�uw8>��t���j��]Y�A��8V�Û���6�!(tW����/�Yn.[��k�Ds�����͙��/���7k�/B�,m�TQ����)	7}<���^㎖���7X�^�o�:=N���e_d����v_G�yc�*6ཿ��a�!���a�[Τ�Υ�L���u��3�ҋ.�K4�^��f"��A�]��d�Uy�Nt�u��.zDf����9fPAe�%ګ6�3c*��O37�&J��f�*��4Z������knq����l�+!�V���(u�2��T���/G26jݗnlo��<���M�m�;.��SP�OR���`�����ZĲW4����aYP��曥Wv@wx�Α[ְc9x�vc���ٸ#쇤\��6����V�,��3 ���7�i'���{0u�����˹��+˔����-'�'2p������o&qט+�P[�CY]X��kr�&�V�ǲ�na�Zz���Ӻ�[��B�5A�7�8�nA�����Rv�[�7�A}�ga�ݪ;2u��7$���J.�k���i��w{E�8�Ĺ�M�t�����xm���r��^
':�{�S��"�K��f[m��즲]�Z:�`�S�Y�V	Tkwa�{X�:Z�]�S.��un�-�t[b�8��n��QN;�1CvWd��7�ecޮkr!�0�#j��x���WW@�Y�1v��_q���Zw�}d_[��U�"@��I�+���nn@�u�d� ����9b�t�*���m�&M����<��e�db�	&�.�]�Z�Eu��;	ŠjC	�[�Gz#/9�@�:��v���z8F�+���;�rp�.���*(���Íp�͝=-:q��������W�w�F)�5�1js���|���e��Ĉ���)�9U[�e3T�cT\�	�
���u��u���}?o��������AK^FEW#�"�2	�0������
����믧�Ǐ������}>_q��#�feT�5�FT�Q��c�����ܱ1�1(*"�̬�����*���������}?o����ώ=�&|��p���2��ȋ���%LFa�Am�]NM��Y9V`�u2(+,���&��,�r2)�
��&���"�1�2"*���$r72�1 ;L��\�0�Č�����*�J(�>�-�D�5[d1��fX�D�f{�o������0T�U�� �cjK3,����KTUTEF�VX�TA3���d4�fcE��0�������.k�LT�USSI��Q5T�SCT4Ifa���Q��m�D�Dl��H$�����C�o{�V��-Wm>���<�t�n�p[@������}n��_c׿���?����M�����:9�3f~�:��SL\|]�Bj}3�h�k��O�[0n�/�fO{��EC�n�0��ũlTV[��跈Ɨ{O����B.E5Í/�Yr)v2���S6�E՝�uu��S WM76��l�VP�ĭ3η���F��\�� 3q4��؛�T���[2g+!����=��I��Xƫ�J�_3�5����SG�q�kj�ǻ�e���:T;D��7]�كΠ��h���0�Q�:�\�M�����Z�a�Aq��{�ly��Mu��Y��#�����k|W	�/�3e%:����-)�#X�Klq�}����ܐ�̎������vW�/h4c��R� ��o�}]��W�F��\��x��҆�O�m�.��v)���k�K�����!1��WǿcV��esޡwF_�����޽W�5���z�"��Q��c��,h����z�C`j��L(ިa�½,C��NZ�+ɸzh·Nd2ݾ��3z1���4Vv}d�6���������@h��ۼ��y��I.��5T:�KiI�ݬ�LZ��W��9�'1����{�����D�6���/�B�-W�z�P���XB��5uB���ӭ�}���n'��X�����Bi�z��Y��m��5��Ƥ��	��5.��5w�q4��UFԙ];���3�/��*>��Ν��~z���x�
֭��6�dӆf�ׇ�>׍V��L]y佂�Z<��o�6�|��#,�	Y}&�ݐz� :�4.<N)��r�s�sl���Xi35�(9�/�O�Jys�>��y���6R(�D �O�r|�?�XE���S�/���9Q8]W��n�P��/\``m���晝Wekfj9O���{u�.�h<h�DB�ab7�8ܟC{ET;F�qqֲ�Xhs���]�Zg��~�KcY���=q��\�nQ��!�Ȑ�C4Ӊ�>f@5��Of0�=1[{��s6��u������k��m��t۸�0��G� b�S���	:�:���ә����F�k�_��^B�eVa6�WB�T�	mœ��\�u|l����.��t6F(�9O���%�����(ׂ�չ	�=��I��Ŵ6�U��0n˰˭���n *ǩ��ʌ]�	�9y�mǺ�Z��8Y�,�)�:��Ю�I��0HϱX�v��k�^ݙ�[�di��zkw������c=�ud�/���9����}����U�k�2�9sW�O)�!��"[C����^�{�j=��
�}ۙr^K~8����h]�����[�Y%�A+ =��"�s�&塁�NEku�}׋_mo:�������/��*p�2�|�{��9����3)�ѹgOļa��.�q|��D�h4R	&�j��i�Η i����v�n}^�W߶�X����MQ�./�ڙ�~帾,_��z����T�j�����)��"�y����m�j�m��c��*KCP��կN�"�㼌������ϋ���&�g.�O��"����M��Q�ʟ1�a>[��vׇql�F7T�Z�,�ɚ�v8B"19��u�"l^����cS���,��	kT�T�Xm�b&`7��G3�/Ç�+�%�|�G�*����O7�؊���Ž'��֕	�5�����S�>���D�X_}�Z��i�L(��';���=Թ':a��B�92t����m4���%�P����j?|Ƈo��l��.�cm�a���`תә��f!�O<
�C�c7)���r����ώ]��#"/�)T�9;������D�VY(��5V�#���C32�p��q�O��Z���D��A���_ʽѭQ&rx��6�}���Ȍ|���.�<zBp�"�T
��ŕ�r�h�a�;�`j�w>Ϯ��Q����$���o�U�5|���\_&B;���V��{�h�9 ~�^D�Ko�+�g9��7���p�U,~�ܣ�����q���&��^V����^7�����^2_�7r�� �w�� �;uѰYX�
�����]K�v�<ݽ�r��=�� y"O�rb����76���KT�M5M�#^Y^�+s|E��.Bm��(V=�Ƒo.��u�A�&-m�څ�zw֐���Ơ��oR�Z�t3�s@�*��T1z/�O[B襐�o���L٧�M�&��-�ۉz�׶0���%��K�(	�T&�a��G�'+����}�*��t�l�\٨TĽ�3m�N0��� P��W��u耙k�plM�Mf�^�Y�Ǹ���(�zs]0�UJn�J=V�~���n�c!ܸ֋�E��fe�w%�T%��r��R��4<5F��4W�̮q^�x�u����ҡ[�J��\Mf��f��!�5P���C�k����z"���ny��>�<ޑ|�%O'!B��~�27��cO9�M���!�}�4˺�L!������J�X����g�(�%݊/����I���ݭ8��B��!W�6x�`T(���Λ��a�m��?[��P�y��=;G��Ѧ<�%^�mMp0������*)�����Kȷ����y;z��Wn2��wf�lha�e�¶����׺���D�-�Z8���Җ~/�3��X�g�I�Ѣvm^��/kJ�P��*#��5���}��b��v]�m�%K�=.�����e�q�.����7�j7z�A#�cO;}�R\�ǻD�Cȏ7��<��z�	v�����·m9�[W�XYUy�ꅭ�GqN@?�@!�[�|}:"j%_���t��:�ɕ����#Z�"��zFљ�1j"�dMm�W%�o�.�J�f�_oVm}	�/;<�c)p�F36˝ֈf|����|�g�`�����9.��1�d�zٯ�.�z-��fv)������Dŷ�sn�K�9Bh.�Jl��k��Ϯ�?$A3$O��<_o6�~���>@���9O�j=T�ì�G�����j�|m����}���Z�jt�N=�.�I�x��@^����8��,<9B�����r��X�7K�J�u�JHnk �2k�������U	�زa�Y�3�8e�%�#DeР�D/t�ߟz��s:��u){�G������/m|+���V�'��)�@��s���vH��t�z�A��/G�Pʌ�N�����33����Y�o	�L��0��	��м�j���rr�C��FI���4�Ø�g�p<F��W��)���,_@N}�ӁlF/��>�C�� �`��sr��]=��Y��,<��+}z+���G�7G��[F:��F8�k�2�y�v��̳j��l�3^�;sF]q����hu�-RQu�N��n ��kr��g����E\ʺLΠr�(��De�4Uqb:���.]`%@�K�i��?�y�7�0���N�5�G�VPv?<y����O�بE��K��WtF_}tk��Uqo9�~�on�)�t�j�!B��a'(l8�x��n�GP���R��+8?�쭳�z�#F�zv9�ħd<�����̋�d�'ω)Mkϖ3�g=�����!F�З���t��UU���};FQ��0%ݮa�����/{:�y�� �k�[vng�x�=эs�'U�އ��ί_	q��{���U
�)��;C��C�x�kO�r��0����k��Z7�R�BX���Cֶ�����yA���_R�ZFsp�;�9�h���N>[��������JW�#a�O�B��[&�OU�^����˶E���U'��9�Y=�6��^�aԨ��=��'��6�c~bIRȎbۓ�����3�LF�{��̣�r�k¬���������3P+(4��]s��GE�+��|3!�6
z��ql`���rTf�C�Ets(za ��=�m�ъw/�^�5��/xJ1��Br������M�_%�ݙ�.5ע۵f﫡��!?_��Ta`� �M甎O�%�D)�����[n��q�~�w�0�O����AJ����9�rh���w�W�yn��c6W�ہ�ׅ���Nך�_V�����xN�U��r��c����@�D�}��Ih!�Yi~�gP�mg�4C��#!�ZE��!����a08$��������i�{m��!��Y��^*�Vj�a-j�!�uC��`$bi�eV/�^��6��1��"��	<㎍xMM�鎿�O׋hiQv���jv,D�PsK��N�9݉Z��ml��&,��u�����S�Q��@�a��M�J��oE�o6ۣw �{&q�>��ip iS�P�VH!�Y��{��m�M�ڻ#U���͗K��J)����d��MNdE�36�����I/>ƍr��`?~Vh�K�~�� �{�x-���x������ b�6�Sͨ(V�aF�3��=�q�Λo�M�1ݵv���n�[h;_:��@�f8��@�\��2gΊ��6�nJ�вt���UP��g%�p�w���7�H�����lZ4*��x�9�	���q�
��ZcZދZs1�R��`^V�8O��ϭT�%Q��'L�����2b�{�=o�Z^�K�`l�̌>!��4s�]�ig��d8�L/�(y��L��~1�������i�\�`��w�N�b�ȹ�۽����u�4��K;�B����bw��g;x�n���1E� _g,���wJgO�؟�e{_Z�oq���������(e�i.8�h�h���+�l{���D�}:r��;�u�ȯ;)X��[}��#�x��<���|ŋd�U
�=�8�h�j�(=~�	��y���A���?,#,=�5[�4�'YuL�+'3�L�E�ǰY�(O�~�8��p��m�-Ojec�#����S��>�#3WN�DJ����E��d��ݨfG'��r٢�p�H*m�q�hO���c���z�Ϟ_�Y~9�O[����]
j.VN0��A�q�y�1��2}�m�<�WP�_�s�-q�s��t˺��ӷxb����ӐK�,��&��'g�+��D	���;e�_{ױj���Q�}_��s�Jͥf��΍��A���.{�?�+s�#ڒ���ױ��,#v8EGű�,�ou#yb�n��ͻ6��{�f���s�tv�AT�)�l�4�T�c��,�p�Tζ�j���٩ec
J3"z�\3
�R-��2�i]�����źYm������s�t¼�Jn�	U���k��5��d3�Q����"���F�s��B`:��3Pv��t���%�Η��3i��s_�c�_��w�� ��������!�m1�����St�x��7�W��i�k;���ف���ߖwOpֽ��^LǑ0�'2F�KM����Q�J��v:5w�]��rC���9�1e��p���g5@��%k~�M!%��j�y�q�3V�|��1�
��K���qkg|�鉈O�Bz^E�1�@�1�or0#IU���s.����pl	�M�Y�Q�a��.]���5�ε��K�0wt���L�׮U
fY���s�;�m��]�n�ርG��_d(��Ʃ�K��Hf}��$�����>��)�����}K�M4�8�&j��B�gB-���W����k�=9�� �Añ�������Qq�ʾ.�'J�X��ן�����BD�P@���z1w�߮������q�f�z8Դ9j�!��*%�P�`��m�Fk��u�j[Q	�|m�/#]��ckXe���3E�a���C��q���Ӓj9s�kM����T���Z�fl��^�7#ps�-�	i$U��Z�6A�J�.6�U���r�[˸�DB��Cc��Z��[��-��-��B�9B�wo.˶�s.���i�c"��Sv��T"w蘚���Fy�Ҫ���;�0�J}[������ԅ���Mo(��mt^�T�F-�$sӸ^�YZ~V���5���������Xt��ƛ+�
c������R��v���P���}q��w�]�TٹN���O:��V찛Y��s{G�}��&���ú\R�kh�uk���Nui����y�)̾g8�����,(��Y��@�EZ�r�隹�����_����a�� �Q~9�w"VJ^��̍��D�l����۱d��jn�20�MX��3����C�Fd��jՄҜq��&�+vA�xX��wBeδ�'�qd��r��熨�~t�����qa�Z�oN �Q���{�����ӿ�OZ�k�/�a���*��e2Y�+&�[hJT��SU��Y*C�3��!��f���(d�"㙢�C4bS��}qʣ��}��r�y��"u��cGD�B�x��`ue;	�|;Ѭ$�!̺ZE�74�t�H�S��W�����U�]��9p��2�=�ň��P�5�=�-���H�g\�.�42D�O�Ɋ�&3of��f��B��<_%�&�WO1Xa�б��+����XW��~�BkyU�2���)g�}��P��|�T�Ω�G�zECL��h�,��Ɏm��{pf�܈�b"t���Q�Z�h����z�,	p��gZ��\�@�[0S��~'��Y�!���ZxŴ��Cd�s��+�#C�5�hB�P�\$N���1}�F>�6���}�>�o��N�e�q��t{p�Pvң���k6�ݗx��n�pJH,���0�E�O���)��Q
��T���l�jvXO�M�f�v(�fk�����<>�2�ѱN�᭽�Z�k��F��ui3��x��Z�WX��v*�N���	�-�.Е�a>[}�Y��]�H.�;I��\�c��m�1F�Lq���CEc�v[s��Nx�t#	��}|o�n�F�4BC7�y��4��N�����h���;�@ۉ�$_n�:�Y����Y݄qvN2'F�2���
L�:�����m�� V����v�|#��6]�`�҄��h������L��&	������.��֮]ەuu���|��~ޕ֨��ayp���okA��Q�R�Wm��1��%�e�v�ɜ��^m������eU�v�Mv.-�VJE��vh������I�)�e�<�#�Gr��&�@��i��a-G�1SkCn��BZ�`��+��a����ڬx��)N��ή��@�o=��w�����cn�TWͧ �Vp�1�R��q=�Z�ьK�Lлl�a�����13�Cq5ս}+��掔1iun��vb�Z�˽~{��`ᆷ٠ҩi��.G�Q�]�yy�v���X�`�\kA����<,�;�>�Hi�i��k5b�Fraaŗ6�+��]L'��5}��A.���j:��_�M%���%�7+�VD��!�d/"M��&���]	_��?�St�\�^�2c��ڵ��I��]�V���}���.j×�hA��_3׸d�R��5䆛�&,���H�Wj}e��R�❻�ۈ�0e�e�a��|��`87�~ԟu�c�;�Wj0�IK���%A�#f,]�zoA��S�\��^:�Z�|��e=�x�s놯�M{����N��A���v�L3AQޜ�lu�Rt�U��2,Ĕ\�##���V��e�1�n��`�-�vr�wT�Nh�&l�ټe���Q�vñӞ����d��J��.�J�Y��$+�i���۝�4�\Ĥ2��:�)�\�s��Z��������C/�}�r�MZ�ߦ�V�qS�T�"������A�H�T�^X*���͵}*w.�{9[]���a@�T\p�*oXчsw`}�;.�rV���x���`��x��N�E��S-�Y���p�B7�54ѵ�ȸ[�|fvf�yc�UwD�7���̷sz+��X��O��~#	� ̞"n�9k�F�͈sqGk��K7���
�kA�v�+2���Yy^���K�L}�v�t]�Ǚ���D�e�6��컣�p���@��P[�f��d�[rms\�Ԧ��g��]�1�wf��,Ӷ�:58ΑV���1ʠ�bM%U5MQ-MI1�e��4�G���OǏ������}>�����W��U�{a�*���er�*�������0��a1x�q׏�Ǐ<}���_�Ǐ��(���c *���(����ʢ,�i�!�JB�j!����u׏��<x�}?��|q���"�0)}�r)���RPd&U�c-)A�`PQLNFE�[�#��MTU\�� ���eM�Fn!����R�R�9XfYD�dcPU[�UEndP�Nf%m�SO3�>f%-�&&�#�%�n$UL�{��-̨&b���)���r((�������!�\� 6���J�AFI�Ud�de��UT�Y��dfaEP4�D�1D4���*h�d�'!2J=\�M!B�	f�Os)j��b��d�T��r����Ͱ�*'�$�>D��ЍYe0
e�DA�03"j&��FT��L�A*E
D�bT�'������]{�ڻ�t׍�)Ý�������xCr��ƻ��|\W�wN�\����g]5���� 5)�PH���$���>22�D%8�%��P�L����bM T��R�p��i��*5a��l��JF�P�q�ߣi� %��0�? ��"�
.(ג��a��~�����:�i�d)�!�?B�m�!���!�q���;�Oꉃ�����|�P�锋�kn�j}{���{3g��0�r��2�wcO\G	Q���K;�ꟍ{�v_ʇ(��P�s���q���O�ug3��\n�����3az�oAf�6ь�
�>�73
G�TO��_h/mn<��S���p�����S��^^�O�-�\7P�ק`'_�ϹBI�y�����#6�$t�㚈�&�);ˡ�&��cy9��1Df\
�4��Ql%:��rK�M�ʤNP�X�����'I,5d2��5��|��2��y�X��p�����%��8��ѹp82hj��ǜ�)��Ŵ6#k���׷����괢�Q܈������>~�ٍw�A��L���r:G:��9�0��l���WK#bLs������E��6h��/B��˭B�����΁)�l��k�V��0�H�
o��\#��̎��7^�E2�8�.ag�׆��S1��!t�Va�����M�v��i�+\�Zn���b�{�;!��!�ok�P��^�T�{S�9���(�/'�]�C�����N7�)���h�ge�u�ު@��V�Y+3#��m7ӊ�Y����>
�7�֩q��vhS��v��K���y�����u�'��a:�K&����"�I.au��,�
0��f�r#��I���2_m������B��R�先�>���;����;�1��u�Z2$Y�.(�U�,�%���k�W��kI|w��Ζ5L��������㸆� �9�0���8��)��=����\ل�
��eIaې̬&Y-]���ZM2.�I��;0f���y��xheB.y�8���b	���X[^⃶���aU2U.��A�{�>v �[Bz�6�	�,.��!��{mW��_��M��L�B��3U���6�mG-�H͒d��[���vQ��U�g!�Ge盖_vk�j�b�i������$Q�,��v�t6\�d21�6���Yu]�M������q�ݞ��x�*�|��.�}������i���}���&Hk�"9��Uq�(5g���o$:���1S4�w{N�����1���ܗ��Sz&|#����$�e�GqX�_��N��9i���d͠U��w�������H{����_G��TU{,��vi~X�KWS��γ�C���,"�ʝ��X��ݢ��z�uF���N�石��Q�]�c#XW�L>���w^��_t;���q!֒�l����ܭٯ��Y6{+/�R��R�҈�ص����o���!�<�=�[T�I�uyz$��i���
Y�z����j��v晙��Rt��8���ݷ�8��z1P0VRR�,��j�%��/T�a�jr�*�ʱd��M�Ix�ڵ��+�@���\%�<���w"�:�6z��sڒ���n���`·���d����4��6��畊����J��k����Z�e�q�[@�+$5����� �V��^@%r��@��#��r��:��#Xh����܃,#��J1S>��T��a뵛��/^�de)��$�]��]�,:V�u�M��-�-�RdDjQ��9���F{�5/�^Y��T涢c�{�|�Ӱ�p�}^�6��Ŭ2K=3S�3GQѨEn��Z��ڷZ�p�ۮ��NG��?O����ݖ;�5�������ܣ�����3�t�se��@1=<���o����+�Y#R�X+u?�Ac�'OlS���Ee�«��,_�s+���X^n걷t�m�w5�����o�$�^:�}�؟}����ϻ�^���b�� /�z�ڍ���N�����K �RѲq����t���֖;�f�GWU����oy��l2hŵ�����l�� �R�>-�m��Eg�d7��EFR�1:}N��g=��y��1����b��^�	��}3|�3�U�{x����/��l��Y�Z�`KH`��XǖZ�%c��L�
��#_�F�u������=��[�6:;*���Hvǚ�ω��T��(�<{���i�ʦ���!�2E+�OVWM�ݗVARnVW���%s"���f��Q��������m�i���6���1�f{���9��jRn%^���U�[- �p[&�g_{���BC�\�0pB����[�,��u�`Il}�w��x���\M۠�v'1�MpB�´ZW�6w#��۱�}�����v��w�org�~ܚ�B[0F�
+���-M��[�]7^p��m#�d���>(�z�:Iv�l2���<[�p�e�`Pl��oG�y&��^Q��K4�`�z��r��H;�5x����j��(̗]�A�\R��T��@��ބ�����PƋ�%�{�Ў��Թh9������B�>e����!S8��ٴ7j]���w}{�����̝ͬ�� wNZ,�B6��ض�v�WP6BGT2�@BQ�FA+�&`!�h��E��������]%@���9P�xc��쮽���Xˠ��2������vb0�N��g�uW��]I��ͻ�l��u5j�v�Ibi�m��wηձ���mv9+������*��ݧ5��1B�C��+�n���.e��=�|��
4*��#8�i��-���ӪM��/T�l�l����^�d�+AMg4�W���<}"QYML��w���u[�4���wWW��^N�1�~�8�H�W
�T��Yw��f=|��^q���bS���w�V�l�kJ�z
�`�N����x�g�	��~}�\;a�fٶ�xb+�����͖�6S�B���r�[22��E�*m�4zv�&*���]�:�5$SA���L���#���d��SE\{�OP�j�Gf����-�q��r.a߶[!�����NJ��1��YG���=�;ρ��S��������)O��A3���^+y��6	W����u��ټb��:��WEf���f��'�q�KH��!�I�>7���7y�!ٜ��ᰁ����εE}�G�:�.�t{pl�omrn�G,@�*�毋"s��3�f^w+��ȮC�P �Fd���C��Vf1���5��~��ȇ�<�������lw}�'uv��v�۲.F�rffw;*�U�U�ȫ޲�ֽ���סf5De�
���-[����Y�����f��uHT��w�4��Sq�Ҝ�S�9�����7E�ՔdV�_���H&����R�]�z���ۓ���,�Έ��7ϳOW����'���%��pT�E�3��Z����;�i[z���4E�h�`1�mɏK��!������v��z���)wmP��ݯ���+����.J!�S��j@��g��ϴwG�=�<ښ�w��a2�=a5�[n���b0N)���Β��o����"I�Ү{��}Ϟr�R�6٫�Փ��6wv4;���^z7ev1�I%H�_ f��4�l:�]��L=�Z�s�[mmճF�+	{UcX=��Hףݶ3���a��hh,��G���C�|=��=ߟ]1�C
���\J�H�m�Zߒ���y���^�l�����M�⩊I��M�.����X�1l�W�5�����f��*�;8Q���b�'F�	�DZ��N'.��B뢶��D7�[�E��d8�o}� Vޓ���|V숳�m�l��~;|�gĵ�*�O�u�j�W܃��iy�f�t���C?�L,zQ3����S=f���|��	5�����nr�L���]�̹S܋�g3��«��L�jN&�'�Q����'e��gvl��'oJܪ��˽����pܩ�%q��)�<D}Yk%���W�e�a�A����q�� U䭶y4K�ʭ�YS�7��%w��\wޤ�A�J[`+�,��Z�3%����P��/����`6�=�3z���/�Qk�ռ������c��=�_��u	 ����Ý*�5W�é �����z���N����b����f�K�b��;@2�h	V�Z�Z�7Ej�*���y<��Alÿv�&���c�ݑ�C���{@�w݀��>��-�}�J1�����u�����o>t����*^�͂�|�=\�΋�v���c()c,s�k��w���W�]&!.�w���y�E�WLun:�:"����g<̵
x,��۹}x�a�R(��,�Cx��d�ג��0[�`��5[1��}� t^�Vq6Ѽ1�W��J%neW盬L��n��uǽ^��]���4�j���~�3$93�����9�\����{�Wz��#��{�Tq��H���yU�q5h��^
��I��=Z�?�j���=���v��C����C�_�3�WFW�Xg�
S��v�e6����tɉ��6��1�h1��	8�R��0ٲ��y�G_LZ*�a�v���~:��dM����ļ����SH\j�Km��ؙ�_>Dġe��]�%�b��ν��Z7�����:h��
�hi�Y猆�R"�|�������qf�R�Ú7$�9P��D�C'�^)e��<t���Ter.��ǐf�3��-5�=]��}�۟���wN�
��gɠUͪw>��A�TyS�3�j'Z:�C�{�����:��m�v�eVQY��Zo�~���V�/C�ti��̧6��â�aєl��^���J��y��D�)&ŶN�2��ɏZ�%ʴX�Y��~�	���;_�Q�޺��q��y�K�R��"Q`��| ���U�t����/���7����+�v�v6V��7h�P����I����?�(�������ŝoq�f8�^���-�Ӓ	��D��?����?P��<�}�M��.�	e�s�0������v��`s(�8�d��"���\��/ �Y��U�K��mf,X����wC宾@'���c��ެOC����R��� \#��)�)C��87�o'X�������I�(��μ>M�e�0�C�{���;'�[�����v􎒹n���,j����h�ߘYU02f���7�e�oH��w���#��v��$��wAƬ׾	r{9�QUGZc��l�a��O���0f\����R#Ln�g�WY�vr�7*d�rd�6�}�k��?,���q��
z�\��Z4ܱ���O;��ÛpM;;��4y���ӈ��ؓ��?pÃ�0$�}0��	��֛�hq��\lq���Kخ���vv�~T�/_�:hl3�1
�d�{r-�2�����^gw��*��z�|����1��I�}\�+��y����K,��]3A�ǎ���WӠ�i]m�G�۵e�w�5�����K���[�|WQ�h+l����W�����804�h��ᑙYL2gO�WՉs�\'O%o4�W�b���Q$��P���N��!�_E[���tк��Q��F^�Vf^g^�M�����r��V��Qf�8�����<�m薮!Ҁ9��o�#���I^gEd��`Ua&_l���[�SY�.OV[*Zm�!���G�?MO�Pv2��(�U���ڊ���ȍ���h�A&��`�i�lX�}V�քC��bQ[Qxs:�n���sS8�$�eߴ��$�� lJ��wVƅ��Y.���j�a�ɽ�=�����ݷ�C��p��^�jz�@�l���2�l�xW߰��Վ��j���z��K��M��yQ\��	Vs�E���'x�Z��5�ױnr4�9]FAwS�vʋ��o6�9��{�#���Z����sB�|:m�kY���f[�s;�g����oP����3�Y�4s]/z�y�����6U���q7h�Dk�]�(��6Pa��e\��Zmi/Os�ݜ+�GVk��\Vi�o�LW ؝� ����ްZ�ZOs4���b�T�Uȵav�Ԯ�A�t�k/2E̒�q�l֞/#�ԥ�,�0�geJ�OiV��Ow|�u�2�h�9����,�1m1�r��N=s�K߯������=�UO�xݣ�K�r�m�/8d�}�쀜Ҵ���Ӎ������.G�_R�F����{�%d�_U��瞮�]r��3�����P]�y�/th|�E�]��Gg��2���͑Ǜ&�������E���M ��:��o�p��(�F�'ݒ+���s�F�^-�o��qcP���ѵ�
�����x�Z�S�b�Wh��:�z�^U�&u[)�pp����������	�ʗ�t�c�Ve;���[ѫG7L���R) ����[�w�����e�/7hhMd7����Z�>r��Xl��#&
!�nW�$����ّ� �y����m�+��#u-�lʱf_�#m�W��k2���C�,��`�Z�Z���ܜ�S��l+�e�m���e�AL��S��B\��B� U�2����7ԟz��i��

7/)qW�HY,&o
����RAG�m픩�i��@����&��E-�ѓ��ne3ڔ;�I�{���V��ʹ���!�(hJ�cz�]3����{//�K�RԵ��x����	Y�!yr��@�����aa�\�}�j�
!�4���N^r�Ŵ�c�k�ee9"<0N2����ѧ:�JK)�k�2�8Φ�	˻8ያ:��Ѷ�R������k�U�OY�FW�%�x2�h��\��f�j�v����W��E�^���ү�BUR��L@��X��Qك�r�N�Cx��9@)��f�����W�iG}7kNS�Oq_w���(R�ED�!�S4P�'�QKu�n�]�E��˘�^�;6^��>�R�6�J+�*G.��2V�r>��pk\*%����3����,�����qQ�Ax0��ᠹ�p�����.yp2� ��7x3�y\�[�Ea���3��t��s�ַ,�����S��`쥢�m������Ed�h'H+�9��e��_��U�����wX}4i2�[v�Z��Z�I�2oWWQ����Ytk�1ڪ��>dOA���D{6�lRK��##
����U��R�vbu�'%zl�* RPY���/�4�38ݤPV��F����lz�iu����&�0�4�������N�=�P'Ws���	-����n�;]�g1���T���&�[mKVRo��G���9�\pX��[�C4��k(�I��V��;���<�h��7�&db�J�Vɶ뇤�|6a�Z(��s���Ե���))c��abV�%�Sδ�f����u��3��{�oÄHW=�l�fAQ�	�e�2��U>�`�*�z����X@Q1�}������Ǐ>޽�3�|B���h���0r����*���r�̐����(4��9jm^FEA���_o��Ǐ<}�>��Ϗ��AS�e��eESe����R�S5�0��TH\�2L����^>><x������z����yw+cuň+�)���2k,�"�jB���|�f4SU�%�������SACAEL^�>f�3,"�� �3(hy�hQ���߼B�9)��@U��
��(�!�f>Y�I�8M-�TKA50TQT�M՘����Hb�n�A7#"!��j�XT�P�SQD�SCIC�1�
��f`P���a�O3-�mMR�Q��b1FI��0-��2����(�������ت2*�9%;T�\��Lɗ!�nYM5�5M�7G"
2J�n�dnn�>�2ߟS�Gojuu�]�'�\�[Ξ��I�\L"��ӫ0p�;׽6�Ћ�������ו�t�͈����9]V�o�$`�Lkx����p�����b5;����bCa�Eudn�Gz�#��x�܊�=�~�W���>��qhlJ`m����7.�#7b�z�sp��w�3a��Y��h�x���î5��΋���R�XeL�T�L�A,�����-�st4�og2p����e�"�AM�?1���w>���C��uG}�.t38�s�5��I���a��*<�ޖ�~>��s$<i�>��K��6n�߹�ڀ�&$r@�!�F�j���3���ls�3O�)��b���R���wT�R�!#<�oY���6m��މ~�[���l�+l�ȉ��w��R�q.7:�ٯ��c(5�{{2r��Wf�4aer���+6�m�=Ah�]ߚ+����rmΫ�u�ea7�_�VgU�Ra%IJ�99>�o�)̊|�AY���g6EN|�fh{�)J�2Ɵ���0U�]nʕt�&����8fo�]��}k��X�i�R����t$(,��}徛�<�yqDIg/�ۙz7x,
�]U�#	ޮ��i]���,I�<�챢'��A
���ɥ���.e��˖�"�2�*�vgZ׼�WdoS�.�vZB`:��'h3�TU*���W�J�ޮ�u�E=g�ܛ٧>�u!�1PdV���6�]�����U���բ��M��Uy��f���0dq��Ԛs�ڍX�6�9�Y���E�v%��z5�Ԣt�|������u{mE���8|��ȇޟD-ꜟ��-~���~��t^�qr��]���@8�]ʯΜ+i��6G�?��8�e�X=�M`���)2���o��e�����
��#N����y�����
q=̶&��ьپ�v�����X�8�w���ǝ��ݗwp�T8 �IӐ��2��>��Y��vĆ��+7g�R.����^�fSQ*�������q=�!��l2ὀ���p�`�Ȯ3��K*>y�������?	�q>����`�� �-v��|�	@x�T,�g'R�/��G��;ۯ�{��CR�rZʙφR<�Le�q�K$�ԟ>��״�'ݰm�K���S�cmq���`�G��=��d����_���Dk���f��u,�dcW�EМ�J�WӋǔ/��=��
�S<���t̖0�ة�]|}��ɗ�)������߅aֿF�2
6�n�~�k�XRiT��b&������D����pޟYT��i�X��S�P�;�ty��R���̭
���� �r�!��2}��ߩ,g�kR�rSL��]�y�jl��WRv�RU"�4rVP+'	W:2������B1�y���{?*����ʐ�/�^���>΅���7$׬��xD$�wp�yk��z�'P�V���M[b�8�}>�I�;u��K�vo7b�����a7�d�Y�[ ��wj|��­�[���ëp������/��l�+uX/+v�K%7�� ��;��68���No3a/�04&��
3f{��0FO4Vn�o�?2Z�)�rAG%��&��6�g��'75�,[gbi~'���,�ٙ޵y	�ӑ��;2.�z�.R�V��HM��vd�@���zw�t�g�S�]Q��1k��uGv����WBܽ�"��,��&P�j1�A������:K�|�.��M�,��)�w� ݼ�J����qg^���h>xX8&<�82�s�ݨ"]����Nsڽ|&!3q{�W,����pc��*��I�cjm�r��C)e*���u�>���u{�v"�KIC�K���v�f;Q�d��C0��wq����91�9�n6u�V�� M�>����_�+����ű�L�����Bc3n2ox۝�ϧO�զ$�{�,3�x�0�	<�2�| 'H��:��ɫ�l'1���z��jP8��r�#�\*�mM�Yx����b2��0ٺ;y���aC%��F_�ڒFw6z�pHX[�K:��(�ܸx�h �fsǦ&�W���/|�d�z�- �Q=�lasy�[�K�b�R��S��r`�4�L7K�gbRYC[ Q������~9[x���[��w��k���vi曏o���Ȩ��k)���V���^����QYk�RS�V�� ��M����.[�p�D3:穞y�'�nۭ�|�k>n��q��6�61VM+�UQ`~��z�w�g��MS9�@�u�,t���>[gjQZ���*5tGWO��l{����hr��}݉�۾Ph��G�K�,qǷ�-�#�62������ApŰ���wH�9�9�;�X�_v��vR�J�H؛�2+%jy��f�	yȹ���Vr���M����"������|>d���Clg���?wXH�#{�����ܑYR:g���Vv���՜���<l��������({;��
�\�t<��px-[c�t���.�
#�d{���(��t���˒�١���j;�#:]�֐�JA6�f{�-���~�;�hOf�1��M���k�P�ӹ��.�ώG������V�1�:Fn��ɛM������D��ݙ�W������C��];�q��>ޏ>�,|ڢ�ꍗf~m�������+8�z�>�0.�����Él��ۥ����UU2�3�5h�>���5����Ź��v�Z{7,p�FAzv�;)n'��f��<e�[a�����#���d^c��w��%��a7���׫"r�:�ﴙ6��P����]��=�Rީ2�/K���.{�8��y�mnb鞺.�ഴXΌw-������Lm!��>��g0�p�j�/�t
��~�&~�	nd�h�zNďv����w]ՂL����y�ӿ�QW��,�:��=Ge٘�۠Yϻu�\ِ!�ƪj��lf��W�x�}��� ���f6\��K᧌
��=5$�oV#�8��vf��yY�)�W2&�֮�<�x�KU�(Fd7*��5��dvH�q��o��0饨��Ah�8��^R�gƚi���(Vͩy�؟8�z��m�:�Ji:�ݱ'����I=y.�%�V�,ǝ<e�ױ�A�wXC0�4�^��r��+->m�J�U.�	V��W�e�%Q���N��䇿V��߲��=�a�o��R��z��5�kCsԵ��v5����-��u)-���˭�6�Е�1��i���KA�����q��B��'խ�X�Σ�ۡav�wY�`cMlխ����ｴ����@��������E��[MΦ͟>��-�os�c�_ݬ��LM۽������ڷRqj�;�Mw�ϩ�
9�٩���kka�,�,Z� �O���=�>�=RO���l���Oj~�O�v�0�gn�)����`*�ct��n>_&�ǔh�Z��k:�'I�|���VT������4�7{�y[�{i�[{�_� m�D��q���V~�88���p�I@L$�<�A$��R	~��S!م��?��\��.K�,�;�����=9�&��F���|�u�^��ud�7�������Vj�է�ӛ�D&���bb�q�~1}Z�Dk�u{����wU��"���X��u���z�xbʼ��]n�-��6�)��Y����|Uw�ә�Z��\2O�'l�k�i����S�(gs.�l�R���!���5Z�H�̜ny5��{ԯUW����C�1H^q>��j��F����(m<FTC�MS�Vޫ�Ǧ_%]J1���=\U`��Ǝ7�es�TMnΩ40dWD�q�q���12��O3� �W���twC羂�WM
Jr��}�t���fo;�o�jU�Zm򭖃Zj�9Y�5�6�$.a��xa1�x�S��{w0�=�G+&�-��c����1�`����k!m}��,T��7qqUXۚ����rHXɒP9�	֘�p;�ᬆH�nl��U�Ee�脲:�b�ث1��þ!�f��� 'ޡR�ё% |��\7�^p;q;<KC3P�뽅�eNMԽ[	�ѾL�����Їnnv;8jI7�=�nWu������n�������ݴr'j�l�ys�����[\�Q$�1a13�`3E�M�G\
J�@��ff-7����@@#�� �m��>M����Y���ߣջm�z�lQR}VxώR���K-�&��ri[Hշ��s8J#�kw����(P]�&y�a�ū;5Ԝʬ|lm�2��WGqiq�8���ŏ��g���d�G!c�®�"�C�˗S���gj^�"��3�Ɵ��� � 3���8U�+�Y3���u��_714v�_k�fC�b��c��z.^��,,$�u���u�I�ua��E1�}bxX�B�������zd9�S-��m��<-�W��;c��r�D����vת�IIkU2�o{:1�Ё"K="YOi���]uq�ٴ�q�1~���S��4�q*.���{��4J��4،��f�ېK~���Ї���I��J8�2.G���ۼ�����L���y�f��a��� +\:e�t�
�;�5va��Uzd�z����U��7/䎞�״,�;�&�������y�]���h�k���=����2�ٓl>��L1�D5��V�}�f#`���&��j��3ǇKly��.���EE�
n�pCe�n˱�p�ʝ��wtz��]�쭰��u�[��׍�-`^�ߟ��q�Y����pљ7>q�nU��듾��*��TM+�T�ulfZ����:�am>=O�S�sk����@�%�Q�ʿd���)��c����ݞKbQ��w�}&o��_t��Y�u"���v�\<.Y��p�E��Z�<�)�{ls��Ź3���9��7��m��;;	B/g%���Ljެ��t�,Z�Y�80eUH��zǍ��H�^�:�����baܣS��s����S	�cS����"�3_��ڽ!-���akN����Cv��Dף�P��d���i��T���n��KԊ2��ݑ�n>c~n���n�b���ba�yZ$4�U���h\��k�Ė=�Λ9���[d�S!��8s5e)�@ԓU1%�<��Զ��A X��}M��' �[�7�)��fn�Pq]�v­���ꆖ�v%ϩ�3E��(��-�-�����P_�3����s��,�ø܁ǛQ��4����g.�l�j&��A��෫vœ;�v���]#�s�@�W��%]ɷ-�Lպq�N�l��v`�B��m���|@���ؾ�j�ӵ�r��jB����ӕ����ŵơ;��s=�|�A��a'E^�^uS?��(������8��]knW-KU�w}+�;-��+��b�?t��x���+��#p۹�:�!�!�!x�|umrY[�X-S�l�{�nU�.�6Uǥ�)�׏�Գ�ʫ0]V�r̭2�|R�v7�bm�c���w*':y�x�ه|��@����u��t���*����k�v�,��M�����*צ���U:��5/�mg������*]Ъ ʖ]4t��3&��q�#z��̆�T�@�P/�y�r���g���k;3��92�ֻ�؃4�sv�)��Q��I�U�X{Q}Xl,�S�}4�L�X)͡�."v��N�9���1���8�z1��r������L{y�Z�u�����W�^M�ϩ��J9w�+gCϗ���ǚ/��1TB�fӶB�n��-Q���9XL�����.�:}�N��
Cwn��<����n���e���̖�Y�����F�w�̳r��(��&�vj�ܕ��%����Wv��f�e��bհ�˦�v�$�G�u���6v�˰0��]j�*)��y�乹R-s��9����g�*q�&�Daއ��]�S5nR-�3{J�eټ�,#a�ж+��r�]�9�Y��,2T�_J6�eNײ��M%���1T%,e9cjk��d�mљ4F2�^�+U聲o�ʀ�zc�����.���e�l��e��ʒ���-��$i�����:��[�:�7by�rN�TB�W,�u5�I�'�3�Bf]8��=�5Y���^�6�[.�z��yK�JH��y�4n5�d#8B8:�R���Oԭ_u�0�A#�.�ݽ.^l�v屡��UJ�5�_rA��)\�j�B{�vQNʵ�����2��O��fm�4�9�U	���J)�t�(��<n#<N���a���S�:��{�>'��E�â�{���s��*33f�2ӗ*�;��3� �Z������̕�Yu��̵�_���l�;b�D���I{�]W�DJ���<f~*����٣��.Ԙa;<NJ���Ani�=왥�G�������ԁ����;����[��qY��[��fa�"�\�uZ�`̼.k[|�'V.��ВYML��U���4�Z],�V:׺�[T��D�B��m��qG-����Ƴ�nz��UR>�Mb��%���c��"&czQ���3���wR�w1�45Q��rsrnkt;��>᫹a}3y���V�����01�@��v��gvL��&Mѯ)��O&Nu]!U���7�|���xr�#�R��h���X5l�Qu^��c媋WJ��K��Bv0���N������gAq�nėwT$+��o��ar�9���7͌ rK��-,��*_j��l�L�N������}s���WC:�೬���I�;��s�VKͽRG�yݘ��e�5�y�0����&ъ��K�����ݩ���W��9���X��bXMm�E�O����X�;0�Kkmܶc�-������Tf����^J�δPGj�W��k�P}Um���[�h�������*���%�-�
m�c����\���qs��t�6�H��;�n\�"-X	M��Wp�/��k�''gfCռVd�VhJo.�%�ew}4V�J��S�*��ܙS��h����"
���PWbќu���Ǐ<}�_��������"��0����q�#s"�(�r�Y�^>�<x��������{�&b�Q���db�94�@����C�8E'#��q����Ǐ<|~>>>3=�]����;�y��X1%�r22#p�b
hJ+c&���>7��
��ԙSM1U5J{�ZcAU���U��ɢ��*9�O$9�y1ne4!��S�������p���QEPm�v ��v	�q��[�(7q�[���� ��D�^�3c �%hk#%�)~�-z�'�AnlDY���lf-RҔP��lR����/��h
�ȣ �9P��66�
",��0˖�f���Xh{���bP"�m�*)�0�j1q2*�
cP�Rz	�0�l�L�#18����WgZ��!Y�q�G�3�Ӽ��,�B�������Pu�iH,���yǠk]!/ �/x�pQ燊7�}{caH���J��BJ"�H�(F��5�~r �d��)��q��!���3#�x���!F�p$�p�1R����!*0CM���hHaM�r(R��Š���?IRі�H�~͈Ca�)��A??��7@��=�
Y��&�}��Pm��Z�m�S���+�Ɯ�]�;�n5O.��!>qn��J΢���4�v&��ڟ��R[6�Ɨk�Sq��'��V�fVD=��]�aP+�e�N8�Y\�zC��E�v�c&K���aW����ݘL�W;x�}\Z�����ѭSL�m�x����f�-�i|�����_�*�:��ˡ��um��*��,�����y�֌<Z=!�^�-�z9�b2�Eٵ������imrD���w�&[���WD�4�Vϻ�Xny�8|�����6Qӽo�cu�i��n����V׵�����,���<d5�ǡ �*zcds�x�S33333gf�#ٍxW$;���U�q�\-o�1�;���Ә͚&[3��g��C2���+�������
7A�h�	�*e i�vGy�䲦�k�M��9L�����7&l�J�i:��ƻ�:��P]�rR��CF�}��w�z��$3�S�x!±wN 0����pm�:3����p3�,#��)�w���c�����>��߄�u�L�f�@95��ҫ���,�Jc��6+�s����|؆��Ϊ���z:m�<7&ٝ�����lL���oo 2QXH��C����ۢ������&����̚>���r��f[��,kXަJ=@XyW�gL�:�3z�~��+3�9���!�3�Em�U�@B.3 ��5�W`9z%��oE�g�Y�ZD��`p����Pd����g��ǥ��uc*���=�!�R�H�f���1�}
�q�+K@�;���s��s���6�۽=���}�W�K��>I]�6�m��*��F*/�`��Fh�o]%EwܦQ�����"��	���;��8"�{��Hȗ��Y����u.Yۦ��x��������cM�;���;$dGj5��>��I4Z7��bz���V��h��y�L�q���a�����0!����0W���fqWH<V�?[�'d֫�ood��Rӷ��ԗE˹T����~��b��N>�+n|Q̝�SFPmԼ����u�2����֖������ͧ���g`��Y��Ν`�*��]�b8c@ĝ�Wm�u�u��Mm�:�_}IajN����ڿO���s��-��Z����0�qC#�����,S�XrqFy��+�Bܚ���hVu�j͡϶h�~S���P��Cj5QB�9!���1�%kc�f�y�����C6�pn���ڈ��
�KwE�[�+:�U��&ݟ<l��)�<����V�xmOߩڇ�v�2C�mp�"��"C3��M����A��.���f��=QSЖ�n��d/.`>��˷���yҽ7��P�c<��T9u�MHE7c��C{:z���ٞμy�-j�%*�$���e7��Z�zz�.u��Fx�f֎R���������va�Σ�1e�)�Vw���G*ؚ��sr�&�д�������^�������\sG����a-�R7� �g2�l�����m�[w^�=x�������j=6��h�J|;���+iڱ�'���L�X�a문��OY��ͽ/Z#�;j���E�W���Wgǜ�q�ƖR؝�1���F�4]S)�dd�K��וǺC���ܦT���ݝ{�Ʌ��_���V��3�����ݩ�w�wMutS������*OF�R����n�g�x��z��m���mS.��%���Ғ�[��[zu�>X��:a�������AL�Ү!nn�n;����%��q����x�,���֝�3[��he���AGѽH��қ6lg�O=��Ȩ�-�=PO�� �����v:^����L� �J}Y��� k�hwi�<�W���m����ChR,"z�^ܿ?��Ԧ���0�;N*�-fGc�O�ya�zF�p<��%FW�݋$Gv�>�q�/D�v�>z�n;�Zgј�W���Ea��3�1Y���.m���6�dvv��=U-b=�֘�+��<p~v�]�BJDM�U�51�]q3<�ܻ{����}���o��Z�K5i�S��d<`Q/\���[e�r7o���ݗ�@^Y��Scx��79�������2*��M��L#��IOZ�*�=�����h�I��$�˰p�y�V�Z� b2ird䲶��U�؇^;5�{��}*�=�w�i9�����l���;��Rd��W��lm�/SXz��f���R�m�F��ok����\�����$}�xr`� �[	�7]�_�_>�q�0�DD�('�
��b)ûߢ%�r�ث��kۈ.�;�.�Y3�κ&��T�K�ʊ�~P#�_��ܩ�R�6�g�R�J�Y6K6�mf��ϖ��GMf=��ُ/x����)m��R��v|���똓���i}��s��5k�mu{كz��ܦ����d���i���UҪ��E�j���n;�\�q%��,�()- �l�{"��p���ݐ����Os�ߍ�R3��+��
;Uy�ܤs��<6�ӳ��fej5r4����ƌM�"9u	��]��͛�g�"�����V�s��C��t6���FEK.���n*�m��C��S33�w����޼���]���G�jѲ��333��^`M��X��`GY����r��v����ڗ富�1����k�=��f����.�_�[�G�B���a�4�/�C��Q�0X^[d�v�Ƽ��=�s�}��]��w5����KUEP�D|���(,����D/a�t�׼7
���Cg[���n�����N5�wo��:@9gmgt��j��&УW�w����{k�v#M�T+̧��S����ӱ�	��ݶ������Od��9�9���!�8d�<��%�`6��k���5`�E�j��`�w�$|��BT�1�S�ؤ<`�p�MI���K^`�teϞ6��J.�q�Ɍ��u�jٴ˫���lK,i�b��Ih3���)���L��^.*���/ٙ��$7�!25Se;֣�P��3.��[�ul3�2[.^���WS�=R��x����%�*��'�9ui��^nh�ng׶�S`�7DʞS�[}[�C�wn�}v�_Q0�P�v��`�}1�@�U��VeP+;�x˵�M]�UÂ��V֮�����o�`c2��]�p
�2�B6������K^r噫nU|���P����6�D=`{Ӓ<ع/+v������������Y�ǳ���g0������_�v�E��+�1K�~ܒ�:.3�3Q�`�Pf^��fR��j=�O���IV�T�fک���]�Ɍd\�Gl.���� �M�oz��Ogo{FXW;�Vw,<�+��}F�捷*��i�G�}���ھ�-��f��9�ݛsK�b�0������o�t�7!���~��.3q�IL��ޫ���I�k9��o7�x�Û�p����p��ίF�;��E�r�j����p�Wʹa�5�e\��\2y���t
�8Ӓ��c+��8b���42UT8�P�Χm������ɓ�9Rbʾ��v~���1�K@���FC���Z�7�߸Bo[4�>$���~���Ɏ��S��k�h�qB:81�2S�qx-�Thp쾅�E^�[b���@�P3Nms�Ygxx�w��r�i��n>�È�_dBf�N����!��_<6�D���*������F�-b���(Ƃ���6o{v&�ǡ�E����6:YŌz*=\�%�֯x+���ժW��|�R������f�M7;Yc`�j���U4��_]+U#K�ݶI�\o��6���㥶%�����l�P����h:�O�)R5�ur�lJ��8��}t�l�CVlN�.�Wt��,����۰^�;�YM�R7�]�|[�[�&�.s�Fe�r������s��-��G�^��Ț��]i�U���
K���x�(�Ҷ�[V��]oj��#32����\�ު�_��k2J����m�����N��!��˃r��2n(�<�ۢ{��n�Y�-�1�YJ�ѻ}��T������uu��Ӓr�ڭݡ�ޥh���O��עx�b���i��~��o��яKױ5y{m�����N!q����5��(�-���G�C�w�Ӗ���A,���}����fn	6�AO}ʟ?8�u��z��3��wx���Z��7��q7�K.;������� �:a��.x�qN����󶔩@ZS;�g��Ԏ:���E��3`�3���$���]V7����6&���:n7���F����S���y�X�DXټjo\(	'������݅���<�T��R0��W�i���<N��e�Z�fY�:���]��{2���z^|���.;��=k 7m��z=�z�R���tZk8u4�8��*��X�A1^���!�2$w�d���Uy���%f�wl��M ����y%35�;�:���������cE��{x�2�<t��=�a�--�xk�X����ؓ���=uyc�x�,T��B"�_W勲Զ9 c��Hq$�E�A#zD�r2U��	"N�k	�`�E�,�l9���B��U
�{*:B�c[�;4mOFj���sP�4��:����᫺|!16l�|AB^�w��]�I���/c�<<�s5�*p�6A-p1S4i�S��e� )X��co�9�\�K����2X,�}�v�U����gpuSX�N�����T�ꌑ5P�z��1�:���E_SW��
��sߓ"�3��f�e��k��C]�:L�W��C/fS0��������q������3S�����b�=�j�j����CP���P���m�}��ӻϛ�F�=�w���qq����J����e������ej�u`.�\^�ѭ��x���,�M���M�~�m�{��j�W�ְOl���0[��f���{TȸF-���n�u��;�3Q���~Xc��m����u��y������1�ڪt��x���y����vB�6-"�7Kߘ���lk(ޞ��9>�f]|ɽ���k&�:���c�M@Y
뤫S����:��5���t���n�׼>6�ɲ��$2���
1�ᒧP�:�8��z�ΖcǊ�e���_{���_�qڧm.��	��Q,�po'En��*�,����3p�8�`�`㩡���|�����:*}qDm�Ι�*�ی�OuWtW@��{�Fj�<Zc՞m�L�9��R'l�&�`s�J�k�CV�}��r�]M�X�kd�9�A�G����a�*��|6X2Ә��7Usė�2z&(ތh���ʶ���/��i5o �l���g 3�:@Vn���c���詧�ō��[ޜC����W��v�ŀ�Q�(9�T6T��V����:���f�)���f�"M�I/�m����]l�s��C$w2�[4q�T��6��^t��7��
=���R��V�K#/���O�(LVf+���|nܬ��ǩ�o"�z�$�
}4�5��{5y<�'���8���M˷^�99�}MY۷����류�)�O���3��\�����s�� �7J�V�W��j�ֻѸ�>�CS-�6�÷�%2X-'�|�m$ЙB�)�f_u�I��(��g*�����*۠�FiҞbL,(n�[*j�u-{���}��4f^�y)�͚�O���ϧ�W��^S.���#�q~����m�a��f�&I�OJ�W�(m�?N��S�ݵQѸ:�[T�=�,%�&��f���y��є9s����K{���y�f�����rъ�x�CC�VօBV� ��uLRڬ��VlfO�5�X�٘-82�2�;��銙��zp����7Q;l�'O,Ɔ9��8u_S�x���3�P��/$�v�e��MI�xޡ�[/;r�����St�V��IG��2�Y��yZ��Bo���#U� ��]to$j񲶤�&�L��@�����S��0ѹ���:�Ѷ�l�׿JB�Q��83D���sW��΋���w*co;��g����[%I����x>�,Ie -auy�t�;L[f��8���[�+v�����n��B�,�&T��2��}���%���r��;)Tb�cf�Kà�^��J�X�K�o1+�f�^7��z+�ZV���4C�1�����l"�=�SJt�M�>��)�'�#zEׅU��� Ƿ�CǴ"s5i��)��n��<I�R��F�v��pI��)�wV V��w��a�[�fn�7�Ygf��<�����JB,��Q�u;�8++�����&������S4�9�B� ��r|�g�TbM֞���8�$X/#�ז�dd�Y�K���g���]�a��%���Xz3�z6�v�'��s�9�ѓ�;���(�Z������w��T;�T���s�n���q<�fwn�l�Z��X���K;:���E�JiZ�	���0�b�^=�ۍS�]��M,n�.CfqR�D�x��]�uf:A�y�qKX���<���`q����F�����9���:üV���Y�v��2d	+wV��[{���p����n�47'Y|�R�w��7rc5��:|�.J��;:�v�M��m;Y4�/��z��y}��E��6qd��X=�
]��7b!S] �`�.��}����K�m]F�[��]�kJkF�{goBR�\f�H�j���.>�c([��r�{���=�ίj̚�uQ����tD�a�b�#�Wu^h|h���R�|{� �p�/0l.peLq�1��u��ۧ\>Ԡ��k	&:�(E԰�hR�ߢ�SԼ�4ݎ��QJ�����4�}F����c2�:�af�m�뺵�X=gv��QR[BE���l1�ƴ�(:\�Ļ3�Z���jx�����VCu�lb���u3�bs3/������rí`af�S��c��u�ǲ�j�9�O1�|콙�����태Ln�@��@�x����m�[�LL����N�-�����g>�O�<x���gǣ����#R�L������ ������l����I��aYefRr|7�-��믧���Ǐ?���>=�y�Pf`T@�fw,6�Ú�mA���@�G3"�z��O�<x���Ϗ������K�盡f9%[�Y9�	�Zh�� �-�~Y��c�أL�,̊��*,�3� Ȉ���,�ʳm-kwt��#�r9X{ݯY���XGpح�:��Q�DS@��0�>s3
��� $�,0(�|
�ϓA�lYt�i����Kl���¸Vf�n�Y4�n�CE�&5̊�9.a�͸fٛ��m���e�fY�YM��`n�o7v7r��A�p��0�r��h,���2(�y;���-�(���V�d��le3Y����l�UaQ��z�n��OZa;g�\,���(kw3pM�2�l��付���іUAATe���A�f#:m溗X{�u�h��JWt��T����u#6�6���@����국��1s��Ont-��xN�������ݯG��}E[�e���5t�s�s#]����َ��wwwt�
]�r�h�il�ٟ5�����OHٽ�S��1�'��އ�p{K5��<^V�%u�t�|�ck�#������=���N����|�aosSn]��ƏP��1/Y��F_�n˳;�t^<�rYexԺ�l�����WoA�_}�?�+W3��3+ӣ�<���ƺ��a!�X��4	��y?;�vK�ͯP�����iޘ�9���+@��4wn��4��kg�Sf;Q�����9��E��bgM���c7��Z������;�w|��1W:�r�y����q5��<�%Ş�Rޟa��ӕ�3���3FK�~������s]ˏ��o$�E ����44(�i�U�sҐM���7;j拳L��TCw.��w��+7d�[u�=:�W���N��\궴���R:�>�]�ٹ[�=v�D���b}D�uf_s�Ni�*sWN��"��S���܌uR��\{�QfkךQr��+]�uۚ^�1����} ��<{+
=�n���a��뵧�A�"&�ܬ��~v�����=�u]�.�;�����hq�2��ڛS>�k-e\Mu��״�ͭsΟ����&�~�h�M,���Ttmr���٠.��a��s����N��Y��{��:��u�Uܤ��B���*��Jt-��~٫-p��]�]�85+Mco1�j/r���K��H� rV՜�J�E��T'��ɇD&�LlvB�k�+;��=3�:�e)r�7*�j�O�9-FF�6e�c*Y���4W�GDy�ҷs1�3�`�Ao�Y9����Z+3���������qX�e��ѥl_H@�M��vY��󵄼������V�R���3O4d1p!�V���c�lz�w���[[��+�H���]�)�*-�t���u�
�q諩*-��tB�>��)^u�2c�Q��i	1����! 
�fdT����0V�V��B��]R�p�.����}��)��w��&��a*�Y�y����b|���4��1VgGԍU�N;w9�gg+4=da�2��]S����z�<��M ��Rf
�yߗS��,�ҳl̈�[3-t�m��\�^�p/�gy���:㘭y#kN�� >�5����-�kϱ���D�]�MG��"Ȉ��EY��/dF_f�(�O)�My�� Up~�@��i}{v�#U�6�}r���kD��5<{ֆN�֋8�y�2�t�~���ˍ�C��.�z��k��I��z��oP|�J��$����.�e��x�����Vu�����+�{u[��,-2we�;7ê�4�|M��t6��j��Z��P�2�c����dQ�T�X��LY���I��Gm�r��-�C������[��U4�6�gPI��!<����(j��j��T����Т���C����>a~�;�u:��(�VtP��bL#^�ko��B��z�w�dk������Ro�~�h���r�ff�@�j�����A���2?f�	Ù����9�o�m^���-u%_C5�k���ܢ��6�oJ�:��+�=�R�I��I4D`�<��X��$�g�Q��R˾qk�z�˱,�D�I�ܘ���3�h���E܄�Ľ�Kv��ŵsL�+�Wﾯ�v���Y5ݛX��@H�|�xҥ��W����)m�劺�X/wF�ݱ�v�G�jIŗr)^oU=񺖷����6���ƨ~����}z�֝j- �wz��y��l%�%,�
KA��f�m��C�(���x�0���	:�4��W)O�i�.A+:�3o�4���n�&tk�̶mk�]�]��x�<z�	�ޯJ�fji�oDzVl��P�.���c�2�܊k=��%yꑦ&_C��Þ3�T�ǟ:g�x�
zYg����X����/�!F��_���r�%�;<���c$���ʇÃsnib�#�<�i��i#�rh�r�������:����u�g��7��յ��y
`9�Ov �����Va���s�$�=26��dܚO��eq3�uc�ωVT(�Փ�v�o���)ߎP��^c�[�4��Ӽ�r᠜3�7f56љw��*׷8�6�_�p^4/�,�W�Z����p�`���Ov��:�aԢ2�p���>����ޞ�v4㔻���vڊf��kn4�u#F�3MC��V��)v������痴/������#kx��������n׭OH��y!Vu�Y%[W��lRz�_c���~�vjNKZ��p��[�O���P�k�SRbu�C��w`���qg�2�o[=t��~g*���x�L�*�4�Ecgh]vM\_�5`�z2�%��
C�N�����^�e`�H�W�v�5s��S8a��r���z���h��eVw8
Ǐe�(�bK^��,�bY:��D8Z��˙�ʼ)wP�;yc-J����ШnI��ji���<1u�B�-�ۼ�Џn��e`��x����׃)�N\m�ֶ�4/%��欴���6PC� CLz�V�N���z���kk[�5C�UiQ���^�En��hȱ���D.3덤���0��T�ެ�ƫ��^A"R�;cVO� ga�]�*i�Q�5��E���U�e��%�Z���P5fx&��`^��\�h�V����_k�
��P�<�B'����j��v/{���'�nN�@F���O�٭�z�b݃+'D;l2-��vg�z,LR��n��X1����ay��ԛ:h]a��'�<�ʪ����Y[�o=��s��}"#�[0n�u�d�ty�;h(�wl�������]Dڛ�6T>�fuݧ*�6���6�O�#�2^��hx�����R����oxL1�j����`���M���oi�A��T�_���\s6V�,lK��Ԟ+�ءK�s$��;<�g�l]�rE�fދq:r���s*�^�>~y�{�'M��
�����������="��O-/���S �������cύM�C�T��bk���ꥊ2m�����WR�ݽf�<���m�y�S��7�UH{5
�3��z�a���7(���2
8
'�hs���e��6w��ߩl�8���Z���S���OX.]ٍ�v�%+Wx
�����_*��;l�����}�Pө�u]�됈q+���|R�^�Y�F�}xȸ���y�[��q�G�[{��q��CN,�H\�2)[&�f�c��B�͊����
�(IG����z(�چ���pe-�3�=�l�L눥z���r��h*J�	�9�Q��������г�����(�(M�@�.'7]U�o般l��D�$14�NHaf<��UF�8��o���ղ�o�����uaq����3Z8F��99�G��m�Ց�t�'4�S�EF�.y.�#�m=�P#S�?P��sۣM[�C�n�/+h-ܞG�vؽh�@�Y1�8��.����imÝ��h��ooE:�+� �NVp�,C,�uo|cbv��LL�.x���J�d�yq��R4�����	��ua���m�����[�Yq���}Ī$�܊"Oc{'�%�^�\M
��9���J�P�q�ГKO�'��*�o��Gq��K]å"l-{�y�O�:b�����4�w26�NlϠ+2,_G�c�M]_m��H�s��g��D��|�=�9I��}f�a�!�x�����f��{��C�#���3ym{�d�5��4�l�՝L��c��1N�4DA�SY-O����'�T-x<i�si�C*r^Y"P�tF�����g+m%���p��Y�Dg?9J���ļѷd�2h��gv���u�[5��Xp��Ti)w�v���{���g*mK��6�8�J%]!ݳI�Xp:�\B�v�[��ig�nj���̼=�7xf;�v!v��S?�#ȪD�9��U�y��u9-�1KG�q;�iY��J;Ի��|I9��뇻�J&Q\�	�o��nr�[��7V����ת���B�Y�}z4�q���uS�Fu�fp�!��+h�{i�����Tyh���~=���R;F�Q&���҅g}��8�ROV�p�7+�W��u�s�j�Wq��H`��O%��Ѣ��7K���j]�8ED���uz��W`%K��E_U�G����M��SW6��[y0�|y��;+o��ݼ�=#[͚u6���Z�v�p�2�"Dp��k\�	΀ G��0��y� ]�v�c;��y%r����ϕ�/p��-w�`��W�]���<צD>��[�����v�BEwZX9kh������^�>��4��ض`�!P}�9�>^��T&v<��#>���CU�Σt,�P�>�52w���E�=Y�8����C���J�iIn�ԭ�Zڎu�㖗JQ�n�m�-{+W_�eN�uJ�ީeP���m�����wyWD��K��~v2;����xUہ�n�y�]�1Sz:^�7��%�axxg^Y��*�^׉G�t�rj�w�p<`�jb��UL���zf��pf������=Þ8��9�yv��@��#�������,�=�5s4�K��U�=�DAէ�2.���U�5��ǯOsHrs��@��є�x��<M����h�0�.����o�i͞{=\[RA�T���ٟ���.����-��I�8s�t8�B0�\�=l����$/���QY�	d���s#r��{��/:-M���glr�u����|���4��mٸ�cL �@�D�8�O��k-�Z
�坜��֦�>?�/w����x��I�s�
��N��o �pơ�&�˜�Qq؆�v���=�ي
��c�R�7$в�(�L3T{�cȺ^v�b�YN��0�6v7t*x��5��z��>��#zR&�j�YA��z��t����{�o��1�d�����q�\ṵ�q�9^�p��I��e��i7���9��wH���ͬ*��󙎸��,�i�.����+��f^m�����/a}u�1�<&}�u��z��/��@��m]���T#�\3�=�ݵMm+Ic��.9u�[��$=p��g7��<��İ{���5��s&����r�^�����6���lxKdAm������F���)�K�61�̙8�Pb�u]Hj���2��=.�K$dx�e<�������u)�n�ۭ��WWj}&�[7���n���~P5d��s3�<�:b��Dp+׫g+���}�G��<d���>j���Ne֞��Ƭ��6g�� �9W2': ���$�t�X����1+�wiʳͲgx���8�c�uV���r�P��7�VȤ�����ԍ�a�UoA��=��Xl�Y����C?	�p��`� %+�� �g{7�0�xh�f����*l��b���~+X��ǲ����as��f&��1꛼�ۊ�����7&+1/qћ�B�Ё��0�y����}�������?����QDW?�*�(����a��T�>��{4=ϳ����X"bC����!���B�@�! ���)!
�2��2����膀"�(b"���)���*(b"��h &`�"/ 0BE �%Ps��� `0BQ �%��	�!T�@!	�!��b(! B!*�B!"�B�!�B(!
�@�*J �(J��
H���B��@ 
 B !
 B !�B�! �B(�@ ! �B � B�B!
�(C@�$! ��(@��B�J�!(�*B�L�CL�HH4"B�0�B$442!��0�C ���B) �	 �0	B�440H�C"���C$*@�(B�H��������=߻�PQQ�AF�@EI��~�x����|�O��������s����`����B�c�L����d�������������*�PW��J�
��?Y U����?��I������~��C� ����?g�?��jI���>��?�'������aY~�AUeBD%�$BH�T��T� �H�JUY�I�dD�D�D�T��Q �	�J$�	 R�U %BRU%�IT��I��H�T��I	D�$B!�HY�$A�d	�d	P�`�d`YXF�`a	�e YY��e�	Q��Dbf�Q@�	
 B 
 �R � �4 %"�P	�2!!H�
 @@$@�B�
�LD LA�$��	�I ��Ȅ��,(HȄ��LB�$JH�$$(a��0����/�'�

4(!@� P�"_���W��߳�
�?��?���g�Q U��X��o�����bW�`�������N��� 
�܇�����>H(��@�����~��*.~C���E U�?�������оh``�3�='�t�><�q U�D?��G�D@p|J�����?���9���?��$������DW����(�����~���R~�������>������@�>�	>~�H��������?�p���|_�w�� T_�x���}q@E��_�{������!�����e5��{( B��� ?�s2}p#���ޢ���(*6�Bh2-dJURSZ���"�}��T��	v�IkJ*�-���UU))T�C*�V�T�0�TH��6�-Y!��6�iQ[5�mf�l�7��R�^�;X��45�ǳ:��[k,�Rkme�ڢY��Vl٦�j��Vw;�٭�U���Ŷ���4�j}��Y�iYZ͍��&V�a4�6��m��YU���[}7b�-���l�KfY5-l����ۛf�e
��5VֶƴY)jIV�	�d%����a@T��  ��S5��kܵ��T���j��V�7X��պZ�S���O-$�{ۗ��$��L<���M��5ڥWmۻmv�����v����k���Q��[^��Rz�Ń1������  �_q!E
(P�C;���E��
��B�l(�
(P��nN%���k��彚��z׽�k�[(׽=nx�n��r��O/bu����77���S���t�J�<<^����[d���[Z���|  ��5����S���v�C�:�W7zwj�.�����l��p�vݻ��Z�������v���ދ^�Mnzt����P3w����-��s���t�wMQ^�6T
�X�1�Kl���  7w�/m ��yӝ歚��⻊붸j�Mu��Pw���E�U�s���e��=��w�M*�=��֬V[���{*��:ev��J��^�L�խ�ҋZ+f�c5Z�  ۷ڒ��b�{o�c�z�����=q�!As�x{��kB���ٗNW��5ESn���ճM�׶듻F���og�ƕV��]vk�!f�Z�L�UM��6�  �覾��w��Akǻ���L��og&����֍ݗ������<��ὲu��:v�d9N�kCpN�6�G�zM6.ڝw5V�ee��   �\}*��}w{֎� �=�  4 	�8  ���  �� ����  7s\
 �Ӏ  ��j��6��5�e�Vk+;�  ��  ��y�  :�0� :��:  u6�  ��4��  �9�  l�  ή� ��[b�� �la��5�f�   ��  <h`  }��� ܠ@�W  u�o   �`  ���@��  of�  �����V���Y����i�3|  �| �{�  �5`  mv㦀 Kn� C�� ��` �W� �ۀ  ��u  |���R� 2 S�0��� ��5OOLMU(қP E?�� �S�'�*�� ɑ��&eU&��������O�>�~�47�o����=X�/V_r��l<<+��`�9hzP.Պ��U}_Wԯ�s�������UE?��x�"+������������?o���Hu=1��#ߡ��y�"�!ܶ4��(ȓ�[�p�p32��?��[�4�p--۹����Z(U�iFᗎ�v�,ڷ6�FT�Z�Z�l1m�n3�@��Y�����Wr�Ԕ�4:��Y��x�-�7������6r�Xt�J͛j�=����mܚ�jn�yQ��Z�Ș��V�C���Am
����[&������+E\˂��:���TD�a��F�Lz��?��S{1�i��D���Ʌ7v=�uS�X�B�"f��ܙB�AC�tq�t�����o�p��?��<�j(�3�6R,���fӊjZ�Ḟu�ek�0Yb05���%�[��7�v�Q�y�@�Q�`zEGhE{Vw7g�]��;�n[t�N�ӈLe��e���M�T+!�=�j��se�\93bio$�� �Uv)y�y��*`&u6����Yb�W���hb�
J	�Y�j�:Ȧr��=+q��������uf�V��0ݤ��(�H��p��1�4�n��e/6�ݷ �t$�� ��j�d���Dڶa�5ҩ�8�A4	Kks��spnӃB�%9l�v��֭��]Y���er�s]d��B����r�ԫ@�V�L��
�W[&��e3H�Xr�4fh`Xŀ���V5a�.v"{u#PZ:ղfiԲ�;��`�vU�z�:5�j�֝Y6��I�z9b��wm릪��1�I�dU�Lf�;��ϣ�UxdMaW-�ԡ����7�x�����E�^�� ��i�e2����$z)�	+%?�[܃S��R�z��J�,,��hI�X��l�o%���i���h��ɉw��rZ�fJ�,yh�yE{Wd����̔���I�ڸQ{@�X ��/a	(`��R�N�نP��mE��d1�-1/�*ӭ��G'�RW�dM�;n0��I\O,�@M,���wz�u�>�VMI���~8�����ҽR:�w��X�z1�XF0�!<����$FoAĕ2�!�1r�I	)�w� [�RT��-S�j�Z����2������t�t�ͽ��B�r���
��n�<9m&ƻӑ�TL(�
�C�Mz*�H�,^õ��ۺ_��ױJ��u�l��EM�0��Ed�M�1 �H�Ⳇ]]�OkQ��Q7�f�t�SE�x�!6�w�b�8�ZSuۦ���
Vے�-u�d9r�h�,��ܨ�_V�x0�NX�ۼ�%�������"��A�:��p�[&�n�ό�C�pbËįn`�xl@�� i�M�)�+��9U��F�'��ڤՆ�I�eZ�zn雽D��C)Z��F��OE���v�jX��ˬv4����q���t�;��3&SoV���v�*lU2d��n6��L���J��{�sFa��j�Z��ڹg1hN[R��vP��]=��Ī4F���;a���j�X����ݕp"�.��d⡥-�Nbԩ�Mj�V�j�3,!�����sw]i�b+�v��f�ܲՋyE�M3�"��di16�$��"�cco���6��5�ϥ
D�Yy�=�eM�`�/l깯e��!:fV�L92��v��ֳy��Y.��VH9(*q��&��a�RCHԸ�9e��ƂTq�ap��R�T�Α�Y��Rʂ� a�J��L�]6B�n8NKq��AB �*mP��`^Fd
lX�ډE�s58ܬ�,@��R#Ijd�@,��x���kHé��ĕ���.��^�����%W-&��;Y�SX�t�Z����4�-b'$�ڡ���~Z{ܛ%����"�95��qQ�[�Yw��@�'5zbK5.�|2���wf�[�gD�/K3%�p�o%���5\DLźl���"���;B�
��Tvţ&jȀ�7�Gbn����/A6�sj]���&�ǈ�JV�F�eJ$P+��Y�C%��5�n��n�@HH:C^m"�X�͠�Z72�R������u��CQ*V�H{���P&�i$3v/XYZt[�hQ�!�YF��Bݽ�ݚ�v>1:���۔�p3	y�8�Pj���2�m�EGa�q�Xc�"�v�"��Je���lC	��]Y��P����V3b%����h�C
2*xn�jJ
�Gu}�ƗG)�ѷ2�����KB��V"�&.��w5�N�W�*V�l����Ge(6J��z^�Ȁ��,�\��Auk�[,�8���\�2�N���sk����ћ�2V�D	ҥg���t��q�5ɜ�]ga�[��w&Z*�,����Ck�&�����eCp�y�Vjˣ�#b�n�����5�I�p�%l�]�G��Isop}%dR��Hj�x��Eh�1;�m�n�Y3c)�f�'T�;����"�X��ayZ4l	�Sy��i����,�io�]���p�9��;�*4qG��$��n1�f��z>\ty���ӊB���Y��Uh6V�,���Yd#x~�%n��!��:��K�wNR3r��IÈT	�7�0U��w�%��Fѷ(M���Э�~����/QՔ˻�������6
F�A�r�����>�p�x���wHJ����l�#�k3f���� �1tz�q���29M�U���� 3Z5�ikc���ˮǄ��Z����u+%!3Ql�VW\��sF�i�,T֫Dj�X����fhLVǗx-�r����ǱB~v�N�J�O[�.����q-9��f(�ux��G.�#5֠�Ld�8U��6�M� �S��F�L@سmm��7n�D躀)G+��QIy���:c�A�En��YUZ3ifh�J͍H��0mK�]ja�K6�8��+%j�V%"��S���)�2�Z-��#ĩLT>�.�h��-<Y0=l��¯R-n�y�Di�ZF㷑��%ܼym۽*a-�(i�F�*?c�"�$��7��gŽؓ�,�j�;�R	WI�FI��r]�Z��[BDqbNF�Ɓ]a�Ch 'r��+v�JSZy�3�)k���ou�-�k4�`����;s��¯��b��e*����Ԥ�q�t֫K8i\R� ��+o�^��K�ӗ�@���u[Z1��,��m=u��F���]B�	!w��� ���n��ƴ$5�x��$<�*� �U�F��y-<h���dt��N��I��ں{M�t�-+�u�)�aٟCxm�2n�i��4��c]BP���u�[�M˼T�d.�
r(��-ӕ�����1[�ܽ�5�X��KTva)ө��.��`a�z��L��ҥ��JBЬm�@��2�܂+б�+N��s`�p�Z���Ʈ*?AP;`�4#��n�K �a��l�y���-�����d�pV��E�Fj���x�ʙ�gl�HӸR^#^nF�-�Ŗ� � p�ˣQ�6݃X
�{�f}r�;�E;�83�G�dlB%jaJ��X��uH ����齩Lm�Q��(鼦v5XiUݱBnI0!� �-�vY�v�*Όm���w�TW�5�.`�0�Z�;�F�<�K�F��X�P����P���@�{@֩J�)[�����R)\9�PWՌ�fFS,��Z��eG��ܩ��2����TbG7tY�[Id�@}gJ�x)����/)RYI\d���낕~u��qmdB�SO���� ql.呇6��	����ؤ(J�t����:v'���(1l���Փ�`�Q��*���[��k�t�m�Q���i��7e[���6��6j���-W�IebpL�0Vh�(���Բ�y
�EGI�5L��*;y������5n�cz�w1�`����TT��r��
����Ҹl]�ٸ��J÷Y��2]I��ޖ�X�A.�u��MK� Ub��G��M� ̘2�q�t�v��"����v�vvf��Jnf�Ě*�݄�&km�ך�rL���^���k��H���",�37Dr�Re�0h�b�і*K�7�[J�#��+D�ޢ���84�&���N�-&��о_&�[y�h@��<,7+76��w!�d�	�
�lux		x.�a� k�<�%Ŗ�!�W͠��E@��lkǷ=���M
"�H6IWF��i5��[R�bD6��%�,���Yv���.�IyWT��z ;w�42��zغ���lI�F��Jf��gRR)�@��JK�Kb�!E�PE��z�#.�S���m�)V;�/i���Elt��A���������m��f��h���*U
�jd�	w�A��H���u����P&��F�̀�KC�ʇ`��r�̃n�]a�jT�1�m!�e�-�v,��}z�Vթ�<���-ص�4 ���Y�a��/ z��ݸq<e��Am䑧Sh��"�oJu�,v�1[D��75b[��)��	��j�Δ�LIPDK��.��kUB$ɵY���g.+l�3~�t��an,�r�������F�]Y�)��8[�n����7 L�*7o)K�J��Q�ѕt�����F��d9�����$Sy!)Y �Ť��(��e-�/,E-N���)����P(P�n�֠i}l�ҸwB�F�;���j�ONJ?7/H��;Y+&F�C�+DyY[�
���T[)R��-�Ҡj���ޠ�������Ik'VVڈ1���c������ll���ݳ.6�{�ɠ�]72)��,�����f��t�b�j�%eBC��Fƃ�C@ݽ��ʰ�š�35�E�yE����hh�7Z�=@�	ތ�h��Q0
)�z�7SA��f�-�YII7��'i&��v·x�غ�u�E7rlh�+):�]��+�� /4\�oX�VȢ��,�ʹ
5
	�ZF�J@�b[M,���-	�!��ݧ�J�M�kkw�yM�O�d7DW���|��Nv1ڡCKX���<s���cД��b�����35��K͵��]�Ӡ�
W[+v0���4��HY��f,��R��I��Y,��sVݪ�u��s��;Z�����*�#(U��A�ئ'ί16��MZ��&����U�YuvlM:V���˔j��6N��rnQWE�U��N�� j�/U�Lj��4�@=11fJx��k���J6SfM�(Id��z�=�� [hc�{aaoe�E���ѢM�d��IG���1h�&���3Sg�l��V���lp��n�"�������F)n�yp�"�u�K	��õ����'�K<ߑ4����m(�4�0}rݳ+nTSJ ́ɻ%m�c4�x�RrFM���q
��e�ë6:] !(�%���m��a�`zj�?�hz�Yf��w��S��lkQl$���dPyxE�)�e"�&fV/
�)S���:�z0��b���x��|���yf��]���G�a��X�+a�5e�ܬ~�Cq�8�B�r!��ё|�S��ZM����(V^S��KqX�n����`Q�4,�������b�4� +���c)Yݻ�@�V���v*��#H5��7&��!Z/"#�жо��gk��w�<У�Ä�-�«;,,c�2��X-#s�-:n�=�4.\��"�ț���u�LOv�aS�8ݵL7����eb�hm��R�U�[x� Y�yCr���xȸ�͉Y�[�ͦM�CԹdiN��m�4ਝ6��ణ`�tÕ�GN��k˦�)QK��;��;������2spv�9!)Eor�S�F=��`�T�Lر�US��fb�'`ʨ5*���m;�*:�B�gwc���VZ,�0�����^ni���[�<W�Ba�2��R{���6�o5+YeYܤ��=yuR ��C �M��.Kɀ�m;.Dr�0��57��ט��LI�[&^��z.�U7r�lv��Or�1U�s77b�ME�JX������|�BԞa�1��JR踤i����9�A5��j*&�a�P��`�-H$v�׶��c�˳5��^�w+V9&_\�{���di��K�����}h���*Vn�f9e��V(� ������<��bk�I���-N=�*��/ x�=8�l674��k�4���2��M��e-��mq�c4sEu�An��F�א	�c����E�F��;�dj��e�j#-���;����2�
p'Q4ح�P˫pʽ���jXZj%��DX��H!1@f-͢�`��`�iC�M�r)�Zu
�6;̂2�uEI��6D��cj�cV[n���.�Bm�Y��W���l�3�e݅RF�ƖZTV�r�$)Cq��D9`Y!�b�oP@��V+�yC5o嚵�HTz���.�R�Ui���\2-�(��ҥ�f��ڒ1��ص꿆�L��l�m%W�(�(��F�r]M5v��Q��{70�
Ѻw��u��+R6�n�bU�L���	v��&0qj�����񌤩��������j-D�y�N�x	����V6��(S�y����CUlz�b�(�ݔ�Y3�v��Y�Dm^<�v�K����1f�kRAP�低�ȱp�̈́�˸�RŌ��Uv�/oj<N�$�a�nK;��a���EX9O��h
�1ET��r����a�Ķ��G,慹[.#5�ʆ�`�h�6�&w�Y�X),f�V��O��
�df�;xtK5+AЕ4��q�녝�8��v�>�1oǦd���<�ǹ���ĝ���b�H���S{��l���Z-��)Z��U�.�ml!|�Z퇨=LVt袄���_�1��L4�y����du=��E�*������u��F�<��s�m���(gW�V�o���*JXN�Y�꾑JW�Ҙ�hJmva����&j��{��®��ۖ��]oqyr�U�m��r<~��c�:83�Y�����?N�-ݵ )[U�#��Vr����G�h�cd]��9թ��v��뀖4����ۗ�i��3��h��Xa�c'���dӓ�Et�^�s��ג�^��A�&F�m����dJؒG�Tѹ��� [�iU���֚�d�4ޣ�r�NJ���Q����^��E ��x���ϬX������x���C�&a��b3/�z��
И������'��[�mCI�η:'x��)N����۵75l�u�"�ʠ[�Lޣ[�8u��.z��s��D4���.��T�fp��sQ��e쓪:��C����=B��"��D��>Us�6�s ��f$��K�^�]�Ҽ�h#��7n����h�v�v��3n\g��2D�X$�9��,�v2Ǟ�t�=��J�[�����oT�a˛����Z{u���%8]��2����KC��Be>;��
�����u�v���Wi<Y+��#�˧�i�D{a���&!�������H�+�����AN�)ޣ�Cj��Y�ɾa��t�Ӷ31"�;�x�t4:0�s�o���}�	�����k{���.E��8ǫ�ZZ,���<�8�r�w�����G�7Z����|�-�(���p�;N�H���5�8=쳕z�ĨPVƢ{ 2�՞���ՙq�VFjNP�yN�N�(�ʀX�N����Ҡ��_ �������=�d��&_C��v�Cct�-�G��ѷ�A�����yݤEH}\Zٻ��!\�V�gF�E)�=�GT���K�һ[�/R)�n��N�g�� �����J��|���v9���ca�t#�,��o`�|!����n���FS���^�=��8z�pw��%�������dt2*���L������<E��t��=�@��h�#�urΤ���qv�p�XK̎�0�zŠ����у�k�4Ɯ�Fu���Y��8�ƃvl�MR���vУ�:�٭t��d�"�}R�5�x�#	W�l�P
�_e
5!�)�N.v��L���YC4�XU5�ç,s��7�%��'5�!�h˜
���^�B�D5k����l�5��q|�	�C���]Z�RG�fm�F��S����\	�}*t͐�km�(����^O5</�31�k.89\�^�O�d�z^䏧C]��-�%��Z��u����l�o��xJT�&�ސp�Z)`�gfobR3�U"}�fI����ٖ�f�ɒ�y�ٸ������������6�f��cLc^�);o��S����uP����k�//{o&Ҁ�+�f�:Ғ<6Z�n��͋��/��t����;,E>���u�
IGk�.l��� d+��8/���}���m���|��o[�f��ڈn˃k�����s���֩2�"Ƴ�>���YEr���E�%�6�Wz5c4#^�7��WZ��ʳn,��!�:9c�%��6о���_W"��LoE�n��H��C����������ME��Mk���!����̩�ۑ�M	Ͳk�q�·�7�tY��X�.����G�c�` ���Żs3��G69�B���Q�h΂T�:�#�m��?�z�l�;��'�u�W,n�>��cl��$'e������;w�﬷�C%޼C�:��ٙ���R!ϑ�W�@��	*'��g6�n���K*�NY�;��2�}vڵ���G�k:KNƨ���W����؛�����@���a����@��j��'E���֦Y���Q5��ic�A�]�Eb�C�7�2���E6� ^侚�:O3(јF�W7 ZfB�\�Uɲ��#Y��w��^�u��Z�.j�p����ld�Z��:�`BGU�e7�Es����P�iM@6mg+�h��V6�`6i<�h�ʌV���t�6�]<C��;u,nf����+�UN����(�����W17*�,RbY)>�fޒp?�̸9�4���th��C=m7x�e�yfi���Q�+Z�g*3s��0�8��갫��������������ں�b�k����jy��[�7O��w�&Әn��ٵm]��stMY��p�m�t�N�wyk]�ۡ�vJ}C�Ǥusd���ז���D�9�������3��3{7��Ӊ>t��h�zB;.�Rx�L@V��!�qeav���ͧ�]�k9M�t.�&�e��gZ]/�!�E��폷V1t�gMB�b��z��/���;�kV�r�۾�1Wmf4&M�̴�n,�Xul��W����X��h���ܼX���K�6�'��4�&�c}7;n�Q���n��{�}�=�V-��3ͮ�	�XAg��<���$ٶ�;$m3�:�S5S��9�;T�uG|���`�Tgo���Wb�ή^��׶��r��4mp��nK��"a�ɓ�*�nq�6�&	2/���j���xfN�����}�����v��`�d7zW��j�m��+�=Ɋ%X
&��)���h���}�᳇4Lݩ�����D�X������k}���|euf�Ֆ��TP���NtzG��a�}Z�e�Dd�PT���QL���+k�K��|߀��<�%�a�ˮ�[Z*���	Ԥ?$���H��YF�o1c���D��U���!:��s%M�]C4nX��Qcip�2�4���L\��y�P8w�
{j7ӌk���u���*nf���:�<�pTCQ�on�&���*U�޷�ws�Ǣ��N�Z����sN[{kt�Z�z����Ff-=�2��z��j��͐��<��U��3��4P:y���v�J��{K��匆W���0r-;-ESe���w0t���!q�j��xv�U�0�j ��O��Ͱt�|ʪ�|l��� �U�=�l.WoZ��ǎ׊\�˷�}}�m�d\?,�������G�9Yr��6��kB�r��r�\�:�=_SF)8���ܞ�q4�m��X��%����t�&����n�����-��x�GC��4�-=9��kA�<�����/
�i�N	�j�_r��IЃ�q�$�[�o��{���n���K\�n�/����@�t�:m�@�KKLE�h�Fnu�Z�-m2�wjrW:H�������� x��m)��y�� �8n5;��K���p��*���'(�Uv��508��[�)�ú���*k2��S���_����Hp�J�ru�y�v�)�v�<p�pnj
���2���]n�34�k�E��S@�] ���T�G�E�?qKI>D�dJG�[{�J���ڥF���7 �hp����9sdKqH�8�A�u��f����n�S�ų�X+���3A��Y��q>9˾�&�;�$�����%�v�7\�U�\+���c2�=��(��<�9Y^�;Z�s_�f�X�\$� F�'Pޟgi�Op�r��%_d��������2�J�TQ�w���� s⛻�w(��kYZ(�ya�#�O��ڬ���F;��O��^��I�{�f�"3��	|��H�g��͛���:�a���)}���eu�:�����Q���:+�, ڶQ��h�N����? :��Z��qus*2�>5�E�͵�u�f�b��.v>M�������5�uv>8]�>�]�`|�U��D{	��Ǖ��PKV$���١7N^D'm2(X�����.`�o�گ�g)fY�dE����fe��5Ct��B�΋*��.�i/0�J9k"Y��� ;L��Z�n��OIQ���tX,uM>ًT6��i��Xq�e�s�w�[���oZƬ���P�0� s�\(�lşnę-�F�Y�)IC��O���sP�.��Gu�̿%|��e�s��G$���0p�Ҋ���V�^=1���uꝻ�y��h�HIq�6@e���&���$��јO����X�7���ӤI���u>���3�;M���^����T��;�m��B���W�.�����Wcq�}וRr3�fծb�R5��x���ۗ���s{!�۲L����e��&�`���k�~:���`4*9��x�]>M�����L��;h(�����I-<)ã>s��^<�K��T��s�r9d�֖J`S���l��ᩂ���s<�`z��癛#;r�뱱�'x�þ7rDu.{z�MK�_tuk�L#u,U�ʸ���&)}�,tx����1���i�9rTX�o ��4-��*[�rR����i��=��l����ۡ��Rǻ��:��(bkAf��`PoM��0D���\��s3\�z6���8�1�k�e�^���Q3x�}/���-�T.]ƕjm_�L��&¸`���[:�v{���z}����^�g�#p׬_��JH;~�˚B�d�"h��z�0��X
��Es���ۏ�/�6�K����۸x�J�m���"~>��Sd��aw]����@�7&��N�xhˈ�t�֯r�p%�z�[�:vM{3m�mk�� 7�q�{�����ZE�����m�f��V�6�Ap*�t�T][�vJJ���C�H��3'O�I�6�4r�A0�,>̢�a|'�徼��.�!��9��+r������\�Ú��c��h}�u�f
�1���$n7�V�SQ�u�z�ы��{�����m�d����-]����kS��m]��Y.2�ǌ|V�H�|����*MV6�&���y4_qRl١��7����J�u/�gJ;\w�F�8��0/N��^(f'�M�wd6�tzk�x�#��c��Sj]]ۇ{0��k�	���������V�S�!�v�C��.�{�рZ}�zu]��{�ש#N�;4F�]���{�-��{�ů�-8�+�]��0�1�e.Ε�eQ�����N#]F�#����q�� ����F��	���a|6��ɸ�WVeX���Ky�ٍf�����9*�ZҥY��3��'.�ٲ!&���>`K��1���85�������`W5�y_�fd���DC�����Y���&�4��qz5>�v��x��ٗ�}��%�,�oZ/YݽG
�穾����74�@6LA�xu:4-������]�ܪd$�K-��1Gs+F�-�`�[a�;oa�d��68h�b�S�w�,+����)ٰAf=u�K��VXQ.U��w���,�8��m��',�/)��BS�Nb�U��e(�w̺��vs�'	��� x����h�OϸC��Ԕ�.�k�c�rnd1���|���<�����'�q!�{ױ���Kaz{���S��d�:�9�����1�f�,��v)H�I`DR�&�K�Qռ&��*�l����i;�c��wK�6��:�����$.���og>ݝ&ޭI��[�&�ݠ��i4J���.���:���FΒ��Wp�ᦾ\�!��ɻ���8GV9�)q��L��W��Y���Y�-��o'���c�I:ӏ�Y룖�ᘎ����=z4j��],Z�ޅk��d3k:5.W6*f�E9�ƫ�6����3o`̻n�<5��� z��m�Gs��k^J)JE�Ql��'���J�U`�l�Ժ{0E���w�H<���+� Ym�h�����g,�e��T1'm�<� ����t��|�$�U�뤍�0>풬�z�qEg���x�fj��*�q?m��	���u�[�F{����ɝ���BK���sە��-��_[n�9~�^�~�!�&�w����g���<�6�m�D �G�.G'i��m�9�J�붆p�6oU�{;И�$������K�^c[|��`���pt���ѷ<,��as{����1��-�sn-�#���2u}˧e��S/W%2��}l<�M���V��nMݪ��j�:�ŧ	9'u:S�h����>�%�:W|�.�]h�{�}}Bǐh����D)}�kVUi�rp���9��ƌ<S���#X�$.T� ��d$�VlnY��<�.��qZ�='*t{�1{{;g-
��)�'��/�Y��K��jB��kf�]��_=\B�q�;%j�@4ұK�pu����;���X��>�F����r��D�*����ʹ�]B'3}�V�b�F�Cvr�+��=�ܻ�̉���];�]/Vvt%��b_=J�e�%�ȹ���J��p�[ǳ1�-ې���2Ɏ�t]65b���ξ�������rr�����{{��n���ܽik��B��H��uf�y���
�}Nq�k�OW���z�θ�ۻH7�o�9I�Y��ʛ�Y� l��v�'���u���K�+`窍컆�,-vS�Ƚ�.�ȺLXl���rL�d7�V��o)��M���C�N	bj�����{5�K)p�CW��jK�,�ۗz�qgP=���8y�K�p�3ǁ	ǡ-���i�]>�V��(�n5@�΁��>��fW%�#{���2Pd	UQ����jб��\X`�n+7yB"��]�b�+���\oj����V�:�z�~Vn���76ތS�w������\�.�~Ȏz-�wʟYD�mǏE��S+CL�޴�*Ջ �F��xƒ�s�4�)�ݘ���2;��z��23�L��S�����咞�:s�%^�SR���.K��<I��9���lou�n?k*��9��������]b���оѓ�)�vb���w�y�N�2�Ԫ��H���<�<k���<͌��e�X<{��@H]���2C�� S0&�vuw������k͓a��gn_��yO'SR�oz�����;��I���Xu���r�����o�y��}��ο}��TEUE?� ���~��WS��W������\��bph�����	��Q
+#I�v���v��쿜+,<q�eSZb;0A��rwnb��+�r���Mo+��]����|;���R�6j&�U�Ϟ-�˜���J�yk��nd����L���f�*L4j�d��-�(��h�z\O��{�c+ڗb���1��g`�ӥ�os4�Otp�\껍]ikvҢ0�N���6�s6D�l���X�p]�����7�f�]�c|�|��X��ߏ9��S�@��bdȇpv؇i4�ҭ�/JF�9�T8V���4ف#�*�t��f���]���=`K�!)�ww�6DU���_Z�q��_S��;ւ���l���j����}��Xi+�'���T�۵����W���qͿ�zj�V����E�"�D����Z�^k�ґd����y�d��y��4�ĲbD;<����t����37;���{�v����Z#.��߹u
ԇe�ʝ�J'�;��z0A�/��*;�c���*N������_j5�5��Q��Dr�W��T�����Ȋ�Wl�(���mt�3/�x��F�4���Q��m]�bP���Ϧ�׽� �	e�4�Xȩ|e.um���Ʋ���@���{IĦ��%��A����Hb>(C��.<�c�o��|��佨x$<�=鰰�c�Wq�����U3��D���Ӧ%�쥧B�|~!.�I�Ɛ���5C���Rż��y��o1R�t�;i�,^e@&a�{\bp�P�}k��GaW�d�ƶ5�M0У��Cć7g��]��+8ow�2�f́��ck���>��nE�N�9�3�}l`����u��w*=O�zm,�p�9�;y���$a�����7�D���w!R�XT�Z���1q��d���v�}H�4����C��m�V��Y��n.dM̦��GrՀ���-{�4�C�WI2 ���n�ղ�H��u5�{#3�DT���
ͱ�M�C���v,m��/�{ �(�u.�EˍgH8R�SET�>�W��[.h��v��:15H	�'>g��H�E�phڍ]��[TV�{AG��_v�I�b�ɦ���0o�ȭ�>��;r�����6�>��Z�/���.M���K�.���@R��{�H8��1f�PW����WLg�WF`kU��������	ߓ9�L"�W)%���WZ�����F��#�Y����h��vN�+.��ńrv�4��a��k�\/E����	,8�����!,2:wK�-n$[5>w���V�j!����ς�k֖
�I9��]�m�՘�wv�-�{�v��z��"�+7���}d)�va�X�9ـPT�d�W�[gI���n`#ӈ*�ME=�;K�~a`En�%�t�L�I��$w�\�;�(�>���-��4t�(?��פf>AM����"�c��^���0xζ�OH������ݮ4`��-�p���ء�B��\�qh�!S70v�k�@h6��,��;���;���N�0+y�����p�ZCmg@��a�U�q=��ذ��3�_^dw���2L�vny#�u��A��e��]
컘qV=|�[�ZG�CSE�T�������\��<4A�.��Ɍ��˙���%�]�vl�"��R3u\���v�v]�<T;��ͫ6�`'(�.s�= ⭷��sƹ��qn#�d�93��$kw,���u!�K�ul$�gl�kRTsa�V,�y�q��6�/�n��Dn4;�2	����/��b�]'C��}�W����N�E�� �N[f�3� �����}�#���Z�1�'=�#m�U�w�WD�M~�������-N��	ao)��#�V�hl��E�yk��6�T�G�@om�2Q�p��]2��|���5z6Y�����#3�����n'���M�1�^��S�2Ch�"C:p4�7�����Q߭8��{�,��&��Ɵw$��S��J����^�D輛X�Y;(u{�N:���L</A��U�b�ێ}��ۈm*ܼ���G�^�&+�+��V"���{w�(�g�μ�+}�M�����#u�:����0X�0�2���%\:��aiP�QYʿ;��A�qy�m��Z�y��v��m=`�}���'�;� �]�5��F�xR8���|���ڠ�hR�Q���2U�������ٙ���df/���P5����r�I��:U���bx�E�i�Sp�����s�VD�OR��#�3�AR\ye�s�ٛ�K�[4�9���PȄ�V�QSf��7��kC�*�ͭ���4L��P�ԋGa��YV�FxV��`�$w&��TA�ˬ�FV�;���Z��N<��c��zt�P8��UJ)c;o�ow�I�s)}���uhཅ�|y��C���Ǌ�5�p*�U���㦄.���iѸ��U�m��Kz���a�;����G9���:d�,�u]惱��&��J�(�	�{\f�����ug"���5!���S���;e�T��͜6p�\0�¶��v,z�檭�$[J���+���ԍb�ԼfXW���F�t�;�ʛn�l��Ɋ<U� ����m��	<�`��>Y�IAW(����͎���:��-���^g7�%ca�|sA!�k R�!eC� ���u.��GY�}%f�*{y�S��&�v�6�Ms[�n�t����k: &E�>`��9�|�Ѿ��;(>��>5�R���Qn&Jo2�C�j��1]G�&�=���ƟQ̝(��S�v�߫��7�a��2u(��3U	�x�@%��-�W*+x�;��Y�5��M5%�\�K�[*^��peM��(Ծsdko,t��H+v�ޜ��ϗ,�q"���5@(u��\熛!��
�s����>P��ӣ8�s����y�����R�V4�a��.�K(��B
bu-o��{2��mT8_J�,�Lnu}�U�4V�
�b��_bL+��/7[�O���|Ո�٭�1d�Xo*�]������^
焫���1C�f�X��m�����C��,��VÕ��<�B�\Zt,C ��b��`��6�H'.��`вC��ʈǈ)R[sX�v:��,��
�5ā���9�
\��v,.��A�V��$�b�Ǚ���]�,L���	��+�͡l�u�F:�;nVM��W����w�b�t!����`��A�`�;���*��y8q��M�<%]�Y�����#ѣz�u�<Ϣ��ϛ��e�4�F��#9qպ#��� ��Q�`%��5m�i�z�A�OfbC���pI-ZY�ܭ=y�t�����bg����k�{�ҫ;e��f���Hb��EaS�WF�Ҟ-��S2�J��86�R�(�YQz��ܹ���ݖ+q@
�k�.**��X��\���3 �اM�`(��p��ON4eF�r
��^�o�
�vY�B�d�)R	��܄����uڸծ��!7���jj��L_�b	`�4e(\\����]�{�ۻ�0F)��)逿��zo�d��ʚ��M�5��8 �o`�u���m�{�Bܲvۀ$y����{��3toA���)M��	�&��mU��NW:�/t��#Z������i"�Y�C�EVk�moآfU�t�-�	g*��;�E���w��
�����*l����ܛI��_wf[�	�>����sp��ǻ�z����W��(�>4F��{�v�5�:�� 냆���D}��D�]�2��E"k-�����.p!�Ԁa��V�1*�܆ڢ�F;���p/���,j�5y��Ì{�c�zmf3�z�rwz�&3�,�3�Ǿi�/���x7&��"&ڪ"[}� ���ۂ�vz���FN�B����̌�쫁OHݫ�<���5�3��� ��|�����Q���wڄ�`�@�Y]�j���9��1���
29�<��lQ�x�#;3p�`��v�����9�k
G�^���z�R@�hGL��ݺ��}�}4�{�Yɧu�e�n\�� ��-�`Vn*8%v��/�{�R͑��KzP��)C�u�h%@�K��5�9y�U�V��z�s���5i�.�{��tQ�8{�*����ǯ&�D�g7�x���+8�Ü(�MLj���%�g�c`T��̳�+#Bq��)>�ك��ݹ]��חL�9�i��+(^���p��͡�o^V[��[Z:��+��H(qUp�Y��VW\ӣZr3�2�	]�y_V5�x٢���O�+�c��9��l�X8��^l�Fc��2�o��(%��DH����ݚq�K��δL��h�u�JY1��S�8�rZ�Z2��ƅBP���
��H�^�ğ��<���px*�ײ>�6��"�L�<l;����lP���g���4	��X&ʥ3�kLGG �Ғ _ V,��>o�+�S��IΣ�9�i���/ir���M٘�:�U-�9.=��gŻ���;�k2e��ޮ\8����C*�I����xN��c�E�g�v���3�b���`ו����=ܖW8ݒ3��,��k�_ω�&N��C��1/@��'�3[&�A��r�18k�R�ҹ���NOΉ�e=��F�YԬ�%�T�Sy�_��m7��t|.rI�Xk����7�lF��C��Í8��*(�$xf#��G��f˴���(({�-���Λ_&?4w�=ި�hl�E��J��M��q�_a3����ʊ�a�I��h0����p��W�1�]���wΆ��k����"J���]�TypΠV��]tP�:q��yG
�8Eb'v*lz�ZY�M�P���0,��[��7mũ"q�޲�'�����X���@���V��N�b�8]X��0�4�R�iv&p"�lE�U���n�{`k��{80�˥�Dtn�%P��OGJT�%�Z�PWXÑ�q��)f\)$�h��+� Z0����C��F�X]fs%��k4_\9FVٜ���LG,S��;�� ���Yݾ2�:�>����J���d#s<�����U���s�jH<��x�J��
}r`�Q�/ZN�"�������݊�8��}������s�j5�E���o�|6�ޕ��Σ�, K��+�o�e`��u��03�,bx���r���3�󾝁��v�ި���l�a����+��z8�_�ǝ���+�.hk�r����x��W>ZnP6��� ӨV%�!kr饸N�nZG,B�n�.���jΏ�e�T���f����c�g]����V	.�������������핚�TT�8W:�6�.b=@��v���9�m��\6๵�PG��/;I=�
�}moT*�|X.n����m���s����T��?7ʶ*�j���1����#�/&_S=���{�����v��7`�viv7��_{rS��@��w��N��'�x< �^�{�8�PYM�	����jCv� �:�����&Z{���Fl�Ӵ���výM��m��@T���r��Xn��rx��[�(��/"�u5�hjz}�����q�V�g�R*���7H��\^հ*]�TOng�:����װ�"K��䱢�z�.U�Js*�b��]�\���ƺ85�"v���ѧ;ȟ0��N��T�CǇ�D{��Q7;_�}�lө7:E�CƗ�w�z{�dqNO^�]י�t�܁ɦi��w9�縀�l�v���$z_LUx�ޖ&��������A�E���9.D ����)��:vj���oϦݰ���
ݳ��P#�Q.㭎�U��]\!�kG`[.�>�֠�w�VVË��Lz7��oc��\��X���Ӓ�k�*�]n$�����R���iC�	GlnsV{���*��oH5��5p۷�7Uzf�g8ps�a�E[�W�=U�6��n���o ���El$�p��RM�<����&�R^�ZZ}��t{"ӽ�����E�c�r�Q;v�WJ�q���6�-�"M�t0����Ě�P&�@���漵�1#xoE�|�|5��1Ĝ���\���_g�3��y��Ge��t͞�h�c"0�[��V���������}l��#HEwv72��DÉ9��U���Mj<�Q���@f��R�ۙ�$�e��}�:�
�޹|�s��}t�0]kA�����hy�l���ٳc�T�G�%�d��grc=X��,�a��c���|�=X]L�%�Z� ��v��Zx7�R�9�K �()���	X��iL֩������72t�����%���h�k^8��ఱ��K���m�+Q��!�c.�1޳�WQ廭������U�ڠo;G[�S{i��X�P�h�nCF�ɭ�}[2�㶔!�@z����ݒ�E�H[����vK#���cz*|��7Xs����LHNk*!՗M�������s�l���#t�p:͵{,��c�Y��sf�k|)U��x0��@(��� �Ms����<��J�s�MO��Y $Vf�*�]%��g��\� Ǭ�ُ�[Ah�=q5�v��X@N��u�۠�v����~[>OQ�!��a�tzFcw�yj�S�������@ܾS��/w�ܢi�`�wk*a��Z�6q�8����a-Y�&�"�hq�[X��[�qP��T̲��V5ѺV�WZ��6%��>�N�����k���b�y��E;$D�7VV�j��� ;��xIbQ�N�vm�l��6�ٺ��O,�Wq��*=��-%��t��ĩ�MG�[�Z�=�1w�h��U��p� n��(pE�u��Sb�7c0`�Nא٘�n��#x*Wj.*d��à���Y����|>������b�w����X.������}�mh��L$shz����a��ǔ��X彎�1�|3�%=���J\�b3o�Χ5u��oD7�4��XJ���4�@b�ۗ˕�����,��8f�VT`�&�U:D�*�s�X��؎��4�޺V�o�x�6��Ҡ�T����MQ��CJ��g_jwq��n���ač��|eq�B�97�畔�BZJ37��DH5��~rOP��F7;Z�]K�+���j�q�.#7rP����VZ��]0q��x�8�{�V�ޡ�6���#�:��_M�[56\7/�4���;v�z�^�Cpթ��-�&jxy���x�V����ز�}nG˹R���W&\��pך��[ѕ��*A��t���2�J�w;�t2�gnu1+��Klm��i퐬��$����ǓL�5�h��X��w\n�tv��Ou�� � dYC���8/3y't�-� д�]/����n,S��K�f	���J�%����:��0M&�7x(qNE�yX��s����ҩ�͘�s"-�}�Stw�٘��bq�L���'�}���57'(K��ck��#*�^ߤ^��|7�B�OT��^������t���+w\㧈���w7���탷`zr,�0��E�:^8�9�U>��u��k�����~����h���
"�X�(�h�)(*�:�	CQ̸�k��(
���i����@bmdh")��TP��5�5̀����&��5��&i�Z��Z��Z���f�h��iY��]#��e1'TW#K\����֚��m��-P4��.p�:qL\�M5Z4Rit5LU��h������K�iZ!�(�ƨ4UMͮ2*�gXu�b��K��4:(�	l�Jk�6T\��4�����-.ڍj-�ւcO.\���l"����I�)��aѧ��v����z����`\�u��)�no`�H�{�c;k����=+��;L�>g-F�����7��A��]Qk)�|�Nժp��ﻶ�<�|��?୉��uƍ-�n�Ij�C;]�Ƌ�|�PF��y�*ڥ���l� ���)�T�Pd1�(��[�[#���^��eV����wq�c�k��>�ܨ�s%�@$n���S�Ѐ���vc��������Q_���
Sg��ؾ���!�Խ��EK�S�ͬ�_�t�t�z��e�+�>���^�o�����Fl�t�g��o����f���Wlt���<|&�z�ŅX�Q�u$1�+����E��>��D��,X�8k��P��<���hW���P�h�-��'<wV)��y\��y=�|��6+�y�3����4<)��@TF���N�F
�Zbwg�\�GP�X48K�}O2�:\����E��w���v,�*eF�oK��P�89�����q­�5o���'��˫�������o]��Q�l��4�f�K$�~+��e«4��r�\���[�U��z��g:v{�]�
ȓU5�@��g�bt�:���~���=��%��N�#�ܦ_l�w#O�9`���4h��`�L���s�(�Y�
=y�U�I�%V�ɪ�`�ˠ���'K<�d�4�.�⾎}�跉z�{N����3u�t�ma�=���Ğ+���������Mvs{8�Rp>���_�_l�8.��n_�R�?i��U��K�ysx�����Z��s%g���t�c��@��y=���7暿����2[���GN3R��1�b�]N]�C�u_#[�r��{y����T*�i�)�8b�{C�PB"}�3+����	�f�t��7,e��9X-�Eh]�{��������U���5Z���X�׹z�zA��S�W���]H�J�2����Wǯ���*�w�b��O(�~��y�D����uY{Z����T|ڰ*���iȣ�N��uF����@S��FA��z��WvS�4L:J����y}�1r�=>����f�QV��(�e�qٕ|/]ۢ�c�s=&�&�p�bb0�뺮J�0ڑ&7�z��w�nW��e{�7��������E����a�y0�ֹ�f�� ;Kq4�f8ạ"nż���f[[�ā�{�/~�m��c����o�d`�ٽ� �J@���C%��epe��fV�eʹKz����(�ϝ@|��2�w�#�E�������[��.Ň�o玹��s�q!:^�ȶ�*��2n�`��/6Gw(.t�/��2r���\����HX�h+]�t[E�,m\7�vݎ���MH�
���[���q)i2we�0�G�4�.��I�3y��@�����;�8k��V�\���U�tSR��n
V�U��.Q^y�f�.\c3P�3�S���^�U�xcG;�7���A�����*�H��pn��*�'tԚ���M0���sx���t�\tAx{ӟٞƴ�+����08(t�$�7����|��!a������!P��/�:Q�҄N�������C���^]����k>���;^H�*�&{t�59�
�sY(s�ŋD�1Cr��J����BV%��s����Fș�z�+��B���ؔ��̪Q��	�{p�)��X)���wP��t]r̹�qJIiU�ou龹뺧�&�D|�q�w�O��w���eA�]�'� �9엃,����V<�t/�ꠅxd�����S"~*_�vȡ�� L*�������T�,$�]NOC1�8SuG
u$	n� 7υ}�n�bQ�V�)ｯ.O ����J��VN��~�*�n�a_zJNr~D	Z��;CD�f٪�E�
˗�����;���H���t�Ҙ�.|=qc�hߵ-���
����j�e��_
y$�_:�SN���7)�*��K����)mh�k��7:��+�f��e5,�g
;�s�;�h_n��e]܋��j�J���은���E��#(:ϛ��ιt%O�L��;���-��8Y&�fW�\9��"�M�Y�g��x����`��c�u���#ʩ�e��/+;�mVGu�Sv+�&�ؓ�,r�o�D�������ŕ�9#��K��7\T:2�����P��V	����߿^t�fR5�ߔuQ[�0���<c��n]�����e���*?pE���uJ9�߫R?g�,�~�&�?��h�_+|.}i��]}��6���(vx]k�;Ml><]V���.�~g;��~�*��{�uZ��wE��pZ�w�r��g@	��\t^L��@�mH{�H֕>1�;�q����9��0Ί�fvй��H��N���%^��g�į���]�bC��.���n�Y��76Ŷ*X���|�M}����h��>Q7�����U�H�/��޷�}e�Qa`��VS��e#�=��%Þ���z�����2+%W��}*�>�[6�U)�o.��Hv���~�}&�I��՘��E%LM㒵_3�MÃ���<��t[B��.�����ջ�g7e�(TYw���'s݃�x���S���C3�tdY���==��(.k$��o2ꢜ��.���'v�YnTj���tbl��A|��z�_U嵱�w��7��qaq�G9N��rQX�C�@-Ȫ�����P�q�U[��m�O"�Äx:�:04�$a4&r#O�)�!l3t䡑D�n�A׃����{U��w]n��[NȬ8za��u�|�
������,��˸����c�M�5��'Oh�0������Tɉ�:%q��2��]r���B*���n�P�e7L�;�Պ���{�7��A�P\58����m���մoL1�ba��i�o���K�p�}�3���>c$�"Ɗ co,
���>(xnJ+��[#�O<E��>fi�*y6���Jeӵ�0[��������h��Q.�X� JwNJ��7��׫�)y���gr�+0�J�<n'Z��I��.������W�z*t�7U�ù4tp�:�e�Į9./gh��f�Z:��J���^ѡ�Vs咨��%k�w����ˎV�I�;b:��s���<gkp5���q�����06����LR Ws�`cU��e�#)?< {"�W���܃��L����ew8v��^���e��#J�����T&�[�ّS�qە��8��Mz�n����Z1���7��{��d����\�ܷ�:o�]��:�`�V�|=o��7|�	�c��F�hq��=b�c]�%��g{�ݿ8�}��]��o�T6+���k���s��8�P�"y�L�4,�U�����#
��C�F�Z��ѧ�Bj��W��P�0���=�
����Iy�ݸ�x��7��s!�j>[yu��7ӷ�k�yA���p3ҺZ\~��}=���SFl⧼�³�v���|<Ͳ�\q�Tp���1��9β�Q�J����?L�z�G������4�W.����Wʾ�+�D3�m�|nU�����#o�QJ�X��i9��;9�aZ��)��hb��*�P��s�������w���CJ��$Q	Skn_�x��M�m)s�sq�G�|~L�ĸ/誑¢y�ÐLpweB�І���qoe4��i[�R�R��UF���RL�����(h��9T��]Sv��ҏn�*鞌N�V.���Q�Y綁[ր!�#u.H�R`@al��9�ms��}0�-����嗙�'�	�C�E��Y@u��X�� '���/�B*-����݌�u3] {�r�j�<��a��p')�`����v�fd��$�E!�ws;ET
ݺ���63"�M�X墸�r-B�Y��Ѥ���10�������D��r��K����xx.����3V:L�oR |ٛܳK��l+�2�w	6�6��ʣ2Aɍ������t��:�C��J���n~|N���;�+��pjc�|�)�,Q���c:�ɘI¨���'�fDwU�B�R4b�h�H#��g�T��}(�f��̗�����X~����՜?J���R�dܺ�F�������<&�+y�Y֔:�hC��k摙FjW�%,u�e_���@���1�P�se\K�K�/�fju��u�9���𖕚�!�U���p�r�]/����
���-�q����L]�����s���5J_h��D׾�/�k�[#0�/+%#�8���}$=ZT�h�X%����.j���˺�C�;N�2�����?O��ߺ¡�~�ŪĶ�S�6/ ����lދ�]��O��/L��ε�a낳�,w���Zp����[/�$	E]�x�4{�58��SY�S�pȗ��K'�2���nX�]]�Olv��j5vY�6y� �|i�u�0ˣ��n/�Ku�����/�*�[��7�h�:wf'\>Z��=g�b��6;.9t�=ב>�5�����U7�=�^��ޥ՚�e�=���/pmf��IZ���ǉ���:g3@~s�k	��g�0.,u!o�����S�=Qb�Ww�qt�~K*�.��-�MKt�}[��lő�K���JsR�����������i�R�@@}��;O)Ok�}�{�lwg��y��W��d�� �ݩuB;�@Ud^��=�!` $x��v�*dI/LsKus�*vr�vn�������=gnT�4GnFor�U��&��"���mڵ��-CO3n�Dm*��z�P�;�z�Ka\Y.�,!�x�9�l�.�k��;�ٺӺ�M�h�=�9?#���= �L��TG��+�MÒ����I�:crmb)AvsZo@��
́u5��W�s;�P+��_�o=|+���������^oc������������_���&ƀ9�.�]�ʩ�����䭠�Z�_8�á�Vz����VL^gfN�wn���)���6m�L!�>�Xn$�^�<�+x����9<�f�n�-a�� gxD���/���|'n}�{��&,C���"r���н���VC��cmgz��S�r����3T���*��T�TP�\�z�D��껠Df�+/Ƀ��>#�d���u�%[��N���(�͙s)�R�q����Z��G�v�}!�����S��L�w���^Iɹv�8�/O�����*������b�/����}|x���J�.,Ұw���A�|`�p3t�,~�v��|�DU�Nr���h{%U� ��/�1C�����4#ƅ(.����g���l�yJՉ]6̯��7	M�¢�q��,B��e���ӟku
��3T�]�z�n��Q�O����?!+���m�]���Aŕ�~u����+������tOl��E��=��:4r˅ʥ���=����)�u\�e���0�Ǟ����m�j�w!�$�԰Ǫy�q���m]z��P��4�Ϊ� Bz�[�UH��i囡�/�^e��1�q]U����ch��T$�#<b��TBr�;.J�5y�U��z�wUju��XOm�t�J����Y�`��/��=��?e��gG�7�;������/�DŶbS"�T�O�t;7�1� ��#z��Y�b(.,D���v�,���̉�Y�1qۉ�<'��O�ׅ�
�R�7��{;6�a��;[��3[�\(G_ŋ uD7�����,�9S̎s�a�>�[��޿��������0b	��f`ڕ�j���F��ۙVm��4֙%�'�������)t86M�B�mYJ鶹d�O(�͑S�e�<�d�����r���/Vޕ��-ho6�7Lמ[��m۲�b���'��5r�C�3�ٷSa��z�E�0���q��d��g�������0k��aÍH�\���j�=���p,E�U����	dKy�;_BAf�**�a��fj4�U	]�Z�1P�EN���<(� �_K��&0wp��2N����RФ&aa�6�Ζ�e*�7��А"�٥�9G>q�퍰��ǔ1MշEI�U{jw�_�T��͹^����P�4���c���Up���UwBy!|����,̻_��v'��h�ȗ�&`�s�!� _�#j�� ;�9B��§���S��[5���Wכ_%rQ͗Z4���Pʌ��hųQT�+y�(5/U4�f�CNؼ0û�_v�NP�p�EpZ@�8���U7 S=+�WvϬ	گ�Mǯt�!�^)�� ���r�C�h�[1��@G���ʔ#V���͆�n��[�_u(���P�a��?Co'���xHp��>4��wI�s��׻2���IY�����m�U0��̪�B:����˯堽9�X�}_8�u%��d�x�F(���P(C.��:�{u>�{�ǽ�Cȅ|qѝP��hy(�dϽee>YzѪ����ѐ�D�R�i�#��q�;4So�>�8>�z���˽��&���]Y��:e��`��NZ:�%o�v�)c`i�Q�݌��]���s'���| 끼7�_cu� h-}8$Aac���칊
R;͝+��CN���7Ӛ����N �eI�5%�矲cĔ��w��ޘpJt���S�73�;D�7y5�4U��Y�ü��-��3㊐���s��Y��]k�z���۾z/:��	ZV����������Ϟ���/�ԍ�[,ӛ���'F��Uv<���� 9��黵9�W��,.�P�]�
\�T�[*h�]���m|{3���Bgݵ7��I�����j�M�s!����vH9wgn��[����zZR=�O��6��bC/����u��][~�L�M����6�o
+�Mr/�j�<-L8$/y� �o6,�A^
޻�Hӧ�.� ky���즊	���f�B�[ٙ�M�|t��-&���d��=��ӝ�;�2�ݫ�Ԩ0郷yur�oe�T�Y&ҷY!v�6�ջ(^k�^i[@�K�]��[�9X�Y]'ne1Ȣ�Uq��}6cۖ;kD�'��3�;���F����|�XsD%�5؏Pֱ����ہ!D�$b7>���S�]w�v �Xm��tK5&�8�� .1��r�n�@��;�����lc��2�É}ۯ�u�M��3$�?z�.�\%f5Mh˼��a�ۦ�"M�ڳ�be��H�T����=R�<o0w
�,�R�]t�b�A0���/��u0��x���J*^�HĻ$K���PFԕ���P#=��-��)g��cw��-A�m*�7vI�gw�X�#.�x�%v<+��+�n�~7���PĄ�]S��5SU�
��ʅ^}�g�f�`�O�l��E�-�(�VA�S��j�U!�6����`�zk������>�u�k4Iռ���H_`���av���2M�k�R��xJWð���YP��=@�rU�¯s��
�Gu�';
�{Aո�,}3
��T�ͬ��u�n�&���f��w��̷g⻺�Qm��&Kn�cS����Jvo��]ᇰ�I�����i4M��m��e!�;�$��B^�!O(_\*mrc9!۶�G=&l\ދ�8D��c�\0�e�ϩg\�����O=��E�3u�g.��N
�p��L�B��B�=�������W3]>컢k�c��K�f+��+<�P/j��t�	��,��.�Ѯyp�6_XA�k����]Z��<v�c�^}Y�Lh�m$�u�op-]Kr�]�7�%��,T���w��f7X�eV����u�q��;=��B0�dy�C���J�ܞ�B����9��x�&��e�m��W�v�N'c�~�3D^�E������)cU0%�P׊�<)m)��8'ir��|��?"�)P�l�[4���te�*%A���Ҏ�ۮAw�y�mg��������AW_�rT��j4��4huE%h%D�����*X�I�b��np�Pr�O6��d((B�����)����STQ�h*��4��ъ*��b�N�T��xN� )MFƊ�X���l:�j%�0EMSE1�h�).gAT��i�X�4%���:�9<�X���[:4�j�ti5N���DTPrB�jѪC���!h��:�5���Er9��C����A����b��HB�䁣F�I�t�9h9 QA�'.\���!֨�ZM6��C\���N1�B���#�\%7�V�h�׌��f_S3*J�JIq_L����� Iʑ�r��Ҿ����'J�͚t=��I|�ĳqNVl�Jh��1@1�X��믾�U6X���y�_ +A�>GӼw�i-r?O�u@h>�a�A�M���p;����ߛ������Ǆ}a�c�D_V߇��99��]��޳�>���b#DH>�9����?��z�OR��O}�����#�7�'Q�u@u�T�}��|�����N��4�s~���Og�9�0r|���d��u	T>ο{������~��z�����b!���}�1b �bK�9�?��~����}�w	O���Ͽ�:�z�I�󮓗�d9�|�Ph=�^Ho��K�K�t}�T�1!����H���9s�՘��Ni{�5
����ur��9s!�������`��;=���`���:���r������t�����t=�R���=T���y��^G�y�:�/��A�|��H��K����s�)�_vh�/ە!t|�����?A��l���u��g�c���'��;�/��%|�޺B!��<��y���Zc���A��!��ߝw>�pr<� ����qx�E�)�E�"���X�p��������w����u/"����h?�윇�5콼����7R��w��t�&��BS��8�F�T='���wR�'P�Ǧ��2�5�#+�}C�c�|D�����8�GRy?��=��A����9	T?���w��J�����)��^A����?`�˨;�4%'�nu����4|>�ǹ;��C� �B/;d���G��/��V} DX��r�_O�;��З�w���)���\��_$����4��C�>}��%>C�r�d��*�����4?>`����>�A�>��?F�NFl%T��Uiћ����0�}B>�"'��?�����u�{���u�����@F��{�}����I�̜�/ە/\��P�5�_���_�C�<�_������|����?�u�^��^��d{�0�v8&����}C�|�א�����A�F�������#�Ͼ�J��&������J���'*~å���?��9���y�׽	���G%������}<R~�?It��l���=XWA�C�l������o�ͬ��YfV�┚eŎe&���/�4Sk6L�+��;-���fݲ�*]��լ��{t�Ϝ�8�X(�C��\i�X���".�+����N\�^s~x�����<s������A�.{|���������盩A���:����%}�e�iuO��/!+�>~����'�k����py��������O�?O �ߜ�)~��x�#����=�^L�1H�Gޜf=�+��wngMv������u��a�8�������~~���r�>��>}�rW���K�/~y������󼧒}�s��b>���v�M$$�>���G����-C�a�85�_���GǼ��4�z�?oa�%�̞�Py����:��5�=���w��y�o���i�.�?��<���~}�������uR��6�;��D1p�#�z���|D�u�?��{��)�~}�GR�:���BD?o���P��h�X���F��ܟ���/�s� BA�"(G�������.��|�����]~��S�'��8�����}������a������`��?u��pNA�m�N��˨��\:�%ѥ�ẇ!+��9���9'�5�;����'��=��>{�����c�ه�ji��>�@H�C�و�� ���'�G�r_����
^Cϟ��C�����	Oq�:���s�Ri5�_9�A�!����c�>���֬�m�_�g�Z�|�^���g��C�������!�<�ː~����;���><�ې����y�����G��9i~G ������Q�����>]C�K��-4"���n{�Q�3� �;�J�*��!�|����N���<����E/���u�4}����l�?�ײu��c��CO��{�;��������e�̼�A�� (��u翺~BWP�>�	��^�Q��4}�#�P��A�_��u��� �~�I�JO���z� �%�w� �'u=C���GP{�����:���\��{����<���{!���!�t�߮������J�.���ޚ��؞�@P�� ���w�	BW�������&�<�P{��c�[�;���>��X>á(�Og�|��䟏�9y&��������<�����>Z^�)�?w����}�=,���qn..�rйQ�VPw���\��b�ɮc4V�g�IQ`*�rԌ����U�=j/
�³7���W󷙗�	�!8+T��0؆��`��m�Kw�`��+��kں|����~��U������ri5���9P�>A�r����t�|�͗�������/��9���4���|?�}���%>_�}���4���� ��D}"#J�]�5�D�_{�?|뮽���G���������{������������?aݞ���p�A�c�y��h���~���K���Nïxw	G��\�
 �c���4}DC3�{�^����������w�k���RZ|�}���z��r�"?p��~BW��y��������:C۹�|�������A׾��;�A�@|=�îd� U`���~UTU¾#o>WX�[D{�w_q��Q�}b>�"�"%>����>n�����!����e�`>��A��O���u��	Tg����O��u'�5����>��rN߾�t������� �:���������3� ���7�y5�#�>"!�#���Ӱ�)�}�:�@{���Gw�����`�N��O��$�k�>�pwP�=����wy!�K���8����� }{򯘯�U?|��?&��(�S�雟_�
�>��>�"!���Ղ>�=�BQ�����\��4�ܜ�{�����	y���}����Oo�u'S�{$��9/��|�����������v{/���/'�}�O��=#&���wi��O��!���h����Q�^�s�����]���K��솃�����/~c�~u�4��y�����%Rz��{=�W�>s-�� ;>uém?��9�=��������xO�>hR줣3="#D} ��ǲr?A�C�=����d�O�?���pƃ�:�u��G�~BP|��ރGu!C���Ηw���y�;��t�<�]G�xO��4w'*�~�������>����1�1"�ѣ�����A~���w��>O��	O����������G*gA�>���=�N�&����罯�#C������^@v|��S��~��g�q=��4����������H�Xl��s�tz>��|DC�;�Hi��|�B^d�NU���A����u�!��{���!�<�B_��ӡ�� ���� �_����y��W������I�#|�������)��N�A�9��%Y��e���U���^��ĕ�iL���6(Ӝ:���w�B{&^��Lk)k��wC-vz�v��u�a�;)�O��5�ڔ�a]m;�ţv����7���;A���*����*���z�M�vNe�&�,�6�%ý��}��#�x�^K����C���X�����?�����u��~_�=BB8}�՟ ��X~��sFz��S2n�v̱ٙ*uJ }[B���ٯ�	]>���|Oi��?�fgq�RlZ���VZ�����Ѿ�Նz�f���p�U�#�^$au<'��`�.�L!4d�]ܤ�k�����TF$�؂a��R�_���T�@'��+�y�S�c�g$.[�dO_.��yzwT�"��0��/�� �ȗ8"�
��WNOP�b0lcp�.Q��Ҝ��?J?DgR�3;����WTj��C��7U�n�$s0B�X��Y�j�-�!��G[�ٹt�d�8�������M<t�I���~�jS�-��	�o���{x�蟴F��*����	�XX�Pt &:i+��#X�@U��Qz1��Z��Q9�w�S͗|lD=�;�{�G���_]�:�`����SV�'H��w���u�Y`1�o��7|"���	�M|��Ӆ�%h�[T�����FA��b���*�oǕ����,��u�VuS��It�s���)g7�.]k�w����є�&����l~���擐�����m���A�\w�� �
zŝ�R��HM�����(N�.�.��s2P�z��a��#T��ի*V�St��e5.�9�0�㟯�g��h��!�pX=qU�=�NÊ���r�jB�v�F?��?TY��oT�W ���r�]z"#�3�y	0T��j�����Lo�&�֬��t.r��[u�xηJ�v��P�L�|K=�C/MJJ�S��es�3�䶤��![ﳩ�0���M�U��`�����o�_Y����Q�m>��u���Sy܏P S�U�B�
����D��>���JT���d���:����F�m�)����g#�j�PB�k�4\	G7L�,%��G4s�㕖�r���{=px˵f��]�qU��T�'��5�s	��p؆�O.�
�("D�A�.2��.����Sy��k�j\S�y�ӄ�4�W���b˜E�ȗ�[ydT[��D .;Z!8��]pp5���\gm��F�!��0�?V7Z7>������#�����
�a��H�֑Uj-پ�6e�Y{wf�R�!�,
�Zo!���,ewU�B�+��c�r���;@��M�V!���!�x����<��-�ou�s��ٗ��ʉ�f�J�mn�^{���뮳����K��)��z��]�-�M9���Q |sb)�T��)QS@�]��h�a[e�)�N4%��LGo���t�� ȍN����ڇ4�Y��� �>\��Ȭ�`�J�V"��v��!ԣ��T��M����^ew;	E��%��t��$1�z�`G���Ɯ���Y��:��4;��#)s=/�#�Ϡ�3������s���@s�Bx�9�CdГ� l&+u�-w��`��t�k%�Ul舾/���2��vab�����=��{Ch�^�� �UmX��[�I�<�n����r�	�8!ξ�D�#�F�b����b�Req�3Jw������*h(���<���?f��p��ʦ3HB��l��$��\wSg�����	�h�s�zm�6�mU[��㕳��~�G��5�yJn ����-*�Qs(sȍ��%��7�� Br���}����m�{sË���@8��t))K�Wd�|�]�S�x��������m�&V�b�_n�]y�� rwaۦ;\��D[��C"I���M������H�:��K�S��	.t�f$A���z�Ds��s�����a�����Z�ɂa�6`�;*`}�T�9�ӡS�n��J}��v����u:��%3�==r<���-�{QI�^�=)ͯ�yܴ�s�,�ǈ���}��M�vɥ�c��쫯q�x\2���au�[�Ǚ�)e�J�ˮ�K6h4�B:�,��^�O��D��8�}-w����
5t���i�k��=�N�3��+��ے�w�w��&�JHB�\U"f��/⧲Ǩ9e�Ψ�c�!U�w��>5�+��NY<+��:?]�"G����i�FvǸgə[��u�ġ*LO�q���d�����T�*`�^�r
��*g��g��ɷ���m��d)+��"�=,h�
L �᳏^�x6����P�MP�
��
 d4�F��;���7��=��=��B�mä���Z��j���6!L�hf�!T���~7��Q�ܧ��lJ�i��VL(�L�}E�!{Hk����i���}��{'�@k9�꣄���~���rq����P�ڵ,dZ�5�Z=st�^��<Ub�(ka�uZ����;W�B�k���Ӽ�c8��鞌[�8
�j�g��
�5��D��_�0���{8 �G�4ejW��ӘpB��7Ӱ�{�F\S��#c�y�p��]���q+��s�Hp������,��sBB®�������cKQxi�ڴ��g	�R��wB�0��Y��s7�rK�/3�����Io���[U���������#��%������F`���ڊ5�u])�U[ջ}Ќ,Nk^N��p:��W���y��>O���h�����C��u�/���u��a����m�k��j;>O�?<�pH�v�Y���.J�l�
k�j�i�3󁨼7�f;"�1��Vu��`V�c��v-��NvMSB˾K�^ւ�b�'i޶��jK�{��e���6ܱ�[��4�gڨ��u����[��*��h��1p�T���\E��\F:����;H�D8�zo쿕HȒܩ��Z�-�_w�yh����o�_Qr�-���k���Zȕ�:�/~��u�	}�vM4EC1��V�kj��֔@�He�~
������zK� ht@Zb�(:�����*�	�Ά^�m)����T�$���z���3�	��y���#f�)+rJC����VmE7�2+�hn�;S�;=-oi�7�B�P�XӢ�����ӛ�J�,�xW�d�/Q\�=�����Wc�F�"`��h	�*�����U�N��M�#u8r��T'w(t+]eO��h�Wʾ��3��2v4������1_6��KS8|Q'�
�F:O�]W:H놎]W�l�2l?k������NO.�buj�`r į�pkV��R}�/�~��С��:9�x�"N2ۦ8(9��-H�ث6F�����ܥ���]b<6!�(s�t%����3}��0��姠B�,�V�fG9�(GԱ{ƥZ2�80*��F���e 7i�0��DW�u:钦v�P-��T��J1�p5�}�̂���@_��ŵ״G��6��\e�uJ���Q�k��{���p�^�7��or��M�`���8�'k��^Lu[��p4R$��y��� #@�c=Z�DJ��Fn	��mi��,uFxs���;��w�l�rU.�P'��,/�L�!��N�7�a�܈u�i���h�[�Q�*p`<�pG;�H��{K�L�����&t�QeF��4�,<7�W�pP;�)�K���*a�X�?��g��R�|(Ę爺���ih����:)��g��r���e,ݺ�}��J"����Z+�O�Ϗk��n �j�\y�]HE3��˯��˶��7o;:�9#:���jݼ�2_X���|���wo ~B�������ςTce��)�(\h��)R�'�ȯV�x�Ԇ^۰�h��9Yng+t���	�T��Xޜ��	-�W�)SŽ����$N��\7,=�萴G��o�Vj�6�w�L ��.����1�Sa���g�����M	_���r��J�Y��E��D�8�: �[K�l9G����t�]�sH��-9X2*�%�s�1�}J�$�;�&M/Ы�&:��L�f�-V���v���]H��K�.!He
0PK���d�41�늖�X���Z>p�wN`)ӟ��}�穋��rK���!۪�����A����M�]ր����Nj!��LͽUm^WeXx��(F�w���Y`{T��J����{��� ���>MV�-WK�uc�^�,x`�[�#¸_���b�Ze�WI�	:ߕ��ܲ+�|~���j� �Q�~�+>Y╇�^��9`)����<ն�;���ڽ�;�=r{B5�"ܠ��ÙQ\+�:����eu��j��g�U3��&b4�坍Mjv�ܿ�0�.��p�T0.Rŋ�#�0W�	:b��;�8]/j���Q\����t(fi���g�*Wj�*�Μ����>��~��o���b�����ЬBg�7~N������K9T�!���^��gYXX��jο�j�b[�7�-5���b��֯hz�u�b�W�2R�FS�%;�ș��Mn�%��3�w�z9�2\�>�v��9�
��o<�3��q#�w�<Q�Z^Yy8I6�\�Vm|I[����u��Pd�U�K�_��q��}���d��9��H6TR=�QkOA�Ȯ���n3q�!���D��EeJZm���ۈ���a��NSp���q���<#+�]��Xv/6:��M8:�4]빳��3���p>�-�c���#jM	�2V,���tM��k�����+�S,�	F�X�;�����?����5w�ۛm�]}P+8�{��yV��b���+��g��5��+wk����l�u�x}-c��|-�OL�&q����XƷY�cl�6���4�LSW}]#0,����M���n���	$v��V�<J|��1�M=�ꕋs����XM-��=p��'��`3ö��+Y��[��p �����>>o��Ǣ��1�]��Ǚ��ו1�4T4��-�`�O���E�tp��ZZK��̥�s�n-ۓ6�N�AR|�\H�ɗzo7]�R�v4�b�=צ��A�����Ք_ZE�@���A����4��UQ����99��o�D������@:F���F�n�i�k5q��=E:ʾ��7l�����z	S�K{���4ԫ�ʌڛ�_h�S{gzjAͻ�FR�{84�\L#�J4:���PW"''Jy�t���*\���f�7���a�:���R$4R2��fn�[���)P�yܟAfh�i���Q�杙9S{Vj��]ʮ���,��3j�[b�M�%�&~9N��ES���״3GQy��W57GAf�@�طie��԰�^��ݻ=P���n8M�Ȓ�0]�W�&�]��o*�����(ԃn$���v�K'^����t3����&�fr��9���'vB��'mD��徧�,>\bǍ��{n#�k����->	o��[;��,X�����,���{[�]mXU�V��)�\��vHt��=Yi/!�;|�
��Y�u`V�������KnⰔ9�/l��7������+���Q5�pc�p��v�% ���\�t��D�V�d2V��+�0�
�ŔG)��^���<��g8��5���eb�$taR4��S�;��̛�5��3+�K�f�yv��(�_C�u��:�1&u��T��z�1�1挃 �ac�f�r%s�2�1��բ�-B��M�L9oXOt�r�]re�zo��ӭI�k�q���w�!�5O4�pu;�6e�8�ݩK�y��ڒ5�wM�Y����j���|W7_��QOe��v�P��8�eS�eCF��%��\DALK���A��W�Ӏw)c3��u^_ ��eA�0�M)�k�>PvǴ}u� �Z��ɹS ���#,QW��W#-�{M����b�h��6��d�>5��LT�,Tݺ��*M�L��r(��T����AǪw^��w�I*;ؐ}��*t����N��C�G�r)77!�l�f$��Iڇ�ٶM&�Й6e�j��+U�s�K�(Ӫm��a�*)ӶV��P�
1C��gB�Q�֐�nѦ��k��nj�IZM8�b
*����Š�slf��UMh�<�4�b���"5�9��Z�i9h) �J�`)��b)*����c��.sq���l�ULUr5W3��PF�j.O**�[��i�m����lc�#r6�E�cZ6�F�͹͖j�5n�ȭ�F�5M󆹂���4P��0UAEV��4ڊ+lE0E�j"b#cDRS�U�[U�F˨ذcb�Z�lh"")�+F�����T���D�Em�&b�C��
 U��,�ݻ.L�A���u��OfRk�δk�`5g4��9Y Y�e�Ҋ�y,RW�	�I��*]A��oef�����c=�����P�zj�{���e*�����7 Mg�L!�2�<�XP��P���= j��Sy��с�n�1�Qa�D�� X����|���_:w0��=ʧ�Y��Ȟ�)�ԧ�w��~�㚨V5Tp�Z%�܍v��WP��uPE S�r]�X>;t��5w��E�te�=f�6\l�+s�h�_m}Q	S���ܑ	����_��Dt����9�X#©�-����%YN�D���b�B��|{���������!Aׂ�����I#r��w��$���er8=��x
:]=���Ȕ����*�-˩=��e\��h��n�}�:�Ҡd�leWS̭�Λ��Q}m|A�e˱�p����c�h��Y�2�k��t��Z�N����*NI����'�L��T��+�|�n��h�
�s�lP|={��3�88��[�B������1@�I��;n�|o7j��K�3�U؜�[�9�x�|��=c�Y������UE� ��S ,�f��0�\O����*���Ɣ�E	�Ѳ'��N�e���z%����<��T�`^Ң�Vzuk��Yc1���	\w.�����;ʇcʕ<0g6��%�g���n������͕u�M[E:S;ά7�N�%&�h�<�NސQ���1�t���힙�_����!#��m���ó����2k�1z��͵Ẃ�2�G���Q�!�ݍg{9N-�z����
W�U��Ů�^y�QXve��+O ��n�g����r#(�Qb�щWK_*��$u�fh�|@��T��U��_�0��}1�{q�h�p$��p��Գ�Ft���85���#�~�̽=b�q0����}s8��!C��7�x��vu6�+����5$p��]����`ۆ�}�W�ѷ�k��ϩ?���ι��q{���`k)���+�
&�"�*��5K��L�˔48�Z���j���l�*�SHR��z����3,�[���S��u1�8ܡ/�V�+�i���-�C���K�+-�T�=�^����']�X��`n$D���?���5,������N�0�b��#O���%��QC7�nz����#���(3�R#�d��9<"
�ez��g\ߋ߻~~�\�J����U������T���:�7Nb,�[Vi{��GGd������'������me%#�R���Axor�jb���[J��u,���[���˂ϝ꾡�	�)ƦZU��xrc\�7k�W>���[��P\��G�T+;-���FC��v*A����`��N�C� ���S�[�Lx����e�8s����}�}��Vd|��{UVi���HE�k'�Y�P�dH��.���� MT��U�1�*��ћ�;��L�B=v��O�1�'����U��^�l�`�o,
�n�a�3���u��t[/��d���<x�"?�R�
ۭ��v�;��`S�x��qUv��ݡ�Y̩է�g#�� �A�ܷ�C�+-xaI����E?��T�jg]�Q�P�N\����]Y�w ��T�x��ǯL��a+~�R��:�7��0�Ш�����ݬ{�-Iq5�����Ȱԯp
��պ����xAaY_/
/q�"�ɧ�;���of�6&�d� 6�Z:t*��MＯU���bW��ߍ�WQ�l!;��YHw����� M8�`���������u<$lc�_%rt���i��(m>����&�kCT��ƣ
���^F�x��������2�����ٌ�?Yޮ���Ù�r>�B]W7�p��?o�a��4�n\��'���]�B�U�ߊ.f#��ͩ��'�;��wgso�h�LE����W��,�`;Έ��~�Nު�.���!��U*�Ap�����\�l�$-� &��*Ԧ�99��o�M�*bqT��yc8�K;P����U� �o�>»}�'� ��ꞩu��r��V�L�w�����D6�5]��w�Y���.s��H��xmZZ=*�t���0O��x�f���j��R�p�̉�J�o
+o��4B��qN�� =�3=TFꨌ�ќCK�rN�P���\SP�Sٿ?�	�;�X%;ydt�W�� ls$0�R�M����s�`-�X�4vZ�A����bـ,d:�)Sc!d@!��F���fmįqm�$Y��=�G+���IǾ�w��-ϝ��$I}�śW�eR��B���"�j�(�.g���{�ci��X9�����o|wNA+$��p�+�0��fKD��Yۚl����r�v2���M�V䉀�a�xs`2�P0��Nc����#�����U�����ܹ���Q� ?��TQ&Mh��t߭Վqxb/���i����n����;��x��H+���y��g�;l�&d�ӒZ;su�Y�0���ڧA�!��&��LLZM�y�h��M�	�EØ�v���ŕb���O��CNJX�ʿc��.E��fg�ߖ�-7�v�{��>{��Ej쉟tY���v��!��>�T�-z�Z�M��Q�+ G�7�sޫ��3���P+Z-�>Ω6���qeڷ��g1�)��Ī���ˁ.Av�d��JŨ�Q���j���0�T��4MT����>�>N���%����C�"�����	E�J���bx�5;��g��t�D vtl�!4Nn�q��z�v-�8t�9;�#Р_b�(1l�J���}}qV^Їe��Y�kASsʳ�n�����oYg�KiX�)�vz}i?e}��m1��������u�P$�[����T.�oy�ENo��(�,h��U�2�QN�ħj�u������y�M�1�´���\�`�)�?r�p�R/M_�l��~��U��ƧQ����B�ɘB�C��ڸ�6&�ŵ���R�8)�0>�/L(e�upC��6����b~�����˧W��%.+')��z��\U���k�4O8��Uj�����;���pi�^�@c�m���Ϳ)�z��X�8�sOk�U��ԓ��|�H�G���J��s�1��U��$���9]��Q�^UrŤv�d/�`�9���_�3��|i��u�i{-�!l��UA�?:�WV9쓒�Uq(\9��*&x�F��V<P��{�B^B/�`˽���.3�6�+�Z6���^��e��춯a��>�巊#%p�)jw�H��i�[6�K59ت�� Okt'Pm�۝H}��t���]m�:+�g3���ZS�Ҳ�b�1��6�vV2+�Ŏ��?}_}�W�Qq^���*}�b:�]�թ�$�蔏d~Da�`�{�� ������L�G�z��&�ӫ$�-�u��=�A��yO������Ծ|�f�t���1W\VO�O�ѫ�:	�[����ԋg.~��yS��T��!���b����P�mP�����6@��tQ�5,v��g��+�/6<�����9��x���l*B!�����5L�6 F��̰��6m�c�5F����w5U�~��ו�/Y�Aq`ؔ�yb��;�}��Y9��d��YΗT��aw�Z���N���]�E���m:�v�g��.f�¬�+�Z2��FP~�G־L����5� ���z�Y��(Κ7^~Y�Uz���xjT}㘚��8a��@fK�
���EU��_�0ꯐ�ƞ���s원�W��l�v�O{k��u�c>�����_Ϲ��1c0��!P���u�x�,zu7�h!0����8c�]Pcq�5L1������3=��v�yV0��S��i�Kq���S����U �4O��TF���Cr���t��Vu��]DG=�%E�7�βޙ[�Ɛ�jvq8�7i�INfI�l��)s�9�z:m-��u1�ټԗ�/�j�ȩ�2����f�u~���[V�~p7�I��]�e�d�l])U��&��Ԓ!�hmX�f�����{fS��p*z�+O����\�	�����B1��R�M���U�G�C��:	���dX�ڈ��+���N^�!�¸�{k��J}hK�<��+�eK��ְ��6�X�'�N��\���*�mD�@U��^:�N�0�h*\W�����y�kq&��-ns�2�?	~�m��[�[5Aa&�=/�T;+�Jθ^}��^��7����fY�W� �w�üOWU��v�>�f���M�42i�h:j�v�>��Ԛ�wF?������Xvt�n���$��"&���D�M�̐]_aO�o=��T��
�Hƚ�#�,k{V�Y,A�<� ��]H��H�7��u9x���e��?p��F<V����|M@�Pϻ��)�@4K��$S%��j3m�̫P���b�䝦n����^Oʋ�6P�2�J��K}#���*QB��Q��;oa�ծ��iP�Q&�FXl�c�+�a+x<UJ6�8���D%G���e���1I1�A�5t��ǎ�^�8�dXj{�[fR?h��\>��J����1�E`[�_i>�S�I��q �
/�2�e�;�F4xPչC(��p�ݨ���vZ�951���`�p���O��q�=i��i��K� wal�ćRv!wwx��V�4n��R;��K��������><�I����l{P3J�X-�����'b����%A�D}}��Gf�7�îu\��_e�:���_�*!����]���F�J����ح~l�@�F}x�v�E�8��� ����@χ#l�7Z!�N�����Z7!�h��a�Eab{}nA���;����6w>�����\f b�S�N3ft5o��4SsD���o�^�R>� �w�a���&��+�&t�Qf)�d.��ە-��Du&$=�=KA��S%㬲F�4���|g���)(9�\^����%��ߺ��u�oP�%5l�3��f���\n%ͣ��L!�K��*m�p�U�OV���½��N���̍������
����|l0,�N���O�Y���'hu���k��5�T5ndN[X���]��=`��K&5;���*u�q���r
f��_7L�,%��&��n��gnj�A�s���<��F��Le�V���p^V���@!�d_�I�#������LbW<��0!�Ĺ�s|wN��BM_��9���L�۹-�^�>`p�ķ2��+l����"��v�aq/��k}]X#����t�[�H
�����f�V,�iԶ�*ιY+nb��pH�^+ʊ�[�/a�r�s5��u��H�M�8r��ԋ�}Vn�=�z���jrU�h�{ﾏ��>�ҍ���3E1L =`T�^�(`�7A�+�|��z��t�_e]v���R-����{�U=y���C�s�g�/+�}����7I�ёG]r�X�U�"�p������,=]��zj���)(1�6a5!��,;F����+�0�}~?{/ް�"&�rWj���z��.�zz����}6�i�FD7��2�K�g�F���̮��;���:z�Lm�0�RΫő�uA:��@���:eU0�`7�%T���𖕚�R������o������Uo\(�$w�fi��K϶إ������?!ПgdW�]%��>�%����P{��dC�s�j���TM+1�(��b��⨾]avw�a�)o:K~~����С{��=�J�w�b�W�fJY�#)�x���:��F�c�'!w3�'����-�3Z~k����h����d����:�EM�X�0�^D�Fa�����	����}�2�֛�;���L����S��Ү�t7�UƱ׼��*�*�Ⱦt8;�iXE�W9W��s�V>�v��}�K7�l7y����E�7��)�d��R�t�^�N������b�{�횢�uo����cm7ʳ�u���<�q@�pmr�x�&�<ݖ�9�>ٕ(�.�>��hcv)�9I)%5�l0�S5S�����>�2ީ�����.���j��f@�Q��h��r5���ʆ,�S$�_M!���ʇw������q'�+K�efL.*"�k䜤P�n�;�
�"��۪��(�ww�h�S�TT�t����ۊ�z_�:^w�μ�w���𐎠�����\��-^$h$�eȫ�v䱦!0`�Jg�ȥ0� �Y��9K������0���)��c�����!>p����p3��U��x��8e�1��E}�X��n��Y܋�ɦ��vvBg���gJ����a���1�A��i�V�[�~;
���]�����U�Z:!M}��}�b��,EԀ����d��cMK��F��خ^���G����nCy�A�Ʉ�DwfZʨ�p F��2ð��7���GL�%���5��f���ɿ���k����~�k)��⓬5G5�W���.�}�ﷅ�y�et-��G6�Z��o[6e{�&�1�4[V�\�ׅt67|�yM<뒫k��\�k�y��Z��GЄ�v�Ѿ��9֫33��&�n���g�t�D�rޭvc���N�c�����j�WRp��ν9DR�79g�j�07p����lV�V����o"�u 7����5��i`��{4�(uؔ#ڻ2�-E2"�H���H���ڕ�^������em`�{֭�U;&�%���޾>â{m��(Gw��ɢ)�i�z�2=u���v��`�t��d�w��N4͑��t���ð�.�{G���E~��+�7ON.�~��iQE���K��,�pIs�^IͶh��`Ѷ�MȢh��ZZ��Q�$d���kM�5G�/_^$�܉+��/�����z�>��7ٗNA�&ڳ�����7�wwXYՎ(���CU�Ǒ�<0��u(V�iJH�\߉m/������v���\kf�8�ƣ��g6�r@.�n�Y!����ں���]�H��p���U�y$��><m
�z1�5�>ԴeZt���V��R�
�F�%͗gsQ����*q�T�੣olCֶ��{�{Fe���i%���p-��>���5S+�f�H���N�� .��뙕EhA]�q%4y��X1��قpnq�Κ31F�.�2-�Z+-k`�8h���F�fU�uėlL��R]#%�&���>�G���b�"�Vr����k�&-w(Y������ä�'�����0�s����۰�.#�����H�ꇮ���xz�/�<΋�M͂����}Z��,��b��05���x�.�u�J�f!�C���&�������sX<��5���,�HpNIpEk�lH�ݔ$!��q�᰺��עX/	�#N�Ԃ���"���[Hެ�oNS���2�������$;R��D�η�I��G/���W�=��6e��Y3H�pR����Ӑ씶[�J��N���˹Ӽs�kA�=��2�|U"�٘�Z��m9y-*u�y����;a��K4����`�-E��o�@Գ���0
�U�����U�)r���2^�6H�3a� rDs�R�љ/��uإ�Li��QL�P���-��]3ii�v�	��Z+f��wb8����C��Z2���/;�T9�-�ʠʯHWל͂�E=�d�u2��rl�P�Ȯ��:�6s��]�U
����o8U\��{�%'ZN���^��[^�C]��Mn5�N� �m<�7���=b_���;���z���x�:�E�X�u,����y�1�]��ۭi�ۤH�U(�9j�V�a5�h@+�+x�i�K�' xQ`tu�oS&u�D�\dʄ���b�}��R�QJ����N�Sj]��-�ڜ�3 ����ګo���i��LW�A˸i���������s|��߽~��������1RA4�Tlj&�!՝�4PQN��i��`�UE5DE4�ILAQQDEPZ�QQ��gF��Y"(���(*�:�&&�"��J��5UDDm�j ��+X�&��b)v�EV�Z0U�4��*f*��cUA43E����-��5m��c[cY�$����&�8��Z�:%�a���
�g�Nڨ&�t[Z5QQV��rP�mY���QEUT�13EE��0TU3�jƂ��4h#cTDAEح��b-kmZԑEUX��U�T�&"th��V5U4�EU�Z�٪�`���"
�*�����)B�p[|�ZL�|7;��616r�
g<��[Y͆�$>�<J�:������d�e#�Rrb�!�ۤ��>�gB3�Ə�����޶��&qN��s�G���IXτf�v�5Au�X�q[� �X��O7ރ��ݼ�JW�Iu*�������EܶbӔ:�����.5�=�����t.�������0j����5^l����3ﴚ��;zr#[�Cq�`�k/��W](���S��'���N�c�u����w�|�`^��w�ĺ�k�g�[�ʹ6,q�Lt��C����� ,���V�fV�+.�Ϧ��(�]Q��VA�	��V�+�ʖ����6ܱt.�W���zѽ�\�HS�T��5�A��mT���U +��(uD06��F���t;����9�^5~�M@S�^��[*�t,���y��@\��@	,97k"���|_)��g�o8,p�Oc9!���������1]��[n$RY����p1ͽ*��P��!<�TN}�M.���LN;)i���fG9�>���������q5�z���M����x;D�̰ў"݊;wklU�s�u�ǽ/)r�q?J�����5c��]ٜ������/�����ݬ��y����ٙ3��A_#��GRv�cn�A"�՟u`cyl�b�В�ɺ�3�v ���xYq��7r����Y&���MTj�nX��t�4�E�W?}��}��}�+��)z��r��ձ\���������F$ˑ�e����N�xWv̥��i����vu�}W���`�o����!�MΘ���U�$f��]8�"Wףތ��R���=~v2�QП7��l[����'a�ܞӡ�&�SS�	=,�lߪAq>}
�͋����R�x�H���g�p	Bǻ���N�"/C'����nE�V�QZDb���>��V�)M���ŭ�\d�z�b�[��o7�<Ci;y��	3��Y���S���\�3:E)�1�;�s�����r��#Sb�y�J�بzE��0�����8;W�E�S�i\�:�jV�VqX|��T�w���s.W���R�y!�oK��;�8�Q���|�$MAމz�cq��j��nd#޾ܘs}���	&�<�u�{�̦��|pX-��ќ�}��r��N�x�4/h�����o*�c
�'@0�� fD���,��Sx�&�|P�t2�<���=�V�|+ii�y�Q�[3%�4��o��Roov���8��gx�2T��p��ߠ��g��C�[)mk�yٕ�z��+r��v,h�(W���>��F�c�*u�C}�Nm����
\�3�q�V�7	���wܷ�O� �{�{����U9s^�)�7^gw��w?3��	�����Q9�O̽�}��.����+L&��x
|���u�; 躛'�"<��.�K�܊��uq��½T�9��Ϩ��U9 ��:K�8
���Վ��
��M�Y����2���t	�AP_D�o-���o˼پ8��o�<m�»V@�w�<���x_D'�w��]�D����������P�;B�;/7����p�b�4���6��%�:�}�m��*TU:���B��fqj8M�N9�3��+�z�8{�5�p�v>�8��UQ� ��d��q�g�JE{��}���g���x&�pH�{qVOm�P���͜kf��n;��ɞe`L)�{��}�ڑn��DxE�SLn���gk�V�щ6c�/G�z�ujծ.�m��U��w�NH����]�ӭ�����4�r���)/X�hn�IZ+j-����8�sC\�*�Wʮ�I�+�O3���-��^���">��r��f]��Շ���m����s�]����+���_H���W�Ufo��4Q{hLPt��t{K�>F���W��oi��p�țߌk�m+�1�x��4��C���U�pގ녱*��D�hGۯE���㞰��{��u��llNQ�nm�MLիk{�&Н\�r8w(s�<���x��e��Zۿ�%uF�T5wZ��q�,�:�M�fWhC	�1A�w��1�|����zY�q<޵8zM�]9q�Ɋʷ<om��45!l�S\]��"5v������?/Mo�/0�5�5��Ԟ�v:�o�
�ͨΨ�Y�R�1t�<%k��.̰�d���[`�^L������ΕIC�7
`;�\Y��oi��LJܘ����j�h���E�F���0�M�;��>�*㛨ϩS<,����U�����ջ�ty��*f�����A՗pw�ݭ^��x'��p;�ŵ��T�z�û�R����bN�2	A���9�����g ly�b!�Z}_��H���F�n;�'���z�N�����[�+Ӛ���:S��ۥ�PW�N�����3�-��b�5�VkA�?�}�}�UL嘼qK5�}��3�,��y�AV�*�oT4��`�N�s}�jxhR'j�e8�FV��<�ϼ����!8~�����j`����n�*Nk�s3{fގ@R�.���Õ����߯1�ד����n�N8.,��v���)�{Z�v�l��R۫�y�qʵg�,����^y�0�k1�G�Td�9��쾕�S�����ס��j׸�O��*�8qv�=�n��͞������9X���A]#����w�&��ڮ^c�Unnt��x�dk!����he�h�_[�Z���}���{�3�z;������{O�CŜz�;�C_�P~��UyTY|�5J��)ҧkq��L���ው�c)��z���]�X=-����No�"��]���p�>�m�J�ܞA��nVf��g)�X���)c��}��	E�k�WL����\��{W$Y�w���^T���Z�c���9c�����
}Q�l�
^�T��b��Gw"����\��]��!��˽f�������Kl�K�:��K�����6w��K�w÷�w��DEa��!�3���WoE]#�>���j�=\��:���r�q��[���*OL}ws5� ���S9����_�3�un˸��>݁Ŵ�D�22IO�}CZ��&�v���?/,��k4�&O��>���m�w���U��3�)F9��L_mEc��Cyv�	J�w�8�ٖ̅Y��;�5�n^~&�v�R�4�gU{��Z�/w��^5�J����54<C{)���)�Bt&�t6\��7�n��Rc�ö���&��2-)q����.�ss�����%�_��ע-+*/&����t���X[�/-l^=�נ�"�!;ͣ�ewS<t?�)�������s�y��v���E��O�c�����O�=��4��𿳱��lilj�g�-�^�+,癰Z�ͯN[�_�'Ҝ�v�g�{�������s������8���G�z��L� ��`Iz���k��_*���PO�b�.J	,���]��ٲ������#��G_#�`��R���xvޣ�����gF�������Ӱ�5��z�'����.�)�0��e�n䇽�,�[����RRG`n&_���#�QZ۰��=ï�9�o�y78�c��K�͊���t�ط�VT�z�n�Q�u<��댰��u�EkYqU���T����n��wFB�=��[�k���oC�{��D�r�}8��;NwoǼ��p���j��#��_���W,A< kN�)}7sK���p��Ob��}�(���s��G.��w��'��B]�"���;<k����:�w����t����K���s��ܢ˖V�Uu�=Ew􉧈U��@��y�����.�����Yod6��	�V���*��4��(k�a&/�BP��W?w�ҵ�ٚ����9�r0��'Nu]MZ�C�5�\AK#�8�w,ƞ���J��	��
~;�}�l��U� �����9Ұ�>�+�G���z��~^I�ٽ��ǔV���V���j��X��Q�(��1}���Spf�tFL(�)���V�4;]:�^��F����/XV�͍��:T:�zS�ul���;��S��s��N�v���Q61J�ɩ��h��Jj����#�ފ{�w=��|�M5e_ȇ0�CwM�(���+��O�sWqG��27&�#�cb�'�嵽��bs��ީ)����C��gA��e��+3�<=)>�^���7�N+Lw�w�Kl�'Rq4I�Lz��-g��6�9�%����+���w�S ��9�M�����*��՟fFz)�x	��ͥ��ܭ�C�T8�|S�Z��O ۉ��R�7Yg���Α��y�lN����%}Ƈ��q���*��e�UwXRQo'���]���P��-I���[�;}PUvU��wT-�H�"j2�3$�.��_�͟x}W���I�GN4���ߑ�9�o�/��TY�qĩf�o���F���O���r�'��`�'F����4��19g��㛐HA���ڞ��-l7ʔP������Pʅ�&�\2-5��b�}	4��K���z6��V�N;�1y�}6f�9�o��Ǐ��y�vm..}���He�Ԍ�E�h�6��u���K%�}�s���e0@�-����fgi!��3�e���9���L ��|�s޷Ү桮�S"����	�l8�)�d���և	[��������B���Љ�ϫ����`K�W�Hת�.w���R�6|ݫ���}ro�R�X���gp��*+���a��+��ekˈy�_�U���M�:%DO5�x���RӮ�CȽ`������+{{)�
�w;��Y���In�s�r.�j��z��/!S�1*��XX��7ӱ1�"s<�7���t^+n=�#9YMC��w�*��6��|T۴n1\_E�w�ZN��{�6:7���7����}�/6�w]������ox`��TՄ���l�]��<�?<�W���r�xL_��&�TGdc.�ق�ot5i��n�&�8$T�N�՗,��5��+
j��PsG��������5���Ξ�Ugz)��=�p�T?g8��5
A�o.�y�t��p�/�+g<�'*x����rW���W5N�%!����c.w�����a��n��B������Cbʇ�'���郈��s�<�]�%lT4��Ǣ�ĳ��iAڲ�WY׬j-�5L���fQ:�6X�9�=n菹��R�.���v�A�pU��.K�� 6�[&
��p��Ovb� *�}}�7�-�Y�l��;�������J���v���C��imC]����_k�ҝ�D�Ul�//I��I�E�ZՎ[_=Ew�5<m>�M�({c��!R��{{נ�d�n@5���^|�W3��c��o�q���ϧ��#��E�Ӥ��r�ھǮ�#��z1۶��e<p�Å���	D�5*#+yD���Y�sO��V�#�߾�]��?I�{�x�;��k��:���`b�u�NW�w[/�r��WI�M���a|�8�=���̖��o9�b�u�Ns��\)�b�n�j̆�1(S��y����_<�1JQ�u(�ɼ���]�𴍅�a#�VԼ8�x��2t~���IG*:��Z��{�f�^aZ�h�q��PN� ��~�V~MM��7��r��&ۧ�nt���C�:����<�Ws��(�nC:ܻ�=�U��������$�Omo�<�[βL΋%�,�qsie���$Rn4)�G&��i�FL�%&�A�xϝ�t��y={>[5k��&�X琬͓n.�4���[[��ɾ����:ܸV2'q�'X�%t�L�p������6�T�o{P;�wGk5q����6�I�̺��D�!}�R�η1_�����J+S���Ko+(s��,	�����x�!]�2��F��N�� JMm(WV�pϳ�l_��gK�q��ˈ���Fv�ҹ��i?;,�̯�.�{��E2�v��j��{WY�솉�9��'1��Z���l���W��n2ճ�D�.���2�ï%�OQ���F�ĥ�f�|0� eӒ�,�ᮦ�v�����V#�t�g`�9��t@�V8�_AtށnK�*��n�0έ;����wt�1�[{Sv<E�#.�8|;Fƫ�=q`��Ę������|g&�E�}2b�Q:|(�oyo��� I�`%o^�1�f�,�W��BF��0b��_�|���1�7y��*�a*i���gV<�*��-�8F�槆�ݎ,�ù}�HS��S�)��Y[��%�k-����d;B|oJ��/O�/�����m�2�98a���p'8�LV𧽼�W�)�[��P�nl4O��Z#��x�td�J���}H��X�lٺ�"��!������kXf���N�����)Vʶus�E�W��)7eD��8�N���fK��� �Dx�S��vd�dҞ��T�m�fsX��/�6��]Kdo]�p��MVYQ^I��)g:<�82P�1����"��xś(��4��v�`e톩�Y�u�%���c���۫�aͬ)�%�n2w���#J��!����DN�V��[��Y�ց�m���(=�DS��XQ�}��WӸc9�6c�t�7fűD��.)�A�c��E�)�¾b��C�����im}�z���7r�`'{��L�i�a�=|i�v�eX�ɃՈ
cj���k:�L�H{j&��1t���Ғa��n(�ւ��y��F�m����^�=㑌���=�����am _A[�k)X �b��-��7�k�7�A�FejJ+��=ZEne�lx{t�f�w��g���G
�K��"�X�p�]�α���bu���ݛt�X�u��v��J�ڴ�NHy���.�����U|�W�Z2���s�V�u�NnM�����
�ԇ�S���1��q��yq��CǬO��.�4`����Ġ���U��!�C�+��Pmݽ�'�fz$N��=7�i���8S��=ދ�Zm+3Gv��ꊜ����UZ�r���T��_,���-��o�,J�w!2��BGH�Ξ+������,`ӹrA��{;��qW*�l�.�.l�5i�U��mw�S�
�����F��ɒGc��vx�����6�}ƺEv�m�n�<���ɠ��7��;:�d�:G�Y�9�v�wb�����voc�ޛ�j֕}DS���u����:Bjj���EF�T�A�F�@h�4T4Di�1UES[h�l�DETM�AASNڒ"Md��M�J��(�%��&�4N���QV�SPQQ%TV�-&"����5Z5UELh�3M$DTUT�k%Fƚ����"��I���i�*�ccU�( �l�4�D�D�E:�DT�U�)A�SV٭+mQN����TUDL�LQ!T�%QD�F�IMlb�bi(b�KF�)�EX�"	��SCAQDTU4�TRPST�V�QPUQ1Ph�CZIl�Ӧ�ֈ�l�PЦ�f"h������PQDEAQST�%4PQ�4DT;j*�� |  *��w\�X�nk�݄�3�93^Ȳ���5�<'��p����띘Q��tܽ�Nn�j�Lw!�+-�yR����P�ʯ����Fd��k��b#?,j'������-���ߊ]�W�����]e��V��c�ѶZp_SZ�q�x�7�5�S�6Î�9���T�x�ۭ�v&&���=I�,�
V<���zp�|����/q���*���橷H�.���ͨ��Q�1����i[Sm��j�WM#ke�oWKxZȸ���W��{�s�>8�H^ߗG*��\ثi��o,��>�8���i��܆�����\��%}���O�~����W�S����i'�1F�`e�S��}�W�!�\����^|����w�zu�^�����{F�ԗ�j
>��}ښ�I7 ����C�	��kN`D�Ys��Y!�`�	r�C�nj����S�C�wd$�ǻP�:�a+�1�U�U�}qY,��D�j��F�Ţ-�{X���'�n�s�����@����Cp��m���f��I��q�ڄ�CP�F�C�����Ց6���\�S����Qt�ΗtFҋe�8�啧Qt���.�\�� ��aab�j����((�v�w� �P�q���9��kn�8�i�*臛,�j�uH�'j���aۮa����f.S��_}�Ͱ�E��x��9ЎY_OL���uէu��-n�y���jD���K�������I�]|�0�>��TO	Z�>����t����z(5-ܘ������F˸����)f+D��bWd�y�6�8{�ѥ*����QG��v�����L��_� ������/?{�)d��ZH��`9�z����I���_�����FD4]Ao��zd�b�B���[3�!�U�j5�8�*��]�=Q�L�1�* 8kR|��v���C�ַ�����V'6�k;�#v��9�zH7�ҩ/�Y������7h��R��}���Z~�����
`���\���/.�0�SN��q�]�W�_���{˂v�{��"�J��]�B�Qj�Mek�p#X�t�d,�\���ux�n-zz�f�����_R�2f�@���w�Hl<�V��-�_	N\��yRF��X��E�V�ۃFph�[*\�q��mq�h��Aq]G�7H�Q���F���҃���-�(=[p�3�t ��]}�Ե٬.#H+���6N��zX-͠`��mF�nI�#19�|��<v�a�����UxOR��i����3��;���swo���;}G���k�,�6
���D���T�؜68ƹ3�{�u�P��s���j�_iO-�>����W�ڨ���2��ܦ�������rsj�p�f���c|�n1�_J��snz���sEt���oL7
�I�)p���b��[	4�jnic��o�K���cH��J2~�t���*��Ϯ:���/.�OZ���m�uH�K�����n⨇�f���C]9a�V��#m�k��Y�ցf�(����1����Þ�š���z�O��:;]�(�[X%>2����5C��P���&.�s��£��A�j_S�hi�*�3w��w��}~՞UȬ���k��o��8'z
���o�����S�VY��0��w3T���J�\�*]�	�����G�ź�E�euwC�V�RؖU���M�<շ�n�,`p:��O���xf_w#�d��Dg:W�/ּ��[�]8\f|��S�pf�)ՕZa����L��v\�%]���"���N,/HYȍN��n�ݾ�m�D���;��tw\RCnfϢ>�#5f;������ӎñU�/�,�����ﲯ1����f1Gq��QKa󲷆.�mM�N3�{^���䊖N�՗*O���+��:�J��M�Ā�4 ۋp~뮊��6u(��gj�����<���^H�}�s'Mޅ�G�{��X=��rjq�k�T����P�g�QṳW���R��'�b���[n9hW��ˌi��w�_5khm��x����:p����'��C�"j+Z�<�,�w�UO.��X2f�R(���ڼ��.?7�:����Ň�>����.f�ZltÁ1|1�V�g6n��k�����o����JeB�*�Q?WsR�������=P�[g�WP�Ky�i_�5�E�5�猳�r��O8��δ'�$�,<E������W���UAO��O8+�?Oc8$2ߕ��>����=��Hɧ��	�I�z��f����#��=����nÚ[�π&l�����7�%K����'��{�xtg�^c��4����)�m��7�P�x+�I�k.>�a�����PW<y��#�Z%�է�l��/��][�뺲*������H{����4[�V��+^����p��`'1۪��7���V�)����s�DէU��&�3�PF���"�[�	��W?w0��v&a\�ڳ�љH����f�{���C�G���/���Ɨ����}~�C��c�șY�^ܦ�Vj3��'�5���q
?=s�|}~�F�(��+���n��ׯ�R�$��j�[G+��K��.�\(�\]�*�&-�g.��R���1���z��Vwx���A6Z�&��x8�|9V� ��ST�k��p���V�C�Z
ms���ͼ��c;���s��5#�EK��W��/u��=��YS�K��%�x��)����������s���5�ޮꋨ��Y(��=��˽3Z��$��B׫���֦�=���ܥ
���xV��d���T�O�c[;k����9+�6��v��H������4�,!ר�+g��e�R��Z���.P�d�_3)��u�il��uiL��:j��A]΢d�z�LY�����F�R{�4>]xs+N	��"��ջpYΠo��6�G���L���N{| ��Z�b��B�S�7�ڗΣ�w�\؝UA�� �3ﾏ������UY��.52��}?ݖއ��ؕ_)�����w���+��&�w�,�Q�Χ��O.��q�����m�u��K���������&'�>6H|�2'���=���A��:������]Z��US:���1в�$���-s�	�^�x�� �~
3���)�����s�ɶD�����CZ�x�s��컈��PZڱ���)~OkW�t���3�=�f��C_r���b3���D�������������O��|���nb�q�p	�]L���F3,`�O����`ȅo=���>�r5���q��^�>IӰ�>���u�uΜ�/�ͬ��<r�9����^���r��';QC�lD��}֧Is��WG�}zS��V����u�S7����,�Sɭfէ���f�ɽ{%�:^#m\{mY*ͩFZz�$�S�|}�Whn�;F��;]�{[��U�Ts�+�ӊ��m<���tU����.�ޏ]c�ݪ@������ٵ'Z���J�
Л�7��U[�m�e����&����̵,�{�N<%�k�wX���\,u������\+����:/?|������|y��w�t�����ԫ�]��Mv�V��x��=� ��ź���j����X>J1ꋱ$Pc��=�����l8�������xv����_lJ���c�/+1a��۬�-g*ڙ��\�z�WͣU��x�g���߇�\?g�T%+l��׶t11����Y|�4��������x�h����?s��W����ta*���No����5՞Ues��j����B��K}*���J�y�ͫq��X���R����b�(�|��J�{�����G<h�ׇ�m>�1)9M��3|ٰ�ᄪP����
�Mf.���´��p~�3��s�&�����Ә�[͹X#���$��}v;�\���]I	wW�!U��I8s����~P'X-��#�CZ���+�g=�;�}�K=l�Q%.�;��^{F�.��Mzބ"�]YtcB:�Y�0��-�
��'��u�_+��'3��0d��żc�������ċZ�gm�"��˷�b��8�<.�O1L�E��n{]Eߐ�7��nr���䭋�l�E������{5���X�nm^��JU��|�i�B8�[O��ʺ�Y��+���R{ĭ#�g�/�\�^��+������{�\���o����U�#M��i�5���Hl�~�+-Z�����6��-��qc��Y?m��&&bP߆溜]�e��q�����������G�Ѿ�tW��`������'J֛���Z�_1}d��{��78�+O�K/�>���ﲯ1����Cj֜�3֖�맚�q�$܋�&k�d�0e|���Z��ޣ�Z69�S�Y���J
X���Q�:�Ew=|1��|fo����m߫L���q�^n�T�zwwpi�{�3�
`ۋ ��s�����9�׼8C��������̝n��ֻ��%p�x�����}S�����EG����n��h�w��d��}<��ɾ�ʑz�1�\5Y�*����tG��Jn���;B��<���"*�+��@�뢞{*K��	�'N
�˫��,дc"��MB{^\4�=ҏ]_7u������Ku�qɂg�7E�}=��E�Q�6N-0F�18�S٢D���
7c՗���l�Ź�t@��	��Y�ֽ��S���^�J�w�fi��Ԣ'>�`#���������z��X��'�8�?*�:��41�����.��xzyl�t�|1f^��5!��ojRw�o*�eB��M��F����ojY�)�9OKǽ5g�S�K4ҿ���0�7|m��гa�)���;\�k�5��޻��^.�*�sJ�4+�	ԩ��?b���dP��y�g�ܼ����"�Y55]�ٗ9���P�[���p�B焚�B�D��P�FO>�BI���	m�a��	[�	�¥�:�9�uwE��
Q��wmˁsvB�ƺ�f+�Ж٥�Ú�3��r�hw�=�і)��9���P��
�u�U�3�pi�ٵ��o���N�.��V4�q�FX���㍺�Zp{Q��3x+l+��h�q�N3�՘TսlɾB�%��7�q{����8�{�jʞvo!�r�a�Y`�C�8EHо@Y��pgn6�ջ�-+fҡȪ���CGn�F�fj��oHK�o�����8���-�Y�Yc41<�;g�R=�=w�+Ӂ>�/�D�;�hm���o7��A��Q�7��(Z)�u{�fN̪�6g%���)VJ'���ﾪ��o;���t�T����X�y��V�z�S�`֜��b@��m�yL���z/}�+��c��3}G�>��.���X_VC��Ϭc9� ���5��vO1}�p�^!��m�q�rʣ�����;X�]l�.�����ctm�|jC�r!��io>��a ��٨1Z�Y�:m��^ME��Uz5�ܫk5�r����kP��L��A6!}כ���׌8k�y�ړn�Wѹ�C��ڭTO.��pۍ��|���;SJ�5���Q�t��D�N����9:2��ۮ��F8�N��B�W7" ��I;��^�ʴ�9tv�9�pj�z�����x%��ܬ���Z���-nh����+��$ۡpN�s-�(6hsxx�s�﫢&�{[��n+SJ��=^+��۸5s�|98��<�4������G,�����]{d�Q�QO�fM
������8��`�R�}G�$�u���C~�6�>�8����;ڑ�O����3��_r�¤����Ϥ��[�$�G�q��,n����]��lj��m+��Fbp��ȭ�i����Y�w[�.q�R�'L�yofa�n���QZ����] ��\�����3q�=}��d��NG-۫�����:#�s`'0���R��\aN)����^�p�K�/5H{�-j�ڝ��0�ێ��칛�>�%�Y'Ną�J�`�R����o�]Lv'�F�=7�G#gN�M��[�a�1�����*�2�B��#��h71��]�;rVn}��3 �I��h�݊��=�++��xx*僠��ʊg��2ni�p�[��/J� S&��GY~d�^���|��P|�:�<UX�</��٠پl���X�,r�Z޼z���b�`Dkq1��-j5�7���r�]�������YBoē��������p�bs7A(ݓ�b���F�g�����'/�󕗒�Ad��^��q�:�S�"t��1�3n&(�ak�ݫWyG��pP����!�7�.�%��u�2�����/m�kNM]FZ1Wi��ԛ)�%��R3.�k}/e�lg��Ux���0ff�3���˫b�E�t�x��]��G.�?���b<z}q{4CW�Yvм��R��f����R��=��N�I���( iuK��k��Cwf+�{��únm��oM0ĸ[��1Oew`s
��͊�;���R�J���g6�h^��:u���m"Ad�Na8
���e2�1#��]М]�fW=����,ݙ��F��a�F��Lfi�ꣷ�$^��Tp5��I�-��tL�z{1�f��� �EO8շ}��ڸU��ѧ�|qu����� UKa�N�0�0�*���í�Zs�A����`V2����yh|�t��5�('pI��R�a��.�"�fu���W;�&T��#\�	�2)U�T4��z�N�����Z�<t���=xO'�<�x�G5L������.�K�֭B���-=�A>��HOe�.���Gz�px(7���|�C��[����4��Ud�.;���.PP��`�F��{1,�w8��Ǻ���-u?^֛�ٵ����f��SMo�j�H�L�Ӄ �. ^Lyo�&원L��m�rՀJcC�u>~e�G���U�l���i��r�˻�6�@��(u:�n&�^|7F*t�����2�*f�2��j��t��y�L���M_$|��Z;�����ރ�+]���'�9�d������d:�u�j����KDjdkY�t�AjU�A���Y֡�8%}��I�NF�Ө`�*�Լ,sz�v��d��8��tGn���[����QJ�8�\���֏N�����]]�6ي�*����UTQ1URRMSU3٪
m��`������*m8!�b4节��%�j���DA�LM%h"��.�5TDF�ACT�T��EQDCIBR�Ѡ�P�4�4R4��i�SQQ50�5ERSVäi�����UQ٠�"�b*�h��v�Eh6������q-3kLM!LE�m����HD:�C��$E45	TME	IDBE�TR�!AKDMP�M	ISlj�8���))ib���Jh�)��l�PCTUES%�D��	AQ1IICMQHQl&��J���T}J>���	.uث.�05$��UIxE��Z�� �1��t�-r�ݠ��Qp#�m� B��m=G���<\ܪ�;�56��V�ቚ��u|���LD��f�T[
҄U=�k�����3���ٹ�u�F�������*` t�z��/Ux�zP`�`�|*n̎Al�J����}�չZ�c����Hu�z��)�:D���;ې8�gb���0,�Z)^^b���F�c�~���jz��_�
��^j��̼���-�:�����+�y�������{A�k����l�oq�v��R��]�~�W�qӊ�R�w�-�D��oj�������N)RC[]O��W�8��X��7)t_E|��f�,�CbS�we�y̌���ci쯯Z��x����W%}�y+�����YY�A��4
n�TY�Qe�+jKy��7�ܕZ���:N���em���Q�*��9L��=��mc�"'m���Ƕ��#U�="������WK����=���A�
��>WLo�M�Zx�z |���`5�ǘ{�R��=�_.����k�)uf���R�.�;:����� ��WC`qA�V����&�l����u}��s��n�q'�'7��F;�'^0�5���Ckf5S�m�Lz>�9}��	֝]^�#�AoY��������϶ko��!R�CťuL[��*
6i�Z9��a+��P���K�&�F.&�Ȫ�Ro�;Rs�/����ܮ1�K�J��zP����m_�̀hs��71�i@��3I�yz^����в�]]q��a�|!,rQ��:��樲��M]����u�{EHC}���不]�$���x�X���ɢ�4�K��1���Gs�	�W�z� �����s��i��}����&��.
�Ɗ�
���b��eA���m<8����'5�u���F��V:���f�y'Q����p���Vʛ�O�S��[x����NVbo5΋@�#')��u�ڜk�=m�=P�t��w��yg�{pw�W������m\n���"dN(�ŹTh�p_SW�užG��SP����u��v��B]��o��S��z�gZ�9����U�p�����%o�c������=���࿖�ܮ@c�L ��f`"���{���^F�F¶��dN�lc�:�>t��������KNT�9����-����c�uɋ]�d;�l�oV�bz�7���s��˽���I97��x�mL7�g߸v���&8�1����5{��x�h����t^�ʮ�a'��d����o`=������<��TLW+{9	�W;�����o�%\��^�)���C�\?g�U��B��}Q����I�=:My��-[�mX��Ev�fg�����k�,�*~+��1u�TY�V_;�*��B�=Bަ�`ր�tgm��K�!��*�.#V���ؕJT-���;�O��M�ߥo�{�:�i��ͥZy-϶���oj
��,ߞ�wc�f�cJBӉ�n��K5Q��r��E;
}O��|;s�d��7q��WW����dR�u�����zkڋDc��������IK �se�)���q]����^�{���n�cg���<H�]�ٖ�հ�[��GLXb;-�M[�oV����Y�e��Q��DFuYz��ă��P�s��)�P�M�Q��vs� �)��<0�f�.��"�����Y�XpC1mJMl���V�7�n�|h�1h��u����>��M�x(�fny1��z��R�6�O����p�Sk���N����	3uZ�����c�9<�è2������^5�ҡ�9YMM�b��B-}���k��d�p�QeSNP�*�����ho�5@�җ{z��\A4��턩O^�6�]�Ng��Wۺ�^rtڃ�N;�l�|]�p잴f�g����|�p�[i�=�נ�b�ަ�9MA�S�"Ý�]n��"�����YW.u���|���NȬ�9��X��u(���.#ͬ�V���˒�}����[�f}x2����x1U��UF(�Y������c��=-M�����ε��>X���ڭ�B�w�h��z�ϓ�%���k�x�[7��Sdu������'ku���f����5+Z�7�\�'x�F�]�t���:����6����l�|��"{�$j�,u�66�u3ϗWt��؟��+��P5<�����W�ڬ螨;��uw=����{o��f��W��-�'�v�5Ö:1ԏ>��ف	�`<V˧c~ڛ���`��%�O�3W���x��Iu�wGer�� ��;���#'I��Y�S���^�L��ux���`�;�N�&��Mz��fwIM�#�*��Z�9�Kh#r��a�@FwF|}ޚtq}�NY�+D��W~7�rv�>'�YX�W�)��G9��
���o�y�^	��ׁ�ܯW�uh>Ƕ6��Z������<a����_r��'��ς컌N��<Kl���u$WP���t�қ��L<��R�x��$�Pm`=V؟�_�6��<!V^�]�i�2��}�a�f˸��;3JY���.ۃK-b�ۼهD>{��j��K�v��Jsf��U9��	:w�z��/ LC�1�؞Vh��b�\��{��χ�x=6�P����5Htڇ�M������n�WM(ח��B�� 8���ݶm�^b���j�gu:�U:�!��c�#�����NZ}9�v�����D�õC��]���{���$Cmx|��v��.�sx�Nw�Ԏ}"���j�pr�����T�[�3X��wy�o{6=UW]��Ǣ_J���A��+j[��=2m�ҥ�5��MМ8ΡE/�CkZ.5c����+f[����?��=�J>�u�`No��JwSU,�zf�Ï6�v�{i���ZlJu:$��I�C��0o
6��lYPX�ǝ9�@�H�Mz���J�V�7����xv�����U}��.���a�ѵ�.
�R��/�b��"�!Q���w�P��޽j�+��&�{;�Ҕ�/����wڢr�%;8���zV�n���Z���+��x-��۾ǧdv������A�֪�+�*�����=ڦtt��F��%Z��Ɩ�N>=|���<�J�C�A�֠�ퟒ��ofm�u���0�}r5�Jgv|¹�t���m��gq���ր�.��<_��a�O�i'�w�dúJ��
����;E�X�)�<^b�A���>����f���)t��&�?qe�n�T>�E��CIv6�#aĮyave��rI�Ū4����*�ꢻ&��VVyu@�ɟ^ؗ�=���V^��9��)��\�;'�F'�g�/�d���QE��vj�����s��%�G)�s�fH&�սaÂu�Y}����0�OZn�i�	ڶ.T/��&x2M��{���l�r�^.&52�/]��+��m��b?�]a\��¤�Ԡ�yæQ�p!�H�+�rr�4�!^C�q�6e�t�Ӿ�|-����5�[�C�O�L������~�}��/c|��G=�S�g�מ��7�c�k���S������T٧�yQ���X�ց�ʹ0�G{q%;�]��rރ��;�
�W��,��=���ʼ�?H�������)pZ�f8��ӂN�\<�9�;�tow�����	7���y��$��n1�=���;�v��F�1�J+���oT>�8�I2���J_����j�\���ur�Ǘx��M��0�^��������6Ԉ��=��g�s:zt�HKwZ{���/�uʻ�Y��u�F�����=t�vU�OF��H0�ڽU
t��}���	UU�����Z��ʬ�vx%80�C�=]�ؒ�7����}Z�ݎ=�$8_���=�7Fw��ޏ|w�uf辝bk;K���7m�:�Z�4�ˈZ�o:
����K�T��!��f�<>Sa���]�Oq�5fP�)�s��l7�D��.�w� �&i<THwy��)�=x����*N�U��hC�9�S V���w��,f^�7�����9]�/k]�]�@@�L�{nm��=6İ�n�#��6&��ﯝu�f����!�ݹu��\2pU��]�knqwS��IBh%ٯ���_q�r���@�\qwC�n��cx�g�]���LV�/��=��J�����b���Z3c&��S V#Ϩk����wve��ulB�o��f:���P:�N=�c2�F3�a��xo��#W�H�zVܭ��9!�t�X���c𨜿[��x�%���>�^5��s�v��Nn�X}k��Ҵ%uت���Z떘:چ¨zD����7�K�)���C6�"��ǨN�=>3�8I�>�z{����!�j�S�
#״�y����v׏rT��xMs����OsfՐ��2k�p9ղ2w��cG���g\̻��w���Jb��^"��7ճ:��^�G�u��KB���y�	8�9�l��[f�������������]��	��L�Z.��@�*oi(8��m����w��NɥLn�m>�'1��bӈ�<�m�c�ٛ����vq���ө�V���	��l4Ьɢu����n�*���P��g`=c��� ��Z���1���R�3���+l��k9a��רT�ʘtZǹ����.�OK���b��}����7�'ruJ��>����K������oU_-EF7ir�n�T�nC�|�
��&S;=sKb�U�H{Z��\��=o��sG>��w��#ڡ6{�e�~�놟�sOHbf*"g�+��s��kO�����}�=�r��lc��3�C���M�yq.;k�8�0�D��%��Wֹ�.�E���x�ؕ�����lS�|[��E��7�R���*�������]��-B���.��I3����� O>x��B���}��M�U��8���;[��j̰�{�;��\�ϵ3e�*|�f+蓀Nv���y�u�h��|�ɬov���t�5���Q��Uۭ�	���>��OՕ��K�Z4�2/=5�gO�[���`�Q�<���f��ӊ("I�w��M�L�O��T���l��o�M�Vɩ��h�y�m�k���ܶx���Z�"2lG˳i۱n�}|D�ۜ������ֺ�`�7V+!�̋�����g�d�##y��q_��f���y�~MC��7x�ߺ�'8/x��g��*
דYՍP]5<üB�)����U�*�{�A�O�S�@!�)��!9J���B��
oqڈnq�b�շ,���<E`	ͼ����x=Bܣ��t򮆵[܄�\j�P�n���\�� ���\w�D���>Ǩ!|4����[^a�c�O�3�����Ίm!&�}��jz�?RL�ˮ>�X#�������V���P��n}�S
f�^��������5ٽ�O.�[9/������yC�#<r\�!����3{~!v��Ŏ{�I�QǪzv�'f/�{I��Q�Z����z���j*j�Ug�E��U.�Jx�1�U\Ld!��{3P�uc�V�����V�X"�:�k@:/��99�)]����X�>SK��[��s��-�'4��ᄫ�eBۓrR�B�5]O'O^�vdW-[ʱ�����=H��#o&)�Y��:��p�w)�Rf�M�(滤�����Y��z̅���˫7H��^G�]Y�E��$^�M�@�5Q��wm:��~�S����^-P�}\!˹W��x#����8�.>��m�Th;��T���_���Fqi
���O}���'���n���wo/Y'{��5�х��i��c�=yP]�Ι4�J��
�8y��(��l2t {H�˷�O=�+�,�]���[gC���]�9���}]�gE�^k���W��<H���y)���X��VgU�':.�Ds�q�ܮ�B�=y������I��f�R����R{G�{�ͭ�}��M<���U���\��T��9�N�#BΦ����+|pٸ�R�A#}�x�
�I�D�Aií��:�([=Տv��2��n<;���[�d���A��[�@9�z��F6H�� ��#1@����Z�L��0A��}�OxC�T����6]r�Jp���������hʦ!�V�zj�1T�4���b��{BTv�a�@�����I���{N-�n��r�TV��6������T����:�a�RoK����t+�7�}tn�&��h�yN8�2�۽�Z�E��u�w�d����qo��N	���.�k
㸠;!Z��op�HFv�D�݅�7i�
B̮R���R�}�ݫgQJšY/]���[�tj��$�>ǫ-Հh܏a�<�V�d2:�p�4qp��ͷ��u���T����5}n�6V�"�@���y)<���MZ��Rj���ͬ����^��k��j�O�
�N
�PR%#|�OQ֨Q����(>V��=��6���Aq̉1�� �Ի���s�>:��o��7�M����"?bs7z�qV���_:/��&���^ث�;&��d�є��;��L[�y��{Bp�:�6U�C��ŵ�?�m�l
%���`x�`��p���2�kaQ�4�G*�K}���p��wW���Z�ְ^��6h��8i.�yw( :#5
v�y��{X��Q��-�k��:ٜ'Zxs6��V��� d�#o� ��P�P)�e���n�tX�4CU�t���83�Q�3���V|��w�k�Ʈ���� b�fQ�%!|�֥��e�2a�Q�b�S�SWF�Ҳ-��ב����z�5&�wM��gu��;��˫e仳�`�:�8ȃ�z'Y�Uk�����S��1�hq�3~瓷.ZÚ
�&bum�w~>�2&GgP���]�=��l���Mnk�4Ծ�ur�9L��g3%���"�k��a�����{q�^��ߑ7���m�8$���'NģJƍ�`kf�N��^��>�щ��éWQ�m/#lس�]��n��]�a�m%�m5�6�4Bj�U���f���U��nﻓ8����͛}�*LūԴ��㗚�� #� 
V��"�4�("�h������+F�R��
h�(����X���4i)�����&��+l[bm�@k0P%USlfhi
j`�Rm�0@5E#CA0�AMD�IAM�#;h��D�%5F�ĕIUTLT�44DQSE: ��IT4�MQE:�4�JSR�Ҕ�,�D#BQ0E�&��U�!C%PD�P�PEQ�U%h-����(��J ��cTSVƊ���%�u�)(�*�JJm��UQ�%`���)h�(�
)(
Z� i)��t�*��
����((b�����t� "��Jb�
("H�h�tij$��$����bi����I)<��y-����
�%l����Ǘ�s�%Ф�OW>wtq�|�԰��s�܂�{��|�K/�s�r$�5K�.s}��J��j��.�&�]���G%׳�h�ޭ35�k1����S����v>���Ju��7���8��2琉�=���Ԅ�s���Z���}��W�ٗ�Nb�w�[�C�p�E�gb��*�+
��{z��'/�U������
~#�[o����(UX�>��V�/-t,�7n��pI�q侯fv���}�L�2+!4�U��7�Z��捤^r5�^sP��k �t�ĵl��O�ͼ��UxȨ���th4��帻z� ��ڽRCރ��8T'!�	e�y��^�L�s��d�������G5s���f�w�n�T닇��5�u;̯��K��7�ki*���{ܒ���n�u�ד��1���gE	����АI3&jK��n���/<�2=EAھ����竨�M�Ծ{�شyw��]���r�+�~�F�d���ֺP����ЎK���ɦ�in��H����9
�<ii�m@�5*�0I�)�иxn�r��"	W>�o�+��������9$1�Yf�H���:�lC{wQ�I��#�s�W������0��]5TgQ*}�m��Գ���]��+�ƥ�����*�4߹����nxn�^�6�ikW��ވ�%QV�_�PkZ���t[��^ȑӮ�f��o5�.��[i��o����T=�T��m��fb���ON�����@d�\5-�}�������O^�N��ad-q.���͡���E�D��գ�����5̑~�|@���m0��Z</��������7�4���<��`�׎�'zh��^�d?M�*�����J�,9�}��V���-�R7�o�z����Ǟ�n^8K7����u`�z|j<���ٺSB�������@�~+�a��S̬��_�c�ޕR&�����
Ͻ����H߭�9"ר��f�W�QN{N��wM\���?m	m%ʬ9Gѭx�<~wt|>��'���޺ �S��EB�;M�y�#��67H��sQ*<lR��%3��G�{<�d�RVn=p�x��Ǽ�yIf�zH
<�%Qɹ�=<r1!>^��3��"H���U�|0�j��^r�0��W{s�ҹ\Z���M���wm�Y�|{qۙ�Sb3�֍�/�:H����k����4}�F��g��$��o�`$d��,ǯNۗʏ�%9���#����5�j���^�=.��C��o�A��=�U�b㚳쌏{�%M�,�ߧn���藯k�9��j��QT}���ǲz��N�ћ^��<�� Lr�_�s�>#�*N֝�:流X5~��:��<���	�e��&���q�U������ �V� P�s���u��`vH>�G�T�E�2�ty	���R�(����b�r�Y�T���7ӝ~�>�{�c[\��O���}~�g�V������7�o�y$v��Vւ�*�ڌ������o�KyM�E-H���[1��H~��)�����5������w��[�ވ^V��ӄ�Ks�����8�Q�~}s����8=3�7�L�^GL�|χD{μ�o���˵q��u�YjO���g��<��S�ue�{x��q�9X�"ܦn2e��ua���z6����uP#-V�~i��b���g����=ޱ윂P�j:7 e�^.��h���w�����z��ٞ�P�$yQ�%@h����b�����!��% �o�2=Rݠp�}�j=#�Ʀv\�=���ʷwѿWj������I��_t[��3ٝ���
Cq���;�(-�!"�b6�E_},�5�B*�G.��pg=�ִk�|-���v�U�4�]t�I�w�ɜ�'>��!'v�w�]�*Y�u^�t�����,��=<r�.r�3m���t���"��l��S��W���CeA�����D�s�>��S�2�P�X���I�H#4�oP��?2m~9�}�<o�G�#
�{r�U��$�8�2  �y�΁&n{v�csէ]�D�;�ѐT�;��TB^�=��W���
�Z���m[����f���I��'4=�W�n��yH��j����|;��4Ʈ���C�׍�_�{�%N �xƩU��ݟt==���ɍ���E\7!U�@'�xׁ�����b�����x�K���c�������X�/�Q�:�{���~]G`׸ٛ�c�E����%��x.�3��n3v��f׸�|L��P�p��>����c���꘽Dޯ0��D{g��~�V�`yF��	(�Ϩ��b���hxvrw�k����LL��rs�s>��������nk�@ϣ�ԣ�̨���Λ��o��Jq��^��n�y����Ԣ����
�q�j��,�����u{�(�z���5Q��۞1~z+������qY�,~�4��}�C0Ζ7��w�}�T�m��lQiW��}����-���V'f<*�5��xW[G��-��S���Əڶ�ή|�_@��~ȏ?����@*����נĞgv6�j�6�̥�,�'�1�ι��|�v�}]��h�X��}PM
�s���l�3K����Sr\Oʼ�z"����q����a�B'���ӅV�'ӆ=�Sg'ӺJʨ��WL\dγq�>	�uHc��~ӟwy߼R��'ǻf{c5��#}�٩��,�ϼ����*��S��ɨ�&+�p��2���e�����TK�_Eh��<�S�>�r�J�^�V�)�,�� K_9��ȣ�Su���C!��AS��N{��W���Ѿ󸮗I�a�{��r=Y�W
��p L�zU �UH�Ή���Mm�;����W���Uա��lǸt�>�H�_{-�<����0��?G���d�Giޭ���R8���t�^9�>
���;t�x���H��˨̸�u�|PP^�g��+���/-␏����͊�LS��9�K�n�>�U~9��`�
��~�XL{�os��,�P�7�*/ԍ�����騿	���մn4��B^5�[�yu�z��`]`گu���W���Pz �� ��*i��
|Y�u�m�/ղt=>�����7z�:��1�Bz��QG͟}ޱP��~vl���<�D��b�	���>�u����m�z��e?׫G�~ Mٚ�[#��V��;Wn�o���O��{o�S�{��k�1NbZt�D�u�.F��#4s����c��k���u{g8�Z�Ys���45���7/���7M6��l�Js̼m���|���|�!���4��ԯN�q��a_��ÊN��PW�|�O�=���.=޻����+p���<ª����$��7�����?ʧ���d�z=!z=/O��8���L	�W��]쁑T�M��~����^�ъk�r�oh�p2wN���!��ڎ��+�|3L��r�㩁0�o����C�AKB�%T�9�t���E:'�P����>6�ߢNaՕP��ѕ����o\����xm�;Gof_���W��֤�t	|�k�7\�e��>��H\=�,�}>�T�b��Wp�&wӃ�9�3�tf=�z�r�ʍϷiu���7��ִ�.�O���F��n�dyp�F�"�sa��������7��a�gM��}��;���|�f=g_�9�c�{NG�/ţ��"]*�؎}e��%�*@Z���r7+Ձ��'5���a�#�\���\d��Ux;�-���矨�~���=E�����R/6�]{��WG�O�U �"�FT����+��}L*����Ͻ�L{��;�k�7%��YRA۟dج�e�٢�
�����2�'�=��� W�Y؂Z>�چ�"븰�ґ1ۗ;�\�odM0����Gr�S�b�o`�4�Z��7=@߶�Џу�H�+��r��8m�W������z���*�ڻ� �������s�]B�9���^� �ea/�vf[���-�)R�g�Q�l���|�fI��y�^G1h��,]�_�eFV�U���������uC}��y�G�� '�t����8KGv?�s�rD�rXr��n�Dfߣ}N��[��߷nE��$o�.���&"����]$'SRc�%f4�7'��kɚ�>�g�.|Ϥ�K�_��[���J�=�t��e@�g̫X�NG�b�s�G{�)�Q�^�]����vLd?z���X�@w@Ty�zK��(]��A2V^�_#޶_�r���+t�>'��N�5Lz�����s�니��	��23�y«��b:�x
�e՟G�����R=�����0�#6����O5�����	;��Dm^x?�Oa��nn�p߾N�H��O��!����X�;ZJ�ە��U](�u�ϫ$�gؘ�J^��j#<��F�۷C��86<��Ϣ}@f���2��a������v��f4}`Uϧ����ns��G��3��\nB��#��H�7S���c+�{tUXN|,��ƴjw��:7�s>S��Bs��f���9�~=�G�w���;���u�6�t���ё�g��i��5��R�(}Y�}2�����@���q��i�}5���-e}@��泥:�|�V��X-��]�����Z��s��m����2�'���q�Ԯ�>1^�w({~��i펑��A����9K��Q�D�-�{�whsvjy+xĮ����;w��ޱ?UU�?\�/��o&|�Ι
���|6;ν��s����Yo������V߈��A�0��E�9'su\�SȁW�L�FL���GS�Ş~��>G���ރTݞ�Y�K&��~�v��������f���D�d	���*ԯY��4j"���:}��(�Ow�tӹ�oL���w���z�-Ue�\ ��P��dz�%�@�d�}���3iflz&���*��
>���G�=N�9��!�o�tT{-�q�W�wd�������L����ER?P�hug��%O�k|����f��������ӜJ9����|6���$
��!S���L���M`��y��e�y�^��i��~>��`1{	z��}�~��>�~�>7w����k��4aɳ���5�&;��G�$GP�g�&��ex���j��ƹ����o+�X~3��P���o+���7�]W}O�*� w�+��5�m�>G�L>���0���{�����|0lr�LM�}�>���gA�(WgşrTY�C<p��<�(���v�8=�7&}�^�|_9���ao����4lMRl!��$��tkw%�e�c^�
VS6Bh����8i������J���ә��]O�?��#�N���f����uωճ.8����7xP���Ⱦ��(>�n�}P�E�]$�$�e�M|L]Ќ�RРi�Ś�bP�oc��yO��}wX=�w,����x׽Tǡؚ�$�����ZN�/c=Z2�	�e<�7G���:$g�9�>�7P��G�3� /'R���ݸ��{l�|zt\D�%�
u�ݶ볫|��v<���iaBp��F�o�V���������
�.��_��*ζ'���&��#���=����ý3�{5��ɝ�r���G��ζ ��J������v��K��v}�̥B�J�2*^��'�,�����ȟN�+"�=����:��ςyR�k��&�4_ko�uݛg�v�o��ye0�W����Ad>�Nn%��"j,	��ü2��X^.��{���g�`���)T��W����9+��_�Å��~
v�=��P���Ȱ2��*��y�uoۻ�;{�y�'=������:H��>+�o��U��2�^i�7�t�~^��Ev�e�G�꧞A�U +���,-ή7���gǳ��ߙg�n�dx�9>~��S�����m��p��Y�
�W�Ð\���gCp�����s��X�j���퓠�4�z�_$�b!�������+5[k���xx�`-��K[�t:-r�f8q�層2g&� 轥Li��uoS�5�i�j�c�U���ood4��y�|B�%5�8��Y�.�*�<�6c�u�&�U8��{g[E:��d���¡ߌO���ۊ�LM>�i���%�T7I���y$z��Վ>�;������~�k@W����Ơ!��@xk�Ǣ�VѸ��{�L<=�QS��oחKs ���d�t=�V�A�<�� +����z�U^��co6�u��;m�}$�"��3�=��;7G��|o��G��l���
⣝V�`�P��]\��D��o�mm�������O�	lOy��n���6P�3ZX�BY�#�Q��ǹEOzg�ܚ+��,�2C��OI3~�>�yK�^���W�k�o�ү'Ei��>j6�����Нw��TG���]NH��<�ǖ-ڽ��ZR��&7�2��Nx���{.#+�X�͚�z���0M2%��j�G@��_��;ͤ��?��W\(~�h�ފ�'�Y��P��emC��u��r��<2��g|�P�|Ls�~�/���{��ޢ�ޭ�xhq˅��K8}<0���,eb��q�;����h�jn'lW_��*V����>��φ�G���s}/�w��4��;�yTZ�}�
Ȫ�|�$�U�Y��eG�5�0n��S�Y470f�ԋ6�TL�) i՜#�u �sܻV��`��-�T�Dn�����m'b�ř�Q��-ʵ%���mCu����_g�"3�=�i� �]hz��I`�sg8��Ȩ*/>��Ye��/�A���ܨ���Ŋ��MF�D�M*�U��{��3PV�L-q��2r��k��M�X�Pް����]�g%�;x��Ӂ��l G�e�/r�*#����Q=,v�Hk"@���vՂ��ӱ�7Q6��n��g�A��i�E%�W{�YՕx~�E�)N�@i��居�Ħ�5�"�q�B�F���E��g�+�3�ڬ�`���t����N{�W#(��F�e��N2���ޤ��90z
�o:��-Kg��WX��ˠ��Ȍ��ģʪ�Uw3ҝ1Ʒ7	D�w��|*�h�em,�^�n�<9�N�����x��u�=�޸�AT�����o���o�.���h=�@c�y� B�5\��89A
���'1@&ݼ�6C�ew=�X�5ϙ��d��(j�؃���r�ןNa�O�2hõ�kyD֘9s����фw3�cd��X;�'u{��G���ltxS�UM�72u��Ԯоdr�D�B��5�n���Wm�qm��\����z胜%�sֶ���1�3FҝC*j���c��!����'
���kR�]�5^ �O��q:�5�W۝wCZ1�x��&<Xv�����Re�%�_C��R$�/�xT��x�����ݚI��o>��F˼;���׃�V�.��J���@w+����j�vr �s�z�w%Z*]�nº�#$#GI���F����V:ٸ+���"��7�\z3���Ӯ��%hu��N��jn�2�ӌ)��E�Mi��Md�2��gQ�{M-�
������s���L8L8-�ί{��nZ�d���S��v$����s���\)
�8�δ�$U���Z�[�`���aa�|�9���A��a��L�$É�$���;�"93���u	]�<�er�7D��	�� ؂g�^��}f��S!p���m6�)	8��N��D	��n���jD�Q�1o	�u�Fij�OZ�8h�:ݟ�T3 �}c����^�Y�=�^I�Y��o�����c}é����;���4E_t	A�����,Ŋ}-��aS�N1d�ƽ���!}���3��yu݂���䏊�6M���nE2@K���J�(ù{KUѥ���Z����ε.Ӯ��B}�[X��	�&��C{V��&]DĂ�N��wL-_J܁��ub��ZM����u��Q[K)>g���.;�G
��M�ՙ3o�7[��Q�Q���[��n�ʰ��`�3�]��g��̣9y�Z�����&ƐL��A��9Q|�Zzp��sYuo�J�tp�'�Y�K8�t�+���Q�����'BB����8�=�c�" 
 ��#DM4��AE-P%3P4�QETELE$@P1V�Ӡ�CM�j�iB����Z���C���lfB�J�������lA�4AM4%��DN�iq[.���PPD�Q@L��LN٤�*Ra��)�j%JZ�AU�u�����J(�II������5JDU4E@��Em���4&!��������Z
B*�
)������D[�ht���5�ӡ*���)tꉩ�Mih���)����
��l�6�R��D�%U:4�Mhu��IAA�Q���N*5��gD�KHDKAAI��
h��E:���2SCZq���$v����J�J(
)

J.����)hJ ���
 
�~��{�Ȼ�u���7{��t��Ci��Y��{Gk�NtЮ��Ju��*�&Y�m���3��R�(�	����o�����Jg����-9ȎsA�u�9�K�h�d�w�ڢ�_��DU��ʎǱ�g�5��<^_���&�x���"����U�t>�����u&��uOb}c0���L�V ��>4a{�S�~�@>Ϫ�eL�@�R�]f�
�z�x?9a���<�e�{t���D�V��7k�/���F�܄1�g�!�ٯ�P����^�gIh�3�j�.��B8��
�>�W��Ĕ��UW���>������N�o�^7Ar�$�n)M �}gIh���؛3������{u*Wp������~�pvx~���n\�Q�+·��TBTFJ>��k<�ٻ��ٗ�yU{���wN��rf���+��>�g�r^P
�������zH��PYޛ�!��[��ͧ�0���W+L�{>������m׍�\G��ǜ윁���>'>�n1^^���&��);D�h�*=����O�I�s��}�ǩ*�,_:�����Z�9�W>���~9��K�@ͩ�}b��,�=�
��K�#�����0�g�{�<�� O+��5y�懪�E.�]�D#��:B�6�z�6�=,�ʕ��K\���ߐ���a�};@���;��%�)��t� �ғyd�=SH�I��q:��=����[4;����bJio���]�Ԕ��h(�w<��6�d;�;)N��;�Gv��;B3[v��!D��OI׮�P��) O��t�ó���q�U����ztQ�&&*i�v�k�#�M =�~�.<�|E���x���ۡ?h��x�D���7��_�[p�f���1�ώ>Iמ���o���΀ش�<z�=�G��Ew���m�<2=[Z
���o����d�E�v9���M#��L�/}!zx�h����O��߬�5��+����v.:�T�U����e򺦉H��{Z
��2�X�u��ɟ"�B���|2=�^g��ey�V�'�iܳ8�g����B�T��{����u8�����"}~���d����g��4<ʕ�D������	gTo����Hx_�p;���P��%���\	n@v�x�ͨh�(����;��o5�[Zx�z29�G��>�}`h����b����Cr��ِG�[����xZ5�W�M��T���ͿC�^5�ƣ�ґGޡǙ���{/ף!̹>�$4nΧ�
*z�6g��*�p�A��>��ә>��w���}9ģ�����r*-�9 �>ښuF{��U�/��$���Nim�6/�T�&Rܭ��w�q ���lW8�+j����fH��E�1��l��W��3�]�j<�=��������<{	}]���<y��Uo$���xrd���[3���J�ʜ `y�){WWHT5ү,��a�>>0|=�Tɚ��:�Ð��z���]T��雗��ڟz��������s��==���@��3��=��W������k�����@��{���j��\ZN:�c�q��QRf�3$�`?]�	צ�=��y70�c+t��OI����W���t�%�Tm�����eg#X<ǻ޻�}�H���Ͻ��Q����Fp{M�n�;����AGG����U�Y���3��/�̶3�Q��'�ǽU��Q�~BJ8} ,'g�k��T�vdiO�{�9)�>�4��L� ��q폛��:T���{��<����L��س���:�&$F���þ����9\2�&�����Zn7�7�qŁ��א+�U���;�W#w�\O��]��^sdA��r\�}�E{�D�FYU�5������r��#ٽLK�����@I�K�(+w�o����Y�ry\�=�-����Q�8�Xߣ&u����O#�G���1��S§����y��gn��^�;�R:�X�K�CF{�)��S��Z��+�N�	��^�U��:|�ېQ=z�ۋ�v�
�F~ռ}F��'e���F�%y]��К�{����Qt��6;5݉.�/��4	�T�������4��=����&rsΈ��=��9MI�/������dO���"_�]&��6蠸�������ѻ<���9��)mo�o?eG�'~��x�ȿ_����l^B��ǻ���(�)��>���2=̕�q���l���=��^F�#}�v9�E�>=�F�_�U��2�^F��G�+wh DW��v^�[3X��UH��]p��dDl��������m�ϼ�]��k�n��u����&�e{���'G�>�n �A��HU2�V.W�fς�����x���m"�{\`Q�eX�7E�_pS�0%�<�"EE��nC1>f��A��T����W�����,z����+�ҋ�{kw�'§ڏ�N�7��<�۸�n|jʠ��}2�__��>�����>�EW�de�g���_���̰��>/��
� +��[��ς�3����!����������W����O�e"����	�o���l��@��{>g(;�K���\kC�=zf�d���zr\��*Ю2w�t�I����TZ[�S�>����f�=�σ�6U��%yfϫ�6��?���C������M��T���4�ްi�?5LU���w�yS�#F�s3ꝩ���J�ٙ�J�-;�'��A�T٫��%Z�,��2�my���EI��K��\�h/��x[;S w]��+#v�P���A�����4:�� ,���6��C������Y=�T$�$c�癝p�3k��I2�ȶ����v+�}������s��.���������Θ� ��!�ڇ���,^l֛�� o���`Jͼd�O����w�R��vw��{Uxh�v��q碻�}>��T�;790�3��u�1�N�Lz���PN$�R��C�~�/ޛ�����{-Z%�h��Ӄ
���V+�{�s�O�p����vʉ�ml�Ǡ?����������?��q�o��~�J=q���eV
�VPR2���V"���j��u��^���]/�4�9״�{��Z;��%Ҩ���Y^�}�b��{��3y����^x�:� �f�ʞ�Z,vL����_�_�T�ю=+O���5C�}u0/��>1]�g�W�q^��B��ag�]�Ҩ�FTL�@��+��m0��Z<<��1���u&Ex\�s+wu���T׽~��ϔ����!�@y�R���Xr	h�3j�#a�=ꙭ�~�T��M���>�@��� ǽ�뱮Y����7� 7�t��A}^��&L�}�������z��zƳQ��p��9����=�����r*�S�/·��G�ߗe�/�,A��]�W9å��P���m8�v{o:�C=8��3��w)��+��-j��,^�n,f��NQ�J�<չ���&�X�$�x:����R^<�}w�:չa�W�U�Q��X��qm��f��GS�;/y����ѷ�z�[���rƬ����'��@-�ӐO��r��Ǽ��G�u�I>�>�%;�$e��tG��)�ݚ�����D�|"���`�����E��"��;���/BVj�^71q�:S�� z�;�>�\z�lT���=�� �9׉�E#���Cܝ��'ä���A���=jh�+�\e?i��(A���Xi���顩�y`���}>G�'��5�
�O@j~�cz�́�?%H���N�J��'���d��u)=q�U	�i O��v�'j�L5�ZL�{T��w�������yO��Ͼ�x>�ǀ&w�(�u1,�{�n���plG����83M��]��"}\d �o=��Q=x��;���7��k���Q��
�Ӭ�����9���qW��m��zd��Y59�4���x6��~�w�S|1�xY:�3�s��|v�������>��*�{�h�a�Q&z�^�}6u%q��kAYV��x���6O���!T�3��3�_n�ʪ*.=��8FF'���Y��W�G��|ag�*���S����2*y*�)��ɖ���a��>ȿg�n� d�50i�!�+z�\�]���#Zf;A^?����{o:�˚8�<%\�4i�еMŻ+/��q��{�ř&��h���`���3�k9��U����x���wes&�)��ܶ뚓1�{wZ��K'�wr����=�}�z��R�������z����MF@���+�׳����f�j��pTm�#��\<R/A����=��x_B���2�'�{7dz��e�9������\�{��ѵF������sސ�g7�:+�n�_��W���Cf��^ڙ��5o����q�ux\�=�������U��KW�7⸔n=�_��F�ځ�r��{fh�m��ˬ����$r����JȦ{� �Xq�T%�C�����c �i�g�{MxX
r����+-�z(��~O2&��JH
��{"n�����bi��:ϴ��Y�Ь��w]#Tq~m����g7ٞJ�>F�����'g�(^7p��i��U�{'*�V�y��5���z8��A��~��K
jO���k�8=�?U���T3� ��+�1%��������ڇ��#ٓ1m9+�l����|ɚچ�By�᜝���1���8'��6k�!%�� �������2u��}��zB��h��N���^=&�V_�=�75� dG)�7�ۊ���ZٿP���_�j�as_�wi�識�aG�S��.�ς�H�(���y����Aěu{ؖ`>�k���e#�w~�J�͏���� ��W0<�U�ʭ�w';� ��a�S��j��DP��v"�;�ǭ*�͏x��wb�7��G�Om%��u�ul���{����ۓ�t�=��*%�����ɭ>���ߵ��M���6�s��ϳ����^G*�u�_�g7���Vxʲwѭ�j1��	�7��F��3�cc&w����:�{s��;l����ձ�}sי��@�+;�YZ;޺Cz#��(���E6O� �c�V+�.2gY��g�7�=�f-v����uvgw�k�p�E����x��χ�}��<6=�P��B�����3}]놭��V�̅P���F[�������sʇc�{N{�x����B�����;E���	i�0Mp�=����~�����TR���G��\��>�٠Ѹ�uC���E�3���������x)��ˍ�~��e���yh���7�R2�Ux
��#�,%�_V�q��1��.7��ە�h��AӺ���{���k�`h(�UH��lYS��:��Њ�g�q�HĮ������4��*\w�P�j��,�r���7n*�1?S���%���zN�3BG��9�7�C���U����`�z����"�׍���A���d���&&�V�v�z��EG���{z�r�Q��W:Y�9�w.�R�p`���8�0A�w��	l��EѰ<�3=
�Y�r����ݫ_ac�:�гۣ�ղ�ĺ��82���4�,S�DZ���L�{��F�P}0�j�Z]����z�6���;��x(���@{�̀C�X��h���.�6�u�8�N[�}H.̞�C�ճ�|�^�T��zU�/O*���q�:��K���.@ߣ�+�]_F:��o�v#�+�;��c��NO���td�3Q��f�K�J�����<}�<��j���kD�v�,��Ģ�����ǏOᝓ�}�D���?���*�ǆ��\��3���F���z/˰��>ɩ�rڱV��:a�a�HGnv���{��p�}qL��7��A�`�ܩu�N��Έ��}h�+��	��Z.<�Wq��:�����y��/i�T�[�93�Ǌ�"���3�ՁV�Y�կ��/]!��˅!p�h���ѥN}E���C��ג��ĵ�n�z3�ϙ�>��o�cn#���s����ˍ��v�G��Q����f>�u�c�!�W^A�ު�&���L�1dϗ�ub�;���}/��Ͻ��7�\n�SI�]^�κ�u
,�^�@R7����*�
<���XY2��O�Q�Z:2Wq�z��ځ�z���&���ۺ�K������p�eE�+�J̭)�D|�)0wz>8e��٫��Ї����=���z�!�+h������;�j��ӥn���.����K���NAE�8�ӛu�3.n2��n�fӾ<�T���ʫ���wج�.�-ɳ��W��$��k�vo�K�g�R2�e�DZ��5�,*����Æ��1/��){8��;��p���w�H/��8�5�CR����U!�*Β��/3�ez�N�&�}�qU��St��:H��R�o��u@{�	ƙsd��fQ�^��T�Ī��r�l���|O#�=���v��q{��ư ����uNH�:>�l�{�Dn�~v�x�uA=�=^��px^�&=������}'%� ��&�Δj�Qjr�s���
>�#�=@s<jX͌�ꋕ�F��;�e���n�������R�9�-Ld{	ܺv��{��C���^���=%ѹ��(��͈��.�'ä�F��ge�o�U�b}����FD��P�/�\\�����OM�M�|YW����|�d�G�U��^�_����h)�����D��#�ӄyW�����_�����W}~�����S�s��t�ó���tM���x��EVy�����4����#�qH+-����FyS�ǻv�\G������Ν���xU}����dX��Q�ү�](��j�zP+��>3Y�ׄ,��CZ�����U��������Դ��l/�7�r�Tv��
��MZc]�7�����+E�F��;z`�=�1���ooa<���������K����˪*�w�2��yH��q�}r\��ըA�'2��/x�I�_?�u��]�r\�ʂ���.��w��i�cU��/V쮭�C	Z���o,�İ�с�@8�&C��g����Hb�nxP^��mH��(.o �`V�M��'ˁ�N�흈93ݴp'�ƨs�9��:ܦ��{7��,�94�][W�m�ڭ����m�̹.��Ԯ��:�[Kt }l^\l��O��G����J��D�/N�~�w�i֫r��1I�Iz��א�W�[ eYZ��j:�j*�zeN�3�2 �*}�v�To
؄ v6m��9(�m�,wUfĴ������fZv�jg�� �&_P�.m�b�����jn��Ճ�&�n�$ۍ�w
�ڇ�
��ջ}��Z/e������s���O(��w=�S�^ʽ����G��N	�͎51�m���_]�}�^W�\�[Ý�ML�ܴ*<�1���#jMٴˡn=�v�[�.���<][UP�5s�\���s4��b^��CFJ���=oI��v�.\��Z̀����d�3�]9�S��,��왊�����2�݇,w.��-����'����n؏g�k��s1�o"V,J�sk�<uE]ʻ��0��e�z����:;H໲�&�5�m"�=�R�(gvz�S>�aƟ3���&�rC7X/fj�X��a����9�|b~/���r��x�3BA��'ڵia��4K�ٔ
G�������ڏ)��/�T��l��j��ۺl'E܍�:�P���̺Nd�ܥ�T�6ӟsaep$�`���h�m4}=�]�0�*S�.zw�����|�U&�hB��͍�y+W���Wz�[K.�D7�V+�T��ʐ9�6j�!�f�2��<I�k���/s����Ca':�۝�+[�|�v�F�0�1Yg�Nj�痷��� ���nJ13t'�v��#�,9=�i򘺟�k��;��q4�^�z<�ћ�C8�2�{�y�ǲ�޼�ŏ��׺o�N�!b �����ϸ�ԑ��(Ӎ�m	q����l�P�p��&��LCw���;�b �WP���82����tg��R���K>���l0�K��h�V�t�Gs�]z��ī�u�3�^��jg;n�A��W����"7�*�	p��Z�&.S���C$��6��c<��]X��U9aZv�q���M]@t���g���q^�o�����ʳA�㌷�%����xf�>���`��T�Д�UUTULDE1&��J4U#li
b(���i�K4MS@�EIAEl�(J���i")����e�JS��ĥ�%450E$I3F�*��KDU�PkM,T,DT��ДU1$BEE%&���bB�
)�
)((�*����"Д�:+AcSHD�QIAAATP�ZLEF��:

i�&(�i*�F����*R��%C�ihb�i�кCBhH������KIT:E�KM1ABPQIM-�Ӫ����MR�h�PRD�MhuBѱ�(��h�ꅡ�Zl1)0�T�CT�I���襭h�M�1,DTitU���߾u����w޺���T�x�[�n��dp���T����_`b�Ձ�����߰�S��+��F9]^<��~�+��oJt�;����Ԯ=y)\�i��>���s�+q;�]�\r6������G����� ���}
71*�d,>�J��^�t����Lk!9�G����7�~+�ǲw���wG���J��DmO]��pc*}	-�G���[9/kAY�U�7=���γ���鐪ϙ�H�=�X���psw�e��Fߵ�vyQ�wE�9'su\D
�L�,w����mU,��T��z3�p�#���J�wH0�Q��P��e���T��	�i���]����q^�9^�B�c�NR*	�]��0?W����(��% ܗ���0}S,a���<r;tz�Э��崙�o'�{����n}Ix�<���:=����^���o�.c�'0Oh�^b6�y.Ȟ>���S"K�q�|Ng�/ƾ��r��x�A9ģq�He�Gz����ױ���H�θ�+މ�7����"f)�x�+p,b^�=鞯Lz@��(����f�]�Hq=�3�S�u�fD�3� )��SW��jv�ƹ��Ő$J˘�Nb���M�,a�O�H-���%�V�{V��~�L��+ʧ�x�ek��B�V��h�m9}c��C;���ĺ-�!��z��û���D����T-�Ymb�{.���N�rü���''Gu�KJ�9��(�c�)�2j"�wru���ٗ U�- ��e<tF�Y��S��ֿ����>~�7�$X�ڀ�zmf|��NT=���0���}���ލ5�u~�%^P�[ב�rv�Hh�v+��9���t�s"�z������d��3'���L{�9��~��񿸾&kj�'�~�O�_{�	���V�E���Q��9�w�=1���<���D��e�ثB�����Ƕd�v/\{����z��ǻv�{)׏d��Μ��;S�l���)$�'�PÒ��MiW>��\���`b�p���x�X�U�o�O��v�w2|�����o��_���O�aՑT�VMib�g|o\���G��^���ɕ{���Y^���$}�\�^����F.��}>��V}U�Q��'Y����(�#'�ﴥ�V����#î<�~ӛ�^g�s���p�>pxr����rf(���K�w~��GX�����w��ɖ9�*��������=�xZ�����	w�1���D8���}�י	f����G ��"����6h4{�0�\����9�|}5����+�=�)���h���EVCj�q}����lY�l�j�-h��cN.�r����Kxc���Ev���w�..�;D��� #W<9�=�k��/��~�{�է����-��bSQ���5��(��M�eޅCw���� �bC���5�LQ��-w�-b�>4{�d��] �*�eK�\��}�,*�ξ���:�9�;���C�4-�-�;��������|ѿ��UHU+�a�_l�*����>��'�s՚�ʩ�^�oi�9��5���ȑ_[�n�2��U"bb�W��-��_���b4U�[3kR�*�������؟:�7�,~>��z��p*!Hnv�dƯ�c�lo��/�]AN�s�>�y�����P�5�q�*����Y� ǽ���H��mƜ�8^)�ٝ����Ha��j�V�d�o�/M}��C���8_� O�X���ڼ����zs��=�6�T=�v�n��rX����#'|f�X�3��l%����uG��<\�!t���
�06��z*��n�¹4}�������=_��d�\d�7�;,���#�V�3�uTY�_v��Wj�'v�N{�V*��+�/]ċg6v���{��p�|=o^V=��ʗ�\��C�/�]l�*����/��V���Ew�!����][�^����Ư��:.1�4��.�ū��M�ɑ0�lĻ2 W3�r��s`����� ��R��
��_Ys�OwB�
��/��
j}��`��޸Dܨw'O�k�d��hyjZz:��ծ(��;x���6s�-!Ɠ�>j@�\�o9�����?V����y+c7�����ҧW��=�df3���<g�܌~W��M����	���cm�_����~/�u����|2<��)N�����ě̝[�}~ʿ�:l {�EU�7޸w�)�a>^�惱�߸�x��=�����rLM{7S�4���2��X�J�\Up�O"*.|��(z�Ux;�2��-�z��?W�W��\�Ze��R��O��Ȅv�1�❛���UHʙl�Q�x�ͦ�%08���V����xx��}����y�l�;����ǆB��zmq=C�)�8��u줙~[����wt�ө6�������ԑϟ��/}@h��[��W����#�@<��9^���3T�g�w�yAͮ�3��c�5��w����\
�{��dnV
��T�퍌*�LR�?]ޡi\�3���3�s�w~;�#�^�]�Q�uW��\珤䬠�0�1����+�};co�� }��H���w&��n3�G��ZdV��ρc*�p�񹍉�rV���ۗ��տE²]��jx�n3�\�8	�L�髙v���ݶ��=].`E��|/y��fz��t������T�f�o����s����p��!*�s��/OY� ��^.[D��^��f�u�+=+���AwDQa`<���Gwa�D���g�E��7Q�Ű�Ms�}�_[(Y�d9#���7�����������ITs��=�9P��K����5�t�c��ӓ����Q>�ż_���%�B�qq�#\ߜ֟d�A@d������m�en�w��8���O
�v��z�EQv�x1�~�29�q�'�=�"���@�7�����<3����:�WM.Ј����o���z{ǧ��5f���w�{����ڲ�\?h�y'�����t{��i�W(�g<G�9<2��ێ��|�oO��M����`TZu�=[��q��G�+��m�=�'�W�l�J꺷����d����h���'S>fp��L�/��!9��#�m{<���~-U^�1�r:qK�M��|�z��*(�C�d�r^ւ�����,nL�7�>E�L�����@��W��^��G������m���v�3}��>�ES6�q�9U�LT� TE�S=}�i�����b⢂����X�}���/{4P���}�>Go���Y��-���^�j=#�4\��ME��v�oɊ$����t����c��t�Y�F����'I�����P*!��~
v�/#L���˨�=�q���p���O4�������῰w����/j���;�%��d~�[�����tS�l��ݼ�4�p�z����������IVw|�vo)Ȼa���4w:��kP}���<�u�t<���k�w�,�+Y.�J�G�_.j��9�E�"W_���h�va����p�{#���_���{3�a[���/�z|o;�}��r<�@RC�x���2&�q��ә��k��w/��#���s��¯���݌�0��u�Ė�ԏE���@n�Q
n�1N{�FJӹ��%�Cѱ4/�7�Ȏ��w��h��1�>�~�؟O ���3^�\���_�u�+���U�o\�w<�#S�LT�w�d)�B����,���P���W�|�yN}.p\G��	5��H���;�9P����0�j[�T7}u�/R7+�'�3�]^u���	b��?H���v7�O���RQW>��7�(H46�̌�J�����7��3�w�^�q��L���N�:��/��R�ޙ��(��~u��b���ܞ�nS+�Q�J����������ǺfX�������Rɍ�t�<L>�|�q^��:}�L�ZTNJq;Le�MiX|'23ң�j��3�]q�h`c����
��s���F�خ&�}�<c������0�ʦ2�kKN�� c�=�}p-z=N� Իβlf`u���pdՆ�'ph�9��MV
jgS��rӄ�D�)�pq|�d6՞��xj��{r�Pac�ut֡��l 9m[|�{Wr�4sc��N#r�-��5�WdU8�Y�������,� ���5����(Hw-�ޅ��vx���N����hvG{nQ���)��>��VET{*�.��ҳjo4�3�޿:}��v/;>�&P~ϣ�Cpׯ�r#|����+�\��4d{�)�&YR�si|�dF����9m.g����.�L�L��s�T8�>��=���d�.*b�S�Y���|���R\V]x�}�LӑG �~�s���l�h�w���)��|{�k�q�Z^�a�#�\�*����^�+�W��}q�@lߥP�H��L
��<��e�Wա����0�<�ꦌ��eyfⰺ@�L�Ft��v�%���[7
o�
�W�Å���>�v�T����ܧ��R�~�~�'��ǼQr�=#J�n\H��S7#�'��(=��LM>�i��Tmy@�����T3�~�9ށ:=Qԑ��R����`��_ �ۙ+�u�p.%E4x��u��~�G����g���<��7��ݟ	�aK�5��_�}��=j�S�X�� =��
�o*������Xo�ph��!����5����o��Q��C��4{����r%�`��O2��xeMFY��I9&�.}�M�Y[[-�`�]7�SX���n_Y�v�xl�<w}�nw{�Î��$K�R]�sYЇY�ȴLr+�e��#�����TBH��J�X'����A�﷡�����$��I#S��ޝg����Y���^'ن��>�����6�;�����4��c�]�7����^ms��y�w]��}���g�ު�7�F��K/	�x匿����>����5��ge�Y�plSW��R
������=ކ=�z�d�*}�4+a�nt�ǐ�n'�ӳ�}���f�i��ڮ��k����rѿW����d�����agU߆��ߤ2ו�`��;�+�1�y9��ђ��l�-��Uo1J}�W�޹]�uH���9�i�{���G/�{-Z%�oG�E\2g��4-�~�Px�&^��pg�G�g]ü��8=2�:e�����;�~>���1��c�}�MS�V!�������T�w��ȿd��W�W?_z��ѓ)�\}�>^��4�]{O�_�����W�f�9u�K��Y�G쇍<�{�����@S6����jygȱd����X����oj*bR��c�^zpz9��H���ĿTyI�,��q.�z] �UH�[ R+��k�0o���ǻ|^����ks�ڤ=�%#��=��ã����i����̐���b:"wj/q?\�]	P��A�r�+�D+S�� j]>�c2�2��ʚrt�V����֫�Ŝ �����n퓻�5n�h�Xp�yӾ}b\��|��-/[y�KUd2�u���vM��,�pb�}�f%eIC��w�70���qy6;����/3���,9��=�y���_�O�C�2<����x�)��l�܏)=���-s﫦�}>��K�a��ݾ�v��8}���z� �{,��0H�Sـk�y���V��rG�z�0|2�j���=�p�r ���/�g�U^7���]�}��Mc�(�����������2E���t�^z��\�2+\�`,e%f�n3}B�L�.L��w�=1��yNO� z��
���G&���NT=��+t����:΃-r�*�.*w���X����Urt[�쌈�zk�h?`yd�VO��%�ی��Dv�*�T�[�����Zvϣ=(���y_��"9�{�I��ު��BO��PGPkT�9��7}t��pq���Tz�6�N���L0�݁p���F}�v�#�ܩ�!Z}�r�Չ�+��3U��s�'����%R�V�En�nV��ۂ�kʢ>�x��&�ͱ�.��''g�_!>�w�^�{r���Dw�mh+*�ʌ����ɝ�Ʋ�{z�k����t�Q����g}����6+8�ɢ^�Q3]��~�Lk}���J-���+�h�t���nrR��n����Y���Yz�.J�uc��uyax�c=<o��4�rr�N�.�����Mz��C!F�3:����z�qϯF�Z��� �b���b����^Q��F���-��^ւ��b.{ŋ���o&|���3/[�5�g:�%H���C��>gr/��7+���Y��f���.r� �Ȁ_z��$���TER͟9��zt�t'��Ճ����ޯ�wh1��C�����d2�{�}S����G�/���8�T����mCF�s�p�9l�����:��_�������]����X"�=�ބ����fP�>�22�W�y-n�4U�T;�^��D{�L�}���N�7�<%�3/6+|�J���D��L�ٿ�gd�As�>���}/Ƣ/��ܶ��G��i�+1��i����m�p;'��,��3�VG�&)�9 \y�����R&i�x��>��rc.-Ώyh���z����2�L{Ӵ�3�O�`+~ˉ�g�@�BZ=�M�=���11MV��<�qQ�쌭5����x��z'�z=�r|/��R�b�s�t_�7p=��W����z��WT#�9���׍���3��6�I�F�iu}^*>�b��uG���t�AuC<s��1%߾�?d�~z��d�guelFgc0 �<�ɗ�Myq���;4wn�6v�����۔�����A=��ϣ�p�3���4�e�z��̆g.���Q;pd1��,�TÑ���(Ɂ��>�}�NmR�w�a$
]����lU� (���1�f����D]//�=�ޤ��T�}��-�7�^7�s�X��&캗Dj�cgC�rbE�;�*�y��$Q���Ks�;��ޖȋ����}�����O,�����v�����89�|+,쫵��l�ӿ���G̖%�.X�mbp^���B�#���#P��.W��'��N��lј�5֖�l�K��Ұ�G�3�P�νLo�t❿Q����	8�{�&���uR�I7f�V�7���xN/��H�[*�ފ��rإ�XU�b���B�5����g���AUǓ�=������n��0[Y�h;HU�I�n�������q�u֥@+�WtwԜ7r�������:$�W8��ˊ��6��F^�cMlkb�}��6pҟ==�N�|�5'b]��Z3��1��:7}Z�
!����Q�0b�������b���`�p���n�j�ޖ�i�Y}����]�\O;(�׼�q�%�Gh��܇9"fl�Q�3�J�Pu�a�S�庖�-�V�����B,���Щ�þR� f���ao,r��7x��m��K��޳�>M�mO4��������y�t\�ڕ������)�j Z��K���`<�i<4+*�NJ�fڢ�W�>}BpVA6�I�1��ŽI�2�|%+u�A�0��~���
��@xo��d��r�,��5�:z������Lu����k)����p���7�5������8����=�T�ݛ�������
���5j��+��T���8#FƽYí/\Ȑ8Iﻮ�H=�=�䵯cEp�|��5O=lTc!A��v:�@����s��t`}؞�����>ll���2����̴M�D�z��� [�G��U�+�:�!��/:�0�A��'`y�SĊ9�n�Z���S��5WGђE�[s�\��#b�N��s������}�`hY�V�� 9t�g(Νi���G�jT�=��p��\�ґͷze�:j�慊�x�G{�{WKbhGrt�j��z��@e�7�l.��]�s��4��G�!W[
>��D;Y�ɥ��<{$�w�b[=�ޡ��rS�`�<[>�=�����[���	�`åXW��E[��bٍ�b�5t5�4`R�!+�Byo��hTr�;�9�UvSj���Qe#j������Ε����89Crk����NS�^�W����.��&�w�+��mG���WN�x!�Q��N�=n�0=rl�Ix^^�5��J�ޖ��u\ȁ�鲶����մ�)��-p���ר�]��\"��0�����3�����x9.Vw%RėQ���t�@Pt�HDPPP�Sm�
j����!��
h"
J��"(Jh���i4�U�T�UE)KB�D�V��cM!IQ%P4PTC�I R���1�HRP�Fɥ
b
�(Zi)*���i
5��h��j���i���t��(�B!�4Z�()hX*����-.-�R5\�)G&�CM#h��0DE�"QF�!��P&��RP�CD@ R�TG-:]4���E4��4]�s��y�l���ЄJ=M"	�X:�oA:Q6ZW�W@X��ƴ\���.���mvӕ}:��b��7Nn����[�����n�߬5��i�ɏtf��q�5�Ƣ����O�ã�uZ+�ܸ���R��0)�*��r��܉��t�^ǧ���������Y^���5� Jؾ�+{U��=�e�<qI�Mrl֟ߙ��&;5��:�Ǿ�if���>��\���`g����\��3۱�N���)@���s7�Tm��ݒ�d<�n}#
YT�a�,o�d���OXQ�s9YA�X�gb�i`U�#�#�y�`
�J������u��hvG{nQ��%�|s	���k\uD��S����e���9�3dς}$1�ׯ�w�|��eH�{�lp�O�ũT�#e���F�N����H��X�}>��@LV�Ǯ0�f�&X^9�*�9״���\�����K�l{�{ޤp��Ҍ����Fb��p�P^��
w�`>��8�7p*���ȍ����*��F�I�\B����}���V����g�Ͼ��;(zni� ��K�Ϫ�eK��<���,+���l�Tq��w3c�����Ӫ�j1�¤�}�����[�y��,���T�J�VC+��릣J�����e���5&~49��w����윙���Ѷ�>#����n�J%���Gc���bA\o�'T�N�A)c������U��Cl�u"fr�nE2�qv	�\G����q!f@sK��d=��}��uq.&:��**	��eFOH3�ܩ_j��+н^>T�a�e7������ض�B��b|������T��X1H�}��'}���o��7��|KGw K����G�U���R�z���Ơ)T�̊7�Z�V�޿ ���LMyVѿ�O�{�ó���x_�����v��� *����;�\�/w}����X/�z@ٖ�>3��sd����5����+����y�F�#�w��z����Tרw�������Xn������kC͟	��cLΆ=�%����y��UQ�ʼش���%�{���6��|=�.rϿ���匿���'t����Zu���B����#66�ΑI.�O9� =�~����p.=����mX��{nt��y=���sbv���W������b�7�ruB�I�>��}}H	YV����DyV��v_�v	��y��O�a�a�BI���ʾ�.5�=0������@�t���t��S��U���뽗����HcMޯf��$c|Q�J�T���w�2g}7��<K���>�����{.7����!C3�p򋞻]c��L��.of�S5�Kk1����.)�uwq�97'�`قu�o��4|GV�j��L��Qjկ�4&�y�N���xb�o�CU�v-��{��3i���t�\��1A���˕}�L�J����g.�ed��k��GN���̇��u��������ü�Nb�g����j8�q�詜����o�ٙ��r�x3Z|�>D�1���/>�uL�:t��&��>E�%!K�t�>����'W%S~�G����s�z}ĺ�G���v}�)ٸ���UH��e��͔S���e�ۦ�'����S���ǣ�t��}»�o��F߫�tf�� �x��qT�V�=�r�^פ,h1�T��̻_mCU]ŋ�^�����y�������p条�='��z�]���y>��У>%���a��rJ��:W�7�<
�zo@21��d��8���j�v� cuď}�,Q����TD�9�;���%�K£����^t����{���T�A���>���_��Xn��ARGz&鍸�Q����EF����ԏ1�-yl�p��j�:\}�S71�~�	RÁ��{�`9>������9P��oC���Oz����§�23w�;޹�>�g��Ty��c��Tt{΄����wD��	Xn}>G�'�=�m0���{�bv2��{��pMw�n-�SXk%�������_L��c���T�����¶�f�VF�3�Ts\ ڎ(��]ڦ���ؽL�G�Ŧ�p�o\�c"��{��}(�4���oQ���5�ƖըDt��uj��g!O������O5���_�}Ψ���;tVG�T$>��㲫���//-��Y�5���x~�;�ض� WM�)�~�=�I��� YN�Ľ]�2<��GݙT
�̥~��'ݹv���l�P�r�>=�>�3LX�.U�����a��JZ�P�[��N��ծn�x��<��&���ýG��"����O�p2ů�kK�ɝ��된�#���g#�9��ob�z{��~@�J��}��o��;��(�{:Kd��uU�7=���γ��p8�|���7�%\����6|7�|��������q��{�<a_���r$�.n*�	��=��,UM5��B�=��轞F�ɖΧ�������p�#��xquH1�t;���z����',6�˝� -z"j.�*�^.��Pѫ��;��$_3>�uh�Q�����߯+�����X��4{�d'7��r�����d�}��mCF���ïZG=��L��WU��nk�������#�=���и�z��^i�"g6�D�>��XZs6_��L2�{}]��Ixlp�ý���fދ/S���n�[��A��O�0r��v�;�-%�
��%�q�x�����*�p�ү0�p��%o�.�9G�GI�5[ʚ������Q�b����g���l���B?b��ϣՆQwh��֥�I�tp��gM����):���Թ�^�|T�%��>�۬n�����6`���3N{�FJӱ4��L�z(\�d޵ޥWg�Ǔ�ޞ�L\9���s���	��&)ω|�KGr&����~��O�{��I������O9Fv���}��C� JQʬ�o�~8|�yN}.p_�7py獠Lϑ�1����G_��B��5pG9��oާ����N��ճ�G-�ld'T|o�@�����9e �_��`Yqy�.����۳��k�=^�3�鿳v��f׸�q|L�mC��/�#�Q��Bx��;� �x߭�%Q�P��l��Q��¢vXˈ��uyU�����%f�=��{�c�Pb�.`u�Ϲ�=���Q�YQ��Qñ�$��O�Pۉ�c/�Ү2|+N�3ҕ?G[�h�Qr�ڍ-� ;�{ T_��}��o���o������]�>�Hë>�c*2kK�I
z�m�?j��N����{H�HY{H��J����O�h{��aC�)����%;��RM�o��d�ҳ���h�)�}��y3�72�}$1�z��|����W���v����R
���Y��S�z�JރD���T�;/J�Wq�]3Y�{]��|��s=���i�ԮL|��5������9Jɵf��<+��Fa�Ep�=��T��f&nT1LA27x�p�4����\	�1�U�ٛ�n��UL�/��7k���gG����IL7��?�N?��N�"j,	��ü2���ax�$�⯩ߴ��+��E�����I���>���=\��E{�V�� �g�jdX��~��͚�uC��#��Y�#jh�z߳��u���F����7�_�7%��L���rފ�R�W,yf�	k�.�^9C=�ڹo�����iX�3�#��{!��'�`-����T�Q+�ao���B�o��l�8]G�e�!�U�p��.��{%/�����"��L�,��"<���L39�\.f֝�=
Z&<��<�w"��Ct������]l�5�;�"~�zɸ!Q}��b�ؿmS+4�4|��1��И�}[F���%�^���>t�s`�xQ�6����2�և�M� }��@�U �����!�_�d֗��s�Ҥo�~�f�;�+��'6e�35��ʫ�y@T>�K�����D��m�ևy;�:^�'UO������j+�����YW���z��QS�QS��ު���<�f��K/NO��������m�mh��N���_��;_���L��� ӸjR��ێ�f*@+��]��!�K�L��^F�u`v��G�i�9[�Vjva�7!���+JŔd�ʬv��fG^��͌3����. 3j�P
���艥e�s�Y��kL�$�gR�bc�u/��j������>�^k�=�ƹ�\�u)sq�ڱW�s�/����q;0�]�G^�#ݻжk�C<���˦�� b��`Jʶ@����3ʴuǻ/��V��=�n��l�b8d�P�7�]ϫ���1�}�����n7����G��:���U��Q�v���[�QWu�.j�;���1d{�9mx�paS�|2�]øɝ��a���ls��N���
S��L�;{U9��{�d��r�|2<��+"P��]``���T�ҽ-.�V�>�n�ɏ�,�������e�R���-����R��UsVYY�)�܀�f���E\�����|�g6�P�;��H�n�^�����w�q.�Q��SA�����zU �"�F_��Y�"��-��7�[C<Qϧx�ͯQ~�~t��������~���9�p���!�軣�Mm]Y�>����~�[���~p1��F��]^Ä�}��R�H���M��zP.��X=����P���/��7kQ���]}ސ O&Q�Ϭ�%���	��_.���* �k�\��v`��Z���r|N܊��n��b���q���p��3�A��$�yM�6IAY6:�"�f㏨�
˾38�}u� �?nܱ�ĳJW��w�q�Րk��Z����ׯh��-��yi�:^}�pS�h��C+`�t�sŕ�Q�����Tou^X�q�=@�o.EE���E�t<X</�)�Ӛ��8K�_%�7X,B�D�
�y}�y���k���Fd�yH
��,u>��5,c�=Dz�V��wǢtx?0��츹���E�&Z�1��51���),�pw@�:��ß�EU�k�cC�MU0���y�V{xzEO��>��@�mpT�\�t=p�΂S�<ՐD�+ϧ��gt��C�ϝll��i�t�z%9Xa{����O5�� Oܯ��s�>"��R���ȑ��i\|{�>��B�Ѿ}�꬛~<��~ُ(ͪ�i~=7z��m��zw�_��~�֫J��ٗq[>���L�'}���o_�d�:\�h�N���
�=E}X���Y���lx�|��ګ��wM+���W����޸�o��qW�nx�C{Dw�mh*e�ܚ��2g}1q�Br}~�j��={��%�wѮ}h���ŜF����l.��Cͧ%��;8
���&�X����ј�/u�V	�Ot�u�d(������y�߯��n%����ό,�ES6�q�/9_�2�X7~�B	��1�tÉmk�-���
Ѥ7vcXw���{�t5�o��̽����Î����������(�/������a9�Ǭ�=�^"��n��ǋ�N�DT5��]WAW5t��v�=��y�`�0@ŋ���ꌾ�ܬř�k�3]����lzo���p��S�Ş~�Hי[��xuˤ��e�p�/��s�r�#�Z�A�Y�/'���K���K�}jW��چ�_����#��O���X��� ||�n��X��ث��)U�-L�_�L���2��NQ����h�%���چ�E�T;u�H��u�O7d�rq�i{ފ�ooף#�>��0�0[;T����0���~.č�س�b���z_�a�S��g��:�ӜJ9�.�ۗ"��uNH��l�A���������w�Ǽ ��m.�����ހtgw���z}0�Js>���
�~̉��z�d�jG�&�m�E��=�55�r��g����1���Tn5K���,er�%�o�~8|�yIf���T�~5��*؝.k�U�E,����"��<�en�y��8S���4W+��Ws�y�Ȧ��sOm]�
�����=�Ig��p{M��C͟i�/��ڇ�I�_�9���dKͅ�u��M�X��G�ʫG�{(ٿ�Q˟PM�챗��������zM�Ł�}�QX���]�m��L�x���=�eT5k�ƥ1Kv���M�q�4!����G�nI��X곮ffk�6�g�^&�4_M���l2�k�"8g��U �I��+
B��Յ����mp�h4e�[0�ev�jЬ�]��츢��A>%u��9��s�u�X<=�n��nTMD{�Ο2I�'�xb����������/�{i���<��#��P2R5�W>��O^@��O}<����{��F�nx�Ǟ��'�Y��T�>R8M#q�r��r=��HStl{�3�o\����{n3��*-*�o��u�>�b��F-�l��=��U1>�ܬ�jT��Oz*���u��L�7�>	��]^�az��;�*���/ca�Yz���$�h�R%O�}8���~��ü2�}nX^9�*�u�9�^-z�_�\T;��7�٘�a�X�ұ[��>=�H�9��Ϩ�M�>NZ����\>�;�M�8k�̉�� ��]߷���;����[������4������$^}�Q,yZ�>�7m\H�#w�!}������/D{ԃ~�6a�I���5~�p��|Kh�����Br{�=C2�n{o�*VM2����L�Dl��/���n׋��ϧI���wW����x��{�.�Zuw22�[�6��ZqU��-��IH�"��딀�r\�W�f�@"����@DE� �����(��`PU���"+�DW� ""�쀈���A�����_�""�耈���"+��"+�_�"+�����@DE��dDW� ""�怈�� ""��1AY&SY!�1� _�RY��=�ݐ?���`�X}^x���QT�DPIP��U*34P��$����TZѪP��H�H�"�U	U%J�U)w�*ӡ��Dk)���L�m� r��+�k[-� 6� �����Z��p���(A�)�k�H�m����s4��2��Л�n`� ��R7c�lҖ�MK�讎�t2h2-�Xi3
k� ��uwL��I8�c2����f�#*�2�(�D�878�J��ղ�*��bj���l��٨�3Z�Qj5*��i��m��XJ�l�dֲm�mmB��ʍQ��m�:mժZlmAB�i6-m��eމA  00�*�  �    O$�T�       ��4i���L=�z&MI�A�T�RO��P�Cd F�hbCLs �	������`���`%=$U4T���y ��[$F��ZR�V-]� ������*�g�$Z���� @ ����@HAUZD��jH�?G���o�!B
�
��/ ��U\Z�@�	T-�������V�����cZ�X����Y��wLU���T�N�e������_䂿j�x*"�G����"(���G�m%�J�+S���l�3Hzj^@�ڷN�\�j�`��s&�/j��%B�P�n�6��(�|�in�Ƶ�b��Efњm�V�6���6�|$�՛G^�b�s�=˺D[�^��[�s(��NƍȠtN�9H�u��;u���H"�j?*��e��ǘNwn�Q�,�$"Gơ97QDl���t��鵥���P���
+ ������Qz�ԳV�l��I��e�;��m޹@��zU��bv���t�۽kq8[L��x�W%����4O��@��w[;"wV�,�A L��l�sj���w�Fn�:�U(Q�q��Kc��ԍfEL��h!�]h���t�t�k$K�jЁAp�li�7��8�%R˂��/�5�&l&ELh���i0�mCe����1,���V�M$�gVa�bZ��W2�kE^�4s��0*�ehN�()ESn��njͺ�9?��}٬ѕ�Y��Jg�X�Y��m5`l+ۼ�bKMGK�VhR�ޑ��۸5۬��kUl ��0�Bڵv�&��)�Ku��aM����%Ow
WHw�Mn���S�:�P�Ϧ�Y�f�يRMa�&�S^]fJ��τ������&��%c4�}yi0�m�e�&��h�̋d�NC:�.Ά�cKv�&1i�i�&=�8Y�v�Lk�-�fTy%���[�yyqӑ�
z+"ޛtb��P'�vO5�9�e퀱�N�w��ɵ���YkS�����{�P䚨��n//[�EY��Y��0-�uWrԡw��f��4��v�K'M�a�ԌqÂ=[3�wh� ��`�+�,�:Ó7u�f-l�k*��ĩ�3�Q��*(5xN�fb��uD�Y��
��4����fU���K�
�5E�B��J,"��c�a�@=�E����b�E%J"�X�M�QE�iYZƅB��^��ӹ�G/A0�V��j����20s\!�R���+%�X��	Ú&��IK����i7��J(��[n���Pd*����#�U*��G!��M�1���R�gz���wd�g룎�5@Ar� r�T��+j�D��e#�aX�دEZ
̣��6��Yo@j����i��$I�Pϱ#,�e���)�m��f#0<xűX*L���2�-*:�;W-\�X�b+�z\�-�ү5ZD��m�b:�	j4Ւ��a����\�V�0D��v�����X��꽫�L�VdZ3B��!.}���*���B&t��[Q"�DQ�R���t�#K/U(2�L1kf `ZХY�c�`�h�8�<����ͱ`�wN3��iҀ�4�X�F)�iaGmV�n|��1��xHX1�
�"�e�E7^"����bGmօi�B l�uzLn�
«MX��C]���ÍT@���(�[�/X.�e��MI͕wv�B��f���fm�
8K�O� �!;�Alml���f3�M�4�MZ�1Q��=�ܗ����� �)b��k+U�ҫ߮�����jT����
����E� V��֌;M��v�T��:Wo��`�Yծň�V#r죏+#`U����I�Ki���/o��2)P�,�є��q�LK��1U��:�Em2�@VU���E쫛Xe�w���qB�4����"v���#K�,͔�Dv�%����I��`R	Y���Ci�LA�իU�kn%n��Ucen8(�1JW�i	&`�kH�p�l�s��r�n5X~��̡X�7����Mޝ�Y�f��g[Iz�y�Z�|g�C����~���q�	�{�J�{�`���,���7���~�7�т��GlÜ�H��Om.��
\�X�Wh�/vA이��1tu��[�厾���ғ�sN�1V>⻷���{����h�� �ofX(w��6Xs4�Z:a��>�ƻ��Mr�GΕ�w�M0)^w����&*���~�|w������v�x!/��(�W�ݻVM�[�y��)OM��H��h�����=�V��C�g���P�.ѵ*�:�ݖjVr�1c̥�����#7���ƹ�%�{��:t�%j��k�k�B(��RYs���z���&[�U�^��k�'[ݮV$��c��G�.�i��;��9�g){�D���T��Z�-���m)�tUo7X��W��\�����Ӂp�(qy˜}��m�8o��z��|
�J�p�wp�%�A·)aC��T鮥�80���GY"u�!�6���\�,u-̙��q�r�SDPѶMe��wjs쩙8��:����]N^#O)m�d�����o�qd��7@T��SY�T�;�q����º�JT�Z]�沷�W7]�@%���b����/3�y+v�pq�(�pv��r��B��n�<��N���(���6�i����V�!���f�P;�{qV�t��(U��ޫ���X,T�{Qp�Ǧ�9(|G��/)ٔ:��z�m��32�*x��W|�kDq_Ù��񯵞�c|�� ��[���)׊1}���_&D/?N�����+�p
{�vR�Pf��+/��#4t�{QP���NG��#{Ώ\�)ɠz/K���4�2��R���˺U`�he���+p(F�%3v˽��Bܢ��u����B�;R�m)��4�٧�)3��C]یe�����=����s����*�T`(�F�Q�ہ��d���O��z�:\B	�f��U1����0꣹s�c_I��:�����IZ�jȺ>�z
y��Y�E����|Ȝ���f_�'P<M�3�Jw̔��9O�ۢ�*�S���ý̈^5O�NB���T�������mf����������ϟ�hq�������ɺ���"/�:]�]��C@�q�S�U]��FG���,I�a�gAk�#���ظhWh�`d;|�XsWbaa|���������JP%��,f<ݧ��<ae��V�Ax�U8���]k4���jjl�o�Q�7VR����;C�����7�%.a���w.������Z��}	��ڕ+5%�1�<��Z�.����#}z[��L�ʳ3*�G�H�u��34�޻��P^Ϋt��	3�Kӽ� �ZO�Ѵ%��z�)'�a4���,�(1�77�O3a��D{�:yL1V����wK$��
yYBR������\���0j��v���q�������Y[Z�S����8�,*�����T�˙^5�Y
Cb�a��Lgpu<i!������N��~B������ ���s3+�7��.������5m�S�Z�E��u=A�B#��Y8 ���M�^�'+�}����WR�e�����.���o�sVf��֒Q�D�kp��6̪ʒ!$i�-u$DX�6�X���fہ�JR�NY�,>.Nu��� b���$�I�"Fn�⒢�u6��L�!B�(��vyov��^'��-���*�]��S��;��^	L�T�
��$t@�֬E�'m���^.��/�*����%c�vf��j���5�B�U��p�;�Y�BV�;�ZB=ܙ]6�7YрC�"�#�{	�qn�)b�v���i�&w�o��O������~!��UUUOhNb�� � >��UTb�|:C���DEU�v��_�d�}�%�;��l��%X�J)�D�58�7�l�����*�ok��ܢ�Tk�2+8U��.�ep-�i��rv���s(�v�1�Ȩ���z����=5*�ث9�[n��:S=�c5�[w[N��U.JK��u�������5�e��kB��U�O&��b��C��tB�֙��ϰ����5�q�'�D 6��J�ⱃ�q��Wb�=1Z��o�{�駕�!L#����S�m�T���D!����8�Q�4
�G��m�j��+�B�R��^��kwe\��K�É�9���V��6;�s�V�7A��1i����b�d�.Nj|���+keի�w$&)y�m)�}�G��xi�T��\�`*һJ�ͣ��=��}���&4q�c�܏ҭ�-�sX��E��Zo(�vR��e�f�3���6s������&]Ny��c΀t�DWYf���ʳ��*Auuգ�i&�:�t�~���(�%lh�t�ڔ�J�Jmr���9��+���-Y��Aj��ݗCr���Yb��x�o���r�}��>\���ݚ���|I���t�j˾K�w���B��+��yAu9�K�ٹ��+�w�D����r;���Nv�C���X�.0TshU8����Ne��	�>?[SV�ۧAݷ	��,�1�e���XV�s�;$��íL'���$�R\�td���ժ�m̕t�TkP��Ә�G���8��p�]��G����R�d@���`��+����<)^�귱��ϝm�Ȍ b�/)J椙nt�.���EwK�y*t�Mp���5V�����Q�<�!��ۙN���g6�,�]��6D�*���\����E$� [�-�"���#���f�q�װ�)_B6�1�U�Ɉ�����X:���8���Kr�n�s�@���nRY�5S[�_Ԟ�m7/k�6��u	��v7�!-��ȻN-��<�ʖkNMgJ9��J�=yAH��6�&WH���h\W��u5qTi;ÒL�i��}
ե_�w;�W���p�w�k-�_��<fPe
}���g�\]�:��'+4�kc��#��7ʪڶdB��]�4���E����/��j��R��t��+�ޱ7b��qg:�+�ٷ�z���nB˧��Hй���؂�:�x�o^�4�����e*��mw�*F�ؠ���j=KG1�F#g�Q��#�.�4�JE��@�����;[��jn|!�-��Y�-yRD�S�����Jm�[�.E��y��AXzu�+s���d(��mq���Ŗ�T-amGub1-�aS��tc{�0�=]_i4�)lu�.�A�wwV�'��M��U�C���ބ`BL�,Mˆ�6\Х��c�`��v_J��q��؎{��L�7��B��h�����{�ፉ�&ҬB��#t�ɒ�����Dr]��i}8O�3��.��b'9 ��Ռc�]��3 b�����Tme��%�,g�!Ü�4����`r�Z��
�G� �S�U���v��^�]-4��Y��T������'�q�O�h�V1�Ȩ��9S��Ԡ3Z��V�e[��-�I*�2X�u�a���3���CTtT�j��.� ��+aia^�1��Ɋ����d���@S��<��͡�Βx�޽CM�X��o�����V���:�@�p���w�8�fm�8�s:�5�lK�;h����}F�tm@e6�YY�@���]�7��v������8۵������+���A��s;��_�-U]u�kl1w`ѱg	y�+=롵,
��=���+I�;����ʠ���A����]W���`~[S舨��#�]�#��@[7b2�Q�'S�ڛ���.��q� (�@�?���W����τ��9㵳:��A�B~����͟@z�rf��(�r��W��]���y��,+���ͮ���=��u���3v+�Pv큰ExiԤ�rm;��{ΰ�����:V�U�#�^\]u���Į��v�Q�B�al(�	�r,ފ}݂3��m�YͮN�V���k
��Lw!*Hz��;<uoY����r�!3.�m�AWwii����*]�YM��e-�1w�8,�L�Y+�Jn�`�n�w�& ��U��d�7airAVX��	M�b�aLb$����0�J�����h �DcT*-$LH]�*�K��ŘI�!��Pnbc��Ie��I!���1�#d�c%�v��"$*w��b��X�
���Gv�K��Ue��c�5���LM���铧<�=â(��r�@^�I/�o��zf��rh� W�
1��UO�[dk'&���Y�b��\��8���{�ȟV�cS��V���	ʨ��P\_S1�>^���^�6Z���/U�sxi�O�n˙��A���[z-jӴB[�VA��*��C��`���O��D�	��hSrd�OU�Ҽ�7�����tK�t&t������=�ʗJ�D�����"�<~`�F���X�r��BI��ۑxrE�:X�)�i����;�n�f79l�>�Eb��=LX���@�p
�)v�@TY2�mfԤ��s���'C~����x��&M_�<�X�x�|I�k�;�Е�(]T���ї��u٫�bފ}�5<�;�'�5��P��Q�nٸ}�Qq�d���·�\��ӱ��*�� ܸ_k�P�zOV���7�λ���f.3��-��`�c��pn���]yo��&��s��2�vXO7`�
>���D	���4#uwPJEc�k"�(�����HLd!J��O28t_�⣍�����8,�Wf�#4�� �?rB�v�6�㗂�x�v����I���=��Wi�:��t�&��T�b�{�`MS̕q��#9f\5~��X~u�?1�����g��o�09^XEw*g�@��MϷ�ל)�.�P9��5��3��ncJ0jz�����*gB ���N����vv�	E����%���Ec�rS��_$J��S��F�Հ>����Ts�d����pM�*��eC�o*ǲ'��{1�<\)5���;���BYݞm��3αl���Fyҗ�(�k�m�<��d
����iS��[���bq���˙IIb�&�X�Q�p‷����hP�}��)DdU����{;ԗ`�=l��ҝ���2�(0�h�)]����Z��*��]�	�T�׻�x��<r]�K�CO�(����D���%׬����
�ɖ,!�7�SwL�*	V�Tve�C�m^> ��6v�4���zwp�ѷV1SJ,���m�5�ne�w7�Q%O�N�ZVX v�U����xٜUY��]�2�@�VkU�)Ȧp3[�M{W��^qm=Wyn��g����WI���e�GF���p�#ᒾ��a�9�y���3�t��T�(-#$gض�S�Z�á$�,�ʈ�c�� �����ӱ�C8e�d�@��pyn�V��,p��.wy-0��gX]���%w�,T/bռ/��ivC���J;�,@� �
���i�sǾ�g:�v��h�g�v�	U.�ʳ@��% RR�>wF���W;L��qP��Y0��c���]��ȝ������s�{`��Qt�q�K,�0�Weq�}�h
F�O{���簰d�ځ�T��P/qiw�.;�jf��J�.����ô���0��}���}��~���V6�mm���7)�C���W��VS�5d��"�J��91��;�vt�f+��������WW�A��׼:�",��CĳDbo	�\=�V��]��2&ҩ�2�`/��7u�n�|��8��}Ğ�9�ݜ�d9/L�E+'kFw'Z�:�4����D�0�jA5[O-���P���~�N�3�,W[�| �۷�Wh,��p^F)�B���)���T��m���d�:��Nڷ�E�"�%\�Q�0�X$:dYAhQV�d�w�n������.��X��XP4&3�f\�`0�iм��X ɨ�TBZ*�1
���B[7"�x(�m��(�FfYi�ŕ�Ck�!���I��z�~F�&��]����E��.B�Y�Åd��w�¸1wm)H*F]ܻKB �i�B -$(�UHPD|�J�H,�MSlčM�F\�V��A��d$�܈4�EDÆ�i���/�nJ0�na��b	$p�h�cڍ�*�T�%cR�Q)L�2g���~;�����2��;���cu��˰Nά�H$n6�7ߔ��7��U��Gr��g�z���̯�j:��3W�R7�Q�,��'8�&���~���1��v<��;i��ب��C����f��1P'ٸ��t�M�>v�7u������`N�U��mߣh���Ս����J&�����5����UġH�ikÜ�Z<�%xl9��Niiu��!�]�p秈�{�j���u��K3k���M�2�xW����WKR�i�G�{O�N:�:Tr��f�t�c&���^��t׸�7@�k�8*K���=�GY���Ԋ)'�^\��p.vmm��D���P$��k�m��(�iM=W�H�ABD����3*�j�6��9��8�4�l{<㓇�'^+-!�X��J��U��:�pv�Xz,�����*֭�LyW~Ke�U~m?������[5V�Ik�����|�7+$�]U˖ep�\�J|ۗ�φ�R^�FLz6b(:�F[������(����WP�y��pj��
�}
�@^eUh�Dj�����ꪔ4Ua �j���G��;r�� u�-
ߍ�_�A���֪IUF���U]h4�i���QƫH���{;�}�U��`��J�)U_4i(8�֨4�D������\}��4�q�¨�Yh��J�4W�m��̠
�U����`q��hQƴ�h�@i����(��)U��i*ƪ�����
�Z�5Tq���y
��8�h�"s�[B�4J��U�g:�>�TF��4Q>�:�U��C����Tu8�ƪ�����Tj� Q��Tj�R�ڪ�4y(2ҁ��סA�DϺ}��ߦ/ӷ~y�������ݦ�P�O�eO��R�%_AK��=�ݯz"&c���
�h��T[X��IA��on���HQiF�UG}
�cAFZ"U�A檫>ǹ���-J%�B��!��*��vUQ��TD���+�\�3���R�GZ
�Yj��Yj���rUa��5Ti��(��c���EU|�GP>h��W���%J5U1�UԢ�(�������ހ�4Q��:���Em
4�e:�UD��UG�Q��|���q�(�@-���Ji��-����@4�O�Tc�w���{�W���9�A_%a*�-R�G�45^h�U5F�4W�}���׺�;3tQ�
�TC� �1�{s�ײb�����k�_6?r߈��w�M�/̿K�5�MNKܭq����O%qj3Q��`�� Hq����+��Fk2;�|�Td��:�Q����"�*�\�"ˑJ�T��Gj9g`״�Q�u4�&z��`ДG;��f����sp4�Ъ���H��譃���ә5U��f����gZm�"���Hxq(�'r�7`$�B*�Z��R��8(���P���Q~m��
�t�Z[�ӷ�����oÒxfL�羉V�E��b�X*�7��ds����lti7�����^�׭ۨ>���E����o����Nf+X�-{f'��xJ/�O�nC�x>��U1C*4V�iY����0���*��[�m��r_)��z����H�����ӥ����#�������/t��m�v�Ƞ���"����1���^xm�j�KE�&X�C�<�f��� �ڂ۝�X���n�s�L��(L�i�OVу�Q�����ca�2�T�
0�i���zo�6�#��6eF)��;��:�.�ـCp���5��\<�V�g��[�1N;XiST�ݛ�r�+k��{��0�V�F.�E���[��h��v�{�m��;���`����<v��ǑKF�h�'�Q�w9rm*����_���E�O�\*������q���kDa�E�����7��j����^<�U�X��˨�C�D>�}�נ�D/��q�;yW����÷����gsxa|��{jXf�=n��-��	�þ�?x�����YJj���7� y������T�-AE�8(5�wu���/����M�4(-㴄��`O��S�-V���s6�vk�=��L��]�A �(�:_9s~�{uB�L���u�]_%� �w�5M�Y��ʋ������h[FQ��P�10�U��S���BG���쓃���
_ZK��񝵴)`�˺�����RõHFG&$���*!~��ob@~](����`�d��Wl�SWw�2�Ѭ ]ZB�%݌�Х+�*;ʻ0�eXr�\�T�%J¼����ڵ
��I�j�pQ.T�u�`�9x%wDE��i��CF��t����%��B� ѓT�C� f��2��@c���A��f�V��Q���$�In�]k�������uo߃߭w�J~���0�#r�ƣKW"� Ԃ�F�hZ�T[d�Y�ԶR�EQ0BU�QX�V� ���"�ґ\B��"4Ҥ��)BH������*��,Hԕd��(\"��"�$UPH�XA�F1j0d-(դ;����!�xB���AZ��D{��Ci��v4���#���bw2����{�'.��wo��o�� 3K=���t���Uh�Kg!���	'$f�l��7�ֺ�/�K�K�Id���X o6����0$�;9��[dm�j�]�Ou���r��Re�7]��
.)o��U�W)
ہ����Dz=	
u$�샽��٘��N�&(~�v�m#R���q�Վt=�F�r'A���f(Z���X$c��������R�Z��I�S��q��[��0�+82�(�]�_a��t�X��ME���D�аn��@RE>������_���v����FqK����-��+�܌y�=��Н��;��^���f�ExSB
�V4��5q��b:�pI7�X������ݜP��Xo+��N�7P�y�m�S�����=U�)b|T>�GSE��s��mȎO%OJ���ɖ�*�J9"�]׽\:��D�pr/��G�9���S�k`��UOԹ�fX��D��q���ڕ�V�9�n��<�f��#���pq�7��k �Kmv�y��ǖ��
�mC�$�ڟ�`�i7u�&��	됏1\��/vR�X#�P�����\���u�dJ�׃Z�ez�dL�g.�M-�8I+��UI �ވ�G�)���k�鹮�B���}��@X��!�����CD�F�S�a�����v�\0���IW�c�L*�=�V
�W�w:��ޫOM�:U�x��umB�S��h������1��y�̋�:{S����ng��P�9ǡA[#'���f�:
�ޏG�M��v\L˱�]��>X3�KsB��ݷ���2��homNdު��(,35&$��A��u��m]U�@�h�l Lrx��U�[,¤Z��^��+l壖��G;TyZJ�jGH�$R�T~�'~SR
6/�d��;�}�
����t��p��÷��ߩX&�8Rq��i��r��i�;k*j���5�7�b2p�v��f[e:��+F�3=U�{p�x���2yfͭǦf?#}	�\Qsڕص���v1�w�+�~'�Q�d�N����]�o4��}R�ݬ���|-u$s��҅�J[����y�����UD�����kM��o�Ώ>��5��̓ΰf�U��q{*_���h�X>ֽّ��e�\��՚$A^�y��2V��x� >M^���[�9�|s&*x�������M�3O��?:����z���g@�5o�0z�D8�?�着��/�{�������п ���G�&�Y௳��{��U!��I"�~��.zڂǕnp��jz��=�KMs������k*��"��Y�_I�mt�oyo�9�����#3 A���8&b��FGu�䏹�՜6�\�;�rȰ�)(��z=";�1����ڋ����=Ѳ�0�ZWzS׼@���6Eg���۵;��S��?�U�Y���0����D����.5{�N� ��&3����z>��\�2k�YΟ4p�U�m��V�ʏ�&D%F>��@���^�X�@��Ag���FDY��|����m7r^loR�ky��98�ճS�p�R�+��%�4Av� �n�4�H�����=D �	��W�cB��%ż57���*7�p�f��7 x���
��Ƿ��n#���nU�����a�]6�r���Գ�
�i���o5@IՌ�l����[A�Q6Z}��G��'w�l�YB��W���Rf�[U��X����tZt1'V�ո�V[7�Y��f��X����\D�d7���>� XQwBSr�|�F����V�C�z
���l�S"k.�AWL*aV;�����]Yre�J�̦�ǐ��Jeڗ���I� �2ȄF�#$e1R21bEcXB��%(���c �"��dE!d)EX2Ja%H�H� ��1I"�T��ҭF����`"�RTRJ��$cRJDbJbH�vAj�X+�H�����?��eDm�#�I�ҿ�����(��ؐ)�k��qJ2���F��[}I��w=F(wb 8WYT��y����[�~ϣn����j׹��ݥ��r���r0z�5=tkwW�M�I���7�Z�Ր����l���g���UDQ7�oje�+�:&9�V��p� ����vW<�cq�f����l��5i�5�Y�j�z9�(q���GeuJ�c�u�5�ֹ����iq9�3�Ew��s[�s�2㙺�ך��Y.�p�8顸a�����O{&���a�
��\+F��}��v�xp�64��y0�8�n��a��ۆs�i+Ha%��ܚ��9�f�)�j�]��+���suj?X�t~6k;�݆�0���Zo0ýC��+��ۅa�q9�^}�PM�t���U�
�.��+�<>T>�U��5�y��.eCu�iX�3�����U/1k�+{>��{���=�(a�t��^l������&��޴t�6�x�z�syξ��\�r�ە�<K�LE8�#�cy���;9p񨉩m��x�'<n��]��L�W���7{��֋�iv#�5�ʞ͙�vh��Ƭh�+�LUk4���K���]m�p�YL���_A�W���Z��[�u܇�5�M���K=�g;�f��&�84X�>ً�0Q
�@�����=�gͽ~75��޵�.�g_P� lݨ�XG��舏���\�Ҧ2'����	�,c����L�ha�'1�L��#��J�ڿnYf����[}����#d!�QPU!Jd�ًX4�C��U��:�Nl�8��^�ך���6��i���9!�v�m�ܵ注m4�7�Za���z�����N��V1	�cx��x��=B>̱�L$�L&k1k��V�6b�.5b�t(CMƏ=7�X5ᘑ��os�zf��ER�8TjX(�Զ�+�G�.&Wˬ��y0�+	�8/��қp���ն'�w\t���{���DN5�S�]�y�L�97ܙM&Z%wW�Ӗ�`"�Me����#�b��(���J���jv�Z�C�C�-�N9f�(B�����c�Dt��ϲb.bkyeoZ�,�/Mg�5Ub�
�:��zt��]�5s.yk�e�Z�y;�5�V�:jvx�gW��Ŋ�j�Ҝ!�'��xbҥM���F-Prt�e�+�7S�$�g2���״�%z��]ᩯ�
�ݣ����?	���^u�XG:�5�ct�<C��Gq2��-��۲�5fn�'am�lp���NZ��i����g!�-ZeS>�[�5��޵[m���B�s��dp�B��^M=f�,V��c�Z���ƈ|%~���i���g��׏֯ma0����[��`����*�]�
�
�L�)�5��s-����,xp��Z �HU1�>�(2���3م��Fͺs���+<>����c�[X�;|�*Ϸe�%��"DÃz���+�����MD}�c��!���¦7kƍ+�r�=�WR���`brJӧ)���1�n̦B���F��"n��D:�����/�X�tAi��X>����٦ �����X��4���|,���
��ג����t�KL��u����w{���hvi�>�VkG�}�U������Ƿ��B%K�ᖦ��}��p=��TW{��{>ެ��[M�iCi�CZ��I]���1V<+�,|�E�X�J�~+�Z0|�����[��t�EDڤ��zխ�o���4�w~kn�����Rt`\kӡUw~ݎ���8�!�>Tj�n�{�澥��0F�z��ǻ���oY5���M���L�1��ǯ�1�_9�v�+XjӨ�br��m4�0�����	�\y��8j�_�M��;������l�d�V P3�VJ Ϋ:j�j����w�O*m4�5��ϓn�����G�u��+c_5�J��z�s6oP<�h�%[Ju-��}�މ�V�4��q4��s![��]gEAO�h�L�,�<y��9��'b��3[�J�m;�L��-*�mZ)���=B�%k]׵�뤉�D���ӷwN�q�`�ʹ���7jt�=��������&��Sf�
�-����Y��v<`?>Z6)Bλ��䀂TѵAd��B�q\��Us]���>�����P�īB&��Kf��&.��q5�]�0&�5s���+�a���馢0p�|��)bs;>C��a�Ξ&u*rZm1�����Ψ���X���C[�{���Ό����'�AT�C�f�{ܨ���U4ki��@�ga)�ML�Ǳ,�uYk-Go�..*��e��9�>�+,k�;t����h1[�ߏ��X��ï>6>�Z��;��m��"��,���S'.^(3����}�Au)I������ԡ�e�D�(:�ZNY������\�}��Y�CZr�gv���xaŚ֝JV��M�و˳��}u,;�N7�R�)�f�Rl�5�K����Wsi#�yB�!^4R{�u)t��sR���6��T�WV2�Z��wxTf�u+��^`�+v��v�e)Y��
e��kkwEI��x��h�n������ك��j`�c�-��uHec�£]�>viP�pe�ڇ{�������V+L&�f��[�l��5(t7+2��zo��7+Xf>W�Ԑ���]�F�!��t#`����-}�������q�vY]c2o39��f�^�V��W6�-3����D�O_5���Y����?"�!� �P�)FfU�Z�1���bʍ"��܈�ZAU0cJH��"Z�,�)����2B2��"�Zd"�FD$�F�֬��V2T�hR%F�Q�)Z�*E��$cM!����!P���:�V{8�AW����8�����F!�!�GPϡ�w�%�[�卵i�)֑�'\7��^��C�p�n�=�q�VP�� ���ε��{����;��#%���1*8�xLn���-B���9�a+���=�}6�ö���U��nUh�F�)�LNq�z���M�K溙C��א�f�o۾h�bÈ�E���0і��w]Mfu-#1��ʈ�L�I\���ơ}�#�.i���O�q`l΁�R��씲u��,D�DG��[��
�&1~���ZM���i�Vj/�Ǹ������~̭:Bvԧ�O����ۦZ=�V��$�ȹ���1��븪i�}¬1��^��}����=95��je6��5�&����0�-��|�kl=�̯:Izg��l4�He��I�+:�n�5�ތ�ګK�0=v�z��{�~߹K���-�������C��"�fg;����oS��OS%m��$�X���H�;�#�a)ُ����:j5n��������ە����FP���߻}x�{�q��aZ<�k]�s��}�Pl58����\�V!��yt�g��O&^�ֱ�q4�<�38�\7r���wR���!3N���fC)�4�Cٕ�	�\5�߶e�e9ل�e�Z�5s)�Wg��'�\:�0�ɧ�wۗ�ֹ�j����PM8s�[�59>�n*�q���K6�l˼\J]G'��Vcd�:
Їވ���g�\�>��P¡�CN��w��fs}��H��u�ǭe�kƲw�ۆ��-�KN�{�`�q���\'�0�C	Q�=�]ױp'q2ߡ��̦�6�XC��tK���a�9���r箭2�N;F�
�H1��Q,Q�����lU��u�
�L��n�va7�h�w���et�0��z�g�<˟w����2�&(`����~g�W��l�W+��U^�utB�p�b�aa�(V�XC�Ҿ�G���G_'1'ن�$L?5�~u�w��uƻ!RKv���XL�<�~FM<B��g��x�Xp��#^�OO߃�� ��:顯{���ogZ4�-#���c�ƻ��S�^'S�ze��V״�ﳛ�����vr��6b�~n�#�󧩾r��u�9�+C��ȄC;Ճ���0����ˎ)��3�P**2_xx- `��z��W��Up!��e�@������Z�6	�興��J����HLf��Ӎ�o?On��tr����֓��u�nwf54�up���[ku0�1�7���m0��Υ�h�m0�3{fg=�էvS�-�.�B��n�7�~��!\<<*��x��+Y�~�5�.ӃZKjWpM$N&s+�w�{]|�p�h桑�)#Ko���y����M�\,}�X2 �4*��D�����׼kp�HVT���e:�d��	��RET�(S�՛��U� �%�,�7�TNx������s��}��Y�����X��x���b9�j�|��-w:�37�k{z�K\r�.�1sO�l�����JTM����f��g��;�)������r>��>�|%,4�dʝ��aѹ��^��x���o��q8�u�iӮBмŨ�3�ci��涙zsV^���Y[Oc���$��~�� ł ��������5�zS�p��J�&�#�w=�4up����@ṹra��~K�p��ե#@i�e;�y���w0�!�D��̬8�s}�n�bu7ل�c3m��i�u�v�HML��f̬*qۧϽ�d�m�4a�5n�r&�#�Mw^s�V�5ma:�M�[�m�{A����dj�n�^��p�Z�9gpM4�Amk���	���]>WN�'�P�!m/طzݑ؝v�=���,�8�#XM�~�k��܇=ow<��y��$���l�h��!{^|L��w��uT��]S����Y�f*����������b�ϳ��]&b�z�mb�7{�x��쮦:������{.2�N���X�O19�`�/~��7u�6���*
����gA�<�DZ+�"�$H�q�r�������.]�j5�7c�M1�Mu컋V.U���L���pVxަ�D���Y�^�Y��'�g\ݪp7bP�S%p=�!�����2k����z#�V����:5��'��w���b���p�243��(5����m�#tU�@�h�JD&=B{��/-߇�4���yE�<��a�M��x0�Td�<��vTP�ِ�.���^:��z'�~�ac�(u����v�_kg�4�kw �+���E�]�.`ѷ�aN��%6�U��n����b��8h�2�[���z��S��ç�	�W_U�c7��C�j����6��q�h���Vh�]Z#�Rͬ�]��>[f�ɹ/;.F��]|r?��1ԥ\�)RN��f�J5a�i�r[��}&o	X��dV^�,��{�_`�2�=�k�Ge?����སF�cE�֍#ºr��+��>84u���'KP�S,nWT�X�����~t�eқf��Y��Q��	�uֈ-�fV»�B���Ud�Ym2��U#&��(0Z1)���V�D���;��:��RŷNE���Щ�>�E�̠�.�,����6��k����;�Di��&��:I�u���y��a'bk�{z����ЍN�����m��{�s[������c�S�JTnAhP�����[ĢJdF	)B$�QR5$"(HD��ahFƚ.�زDc�Z)H�i�H��r҈�*�\�R�$�AcV��mI%�\Ei�Ei�%�,�?�]�|�w��Up��U� �"�+��zL7�D&G��޷�H7_��Z�A׹�p���k�p�L�
�-u=�qV^�ˆNy���'�&
�mzT�'v������� ���X��oK�v�W)�u�D��@�u���n�E��F��=����8w�(�tq���\?G��R������T#c���-[��'I`�\w^�	�vR�6d�N�����5��;�2I��F9���V��C���|�mlu�Q�ޞX��̮5(�/LxP�u�gf�|�PX���O�zO���:��h�[�4c(U���*�R��:_EM��K��	W�u4���t�����rI��~����H��Q��[����Gt1]������C���\���4�ZbW���<e�;�5��r�B��;%��۰��<�
���T���)��`Z=A���gz�f�я+h�Z�ȳ�.C�xƜV�7��o�u'�M�sӫ7#f�OE?��8��Q�/aK�J{s�5y��'6���_E��ڭ׺>�:'n�g�y<��,V���ҵ�s����'#K"o��Ԏ�a����(z"��v�f�et���NQ�.N�Cy�8��:��g��Іʂq(1\����+PҾ�����l���mf�#[�f�{'_��n#P��6u���]�0�j��:	�ֹ��
=UK�J�,N�U4�o5���ne�F��N�ڢ�.����	��#�VuEh�:���X~��1��1���_	�B�yQ̈́���^���;L%!W�v���J��U�D%�G��F�>���7��y�+�u|�Ⱥx"�8T�p��6!6��/��D���v �K��vVn|�>GNd>�	���Cn�ځ�q �3��\nn&I�f�b�B�u��{'��p�<�ݘ��?9���*�����3F�wP�n��v�J,S�h]�ME�dnnD9�l�7?UT��3���
j�������O	���6���>��62�q�^���֦��e�+�:�9o�Fz�����F	D���8�h'�Ӝ��	�宬�^��ގmH/��@�W�jA�x]�ٵhq�#*�V�R��u뤫v\�:���߫Ǝ9�z���K��G饇��	��Un�N�9k�<p�ê��wy�FW�YX�ʺ�X��P�:r�}h��Ց�4���ǈ/.}Lf��ne[y�B�FRN,�����k(��L��^+�nw=�'������@��,�ք�J��j�1`�9�g%�#��������3��?m虪�07����:�2i�?e�=g:pα�5X@��k#�;5l�-/�r�t\YӇO,v�y+H���B�]:8�/ئ��8V�[�8���?x����v��C�+�R�p���5���o���f��l%V��
a�:�<�����+�qwg������S.��c`E�}f&D�V�b�.qpE��7b&�r����'"�+8�W�Ɠ�5|�H������m��A�&\Ɲ��l���z���;x4��@���2.UgR��2����;�r�;����t��hz�����-u�:�Q�:˜	Z�% �:+����Z�yf����ň�$C7��d�[W�KX�No*���o�X��P�,*	�wogCvM�u���'�����h����U�Mw�w�h��q\	x�xb��}pըW1d��>��J�n�@�W�$�i����ju��՛��%t��m˽�ne:(��V2�J'Mf Q�I��_�-����O>[��[T���(���bC.褰�]]�eQP����YBY��rH�M��ɀUܺ 1yIb�?g!� r���j�
v�"�,�L��d&�H�ܵp�-'�nf@U]��V��9���k{ǳ��4�Im[JTh�r�TR$�"[P[�E�����DP[�"""��.����
�4�I����V�[�B5�eܵ	�;ε��3��6�Cm��NF�����t.�ȅ�t��&6��z#ބ�YG�A����u�oN�ok!Q��P�k5U��ج��XY�K��ĭ9��w���PF�ҸԔ����:ա %��[�)-Ƚ�U�#�� u�|�b��z����`�c@f:�݈�oaUQF��Χ���ޏCܪ�P
ˋ_p�'�=�U|y�(N�O�&^Z���m�	f�Һn�S0Ȥ�X��:b��(r�D��H`ɪ�v�T��]V��ö���z��	���d,epg�\�q�%�kV׻�\�.����eս��a�RW)M�+n,j@i_Dx��߽�뱄2���f���)�2�L��K�.�����s�'¢��w5m�l%/s�g��ZnJx�q���ys����e*ɔ��닾���!R!n���<؎ o�!T�r�
�nh�����2�qWK�ك��$� 	eU�gr���6a��5��b�N��y�F@ȷ0�zݡh����E5�{�\�x�F��v�Z�}Y���O���D��/v���-���H��KH~'h�]�n���_<���r�ڞ����(�|r��j����g$EN���	�*mB�`櫞�R"�>�r�_�]�0B6X[䤔��y�m���$FXp�p����!�y!�+��sT-m��̌�x7L���*�������e3��D̋^�>v)�a����}�2��Ќ�s9+�(�@�(8s&�TL ]p ��F%�U�*��G����m�ڻ�����:�&|A��*W�h�;���W[t���2�[��MI��"6�[X`л����[n�i�xR�=�����.��)��5A��v���E����T��v�1���U&5~�5�ݴDj�w�8]kv�්A+�r���'�v*����}���c��eJ��1Ô�ai���p��2ǯ���zS�v#�{=����?`k���a��Z�O�)zj�qp .��y���J��W����=h��w9˯0����7QSE��2���F�>\6.t�\)��7w3��eiK�o�u�O�pl�ˠ����{�]a�	K���/�{���ޏ.����敫��yܽ3-���{����;I�dl�v�%Q��3I�Oa�7@��:�˧[�o��5�J!�a[�������fp�����'�ƃ���R�4���u� �	RwAl����Sb�D^^(s�@��;�{K��:��;����<BS �0!p�$���z=us�I���@=(V������ 6���A�>�=�����u��n�ⶲnJ�&�N)�uIb�24$g �T�9C�؊Z�Ւ�z�b�0�]ni}�z�d�܅bIVZ��4+3��ԭ��r#�z"�2�tv��\�����G{^[�o�_dmI�ZBczS�J�M�3
vg~�ZCv;宱ec�I�n�[]�U"b�'�$�<uw$��Y@�]�i0�®&��3�L?m̚�!����;g�u3OW������\Z2�W"��<���A���
�,��	\@��HE�q4 �4w5��{I�>kNd�s���3:ʀ�۬Dgh%.�+au�<!b�]=j�v���H`װQCc�j�Z.OsWF�,�m�&uK�r��ޮ��s��w(Zs���qHt9P�e~���9y.m�BC%\����R��Q9i����N�ɗ
3]�4r��&]v�8�x/�_]:�VRA����Q�tb� LM hU��y��7U���w,,5vr�K�J�5x���C��52�b�!�T�3K�*��q����wf�3 RdM&Jt���)�19j���.�o+2�#W"(���Ϛ�|p�G	.��Y+d��\,���[�2�Fb�E�H�lm$$�n�m.��-��-��7q�����IV�%�Aj��]�kwl�5"�"�[)D���n��T���.�ʟUW��**i�-"���e#4�6%��wsio�q="�f�a�k[�;�ޅe<�j�9H�5��n�"\����Fb�B��uV梁|�䨩�׹J��;%#�5��+�V��Z���$L�q{ƒw<M�t�����q1�i��!����M��4�	��N��t[�1�1�G!�&����B���P����\QX�<9�ב���Etm���&�S1�v׷��+XȋYC���8���^gu�L��ݺ{oj����K�E�!��d']�/<A�Z~{����o�$�3���b�3ւPN��Y�}:uX��^�#8�u�g����<�l叧7�)>MݓJ�&����wxqJ^K��(�k=��k�Q�RF���o�=e���x�z�H�-�@�L���'T<"�������a���y��̚����3mq�=]�ڱ�c������-RU�Ӣ)H&TO��R�%_ĤA���b�.���Lo���V����`�Lnq��ݗ7�)�}���ݬ=�����='�@��O�����P�~��#}u����&�^z�L�d���ȼ�U+O�zm��R0;�gn�����:�^L3hQX/��v�MqO�cs���(��&��KZ�@'Z�z2C��z���{Ɛ{�.2bE- ���@�q�ݖ�^��q�"�ina�Dm+��<o��{Vt���l��LV�ٮ�d��qm(:`'jw���%
��4�ގ�,�%\�6��,�v|�E�Va�k�G��;;:��=���vv�:E�Ǳ�*l-�ѓ��w��e�Ѭ�~�'T>�t����%��k��X�����2�PBֹ���,����9[� ʍd/B���ʸ!�4�L��]7�F��< -���Zk8���b�v�ۺ���}(��T>/� ���/����M��g��
�,�QI��ht��Eb�Cq�%���8��v�c�H7O{ۉ�M�5�{[VS(��=דjdv�p�+��o��]j�D�k��ĐU�w��N��ݫ:�������Rt���}�&nn��*onh��U��.�;�hm�1��b�r�Kè���؄��B1N唒���ٞ�� _��5D6�۫�Ƕ��Vz5��ѧ�8߅��]e�#��"Oq���j'(AĚ�أF��rA�Eݹ��(���
��[9�+�>)U}��4���غ����n�sk��GByG�7ʟ���)��r�y���S*�Q`7-J��[�%b�F����B��8Qi��J�"��$F�pe\*�����vg����-hT�3�b��O�M���)���ΰf��c�k���0�{J��Q]���ݲ
h�*s���6��܇��F��i8�\�
�gd�@Z�"�:�aM>��'�����[5�!`3.���O	�Vc���)`ʂ�_����b�C=:)�P]Ů��X�BOck�+�>(���qP�����y�@���eQ�:sR&auvm����(a�x�Z.�?���e����	'-�_�($��5�&�(s�\�L|Ռu�a���Hf�ܘ�S��NTR���8NgZ��%Hta��\w�~-�of]V94�V��`�@x٠�ڮ�+{�϶�pu�_4s��o���v�VCJ����4���qX�>�d�Ɯ���L4Q�`���&V5��]+{j�D��9��Q�F%��Lqش�Z��o]u\
�'q4��=��L*OVކ����,��(�P�3j��̴���s#���g�#yVP�Kaϋ�"�V��;�W��\j,X���K9s/>M�Fg�ն/2�fU�%������j� �J�ܺ���u.^R�۸J��D�w��VK��d2�Y�X�� $VAR�
X�]7l���3�� �!b�*��b6J��6(�G
\G8��F�6���,Ti�Q�~����H$Q!h���"��6�?E �T�&�%�h�샌�Z�D�.\R��V�GAQg��@�t)��Q9�z=�WY)N�\��һ_��p�6̲�STKM�22�@�J��v�@������u4Oy��2��$��#���x�yyh~Z��˱���ԯ����Mn���W]uec�Xa�p�5�)#�j6�9N����,��\�^QRTɂ#��2����gv�Ɲ� RRަ����W����g�bh�_Y[�7(UE\���27{WE�򷵎D�/���lvjޓ�*C�"��ޛ\3%��wT��q��ܔxX�zM+�&T U��A��uFւ:�w�i�w�AHr�ZNX�,IطGGJ��v�e���q�~k�������Ѝ�����-��^&.+�������WJ�ʄ��j�!�,nC�m��usΆ���Ihnl#�����p�)�pV��#z;�~������9�V�����l��Sx��&�5k�l��M;{�'~�tr�ʫ�lj	%m|�Զ�Z|�b�H��2��_� ';�a�����h�T)v�1�W���b,\�Y}��'�[x�86ɯ}Y�}fj��u��-*�T~�xy�Q��wwm���|6=�Ys|��EV��y�b�#�YP��s"�\��@�]À`-k{�ڴ�Q��,�Ӗs��!e �E'�V����{�Qضn:�k /�H�fm�ߊ��ވ*i�u�aw�PY#����u��؆ )j�=[�z5��c�Ζ!�Jy"�.�Ժ�z�����ū{=ΡHW/Z��l�B���m��Y8].��ka�8z���
�`)��ToP�&�q̖7+
23�&�H�ۚ�-X�}�'Ym�gr���۔:��Y�UM��+(��~�p��K��/��U^η׽�&f�5�*�E�S2g�������+���������K.9������V\9�F5��7i?6�)rq����0��D��lh� #)��5���kŵ���'E���a;���6��ӆu/]g�jU��a�>�ڙ�)weg��do�<�x��Q�~)�c@r;}�Ip�ܺ�A���Xv�f1�P��s<�r�pq,ю�e`&�讧V�tP��A(���[�r/�Z	�?a�O5,��l�QZ�H���U@�N��>��y�Q|�UJ��g�c���Co_D�|��s�Fʷ�.Ŝ��vZɎ�]�X&�]�DgjcouT�T���l5Iڬ8)<Ħu�wB��S���6Ң���;qԕ~jؗB��v���g���-7�/�h-~V{�Q��5XlS��vou�>r���7��C�1(��d���*,���5O����ս1)� �p��Vg ����(�A�T�y�}�[�3>���L�r*��hn����J�!)"�8D\�p��s@�o��27gυ1a�6s��VHS�f�d��\�&N��{��H$�t)����bl�{�{��f��1w��g�h���xo������H�茬��Rr]��k��4�����sq_F5��5�7�$�yf�u��Gf_�{ںӬ�Z��U���N�:;}���V�Xn���n{t�偕�����#���u�y��\�:���^�2���]z/8���.o��YD{�(�6��v-k�]���R������M9���]����OVsI����DY��(b\������ηV�X��|ޘ�C��OR�T�y��ʌ8"J�g�FE��%�����=1���;���S� ��=�y:�6���2�Q[WwL�W�Q����̳��C6��ܽ"J���\���$�[�4)�� U�L,T�㢰қ�x�v1�V��R���V���ͮ���ʕ{Ж�����Q[�Q�8V�	�2�%PO��#54�	x�AE���qL(�K�$$"�cw]�˃�^"[�e�cpn��-.�HY11f��R2��]�n�e��K�Ĳ�
��wE�-%�!LU G�a1�� h��d �TҫY(��qakr1p��80K�v�p4+�.��YrT�-%���j&ffa ��F��l�Z*wB���7�?Fc���(.y�Pg��tۚ;uVMC�(ijt���ZfS�.N�m���y�筙��h��;�Tc�)��������!b�~�u����P>י{a�ף툨;'N��h�k�5�� �E�������Sr���ރf�;��Jԕɱ��K(�I:�����|͕[��3i1�����6�u�,�Wm����j޸�^l��&��"&#�j�W�dYW,;j��`��/��vY�������[^J������,��c��c#y��j�fl���(�XBG� KI�=�\*٪屳V��m���y���:��Š�6�V�.㏆G�]r:5�����g���C��K3�\!+ue<�.!_�����L���;�����p׷��3��+7j�ɶ:��]x5�U����Ҝ*"�2��;�tK�%R�^�o�·U�O[΄:{6e>q�\,L��׿V�'�Cz����l*�-�:�3���'���ɏq].4���h�=7�aD'�Oz��1�%�+Gx-�T�s/ZΌ��)��D_6��jo��:wm��쥒����v;wl$Z��Tc05�V�,Y�#s�|xR�k9��E9J��x2	}ii��t��˼���;�89uo�(Y��i���ocv�C��� ������}d"��#@�w0P�q{�<�d�j����4�+JS�N�������zНÆ���0����f�C�~F�WYq9gwb���/[������8K��L�G�/��7��(�Yd�*����w����ᚆ�>�c]�3޾�)Z�1�[1�l�1�
%@E\���+�Ef�u-&(�3��2)dR��7�f�[t6�����,՟X��-�I9w�� 9H7oW�=�QY��F� �K3R�qP�Q��+6��ڲ&"����:+U����M	V�]7��cU��ʞ=G�T¿����W��i�����]E}�R)󝆺�'0v�L��rN9+�?��"�ݩ��������CЭ��6�=bu-ɹV�wvb#�!�y��{ф����=��l�c\%n�u����l�Z��)�k���qsvo�|2��4V:��x`�E/M_z�D��^�v�h�0.
[^5¹T��7�ڄ�zl��5-�]Ɠ�87�Ƨ�$^���R����qI�ll�:��+ظp�e�vR�ָ�U�^a�e��J��fՊ�z�b���
�4�����b��eaV��v'�Q�e�%0�]�f��9Gr�"��dR�r�P�F�:&D���vT.(OGxd0'ß'ݬ����6u���C�� c�{Ѽ�K�������H��������E�[) ��:�<�qf
K!�x^h`�t��,�L�s�ݺ�}�U��7�N��u�q2�{��c�~�W�����b���~�*��GO�����IԨ*�1+6�J��`�7?.Ɵ����83��q�UPUUU%G��XC c �P�㙀?*��G���0�ɬf~���	��3��

��@�e|8Fq���>�ah]�I�jiL�ֺP��#:Io���6m ��>�U����7�UJ%����V�jTW�C��j�M�X�  .C�(��1�,�����	%�������A����Cڤ�����Mxz��G�K�$q<U������(X����Ě�x� ,�d���l)T#R�Y���ӌUI�oT	Y�?a��{�?cK\O���Y_ɢ�R�p��O�UAUUT�/�1۟��z�UUUV(��a��WJr��]�ș+e+�YN}��.�P����ܨ*����Z�C6���5��� Q$�9ɼ
^�)8�B��������BO����R/��Yqd*�y�p�D����nH���6}�ؤ����SpR@In ��o����"�f�T���v^OZ���x����tTWc����������5����"�$ad;�xHL�UU��ך����� ��)�s�J	.s�����o.*�1*������UU�X�8�F������� ?�8��T  #U�Pdؔ����X�~��P:�Ĕ'�vU�P]���h$����.��
 ����u�s;�nMU�y���6<���]k��a�����~3���
�:��I��uD���V<�x�'�x�{��?��Yr���I*
���s��8�V#�	H�Ow�/H�TVK�T-�1{3��C�՞'�^�X�n`��;��!b�qdI��òT! ����2�_:wc�+n�j }ߖ���|˝Xer�\��*�.��5r[��"yK�%�;�$A�R嚘;��@�wKu�B�� *!׈HFEU�P��&��{O3cv�2W�� mH[5�����b�%��+t�&���Y�" :��!x�G۟�.�p� �g�