BZh91AY&SY]�E��ߔpy����߰����  a
��� A@   �  
� :( y�                � d B  G�ǀ��>��     >���]{�v�=�wC��鷡�۰{��]�G���O{p=i�8s��J��Cãp��	:^�g�����U�#�ّRي�t*������  x"����^�ڻ�Rz��9ʻ����Z��v�N���I���PѓMp8���Do�ޫ/q�c��UJ�����g�Uݸ��zh:0�W�@ @�� g���n���Wm�i�'t��{3�UW�W�����/xk�I�8(/ f}᝴��|G�[w{��c�Hm�2wyU�Jz��n��:w�U��p��9�^�#l���n�׼���'gv^�V�]Ǘ=]of��@�3קg�*�zG�����w���u���=$WO]=7g�!�� �y��ד׽��ӧ���sޝ��]���ݓ��xy���.��Ά3�˶�p��,�ۏM���kKׇ��$�{��݌_(T     PQ�%T)T�J� ��)$U@%�     	T��*U(C�@&F�!�  ��*��&  	� ��10�ȥ �S@ � @ i"hԪ��     0��$�	�M��S�3*~���f��Ԙ(
��LR�(2h�h� `��M��7o8IĠj�פ-j���D-#��ldb�I�AQF#P2�x���(�	� EG��������(��uE�$R������E�[�!b�� �B >A����q��/	TUHIA��QQG����C ����!��B�����!��^�����ÿ����x�S
��W�N�$�n$DÇ^�=���$NY>��D������f8$�$[1����a$I0�ɉ(D��frb;3	<Ʉ�f<&b��Y"^L�D����$@�Q��#jG�g��G�ç"$��ǆ�1"=��n�8�t�Q���)G���:`�����71pϱ ��Ἐ�Q)���=,�Kɇ�A����G���2����>�F�,��(�VDP$�Ȓ�H�E�+�{+�ݝ^�2ղi�KFb�:�3H�1��6DQ�F��L��&�X�;l�Ɏt{3	"`�f08t��L'�8tf,G;0�'�1H������I�Lx���ĉ�\�X�����*�c���"9ل�gO�	bYTD1�	�%��@�#��At�x�F#�H81ي s&�ra0�f�JY�������:#�0�+1aB\3x��|�1D�"z��$F|ODys���0�DE�9l��a�f$Dg�	���I���@���U�&_I���,f0N�}�H�#�x��3��`�'��=:9.DH�~�Ӓ��y��(�	�(��F�:#0�)��9#�Dr1I�ÇD�ǒ�=i8baӼ����Z>���w+�]����Fk��n���Ϧ����dH�a&�D����A�,�IO	ӢB@���&^&D�f0��ID�3&و�f��	q�}BI�p� �b �$�T�ĔLGA	� ��A�]u'nZ9&Ѻ��_:�n��i;��N���1�rb0���1tk��ǄN-���*���:X�!,�#�DyوɘN��53�#1�DNv$D��&<��G#䲄������L"a_`�5��I�N�Ğ(Dn�ȁ��DG���Ib"#�D}��1e0�p�"9	'�;0��b�D�D�#1D��:ISR�LfSr8X'�DE8x�G��3"#qzc�@��(X�ℷ"R�,{P�@�G䄗�)��,L1�J%�p{	|G���P�<'��L���'��TO�&@�W��D�%1��	b&5b�c܉������xP�����8%�tC�	�D�"RΝ,n J,Fc��G�G�?5��y�#q�$�	�z&DF�$q���K�N�1$�%��Dy`��O�'��ĥ	`�X���ȟ����$D�":%��%���'����]����L�BSȔN	剑�O��CW�	�>�bh����)Ԅ�ID��a>�ve?�;x��\ƚnF	�1���T%��(��&rfNT�AO�RD���Ç�:'^D���"Q8/тX�"z	��̧Y��雦c�`�D�Lt��@����:>��ȗb6̸Ea�����sݘF�(m����ȁ0j0������Q+�d���KS3P��"SY�@�}H>��g�b�9Ꙛ��%=���H��Ja�ߡ0E�O�0�̙r"(��0=�3?"A&~E���|Q�3�������f����O�f���||���|z��Sr�8#؞�t�:�τ�g�	ɉ�EGO{3�,���DxG"���D��<�I�l�ע~�".%���C�Dϖ% �:I/Љ<�!������DrK~��I{����D�WϡG�D����1(����� ����(�"�pN,L�">DƢz=��Ȟ��'���0'D�"ŉB`��S�w�OJ��
�D{ �s>�9gx��"#0��&rfx'}�D	|�����Q7<�G��=蟖0�_� ������J>���=*b	�&~9�N#�f�87X�X��2�tK*�e,�Ӥ|�J(����.�=p��O	�"Ą�#����O�N��0y�x@�q�$IȊ���%�J&<OJ���IOН0�3� �9ء��٘�"p��	>��xH&0ÂdB"e3%�))}ɜ.�JQe��;�Bx�I�G�~��ô��q�JQ۸���Ğ��1�̉���4O�Թnb����O�ߊ}=~�0�:)�_�$����G�����	&L`X�@��R�x?i^o'�^?2�(�A	-LВ�'�tX��:�)"(��f����B9tL�3�=獦��>�ߪ����q>�:	c�8g�I<�����q���\�A9a�2�S��H$R!�}s2`��2�&�F��	"5�)E���=��#ߣ�}�X�?��'��"R����D_D����ЉɄG������Jt�j<�B%��~y��"t�bl���Tp�=#q�N?B%��ti��G��L��Q�8A�I{���=�LybX�D�O<bh�NK�
�N�'	z���ÏН�bR��!����%��'�xy`�L�`$�'�D�}H���cH�BH��3#�D~D�� D�a�O	�"7�!%f|rb	=���[�F�߮�J�����f�)+�;��%	^D���'D;��K�ĥ�zϯ������U�GP�ޱf&�n�:@�գӮ�֙q��M�-îȝq8I_"u ����0���c�$�%9���&D�1	~����H�{��4BAD�,�0�D��nq�_�x���b�#��Æ'E�0��c�0��$�=�TŃ����,N<��ǉ0�B7�c���D�DQ	���䂮(I���ŝ0H�=��%	]�d������f(�$�Bpg����ϣ�O�Ĉ��&'-��'&b���$=��Af<IBP3DȉBP�pN�	����������XISHW�u�B�pft6|�e���ӌL��c1
t(H2N��*�p֋̭1���\ӞL�L�*b+�����d�e��޸����tYs�Ξ��:|x��<2&g�c+w7ė|�*��h�5۟C`�����3n���|f��>}�uyw��:{�_��o"����=��|�|s� �}G�5����wYA��J{~�×$�w�W��R���u)��X�	a��W��ѧϯޔ 2T��X?G�=���ΨO�S��ɑ��07L�4��##����a�\��|+v�z�����|~$��5(�,q�?�3�ǚ����O��7���~;����P����;>+�6����g�(��k��N�^����Ս���+�ɑ�t������5��r8:��k�e2����6��;K��0�qIM��_�=�m�[~h���a�g\"{{q������CR<e�5�����?7�;�~�����~}�tO`��dź���E��ƆNG�(��y�6�}xJ��W]�A���T�~��c�s�ۛٺ�w���S���ս�T�]��o5~P���֋������s�}�|��S��k�������{�7N>��&���:2���;:l���&c讝�������޼��WA��ڛh�ҫ6��1���d�>�ǿ�����{5vt��d�8��>�|����W_���\ǆJm��ɨV�A���ǽ��9�	���L�J�q\�Gd���>���k����/��9���2|���Vݔ/,�+=QLĊ/�7p�p�g=>*�Y�����~=���B��w��qex��q�6������v�Eicr�+\�V�R=��)�Q&<��5d���|H�;@�iQ�Cc2S�dt�ʝ�����4�Zp�u�����L��ݯ�ݹ��7s�����~h�Ŝ$&_�m+!>M��o挤�OEك�:g[��fH�67k,��&�D�&�~���;,�#�VNϳH�fǫ��ww�p���'�S�E���6��s��Xdxd��wqH��1��Ǥ1��]8�M�n|�篫�����7Ih=N<���)"�;]�\À��(�j����wt�`�}��Yco}�J�;�����x�4��e�wv	�Uzl��޴u{s�v�o�}�P�{d��;��E�9/pS��������7�q;��0j�繪��=ǌ�̝��L�o���y�_׶s=����t��gޫ���ӧ��=�~̢x �����O�Ǚ�+��Sf˸~������Gfo����#�o:��Y�]sL���[�)2RL���)�C�33�擅-��|���4�<�73=$E�۔w��y������Vޞ�/�l=�;R/3N����"��Y�uHoq��	�8l1�,p*1iņ�u2����ʷ=t˓��ޯ�0���eo���e=Ҏ<z-�}�ڶx��Xmf&U�s_oX]_-�.����rS�a�f-'�2�Vn�O����}B�9�?�D���\p���LHjZG��˱�%�~�w�N��,��
�A��^6sk'J0�����gF��=:��tϻ���JG{�
A��gm4�7#:~���J`�������z�5�?v��6����`�������z60r��(`�t�V>�ӧ�\>�f��=���g��qӰ�}��a�]��T�!�W	"�h�y�������4I拾	#�.�p�Z�p҅M�ok�z{;������ǎ�L�Yކ������R=>���|R؏��B�/�Iӈ��,�z~�zL�f��y���p�r;q�w�V�������u�>�h�c����g3V��	���Ù�*G:I���ޤ����=i�ٱ�y�-��]o{�s��z}	�s��v鹏'٧���̝+�O_�6ʐV);��������}r������k`(��5����C��,�L���0
�0���ݵf��2S�OϽg�\,�Ck_�d�s�]6"�xr�_���ՙ>�Ϻ��Y~�|�>�Ղ�W�(���=�aW<�gv7��ٮK@�N �ɠ����%�\�{�`X������H�D������7�OL�~}�q*��C!��E��:��8]�D�]$��%�a�&8��&�cGF>Xfٶ2�����08y;�Ӹ�α�xu��/G{�|��������U��6�z�_���w!,�D��np�}��`�e
v|A� ��~(wv3��[r�T�c�u6�'���.���������:��RDŇ�?:j)��f�K�N���E8�@�1N� }9��=']��d5xio'_��U��iY��}��W�=0�%���.u���[�Y���Fk�W�{Б�Y��_���o�=Q�M	���z�^c�;%B�"�-r�6t����޻�������Sew����։ok�;��TV\Au�;u���״����{`�K vw'����hp���^ŉG�o&6��I�0�L�	/���v��a��p�?n=���{��<:������~�}�K%�}p⇰��v�>x�h9�?���rB�
oK=�|ws�{�r�s��ޭ}u��ǧw�
l�s
�[�z#�;Oۦ]���h�ۅ��,�3E�����;{Љ�ǫ՟n����J(�����d�(j/e�\��$ܝ�Ϭ�}7g�3V:IM�?_�^�����_�꺂�l;|^v�s_��՛{�������3_����n�d����kdA�zV�Xq#�_������ݦW;��;�d�؁bt�2iY��m���`Y�w�,��D���f��~�չ�c����@����3[�c�;<�$a�YLφ�D-��O���/m���[�s٦���]h4��gβB����i��x���o�{�9�~���ny�i�����s��;��+;p�|��޹}A��z��.�'27�q�h�;4�8F��als!}�.�����H�������I�{�rg<��[�/`�&Μ~~�>���#�wo�2��3�W��8����N)��������x��P�gL�1���f�<���_�(,]�_�32��~����p}VՙL�g�5H���B�==����W�ۙ�o�h��2����
�W����E8��='N�O(V�f�-�ᡐ��z������S�5��Eޕ0�³��qz땁*P$��7��>�9���4�c�C��dz����{������Jo��L�tÅe{�2�L�^�I���Ii��'�p~�|*���ؐ�*Ŷ�6o��3=��>WG7���%�A18'=x1,j��Et�dc���{2�b�m.�f��̥�`��[,�6e\�L�X�gM��$�m�SkN��4avwm��5��� �.%�����ڏ�V\i�Z�,�0��]IL�1:�y�X�dy�����!�ٶ���2�&�L�^x6��?g��'�{�HԾ�."/������-f-�cv���9�:��J]]�}m*zP��֙~�cV�驦����U�[�n�1v��͋�����
�
rHt�L���C^>L�$�I�n����D���	��LB9��+l���}7�*�X��o�	��7���4/՛t�e�Z���K	�T�����<Ԃ�h�AXv)�dފ�}�mt�.�j�Ս��ڗ��B~�)򜍷�%4����i����7�Fϛo��'�_\2�O��+�$<𼊰�/zh�Gq]��r���8��>2�kHеm�h�:ɼ�&u���l�%?}|:O1��OC�����q2�\7�X���z��Ɨ9�cv�@��e����O=�=��o��t}{�7�� �me�ml%T�"L�Ʊ�\���(x����f͇dx���τ��_����8�m�����Kf�cd0�BF���"2��C�DÏ�i�����m�e�n��`ij�J�n�]K�vt�h�Ku7���u�*Jm3v��K bq��l#�r��Q��h����M�X����E��P)��b0B���0廏1��HD�FAh)�2E���&x�77BM7�#v�J�(�b?G?���,��n>{�a�o������*���}����sԗڙ�A�K�Oa�2�b+-��-����+x�bA���LiBj�tz��JLvm4�0:6��k�\̳7@��v�fn��sB���~�I�y�Ն].F��ډ4��[=M�� l$vw�?~?7�m�zۺ׾W����;gl�[(bJ9>�S�[�-�)��m��][bا��x��e+�4Q�R؉k�5|^�_�A�Xf�Oμ��J-��^aA��M����x�ı��W��<BD⯅k�q!�3&\OHU2��Z��F�&FN#�E`F��YP��.�\��INg������9Vm���W�cS{��ұ\R��5���@	B����I��Ź�v��t:���Ii!ն�DP
ٷSl�ݿ P6	��yg$�DH	����������u"�PeR��CeZ������]U�*���+�maUWUV�UU\aU_{���ʭ�*��*���*�|�*Ҫ�aUWUqU\aUXO�����`>�*+�����U��W����VTUmUUaUo����*�U�U򲪭����*�W����U��W�ʪ�����|}�D}��}��A���|ī
�����0��k*��^*�Uz�J��W�����򶲪�U��W�ʪ�������k*��ZE^*�V���{	=H(A@�a؅g[��ݭ���
�����������U��W���v]�ڪ��������W��VUqUUU\aU_+J��!$IXDYAP�@\ #�ݿ��AQ�HĄ������T���gC�����hfdQ�����ӂ@�(�BI�A I<%	"'D��d	�	�����	bX�'����N�P��Έ�H�I"�"Qb'D���pK�?x��$�:ɓ,�2�:t���[�u�""&$`�@��'����H<���	�&	bxä�b`�X�%�`�Ibt��D�$���'�Έ�Y�:A��$$��(� D�,���N:�L=UXJolw/�i�b��]��~��-s�c�BV��ZSb0݃Rֺں�6lZV��-��Y�u�k�KS�-Wy�m6mq�z_z�Kj�jV%�RmeԒ�tִ��kB+[Z�o6�ZB퉍�-�\��љ&���p�OT�KaY�E���t5ZM\b�Z���Ѩ�hY���[�h%.m�6Ņ6���9&�"}��ǭ�ҨҖ�����U�X�6��#�a�ִv�X�2�K���b�[b��!mL�Xؘ�[h�Y���շF��0X¬�xHͮ�շ��u��f�;M*�oWr[6���RΫ����3hs.s� љ�E���Ֆ�e���t���W�\[B��a�F��my)��ȶ
/XWu~��aXB�lz�}q�6:���..�����m)��ζd��-�kfآ�����|YtΕ����}�-a��^x�\�̄jG}-������F�%j�غ�Am�Im���W���\k�i�'zq=���>hU� �&��K��]u6׭qn���i��.�T.]�m����I(}�I]tQcz���cL�Vfഷ6�z�Z;[ ��U�f Z�C6�t���,˝!�2�ۊV�0 ԋj�l��,f�.����mX�8���&��l���۴�K���[�-y�f�-"�q���F�msJ٘Ͷl&�WH}Y���f�u6�h9H땢��z7hʤ�ns��aՌ4�Ҵ���R��ĥH�%�6Y�h#Hؚ,u�M�����j�iR�ű:�� i�a�XR��a����k��RkX���L,���W�kY���ݵ���]���S�αvV\l��`���88����wws��>��7wwwn���ݍ���7wwwn���ݍ�����ۻ���c~� �~��Y�&�����%	Ft�<<ԟ:�@9b0x�ʁC$$CK`��]�/���o>��Bb�IK�Tj�f�k�Ɏ��im![ӭ5�IU�\DX\�c�z� �\�\E��ę�&5U	=����ř�=e�1��x;	��6�Ze�c#~{M7��i�G	Y�1݅f������^Д�Į +cZ{װ�m^[�C����z4h ���|���%g(�q��O�y��{�E�?ás��Q �}�J��bxrN�jM�Rt�=ᨗw#m���!��8�������j�{(p��ò�5���
K��'�2~\��ik�СtX����M���a�}�=���'�?~0�,K4M0��pD�(��u�O���DĻ�#ILS�O���zY�f�%�ˌ���4��d��VQխ�y�e$�2���.�a�e�m�#A��)(E�G��{2$�衮���i_�����ꮛ�Ԧ����\�{d|t����"agD��BQ�0���*|_�ފ��������J�u���@�ѱ)���33�F1c�"!�8P��'��ٵi�Ï����\>>�����۬��uF2�ׁn`I�b���^�]?Y��mӓ8�W��1�9����E���F��R�'ӓ��f4�utrSO�ƪ�l�j�ܧ�͸��[q�D�Ή���:`���T@��&�	��X���l�T�>�?gO�z��xo�L��#���k�i���/ƕ5<<��0�a���%�"�<��Gi�rϏ	��V[�7�&���l���5���SxaM�m_�V��xr�3�6�W�c��"4����ڥ��|Qba�����%	Ft�=?:g}��ấ�0v�Om�^\^��ͻ�xZ��'3+t�D+����#u�B�(
Ԛ2���
�\O$`%��XI��/-b����ŗ2�!��E`�i����L��0��ًkZ�"d��[���][=͵��Z�Ϡ���Ξ��Ϭ��8olX�oR���f��4�\���.U/}f�Ѻf�-��.�Jj�d��y+*���B�U��)�C)�Q1�2(p�-��y�l��B�f/Ǟ�����f��Y�8"P�a�L�m��VV,���f��P3(�ł��n�yOf͝	9%;�V���e(t�tԾ�f73;΁9�W�r��<&���B���r�}�����3�.�#5�kW#��Q��q�6n��馌�t��Ç�g�i�v�a��M��u��7ǹd���#M��o�<�L,�(J0æ	�Z���S�S@da� y�m:HM���`J�{�F��CE(�p`0���xC�p齖����[��-կ��eL�^x�ɲ���]��ˎ!������g|�����fa��'Ni:(�@�����zPf0�JHВ��$������Ge�]y�]q�.��:Î4㭺a���(ܶ�a�\���J�{����lC�C�Mz;mq�W.�-��$(Țm�Tp^2��cF����J�4VR��gI���Q�3+Up�><G�`lb�X�����͊h��p�y�s�8�:�M��Ifk�f�U_��e��<��]`���'J�0�xA�\�/���Mu"lƒ��č�TD�Y6�!��@z����<�BD�i���-�u����=�p�0<Uq�TH�h��1S1I�I�����"WOM�
J1ܔ��(�������:7Ӧ�Z7�ލ�{�ѭ���j�8�i������a�:@,>5���������>|>C!�,9"t9L�M�TQ�ل�-퇞��r�m��U��;��7�7��d0��=xHl߱sa��G녦
� ��%�������wDމ���%S�u�c���!}�ZqbX�a��e	B%	Ft�<!�QՊ��f2z��a��컫�����dj�G8��w/T|tW�I�����Yu�p٨X<0�ГP��j�4{9��t��$�ܝ���'֧�B_����6m���Hap|O�h�C���:O+J�L��
p�N��z<4y���n
��_6��u��??/����˖����q�M/�^�%���a�i~&Ǯyv�|����ˬm����8��W��u��:�yzN<��ϗ��������y�<��O<�-��<�<�O8�O#/̤��Iҍ+N���2��'DҴ���<_���~O-v�'�&I�GC�(���ؽ/J_�-����.y~O4_��\���y���,�~'�~O����qz~^��������~�'𒟉���	��F�8D[O'S����q<����<�q~m|O�ry�-<�O0�'���ǜc�[��:'O��x=^J�U�)O/L�i҈�Q:az8t�/M���Κ�æU��!�ݮ����?~��3b�\}3���lT�'����(�� g~5�vq-����t�l���p�۷�)	�tU���ڛ��f.ݑ��ȇv�;�RVZM�L�Yy���
=��0D�[�|gƕ�NU�S���A�.}�?�9�wS[$��A?�����G�=��ۻ�������������fn����ۻ���t�����˻���7�首i�4�4�K(ҍNpDۯ6񊎒�rI$DGc��.��e(9H*;j��=x��ucz"$A m}誴�����I����5�Uhv�3��{����K�$��y=�"#u�SxYp�R��R�d&�A6v�1[��msL���r���G�rHg��~�����UR)�J�L"�$���C��\�����Z"P�֯��swy�pm(�+�Ϫ�P�J"v�9�[if=���.�q	�C�D�

,.��Hv���o�����:�6�ᤆCv�C!����L��>mלu��ǟ<�-�|�.�ۏ6��둜bF�ץ�UDD�x0��Boq��d�Ka����`�H� ��F���ۆC�C�O�$@�	���[�ym�gӻ2�����&x���})U	UV�V�WQ\>�st?	�e�I�߻t�5���4{"x�6����F0��@(��ٰ��a��l`�{z�?~cje�C��8�~����嫑�?��""�aX80�Hl`��J"0��?g{m��Di)_A�����U�U�R�����UP��J��0ZUu�y����mמqo0��6�.�ۯ6�7rv�s���FcDTSm�g8���
 �"b%���D�f�5�jt���+�!�r�P ]i����!�#2P_�Ŕ�D��N�P1"�2X�E���{ϼ})3,�u]��0�IE��{��" �P������B����.r�C��R
"B���������M�̀�|�:@�� ?�s)(�Z �B�XFi�lCt��1��k$���\̦�m��B�@��0��7�4�hVC��4n�T��4�}�R���5�d��Q
$��h�P�G))ȭ�k�DE5�kZgdHE6\��qn�&���Q������2�RJU6d����0D@D؆�0`v��ܹ֚3Ȱ�H�򅲈�ti��F�0,a�J�' �P��ɂ""w�����Z�fc]f3d�� ��3�a���i��b"`&���|�q��AeuN%a��<����8۽���/<�/2뭺�o�w��$�
��Q<������MA��Y?DD3
"d%�����5'� ���DM$�B1A��=��ċ$S\QFI��0�0�H�J�1(~0� y�kR�2�Vݝ�\��m(����*����F�'D4��~��T�ԛ���VN���mW���evT�h��TI��o����!���P��P=4�"0�D�FSP`{��ȇ���paS�"vD���
�~��n|$����FْbED!��-�VMH�S�E���.��d���_�q��iӯ<�N�h����㧆WR�-���U��	���2	�N��l����6�=��sROD����IDF���T�jQ�DP�	@#!��O�lٲ#$��J��Z��P�l�w��|�F�"M�0J �z$�2-N��&��߰����In:��j�n�dͧD���Ԟ�>�;T���i�5!��/
ɐIb2k�L�^����xl�L��Oa�@bm��D0R#=)�f�K�)8t��P��HM�p>���{�wsF���2M2�~[O�Hh<< Dtp�4QCC	SDģ�7y��ID���.��]�f��M�ٳϞ~u���iӯ�$�J8i��i⛸�y1ٙ"b>���׌��&_7�=-&}�UV"!?��!bA(l�{m�A�DHp'�&$2J"2J�dP���Nc	�%�B�KB���A�������B��ul��m������H��S%9�It�(�}H�M.����pM2L0�BN�a�� P@3"��F���+�)4RCs�i62E=��t��/��-���QP�T��C�kq��7��%)�M�Ģ	^��IхE7{�SXXi��8���x� �,��3)�$��E��!�a?���2z�j�
���Y���2T<�Ƶ6`�iJRpB����)�ضO|�RWˤC;�'D�ȥ��0��$�05�!U���:��?8���&�I��pӂ'���؈����ES"2$�ϔ���V���D�|�C@j�AY͘Dc����W�r�`Ҽb���I�X����I+66J�v�_��y-��z�m�(����EqoI$�'>��_�|�������RO{7&b]nSGe�B]z(���V�ނ:<8�PC6���}��p~B]��L00B�1z�JDI���{,i�R��1�C��l�F��	��;2CX!'ҁ�8!�����a���I���8��3�<<7���͆��	bVJ#�ś4C�fLK�����w6SE �Ja�
T�H������L��=�d({2���}�6&�NE��a�-~ޓL�H�Oϖ�]�i�ںzC�iI�d�����j��O���PJ��є?|�f�I�8�0�ˣBSE�z?�/���SH�I3��μ����iӯ�-�y�]u�^|�\��� WL�y�nc�3Iu齼Ϊ�H)����C�LF&�B���R���͉Na�{)F&��.Z�]��"0��F�\�ߴ��Q�d"X������0ؐ�vc�=�J��q���EŢ�jf�["�#�Z��Túf��]�MvOX%'��:r���J� �@N��ԣR"�N���~�1l\�1x��qe��-_m,�[���YdZ�<��1�FVZ_4u33F�Л2~6h%�X&	`��>�4 Ȓ�ۆ�mz5����Hza�N:W�q����iӯ�-�y�]u��Nؙ�u�Y��{n�V$? �<-2	���T�.�D�����Љ��s���*d��x$LO��w�=��p��)�L(��2��#�qmRQ�~~�Q,��!���ȥ��)��,r,H^mmK��-}8����<�L,J��g�nY� M΢��9H�ž�i���um�T�k�e�g⢹H�2�5R-�}A���2$*�5ch�4~I��-2����Ec1�Yv����/Y`�V�f�ҥR�v��ZE.�--e����*���~q����iӯ�-�y�]u�^|�ܻ���4ZZR��:*��I�ц#���8�_�;����="MC��Δ(��d���-���c	����wi��6˷WB	�K�`]�\A3�C8E��Ւ���>"��H�.��H��-���-MR3�&�TW��u�d�i�j�항��K�I�q�ی0�Q�F�kE��s������g4�!����E���{��G�����i��k�D�mn�Ulڰa#k��њ-zu�O8ǟ��y����m<�O8��O"���a~av�6�_����m�'�_�4��N�'HM�IH4��:BA�	醔��4ǜ[�/�/ϗ��y�ش���y<�y�<�O:���O2�=s(������y���K���<��y6�8�e�[_�_�]��\�4�5U]����q���ӥ�K����z=7^��z^�Nק���~G�O��&�2��y��o3�?�0�H�Ri:x�!4�#R$�#����:��\�����弜m�8���9]�gJ�D����:;:~3���?���^���?/��V�L�^�N�cD�Q:_�E;\/Dä��N�4�JXh~��G4�|�&aΑt��9?[�[{;ܰ�"ݧEʔ�:�]˗r5^���f��.Уib$�.�#��ܙT2�(zW��%���	���V$fDQ8�;wFAH$b�@ll���w��C�-?x8����l��'=�d���9:^7؎����rLn$";�L��d�����2Zw10�%�C�X�xX��X�#j��ffqd�Hj�B����Vf<#�x��F)�:	s���o^t��9��įp�b<ӟe�]���b��V�QA�٩kc_t1ٽ�D�n��pAe)�F�XHq����{���F�������u�"<'�3��5��v���s&�j����oT��A��T�WK�V�#&�����o��v5��yQ8��<6^ղ�2�ԌBD�AVD��{�3��5�I�������/h��@���q��A!��g�	��ĻK�O�7nn٧[kg�>�w�q-۵��T�k���VsJ�]�x}�!�ݮ�eؚ�>���~i�f���e�a�ѵs[Vj��MNڪ�F�$F(�Z�6��`�}�$�ep�H�N���
�E�!D!�ɉED6�歫�)�P�۵�ƙ�h`�$ ��:�N���mg��s2�����Uww332�tUU������UV�3337F��Y�i�: �i&�Q�N�<>~*�Θ�!8�
#j6䐚m��V�b���xZ9$��ъ��룼	�j��`����ވ�򞥭̴8���&*\B+5˦t��B�nfլluXG;TW+-�5�[vk�RZs���n��[e�h]]�T�y���U-�ЬtK36��t4�Wm���;Y�b�nҍњ��7��ǭ��.�ʪ�l��w�Ѯ�i��>��{y����G:'F�R�sr �E*���F�Fs�qH{���	wL0(�_&�f���b6
~��=�7&J3ϼm���� �����c�7��O�D�xC����g%�����T<�`����Y�Fr�ޢ�?�8Jm�3LR���"V��y��J��D��v�0|�Vm�e��v�ɿs�?$bC8S-����3��e�v��cm�)��:ޫ4�=I���������~4�a�	��My��e�[u��1&��'�$�D;ş�,ȝ4s=���Xo�M*S?uzl�D)�zUX͙
hv�coa>]ܖ�,��ܑ��WYp���r�[���R�e��ˮ�˔��z��.���f��ho"jBX�*M{l��ˈݝ����X�C�J�/&	C�Z��.|�>�L}=1��?U��M�b�N(2Hi	<;�]���)��V���P�o�8�?x�i��iF�8"xM,�Ot��֙��Q%�RJ>66��IQ��l�?z�d"C�~����2p���$�5 �<��I�Iӿ.�ɢ�5O���a<�g�\
�������5�+����k�k�2�S�==>������ǂP}�����ןf��fj�Lrֶ��C��f$6`w|�|�|(n�H���w��+i\��\j�h����k|)�ۮ4񦶆��SZ��51TӋi�\fm��q����t���y�i�]mן>h��"`H2��C�UTC���W2NCf����&�|��!��2~~�ى-Q�V�F�a�[��"�H���_ޭ�a�~�tcT�Wy����bf2�-��Y�+��i�g-��d�U&�����j�_{>���7O����K���j����sy�S���C�,=gƌ�h:�+�S1�V�S�6˕���Fڪ�j���-�i���^y���t��-�y�]u�^|���oҮf&��m��c�l����F�u����CO�xѰ��4I"��1�|�}�L*�0riAY�6H'�#��pd�7��k�O��@�F�rƘI���mM�K�עJ��-�ar�]>X   ���<gH�L#�`��m'N��XZ���.cc0çq�t�����#Z����깯yN?N��g�kz�~j�2��Ð�D:h)��n�j����9��s�T��|���[�T��v�9[}�j��.�m�{�&3x�Þ����z��h�_��ɚ�6|�V�J�k'�I��t�!)]}/����B����ߜˎdRێR�����{V�I>N��&�����5[~�%����~h7I��G�y�ǟ�m�N���y��e�[u��V���Mc3���I"��Fa���&�C'j�?6������j+^�4�����1_����"m�6�Jw�U~,2y�d.�D�3��;�\�}��MU�MS|�M���In��̟���z��5���묑��u���&&�l��dH�����Ӊ'�;L-�f�ƈj��2����k���7)2~)ӧ�I�j�������m��>n�N#�Ͷ�M?	�	��i�Q��ig�S�%�2�;�UD0�?���p>���֫CA�;MB���x3�CV,�/�����ʥs�a�����>g�uȓo���n�������WZe*��-iBZ�]�4'���M���o�fһL���/�Soϩ���f�`���vj"l�K����M�[f��N5��n�K~}L>���g��'İ��8
U2s��	�X�%b�*�c��xim�y��^: ���i�J:"xM,��ݚ�
w@���ZR��`tCZ�n	�+���
�� ��ۙ�xm���>�Tϖ�!�u��j���<������u��`��JR�w��{%��s����f;�H�}�v��0qh�6k.�Jr�)�@��~�i�&i�\��O�|�g^���g�)����|����<��+�0��|��VS�S��|�?~�z|M���-Y���.d�M���[v�2�D�a��'��"i&�pҎ���ѝ��ɲ�&�lx�m�(��q��>P����5��L_Ret1c7^`X�֠_G���ꦈz����3�U�U�  ;R�B���&�Qd���A��'mI�i/q�ֶV*�"�Cۖ���8
���M�
~���C󚪗u%y�[9o�/>[,-�5�ϧ�7�˖c�d���?Cf��ٔ�|;s1��8O��ӌ�!}���91�vH��W�޹��3�1��a.�g>�#���yb��Y�ӣ�Z�"�#���
lء��	.�����޺�4����~ٳ�L&� N�h���<tAI4ӏ0Ӯ��Ϟs�E��!lc��bI$�6䆟�V�U���ukk���iv�䔔{(MS�e:���g�M�6lA����oe���a������ьbSg��t�F�5]��>`�zr��wҳT�t�i�i���|ˍ^.��1�����nVj�G��tJ"��{	�͜�;a�B	���\i���W�}.��5/��U�i�x�/N�c��~g������qm����w'�������L��]���<���Z��d��'�o/M>c��W�S�	)@�M��1��M��Q��������<���̸�b��yzy�7'����y���X��<�����e�<��O/�/�/��ĩ���)�0iң՝)�v�6Q�tS�:R�����Θ\0�0����m�c����k���<~~c�?&�7?4����~a���/��]Č4ڎP��ai&I�Q���VI��վyn�y�<�����Zi�<��/-�����<�1�<�������&җ�?�~)v84�'��-<�������<�y{y�4|(���k�8s~�����(R����M&��,wur�jX��Dx�q��$r�'�#"6�:�u��XRD��M�'��Pwas�	�q5kh'Go������5���j>�gV�o��2v�4c�!FE'V���'N��PG��"ٲ���l<k�Ɉ;=��������333?i����fff�ª���������nfffn� �K4�M4Ot�-�y��u�^|ߤ�I�v�	��i��{�0�dү�՚c�O�&�P�a�1R���6 Æ{ڗ��sx0fA _�:K�\
�I����a��eZe��O����}�M�B<�1����m�ֻŻN.���s[Je5�[W���f���NW�Z6Yxn�ݮ���˧���/q�fZg'�а���XS6w��������y���t���2Ҏ'����ѳӜ�������\����0׃��ǐ�E���7��qz��U�1K9��.I[E�	���e=�x|2������������Û��m2���~��ç��Ζn�ßzh�D����;;g�Z�?���u�Nܨ�i���z��ɸ��Ϻ�2v��y��������O�E�.�[�����2뭸�a���H4�NQ�D�YK��m��g�z[w�>���X������&�b|�0��V���>�lItz�©���D��i�"C&:y�9|/��8 �K[jM���mcHR��\[�#X�uƮ�C��$=（G�˾�D�9&��ir��N6�́AUr*M�&hгo�t�6�@�j3a���\�EVjy:�z�ן]˼b�0mv|�ND��D��
"2ӫ�l��g���z��1D\[$�>)��b}�g�z�kS��5.L�S�S�~~�'b��˯�my	7����|͑F_ �(1'��A8A.F]��?^�8`�`��F5����،"Iv�<�R�Fu��4�<tA4ӆ�p�<&����UQ&�}=0��j	�~��C'������r}1p�=KJ	F��s��ؗs�HS�ϡO�m{aD�im0��k�i����]>J�P��������~�ߎq�l��奼�Rn�˱�&S���Ӿ���4Õl>�2JG�~J~�L��E�j��6K�މ3M��{�WnEr���i�Il4m��m�矜~m�$i�(�xM,�1�}��j�V��7mӷ<|.|���!������g��K��P�ة���
w�`f���i�i�s9��W�>u)�uY����a�O�(=\N�4��\mM����?D�G��G~-�n��Ye;4S?v�̸���b�t��Nɿ�؍��"Su�x�֛,�ҡy_���\�j���5�&F���e?3l�?S�����~m����<��<ӭ����@��	ęi�eTg}UTCe��s�#�1IO6�.�����<?kRM���KL���S��֛p�E0֮a�Z��kO�O ����!O$A�ݭ��b\^��i����k�9�S'���f�r�f2��g��ř?c��5K�z��M:�\�i(�E2~�9�k2����~Y���X��V�nn~906h��~�uzp�M�X���a����NpӢxx|4g�|����X��B�.6�Q���dWm��V���a䤒RbcN�.�B	�$��4V@ "�ֹ�V�KU,T(*H�n7 k4�񵞪�VUj��J�G�>$�H =��h� �~�Z6�E���{��p�˞�ۙ�}+�Z���{���|�Wr�W�ֹ]FHn�0�L����ӌ��1[~�Ԑ��������!��C�!��PKþ/�kͯ!�G�x���^[��qoۮ~����+�$�S��Z2~<��
���d�o #@�0�d�2'ș|�)�s(��y���,;CӁ�c��6�C�&�!�֘8�C�,�?~<t�D�4ӆ�4�N�>Y
��ћ¢�M�kNe�L�Sm)c�W�UTA?X�5Y?n��1]�#߷�Kħ�UD�����A����K=4ja���<�ϩ�q7T]�S��|��]�����7�-�"{Ȧ���)�_��q�VÄ�P�C�'���s���{�$��}u��ǘ�� ��6l��;����6NJd��Oz���e�Gͭ���y��iî��<�̼ӭ����y�.�qs�I$B������\W�4��Q�닖���(�=��ޏm.{
v��a�Ek�b ���7τ�~�g�'�Xl�O[1��ksZչ3K�KN�f)C���s���I�f�W�r�0qq�0����'ԕhb����w�|n�z��s
��զ��nSSP}\?j�%101YcRL�Vi��u�j��-�q����:�:�<�̼�m����1�&&[Zi�m�)�UU�TIO��w�����it�R�7x���1�v���].��T�,�O�m�%y�i�FK6�+����/��l����1K0����Wv��V��>���6S���=�h��/�ɏ�;N���m�1O�J�r��6���W��ihp�qن\�l��#)���<�����?1�ky:����'����K�y�������yq<y-�<���+�bm�2�:\Ɠ$h��	)��YIiF�W�nW������~q{F�//������Ϙ��1��Fה�+��LD���m�痧��c����������N��:fN�0���7X�ե�tS��K�
t��^�.^�^�Nץ��ze^�/N�e�J���S�������n��l�g�����p�aZi)��i�4��2b0�r#W��7'_��k��_\��19sƼ/�v=ץ���z;:w����<�O����.=rqk�??0f����~,N�S�.ˇ��l���������Q��p�~u��kg~��i�I����VzDBD'v٨,R2��(�k�0��T:���qY�}�v̰����R/�3BC}=�i��y��R��) ʤj꥔j�71�ǘI�ك!uL��EdBB�ą�ws'&#\�X
HR�itRMh.����Л��݅��JpӉ�6�ڝ&�b�{��"��L�<�Խ�8���.�uf/�3�����Z��ͨ6g�q��J�j��ڰ��0�1*�)��wl��Ȅ���IESpj��A�0��a˙����xh\J	;a�23f?^�4n�V*Mh@�<�%jy	(���\=� �6�պ2q�\RA#2�Ĥ�n$� ����]�X�^��1�J�uC۝����fa0��
18�v��LB� �M,-)f���E0Mf�ٷK �,���J�5KG�溺�А�ǳv��[�|�=�����L7��lZX0�#m	H�s�lݍ�YU��5�Mwb�w�!-Ɓ�ئ��m=ld���RLK%�?�a#�g!�����J�����:	
�0�]��#l�_�}�����B"�i&���'�
���\�~���ٙ���cUW/s337v5Ur�333wvUW3s337~ᤚxK0O0 M4�Ǆ���ɫ�W����;~�2�m��Ԅ]vfv�icf���Zo)bm��`��&2� ��R�6��EIj0�se.�ph�;c�L�H�J6���?+�c#K�R����e�����[u�W�Ú���x��>t��&5��c�3.���i��Zjz���fK.���1�ff��}�	>g㞝A��AXn2bcDM(PȶNk/��ۺ���Q7h�����]������+�Z�#K���2��FS��5Z����Y�Ѳs��4�S/b���1Zo��p�٫�ߛNVi�W���j�.��?Rg��#����Gd�Y�$� l�ՔH�?�E�������)2�N�ϒ�ɪ��:�J��v�q5M��[�>yל~m����<pӆ���id����C���|�b�<O<��f|�������bh�|R�O�[r�4a�B�xh��rS�����XZ2Rl�ߖl���NyxZ����1L��m�����;�ܘ��)�:��.��V^Z�]:�a��o��:ѕ�t���ݗMUz��SL4�:���վYg��:쑧�D�ܻ���&<�?<��m���0 M4�Ǆ�ʳ�fOR`��nD着�{��-<�ߚ֧���tȨ����$�5a��!�}�[l���=)�"a��<��x�~u�kK�	tR�.�a��5@1�V�h|/��ѺSA���?/f�am�V)Ŵ�2��k��VԺ�3�!n�l9E���NPPXC��Wߛ�2B+3]H������a��8IG���i���LH4�g��N	�N��z����*� �1�$�=M8��̺�F)�ݓ&�~� h@��~GD.q�!�F[�]�8��.�Kn�n�i��Y�?g&��wH��7�b�Ff?Y�i��*���k���d�KDn�~��m��g	�>�aݾ�)�6��uV7��G�E�B�{a}�y�n���̲|-e�Z���XR8��~i����iî����̼�Ll5�%�&�i2ɑ8�V)�&�\�p�H'VQ@��*�njhML4����d���6�����o�u4C[��,Է�Uux������  ��V�T���yjZ6�`��s;�:�I�!�	����:K�Z��f�3g��.aI��8j�(n$Kj��H��H��2��̲xb���x<NF0�F;��|�ٱ2a��*E;0��s��(�5�K��e�աջ�˽S�j��?#x��ODC��<-\F���~�٨{G�^Yl���#%��h`��~�yg��..���7\���4���wӰ�0���02�UX���"�S�D���<������{L�H���?6��?6ӂ$�pӆ���ifl}�L�DM�D* �'��h�Wz4#0�����M( �6����9�_!�ƣV�/��̒~J�������nU�mk�����~K�����?2�<78���h# ��!�b��G�y#)s3.k�TEO���r��n�e����a�Vq�S{����bS������F�G?v>YKy*g�>[N-��|����m8u�uיt���g��NOVx�[i�[L�B�}$�D8���H�5��a/̿L�_�ڍJ\����ҝ�.f��N��[m��!�N�T��+-h���>�!����aLX�m�3l�(��n<?N͚?G�05���}3�Dm3�<,�p�0���aXCC9�pa��o�^m�ڹ4<ó�p����'뫣�<m������ǫ��f��?m�m����x选&�4�xK4�f
���ј�N�/U��a�j�p,�p4	�lZ��C�w�@�>�Y���+��,� @�Ļ�Ķ�2�0���8���4���6�s���I"�j9�q�*S廟�5�B�eEFs�R�6~�p�R��~V������ϩ��J���j2��3�q8�H�a�$/1"I(�W�>�k4�S=��X~Gu�q�i�Y��0 D���`�h�4�}vC��Y(�ۍ�����W��G:z�,�o2�?\31��:H�%���l��=����c32R�.v4C�_f&���Ŷ���Φ.0&�Ap���� ���y�|al��s���E%,*�xT���en�|�]�f��`�OHD��UY���m��b��ۖ��S��e�Q��`���t��*u)��:�Q=����&O�$�b�n��`�5˗ƚ>Z�y?Ti���$?|���:��cH�In0Z�K�IN�p̻����fگ����LV)��E�4o>�4J0��L0��K:�:��2��ϟ+��qW%UCZ�hU*j�x���l�'�i��Ugy���i�|�&��tv�q�}L��#�ěZe�Ҽ���<7�(a�;�m)�d�N&C3�(l=�6w���.���t��m3���r�t&��'Ν)�"*}B �>��5u6lݿf%quY.�Ħ(�5i�����dW?SO��;O4�2�&Q���8'��$�,� N�BpH8'@�	�H��<$�`�&�	%��X�I�,K�(�A�""xDL�"Q$� �xN�:"""Z�:u�uh��Ӭ2FYDdA�$�(�D�<""'BAM(ӆ�4�OibxL$L�,�,K�腉�����0��pA�8��� D��DH đ$�H�y����=�4��4�O8��y���_n�3�zz��BK����n:2�N��wA]�����/� �ˈ�j���Ex�s�_u�	�PAd�yq�Cd6���3�����.����=�>#s	�KHtn��iBz'��w$έ��,K7���.�i殬;o��zy�4i#�����!�;�Z�!�a�(��eB4PY�C0��Ukͬ͞���R?r�HJi�wۿ}�{�������e�ffn�Ϊ����������f�ff��4ҏX��x�c�����̼�n����/ْI"�%yf�_��O�<|�����n�D�s,��չ�i��26Q�i%)�G���=)=]T��`f[�h�K�.����Bz�)�3�{�U������O�l<=�E�����`���m�l�kg�ٲl����<��6��WL+M}�>�D���:E*#�m_�8�:���Ϝq��X"@�F�p�<'�,��w��������UQ	�p<@YE��#Y�"�����o��Ӯz>������:s���W[��5�Nc�Xꚋ�j��p�||S�}�����m�U���T�5���W)�u��)���-��%.�����ϓm���2uK�X]gy&JC�_�RUѐ�!��h�ý��~�n��)]�%G.���F��e�֙e���i��, D���x�h�n:W�&��e�,�1���)v5��hJ�0�S28RE���>F�][}�5*>�7���R�(�]��ΌE�A\# Fn1u�f�Kl��� �w��娋���N���	�c�@��QF��GEP-�0���q�f�n_f0����z�0�"i�A*w�N�9���߻�����0��o��'ꎬV_��[g?IQ���n'�=�\��䄝OX�7LSl/;��La�n�k4�V�5�΢�B�4�����A�����yCR!�a��Ӹx"l�0��z��>�V��0�{���޵��1���>bޥ��Ry�iז��JZ��}ӥ�`��?~<t�J��������KC���$]$�b]4��\z�l�F߲�yؓ�9��A�S�S��l��VRղ����fof����[uY.����ӿ�W"GY9kWN�֮H�=�����0��� ��L�\țGљ��-kh�r{:d5;�$�9��{�I�ȼ��OA:2K!�`{��r�UC��5�a��O���X���-�H(O�><>6t��Xu�jFL:�M�&��*� �p��߽�ĦR�r,���g՘�3P�C<�y���Ӡ��L�$�~I�l�~5>&��	<��U���g�85��L�c�?%������C�\aZ�$g�#�y��Vd�d��]kU*%r���d�=L���!�ݰ�Gk!�+�n��ui�me�a����H(O�,饜��X��
�|UTA0��ܵ�v�J�=�n�V%cɗ���~6�'�ѧܫy���B���%5E�ɚ�6��e�ʺ~E����=�I��\�sՄp��G��m�e��l��P����i��!ѣ�ق�L(rv~V�S`�f��[lѣó�2|}Xqե_$�5M�KKD;W[G)����ԏ����e��]p�Y�0I(M8h�gM,�<�
��?+��V1G?592��j6.Y>R��Z���O�zh�ۥUg2���Hby��k��V�rY%	�%��C�UO9޾���2hW�*c�5�	��]��I ��|Ֆ(�A�O�R �Wz���u���CF
�IQ�FsP���\��	�&C��TYX(��Ԙ���2Ǿ�w_�n?9]���g7�e�'�:_�:���FP}�"?2*Ȟ�i9C�D�F��ɾ�Iv�}_��q�0n�બC������Q�~)��	��Շ��C���%a��\�\��7��~?i�,�&�:&	"%	�>>8l��p6���X��UQ�����Y��<�?2̚��ۗO;�<��0ؚ��	���y<���e�5��������q̦W�+��Je�;ϫ��Z�^a��=z�+�;�~Tf�{Gĥ�=/��F��K~	����0=�rO���.�g��th�ry_�$�(	��Dӧ!�{��*�V)?Sty��Y|��	gD�$D�?4D���d'=�ռt����!��06j�o��pU�G�N�i�w�!����#ㅾ뾒�F%�m��]��M?[-�h�s�t���U��}zc�s[FP`\��2K�x�'�����=OB�"��j�Fo�����>�M	�z2,8Y4 �C�w��z2y�y:pѣA�Q�a��0N���s['��|Z�;�j~(��M?`�tLDJ��O��:p��|b��\�x���զ0���UQ�F}��Lk�ᇂ,��]{�L�h�K���δ�����$[C�ҋ��"��عLdSY�.h4�َ���~2��C�����=O�v�]���b��|o���O��z��#�D!����β���'�F���5s�Ml��ha���#�q�0�������q��\�6��Z歶M��'�"d�MO�ف���<tDM�tO'��8'��
 AD��N�,�`�tDOCb`�'��gO1%�I� �DDDO�!�D�IAJ,D��"&m:u�uh�Ӭ�#,�2D�$�0�	DDD���� �D�J4��Oib%�@��`�X�%�btK L%�%�:P� ��	�<X�$�g��'ɂH�Q$$ �#Q4��M,�|F4T|l�4�)J)feL��Q0W��rT�v�����\�-�Fk�^�����"���b���g���О���0S��;�;!0t=6&kp�n=�\�3�m�(kU�1� � �D�Z�U8�UF�AX�V��.�w_s{Ah�ѨCmXТ5�����Q�2[4�e����)と��yz�VnB{�����-I���{`��h�fn{,�f�ŕ�q�DMz��솜x�c�]�����0�jū.Y��a\�� �`���:�Kٍ�"�����rU�j��w2-�0�{s�I�`n�Be���@J\H6NY�B�����/l��\|[���ՙ�4؄�>6j\s�kj٥N�u+��/s�t��&�=�7+�h����@%УB�@���i�ű����IEl�Y��v�V�������]2Sѩ�B��-14z��a�Χ.a��s�4�M��F��َ����c<��<{�\u��+/j�H;#,,ɵ��Ԗŗ38Ɲ��W�Z�D6��b�P����٫����z,��W>�i��n�MM�)��H���!�}��������{��}�Us2�33wwkUs2�33wwkUs2�33w�i㆖h�%�������G����ֵ6�- �&�(����K	�n�4!H����@*�;:�v�m�i5���-�ˡ��b�#�ƕ�c��)W��+V�Z䦴b�ta� �i
p��%jmrļĎ�'T�v���J]x�!!�Q��.�mM0�	���9&���ݦS<_��@��ea22��o-����X��q*H�!�m�A���'8?x]1V�Θh­^~Z��Q��L<��h�����Z����u���+���<�`},D��)�}.�_�f�yfݤ�I�e����~ݢ%�����<��Hjv�h�A��|���fi��9���9'ɱ48a��+q�K��-�u��e�ϟ�ub`�&a���if�,���dy����Ʒz⪢	�)D��Қ-%VL�鸸���z����Ր�
�)$���V��ZqĮ�,�ֿL97:a�CD����m��`����z3Pܥ�c�&\˖���*�-���Xs��K��0^��?5M��'���S�S
J~�k�H��DJ�%j%}֫&���/μ���&	"aF~,��>�W�TP�l{�UD=�E���a�sXq�_�˗���~Y��i��F�����8�O\������Ρ�,	�Gc����eg��l���tb��}�$E"����>c��p`�B6�5]�uU0*3Y"!ĕZC�L�Gk��Fr��ð�
~v��3��%�L�X��k�ʹ�M�ˮ��>u�]a�e�\y�ϐ�����$�4ʅA.��Lm��5�UDg�Q݅o�#���A?�~���	<��k>:���l?��h�<#2�n^s��q�0h�*�����ؕ+����A�~��8A��n_%oM�㿧~a�L8OV�l����a��7W�j��MS��-���5�d����|��XjOߡ�TP�O�9	ᣧ��~4�KJ0�&Y��fb���w��ԟо�*"V�6���y_mp��4��<2eY�7��=g���>���[�
a�[�ǂ��v�M���Z[,&Zƛi5��� !'ϟ��>P�=���K���Nh�9���<�YݑL�C8�ȧ\p�\Y�2O	'�RGR�aS��1^����.�z��<j��a��״�t�}H�ԷϏ�%z��~G[��:�]n3�Ja�R�~s�L�v�a���j1��|y3���tk�4�MY4�1��FU�pA�)�'��}���J�|�\Ėa���Ym��L?&�aF0�,�Ƣ�@��B�9F)ߕU��zh�>�O�M6mV�/��2o��֪!�ҿ}䬴�u�H�'�]q����Q`�����I�r�&���ɨlC�����̙nh�`����h��ؖ�?'�����!�ը�n����߾��c;M!�j��ql��T6i�Evj�����饉�X�"Q�p�L4�K/w��r��dU)�Z9x���w"a�=r�2Z5蘆ۍ��]5H��ؒ{:�fL�gk|���󆦠�6}��ߪ�lyV�k�LqB���|F�*N��ψ�)�~�2=4a>���2,K#���G�av�mW��w�\~Ñ�lMZR�C��6o��hD䧻>����H�m0�M??<�ϝq�Xq���N��8t�ɉ������U���SO�v���->��n\Ϋ�>F��:щ�E�̊3���|c�{��	a&�]�3�ߤ����S2�Ӂ�{��t{�y0����x�)�ݓ�﹄i��ˈ�OQ�a�;Y���Gg���);5��<'�5��Ɲh�Ѻ�晦ܦ�V���y��h�~,L(8a�Y�NǺ��`=l����Q����uA���ތ��"�J�)3-
SB�0�!8��=k���a�$ho�X\>������ ��o���RyM0}�\�C�h`�jdV�	�H�'�&����z������+M?�q�Qu�2�N4���rD��~��e/(����ҙ}_���C��g"S��������r�Sݸ��?S\V�M���z�i��o���n`&�ܒ��[�ǐ<����|�K*��=Iu�T�����vw|>.����f�����Ɇ&/t�>|��e��m�]q�άD�
0ᆘif�wrp�T�DIU�Q�Ub'D��0O��E�Ws�c�4n	D�>��F�/��M0�]�Gk���[I�Qj��1i��(�����D�?w�Sa~'�`�6�p^�̭D�fj�)�љ�Zي����0�p��r�s�8'�Ч��߭��I��D�G��S���x&�2�i�0�k�ZFp�0ӏ�~qםs2m��F�4�N%�p��A�(D���Ď��a�,�K�<'�<'��
<$�DD舏""HI$� D�����'�A�N�[+FN�uZ:�:�u""%��� BD Dӆ�4醚x�K0�DA0K,Kı�$L�%�%�:P��G�D��:'�J,� O�L(�HH D��N8pD��P��e�&s޻b�$�93\&7m{x��6@t�4��(���P8���:�<o��p9�uVy��w3���YYgf���N���R�ЫYJo
����M[���*vV	�V��Me,���p2)�u_nXﯗ{�}��]<��>�ej�����;�.��\�����Q��
7�{���-#A��nfN�o��*�=G`ڦ���PD(��y�b"���r��z���s�k�ᾼ̷f�6��&�y�������ww�����ff���s3733www��������4�<&���%��aF0�,�{����*o�}�z�e�oU��eb��"�L��s��Q�E��ӹb�4'�'�ٗm�GZ��t��u$n��G̲�#�V%|�����~�����<9~W���t8pL�gq�;��s��T�c_F?-��Fj7Y�^�ꙥ����#���4F���(�æx�,K(8a�8t�>W��7�]k!W���D��v�5�AR��(��o/	�L���\N�Kd�I�g	0�>�*i�����U_4�6يS�K
nŬ�fg'�vp��<�8���8��up�t�=ͻM�٭]�ؔ�����Χ��<`���<��[E�W�C�jV��~y��_?8��n?:�ϝ|�(8a�Y��Ǔ,Ep��O9����:��
6oOx�Ԇ���@0�1�e��*Ġ�	.d���qu7��i�*�]ʌ�.��sKCE���x�I�@����K�G�3�}���W5����VÛ����ĥ>ٞ�#�lV��=щ0�<$|(\��A��pj�������'�yٹ�����9Dd�~w��>��
#����:i9<��Z�0O �g��g��O���0����mkJ��a0D֖�j{3�W��
'�j9ie6]f�t�3�6�����j�x����X�0���ibY�Xq�q�|�fIJo�a�fZ����;�����,Vp�8zmlB��v[�M��|��NN��&	���X��|Y�GV��4QG��7'�R����Ji�y|�����	蚐"~<�tM��v�L�1�z�B�Q��qw����!��Gi�D!t�>��k﹕�#�!�l#D�5+S�K����ͣaf��<`���%��aF0�M8t�a4��R�;��F	��O_K畡���5΃
'�n��O��0J�?r�l�7C��4pFpZ�}�z��;ϻ�?�¡M,�{�}*���O;��z`!��#�|�2�B8��\��R6��N��E�4��wg�~2�
!��\��ц	���>�k^��m|��\�a�q�%����|~0�<~4�&��J�8zp�ӇNȡ��C)�U��?~|�i�ڭ�F?Wj��m�}9����]GEL��!&�ⱶ^�'�}�0�&1l2�����o��c�m�<��<Bp���EW���'>$�[�m����"a�E���e0�d>w��>B�Oи>9Gra�Df�MS}�T��Ym��ŉb%	F0�M,�2���?{Sz��+N��ޚ����%��bf$�5O��ASk,�q^Tc+�*����*���"؈i�A9��t�l�h�m�	
�OX�\
@@�.C�I'�\�����{ !���f+��n�(�,!e5����7��r|w��a҉g͇��_ �r�6&��hOߠ���|��_u|���r����~�ذ�⿏���5L�\f�VF�B����ы�V��8	��r�<K��?f��Zc5[��ۙ�c�O�=����ᫌ��7�f�K���~u����u��:��Xu�q��>y鄴��oq��j�18HS��0�a�1ι��ɨP��,5>4#� ��߼����������9^Cf��Ʃ��W��/M4�֔ϑGx���?h�G�_Wz�:h�趘{@�O9��)-m^
�|��/c�����_�=�2��O	ΰɆ��K���u1ְ��ύCE)Ft�,K(J0ᅚt���<��s3Hߛ���w�U�7L���a�]�Ŷ���%3WOՀ�}t��S��7�K�1��
"~<0�=�;��h�?`�^fbeL�[A"L��r�b��V��~ҧ�԰�L�J��U=��4D��0���5�}4Q2O!爭�k1f��V+9ZѪ�v���z��(�e�,���ibX�BQ�,�ӇN�;��&�fj���+x����m���Ӭ�8S��o���П_	H��(k���s(^t�I+O��ɷ����"��o���v^���Ӂ�3���F�$֗����sf	�4���Fk�4쑪��N��P���ѣo����������<��:��'��6���V�8��<��u���O<��0��Q����#�|�]wR'�K"P��,��,O	�F�(�H��8`�CDAD�H�$��,�"X� AHHA8p��@�aH�$���&	D �DJ4ӆ��4�ƚY�1"H�	�D�0K,K+"	,N�xO$D�8&	�D�,D��N� �"Q�$��H�'N�,��3��x���ۖHl��VZ���V�ˠă0�nEɛ����^�3������N�6�+����WS�2�G	�Bo�����{���H�ӭ�Z�E�HA@�R�YI��Mi@__��>y
��y��LK�#�i����Z�K	0"6 �6���6h��E�ҁl��RNC�|��wt����(��jdF4�qM����Ev��6,�N�֚rUn�s������	�n���:0�=Tõ��:�|��1�tW�r���͓iG����ߩK���d�]}�1JQ��T�ڳ
,X1!��kmĘ>��f'�&M�LK����4��I4�,,��Z��Q��j��D����nl9�D�=�AOO:5i�޺��Gd�߻T�(o�FTIX+��!R�\1���3��\4uXS[kQ�b����/%.�*�L[�c�z����i ?>>�c�/!�Ͷ���m�H�e�1��O	��J{���{����ww����������ݻ���ջ��������������:x�L4񦈚X�"P�a�4ѣ���oɠ���H<2���]n�D�%q�X�:�θ�S3L5u�W�!m6YB�YVn4�0"I�an"�i�&c)�1v[ģ�vf�fɃ���F+n����\���-ٺ���a��h�+v�a���l]��9Z�1*����y��kP4�F�Э�Ǝ�Ɔ~�Ub&o]��:g���
�q�Y"=��!XaMi��;p�7ђRD�`R�����?qs� "�Ǜ��\N8������u�»p�A�j��V���W[i���<���^w&\�����ߟ����SG����}�+ta��m��O��ũr��|�a	����/�	�e�k2뜌��#��`�X(���ѣ�مa�3�Ϻ���Ӈ��4��"if�"P�a�4��5���!�`�P�W�f�UX����3���?BFjs{���q�sߢ�is-��j�PӒe�1�b��0�Ӝ��h�[�>���e<�N����jQ��N��q�%�6�%e���ee�i	u�>t�����~��0N	���á;ID��f�y�Q
H\>�����:?p�e�DM,��J�8af�p�x�=�C�E�����Sp�Y[�I����H�%/��ǝ~��Jf�!������i�U�'&j�2п�<�% �٨�������e��U�͉a灇�lN��\S���{������f���G$�,83��F��p����Gg��o�����cq���M���>[�'�Y�x�DM,��J�8açNq�>�L�]ndǾ��D�=8SY��}�'	���'�_!�J<I���D'�!�P�J��6�y��siFW�h��g��菁������{�+-��ϤJ'J���y7'�Âx!ɡ�}MO��L��+�;���C��`�FC���ј8Q6nb�;�78l3?}�Um4�v8Y�?�:h�0�"if�"P�a�K4������O߲>���Yn��YB������=�=���w�i<�T}�M�:��QIV۴��D�̭0�����n	W3����Rc4� 8���,C�
PM\��K,"{0$��<u�n"�*$`;�YI���=O0��#�m����\\��v�8&C�va�>�����~�OD��Q��I�aY�#UĮ�4�1O>�>n��l#t�������?bLJ��|;9Ո1�
ZL$��$&;�[Ku�>�o��M�j	�;��2��ӿ7Ki�i�u�]y�K4J�0�f�Y�x�4TMMd������D�d�˽�=:`hOgǈ�*�Lؙ��0�l�Vi���]�WQ���RDGO�S��x\6%B���Ç��D���Ŭj�e�(��-�P'�|����?2�h�U})r�$�M�=<�\Uf]��V��DGX�Xm��R<히�����h�9�ɩ�,��4p��~4�DM,�ƉBQ�,�K4N�Hڨ�;f1bɉ�1.�Mf�/��>��5�&#=Û��y4���_m���!���x&�V�]���5���6z'��U���;�n��ɑ�IC�Rz|��i�y�OmkEӋ��&�Dw�Q_W����7���I}]�j):'��z&��)�>g�ny�_(ی��R�+��-��N<��]u��6�:Î4��<��ȸI�Vg1�PQ
�m�tw�U��5�Ό��v�Hl��<�B�9��3�>zd	��.�U��N��$��!!y�o�&�3þ���i�a����$��+7NS���,�i��F��ZV�0�lO|����nC.��+na|9�m�Ke�|�חQ�L����|"&�i�D�(��i��pr�14�j~����U�*f��Q5!��b>Ա�+�}/�u���c3}�"���oU���[�#nI��X]p�Y�� 8���2I�����)�䠜h���N�#�� ���ӕ�"��ƞ�A��>�7���k���gȝq�����b0����2��&��"~9°O!��=8&�
`��a�wt��Ͽ&cLpEUtX}?	�-m���l�hޱT�i�a)��hNS���8��%���<5
k'zS�?|W���c�YD�OO�K0��,�"if�4J�0�f�p�y¹�`kF��UX����P�0���Y����qt�Z��U�_�|sՇ��E�s'�uZ����8�)|/����KWz<4#�釰�4�@A�G��ZM�Dq۲Mi�4k5��3/�̭�<���8{4a�0�����CݔM�b���54`��bv�-��M�N�ONp�"t�a�ae����H�)�-��x���x��:ӭ��&�ȏ�����X�'��a�<t��#Q�,�$�D� ���(DN	� K,N �	I'�ÅI�A�0�$IDDL�D�"'ӆ�x�K4�L0L���âX�%��%�`�Ibt��x�"$��	�,�� ��G� ��H
N�%�+�زc�i�p^��{1ݨv�ԧ���)2jC���l�ڟ	�N��z���U=��yl`��D�<�b�=|��b3��z#:��z`��j�ڷ '�=����0۞��Gϓ[�p��� ؁"�sk�3�F4���y���yz�S���5w�o����ӫ� �Կw=�f]�߶�t����www������n����wwww������M<i��i��"Y��4J�0醚Y�~7���L>�Eƫw"&10�t�n�5�kᝰ��D��[|��ӽ�Y����I���[uG�U�I�#K�p�r��"��%4�U�y<־nf���:~��cL���b���n��ɛ����6-֤�?S_�y�|��q�q�κ��4�P�a�LK4�a�b>����V"l�!������kQ��|�8�;_SL6����Fs<��ܻe�2�5k�2�Y��ɜ2�6~�j�r��ߢ&$��L����i�C������m�Ty�e����f�Da��lЙ9i�|?-�nI�w��qr�0�-�k��ST�H�K����S���ύ4���g�O%	Ft�4�L�����U�d�$S�k��Ձ`��>6�M�������|���W#����|��IR���)[-n��&�ң��
�4v���$��)�Y	��R��)S��!a
�Y Вv�)�&�"�l���0�!�H%���t{�P�E"�N�_��jc���^�0�O�٤�R��a����SR1$_�b/l�Ke��2�K�R?2�-z��Cӓ�pN�A�ЏN��(���>D���.3���y�>dG	��&�3���AA���|��=��߫q�U����^uǟ4D�M<h�%a���+�!0>���j�҇��kb�p�I�D{2a�J���Gk�����1�\f�u|���@R(�FՑ�:s����/W����!�;4C��̜�ϰs<<8z0D����t'�Ѝ����GF�	`�L�TуN����x]��Μg�{�H"Y��x?xhO598n��E����\�0�j�q��:i��X��i��4�(��&�i���m-�N����a����ߡ����ѕ�j#�-����5�c����1+�S5�~i�>�n��]�<��:���4u�k.�J9��8 �����(�g�7�?~�j��׋��63hO~��7M�:���a��I~��)�DJ�2�r�S--�^u�:돞y��a�q�m�v�ˑ&�0�F�(�Y5��UX���;���[�8p�OO�g7����6`����ڜ��,B�tD��(���Z��ҭO��O~=!#�'L�����3O���[��e�8�!���&���ys3_���>�J'��.�`�4"~�E�C�ׁr)�4��MϤ��#&�}L��M�˷7�b}_x��(��4�0�Mi�u�i�[y��7>��8g̬�^��c�%�.��mʆn3UM��Kl��#�E{'��_�>��lV�Qe���]���K�6kU�fu���)
��"`���$����N���<�Ҍ@��iń@�w[9~A#.	�1+\�\]v���w���
2Ƥ��_T�4��b���)�����n�76'=]��zrie���kwZz���u��|�z��yշM0╓�1�%<�MS:A��eZ���#�<ߔ��T֊�YZ��ۭ]G������=('e3��K�T�m�e�[|��\u��<��0�8ӎ����˒K�����S�\�X%Tڪ���7�3��֚t���wk\&�F,��b�����3~��t�_2��-� �6�|���l^1st����|�� �� =�(�	P�H�D�P�Kj49�gA(:I�
f���o��Q��KGP�H{16n������%ie�Y�"ag�NiBa����çNn(��
�Z�(ƉD��M8�l�1��N��:��ӆ�m�S��۲['��Im��%��Ӫ�O!��	驁�����T��V�D�Q& |��X~��I��.�h�;�sZ�R���CG�}��������A�O�T�'1���S~�s�a�s�wa��W����èu�u��8���4ᦔ%a�����O����TS([��=�!���B���Ce����U�氺4̧؆Mtv��=����!�=0s��iO�n��ｋ�3�nL%e��-R>idF�������V��W�u���q���y�K�̹����7�_I��s��,N:s�sM�OJϕ�_�\�F�icX/�>'D�a!NRE��I$�(�G��='�O�f]>,XG�l�BX��(ʀP��	%�a�;���桑&�29�*�EILʳ��1P�BUB)	HEBRP��*)�%T!	UBQZ��B*�A"�	dH�R�A�	HB��JB���!	HEBR���R	H"��%!�HD% �%T�HT �B��!)�%!D%!	H$!R�J�D% ��JC���%T���A��"H�"�J�EBR�BR���2!1A� �B����**�����0Ab ��A��0D��#AH2�2"1FDH�D��#H�"0D�""0"2"#" ���I"0`"D`"ȉ�%�D��"#A"DdH �@F�0D`��A"DdD`�#@F	2"0D�"� ��FDA�#D`�`���"#DdF	���1 �""A�����#"A��0H�`#b$�F10DDH0DF� �A!��#H�A"$""#" �� �`��DdF �AdDH"2#" �"$A!0D����DdDF�1$D� �Ȉ�`��#" �dDFDD`�`����%���#dH �D�"0DD" ��D`����"0dD�F�#H�b$F"D`���"A"1#A��$�`�"#"$DF$DF����`���D����A�#"0D�Ȍ�FDA
�k!FDH�H�dD`"D����0D��F�#H�`��$F�FD`"A"A����FA"A ȉ�FD@F�F2"A�D��"2"�FDH�dFDH�D��#	��Q)�DA�0��@F$F�#" #"2����"�Y�D`#"2#�DdDF0D����$FD`"D`#��
A���	������"%IbJ$%$�� �`,+$ � 1$$�!($# BFH++�
�	!@D�1	��%�I D#��0A��z=0D��5aB$@PD�Y�HD% �BT!	P�4���J���T"	Hc0��"�J� 2 1�HR �dA!JA)AhD%T!	D%�JB!)b�J!%!JBR��20�
0AH�dC�`��2BQBQ)qKBUB��  ��0`�K�2!)BR	U	HD$�#
�� �0D ��J�B�����B*��"��-�B�BRP�BR�J�!)�abȨJ�TAȂ2 �Aa��"*P�P��B��BP�D"�)dAdAd�i��>��HEB�J��dA"��"���� ��BRP�B!*	HJ�J� ��`� Ȃ �" 0Ad%T% �%B�BUB�P�BR�JBTR�B�J!(�T%!��2 �� �" �2! 2 �D �"��T!)B!*����"���D%!A"�0A! �!	D!BUB�B`�D ���"D#"�" �2 �B�P�BR�%T	H�	UBUB!)�JB ��BUBRB�!�PD%B!)B�P�% �� �!)@��B��BB% ����%BR�JB�P�%!%T!	HRJB!)��%!�
�%!��JB�JB�P�%!JB�AJ�B�D%B1���$A�D	HT!*��HB�BA��2 �D�A	P�%!P��B�"�"�"� �A� �"dA`�D �2 Ȃ2 �2 �,��A� �dH�R�J�!)A�AdA��dADA �Dȃ!	UBQ�J�EBQ2 �"	`�D` ȃ�$A�1�J�!	H�J�BR��J�J�B��JA`� �DB"`� Ȃ1b�F
��JB!)�%B��A*	HD �D��JBJB*!H ȂD �DA� J�!*��!	P��D`� ��A�%T*��R	HD%���T!)BT!	P�%B�B����� ��"�j�D�A)	HJ�D%!J�@�A� � �1"�"��J�BT!	PD%���!	P�J�A)	U
��BT!	HD"��%!Q	HB��J�!)��BR	P���"��%T*!)B!*	HA!�JB)	HA	HEBT"2 �B0A"H�H �H�FD`$�B*��%T �RP	�_^i4bld��a1ui��پ'6���HH����"�I[�o�k�3��g�}�ǚo��	�@�\(�8��tG�����CS ��<���n2ۂ,����LvM��<�a|��B��Z�8P����_���k)�nJ=Z]��jnEQ��n��+��?p'�a~�`��?�@�_IE|���� �F4�z=C�K��>��u�yA������/�	�w� ����6?�`v���d|�E`nG�=t~� B0��d���8���. ���ᚗ��N��O��II�L��x S@ָ㑚�@��8!�n��%�B�#�2;�M����%A ���iK�T6hU��T8Ao �b  ^*(� �z�h����l(�	V
l�;�N��v��z��q�1B1@H@���B��
��B�!�"� �V8�Hd���:�������>(�#�r�����D�H4�hg����G�����<�$"�(�u�����|O�L��.>����o`� �9��فZ d}���;�V���|ĸ���7�8����+����狑�9�r��<�R4_��`C�
��<憆F���:���x�ƕ@TaOB���:҉�Ӊ�X't�Z�u������]31
7� 	F
@��A@�D	2Q�$��Ń��5"��JӈF�8 y���@�l2��'ؔ��1Q�CA0C,Z{@�b�\�>�$pKL�I���j��4��:s!$�<P	��\: �(�}�+�8�w6�a���4��t��>A�.�K �Ԝ�PN����9@��{�`�$��C���Ϩ~c�z:��Ew���D�@����{�Er��;uf}a����/ppM��8D�)��O���i3��1H�:xe�70 ���.�P��n��Gy�] ��}E�ܚ� X4.0Ǡ�)��0�q����&("�0}��.�vbޘ�Ni����Z \6}����Øn4tL��D��$(���)@� l<���.�� A pb�-�8���	�>�~C�p��" �t(5��z\N�q�s:�- �����jH�֔t��]M�������"�(H.����