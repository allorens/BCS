BZh91AY&SY�,�k�*_�py����߰����  a7{Ϫ��   %}5�   R� �M���  �\È
  BB	UT)@
��R�� ����]`4�Ӣ�*�  � ���� �
E    P�Ǯ@����lͳٝ���4�7m���z��8_{p�@�: ��������<��%}4Q������U�0h݁���� �=i� ����P�p> Q��(6`W�GZ{`����Q���z�w`����n����� = ���:��<�;����2=  �wF���� � Pp�|=�@� �p;`(���;�hkF���@	���A��X4��05� �@������ �p �Mǻ� U��iJd���ppQ�P@JA��`�]d,(�����4��x h�h< / ޷�n=U(PX8�Kjh(J��Ѡ	��Mk��@8� (5�Eu���Pn�4(�T;���@                 �AE �P��47������&� � &   jx@��H`�&L� 	�12`"{J��Q4�d       zJ�F	�0&  �`*j�"M�56��?(��꟤�1R�@ԥ��&&��MS�z�@z�4�6��������߻�ϝ�=ٗ۸Cw���������늧����zq�|����]go]���ca��3fa���0}�ɼ�@� ?��f�AZ��~������⠇\�������6���lnG��_�9 �n#��I � 6\B>B?��%��eUTg�y�3f����>��?��I�h���#�40��sL᫧���_���;�BZ{E{��&�:�����l�FĴ��O'���Nk{$�f��&�a� ����9RYқ$�#d��;�LGd�D�넓�M��e���dב3{��!�_N��i�{Mɇ��:FD�M�D�rx���]8Y��֥2`��8���ã�N��'GmW���-�a²%�L��{)��6X�\� �$�ґ=S�y���Jӯ2�lw:��YB#�<"wl�<�'{��r%u�#���:D�w)�D�X����bm�H�nR"ܮ�*�'JjR'<��΢#��Åjj"[�H��P�SY��"Yo%"y�Lr��ﲴ���M�r�%���k+4�9w+U��"m��N�+��u0��Ҵ�epٷQ��"cr���SY��"m�H�u�$E�Vtw�Zt�R&��\��D���/l�V����ґ;��1�Ý�M9��U�W�I8S$F�Q�*�'�ʡ�UK��'r%k��u<rN7r��#؝eRt��]<_Y\.K�nD�jY��rt�D�[&�$8H �O���j�Hx��j��Dy,K})`�������JÙ7��57=D�q=��r%�����'=��-�V�*�b�i�Dƥa��	�����#SǤ�d0ʉ��:��T��a�#Q;"5,�ZE�]G��b䫡����rqb���.X�+K���$aY2;�IM� �!�WqsRs|����tm���[#�ʡj�S��"�#�#�)�v�]jO�*iO�B�Q��>��=���B�	s�?�=�v�q[f*)BB�C;Ī<�Ow%\l:ԟ�|��K���dSTVJ����)��q7뱞��X�d�0m�(0[�,��7�tbx�t����9�$�z�y3��͜Y�	퉍��9�:��%��%�N�U�n�m;��N�<�t��7f��LL��3���9�I�Ѕ�"N��ͤ�g!%�N�i���&k�'t��d�nOlJ��,�l��"��88+�/�̜�I�w|���%�9�2JN�'�3&k����N��&2b8$��t�eo$���N	�2pG�'����Y���K;by:e��	�Y�퓛I�,�"bA1��9#�W������<Y͐撼q!�'8N���1�0p�(�I�ܗ�:':p��,vt��Nn��&�M���'�6fY,h�x�E\�/MȖSd��&%zB�7�&���"a�$Oy"x��Q`'�D��	C�$�DM��M�H$D�'��69�#�i.$��DGН:Nt��O:���K�H���8Q��D��I�Rt���D��G���$D��M�a&$Ç&�|��J���K"xH�Ģh�NĈ��:l�$D�$N�,��6:�X��"8p���I;Ԉ�Ğ�B�k�;�Å�^$�z$��:lu}IpD�;����H��'�0��kh%Ĝ��M���G]�x�M��� �ܔ5*Ol�lٱ"ZA;�1!�'�҈��"X�l�̳fY`�7B]$N�^��9$�ӄ¼xKM�8t�u5C����"Nv�5<&�2x��9��Z9"F�Q���tLP�3��Scd�082t�:")I�<D��z%�TN3���W">���`�{Vn]M54����D����,���虜��&�!'I��R�5ii��Դ�'�}·J	���A1�X���z������#ޕ������/
ב�I6n�� ܇xp}ڞM�����N&���}G=�ŏ���9N
\���Ʀ��^�������F��eL8�'�R�w)*ӽ���",�w��.�X���Һ��2a���Du�թ������{4���:q�J�Oz��鶪l،�DG"&�Ԣ�M�dG���H`Ƣa[ji�DFL:;�DG��Z��!w6=��:tޚ�B<�DG2�a~jQ£SH�sH���	�ꈝ��,���S�7ʈ��Q�l��"=�Oi�*&mL:WZ�A�'yR�zH���p��eI��H���-�J�L8VښE��#.����">j'�asu5��T�������*&mL(��B-TN���B=$DRL8&�0�ʑ(}u-�J�L8VښrP�e��/�VV�<�Dk�<���1)�jx�'L9֠�/��!��J�_!Y�SP��_ej �TQ<I���A����אߦ�٭���]F�Q8p�����85ʞ:7ʉ��"90kR�H��N��C��H�=*]@�V	�w��6����1�ѩƹ1֛�O��RQ3�%��>�u%����7(ou2=J�+�:m�+ݩC�Ԏxf������CdL7iI�JL'Z�a�]��ϖ��F��̾2xʻ��F �#0�0$¦a�,9CmC�C�5�MvMrMU��&��NďkG�����ɠ���H�V�^#�aA�Ѯh�h��G�G�G�����7����&�#ă�zZ-�yQZ��)���j=j9E$RL�K���q+TtI����Q�*y|�W��� x1��i��ϼ&�Q��,��m������x��aH�xZ�]e��xw/����Y쌪�$KI3G�N�/����Iv���g��KF�#�h�iu���,p����5��}�M��zfM'��H�a�H�S�#�H�H��v��G�'=�pW�P$�<�E�#9L�|����p�V���0_S>�x�:���xX�yB��l����ʜ�e&�V�y��c���H���:�N,��3f:�6;ܭ#�(ۨ�5G���'���D�b#�%eJӯT�m�L:ܤE�]6UΈ��V'<��΢#��Å�K�����L(}���R�6ܤN���Xtw�Zt�R&��\��D�����[+U��H�})���L8;��&Ȳ�lۨ��r�1�Xlw���R�6ܮ�"yԱnV�V�>���nW���-e'K�+U��"m��N�+����S���iȞ�Vɮ�N���]d�T:E���]�ʞ�O3��x�87r�ޑ�N�2�:{�W��WNIcR���MԳ}��鼉�2�Mx:Hp�A*�Ui��k���Z�oQK�JE�&c+��i̕�2o�dgjz���A��":��852�D��U�1�WLz�68H�9UI��Odx�9scs�$F�NH������W^6y�r%	����V�3q'�IܐrCrwH䃚����s%fO2^J=��h�	pNC|�POA9U�EbAZA2�.��RO�'�R��m�YV��$�$�$�$�ҡ;��>Գ�"C,I+I.I.��Y]�����H/��S�=�z}���B�5i�sP��of��X�[���,|x��Jdp�]�-����6{H¬�0��62K���Ñ�;���I�=�!�j��ے��¨P���H��������e��
Z"Lm���7[s��������m�ä	I͔[�A�R�:h��G��Z)r�W>��:���ȤQUơ�c������o�W�$=͒̬��2^�s�х{��U�f9Ai�9tԧ�֔6�^�<�e��um��f���n�o�8�ל��ßZj��bSoM������8bAJ�K��:���
7Z��uL����e6)��e�f���?|��&��l�0�%v?��R<{-�鹗�u{(ʎK5%�K!ߞ��=	rs_W�(@�X�t�L�G:�ui.���xYd�|$������$��G��%2t�w���[}ur��© u�N}�HC�ƕ�9��ތ.���r�uF��!�ǭ����+�uFΘp��#�f�0ά��i�9W\�=U�;�e����
=T��i����4b+�v��
[n�:=���*������V�ٵ_00ժ���G��(q痆M$����>*\-޼v��i��^�m���f> ^,YwF�]u
��]�>)��/ٴ���I$�]�������a->���F���G�>J>v��ׅf:�裄F��9���D]dQ�t���&LSN:l�4l����l�7�����C��6L+5�[��>(��)��#��%�>�gXlù4��������fq�g��Um��f���(�G32�3UTa�����̷pK�Tu��,�Q���4�]Uc�gJ�P�=��:I�E �8@�i���>�����K0��1�><z}��@����4�����8b��yd���N	n�1�4�M)��O����'���p�}��t���g[� �b�O>����=y�2~��-���g���u4���OI�f�6x��[[i�Y�1��h��C��o����HrH���8r�|i�T��4��t��p L\� �GyW���I~�<pf���}��Ld4 
8s�@�3�6y�.�x����9��/1�Y��Q���6�a^�N���QD��z��MN��MN�I$>��NWӪ��υ�YD	I�;#����>G��H
,Ä��mB�D��a�'[1�D��ӦB�Q�}G������d{! \�j������A��Ԝ��$
Ň	>�����i�t������f��v��O���odu�=�-��çO��ڧD�:|:|xbW�}7M~��׼}8h
�%�g��Y��Ə|(�� �<�D�6G�4�0,�פQͼ*QC2�T�7��#մ�a���iV��Ɛ��_1|i�Eú�d�\�>h��᧷ [t��E�8B7�^�*-<S����}#3с�،Ym����Q�6t�^�[����5=>1|p�]���E��1pӅ1t܍�G���/o,C�I����%��+S�հ.ښ��5��.~��G�U�/��d|r��12�@���emCN�N��iK��;�M����_��߷e 驰K}͠��x�t�<tK���~1|~:b�[$�)�>I����N�**s��-4��9<��i����<)7�w�0���@D$O�2���Si�.��0�9�(����"U��8��=4d)s��I~�)��vO��<8h�;��y��S�Y�@҈ێ?0��ں�����|1ag(�����O���m��e)��:� �js��YMl��ɔW�+p�0��sM�h���&k��'�=F�o6�I��Rոx�T�J�.��Tb�wZp�=�nca�m������&8(�%AU�(�fU>:oq�a�Ó������5��k5n��5W��R�0�S�π����AqÊ=,�|I�	#eys��ǌ,�ZJ�k���K8�׎���}����e�Y��(ی�@AC?r�pKK9__�/�X3�4��t�|��(g�c�}j<-ոT6��Bᳰ/��Nh�1/�����{�>��(����������|1.�|Y��o&hZ��hR�)`���s�On�(��YÅ���/k��\I�Ң�@�oG���Àx���8bG�_'���{
��0ѫ+�4�Sʅ-CU*��dh�
�4{]ue��fQ,ٲ�\|�d�?�m̶J>�,j���f�?hDÄ����ѽ�0�
��8x�H[$83�ѽ��K*m����h�g��`ń ��x�1���8n��Ԏ���F�ᙎ��6h���lvWg�dv�����Ĝ5�Y��>7���QE�4x��%צp��`i�8h�R��K��'$�M퐣4 ����|i�	�<S�����CC�&����C���~����p����=�9Ҹ�h�'_:�����E�D��x��H	�KƟ�:Y� ���M}4 �t�2w��1(p�ݞV����8zʃ��Mh����FOzCƚ1���4���b� 4���ri�΍o^txI��8�<oM�Ym�q&�::uIO3�t����)Æ����a���8pĩ��4��~���h�t�<b�?�f��p`t�!�=����f*w��d���|���d��OL��!���Μ)�o7���G6iF';>�٢G^d��x�gH����4��R��f���Ã��~;;4��D��<CFz��q��2v1��ʹ��Ir�*>��pޕ�<t�w�t�6�J}�RbA�7�����O��x��8��g�8p�<C���[��O�Qb����zn���T�� �!���>�Cq�sBG�F�+,颞��Ym|V\9R+l�Rޞ:_7�O,h�� g	#�s�2��Fcpٺ�G����gV��C6ya��xˎ�5�T�V1"� ڲ�)�۾w�����t>��J{��d4��K:����ύO�O�(ĴŊ(�~�w�>,��A�zY��h�?|��(ޔ��F��"��v�=;O���C����s�[��I7��8~�޵�Hᣧ�m�p��>f��g&�$�>��d;l�zG��F8_�чM�$��(�m�;2韷�Ncnq�͝4t�@C���>4wJ���rPP�����md�ӽL�"�M�,^�M�f�QH���gI4Y��:v�⚸��Q~1{��>�8R8z7��L��v��ӓH������MEF�*c�i
�|��$[�ɇ�
Tp�ʷ�ay��q�t�,��������p��Ak��<x��=�aXU����;�iSK��|p�f�0�=�N�0�К6r�$�T�`�h�M��d�
s�:z�0����(����	+9��y;)�g~�V8h�N���[8I&���BՉ�p��ֶY�f�qs���,�D��zl�7�^,�F�$��x�b��޻�h�F���uS�ϡZ�>��k��q�*�]�tG��̎�,��ܓ	�o\	#�U��V)z���p�̎�����$]�k�1׵��޹e�6�q������?���?���?�ԣZ?_�~���ϳ<q��]'����u�)�������z�_~���Zl����h��c,M'#����J��cp#ȿ��Z,Z �5��!���#��*�����T�e#m�e颻�AZ�J߅5	-
�$�E�LL�(c��u���:�Ɏ���^��y�7�����Z���21��,�7�x��0\K<���ٍ�]-em ��<�m��Ė���1��|�v��ED���ZV\b�y��X�۞�;8�봝tJa�w ѨH9�?l5pkd�/WW[�[���|��~#�Sé��*ku�d1&,��("<�+y,fe�8F�G#.�(���Ԉe1Z��L�يk5�1~����
`�JV��I�/?�r%���eLT�vO���y�ʚn%Ep��=�V�\ؓ�,�x��<�f1Q&6�
q4q�T�9��Ȉ�A���T�tA��)��,�uG����ĥO/�+��Rc5r��+wh��{v�{��Dg�!�F<l�a!��+7j��Px�fI%BPT̄qOV���BK��$�y]W���o���{x`����*�ϷfW�&)QO�V�(a�_n�B3ZzƑI�1rij[ZRDP�QTP�oJ���Mod%��i�5��L��[�c2G�F��4풦�)$���2�M�

�H�1��⭅f3Rį F�f�M�^z`v���4�a�Q��$xf��<0��vd��v�G����We.h��.vu�h���]� -�S��c`�vzf4�鲀F�kV�6$��S)��.�ht��֐m�@G-GoWhz�6����k�9���6"1�7�:яom{��-�S�V�1���R	��Fٶ��.�m�掴S��4�X��`c�mv�6pb�+�Kl7�v頍�撦J�c�D���U3���q�KL�+|a��md4�ĭ���\h��ln:gX��ͼ�����y�����}��7>�u��32I �f�T�b@���k�4���g��������;Q�l}��?>�o��~?O~{����ק�J��1UUQUUQUUQU^��V�^*�mWj��]��Uvګ�UWUU�*��v�ګ�iU_"���UU�Ҫ�Wj�W���U_-*���Uz��v���b������UU�UU�Ҫ����zZ�
�=[���e(V�[c��Օ���+SVI����m%F��-M�6��ͫ��l��Z����m5��i�[�\LUUQUUQUUU�U|�*��UUq���]���iU^��U⭪�mWj��iW�^EUW��U�V�^+J��UUU|��ګ�iU_"��iEU_-*�wv�UqZUWʻU^�UU�UUTWD4kZh�T&���f�F+-lճQ-L+6Sm�jE�)����E�L����$�f�@
��jkZ�CZ�ڪ�J��Wj��iU_*�mU�W�Ҫ�EUUEUUEUW���U|���U�V�^+J��U|��W�Uګj��U|�UWU^��]��Uv��X�����s���V�^*�mUx�jҪ�V�U�ű���jjͽCn,Sr��M��P$�Z�	|��}�>�mU��V�W�����Uz��[Ux�*��iU_,UUŊ��������1U^��V�^+J��U\b��Wj��V�v��X��-*�mUx�j���X�˼����iUU�*��iUx�j��[U��Z��ns��ޡ��j<�i�(ͥ��6�+cy��Xʭ�1���[f�M�Slt�-���92���!Z�fݭ���m�ئ��Jo�������l�KD������_���!�lz}{�}ϣ��vv}ݞ]'�}��"'DDp� �"P��<"`��x����A
A�x؛6"X�8'D���0L�6`�"pL<t؂"&�N����Hl�b"pDL,D�N	�,K͝6AH&�DO�Mp��B"pDL�0O:pN	fĄ6%$,M�A�`�H"X�N�'D�6Q�x���&$��"%�pD���&	�p��AA4h`�č�����t�j8�,���n7aZH�hr0�^ڌ��<��U�\��ѹ�=�Zz;9��'�4�}��ns�cy�[�V�^��/U����&�����lu��~��$�p|ն4�wI��^;a�[�-1/�s�\��0���c{$l�ŝ�c��U�9+�G�VG��m��M�$$��
Q�s��b�n���o9�M�ۡ���]Ñr-j�51�V:Krҡ��Z�=�Ƶ�����g��{���2�/�4�� rw8M��M1�6�<�	<k����<z;*���%MKP �
����%(�]��������|�`F�}�mӃ�k#��ձ��m5�ݞ��T�n���iN�v�8�:�k�3mw4u�y�E��ۏm���_����ag��x��ٷ�~����nA����7;٘���R��
�\�Z�&�&8�;Y7i�_�Wҟ���wn�s�E"��7���SlrB͝��t2A��=�<v�z�}v�j��U�;�MEu��6�q�vG�l��=������p>"}���wL:y��r��Gmڪ4s�N_k!���n��rq�qcJK�C��6�%uΤ����M�5�X�6�s����ݻW3��L�g�2k�hw�ۮ��t���l�9㧻�q]�꽏]�����.s�g�a���U�w^yۮk,��n���t��Z:�@�J	�H�E1�Ex�k��cD]�ltl��%|�0�T����4�nk�۝l`���y@�6�v����]ـ%��s�ö�nUG�W5� -�)\��֌����F��鋮G�򞶭�[���~����j�tr72>����e`q%�y
sqּ[v�Pp���Z�N�՛B=���Rem3�������d:�8]�*^c����CV:��;f��9?\X��K�O1�cu��3玻�&7n����5X�R������U�bb���� %=�GP���,|0N�6�w����L^7kz�Ǚ�7 �;ѷ%�lp:0n�n��<k;�v�ý`�����nͺ@�iOY�۶s����=��tS���7e܆��ëm��"�=v�����{�IG�%�����8ۇ
n�p�+q#��f^�v�4�R�l�B<gBn�7]�>q������N��e2�G��D"Dm��Aj��17�?}�����<������mD��K�k�w����0B���*�����Jmۊ���g{r�v4s�u�]�>^����]IY��^�8,�e|��P����1��m�C�.59�	��.����n+�n��c�uq֑���F6���)�]�_n�I�n6̣����햶�x��kwGc��øv��ۿ%�>���tg\q�}q���hM��nb �����ks\<u�v�$�����lͷlGA(�:���d��e lq���:�e,�����"osX]���m�(����:�Ư�� �^-ny��D��4b�ݪ�K�.���7&�-n*�z꓂�k�ۍ��Y;$�k]p<���rv�T�{e��v�F}v��Nr�gd4��x�:����8��m�ػN�q�;pvg����l�ǲ8i�nI󣱎��k���[V���Y�.;=���1��#g=�lwlv��`�z��v��r�=�m�s�7��#���	�9ʪ#�d�8��]��w�u���O�.�n���n8��]�l�܆�.��+^w�b1���vݷA�=z��d��*kv�թ�b������;�k��ύ �{����.�|�g�u��㎰����ש��6Ƌ�-����,�ɷ�r�tcu�RB�����j��%�_���j�7g��n�b�DG�jR���z��k��U1��D�r������]b��V���Ⱌ�ͻk'�V�b�'(�YOQ����]�ܯ��K��s�;\b���:�l$
[q��" �����������EV���� ֍.�W�,UU�Un��πѭ]���X������۟ֵ�.�W�,UU�Un���� 0H a�0(��0�0L8'�ن��g��'��R�\&���ǁYg��΃m&���QU�[��L��v�ݭ�� t�t���v��v�a����dw�i�n�k<[<qy�u���5�U�����l.0�Yr�����N��z��f7vD�a86�x���Z���0cͻJ�^.x�WIōz�Nrۋ{��e��d��ڛlh�֮��Y��>�ύ��	�O	��Ŷ�(6���i�%I���D@'X���L��Jh��w�u��|K=m/rw�E.5�v�tr��r�y�W���ݱ+@�48�"B�ESU0"����s�G'yU���t���L]�n�'uƞ�Op��;l;S�F�8㞞,�������$�Y��7�A�7��yQ��7��g���^%�,n��,�vƦI$���C�L��8�LB��.�v]vK-I����+oiZ�t�$�KuV��0b�B����nm��FDP9k�,9uUu��[Kcn��B:ijv��x�IuT,���xA�V�<F��GN8�x�ׇLj��塢��U���m����^<e�I#�����_b�1�sɱ�j45��f��#�
P=G�#��-ҳ����F·�rr�y-Ǘ>�h�/#���V1p��ъ_��ޣˑZ���類0�
?<a�l�ㆎ8X���a����$��h�婡§Z � .���_.��D�h��TyF٦/�qW�77N�ܻ������:��m�	���躟0��i�yj�)����6�%�ԒI�Uj��Ay��7yѮ�?�^@.�E"ѯ�l�V���%�o\(�m���p͜e���o�D�P��(�Fx���D�0N��0���.]ʆ�|. M�1ǔ�LKLZ*$ŬVh 

	�V�:,��ߌ��65���c���=��F��h�����m�qUi
�6yf��#��� ��b_�)bJڗt5+��r��|�*�n+6�o�7��U"��h�2�F��1���i��gW9,�K��Mm=��m8�T�OGL�6���-+1W��U<`��S�(��<l�f	�0L����A,1��0�P�t-�P:�����L~ z�ƹ�����]Q{����&�,W�s*�r���������sugnOh{��Y�	�)t����PT�UVMdǕj�����;�؜�=ݮ�8ַ��q�(�o!�7���ӆQp8yt��lQ�R���+t�)��;��R����e(�f0؈�&	��Q���z�k��\2�R�e���Xʀ�n��,b�1ƣ�ѕFख�ا�9i��J�7f���HGX�  ��{ǃ��"��.�"�-9�-�6(Z�\��X�v�2�VvK�v3k7:ҹ֝�s�;8ƫ7K�(t��'�o$ZƖ�krg#�L��T>%P]E���8դ��ݥ����0H(5�d&HL��8l�=����X�wJ���!��Bb�j9��Y��և�T4XO���P gQ� �Q5�64��<������4�ki��-�/#,<��7�Z�mDoV1�ڼS6�=��i��x��{��<����l1Fv��j��Ywyc|�	xp��]/E�Nk��ΐ����'DD�0N��0���]��(�i�Զ`�g�  ���B\E#��2�Sc�q��j�zQn�S�l�*킦k�8u]e�ň�����JG	���r�
�����<������zp��Q)�M��C��kgQ���ΣH�T0k�qjh��eB^80����[ӫ�@`�8l�Ϗ�舘&6p���e*t��T���EG$�G6  ���>h�6��-�a�8��^ �^�n=����4g���m���8h����K�GWN���-zm�D�3��ӄ1
�f?7V~�m�E̶la��j#QҖ��T=�1\#e��Ѣ�m�-#d:�`֑��=�t=��[4��F�Q�k�"���`y��Bύ�l�g���DD�0豠�����AÆ9��Z��Ƞ��)�$�F�W�C4��1.M3��6C��x�^�j�kF�zȝK�,��k�k��wb4^�� 8"֍�m���y�-V�(���4�Xj���lz�[6.�pﮤnH9j��6=�8�l��0��\�|}tsn��cx����ma�-��f��B��٤�e(�gK0�:"&	�L<<C�l�6�y��e�(T\|g$�ww3���D��N��X�b��v���S�p�I"���/
���&C:�7{�"���IRWR�/���tY��n(���cUOUTܼYD�.�ŵ�6���MYjj�)��#��l�P;JM�==j�1�.!��gXV0\���_0��Wnʔ���=�[cm�����Υב@r؄��W@ 7il!HZ]P�4����[͢�m���t�����m4�14Yè��cmYkH��Ze��qDD(�EC�6��^6��Q\��
g�7O��ci�1��ʤo�t�t�j�Ic���Iӳ���,DN���a���7|���U]���b�c@� \�gZ�;Q����h�j��GC�n����e1x�3��!�m��t�iF�� uES�лF���0�5Ӧ61�qQ*E�K�9��ۇCA����gWV�?c[��5��}{���ҟ*�9�K�/ZUbx�� Y�2/."�(�[,���WM��:Y���i���=/R������Ylf�O��0����0�BN�{���d�#�aD��<2>���0�$xFa0xQ0��f�#x?��a��ǃ����3�`�a3l�koL��5�:\tCEf`�c��3f0�Ҍ��l��0~!�I�|M$��>"O��>7�,��N�����x<,°{0��>�������D�t2�G�>�L���<��D���͏p�|?�>�Y�X�>#>!��x�>0�>�L��@x6a0xQ�`�{0�<<Ca�
0�M��le��	��<,��83
���'�w�IorwRޓ�q=������x�P�px۱��o#�x�x~���t�<�&�#0�>YXdz&�&鑼����0�ofc42��3#L��#lk���3��`3C,g��2���J�-���A����껆�ُƚ)C� ��&��Y��0JK���(B��Ô�]Un�d�P��
��XVI �i��U��KcG5��³E9mq�o-�����L��Wٓ���A%�����Kn����)P���7k)d:k�c��0�Q���{�7�Y��:�H�S�n,[�L���y���t�
����9�5*���m �߿>��>�?9�fVfffs{ު��vD$����{���ޞ������UU{:�K�����}�iW��>>�﷽��h�f^fg�uZW��gp�̪�����ӥ(�gO�����a���(��jj����DA���U�	��TmY��4(���m.�uG��F�2�%����q	�&�k(vE6VrwoU����ߎ%V��ἐ���3���I�Ǝ0aHb�ҡ�hb�F�����0q:�[[�#�c��	���s�>�!�N�w�<"L���A�TGZ]��l�G��F�5�(�m���ny�ɠ��@�·^�)���Ige�8�D��g�*J���+F�iq4�g���A>��.oZ�>b�����h1��"1)�H�CXD�f��x���>>6t�ç<0�`ņ�=6���P�BH�1���b�����Ax4�R��E3�!��(�Ĵ�����i�ZL<���������[h횳sH�"F�!%äF�� ��d:yR>ia��I��{Cjܹ-%�N�ںEH�:1iTDi�Z�f�N�G���s,ݻ����Y�='w\��i�5U^=UI�0Dt����#�E%9;��RL`�#�"�,F�Cѻ `��o�]U�x�X���Ĭdf��<2:8[G��cM0���=�JB����t�.�l40�B�x�>����0D釃��x����z����|�Sׅ�|\�6�J�\׶SZ\�����,L�X= �u���<�H$�HnU�Iy�-X��[��j��P�l��K��MUO2��\��7y��ݙr�{�|�#�UX�a��,^�Z����n�Pc��N�3dҹDn�ڵiv0f���U�i���2�'G!S�B��� ���"4�_=��h�:�4�1`Fb����.����m�GZ�Dw17|��7ڸ�6�{'i;#,`�	�DxaHa��i���=#���YN�ol�����v�5�q���qs�:����Ȃ0��^�5�V�����ȅ��rCDCB���-E���xi(�D�i���5�����Y�O}�Ǚ̷���yGw�՝7;OZ�[r�D����r	��6q�5�
�V�e��
�W���
�GXSм�V�zө��}GH�����ų4�Ac��Tc�
��h���CGf�x�a������"`�ӧ�!�
K�o{�ʗp�*�Zof�	!$$�!�7���	���Kd��{Gi���g}������c>8t���B�H.:	�$�r��d&�L m�=ߤ�Pe��4���4&��p��7i�-�����yOHt��&&���C<11\B}dH�h80cXB�)Z���W���4�A���\o���ƯZ�E�q6Z)��,3���k�@�<���[u����m����5���|�E�dD44�M����ZaP�pL[C<r�4������m�3�SV2��4�a�D-%c��)+@���l��5l4uE���l�a�����舘"tÁÃ0��I�U���ݏ.�^��I	!$0�68+�_j�0�)h���>�DRe��|D8��^s��t��n��;����j�m(��(0^#����a]�u~�M�|�]0����l�օ��ui|�.�(0�CH��cK�B5���2l�-��X���ې�)����Sy��֯�J�J�
C>LA)DJ�A���1Jw�x��ێm�;|:R=;���l�͌/dM��� �[p�R҇Ʌ����@��������6P2֪�C�)D�6c�Ɇ�#�ꘚ���`��.����XКcR��Q�U$� ��)/����0�G�~?��<x���Μ��+��+�2�t>2�nS����^�eJ7P�BHb�DP�13��
M�%]G:���=��u�;���)с���a^y#$#�rP>{�r���q5�f�P�������9l���os�v��Y����.!����$�L��p�cf�ێJ,i4���*"���h��A�y4R,�)H��KC<��������B�6B�I���D�����-�G�Qq�;�N���Z
C\��z�D�aHD�`�k'S�r++:G-�gI��Q
��E�i3ْ��6�5�zF�V3Q�R�H�dM3�6�[[,f͔aFh����ǎ�<l�����0���ے����z�i�1/������ۜZ��կ��ʸj�J�\��Z4�H"�H9����R��TC��6 �	 �C�������e�
�TL�
�FʣJ�X&P�����@�>��qV�$�dЦ��H�Yë��h�g��3��:��7B�-3+TPj�uØkm��l�AS����z}��
H*��:.kD%T\<��`������h�K��cD��4�Y���qR���l�HK�s�K�#E4h�1����PB F���#0�l���\	�s򀢸���1*(�p�CJ�4D��"�O%Tt�US:h�I��h[C8��o��Ж�"�iu��j"�͛Ú7j�0��^d�841���G"3G�������*&�΢B"���qL���j�y�C0c�l���+B�֡$]E���q4[!�����
���V�2�4��H��6�5���:l������tDL�`a�<|x��������rA�ի�{�E���I	!$0�������H� X�C�E�l`1q6EH�MuN�V#��
G��h�h��ե��il��[F���xE�h-�����'������@�JƲ��*E���ilta�0�h��ZF#h�`b��}��J�.~��Ņ�P��~���:����R��ċ�D�ub��#k1'H�J5�Ty����'E��Pq@cS�e#�\C
"2��R�)����y�4�þ�}�X��Ə#bf���=ҫ
 l�<lO���"`��<t:tg80ٌ�3��n�lZ�"���(֨��$$��a�����K��&�޵�w�u��_i(���È��Da����ZE)yj֒�*A��"�t� �DQY�R8R(�����)O�H޾��Թtᣈf(0��6�t�A1ƚ#MT���,��uQѪ�kk�B45��:0�;]E)��"�����J��-s�Ê�
|�W�cm�J^{VU�"_7$������J�yZ��ϑ�a��)������m�B�ц��v<�È�PXQT����kf�6���V�qb7ih4pgNt؉����0DO	�����h�U1�8� O�2K�fŧ��N8�0�᭬��Q���m�GQ��$�a�F�n+Cd��Q-�9ϟ]UU��f9Pe��ϐ�9����H�H�ޒ��I��E��C%�)�o:����Ĩ`p�E�8JDEb>E-&���P}kj��6��F��QdE���J�Lj$�����mF�U�Gv�1h�oj0�0��/��/T��b�ip��]>��0�� ������X��6�l�SO�>�R�DL<4�!��[zU4� Q���j�J�tg�2�Y�0��X�c�F��<*<&ä���	�f�O��D��z7���xx��!�	���#��l�ݐ�f&ى�`��\.6adVa
0��`�<�6a��?��^��XD�	G�I�|D�I�|D�����t|���xa,�`�a0f���x20��Ƀ0�0f��o�x{��v>cpÄ6<��t�2�&�������>0�G����#0�J0�<�&<���N�78=�c�D4L4F;L|U��ӎWÚ|8��I��R���Ã�ٍ����
��x�3�����ȗQ)�Xa_�$��J+�	���
�ل������xx�!�	�����3omb�ܞ�^��I�]8�|��\'��^i<b9��-.���X��R�tn�e�i�Y���k(b����QgL���e�C8&������9�&�ե;YƖ�� �Tv�w?1Xg���Ku%�����	ؗ�*���4-{�ìeZki�L̷z�֡dl��Om��ѨU���:"fg.�;h���o(儖Ob���^w�(L�-X�\�7@�:٬1
닑���!�_�*��fk�
�����^��>և�Zh�[��a��鿷{p�{�F�̲��s�"����̓J�3gUˡ��m"M�r���e5�\o&��hR��ϕ�߯������s�.��[5��2���G�c�	�J��6��K	�\��&���E�Єu�"	�vm��&*t���nI�8
Ǻ��R�hH�7�m&�	�|�y>|����������Uz��}�����C33/3>���U^�~��^��ffe�g�qWj�Պ�˻������Ͼ��W���w� 0!���l�>0DC�`a�<|x��h�vʆ�{��Z���3BK�[��t��F1��Z�y5t�=��ݮt�zx_H�j�ɴ�&8�n��g��n� �b�;��=�X15U-�P;jBU
5Ru�=��w���|�+��5?���q�-�ܭk���n�z�Şg������܃���Zݞ��m�ۡ4�l�xȼ�,��_A�ݖ6�=F�1��ȇ��ˋ�W���'_s�j�*���`{eTJF�iЎ�5]M��v��c�غ뵸�C�5ej�*����FmOwϑkoSoc���Lш�ݳ�w`��$��x�3^ɫ.�ஹ/-d���zW,\Y�;t�q��g~���m��`*�3u�m�4�t��KF7J7j����W�_�	�9���`[" ��y#/�ьcĚ'^�p0o���nS2��:w��.��9�V����O;4�w�4�Sn��6�%+�woB��u+��Ϋ�t��.�mS�}�y��4�H�;���8�2g<��̦�{p����H��K�����)5'oKoj�B�W��)R�6���N�Ǝ"��}ځ��j�T�&��RK:{��9h(`����g�#�m�j4|�_�XhhP-(����V��DR;�1A��&w��*r��|a�F�#��6�c:Qj�6*-k��m�|04&ks�GzE���":"����
K�7E#�m�m�7&[~��G�j�ZA�s���MD����.�*Q�����\����Iʡ`�(Bnl��Z�y���h����}����lc"��� xa�>�:�7��RZ!�[�C>8{��4C(���Ə��O�L�a #�̄�@��~q�q�`q4C�5i�TGưlce���((a���4�Ç��6��/v�P�I}ϫ�0�Ld������3W8�-�!��;=cZ����+:6c�=�h�N(yPE�2��.#��40�>���$�C�"��M4���~Z(�j* 2�8V��5cYOKE���1l`��%QN�DL�)�[i�^Ȼ��z�/�L"1��"c
E�!��o���Ŕ��{ll�y3�C8�מ��k��C
�(5�H��I�6yr���A�#EPb!��n�!��qX�"*E$���4C��Q�|l�ǎ��C�`a�<|x��r��RMHD򼈏 
	F�7���͇1�chK����{��첊7�ޮ&�|����H�8Xx�`B�*���ik�C�`Ɛղ�"� ��EhqZ�G��[I0��ҲHh�X�j�	��H܌�Ң)����8��� hb)�4>(y�G
E1�E)$#DaC0{����H�O^%"
i��7���D�f��\ �(�-��R����|�ȉh�ޖu<g�z�Mӻ���v��]	h� C�h�%���m��u�XѠ�9�� �<3L60zlq"��Y��i�M<�G����mJ��G����k�I$���#�Mx�l��/��H�8>*Vl숱�[�Yj�#E�Z5H�4P0�eabl���������c$<'C�Fpف�r���Cw��q��"�ŷ��<9��:޶����D|i8�0�1S-DmZ��1��hf��)�M+accX[a�� ���Ԕ�-	$� ^�5S����R�<xs:�γ�� ��Q&�t�T�������4RX4l� k�#d�(���ࡡ�E�A��"�Q{�V�-TRj*s��i6y\m>��8ےqsK��P��DΡ��T����:v��,���;.���Y�F5�#hf�&0�h���6�Yh�2x���"�P`�Ë��G��DD ҳF�E@���!gK>6"p�~:|"`�$<&���0�λ���Aqԣ�^��di
L���R��y9��R����֥7nKm��	ɢ�ʣ�� �1�Q�B�S�SׇՈ�z]�� �R��՛�/�ۼ�t�Κ�����Ϋ���Mu3}�{lT�l���BkGt�Ȏ����>�,t�˥��y6�˸g;h؆�"c�!µ)[��hZI��I7�[�^n�;����
:�{��w�������C����-�Edw�n�Y���[�v@|�Q�h��Z��"�wI1�҃����Z,MDTƭ���E��Ӣ�c|$����#��(�Hh�G�{,�<}�0cp���\��Ξ�yG���N'�c��ZC'�"hߑJ��lb%Ȗ��^�㖍�6�>ҢP`ն��Ým�l����SC@��2'������y�?��J���M�j\&�é�t�"ъ��6Db���*x4��dT��{�t��ʹ�h��(<`�>4YҎ�>?>>�!�00�:|��~��Z��Z�R�Nc�$б_�R�Ůh�-��T0=�b4Xw[nR�np�[{�g4n�P��BC7��HX���W�gW�D,�9#�p��k�64�٥H�1X�ha["��C603<8�Zۤw���6����:"*]����ͥ܉�)��H�;s;�8�Χu�5�RP�o�]��/[��}Gd�]]�=�f�ޝ;�^~F-�|��0�`�D)2%��LdqC��)�r�ш����@c�C4��=�>MD{gSև�伭������+`t�)@j��R��@��8Y�g�>>8~?>>�!�00�]_�>^��"��a� �1�bM0&f7$�
��B)D[E����f�Rk�60�@���Z4�)�>"�ҾD��&�C��)us��!�Z4����iU�F��a�i�a�4qb��p�F2��*	Ɨ�A ��#N�����\�st�.�՗r��8��N�F��U�6��'�jaM9���|sx
W�����i1��9UkZQ/����(�T-0 b�"41P��5�4W����Æ��B����m���%1~�4D���?�R#�v������oZ$7&�j���v�y�V���
G��XZ^P�꾔X֑�T�R!��������������͌ t��ŉf>?>>�!�04h#��mz?D�蘕U=UTg�q2]�sM�1�I�<BM���13����4.����`�ѣEWU�����jcmwP�n:��� ���Ĺe�z߃�������{�V�ZQ�E��ɌtY�l`�1A���q�h�
�h��dGP��բi��c@B��H��ѫ!���3�g��"\I�DBc9~;��r��Q��D��PAA����R9�h�<�š��E$��A-�R���=h(am	�,��Q�3�Ȉ���<n�Ҥ�{�P��G8�8�82�9H�����*E����K0��b~8~?>>�!�00��~kq�깖[ʭ�5z�:rMQ��앙�)ۖ
'�Ria�J*�H��k%�z� ˽�� �"�(����ߴ���A�5��t*WF�m�{F�nt�LR���m'[a�l����7y9{34����cF�ז0
�霡�u�o�s�y�
�5cH��V�]���7���a����?seӕ�5E����39��|�A�54C�Hi���"ac�����Q�����0m�/��4ha�����Yh,f�G�aW�Xұ��0�hi��{�uF�wH�a��	��0�jBh��u<�`m0����F��������-�{8�8�������фץ�!���&�к0����A���x�:Q�"1D,iB���p�M%����ǾY�ӀҲD�FT0��=�����n�=�����L�UU(��g��%�`��gi�8��[u�㶛�7Z�Ԝ"悒�dL��h�H�X�S�eu���g�6Y�0��O<3���N�ს�m�$F#�J$�y��v&��V=��1��Y�n 晿o�#�8Y�)+�t����uX�����)<4�3����m����<R)��w^�t��c�r�mxdh�Ϊ�l���h�������"��X1�1�*��)/+�#e.,�۴Y�(���,a���3��4�ҳ�r���Z�85<b�j�L"��)q�R�%mD0�8Du*������ݻ��K�*�QɎ��ݭ5d֬��,<�l� ε�5ᣩ2��\��b����vil���DG��)V��#�0ᡣ��CH�'d)��8Xi1�l���-#l,a���AcGQ|74�X���mg�%Z�Ό0f�Y�-!�hv?�X�xFa0xTxe<&���xh�B`ل�#�
���a0xz<��<L!�n8M���&��x�x1�bm���ɉ��f���.6��+0���j�!�6a���cu��L!�	G�O�|D���c�	���a�Y�X���	�������0x>��ǃ!���F��h�<m��`����<�8>E���px=�M��E�f�+�0}0�XY<<4H<!��(���	��0����'�p�lvn7c��=�!e&<(������&<�xlf���ۣ#����l����3��FFύG�S�`�t���ᢠ�c0�dtaX<�&G��"���&�ht<N��I�^�I����F�����n���/��v=������?%�:YBʢѧgߍ�#�d��jt���1�N�T+4:�i�}q�ZV�jaݺO;*g�����T�y#m��xX�nσŤ�L�p�Z�mV��n����⹙n�^�k5��v��'U̘��������Q�U����;��V��$��N�]zvbF���s�v ��u)w���{���HZCBp��Qݾ����Ͼ}����Uڪ�b�r���339��֪ګ�io�]�fffg3>��[Ux�-�˿�Y������UmUⴷ�.��Xa,��,�>>D�ad�R���C�6�4%��q�������Q���/��G�DKcGȲ��T�*�y�#FώS�>!J���Z:Q�"�5��CW��͛U��Ѱڨk�1݁у�����Y��uZ�t���	;��Z湷�n�d�Qg��EE*�gtvX�;�ös:G���7#�<��[�ʮۺ]���z�l4М�uY�1�^��4���+��C��--g�e)N�if��K�֬�*�ѝ1@�u���'j�n6�P��|6R\V<��5���>g�u|r�ȫ�Z+���z5�u�ܐq�V@�4��!�1��8p���	������0DO	��0|
�C!Ye��ʤ �z�A$��e����CG����9F�l����Ͷ٪[hwf�?��FsĪ�S�7	]��%�o7x7�C��n���d�b���/���Pk{m�H�K���Y�(PV�q�q��lkC�G�U���DG-(cK�MDlh�4\�h�G���4�c"6M"���5�W۪����/{�t�SZ{���#D*�CG0{T+}H�G�b��h�[c���#��4��R5�4��Z/G�m�(Ǎ�-F�nцHf�΢?�4��,�gN�Y�Ο<|l�0DO	�����>�%d�ݓ' ����`A��w[$z^0*��X�U��p�y�+�X:��Y�Mcf���&�k�}֛i��x�L�Ɲ�}��l�]Z�lS4��ث�g�-\:����S������ة�9:ּ���{+	�ѓ<Z�('�\%XS�v�Hu�Ӳ$i���z������DFƎ���ZCCD45���|F�+G����{L=:�l�1����Ũ.�4�D��R4QGM��a���7Ӷ�#x2��M�F"ʠ����هd�(u$*S���*qohh�e#�����4+������G�=�v���y��;%c��#_P�`6��4arQM��|��c3�0m7���>�DÈ�Z��c�Jpg��**�O��YA%��us�|b(����ٖm�A��EYe-�"5��1��!��Ŗ7���(�G�������|"xL0�����	H�Kl
���rBHI�۲R�g�cL�Z0�� 1�6��*:�l:xm��kf�.#o#��_y��le�j�M�䍷">Z^�iDip��F�,llgu��lg�/�����h�kG�j���M��7�5����9�m4H�f�l��|J�������܈�����U}]M⸵{hȅsjɋ��[���Ƀپcx��˩I�̈˲'�ip�ȅ�c9��ζ6iZ�,[�ۈ��t�3ad6Bϊ8Q�f>0�x�ǎ::3���2F�7UT�!|��n��e4��Zm��m�hGo����Tk�|��Z��>5������@P�tk��"��7��Q��h��8��{���\D���um|PpgQ�EC1DP�F�����y%�<�:��xĺ�*�����m��OR4�iR�C~}V�������H���z�C8W�,]:R�cG�#Hj�s�����bkaD�E����)X��i3gk}��W=z�]��֓8��:�|%#Kql�Q��(Z��j�aIZ,�}�,4��p�GJ:l�����0�<t:tgs�B����;�I	!$Dh��_Dg���Z1x�@�3ܦN��4����\-AΨZ�i5�e�i�?�*��vDlb�mDDip�V���۳k��e�KԊ1�c��*4�
i�#ƇH�6�T���H���I�)b, ��f}��Ɋ�\K�D=���r��chÇ"���x����È�c;g��"��x�:��*�"!�戸�J� @��!�<Q���p�<a��::3��z���,�}'Z�H�J�Z�KF�ӻ�n<��nf��z�_�߃��8���3b˾[����t�)�X��p�K�ws{2R	��&�x���P�*,d�h�;2B�n��f�����q^) ȠAip�Xf�Q�AmiV,e��A��}ۗ���]½^�h��J�=���nj��L�<y5�գY\_42"#��}�1�A��a�C�p�G<��FѰf��KC5���.���UP�J��E��h�\E�͞V3a�.ycE#��r����c����UGYLl���ּx63䗈�;����*�=c��(���sDq�����n�M�Nۤ��"Κ�=���岑��ƴ��H��D�
(��0���<|p�<a��::3��x�5�SΪj"�ab
�Zj�@����BHIb�,��V��͟l������h�zFա�S�E�3kw���6l҈�;�q�(p�Qk��x}[:d0��޿���k�7��,�m�ۤx �3Kʑ�ER��I��)�HOj�4Ə��2�j4$)쉛<n���K���|kM�P��)h��{��΢43�C�E�^���0�Ȗ��䊣����@ᡔh�p�����a�<p���ќ
��9m��6�i��x��&�ܵ�kj�3l43Z4�MZ�m��)X�d�^r-h疑h��E#��A�F�/�v31&�X����ߣ����s��I�ͦ�lV
�֩��:5`@��Dg"�Z�[�|%q�4�DQlzoJ���#�l�h���E���ã6Q�4b�i��P��Gڔ�ٻXxV3j0E��;>eCt�$p�8������ȥ�R A���F�F��h(,��t�0�FϏÆa�0�����<���	Qgų�F֚p��s�8�`)ǹ���n:&z�$$��f�&4a�YK6�V*�!���((g���V�e�Z��]�vH���q�5����P�8�c@�V�fR!��CG���Qq��a�X��������p`���ޑ��l(cE�߲��uwQ5%K<�N��R:yd_Y��t�0�4������c3>^6����D�T/7K����CYCގq�"ȅ\���Fl�>"��3F���6Y	�c���0�����ǃ��FS�a�`�xp�7��0��"�70�p����/t�����{극=�^��e��Fʹ$��F����f!�8a t�1�f���0g�!���a���a�txt�8K&l��Ѳ`�xt�<Gc�fF�D�`�x<�I�0~0����fهJZ�	���>Ơ�l�t�e�0x<0��va��C	��D0�0�tx3G��0�t��&��Ȱ�4K��	e���l�n� ��$�I<�弮/��	�����5�����|>������od���S����|O'����|F?����L4C�ÆSx?C������4A����`��M��`5�c���33�e(pa��y����B�?���VmjY'_���*K5�6�fm]���@��/�wv�Re(�0��y%7Y/N|]�鼸}�2��G�B���=ٛs(U!Z��E��"�({L�n��J����AݬB�R���z��8���7 W����F����9�3	�.59�F�aP%�㠛�]O�\�T�ֻ���(����4���5͛�.\Tx��nT}�.��E�:w[�9�Ԏ��#��ǅ��wUUJ�5(�G7c5�`�()�(p�bI�8uunǛT�R$t�niz���|\e���8EDKD��NH��d>ղ��;�ѧ\h�d�I����xy�Fh�J��)[����]r0������"54��+,<zXۣ���*z}MQ^��+�����Z[��^fffw>�j���U�w�/��ffgsﶪ�U�]�r��fffw>�j��[U�w�/����afafp��0��aÁÃ6m��%l�M���3�%{�X*�u44*�P滭��U��qQ4;WQOE��v�����'t{J0q�f�j�ۗ���<&���?m&w�z�lgK�r��ܠ;u�m��y_qv����i�X�@�E��gy�K�Q�����ajc�ɀ蔕DQ�Rq\���T����`�^Z�v�-���N���lolK�h��{3�����.��4Rk�2[m���G���=��v���!X�헷��<n[��}�n�`>O=�9���v�n}s���[nx�h<2S��[s�&8;tq����+�zݩ�඗��Uwŭ��T�P׶��T���v�Վ�x���i9�:��=�F��/�-Gl.�I�>�����8���}zF��,�%��:r�\͡�W��ո�Yp��Åb�ʨ��!KpQ<���ܮf�G|)ѷ�i�]ǜv���V�ry,Yv��j2 [4�yt��'��Vsw�9�;��v��w}%u����E�.*4f֚�i�e�K9<qumC���-�ёy5��>��rHQk��G�P_6���"�/��Ï��hgʑ
S��B�c2����MZAC=��D^6��؛#hi�è�2�HBp֩���&$���iϟ�����IWQf+S,L��>�	>��xy�[_\)>43�ҊOE����p843��,�g4|p��x�8p8pf͜�GUTl�#�4�����DA�*P�ӈkB�F�O�(d�S}^]8�-t(g�ߩ�T���<�mS�DD��y��3ˀ�i4�k�A�gɗa|7����H��4����(@,괄� �B��}T�4�UI�5�^<z�s��^8t1��s�Z:������yY�p�>��Ƞ1�/�-�E��a�����gK0�4|pÆa�0�����!p�d�\��UB���I	!$D=��m�,��6�����;#3z�H��G���k��pϑ���"�����$�^=�p�j|��{�l��,  F��B G
E9���߫3+�2��q�M���U�[�X�wc|	
� ?���-iY�Z4�1����N3Â��>Z<��4�c5�B�Un�
�]��R���#�#�>���A�p�|ǋCJ4�'���ƶ2�CKA3Ş,���Ə�0�a��FTg�6&�ʱղT��MBHI	" �i܎89Hh�Ťp���������<4b��b(8�0�����t�8�T��0�m��j������{���+�h�#I��g�@�zZF�5@�|ͯ�|>[��/6�t�|�X��~�ݎ�cov�����s;���]G��Y�#E�k��x"�c6�>����+L�%���h�3�3��[]���g��ೃ,���,�p��x�8p8pf�o���*���U�v�K/*�rQ+*#Jl�S	���� �i8V�j����p$�#���CG�2%?O���X��_��'���*���<� �Z���-U�5������_3��$9I{��Q�
��s���ۍ�>�F���W;�`b�u��;�.ä]3�F�1�]�i�@��-�EX���ER�.!���Z6���c3C_E�;��Dp�x, ʹp���lltmquE1wT���.ڭ��:�`\,��C���q�#t=�&���d[_p����:h�Q�M�Dt�o���^F��)Qe�����V|�
3�UXW̪5�r�ݕWr%uv�i�<mG�4O!��ب�1��Dg�ض�c!	TIC��!��ٺ)F#�mR@��t���,��_��0��x�����/�v��n��J�TT�#�u��m��&�b��KC<hZ�1�F�w�F�����h�+�{��g�g�~�쟤�j�m�����#�VGGM1���!�<Z4�i�鯛�iWG�p�h�4�Z�=��E���q���!�V��N�
n�Fd�I��0��r��I��586ứ�3��lk�ƔF�+�մ��Ó�˥�t۳f��+ž28��m2p���^ӳ��PΖ|Y��0�g�a��0� ����f��.Ih�dQz?�a$$��e�\�H�Bt4/��t�w��h60�p��p(f����G�67��ϳ�Q5�}m6�1T�.*�UBBӜs���b��3�4p��Ӂ�G?� >��"󞒑���#G*<�u��Blg`P�,<����c8����AC���-�h頡�효S�UB��ӈ�����������4�!���K�V���N7H�4hf4Y��0���a�<p�p�͒�M� 1�b�3��m��m�i�Z,�Jpi���0aC"���A���w��T3���4�g���j���uui��A���!_Z[E�����<O��41���l��<�"-�����Ep�8�,� pg��2Wj��D-�U�g���,m'�||�G(�a]G����<t�h��h�����[g���l62Z!���443gJ4p���>8a�0���}4�6���L��9S'
��h��ͷF9���6a����H�0�DAY-���i�A%�����[)%ܯAU�e4/3t!��]����
�WSb4)R����������Tf�a�+g6����Ey�Ó��$80�*v�����ZԎ����e����{f�u�v���[���+��E���yEg�M����_$��X͢y�f1y�83�H���xz����8�l����������!�~�Ã8+Gm-#X�"q��6x�A���,�ɳF�@�I���|�{�y�&�~7A��˲YQ�]���᳅%�8Z�iE��ӨF`�P�@ʁ�]&y.�f��:Y���8a�0���Zh�3�1QS#id?E�p�V�R�s��BH�2��4��
ֆ�aM�
[Vy8��.���>I$����}v�Ƹ�/��<��3��,��#����� �Ps�I)h��A�4��#�KH�:������2�m ��M%"�*�w٠���;L4��f��4b(�-���a�����q��Gz���p�c�����e�漞�H���8xV{[�lK6l�>,�Y��""lDD���b�DK:"'�DO	ӂp��AA<"l�bYB%���ĉ�<��0�`�&	�0LDL<'�"!B`�(DL<lA	�,D�"'��'�	ât��� �6""xD��(DK�a�(�:'���bY�6%HFM � �� �� �"Q���(��g�:a�:Q��C0�0ن<'N	�AA�0��{*�N7�1glvv?��1D^k���R�6�FFN1��J8�]>�B���9�[��`좺�����,V��D�:X�mU��Y�/ r#�u� ���.�tA�[�u�(fK�]��D�k��z��ǭ1&t�8��zN�P��7�#/��dS�z��n��׽)fN�;^Z��4�p5("�賩r��S�Gaဃw�t򳌙�(��w|�F��w��Ux�j�n����333���U^*ڮۻ�������}�*�mWm��Vfffg���W������Ϩ�C
0�g,��p�x�8pgl����jBHIl�_Ҥ�U��F�Δ�
��0�:j���
�S�wHѲ����lc���)(gEGO�qi[�m��(Y�ÁC5���J�6�.+�I�)Uۍ�Pj�BA$��	Ѷ�GJ���C 4E�����!�he���6�t�ih�ճ�&�K��ѵ�C�T��k`E�M���WC�.�G$r#H�uYHhB�]��Z�4hgHl�F��:a��0�a���n5����q-��$^��m��m�{:��3��L=-&��o��Cm��ia�h���qW�C	ӳ��-���h��(�;U�}���e{\�x��b����M��-&����kG��ٱ�͋d-fY�Rz]�(�eآ\��m�����F��l�hZGzY6���><�2�Ϧ���6��t|�1p,g��,���<�6�X�b�%��F�=,Xg�:<-�3�>4Q���>8|p�x�8pgX�A�-��BEۥβ�EW�*N�����"n�޶ֹ;TB�aI�T�:����	 �	/�7��>����L���Lὂ��IXNY���a7�w�$z�>k�pTX¢��˲���oon��r������܌Wu�Un|�c/z�RN���p�wۀ�~͛�����pYO&���wͼ�������֬#˄I��q���|�����6֑�`ϣG��΂8�,3�EFÛѳ��f[B��H�[��{�6�͠�2�G��۟G�H�G��"t��yZ:t(:u2�ͦYi0���u4J�a����\�ݶT0 �|���ϲbԘ�Xsd�X�rI�e(P�!���	f�><x���O�����<R�׽�QsdM�\%�q'��m�!$D<��g�͌Ѷq�ؔ`����5����6�O���F����r67$��QJ�(��E/�G{�9t9J<�t��l��6����x�p�Hw����;�t|b�/�F.4s`�|����.�ﾣ|5%�Z���Տ�nl��1F�#�͆��m��Z>�f}�L��~L����%�(,5��5�-��C�<����/����h�f|pÇ0��x�Ã8Ci���e��"�M(C� �,�}kM��M�M}� eUS�UT:�����_W-,����"�G�|L��)p�:�d���fT��Ca����s�p��M]ު�&��<Q�h��C����.D6|�~�>)�[E�:ڷ�t�j�#_�wta��e+ x6t�_/0�qE�ђI$���l��6i�h�K���6�Y��Ţ��6p� YC>!�E6Y�8|l�x�8pgm_2�5N��	�CekZ�\�P�BH�t
�W2�Q-(�����H5��š�G�	���G#dc�Q��7kmHWAשqy.��~�h(�_j���&��l��0g�gHkŊ0�Y�
.���U��#Y�='ݭ��g��u7RISZ(����Z
6�ѲΔb1B�IÈ��Q�Hv���|P�\6}�����H�F$��a��h�(�e�p�g0�p�|8`���_�U
R�=x�*+';*���a��*���^ ��[�#[��5x[��'��kM��M�H_�c5���}�:�aHpk�P��_K�6^ ޜ�C�'��p�'k��'b.�k�Tܚ㵕�"(Vf����J�p᱊*�����e��P��Xm�U��+2Ez�Z���0�cz��08l���#{,�S)yb6RX)G�\5�����&U#�֧E�~<��� ��A�����[w;�"����6Y������|�])��dT�m��k5Q(�S��O5����6�U��v˒����F�]ז���I4Tߊ���.�E�E*K�G~m�ƾ1y��(��>8aÆ`�	���GD犓�nH7�r�/׻��Ip�5�~���DB�34m(���b l�J������ց%�W���ɾm��]��uWvT�8]����w��b8f�^8�-t�Ŵ�!T#�_SqC4=��MGQË@h�6�m���p��:bV���������i����%�����n�^֎��|5�����0��x�g4l:ib�9�"��d��HV7��og��ԅ������(�e�>8a��a�<t���!��-ª��%�ME^�UU0���H$�K�����ܗr�.��o�����fέd�r��C�K�Ѥ|�@��l}4��G�}G��>5���G��&��E�/*Cz�P�Q�J2H6�6��a�GCj����F���ŷ�pᮆ͡��Ej���i��ż����)!�]=�^0���2����V��㧏�?�GC�[�{;ϴ����0؛:~>??><||&x�Ӄ8Cf牛��2V�t�&�${��(�Bo+J�X����6Ӑ�"�9F(i���6Z�83�3F�4}�h4�4�����Y}�?�m� ������Ƨ�KUQ�v�Z�l��|b1UAD5��{����E���YW�ֶ���n�K����8`�{a�Ӣ��\=�a3�
-:�m�ǄD4O��G��.���f���x�C�}�rI�M.%�Ѡ�f�6Y�}�Y�C:���B�DK�&��<>'D鲎�	� �'�f͛dM���'D��`�lL��&	�"&�
��,A�x�H"lN	�DL:"&	�,Kı�8B� �6""xD�H"xN	�:"`�"'���8A,�f�ؔ%�HFM �0 ���(�Ie�a�g��0��O�(�>> ��"&�0��a�L��a�����A�����r���a�}<C|�+Ӝ�>�u�����v��Z��#��օ�$���Az���5��[2A�%i�̤�]t�9	E,N5��)�啮�ck}4(�[�)݆}t*��֪�m:����d�c���*�K߱?��>G�_?Qq�����D�"���z�+�Y�b>�u&�0�f&*d�H�T�YU���]d
��"�� �.7۸o�*�+�:���pVǹS��Rb���ҟ�&6�������jfl$�IꝌҀ&�K�P�A����0�!WS[2]$�fS��P��{��/o�9U1�)��Z�&���u������1���q�c5f@-�8��۟�vƆ>r��Z2v�H��R��&#+gt�BT	�a����:T3�~k��|�J��]��ws�������R��Wj�����������R��Wj����������>���]��ww��Z�a�(�FΝ0�8a��0�ӧ����Ǜ����c���(0�"v�s��w'\���z���6��'"����r����;6���}�8y��8�b�hp�N-t�ܺ6z��K�v�ɣnz�����r�W7~��`�����Ź=�Ѳpv9v	�r��9�.��Ov�m(>�m���;�a<�<�q�ru�P�n(���PI�M2���F�g%7X���4<�A\�1E�;����F����v�70�C��[c\�q���}5�qr�^yƹ���x���w��<�v⸮���笅X�v�Nqf��ɴ�y�v:tq�x8㮅�� ��pv,��۵Ν�S�Ϥ��:C]�T��yc�lq��J㭸ݱ�iUy���q�J�Y�7[�ݍ�^簾{e]�g��B2���n5 ��U�,�Ś�瑸j���ۋw�v�	� ��-���6�m6�!:�dP�ǭP�]��7Y%g<�Zt��]fd<���׺�5�НG�m�_^*�gGJbgU�M��E�<�m�]31��e�ҥs��=9!� |��^�2��Fs��'�x�z�Q�D����[�7�#kl�Ʒ�٠������%#b�Y%����G�#���ylь�l��3�����t�
�Ɛ3�dG�-����aHt5�U�j-��#�o��RuF��G@鋧آ>�m��i���I�*�/��Z��x�6�k��+L^������-X�rO��a�顜!�J>(ه��0��<a��83�\S��v51�5�2�0���l����!$$����<�@eSr�vuNϬ,��#7	�"��&f3L��V�����{
GQ�ͱң���|U\�3���T|x�Ph�u�4�9Z6�;�=oq��^lX8>�e����L�N ȟ��܊+A(�/*�&��3�5�0(�1t�9��"���f(�7������M��#1�2��F�m�Z�eᢏ�:p�����0��x�Ӄ8Cg7��t��U�C"�J��	!$$����H�#!�_!y�q��>��#dW��CZ>9��#�\\4�G��:Z<�h�C߁$�(A3>#�<�ghk�#�R�64�d�c8m��>�6CB}�k�����~cG�]6<�#�x<Z�\�����Т���l�n�l�H$H��٩$�tT���Dq.�/p!��!f�0��p�æ�0�8t���^�S��s�[;��Kh2�~w��q"!�}g9�>�H�E%��|�hk�ب�A&�T�۽��w�_��*�J8n�ʼF�E(�A��`�4��$ƥI�[&�Xx( ��|F��Őe
Db(Z+�ԭ��+F͚L���̩NRp���8||��:Y�h�^G-��3�0�������a�M�1�o��{$m�m<e��b��&��l�3c4Cg�<QӇ��a�fx�:pgl�y*��n�0{uUv[/�J�%�S�����ȝSv��Z-q��X��,���_��)�rH$��+��6{,M�[����70'�c��Y9[���<-к�%P�l�����ip�q�X�=&�ڦ�Z��u�q8����A�8ǧq[�Sq�1˸�˜8ǯ*�J�:�D�,�#e0��ECG�E�ɯ���g[�����٢��iR�b(,�?��Xǳ-�#Agx���Lp�M�����Dah����"�1�p���4gEgۣ���<"�7�{-��� X�m�����!ԎT��v��_5�3h�R8uJ|�oM78������Yp��(�GN>8a�L8a�<p�ќ!��N=�(�J�bl�D�B��!$$���:��}�鈣�k�Ө�Y�l�/Jo�h���A���{r���+U��uH�:|@�д�y�Ɠhċ;C0�8���Y���k@R,�-����Cg���S�F�8��X�X� w򸹞��`�Y�l�2(D����xm��klm�8����h�n��[7����V$��8Q��0��:a�a�N����{�wD!m:�v�Y�BHI	"!�?rJp�����:�����pk�R�6�F���\Tr��H���X3���E� !AcԢ���x��I�i�:��S��u;����8�Q��Q�ɇ�p���H��f�t�uha�]�log��3˰��9)و��K���q�R�W��2涹CM�:n�i}�s��h�P�]4�Ѡ��t��>:a���a��x�ӣ:Cdz��EP��z�:��BHI���c��j9挎GذW��ڭ�q(�3ՇE��?���EIAv�2ȩp~$��E(�m �㔗�ڍ)��;m�H�o��H��C�F��K��/zr-���
b�Y�GC�=��kD{����)�4mq����6�h��)l�a�|�O��oH�5�q�߃�>��Z���e��4Q�0��L0��<p�ѝ!���nn�4�)$*�Q�(�Mwp5�b���0�aL[+	�
m��uaD�DBʲT*���z���BHI��!�K��G�gB�H�
h\ߗ\˧�T�a�c&U���UNh^Z��*p��i��z�(����osL����̂���F'ȱ4�!��[$t`�Dh�c��ς��$yN,�vӓ+~�]�	Z��4^��/�����υ�#�iR��eil�>H�;ޜZ�ţ��p0�h��o�Q��8�bGÎ:hڃ'Hmͻy�x��ǑӨ��iR�Epp�ٰ�I&��j�.qu2��ۑ��U�n]߷Z�Sn�����PZ�C��j�X��8��=K����0�,��aG��O�a�8x�:tgH����g6��eM����M��NDB(��G��ē���ӿ7�F����|�\Gǂ~Ci�nյ*	�����x\��TZ16>����p(��١��T/&=�&:��DЏ�l:@��\��gJG�*�:-:��<��H�(����IGu'��B�ʬ��fd,Ը�P�WHX���<�0�Xx�H\<m(�7���p8����Zڤ|#����h�+���q2�%8l�g�,٣g��:Yd>� ��""&	� ��"'DL<pN	�,�@�X� ��؉�6"pD��xLÂ`��0DD��D�D��N�""p�"lN�L:"'��%�bY���4#$��DD�<P�$�A:"`�'D��8'lN(M��,M�A�`"P�J8"Q��Q��<x����>0������%���D��ç�O�
>���A�`�%ɬ�oU^z�꫺�$3�P#�mY�kiP��� �{8m���#��[�_|a�����$�S�n�v���ݤ�h����S�?3���Ȇ��h�+�����s����|�p̨��F�x�۾�U}l�ʵ��;3�9�)�B��^P��6��+#�����m���+�~W��G-n;�r�:j������U�(�"��O�Ӕ�`_��ϳ���V����ffff}�EU_-*�wv�ffff}�EU_-*�wv�ffff}�*��iU����XtgHt�GJ:t�0�<a��:3��{W	!$$��1�7h�6b�0��넥\��dk��;��~�➲JGA�kx�g�&�#����l�ծR>R���]SQ�)������\�-����,t�������rgZ=���/㡓�*6@Ϗ#�Ax8W�G��C_5�:޺""�I�-e���DyY�����d>4QҎ�:x��L0��<p�ўO����2!H ��1 cx�����b���4�M��E�S}mx���il8���Xw�x�a�~�#��]���f]Qe]��L���n�|�[L�#�I������7W�$�FÊ�Me.��AF&�F�l#�JY�t��#���x����\�%�WUm�F�X������s��u2��h�ڹA�h>������↶uC@�m��	��g��D"l!��!�e(�O�t�0����m�hw��!�)�<Xn@�eF��qT�o"�ҥ��)�C\�M���\�AUB��2>�~�m��m����	]�r����M/q�cc����<���M���uN�+��pb�x��sX�����FP�/�n㚒y��j7��yսw�0�Cf�f�(�'����6�wې��qӕ<��0�8/��hi�����&k�R�"F�x�p/��΍2�n��k�F��u�R�T����Vh�Z6�_!��]>m����k�J4y���hz�E�^@�|�/������i�Ӳ��W������f�
Ge�h�kJ�|y��6���c<CgJ0�0����a��x�ӣ:M�f�G˥�T��Z���7���B���g�$$���j���l�������?%�ⵣ���"���ލ�1a����m"�7��A�x�9�&/�h�ӧ��f�&������ ���H��]3�C�H`j���U.��N/-S7��~��#��ol ؙ��Zޛ�w�Z[lm���{�Z��ةY�<�������d�>(�G�L<p��a��p��A�C�-��I.$�Ct3��$���#�⥣h�:�8���5Rz��Q���g�������c�G��K)l��x���;��Wu�c����/b�]FxF��ž�3�ы�7�ԍ�@�x�x���3�O��߯��Zᯠ�?�Χ�qv��ա�R�gٹ��ێS�O�[m?��F���H��~FÆ�Q>(�G�8|a�6x�4h#B�o)|F�*�4B�T.�a$$���>�E�[�v�Z,�h��Q���iN>�C�J��F:q�c�]jִ�"�4oQ�5�5����>��hb�gC�����6�abI��m�q�1��cY��4tW�}��mv��EV����)�dc=���uD�<��1oe[G���4:{���s-�ypͦ���8�k�3��C���%	�bl��:'��0�<p�ѝ&۷�z��r�l��	\�dr=�i�y@��"�\�r�M3�v��-1S1lo��ݤ���Ws/Kg���6�}�}z�H$�K�K���n�"�8��f��M��B"ܭ��w}�q���ʲ0N��1o���t2�xΣ*-ݳ��m�MU��v/��$]WU��Ld�����FŸ^c���j��4+��x3���ν��w:��I��0Z��X�bx�<�h"׻{�T�)�hF¢lƆ�ш��bg6ƍ��#G��Mw�����Z��StR"=��,T��>�{F-��?���kL�,ME��Á\��<x��G�@�0�Ջ�W��V��^w_6Red�M:Ur�{J��1˪`C���;4�_FȊ4��e��<Q�G�6x��a�fx�ӣ:M��֤%��(�EUNE�I	!$F#�T�-,V�h'ZM�6���p�XQ�U�ҤR(�k�i��Ⳇ���I���vDul+�o��:tͦ�Q��VI�H�c��Aq�|a��٥�σ+�
Ə�e4*`Y��}!�"?~�4��T��
t���C}�����%�q-����.8͢���������t�4�G��2�p�G�8x�����a�fx�ӣ:M��[�#�Ha��<7\�Q==��M����+J�#�p8�1��x0� ����oPn2p���m�t�4a�Ű�q-���>e�\,L�>> |���<�|o���8.�ڿ|�L��][�G'��x��MC ��E���E�I� y a������=qQ����u�6C#����]G=��#���q+�8x8���_n�%8�"��͐��t��a�<l�:tgI���݉��7(��~�p�e#f��5�����N�:�_:����l�v8��	��i<���ȇ�iQ{�:��Dcn;��Q���WN�[\�l����-m�q|�B�H���5Ђ�H.N﷪֞�c���[t�tx�C�gL\GH��h���ʦ���`D@&���w�VlM�%���:'�p�0�"'DL�"A,DD�""t����H �A��6&�8"xN��	�`�&	��&	�&	���d�D����"Q�'H"lDN	�D���8%�bX�l��i�"&	҄ ��"'Dؘ""a�����b$!bQA�%ܚH=�:&��͔a��>>>����>>�DO	�x��f�<h��00�� G��A)�}v�_J�IU�+��S��ZFa���o���i%�'���UdGTd(��9eh�+(��Ωt������G3����ާ赅9���/Xi>���n-�YE�R��u���
˛ۃ�����a�y�,:l�K#ݣ�(�8�ۺ�d*���h��V��/��H�_	��ܼ���_DEgd�v$�V��ϕ@���G��S)^��k���Y��8]��W�LK�X��4�L��ta�t�6�4�2釧5n����p����1fjƭ�zV�ow�BO���"e��p"%���p��Л+
I�7Q�b4�k�Вnq�g�����p\���Q�ʙY])����Al���w�T��l�*@W��7L�C�ˆ��]��e����^��/�~EU_-*�wv�����ϾEUW����񙙙��Ȫ��[��~�fffg�"���Un���K�Ft�N�t��L6x��a�fx`Ѡ��"\h|�D�B"#���<_��8�.��棕@��ػl�q��n�tS���9�]��ڜ=>-լ�q�;0u��4��"��&F���3��<v��Ro!�o��� ATc���
�"dn܄��^�{q�=s��ti�*
U#n���7l�Ռ�A��Kn��Y�x�%$��p�k���c��n���]T/f��D�%M
�V�[ N��u���t<lt�;����sI��e��V��+/k�r�g��Bۤ-q�{����p�ݳl��"�(I�$�)�qr8=Z��2��'���ף[l��!9�o>;���q�;ZE��]q�c���+n^�;fݡ�7����G7-�p>0��bx���i���A̜S�	��*7,�[/��M��M�QBs��m�Ŏ�|w��};T�ɦ�	�U�՝C%�i��s;R\�t�υ�X��j��e�y��E&�T/�"�A~�[����7O��Yᚇv���&�^�Gj��Y7�+=@�>+:텛B�s�)����,ш��u���Zn���][)�ٳ��:F#H��/k��Zh���|�Z�p�K7�߆����V]�t�[�.��U�!\\S��_��e|���8��h`��4@�M�4{�_4}��c�`l�۩!*UP��*~*���D��ط/ ���(��{ý��#dC^6uu}��g�9�j����t��<|a�<a�4h#F-@�4$V�5k��T���7^KN���1O���+q}f"P_�c1b:�8�&ͨx���H@�~ŹDb�8�6�(��o�m����	��h>
P�J�	��˴4y_��Q�aM�m�>��\��8�ܯ�,�.��|��yCA���gLP����c�qσHŇ����$�v��mQ�^M/a��t�e��g��|��(���a�L0��<p�ѝ8Q�y<h#D*�eB&gX���,�m���"l��FRد`"�/�bκ��[��8�I�&
�/-���Zf���|�lų�5�NrUTsG�wp�W�lG����G�q>�k��M�c�дl��˨��;\]���ni-�#�s��m��F�&唎hٺzCG����|�i�y�6 �M�G
>:xنt�l���Ӆ��e�W���jj��!���������1}�h�4M1�����ʥ5�B?�wt�Ti� �"�/->��<�#�n�Ix4�G�쌌�#���x!�庴b7H�kA��M�<���Z����%�}B��X:�_$��&H)Z,�m�KF�F����u$�IB#H�B���uP�e�-Y��D��Q��a�0�0ه�:3�
'K�	�ܳ�TA�5դ\��="جwoQ>
��v����l�� (��t�Rw� �O��
��s/�*����
�bֻ:ڭOqn�
�.��Cr۴��Z���kxmT�D�ZE����P���DR���,������A<�mզv����:��
��W*�Z���^C��>"� ���_u��:�]�壣�T>8F�[+�E�ab�.#���,C:��9������߽5��3RH9�h�7�:Cc[<��و�'�ٴ�zc'��l�WT~n��z��M�k�e���F:Fϲ�6CE���~#KAJSM����ҍ�l�ǌ6|a�L0��<p�ѝ8Q4wn=M�F��ۛ�Ɓv�^b1o�	��f�q���]GB�����E�F��4��iѱ���t���7
D��|Ê͡����0�Sm�:GI��[�|qn,�����g�}������jQ��(J��rP��?x�b��f4�0i�hl��](�����:�8�Z+l������R*��O�GP�-Y	3Tk���� �6Qҏ�0��g�t�l���Ӆ�r-H��:q�#����J/��]��
&�M������lf��E%��x1������Gв�t�@�M�
���֍���[Gy���ɴ1�G���#�@N�ub�ʫ"�)���M��4kUn�]�6��x���q��hi��}���l�$�Z>L,6��ϖ�h�ȶ6�L�]
mdf��Jd�����{��#K9��]��cm�z-E�
 �8Q⏋>:xنt�l���Ӆ��ʦ�T�ýccchkgO�c!��9����.�||�=gC{6��NEEQGg�~#ZJ�&�c.�Tu�����ČpYc�f����[l����[F����aiR4��
�-*jѳǆ�yiuu{��P�+����Ҍ1m�I|�m���< �׶�-l�� R��6B��?}c[42�|Q��>6a�0��0�F�4``�0�n���P��2��1
���a��W�]3�{'�e=������������9�{��@�+��m������\��;r�.���/3��v;�r��m��L-�	�Z�rc��sY�&I�c�uÙ���9]`�t���㮅T�N�T��c��m"h��!cs���;��2���@���/�����b":�C���&Z�4���Kh�����""��m�'čɤaݣHl��"�CE#x:-0�����h����e�]������GL����˫�|�9���]ӳ�J��f��m��p��+�|���6�e�>CKLo�iqyP�8Qa��Ϗt�h�g᲍f0Cc���E��%5��1u=��iR��a�����43��1��'$i�5�lv����r(l0�-i��6�� am�֛d�m:�9ѷa�l���{ZF����X����|�ERR�%��`!���i���!�A�d-�s)�k֑Z�@�a��a��Vuf�#I�b�X���<Z4|!��aÇ��<l(���0N� ��"'O�"`�8'ᲄ� �xA(J)&�Kb%�<'��	�`�&	�C�0D�x�A(DN��0C�$�B&�D��B`��8'D�,K6x�(��<'JDJ�"a�0Dâp��,�X�!�(D��&� �t��$,	�:&��Fx��Ǆ��O�|||'O�"`�8x��E�a�fІ>�����Ջ>�R�_R�!�^ݡ���-�O[sz<fήё�v���Y�ƭj��*���� +[xh���g�*�Ӧ;`��,#e���u��R�V��j���ށ�(���-2e����/�����a�>��ˎ�c�����w,9�ݪ���UP�#aH���|f��az�꩸�����2��n��úԤD4
���5n�~6A2�M�fmР��э��*S{�Q����GW�}���S.�?��:�������}��"���Un���������UUq���ݿd���Ͼ�UUTUn���&fff}��UU�Un���t�Ν(�GK:t�f8a�0�4�:$�+l�A ��x��%ʔQn.Fp��Υ�cn��2�2��M�mZ4�0��t�����Kh�(�a��}����I욪ԕx��z��F�Ai(=�wo��D����;�I�Q6�����[Z-!�b�uA����o�V����s�9�*Fր�m�6���予E��|� �(t��x�x��<p�ѝ8Q�y��-꣎�d��m��4iR6�uFp:��|�b���0k)6�)��1 �L�%�+��t
"4X�Хe#e���+F��6!��Xͭj�ş7���A�Ͷ�|w�6��8�m�kg>WK��n��#�2�C}�tI�/��u.��Q;�$|�6��Z�[6Y�gM�X������>6|x�ӣ:p�wOt��&�T������n��gtkKȭ��gcɽ�1��0��뮴W\M4�J�o��D�I ��O�#���?-ƨ�f�u��GNMY�a�!�S}��^lZ�����q:���LҝP�ݪd���V��Z�0�w��ʪx����\2�oZuD��5��}Ӎmh��h�+E��"-z�<���
G�n}����"�8 �����T���;���9�j�M4=[��8϶{z�`�h�>V���y��-j��B�k#�K��H���G܃i�/0�/����"a���vB��QH���Z<����	�h��C[Մ(�x��bX�>�||&x�çFt�Ey`*ho���ְ3e_@ �y�sqE���֕��^9$�$]_���/�h[�mk�m��5C����w�xݜ8G�mu�ǯ��M�G��~ѦRۏ�S����V��z��?��M�H�i�G�\��Xn���Ǔ٤�����	��_���t8�"��,��?1��6ܐ��SX�o�K�ؐ��a�HՐ,Hl�gM�X����O0��x�çFt�E��::�1�;� �^�(q!����������|����x�)����4Z(�i�$%l�ֶ�C��n��>��T�E�!R���U�r�+m���Q�FiZ⮮�����H����ƍk	:i�R-Yd(wDlc����B
}�8�1�/�#
��bk��h4 �(�G:|a���a��z:pg�t���$؃��5�л@ _�I�����c4�3��6hh��̢)[����f׭���WO����1D�>_a����,�ߗ�Dc�VuRhh�k�|m��m��3����:��!#���"���-��P�^4K��-[X4a\ccڇ�QF�u�>�`Pu�/:}�Ë��0-`2���bY��N�����|Y��,1Ah�҇��9K��B�;j��{����s�o@[��K9�+R':ඵ��%uH�U�u��$d쩣N���U#N�n�ˉ/�![���*��>Ǣ��~�}F�;�'O�,�Z�q|Er���2\��v���9��Ɓ��Q��㦨Wc�=�+bߣ��V;�YapF�j�ޭ�m�C,�t몛���#��������z�*m���Ëa�D\m�h�K��I(��L�n��\��{�j���T�yV��s���mᵴa��x6��������&�*8��MF�\(���r{�[.訫r���'�wV��1r��������3֛�����Q���l�0ه�<a��YӃ8l�AG{l�붋��Y4��$�H#�傆#H��`U�M���cm��ū䬿�R�2Gw�\T�4|y�,��|S ��<o�Ńi�#���!��I��DFJv���J����s��wUn1�#P7*L�v�T,@���i4>�����cZ5M�FHރd�h���Ӧ#�GZ8lg�E!��vWG�/9a�SM������G���e6ag�?>�'�|a�f!����Dc Ɔ���;�M[H"��$�H�[
D�H�z{<,w-�կX�@����i����P����.����B*M��\�\�[�De�,~=�4�8�/�길�C��#�GD�Y�I�p6��7�}Q����p����4qa�C�$��zVCh�|�F#��$�K���v7����u끀�K�R�*�cM�7�O����a�g�gň���0æt��(q�cp�r�ITH�֛m�}�m_Aפl�A�J���A��X�<l�C�>���]7EU�i����Cᾓ܇���/I<C!�A�G�޷$>m����ѣH�4���YȄ��"��SwW�-˗���l��b��q3H��8��U���4�Xy���ٲ��n��� _п���M)e}�UR��6���/�_�ȗ�'K?�����������B -���i��]"&_
U`�l��Y�����3u�Qi�E��i盉-1h��Ih-�i%�-�i�1i��Zb�i%����h-5��Y�ȴ�,�Z덝%�%�d��D�ȴId��Y���E��d�E��E�I6�Ii%�i"i��K"�E�KM�����%���Id�4��%���,�kE��е�CsE�I-"Y$�mK$KI-��I6��M&H�H��K&�Id��Id�d�i-"Y"Y"Y"Zmd��Im$�D����K$�Y$��&�I,�Y,�Id���Ki�$�KM����I,�-��ۮ�Β��%�%�%��I-����I%��k$Ki$�%���ki%���Im$��mm$�D�Im$��m%��4��[I$��Im$�D��[I,�D��[I,�ZIi��I��%�K$�ZD�D�Ii%��Cs"�ZIii&֒ZDY,�ZI��%�%�KD�M�KI-$��ZId�iȲm�%�%��-��Y$��d��%�M�"Y$�֖��%��Ai%��EM��d����i����"B�"�!4�E�h��&։-"Ih�DD�%�"ɴKI�ZH��KD��E���K!h�-&�M�ihSZb�"ɬ�&,�%�ȲbȲI%�ɋ"�"Ȅőd֋&,�Ȳ,��Ȳ$�bɬ�"%�Md�X���#[hѣF�6�1؍i���8��m25�b4�h#Aևk4�mlF���N1�Y��#CF�#Fѣ#[e���gN8�4�Im�kb5�̍m��h�����h�4؍��5�5��m��#Y��M��dk24�@�fѣ��m�X���؍l#F#h4hdkf�f#LѠF�F��M�ml�cF��[�Ѭ�4�ͣCF��5�5�٣FѦ�4dh�5�XF�#[4i��F��[4i�5�ѭ�6��ѦF�h�؍a�M�Ѳ4b5���,d,�fBcB�Bِ�гd4ƅ�Л�h[4-�	���	�	�v뤔���Bm�M��BlB١3Bm�`�#i�i�&�Mf�ƚl��&��bl����2i��ɦ&���km5�6A5�h&�M6�m4�5��bk	��MlMa5�4d�M15�4�i���&��̚�Mm��ɦi�&��g2�6I��Mm5�I��ɤ��d�ɤ�k&��4��i6I���[M&�i5��Md�Y4�Md�ki�֚,rYMd�kI�֛"4ɤ�k&���&��$�M&��Mm4��i4�-��Y4Md�5��Md�l�[&�[M&��Md�k&ȚMm5��i5�D�Me�D�Mm5�D�M&��&�&���&�i��h�ɤ�m4�Mm4��i5��hM�5��k&����Y4Md:냩�&�h�ɢki���I���5��hM&��kMd�l�4��[L�m���",��MdZ2ѭ�#-$Y--FDX�"B�"ȴZ2E�E�B�"��,�����"2ȑdDY��"���d�DE��"D��",��ѵ�D��HZ"-
$5�E�E�D��2"Ȉ�"DE�#$Y-Bh���D��Bђ����DCZ$Z"$MDC��4$Z$Z-�!d&�FHYF�Z �
-ѵ��5��6�5���0��YB���YB���Y��dK��5�̍d,�d5��,�dmdZ,�E�������5���dhBѵ�hօ�kF�-Z5�ZFݣ�5�ZБh�h։�ۚ5�Z"!2дHZ��kB�� ���"дŢ�Zb�Z--$����Zb�h�Ih-4Mh�Ţ�d�f�� �~�u�j~&��(�l�k��~��Y�0��ʦ�f̩li��d��g�'�w�;��?���������L?�a?�k����ٯ���o�������}��^?�\��Pͳ�g�@����?��C������
����г�������m�h?�_���Y���$����_�������)�����f7����Y�l���������o�v���_�����{�mg>���?Ż�#�~���;?Gԟ���>m����������G|����M�x�g��Svߧ}^�:�~9��?�DDG�#��l��ý�g?p�����{�>ϻ���i���w�����ws}|�0�}]�m�t��6:�cq�5��6�������3X`Ep���OO1����=>=go�k��������$62��l�P�cZ���`P�fP��`���=�#��i���y��x���������7�{��������8�ӿ�߼[��������&�63�=����nߟ�o���&��'��V����^>[��폎�zf�m������>����vo�e��|����~�>{��o��{���߫6́�7�m���~;S�|9������������>��͛l��~��6������~����\u��v;�������w�/�=���/l�8�?�|��6n����jO��N��ط�:��m�������ku��7��:h���ۅ����ݴ"lG�����T5L,��UĴ��y���?���`s7�{��T���~_��_����fٰ>�����#_�>������n�����O������ٟ���-�l���o\��O�~;��[��������d����+�����|���f�����>����n��o���ͳ`y7��~/^_���������ϩ�>�׷�v�u�m��f��i�kG���7ga����6��wɿ-۟�~��4�����@��h?_hE˴o�+U�V.�{�|�6��+�o�|�;nd埆}{�o���t����cy7�}�'��>6y�>�N{xv9�n����?nxl��Y�[0ٿ����>ͽ�g�?���7�����0پ�����~��~\���x�{9�s��ާ|�g���Oݜ�di�����~���"�(HXe��