BZh91AY&SY��hW�{_�py����߰����  a��        �       ;xP��UH(� �B���"!@IAU)QE/���"�$�B��� �
=A�'���*�}�^��n������wxx{��n�幷�3��ޮo.��@��ozǯ>�{�HK��'�@�)
餀U��3�w���i=�J��R�MVo��Ra�\��{ev�zj=���x��*��֒���=ԏ ��L���7l0��z�+OK��N��f��zpz�i�wiUn�C@H� �%���v���l��zc���{j6�ev{��ǫ�K^�.���A�=��Ux��	��L������^�G����Z����4�a�zZ�����{����u�Z��7�.����{�˦� @����i�����ڻ9����MǗ�K�'D��ӳ��   P�Ǐm�;�л^ܮ��κm���Ԭ���띧��(�֨T箳��j��y޶J�۶��6���x���j�n�{ؽo#S�@        h     4         � ����J����A�M=L L��2`�`5?B"JUM `4  M h j~E"��i�     L10�H�%J�LF��4�
���!4OA'�)�h�S�Dl#DP�jT�F�L` i�o#���㇜��pr����uwON�ٳ\�:���ffٺ�f1��fټٿ��O�\p�^�f��nٳ��o���ž�듩�?���jXo�F�ٳL�'�t�Upq���6͛�l��L�*���l�V�-��u��c����'����~�f�=q�������O���8�1�*�aOG��R^E8R!�S$d�[�,��1�c(OvC��3FM2D�3��@�h���f�&AC8�B�Jc6n�*;�+`��I�
ͅ8�:�`�|F"]¢�&���/����D&Y)g֖E�Bd�;�L��¶Yu�(d#	�C$�da�2	zE�9�+8��ߙ�л�P�#
0�p�xYE;���A"�/�J�0��^&i�ffd,$�X��b/�l��-p�ax%�}�ʂ`ac��X�YqP���ĸfLd&?�cN����p��I�
�AXIԑD� ��B��1���X�Q�d&H�+R(cJ`K�<�L���,$��d&`�}
�p�3���L�/��!2�>�,g`�K���#F3�o28��^/�8L��6\,$���1��c��3�fI3��f�Kp��K)2�37H���(��rp��K��50�d�BLe�q�����c �p��I��S�P1�ZN�-��2�C6�Ӌ���d@��ZFmi؄��Y&�*�qc#p�:�]�Y�?��ߴ����d��ԙ�o��1�f�O��UBLc��wq�Ab�E3CK�D��,��wrVQ_�aض�7��
u
��B���`�+?�.Y��Zd1��4Ƒ��ÅCeL$fs��s� cW�.Ygc��8W��3�B�]��"�I���H����,��*R$��9_0a�$>_2D�便���u�f��*$���ƌwЙ�n���.,��B�������	��<�Lf�N�$�����!3J'�� c���6�ƶ"i1���g:�X2��i#%,��ɚ��i?1�`�1�2ũ�E�Hc�1���	�xC�a3,,e�&1��(4�4�A��L��\..Yc��0C�"��q����1��3�.Ռ����Q�[����Di�E-0`�Gck$f=P�����H����f�3�9چ3	�#�5A#��e�f>P�2�!�X�T|���1/��-$�nT3F3��1�h�`��j0��$�'
���1�3R��!��b|�Q���L��r��(s����ʆ1���� uJ�=LgmDc�c���F1¡�s����9Q�$1x��9ʌ$�Lbz��d��k�3$s�>a??� c%��C6D3^(��3��a�$q�>a�SQ$d�P�i}dڈ�>�X�j��?�Q�2]�c0f�!���qX�\C�����F����ǹp�8���L���#1�P�"�I���ڋ(��ɖ2�(f����م�����(��:؆[�M�B ���,e�23���0�~���w
F=L|� �z�d�c����F�⎥����Js��ˆKHӄ����&2a��k�+&!*�Kȋ&� f�P�(��gn�q��}��R#>4�	@�C���ځ��=�z���[==|l�}�S�Y�>���b��3�Í/蘂T�W��e��"�3Jn"�0��2�S0��`���i����N0�
,a��3��F9�h�|�FN�H�1�ڌ��"U�C�1�:Le4��d9P�>L�_�E��1��C�cJ�ǉ�ck�|�&�a#-1�j�4/�ɉ��UI-
F2FKj c5ʆ;L�z#�Ì%(4b�P�x��c��Rh�[���3)E�ME���b��[؍��Q�.��1��3�s�8w��(�f�P�J�Hg�����<�SHO���(�v�ǋ�s�L/�G|1�S�4�qiC�'��>���C4{�0fI:BaD�1�Q��0`�i&`�i)I�f�L��c��P�Q��c9�FU�`��|��qD1�������3�XD,���g3
$��e�LʈX:H�V3���k�RY%�2�d�{��þ��B���3�t�\3M�C0*��Ic0�
��"-���a�p�e:P�)��H�NpD�V1����QD��D}#E}0@�s4�j�<��*�$�bL��j(�AOT`�)�E4��CꈙđD��&�E�(z��F	�E����$�Lҧ1SJGjtX�]dĨDؔD��LB&>L��I�DI����I�D8I��P��1	��!w�)BN����C�	�q�. lI�i���Ac؈f�3qi�XH��C$��J�H�6�;�|ǋ�Sj0����P�أ���C$3��1��G���1�d�1�c9��
(c���5��e�>t����gq�0���@�C(ck-����P��@�X3�r��c�c��Hg��f:P�Δh�r������D5@2�������5���(��f2�(e�sj�(o��8{J,f�R2/��}`�x���$�8b��|��G�p�1����Bc&v�ǫF3�YC��U��4��#�;�I��Bu����6��1/���p��2(e��r��ԡ�2ިd�m%���$p��S���,�c.�W'i�c7�+��
�12�.�V"�1�&p��O
��$�"L��3�%�����(�I�0�ई�8I��Y%=���+"Dɇ	�+* �1�4���f��҉e��B�~�if��t��n�k���%*L(r�c����+Ia��3����1��J�J)�;_1ꁔ>�L吸��i�Bdc)�Q&�!��21XI#(qdQm/������l���8ᓼC(��'�A;_0��L���#��ä��(f��E��Oc��|8'G|���8v�a+���+;�%3����H���Y��O;��������l�$�s�e��}�����:wj�7�����{T�����쇬æ>��!e�l�I��M��ݿn�|���·{m`>�0�����������n+ׁQ�7_fnod�wپ�da�5� Ic�b�{�1�j;���_K�����5wX�#�M��wv��}��z��N���\E�sy��*���Ǻ��V�l������3G�����X�����U���Ȼ�I߽�c�[t~��ڝ���L>Yu�c��T������9\�QqV�]ȵr�����,\�Y7}TS�ʟNι�����F���^���n��̠ިy�F����퓜�^��WB���[?)�̋��d�3}U�>�L���.f�'՗���FFh�̍f�t��vozfy��2�����=$�vN��c����M�h��Ĝ~DWt�T��g���!w��aᤤ��N͝F��!S]��zj��+1d�U,Q��N��E}u�W��i��du;I���jz�.�ǹ9I]�VE��^���M),�\5u��Z�}��ro��}^�U,�����{��VZuJ�%�T~�+��ߧ}�w��gV)^�`H���o�i�{�	�����w���7tp�l�苝�6����{�է���;I����W3���Mх�]����z����v_7�
���\���������f���|8�XX��)��j�V���0�&np����Q�3&rzL���ϛ������\����~뎵�2��5�tw0-C������������}7�\�-�vl�3*�5�z�3ff���խב(�fL�޲��g�O�(�3����}�`R�=s��!dӗ�p�r��_�]��݊������?r�6�����!M���ӱ����V]"=g��ޞy.`�ٗd��ly7�of�1�>ܹt�w�z'���8e�%~��e�t�>���e���]��˰�N]�=����/\�cS	��}g��_`����{���T���]�'W9-:���QT��fB{Y�_����L:0��.��,�i��<i��V�ˇ�w�'s���>ƺH|;���m�[�;��߽�ꭥ޹p^[./����U��U��!M��}���^����U��Op�
��K�s��g��X׹�>3�t�|�{��Y��n�˓��v�þ�M��R��C�nؠ�Y���}Hg����(�g�����}��������Kw��W+���+�]K>}7R��.��360T�ӧҔ�:c�R*����fG��{3�:�1͖��o�z{��4^��v�O�0o����ž�������Q]�gf׾��;{g��+�������Cf����%}�t�nṀ��:Vkss�_{fn�L��}M�M�ʙd�C2_f�����_��r�Z���៳Ù�����݆*�a�ȩ����)<�iծo��xf��w["����j��\�v������RSJ�g{��[��Vx�������7f�ﭔI�-�s�8я��_-�.�%��f_t�}�&�n�ՊR�O.e%s;�F��}qw�^����ͮ��dl�ݤ����+�N�*��wv�:Q�&9Wm���O�lֽжt��ɒ���l��ٞ�ݙ!��;�[ٌ�6�\�¶	&\����l����7�L���']�#�K�vY��ϡ�*��ܓӳ��Fy����a�t��dq�ػm�=�w55�������L���������a2�qY3;�o}��O:�x-�}۳y�;�����#��N*�x�v)�y���=<~���>/{})�d��97Z�c��fIp
���vw���w=�/�Y����OxrI��mz���1�c�;�a7�՛��y���m��i���(\�k�B�){N�g^j��ݹQ7�}�*����>[se�Ϣ�vA�ٿ�˽�	����*����3Tza,�Sl��<�=�l�}~���7d��}��|2�D7wc�s!���Ven���2�r�)�kwn�m݋�'����ƪ�z��իD;�@������*�*�)ߦ�eaY����޿.-V@�$�.d�>�w�ݗ��О�6!�,�#��cy>�Q���Sq.���M���t~��R,�J�6L�w/{#�Q�S��U��e-��s��u�Da�<��4�vT�k�}��7�b�$�ɍyw�T�寭m(�����Vaw&VN����������V�}�~~쫴�ݕ��;{�����if� Q�����au�����"}�^W�9�s��Q����`w�v��ٯ�N���9w�1�ʫad�n�v{
���m�͋٪�����C��g�>��Q��S2'a2?�B{�yc�_d��������~�_[�rf���~�%ŝ��<�'}�z�g�L�M�CLݛ�;���۹ݖ�LV=�נM�r�^Ϸ���S"r�=���7���ϧz�o�Hk��߷	�a�j˛����oX��˙�����R�����٬׽ifi�USɕWQS��5���k׽nR":+���}���v{ݶoV�s�*���n����K�����Bx4������;�/f���WT�a�Oa=��L��'�*���}��SyrR�&K�����%�d����/��We=:X
�;��N���{~�(�����]�K6'ҟY��xd�:~�޽o=�s���g��x�����;��Cq<�W�"�U�8�ڔ�!Z�ΞǙZ���͟�N���w증�y�o�~��e��e���x�E�n�*���r
��oT��ڽ����1�~���̯:M��oF$�9�q;ңW'��8�ٗO��y����+z��\V4����O_*���[dZ6��^��{2f�rgg���L�?]\�][����{5��on�9b�xMڂ�e�y���T��\���]���J�m�@��;6zqFY�6I$�fgGߡ�Z廧�����=�$a���a+���g$_?��gc��~�7��˶�v,c�a~{�;ޙͷ��,�ɰfd������8�Y�'�(�;�ɼ�;0�n�����3&��-\�֕��]�.U�3c�d�N��s7M��ޗ��:����(B�������#:����y�v7�ϳ='s1���r�4���X?��֦e�3�	�ᗾ���Z�͋Vl�Y��'���6���j���s���ƺ,��ȝ�sӧHu�� ՗:]{v~�W��w�b�욻;�Lgsn2�{6�K�}��G�s��������~��p����y��3�-��4v�[���7~�w/_��W/2Mg�<=^����ǗmÞ��������]�җ�-qy�����m�6�ŚK!w%fƥ�/7:��M��q�Lն���KT[�S7M\EƵ�l�F��o|����+�M��e�ڹ��o	Z8��i3;�n��Hse��r9rZ6���=����g*��.���Y�j�:�F�CDM,�2��H��V��6<e���i���6��kn���=�<�1�lZX�cF�j%ە�jx���b�t�@Kb$V����`s[4͖�,���ׁr0��,6㥕��a	�l����wë�O��=||��Ce-���'���Z�9#�1����3kל���'y���n�$Gh�5ƻWBc7jJ�u[���9v��hAr1K,!=똿z��ռVn�ssvt�c��w4��k��n�#��Y��f\��.%�ku�e-�ڲ�!���Vݳ�k���4�֎��W��{H����.`�n'!��S2�TȰi��W���]F9Q]M�DI�KG��2[m�jʛD�U�ͫ���R;%��G���Q�̂��Ě�T��w�@��[)UH�F��9�s[5�]��뱝\|*�������ڵw��]�{nEH�X�1�n/}��zR��BoX33屧)�����a�e�6�`�g�>B����\ek�y��]�Ffe�I׆�u6�S#s��me�=�3�W���곽�ȶ�#������S��P��zdf@���C�J�2�/tI�X^���m�bp������$����+�k��w)��\�2���+`�3LSOEN���������ۆ�.�&�cmlcD/���	�dc*��Ћ��u}&f)���>:�9T8��9[8Et�g��ۙ�������c�m���.�\U�Rlc�Y��LP�4/E���n�cZ68MS��{<Z�%�].J������rKdW���ohк�U���e��!xn���x��F)�N�ʗi�x�k�9,�k\lg��;{	�� ^\,�],�kK��kY�eB�Uf>�Q�����Ϫ�DE�����|Ӣr*�yU��nyl���M&�M�bb'M��Gӯ�26d���_]��Zg�@r<�kS�ﯷc�޷��ۯ��_������e5�\�x�#�����o�q9����Z��b�����b77eǐf���y�B�-j8 �����ƅ��;����$�k���8r�מӧ��=�q�׭��ޞ:�lv�ފ�7�]�x��n��uqn�����y?{�{w�{��`SfPel���������������m�m�m�M���[mͶ���m��1��m�M����Ͷ���m��1��o[�ۖ�m��ݶ�6�v�t�n�m�m�m��m�v�7|b�6(٫5f��Cm��m��m���m���m�������&�m�i��]�۶ۦ�6�o[M��|��n�n�M�����o[�6�xۖ�n�n�p����A��2�VH���j�ܶ�x��m���m����m�nm�m�m�M���7�f]���m�M���6۶6�orۆ�m�m��cm��lm��6�}��� jI"��!>d�=g��w�M��r۶޶��z��m���m���m��-���ř��|��m�n[m�m�m�m��&ۖ�op�m�m�m����m��m����j�X��Xem�ji�+m��^�6�c6l�%TRo��������=�yy=os������{��x;8јIc0E���H� �D0`�!�3��Y#0d��p�`�3�h�p����a�0�Q�$c(c�8f�A$��C#C�p�i#by)x�	y�,%,x�璗�!�2!�c�b�!�2�HP�,c1���p�3�#Fq�4g�&��i�8�	,d@�!�e2�q� g�Ǐm0��yL��$��y��e��y��oL{/ܘ�s>�2ʷ�b�c%�k�+	�}�}��㽝�#�U?_��A� u}��3/f#f���3������[:���S���hgm��l��o4��E��K�n�3R:�pU���krk����O�%x�pU[���oZrV�l�V�a��]h݂����^IU��D���L��2�!I��u��Hj��m~G:�m��l,]iYv�ծ\CՏi�Xw=�W7%]����="_��t{�xQJt�Z�-Q�e���Cl��p�;&�<��2V���b�ǖ�X�Ƽ��I����Ny8B�<<�J�4���
�"���������e�g�b��8g�~-�.�/u6�u9PY�N93�A5T�v����;���O���>[���T�1AeK�(=���5+T�$�{mő�U
����WQ��CJ@���v�x�di��PS
��e6:����ͻlD�֮��컬˸8֐qG4��eܶ��uQ��X�u{$�͹-E~���nc�/�65�E6ڦV��{$�C�g�{�_w�}����~�I$��{���ۻ��}�>=�{��{wwu��|������s�߮l���A��ź�<h�q�����qŜp� ��j{����R�tp��T,�J��X�b��]{���i�Y�m٬$Ӱ�o�y� ������pf��\WN���8�s2� K�X&!�.aX2�7���m-8�&Z�3�(zp�Ρ�~���>-+F���6F2s09QC�}
3�cS`w&�F��!=���Sm��s����!aóÇ���Rw/B�<T:1g"O������V�8��Ym�Xo|�����d�G����M4ў4�xg`��'Y��GtJr�V�
+�1�Um�۔M>:��E�[9���{:[t��<:�!�=9�J	ڥ6{8�o����
!N�ZK�>��G
%�Ǌ�d��L�b�	�:�	5&Ȼ`K4�2�\I,�GbM`ޓ:�+ɪ�OJ��sm�3QE!�zwI�a�i,C��e3Fh�q�����qŜq��h��#�b�s����vn�,Ib�"s��}��|����,m��C�J	�f�!��Jԫ���o�YI��<��Z�,��Y5+���aiK����pӳ�Q6$S��9��bv0��Hw4LN#9�	��G�����au�&�Yj5Y���#�5�����4���4$O�IŚ1�3F3�0fd���,�iU��tܠ���8��>$�JF ���_�3��UE����im��E[�[�V^(��!��ܕ��ʰ�}'zpksчq�*/��7��9φ�8N���ò��a��<
�a~|��JR�a��P�SP�-���:�<�L�#$�8c4Ed�d\���X����ӂ���dǚ5��� N�A̵���K亯�s��_MG�/:���i��m��T�� ��@݁ZKń�j5̠ȶHҤc�.��Q�V�M�r�@���@�y�
u)�f�2��޴�r��O%���p(�o����带V�aD>!�2C��a�u��$��!�a�����O��fxi�C�+jMM�k4Z�g!bif}�@+�N�X��]-ݦ*n�M6���}N�s�C�f�����a�Xm�uǞu��m�'Y��&Wצ!Oҁ|n��N\��&ˀ�k�AI���}��,,4�凐�BXyпߑ0ˆ7آ�U�b���m1��n&�$�S����R���V��ae��4��S2��ȇ�/��}��:;���h��M=��*j�[��yh�&�z!�@ԑb2`�絿Ca��A����3N4c8�`�H�8�����QϪ����+������9��}$C�a�E�z��!��B�T7�lR&�T;�7	f%���F�T'UE�X��-#�U-@W]�9�o&����ʴ�c���6�Xz!���m��8��30��p�Z�&b��-�#f�x�N<q��q������qŜ1�"�#�����(3�ƙ����|�D� ��~,��\��D�3ǭ�#��D'N�f����y��}=���_�8K�k����?�S��6�&����2�R;�kѤ8xw�;�����;s8�Η�w��=6@�-�.\|H�>,�4pv��"0�gxgX��'Y�0`���]U�]ޠ�;�|3z�r�5�l9P�8��5�Qي> նk���X�]qi����$}[r���e�%܃T[l��"�`!B���,�'b��� U[��lp1Y���m��ӭE,�U!'U�I�E' R�,�����a��f;>���j�<��Ä$����2֙�0ܡ���J��Q��RS��ϱQ%���:
�O"x?����J��;���R۪��G�g!.�%�76��s<�-N~��3&\qB�FDɍr5yQ���^�B�u^{��p�yܸa��<k-��Yy����Y�M4�ǆp�4��1�2N8��`�s�H�
���ȱf�h��M:�99�{^�6�p�SUXy+r8b|�c
�LN0"$�B��ER��:��4g����\��0����ł)ܓ���	;�s���1s˵ၒ�aja\�zS����hxl�gr��O�\��TTh��&2%�ɦ}������ȓ�3�?��H�q,�^#EFB�5S<M��\�2�1;a���&˩�RՄ۪��kV�[�:M��-XNSi�V�Z�M��uKO�4�8�6���)6���NWSj��Ŧ�[M�
a�a56SU�l[*����q6�ylZz��]R��h����J_��SK�����ɖ�q3j�+�*�4�
�*mV��*���mV�[�L��,R~'�~O����->V��y�J�n�i���kU�����y�|�6�^K��?&�<iT.�A�q-2�0�-V�NSj�j�nT�ؔ��<V�iL��M��LM�ԥ��0��
RSi��l1i�m6���iV���㾕��>N4�ST]ʙ���zvWu!,�������S׼}#2�X�>���^�Z�1��4 �o�Bu�:G�̈j���=����@�>����@
��6����z4���;�ѷ����^�z��`�����v�o;�)z�B��'ݴ��\:|N& �����߇ ����_�V0�(���3"�\���=މ��.�Z�|��~.��֞_��~�ԕݛ�i���!}����ݏww�������{ۻ�����{����������z=�{����ݻZ"ZZ�[n�o-kyƖ��YG����
���T�MZITDO	@�E'�tY9�u��hIP�D<�e��O�CDFC��x�����qtI��w�X2	�[Z�:���̸i�0a���BȈ�u)	��CXl0�,�DBpD���qI�S9 �@W-vZ����jI�S5ZNaI�A�H珡�G�8l�,v[N��Hs3�M��U���Aw��$��|u
0��bQ�p�1�L+��I��@�d��@� j22��cd���o�n!�I�4&�D&��:�%��P�R�I����ʅ$�LA�O��Df6��yן<�έղ����u��[k^.�U*�U+2��FI��?���g����!��u�,!x��0��	>���L!�&&�)S��>.�W��v���K{4�BͪG3.]��v�A��	50DO ��Z`�T�2T�%I�~r�8B|�	�J"1  X2�I��`�NDM�� �x�TF�i8�t T/�J��h�q1
LJR���"P�r�����G pCS�.I���$�" Vd��a(!���}Zd'�}�@�C�԰�"xc`L&�<(c Y4�RjVO!�D@�"��BM&�Lʟ6�:��u�8�O,��J<P�`�{���3J����كC��J�Q#i�d����c�o���Gǽ7umzV=�0�E= ��R{[y�2,������K�P��E�圶9XBZ��Y���f�1)�9g� 8B��,!�N t�ׁ�61&u���sqnB~�x$�c&[`����`�@�������HnX��YhZ%2��#
�Ԉ̑�I�ï2���e/���C�4B��%��v�I�;?"em�M�m
��2χ��8� �&0�=�,&�zÎ�I�\���������XiC�r$�����h��%ē�&�,`}yAUKѧ���<r-��Ј�iJ����2�;PL�f7`Ɉ(,�@�����F>���2�\ɣn6�p����!��Na4�=VN�D�PȒ����$��yȖb�d���b�	i�[���zg�0������y��[k�귄�G���1$D��� ΄�2BFSI<�M�BR���G���c��e1���c	��DJIϥ!�d��a.B�dgBk �>�+�M�`��aDD��;``��a)�	�����e(��!FI���h���pB����r&f"bV����i��[yL�SپO+M9a9�N�
0""���Dz�i�k�,RZ�&.rd����a��L,d�[ Q��,0DK���h���v�)���k�zK��)'�:��q$�o��î����`�
ihh��;�~���I@�2�2b&c3a/%O<�Ϝ[�μ�0������y��[ko
}���3��:��U��a��aȁϻ�rC�n��`��"PHΊ`��bT;����2L�� �ޕ�>��¡`��#;D�$+"'�K�2x�S�`DO~A������M\-��5+����PĞA��<�M2���(=��)K:e�`�p�ⓔ��m��2ۜ�O�(�#I��� щ�"III!��L����(a�&��u�*\k�g|�b�%�}/&@��R���:�"vY<�CY'^-=�;nf�����s2��iDa0a>H`�e��9,�	׍���[��a�0�֧��~<�>~�:�8�岵���y��|t|vp@��1���I=zz��wk�o�U��&��0��4���,���_��OǱ����FAQK������"r0����d�)Ԉ�ʄ!~��e���\��`�Ʀ�8f��7��o��O�K'�҄DXzm>�J�:�"O"B��A�	��Y�d������C�!�kт c"�L�m�`��w>�d��yG�m�c��K�pJ��AH�z2)I%���G�C���й��O�r�p�\�v�N�?D�Ȧ	!P?�p���0DHh��!QE<�$��OO2�{4ф�A?~t�$�C�'\(uA|��>R5܄�Fa1�PL��o�q��>u��qK[+[���m��j�����{���q���%��kˋ#����pݶ���3���ym��3�IKìs�9a�ck(HׅG޷O5�$:�����S�spc I���]��٘�bݲX���VS�U�c�\�(�,��r�@�S���S��b��=�H�<�re����3x���SM���DIជ�9��n�՛�,ghݣ��Д� ��$���m����I�CJXwb�0��0�D'�K�d�� X'���Ӌ���.$�a,)HJ��I�T�J���~�E�����bK�E�ʜ��kZ���RRj|��`�Ҟ�E;?o�����dM2�$2�J&���G��KN��C���}y�7�i�y�m�p]��L9I�Fr�����+%6�	������,R���N�am<�-o�m�S岵���y��񇇽{D�OВ��ju$�����B�,��(o��L:"A�]��L%Ĵ�0Ҟ��W#���ϙܘz!D<���i��,#iN�(�D�%!����D��FHC0�I�L#R��f��e-���Q���rS4T#*b1�pm#	>��Y�O��l!ˑ�X��`��u
w(� ���ha���̡��
NA=�ġK�T�~�����P�m��4�d�)�ې��$�҉��E3�{̸p�bX%��~:9$�v&��$�*q���ζ��)��Z�el��o-��1U�+LM*���8�5UbD�����L:J)*sDnI6�!,�Qp��4ttR\\10DC|(��tj�&�*Ip�i,�2��S�\���&"�h�QP0�bl�F��7sL˜�:"Yᅞ�F��H������n8S��t{�{�6�)�vS�>�i�6�8��d��~73Xu:8��xxi���0�y>U���g<��:2D$�v{)���ڒ�E2�T�a�&r�j��-�|��|���m�>[[���m�|w^�ۅ�l-��w��Э�G/<UTH2iO�=�b�u��ڎC'Гp�>aHi/�Թ+m�	�B� �^}m�����0�˗2�&�����'BN��;7��O��Kqb5
G"JK�&�ҕ-)o�ӈ�4�C���aԖ)Q܆'(}�Ҧ��~孵C��~�☚\0��
A��C6a�=�2�=zS��P�a٦.PL�8"<�'g�C��J\�2�YSLDyc��y��CJ�
��q?-�|�&��<�O��6�)Vҝeli6´²¬�-V�[c�����km�uV�����ʴ�Z^J�V��&V���[�[���m�y�[
�mj��i�kU��&�VS��ɶW��ͥ���U��M�lZz�M�g����p~0�~>�Ng9U]*R���v�Nl*��R�­,-V�j*mx�U��Sn�l*���|~����I�E�����)/��I��5yj��i�m:uY_�������ѩx�:Iҗ#�b�q�L�6g�JU��S��婶n*�^&�)������~�ڏ�c_�'���:=S�X��Oվ�~4���p�<N#ƌ�{U��ˡU��vE}H�'4J^ڛ�M������35����ަ�"���PZ[S�ߠ�!2��+��m���44R<n-�G��w#Ok�:-n֊ n���.�يb���Ac��)l��]
�ɑ{�{փ��9j����H^�3�^j.H�\��{"Ǚ�
1�?�ܦ�ƀ��,t�W���~۰W>��)j�yú���wm�rşc�!�!�h=��߳1�6:�LE���X�kbd����RԺ /�g���'��Yb�X�2��s�[�J��f�轟{-r#���mď9\�I�r�5oZ��C6nSuB��b�w���ۤ52,����7�YvH������cI��	*|){����꽗�����&A��/7���Ɂ	�� �ߣ�N�c�d�����+���}����6�xt�q�ڞ�ug2F�m�o�W��lRi1�5��5"��I��ōV��+��o�X^�bz�O?5<dF��6�8�rW[s��Wy�q��>��y��P	p�e�?n�oG,LDҍ
SUd���dK#�)�x0�O�b�i��ǽ�3��M�C����m�V*5h64���e�[ ���9�ƚrN	����jw����G��D�"}�"�aT@n�b�K��h�`?�~���ϻ�ww���~�wwwo�6�m������m��������4c�0g�x�'�(c0g�<MCQzUUWBUu0UAL�Β��LD��'kl���(ԣ��r�ͪ�!�C[!�˥��`XM�Xwv��f���q��Jp�����t��Hn�YTR�Y�T�r@�J� �(��(����� %��x����(f
K��k�t�r��crøl;�1?~^A9aL����=�9���nC�|�xz�3����̇���f5���QM�����aReQN[uJ��I�a�ķ�'Bؘ���gUC	߽N�)J^r2�Ɣˌ��>��(�s:�-e凉���t��j�L����� i�=�Gg\\=�R�D�r�Ɲ6�m2�N<���:���x�ǉ<YC�<i�^�Ip�^�^�� �O��6���b2��\S��E�3L[t΢:I��V_Doi�l��;RΗU3X�gP�%!�O{�ngG��.fVei��[
���J���ħ�'�\=@�vO�Jǖ�FSW.�,]���7�~=	��Oߖ�NpO�u�P�%N|k>b	8W��)/�tnB�&�L�XS�>)��џ��X���x�'�(c0g�gǠx$�@�k*zfUUDΗ��id$OTDӖԼ�:�}	�*yȆ5CޔO+:^S1��P����Ag�C
z~�w]K�����1䜑AAT6�-bd*j���S�?O��N��K�<2s���Τ����'�)����(ÿ!�\�a��\�Ͳ�-��)Ŀ~0+Fp/~J��g��Y[�[�[i�ϖ������6��q���R�uUz��������L���&c��j%�D���}�8�>o���C���O�M[G&ծ�vs�h�U��D�a�$����=��a�'R��c�e�Y(�z1���~v9$�SnC,��7�9�ӈ¡O���jW2�s!�����{�?B�qi6�6�F�Q)v�H��1�)Ӟ��ڗ;�vt{?Ca��k<,�}��"a'$�i�|�[i��Z��'�(c0g���HBPX�.*�Ԉ+~@��d�4��o$Ǳf*L|���7J�%`���E�h��	pV�_���tZs[fr|8��v��.v-��h�KbV��ho�` ���;�*���W�q�QS�R6�&5*�z}^�=��A�p��Rh}���ۿ*UU2�
�]2\=14�Zs�"�4y1��L�2�Q|�dڸ��[Ҟ��P�%5T�U&'aS��zQWóa���;0��%<�Q���f*i��7ߕR�\6����g
$����i����<p�>c����~/������X�ưZd��?M�CgХ
�:��~�1J���0�j��2ۋ[�m��>Z���/<��q��V�>MT��̸̤�ӳ&bKq�
&�x�*��w9z;��	��-g<�JԻ�������✎S'�F��I�7��++N���f�DC�6�62��d�&n8�nk3���Kh"��]�V����p����(i�RT'Pʙr�G�d�a������Rr�V�m�>�N<��y��m��>Z���/<��qý�xou\:UT`d��>=���m�J�I�Fq.uL%�R��X}�m?53�;<H�_ȃ
y��I�f~=:�
P¢t}?]٦fn����
]ʂqvX��Y�r����?K����&>�.w�a�}隖c���e�R�\NX2���-7��{mo-������N����[�&����Y\�1n�S���3*���塌C�r9��6�ϖ�ζ�ǞZ��V�/<��qq���ۦ���p�5UTCa���?rk�cx��̳3�>}Kũ��lr���4��9�m:[yHAA+	m��q�H��*X���Nj�j��>X��g�~;��f5)��rxt`j��\�ݍf.��J�ð�C.q�D��XO�Wz����p�MD���rD�EL>��)����L`��n|Y��$��P���Yo<��|�m<y�kem2�ͼ���/����_\�"�B�kq�+����/��:n�)Y74 �6�f�$-���-{:�mp�����P�XM,������Wl,f�6n�	} w��xM{msj�ˡwb�m���GP�	�Ly�Ӵ�_��}ST�.�[>��g����P���"�\J{���\���Q�q��v0�L�����K���c��e�4dk�|����k|=�S'Bh~�E9�_O4�u~�z���w
�E=����G��vM:���zvd�LӔ�0�7bTN,�/��g�O�<1��0���(�ef����[TX�i��o.`���q�R�?n=^��*��a���$ӭ�D�ߡL��Q�6!�L����񍬚U490Ȉ����2����"Y�S���`{�_0�ōu��f"4T�3�ku��r�94��>��Zi'��3�n�0Q0�lK]B��K@����u{�T)�&���˟8�9������cΪ�+ɷU�����-��U��-Vҭ�)�K*��+U�V��㉶�Ÿ�M���Ӆ��^OV�-�<�f�YZ��y���ۊ�U��iӊej��J��mZZش�kan�I�U���&ɵ��ղ�[6��3���kU��/e�Զ0�Z�u1�tS�x)��O�|R�ej��Ű�0�aV�J�^&�Ŧ֫M��aT�&�%���p������B�~'�B�</�x��=)��p�<q"<i</	� ��(�8\x�'�+�W���'i��b�k��aj��iU��Oas1j�x��MT�R�'�TZ�m+)�JJ�JV�T�T��G�?
�?b�,?�ZP�+�k?LS�n�Ѩ�߄e��uέ���~�\�`�=�K-L����,��f(�$�!	{�S���}�*�Si2e(I�S�:�7wg#[�$���z�ޡϥ�wE���,>9�a|�����1g���'���i��-;˭S
�e��4�������o������Ͷ��wwww�y��{�������m�������1�<i�<q���x�G�(c0g�7�脒Q~�UD<�?�Ɲ���(rS�jCN}=��Yl�L�b�؍��!:Y�$X��4=���}|�"�O�ߜ7r�3��C��q<9C�4�PL��f�ڧB�ɡ�d��@i�9�d�)���30p��C�ß+�Zp;����)�~X�0,��Z��&=0�i�ri��qk|��i��-K[+i����q�n�U�E{)\����N���T���J>�<����-���2�̻��:�aD�*h��:UUɹ��Y�Ӡ;l�.�ᙏa���0Ϊj�gJI�x��!�C�hr�.EO'��C�}����Kz<��{J��hZ���s���}ق�񶓿C'�G���1�q��ٶ�q��<���0c<A��,��0g� ˙H�P�r��&l��4TT�G �Ns������U���� s�Fq%i\|�T⿟6I��Y��̚���������'_6z%�8� �����~[��D�1)mM��,%t�2H���*��tB�Y2��o� !.���>MT�V*FRh4E�tu#���,H�4l�-g�1�L��!�|��D��u���NvQ
~d��������<��s1)��i�(�n�̥�Te�Z���$��9gg]Yl�N�Xt{��a��'Hp`����p���)}�\�/�SW��v�F��lJ�bP4y;Iؔ�"̨�)īq2��&8�8�ĢaGa�q�6�ǞZ��Vҏ��4�IX�R�)$�i�$����0�j�3���L8�*�\�x�g"T�ۨ��%��Q��E�s\g���B�����p\q�"%#��@>����%<�C}C�_�m�������M��ͬ���<�M	�K�����V!��uȘ`<��0�j��0��K��o�f#P�m��m�[m<y�kel����J�2��T�T�I$ ������c6̧)I�a{L�b-*`�0��m$�^L�~��=�R]eU�$,�%l��Q�O	��g��}���4�M�<�b�ê`�%$�^�a�T7OL�0ѷ��bU�#��܆�H�ɿ�D�1ٚ��DqM�(�2��%���D��V�����<�_-l��V�o-�51,��]��UD===�x�¢�RèT=4j6����V�1t�)�2|�K�_#��BR:R����0�̙[��=���
 1�/�R��}��tw�5�?Jp�L%(�}5\h�ZnaG�'
�p}�qwWN� �FL
<9�׾K�c��q�������<ʚcS9��\2mKen>y�ʹ���Ǌ<QG�`�wx�#�W��o��TU�m����q��T�;6��El�n�6t�5-��[�4e��o{&ؙ�i�sl�ۜ �u�[G�3X96�n7:Y��r�4tj��	N�Ya���q������YXw�����b�[�x�S���&�q0�r���F^�v%�=آ-/7
I��un�;h��N��ۆRn��V1����e�p�f`�Ɣ�����33;��7I�]�
���7n�M���Tͣwu�I��:)$�$��S��NaK��Y�`�8f�0���x�G�(��=>;93�Ȱ�`��&3Y���ڪ�u����,�NC�M��>�g0ӫK3���C	wjy,�A,�DN�m�����'�E�e�􃇺P�_g��6�뺻���:7j�)%i�@8��Z������{m��S$�	���!Ϻ��泭k<��R�qKa<�GY4`�5Cx�5�c[mQNC�l���un<�O�x�G�<X��G�֔��D�
}UTI�rd6O�8ys�|�W32��%�YL��K�J�V�V��+�w�tvHɎj�?�
aȈ'�>��w����8��n��U%Tʕ3-=�q���X��~���<�{��N�Rñ�O�0�Q)��ķ�J>��bg1Ԥ�eq=�;�z��w�ˎd�� ���Q��,�~yo�~i��%��l����<hЈ�iD��J�i
R��g$NG=\U7ۥ�9���� �!O~]�ɰ�>cp�!���)_i�?�ᦚ��梒RȻ��X�Z��+��Z��'C��ӡ(��!�@�Æ���ѯ�ߡ��bXaGtp���R��≯�4O��A������Fw�u�����fa�:�4:�?qDL6M�T����_}s�]m���\�-�X�;U�6���m�a�Z���<J�R�i�Z��0�K53e�V�RضU���l[�����ԥ��^K�U,��Q>�
O��i�<i��.*��l��V�[�Z�ժ�VSi�p���-V�ZՕ��ml�Z�6�v�bV�Z�Kc	��V�Z����Jj�iI�+L�V�[
[6�eXaV­6��V֚����k�کj��ŪV����Y�����>c�bk�>uYZ�y�[Z��t%ǈ�^4����a�IF�ǉ��QҼ9ZF�b<�'��YN��M8�z�6�<�'i��ʕ���|�aV�VRV�L��R�\����m8�V�>c��:���ڙ��ެ�s$��U.�fF��޴j�(��:V;(���q��6F�4U�M�Uo��	�����qc�[q�fR��L����ne�^��4�0n��&7�k�+j��6dN�0r��S�J<k.+�O^�x��S�ɋ&6�Y��*��m֭�a��7)*�n,�5b��	�J�j�n,��ٸ���mO+�d�j�-O79�Ӎҕ���B�<LAoF��1=U�߲����f"�2\�׬�w�2��E���}4f�ۮ�MM���_�y}�ڇ��=�)(�>7���>0�o|�+gr}��+���b�vd�ͬʬ�fAU��n���f:`�1�&�M��2��g�j�٩ڮ������{[q<�r"�*q��Ʊ�%�ne���u�SVS�����R۰�P5�+{�N޶X�͝��Y�SY��1{�wUWW������xp�ED,4d�?m�*�e��R7-AI�����7$p!&�%r�!�'!�I'Wj�[%�1��ƎlU���3��Y��������W��̭���@�ޛ��CR8�-�rf�:%�ԭ6�td-��)�$�U�!�,��JYe:#ٴ�kXSJ���Z�O��_����w�www�yy����www����o��������m��www{�P�0f�g��b��(�c0g��ԕE%bC��R�ZӘV[.[̵,tQTYN�}Uc����j����1� r���Wa��/Q�me�i��kJ��љ��%j�(�py�Z�䏌VI��?� l{��h�®4���X�0��1��J;�a�r�ɘn�j�~;��2�1�S�v���9$ᘮÚ�����[�m�L�!��l�ffe/77�c+�a�{Uӄ��v�|���J�i�r�J���:���.H ^.Z��J˸q0���4S�d�ia�Yn8��/�>��(0政�t`�<8h��.��o�y��<�^Z�[+i���u7�g�Z���
\�S�c��xQI��W��<��M>�b:��mOd��,�?R��m>{=^sR�Ze�6vx{6Jr~M8%?I���H�Y���g��CEo���!ZLͫV��-����Y��QÐ���S���Qp;�����3M�5�"\10ӍFP)ӲL�>����R]I��3�X��C<x��,f����F�j:���~�UQ'�2ta����G�)�e��ɷu5�J-1��JfTç����3��FM}�V��כj�iqN����K�P�"��0�R�����4y1���Rf1�'�eE}��ĘI���؈_�~6PO�]bރ�d�W�~���<73iws����eJl)�М����>q�i��%��el���yn=I�UԪ��333)7
T.Ogx�����+a�y�x�S�$!K��I�K8;9U� }1�!��K��>�G��\����)�4�_}ZF�o)щ��²�$�iRLB��)ED.㪥/-Sjry�C���
b�җ�L�#Q�J�iq�[O����I"8Ӌ��ac1g�<Q�`�G�RsV����:�b�n�ɋx�K��lBA]܍��+�rI�8Z䆔�<�#����e.ܮ�%e-M'Ҭ�kP��.��^5-j��('	dr��  ���b�KGd�m5!��l#c4�&������NCҘ"aD���i!yw��_\�u�?L?;�O'��-15�\L��0%��]d�^ϟ5��S,#q���a�t��e��m�UU)�3`�����u���c}~��#���Q���.�74�f���Jw�(p$;AcR2
�Xfy�K���fҋ,F����3�ac�^yl����o-Ǖ�&%)��⪢D�~�Z�P�'���ˌT��6����NĲb��^��OR�e46z���ߦ��՝����P�pL�������N����������~��0���v����zպ��ۉ�m6�	a����_���r}(d(��?JgQN_}.	�d�R�C��3��ن�JI�K���UL�	 ��2�i����,`�!��G�<2��K*�©LTDQ>�UD~������R�g���i�LF^�ZXI˟���暄���ƶ1Vr1��d6N�(�;֖��&/Y(�
|�$\l�PEE�,R�`�ߌSؖL0��(�fe�'P����q��2�0��)���pg���2���ӫ,�즆������P�c���>�Ð�NC1N��uJm�����1g�<Q�`�3��'�U~����Z�?*� ��F
�~a����0v��y��a&6-�i��h�0$N)�ʈ�%�S��%��ޮ1LV�\0�ģP�������f}�F3��f��itv0��dwzi�P�v����p<�����٥ ��	GG�[Dǯ�:>� S��l�c�B\aL>[ξu�m:1�c<Q��x�q�P�*"�"�.c�ʅ31K1��&��9Vs5��̍Ac�`�cgM��0w7q��1aC+`ӎ�����R:l��q%h���[b�ِmS�k�J��d[� Kru��f,�l҂�R��%�4�Yv�Z�f���N��c�<a�p�;5���v;0�������X�v~�NB�b���_CN��F�4��l�g������Ъ�~�0�e9�ڨ�xQ,?$�LM�}}:��
�j�Ḗ��a�C\��7��O�}��~¢j��v��`�bk\*<��i��_J��L���'��q��38�1�(�Gǧ�O����֖��1�ɓ2�F)$�	���Mwr�3n������k|�������ǣ�y&���檻�ˌ�)1�gP�!&ۇ�JS?iil��%0~9L
\�t�R�c&䲊<�I�/�����ؤ���i�h.
`���?�;�L��4�<?�GF�r7���N��j�=�P�ODB3|�)*�Dq�#���y����[�V��eո����`�R^G�4��K�0�̘��4b�c
8g3�h�(f1�Y$�8�c��d��0c�H�2�c$c0��`�@�!%@�b c$�@�1����yIx���Z�[ek[jx�,g1�3�i�4���h�0g3�8e�ae�LL��o	��(a��#�I����1�d�
2�X�a����:�׼{n���L�};#��3w�"�45��8�2Xƻ����?��"Ԩwd��;zE�f/nw�ԝBâ>�\P�w����?����[�΁8��M��D�i�:*4����ۺ��R]%��'���=K$�5�D��*�v}�������{�Ͷ�n�����z<�o�}�����m�ݾ���{�<A�1�38�1�x�G�Q�<i�c�J��)���Ԧ��C�j'ffÇoϴ�bYa��&N��L�μc�fe������JP�Չɧ��Pe�%2�y��{z)����-��v\g��p�^l��n|ry<+�tȞ�����C���f���'aًa�u�N�r�VӤӹ�Rs���x����S���Ev�'pN���ø2Iqy��W�AY�1�3�Y��!��Ǌ<�o6�#}����e�R�/s332�`��뙐�n�����~:�G�H��HN���1�Ͼ�v���K���i����v�.�t��!�3����5J�Ű�%�m.Í�W[T7��g�u�\0�T-�*�,��R������lц�_3F���!���c䶘�KF�36ܜ<.D�d�g<�՚rx'��:;in�նӧ�K�0����y��������^�5�8�@��թ��ӷ.���4.�u�n�e��c[m�kV�j�5f[�d�Ԍ�-�\�X�Բ�pV�n���jw7�����]��].1��i5��� I��V2V0`�*Y+iex$*�r�����3�O)D�pM���hu'����L;B὘7)�G��)�L�e�;ɇ�C��'�ޢ��G�ӠO���Z�h&��>6�U(y�6��QC�aߓ����D���C%60�����~yx���wP��-�Y��J���r9{
j<�C�;
8�.j���a�:ۮ<�V�N��^'�xf�ƞ/���&fKԒJ!�g�/�3a�`'�~{�h�f���a�C�p}�:�$�L%<&;v=}J�����P��~�~,�s���9�Ɂ����b�"9���j�Z�CP� B^N��� �Jl�t�-����)m}��!AN�C�,�4�8�����Mo��m)�ͺ�ξm�}3�����m���Ǒ&L�\�G)�+����n��2�C�PN�c}��'[�a��m6	d�"]�1��*�����p�(�z#�&5����&b�v�aJ�3�����
��5t{�����Q.f�ꪧO�%��N��-�&D�w�G���)䞅�Xa����Y:*3	z%l6a��[��38c�H�xc4�Ɩ!_�ʗ����I�Xy0��5)U����$��	C���b+��T\-�5��E.Y�aèzS��C�"y�C�O������X<ԧvgc'F�0>>�*&�)���ty�'k�6�
:�#�b.���q���yv{�P�r`�Wg��Af�i�����@�H���X�.�G\2��}Hk�Y����"�MunZ�C�T�N�WM�u�l%~+{x���wt�S;$65�c�V����u�Kn����0��qY!0���U�u�5,�Dk�{� #)���TL�e�b �rÎu����CNq7��c	Z\���N�ϔD��h!�7�S�wmf�����-;����p�¤l�G51�K�9�rm��7��o�Le.�<n1ʆ�"!�0����Uݹ˶�[*��Wm�V��Ft�à䒓�����DZ،�h����zx��<ac���f�x���_���ʟB	��؜Z�U� �������P���y�)�7�8L9;L(�=,�L��&'pӄŻqb������<���t�}TE�#N���m��qf�D�F�NS��O��	��h�\54v#6n-ilJQ��p��R�*R�3V�iԸd�BwJ���}��-2��g��r�|��yg�����@�H���,�wϩ��:ҟv������I� �}�u�&p�ܱBND�-��K&ap�bf"��Y�1p�z�9��c!��N��G�B����V�%]��@e�5�D|���!%8-H�u��7N���a���:�I�E��������0�5zԝ���*�RzS����~C`�G�fӣ�$��8�q���p������-��S)���a'��J�RL�E0f�!.Vڋ�r��2**�D��/^�� ï�c\:4�a:�9��H|T�43z)�bJ)
eˋp�1��*������񧽳�RјTf�̣d��$�To�R�m0�Q���K*��&]����Tv�;�%����0�2��f83��-I��g�!F���*f<�Ƙ8���	��>}X��J�e�\[N�םm��m-�m-�a�%e�����y�y��m�4b�c8�iH��0��c���8`�1�gg�I1�c$cc�3�e�<x�IyIx��2ʒ���!�!�!���c��3D�x�疶��Z���ˏ,g1�3�i�4b0ќ2��4e1q3L,��#C�0g`�q��0�c�����3�4��&1�1�b���.������f�$�����pi�p�[;:�Ae�Z�+�{B�-#0j��y�a5{�f��e���K�#�m4je6����z\�⃩�?qan��RvR[����\���1�� lK��˂�U����5��H����M�j��y�Y$b۸��Y$)��Z�F���f]��[C��BvY議�AM��^Y��&�����+���e�u���R�gLB�#G��E�Ѳf\wӱ�����J}���f<xsdYT�ܳ*u��O���~x��U5�$R����!j�a�lB����i�rnt��^�;�<��d����_`la}�W����$�r@r"-��~ܹ��}p�S�`��9��Ȳ�F�U%���~�U���vN����9{�"w2�o�U�"km�f���ںf)v�r굖�f�l��Ҟ��1�����ڼ&��+i��T嘃Z��_k��͑�WSf��&�Դ�m����%�C�6.���͎Ԛ6�f�i*�惼���i<Յ��z�V���U��EL��jKD�f#t�5#aA��h�!v�lqf�K]�����ލa��%UEx��NVn\Y[)rHDvP,j[l�Q]jAP�'�g0O��܂��;7��q����~���������m�ݾ���{�������ww�������wv���{�<x�xg��p���f�xҌ�5;Q��1C�9���ț��5�/5���X��/
)k�]���՗RA��Sa1���5���*�e�i��]7
#5Z��&�Ft %n�BY��M�*�x�Q�;iV�X�1g!���yN�8v5e�a�)��Պ�c�[Q�Z]*6�QơL%G[u�أ�j�a�(���������6M%&�=72�X��L8n����UX�&K���uX>G:^�C:���(~�~�ơ�<��"�����JQ%��`&�����ړ�04;)a�N�T�x&H�?8�3�@�$���Ɩx���y!X� �r٬��<���r�0����UD2(3؞{m|�G�D��������j��}J7,�{�CO�I�X�P}�a�	ih�!�<��4f:Ð���C��s�޼�ƥD�v^ZES��+\�?|i���
e�A�}���d��K{N؊i���7�f"S�j�5��+0�}��1ɟ0S�X[�-n���2q'�Ǎ,�x��"T$Y�@ BW���� �C~Ǆ�3"��ӱ�O���{����0::T�4��ٍ��'C:���e8s�wߢ��u�Uy^��k�	�y'>O�NCl�a*T�b?1&�)�ssp�M���p�	d��=Jb^��cI=a��U�6���d�L4ҡ�e�������u�8��3�Y�E�~�R	�Qr�%н*�!��w/r�����<<
!a����,>0�s+�`��bk�Sq`ѧ �g�47��}���������<C��2h_�4��6p���8vl8!�<�M�0��9lz738���X�z"aM:r!�0�����c������μ��d�IǋǍ,����
�IEѼ�S�z=���X��L9lf�y��\,#��{*���Qh��*���a(�-E��Y�Ƃ�)V�)lf��xC�b�@���B3WmZ�Go�� !%�����,<��AΫH�Wl�����n"�ÇBr�SO���2��UTgn�㞘L���q��e�}Q�L̢��8�\�����*��h�&&ik�ky��6��p����:|P������pC�*��`}�߸.e��T���#�������t��,���~�m)�*~$�N,�ǎ�8c$�N<X�<i��ِ����_nێWkҪ�#
��Jf��MGg2�Z�|��O�vxS��q�υ��h�WC�k;Qu!ux�U�ԿC�6�b��I�q��-�̚_a���}��w�^)�p�k��~Ǔ��.�K0�ffwF�S�J���~ߤ�X�
~4�Î4����'q���x��^�'H�
_�2��J��w#?S �{{�a�h��!�N�������~���qo�C&�~,���o5(��I���`�(HԎ��c��6���GG]�R���Ä��Æ�S���uSq�5�e��Ivnv{ne���r�'���0<�.���zi�>��N_Ng�p��UA2�(gg4gd�IǋǍ<_r���%��4�K� ߢ-r�c�DJ\���2�m�v&q��>�~�^RX�(�3na�YL��r�'��
J�")xa{)�-���faKjfZ�Q�S	G���
�Ɉ�`R�OQe0C����zK�DyN��|[g-	m.�jFѦZ��0ӊ<x�Ǐ�ƌጓ�8��8������)a��(�>��M��0`63�X�0��k���;�����۶7�m������T6I�d�2� ^e&�\�n�Riunf�����M�E�x!��Y���!X�,� !<�Ĉ�(VU B�BR�3+c��m�p����{���b}��\�����N�=�i�N�.������dX�SA��~�W����N��4Fw�ķ�3�9Mw:;`�`��/�v͆�H���D��R�Y���\70��h�h�̍t�8YJ��������I�Sm).��E1�̶aFQ��ƌጓ�8��8񧍩���H���(�(�"�bP�)�n�pw�z���}�㓆	�/���&R�q�øtw�N�FR˭C�f���ʆ[�#UU>m�잘�	=�D�K���&S�&�>��{�L�j�
��Za��E�й��3B6��P��n��w����G�C��-?	��#�ޡ��w�csC�Ԣ'IŚ�j��=S9f0���b��R֜/��I��4��4����
,ag�y�0▥�Zҵ;��[L�(f1�3��p�3�4d3�H��0�ad�!1�c8c���$�0`�!��&2�1�3F`�0d�d`��IDP0c���@�1�f�cB@��C<x��(�ǌ<xј3�$c$g�Fh�a�8e3�h�q��0�G�C,c0f��3�4��"��C ��Ag�b�$3X�H�/�=[�Z�L۫���ϑ�B|0�)����1�Z����j�V���b�9���OIF�o^p�]�DBE��=�v?��,A�~t��f�՟;}f�>��m��k%v�n8���7�8�κ�"o.,�x�grڕ5��o=���sq��iv)�}���s�?-��L�*���ɩ�7ڠ��y�������{������ww��z|�}ݾ�����z�o��������8��<3�3�2N$��ƞ"I'��V"Y���Cӯ���U��=��p:��4O ��?�1�t~���|O$��DȞ�ΊQ9ã�X�wb:f��Z�d�Ӈ�𧐵)+��[�i��LR��Y�,���v>X�p�gw�aC�	�����;��eZV�*<�)���0�#-�8�m4�O���?3�2N$��ƞ&� �Ԁ<E�2)	��T'L�@߼UX�OTOz��vQ�`�'�|gi�[�1kj��������r��>������93T�;�2�W)�C3�a,��z�����bp�v~�L2��囧BauB\�B�K1��2�X�*��o�M|�̥�QP�MbgP�-2��q����?3�2N$�<q�OK�-�8�~{n���[UAB�yih=���'n��D2d��pA��)0c�y�hDi�2�^�,Hl����a�(�h.�f�c`,4ۙE��� �pV�l�B�����5Q%M}4�D�E�oͥ#�9)�A�)̪�PV�#�������J?C0�N6�q��[��a�a�Y�\��Wϡƒ^����%G��W+Rı,L�n�D��u�C�M%N0��jB-��"�I�E��mi�/8�N��鹹�+���]��OP���?��8c$�N(��4�&�i?j>��	9�U��jw�;�:�y�ʫ�߳Ga﫸�8㉈���E�-1IJ݅1�����幡��z#:���h�G^�r[eO![�������3O�������M,>�>���!0� a�¯�L�&2E^`��S�E�����U��G��Ӈ8(�N4g�4��8�8c$�N(��4��@O���בVFTR��ZIX��a��|
��0���s�<�ݻ������J�"'���}�d��f�	؟�����8'\վ��6M���P�*���i�y/�M6�93ؖ��c�m)50��TGZS��]��\Kq�LJ9�N���i�K�+�q��+�ں��5�f\aĥMa8�T��e䲷^|��|���Fp�H�8��x��z"�0Sۃ� ���'��):�$�[�|$��c��&�����7����\&C����rQ)*Q�"#�1��� s��K�4�y�m��)�a�7a��m�}i,���|�$���'L�p������aÓ��Sӆ���Ƙy�oDm�a���%F�:L�a�ik)�s���Ze�qo<��x጑�qG8�4$����##�sfM�׮��7"Jbx-�qd�*��j-錋M�(݊�Nț,�)�.Mdaۇ���)'�n[0M��ț.�[�� ��ء�#W���m�ᘬ> S�4�c����G-�ဢ��'�SNy�%6���y35Q�4�nK��Gb{8��!�NH�ɇ�>E��t�[�)Ir>�V󲡆a/B�I�L��2�m)���q1�u�*0K�DذV��}2��|;�1�8k��KZ��~"������J&X"'�^rei���4�Nf�c8�8c$d�Qǎ<i�
��I���#늢�f�[���o��)�2
&`� 
/l���g�l��>�p󑖞��u�N1ˉR&*�2��m)r*��������Xw
'SR�>0�N����#��'0�5��y����[n��`�a��0�)�L��=�ͺ��Q�g,8��=)�y�P�Ji�ϚZ��q�^y��qG8񧌌��Hm*���$������8��){����D�F�|D0Niߋ�HW�{=��ޑK�3�0ó=�;��L�ߛ6���D����t\r���[Iu&��ҭ����1�E\4�,y��:4(�ȝ��4��ÁD�vfZi�a�&�i,�c��K�p����ΙKDK0����qN���qo��8c$d�Qǎ<i����w�KoR�\[Lq������o���+:�l��,����<2���׺y�iH���[u�0���}�gF������x��g�-����O���Y�ٛ���+�y4��`bN��u���\̫츗���������e���tt'~���{9�ID~$��,fq�8јYe�,e��F"L$Cb�+ ��ږx�ǎ�gh��C0f�L��2�@�H�P�1��G"�1�cC��ic0C	220`�	$�(1�Cp�@�21�c8g�H�!��G�<^�ǌ<xјsKI��8њ3M���(ќ3N4g���Q�1�3`�c8��c�} �!�a AC>c�Id���1�5~|��nv`��ߟa��\�m]��wS�٦�E3$�c%�Z�M�$�O�f�l�2�JH�(c�Ee�V@x��T�;{΃�<3>��7X/N���Ö�\2v�����Tmb�w%+�f7C�F���Ol��Wm��L˕\`�HH��i�P�GfL{�F�\��(7�1Yd�)�Ԟ����c�2VfWl�.+�e�����{��z���������F����E�{6��^u��<W��okC�׌��}����C��%�VKHО��O�{�O�b<�!;�=P��M�u�d+q�cn�}�ܘu�n{�fu>��Z|�r�J�4y6����欲3�1X�ܣW�!��?��M�9�t�"������%ۘ�a�"�/�S�U��9�zχ�����4mY��>;�����{{�z����۝�V<oT�̍�!_vדh�ȰܒL������f�;�,�'�q�+�4QD�$�݋�Kچ�-�ڕ��V��*[�v�74֪0׈i�(+v3�I�X��p�Ѷ���Zǖ�Ik���k�5'���R�2�,���� tU%�Й{/[[4%�#D�&1[O���{�6ҍ�D�~��� (�.�CLj�r�)e�v�X��5��L�s��gz]\�Ѭ	���Ep�Yۺn��l�b0ݔ�[M�v#�ݜ��'�z}����{���������{���wsۯ�����{����{���^oww=��{a��Y�ǆq�Fp�H�8��x����1E3*&& ��e%������^�Ac.j�&�6]�5&��Ym��ٱl�wv�l��K+TL����s���j�BƬ��Ѐ�*��R���b�r�bo> Y��A�ܴ�4��Y�,�F�N��s3�aL:�B���|�bp��m�Җ�d�\bc�8�0�N�e���-��ci�Rjh�\
�
m*�����7�[�4������Ç�pM��c9&��uDO�?uK���WunV]q�K��b���g���"��&N����uh�:�����#�ŜY���ƌ጑�qG8��s������˿�&@�k�(��66��ùm����{�1LK�N�F�0��=L�2�4�"3�Ҫ[N%��G��Ė"~�QLV37�F����q�}�Bl�~�W�l������p\u���h�¥̆׌�%ۙ�C
g7m����s�{���=2�;�{<��yU���J��Z�)���䔭-=ꊒ����9�a�im���X�<h��'q�xS�b0��� ���SLUvB.a���Н�w1t�a��9%�1쭤�u�by.�-����5��D:4�ba�z�i����f�v���,�P��e6<�R����ҰXd6�Q;��κ��#�"w��������4q��,%�u*�cq&H���[�2ɦ�a��ƌь��qGx��>>�����U���N�0����D{�`"���0.���WR;��zܕȐ�륶3mv����QO�M:0�,�as��Qs�K��Xa��y�RR��ʉUa��JO�`�U���ڽD7D�'}�aق3�.<�~9�"`�Y�S��l�˭��V�q�d���,�Ǎ<#�̻!*�&澕L���"�l㬹Q5��f�Ki�;���8��]\�xV�*�p.@�YNS��4��4e.�%NĤe[c��Q���� �hmk8ݙ4)w
j�te>2f
�C�1��\���4�bs��fm.�ȣP�z��M0T�8pJXS)�S�b���QL2|'ByW�69��6����i�Nj7��a-�Ҧ��=����V<m��b��-��Zܳq6�j]V�م��:w��x|?�ߐ�Ð��+J(��JS�����g�<h�H�8��<x��AN�������z���/ީL�}'JYO�ԥ	��ڙ�98'�Ugp��M�a��>��E�Ì)ؖ\,�	�yyv*6�013m6�F�n%Do�gǁ�=�Op��Ax1@��k	�S;���DL�.�D���)�2O���v�X�},U+��o_=m�>i�^m��xь��qŚx�o�Ak�ΕV"e<0�N�0R��}�qs:��԰���&�Sh�\L[��&���$B+h�<�)Ar������X;�W�N��.v`5��þ�O'f' Ϗ�P�a䦥�%I�����O���6�R�n7G&���t&��,�'P����Ii�p�3��':Ӌ[�L3�K��*�:��L�fffbR��-9��栙v&g*KH����~�A;oOώҸZ�����)���wgUUGͥ:6�������xs���v&�Nh��g�r���ݜ���艻>�0��L���S��L�Kb\s�:�T����rw��Tͻu�0��&NOc���$�tx��Q��0����'Y��x�r�zeJ�"'$����R��8B-�,WTlM
Tб�LN嬉��L {�L���>F< �C����Q�g�R�vmS���Z7�"�	�+���ݙ�K�nc���T�m`�V�T��'~��#��;����4�+̶ݕs�n�nz0��<��DJh�'Ӳ��a2�T	H�_pi��;�����?/��E�DNC�~jV�C�W�����2i���sR��4�؞i���%�%+F��Īa��vy*J���l󝄳����oI�&���&���-p�p�ju�6���S.�&_3�
_���Y�0g�3ƞ4c$d�qf�<i��P�p�IK>���SL18����������`�	K��t����ʭL�IK]T-�Řc�� �M�Fd=�QM�i�M�y��.���	��{��*<Բ�;��F�;+�!���
�Q��}����FG��~�G�m��A��'�>C�TZ�]�����F��L�Z|Nc�ᶶҞi��8�ќh�,��2�Q#&!�1����\�0�3qiZ�Z��p�^q��my;pf@��&H�1�3�qD��!����1���c4c4eaǏ))y)x��0�T��ǁ�����1c�p�"0e���G�<i��x��8g�dќh��8��I�8gh�4��1�cG�Fh��0��B1e�db1d�2���&�#���D���-ݝ�ﯝ>be� )�n?6��}����&'���TP�o�>ຶ��חb����goEɊ���`�gk�'F��Y�,��+lZs��X��7�>n�6�ǅ�c�Ow���x����LHF�>?E8,�OV�r�:+|���XZ$&Ro��8E���&�Z�1i�{��`��eZ����nd��*>��=��-F�ܐ�u7��}}}���ov�μO=��=��^�}�wM�I�E�UM��d-�0����~�z��{���N��p���uoi\��L}6�4`{sr&���wu6}���Fq��tG:/�s��5�}#����G�~���^�=U�ϗ�~���G[{K%f*-\�q�$�A�fչśY{�U��=�{j}�:�������'.����VF�����=�����n�����[{����{����owws��{���~{���۽-���V����qn-�a�Zqkqj��fff%-G�ٚ�ɟE%N����V�҉��>�!��<��0�.\y���UTJ�����qĻ	g�[�!�z�[�V�B�TM��{�G��a��S�|�~��V��=��%0OЦ��6z&��q9N~�lM��!�Ʌ;N
�D\<�RD}���#������V�p���<i�c0��O��qŜx�����ww�x�� ���9�0�JT�={�ͥ�7ى�by��0�n-K��&Jkk�&�ST嵳���(�gs�����z�"e�Ԟ�Â'��{m�É�a,���L�>�7i�UUm�R�Ŵ�4'^��*w��nf4�L;)�M���B{3,ña��m�y�m��<2FI�q�ƞ#�&#~�E)� v���{�Xp���^���Q��$T¥TRZ��բ�d���&��e�ѥn��[l4+�Ь��nt��Y�K�O� �w������V%%�钵�!���P~�{<
&�SM2l;>99���a��ol]�rQC �	�o�(��i�;��(���p�0�%��S���X�be���aC��k�&Cߍ>�	��U0f�14r��2g�����I�a��P��\�T�J��6�-��6��mkqo0��ӫ[��TĢ���C-�O���x�d�,ѓ�I�G��m�.'OIs|UX���Q�I���a:95T�M�N��[V�X@)���B�'7�sq��q��Jመa���Î��5ͨ+ϸ�Q��z��,���W8�*�8�sڢ�z~㐑�xJ`����l���4�8�֞�L�1�'�����yŭ���a�ƞ#$�8��O
Ɍ�S"O�UX���u4�<?`�O��}�e�m,C{&b<�����q+�|�(�b��me>;kA	+���M�53nff�9��ɥ0�-���3�}ϫ(�̣�o�3�\���Ϛ�ܥ,D��>�'�u�&JV�*�"-%�1�����,��1�a��#$�8��OTyJ;��ΕV"u�g!�"�k�J�n����KLff|�)O�<�,����u22�uT&�iL2�f~�O��H�a�t'�G�ۏ73�R��j<�!�R�S��j#�R]Z�����>���K���9�G�/�'��(��N�Ե,S�V�8��KP6�0��4�p�Ǎ4���4����q�//�����Y���,R�l%!�d��,��.Q�ˋ�X�2�S�8Cb�K�/<��i�)b��Q�2�����C��,��R<�P�Y����73�fZ���3DkVRZ�6Ȯ����﯐ ��ӫ|�pHVhl����Sr�	�!�W���t>U-L�Ym^`.���S��a�d�['~E(�K�]��f�i�f;ɝ��F��[�3�� (���%�M��D�݉����!��C ��Q��n�Sh����f�^3r�L��v�;>w�bp:����'��K��?��wᶟ���I,e�Ï~Ɵ�xd����������YSt�bc�330�,;����s�>���3��V�8}�_pK̽�zn��X��E96��uLh��e'!��a΅�ڟ,8�gw)����g�zg�ai�ԧ��U��l��RA��x�� �_��~�p��Jw>:��t���z��L4����6���e��
X�3Oxgx�H�8��<x����e��VE�l�EUZ��B("�
6�X�f$q-��ڊ4[)c�S"-�
���K�y(,����:`�Дq�ң�[��Ve��)1;�IC�!}�Z�=g9�K�[9�p��c�Nxop���0����5g��B�YOg%��G����x}n�GR���4��b�
��B�v}%�����(�I0�����-m�l<î�����T��R_iD��#ice�B��iImEr�؈[Rp' R@- 9YR���G�-�,j$�92�����p�~��r)�/���v�����Se��ٚ�L��Gt�R���9�|a��}��O#:*�uU��5�0�^Qa�/F�(y׽-�|�[O!��NF����2�����b���ñ���~�3'��Y���c��N;��:��V����V�o~SJY^�YZ��ѳf�Ç��&������{�~:�[�z?r�<8v��ܘIap�/�A��2$�FG8J�@b�t���D�mE�,D"�"5�dX�d["�";�ۂ�F�Dh�ș"4Y,�!d[E�m,���m�b"D�"F�,�B�,��H�d(��,E��дD-�"�4�#Y�h�-�Z""E�!�2"&DB�-,���",E�DZ4E�M�"�"Ȉ�5�b&�h�,DE�#Z"-��[DE�!E��-�h�&�H��ii�#I���l��im!2�4��KiĚX�&M,K4��KibM-�L����%�%��[HGn2D�&��%��H�e�bD��Kid��d�d��%�%�K&M-&�I,��%��Id��D�D�I�-��K$��Y$�I,�,�ѭ"Id�Im5�$�,�[E��#ZD��,�Y�&�$�KI���D��K$�Kim,L�"ZD��,H��m2%��m$���$i,�,�$�����$K$KI���Kim2K$K$I-���m2%��d��ĉ"Y"ZD�IbDki%�K$�d�d��mƒIm$�m"Ibd��%��D�I-!-&��I��ii�KH��K��&M-&�I�Ki$KL�%�K�F��HKim&���M-�Y&��Kd��M,�4��Ki4�Ki�D�d���M!&�%��ۧ9�id�X���%�,H��%��,��HL����Ki	d���&M-�K%�m"Y&�L�Y"X�,�$I,�b[H�H��KH�L�id[I&��il�m,��	f�HKil��Y!-��B[Kd���L�Kib[KK�m&�Sn1,�Kim&�I��m2i6��ib[Eѩ�q�%�ș�1&H�����dn q�4C-6�F�Y6�6Y4�$�i� �YH�Ѵ�Z!�mh�@�$ؓl��gi2��L&$�L�:��1�Qd-,��DF���!h����dH�DE��מ9""�$X�E�8���pH�m"�H�$r�"m-��m9���m�mЖq3����-�"m�0�h�mȱ-�D,�g��DE�H���.x9�;D�""ȑ��E�L�""Ȉ�",��"#�8�dH���"�$Y9C�YE�"Ț,��h�E�4Z$Y,��kD�b&�mDF�E�D[D�""Ț,F�D�"h�&E�DY"�[DE�"-�E�#X�D�""�$H�E��"Ȑ�H�$Y�d$YD�D�dY	-"Ȉ����dM"h�&��X��dDMD���g��-�"Ȉ�"-��X��h�,�!E�4,D�dH�-"E�"hYD�F��",��dD[D�"!E�4,��F�"�$[D�DE��,��dDY$Y5�,BE�"�5�"�dHY,���"��-�dDY,�"�E�DY� �(���h�2ȑB!dH�C��6�X �H�2 [DE��-!dH[D�Ȉ�h��$Z"&AdH�DY�h�DB�hD�!hք�Ȉ��m""���f�h�b-�"�MѬDȴD[D�h�"-�[D�h�d[D�m�f8�",�""�$X�E���"ȶ��"h����D�dH��h��"!E�[DE�m�#[E�����ȶE�D[F�E�����[D"��E�DX�h�&D�d��"Ț,�����D�"dDY,�#ME�m,���$Z$YE�E�"ѤY-�"Ȉ�h�h�&D�dMD�di�DE�H�,�Ȉ�H�-D�mDE����h��"ȶ�"ȑdM�dMhH�H֎���dH�H���dDY-D�F[E��h��H�$kh�"�Z$Z$Yȑh��"-��Y�di��D�h��"5�"ȑh��-ȑh�,���A"Ȉ�-�2,��[D�mE��4[E���L�l�dX��l�6x��o��[���ѫӺ�λ�q��u���=��mhljV36�Kn�ގ3�,�_��������z��������g�Ǳ���<�����?���gD�����C��ۣG;����.���=]���{�_��y8?ONz���7����Æ�;����o��vzONpޯw�M�Q��͛6o�g���q����/�g��m�;s3��xm��c6l��8�"�n���3|�?���|�{�o��8l�o�3�7'�o���_F�}i��$��+���l٣ٛ�__�>TI���;m�o�^�}�������nZ2�u�&w��~q�g�����0�pn>z�w㫴{��g��y}�o;wgIݮm-�׶��^���t�\ i�src�m�6��@ms��1���h,�:[lB5Ɗ��R�D�>S��`����|_Ws������}o&�ޖ��Z�`�Q��$l(��Q#���3mF�ۈ��6\�߁�����i�Yշ~��|��~�ȷ˻v|緎�o'l:8p���}��ط��~w7]��d,ٳf�>��g#տ.��u�;o�ۻ���vC������,�:�����?�|Σ�=ǣ?�:���s;��e�������}g��ُ�z����s��>3f����m���gʹOW�z\�o{��x�<[�!�OGfq�������l�u}8͛7�=���-���/Wߦ|n<��9;���[�'����NE�!�9wl}���c`�w\�{Yj^-ʮ7��i���,lm��������6�f����ټ��3���g᷸�u��gv;u,��	0f!������!�E����߶͛7M��_���|=�n��f͛�s��ٿJm���=�6���Ǵ�����#������=G93�g��g�����n�{O���?�o�F�}y�O������7�՛�:6lާzY���6�W��v�f͛�������y�������z��������I����'{<�ÿ)�f�I=�O_�w;�[�ӣ��:5�����G?N:dϛ�x��|������xw3�к�_C9n]����x���͛4�r�m�m��q�.,�g��7�����:����ۼ�G����Ў�����&T��#H��D����ݝ��^�󰙘7���nw��6vw�3����n��u���3�������'u|�zݜ����!�?��~�w͕�ל�#Fއ�����.�p�!��Ю