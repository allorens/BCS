BZh91AY&SYcӭ��{߀@qg���#� ����bJo�              �T�j�omTQ֢T1d�M��	��J��
�jlʊ���B��֔P��C3(ٔU-2�
"��4�()Kf̐$Umk�i@�J;aRH�J m�@�֡B����J��K@Ҥ���UD���jH��$QP�� @U(����h' 0QU.��*"�L n�@Q%d�r�*��v͘(������Y`�	TJJI*)�UJ9�s$I
Ѐ>yJR �л���"���{�W�=�]�vF�R���4��Lo^z��7Oxi�{�W:)s:�1�T]��@�wb�vӭ�v��zUEH��4�%T���II s���T�R��^��*[jT�����O@5vn����l�M�t�ޝ�T�^:��Vƨz5�oG�F��U/8�m+[�vTwN����SܝﯝTzeO�=�޵	J �E�JH*KW�%$� o'/���
��[���P�nמ��M7��p�k4w3x�z�J��<<�J�킓�y��k�T����z4j/se�x:�zew/=��u�]��(HT����C�ϒ���9����UNt�=�5Y��^�U�5Xw�t=RTϯ���AJ�N�]�3�V�
^����;iU��s�{c�[j�<���)J���Ҕ�=m�j�WE�%"P�H���R� 7��2�
�o��T�J��ס��T����QU;��׺�U-��Ow��RJ�8:��9��(*�Tw#���Uz��2��^��S��4`�ΒUP�_|�) �ER��{�҅{���+.�P*�5�N��U*s�P
�����[����րѼw� ���p: �{[�@ �)K���J�d�\@ru�t �F 7`wm��t��r ������ ��{� ���r;׀ �8:tJ�J��kTJ�TG�)% ��@}0@ �ܛ�  9�{��@�����{� 3�kW 
;�`N�S`: �Kr�:��P��P
HJ1G�)T����  3��� �n�hR�w3o^P�yX ������-���^���� =��CL)%4j�Z*$�>�JJ |�@3}p� cv��:����@�� ;��@P{�/o vE {`: n�8dh��     �  �P  ��2R���zP��4�0��1%*�       5<�%U =M     jxBi%J� h     ��JRF*�� � @� !!�I(��{��Ҟ�M���4��6�H������_��~��~���8�����L�5m�o����Ӯ�ʺ9��/�|� j* �T��
�� U���}���3��?��O��W�>�?� *���I$��A ~��̂Q: (�����?Ӆ1~�?���`����.0q��L`���ؘ��0q��b�8��8Ŧ&11��bc���&0#b����&1q��`�)��b[���$f0q��`c��1q��bc���%38Ķ11��L`�8��201��L`�8��11��L`�8�c�`�8��&0q��)��L`�8��11��`��11��L`�8��0q��bc#8��.0q�c���&1)����1��L`�8��-��S8��&0q��`c8��.0q��Lb�8��.6���c0q��bc�`��8��11��Lbc8��4���0q��L`�8����0q��Lbc���[���11��b�[���11��Lb�8��f0q��`����&1c�&0q��\b�1�c�$b����11��`���0q��`����.11��1����.0L`c8��c����.0q��b���0�.11��L`�8��.01�n44��&11��\`���1��`�1����.01��\`�8��.1�8Ŧ1q��`�8��&20q��\`����&11���1q�l`����.11��\c�8��.0q��`��8��0q�c����c �0q��b����38Ķ11��Lb� �0q���`c���01�l�0q��b�8��&01�`c���11��Lbc���8�1�c���&0q��`c8��c����&11��Lbc��38��.1�0q��`���`S��01��L`�0i�11�lb�8��11��La��.1q��\bc���.0q�1�bc8��&0`��.11�����0q��X�A���1��b����c��q��\`�����im�l8���\`S�1m��C�0q�c �S �1`���h�1�c �.0b��6��L1`��F�1q�c �.0m�0
`� �.0q�c �.1-�1i����1�c �0-�����1��\bc1b��1q��`��0q���!L8��.3��`����1mƖ�8���\`�0�.0q��0q�����1q�c8��ŌC��1��\b���`��.0`��1������\`�c0q�c0bc�b����.211��b[b�&0b��c �!�\`�HA��C&0`ƀ�.1b�1�c��S��[`�Pq�0 1��0Y!\`��q�.0�
8� ���G�`��q���Eq�!�Tb cb�q��0Rث�i�.1� 8�G��\b��` c\bS b��m�.0� ���`��`�� #1�.01��0� 8�G�� \`�Qq�%�bLDq�0�*��G�� � 8� �\b%�G �\`��q�&0E�
��G��\b��0�
��S�b�Dq��1T�*��S�`#�Dm����cb�q�0�*��*cb�
�[`�c
� � ��G�c�c�8��0q��`�1q�N48��11��\bc8ķZbc����)�Lbc#8��0q��`����&0�$`�8��.0q��b������.0q��\`��Ŷc �1q�c��C0q���1q�c �.0b�`��1q�c�,q�1�c �.0b�0�!�C1q�c �.0b�c0`�1�c��#��\`��.0b�1��11��`�8��1q�0#���.11����1��i��`����0q���`�8��0q�o�@�$����9���ίg0��N����6%!4�D�&P�Z���䲅�^z��["8G�n�4�[d�ݗL�;b�j���)��S��Z�%Q��xu|�i0�L��Q���  (��E��,^�vE�����1s8��a���DlِZ��W���nS��۠qٷ�Q�n�Y1U��eږ�]Yx�`ƝZzC��
߳�Vs5��sz�S[�N/������i�4���c�:�T���c[[�(nC���iz8��ᡢ�"�R�N�pp��5�`�(L���<��v�;�۹��4��0��z�oIҮI}±���I�1G�Z1+Ur4����m�E��������x����q�e�/�)"�FF��eLV��*}�"t�!�}�R�JQk@݆C,i�H�F{l�*���u�J�n�]�o�/���
�%�y�Ѭ�mb�^Cw��G��=�;�ug�<��=)M�ۃ֭�wn��ˌ�۬V�b׎%2���nJ	>��ηc{F[Xf�eH4렎V	�]� ��0��rn�Y�cu<�̻[�7S�2N�5C/a��=�V�`Ú�Orf�pCY�`�eZ�Ъ/i��&�^�t�8el�*��b T���#DҀK5�{�͂Z{�^P�Z1i�B�7ͧ t�y���븐h^�o�$�ʞ8K��cʀ�#��f̓^H'��~������'U�e/�xl�O^�y��AAC]6!6�"2�7�f�0��b���D�')���a�O�I`�L��;�DЖ�o��ڬ������:�X��O���l�v<��!�I�x���Z�0U���mǮ]�Cp�f�2n�N��d��R2�yV�8��U�9k�y��X���r�����f�Y$F��e�W2�x��w��"+rWm]F��Ta�c�����Y��:Z��P]X��$�5��{+Rz�UO%71��N��H�ȗiI�ƭcWn�Gn��[�dU�e"+A��x�5P3��%�����*=λ�y�f�S�A�^�1�i��%
�i��R܋"�1�Dܙ�����gF����L)�.8P֚#u�z!�b�3�+U2Z�ó�%Ҏe�'������ҥ�떃7*�~�a-Ę�k	���ެf�8+���u���͢b��b�y�	��eNa�n�T�+,^�H�c&mMO!ׯ0$�we�Ш�F拁n��J��znm�G�z�c�{-㥵���*�d��ŶR�<gV�!�W��5�-V��������/66�n�����L�.XV��%ҹ)f�U��t���`S�lꧦ�/�-�*�(a�㪁�L�֮�:Um��M6�c�Ahj*�݃9���s�"
ݫN���(P��S�id�מ�L�E��.տ-�I>�'�҇."ŰK�����!�Լm��x�ˬqhl�/#�l�	�,�4J}',�T��u���C�SW�!{���V
)�S�&��nɲb;t�U�����{{���`Di����$���Q�#̕E��9[�+��bP��@����L����B��2'�;��ۖ�.�6���Zr�bj�7�q�㔋2���#z
3�AyY;]�W�>�*��$̫Ռ��Ȕ��D2���*2+1U��c��1�`TN���_4�����d긶��&�e�����1[vN��˖�s*]��y.����8:C�e��r�̰�h��U��IR�:�7L.Zb��R�=�c'�1Қ�g����ԝ1OV�j���s��N�A�ww��Yscx¡CV��pt[�e�	�c;��Ԥ��:��M%
f�yh���R�Zn���-��`�g�Žs ܎�P��e8�t��Y@ɦ)d�����)z��1^y�56��B��2b�.�^��̧tm��Cv%;uX��U�u�XxuI�y��YY���E��lE��Cj�m����.��$��)hȋ:b�h��r�]��ڐ��;,��(��Zt��0�e"��+�H��#&C���ln���IZ��R��.�W���X��;l��X���]�us�ˉ�H�Ne�x��D�H
ˢ���H,�����K�������*խeh���c��[�M�9LQ��Ksc<x��R��Kf�'��eTq[�L
���D4���H�o׃6�Z���r�<u�����Y��q���6K��/�7&-�ރ
Ӭ�e��-Oq����9�h
���Ǫ��#%��:��)��& ��Xѵ�w�e�P�FX�ٔ�n��l�F�\��52m�8��0�+iw0;`��VC��)�G	�WO)��K.�I���ܔ�9.��
��J��6++6�R ҩ<�w���M�a�-V9h�0�"��-�x�a[ɖ�����%^0p�M[w�I�,�r�|�T��b5W�	�|l��=�x6�ҦdPj�V�!]�������J��1�r��u
ɷ���h�{�Sd�cm\b䉫`R`ԕ�4C*�wD�xm�V�v�en�-ת��Cu�8n��4ݦ�!n��#v#Db�0(ü4�2;�#*�S��a(���B�FV���[W-�P6&R�ʒ�'b���(hi�ŷJv-fj�[���*"ɧ�>�ݲNۼEûj��T��̖�E76�SK/k�3*��ج��T�c���Իj��D�N�bn}�Q[V�l1f<܎�@Un��w0�ŕZ���r�^me�pc��7�*TRգN�J:�ze�{�)� Uj�no���l6��!���ǀ�6��(��1^� Ā��x����x�H=��]���M�V���m������-��#��k��u1��;���C�P]�+IbV��:N���E(d�EPRy�o7NI�Ma�7�3sh�h;��Xۗ�ChL��V:̢}xU6�Tq�A<[ZN��:�6�rR:�(ƭ��M]�U#��o
1�K6K�ʦ��9��v��hfM1ˤ����lN �QӵW�ի�ݗ@Z-'�@jKoZE����p@B_2�Ƿ����2X�"7B��m���ٻ�����Zą]�mf�L�J7Qڹ��9y{tv��nVF*�|�9:�B�x-�[|�����F�w6�����f,�M��86�e�t`�U�갚כ���r�1�ܩ6ܫ��2�LÒ�c�7y0f���^���ɲзb34%�C�)��T�ac,\-����]�����f�`6v�:�j��n�R"�*E�Z�6�XÄ]eEJ�A��B��:�J$Ph\i��N�df;�nҏc!�m��h[�����n��k �˹�	x��������rn{#mF���Y=���nl�O�-�Y��� [V��bä5ޒ�̑��&LZ�Jw��kt4�uX�MJ��o#2�\mWoP�卛(�,Ȯ���E�雩[�R��i]ɉ�m��{��YfV톶Rz��!�&hkS�kE��(2R����5.�*hm��賺j�ٍ#�<d�e'�,�7	'�k,�h���o�O��y6��b�Q�����%��E9��U��kl�3*��B�(ދ�
�#ꪛ�Q��������04T��-�s.l�A��j:��'�lk��n��,T��b3����zt���Yp�*�z���ǇT�UT�d�f&���X��ӫI��	�2�T`��u^�g	�U��t2�\b]7v���{&F�F��(�ǹfGmڹ��Ov��8��6�Ѵ��6 -^(��%c��n���D*�\�z��h�a��躭4:+CX���)9EX��d*8^�W[�<�ǥ�e�(�^�T�����;m歠��A��]ᡥ\T�2AJ�<6zb�6#�r�{n���W�+�[/ m�m	�*B ����oq�KuU;��U��w5N��6��T����ۣ����-=jm�-���H��:���S{2�P$��\����b��KJ�J��=�6cr�p�9+r}�
J�fB$CU�nX�^���Uj�aR�+�r�u\xh�[���"%ݪ�06i�����u��bM�W���4�^�44Jv�btI-�2n��S.�е�Ch��׳����-v��FfT��� �\B�VS�*�,ŗ���W��;�^C$��r(��uuv�1����jict�ͷ=�$�l��ׅ�ae�Z���0��fi?n��<��a��,��G!����oi:��ͳ��Wq�B�ѽ�5��٣�H4r�"��
��p���U	sFb�2�Jܳ����)����	A̅�JF���J�#&�9M`���
��F��rT����#t���#Ƣ�����hZ��㶆��K����� o]��4R�5�A����x�<-���E-.��tKH��*hP�3j �,1eQ��]օ��w�RJ�j
�`�^�	�kT+$d&�̱�2���&�a��HuK�d���V���p`j���E8&0Y��#07}|�����2]�l�xX�l�
�t�%���me����T�%�V�Ȏb�m��j�̘2��f���j�/[��pXq��Z�Oy7��'��;��;N�Q���f��[��
;c�PxJ"X~��z�U͹��^fF=7��y]�1ڹ�Wך���,��	k2�%b��us̊*Ů�lׅ��f�S?7[Z��A(���lB++x���ȩNct�;��Զbq)RM.��<W��N�ے�1���y5�7a�:^�0nV�R�N������å�G�U�0i���ϛ�F�8kBWO.��/��Mb�f�\��TS%�x�\��L��Gr���`i	�w2!4ɘ�̴!��uʙ�Pa�cAtQqnJ��,������R�^����Ŕ���cWQA�����ǅe�E��{`��@�X�6�fc�웶����RU:J0�e`�c`��wND2��n�e^����7&G���3��f���6�K�K����m$-"j����n�M&�K�gz�ع.���5{qFZe���$LP�%����E�Xywۍ�ÐZ#���s��4���<�A�Ⰳ��mc�Il��	+�i,k_׮��t�:A(��V���A[}�}���wbmئ�w�ǒd�5����Z�*���Ԇ୛q]Q�4iW]�&'>kp���7��SE�.��)l��jMN#W4�b���Z�r�2��3A�^��P\�#��w�,��e��`�/-��
Q1�$��6��+q\M�Y�k���nG�֮[V��-��)AުR'eޝ�
����ڃn��e��ՌQk����`��xE���Lݍ�[R����.�������#X�3%��U�<A ���NTUKJ�<�f����YU2��u�i�R��(5�@3J0K�p���f�f�N�Q�����h˘b��!����B,B�(pշ�T[,�Z ����P�����P�V=���0�܎V�a���`�2]2(�"�fȸ��w�	r����9d�V���Y�фATh� >!�TYF����#�� �%��Pg4U;;T�LgvuԴu��'C��fk2���+#����7@Z=�����P'��
��Z��ET��j��ѵ֍δ\J���u.w�����J�5��$��iSV�m8�Uڬu��jv�lZ D�
�՞�a��rض�U�]N �^]�m"e��Ar�:�֯Uu#�VH�$#�^S�)n2j�VC˜�:��F-�uV���<�Z�6
t��k-�PjY�)T�J�@�EE�`��N���	���1P5���;qn���$!��˴-�F�k�Ӫ�aq��<i�@�[j��cn��R�� �f�SmmY�>$������@�R�Z��A�Ȅ+Vj�-J_c����QTn�3{kb�T���0M��!�3���B�ŏ)'kRTF����-HZi2cq)F��3$*��LH�J(�EX�M��A�$�Ś�ڪ\��2ɕ��}�֎!���K^{u6D�)�Ϩ\�H��*#N'����4��ЭB�Y�H�k�D�7^u)b@�KR�+J�G�̱��*�e�x�8���B�>�Ē�B�ۦ��g"�Q�Smj��J��A4�=7���B�;��."⤨��5��"��cȁ���#(F���*�`�������B��^�z_(m�)��m�N*S`�H����VՈI�)ẗ��j�5��^M��c	E<[�M2-sO��ݪ��`�Ka�M<p�(�o,�}��Wid��V�|$�I�Y&�Z�� ���A+�A�p!:q��je�hi���{��K7V�#!�^cl�C@ZR�
)��|��h\J���+��b1w[wVbM����8��[�-T"�v�jE�I��pѽ����w
�k�1[屝5k��Cy̢��hiGVHd��6�+�W�I��0�K�)*L�1��i��vu�j�C׮�"!�2�PB�Zb��Qδܜ�Ԗ������4(�L�b>�����5P���v�r�䳨�(�$�B��#�����iQ��
��L���os�D�Yj(ϵ�L���dB���c�.��R�&�泻+&�{���E �&���%՝U�l(
4�A&^GNT�k�Ju(Ӌ��%$��=&�4��B�[Y�zN�4�,Ո�+��0�R4�Ë!- ��,�Ut�ܸΑZT�������L�"�R�%�iD��M`��CK̶knWH�����	%d�{O��2����r��,� �&K�tڻ+�ҳi�8᏶ɩ�/ț�φ�BkK�x�����q�! ��&�b�l*�ٝ�bH�X�K{���9IL�i��W�n� �4�v(�"7s��ҵdp���i����Rq�c�L{���� �b�Z
�c�ah,PF�%v��#����9.�t�d_E����y$ȭ��-2ZJ�X,��nb�aRjlP$g;.t�����ȭ�h
��G���EERȡ�g��Z�tN�@��^6�K�۾����������~�����������a^g߄�I$�I$�I$�t��,�w�I�X�I'H$�I$�I��$��M�g�A�Ѝ�l�s�t�&�.�q�����
��^�}/z�Wy� �W�L�_!s��e�:탕����ٞ�6(N��9���u�x8���U���Q7{̉�w�Ү��+�����Rm����72���͕���tbj��:�=v�
��U���q��0�������k�y˱����s��	]�X�2Q�8�8�mk�6�x�=�Ǔ�;�U����5VM+�ì�)��P��k�\�0�oJ��ζچ)]O(�� ��9DVX�B�P��\+5��Gv���:�eӜ83�ow�^^^���S��qS-N�%i�Y���^����jhY�s�_-�r��N�{��n�����c��7.��\k�Wɋ��u�>�Ou�FkC��{�j^-:�K��
=e��q�:�e9��c��A���־�]/�`X���W̋JL����S6Ŏ��6ÚC��|&̣���t�h����ʾr��J���[}�/mV�\L��@�EFu[��T�f�}�)������F$��]�i-y&@і)�����Ӻ��"b�:�r�W���Z��m$g�W;�,��;�7ZB���V接b�؀��Y����iRc�I�>��gY���p)v���M2�����  Sx�_My�eS���|�e�����}�ֈ��R���q���0M�DK��×��f�I�T����`�5��W�N�Iᓞ��g���Լ}Z���g�c(\���P=����9U�� b��������0P/v��0-y��`���f��.Y��[e���ȆP�;H|׀<o]e_�^��0���@(��.�{V�]��C�W�g[��YaZ���M�v{�d��T��!��;�n�T)6����0(goױ�#��+4*+"ڭ�ab��u�}w6䕭E9j��93��i�Ykvs��;I��MC�z]�7�r\��u Ŏ��Mve�S��upo*�{��]`����{z�.�*�7lm��o�pV7!��HV�weP���{�������m�1�xq�T�:w��'�Օ��i��]��T!2��Q5����h���:�f�6+0P,���U�iJ�l�;Q)fQ��F]5$ٌ�1(u棇�J�۷��|i����;G"�ʴ���.	Z3�r���X%���ۧV��TPu��g�w%O;��n�<Vc��2u^����e��Y�J�#6�V���5%#\%���7�sǦ�(���hJR��ubţ'l���J3yn`Sˋ��vKŵ&-N��yn,����0�����ζa����7ML�����+�2�3G]�D���F��1����l������3";Rn�Jы���g��̷��R�	�A��������+\1����x;����t�*˸;
���Է��e��DG�.�yZn��v.6�s�rod���fR��:��fL���gi0�b�*I�)vs���\��ou��a�ņ�
�3\ݏ�=L����ƯOa影�۬�i�<���T�p��'\�N��i�#Zv/I���P�-�sڹrݮ��-qWF^u�܃���g`�Ǚw�U�v(kv���޸3uA\�s-�j����]Ү3��-�Y��9�X�>���\��K��u+w�-�]�Y72A#��l���[�^���}�ݪ�u��%�6�7wә��`�͡���52D/��Ȝ��OM��7��-w9h����W�9u�T�]K2f�Ư_q�(�&�b�s��\�e�ə���Dz�xi���4Ao=^���+�'�d���<oF�f�9�Z�1��gC�Z���,�x�4�dٰ<��Z�ֽ��f]5bj��I�HN;=�Ul�x �V^-�Ȝ��@ڙ1�B����M��V	�z� l+J��6Vj�1�;Fr��zMc��	����.L��^<օ��ཤ_��AF���bꀞ�׻z{���D���t�ȫ�]��r�m*N�F�=����mZ�¶�	6t�.��^���iL>�l`��[��b�nT�Z�u���]i�!%��{�����u��	}{O�a�k�wM�Ә���G+YZd��s��-s��ث�-پ����mgv�-y��%=�q`��o�Z��nˢ�Yt����Zz��cI�8�SS�s����H��"�{Om�]���{C���U�S�Xd"���nJ��S���}�TQg4�r�ee�E
Ê�j�[뮷�Q�����j���,�(^͡9V��N���v�Z��m�%d�oze�Q�n���,���]�Z�N�[�6̶��Vt��b�қ��i�ed�Tn�f*�9��n51�С�\�
�V�]�
���w�>S�M^��;�O��i����傣�R����2	�C�w۶n�nK#6l�2s�O�݌������+Q��D�v��N��}u.h�U��q�d��!�vv�5ڝg�fBf��<mх�g���p�����S�7��cy^;�smӛ��=�gsJJLl��=�cp���ϐ���uxr��Ds���fn��$�uU՞�ܴ%vx��k�_Mh���q����3�I�u�\mf��_.�.�O�a���B�=�����#z��⤡����_lubw����lS��Hh}�;�\3bf�w:o�����0�J��S⦾�>]�yNvDe�3��T��)�l��;(ǽ%s���.��u��x)p4 ����}��u]ay��َ�� q; �,�[j�"�|���C|�����c�c��ࣛ���O�u�Sw2s�	/�潘���'��Z��C��y�;����J��.F�XrƊ����A�j͗J�=ע�t������d��!�n,��P�ڈX����Y��"��t�Jr�4�w�tAoz���+B��Ϛ���w�Y�ԁhY��x2>�2���{Pk��E�=PYW��>��n1G�
�0�Y�vZ��cνo���w��w�՛^����z��=�����f��aVW9�ƫ��_=!���1hm̳bi�]���YI�OLS.�N	�X�u��N���n�d+ʵ�%g���&/j��F��oz^�=;.��uoe�弶ň��m�զ:�
I�s��|f�bڼ�Aܥ�"��|�2�Q/�1�(�,�뱈9OU�z��u5��7OWBc�S�-1np����*��c����S�;���哢�ݼ���᧾�j騆��:B37�U��r���*Ng��8���u<㘜��Gx��:�e�iC(J�k1pN�`��Sx.�5z��(AE}��Ȥ��J뫺�n�=���c�>4�C�����N묠��6�N�g��`�b�p��h���2��0��SK����U�-��o�/���l}(��-Ym�Oh��8��p����BΓZ4��Go�S�7:���ͅS6�gH�NvYM_u.�'�ݑ��Z4���0��,��a�r��ca�|�C���G���7��vf`�T��N�i��h�%��z÷(mȌ��q�9U�Ìf������(u�Џ9�jh�:v�7��%*gi�n5�5��(]t��ѯnӨ��dE7�u�n��a�ą��$�����	TW;,7��t��>�;_v�-f6/�T�gmAsx�J��vR�5Y���:d�H͏Q��f���^��/�u���$˪�һ��:�成ޚ�I�_҄M��ħ�^qޚC����ۜ����vwFV^O�3�J��Ꮚbu�j���c�kBbݽ�d�D��V���_k� o0ER��]�@�J���d�Վ����vCzk{�M�F�;d�����hn!��Ad��!�>#7�ѡ������wcX��{
E�	�L���(AwL^͸�#�W]�����P�c�	����|{A�����'�0(^����9��l8��c�Xm���4]�v1Ԟ���+��8n�f-#t���m1�נ�L؝\KK�0��z*�f�Y�9}�{Jdײ��F���Ω�wU���r�S`{H�8fA[��f�xWG[9$�n���Ę�O�l�UяdTُ���X/��sk� ���1�}N��ޤ�*D-��W;���ƱI�lu���.Z��'��meHb�P)�槅k{/D���z�Ĩ��da�.�eEX�`���9%v�$B��'��i�@�ԓ�R��0�Bs�Nw�N�k�I]`��jN�³pMv�Y�6��Q��ʬR�m�*�P��HD�*JW������X�:Xާ�v�_Au��-�Δ�E,!c�mf�Xӽ�'_*y��p����IڀW��Mv�'%5ʛ݊��TO�UeZ�ka�\O[�l���P�B��00��U���G!�G�+�97��m�m-OD:�u�T��â�ܬ2ܡ�3��>Ȅ���U�%r�_w$ԩZ��w�P;X�Z�l�����x�Z3��z;d�}�\��GM�z�7��Fk4���l��s{v�S:�L�����/.����w��3�F�3s8���!E�V�����2n��|/4��!�I����}u��3v��x�*�1ڏM�D��*�4m�w�*R�o}�-�:~�A���d��n!���w�X��l{��Q��n���K�z�K!��vR�/E[�d��+jI*�wW) ���bMu3՗&�_6]��O1,x��v*È3W�7�S�O�M�WG�\�4(�v�)��1����OU�L]*q��
X�Mzb�����W+)��*��#�V��\���oIj���z!ְo<7�q�FgǠu��6�/�^k;�s�G��8������2�}\��f��G!���oOZ��[��![�:�IAAl�P��<W�@k��l$k�(����ʛ$V���G{o�m��eO=����p�{�9�1�!_.}�ի4/a}cB�g.���`�)���=J�\��y�I��*t�3�����Y�Q��|�3��z�Y�ֳ��:�g�]��%pY[�yq}/�t�b���̴x���c�Q;�2j�9������мx���g�Vy���Z�nr:j�� ��laU鷶�f��Pth�N�Ϯ�mү�@D�|y������^�,�`賞ˆ[�Y��3mvp9I�����dݫU%��dW�t�Q@������k�%f�+#5��x9����Ț����$�u1Ɏ���sMﳕ.SvԽ�H]�i�Z���P#RKT�kS�-SD��Ԯ=h��]���;�^3��\s9�,;o����Ա������k�J��p�@m�۔,��I�Ve�-uܳժ��w=����a����5ح�&d�u�Q|����E$�Ι]|kw�����k�)���Ui��M��2�F�"ا��X�p��o��¦�Gz��m��Ǚó������$��p�Z\����r�۸�V��`VS�k(�VHs��{8;88t�t�F��u��=gkaW����؇W/w66��*�v���D^Ýi�w�3�rt�U�^\l;���;9�+�n���.[ܻSK�>�Hj.����V�������K;9^L���Y؟t��E�
�{��r�{�������!yPRE�!��DБ�	 N4SA���G�.�r� �E�}(�*�AED�xB@��-tCA"�A�*J�Aq�I% X������n�J��iS.a�T��I���n	$ieC)
A�Zi��\*NB����&��ɴ
�@�S���r�90�QrD$p����e���H&'a�"��o�l:��I#�R�
�0�,�̲�2C�B��(�@�Q��J��+���8؅.�!t�APg�DbC�L�TM,�xS4UT|q�ULQF�E�#(�!2�V*Ȓ<J��T�m)�0����"��ā�J.E$� PpNF����C$�@I$�)�``Li�A��%��U&�'��v����L�8NH$	 � ���� R
�t"$y �)�`�I���/�����vPҨ�-R$�s�"Ha!I$K��10�i�0�e"���,�\�I
@�N"�j�b@a��F�h�O��[�I$�e"*�H"L�LB�H�FPp����N4�1Dҡ$ǣ��	�xd&$8��*�ʵo�A��ܖA �j�J�d�
�!�P���l0��G�(�q�`�"pd��Xu,�G�(�[�p��1 ��A�\��T�FE��ȁ��!#�@��,�6M T"�PT��� �-4�D�'"��׀���p�#1��M�=J�J�-��dv9��ڳ6:�bYa�:Sh��ݻ�$+i
2ģ��L:�.Q	AZ{i�A�E&d�~is��+���$	��u�#*�3l��:tʻ����(%��d2J
(\�&�;BR�%LtɆ���)�Roe	��!@�I�Pj�S�"A@��NnL7dE\LPUP�aq��)�ٜA�d(�	�A�DPP��p�I*��r��]�a2YL.^W�
����?��0@>��'���@�������>���G�?����<>�����U~ï��_�w�m�����]�t,f����A�[e�
q-�˖�[�ۂ<F�b�uk�Ѷ��)èb�yu�����x]�/XA�)-��3\[4�Ł�ܹ���B��x�$�JmXP�p��.�<�5�u�{���ls��d���AD��f��Μ8'���W�����Gs�f �o�\Ng1�5�-�6�^ko���*o[�m�ҍ�n�H�L!cU�ۃwu��Õ5���_WU�u
�pjÅ݉��sr�|������%v� ��F�h���f�J8wm�3c۹����0�p4���7�!'f��P���u�[��,���_Wwj��˩�}t�Mpٳ:�S7��M75�.�kz�Q��Z��-h�q��ᝬsN�w���t�������7���.���%ؘ#�
86��*�~XV���K��M7��,Dܾc��}�Mv
5���ztZ-A�c�)u����z�vc
`@���5��LT/�Ã��[��f>S���]���t��v���*;OQ��J���+j�0n)ڡ"��EִS��m�sٳ�������w���u�]u�^�u��u�]u�^�u�]u�]u��]m�]u�]zu�[u�]u׎��:뮶뮺�N�뮸뮺��]u�\u�]u㮺Ӯ�뮼u��\u�]u�]zu�]m�]u�^�u֝u�]u׷G]u�]u��]m�]u�]u�]ztu�]u�]{u֝u֚{m�[u�]u�]{u֝u�]u�]|u��뮺뮾:�]u�]u�_c���u�]|u���뮺�ۮ�����/4��.ʔ殰c|`:o[߾�%M��8�+�s��]��ﳺ7�hX�
-�k,ʋ�K�Z�-���*I�A���(����z�X: ##c�%)�vs�}�4~f[���Ji����;�Sb�Nٴ έ����q�d	{����u���n��E6�60��Hw�9<в[���5ۼwï�r���C3�aʼ�&#������[��ޙ�eN�2g.
�Q�z�)w	ե��x����z�_k.��
^.�t��}:uZ�J;/f�F��z˻2%upqz�*��ޠ���H��'���}�l��ti��,vٳN�G:��_fN�N���.vड9ŕ>�b������T��t���k�]����e7���(8��H,�/��7��^�h�Е��V:���yA������ܪC�B�3.�3�*.��6��k"So1|T굛��ˆh�'��Z��r]\�|q�J}�1%�'�]���7���b��%knd�A��KK�����k*��Ur��w�ݭ�Oh�� k:7Y�Vhhu�7N�ݚ��Bsۼ��i�%�P>B
=��f�f�|<M�z���ӏ��룮�Ӯ�뮺�:뮺뮺룮�뮺뮺:뮺뮺��u�]uק]u�]u�]u��]m�]u�]zu�[u�]u�^�u��u�]u㮺뎺뮺��]u�]u�]x뮺㮺Ӯ�뮺��G]u�]u׷]i�]u�^:뮸뮴뮺뮺��]u��u�G]u�]u�]tu�]u�]u�]c��뮺�㣮�뮺뮺:뮺뮺룮�뮺뮺:�P,K�6�-�=Y-��ib�4]��6��B�hU�u]�D9���JG���/�:e-��l����ͳ�"7!�;έ���+��ج�r&��JN���՚��������h��p�D�kWR]w ى�� � ����I���g%��*����^�t�)��E�msMS�����frWh+�Qc���TﲹT��寞WM�ϕ��24��9C-7�k����4k	��w�TOZ���������>ꏂ8���J�+��y���HVI5�W�>z���Zx�7^_�I�'`*W-��B,���j�P}���܎1;]�@�j�8��S��h�X��[��֙J�2��6e�U��@��/t�=�.9tv�37��=�ͥq�v��d��EG�ێ�L���r��	�X��l8�[���
��|T
�� s�]�r�X��to�8-�Xe ��IQ;��m)�t����i�:[BpC�V��;J��W�����+5efH�4.��z<�ݮ�UC��IΗH7ոr��W%��Ta��Y��������v�㮱�]u�]u��]i�]u�]{u�Zu�]u�^��u�]u��_u�]u�]u��]u�]u��X뮺뮺뮎�뮺뮾:�]u�]u׷]i�]u�]u��X뮺뮺��u�]u�^�u��u֝u�]u׷F�u�]uק�]m�]u�]u�]ztu�Zi�]u�:뮺뮾:�:뮺�n�뭺뮺�Ӯ��n�뮺�뮴뮺뮽��:뮺�n��y3w��-���뻜;��:89q� �6��'�+�o�Y*�׶�佮�*�نnο(F��ˍHFm�Rr��<�]se�����W;	�ZJ�g�^��*�5]��N����a�7�[����U
�u�����H��;�;;v�q��H�n���N\�⒩����Wº8�r����i�`�lͷ�c�NPf�t)�}�
�WƩ3u*�#[@���Px�i�EF��S���u;St������W���"�B����kU���ۣ���y�)g9���������f��{���Fnw80.���Ds�yJ��l���Ф��+¡N�c�`�z���ԫ��`��@E��sC�������w.q��m�]�O���[ǧZ�8j
˛�����Y�t<�3�X�<�c�)5���|��[��p��u1>��ٜ2�-Kk4@�@D�\��>��ra�,�%f �8r���׽��KZ�]�
�c��Tb�Ѽ\d7�ReK_���'���ï��7{j����xc|��-��U�q�3u��ن�/D�������#}�a�>T�y����D�PW~���xIo��"N��D��קq�m�Z��e����W������{}ޞ�]u�u�]x뮺뎺뮼u�]u�]u�^:뮺㮺�u�[u�]uק]c��뮺��i�]x뮺�뮴뮺뮽�:뮺뮺룮�뮺뮺�u�]u�_u�]u�^�u�]u�\u�]u㮱�]u�]u�X뮺�u��㮱�[i�_u�]q�]u׎�뮺��]u�]u�]u��]m�]u�]zu�[u�]u�^�u��u�]q�]u׎�N��7&Ug;MgJ3"G�`>��d.�}�۫_I3N������vYk{OG��}J�����弨84�<B��K*��V#��Py��6T�ݱme&�g=�����ؼe"�y,�76�i�j��*���k�F���F!�R�u!1U�l�=��νR�X;�޹J��GF��BvT
�w!k(1��%��1�:�kV_^�{\�NAP��鋤�P��Jt۶�lžS�W.���
E��u%�ە�]��4$j�����LZ��V%NV�١<�ʬ,*Vͱ��8lQ�.)y�
�v���VЧ	���a��� -�2����Av�Q�Z�Y��(x�q����`[[�0A5�.�5�Z��.�����[zk��g�R{���$�&vޥ8��ӷ91Ym�E o��zwWvu7�UY A�����s��;ժ��2��t�{��L�9܈{��U�+h�J�� ��Sj��ق��Ǻ��Q�ܝ��w�ߤ��؝�t�B�ꪹ�,�E��.\�fR��B��46Xݷ�C,�a�*�J�oQ�3�x�V�"�d�]u��s�� �˷���Tm���<��O��Pi�}9^S<B�$j�F�#�������ɻr���sk��Mm�Vq(�{�,�;�.���O�(�� b���noK6���n���3*���L��Q�5e`��tg�˃V}��|wr�uWw6��ҊVJ2+�y�4���]}�/�Cbň�3� -����h�i�f]����T�ǎ<�3��H��:8w^Sc��f`�2�H	��k�nf�B���P�������L���ӆ�~��U���
�E�]\�n��u�c/��n�Ŗ�O�)Ei\��5߽�`�%�.�n��u��>=�������V��1e栘ۡ]P�M[Vm`����� �>�[�O��4�ڵe�WPt���O��뭦�u���@SB�R���^�S�W��]���𺕄 %%��]i�q��2+c�p�2B��Y�䂦egd@�������1JYyu��Sf�0>�0Z�]�7������UL� 8�ż8&��������ڬ�:�j�cEc]��	�mⲤ��3["��N�k/�*��|�ej�Ze/b!��1��=�|�ޚVw\��H�����U�VLTnv9}}V'j�N�k�l���M�Jg�i����qZ�0�5�=V�B+��b�1�	�-ї+/"�ۥ�Hs�5�]�E���]
�QY=��0L\K��k�L��R�	lx
LwW�uX���H��]�.�\����:�䔎*�J�����r�=��6���߽�Rw԰ޮ�Ą��64_Ew�Wg�V���
�I�
Z@on�DA�^l�ur�P�'Dyn^���t���ҹ]��r��yr��R1�M��Z2�_`V&�3;�鋯oS{ �;.����������2�v�}wvp��znkU&�^Q��j�W���W;y�����_�ӹ���uG�n����}[�)���³pX�k��}��9��u��E�3��md�޹ڴ�"�{tΪ�C���-�nj�ҹ��K�(��7JE���B���!��eݸ*�e�I�r!Қ�7����Ku*�N�+�SeD*�h�ݷ�f���u|��M�T-|%��Cd�}t��Y"l
��˕T��Bd|���Q��C��b:�׹W��Mܺ�_����7[�4�#Ep}wT�Z���i�h��,n^�uUR��lC<V�9B1᳗T�K.�ݥ�p��Uй��m��.J�DЭ�lZT���Y|���J�n
3"z�O]�����dwC�Os��66�3�Je)4��q#��+`1�!�+R�s�L��z�}��YO���1�K��b��K��x*>���/��m9�=�B������8&-�+�{{���3.�`#����p��sk.b���v����}�j��6��Ͷ�A"�(���x��1�l����
u
N�߇���c��s׽��W�e�AQf�u9{}C�m��[�芢��t�3g�	OLJ�	�xr�ŷ�)��i�	+��}��y��2�L/�훝�� LN��������н�2}�.�+�˓�M�"�>��]h��7�'U��v��))�Ϫ��M��$�.s��J�ZZ{˜|�7���VX�Ӥ�[�9�����5���E���"������Dэ�-�h,�g3��Ac��rՍ ��jC�5�V*S-���PHA�$k}$��\7}T����Z�J�c��庲����5{��X��(n��*l!>����|��m��,�5�]&���A��mvl���gLq��N���)��3Kn���꽺��Κgcb�� 4�cZ��]K�w��WYfr�����;[�����cEo!�:�{�ŭ�7�.Ίi�Z ��b��gB%�-lƯ���&볜Ӎ,q���c2Y�$��o[6z�u���^2�ei�b�csB��^��N2��	��NX�'ܚs)
:�\����m�{7��h�ԫ촡9�v8�J�����շ�6š����X����Yr�!�i<q뇚���+��)u��TbN\�c��ȎQ}�q��nDO(��g��7�S�T���0]����$��$����2���2Ue��p��L��)�6T<g*���|5�R�GG�rԻf���Q+�<��
���+�qʺ�e�Hc�HεB��֩�Y�N�>OS�J\�dt��Q�yo���D����zб�ە1�l���[�B8T����[p�:��n��=2�ar�fZi��"�<<Ι�4k�1�U&Ҹx�+0�����Z�;Q��kW�� x2fյ{����0$�T�sᯁ�r���nucwT�t.̇�5b^qM�W�S[|��r��-�ർN��|��%\�������@G�N*�`I�4p^W��lǡ
�݆V��ï�ny��o"��Z��E��J��*��b�#���R7:��y���ye���rVwV�5��۲$���v�{���(�{E�x��ifW[U���3�xi%gwnGa��b��b� iCv���7�r��ӂں��y�m֛�NdJJ�NKu�����\�:SL�����bq�}��p�f�<&��]�8�>���[�oR�ooæ���ѐ�!����֭��Et���o5Um���C��'.�t���HL8iu������F�������M&w�u�7B���޷{���'El7uNggs�u�$���D�FfeM��w��B岦��ŀ���
�lu�[���:h±C7R�x�&>8�v>ȥn����;�K�j�ꄾ�K��V��zu1�M)�Ϊ׵lv���\�k���Y;*�=�XLg>x����E)�b�,��1��w���N��o�Z��}��צB�������e=�L ^l��7�:_!���z�\��uܩ	s�Fm�UU7QӮ��H�O.�;ڷ#��f�i
���l/�H��_o)��[�2���9t��ou��{D ���uz�H�M��|(�w֧�,闕�O��wV!�X"ے2^_;雷p+�y]A�X����/�o!;�nB�/h�	��A��x�u7��ZGa��=*T�WA�s�i�q,�����b�^2k�Λ&
��S�wNI����i�=�`�����j�W��\�UNJȆ�f�ڥ(
:+�*�<B�d�ί��Uf��� �������o������?��߿�E���Q�/�L�]��+�VJt�B�9���B��"fN ��!��27��K��4_�H0�,�l�ˬ��0JDTl���e�D
l�`|$М�+�9�/Oe�k��5����JU�YC�m(�s<7r��L��غ�^l�}�^����f�j�}d��O-_)��Jt�
:�5Y]�:�����T#z��&
�����5볈��)AIV��ELf;ܙ�����Ʃ�@V�Y�X�N�u0ol��*�Ԭ��Щ2�t�qTٝ͜4{!�l��Uf#V�2���3���7�i	�����u#jd�r���v�w�*:7��<��֘moS�W�`�DR�%$k��m�+��N�.��CK����"�fX=�O9GF3�aYU�Q������f|iX��bO��N��bB�������5[{Ϩ$�
�uu��W��hh���k�_�]�Rh3o�yk}z����Ϗ\�&V8�=�3�����X�K+�Lu��j�;�����R{W|C��rS;2�j�gu��[�z��[q���Xѻ1��7C��"�86|�+.���S�儎ͻ6�,|��(�Gx����|h�ŪȆ�ú�\ח4��h�׵؅�ڈ�H�.��ެwn*�v�-�����Y�V�1C.a�f���%�e�.��4C2�%�X%��j\&7Q�AQ�	��N%�r(K-���Y	�Dˁ$Wb� �䀐A�$0$\����!�ȓL��D"1�j"bJ&H���IR�5!��ND���FDLJdIH[\l�[d$�%�	�����aP0&"'���^m�Έ����;8K;M���R��i�L����$�LcX�M��:�뮺:뮺�Ǐ<x믞�"F�U����(�ݜ%D.��$��QMB4�n��㮺�뮺�<x�㮽��S*IARUB�3H�K�m�krS�	TȲ�i��u�]u�G]u�]x��Ǐu��$�� �TEI$K�Vy�e_;�_��yˎ�	$��-�T���$1�m�������룮�뮼x��ǎ��N���z�Cr�k��wf�u���=6�r|ml{��{I6�l��v.���	��������׾|ޭʯ{^��/{U���m�v�=�D��籶�y���8Ȯ����[wwa���uW�/l�w3'W%�����*��꬞��eSf����[C]��kk����T=^��k�B��UJ��2�L�]�"5TH����3/������sz�wY�\�kwvɮ�ib��l�v��owGev��vm��w|����k�v��V����3���v������ͩ�Z��u�m(�{�� `0G��3n�IE�"��ŷ#u��cm�M�nF��u{�J$q?��=�9�Vk�!=�ٴ��rS-��y��:"@��d���h�B����Q��K�o��h��_P��v+���v����rZ�̒��X��K�I��hU�t�f{�fc��37���`���yT�&D�j�m��+��U� �u����cc0o�sz�y�u��y]���W�^��B	�����<�,��l�`/�>�9-�����4ߗ�9�C뚾�"�YkeYpi\%��G3=Y[�k�N!�ê�:����qlQ1�!�OV2=�׊*|�(�/�����l��-�>��:5x�w�hR@U���#{B���DMo�(W���4Ĕ��n�����Օ��s���$�+0�f�G��Gŀv\��'�5]{�9�=���_�Ө����LY�*Gͣ,�&x���������{���qP&�P��]&�Q��A�բ�mY.r�%���Z����I�|��{�g�侙]��/_OE�V��vz�7������$
�CD*3{1	�׹����MMR�j�[elQK&�{���==G=[�������!�,0�\{.S eS�@ǴI{�����cQ$a��7M�d��-���5t)�-�Z�Ƌg�t�IB�9�ec�V�y-���G˕N��:�nE3o�A`g��·��y��|�!03����R"ful��)���|yV��txsf��;���1���;���ی'K����`a�3��>^�Wt#¡���X*�Pj��T�' ����	�
Dw��X(Z+��{�=����4f�R��k�7��k:���4��pS�s���O[Ѽ�l=�~�J���<�Cn��e�jW��^uf��(j?M�6���#k!SL�J�Æ��9djk��E���7@�����/�wD��7q�r�njJ�ZI,VK=�qAl=Dm>Ȉ��>���0�a[Q ���zq7V�k���A�TK���we4ܞ(h��� 9�7���4�!�!EM~�}�5y����L�i����`����lٕ���mJ�F��PN�M�1�EJ��UA����u;�@6ʝ��x�>Dv"q�����x@���w�����*R;>&��5ϟ�I�(lU�LB:��:��G�B�/s���I{m�s�n�,P�c�.ۊ��«����:�]�$t�~��#+��ܡq����9꾹^��*��r����Cw��Q�y�u�nS���������J�������|@>>��{oo6��s��Qѐ�� ����l�,&�D�EeV�^��E
�o_��D�~���������6>�5�ڏ޼���\�C�ǵbJ�%�~�z��Y���l;�y��-3w���6�R}�T�A���7
/U�8nvVӃ3s������`Q�#'��bU*����:�bu�y��{ٵ����D�|�lߧL����z�t>�4�H�׏��ei^^@�ͭV�k�ct,�N�{M��ݟ���zц�N�evuI�E�Aૡv@�o����	cW�m1,�f��h�rs5N-�e���1�+_�g��m륗5ݓ�M�mQ��:ǹͺ�9�lS܂,k�"�5R//^�����gRz����V�}�V5���9��|�����W�ؾ��r�xfX�3>���]��T�3�^[
:�'�+��k����3@�%��]F}�4@h���U���kzah��V47����LΖ^���	ְR�g,gbwwvWm�����eЀ�_��{+Ҭ�ۢ�ȋ#�Ǳ]��zl�||||@�><���nom����;Z���f+��e%D����/h���A�w��n��g]^�l�����-����B�ڭ�|�gܣ1yc]�@��Z�䧟�!Ě  ` �(��q	���}���.��K��/n]9��x��
4V��FbN����E��'"�w�0���R-\�ǔq�� ���ʳ��\��=��V�q���%;�*1Hݓ�Q�tf����-��ۛ�9�b�OQ�U����4����9B�O�C�%��r��|TC��:NN��đ3�I�/C�w|���E��{�Z�y�,�s�w�U/H��&|ui�T���O���זq��_ٲ�R�QU��i�}�ݝ:�څ��S�%ᙼT\��
v��f$ml{k�C��c�@��QӚ7�F�	0�m�J�K$k��I;:ml=;�˄ؽ,S��*�]���o��^�/q2U���|r��x-�����vNd��h8b>�-��&��������J6J�0��ѲI&���*��7�B�^�W��"P�(����eӍ��^I{�L���7��[3{��r����ɹ5��0��2z9m�.�.�V��x�G��W"oa���9�4te���[)6��H1�8ɉ�P�ʗ�WE�.Ve��1#�L�!e�O+k�{]ފ�D���e�����BT�hA�r��<�����s9,�k(�2ىlA:c�[�����e��1{�d�r˿�}a�fV�t%��.���#�%�	6�ǭ��E��Q�=$ޑT����������m�w0��q�����2���S��g���BZ�jS�:��ôuT߶�C�L����LCB�\�wY��!�ܢ�ǿc༵ԓ��X�Y�|�Ve��g��93���Mܒ�?�M�k��w5��B��MKeG���ޭY��QM���B��5�zq�S{�wn,��Xa�(>]�4u� �1Ho����΅YL{�z�E/y7��v�<�)�1�N3
5��f֤1z���z�pjC��={rی&�`݈�N�N�p������)�+�7��1�q� �F9҄�����c���d,(7Gĺ�]c�bw�z�;�,�ΰm�Ρ���b�lWQ ��9�2�ܹAL�mem��Hq�*���w=�+YΛ���m�vbv/�u�u�g}�@��x&�vr�ڊv��6�1�c<�����|�<�����z2  ��ԋ��1&�P� 1�J�9t��D�ၡ����D3�0lډȤgu?��G�J	/f�ߧ
��|�#gS=!Kjwij:�u(0N�>��*�V\o��{��n��:������qg�������C|��3T8ʁ&o�P�=��je)����.�ؖWnsu=�&&�>v9�(v
�$�cM=���z@W(n��5�ͩf󣔊H���TL�
�u�����͞��al�E��]��;��Z=�3�=��6ۧ	E���|1�ʷ:1�>��b� :@SYh��}UQT�����Rگ(�^�-v��j�f�ZPo<��1O��@���Z�Z�����G���Ϊ�13Z�7ۻ&I�m�7fL�xTF����eAF��AH�r���r�oջ(�>h�/���^T}��$�ޠ��V"j�ݛ�)������0+2�X֕m�]���z W^��Ƌ-ݮ�j����,T���*� ��[M>X܇����K��̈�r��cV�Ǐ��|2�E�Uk5��C�����yo����������7w��f�ov$���]���6�`��U�[S;6���Q�RŁx*��n���`�"eP��G�w;G�J,i����\��Ҟ�#6�T�H�{BI�we�4�)���d�{r�Ƴ�Jn`���K�5�Yw���bu	́�����6�HϷA8e�����_���Hfb������j�>2����7�� ����%lz� dKU�W��[g!U�Mz�B����;(�����=|�	li{'a��^nz�;lp��ޛ;��.y.��"�{:v?Tc�p�17�Q�k�8����|ʗ���!�b���i3~L�����`��j�%�� ����b2��Y�[�,�:N޶�Oz�؃�vj2FFy�֪͢4����bU�ä��r�Zpl,n��������A�^/g�������������Y�Gcǫ�;�^�c�S^}��Y��uf9�Vm�IW���zը��B�:��q�-#U�sή��w����0-��\{�N���&k��\]n�[c�;Y��A�9��-�N����x���|*��蝹�Z�],>�(yq�ҽ�E-�'t($?���-����Y���N��"ߺ��>�*_@����O?12{���_�T:��X�2�̩��t:�`��Ƴ�޿;���^�-T�TDˍ&6Z�z���+u�j���l	��
$��� �(�g�`����o2��bh��������d��j8�+ͫ��ӫ�wYc�}�[��A���(2��p��y��N���z��S�r�fnQ�4 ��o]��ħN7DQ�)�0��z�JN�ȃ�+C�j}E��1� �B�A�Y��k�Xrc_1�lOg�b�Vc��D�|�'4N�u�����Gw�zDM�r�{gF�X�nJ�;���B,�>�z���Y*��,�[Rk݃ҳ�C��S�ّxI.��\?:��_e9�(���Psu�rd��>��G�q�}l2R��V�3E���$7��y^����VR�_�����%�5���/�{j&�,�^�N�B�-�D!.��ݨ�\�|�1�f��/4�+�']���a�X�E/m�pu!Ѳ���7�NnV;�:w�I�a��K4��Ww(��e̗|���c�0#�(���f̙̾�$����r6��I�1j��4���+ڀM��mp��anͶ$fl0�_6ʤ�-���^�kպr}�Of�^𫯖����]:�9W�V�ڽ�k~�%z������fjI+�'vsf��!��F���I"|�|�cݙ&�܀����>�Vg���+њ��#~�!�Xn�m���ۭ�����R���π���WL�yaF�h�����V�H0���6��Wי����W@ N}�X��27�e�����ܧ��P?o���n��p�W8�z��ob�`���Ya����j�n�<v
U+�>�a�!CQ+iO�S�C=� ���et�f�$Q��s��s������(�:@+L�k�+����g2��|�u�̼��qu������t�."��Z���CA��Ya����%C$�"@��m�ϗt�g��le��;7�S�j�=H�p4p�������k��ޮ�zOF�ɨ^h�s�=�Eڽ�6���OCl�Eef�׽Q���ݯ��&�i�u�uЫ;��2���M&��z���M<9T���_f��;��h^�������x��wuܩ�Ͻ.���(mJ��C���^݉�jR��fP��)%�w^���A P@�3���
��[���*�8 }�&���G���.fU�o�>Ҕ�����{��Z�p�����U�膆�wˬ�(�Ԏ����@��6�*V&��4�A[��mhõ�T��wI!��A0gզ<����p�&�D��6z��pm��NR�wn�p�:�}Q4F�^���̝�xfwVăs�SA+��Pl��a3�])���C���ˁfe�f>Hv�×~#P#s�7~���}�w�~Kvfrԓ�yeU)�Zt��l�1�����.��e#Ǟ|���&M��-�[s1z��J�n��H�4̀�Fi�k`m0k9ǟ/\+��׻&6
���ν���$ ��,��@/��:�`*���p_���G�+�����B��w�;�°]~�6�%Y������[:��^=�i�:ʹ�h�B���.Kɻz�]��I�z�{���p���`{ӥh���;Cuؔ��ו�F�]��5`넞};:�D�
�FWK�L<���7NLȐd�c���f��v�k�T��Kd[�ˎ�$�'!u�㡚��'�Q2+��۾x�]Ý�%[��].%����4�-<.U���i0dƱ`�WN�]I��)V��jm\}w6N��K���������1n��UM;����0����e�cQ�i/z��1"�;k�a�+�����=��Ji���f�V�T8��wG4f���U�Es4E��gn�ǭfU<�:^����1�C�e�g.�p��[x��1X��V云��V���_=�ݧ�y��]Z[Gi؉^5/D�l�.��qYO<���P^�"�X�֗N�;�+��q\����Z��y�%�c)�r�Xv���1Q�T�XǾf�Wg�:h�$��(DБt�3�js�V����y�_��B�f<#cI#�U�۩Ҽ����t��j��{�&�z��M����tg*�e3��[D��;�����eu����vܦg)6��KVu�f��U-�r�S�:�l�
"�<�{��۲��'�ݯ}^�M��>��AH�gR�����*�6�Pqs�����B짱���x�t���]�w��2�[5�4��ZlS~U���h7�8�Ԡ�{�U,$�>�n��<V�nV�xA�x�fGݸ�S����EvS�m�Z3�WV�*1[��[8�u��<�ٗd 4Lк�Yr�5*Vކ��a1n/b��r���6��z�o!�8mmA8Q�s���jLUp�¤�uƍ��{�A��WwL�ˮ��.	���VP��Y*�W�:l��벡ؙB �m�>C�Zͽ�9Չd�(�V Y����*[*l]���EV�j�ʍ^�T��1�X5��fTe���6[w�{��7{ump������;�w+:�b��q�E[�s����z�]onQ�"�w'YͮU'A�w-S��;��ݸ��K����JvUݲ9��`v1{��a7UV��m\��z�N`�r��yכfK9����f�To�<�b�����>"u�����& ���}gk��Z�w��A(������`��Ʈ<hP���,-�0_B#*��q�[��>���������71�e^.�uv<f�e�o�9�R`�����}c�xI�NA�,�"BF!$c��F3����|~>�u�G]u�\q�u����Ȥr_x�#�N[o��R�8�{X�7n�Neg��S׏�mǧ׷�__]tu�]u�q�]{�
�#!"�BB ���\�@v�mdW��q�co_____]}_]u�q�;����E�Q9�~]K���Źܕ�;5�aBzQGiAP��W*N�i��>�����믯�}}}}x�8�Op�	;��:+�����!á��U�̹~m�ҬN�Ȅ������?׬G�J�*�-q$���ni���D��sn��(HN$�s��@����a�V��++@r�裤�3.�"I��{n'2��U�{؜�|��6�-�NA�gmY�3M��6�e��Y��A)9��N�收�[Y��v�8�\Ye�vu�'�D�O�$�H>UB�f��u���B�g=)o'����1�;}n��棭�_=±ngA7��&7b^Hzo�.wav�W�����cM4�M'I;����y�o��� r�c<0	��2i�$	��?�6c�p4f�=� KՂ�=�J%rK<�"��\��A�Q���l�� haM��a���2�ٓ�T��r�;�c�9�Bx�I�`-&ÿ<t�R��=yzgQ�<j�g�R�� �4y��F@3��`��'�Z���&�`'�b�&O�� a�q!�n֣W��j[5�ِ0�52��*�ܰ�!|����9>@Y�n��M�_+��W
7{�ü<��ija=Q�AI�?s��X�`�����k���W/�;�x��|gʭ>$����
]���qp+�O��ʀ�"�U_,�����1��bX�\�[��W�P��xo�A��n��mP��S��w�d��Y����=� ,9\Ql�Ƚؒ�k����>4'�0ձy鍳ƻi�8�U]�U�ݼ�=�!�x�@��SL�����=H�3�=?'�0��������(��&�����s��[�P�2�~0a:=�<1s�_A�5�y�z`����Y��
�u��c�s�j|r�S��A�<����<>` �̛�^�?���!�p)�~ ,~^�B(��s\<'�/�$_bށ�ψ)I�W�������C��Ƹ���lYZ�ru1J��];��;GJ��Ƃ*}z��N��Cy"�
Z�M�a�S��]Nn]�)��v[^�9��CĻNJ���]�.p�]��	��ƀi��i���7�{��^���Àw˂��)�;��T�W�i)x[EL QR�����X�M_T|�� z�KrRZ���NDv��|�^y�����y��9�j�p�
�V�#�Oˤx�i���MT�:�U�YV��{�g~�d�[D!
�_J�R~r���W��� c.{	�PS>���A������Ƈ8�Je�D�ej����{�0l�i��B ��+=C��������F��4����=}@&os���w��4uPW���ٻ������S?��p~|a}���j4>?���mx]z	��Ip	vd�䡛��	�n��oj�����z� �v���������)rp(�PA�3� �N�ߕ�߸�үM��P��ŧyY�� u��QΣ��7�8A�i����y:��_(/�,��h��Eu	j�� 0*���+���Ws<�k�i����I�=� <�]8��a�L ��,��3�>��Y^S�� �1`�� }��zg1��lC��
���p� 3{��-�^���-����{ H/>��8�e{݀Yty�!9q��>��.
����3'�\�f=��ff`���hr��&f 4����C�u|�7������^�OW��\��3��9rdO���h�������a���W:��:���[s�ϓ
QRs��[]nM��Z��7�"���$��mў�%8e�$$4o[�v�{}�u�D�>��*|�`�qf){��)���:���%�2D8u���u������t����N@�	��L1q����m�Ȉ%Y�ƚi��iF�h>�^��E��n����ˤ�BE!�8"q�d�~�1�����-phb��gǿI\��1<��>���`��u��4:I}�9M;]gj�����7�p��kh�3���a�$C�^A��|m5q����F�A���I��h�������g�����sg�Z�Q7I��χϦ��Ԇ����Ctђ�Ip��wXXY����xe��v����9�e4�l���/@%�n{|�i�?0�?/��q�GBu���s�Uuf�� '͍m�M9oc&�<_��L��S���;��;ި/aC�h.s��7-�Mʳ;����y�]?	�Es���:.
�@��z�,-3m�c�����[O��O��w�`�Ӗ����g��K�� �����`���ǆ0c�]�;���x�P(��7s���I�xH[}�<��l���6Q�ď  M�B}ΰB	@x.x၅�Q�q|�*K�}Ҽ��*�����՚��Kʩ�MC��z��ov�=%���)�����3gE�tO���IO��J������7����2�n�q�s.���;��n�r���w�S�� .6c�J``��'�5�+�����/B�h	� �_{+��("?6~��j�������un��$�z�������|�h�mC��_M�4Z1k�}���G���l�#*��􏭴�uk�}G���:wX���p������N���z� �#�n�M����@�y� ������^^{���.�G��p�`��Z}$f�����ǁ�|7���D�qsᯂO��@��u��oN�ow��.��ynl"�
lO4��U[�aJ��}�����[	��K:�$犔J�;Kx{��ȏ���!�������TX�>
�#�Az�û�'J�@�&M���8���Z��66,ξ�(�����P�S<h�/0���)�+?}�r�y�
���2�ޠj�b���r[�8I  $��fo�|;,�9����n�lc{��j�6Q���D�G��b!%����y�����S��\�6��|e�r��|oqQ�?wH�c]��{g���Hqm�O�09�_����i��={&�RV����E=hbu�	9y����D3=�X�\Gc�c���[�M���#W]��.��C�&<�����s����f�ޣ;�l�.�-!���o0��������I�/-��f��Q�> }^��C�,vd��W��w~Z���'�$mDŽ=�%U�'j ��!E��	�U����7��K1��<�^�G���|������ fE���z`=@}Q�t�z_�����z �MwP-��w��
W��5W�4�t\����	��ͻ'�<�vǶ�w4�3$����u�ө��T��-�љ�4L�(�R��|7�c����
�yd����%�Au�n�yI��Z�݆gw�v�opgr
ЈNPf�LR��}�����^^�������q�Y�If�����)���
��H�!sǌ ���G��n}�7�s��Ux��/{=]�������@E����@B76������/D�����x�w���i���.�KOf�.�չow(��倹��US�pܮ�f�6�+L􄏼L���>����ԬƉ�W4�/8��f�D9m����׏K{Ӻ vQ4= �K"���.>��K�->��}�^V��;��(��9�HU��:�� ���2�\����~պ�����!�Jw�G��f����rqn��y53����M����2��d�|9� Vؕ{ &��!
�'��2�qOP�kk���9��3�K����@QN�����a\_:���/M-]�>[3U�qBu����!����$���X_Xg���s���S�����|���f϶�O�������Ɲ�έ���{,?��](5x��9�%8��f_����<'�f���^�H(���P�}Yo���yK�߻����N�X����ĲN�D��=�*�{�7���W�
\�5(S�>};��v�_�v��wf�GY���o��z�{�������;C��Qf*�K$�֠y+U�C�7����͕�m7)�WV�#j��pw6��
��%�5'�L��s����쓚W����5��4�AM4�O�rII���v���������Q~��S�X)��y�g��t����E7w)s�L@��c��uNe4�|v����{���;�@�u�5��E��ҟz��O��L�P��`Ohn�LXn,r����q�$��;U�}�L�)8�$�3�?��o:��v�ok�^�88��Xt��Lhj��o_�
Oy�o�Oމ��'�p+3����궤L˕�����cu�i��f� =@%;�4k���C�xF��gs/�%Ol�����ے����{%�{��	�^�{��|��6���oB�I�Y�����!t�_�H'WһR�*������y7�6����5�½\�L,3��c�G��kӸ�`�S������̌��wW59Yڧ������ܿK�Ń����<�3H/ڞҏ����[w���# m�	��V�~޷H��n�g���4F����$�.��6`��{� ���4� M���b�׌/��'`�۾4������ᩕ�iD
��*$J�V�ָ>?m��;�������'fLz;GvV�C������'��9�"G��<:a���"ZD	��L��*h
7��.eM����4SM}~�^W����ݧ+:������ڬ�:=ݷM��r�mj��BC�4�у��<aI
Ɋ����E����7x#<�.Y��{-���'���FAJ�,({;*��Ɣ�,�v��s�f�E�o��
�
��H�QdD�n�&���
L�� 4�~�x���b��m-���m��$�H�H�匘�Is�{�^n�%>�b�A>�[M�/�g��@��d��>v:� �@J5�<CV���qr�%*��Bi9�ՙۋ��m�?<�fa'�W�PHσM��ՃO)��,lx@��wK�7b�un��������F�r�'MM"�  �Y�~�VU��k��*T�}{^�~IJ;}��eZ9ư��n|��"S�J�N�M.�mnc�rѮ��=0���$_*�6%Jf�S#ql��2B�G�[]���=��~.Jz�������>Al��b���gbS��r�ݵ�z�WQޝ�=��������*/ٰ<be��}�ට>
E�{�����x����ո��(=�5��&�vҝ��Sa�R(�EO�s^����9�tE�r�c���Ԇ�����lыKr܇fˎ腻���OM�t�o&I�E�`s��4���r��`�[W�8ƍpbnu��^j�R�-nv�r���-��2O�r3���vf������;�	�������O�*q�Q ��|\'	�x����Ʀ�e�����5���rzA������Qai�`�O�:�X&��k���߼�ֲn*$���ץ�ѨV�{z��5W�%�o���#��Y��i���d�F܉��ܻWt۹+��ӆp���cC�W�T6d�K]��d\r-��N��S�ۉ��K:S[��.y�6y��ג�W�FE�ǦĶ�m�F�m.m�m@��� f��f�r\�rG��`���|�W��0N1����j|+��S�'g���`��U':���q�;��UE%�6�/w��fS�֬���`g�����#�PR'��G����~w�g�k�)x}y�u'9��g��N��ґ�ݰ9��Qay@� /F0�C����9v�q�k��K��P\UN���ջ���z�R��l`uC7k�J< -�^v�Ξq�y���2*<}D����ww]����yk�-���S� �2��Ǟ�O8~}D�ЙJj�˱w�^���=k�\ǚ��x���<�q�`/R�j������@3/��1�y��M���}�����'Y�+_a�9���ON�f��?��@��x(x>�]��`�r��P��q�~��x�pM�q���畮��	���p�{W�u#�|��@a��h�k���Ő���h=@@�~(�&����~�A�<9��,@����!w#���d��E�+��q�����2��_���|�J�}����s�Yƭ�O��g�����V.ռ��CKpFa9�
|��{�����c�E퟽�{w�Hh��~��Txsv'WlD��w���w�uq��{N4t8���<�__V]�5��]L�i0'��z� �*��^�v1�������Z�V�Ē�+�����׹}h�|-3�sF,s�^5��G[����n��� \����8�|m�p [m�p�m�IH�	}����_>{�n�����!'VĲo��M���o�,������Uֻ��W����c)�{	������y2o���V�3Bё���_=��\��S"����a��=��������W]Er���\���!p=�L@��yݚ��\^O'-@]&��L#���z���A�[���O�K�T��Q�H�L�in̏�����tF��x��`�֛�"�� �VF�Kz��h���,�7�盔�[�-4[�G�$:y���1fsU$���^]#l�|�0��֙��F@��Hʡw6� 9��7-qV�
a�{R�PoA�{s��S���6 �#c��?�s�2�C�������L��J5]��%&$�;���"��� ��/���פ��5�0:6��<B������KAj/�6��w�pM�O��t�c�ϙ�)�8������u��N<t�	�P�h��G����˾��k�t�TO�G�o��8�ЁϠ��{r\���y�ڴ���I���hSz�U��Ѥ�ݮ?�Emo�`B�C��?|�Oq�+��y�����@<D����w��/��n�e7��=������v.̱֕B>��YQ��w��̖���L64ڥ�U����ď��/�h
�w��i�e����Y�w�M��Y
l�ν�v�\b�ۏ��bl��4<kTas �X����x{����=�m��-�۸	����=�q�GqTW$�E���$� F220��GK���|������`#���<��<��J��y�,�_�g��0���O�Ղ���u#o��4��9ǀ���Pr^���r�����A�Q�,XB�����������$%s���1�U����3oH��*3!P��#��z��+����$����𰢽 f>5[�sa�f<:H����D�\D��Vnn���&_��7�1�o��I�%���vk����,O���iK��), �#�����{E?�gN6ýYE=��Y1\�ؒ������jc'��9��}j>׳�߷�9�[U�5���I$Q��:l;� k�, ���������ȗLRs��s�=o����I���8j|#��{\<|]@a\Ĺ�FN7�s���Ɉ��1�:`;�=C�.i��?^���=�������4�����K��4�����.?�����Ϙ���s���mXr�vN��/7���X<;$|@�/�w����:��4�Vx3�H��V�vY�uW
ǀ�zO^�\�N[�%Ķ���`�a�8y|��{�Xo�]�wT_�	��Y� ��{�����Wu���n���� y��[B�.�}8]\�+������mdmk�i����R�fIb����v[4؛=*�%u�[je{yI�_t�]-�¤I'�˂{j�#�/��<�w�ʡm�U����!οk�Q�����Fa2<��w*�r�3W]�I�\^�O�_]^@ZWЖ ��e}��^,w�!�&��F]�5��v8�c��n�Nmd�X̀�E�r%��Ӭ\��Λt-7�&
�<���a���'��kIX���&�!���{o�T��9�t��C�2nn%}��fG�+�^)j����΋	����Y�(��w��b�p���ǲ�2Z���׽cQ�/GFͧˣ��b��73J0��C��^���>V��DJ�ańN逹F��=�W�b0A����n��#���&�{�M.�oAݽY%�,г3�L�o/U�vc�f�y��T�����V����Z{��.�`)p���yyq8�Y�MŻlN�-����=� �0�%^0$���(-�$5˵ڮ:\�3�{ٜ������[�B��]���6�At�'jX���d�h`ͮ��[��u�f�x:�h5t8'����"�k����i̦6�07�����T|$Z�w|h�*����)AI�ڦ���D�(�q*-������QH�
�,]�2���D��N�eJ�Z()rd��^��K*��t1� �4�Ѣ��j�%Q5�iQkOq[�S׸�af��TJ����!z\�Yx��.]{�{�V�a��q���}z�������6�iX1湜�mZ��N�]z8cTUUy[	-�v�h��������X4n�v���Rz6�b�2��:�#��9}ǫ_Lidj���
��#���v�b�`�ʕN+�CY�-���s���{����uv\E+yJ��^u����!�.m�2ү��޵A�j�榵c�x��u��!��7-�m�Kd�7�V�y�[�o;�w+�Wu;;J=І���iJ<���1Q��s$�����*���_<�C�y�w��s�SB$by����(�X��ٽ��!�mi1ఱg1�����6w��z���T�͎��]˻��]d��oY�:����+�q��z��;��yaO�����2�ҨZ�����]��\G0�W&��T4bM�i�wk�U.ʗή��2i��zKTo_G�������dP���.�]uƗi�#���;d��u���oseA��Cx]���{��L�s?��q_#��<ڀJ��[=�j�U�Uo,��g3m�����0�ƁC�D�fH}�%�А(�ޝ�\�4*F)�G�q�}�Jq!�T\�AQI�3#j%!�MP4�$	��d(�L锢5P�JB�!����%b"r�)Uin�*��%I��Q���5	�PlH��
�Q�M�	E�Ad1A0�d���$K�C,�RXp�4���G���g���4�(�PIDD: �4ډ�T
�4��6?p�^ۢq��h[�o��^��,wm���LM��<�B�'�6��|}}u�_]}}c�����q��׾�$'uR����!I�""88��M���G$���~w�����뮺�믭>����8�>���i$�$)�u���B8*�����5!��`�$�$'O�6�Ӯ�:�n��]}}}zx��_^xvU4F����ATU	s�r~�̡	G$�I�!��m��N:뮺�ۮ��]u����뾻��{��N�v8�#�f�
AC�b"H	�H(�8���wV�s�嚶��9:I�D�v !�k��!A�	�'ݻ�#��NT��lI:���okrpRs4��!P��W����P�kn�����&�t��(�)K;X�ݸ���grN�ډNRB�ۇ&b �Gwϛ��v�6��8S-�\G9(��8�"��Q
r6�.*QPA<Lz�UbG�ۚ�]d��<��\��s5=�<H�}mX޼|���2���o{w��;��6� ��Lf$('M�����I��E'�� ����Z�H�m�$�m��m�7$@VE�w���7�{�:��pad"��'�(���F��ƪ/�7�_H��X�,6<^ -��o0�6�S���6�I�[e��ͥ��D���A���ߓ'���K�O7���s��ɭ�V�#��u Y�	�1<��f��v@�=�m�נ��?��5�Xi��q"^�����U<�{��q4Ec8�,��n���<S�&�p��#�Ӟʖ�%���xNF�>6�3Lzc�ǟa���xD��;�$�� ӑח�Q�=�p"L�}	8��z %�V��g�5�@;��J����Op;"<��r{��b��b�q�<��w�X0i�u�q VƆ��0�bF|of�h�5�7�Qzw�
<(QP�c��͇j��b�=��?��\�z��5�����F|l؛�O~$��zŚ��x
�҃�&�}4ޖI��Φ	����O�� ��.������Y񖰀�hj���,o��I2�6�ݛ�Q�eޤ�W;+�yW�� ��f'�r�y�Jܰ4����(��.����|��+���
���_m�*�$.�����A>�w�{�ΧU�f�̌}�/�\#{լ(�a���@l�Y_$ߐ��7D :p6]k�������;�{V��0q�ha��G�ξ��c[�0���z%6�Wb���n�qS���Iֶ�;�����!�9��|hwu��ʻ���[뛤�̨�@�4�r�R�������DB�W `�]�꿅}I���R���ln$�,m��m���b�Ȣ��9����|���L����9��3�\�;��A�[x�;ݦFb���� k���π�<�h�~O�;[K{��8�=Ti�L"�LW{�p;���ś��b��w��Spm�c!G�㫦�](;���0����%H�B�7�Ȩ8����5��L��]��W0�&Hڇ�p��c7G{�5�J��7��`� d`z�T��2.58�zKo�mn�u�[ |\�l
��.�JъL^c��=�h~������hPb������:�����̱��Oe�pW����K`��Gs�=3�Y3�ە�Tei@s|��̦�k�<���l��m{�#P�ɜ6�4y�U��6y�W��A~W��ySQ����L�2ϩ3��I�#BS��M!=k�`+|�� tL�{��f�a��7��Q[=�����&fxi�a=�%��p=%������	�߂z�z����nMUr��\���"}R�n�7���Y�rB/�G���T3G����3j���c.���[�{Bp��S�gfarְP�j�0�>#i�c_���|'��͵�^=���#ç��-Q9�X���Zs��y|��+�qC��.xn�;;|5ݸ݊�v���]^ĺ�O9�҃���1��r��1�������q�)��{(.��qAqVݚv��37@h�M�k��xy7��{=����l -��Dm����� �~|�~o����y^F��u���᠁� ���ȸʂ�|���w��܅5���d�267��Y�=�ָ~�@0�.:k�P���|$�����5��qQ��G� +q�cu�7^'�����o�y������� H��"yن��(�cU�i$�9��Z������n�ct�q���y3K�`5�};�L#�?������UΫ /�J���?%�Z�m��ͭm-qS�����1E5W�p�a~�M)�@���:��X����eiW~��U��ŗ���O^���:F����p!?��Dki�A��<9/�<���ܟ�\���Se{�P�7��Z�ˍ�4��j����x�=_%�叜�\0/�@����<Q����W9b��v��Mu�Ϸ�׽��sښ]?Z������	��a���'Z�8���l�H�'�ˁ�M�sҦ��o��@{S��u*���4�p"]�}�O����и
�Z�l�O��z#����%���afGI��x��5E��7�T��
�#͗�-�6s���[�h�|s��y��Q��Q~
^��c�+�'w��P_\��ݽ[ra�5X��`ޝ��0�p`���EV��fc�2�Ê֥@���ڕxx7sk�'P���T�ph+��saJ�э���<9�ֈ�ܶ3��-�w"�+V�/�_}����o��.H�"$m������m�����Ȁ!!��o.�\pL�:��>�6"<XT��'���
�y��( ��r%=v�8c�X�<׎�]�����+�:R���Ԫ ����6�L�@es��;���
�B�&�Ɲ�"o��9���.�~8�'s{���-���">xE�xJ��r� ��\LMyS���屻�o���oh݄���R���o�=Y��ݤ������]�K����88���Q��_ߔ��
執���;��%|Frݑq��Y���K�ֿ��>��"�PT���LL�L��
�:?8jz�P��\�zhX��I�~1N����x���PCG'0�į(>lZ}�)�+�2W�p�PN,���g��}={/�Iv*{�U�ɵ�@G�z���@�a{���p"� �yS���o�ޛ���V��8t�m�hn�U�9T��{kxOD��v�dk]7!7'\���ݼ��s�w�X��μ��p�YA�k�����X8�:{5�O!��C��-U$����~ w(ߦ���SuouslB���HS-W��V���ʁ��u�0<�@P�"�OHv ��'=�MF��ttr}s	�������-��XDY�zj}�j�%e�]�]�'Efň�j�� v�z��9��o�з[����-�[C �31&@*P$-��g�)T'��I%�`Q�^�S�(�������M��]�z��]n7�!\R�=�'k��i��ȒOE7�ŠΤ"5�v�� ����^r6�1���"�8�lF�B�dA2�ѕ�^p�̒�7�>�:��z~�Am��B�m�P��m[�� "� H��+�g:ܯ����+�����O�8W�|����*y�C�9���^�X�#�Ϣe�]���j M��k4�Vb���ŋI|/I��xkvriH�0�Lx9��sEn������?�~�ջR�U]�K�'xlop&�	{@���9�\
|�Up��N�𛍁qaD?�y����
duE�!r�0�;��&�2%=t�����MU�=��n�	�M]P=ʪ[͚���x�.W�3--��=��)_>���*t�����t���������l�ʪ��[=�z���B蚽~�ȣ�|I�<�?�^z5��3���5�ڨD�d�Ao�ψFi���~t��Q�}Q�<S�o���ӝ_Z����,?v<�K�[b07����Cc�(�������4�)�ȵ����OB��8@��Q#�.`����a�_��⃣����v"�|�y�"xD�HcN�E���)��� 0h��Θ8�WNz�&�J���I�f �/=s�/8��U���m�k���%�_+0����O/z�.<��Kw��q"�a:�@A����Ty���7W�x[g���^���Q~i�멍��j��׊`n.0� f��9ޫ�^}��_��OS*�c}$�ߺA�N����Ν��W0��k�'Mq7z�\ܭ�����lu�o�Qf�X��U�� 6�E�`�M�^w]��rm��o<>�C�o�b�6�hm��"[m�őP<_^�ugpE�3�}��<�{��0o�QM~�	������+`TS��Μێ7��[V�9���Q�<q�zr�����)��Nt)h`i�A��L�[X��A��8�E�J����]<wCUv�Ӽ�:oݛ����t�[<3�ǟ/1������CE!f�-�ޭ�K	i�L�cM�(BuO�T�������'g+���s��d
���x��/��CX� ����z�ue�u��<�������G��Y��5x1p(�;ݼ3��f@��@� ?6��S*Q���eJ9��8LSqu�`}�M�}�/uD��A&@x�@���|K�:&\�ϯ����n��^H0v1��b�f=�ni�%"U\�xM:�M�.W8t �P��v���R"l�9�{�t������C��	�>K�~�&<�����B2Ӎ!����^v�����omK�gWLܻx*��Ž���0�U���3�&>P���-!����_�<1��ԉ�v��O�$���)=�٤��ي�-���O��_X��I+�`�@5��xx	\�u�,�F�'낦���ϵ�Ǿύ�Kʬ"�_U賦��:�s�~skxpaԯ���\l�)�o��������2_�+%�K�H���L����jr�O�4k��;t��|�N�IϹ���fRp�wDk�`�>���+��O7�<��;w�`D����m�@��m-��Q.2$�$�"+����8xi��4�_����Q��|����lx38з� �\'a\��9=޷q�9�T\3)��8{��fg�������u�<��,��S��`p���XN���8(���"vc�o�pA����S�����q�H[~ �)�1��px�"0ng�p)R�W%��M���<�3p"�`�|*���	q�&e�!�h�ӥ�L���\��8<+ϝ���OW}���c����p�*�Y$�>���/֙�b�8��1a��\��1ϓ<ݩ\$����Ø�:����NW�=����n� �>n�-���(��!d���<U|���>*�y�&�q�ҧN��Á~e޾���y�+�sޜ���y������� Ր3�P��-���@���������㬪����<��7p9�pލk݉/���L9�w/u�s���^����[��z���O;�=ۖ�W��޸Lo4ځ"EG�(��c�y�ע�������N1�f�.N>�L2�Os���p�Sq���x<WQ$��lAoǞ0uD��]���P��P=O;�k�&��,�>fT���wot�YY��ڹuCOC�)�?t�굞��f53�JHp��%��У�+=�kC�L�y���ޜC�9���a\��u�y1WN�n�e%���*���T���7�SJ�{s�|�n�>��~�P[m���m���m��Ȁ$ �(ȃ���c-.<�m>0p���0'� �" sd��|%P<�Mǔ�{J �}f�����q�{}�u�)�<z,������qw�@�߼B@��\w��Ό�o�}�)t�t:�^k�4��^я���ge��O��>�yG���|}3�������w�4��F;Ǒ���l`����~�1�h[8�~�lvV)���iQ���a�� �߯�,r����5�'�{�C��A|8�	�GX��(�^B���[;��U�����fOm���^k����F�1���z1�PY�pXE�<�3o^�x�s�wp��5��q�d"���)q�WV�6�:�j��!���p���g���4�Ϋݮ���9�SI�]#����nzXL����@q��Q�f?j�����{��[�qX[U��~��>D��-P<{n��L���A�����~�_/����>G�8���!�o7�p������e�V<���AC�P���- 3ง:F�n�u`�S�2�|�m�֑�s{��ffn�P�<�[�;�+_Cg���<ɬ$����9�������]����)Q�o��(b�6 gZ���7NZ��\ò�q�&�Ol��V�^�Z7�`۪�nN����[�%��]H�,T��(�6����J$N��xwpt6Ξ��ȭ���na�g:�q�b6o;�&\�L��5�m�.��u����Y^-;��e4J��1D"LxK���̻�WEK�s*ʿ�D�����l��m�D��lB⧀�a3:�?_���l�]&_�<a�At¶��%L�EW�$�-^��%=��y�c)�[ռ'�veg���W59�k{��Ϡ_,6D@Ec0i����z�0�\k�)�>�i�H��8�ٶ�X
2�J+kwk��,}\���p x..��u��s�����x�7Y���}����/N�Zf{���4{jE��d��$W�ɑx\C�,������G�>�	�S�ɖ4pvMí��ڷS��K^��T�I�>�G��fלpw� �s�T��D6ÇN�+r��M<9�j��Z��n�L���=�9�m��� ��&����	�s2�l8672#q�	��+n�o�Zs�+bZ���N���dcx@MѾ���������W�j;c�+7r�k~�9�t'n���2%9��-�%���������@)���c�Q��a<L��p�S��W}����-�uJ�#��(C�B��N4u}�8�R���z
��,p�k�7s�1�*gZ�5<�R��M�����-w�[�.��|>Ǧ�ڨM#HD"�M~]~�k����l��5���߸���qZ��e�",N{�ot�S�w��8��v�֨�)�o ������*^��ZjŃ�����CL�g��m���	�:JF��CQR �M���6��lJ�p�|�X�6�}���e�kU=w*�S��:��i�o�U=�v�����Gem����(���`	h��� [m� ��m�� �P$���{�|�v��O������g��mA�5�^�`���3�R�rߢ?z�6���jtV.�1Q�9����c���Z�Ļ=K&��fB��PW� �1��/���	O�$���9SUY��kBr��*vDN�z�=�?p����S%�WM|����f�D�h��K��ޝ���1����Xpu���=u���K&�o8"�`zX�3�z�D���7%�n��m�(���-���ܙSȢ{�����Cݽ0�����q�sKUd^x������Ec��r3��fuˎي�4nŁ^��^1���X~�{=+AgqǾ����C���n�H��x��!�x)�=_G6ݜ��&Eg
σ�?����4K�=�ODXf"�MM���[���~bS��g0���q�q���h=���
-�ca�)��L?�S��9��,��w[������}�@�%����[��rT(>���K��Z>xqnm��JͿ������V=FKM�}P\M��B�9Gɽ��a�{�|e�O+��G͢�zW��=ү�|�WFݷX���هS�7��-�'5o(��
=�˂K��nc�X���.�ɒnu�,!�-�[��:˳m����ƛt]vj
�����u�s唑���C�|�Z�O4Ș�D�Vm��α4&��J,��5V�X�9U����	v��饙�Ү��`ي�n�w=�Ex���i�%A��j������#[�MCE-����ld7��֛�;T�1.���a�8�T��l�n��^&����Wd��F��;3M+w�Ou`�n�]�\O�,�N�{�P�J[쫫�In�g
R�şn��v5�Ϛm2_-O7i�֠�}m�v�`Gf�c����yd��Ң�޹�^GTn49�I,��4�j�7u3o�-�R�*s�__+�������hS��t�[\z�D��Lȉ+^f��<q;�%�3����|r�֞��C�2;�Y�j��$)072�[&SB��4q��C\l։9�d����.{&*D�o����������oF��*�<o�A�;�\��� ۊ�,8��a�2�]��N;�o�[�ÍMꦝ��Q�P��/_F�Zf����^���q�H츩��6�w�w=��{;�h�`�o���Ŵ�c-�f���u��n�b�b�s�F]�9�Ď���>��D�륅�c���B2��nP�\�Jݾ��'7��eV�"L~_M���sֳo��>Dgr���
���agwyL�Eohy7�Zj�H.n=�k�-wǰorFcw���k"�o�f�6�W��1757�,=�EMk�n>�� Y��<��a��M�p%W��VR�1���б��͒��|�0�����	�s5��S�{��&Q��CG��ȡ)YB�56�JM[��v�vn�>�ӵ��@�q�6e�3]?� �9s{D�e�Ƒv���W�+�NE\T��R�m�Ώƅw(2��|���_)7(�jk(�sr7P�)G���}��:s\D*s]�x�Տ)6��]��v��l�#������$���]�m�G�[�5�5-gU��k��c�ˡo �|	v��u�PC��ec+�()�R����t7��M0Պ�ؙ�kh2#b���m%���YJ����yʛ��S��H�R �J��ɢ�{4J;xCb��6N�f��juDю��V��N�y��z��ټ�0�flś8r��ds��յ����^,�޽{��ؼ�!�\��Z�3�@�X���3"�O�r	�����T�n�Ťi9��|�-B�ԩ���}?�_������lE8�%}�/7I.�8�$N�T
�C�
	.��B�Zm�|u��׷]c�����Ǐ>��1�A���@�$���(R:T� ��:������n��뮺�ۮ�Ӯ���������öH$N�G]��(FI$���Y$�`����q�]u�]zu�Zu�^>�<x�����I���2�?�q��8N:ߞ��t�~�[rD�/��4�%�m�u���]zu�Zu�^>�<x����<�@���BwEN�s��[�R��P�?=�9 ��s��X��;��v�\w��$�]�<�XV	���y�������!$]��9����tEP�J���)���rRRm�$�8�J�Y����R	�Im�$Y�qr���9�?��5����;��O�i'_k*��vs���@ �> �3�q��37�L��̸d��c���Z����+��G	||�Ք��Ÿ�w��vZ�;}ʹԯ������[m���m��\$�m�� b17����s��>s�7�A�67x75����"s����9cu�ú-�`G4����K�ܯR;�H}��8�8�����6qm,������7�|�fz�
��7��Z#��=���t��~��81��B��E����q��hI��Y�ڤW3�qpk������oa<|���=^��T��MsU��X'�|%xu�5T�,��D��8�0^/9(z}D
HT{O����(�QF)1!�G�~�l����^����0Jz�l�<{B��4G3����y���5o�o}0̗�W�ٲ��7c}F �2�б�;5z�!��(�|r������F��u���96�!��d(��{���L�p;�uW|ǁ��2p-L����4��{W�N��o{`3.tu�<��p<|�EV�ի4}����}�R&zޫ�P��Z\�a��T�~��1�:�����t�� ����9ո��c���]r����2��1�@{����7Y�dg.:��|�C�����>V~�h,Yb��=�'J�{[�r���ژ9�3�q �&v����X~����}o�a�:�c���||H>8j�����sG��՛5>N]c���gw\��#� wbr�/B��5���bB)������&������ڭ�6�jpH�m����` �}��\ϛ��~|ߏ]_�7�N�п��yZ�e�j̮>���0Jw��3�W��%�c[q�&�Q&�v���L��)�F����~�Ja�Q��˹��U�e|��iy:��}����\�$S�b#��řG��w�R8�|lT�h�?�%��lOyӽ�{��篻��V�����r6�s>J˓�i�k��֝���������� o�;�B�C0�5(��=�z���.�T��M���m>[�����^����3���n`sl��*�kܠV(������ԛ��gݝͭ�eM9`;Ls*���ȸ�V��Ec�(��g��m����;>?l�a�I��l5'l�W=���Z��~�n��K׻ ������v����x�ϕ#=��M�|���j1���ΰ���ϝе���T�okS��2.$^k�t��/;z�t}��h�|cD�+]�	'�;�O>u~J}:���#r$�vr��B�[�����>A|����ϕ��%�M�'�g�5�� �^N2y�깪�X��k�1����^ї[1��&AC�#c���٪<��Q�|����|�����K�y\(A��\����d�H��g'���+s;�9ܗmck�fdڧER{SW5-F�X�:t���wpY��د�����t-
��h�!LF������	�$�n20+�yu�^Y/2u���_~6�m����jm�بX�P���{��~��w4���"@�%M��[�~�0���1�{C�p�����O�yA�,�D[w�)���=^׭e�v�Z}#���f�J�;�"�.�lK;z��Z�mx��Z�c��?��*Ϯ�NZ����*xGR�a>�R8j�a6�GT���-�'0='�K0·/Ou��t�eJ�"�>�������Ѻ�<M��%�r��w��?���`e_.�e|���zËg[l����[v壆��iwO�.09��˃��Q�A�bx��;��M�|��-�=u���y5�r�I�f�:��������?�1���YW�.3�f��B�wD�+:���염�S:~�i8:��<G7���rW'�K���<=�6�LhsO�%Y��T�dQ�B�8����U\��O�lc
��-���O�A����I>��IDx�S�����I��.GA�Q�;����ldWwJ`Y��>G�Ű���t jo~��)Mͥ��՘�����\�6��'�k�-l���Q|�7H-#93�x;^�dNn���N�_{�|�}�|�e����Y���B���FK�$�t��4�����O�}���X��--�=
q���U��P��|OA��V����;q"b�E�r^r����x�"�anْ�:������gu��:�7s�es���W���.���j��b��`-��j��Q$@ݼE���W�q�7S�xc�dM?c�p9�]'�~n�q<;�[;�r�8�f����/��V���Z9��_O:�����s��Jz��򩁙��[�)��o]{��=N��p��4����vd�}��}o��Eu<k�c��:˝{�H�5�)�C�zoM������[��Ֆ�����AX�S�J/�������	8�S[�oI�2s�/I�z�jf}��i����	.����!�/{�4?c��x&
�K�]�Ze�E�$�m|ڇ�?xtGz�$��������}�&�{'aX跧7��� �0.]����㹗����3za�
,�P�~�$`qg���C�G�(;��[�����5a�������c`p�[W4Tu����#�3/I���RB ,��s��z<�x�N$V�'z�H�ml<1�fVH[KX�=״Q<5�_�*I�0����Wj���m\����@VA"�e1"l����LZ�{Y�^A�}ᰅ���4��j��|���\��L<��m�>��W�(k����SV'�v�ֶ�yU:rY���Q��_*���I��:��;�H�ǇD?uE%�E��Ү�R��fͅ���0zV��"J>݈�lO�8���m�,�w���F����!�fvq�|�[�31�*�=���}��7ru��є�kSs��p
�y��K���R���-��P[���'�y�ν��>^���}�����C�۳�NھP���>ǖΤ]�ݘ
��F����d�;ke���Ǆ����Kߞ�K� ʇTt�8�\��;j��va����{�K�l��WW4��/�oVv����=5�!A��h	o��@�~�w����������*#Y���V���=�/�\���a�Üw���&�u�A1M��1����Mu��^E6h��fTGeu-%��[�FT���|W�%��!\���0�[t%"M�8�/��-�����<�!�)��+x�̾�ۇo��Sø����縂��|{����QR����>K��D�L[����5����������'>Vzf�I��gO���] C��{�e@ֹ�"��8D�}l/� {iQ9�Q��:�����{�.����ε��T�0O�h���.᳞�w8�9Ws&�-�$�4a�a�תF�}��tbQ�'}cݱ�;�*VI� E�y�/��t��q��M�㵺�������=w�<�^�٪t�y�lD��Y2��E�-��
TV����&�Z�҇�����|d�npAU���E�:7�Y�������v�6�M˥��@ۨR#D��K��{�y%ݙǀ���7��Ӫ�t�`����3��{�Va��-
��V�n��ҏ�H�ou'ջ/�?�899����m�څ�cm�[m���i�g��{z]��,?k�<��	�wfh�H��Y��i|ހ�^�n��\�L�ͻ�~̡�8TL���+�H<�	R��&f+�+6pZ�&g+��,_(��hD�^hH��g�YZ� �H �U�9{_�?�O�7k���ݵ ��|��������[��(���1L�FoU�����&�r�*�����L"\t׫���88I�����x������K^�x��[ç�P�3��	�Y�'�o�W�udPZ��h������[�����.���6��֞b�8@�	JK��X�k�i�WܝD?���#⻺Eo�l�=k�?=���r�u8uJI�Χ~!��y/^댹����^͌�X��:Q��m�i�=�-�M�7���<³�Ƣ{$�L6;1U��������,�k�n�5�z44񀀐*y�<��](t���m����'�[�4��q͡���6�`�A�U4�Ty��|�l!i�X~���/�wڻ��坶=�'�*� ��ޢ����_t&U�<�@`(s�h;�Z���)%�(x��?�=[��V���(L����"�ݐޤ�L�:V9�s���|J�ߡz2B�D�׺Ɨ���ؕݧ�mܙ`uEPD��\�$A!��Cq"���' �U��d�3�v�m�� ��Zq�W1� #�/���ںbÕ}NO;�ږ�L�{Z5duw�\�i�%�JeAa�J���@�D	�QQ$�(șJ�Ϡ^<~���l�m�[m��C<�89h]�(w��z��u�&0��b��8w�co�q�U�ї�,�n���c`T��q��ϧxM���l<d��j���#�<���2&��R�T�'t���t�}L���9]υVŰ�p��:E�e����'qc���O��Ιٛ-�WE7Ttכ5�9֥>�z���w!�c�3C߿����$��B���D~}��A!6��R��Ӛ�D~Y-�m���:W!���f���a¸lk�[��ҽø�uW6�E�~�s�?p���*_�8~�No�ƣI�{�d#��y�o��_V��=���q�P��C5���2⏦�����������E��ə�}�w���G=�lu��xg����"{j���r�o�!��G�k�R�8Y@U�����tG.|��X-^�Ӟ{��~,����e����C`��2F�=�Z{�=�$�w1O�ÊŭOZN�t8l)��>����Ϻ#��tǬr&w'G�wj���S�)�s��*/��mU�oX���p>|,8E����beO�4(�M��a�n/ܢ[��ؙ�I�[�%��>�`W�J�i�ot�^s�0����p�f��{�S3��O^�}Nq�2�[S媥[��FvCy�t�Idf�ɇ��Wu���;��TZȝ��^�m����;����l9�N|6�]�{���Ӝ9��@��?M�[m�#p�����iq"0���������߇�Go����Y^Tm+��|C\���
�������$�|wR�|��߳�)�	S�����͍��"@9��21|��vG�B�@h/��HK"V3��-z5�.WR����.;�g��:b�^}bz�Ԕbz|�<�k�N�s�f:���O%	ynu9���ޠǼ�BzO͖�=%�{�O��riJ<Z���\�,n^�C< ~�os?^~C��~��"��5���p��G�JR׉��/����;�`@�4ȭ���ά$�z����Z�=	���%�C���v{}�,-R���{s�C�98�������ޏ�#Ģ	�k� L�M��H1� �]!�<	�V��}�Qt�A]O�'^1�o����[�t/��]�6-9�=��:g˶�;ZH��kYA��>Dhbqu�~/���C��͟#�i���a�6D��";�ڔ������=��&U�-(��.m�kt�{�d����ʎr<����#u�> L3sJMq"^�zgU�&�jp|'��kh~ԉK3��/��Zmk�n6s;���3_Ugr�p51���7�C�y31׺���[��fwW&���������X����W:��]�ڧ�;��K
ٝss���j*�x%��8�w��WW�����ԟ�����mm��m�Զ�lT."XW׿^o�����w���&����>^@��"&�y=���o�ȍi��]�'���M��o��>��f�{��O�<xĔ�Vs� ��)KW���M�`�w�PjH�b0]��hІA�nT�+3n��p�ΞBzw��� A�a�R�Wƻ�DPv�ޫ�^�ji VA��lǋ$��n��sO�s��Ƨ��w����u���@��<�i�+'����l̓� �g���,���m{{���P�$�(B��7xOG1�2'��L)����Qp�N��M��R.�;��+x��Oy�Q�����;<��rļz�f�����a�GO|��H��E�e��0@�ӻ?|��m4�o{x�������ؿ4�=<�5�n �Es�rT����	���s5u��~��~)aɉRm�~p(4{�&�P���<{v)�\��ӝ���
0�Dw��j�j��D��[;0k��/�A�|{��{O�E=Ŧ�,�����+���X���An��ô��<�C��W#�G�b��C�U���=���o�?��:%�ޒ��t|���y�v��6�� w׉8vZηu
[ ����ӛZOI���R��������R�PԈ|�|��� �@h�[���{�w5�����د��k�Wg�.�=��hj�%>={X%Ƙ3�+�/�ɧ�s�y�ez{~ͣm�ڥ��b�m�\!��~��_��熏[O���y��+��A{miI�����g�k�-!����1��vҭe����{<�Y�w(����	w337�Y��9\�ML�&/��A�3?�R�D.��'��j�{_{ߖ�)p�K<(������;������ĨNf��q�*�#2i�`'xo/&�V�]�9�c8/����ڵ�/����6J���:{�!������0̋�0 �·��YD����VU-<)�_�˼`0l�)Y;?z�xU(�Ypn����U���p�ᕸz#V�;p�m���&��{�Z<��S����Z"�TlѱKގ3Ums8�z4c��g9V����3
F|d\m�51q���a��ƞ����%�,�/yY�����<5��=�̯V^��o���ւљ�D�:�F�b�ϸ@ƿ`趌�g��aS�ַ��-i�~�����hbLힴ�@P�W�ۂ|����vyĠ��0��*3l�`ٽ�~�[9{�z�J��s�m��L�� �)�Ȇ��E U=���j��w9���k x1���e)�a�s�����:�U�L�k�Uˎ��$�TK܅�ƙ#���%�2W�xm�΁�d�v�u�\��8�m@Q8�{�z�=}�Yq�f�H�]�\٫P�׋��
4��,b6C��9΃��h_b��:ꚭ-���,�w]sJ��1�|z!%�؛�<�ùƷE��[��9��9���[�+�Q�)�-5�Q�=�i&�@�0�yY,�*��q�5y��T�t��w�p��8�c���7e����}�DC���^v>�e��#���Oʃ������J���w\�""�mq��do��>z�����B��𴮔~����駗	�Ή$�����R��Du�GA�!M�s!=��Cۆs&���v4u�2��i_q㗶�6i+ݔ�5��k$2��*�����Ot�ңOzH����Xɦ�����f�Ô�x���V�6c.]�Z�+2)�WPUu��Du04�:���gf��b��f���2��nM,��j�dꢛ�1fL��ȝ��*�����;J����P_��{[���3�V�C�+�8�W���}�{�g\�6C�3pjfS�y���vQ��%ҽ�W�/��A��z����HJ�{��t��虴G<��Z�$2���+�Gw+���\�y!W�֪42��ՍC�y�PL�Po-��0H�X�I���T�;��m5Y�T��ڰ�#����E!M���U�`u�\(�r�Ғ:뱑�n��sU�^,jk�O�1�Y�@�U�j���̗Sz9�Z��
�V���Ů�c��pͅmԏ8ͣsedJֵb�ͮ����o�	�c�����5�xΌ"]�N�S�Z����ci."��9QǷ5�΄Ӎ�0�#�����Y���{o���s(�/�Tֽ�݅���smqm�Ǯ�u�ʠʾC(]�x��<�;!SAޫ�Q� �f��%ͫU� � ㋯1��uŇb���fU�ʻ�&  y�������]$2����u��Z+7*Q"���(�n\Ѳ�l3A�Է��|��O<�ݱsF��X셗ӡ���3�.t�q�<t�r]�A�'
�sE>ō	f�ɰwegsj*R����n�_gw,��iwc��wj�F��Y���ĝ3�\W�s��L[j�I�.���\���lu}X%k��T8(��_�����_N�z��ry�m���V
t����0[b�Ï�����2���U�m����	�r��D:�Tx��9����T�9�r�Q5��oq�f��=�T5���&_,�/��m���܌Syh�3ja�G�t�/�3%��qdm�yA�-�k2��YU����{ڲ��#ZJ����bp�%^�Vs��*�v^���l�:�*v2��������|�9YBI��f��:�V�we��7��db�ڋ/��³�s��U|���jfɛ�WN51�'�L�����E8�2t�*���+vT��^��4p�Wz���]�ΩSX]\TFW*�(�,��\�s8K��T�f�4��)�6���#k�F�ƥ�&А�kx�s�����=�q�TL��o!T貶p�2�H*n7�[�8�ғ��X��ȂD8|�3Ɓ<��P�<]a�I���R0�QD�! ��Ra�NT�J	BBe5
s�H�Ad�c�q���I�
M�g��$I�$ё�AȧA8��"����0��ae�Q��	�dv���J�L �Nr\R���Q�2TH�(��i�[�ʈ*�JNSu)�͟/|���mkl\��u���YF�t$�w H$�'�m��{||uק]u�]u�������׿$d=����"K�v���)�h)T%�U�8�n6뮺�N��N���ק�>��y$}�C�S��ȜO:���I������		$aMǍ���u�]x뮴뮼x����������!$q��S�w�\����(�H��1�_[m�\u��]x뮺ۮ�x�������=@��9��D�a�8���?U�]��q6�g N�9������I�)Ht���͵�Y�_�b%�IԊQ�qȑ�_N�$�"C���8#�"�:S���Ґ��hIt��v�kĨ�;�ŉNr�@����pq����VIwu��rW_޶�;))Clge�]��n,�m�D]�a"���%o����m��d-��5b0�fq\��ۇo/�妻����d3�-S�]����(b˕���Ɉ�z�X���% �t��z�a\K4�m�B�䐮���R@�Z��H����}����cm�ؖ�m��ߣ�ކ���f�I㻕i;2'�"!��g����[G:NT�MZ}�)����m�c��m�3Gq1۷OxlV[��h�n���|;�(+��t�|ť�0��\_b\ۗ��߈�q�?<�}�O2�A�X���SZ���6��ׁ�)�|�a.h"�lx����ګ)z����%Vю��T�B��r��	�oO;�<��lo^��O���MI(�VWe�_j4禽:�5bR*��Q�X��=�7_�d������ G>�6G.=�Ӎ�Z�n��b�����~��d�dK��$n��{�� 2��lq`l�~���n�T�ea��'��q���;�u=)29j�s��˖�vj~�>~Ͼ���wBly�����UO\>M���r�Tp�k��������5ӞU��Ȯ�V���S��c�[$��g��zc)��^�퓉D�/P?W�����asT�,Zi1෼Bо\�I>��q>b��`�]�ʌuw4��x�cn�1�q3�P]�%����mԥ���¿�]qL����|`�����C��T�\���@�;�yǳr��9N3j,�Kl�G�u���aBsb���<�k_b�hT�\\���"��]�w�p_op�gZa��%�wsU+�"0��OS�΄��΀;��^h��V�̳����x�������m�H�m�c$D�9�9�~|�{e�G�8��>ܒ�F���j�aX�Z)�Y�� ϝ��M�w�ToQ��Z7����+�\���/M,�@�y���:b�&�-9@��cMjz׶}�Y�]6�MO$�w������^�"�o����׹=��B�9(2jbS���ao���p=�n�λ\�+��}�S뉧�N���������T������Aŧ�W�=�E�磏:��|w�([>��{gN���<���Q�C�c�r���޻}�S]8����z��bz=���z;�O�:�H�z��1�萤cH���7o]�u,��s$�]g~�>v��!����_ �zH�N�s�~s	��t�����y��p����ѾM0�7(�#���T�L<����I�(�t���O���a$�=�xqJ^]�n�8���Z�N��e����B����z� Kmzԉ��s��n��sɄ υ��?)��������7���VG�?A��<�x��$����ʂ���n�s���qD�e��8�Qt#�� p�[S'~^����{;�C-^K*��v���n3P�/
�<5��˥��].�*�<�lj��>q&3�h��)[u�pl�]���x$n��0S�b�>X���]�k���N��.�{d�~�m���[m���~yƣ����ە#]0��1�����!Ψ/��WȺo��G�����o�q��~J7 �OmlaXy5S�����n/����CuO��}C��~(���ƈ�*��m�٨����\w��@j�٦�D�I�)3��b�,yg����s�Ⱦ��[�+��u�����&&}�.���b��P��֤�|�	c�婖���
]��!F> ��gǟ����;{�;G.1�|,����������r<���>ܘJ �xpc��`�5s��O��������OM����t+"·g�W-�Ne�|�-���h^�J��f�q�ở����.ma<�nY�4B:�V�JA����Wj�V��GFN6�z9���{P��u\�u��0zCp� �脠C`*�Р���Mz�������1V���j�P��Fox�Tݝ�'��Sn��} �^�OW��^ܘhws�I��)	����L�NޱФo+��4���z=9�P1�[�&��k�{�j�>����X}�a<�;/�ٛ�ʿnK��߾�\ڬ+���M�8c㳶���$�lvs�fm��-/%,=������ {1�#fN��!�X�.�6���:���fK�4+���$ P.�2{���2%�����:� ��s��y\{�o!��#��m��v�m���[c��*��\�s�8����� ρ��ٍ��rC�,1�\�4w:�Nb�ꀩ�/WZ��xa���tcULs�F��i	���u�*SM�-z&)���09����V�n����N�`�n���+�yE���vcY~ZLkǳ�A6��0��8�|�Ѱ(�-�����5��1�_���W���'�������v#��@M��K�~�2�4Tgwflq��դ���~�,8ے�V:�X&��-.�8`��o�XPp���`�~�6r�����n�>�'eu�z{�В���zD��yD����A78���O��ɞ�w�e3�_hΦ����nEI`Z@����V���4�%@��`IffQ~���+���*nl��̭Z����
aA|E&����˼�6�}<D�\��W��eG�j jnUl%CM̻�9C,xes�\TZZU����
�H������
m�<n@6�.
�4�페�F�w~�:��N��/4	��X����Go�2�P�4r<��9��me!0�`��f�"v/t��Y93��&[�۽X�ў�ڜ�@��%=�wbs0f�Ln+��L�Bjd�,��
��$�o��<Qq �L��(��t��M�5G���kPњ݋�{�SX�ӻ*]Lz�b1�.��E@jDzU�ζU9j&��ي��8묡[ �"B
LT�q�4ԍ�qJ2�ʏ%co�rG�鴶�n�m��m�D�G-����]��҅��%�����O������p���"�m�z���_
�ߍ+K��� �ʛ~�*����������i�CV��L��@��^ل\ug��eP�w��AZw*����D�Q�;���f�q孎����B_����j�hR{���y�t)���E��76���c���
���: ,XC[�'z|�S@����DkM�Juk�o�sGuH���k-��5�+�;�쾚|jg��K�t����:/���%�Nߵi�l7��D��s���S������[gk�U�b��˦�c�Z_�Z�ڃ��_+��d��h���[��^Xp�<޾�~�{6���=��x���k���
�;�dp�͐�>���䕎.�`�ٜUڋp��$��O�	E��t�oO:��x�u���ḻ��沾�|(��R��7�f�0O5n�)�B$�hP�Ο:cX�,��OQ���5�k���_cg���v�S+�Ǽ '��o웝ۦ�o�ݳ�No��%�ȖS��/u�Ws�	=��8�T��u�l�\�G�"��w�o�TY��T�/4�����sEMoY�\(Y�ۣTG�@�)���N�pWg��_Yc}�2t�V1����r�u�}���ZjQ�m�6G�uϣ���D�gB)d���\��~MﭮA����m�۶�l�)�q��iq=,#�3���G;ȇm~hD�Z����xw~I�W}����c�!Gs�S<�<�Zy��=!�&a�ξz>AO��� �Nj�D~Y-�m�dB�Z�9��Qe,=�`0�y��: i�h5�)�Q'�TC��� .|������Fer�}��̮�U��b2�ݚ<%��ro��Pcw̝6.�k��
c���⦤&)���2�<=��m�͞��MZ�/E�,d�0��"'� \;�֯1�����,�w��_5LLΨV��W�}���Ǝ�����G�=����M'�k�D��!�LS��Pz�^�wos6ە#RWB%�?R�ߧ���CJh$�lb�E/�^��){�s�,`��%�ǂ�%^�� ��ܒ�Y��P�Zgd�`��gA�$�r`�����{��5�Z�&>�\�\"�	 �w�>�x�|ع��4���8/�ҧ|̘�^�4v�ɫ��W=��k�D|jퟞ��z"�=A@�t���/!��R�yt���%Kq}b^��q4]b�����L�p4n0-��|@1�,���
���ߘ�Ov�G^���taR�R�����=��v�St�S/.�[=�T���0ޥC�P�-T�H�<l^(\�;�YI����Щ��(���vCڱ�K}�����p�!�޷�V���}>����~��=?�вt�9�۞��=Í��zn����)y�����pZҍǥ�G�L�0�Ey���Nw��7�A�s����Co8r�]���[��1(9���X��A��r1%�s-r/7+J%�>sG��u�W��C��jrk����
�}r7K��\�L���їw��qe�I|5x���g��k�k��H&�P���M��s��w�.��9�k^�ǻ���t�3��'I$��_�\�ʨ2���o8hp����/৔�G���K޻�oR+�WI�:��ۼ'M�L90��m/`r3���iNm�>�5���C�<!
���v��>w�R�07b&�:֣�ＲA��N6�}�`Hq�~ԮZ�^PY4��kC<��г}�J�OY"���
�����1�!����݀��-��'���&���ܠ�eO�G0��[�N�G���`�4������ӫT��4Ќ���x��81�����S���xV,�W\�g[J~/6� $Fb}G���'g!7�b[���ޡ�-vO��(?Y�������}Cv�o7��I�;vb���t.X>1&��
��m���3�+?��ￓ�׾�����B���pb�
>\���pL���J�[�8j���h'8�e�Lmdp\ɜ�9/XFm��lC}֖pzO[무/���^^^^^?���[�{����`o��!�� 6m�P��SH�u ]��'&��q��DPwtn*�͘gu��$ܮң�n���=(A�8Mڒ�gNm���u[���rÞB9�5O��o�Z_�7חڥ�����8v�X?�dݯL�����ez{{(W_���Pn7�^��S�<!7��k/Lh�LI��W��}s����!� ���v׎u�.p:�ף���؍�`N���z1���|ɸ���r�k��)�����}�7��`k=%*������4��1�k�ܲ�t2EA�f�9{�ʬ��}X�K֙�A�`�
xc^=����p�꺒���Ex�۴���e�5緪��+�� 5�YƑ��h�7�k�w��Y��=7Ƴ�J���#y<,�n�kU9�1����-�\�~�L�����a@�Q!�B����Ő�����4N{��uS�i�N��-qT4�����@A����1+@����"��2ѷ1[J���#R�=p<�м��Y�7�JFz�8ۥ�F�Z��`�`L�أ;{_�r�*��gz6�}��q��O������v�� 6��[�2��O�J���PV����0�{}��W|� �EJ���^��v,�3�'�G-�T|��;�u��̴�+�_V	s��ö��(Z�"K���ޮ�Cm���:�c����ܫ��O���18��2bB�QrW(�	�O�4�M4�[m�v�w�2{�����A�D>�gZd�=�=2�G���r�sޙmr�-�Qa*�ԤEƶ�n�-r)�&�mR:T���&X��p��삖Z|��'��P9UO�Л��� D�^	�e��V�oIve�z��+O�����x/���:�j�j|���g�^BwLVV�7pUB������*��n�e������Ѫ���x����+��Sb��˃6ʥ��'��a(����?��::P���w�p��}��lv֖T�,�A���$N��j�|ֳV�ީ޽~8�h>�؆��޵z��O}��P�lc
��oT���L��x�	6�_v�c��~04��c�`��N,�ă�cVM	�~�������U�U	�|�����v'�����)�g��1��� �>l�ȍ`$nħVJ��C�"5��[�`l���Fu�42%�a�?�㿃�ܠ++S���R`@��51��sJ�?����_��$1x~*����MX�<TS�\ŗ�5E��=t�xǘ���#/���/�.P�AC�AmDy�1z��\ם�C휼������l$����u���.?�/i��9p36L�>��Pҟ-d�@BȒ�R�A��a�8Ex�DR=q��zz�<�'�������k�j����!�S��{���+E��Z�tқ�t����;޺��|�:�|���ƚi��~���9�̴g�����9�_�W�Tߑ��]�~� �5;�ׇzh��;�0����융�}�K["U	���#�����!:���r��%���A���g�%u�����#�i���Ba3y���s��3@��e�dkt�u^�`6Ad��*��k�貟9�-%D�������0?Z��ޗΑ2%��8���~�t]=�G�|����VM��;wr�p��\0j�bx��_Dz�(����O=�/����:�`{Z'��WI�����^�osg�[��z~��Cʁ:�
?i�+?���@��L#�J���}�c[Eۏ�n��UTRG*4�^�-���3�>ϻ}=���=��J��#�_���7�5mʕa�9��S�����i��"��ו�c龅�8�r�5�xg�~ig)5� l'���W��Hަv�2�7薻��Gd��@���6�\�*�$:��Ɏ��Ͻ���g�p߱�K��{�
Y�3� ���~�1�/4}Һ�V�6i�`��^[a��-�~{kv���2�y؏	*ڋ�`�hԦе>�C�۫YA�F�*�2�'3ov�&v�� �r�k��mƙ��un*�`�z�MK)$���$��ٹ�����5v�u�j�@B�Ǜ������կ!���ʤU�]ڌ��Ż8�:%\�R�Ҭ��`��,��ۨU�v&W*X��+7��Ն�q�}/อ�����[쒸����5V����3qM�}���m�I�R݋�|�ǒ�uX��q�+�~8""���뭷�\͔�Z���9)i�,�q^���6��TȆˉ������ÆX��,���R��4 ��!�}e.���ZE�;�<t�b9�Uܗ�!��;׋N�ɨ�t�^bͶ4L���5av�oa���7�N����U�wjR)�dfw�p7�R͵�����9���^�Y9ξ9|v,ԡt7/��qO�eNջ';�[]�$��/p-w����m_w�wt�t�K)����d%kz<��VECV�#L�Q�8nĘ�}3_��HӸ�9��:�u�5yAG��T�P�8��x�%؂�6,��-x{:v�)ݻp�����t�ҝ�������sx����xU��,�=7l�����*��4��I�:�� ^/L*ZE�1�6�����1�u�B�^W[j�D�v�'icA��A��ܰ!��y��H�3X���|@�|��(�.��ݲ��
�U�R|��ik%�*�vZw�U��`����*�WK|/Ww���%w'����@���ۜ��*[H]!|��V�ɑ`�ct���}�d}ɾ�V��&�5����	C7Qy܅;�S�=:�^��UY}�q	���S��,����[�Ņ3�M|��wph; \��6�WPjѻ�B�Uī��[�W�:�f�N��k;�v�p��Z�v;����E���y��LV�+hbGvU����U��0\����k`ڰ��$�0m�v�0�h��J�-���=�Q�/{��ytJ2�ٶ��XKjq�V����Wo^N��	n��vLz4yM���(@/t���-{��6׻��{�~�7��2ܝ:�3y3���T!J`=�[m>lvv�qJ���ʶ��>��ˌ���Z�h:����^�RTw+�������n��[vkgu��R����L�V���v�G�J��:5�W�*Rft��:m�i��q�L�|�i��^�*��n������e�W�FSӼ��UV���zY���.7��;����T^�nQZu'_�p��-��m��N�;.���q��q��__]x뮺ۮ�x�������y��FHD�mY��S�R}�����FA�'����ӎ�뮼u�]m�^<x�����ߌ�$�
��t�����9u$�H;(�$O\i�\u�]u㮺�n����׏__�2I�q��QȽ��8��2H���@����x���_u�]u��u�Ǐ�>��I#HA���R��&���;��ۺv^��z���ۈ�;���+�䈉�v�!@ڲ�̐��TG{h�::�'\��uynu�t�K�W�򹽻:S��8��P�ĝ��絧ͷ��.<�.��ʼ�l�	�ܖ����'+Dټ��"�:ͷ]�9J�������!��&-���X���p;�B��Q̝���/26�����3�[oo��h�7yߕ~p�ަ��֚i��i���s=��V�wfz�S��r`K���`s�>�>�U�a�q��_���y��Y������oo���<��;�k
/v�oV��v��x��,�V	���p�ߺ�Fײ5�+�텕����:w8�&-�{�=o�}�C[���c�ǅ�U���4g'μ�T���]�Ε��Sp±�M�q~1	�w��z}�.�� 󷼺�z�:3����B��.7�����gJ�hM��U�-�Jos~���D�P�����p�!�4z]0SP��S����&*��Eu��L$��_ /4G���Z���b�v�RZ����{�K���_��d6H��k���c;4���=s���|O��g��wN��;e�z�����T÷`>�=�������C	x�UMp��a�����>=/o3.��B�ףD��xc���7�0bjr+(�����(��_{��H'W�$	m��j-y�2�����:�s�r��.4��d�v�/?�����T��(l[�y������]�8���ʄ]8e}�#�tU�4�x��z�x-v����u��NЁ�6��C�!��,_$.ޣ�c��
:Y�?{�we����evwl�N+Ӹ�q�ԧ��s�w�`^�I0�ŋ1��wm*��l�]�c�Vʿ�3�Z���A��l\��K��8�350{��Kos���$\L˽����3�g����Q�oƚi��i��>�����o�����}.��}�|�Ota�7y��$�o���Ԛq�&���� 3����z�ǩ�[��c�����q��;X����ґ>݉/~&�p�#�ok�����6���wzv/y*��VBL�P< ��y_k&, σ���T$���}��0�R �b}=�w����s�,fr9Nf���}h�{��(�:-� �xA�g�,[�E�??s���c����N�5�1،oHa�*����r0�7R��Ƃ����2X~����D���w�1�.$�#�v��%����7���}j�l`�❭@Mu�{՞�v��\�%��u�P�Ằ�8�`�l�ļL�ss�NooU�'���à���_�������~����H�^!�ZsJk������I�~����+>^�#xL-y��B�[[knl3�Juar�i�7eMw8�f1œ�cbZL�;={ZN�aty��������"q��6-t��F���F��'��U���3{��*�5�;�EnPÓßb����n����(W>;3�iԫ��ߗ5ʝ3�G�+������Ȼm�߆k��ܮq#���8Q�Ǻ�1�^nҕn*Q!�v��od��îY��l̘P띱a��L�I�2�z��`�a�*"�ݺ�iPH20x�.����F���U�\�<�c�)=��zYZ��j��i���7��]1�g�1�h��B�@x�	5'
\)(�IL���E��є�ID��jaA�3�qyyyyyyyyzS��w�����gO��^�"�st�To����x�;���6�a���S��t�]7އ�lϵ���ub�xd�r<�p�\���W=�Be\��R"s��c��"Gxa����r�_S?Z�n��u�Z�4�; ��O�TJ����s�����3��L�, �sya>�B�8i�������\k�s��?XR�ûȆ�-�d����=���=2�Tzt}k�{b�uF��[�����ʮ&��y��;�=�k�������3dz�]ؽ�>mПg O`������Tu�j�`�)�۾չ]�h|`3p��D��댟|������x��0��O�К.q�qV�O3o�G�#�q���ޘP.E�)�0/���E_*"�����.�Ԝm��ś���c<oÔi�����J���r�%s> �'��Z8�����-���r~��*�G� H������P�����<�|=��[�A��smtQ�si�],��􃾫N�N��s��&@�n��Z:���nϭ2=ǽH�W���u�l�ⰶ=��ׄ;Q.�}��2��f<:{T3��o�hݫދ���&�᥼}��ض�\���]P�;��]pڃw[�����4�q�����8Ɛ5�^�{v�N��k[�n�wTX[���.����{����.1�э'�J��^Xpq�8^�`>�/?�������?�xӻ:{���hwƺS>�)??{��P�ߠ���G2�R'��IeX&#�zUu�ՙ^�8�긙���	|����A{ŕUǫ��=�Y���xN��hinQ�}onC�g�s�p�?U���KH�J�	ЉX��@[C�b�NA�$^�l��1���= �'�\V��e�c��ֿr�n�����[>Mz���
�އ}�]��T7G�u��\ �'����L1TXB�.'�m�weC�����3>�7q�yaV���[Ӆ7��@��������ъ%;��Jo��s�L3�;�w0q->�d9�q��Ҝ��<�N������4����TzGM����ղ����]�	z�dts�4��޽����f0����
�..�r��J�r��ꭶvj���/zx��� �����t�T�L�;	��kOv���m��ް�.��n����DU����?��RI�����3F�3�
T��oO���8�}��j�F�5�WBx:絣Q�� ��D��;�|aϾ�`�\��N��ʒ�z�B�~�Z+tQ۸>jF�=Ku�V#|֣!T���q��7�@�E/#������xq7��r��^��4��\�=�A-�{��x�����o5NO+��{����=XF�Wa]���)˷�s�u��K�������������)�	B��+��A�������#��ݜ�7�i�5i����)��C�B�8���<����S����'O]�.�n0r��K��j��Ǡ��EX��3��Q9`�4d�OG�6����vc3�������i������O`s�>"}���@���<���T�x<!�mfv�8Q�D��3�#ZZ|��p�W�����d��5ߝ�㝾ڶ}��y{eW��(�\I��jd���;S5{��Jp}#ŀ�r��%HOJ�Ja�#��#�.����sg�J�ݮyު��L"��6a��qĺI����� ,<��p������L�-S\i�ǥ�c�a�y���?J�nS�Bj��O��孝�^��z��+�_c�l�3��yxp���}WN�O��ϬCħ������l�q>l܌��9���s
i�5�~����ztp��P3~ާ� �, (�%��r�2+�]%�1.����6���~2s:���}u����S��b]/X)���ֆ&~0n��w�@�o �zF�ߡ�!h��M�fUQ�t�i�Z�Gm�V˻V!��J�a��o�۽��s&�������uidq�+�>��Su֮�`�����,�t��������Uur���⨓-���k{������.W>�������?���6��[�m����%��?�l4Q{�Y|��CH{k��N��r��W��Q���gvJ�2�<)�w��OO<�׊�<�N+�L�p��l,,s�^���sFeC�G@�{g��������0����1�4������MW*�G������`��T�P�u9�I�^N�'N����{�L��2�t�Z����0q�|5�QSuY�V�d���.��k�3_$�&}>Z� $w��AG��͸G���8�gy`�9��V��,I��9���JZ�<9��E�_e�%�B������q��q��s���J"r��ݲ�ٰ��U��4��T�=>�O��-5�g���:a����ͽ��׵f�$w=R��{���i�6Z��_c��6��U.�ގ�i�7i�+Դ�-���M�]g)ͱ� U��Ű��~/4�劂�r�e�)��,�r��2 �6f��R��@M]��<�`vD�u|5���Ƭ��{Cj��'!P� �ܻ�Fy%�PݢM�NJ�cR�����T�VU��U�v�H^e�1�/�[NK���|�Cؖ�K��WVdv�)�w%l�g1�)X�8jɡ���		!��	�"�Ԓ��Q�n?i��i��i�޹�UW̹�����[E-h�K0���?q����f�De��l-�UR9�~cV�f5݅�%}7�NK`=�<v3꧶ͩ�n�K�2$	��{�k.�bL^��^ne�d�ҡ�N뾏���F~�gU���I���(��'��%]�]n,y�kOz�<	�;�ex=������|�b/��`h��Q�2��I�h�,��n��}��9�9p�[0��a�@~
��٘m��F���)�[ZIg���^���M.���&q&��9^|���-�Dķos3Y��Y7F4�5����آ�F�XԳzv�^�2��%���qS��gP�&��wt������5�6�Ss���1wRD���é���ڼ��_��b��@��5;�{pQ�s?���y�Z�<y����a/�T=�>F�X���a���i�E�^ȿ&w1��36����Ww�9���ۋHۖ����{1�o~%��ǳw��.V���Q�xs��.U��T�aUbJ�⭫k�z��{�8���üHqb�yv=�X9��*G%B+�'�,vdlm��u{���;�9��w	oO���i��i��swJ°�Ol�$c30��`i��vp8�i�"4�s��h"��D�4p����͡��(�D�^\ͱw�
&�\�_S�f�2w�kժj��veR� 7�P�a@O�VZ@@͹v��ȁq��\Le"M-�{�j��(C�	��JsE�n����=�Ot3x�R�����K�FIb�YŊzql�@g.����'��x���hY�xzV-�[�A5zzY;���Oz���h2PǤ���_Wy������h��Ix�$����fw�� �Zl�aj
I�����2;n�m7M5@-���D���|������Az��_i^��t�m����WJ��s���L7#�S�Dy���+9}s��Մޜ;$���
�+�Le���vA7�6˵�@���嫪���h1���b������y��yG�5�*����c�ɟ�*�l?6MT�&��.''�5O ��Kw�K1��KL���@W��6���@�[�ͽ��\g10t���硐�Ф�H�VS�7��#*�y4��I7'1}�݂-jQB�v"').L�Uy*tюu�gh��ǺNEqH��Zi��i���|��|����'_S데��c����Ί��l����J�p��]T]#��](���dy{Oi0oH���d�\�/b���~��]]���ii�I0���
�f��X��}�E�8\��.dߨ��wT�'���Z�6s{ǀ��U�e-�a��H�����96�0��պ]�/�MID�ɰ*Y�4l+,��p�wG�[{@���L����h@��m��gz��S�j�����=Fi��eL��>�bb gT�>�Q��_��\�fΝ˩Gw�z]hw�`��G�;�:��@[z`��w�k0v@�3T�S}�u�fTT�w
:��H�F�&_��Ȭ��ЭE٨=ĝ��'{M��$��L�l6PS�95�WZڲ)��6��ؖ��1�6��o�8½�/P��Y�@X�������w5�T��b�Ӫ�ע�F�Ŝ|ơ���D��Y���e8:�;�q��7c�⹉\@�4��u��:_V�.OK!%�(PH�gH�2��L>"��uvz{O4jS^ɷ3I����z�9u�,[ې�s��i�[�9�t{]N�n���.�.gKwing�������?����F͗�I�]�P��H�I��+�s ���ڭ曂ͧ��71\��5YZ�Ԩ=�M@+pc�c�;�ww]�\x�z�;�w:<hbS�;�����M�SM��i�O�Pa�*�����oR��X�[� 6��l�3��h���z07�ɫ����~y���\�����u�0)gH�=���Z���|=׻ت6�ӈe�2�g�!���.�~D=����>��"���w�y��ȫO�O�I�崓�nɷ����C��c�0}+�)�Ϫ|^�{U8�=���_�,���WJ��������3^7��W��MM�?OU�n�6��nR�N�x�ܴ��"j������5��q��a�-������Yy�/���07s�+�5�@Z���8g�Ȕ���<�o�f�2�M�%����5�I��3�9�=�ՃWT{p27BHxR�w��6������؋[�QJjͪy9.�Z��<�T�erѓ%0��t����6P
�P��S{��E��-��f�D�Ū����;y�p�S��BN}�A`ų��/G-/���چ�7:��:�Q� ��@_n��=r �0�v�*��K ��ܽ�YיU��m�w�ʨ0L��1e��P^nmp�c��ms�J=̾�hˍ�	E�SgV�VsUK��Y��E��ݎj(f!ڶq�>�˅�ڷ|;��.��ѡ1"u�\�
���Ф�b�[�Pw�k��K�o�ev��%��}��$Тo�bΔ����b��4xv�]�E��a��v�0��bL]N(/�ю��PP}�ڎ����ŕ��R9��^*�1Ւ&��9��wPХ,�'�T���z�o)�b��ь9{���Zz��8S�JIK�0,��4]�k��9��|�mm�(4c���E�}���;b�����j}�b��:�j�N��8�r�Ƞf����˰���3&ښ��y�!�;��n��Mqv�|��f"������u�tk��C���.�V(���ko��Kv�P������(����U�*��`�(�	�Ԡơ��%V���������<���qc-�f�n���*�A\1�)2��.H	�\p.fع]�������$�TR�|�2�݊��%�lˁVjA.�`��H�_]��O;t��,HՄc�*[p�p�Mۣġ����h��ʼ��e�]'v�����|s���vwh���Ъ0܇��6_x��!z&�wbک�S�s��H����&�LŴ��ʜ�	�|8��Wtg:�fn�}س�^ʸ��YU�DwҪy�Rv;�:f\DIhK���c�ȝ���ʭ�aoXkWm��8b��6jX+ۮ˷ee`�����;\�n��D��ǂҙ���]ދ�|��%y�K2c�X�]���MEpP��n�����W#�ބ���%:4 T�O�&�T2�܎���/C{�}W�i}ƒF	�B5��?e���e�w]R�O�vd�E�}����-l�GM�en����Q�7b�@Ri�q�݇�f��I�݂����p_R�:�����U�]N���۠2Kڙ�e>�#�pf�[�5�f��)Q�X��;r8	��5�u�*�����$�G\�B�L�D�69�o*�w�⯄���;&-��,����t��(g)�us��Wm|��ѻR���Z]�X="3(a�z��ۻ2����G��g"ٺ�����Z�/1\'d���=k+(��w��&Wד�r]L��z_iS4�ŭ�PH���e"!��q&�E>HӔA�)$I�L�[+���|f ȋM8�m��d�D��@��M��
&`BB�\Epƛ	��q4�(�#���QB�A��T�<aCP�@��A4����H����Z�6
�D\�2�&7X!�\��%�\+9�ZuHG�q�w{iD�eQ5�6���Ƿ]u�]u�\u�Ǐ����׿aD$�UPԬ�ݽ뻶K����u�P�I%QQ���}}u㯎�㮺�:��Ǐ�__! 2&�$jHpR~>:�9�ݙ�/��[o_^:뮸뮺뎼x��������g�O��0��ב^D	�]�f�ɝ��W�[M������뭺뮺�<x�������?&�,ÈB��W����Å�u�w^B%�J���k���FwiGE��y�x�֛Gm�����w�R~v����vu�LADA�m�9��������H��ʶݗXu���y9q^�;8�k����\gVm����m�X�Y��gPQ�g_��eڴ�;��E,�N��t��;���D�������y��yݐa��{(�,�����R'A������(p�K���x������t�K۴&���c��k�kݧĵU�v�˪�pt^����A�� �Q�
m�H��R&Đ�$%(#I���/&8��M4�M4�O�Ծ�U��ι���l��dB�RkB��������zλk�� �#�[IM3��t�e����f)�#���co+b�$hi��(Z��SR�i"7v*�D�N��8����m�W�W�"�z��o��,�vs�g�h�������S���_��]zǛV�w��S��c������fSZ��_�q����Y�!�z@��kz�^�"�}���l����j�T�J�+א+N��G/_1������O�H�n�l���R����}z������I�ÒO��Y_��u0c힩��9~�[c�����"��R�ț�\�z����Z�Cmmz��N��Ϥ�!z;���]��4�q�I�E��H��0c�������7}܆wR�u�zAe{�_���ƨ]v�CtuD��񵱨����A4��s���I�$�?M��K��uH{�?o+�
h���V�U�A|ug���H4]�G8�M��{="5��P�F*yvՊ�x�ޟ}��8]pw�F*�K��[q��y��ֵ*(w�oSU�p�z%��Vk��x-�n��8�%��A������G�������J�=�ًC��s��-�|�|OioR��ݛ!^ǌ��`���}�=:ipo7��`��>��E�sa�nt��<���\v��fk5Q���l�'n�f���5�0]�M��$�V�}�:��۞7����g5�i0�d 7�[��0qã��S�� .�A��*nom��E�e��Q9�^���GX�u�������ў�k��ʞ:�A��L���Ҝ��X\�T�33Ff��3���}�+�����~7��G�e,_��y��H�;Fn �}dOj}ϧ�gREEe-y{�͡��Ov��D�o�!�SUo;��ú}�]h*:�-�9��Ĩ����Y�}爫��� U�k�ǒ��a�N�"Uk���\3�x[ʒ�Y�4׎o��w�1{�3O�+�u�ۣ}W�0V���Av��MYɯ/�vW�ziX�R/�d�΀�4���K���Ls+2����QGۦ���*K�����uɘ�j��M��R$��k����]�5|ԥ�_Z�ZbDC7v�z���y煴�4�M4�M4���]R'V戌}�a�I�?�dW�iߞi�@/<ÀYQ���Ʈ	�}7���{�����J�O$�{��,�WN���S|���)'ooQ=��>�N�v��w���n�]�eOq�$�2ɢ��s���Շzٽ�S ���۰9�	��"g���03�l1�n׸hMn�b��͖ܽ'rSL�D`�"~������3�Q?{;7���&��Md�d�+v�֭3�}^�M�s}�'vwg>�z}��xQ�� ������o��J�7��p�&w�j2eI��]����4�\_=�y��bi0fvf'�O#��9�*6�zR� �l��}�����[Y�j�Y0o�V�f\S{+���B�$�}ӟu���,5շ��5�l�����ҟ_�m��4b2	�攃�\N�D��[�BɾQw2�l8�����z������
����ۙK�� ����@+��;������틤�6)�5��Xɝ/X��=��\��}��wd���X��KĤ��*��ri��G�c���7'��	�bw���?�������~V�q+q2��2�G� "�ޑ������笅��
#/�ÍH>y�ľ�j�� T��x�ca�}M�����!C��7�b#�qXnU�G�>S5N�Ǚ�1�q�����z�8=�J��3����>�i����`ܳ�W'���,ht���37{��{�X�\�,$ڠ�#�0qԃT;ЎU8�;a��]V����ӫ®�v�'�U�E�3�����=���Z�+2�b�6�Wa�X%'[F]�;y���lӝ)ݙ����U����n}�����-�E�yC:r9�"}7����xCろ��U5�s�;U:U�#���=Ր���-��:�p4dwz}=Q;OW��]2�/*	�~F��3;i�E���La���>���{_JcS��f�����T%*�^Y�݅�^%�4wC1�\hS?�NN���t�1�����I���n0r��0����,�Q�r�4�ˮ�gMl�����R��ˊH��غN��8]CW�
=EB�V�W��a��S1j���\�H���s:C�^5��aV�y�WO����\�P���L��Voe��eKL�y��ݫy�V�]�v�(�@\%�Y�e8HE4Q&DD�'N:���^^^^^^^^^i˧@��.���%���!̻C�F˥ޫ�n������]
�6Z����e��e��9ĝ5����%0@1FKg^�O��G�A
v<	��ku�&j��^���#��x��!&�����p���IY�,RSy/f�lݔw*�H�4QE%C��Pj}X��9�ϻ �_y� ������{2�<�lÓgm��{�P��c��[/��0N����S"r�,�|J;��1�k�����u'2R�oͽ��g�[��pK�\3�R��"j�8Y����3Xw��yw��Q����
�-+)kyT^�8�R���J`�ݜ�X0�%\��8ӎ37�3N��v��sN}��:����1Ȼ}�&f��l�Ba���3Y�34*]�*l��0Q�NJ�u���]�|NeE,�y��3�@����"���'`�{�Zf�Z��3�%(r^�^5,}�h���^�Z^�k�tE�͂h�cČgkF�j��9.	��̬�b�s��<�
49&��uw�[K\I:�,v���F�s��{��M��ﾰǧ�M4�M4�OU�K�Ef�^ރ�G���䍦0���=k�du�[{XG��������f�k�y�N�̦��v����̆�~>�X�������}��0&Q��U����o�e!���V��ϕ��}ÍQSr�VF'�5\T-�H���t���[�����L�M���ȗɷ��eNVVVI�4��R��6
X7�zS��'5PX�wl�n4�W^��܉`�aR�m�ZI�|�ƽ��s��l-����	i@ʹ��ꎇ�x*����Le%1/��.y�qW��y
4�:��u_`��P��I�[W�4�U7�"֞�ϧƁ���C�q��ǯ2�lH��ܽ��Υ��CMߺ����W ������1�߆��]�u�*��ɲh�:k�Ж�lgo3>g����i*J�k_g��%�{k�����V���h�y¥�t�J������U��*N�����FN�౗r�UhD�"�z-���2�:�nz�z-ҋ����>T�.=`6M>2	��T7]�{�ݣ��M���h��O&�f���oS�W��u�p�O�n����}q���%�:�U���i��i��i�O3�wϟ:��>ƞp#Ζ�z@h��"��}�:/5�B�̠`i��*��)�ĳd�g�[x���'j��V%�ze��	�l�b^����c77������ܯe5ǶY����l�b٦� �+�Xq�c-'�vm�1=7���l�%���ji�
o�������WY4�;�ٔ�=�R�0`<8xh�W���݌%����L����tI��H��ޟ^��v��ܼ���z����CkzP��>���&�p���3��d�FU��X7����6=;��):t�v�!k���%khx�M3�k;��X��=��� Q��M���-;�so�[٧7�N#�؅tߗ3�p��`Dw]>��"��dl��ʛ3����U��[��!�V�̵or�+{7�g���\G?���mk��*�k�I�ٓ��wqx���aJ�$���&�M�W�i!�64�HغӔ�,(8D<|(jd��e-����e��y9H׮��*�}���je�S�u1��fvKnaVX�`4wF��\�nC�t�?���l�r���z=��������?���l�Z��[Z�����f�f��F���31�m|k߼�Ɉ�|96\���N�q[�k>ǲ���;��}q�z�G��������eS&�c��5f%��;�>��V���
���ek�H�>9��<d=�6i�fWuz��ça�+��87WP��������!�Մ{$$:���N�b�+e�K2�p�j��
����y�Uo���C/D��qF�xU^ff�s�|��*���`�����B:W9���c�����5n�CT��m����Dy)�H�r)_��]��PWێ᝔���,K��35z�/8��K��9����{s�|�q���­�nK��m,骽�j�uy��o��3x�;D�D#~�;�6����E��yA'V,�� ����O�zhq4V��H����
���h�g��Oe�r�a�s.��9�;ܯ����R�V#��^L
B��Ͼ�wk9�A�A��A7r4,�K5���u�r�NN�Uq����)*���0Ue޼ެ��ͳ�r��}]x��sOI{�wD;�� S�L�)�EA�(��J�DUT�����i��i��z���=���~��i�!H~��}��Z�����!���?q�6;���5'�����֚�ờ!"��W��wf�l���S]M��sgݳ8V��XAT����$k��-��lX��zޭ�g�.5�=�؊�wf ��nr��{ʼ6HM�|���v�5V���['T�*"��'�^�;����w����� dk
{�e���)ߢuwen�nS�����N����^��a�ȍ������ʂNM@S�g+���vE�$צ���paS��wnn���P-s{Kd�+a�X�����V�lj��Z] �y��>r�?����Z|}��v��+�wR���$��u��M��C]6��}����W�X��l���~�^�x]��/l9'���qb��\]굄�f���5�:�	C�������`�p�>6���_E[���2h�d���;�L�dCM�SF�#L�[�#s�1��nFv��n'-�����DE*)��N�$ƃ-�AU*��ˈ�	� ��w"�ܭ��a��p���*
��%\�O]wD����=����ޭ�Y(?��//////?����K3uWofμt}��]z�@�v
�ў��>��oy�c!�!J��	�*ȧp�+�[Q+�
�� N�)in�S&�g�T�b�D�r�3���qC�=z�|���h`&,kxO���Gl�N����K;m^�gl���e*���p�l :P0B*���z���jճπ�j���6��|TBU^|��n���Š?~����i��� ��;���_�H�h�=>�k����Rі�|����r�Lέ��\�K�u��	++���Ƥ	��~���W�z���a�t�3��4@��p�xE��^l���(�ztr�m����Tp��\_u�%#57H� ��:�����j~�ޭ�u�Ϝ��ֶǝ�dv����X|zk�u��jQ7و�h˛�]3���{�����:}{����wO��b��}�P���ҕ%+��jb�i��[Cy撦g
7�I�/)��ͩ|�s���t�m�+e� ��*	PжbE�iǜ�6��KW�ˡ���@�\��=�_��aQi1�ɓ�[�-�A��q��ڻ���v-4Wܝ%{�H��;SL�.u��Q��7J���m���'<�6���eRsz��Z|w
w^s��f�[4�T���3�k�����}Uf��UN�����j����kt{�'%B[�J�d�ȉ���l:�Uˮ}�dW�V��&i�7/�T1��ήI����o%��yr��=�Crrr���w����i�ܲkff��O��~�r�x�*����s�i��"3kH�q:�w-��s7,u<�΄:z�S�YBe������g�Y�":^@Ԑ�GRl�
��W|N�M�;Y���l�MWYA��ԩK#}��J�$J�-Ԣ��F�L�k�Z¼{N�,՜mͧuֳ���0��bTb�,n�x����w֞Z��~�ڃ"EWX�W�8Gi0�`���{���s�a�4u굺@�ת>g%<.��OUzJ:�|��)�aN��{.v�:���6������nS�}�D��T���^\H���+荎	1��
ټ��6�9B�L.��uw;;�!�{�)M�J�g�Z^"�>�	�Tt�_I��B=�&ei�f�����r6k��`���|�;w�g
މb�x�o�N�ڴ��AZq���j^��C&�-:Yr��n��ͻ{7����Q�N4e�pw�![�g1�:X�-8��*�LھuX�=�C�a�5�4���B�&pŌ޽p��UD��*wT琲�y�8O4	s�.�;�,D�p��ڵ38�&�G��u����Y˲8E�����Y����̷�P�-�a�ېwh���`�٪�c7��+$Vyʞ;�p\7�
�N-#*�Tq@�n��2��k`��.�>-��B�� '�4���(�1�P.��=��0��Vk�ѝf�2\z�Ѿ�zO]"�;������m�Sn��UǙ[]���Gq���ޮ3m��^j���.��Pn(�Tjݗ4�����o�v�J=/���;p�ڗȲ�Tu�ym�����+�M۱��V�ar�7�Ƃ�Y��51!b����`�P����R��W\��.�W+��]%e]����G�H�d��ʖJ�
�pM�����T�Y�s��݃�3:����c����(n1���S�K����[˛��I6*�6��X��ۗ�V�f��I�A(��G�gd��n�७�F۠�A!TRTG��m���^�]u�]u�\u�Ǐ^>���l�Tn�VU�u��w��^�7q�	 TdjB�H��m6�����뮶뮺뎼x�㏯����*Wwam��p]-��4�8�cm����,n��vXm��___^�u��u�]u�Ǐ<}}}|<�UFF�HH����N���K+�8�3)
�J�]�R�7�cm6�������:뮺�Ǐ<x�����Cd�a3mh]�Grڳ��Ӭӭ�D]��E�5�����U��h��3��ٳ�e�n���<��k���]۳ô�:�"β�DQW�ۻ���ov��ۋ���Y�z��_k�{Q�M����z��N����ٶ;�y;�Yu�����N����^ͩ�TYgY�ӫ#�����6��sn3��Ӹ����.�Ύ��W����c��R��R���b9Y����Y/n�=�\�#��BN��9jj�2�G��yy���^^^^^^^^^{����Zo=��7~�1��k����i�(���(9�I?���D3��l����&��c$���`N���������7��;�Y��p� ��͏���7f<�. ����	�Un�ࣥ���NM��".P��5u�R,[y�G����F<�^_.:e�{�d�@20֙�:b[f!�������0���ԛ�kѣa@҄�*���ekӵ<R�,۵��t��w�A��>A��o>,HG�=Wn:��{D(�9x��3.��h��^��pͽ�t�@��R��^��Y[��&�#k*綳4�P*U{���y��ĩeTh��P���T#8i�צ���7�O.��	��k��=^<{�;�{~̮l��Q��%�C���,7��|z�bZf{mn�5= -��¹���f�* ���lܿt5��.fj͘�m�g�+G^3ٽS,�&X����	���4퍾�U�t���4ʃ*���чC�o7 ��}ݑ���&����G�7X����Ʃ��r U�@�t1kd5�*)���)�$\h�]�<����߾?8�����EB���uX��{�ؿA,7Ӫ�߻�"*���;f##6L�FޤNM��ʞ	z��{gD�Vx�Jx�i��l�p�홬z���38wb��^s���u�CSy	����g]0V���OgTd��ؓYڴ���l%��5_B��i��p�����P��"���/��oW����8��==<��� ��;DRR؞���n�7�l��:m��Q�9ȷ���2�{d���~[e6����w;k�b��2���_e�p#_&}�#�+���0�`���ܟ�n*�-��2���v�����!��{������L�M�Ⱥ3��JU�3�V�m`�o�O�f����/a��C����ao�Kq�;*S��4�>��m�s{�ڈ¯	��K��y�s^\b�N<+�>>��/��_��U�JU�����7p	�tm��-�|[�޹4��9Z�%U�f��G7*����=!�{�$�5D��Mufng{:��Kvk��>���b��g����\]���zWLv����FEurُ�=ǩ7�Р��$-2l�/�Q�	�����Lj�V���M%4�M4�G+��r5%������Xgm� NX�H�M������ݞl#��-~�	���&��>�ه+t�(����3F�-�j���t����cf;7�b�R���|���@V�p���RoN��(�?�-�]��X��s���?Jó>D��u2���W��E�.ڐ�ސW���T���6��rݳeNٹ(>]�31��/|�*����<f���p��1��u�wq�ը�"�U�+X����y2��,o^����jHط@Ņm19�7�b/V�f<{O%ޭ=�_�N���V�H+�g�t([�휢o��7wq^u��@����6���.�&��N׌1��������LR���{���|��9ga�7������ ���;��ft����{��O�����?��=f��D������l1�*�v�Y;��ȓT�x�KWh���مJK�n�q��P��غ4�ؾx�T�ͬ4�iщV~HVԭ	��v2������.�Ss�;��gC����sU���,sE��x����LR���ܮ��N��Պ�/o�p�jP|��n�u�]o]�no�����M4�M'��l��z�-��S7�>a�dc��2dU(��3[ ���2h��{Ņ��1��PX_�[��D�8���j�ѫ�ŉ;P�C�I캺Ӻ{uɍzK|O�s��1��~=8��g"W=�U+��DW���n�q�%�R��7o����̛�6�x7���vk[��t���U��Y�� ���Yx���Z��;to�z7��JZ+%^�t4fCW,軜�$�v����U=Q�)�0o����3�M˃4}�=��K[�]��ʸ��q�%:�O��7�k���=�b�C�-�茳�Kn�L�Q/<�f����:t�W7�����f��"�:\E	��������vn.�j�b�FqUk�G1��.�*�>_H�n�n�E�蹎�z5,�ˬWu߈���}`�h|�ϏR3��%-��kH ���/����P�6>������1�1Kۃ���.XuFŚް���Nb?L�d�k.r�ׂ�q�k6��zm��p���H�������&�
�Z�&פ��`��LZ�A���;]� ���<����T��\^����;��U��3��Π�_~����?����&�V�:����_��i����ս��cM���X�G+wM�u�os�qt�r�G	1=���21&�,:Z�V�SB�Q���e"`	�k!��z�aȳv܏
�3�ڀ���T���lّ��Ҁ�q���`�����s��øȃ�=��,��Tt�����t�M��L��+���Em���[0�������y�zq0�z�M��;wb�5�nQ'x�M��R1�4���bz����Л���a\%46��ב�Q3*�
�szwf7A���;�э� DsH�E:�Y�{7�F� �,��n*{Ϙ�ˤ��,*�d��D���.;H�3o;|���
���{�=�{z�r ���\����Gfd���)8��?������P���W*kX�}���`�ϫ�wiq*���JQ�밺� ɝ:|�߽�<<>0߯�OsϬ��.w��a�W׊���u�T�|��|F�>H��^-�(��:�i
+Ͼ>����jcRj���M�rm�����CP�Z'.���N��W+ΧW��xa}����4�i��i��h}�85F�P`q3r����pĆf�{�j�v��������MK�o�I[��אk}���O�W^��ۙ.��p[�����}�q�=sy�Q����xbXD�30�,�p�������U�ˣ�g��e����ؙ�x�El���f�z�s�Z�5�� N�v�F�b�zzRK��3\pYHꇺ����K���p�<皽���;����Ȣ��9��ѹx^3go+���޳��	h�A;p��YC����Ks=e�l��aa���N�i8�n#9��m���-���T��/U��lؾiv�ɇ���d�F��AZQ>KvC@�7�km��؀Ëv��x�,�7w.�s�gz# �����u����/�fnF�Fyo6�1Ű;b3�*�F�	�+�T�k��ɍ���)<����3�׈�VVh�HY?�t7ZӼ^��81\�^�O�l��+8�;��>}O�P:�.���l��qL���馊a!�$�p�Ф
�[.�>��&�3D\��K�ud��[�o;rIR�[��S=����H��['@���5���/:��%F��J(�D)��!��eIi����������������-�����ۿe
�s�2�$#HZ r�toX_n!>��ЮY����Ex��N�<VL���l�WgNeR�ޏnX�@x�]�+jLZ`<5��'٪1�+x�̽�c���B,7���Z������\m߰tʪ؋;�,��/|ȸC>�:�E��c�9ڧ�|�Z*�M�Ư}�*�͢�.
g׹9�F�=I�6ʳL�Y.����_���TMr͵�5��[5k�F�ED�Z�ED�h��z���JĎG�h���i���vO�5����UFy�`�Ǭ[Y�VU�Y�뗾���=z:�G*>"j��:F&~~�=��U�D�S_o]{w)��"C,9��n=��������'�Jq����" ��4o�@�:�(���������b�^m��34��J6Eۡ��5z}z:�p�J�P�R������!��~�3�X'	����p��Jș�u�o������U����Y�=��0.�ʛL*�]����Y��"��5;Ɉc:7�����B�ىj��7���s��wM�"��gG/J���.E�G=/�����;4y��?�������?�⹢���/�-��0��c��k��+� \�/���ޝ�%�F��^�+wGsדFll����a5}��L�&LӖ�y{Fݼ���@�qh��&c��"����J�ޔ%�`U�Ȩ�|���a���t��o#�H����7s�����9���O�Ҽ�(�/~M��{}��30(A��9�]�*+���/g`k\e�ݫ��~����+��q>�գ�<����t"���!�x}��������.o��ֈI����bv�����W���0�A����,������ow�N� Fm�uKH�����U�t�[����ͮJW��Sa�<��G��,[#�7��}�}B��ES�9"�l��P�%�>R�.�r#(��a���~���x���YU%�ʯT���fb.�����r�'�cb�op�9{.�:�̳�tr��~��F��4"&y��*q��C�Vh�M��)11s9���Z���M��՚��i��,6L�`�	�f��=/�On���H��nVr�R�0h�=�&̭�M�+߼���?��?�����)E�'ꏺ�_۾��y��^y�W�B���_S;Э�{�A���w�#w �<M7�z)���"�������l�^vj0����U�˟!DJ��zr�M���]{�ܟ6��Z����,[��i� ���6q�E�=ܖ�V�U:���;KKfi^�j�E�~��t�h$��H I+{��_s|��x���j��[(�E�9��<�F�Jl�[��pzs�Lt�{wf�Vw�wv���M^tT�=ىn��r����� �l��t�؊aʑ<���\9j�T�zNY��;f���z���y=�Y�n�0r.s���������}�ϕ��D�X�[��6� ���)�3����J%o<0������2��r2E�F�.�c$�:��00`,�S�{_��܋'���J�w)Vy�^� 
r��KJE�l8c��n�vl��ju��Yݽno����@U�t(�h+��4֎�l�@oU��웸g���u�I�0�~ɬ���P�y�:h^gK�*�uohO~������?���VwvM��\� �)�S>�6Lő�$������{hmi�������bӰ�hjj�e�k�ba�
�T1y���ٚN�C���y�l5�V�~��O�s��0GĒH[�,U�{���=>�Y�.��UN��/;�<���%��Y���~�N�`|���Ϻ�<e
돿&
���k菮LF����_����=NZ��N�A�ܧ��l�噺`_��(S��ϰ��#�������� �w�����j�rJ�����i�F���F�H��1^<;�a'�Ҿ��ŲTU����G�����Uci��>�m`=Y�eY,�s�����w��я@TtS���Ғ]/�Ui,�|�<VnU�;�7��#�oN[��������+�n����v�QAL�U0�`^�{��ֱ�i--r���p�q_�^���?v#���l�	⇴^�u���2/�uц�mѠ�#'t^]�x������K��%�I�׵Pf���_���U\�gUm`�6�"�yKwj]is9��A�RG����\={��ዎV�d�:9]�����Bbކ�Q_Q��͑	k��#Et���e��PM�4S;:wi�j.W��t*�v\Z�rv��P��p��<b�����V�E��#���d(��\��Z��[�X92��o�{�	�N�a���bZ�������O��{�)�{<��`��X�bȳ2ݡ��=�SN�M==���ݖz�6K�W4Xbk��]�����r�'��!m�$�z��xIJ�D0c �A��#4��7��/e���';��LhXE��r�<S���>���CT8;q:�[���Z�T³C�cS���u��|�Wݢ�a�]�����Ս�]%L;�|�M�]�x�o�e���	��yM�.ܵ++�t��a�-���`�WF��/��(\����3�������!w:��oS��9�����.v���J\��[jh,��yi{i���2�����ՊG�CD��z�^�2H�1E:��dCs!���K����2;0�L4��z�8�Ӄ>kyu�ܿ��f�K'��x�X�z��	v�a��	Nv�[�/j�����ySez^6�5�̱J�	]e�e��y�]��r���S6�ta#�	١y����ܸ+ �߂���	�1�3�L��� �U^�t0��u�S��"ږf��:��VF"��vA�r��Y��nn�p�驾u����]@���}i䶍���]p���B*�T
o�L���ɚ�N�]iN�]�OÜZ�K�홲ef���u���c��՘ʺhmK����{n뛿��bZ��t#��Z�F��\ b;N%�yepb��7k&B�����㽡H)��v�d��V�p�G̙t�v6_	��|�:��jVs����t��z�� :qM��S��ݽn���]���W� =�����oj�h���C#�妩�G-"%k5���ڎ�����#\�P�|q]�y!X9.r�f+!�v4�(h���Ma��Mu���v�*�A�X+�R\�f�y�;JS'76eC�D�z.-~�nh�L�p4��muҕ�/s�� f�8vJ���w�c���ww�˹���֧b�%r�nm_B!�97oqƺ*��5�nu���9�Z1�Q7+w��Y�Z,R�ϱ�S��Q�{��M[6AJ�x_h�27ZA�]�:��]]QG��2�^5w3c7��+��+��L�8��ڢl)�mת�y�?:�ھ��օ�s��J���G�d�T�-�U�Yv�oMT�B�K �꽡R	 A%�Rl���)�$1X,�"L-�,�!pL���j��(�T)�fIEX���Yd&��p��ʒ+UQE�U�qB�� ڔ�2am2bN�!j�bE	���b$��Ik�(S�(CN6[$Z�*�Rݖ��}�N��pC�ͥ�w/���w�maw�qDQx�� � Q
�Q	�4��������:뮺�Ǐ<x��__����u���s�����*+.;�TnRHBOZi��ק�Ƿ]i�]u�^<x���___��Z$�$qhtw��ݟ��w���{�����Zu�]u׏<x����|�k��Fi�~n���dV�T$*�$y.
��*�M�>���:��u�]u�Ǐ<u���XW�#,��pw���s��TnE�s���e�GDL�����K�Ȭ��4���u�aq-�����',�gE|u�ۛ������'!��n\g�y�}.�{3]ͬ�m[[��m��]�u��ᵻm[�歶�8�",�v;`�$��e�!�%)������Y��8�˶�_���|V��9@b'���6�2�5q��8D�Z����h��V�uؾ��;�sW��q�mX��]�f�z�����u����p�+i`�޾���.�%LAe)f�0i�1�1�8�wM�8fUfv��i��i����β�w4�\b�yY�X�&{k�,�=`.1��e�m�5?~#O�D.����}Ϋ�������
O��l��Ж������(�r�uYs�6
[#��v�I:��w=�靀��w{�'�����W7��u��)U�v��C\��vvg�B���[g$<$�'�6'��]ު
6ڛ�gr�10�ٷ  ���\�D��Bs�x�8B�<����W\��ffm�$^G���:g9��Ν=���B��4���V��,g�O�j�͵&�u'n*aّ=
&����|�P�ltDc�j�A�&�wB��u��0�lV��3Q�I��$��x3�oW��}�<ܩȧ��c\w!UB��3������0!�a��ҽ闾�;��"��g_r��Ku���%�f�ւ�l�Ń�!��du�H�1�:�V��$���f`���d���G�s����*򫶕���/����ohg�oԣO^`�쳷"�%v�u��MNԮ-�F�]�1U�i�[+Oq4_v\�&c�[J>�8f�&��f;���7������.��7��&��{�~?������ŰQ�.x�Ш���zS��V�����5�������|F����>]��K�d�%/�e��n�P�a ��.�}|����=�n���sW~��[�7�93kO���[R�����w�0�&��;01�K�ۥפ�׺3��*R<��]�e�G�v4�J#f%�!�7��x�v������nzA3ڭ�E�l�v@�4H�Y�'���á��=c��s���������ws�E��
���/�i�X�Q��F��w�� ���Fx��'S37u����z��OUx���W���+�-l%��=؎��Be�Я��F�`��n�vi�à#�������)�/
�6����q�x�ᵰ��0>w�"���#Һb9>�I��^_Q�'k׵z�'���yI��z���AlL�ZœK��O����D�����Sy"���z^+ޭƼ�S"��KX�|�����D��IM���,늷�l�=��#�aֲ��u-��Ĩ+�]����}�7bA^��g<t�8�9��¹���Ef��ʿ�y��`���{�%���ǟ~yո����L�pE��1� ��p�O�[>7*={{d���T���B��Ke﹬jB4���c�����;�:wIh1������	{���rEbބ�j��qr�tjot�\���3�3�_��MFy4z��t����+�����|K?��M�{���XA UDz��/��;���n�q�����б���W)������Z�u�i欼RN�ݰP��#Gao������̣4��X
~��P*a/[���*���*2�D�g�s~�����}��M�n�E�Djn��<�o8�n�k���0M~i��)�OPFz}��%�i��k�I]Ecƛ�k���"���8]�������`H}p�{���-�&�=<�-1��:��rm3���2Y�������\�зٜ��c�"R������S��ɧ!}���$/��>Ov���s8�[��wR	���u9�>�G0r��[�v���2�8�*2�J�ˆp����q�ip[�� �35%����@_k�b_|��C�|�'�)Z�~?������y�'0�OJ��7׹�=zw/�&o�U��W��:3�2�l6��zu�ߦj����:L��ݻB��z�ύ3��u�5�3:�ƕO���v�{�ݬ��%��A-�K�+>:ǳ�����k��@[S��3̌zF���31褉�ä�L2Ԯ��`�ĩ��m)���Ph���;M5�ٮո��6�T{�4�
p'oݨt/,���A���:]v�<$p�������_s\~vSI�n��+��7X�3狵�hd��M�6_f�)7בp�*DƼ��{9��B�4^� ~�#�.��\�j��GD���"��q�  L�;�Y]��2�Cv #���;��t�F��'�D�#�<ɝ��Y�6��+Pf`��߇uF5�[�x�����NszJ9'C�i��$��pE{w&��P���1&�;��f6`�W���w�Fj�~��Y�f�a71G6�FA���֤�vX��P�<��aGz�r�Le)t�� l��[�i�� ��n���9J�$���jfV񴄮���r�ݼ�����I���:������|E�5��+9�zs�L��ݣ��� he$,����܉aĔ��QEp"a�B�Fr����1�b��̄���ߝw�{��Dd8I�\jB"!��~�kj*����܌�V#��u���m�9�c.k	ń��wZVa�Ǥwr�ӄP�h�J<��-� ��V�>S�~�[J�k�5j�w(��r{��yr�ƘL�{#D�j�Q1йm̶�*S���c��ރ��p��M�}�n���1ز��$,�����<�w��{I2wJJ�߻�r^sB�.`��4�t<�U�`=���eYݝ^��6�v�vtif���G_w��L`0l�=4����ڝ�z�#��w��E��{ ��])��~37����W�*J�\I>Cm��8[�#.(�H~�Ƕ�"T%�������ĸ��}ﻙwcrA�<������h�Z|ύ@�W�U졯m�������*]�x0jA����K!��{�{����pv���U2��c޷C�3 �k���Z��+�v�@����S+X��$�ʾ�d=M�Dm/"����(�Di�!_gv�f�(�:��1���ݚ��s��tQ�)b��6,m��`�|&X��َd��c[Ϟ�G�y��o7�y�"��[�宕�<GG�$:N�2X�@���l>���
7���sj��3샼�E0�q��uǸv��F�,y}���{};��S`̎h��u�UE��Z��K�E�MM� M��*���m)��?LVN�#��x\)3h��� �8;k��z�q��W8��� �>�
I6��欓�Oy�wkNeC{��/��3��A����=}5w�b ��%�d;�}=�'J�:J����2|r��E[:�T�(��4"��<��e�����W�wwv�GAq4�����j�U⻤wwUۍ�~�xi�S���f/p���f��iF;zy)1�ͅ�ؑ��6e��o�f8�ز;%;i��{VQD�޾	D�Q1�S.�-�vz@#_H�0"�ir{v�{z�nn��o!̍y95�={�g��q3��}��3� ���AVmX�`]�h���W(�h�ۢ�0���Z��x#u��W��'�����ԫ�s���έ��g�W�Nͭq��6��o-}R�s���J�C���\Oޤ�c1Z�vw�_m��s�'Ϯ�}�N�בo*�F=X�	����zi^������NkV�ᷠ*��_�ۗ#}�k�9֣��d��b*!�	�1��k�-��UPv�c[·}�����:Åa��l�5��f�q�Ԥ�{���U>9�����ɩ��v�0���h-�/*��7�ӝ�C�(��P�C��sw�],�i�h�,����R����n��tr��a�\ қ�N8Ψp�j�V�rP�t��м�Ǯ��ێV�"�q����|%鈓�����&)�����\ԕ����#�X���;]r��$�dq½[���a!m֐8
}v����O���Fģ@D�Nʸ��j����o�lI���Γm'n}>��3�����X���y�G�����i��Vn��>]�V�O#U`�<�W��7.ts��MW�~�j�p�x�v��ӷ��݅Z����KgD�g�_
�NNz�=�Ɯ�P���]3���X��;����kK�*\��k�η�wb&hw��%�n:�v����A�1�!��ϴ)�-��|<�o0�����ŋW� ::m���"�\I�\�)w�Ώ>�q�1_p��7b���i�:0�]��9�t�����w$��1��3r@��\�>�݌� 2A���[�Gl��IȺގmߕ�Y�Ѳ���F�����[�K+���Y���]z��e0�W*X��U7lċ���+z��3R�Q�I���!���v�fW��*g[3.�tnϩ�7TA:I��-F�7�!��/o[���#-�o��.5�5֛7nv�n��
;��H��@H%r��M+N�r}������	��ْy�#7����VUYђ�b`�ڨ�3}����#>�'[�Vx�1��%wn[��erӃ_̄	g������(T�*�˒�ew�U�S�J���k蔜���flg�Trv�G�_�gA�~����͘b����c�P~{l����zc	-Y�5��a6󷷳`�N���54�Oಲ�X��A�Z;`P7�?o�� �U��g����#HBz�d�H���[���Unk�V��Ev9��f�s��Q����J`n�l�G�Z��T���9�N��mt>&�.�%6�8�`�)�!����kĖQ�*O��#���ۇ}w~y�;��[u*o Ĝ{��C������t��!���T�S�A�&©ݛ�̜���;2�]F�0�d�ا��Q��my��}��Ã�+5��N}�V�IT{=C�ǗtA=����0V���7y]��Lu��Z����$��޵��X�<g]n���\�S����/
����t�n�!�7>}��מU��A���=��f=���k�4�;6�s��W��.)�[�ճ�諘����.;��`��~x���1$��V�t�9�7N�5�Y��B����1@��8㢆��E-��������1�����L�OÝ���0x٪
�p�{뫬��,���;Չe�J�k%��nf�l5G�^7����L���ux��N�N�}�LX�v���*����
z<��e��=tָQ���1w�5�0�/�\�)�bCJ������c�SF�4-o�Zҳ����?i@x�aq���@A �	��r��7�.����JW]gH`�S��LNnM֘={��]X�)���Z���{�ٳd�~+��-o}���x��a���dƧ{k'F�V�3u�A��Nf_׷8������n']+�D秸o�λ�O�����y�վ{��F9=�c�*%Nf-�A�D�YRf�{V����sP�7�F����`��m�]¹�V�\��E�p��x5�w��FS0{���H#���_�eTN�@��x�͓��f�v�$,A7�8�!��g��FS��*�p�V��L��ڣ���������GF�#PۅY�9�bkqS�8K�34��B�@S|O
%nh������E�y���U$E쨢�5L�E�*%fΩ)���u���]�������0��Ve�m��ӰD�Y�l��wxn��ni�A
d>���gefz0��Wl�zT�ˆy�(�v}3�^nk�\�v�z���'�:��K݌ ��p68���7�V6���9�M�`ռ�Y�����U��u3�/9����9�!N��⡶���*�`�u���)'q=��m���/��ct����n����/�L(cU�Z�7���r"�.�]GgZ����-Uf���k�h֬�%]H(in�uFwq�����[�ͭB[!yj�:I�������$Z�̫މu��_*���;��&�#�h
?&��}��У����J�*��$�Y�;5�*��Q�PN���ǒ̺�g�Zݪ�v2_.�6��� [w�K��d���\D� �U[Ow�A\t�:�X<z�l}"�]K�Q��]kƣ��/����\m��9p���J���ӕ�W(�k`gG=̆Z�˵�m�rg\zn�S��ᦅ'Fb���J,M%]�
)h�|��p]dX4�Ŝ޽Mn[���\+���%�><�ł�����_Smk����nRK����U�6�WU��v�;n�]���ni�^0̶a����X\�lb^���fި�z�.�W�[�7��IC�LމRz��K��C�wUٗ,lh[�)��y|�=�M�bT�;��c�Z%�my��>X�1���[r��2��p�EU�fu����Ɛ�1LU��r��\���D�	�R(D-E����-��iH;6�0L�ֱ�/R���9��`ty��r��,jF���"]&� �=#Cz�H���u]�ʐ�GUu��(��$��v6�h��2�ai�X�;gս��ەI�"S*�%roG�5wP�5�;���6��wl�͏:Į+������y���V��T)6�b��-[�G*�ʦ�7-�t�ҳF=�y�
��K:�\Y[&աD $L�=u�+{�o;Dab	n��,a˪�\�=�N���cB�f�ۨꏽ��\���鱽��)�/��V���\{`�Lq����5nn�T�mt��}eE'j�d�\g	��w6m�b�9}��=Wcc�/���E�~����x������-Sl�k�,��!C��9{9���@7�G�s�֪�\�7s:X��٬}�f]+!+G�6W5[�-��y�w����CBNُR;�*/k��A�H��m]N�y�8H,� ꦯn<Ý:c'��ɂ�&��o�l�!��\We�LF(-uǳ��R�I=��ݢ䧶��w<w�le�)�,��2���J>w7\Z��l�t�ʞ��W�ȕ4���TP�������h<�޼���A쮅Rӌ��NL�H���WL�\�Uů� ��5:
���o���Os���wM��&�O!�F��fFsx��:�(#�K4J4*;�0&���j���s���}ɒ���l5J�쭝��[n�?�_X�ګ�0D�.3-).��Urrp΁���x�����3gvT��vr���^=wC��W�E�4.���y.m�"ٵ}�u���E�c��WA�RȡǗ+r�����$�z8%���Q�f�b�:	$x�B@����o=����u�y�ڒ8�Ti���z|u��X뮺�<x������b��!�$��H�8β�39�����B�J�T*2cM6�������u�]u׏<x����wg%��IKl�f�gh���92�Ԩ�T2D�%Ï�x�������u�]u׏<x��_*QR���.�7y���H�mDۍ����E�gn�}wO8���~��8������뮎�뮺��Ǐ;ߝ������3m�@�3���Q�E��%S�#�Gy���}>�6��4Pw���̸#������ݵgVi3e{w����N�����{\�qeg)�g'Y����w�i���.ҖM�v��^sk�/7����u��q���Tw�e��d�B!8�n����d��+2#����,ˠ۷wʧ��C��޷%�m�D9m��|o���O��n���!���Z��q��k�wgQ�J
����Mb���Dy�8E("��ݚ�����y��o7����)�0�Y��3�77k�6p�\g������t�:]�Ӽxi��<�3Ě֫�h���퀶��[i�;�����)��#G�l�9��L�'gVo�8����#`sǌ��w���t�H�=�.>�-�o��gZ2����u֤My�m	$O��1�ٮ�z�v�u�N��������0�*�e�w��w�yip�����H�g�;Zm��1*7�Y�U0+��/e���E�;�[�_{�g�-�鿯��`+̯ ?y�����
S�Ufh?[�ܻ�&��9��J�k܋S�v�v�4y����9�ζ��2�[��>DVFNTb9٤��sh����<]��yH}P���x?C��3D��R��7�40l2���-�=ێot%)g�$��>O�{�Mb�@��7J�N�[�h�X�o��Ӿ��\TǞ���t#P6��2Z&���Tݸ����i��{<ul�nwZ�z�R��Gz����X�!���1�m�C���L�f��ۜQ��n:�[�fl�� nwB$��E'�7��^-��5V��鋣�4�o�[]+�;�Ɏ����>o7�����h��Vb��c�ގ�=����!P��S5]�,V-�R�7����*Ӗn{6��2r�o[�]����^z�.��,���u�\�gw��G.��Ƴ�dD�*r2��䫕��Z�`�ۿ_��wzviԣ�����C��ry�3�f����˴�|Z�{Ydv�	S�	��o �< ��8q��&�� yor�pټ�s{���r�ݎT�s$�<�};Q���v|����'7{%G��F������)�"륄��v������rm��ZjhՒv���cOӬ8uǝch�wc�� ���a���95*��e#���gO2`���~�aCd:��$W-��=�NK��A�''_ٮp���d��cx{�P,��S�����u�	빲��&���ַrN��ycY�3u)ݺ�[���҅w�ܽrlsi��� �
H��k��J��i|G҄�.�5�a�b�����pa=	]tt��-z��CT`(��J3@���&J�G�S���n����u�vI�6�wf �j�*�j�/:��V]���Q��{�p��׊����i	�>�Lr2Q ����*.2�QH�(AeBZ|�q|�|||����p�������h�H*����Ι�nm�}�WV�Mu�8[9;[��������庵�6s�vÃP"Xq��{w�G_çSuP�a��T�坹�D�t00�m�ٙ��N���m�^U��� ���7c$o2��I�[�*4���a��E^Y�=J��eb�f8ێ�Ɩ)�ͅ�V��=��g�o�(���z�t*�� �M{�}��.kC�������9�J1��"V��;�m�X��2�,p�b�K�jw6oM��k>Ln�	����7�v�o;ز�`2��xμ[e��9�{,�b��'���ff9q.�)U�RVɆ�C�]��d�h�{������pF$Q�����|(h냓r(7�t,��t�=�ov�A�O8�[k��U�ܚcW�=#�r�,:=C�ҟ�bp5ɪ���Ș���ۗ��ҋ�(9��C-�]:o���52��Z���V����-j
�yL�w�}�w]^4E��*[��I�1ӫ6�Vҩ���&;�¯�Z{^��Z���6����d{u)���t{1���}�c�s��ݬ�}��s��nS�	%͔j_�\*������_�c\[�:9�;]���wN�L�(�3"�T���tfC&}��akhڶ�w�=�N��+����J��H&�{����}S8��4^�-3D��;k5v�F��c��S�׮ܾ���y �tG��n�΍��&�cCS]w[Zx�2u��{��Ȍf`Ӝ�͔s'�r	N��X��uݏF���+Ӊm�Kzf{���4�p��c3(�	�����|s�0=��ۧH�k,��	�l$bd�	?z�_}��8�g�����j�q�*=L3Gw&i�tѱ6����E�j��#��8�$�g��<p;����;�q<8f��V��5�w��vfi��%�;�Cm�_T
��9�����ͫ��D?�S��+��ׁ�㼆����S#f^��CҀ���Nob�x��x�,��>�p��b�2~ˁ+�m�K}�M�P˯:hS�̚7:vd�X�a �+�=,h�o�M��@����V���S,��I�5>����L�Kz)WAN`t3#}�y�Ϭ���l�+7��g�1�c��]�ը��� D��j�/�R�m;��WI�c�����wT�+2���2��@����_#V�=;���ޞx�ל)f���wr�����ưg:�>�9����6�є󓗏�R�+N��H�#=^�f|v�u[��g���G)��ªe�f(Ǌ��x��Q�x�p��	'Ø1�»������6½�[��^3�d8�«�}����8��kSw��Q�3���՝>�d����]�s�����+��F@�D���zI��a�_�7��2��l���QI�ޤN� ��h��w���	vdl�D��=���=ҨlL8����ۯF�i>�^�Z �h�m��[�Z����Ì��*B�C��\d�j�}��3��X�Ũʞ��#e�^��Ǎ�4>��}��i�۞��(��R��:���v��g�mAQ��;�
�8�.0<cʋ%G`�oh��t��9y_������q�Zt��%��DYP6X�,j���ܔ�v�M��2r	�n����~�CV���S-W�:�o/j�h����Y��x~?����y���;��qܿo�D���F��5Bp�����tl�0}�t8�6S�EW't��:�Z�c�ޞP+6��5�M�|����@V[s��w���;�f]��{�2#�%"p"CG����B9��<0d���!H���8+�n�K��M���i����|�/ <���A���D����_w�g��iܨm�U�Z(ZLF�!]TZ\��
��(�����sܞs���syd����^��f��k�f�!��>�H(ws�&�6�*3w���3�r�e{�<��M��oy�Rү��8/�{���� �����ؤ
]6ע#,����Ux��3O@5������8'��a��g��a����.��*l��M�9�s��{�F0�ZN��8k��G7�F���j V�o�W�ǣ�ƃ^���z��3o#{��>����U����c��t6F%��nr��&�q��߭P����}y��,u�Bчi[�d�W�CR�WѺm4�G��c���e����ض�m��3J�Դ�K;ܵ
�t�7�N*��B�p6(`]��js&���R�o��$��J8ZM2QL���apƢuU*r�s*�U9Go��b'\��wߏ����l�͒	�I�x�������˦�D������=Oj1���b5_(39����j�F��W=F�
�wf\��8���Ề�a�����w��-��۸Kr~��d0��ѹ�i�2&��e���:��a���?�W��Mu,މ�v�/�h9�7}Y����u�
�^Rj�����X.����}�]����h�6Xh�l��W{��$�9z�&9¨@޾�k�1��{�M���4&�Ҳ��w��n��������
�ȁ;�g��Lt,�{�޵�?�!E���n����~�֟#˘q��it�K@hx׹+3wx�}����a֯da�%8&<�ϯ=����G�H|��kn��t���N9��_�Wk���XcT� b.W	9~��i����7Ԭ��@~EQa���Q�����[թ��l�}}{h��b�6\�R���F�u��M�Z���V�s�KαL ��)3;�9ϧyS^�2�����/�&�zn*�ݽR�L]Y�Q�J��P=̝�v���:�8A�^o7������K+5aţx1�k�//+����r�WtC)5شu ^ٛ�j�O"��o�#p �}qӷق���z�Y�J��?��5F��̨�2i�k����T�w�f�~��4U����z�����]��j��-?'ǵ����WS�����*�V�_��iD�kw�����9�w�����[^G�]�ݘT�����H���)�{���$׀�[�Y�`�����`��$U3�݅�g}N����v9�`���b,O�S�g�0h�4p�:~�<�(�D�o�}>a#96{V��K6���x{��y{9�ipc��v̥b)��gk�8%����_3^q��MWxI0�.��o�-;�1d��/D��Ob��dor�4�5��	Y�����{��0�^��pF�@df2���h�l~���M����'�-��1f��h�=�����f3)��:� �{gEi���}��<�gכ�*�¶�}�wg� h֔J������.P/W�z�4�Zg{��ľ\g�/un��[��
A>��Fʳ��;yFs�)��[1���o7������U�)P�j�����(���O�h���ͣ�7��zą�&��wn���*7��<~�a�W�����c��8I��[g�~��<sN"CМ�UWw���v��vfO��HP�>���m�()ݟD5�]��n
����~y���ϲџo!P�m�7�Q�ó�ys��v_ם�{]xzQE ��m��;���nlF�v��Q�驡���^t��Հ��,����k�8HYU�i��8��u᪪��M^�_]ц��Q
�浆0�K��#�[>p<)���4uE��z�Hj�Y�ׯ�+2v�oB�t�!�au�P�S>[>���x�� �7Wn�:a
��KiY8�8�uM�Z�[!q]ǻ��j�a���WW*��T\�������I���^�9["���0���=)�l� ��꽌a�:.������;�;��6ѕ�{�u`un�Y�pW���֯�^U	[�9��7��Vƫ�&r��M��}���*ej�Í� �M� �\i*�����Q�$ ��*��)_�&�ر��{zgA�gM�nM�G�:�+��n9AGv9��6�Ks��ǜ�9@���4^ٛ=�o7��=��xbҰ�(�'�qN3��Ǹ[K`��my=D�)ba��2�[.����Qw��7��*�V�6���i�!y]!j���$c,��6k�'��]���|w��=�ݮ�i(��}m��߹�<��g�� ��Ͱ>��wi�d��@{ۂ$LL�u^a���MI9�+�SJ�<�#e��1�`�P%��82c�����W�a�͸ƾop����N�\?s*}6\��O��>�Z]���,�V-�.4c����;��Bo>��ۓ���I*�#kyG��W�÷�vJ�Ň�jg4_�o�[�O(�h؈gx�@���Úܱ=��ۗx�e
��<��C���4A��|�V�Ɂt��0�[B���/qZ��ƅxlֽ:�����l����G*AU��p.t�z]v+�:�"�>����ʡ>8&�װ��v0�O}�\�y�w���%�ʤ@V�� T���_�E��TG��
�	�TYQ����aHNP*F �!FFF
F*��A���b���BF �	"���d1��aD `)F(�a �����.Wu8�]u8�9�t��A��da(���d�@b����	"��`	��$D�`#(���b)0`	A��(�d �b)��$BF*��@b���(��@`)�$ �"�@`	�� ��@b	�� �@(@`!�$�@`��$ ��U@���*�@b	�� ��@`	�� �*�@b!�$
@`!�$
@�@`��$"�@`!�� �@b��]�@`��$�@`	�$
�@`� `	�$"�@`	�� �@b��$*��� �@`!�$"�@`��"(@`!�" @b!� ��@(@`���"@`!��"�@b� `	�� �(@`!�� � @`	���"(@b!��"�@b	�� ��@`!��( @`!�(� �`���D�� H4����� �� ��"� v` �����*��
� �T�J����l��������dB"�@b	W`6�@`��� ��@`)�
�"@b!T�H���]K��]:���:�H�@b!�$B`��%ݫaF�1�$*$`���B�$b��`���d,`�a�U ҃��0`	�B
0��(��`���dB
1�b	�����;�GR~�(!   �*��b/���|��?P~�Ϸ����9����l?�������ug���v�?�~Y��������������E��$E ����8~��"���>��C� _����{����i�_�;��a�By�W���~�D��E�DH�@(EAH�AH�EH@H�@ �b) b!`	
@B �`!
D
@�$B"P�$@ )�DXDH�F� �*��D�$ ��`� ��A"! �!�ҩ]EwK�]t�P�`)"!��	
� �F*�  H�!��EER�! 
Ȩ���"�Ȉ@��`�"�"��E��@b�" Db!��(uK�]*�T���.�t�(`	`	��V �B"B ��e�p������g�O�@ dTB@	 @$��:����_`�=���0�w�}
 
�������}������H~ g�B?��'����" 
���C�O���y@_�@W�!�|?���DAs�q��
� ������\^�{l((?����Q�h������c�C��s _�?#S�.���������O�3��?�A�?p�A���"  ����D?w�D P�ÿ���D���(�@��������x�����@W�Ԓ1;{?$������|<_�&��dA�`P}<�A���߮?�������e5��|�@�m� ?�s2}p$@���*�j����"��ђ5�Iv�DR��Q�&���u��V���B�]gm"�DT�E�EQ	H�P��T��ъEjً[CY�#�{�;Cjƴ���	��*�YJZ�;�lZ۱����B]ZVػ��TڛY��i-K�����٣��:�ۻ�R�{w��,�KwnL�h:��l�[a�R��n����m%֫�M������ݵ%P���˖����ksn�ӻ� ��˺c��V�V6�i�ŵv:��l6ڭav�JZ��wn�5�   n�}m϶��oo��mS���g��y�w���O��k�ڽon�uV��޻ۭ֮��{m^�u�g[�۷�s^�n�ov��w�����w{ڧ:��{��u���η{�ݣ�.���jԭX-���a���vg�   ��/�6g�]���[i�[\���Q6�m[lU4LϾ}NK�Zi>�۶gW��Q��ov���kz��]۷�[go{��]<���^�׻���9���M^ͽ��;N��Ѷ{�����ۏZ���׼�����ը��m�gg*��  w�N}�{��<����Sͻ=����m�7m��v���w�����{��{��Sc4�+[m���n�kZ�vr�KJ�&��f��(�w,�֔��)���[=�v��Sw� ��iJ�l�-j�Uu��ʫ�C�S��kf���U��kV��;�s�M6�Y�J�jFε��K$���1��;�T+����I3{��E(�����o� �z��)kA��E�Վ�i��hG�;j�Uu�,��u�K�ݪW]`;n�k�����O3m�9�;CI�T�5lµ�qS���we�X��[A�w�  >}��Lwip�3�F��62�w�<����Z��WG���Y�x�<��P w[v�PR��۠��Qɪ� w��lԊKf���j�5��  ��ҩ��7 
6�
M�B��À�K\� ��� t�hun A1��t��RΥ5F�M��.m����7�#�l[V�;���  ��TP��p l-*i�wY��	�c� hk����m� ]ɸ �k� 5G7i@P�;��7=ݹ��U��Y�bժ�0���   {���L���� ]]n
�I�\���� �7:[��A+�� t�
n&� ��)A�G;���:gUvmm����6ٛl��ٓd�   >��� ��u4��� t)Ja�s�R��{{А��`�@(�v�� �� V�Sv��	(h���  �M�2R�G�  "��F)IT& CA���JR�  *�h��@  L@IU  J~�H���  )������?W������"�o?-������lVԦF�;�g[��#�J���U� ]��������}]w]ww�u��Ww_���뻿���u�w�W]�]ܺ�꫻����e�w�k�-a� �g�i�zǧ��Oo噎[&),��ZӒ�iGN[6��y)�B��O�NA��Pe�9�0��{x�m�R��U7.�\�ͩ*6e1�)���]fQY��Q�y�I5���u4����G@ӛ�%��q�
��:-�R֌���)ٲ6嘆ME��3`�	��S �[g2BB�(,P!5������)�t�`M�4�kf,�R�z��.�5cNe�2BYJ��[�w2'B$�u�0���<�"���{sSn͊���;-����T��,\���Lf hz�[�AT՛F�ɨ��h�gq�^RL��^;�a��(�R	�����ݽ+Z�f5m��G�86�~��!�³Ry����n���ݱ���!S�3(0#����$�KP��83sBu�QK&D�K��1��Tͭ�2,P#ke	I��K�&����-����4BV8u��-�R�V(^%�pe�L���N���ۤPX��0 ��P�����.n�Q������r��5t*4� �b[#��jl{���b'��Ĉ�wa���;[�hX�m��L"=�V�f�j��m[����]0�g
�J�y��
�[B�'s-��d�rˁ�-I��[�AL(t;���hsJdL�r�.JC�&K�zr ��������7uu�Û�l%���>��(BR�mV-�zt��HX"��Z��U-A��̭o��2�J��Y&˰�ŵ����%�(%یN%���!L�w��n��b�/+s]f�P�i�zm�?����hRF4�v�%��7!Ysv��YĞ��#i��9�r�nVܗ)�6�ՙ���%^k�\�3 h�t ܹ��V�d 1&�teRb���X���yWh���Uuv�]�Q�D\��(����=��rK�+)⺋E�h齣Z�S��HH�v��z#���=��e)r���µ��ҥhz�L�K���͚j!��V��f�m�
ɋ$$�y�Q	�ǖ�Xj����E�b�9������~]#E%][���u$�!X��tɪ@�W��@�۶�Uؕ�[ ^�ص�q\��w��Z\,�	��)�. 
N�J�2视�VַB�@�[X��F�EG�Y��N���v�gF�gh	�lIY�k n[�h;�,�,����w<f[�YC\�=U�"I�z�uĴ���'sn^ѷh�[x���PLằ�� ^�Ƥ�1m�*Ʒ�ViC�w��f��Dˠ�(�M{p�(�����*�!<ӆ���q���.K�NS���F
x��5��6ܬײF�$�f�iiN��( ���%Kؕ�a�n�m�9�$;&������MbqZ��������J��D�\�S�V��Ec(�5d�ʰ��+��X.e��(Uh�4�纁nL��R��$��en��,�I���QT�����PL�`�2�+EfPwz���bȃ,/��ˉ�xZ��{�]���{�@ ���وR��9�Z��?Z�D%x�Ƌ �ix�.b�z�ZJޢsV;yZ��xU؀��YNR@�x��=ְh�M7.�V )��@��q��N��[b�+���c��]H�K.�Գ&�LK\0&��6�GOhK��CA�9F�T�٫�2L�AM)T!*q�T�5(.n`�J�ḷ��L;�f2*�k�1��KjK
��m����l��J�(^^�*]�z�M�L�r��5pMIU��#E���B��{y#Cuڛvq,���4n�~�֛�Tk���p ��y��A�[Y7f�TwzUȰd��d�H]:č$�R�[�t���K-���0��ƍJǴ���4Lt䳖�����`�X,H�4�k�e��ݑ˳V`|:���s���J�WV�
�X��3*ֱfDb���� 
V$�AjF���9ww����X��y���N�.�S�gB��(�S�4U̥sFB�VT��\/!�J�n@��۸1��	�qZCi�^���
��@ 9��$MF����f]hw$ܺm�a��Ɍ�<�
�.�T[:�S��4�1E�����3�+U0^�w���c,h�`8�4�(��"x�]�X0IVf�.�,X#1���M ��v�bN�7�JbQ��G�H�(f���=B�m�Ku���t�Z��V�V��óH�'.*���t�Ī����c-ӆQ����)R��K��yneEa
���n깴Q��U��M��|��P���w;Z��S�%�
N���zR[��jR�S�A�:��m�Rjv��S����ܥ1@�N�3�*ҧV,���t����9�+b̡Rᱲ�r��m��)B�X������O4e
���aa*���ҵ�ۨ+�����zַ��fh��*��5ֺL�CZ�qtN�R�lj��;*����N���t�;ۈY��&\*M�љ�Z��Ld��(�܌��"*���F\�5mB�&�؋k�f:t���?!d��G�`cO9�R���4d�a���:U���S�rʉ��[
�����\�	��M�J��+��%&#�үb�u�̤�1n�"�r��J�6�iwD�@�8��K��+f���/b�jJfڼ�����Ի��H���І�i�F�ɶ��"�V/Y���ش5h��n�ܛ��V��u�
�n�CF�w$�mQƜ���q��*3�:���CVx�)����G��(-�JA�n�ןe ��憅��@�]�ڛ�]�Gّ�l�.*��S?f�[�^�t�q훻�*�Ij�؄Aˎ������``iI���������n�%�]�-��ƥ�� �������Ȉ���n�����7c�쌪�HN��Ck�%	N=��v�<M�fPIk��*&��t����$2�kF[�˃IE��,�ćt�R��]�ńdy�N��q곱ǡ�Ӷ�����t\��6R�&V�M�Z#Q��1��jMa*&�0����u��QT�@dT��SV�L?����7X� �Z�e\m�@-9$���P�i�Yw�p
���ЃU(�f���� nҏ)�
��j=�ХgQ� ��
;
��<�1�н��/�u�Jz0��T�K�v&�6	ׁe���wN@_�jڱ���Ӳܥ���C�ɲ)�65h��e9)�T�N3�{rr�l��֧d=K;����J�p��O�62�p}bDpSth�&�z
��"L݂�U/q�S� �x�ʡw�f�7-#��Y��B1
ͻ��4��K�Z^�c .Z��)YF��£E����3b�[6��S��,�@��	�1@��h���.�o��e"1���|��%��o�DL��k+z:�`�eN���QV�����3n�����(a�n�m�J��Q�1[KmR�S��];:��m���+԰C�����2�7��.^�pblej@]���9�L*B��bSn�$�Ta��Xh�DiQ�أ������ę�&�.f�f(�-25�����#Q����*�
� ��FP+�n�8�OF��F�Z�d��A˒�8�l7y� ��٨�:Ɣ.}���O
Yn�eM+Q4AG�T.鐍�R6�D��v�T�.�9�E�,�T$�p�'Ҍ�V\{!J��1Sܻ�Z�ڤR���7l�Cx(��PTo`E��!1���ɴT�5j�L�v�^�A�i��ѵ���­Yn��}t��k�oE��)��Nl� ��Wm�	I#WZU�"����7(J����b�ɐD/nZ��#/4ԔR��P9IF��͗.��7`�s\�sRrn�0��Y�2�X5��YShM_ѣww�0j����""��@uJe����S{u��V]���&f�]fn�
� �ALQY7 �#n�Gm#���#R6�Z�nإ	� ��*��-���f'w�-̬�r�75�[n�,YV7%Mb�]l�x@�k*�Wx��$�s%�_�CT�D$������/w7�@�܃Uj�1�[�wx)�ZC����\ dʼ�)� �F���Ւ���m%f��(��4��Ƕ;��m�Q	��֮��l4�C�j��k�R��m����ޱYQ�T�M"�	�m�Ȫ�]�XF�y�m,��4����\� �,�K����x�����OS�
�&���B`��jn^���emM�o2�>:���Dz��u� l8ŢZ3,4�����&��p��.�?g�����'��4E��u�]��&oN���hQR�nr�U-��d*@�0E�&4[�/-�nhYv�W3*�B�X�h�S$ �`��HY���Nmꄆ�Q��*h�������Y�-FKe,)�zՋ��`=4M�w(b�lZwn��C�a��.�K2�l�
��J��"�13nRy%��*#7]6�6���q�ׯr��U��n�:CF�Wjk��	*��+]H3L-!
���%m�hF�wB�&����C*Щ��.V`���LYZ����sF�[5�%�X�o%޺&����+)V�׻���$���Mͪ�B���MJo0+wr�a����Ѭ�y�����.��NJ�-D�o0m6�$��:��s��z�`e��d^Mvb2�H�*�����`���C&,6h�J�����KyY��{�����d�b���V�X�M�;�o.^�l�Z/)��Z�]�L�j��Fm�}t_S�.��av7�Xmt���Ū�B��tW}v�=khfa����	 �oȏ��z��M�^4�9w�.���QbMȁ�j���a�ݐ�)�ĕm�fS.ݗ���ȔT��̶YsbE%�哉b	X��eʛ�n���k�i�e]��R��e�Y?
��)c6�� �鳗���5o�Z(,?Ihc�1~ǻ�M)�Zg댥�Z)ņ^�#c԰���.��e��1ɉ�x���f�/K�H���=�6�!o/S(jo���V��c��- �j"��S0�c;�t�YWn�"/+mS*桉JE
��	ab�aP�X���\g&3um���Ë5G/fի	oS#R�U��!��.�h�92RRZ-���#(āb�ں���V��H��@w%7���e9��oc�N�0��lpM�VS�JB4ӓ5���v�����-Wpnq�و�"���Y����d:8��� �3j!�7@��#��ʛn"�y+1�Z��k���-���T�X�SN5d{n�]�KC]�qv��&9�j}�,%ỹ���\.�ݍR�Fԧ�n���k���C �H��R�kj����XY����M:H�Dڊ0�W�S0�IK��U�J�W������+�[�ϕ��4Р���w��eF�T�`�����ݖ[��^��yO�gi�Œ�:�MFbM�!Z+ZM��3v���OZb�j
���LB�d߶Λ�m����XYX��2En9�����C�d U��R� �\��BK(�wc��z��YT5W��w������˳k�l��t")Ikv�P�.���e�^���j��*86�ui��]�����d���:�mT��ˬT2�K�e3�n0�J@��yy�����9I��;���mA�j�JEfh�6��C�@nhA����3r����D��KpL���� 't��u��г�u/�\�U
��H``:8Y�!�����5� �$b���nV�|���m�o�lB��
u�BAV�Ϣɬ�RQ �f*�h����zJ.�Q"ƍ�
�7ٚ��tm�&�jXwH�#;�]�B%����4Av��m(w7'�7������R��P���E�M=8���ҕ�U���7Aʗ/ŲfQ[V@�a��\�ZA�[yӲ芵�D���+6D[1V����� Vr^�!�)~���T*�ŗ��Z[:F)-5SL� �v;KseG���]c]�ۓ(���;v%�����֥+�
O�L��[9u�l5c7k`\����VBO5�4rؔ���ˏ��:���Z�^ڙ(YXiV�n����qѢ�HG�5B�N4�U�*�*�X��Rb̬6��USq���*�ԑ�U���j��fň�ژ���m�ؖ=�1ܣӥ��Fjz�f]*�6([�!W�a��7 �46	���QPN�A�j�[oj�QX�����+ko#`�IB���,��QL/I��� �2�n�yqa�q@�o��oJە��Z�CP��Җ7TW��+��%��y���e'���ɘ���}�� )U�ss\�x�V����(����Ց�%�V���K2)4	�6����n42�VZ��wjڱ��V*�ZV�N���6µ��m(eEN��el��z�H��D�Ҵf����s�έ�� N`��-�����Y��0b�ka��DP��?�fXY-M�wt��%�ƍ�PM���R�'�(�:�ܻ��P���Z��
u,C0$j��ǵt�*@!�-� �0d� ʤ��V�r���@���L2�V,�Dɩ�7�wGn�O裹�Y��9V�� �$�t�m���!%�w���rF�(wVfMP�d��e9x�b�ܷu�cOA��Z0�s)R�E*�jq�5
meB�X�X����
��) ��;�� ]5��%lۂ'35�7Iڈ��<J��M&�4�]^m�2YhU�������9�kC�s)�y���aH��h���T�YusIƳE��Q��w%	[����X�v�8�&���"�ۼ,5	� ګ�7f
ͼ�6ޙ$oR	F�h�+nA�5W.=ѱ��v�էv�˷p����5����V����A�,��<Nmf.��{g빴e��:M;Ӹ3O4�ȪU(!YF-��jm��"������,�+�-�x�];�L%�ŉ�,L��ERX��%9c&��:��r��od�=C_2�*_��zlh�H�ˤr�$�F;Xr�'&�:LL	13E\��1[A>C��1h�tq�-�ue.H/��CcR ��s��e�i�\͇]�|�Y�\n�]�bf�@wa�C��2j������1
��}·����P��rY0�vC6;5,�Xi�wb�\4f�x���`��QmT�eYNF�\�Lq�*n�2��#�εG���C�&[��� ^�b־[֣�j������+#S-ͽ�O��3�F��ꐬ�9m<Ձ�R�CR�L��Q昨������|Tϛe�j�`��4�f�9�t�]��l�b���ݾ2C��_ur
���}^�J,��������P�(����ۡs ��,���ٔ�ð=ﰼIe,�WOn(�ᙜ�v>�]��C���IB�J�>|���zӠ(ܔըye��i�֠5a�7�7���rխ}zS4�IO��e�r��b��>59`Jŵ�djH�LSl�{e��Eݎ�!�7Z9��ֆi��&o)�SQ���)&�AY��Y:ű��$\��p,̒�A/;k��>�@Cg)��G���$�Z��*A���z�LB��|&V�++�f�ߒoS#�6�d��wX�ݮ:\]�9��eLl��5ܖ�/ub=�)�U��XR�h� U�pt�6eY�S�`5lw(�d�_�Q����{��<éJ���\���T���囕��MGsN�a��	�p��L3�tv�wV+<���}h�4�9���d��k��ST�ٺ���s���{�,�۫�8���.���7%+����KS�����7X���O�/l��MJ�(f�f��t���f�FY�B<���
���{c�{���L�g
ՐQy���m�Sz5�q�M;1ջ;X��¤�-�f� n![8pV�v��L��q�}I6��ÎY4�N�[�fjM��x���GNq�,����|7+�!.5���~q�	�z�7c����w�����rfU�q����<�bSXU�9\a	��l8n�1�<�|���)xp��R���	:��Vu�m�XS���B	����BQ�%j<��-���n�u��A�Պ,�]�|&.WV�!�W�����Ǹ�c���dښ3�ӓ緹��jv8ںc�SO+=���{z�GD�Is���u��4������z�*�빶�^5Mfգ��th����)�3J|;-k_�\���$����FZj1�i�wh���Z��ȓ��%u�M�u7��:"v^�l��f�z�Q!9��EZ,L�t(��SM��[��G�WJ���늫��Y�9U�pw�j�\t܇2v�-�t�#��|h�b73���J��$W_dW�x�-�k�� �:�\]XW$n���:�K_SmNNHCO�;y[cp���uS&�u-o&F1Y���Li�w"���rܵL��|���O(��7Y��9�E�+Ӗ{�Vfr�0�R(/)ÏXU�H��p(�7��'�}Ps��t�#�.YM��k�y���ɻ�mnH�r��G6-ɂb��-J�������=Np<Ă���LCUI��E\�1��V]��[[O��u#� {( �	�=$��x�vA�-�u��V%�nݢL�
��j:�ݬ�S ���ȞP+���Ҡ�F#�}�Һ�K�Q��T4f��J&P�ĦL��u �6h;=Y(V:21W��v9v��3��׉;����.W�R�GY�t�S6�y1�j�����}*Ԁ��PZ�u���+]�W�����FwE�V��j��pV@�=�+-lx�@%f�p�ZD�IIq�b� �^ێp�V��u�K��1�Z��
n�Y�JM�'9��Ŏ��J�G�������JY����`
��/:AL~�e�0�,�ө��K
u3��C��廱��0VL�2��n����9-¬�W��U��ra��}	c�3�K�*��x��j'X�ul��i:����ڷ[(Hze�ʔ5L�`�"/��zVN�9�HaE�N���?�F��L�	�@�_9�w/�՛SvqdI���j㿒��5�3O=�+qܡ�2-��9��Q!i��A'V���fH�i��.��q�U��u�n�J�T�-&����B��+����V<x3:��+� f�6��vpU��؀���"(�C3��bͮ�Џ8T��+�Ͳ�ھJ�['/�׈��Y���+�ki�(���T1o3%���.��5��fN\�Ԧǲ�W<�8�dxK̾ �������W���..�fq�Җf��fH����\�]c"T� �����t�26nV��'��A9ؙt~�b�d�Ζ��v��;2�T�A�O8UOa�-����K�v���g�yoD��\U�j�T`����L���@T��3X���Q2-�*����K���̼�IlSr����	��X\����v���uò��]=k{n5D��O%)��O�^t9EpP�|5��r��+δ��Bhc�ڜM� �V/q+^kW��UyD��M=� ߉"�kc���Q@~xmaF��:�����V�Y�0�u�y!���s(D�q����3@�P�_.4����YVFͺ�6pvĲ��C0*���ZC�Ȅͤ���ӗ������&��2�엹��.�W6i+f	��2��q��P��e�dԙ��2-<�J�~�/F��{5z�.�)y�'4��P/��,��YRuLܸk]�U���`����W�P��35�F��IsP[�x�%GY����PE�7E�9rB����V*p�W��<MmY�����pf�����G:6Ps��}#ŷ���7G�|��eu�v�c\^^es)ڵ��Ev�ԚbpLcGI-,U�W��J%]�:GC�Y&N��(H���W0�����ȩ�ӥ��X�#5�S\�{�����m�`�e����Y�V�S2���B�+��tk��ob��,v=m���b�^������	*C}M� #��S�U�1�m�1�i�ie��b�(��;��[k%E����P�/i_��k��3EN�;·�������q�V-��bX�č�k1��
���ߘ:��W��ߴ]��	T�{�b �;���A~�����%^;�<�H�Nz��::,���r��}65�\5j\TE4
u9e�d4�/�j���1��*��JBj����]������)�)X�J���3��-
��
���M��f�4jÂ�x`���Ʒ{Kp�� ���U
W�"#*���9�����y+��۵��S�9Q�6�����c�h��M��:U�p�Y��7g2�ߏw���V��Sɔ�-WQ�U�u����ŞG)����! E
&4��j*�y��t�Z{
*`1vEY���rR�fIb�ݍ����'�\�To���$ݷ�ƨ�7�3u7'ٝدJ�/��*�X:�^�\�X�T�>��&��\��b<�{��A�tP������S\�[Q����ݶ�j��ёT49���qV&�ngBfTt\֚@�];T���38�:t���M��a�@k�-��/�Y���젎`�ymR�R�կ��_��	%J�U�lt%ӓ�]����ne�U�6�$Ԭ�4�+H�d�+]�ġ�\��>݄���ńe�6�wk�[k�!������(�K�����3Q��uI6�z�U�P��h�aX/;/	�(t�娟uV8����s�h���Ht77�{2k�i]QF��U=JF.��1���I�1|9��v�U2]�����wv�#��%M�$�mlt��*#ݚ&
�?r��k���n�s�K	+ԟU���9���`0\����`�`�f�F&F'v���2��ُr��[PRz42f[U�f��/�G�[��[ܽ(S�,��s��I�N�%��nqs��/VV:�ގ�����cg:5����\�wy��6nh�/���^&�攷�˲�U���i���Lu#:dOSN9f�,�wXzh���%<���(�v�À6�	�{�Y*V��Ȧ���v}�*wc�ty�PM81�$R�Osdњ�I��[B��;T|���4,��_)G��Uf�gS�)������1�*"	#!0n
�h��T�MR�uם��-+wtk���ޥ9�X�#+���H3vA����=R��u����V�:��%�Yg(\W3��*;%��enÙܬLQ���w6.�)
�)�#yK�7'3��[GU^o*��ʹ�fvm�V���T+�#Yv�Z�`���ň�[7y�]%��P�->[t,�Q������nq��0�&�'鮨(�?N���U�F�a�hA�ǻ�vk�7��;F�zM×¬P�i=�*f���u$�t�����X	ǝvތ�c�*�r�Է����;2e�n��Ř�nkP�Wj`A��q���%�&�:�A,�y$Y�)έ�OE"����j�}�!�`{N:�w`�km��8�jgw{4�HJ��՛)9\j��0�fu���[�B�Z��W=ܥ��ח��welg8�Cj��K2E��4�q/k)�Gt�W��R�r��K+��獑�XAAܙP�![�4/u�eM�f������s�s���[�m��+�"��O�5v�]wm��+ư䓝,�tT{,�w���Q��bT*/��8���u��i�8���L�I�'n�u��^��(�e�#����t8�:�h��#�&�J"����ؗr�T|�g(h��]D��ڗb�Wl5�2�5WGgB?/�����u݁>�]c{(���R���j��[��]t �_<��w9W>$�j-���aH�6�@���i�P��8�KF�̰IʉPjk[Jr՘ޤx=��c�2��.M��G��a��D��Cmb���c�}\k3(�x. S4�<�݌96�S�^<��'}v��1Ea�}��d�4�=WX��z".��4��;��m��.ZA��#-����E)�Ow
�ۭm���E�z�����X�Y�◗��Ξ�5��"��R�*�`^u5x� C*��ų��muH�#3��+Pe��B�=Q�f�:�m�࣫���7Q��4������rZ��kM+uwd��L��()="hq pXׇ��X�&��7iu,̺W+{�;9v��)R��6���b5�J�]��7�mX�]�����y�#���h�;|��̵�5��y��!�;��TT�]w��@�7���&���$6��}�j9�V��ʏ�E.!n9���� ;��ҧ�c��+��q�*᷍\��	gm���"��4;+@�0KŐ�ʴ&�B
n����Bap[Ty�I��}}������m���r(ĺ2�+��r81R�lSIp͠��/g^sinWT�g�d j���hL'�� �)�����vLŅV	�ʡ�\���g	��o�Mg]<�����Ù�k.+锯�7�1]�P7�P6 8��mw/�\6��5��F1�Ǫ�FhI�i�!����Nk��̺r:�e�%������A9b�V���j���RjJ��ҍ���N���H�SV=��I�;2���I�ֻT5>�6�MH<��wd}
ս�:B�+۰o-X��F[��t�I.�X�n�HHc);��`���p��W9�f�����
VT%�"�1ek'/P� �}�s�����]p���.R������y�46��HږfJ{YFܼA�7[m�NU�A}$5S�^��'��f:��NQ1r�G��Y��P�l��]1�e�8u[�EΛ�3�*��$ӣt��5z�혋��e�x�����v�L7��y�V���ꎍ0�#W���DC��Oec���|�>8#x�	y��������P��a�����f,,cΠ[�]u�˲�PT&�[7[v�"Ǚ]��ޛ�Az�X�ԡfG�/���u����� h��6P�s�Wv#$�!�.��E;<:��Z��t�^vM�� Vx��LN[��+uL�깮�C"�	������Evj��␬A����k���g�f���x�e����D��M�yS���(m�������p�4\"�_�|4V�l)��!}6�5�iK�k���yq;�r��I�*7\���U�!�:�n����X�T����k��SS
�8��ywK��
��;�<�D����0`�$��8��Hܾĺ�u�����-�����nl��]x\\c.+��t,�v)7�@q��j���J0#�s{x�{�`Hۭ��n����Y�rXD�t��0���H�8��@��[���R�q�H�B^r=���3�^��C3M�Ŷ��
�|P�y���% �6����s��k,�Z�3�73��,��V�֙��oS��m��e�y�9�o૥��RE�k+��rm+z䳯)%.3��"�+���'������y�^��:�a���	���=�T��{zK���u��KFEqX �Rp�4@���nF����a����&�W���r�-�Ժ�D��K A;���G�/جMc�l�[�����N�� L��7z#D�I45d7X�h�3��G�����9%�c@kEҮ�ܠ�U��p����l����6�٠u2�R��q�Q�`��[\��ie�=�t�S��Kx�CdT���u��/�lAA�m��5���\�e�ˠ����3%fz�=�e�41� y)�����=i��r�#�[|.�5��@�ǩ!�p���k�Mަ���E�ZZ�%��6����!.�7�c&�X�ӫ
W#�.��i5�m^��m�%���9�6Ʃk��VN٣�V/w��Ѽɉt�-�S<6#��Y���x�9��Z�k8�y�p���$N�3��s���ᜮ<ȯc���������t5K}�yN��w�.�T�S(���ڤ꽆��D��Ww��%c�;�k�Ԛ��^��6�j&��gYp\�u%��T���3�Z	���rb��f����9N�Ta�p�����[��y����7���oy����5+ߕ��n�������e�ic��ں�z�۱hñ�W�;)�fw*�	��nsnr�
Ȧ-Z�(soަ
���2!@��A*̋��W\�QK�ҘƚA�b�N̼w2<[�s2gRQ�ŋLь=ZO��)��ljum���\~J��^�XY"2#6I��ُ(�2[}>9W1�
���\ix)Sz��Y���cƱ�+ ѣQ&��)�
��	;U�ԛ��qY4WBK�d���e�
������TV���R�n4�_�W*�Jg9#��	�Rp�*e���:+�/.JFtT�ǁ�>w
UbqR:3W"D_s(���gn��9�q`֖�5 ��=�VLz怉X*7u���vMa��%`vs�@��7c�杲d��Qُ]2QS�f��iu�c����AV5Ӝ�8�>�����
���q}�W!�ӴR�W�VA�(�N��R��
�gF��.F3}�����˔�s��Q�\����:�M�v!*ɕkO`���w݄щk�
X�F�t����C�t��h��
]�PIɫB�غ諽ZZ���v��bӉ�bx*^�5tu۶�'y��U)�<	dc�q���:sC�B�җ�N���6F��w&�a�$[ɔ�"W�ĩY���[-reԉf޼��y�pV-rƤB�x��P];J�Z�|�=u��LS��QWv8�;��)5����v���-vt˲�an�:�m^lh�Up&��u ���(�f�Y��R*]������Z0����F��~L^���-�'b������/E0_(�L�׆�w��!�[q�-rpq"���8��n3��5��2m>����9:GU����8b��mZRWeD��zٝ'<�\��7�K�q��g�$m�U�/[Ь[7(ݹdQ0*�t�XKJ�q��Un�a����r�\���k7BsW�	Sm��6��o�9.T��-[O@��3�Fُ~8�|��zh��x���¥Ѧ�dQi��+9&5���Ly%*Ѝfeuh�v*֙v�&����+2��̫�k$�k �n]۽r���œr��rA�B	X:$d��U-�ܗѩ���"M��'���,ݱ���yk��@�iZB|v��e)�>`�Z�c[�*��툮&y���2YU�R�1�>�;�*�ޕ6�Q�6�]�i�t�t
�!��]h�Ñ7�|�ʝ}1�3]��켏JIHm�p+���q�0�'�T��b'�0X��yPE[�?�Q��Y&`��j�Jj�u��Li�sz�jdC�kK��2a��Y/:+R�je���+�wx�bb��鼒�U�emdި~�����jhP��Ƌ�&��pҦM�b�V�v���6��sW0����.�)z��8*����T�˷�X���T��;!;�_Vn���*t�rF�B�˭t�B�.��ü�lЛ7\Wk�t���w���J2�ax�{FN��ЩT}���!����YQ��f���Yw��� ��0-�1@��{V�sz��Wda�<�X/�r{9�N����.�b�#[%
(n��3j#put�M%����Q�Vw��\�hV�J�O���[l�2�v·@�V�-Y�����g>���"����m1[X*|BՔ���p�ޕ�6��_�:a��ͳ� 0fof�ՎWhz(b�����
�z"�Z�J���t�����YǙoi��{M	�B�ي���`��x4��΂O��w:�&c=B���ϴ��BY\f���'Mh�������[u}g�!ֻ�pg��o�`���^Z�Ge*h0�Z��CTK��֛Wz�i���!0Lx�6
��{+5ғ͝�"K��襄C��J+MԾw]"2��ď*�{2_CzSU���,SWt�N"��}f���&�|�����x_D*f�;Wo^���$���<����
Ǒ�õRĐ� ;�+����ÕJ�4���0v2�TR��o�.��V�nm	Si�����ἳbR�Q'Vۉ�2BTj�������7�=�e����c��NU��V�{���A��q�����Tth�X���n �|,��;��BV�68�����r��,�XA�P�fsܭr�k��vƱZ�m%&q�5��3ҏ:U�q�[;hl�Vc�����ۤ����ΠtT��h�j�Gkgth	�ٵgO]d�#���mtW˯�/�ޞ8V�������sD��dЁ8���[��m�*�Ev9�Ki%I|͙b8n��fQV��u��5z�';z��l���\n.���qJ\��K{n�:����Jqc-E�k؇=R;�X8`C��Hk])L#�wx�wj���V%+�������)���Ak
�'0�u_�7s!uے��)}ڡ�1d�@'N��ɑ�v2����v�&����ur�:�j����tYn�h��h�V�·�� ;�e�ᢡ9������
����빤�Tj�iT+o�ѽ\�-����K�N���%6k
U/�D�<��ഃ�vYw�m�j����B�-�Gdu���L�Lޱ��v]��9N�Ĕ�hT3a��������j1e<[��N��K@�R��25h`AZ_����ޝZZ��[`��%V�7#�;�C%H'-Ź�U�R��%䝄j���ʺY%�Bfe���	W��6*G�<aۿ��+��X�r�cO箝�n����m� �����I�m~�4(逼�%���*�[��l�f1��Uۧ��xYY|��bT�1b���1Ð�Nd˕��zO�7��T�;n�b�xs��V�l]�LB��N� ��(�к�`�q�T����W���KZJK� ��5����s�jf��P���;A^�]��/Z�v�U�U(��ޮ�w֯AL�ʉ��:+{��(�[�+�	_�+bN��*��&�Y1��(ةu*a��x���5]�I�����L+ɲ��_���D�j�gG�\Jn&ej��ޤ���P��t*n�8r�*{��[�y@shv���`������|����r����Z)�f�Y�3kWR�`�4S�"m�C՗ap�ػU��mU���$1{}xCvP]�"�Yч���L�o�m���@pGj��J×be�fh�B8$��7M�<Bq���Y�� w��Em�,U{�B**w�:e��+X��kR��[7��A;z�em��	ES1̭�k��Ld${F�)h����ӵ�M�I��,����iV��t��x�;U���\��WN����V�eZ�,�S�rGQ}�Ӷ[��ԬB��u���{i��v��Sq.ګb�l��f��8ٴ��G!`P �-\����BZT�Gk�r�^f�7�Fm�*<):,����#ݥ�Q*`�W�V	���X�)����H\7(���sF�N�<����;\�&\�k��,*�M����|��i8v����K�������i��F�X��IN9�Sbd�s�B�I=Xy<p?��-ޏK/�����x�n�N�e�dL�U;2����
�1vc��`c��@Q)�!�$L�/<��.��VR��&+���!Yu/#�Jv��x���F7teɔ�E��Y\���7{"�7$�{�J�9S�"�5�f��$�4]�:�+e\}:l�&8�y��Da�#1��ٶ�]	��P*�'9��X�#gXh��bSY�Z�5��7!��5�
Q6�]�����3��O�z�jb��',�1l����f���4�"�AHm�7S�����ic�@��W�aڽ:�k�4E,��!W
YK4�v� ��HӨ�'������X)B�i M�k9���w=�y���Ԃ2ɗ�����.�]]��ᩣ,
�(����P�Zsc�E\Ў)hyI=�O�d��)�������횐�,���V=A��c�:��]�?=���R��vs�:���M(t��k�h3����
�$��������*6��"��4�iءZ��Z���'u#�+:��{�Vm,�6�Y�Wtb�-UbC�q� �S�tea]���m�]�;�Z���Hj�+�m�}�%���;@�5q�U��|Χ���*���N+����i�A��wfe����u��-�=%4�Ts�U�/R�j�B�oM�ƛU�9�I�R�t�аro@�sk%et�˵,&�B��)8B�۰��Eu��/�z�{�& �Wh+��f.��t�8�^�K4�m���E0"S�t�ญ���k�(F!�xb`��uiw�5Dk�Fb�\F�;V�Uțj��uԌ��F0u:�&.��a��Y��es3��o����D.�N-��ΙRcZN����j�R7|�Pힳħdj��A������s�A��+ ��Pe��݀ۖI�z�`?����]h�2�Vv�Et��g>ҹ���v� BF��ܶ��R�Y���BE]X�gfe�O�!d*�*O�X��+ٯ���YP�)<
��Zj��k��3�YC�n3����N�V�Z�bJg�K����	��Ԯ��-�n�N��I�-=�u�����V�N���t��w�0��Ԅ�#���T����/�jF��+�U�/x9�l�z���w�R���ז�"��Wr�P��si��(��[�7��4�f�������L#��j�C�ř�D��ŗ;%����$W�d��m�� �(>Źlg�S$!���x��۸�Lvg�-�!��#�XJa���(I����-�P�]H���]�R��9��z�*�қ�S�ֆ�,��K���kF^E�	�#��c��nM]wF΅��K�BH�Wg"UƎ���դ2���L6�����Ig>��}��-J��QN4�̗��1�	C�1Jn�;hmʽJ*u�N����X$v2�1��!�6�=�<pujI!V��N���ޖ��{�}��B�}i��C��P��mk�����ic��u�&��I�ɽx�J}kh��5x���2�Sf�Z�����tg�nY�C��uc�U˵[̡J0�Z�fb� ��VR��Rm�A5b�ؔ1�nh>��%E]�Ѹ(gl�
�Z�k�v�jR�4��Y� �V�6��j�T���3NPv^��H�B<��VFr$3�����rE6�����3��	��4����N���!N*G�Iĩe�
c��%�2���Z���2ɾڲC[�
���Q!kIz�&YFն�b�xn�f����{ʦv���,�N�C�;f� ���	������/��C;'h{���� �YX�`����ͨ+&��`���VK�B���n����:�Oa7-AƊIP�³FpNun���[�d�!` *�J���SoEn��}4�V9dC��n[#���9fj�yoeJE�z�*Xy�v�94�dyձr$���c.�:D��d4�V����R�+�Ѿ0�%d�r����s���Q�����Dfb��AP��2�����9����Z4q�S#�Ö\�%
wQH�Q���x�ր��i����쎅>����AQ��5�E��o:�@�M[�:�ŵ8�C�7w��t*GV\�t���ضb7�{�Aef��sLx���F�ݎ��Ir�v�˫=�����/L�a��ϯ�k)P�Q�g�j�],��[��eM�����ls(e?vl���\����mw�����Y�t�
�b���.|ř^���Ep42�TO	�*c�0e�KMK�/��a<�.�ZD��Y' ���77ub�ؘ��Q��r(3�Z-� 3b8��	A��l�/9�C0�֛�7���tź�euӚ��*�ڛlt��Ĩ�V=[�Y��v�CI :�O��4_WT`��,�fR�X�ہ	��^V�ݙd���B�����m���m���u��������j%N h�:_M(��[��ZFws�z�{�2�`@^Wnl^s��K,[7����|Xr�r��9��Jt��w
]@���/My��s�o*�`{ �
��&`�z?�;�r�Y��̎��\I��pr/�{���F��M\�ݾm��ĕ�eY��ڔ�<-���j��r�d�ι�%t�f5�]h�7�8*'i�j���I�#B}�5ۏ{�e�Z�yWKT��ղc�(�[r�ֵR�H�D�����Kk�o�j�A���oZ@Z�.b�lS���е�#u�p5;�C�c'9��à����9n��:Y��Ztis��t�ƭP��.S�+Iįa����c���q�7��Sz�i�ك�%YlgX�] ە�������jg�G�C����RHv��T�o*h�4�\-���ᒯ1Y�;U5E���Bk
k����Z��P������q_�S�E1Q���N}�yA��`�`e]�n��/�����k��6 N�he�G>/�p;�hd������ U�
q4ky�x%�+���$��5Ko"2v����B�|wiѣ*�9w-��������F��w,�2c�-Z&�Z&��j.:��x�t�X3����o/r��4��k�OX�˕}Ҙ.U��,2 o5R(_�f-[K����L�f�a�v/�Tz��e�A�OH����[�g�VF�C3�<�$ڳ֋�^q|�2�N�Sj�J�/vZئ���^6�Fr��K�.x�ؖr�02����4�õ�,���]X핧	tQon�ҎBK�1m2�C%>�7�wN������i��rP�X��
�
�0�7�^���n�b�Ԋ���*�T�؂�5�;@~�=yoCyQ��c��5�0)�| P��:8wh���au��$�ݷ��¼��J�,ݧW7D��2�F�ڎ�ټqp��7���k7eCN�m�s�R��ہ���wL��8]	���ձ*Ygt&���J=1�L�X��[s�Y�ʳtS]Ҵ*F�9!i����[���Q)6�J�9	+�a�Kx	dĦ9��+�0���Y�VD]��˨c��E�u�\�@�΂�œE3y}%����7���X��oI�Nv��K��d��[� � DA eՁ��ʆ^�tl�rkꋖy��u��_^�`�G�3I�u_	�(�.`
�Z�^`��̣٘-D�@��r������F����6K�� P�ԷiR*�V�m�4�:�U�w\6w
��ƪ��י��r�i�p�"�H�!�t"n���#5��q�9']}��4��L��P�e ����5�l%��5�a�,�a�����w^����ID�Hؼ��Ż�\7dБil�|�٠Y�6r����;��/sZ.0�/M:/T]�[WQY��f��
�t�S�k�>�W.A������a����c�q��q��ʞ�"� ̪DE[Ed��s�͘�?�Oe/u,,b�>���[�X��?�K��S��6s(���H��u$�F��7/��[j����b.XCzX��K�nݪ/3j �SG*h����_-�D�Q�ݦ���+g���4f苒82l<-
9<�3*����a8mj��n^>1�7�ow��FU̳:�dE�r��MV�jS���dC+��[�('��*fV�̝�q+��PU�7ƭ9�9�y7��Y�u��[��]Nu�����G�jU|�td�Դ�Z"�Y�����:�i��A��V��ɋ�S�2J�h�)�����z��d��qGz�'���ᘻm��ss/�9.��9��na�Q���l�EW]�X[bJ�wr���H7!��L����(~�G''+kr,�N��@"vd$�4t����8mhR	I���nN���sn�#m�h�	s4IΝN�"F��8�D�#�;m���f�Zڴ�K��!�`��3H�NR��3���t��s�X\pm�r#�Jgi'9��w.mi6�p����(����S�rC��vZ2�k�#4,��I	[�Ns;eڜVu���RC;qcVNI2�����8
"�δ�q��À�&i���[(��p��H9I�f�f�"t��D�	����*���QI';+ �8Gٶ�@� )ٮ9,Ȏ�3v�9$�V-�8鵒$�R�-��$����:I��n[nP��`�]���ݟ����ܗiȟ3!t�v�R�*հ�a[ܭ-��;��-��=*����~�G�����
UkR�h ���aAv)a���!�0m"��tL��q����g[��2r��r$B��(�Vin�mކ$S����U��ĺ\�j��[�Ct�C�m!]y\�n��PH�A���m2��I�81�.�5��풔��b���
^,��G���>��]����47�O-���^ew��To��)�2��s�S��ޟ�Hg=�(ɿkI
�<�:-[�����2ĶJuV<0P��9u��]��O�{�>�y;��(a��@H�E�N�˼�`���+��P��ea�qp# �` �]\�<n����V�,f��M�ӯL����K�o���ӵ�4m/g��7	i*��3̟m�~ R�@n�����ƺ�y`^Y�#�s���
�b."�-[^���MA ��r+\SCڤ��b���gI1Y3���V�2����N��e8+��e��"��[��`��f��s-���pn)S�&;Z��s���=޽�ZfR-���i���A_�E�"����:MzU����ݯ���8&�{����E��Y��k��8�ش�-J�YIf�t�� �. z؎VűY�e]�
��w)�(�s0J�)�i�V�y+��>Ỷm]<�R�3Z]�;�S���١'�]�%�Ιf2���z����z�I%��y���M1�)�x�2]=�28���5���,��y�T�+�Z�����O�L����}���� /�ԅ]��R�r�d�z�E����N��SF�f�$xkL[����Eƫ1�����,HP���Ш�0��Э��=�_vi��¶�e�v�	����̥u܈V��f�)�9!����D���q�_�^\�]x���#7� �F��ɵ��]S�M�qӇ� ���~�;�Ut��n�����潦3M��m4[b�^F�p�Ǜ�D�>y3�`�
1J]�_��w��S�#4� g�+Vo2b�����S���k=�Zާ{�y^PpKdԱ��5P�ǐ�Bg3|�ɾb+Y�.����������x��W�;�R*a���Vq��xc����n��kf¥�<҆N1)h���U����:fOWY悛q� g0?P>f�w
�T�v�8`8�������<��0Z[u�J2��X�S��b.#ڛ:��߼�,��!Z�Y�
��`5�Kh8�^�⵱Ă��di�bүk+mW���k�pZ���{�/�a�݁�n��}�R�|�lU��nZ̧��+��`PW��`�tӹ�U·r����2��W��Pk9�r��.ު�]�-��º���=@�6������5p��L�N���eh�:�53R��`�.�e��$Wf�	nD*5�~��(�ߜ�����c57�C~"���*�)�oJ7��(k[ٝ�M�P��=FAbg��r��V�ӛN♸��" �Z�%����/o�g�:U\�o�����ku-{,�!$�(iW^��/z%���R`8:�"�R:��׶��q�Oy>��Z<ڝ����U�dO6����2�18G�;��ssw���=���&�V�C8��iW�J5�[T��Bz|��xD5yd2�Ck�
_���=W����ӯ3\�J@$�=��yU�ↃAu�'˹4��;2��/i[����{��ɮ��/z=�w��܅�^.G�2��$��R뚳k'�mXw�\~�n�~K��g�wM	����#�\S�����`�iq��^�I1֣!-�~2��'s���
]%�8t��	�xl�Gil�]��y,�=�.�+�B/7D?�Q#��& ��i��1Ҡ��˓�L=R��tW�8,��pQn{G�{2�{`5�~�#����l����BϮ�mv[��Z�4�,����W]�^�N]�*̻#C�/1�f�4�ɝD�+�0������=Oi>b�U|]/�0;��9�:@�;��mI\�\�K.],��.5�A��k�V�Ռ�)Pe`����M��p\�\A=4|����-�T�7��"���J��:�k����\1g��	��o�{��_�3�;��ʦo0�m�t͹u%����D>5���Du׵i�vj�����*�9�<Vu��J7�k��_����H1j׾�׽K>u�3"��y�n��E�h˧t��<��������������BGeݓթ���V�K������(<wȲt*"~G��%݃���g'U{�==�xTb�x�]>�x횿Y�]{^��BE�!��P�2=�r�,���w��~x��� ���)��Ѧ���ե9a�-�q��kz��/Y�X%�
�=��$���d�"]�F�\K��a�w��C��0������ve�6���V�EcNI}���F��0�P	�����"y�:@�˷��;f��ׯ<�_�u��{��zP��r�r֐�Sr��̔q�Uj
�Fws=s�Y�tk���q�=�DDy�"+�����0V��"�^Lö���1;K�q$�9i,�0���"F1<*[�`�ݎWk/���q�����
���*m�J�qX���؁ɏ�A	�w3�m���o�j���x�yQ�k�γ(��-)��۸h�ǚ�
��n]f��Ȼ\�|zJq[8ƃ���m^F;���%�M�y���Y��)��)ش��n������N��ר#��ez�^�.��������g���u}Hi�HC���/�_������Y�S���{:�z���jطT�d�!���,�J��h�UT���H�kެ���6�k,ξ�@w��{�'<U�fC������F;F�N��h�B���RU�
�4<�Fní�O%�-bS����h��6D��#p4S(.���C��шz|J�Z��)�չX��1��t��M�_ƨB^���9,�:#.�k3]u����l���}`M�Z�tɥ<1I��鰝�B%��Pg�e��1�[2)�N�\C�?���E�޵N���ܶS�4�i.ؖ����.�z�wv�Je�y�n�yVZ<Z��B/�t����b�i��	1'r+Z���� ���Ԏ��7�p5z�4��e<�iCS˟-�Rw-��wS���Ż��c��9�|s����N�ֶ��7��������Q(i�Uw/~Cxf���S�Eۭ������%`��k�� ���3Nm?/h�;Fq��F-6�5!�G�lm;������IGh�E�����&�YS��uP� �����Xk-'����h���g���wX�1V6�b��,r�����OvV��)b0l���);�LԸ�����(é&mUbW)�c�9�)Gj��^'���#�Lx�O��˝~�<�<:�����~�4��������? )VrV�=�W}	��N�xy�w��'Z<)���]<��.�gtu�$�SUȭp���p;�m�-Ժ���'��IA]��
vy�pV�Fe�ȵ�Ґ��ܖ �Y��*����̷u���O�J
J��,뭞�9M�H���{4��T�
E��|H�'�1��V��C�N�M+�=л7��')ا	�m�5LCj#�LON���	9����צ�G��㕝%=sJ�U�ޙM_��\,��>�t
�Bb�S�0v}�Z�~Jw@�X��Ft�:�a�=���	S���m0ςZ�;95A�t@]U`��t�=��=A�[�.e*W�M�DMH���gt�4��4�<o��>�P��}��z�.��^U'y]%�I�NB����}�+ksMD� ��θ6��L�5��2�X}5��(�ՉF0{'�Z�������K����_�ƽ�թ�|���7(=��@@)C�"���z���P�*�ODj�w��7�TA��d�8mn�v'0�s�n��+q$�],����'i���*�|�oZ�ߘ�K�Z��E-|��.�j�` �W`l��i�wgh���[n�+�J.�,�R�<���#R�����^��j=��r$I���Q��P"*M]ۋ(�].;ٝvd�ɝz������ TԱ��UP��Y(L�+ͪ��K�w�����;;K���*V"*i��xb�4*0���?
Z:٦J��!�t�{��<҆N2������!��,�գ���YݶڲeFxv�P�=�q����Q���j�����JC�i���a�������(�&����ٷ��w�(R7n8:b��[䶃IB�������
��;I'4�ζ;����2W+C"�m��DV��k�Ĥ6�3S~(�4��Am'���Y"��n���$�W��;��L�~�)�=:��u��\ኁ���5u�`ˠ������%u��׭x-���48��{.�f�W���j����ĩ(���k���`�*2��e랞O.�q�@���J?�׷��B��3^��ͨgC'�e��'�S*04�*���/���! 5ƻ�z�ZC��oN������u?4��p����ij�Rj�&+~'zHK{镔:�\�Uj�Ƃ�u�2��U-�.�U�����z��vQ����s)z��b����Y��bl�˂h1��"hY��%�Z	0!�qB1C�8��w2Ey����t����dT��m�����a1Ω78d��*�庛���3���Tܝ�v2C�����jd6�B�CY��L�˻�'��E��T�Z�|���"^x��y� 8:���:w�����%�NԔ#
^R�.L�$��y1�'E���e���ɲ�{��ПM�ť�}�+ݝ@]и��9O��O�#�9�|_b�Cwc^W�f�kǆRN�"�D6�'�e~K�<�	�=�&i�d#'ZG�W��Y0%�����O$�.���쭼������
�`�C@���{2�{j]Fx����q%�9���c��3ޒ�}4)��k�!�CS�B�bk���z��;��hX�#�?yx�(�vZש;���_�S5f���d_���C�Y��˗^��#/����7�Wq�/Q%��-��H�q�!�.�!!�ښ��E6� �v^���#�n}���dY�k|�F^�d�\������F)�;��ǿ"�ᣪ]�=����V�K���@qA��胋,J�ͣR��8c����y��	!y�frXףbqp��d�S��)�c�٬�GJ��ɳ��޻�)�֊���>_��.g���=���b��<�
�������u{�Э����=XU�N����v1T�<;@��ŧZ4�UXґ{W���9�����3��ǫ��-u^;n���t����y�^����Y�����Uż�x��D9��ZzRF�b3k��`��wz0�.�Z� ��i�=���;�]�T�O'i0����F�V_�'�.�\x[��uK�㷉�m�N�WE�?��EA��^��/Bh�Ɣb��JZjQ�7������z�^�t�\�!�o<�?�8��W:�E	՜��̨\�Zuľ��Nז�e7:��@#<�q�*�q����9������vԻjܓ�H�����]�mpV��o�����Q����N��A�|{�VU��F⤴���E�ۥ����TT%�LL2s��lm�j��Mm�Gee�6�.�&a��zsׄ��\u~gx<ٹF-у$�./!`����|��^IxYĎݛ�y�؟���"�'<WZf^l�.��;*�s��i�q��K��(ߒ���P$רYh^ٝ(�{&��x�Vz��sċ��۵@"�;h:������՞Q=ޝK�;��v���N���ޱ3Hv�r���q>� �=��GC�e׭cf��>~G��_S��b�=�S&%$���W��(���������^�~�JC����c�N9
�?5\*kӖ2U�Tn�V�Ñݹ=i��gN�T��r^��9W1��� �g�~�M�[�sk���^���m��GP8�N�������0����r��@m37!��#���װ����H[�f��z��w���t͛��^�͘{1k��G�N���7P��Z�7~������S/u�_R��^TT�7����T����Ī����Z���r�`�+�5��uW���R��o�v~�����X,W��� *}M���oJeg�׋	W}깞�#���y�x�u���w���;��>*~޹{-øO���n�/����{��s(y�E�E��0���S��C�<�=:�w�γ�E���E�ZP㭽�ZJ`=F��ǦZv�+�F���qD�#���g�>���wY]2�,��{���_L�}�9ν��M&Jn����Vץa���cr@S@��~?`�0~��n�q��rZ��}��c�u�+Y����_A^�d4୬��}�k��!x+}�,71��_3Q|�������*���#��/��{���B�UoLuL �[�|��2z1���t�,^r�Z�V��f7%�w�y,��e`�D|�e����{d�``4�/G�Y)d�zKǝ��&)z�S��oV�gOqZO�Ik�:#HjB\�1�����%;�?�ޅ�)�p���A�(L׌����6)�4Ь��GMs	A}Q�
��gl�tsh��u���K#���:��8�*�tf��Q0 �$k�h��-���;\OT�)��˻�xK+�KRZ.>��W�ܔ^WN�x�ud�Q쨮�k�,7}��f��sީ��HA{	4�7Nu:]<��Y;Ѵ�6�6���1�H.řDD�P�Z�=�msU�N�`Q�:������˳�߭5�ds�,*Ef����W;W��N鼝���Nr��gt�Y`��͵�β#Ar�=�؝��Rk�Ô��A�7�3F�X����I���nox�kj	��7�\�-xW��k6v�ׄ�ڈ����ap�4`�r7J�gx�;$߬s��G8���ru<Ӓ%��>̷�,|񬰒&L�;6��t�]��������]��
7xp_�GY����}j��d��f�R�%մ�J9�]LV,��LڜR��3"AS�Ƥ|�Ч���$�f؄���T�y�
ᠸ{��o2�>S�s�j��ML����]+Fu�j�X��s�O�˭�{$�9V6
�X��[��R-q0�ޗZ��͈Ʒ&��.����O��gpZ�Et8�9V��2��n������&�	e-M�&�m�LUʶA�~5�R`���^���d߆4��N�w`[*���X��z�����{U^�ۚ�;Є�2��C^2�-��J�;4�h��h$�mIk�wn�����W���.}Ջ�����]�F�:�p��"5��Pn �edN�O�-�@�'T%Ӗgjk#�Q%s��<GFNg�\����P�f��ѽ����L(ب~���(�����(懍�EJ���'�N �GOKջ!V>���S���&|?E��߭c
��]i��%�eX�ʆa���ڶ�#����GrҌy j@�B:��I�NF�
m�ok,f�]X�l,wE�|?�* �h�}�M��m������<?J&�f�r�{���\�[%��a�W�����n#M�;��;h�r̨�ELl�Ji���ly�|�ǊZ��a9tY5��(�]��aV*ʁ�,�r-
���I���� ��at�މ����\jM��#:��\�P�x��j�v�^�v�+G����%7�3�1a-��p�պ�%�"��%��nr�	w}e��U�c2�
u(���ŤF�S�9���.g.ɴհ�j�f�v��+�M[j�����Qܮ���c�4�t��գS
���f�ʮέ�x��tTuͫhZ4�b]��祗�6⑺�����h�R�]j�	�'����9f̛к}�1h]%��9�$~=�սx�Bl�]��P�ɱº]	}%�9F���Ư[6G
bZȻ4��+w��0���Ҷ+�H>Q�+�u�v<�Hι�l9�'v�ٻ݀�JWuelX�M����;4�-��Oθv���{}wB��z�z_>��IR	 �D"941�mGZ��囊���'#��mۜ�,��6�)Va�۵:N���ά�)9�D�ɵ�mmn�9�N�$s�	A������(@:۵f��pQ�w�;�Y��GqF�(��($�mۈ��ΎrK���rq�䜐�;+-�j�rDrD��!�Iܜ�q�:"J:@8qD�8��a!8J'%;2$�B"�I.3:G�8(a��H�"r)$8HH�Rw[��n��IѶ�)�9N�,�'A3r���$s�+f���7jA�C7�$��۷	q�XI�3"e�s��%9	�g6Ȝ�N#2��
2΁m�GH�BPr�'$���!ȤI9�̓�N�� �A8�Ns�����-r���%��3�VxwFګ�n�@��;�5V��O�"�����o��7�K�G�ٛ��[�;O�Zf�ʠObW�o+k7�����LI��?�{�u��k��^��u���x���W�w�����kҬ�����������,�~k�^���˼��O�}�2.�0�B !�|�8ю1�9]K����L�����ry��[������ qwڳ�����|���׷~;���^�y_o��tw�盧��?�U��^
�.���5 4�,Ŀ���HDE(qc�q���"�%$@$���GT��T��5v6^�E�^��;5�y�C7y����^;�w{��|^����n����{U���;��>����e����+���]g2ϜQD|d��N$�"LG�bᨆI�	���F�D��H�v_M��ף�K�S����PUX�>��Ɛ4�1@o8�"$���(�jί��z�����N�W��;�/n���_w�<�گŕ�����ue��_<�dB�I���Ef�0`s���W](vy�p$����'����#���w~;����^]���k�ս������~<u��ߝ�����u����ۯn��]�޽w_����|����vw���߿0,�(�b4��TC B!/
A��M�MF�%�3k�C��?���C[��t��󯽯C��W����w��}�����������w�����Ϸw��j��`�O��5^�9v�o3���t��B,�DP�`I$�DC�5���'���~��oss��DJ ��jF@B }��"�I`24�a�,�n��]{��ۯ�x�k���K������_�;�ݼ����zU���;�ߦ� H��f#�q�!�?a�;��늳/�Ii8��N�����٘�����û��y��端C��^��w��_j�!b��0(��@�d}2(��Wۼ{�����t�k�^�}�.�޵y�������
��u�e������򥋎ݜ�ȸ���,8��]���;7zr��N�y�;x8C�ٹ���?���O���s���3�r�1S������V�z�&"�y�"4�,��Ճ�p�#K1a�&8�"1���F��*��?��גpd�^�ߏ�I�$�d~C�у�w�s�of`�ކ'���?7w���y�w�a|we��y^��m1}��c�B1=��Qb$�{��ו}�O���y��]���V�
�L��ro.,��yA����W�^��UL�|U٧ޡ|��s2CȨ�����Q�¼b�)�����N��AV��Ǻ՜}L�Xރ�3���4����r��	�* ��.4Q���xU�����cB&(+�c&����49������}�Z�
BeDa�DlRb%(��Y�n���e߿_�W��n������;��׊�,����w��������<����+��^y����^:�|�jˏ?���7�>llʎ4����6n�s���|�۬���_כ����w���Wڽy��/���@�1v��v���3C��ٵ>��lϚ������~A������v�J���������۷����$��H����O���t_�W�eߊ����z��x�����w�_�:νo<�߮�,�/x�ug_w��^���~�ﾾ���O��2v�W�s�?�����Q����O�v���a�f�$��F��������߫��'���w�ǿ�WӾ/����y_kۯ��]���TE~��{�ޗO��v^�7��w�Yeg|w���Q�lR�$������ I!+�f�G*�m�pô���[�a��w[���Ϟ���~��<w�ϟ<���g��?���dl�8C��1C�[����W�����gvۻ?�{��:�Y^W�����t��{w�ӿ��^*�\�XDw[NX�3���In�vf�`��k0w1E �*>�H�<`q�����f�w�d��gL�6�S������d$#D��M!��D��_��=�?����׋�?�����݇_<z��5ں�#^�!��:�Qۡ�����nf���a@�!RĠc�0�����;���߾���/_u�מ�~�.�����*��������n�*�Y�_�Ϟw�����W���|�^�{x�F
3u(gw�D��j��7��@dDo����u�����?����vw�v}�Q!r���Q��"+5�-���w����u�ޗ�������׎��W��^]�Q��>������}����Ɂ}Ĳ"���ͤ�s�z`r.އfl��~��۽�����ן7z^�x���~v���J˧�Ϟ��w��n��[���|w}�w�����gۻ���/k��M�Ͻn�!���`���{�]������;Aƽ�j��mn���������8~ܑ �
4>��8�� ����I`3_y�@�c�<`b�8���]����ޟn���N�������~w潪�Y�n�y�ӻ�_�;ϼ?�w����X,��,�Ɍ�W��o:�OTG}u�f�Sp�,�9ӌX�i^����]^9�d�V{Ɩ	{�g�>o�\��5�`Aޅ6�{a�r�xܭ�iM�26���ԙ�;�@�L9{���ņ���V���5Υ��3�c؝Cy��jT�G=X$�oE�ţ��N���_?�}W���z�}y��;ۻ/��?�>n��݇~~��z���~�������+��ͼ��Yޕ��_j�^�G?���{w�_��w׽��ՔaK�PF�����5_^���i�#��b(�8�`X�3�!��zoj˱�uo��竽�ھ.޷�������ݝ��}|��_S�ӳ��}w��/j�I��0ɯ�`	"�,�A��	� #e�h�݀P|L����c�o����;C�zg~��^:��k��5^�+��� Q�C��Li���S���w������]�z]�X_����{]��@�!f!�cB����Q�ig۷�Q�=�Ɖ�����D/{���:0>	"I0"4�J�f"�x�n����߯��_]������w��^~,�/~�"7�D��<�<lǈ��fJ$�@�YF��qdq�2 �]\�2�>�V�kx����v�x6;4?�kq�'�<E���� ��0- �G�@���!�F &0J�^]c"_�b�w�,����1[m�Z�bf�87kqp��C���Th4��N��Z�]4��� +���g��0�pۆpe�uU�&��5<-�N��W����R\�=��.* kP��r�o�yz~�~���_gTN1��{�X2�7�d�rC�sd��B��` 7��t��,Y�*:�_���2�Ց��u�2��|�K���]�^��h٪�C�J� �n��C�8�U��jZ3�	wwƋ�vv�^vK"iE��2h����JU�h��%�
3	iz�����nIIBg{��b�"��kk/_	���e�Ӂ�jukZ��y��b��i@j��)\����7u��kR�:%��i�9��c�v�E�F����19���OWh�A�V\B#kw�����R	s��+�ܻR]����4;����c��?{���x�SԀ���z�2�x�x�f9�����Լ*�x}�'���Sz�>�[��k��Co���\��u";� 4"`!#�i:����E�v�>�OqOe�S���9�1y����!��ᒔ��fT� Z�T#(����nT��k�!�T�N7��y���閙��`�p��Bw�����	�3���h1�[�"�FFXر,|�.�RK��ÿ���$ro0�7:�������{͌����ՓPo�QR�ыT�����
*�9�ѳ�p"�A�����W��������}y:��#��`�Z��å컅M�����Mw���,���������,��p<�?�TZ	�D����[ѭ���U�//�e3�yP]rtB�x++S��C��_(�=�� >򫳾������}'Y��C��=O̫�8� ���"�a��B�:`+/T��O��O� �J�Z��;��D\f��;�m�"$L)�������;r�܀%`�,<�~�^a��o��ifv�I�P$��7�mU�r&���6��lŪ�ߘCy����(�q�_���{�{@���cx�{E���0+2�[�l�s؇YI�%��CK���V�GC�R�Xw3�R����e�Zc#U�����_>���7U`��<Z�k�z�,䟙��UKV�V�D�c=��S3��I����¥�������}��`���u�9}Y��G���j���?�O �u�+��]$^;j������|�$i�׌E���E� �|���>#U��no������r�>KI��8¡�bP���c%��ב�D�d``�C������ҝ��r�wM��k��;ԟ�L�ǾN��BkΏ�cߥ�,۷��a��<WI΀/bTѢ��P΅������p4���n����W�[��+��m�*��Q1V�\a�ǰ%%8�M
ղ��R�P�tHҏ�A���cOv��1Q6�_�ZY���l� �W�yNhB�q�Ux���ؠ�#���ʆU�[��C&��mɛ�Y�Ȃ#P��/>��[��0O{.ץx�_��v<��Y��K�r���5.�Z��n@E{�vl �}ՏǬ�ݑH�^l�U��y>J8��R�r�˖�Ͱ^_�����$\���z�{l0��|:��gxR�{���l��w�x݋�r�$�u�'��~�UZ'�(�7L�J��Ź=l
����í�򠏝���X�����A>÷�wl�΂E�By<��x]�J�2ڋmi��=��(f��@��d��=R�_K�r�o��cu=nu����C��m�RU��N�]��"�ܬw��+k�1k76�~�ﾯ��=��o��J��R*:����ݧ0mBT�A�C�Š�E��c��#��H�6��f�����c�z���.��O����&ͷ���$u^�A�7OƾŎ�	� �dx<�睷�ord��{�`z�1*�=GG���z���x.�Т+~s
׳;��������s�M��x���h)�	��ϲ���:�ߠψ��B���i�ΛkM��A-�H(��w�;�����b&yT������'���g��.��T�*�f�/z4�Bx�*|�H��+I/{n�Bl�!�!��X����e�'=;�e�/ƫ*� �yA�*o+�z/[p��n.����Z@2դE��yr钂 U����tҮ%�}�n��წl�u��s��Ձ�(2܀FR��'�R�W�W*�zS��$���M.#vq���.ˬ�O{ގVm��_��q�2~�2'�EDc>g�u�6|�9 
�{Bq��ƽq�v=�Ӈs[~263��	�?��@���ۯp~�.¯{�.#�b��x"x{�>���j��@<Ț�q6QZ��gk�u`�����[|rR��9^��z�ܺ������ͱ8 �ueҬ���>���;P޳.X���|Ѹil���S[��yv�giL����-��� ��N#��Q�2U�R�&�wT�,�x�\�k��Һ�ͧϩ+ ���{��l@5��U�p�	�ٜ׏g��"��DL�㼲S~}ϟ�"����qUߴ��9%�/���o�g��Ξ;hH��Sx��[�`6�R*!�Z�EL^�ْ�WqM�w$Ə�6��z皠�e��*3�E����X�~_�6nݠ�U*���~���KI�����'w5�#��ؚ�Y��H���d{�-��ҋ0�½��|0ژr�,}���*�h��+�yC�[�?1⇂X����U�����[<V�����g��V��U�F0I�ާ�����Ä�k�P�7��|����7�+ΎOz�3U�EZIj3�Y��8�0�X���zc޳�ɃH��CP��jn<+�6^7�^�ψ���i:ҽ�Ā�04�GI�`�fCܾG��T�z�Cڮ��b��S����r�<2q��tҷ�/�$?kRYO�6:��En����i�q1N�!�o۩�A��ju�MA��]j׀d�M���j�z�:�2��?{�n1Ӳ��2�̼'�W+�7�4�o���e�
C�\���$�K�l�&�+;�r�ڕrޟaqFZ� ����2��^�Z���C�n������u���R�O��v�Q�x���^\*r�آ�Ζ�i��\��&v���"�i�ڸ,b���rn��Ś���[ۨŝ���ucZp]�Ԝ�{�����38R�Y��sD�x�,��aO�3s�]�1( L3�^�P��7����}%N3�SN�G�1](v���v�E�6�f[��Tz�;K�ē���r�7jD��1�/c98^������Bxv�;�b��NtZ��>V��D�w�E�v�����Kk����zoD3~H	[
fp�K;iȖ����C3��X/�Ccϕ�h�Cn�G+�{��t��jJ�կ�d��(�eu�Vs/\u��o۪���#A�U��-e�E(�=X�>d�h���W�fC����;���.�28F����g�Ui�Qf�cV檉��΀mN��H�W��?:<ߑ����9E��k���yGh;ρ���5��J�׎�.����t���%	��"_+�5�x�#,��1�[�"�Z�1[^�&���H�|ϡ�7`�k�y�;Sy��o��i�����#B^�`T�ziaT��u<*���Ŏ/@J۔����_`����e���4��e<�h|gJh�+�
����@`�c=�����D��)W�y�6V�XP�u��g�7k^�/��ɐ� G������Q�ϗ+�aX�;UE3:-%�.ҝ}`� D|b��@',�HV�;��x�D,�J�e�|^�*Ԣ��F/��C�]y.Y�����y��L�3�VV������0H�*�e�w��������u�|��36��Qh�3�U��NZ��cy�kSNM����r��b(S2P����X�B�ON���/0p|� O;ٕ��ixƤqL�������W솟���ϼ�?,�u��o@�������K�u�~o�v]�Y+�o�agW���pHwvUp�L���M=�^��J�u��� �Y��ώ��4Y��W���-Uf���v/,�"�㵝$�|�?Hi�B<��Ցk��!x+}�,{Sf_�5�^���Oc��ߪ��[�̿]�z�t��v�5A�u�摦OLb-d�D��7]�e��-�R�9����\OJ����	lo�Q8a��������0!��v�;���r��WSi#�zV]��%�P5�F-�V�W�c����}�[�ōI��2MognL
���/o�dL�Q~��`W2���t��$�Z�lz����Ի�چb���]��E&��Q��5��`O�S��
մSD49tC�;D�(�4,Zz:����Z;w�E9� ]L�� ז�W�}d:����l:u� �ug�u��QM�͋E��>�n�]-	�/���7i�L�w]�Hn�n��C��IdF�	�g]��($�hK&ntƬM�S	�m�j�Q4���� �Ӭɼ����rX��7��7�"��q�Q�3O<{��ݖ K�\+BqӇ.���p`��Uh�]��7�l��q�M���_N���_�vw�9 Dm!+ןbh�-��{��y��?L�]����ʏ��	����-��g�)U�5����e<���\���R}�x�g�ƅ%e�KJ�֗�=��u����8����}�m���;?��[~���}jC��fg�{���ߖ_=��+=v/��z���c���w�y���خG+���c1p����{�<]5[���J�VbV=��{�����O��M�o�`?��/��uJ�h�g�z�:��{�T��ǣ����eu݊֋��dԻ߄����}?t.���"����wG-ѳl։c��NI;Gc"��M�ϲ���:��A�잝HOy~*��ח�`w�+�e��7���TZ~�8�5��,�\2�ڪ� 4<5�ʃǆ[~�ɧ�ܢ�=�W5�Y���ʏ5���\�=](�*N�)��^C-����2��U����>��V�/��M-�D�}y]J�ܤ��
J3�u�R�;o ]�ऋ=���_���;\2�`�&i�|��z`|��O7�b�L�����u�e�gB;��|�B�ۻu��#m%.�toe���qZ�{�\4Z~}�::�_KM�j�ׅ����򴦉�]K��h��z�ȍ\�WBB��-���^ b�1�+�� ��U�ܱ�����Y*I�Gi�kG䥸�\��n� ��>z��QD�d��V+�k���Q�/���2�avu��4[GH�)�G�ЬV�V�Xq*I�6�/��z��:���foQG�N��<��Jܘ�(�3B�1Q5�kB=����C�DV����޼WN���V7�sb�vR��dg��{��:�n��[����L=v���םsG��h�9j)_V<�yb�ckt�!��=f�g�Ў�۾[G7I���B��(�H�z��ֶ+��Y$��{�s�Њ���g��
�I�١=�i�;�����;{bZ:��İE������4�7��S�enqLՑ���Y�
��\k��`��騷,�Ѯs^�Z�%�+{&s�:� kB��l��n�E(�"�y}��K�X�0u0���MB�݋���)��ْ�d]a�Je.z�=7���:"@��zk/w�|��cyR�7��*���O�>��yMb�ʰ� �䳸^t�A."�h}�%���h_�Tͫ�Y�:\��[&�v;GnU����[nT�
me��{�8�����or�����Hk1i7�r��I!�R��y���ɭr�L��+qV8�vF�n>���t�a皪註�u�y��b�`ګ	S\M㛶�+FA�'iڸ�171�*�{��O��҃��L�y�*��k��}�B�9��s�ݧH:D�+��uyW��ه-�z�+v�ve�uL�X��YV�5*'v�˧�S�ʹ(_�\�+�L'-�Q ��M.�-۫�4�W���j1RT33-��r[�]S3�vK�J36�D��¹��ךQ�P�q�@��Ao ��O��ܢ���m�z,p8����o��\ֺ��a��*�P�x3���y��YۋdQ�4�v�r��T��HV�p}��8�%(ͣ�{RZ��h��D��u�Q(V�z���ˠ�݈��5�`����%��cb��k�?
���՜���:��N��⳱j�ֶU�:m&Cv�Z�Rp,
s��:�T��M<��0�n�Hw2G[e�J�#�G.]J�VӃ#_Ö���zS����I�g����h�]�\o����\����vl��\Qd;(nn�sK/��X�i0���؜fI9�Twm�Z���j��&���4s��1�=��T�ɮ��G�{�ع�����ł�,�� q Sve��|��w��E�j��牣�^�&Ka_n�Е8[��^��Y�[..�/s���̆�7��������>�]$�ĕ��ӝ9E�)8t*2�8�(�;����N8s��m�f�� ��N�2� ���S3������'��mm�f#���B�k�f�#�8Nq�9�D�6��$D��$�:fL�Ah�8�㓣�9$��r����i��Q�rKmĎR8��$D�T�u�JY�Hw9Dp�8!Vڈ�RH�#��Br��d9$tEe�$��t�I��K;t��)t��6Ӝ�rC�k
Sn�8�
�D�q8��p�����㜎��Y$�Jq�P\	Ͳ
;��;,�)�`RY���A�I����'`M9���m�5�ڜ1ӓ�C��fv��;N��� B�s�q�n�q�kU�e�=X�p�zҁ"�9������EecRR'C>��7)��������.I{BzK*�qi6���~���4n�F�)Ry��z�����q�,��S(mqb|�*ez.A�<��uyBq�#� �:��Str�*z����)k�7��Y�~����%�j��#3�:��>W����?hs" �Sڑّ+1(�YӨDE8�:/*=�
wE���dB�U��]����m��+�6��[�N�f缟b�~	>�-9	��-׏g�N�"�Ck�zQ�/��y�߲���nNU�<�O^9X��Eq$I���yW���N���Ȉ�A�pQn{G�{��ó��2IZ�|��(	�,P��&�2#���S�F�)�2�kz�
��b�j|��7�'��M+5A����0���D�P��Q�y��jϹ��k�ȿs��!����������A>�<g�o�mwu[�~���e���j��B('�Q���l��>Z*"5X���CLrL��o7��#m7�ί9zP�,ȵ�S9>4Q����G�5����u[�2릇�or���+�i��T����Ol�p���4N���v$�{��-�]�T	>�©⳺���jvHF�i5�^w�DMi)��j��N+���o�%�#:�o���LYC�3vNT |zcx���o��£�r���e���@�#`�]�@:�!�sv��A����v1������rS��N""G��V�'��j��:�Z��R>�y)��ئ�Ln^�҉SDZ��v!�k��c0��dc��t����!�Pp��<����X����O,���]��#G��{�qj��h���C�l�+W��������hgP'�ۺe�"]��M�t���`�*(�Z$3M?{��9ب
��i���D�L�����=vbOxjngZ���nz�;g�	d�K$�ە^Z+�f�\�@>J ���U4�(>�Z}{���r��PMh��:-�!;K3NqD �|�d:�M��>��g���C8	�]ݹ�WѤ�m��a��
�n�����5�O�&D ����sBH�L2s���v�ej��I/ӯj�D�D�,c��Ȋ'���bhty��d�ˆ�=.�r&�[�c&��=�h{�[ts���t��L���O5��VHw�)4!�����$t�Q:��2�ټk׊�u�A�ݕ'��mJ��On�s�g�&��R��<P��} 5�{~���K'�n��GvP@h_���KˡB�T ����I!I�;�7U��M�Ɏ�T �*bҦM��U�W���3����Ն�B� �2���z�����	vf��!v3S��m���5VF7>Q�����^��E/����{���:��%oM:�j	�=�d��N���[��X�=?�UU}UG��ܲ���!���G��S�$�;�>��n��JH�|�=r�����YV
<�޷<γ��M�.����;����B�&=i��P��+b"_(&�Ό2�y��f��Y�G�{��vm/a.�<\4��u��F��ɱy�O48�+����Z�b�m%)f�o��X�;�q�����g��DH?���7��+y����Je<�lmǬ��hԨ�9�4��1�kuk�g0SU�Wr�wΎ?���`5O:�+�����	��Ǣ�;V�nN�R'��LJsͪ����	{d����D�f�N��o��|��r�i�,��+8K\:h�J��5(�͋ճ���/�6�g��6�������&W����8�R�/���)�wk��^�S�D��9�;}i��W���}S� @,����x��B��II7�󟼍^�*P�,���]��b�|L�(5�2��,��Qe�֏G涝����r�'	�z�y��Hh�H��7B��y�a��e���׭����@�ޭI:Y��j�^����;Վ��i��]ck#{��R�v�u6*������z�<��A=ɶu$���5,)]u��dC;5�\���tp�w�t
�Vy�IS��$�i��^#X�K��LcNX�����sZ��:$�����!���U_}M�����$��3�A�ބX�Ii,zT����-��*7������� �lv�=�k�Ǘ�d�;�B!���H��U+��"w�>%�,��=�a��QN]�1�8qP�+M��:�<E�2�>ZS�yb���$�O�(gB}F��� 4#р����]÷qJwڷ=�¬�c���v֛�N�f����8J�z�H#�ځ>�䎭#*�ɮ*����qy�z�-�<�Ux{uW���\$�n�9v�r�U'iD3�-� �R�p��E��#�B��N��L-"����bx�{7%��n�@@)C�"�]�����>�VB�o�>w~�����ȏ
W�o>�f���e�c~ҍr���U�� �J[%��%y:�y{�������.��!��D{�#��<�k���Y*�ߚ��� �zlyXs��;��2�}J8�J�pS#yVn=�-���F�*���=�q����~�Q��l��R糄W��g*Y���ª���:��t O����F���A��n��c�ߓ��,W�}+��d��-����HqEb���q��v����.�{)ߋ�S��>��V���e��>����r��;b9o�Ъ���x/�7KV���w]u�$�q������V�:��"��zc�y�R�����W����U������jp�@�N�G!=�&�ݻ�����+�ў��gI�@+[Y~�Cpw�&�l�xI$�]���E���"���5���#a���>��k�������Ͷ��-��|���܌��ג��і����|���a������ĩ(��)��22]p�fMar�oq}I�{�>d`�)Q�]c_�P��ע�^�Ye
�U�u[=NM��ν��L�S^�;c
��|2R4�l���`�b��A *�����KәR�fc��cR�����ߖ��6�y���k�"��,u��E�R�`���9n��Y����4��J�[���rrs!�U`��\5oj�]��|���<x�{/Ɨ}9��P�1�Zǭ�͒�V�v��X��z��MI�l-�b/�2�RC&��3>.�K3!D�KN9X��S;h��2ͫs��t���ýso��^`7�Y�3_"���uy����.=��T^���Or��`�<�}�&u6F�r.��2� ��Gr��қ�N�t^��W*�+]Z���4�dh��gj�d�6-(�p��1�FԼ��9& ��u�E��'�g�xz�{0L�)�\�6'ڶ��|#�P�#��JT��J�>�,]>W.���2�[W���i��UUUU'��A���讞�m	�א��)��B|�a��3�C9˺��%��v�,@Ll�Z�xQ/GR�"Z�2�&�LD\�&��F��F�m3^���U��]��X��Bl�[���e#v#wL^ަBZ����d�k�������Y�,Լ�G}�q��}����W;��W�BM�VO�R���5p���a����?pny��o��;�J���S��*߷��mM���(�0gYI������{�P�z�*.}�͚]���z�֎Õ(ܲ!��s�[o�}�p�����oݝ����=�c�,� ���'ln���Vt&��7
�ы�d���cEܼmyƙ��ǆ������J��d�����Y��ٵ^S�Z[Lb��˔��_�z�j�¬��R�ՃP����SL^������~���Q��h+�o#k�N��v���5�r�h��&c치F����ڷV��%8{ƥҁ�It_<��JZ/���I�ȹ����F�en���=��DD%�C���X�r��f1��!.�ǃ���4)f�����c����v'��fp�\ע� c7��oz�$�Den�������֧�=��j�N�S�;����h�ޥ�Jߍ:>�X������)��Օi�S�V�}m���oPT��<.7�b�v�^�E�S&%��(�f���1ͫsq>{h)�0��[�j&-3 ��2�Y%�!R!#a�Ӷ9�dau�h�ԭ���Ӫ�v��=ܵ� �zd�9P}�2���\�;v'��K��7�{'vtޮ�&�:�K$�8��BTk��)	5��\/����z���s�a�|�����S�HM$ϒ�[�;e�Mn)��V]������������O�69�n{)��Rg���Sb��80إ�b��(�U���-%�3Oy5�Kk�s-�8��<ퟟ0jX\�uwڠE<�v��,:i��;��BͿb��UqT�c�R���ޙ�����T�r�<��ϫ�`�uK����>1���㌜��ߑ�$�p���1ہm2J�O�L�2�wކ:nz&o֒��vu�	[L�=r*���m��sUxE��9�ų���-cܝ�NᷭJ�`�|i
��Y���YQk9(��C��=�H�qa[��S���foYW�iU�B�l�3�-L4ڦ^�'�?>5�{7�-�gu[�-p�T����)��#���ٴ�{���𦂊!M^j°����d���b�Ae��E�h=�[5X[-e��"ؔV�V����zٳR��m�r�3��K:��j��(}V����=9Q�?��LQ_��_g�N_z��v[/���!~�r{Hm���w�����~���������ݞ�����v�����y�������6�kg��}s�-?n.��@*D��.UZD�̯��B�奸�мS3{�~;>�7LUΧͫ����q/gdk=ع��!�m�_5ڃ�����%��P�ạ.��
�7�b�f���'Z!�Qˆӕnc۸����!i�zd�>i"�k]z%�ݡwQ-;A0P���5����=;+�sD���R�"�w�y��K��u�6�"�R»�eַT6�cT�]G:�^�c�Wyu������T�1��Ɋ�A�

�W�T��N��J��sk͵�@!��v�g���7qs��������PI�d��`(�c+:
�&k)����Y�*�jn�2㫓g`���αs��ꪪ�2r uā����%Za��%�]_����>lg'�"����uPMH��{�p5��W��[Q=�綗�V>�Y9f*���Fa���;�F/]��m,��z�
P��2Q����2����{�1JG����g��rn�����~�oo�^싌/�S��ň!���MD�dq�)C�ϻ`�T�M����q?C;=X��Kg�R�ccS0�j���l�ܵ���8�mֆ���J~��ۚ���ǌuzk-��-��63��
U�c�ZUε��{Ď[�!z�����}a�g�,vZ�l�`�d MM>e�l)8�mS�l�$��n�����R6�w�'aƐ��y̴��������?aȤRU�R�4�,u���b��
s,�wR5�֙h���h�Hi�J��ݙS8eIWL���厲Y��JR�援�d�Qj�ۊ-{���()%3:�?���7�J�KȾ*p���k;��Gs�~�lx7]��������W�u���M��]�JMnNo�R���K����yOlv��Z?�O^@Ȃ���L�AVs��",��㯅Z��7T����V�0�sr��fo{��!�F�V�:[�:��1�I�'v��[���YZ0�����>�ۄS/���/���nR�6
q*��~y������x.��x$����|��&�?�-��T�6鋈`q{�e'}�&�*����ӽ{�u��Ҳ!^�.&�W�E�RE�K�;Oq`�s�{+�͚��%љ��	�倵�yf�db/M~)��BXl:�g�ʾ��w�+�'��Nx����Q���s��Ț��JI�~������i��y�P�v�� N����E"b��Fכ6�?I��W��x�j��L�2}]3���3�M�U��Q�DH)��h�s��V5�uV۩�Zf��X�n�1�n��Q�%X���s}1z��l�.e[~5��k��J�)�╡���l5wr����ԡ.�n�'����yC��y����U쵟U��X��ίCT�����/�_���R����V�W�K��b����Wi�t���Tz�˫��b�t����XqW;�:�bӈS�� b2��T��p��.��l��])�/�d�ֱ��Z�������Q%Tn���F@dŰ���yo{�S�W�qY��R#�栻���ȕ%�\0�C4�f����Ԇ���!����-��{��a�-�UN���m�\(9)�K����4`>�]�3��Neoy\��Od��ނ�>��]ҿ��ɸEKD�m�E���,�e��V�f��}���]��۽�29ܥ��b0և������t*v��<�f)n�lw;9)sۓ9�C4�Y(��F���O{fEXk��#{fX#�m
��H�0҉� �}������O;w�.B2�{�;S��t�0��]� ����]��3l�@2Ȗ �;h`�+^oK�d�f�'��M���dҨ�v&���Y1j�<����@˦���:���Z~���2���hu��.Z���T.iǓuV9k�h���e��(b�j�]�u�18�X[zb��e:U�]E�h�]��=�˥F�~᫰Q��G:Z�A>����QaY�7��^�,a�i��5��f���
NvF�0��k���	�Ƹ��oov�5�3�A]�ٮ���	�:�T՚l�U���P��(��� h���7W��ڌRa���)��ku��+�,6�|㥲ݍ��:1%��Y�.ù�Ocx�K}d�}��F�o(��Z�5"U� D��-yw�����)��JfB��K�>ޝf.�ث�/�^,����TZlZts��>�Wpf^>-����c= �T,��L<�8zP�ܬz�o�8�2���v��bKs:�bG{��|� �1��-�n�O7M��-��������[��9���'�8�:�\��L�8�Z[H�Yq�:�U�5f�&�(($�*�siL�|p3�P,����IK�7�՛��jWO���g{5��4�s|�<��EE�HC�&r:4��vTe�LQ���K9��T����1o۫)�@Ҭǵ�a�ȼ�[3�����f�{W�湣wVӿʏ����g��X��n\�Wp1v(�@��+7X3^3k�T;�n�P��\/�
1�c�ImR�4D@���e�i�4�+�Z��%1�F�B(Fp,�9#,�ժ㸩�H�~��/-K{"�5�p�,�j��X4�.0+z��w���K8�g	��R�	p[V�\K�1u/,MXQAJ�*�u�4������"N�����3��ƥ��7�"�Y��ݼ�]tm�&>�&�R�*����S��Y0�m�"򲡃wq���dA���l�Se*ꜚ̹۫"��
˵4L��l��7��s���[��֋0,�:�����q����Ǥ�mǝYd@\f���޽4�S��W�Xm���
]��#L�eN��wO���/s�����OD�+��Ht52�[e��ټ�vOM�0	�(�:9"ʬβB�B��":K���2�ˤH�:#�;kH�PE�GEfG\�IGqNB]']%�%@۱.H��.B"'�"N.��蓍�DqAS�Etpu����'G	�EABG'9�Hf��N����s��r��ӄ#�����8���q(:$�.N.B��h���:N��8�N:��J�����-���gmڠ��<I^5mx��De�� �A-	�@&��y�2��9S;<�CW\�gk�%�j8�5��\6Fu����u�L���Ԩg �r
�k[6�vƶ/�m>�g5j����諭���3YŚi�q��S0R�-�۟,86�չ5���V'�����v\��gP'`���0wu
�vƷMm�R�c���.�][�ʼ� a�dƽ�7g��'6Z�v�^�Eya[^�Vы�M��ϒ.�Cb�H�t_t��[;��!ת�����!�QM5���;���T�@��,Q}�SBU�Z+K�</^�l��Z쉿4*�3�L��bq�y�=��X~�b�q���,��U�y��Z���0m��5	����R�,`�<��{۸Z�B'��R,y��FՕhb�Q~��w���Č8���2b�DKٕ�//��:�k�̅�I[?�����-g���=��}ws�^�h�rk��]�L�"w��+�I��w���/i��J���-�í���2C��`aQĠ�tv'�MŚ�Tgٻ"kJq,�&�Dc5[�t��@J9����i�x0mGK&0=���/uj�՚���XuE��@,3�bGM�i��Q���g.����!w:�jy��@��'{"���g�3)�3(�\g 7���#�2���v���=����.B(_h�]H�#%����d[=������7�s�"d���(~7ܪ�Ú٬���)����S�^�ޫX�ή͢�L�ܘ����ƿT���������|k#f��v��y��Rg�ι���K��;/[Yjl��Y��bkQ��]R�����4R���춽·�P.���ZY��
��:�P�=��<K���^�Ynq�?lk�o�'���N]-Ox򍰬ǆ�Z�i�IRͽ[r���cV���츝���ʋ��!n�2j�Lь�l�Ǭ��:�4Q��o'��p~H�EMUߡ����g�
���N*��k��A'��󏛂@�k�>��f{�����]�
�p[}��2��c��G�j{�74�2ʌ6�++Q:u3aŔ�-*l��wp�B��zN�߳�y��{Xfb�W�vgU�.�gn��ǬJ�\�)V
��:s�*������f��(*�XKg�`WՈ��T���z8b���]C��W�d?g�Lmxt>���-�#eTyE7�*��m�8KФSo�'GW�*.GxDO��ï5��p�ޗ2;P���J�9���.^����gi�SE6���hj-l�Y�U�𕮄r����s���f�{�T�cIn۞;FT����-ǟ+C%L���Ե#.�^�T|�&����ut\�ҷ?9�׮D����F�ݯx����$��*A�s8���{j���|�����%��]Aq+�fr���n��V��-:�m7�!�ˈ؎��۬y5y��wk�e�Ap��t���v,�����2� dӾo/d�"�mx�h�MM����i�_���w�>HgR]gŕp��׻���� %��Ky$Ϛ�[6&���24�i�1Lm�������5�6�Me�%��LNK��zY	�(bB�̍]S-�.P��v]�c]�X�8�.�j&+(e=U�k����w��x=����{�Ei 喻�V���p�z�];�Y���^�zPjX����m%*�Q�`�qT4[����K�	I}��=�=]�I~Y�7��,k�l�m�Y`۫S9E[xc�%�^b_n��ʆC�ד�N�{��䗐G����t��'��r���C�C��Xڴ�S��b�:%���O\���ǋ�,/>��/PO�B4�f&�����c1��r�n�Z��X`��N4�����
�'n�\ݶ%���4�Y�������{��ɕ�j�mk�[|ܴ�T7|ʭɪ�n�X=WD=��T7�>kp�4�i��c/4�hT����d�Lʋ� �����������^]�ս[�/VصTq�+ra���R�Y)�b�����.���N��g]�I�N���{|K���c���w�55!�~Cn��%݆�$�^1�3���z�ʨz̘	dB8�N�kr�'��h\<�̛u�i�l��Kk�g\���zN��|�P�>�����5�>C-�� �0R����l� ébe��;hs����U���ť�\ւŕM�J���i9W/I�YsL��R��H�s������Y��}�Sef������_���w��sdJҝ'MkH�����$l:�u阖���9�y��~��3�����f��id%$؋��Ml��L�_��N���G��η��8��2��B��Ho�M�
�4}D�Xռ7����1.�E��_�O$���=�g(�T��&7��;:<z�����\��:�)W�`U9P.U�����]�\� �)���a��krI�Er�m�}�xD�y��ff�R\Z�)�cr�ѾlWq'uE�^�B}JP�d�55C���%�፟b��ڎ@l���r��4{�^����^�lV�D��eU*v�T*8O�'�UlWs�V(}��3�X�O�����Lޫ�+ʵ�'��Z�������9�Mx��{{���߽��|�k1�鯪��싴�`K���5��t+	j`QT���d��a��ƭɪ�cus�E�ֵg���0֝t�����z׶�
��7
�������5.����Nݤ��3�fg��2j�F1R�7e�Lm�TS,+kЊ�f1zq�q�{���^n��g{�FQ�~��J`-5#L�5'G-k��W�V=��*wޒR6ג�ď�u����:^�ʫ��ߨ�1�ȽV
Tk��d+.;Iʦѳx��}����R�2ꏴ�cu�P�����?SO�o����[t��[
�Ed[���M���cP�ǹ'��}K���T��ty���ز���9��P�xfm��/�ݨ�J�D?l~��)��X[���Xr�Z�z�Qw���N�D�"u��<;J�,��Q�x�O�x��������������̅*;p�n�e���[�>ehb�Q~ϑ�2�؁�)���zI�3׊����Q�����ݬ��Z�i�%�>
��H�s�����lE&|��.ʞ�����"�;Z�Ur�b�B|J�T̂lT�E�%I�BcY��4'�,��*�5<(g9q0UŚ�'Sd�=`��z���dg��	�G��y��N��hxߞ�h��.㓽��e<<~{�ίN�+1�����-�6Iy�g�M����׆�o֗��oUs�vX�,�[A?�t^��䓄k�2:ح3Y�FO���e��(}�{�,ؽ���wsm0��K�{���Аm�ۧ{,��[>�W���(z�g�1v��У_o��L{�w����m0j8��1aj�6�*Y�ͫma��U7�+��ܜ��<ζx/I/6z�C��LvZ�l5�mӨ���
�+ڰ��|ixc9��^�r�1�C�ː]�,I��:v	�ٜ�,:ӆ�;�N�W�V1��_�'Ms�%?��ez�\�(�/	Qf��I73V\{*�
��c��@%q�--�C�w-��Α����_#}1�PT��Jj�5l\Bf�3y�;�����{��I�ȝ�q�:�[I����Xm�D�(�׫�i�B�]��tp���F��eܵ�RU`l�Y�s-�]�\��t���g�����{Q��i�++�-*l�h�}j�ֽzAm�O^������ËG�jJÞ�m�#��׬U��R�`�R�}�����l�6�V��rɠH�U!��MA��l'��j�2`����uHZS&%��T|�<j�V�u���Y���[�[Y���],�U��ŻLE�V�e��%�>
��ѝ�f�өo^���߽%sԼm{n�����b����!��t���4��bЎŲt��j�*���!`�yq�]q{g�a����h�Z�a�d�� �)�6Nvn�-��k�[F&�FP}�Y��0]�AWf�͗U�L�QC5ռ����e�Ejd,���.q5��}�W�[��V7�xz6�J>�WB��+�%��v�uCMfZyX�v}�_���Tj���-̻��I�z�aI������.�����mH��Vbç�졣�@�d�=��I��b����S���f>D�c�7�d�s�$V�eƌ�g[�)�O�ި-���+�\]���9by��fo5,�}:�Xu;ݓ��q&[vS5�d%�JIFJ5uKl�B��h�狢փ�����~���{�ʏ\a��m�۫{!�j�J���%����ݻ��	�i�@:�{痹}�9Qs��kjX�F�mW������y5�%K\tk}�"o7��v߂U{��<g:�Ϫe>�U'��kk��b,��F)�&�j�PFr��y{��ۑ��5a�g%G�̛������qy��7���o�dQ[~�K\֥���dNÍ3vr�]��J��Rƴi۷0�y�f6�*)c�H���4�)̤]��k&��@UWJ�(��Fv�<ځ��4�*�.�S,u��E�2R�`�3���p��r�#3w��~��>�V��V��~�wi���~I�e��m��-(ˢ�b����������`�ʹ3�B|���i�ߠ���wkB�O��L�E*՜�{�Q��:u��1ݧ³����e�w�e��Ĝ�\�㻋����,�Jdݚ+�փ7�jJl�y���&V�d|��L�r���( ��y��9]s�H�u�	�by+�R�.�Z`<]NX�]D55i㱠1d������������UX�d��RD�eC~�t�!n/eyM랇��d|�^�3*J��5��S�s�[BT��0���s���qD���;kI��$��Q͋�T������9�RuL�lTE�1MM��aְŏupV1��b��$�6��b��n��&kT��vEid-ex���^��Bt��xHd�.G<�N7��U�㋸�d�N��0�⷟����ӛ�g�l�a�d�ao��;L���y�G)X6�mz��e�º�M��ԥ��K�QI=K��'����o������w=�vm�1��6X5,4�4�]����ɜ(�y6��r�A^Z�6��U�m��YuV�ՋίL��YS�!�Cz��JQ���jV�r{G�^Z[r���5nJV�5\5��LX�6�J�ZgM��mV��u QZ�Lb�|���h���aTW��μ��5�,�s������n>O�*�QǏ:*`
�T[��xNei����v�r^�Ӄ/r�.���n�gr�Ymr�kWj,0'Xq��J��0��o�a⫰h����4�I	.L$ԩ�^��O$h�&�TR���ٷ�E�:>o{��lF!p��H��2�)��f��ژ� �XV�V��/�vn����%S�{�Jw��(�xtv���{�s-�Uؼ=:yߐC����V���̅���M��v|��뼿Hp9�&q�=*�~��mg G���װ��=�b�x���+B�I)��Q���m����5n*���^̭�XK�zI,���H^,�Kqաx�T9m��2���؇3zl���3;7�,���[�1��u��2�RX�! �6��36g8+���6���z���zz�̮W2�HK1+]'MkH�JS��g%����$�R��Ӵ�:�����Wj����ZS�fI6!-�e����@U�j��[BTD�.��%KF]�Q>�v2o/�o�fyɺ�2G8���h�Qk^��m���)|�-w0m�oR�����UQ��Y�d�H͙Of'P�^T��ha2�M�}o��vYa��M����r��)�W����cO-�8���eg���nv_F���5ϻA4u�DBk7AdmM��٧�`"W;]���Y�	1fZ&Ê�Y� s8e.��U󧰸dV� ����eEfAyZ;H�OnY�V��\Is]��7�D���j��������id��ѫ�oWr<��9:��i9!|&�*�������)��{����&;/�/�gݶJ-L���-φ`c/m�r*{�U*+V���6�Ku���x4b�rF7.M��-�c���ڨN"«�ֳ�K(F�f�����:�"{�	��긡C�������k�u�{�2FgH�+6���k��#�(����v�:�3��-�T�5���r�%#��:IR��@Y7���p4�/2�]AQT5�8sD���|�c\
тXeΣ�t����r���뇩Dk�WQ��W�����v�*z�f­��R�}�u_fJ�ՍU8�r�'-��^7�H���`�GNv�S�q0�i��C]��̻dVq귷�
ya����J�E_k�bC5)MV�tсAV���F�V?����Cz�F�킆l��p���֜U��vsj���M��o��b�cAj�3�bE[;����3�5��fF�bכ����YfU��{ U&�ʄS��C9��D��*�H��*S��;3$U�%�V��գ�r���;�T�Ir�FC�H$�S��2�V�r�<GVQN����o��e�(,ކe�5��.��]uq+A��'V);�$�c�eѽyRA�C������Y�Ⱥp�p�U�)�Z�B�Ի=�2�Ʋ�������`��p-U�ӜVb�ECNY0�[@�x�<�W9^��/E�}��e�	�e��wJ��;8�B���Ԣ�ևWt��Ԫc���.�}i�Pge�团�^�D(�P��a]@4ڥ�a��<�e�?�L)VӘN$0�!s�J�k�KT��wMt�l�}�خ�3L�p��Zt�}x6X��gUEsb�o,�i��7�G�n��p�V�m��b�o9ѩt��7�h4^ΡEҕ:�O1���uk�:vT�Pe�O!p��8GW��PVw;�7nb����;FQ�tR�u-�IL
�4���iP��dݧ�,��ù���͇��@ʝ��K��ڴJ����V��X�/��.�r�k�8�I��Ze���X�\��W_7���MZ�Dz�*�F%�l-�{���E����e��p�����S���}i��É�Ⱦ7XsV��)�/K��AQ�+����K_U𧕎�*-H�}�<�dB��<�Y����+f���p��;�QB"�.�9��=.�]��eI�eQ˾�r����i!Q�w�a[k0u4Y0�tf�<�M5;��t�B�!{mXd�2��ź6�fJGN39=��j"���$�N�Yy�q�fqىtdJ:$N��5 �y;"�8 ;;<X\\۬�K�Q�j��Ŕ\twft�B��	D��NQ٥s��A�Y�x��+�^.�.:r����r%'qua%H�M�:��uwGqV���䓺.����(��.�`G�YԐ�NTqx�H@R��;��I-�TAHpI�0�ࣼeM�����"��ζ�w%9	�vvZT.���+$���rp�:�Z�蜼X]��C�eeJtqGi�w��9)(������:'�Q0�EL@F	��X2�<�s�EӋ�퓅�iޛK���{{A��vc�9}�;�9��(a
f��S3�ۛ��r�b�v]�����}_R�kw�'��k���ש�U�Cj�d�WT�����\ʶ����]�2�����u<�'���V
޷V*ob��x�f�\U%���^��a��<�L	7E�!����g������yJ�7��[9�Ka����3s4�9�e�M���ڹ����f�l5��P���6�
�1=�c@�q����p��Ss��q��갡�g��g�
��A�՚��c��8Q6�[�7Q��e�nJ���a��C��ʈ�� <�Vh-��q�m�	���LS,u��YF-*l�Z���Aнw^��2�Q�;��1_m7�c��2�g�IW^G�e�z�EbR�6
uG�_�@��}`�aŐ�J�*t����s(і0wK��ԷU���LO��X,�&Ԛ�����X��m&gmsm��Y�ʷ8ۋv��ĭ�I[��,TF^�/S�kE[e���f���<64S�����v�b���*�x�%�ˠ�epY��Y6M{5tp�w,��C�g�����Fv><��"�\l��͚���R*������i�qsy���dY�(\2�w~g��[ͫ���mjڴ5R�dK���}_U{Ih[�}�����.M3;hu���E��V��q	%k������լ+X�����-��/,����i�!�‶���ǭ9s���*��q�k/t��y��M�}����/r�"�W�(v����T�߰��6Se^�����i�1;'��,����uE�jk[@B4�i�1Je.�;
��^�u	����� Ѵ�͸�����oK��W��~�&�z0T��%�G�^��~R"z���M�}=��'>�[!��U��f QE��[U#l�Q���L^���U쵕m���~�돩�/o�x�hs�-+�i�nt�Io7����j�?7��v���6j���y��_T��K��D���?l�3�|��6������J�+	e���*�&�b�\mK@[0X�и�&�Wy4���槨+1��YO�Em¥����$p%%��	�q���,��v+!0T{S��{�탷���1�6A'g��^<���Ŵ��[V��+Zw�u;��SYW�;�Y���M�cj�8���b�$z{����6�:�I(,��`���;���C��D���ɫ�n���ec����%�.;�}2�d|���0G}/�R���O�$Nj�s�{��͙�� ����"�X��l�"�e:M;�ܵMF5J$�d��v� �ӌd�EѲ�d��r�JY��N�y��m�E�/�g�_Z��C�C����&���[�=dV�ڭ�k-^j3u��&ģ���K�מue��m�~��i��ƶ�\��w�=�Y��v.�-4)BXs(ˣ�cc�ٵ~ve��%���/Q	OIf���Ak�d-9�B�*BA�$l9�g�c�2�ɾ�^�Qh��~^y�Oco=^�Ƿ3r�NS �mSSG��%�l:�1�Q�EN�@m�3�j�I�,��n'�n=j��7dMid%�M����lMl,)����E�eVYh��a��(���rkφ���g��yk��OT��{<+��	�d{���)﷩��0'Y�V�^f����cy�Bg�/�.�!�����,�j�կ��F�n��ٯb�)�(�M�% 6��Ѭ��6u}�٩��n�N��lNKh�ʵ*���-��0V�/D�H�C�Qm���ֱ-}s���"2J����9�:VZ2�������H�j�J�����4����}G��e���E{M& ��ud��M���[��<�dP���,o\�9��f�b
���m0�%���T��ܞ�y��.��$�(f��V�.(�%MΉ�O^ꣾ��G�S�}�^�d��J����a��jܚ�(��q571�����!�=U��U�~��J�� ��¥�b�|����@Vs������'�>e�3X#?d�:�U]㏠*+�
ڄV�z��KH����R���Iɝ��~����?�ͬsHp��M��Ӽ ��og��@ͅ�Z܏-�#�RZ�-����φ��ּy�2�4�i.*W��Y+k�1+ڽ�'i{$��y"��k�ʴ.aI4�:�>���6�Ϛ�ṏ�ud�U�}�����~�F���Ŗ�n<��1D(�a�>G]��Aؗ���}�Z[���b�1;�����e2�RXΥ!	��&4k]���kz�T>#A���p͝J�@!��.Ț�.g������U�H��uױ(��
x��u,���]DK�9[�Ic�{�Ďtku����*�H�ǜ��WC,��'�9Ʌ�N�hр���J���*q]%�P}_P�� m#�.o��s�<�N\��c7�V��A6*"�i��cc�ř�[�
&�r�wk�e�Au_�a���ӻ�u&�5�zƘ�*
��}Vq�\�.�9��m1i55�I�:�|�-w-�O��5đ�,,b\�BUjr��#S-�Bi&|���k�ϖ�(R5�|�1��;]�Ϛ����Z�Wx��j��)>8tԘ��O������]��}�b�^o!5۽��O�qL��k��Lաm���#`����X�f�b��UqU��yQ��KoB>��X9���P�P���х�}e����Ņ��M��^n��e<�Q�m�Ų^c2{��1��;���6jƙ���Ae�֛b����)���=e���X�{_Bv�gw���S�g�)���v^6�a�e���u��[l��1d��DEÕ)Nm��	n��Њ4�Z�I{���\���	�l� M�fPk�5��j�c�<n�y�,��f�׶�F�[�����h�R��b�b�z8P�5켂�ik���6l�Z�s��V�'fR���%%���nNw��M�u�»KS�H�s���ܮ���c#X�n��S3�]kn�ckW8��HZ�W�Vfd��l�,E�#�.a�^��^8�'ޞ[S;�Vn-��[��vA�-�i��m�0o5A�^�{�钥��t��;~Z���c�������/�λ���!��GxάE��4y�2a,�'���kr�+�ehd��ن6���)B�����r�yC�gU��-��ʳ����F�����v�S�8W�,��[u�"[��}�P��B����+��W�����q�#$��Fo9W/X�_R��R�g2���;l(�t��K7�������	ڞ݌כE�������RlE魊jhF�"W�n!͹��V��Z��d�^��m����כ"kK!)&�mQs�����X�����X�������D����+)�S!4�HZ5	ಌ�
k�:����z{��OSJoA�9Z*{l"g��~^6%�o��9p��jZ�՟o�d:+��up֝�m�5���+��<Z���5f;����Z��o�u}�Y��3:��&5�F�ܻF;z��b�Xe(��|�wV�7��;u�3��N�.��3RL�7[ �7�ӭC�ͥ٠��w��?36�eeN�������W^I��>÷ƫ1=mu>t76W<��Y��k�ft���f="��o����s�����T=阸���g�[���%�R�FM�`��,6�������ylVǕ�U�܊����2�/Of�W9�vc���W�-Xn��4�c�����ybQF�-�9�ӂ�ݲ
�_J��xL��X3�"�֨��¦��Z��m�T,W��ZM�`c���߲wd2mƗ�I��W�4� ��VN�8U�.�S,u��n�rfnA�yy�Δ���	�������t*��6-?:'���N�I�����r-������N��l$\�)R�:�>�E1s�*�z�>���ts��k4SQ�D�I��T&,�Y^K-�$0(B��2Ȳ'�*�
/abՎ�=u��W�+�V/n���;L�-t���V��	���jֿS��O��n��ĳ��-�����yx��F��|�,��N��r�Ee�&j4/'Y�_'��r�Gtjn�*�{,�㊺��į����2@�M\��ld�n����+�N!���T.�u�Ow��H�ں��쀊̴����}��̉j17�.�+7�׎/,���N��ب�hb���)���hE��#��U��rܩ�j7�F[7dO�R	&��"/2��z����� �u�����N���<o�~�a��rw�M��0�ⶹ��w�rq��V��R>��x��Lf��d�F5ࡶ�����v�����=4�c�i-v�b�b�,�5�#���C7��eҢ���ct>��	��M�he��t��w���7g'W��f��G��{}��k�c�xk�v���k*��2{I���|�{��9�$�֘Qǁ�W��)J��Kx�D�޹vu;���$��>
zK8ܘ�RИ�Zز�t�m�d��1j���qu����f�Q�⤒�X���̰�gR��kf�X[j��d��K�(jt����ͼ����E�k4�Y"�_Z���@�`l>nڝ<�dnF��-��+.��} �+�bG(�@�
�#1�.ޜVm���ȯW�u��F�343ҵ����3��U�]XY�:W0�r{ت?>���s,b~V�����e��&�2�dȳn�+vY:�t]�/j��,pМ�7����.7�G��%+�����4�7���p���sr��uIk`�3E���=k�:&Z�r��<U���8�3�ΝXO���{��m���zJ	�B�Mi}cM+/LݵĔm^MB��l5]�5mG�nf�%{�YZ,�D20�Y"�e	��(JkQ.؞��S:ʷ7��k�bṪzϽ�D{|�X9d
���zIE^����>���]4�V�w�%k��ջ8ZB�v���ed)�XIn�ya�-�o��{s��gzbh��#Vr3o@���3\2a�3�a�\�^���Y��x�7�N���a|�?�v*�L�w1\ە �-'�3���$��x.���@���{�?do�(���9��q�c�f���r�v[v^�R����y4��`3^/�W���yΉf��NH�*�F�V�6�,26�n�Tءm��Ⰿb�je�z��SlV9���}���=�ALz�g�ʺ{Ξ���3�?^_m�N�f��%ٖ��/4�&�vM%AU�|$��	0ܔ�Vަ�f���)����;���N��{¸�W�P��j0Q�c��1k�F�{^�G-S�/(�Ϊ;=
��B�7F ��n@:�!g���sNIh�:�Z�no���N4���[�!褲��pf���Ƭ8~�̡+�쥜�7�┾�VF;�.�w�O"M<Vjf���+�N~�R]Z���J���+/�	!��qe�������:Ihl�����-�[�F:W�]�}jq�'�K/����nW��o|�7��vUj̥�9�Q_�����3��m��ܷ]��$��{8I�/5N�a���3UL�2U���s�^��JR��NU[�5E���U ���U>�C=��υKF��Td�ݯ1�-+�V�-�u����P��PGi���/o�_i���o��y��9zQ��N��a��35n������0�Yti�Cy��6�:��|��ʝ[�Kܑ✦�,8��s^BӚB�)V�e��s��[B�>��f��}�/����,��T�s6�����R�Õ��u�e%j��ObVRr���<�Щ;t��c;B|�+"�<fX���Z���r���=t;v��s��B�R��j�KI4���1���Aܾ�����3K�'�bk(6p�"g0�ˑw%�-��»8V`tf�4kXA8�-�ܮz�-��#�kD���2n�+� ނ"�U�ope+.�t��v ��n�]���*��y\�*�iL�x]$��ݒ��{A^K[�x�;YJ�	�\�'��+�}��c�S��']��� �L�w���\���-��}J��V F��q�[����+.�.���;��:�k���B��ͳ��b��+LAQ3_PE�x��E��|�I����p�����L8�嵊�����P��>�n�u:A#4�u]�X���\;����g!I��$�O��a��T��Č6%Y!$�p< N���r�ۻ��O�rĢm�F� ��x5�wӶ����WJ�=ݽ���@��
��G6�X��iF�EJ��]�*鮴Xۚ8/D�bB��r9��LwL_\'!��u]��f3l��Z������`�������뛵]�/��̹�`�:��ޑ�5��A�[�Kn�aȤ��i�-	׹sa��:ļ��6�3۹8H���^8�����Qڐ����W{��oQ��p�k�8pV�4�FԴ��tKU�
wv�<ys0�y@�E�t �1��h]b�M˟�<�vE)��E�����!p0cKô�@�T+f:�ib�Am�]pn�~Z�8�#؄�o:ژ�G,�Jm��%1��Y)��k���L�[�f����3X.�MꚲA)ה���.X�<�4�f艅��H�7�Mi��
�p�P���y�	[�pA�3"S�,B{z�D��,��Nzزw.6�<Yd�܇Z�k�5��m���V�P��l��%��Z��Tѹs����0f����(ʚzN�mc�Ӥ* ;�җ�g����N�\f��t���+�ƛF򝻨W������o+�t�/���!�fN�"��#�Ɯe��P�ų ��]H��y7'T���;�c�i�&�v�;�pgW0Ȩ�V)1*Ex�:9c��v�����۪�T2d;}hR6�Y)��{��;�[��S���(�}�U� Wb�h�l>Řp(i�P���ln_�9�R�@cA�d�ݔ����i���>�����i�Y��R17-5�Mv�j�{��/�ZX�[i%�W��Q���.�rR��K%l�7���b�Z�oK��+��Wi�H��q�K�;L�cH�����۝#B��0��8�X��B�]D�wi�J}"��r�q�πKh�[I�R]D����t��#�H�+�N���b][E�T�	�N�]c�����On�I�Y�\�q���y/��L  �@&�*Ӥ� �(��,�(�8��ͭEqI�Gsn�N���#198�@E8\��W�9�U��Z�;nЬ��"��Ѵ������ⓝ���5�mZt��'8��:	"9L���m��!� �.qe�H�m�#-.9+;9%�<��۝�֥�2��m��m,��7E��v�2�8��Mk���lQ�'A�^-N��H�x[�q١GGA�e��aͭΎL���Bp�mn��&h�,�'mnD��QN�#kDtvՎ����3��6�v����r
N�Ð�u���k��ڱm�dɲ#�A�Zs��r�w3\Pe�]�v�U����e:����iN9a�vX�N̶ݜ�����)�1����iQ�1�8��
Wv�÷#��̙���ed�2�M�2�,}���&d�90fN��a�پ�����Ν6)W���o$D��3ޥ�f"�<SSG��Yn>K�k�\j=���yH�F*�^����d�(ZY	IT�����u��� ����^��V�i#�M��׭i���)��É{�y��
����f��:Q�{�v_��)V�ӓ���Bo�/`�hҞǛ	�j�����A��xA{)Okޞ��/H�׼�%^�o��o�b�'����>�����s����㸐�����m���-˛Wq��>exHz�]�[��u�w`<�h�G+t�7 �5蚕CIT��+a��f�wYE�����T�@�W٦"kt�8���\-�,=�S�(�~�Ki���H��:�'f��u����OH�X\j�/8�����E�d�Vы�l���6%qBT�8xQ/��3��A�n�M:`�WH��^���n+�K�j��7�,�b`_ryk�+z`�N��FVؕ�M�5��:���S6�F��(Щ'e]�d@B��K����ܜ�W����Y��O�]��㬨��O���c(�5Z����]�%�Y��E��|`|:-��>VƇ��w4,]kޒ���:�ϜuA�����`Oٞ��cpW��=���Kxgro}ۓ�WKp����x��T�}G�d6�sm|O�yEZ�ۆ��f�*m^g4n�B�RYo,�-
P�gȲ2��l3���N�%v��e�`�d'�4�34���!i咶JP�3�ظ���[Z�כ�8u�1z��Aۋ�V��yhn���ب�h*��nk��K+�lj\1�9%����⨺����Te�vD�jA$֣!�՛�ŏL ��Y%iD�z�Z�*ra��%��唰�����J�5xo<��]��vi�T����u��O����3T�:����lYCk��z�༦���+�q�^Z�5�Ck�B���U=P��B�Ѝ�g*��b�v�di�޾N���Sb��~�[jj&���Aݓ����ۼ1�����_ػ*p���Q��h����ā0�w��[%C�`ݩV�ѧCj,���5��]���B���x�W�	�(V)��E��ӛRt����VJ���Ơ�ʊ&R��Y��X;3�핻�i���p뙆[%��LOr�C3=P`ϡٲ��q�b���M�d�fߵmϖ
����/����`[��T��S>��f�lYa�ӨW����^9H�ՍU�xI�_M~p��78=����^U�1)Ϳ'U҅>��r���o�>�|K�qYl.�^���Ow�P�S�`��Y�������T�>娻�^���+�d�"��J���j:�e�o�^|�n2�uੋV��1�=�4���%�fTΕV28��׽�ez.|�}�Co�g����/4
��:��<�����'1���@զ��F��]^�ǖV�O�ɉJdLܭ��/k�X��f�S����t�ά��6��S����2�RX�d��֚i2WI��������m�>���r����n��t3ǥǴ4L4�9Y�Ƥ��k��VOly`e	u�1�n'�nә��6�-v�	Rwd�2��J{�%W�tbPӉ��]r�41<
�F�+z=�Й��N�����ب�:�(��{űB�.��r�N�n�6��H˾�u�F�sZjL��\�6��Z6��%�5sWκ����s�Q��F%��iҽ�Ņ�kn��Ӄ��݉d�b�b-��5424��l��ȿ�u�;^r�+��f���^~�o�5��ZY	I3�ꋖZ���hdim3�-������m��X��ej&+J�k)�6�B�
��2�ģ%���[`^(*&��<���l*^jA�%)=��{�ϱBN��ދ�����g	[~��E�Z\����k�6Gm��j��X����~���Ƅ��Bs���:2��N���麒<�Q��[r֪�)���W�]ˍ2�-�-��XZ��d��-u�#2��zm骴�����?E8=��rhݫSj�y�4;9 y�[��DVX�4�S����BؔV�*[L�p*�*.�D�8�
`�:_��,��1��f�.���sW���;d��JEex��l�R.�P�Q����L،�9-W����l���Ι2Uבtr�c��+�r���D����B����=n�W�C{�j6�y������)�����g�ߚh`՗����N�X�g�����2�,�j���q����+�����Z�} ��6=:��4��`&9jKra�N��6&H������ӳo*V�i7vQb�*tGGp���Qr��x�=��ބ:;�H-�d�J���O^�̷��vΗ&�o���7#�?P�*�VZ��G{ay��\5,�Y�mx��e^�Ӥ�Ʌ(Keti�C9��N,ڿ;��]���đǯ�GOI/m>MK8���-���4l9�g��8��3�g4a��N����ݞ��Y\��&���I�2	�SlSK#(h�u���0����{2��D's邽�e�j1��5�Y��K �kZ�E�jjPn�42wZ;��~��ճnM�E���=��evi����}�tX��̯M�sVMgc�o��l�y�:Ȏ���b��?��1���?=���~j��s�/���zmŦ�SeMD�w�L��<�f|�Qs���+Y[�_��>P{2t�U��ܒ��V����l���UE�#��^��ze�1��C�5ۜ��T=޻v�Ё*�֩i�%����i�j���z���Z4iU�${�T�׻8,]i��m��͛Z����Eb�^�Y���5u���F�)y�7��C���ѱ'jup�r.]����C��YJ.w�e_-Cz+�u%V-1�'A\WVj��[��>ԯ((�[�҇���8�k�p{7uזe*ķ�ŰӞ-墲Ow>h���f�쵖gP�I���ӛ�mAZ��Ɛ��cr�� 
�X$B�zi�$Gr��0��gM<��%p���m��?�9��t���:�/���z_y��W�� b�,�*�HT�s�$�V��Z1|믅)n�Ԡ8{=�b�'c��;ڶy��;+���F �C���xf{2�_�!L� ��ڪ/y��Tu^u�ɻ�;��.��3BН�f׳ք^O��^��4����С�4wY�;;�ecq�)-�ݙPtS�t�$5�ͮѝ�t
nΦ�����P�Bܚ�0w"�^$��׽����;tC�#8D��;y!�I�.^ٔq���#8��}h��h�Q=Ļvrj+q��KA�1v�	�xw瀶aì���l��N���� u��s��ykw�����2��h�6sz�0R` ��6,���!pɯd���P�I��^���CkR��Q\7�^�ι����f��Չ��ҟ+d-�R��ޕ����x^�>}�2��y6���of��{`[:���.�e���1��N;���!�G�oc�dJ�r�o�$�µ�Qn����6�=s�?yZfQ1���V�*wLz��er�"&��V�77gp_`g�S����������`��ic�Ctϡ����MK �����0kc�Q�뽳�,u��˿@��w��/���|\g A����Pգ��	mz�a%��*z;�MV���X*&�8����~Ι�m��/��M��@^�d>�3�c�n�-�i�1���+�N�c��`_d'xf�����t����B�ͽV���hg��@ݭ����..�(~\�7Q/�sƑ�Sq8+Ӱ��N��\=���g��+:/��o�c<x�<LQ..�Th���ǈ�ZI{����ی��%�0�,��&H���k�<��;��xB�<�+��j�9y9����.:=���ݫ*�� @�
"XF�*��!�9B����R�K^�eM]�n�+r�Q6��"9�KwlGO�NQzlFr�n�N T����( �l��(d�P��n6��-��'o	n��v��T�"۶�w*n�`�8v��o���l�Ɩ��}�2�͵��OB���!�܉yr��+���+B��vh��Ŵ\��M�[�fJ����!��Zg��5 Y]�
]��|Ě��@W��.�]va��S�nq����j�� ��J�ũ����v��w��O�wz��O�f�wɝ��{�R�h���`y�g-u�1�&�;�%�3���D�p�4����]D�&���2�a�2�������a�Y�������OJQ���3���s�&��]-7_]���j��/);T�dV�n�����oC��0w/c�]�l-^p�&�����%и��F��r�Em	-�&���$�w�6���
dtW�(�9�C��=4Z2X2��x��I�� f�ɈTV��ު!M�'j��g38��_������SB�� #�˭�y��#$S6�eZ���#��U)r�mi%�������M���t��[y	�yޗ��x>F�u����:^[O���j��s�.�"��R���>ן�	ɩeL٪�SY柠wg��_)����,�nb���q�Y��9Y�wb-�E�ӝ/p7�4��6����:zbg�����DU�W�ܯ*�L>�����Ӥ��H�T�ꠤ5������ˏ���짨2�_��ދމ~�eP�8�(�WR�*�/.{U����N��l�XX��5�x�7L����~ *ϵ�-s{�4U�f�c�m�ֽU�<�;ě~�Dw���~g�|�qD>�x��ٝ���������l	��փ*{�wxB�d�&; g\6@٣��^��&ց��d�k#$eO9�Y K�U�(P�X�����Vxf��
�����`6��h���a�n��ڝ+N9yHCuf78^Gw��Zy����y)f���|����C��Ǯ�����[kY}kB67�֢M:�����_nwX�U��ش�73�����oe �
y��W�V�zZ� �Y��%��z��*�@�� r�l8�ư���p^,.�,��:��=3%Ҹ��,���Z#���xE9�\�[\r�Cd�i�l��_�cWEЇ&�����
��ٻdp��r��Q8C+m!	���P����Ǻ8��w�k�=�� .1�LK�5�.�{���ol{$�`�r�{��YY�1�}�x��b.B���穄1gu��C�!S]h��c&N޽���F����{gCwV������I�A��jS��U�5�2:(_�'��4y0���~�:+��P�!Mm�OI���;_`�W[����zpwDf�C=ѳ�+��jzk�|nU#�[*�I�K����s�.��`��Wz-Y1�K!"��_q�D[(� p���_	�y�t�z�3����K�jb5�K=�y;~���,|�H]���\�G���	]C��G3�[!-�,�^ü���i�;%~+}m-�{�s��	�U��pBbu���M�=6�U^���"������x�8|��_+�۠
���(�;QT83�\�6�Ho<�\�ןb:�]�YԔ��;�e���P��W�N����x.�s���f'0$[얙�.(���g�iQ��b�Rucgg9������GT�#)� �Y�+�Nb��p}�J��%'y+��b�ɛg���L�o3���ˮC�u�k�T��?nk��&�;�N���*[m��Q=t�r�n��Oqq�ľ�7}R���q%��X�du��2��&����O�M��6�R�æ����˾��x6͝V�L��$]��W�d##E�`�<�����+���B*��!��ՊX�#Pw�AS�/��<�q�ռ��]�c�r�4��|��'�;T����p�i�b�g���p��L�9�-m0�ޭA��\/��<���GSv��"�\`	>�Qd��F���\u��F�4�O
i�tdK�T���h֕<�3OM�f
p�Ÿ����F�LD�q:I/u�,s6�p8i"�穈�)�C�U�r泦�N!+��7l�㍂?��s$���9>�9<��E��^� U�Y��2�	i��([TAu^Z��S�\Cl �!���U�i��*/��d:�M�e>�Ges����Z�w*�{{2�|�	pB�F��M�*r,���+KGS�*4p_�F�DqƖ��ʞ�As�q�Z�C��!ܲ�g�7��-u�����F�ɍ��% M]Y+^��G�P�S�fx�ue�`󾒂#�
�3%�Ɛ�u��IpJmd��1ς�Ħs�z`�+��^�fӧ\c�[�g"�żd}c j\��bN�*�NZ��3�Y�IطZ�L9���
L����w�vL��]�����Q��{�:2��{��WVO7n+(+�;�Z��g(+T�]�Ls��&e�ݷ)�u�}�=��.�%մx����M;D
$$u�m���V��Q㣸yr��9�*\1�b��Zԕp�j�t��c�(���o��������<�����KT]�+,�P��SĴ�=,*�,�{|�=X5b�B�6�U�錬���xtԤ���띊F��k6IyZ�u# ��U�����0A�XT�k��NsT��:�r�&��W/nT�ͽ����I�L,թ��Rv�	l'e���Q�l
T�&�n���/o�y��x\9���)In'ʷ!/��2K�4>�F��<�:�vE�vZEL�5MM��;�.��U��v��X�Jn�8�Z�7��K����ĭ�tfl�\ �B�&��lv4)��v�����Wl;V�V\��[};e�����H��되�3r��dWI��ʺV`���<Ac��C��u�1����;�����A������y:̈́VH�&넩P�&��> ��:��[g����V�U7!�?����Q���|#���&\�K:�v�uT��)YyD�"UKWu�A#��Fv���!eEg�O�S��_>tmc�j�4��T��(53hv����l�I��3)�喒�096R���P],�xU��J,w�	�;7�j]r���`���d�V�K��Hs�ԡ�[o#�D,�&s�w�Ac0#�GMLзxi͖cqY��:_3W:�r�����+7e:ץ�㩆�=�VГ��;��e�"��ɑF�J�F����.�I�@0�A���������]��t��MY���構�P�����G�Y������4M�E`�F�/ڊ{
��AVs��m�ɶ�b˅0��;��0d��E�8�}ǒ��MJl>ɚi�'q{7(��T��������!�\"�f$�=�g0y��*Dtӵ+���+`��C�&���w=@ �YwP�r��x�?��N�5^��BÞ���-�e_+�m����\���e,����Y�3	�P/�U&�u�f�S�f}�u&*v����p@c��Rp���n�R�[0���:��*��N�V�����٪gn��뢳���(M��3m��Ќ�h]1W$�(v�Sv�e�1 �/	��Ӯ��O5a��wF!�'k۪]+Pr/�6�ˀp�O���yڲ�vN���8����I]l&R�\lX�N��tٚOQ)k��D���k��XPH�=��o"v^f���å�W:��ܰ?:L\��#���r��@��}]h�Sut�v;D�ވt��g��QZ�^K��w���'m^��kv�w�.C�Y�oqK$�����o��JJN� �,̩�-If���n��D�N,�k2�vV��ƝDXD[k����kX�3�6nڛiZÝ��y�gL��G'9֝Y�V��D��ZVYdu���m3d'3� �Z�ô��m���F��-:Im�r�e��YY�Y�MhK�8&h�#��s73]y���B�М�,�v�;l�#�Y��r;l�K����N���Z��ͳ��9��e�mF�&�m��$�3�x��!m���t�Z�$vi^y���,�K���6ٸ�;6�m�۶�m6i��ٵ��&�hX��vf�2�l�e��k�����6�m<۞e�m��Y���,��ز�,L2�KN..-:܎��;s#��:�m�2�s�6Śh!��%"�D � �ao+/l�{�c�Zy"M�W�<xM%�s�iʧY��4��Xٮ�x�Vn��o
�m�>䑄��l�ژd�=�m!�"v�j+sL��!���E?k)THkQ�]�;�����ѵ=U��L�90w�sݕ\�KV��4l��_����h�cxN��3y!ԓ�\���C��Fp����Q�����w"�;��y��0N����Iiθ6D�4�G�'u����dx:�߭=%�@���y�K�}�F����N"@�.��o��4uр�8��2B��ꎽ��?��v�묩�y������)Ix�7��9��wЭ�D�W�~�t�y�V���,}�\�C�;P,��C@����H�N��y��Uh�=.�����mwT�V��
������o�ߌ*�ǛOe:�)&���'{����ɩc^&%hkl<Ӽ-��y���T��}7��� ����+l��0��X?L *(�������рeds�5��'��=[���xiޚ}{깚�T�՝f��f6�� v��bX[C�=7��=��Jw��:��{U��A���`lj��1plR�݉kp��V�Jڄ/�0��-�(A�U92EzT;���q�<����y14�p�VJ���ܬ�u�	�#G�ƺ��ZiT�/���-2�gu[�f�`�a<��%y��Cu��3A�/�o�E��R�4��z\i6�����)�7_]!�Ss@��������<]?k����b�ԣ,s�!`ͤ��Ԧ^k��W{K���x$�m��~�V��l�i=v��sl�P
�DH��U��T��P�9�N�9=	F����ɜ�V����sf�n2�lB0�K)�/M��@W�N U]��fYT�Z�]1�����u�Z[w����{ݪ����"�`p��Tݮ��q��F�XAw�]�,�KneZ����޷�Y����S�J����Ε�7vh��Ŵ\��nܕ�U��S#b��(��z���g���\"��
}��J4]�/��N���тaH�U�b5��fۺ�D�q4�4U�;:UA�~>�GW���k��#���}��<�w�]�j!=�V6DME����:�^��m
d(�$@��@�yh0�d�<2�7���sA�
�YD���an暉�ݪK�m�q��[!8�>����%WK�>儱�{_���g�SY�*~�v�"�묖Uc�^�#�P(��.�w޿2�����yM�@��R8�.6��L�~n�N��!?z{gi�	ɩe��0Z�i����6�z���B����0*gw]��M��T���ç��j����P����ۼ�bƛ[�\Y|�Ԅ.��[x�ӔT�Gƺ���1٠�6�8Tsz]�#hɝ`;�ą���KMp��r��ىwN���ːZs:ޠ�ʆ���(L���X�&����u2�d��RV����k����|w+W�q���u�;�~�����l��ӣ�f�b�*��U��;���rbs�4��`eSs�SJ�q����͓�������oE]Q�y�]3M�����z^����{�S�n�C��ё׮��p�3��Q��j�2��R=O�:-n2I[�e率�2_8[w\����c�\\�ҧ@�ވ� �*���M!3�/Yh���U�U��(g]y.��*O�B�u��:��/�m��Z� �������%��t����}��wPUj�5�l7zn:1��R�qTp���W��M�"��Dp��!��zD�A���{�0Q#��y�hǁ�ύ3TK�&�Z\�AW<�l�Mܩ�P�!����7�Zb质�qq]�K�p�͆8 i�v{#��!!S\��Ӕ��}���m����a���_aM_%'�;�ki�����z�;9T!�<0Y.�á!M1���&G�㚕��6Ee<�7��?doM��FC�ݝ0�]UI滦GE5�wr��9�d��>���p]h�g��(}�d�)x���*�P��\9;z��Z4i��Cl����XI^�79�ĉ��Ry��r��tB*�@6�kq��{sSu���ع�>��1[�
�Q�)gp�ں�$v����yU�jݞX��n4���Z���{7��9�l1��^�1I%����H�n���tl������
d�ʤr�ܲ�h�7�Y���'�v�/Q��c^{�3D�^<2�v� p�- {�'���C�B��d:6h.��Vgv�^�ގO��Ј�����k��h�N�@bWH��&|\��4�����Ѽ�q3w4�i��:����ގ����o�<���\>'���ou�Y�o�����˥sK��Qw�)luȒ5��[%��� [%r��m�i��!`���R����ֈ' O��٪���D�q�>�&i�6/�%��\��Ȉ<��Q�ז/������k�������q�a.���2p#��gL���gU��묑vܤ8��� �f��P�}��t��__��K�r=�Ɂ�����l��h1;����}�3ϧ6i�u�c�-��mL���ԋt�7rr#ę=O<�
Bz��)�'{[,-�z�{��p������n�8�V��.������X�Wg���Й�UjpJ��8�
f����~5����=Mҧ�B��~���˓9�r�t9�z8�S�5iÂl��h������J��.����Jŵ(o:=c0q�9��B�,U�fL��A[����W��#ri��5}��U�q�gSB�B&5@����7�=�!�iS�9N4,,��"�u���9����h�[����u����0��;�H�d7���n�@^�C�	�b8�Aܭl�r�:%����wt��ΦFED�p�D���rzMk�Ӓ]^���y�� 0�,��fYSH��LG9B� �Y��5<�sc;?Ws�YW�����n@*2�d:а�|>����q`-kR��Ezw�g�,�AηkKXH��6&8lޖ�#(L�s�Ԩണx"1���k��+�=4���ㅦB1��;�@3�4�D�2&�R�<��sa���N�z�[�)THkfQ�]���^��h�n���
d!�85��ƫ3bVv!���<;�p�CϣL�l��������q�����WwSk;��n5[Ņ�Q���h�����l��������ͳd:ym;��A��
�uͳD�Z�On"�޷�E6;�wZ��W]�$"�Lk�[9"�B�M���\�I54n��O�1U��(t��v�.#�y�S~�t%}�%t���,}���o�+H����ku�'n��n��5,i�UZ-�
�~�M}��7�a�7��U7�W������st*w�}oU`�����L����Ҷ��N�.4ƃit��^6�f@7����d
��E�ͻ���N��x�h��_Q�F<����f-�v<�q�P��N�U�#Wڨǔ4̧gzqz��J�8�����_]R��RW^�;�q��l)0j�[I'I1H�酀`���'͓R�D����a��~Ι�}R�M�M��@�m���2`\�-�p�:�1���#^����vK'0ee�'�8&މ���ܽ*���b�;=M�B�Y�螜�h����O�q8+ң�l���:����g�2��I���n�G��[��2�"��dswǯv��"�\`o�[0�ʽo���ڏ�:�`[�o�Ԕ�>EMT)G���z����#��o��Ƕ��7jʇ6̮P �C��Z�#��	��!����W<�7�-Mn���v]ᛱLp�d��ض�e9�S�^�����S�Dxg�,��4Ò�����W�}���S�܆��9'E��!��z����"���׻�7m�)�z#!V��
(wa�}�7��_N������.%�Y0�1T[P�*�+�Ǿ[Ԉ���2�{���W;�֭��ڢ���wdEn�/��m�~T �ǜvy�S���_M�ze(�{Q�E��7 ��n��d����f��F�cU���@ᶡ��W���@Y��*������������ߘ9�gTq��GoMu�����-�ír+�L#�����ss7BYҞֈ�3L熵֘���ŹN�]���Zv�j]�рb�J���n*d�^Ibu]tˤKײ�츋غ�̩\�\0!]���c^�v��]���"��T�%�[x��M;�;��4��NN�h�B5�
n�w�����hS!G! r�r!�lÂ����.��FQę|��Izt�̴ҁˠ�����:��㼳w]s��z!��`�	}�u��,q��-ӹ=S��G4�0d��0�c�v��@�]��hN;�oK�y�6� �k���Ԉ#`r�r��5���Ot��6G`�l��T͛�P��i����kǪ_8���R�l�.��K�f;����y#�g�׽�5����C��gО�&i��3�m���!z�+�k>v��U,��}�����?wd����K��k�T�����@d^���Z�����X&J�U�E�f��G��LD:�����UԽy�3-D��>��뮞7
1pϾ᫵N�Ծ͝�w���s)
9�uB����>u���*t}�t�`�2�2#vk9~2\Bm�֊[{��϶9����w'��p����GT��[e�(�ڼ������v����Fe���LE�j��?�`�b�s�c�>2]+���n���p{�ݦ�7B�aiu���|_wJ����*��r��<�V��n=�*���l��>�U�4g�Y��,��C�!2��(�|���Ak������)<{�[\ӿ�<�78�ln��|�Γ&QUե�o��[�f���8��+�P�L�t�����Aϊ���_��2��0��f�M3gSS�x�
��=ʛ��_F�ݱ�ӽ�ͪj����`r���\�+��� ��8��4�$*b���r���o��9�*WU֋�x�:[ͭGc�ͪu�3.����r���Ub�d���H@֍j�b����H�f������u��%�G{��)����{�dtS5�wr����%�|��0����a���nǺ�ܱ��D���tl��wT>ק��@Q '�U#�X�[��[!ň8ɧ.�"39���/7�����q;<AQ@�m��+�8�-�7���@9�I>���YGn,�"3����/��H�ƕ�d.�����T����Ds>��	lmڂ�R�08�-̶�9{��s��̍ʃk�����b�o�.~_B�/	>V>x�C�P��Z�FhE�SV+[��n����c��%�*��m��?g���S��)�,��)���5)�mY�a�f2�M�=A�1[ًM��#������Oѱ}�/�Ǜ)���DA���E�e^���^��Uu�G���[�+7��B�mC9�e�X�SY�/�Ɋ�]���'�-��B��TS�P9,��m���`�ps
�[�Q�E�K�RJ�2�
�3�6��zԡcW6ffF{���ڍ�1����P�g_{�Lư4gwZ�\�֤a��q+AK�N�-;%��:e`%C�pY�<�m���kˮ�E��ź�H������PW���2��햆�nI�c��,`L�v#w�|;��<�sf�=J:�1�l��s^�{l��6)�s<D�pu����.F< ���N�ki��ѽZ�=�AT�[GT���uA���Mޞ�&�Fm"K��Fی��'�x�%8��~CǮ�c���@t�u4l��Э�9�Nh�壢ﰗ��)�]�jTj"| �x��i�]�,.:_�ٙ���K�t���f�M��H���<vy��OR~"�NIu�P�� T����,��!!M1�w��40=�m�£/xmΛ�Z:^ynսv��l�C�'���ע0L֥�ʊh�̰��k]{�+�r�4�5A�BX�U�J�a!���X�nΨ|��As�q�Zhr���ح�X��/f@�=�K��=l�ˋ݆����O��U��6�FwA�+���i���K�IݺOs�˪�66�D��;y��U<;�g�Z5N���}y!ԓ�\���C���������i�V?D����2��z�^��}%*�`�,��v������,��yzs�4��LGc��Q�[z���0�L�3Pq�e<問Ǔ�aN�0otօ�sEE�,����Vw<�Q����w��7�})n19E�����ݱq���z��/�h}�vz�_���\���Z������5�����Av���{�O~Nm��Xٳ�v���"9�W<�����a^���7�rd��#�k��3�wUz'm��6���6�o7��z<]��q�\���l�ynS}P��q�f:�|�L#-��|�4���}z�����`����0�y��E�
�~�^��w]�/��/�����5�.y�n:�n��Ƹ��#�W��Fkh�j�����d���a���[��K�}6L�6k����[o��{��"�X�����y���L�����z����O5���\����"_��߯�N��O��ʛ�Ѡnډar��'�M��Q�z? �g��߷�C�|����Y�[���mԣL[����q�mA�q�-���0�u��@��� ;�,)�T$�X��Ia��sg��iS�r����c�I�U�9*� $[�e^�D}"�7�,[�.�t��������G�f�.�:!JVBiFS�S�^���@]P� ��t�yس\���O9Q�u�U3x�]J=Õ�je�J������ƻ[ӕ�Kq���3[҆<�
n�;�Ӽ�,�ə6 1���QL�8�#�<��hʒ�����Gs�۲��kH�d�*z��ԦI�9��ݣ����#$=�O����Ι}E kp��tS�[6l�[KX���v����zd8;��)F<˵0�ۗ�X��'a�0���� v䏜�J�+���:���`���D̑�%51p\im[cVTD��K��}�=�F�yG�3ћT��;gCN�W6$��N�.�5j���i�C]N&%v�������G:�\��ɚF��sh�S���m,�;$�`#����ˬ�����PV�6,©�\�I�ʮ6g,��8�`*��s����ݷ�I���u���F�����Á��6,Պe�鑮��+^5����dv1�&����vD�	��������s\�,p��K
y�Q)���RQ��\&LJ����_sD�xS���k�����V���}oh�*̗C�C��0S1�)���%�a۾����yvi_R�a��a�X�v�fQﲂt�r�q�Ō���󤵜��Ӛ�B�;�&P�*H3����"%)�p���/���T�#�J��}���K�Z��)�v�~T/9�A3J6���ZظV^�V����u3)��'�;"R�>r3��u5P��f��e��xqn�o�u�4.�^;M��6��y�f�h�ҍ#�v�����IÄm�� ���=A��h���;�!�0�
���M��v�gH���KYz���KXфr���u2��'�<��Q�S�ם۠"���Y��}�h5\e����7�
�s��:1/-��-���'eHf�0�y/:�����t�f$���'}W�"X񜾨��ku+#�Ĺ�/B��X���i%Z]0�-|k�����M����iU崍��a�1��&��Yߗ!�?= `�/���Ē�vy;��m��{J�,@m��m�U�9�r�CD�q=�r<ʲ�l u޶��v�0<��R��Xss���(mBr�ۡs�#�2.��b��xS����@��[Q`b9��+��y��A̓��XNe��%�@�»4k6s�n��ދ]5X�X1���N�B�L
�����AXdB�u�V )d��.��p�͔�gk3����f�d�����qe\#S0�ɱ^���չ�Wo�لlW�nX��b{�s��v�q�˻����]wMq]��l�RR_&��9>��u��*���>����[e:X�M��rޣ���f�\�b��htC�ׄk��Lwƀ�A;��v���#�5V��t�$��y��x���Z�ɽz܉��ͨ�6�]�Rp�B���P��R�U�=ڙ��nQ�&�wer�u�K�P6���^�u:�[}!���r��r��Z��
Z��j�n�.�$j,E}��^^i`́͞��;�� �(��$� ��E�X͙g6����vxkki(�̎9m����ܜtvn���nS2[Drl��ge�Y�ǋ�5�k���6���h˲rl[f�-����63g6����βlSYc���a���<����l�6s`f�mx��c���ͣkl)�MfͷiH���F�hvŨm3nib���f�:�y��`Rcu���-vp��ݛkm�q��v7kf�Kh�����i�٭m��mi�b�mևYֶ��kq6�dm�o<�y۶Q3Y�[qf��C�$<��M6�j9mbF�q�C@�n�l��s,��6�ͼ<ݼ��Jح62v�δۧ;�G�x㤳�y�x��tvqe�]���ѶK2Y�6��5��l�y�I�}�~}}��Yj,n�&�a�Z�S��M�ݬ�8�P��7����L�l­��rLe��M�)�������$ō9y�v�c�LF�ji���ڄ�oU�ވ�&�l^�Tݶ�s�[h�p���Fz�!{���~�A���PŮ%�j�j���mB��eJ���oR#8��{�\0�I��ܷ:������Z\r!�!r4W��ʦ]�,���S���E:}e(�{Q�E��c-y$kϕC��`���v��ؕ4h�ꮦ��tH�h;?&���w���E8c�WA��f�&Y2�R٥�-�wEV檉���n��౸F�M�Ӯ㫩�(����Pㄎ#�H_���c�ڝ_W�}�☔��{$�naC�^�P5.�㯄��O�쿁��%WK�>�D���V�^�����;�t�����H�'�N�@$.o.�w޴'���?(��2��Oe�>�7fA51q����	���êZ�3�>���/CU�6�vri�����h�K���D��x���ҭ�m�:���Q9�\�g��T�=4���=�6Lӧ�&{m�K�@��fz�̛Ы6�����M=V"���i�L��e}Ѥe����AHk�O�n�?(�������h����_f_Brr�B]��;�Ӻ�V�9dy�Ma�������(HDUǼ�{���6��j6�To�=	e�*��w*���8�r��*�[8�!�� �����φ;B�A:�,=SS�H�X�7�o	/L�eJ�M:�sՂM|�d�i���㛔��oD�A�l��]yr�m�t�f�%�d����x��ƨ��!��\r�DѻS��b��gPpa=�>���ͽ�����N����9��A�U]��g����3���7���L���g�lR�OI���Sθ[4uK^Y[e�j��^��"Y��SF�ƃ�*-��![� ������ъ�`���Y�)��t
���S�MH��l�����mm�O����DP���0�s. �x�*P�&��MO'U�7��7{rj�����3���'3��i �Y�����\�� 9ƻ�qd'�i�HSLAs��r�2�Տ�!9�9툫�7;w�p:��۲�n�/;����h�SZ�g*�Cx%�Xt$)� �Ѣ3;ܝ�GUƘRj����=�$޿�#.��E�������}�g�u�@�G��:����~Ź�8g��U�h~�\k��U-Df�C�gSwuC�tO�S '�U#�uU��K�_3�7�	Mf�nw�f|�h�DY��tF��ᔓ�� 8��7Dg ��N;�7t�~��D،|������!J�+4���b������,�C5����oM�\]m�]��=+I��=���@��DM��u�DP�/�ZF>B���VtrrU��Nf��BT���/ aXK��"I] ������9`Ϗ'ۘ�glb&8��v������؏��Ȟ�	�t9oŅ��\��5罷h��{�p���}�U�����S&sb��$n��Y��ȞH�u+w�.~_B�/�O���u�>yDր�_}-��t؞|��c��_
i�����bnW!�ߞ6�tle���v��|t�C؊��f���k��	g=��ڦ�^��}4���G�)��\D��ExfK*����=�FT���b�wZ�ku?f��}��;%��`�z]���L�����e�Y"�ȃ�>H������[�9g��o��}&e
�H�~g��d`F �Q�=�ۺg�Ny��[��]�c��X��uL<��;�Nxÿsdc����0O��}���
�m0�ޭA��
���y�k�����*p��20�a/<l6�ɂ;�0�E���9��h2��4͑/ƛ3��z�!���H3<�����K��齃�fߍ�t�^�[PE��@L���e=4�q�P�Ud×2�IJ��fe�W)���?6�(Ol'�^i�O�(�.�h�Wt �ŞY�T�!!W��N��v�2:�Ú�i��Y�Mz�eL�g���Z���aQ^g�����gDr�A��o8l�|t<�����z+��}������[Y|��JΫ{��.}��d��t���ˎ����\���ښ�M�9-őG���{N���[�]m�U�sBol����ꄁ�y�U[���d:�K�ێ�������wr��.��4:�`�C�rF��xL���c4C���AuL�Q�l�oF{����*zi|"�p+1�ZXF`��yȬ�$Ksо�w�s��,�{�����k��R��֣6�F7t����k����1X�۷|���1�K�,s.hwJ����8X!�5N�t�}y!������G2�M�j�ڃyC7YDu�E�Vڕ6к��z�Z�#�6G��%k@��}	�sd:uwqx����θ���չ��c���T���}�B��_[
hW]�ā�X�א�rEH\2l�U�X�V?qXb���-�V:��y5���wW;���/��͔��+�2S�1~� ������:����k&+��;H�`82&[f�V�l*]��C��n��ޗ�T�g A⚼ �+�y��p�N"U:�s	���>T��0W�������3��t�<��|/��/�P���!�N31�m^7|���& ���5���������>ۯ���(�|��0:|D�����_J� ;K7�`~�]B����\����y�������k����I�S�5��.:��s��1� >�%��RoP
�(\���17�\Ue�|.u��e:�뫬��'ٻ�-au������[t��*�u->۽u�a��'M���G��Ħ�_��*l[wF��}���BzoM���9��6Jw�5���@s�Mɡ7&�I��O;���Nt_��ߴ�1�8�ڶ��B�Y�ق�eLӓ$S4�w����煰X�F�\��Q�t��w]��w�*O�J�C�OU�>ߏm'�Օm\���q��/sy���̌zS�5V�Un��Z:F3���ױK�1�0�%VA�e9�9E������8^���F���y;��Z�ƭ#��y��ezb7���zJޡ*[�oL�zc��}�8m7r���:��ݛY�q�E�:^:�H�=!��]����8䡩� ���NU2�|��ܷ�����!�V�ū]FMYE��A�e�Z^����r��xg����)�6���=2�k���q)rr[���^M�z�[	���Ѣ�=J�+��8S5�v~T���d;��Z"��fR�X��A����r�%��&u��2w�s�{�������^�2W(�9�Dه��k��yK(���]��'��?���W��=�
d�K��p�~qք��]s��5�@�g�Vi߲�~φd%8�d�)nuJD�b(���(���P��jF��6U�'���6	2����zTR᧭_EԽ-�#%Н�,ۙp�!X���ỤSh<�����LG �*�u՜8��ދ���])v����(y5O�#��;Ό[{;����C��x�n���g��TB� .�w޴'�����&8y��L�Z^;^�0<��
7=�t��6B�95,�zfo�����9�aƭV�G��W/�� 7�Qq��f}�4��j���}mt0]S�����H��\��mJ��6'�jK�7���ʨ}��IǞ|��1\#m���tSr��|��H˯�:]t���}�_�\~�!ڰ�VOMb��ђk#�z%�g
|�ח/v��t��tK����p"��ЧՉ�9��Η��(Ż�Y�/Pfu�A��ú��if�k��rF�S�k�D]��;܊��z[	;�MsOzT�#Y����̶)w'��}�)�\-��Z��j��]�;�H�~{�[��/:ӄ�B�`�h�{`�i�F�C��'���,�qTp�K�p���M�i�Ț��ڲC��KE6��RR;�L-�R��Ne�������*.�99����q\��uNl͒�(֒tp �6����!��E�B��� :� �Ë!=4�$+�\��Ӕ&�mm3�>h�G��:����3�92�h�ٓ��O6-}mu��6���:��kuō��'ˆ�s�|�_t�
�����'��=�z:��]���ѫoO*-nI��.��F���
�JU�o���*ސwy��(���j��X,������ܞ������b@w�}_k?��/;���� ��;9T�!�<0Y.�á!7�V����ܞ�%��!�7I�׳(��]!���gL>SOU'��t��Z�w*��ب�g{:�D��1����B"˝yr�Lg������q���P��2�	泯��<<b�M1Y��A�8u�-�lsͳ�"��,bv��8p�=�q��M�-����vU4tuf�qĈ~�2�W��C�o�/Ѽ%�T�p�̀�t�T�WP���*q�E��ٝe}&�l����4�t��yd�z 1���mm[��m*;�d'�fΛ~pƟ;��7W|ٴ�cjib9B:�v]DSwG;�Zӂ��%�}��{v�k�z�(z������{^����]i,����jKבSZ/
��}4���/�y����g" ���)�d��5��o˙�&���a�LWj������禃3�-��w��3���i�]d��R`�F�4E�ԙr�\arq��Ss8*F�1�=vC ��w^�������j�7�W	�W�ݛ���a� 3��� ��5r&�֋�7���A�\�ec��ג��l:i�qc�M�ǗRً���
�(�z<]��v��ۇY+x�Vj�Z�=�&���xx9�I"G�!º��*S������S���k��wr�ƌ�x������?#�4m��{��.��.F=4�~1X�Z�`7�Pgւ�p��捭˶���Mw�[��n��ʎ�յ_�� ���q�A�ӑ$SJ�@�D��L�ٶ�%`�Q�{J��{��i�+�d���8CSw-�"�\'uB��S�F3J�r�q�x��|uJ�^U��O.�"_����7��O��?jrK�m!
n�@L!�<2�i�P�HD[Y��*	��V���s��Q	���U���+d:�L��}�Ges��SZ�w*7rC`��t��JN�/��ϦXK=�"�"8w	�])S�Q��``5�Ψ|���AI�u���#mlgu8*t�";!����w��?t����h�8+b��-�B�C��3����46m�e�s�^T���3���B^�L����Ɲ��K��5^29�﯇ i�xn5N�Jټ$�\��b1�Υ��}t�����͑���Џ��GeD�B~��k�uyx�o7��z����T={�I��s���M����SB��$"�Lk���-��)�^�m�[��~o{݋������5��^�����K�8]r_.��m��މ���e����O2:�|��o*\f��ɇn�%Qh�Q�CnK��{���X8�U�5@,�'6�{)�w�P�&�f���{�Z�T�2�r�[/P�� �nig��i���?��ƒN2��w�O������}~B%�)�}�o�)�E8��fX N�VLqp%-�3\�9�I�M!`���dL2�ު�xT��
f��wM�R�[��*�o�b��5?<69S�$�������ù*�*� 8$'�i5�'�5���m�3���U4��B��n:�q�>�Z��S�ﾀ..��C�F:���kԨ�3wƾ�d�V[�쇃C��ؔ��G	Ǯ$w���7�ܾu\��ZN�|���|~_�Q�	]-��]q�Y;�b2�IhEÉ�i�V����ߴ�x�z�rڒ-\`m�%����&H{������!k�j4�S�;��)�w��.��
8�0���5d�Xna���B筽�M]O�p�E�0g�zDa�θVDs��.�qL!�K�r��6�r�ױ�
����8BsC�$�}��p��3�[t��*�oϼn����[�ޘ�[v����MۚN���u�st�/��	���p�5����3��9(h ���
r�R�|{�-�Dt*�����t2�>���+���=aw^l̺����)Dڱ��´Θ/:�N��S( �i;���#o�Ǩ3:�@�C�T��Q���0v&��|^��2�����6�sA�ٱM�PtI�s4DF<��-��[�0%�a�}vlW;eFupz��[��sm�f����m[M�g�qm#�5��r�Aw�p�;�0�<"�6���n�2x��f�+j���8wL����Ϲ�'@�Φ���T�]�#�z�;?*fxw/d�φ��x�|Q�Y��y�����5W����/~Q��;�F�^���z����hS!E{�P��F��[˶�
�j�jiG�"&��n�xb���ḝ����K���8��	�y��Ц�!�_t[���qVm��16�1�_���K�"�c`X%��N���H\��s!8�ٗ���э�;m=��j���ͺ�:`p:����Ѹ1�ҹ���15^ʛ��5yާ�2�bzދh�w�S�mKl����+�MK�2��ZH���_vz>�k��ߔ��j�&<�G-�o��N���n��[��nF_�*�+�m�SN��yV��& g=CAǌ�ʽ7<EJ�q��+�gQw[Q9�j��x*|~�R^��eV8&t-��1m��^]yr�|�@ݾ�aa�!���w��Y�xzk	�2�^��c�,�9��l��A���S�n��s܍c�vNH�b�@ۆ���^��i6RL�-?�.�X��2��eU����j^�h�ھ��k˽�Cت	����w,���j�,)��$$��{Y��Z(%�fv*�}�ϳuu��=1�4�;�Mgn�:�� 4F���T��z�	$OZH������9���n?�%�'s�/�f4�E��Wz:WL�m��=��iݘ�aP�aL��[6*
�u�֊�ڛ�n���&�<��rGR]�����`�0���"l�y ��]k��]��C����9�\W!����P�ֲ.U���Rw=E���CԖ��f��M��'�8�M����S�oYˣS$P�a,�N�l��u��,g!u���0�'�����늭Y�_]m�xPR9:e*F��c�̦�g<�| �B�/��N@��wf]���ܱ>u��]�$�I�ͤ0Ց(�v&�yG�.���qZk�v�"��vWs��҄���b�7xe����v��:'YS]�%�Y��W0L��-�M�M�v<i���*mDeֽ�6���t@���һy����4� B���"FMq|Q��D�m�X,R.Cm[{�KƗ
2��C3�q������}%^�z%����*}�;8Y�Qe }�9Z�jC=t�׷���3���Un�7MΝ���n�ƞ�l-K�ٱK�X�r���C.���\(�@�j9Oqu�G�6M�q|\�T콕-�@�w�%��
���+1���V�5r�Q�p�ev���n�ɉ���SY�[;�N�芀pj=�������J�N��S2�W,`�8X��H�CŻ�8D���������E�72�-������Yi��6-�>���9�N�^�r� ����on����g�kp��n�f'�6��+!�|r	�x@�Í�p
�[��S���W̀q4aŕ�uq�=1�Q ��T�ޭv�;2F����e!��o%Ӳ�V�%�97/�
�>�2c3���;C�L
�f��+�G��m����ie^'�p!+����ˮ1X��K�}Ǧ�4�֗"Ģ�(�^����i��́��،�"z��W���Gw���#�5dW��4��9O�'�X��a��/�U�t����W.mw@-���I[��L��|��.�q�EǸjR��^麺�bùC�vI��t�,�9���U�f�)k��%��c��gYP���%�m(192�<3r�˹/��WdZ;?d3��)E�����y�fwG.� ]��Ö��=,��EP)u�����Rx�e���*m���ح�L�n���d�t4��tNH@8�#���YJhthj�c�Ej�V��x�te��̩�%g0�� J�:n�n��������������d8Q5"���-���mQV{L�;���5o2�Ѿ����i�ꓫ��������t����	�(�'v��z��Ҿ�����a�$����fK�Ym�����,�"��n����6�ٱ�wmhM7�yxh��-���m�m����4%����݌�F��t#�ݭm�E��۬�Cl�ff���em�f�u���s��L�a��p�ٖ�9�ҳN��Kqٵ��v�0j�X۝��`M�-��l�6��ɺ�-7�&e��kY	��̱ikm���hv��۝��Gm�ӛmm�ܱ�ƶ��,�fH̔њ�ͬ����n7l�sZ6�l�m�ZŷZm���Nj�fݬ6MFC8�f�����hśi�d��,�-���935��8�ҙ��45��ͳ����45�3dɅ��Zۍ��m�X�6��l�,�@Jm&Ȗ�79��ihlф�mJm��fm�ֶ�j�ݣ�[6[�����'cV�c;a��LI	(H"�QD�)'&�nvyol曁�ģ���=�)��{Uw�R��N	\���Ԫo`�b�n�S�u;�*u�&����dy�|X���>�l6}�ɜ�9"�&s8�������RזV�u�2�Y�� I��I%�����D[ܳ�k�4�q��J�F+�4إ���L�J�e�ʶ;A��/�w]��ۜ�Nh�r��8[7Z��P�s-�Bz�2^�c��j��KK�����ާ�Ϋ�F��u��@#;�ʛ��N��E�B�� :�Aw�qd'�i{��þ��,������`���ss8�SԎ�5�|�9���i�$�`�wWSu����z�;9T!�<��cj�u7�f�^i�Ղ ��U����r.8�+�>M������^��jܨ��)���Z##;f�H�>������q��)�.YS�$Z���tl���ڞ��z��"pY�j*��^r%�����#z-�w-�V�<ێ"Z�ᔓ��[(� p���3�A��� VQ����@X��͡P�L
�2	�c�~,[��]����F��s����ו���N�������Ke:��a�}�#k�#���1K}��ʧ��.��>�C��ǵm��e�~�O+����WQ�3v?yS��W#�oUߊ��Cw�I��{�.��yQR�����$�γ/���DGU�V;U �%��&6�zg;94��3{vu'26�ܴ����o`��a2�9�W�����7{Q�m�:=��salӣ�9:fޱ��:Z�9~⪡��K�E{�9�zЦ��pόܮ�����h7T��
O ]�9�����l��/�.n����5%�Q8,�?���ضn��<�MU�3�i�E�i��饝����Ea�2���Q���y ��<"ϯr��?}�m�3�ٳ��WT܊�쎥W툈�T���@���K0���i������3�dY������8wDs�˽U�L�{gg�<dt�{]�k�r�6�K#�z�5��t��ܮ ��t_�^��2p);p޼�y8I6�ף�jS�绨�j�[PB�`$[�q���Ȓ+ҡ�4��y'ڔЎ�n���3D([�KG3��#Mҧ�B�OM�Qd7qɍ	�\ ��D�A����)xg�=�|�b��:�Ҥ��;���0��M�i�p��o�S�OR~"��W��!]Ѐ	�{asC����H���ӵͼ�"/D�xmDT̵U�3-��e�l�Z)�O���~��!v�w݂ѹ1�s��;���v�����"\.��*M�d�x"1���k���n4�]s�-���-D�++1@��`X�n���N�O�1�F̱�)�b�T���;��
y���_n�d�W�I��ye���VܐuF��֕�M�z1β�yM�ڗ��F*Yl���2�+sdgB��O�ڼ޲�q��8�o*�)Pp\�֣��[�����=�x�E_49
��a�K<����^pV�5�[�)THke��(�3�.�K$`��Cf��;����B\(��7&�~L�:���S�&��s-y!׏=;sKF�E3�����5����8�B�#8
n���Ϯ���"y"=���h4zdOK�kʪ��Z����{����p�?%�@�n��օ6;���aM
�T�8��������̙���5��1W�GzB��Y,�N+����@�k*y�Wus���d"_+�͔�,ܦ�"[[:�aXݕ&cL�j��q*9��?T��
i���\L2����T���q���R���:�I�-�k�/*�t�'o��8�ň�*�g���f�8�S �M��ɩe^&'�5�a��E���v�j��~�-[�{�Ze[��7ƥ����..����ϑ��b��ң ��N���d�+���S[��[3ǎ�����kx^�O2�����}����ZN�W�����t�8W���ޛwZ��RrK&x�{&���.�N�g�2����ߴ�1�8�����W��cd��=R���"i[mF��P�g��GӐ���	]�ȾC;�v:�աc����x\*���%&F %�,��)t�|e��ZSY^�t���}�O��镯�<���u=��j:`�X4��r�iS������D��<����owM4Snw6��i�}E�<�س;�f]�%�����v�1H��C��=�s�Ҟws>�.�J��!G!�4�[���O^�YP��� !��Gf�GgBl�H�C�)l��*G3�)�#��b�s�!�%,V��Q���NQq��k:��k�Gf�/�sm�8TAw�3ٖꘂa��zJBT��ޖ��"�����@��|宲��i�y�{�sA���
�d8U����g䡱� ���NU2�|��g3��,��螜��X6:�q00�-��U�X�r�T�2{�q6W�uw��+�6'!چ���ʌ���%�S��2�h��gQ}��gSF�i�T�]�#�Z�g�L����w�����9Z/�qA��Z���v���[R4^�FN����7wN��G_[Ez�QM�(B$��_[��:j�}(
餑~}�8�<�.��g�(M��)'k�%�\w<[��	�yf��4����l��;���7��鑜��c]��w����n�B��W�om�
�0���.[{j�]DD�@\ݬa�F�u���CU���1����zQۯ\߮ѩ�u�?�-�G�+	>�����gQ��Id�	�뚚��۪ʲ6�&���%����+�O�<�v�H���������d|EJ]{%7a��wX& �7ut�&pOz$4��0+�r7;xhF6 ���=B��N
}Z�[��aim��e��#d��ķdF9�mwT�W��DnW-���:�M0pc�J�ᷰ�ϔjaD���Z���F����|~e������DW���F�u4�W�om�& e7��L�T����&{�`�Zk������st���6N�z�=X�ؙ��މ~�5u���(�38C
.�v�9�����	2o�y�L�^��Y<��}��Pfu�A�����{A�r5�M���4>�u�X2bfE1�� ,q���!KuNL�	���	��{bzO
9�F��<|\k?V���~7�O ��^HA_�-�Y�#]@a�[��V)g�U!�����&q#�񓜉���zM�q�ӄSwB�/�Hp�E9�Bzi�%���֞��gAvKѽ���1��Ig����ͳv���ʛ���p�Z�� ����,��1	������93[6�v��/U�SO�Su.�~N9쀆wd���]M��.B]캹�*�+��?��L�*-��N��њ+���]T10v����O�ˤ>��{=T�+��#�Msa�u��5E�(Y����
�z1�u�C�)m,��hV�k�L��y�Ӥ�K1�yi��o;{������kk�;u�us]��$�;0e�_3w-�HQ����hmE;�LW�2��֦#R�3���3��f��i����,�Z-�`����!���Y|�軈E���*0{5I�_���#J=5w�����Lu�3�H��9n��q�����ԖxR6��!�M�#���2�.�	E��a�l�KD��6�8������@�Y��M���
�:�l�%�V��'�t���S= ���<K쳨����9�.�j#��=ߛ1-�g�kB�ߑۛ�n)L��h!m�Ͻl��4�.���>nW=��~7�x�h���ǹQ�&�Rmh��ș��J�n��ȧ��"j��ʗ�n��}�fB�pSo6K<�+��>�r���
�qQ����+ci���LW:G`����5)螚�xz_�_D�(���1�]�K���ė!w�GޅOh���ׇ8��xC�
��i�X+���	��������x���o��F���/{#��m,Z���FC�M� �a���73���-�=��@�����8&9t���;�7q��]�-0��r귛�f5W��t�"��_汘/��r�|�mѻ�t��8��li���Λ�+��~�ip�����ŻV�j� ^��(��\W��߾z��Wz�:���v	o�R ����X8�G����V(%M�Ҳ����\����Sym~�X�R�d%\�M��: a�����[ۜ�g]�`�cJ�}����������9nk���puM���Sݴ�
4��I̥G5$5E,#�׸��"u%����>��{Wy��G��r�)�zm���!���j�W ��5"�:g Fv��[���i��G4�;��ɇNi�M<��%p��Oښz���$���r��@Hj��}�t1�A��HLY�a����i�NP���i� v,�8�)��;+��>�k��Bwl�`gk�y�E�Z^:��lR��`9w�=�a,�	
�.U�2�G�����ʹ�)�f�Yr�su��}��]��`�w=Hq��!��0w�T�r�־�~�*�͛Py��(�x=�x�F�f�F�]�M]U\%�ЦBܚ�X@r��A��=����48�8{��͝��K���Rr�8����3�����hZ�>�WK�����mP@hԅ���ӌ�Cd�[H�ޭ���1ٙ��-�!��i�P�t97�}�B����T*��M$#,���h#��(������搐ɬ�X':�={I��L�T��w�Ő�|���g���8v�7�ף_{{��ۉ|��yg�:�u��!�;H��MK*�oUh�*]�z���o'ᓋ&d&���ێ���q{e�mX��o"��ɢj�ɮnK]]_(q�@,�4��+����*�n���K�79[`���|��k\��N�]����o�^b�`ˆ��Ŋ�221E����iT���ѝ�}V�ufI�fY���l\���:7%���O����Ӑ �e<����1�&����c�^����H�[�q�y^��v����ݏM�F����}R�M��|-�� \]{���Pz����t��2��׋)��ޠl�kX�fAVt��6?E��`�Np��o6�[���ʛ��D��B|�����H�Q�7�9u�^ָ��w���p�N�g�2������0�znյZ���tKf�̽|2������sQ�<�ޕ2E3Nÿl���qK����Q�qS�o���=����eC������&KNK�(�� P88B�0��9C �;�]��B+�K�r��#2�a�D�9	��l�˙(�=/�J����8��[��d�=%�!-��-�
GJ�YMX�f�h���v8p��"�\�"�!V��
� �Ǟท�5LA=��W��X*�;���w3�zK��z~��\F{��4e7uW��r8W�4;�L �������-�Z�F榢״{p���ͺz�F�ڌ�/��'@�7gSF���M��#�5�v~L��y���U���KA�}�trq�HZ��5^+�F���sb�ا�-�ԉս�us�N��`	�����m���Z5�U���ZJO/�y腩/��oBw(�62��XNqw2�����U�d��h����Z� �pmn����
~���nl�KTf�=.G/���1�t��/�}��B�xw8ǰ;��]飯��(�����,���-ߊ�rOq^�>��tI�'���\%�<2�'k�R]%�_	��hN;�ޗ\�zcn&��B�W��oS���g�g�X�C�t��c7�m���w&H�ap3v��uu���n�Zj��î);�sp�w��{�S�h5#���å����8��\v��+-yVUFë���h�9C�s7n������h�K�7���	�r�oϳ��郃�*3���פ��kgS�^��`�۴Ku�s5L��ב��ׅK�E5�W�f�W�o����KA�<^J�Dl�ie�MU���䙿�����E߬��>��*�œ=���-�:-��^\�߹N���WƷ������N�����^���M#x^�N����3:��A���ۺ�[6��nnla��"�"�v���Fnխ�=g����<7�"U���[Mf]�T��K!Nì4dҞ�7��\�������m���9 ��\1�O�z�8�B�-��)gGmjU�)SC�d��pc��\xb0M�w�ܮ��*a=
U�Aʺ��]�tQ�)�K]�<,d���dP��-O�\��@e۔Vk��Y�W*ls*h,����'�R�M����=�J`	���Άl��p��n0�i��BFef�y"�����Zm����ep9���aN���`8)�S�pB{�2^�c��O�vo,�b��7�[��S��;MO=�usͷl�]ʛ���p�V�.B�ЀB�38��5Zս&��ȣ��V��c����\��}���ol|ݒ^0W����ٴ\�-g*-�8��Hܘ��L��_�U��(n�y Ts?_�Y\k��׶1���e�������Rxn&:s_M��aO�4ɘ���GoC��hD3�gm�3�X�.YQ��E����gF�8�B�����#.Ul�]}ȁ�C��f��� �ĪG�,s�e�Z ��y��~����������k����9]��c�m�qߺ+�>4)��Md:,!��o	z��B�|�9w��3��\�[���^�>����\WP��s>qd%��C�w��s�*�~7�v�jܬ{m�v|����v��Kev�w��<�я��fܽ3i5P�eK�E7ts���!M0��Q�u���/�c#��ʳ�ۂ��8���A��I�R���|y�MJzbzkF���.�#��_i�6SV�4��^��x��[�䚿�:���'2�"i6kv�uI�ͽ=�E�$�dJMxv��v�Y�V�^dr%h��3Fc3�Edkz
<��Q��}���.]�30C؛�r�oU�ح��_���j��_S�d�M"���~If��@xw��2[��Jt��.]��5�Fe5E1P̐����@�
��/f��=�w�XY�%�g(��}��Ҕt��۱܈�Q<���;�;�N8b�j7w���{n����qw��T�����w1�,t�� s^nJ�"��W��H�+ �m�WB�:�	'h�x[zpP(���N�ͷ�Kt��6�m�W1a[m"�I��/��NY��)�]�ˮOw�,k~Y#���s(Tn����f~^�y��4�Y~GJ�	.*ϱm��Z�#Ua�N���er�)�N��»)�vD��s��V��Z-���X��*.VMOw{�H�Y��Y]%�W����;�2%t�^�������k�\�J^7-�7�����r0\�Ek�+�g�n�UZ�2���Re�3RN�l��hj�����5+KB���da�e��4��ẇ����R�_l����I��h�	��mu��3k��1n,�J��:^"��@�
�*m٣\���?��8�����o�.��T%���ށ6鎕ΠK�r�;�ui��L���@k�_��S6z�E#2��n����#�;�f��	f�Y;�^˥����ՌV49.�X�`[/_l�jcem�β��	�i`Q�dDh��3t
�Q��:�/�����������ogR"`�/�_�n�!K�R�,��N��%i}:�w�ֵ�!�,�$�PO�bĎ� �����u�"�O:4Ѹb�lgV^��q�j�ҭ����ۗ��ɋ #�0�N���&�X�X
MZv��@m���O8�ݮ8��&y�C���A{���'A�q�hb����V��'����$Ю<v*�"�k��
^�u1�[v�?�c�{��06�{���],��>D��R3Et�-��aͷ�9��7�� �2dV,���
/M9�PisPEfIay%1������Z&�O�����mJ��W8^FFm5ӡ�Z��b���Ihi�9��b�XT�7#JVdZE=q�&�u�۽B�
/jns&A�c�gs+5��,��P�&�7	!h���(	3�UA�ۤ#�1lǔ�U�N��5"fӰ�� 'g)#C?}��z3�GP��^<F�V�,�PV*���gi��$,�4�]\���e���(s}��Y�c�����eK�:m횾j�˗�+0҆�\�:�[�������t
�rە4<t���<�;��|7�=j�E��3������Q>��J�7
9�4��H�I�	]�hvյ{���PK�m�0�Cj9�	��R��'e���J�x�5}ˮ=��i�Y��3bR�wf����<gps�r��E3���m(��Z�	�j��lf�֦�:Hkim�N��4�ٸ�L�31�f�չ-�m�B�Y�3V��`��s$vM�t����m����jڲ���E���dka��L����m�m��1�fێ6�۳M�܋e�G,����ZqIh�@s;p�n�8��A�n�fYm�e�ZSn-���e��f�mh�v#m��6h��4��c7$6�#�v�[P RC�f6�٫2��r��6���!;mm���vn:����m��m�,�t���9�,����Ӷؖ���Y��Z\Z@�N�E��:A	VC�@�kX]�N&q��5�H��]���D�88E6�Yi"�p��������l�
��4�%��9�Q$���5�и�d��@��F$��A�S���{��v�<���y�1#"��f�;�뙢�j����Q.j���Ef��|j`9��פ*������фG���陓�m��4���~@pHO�rvS���d����t�<�'���<���c)a.:\��]d����SW��Pz��zm���nPY����.OPw�E�
�R�t��<H�y��r��w1�|�F�Q�E�.F=4�~1M�;��ܐ-p�3ƀ�̴�FsY$�~�Ը\uO>ot�>�[PE�\`	[tN>W�A�9E��=WXч����|OB��D�ua�w��z�!G.���ߋ��}ܶ��ep�	�I�N-����+GT��1E3Nú����M<�BW	�v�~7=I��e9%ֽ@Be����d���Ni�� [��~��R!p���r����e���lc�u��2�j[8C�K�����qpy9�# T���碠x�ٖ�А�B�l�P]R�G�Q�z�U��l7�N�gjU�=5�[p�q­49r�᝟OCB�*�-�Y��k����{.vw7L����^J���tΖ�ު��ЦB��@}�_��(:��{�s�u�۽��/�I.gWZ�<)�� XQ�m����A=ƌf���l�p��sF^{��]޺~i��9=�p��^;�"��e�`]s�E�0%�ʹ���Ǚ[1\�B̒ ��zˎ��a��-�ҝ�`ᮈ��2�8�NT��g]�4�h�
��p�'Q��׭������G-�#8
�wSk=4u�4T(��7섋��˷k��!Qt�~|yN�;�bo���2�&�Au-�!��N�Cג� w8�|��Sc�uu0�hU]z�t���gﷵ}*5=&�/��E��=�2�p���e�s�S֓5�ʞq�\���OFGtp錙�M&�j�m�~[9���X?rêǮ���>��o�>�'�7��^.�3vA���i�2�opW��3�C�X���kþ��G˖=�V���"a�5���T�Q8��(��n���C#��6t�<��|�o���o(�龙e�#@���!`Xnl����LL截��ñߙ�1z�+-���x_���NoU�zl�ʛ��D��x�����1��#r����䇽,B�s{'��F�q����Y�m���3ǌ�׻V�j� [�k<���ne�.9���-��2zѦ��w3�R�J��7ҧ�垞�|}��I��-�F�b��i�����t��[��ͷ< B���_ ~��񺨗îy�����WT��[����#���;v.�;M��,)!V�eZ�K��J�jP�׎B���fq�
D�V�z�ƚ�N�O�-�����]Z��y҃1�M�u�F�2e�iֵ���iwB�5�7��gr�J�j�c�$ݮ)E���YcM�����.�=-��Us�1p;���հ� ݆S=%jB��V�@���T�윫�&��H����TݨE��-��h�p�Aw�{��\rP��OEUj�r6y��M��哥��WyV�|{�H��vh�n�������r��xg����ɡ�0����A�ރՂ9��hڳ6�锣E�gQ}��:7gSF�f��M�8W�C���r�Y�g�ȕ�f�D|���㋴��^Yo�u���;8F�M�Ӯ�����\�.]�ywI-+B�B@�9�"-�y�FM�2�7�����It�m�q��[�t���T�N�/U9pd�b$�~�7\♗��Ty#�[TK�{_��_q��>��xe-�j�-�3�]qQ� ��'g����OK��x�|m�{,ܦߠSA�{����`��a�|wծ�=w���;q2�o7�t�b���n��=��9�i釾0,;�71[��q������ז��H[��R���}!����)t�L���=/�}�6ۺ�tS7+ʷ�91)�\����,;*[������Im	���1p�X��Hp�W\2a|o!Y-T�89V��S.���/ ��`.�j�S��P�4�gݯ�$3R��R�s�Xi�U�3��R�F���s�%N��20oQݬ;�Xˠ�u���)���nA�>�����1�y�G�»��/��?�XZ�����N�z�*��1�н��3�>j�˗���� �-�24I����D�3tE?|�(c>�=u�>��\���h2�8[7u�h;�[,�A	��
l�ŝ���[��=���Iѹ���7Es�(�9�	�����̶)w�zO���^/6�)�zZ�<���M:��ѵ-yl{l�-N#�=��g��XK�]4��WO�{�����NDE8��5* �n�-��6��z�.���z��0S�SwB�/�j@>��X�@�>��|3�gpn)��;�j���椩im������MNs��y��2�9�N��E�B������~Ã�s\��ѹo	�lk�LE�i��=mSNP�*]X��r��G��c{����E�B�k�|���4�uO;<ۆ�~�9.�6
��Z.�ɓ��lc%��C�������zw�p��6��r����26*���S@r!��g�>���p]h��e�z��#4r�N^ta�L��[��*�MMv��f!D�
d��( ;�fu��,�V�<ۏ����g�Fg�^?��-R�՟3q��Z�7���DZ�͡b�ol��V��i^�V;4������Z+*X�fq�DhW�W)WM��4��%���E�˚5�W��+[5�M����k\��.��ଳEb!i=�&blⲺԪ�5sK����ئ����iR�����25����Q=89�#�_Dg ��N;�t�K����l�vPLmx�ŉ��t/��o=��:�Q�V�an9�`9Kf`1=�@&|\��4��{�ܮz 1���m��xa����6/��V��b��~���4��9�oϤ���P�����օS��o����8�� �S�G�>ku���?��}Tٯ���>�ۚ� qԧ�'��[a�~W�Oѱm��}��Z� ^%L���T��\�g"#��E�C2YS4��
�����짯A���z]��n��˪�͵ve�ii���ݚ|���D9��Q�[���=�0�>��,��Y@ܴB����De�q��7t�>�m귛諘Ǿ[#F�)dc�]5��o�}�ֵþ�1�}��5'wP�w�2Ú4֠�mR�q�<��Ӷ�jڂ-�� ��N>W�A�CF옡ݲɥ��q��7������p�udK�b�w�8�[D(��SOM�Q8Cw+� �� ItIi��AA�$���q�o�1½*ʬ�r�:%����{a?lt�Z9��D�ti�rۛ��l�vtew귮.ՙwa�3$,LM����WuN��-�F��dz;���s�R��>e"�[�z{9��	�U�91v<z%ZT	��|�@$'��W״��w�1�fH2'�)��j���ܔ�������5���傖�wpS����68 ��1g�f[��C=1��DKT����Z��Ln�c-f�U�{�7|����;+]^���wr��.��fXO��!\5����T������	���;|#6��2/ygL=�D�W�~7��8���GA���t{P��2���8<*�2c-^z�yI�Cp���{��ݝM]U\%�L�)�4;�xw0�`��j(jS�&��.2�T[�Y����*���(�C��Fp���K���]/'�7K�#�{͚��@�Y� ^M�	�_�8�8tj&�R�͐��N�C��@��9�z�
lw���a.m�p�L-~�sd�$��\�tH���ז`�rE4��M���u�}&&��<�)����p��W��r�^N���$�<ĶS<��mD%�ѱO����!`��	l��TٽU��= Ó���t�ә1���ΒM��@�1=.�{�񷘆��q����졫G���_�	������J�U��s�<�����y������y�x^t�<o��}����om�..��[:ɋ�k�F\7;R�:3}@��e�l� �"ʕw�][v*[�]�q#gHx��K�+��) �L��V�����A��u�I�C2�p��͒Hn�`��V��,w�c n��/V�s�t�y+�����I����i��g���s����)���ܺƵ��/X�4Y����i�k��M����᯶�81�L3��ofމ�z���U�g�&N�:8�.��� ��� 3-�� �j3�D�4��)��85��N�ju��oj�{�Y��)�63�Mڶ�����|�˘/:˷Q�\�%��n���"w㭓��qC�����iS�rƞ�|}��D�Uv90��֝3����o�r��l2�H�"�Bg(W�"9�b�xc�a��\H��^�]EFk���:q�Y1�vy�E�}�g +��Qݬ�+i�&#��.Um��eMk��5�Sv��p���sfR-�`p��Tݷ��:�E�Bр�0���p\K8䡵t� _k�W����n���j��S�]J��훖�"3�``5�i�)����v�@ᾴ��U0����xQ��ך�ؑ�y�x���f����Z�t��.������t
�gSF�i�T�]�#��|���|��}�����P@pGрήҨWfz����j�Eи���#_ ����t�bN_�qE���n�����dlS.�!l��a��ђ��f�xe$�t
�]%�-����x�;��)���r��\B\�&����|��9��+ޔ �^��o*�	���\
��`Q���E,��Wm_nCq�ٜ�b�z�t�7�.Iʵ��K��^I�1lr奪�[٪+I���e76(�ؿNck2�H9��S0B��(�6w���X߽�_���%V���X�,ζy�c���	�s�%M��@��YT�rs#b�;VUt���$��}��n����}�m� 3��اn|���y�2���f�$�u�ݘ&&N��e4�
n��q���/�`Xw��s'��q����=W�O`9�ji��$�d'���m�_%�f������k���^���}�Ӣ��^U���L@���|u\_@R"����DEsBa�2����*1�VJ~y��OPeV8�=���`�:-�T���Z�vq�%K�2S�n�D��>��t�n������ Y����\�����>p�i��ݘt>�m����hZ��X���C���v��Ĥ,L�"�C/��x9�R�ÖN���ݭ1{ZpޛzGC�A��醫++]a����^HA[)�|����ܪߐ�,�KB]C|O�u�8��4�����<7b��^K�p1�-�X)�+���Ԡ8N%������bͯ���L~n��ݛ���>mNՖP�]{59�����k�ʛ���r�n�@�up�i��l�5����g�fҏ�	t�f����4��Y���Ν{\Ãإ����t��J��TH�e�ö�%���;��F!v��cNN���鵆A�e��9Eҭ�{*=8�Խ䤼���vF.��bLkOfa<��swuցt�!1Wr�;{���4�zi�$W�!9S�eK��<rm�#��vIx�M�]M�*0�rg]d�|����}������#�C��0�,�K����zb�Ue����"���=�"�|�)<5p�Rs_UN���ӵX�^�2:-w*�9K;h\#Z/*o���޲ʞ/lMť���;�<dn2-�Ja󧦸Ez�	�H���3����+c�o�8������E�p�{�����sd��������:������=��-����etͨ���'ݺ��ɞ�W����.���[N�@jb{�p�tG3�'��]AߍG@mb�Ba��øWt�E��IۿT��1�����9��������1�W]������o6K=SH�^�磛�3�ĸΈ�j�:V�A�4��
i���S�ϛ&�9=�p�������.�6�V��a�Nqq��\��t�Dd"� ߨ$k����#����,��!?��{�EE,��|���q�Ύ*g��u[�2묑|�8�z�Dxdc�f���R��&}fh�����R�9�dF����{ZO=�gU��H�Z�8��5��FfR�q<=e�늵����-��J��Cq�@��(PҺ�]��;��X�M�m�]/��L��-_+����q�#yՖf]<��Ż:Z/�z����ά��Ji�6��FDn��ϼ���=�����{~���x����;䈺���Mc0zlŝ���`^ڸ�Ei�O��q�C��i�ƪ��
���Sϛ��p5v��!P���xP�8�B7c+*�B��g�	~iQ$T�?M�.�b�w�8�[E���вzm��2����T����/>�ƞ�8I�� _j�":Kצ!;��ɇ.s�\��O{�S��O�%#K�^�i���}TN�����E�"�� xCxafYT�O0���u]S-UoL�1�Z�+�J���d����[��prG{V�>�vW?[6��Z�w**w�{2��$1�A��.�_cXn��n+k�0:hsv��cq���vuC�OM ��E��Mi��@;�W��z^el�I�E��zS-��qʎdb��)$1Q�]��n [���i���K�)��3rhw�O淓C_:�i�è���	N6๟^H~'��s�hp�/���lg���h�Q<���w�v�O\T�X|���#��x <�Ѡ�#���^U�����2r�[!	�i�����o7��o{����{��7������U�u�w׫����u�u��竮���]w]ww�j�뻿�W]�]�������u�u�����뻿�W]�]��W]�]ݪ�뻾�������:�������u�w�W]�]��:�������u�w��������뻿�b��L���2R�� � ���fO� ă�Ǽ�T��!R�"�
R�$�()J�@��D�U$!!�U$)���%J)�PHUT�RE�6-��b�E��Mmb+C��сR�5�m+Lō�P�"�k[f�4!�!	���Ju��f��m�QT56͍[e�%GCUtj-aM����W���
��f٭���e�lk6�٭�j��m�4�Pf2-��*E�mT�kJ��J�����lŶ>�U:m,���lͳ#��  �����:��t��@��UA�r�ɛ��)U[�G��2�Vn�6X�M��ޢ�f��������X5���yצ�sZ���'��%4Ĉm�*��  ;�y|װ�]���6�^��=�N��(��/�•�(
(�ޮ=QG�F�w/7 �E��w�(�Ѣ�(��� ���Eh�n���EQ@QE��xz=��/Q6����-aPh��  Z�ꪊ"���SGg|��ևc�3t�l��u��QF����뭻��N:W;�\�˔:����ݷ�w�����ٶ)�$��h6���-�  w=�i�+Uد���z���s��ݴ#���n�:�Gn��]ڵ%ës�ͫt��U8��^�UN�˞{6�hۨ�]��n���z������(�E�lm�A
�  1��[�\�և� ws����m����V�wni��ݺ��h�պC����wvh��ν��wn��������zn��]���IL��*��e�_  >�{��]�wv���S�����v��F����*4{������J��=׽�۴h��^�v�˻�J����X����s\4V����wm�v�H���*B�l���Uv� ؾ��_bv㺏w��������P�O=�zSgH��j���9V�Q�hw^��^�뫱�K��`�������]5�Z��u�݃�.��H�4�a�ͪm�JUM� ;��� ��N[;��+n�n��x�X4kKy벀e^�ޭ��hh��!���j{upw��)k'^���y;��-���g��]kl�t���5T�1����0�O� ���t�v�x܄	�鮹�+T��;���m��3���4�m��������=���U��)�һS�N=��l(���s��ۣ�^
�f��R�ڶȋёv��  .��}u�n��æ�AC�����T��S��[skJ6�p��=m*Ə^�x�^f磮��:^���v����S���c���ZSd�S�	��J@  Oh�JR�  E=<LU*Q��  O��T��414ʨ�  �OI! h������?���HX3�/�}���ٵx��<�~�=���~���^���?�W}�ED�T@QO�"�
����+��TAYAQ���+�|�Q����C��'����H[b�3���	�l�B��#�4C�$�5�vl�y���5O�[�H��VH�9{8�p�����2=����������q2�썚U�����V%WP勥Nи��� �T���@��T{�.�;QUAMF᭼�*��itD f�tY�kJ�v�RԈ�j��=�&	z�"�4}*���e��+���ۏk���s6k
�1V1y>��H �-v�A��uc�,Y��;1�4��Ӕj����VM�
]�svL�`2#"ƹ�չB�]� �wp*ZՋn�W���$���]��G-��)0m,7W��į-!l`n�H#�<v��7Z�V���r:�m�L"[ˤn�Rr��n��q拥0�A[F�#P��M���m�[TnѡK)�W>X��B%�&�u{qӅ(�;ֳr��#�T�6	i`�f�̻(iL������jAmh���Q��UH���J�ۙdf��Xߖ�K[i湲Ka�oo�,프�B��#n�	&�t�(M0 9N���u�Rm`�QA���S����Z�Q$NZ�Fb�(�75�[�Ú�-y{a���5D�W��Vu�Ta$\(�WZ��7�T�±��4eÈb�����Џ�Vf�t��NZ�*2RfY�)�d����Y{aT:�b���XO(m �-�e<Q3��&Q�&f�f$�5�7��շw����93db�nQ3l�M���,�H�K2�n��Z�h�C������lŶ��N�a �ux���G�vG�@��eX���o�n ��R��UJu{A*ܷ��V�e5S
�h�^�A��u��3m�h�n32��ҕ˖��4�
ToY�R�.�Sj�z���X�ҒY���e���T�V�[�jupB햨0����n�i�y,��Cul2�X�
�ʚ*!�� #��h�I���1d���k�=���}��)b�@j�e5����t�,���ա�l�X��R��&-4�����3Z�wm�F��Y6�8�����@�&�ՍM��ܽǴ�+%nZ�6I3=�*M�
�c&f8`���� �Z�N��`�H}$���u��k��MS"��[����m�$f������*^Y_;�P�s�˫��v��\t͒�e���u�iL`=U,
ȴ+3.ºˬ���l�K���-r@��&}��uD�r	XK�eJG/hb�{�J�x.臭*+Y���NૠEJ��Sܭ�YkM�-[�
7�PE�1��t�m�u��D�w�������]*�e:�Z[��W�ܫt�oX�i�o4Fj,0�J�וVv�?V��[��m;�i�u`��E2%L���{*�l�� �8,Fb3C�S�� ӭ�N�r[дP��d�4�j�VVT�u�|�e�˶����wK���`I�/ ٘E���Wj�<�2 �P� U�$0�U.�i0c�,�6�X*��NMX�߶!i��7�:y ɴU��
�":��qS/i����{�Ѷβ]�ͺq��+(iP�2Q��n#x0e���i��Z��Ua�2�Lת��&�6��c��"����>���x`2�ٱN�	)eԼ1�)h52���VR�XR B�ˁ�5�u�iM���.��JJ׃�n%v-
�͹-Õ.�$�Ӛ�]�
��xHFS֮���n�Y�QLZ�L:�[�$&�e
u��.����1Rjx�Je�""�@v
�h؛R�f���U����rxt�Ua ƈaV�-�j_�7��Qi	�^Z�I�U���
t)у\��n���-kYW�Ԡ	,�}b�R�yL� �8�o&���n<	�x�9��*ƩF4XN��'0�iJ�%�6un��pV�P9wyc!�N��Ir��2��!u���-�M-s)hU��gU�*-�s��f���'b�S��M������t
ʴ�����ٻ�Y!Py��l���"ݱ{)]ظ����-u������3KZX���)#�7SN���i*�:�Q�5�U��KЫSn�� ��7ELQ�vb��)�mkP�3Sf�Fj�B�X�PV��4�=UG����ݴ�vNl{�K"ˡ���M�f����Ζfl����O.]f`J'F�vnDcvŴ��6���cM7p���m�n,��Bs&';�7��T��M�*m�@4�
L�JT���5�/M+4jE�]��n�-�eX�CoZ�S���@\�x@���{�4+�KS�^�RN٫v�ɫjQkP%k�u� ���J��7�j��	٫ѹH-R΁�M�'���b(��w��LXYz��"-��O[[brQ�lb$�h|����E)�����3A-eI�f0n��Z�'h1��-ݓ*�&�(b�]n��{)}lR��cȖ�r�KT�6,�+wbJ��2o>��x�`t&�Ӄ�(�P1fd9��ndP�tR��2d@Ն\`�܌D2�,�X�C�5��]WT戅m�**�c2�d�si��Z�Q�oC����h�Ӻ�ڦ����T���-U�e���bA�qP@]^7�����)�Y��b��M�0�Eb޳E ֭�m��<Z^� A��F�d�e������,ϋ.�vMk� �[qÌe(�.�c�ZY��Ħ%�1�j��qm��F���n)HR9�k�NV�;��ǖ��մL[&>����u�WÊ�����3`ٰG*�omTDj ��K����CHZ
���<�4��y ����`J慱�h7�13��z�h��!b�3Ӳ�a�L
ko�V
;y��]^�I�m�ӷ��ݓ�5�fn��f�h�.��0����3�Vk�C	�DnZ[E4��r!y� �Q`�N�;��Vŗ"�7��Tp�����M�WHā2n�;K ��#r6�xZd�ջz.�@���wÁ�B�Xw*4�n/�m�íI�jm�ǔ�&]�w�"h�j��1��ܑ�	��h���F�KYD�V��FηyO[y�+-�Y��ke˥�n�Ƒ/[n�'�ʘ2�-���ڤ�7�i������8���M���
j�6:E�Տ .[���i��e��6w���<�$e ��L+����.杖ĚX�KGԬ�ւe�쬒ջ/5]�ӖK�f��2lze��X��s^B�A�����(�z����kY"�h��:���uv���ǚ,�䣎��Vv�J��,�ב�OB��SF��ëݳ��
ks\Z):˕!n�q=���P�iVj�Q],y���.���pX�E��=�B^��kD+"mh���,���\���dVck6��>�ӳt(�M��K!�f�q%-]�㲣˸(���[���y-�u�x�7
��ٻu-,�^�yM6E�TM�Y�ӱI=
f�.�LÒ�]���.��f�PaX	�����x�]}FX�������ؙ���e����f�	��h�-�W*��f�#tL¦XM��z!srX)�^O҄�tĮ�5`���4�&ڭ�XÖ���MZ׀j���Z�]�<V�i�`
���o
Ea�!�/ �a����-M�l��a�{n-�ي�����e=f-$�b��W`CcaE�#cf�8��DV�Jͷ����Z��ӥ5&� ��R6ᤲ���V[�1i��Y5*X:ਜ਼��ڍ鵅��0�V�6*\:%=-��2��n7�v@{"�?4�t���$֭��͚�P>�JI���\Ta��k�K͠ƶ��b{(��y�Z@�li���:���:�n��Q^T�k`�E��!G�P�Y��0�zd��{�6VY�P��Au�V^���n���#e��*�wp;�(E>��-�q"6ek�0e�*Y�>��u�h*_ v��ԓ�{���Z�2㛊�Ȗ;��LmZ��b]$0�УK��Vie��.bm���պI�G1S�g0,�]�4b��\M�젋�0�)2�� �2��2�X9���(�p���MH�hMծ�#gn�V�������ҫ @L[���&7��0+v�}�M��FBܩ[��6
���Qٗ�5���WE��GEf�0[DA��i���y�c#^H�:K��֥ �Gk1z�f;W���q��ե�֕ �̔��Iݬs>��n�Py[�j��mR	'�*����DT�;�IGQ[�L�������_^R����Y�p�Q
������Q'T/(+��:9��c\�iH͹r�2���ʙ�s4�H�LS{y��
�/~����>�V(��;����AQn2��kF����Y/J�s5��N�)]۽�K��Q��$�r�/]짃��@4)15̴�*Tj���h!q��Ճ�%)��q��64&]�,��扲$).��ƙ�;���z��Cp�u慦ؘ����.[;j���F�=�z��cd�Ŕݩ�7jYV/�[��{���"����E�P
�Ȩi� �� ]!J�ܚu:���vii��w�]��Bno�0�QѨ2m����zY�2X%�:���/�^�bX�l��p㩩d���9��l����`�.��V��bP�$� �,C�%�y��sM�Q�p'�t�w�J�k�UIVVI�n(����p�p�Q��n�b쀓�)̙�
o,�f��V�8c)���u���j���^�ͱ[��,J;��w�G�
��e�i&�Lh��`�)2�C����7hmJbN#R�� �f��p��n�W��%Ne+�0�Vm���H$�,�vŇ*�qf��� �����Ƶ����]�/"�����eV����m�B�8���J��
E���+vuc�@M1vl٭-Ś�"�KB8K��B��,%	���T{z�B4�2�5z��˥HN?�Ӗk5���6H���fO�8֢��H�uEW�f��E�T�x�2X�������g���L�82;CQ�*��%HT��YY�b�7&ED4�ʴ-ۦ�!H�v�U��Y��G�Lڔ���%�,�h�*V�Q̕`�\�o]ݛYp��^'�%{����]͐��K�Xu�h����@R�h��vڳxU��<n���`ѷb��<I�^�P1Pj�jMͦ)�0�Rz+h�۔�f��qȮ�\���l�1�퇯E�ˎ4�Ww+��B���VQ"J�Cku���l�I*�BSL��SSP��m�7pV���b����s1V���ʾ�`�sFiDv�J`��H�YRT�p5u)c{o3n��sE�!�Z�/jn��U�a�XX	V)����u{���m�J��+5Q�Cƃ�K���YX�G,��@	+&�ef���&Ս��07�f�ej:�U�ôvk�Y��7kV�7�x7o�V#o&��e7Qӵ�Z�ݭ�NE����2[U��zi:�w�kMeiJ�����f�n17�I�a�v]n�	�Q�z*a�鈦�+�6�2h�Y�KҲ4�t��ĩeڠS�$�E-B���g.�
^.��u�V��ި���j]-����^���Ɗ��.��ѥ"Z��
�`wp�� ��nP�Ʈ�˳�ۦ�60�z�֓�4���,�6��6����Y����& 0�A��n������L@��z�)4��,YWF�l�j*�Or�QS�y�a�W�`Z��	.�`��\<�My�2:9W>eHp��Ĕ�[���nҟKf���2�=�X�aɈ�.m�nh6�[+Cp�K@��ݭ��-=�cS\�������hSVB��8�N�謢��#t��Ų/M�9����n�<F;�W� I���[�/g�`̰��a^9qH'�6/oFA�2Hh��`�4U��3n|$����-P���6U�5�vݦ�"�(��b��2+ &�^դ^���0[Ki��WR��N<ћP�mӵK�b���2d&��"�˧�N�ˌ�b-{��ٹ�7Y#��Mk؞P��k6j,b��pc&R��h�Z״���30e����؛�J���qj̑�[W�DƉ��*X���K��'%cj��j�� ��S��e�� U!���i
l��0���x7�Y``��f��F�]���5��[q	zZw���
�Վ=a[��o��x���Hf��JŤ�*�^�^�7�qZ%ܨt�oP��� �s�u˺�jH�uf'�Vv���Gm0��Tc�
45h��2�f� �MX ]:����[����Ƒ�2�Z���/,V���)E�u�ى��sR��:jbU�&`f�d��1��אt���t��esú�+�d���b��c!8#���ܐ�`�$7(K�% l\�zd,&�Wr�1bF�0��RҪ͚7aw�N���bUyA=:5��#�t��4��Rɴ�e��8ب��^��5/QT[Qɗm�f��o�2��P�>5�Q',�gW�^U".QJ�	�d!9+[��Sg0յ��j�jK�ʖL�(�&�r��F�47fb��\��[*+;�F�Ph�ݠ+���[jc�[na.Ԩ62�U�(A�#���Pl#!�Wtr3@24�����X�8i���#T�b���
uDD�/T����Ĭ��j UČ��^/���V���fV[�y�.�m�E��8��ՑT1a�oXj�I��Ƶ;�� Y��WunYnmע}.BEɴ+m�,�*Śωj_w:G�J�S9�-[;q݊eXMV��8��;�AR���#P;��@Jδ�Z6�ld=��H��ձL��eG��P���{rc�C1���YY�[�RɻU����ˡ�EF��N���̬4r�5�&���X���9�u�&ĺ!��
)�Ym"R��0�(��(:[ﺈ�C���nQgQ��n�vܮޟ?<�U�xN۪���4T�6\�opG�Z�0�UKi٧�j!�v�qQ�\��ޢ�cΥi�=��D��N���U�n7:�R�,�3����w:v:��{'�ųodv����f���`,�d6��g�COU����vM��l���:`i�c#;/^l\�������T�fSL��ܝ��0ل*����wY�	�~ﯨ��=z�m�[x�z��ݏs ����X�FR��ئ+�z�*��#��8z�n�3_���ۢ�1���Qń�a��=���Z��Y�x��Eն�Ck5p;��+	�=Ý�Ü�$�q�9�T�Q�[j>5 ��b���5Rn�i�fod��;�`�����ӕ���G/JQ�V�+.qWCW�][M�|�CW��/��`�@˫�u1��J����nSj!�aգvM`��;�$�hS�C��� hT�3k\��`Ӓ�ƕ�7&�/W1�ג)ǛW���1�&�׸0'��8[{�u�$���}3�pm��!�(Wn��sY�y;�F��5Q�t��c�|���q�2+`�	������j�Z�R���%f�JKص@L�fXjﰶ��
8;7�>8�)�7�eX����S�^k5|�Mfi+%\m�	�ۨEw��6�Ś�f��O��u�D��m���%�O�9����5Ϝ��X��|�N�\z�e`�oL7�����Gj���!�	=k}Vu.<�������9�ۆm�<���qQmk�v���(�j�IÛ�v���}�r.�9	ì�V���o]��UYz�A��x���`w.&�S�@�;ׇ*J5;Z{�VgNj���S�̤��ۍ6�)�u�1�@�פge@�_eҕ	w,,�]�<�R���h��RGY��*�s6; a��U�T�u3�դb܄_r6N%�\�,���¥ZVh��F�.;�Z���@6Ͷ\#Ǳ�BA,#V�n�<4�8[����r��)���o�w�YqX���X׏���* ^gv�4����cJۑk:���A��r���ʛ��U%e�����q���z�9��[�����;�#��Xe"qкآ���wn��#���]"]�6U���<U�e3���ƶ�oQ�tR�9���s;O^�C85�x4p	+wd�_NS�:uJ�����n���k��f�`��k���D0��(=���rJ%�Y��{�ܯI�j�Zge�5x�/Y]�b殢y2�2���)��쐺 �t���%�Rb5v��h���d\�{)��˝��e+���>��)�]�u�}7:͈����go-��5>���t����fF:n�fb�\�U��2���B�e�fu����F��`�I�vńŢ�c�:��A˫�xܑ�h��m5v�pFkk�AH��s|7+s^n���Ô���>][rZّ�g7F;�Q�8S���/mpĚ��]�j�o���4�v�o*\��^)*!M�f��Nx�
`����ܝ5���v����(v��xu��[��^�r4�&�p�>��B���m��=Y}Rѥ H5���pk-9��xV�5�u8�8���	Z%�:���{���#���
V��/�,�!]i⹙�P ����Ґ9P��_h[o>�-��֔5��B�����;z� w\Ue�������q��y,<��Qռ�Q��F�B'pB�]�fKq�\�����s&� �S{L�7�9��]�8�l��J�%Ѡ<�w)A�.�x�4�샪�EqOAG9�rл� �hP�w���$Ŵ���32���lV����sH�%Zten!�{+��Q�R�L�Gp���.���4��jս�X�ADLL��	xYu�X;��{�H7Z��M���͕]tC�
Z��ꬄY�[�dEm��_Ө|�K):�Fb���؝�o*ܹ[ӵ�uY:�7 �V�� [�Vݛ���	C9=�$�J��k(�OQ�WjZ۷����Y\��Q�K��m�a9���d�Gi�Dh.Te�<J��i�	�M�����ۈ;�Auo�l��䫥�����l��	��d(���Ք��戽�ilK�sRCw�y�k��O=�V)�`c��y��KVB��6�lto)�dK0���"+/�8�������u<�(&���2#��9]e<�b)�蘸�7��\��o�����*��ҧ������Lp�<I��֚}�Ж/�m��Q#OT��X��u��o��H��u�ւ2UдZ�hhvY2�����=��2�Sx�u�*��Ճn����8-Ú�@*�_hY�*�vWiֈ}�-�ShI:�Om)Iu�X�YX���"tyU�g.�)Y�J��xY;��b�J���ے��Ƿjg/��B�1�wQ�|c:pc&-��.m�2>.��܁/f3�y�W|�U��=e�40:��V<v��f�q�Cك�a�o��B�̗Jˇje�w�vx�q�w���Y�jq�xM��Z���a�)5��۔�] �V��{r�'0������󝴷ygZu�3xZL��_ql������Uj�٪oD�-����^�U��V(�oQ���.
(�ͦ��Ԧ�>[�K�su�|3�0.�1�Ϛ��*���u�.e^�.X��#z�͉W�)���V�N�`�J�b\9fֈ�hs������*_I|�-�iq�+�9wXBA��x�>��7V7��*K���-1ɰ���ƕfY�)k�CZ�k�f���6�t�򒕽�?�|H�]��Zɫ9] �QĎXu���E�;7�������ob�8��T?Z�|���#�gZ�];79-�#5���gM��#���ٮ���"�qY3�L&�D���gv�JY��h�cti�q��,`�SaY�̚�u���(��V5/��+�!����8*�e���ػk�2��z��0Phɼ+��m1Wg���������kw0ʨ��0v�A��Պ���q�(z.��̾�;g(���,&�c�5��O;fԍ�9L49*ަ���	�7)RQ��t́��l�Ž�dK}~S����p<�.�aӍ�Ң�!�Z�SWӞ/�@,���7+�9B����/T�U+��H
��f]V��u��u���]]W�p�g�­%�t��j�x�֫GS���W�cB榝�w�8��C7t�f<"Xu�#sA-)���zc�b(�W�WE��tz��[.�=�I;o�2N��5�ŋ.�fL�"��m��R1�(*V�T�W|�1�3�*�)w������Z��Ծv�啣$b�ض�a���<}�eī�7`��r=i�):}c�,$�n�z����YpHAyYe���4]S',E�j��޴[:ͺ� ��ԴqgW���ن+� �N���R���6�ʩ�^ο<��Y��9���^U�
g;��2���z�.�m����j�{kn��=����@V�h�"�AG^������v6�R*ԒM*�P4��˟���6���.��t`ũ��xh㏻X�w��&���t&U�U6薺^c�|�q��ƌ��/�s��p\�W�cb߈!�HWm�Cm&���ECʕL[/^�W�o��8,D�n��;JF:}�
�|9�/�)m$��t|�]s�c.��*�X���*n���b5`�#}����COw4zc�U�B���mV�;W��uF�4x:E_-�LTjZ1K����?�Ϙl{��rg����l���.mͽ{ƮYꢘ3����O��lk{ٲ�p�un���gf)9�58c�fT�f	}�N�7�p�KB�nJ�	�!�X�qY��{B5	��lA`�[�︵[8����L�o0[GzqN9~.�/��=�b+�Ƞ��}�v�VЫO�{�=�Wn���E]Y��G��y�3���@�Z� 5���Ccn��4��]s�G��r����Ks^��eH�E���m�[P�hx��.Ż�m>�"�l���T�>Q�L��*	��Me݋t���wuo�魵V�M\70S�m�kc��ⅎ���n�D^`���Jp$+XM��BӤ�m^���L����s/�@Q�-���KW&9�i,�w�6���r)92��ћ���j��f�D�cWcs���U���vk���vnJ��p]�����3g�\��	�&Vj�f�z�!��=�>�y�C5�GҏILsONk�8ޛ4Hx10ɻ��)� ����u�!�6b�Z�u�m�;c�:+����b*�Ҳ��\W;����\���l�/=���r��Y��\���3�t3]e.�Ѩ�8�nb�j�N���otfM��b_
K��Hi��rL���J�#x�n_m�jQ�hvx�iJWBaSW�������[\pf8�ZH�.X���Uo�A	��%���h���)�P�����=s�j���,��e��k\��^w:�r�C�94^p$�U���r���G]
��l+����{�;O���a����]cqUƶ{8����Ă���(��w*�%OnRl�:���sR�j�~��g�A����>�����!]Z���x���ɦ5<�N#����98[��X������x�s�g;v�xqr�6BX�h�7�#YQa��x�Ux{�`ޮ}��i��{������S��rp�/�,Ut�_t����o5o Q��^��f�f�XΣr���Q��`�&6��� q�����мck#9|�*�Y�N�^��ٺ�y��_���]�Z;Icu�Ҵf�Φ�Ď%�zJ %��}Pۣs�.�w7Ͳ�Y��83EgQs*�B��gu��3��"eE8����� PP[I�ta}¡��֓�6��,H������z�gc3��L����^��d���� ���o���U�(F�ݱ@؏�$p�7����W�5.�#v�YQ�t�v��*�����j�Z��ͭ�}�Q�)B.2;A���'�>�d�:��
�*��d��t=z!K�37V�q�io���1Ɉɢz��͇;�Ev�䐙�r��>-�Nպհ�}�����W�5�9�nn�te��&'�
��x;aq��&�;Y���I�� �y��+6(��LC���NZ�~>�h]r7��}��>嚳(vIr�K�z���"C v��vR�I��[CG��4ћ["�F����]��Y7��.r��z����vZ�����c]��+HaN3�[V�YYAd���αD�t����Wv3\Oz��hU��Nn�����c=ua]�+�P��\+,4����{�.[j�e��e���B��ኁ����
�{�N���U��l㽇�g�u��obk�]+qHr�V�,��L��G��j@��c"���|�a�:_v'���.��Q&�5���'jb�h��
�\����׏%��GZJ�K���٬���&]��E��
ô��+��oq��b��ސ��1�z��H.���f���Ž�^5���q�S�eYɜ`�����ɼn�NOR`X�b�6U��n[c["�N�1JZ&�=�ױ6 �CV����g��W�����r�:�t<�(�~��dk$gB�|�i���np���,��oVMOy43�g�sfw����y�R� 0$r�9|kq�]��g�uh���1�p��ur�Q�s;��lo ����.�<�N����g^��&�Q��6������1�N��9  �������Vn֬BS�J%��W�(��K��L����Fj�dҒ�9���S8������s�*Z���!T�i�7R�jm�]X_6�T�l�f�(�*u�=� 埞���#��tzN愾7���̻��*u�m�l}��ԜŚ�$ʷD���O[L=����UtG��*��ި�p��L�����u7G�F�aϭ=���ۍ�X'�qx���tb>2<��v<���Gl-�c�\�y���K�j;�#�u-wQ��:Vx������٨œ;x����5��-�SU�j���%s�|���s0�B̬GbN��*�K��e���M��vX�DU�n��a���8�v��_kaR+6�5�{S��X^�D�=<F�q_+�odÙ��S1T-5Xr�r+�2��H��-��������4��I��ʖq��7v8��E�h��O�}�2盢ھ~���^ms�ˋ"�M8��SEF6�r�˻��V&�ܒŒ�f����P�*b���rl�xٴ����ZUY\(^u8���,��V��륓�E��ö3��Ϲ%&l:��̌��W"��#����&�k����7��f,W�ͮHʂK��%°c�����i�h���`�YM>��7W�Y�[���M7�Ei'�����j�<����Ҡ���3���K���!�ݭ�k��Z&T����W5�p�> �4�**���u:g1d�7��̹/�u:�R���s�3{'\�¨C�+;�!Qg1����f�rc���<(`l\�KVk%�y�z=fjfueF�
	�޾�-�������hn��U���!��3h�����G,�s_>��w-��ޘAԤސvp.�7��|osy�ױ�$Uʾ�ts��>tq�uz }�+�)'�q��x׮<�4���E�ԯv%��C�/ ��#j��x�+�7��r��ð��&��ϔa[Gr�]+�����nCd�W �j�4��J"M������� X{�@��ꗏ�\8��k6]YA���a�W�*�r��21�q�Yb&�=�e��(���M`/C~�iQ_0XW���zz\�w���E��_��p��]Z	S)t�\��Z�D9��V��$������GM�R$�d|E�gzG�W]d��z�Z��I��3C��]\1dp��ܣFҔ�a�~1��G����>��
�aW��m�?g������S�c hnt�M�v��;�[����h�Ǐ%���iT�:�`h�����]P��Z��-�&���`맗B�Y,�8�tǩ�Q�b݆�����◩@g.�l�V�:��ܫ��X�YZ8ۦ��?%��-�o��J�d[�w)\ީ ��j��U�z_Kog]��S=�����z�����nvH*��ASXܦo�1P�6�u3����p�,	�d�  e��]w�����fե���j�o�GF�l����W�m(c��.��xV)g�O�vf��I��j�
�/0��J��nL�����*���F�%��p�^����j�鎖�4��Y����P	:��e9��B�ȁe.�t�J��x�+�sr�}w)7�U"��b��*�H~?LV:zZ�ҔM�>iî\���^n邷:)J�Xr��5U3�Q�ӭ���O_v +��f��ndz����U�U��:\���/����r��/0@�G��y��]�:�� �G����WG9���	�n��sV�5%[jf�)TIK�f�����`u9��t��Е+�����J��� �G�n��E�.��j�*,(��wi�F/Y�7��M���+����l���koxM��ع����1R-#��{�6�`o_rÔn��!χ�����˓�R�Ӭruʥp�Im ݯݞ����Ha�i>=G{���֥�fHތ�BB-�1�V���՞�4����Dm�̫�x�'[j�]��ƞ�Q�K<r�y_%���^��"���mc��3m+��N��U	!xs�!�X�#�V�N��F.�f�+�W��qHo�{E����EwvQ;� ���ek�2�a�`d��A��x1��QZ�h���}Ix�j:ɴl�ܧs*_%A�'i�u�O�3if�
,��$d��������W_eⷢ��/iT4�!t0�28�8^5Ə�8��7�'ܳ�gR4)]��qx˘�2f�S@{���5���['sά�ov�V�3/w�_$n=�����x�\����k�k����H@ә+]i��Em큃me���8��5n�|N,Nu�#+/�-�8K���M�Y6(g3I�y�L���y6\n��'2�m	ܩ�],�3} 3CD��w�������F(�	/=Ĥ����ov�fN�#:�7J��Ԗ�����xA�
Ь��,��Y3tH�u�t�'K�4�4�r D�w�՞0��,��
� �f
i-4uv2骖J��;5�6˛�ǥDnZμ�\��L<gZ����<۬K/Q\Pݘ��L4m2p2�V��ɗ+���cxK&a��}N&�̣hJ0I�wN+����3+�'cB	�͎��9�2�
��� �%�g;Ml��v�s�������pɗR��\�;�0bg(�W�w�kZA7)WVA\:39D��Hު;䚼V�wVZ�EP�6�(<�J����e�_,�4f_Z
5`��	m�Q9[ӯ�x�R�j��5�7^��7f�=&�9T 9���qj��f=/��$b�S�SqZq�XΎ\$W/YEˠ;)y�x���=+]q�{��)��U4 _.�	ن�+�r涮�&�7"�{ѧN�L]�z+��,�Å��Ȏ_1�� ��o�)[V������utќ���Vr��Ѣ�cЖ1���b�G��
la��ϵ����
��sk���2��oT>���j7_@	�ˊ�����%Y�|#���'� A1s"ۺ���;0�Ԑ'e��x�+su��(����D�Q�VEܾ��K��:7.����dJ��
����=[L��jL ��{���m�j��VZ�\b�n#�V�X�F�Ճ8�����|h���������-�&��ڌC˺��|.�="����9������*e`{)s[��ޗx�*N#ST�zj�ۭT�8]q��m��35�)���1w:��7Oڥ�|WU���wH�=Ǫm�&�lz��r�Z�v����d��Z6y���K�ەz�Ԯ����[�����H �-�� �7W�Ŭ����DV�N��ΗM�%��E�D��۰%;(g'{�p�s}�Qn[�ߣ��Pd�i�<������Q�Y�m	�W�V�������#���$���V���04��n\�"�3N�ڙE�F'Sb�lR����4�ķ�j�������.�j��0�]�wb���/`&-�!4V��80J�۷WL� C/[��`^s��з/[0]�~�����B{�J��0�X5U���o��_k:k��7���<oxYp�N*�'�`$3 ��1^uB2�^L�ēœ_�^�e+�M�0����odukW\*:�1R5٥�V�#��Cz�r<@u�n�'wlҷV�t���Ռ-:X��yR�i����|[[yJ�F9WU����Cdh�'�Bݚ��v/�]`n�+'��%�G��Q>k���Q^���ݥ2��j' �52S�lYs����xU���B�zh��~O2��t�sO��������v\}֝��M����Y�Wy��inm��>�r��R<�ZFg�r]�h}���_P��-RW·z�f����@�Z��@ݰ�W=YN��g�~;�֙����kn�a��Y�Ľ�D��-T[yv�tR�6GӮ���:a�56XX��Y�tH�r�zm�S�"�6��=���b��N�q<��Ț4���L�b��d��6��:L�Z�s�1���F��)BŨ2����c�"+�:Ai٣[n���u���]<\h����T�L�	�f�;x\�s�cbK���rI�ӑb���:p4S4j�1O��a�sińv�S{�:���Z��1݅�v��j�z^.!"��S7&��+�m�m1%V�x�.�!u�\z�t���7��x����IS�N��8�K����	fb��,N��Q��M��X��4�	����z9���Ӥ� �*d�6^)�4	Z�i�.d-�ՙ��`5��FԻ��<:/��&8Ru��wer����p���{)PaL�YkL�g5Rt����ß P��X��NJ���SXw}�b,�R�:�Z�%���9����[�!�uyl���2� ��:��@�������3k׾+U�(���	�6ppU�Dm5�T��Y<��=M��������:�I�S@�7  ̭�VJstCJ�U��]��dx]�"�t/GP�m�A��9�vL{]E\�8Խw�\�Wr�L_xfY��2eĪ�xr���>`�C�6���em�+;��=]�/�T��j�TUx�G��I>9�.��f:,1���.
�3�N�0�(�����N�p���lg$Vm�⸷36IoU`�~g�YuvȁM@�F��IY�3:��ܻ�i�ũY�W@�����ܑUК ��r������d��w��\;+/�����`[F�DjF��]Cf�i�yX��܇���z�����X�ҝ�ݶ�Mu�z�X�m(�р�S:]�s�>���Hw�ľ��ˢ7�p�T�N��i�~�[d�7YK@{����y�z�T����1+O5*�Z��,��V�'[z/�'�V�:Sk&��q�=褂�<4�ĉk�8(#���E5�<���-���ɑVuc��tl�K�E��x�Vٹ�W�] ���6��OΈ�����f�	r�h*�26��;&�LXLmb�\�[����f���aiy����Uh��C[�dM.��@���F�	�p��D([r�`���PU��9W3�b�D�r���k�����c�5�f�ˮ���[4��%)ÝPᦄ��t�}@S;-�J�2/2���P������՗��Kh��1����� �� �%c0,U����+h��]�.*�r��D<'���"d�D^S��R(v�#�����W�8�+�w-,�wi�ܢ�J9C�b�N\�{���nooh"�� ���nTЧp�	L���	ǞI�K�sZ�xN����x	�+d���>�x���@P�fo7�.�@ p�[P�bK�$N���˖������㼋�ېVe��y�d��;eVj��Ar'��ɶ���2'[�XO�g��m6%wD>�znHn��u�V�c��|��vu��Ўk,��}�	ȸ� ���3/�����a��[�F��X��$�����
 >��`�\G*�Y��r}�{���v,&r�+/�7f��@�J�����ڼ��@+~��
��sc����M�j�%�סc�V���m��Y���F,L���.�Mx޷;�΍�8�E+�=l��f�ĎH�b�I	l���s�c���8��{�S6ۑ���K5h�=ҹ�en䧅T���	>��x�m�6�tpl�b�&��høAN�Q�J�68l���ŗ�u���u�Ȯ��V@��Μ>�n��҈�gL�	��nx���..N
��{�	��c#��c��+Gu�/4'-�Ӻf:��Ŷv�uLVwr��X���x�7��YC6cF�Y�oHĩ��G�%齩[�b%I�:��n��Y���Ȏ�W�m��4���v���WH9p%J!hugl�=*t���j�>}o�;k���77�_m+���幊���S�)1��7��Ѧ#3�QM�&:���u6������UCk�G���|����.�p&��:���Y N%�0x��Yl�4,;/���{W9n���(�iV�,�)��`T\���+-Lú�f���ۖ�.�M�4�+o*� 'E
]��8%e&����m0�]�����%�s�} -��Qbj�v �B��3l+v���.���[{�kwx��̾��f�5t�&:4�A�*��݌�8s%mK�����_}��<��7���tR�R'�������s�u�T�Znm�B�V������쳴��tY�{�eZ�5�\��vq9�;�[��D\9%"�os˽��:�dOi�R�f����Aз6>��v���������2�]�]K����d@�յe���T����d���6�5��p�vI�����;'t�un�>���.�&�r���v�[�s�������Nv��ywN��
��3n��5�>sxz���,(���D�d[���a;�2Ja�O�j�ꃷyS�p�j�2n�nj|�c�����JI䩁�h��8�t�ZŲev�n�`]�TKqZÔ�}�\��׊����h�<�Ff��<�cǚr��')�J3��Y*,X��V@��˷CA�K>�W$b�5��X"�aZ�����ո�]-�r�C�le�R�4��U)�h ;����7��p�j�`��4�R���ϻn�E�Vgy=J�eo5��^E�������,��%]�]��r�v�%��C'�+Eb���7V�H��U�v�8�FDx�b���Q;GL=P�
=�T$>"�P���]p�|^�k�o��c8�d�2gs��QT�r�8�b����ő�ذK_jn��xxf+�X7
ؕ�;[�����[��9{��݃�=@9�������{�l����"޼O.��Գ��H�;�.U��1<;�!�eRj���)̒"������i���u�Vλ5�n2�#�%�$�DW^��;uY\�n�8)��|��g�2��:J�;v��C�/���:���P-���җ�.Zy�W\Mjۗ.���	�LFM1ѽ�Ѧ�ȓb��.����$�F��,-ǹ:J��Z֨b�g�վB���Z��G��9��i#U��F�c�\�%WQ�6���t6D3�֛����@�j]��*P$;;��cv�؃7L0�3�L�;q�
)���n�Нl�΋3;�q����܋����N�[B�����S��-���z���Lm�����N�Ng������]͕�<�Ԁ�"5'|5��P̲lP��Vw3�h cɹ���ۗ5V�#~��	��ݺ���7`�)Z;�3��f\��fyA'�k�ε]���V���1N�����I,�h�����s�0�:xwe�d0����*w7u�E�LJ�s��j�H
������{ob�-�Z�g}�&%d��|5��V�=;6QE�.S-S�L��2��.S��%�A����,AGz�F�QWW;f1�aT�`⊼���`�cYu�Mi�c���*j��Ts����Do2[îs�"3�v%
g7(��on�+የc �ө�����nnuv�#�������[��5�uLR��`�f����U�����N�d[��=ms�uv���W�Y��$]r�Z�jQ��E#]W�3�op�p�9�qSV�bj�)WG�7;ua]E]��>k��'����p�Ћ7���9�aCJ����x��z�n;�	�&���1��wF��X��rʢ�ҳ^^�5H85Y��C-�̤6Y*E�����&�_A�Ɔ@#��r�K}w��`�E��S�sPP0��K��ۛ��O��a�LNN-ɪ�(��{*^��Ҙ�Z���F8m��9�q�2��T�I��y�����[ML}Km����uYg�,[��u�
͋�'U�7rV��p����J���Ww2�|F`W[�0� 4[��0Lx�&"�(����zM�~n�ΏB�ʄ�P���D��
�}j���l֪A:σl�$
���W�h>��,+��bF)��(����Vӏ
�/�ͧBva�lq��.]�}o�|�l74���lG%��_>�7�ѝ�Co�o]����F�
���2V�4�}�#��^M/^OUۓS�A=�������\��PrvNYv�/��X���M�j.�gV�yf�wC1�H,XG����Ⱥ���JP'��gd���Sn��)�(Ҿ��0Tƃ��=�����<c��f]���n��J�keG�ZvR�6���wz=Khd�j`�lCUlJ����K��s�胪[�����"Ψ���*�#)��z,t��j��uxK���W �q�	�K�&A�'[���*�[����K��D����!�� ����9���⋒%e����k6\b6����~wn����w7�J�sh�``6��M�=�V��҆�w�z᤺跮�΂��Qr\Y�0pҸe�!G�b��lI
�wN�^�oy��'!fA�bi�z�s�b0�;��(��C*���nYEV��������2mq˓����k��qn ���`��mo h[t��"��rJn�^`T ���+U�[w-J=M�N�΂w���ݼ��Bȳ[J^>iC�eޭ�n��K��}[�n+H����DM��u�%��¹O����%��숕y]Xkw����}B�O������avv�fP���,1Nw��Q��X�w1�6�!�dU�!!�r�1�Z�a��N]�.Fޭ�[\/r��%i�M�U<�R��d��Z��yXw�_h��S�1bT\sX��]m�q�X>�Ł��_>�3�b{tq�Sh���:���Z<k&A����4��(ڽ�k)V{����ݻ��[<��@*P������q�{c�Y.ZUw(���
��6�C���'{�1��<���I��II�H/�0����3�K0�"�����"�����bJ�1�"��((23���rbJ�)����
Z�2�2�r��Ģ�**�
S �,�ʫ'j��� �"���2��*(��������
�,�����b��""�0�3�2��*+'*�&c#*��+ �"���	ʊ(ȳ�r*�j���
���2���b�* ���"�1����02\2����J2h2i'3	�#��*�bJR#0�&�
���(� �r�s1b20��+0���2�32*��'$���K33"��	�,����,���r�������0��L��r�+��2�l����������¢���¨"&�$�"��c3(�"��3)����2Ġ��2Ȧ
�"���)���*,*ȃ$?V�n5��A��c��*�ϦwӉ�ʴ�M���Y7Z�+�H��x���Cn���k�����_w �ާɽ�!\�vW1p�E�Σ��r�n�G�־��]
�^
\�p{_s�ֺ����=��z���Lu�ੂ!����V��+���5��}\[�ic�(n�JΡ�z����=�:�U7�Z<s����H����kN��B�`�_Gډ���'ޥ;~��c4��_oIV�[ޮt;���2���Xt,��8М|�y(de���e��T��ng�	[�'������a�W)�NNĝ����О˫�=;��}��S��o10�;�6wT�X��ė��s
�sf�a̜}�y���P	��iY7%^�:%��9M[�m�*rP��zz��sj'��џEo*]y�+iy]E�O��#�Ι�l�[�^�m)�'i4���3�#�#�4pV����;41��`��=^�pճচz1|�{җ,@�z!��a�v7m��j;��NT�g+4-Bt)��[n��W�U]1�+)us=�QC�?}�46�ɷ�d �s�*�(�1]�v�Y�խy�I�>�3�}rM��{&p]yV$�}1ɺۥت>�¢�Q]�{x��ԩ:L��!�P�4���se>�]����zvÝ�Ժo��A�'�1��9�c��c*n���N�¹�$�Q�Cl��<T�J�*��J�����7�]�+&_*[�-_2�<�s�ߠ��	�z��,���_m��뫮��Kg&.�xI�g��y������9�9���c� �/�;m8yߪ���ub�}w#l�ʖ���{�,9�J�y�3���4��H�ϡw����w���˷���r�;�)�#�oL�xpy�����X���'��u���t�!�s�k�m�6�m_��_el��.KƄ�o��T��k]p�&�z2�#Xn��w���ð^_N�"=nt�:�������l�Ep��E{r嗍����W���$�d���~�SP�P�u����oW�<�_H&�>>{�wX^�����	2�<9�)��Ц;�_1L
��F�y�x�J�b�I@e)�YI�;2�bi��U�U1_Q�7n�5���<�v���>�������C�% ��)�=�xa|���ϗK��Y��W9Q�P3��VmV�*p������5 �=��S����*��9v|��~��Ca�6���U��j�u�9#=�A�X�'�������~��3}LX������'a3�O��M�Y]T%�em���Ҩ:kU �x�j��:��,f�,o:R����#�o;w�ԯ.r]������s���:�����f�����o������U�D���(����C���m��{�&E���t[
�ۗ����x�/"�=���r�r_�yBy�;ȯW&j��l�j��9�����K`�:�v��W.�`�����kunz`js��=�N;�$�,�co�;��m	zw�Ƅ���]Ob�M��DjW��Rg������J��uS��H��.'N�{ �^�Щٳ;hz������/ ��[O�"3�D�ݼ���i������5��q�O��C�_B�6�����+�*�;	�!��&ㅋ�ψ���j��Zb��⽊��ۦ���]�].�::#6�i���Lrjo\#)ʹ�5�`[h_Y�^v��+�`u{S~=�נp�O%j� ��'�%�J��6���U�Z1-h9%��{�*�k�&u�LL��㫰\㉇㋇A�;���b���R���p=}�-6.7X�Rto��v=���R����5s���T�J��gC��Nں~�0B��c�w�L��6�C��~{;>j��xI7�]��0p�5;�,[�q-e��%l��R�>��c����Y�W���p=6:�2��x:����I�vf�di<ɩ�r���.-��Ƴ�7q��$�����a��G���9�v���W��ٙ�;6M�;7)��4(�hw�הN��	9ףjF��8�Y/P&G=/�Y�t�皍9/I���1f�.��K�~\=��~�C|�y��	Jrl�CK{�C�굱˦���7����RnM�8}�hM�v3�*_���W,SdkO��w�f�yզ4z���j�5`[ѷ��88��6s���\�I�|�lF6H��B2��1uy*�&<�W���F���"'���p^9oJ�Nk�E���iI1�*Z���g@1)b�=u���=+*��g!�g�x��s^�s)�~��gwR+}�>��l^��-��5k�h�9��u�;���<s�nU� �\��f�͆��ێL��}C��K�A���ټn�s��<�3}�:�P�����-_`�d�J2%v;Y�:^�#������^@�jgHHX1ś���y���Ϥ��(����v!S��d߇�ھ�;�&��Sp�M�1r��{������v��e�@<k���l!���i>ڞ&�{�3����P!;o!>\sk����{1y�zsԻs���=a��wKq�9x�BC{��cS=�I|0K��X�4�������'+r���f��#[9/�N�#�6^)��N�5Sps������"f٧=�]hj�ڑb�����E;�b�W�z��~j�����ij����B��$6�]�{��vnx���r�޻��cѮe�v�F�0��.�]q4����s��ѝ�����zv`<3�_f�kW�n���w9y�[����7М���Cc����m_a�R��)ó���a��|�z���.��,�t[�.���Ll ���uN�;.�<ԯE�����W�e�r�'��c�+�r�� ku5�GJ�yد�P�ND�Ur��߷�+<��xy�oܔ=�
�t���#"9���z����Q�"^񽛍���M�D�5����p�?Ty���T����~s��w�hv����{�9Z��gD.�ukh]��PSwɋ��y��ɬ�w�f�^#�t�{�"�ӣk���,��1��<{C��V�~�ߌ�^��;x�Oj�X%j��ꒅ�x̃ΰ��ȕ`o�@�Q��T^z�YNtrR�Jp�gZ�6Ɏ���jx��D���I=2^K��_�:�y���|l��=�t%���uf��|����cy=^�9���N;�Y�Bŗ�a.y�{o�=����E��:�k���/��i��ͬs�����"���Gj�4���}�f�9�Yt{ս��mt�o�9�غ�g]��⼿𻫣-�"#zxڝ�9�����.g�u=�OI+l��OOM+E{N��C�Ն���b�Jm��Vsz(�7��S唬�:@��<�:r����-���;㭁iT�K�Z����;�e��T�t�گ���vCYs�fNۢ�f;Y #�:�5�2d�������Y�i�rֻR�TV��פ���j��Q�����#�b)�6�UOxh�Mv)�����K&��B�fh��6�8p|����ٌ�s�X��jt=���O�/]�>��$پ�rj��i�pJ}U8E�����~ߤ˘�e�ð�^mt�<�V�xzi�s��ntٯ3Y+u�C� ��>��}&]X�N�<=��u�G�9�"�,�ژ\E~�K �����6$�ム��{=Dko�.�3h����5PF5�����^�~�S�(y���|cnx����9ʼ��X�Nd�s�F�o4�mwRu���YմW��N�o�':5�'d69���w��I�%�]��x
7�*,�S��`�>���k��ɽq�k��`w���tt֚}7�2{n$���R�
Տ3��zHޗ��(�'�5��<�%XH.;}G�ut�dh|�ݛ{+,0V*�^:W�ʴ���c������_��U�y��]P�,зg�^n�ckv��Nya����4B5f�0v0���NrK١�`�y�:4����R���`��V\X��@�D��bG�Ф�6̻hYW7Q������fX];�u�=.CY��Nk�59��� };�ؗ�����qgR';<(�g�{IsjWXO�}7�oܓ����!��ѡ:KsJ�m�j���n<�9о�aN����r����<�}�nM�m��q��<��j���pu��}�t���_��3��W�/���=�e�F]Y#u����۱���s�>O�����$�ٞ"7����;#K��pJ{��W=�K�*g����k���3���r9���k���oo���ڝ�9�]Ac�������K���3w*�T�O:�ɔ&�&�]1��;yeX�W����J�U��-���A�ڪs9�=ٚr�\q�³`/<<;�ͧ�Q���5��%EX���*�V4�I$��j�K �C[:ǕH9�|4Z���K���{�1J,��� ��Y��ŧ�T�y��ġ��!��K� �g�ƚ�~��el���p����K�G�{6�8��C�yHf6����	��/��+�uЙ�;oH�PW9�G(�c�-�B��\{��N�;-ۖ��Vվ)���"){�3��J쿱�t���#О��}�y�Ȇ�ND�$Z�^ڋ�pg��ݜ]�M�ּ{a�� ���ܨ�m0���z��,��Y�&]����lW}t��;����Ǿ�t�`��5��c�!f�yղ�ʹ-Seǵ
3�=>��W�l�~�TguꞺ�P�Rz5�=��(7�e�9AF��o!v���䞏�w�5�ul	z]1�n�9�c��L���i�k�ϼ���z��A��;���K�e��}��;�u���<������Z8g��8x^o7[�S��y��=Y,��&xY���:�4z�1���mr�?����ջ�ɑy@�ޗ�s̝��Q����H醲�oA�5U	��e-�LӀ�rW:ۿ���/�{%�9���"����WgV`�5C���6�
��d�{E��ɞ��[�ʙ�m��Y���j+#L��)���ݹ�X��/�+���+ 5�g &��Y��ց��w�@�{�)��J��ud�SK{Y����^��{[Η�s���(�v3���U�n��̾^���8Ro2vz��-������Wnd|%���\4Y����x
8{���g���m]?P�=B��z��t�T��+�\8/̗K2�o�g2�����2�����]�_]K��hޒ�`��Am\��fR�N�2���pLr���b%	OG��G�;�Ճw'K}Yȵk;����ot�É��o��1������dzvaឰ_f�m��%v�j�Wf�ޝ�6�5�]N����799��3�t�޼�;;x�i�w���:=`bv�s�+�^���X�=[H�QO7�r�=D�4{<��Rq��6� ���sm��|�o5X�*�����:�s��^�;�dʃ����Z���L�C��7���f�<{T9^V�c�R�7�)s���yt�*�+��>t��|�G�%X��4ٙ/}��e9��ɛ��ط^�Lxl�0�:�g���Z5��!�XxB�(�R�Ȫ垷|��l�z�q���Yġ��.�`sm���35Q)޹vܒ�������xN��%@Ɗ�18�	�,�۾�&b'�} �t˺&�.�T˽@r�Άn4J��T���5ydT��	��@t82_	��:�-����Rz�+��.���:
Ҍ�e�A�u�/\��4��/�D*�m�<Fl{�s�Hł��l��;Y����n��`���'�;�������U��Fj48Hge��ȩUˆB��,�|1 �o�B��L�Xͦt��ou�+k�̰5�I�l:Ö���R_a�k4�W����O('%:�vs<��ۙ��LV>yǒ%m�@�트�ػ/f��jt�8�h~��¥������\^�����3����I��7��R��'lT�M�ھ�úֽ���{�c�5�MΧP�����&�F�B�O__�ik7S.��#��Z���Ȫe��c�sFHo�[��0g77�L�AV�ռ4w[��vgN2�*Vf«��L���$�	��u;��]�PH����7��A���6����?mE(T���*���4�9�7p�"$ofqޖ�5XU-C�gsujA�7��j ����/]���x嘀�)�YL�p�D0g^�9�nE����Ǯ���q�K�������b3�՚�:�+];l�ֶxL=�jJ�Bl/{�=6�.r�xl��і3�]�3���%��-��nyX���%���f�f�����i��ep�ۼ��Q�jV�B��}��e�ۅ8��ݱYٯV��.���e�RE�,�kX�0,a$��өYʗh��8H���(�eV^3wAF;�W�g�+�3�Q��}�"�o[�{tR�/�x.�L{�%��˯+��LզD��m�$e���!up]k������Zb+�	�.�5��U��"�3��3xuÁ�"�U�tZI�4��v��07�ݳ����y\�ƀv�wG�r��*H��pa���J�����Ky 6�T�G(tg�*��.���Mk(�rbŧS��7Z�T��v���X�h.�t��XJ�Q�i��/���oz}�'u���#���Q.�	#�<��6��N��h��A�U�M��7hX�r�\�P��|��n�Ǚ�t�ٔ3��wK6����x�uA gӀ�π�k����Z<�l��,� ��e^[��9�v=��ܩ�}�]<y�1=1�/��J}g�f�C�NYL<t�sM��#�r�M��w�-/�,+�+�j6�_Jۗ-_[j���)�ﳝvQ ^����;��+����)��/Xxn��$eHz;�3�nS����̊]��kRj!ݺqh�(a�ԯ4���\��)62��Y��m�4��c�Cw ��=ž��-����aQ
��=�/��p�\E.��[����jj�7���W���xe>�פk~��H��Ă��MQ0DSUEP�3�QUQHP՘��MTDFYUSEEAFFAT3�%SY�d�C%VNCDT�4�fe4DPUAX�D4PAUT�ERPY�AfeMSLAU13D�E1QD�5��M��MQ!1E4�0T�IEMP�DET�MDMEUTRP�K3�UD��T�!ESIMU4QE-EEDP�4VI�L@P�$�@�U4UIM���5E�EQUUD�U#UTSUTEEDd�TTMNc�UEDADMQ2SE%DUPEQ-RSQD�)��U4�E%%4fU%DdaP45D�eA@�fE��|� �>��R�P�m���K;���wa�Ϭ����N�餮t�ܘu����lYL�{�6����мX��F�~P�O��܎����!�.�j^ݓ��꿇I����8�Ify�_ϲ���w\+�Y��J�y�2�5�7�zx��[��s'zq�BE��L�5z��c����9�܊��:ԗ��7�\�'ʳ�X<�ݘ�MP��Y�M�>oH�p��Hso�����#�kxB�t蕹701������߲c����X	T{m˞����v1��k5v[���/�+��f�-��M�5:�;k��+[�y*�?ز������.��	������Hsd˘^/�ò��jp��=m��`ifh�{<���{�t湚E^�����N��b�םC$��\�9����Σ|E���.��pfT��M}��\Nq���s����ۿvT��L��J�����0tZ���j242��ސ��ó��;��b^!k0�;��'���=�l���bV��K�ZH�����+��dW��/u�mo�K����u�^��M2���]lPЄ��`��%���!Fi�1��0m��*�;<��p
���YF�R�"�{Ù6�y-�t�?[�x����s-���|� �j�������,o<X�~�S ꑍ:��I��ꏫ7��U[f�,�����ViJ��S�{��N\1G�titƝ�;'����Bi�����B��l:#M��S�¦Z�E�Tڵˆ�]J�N;L�f�F��J���y/W;�o��Ûb��Ԑ�j���鞾��S�_��U�5����[e�O��H.7���bpBPh�}9C��=6��T����n��߹e�z�"^UȢ��ݘj����g��D��p3���������q�~ca;m9Z�����x}Z�5Ϲ�}�=z��q��l!҅�u��oL�B�YD���_�s�ƺ�%M�ϧJ�{��IX:��(�x�O��S��y�TZ�A�o0�������>�8����^y:�/�	so�X%����x���U�O���x��uF�=r.%�7�z&��o�tV#��9�]3� #]j��=��`��X&��lM��mK�cw�aٵ�t�S
�p˝�[�)~{��_+���$8s��Oo;u,h<��]�,�J��+O �v_nT:�s��Z%��t]�9N��Q�6����T���ǰ76 ���h$�	$�v�zǲ�]�%e�ݗ��T ���q�N�o��e�u�[z�39�:>�=�2	�ᵰv�.���:�o�ٛ%E\���#'T��>�4�>ȎQ��A�kgZ����B�q��r�`���h8|��T1O_�R�������w���������{����]B�s}��19!���zw�nG�}���h���ߗ���n���]�2;�pR�� ����������w+���y'%<��r�}7�@~��s��#�Cך����/q��h5��|׺��x��7���Mm�����~D~����M���������n^FG��#�7'}k�q䯳�������}΍��u~��9��CP��ߟv����yh�ҙ�I��/wb���t��� }���j;����<�����(^���r^A@y�&�ܻ���I�;�]�J�O]uѹy�#��:5.��Y������������⾨&��~���~ws~}�?�<�^v���ܟ����=��|:ΥA��M�H��<��<����MC�w{�n]�����R��������'�������ؽ=��z�����d�}����t������<��f�M�R�
O�7��r�]A���NGr���p�rC�����>���~�	P�)��Ȣ����_��1ԫ�̓N�7���9ܩ���a(�w�[�����(t6i3X�gUX����O҅f4���ǩ�\�d�G]�s:�і�(�.�V@�V*Fs�k{��@C㭱�i�UgHN�ֹ��&+�;vR2��÷�8ߖ�o�Z����c�<����3>�Q B{[��^o}�V�}��A�ܾ��C����y�k�nS�uѸ2]AI�' ԿG�����y���WW��{�(����M_~/��?|�}�����w�{�!�����?Z��]���\��4o�!�7��5���Gpx}�;\��߸n���� �:����Y���U��翹�Y�}󟵠�'S��Wq��M�ϱJ˨|�I��}!�A�tj��=9�F��{/�=��{�:�!��>�)]���>�r���O�~y�'��lJ�goλ�/̏�{9@y����w/���Y+���O����ӸC��Oƻ��}�7�<���b�;��)�s΁�#��s��~�+�N~������~��5��\����}n�S��<�R�w|�;�����:��9^�~��}Q�<ֺ����]��>�=�gM����>���<�2�|	�Y ����}/w�g�����ݮFB��u�r]��{�%Կ���r��p<��ܞ�}\��ܧ�uIԶs��W����o'y����F�~��)��R�<5΄��^�s��%y'��{\���Z]y�~z�ܺ�����܇#��/�w���}���3�N}��9��\x'�ܾ�ϳ��9G�tj
W��ֺ7/ �<�:a�?� ���!�^~��������^zZ�h}�Hy����>�Oy�hS��V����Wg~��~����G�A���>{�{˨+�p_`���tr
W��=�F��d�9��;����!��K���P��y��v9}#�k��?6�<�{���s�q�|H�M����B��~����	����{�rru�����/�n�o���������>��w/��?'7��Ի�]�om���Ib�5��N�C
�:��I�D�V���	�ni?��K��K���B֌ӎiZ��=Y�v�Q�PoXgˈ;B²p�'5_X
px-�E��h�[��,s�3�1{���BQޫ�h�2��Dh�n{J��{���(H�t���Z{��M����x}_\�5ϻ�H�s�r�����u>=�r��y���w/���A�yy��wk�r�O���r��Ǐ�ꛏ�7�J�"�?w�7��w����k�o�>��?�o��C����:���>�b�~���;��r>�pR�w��仂��pu���x}��#����D��N�!cƝ�^�ן��܏�8뮎K��M�r�֥�������C�o��s��>��K�~��A���pR�������
����?���~�� �H���%5/�9��r�/$��]<�w�>�p����_Ns���9�����'���79.���X���_�ΰ�~��!����=�c�J��������2W� ܺ���<�r��_�M˹7��H���!�jG��t����/�5�d��j<�=�rBo1�/����t����Vo��?��T��}�ΰ�G�y=�j;���X�W����u/=���ܻ����P�K��}����wΐԛ�e��v�J���a���B�?,���n��� ߞ�~�%��!�>��.��v����Gs�~����f��>ߠ��t&�9'��֭��/�<��'p&�OIV#��<�ggM�'�z����u����
Wpy���r
�5��2]FK�X��?N;��ܚ�sܟC����>_A�wЛ��n�/ޙ�>�Oz�����e~~a ~���O�����^� �_��aJ�s��#${�]�%�d�`�R���;��v�r��ߘ��/��_����-�hz�t��r�������$>Z��\�J}��ty/!�|��:��)�o�)�?K�;���y�:\�����.��=z�亗�xu}_x}���?]��₥����FZc/<�۬2���)�/�&�TܥV�75?�;"D�GHZ�
Q9���}�k{erAbX��}	�P.Az�e��]�s}Ga�d�uǚ�LF���_�:���t��#y�$�Ka-��#U��8���������ꇽ��?^�����NC��;�5	��GRw�������t� �<�:J��
y�!���{|��>��{\����yW�}�U�3�r�^��T���[�G�~�W�Ǽ�'��|���{��N�<�9+��{�������<��P�s�&A�~��Û�L��{9�{|��_��~���ν�g;�;?�sz�����.�f�Zװ=bnCP�}���C�����;��qg�y��$~�$��9+�}�7/#%<�:dܿ�$�wz����g=��}�����[�����P�/�y��{���ݮ_H�o}-��3�C��{�	�Oc�0�<���O�Aܻ����I��}������s��k�}�s����5�Ͽk3f��2S�o��O���C����Լߺ�^����v?��{�率��!Op���uI�7#��>��� ��� ~?}�ʫ9���?P⇳�����j�=è8~�s�/�{��7.�%<=�G%俯��o�>��?�y�݋���=�uw�y��Zө
{����_@$}�C���e��~n��׭���y��
�������������ϒ;��a�y{#�|�p�W�~�/$5�}�о�|s���������V���������4�\�XD�)ϵ�xm����x���;��r]�Hx���7.�'��P�εӿخ��a�y{#���Hn����/��V��Eצ:��>������ErO�A2g����fl;���g�`���_��Xu�O�x���ߘ��Q����NK��=>�7.�߸��+�4ﮎC�a}�߅|�>��>����=.�����9�Z������phO��8k^��&�<7�A��w'�`��R�u�R:�q��'�]^bn]FHv���u//���Sr�O7��B���/5�����	"xYB�F�Z����HEBnw��z:Z�{m�E�v����Ocy�J��ݕ��@�� i���.��mv�b(�L��趟c�/r]��g����$�w�_�]�䦞�f0zN�9%�1�����h�:�%��=�������Fz�~_���_�B>��|�F�t����_y��%u��;^��y�wC�(�rK�a+�w`j{������u{	�`nP��]��1]
Mh�����������(~����^��x��r>[��=��|���GPx}�;\���׽<��u/�X�ԿG�F+�y�������~Jr����C�y־����z]]�p�}��m����C�I�֮@��yӨ9��o��@�%��~�.���>�r
�g!�u}�R C�g�l�����)�ԍT�vs��|���b����9{)ϱ܆�����9	��݇r�O�?o�'�u<�����~��!�7�c��}_ZU�k�a�}���Y��/j���|B�.C��K��u#�~�>�y}�<=��9~����}S�<���䮼��ܼ�����J��;�����Xӻs�F�w�ϩ�_��u߽�NH���KK���y�����ԇ#�p<���>�}������>���9#�~����H�M/+�Ǆ�֎A����~�<���9���'���׽�J�\߽�{���-.� 2M�~����SrF�0<��|}����y'����}�����T��3�~e�ǫ1o9��s���PP�:�O��_ђk�%'��9���J�/��ݮ}���7���~���NHjo�Ӽp��g�x�?}��!~�+����?C|1ރ�x��C��>�\~�}��v~�Ѩ)��c�y9)��t���&��{/����~��]o�ݏ�^�Û�h~�H`K����~�()�^�SB�sg�c�������~�>�P�
���I�xr;��~��C��Oy��y/��?o�>���9�z��!��|���G=�<�mg�,?-6*���u��Ux�q���*�fǴ?jAL�Q���1��-��t_������j��c�Oq\����
m+�U�n�{n�n�S�d>����m{�Z��c���=b��}&��@���\�(\�Pb�ޮ�쮜]G���������ǿ�o<������d?�0<��9�brNH�����y/���n^FG�:�r~:�F��_g߷��y���n^K���s�䆡�{�<��y�_za���οk_��3��!���]@��h?Gr���܎���M�B�w��伂���P�]�G�؎�䝝k�w�]ɬ�r��G�u＼ן���q��o�L�<_����+�}�ӗ�~Ul?��~��?���qԻ��=b���O�Yԯ�?��x����ߘ������j˸���ܻ����5��X�lP�r�/�#���������2�u�-����d!��/��K��ny߽�O�o��u.ड7��r�]A���'#�]^bnNH~���}��E�=�H�̜D�:���ϫ�S��6��<>�9�;7�F��=˽��unGg5�Hj���������\�r�s�����
O�9��<:3�g���=������՝USǛ� Dd���9.��<3r�]����!�����jG���?�@���Hjǲ�s_��w���(��F�~��	�9�������؟��������~���F+�NO~`r�]G�~�~�f��>ߤ��}!�A��ѫp:���tjNG������#���h~��@��4{��Z��y��mr
�����u9@rK�|tb<������%wI�����w�~�I���}��t���9��~�7����D�z��2��O.���_������R������r2�f��u9/�K�~��{�w�;��$u'a�!��Nϱ܇�u����>����d��4z���~�{Z������k3���O 8�%r���o�K�����$�7�k����]r�b�`�]K���r�����G��3P#�����4���XX�F�9n8+���7���L�q�g�]Q���@�)e�*=�Y��"�@���6�Ǖ1�?CZ���ǜ/
g��o��y��E(�=��l*��V����*乜���t9M���B��OT`���	��3x ��+-ܬ���3B�)�)~���#�g{���)�}:}�ssI�;���H�k�K�)�ܿAN��P�/�罞J�Os~��{+�mt����w.���>;�w �G<>2�>�(*�~��n�������~���$�<��z}����:���J��]��R9�{��9��Bd?K��tw#ܾ�7�k�Ҽ}�#�<~f�uv�V����,�}������O�O�=��0�w�|=�=��������~���Q��7/# |9Οa�?� ��:C��~� ��l��� �<��Ա��?v��~��k89w#�k�-��9����G��;�7��Or�NC�AԻ���������y+��}��K���o��H���C��{�jIj�vL��gq�}kZ?qe�^��z��!���c���b��nB��<���z���~f��]�K縿A�yx���@�u�#�}��wߡq��Ɵ����5���y��fpܿ_�y�}�r��Ϝ�����\�ؿ�<s��Wp?���Q二�%~������]��9.��=��;�������~߿k���;�����ϰ�w#�>�5.�dy�tn^C�Կs���^�ϻ�o΃s��~����<��A�Q	��~()0��U���K�曁�����~��;��=�9/$���^I�ǐ��G�����]��K��r=���!<�]�%ܜ@G�!��i~���f�a�&���Eo���tp�+�<�w���WW�X������y.����ܻ������p��[����Hj����t�)�����D}���������=�s3\�~��K���5�~����<���5���9.�%>3r�^{���)�w'a���j�|�}���>��O���!~�?9��^�=U���I����,���P�-`�r���)��ϲL��OA�����W��BuhG����_���Y�7��`�iړȮa�xvS.���u�nq�;�_?M�lܦL<�Q"��v_���ᙈ�	�%s���v��+ ٙ"9�ϫ�5��;��׿��{�N�|��~ם�PP=�}<�%��`�P�>t`��q�y���Gs�~�����P�}��Л���Z�Թ��\�u��R~��+�v:�x�W�����yC���+�?����(�5��2]FK���u��ш�^G�j�]��b~���O�r���ν��(�)���=_��W���}U��0�G��C��_�y{�zpy/�����ݮFH��9&K��rp������#�G~�r���~9�����{u��DO���~�����5��_�p�����V��N���U�:6�ʡ �r4�z��t��qO�U��L?�2��4�e�g�>(r���"���F�Waw����3P����7(I�S�88@8`:v��\�f���[:������DZ�o =���/^�|T=�V7�i>��|J�ݹ�o�R�_�Czv��75;�����1cr
q�P�o��od��7��*��Η�x��y�q����Ԟޔ6�ݨup����&�8��h��^<#58�X��l�Ct�d��vV�轗�MKN6{�i�}�͙�+�M�L���woy��R��;H �O�����9�dLꚡ��(LԵ%)����N�%;��9$��R�Vw3�>�-�vx��w�i�B��oJd��r�tt5�^ֽA�U��n�	7êv$�����}Q-���b�"�d� �箲@��Z�:�4fT�{��аӡyg��=J���F���6���}Ƹ�p%N�v7H����PP�nS�ܢ��d�G7����5X���/Y�|k�g~�{OZ�vYjt2���I��i�v���ñ�M�
�]��,;�Gw���"�^Ax6�4�U-J{v�7a
�"}e��Hwy[�W\4���[D1��-�=N��NX��ugH�Z�vm�YKbĩ�]ܻ�º�1RuwQ��X~ld�%*����n]��M���2w��]��F�
������d�w�x]N)jVP�"�����]f*W���ZT�.�ޔ���q�juۼ�4�;��� �Ku�J� �@R�mFI��<�n&����F�q^)��u,9�T��E|{�Vâ���[��HLU޵���x*.Ky��V+�1�,RvM)͉}}L����sf�����ȶ��f���f�G�&��q��ՃN^7Wim�!v&[!os�lܵT�C�ۃ�ՠp#/�� r���խ��==ȹܳ`Ey��)�8m�.l�}�:Gi��.���M��]���̫��ۙ����i[՘ڮG:c[Ȃv�i��9P��c�/�5�|�ݐ�.�MQB�=��{v�j�@�敏�8fC�|�|�M������{H���`M]�ty��,^[=¸rknuk�Z���{vf�+Ƙ^�R7���I{nMc����EYʻo����:*�h�oVuά�u���ZH]�gN��}���W6^���Y�i�@�.ow��٭:���q�20*Kꏵ�H褷j.!s���N��b����q�=GBqg� �z���ݼֳE��Ex����=ٹS�nÔ3�mC�ݾ�i�"O�J�N[��˶ғy���+,�j	[`��N�-��kv���� w9r�ɶ*�Q=932`U��ox�®��%l+� v-z�enj7˜[AW؊8��T�lrymn��om��m��sm�rt���ِ�����VF�
|.	�`Y�'/���c����V�x��|���k(>�39٘�X�[p�P
�d��]��b�V�eɝ��-)��u��̼%�&@���ҡV֕�Z�V���a����5?�)��P�͠G���Qo �g�*�v\���/��O=͵�Kw��Ѷ���q�<�������	��5s�z��\��H�fV���
�9�7���b���ґ���+T4�RǨm�d�G��m�Ԕ�^n[X,T�� �������C��%v�F3fM�DM�������S�`�zt43h��uɷ[
�tM�� �����^Ǿ�^�UPR�bP��3C3T�ULUIM5UQfMAA$��՘af1�4@EPPT�ESPSELTD�AQ5PEEK3TDPQ5STQQA0D�UUU1TDST��EQ2S%1UQET�3QMTEA1ESP��TTETU�ASLQA5�$P�LALM@LQQEISLT�4QT�%Q1EE4�TRT�2�E5A!T�4�DLD3QLD�AMD�PDQ�DEQQQPA5SII�D4�EQEIEP�4P�Nk�Sr���vǰ��y_���:�Q�-)am��RZW�k�ڌ�՜v���
,���d#�ĩ��T������ n,�rK3ы�7��?��4ބ��m��Y��:��ր����(v��<���m�x`�
������*�:���i	�_�g�
��Pɾ�:�F�'�N�izX�:��43��mc��>QU�h�d�Evا:���nY��X�_m���WZ|k�}7[�'Ps��������4o�%'����tFH����s�}Lζ��Ǯ�`�1�w�X'{�1��kt-����+��^z��q��m�J#�3Hu���=g��)���pnz{��`�.|������ri/���ͼH��{d��=�Ы����.��M�uM�\�%��.m����7g�0h��=D���_e�Z"����i��!U�ȎPLK��W<���q�1<m>7�*���#�D�dOG��v��f����L�7f�q���l���1תƻ���/,u�0�X�B�;�tI��@r��E�m<H,��4*&%�)��!�1(���^Q��
�Z�WM%>�g��y��Z4Ÿqեkb�}�ed�f�p���V�����s���oH^WTę�}_W��t�J�>�I��8=��1��szr~>��O(]�ݹ��=��G�+��z�q��(1�/�1���6��z����X�Y����?@�sW��uz�OC�	�����#��Jw��b��Oj���1�^�NҺ��������2�T)�Z�D���mx_����짚8�!���ŧ�!p�T9��q	���j��AZuξ�,f�w��\�3\�϶9�0F��o;�gZR���s��p;ݶ���Z|j�_W�3�67� ����]��-o;󓶕�g��'�D���6H��!PT�ѳ��/"�u�r9�s�4z���:���]�C��U����}�����o�s��/e���}��b�J��6BF��5~�-z����������<�N<�N=Y,�3���1Sz�xwN��\���?UM�������[�'^��s����'�R��}=v|��(]7)�aLdfƲ�t�����fݚ�l|���E�"�/(/|9xbu��G+��U��̪�xIMG���X:�d��M�{��+��}gz]�52i�[�x��e-�0��i��/47��sL��["�Qb�{NU�A��V�&������ >;�}$cؼ?��퀄�|]_����u9ns�]/s���rp���f�͋6�-G��C�="���NE.لw��3���ᵤDu2��<����fy�گ[�X]s���G���QW3h�G]�^;�V}��O'��Sa�=�U{s�¼/�碪��>�{�n'K�Tw�{&h�ʵ�vǴ�ϫ�C��)<��Py��_A���p;7<xvZp���{{���E�no;s�C�w�����N�;�&?�z{.�G�e(2�R��vR	hrIs��P��O*���Ss��9�bL~=7e���̭�����u~���u�Tp�Y{��hV�|iG{B��G���]2F�w�vo8�8Z��s~���Lf�T����[3�j���~S�㒒�	>�K�7=�[����'Dzs^�&�t�f3Φ��y��������N�� T�������+�._�U���+��t�}�����c��B�]��.S(�M'� �f��֝����0ыrĜ��읋����=��cK�k�t��4��jht��p�Բ9C@�ϐr��;T�}`G�a���3����}���y�ksHog��x���6����V,U�kTUz6���T�c�����O��/_}��W�Θ�{��`OIW=�L�L׵�z�e�la,�o����<��y�}43���[��z�No�A��w�i"��aС�^��N�z|֞{��z+��)�O������6
ٛ�f�4�*��tc�k���6�Fz_nTr�gZ�/A}���e�/��syRy�7�[�[��4v�#~�����h9B�����g�o��N�Q��R�gxp0��y��g9�L�/���uu��O�3x<�v	��}C{w�t�Ʈk�l��;�҄;s�I�=��`�r��Җ��۱�����l=��-��*��~�jL�nnbW�D��,ݔ�����S<�*�Eq=m߳5`�y�j P�ᾐH^�DT';���O�ea�e:)�m"�n`��'8|��w����+��L{1�v��0�l�۠%߲��ג�����M�m'�t��>ε�fzcU�ݜ6��(�Zp��eص\�r��#�n'�ˍ��a$�s��.8jmj��"����U_UUQ�s}��+��?��:���md�j{��J�0��j�V�ʼa�];�N̜	��n�/|�i�KѴ�c7i���N+��7�gA���͛�����kz�!�5x�i�N�i�C�����;�!��;��l���uK��rl�Ť����[����h�&��j�������x���:z<��q��I��{�W���d�Z�)��wʖv��R��L��9��K�"�\��o��3q�.-��0\�kz;��p)�w���n����E��Ht�t�z`���tұ����\2��c���Nl�����<�g�
~��֥�Y���'�[�Eo�n�=%�.�$ ^I�����8/��<`�y�yCܱ�\ӎ�e��l�1�ȃ��u ���^�Q-�v�nmgt���I�)�no'<��g\"��v;9�|py�l=�� �Ax^;��n���_ӷ;������c��+ٸ�Pa��-$R��u˖�����B�.��f�{`Q8�;��V����L:�C��!5󃯍��aD
*{iW_`ީf�Iۉf݂�mQ�3��� C[�y���x��k(-����fN���}U��[�«���? ���Ж��W�P����ԑ��Hb�����-�v"�dTM�lV!�.F|�׃mw?/j:���^]�����\����7Ճ���o�fC���-p8&T!k����9�YwPNr���I��ieJg�Ub�L������������'$�ʂ���љG�ˡ�hΡ�뮻"O	�ؼ(��ip�˘�'�x�S��D�Q��`�otonR%��5VLmщmE�T9�ɗ�fN�!#�H����3�r�no���3��oB@�7;��������mb����bg�>���λ>ifG���֜tt���	-<��λ����,���<��z
�y�K6V��hi����?t{0m�)Y��U�YQ�.��C�<�[\<O��j��1X��!x�sP5�;��vz��ˋ�d@r!_?Iԝa���V`�Ȱl�T6�V3��|�KW)�û�by�#{Kmv������>�V�=�&{G�3�x�>��:�`���.���X=l��
��Ø���{�'h�R�P��("�L�U���J�V�I�l��zn0}4&�\:�S:�^���I(����v�	�O��9�R�)��fKr��֧͑���oUiu³�m�ƥ5��җ
�W���z��r�i�e��C��evl2��	
�W�}_U}^���{�z����?���Ӏk�~]�uM�Jز��]k�C��)�&bQ�:�����|s|�G���B�\����\ꅩ|�C�i�)*��r=M庑4����)����]�Ea�Y����,+#eTeY��>�ڷ���qsLN5ő�q�ד15�S�X9k�s���3�_G2���PP^2�;�hju�kA�~��_t�:<�N�C������[EA��|۵h�:�L��)�`)�yM)y\F�	�b���l�
s��|g���#ܧ�:�c�I'*x����A��%�>^A3�ʉCg`c_���L޵.�zb�@T.
��&�&�tW��i���U��g(����
�{�t���M�iw�ps�᱗̌���MMN���`_C�%M�}fc��f2���<0ﾗ��	��6"�=H�ۖ}���S��b��]$-2�2���^������<�9E�Y>7�[�B�S����%�xN��׍\S���ΠN�Ǘ����w-�uU~%Ŋ��@nJƼ���y\�̲�S��R�њ �7{3��R��pѰI�I���$s��X4WE@�4kW{C���
��
l�E$��;{b
�w�}:=���gA�/v�ۍ̽2�����R��9�����p��yj&�R�<��8�s#��q���r:�IV�l��eN��J��`OE�)|{ޏz#�T҅��*O���;���r�9W�87j�:��>�Mk�I�-�������Vn�,��%7)�xF�Q��Q ъ���Rf�JE�w���K���=B�L���V.����i<�`׶=壥x���q�����>��e�`a�W�llPm.��{��$��3��;g����O�/S�=�/O��z�{����:��{�V�%c ���z�V�n'��<+Uu[���>�3�OZ���a�>�2���4��(��W�!}�d�ʞ��`����{Y���&���&�.-���W�&5-�oނ��-C��s��"{�לU� �h�eP�u�g��*�*U��65�z�je���,�9�~���[�]7I�)a༽^�od������\I��
U��v����e.%��dЇ>��Wr������|�y�.|�S�����P���-ϨP�c/�3����R��Xr���)�}ںS�K�����y�扖�E��>צɱ�-o��!�
�y_�}R��{4�e]�E�i��v�@dct��Z˻�L[�0��m��[�0� �vWn����f�E�t1�yF�6N��H��eqTo���:��<�5��C쏵-� ��#:]'*U�9��]Y�|fm���r���"�nլ��:�vH�����>�V�ضAgs�~mx늡��T<dR���8qދ�ґ���/|�
�r���ػ��μ[�@?=�W���Γ�5�v0��k��9d��DSܪ�<;9Wu��sZ�=md���V�N�/tX��Qx�W�V}=�]�s�(��nJZ���Sɹ8ɦ�;}Ҧ%x:��gb��+��n�j�3��v$V�ׄ��������2iEs�����f_����ۂ04qy	��]�Jg}�p鿳��1e����ծ3'�"j�J��	'��M����l�K�t�D��ŝ��`���W ���7�Kj�&��j����4!�M0��O)?IT!�ƺ�����P�o��R��������ȃ�B�i0^%�?m�]�S���v�޳3%_��3��Y����N�V��u�t�ï�C��ޯ]�6/���Z2kX۪-a�eq^�N�T��^0�z����=�r�<� ��+��|�3A��cXT4:m��L��W�{ �|U��_S�jD��L�\���NmC�6(9������~����^gޠX�������.��Τ)��S}�[�Rw�e_Uʲ�[���q��cU��-�v֔��"p��>���HeNcrs�2f��]p��7��W�4��9FG4)���q�}rj�ŒuwJ�-���2�o舚�vF�!PX�䯈�G�#��U�,m�d_<��}�y���X��Z�8]�x��4��f�����;��s��w�&߅�=Nc:���oꘑ��t���l�[�y*��I��RRᒏf>u�+3S�T'���.p>B�1pz�(k�{�v�7��`Ɨ#`�x�A/G����ڥ���`8�~���bS�j�����9�:��]�Ł�+�yh{.�M���Ǉ���1t��懇֥�U�A��L=�]�L�����+���-K]/E��r��y�%���8��x��ԏ��)�^�{P%��%��3}Y�P����{D�-p)кCں��<z�rz�m׎�g�k@ӯ8	����C���&p@�P�[J`	�y_���w����W^�z%�Q0t܎|�C�����xM�8.��O���0������ ��5�h�o`c������C�Vpi�?%����
b�|�U�5�G���϶,h5딚H�#��}���]���%�E���13�t�|nv�Y���`.�,u���^���xn5�f�K�y�j]�7�н�������؜K`�q�F����a����7`�P-=q�`��v)�J�.��3�{b6�8qU��GR
@N!kj�>O���Y�o˹�T4�Fm"�:ouo��;�=��~��^Vu�5Q�غŹD��J*���LY���v���ئJ�e��L�@���Ҳ�1r���1�E��iq��ex�c;�R2����U.�Wju��Qr=K�`2��<�:X}���&�K<k6mw}�Ҝ�e0eX��)|Ŭ5�;3��mJʃE_�9���d��Y��(�7�*��@Tz����{>d��;9���b�T�9�1S��2�i�$�r��|�����n�Ӗi�b�P8�W��0Mk�tY�X;�7t�_kYɍ�{�����[4��']�6�d�����w��pr�91��]�AȨqM�����dj�4}:H�R��fRwX{��g�J�r�#���gFR�{�-�g���c�8�e-��{]���,tN��k>��W4�����y]��u61�dA|��D-gl�0����)c���; ̦H�e��1v�\���e�P��/��kKc�t���lQ�C,`��wN+���&�kTѹ��]��q�u�¦P�7�NL��g��/��Gt�z�����yXߍU�!��ȵ3��1��ߥ���p�)ն�A��G�	��;j��O��xH�N������}�M�8A�Wk������a��0-�=�d'*.�4�I������;z{{�[�a�S1:�-J&�]���|^�R�yv�Zc�o��s^+gf����A%Wj����4b�g��]�]��9�z��:O�m�֮�rG��6dW��a��u@����B�cD���f�ġȇK�5�fA�TI��w�i�Ώ
����"���B���
��4 cE�
��*�F����V�Y���|ǃ�S��x�ѳ�%ۭ�8�=��wKyږ\��1e�#Q�`��f�ef�o�o������W\=B��ڈm�[�=]f�*۱F�[X�\y��J3����s��Nf�AGX���u�]�V`���f�v��P���,��/`��|����+6�w4lAJ�`���q�Wܯ���%wg^꧒�뿢������ɓ2!C-�������S�{�T���VX�dw��;k5u��]p�5¤�֬�h����@J����2b4��U>�er����]����[��ܹ.�E�.7us1�EY6�Z�+��Wh)w݅]�c�������R�z� �=�U��A]ghU���b4�hb�����{W1���J�݄���U�qy�B�3�#pe)X.KᏃ�b�)�	M�`6���[��&�=z�2��Q���	6��X0}���SA��ܻ�].m�����IKVo1�W�[�����秠�ɪ��0�w2LA�ELQ�T�E�QAS@A4QC@D��QSQD��SA�ED�UT�ERQ�P�ED4AT�CCTP��S4�R�Q-1SUED�ET��IT�3@D�E$TDQ1ESJPD��TRQKEU�%T�4�UEQPEQM5LUT�2ID�RUUML14�AEQA5%TQK@DRQLEDD3,TPRUMUD4UR�D�E451I%R�T�EP�DLSIDAU-ADDL�U$QPQE
��W��ě�y�q����k$�v��̽��&�
M�ǃ&s&ni���}M��86�ʾ�h:��\�q�e�/ȷ��N�6����@���L�޿��S��@�[�g)ă[1~%�F��Vl�k����{(��)yqR��dQ2�8��p:b������CB�V���"/զX�vF��\��&w+=��]C��uE7�T��Fb�W��q�S"͑��܋9Q`�}N%��̺s0�X�����XL)�z����D��A��w^:s�0v�c�̈ړ��WWA�z\7���h�\�q����M��*���n(Z�0�η���%��SpC�VŐ��WZ�C��������2ά��/����N[��m��:���_5�q���������Qaz�w�1oά$���l�����B��z�jm[��gP�S��Ȟ(zd�Td�aNf���;��26�a�����T[��v!i�M�?uv�o�藺ڿ\�3���?P��a���7�>�@�u�KL�)�c)߶�K�{C��M޿����6̊8_,�Ю��R�]���v�1a�v6]
��,%��nR���/��j���/��pN�������`"�mg.Tm��W1����u�� ��u�T�D��&$�NɎ�XK��6�gt�S��7X��*Ǹ�G�zǕ﬋Cmb��8�]Hϑ���zOZ���uz��.�/���a�]�Ͱ�oޝ|;�mӬC�:�����៪�ꪪ�,^�8��^�Zwt�>?�����u�Y0Ä���,�fT`��^ҽ�� �⟏�ɨ1{�����j��£��0�ļ��(��G��l8���D������h�9\���N�@6�ukC�U���wpQk�>r��f]B^R0���l�v��]t�^�����3���2T%Cޔ����Z��3�xGKVt��=wY9(���4��#�,\<��u��
��C��n�Ś���W��$m\���5�UO�Yn��-��������o`��Ob򳅃�V�i���MP�o'�x�ˁ�rg�k��_������~�΄Y\�����q�z(i���(b�������l�Uʽ��ޞ�0=������i��ldw��[�>��'_鮰d�t�Ui�Ps��v��_u,��b}�A��Ǘ�x����t�x�CT�F<s��Ѳ<޼��&�f��夠̖��gN�-O�i�u�W��8x�WP�O�<��-��Ԟ�t�����˷���p���d���/빯Opǻ�<zy��RF��YS��쭾��T�Z��x���w�n:A[��bR��؛��N���<����od�8�&������j&ļ��H�_W��m���z�t�9gWە�۾�]u��� ���� ���:����U~[N���z�eF��t��˼s�`΃r��UR�>�'v%�GT=�+���Ր�uD�NḊ���3�R���˅Ik��6�B�q�,�b���bX�/ճ�ʕD9�Nڣ����X��'���B����:%//Y����t�%�ޱ���y��e���9�~��K�7%iu�w:Z$����P����Z��Y���頟
�]�.�w��t��<lIS�f�8]`�|f�/�.K���aZ���ݳ����*�a���}k�j�B�+i�{��0iϜ�>�<�^����¡v����Ⴣ�m�� ���a:�)&}�+:z�ʋ�,j�*��C���@VP�)�ޖ20��r���y�C�䕷Cm�xO�R�1yh��\)2��(]�WȂ��)H��X�'�����Z����H;D΂�I���v�����B�¥3�߮��b٪R�\g��ї��p�=��|8�Pw[����dY(�y3�#$CFH����̹CO�!��6���kث�zO:�x7z�m<��}�X=�l���_{r���^���Vۓ3f�U}Ժq��I���r���Z��s�4Ņ7xVr�E]�����<v�cz������X/����a^��G�wc-�d)Z5��a����ɚ0uu;��iF6�GaN~�������r�y�[}���1�<��n��2���m�{Vv^D�1���D{��h��72��g=U��j�^�g�]���^Ip�/~�0��ro7�LQ��Wy�h4���C�ex��|�G�k�lj��:���\����51�hm)��ԛ�N���U�̞}2`�i��Z2�J¦r��=ƝM]ė���k�^u�)����zc:��:X۠��PDف��#�k�����ʦ��Ψ���W��O�D�&N�3w���f�g���gG����C�*bFtͰq&F�D3U.ǧX|�]�r�z�ݼ�{ �=iA�^/�=p�`dv��{�8k�z#�Y�f����l�x��d��˛��m�y�7�.�С\i�lnr >B��_��<��W�<��%�+v�z����_)9��V}D��2�Q��*����M8_ԭq����e=2��3^�{�3�Y�zG~�ß9�@��-�}R��
�z�.���Zl�7՝t7�e��1"7L
��^\4�`U�������v��vZ��:�^h����]�h6�yW����P��&�-~�+w�����K6�=K��M��Wǖ�������ܯ^���J5gJWD��<+_n%���2�d=cG:c���5�I78o(�Ԡ�~=�z"<��,��n�V�ex�V(`om$'CM.�L���v�pu*�+G�-�G�'kܧ��\��,�Z�|+��P��*����l]{im��iƗ�xo����ͩ|���º���?��A*��w+8Z�ۂ��Uo�<��f�XFDE[��=z���<��7!��]Z���٤9G��hn�b���-3�æ�s���d]��e�1�:��\tR��r��ڹh���ʽ�fh�z����Ab�s���UuV��2��Qn���/�o6��}�z!�h���]Q�xr�kC¼tY���L��doz�(O���p!@�暿9����=���u��=��'e/�,�����R&<��D�^�U���N'����F�Z�M�㈈L��|�O��}t-:������:���n��gm� ����=B̗�˞�q�|�b5�<sݾ�w؞�z���E���O����P��k����"�y*�Ӌ��,�:���[8'�}��9���{Nz��u�Z ���9d��1��bb�Aʲ�\H�e'�����M���\�5!;7I��XIYl���BGumK��ųM
�ғL��C����|%p\/.�a̒>쭴{F]da9���]�5�Z��ҕX �r�^6l�d�ή��V�G���N��������^s�c����䕏O�B�����W�����v�#ʜ���}>�fn�dc�zS*��֚i��xO�e�e&e��ݖ��C@N�mi��v�EgeΕ�����<�ʊ���L��S����u�=v��4�	�>�B���̼�#��p�����y4�fZ��� ���q�:�0!��"��%b�yn
�^TJ�gW�l���Y���k��~c_��	W��p��7�)�c��`�6 ����2��i*�;M��66:U}�;5��3җ���ܡ�T�b���BJ��OM�b(Gj���I=V�ͦ��ۺ�:}����v����c���׆9d��3.����Q�Q*Ǆ������$Y��ط=��9+u۝.��K���%��s��$���B�R}��/��(���b�l���ϗ������.��fǭ��k�]���F�]����}̪d�<��f����y����k$J��Y�H��4�Q��ޫ<@�����JXlLlw<�==�V��e�=n��&�W��MѺpTו$��V��i��#̼�/��%�S�e�fSYl��.�0��>a�|�]�>T�I�x��
��,=��br ��o2wjwBXН��҆Ю�6�5\8�3�Q~����fI�g<j3g�t���)
��r	�N�����;y`�(�YC}X*�"�{/d��.����ح`�'��_����N���������k��t�{��8�j����QħAB���V/�U���6��D�Nx{9���;��Qr��`݋O��,����_�hzb\e�hꄛ���_�|]MPz
g܉wv'V�%��yl};(ٞ�l:��ymuY�+���it��w�9���N���[�ouM����lW{�G͚y�B�'�Ի�p
Kʦ��	T��:�.366ܮG�k:��s5�ñ�E��{!���="�{m!�^�
~>�8#T�5�x·�솱^�����k�E��x�����(�����2�Ȱ�>צɼ�h�`�{e��C{�-i����`�1�%=�����^92!��8ݱDkФJ���Pb��e=�p��x/dO����ħ�ZF���nq�_Z����l���`�⣣���	F�^��W�ŏx^0e�OB{�~�,^��Z_�J-�5Z�]�r���p}��dy�Ms>�()�]f��Est���/P�v��I��x�>����~����-���W�a��W��<t�x=)�o-7��BNe����W�}��כ�Ǥ�C�Oe$� y�x�R�������:z�ʋ�/V�C�C����%�z2�E��_���UY"��'V�������P�Ģ��L��8wT65�+��l���v\�/{ҝ�ة�ț�d����2�h�mjAb���L��7�3Ɵe���UoQ�o�d
*���h���0E��,��*{=��G����\P��.�	Υ�%���H�Ʋ2c�pj���D:�9�K&Wx�X����� �A{\��,�������O��V\�lg��8�Ơ�`�n�t�v���Hy�W(�5Vxmb�gv��r�%:�c��~v/���mx�N�/���g�����S�Q��m�k�e�qƳ�����m���xb�[����\_T�`�R$��v�����[���qA}Vѡ�ҧ�����7Y[V4������b�3�:�S��𐺻iР޾C�.�]�c��c;8��WD5�����tͰq&F�D2�n�>��������z|v>��)a��9wz�;3-�0��,,Xs �;E��ۚ����j��X�b�S���kKZښs����$r��}�z$�9�<uVo_J]��u/6�i�&��̺��h�����1�%�)�����;��}��ܧ�\f9a_�*\J�ʆ{}p�y�ICܰ8k�{����b��.G|2i�vJ�42l��~���y�머�VEUq��U9P!r!��Zw�|�/@��J�K�V��H�.�x����f�>��P�$#o�aM�G�iyq�>��et�W�dj���lx�cvJ�!\���c܈���Ԫ��|2R^��a��R����`�K�n�� @�v�H�tb{)L?;ň��B��m��)�^]�����f� uy��{K�Z9�c*�12>n�t� �\C9��G��U��'
�H�[~l��˰zb�xD5��6�F�xΕ�c���qYϹY���
~Y�o���<'ǐ�������K�7R�6�;����X�!ϵ{�Cb�n�b��d���ΘO��;n��P�C��Wu���cq�E���(�<6�T�j^�9N$ً%�FO�ʮ�:N+�r��;kV9��wV@���/���^p��ba��%��~��X��!Pn�����Q[���d�7
iLɉ�R�{)�"pF�*��W}�,d��q��.���g.�AOj��ʰ���՞m��=m
hй���]���"��m�l}���4���\�.ٕ��^m:I�b�[��7y�4���x�?�ﾯ��[���\����(�!���8+�b�^�f�γ�T+���aChK>���s�j�f�ʺ�Ҽ��3c��^(nw�U���`�F5O�ʂ5�(�{6���Y�T)�����q�[��\b��f_��p�c�OW�K��E�o�ا��%��4E:e<7Nc���/��fs����AB�1*��`|a��T8���߆�L)*�m�
�q녝���e_O^u�V<P��,�%�ҚB����!�X{�d��mC�d�\~ٷԛn��m����M��MF8� Q�
�Qc
��"̷T[C��L��
���Gu��E0Z59`	��T֭��T��N�E�h��\'L�
f^S3�b�-�=�/J���Q��\��7%0�%߱akzt��!P�T �&&:3����k+%���{R�n[UĎ�u�����<��\<r(o�Zgs��<'��)S�3��G�Ⱥ���v';^LӋ�[~ءXf�XWF��0`�B;WsTaQ��BJ���=6�������f7�s�����k�WY)�;2��yCRȒq	}�5�8�5.��sN�Qu�VRꐥO�yU���f5l<oa�՜)n\WRL.�pN���٨-��I�ɝ݂��Ž�@o{�"���D�y����5��:�<Ѽ��`x�	�p�B�.���6U:��o^TQѽ;l:t+�\�R�7�P��aʡ��Npבq�H��_=����#}B���ɷq]�ofkl����0D5�+F�$�j��]�7���4�[�����tV��3���#e��Ƣ�D밡�UK�u�:��鷋�ۗ7Ç��re�m�[�M���I�g�#n*��,ʊ�f�����M���t�[���晪;���!S%�N���dC��5e�����=�k���M:in���*�f��s���_#��pJ��l���,�2̱�l�VM
��Yx�X�5˒�Vo_���e���|���]u]��t�H{��0:��ix.l��hmҍ��W+m�%]��Y�u����'#ܬ��}�Շgv\�c	]��W�C�i�5�Ƿ=�)�[@��zN4$�T'F:Oq�����
��%Zp+�(Rx�鼕tHڍT��]�����ҕ��mb
F�c96�!"?;��eH���Xb8���^�e�#�Y1Rw٘n��{;��@4��^��e��rQj�1��<)u+$%�l$60i+K������^���dז�).��%��º���IMB���]	�K�G�aΦ�aS�G���jd���yr+�髫I��JE�e�)������[�Ѭwۃ��նT�����ٝS��㠳'M��5��Ժ�"���l�����xRi�5��L�u���
�{4ˤO6'wj�-+M�]��,���Z�u#Ҿ9R�0}��z�ƅ�4��;��_/h\���a��Bj�YL�eD,�r�v�Qm<�w]��
�eZ{��2,R�jKjΨ�S�Dٽ����+����e6T4]�.u"��{9�Jӵ��iH�c�3
��aB$m�0z�W��O��Y)�YY�N��T-|�T�:���uڣ$$�Ӎ���ѝ�q%.}���먻�c3��r���d��:ͻ�2�xq��v��(�C��� xD�$��
�Sm\���^�ρT��@�r�+����d;����d��͸�u�^��1��jR���3��fCZsC�N��Ŭ��6i
��S�� =ϳ.���-�W����V����k�1m�I%�@���1�[��P�� s���Jmt��]\g	�d�1��X���R�Gt�o��V����S��8�yr��	L�c�}�>�����\.�FP{0	S2c(�3E�� �0X�˭9�u�	HjO)�w�
�{���})f�'������@ɇ�<9X"����v��9�sp̷�@h����ˍ�.�4$k,%ϻ������|���b��5~�Ou,A@DP�SAM	Q5E5MA4R�UTSSQT�T�EP�Q4DM�11T�Q1RT�+KASEUUD�ML�3!5$M-D�DT�DAED2�-5QUE-5IACCKT4IBL4CTD�%PUTQA@RSJ�D%A3DEUCT�E41DEE%%�QHD%D�5T�JT�AITM%D151Q1$M4T��UQ@U%P�TUALBDDR�4Д��UM-��ITP%�1Iy}������پB'ȗ����WT�x���Gȇqv�!������,oR˥��=O�'1��oM�
N�}�UU>elr�������.=�#��^�z���eUU��G:���׃�N�����e_�½}��®�ϓ�E���f̒+n�Y ������wUW�\d^G,�$���E��n��]�m�mwFر�M�V�0?'��S��]��ml��Qm���j@���x7&m�4�GK��{�x����{��,�1if��Q�����\�T[|����D�2��i�����̡��Z|���~�;y`�(�hf�@���;��#�C"}�\��^�_�u�Zw�0��#�FӬ;���:���V:QL_%t�M~/���gG^/k'«KJ�AB��@lJ]d_�����M�f�Z�<=��N��T׽͑8A+���^��̣���|�R�2Q;}P�x��V|5CA��}���5�������7��ߺ+�✡���j�:Դ��t�1�����\�/rF��A�ϵ2�� �/+~կ�
{�}X!�㡛?uh����xD6PA�;��"�lk��><7]��^_9�w��l�Fqm��.g��Po��X("|�-�{�&H�XOf��#q5�)��AJ���åVQ�M<�w{�zi����&o���ҿ&��1�F�y,VA(�]�\�;�%���x�p�Co��f�(,�&�*�&M�3����}�y�D<�v��mB�����s��}Y��]�'fP"C�%�B��9�kG'M��m+%�����'L��p�9�(���q̶s�#����2 <�q�;u�������B f�C�g���J�{C����<nJ���&�8p;�p��h��G|-v�����oBݯ%�����}�У啺��J�NX�س�r��bo�����3�I��^����dE���.^��E'Ip�����qS�gʳ��W��Vދ��Uף�B�X>h���δ�wbx���8b��+����V�8wT=����y3<7���}ڊ�s�V:�4M�)�lGH�V#�X�e�z�T�w�P�/��������x!f�R�*���F��y��z��K$T�{���}�󭷘��M}�,�p�y�;킭��{0q���2�Eg�Zw�D�f�=�(t���񣣞P�o�xm�,h�-��N����J$o���oj�8t���
l�n�Rt�x纸e��Q|�j�uY���FL�-Y'5�L��������M���z����j��-Ս�əl_����Q%to&cV��W>�
���}�XM��}�ݶ]&Eb[�P���R'��Ⱥ��F�U���Ҋꝱ���+�Y�`5�Hɱ�l�U��Oԟ�}�b�:u�C٘3b��%f�tp�z��%Z���|�v�@V�ne!��`�w��sT��*�ZΞ� A�9>�+r�DZ�U���H���R%��iÌ�D�`Bos��� �;�7�'�Ouh�C�g�.�T��8����U~��P�u��D��En�=#��k���ٖ#m�����S���M�z!�LH��4�%��՜֍�vQ�3w�AHz�������\g��9#�%r�sN:E��hp���!5���V\����X�+��A	/+���)�"��=�*��@|��οYX�\�#޶�M.���t{֯�u�|�]4L/W���|h;C�j�H{6���>��n]����ѩ�v���i>�geY��X�Ob�9h��T�}��qP�b�^+���&|�G��u�W��^��1���K\����m$/���K*S>�p��A�P�����۵��$h-K��)�B�5Q�w��B]K�!��'
�X)>^�%v8�<��F���kW�o'��{�wy�:2�WmfK��O%���p�ƽ�ɥ@��S���A.�ᩮ�Z�%�Ƞ���붟L!�n�N}�3�;o����Y�6bP�X���1V�P!!������D���[�y�(�e�wT8{��������TJ���g��v�҉���+0�N�!{^�Vs�lS�g���/#W-JgG9�!�5{�C>�@��(Wt�bg˥���6۳�i��[���vk�Y�0%	7"�OO����6r�H�[1d���;|���&�=��I@�=�{���O��Y�95�<M��2�H�{.Q:BΎ��˽W�9�(��O�lw�-W�a���w��Y~E�eƯ=Vxٓsw�O��݁�>�Ξs���Pj���s0���<���u\C�����V�'j��:�ҟu�K�(�-:�Q���&z[6S-`��2�9s��2O��F��&ޏ4��s݇�]zZ@��}�&��H_�V)��HpiU�r�����:��	�_f��c>�)���JU�����V����Q<;��F��iv��W����/�lbW(y���f*4����[PsVW�����15�����~X)3/�we���ex����i����:i��pn�*��3y�mGm��ަ*�׽����s�[��W��Ι�k���LrS�nC���!��pgjС:sb�历T-��س5
�_a��@�A��-��C��A�R�ʽ�hP��h�iL�3n��4�̈́弾\��d�q���xW���T��:<�u"+%���q;@q�x�p󋇡�L	<�dG]��OE�.S��+��R�S�~�xZޝ16�!0 ���^J�.��+���
��8e����U��h�:�������]W�5�0֨&S>ϝ�E��W�z�xj;ِ=�ű�3�ʺ�IS��f�Ɨ��+�X�T#����Db����C�Wb���w\�9� ��v#�`�Lue��Z�����[Wʱ$�|�5u�����E���{w-o�C�$k9l��|5LW�3-�rd���nw��U���Vg%
���S��b��G^:�7KU�72��-^�P���\"v�4K��q���+=�,>��5����;�W���H����+�vu��mj��,�+H��d����5�v�o��y��A5qg��l緛#�� ��N��Z����z�^	,�Tu��Vתfp��|�
c�R�2(]W����Pj���-ac�0�Gp��n���D�|y�-ک[�Χ�μk��Գ{����%8��kM��g}�[Ÿr�q��B��4���D;��^�)j�/��$E�y��s8ǌ�x#W)BӻL�{]�0�ض����{�S᭘�� ��/O7�7z�oS��磺<޸|��0�^a��X��ġ��R%�k7�ߗV�󮂫O���A�e˧~*�,�;�3P�9'22�ٍ�u�۝%�������=�z��$x�d�j��'������9}��{v�M����I�i�\w������T�~Z)՟"���K��F��z�t���kiFZ6��ݾ_BQs�懡#9���T���!��L@�`�}��:��(�z���M��۴n0��4����nmB����=�D���޺=��(E`�I��Y��z���XF���ߧ��^S���j��3۠y�?d�tzg�3�&[9x������
��ܛ;����2�HB�3�	c:�)L�5P��v8��z�^�� dž�<	v���mߨo�Q2۵�eS#iX!�P�l;\�W���Rr���Y�O����X�:'j{X�V;,w����D��F���墓��c�ōqx�|�y0�ϰ��u�]��Yឬ-�	M�#�ؒ��}S3���P�LSՀTZ1��R�����^3� &�W=,�J3&��\�Ҹ>��� ΉX"c��j��	�I���XP��u]�ۮ_3M]b	�#s�Ňc۽��w�fuoq��mcu�4GZ</�h��̺�7�Z��hwY�]� oP+e�𒳭���,�/&�Y]3��"r���:�||��)[��o:��K�2LibM�K�Z���=X*S;�*s��J���C�l��7�-xÅoz�4loI���a~K:Y"���,ǧlN����P:j?{�\�{��:�k7��{��t��Ԑȼ�M�;�fͶyh����v�#��������3FtהnJ;��(}�[yP��]�t��1i�9�=�z(�:��l�Ǜ�Z��du?s�*ޣ#ګIN������~r~"U� 4%�)V�Ty|�#f���_�����S��}�]��7.��A�c����`о�%UN�Fl�ܯetshz�U=�1ü[V����>VEC�B�*r�e`�	��Ug�a����[^^�cP:gޔ�ء��ۆ\�8ß:���ӍOuo�*��Č6�m�)R/�����%p8��3���̆=n�-j�=pÑ���(sX'��h�?X[6wu^J%�>��G�Aļ�q�h!��]Hr�ش�)�@��o=��բ��z�w������* ��H+3��h�^5R������'6i�m#i�4������ާH��+w�i��e���nU�F�8��[��
�;��rq�:.�{/5Wl��Y�W����w�#0�vPN�^��+���b�����U�=I�p�� |�]4p�_�}A2/�~C�j���g_�uv��W/uLf`��lK"�m��B�P�&c!,���	�O)ypȩxk����`*;/=cV �<Ɨ]R]C�E3Oh�%�&T"����Ϥ�$��Cm,)�^wGE�{[Z��q�� K��U���,ЗXuqi��U�Ї�R�K�hN�� ���ݥ�aƭrAN�n�u[7���}H�h%}r+<>�fn
~DG<�9�买�ኞ�����2Q�: ]m#ǳj�2�n5{�C�	*�X���f&|��8W�c�k�[��a}��z��F'�����C�\Oh�[E����՛�M���=�2�!u���k�sI�JzV�����/x\�\r�c��hӽ�;�������W��7�����[+ݹ������7<q)�׫	�n�P��fD>9�Y!�>�5`ۍ�0�6��x��aNx�b���+�>L��a�,O!�lw;��)܋��U.����!or�dRR�Sۺ=�b]x$�����Ë�w�'��}f�:���zt{8�K|����k0�.�X�j�O�ı�3vfH�l*"rL��z7���I;�2{�7��Ӻ�׽õ5hq�{�ձ����f
D�2V���/_�3�%-�]�i�{{�c�x�/� "��w���zٗN�(tuKrGs˽�����5N�Eo���f���w����`��]Kȡ� �(Q�Q+������.uI��5���L������m�=ĵ|��z��R]E�*��,US2�#�
��_�tOVM�{;,��=��;uM})3�A���>4:��QgS�X�T=�|����īa��}V�ػ����I�gt���V_[�Vt��+�Du��@ܕ`�ϳ����L�βvwh� �c��ˊ�"���,S�B��G�veu�Ѓ�@�7��o�ʥ�{Va����Uve����-U9���~G^)��X�yӜ5�����&\�:ٙ��QGE�e���]��֚N�M���}�m�@WF��;'���j�j��<0:�c�U�.���ٞNA���P�,��<+l�G�q�����-x�w�X�v�
����C 7��S1�V�xc�GUFՍ�'L�^��O��5P:2�֏?��]7�V���)h��7�uݩ:؈��W��{��{G-��'5��D�u�|o%e��~�&�X�a�Z-���E����*"�a����]R�N�)�RaL��_vz8�v��~�8�p�0��j�S�GS6��
g�c�w��mdק�s�6���K��;<PE�'�:w�<+��X�o�t�Ժ#�L��ì�>�CPf._K��D��p��ɣv���Dڀ�0�����x���5z�Eɖ�V�ҏ����y'�yY���+
V�=�xž��^w���`��W#�en&?T�c�~ Xw��"U��a����h������0j
�	u�;2��};�lk��@����U�E۶�6���-a���GP��w��[�"i��2��e@��]t��5��`g'�n��>J�AB���Z�X+�j��gZy�����慹C;'��Y}یK��pS�h�l<�;Fl�z-ښ�w:�&�.-��j�^1���e�9Ӈ�,�/}Hl�w�Z��}�@�`ya������ugȮ2��ʍ"�s��^���Y=����;�j��9�&�g:6
~���<��m�4�8|�����M�������W^���*׌)�z鑹�˱��Ǝs��I��s�t{>��@�����o���o���O�W(P����2�x��{w�!�';��,)b�����GY�ccs�����(�b�u0A*3�3z���;:�>�&	��}uS��tuGx�A��q>�@�S��۴[7� ��#��|���v�i%Y�n��Sv�y������G �s�%?��:�r�
/���kj�1���q���}�eX[W^)V���MvÆQ}S�}~KM�|s��|*i��f���+7� ^�l.[�v��r�m�U�霰D9B���7#v8W
�V�</J���t	H�R��t���l'���Z��R� bm���YWn�\`7�l�n]+���8�%7� �����P�_tw4myT�����G��lm|��w���z�n��=A���jnw.*���:C���l;��R�3M*���=Ӏ�c.�T~34K=`�9�91�\;�`]44�&�ȃ:�θ��-E��:�!6��y���,酹���A�{ܺڌs�|>�nt�4�7�mk��.�SYCMy��V�`�{��AS�����×�/]q`��L�`6ȥBK�5PR-�.�,P�֝�Ki_Q����fm�u�T^��Z���|�cᆶk��ܓ�f�	hT�R]���`t��*���k#;$JBgr)^�q�Yt� ���X�}*�A"�!��>b*�K�^b�R<=nhޓ�)]�ӈ�)����6�X���5*(�5�k��6��U1��6J�=ٙ75�Vֆ��5HY�c���t�S��V%�c>�lF{�Y�H��f��f��ݦ�kM�s1��k�u�s��*�(R���sD;��N�(a�'Y���Ա�v8�����-����W�;�.����[W}��
H-�à��{��!o;Z�����#��lhі�қ��xتz�����Q��V�d��L�7��Rs=���:�_]ѫ�12m"�743̓{5�8�W�T����6������[D�����?�f��4�-���b�_`EE�˭5�X�A����ӃR:C���$���e�R=Z���}�lԸ�,��R�*�:g��5nu�7�	�o��<�o�`pa��)%�k��w��I>:&����#Z��竊Kf�;.�D8m6�����Y,�l��]׷C��w~t�@ok=�U1��a���qIj�U�%����1�3\�BV�ml:�	��쒧J:��!�@�&��������2�G��[р=�������[�b�T(G{K�8��8L� 4z��k�MXdJ%ZP#�a��4'h��WuIF�k������m����z�rX��}�A�0HM.���E�LX�W�(�Θp��&Z^,f,�i:D�}Rd��yN�q�oi���`�F+%`+�t���-���`���[�V�hƪR�,�G��w�D{Th���F�V���6Ɲ��w��z�қ���[�w,�R�uX�{�|��[m��lu�tZb �JJ("�b����&�Zi��()()����f��������(�(b
i*h����)��)J�U,IMP�`R�KSDQ0�IE5T9�4��RPPRLCD�5IAEATM%P�DM--1IER�d+E%,AE&`bS@�L�T�T,TRDҴ�!H�DҔ�AB�%SUP�#MUE5AQHP�HV@d�E	ACUAJR%%P	@P�%P�UIMd&C�����D�>���/y���sM��.!����Z�@;��I7�"���y�=��M������Y��E�ƌ��X��Jv"nJ{���i�p����,��7�D�"��
��q��j��S;��x��mdt���	�kk���P�sW�1���l�gI�p�E��������y3=մ�2��n�����N�gg��~`�b�,O)X*�>�I�#It��Rip��bƸ�s+8����v��e���)�Q�vS![�T��Q#�ܕ<��f	����%��z�q��2:$z���>g�z�f�-N�[��53`k�Un���\Dۂ�&�t�ܛx&�^��&�X���lw�z��]�h�m�!��l~:o2�6,�3��@w��F���p��%҉��`�ʃ9���2S�����#�5��e��$��m\#s�a�[i����<uC^➨���5�C���Yy�Pf=��!�1���	���uN/1�U�A�uj�<6�x�p��d�tOYN�@�U�C��&�g:C��2\uU�W[xJ1`/<�'�2� ,%�x<��e�9�r�S�x#Kx�?A�N��G��q}ŗf��ܺvPz��ch�Q�v�nf�>�;O9|��lX��f�W���Ƥ��x��toyӧ�Ԟ����Գ�3[���?!�����Ɖ��S{v�4���pt�LI@�s"��>��d)�g`�����L��:C����֤�����u�+{
�>{۳���h�pmL]r"�Zf�l��I]��q���b8��%"����ޒ�����"�{]Cm�$�����N5=տ��W�SOŊ^�粁�<n�;�݁�(����ԫ<)�%c]C=��a��>�9%k�\Ӽ�x��jҞ➾�܍��7��#����ຐ�}�>I��9�������b0��!ȰA���>�1g�{���� }��t�g>TxR��U��z���x�|ؾ��͞����2\Q.̄/��	�1}��Ob��E���3�=�	sG�K�|��Z����\vAԙ���K�}�S4�BR�=�ʄ_ҰXy'�$/��m���3�<�$�7�R�]T���>�r����Fj���Oy�Qa��S�'ܫ��b�%Q����_'k~��a[���G���P
M���e��T>o�Ci����+9�V`.��M�~�Wy��T��B;������C](jh�����'��9�T�*%P�b�_�� 7򷉸ro��W����E���X�tC��ZDQ�z����V������wN��(�{��e��T��5L��~̽=�0�ce��o��y�t�K�'u�����vi�5i�|��flބ�*���s�X���Z,f՜�RYc"��Ԇ'���NmoE�33�&p3��[�#��Xq�9D�iOi���S��X�f���쉋5ۑ�8<ŨY8���~<��޺����={�v�8\�.���˦�&o<�����	�Φ��3ƥ�oe�,ɍ�m�@{�M6�	[�dz�;(جAh\22�2����Λ�Zx����&���.wg<�=CS�������U,�p���+7{�k�I��7�]��)C�����;ɘ���,
w1C�P�'S����+Ӑ��c��c�t�yxi��i�Uu�E#@�(P>j%x����a�\ꅩOS�:��ac�V����>�w��ϲE/jR]E�*��,��f}uDrO��GD�f���'��P��]��.��o�b�=ZxưN5��d�ZzL�Rу>B���.\���*�j`SK��
�*vB~�ᳺs������+���ȇ���׳1IQ&	����)����<��kF�'Z���j�i2,�^����`S�
73���	��	��X ��I�g�c#5r�%�Ȱ��/o�m���ڏ��[�Sƍg]-{[95��sSKL�I�̻��!��G��z$�ƃ��(S�u	J����W������%�d��Ũt�����&�ϼ�m��.�Y%s*�X:�*`7���y �����+�g�������hS�#��l*�=!Ӝ��޷�Nw �V��~z({��L������$�۵�`�9z���^�P�خ�avdȮ�;=��3M�\�ùW�t�Ͻ�����l���@0J9a���¶�G�q��\�]>�^:��V$�����I�«�{\ެ�u�;�'�q9S�``cѯ	G��}�*8d7��&J�V�<�,�CBLfhw^���gI)���c���)5�`�G��둉T:ɳ�5�e._K�*����M�Հ��7����6f�[Y��UΘMk�I�-�����;{��Ob򳅃�G���J�5��Ik'tAޞ2�9hnQ��y.���s3���ة׹և+ǲ?=uS�mx���aˋͶ��q��JŔ7Օb_۶6&,mqv+�b����#�G��N47��^��њ�M]�Eg���e���a�?y����''�R�������ϗ��Rޓ�4�ÙqY���	r�@�B��:�|G�f��ޱs��}9�N�р�f�:�����v^iso��d}�K�M�@U��1
n��">������@��n���jە�6�滖�(���yֆh�ha�o�����N��[g��.����Mo��}�z$~�֦:�o(+NB7��.�k4<�v�oh'u�ܸ��׹��s������j��;�[�g/��I�'SWz
gܴ�����Wn���:�Ȯ3�,�/}�%ѓq�e��������i�Bj����4$g:6
~���<��Cn���ğ/\�u2��MTr�h��	-�t�*TJ��L�ͦ]�1�8ѧ9�qϫ�]�w@���\~��{+/m�~:F�]�r�	2��>)��)��;����L��.�Cm��M�1]�Ss��E07�ɿ�9h�d3�`!C�����SQ�����^&z1����{t�5�m�n���+3�f�����&|�
�~�<s�N'���R�Y�^���߬�{��gW�Y��=Φ.&X�Y/Eß)����#�X�\):K�,ir��ܺ���Yg�A���X{S<�T�Q#���T�R���{i(q1OVT�>��Y=�&��j�$=�-"W�ux�H��y�P���2M���&�	��BHs޼�Yx
�����&.X/-��*�u-h�.vh��&�7�!Дj�<���oB��Of��;nع��7f鈸���d=S�0���od�h�Or�����ӽ��4����A���9���Q�N[�-�݃��"#��VVp���zv�9zGS�ּ�9���ˋO˷=�J�n�9gTh5w�Q]=4_Qn�6����W�]��.���U��fsV�c�ج��l�+u@�����dV�����ȧ}60:�Z}��+��j��f����H;��+xcw,T�co�|_���m�N��T�$�x#�#η��}q���[xJ1`/<�NO����]�xs�{y�"��� �Ǭ
�x7@�9o�Buƶy��e�OLl�lQ�"�qY�ᚼ���T��6�ԫ�#�����D�*D��ȯ�?`z9S���z;�����Ǹ�k������\��EV��ǹ�Eky+����Ļ��Cò����S�q��{�ϟS<�=�r�Σ�x:,��:�G�u-��26�#�_�.�ϩ�%c]C=��a���Q�(sG��r��S,Q�]��U�x�wZ,�ن������a8��ߪ_j���5o�B���ow���r�{(ϻ�/>���Z'r�}.�3%W"�P�,��d\�\�?,��AP.%y[�#�Ū�})���s�ŻR�>VdC�n>s��Ͻ=�r�iuJg��
��;�o6�>tP�^�D��]c���Ѭ�ȱ��.�dn���$�laNIeaϴ2�n��N�r�4ߖ����N�<ogI3�L�5���gc��ha熯J׻2�=�yAw���
���4���
U�� 4�f����'Lq���j��7�_a��n�������κ�ݡ��{~�%�&T"Ĭ�`
�����p=[��b�H���u[~nƺ���
�U_+GҎ��W�9��G}u.Ȇْff�#�s� *�вϑ�:���1�J�DR���U���+9�V`.�cE�!��k�M\��"��^�0O�!mi|��i��R�� �"6�5�UU�ꌋ:�:7\�s�sl��4��s���^ۑ������CP� <6�[<-��W��ǣ�yY,W����Yy��R_o��Ŋ���V��3�N�����(�;��YN���e��18䭧z{���R�B$A��8�DA����&4{�755�;��wʄD��2!�κ�Œ80W!�P�h�wI����w����87��8=L��a�����0lw;��f{����NJ[�,�n/��[2I-�*�]
P�t !
��}�Lŀzٗ�;���(a��.���:e�;U��Bk;�~�v������}k��"���X��5�l�eΩ19[Bbٸ�4�o-��Tp���s'cI��N/xzy���$�Ӓm6����&���u-)֏3w��V��ޒu��b�0:�9��2;#۪7c������ԇcGx;m�w�ɑg#�_n.������yyx���$��C�վ�!6#�����1��!_zJ=E�F+�����\&J���5���fe��>+��������@q�j���yݙ�P�Y8��q�=�n(�����ڟ�T��we���G⟭���9ԯ�ϴu!��k@"_[�h��s�:a畂u":����$���|l�z�Y��'"^�����5��r���N����f`S�
73���M��Ѓ��B�gpg��>��=���`�'����/��8:ɡ���Z�ܫ�u�^	��U��߆�Lˍ�u�s���x�֒Em��|���톡����fL�W[���*�Q@[��U26�voEY�b��l`Dz�|+l�|7C��̕�׎���V$���d�⼗d�.gr�V{��Е�CNT�d��uP����ȑd3����2�g�&����U��L
j+�u�	�(��e�U\x���N7t�j�;�Xށ�=|�C��!���[�۵Sa��a��;�?X^��h�v��~X��@�~$�.���Nv��'�yYI�R��יe�i�m����沖v]����V��Em[��Bo2It8	k�n�":����������y��m7��nLz�ZΧ�]�q��󡝸��;:[lIf���"�&�����K#\%��́�tZ��7i�(
�n�*M��`���v+V~�,�
Z;�z4�J�oe�[�����b�{^�[��ǵ�e�d�֫oԶ��Iس>��\�w��YC}YV������������f*.�g�y>�Rn�E�@�v��u2a���M�jyv��;�͓U�\gT(���_�W�{hX>���a�ְ�-[�ke�s�`0��X�=��Y�����g��x�ǺLu{w���423g�i����5GR�h��wɈ���<��UN���ug�R�1e���Wz�j�Ȧ����;��6�H��V�_c��g:l�ձ�x%��Ω��3Z�s�j�F�I2���+�"�z|ֳ�)yq.��U�\9�;&�Nx��}X'z��/���;l���5��p3他�
�쾴ʉ��
S=�<��'<��L��p�ɀ�qp��'��sO��?U�puW�0M� ��ߐ��X�4��s� R������-�9��0�!t��/L	gv�j͖��4�h_K\�U26��Ϩg���N/7$�k̥��/I���u��h���J1aZ胖�T�lMġ�e2&a�F��}y41k֍��ʈ��Ų;A̝,y��l��7�lua]e$0U̙]��.�Mm�I����؊�ʑ�]�=�{�#���\QIC��
��G;����	���(P�~��k�#d'lWF�'�}/EÁM����#�(��I��ې��Co��/\96`�gӪ.�z���>=�f��$h,	*yeL�<��%�ؔ�V=oS������~7p]���z�ú���H��!�B�%�����D��&��KlR��z6�^'s���ht�+�&����:o2�9�-C-X���^^Ҟ�>���[��b�ś��S�L�^�l�%{pd���_V%�*�e��g�m�3hlV}ӥ��9���E<�:�\��|�\�E���>�ȃ��c5O����t��ڼC�T�S��m�����������|Pv��U��s�F9�oQ��P�\�v5�}x�f�et�ʺ�����]�W��C=�L�&\e�\�F�a���� �t��A��������^Dg����n���O���s�����DN}��Kɐy�r�=CG��N�Ez��'���ÇkK���?K�)vN�J��3�/X�z`��񱎢W���6�%�0�:�s�OuX�R����a'3´���/�2�c.v�;X)�Ru�j� �.�F�,�U�h�(wjF啦���14�x��z�Zդ�>��@��?u�H:�t�f�t�oJ���v�&p�Pk�3�������H�㼽�
�\ǹԯ/���mJ���(9t�碨��Xw��J����	��ՒձSf��ܮ����V5�a\���e'u
���{ѯ,�b��0G�k���}��;Mr�XU��IR�**�e(�b�x�z���_Eo��t���J��������Q�v�ͬ���;��F�^���;wArw�U���-��%M�[X�.]
��gL(���V<ޭ�l�!�"Go �+g�97s�뽦Fي��Tb�8)c��"��6va�o<(�`�X�v9ut�U�ν( �#�9\W�.���vY���!o<���ͬE^�)Ѿ
\p
��WaĪ�q`]8k}P��K*U�X&io{J��]F=��p�h��Nh�)*�g(�)���+~ҳ�X�|1���LR:���ѥ�*_
*n����qc���6���:�w ��N�t�޾��*,�k(��F��I�
�j�1j��$���Q'#㵭ަ	$r��0��nm�ό�޽��7s'9���SO�\;:�j�v"�سK]�t�t;SM�Ys�g;���#ky��bۀ���L�o0oY�Z�>��4޸ܬ䖙������I�v�V��Uס��o�,Ϛ9m�V��Jƾ�E�K�Bs	�1�1��.��,'z��`pQ��=�EMg��Gk��+(Z�\6�+�j�T7)�������ŁO��9��@��M:�+��^`(C����=�>w��<�Hj��.�ۑ�ikXN�@Y�۵Ѷ ��o�׻�Vq=wJg�J���3�nZ�>���CF�uTbʏp:Z�!h]Q`�uql�48:i>�V�3rKn���07q]~�R#=�N��U�O�k��x3�:��a� ]%��sM4�Ԏ|�-��Bc�����gM�,?��W@�}]�ժ.���^�9�a���6����-��[�����Efn�-G�Z̙E�^�]wK7��;畣'��H"�k���Ong^�jq�vz,]���I���Z,�U����|M���"���8�a��nc�]_B����R��L���f�n���Ѷ����0{tZ.�V^�ת����j��V�iVb�9��8�7)���d���к��-/Y��'�-k\��VC�X�M2����v���$���Ȣj/��ڕ��������{�{^��T�{+�[܈�u(^�u!At�����ܹ5���gAU�N��������ի@�a�B�{s�v��U�i�ܻ�r�$��{�+��I�{��N�zw�������:�,o���+�U�#� 1-�U|����#|j��j�t��3�ٻ�e�S$�2 (�,�*���)(h�$��!2����p��r�"�C r��(b�(�F�!L�31
@�
�r
�	�R���i��!(�30J\��!2���������
�i�2�!�J,�
rr
@�\��� ��2�hD��"*������*��2̐ɥ,����0�i"\�)2�r��2�)2r��h2hZi��ȳ s1""B��J��rh2'���e�n��{H>]����>gC��m���|�;�܋�)Ou9����3H��9��Q�x��Z.�����}���`�
�w[L}����{^���q&F������|��g��7���/�F�rFN�F�@`+/K�P
���o�n���#��.�:�K�X|����bc��*�@q�9[ر�K�/�f˭�d�#͌���h�.�8T/�>���>*��ʝ@�z�}����7��ӹԚe�9׎|��ہ;_
��d"�*$�O*UP��g�u0�ܼ��عS������K�u�y��]3�ߚ������T#��B"���yݣwM�N ����5a2}�\o�_ְ�U*������Xj�-<¯#΄>�P��'�6���su1*#�|�b�|Ϳ-�]yw;~�|��֚��Ya�0�Q�6�pn��*�d^�/�j��yk҆�������l��'���K�M4f�B�Fd\u�^7��Ueg��U��bg�L'���̳�-#L��q{
g���)N��KZ(�T���%$)?pU�,���qy�RN��Uo�l�,v\���(�;��YN�����gWW;��Ѯ�Kf�,:0ͩa�4�\078�Fb1�5�:�77�:���V�VU��Vj�)!�� k���ٗ;�Ǖ8\>Su�6NA�v ���Cfq7 �����`.�߻%�ʉ�� �ʸ��ޛx�E2
V�KU�Hl�S����^�i���K�s̘����z����J޳"�V^��ͺ&X�|�ƅ�8v�]������H��3��úK�lu=�c%x�v׈f�P�xes|�-ayʼsQ��-[�U�l��^�gS����XҦ�np�U�U�u�p���:��[��vk��
��&�iP�,S(5���k6ه�S�Y�ߧ�FU�0��b�<�'՟'������L�Q{���,T��.�����S�N��dн�������ƞ�Uoge�jk>�q�'��&�>u-0��UL�fz��ԙ��ju*z{����!ք	�{[���߻Ee���΃<��׳1rTI�\�*>O��V��{��Xf���\�D�T��ؽ�����:ng����x��j�,3{��-Ԡw9ǈD��7�g©���UNrY4)߁׊w�ۓ<���=�س]& 2�[��8���V� R�{��1ӎSu�]_��u9/<�`�uxXݴ7�Q��7m<����Y�&b��;g���_W��P��yt`����P�Qe��>�K`���P�N�c/��q�GW��}����T�Sq �j�]@�^�\�X��u�m�݅R2ش#[{Ò���R5���V�=�ݖ؏n2�Q�n���5z�Yj�=K^����6�uK�a=f����H����n{ͷ]iVmJ^�0�}�]��vf8|]�����'O��u|��J`=D�6>Źu�"�v{����\�_�߇O���i�I.���V9؀ؒ�Z�w&��$D���c��2v��=��9��Z=ap��͐��jn^�,�۵q`�^*����I&[�Z:Q�;{����i{�	`��m��Y��u�]Zt�&r�CmF�o��Xg��'M��&#�f����Ӫ��ig@�N1�M�y�;yX�Y�Q�7���"����lLj��]s����x��6W�q�<��S�]�0v1��4ٳ%���^f�:���O���A��b֢�w�u�n�r����v����@+�1��;~[-S�:s�!f��ޱsƺl�zݩ�,��C�:���j��ܻ���g->e`��"����j��E���m��Ô�1���G��@恓�܇��K�OXʑ#��ڙw�v��#9�϶
~���9VD2'�.���(ɕ{��o��ΩX'>�qb}.	���t�ҩI&��ܵ%?�n� d=��J;�������ݑ�f�q�v���a�"�cm�uO��r�><r�0���,'�Ձq�N[�[C�Eo�Lvr+2�8��{��Yat��w	=�#4*�%��\h��R�{-�)�Uf�dn}�˼~�4s�s��ϫ0D3��q-���nonQ���2��!�i>[�(s��֙υJz�)L��C����QX7��ݮט�f����7v�vA�S�ޔx�׆�Δ�>!���!C���A���hE;S�9g������EP��I�=�c������nC���4�h_K\�U26��gՐ�a�t�Һ���}���N��������E�4�1pٖ'�K�p�i+ �H�WR�������]��y{o|�~,x[�-8��z�p=�Ʈ�8�<�S�K�<��+��ֹ��v�x��R>#���Z1��R�]����wȂ����r�S��
d��D�=b�YI-qUm����+�m�BĢ�U�A�ͭ����Y8�nw�ɝ�ݎ� �GY$����O�X��ɒ��X�^߇!z�>yi�U��W��W�X��V��z��g��*�_���\���6�=�B�� ��^�'�7Rg�*c~���˱J��Ou�7���:۰b�����(`��l��l7���
�9%ϔU+R��P��O�-T"���7��b*�9s�����o����01��)Jb�ZY�J���ejk S\��3�"⡙i����[�s3m�\���wLb�:��;EӪےU��"�^9:�%V����○�����MMfL~�t^��O�`��=+/�Ҟ3L�'\k�'��:�j4V�A�2�/TP�h�0G>��X�r�U�0j��D���D�z����ʛ7��>VEC�Ok*��v�1W
3c�Y�AՑ`��G�z�P�˶�D��b�e�,q���έ�i�}g`��jIU��\=Ҩ�<�T=4
�H�a�6�%����\��S�J��P�i�.x�ʪ{5�Ђ]�&0j�zo�{�)8�4�;E��f�
ir6T<lK�M�l@�u�)��fz����'�=*��(����[���s�[>�H���eB���dl>.��r�"��ˮ砛C�Q<}�S����:�et�vev,s����@��Z_�,9[�\������3�:�7(V�y@��䴈fmw]3�֦i�%�>�P����Y����S�����t��i!$��X"gۗp��$ϱ�Z�Sˌ=a������N��K;Jy�#�/k��y� �er;o{�$�!I?a4qt;���[3�ǌ���BE�9,x�u0��m��	�"��Ko���u�N{��&v[�Uv3�Ls�cܸ6�iٜ�V�4�z�j�����T�k�Wå��v����[���(ج�������:�7����~�S����yY�'��m��-��Ҿ��2��`pW��:'b�F��L���,�m{�xy�&O	Vs"�(<�Zc.�g�O}�]+�0����M�`�13僦�u���b�z}CP�(p�k>g���1�nS��)�r>>�]g����[�t�%FE�X�;�]T�Nΰr�q�5�΀�/��ʿ�������h>�^�L�Υ��qԃ{/=�2cGnj��uH�ɂ���kޫŷ*��p0pyz�F�:V_�O��;WvⱝVX9���fu9�wzX�C6;���/34\��ً'�<@�7͙�Y�UwER��;([��V(0B�K`�&b~�eӹ���ۙ�o��2�le��9Ծ�"{:���h�s"�>諸�"���
>j%c4�b�R��������7Ϥ7�ʣ�D�v�y[�h���L9.��r)��]�PߖUS2�#������}������*|Fꚰj�[��g>jk'��3�ƴ�I���RуP�+B�ǅ�>Aܠ�PYz"����k���_g����5x�B�gq���V�T*{]�� ]s;��jfu�������Og�3Mx'�)��_�����<:�?k��ǉǑ'P����Y�,�c�h�j��uyu��^��3M��U&wc�fN�O�ss��6}�ll�*�i�yo�_¸r��(��٩�ze`�H��v��6{�ɚMIN�՗[~>Լ	է`��C/)ډqt']��]l��Nt(ؙ���fS��~��=��TT'@}��U�Y=�z��A5Ⱥ�ñR����j�0�}2j|/o�/�A4��]d�3v��G��X#.����p�pE��})q^�/^]��dӓ].�쓱%�_M��k�^�烙��Yo�@��r�_�3	�xm�
�1ƥS<6ڮk�õ����^��V�L�:��ҙT��<�09d���̺��IL��0�}k8|3�;뻝��*��4�R����� eR�C܃[��R���M�Ѱ{/�{t:%�v𐵡ԭWA<k�&pӵ~A�߯m�sv�,+�X}0��P�<����ri�U�q%�sɵxP|���[�m��+"<#5l���LuOV�c�t��zLG�����Ϲ�W_�$1����ǰ7��	���K;Ջ(oVU�E^ݰ~ؘ�ź�f�I�jeQ�Wz�2��^�W�*y����{�����X��n[�|#ݯ|X�k{�R�z�AMÛ�<.Ӣ��{��w�dڷ۰�3:���]���`b�	5J�]=[7�7�5����v��н�%��8�}@�:�[3��yǜx{������Gcl�M�2X��Ƿ'�U	ڦ\^u�r���P�
�	��H;�R�ڥ�N�x�CT��9���#��6�hze/.��$�/!�Jj��y���$�g��>j}I����-��S>�C��ya���'�gNܳw^mr��͏����sϩV���ɖ2�H�A���˱�v��Άl�ձ�w�J캽�����GԈ�TI��'�'ȭ�y��^\K�.r�p�;&�2�碵AbH��>���-�{6��k	��A�z��ٔ��'�p
9߆vR�n���S�=�Ps��OA�I-��X]�.�8�|�����K�o���7��6M�KD�3�!C���h;�Ҏ��e�z���]]:u#׳�u�$v8�����	����
'~�� �κX7뮶n�����V�r�8�Q�[ș1lۣxk����
�:6s�*b�.���K�p�i+��H�[};y�jYk^%j��*͊^�(5�b�^W/PֽR���{Wp#A�T4"�fP�Yxy���vGP���G��*��_�xhr)�K�K]l��e뻡� �߅�۩�{Mdfʾ[���zr�=�� 땽�J.K �#���ĮQw��ב�B�1L=�t|��G���������yݪP7�+Y��`�e�oe���F�ཊ
u�חp�5����lt���fCx:��M��Ig�.ZА�t��[~4ضMfeX��=,SՀ/.�߅��p�j���|0�c�Wd�w�5�_����;�dX}�vH�d-l�C�J�ޱNV����g>ն��W�ղ.�]����4o(|��cy�KͶy(p��\h�g���s�Q>���^Y���S�t��eʘ���T"B��9�=�z'T�$�x#�!��}q�W�rz��TN�ǒ<](b�vw���J�.��>^0�������n�̜�C�ڟ�$����.�;��}�G]	Y"s����r���R��ʀо�9��Kɑ����i���k+b��b���Zl�׭�mǛ�!��Ɵ|G�y=4]�x�:�kPŕ�X���*���J{���:O9��p��V�P�U�|�`���	�UN�,j�x��OCc�L��|/��<gỵ�P��t�G�ن��SK��T<l �y!�;tгF�~:TCQ�Z|!����tVȟn���(uM�&�6��S5[?lw��t�^�G�����یT��l1��P������c�ު��}cYq��%�B�"�5���⻺B.�]E�u�MEBJ)t׽�9�^k����N�
]�9.�]�ou�ǻG�	��J��NyG>���^9|^��[>�H���eB���e��/^���{9�D~�	h9�K=���fg�s�92�m��b�PL�B�Q=j�n
IE�m؞��9dY>�kEK���g	�3}X:�v�3Oh�%�Z�z�?`;;Q��L����_���~Đ��m��&}�wX��L��:�]m)��=mUŦ�37��T�Q�
���̴`�>��!��b��m�h���w7���֘N��+�`׺u��o�5���/3Z������J'|%a�	h���m�H���l��'��Ԓq`�����Kb?�yЀl������_s�13�0����r-#L��q{L��$TT3k#�y%���_���v	7��9J$x��Y.2/<9T!;�]U��3�Z����X)KƂ�gok��U��xq�>>�Z��b��[��\�N75���[�U�}�'l��/�U�Wj<��o��,Oe,�1�߸���8�}R#�z���9�wGK�1�-���L^X�tN����6��ԧݍ=�Х���u��`�ú�Vݑ�w�shL7�d#���E�>�f��fp
� �
��
�R���-���zJ�tT��C�h����]��ܓu�\�mO��%#����l�`h��_�Y���tr�ܡ��O��t2-�3r�df�w�ԗC���5\����%����鞔?UE��z�⢽P: ������Z�Q;�&:��
��vĤ�弨*xq6�B�9��6|mT��:���q��Z���tu�&u��Vt�c'
C�y-���h&�ǳt]r�-0�#5�+,Y#�j�ʙ�Γ�jÚ*�e��즷�- �m��`�U�*µ�����V��u�}���9-n�S�5�7���ve�ٺ�D��ٛ7�)��IvR[ם.��ǐ���WM�ޮY
����I�s��Ђ�uk3k�,vsb/T�`��~�0�v�.qV�2��Hੑ�����d�
8�'k+��x��VܷA�[F�Eo�H{�"�f��E,o�]_}B�����r���$����WA�yP��_?��'�vK�~��C��G��zq]�Lc�#�V1�#&�������W���e��*V�;]�ݩ�#��_�4o.�m:��P����{Xes}S�{��x�ح�k )U�vk�Tƭ� �4a���^�3�-ko�KVi�'p�:�������Ҭ�ا����a�35DS�fp���q�ڻ�ˡ�c�f�u��'T|�:�k�6೉��J:p�ҩ��/�U�쭅���pM�I���m��\Vk
wS����������#|e6�q�5����;ܬ<Ҽ��z�y;]����U4�s�ݔS�ke�����&Oz��J=<r�D_!N�v�
����K��G2y�u���-7O%�
dr��p��l�t�V��Q4@�O<%Q�hm��o�s���Vl�Z@<-�Ѷo��vq�ہFԳ*�P|"��u�{:`���u}��M�O`m�t�f]ܨ�]���'QU��f�!�%i��(��_uM����X���Ĳ�cp)Ccʀ��f�$҂��pS�>��`���,0��c-�8B����0qXoB���J��(�����#l77ɱ�占�黷/��RTk��]�x�͜Su��0uev�1��re-Xz�b��v�`�Qrdj��C����yF֖`!(�&we����͛�����iR�N�8�]�����!n�<U��2kj��a�m�S�͚ഫ�E7lNR������yGU�W3�<WRڍK)j�Mt����\-6�.�.���Wwj5h,�a�����+�PVk��߅�B|���$|�Y�.L���hJ,5�g����'�dѪW:' b=�[wf��˧�v���v��7,��oqm�H�t{����q��\Z�AݰdGrL�衱�Ӓ��N>��V�T'��^�~<��~��rJ��
� �����,���B`X���q��1�r��(�(h( 2L��!J3',��)2P�0�#
�
,����2J#3��K0���2(ibr@�2r(�X��(b��02(,�rrp�&��)C 2A�
�*��Zp�i2riL��,�2�2l���� �(2k&��!�2��,���'$2
*2r� �ɪ�h�#rJ��S J%)2@��"��22S!Z�p�,Ƈ&�J�rriS Ȥ�)JL�	(r����G'!�b+�+�+�*���w|���P}�a��_]��:��W�:�W�n��W�T|��:��Ӻ�o�S1�� � ǻ�-�=9�E�o%�Ӣat�;I�*?��+ǻ~s�q����^85]�մ!/N�)t����i�cLƱ���kFM+�-5���{����2�t��KY�T���]K���{	Ŧ�վ��O:�e0"��S�➜����B��֗�"K�`��o-�U9��wl�G��~�=v�l�3�XVFϪ�*ȍ=Y������8�<�����Z{$�Q5)6�,彄�0f�k���7�mJ��n�ćZ�t��t-��Vn�:��yX'R#��V��~@��ѻV����0s�)�g�)�e;SW��uؽ��٘�:lL�{���VY���c��ǚʻP��]y|�%��8^�����[��jC�RwiĪ+��e-<�霗����,�&p�+�/ԟ/^]����^[\:�=G[2�9��y�0)^:{CYs�dg��0�U�0�OM�`E�Hö�0�}��кH{��s�J��0�ڃ]UU�:�v��8�^�|D��u=���Vc��@���۝��}�xbd����	��W/�Ϙ�G�D�f(��}�\�)`�~���0���j�c9�u���t�vn���R}W�+�`�9S�t.nE���묎sOĖ����H[��:�;��i�Yip�T,�n��V��}:oPn3�%p'Mc�e케�#l�{:]�Q0P��bII�KJ>Reݙ��S_�ȬN��T�.����כ�r�npn�űiO�ɧ����re�u�]��:wl��5&����"�d�^�Jӧ&r�j5�o��=Zg(@�݁@�n�L�j����dM��i�9ٞ����=b�ƛy���`��1�F��˞�B7�`o".s��O���iJ���9���6I�o��}�]`��y�����P��f��#}�	�ty�mu9���`��r�+�q|�S��3[-S�:s�!f���˓��s�n�P�h*���4�Q����2��M_�lb��Y���X����K���Ԟ��NL��B� �ȭ:]���z:��Oo��h�>Z��H��?0(�>�A����c��g:l����k�GD�~����Z�v�4���n��uM&�/gԫ��u-3�)�{)�����������_�I��O�qr�D��ϧz��	ٔ��	>[�(o:�Y�|z>\6��%�w���&d����b�9�u_���'m�Sy�1v��v�8�yLH��إO9�-�xr=0]-�ܙO�A��vMk��������9��$����v5 xA}�ҡ~ʄ�t�YX)��\�V��z���}k��l�<x�JҶUa3�K!Ñ�b�����a�o��h�`�{HC���A�ů�ܴ�}NM/z
;�j-�{���� ���_\��2���p�__K\�U1V�u���n�`�#E����U ֋��[�y��׶�ANs INخ��2�b-Ɉ��UD��f��Y�r`6�oa�C'�
M/e�qq�O��Շ�C����G��%O'����`v��6Jx����I3��z��q���"��z��wT7��[��u��̇����n|�jz�͞���҉�vU���Z��X��*S;�M��桔�S�5�KV���;26�'9�~���Ɂ�/�`,�B{=��G��Atw�>J�U��`e2s5����G!1�.k!��Xf��|4��׵hA�e�A�s��B+�f���P+��;
ك]��ўۀ�
`Aآ��g�x纈G:G�o/�C���SŞ�te��d�mcn���,�*�.�\G׌$��Ůw�7�0���'\kc����IMa����yu"GV���^w������.�
X0>�����Y(�w��[6��Ź(�,-�r�AH��5O�o�����%5�l�Y�s"妍3���#���I��K���ź02z���lYo�'s\Ws�#/�v9v���[�e���q�
��)'@"�@n];4�=�+~��:ԉ?S"�?`|S�C�1�mN���L���P.p�g,��l���S��+��q�*���������X�PŃ�d�b�����i�w��o���fqS}S�>r�R0�tͰq.n��]?7[=&0�-�ӈ�[�9���=�L�G�G ��5�N5�=�,��0�8SK��������:�C��A��Uw~�`8���ޢcO~�ld�pL��/>r��S���閁����$�zO}ٛG�����Z���+놇Z{VL����0�uxɕ�ha�2�|煆�t��]^6)yX�sq�m�<�T�}�P�{%�`uW����ηp�W���U�R�z;�&f=l��(}hm��
�ri�v�υJgחp��$φ uV��P�x���7ۆNa<�}�p�7Ɡ�,�B_�.ȇxM���-��˸Y�F��F���J�Y�e)iP��-tu�U5��g>������O�}+�p'G�z�m"�f׾�� ��X���gy+���)>�5�J��iR���Pulpvb��,�{�tV/]�l�?RÕ�Yc�-h��D���[�V`.���eq�x�W����ofǲΦ�F+��z�x��%J��eD�ㇲ��2��Bs
ї�i���lFv��q���S�S�������/�y��T�J��*�t�����O����8"�4����{��~�M��y�ЊRI�FwCeۧ�kf,�9c�;ؼ ��{�z(v��W'\wTQ1*]��>m�V���.�����긣\j"ǫL��dn��P�6y�r=�g�AYf���YT��%tS��fB�J��Z~�g*�4�uY`��%9�w7��qB�y�����w�Lo��z=�1��;�Wz*�k�vP��Z;)�!^���7������W�qn�_+�srA�*�[]k��v4��{�v�3�<p6,�ު�]��q)�p6@;s�[�yK�\��j�>ۆ�S�N�kTW��&�Z��.�ӣ�v�W��9�.?:I=�7C[9>��:�T�}�<^�Sj���,��O�Iƴ��j-�c3.>݆N㙏���棢�n�������a�yo�X���m��w9՝0�ʬj�A�K��i%��{gM�D\�1a��0p)L� �L�N�ʮ#��{Eu�0)΅}uq�z=�p��1�l�n��\w&MB����[s�x�ǒ'������ 4��iT�����A�:{�yi�V�<�!�����w&���P�ѳ�6�tJ`7zJ�҈�.7ף����������O��(3X\b`�[o#�����X��gi����kܷ��*��B���|�3/)��W���{>-Y���Ĳ=�{�z�k��{�y\<s桿+�L߃��a��E�h�`���k����[��$q��e��_�\�Do&��WR���˞[ �<3�>��� ��F��ڲ�=켛u�m��룽E�e�~�A}]V5��U_�Ρ���9G��9d�ٙu|��Jg1Y�a`��7��ֈ���"�z2̬ �[G]����s��)5�gJ>R��]M��MܾV��qǚVm�Ե1ȟbM}y�
�^�,�ݫ� �^*��Ձ��$Q��8�K��3s�Og�7�����ci�>�ؼ��,��:p
L���ڍby��~x��״.R&�7�"����wr��B,��m6;�[�{�*�>�Zk�c5C^(�p�N������zjET�7}�:��֗>v�i߹C�x��,�&��Ξa^Ft3���}w�R
����sX�ے�M��oWU{����o��j�����-E_�}�m��sB�d�g��z�g�s��d`�Gv�J���M�����Zc5��=�맵=5��7����x'w���UX�ҎI��?W�À�ғ�����]ۥ��m��]vكnŀ�"����w��*��.H�����;9��v�j5R�ه�?,�`'���:;��wţ�k��~�\R�4�92{r���.0�Fz�]0:�����:��)W���F���V�]����B����4�h�潏r��Ψ{�Tl���xD6�i0p$�y��]KL�M+�L������V�)���G3gJݯ2�ǣb'�V	޺=:��(C�I���쾴�
��+���s���^�'1~��=l�B�6!+�t����'�V������o� ?�p�f�o��Go�m׍Gpc�{�A>=-����W����	}sWo��8r^�g�Q7җ%B���9En�ӽ�I�w�6)#�Pj�s���x|=�w,y�v4�*b�.����\'e��[j��c������$��*�.�,X��*_,^U��n��Bs��1)�g4f-�6����<�̧�]�+lm�O	��]f/-�|)B��}��U�2�/�]T���:��[�4��Lx�|蝱&�	��BļtK��,?�U��W�}E��w���͡�\�E���w\ ;�R�z���r���z$]��;��o	R�yI�.ed,�,!Sx�z�{U{G$E+�Y ���o|xt�[��t�=���
��`Đ�NY;��,�`�Eob��gV2�����e$�k �qBi�+y�N�y<���w�7�~�n�t%��y3�"2CFH���w�U9Zv��m�V��F\ؘu���:�"�FH�I�C9O��Zlo;�`ٶ�-����s��We�A���Y�+GN����q����&wv�׌�]�:|D��ǜ�нJ�Ip�/c�������VP�{c���&�o�m�A�ϔ8W������86�a&Ʈ.����zc��8��<y�|f��-:�&��}y����じ4V	���r.z��*z�����=L���;sԖ���Y+r�y󥍺Is�Y����F+�cN6��T=2���:�_�����Ç����7|Ϭ��}bp:����S�[C�~�Ԍ63lI��#�T��÷���I�iI��v�׊���}{�k�S�v�gk#C���}@��P�Ƹ�U2���9�*[A�맱��6Iz�,	>SV�J�';��:�����z�w+g=2�$E�o�]�����E���_W#
��,����M�I��V�:�g5�k�o�T�~�䍼FW�(�]�TN���Tj��6)9��M>.�|X�x�e�6�.��۔wE֋��,�zz�����h�׻�w���l�]�x	�YW�LS��Ў�7)��=�2��Z�4NK���A�;u�"�.�N�j+gF
���[\HN�{w_SU뾳��~��綁�%��ʔ�JT�5�@r���lWLY���6돥�[�\�^�:���OJOV=���ZA����I��K>�L����$Æ���h��yr��Fƭ-��k�����U~Zt¯��B]K�!����m�#��C�/j��+s�S���MMx�A�Vp5f�OQ�D����!zP�6ԯ�᷋��N9�NS��T��oճl�m.�����Q�y�É�)I��bd�y���l��;b���Wh;B�9S�tҸS>�Ur�`���� ��Y.2/ ꓠ��)��H�\��n�j�f���!����X� 4�z�ғ����Wӎ�A����$n��PбE�[�R��u�5{���X�L=�4��^����'e,�1���`��Q"4�u&���>�]�D"OK���D�O�)�y��ku���/d�6iX%��S��-WP��Ϩ'FIXg.��{�]�~㓤�;��m��k�;�!���c�$�`����7)-geR*�Pj���y��b�0?F-�փM�B^P����7�!����+R�����f���e�����<��l.�Z�Ecr]ĳ@�5�z�)�=bt�nT\7�)'+Wx^�k�|h�X� �:���������{Br��+��R�����-CI�e�o��];��݂,C�W�4�}��7)����4\W��a�u�r<��:����d�ʫ��6��FS���2�D���}�<^�W���g���W"x�>�6��\���8{[}i��ڣ�|S/�U30[�/>���ex˫n*�[��ٷ��H��{h�DVd��m���R#�ݠw�*$�ς�ϳ�̱���RZ*��������<vO��2CJg�Y��Go�٧{+�@f������{ 8:(u���={��+燓V&�^�s����Uý�Ep�ȡx\���`xx@m=�:G��J�I ���i�2��M�*{j�+���ߜ��uC���甁Q�0î��f'�ѿ��v��B�$量S�os��>mz����+��:��V$���·�^��(�����e�+��%�R=i;�>5�U�]L	Ȟ�+F[����.�w��U����C��7t�j��nh�n�(7���cQ�n�$�V�GT�������87j�϶W���L&������0�v��Y�)�Hm�}�v��뜝2c!y�:�)k�5 9�	�&n��K�����Zo��Vx�eoX��eˮ�T�ՊZ\��qy��T�q��wl�����r��}{�A�"��zY�=�i�kp�u��n��W@ͮ�Nҽ5Di�2t(G+3(_RZ���j������j��Z�U\�N�*�Qu�U�힓5��t(M�{T��d4L�XGi<�Nլ��^͵�����~)y�z%��z�)Nv�V!��g���>y�*�Ѻ����7�t��`����4��j�����ĐG�����Nm�`eد�c+��lC(>��f��m���y6�U� ��2�[U�Q�(j	Tʔ]� �F�X�N(2��=�2���c�౑�RH�\�-ռ*���tq�T����a���,���+���	���zh΅�xoKi������=�n`�Cc�[� .V��]>��tU�z�����PS�㽬��ݤ���8H�����y?�Z)q�3�D�I�z)��seZ+�5<{\)�Boe�Z�>ޝ��%�Y��;5�{]r�V���b�|X7 �f�$�����b�c�z�ټas,֨��� 4�+S���oF�E.�TX��3�}/8���mXȗ�ʼ�\���9��ܫ(4���9�n��u��
|:�V�[��jcT�i�b���0ZYy���!1��nϖռ�m�wYo9�z0C���=+N"��$����F��!L%;V�}�bWw�j��wP]$yQ_ڑBm� �͕���Z�R6ƥG.m����	V�35�܄��Q)w�;��qF�F�d�MB��[�m�U���;��+X�KsLZ'�{�4�TP5ơS��/n*�� �,��m#r����+F�]��},�y`�S�1]��w9���V)�f��`f���=�r���M�jb+Z�9�����:�RrW*޳��|�콥�V���ygo�o�i��Z��\<>�'i�|��o���\�֘|C\��sp:���/�D�����G^��Źq���rvaAW"��Po�]�}��]@����'�fr�ڵ�����+�V����ݣpU����z��o/z��#�g���S��,�rr��w�:^�8||�
������c�#�p�U�v�fVs�h�L�Z��\xg:��v�]��U�m�|`r���L�«]Һk;v$6�j�It�Il�ɺمӤ3F��m�8v_
̏g���b�����.���ݦ4��݉�Js�C��*^Y�%�b�&`�Ndy�L�A�[�y�ۇt^�O�[��u��U�Ǜ$�$��� q�z���Ct�HR��о�M� �8�(�*�1�����%Mr�v��;���YIW�|�kv��E�}�c"[$�гl��{���jJ���]���{��vJ�^��bRW�E�ˀ��N��k`*�W+���ޚ��{�z���B�r��*�%�&���\�2%��C!JZ�2$,�
P��!��22C$r�,2���)rq���rC*L����J�2B���,�30��#*������)(C*ɠ��JV���!�%)rL����h���2"��"�	���*(i(�2�h��
����22i��)����
3)+,�p�������!rJ!(2���3!�

JJW%�C'���h0����L���2B$��Ȩ���(��J!���&���2Z�i�� �0�(,�ɤ��2 ������*���L��Φ��1�f��
.uݹl��j�u�h��~��鹣���j�6<+\����[����ꘌ;�R���I�3��S#	��S�����ȣY0�A��w��&r�CmF��Yaؤ�zV/yꔞ�]ǫM�L�W�)�E����a}��6{������2����P�W�'\)��A����Ud5��s�Z���c�AٌV��9uY��9�j���f̯s�b0	�<�X9��N���>����8�
�A�c�
���\��50b�<v|B�"�mMU�@6���K�^��^5�>�L�,���I�Ų�6��]#P�u,f��ũ=U!�0�,�j'd#�XMi-���O�A�Wn�mW���U�T�_��H�A���˿���1�y�֛�⮲�{X��s�^:�]�l��ϥ�۪i0p$�{)WJRg�)�ce27��I쪡��<̺.��9nsѢ"y�d�]�ٔ��]V������:�z�~�? 27e��-g�q`�|>T�6!>�<%��g3�ZQ���gKD�!���R�<��ἁ�Bn�[ܢUӀ����hT�w��t�����M�p����ό҉�Y�og�����?��v����
��\k�kEG��_20[�S�X�v���:e6#�s��bk�/�+�8�f��w����͊Ye�j�m�ժp��1`��8�f��v��$�,����X�����[ԆԹ=��ZW泖H�\̼��()9�,)�-��l�|���_¸b���]�YXxOuk�c�b�8����RO�Vm
�	�����g��C�g��iJז�N��ύ����b���>�/PG��B���C���s�i�J�ٻ?��+�tD��h�.���r��������_">2����)��O%��y��s�_"c	�}�J'nM�K�Z���=J&s|.��fPg��A	g;�_�X�o�ׅϊ�Y>P�������%��a~K:Y"z�b����K��X��=�%��:���#��m��2y��[k�m�z�w�İl�g��:|n��B�� �;ޡaB`.��M���x]�8^b��/1�P�pWS�S��;�Q�.�V@o�Q�Ow8&y1��]�p��o�:�X|��M�ɓk�h��oᎮ#�mx�M�����9����d��5ٝ
j��~��6Lv�\Yv|��84/Z�N���`�)>�D��Ȋ���F�^2h�����ǧܪ#pZ�z�aN���`+
��L�����l6:�aN�k�K��P[�J��V725��+�t�v�hd/r� ����X �
����}l�� U���U�%2"��U��퐖f�T�y"m���~o{����C2�z�5qkr��`I5j���/�o�*�dR��P�ý%)�2�ykkG�O=�{��Û�7�1�k�p�X�S���j{�c�zm^�a��`���	拪���^݉�Y�8����ʆ{~��9]��58�k�R<g�0�8SK����O)�3ڳEh��G���0 ��k�	
�ډ|�.��>Yr�٘Ğt����X��K���;��g��^	���� g���/R��_��W�L���u�3>S�q�2�m��v]D(f烵���T�q���m�Z-,)�e
��(�y-C��ָf�V&I˷�>�Ϝ��������p.�#�J�a�Đ��m��/.�~g	�г��
�o���6�J�x��K�҇�[Uqi߹��G}u.ȇ>	�6.t6���Q���Y1�׼+��!�������}�DR��%}n+<��?#�,�\�6a��A���E8W��w�]Њ�8W'Q�'��Q�� �"6�]�U\n�ȼ�w0���ϖG���˻6]��ׂu�Txl��\.�.��Q�<zf���S��[0K�����޺��V5?c�Gx��[��KN� �y�d鷢��9�e����qk1hR�Q]u��I#�A���ۮA�*�;�C�m�疞�l#Ԅ-���_5�k�O���+zV�f�O���h%ƕ%���;�3�Iv5Z΂={^vEO�u3y~��;g��cMvU&/�Cx����}u�C��?�͊������;7�`���.V+Ϝ2]����=��%vR�N�Zm������7�"!^��Z�;�o.��͘���==P�d#P5�}׎�IL�2�<:��#�yU�J��4j�u"��`{%^�M�B��1��Ş�bu-C�T	P��k��{�!��e0���tB{s4!���T*k���D���Gb�X��5�m�l�T8K~Z=}��2:�9��fCUr�-���B�������TG_�O��螬Sj���,��0'��2��wNo����[�L����qr��џ^��1�n���vTJ�b�����wg+���4O6|���U�Y�9";�f lIQ&+�O�.u3�tSyl9�K���ѣ2�_B+e]�%��w9�ZgL=�*��`�*����O��L�M(Edގ�Ʌ3����b�Ago�@���C���8"���>�l�;�&�I"�#��#�q�>z��CR\R��~���ڿ09��n���Ӭ��FE�u�+��ӅsNZn�����/r 0��\��ª]_c��R�<�Xy��@�v���w�?t~6Н���Ud�)��Mr�5̶�E��
�V�U�L���@>�V_u��Q�']&s2t�-�Ž�ч�4,�#��r��i��Y�������>���'���D��^�~��ɞ�j�X�`�����"`ڋ�����}P����>r�\2KGǯ7�d��Em�r�%u� ��I�$S<2GG��]��<�]g�'3ԩh�b�A�k�*0��S����yZQ�>V=̳��KT��O�`�_f����T�t}���$�#iy����x7&mƜ陎ykf�s�4X�>l���B𿏕����g�FSs����(R��u��޶tOV�}L����zL��r	����5�FOy����=s�W���k�sº�45[���tk�=Kh|{}/;1��ާ.� 7�`�,�&��u���]`�aIUq-�A��w��u���
�-,�
� =�Z�}�P�1��o��j���ß�oRR�0۝ģc(����uV	~+X��]6j��Q2��&�.-��WEb��9;�=R����cئ�K3;������cz�q�:�t���՞�J��,�c*4���f�YK*��?���@��-;Ҙv���d�ZŦ!hX�)`�O�@:��gQ�rwG]�ɻ�OO��=Sy-D�f[����kjm����܎�J����{+M�S�]���f��>m�AE�(�q�j�"�3G�����棱0�ؠ�mrw6��-�}!냩{�n�Ճ�"㡛?uh����xD6�L�'��)WJRg�)�W	��^���;Yw��y��#�mB�~�4r��~ϫ�]�ٔ��%�g|(P�g�4WU�h|�R~r�,Vg��xl����}��3����|$�F��_@�M� o�N��%]�ۗ���9D!�L����o���w|��������]�.2�WZ^+�����؜dq�(�۵䲪��g��Ca�����f{�C�c����9S}����X�+�s[����~�3����*��$��$i-~Z)4�c�ōu�*u|�yJ��|6���q�=ѫں~�蓬�H�<���f`��IC�1OV}R����@b�L��
��k���UcǠ�=�s�ڊ�����[D�
d��D�ɷ�h�f�z�K�������1eL��B"ً�a�Q���������'M�,���X:Y"���,�~>�45Kz�R}���jKp��R�;�2;킭����R���؇�Xto;�g�5��t�,`~ա�������sA����d��p{q��y�5I���I1����p�ڻ��u��B��-�8��Ŋ�d�
�<�wd����}u:d�m����:��&l�^�w�H�bv� ���� K벥Ë
�������b��^�5�O�1�ܭi�m]Oi�owh?}��yBxf�L�g��	[FaFDm�U�0 �N�7nI��.t����c�t��	7,���2��rۃ��ŀ��?S��px�Vts[�U�I�ry������;�u hx��. ����#N��:�\2�4/�DNu"]��,��XѾ}���=d�a�ʤ���:�!���u����:���e?ޫ���~�pr��ʛ7�!�{��ۆ\�8Î�c;8��TjEX�g��bL��gׯ���,.�����#�O�]�Ϫ\KZ�o}��#죂J�⹮`Gh�{0�8'���R�K<��Vřݲ?K�q�a!�R�v"_)�bf}��QϦu��_���z�m��V��#e����*�<P�,��/�aM�I��V����=;%�c�V��.~�a����v�졇֝�$���؁�r�i`�NME9��q2��V�)cn��s9H�/)��}��p���/��I��t�z�1�ԧ]>��i��|L^\1�o�]�'��Z�faj:N�Nx�F�q<*z�j��v�Պ��(��]�!�̏������[�yG6���Wmf:��п�b��ڃ�[Z�ᘬ}��;�P�ػ<��f����	R=d�������M�0fuK8��enY���,\��W2m5�A���$NQgyi�x]h-A{^�3�A����Ӽ�_#�:�UQ��О��R3��Hlͭ��<�=�I�i�7%���R#"�U�὎+8՘�=G�t�}bV0�tq	�1ٱU>zV{�v΃o^z���*��h���E���������aĈ�)I�����yy�d�}��� �p��XSo�+�}P^��u��h�E�M�<z=Vi�1~%�E�X�y��ǈ�:+����,������"�l�tz�
����\��}r��D�V<�^y��|����8���X���P���+z�J�n=E�]��|���������Ψɓ�hr(�r�{}+=i�;��!���c����rdA����#jNP��^��[�~Py�厧K��/]p0��^�gS��RƜ����d�{���#�롳�{��ݣ�'mM;�C|b��*B��4ұ��k�0�:����F���ބÒ��ى�N�Ѝ���\�U�:�������I3)";��|U��=Z[\��8�<��*P2'_6w�*�Nu��kbb�djjZ�/��\͂�'�U�y`�[T�ngV�:]'m���B^J�%�w{4"����2� �YNm������Zx9���@���gNz��ׅ���|��ĝ\�	�R�{�ͅ���"�.�u��{���-��ő �5��sqD\�0qP�$�3��>J�g��Պ���õa�.t�s���η}����*Ώ�<�$Gd�@�%D�&&u̵Ԥ���Ð�%<����]��Nc+ms\\
s�F_��;�m��5ce��|��Y�'��B���gC,,UњT<}=�UW/]���{�{CWC~W2��|�p�a�]=�:�@?L�9)-��=ʹ��̍U�iI�WF��;&=]nv{Uf��Vxg�C�K�&ĕ�笃c��G���L�՟Rg�u��={���mE�{(z������(��9�.��
������ڤhÙu��i.�;.H�}/ "�%�ΗuUd��x�Ea~�n�#ۗg%]t��������+ne��Z��O�&��A�����⨷�;��<W��$q���	^;�7x�U*�݊��hs/kz�������:�-q�RM�5b�6[��ɓe�]�]j�f�i��	:ozLG>׹��;3�+c$>=B1���ˍ\�׫ӧ�����2�Zo�%��U��ɮ*�V�0���ئ�=��/F�׭�g:�ڶ7�_�]0t|j���4=u�Xeb�0�ri ��7�w�V�s+#�et}��a�"]i��A������ȫ6�4��d	=y*�Z_���1r<߹Ц=�>a�W�~�P_�\]��ŧ@�J�K�{E��Mo���rr ѐ*�>���e�Ү��n��d��O���P�}A��Z��}�W��1��K�ZcP���LUL�Y����r�Y��{�[�t}����(�^,���P��Y�H���\�P�8��f�v���s��b��-E��,3n��'䚣�W�b��eF����z��{��ﳳM&��]�&���4=	Ά�S�V���^��L_-Eql�i���b���7m�'o�k��J�����_m�р[��o�"y�Nڣ�'fP"�0m'�{E���^�e��c���w6�pS��>R���?��؄����_ޏ��yX#C�����G�w�{����P�'\ӗw�'t�$[�hK�<�Jg{]\>8$v8���k��=D��8o��Nz�vf�j�CxρzQ4-�\�U26���~�l<\�^�f{�~w,y��fl��"ɦ��]��}��;��qM���z$x���R'�],l>8�/�/!U�'����,�I��q6hq>��ܱͨ�x3�]^�&�}�5� ���ӽ�6��Oe���wJ�xS�T�_;�l͊��eF��zk�,�X����h��؄ߔ�NS��e���uw:�;K�Q�%F#Lf�2�d�Jo%�Pm���F�H����7q�ƺ+�z;��3��T[@����qn�	��³j�Y����SFv�_"�b�����͈<���7���B�b�LP�tÓ��)�4����س���ʑ�:���O]��`6��
�<kY�|鱗�{��`]z}j�)}&\$�9.{5s���ݺ��y�'$�8۱�m���>]���e,�
燖����+ՌAmf;�M^��f���-VƩ_Voj����^IP+�%�э$�F�A�`]۫�۱���z1�����}�֗���He#u�{{Bs���/i^�x(�1i}�L�	c+��M0��X�*�m��`%���u�o{�'��tE+�@��q�O���=�R*h��ݰz�%b
t&)u��)��ue���82Ln��IϞ�|ƣ���3k5��b�nd�iI�5m͎֚En�)�ӝ�����mMi�x5�$���+*f����F��AL=�&\��<u^]u��"�cT8n�L'�G{
��������ֹΎպ :f��}������w{(.���z���h's[�n'�p�J	.�*]w,��ΥԦ�s� Y��eo)��=e:�Խ��6lC��HEV��'+��z�.��,��p��^r��\�楌��S��i��ݍ�bY�����遉[�bhSD������w�]�I�)�*t�iz�Xf��ras3�dO��4�餗[N�u��"�h�jȜ��<yD;-d\s���s�\@�n=j��V�u�\�3lD(L��xKm��(7��{r�r)��vT�ޤ(�fY�s���b��o����Aˁ����Y�D����ۻ� ��ʋC�eNg���g*(��.�Q�N��u���@�H�1��Pٹd�E�܃5t3Kf.�����K�b���1��˭�](�
�x�+f��"T�]6{v#�u����O��(��c��f=m�#����WV�M[�k]]o@т>_G�,��*6�_UɌpr]G��� �H��ڎ�h��h��Z礱G8Y�\c6��"wN�Yz�٨աz�u}K�-�er�L��m�2��̐ .ͰE�++���Ɗ<���Op%���)�Ւm����8Z�/,��a�R�����Ԇ����qq�ݱiN�*IG��[ú�U˩d������b�2[�Mq
@a;|�V�pqѭ��f]�X���O3�z�t���K/��@�_ �z�r�nɗ3sտI�%�c��N-���T��b	"�R]���S+A��n,AH�.s�2�m��WQ^�ިFƜ�^�S�
�sZ붷�מ}�u�����@j���ɣ&�(�L��)()
��)iH���+,�Eȉ�2��'$ʓ$�G$(h�*JJh�)(���V�� 30(L%�L�!
��)��&!�)
P�j��
L3
i�c12i�rr�3��2((2�������*(�����H����1Ȣj�0���¢$Ȥ�S',�'	\"�����h2��Jh��̪�+*2\�++$�B�)(r� �"�()�#*�ɥ�*�2J0�ɧ32)L�h�L���)�i�#' +,�0���,�#'$��L���*�',��(�
h)�"�'0�L��L"����#!�2�
��*���&i
rL���"��²j����3� ��rj�"������eDg �d!�㊹͇�ue�Ae�b&���[��A�ԓc����Tz��5�H����n'}��1����w��.�S>������#�ؒ��^�W�u�O��=|��c��
_B��h�a��C�����ߍ:c��ɘ2R*�{8�u��
d�����x&���	��=XJg|���;�v�c{�J�rZ��9.4\��v)ɚ�qD�緤�s谿%���*{=��zv����H�J�ei};]F7s�u��l�[�MC�V�c�د�����Y�m�[P���ئ:�/[@_��W��a<Κ�s�%�u��ו��85x�5k�n���<B+S50��b<��6`թ_Of����=�x(�
�d���f��矃�r~"}k�Ύ��4�V��6V�҄�oB9�L>��N���6�o;v2�`�X%U��p��r��
��:���o/o�sڢo��n�T��f/�̈]4��/��IX�0�*gƫM��f 1��mٳI<��:`����b϶�%�0������uMz��æm��0�*�(s���fbߪ���{o:�#U�gNCG�FD=�}8�4�Gh������+�����<�pvo���8vꔟ��c�-���]�g
#3�W
Z�VI�ծ1j��S.���]�-��ر���:e�������d��F��&��N2;p���Dh��"hob�/��N���¾a'��a�8��K��ۭ���ԫ:��'M���ڱ.��u!�Wbߒ|��E�'<��:���e�=�����
3o�
�H�\8�Z�˦�0�HEx��ٕg�տu�2��tY�L*{).�G���3�O��<�Ł��mnR<�R�ᒕ/uɬ&��4�����r�{Ƥo�iu�%�>{�=�C-p9�P��P{'�$/:i`�L�������t��Ax�H�K�rʀޭ���!�UE�G1W��΄>��ݑ����m�_u���*+��ݩ�B����h��D�EeNVu{=����Â������VhÞ7����jwp�%X��s���:G�Y�.=��0���C��졃e��,U��2%�ud���s-�,����g� ���9�����E�s�or����5�N'�lŗ��ũ,X+�e���:�B��LP@n��;f�=i��T���P5�ן_��q���n�NӴ.m���&e�K$�^^|d�{'|�;�Y01��K:Ai�~�z�TP=W�D��R��W��wM�ͳ�-�ڽ����,~��74Ç��r���i&��&�����Sz�{�F�]���O�6oc����<�A���wVJ�1� |��<es�(=���ɡ��WR|7r��EkY�W7K ����m��Ik�\�;��gJ�z��)�ú:X�~���I��Ȼ�T�W�or�.��Em��)�h/��0*�D���p7���zٗN�(tuKs��.��.���ǹ��LX�Vh	����Bv}Uֹ8��(Q�Q+����a��}nDB���q^yȬ���ڲ.�K�|�׵��j.ڨo�>��f�#�U>*�螬�Og]��]s$B�Â
�di)=���rõu�^+�&∹T`�~YUL̷v^
�؅����k�/�(/�x_Bu�2�cA�w^��}o�Y�H�M����LR��
���M�ɩۜ|��q[e��b��"���,S�qs��Η��3B�X ���%����e׺�3�ٶ�M���$NeuR���J���;����kU�m���8Iݛ�ʤ����(��w�֚O�Zh�̅������K�����=�e�-
��������o"\ːΫ�g�+U�c�l2�e#�����d���v���+��p��=��d �7����PN�����%=
v7�˦�����V�b�����u�j��YY�j�#�S������2�@�!��7�p䋨��<�PuЪ�[Ƴm%���f�=�nJj'+��y$w��fh�&Qy$y���^��\�_0��ǝ� ˯Wk#��ULD����Rr�����!��<\����DEmyjۃ4#7��*�-ף/OA�$˫=;3���i�jw��������UX=;O��٦��
��l##�m�����y�Ӟ�z5*����:��d��w~[]����O?V��)��܈�nrN�{!���gM]�2UE���u�D�==���j�n��1�w��S�Ss�d�b�xF�ܛh�s����o���w�[���q�+�Z���y���&�+h7�#��Ύ1|s�g.*��l::kLS��S���@�Lu=8+���3g�o<Ӛ�.��P���#�5b�T�ҳ��/-���pﬂ7k/u�M���Rq�;}\����`{��qޒ��2ŀ_nEW)a�)�nj�����Ȭ2�s���~�S��}��u�Z$,p�;#��@D���[�'[V0��р�&���c�A,+{^	kB�Ů�{�����lp��# ��<��ɰ���]LmY�CWo��p�J����ξ���
���_U��#ν3��U�q���hf��wYWD��t`G[�Z�y�E�z��x��x���W�������5�߹:����9�lweG������1j'��N���|*{6_k�W�Y�������{Y�l���U�·Y&?I����j{��ιltY����V�K�\.�eKEͽ^~��rf��v�.6c��<�&oϜ��S�ͬ�uM�����N� �הC�X�wk���cU���}�s�e��{����j��pWnĘ+�9����Mv5�����p==h�.`/Aî9�걚
�s�ݒ�(]�y�o^�%EX��Ȏq��7p"�Ҙ�7�0k�����@{�pS�ڏ�v�f�~%��o'9���a�nի��%����4�o�c;���Jf��Ծ+�[H�>��X*tŇ�Y�xz܀�.z��ˤmV�=��f���vޫ��g�3�Jp�FȺt�*^���C-ؼK����i��p�Nj�3`��dަ	�4�֚�\�ʽ1���ڻ�]�����;LK+�6'��#��wG�c�C�WQ��\�+�P�"�u���H�l%R�YXk�ŷ��t�:V�G��g�G��ڗ^}z��&�����:+ ԑ֟�7�,���Qc���WeP#v�tF�o�S��k%�΂����᳟�nO{붭��峍K�ڇ�*�{��c�r��tg���Ljs�37�?<����'j<�n�{;�͆{l��S����8��o����N<ٚ���૨���#�7>�Y����fv�C���
v��6f��}A&�l��v��=#��rw���E<k�}��J�ߦײ�N-�]�nJ2��q��9�:�=�l�*�%�hA��7ڧv�������Ĳce8�uoyK�-���;Ʉ���&vR)�k��zU.��ύ��_��N��Xj����x[s������>�2+�.SG ��ed��\||o���]wPz���1�Z7����~:����^�n���:�>���F�(����X�!��+���sLwN��.�v�P��PL�Tï�1���,����w^7�f�ѐ6��n�x�Q�J��R�n���nq�R�S�y��Kjr�C6�2�ŵ �9]��s�4u#�oS�,rUu���#��N7��[��ll�[Ï��N��r���n�̈́��XT;��ٚ�H�DMZ�����y�����5;q�e���"z�J�м��]V�(hs����O�s^�o�b�~�4�|�2=̜����Ggo�9/xҡM�X���ij���
�����y��r[�=�kx�V���U5t��:	��n-���m_z��ZT��?��
l�L�zH�2_gVݕ���[�_-q��N5��^�ns�������Rz!��n6N>8�xd�Jȅ5.}TA�;�6r���QVS���N��KCf	�5C�n�vm��0�Y��=3�y,4��k4%��J�	񯳣��{���1���v0#�lݸ<�.8o}8�\�e�\LY}��;��u�z�瞜�K+"���_.��"���G�-3��;s���Y$��3���z��KJ��Zǹ֮���q��S��`�{ݸh�θ��=P�	��u�]X���l�۳�2Y�Kc]eV��+)Y��gu�Y���=iU�H��\�J��;���&�[*�LDj.�,�<�λkKku����[]ۏ��DU�0��U-�����>=m���g�z�
vY}���KsR�d�Shv6i|��6�b��i��u�z9B��Tx���lַ��3��8�Z��2M�;-M  ���R���L�t�S��C!u|v����;�j��
��ԋE�g*�����ϯ���b��\��C���L:�h��@eG�H�/r�q���zU�s��v'à���gjL����?�������ʛ�r�Ӕ��\e^"��Ѿ�q3|¯>bą��3d˩�ϝ�ght(�q�l�h�T<���GV����m�99-�d{�m� �%��q���n��5V珼U��2��O*3p��i���w���LBg���Ww(�>Ƀ �`��MTce��WN^�761`o>R��r$��(����g[�sڧw�ѽ��fo*pޫΡ���ῷ�.v��M9�=Գ]��������\pr���)��S��c������6b_�h��������7���kj�>K]{ V��|�p��d����>�a�s|*�jj<�:aP����_�; @تla�������332l�,J�7]OGx��7�r*������7�B���֘�g)��W����yanjr?;1����+�μ���Sc�M�C{ɲB�Y�#���UN;�q"�+���5�>�ُ���4�͒��=059�7����e�/�cϮ^����2����5�/,t{��.z#R�z��xBs˄>��r�02j��S��V1pm� 8�o:��>}���P��V�9y/��ł�zCS���z�F���\K��:U�u��-�B��[�=;3��J�`K�轡�fO�:ڱ�&�W���i?nB��|w>]��y�ʿ]n�/R�q����z����/�K�bV	e�4�xڝ�S�}��]{7����W�Е���ʱ���}�T�~$��.�|^/�ò�O�E�i�\VՋ^O<gO��˛c7}l%f9W���2��'��NxYo����*u��^W�B��6C�e�Z�� �{�������8h�x�z`3�xSq�3�����9zO@�r��rQH�|7R�Ѿκ�E��w)ZL�/�_�K)�Y,�o�G�ǯ7u��i�5��Q�mNd�.�u��&f�',�&t�+_�"�^��/7n`�g�y�C:A%�>�i�͹��s�u� ZݚV����8O�p�h^n4#v�dhvK���实'[C�_Jz�k����tOdS6��c7�u'�~M����YմW���{����v�K#�oM�����S��N�-8���z�!��`ޚd�}LLk{�Jg����yѫ�6yt�"_�u�W,56F���c|U���[(�(V�l5;޺W����|&F́���o�]7�~�w�j�X����d��m�7љo�A�Y�x���V��>C���=��jHw4U���fr�G����z`�/��.�u���8�[�}���2�v��ۋ�U�;�+=w�}1�vL��Z*v�/�g���{�����Z��{3wl��3�JOgM<���ЛT�n����W��0�]w�����TA_�����PTA_����"�
��W�����"�
��W��* ������Q���+�WTA_TW������ED��* ��QȊ�+��TA_�TA_�1AY&SY��3�}ـpP��3'� bJZ��{mSf�UI(%"��QJ[j�kR�0���i�l)h5��"��
�P��JEUUA@$*fԐ�P��-����UY�f1ljZ�k6�j�6�icd���LBlY-*�b�I�k,�mVZ�t��l�Q���i&�I�k#[L�PV�fZ�ślb[[T^�lj��K�ic,��M��6Քce��k6��6�l��eMj����kjj�+aK[5���d�kl�j�Mi��McL��m���޺�����T�o   �y�ʔm�Wm� ���:P�U�����m
�i�wt�[*�H�.����KmR��]��U ٮ��F�SM���-�5m��m�V��V�fٓw��L�  �B�=[-���QB�eG]���jg�E*����h���jU5U6���]�:Q�WR����� S�F�ׅ
 �B��U�[-J!����a6��^  	��B�C@H�y�z(P ����B�(Q@ ��B� 
(�=]�B�
( (^��B�

7��x�5�1��Ӵʫ8������ �U4�%"IU��5����5�  ��5M
�n�R�f�� Ҏ�)�]�nܮڔ���v%JP�t��Kj�)�ո�h
n��mZv�hF�u8hU��JsP�նʹ���1�f�O   l��26��������i�R�m���m�.�8:6�Tc��
timmcV��k]�Ҁ���������ji�h�wU�kUR�YU�6ڲ���[x  �=�-��&��ҕB�\8���R��V])-ju��Q�CeBVjT��s��5@�ص��
���܂����ͯ@tW{��$
Ū��6��ZK[il�   ��TjZ��͛�m�
�s�N�D��p(��Lh R�0*�	��v�N�̘�'IT*���i��V���+f�YmD��  �= e�e���� tZt�h��+�;wn� 5������S�;a�P
�v�� ;�ج[m�RئTl�*M���   \�U`݇  l����U ��m�h;L.��Pj�tt -t� iMws�@;.a�QJ���m&��[lmmU��&Z<   fx (^�����H
�Ε+j�k[7f*��5��uѶ�kF:nF��M� t][EΜ�Tu#c]s���@o 51�ʒ��@h�0�{FR�   OO�R���z�F� "��	QI &�CFM0i"&ʩ@ ����?����D~�K��]~�q��ɹ�5[��a�`^N��T����{��{�{���$�	&�! ����B���IO�H@�2�HH{�������,�7�  �"�U�����R��Y�<���5��Amp7a	b{1jx�ỵP�4�ڹ�۩R�����yKm�Yu�V�I�ŵ���'�dwBC&�nÐ�>ŷ��d-i��< kw�� �wj��lXA,/$�zf���Z��Т&YVJ$��h��d�p�8��Yǫ����!a�[��y�-{�����W���t�˺�,��+��4�)�s� j�%5�4���y��d2�w��v���T?����^0�G.�iH������*@��(��O��k�:C��'��Jv)����Ǭ���h|��H;qL��H��=ɩ��GbEQB�70'��B�-e����]Ksi�H��;�Mq�J����&��A��.�3�2]ԌC��I��i'X��Tb����̙U���,қID��`%=���4-�oB*m����$�P��%�۩r��a�z�)T7��t֭���N�T�$b�魼���圤�d�B)�����Aк;+0��LRbZ]�������Jə�O1��P9�-�F%h�b����R�ΐ2A=K:X�B���n	�d*K
��R���!�!�Õ{z��$���P8���YEӔK�7K��J8>�` �7Pz/JX�F^n	�Am��7�r���I�1����zU$)ɠK�-a܏o+T��WgS2]�BM*e���M��T�h�,��D�B��0e��Ѳ�fX�R2�4�ձ�Pg75[��^�7��Y�܈\I+	n�W%p�Q��X��hn4��-�5/�MV�蠎��>m�3�%�f���Gu�E�n�hC.�4�:�ʱ���W�Pf����IՉ��u��5<�%��D+q�6��-��uV�@�Y�eE�9Ql��b$L.R �T��� ����)0����.��Ml����$j:Ki1	L�Y��5���'��ov��`��4�MӾ�8_wW`kZ,���эɡ*���XW�n��@�,��"��4�*H*m�L��U#'�z��@�.c�1{i��PR���!���eŗ��p�4�jh�mLڻBH�yB��gU��92�sq���5�xCL�M�rX�B�,
˼�0c�[�Ey[��ۂ��S#�p㬷^'��&��� ��Ѵ�Vڙ݋M����H��?b�Z�ܽz ] ���1Y��pV6�0e�ө��lq6Ѧ��-�a0m��q�5r@�lpyz�'R���\L�	|��V�ZU��Z�$mq�^�y��A
���e��f�)�GJ��aZ�"�z�r�,(�(e��{K^p�R���Ol,������`���T䩰���v䂣�Ѭ����Ƣ%R���������e��W�8(6��Xې�ifJ̹	���"WNͪ�Y�,x�,��F�T�ИH�jv����ʚq����J
A8�u���F��CTd��9V��WW)Ȳ��c�T��B�����0Yů�Y��V�S'&��E���)�[+n�b�'^U;���e-�ɬ,a:��j]����$���V.Y��YHEz��X���Lm�Ta*�x���W�L̳K�]��Ae��Ț�FJU�e㷭��E1 �P��/(�ֆڙypǢ H;f��]��Q�w��)�]�QYx�a���/V#����sUA�f�:�@�K+D"�̭�&�zH�ʓZ��uoPL|+.V�%m�nWr5��X��)�¶%�D����w���}�q��{�9:g@�i�:傀W�2��VPY�(r]��N�\��Q�r�Kv��.�%�̽�h�nÌ��Yw�v�e�[��2����36凲K
���fQKo1�E�i�@�j钨�.ĂSkRI�1S�SQY�f��5��V�Vc��p����6ɡX�a�Kr K�Ai�I2I Nj�Ҏm$��$����h	v��ȴ�q���`]��20�2.�n��"XsF�(wQF/p�� �xq��)A�$6�ǥL��ӥ�=x�]2e��;rE�6���ǁ&�Q��cn!#GF�{�B��b��K�r�J�Kp��eP:���zl�i�G/�.°��Z�Vњ^޵E'�l]<�3U�<���`�<�r[�n�Ӛ3�����V>S�k
��:�߈Mb���*����+6=��.6�O`Y�.��ǆU������s*8�;�H���Y&�͘�=�xq
�n�.� h�33:7��*�F-�m�f�]-��c6��`��+�#AHZI��К�.�U�֕��%T7��n+Z~˫qfl�y3F�"'����1<"�蔭q��:6�;X#�����*��1���V���Q�����a'SfJo6-��Я(gi�U�sh���Ƭ�y�C��;ݶ[wz��B����f^fȖڣ)�9H[�nI��кT����D�ճ
C�݉WT+��R
dщ+o2`�W%0d�ef�Ҍ�R�M*�Q��K��#����� �@f�H�^<�u�x�3���lMܣ(Sr@�?h��2�5�u��!��U�X�XSE={ݡ�kjP���p�X�d+�iݓ����� �8��
����.�;YyYf�E)�h,X��VR�-+�d�ʳ���(��b�*54)Qf� �Y15��{��3.R�p��>r\x�k�,na��"�	QyNk�4��a�C7w\@�@H1ve+�r庹s.<���^1ͥOp�U�*ǉK�m=��D%b�"��	,Ŗ�X�.��i��2���&ہ��ml��ֳwR)� 2ٲ�K�"n�0*�/coJTڦb��
�ױ*0<��ӏ]���Hn�D,b���7���:Uq�Xr�f�\b��ba�n������w���s�t|�>�蓎t��n��0�����������"�g��yOd�R��c��y�c��(��@�#߱=��0m=Ӱ�B���v>[ri�d�xݢq��і�FQ�D���vPrEtj�m�`5�(,2H�p�V��v�]�-�5N�%T�7,(�Ǖ+�G��XV�wu<!�+�g��x/�bzw#���,��V�j%���˰�A�B���4�,��@�܎M�fX����-��(i��1
V�`z��(V�cY��A)㣎�uCv�:��Z�+�l��A���MuoR1�t��۟*6�2n�Dab�\IAu.���n��uyG2PƋܚc���:	��,I���$�_��oj�˦�ۡ��ڽ(����-!�,�t!� ٵh����,�f������Â�n�0��q��]趝�jN7.�	ИjnP��`/t�#���Q����̻+ �4ՙ�����b<��-�
ɹmo�l}���u ����7	t,Dukڛ�@�6��6@P*�Uզkf�v�/):YBiȭfӆҼ�Zw�p�q ��4F2	� 6���^��̬ã��v��;�Ye��e -Veh�%Ʒ����E��	���Чj���l[d%0��%�*n�YBjʮYc��)��K?6m��d�V�9J�-ܫ (�ύ��*�����f�WY5����9[wIE����w
؞�F��WJ�l�F��Z���yTd���E�G���#��=96h����n0��mH]��A�nj����ta�@����+t%�m��VnH4c��y�A*0�Ѳ�� 
�
�Kw6���v5���ʙ�c�^����l��XpYYg wp���1@�^�"M^R%�$�,ߜww���C1�@L���W�ofݔ��Wѵ�E�Ό�V⠄�u�V^ˬ�Ukp��5!���̒]�l�KvG�`��P�F�]L�R�Ƣ�*�ͧ/l��b-���C�(i�-۳j�r�`3݄��p0e�V]��XZT5XT�u�$n��ö����n��r�򈬃2��x��(scP!b��#I�Y��r)2�j�h��̴.�#�,R�Z��*r�n������4VM��rM�Z٥V�M� 8-�Qމ�����<��MЃb�Z1l�u휆�/gٚS�'I`�WB�"�Vj�$k
��A�ר��pՋw{���u�T�)���-��k��z�;��텁:7�n�wIY�)N�*#*��*�ٚ���܍�t�ܚH�L5�6� PJ`�M�� �ؙ�Ћ!L��:.��]%��ʱ�u˚���U(J�Pmެ��N�ڕe���5Q��of�[&���h5,^ l��fk3F�5���Yt��p�
�����J�#U#OC�nTT�R�u�1a`-��X�b��i-��[Tј���W�Q#���S9�m�Y����H�E:��Oc��6��V��T���.!0+�R��(4��2(��R�.��t�l��M�6�iԮBlV�Ʋ��x��Ujpma��"�4�U�FYa��h�3[�yXA�U�MR:�iV�
c��$4�m��麯��W0嶠�S�R���[
�wxb�6Y�iML��ieۏ�i�^9,���S��Tt���*�ތ$i�Dܒ�GAd��6w%����e0]݂�c�$�^�ǚIYt�I	�/ig�Y�ުd��h��؃tԼvB�%ό�Z����QPX!H��1�@�Z!@�@���[Nޣzks�9=��	?A��n����̋KqB�������2���u(�u��ehT�)����X���i؂Ŋ�����	RT@�;W[��Qc��Ɇ�7"���;�aYN�WwH�.�6�(Mf�[�Ѣ��r'"��f��i<�����2%���������L��J`���T�)�K.���z���0S��Gb[�5И�i�h@�*�q�-mn	d	(�YOp��� �ĵ)F���L]VC����X�W"�N���aٖNT,zr��(���X���t>r��n��v��u�g��B���6|��Ÿ�
T.\�X�0����oV5d٦�pJ�yJ�0lbrf�f�n�	�,�,g�!Yz���&ұfa�HQ�2 ���U�2U�Y����`�sI�jPt�r�	���ю� v�b�Tsf��vFů�ܴvFf*�q k,p�f��K$t
6��+m�̫���%h
�0'�t��Y�)���j`D�6�^K��U���tB���Jx��֐�F��
7Q�F&�m+S�U��
6�L:�L�
��fvr��~WsDfd��^(Em'1��:�f���M4������z��@�U޳���=�Ѣ�KJi�)�!���D4I]�$\*ZjT5���Ʃ�̗ BQ7�*�9@*�I�h��m�z�q�F �'Ri����5j�̽�@�r�MQ9���&���`�s5j��݄�ǩZJ����ylYn^]'�
f����6��̃*-��ȭ�K�`���ͫ�`�NY�t�2!H�t&��)��Z�r�n�\w�#`�f��l6��V�7+F�̭�m|�z`*�� ��-i��V�n�)-��K.��!L����2�ko���w$��2�X��
�)�)�(
�J$Dc)ʳ����V6��I�������ei֌�Zc܎�r,�_Gl���i�j�C	��_jյ�{�S;� c�q]�$�(�@��U����� ɵ,ة@Mn��T+d�A��*7��j�,v�ୡ`��.)@�.��������\�e寄�j6/lh�޲��Dk��lFؚj�j%lA��w�
u�Eم-.��-�Pۺ�p�f��Jn�Xi{'n��1���L���[j���#I��)\b�o�(i*�D�\ݶV�$�ݛ�PU��Kw�m�$��L�795mH���:p�N����|8 �4c2d�<�(�8g�Ï4wh���,\��i�"��yz"�aQ�k�	��&ov�g�.�!��Z�h���ƃ�޴�k�{|E���I����Sɢ�q��;U�emn�2��аc�)j�X**��svH�AĀ�&�y"E�����B��7�Jŕ$��r��>����W�����������U/2��ہ��,��i�J��,,Ӹ��_X�ʩ�c.=���gKXeR����ZD�iun
p,{X]ؚD0)k7�6S��wPd�XHӥ!I�~W{��"��!������6#�F��س\���.�GKf@�l���N��rɭ; A�`��Df�o2���F�]ڊ[�&��;���_E��`hO~Żmk�kyGtI'�
��.^��W1LQ ��v��m�5+&Sgjf@�r�@):P��h%Wf�N�V��Z��%���ݦ[m)N�m�	^ǚ��LM���ۆ��l'Z:&<	��S��WYvtl��
�$˸��j\���+t)a;.�%�����ѷ����Ej���F�U%]�`sU��YX�9vȂ��n�F�z�h3@�Q!�h�'1��9q��+/E�V�y[t
�yZ��R0�i��Jգ�i�Z4�"
X�ɵ�Ee�9����oc�pTܫ��B�e�0a�o�^�)+��k�֐V63!�[5u��V���Y�Y$�	q�x\�qnӎ�f��;�cSt��[VN�KZ���˵.isN� �k*��Yh���%�Z;�����U�N���H�͏\��m��CHQD�ۅ?���ɠ��D�ԣ��te-�.�	i��p����L�H���	��S:�}����v��� �G�oi}7î=��3�P;������2�:�$��W����6U��D @���ѯs�X�-� 3{#ZOnyw����֪\7ZM�-)���(��2�U�B	/�c���x�9f��SV:�xV�r��;������*�N�>�i��x�w�j�""s��T=�]��ԥ'g��^�-�{���p�_N~�	+j>.j�"N�\Z�p�P�IY���W�ǈ�8hҞi���A۾�aW�\iu�F]]V;z35f�UQ�/]������>�_?k���.*���y�:�<U�Y�ιu0sW��F���{vb��2r�{4M;:�[Њe��:��X'\���);◣㸰^V3:Y����n����Y�?y��2�-S"e�������B�\��Sb��><:t�
�=�9�,���žk�.ZZ���/�I�t�m	A7&^.$qm��"r;�7�U�����0ٗ��C<i�3^����C}��<��:W`[�w���bALS������>�lR�O�L�}�	��dQ��E�7�iwpnYq9�qEt[m��������*��ݾ�I�X��0��C*�a nő�h��Np���l�)Ǻ6�`�ӛr���eq׼��;����a�k��R�WR7��Tve^���O)��9N��h�k�|�l�r��r�{��a2<��e~X�:������>%�۫@O�i7��>�9O����v�b7�n���\B��Z�.�"�IK��/�bEm�f��۬qCq��^W�M�
����j��҂���)V!W�(l:(\�v�>��|�K*�����=7�S�[5uCe����e���5��-�Հ�D�7��%*�l��(F�貉��h<�����>A����N�2�=BS�p��Fy�Z��{�<���xG�!כ�{l7��Zs�������]�vWn��%�z;-�r������A�B ��h�)���e`6c�MD�g5�^G(U�r�{6�t�����4��;A6&V��0�EY��G�@d��ؕ-��G�{h*gL0ۨ(�w���CHJ�q��($�.�7�z���1�!]c�zE���Ǥ ��$�H��x3aMYw`��Ac�ţ  _8��n��aot�e<�0�u�/&v��+_:A�m��x�9�W���P��իR)S�w��]w�m�:v��'���}n ����@j���p�g����p��e֏x_��Ozk5t���\��{�`'`�ë)ڸ�Y���+�y�p��fX��9r��6��<`3X֎ξ�P���}:{�d/A2��E�{;���7P;]7�]Y)�H��M'Nԏ�=:�e>�v9�@f.���l��^Yzn���O��A��Tt=�l������9
�rEq�Q>�i��+q��f�6���vh8ἡ)o��;&ު�Vb�\� +��'��P�P��ڗ�V��yA�[���X�w��)H���rf�<Rp��:
5ۊո�R����Қ7�
���,aVy�es��%�Ok"����`K5�iQ����V��˩nR����r�:=�O�q�ԟ��gn{1�=Z��-���(/$�[�@��M�-�ɼ�����]�ug���[�vr7���N����o=�gB��WvWV�u`^�n�@
�Ն�O��]8��<sU���7��`���O ��co�2�Ϣr�S-��X�ӗ�%���	9B{7OL�젌齸K'xb�u'��{��f,B=�!
�@�z��9}m`AL�L�)��q�����A7�u�R;5��p��n��H�v�L�\�A�÷/�Gy�0"H�P��Ù	n�q�x��Q2�*��</�~�P���N��X��FY���]�u��̠�$���кoC�pv�i(Y�nbU���^<*�������H��L��T��yU�萔߅��坬{=��1Ј��n�=P����hxŁ#�|�c��5�	cd�ܻ_<(�ː��g��9F9`�����|��%��=]��q�����B�-�:z�wI<IV+��@�Cg�l�p	�~���z��f�DV���X��I���yZ��(|H�te�E!�����X�g�zM�<�KĮ^�qd'�]�d��G�����)��2b6���x�븋]v�A��u��eF9R�fڼKt�C]t,�����,�mK����D���;�=@�&$6�it���n���|�Vm��	��i	L��<�s��ښ�3:���������s��ϐ�gK��G��66�^�L��r�x�`������=�O��a�.�����X� �ÎMђ�U��.��.�(ˊq��#�x���W�!f����ǐ�^������k�n{:�\tRq�«�{�뒀cN�H�*'O���.%����G����Y<p�,�[|h�˲�G�n�:�'��;��rM���dㆵ�(Z�y�He�>���P�<��|Q[uֶ �j��@ݚp>2wF8ۺ
8WEh�mXDoJƮ(�,���א�\6��b{5�u�y8�l]���H�`�ef�Q�;�����v�JJ�r^X�P9mO���ӋOp���C�D���0e䒥��Xψqn���m��!%7w}I�_)t�3c//::c�u�40v/�ʼ�����{�J��{�u����Ţ���$�e�o^��t|;�Aj�敎�����P�U��r��@
,���}����@S���P�:�9�E��p���w����M��V�f�g�LȨ���!�A���F�2����&�F�1h��,��@��ھk���-��,O��PAx�"�q���ej�D�z�u��\V]%蓛ʀ:ܕ�u�&��3����3�q�wb�t��8K~�l��*�!wއ�aRȬK��w��f���,;0��u+���K�";�0��~�M�Ul��"f��I��al�!ӧ>TD��7W���8���uVq�Sn��f�J\�or��)M�����n�/��wE`�&�[8n���7���7$;ۃu��g��)�+w)���b"�;����U����o
��S(B)��d\���]q���ۣ�R`h���J��s|jl�&��՝^'��S�8.̃pH���,�a�{3�c�� 7���b}�Q���F�����B�ф.�U���v�/}�|k��OL�1�n8�a֬�Π(l�9J�@'�|֑��>�o�G�ͮ�PFwx"bẫ�<����J�����``5t��y��M��Z��#�,W��� �3��[k6<�2Q4�|&�<8v[��oCо�t�\�%��gj��*Y�/7���owj�y��;�uc���q�d�"�x��Q\�Lz͝��J�tf=H��5du��ë�Ι���0�W�vJ&�S�#��Nh��ǒ9�H;Lϖ�f��+z���/�,R��<`��_|�<<	�&�]yC�v�|���ξ��ĉ��!�3���y�ysA=����^� �"s�L�YV�M���}�2����r/J=j�Jw{/�o}h��Z�B[<
��FaS�'U�؎*��vv\���#�Y�~��2M��ǂw�[�f�L�pPq=M,̊���u7�|8Y�79_6\"�j�.�Y�'tP����e�ك:���i:_t���`Q��CY��0R�L�6�����z`=[�T*!�3:qv�e�*��S��YA���r��r*=|�s�V�D>���]wb;�<���S�@�C���3���%�s(�t���ᑳed�[�RC�llHJ4����e]�QsTrEC�R��xdK�z�j%֊��'�۝����
o����^!��
���z X�;ͦ��^�_E����Q��&jtI�Wd���5�RF��^j���`�>"�� ��6�Z��*2�va�,�JP��+���ӎ�ݣ�)��E%�S7H=�>2i�V�t���lb �u�6��2�	X���Q6:_D񖪝�jq��0��f�p�-�87I�lP�)(np.f���f��g}l��݂n�eX�!f>���:�V+r9Z5�;0`5rQzޓ�;4�&Q��,����P��c�����1��� Bp�v��1�v��3������I��Qm�}��OJH|��hlA�tb��ëU�^i�:������o!�CY�qA�4H��ܥ�&-�Y�+F��xyq~��r�G���e��1T�n��+9=�v�뎮DC��i�X�;���d�N��W������]\jټ�Y���0`��m�*�:	Y�a2�����Z7��C�5���[&�"74��C��<C}�]�S��b�8�w���v��X�i�ĩՁ{%���8�i*0][�,����3��4od<��s*��5��*��h��s������ͽ���Wn�6�6�������B�1�U�����p�5d����o3�X��*�v�t�/��\�h]M��'٣��Z܂�G<Ok�ڪ�:݇ǋ�Z7|��*X�=@��}�(Gz�Ms'8�&u��&L{w�z�xT�%/p�Oq���ڈ9|��Ĥ��xEoaj�K�%vJb��9Z�S�K)���b�#���3t�u�����Mhҹi�<�l�U���֔�L�1�v��*�j���۲1E��&��D�ˍG*n�e���>�/�lrb�3u�[��e�{��2��u�%1��Zhh%�95V���WGO	_>�	A���v���0*���fC]}>黈�Wu�H��A����$Y��<��%�H;v�:!�>�r���ɶ�@�s��2\����9�P�:�.h�w�u8Ö�n%5;M�[�L��W��ߣ��62��xaɎў�Q\;��łhq�t�j�r�Yd�
�3�֞Nm�����Л�y h��;�2D�����aqڥ�ݮ�&�y[���v�;XbW^�@�2��,��/���)��x���tb�N��xz	��Yݑ\�����[[�n�H����e�7�i*+*���#�b��O�)ؘ���U�7R���vLhֱ��-��=�
{�~��/��A޴�_���š[�M���������9�����d[9�^���zw}
�;�س���7��[�82:J����C���o��W��'ڃ�d�C^�ѝےq��X�l��!��z���p`�<Y�@�� tv���v[v\z3WK�0�a�8�KV�]ԏ6�KZ�\�rBҵX����cB�ah�"��u��g��Q�l���
�|d�7O(���a�*���'�ʗ����J=S�[�-�&�����	F�<�=&Բjn�^�l�	��h��IUȷ8�� /VT�������2��r��ȭ�����+a���Y�~s���/�Q��u�%����M=.x�ps��P��N�+��O4"�����}�/*�8OH���<��M��\�"���ipB�n�t<*�B9�:�N�f�v�5�F����wJcB	��N9d� >�G3k��_r��,nJ�_;mm��'d�5� �Q��g]��Z�ݑ�Lҝ�Pwjؓ�<������_��|�;֜�5r���k��wIy�\YB����&f�&$�a��v�Dݴ��}����#@�#�����Ƕ�u��Q��[('�uu�O��T�7o:�޾���n�/A��0�Ӈ��I'dwW��ҏ�ۻ6��n]�|�;��vLG���^�C���\\���(�G�V���gjal�3� ��-'�{:U����ܔN� w��eՠM7b�f�[��3� AtAh��x���O�dj��ef^���Nb$�a�"�ܲz��QZ"�G7�f�\,��a3NW /.��C�e��;�a\���-�,R��3���i�π�(��=��Q쯩�� �Z&Y�B/[���o,
����zlgpz�!V>���U�_�,�GN*E�]�apab�"*n �Ҵ2����k�026�p7���bs�%G��*�/�ǥ_9����%˞a�@��{۔TT_6K��K�bG�m��G�'(�@Y�X�B�k��ޱ2�N�S�7Gl�E�N6:#DMu	ޝ>`�ynyG�\�F�m) ��-:6wW�{�Ɇ���%��W
͜�m��u�^Y��k�L�׺J���PGg�m�X:��۩��ܾ�e��O��%�凄���U��P��aV�	Ü�-�F�nb�z�ܤ8'W0�1��j����n�� ���gDa��)��6��]����3d��5{x ,�@�����3n����K͚f7d�]̮�Y��%	�{1�ԗ���An;SU�y��ԉ�����G���4�\M�wƺ�=ӹ��U�w]�w�w�7Y�u��e�;ӊՊ��9���j1��Q��������23+��W51���S�T����7&��S���r_F���"L`e�{�����~�Չ@�L �t{6�P��{n��Cm�<|Š ]<70�%-݈�̜���)�y�*��ŋ�sz+Θ?GZq�Z�Av�=�(в��)��F���*��ol2���\Z#5ȶ{�v�;����z�zn%n���Y��<�\F�ozv^��|�-.hޫ�Irٚ���[P_.��w���OIkv���S\P4F���k5�pB�b�WZ�*�%���r���ɼ� �:�.�".�=�z�B�>:���$`��o���%����J�Ú`���;r�GL��8��k��)��Τ�3bv3�2T�/RX����C�Xyü��6��j�Oh*��u���hw-ӎ�Y:��N�C}sRYLǺ�q�	r��x�>�HY�����3Ghn_>,�g��W����~�]��=�3�;rz[�ޛ2�o���ܷ]��i�}]w��z�ө��V�KǨ�(�z�E�m�S���Aػ�0���E9��5_}_!!�@�$���s�3��ןl�|����uha���YL�½�8�F�QQNR����@m+����0���6Ut]��ePh�t��]]u���h�C��Y�\N��_qi{���t�fN����M�\�A,M�`Klf�9���׉�c��;��.k�p��"�����5�s�3o���s�sx��<�\i�(�iLư�ظ_�`FJ�޾�/�垹�������}�u�z���vR�ҞV��cM���r 8���=���|e��MZ;��o,������Ac)'�2]�olkV�)�
�-���% r����ul��5�� Gp�|~;VuP�l�W�Xv�R�����}��.���L񹄃-��%l�4.�X/q���HE��<�/I���2F�����`c|7i�ǂ�Ż42J�^}�}M�˥�������R�f�c�ur��W9�E�5�(n�7Lz|4�t��qi�o$:���n(��\5+�D�]*�ɼ�,�BN��CAL쵵k����)��ȄT1���������맴���Z��pE����L�7$�L��/��s$݌�K5��z���}�&^��c:��#�(A�g���8o�93#���A�v�'X���e�yy�*!yG�x\�/��LՅa�+�.ۘ��V�J��;�s�SY)N}�#��&���,Y���.��W˴.�7i�/zp°�����d��O����>�ݢ�̥X�N�r�)1᡽��G,��T�x�W�d�@�PHᜃ�����M!�����A��P�mG��-���]h{�¬�� �M'��=�X#=���jZs=�V����4����(I��g��c�3�<��g�b0�ޔ���$�J�(�˦�b��(!���uk�R�V��ƴ��V�����̾":�oE>آ�E��Մ�=���=��9F��(vX�R�"�/j��Zkp�N7W̉$�#���k!�3���R�AϺ,q�q��&>��x���[��ٷ�}�X>{�����;i�W`-�J�ӝ��:��c��N6��[W�~��ח]S�&�r�]G���3�i���_$&��>�ao�ŭ=zn伴�xep��יJI�s��xJ��eJ�9^A�ix�㶞V�IЁg/^�k�;6�	���{)��"d�=+�i�^��k���a�X��P�V��PHS�l)y����3�.�<��\�ۈ��*�q��Ĵ/4�;�7�+�cLh � ���;��f����͕��s��6�>�ټ�bH��]=��QB�1��ö�������#t-��r)�E�gb���h��!�{r��P�&jś��k���c�s�NR�ͧ�M�gH��f�FW61�7�'%Ė�T�MF����:��\�0	�T��W�J�5{Z7׏�)���w�	��Q@R���se$,�`�n�K���JG��fE�.f�X^B9$��+ e 	.�u�����ݡ7�#���k�E���>��O��2n9���:�<��qP����i^��f��M{�#-�7�u�W%��N�,�a�ն��C���Ŝ��5rjl��p(�1���p�-%�*ŬU���AXs�"L����� �vE�>�^���� �2��	���OR�7�N-�xS�|�#��(GD�L�0�:m�g+O�:��B^������3V���Sq5�HA�Rs��&!-;��7��>��!�"I����rWl��U��ZH�l������
�`�A��&F��a�o7;��@�u��sp�r�]�N?C�F1�
�7����.U���G�G&ѵ�v��i�l�(!�8n��~C��{���=��9o�ʥяm�$��=8�xtN'gS��-Wt}",d
���������9��"�Wf�v�.��Ț�����2H<�]jKr;�F8M9ه/Y�Ris]±A�E0Y��H�I�C�VF�{���A�7hP{��mu�]��7�(������CX�*��s���4��p���&@�>>��óI��	G���\���d1xW�˳��]
{�(���IX�S�a��#Be����l:|(�T%jQt��8�qH��m�F#Dq�j��r�e��r!��Q�=���]�Be�2�9��.y{����^�%rQfh�*GY�9WyC�SkNfq�c4^�ӗ�2g+�C��������=�D軣ڔ�+S��IV�������� �ŝ7��etjy�>c��,_WҶh2�yN!ۊ�!�=�:܀��4oh�X]*2.0&����T�bH�,8�����k'�ڤ��<&��ܳz]++�#�����ª<��:�y�G[�#�6�����_W��.��t�a�|;wx&gۥwc�:Ǹ�Y��;�o1���f��`-���M<-� �SpVл�T)U6�a��V�/s��J�	h��FhA㇡��9H�^&��%&���;��VR�8��/�g.�n���+���\��^l7V�BHR��׵�9�)^�;z�������y/R�Fq�[�i� P��W������(�9M��X��v������^��:�S�<��� K��� ֔��4�8V3�r�&��5R�a�nP�$�3[�r�x�9�r�Чo�=��ӃO[PF�r��i�J�3.%v�	�j]t����������\�k���}D�L�xѳ=ޯH��Vhh��;�����wY�܂t��q7ۑ�Z��xnm�x�nv�<]�iAF�eJ�&2��7[���Qeq�\�෥;4]�W �C�tz�N��w�#�tVej�aG�wZF�!�X�:K��
��\��}���x�\���O��{�YM�th�S�
���0�w<|�93�}������$W�Y���R;�`$��n���>#<d��q�P!�x&������+.�`	˗$�a��Mh�UfU���X�2i��:�e,�q�@l_\���wC���J�� ����C�l������Q�pt�'px���w��Q�rC��\��F��p��+�Z�����}����;1�ȍ��h�؁�ۻ2��k�U/��;�y�
� w-�B}�R��	_xc��Xe-E7�3�J0-�:"Ҹ�J:=(.�|I�&�'����͊	����]�TD��à�j=�[Qv���H�Mtݹ�����w��Mss�w_� ��I�>��3���Ѭ��.��D�,�O���r7'Շ3_����B�^K=R���S�Kj�R��6�2f�DZ8wF��l���u�%�F�>1�v�9K���b�k~��%Qc�B ���2�o>�c#��]�W�v`!�4��좥k&Q�Y�2�z_*|�3�N#�Hv���{%�0ʗAK��٦Ώ3�<�����}-p���7t�[�p�|�ҕ��&�I����ӑ���M�\c�]�б+�hd��)�]��4h�{-��㢵�ɵ�+���U�������Z���*&%0�w]py��7c@f�b�v�bB�έ#�z���ֶ4`��q}���70�%ǩ�き���x%*<?9vMw�6�Zj�Z���j�Xۢ�쮂���Ɗ����N��&ĺ���g�Y�YL�]����Y8�F��&��LOk~��V#�{9�q1�4��C+\?-���,ꗋ�"�r����>6�Z�����]���H`��侕%���M�f\����XR�O|tF\w��>ZZ(��7-�m����V�ّ���ҏZ*���Qy�f��Ћ���=�q�P�%~-�7�iKI�F�Be���)�{�Vr�pNr�t����R�3�Ux�T�phb;��Y)�"�k!f�7�q��jU��s��k��v�;�n���8��DJCË�x|m8�[��g3pw�@һ,����p�S��f-�Ὓ�!�{rd�.:A�ۃ҄���7kb-e�c��Bp�J֍D�r�;�L@��%;�k川jY|�Ұ~���/5���$V�ʘ�]�`㧛�.nh�w6r��$q.r�I}y�#t���-*��a��E��s�KLe7����v� �B5��E"kM�ےa��2���G^R�ew^ӭrZ#���ei˽NJb�J��u���U����]DM질$1}u������g�v���OsCf��z����=3w�C\�gG�9���Ʃ#O��3j��(��`�kf�tS2�9�[έ�$��om�=���>8�Şk;:��i��X���j�M�vf��GH�X�j�
��
�q���#���l�
͛س�����v\�h�Wz�����0'*S�ܮ,ԨJF���������qχaWG����VCҝu;��tC��w�K0(�^8��g�Ȭ��è+`�e3����^Mz�J�J�:_}�k]X��_��Yf���Z��F�}DN8���;=|*#����(;�5k] ����2�#!�f%�ָݫ
��$�+�_��do�V�L�G���Z��6�j�Ũ�)-�T���7w�XY�a�g�s�,f�-�O����ҷ������i��yus�9/M� ��v�]�0���8Z����T�F�C(�x�.�[�x�l�VaZ���y�BM����|'#�ϝN���I�����w^�/�2t��(��d�r�i�l��6�C���Nu�Y���5ǖ�66�� M���ʷ= ZQޖk��u�0]�l�e�A�
#v�!DnX��{m'��1�
�i�Z�w��Xܵ�ݦ��+B�%��YC\ৈS�tm��S~tz뇎mg�۝"�q��{@�=E�����#{b�ޛ�Ҟ�jSZ]�o��1�[idӗ�:ɼI�-�1�6��Ѓ�-��_l�Z�i���Lr|�Z�����	�ҳ�:��f4�o4캱�<��,��k=S�����Vu
q]��'i�.����
�&'��ճ�J����ATGsX)�u�j�{@=y��֜�n���-���Ȫ�ī�A^�Y�=9��p��Y���)��9Ӷ��6t�����r�,�KU�
����{4��o;���qbU�0e��x���~6vw��RY�{��˫Y�2d��8�kja�l�J	��\+�jvm���um�c{�
��iΝN#���w}H#}���%�Q��]lW�.���L_oi��@��tbܭ%`���)����.��#,�۞;���۸�H~p�F9������+�7��%D���d�eCL[m���f�%W�|�ɞ�]y.f��X����&�ܫ`*��� 
�iP9�\�}�m^�7w�P�\��K�C	� m#8_7����L��a!���I�o 0f�(�DR��f�XsS��#��9��!�y\)ކ������2��%KON�O�u��s��S
�V���v���Q����t\�6�&���8i�]��/m�O-B�X|q��o���Dz\ޭ)��<6}'��x�����K�-�c���r*ܲ��=5�9�^ r�g|����f,�x�]쾔����o��g��n�^ц��b��E}�:!��C/�^"b�%bѽ�m�}�v��w��N
ں�V(z���>�lި7�j��5�u�x�傯l�x�d�{��Ӯ��s��,<[�&�Rq��Tq�ӲV;,��n�I���	5=��T�z::���y��u��7 e+ڃ��zh	P���BR}	VE[kp�B�Մ;��Xzgr
�j�z:���=sQ*Y�����fD8>B��ԏHY"�.���s+{��1��H Gi��(��;:���e,�)Q��K\+y���(�ph�-Sq�u-����0�vc�)���#�N]��Y�����n2�_�����K��1ϭp�+Yb����*lX�d��FΨB,X�� �ڌ�?���.@e�u�Z6�U&�_C�σmћڦ�7p�h��`���8�4�2���;��3��q{u.�_���*ϯy���|w�$R/R`��|�m�	�Β�n��%��]v����f�0�����um��k�tVya��w�`�p�uzP%�6�_�}#������G���S1d*gN˨5�J�b��MwF�a���l�Y]��T�G�9��۳���ǥ���!b'����9G4��y��XB��͕�. ۗ�m���x_wi57��:�O��I�
�}T��x��La�}�}�,��_M����x�LW�;���|p��^�ee>��x��wc�+L���mۉ>ڮ�z6'����:��>�HL�k�^�<n�k�HJG����y̸9)ŗ��kqq�z/`�4�!��՘[����2(�����'u�wn�Ā�D�z�G:𭮎��-�2x�h�A�{�'�T,tzzA*�@��I�r�phAK�.�8���42J�ib�v�Q�=��]'C��r�F����}��;w�i�d9gF�`>��D�-{�9��U��bS�S�T�	�6�'ip�n�����L�z�oگ��2�23�/���Cʇ��6���H�Ђ����lݡj�������8[���&F{��5(4��8���)y��c)�t׀�6/GML曂ȯ�E��{�H<yw��������FY�Y�eEF������d�_<j+W�-��zy�u��w�oH��|u=n�N�s0L����#�X}�|�0�>
X�f�U��#[MY�l-�i����D���(Q�p*Z6evv���(8��DpP�CԴ퇽*�^��&�L��GAs������1�<���=�w���8�nU�_�Ȑ�h"�&�昼�\ݐ��	ߎ����a�@��m�5=�Ϣ�8�Uض2��k��8�
���̷l�"������P�C��	�^�#\�k��q{�A���4��<�P�č�dfj�P��M�U�T�h:Z��d���tKD�����o��v��G�т������/��r�	 ��:���'�u��Y�Y|$w�f��x��P�+��	}՟�w:ϊ�'�VP�\M��̥��)]�v���]�@��H����9�C���P�wrO���=���������N��Yp]��ޡ��r��Z��Z�o�Q�`�<��|�]M�;Yȍ[ܓBF�vf2ڋ��0�+�kU�H�4�H��9�cG7�h;��qI*��e8l���p����p�[�C��<�fu�wU&�;���|�����|�Q3��T��t���

�D*�
u��D��_������n�Fx�-�=m�^w��U.��|�J$��I�At��9;�[ "�^*9�a�HS٦C��r\{3Q��l�巵pR�nt,6�$J��� �v��F�<�U�KT\adi�BS��"�w�:TXo/vK�3�mh�h�J8^��y4L���ܻ�˓ bFe�K2>4'(V�\�9�GC�6[�R�tG���7�ݽ�:�rV�n�WӠ�H Pƀ�QV(�Zұb-��V(�UP���YZ���,���"�����X"#�T�j�1Eƈ�R�Q��J�RP�rЭEZ������6Ѵ�"
�V6UH��Tb"�aEE��a+"�"��(���F�r�Y��.%T�@��[ej��EQQ�QUe��UQE��1@�*9q�b�KaU��
*�TTEADeB�""�`���"�kE[IA�V,1����[J�R,c�1U��Ak�Eb(ȱ`�E����b��FT��EQQc1��QT��m�UAX�(��"�Ȣ��FڤKiE��2��V"��PQU(�TV���
�i�Da[Ub(Ȋ�0TTAAU`�AX�Z �RcUU��D0UAH�)QQb�UUEb"����**KĦ�j���o�R߾��n�8K8�v��~���K0p|\�3��x�&��a��@]y3��}��v���G~���+nv���@B�*�F���u}�Gaeչv#�ϴ��v*#�_��:\�2ә���m��+<���>����>����8�)�����e�|�3s��5v���ݏc4��*�;�P$An���N���T��T���r�r����{�rdЖ�1��1v�Y8������F�U�5ˁ��Z<H�<z�T��G]���t���:=׼��� Q�(lW1��H���9���R��BRv�w��s����E+�ls����;2�1zn<p*��L����)�#�M�!���|�㣊�H�6�xZ��tV�=H�C�样|� ��:S�����S"\��5Ϫ2]�>�o��0�i.\�#�'LL�ah!��llc��F]��x�66�F��q�	T���6^�S��{r�G��z[<�����4��}�VKC��S�Z6)��U�Rs�ě�͠�eI-�H,�]����gT�#q�]!\�Nl��-#��T�,�	H�5���vq����A�)17����<��w��*�������yݹ��%�c�u���� uI�;r�$�C�h�r�$�b�h���C���f��ta�qu۪p:o��Њ'���gb�zW �<x��ݨ�l��v��v
���FPiΆu]{����׸�y�i��d�pxv'����ы�L�+����5���)��t��T�Єtu]���w�Cr���خO��^vb�`���H�x����e���}
TpM������*zE)z��;q��jxU�'���{ѓ�ȖV�s�&��)�+M�3��e�Qp��j��ʈ���PGX ������x�.�#rG[�2Bp���zg!�������_��l*�=��]�j���ybYc�tn��?b=�M˃R�������؇$R�E�T�B�̽�t0�1�~�z��m�	r{�>?M�<'��;�T}��l�]܅a��OJcu�a6���>�w|w�OX*¹�=띀U���v)����NT�'&(TH!��s)]P�عH�j����ϏN���\*�"ƍ� ���:��]��J�*�k/��{�-��I�=��]P%��F�¹����2��	��TAsi�P!�A��R�������b��r�f�P8&NJ��\.ͩ9[�Ȋ��}���CB�����A�;pf 2�M���av���S/����1�U˙(��\<���	��	bn�a��wl+��7 [����oW�7$�7�]�c�*j&Z��»njՑ��<QYR@lW����r|*NHV*�2����T�)ܻB"�����%��;�{��ӳ�H	�[P��d4_������J�<m���9�)�ɜ호L>��e��q�=�F80�Oh�l�fO�QWR}^�D7��=E��`�T���RŤy&��tw(��]]���9EC^ˠ��v����[�"b�h�(>cN�=5!�mDfS���Jݻ���ԫ�yUGE1h��@Ì�/eD;
�Ǌo���񩆓��oϸ�bNՋ���M\���5S;8e0ly$tn������*P��g^���mk���b�~P�Ո�w<e�>��K��G]��{7R*-�=�d���8W��ϵ�Z�,!K�/�vnr�잜�F�a�Μu]�P-��@�� �J�h��z�Z=�\���%�i\�\n�G@Pފ�cEBL���L�FR�3�-����DU��OJ�ӛ��ֱ��w�Y<m�;fK�A�t	�µ�d�_o����-NL�K���ы�"� ��E����������ĵ�O*�gw�$C��t�:� �_�
��6xG��}�k3-�$�4����ܚ�	W7��rB�r����I8���}W�w*ܷq�Y�N�=�9e'���{�U�͸Z%0�Y���s�-9e��b���֟Rj�c��9������Q�veGc�7�TJqN&��M0z֫�����w�BǾ��фU{�K�t�(Ѷ�9�s�7Ur�������55�a7g'�cƷ-lP~z�v��:�2�F��N������x�2\>�EK����B�����g�lf�<�0E�w4#|S3(W@�37�P�c�T�{�|>��5 .�7��S��9i���\�|\]���l ZgM�)ğR�ة;9�S5��ۼ����4�E^�/�p[4�VE��p*������$p�����@���	T���S/��3�������2�Z�����V%9��7B�>���[�J����"�q�������6��}2L1N�e`5��f;0��9A��,bG���R��a��,9�Fh��6s�S|���Vc����ѫ�y��6��z�]\ 瓮�˲�N�
�{S�s�3�y^�)ޡ��V��]n�fkյ�k>��[=�����!�b~{��:A�L�څ��j��5m.�J�]�{t��Ɗ�F�����=N�ߎc&=�N����Z$w��||�lU��zk{���L[��K�h���k3�L�8o�+۵�X6x`���;/��j�j�Y�W�������{]"��p9"<܏�'~~��b�r���h�R6:g��W���FA���:�����R:�Jox��a�OrP�c�o*�l�N�9��9�[S�k�\�R8�Lt��б�:e{*C��	J���!���������V��NÅa����dN�*%خ���ݽ��fWc�[p��}D����q�:(�(�9�jU��ӊ����nm�9��ɭ�-j�ѹ��֮�M�D���U�ʏW:Q�u����=�?�77����t���[�<���fs��_�<�WX\]��ʫh��:J�G�.������U�#c\�`��\�/&[��k�fJ�o{p<@�-R�"n��P`�iij�Ԕ<���i�[y3�����W�B�̖�8*��C4��;3(Գ�c�p4��D���&����>�9D���Rx>���wt 5}����P�\X�N�gDU��p+�#���O;��b'tt�����"�G?�5�L�7������&[�'s���!�؂�X�*;T\�Ѝ��E�U�^Ĺy-�Q	�5��<�_�Ҏ�Yua3z��`���p���t__qf-���o�h""��GS�v1��-<-b���Jh�Pb���v����]�ҨwG)��V�w�u�΅��Pw�r����]_v�h��+#Y"��_��Z �ӑ�3�䦁����XrNvMv���o �tӞ�T�J�d@�`�~�7��Rs�/��9�'�]g+	�KUޫ�����|g9��|�B���׽*�ch|�{)�$X��J�x)��M��tye
H]�P�l\f#�6z�$ߞ�٨-U��GG���*p��K�z�
�^l_k��珏t�>5�%G��	w���+���h�j�%z����l�s��׳�hݥ4]�ΡZ��N@�.hi�GA�*�.��a�܃�Y�61�z)`�?_�����:��3�zV#'���߱;)Q�6*z.}�@�ʅT���`'n<\�N)�W�#�iP}x�m]�ii�K��0C���T+�UME��a6�A!9V6�OB��s��#��PZ{��[=����c�^@�#�B�4:d���(O3���
���Catnq]�.C�o��U��[_g�K8W-��c���Ӌ�
@հ("���؇'ޥ^�7V��F%���Z.���l4s��f��Nu$�i�e���oEB�e�Vb�=�IڡMA� ��kݹ���F�^	��1���1��S�t��?lg.x4� ���F��O���8c�<^pch�)ct|��k`4&�G&�}���`�F"f4�}�I����Q`�l&Y�rgfT8�5*4%y�q$mx*
�l�%K��{���eD��I�X�D]¥"�S��_C�L�O�͓�6!91@�TH��L�u6�{����`G��Q�y=)�!F�N9�#�lRyn0K'5�S|�Pr��d�w��% k�
*�VM5Pu��:TT�\X�<UX�S̈́�(s��x�v���[y���X ��]{��~�/�3��f�RPXt=��o7��Y�=1Cʷ���\���,��Dؖʘ���!������hA�}��P��B
����߼�u��bح�ϺHa�G9�>�p�*����{��'�G�D���Qh�)�����R3ϸj��tn�NjԽ����Nv0EBYt1c��*CYF-�1D4~�L���K�!���`��y�7S�{X�u�2�v�Q{*!ڻq�*�g\��Xr+��J���eJImND��>>|(ԑ[[r��*�H�6�>�Aʱ�z-H��gk�L�s=[�w�'#��u�pL��Q��9^��2��]@�C�[,#	�ݦ�ΏY;� sU�-r�4Y2��95��=vu���;��\����S��~�����H�V�l�4j�+w�����W�K�<�)p9r�oH�sŚȐ�Rs���{�0��W��u�h��z��*��'�Їe��Υ���_w�A��n�#�r�ѣ�ْ�V����(T�yi>·�,��BP"�;�d�M�=�'?o��Y%:z�"����pb��ƭB��[/=3J��D��U{�;D@$���L�<��f���������띂�b����C�]�<革y3X�B"8���/�Wb�����,H�rz&�|S�c-�fNKx���u�*1�]Ob�bTe���p�gSpO ���X�wW׏�ﶳ=�%c�aE�m�s��n/�P�6�u��ӧ%��l��/z�z��7�~(�"�~�	��U1�9J<}eA�8�����u	���R�w���o:�d�b�o��#j�M�S3}H�%a"׮TL��%\-�mW]	�b�fSw�|b��s��qvR�[ 4��N�)ğ
@����1��e��{�:�M`�(n�W:)���R��a6��0�B���.Q^�h	S��h���G]YJ��XJ(]����������j;�~*��X�^x��82���Neq QA�\�V,�4+�q����t�JF�<���U�u"�7�q�P	�i[-��H&���[�=�S�f��0yu�����j�ײ��gkGK�}r�]�IMpZ�5��}���ͳ�o��]���\)][-��i�C�󧧄T7�U�b
Jm��h�z���fE<#,Y���#Nc��xY�d�"�K��=J�����M�Y��ڌi7��%��(i�Dlc�]RjFAVNC9��Ō(�����A�^f�gv52z�S��]�U�v��N�轚��̐��5Ϫgb�:鿐O�z-�kد�VR�}Ԃ����v�c�+�ذ�+�Z9�q�4��~���Շ�Fx�z��O�}���T�^Y��{6tByN!��l�N�puC�v0rG�V�D�6�! N�X��Ne]�\������h�9���[�r�^�)���!�u\'y*�roN���v"�����S�a����5[�L�0e�Qnz
��PN+s#��-�[�w�[6 ��Ǽ����Q{�
2���߯#�Y������D3T�ǝ(�����������N���Xy�{���ڶ{����}sLO��)|���s�J��Gτ��k�t�'w��&�4n���̙��;9d̔7���pă�L������h�=+9���<��W�����WeV�0R�������heT�ڶ�u�Y�n�����YQ^D��I�������X	��C��i��Rz��:�;�mf�N^v=|7�8'[[���Υ�M�/
�o��]@��T�H��3����5ZZ�u4#��j�c2>}�̤6��Jodl`R��/�kf�H�|,|�r�i�x=�$4ߎbܫ�m�U��b��mx�]ӑ%N��߹_��ܸ�d��i�V��dA�H�@�"6��I�	N�C��C�jоdQ�78gT�o<�������i0R���y��9��4�b�"�W�8A�V3릠�~~9��9O7¶��u�ݔ<���ʸd����AT;�cf�Tz��V8�)9ؕ~���]EyPN2=��˼֖Ѩ1��ژⶺ�-�;4["�F��������\8�]��͠bW9Pn��P���}�\�
�!nab�A�,�oNl�h��#���
����Z��,?0�/G�ii�ٛO�.�2vB�+y��P�����7�]��Z�#�xt�l'0)z|��I��K�R��]��<:����>�s>.�!�s����=��zb1i!�A8}���"˄\���Sٽ�{�����s���:p3p��G�O5%��>�SS�0r׬z�}�@鴰���%�i^�qus��ɂ�2vf=����x�B��֗� ��gejo��fm� �Y��ܲ�D��ƑA�N��֐�9b���J��'��)ꇗ.�k��1/�N.�b4���t6���>�9���S��V�����3�v��5̋nL+=�F�wr'ཞ�e@f�$�Wui�1���u����+����}�A��im��b;x�}��^-���8�+]3"���}�P<lu��{� ������$bھ&�1�^q;�Q]�k��ZC d���}z�gm���]#�rh�Mik�!�Jn��Ű��{f�Cv�=��ӝ���}���ݏɱq�z�BY�[n�i_�Pٮ�J1�d�NJ"bh���3��oX���r��)k8�s�pj���!����JՉ���{��� ��7�+#��.Q�T�κ)�I3�0�\x+e��"_Z�ܽE7	�jƹVA�|�.͕�m���
+��t�x��R}w־C�K�&I���٢bX�ݜq�@=9�N�@k�h�^��n�]�춚숌-���B�%�f��&�f��]�rɠ ��< <݇��k���Q���큖q�l`�r�oaSƑ��y�w��r�/keɃ��/���;`�k��f-Z3r62g6�bj#�a`t��k���E��z��Ӏ�(�����o��,۾�a��[�fܼ�7�e�/�U����FS�ԥO���M��{Nnl�ں�N!'�U���ɣҋ<5q�KoWm�2p�����4��A�t�Ep\2����%)٧s
9��}�)5�u"GVmiVU�aw[
z^� pą��w���Gmj���py���vԔjU�%���o����q����&5���'{� �5}|��A��>���b��O������+LwT�#��X9����Ƴ�n��q��zE�[#N�;�P|0v���8٤��FJ���o�8ު�9=����;�z%vnٳ F����N��7�XsD	2'*� r�hط�Q���X�ܶV-�W*o:ˡ񕍅��-JZo,��Kah��w�Gd��p�[9g+���ܸ���\6f�ڰ$�gz�ڮS�zsװ^�OV�����X�q��.�.��0�Xy@u�I�P57��`Q�k�tZ�y�R/���A��,�wz=�	��EJ�����T�Y�Np�-o[�:�(}�k��'�m�}f��M��_{�th�v
M����%����%�����\m�����W#�pbͣ��w�njĊ�&' ����9�Yq;�P3]f.W;7%���e�Ύ�v]��\�R���'wJ�L�ܜ5Jh!�jW��2k���8b��7��������Cv��5l�)iH�(1�J�UjQF0QU
�ER"� ���PUEQUUUV"�b�*����QEQF �L�EEE�PEU`*"��1TPV ��R�b����*�AQL��AAq��EDPIR�1UF*����UEF1�E����H��b"*�EĨ�����T�U��
,DQ����Ԫ�*�DFEX�U�EQU�"��X���A�""(*�����W,X��*�1�������!X�F1���ʫUEDDUE`���AER**�X�Q`*����DEPU��A"������)dDU�7��z��7�Gkf�M����#y�%���i�i�)҃_��^�o��Ʉ��WK��
o���:�6#���ڽ����{sKN��w�87i���;�����}L�Y"��b�z�p����Aw�[��{��̗�J���D�x�=r�j,h[A�J�Br�J��:7k9e��%qW���븈ޖ����7���!N*����%*;B�c���:���k�`E8�i�;�N���������Nf;u�kt��E�H���B�B"�b��<ƨ� �w:����9�`dې����y�w�!3�*ĸ뚃i�6t�O���7$��0N��ҁSѬ�rEww
��I�nLl
\
��`S;��ꮧ}	ɊN�w�o��Y%�n�=�Q!���2��tׯ)�؇\�^�� ���C�Qs)�pr�@96���	Q�|mIVX�b�:�b�u=�Y�W
Ā�Ҋ��e��*�ڪ`�<z�wtrA�/��c�F��@����`"��_U��t��])(,?��>��Rd5Jx:�s��#S��K�['gXT"+���L4���\.j�F`Ԑ�������*��lWUR���dYj��7R�/J_z�G҇L�q��&�C��ݗ
�"�^`�7�s�kbe�NYw �21!��z�ը��� ��go�����g5��@3p�-�σ�W{[E]��:�w��PFm'Oz�j_f��mN�)#�*SJ�N�_�

�rj��F�B!מ�Pl6}�/�h�W��|���0����?hi�g�pWR3���[�7���B�5\:�q�P#�YdLR��rY$�	�.�WS�v��^�gJ�'�����[�A�����Q»q��ʼ����r��
<�r�s�ݎ��^��z�b����[[r���W�:�2Pr�ۧ����QU�ݹˉ�y��+�Ij�&�����j�f�}�4!��Ĝ�����c����:��g�n!/���%�'pƺ�I��Q�q�./�9ՊT�l��f_��� �J�F0A�������F�����]C�Qʞu\��W�4T$�[/&c�)R���{R�p��W��v+���%�=򋀘�V}�+�q�ɷ �B�:�2��*l:G*TD8���u��/[���_ҟ�컪�0l�:q'�Ź2����'aA�[#�za��u<��Mc7b9{�t��i~����i}�������&O=�t�*�yJ�M O��O��6���n��,|��=�N��&q�3:���U��.�/����>{*��Aț��w\
�;�+�&η���{e+��@T
�t�I�������m ,i�(*�4x�}��Ҡu�ub/�i�����S:�^xl��(���w]�%`+���oo��8B#n��QNR�{*0F9sW����͗x�[����g��०+���m��-K���LB��L�M��"�ʉ�˝fukǣ9�����*�K�{"������ˋ�U!�C��LੰP�i�lT����GX��1-��m��#�����.�٣�������N���$p��梽4�.-\������v�����;S��p�9Ӏ�l�3+�@�
8Ks~��p�J���{*��閳<]Bb��'Qjz���Ӣ�7E�^�Ǭ�<lyV⶗m+c>�전PΫr�$zJ�g1^]+훛�����>�J�����KQ"�)g��df�6��yմd^<{������79L콨$�/����w,�������g�ȓf��o�?y�ɛ���aT�sy��u������q�]�[|��hh�S���*��.:�|	ՙ�,���3a+��{-u�c��v�����sup82ˋuC�v3�=R�zoX�\*.��CW`�	z�[Q{��eu�yK�wYǂ�9�kL.����ˈ3x8Rbi�N���~���c�2l�WdAθ���+���=k^��s�s��JK�{�Vm���{{&��{���u}=k�Դ���W�Z�*(#���*�5��9tlt��T,G����������@�D(���Q�q���N󂡛b. ��Jj�Z��o���k(������p�EҦ�mJ�u t�V�Ge�{
j���|���S^�f�yگ9}�] ��J�'Dq��eG��(�>�z��{��_Z���,c&ޚƵ3�,���c�B�lL�\�����/�W�'D#�������4��Ĳ���wa6F��4�~��)Wl�r}�ȫ���P$An���?S���ND����BӰ1�5�WU�9��)��B�u��r9͍��U�Q��<�����`d����D��x=�����)�N���]2v����Ú��x��Nr"�т\c���*ˋ�N�����P��X�Od���_v�B���'n�]4<UM�I�p|�隖�'s���r����6��s{=b�P��B�����V*��j c.*/� ��.F�����l�W�;�7�u7{I{��*Q��+�4�h���}�Wh�X�e���u\���y��/*�l[�@�Yh�_:F�Lnbh�oa�c'���R9�Ǩon��z�Ѿ�ֻ-�)Ć)��ٲ������2.�u�U�pIR��39�{|���l6즋��)c՞w��d
�Y!z3�[�P��㇌xt��f��NQ��V8}+�D{�<r/Cf�h��ɓ���Aڒ*rWC!��2U��.q|���^n�\��A��!�[du�A�͚�a��$40��O03J)M\���͹��jU��LmK�z�L@>�p�dl(�I�}��Z4_�V�z�����б��ʾ\��ǈ���G$LdbFl�B:*�.�3��܂�:��gp�{Lf��I=nw{�u�S�gO��шpJޫ;]G�OC��lQA��RΰE���yG|$&k�ӧ3��V�,z���'�*&;�>>T+�V1��l![��'+{E�Ҧ#�g<�7��)��A�>Ơ��ۼ�nGd�aM�)�..�������S�;I�=�H�����C��l��&m����>�N��Js1�뮩�pjC��+��$'D%k��$��`5�����bLGKu��\߆M�
/�ka��~�;2�K�����НӉ��r���G"��>j<5�P�mMt穢,)�rܫ��U��G���?Oy�G�wt�H���~j���뻖;���sYӶ�:�ie$kF�YaԀ���70�K
ٯ{U$�!�Œ�p�䈹]�8u�i��ٶ���4z%�@���ط��^�}a����S3�WP��zU�b�&Ozm�u������*{%�L9����9:�^�g�d*�x�>�C쇛CL������X��f�k��[7͒n؎�o��ױ��x�m�ȐeCՏ�F��U���A�/��hj�e�2&����m�T9�n��*凴�H��a����lO���Rp�J����{�豱�w*MH�I��^ﯹl�m˾�LJS0�2x��BG}�>�Z+	Vg��� ۛ�㛭���W"�C5	ͮ�p�B!�{EA���̐�UԾ1SI�4���Q^RA׹�IOuK��{��5���z�i%9��EB^ˠ��#��B�Q��������&mf'���:k�ʬ��j3�Pkkm�x��"��\� ^e>�c��x�]U�<�BC˃�g�s����"�E<���ٌ�I���xlhmK>E|��çG�O·�1�u%��~�ɔ����2��B�����K��J���L1BzSz� ٳk|f�=������������c��X�z���[�
���]x�
�T�E	Wٛ�v*1ٝI�3�<&e`{0��Ju r�y$�m*c/A�'�7(;��<X�&M�E|9�����#��9���T۬�Q�&q����TK���[;95]��l�eK���e�I`�94\iq��9ζ0kv��r���#uqRG����3��˾��Hؿ�Ml{P�.���7�Z��d�� �-���S�F�z�@xߢ���#��G�@/ԍ�>�����}sJuN�r;څtv�s#��E�r�*]7biq�l�ɞ�͌��!D�w�#�:�#��J$�_�^Z=����y;
:ّ<��on=��oc;�sdTO7%�ÁC���psK�T|87CV'��3�����!g�C�������g��|MԱ�TbADW��8B#n�����1�:����TDd{f(�g���g��26�'~����y4"ʨ�hW@�36��E�I�Q��HQ����ͬSb=�H�g\¹x�qwT�0�`i��gϩxԴ�]�.$.����O-�*ʹ���<���.H.
���P݄�`��B���p�O�+��k�-!ַ}W���Xg)`�V(=H�.:��d(G�����B�G�u�*6�h���!����uZ�9T���HT��5Q���kv^Ys�"�>����uOSŶ�pT=ex�y�S��1�(l�B�ɵ�.��s�M��0�D����^{��d틞VE����4�c�,���ҏ��pi�����9�+�n ��ɳ�q��0)��c��O��$bU��7�'l���r> ��޸\�-��  ����+o9-�����vh�j�I� =�7R.
�rfu�9�
�2a��Nݔ��5חz�>ʸC�eCE�����Pԃ3��#n��d�F��"���;'�w_��[S�1��
���a{�+�Z8��Jޥ��Ԫ�v�����n��|���3xPgx��2����g@��W6|�ӍuCrvU�<�u�9\�j�'C��3{
K���N��g��5eT9�2k�����U�jj��/�^aCƊ$��{�,o�2�וo_\���5�,"pu3�Ä\�2��;1Uo�s��<��M�4�m�:sր�S�İw�V��_o���R��5�X<�.�W�2��u��&��}�qݯ��c��jSHnC�ixD���4ڒ")l
��8�dC K*=>���p��Jg��:����y#�FƩw�g�����{C�E�P$F��̜~��#d�q(d,�Ǿ��wAIά�ǱM�j�W�Z��1NʺQ�ϩ��v���q��R�F�Z�q�V�+���3~U�Y�,6���غZǿZ�{!w-�J�[����΃�b�����v�C~2�37��Ա�vl���ibJ�
��trͱ�+l�G������C�It5�i�Y�z��HMs*�~G��v�N�r�;���vIK�������*��|�?>Hx�h�.��P��3� R��σ�ޟ1���%(nz�w^ �g������v�l/5\)}�:"v�u���SU#���T�o�m��KA�Ó}ׇW=�" ��!��Z�D�R2�T��ˊ�}dQMȼt����j�9̳�ն[ə�a�"zZB���d�ʏT�W ����l�}qB��c��v��a��gsZ�D�j�I���q�J�k�b�͛����p�U�ړ꜀SS�E��=�U�w}���f.�9��юw0�y���/�,�~zsf��G&KB�C={U�Ļ����y��ȍ��_HȘʐ܎���@���z>���w�`�+ت�Q3�ܝ 't��[K�lK�#l4b���u9�D�BUV��.D7""�	u��
G,m���';�iߜ�b�шpOuG��P�#���[����E)fs�Q
�R���in\��W����:qNyUt	�؈�c��P����X<�ˀе��z@�6��F��M�y�,&"si���u1F�n�]Р�`0���#sC�K+z��Õ5ع���ߟ��W���E~��&v>͋7����U]��٧�ݝhCU>��ҏ���kC���4�T�hT�8e@���#n6U-�<=��Zc6��O4q��m_J�q\�h������!Z�2|�D@�,	�� S�Շ�]lf��$�Ƨ)(����6k�d�����)��g�l7N6�Z��(b��vOܲJ����,;�F�=���|���� �o?����>
$n��;!Ɲ��B�;{'R�*?ƣ���UH)��� ��<ayO�4�l�1��܆�6�e�!�
�C�M0�1�P�m��d�Y���|�� ��l�p�?{d��+)���;=;x�V+�G���@ m��VauE}CL>aP�;��X�d���(��<LN&��4���Y5<�&�HV0{�O��?{T��IԨ��{a��'\`�K���]�ާ8�Я���|2�t�6|x��l<H,��m6�U%I��d�1?�*N�Y1���'�,8¡�+M�8�fPPS��7�m8�Ri
��ܓ��HT5��忞�3��z�gy�����V�'����4�d�>�y;�h��@�o;��f�l<��~݇��@��0�ֲ�����"�R��`�����7��Xb,��ACԕ�{�y_=�vR���cj�-N��Q�T "@TM;x��6�{f��O3����aXVi��M����:��w&�R
u��1>Af�a���4�&3�Qa��Ns�*m���^����������Ph�o*a�����@
�\�3�%b�y�0�AI��
�rɈ�.0�
��>�!�������,+
�Y���6�Y���sh
/�����I<CYaޙ��{��w��vVX����ሏ*��1�Ϥ��*B�=I�<J�;�&'��q���� �@��xm�{a���1+8�+4y�CH�u�:�y�06�����wX��2{���}Ϸ߼���y��}��+����Qu(-Ξ���7�>:�z(6}��=��uȨ�F�-�����YaC��3L� 35[RO1�B	t����@+ �`
���9�o����tu^A���Q;ρ����(36$�$����.!������/\��E9�q�؆���$��wYxv���K�;�"18w��BJiQ+�J1��9s�fY�V��qwkăa놻~����8�՞��������{��I\$�u9+3��z�1[/V3y�-`�4�]�YٜsD�� �3j�v$Ē0�y��N�)�c���������ۅ34�{�Om��7o �GT���,R�zc�C?Z����洀{��.�m]<�i0�6�Cz[r��ʲ�6��]wSU��=�{�c�	\^K&P%�8�<��
�?V���j
���*�$���u
�]
��=�[�Kh�ȩ���:�Ӷ�᜷%${ڣ�8M.�ilv�=��jz��ʙ�ꁃ\�pE�z��&��ǧr+�%/ۛ�}�]�珅��ć�,�np�[�hv�<d�j�6��깘#�~.z�l��b�m�+x�,4&�9c"��2�_Ec5^��@p]��(̩����-����\{WғȤTL�m|��F-�bz1x��/��u��g(�sӋ���ܙ̀&4C���R�"=�!��/��Mݤ�=����᧾�VL���}��P;8=t��}�Ʋ<��1�l�S 1c+�ԃ-��Ү���!.}v�fa�Z7|&�zͶ3�=<�R�������A��X�s��ian�L7.��Jy���Ju`�<<��j�u睕
1�F��5��Z�HṌ���6�S�5j��$V+�9{Ox�ꎀ�hФ���Vk��ym�B�!ۚ́��Oe������}��͞[A%�i�@iE��	�2pd'�'ϻh�+.�=�ۋ���V�N��cp�;��r/w)��X��^o���{S��s̞P�F��m01� �'_ƭK���!Z�ި�sܰI�z@���a�g:y�U�L���9m���2�n��h������2Y�b�Q�\y�3e|Z9ҳ�Éջ�-�t �Z��q*�S�Y�A�]�׫L���( �ꖰ������0dġ��U�I��*�R�cop�_����ڡ�P�< ����k��z{N��X��퇞��7�����kɽ��56[Ѕod��tV�ܸ�D��ş~tr��l��n^��X�ɲ�k��y�.��Y��8�����-��T���m�b� �+_Tv��u��
�L) ��ғl�|�u+;��qث7�1 ��SG�t�=~�	��,�F�Mn׫3͋�[&C�*8)0��')�*�=�^4z��xt'[p��E�-�ZB��,�7w_XHgB{_}����*�(�A`�G�"���j��V�F#EU��,Pb���6
�,A�bb�-*��QTU��+��b�ƈ��"�"��b5���U�)����Q2�QJ����c11�т�(�ZQ�cU\�"Ŭ��	mb�+�� �̶2�U���"�`��H�mAb"*
�6Ֆ�1E1�QD�Ƹµ*1YJ#J1dU%�QQb�"�����1"E"R�F"� �H��"�9J�U-��*���ELj���PEQ�*+JAA��X����"�`�E`�*ň��dQ2�UĪ���� 1i�T�������m0gb���㩬<m��psTΨMi�˫���t��q��? ��H\�������n{ы�</e�WV��˺_���� �n�����t[f?�7�h
)Xk�`�L@�?!���ь�9�B��Y���̞&0�V�Y+�M�;�
AOP6y�	�eH>ٹ퓻��Rn��Xk+:��9�WS��F���)v�=q�0"�=���>a�z��1�s�a��"�;�H(V;��S�L@QM����N� b���~d�s$�n�0�³l����2Tߝ�iU ��|��p��SƔ�F��w��1Q��t��o��a�:��;�u�$jw��'�~B�����i<a�1'��QH?Y+�`��6�P��pP�7�bTXc
���wi?!X��
��8�P���ga.��?j�U]Q�T:}�&�0+:������N��w�@�=C�ON���7�B�o��I��S�'�i*<�tCI�&8��0^!Rԛ9������8��)���ŭ�f��o|>P �QJ�VLE����yi1'�VO|�M[:��Xq~�H)�5?sM (�Y����IǺ�I�'�r���>a_Y4�͟s$�>d�!�so���oϿ~�u����������Si;<���ʐ]��?n��B�f����YY�}��>aQ`oˉ�|��q}���ì1��b�I�߼ɷ������sH|��<@������׺��Á;����9.���������c�����X�Y�Oy�*J��S�)�:�5̆�HV͞}��u�H.���|�C�y�&&�u�@@�_���}�{9;B;���(�-�݋c�d
�
����k�@�>�!��`iaS9a��ɴ�B��7��h�VaS\���
�&0��O3�T�I�6_��?2���Owt�!R^w]�~��s~/u������מ�Ά�Ěq'�zo�H)�O�|�p4��H<����'�=Ն$��`iiY�ü�@Qd����L�I�*�2����Xq<ݚH"��|�ޘ D��d�s�h�f�1��^�������q���Xw�P����r��c�W�M�}7p��̕�o\�w�)>C���'�ʁ��a��冕
�7́�k+��`��|¢�s(bVz��8���x��s��{�"|��{���Ȝo¹{.�<�+)���f'�Y&c���i�{�n��#9k<A�F�]n
�+��]y2_�	-[�j��������눥wxD��Q<ι�N�V�G/���'������-ff�\�H´G�uE��eC'#3�}�W�U�9~;���R���'�s2q�H(k~�4��2c"���J��>���&�w��6ì+<Ok!�H,�������N�GP6���N3�|���	�
�����/6VY�s���A�XT�Lf�q1���1+��4�CiVM�5�fӬ1��n$���������
����b���s�7�(�Xx\��믅���_ߋ����Ьׅy~���I���)��I�y��;�~e�!\CL>�'�VzjɌ�'�$��i��ɾ�0^!R���6�a��b���%g�̕F=�!#2㻌J=[ouw}������B�����[=d֬;;�B�L��Y��M�VO\N�VyY�'�O�v��va�
�d߾ᴂ�Y+������}d�'�'~�3��Y9����{��FG���tDyt�潗�g�i�0���w�M&���&����d� �a�o��V �QI���&0�՘�$��0�ݛI��d߾�!X~aY�?v��������͋�������G�G�{� 	%U@׾a���PY�O����!P�.���XT�_��a�bB���i ��1���pS�6�P��E�6��1�'�Vk�N����S�E��F�n/�� �<&�{��|�a��k�P+����RW���u>d����:�OP*O���yd�����a���Ri
�_rg��>�
i����>xy����}���{�Ϲ�ױ~`�!X-P4���l1<7@�%g�fH
,��2i8�J��{���[gY;�y>�N��Aa���wvu��y�kB��=q? _C��8���M9�/ٻ���۽�y�}������~�z�a��q�L��� ���0�Y>�)�e���'�ʂ��Hw,8��04�X�3L��ϘTS�
�Ϙbu��b���O9ܞ"ΰ�o_�ʜ�p���|��<�w���ކ�W������ERW���2$���d�;��8¾X,�e ��5�i?$��*? T�<��a���w����aP�~��m�Ɉ|�y���='�W��?]q�@ؒ��!s�jkm�W�o��^0"�+��^�r(���Y����� �� ={��2;�t7ۙk
J��	ޟM�<�OlyJk���*�)���2[qWWe�gJ�� ��e�>��J�]�oM����ǝ��]+		�����1��3���X����<"G�����@��)��i�6�a�>;���x�fr��fM�����g�I�+<���a��d4���&�M3��<"����p &=�C~��a�ȫX����riY6˺N�CL<a�)>g����8��>}��R
|����.!Y;�3��0�h|s3i�M{�U&�}E�������c=�����P��Nrq�W�=lU�p��{}�<H2m�!9�=g��=d���|�O�?3p���'�l?2x�kd�$��A�`HT5<�*��k�!�̬rt���B#��ǌQ�{���:�s_�?!��凗솑gXTR��J�:ɟ�!�~I]�|5̒��
γa��{�B�����g����_m:�S�J�sy�<�~���=�.�����|=� &@��0c���M]0��1��*nj���>LC~�bAM0�ɤ:�C{�IX�I���T�B�]�ܰ�Aa�_�S��bN!O]}����j���72kD�\���W�c�zD@c�j��C�J釛�βT�q��bq��H{�'����t�aXw)4y��1&��ͤ� ��K']0^!P���Mei�;�\׾�)�㜆���Ҵ�ݵ������ϜDL,�_�?3�RV�c'���0�w�>Xu�H.˙�Y�J��ɉ�'�'�t4��*z��n�HV`��U�d���%x*�tl����s~��������OɌ�~ɤ�
$�Sg{�H9Hw)����Ci�{C��Y��!�r�$�1���4T1H;�}��ΰ�6[RW���t�ACĕ��.������s����~����@�N!Y���o�B�������N偳�3L���Y*��@�bN���3���_,��a�~La�>�6�Y�LM��� �����f���C7���_ߏ�k�ź��Y�=�ﳳ߬��>Ot�H):�f�u&�������bO���i��_��W������J�=�rM��J�s�`i�'���O'f�z��i�t�����cª@�)Ɋ�4_p������\k^D�n�7�[��÷^��/:���e�S]���2���ۦ:�5�T!��AM��W3tƞI����u�+_oo�����������r�!؇L��-�
~�)s��{�&�'s}(<IJ�W*��v�*?�� ��_��|��m�$i��R~J�B�m��/��MP3��=�C
��g%@S~fI�T�)+=�~B�|�l�>��}��� ?�T��ǽ1�,�Ӝ��}�7���;&�OY1��t��&�|�LCs�Ȼ���>C��6�O
o/̚~d�(��*z�D�fM$Ԇ�C��H)�哎�Y�1�Oνp"�@��AV'����ϻ���u}��{�E6��ă����|��Y��g�y�i�+��<;��*9�k�$��|;�O7�T<5~a�m�ܤ��g̕:��<�R
~@��|�Y�l8�����;��s��S���ֿzy�~�3q;>��i�0�<�|�u
�AM�纇��=N!�=9����V,���w�x�RT+��0~�mE��X,4���bO���m���&殘~aP�J����9�כ���My���9ݿ{�>�����d�~B����bq�C��I��'��s-�+��S~��m ���hu�OR����dS�O\`�C�f�A�����h��I��)���*�7�빗{�ZϷ�7�k�{�~:~d�*q���'̶���I�,8¤���$?[8��
)�O�?����|�O���C�e!X|���?2x������J�d�R `u@��"<&q�m�Uh�w�'�<��|�Vx�}�t厬:�T��2�eg�1�5܆�H)Y��N!�1���,:�gW����+��;�<@QC��hi��$�>3��{(��m�ú�hf�l�9;������?0�?2k({���J�ÿ���AN�jsXT~q��/)��m�&0ٮ�4�Y��C����6ì�:�C�<�g�%bͧ#��� {��"��]�7�)nn������~�Ɉ
/}���Ou@�<9�u
�l.���|��0�c����+:�QH��d�bq4�T>�'�=ɮR��<���>B�ߵI뤝J���7��~�^o�������N2i��w~ᴃ���k��=�� ���!��=T�'���H�zʘ���:�d�[}5�O�Xq�C�RbC�g���&��N 	�� L���L��~�����Tk��3'�J�29���N�*�q.8g���ɱ��� �����;���X �|W�Ȏ����+�f����gNw�I)ح�\��ˋ���k#g�zǼ\;�Ӎ*���E����̻6�l%� ���cV��k���};��{����U׷�O����R<& ��Xc��i����&����'r��AN Q73�Vm ���܇��z�T�0=k+1���,4�AJ��`�����7��Xb,��7�R��g#o_�~� (����̘������i��m�{f��O3���b°��'r����:���M����ܚO�Y�4�ü��
�l�c7�`��Af��^s�ML�&��u����1����0" t�bi��b'�c�=�V,��~a�����
�rɈ�.0�
����~Cl<ayE=��aXT:���o�I��͠(��bb7kc�+�ɒq��߹v����Xw��,�R��g�d���
�����'�z�xjɉ�'\a�38�H>�7�����
�T�⤬�ϲE����S��`m'�+'S7���G�A�gv��mw<�>���υǄ����Il�]�h
)Xjw���
����z+'٬���Y���̞&0�Ն3�J��g�ޅ ���F�ʐ}��N�Ê�H��Ͼ�7��k|�JՏsu,��	� bc��%C#�<& ���m�a�z��1��#���4��H(V�6��Sg`�ӷH�'�1��7��?�L?0��&�;�Y�%K������{oF\o��77�[q<"�|��`r8����k�B��8��y�Ă�N��C���TRzw�O|�CI�{;�����y��$<;�4��dĞMSa�<��;��{r럵���o�g8�HVaS�@�0�o�&<`V|�C��@Qx�����h�I��{�2f�HVK��j��*�s3�8�IQ��'̘�7��x�H?R|}�ܹ��dg�{w�7�����s��� i+<T��jɈ�zʟ��I�?!Y7�2��N���?8�R�8~�,�@QN�a��q�8�Rq��ɴ�'�;H{U��cc�0*=w}� ܆�8������4�2W�����&Ú�|���a���<T+1��8�Vx���
�Ʀ3��C�c��<��E7����AC�6{̗@��� U��ܗ��2s&DϰoК��n�4`&��)"��F2�RΩ���lzU��Z�d˄<�2~�z�H��ա	��oU�R��Z����qG���������{�HݳHW7=w�<��3Ѣ�]ִ㣀�6���_\C��zm��+�=��w:�%��W���xl����q��� ��Q���}���~d�w!限�>aY�k�dwH,�&�5�IUR
|�E=Ag\a���R�3��a�aR�)�&���E�nɉ�f!����G�'U\Fe.2���|�>`xC�z`}�i�&0Ă�ϲ��<Փ���,6¦r���ɴ�B��6gr�(�T��)1����nj�H
/̚��*q��/�ԟ�yHVo���"�/��.���_m���
�{ 	�� ��O�I�^��$���';���*A�?w�񇺰ĞOy���f+�y�@Qd����0Ri'P�l�2����Xq<٤����u���c*/��+��~q�L "@Y<q=@�:{T1=d���<�SL>a_�<L���?2W��\�w�)>C��p6$�YP6y�5�Cܰҡ]r��k+��0P�>aQI�/_Sn+��i�[e}ʾ ���ǅ@P�Ӥ�l8������H(k~�4�:Ɍ�Z���+��=����'��=�p��
��Z�r�:�w�i?$��}掠m=Af�e��y�?UumP|�����{���Dxm������)�0��Lf�z���T\`T�:�C��!���&��E�N0�����Vo�LG�J�aS����x��6��ro�P+����ӎ�ڷ�f3g����~W_����������I���dSi�
����0wd���B���}�O��VLg�=q'��"�S5ۦ�*A���ɴ������HJ�+���߾#nFn���v�v���0 ��'O|ͧȤ�4�M������~d֬<;�B�N�c�c%@Sgy�������O̟�퇦�4���ɿ}�i��W��;�)4���|y�����}0T.��[ӿo���Ȉ�������)e���N�6�Xj��3�4Ͱ�����4�g��Co��O����QeaR
a��)4�M2c��Cĕ��f�z�gY>�8��%}�w�(��v�Zv�����c�ǊΝ�I������N��������
�Ag\}����!P�.���XT�_��a�bB�;��AOc1;�)�H?�~��E�6�V_�Oe1Y�F�=F��*
(�©�	w�{��ŉGv�F�v�4r�G5��	�+����݇�{�ٚ�\�s:��X�aM
��Y���:�CSl�h.�I�u]�.UV0�ǽ� �,윳�y��k�Aͭr�6�����ȅ���o֜�vj�����}����3��������� L{��߮�"!�4o�4�~B����5�(��y?SHq%z����̛@Qx�7��x��*O;ߴ���/(���l=a̤��K�@���A�k��=5�����o|���~���R
x�O>Ȼ`��X�����v�H�������&��&����?!���1�Ձ}�}_��Pܝ�Ժ�1�s�Q[nͦ֔�M�����s���F�",@�*�E)�=�Mt���aF�x?YU���jv�|�}9�[~��K,/%VJ�N׮��
��4�|��CÇ���x��29�=<�Ϋ�Ո��؊���-ͺ��V:O���g�C(n%�Β��]�ޥ����M�Z푛���㇃3��������h^׼�
��t���(k@3�6��d��;mrs���g׋�^��q��{]trzB�r�J�!�s4�g���m����uO^k��?&��[$R�.��P}�����\)GC��㛣�'!np� �n���ze�u���ݲ>����U��$i���>v�o�^�@���/��,n:��Ƭ�i^�[�&�'4�"�C����eE�Ð��7�[��W�u�(�`~�Ol:�;����^��X�=��=�X�dU�gY�p`��b���2Xb�T�/�,��7��	˃�����n��uԥJ�&gD*.�ke�������Gk%����b���ũjr���:���F
��6���?_fg���b��f�y57��	��x�ٱ�EdEз �츘ea��#qQ�C�b8��vui��y!OʱH:�`0�	s�4-�5~��4���-
6E�����ѥ:۪�����nO�0��Fi�&��U���L��=����7�W�ȹ�#�z�A�tE_D���	�3]򥊗 ��%�\�s�� ��.u��>��M��6j��X��x|��sػ;�������%\��
Ŋ�2�S(@�r�9;짛u�X��=�T��[�{���u�����S����CN���5�\�XχU��~P���u~s���nGœ����kL�V;����O���C��MX�Z��H��p��HV��)"ql��e�x����"�Qȷa;q��:qN*��=m؈�c����=��`;5�c�iy��1��#���k�{�G���4G_�w�-�쐔H��a�iF*�NhÙ���Ǻ��w�ЯQ::�Z�B�Z���Gk�g����)��c=�~n��i�i�K޶t,�imw%ԟ��t�+��ƹ�b5 �n�ƅ��*��!�E�jQ$�v�g��̭���cB}�f�rN��{��|<1f�.�.)3I{gg'gt�
������h��}J���G#��׹l��mb�nK{Ar-���6�{��Y�X:PV~��� 729��f�p:�}A�"2!͊��Q��߲m�Qfr�'~�gfV��)HH��9��C���kb7f��u7��8��r����ו65`��/��7
|od՚ܳO����5kkOd��D�L��§����y���d<�UK\$��dt=�-J�upue�|�Y�-����7I����q#}*LE
CmE��#��2՘K�qA⚱��w9�QP�ե��3�3	��(Z;��[U�-��d��C�J��U�.�o-P�y*�Cx�����Z�=5P��܈�yU{(ymB�Ȅ�Q�Fa�qN�����@��
�;%�9���┃sP�߻��!�T"y�QRw$�E\�K��u�~�����IxG�Ԉ{�a9���X�S>��ƥ:����=Q�U��&���w��mˋ�hR�1~�j"h|�����1�όt�[[s`T�2-�a�@�,�VZ��79��!�2Gݸ�	�y��E�>xD7Pg��5;X��q��R�u��R��,�%9�z�d܋6����b�p��O0v�v@E�-����GP�w���6_Eb�3�u ���q���R��ڏ�L���̋���\�k��{���y��P#دc[o�=xv���V�4��]]�T��O��;n���<�쫤s�ycG,T|7��AJ�7OE��Ȧ�`cu}5�Ϻ+Cbj�2��UIs���6��=���%��ȝ��8W�&uڌs��..':�,U�5� WƟ����;�����;�u��������k����C���UhU�K̄ըX�[.�HEOv'�sv��.�]p��Xή�!�}�*�֛@�Q= ���jv�څ��)/�0I-�ɐ�e(��.���FĬ@�� �ʕw��>��`ۖ���vZy�y�sGj{�8>�[2�7SmP1*ܗ}. B�N� U{�\(:P�5;|�u�����IGC����gv\X*���� +�����TbA�G���N��t-���hoV=�5����P�;����R�utùdl2);�[d`���U|���=�;�t]����¯z�gJ��i_C����2��:����"��U8�u�ᣬ�飒��Ʈ�\��wm�t��:�m=�f
���M�(��T��M�:Ci���xDvT����E��͵��)�p���]8�qɗKB4Z$A��.mqj��ǣ��Y1�z5�=$=[H���unq��YMc����t,��6L� �/f��A�##M´]5���7Ĝ� ���',� ��0]=�x���W�v�p*�q�K�:�[���[����޿;�ܖx���sV�o\��U�o���冂D��V�P;�^U
tof�B��/GhO��r\�)��GNm�	��9��֎���Y��m��*yܹ|�P�f�U���:��.�s�d��Y�G��
��������Gq���+��t%��3��*�������}.��wʒ:�/y�X}��GrZUl�o�R�6̣*��עz�pS��j`F���`h�| �mɜÏ���,f��2v�h��¡��d�᎔��	i��+�Q��z�Oo�sG���m{�J�<}��N�s�W^�`;��e�ڤ޼�˷RE�R�����]7B�^-�m����ˢކ�Н�s��>�ӡp�e_A�[�ĎԺ�vu+�J^䢦���nՊ�7����eH]�;�{�.}�^�t��m �nj��y��N��ȑ<�ef�6^!�� �%r6�$D�$�o d��vi盞�w_5V3��{��ʐ�$Ԣ�b����w�%������R*g�r�<�?s7�,���=�nUɫ���;���P%gn/\�r�H#먀k��uv�nnZO�K*���GGٵzuQ�S�x���yWȬO;w��ۃ�h�f	�$<��V7�i*�d�H�&dɜ���
{��B\��o��'Jet�˔���:�L��n�o.�>������qwnX~�[�j���a�OfeL����W10&yݑm�Pv}\nS]΁�Y�����v���г��Sv�D�/M1ê�I�d�kIR<�g��@ӕcKNʎ�C��{�e7��kC��&��u�Uv,\V_9�:�]�_kx�9�x�.Ӣnf��y�֤��j���ɲ[�f8��[E��_N7��E
�8���uܜ�^p��ӡ�xL���t�:��Kިs��TZ�5��s��]�(��3��+����׏�iI�(M�5{��z&·���6�3�E�B8��lع������Kv���ݪ.�	��ug��Q_v��0�;���o�fuO�R,���;�� ����1T��I�r��{}����d�u�h������EZ%͆�G��J�NWCs��	ٲZ}��߀��q�Wܼ��gc72�uk;1�*���m�1�$���=0N���2�tv.(3�n��&�s�{ơ�hT�mv/X��*�ه�M@WfT�s��k�|l�[;���'`*iU����vs� ��{vAO-H{���#բ���t�5'��w�Y脏�M�t}u��w�P����Q�27w���
�Ƕq�AD�QQQQF��-s
F#DEEQDV("��X����D�A�1Q����,1
�����ň�A0QUU�(�������ŐTD���ETEE",TTƌX��.4�̵TE,b��X�B�"���TEF",D*�UXȪ�*�
�Ҫ ��1UU��e����X�
,d\KPb"1��
1E#Z�"�h�U-��UU2���Ub,TR*������T �DX�Ī�*��DDX�0U��\�V �,QPkV���F1���ʨ�U��UEb"*FT+Aĕ�X��EQb"����DAL�U1�*�bTUDU���(�DD`ֈ���1҂�b1D�V����EU"1EEDb�,�~���z�ݾ'����o.>�C'	��d��(��F�Z�]�u���-�h��G�po	��
r$r.蠈�[���/��^�� �ެK4��v �#�����4�� vX���FYs��~u���׹ş\�^���Y[Q��Ǻ�G�T7�6��{h�[^�,�9g��{Wn�?\��Hر2�����o�W�dh����	Pp�����~�tvh�j�I� Hz+jH�{�%�W}��!�Xx����o��j?m8���A�']�[�����PЭ{Զ�0D�h�zU�x4��c��'`ݓꂕlhk�m�����W�]�Xo��-h⚈
%T۔�z�)%�&]��iՏ���l���~]C%�ι�� �G.�B�R�I���[����J��D��k���'hX�k����ET9�2k���(tK���y�ܱC����|�-NT2'm�Q$<B*�UѦ>UD��t|8p13�w%/kONP'��K;�供R��;S#�6E��:�IEz53*\X�:#�\�m�q}1���*I᩹�{�TX������y0BS��{��	�w4�'�C���0�&����l�1S��r�Qpp�x/g,Ҧܮ�1�J�YO����m�b��K�����*��R7�ݞ����R
�Φ;&����k,�1�n�*�M����o$��P�ؽd��Wn��I�u��(��ʱ!J�]�f��{�����MN��_ ���z�wưg���Ѳ�>����mR�""D)��gD��P�mf����|�?���a�4��yS����#d79둰U�R��@����O^��s�ff���.^c�x��Pc%A�T�i�x=�$4���,�d
\]�8��3ˢ���-9��u���[r:��J^�<DF�rG����ɼ�9���f.9�i��%�K���}��;&jw[v��b<}f���"�h[�t-߭}��w��'�S��i�ie��ʰ�T^� ����L
DK�@��KF2j�G�h5q2	��^Ғ��/x�y!�'���MPNk���-Վu�q�	T�/k�b�}5a�"�IvWm���ؾ�ܮzؾ�f2,�p���T���a;�[����>}��j�&�l�t��Q%t���2�Իl�^�
�����vk���x�uQ��O�>A���yi�-g�W�����ۆ7l���}Cfh��ؒ#��5CkV�R��\�U���P�̌��yX����0V	���+��mZ��u���ʺ"!�G'vR!�(`ɹǣh�	).6z75���c���}ƛ�u�C�\Ո��1t_�YO�R�)�3dqR޿J���?o�
I�>9m~��c,�^��g]b����]�a�� �9�G�
j�*{���d7 ��u��n��v>�B��;س�u�q� eA��x(z�贺���9�C���C�"���X��q�s�8�W@����L��Wd�B:�I�(ک�=�����57�J.r�J�BTD$cJ��˽��u�\��L�(J�8sw.l�5ى>��p�J(L�h��q�h���Ͻ���r��\���v�Z�A��g���Ŝ���mH}#�v�����9�R�E-��ڐ�ɬ��>Su�|+�9D3����R.vH�
���U��8�ׂ���¿=&�"�t��\��1���$n�W��7yhkǐ�]������>����P⢆�Q@�z�X�_�44���C�8����|����-eZ��Ҁ}��!YDu�K�sE��G�%�U�L�� /�VNQ	��9�/���
�M�OØXTT�z8GR��S�9
>��[L��Q�Z�Y[~�η���p�p���|�ø��v�MT�������p����]n�8M^b��uEߜ4����j��y{ƻ�'���p���:�&a�e�!70�e�r2�b�&��d���nv�&V�^�7sp=�Y����4,�t�"dO��<ɏe�Ʃ�+ü��-
�=6B#S�@gR�^���]V��I�I�����{��Z�r95˱L���Ȼ��2V�rsA�Ƭ��wuʀ�Y"���M�O��ٿ� ���?��/�H��|v�ӂ�#,�xU��-Ɂ0�>��b�f6%�I-�ֳjEE��c��ؘ�j�^�?��m21�{X҃�ǌ�-��|s�$��Q��D|A�}����;7/1٧N��9��ߎ^%?QPQ���/��,��E#kC!�v�r�;��Vi�y����&7��HrÕ��E�� ��|ޫ�����<ϺyX��dԭ�F��.T�}��St�D;`��+b����^L�v��\\10�gpˣ��t���&Ů�ޝ�}Xkk��=�p�(]#^���-T5KQ�ѨO����y��n`Ŏ̜&k�ݿ`.�FX�{��x?��{�;DE�҈"�P�)nplڑm�%s�'��y��.���"�An�[�+G�D�_V��IU���e.\�ũn'H�H�g&�(��3�m��������u�=��Tߛ�bZ�q;,ët�ۤKؑ�.'j��T{���q�nz���
TA�L����	�w��5�r���6��"�N.���#djM`�W�K]�)]�t�|�M�Gݴ����5LZ �)�b��A���]
E�zv�Pİ=�$��X�Z��uR�D���xx��ñG:盞�g���[�϶pTD�מ ���u�����H�P���F?K���T��;�"�S�;��PQJ��Fzv�<}����_OGF�b�_��#mSɡ(������S�(?+aO�}���ծ�h`���iU����X]h#��y�;�������W�V�Y�Ϋ,�8�B�N����.��:ȫ�Jp`�M�@�m�'����'n��W��"H��Ьd�~>�S�S��>���&������R�k=��=�m�E��Y�oK}a�t�B*o�mU���/�����C��X����լ\p�IFS�+hfd��]]V>v}G(1u[�3��F�V@���ѿ5b˯?�AW��#�#dݛA�x�7,�^�U�c�����N2.�#P�1��]\ 瓮�ջۜ�{55B�o��7w�Ya+>�L���*�|�J+�M��x�z,a�#oi�� nq�"�b��}E�Dڱ����Xgm����mQɣ/���5�{K�FA��6���0�'�����/sf�g#DDP�ufX�BUj�:�ڻ��g�
��E���{�4�}tJ�̂[%08�N�"�]ffH7�ʜU:��F��	��t��0U[q��wDص�1�5mb�^Y�~g_����5�����ϫ'��5b䀼Y�г�M��O,D�=�x{ë�.�Mj�7q�ڡ�;*ڞU�|2��u��?:8�P�<{*��9������ȝ�^�LG��S�݇r�-J���ډ>x
�"�eW`�����_^�C��hf�m$z:1�
s�tڕc���jdu�E��:�K�Bu*\H���U�Cp&/v��zd�{�W�J�<Ǣ}�<���z�%=G����L�sO Rz&(�VK�1v�e̕��(�y�%�ƕ�����C�ppu{J5�<}*y膻��x�<�EsHJ�(�Ct�Fy{��`H���s';������H���M�b
�kq_��xu���k��â���,ެ��籙���7�B�K�>�J$;�������>dq�~Pyg��.6n��0��mO	��6ڴ�3N�Ttq��|�О�<DJj�)rG��t��B�S���ҕ�l��ٔ�gj�>AAI��;Qr���{6 ��CBx�<5p�^�ҏM`��Y�p�f޵*�⢢����rީ��H�r|���Z1�P��-�y,�ܖ���B� �Ԉ'�ق恙�K������sT�����Z���Wf��i�^w-�w�7�;{vb�md�"VH�hK0L�,Zm�͡GO
T��ؐp��	�7�;
�~ԺQ�s���x2�.wuω�vw��s��U�suiL#;ں�{�����j5���o�e1��6SXRc�*�>
����X �w"<�ض`��9�[U�'v���ӷ��G�2��}�Ohا�T
���uM���!wM�?&z7��G"'"%���V����A�,f�٨7�L��P���#2B�8d�nr��K�W��=o��%�i��S�a��~��l_��660>��4Cñ$6GXh��KV�Q�Y]C"5�����٣o-�B0��K���"��8��n��v>�E+1s�~�;utMNN�m.�i����uu�tQЋ��)Kֈ���ǋ���*g�N�n�&x��q�pf��H��;���~�`5N9M�*����V��Ң �Ƒ	2�`_���
`$^Yބ%���U���5����Ǣ|��
_c�5��u=ӄ�Ca_���N�]~��v�Q��OM���Ķ/7i���mH���K`PE
�j�!��^����6�(�k!��.����j��L�m.Ř���OL��sP}i�X�I��U�P6n�G���"�Ы���UX�����:1i�U�	��҄���Y6H#�Nv�Bފ<��t�ZpC����|�+\�D3�J3�Ԫ�F�SG�*����]�;���S�V)t�W���<�}�v�(��/[m�7�3�,Qu�����I*Y|�<�n��(���x�¡R�x{�މ]�;�1_<��ݟ�\����nO��NTڗ(QQ'��bG��j:wc�X�K���(�r����
��XѴ����(���Ry}��/��dH"T8���ڈOJ��_D.'�;<��#���x�ب7����x��U0�l'A@ K@�p����L�EH�U1*:eLԷ�wW>�^���.�vk�@XC�~_;O���J�")��7S�@n-�=����@�xZ����YF�1�fI	Eߙ���Xg�UԜ�c��ex���P~��n�(jm+ζ�����S����P�.���n�|��Gt�H�0p�����@Y��rڄ�ZC'�>{f�l�7"Uэl��-E>cHsn��ǌ�/�;���tT��"v.��&��ee�=�n<|���>���L�y�?{h�Rܩt��"�N���9{��]���|�Q��@a��Aʱ�z-NA{@��_@��}5��}�4�Y��]9Iõ�V_U�K`vd03�^���/=D�m�b��&uڌs��~/T��,S!m�r�_��K}�k]ċ<�D�<w����|V��T]��EL&��gięEf����W�E��m�U�鞃��q�*س|������(����A>r��+�KL�9Y�i[��>���g<�
XI5�w�u�=�����w�wɭ2�j�:���qDɱ[F0E��8Dz��9r�LV��?x�W�:�7�薛��z�mڸLK�X&c�+j�ʔM��v��� #�ZlA��m� �Җ�$��p�5�c ��v^�o�ԇ碌u�S �J-�:gj^	���!��@����
T�c3t1�!)ue�z���!��J�fJ�x���fz8c�6tK�%ęqPmD.٣1ş�1:a<�{�qpH�����)1�..�t�خ���]�o(����*�����r��pИy]SP,NWG�=������R#��)���6Fڰ�An��3��q��iu�3B:���P��3�P�p�a�^������>�o>d�����y�pk\[<��b��˪��i>��Z�{�R/����O<�:��0K��7���tq�9Z�Nҡ�����D	���.���H똂�W���..�H�(��8g6N:�ѻuR��#��*Ӌ����T≨A�*<Ӥ"�z�%<@B����#�|�f>���N��,%K��*��S��q=��4m��pg-��*�3w�2Y@���o�Vdmg�`2����́5�3\���f`�һ\��`Ț��S�����pɹ=$�C���!�ew���L��3�yoL��������ӯ�&+�C�Vu��� G]�tM�7=p��s���kչAΒ�	�ѵՐ-�;4l5c%ע&/Y9ur��o�-�b�t`��>�.6,aN�`F=^˫���K�q�d+vX�6+���m)���2F̼фm�^34*�"�x�TQl�^B6��sw8�Z.����M �{�aI��r��gs�t'��226gG!^�26���9F�&�E��2�Cu���bw�̢g8�%��Tٲ�ݙS'ch�J��DŃ#yT�	� ��=�c�p�<N^ြ�}�s�ۀ�y��V�E�NÇ9]�L��֏D���Qb(vPVh��r7��bd�}-���r26�Z��M�W�>�jdu�E���E,
O��fT���lt�1o��S����w?IQ�0�WG��*?]]_����	M����}b`���Ӛ��j�e���r��ϳ�A���VD8T�c.v\���	�]���~b����(xˑ6��lW�O=t*��s$c�((Lt�R+��d]��
���k���O�m"-���Wk�j�wV��c�ka�mJ�둋E�D�Xn�`����*;ØL"�%���&հ��<EG��h9Q����A�����+�7H�-�Z=|s�6���+T���2 �6�Xq��L[����N��[��/sOL�
);�ڕ�l����x򩀇��� W|��U�P�d$�>�݈Mt�H�Ј����y�5�k��i1M���K�1d��E�5Js˫��ꨚ읷��Uuӆُ46-�}oݷ��ۡ�C����&�}z�٢��{*�H Rg�:j����2ܠ�ZTb�C�hs��@�:yG<���{�X�������=M����O��v��{�����o�Pd�^�L�������E��'m�:j�01G��|<t��#$v�ݍI��]�oCH���Cc�{���ooU���	)�Ӛ��M��� \ܱ��V��\�1W7{\oᡮ�÷��0���mo��oB��y�t�W;})��x���j�iG6!`�t�|9�#��qGw]��F���g<��0�{]v{݋�"�<U��9���zI�4��|�*"U��h���C	�D�ZεAu�c�]tȍ0�Xnx�/ފ{T��b�-o��
;����4��J����X.}��a�W+ON�)�{��кȰ7Y��5���77!i6�#���)n�sl�h��!Y�͡�E�p)ni�o*R��NX,کQM���u��L X�wPb8��aH��[g�	�T����ILtum�PN�%�%]��G������w�����:t)��]�|����Ū���k��W7to�����R��&��a�ྖE-1gj��׵��L��Mu��p3�����x��;t_��mnC�sa�q�٢�q���oo,^��*Q�+�����y����ä���0d�-�_ ��->�EJΣ�^7
�z�.���l�A1[���ZUϥ�՘s�Q��KIღ�����GL�e3�*n6ᗿ
�J���6�u+9;�e��<�; /d,�p��3QL�u�
�"�zb�{����v�z� nsX���+��^!�%��hz�K���-����Y����ٯ%Y�$h��Ǽw�ト��>h���L�g�Տ�	
w�GG���y��=۹��p���d�;�yZ�0�z</=S�n���~�K2�לX��{}0���E˻G>:&O^�����c�t�+���sO���p�^Rk(� w��j���:��sN�����t�D�v���
�pum�K���W%�|"w�iq���Q��#�m��G����S�e�a�[��E��:0�=���}�9�V�{A�{�f\�f_lM�{��VvZ�)m���CWizC�A�X�� �M���<�mY�+��7&堡�Yw�Y��J����@��n�]KV��ѽ��;����y��Eh_u��v������[ן�TX�"Ȣ�"�1b �PAX*��,b(���Ň�U�QAV
,� �Q���Ab*0b*"�,`����*#Da��� ��U��H���[KT���"��EQ`�D��b
AU1TEE�EQE��+��cQ���EE�(�TU��b�R(1UQk,Q""+FEEQTU��R�E�"�.4DDrʈ�X1���"�!Z"��QX*(��"�QEUX���%�EV(�U�J*�AX��**�QF ���PT����AE2̊��+�U1V*ETF
*����*�X�Q[J�QX�((e� �5�*�E��b"�����.�1�N��}N?D�O�^��f�����,�C{�b�efǭmM�s�84��޾.�d��*!#�o�d�_�� %�EO8���Vm�<h������r�i����F��UL_7C�<i]��o�h�_�n�����`�~&T;�,�m3�1f���geF
8rP�`]���[�٪!C������x�C���)瓵t���zep0��G0xe�ȴ��T�:wk-�{|�M8�1hC�g�9�/CO����'ɠ\CU5���&�B��14�ϛ�N����FD�,�C�1�^�h�X�eA���s��ЕL3��B��y�'�˄����s�G}�ߧ�lҽW��E���^�x����O��U�>7T���Ass�n�*�[OdMң۶���d��;$�ӛ5�6K�uZ���J���\%#l���l8�+���#��K�iEQ}����zB��b��660>��4^�!�r9��T6���LdrZ�}��CxM#�!�h�
��p���J�v�a܂�:��f�+^�B�Vb�b�b���0��ީ*�y���U
*϶�.�JY֬c�v���t�
��O_�����L���M�E�V- ��Gj�f�H�Ѫ��,z���;�ֲh����/!�XS̀Tnؗ0�GX��3K�����m���R��L���T�e.+sw.^����&�'�ѫ��s�
i�c�N53��Wo]�p�t^���S6����<1���Oe���~��v���Ul77�J�	ʿmZ��*"�1�a:g#�P�V�_�(�LS��)������*�@�&r�]J �V����V6��H�ts�6���JVm����fc��aYՎ��ԋR:�($'Dv�lC�)W�z��,�5�Z�yf��;r��RJ�q�����veX�sPm#t�<�NςS$��G�Z�fx�F��mi�N��ע�P�,R��{���?g���7ρu�S���9�/���y I�|�,,�b:��~Ѵ����Du��y}��1�Ȑ@�&"�������ot:.�:N���N;��U�f�N��@���=/7:�lE�����5x%�X���|���e�vk� ,W�~����Z�=>�@/yJ��qh�S8�����e��@S�ep��h���d]��= �J�<P���9�^�@G�i��ot����F)2����S�LX}B#�=WE��%׸(��m"��2��8*#,��v���N��W�;�8Nr��]>,�����u�y��-c>֍Y�i_��ź�2^ɂU�V��=m�5l/VY�����δ��G+���; �.��h��{\���_l쬓.u,��̣�@��l��O�R��'���#|ʾ����Wֲ6����Ѯ#o�y"�*��ÿ:��[�"b�G�@{i���Ɣ|���u�v,�>�b7���F������U��������n<C�6uȽ�D<7|ٌ�mzDK�?
��j^����������Ő��k`�J�)*���9���_@��}5��f��P��$�8�<�����ו�]��H�қ��K+�f!X��g]��,�qL��um\uT�e�k7{��͗�IM@���d�
i�KBR5����=ˮ�1Z1�:,;Vws��[�;��u�,d���H�k��������/��s��P8xʁ����F<b��u��黗�R5���s ��E��L�K�L�D���]) *�U׊a��QN���ތ��qD��E��/�K�x������u=�7@ĵ�tK��g���1�on�[~��K �R_p��A����LwK���wM�:�
ƻ��Ĩ�G����'�Gb��o!z!��8#D��;�
����F	�/����a�S��_��(,�;	J�	-�37�=@ �THIX�9=��Ѽ��C�v�u����!��R��9�d�0˅ Y��U���r���B!ѲO3�d��iW�>����L�9o�C ����O0�ق�r󞛀;-L{,e�xK]lt%�#����g�}|x"�I,\����ەx�^;�#��,�`��6
�fcf�P���ʃ���{"�C2�Iq^�����}�`�������S�y�#*�R�-u=�)��DG�y�J\W�j���3�^<���^{�s�nAJ��Fb�WLD���-Ezk���ԃ���|m��N|v5m�x����6���0���p�\��(EAo�m)^ !^�$T�r|K���x���g`�oy�N�� �C9�����9AΒ�H�8>����`7Gf��c&�U�f��˺</-�w��`_
�*FAW�r�aq�x[����e��preA�A�p��=�{�{ufj�ė'�޲�����ڷY>����Ebu���Z2���-�Gnq��7x�Az���m�E.�=p�y_B֎)�73@r�!�##�%�۴�O����P�Ğf��W�K�Z�qS�r7�,�s#�r7��z�`|TIb�i�b��	� ��\��muLi�Y��ל�#�B�b\�X"ݧa��=�|�����j$���QaVڮ���@�=	e�0�/4��R}�=�?o .2H�nJ��-����kbOE'�̻k�z�(L?;��v{��� �n�q���\���d�o�+��q���^�c�lZb���'�4>��
y0�H��yѩ�&��Gf;4af�� �R1?}����/���D(C�OC��-Ntڕ~� �1ڙm�nl:�K�r���n�����Y�����H�#�V��N=@�*/����]_�֘!)���{����V����nt��KOoMs�`�_/�WQ��+×/�pppװ���r����8��d��.a����z�{����W ��P$An����PB9T��>�Ȼ����5��Ǽ��N�ލ���z�x͔/onZ�dE[U]�^e+UztU��$��h.�����Y��qVz�e��t���]'ٔ��z��e��'_�gjb���W�T쨺8r�&�͉1}ҨF������Eң�F�q�3R��E���!�؆�n"��n&�q1j��/s_ ���R6�LfEEGS��6��;�0>H�rBh%�5vz�.��T
��&��^���>G�2i�ܧ\B������+��*M7\9��Ǭ%Sa�.a�RVZ������D�k�T���/�>K|"E�]j���U��^&:���{jݍ6������v��X��{���->�|��{vM�*�n_X�.�bsnǴ@F{�OzT�	KĦw=s73��k�*�~���3'S�0�%��'��w�x��!����I�u&����W��g�l�H�Y��v�~�s�w���T����B���xPr���~�
�m��e#l�Cs���)�nm�=��Y�vr�� ������lXN����>��4Cñ$6G[F.�OO��|1é������U�̉�# �r����w�����]��Ю�������jv�b��O�u�:Tsk�0n}�E�T(���-�ۏ�:qN*��=\c��Ho+{���jW9�0����<�V����.��`����A]��X��x ܜiXM	Vn�*�j��0WF���[� ��9Ď�lul!Bx@���"`�}Ǭ��wƞ}�2ϊ��bN�µf��o�����G�U�uN6�XR:-�A!Z#�V�94��@�nnE���3�;�+^�3�d��0ɮ��	ߑ���z���qr��^���W!Xd+4ziq+e;ۘ�֮������oѵ��.uɍ�K���a3�>�d�3��
�.������_�IC6^m��S�F���@��~^;5�p��箵�����N�G7gDX�dH��ƌ=㷺=�#|0���Y�!��kgu�jڷ��t�ǚ=���5�n�4JW�4�f�v�4��Q7|Z9��H��1�o��<O	<�
�ܭkOjڻ
�+�oj��)r�շ�`���i�7���d�\����zWZ���z[��;��s�+n�;����B7G����D�~�-E�.8�H�8��xˋ'�����w)�P8	hө�����M��'һ�ի#�U�,+�R�k���]) ,*���\\>g��P�V�
4��)ye��=�T�N3��i,�����S��h��ʙ�,��3�*��z�&E�	,�0wq�xO2m0�(��A긊-�d�E]I|*`�����HѪ�P�G�l�v7i��.�>��	�N�1qP�P�1as��=����_e"/��cJ	����bOk�{�F��V��:���`�y��2�z1� ����r�>|U�·"�E�N��Lt�"�,������0/��+�n^x�� [veH�H9W���jr��;H۽�o0���Vv��Kkof��O��k#{6*EE��Y��وW��λQ�{+i���G4z��y�E�Xs��e���$!@��gf��g�Hp��tj��NLftS|#pf��)��p0�W�����2Vˈ�����D�p}�W��q��<M����i*{���;\�HSγ9vE�j�v���VX��m�D�X\M
�(T���e��.!{�2b���a��P��s�k4L�l���:��#�x��8�����T��Y/� ���E���&�<�#1��sv>�DI��}X��f�~g��~鬕Ӄfԃ�Q�����Ct����}č���g�U�7py��G��TJW����)����ޑc-�~2\���(�;3����M��%�
K�H�&��xK���p��� OR_j��x1Ӱ�|6��&;��9��u��wyR�e�gru��ܩ奉m���>����P|���+4`FJ�X�����_OGK�#�䈑w�f��@�3��+�q��yB�1j�M�����*1�n��B�A�')��Ȥ��QW�&�M���3�m;ȉ������R��:0MJG)�/�S�1��JDx�y�H0���
S���
¹_��NASp�T7i��!2�;#�bj+�M��R߬�l��yV��)٘�^�N�oi��{-uzh�
��=�j�Q�I�"���k����Ez�(�zǋ��Ww��ac��p�0d���ߣ�;U��>��G�|1j�S�O
t��5��OC��c��뼾t�
W�ku_�εo��f�؎���f .�ؖ�ޅ��:Ӆz���ܶ3pv���L��\�ƺv�{�j�,��A�[�X�0����,>��&;���vD%[��4��e0���ᘦd}p���N������`oX8�M�h���ܫ6E�l͹|\�ZzD�Gbx�u�܍,����Ŝy�I�{�ɫ��^�P�mEY���%|��:��[�l���ӧ�𻻍�Q�4���ڜ�Y��i���;�8�����5�W���:��N�,����\��y���cg5-�B-��b9U�f�[,�s#�r5�z�`|TIb�i�\�6A�p�K�̕y��Bvq���"��K��*_{X"�d8su�})U��n�Ix
��Y͡]k|H1�wh��V�x�F�'�,���M�W�8�L�����qؤ���D��\u�a�Ocu�^�df���ig�ip�=�����{����mw��)`��=O(��si3<�4L1�J�9=ڽ^�'D#U��G�5�=`�1HY���y�Lͳ�%س%F,�!=�� ڥD�̑�Ԡ�	���*Et�M�w��
/ڹ�%'hBR֘����]��C��S��i��vy�{T/%��J�3���wY��t_�I~�94���R���oWs�^�#�:r"�љJ-�}Z%C�qbY8"�gjb�8�U;*�ᑊ�t��l�m]��]�wjY���o<��%�+i���䑋�*�3��t73+�4��gT�������k�>ה���²'ֵ�g��=�wu1�]G)uaF'�V����D�����iq��h������bL��CcI��F0�j޸�S��xyͭ�E��ԝ�siP��ǈѴ�Re�ʂ�2�x�{6 ��y��l�&�WVF=��v�s�Y`�h���样���A��ҞK23�` �DK�@�}�6�el�&4a0g����K�N��½���=�J}�^�'�7��';�1?yM��o뙽�b��_{��g�w2��5��.��iS�x:��C����F�>�*��I����r�KԺ�)^�Gz;����+�1��_PY&����A���_���CE!�Dw���7�����j�ǺT0�h�FK� ��8�`��vF��>��4^� 6G[F.�aN�z,�^mf�;m�W���q#rT!ت���.D7!�q�ȧ��~�� ���H��ǪbRy۸�䅝��Gg��1q��(2�d�Rεcv��y�t���T2��$�W�w��:�Iy֢`��)�+|h�	���j������)�gǀ�g{�vs;k-�ek�d�c���nGd��GL�a��	�#!�+�D[EEԌ�>������A,u)�25�N������r��v����F_.����o�V����$�7�)DiOn�U���gT &�ٶ1���fE\uS����{f��.��󗔛u�λ�sٺ����oI�1��l�x,b\vJ鰺���h�E�:=�t�s^�a6]~�]�	��y#�1s�"oѻ�,QÆ�ֈ��/��Q�Bi���Xk3���f� kr�L�����%�����-�vU�J�vwP$¸�8��}	xw�M�Ow��T�;��I5p�����&�wbc���F�fWA��q0�����vb����ݙ��Vc�6��[�@W�֎�k{�4V�[]];������c0�x7z���F��ѕ	�ˮB "�o<|��x�ii�7\��_�!�(�M5�|����!�1�E���.�^`�UuZ���	�z���!�2>͋q��0܆���]G���Ĉ�:(r����V�or��
���{�:v���"�ř�v�T�;oP`���q7Z%igE��p-���V1SiX��I������[z�dDR�;��Ȋ���N�"y��֪���;�*����@��AY�S��C�n�������_CA)��`c#��՟Ot�{ׅ�/Qp
@ᠻO%�c+� �o����]oX�A�'Y��h���a����Iwl��<*�&hX��^�Z�9g�Wak��s����\�ca�Z�]�kF�q]��ܯ���;~G��3S`
�E�k�miE�7��Z��e���<ݬ��YL@m����%=�=�`�t�J��/�]�7��绝܋Ww`���1���)e���B�A9.֘�T�W�ь9�f�o��ĭ6�����VW��^��]�e#��R3�������W$7&,�7�c�
|Kk]刪
�N����#�A���X�]�Y|�5�Xlؾ�(֥�75�2��\���j�W�9��V���ܴ�B3w�B�=�:r��^��#�f!�
ƨk$v؄��\����2�9�KqJ��m=�v�;r)v�dY=j�V��)�i��yg�lux�I��Ǘ��5A�ڭ�r��J�\�ݯ����Ԭ�x�3U���P�K��h��)��n�$@��˼^�z����m��+��XҖX�����J�N�[�"�TW�mӹ2���K���eT܂�wkO1�@`Chb�_X����XN�g�{cw�[tj����uh(,�6�b�O�E�Y}�7-e��u�f�*�yw�u�1f`��#/�m�Y�	��Ԣ�r��}w}����m���:�w1����ΛX�=��������������l��ĸh��{���z[��Ɯ|�&�z�u	�z]��j��t.� ���k>��Ej���
���^�
�=uyV�rݔ�=�����9���^��:�5ݏ��.�V^�����_·�P�Ȃ �EUPb��mPDX1_��(UQX����*"+X���1X���F"��X��E"1((��֊"
,QE��Q��*"0TQX�b��.+X���F*�Qb�#(�TTA�QQX(��DQDDU�#����T��V2�Tul Z��Ld��PF,U""�*��[1UQX�Z"1TıQQQQY-����TQ��ձT�(�c�DF"�"�
��QTQQ�Q�UQ��b�IAb�Db(�"�AQE��1Q��UUV�ejPUF"��*��
(��QE�bF
�Rc����,E�((�+���ȹeUQQb,TRETUF# z" ���rsJ��E�OR6w������HA�ho<*�35����2��i,Gb[�M����N@�Z�nR�PP�������u�,�1>�J���
幘��*��mH�#�R�
ڹ������O� ��J�~d?t��:�Б�{�ޟs�<'��Q#t�S�;^
��7	J�Z�vm�@;n'�|=�ms%����~
�w[�U�;	�������.P#��G@�VRv����Ij�Ux���?���W)�i�;;�����_F7gD���:["�9��\��Q!��Q1�ѷ�b���d �QP|/q|'��O�_�?w���1�A2��[���f��LR����"�G�g�g�Eٮ�b��Y�*NK2���Tʆ:Y��p��"$�,��m�\.j�3���b�Q+�lR�9���Ɨ�������}ЪGDƩa���3ʄC���)����j*�H|*`�s��lT�N����3E_cO"����*q�OTo�X��
���,$v�B�Q�l��!����=�^�pw6nQ��'�v�_�=�}���a���>�P�r��/���pH�����e�T�Ng]�k�F]pN"�u��P�C!�ʮ�CV؍�eY�o�m`�^v��t�#�����*O�o���5
��}�M���`{_�@S�F���utwuu�[Wt���R3ָvL9�:���[	��ڧ�q.���uq?���Tn���uV���c'�I���ᭃm���@�H9V7OE�����:%M�n��O�sǶl���Ϻ+ؕ�R�H��Ї@lmOy�ұ}�p�e���>9���\��1_p��oY':�g=ʒ��~{]2C��qDɿV�.�����>f�s���s�\�V�k7#����`(>�+̦����[/ �����R�z�qU������+9Otwq3 �^<��q���i�R1�"�Aҋs��v��GD��XG:�<�]���0�Fq7& 	~��JV�����碐^9��������Sa�%��W��R	ޜSb�'^N�<��8ea�/�||865`�+'���=��ˡ�6�d��㨧��9/m�[�Տ#NԼ�n(Xl�"�?S��ܥ~4`W�)@eF��r﫣�Qo&��j����c�gYb���6����Ќ}́�R�YD�3�P�C��F׼xty7}y��R��N�o�]���a���܇~�F -3����O��lT���uX/'�v���^f�3M'��#D֯z���f��=�%�h!B�Zh�rn�-�EsiL�آ�-Ԍkqp%��~7\j��L^\GA��ד]�"�s�Cv�otY%S�F��(��=oQ�k#X%^&�͌	�ʪg7}��\���=~rԱ[�I�}�g$E�GFsss��@�>�*H�	�w0S�!��G\�5�Ɓqv)����q��1V��y.u7}���s�}5�
�%�7i1�(������{Xĥx��0#��(>�4d��7X.�Fe��4=��#1Xر�Ϩ�"�Ϋr�$f��LW�m�2F��!I�:���+2aOײ�� ���#t�X|��g�o�b�c��Ǩe��l���۰�q�ڤ�[E.�*��W�8#b�jj�̐=�n�}��%R���"߼�Z=B��9��܂4vC�����3���~e�ņ�_Bj����FF������}jm��1�������{;UBLX�eg�y��l��S�n��7�eŇT;'cG�V ���&���#>�abX*7�饺�O�f�YC»�\+�CǅO���z��y;�tZ�UCbz�v�^E��/=s��d�ˎ���Q����ӏT��\(P@��S��Ԯ�)�r:�d[�u�ɻ�}��g5֭Ek��9T�q�'Dq��0ER�Q�TX�l�<�?��VWpCm�4���#��c.fS��hr�}���h�yW������&=����]�S]�}C��3�w�f��5�b�1xX���t���K!���.�ˮ�:(Zi�"�J�4����1{�Ve'Z���ǲKY�#����G����+V�7�w=�_��X�j��I�>���'D"*�!�%�aA��{+,���֖�m���ɶ/
���E��8��j�	Ct�H�JBc� ��]$SdX�*�cn�#��/�W;Hl1���b�R��E<�����P�d�1�R�F'�ت��5�OK�W��V�S�Q�=}�o'M��
Rs)ż���2�ܸ�,�a�q)���*&������:tz���xjׯ�E�q�!F�:��xv��S,G�=��ՙA���M$�*�^�����C�l�%ߟ�_:y[N��S"\�"��w������As��MX��4���p�'�7��Rs�*�*�?yzF"�N=�����݊ �ޭ�F�v'��� �u&8G��9�ړS�
�a�v�曧�v�w��-���9跈���B����&z�$�ӛ5����Bk��4R&��a��`���Ǘ�\���N�Ԍɸ5< <�A��Qռ�+�X��5d����z���3�yw{�XU�=��6��c����j]�J��=׻m���v�r4L�z�S��n`�p킌Ivr�Գ�4{�dr��yr��A�}��Ӏ��5�n���ia��Bj�;R��W3�k]��9��uz����A��t��v�Hl,J�{��M�x��ڡ7:dL\�\���B2*�*�O��"�]gX�l�w��C
cD9��,__�=�=}ո�k��T \�b�
�Y�H�,�j�yx�]PKf�m�7mw5�з';�Kڥz۾���W��ەSQa
����U(7!9V6�OJ1�6���d��g$�]�Gt��͗{܎�
����G�Tv�"lu�p�{�]�{@�#]�}��V��өop0^׹N�=	�ƿc=��ˌ�
��#�B�G��s�5�Kz��t6�en�}�2�Ԟ�
�(�Md6��\�̫�j��ҧ2�r|����GV��(webx�@���$
�E�=FIs�s�; ��*���l������.P���Χ+&yN4o^w`\�]0<�?�T��%P��]<�ְدgeM�;��9˲qp[��cg�x�oˍ�*�lW�_�]�ud�)Q�8UyZ��K��m|�g"=���������p̑�u�ո��y��Q��~:��]) ,*������W�;���0VL*{ �}��#3� 0#]��T�.9�䄬tM�+�;�����h�Qw�o�ZB)7N��nKp+���,Y��b������\<�9V���WR�合�Wݎ�}QVͰa�oC�Ї+��0�|�n᣼�p�S�g:�l����vjwu�W�d���*�V�L��u��4fIh2.�L�D�lߍ�b����WL��=��cݼ�����5	M��7b��=WD��K��E׶���=�Ad˺*����ܾ��nw��:(�Ŏ=�%�Π�	�aХ�b��>��ѹ��k���{}"����d�H��t��c(@�*!��n<C�6OJ�u"hj�K����� �yFꋟ`|E�Y[X������v��zf=������)�]���l�'s+J�u��§/�V�u	C䨌ڨU�;�]t��ti�U5l��fT�l�w�rp�8�"s�6yJ��k�Hr!{d�BP"�:�|���.[��t���Q�1�I�u�B��%j2V��3[WʔI���U���ӽH�vkl��@�9ש
�!ӧE�p.%�s�6��Q��Ĕ�AsΙڗ�f:'q����>̕�I��䂍��
��:��N&���eV�FK�xvζg���5`1�_t^��n��j��A�\��hVVWn�q>Sa+��F'4B4�X��!Yb %�n[�[�,�d�UrAA���|v�$h�y������8/|��y�}�Y#%l��$c��{d�����r�U�ܳ���;H܈�-��J)�v�~�v�	��x��n��w2wvL�=���]j�C�ub���K�t�(Ѷ�)1�.t;�h&tl\�F��S_�o�y�w]��X
��yV>�����1�J��X�� =�	�,^�N�qZ⺲�]BK/F�W**8���_�d`�j�M�R3إ e�[��C���y��A��G}6=�Ȣ�\{"��FU��QvS���N��wH�Լ����u+F�!匘��ƘF�S������t��	P\��0�fb�WN$u�Aj+�^h4�7Y����QC���'���ӊs�sg�p!@��%��P�J�:L��1�WDb�J��k4޾]� 虀��l��V���#1Xر�ϫ$!iL>�ݢ�gָ���Չd<�9�d����ɢ�j�I�DTS�[R}R2
����F��v;=�c�84;k�rd�iq6��S;/jwv����Ő�ؘP~�P��u������Ebu� ��z�Ջ:4�b������L:�1s����b�|��hh�226g}�W���# �SnkvU��]kC�]p�ų�jQ�Уx�yලxA�zj :ǡ��۠�׋���3�eL�t�b���zw�b�Y^����]�Y��횈��ټ�=�����u{t�|3e/��u��rA����z������=�r�>��n��C�C���1ĝQ�{��^=HG^S�n��082ˇ3[����=~���2���ʴ��C��Wۭ�dt�ʡb�=�"���*�җ�P/�NÂ�F)�T6'�7D���4Ɂ��7H�z�Ψ��B�(vPVhǪga.(>Qjs�ԫ�P�'�I�=�uI^u���G�֟���Y,eiخ���(y3*\H��8�&TyeE�l�<�����H���5����[,9����L7,�&��L^�R�sJ����������[;Q���J�>۝K,i�ć	J�g��>�dq���(!�s;�~�&:rH��a�}���f�`lQ{s���b:��k#��#`��(�dS����ڡy.x�T�Bq]/����u,��t��=��#�M_69g�� R��ׄ��N�1�̸�d��3�1ԗZb8�>�.�,�υ!^ԍ�����G�M��?�VV*Q�3R�'j.�L���1)�D��v弼�u�9C�4+wS�#<R5p����W����l�NV/CN�5]H��3�LQV-x:ܮeMAr#�ƅ�Ez~��N�؋k��F�H���Z���_��Ӂ&�o���5�q��sr��1������Qi
Ø��mm�YV�jR�$|��c-��GԢLZ�+|��;��΂s�Oc��eH�	]�o\ξqԂp��g�K��ܲ�bqM��sޠ�R��ûm����m�Y��C��ȷd�"��ȱ�ʂ�t!kPY3_�Cke�ѽ��/v�}=�G�{����ҽ੣�6��}�hا�B��h�M��ST2��亻���\��F��s	����$�zsf��W3����:��/U�:晾ԫ{d(u<dr���L@9.����+y�i���6f�V�ʛ���8��X�z���Wh�}|�J���F�y«�B2�T9Vi�J�rޑ�v=�m�َ����e��Ѽ��7��AY��������:�*�lQA��Rεcu���z*��On_.[uq�6w�:q�t	��w�0|�#��Wd��V�sc*�\�J�64��ɬ�g�]�R�����F4�,����
����H�0L�!��@B'���osC��5�p�R=�a񠣯k˧P���%9��1��XS��
@�-�A�h��Fi��~R2�-����R����M�ڐ��5��'~Ds;2���j�"s�{3��c�ސ��ڰ�a8�P��)���h���b��>�S��AQJ�h�5�
.5,���4�����f/G:�Зy�������]�[�(zL8�ڶ�:Ac��⴬ɽ����53蹺}�������fI�e�����U'�_Q�ک��Vw��qY�n%^r��_�@sq�h��M�w
��.u�\��{�g�}cY9Rj ��/=����=}�;�X�R��묻�����.Vu��*U:y�a�^;�P�-���bƼ[>��9�����:���U!���H�D	ɷ�/��m|���x�egP�wc�ZW71W/�h8J@�b�Ӭ���̎_��Z���1|py�<�������Dg׸^���IaVܻB"��n�	2"p���RZ��L�}3[6�4��&��nv�,ڨ~�T��P��v��0*�z�"�l�&Z�58�T�˒�u�h���r��M��3� 1Sy7咜�E� ��w�B�Q�{dLT�!UCYE��3��Yx}7ӡ_�:�o�\o3ش;��a�] f:B4Eܨ�|�ǭ�V��o��7Z�mw-�ovX��(�7[1���j�mm��k`�d(ᆀ̔��E���S���[��o�r?&R��cY^�Z��c꾚��>��YȰث٘�z�VVU\c�������Ǥ�#8�l].���e��w�W��p���0��{k���k���Td�����ᝁm#6y@���Ύ,��̾�\Mv�֙�t�tV^G�-�� j�Ʋ��e��X#kg|���F!��wc�
ʣ0���I����CM���l�q�K��B���Ո���A:�fn���`gf��'8+\��S���5��W=�O[�:���㽉�m
�>���7�u����`�#h'Թ�����oj\�H" �)h����-���]=�S��On�|�z���Ώ]
Y@Lb*� ����z!�u�/JO�wx��Z���J�^�G�<��YiV,�V��Z�fT��Kr��۽���;��N�5t�� K:)D�<X��B�+ �� �����V�4�Ǽ ����J��Y�H7hu��tf�U�{�)SKvx'@�r��WN� g����b��i���+�h-iEӗ?-��=Z�qMȺ�O`�D��X�����(ʔ�K���r�T�z@@Qc��luYyU֘<�����'z����!t��{j���Y%;����wW�s�y�z݂p���l���
�c��a�bN����V��+(��}G/�����i���8LcA��(k|w��e�{'	�Kp
X����yDy�C�)��)��d�����#{/;\q����|�O��W��%q�QO��Y�J{{�E�dA�D��}X�c�e`:L�M1��qW,w�[�\��-J��e��=��z��QF��h���Ŕ�L��{BL�Jóts�(#5�ރy�����������[n*��N�8mĀ-��|�:�qS��G�+:�/Y%ܟt�ʾ��]el+#��޽b8�K����+|�`r�ڷ�9$m��7�{ z���w]�
B�O��V¦j��pj�R��K�P�/�[8rt��p�i���|U��c���t��]�:N�<��Ԣ�f�>!T�z$�A�V�����(�Q���7jӉf�~f2;��_�N̘O{����ޥ�ˬ��E�@c����a��p˳�e�;Gx�[�J�,>z2�yиX�F�1�z��G@��ˬ�R2K�zRJ�n��8:dX�Bn��{���5��l�������W�|�!y1�Ν�(����u��J##Ǭ��e����WC֮���v�� *:�Jr�"p��	���+-��%�X�3���3(�u���9���]�5�фU�MƉYb�R�M�WR�R��q�t�p���Zm�u�NC8"bk�iUk���wmS��
}M�\��7�m�k��[}����4�h
�oAcY��m嘺vcb�����^r�vw��e�� ��x��t�ӽ�k���	}�X�p�ke�s��5�RD�W����w��G'*p���Օm�o�
]��٩Ջiᖗl����ih��(�CX�.���o[���%���5UF1VDb��	�k ��UW-T���
*���6X�YQU*+��dTA��T�QTR(1U`��EF
�J��*(�
(*
(����QX���e�kQF)UTb��,`�TJʋDUAQ����b�"��X"��*�)[j���(��X6ы+rت��(�b*���QQQQ�*������b����P�F" �b�ZQE��[�R���H�Qb�-1���[-����%b�Ę�V#EAE��AJ�҈�F2-�AAH��eAVA�V �LLU�V)UX�Ae�Db�+R�Qj,��j,kb��Z6��QAA���
Z�mj�[amUDƠ�-�V��j�ZP�Z�D,��5�F�k��Ģ�����Tj(��"#o®�D�G���{���)��NF{��P=�*T�{�4����g_�y�8\�f����p(j�{�x�k�֝}�%[JҔ�9�vݟ�L�v���^
���Fu^N򤦠=���9
�=�u�cE�wыV���n���{M���o&��Bt����:�y�˄�%l���+Y��S��� �/˽4�Κ=�U��=�t��>�[@�.4����jF�5�s ��Qnq�;R�j,hD�������������H9�*&�R0��d�ׁ;
�[3�W����֒��Y���yړb�����@�l�,^���PO�ul(�딘ݗ'�
�Q����Z\�b�!d����WySx���m�DW���!1�J�LR6�|��¤��6^&�D��lN��|�^d�
�;t`t9v}�6F"�<*���2�z�
tH�=>n��Čs~ʈub����| f�.�#��}b�܆��i�4���B�M쮓"3�bB�i�s|\�ńK�`����*�S��*n:Cv���!�H�~��s��br�U������>�&譅Q�j/gF:���
 a-͎�F�{��Qju��t��ٓ+�r]���E	�5)f�1�ю+��^�`]�\���y�e{�,1�#hf��1u�G�yE�"���P�\���u�#���V�:!���e=��{�	dY
Hi+d�W��;s^��7-�5͛5� ^ˎ��y���4��Sv^t�ƥ� !J��K܆�f#e�J�/���Z����S�ԴV����~�J�s$Y�U���>�ɢ�(}QA譩>�Ud;�Q�t�r�滯Rx�rQgCZ��{�Lp�IWB�\��PZ�s'φ���JQX�m����ō�s$����wp��Z#lm%1nq�]�'��r�}��~�l	�>kҶ��6�)�
�sҟ�v�Pgx�P��|���\���ٸ�8�y�����=R�R�2V��cjS:��,��	�>`OP�@�,�s[֪��J^�@�	�p]a��1�B�Rh���%I����X�����oB�4;���ji\��J��e��Q��{+W-��y����ʰ����&dh�b��h�����&�:�.`�U���}��S�����>�-�.����r�
�}קmX���+��x�޺�}�ƜJ��v_r{
ޙV��[qC=�*��'$5ssgÆߐ�e�({�pWg�O7�Y/ޥ�	�ƣ��	-���d����Z3�C�X�`T�AR�(,�Y��o�az��ȯ�u�����ͭg���b.�Ylu �P�/p��9o�	��VT;�t���6�@G��:W�����=���$3��?Gs8q;;�Y\̼����"�2��T�w�;۴��fޭ�����$;�C�u\-g�2��e���~�VuAp�]Mn���w)$��:���k-]>:���΍���&� ���� �V��o����e����J��9��b�+���:Uc/�dS5�"dJ]�v�Y6��Pia�!�����_o�y�sҔ�']�7ȑ�QW�\��'sS�UM�25�A(|�������ʯ���+�v��x�[ii{��w�9��w.S���2�|�������f���U���(n��9�t���z�ʠxn���hV^���&Vn׳N^�e��W������Iud1�/�5;�߫)\n�bnu%Mm��)^�d�����������E�{իC��Y3�����f�z�?+q�0v�z!�x`�;,r�7}n�{WtP�ˋ<9Y��C^太7��-w@��`�֞�O{H�|U:�n!p�����^��Bȏg�f-��� �A��C�ݢ�8!�R�tg%u��ש��z Vx���Tt�g�wj��Wm4{��y|d�ɸ{�'���M��LJ;'x7�A�\�u���S��v�mU@SQ�i���򷞰Yƒ�K�=��t6;``���.��n.�i�3G69�\nu�������N8��V��aOE-������sj��m���m@"_��Q�,�g�V��o�H��Dc�Ku�UW��^�K��A�7ׇ��ϭu�-#����\V��B�"�9Д�r�}�;x�^+��cqԔPo΂jGV*�z�����.�z�;��-f���o��F��n�8��A�'�P0�����;n�v6�^�
��3O_--��z�F|!��	 R*P��H�s��u�V���*ɖ3��U��)�˂p�Y�Qs^h2D��DOL�/���S��rW�ԧ��P(�9M��(ZP��M7�'�A�U�}]bex�u�43,��4�� *8��v�s��#��n�:�gC�~�w{F��b��ŗ��ώ���U}F�ٺ�=� d� -~��B���	�P:L��܋��kySP�c������wex���N��S��'c���]կt�۫G[Χj+y�;�����|9�;���yWoM�HVu�--o�Y�֠�^�rz����,���d�Ӿ�����æ�0��uv���0��Gz�S�t�r��5�g��3��Kbj��٧�1�zC�f��94������n����3���Yf�ϬK���^��7����{�@+��r6K�]J���Bct�:�a�s9Lopg��>ջ��:�G%Ҟ�s���C��ji,w+.;R7E�kb��O�;a�ciq�>M�n�;{'oܔ<m)�����'�ff��4�]4�;b5�-#�������N8����f��ܞ��9��u���l0;c����	��yQ揬�VK֚W�3&�Y��vN�-��ݯ`�m�ʥ0��y�^hU9�%�}���>��8/&�t��3����1���Ů�tZFA���΂��5]Bq�4�M<�޲ ���D�����)��q<Jq��ʷC�=X
����ṥ��Ä�<d�T�H=A���{P˻�a����ܗ��R����F��<Y�fy����
���w%7f�;�#&��5������<wV�1o��PkB(��gV������wm6˲��%��ucm<�)@��8]�`�e��	����i{�����2���3ˌ&^�u`��	����#����؏���f��j�C��h�g�FtSv�Uy4��+d��:f��c�O�lTގ�:5�5���zۚ�ҫ%��]]��c�,e�f.�[}'��j������*���D��W�.�l�9H4�)y����?zF�-�s������v��-\S�^z6js
��^�Y�T٪ᮻ�7y���O�j���l+崵�/NMkW����M�On�D񞚪[KM�X�y���lYė�zB���c7��N��%�ם��B'����6�Gkv�,VR7;E!�l�E��C���mt��/�Zp�T�E�ɽ�Zy��E�H"v�N�q�
+i=b���@o��;��bk����h��8���u"42+r#�;�E�0�Q��-�^N�08,�w܋�y��[,ڦUwח�}�ú��2����sp�el;ܧ�y�]�	O�83��# �k[�]��[K��M�yK�K�k5���|�j^�;g�Q�v�v+��j�|Rj��vn�o=u�@s�kQ���u��k�M[q�+���9d�R؎W��sJn�Ny�y��i��'�w�û���q��ٗ`)�b�4*�����͛���7�[�s�O\^^;/U���>��{�}r}i�?$�ևlK�	�R�,�޷^��T�v�Gk#7[��k~����ɴ�F���*�ޒ�ڭKa@yp�h�R:�ցYR#1�~*n��z��2���M�����u�]�_��)��ُ�h���=uRf̞=iZw�y-�no�";l1A4/*�q8Vz�*ۚ:UT]�KMb����ږ�ү����p-ï&�>�������Њ���Yn�W����¸<scX������S����6uab��:{]E��j*p�*���JD��1�`�R��bZIɂՊ��[��"�ےn�Vz�ݦy���A����� ��Z��S2�5��>`o9�-C�)WX�wɇ{�p�we�\k�\ޘ��-��c�z0g�L�� �g��Át<���~�Y�l��e�w�W���������4Wo*��~n�ٖ����e�b��h-kӓM;1�bh-ҩj���K���}q�@Nas��-a�C42��"���7��+DF7�7f��Ӗ�[G&��褅��S�wK��W�-#h�s��������&]�O;-&�ň|��/kޭ[A���C�(>@��nt*QP]ݝc9��}�Ӧ�9�Ŋ{g������2Eη�}�/`�ܣIt��YX��g�����v�Y�V,v�J��=��#G^�T�A��ѽ*ܐ�������M8�_��>�;���>��ܾ򞍺̄�:��*�*\_��c���Ōb[��שּׂW�q�M#�ac�&b���yOL�Qeݼ���5��:���;�{^��Hڎ���VV�W1�%M��n���n�籚��$�f�����!���"D=D`��t�v0�Ɲ���t�y�#q�2|� |5!}�bT�j�=��"�:x&/n]%�}�m���=�M �Ц!҈�1 4n.yQs��v�S��s���k��Q]���㮩�v87�D�
��)�z�Uvf����|��2������NM�R`�8�.�C�����*���+Sx��a#�g�H"��BP�D��!�8������E�n�%t�[�uܭ.|2��2�ɣ���i���R!y5��v��Y����U���F�y��t�ô}��7���7^Ma���h2xL�d�U�3#��������XV|K[�؇���
�7�Ny�����#emm�Q�����˲.^p���k��roE��t��(g[b��u�+�f���>;N���y�~�f��W�ç�~���yԵ{��QرS�"��7����Z�y�T����⸬�}{4^\W���3S�U�U� �W6fknd�g��K���*zբ���{_O[ޅ`�6F�aV��%P"v�n��<J�eưu8�#Z�l�\�f��J{����6%���xIG�}��O	�����"eo��{K��>	��Ζ7s�4�aq޽U��*�R�5�`w��:�u��^����;[H ~[����T�x]�S;��VĈ�$�.�/{s����{���ˋ�kJl�#��t�ߚO������s�޴{6�A<��	W����oJ��T/�9�Z�q|�.� ��]�;+y\(��*��S�Q}�w��}X�.���ys7�*
C��׼촮=������߅:�{>h�ĉz�9�x׭�)v�ye�a�B8����e�p�A
��T�H��T�wm�k�jx�2k�<��Β?�B{����J�kn1����>���9���\U�+5"p�}Wߕ)����V
�kg��D��Rkv+��zk��ʁ�t��DbgR������v�C�;ޭ�Q���rsF�}�9���b���h�X�����W{��e�����E�����E�y ���&����nh*�Sdo^u�7s;��Z��
yS>��3g�A4p�-EM�)��3-�������xhBg�=����צ�Y��t���vi��F�zs
�V?yE^$隕aV���dͰ�-�5P]r�_����h`Hǵ��kLѧV�l*r�U���A��X����p:��4�mhĶ�����N��[\���ŧ�.w���=BT�9okTh'6��g/��"4�V�Ti�;�;j]�ѭ�A�t]���L�67��{��$��(�\�4�N޹���
n�y�F=���4Hb�q_P�T���k��U�TZ�* ��lu�,=]]��4>��v��{����w^*�>���bQ����=�Dr����c����J�c��N�&U��a��6���MV�w7pX�w��Ϋ�[v�%� �dj�K���\�#u��������M��h��o�v���2l��}��0�-^�7���H�*Q��8�a.���L���]e�5�	������7ǁ�p�~]k5V�lA�a;�W��s�^�qE{�19���{^�:x���1q�W��mv�W0\Pe�ﶛ�%�c�6a�7���}���=��OXGd�yW�f��m�W޹�u� �C������u��
Y[c[�z�|�y|*K��[�b��Q�}� ئ���t�rkn	.K�i`{>MK�)ASx=�g�]{;i찞j�Q1��)�f�M[�����Y���>̅Ȃ▓��w�-=`�s�dAs9}��'k�-��
�#��v���6�r)_}֞yqG�zir���8�1t�{7d�Evx!\=���kf$ȑ\,���e�,ٟv��ͼLm*Ls������}1�F��?95뎎)�آ&��f��nķK��cv������ڹ��*�*w\�t�;Ɛ�\՘+gM�[��cy*�K;�^tZ�����OTk�ğgp�O�p���9� B�;*�vB�^+	�N�_2�m��֞�y�������`0z��l^S�Z��u���'�J{�I�q��8(�����`�J���-������"Y��yu�h�fn����+�����,@Y�u�"�
zK�fM	�����NBn��"���2�l����T��}�jL(J�:p�[�@��X7}��=�t�bp(%�W�wf���VWwp�P�vqY�H]����:�v&�]��sE5l+�O�Wi�L�u��������+�w:	���ۊ����N��@�i*ާ��:i�	l^�Yx���xA��e����A�c(���b�)��pj�P��r�<P£ꗂ��mrع�us����b#���=\p��Lz�3������z��9��:��FFAݔr9Z��d1�b�ui�a�ٴ�!��o��]�{�ݭ����ː+_���������մW�c�N��^ݘnOgj��C�z��<�Κk�O��-d)Ow/r�<A����[µY��[]׵a��H��`��eã�ݱm�.n���a��}�&ޚP��o'�%Y���Ah|�~�����_k﷯��X�D�`���l���,E�*9j���5*��)Z�֡XZ+A�mm`�m�[X���J�P��6ԫl,����AF(�*�Vڍm@��"¥U�%�#
�J�AEYZ��B�EJ��Z\B�[�%QE��K����bԨ6�ʕ��YP��*�sm
�1�cV֍-j*�����mE-�2Ҫ�Z)h�h�[
���Ԩ��U�KJڶ-�QB�*+J����e+U&8�lQT�%��`�D��ťlZ���,�"��QX*��*��U(�TPEb*,AEKm�V)YU��XT����k�1�j
�[j�(5�U-ʪ�X#��b1[q(��c[�Jʊ��*���eZ�m���-��֋mh6¨R�A�Dh�V!Y+*�+YV()Z4-E[lVҎP�)�kF��߽��g�y�2E`��:��Է�c��@3��c��lw3�\����9R�7��d���z��kx5y��=M�#neu�����k��B�]��r�kXl=��!����|��>hgkwrℨ��&�<֏_)�`}r��c���*x�vj��0�^�����´6�ZMR��`m�|�u�υΖ�n ��vl����adl�^�7�-+���J(;��\l��u�.t�����jo
J�Pl�r�I�̏?Nd滛qEU�ힿ6����GZګ�Y}^)5��N�2.��i��1.�L=�5|ڷa�d�S�A8L����'����.J�ug޴{���ꥺ9����}r۩|�b��4%�2-	2/�DF�͘Y����I���l�V�v_qOa��O�# ��I�q��M.��]y���k�􊮯	h��G7`�es���6rx�<Q�Tb�^;/4��fD��BCJ�qU��pe#�˲�ڤd��}F��3n+z�4�P^�x���!���՜[I�� �}C0�IW-+r�q��B�*Z�P39��K�!^��*i�Bq�u�t����f�*I�Wz1TVn��e%x1�C�-�U�jׯ�{�.u����oh�w��gUN�Rj��fB�����Ck�^�!C�j�#TN��Rq�Ѵ��ݷ�6!�J��6��a �C��E�h8�Q���_aG����S�f ^��;�oT�9e?vu�0�=Ma�-EMy��5��h�	���ܢb��o9)f���Tr�>Յ�Jy�u햢��$�d[������'aV�����/��U�۳)�m!�[�V�gC�٥
""{je�IQ6�:���b�F=Q����<[˕E|�՟"��{|ߠ�H�5 ���fN[��٢l6�1�NnV��h�0���B�Ю����Z��כvu�=�Nvny����ފV/K`ᝫv+�c8♝���72�ͻz盨|���j���˜�X��Xo����ʇb��F�z�|�,;��=�`g� ���=�:�gJå���J�=�]���n ��ϖ�=�<	lE���-��=�-�t��=hϦ_/y�ePL,S����w^��u��.%/�ؑ�3�2W|_�Y����w�z�'�g�<�����G/�+=:�R�Ԑ����ךּy]}HW��\�b��B��P<�KU�/��;��㏱������@�x�cv��jWn��GP����YZ��m4���"_��'�'�����ݍ{����l�f�*ܸ�c��U�Nt5C�w��v�\��\ȱ|�RZ�e�Y���rO�3@�J+����H�8���������t`���|�]�m��_)�Xl��F�p+҆�VPsM���n��y���6��6����F�9ЋMT>�{)��t].�G�<B�R�����R{] � �t}���݆�&�"!���g�3E�u�<�s�[ �<9�5��*�Mʢ2�>����&��Fv:�I��W��^�+ ���2�����;��U����9Hg�z�x�n�	�<{�~�|SY�MW�f����F�8�~�uv���앑�u�/�j��u6&���o�=�ڦ\�����c��=��K�i��
�;`fT�Jqx��nM���<�D�
�qr�
�΁��Xe���UmU�Qܔ���Ӏ�����u�=g���ꏫ����V��{uu6�t���lA�H�tI.�B�{{����]3�ˍ��hu������}{4Cˊl^���N�S��`��a���w�_c�Lup�An^�~E�oV�㳯6V/z�eO
�*�*�;�DLS�"�h�I�j݆[>s����J{з{��r�'�T�9/-��]�XG����l�� Pi_����i�Z��q���]�&��Ic;�������^�B�H�������t���TN	��h�n�&���m���/%ߔ�W��(;�q��4}eo/3�;��L�%��y�c����������2�K���
�Ъs�KE�;¤��Ĝ-���xqun��/������H�-���{mEwn�s�Oh�0�>c6�;�1=ݥK[����6pZy �Q�*oK�9XV��cڹ�}�@݀�H�q1���)`r�ܸ�N�ë�w(���Cܛ��5}v$g	gfĲ��s!˷u3��w����0�ca��S������4A��ʲ�1CS%�W��x��S�8n'\զ�NC��toc�u���������Xګv�!~���SU@n��x;���kҎ�͵��C'�V��ѽ�g�9��4p���9�M�qP�c�\Ej�u��N�[P�!�4�d���ړ�m�*��mf5Hm�q���\wy16�c�4�כ�CQE}����2{�Ru�>˒���R�m�����ܪ���Cح��>{]��;4@j���l��!�mqIu�:��e]�iM�����{����A�ŏ��94�W�^�^��������r���U��0����ԭ�'�{�¥��Eu�S�s�����c�^T��N��[�+)s�C����|�o;
��lO�{�rs���΃�����V�`�֏�v�(4�m'��dv�ص�c-G��hԒ7�]�s����@UX��+���[1SO��b��	^h���x�y��Gpm[�9�~S�I�p4vN1⫑��U���ͺ�z\i#��5<���]���$�\�S��c�����GT�/�>W��O���%�8�wG���f��f�����v��Dt���4�j�Y���P�	c��=2���\#��/U���\>�)���ͯp�㇯c�u���9"�c-=�5��I�����n�#��}`����_��c�f]�)衋�%#�{;�uj�v�"��O���l�Vw[����V����Z�Me��S���1�����]B[$�G�q�t�+���ʮ��]9A�����{�����(����:N"�+�c/yf��no��V���m���Ci�I�*�Fk-X����8�ǯqE�'��zo���}�������6�4�{`�&�ƼYj�^r��#j��W���ɗ��v�z)��Ma�!��hD���d1���u���\I<����~�t.�����Յ��P��V7�%�3jE��'2���ں�-n�w�:hNaW�V�]�7M�� ����<�~己�2�Y�a���%wy�l����.��'0����]!��Ы���'�<�'I碧�84�b��rVۅ�͍\��|PT�5'�9Q������e� ��,��|����O�jC|A�x����Jeؽ���R�cMt}�e����kl]�Ѻ�ƇQ7�QCJmu�'��.�}Búa��vm��6V�6�D��ٸ��h��b��jwK�YH��h�0m.�.g�N�6�-u��ڊ�[q�y���=��+�����[��N�LwK���[�<�]u��r9Lodcl�Z�l��:ҍ���E;��ة�Jn$v�"��fp��hS��[kiw@��%~t����z;��:{�cW׻csI�]��t,]4�v�zy�-#t�_�� j�ڜv>+Q��L�(���Ӌ9���ݍ��R:��t%(�y�ej�q��iV��TE��j�������{���#*ܸ�~T�W�:���n>վ~�g.�,�}hr�Şw˗Y��7���΋LȔ� oμ�D
'݉pw���Rg"5�;�)�E-~щ��Y\H�;��I��CQFZ��4�=�B��;�Woy���4wH��e�M%��=�ӱ2������jz��8�Q�9Z޵y���xP�ҽS/F�v�Sb]�v�������p���j�M�:���i��Q��r�C�DS���CϷ4&b0wG^oJ�­��@c9K�겵8�,�J��U�����q��Gxw܎G�o Ν#�N�|3��ot����+z%��Rh2!�3=���;eY֚�='Ex<�v�O��aYTmMʣ���v,%j9�&��������Bj���� �EPhk N�;yD�Ӟ�!�8h�E�Q���1W���B�Xm�٦�>��t��~���R$�uV��\mf��A0�
˶���������\
����e��O��{Ռ�ŉ�L��/0�/R�^�ϓ��|��(U�[$e據k7͹�z�/".v�lq�#Z�l�\�f�%Ҹx�2+��.)���ëz���N4g=�9��A�{�1���M�Xm�<�y�Ŝ7#ޒ.w���>�v)�دN�ZZ.�{K�)vK���Y[׸��H�`v�qm[�/%��ձ���сߧ��f�dgTEH8�m�H��X-dF����C�����s�XGh�82�ѧNb���wNj4(9���'�|�^�C�Ɂg���p��b���8Il剏;���}de�-�^�����~�6�ޘ���w�A*%X�,<�í���ˣ͖�_��w��w��%�����<�8���ٗj\P{!�`��8��t�ӎ��+��z�e����[E����W;�H�-���8@�"�o"�f'1�u��~�t't������`�f^_Xl��E�u�8LM^Of�vk{
<1�h� �&1�+p:dr�e;g8���w�¼v6�����;�}K��V(9\�����gE7m�l:�)B÷mZ��ڋ�������(k�Ҥ�zۚ:Uv3]+o�,:a�˩�[��=;�lW���M	o��54�����v^S�&�1'E݅�1i>������b���iC���m��E��|"�=)�B=n�7���5��N�zحwn�齰6���A�-���/NMhj��񓡬��dA΋1���o��@��A�]!�cb�^�h�!=[�3.z��)�%��s�l��7���+�ἀ��qJ��SC,�%贺��3K7Ǽ�²CW�V�z��� Ky�m�̕`�g�t�W��k9��]:���z�v�\lՃ�\�eg�戀5��=�ܱ�]��Rt[;�(8�4��k���Y�I��aj����|��eB���ڷ9+|.v�hq�:�u2�˾c;�]n��6&�w>kw�8�����E;��8D�X3�\�A�qp�c�]�\1>�Mh<|�d9�ŞS�=m��aqT;�X�:�ތ��iqF��=��ďKV'����Y�q�v�U�=	�{#G��TeӋ�{Qu}y��JI���S��O�G!�u����m�w�=�fb\�i���vd�����cjpm-�x��e곺ݗ�B{�}rV����;�]B�s�j�[{��q��^�DUt7C�vn��*�;ͽn!�iQޮ+;7^r��W�r�3"R���CJ�qU��F���f�k�*�b^\b��M���a"�C���%8�Q����!֩R6�,�-�n���R�|�E�7���&���H��X��A�Q���V�
xK�GM�r�v eH�:I69��J�3�ۖ�K�'u��srѨNM-����rG��r;bҡ����r���=�M�VL�#sV�M:h�_;9�q?Y��s��e�6�Npμ��`�v]$�C�%�ݻ]��qE�䠌�{��*N�k�+C�k�&K�`��YN�O��FF�g:n$tT�H
v�8rsǢ����r�og)�Y'u=�q�"h����A�:gM/-���vct{6��=r,�0�h���Ϲ��,/6o	�v˼6��a�6/=��I���ǩ�un@�2��AeX����.ή��:̢��hX�ܸ���;%dX}y����*&`�M`�� �`7ЦF��I��B6E�YAt�龡���S��I�=o
�u^>��q��/���%k�]�;	C�B=(�>�˺Xh+"���R�Z�iA�$ov�Tch�J���n�X�T�p�I�F��1uD��'-q��|�32Jߤ[��wٻ�m�h�47�������=f��vT�J�#�G*�U��VnM}�k�=0 #�4�X@v��d�tIt�Jv����� w���<���gW�s2�w3�FaB��C$��V8�XuZ�:�,ݬ'�t֗�v�6|�#8�m��bj �ƫ����K,��O&}z��&��˓<�{$�[#��Փ{҃�U��i�e]�p�FX�o
��Z{Ji)��=�k|K�z��	��ځ�0��l�/aw6�ZA��'qz�v���tTy5��x�gT��F�R���¥�Ԯ }�ҧ��{�+��;�臆8�����|�̣{f1�[��uo��Yҍ���W�AC)�TAaד��V��.���f�j�O??�`]��EX�{���#��]��t�v{w�F�����kw��pO��oo',�%)��!d\L�"9�m�����w��Rݘ��ݪ��MJY�<�KoV��u9�3z��ܿ��6���K�J�wsGR?/��mcR�+vn�W'E���(gU��w�� U�`ݺJRf�Հ�c�	zf����J�
	g"k\�l����B��͝�J�@a��a샴�=��M�}pf���QM����_f@W]t�Y�����#���J@-�Z�����N�:��-I��I�+4G区�{Q�Ե9�\�oMx�#�;l�����r���	7�8*�)\c[�Ol�Er/������gv�ūb���YPr(-|�P����NoIKŻC��`�8dm`*�������P��+�>�w�AhE��S��\��9Z�|S��Y���.��a"�ږ� i�eWe,us���o�Y�9�b��M.Ә̴�J����YR��#����8:�3������ϣ��c�U>�1�垮-������F��V规g5��M��S�뎡!��[/�ʼt���z��Xj��K�"C-k3z��q���tN�.l ۭ[9�Μg��*�4@ }T@P�*[J�ъVZ��jR����h�[h[Q�U�[J��*���ԶȢ5����Q�����m�U��9iUkZ�J�Q�E�h�H�h���P�S,Z�(X�maR���k`�mE�Udm����V�ʃe��ň�*�����j�QU�jUbT+ZԱ��F�m��+,��Um
��L��a*T�DU�f(奰Z�EQ�ZPQTYKbڴZ¶��@��m�Ej(�ũXV�Jڢ
6�R���2f*6֍cF�R�kJ��T�U�ʭQ����)keR���1����0�F8Qj�X�**�Ab����YT*��-�A�TP�«q�m
�,PX����,QV*0TQ`�VE*ւ�(��5�ڌĹTV,��,��5(T�Am�
5�l�((��XVfTU1)m�mJ(��XEkB���$m%�m��TU[i�h��4*��>�)�a�/V�\�T�w���N�Y�c&1js�W��S,����Z yF)��蒜ڷ|���,�OI�"��{������&?V��8�#z)�:Ma�>j*h�UbK���=}�7��O�R�������6����XX��7�Հ7�"f�.R�S���c��N���uy����	j�U��a齱���lX�0.A�9Ykm�<�t��{4|���6��:hNaWYT[��0�hMv��9z�]L|�曜���2�P�W��z��JЎc��k�8w��OK�ج{��w5���}h&Й�U��s�q���z)X�-��v��͘W�N��5�S��}�|�{��v�i�jۦ�9�Ŋ{g���S���\�VOQ|��)6/��>�݌UX�/x��x���\u�4���c��V�f`׳uV�{��C��*��By
�r�v��C��N9�O���LV��ۙ���n1��U�蠶����8%y�,�UX�;T��s�n��N���ֽ��Z'#u�(Q�&.P}����Xm�/i7qw�Mx�+����<�Jŧ�<Dv��C�ڋn.1�&C�+�7P��ʎ�[�+^*{c�n�:Y�H�pR!rޛ��ٺL�S���p�u�Ӊo[���E�ܦ�$�3������]�<��4c򠽪�:�-چ� k.��Gg���,�e���=���P��)F��ҰP늪���b��:r�9:��#sH������ĉN������A�
���#Qw9�]Sڍ;:��=�=�G:6��Ά]�4L���i��qQ��]eg�d�73��Dh�SYjF`-I�U��#z)��u4�Wr�w�W
�T�e��Z�,k���H2edMm��^P�R]*̦�vAo/f\\��-+�ږ�[��5�ݒ�T��A��7m��k�u�a�]RaA�pBȥJ��zl?��7���Xl=;4|��y���æ��u�sm5S<����z��w&hÍ
�]�����f��٢\6�|���sg��Y��LV����qYz����f����h��;z�)K�O`av�;q�D��CK��XL�Zzشm�;�?Owr�u�����jr��%�t��;�m9u�4�yjL��Z7W��7+�����
ehwm��Փ�@Ͳ�{ٽ}�Ũ�����ޔ�]a�K�XG'R��䖢�dYRN�^$�[�#���f2���3�[�[.s�v�c��][�^v�sq�n���5�t�����
�av�֍�QA�ciq��#��̝}� ;}��r��N�!~��3S��k�U�ء:�iM�1y��\�l�ὴ1��M�<q(��ջr�]�=����'�[j�b��w9ZP�ԏqc�.�����=���[u+�C�{PCB�3z����j�t�,\�s�ݑ��
�~;����Z��m# ��<a����]=ySٍsQ��#���NqV���U���^_Xl���8�FQ=}�n����N(Ñ6�:A�F7����9z9q1�]�\���|���w�k^�iq�a�bv����5����s@�G�*)g])6�w��&�y'{^i}��\�A�C^��<p�>���T���(�ϩR��d��l�XZѷ\���0��bfNɮ�3g��7Q���>-�t��&��@�283�J�q����t�!�Qh��**;d����*	�*w�]��ٮ��}��Sɽ^�낼,�J�C���/�mֆ�O���f0�u�(t����g���CY��y�=�����fi��&󛒚������!Y�ش�������h��)�����DGH�7�/���%�v+6���t���B�'�ӓ�~�̱��n^���~��\vh�\*ro�YE�ۤ0�b����o�_���7�/�51|��sd�!��r��8gj����;@�8�lWs<OG���:���7�����ϼh��իh<5o��!�3$�x�=y���u=����#�Sl��Ŋ{g�Q��\|�b���ҡr|�{̗v�R���y�㩫Ҹ��j8�ջ{%XS�A8L��.|�q��Y�3���S�B;l�G���?i�!�F���>�!����}��x���K'�9����yӮ�	��Ҕբ��gu�/����lj�:=5G
��7=�r�y6ʽ�t\t�V���I�%Wu��K�:��W%�Z�xq��v���a*�6���+k���'�^�.�7gV/��/�w}W�$�@(�B�X�}A���{r�`w,�'�a�	^�0 ̜�{�s�{����w�G�\�t{-���P^�D
��-�#���wJ��fN�=U[�ܳ�����<�9$ZfD�<�:m��'"�����Q�慛�:����m���_�N݈ua�b�#:諝xb��
C��v%�f����^v"4mwh��&��f�!��4�p�5�[L^���'Oq�Z\�o���W�h�tF2��H%@M}��j*p�T��W(eUwtg.�"�ds3Yn�^U�����6uab�P��&|�����``��}��`�;�%[�]��<��q{ه�.Oz�5F���1��p��=��9�TZḵ��7��V���ʠ��C=�u+y|�^��I����cs�VzBef�94�!���S�wK�VR��ڍ�k^շ\[�׍��� ���a˜�������̓�V�%դ�S�W_;�QL�>�[���SW<���mi��t &�JsL~����O�޽��{r�zg��ۅSYV'�y׭�;�����}����V9ϊ=�g�q��ǭ�����k		�pu�^1�|V���1��]�4\bs�3��Oz�_~��7�6����1&u�v�g�s�`S�=m�r�h!���Z�T�2�{KAf�U���w����\u�4��X��kd"��C�G�.�6��N�l6��pQ�_��ZF�j�/����T�nK���Wf��֒ڸ�:ܼ�jz�H`��)Ex�dYZ��Y���[�7�$�-�h�{�Hʰ��c��Q�bZ>�"��M��=�ݜڸ�a����~�q+;����=�z�I��E%~u�6��غ�$dI�hI�Z
x�{_#����n�vWL��pi�'a9�����j㬖b�\��y�':hL��Y����F<#A/
FQ뤜��X�-�$�.��ZW�F�5��P�-�x�TF2��M��L���K'U��ݽ\���Ϛ���A�%fkg��Z�8�~|��z�}��!y���7�E�2��>�5��Z�53T�%�ZY:]kHH:
�)-�\5 �����^Pa}R�\v��)��g@]�5��8K�N���>�Se�}ُyx2�reo�U������m�61꽤cd�Z������b����
þ�	wuB�ҕ���)ʫ��P��}e׸2��A*�VxfOb��N��u챩�Z���7k5��T�W
�m�KY}K�;4Z�|#q���Y�b�b�ҫ��nm<���t�hP˴'���cU�X��7��WC�GzR���m��kdl��998R�t�b��+�-������Ř�(�z�v&��E����~��p8};V��-�8�>֭�-���v`=��E��mfos��{��<��Pv)x'j��h��V6�lW.o�����g�=o��������cq�9���ar��/Nؠ'P�ZC�X%�jr�)!��gq,<���N9�_y��v�R��D�S��wGS�鍋�u�yPJ��终�/]���i�c���-����`,�w�V���=���k.��"���gS�-daz��O�������{�V�Ґ�/or%濬*Y���lz\�2�7Pso�����m.��|C��"�B�nm:�ל��w%�PXi��:�G�F��I�%u&�/Dtp�xWX޴�[l���3�c�s�M���:�9�t��N�N�� s��\=h�m�.p�%�yȻÍ^��g{�* �^���Բ?��s=`N"a�81���*��D��͉"�J;�Of=׊�t�=�ls26�:A�F7�R8>0Ƽ�;i�+�oTZ�屶�:Ո�ӱ2�G�<�'\�����%�=N�By�z�h;��;���Rh3�5p4�5��]W��y���V����F�B|�fX�=De$F�R(u�Ж�\�QS^|"����6��������$��:�뒘�Yn�o����lZP��Yn�k�WIg[��<j�����p"ؾ4'0��t.������h;����,ɼ*���n�E�[�{�g��yҋ����¬VQo���8ج�J!��g0t7ȼ�ܱ��m��7���w�����,�!���g3\�Ɋ�jqn��	5bS�E:o��f�k�_��;s�8};V�P=�ffe�|y�UFed�m���`]�橎,���Y~X�Q����
C�@�7\���:X0��G�mv\�//�X�܊f6�EN [YQ�u/3���j1:� \oD�θ�{�=�x�f�j�ʺ{��)����y�f��dH�z
�!Ƨ0p/�}Yy�qf�M���G)���6u��M��;)ힶ�Pv�v,�}�黛i
�==��A�lQ��R�F Y���ݾ����	w~�5��Bb�Ɠ�KX�#�М��h���`���C�_�ݏ�M�NX���#]gK8���͝}=��*
����WYz�����"\3p�q(M�(3ڜqH��o��,_#!��ʗ�Ѫ���[��ꎯ�����7�S�ǁ>�飑��{Pڴ̃�Jp�6�8���:�,�y{V��)kѕي���%;w��H4�T��'
	�}w7kg������,ś�O��)�qq���Gh��4a���8���PǷyԲ�m��0�jk�GI���8UEoD��%˂0�\�W�Gw&�V'��.]�R��U�5�Me��˵yl�9M����%���fi�^2P��ʁ�����ly|���G�c|i1��nb�y�Ft0��Y[9�f��"��L��gS̜�>�4���Q�;�4��_Y8G�Ù��3��MX$#:��x��D����:\>�J�x���n���J��h�Q�s��犌o��zU�=lg�-�_ȏy7�Bc�\��٥rl������#��u�y�3ݶ�ҭ�\���ř[�+���� g�>����A?-B���h�!2�p>��>y�M��4���DW3s�?R;z��V}�ǘ��#s��m�u�{=a�E#E���s��wtQe9�*O	��g��a�ęZ�a�˜�J;'f�EU#ד�A�v-�=8�U'Np�x�5��V4�#P/J��\�a�����Wv-���N���=�T8#;b9
iw�������z���l�q��x�9t&���yt<~�!�o�w]Hh������T[�*���R��gym�,���<���&�2�9q����){�4F�*�R/V*�|GwM"��볺U�����k9&�2���8���j\��7�e�s�߳0%���ı�.ۭ�������ta&�i�(r����u8.�T�<+k�5�B�����G�e�
S � �QYȪ��.��p2{{�8��e�sj���-�������R
�.���Z��x ���G�y��"�F[����E�0�;9o]4'I}�.[/���������Ss�������.��g�lT�!�}%�	�o,wuIqQT�������:��e	��jȨ�nû]̇�ӂK��쫴�oh��٬�nKPrI��8�I�3yX @�<ũ�9�ӮK��Tچt��-���z#�r�]Er
�A��]�:��͠���uG`��\��kp�])wfWD{��s���0�|�UM�=��
櫠���5a�9��c]K/�j��z�0ި��B�ݣ�����t�s�x`eMۧ���� VT��"�\��������ʸ�Io���-s�S1w'��6JMS���U�.��R��o7�>�f�8�oj�s�!�*�i��+��1���$�Χ��������Z�?�<f���5�Z@�/���J�H��:w)R��2[|r��Vnu�n�7����I:RWU�TO�h���8k4��O�~�w�c�8��%#�.���zOaԨ�/s���'�]̜��'�w�<�^��ީ�$�]xm��;!�1��})��,>��Ӗ^F�@���מ� (�땀F�,<B�s�[���\��\"a����n�)k�t�]�m0���ڷ!��Lb��R[8�Z�Bֲ_S��R�ob�q6�o�*�L)��x�݊��O��2�q6s0䉭�����E����p�F}(�]��j�d�5���O,Y6*�.�@"�p��4K ,�̗6ڱ7@�F��<=�ç�f������X��$ק ;-�r���=5�AfXv:)aw,ku�@rN�E].&*.���=}sv��	�2���Ɣ�S�5ɾ�{������:��7ɘ{L߸"���������н�&݌=�<��[b��n���Ζ�v�.�����Bp��o ��	}���e���_K��0�#�/A�T��Ӱ�N�{ �vL2%K~V��	�'��G:�v��o�$(m�����hɛzNx�st}'�������g%
��g!�q52���F����j�[�]/F��;�N(R�3����$@��K
ZK��n��7[�F�����#�����'�'�3+�-����ؑ�A�b�'b`��_S�j�c����mnfU���gn�(�=��L�(I���42s�	FGn�XGT��djN\f"�Lmoﲥ>��h�Ŋb�lvB���sT��Ҵ.aAz���$�I����ҶB|9�Mw���p�0d��Q%˾�'T0\���מ����Z|Qy��7e>�NJ<��Ŗ��C����[�� �X���[E�+D`�g��0`����aP�!U"�+U""1T��X�XVV��R���1*�Z��(��UEJʶ�Ȍ�T����+X6�b�j"(
"8[F�T�V(Ԣ*�*���-(��%E�mh��E�#mE�,m�Ŭf$Xe[
�d��`���$��V�DJȲ��VE*�
�*$��Eb�m��+F��m�(V(*�e��2++*,+PQJ!QF�@QJR�`�E
ZV"�b�EPj,X�����X6ְ��ԥ�-cJ!r�QI�Ő��iP��m�Dj�mT
��i\J�V�"��X���U�«Y*Kh*���Q�H���cj�,H�����R��0X���jPV�b�������Z�V�R�3Q�EG-Ab��F*���%����������ȰDbT�(�"�֨��}�f��{���6={'Y���K��۸
���Q��]M��x��Bw{�u�c��e�8�Qf��Hu��N�C�mgDNrQN���v%����7�wK��	�^l�"��,��W�g���gu�{��L�������5���Zt2�&���r4�i=V�
�կ#41|�I����&�Ԍ���¨�DoE6�Mכ�n�;o��|�Ű38"#�[Pe��	C\N�&�S����* �s�j�VeO]�z���c�:z��o�Z���U��ݷ�yѕZ殇5�d�{I���02���lXKY}K�ɭ\S�O�L
m#���Q��뷭��ݻ�.�Í
.�v9>/���^�\L+�/�����X-Z֮|���~����TR��R/���׼��_f\:T��ɾ�W5�rM��V/l3�nzV�s���1'�P�^�{�'g�^��Ij�%����.�a�C��U��ڱ���[Ŋ�ۛ��c�Wi!��6�ٓ�n���5��V�e�BيZ[��5(���4�������3�r���,�0��Ux�e�FU�B�k�ʼj�Wl�Nt%��d+�����`�Qe�����	�͝��d&7O�����c8i��;۽c�����wd�:ޥ��m�a��n{'lrQN��pQ�_�P�I}p�m�U��w=��bW�q��t��>m[�9y.�[��W�{b�7�򳹂����륫�/]����1���.���Gl��g*�cC�&�k��NfjA@�c*sk��1ڏ��Vw[����X����Ue
���
�qw2دI��>���̘nߟm*^����Ξ�#��,ǳ��{$M�屚��N�i�I@ls�H�r:�q���RX�^�|%��m�m���)[�u`��	"��U���ՊA�+�p�p��^Z�x_,�.z�J\�ypNX!��h:�1��JQ�ѝٷ9��N�h(�\��f�J�2�;�H%BhMy�'�EM�)[��35Y�p��o�i����yW}�[.��B���`%���l�������,�}S���u6��N��CAڭ�g�e����t�]�}��#~:Н7��w�w���o��n�(��ʺ4�v`W}��Qt�[��M�սK�\E�TC��Β�ȕ�u�l)���!Ԛzv�9tDȮ�Y.l*��8�,D�|�X��:��tť����'��o:��OW�����W=C�
��d�y�'('Kͽ�-\>_
��§'o���Z��ܣ.�pה�d��[mw)�_�ǿT��/Co���E�VY�D5��&ر��c9�����ƴ[��9�����V�Pv/y
����4kP*�ư�'��)T�\m`���I��6�s����[j)�]v�3�^B���p�o.���UX�/E�^-5cJ�B��j8��nÞ�Z�mtͲw�Z̺�Ѻ�6��@N1ByW�4G��=��#��]�;��׼�}�3���FU�=`,�`w)E {Q��_��eZ��M>��gq�]�1c�ކquɴ��ۊ�佥`����W�Qz|ҞR\�=F1ZξWݘ�eY|̼���I�̃I@�ä6���pL�F����B��6�)=�4�O���� u�<4s�)���_���_� ��(��U�+ {��[�Z�ޤ��H]����3��NUx���Ϲr�0���Um�@���u�&�=�}�"�A�[Ӂ�\����i�9�;��E#'NJu[��82���+�&^�Xi�H�*	�Cm@|j�Y�F��k���"�E��W��^�%����U��\�N��e�Cj�5q<V�jR�̓�ލ�\�z��&�f�|���S���Uk��M z�)�l&@{GiKo�$��e�����
��H�������� ��A�<�G�s;�2;��-�''m��KlD�=���fO�����S��=E�9�
��P�u��
�fR���sƢ��}��l��*[�Pl����=����>cH�g�/k3ثC���u�_8N|��g�O/J��� [�2����v��&U����S'���>����<��ҴjCf�vY,w�ܗ���,�$uxwS��jpAn�u�{ n�f��@�|�wn�k�<��v
ۃ״�(��oC�~ɭ�-
p�kɑ��c��p#:�Hǰ����Ik�,�ӹ��2�Ԧp�� �J����1;.Rt�L�K�]��лƹ���*H���Ʀ$gu@�*x5����
�jz��H�g"��.CYˢ�s�t���W¦C����ҸҚ)G�����V��d�,{r���y����\b�a$0�a��J:W�B�c;"�:�p��-��Zr�^.]�p����O�}�^ʈ���]�U�$6�O�@S�Dmu(�l�\ҝStF�SZOb�:�1�[R��p�Ys �u�jp:gj^L�D��A`UW�`sB�(��l�e���5Y�/y_�u�P/�NJx��s��Qc��"�W%�È���%��`'`���]�z��0�CV	�N{���ci���b�g��e��
�/�K]T��.��Ƀoa��7���G��tYꦀ��h��������V��LV��N��#D�@=v���nu��Ͳ�z�k ����g%C��'k�N�?�"�G�����9k��w=�w��*����b�
; ?$�
�(S�4���/���)�Γ�*|U�ĺS�k����S6Sȁ0q��0Z�!� �U{�����O�E��xD�ߊ���Ꝣ�,Y�է=�*1����7B�>JP@n�j��A�O�L
j�eİ����	��sA��7K���H�;�{>�전W��ܰ�l8B:�dh�O����,��JP�62G�S*�31����f*��7D�:�3�����s�����ӨK�]'�ar�7p#{�;�Q���g��NM��T����Y�p�r��#�yk>�s������T_u�7S��X��P�(ob��eZ��ˠ-�~��dm�8ȺB�-����A�reE�����
����ix�qK��|��ڍa>4a~U�3U��o>����ʔ#7iU�ڙ�v{U��e�G��t[}�4�H��]z���\lt�b��6�06����0�&�@�b:�N���IZ9q]<���Z�2�T���vN�rG�S�Pz��5������R��<�ZEf�:�k��z�m���onu�24�[Gɐ�/2Tc�����v+��z(p�Β���El���<ڹ�w�!� ��Qnz
��e�s#_�"ܹuqO��蠴�J���O��@�2��8��$EL�u]�Ȩ�AS��][�x��ڝ�q���ӹ�E�*tf9j�лe(�Hj��6�W�`��Fv	eE�F�c���q�ˇ��C؈�*T��[ROJ����7d^J�"��2q�� F�Q��>U��ѱ���>����e���8���+6���c%�G��R���}U8�཯�ܞ��f�*ݼ�7����J��}s��Zf���εx��ݖ�[N<5��|N�:Gz\=���u,������y�u��!�퍃|�Ⱥ��r^�*�5��$�ɒ�;Wo�5��pN�I�o���@*���*w͞����dM���]�l3:���p�|:��ƒ��q�XbT����%C�q~�N���j�)rG��4<j+�.��4��{cw��11���V���,���ЂS,G���bQC(�����R6rK#t2�q�q.U"�u���9�EE�D�r;z�"%�hUC}Q�HJ��QX��{�.�d�.I<mX��#"� �dP�G#���BuMÏ.����]��]�B=�;�7Ǖå?_J�_è|�{)�-�U*��D|E�7;�F�ˤ!���̓3j�J�<�l����%�9�Pm��'���u��R&Y��m�=��F��$�-�*����>��!���w�����^}CI^����;+���QjvjU#b�L���2���O9��ccD(cC�c��w��nA�u���h�R���;1s�ʷ�^U��m�����u^k��~�s�å��JY��iۏ�:qN*��<�Q1�F鍲���s�i-���]
Y;��`"�a�"�(�	��6�O_�DArF5u�� lnX8z��ӓ��^Ͷ}�|}8�*%4ӻ��^�~Y�lƷDToyFpg`�{�������d	����t:��0Rv
���&�g{k�/`��4�T��2�&x�W�d�_Sg�O�q�<���'V�=��]'��v�׼Tc�'	Ƕf��p� X�O2�}o,��?6ht��8EŊ�	��"zB��j>2:^�d��WGK����u�|�Y�J7��{f�²�گ��E�H��B�[�U�:� �
eu���#�ݵ����ܻz�q�^߸�6veC�3PR�BPn�NςS$��h��tF�����ۚOM��)ۮV�@cd�&6:Gaʬ����6!91@�TH!���ە�+&ɽӬ3w����ae(����_�m�r�G\ߩ<�>n�J��X4�����"���%#�����ot1F�;��PE�.,p�*�LE9��(K@�b�V�q��|��%z��&��ꈩ~���x�.�z|�+�?]<O��U�C骮�ov�ȸ1�;�1���y^Ug�ZڅOs!���AS}��S%Y�7T͊�{U��^�2��i�M6��W.Gu��$Ň�":��=�>ْQWR_R!����$f(����3oǹ%�J)H]J����ۊ硈�B+.��/��>R�1a�1D���1��zj7¶��+�ˍ���y�[���ξ�`��V�	�6����R�E�(wY��3���L:���uz_��֤y�];������T%�J�[S���LmEpejb�.*xzp���3��嫼�Tz�[L�$����ޯX.+��r�.9��}G������Be"/eD;]��t���{"�ğ6c'���#���NR��~���By��{G��!��Ҟ��R)�g^��7W�]������I�t��ײ�z-!W�b�T[�z+�MlB�+��g]��8�\C}fG�֌�=�rnNw7�]{�����A앆�`�R3s]\��`������;7\I���5>��w=^�[/<&c�)U�U�$��^�V�k�Dl�
N�ّ�h�Z�ө�wMܱ�jF�=ڋ�c��S��;R�Lƃ}��V���&`4��CM������w�Xl�
��o�����XO	~�hϯ�0z}����
j󷹓#©:���7���������,�6��&;��x������]�T�����7+�k���ۭK!z!���1�N�j O�S�eA'�]n�/v�;��w�3��;8��/u�=1u�BS�2�Z(�n���/��x��ίa����7\G�PĮ�r;Xe��\k��f���YIn��tly���P���#q\C��@�GMW��a�y1V�磓��o$H�=�|8�cp����jOA�n�ɔ2�06�]�t[3l�h�4�P�5%X�[��%�]�M����CcΙ�s�ܡ1��>v�]OU�wU��pTߊ�O��n������-�F�V����b�������=V����P	���#D\>���)��+!��6j�Z��u�y�R�W$�A�`g�(�)N�Q�;�Ty��Q���+�)}�E/r|5�9/{$�����N�w�٬�s���ϫ$!�\����q~��Y��;4l5c$q�x���n�Yu.v�A�z���]#VO���vTle!C4	q�]9��5n����כ�f&�jӦ�$��ɨc:�̐�a~u�3B��-`���]2P�;HC���t]����B�����oԜ�!hSJp��b}��# �ڛs]5rk��އl��r�A��[s�n��"ʦ;���Yqa������Y��D�6�!>3�,G�ʦ\o]�wo1������P��)p/�4�
�v+������瀨Qb(p���qrE�h;29V����P��48���0k�Ujk�k%Ws��Q�}���=�$ I?���$��H@��	!I`IO�BH@�HB���IO�H@��	!H�(B�� IO�H@�r��$�$�	'���$�p$�	'��$ I?�	!I� IO�H@�i	!I���L�b��L����6B:� � ����{ϻ ����y��HT�J�J�	B���J�)T��TUPEB��Q!�*�6�Z"����Q(��%UR*��H%2iGp�v�P��+RSkmV��hd�h(Mj��\�f�Re�Cl�Եa�	J��V���Q5�-+���PUh[Q�Rָ �  ��Z2����rj�L�-aD�e���Qm��AUp�S��da�D�¢�Z��Z�hUB7 wt���4dɶ3V�kmF�eRmkm������u��b��l�6m�����%]ۤ�,Tm();8���ʫ�R�[���ҩ��Ӧ.�:�-
�a](�Fn�:�v�)�-��k��e�&UJ�5�̝�S5��Dl��d��4��    ���R�MQ�40 #L&!�� �x�%ET�       �2b`b0#L1&L0j����R�� 	�    �2b`b0#L1&L0I��R�&ML�2b��O)�4i��~�S�w��������voZ��Y!$$��͒�焄����IA&@���B$��@�BB@�#_������A��Vm$T��! %!�d�	$$$�.�Bq$$���>�ӯ���������l�$$�ʼԯ�����%~��f�F��

(E��/�u��U�>ŭV��x���
�T�l�i�)�ӛ��~�����;�bR36R5�az�vn�e�хYK�<��X,p<�q���N���Z��f+��7in�D@�E0�uimtZ5��%0�'@̈����N�S�F��w���G�m�:�ؙ�t��a�V6u)���=0�#�"SjO�1͓Ec�˨���b��騞^�B��
�Se�ۨ������*�Ћ8-(iF����c��$�=*��L�᫋v��"0�AӂJ��H6��#f�e ˁ�Dfl'�D ��[�+�Y2^|i^���ZB`�@� �5
��GG��T��	h*�4�efЏt�Ȟ;T��sq�i��R�i�pf���-Y����)��nGw�w/4�$�z�&^�xu貞'II2&�bȲnj�lSjL�3rl�#�j/��n��豠b�s0$Z�m���u��TX9X�R�h�*̬(UPƩ1�I�uy��˂���R�+ (����M�si�������[uh�u�4�"H��&|��{HX��ڄ��EP�aP�i�J��kBW��r�+�[` �Ӣ#l�Hd�Zp
�u�9knұ{f�;_Su3sm0\�׍�.K�ͥl=�3p�j�טX�3aHR�M��^�ǻ/e3�����#�R�^��l9����b�����iV⥉V���G[�m;r�n*2�h@���Yy��R�X��⼗qJj:,au^���p;����SMc��5���h��j�uo_5X蠪�*ѦM*72ɰ��D(e��լWe4���q�R���cS�w���n�sD6�P1�ӊ;�L�\�dƪ̂��̧Z�F.mi�j�Խ���C�F�RJ�GjI{��Ř���9�IK7�jU;Ѥ8����CvH�֠��JDZ:��#Z0�Y�U��K�y0��]��Ù𴱤2Lٻt�%G�AIX���ٰ�dk�NT�
���3
	I��c�I�Y45�`�7v�#%Ă�栣[v�'5,YZ����;w�"��Fw>{�eA��k�����+�L�-|i�HB�>Q�Y�C�e�k�8&�n-r˴q6��N�]���h�*-��j�wz�S-�(9�9���n�X���`<J�p��ͺd���`���*��&*t�Mķ1Ԩ܆Y�u�K6"�zh�:��
��o6{��ԗV˫5C��i;Zu:nci�:]
M�*��2)UeV�NUh[o,�2�H�{D^�p�����0b��(\��St�o>6ග�T7&.�5.^K�1�Ix�৉jzU�ЦG������>�5t�K��5%�/Z'~?%X��=���(�.����ޜ�D�Q87]��G���4NR��30�]<-�A$P�4!��Z+"�'(�z�*շ�ܖh��`2��{J�g�M�#UY�B�+KU���v5���C
b����0���o+i�T��&��J��ٚEd��ԕa�RXJ5@�0rȨú�t`.��
�+�;�Q;�vr#�\W2 ��i�O1кL�)O�c{��VHF��(�b�p��D�5�^���î�ֺ���)�6��X�.�FX�E�mK��VH�s�v˚�/�o�tʛ���,:��J�`&I�1��Nl�Ԇf�ma�d��Օ��@z齢��țǵZh���ml�YD�[�B�eX�f��-c�Sy[&�K[��SI����7�p
cڣffޫJ�:X0�Ʊ�X�f�:+S�T^]�y�;�i��WC�p<�*�CdJ
��E)��N�T��k�fGB��&D�P.����N�,��ت�*���W���8���ǌ��%U梙c.��g׮��h�{�����P�+�Z)����7�V����5Y��-�9YtCߋh�� �*�ݫV���w%��)ܬ�W
wwYGeQǙy�7b�B�<�&]I;���i3�줌h0(^� nmE���!��,M��*d�X�n��k>b݅*�����:���t���Vыsvnc���̏)Q+05��UޕD�E�%[J6�Svf���L�yGe��%CA�ɀ �:v�4�h�N��ZI��J����}qSMʢ�g���&l����q=N^� �I��7RY>����A�'�fT:��$r����e��	f�m�H�0n��ӪY���m^P��[E��e	�sTq���y{e���+g�Ƴ�QM�~���o�?@c��Б>㮺����}M�i��2��ξ��V3��K'�QJ�n�IV+�IU:RP��s�V��u�N����u�"0V����͗��Cμ9|�Q��W�j��6kW��L�C�T�گ�E�NVr�]��t����������tچ�R�V�\AgV��9�54q�YW���ԭ���ޖ!����;&>��9B�X^��6���9���#I�&��0��+N��Z�R��խ�[؝/����G��jձb�mi�J�E����o��B��wՒ�a'�(�Q�B�����NRR����~GNg>�헏��cⵎ��=��*|I����+E>�n]:���I�T�5�5�r��P)-��� N��H=���d�-�����sٮۮ[������l�;�v\y�����/�X�5Q�}/�i�|kkb�qb��l1}[��[���)	ὕ�:�V8e,R{��r�T�#3�&uAq�Z"��x��e�PI����$ܭ;�np�N�H��UҸr�&���%:�q�ܝ؃��Bn��������i��I ���\ҡ'����o�eG,�
��R�*Q�Y��2m!�[]V�5�:�І�g�r󘕭�՝�[������`�K��MWh��H�Yz�G�N�j�Z���W�c�׼��n������XX���b�j�Ѿ�r���;�ON�S'��n����ݡMWb�M�9����Z�IP9�M�6��N!9��:�nm�e���q|V	�b	���;��v�x�t׺s��H�MfF�����n�9��Z9F�c����RgJM������R��*q2��t�l���>�<�hG�3~�s��޸}�(f�]ע˙d.7V��w��l�nT�$%�X�Av�3W2�����=���NJ��-�e�2�5N�슍i�yX��WB1�&u+��y�)
~�t4� }�]4�V�+�nN��6� �Ab�d�s�-�cr��IGx�U����1RjqdNQg.��If��#;�1sw��olf�&ɤ�o�VUᝁt�Hm�&&�kz�e�/wz�.�%2]g.�?)v֏*0��^��|�:�u�^l�X����πj�A�.�gE�uqV��5��͝f�\v�'�+Y�v�Z)��u��Y��<�����_R�\�yu�,�ʩH^`��0����uF�TMKv��+4V�.�s�En䙑�[�	��K*pގܙ�N�o�2��T���w6��e��e�Z9�����I����g�|���S7`=��*�F�}����Q:w�Z�:��K�^�$ȧf��.u��K�Y���#�-�aN������P�u{+r���Վ�p�ڝ�f�Ӥ4M��v��U�Z4�պ��<�/V�o87�6��f���-�>���S��]�7�yyP���[��q9�U+t��ˠ��vF$���I���pոʎF.�]�c���]���;�f��m�=h������5ӦZ؜fv����d˻�6��� t�J�\b���yS�i��Cb=bθ��ʙ�����7�=]��7�A���t�\#�,'���*�ˣs�t� ��tx��p�čI�{�	�~��I�*t~�m���)ϯk
l��1a��@NV�1u��mZa��x%�� �Ý�*��I��X����΅�工�G/9�ꝅNZl��ѺɝܛEL���V��8Uk�9���_vͽ�T*��GF'Vhs��@�Q�7[��]��}7��0���z���5S�A��U��zR�J;<�rK7��(&6�k����X��.qoRgQK)$�%չF�R�!|1m-Т�*�;��P�m����s<�Uf��}ee���7�Y�Y��H E�WS�ss�"�Eǥ�����q�EI�鶵����醵�7�z,s�}W2���P���{6⋺gZ�θ>n�Y�GJ)r+�I-��RI�$�-��Cy�rWi{�'R�5�]zpc���K�k�k��3;�1�13��L�ĩ9O���uCM��>��9�×q��L\�������X��%�ٝ.�
��E�Y�);��_wwUq紥E����!��)hU��坤*�k�+���EU�r�7�2�J;ӽ����gI�u����!N��"n��:�Z�g2���Zf��[;����J�.L��st���5�?\�v�>̓�x5�;U�9�__u�o����I�K�U�r��l7ʫ��دTSw�>�����l�Z���F�&�J�u�N�E�
�;y���{�:�o�;�}���<|~������5�RBӰK��2@$�>k�擇�,$! �hI!�����ג�U���������ky�Ѻ��$��QQ�]��Ќ�ŋsl6x�I��4�����s�7��;t��;�%�w�RS2��# �dO��o*�]���Za����*Ps�pY3��N�1amǧ.{�Hj!n���Kpl�R�Yy���M�WRAܨ�V�}du��u��+zkm���2�9��l�m�Ϩ�Yh�w�a�����z��p�B]�f��;p|X��I��T�U(�]���5]r��BImb��(�$m���jí.��3���(�]#Gܡ�cI�C=�V�u�*��͐���I.
��r�wܨ\?h���Z������qÝuj�k"���|g���f�4������d1��g�]wjmN]V(�h.	�F�J��9w�8�AĚ�:h�Z�k��MV̰�e��MT���j�kj�:�6���]����gF$-�f��um5���V��:�W��e=�XwV*v' �[�ݲA"ަ�����Mn������;l>��uv#s6�2\WAR��<����͕xcŖ�γ+���BӮ�Z�^�6�����*wA��ۦ��i�˥e]����9��c��S8��C	�C���ZM/��j٩�DzV����h����X
��|XY����u�/�ZB�er��Ǵ�eHY�]��se�e6QܤvG���_a07��U�+��:�
s��)��hT8"����=u��Z֜��oT|�r�uʋ�ؐ�O���Ĉ�T/���e�pWC�����o�nөO�B�f��N:Ưu�}�]N"�����(r�[t ����33�nȖ�\6
\�*n���tҧ؍����n�SW�Ĥ��1
�f�5$[Cfӧ��p�/!NR
�q��h�Z�U��@�k��ŵ�����]¯w7jS��.[���ZŹ��Jn�T贻�B��!������8��Wlnn|���3@���$Vܫ�rG���Nql��:�9���)C`ȸ�/��L���V����i�a�O�sX1-"�7"���Q4�1+��{N��ؙ`�>�&�1�v]�V�r<�Ln��GtE:��F���r�*�W07�����E�"G�z^��ً��ϊ��(D/Y����j���J*�Y=�d��I���<rX�]Z��p`QT�#JNX^��W��J�R�8�A+j�4�+�r��H�wن�#����T�)D!*ihijm7����^�j�=&h�nkqgv�!�;�9��<ڎҎ���tFܛ+l�\�q�(�g�j�]�osc.�ɚ]���l�K;���jۆ�r�C'�,M�ˬ�X��2S:�U)�����|�T�5TN�����vq�N�$V5v�r�"�\9�T�8���&��T+d�-+�!����Y�omV�5�B�$�Re���:Y-Х��/��aՌ��2����cD����<9ݪt/�j�dN�����u�6]Ԗz#P�f�Z��S
ru\�l�'�9����,���Ur�=4��\�q�']�"�G��[a����֧�76��tї�ֶ�u�M����ڹ�j���'�'��l��ѭ�!1,�Uo2D;���R�竍�*��vu�8:�ֱX�0;��G�8�A�8��C��f�#.��7�����VծU;e�W�3V�J����'���i��x�q�L�@���_fVt��Ǣ��hP'm�i�P�w�W$-�6��k,���ݔ�yO@��N�)o���F����iD��vҬ�˖ҍVb/VY�v�G,�����P.��k^���)�L��d�-�<�Dt�]�:R�Ief�)���0�	��ֶR�4EDF��&�n<�N�m*�v��WcEws�X����k)�ʾ�o����d�|&+/�c��
�V�4�z+MϢ�;��x񽂦���b��Ts1��]-��w=�qgU��
��7dy�#�u��ؖCgb鱪�����a{�o���{ٖ�[�3�˫�Y*;��'hJz����u���H���k�q-x�-�h�)�pi��cٷ]ؒ��k]ge/U3��\�"�,n�:�u��w\e�ڞ]���P�=�s�f��ے�i� %��7��?N��������'h@�	٧60��@St�B��f��M���u]EH]���d�ݤ�K�u��X�gL{��Ni�� ��m��C��ђ�z-F��?�����������ǝ�:S����|'�
ȿ���V�9P��X����&h_�S��#�:�WXU��弆\=Bp֌�B�d�����S'O7�}}y����b���v�s�3(�z�ڠ�b����薾]�Z�����!���:��;��֫"cq�}ff�)B!���ѥYu��4�����ڢ��l�TC��a�R�c�^����y����Sl=�N�ʁ��n��6�O��'N���N������9���;�������x樤�"�)CR�!����Q_}�LD�JB�B�Jd�0�`�XL)�R���II�L�@)�
Ha�� ���q��0����KB�,�B����]_���B4Vx[�x�(j^���@����Hj%o�5i~��܏v��]z�mS���!�7�9��)l=L*�~Ѯ�;�=oޝ5SߎU3�zrF	ً�<���.B{���=mVܮ��6��f�4�r��c��p�ø������n��嘴=M{���N�x	��8n����nnG;�s��>�%ٳ=� |�V*�*�R����.d�� k;l=Z���S�;.�J�IU)�|&ݾ;�5K�;�Pu���ߣ�οZ���c�h�h��O�r�a�_>������= �������Ift�^OS����\�j�t�NpM�"�]-V�E9����G3�@Êt�G^g];2�h��}�b�cu�F!S9)
> ���1 l2������|�hu�ul���k��6�l/��;C��׽�7�콂sU�[�s��%���*NC�����uϷr�U�8��n�/vlSCs9���9w��^-v��:�o�5�'Ҧ��*�z�[�Ĉ�[���~��rRz�d��K����.��%�qLi>�d�^S�>��ĺ�M�U�vZ��NU��5�ZN:�e*�Z
��>8=��㧥�T+6�)�u-@�W4��h�t ޫ���-*��e�ƮV?!҉�<uo���	R`s˸�C �y�%�L��M�s�� C.Ӫ��Yz�5')Q �
Y�v�e-����
^�m�O�񫕲8�]{=)U=+8iɵ:y����W^��s��qM��
�T㒂�q}�a��.��-z8��	�f�����ܽN�Fr�v��&�V޷9��3	fQ�l����������[�r-tI�aN]�Ƹ�7�Vp{��;�F;��2֙X�&܏|g�j��\gt:ݨ>ڍ�Ū��}y�-{j2;�����{�7�B#ht�}7�uK�/�Ȋݭܨ�wb5�c�0j钔K���At<���K��g��X닇%��b��0z�TL�m���r��
���۵��a�ۚ��o��/U�;:�m�qd<��eSq%�r�y85�m`K�8OsZ��2a��8�]�v�G��?c�vwv>%���0&�mZZ�f��A�6��*�arl>�ƺ��m�<�]ct{]b�\�;�3�#1ٓ�;,%Gbİ��RT�X�>�1�~>����yU�7�a��ϓ�8X��g9��!M�r5�v����ʸ��¸�I����WCC	��fy<�/�{[��?�i_������D���a)ֱ�(��=Ъ�G��>N��������w���F����eJ�u���*�璚�}�dZ�
�
1e*{p��=2a����<(�I@��9Y#�Wu!���y:���_�J,j�s\����i�m�&o�j����r��aL*��x�ˌ�m���L��u�`΀�֎�e&�S�5�o%�����3|*a䫢��R�B�T�F�byF}
�P��=RO�3��xMgkS8�KBZG.J*��������$�JЕ� fjK��m7SC��,���Ss�V�:���Vӵ���v��/xd�ܨ�����ts��s��&˃*nu�}����2s䖬��ɉ[{��?뱚�!d�+���	�=W���YX�S,�ɼd�L9"q}X*�G���8D<����W�ߩ�}#Sn��ҵs���k�p��"� �r�pz��0���"�E��
c���=��de
UF��"�^����h�N���i���8�U���11��׊����3���a綪�s�o���#Ol���rm{0��MV�e=m1q��Z�S�_����ܿ��)�B�+���^��fT�KX����r�*�eJ�{r�G	ˇP��KgI�`���wt(N��9�x��M��to�[T	���jރ���]���,�N��jj�/o�q)��)��U��w=�OAS3z�@��B�P��
�����w�5zù㿮�>x9���O9�+�+�ɕ�n!����
%8��[{���
�"/S�b�mi�{��s ��vV�}\�r���@�9���S���:�k�D��5�@�F�i&�;�����/]��Wn=W�ZwQ��4����w�J�j���5��z�p�>�u�Q|�\.��iWhł�4Lp��XF�r�bN�!K^t�*�}�4ԡD��^�;�.I|�U�l�;k\����k6����e������C�*r$��VWU��a�.��p�6��ƃn�X�C]����i�u�bs���Ӻ6��ۇ�>@�I�ӫ�����������u�Y�G9�����_���AH�y�����R
�A��>�+#tILP�����EYTX*�A`"��hRBS	I(H�"�R*,�)$Y-h���X
)�$D"�b �"�)�Z0d���������'�t��ו�K�WN�i�/o�rs=��W�5|��tl��w;վ>0zU���РO��w��6җ�R���?d��,r���^!��w��Xf��N���~cP���f���'Ж�D��1��~hd�~�_���%�8�����GewP�`���y�;�a��ˁo�ό��	�ۧv�5�68\�*{���Nlp�P(@J�G;f�ø9��kcv�y�8~c=�����}��
Lĭ�ǎ�A.�1�8#!��N��t��!9��4�-�������Ww�j�+1�B��!o+����mr��ھ9[w������Y�2vן�cxM)0��(�H���aݩ'����ُB�I�'�.��F�2rohT"�z:� ],��j�]A~�2�U���ˢ^�n�3&UQ�j���O��ܣ�䤣��K/�c�s=�f�!ECcPS\�o;G�S]�+��I2���'�X[C�^ڂe��eQ��s+)�ʨw@�mڑ�ۺ���m�ŵ��%fq�3p�ld�ځށ�Q3m������΍�*�T
�rU4��=���M먼�kB��88R��ͧ&����aeHg�AG���{F-\��N�1@Sy���Ҧ��n�'W{�ّ����-Rk����Y��b�ZDF+����C������Oo�<I������0fQ�o���x=���'?c��[MIi� Nc�N�
.��/'s<�h.�\y��K<��SI*>��5����C�3s�,U�&)�	��1ܨ_�?[�������mG���^V�뵯����`�G��k��n�j����θ���$�F=~�KrDnj�=������E�U�IW����X����S6��Jgkm��;f9{�q޼��������1W���暈p�����ޢy��)�+�&�jf��|��v��[z���;-TKM=��OV+�����>��c�+o/7"��/����Q�
�f�~�ӯ&ѭL��>������6��/�q�"��6czik�E���<��x�u�.sw��r�ؽ80�r.�h�����Pޭ�u9�mԗTt�5������^Sܯ�.�d�&N�@��Lnd�����[ñT�O����%0�z˧��y��mX��5�u����m�Y��i��c4n����L�+�Rg���\�ܣ�j"e�d�C g,Mjl%���ͰrE��2'F��le^Hq�G�3T38����D3}���n����֋V�>��R�G�X����A�a[�>���m	��{bƸ�[�����Ы�Ȼ��B $T�${Ǯ7�L�ۙ���B��*��;�/�d;g�f$;���*��d'�%�٦������x�%�]��!��ʾFgU@R��g�s��[tr����n'�d�<���<��W5��nwK"̧�U{��9���R�fµ�,�T=ӋR�0��3���n������T�(t����H�+���&�s����3��
c��A1f��m%{˫f,w�ǅs����7�l	i�::fv����}���t�a)eW6��y����<ڧ)�gzS��n0�W�=�3��ٞ����˫-��z=�:[b��K<4�[��j�(wp�3�x�����}���l�免}CU���zG��|P���ˤ�E&��m������z���3������	���/?%{^׀/�nG��Ex\W!g���Gv\��\=3�Vl��a�2�I�|F��h�j<���J���al��+(YMᔝtK�b�����E�M��+b}qÞ'ۊ�r�4�v��E�����xJ��Tk�Bꉘ��d���te힭��>a�mx1�`�e�t�>t�΍w
�z��V4Z;���d%�͑3 s1�QD[ѯp�1����ű>�ת�;��lV6"��Ѐu��v�
�G�V�6�g����|8�J�aQ�,��b�y�ѝ��A�VsvG"�L�)u����V��o:��if�v����4���ki:$f!1��&��aKY�����?�R���%���������8*c��.���ʹ�����m�i9Y���M�t�]�R�+,�p�%vU�(ݥ�Vi��B:ͽr���b=[dpծ�U�G+�mHS��h�?VCQ��7�.��M\p�K9M(\��-w_*�u�5"θ�ԏ��Μ����eK�6f��v�j���M]���/5[<�`1���hi��X�A�Gۦt^���u=�+��Hwq*�X\�����%kj`h��
s[Vﻲ&�.�s�����:Ϫ�FN$IH� ������#)n���B2�`����(�,X��TQA.�LF*+MD-�Ī
ER�RRT"Ŵ�
Ji���`��U�)!L�t��Ƙ�H���-*1R���U�]SU�
TdUQU����b]U�V�e��g���[��^�t��vт�#
�8��/����n�?Z� �o(�#{!����jZ��߼i��{O�ȕH�����@�+���N�쎺#�\}�vjI�}!�Tr0���3$�OI]i��s=h��H_5�G��4�8�ֿ_�8z���ԥ����M����ǹx�C�[Q���-���7�kry
�̮��^v��A��v�ְ��Q>���}�1���:�g���$/��������>"$#��72^	��Y �ڣz�4�\ٔe�[�;�zf� 3Ր)��غ����y?�A֊V6�2K�ޭ��h.["���q��/B�xP;����1�i)�������n:b��/^t��6�j�N髽�Ft�?��w�&$E�R�enJC���U�ۯ.�p�B<��֕��q	}���ᅞF�n�V�:j�J5�o�%�C�{�rܝ�xM{V��l�;1��`#�U|���������3ۢf��mP����'�yE���R���E]��hLg5�~`#{2�tM�I�E�k�si�]�L#׾����Nhfs��N��#
]K��igS=SOv���ڂޮ=.��x>�H.����}�K��{�mC�^W�\�j�U]�8��zԶ�Eu�;�����M�1z��K�U߇j�k_]v2�s{�`�z��o�/>&����"ҎdeU׎
�1��|l=hF����5ݷ�c��b���h�L9�Z�SW�^B%�r��y�>�&�P�"�*�#�`�g����j��L:}��f^�������}w}b6��*7%��}�}���[1��^�7potl���A�?<�t[�2/D����Kv��ٚ�U�c*Z���6��Nt�G��E��3�<�p�Rڧ�Z��b���?�С�+
p{�=����'�K'3@����T�T���U��z�tY!�9�����g���D:}��WQ� ��Q�f7�D�=���z��L��0.ЪW�t^����m�y�G��y���1F�0�Ѩ�%��Ь��*�ё^�`��ż��v�˃{J![�N�
Z��|�ּ�b�]�Pn���S�֚[\���x����*�!u��#}�n�����`�=���X�s�F����I�����]�AZ;v�
�i�̙�WRhupC��K���R�,S�k�.�ޭr���T��÷PH��~#�艻nc�ag��71}!�y��s���s��>���I&L�η�j���I�E���J�Ij�
i��)��jHu�� c&���w&L!�9�)$�&�:ɴ�i��ˆRC;�Ԓ�]c�=\� q	�&�(I�!���@2�N�P�HY�\�α����ChO2C�I)���N�i�>$��e�IĒ�I2��I�w�w��!�$�y$6�S'ϕ$)04�i�a'Xe6�&P�f���}���y���R�I�2�gt�k�BH����I6��wY��� O0�H�P��|C�CI:�m�ē)ި�`�)/��;��|�@��y�>!OĒ�-<�)��B�T��CHL�l> I6����oXϽB�C�u�b��9�Y5s�Xώ9���I��4�A��m�{7
j��z�#�=;�꯾���^����Z��}��I�I&Y�Q!i,>���O���1�|i��kR["���<��!��iL��!�2��!�C�����=�;��C��(ēL�N!8��|I�q���i$�ian�9�9��; �O�	9T�"ɶI�@��!��8�[a��C$�$����o	Ii��K� i�j��l���O�<�XN0:�RC,	�����שe ���2Ȳp��RR�N B�a�9U$o���� �N!L
a�!�He"�e �%k6I�v��g*O�)��f�����\$=�i$�Ha�>4�d�P�))!�(�u�l�u>c���	%3ܩ4�Yڀ)+�@��a�$�Cm�>0���>$�&{�+<���m�ܨKH{THg�!�'���I f��,��N]fL��Z?4MEY�	X��y�����X�e�V��Z�#��HI f��}2u$�0�d��|L��!_J q�C�L�d��$2�B{9�9ߞ޺@�&�N$�|a
a񁔐�L���!��!�hCI�T!��^�վ�4�I!��Ēa�RJz��I�@�1���I����߳��!��h�a���|I�HH<������c9��:r�ł�XO���ۨ��Ux1��Lׅ�|��ҟ�ַVc��bn��H��˥s��d�KN<4]��fkK"w���A��qպuΪ�߷Ƥ�H�Ր
�F���(��^�Nԣ;fܓ��gF�<��ĳ�_��������{�/��Yq��8At���Z���	��:�״ˇ��#f����m9�
}�ɮ��/�/.�������z��k��Z2s�J�9+�`�S�K3��#=	u���D޿07�׋p�}�g��:� ���I'!�/,]b��',F���t/޹����C��G*{䐵����d���J�V��� O#�T��e���7m:͡�v�t^��	�˗ưY�O�8f�<�J�j��Brbko6�[M�چ�(]�ƺ���(魵E�Έ�V��־�5Iwm�y{`�o7#9��+Ֆ8���;Z3��tڙ%f���ާ.H���@�]<��;�e�ݸ ̨Q����l%�࣏��K;D�C�U�,�ӕKLT&�kϲ��4�.�2D�ǹ�!�w�N������9�{� �~�KM\r��m��
�`���Ed�}�SB��H�V�eY��,Y�y]�#SY�x����܎�m�I"�샽�oum���\��A��g���������]���:�u�Mwv-�\+FI4ݦ]U��)H�P���a�H�����	n`�$:��ha�����І
gh��II'S�������%]��H�����QP��e1�>�6n3|;>oF���]���HDc�!B,��2�LD�,��-j��e���[ Z�S��S	H���[-�
B�e2��$��������[L%%�)�����7�k��<w:ƨ�nt�sX�B�H��DDDD�o���R W���	�_]f=R�7(���:*�U</S|b]�\i�v�:ݳ��{�s#�&Rs���w'�$dnf�ڠ^0ڒ]�#;�u oݵ���Iߤʳf<섦�BL����%"s�����z]ە��i���|��~���d-�~�i.�ڿZ�>��nmEWX[����T�tSd嫴��@EQ���Gr�G��U�UDEշ7�r���u��i�Uþ9�-�ro2 �ވ�9Meq���MHlt�	j�{U�݇�f�����^y:��n	C�D:�b[���ӕ�^ 2����4��뾨������2�y�e<�Ҁ1w#ePr�G��r�V	�֥Ϩd��,��k�(A.U�y%=�W��bR_^����<8Iǹ��:fI��	P*rdu�>=;>�����^������po���>޽��^L�:JxI{s|�Ľ׊c[麞�u�Z��)U��W-��<J9�5����a�x[���,�׷����츒R%�#&9v*�P�'Yk�v<z�rG0xC�܃�*:�QI��.9^��£��qC9��z�Z��f�On���hu���àF޹/rt��@���|���U_}UC������R��5��F������Ս�R}К�e��p[���f��@�U��}��ށ�T��4t]�7*r2� `�9��xeW40��
�|1$s��k�J�S�՝ VĠ�g��Mt_��"�	�VNm7��:�P'���r1�Q��>.׏�3�A���� h�.�Eα8�O ];e*�!b<u/}�G���r}�7ډcY�X�$���=�{p���K5|n\��G	�����/�KY=��F���ܣF�f+���,�����;�΋�d�s1 +��嗈����u�_���W���f�^U蜅J~jw��!k���{��5R���nGvy�p8�r�q��j{�;��Lj��.hf'r,�REM�\�͞�H��@H�>���"q��:Tf���J�ت��wu��ڄj�J9�^��MIh@�h:a
�y��S��/�����$c�Gה�u߻������j��ZE�x����t<1[η^:'i�,��ŕEtY��+�737�;� ����㽇j)����z��pߨś֓�����	�,"����_v^�訋�_�w�C��{V�S��x��/�D}}7m�1����61W��6bM�0���u�PЖ����{�����M�b��x���Ξ��cn��J�|�3�G����x����k��*�0{�Q�~��a6r�ey�1Uןd�ٞ��7�ēiߛը!��Q4a��=hQ��G�g��a��M�h���[�ӊT��8
b�mp��e��B�^�>���m�/G�����=�yCoҹ�F_i���=[��=.I��q%�6C���sk���=Γ{��&�oPT9��-<�%�&�;ŔT�A�O��(Һ�ׅ��8���F�X9r���Q�������A�;PY.{b	�xm����-��7���e}��4���;-V�ٔ�qު3�V����Ds.țc����O�+�Po�a��z�{���u_�we>��L�DQo�*����� �躴��e�nܚ�<��ma��vF�MƻuAK���W��1��M�<\Vp܌�v��[�r�bּ-4��e}<љ��<�����7xB�wmU������w�<*�.a��Z<�΋m�Rv�/ ���h�:�G%��#2۞���bυ�~R{�_=�1�������m�r��5ͿNy0�',�c�y3uK���Z��Y]����^�5�16�f𸴇�k%�F$����BI*�R��G"M��Q쳥��Z�ټ�{��V��;{�� ��ź���գ}���tDs#�x��ד2�wfJ�m��HP�����ESgdp��n�3`V�PT�S�F�'	��sǲ�It]Y����1(��[��!CE��b(88��Y$֎d�V 4kn3ʝ5��͊��gx+yCZ-�1h�'a���m�\�ּ=x�H:
zl�=M�]U4m��]��Y���`�>�gv.��oRzN_$�F�*,����v�y*_�&�J=\�[�
u5��3Eot˰�Go��t�B:��;��zx]V���<��GȞ���+X����]q��'���N����ܯ���e*)��6��T�׼WGmu����c��U�Y��Y�*]J�ī�R"��N�J��
%��ַ�򕁃Z:� &�@X��Pj�G�ܠTt�E����֛����\���	Ii�<�1hJJ����G�p�'O7�%1R���ϡ��#��ApU�P��YpU"�-(TR"��]ܴR�����R�U���鴶UU�Q����.��*��uM-T�m�\��)������EF�(�j�R�T5R�
U5J�R""Dm��*�JhU;u���G����'��m�V�3���G�|��C������Zk�̯\u���M��	��m�۬�+�7n��*�N��%�i6�{|�˙¦r;�mD�5^����p�Ԗ������ދrI��7�q�9a�k��2��\N�ʡp��9O�l1�N�R�YO��ϝu��1V�w`}�������(�����G�f�����
Aq+}��}V��y��^���tu}����_$ȇ=�ɪ�37yp|U+��F����!�[����π��ԧ�^yj�r���3�+��Gَ\����
�;2瞚ޞ��Qgu��K����L��wtE+�¼�^z�\��N�>]μ�~��	7�����z"\����<UqD���6���2[]X+�����Éa%{�>��۪�b}6�'"�*�_)<4|&�j�.�Y"5������e�Vy0ZM:�awl�j�N����Ww40�<�e��k���|'����BoE�ՎȭL�[;l�ED�]$7�����޸X��ۈo��!k��+�A�q�7�=Q��_]Q�w��N�)���_@T7�*$�&�lҼ㣹z#�a��u�ehb 5�+�MkZ��I�LE�C�y�����O���2�^�\ʫ�����F���O�*.�8�_ڕ������P�E�{�68�utM���t�y@��\6#��x�Z�D��{{n���^��23��rχ����]�W �� rx�|.����v��rn��w�[��K�¹���J��}um���ȵ���fu>\=�Ҡ�o�%X�$I��8;����qFBv�ƍ/\w�CPG<g�P�]������P�|3j�TVQ���Ѱl)f��g��#�¨���+J�WZ{*e�`�NM-�[G��g��0�љT[��JD�Ր�'VR��X�J��MX�p��d�v�DA��hS(z4�"B+��}L7>����+X�F��|2.tKqk��u�]���^��!��,�w�z��PgF�Һ���>��Qi7�%k�Dl^�`��U���2��Qtҷ��ǜڞ*I3^��?tl�HFI/�<}|��>K_�9/�Q\+j���w�\T�蛌2�<80
ۆ�ނR��{�h.������X���ϲB$y��%��lWU��0W������%ʣ}lW���e���Y�m��dN�V� =���3FjK�<G�r�%!���%�+���N��Ti���Pԉ0����%������4\i�nE�,�A@g�/=�Z2nw��5�p�}k:��d-��]υۭÄ%&���vޕ%Gbİ���D}tח�FA�3�ja�Ւ����B�ޢ�VvUO��ܙ���{�c��au�R��`��ْ1����!��=٪�y��л#k}����RO��1D��R���<���m�a��^�[�O�b����%�e��V��wEl9������k3�eUX:E%�Ǚ���
j�o$}Y�j�LgA��3Al�`�
>�>��{ދ���O��nz�|��xڝ��:���'�[�b6�Mʇ%�+�c����4�p���	����Q���P��j���KJ�uW��J�=JY��u=c�v'EA���x=V��Vr���2�y�k�9��� ��9'�t���j]��Ҥ�h����1�'OT[-alJ��T,n�9�7�i�/�D}�շ>rC���{��;��y �R��agl\�,0�i����N�S��T�v'˷�v-�&Ѐ�zk���v��(SC��9�+5�h��;G7�o��"8��:QeC<���ӱ�)�/Ñ1ts�2"].ŏsXy���Q���=��r}���0�U��ot�ҵfrj
�v�e���D-�mѮ��
.�Mѝ�;7:�Uf�����L���/%��FD���B��n��v�p����"ҋwۗ�����u���DZ�m�6�Ñj��Ӣv�Ĭ��JJ\�;�^YE�c\{;�H7��*���]�7E=2��/��e5l�<�e��5kO ]��s/�;��]%���@��H`�'��m���T�������lԠ%ɡ˺��@������xSCwP<ӛ��Dr} ˮ������r�P��M.K;����/:��t�8���v;�k]�R�Mƥ)��oVQ�ʙ�-擋�T��e�)�"�W�x�h3V\F���*�OTғ��_K�� �-l�CI������o��_YR�����y@G=+͞sֵ�0`8bnq�仧�}��R�\e%;�)Yx-r4"̠e*��N�9Ӽ�{��k�
�DJj ����U�7H�Hl������R�i��E4�)�EZe0��%����#R�i�USE%%K�X(�҉TSUER���ET(`���h�)`�IT�WE\����(RP��BTU4��S*�V��Z�������K�R��)��dX�E�)�	$�ɶS`@$R$��_���^_z�R?���7��]g�$9�ӿ�UVy�~Q�����w/_���N�{��-l�U��L]��hW2����y40A�x.0�������V�b�9)�K3U�X�ՒkoGq��*%̊*�Q�%gZ�f��n,�gD�]��X��+mJ�W;�@e�F�������F[�+O<%<ƻ�Dkt�]c�jT��T�3���F������Eww���g"�+���,L]�G�"]��Y�s�x7�<Q���R���J��r&�th�Y�}��ݨ�C+�q]���ԦP�����YOT���:[*���;��Ԭ��I�J�A�>�Nm�MѺ�I�I�4g�*�s43���M�z�5��f��n��5��Яv78�GX���"�v�#=s�;�=j�L�+��f�z����j�&yf'{�yS��fOH�N�y� �Զ�k��۹�i٫���^�ƪ��v��	�y�[�n*�g�ʋ��մ\�K/�u������_lV�{Wf�V�I�nH��-�Q��?m�{�jD�)��\C����mm,��c���������0d��(�"G�G��������#5W�&;yY=q!pp+���%.T�����<��n��@/��[Is�+��L)yZ�tȟ)�Z�õ'��=˓;,Wf�bڸK����*\���ev�n�,��\�eZی�6��nڋ�[E�5jع�i;o,
�|��i��S��X�lU�L*(N��(�FgnңU<��K�}���շ;�혤.9 ,t,�4����v�j��K��8�Ga;r��� �),�n4{��hG�}���.s��X�˦`�v��,�)T9�w��_U�Em��/���v �/'�*4�]�����O
 ������uL���px3zgף����B췜��n�ő��s��D�a����Ѹ�e���8�">�"�%G�s�ڇ��^�n��r���r���D�͑�I:�؛��y\�x�P����ajG@�h���q�P��V����-����<�ֽ�7+���u����Û�y��ۮ{l���:ȕD�l��<�"��� �{���fV���%RQ�MbN��<�gY�;v`�r�=m��r��}}}�ۧ�*�`�m�v�d(��U���C:(�v�u;��r�������ʩ�'u��Lc
��I�srRb3�|J�R�/^{�n,,�dh��s�9W��r��W�x	���ptn�oCU1S:D[=�${h��(d����P@�����Y}~�I��Y���󒽎���P��ټ�ʤ��(�$������v��2=ӳ��L�ή���E��M�ͥy�����ĺC�]M52��V=S�u~/�K�}�7;3����Ă��tu�8�a�u���r��2�����<��g��ۥo鬨D�Ιx���Z]��b��?TՒ�F�Q���=św�2�^>yڛp2��P�\w�[��ܛ�;hN!>�Xme{ΎTK�l=ӛ3�b�֌R�l��=W�u'⣮���嬮��ۗ���YRz�1���$�`k�9ؐ���ǦtҾgy=��E'ϻs�,���,�<�[a�-4��\v5ڨf����ekN�TX�m�r����p3*�+¬:Ğ��G5��d+��QD��+�v�O����4�uӶa=�!�a{����\��f]�e|���Z�\���ήv�!��N�U�ia��~���m1��"]�ï_�u祂�1�$��G�����XȬ(��n/��0&z���I�\�K�߅qxo����'�w�;QU��o]5�>��]�͜�m�a����R�TH��3wh��i��Θ�z~��B�ȼ�_B�:îv�⛌��R�弫ˆkf���6�t2�x	q�ؑ�����B�[cr�Ug#�s�WQ�|*廼��?\ ���d�n?��Ꞹ��N�WQ=/|���FBfxd��=�V��;x���M7�����)K6N��!鮾y��e(� �E��2����7��[
p�,�J�ы���X�[xkuz�i4�xsF@�@r�+;u��'ձtV��u�>/C7O\�����ē�f���	C�}9-QVڮ�6=�o]��˹���p��	�<r�쑛��o�;�86V5��f	G���c��`�<�_;�����j�٤�;$�K��9�������h�uV�8��^�����Wt�jwqI[�%eZ��R*f���Z����X�8淎��9�ȴ<�j"�S*�h�4P�BP�
�SD�*��*1*���Kav�L�mڔЕu
-�TQJʪ����Q���K)����[Z���B�C�R�D���U4����%U,*��)LP�4˫n
P�EWumT���jPUUSR�YT�]ݵM7t�*ۅ4�B7U(�ڲ�*Ү˖�Q*�����.�TU7JU�uM�˫��w'R{ǥ����Q#��Ss���7�J�Ɏ��t��&�Q�~��W1'-��vI�b����<�3Q���`�a^����aqz�Ӻ�o�	5Q�:7���'��U��8���dyL�g�r\it�t�(c�⒈�m������?k���^Xz�d�b�����n��Mzk5|�+��뫫�6����vق�#]�I�����}��|o���*A͐�3�%.���Ր���O�4�d9��}�ו�7)�+ ֽ�
x��h�U��q���j��ܑq�=�� Yш" ]��y�ȇ��<a�@��y�Y�A x֡� v�`Å�c��)���A�|ȬD���a��A�oX����|b�홑��mW'H��r����3M�v�����n���Wq�GH�!G��G�&���i�_g��{�Y��F�x�Τ3���0Þ�)���o�?ы5w:�+��í�ЛO�12����	�OXDYh�?.�ڥ��8����"���������`�$At���</����霯.�>#Tc�ܬf�i&b[;�w9������Q���iM�s�2������>x�]&Nкz�5�P�Ӝ�:-9�)��v�*��0�qG�OP!R����R�n�f�Gw��X�Kv��v���Ö.���]�;x�w;�3�e�DC5Y��_g�9�-`<�� DJ�3��fsE:L��j��fӞ�b�9p�:O�G���H#1��bK���^��}�ގ��l�z���c��aه��˖86����GLi�^B�Y��μ�qao�#W�#d�JA�F�9��{��_(��"�F�ha�Pȧ���m�:����g��0�d"1*��v���	����Ԇb�(�G�G*�|�{��хГR6����n�ɖ"�Z��V�6?d��s�P���ٛͮ�Q���Ĝ<E��,���?^O{6E�H ��:l�C���t��rs9�3):���X�����u�[�8�Q�0ԙ��[���������{N�o7���4@Z�:�7X�k��(��8�:�����NӚku��_(˴߮��Wl�u�dz�����gb{�CK#O�p����+yx�ӧ��(�)/���?V�~�t��:G�٫� �=�!J9|=^�~�;��Hi���2�ĺ(�3fX���bh��v(�l��.s���RTn,K	K%%VeLQrꢧ�0�B��n��e��ǎ�r���QEי�I�r�b�]]��=��a�<ş��FOٝdM����0���jYW̞�Y; ��;?9��\����Q�N��׸q��-�W��
��u+����7�i�l����0ؚ��~ϯ�#������g�����^fn<9�\���\m)��`t�L��k��6��@�,�ƫ�]a�""`�۽��S���a��b��I:&}*�<���j�с�G���+�tb���x���Xl��g��	P�<�e��&���Q�N5AF�׻���`�,���i��r�������֎�N���KLf�)�W�o5�V�\�F�o�Iz�)�N�6��o��q{���e�u5���s�3���{��vu�ݰ�Q�ßQ������7�꺛E�Љ�ґV��6"}Ay^�JB9��D?Y����6J��Ώ.6~f���?ݢ�2��6���W��7/�UY�T��볂l�����s�ĠM�Jt� �pH˒���C{fb]B�j LJKg����i1�S~��yJkܲ� ��=O���/P&ʋI/�Y��5�H�2]Ӫ��ۼ��Fq�QY�CO�>8wA��7��P�A����!�����'3�j��@�a�@x�C�{U�����y^��Govu9�6�t#�°Þ<�V��>Mg�M�3{����Cɶ�rٸ�k�!�{������^�γ]�'Cɛ�hQ����7^f���R�<oJ��5)�2�_V��S��V���t����sQ|B*R
ȘُD����˘�1DSP��E�X������R�T�Zs7F9�˽��GqZ����Sl�_��;}(��^!��Z�ㅑv�� ��b��z�t��ظ�/���cA)V�Z�W���M���m�F�S�i�c8�=���Ì)2���(���̅ۉ���?e���x�t�˕�ߜ�(�T�y�6�8m�cW����݆��}u._���]m�Rʺ��)�۸6��N�Ԃ�܌�%]��oJ``�����Q���+�P��}Ae^�����2�o��Z�tX�Q[��M9x��a��Å�Y��[3>�f���-}D]7�ƍ��p��^0�dx���a��ö��ƾ���B=b�!�5G��5��ǜ�o�tv����������-����|~g���5~��)��R:+W�V��m��8�|�q��(�
�q�m�N��8�C^�ڥ<�c��n�Ϩ[����&3T�>���i���zc��o�h�Ȗ�L�f��L���9;��\�.��b�*���O4j�ۙgv|:�L�I*N���,,�i墙Me.���m��mz��t.�V��sͷX]�����+� ��
�Pz�p7�N0t7ݴXU�5���x��ɚR)��J�ţ�,�`�-�)%�^gj��y��ܩC�V����oot&�ŷO;�\��bᔟcl�Xz�+jL{6��ݖ��P��Z-��&U��a�/[��M,M�%b}�h4�i��鷳��G����Kq.8�Td�J�ۗ� *>�Pw#C�6��m�H��םiF!v�.Ɍ��N���Vөs#�F�^K������!�
�OqZ X?O����W�ȕ�5*{U��2YM��ԭ��^b�|�Y�X�����]M)x+��\e��r�2�7Y���M��Gn�Ø�k4 BNu�<����;�qK���R��m�#�ILЬ�j�cI��
�E���������A��mI�(&i2�L"��CA �h��"��ō]�)E�t]�M�j�5WMRR��EX�t]�Up���V]ĻJ*���.�j�n�����T�*�(e[ut]��JT���lh���R��T[E���2�X(�,j�Q��T� D��E�?V-���^��W���T���ŉg�RW�a
S�UqFc&.�@���t�%��vF����4�����C(�ֶ�3V��X��?�x��O����(�D4]uL�|�a �0��}U�v��+Z�O3Bq�{U�s��oSj��9��a��fyFyZoUn�=]���Q6GHh���m}rg}»��jm<�4�ʖ��(S��Q�޽=��i>� ���P?q���L���/f���#�]���5hdB��U]����vo��I�a5����=n�����;X��R�H�	��5�+R��� "(��\C�Q���u{����}g� Q��"��^�纔&ǐ�~���D�:��3hMn��~�@�N��b�6�a����K���gSح'
ݗ��+�-0�=�l��]�L��q3��D���x�t}��	�a��U�iN���n�Ӭ������܅��M}�a�G<�>�Q�{��Pۄ�cծ��W�g5���<9e24�8�v��Q;X.���	U=���]��n��Z��n�X���6R��c��3�o����k�l���i�zͱg�Ֆ���vSG��\��.����1�"�����u
"��!�ƈV����w��w{�Re6<�K�Pq3�<�����wJ��(�>�� ���:C|�]�����M��?d_Q
V��ɷI�QnGɟQ�	q�uS5�-�v0����|��ya�3̋K��|�Z�ϡ�6~�Vt%��f���X%z��x��HG�<F�e�a�/�g9W�U���fn�*D����^�Ӯ �6^��ؒ�f����PJr`uT��ӷ���F��a�#�d E�o��޷����>�<L�a���W�x��럻����w��1nw��C�5[��ޯ���B.�O_�^���BΤ�c�"��B��t�"�5���W����Qx�s���?+;��֯t�c�)�g�\r�1w0�p���v⿯�,��"�޴,�
\W!�ޡ��۔r�r�yC���Hg�F��+*�o>毽4n����^�F�ZS�)�~̀�9}#�Y��	�7�U� ���4�̌��q�W���/y�+����{�z8�g־�r��nc~��3�i�2�t�	�&��j��8rs^(�6^��u�'#ƚ|�0�&P�h�wd�F�t侞C���|!��e%gH����VG�#��#-iR����ܹ�7ǂo59Ҹ�v�t����~K���>;�I��↝?/~w�cө�o(ߨӺ������o6��?P"�!e�?P�=:x����M�|��r�"
��P�f����̮�ՙ:���������hgl[�`���WøNQJ��X�:�U�;f���5Tr�g�F�/�k:5�q�����R�
�	�k��g����+Ʉ���w�.Q�-���׹�sn^�����9Lr�\��&\���޲��<E�x�3���F]<�w>�U�K�N��i3tb���r���۲�~��:�-��e�+tg��޽�Y���8�|��-ӧl����aƱ�9��Խ���(��Pe����J�����)-9�ڕ���ܬ$3PF�[s/�Uz���t�^���t���Y�'wV�m����q[u³L퓻C����4�V�I�-O���[������L0���S8��g9�)
>:x�r��8�"r�LwV/Nw��`��P<� ИS�����?k��*���1��K�(�3�<���w�6a���c���bH&3'r�#�+G���2���V�����ݛz�|���i�P�f��h��ݼ��u6��oɖwu1�)����s�6i�oնeXe<�F����^�e?C���w��<�G'a���*ݐ�Mc׶gZ�a�+�R�8bKj��Gw%5IM�ui�q���Sb�?q�X\�Uw<����CH����<:p�!��dZ�r��`��ʎ���	:w�f���<�]���V�Q��@�h�C��͇��9�����Cu
?a��u-0�/��/{����YN;x&Y�:h�*.�5[�8��]|�X��!���l�k;��ѱ���fɇιFݲ^1���j:�i����Q�)�]�g�&�͜�l�c���(�A�(��s�C�`�Ko�x��c�*i�nWKFX��۬�3A5τNiL�Rƒ�K��bNΝ�_w/���x��g�P0�K�*�����o.���n��us(�l�Ŏ�uZhn�:~�FD' �?	?5o5v�������L65��H&�J��ξ��#H�
_*P��o����}r���A?6~hд8���i�z�x�h֪[��̰p�5FP�z�V��j�庄���=b��У�(�C)+)n]_T����Ogh�Ĵ�锘N���o=޳<���q�gշ�34�3��}~ڟ2w��W�U���1�1�t����*��.�2�	�9���k[�_;ٖxt�4s�7ƍ�x����i�],�d:E��� ��!�Y����U���CO���⾲��@�����G�j�*�8�ڀ���qg�z����� oڙ�* H0�?tB�>�W��:��oTy+u-1�PߵHs��H�n&-��V ����`��V�ȹ��?t�Ø�,T���Ld�Vz�A���������Y^t��j��j~X���(�A�[�/me�s;Ղ��Wj�i���s��Q�S�U��d�������{@�(��Z͵i姽,5F�6�z�X�i�ҀLAF�,˻����ے�۩i�Κ'=|U7����U���eqk�.�|�ѻ��'�<�A֫����vt:җ��A�Gl�9oj^����U����;Ņ#�v�f,�]pKe޸����v��7X�*�Wu��
݇�"�t�u)Ʌ@��̣ٷYs��	��Q��t�Tz�m��}P�ˣ{�F^�:����f�u�DvU*���X�����UE�n.5ʙwJ���U��W�]��Wie��d�����f��scRWG���vmY�|�ɯ�����WKe^m\��=�MwZk�Ęi췊��C�2MұV�V�p�Ъ����IkZ�i���Qo��Zi���y@D�m����(�R)qHrH.&��$U��y$��ر];Q}Ȥ&���T���l��ф�H$�%*TX"�IMQK����H�,P�T���H�B���Km"�-�Ȳ�#T#V,	BSA`(AJJAi!L��>'����\k�����uUQ���^�n��H�m)11�S"~�����W�`����S�l`�`���@C~Xl�T���kN����6���]�qQ���Pi�D�p��؆���]"F�z��#9E9�w����6�:v�]&uB��N��V�v���(KM�uۇ.��V+��{'\4�Ӵ﨡�e'�'�%���ݼ+mih�� ��t@y�f�.��s�g�A�f�o��i�Q���P��W��D��QF��wF<cO�1�=���܊��Ko�`�Ω��U��Il���d�w
��1��NKGs����N��ӷG��QQ�d3��e���i.����W2ͧ1[m�5���hP�g��<5�rM%괘g�S�N�.����}þ��&�3
��4��N�u��.�fc�<Gb�x�E~��{p�~� �yq/���Z��C1}2�͖�д���?uQz�B�᤼|Fj���w*�$��D4����}���㺄v�?YQ���V���Q���%��M3&�a�׎�vY�]X�Xh��b�Em�2��#=��=����u2�v�et=$��J��?iw�p��_���%0�w�����v�s.��u�q�}������Z_
�h����H�MT���0��&Ɠɗ�9G]��ǹ���\�:C��-�Y���]P^sX�����mp�據��}��ףΓo3.�' �"��!ف���C����a�pÄA���+J�-����x�!��5��t���1g/�JN�ׯ� ��4~
*<Eb��^��Oʅ;{��w�ʺ8M��R�y������bu��7��k��w�wr�ϼ��o�,p�F�<�,�H��m�bǣ$q��X��v����"�w����!	!��=��gHߩ}e���)�a�������E��M$ӃU��Z�	��m�(�Nܭ���!������[<A6��t]v;�L�0�E:!����;�P.�y�v��� :����VAY(�#�90��½�=Ooƫ}s�[������U֊U�5���x��8k�������
��B&��Gx���1�����;�CP���0=�����>H��Y7�d�w�)���k9�9۞���"؛R���}��0�^+�=/�\����pؽ��Z$,Yuo��ti��U���>WJ-jw�$��yM�<Ҫ^��
�����tuݑ����{�x34�
.��窽�o�W�b���Va�d���Q�S���%�goJ*��p��\��p�z�\b��c�|�8�}���qT����@����� t|P*��g_�j�]��f��f�T��u#p:�fv.�c^�t����}-T��C<�אە;i/#嫰���,r�eM���
cs9i�lnx�����n?b.���wɜ�VP*϶��C1��y�HR�u�^4w�C�Т8%̎�G��F.!+��`�v\�r�T��qs��"t�[���ٺ&��Q*Ds�aY5��vGm�<���=j:����~�q� 숩>�]�������X.�'�e�.�+)X�D���Ť�����lZ��cZuM�2�;U޻�qS��.v�,���iH���R[hT��w�Ve���PD�˳��]';o�my�׽d ���ӚF�)�W6	H�*I=2��U�r�3_���QDu!��݅�M�ڮ�O�1չa	X��:ވ���[Rj�tc=,���^蓩";(�{�]F�[�]��YFt�uOr���-��U�a�7��6,�{5+Vk��͏y�I�i��xN�h]�g	��4���:������%��Ñs+�~��:ϧ�n��x'�<X��=�L�<�ƌ�/ťp�#��f�*Td:��=�^�BK��R�7�!�+�ٞ���*�ZG-�CZ��9*�FL�[��9}���b,89W>�%�;_\ϼ��e}�h��=��~`k��Yz&�/u�и^�eM|�p���l��3X�B�H���q�གྷ�����J����Y�Fjl�:���b�[�٧�ֵ�Q]gf�\�Yi�RJ�H�n�Tei�fm��]�$�4K|qT0&��v�v^tu�@�;���~�W:�����3q�S�4���`�p��&
�yF��^��5�������ܚ
TU��[�r�s>�Z�<����z8�a�BC��S��j�C�wIm�]�����=0iݽ�2Uk8�C�c��v�^���٭�d�!T�R��1i�z��w����57�~�x�۩���qf]������ޤUe,��;8�٫XƂ�e�|�0#�4�Ҭ�Ç
�/cO�i��D��+����JsS��Si!���G�Ty.�*��cbSw#	׹έ�Et�kȦ�!�JT/M�r'b��;}������B�	�٘�.��no�_��-�Q�����վ&�j���wSj��3m�L��<3@鎦{s�y��e��H��Xv��u�L�B��-��g8f4��;YG�A��u�5X��g:�B�X��u�.��YJ��i���==�����L��-9�r�Af�M�y#"�I%@�R\��vV"���c�նB��]ǘڄ�R��{�{�|,��E 2���JHRj�%$P��YQQ�Qb�-U �X*))
cU<�M�SiRB�E���
*� Y
I��bȤ�I��5�{�3����8�q���#��ZF�J���>=n��=��F�[&����4�k��R6�q���d�,���3�c=��^��#̙KY����Q�����Y�U��F�bl��}�X��(��^W1��.T��H���52�_9Ӭn�J��'���j�8u���Iq,��W�۬{�3�c������]-6��h)4��9|QSi*�z���� LAw_!m�SF�3p�E�l�f,�Ʈ�A���7ےx�v3����Ѳ dm���%��xc˛0�aM�����=7�Ǝ�5{�<�!���;W�CyK�X|��\ ʕz�x�ev`^�}iZ��P�����>�� ���C����xpB�e�/"�G��+���.�	�ʳ5g�4x�p5ue�����/���h\��r�u�2�t���������U��ˑ
z�]��.���'������	��y�;��F�i��Ħ���+�Ƭ�e�ѝ��u����/�y`�x=z��y*uxVq[�/�"%��G�x�EvZ�vY�ui)�a�RgX.�+x�^��'��Tu��b�սײ ���mZ��K��i�E�k�����-L�f�45��k�t��m��v;q�̽-��XU����g���aV£W�#�d���>����.��:�<��%:�v�EvV�S�ga�����;fx a�VK\��tԫ�l�� �ߚ���/$9���x�����c�R�L�@H�ĭX8s'N�G&Z����`�<�kTz�=����`�uU�6�o��ڙ�෗h��U��9�o-_D/y�'�Fn�e
�u���w���e�]��yH�q�nB��#i<۵I7Q׋)N�a�-������b��K���V�L:�ԱyJk;qTg�8�R��hN��:ˏ�o�/;��w�����Fo��
׼+Mכ}�P�z�db��@o%O���Ug�ʠ1�űZ��e�u������U�0�V���dL<Vgrxs�V���Wփыt�7}�C��W�^��Xz�i�UZ�ez��|��I�a��\P8/Hu�#�!X=u*��fު˱ɩ&�]8�	P��ᵕ�uڀ\��4��
�*'�;��p�˽+�s��(j�=��2���X�V.n��k�}��{H{;���c�J�ݿ��jvH�r��m�Hs���߼�7������W��ε��j�u��xְ��u�W����{�[%�b��89E;������'di�$W�����zB�}�\EZ1�@���ڹ¥s���'gf��k�C�L�����&p����g-�Y0�X:ڛMa�Z��Y�p&1bo]*޸�]�9m¶;�:�����V���>�o��=X�Wg\�X�o_�*��/�[��;��}�Ojm�8�t���E�����8�m&�x�|��v�D�^ ����:Q#>�xk���'ݳtf�����V �$rUj�kXnOH���âE󝆲wJލ�9ԑ�0�:��"3�w7+V6v5t_��nD^�Ч�p��k���fW���IE��R��D6�L�[M"Q7�sl8S��9���A�,�f�;q�##(i�GU� �.إS���x���i�p���ܼ�Ԇ����%B���{�5@5�hN!*PG=ʺ���D�9���l�䅐�h��<����W����s�?���^qY�X4�j�T6nw��Nہ��j0�&y���,�2���>���&{��m���[sH�M��w2C��[Kٵ|�w�xƳ�;�Ѵ��?����?�?W��*�EUU�5�~��H���T� HH?�A�J݅�R���������|�qd�ʭ��B��j�!P��Š�9�I]���}l HH�A~��u��ڿ������r|������5������Cr�����ٽc��w��>�$pt>x��vc}����Y=��~���?�!A��HH�:B�a��aRY����p~�~j���̟�K�}z�����g�2����$		������O�@��^�p�`O����r�����L��O��@?�
��z�}�q?o��Wu���l2k�?����		���.�����B@�z�\!�p�	ܒ�+?J���-��~�$�x?�������&����$�'�}e�'�\?gڋ>���!�|����O��&p~��G����-����~pe���#9Q�O�~�}5�9?����}Td�����S��(4I��?���}��������?���g�O������ϰ�0�! }p��A�����������,�	��""Є�����$		�����D�����AR}�:~��8fB}F`_U�B@���Z���\�C��G	�;�I! 1�5&M��~i���ӤL�J��H�d�5�?X2�P�0g�����d�! x��?y�~� ~h}��! c�G��@B?d���>���o�������O�����Id'��l������/�?�柗�����?i�B��������@��>��1��rq	�d?T HH����g�e�����s�_���	������ܙ�i���ƌD,�����$���;��u��u��O��Y�59���1��aB@�ϴ���g�����~�É�nR}]����A�g��}�i�Ē��!����$!! �I?���,�� }��?��o�~QHH��q����4���?
&�9I�&wu?Ec$������@�~�G���H�
Ǜ 